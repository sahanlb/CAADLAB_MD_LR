-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1uw90AGQJfUCdS0bHrwaI3vPmgKquOEVltTRU2P9na9DUeeT9BRzDKeqSz1g4hS5
b9mEZMR5KFIiWoFwM5CL3+ArqBFeI1EoR6v+Rebl+cL2oRJ0+MYyCWA/HiMnrtWR
ARifPU1XIaI/IA6ll0e0uHBUKBZ6gGRB5zWFSvw2TgE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7712)
`protect data_block
7YuT/EdLscFyKkzkxrzf0138+rSTd3/lWSezAalh+Qg5scKdfJCLlFL7UApf0YAr
WN6AYyXSbgSQxl7J/SdwXz4KpIIrJhY1Rc8/m0JLkhw+NKX2WIGXNxDlvEnq7ty7
BwOivfw934pSIiEAhg7B1M7RFxC47YBbPFG+NzhjDnwcSEl+KJKPlpKkGtbJ2o2m
NEfuYmpu84G1DAHhVM+40/iAm0IpzFVDhXVtNE1hQ1EN1Sq18tCdMi705Pt2cwGO
KXC6NfY3e0mhQjieA24p9eNGgH0cTl9FnKmSoCeBHZFubtSMXT7+0bTGZ4KmxSNB
bSJRXnyYADxM2Yt6DdgY7IOkJtvakJuoXO8arMBLzJqci8rSCvLcy1kqhXsF8+6I
1lwMplJ7aQLwpnMxFONRvbRAIuTImXIJAq+hcDkiFUgciy88cAHX6svkJjo+CCzl
Q82sFeApApru05kMxaXct/mlmE7DAoGs4WN/85mgg4wwlbVCbGkgaIbXnF73mn5r
3uqhq8jVuqRFDq5LaT0E2nydLWK4AmOCDo90OeM7lliOkv2e6vVyaFDUak1EWQvP
sFcn4nq8q2OLc0YzgTYgRfbNeQp3BfQHptv4IYeKxZho62l0/8OUmxbtI1NvJNki
KnyoUxQ8YKvMXeS8rPv34GLUaTjNEx6Kla2l4FtuVhA/Q1QXOlTVFSMJKF0akEQt
UbbKEl7Ini0Kh3mh4Jt8HqUxDCEvvq9RuvMBFi2zTL3b0hClazdQjmR1bIYGRome
ucNn6wmmhswdFmoWqFPidKKXNql9TYC7ObFGdjM9gZGOHmGp7SRmuqrXsHTCN+0a
rmTfTGeMMcFhlobV2T/hn4puB7upYJjgX8ch/5dhCXXrstx+TrqMYncOv/zUNJdp
+wYx4SmZUIBVOgJA4boD+WwM5OeMC6i/uUpFxTvK1Q/I7muXAMjsLuMAucquxbeX
p9TCHk5GspR4GPbpYGrvzChjaSXCeRgkD9Hjw5TToTGiZIOtAIv1LsNnt4gruvvf
DGZQP3aLarnJRZfABJEw3EyKeovDIWToaRRgoJlQHKSMnYkyRXAcul/ixhqU470Y
StoSBIcrzVU+HK5C1Ju8yc4V/mO9Ib3ajyHP/xGW2Zk7hKPvkJ3f2GHQarNYQxpQ
dLv5CGZJMVRI1tALa4xxdNYZuoNUhc/jfZG9Bz57P+Owt6v2vzUnpvZOhokWzITU
WkMeYtFAXbH96RBRArH7LMvhzpv+QU56SkBYrR/djubebhQG03Gt2TPT1Fkl/ihi
cDIHe8Jvyj/6zpQn+ftnKq8pfM6GJvEZ0APIA8fVzOUALcMW0q2yXOXJrD4xytDU
dF63sEUZJ7el/ztr1DsyZ68gt451pWFRAS8S6tLTRcrOEIBXJ2rfshR4fiMWJq1Q
hXvMeNhGpRmXlM3cdbXXSkWcIc84ZbM8S6bfk0md1MHINDKNrsHprNNxNhgOCzZd
8hZYdmenCQ7UdjMN6y25vVcZHnIHEB3xqbDodhYvf8VRStZclLV/jrhfikr0sLiQ
fOAY3JSMsuaMEkQeqZSq8AB1iEmMxe/ybXBNS7pzyOBYmXKE6OBktACghKJvxLdQ
Wzhv0HKlrTId5twCGZg1nltbQCZD5V/22hvH/GYhtzg+FS9qBJGy5spS9vmioI3C
x15RC65u01QG9tRb3d50SJCFMgNs5Pxi5zmFnbLPzytWDHGlEG5tEABzYbLHgdWp
2SoABOABbBfmawqM7JmOb6zUqNMXY6MHCwlnZyMwl+SYy6Nx7zmgIr+kD+hRcwQ0
JDHzY8EvG4OThmHBkvO3pydB0jjPfSmIm/4QUylWnDWwER8KA5GMtedssANOsXGV
RqASYz9wu96fFBr0xH/AtU9O7gT/E6zz13/JshPjYqUD18brRiD48xXGKpA4Ffj0
kIiQTkwfxxhmjk/ciKRby5ZxAmrB7vTEHMcfRNNAN18BhZaIa6sT0YBcWzYdRlRi
hqshUGgs5TgfMVWaQZ8/2Cso94aIBUdZGhw/Ibv4DqfURKOI+PF+5HYFDLRzCw+S
y9eaGfdJr4CiZIP8rnoxBOV+3Ax7Lkuu9hghscBeqpvDGhTfJTc/KhQZ7zHEpJKb
UkDA0K5Kqxkj/+hpRXhkHW+zYhthdFtv0Xb6JLUc/U5ifx88UlTIJLgjF7LUKoVk
N5XfDW7BwWnV9NVxUu7men+QWXVv+ToFEFQuUlDxi6zZnc9prQgN6kXJl3kmg8fB
gfHjSLf8V2ZFu6pJwj87w32f9FIPCQAd+3tsZNAcJvSkSM6/B46zL7GX+MsXyUs1
Er7QnM5PzWrpKZiz36odgfm4XBeaO5lj14OePiJd9BOf2GSrLNIETUls+edlhpZG
H4+gxh9AXGa4V4eDg5nXhnHFtOXoh4pY4niNuWkCMNMydndlLyqovIRZ2Lmr5kKr
lf2O0nMiRAVGyRmP8i9LeQNRClJotVh4qNLkpkqBBiqOG5N6+JTED5mpb166yZcT
j3/QOYRHmIGS+i96CKrwAniFhvMZS40xUNifNoOmaHjYBKQjS0QavRS8xUB8Bkfv
fATEuJo7vP7Mm3ITdy4Gb28mILpW9xCA9iQUdbp5/igJwieKz1XOFQtNgqCu2lx4
PFAht2yrz7Rb3qUd4tUZnU6itwqf5RGTH5NGxk4dOV+/LuxtjVrvFCzyGxW6jpKa
shlyoXZnCCbGshMSUmXTyd96HMf/2BFFa2vJNBfDh+IOUuSNwPuquyAdOqVaP4UQ
zw+BxNSJHCh2W4x/SFMttCHwzwHeGNqTfLFLT0MUKCCJeX1Smo76F9rDNmnrrgwe
Ne0NMahqXFVhIB7bNP3gJd/BwhrgPe+QLdbOoH1RZfs8GtNmFUMwm9LFLa97y2rd
5RfQluiWs5fnpJYtFSmJKwuLsI5f+WMiNxc3wkAhs9wlqu9vPeG/hNaXzgDXej+d
17n9RHijqCGt1dYLr2/UgH0Ys+TlmBmUI/lgdzWO1dNSusaj57TabM3T4RK6Hsik
XFuETlsgLWds6TPCm0PlL0aggqeor+yDvlSNLoPP/brbj1Fq4bYgXx2TiFC1PHZx
E7zSydT0bKxUsCHcrGQN6tE/7jMs8eiW4NZtmp/aYUIUVtQYcZeb/sUWPj+D7wR8
wWzna8saQ/nvP9G2gxp9lswiWSo76RueABpHJm63wlhUqVFmp+Pf2PSr0ZqXIk6u
UaO7lCQha8kvrqTWAg19RstE8jz37JqJd2fx/jiz9FlC+pehBdSoB7N5yiy6LKO6
26972ipX6vUXal/0psZFrI246FIfTuYe4/QnRb5jZp6Y+FPklj8vn7NA+J/cVhGy
BFyc2vYwKsikUZFJbgNp75UuAciyR7K1W9k31+t9kEwWqALCG9xD7p2rAuRPwjjP
1F414Ht3xi/MKR1wY6prDyJEQXF4ZWQZ2zihWBejfXjPDF6e1vRQxdg9y0xFV6uZ
nT1Pve+WaTgIfQecUadFr98AsQfqyxIHYfj/gg9LKTalTTJxU5g9wh/4cqI/7ZXD
zizcC20oXSfyuYn5kjVXeHGOPlY+BKvzyQh8RkIGmCGYZlsP1oreM+qy3WGPZb3E
bMqQ21d0s77Es4/KM1CIaTSDb4q8lBEbZME+xlDG/YJ2A/oiXjgyPsmIFaaCmEgD
ijSPUe7qq5Z+Ws0aP+XBPWgym3j53JT3mTQFikbRWjtJmPpF5GC+3ssszFSEYsO0
RYPB7/qSNGIe5wPf7Y5TO3Hvou2rzqel6eRnNap9FlGOxE1WnUPGEHbLtMUDQIGP
I7ZKdkmvxVDo8w1NTofQUkcKO61763LtpKBErkH5tofdhlStJ1CvkpLpLWLhUJVg
0pe2dfUkVAukxeA/ql93NV8RktYTKAwitU3O/75oCYYq9GGhYnLRH8ucVYIpYLUT
DFzEKKOM+ulkFCE9i7o7FBA+DkDSrbV8ZSXKDLnHHUBdZdACRVs7S6SwUlPBeE2w
n1JFxyWKfXGqR69MeLTKE0QXiv2GHX3usq0HXq1pmTr8t5ItRYoqFQGBuR2CQoFz
c9njjnwMQ2C+mQqSJEtg2HrjUW/jSEWitXeLWWfkFRpRXa3obYhbQ252+5Req0Gf
XF2+0+eKKJLb2aCWlwf80boq8NjaKc7QIvGnK+RWdxRq/N44DRW/93ZZsEUMRETL
XetFn4UidJDNm0PmDptkjE3kzMN+nxWGh2i+Mhlv4sdHxCfueze8s+CIxbP8WHwD
xNiG9ex0HXSWMklWLDPxBVaOsQRc7ImsxsgZXBSsuz5bsUq5cxsr2cNJaz+7BnQW
3chOHlqWdcOWIG8snfzrSEhpeRnb4Tspi+SXIHLS1uGZyrJtN5maJ/8HDv8Do1Py
q5Bs8WUnoR2J5ud4BxODcQUyOZCXnsBqU12fTIXMfbuy/yGMthLGNa1w04RwNaRD
Fx4OM0ai15VwTVv+XvVLHNi8hW7f6iX0387AoRNeqGWDhzLTluOHNxzVusxtRStd
Ys2kzYoP4YyqGRwug7+pjmPx9tGxPSNX0g5qwl3CWQcNyS+G/6s/MhzwhZQYLpES
JXoLyXke/TL9C+ikNfV9dswYg7c1ajEQDAtNKPeTg2IdWrsTmiJOEdCCH5SpmUKT
kiyxvoM61mhL9KiPd0uFhJ4qDDD09Nx0BFZ7Wv4N6vAGtq3DLMm6nWyttGl97WXz
el62MhJEuWgmDUszUg8FGdZduhEHhp7p8LbWl2yomGhbRHbfhTU2GN6C/cFeSBat
bzqPXxnzpry6pgga4dK2qCNcshJ23f8GoSBlnqvOqP01SDhe15cUIYasMYlPMLbT
6csh2Tj11l9bjv0AV0QlXjPCbbEOt9GcuhHprAm7ceK/x52UBb+AQl5HCxUQtU35
DoB6P9pgQryuTuzZcBiERCZkJarevB5CietIAlQgub1TU/1U9DaxeUuwCYvI4b98
RoeJKi61GK/ZNzzuPhZqYWfWSa7/qnSdy8V9AZWV46VxJAqd315381ikhHnD52W1
vqADt01ZfhG0ncnKFKoNiZfu1KVwDehR3PxSSU9/8g35IVgeLTj8v1XcpFhyOp3I
NCjuc+lFbxCtV19jsZmAJaqPGgnhGRKJlC/1wDqdS1AT+TynDRkR1wPDYfY9OyLk
OQhY+NpZ/K6SADG7erJzO/UuPFpaeKRWC2xfMA8P9+d7R78J/clHmPuTZqZ34znJ
u67ojWWrPzT8I/5eUAF1MOX21QRHBf7/SsOu9N8DdXQrClTHhWRRwaBQcqgmvgYZ
g2PcyezWf786pxHc9gL2ybe5frOzg0bSfhAJumgcU4E+Swo6sjWXHmfpKFB/P1VJ
cq+ysl7Hu48pws33aYc71r/sWpC9xUTBAa+0EUmbePjiNZqo5e7NHsdWlI0UwVqb
jtXvaZBsUoQNHYns57vD3wsvzEhnbeaqoCezLYH4xdlCom30O/rgxLHPTjMaSbF/
Y1hFlAq9Z3OmqJBhMpUoflwUvQqYCt74eq1iiIwuO9c75h+2VtVv711uYP0FE5Gu
hiSu+94lHyFA6Vx4eHtKU8SSksPYuH0jPBlb7Y1o59dK8uoPbpWHuNNkunmJV9RZ
zDXE83o99lc8if/y6oZykTj8R2Fl6i+zkAhM+O1E5shFskUjCPR2a6qEhXnV8V2S
G6+TPXUoXJOjhWXMtyhbF1Nx3bJsscS2Vumdd0L+2vX2WNr7efm6lD1+ot3I+E45
Sz5gOFLzdxRn3J62MMLSYRM8t0cWIyOtSJ58b63P62zknrVZDhNIiYaCdSiyEwSN
VgHaOAKZIF8Gbbwc322BWDSQrztp8DPzRZNB6RPavxli/9yyNLfHxdqk7qVS/e+u
2ytkZdZfDjoe3LDhM6SNrjpgR/TBVQU1shqV/Pn4fdw8wc+dI3tnNZQ7EQIUyW/R
CnUpy3m7o3CHjtzmOSt5ZitqyKLos2Z6jhE8+ywHRqdHJ37HeMnx41lRCPjQ4KQB
lRHe4s47prsySgsG9maZV/lcE++Jhc/uBry82tNGqNE1fl8bpriWQX/axvt1CFMo
L0u023htzMOotb9myjjvM0uTFtCEYZgUHXUPf9ngqoob4VeZknxmtKywcrvneUVj
hu1T1n8AMs+euX9OiQ5dTU41QaH1QJKWavlI9gIpprX6iGnneAN+JEvPMbUWDmkR
6sMNPkD4NPCZxSq1+2Rqcir4ovNgFCt5dC8wOcq7hPvQDuFfmO9xSR22c3e8j9ZK
gWT0hFy14XoXWJ+GcrNlncfJ8cuAIARECcrk+XBoGQ0AJ3y5spCmqEsGVoygOBD+
6XdyAeNcUZV/JVsnBJhOxFWVbOvGsdbgK+2vGuhTOq0TwqAhw9wmyaeovuIVo5ec
Dmhm7O9l9uQjsoVyqkBaG8aI8mylDPwxMVvQnf6i190ToyLy++r6jva4WFbtVgjA
NSfPorYyOJuddfgF4tr7ufATLOtx+t9LTFWKEHpLB+SIDpZqsdXFPcB7AcY1hHpt
jrx5rtNuEmf75OsM0COR9WojWJG2UxgCLSV6ZhX5dS2tUnXbu/ytCi72dXsnpvLC
C1Yj9eK5DiSa1fD+G/Cf03wzLPLQjeIyEO2U4RqvXFi74NGc6lCcFBQaDXU03LNa
1uw1TOULhdJ5NV7u8Z7LrHGAZFcY9ZSsodKA7TZn8j0z98OVBKlqvVOmEWC5z56/
+HQd3NsFbwdUEKZgR/j3XFFbF519N2GwH6bSEREi4ixjOft2CcqA8VJaeJK8YpBk
oXgbBbClUiFkWw9MsZ93rTIXW1U4hkfb5LIGYr0OPbj1qb/TDmSyWXZsS5VVN2T/
CwSIEkBD9wxNr3qMVMV0AR358xOU6rWc9RFV+A/d0Ipzpd0Yitid3ULOPHSid+yX
doaU5MoAADeFvCg7zcGR3TsUsUwKGLbkYRsec+Rpmto7vlNLRR2Fqd8y2OXeAtoD
8eNr7lRC6gko+fvRxgsqPnZ06Yfhv0MWFnH8R4iYg6a7RLf67S5YR2btje7NJxhn
FWw/70hAStG4NG4WQ8ZmUC2PFy+KyacQbE+fQbbNDHgjdBRYCEUXqIpkIX7EBv/1
9QLP0flzu4y+NIkiUyNUOsqFFINefMuAnIaFnlxLeaqPI28tM2R5Xbz79/J5UH93
BT26W6koDvKlqOhtFV0zG17mkMYgvz1AioWNidQs6B+mciwcLxsrCU0qG0bY4S2u
u50cUgbXbpL6gWqQpjtr7E/k/aEdwqmDhA67WtH9nS4P2CgD+vyYwRHGKeGRqgre
LUpa3kwxDyUwc+yenzVmiv6hptGw5kqCHBGhIsmm+Mo8jCO3MJah5KfCALwEjIPZ
TLOii4Xbv6c6x0LiUvyF+39T9zr7HiiUvwLOe8SQaZUPXVpfYGkuairPaes11ow+
8F53dx7y4tRsiaZceYiZpU5/bfwjjfCjZ9cIc75aq9EQwrOeO0IFJfXsfHVr/9pL
Vlz9NKFvYAKnxBcItWu1ScLsc4qRJ18iUqBTuURnqSsRKJBAOMlt3QG7ts7CvoP5
SRKNsO8l/9Vu78Ypt9w5uXjLhyrW5wNhrBxkYX2BF0GVLiyY9+z/Sl5O52suiuLn
GBjagNGp8jyDoyOqf/4OZBXK+9yijh4fgT0V7n3KukHP1ircEhQosfgpHemDLFgp
spmoQ6igd6yFAer4zg6LT8jKKnz6+s2vNZMwB0vjM3bYwnUlleltFT9dfM/lwdWW
AmeV+8cTHj1nrh+nbQ3S2OsQskhti2Ifr8Um3TXMHP9Z1dSGet2+K2Ve+JEAUgCJ
OyCvTrbY3hfcPcJj/jiOgLX/3no0wOniQGyYx3eSwzxRfdHYOVQyQrRbJ7C7h2fl
9fvvkJn6XsQ4IX7SmBAbJ4/5jNFflt2xKCvkZlX0nf0MNhOTPKvYFNMAS0mIPL0G
Krue+cmu/3GIBvliRYeovPR2iOViAojwE44ZlDtFthKBuiM2TFF5BlFzjn+si3hl
V0BNtQ32lZmnX7QVm6KxnPrRFjeMmwjT6JAjuodkRZiwjPG8BRoGj4f/f0vyKT4F
w8av/t87JqQm+ikfJD3UJqUGVlW+3IvmS36nVNbHAmEzzcVMOMeVoYhuaUqZJvJV
CKohPZcFiuqE3HfikzQiIYgk5u/EtrLThCU+j8b3BuAiQGryL93TObWCOBksVDQP
DD0/idIhL0ZLAzBi68v2llq70ZGjZTJukMV+YvSyJyUD3B4pdqhx3efwbYNwMT2i
9Jbbg4/kpMYmDwUzjRmEMDBiAOeOdElCMZnK7WRMYTnMsOZgG011eTUDzlQAoDnu
7giU+xiwefDJ9RsSM6lyP9t2OBrSXPXDhgF5D6F6GrtM/bA252yv3N7Ym3VPiX/B
2fMJlX8c8mSO2M/g42W+TxunbGzVwBL50g7GUriFNGJBr6A504gNQCKFm0ydsDiz
G6YNhgIAD2vXpgWRlF9Olh1+HWNrx8np/pIYE8nmcjZAzH+UnMueYnhYQaVMC25v
y/FFCysuEWE5IUhoUZF4Xml/9kGYC5CR6EhcjjAZosQtVHzIbRnmMY1zMdSy1+To
yHeyJ+UT28hsBm8TiPeb2T+9S529VOe7jXM4PHSE06DMMqwJfgS+H0dcYpOv9buZ
4pNmF9xRXlLLm9NqTxjZRzuTq9KG+C+2NI9WTwEaILdRxsQ53hgwlQt1jwY1e7Bc
spun5B2NRXo/RR4seXaQMKAD3PGFnGl4dgaaVYPHXQMSej08wP+1hQevDU+BmGkP
/L7iwnwQNL1+Xer0fhlWBMeeGZuyuAJ6mocSn09nQ5Qz+OoveRycr9JfL0PMWRmG
FOBQpa0VcKtIeClI87z+JxuBq789Is88if/WoiuXCHr5dxDBW6BPNIin8F2a4pvg
8RR5gsFntxXofHBL5r9I88qt8JjhRPw+ZofSNL1OauIwyywptuo67i+IqU7O7yB8
Rd/rC4JHhxZQHP4hVYQ0APH6nCpTnUrA5BdIuN/9v2/oCw61bSHWXtJQZQBBLI+6
tJZAGjJZ1OOCTwThdh0U+3E5TuKtIQC+RE/CMapaZ/iVWJpMow3VBXttmN0J4ZO6
+rnUp0Bg8OxCA0wQ+n/uvg+Eaa4m+seqmbC19hgICWmrnLsRGcRRjC15w3/ZLxiT
opjHfkV+bOvGoli/1sdHxJMrGFTJrEk11RfiVUR/fBQbmDh+aN/rbwntj/fXwBbe
PuU0KCnF21dTSlqxAGQvS5gqI27C6kak7TFIx7xgCD5SDN3hL0kGiKnbv/8CFRPP
dp41ZXkzRKA5X7HbcgpfeRPirBo8t0Gcz3SuPbMtSdmkWwwv0gsjEgtprVz5hKLw
dyKDh6bVqGjMuYyIzXS6XHi1ydW+jypMRucMAxARQnqNk1Vs2/JRpdyCqf8j0IWB
cNJkqBB4uN0cpdtoJ8VbcbBGO+RJfUV1tz2XiAIdrNFnB80amZccKgG353kFSW+A
oiRBteV3j/5ZukFXhsHyW2wjHNdW2JBJBU8qfDtBgaZRxeDKMc2w/meau5WCe/h6
IMtVNa+NRjAyMCyTfiTs2AOh2gpXa4NW3ogiil/GcDd/igLduUsQS1ju9SA9bm1n
30dIuS2cGQ+WD7vgdd0LEdj6Q3dP3sxvJjLtb1kW78GwcB1H5fSqjtuLrCMq3NwU
St4IGdpXXdzlbLsZzqUAwCt56j8xA6iOx2hIrfo3yW7p6VvfzT75Jv9pHplWXwxj
j+cNYgeBAE48+xqxxcY1kZjVhbaLlMeVihs2cuOBeCJP0YA4SkGe+g2i6rxL1LYW
zH4HtIIsVcKi5Sn3MJGPpvfp8bQ1WaLXxTL4Y487NUvEQtSkRxQeOoP3j1CtSVzu
TsOOrt2uOx7uB2wUegcwGvl9W0Mp+cbz//0V/sPyuOkS9vzYsuNKBBPUW0v1lYJ6
xZuKhUNrpznesFkNMdh9tHT1tI5AsDOom98phvT+tahMvm3PaSoszNMurybBXg5m
1h7Ne0TGSvxzx5TvJY2F0oJQFgy51lF6xJVwESW1WQp+JwMLTqHcumb0mCr2w6g/
g6AAE88pwWbtEJ7S2sq3QaQHebsWshNaLb3tpC+bOf8Tlr3Gw6OaI/qRcLD7hA5y
m0Me5Iqx/EhaOF4vQaHtDXoc2ASjCtKOdUNws4UKTuhIZH18Jxvt8pPn1GQ5eZTe
xWAmijLWp9ZfFyMPq+ZrjVHtz5E9OcdS2D5mTYOJHZCCTAtu6YUvTRSBzorNrst+
WyeZR7NTKTt6W/aKJftumyt6Q8XNpEkvJI/jE0WCI8PSfkrSNju8zJ5JV5MgeHGY
6Sw8Y07OPinpv7rOKC7Kh2DJxhd3/Z1dgOQPc5FlOMU=
`protect end_protected
