-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QVtWt1GhQ6vk69iXliubtH/vGyebh2/YtafiFaYCZknlxNsXLMtwObJTylt5fHeEnl/Z72xNcBHV
en0Llit9YYj9ekAi8xxN4/eisGUeJtVHhsYgOzvgNJtVXDgx4p2RAhqxh1JmqCRjEc3o/yfbULVg
GQCP5DukEkn8twKkL+RV0J224AT1Sfx/bKHyl55mfA3Qc65tQr6tr0nAKpyTRDdPtsfF7gXLEuWZ
oa4cs25Va0w4uZHmSkqdz+gVHYSzfSf//lRVvKHY7aSbpR/YJ+Hlp/muRmc0wxrNcoHEv1JUL+aW
Ba0YE5lwfa5SQ6ftGkic5gFwakgq+q0DyEWw8w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21408)
`protect data_block
S1RYn+MUhUVxHBLVzvaRjv1IKEEPh42f5NN0O3P9+ElN6OJIMwkIl8cEFc5VH5WKXf4ut62dOxHz
F793Mce/HHByzfbsQPfBMn4w6zXaTQYcCSeQCjDkCfFQP4RRHCxAJSVAtNjovkP4MtTxQya/3Dri
eKg72aWbg1y/jE4C5ti1I9qZ2YdTAXqbI66VA72/uoRI/Ur7lRBM11rQnT2iFEicKRtx41xOwpj0
/92ZrdmBBA+tVORKQWhR4s/o0Hm5C+FLWp6YmqJlO+aRK4cwDuVoi0k58PxIjhFM0JRpaQCfzAaG
2fCr2eblJD8qomF5dUoY5TUJ++7VsCzSTuberC2GaDaEhKCD52+Dq033gYJdrcTwkFkgdW3kzNOZ
ciMFlRGRR9Orbkkm7ZPpmmtbi6Tin5faazN1p0Zyagl1Hz9XZhbkmA60UolFfT/SG77FCpmdb2Yn
wcwIqyG5jJrE9Szy9eSZ1gHqjwIbq3UOS79TKD8yqgV3XQqiOpx4lkKGrthhBfGkDe4QV9+/1hsR
Rc9+61sVu+ahBnbrxYlYFCxYWmusYKnz/CwmAYQ0bwV7u0r/A2UYrFcBOXhwTqp58HYrbBlciiUu
t81pHLTGXwDAoUey8YlFHEyRfVmlyIyt+fU4HdadH18gTSrt35OCni8M+ThYMWIfnC+SKsEeJ9z2
+n5z+PAJ36OsawoWJEh2TPCQfOB0I55YcOu7KkoOQW3yj1kbAqcW6PIo7DNITu/UvBjM/9YWEuPZ
u9f1pJzTzLdonqRopiSyB81dMDulxhhaIcb8kMLL68Wwi2yC7/f8HzYuObM3qzyuMxM8ipBOfi26
pmbTNYM8V2gAO6qnyOzJn4kHNdq+zWQymUNDrIMAHAwD0ThqOYsG8vj4y8KZ2avMOsl/U8q6iVhG
IMHEYYb1UMiu2WDe9N+HeClvgtdHAUvISBSJvS8HbhAYsdyga/oE+uLtp9sBdyBWgE6LY76D+jrq
XZ/N9uwgc8h8mlirU9OEY4De46XHrKFmvF9cV2c/pvTFuh+c3Psiqi/PJ5JPxEnP70CWG6aEbJea
VpnfFVxXdRZd59T/392dxtGGhPCP096wBn/TtwFewqqofGGYa07wz1JYOIj1WxLFiUWQ13QjUQXm
LTm2Zdt/AcbHZJ1R9objzIlzbgDOmC8gXcwRAoE6PW/0O3NJVGUX/GWH77wR6KYQ0JFjw/18z70D
pC8LBi8sRfxYahSspNnUUloTwAsH07Vr+EKvrpZABUJPWKpAq3Fk907CYoL3QPGZaq4ICugzjRza
Ari4A9spHD3L2j2RUXnj5uG748h7L6aVAaafKk+f5KkGv0n07MNrRjRYx+R6ssqAdMFZqb68vISx
3u6v/IyPgje5uUeOAqJsDO8Io9wuBnP07SkirH3NT8+1Q1UK+SemTDNQSog68cV546aVBCsgi4k5
35ysyoibSdnxXBaqnRaDetKX6vNnBC4a5qgBp2vK9MpOQk1AaDAftp04W/5A6Fmgp16DPZF+KFOv
4y9aY0S2kB/q62R7Ajr/qesCk219/o+H4VPqjArm+pjZBgGqdjhxEJKOhNNaEfgZnuklbJb710dr
ghEh8Doea28c77sEjoeTBWkRmlpaCqVAcJMJgtOy15qVjqI16RCj5kp/AKGRbbZPsS5lw7NYc0Qu
8F31fcjKy9qCBGLNI8wUSkgPFs5F3pjdHThl16wyl6HetWPiL4gAAwzd0PwScJNPOG7QDdJa8LLN
tBmHLN1DHodX6LHVp+8r3FdCcmljAKVloGCUJTlgQjozg3k+xfIrbS8TPwC8zk0bvegESD4IPZAC
qnkWKRAKlQvSydeMW2jIhgZAMLBEHnyi3wPoGihp2BWoNFoKPKuP/VOhZmnwBtSFnFnYFFDabkGw
55m/7sMHVJZqG9ZmWIPilb0EIdWM7UcTpN+r6tXzIdKHSD4V8kkKga+l30HYKukEkUt1wmUKHdBd
K0sp/Jtrc4iKvyZuLRxhSGn9zb6XEvL2TPQtgKt9WS21Yo81x/acBWby7FKeX0OlMriREihdVINN
Si64qaYIvIKseh/VuaE3qTlrG0YqdzVW0PzjCJ211u6Wl8d/M4Lw/8XginMez0mhMlS0CoLDOwDj
XRKsEKIJc+xKtoDRNvBLnqQY2U66ajoKflHhP79PbF4rFKnh462UtYCcHArgO91z5AdpMXbzluFP
rpDGsH1rsS/L6wJ+5FisdiQkVRDGKrL5ot4N310E1JWNbaTAMDTEQrEWImEulJbPvF6xHvtIEEyO
z0eOTZhhdHxRhj3A8lmIAAC6tVzo0h+G5xY9g1OONzLQhAL6YWR07fryK21IDk1Nmm6lfdA3lYBr
S0IBGqJul736ZhQzjhzC6GXRGtgOnb7xyXyy1yLo8Ap6kJG693ZNMuIdOKfcw4iga98lUfuK0+Ir
0OPPUHJVVHY95TeAs8UB6gJ8hF5f8s7pbQjE/AOOPcq9XmZOWhi4wNo0RfuwB3KM4Ddva/qFJU1c
lzypuTa2p/dUKJO3WYvsLe5kWSuIBcz2MZV6Y7DYEVnljAc0+gKYtTxelwSOejbPxu5gtPFEn78u
qJGP9JXawXorkKjvdbNpZ+G1FRARJX+q9AVm7U5t7pZuMKnHRib/HRGSj7eoGZ+ahBzo2Mo1S/MH
s7j1yPeD/TBWjD3QWwt7cBAJlTzMwfRml/drZVW8VYQF2hKD909yQCXTLgbWGS43I0aOOiJkbqZ1
bx3HKzu6UiPsjuPFBSUjyVrDESElhtwrBugbxHOmrQepLZfrwkXvHavQC613NT5l3odLZD53/BLj
fiFBJEp0wiFcgLXrCfud53E3BRJKdB/m+uKQUA+SbqAOTokrwNHi9QxZ/K/8jup0cJHsjkz7BUYN
hpRyP3DVvVxdJLXj3pJpXxIWciJdTLYeWwS5THJwy7h7vFKmyxuUHxPWNEgf9xNh0JUz5lvudmhF
4jCqbUlBUDKLAO1qr6xNLQgArjB42G+gM6EMRPMqjhv7Quy+eSIUXUTMYR4rduxvx795LILf1s05
0UC7KtIg218++dOMBTKci+/WnCGQ+n9whjoZ7O6spfwkOH3Q6P3DqkiIAuJQgATQwZN4N302R6Ay
UMJFkGkNMTA1KTA0/LAh8PHNJ781GhVp4fPQoMIXsAfwywHTKKsPto6wFKhsn0kNdlG6XpWLlUtD
iT3eb9cVlHkkSspFMZB1L93L6sl5Ahfdb2p2oRAD236IKguFfgg64ZiZEmVXKBWqynyAxgqCTbv3
oS8LSU3r/dYoInI25H7uLKFuUrzJWcOc1Mu9IJd8r1ln/zQr7iKLXa246LuOzhWTMTA8Qdmzcjug
csheRq90NjkvRnnlFGNwSqtyObc4rU1kPrfZGe1D0Ws+TjgGDw2ISm3qwstxhSWJC5PyGpdXgDjX
FN6TXP6BVIJDRATCgQnEgUEpoN3JOKAoWznUtPSi6+8m8T9syN187K3H+jT0BMPDluUNQbGUoviw
1tYf27dlu/SQ6AbqFOuVzDkIm2TwmqM1RnEJ17T6svdVa5v15VyAWClJLFAcFq2yT/O5VMqbdWTc
jHGhxazPZAqopAEe4KGH6xycOKjR+r3k3m6lfTeEvVFuVe3sYjQteRgxHAi/h40/Xx8VoRbzVHbn
lOozcyYG0nKGC/DDJHUUb6HfLdBDaGrDSxgmyJOK3N3ATSuX6HvVQ1GmE57dxIbQdoGF3yCi7YuC
Hu1YTnYP7vF+0Lvjza06RxoXwWlB3ioln22BX8wOS9e566GwRKwgmYHxlQc0GN19vY1cxaJl/MAU
qzpsoQZSPR2vekrUT2ReadSyFIEnuyu5cSX3VQzLSwzTvIln2mgboWTbd9EL3eOgwdc/JuLfi9Iv
GvNo7ZkrT+wOrcMIoglDi7p9fHTS4tKza3chWt2QrY1+HcRDh3FUs84Tyd320JGhMcOuFSBNwphl
p8gHZIopigC8xvG+yGkiBoBHNPESq/iAOP2IFORjChGR0+fis+YDzsMesMWs6pViRWLna+TPqF4j
VosdnNb/fXai5mBjSrzXDyUaf0rvbLBLuX0etesreO70U05bRb13UUJuVH9AVLfzEh1VxLtxTnvR
ZcHm0TP8/uzILqrX2Kcl3XDoYPrzAeq9rfLlOxPCGQThWqL0JS9NrkMim8ShG7YJdICmazw6x8cU
JI1HoVEgRO5738d+35DOeUeceOTCpPd0ar0KGCrh/Qo5mXK5YDzkV5+QcCub71t0gBHmV9kRAwz5
baffAPTMPew8xa36D3pLNbKhb3bGAhBHBBn9mMLFpaLb6qyPcunq2YG6d85a2C9ETUyyVQbrD1EY
aIkcctNfpvDjVTcdIVcfHgeokz4ANhQKh/b/NCisM/qce887kioZnZjen6Vi9+RbPFkv1nOwnKMi
JWn68nBTuM55Pxas955qHEeItcgNNsf2rBiDKDr6BKPDzAfirVzkE2yPoU1lu+kRlBXMATv1pug+
H4fDVjqYvyVVp54Cq1d0UWwInXBVYyN9TkFmAewfb+dYe6SSLMwMBCWbDytg3NYzoczVCBGBLdmK
ZM3tfljviNGSzL8CNII2qnJnDfAyKlWoMzmNhNlELJYAHcnX69aNH006sGUGZ6fqPS/RZDeU/iGH
oI/s1hgA6wNjH4MX1AG4IzS+THoAsCZkNHprkr9lDAQPKMduZytdF00AeVeyWmCO0wjNgXHG85xJ
J11JnwXfylEPRtvxWndOCTPKfhkGQuBf/+wNoWjpZk9MC/Lcecd7IWaKXeYM5Nm5Ghu+fvdaaZkO
VXvGs5QPI6yKb28HheaaDRF52GU9D4uio4U8r7It1zsXx+5RsfFscmS27Avaoou8WH7c8QHb/fzF
nXVJlXG07YrpYR8zMV5KC8LmP6dYhsQlkYCC0lO6N14QI91VWic0kXbyWg0R5HoWeGUDoOrDJBF4
1R4D087k7Kra4/BcnsvDpQbdPFFjN/VhgGRc9978G2cAz7oVquySCqFayyzeQ7+vXViaDsYzULow
pYsK8TxpWeag1G/SOCAjZ2bDYOQDdOaNC+q9JkERQnSTVG2m6aOCVwltXeCbCWOQEd806UqnnigK
Kfcbm+CRSPHjzL6FCATEvy9ElIh+Q+QPKPXFBtsZT6Skv2es8MBgm1vPV4ov1eePK9/2MWzI/eMs
wamMrMdD+rOfV6rvBGhkCZXD+chtc1D8nsFff1Go7lsIrGmTN/uwvmmPmzhz4w3WiAZ+T8yng4DD
fH84P5lgiImNebmeCRZv+E1TI8UKNnXTMoBOQa/rzs4U/0Rqa6lkcRlDWy0d2BZ+0QRAYnTGVlu/
SKhwe84UBqFM1m2jFfYYRnUS8NMs4ZoT5clqNP/C1wntJoDqPTxEz6QTxrHOwGOaKVXEhd7PvFsw
U4xBDRTqpXehHFQl9DltQqhBs2yuEfcvu9LTD+3nfdw2T8pZZRI+5cOF9uqYukCJ6P6V2eQBW9SD
GTQum2bxCWMfel5F1uti/mh03pgQNMOaZSrUlqCGUHBMDLe3W9oXS1prdjElCOohIFSPmf7/RPnt
8ng1/Ydy4cWdaNKmsP0l/FzuwRWFG0ObPpZnMermkH5efp80/22JBnegVZWM0nVz/9hpXJCg1jWL
g3N4gP8q7Vmbweb+11U5YwvEew5QypGNHGX3D3RotpUPAQzYb8Ua5sBlUMAfAh3+8mZNCgl41ele
5DnC9kyAr+dx0sPSYp7woF8AllZkY9hyKaiuO6P8NFbThKWaw0dChSbKmDEY05mEsHCTFYFJY1mT
h9a8ULz8lfsBWqj2U/kH3ymTUP/485o1QaoZ2kn6hyvJbsMobjy5sjYszPQNBOKU4gaa6BKQEHSv
gMYBMgUZZvbFxHbx1bgYCOo6usCFNX8LB621jnvFR/JqDVCAF9rimSbT7w+5o16QseeQ9Ah0LdgI
WjCmDjHE7EsihxwFdf/f3WJWstr9kov6Y2KfdS4wC3yQZ3H/3BJCJJYc7l+xN1pJsXqnltr+eD2F
K2XcO8Xpi8jJWwcfQycg354dgm7QJZJ9OTtzvsO2sOg9dFLTZKgmgfhQpnbsTeGE5PkCWC7RwceP
Ju+jVbYOi43VWepQ9qfadXSDJAcIVCMsSpr7vU/NcsaU8az2YnnG7jE4cw7yFK+1xm0tWTpBCetb
pejOs5nSw8a9avkXDNVhgCBZcZIFFODWEE9QxVVrhRuqfbGrgw8rD+48fWHQEh8yW/SD81+YV+HN
8xHgp79y0YKFWlt0rE+7tTrxKrzmplezWpT4vC+KEx60hKyLoamJGY691V5FSEEU24+Zv94tw3FZ
HGxgyE9A2w4h0y1KhZsjAZmIm4afpG8FkeKeBls2VhtFfyMTH5/7CIQaj76E/qNwF2VJ/qpFEety
hAW++GoVzADDq6/h5/NhjKvHy+UyEnwINf0AVcvzv/bp3K/zR+4KDruCGernR5OuEshXf2JILTBV
obyssZzDLmLafafx59cO+mOx592KPOWvC8tx30roirwXk8fwABUtncUxWpwvUjX0lRz7o2gk+4Ne
/1tBzW56RgfTcgE0SRT1lfhF03dLHmMo5bq4ahUffFkRwW68GQU9k6GMhOL1sTcIaT6djtjd2NHO
IhOT/c6pATf4gxHwqaAg50rK3BWTrQu0u2s8CFzxpbhiIBZfF0MBFyChOoKw2GgQ5mdcCb5LZjux
llMZ8EBIXWJCz7Jxl6IJYqROy927q+/2nqvprGMtSIfsVGGoSDQmB0sk3q94jlcqQmVj/Y0Bvu5p
6+uXTK6YK8I7GM/JDWw0a3meaV+FooYsBYZsxsecAAG86Q/r6HOsmG49ElXZjwoL733D2p5L6PFN
5PXP5HXgUjprwnFaVhLJr1KzdttslNSafy6bcDqu3/M44T+VuuiL1KHqTYj0qXA3GasBaRg4aHKv
GDUVitPkttJbsmeeC57XLd3jFbFemjuw37YPpPV9l7QdVKTlJ/KLcUCDeJ7K11AeL1PlCUZomkd6
E8rzKq3D6QXx5RHAKyrXcYw9q7attfGkYoCGEIQDqiaYfyYpuFi5v64Si9XhEtqozvGwiXSxOmoL
x/PC0ufVSI4tH3qWdJhcqAWDhAEZDYJg6iAs6zuZ2BnRRjb0LjMY3k91DboG1BCc4QI6an5xbwrZ
KeWG91S5VnlCpjqwlP5yms3arSD1/Olj5RqJUWh/jfa1RvqurX8cVHiTyaMMJEfVbzO12ocDQIlR
+ccEjVMEmJgCFysrJ0LWdQUAbgbjgYx131bO7LZ1yjV30dvjb3pV/c9oK09CrMFrf67EazswDNSd
TnCgUrlJ0a0BBe/uWxR49AUNM9oNmVsKlxQ03ryRC93JO6HU/hAJ5wMqgDGRWtmLEm/cGilyarBq
b//2XUROpyr8FqRO0NGL8+52JI3ZqZ4mynEwsOg4B5UyUlpprYPliIOPaUXS5bsF1vdhm8ziw44P
3O5Au2nDtKuc7/K8mGEfRqOrRTRNz0/HiW9TNweysCfq68vxP1oXHrnbF30kl804NqG8R0GjTWH6
5Pt7MN4yZjE5Ojac8fSM7qKW1DFBLG5I6PNA6iqE3vdi07EwTxMyvYbsFSWHJcHSOy+ilRQZo9gw
F5/J5tjmAHKztlGXZzkrkGioILbf+ErebV3HWbgi0j7r2/L5tbcnqnQLBIokWzVgW3mqU4cjFfmj
QTqkhGXYgg0FmXrAb1m1ar2kWqt/BGJLLNKdE3ON/UlalV5XixlHG3jUbomwE00ZoqCF8xDBMka6
G3ZZS7paJK0XaDg/gXOPdMOdvVULwYpn3CGK+Iw+Mh0U54ZxllyZ+qoe411YcM47540V2ig3qFny
8yjvDXxbiqgwc65TBpCPN1VZ9b/1zZvIfWM1K65nLf9ec0UsF3w2+wkiO8RHethFq6gthn3D7F03
bKlBygHCKV/H/yey+mdrHY/gvHz+yj8rFOPPloNLHfEr16V6ce5AmUbDYw+UAPKk05kA4WgjO2NT
+H6LebsqD4vSa3VQRvA+MHFdRqYTqZZ2YlYQj2orTGUcMc4bAFe3lqWAOTz94jvEJVhfivScX2ST
NPOHzZLrsdrfyKL1nqEGIj5R04E9vG+Qhf9Pl0oaZpPCcAkwEB2u052NfV+4rNWWchmkfchp1xST
hzUeTQAykFY0zYg2g9udUFEN5gQMq0t5P2aGLTi/sBkRcHomi52CjeQm1rRyWGLdJDEx1GZtwz9r
GuqWEkn5HNTxNFEcOE0pnXYQzWToJxlJzkN4J31pMQuNkj7zuODd5Y1himew4BqJczaF6bRxUPEE
qapSHc8dZ7LRqPPLNgUREIbJ9X7kHMSQu669x3Xes0anaWDFq2aqPYStPtGrZ2Q+NKrFkqlDvhvM
Ta+J1xh+vFV4w8p8cOVSAgtinGVQPm9fbUY3sDmiQanjj/+QA5SQtF3DLyNVWCi5rGYUXokG8pgQ
KxeiPlgCbE/i/o87YmtyaRtfchKBMr9wA40JqbwenB5JcPh4SNjVyr+Tqr1QJzE64DjIDoo1x+WO
d70vwPxbB1UX8eU0w3Nn+hnJDxKj3+d3I7pUpFCmChioeMRoRwabxXI8lRhwQzrDfK/6IBVpq27P
I0H90VwOE+D54tKaaKwIBgS3uSIzEEqg4mU+cmU2aiQuwv1oPFi1avLJ0XCmqG+3WHJPLnXS10rF
TlqUEzLWxGHRt+yp1NNLALiKR8cdiudyDabdiZj5qNDKoZx0nOGobwtEL5Q6y1lJ7Y05m+y3pnpx
OYlB+IzNhPBsGn0tvud+s74U7/yrTYdJ2zdCYDQye5EThVfbR7+g7rtfflBvka9Rh3w+8KfUpypc
mKn5eGONTLUEQUPXZnSUiwSRR5ISE/W7ZI7N3xCeUxTilBTv/OMU7uHOYZRODPOSDy6xBvF6Hbf6
WGgFIf1vaUgt04ugWgCKEVkicZpd0RsWUI8H44Js6NZBCVqG4pV6m6SGi3s1NAbxPzGmDWyiWRPf
66dQVxPVMNoetOPdJ9DOexHpM3SwvUCqZXYngHOtrXdT5+Fi/AjzbOKmjHsuk1hpSdAU891ne2Cj
JVhytdMhn8vJcw/Uj1FljAshht0+o1zz1T+e7cL/nTYzmaLqYZev+td+ftzJN2/zgbZoQZWdpL8G
zV4XKqNJqaPDhy1FGThFvmkN9cZVSnPgKd/6dmAN4mruWw/irPTjE1EMNEjGBQqZXyTNYtMDpEDT
fpq+w/C/IUjQV5W0VBKPNKUdXp6PC8Fw2S892CP163Y47ef0g1M3R7poLhU5TKpumpNqSGW1XkvS
6yE7Tn1BWbKKTGgvCXq77JRJMSvOmV9MGraZRSJCX3m7iKpwsjVlfOlZwEquOuWQPExwm2BXFB0D
y6Uy9tOMmjQ4LlOPfFF8Exo4seF1fAOqTyjZIu7rYKk6z/RYo5wS16h5Byu9IOI5oBjvRY5bEKIE
qQNS4KvV5p3fswt8OTxghXMSapD74PWQAcoyUYVmyAqrhW+VLnHG4XX3z1J6K5adqy4VPn/JZpGJ
JLedTXLV3IPc82dh7ZzcA0dBWfqLpGneZWI7Pbaca/Ub2nkGtWaeWoNjyW0jJrC2pt8Q/CtAw+7Y
mCjFxDdLl7XDpNZgK+BbN4GmasyQ70gA3Pex4ZaMB/YYoUMQ3fce8KSkBPlKVtfJ+a95UBQLwmlx
g5Ub8ky7BuU3ubQyHrMLuAPwrxeK16qpkpgh447CKJKYoHCi66cE/255qhMtcCM8cF7yh2T3rosk
kTyhN+AuzW5suaaspTHWCOyObOJP62kBUE8MH8uU+rXgEx72irCOofLmuO2l9/L2TO+ibZlZujhU
hVYaRDQHTfdbKRDarGXB/s+PbfbesmZLG0sDmyopzoVtRRpnUVk+0H0/3Cv34suYrARqrneeAUKT
PhW5AQBh2wiyheizDzJVLWfLw472T50pnQC0oJxq3VFSDxY0yN9zfjjBZWWkgFUHNzvRKUNBbBZW
4poXZroN1onzsfnf/hAc+x7YLz6GDA02hRPLjETdo8fJAecTn8cQNMI4dWrvPGOe7PZMz8Ti/xmB
0Zsmp1xD4ni4tMwyy9pvQWkB0n1V0MKe3IDVt67ZwGnvMqp3IqzyIjKzIrtlAqCcQhKxU7DbOJJb
cpAEc4wcX2D8ZSauUlWOWpSFlg78i1/8VkCWy1dPHkDPE3PhDMYeU+0rApu4OgdlPyafPFMD3QpV
W8PCpUdBxRIp5waNf+Hlj82eyb6lvmax+RcwpsmKCGakDBY0bxrSF6IyNtPLfmMOr/ZfUvTu5OkJ
DRKaFhM+Y83AonaYinB+iVgfjVHTNToGOPCc5MTUOrzrB/nWxTSkz+jM6VZxRinT36NU6vFAetaH
Bhno56nvh3lJMqFruXllLRzsRUMPW/T159DY0zHy/vblti2skr/GjH60b7kv9uukL34NJ9i9wNo5
WpiEVdqscKhfKL/VjSjwpj3vLByZYKpx6iMcliTNumlJ7nkK1r9H7V9SKF6N01tvOXRCdkJExPH8
kvunJa1NlMOkBd/PgPxWCS+REmf8urnKhljvkFzGFC9rMZG5hKVTYbvZdEU4f0nxN8R60A1A+Yg0
tFDfmuPtEg2WxuvEVIjpip4jxSorOZdQb+ql79k0Sto9jkuwizXnH1Nq8bgUJkhuZ1BW/IqUB9dq
iimmqUZ+ngu+GXfo0ByNwzHI0aqlgEm5VlijOA9U7c7P4eeUEcngqFOHLbmi8LwjA3As3IdkQepQ
9pjLAtBKyNzSVsMuUqrH9/FahfGHgTbnIhJUuUpbIMwYvdGCURjIlKeb3GLzYc4k6B+7MT6GZsr+
tVibeGNdb99e3VTpeYei6ZBFvBScKXDurDGW6/AdSCXJw8pzXnn2gGBTMehdqwArVQ9gB9MckiKr
w1OrYlZ7wb73Ja/DYBeU5B51b1ShPpALTB3NvXtDr+I5b0Ij97OfXPd2xG/sba/3spUGo0ImK4tU
yF+reAB6js3NtDICcQriaeMOcHWWjaULS2HvEhZOWIofQ7nW9rpZDSkCGqF/Ta5ftPOt3ROoDDl1
Cr47O2Ntl7HZnCFOr1g/QW46cIkUoRH0F1f5Shkrn7RGmRKZUyxpvS+o8baqwYbMo1K1AUaDWdOW
sb07Y22V39dXnlAAYGizeMYCyd3Vf0PyyxegA9fsnqXqAH9P5QHx80n8Haz7NONSk6m14HZiGNTU
YgQp0AKXnlKt8HFwuZHJy+3bpVfvW0gIE1ZHYEFBKSOnGWHvCtDV9PKdQMDm7/pF4FG4xAV9XXXs
61vshG14Na6LPmo3wL9skXeDN3tgFDb/2vBwgEiCvhGTUBnbeoPNZz/e0KRyVRHTA2mWglTbfPUO
y/coO8T/iCZ25qJAT8wafe0AzqEioDBJ4Q68MRxUtKyR61dxc+kAbfst332oyjfJiDQUXCQclhlZ
Z/w1H3KN89Iuzk34ZpR0nfNkCqF/awDo9STiuEaVfQNZFcWGqw6K6fT+0rlwUOD0CzPaUo7QB+gp
3mIpMn08EcYXwLLtyxeAr9zhQE87siNbaLKR3f9wQp20twAh1jEkTZKcyUYJ5C4om76e1Vx0Got5
t5kxWshhbxdZquvmo0F6YpV1/PDI1TH4kWs9rv12xzeUQDdyrWaY8lQWvk11jh8CRY1j8Bblc2Om
aJNOa+d+bPf4V0sb04IlcApahHQbgaXl7ugUhrShKOGCvfVP5ELBZthKFQdkbSypDh2UXdLeZe78
fZ04Mzq8fuXYzbUqZYK8DC730KGoNOvNT7E0PWb3RvBMvJBtzoaTGLjbdah9Sc2OKrbSUivGA31/
whuXDzLGHkgMGOpAIQGSrMhtoWigUzDVj8Gf5KkNyZI0bhCr0PWmJxXQDwQzxYAaD7A8gDQKDAen
5jQOiDeH9gbevM+ri/47WUeNOT8PCWVOj7wRTpA/Y8u+wm9yTAOA8Ih2rW+8IL8w76SAoNOFKmf6
lqFZvoqcabJD0ruOs1U+7xdH9+gV9+bBvetCXzoZH7O92jq24lKv0utYWcuH8BiyMs36wejc4lov
OCvKLFjGh+YyhgSnJ+czs/IxB3AO34PGIEeeMq9WuClq4Qs4nUjKeS2ONdgLhm9yBqd55O8uAnC9
9sSOh3iIMyKUnxbvs7YJNshSpyQQmucCvmuegVHluHNn9UzwFuEd9Zn4JH6t5kzj4CJvUmjt7XgM
7wnDPomjjDpLEZP+ThauvCUsapo0TBUcMh2UgeVH+tlqKlBbwm9bwTQOYzuNtqWT981+vgaYOb9X
5cz3F4RvGHF1EdD9EKgs9FLsjN9XsQlsbuN/JOiKeGdkNuILXEn0sLo+ROrYA9ELEmYWC3hSN3dS
32UWbvhDS2EOoZRjIH/QXPCIWku6D3pIVz8Q/5edEry5UoQzWzOK+AGAsgW/WS5preKMMSE8oNjl
GZavpf3Z01GBGOBcCthOySsjkVO83wGNdjYyDWdZfQNWGeYLH6m+OS0w1IxGfzvoazriP/xCzgyf
b28RCvvBBaelgUbenmvqa3Z0rMecpqPS8XDe7hNrtdT4KLU6+AR+xz7u1jpH2wfLA8ZhTJjEFAH8
Qbxg7KhSjfmJlGai0UXTCuByUXbfPu+IWCrRaELt+L0meSfHKEJK36WY+T7R4gNmpETDJwRTxOli
G4QlzWBUcRtzAfqOH12LJhjyQY6FibCEYbPiTJZ3An++BGkmbzfk3TZ4rv6JjQP/6GIeltL00Vmy
PzlJu+2NXnUOw80Z+cCICxV39GCs8V5t7b0yk5W/aI3ZtfPlUtRnGaCAvQqA8llnk/biPauVRXI/
ALfmaHwJrUlPKXuKyzbVB+FSdWRVA0scbF597kN0x1o1geTZsKRfXAopgB6rgMDpKSmQBqfbc1cd
E3Q9/b4Xu3BeoPOcMgR24yCTZVx29gC/mBbDyK9L5I6bW5OoVuIXJHrf7bOWR8XnwfQElO7AjXYI
aOzvVOs5UeV+EoiOnXwVBXrDCT/96v0+hZgwQd2QsnwLcawAZN+1FwKJJPB7BSiCjMhS1VGQQT2h
DHClqLOXOiGP/NARPvVkZTrnu7h8VcZP/jKudqsg9JlhJoC+gcRSX99ZR5ZB8QnXIxYkp7x0kytO
ZwMt0xtovv4ZkrqvwnzRuL2FSrxnu/di7lf2wiCIuxFvLJBZvWm7jV9PlKUYdKSYSBqaWFZffd7J
BvwkG6NJ6fYPEtLSZsB6F5MLwzgFPZLBxasKiOIrfeJY3yt5k3g1oDbNt8AWizhNjszR10EB4c2e
A0sdr2wFTVrnqeeaCmkX1xKBpIwbQpsa0lASu2TTRCmd6vzho5p++1pbWrDX3faM5HqEadFMq9eM
/Dczv+DA4tE5edm16YwGnmUhGDwJeqHogkUbmyWComC3Do2Uxd/WefRZxDgqphx9X2VU5GSY9ZU8
g2/1ChAmaGZLNAKKN2yQQiBp1p3YZOMI0ovPc+AU4naZ2ZX0Y6KtrFYmNh/S8Nd3HQrUWm/MMjfL
vblHMNi9V2q/v+HxDyBeBdM+S4/8QdYctOecBIZWE0d/oBTLFVUz8HSRfPBJSTZ114jZygULuTHF
IFnwOi5VAawSfxfgtTM9f4PzJrzYk9pHFOrkQn1oUi2vzZPGTmLKUR0hnWN5RRahpLvEyUaNCz9z
lPzK8bPeefuIsbSAKM2V5qWm6DWfUN3S66z5pbpefDileB38FwgJXkWubIWjqtU8rzVoE2K/cPpw
mpfFAsZlDeFmarOFsaVY9qtZIuPHuNIERi5wc93vfo8oEeFkw4h19RglOUtTXnYkrL+TXn6bN2jM
0NS2vq8wZnet+EIthjcnW7t7f82yq9c+fQEGey+9gibOsWO9rgvCwHad4En5rrAZdQD7cD2wW+XR
8p/daW5HEr7nwj7PPZltzWFz6BZCX434jEkVDg/MWKAEsixkFwWl14lZQNDJvaf7O++iyzEZ0S21
0/n4lmhp0iOVe89+pXOw98BiH9671Yd5mqw5Nc9nhEAlxXWBRHqhSoNiMClFf3/ui0CJaouE6InI
u3wy/UjE3ArBudmMbfFG8COiWHNZ7Yxd6MjZ3/35tfCrXAzHvXxoZE/PaBWNQ2wtmoCZreVuIfLn
CrHo5cp6zTKOMmT2mytSJctsGm/jTyyjOPJjfDa+tizLE8KwtoTUEHdjjCPTnC11Bj7E3l7Y7I3f
NUzvLwI3B3reQ+NELPVbL47NRx8Ync6mz9ZyUtTjVU2y4FwvZ8lOYNncBCTJ373OmrQtW8aFaWTY
Hd1HrnAmg2mzONK5u5yo72T3Hz5jFdHfIe35qeqLgbjKOOKJpXTAcrkiBwmTg+IjItnDUMPerLID
AKlcmN0bx494/2sHQOSMSuEuWGZftoXxCGuMedNY1L3s1EawyIC3QQ9ZgeV9Of2T3X+4s5p5O/bq
iOHcV6hKB0/8jM4yYMyF58zkzvzssHisquvX3SgaB1yq1BrHATRTZWpMWv6BrERaScoX6h9hL3MB
bj6D/p0VCL0OOp/2UFBjnwoe6z4mjCPYo6+ArJNqHjBVAUgKCfcupANMEbR92u9nwzdKEiWZZMzj
nHzWFgCY8kGr+5BrUOZnRX/rP9Cjz+vYFHQHprchcx6ueWKpCxQm+PJ0wnTSJ/6bGnd2hpms2AH5
/EZ4niQdy7ZOW6tWYbQvkOAhoH9fMqjvzFbB8Jr2iUkZ9ErWk8vt6mVSc8FW/sVU53cK5cf/kM9W
MI+8lg64xp1CDq48YWGJp0SHHakONQ4y8j2Hz9USu1K8C2y8AwpsqIKi97fdmlhVG8T5FAZ70ZNB
CHfwMMa6DgUlp3XKPLe+4IN8sQzf6R1/1rMQvpNhT7YDBoOQxRn1vil8ocOsNL2OZq2hx7km09rf
aa4NT1C3CleXaXKAA1/JBdhkJJCLmO1dpvElAIbVx+kKPT6Pcqd8x/D2tRI4rIzVGuSepdtZw4Sh
8whdvPYdio4lhRqFbpiJzYXty9RDgOQsSl0+b7i3pJRqskIH8Mdua43cX7niRPwR8D563bPJNjMB
KJRna8YrTxxSk/6ts2+rwTUJZZ1F9bZrXmikg7xo+8hZKMsEhndrcZ3WGjOHO9g2CQoktU0NnWVI
38gMOzGmEtXqodiCgIK8WJyufvKeJBUdHX7M4X9eCfahE+SR3NvwBUUMgQmauDAC68gtBlv7OwjA
510wbzwUDmgj3UXq340kh0Qo/54q+kOqbth+QZhBf4pdyNri0mlsr998cmgCySk4lCial21a4d7n
/uGsr2yRvxu4DGAfcWfDDnqngay7+ITn657y9RpQY7ZNXzyYeaminQ9CBEeJatP3V8aKlsWNpDwl
YxwXSMnuSHcjo9u6F59s6pr+gZrXsj+mSp8CiJAhIXd3RbanTIc49p+hZEY1EKFDYP3UKgUS1fAV
HdIgxeRAS1u9wys+UiCmhNVknz+LKCEVPhoJae90QS40i7tT8adiDsdvc6AlvGBk8lIXZCZba3YZ
HtTsX4EBAg578J/n5R6zUWPr5UwjOJIH6fcsLg2zZk2Vk3USTOtxc8WIpa9AflZdCMck14in7Y0G
DDjEc0k/4AyCXp8PkyRlH9UxVKRtpfDXn3PUCTUPcuMnHSXGr1JpoTT+OcYhs/Z9cSA1cnjEzcv5
6PzFJgb2Ebm/sfIjAI73+zwoXcSEA4gISxCafrCg0oyAo81tSGHJMhsb+/JSGCwr+9uN14qpVq5J
sUrdv10Xzi42QlarJSKUiLhZUdE7A+Uo2htc04iS4iDfoMugdihPelRaLNVgIV50PN2guwIYM1tZ
nhypPc9o0NH1ASZ8bdnZNQIj8hECrOtNvijQq0kNsrRBnW1apcmF0xCTjtMEsSqFbS82AOkZbPiK
icb4utzfIRBDN3rXGi27N4TO6dEFRm7J/TwsAmV8uqteEuP0g8S8rrs15t8MpeSa7vb+qUb7Kp/a
rYSP+5bwlbFM+a1DyaBHHLufQrY3xjvWW0kbAoo+5o0arZSOcgQckotJZj+JvxpQhKILxXaPsfEQ
ttpdpdMYgvVA+IX1ttQKYvZkU/tVSnXUeKEQ/FTveb4wXlOGNogGu86xz9Jj6jA8yW8Y3V/fhZla
Q34xnvLR0RE/xUyeEeDVTZZDfK20Dvp3kT9kaMEDjehSG/iO/F5eVBKlBDO0dBlS81/5I+msg3U+
5lEct6Il1x68yBfVnl4qJBYeCtso2x/7nha9PL+hJmkj+MJeEDaF3M+W9SDXgC9UUXqjsCmIPCFD
SbckjLorz5iW2vWSKazSmQpLOxj9PAgFuV5N1fzG5kBuIYfE+ArlE/00Pe8l6iCWuh6+8PUBkz7T
jSHWri8DFi11rmhurJdXGvxalg3qtf3Yh/TrDXkH1b4oWc3NWIgJTuHXdpO92mbTv6wORu4sBKNG
L2PsMwf/Cw3QyoPV0n8i03BXOZC4x/uYhUQFcs1mKX9G4Oe7JT45bS5lKuEt92WZNM9uQ6tQFQ+l
2mRW+DvMw6VdnDr8LSwo2JX67hvkWo0qImlMpphsKW87/WldlFg00rJ4qV5uofWooca0bldr0CBw
+mJtQN9p9ybQ26ZwbjUuiEx16Rtj6DLshvA++szP/k8Omq+S3sABtCAF7DED6dgCmMio3ck6nnhz
90v/X6WsAEjUNt6sgFjquGv3UhyWgWDlarZoi91krMQ7SjzQSoMr1ct0GmwCc+8OzZKqTTA2WH+u
2p7UqujiNAFKSwgYrvRglONXqlcY2eaA0TbDu8JnCI8FRUbmePtU1zfbMhMxU44JifuJvnGTUHZr
mQM7erQfR3qKAGNnNq0I7wwgau+EUvNQlUW5Q0cn9bXazpkXdZlJWMc3wltvd9qlS/Cb5eNfWuLH
v9aCBI1J7z/R08jiistn6Vm2XZBiieV+tAB6NtRernCSsYKYei0J44hRMybX4dwIoYfJxD89iSHq
zqARwz84hUokCw54wgNtUNMvtngtTkMp+dd9LgfQsr0MFy8wBzHOB4aWuUUcvK364OzF7Zl2i9KF
PSRv6ZpfORW76QJhuc5EN4H5n/2FDRUS/8nBp+H0YqUxLPINJowjCeVScYiXNmES+HCFrYJDsHBC
Rayst5vjdFnl+EvfiEnYsbTjVVWKHOp6aIO43BIUj4L+vMNtuMSEWKhT9kjGDpu9HFYnxQRVzPL3
vgSE0tLtTNxBxIBxuuzW1x7C5bOdC2mh1r6wLSlcqAJjx6spQx6PMC8EWjsOVlOHEP4cvuHmLxPt
4ftD3cbxZGlHX9hczOUphATsoH1LGAUxV8tt+fLb1qaZHzJyriIThRDU+Tf43/dfADOtD4ZxlifB
ITQwx8O+g/Om/SuUxMLjm33EmaKbBebiq9781u87HkYSWfFRMG2aPStc/4P27LOAkb5fme7pfARB
0rJRwB0+7IQK+ufnA/I/nkSBFENw3Onw5oa4mVVrgQNst58K99KcWzfM8oHgCDpBx3/yEsWizAmR
HGa+cgH/9hZNybcKfUT40LGIP39CCMU9Hh1XGYWoYeWqCPsVfqVgB5or/jMsQKnj+T0TNhV+VZjI
hmGRiWwNsEP4V32ZrEKzVZ1nujFlmT5zg89enP2rpyaz4MT+A0T/qv460t4HAgaDGTQF68gq4xYh
Y7MY6AgNgAvukXGVx6LfMhBlwEiEYFUxNXJFxtrLxMMWjk/7gcsjtPUz1NYTO0fvmshqXONdkEPX
ZGLpvJhjGQ5x19Un2PBz9hjhZQMkx6bYB+Do45lLLWrKzCalX71LUAfISpkVXtE/JQL7eJsvuZmr
s/MYkZhmvwna52RnqVdtQPRlzU76rT8i9aYiKXKnaBqnNcjjMGKwuPVamSfR5eJlV1DVpVoHYtw0
jaXfE17Kze4hBMRzdv7v2XmIuQLTjKq/UysIBP8YWco8DQevEHoXsd3u59hSc3TmGusRTKP2K9II
FFRJuOiEOEokl4HmkrHspyr49EJ+z8BwT9XwEkip8e3gR4+v4qHTVE+LAjCVNT4ZHinfSNdjWKas
LNn7GY70EV90uk99PLBXu5adaJRvpbxE+wbVG6cUYr54l3kAhT9EVBPqrRqBjU5xWr6P1ixRNm2m
WNka+VSTFNLWnSd+Zmocu+Pqu/QEvB/QLlAHedpNJ7gYPenBE5FwuvOR35wg3BvWa3YNK/VyBxhM
zvHR0Grm3xn68TMHqrK0iQlcfUpSJJ0MQLzZqavw93sG3CgDwsbsgrBx6wPV9wEUfr+kazfbamQ6
iRFyIIhLzplL+lO7wKat/oAGdfwHGN/0n5AGcOouUwL1dXfyxt4/a8wL+ZuyAANHzUQ4l6DQgFd4
57mRUzLxFliYfVvjZ+Guw/BCjgRrC4icxSFouSsPIsfA34V4rdg5itdJh5E6ygkdWshdA1YIQLr2
vwa6OiXRquwwkv7gS3OBUuq0KIrXIVFr242mN4Esi+cMDIA1IpX28kF1VUdontRqA6xzRsGOnlwb
afbLxacv/C/zcYCK+HfIuqfW6RETs1wyQLDjrUl+P2loMsW3sQBym9RyTf7Q8fI46AbFaqhc9MfF
jHXmWPwB83vvl7Y0A8iZ6mq/TY2aDtLcZkf1DVdx5B6QFcW6I5vyU0UceMXE/rKM6f2bfAhnb6WL
iupoFRRjZ6ujCOqNCBx4KXUTe2NaBonhEdH7URNtBuA4HRaER/mmB6ZziOZ1z0KP7q0e7qYdXQ/w
plcaClCMzjSZrPmpEyahryqD96mVaxExuTqBCde8l9ba7AI5hInMs+g+qW5r11V2NJRAwbUl7h0g
w4YY8GWZ0PvHePzgB6yD6vSoJJThHSM8h2p+bhiEyFZH+/U7fxZg6a5k1eHR1ExBMtSUotvoG+1z
pClP1Onr5LWdbhPACon9T4Sw8bKfeIz+8C5vXrq3qP8xbzi+dJ+zl7WSon3Nagc825EGKEm4ors0
P5dYbw0BCf/Us687aoF4GqmnDPJJhiKznPx+tx250boR5MY2+143zFez7fWZdv/Z0ETivrq0EErF
fqurPBFLJzFEkatX+p0IVObvx56LOhBypuePmfidCJaY5vzcsaxbJcWnPuM0B7q5Y8Lz0kynYzTK
DYQLcvdTeW6X0Z5HvkXsy91Fv++SO4cLzFDsUU43juRW9tETKfurEDbm6Nb+8ohLMycz60+s+nv8
2dWRiFHL40YiVwYVQSxuod7UWqycDGYegFW1XIqAAZ90uVt/xFaTsvE/jt6fTiyfecJB60pZtTub
ViVdhkawJtNdmyNkzMv/HmB4WzhrvzWi7+ofFLTxWljMeGVvHz67zmRCJ5ngcqlMsdaOsZRTa6h4
KKMl9T/tJ2svDjcSVLRZ88RJDpA83hGlzOcfyf4sQby2220Vm/h20H1+O0G0iVqR2DAzDf12YX/i
qbum0L/JThG5JLbEIW+msvqWeZqZ/RpQUOXDlCe7koO/7RXtVuXZ6g8qSgaApxHcpFdVO6EaxMq8
PHxfqsw/iubFVefX68tgbuJ8nilWYwYk4Sa4ukMun5+v3kARemiE9BpzslXxzFDCX4lcoqenEIo5
DgTAmHXkyY9LZ/r9L26d0w+FsBDlW39V7Rwmg4BW1cRJKux4lmw+/a4ZFkLrcz+2sQBIsjLc/idw
fpZzk/xMiRHHHu8gSiY6fxqIlz+I8ebQNFDStMuTE9gl8dXeOfF06tYYm1R/RXSlUsfY8kbwlXVf
DuAejuMUgDU1P9PWPvFm5+I2YLXmpTbW8hftp4AXAyK80edETqUSGxdOT1dZ3iKny57IWLQRCFDo
6GOeMGb04FZEh926vryqHytNeATis/y6DOWP5fHfcmzhYb/50ISCMADtiPwi48hBjG8yi3AtfhLb
Y1+yA6NdSxcqROWyd5HiBB/n6rG0Pa2wG1cwc3Kb3/QMhpRgZUymcAM/fchwzBm1/JSUyGt02LuZ
ih8mbVwap7EcjGm7dOvpe64XUCuj4rG2URumgqAvnfQzFZWSqb4fzH8LJWfFU50JWIvEkq5exTIh
0EDOVaW1q6ACfSnvco2klTvz3BRM894854T2OOUhgRTYkC57qM5KEzyi8JG2UyUDudG3rOfDLPKd
hmhrc/IbEkUzv9OW5NJoqtjFcrxwYkinrC4G+P6lY9CELc9BskMBm1A8VjsCCnPI84yAzPyXQM3A
N5nuA3T74BjtogThDc6FsgkHkN2y4Truvhfr0EeWAqhdTVMoljttjIws3K2yltGlX6MBCr+UvT8N
qixq4RuNcLZqSSxE+TGkM6/2LqAE5kZFdOTdD7aDnnMkewCx1ZiJLBZl43y2p3uy2PcQ99j5cnnK
gHqOTSXgRcaoW//n2tnr7d/2ouvrVim2zzSJaFvsV29p1m4DjEkoCWfSO6HzsnhxwagfOyw9WWoU
UIOuiGei1S3ircvWZR+B7zN5OC+RGTz9b4431Fmmfq1IHiayjf0bFUrruiMD3s/4tTKsrnTFbY4O
jq8dKQC5EwC9tYK5wJVZtzDhX/3LaG76Q7tnW8DTOFmcnhLwGl/sRzKSlO9PwH6fZW5P8fgFHM4z
O8qZ4BslIB9OCQsIneEx0DV/R2Y74Ou/jXQk0UzW1DGmYZ5mnfZ4b2pnJxophKyrYRkdkSqXMdy8
ZgnDvm2X9ZM9aVDNwCIL9P7F+WFq3uVnH8GhAPYHuRYGX/z0p9t3tPLPHjNsADhxFHk36vxpwSgB
+xWVoCLExKwp/qh0qg3xDqfWmMQOf24nfiEbajnIeCAiiYa0qBVqI3yqATcIhWY2Fi3PCIp/A0n4
Ry/U9ny2AagAf0vZ6Wi1ULPEtoMZji9t8YOtSdJQm52W+OQb7kpkfCHf/ZQICixTup7xnCfR+ow4
Zya3pYVHjnyOmbMhUx34Z39Bl5QiNZoKV+TZ9Ct1WlhbYltfY/F6IJCiFbe17JhTv4N4KVIbwz2a
ZmnL63M8pQH0FiNcBBWFRO4x3k36oSHlqiVj5XfzpgWFGe1sLI+iAgYGJpkMnZNeLLTjtccgVuBg
hUftZHFwLK/BCrlgdsDXXMnmjIfUjiNPlAo8GXMfPU6RnziDw15UTRRkGn8K9wMqIGhXq++UfYBN
0/Gr4/wMp7tK5db/Qku0GgeBtGmCOQYjOiXp9d0N1/CDL8sj5sGV+VENqElOX/1LsgXIoIWd9EZ0
xETaZNKgf2QhEjrYfsQDr3zXoPCTy9TafmvSQ0WXlE5yG6PfR4f3WawAALMmCFlqSHTNdY0GLgNA
30FqUtbc28WPSxrXRKjbqLFwjWwtaawc88MFU4+S1wwMCwv0yPXqwvH9yfDYZ3I8qxk4J4LyXAk5
rwsAeFuH0q4EDRPJQEGqX+zXCE/RIEAsifQcX7hpGsu877oh7a9plPmIvRp2eHQmJcY2d4k/AC8o
W4kPHiJwg6yJOKU6otnIRX4jPXYP8xa9wfU2vpNjDdjE5rq0yOiD2nIt6PWeXn77qrXAlvhpMWJ6
ApnE2BdOp8N4NScw1AhSODW0kgd+mb4Hxo4Qb0IKG40Vcx7EoAvkicMCmv7FJyRe3cn4b4KbQnVY
tZYMxK2QaX/rbAsgKnxHPls8zeAWBQdC9f+3j8mX4pBlLTW6opUjceY3sbvmmqVOiypKBMNv46S4
RgObNiTWgG+wFI9CTxzb3S/tW7hubyQFqwsuH+Hr7g7Ljs3kbPnZ9XGUBbxoftxRmNuhUZ6UqCQR
alhRLZMRr7ZcuRatKyeyNbEF8P2Xm2dxTzkvxcMz4HkxQQUsnu++jDcvlvaMAf9dSOGykZbnsbjN
gMQIRsRV8euz0Bhbvz/oBjq3sjuPJHZFZVOJ34YI5af7coR825X7c4UM7nQkm4tJISpC7ohJnig2
VP70ylx/vD6S+zUNdg4eEpqe8EMLNa2u04y6zB3ihJnWwYVoNylv59TeF12CYMGasBXT2XRKAxvy
sqHC6Q6F5OCi6yx7baG9nTMAWfz/wuN3O8V/EWI8FHMKkStHz9brojP8fbX/CdCMrZHNyVs8el59
lssymVyWcExgxK7qamnrYbV2l4C4p2ooOgREMrpWw2bdYhcA9oNm/HIj5CtXlJsDBolLoY2KaHk5
GAIh8hFlQSPZjNafwLbPWJEjWp8akdaA7vwgACpqOiBUUVcU8eACXB2X3OJmuIAvJpyoIu1YiAza
jkZJiJ62Xj/NuhW8TcG8Poi5thz4fyHzVMiyg+xHSzQrrzo4YgxjINKYbD0/hrz1nM49yT2arS4h
n6RlsPsOV8qjAhu4IRPalOu3sy1zA4J/YC/tIvkbbwbBlm42z7yujENVqcRjZycitaaHgPmqgi57
a//ZCbvE4adeQ6cEZwuqH9nydFsIeQAeaNnOe0avHUO08rHUr71TdmQ6wLBns65BaNqC8316NYqY
5AWlOYtJVcC3PvDtZkCynFVmXF0d0gzhhjjkEh37JkLR0yl2Q3VeaXKMI0+JM+n9RuZ2nAXabJZC
BS/lWw9RPAarJRRaZ2mMbFIGB0PplxR4klg4iSms7fywp467z7J3NVSwga8RhLf7CLcHZXIn2JwP
AUaTcbMa6N6wl/vFrDwKdGIenGc5+yYBAMiCtCXMEYKuMd1+J72h09cvXxyfCvCt2mRvC8ulQ0P5
0TkOFsgosr0CNs2SsPtRoMsoTvjPSYViCq3fdMSB2ogygdB2S/WH+2NGAD4aaSdbJ6byX9IzRtBZ
LbWa7lgX8N+KEV87cPcvO7jBbJ/BHRnNTRm++Mdt0bk/NgAEy3prK1gpiPs301HyR6H4KWdX6Ljn
b+UiI+tKCljvsrzjlOfEa2+/57Muas+bQsePbQ5OlLDA/0DxjsExkOYVyPu87hlAPR119tIRDvjH
vOIIb6rJ0LHId/n0O3tAA99zs3ko/wD0Y8E6rObDSse2dStT0TYk/tZqEJOdRyha7EZnLEnKN+fC
V6c1r+YCheAh36htBwJ/D/bS/XKhcjaRZECKbk7noW6UbOOBLQO2Ftzr16E/3e9tF9WkBzAuNBjp
CwhzqoccMF9VhZhS/xgKlTF+cmFKj/b6uECnPwzWY707a90kQkcaLrL7LdjrSQGzFi8BT3oCBiOa
/xUaQU2HUyKnksEKy5ed3hHgMNxSv43spKF95/OFL6kICOlZ3LPG7MyvFUsgyc2+405kVw+SZeoc
N+Oy/dMKPDHw4jTj+0RmkHbaA7wnqKp9ERsh4voCa4INHcgj06JRYj2j1Jrg+lIGAit+ECle/gEK
Ko+6TqLcWeAeMst79lXZ2ZgDNhxHFjnm9cDQLdl86TTJAlfhA+jMtMBAcUJVAmnzmwdYAn2PtJn/
Mha1386XB5BktTNhd7rpEwPWQ4qFxyqgp7x6qnTJSAePcQLaXlwr4au1LnJhj2jzsdtFAx8gzImU
HBfiCkj3fNtV3S6wmRqKUUCX9TM2xm+V56aVAG6rmUNvIN8gs0fLjVLVWDhpgmVAJ+IDNhcxKs3+
0SH+iCzkb+fstXoVENYGJzqFpvXEPzsGlCT7vfEZP6kg9LCk05xOkWDWjy4kIh7iBRp6C+KgH5jX
Mfne68qSFQcY1GlT1bZSQd/lGBtWz8eaJki/bZ+z1QSk8IqKPAXMJ+n2iLdSe3njBQGamsDlf/4r
0XN5S6EULO+egnlCZ55/aG4Pg03nTqoXghsDin7r9mVB8arpuTjxniLVbnDzhLWf6GnmyIROhGRS
q/3LNZtR60cYItLOeVeQzu3y4bjEvy/OSBXf1s/mbkWJcmvMZsdUH1jvExTrAQNfIi8AW3cnXeoR
9DytC2GoBu01R3b9NISXnwmNZYHHSQ853T0YnrdxN5/xdufXCMPNNRCRnRqkyacwr7WPWpjKnUSV
5PaFrLI6SsZfpZ/TQb6Qj8+BAXz0O2FowmVtuGlFawDT4KF/JrEf133Y9IrMxeIFvyCn9C/5YL0E
Bkq8uDf5MwwUYgSS6m+MF/uxa5T+xd6+f96TyQfBV3FeYMFqeM5Dde0Ly2w5aC8Ane0QQj21qfOY
Qp7g1Tia4HMljIBxCoi1ST+pXdVtT4+duNG6+WQ1WvpLFk3GJCV0gXDH5HNUpJaW4d+4JP8EKDF6
fLU6K+lKtyX9/FVyp3L/JPsFKdL2cbfyqkKzGeJWC4RADFRwsdpCxan5tOb81u5285BD8XpVl5uD
bztQ6x5l8eSeDnrEjC9LAEFQDrtwPPW2OV4rEVkQ/nfl6OxpWtX8Dg5givVovJ9Z7LROd81VplR2
n6ke8v406tr+h0WzrSTPQaBHV7LBD47EApM4JEZs3khxokJJYIlWE+TXv/BBLDic3fqpBAKN9g2T
zpXdBrXpBO0XSjD7XUiwfG7f0AhjMwrsJYnWNQGLXM2CTBoF45JXmbujuPdi4vyS7T+T6Qw8Z+iw
O6LTdbwc/MCHtg9g4CUTpPXFuC7nFRrWW/eI3JBofDLjUBVaG8c86SXSmQbWR5oBD/vuPCGTcAR6
tEJDJSyN1gCLbiEv1HQTJbkewDgx9I9O2xiUTsZbKMANmLI6cU+MtL+/nRovNn1Dfc8EJp4qJsbD
+tpbidKFoKzBIIlT7De2iLpYWvRygzj7Nf4QnTso4wzgyyQ3UM09o5CeJir6+8pIR4Wy2vyFWUUV
jlF5O/pHb3KxuTLNBBqTlTmLiPWM1yIw12komhg2CIXk+W2C3oDT2IZdLTcfexAt+UdBLqJTS2nj
CmSVGqAfFb64L7/Hiuq5FtaZ4ka26RLeyeE+InlHLgOSVsoj4udSp/pPWsleZC2/E+SP7PYFgfFP
4k2JfOqS/Pqnuw9jE7LQIl4adHcG/iIxC2ZGXwLCnjDsCX1E7Dsx2pszgz8kGhNktWX66QM4SBU6
AN0jJsaquQcecWzw6j1KLnzqCiXcSYxdY3ICOf1CZGNHBQ6OoYTAkx07KBaUet0Knr+H556g9sCt
oCL1Wv23TgIAyi5flGF6t8+FWYhX+u6ViYWO6Ew+Z9TKowNReHCvccjliI5u4nRZgDIPlccV6rbG
rDg4G1Fe9WckMhON8p4dwiI0nGIw86WZ6mxInY3fWFjfqw9uOg0jWKwkEnbD58sPipwEqpcnf+e/
U4LAr8larTBNyusduXjSRAowQDXeVXgpXZSYCkmlngcXzZbJEdydVmAwT978dExxOdU7UZhYmxgJ
gFiCZRlrBoVrFaaquZdh6bf2sJB6MdUa+nURbgCI4yvDv/crz/7aQYHlwq4hPulv8erQPfMhpiFL
rmtzn+/nzbpAq6pU9TiyEaWoHWsKwYBRRDhmC70IhHGqGgETNNEo1cpa95CSOFulK3piQt0wFEf6
+wORw6eMzn1bdKpOmn6xBUEmM/zc6Pn01iMSbpjxgtYEKHvRG0D6YGCE3uEUPpoYryQiwxgjZKpj
ijZTsAGP1Aufea9BjAFicXBhMZo2cxQMcBajjucQ1NfE3MrzJgpZARFj3D3f4FMNS/v02iv7GJ2w
mP2mzXGx5gNmQ16QcVRopsdhQ8GTJSTMiaPCo6N/Q0IKnXhxv/12KQbZuEAORtJ0MZo0Mwbi2OZ8
Y3qmSfDixtZMt5Cpwj+XOGc3CV5l4aKUFW7MALAHfdXx60LF9RZ+dzYD+iOp9ToaR21DF5s6H4Dd
GsNdmjxDyuQVxueNmyEcwpA0HZ5JFYv+jBSZigKDEqVqgR/UOPrbXOxWJ0ldOBAOBIc1g+RBpnTn
5KeUm4WWhciCm2n0+x/XxY9DSeMaI7rhOnMduLrMm7MNwlboEvTaiYFWGC7sV09sGtENepz176Na
MG2p5KCwsMZZZtOv4Us7Y/m6pfylcA3HoquWda/A1Dt5khmRluywtu/UoOkbZT4gzJ3Btzv3wyq3
TPQFeCBWvKLybLrDO6V2QqroUxukyw0LEcpOapLQLm/LfNMaAveaaJRjfj+y679M7F6Rbh4Ne0JO
pa2lBBeC7dlesGp1ZeMMwQ9yUYFuqv6Aq4Chc1SSNQ2rbsrLeqhTqN4JW/+RHiJi8op1O7Z9gafy
Ip5LtwxUmgCcZhg/iesGmsgrjTE+R1S/xw5yweQivuMOd77eAod5eWQFhkh9CGLiEtrdLCdXZG3f
CJfZI21Qn2mRv2IPrmPvOwomeKfB6jFYcofgPWlB2TfD4B/zTs9WeRu7TGlzRqPsRxOl3LoPhrAm
bNgklVY/j5qGCyUrj+rUi7FAIb1ZOJYQdK4O/m2R9DedPwfRnTKGPRW05DyOwaV7kMNoxPGbBtFS
ecEWV+p9HFJ9P7d8RGDOrXvUZ2y7YfpidEkH6HIpH5BMVN0/j/BqOLl0lE19KW8kc+aCypq4pISe
VmXg484ThmcMs4XniWCq/TC5RgCf6x3A9mmO9d5joDKlYeFaizo0Dq9llm55RTE/wC6NgI+0zzUr
SDOwcxyESlSiqcKITpSOWyoyWjPeCghPmuJt8e3sS8G3tTiJlNjKrGpXjOE+h8LjAi5Yw5ziMmyj
lwpqQbRWJJukze9Pqf6mPIi6K8jSHTI7gRmAawCopnYIAQVie2HIO65hLljtR1x5M45/EXFGcsoi
LWGMNrr6WjZqgDPmpThpKlceg1zWRY1OIlQT8P8YXeuRkYkX1RHcnd32vDWoQ79zRfix+JTTdfha
3Wo1l4pH22PphvPIyIs6j6/dxGGq1K7cLec0UnEMm8gvJn5RiwtxrCFq5a2Zqs+JrcpOITCAe126
++uc8ZHGQhzywNOuCYKOK1kt7AJkya/Wn6tpdDoQofsmnB7vBi0oPaFjyG0nu8fV3WqRaCEwyrXW
KsUbxRTp4qvOy/InkXRy1AwIhG01QWusiEpcpDoBXDGZQaarH7xQ32Ux4019v0xs9uWrcXBYmWGB
+EV5KLqu4b03PZIsSz2kd3jSg0FbVepQhZMQYFhq8BaWgCpKoi2lDoVABvDtg3G9Qzo1E6Vl2a/E
Nxl56Uo8jRZnTYkX3oykqcqoXa948WnStr9Y34H4RVb6gHPFHBS2dCY5Rq3VSKvYyvzAaVI4yvtV
MtyueVo41zMTXMfXQB9bN+t/ARHGTFmP23aDv14KO673LI8wvfOwFwzqkSV4Nwv8mg3CP4Rs2lmb
gL2KZtdfmj1biDKOh9LbLdvgiFmAubOrER11Nm05hPo/Zv6xOCNn/winfCKAMSOWhVEjvxA2puMH
+FKSh3mXhhMloiOkV5wlOrjKzAV5oJ1ooOpd5UjPKnqA1tcpOwHy00O7IxE6ssHhk1ZEm7nTArt0
bnHulH2TxEbI4KsRITCi8UoMyAmaC4dOE4Axrg3YRpmn0M+qBjEHWQVF8Xza4qmuIGImTrVmBsp1
JrTxCZjaRnHFiMKJ/jfwUIbcbHIi9nvIszu9Xes0dhD7EY3XYBfIiihlgH0Onj1jq98yPSocbbjw
rDAkEQpBKh9LeyF6Z5WVAG89RCgok1QGQP144f0vuc3ACRkVAQVkiJchZx7q5TFOP+CU4puih0zI
+BXPXPXSKr9lkmq6dc0D3gH9z6YxFuBu1R7jHI+BGsq9x6CsCOsfLScPgFugQD8kSf1v+7UWVIxL
7J3ln7jgNKYDUqQ6HFwlQgw85PllWymIa7ssBAzpw5ulEP6iw1ICA3QWEKCm/zo4aKEgjqXmTEDv
zLSbYd3QcdRSEHdPv7p7q12c33X5yESRi8/z6eIlFrN3CQefM6v6/KSVcvShRZfEE1Bz8e7CBNb4
7OjTEe8zc++fo7Zk17YTQeykW9mxnKQmI6yT4nazytWUxN1/b0Mzwsc191dWs/3nlLaH3OWqZJxH
/8MjVBtQ1F18+9c6+FTGTIWT7Ph/cPUZiuTlSyTfT6W8kVMOB/YU/Al5hArSKJvsJDSXCX2VscXF
nvPd7xRmKtGR1nIkytMU3W8FqxPxP+jZJ+mI4Y83nSnD4e/9FmKrR3TjCMS2T9FOVsct+iefst0F
5NQnN4ZHmmAV+AcW7E/7UmpQjcjvvz5yuJX3CpE0BaZPbTPdOQ8XGiSGAwGtWjCpFzbz80BXiTrg
eqas5VQlNuhh+9CWJ3ziSFlolNmi+xh3iwkiDR70+t/CbfhdkLO2UNbW46n3go7k/BmmslWqLDGR
xem/0ybc1Lx3PQ8SsEnO1bMHvoHRjg6gOllbjeDV8WeAGobkrgjhKLqky8+147JYP8FY0nU879i5
9NM1mLdhq0sFVAM8CoBbEFUKCkjZRZyuQVqggbOKYikdt+7kVS1R69uaxI/H/0LU6PywQ3HgA4hy
GKKLDWMw3fIBTd8ske7JRvgi/0q+ot8i405sKvpIAWFrs/ov1REocEaHKyp5yX3e4MrqFX5Qi1s4
VyQIVE2cNk4G5Cj3BEbmMUBwhuRLGkmkQOBsT5R1x3SLoiUI94moLZY6cVst/t5UCHhXVIvKRXII
pG3dh+EWckRcIrjTFRl4XYyh03CdMlD7EsTXy/4UvOnvZGZSLiKoWLrq+mQr1Ti3m55IQ+0+VGCG
mpT+0H7+77DDl36OZyAOTgyFiNJk/R9ZnhF09wqY7gh6w5x/FnJCH6rJD9jpzHAHA8O6riS0kGJb
fcdoD6CqFRZmvxGmzMC/YElHVclKoaLnT/Yhk+cI2kpovvgTvFry+GllBHhO8P/B2DQufOI+bIyj
Axg7Pq8AN+XPsWOEiFUW2m+UsB4QSOUDYmkArpFFBSrwwqq5BL5vVorm3XIC/bFIPuSIyyphICuC
YosoDRUZFygRSSWzNN9F4almUCeGn7VPu7SZx4ISvVDO
`protect end_protected
