-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
VAddELz64gtIetkxD68pdXsx4R6vHIL57Uo2DnV6IvcTPpaWA5kKnM4Q4+3hSrkN
2VWC0x8A9m42nulr4bqDBcrrrwQ8juOy1VTxW6Kvd4j4cVlimCp4Y7StFa/N+Jy/
dtNTlsYxwWbU2j9VT8qq7qZ7JsexLmPzfigJ90qRXyg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4810)

`protect DATA_BLOCK
v+wFg9U7/YCYtP2r+YV8IsUllq9OqQUo8AFvlOEZfZ1ok7/r8tNANp7ikaOa1QXZ
I6hbss5IVycoq0k0r43MDbo2Sq/8YHJ68IKkJRMM4/DIB3bMskKB4RfgvruZNzEk
5d5oP5hUdzTkYTdFiNW4XTla0Mez+1Ah2oOCu5Loha6YcZh91DCp1k5ukq4PfJpB
x48eOvMEy8U7GqQ3QtuNgnJ7xRGfYCLs9AnSEKnX+GXjw+Vay8Iat4HsO1+Ez5I2
t4+RUV+VB4eWmahMJ/gd4+cEu00sjNmHQBNGwX8jD8IRiTJFYQARaNOIJAooebvT
qG2DY+DCAZ+NRJ/g2Of5wJBaWcBIuKOx3gjW+Xd8TWMUA+BYAjSNyRZngvXwaaUd
2qrbmuFjrmL84IOiLl9a2ubS+UgNDBQY9qCCo+2zjFs7aaBEpQXzDtjZ4cL4TP/G
F2k2wbPCh87YLZVkuArrzlK562BdjyYjSRJa9sIE2p3myReWfVUQBCvtYyUrecZ5
0QaCqp4HpfF2+ezGCPzpTXi9nUD04e8h3HISPyPxPwRBbu7x2Vl+iJw54WULNYVs
QWUh9zqlufGZahBjTXSHOfztrb0spb6KB42ysA+uI89935MS+3z28fcvmjbuOqEW
nUNzHAwoObh7Doyw+LjAqSXUb9AYrT5eRG3oS2Xh+M/Zrb3jUDZOesCScYkIJ8lh
4BqdAJKinDzwqII0HsZebtzcXnwfQny++LPY9gYQKRPAi4UGbJ70qGzZe/yewT4H
do8VwK/mA4JAIo/t6VlQWuS4NRpVGRu6UsV9Ttj/sl0DIidZ+VZiCPPrtw44i3hI
Oag7uITNFlOFTZJrf6EOrn86KGkwl0GgwiuTk2TE0jhOUAZ7rHGj2dQEvUBtc0p4
vXpC3RXZyxBNa1OuH5rHN1AvBqRliK25GTvdh5UyyRXjQuIodbR9ncwQ6vU71cWR
/w6TXuk7xXos9NEI5AAPI2sWOqbg7ALmN5TBJQR2RspvThlLB3m/1yj+xl/6yURX
VI3JukCYJwll6odYT73Ls7Rb9vmYi+dR7Wf4h1u0U8M3GaYfw7uvr9TeUKgQPXJB
0iQa7UCPHrztiihvb+WwHI7DaqO63pa9CVPwiZmpF+Go/Cs8ld8kGK8swQV2RAKc
ETkhXuADqhKI06wFoFj5yE8shleXjg2gxqpzNzh/cxMkSDjatpdz8dVEma7UAuqK
GCZdl6L3JuYMvGr0+dxkHFfCL3YjTXHpBHRs3t1tQWfLJMlM0odg8KvLqYYZVCr5
ceTlF76GR/3Vly1qiCVLoRSf4UEUdX7sl/rxRii55z7UAP+Tdus3nS0rAs4SV7aI
DXH9mhi9GguXBrGdVyQlPtjh//9Gs7BwRKIsDf7SdWnN8wfz9X/SF/PCxW0J08P3
kzScHN/f4ErvNp4FwBtEXvZfJ83S2GlLiqEtLN2MQVxSZ2mdsfiDneUzPUKusxaI
N6uBuvhD/eHYN13uiqKxBE341GWobfBalEK9ujzLKeyLiGeRp7V4onw9uNqXj5YQ
qhWTMMoGbWsJxBbOYbHARWPSgt4fOqQ6CNZMzGFawDoQudichU31aWm1byYkMEaq
M4yEOYKno2NGFz3qs2d4npTQmuIo8kO9dVAILZy2FOHjKKld6ebY3NeX1j3GmlRx
ZfAwh4OS+sk/2Xul64GRexeiSWfzb0U8IlrpF4VwKlNZhsdq+9UzTWiU414HCfcV
W/4y3TdyseTGZrwcoJQdINubtgP/b42woaX5iekAWh9wP8BpKcDJ4o68gjVhW2Ad
uSu5ThnWwEZEYwKPNGhBZH4/7IDzeqNaMhFtX0W31kTNOMgxFWoJtgK2s8E/UoIS
fXS2JVyH/YN0L+A3GrS29dwmqIoP/P7iL7DU2f5maXhI7PnGphgij8XPufDWvmqw
MRKBuMlZTzpVRWd2Fpp/IpMh2hb2nIS0OJFZKEY1TNJ0q7UP/6L5rUnnKIhsa+zZ
/e29zpxxWw0SoRLCiWmfI4niAuXUM/x0kB6S4qgs/LnsKJNncNh3Izxk8kB7Mt62
1Pi6CIAyRuq8kAK3RkQ7d0Wvw3FdirJIJi16iEQa/mLBKlAtuJlWcG4dm2Lb8x/0
grj0UW2G7NoN15l5jh6ZBhbKACKYpLy+wuj5nQdC8tmadfSDqP9haC1FkMMI/N95
qSC+hrv3BbAEfFFskSfdXfeAFqueTAvF1htkdEqOuZlR822KOFlsQDrtxT26ZPLE
+BdUgVfxwLpyO9yHM36WrMq2PaQkvpKJnYfn56GZJ0NKs3/BqnBy2gpPpq7liSj/
IrS3U9mUJH22ay+3y0eBJJCvvZn1UJ7j3TOrEeKeOjxrfK6MOpCjpW8FfSy0TZdy
qrjMEN8VhBxq8fVM5ZtNpX7fxqMPYI7QUwY0Wy0nRT36s/V8NXO8tiAPC9bN4j48
81u2figFqwHnV9lcEaXG6Z795bshWjEtKO0fm4uT6tCzcjdvMhHcLiAsfyrmlhdM
QlXl8arqheMYxWcX1U4aEe+ZOUZLEzv+PtYy4HGgwhZqOVdze3FZDa66pFpk2fbw
EsbBbJmbFh2QwJvNc3jbmzLL/T2HCa76IggwZ5BGdB4gTEqAqvlJcHNQKnTfBws5
cEWnYJlf7fHBq0+4wpdeRdPcUiM2cVP9sdUxkC6cx1YV8JWXngvvUY8tXRnYtZbt
AQlkd+uq3fl8LReNhmqPC7cMQkTKYjej1NsdvjdI4TFq5fpBsaQUOCiD9SQWfl5e
UDGBSinI/BHCKAaXRi658oUkrfqway4VjM0kzZSPyXrE4X/6v327+WSGLSjG5cBI
jGJDld0ug0tOgJoV038y4W8ljBGTCG10vSx1JvTnFuXYCTNcoyafMI6ICpK5GlcQ
gk+utbLwLKypsFnpZUxmH1ystAgWpwXIT9Iy6XZiMwlwHwdBsw1K6JK3I9uFWAEc
pTv4qKM03fC7acqNIGz5axoDZod4j9kxxtvYYwwB5NaZEL37dhdx9O8n0h4AS8Ka
YbXLHeZ5SsT2e5AxAi2DkCknMUU/gq5aex5aLBDxtwzBYxyU9jS5Nww/lPc9bmyo
tyLwpb08u62yyaxu3tQxP6/HXSLCU2ZTo4GDGDRWjQOzpjxnkVQDuvXQhBJysQCs
J2ENb2GtcLI8tCF0dnGD1E3lrhgCTwFa21e3B6z7qDIT+0HWgODT5JR2++TCUWWw
f6WsUqeh5ezUW/MClHHjd0Z+V3sY0LDw2B4GMXzXNxSAH5pUnTe3CJBKhNkzmqVP
c2rO3gshpn1uiBGFwzQ4rvS7Bt6dEO9Ew5rVtvQtdE6rEjiQnKubgDvnYfliFSkd
j9NoNYdTBMQriLVSkdJPqShsPkAqSadwA7iKlKpwEM/TUSnnCdVHRGcDZWujC8+e
Rt4yKxQlJS1hYl703M8zaSHaWEldHcxkgLA3rh3GWaxZ5usrqna3K8oxh/V3A+m4
Q7Hj1f8P8ZxjVtPBWer4i6YZcEd++D8gH1cprcVF73+AG04KUiRtDrvrvBeZf2ZB
mDkZbH94mY649IRFT78zIokPx5fYtxG0LLQeeX5kCjSmOw04zeaMbeU7MH/0po6G
vgQhwroVIiLN1RPePOgviX9Ohr/ONlY6NkYzDb52khwR95V6Z4E+q3RB5m1IIsKA
tGKl6gjUHfa+nwc1Z4B/F4KNBFgiaVyU3wHFOF5VIpXxKnTFHHCh7jRqUVw2sGIp
zYzHEJLwbNcArtBmOUnweaHaJRlCv54UklTGe8Qgtym1E9vRCtNh8Qwg4oC6lTV0
dICajuzf4p1AAAChpkOtR58pA/eV9RihiwV7TAvW0rpxu26sWRY0Fbe12DsHivxI
HQC0uzb1phX6nTH4g7gAIC3YJR19QJjXdRfSGSuolqI3vVgTHfHxHfTz3oiW7k/5
bQ4HbOLKEm9CNGYwr0tgJ32XUrQr6WRIJXL8YGguX9WM3FgYWx4cIk3bO+I4a3jc
ylXG+fq3O5154QyYAqnOElOjTT2anCqAXC0PlcisrtWprwiq3+Vr2Gc9p6vZZEtF
eF1SMORn/JD8E/bd1UN1GkZ8b/nnNoaucCo6pVDoaLS4ozDd3WBbCMnE14z+jMXJ
bJfWCpx4a6SofZSUmbHSfRtgjhrOBHiyDcNw9SGqlUs4nNyjtlOAsniTVxulFTpC
tAo1NGcquO9h9e3fKmmuAzrIObXC70CshfA3BF141LHmPeVw0DkLAZ0QVTQWr9aB
3aSA2EvtMVt7yLepRDmyVvEd8bD3yyHnZ421sveZiWPn2M5ThLJtrbSgp68NRrxV
WIz22IAHjBZlLpHzO4mfXUv0L8thGIKrTP4Qk8JeTXMqR40rUf+BIlmSTOGKQTBS
eewmFC58nhNtMHNGja88IOfFUAkUXqx+B7JHfbmBuubS5e1ojm4ov5BGQNusiMGq
W11MeG+Jp+mVgYCSxyQqQ2IrRaQpDS66UiCyMWMrOqve5iVtb/e0RYVsCrZAZhyk
5ovv+O3BSYN/aYPy61cPvlxiGal6h6MQj5ABW7jstnTInDRo4QtoJTaz3RLBrejp
DlY8/DgMUhHa2iFr+7yLeOTMIA8Cg5dif1MWLs0U7KA2GCheG/wI5aaCznSvz5Fg
39YtWboH37hCISyo0cZK1SRuWIGVjk1M7RiipRaCaqZehZND89NopoeBLBOTT8WX
NrmPehaman5uA2lZvZihB1xXVXOteoe1jeM+EZnxyUbM6wdQYuX6EF2O3nRKKmrP
DNNWwfgNZ9y8gXYsQDrHnZeaGEyZ3Zh7rkWb+DG1LtC8GdksF6EFz9N4HzwIumO+
FZhOIZDgVVV2ZksAaQp0/I+F8eECPZLsAdIh9ghhQ3zqWLsCxEMqlqkKI23Q2GKj
FIIr7quB5mib8IvQDcB5n/lB0OUNhf2tx8r1j/31xYOZe1PmXNIU7uOrfVPKL4MF
f1K3tGQ5GM0R1cIw/4tiHizG2pO6zHU06D+DRmyYUO4y7ZpGxnkAacmn2fGKoAOm
S7HO/xvMepgCofrF6tQ54XTyDCPFSoe85FzGSL7pdguGAjpzrk0r72bXoaGKEM8P
RRwqF8BCDLTaaT157RFd89aBs3qJBmOQfl9Z6U/VI4kzGeOhdmgMAxKmYTXdBSYO
ZSlaDZmUtlD1RtVdOxfhklKv0eOIEmc10EihIoTwFwZWxJO8Bv6goaS+lLpzIHXQ
Ju0ELiehfuF/gwL/FpgKawaikn2zHFaqz7vwqPvhPMFpJdNz77wlv7wKRFH/vFnF
lDLPGaa2PQ/911qul6BBY7WT2UI8ySndpjE8KB/eZ9xrjbj/15T7HLpjrjKb3ev1
Yy6i0UQULvftpLjuIDvIo3joyXQZrpj8bpN75cskLIL+SaATYHjc2wvXUhPHkNdi
3qkyziVVgXbBMqmhoco6XAj+GGjdcXJLzACr+VavyDHdvcGL128WE+CxB9tE7Obg
KUG3PIUe7itUSZnaoUFvMgaNb/ZlX/3S5w8RYIW2b7PGpxkNPa2l+ViT93wZHq8s
cMjjk2xjFtFwIwAEWiVK42UbPs0WzbQ/GnNuBt+tsoZ9V+tyl4gGln9v7bi+fkHl
tlaTGB3LIidzRK1eJNtSl63PA5zRn6i7G8bX26YGIhbJTR0E+O3huSGxzlBBN6Tm
r6oZdiywvsQrpHSLRCjfZnhq5MKFRA0l9GgPBCkXRkVTk3wP053UBaslx04NGvMo
N7Svnb+i/X0GuGaUfLmw8f+wTZYq5kBaooZyunxUvORIBtDi6s/mYwmlVE0g9gpr
I7eBSSORRM2MH4eHSFbjz1GVerMgLULFLuL11/xLBQH1aBINoVMazpj3Xa22UHWn
i9gjNUPa2+2QRc4dAXv62yxFlJDgfkH+wGUg56T18zzvel387aTDpS2SO+7DY2c5
+iXV72uRSXJehpN5cds7RGk1maZkULgRwmPnL4IajIqb/jdLK1G26rMky6Daxr9h
SsSjMSZmLu4e1Ng0fFuboJ9sRjBLy/o25KPVqH2f2VBkSQTFl82pWYLFjEOtNaK1
kT/iOgwXpJvazDAEL+i0082viEy6jD0Ds/g5oYV2g7qezqmRuw5WZKWotvLGUjoi
Fz2z4yqiCtrERnOaAO/YH0Qgg/A7xA2Udkxml260eP6u8pdP9NZYGnjrFBh6MhJL
gD2sVyGZwARNrMVlSkvhh8ViMyNNQVpHCXIlVjuzwpM5/UPGT+SW41i+KTNOr7LC
CGqtH8cI3bvYI0R22l9IFV9I+Hv93PBdY8Ujq3hYQjL/oaLm1wqDcnnhApfhKyCx
qBAiwK0IIvBeFmD3VJwgRL1qSfkSe+/+e7uLc34NCngrHG7JkSXD3RP+8vOMWU9N
rmoXwfP38QzoHjXt5J4HcqEHdTiQaAB/qkdw22nJN9EVnHOEh4MNqSayM3J25Y3U
4VW+nn8mGB5J6dWRhEal94Gx85KJQgtdNON7AWFYxPE=
`protect END_PROTECTED