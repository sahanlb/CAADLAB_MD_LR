-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
gvmIYhcG73epdlZtGN1H4hHAwwo+44zPs63QPTdQ13lYuBJ6hYGVaev4ZCWUSJIe
MuQ4pPMmwgJzYSQICMVohh666xTarmpmEIT8tVwllYho8ovhJ42BMldsiB6NDSHA
gPYhkbjbtmw+sCmo2+rrYo+sHQ6NG79K8nv4xNBDjI4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6880)
`protect data_block
erNiwkwdqKwMH/OCV6ST/9s1UsBQUIVYaXEIP7fsSiOO44SsyCfOHVlnkK8pCrzY
5Y8UzQeck8fWJangcv4I4gwJYGdvB4Pax6NIDyCyjNbRpZpX0U2hOSsfKO/uZMu1
dDLcldz+3XhGZdTgNiUIImeTY7f69eQfcs3PdBO9Xbhkk2ljnNo0dZ/djYT1QnrB
w/GgB4GRetK9ugMBxNxBFMaiaQx7ntt1uXCSY1M3m2k/2D3wfn+3H4yDPio7lhAk
B1iwnSa0F9xN5IOPq/IJ68K2hc/cQo/J2uubeR9hnj5HYIEmCkDNbkAsGH7d1dRf
uUljpnsCeG7e/071ohdrQqGKFSh0c63xgipEjnhTVxgB3/s8CtpAZDZGBq4bRmZC
8jYUHr2aELYAqxDARWXE9K1qhuM/dVI/mTBxV4LSmsi/fW44FI+ij2DygctIe/XK
4I0G5MTzPSo0uUTsS3hT9FigRJGmV+bSAZTVBqnIaCWmAhCQdN3xlkIyXN2aVila
AL9uTovjCYIcm3mgTDXDyZzVJLafQyNXZXxTiFQfTNMuGQODJZ+gZJQhVpqqWLHV
a83Nj2P1uIbdRE2a1WyKm/sDn59h0yzWefl6taTaqvJpMDrSaO9BoCWeCcDScqh0
NFXvoI+3khV22gMzPYm0vBnaX+dGn0/Su5tHer+91c3Co2dbowThz3GcNE+6lUFs
jrZHPvpD840t+zm/1EcWyjkrx6TEwrIRXwGh1E0Sbn7Yj5YCmyUlb9ldHWcg4bVl
wvBRCB/uNQK4K5L291a2Yv68A7Sb50fFjvpTHV30xPvwv0F9HLVPVDKLm01xd7xM
908Lil9UJFqgz45Ibs4THKh3yyfbzrGuqVz/6sca4hSrWJpqzFQa1V3bw8BTg0sT
hRoJ9ipAMET/cMFT/fgH5mJertJ77jqEILiFBEZGbc2LuAmSsTnNPeov50Pubh45
pxzTlk2Poq9cHJiX7vaUUclOvcEK/6alIBfgVMuGNrj7c+LWxBu4qR/y3XeqZonP
gzCnsBWbGflnph5qyCpM2tN/Xf75USp1eXSfAvxd9L1Yak6bz0LPhaIXz31IlP4e
VOCwi1q7msX/WfZyHRuhDnPUBOPyhh3JIuR8K56RC3eIGqPSAlZL30GvqCn1cngQ
6R/HxuYxTbv9SBvjWp0DsYv/lGU0/M1HZJfei2FX/TcnPP9ziMjmHyQ7LRaLWGmL
37G6/nXrj6QkdfxsRrrJ7OHkAdGQRZd0NxkLf4q7LAH3s0i0qC5D0a1aKyQPzpYv
ubMOIf3M7OK4GgVAZ7cqfwUJB8TzP0XgNhaLWo7KVidkUIAXEaZH6f5uOYP4s8GO
h7vz8BPqTgmW5urwoglFyi3IYYY0fBaPkj5ozdG4u1pRuP31h+MM6s6KA1CxiENU
4prccL0KMDM0H+y5WXhRvegJiDdYwWLOwvHXW+hBZ2EMk6vsMKUJmdM7sRGGiIsl
y66gUbtO3C0vS+RPTLj4vNKuzXq4fQwJ8bM/AAqmKY5nbkM1Ja5U2YhaFTKWsHCZ
wi61ZxbqpqFv+sYp1AaRheOZW7w7ISadgfVoJN1GJRTjH3WzRL5Kk92V3C/IkQYz
e7n9wKiugNrkLIdfssekI1ptXm4npRRMnJUAiZvseiVXcfm0O6nfz5fTP86PchS0
pIgYfnQM55j35Kdx1HV8ZsGmmBu8zaOezH08C/OhK25pEteYfI3mPgWR+9936yPx
zB/uNtQWbMQF2YfbPIOXn58NemoSGg91HbAZaz+J1CulfXSjDOFSXCGlgCtsZy5r
x6lqIOwIhysIOXyzZ/QN1BchRIDgul29LS6xcp/TZUkyDVlvY0u6cBt8F22xfoHk
VPfQ6aQ8fYsjZpgs77MjaTJKhLXeasAQ1VkBezYWvxrWLK6YbGvFDnTVrQZmLI+Z
FPHK6iZVpylXsTHiP9x03gVyRz17mNpqkdq3+MsjYqI8NrRLIuLh/8ECz3/0hVSw
85BEaiZIcmQP70HwT9FTll5XdUHqix+v4SB7Y1DTxLjItgr8EAvyNbQGELIrr5cA
EbjGvYjB6PZCPFFzCvcqRGE5XuSUJUJQnruLSjdbCbXnXgxGwTcQ1rwLMFJthxm6
xU1imM3aQqZ8RMrnfvb+fl36kerayBZ/StfZkopjm/iPE4ab9+ZUX53lVmv8E3B3
ZF0l/YF4vMsnuw8NbKX6EWqkVRYPW59ReqQS21yyYxdVXnoa9z5dBpFkmFqZSXJ1
VPzj8ETpNjWNqriQfYfiM7wd5Csfz6BePatFzm+tOX05oSyM00NWbSG5vkcAlTDI
Yc4gsgsIBDNCg2AXpHvWSU+VB1cY2LLBBpiOeQRz9V6JiTr+xnSB/Yg9I71Hsgw/
Oc59ZRDizuDVZMwns/vM6wNSHNEJ69NFtrDe+AIElqsJbNySm2bpv44doFYBQaCA
XUliMFc/F67iNGEb/fTvhdBGMCeQQgCmcgvZlZT+pr/tXKXvVYS/lMIBmmjthuvC
Kd+wvg5nkhfGitFFEbUCsFKQevxDVABYlItLGpFSM00oiY5JX8mJD4pKNAEvehOu
yjgUm/0Nj/ktG/L4jJ7YZ1l2ewtZWE3ifRaObSlbTiPuIj4FumSXHM7xPZlycizX
I5c/VvuZcXkx9V5C2ifJluhKRyaTfvzIECXkCLOgvSjOZ02lgibkIsHpcvD0MAB+
ubuXFDG1aoKCVFFZ38QgHf/Q4cYCqnTmZc2idn1OoNAsBzewUWMnChUmlqpXUvEr
MX+UpuG09P4QM3BVB70W+WZrqFB0+nGoNReqLfU3oqxofTZ/49oVmAyeKbCWjmJu
TEGdO0ysGmcgskie7ng0+nbUKHUy2ZJv5dCBj2mxxthLKWqTbx1NAqtWkBdSscvI
7ZcuV5ViypvrCH8dnKG5aGRCDTpo/xqEJhPHAflOffl9OHvhBLQ10WJzeK3/ji+M
/F654adl80aMIJ5cp4XQSAQFyfn58OqnhR6hmyAtwslweaL8yUf1yr0/KcO8+hXO
30RPGfKjc2ghjBVvwscoobTfEyKdakJ3TLyjBGjss9zxCt6BT8fixMU7JeHRhGoo
kQJ/pUBdSHaLCEDEcVRnEJyLolUlQkAdssuC1FHmJPSmU9Ebs4vSCM22NlO/DNjf
ixggINB5WcQ6gKRVCosp6N7zZ22sCPlzkT4EhoU3ooXdvYboF9pNZkM+0ilfUa1r
5YGrAvsjXKw/iH3V3rtEnjKS6O9MDMVWOG1a4XTZLPwn6OgHGkK9xXW14bTjIzoP
Jk+r9OAcBAi0CiOcC68vAS2FcIKqtyiv9D4ql87O/0q7mAaJJlj1DQwt6lFQ9NRS
YB0jMxCDmFiMpRlwafF30wQ4uOTmokodc0PfK1MP2SE5QxcmIpgiF8IP/yAlcFuE
+jpseCjBbexNDaY6/k3LE0Y0yoeLZXq6KvLuYUI6NJAiz7B6fQ4+WX9rjcCHIbTv
DTZn5GVD91zIXUo2QNzmxPJDCGQ+Bz5vbFP2PeX2IttyF+E3G4O2kdD6FS7Cxaog
t45j3X8H6IFulK/3fOmfRQ2hXgzpj2kmCEIqIdD9BHIOgYOlnMHsK1eYFFllF8JI
QB6uEm4WEhwbJG6LxO+ZGMk6FvJ/RRutD2OSVQfH7QaW7me7sceB3uObyuuomzmq
2gBc7Lynggmv7InrRio+raWtYDbV5JQDN8zyGtY49b8CMCFPZffkBgf3OLp4FxZM
28ofmPb3jrpZILWWq3YvL5qZA7j4yWbF1rlLvMEaMQ/WPJjuTWt1zpqxIud34i4C
hv1t3jCc4Np69X9wDnD3fbZhActeRIHJ991yVert/vflQANqeweX9WpqW4STcbKr
KYJW0dSJTe4cyEb8HSW62KwWAnHRLwejCBIUw+rXddZRHRYIxs2GYQQ3+51DPVj6
/6CXjQkNlRBWxggxzgFkNObpIi6bUBa46fyQ3TcwNHOaPb0xP0hrG2dOn9LI+hsK
DKndQRKBt5adzl03ZDsQP/NtavMlxPT4wIecDFunK6lLNN9wwIF1P7+bC3JMi6f+
qRh0wWQDinUFW+/+UhphpvZc5g7K3NCVVAmQvfkGnHrTP05oIl1CjHOAp/ckpwBY
oFjk/esPyp0NKTgfYgs71tgzo5Um12WlXOlCrGUJUrzRMNFfNRKftdfsK7wBK22v
ODjnRhrLLhkqLU3mp3+Dx1ptS/McFhN0r/hoh+qgDqmLIFp+VQm+NW6ah7AsVu/s
xuFe3LDJQ5ZUlsV8SwuofOBEsktNCNbxoPBnJs5YmjwAhTbmrzKj2nO86X1G1tEk
NVB1dTMJ4/Mc1+cnw/IeIAQk+8vbJdABAh0wMIPaNiSusFvmrQToI0IRRI9cg1lD
DsWvfd9+QYFmtmUL8xzduuNrkOVv3K8MMRqIn4mrfm5fDcQEDqMkK6HupsN0ShfK
635inryPd3eTv7+2MHfAZKzDlO7i+dtng64dAET6GtgQa6EtaXr6qra9ThbubM6V
jNtCzCwhcuSISWY0MabQEpZIplb1Dx8izNRNxVxA0vdM1Dt8tufBL1ktHKbaPkCn
xThoF6O1Ysf7PUbyaZt+waSpsIZzp3YZLmyReszw0PuwuV4D5rkwFwbzXjPgs3fA
tyophQapOuKRtadaEPGW6imudjU2xHNgtvKmZmoNDQAsUDmo/AEnflENI5bWoBRP
Ls/uRaOdrAvj9XcvkDe995a6iXfj2vOviGDq2RjiILOJOqfurSDs1PajNALVPnso
MpBtdb4v0+0pYDPW+HiaQpQ1UR0MBShMoEgiiAA1Q5zDYCs/zPIL+sY6TTK5Fzpj
fuR7/QqPzEsViZ/QCL1EGDBMeKATOD0Ew5VF1CCHo9plTw/LbkpSO0TsFfRz3S7Q
ozRxcMISWKJNAKQ9cPzsyYQlQmdQKwpGkTq5/b4BhFeniFc/vAWea8vm9FSO1qyT
A6jTvqGaAfAcwqA/kp4MXMnbaR5uI5TVL1C5Xfucf1rgtaak0/FfAszC6IpKyNB7
n/Y5SaL9ZpmraKSLANKWGAGYZwwZgCMy2CrSSDIeEhExQDOncGzgPBCc4aemXrtX
pJtF4UHhrFqiuTyhq4xxMwyfwilpi4eWPWgT1TkmrtI8RdpHz/JDJs9L19l/o5Uh
eBo7x5+c1J/qsVaazgZGVskygY552x1GUR/I3TdoIc/0tV4xHqsR3aPZNSaKfVqn
ed12W6sh9wbrcjolUTAzpAsrrkhD4hPLxOkfUi8zi8R4uDd5IWeEKcY0OjOseeSR
4lkzT21LIOHocHEsIJKUGvrynmYKVZnm4dBMI2fX3xuZmNAbOWEaJnC89huVEbvQ
+vDL4XAefjSY1lCoqMf+tDnjH2EeGOxRIyGP19RbzPvyySpKi2ZF5E0qqptKPtHM
eW3pN+o03iHRurZb5WWSVTpghBsafvlP407H+18/94NcO5E+Cpe+/rUg6D/TOji2
njFC9t8rVckgGMjO19oixypjeqX+d9HyveXwv/8KoeAJMN7MzcvpHYDrHn0Rqo+B
FSBg8b50wZDW0U0r0RZ1HFhMr2+7op5DdoB5IPYKHUKpqIhV572ArT3mXfWQpGF4
cLgHpb4TrQXFYtELPyBOOC+BUcR9tiKtvzcuh/i9Ie2/gXBAvL0fZo89YzlAdho8
Gj6zorSPdNaJMYk0n7CvMDX5BgzJwcyLVhb+RT7C0YRKVZWQWKmi5Oy6IIPpOCtI
iKu5ONQM5tU8SjUJCnoly+ZjrBKsVeQwp4rov9jVQvPbFPcQp0q7YymtfqY+ZSre
CowHIgDNaD+EhoMSIVrmuJhEV+FZ0xkptaAf89zPsUOyebkH7JSUSFp6hLejmPxm
y2OLWXjSyE59qYNhkb/AL1UoeU+LPbZqiSGcjyc5B0gL35XM270ukbujSSBLEdYk
CXrXeqdgNQRZuDEJ8NsHUT8QbNVFdn+ByKUQzay8WckEaEx16xtmlJgTtZ3B/6OJ
Q09ILPyZ9T1x7sM74RY49oo//s2QTbWbmB3Bpy2uuwfA5dKZpOoByaPFvB/Ptsp0
PDBuxADiqkhBQkh+wSig6X2Vk7RHkjVDJ+ZIum6ika2u49x3ZybcfdlAoJ6C0FE7
8NccBj7xMJOkVq2QceWB/k76FjdAunpOTWK4MEtwyMp21FJLrYGTSt04lYnWWEdk
cKLGN+6IhUBcNwTuxMNVgdvKeb7B21eEAMhqbIgI/in6gZL/Wan+KflTTUBlgBAl
1suyUOb9lXk5LUByP89hqQNMbs+hFLKtsaAK/p/drTaQEWuxbFsbZY8/AmzrgPAQ
gx44YER1+QITIEe9P6Oia9wwgxqFRoJb1wrNZ39Qt7Z6E9QF/aBnet+lGhbkO+Q6
gWSqnOHIJFgK0PI/4aumhgoYJyCwBBtcq0PvRkZOTaKYBFS3QgOHNTzKS+TtcUCy
XKcK/1+OLTEolTf8CV280SOiOV7a+MPM68jKYmOdyN4kcwcW7k8FqkCghzpZOXLY
3NQLHzEALBmJNQGRUL9Qah6LdYCO9A3urikjEQubVQ8yJb6Fx154u/kFGI7C8zkk
Y/QTTR94Jz1iqih0iU02qPjrrvBs7tJIOV19zRkVdQiZ9OGo1He6TEt8/3ZijQSb
fsw38rLncOgrxiuaFKLdMhzWmboH4khmaWHVQHgq6GFc90e6KQv8kGQO+9e/pynA
pAwnwHOGiGtHRkZmtvzA8UcVRSUeQahTUn5wEBjDKFivHYasJjdG3LSkllJqE6JU
GsMrzGnl4eqUTIk4d9bXZlQoZ4QCgAruhRb79QEiPbZq+MHCB/G5jJY60pT3ZsNS
Cfv4v0HK04tjiL44pD4iC6tukyS+2y+aScKk164Ic3bqYJ/vzFRhHFekmNT8fspc
U67zAcd4Wy/BY4m+KEYjJvtyRwc7lnB5fP1p9td3nj45JBkRFgvl2pyPM5lKU45z
QGjNRNkPeHtqek1VDanAC7k/w+o8blrGYH6vcRPVIjqUZr0iEtCYJ1zzVBwR0VCM
WPK0PVRC+FheGfW/vLRz/0LHGpkDNSRMFXXGiMDgP3rqt1+lq256HlksA56OkEAC
Fbl/sUeIk+Nk0JKaakrrp+WxMLaaQrIT28IqgcgsXJ0G4UflZX5YyPKWnmWrw73l
Ca+MsGOdQ781duu7PKzn5mraHY98Gt/UjbM63LF1bAMbCYKlobtzFk4R2HCF7S7D
y8BmhiDXoKIwTGHhupw0dtqGBj6OlNnN1cXsRW9kHZSogNkSzvBqmVSbQDjbtdoZ
DkjM8oQhecMXkikm2qSyneV3cujQAnZWyz6hlmLXIR0c0R8qeEwu+YiBI+H9Mai7
MGodd5lT+cs6pUnGnYCbVi5r/PT6pjpKEBJXsMbcd3hvpBg96FCbrWPgEmsIRqMU
20oBs53D94NA7HVlky2JDLxOzxfSRSK+KsxUhtrDVC0Mn5eN8NCAyUb3B0tgK3HC
rYWOIOquYtQGaUVHjeAPqEUdbmvt3DsuoRDajBvCiVN2pFmar9pHgAOAAPsmyynN
SzZzhwAfJ5QPnMriiXa48eEJ9xPPNavDg6og6g9D2ukk6dR7pYpT1suTCOlcw0ZN
wOBpGAm+jdYgGuiiZYs5v25XsU8I30y23oJ9DHWe+ew1FVNd3TYf+s2DSZfhG3J7
YrsjBS6GholPP4eIxMpKlZ6WOnbRBF4izkIxaXRWETmgCcO4ChMSntmDTi2F80OA
oOCyAwz8xXeMeqTPTSmPO3lTvujmQUem/mNHeMJ00amAhQR8GsEVvlzTUncH+7R0
ZpsuqdT9JqXJ7A8beeMUWp0xr8ROTuRaxlBt3UQjv1i6Pu7GmUowTewdagX30pKo
DLr5Xv9jL25jJjMRqrcpi+dBqTzKScC4pTfRum6JYXnRto3q1T8mVPR0CE39EfAN
zRke0rBrtQbqp9cVuouG6QZ0LlkEfBEOiZ3GghvVFrOuWcI7Hu6geVv9IvvjSqtW
8VgBg5B3GtPCttZQJJQKZ++oeVTVbmQpHthCokWgs/bw74+vEEx7gmxbpLLWdLy4
cFjs9lvC9Vchm7SvhByiYFXp6HM2RJlUm5WZuxaQgq0xR+p4W/46VaOkg5aTrRtU
q6/uZbD8pfhxF3uP4szXmiJB0faV3wDT39TzRepaDwOnyimvLA2N2yffuEDj6RCN
/5MeOs2mseBCGJCVsOhuX0uxCnYqRfbdlLSxWDT3QVyjcMlatphwLi7dugZ7g3im
eruVZJBCU5JLNlxZrzd0b7OqPCh/P7eCijkDl5Rpp2dvb58+Ykv384vbjJM88QBG
nM+Pfwf78oMb2gD47rW7TOMcrOuwcj393XuxAGKSGpTiPXY1/+7sIy+047QNoAM+
lpzm/sFAMhnADO0hHd4uIRkSQxPREbVqwiGtkCufESyZhsuihiW1/ChPhJucB67k
3cEIMw09AbaS76015HkejwvGAd9CFHc4aG3cFKGWJhFGwtdCm2A1VA6jbn7qxl5X
kzmbu1gkcDnCDG7xZ8NeRqDobhGBxQqMoHdVfTpIj678Jat2IAyTJ8Pm6NBoL++Z
wVqR/kJ+vG0m82nS6YHIHKNnGDYMucldodwvRyMNPTz+oh0U+F1+Rzr2/WGcTXJp
HiweEsADqZ2iaTpuMCJZJNHxnvEg16fX44Lwg8a7UR+Ul1Q3UeGT5sqKt75eTy2P
H05ousjCGxTYlp4RXad5S79Azryod/SYFlSP7rze+e+8ONjsV57+5L+am2duELt9
sAMd5CUXnQRnN555Rd4juul8BkqHU0SbpyGjei/psDE9dF9NXXHybeCKgiPjLIRf
XDTUeG0dFGO0VRtLBr2RbflbFx/ASALsqNmd/vvUuGLTs/VyXMle4hLTfBXwsbXw
VPlWyKe5NM5Wlm1QjklHmPd1x4dxLxlsBJb9aCFoshsDLHozzXofgSscwik6hS6j
No1Dc4flCQl7ZFI2JnZAG7qBHaKErIjBcCsVGBYErVjN7XxN3V+8V7t2RJc8Ic1F
kydcHqWeBDd0lPz+6u5mlMuax+0w1Ewyq3VF2W4LfA1MRke+NB9mNNInLiGmT0Bg
pLDy4R2aUAASADhJmNJzFloF4AMJ1BZSs+Cd/E8ujRdZxq504Gx7qzgKsDPmM88y
MM47BQTqBJALUztYHQ1fjGo4C+6pxSzL1h6tLNDCrMMPEZTRIOheX6nq6s3t+U3c
jkv3vPrX9Bq/MbBC2+ypzw==
`protect end_protected
