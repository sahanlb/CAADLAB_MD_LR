localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTZ_CHK = {
  {32'h43531850, 32'h00000000} /* (31, 31, 31) {real, imag} */,
  {32'h43e54e34, 32'h00000000} /* (31, 31, 30) {real, imag} */,
  {32'h43dc0070, 32'h00000000} /* (31, 31, 29) {real, imag} */,
  {32'h440ed220, 32'h00000000} /* (31, 31, 28) {real, imag} */,
  {32'h4467bbe2, 32'h00000000} /* (31, 31, 27) {real, imag} */,
  {32'h446e2458, 32'h00000000} /* (31, 31, 26) {real, imag} */,
  {32'h44af4751, 32'h00000000} /* (31, 31, 25) {real, imag} */,
  {32'h44a4de38, 32'h00000000} /* (31, 31, 24) {real, imag} */,
  {32'h448d5e25, 32'h00000000} /* (31, 31, 23) {real, imag} */,
  {32'h4475e80a, 32'h00000000} /* (31, 31, 22) {real, imag} */,
  {32'h447cc0e2, 32'h00000000} /* (31, 31, 21) {real, imag} */,
  {32'h4330bfe7, 32'h00000000} /* (31, 31, 20) {real, imag} */,
  {32'hc2a8d9bc, 32'h00000000} /* (31, 31, 19) {real, imag} */,
  {32'hc38eca5f, 32'h00000000} /* (31, 31, 18) {real, imag} */,
  {32'hc41e4b22, 32'h00000000} /* (31, 31, 17) {real, imag} */,
  {32'hc3f694de, 32'h00000000} /* (31, 31, 16) {real, imag} */,
  {32'hc48e751c, 32'h00000000} /* (31, 31, 15) {real, imag} */,
  {32'hc4e1a57b, 32'h00000000} /* (31, 31, 14) {real, imag} */,
  {32'hc49de363, 32'h00000000} /* (31, 31, 13) {real, imag} */,
  {32'hc48acb17, 32'h00000000} /* (31, 31, 12) {real, imag} */,
  {32'hc467b656, 32'h00000000} /* (31, 31, 11) {real, imag} */,
  {32'hc361a402, 32'h00000000} /* (31, 31, 10) {real, imag} */,
  {32'h43bc1cac, 32'h00000000} /* (31, 31, 9) {real, imag} */,
  {32'h4443c835, 32'h00000000} /* (31, 31, 8) {real, imag} */,
  {32'h43c2e2dc, 32'h00000000} /* (31, 31, 7) {real, imag} */,
  {32'h43715ac6, 32'h00000000} /* (31, 31, 6) {real, imag} */,
  {32'h44509c0c, 32'h00000000} /* (31, 31, 5) {real, imag} */,
  {32'h4424730e, 32'h00000000} /* (31, 31, 4) {real, imag} */,
  {32'h440aaaa4, 32'h00000000} /* (31, 31, 3) {real, imag} */,
  {32'h4463ea64, 32'h00000000} /* (31, 31, 2) {real, imag} */,
  {32'h43d30864, 32'h00000000} /* (31, 31, 1) {real, imag} */,
  {32'h43d95d14, 32'h00000000} /* (31, 31, 0) {real, imag} */,
  {32'h441ace83, 32'h00000000} /* (31, 30, 31) {real, imag} */,
  {32'h4397c48e, 32'h00000000} /* (31, 30, 30) {real, imag} */,
  {32'h4338ac80, 32'h00000000} /* (31, 30, 29) {real, imag} */,
  {32'h44407771, 32'h00000000} /* (31, 30, 28) {real, imag} */,
  {32'h44ac4b06, 32'h00000000} /* (31, 30, 27) {real, imag} */,
  {32'h44662c5a, 32'h00000000} /* (31, 30, 26) {real, imag} */,
  {32'h44e0493c, 32'h00000000} /* (31, 30, 25) {real, imag} */,
  {32'h44d5017e, 32'h00000000} /* (31, 30, 24) {real, imag} */,
  {32'h44c8c08c, 32'h00000000} /* (31, 30, 23) {real, imag} */,
  {32'h44992257, 32'h00000000} /* (31, 30, 22) {real, imag} */,
  {32'h44b8a944, 32'h00000000} /* (31, 30, 21) {real, imag} */,
  {32'h43d3ed18, 32'h00000000} /* (31, 30, 20) {real, imag} */,
  {32'hc46a696d, 32'h00000000} /* (31, 30, 19) {real, imag} */,
  {32'hc47f6075, 32'h00000000} /* (31, 30, 18) {real, imag} */,
  {32'hc4891bdc, 32'h00000000} /* (31, 30, 17) {real, imag} */,
  {32'hc49c574e, 32'h00000000} /* (31, 30, 16) {real, imag} */,
  {32'hc50f31d0, 32'h00000000} /* (31, 30, 15) {real, imag} */,
  {32'hc50fc44c, 32'h00000000} /* (31, 30, 14) {real, imag} */,
  {32'hc4ec87bc, 32'h00000000} /* (31, 30, 13) {real, imag} */,
  {32'hc4c39718, 32'h00000000} /* (31, 30, 12) {real, imag} */,
  {32'hc4853112, 32'h00000000} /* (31, 30, 11) {real, imag} */,
  {32'hc41d5e92, 32'h00000000} /* (31, 30, 10) {real, imag} */,
  {32'h438cf89e, 32'h00000000} /* (31, 30, 9) {real, imag} */,
  {32'h44431b1f, 32'h00000000} /* (31, 30, 8) {real, imag} */,
  {32'h448db6dc, 32'h00000000} /* (31, 30, 7) {real, imag} */,
  {32'h4407a960, 32'h00000000} /* (31, 30, 6) {real, imag} */,
  {32'h44957c40, 32'h00000000} /* (31, 30, 5) {real, imag} */,
  {32'h448c975b, 32'h00000000} /* (31, 30, 4) {real, imag} */,
  {32'h4457e963, 32'h00000000} /* (31, 30, 3) {real, imag} */,
  {32'h4455c573, 32'h00000000} /* (31, 30, 2) {real, imag} */,
  {32'h43b4e407, 32'h00000000} /* (31, 30, 1) {real, imag} */,
  {32'h43e8bfea, 32'h00000000} /* (31, 30, 0) {real, imag} */,
  {32'h4411eea9, 32'h00000000} /* (31, 29, 31) {real, imag} */,
  {32'h43ac6d80, 32'h00000000} /* (31, 29, 30) {real, imag} */,
  {32'h4464a116, 32'h00000000} /* (31, 29, 29) {real, imag} */,
  {32'h43afe79c, 32'h00000000} /* (31, 29, 28) {real, imag} */,
  {32'h440aef3c, 32'h00000000} /* (31, 29, 27) {real, imag} */,
  {32'h44a9d508, 32'h00000000} /* (31, 29, 26) {real, imag} */,
  {32'h44cbb520, 32'h00000000} /* (31, 29, 25) {real, imag} */,
  {32'h44b785fd, 32'h00000000} /* (31, 29, 24) {real, imag} */,
  {32'h448cc111, 32'h00000000} /* (31, 29, 23) {real, imag} */,
  {32'h44e5041e, 32'h00000000} /* (31, 29, 22) {real, imag} */,
  {32'hc319da74, 32'h00000000} /* (31, 29, 21) {real, imag} */,
  {32'hc42bebc7, 32'h00000000} /* (31, 29, 20) {real, imag} */,
  {32'hc3896937, 32'h00000000} /* (31, 29, 19) {real, imag} */,
  {32'hc4a2a60b, 32'h00000000} /* (31, 29, 18) {real, imag} */,
  {32'hc4c45d18, 32'h00000000} /* (31, 29, 17) {real, imag} */,
  {32'hc4b18170, 32'h00000000} /* (31, 29, 16) {real, imag} */,
  {32'hc4f00d16, 32'h00000000} /* (31, 29, 15) {real, imag} */,
  {32'hc4c3bd14, 32'h00000000} /* (31, 29, 14) {real, imag} */,
  {32'hc500f930, 32'h00000000} /* (31, 29, 13) {real, imag} */,
  {32'hc4a3f4c2, 32'h00000000} /* (31, 29, 12) {real, imag} */,
  {32'hc4b35c74, 32'h00000000} /* (31, 29, 11) {real, imag} */,
  {32'hc40f2a9b, 32'h00000000} /* (31, 29, 10) {real, imag} */,
  {32'h44165881, 32'h00000000} /* (31, 29, 9) {real, imag} */,
  {32'h44607246, 32'h00000000} /* (31, 29, 8) {real, imag} */,
  {32'h4453927b, 32'h00000000} /* (31, 29, 7) {real, imag} */,
  {32'h4471c0e1, 32'h00000000} /* (31, 29, 6) {real, imag} */,
  {32'h447b4fc3, 32'h00000000} /* (31, 29, 5) {real, imag} */,
  {32'h44e34ea2, 32'h00000000} /* (31, 29, 4) {real, imag} */,
  {32'h447f2f4c, 32'h00000000} /* (31, 29, 3) {real, imag} */,
  {32'h44ba44bf, 32'h00000000} /* (31, 29, 2) {real, imag} */,
  {32'h446257fb, 32'h00000000} /* (31, 29, 1) {real, imag} */,
  {32'h43e98f9c, 32'h00000000} /* (31, 29, 0) {real, imag} */,
  {32'h4417cf9c, 32'h00000000} /* (31, 28, 31) {real, imag} */,
  {32'h446dec18, 32'h00000000} /* (31, 28, 30) {real, imag} */,
  {32'h4457bfa3, 32'h00000000} /* (31, 28, 29) {real, imag} */,
  {32'h44863dea, 32'h00000000} /* (31, 28, 28) {real, imag} */,
  {32'h4416d5e9, 32'h00000000} /* (31, 28, 27) {real, imag} */,
  {32'h44c3f028, 32'h00000000} /* (31, 28, 26) {real, imag} */,
  {32'h44bff62e, 32'h00000000} /* (31, 28, 25) {real, imag} */,
  {32'h449086f3, 32'h00000000} /* (31, 28, 24) {real, imag} */,
  {32'h44873538, 32'h00000000} /* (31, 28, 23) {real, imag} */,
  {32'h445820ba, 32'h00000000} /* (31, 28, 22) {real, imag} */,
  {32'h436fa9f8, 32'h00000000} /* (31, 28, 21) {real, imag} */,
  {32'hc4ac77c4, 32'h00000000} /* (31, 28, 20) {real, imag} */,
  {32'hc480547e, 32'h00000000} /* (31, 28, 19) {real, imag} */,
  {32'hc3e7d5c7, 32'h00000000} /* (31, 28, 18) {real, imag} */,
  {32'hc33920ec, 32'h00000000} /* (31, 28, 17) {real, imag} */,
  {32'hc4a3e1bb, 32'h00000000} /* (31, 28, 16) {real, imag} */,
  {32'hc4bec850, 32'h00000000} /* (31, 28, 15) {real, imag} */,
  {32'hc4cec7f0, 32'h00000000} /* (31, 28, 14) {real, imag} */,
  {32'hc49a0df2, 32'h00000000} /* (31, 28, 13) {real, imag} */,
  {32'hc4a38200, 32'h00000000} /* (31, 28, 12) {real, imag} */,
  {32'hc445af93, 32'h00000000} /* (31, 28, 11) {real, imag} */,
  {32'h434a88dc, 32'h00000000} /* (31, 28, 10) {real, imag} */,
  {32'h43f548b8, 32'h00000000} /* (31, 28, 9) {real, imag} */,
  {32'h4496e15f, 32'h00000000} /* (31, 28, 8) {real, imag} */,
  {32'h444e842d, 32'h00000000} /* (31, 28, 7) {real, imag} */,
  {32'h4466060a, 32'h00000000} /* (31, 28, 6) {real, imag} */,
  {32'h4480d8e4, 32'h00000000} /* (31, 28, 5) {real, imag} */,
  {32'h44363d8c, 32'h00000000} /* (31, 28, 4) {real, imag} */,
  {32'h446eee45, 32'h00000000} /* (31, 28, 3) {real, imag} */,
  {32'h448ec922, 32'h00000000} /* (31, 28, 2) {real, imag} */,
  {32'h449658b8, 32'h00000000} /* (31, 28, 1) {real, imag} */,
  {32'h4430a3ee, 32'h00000000} /* (31, 28, 0) {real, imag} */,
  {32'h43ee7a84, 32'h00000000} /* (31, 27, 31) {real, imag} */,
  {32'h4471ee86, 32'h00000000} /* (31, 27, 30) {real, imag} */,
  {32'h432e006e, 32'h00000000} /* (31, 27, 29) {real, imag} */,
  {32'h447e8d4b, 32'h00000000} /* (31, 27, 28) {real, imag} */,
  {32'h44a0174d, 32'h00000000} /* (31, 27, 27) {real, imag} */,
  {32'h44fddcf8, 32'h00000000} /* (31, 27, 26) {real, imag} */,
  {32'h44ed3fe2, 32'h00000000} /* (31, 27, 25) {real, imag} */,
  {32'h4434631a, 32'h00000000} /* (31, 27, 24) {real, imag} */,
  {32'h44744356, 32'h00000000} /* (31, 27, 23) {real, imag} */,
  {32'h448bc4fb, 32'h00000000} /* (31, 27, 22) {real, imag} */,
  {32'h4466f8b0, 32'h00000000} /* (31, 27, 21) {real, imag} */,
  {32'hc39666fe, 32'h00000000} /* (31, 27, 20) {real, imag} */,
  {32'h4387d69e, 32'h00000000} /* (31, 27, 19) {real, imag} */,
  {32'hc40114aa, 32'h00000000} /* (31, 27, 18) {real, imag} */,
  {32'hc488c635, 32'h00000000} /* (31, 27, 17) {real, imag} */,
  {32'hc48d0d10, 32'h00000000} /* (31, 27, 16) {real, imag} */,
  {32'hc4ccc8f7, 32'h00000000} /* (31, 27, 15) {real, imag} */,
  {32'hc4c485c3, 32'h00000000} /* (31, 27, 14) {real, imag} */,
  {32'hc493feb1, 32'h00000000} /* (31, 27, 13) {real, imag} */,
  {32'hc4026d6d, 32'h00000000} /* (31, 27, 12) {real, imag} */,
  {32'hc3d083b4, 32'h00000000} /* (31, 27, 11) {real, imag} */,
  {32'h4425b1a8, 32'h00000000} /* (31, 27, 10) {real, imag} */,
  {32'h43888fb8, 32'h00000000} /* (31, 27, 9) {real, imag} */,
  {32'h44a72273, 32'h00000000} /* (31, 27, 8) {real, imag} */,
  {32'h44841e87, 32'h00000000} /* (31, 27, 7) {real, imag} */,
  {32'h44a5e1e7, 32'h00000000} /* (31, 27, 6) {real, imag} */,
  {32'h448d136c, 32'h00000000} /* (31, 27, 5) {real, imag} */,
  {32'h445f257b, 32'h00000000} /* (31, 27, 4) {real, imag} */,
  {32'h44977ff2, 32'h00000000} /* (31, 27, 3) {real, imag} */,
  {32'h443b7244, 32'h00000000} /* (31, 27, 2) {real, imag} */,
  {32'h44061662, 32'h00000000} /* (31, 27, 1) {real, imag} */,
  {32'h43c7f649, 32'h00000000} /* (31, 27, 0) {real, imag} */,
  {32'h43e93a74, 32'h00000000} /* (31, 26, 31) {real, imag} */,
  {32'h43f04aa6, 32'h00000000} /* (31, 26, 30) {real, imag} */,
  {32'h440248ac, 32'h00000000} /* (31, 26, 29) {real, imag} */,
  {32'h43b714c5, 32'h00000000} /* (31, 26, 28) {real, imag} */,
  {32'h44b7508d, 32'h00000000} /* (31, 26, 27) {real, imag} */,
  {32'h44e75480, 32'h00000000} /* (31, 26, 26) {real, imag} */,
  {32'h44a854f7, 32'h00000000} /* (31, 26, 25) {real, imag} */,
  {32'h44f5cd3b, 32'h00000000} /* (31, 26, 24) {real, imag} */,
  {32'h44b998bb, 32'h00000000} /* (31, 26, 23) {real, imag} */,
  {32'h448f4310, 32'h00000000} /* (31, 26, 22) {real, imag} */,
  {32'h449e5d24, 32'h00000000} /* (31, 26, 21) {real, imag} */,
  {32'h437fe23e, 32'h00000000} /* (31, 26, 20) {real, imag} */,
  {32'hc3487a2e, 32'h00000000} /* (31, 26, 19) {real, imag} */,
  {32'hc4a938ba, 32'h00000000} /* (31, 26, 18) {real, imag} */,
  {32'hc4196623, 32'h00000000} /* (31, 26, 17) {real, imag} */,
  {32'hc4c41785, 32'h00000000} /* (31, 26, 16) {real, imag} */,
  {32'hc51e31b0, 32'h00000000} /* (31, 26, 15) {real, imag} */,
  {32'hc4d1a1b0, 32'h00000000} /* (31, 26, 14) {real, imag} */,
  {32'hc4a5dc82, 32'h00000000} /* (31, 26, 13) {real, imag} */,
  {32'hc42646f4, 32'h00000000} /* (31, 26, 12) {real, imag} */,
  {32'hc4328d66, 32'h00000000} /* (31, 26, 11) {real, imag} */,
  {32'hc33cf100, 32'h00000000} /* (31, 26, 10) {real, imag} */,
  {32'h44853d43, 32'h00000000} /* (31, 26, 9) {real, imag} */,
  {32'h44a9afd5, 32'h00000000} /* (31, 26, 8) {real, imag} */,
  {32'h44b9c2db, 32'h00000000} /* (31, 26, 7) {real, imag} */,
  {32'h44d95db8, 32'h00000000} /* (31, 26, 6) {real, imag} */,
  {32'h449ae4e4, 32'h00000000} /* (31, 26, 5) {real, imag} */,
  {32'h44805e3c, 32'h00000000} /* (31, 26, 4) {real, imag} */,
  {32'h448107fa, 32'h00000000} /* (31, 26, 3) {real, imag} */,
  {32'h4492c326, 32'h00000000} /* (31, 26, 2) {real, imag} */,
  {32'h442b4287, 32'h00000000} /* (31, 26, 1) {real, imag} */,
  {32'h43862c44, 32'h00000000} /* (31, 26, 0) {real, imag} */,
  {32'h438897b0, 32'h00000000} /* (31, 25, 31) {real, imag} */,
  {32'h4403d7be, 32'h00000000} /* (31, 25, 30) {real, imag} */,
  {32'h43ca7b20, 32'h00000000} /* (31, 25, 29) {real, imag} */,
  {32'h43b4df78, 32'h00000000} /* (31, 25, 28) {real, imag} */,
  {32'h44891a88, 32'h00000000} /* (31, 25, 27) {real, imag} */,
  {32'h44b45b52, 32'h00000000} /* (31, 25, 26) {real, imag} */,
  {32'h44b51662, 32'h00000000} /* (31, 25, 25) {real, imag} */,
  {32'h44c2df04, 32'h00000000} /* (31, 25, 24) {real, imag} */,
  {32'h4479825d, 32'h00000000} /* (31, 25, 23) {real, imag} */,
  {32'h44e54d35, 32'h00000000} /* (31, 25, 22) {real, imag} */,
  {32'h43fc8608, 32'h00000000} /* (31, 25, 21) {real, imag} */,
  {32'hc3d4027e, 32'h00000000} /* (31, 25, 20) {real, imag} */,
  {32'hc3d55b65, 32'h00000000} /* (31, 25, 19) {real, imag} */,
  {32'hc46ca186, 32'h00000000} /* (31, 25, 18) {real, imag} */,
  {32'hc4e73b46, 32'h00000000} /* (31, 25, 17) {real, imag} */,
  {32'hc4c31918, 32'h00000000} /* (31, 25, 16) {real, imag} */,
  {32'hc4ebd3ec, 32'h00000000} /* (31, 25, 15) {real, imag} */,
  {32'hc4bef11d, 32'h00000000} /* (31, 25, 14) {real, imag} */,
  {32'hc49b498e, 32'h00000000} /* (31, 25, 13) {real, imag} */,
  {32'hc4d342f6, 32'h00000000} /* (31, 25, 12) {real, imag} */,
  {32'hc446663a, 32'h00000000} /* (31, 25, 11) {real, imag} */,
  {32'h43c032a0, 32'h00000000} /* (31, 25, 10) {real, imag} */,
  {32'h446efab0, 32'h00000000} /* (31, 25, 9) {real, imag} */,
  {32'h44ca87e8, 32'h00000000} /* (31, 25, 8) {real, imag} */,
  {32'h4503c8bf, 32'h00000000} /* (31, 25, 7) {real, imag} */,
  {32'h44bc5d39, 32'h00000000} /* (31, 25, 6) {real, imag} */,
  {32'h452c7604, 32'h00000000} /* (31, 25, 5) {real, imag} */,
  {32'h44ab0f70, 32'h00000000} /* (31, 25, 4) {real, imag} */,
  {32'h44af4c2e, 32'h00000000} /* (31, 25, 3) {real, imag} */,
  {32'h44837ce4, 32'h00000000} /* (31, 25, 2) {real, imag} */,
  {32'h4400741c, 32'h00000000} /* (31, 25, 1) {real, imag} */,
  {32'h440d8773, 32'h00000000} /* (31, 25, 0) {real, imag} */,
  {32'h43ddd5e2, 32'h00000000} /* (31, 24, 31) {real, imag} */,
  {32'h44c3af72, 32'h00000000} /* (31, 24, 30) {real, imag} */,
  {32'h44aa7376, 32'h00000000} /* (31, 24, 29) {real, imag} */,
  {32'h4434d96c, 32'h00000000} /* (31, 24, 28) {real, imag} */,
  {32'h44527e11, 32'h00000000} /* (31, 24, 27) {real, imag} */,
  {32'h44a873d8, 32'h00000000} /* (31, 24, 26) {real, imag} */,
  {32'h44993ff1, 32'h00000000} /* (31, 24, 25) {real, imag} */,
  {32'h44c65789, 32'h00000000} /* (31, 24, 24) {real, imag} */,
  {32'h44af1895, 32'h00000000} /* (31, 24, 23) {real, imag} */,
  {32'h44f29480, 32'h00000000} /* (31, 24, 22) {real, imag} */,
  {32'h44186775, 32'h00000000} /* (31, 24, 21) {real, imag} */,
  {32'h43a60a34, 32'h00000000} /* (31, 24, 20) {real, imag} */,
  {32'h433f7244, 32'h00000000} /* (31, 24, 19) {real, imag} */,
  {32'hc3c25643, 32'h00000000} /* (31, 24, 18) {real, imag} */,
  {32'hc4e245b2, 32'h00000000} /* (31, 24, 17) {real, imag} */,
  {32'hc4e0105e, 32'h00000000} /* (31, 24, 16) {real, imag} */,
  {32'hc4683187, 32'h00000000} /* (31, 24, 15) {real, imag} */,
  {32'hc4baf8b6, 32'h00000000} /* (31, 24, 14) {real, imag} */,
  {32'hc495040c, 32'h00000000} /* (31, 24, 13) {real, imag} */,
  {32'hc4a89180, 32'h00000000} /* (31, 24, 12) {real, imag} */,
  {32'hc389fbde, 32'h00000000} /* (31, 24, 11) {real, imag} */,
  {32'h443d3a70, 32'h00000000} /* (31, 24, 10) {real, imag} */,
  {32'h4496cb63, 32'h00000000} /* (31, 24, 9) {real, imag} */,
  {32'h44bfe3c9, 32'h00000000} /* (31, 24, 8) {real, imag} */,
  {32'h44b870d3, 32'h00000000} /* (31, 24, 7) {real, imag} */,
  {32'h4500ce4e, 32'h00000000} /* (31, 24, 6) {real, imag} */,
  {32'h45238785, 32'h00000000} /* (31, 24, 5) {real, imag} */,
  {32'h44ae6af1, 32'h00000000} /* (31, 24, 4) {real, imag} */,
  {32'h44883762, 32'h00000000} /* (31, 24, 3) {real, imag} */,
  {32'h44908364, 32'h00000000} /* (31, 24, 2) {real, imag} */,
  {32'h440c5953, 32'h00000000} /* (31, 24, 1) {real, imag} */,
  {32'h43aeadf0, 32'h00000000} /* (31, 24, 0) {real, imag} */,
  {32'h437afce4, 32'h00000000} /* (31, 23, 31) {real, imag} */,
  {32'h44c1254c, 32'h00000000} /* (31, 23, 30) {real, imag} */,
  {32'h449ad582, 32'h00000000} /* (31, 23, 29) {real, imag} */,
  {32'h4448a4ba, 32'h00000000} /* (31, 23, 28) {real, imag} */,
  {32'h441372d8, 32'h00000000} /* (31, 23, 27) {real, imag} */,
  {32'h44984de6, 32'h00000000} /* (31, 23, 26) {real, imag} */,
  {32'h446e6447, 32'h00000000} /* (31, 23, 25) {real, imag} */,
  {32'h44508303, 32'h00000000} /* (31, 23, 24) {real, imag} */,
  {32'h44fb79d6, 32'h00000000} /* (31, 23, 23) {real, imag} */,
  {32'h44d003cb, 32'h00000000} /* (31, 23, 22) {real, imag} */,
  {32'h448411ec, 32'h00000000} /* (31, 23, 21) {real, imag} */,
  {32'h43baefbb, 32'h00000000} /* (31, 23, 20) {real, imag} */,
  {32'hc3cb2e22, 32'h00000000} /* (31, 23, 19) {real, imag} */,
  {32'hc43c6096, 32'h00000000} /* (31, 23, 18) {real, imag} */,
  {32'hc4360b66, 32'h00000000} /* (31, 23, 17) {real, imag} */,
  {32'hc49f0461, 32'h00000000} /* (31, 23, 16) {real, imag} */,
  {32'hc4ae102e, 32'h00000000} /* (31, 23, 15) {real, imag} */,
  {32'hc4b4f638, 32'h00000000} /* (31, 23, 14) {real, imag} */,
  {32'hc3d8e6da, 32'h00000000} /* (31, 23, 13) {real, imag} */,
  {32'hc32b9148, 32'h00000000} /* (31, 23, 12) {real, imag} */,
  {32'h424d2718, 32'h00000000} /* (31, 23, 11) {real, imag} */,
  {32'h440fe46c, 32'h00000000} /* (31, 23, 10) {real, imag} */,
  {32'h44bf1e1e, 32'h00000000} /* (31, 23, 9) {real, imag} */,
  {32'h4484def3, 32'h00000000} /* (31, 23, 8) {real, imag} */,
  {32'h44c5bd08, 32'h00000000} /* (31, 23, 7) {real, imag} */,
  {32'h44d51329, 32'h00000000} /* (31, 23, 6) {real, imag} */,
  {32'h448b26d4, 32'h00000000} /* (31, 23, 5) {real, imag} */,
  {32'h44aa4431, 32'h00000000} /* (31, 23, 4) {real, imag} */,
  {32'h44fcfeb4, 32'h00000000} /* (31, 23, 3) {real, imag} */,
  {32'h44c61c77, 32'h00000000} /* (31, 23, 2) {real, imag} */,
  {32'h449458db, 32'h00000000} /* (31, 23, 1) {real, imag} */,
  {32'h445bd276, 32'h00000000} /* (31, 23, 0) {real, imag} */,
  {32'hc1bcca90, 32'h00000000} /* (31, 22, 31) {real, imag} */,
  {32'h43b6a1da, 32'h00000000} /* (31, 22, 30) {real, imag} */,
  {32'h421a1748, 32'h00000000} /* (31, 22, 29) {real, imag} */,
  {32'hc33d1d50, 32'h00000000} /* (31, 22, 28) {real, imag} */,
  {32'hc0c931c0, 32'h00000000} /* (31, 22, 27) {real, imag} */,
  {32'hc229e510, 32'h00000000} /* (31, 22, 26) {real, imag} */,
  {32'h4411ada1, 32'h00000000} /* (31, 22, 25) {real, imag} */,
  {32'h445caab8, 32'h00000000} /* (31, 22, 24) {real, imag} */,
  {32'h44ff26cc, 32'h00000000} /* (31, 22, 23) {real, imag} */,
  {32'h45017a16, 32'h00000000} /* (31, 22, 22) {real, imag} */,
  {32'h446f0523, 32'h00000000} /* (31, 22, 21) {real, imag} */,
  {32'h4316d378, 32'h00000000} /* (31, 22, 20) {real, imag} */,
  {32'hc4801439, 32'h00000000} /* (31, 22, 19) {real, imag} */,
  {32'hc3dcae44, 32'h00000000} /* (31, 22, 18) {real, imag} */,
  {32'hc455c97a, 32'h00000000} /* (31, 22, 17) {real, imag} */,
  {32'hc4ddab13, 32'h00000000} /* (31, 22, 16) {real, imag} */,
  {32'hc4538b58, 32'h00000000} /* (31, 22, 15) {real, imag} */,
  {32'hc426d3bf, 32'h00000000} /* (31, 22, 14) {real, imag} */,
  {32'hc3581752, 32'h00000000} /* (31, 22, 13) {real, imag} */,
  {32'hc2acd878, 32'h00000000} /* (31, 22, 12) {real, imag} */,
  {32'h42765248, 32'h00000000} /* (31, 22, 11) {real, imag} */,
  {32'h444fe25d, 32'h00000000} /* (31, 22, 10) {real, imag} */,
  {32'h44e3c512, 32'h00000000} /* (31, 22, 9) {real, imag} */,
  {32'h44afb7b4, 32'h00000000} /* (31, 22, 8) {real, imag} */,
  {32'h4472be3b, 32'h00000000} /* (31, 22, 7) {real, imag} */,
  {32'h446b4d82, 32'h00000000} /* (31, 22, 6) {real, imag} */,
  {32'h447d4cd5, 32'h00000000} /* (31, 22, 5) {real, imag} */,
  {32'h44ff19cb, 32'h00000000} /* (31, 22, 4) {real, imag} */,
  {32'h44ac303f, 32'h00000000} /* (31, 22, 3) {real, imag} */,
  {32'h4500ab24, 32'h00000000} /* (31, 22, 2) {real, imag} */,
  {32'h446879ae, 32'h00000000} /* (31, 22, 1) {real, imag} */,
  {32'h44476f32, 32'h00000000} /* (31, 22, 0) {real, imag} */,
  {32'hc38def3c, 32'h00000000} /* (31, 21, 31) {real, imag} */,
  {32'h438ca115, 32'h00000000} /* (31, 21, 30) {real, imag} */,
  {32'hc2b46ecc, 32'h00000000} /* (31, 21, 29) {real, imag} */,
  {32'h434134fe, 32'h00000000} /* (31, 21, 28) {real, imag} */,
  {32'hc406dd64, 32'h00000000} /* (31, 21, 27) {real, imag} */,
  {32'hc336da4e, 32'h00000000} /* (31, 21, 26) {real, imag} */,
  {32'hc2323d38, 32'h00000000} /* (31, 21, 25) {real, imag} */,
  {32'h438c9988, 32'h00000000} /* (31, 21, 24) {real, imag} */,
  {32'h4474f039, 32'h00000000} /* (31, 21, 23) {real, imag} */,
  {32'h43ad8e33, 32'h00000000} /* (31, 21, 22) {real, imag} */,
  {32'h43f950bc, 32'h00000000} /* (31, 21, 21) {real, imag} */,
  {32'h43bcd491, 32'h00000000} /* (31, 21, 20) {real, imag} */,
  {32'h42638220, 32'h00000000} /* (31, 21, 19) {real, imag} */,
  {32'hc3f2bc64, 32'h00000000} /* (31, 21, 18) {real, imag} */,
  {32'hc47f0dc2, 32'h00000000} /* (31, 21, 17) {real, imag} */,
  {32'hc32e388c, 32'h00000000} /* (31, 21, 16) {real, imag} */,
  {32'h4258f004, 32'h00000000} /* (31, 21, 15) {real, imag} */,
  {32'hc3856a7f, 32'h00000000} /* (31, 21, 14) {real, imag} */,
  {32'h43ade8ad, 32'h00000000} /* (31, 21, 13) {real, imag} */,
  {32'h4465ddc4, 32'h00000000} /* (31, 21, 12) {real, imag} */,
  {32'h44002f24, 32'h00000000} /* (31, 21, 11) {real, imag} */,
  {32'h43d49f8d, 32'h00000000} /* (31, 21, 10) {real, imag} */,
  {32'h444f2b66, 32'h00000000} /* (31, 21, 9) {real, imag} */,
  {32'h44025091, 32'h00000000} /* (31, 21, 8) {real, imag} */,
  {32'h42656bb0, 32'h00000000} /* (31, 21, 7) {real, imag} */,
  {32'h440aa9a6, 32'h00000000} /* (31, 21, 6) {real, imag} */,
  {32'h438e6942, 32'h00000000} /* (31, 21, 5) {real, imag} */,
  {32'h44397e20, 32'h00000000} /* (31, 21, 4) {real, imag} */,
  {32'h43fd4fac, 32'h00000000} /* (31, 21, 3) {real, imag} */,
  {32'h439ae1ce, 32'h00000000} /* (31, 21, 2) {real, imag} */,
  {32'h429e1064, 32'h00000000} /* (31, 21, 1) {real, imag} */,
  {32'hc4206176, 32'h00000000} /* (31, 21, 0) {real, imag} */,
  {32'hc4310f4a, 32'h00000000} /* (31, 20, 31) {real, imag} */,
  {32'hc45a3acf, 32'h00000000} /* (31, 20, 30) {real, imag} */,
  {32'hc4a78a42, 32'h00000000} /* (31, 20, 29) {real, imag} */,
  {32'hc3d5f5e1, 32'h00000000} /* (31, 20, 28) {real, imag} */,
  {32'hc46ffd8c, 32'h00000000} /* (31, 20, 27) {real, imag} */,
  {32'hc40ca3da, 32'h00000000} /* (31, 20, 26) {real, imag} */,
  {32'hc396a256, 32'h00000000} /* (31, 20, 25) {real, imag} */,
  {32'hc4c2622e, 32'h00000000} /* (31, 20, 24) {real, imag} */,
  {32'hc48575e6, 32'h00000000} /* (31, 20, 23) {real, imag} */,
  {32'hc3466628, 32'h00000000} /* (31, 20, 22) {real, imag} */,
  {32'hc3f11c48, 32'h00000000} /* (31, 20, 21) {real, imag} */,
  {32'h440e0d7e, 32'h00000000} /* (31, 20, 20) {real, imag} */,
  {32'h43d46cf8, 32'h00000000} /* (31, 20, 19) {real, imag} */,
  {32'h43b8ebd6, 32'h00000000} /* (31, 20, 18) {real, imag} */,
  {32'h42948acc, 32'h00000000} /* (31, 20, 17) {real, imag} */,
  {32'h43938b25, 32'h00000000} /* (31, 20, 16) {real, imag} */,
  {32'h447ec370, 32'h00000000} /* (31, 20, 15) {real, imag} */,
  {32'h4468b3bd, 32'h00000000} /* (31, 20, 14) {real, imag} */,
  {32'h44f5e13a, 32'h00000000} /* (31, 20, 13) {real, imag} */,
  {32'h44b131ee, 32'h00000000} /* (31, 20, 12) {real, imag} */,
  {32'h4431417c, 32'h00000000} /* (31, 20, 11) {real, imag} */,
  {32'h4382d1fc, 32'h00000000} /* (31, 20, 10) {real, imag} */,
  {32'hc33f7d00, 32'h00000000} /* (31, 20, 9) {real, imag} */,
  {32'hc46f6f3c, 32'h00000000} /* (31, 20, 8) {real, imag} */,
  {32'hc4c7b7d2, 32'h00000000} /* (31, 20, 7) {real, imag} */,
  {32'hc4e1b2e4, 32'h00000000} /* (31, 20, 6) {real, imag} */,
  {32'hc43efa5c, 32'h00000000} /* (31, 20, 5) {real, imag} */,
  {32'hc47239a4, 32'h00000000} /* (31, 20, 4) {real, imag} */,
  {32'hc48776b6, 32'h00000000} /* (31, 20, 3) {real, imag} */,
  {32'hc489623a, 32'h00000000} /* (31, 20, 2) {real, imag} */,
  {32'hc46f51c4, 32'h00000000} /* (31, 20, 1) {real, imag} */,
  {32'hc4a194a3, 32'h00000000} /* (31, 20, 0) {real, imag} */,
  {32'hc47e4c93, 32'h00000000} /* (31, 19, 31) {real, imag} */,
  {32'hc4c1a437, 32'h00000000} /* (31, 19, 30) {real, imag} */,
  {32'hc450ba73, 32'h00000000} /* (31, 19, 29) {real, imag} */,
  {32'hc4ab7e54, 32'h00000000} /* (31, 19, 28) {real, imag} */,
  {32'hc49f1580, 32'h00000000} /* (31, 19, 27) {real, imag} */,
  {32'hc4b77922, 32'h00000000} /* (31, 19, 26) {real, imag} */,
  {32'hc4c9b1d3, 32'h00000000} /* (31, 19, 25) {real, imag} */,
  {32'hc4551b81, 32'h00000000} /* (31, 19, 24) {real, imag} */,
  {32'hc4c2f41e, 32'h00000000} /* (31, 19, 23) {real, imag} */,
  {32'hc3ea76c5, 32'h00000000} /* (31, 19, 22) {real, imag} */,
  {32'hc319a044, 32'h00000000} /* (31, 19, 21) {real, imag} */,
  {32'h431bc4f0, 32'h00000000} /* (31, 19, 20) {real, imag} */,
  {32'h447eacf8, 32'h00000000} /* (31, 19, 19) {real, imag} */,
  {32'h44e2b92a, 32'h00000000} /* (31, 19, 18) {real, imag} */,
  {32'h44355ceb, 32'h00000000} /* (31, 19, 17) {real, imag} */,
  {32'h44adeb7a, 32'h00000000} /* (31, 19, 16) {real, imag} */,
  {32'h44ed7784, 32'h00000000} /* (31, 19, 15) {real, imag} */,
  {32'h44ce233d, 32'h00000000} /* (31, 19, 14) {real, imag} */,
  {32'h4508d34d, 32'h00000000} /* (31, 19, 13) {real, imag} */,
  {32'h44d85d62, 32'h00000000} /* (31, 19, 12) {real, imag} */,
  {32'h44a44148, 32'h00000000} /* (31, 19, 11) {real, imag} */,
  {32'hc3cf08de, 32'h00000000} /* (31, 19, 10) {real, imag} */,
  {32'hc4c19541, 32'h00000000} /* (31, 19, 9) {real, imag} */,
  {32'hc5009f2a, 32'h00000000} /* (31, 19, 8) {real, imag} */,
  {32'hc4c3ca66, 32'h00000000} /* (31, 19, 7) {real, imag} */,
  {32'hc49bf367, 32'h00000000} /* (31, 19, 6) {real, imag} */,
  {32'hc498ad72, 32'h00000000} /* (31, 19, 5) {real, imag} */,
  {32'hc4b7e58e, 32'h00000000} /* (31, 19, 4) {real, imag} */,
  {32'hc51a6c4d, 32'h00000000} /* (31, 19, 3) {real, imag} */,
  {32'hc4981692, 32'h00000000} /* (31, 19, 2) {real, imag} */,
  {32'hc4ef48f2, 32'h00000000} /* (31, 19, 1) {real, imag} */,
  {32'hc4eb3312, 32'h00000000} /* (31, 19, 0) {real, imag} */,
  {32'hc5013eb0, 32'h00000000} /* (31, 18, 31) {real, imag} */,
  {32'hc4bd8201, 32'h00000000} /* (31, 18, 30) {real, imag} */,
  {32'hc48dd913, 32'h00000000} /* (31, 18, 29) {real, imag} */,
  {32'hc4936196, 32'h00000000} /* (31, 18, 28) {real, imag} */,
  {32'hc4224777, 32'h00000000} /* (31, 18, 27) {real, imag} */,
  {32'hc466b6c8, 32'h00000000} /* (31, 18, 26) {real, imag} */,
  {32'hc4631ba0, 32'h00000000} /* (31, 18, 25) {real, imag} */,
  {32'hc4833725, 32'h00000000} /* (31, 18, 24) {real, imag} */,
  {32'hc4adc5b7, 32'h00000000} /* (31, 18, 23) {real, imag} */,
  {32'hc38c50ea, 32'h00000000} /* (31, 18, 22) {real, imag} */,
  {32'hc1b43c10, 32'h00000000} /* (31, 18, 21) {real, imag} */,
  {32'h4489d3db, 32'h00000000} /* (31, 18, 20) {real, imag} */,
  {32'h44d66dba, 32'h00000000} /* (31, 18, 19) {real, imag} */,
  {32'h44c15ece, 32'h00000000} /* (31, 18, 18) {real, imag} */,
  {32'h44a2e9f4, 32'h00000000} /* (31, 18, 17) {real, imag} */,
  {32'h44a15042, 32'h00000000} /* (31, 18, 16) {real, imag} */,
  {32'h44d5b202, 32'h00000000} /* (31, 18, 15) {real, imag} */,
  {32'h44c9a52f, 32'h00000000} /* (31, 18, 14) {real, imag} */,
  {32'h451219a6, 32'h00000000} /* (31, 18, 13) {real, imag} */,
  {32'h45042542, 32'h00000000} /* (31, 18, 12) {real, imag} */,
  {32'h444cf025, 32'h00000000} /* (31, 18, 11) {real, imag} */,
  {32'hc3d3b3d4, 32'h00000000} /* (31, 18, 10) {real, imag} */,
  {32'hc4b4e174, 32'h00000000} /* (31, 18, 9) {real, imag} */,
  {32'hc4d6ea6b, 32'h00000000} /* (31, 18, 8) {real, imag} */,
  {32'hc4f05b3d, 32'h00000000} /* (31, 18, 7) {real, imag} */,
  {32'hc4dad598, 32'h00000000} /* (31, 18, 6) {real, imag} */,
  {32'hc478e39a, 32'h00000000} /* (31, 18, 5) {real, imag} */,
  {32'hc4a508e9, 32'h00000000} /* (31, 18, 4) {real, imag} */,
  {32'hc4a801f6, 32'h00000000} /* (31, 18, 3) {real, imag} */,
  {32'hc4ecee76, 32'h00000000} /* (31, 18, 2) {real, imag} */,
  {32'hc4f92b5c, 32'h00000000} /* (31, 18, 1) {real, imag} */,
  {32'hc4974458, 32'h00000000} /* (31, 18, 0) {real, imag} */,
  {32'hc4b99560, 32'h00000000} /* (31, 17, 31) {real, imag} */,
  {32'hc4b16cb0, 32'h00000000} /* (31, 17, 30) {real, imag} */,
  {32'hc49fb55e, 32'h00000000} /* (31, 17, 29) {real, imag} */,
  {32'hc4809dfa, 32'h00000000} /* (31, 17, 28) {real, imag} */,
  {32'hc46a8576, 32'h00000000} /* (31, 17, 27) {real, imag} */,
  {32'hc45b4322, 32'h00000000} /* (31, 17, 26) {real, imag} */,
  {32'hc42241ba, 32'h00000000} /* (31, 17, 25) {real, imag} */,
  {32'hc4324dab, 32'h00000000} /* (31, 17, 24) {real, imag} */,
  {32'hc3e5472f, 32'h00000000} /* (31, 17, 23) {real, imag} */,
  {32'hc422b03f, 32'h00000000} /* (31, 17, 22) {real, imag} */,
  {32'h42e1f960, 32'h00000000} /* (31, 17, 21) {real, imag} */,
  {32'h45042c19, 32'h00000000} /* (31, 17, 20) {real, imag} */,
  {32'h44a27726, 32'h00000000} /* (31, 17, 19) {real, imag} */,
  {32'h44cf50f1, 32'h00000000} /* (31, 17, 18) {real, imag} */,
  {32'h44c55da7, 32'h00000000} /* (31, 17, 17) {real, imag} */,
  {32'h44a46d9b, 32'h00000000} /* (31, 17, 16) {real, imag} */,
  {32'h44d9b9d0, 32'h00000000} /* (31, 17, 15) {real, imag} */,
  {32'h44d6e18e, 32'h00000000} /* (31, 17, 14) {real, imag} */,
  {32'h448c220c, 32'h00000000} /* (31, 17, 13) {real, imag} */,
  {32'h448d0f1a, 32'h00000000} /* (31, 17, 12) {real, imag} */,
  {32'h4431872a, 32'h00000000} /* (31, 17, 11) {real, imag} */,
  {32'hc40fcdde, 32'h00000000} /* (31, 17, 10) {real, imag} */,
  {32'hc4b14749, 32'h00000000} /* (31, 17, 9) {real, imag} */,
  {32'hc4dddea0, 32'h00000000} /* (31, 17, 8) {real, imag} */,
  {32'hc4a6cbfa, 32'h00000000} /* (31, 17, 7) {real, imag} */,
  {32'hc4a5a07a, 32'h00000000} /* (31, 17, 6) {real, imag} */,
  {32'hc4db55d0, 32'h00000000} /* (31, 17, 5) {real, imag} */,
  {32'hc4bb8484, 32'h00000000} /* (31, 17, 4) {real, imag} */,
  {32'hc4e7ba5e, 32'h00000000} /* (31, 17, 3) {real, imag} */,
  {32'hc4c9e033, 32'h00000000} /* (31, 17, 2) {real, imag} */,
  {32'hc5148b3c, 32'h00000000} /* (31, 17, 1) {real, imag} */,
  {32'hc4d4d00d, 32'h00000000} /* (31, 17, 0) {real, imag} */,
  {32'hc493b536, 32'h00000000} /* (31, 16, 31) {real, imag} */,
  {32'hc4bd6c4a, 32'h00000000} /* (31, 16, 30) {real, imag} */,
  {32'hc4c0f51a, 32'h00000000} /* (31, 16, 29) {real, imag} */,
  {32'hc4506f5a, 32'h00000000} /* (31, 16, 28) {real, imag} */,
  {32'hc43cc857, 32'h00000000} /* (31, 16, 27) {real, imag} */,
  {32'hc4588824, 32'h00000000} /* (31, 16, 26) {real, imag} */,
  {32'hc47ca324, 32'h00000000} /* (31, 16, 25) {real, imag} */,
  {32'hc43695ec, 32'h00000000} /* (31, 16, 24) {real, imag} */,
  {32'hc4476077, 32'h00000000} /* (31, 16, 23) {real, imag} */,
  {32'hc42dfd2a, 32'h00000000} /* (31, 16, 22) {real, imag} */,
  {32'h418365e0, 32'h00000000} /* (31, 16, 21) {real, imag} */,
  {32'h4497f3e3, 32'h00000000} /* (31, 16, 20) {real, imag} */,
  {32'h44889a3a, 32'h00000000} /* (31, 16, 19) {real, imag} */,
  {32'h44955710, 32'h00000000} /* (31, 16, 18) {real, imag} */,
  {32'h44a6118c, 32'h00000000} /* (31, 16, 17) {real, imag} */,
  {32'h44c84a77, 32'h00000000} /* (31, 16, 16) {real, imag} */,
  {32'h44a1fbb2, 32'h00000000} /* (31, 16, 15) {real, imag} */,
  {32'h44b4d2d0, 32'h00000000} /* (31, 16, 14) {real, imag} */,
  {32'h44b90aa4, 32'h00000000} /* (31, 16, 13) {real, imag} */,
  {32'h44cd64c5, 32'h00000000} /* (31, 16, 12) {real, imag} */,
  {32'hc2ff3c78, 32'h00000000} /* (31, 16, 11) {real, imag} */,
  {32'hc4875d61, 32'h00000000} /* (31, 16, 10) {real, imag} */,
  {32'hc4e3bb3a, 32'h00000000} /* (31, 16, 9) {real, imag} */,
  {32'hc4cf72ae, 32'h00000000} /* (31, 16, 8) {real, imag} */,
  {32'hc4ab6aac, 32'h00000000} /* (31, 16, 7) {real, imag} */,
  {32'hc511fd28, 32'h00000000} /* (31, 16, 6) {real, imag} */,
  {32'hc4f09eac, 32'h00000000} /* (31, 16, 5) {real, imag} */,
  {32'hc4dc8cf7, 32'h00000000} /* (31, 16, 4) {real, imag} */,
  {32'hc4c152ec, 32'h00000000} /* (31, 16, 3) {real, imag} */,
  {32'hc4c6603a, 32'h00000000} /* (31, 16, 2) {real, imag} */,
  {32'hc4f94416, 32'h00000000} /* (31, 16, 1) {real, imag} */,
  {32'hc4e58a5b, 32'h00000000} /* (31, 16, 0) {real, imag} */,
  {32'hc4decd64, 32'h00000000} /* (31, 15, 31) {real, imag} */,
  {32'hc4bf1908, 32'h00000000} /* (31, 15, 30) {real, imag} */,
  {32'hc4de29b8, 32'h00000000} /* (31, 15, 29) {real, imag} */,
  {32'hc463494c, 32'h00000000} /* (31, 15, 28) {real, imag} */,
  {32'hc43f49b4, 32'h00000000} /* (31, 15, 27) {real, imag} */,
  {32'hc447ab52, 32'h00000000} /* (31, 15, 26) {real, imag} */,
  {32'hc42a9a17, 32'h00000000} /* (31, 15, 25) {real, imag} */,
  {32'hc46cb436, 32'h00000000} /* (31, 15, 24) {real, imag} */,
  {32'hc4a406e1, 32'h00000000} /* (31, 15, 23) {real, imag} */,
  {32'hc39adc46, 32'h00000000} /* (31, 15, 22) {real, imag} */,
  {32'h411510c0, 32'h00000000} /* (31, 15, 21) {real, imag} */,
  {32'h43b1fe70, 32'h00000000} /* (31, 15, 20) {real, imag} */,
  {32'h4464f8c8, 32'h00000000} /* (31, 15, 19) {real, imag} */,
  {32'h44755f19, 32'h00000000} /* (31, 15, 18) {real, imag} */,
  {32'h444e62dd, 32'h00000000} /* (31, 15, 17) {real, imag} */,
  {32'h4483d60c, 32'h00000000} /* (31, 15, 16) {real, imag} */,
  {32'h44c38e5a, 32'h00000000} /* (31, 15, 15) {real, imag} */,
  {32'h44a79c28, 32'h00000000} /* (31, 15, 14) {real, imag} */,
  {32'h44a0cbe0, 32'h00000000} /* (31, 15, 13) {real, imag} */,
  {32'h4418d548, 32'h00000000} /* (31, 15, 12) {real, imag} */,
  {32'hc2b22edc, 32'h00000000} /* (31, 15, 11) {real, imag} */,
  {32'hc4992bf4, 32'h00000000} /* (31, 15, 10) {real, imag} */,
  {32'hc4c55628, 32'h00000000} /* (31, 15, 9) {real, imag} */,
  {32'hc49782c9, 32'h00000000} /* (31, 15, 8) {real, imag} */,
  {32'hc4f1fc3f, 32'h00000000} /* (31, 15, 7) {real, imag} */,
  {32'hc4fe3dea, 32'h00000000} /* (31, 15, 6) {real, imag} */,
  {32'hc4c3d0a0, 32'h00000000} /* (31, 15, 5) {real, imag} */,
  {32'hc50ae154, 32'h00000000} /* (31, 15, 4) {real, imag} */,
  {32'hc4afefd6, 32'h00000000} /* (31, 15, 3) {real, imag} */,
  {32'hc4bde5e2, 32'h00000000} /* (31, 15, 2) {real, imag} */,
  {32'hc4f164f4, 32'h00000000} /* (31, 15, 1) {real, imag} */,
  {32'hc4636fd5, 32'h00000000} /* (31, 15, 0) {real, imag} */,
  {32'hc48b928c, 32'h00000000} /* (31, 14, 31) {real, imag} */,
  {32'hc4d06802, 32'h00000000} /* (31, 14, 30) {real, imag} */,
  {32'hc4bfce6a, 32'h00000000} /* (31, 14, 29) {real, imag} */,
  {32'hc4a1a424, 32'h00000000} /* (31, 14, 28) {real, imag} */,
  {32'hc4a9b42d, 32'h00000000} /* (31, 14, 27) {real, imag} */,
  {32'hc46a6876, 32'h00000000} /* (31, 14, 26) {real, imag} */,
  {32'hc49b1d06, 32'h00000000} /* (31, 14, 25) {real, imag} */,
  {32'hc4640d4e, 32'h00000000} /* (31, 14, 24) {real, imag} */,
  {32'hc4318ae4, 32'h00000000} /* (31, 14, 23) {real, imag} */,
  {32'hc4845fd3, 32'h00000000} /* (31, 14, 22) {real, imag} */,
  {32'hc3c39550, 32'h00000000} /* (31, 14, 21) {real, imag} */,
  {32'h4458340e, 32'h00000000} /* (31, 14, 20) {real, imag} */,
  {32'h44152b56, 32'h00000000} /* (31, 14, 19) {real, imag} */,
  {32'h442c3fac, 32'h00000000} /* (31, 14, 18) {real, imag} */,
  {32'h4487c137, 32'h00000000} /* (31, 14, 17) {real, imag} */,
  {32'h44854140, 32'h00000000} /* (31, 14, 16) {real, imag} */,
  {32'h44aa9424, 32'h00000000} /* (31, 14, 15) {real, imag} */,
  {32'h44186399, 32'h00000000} /* (31, 14, 14) {real, imag} */,
  {32'hc1d66880, 32'h00000000} /* (31, 14, 13) {real, imag} */,
  {32'h431c1d98, 32'h00000000} /* (31, 14, 12) {real, imag} */,
  {32'hc39b17e4, 32'h00000000} /* (31, 14, 11) {real, imag} */,
  {32'hc487028b, 32'h00000000} /* (31, 14, 10) {real, imag} */,
  {32'hc4a9f0c0, 32'h00000000} /* (31, 14, 9) {real, imag} */,
  {32'hc4edfea5, 32'h00000000} /* (31, 14, 8) {real, imag} */,
  {32'hc4ba1778, 32'h00000000} /* (31, 14, 7) {real, imag} */,
  {32'hc4b390d1, 32'h00000000} /* (31, 14, 6) {real, imag} */,
  {32'hc504a7bf, 32'h00000000} /* (31, 14, 5) {real, imag} */,
  {32'hc4bb7695, 32'h00000000} /* (31, 14, 4) {real, imag} */,
  {32'hc4affb2d, 32'h00000000} /* (31, 14, 3) {real, imag} */,
  {32'hc4974d7c, 32'h00000000} /* (31, 14, 2) {real, imag} */,
  {32'hc4446b5e, 32'h00000000} /* (31, 14, 1) {real, imag} */,
  {32'hc47696f3, 32'h00000000} /* (31, 14, 0) {real, imag} */,
  {32'hc479e231, 32'h00000000} /* (31, 13, 31) {real, imag} */,
  {32'hc4a65208, 32'h00000000} /* (31, 13, 30) {real, imag} */,
  {32'hc4966c6e, 32'h00000000} /* (31, 13, 29) {real, imag} */,
  {32'hc43f7b59, 32'h00000000} /* (31, 13, 28) {real, imag} */,
  {32'hc4414128, 32'h00000000} /* (31, 13, 27) {real, imag} */,
  {32'hc49f2371, 32'h00000000} /* (31, 13, 26) {real, imag} */,
  {32'hc4a5bbd1, 32'h00000000} /* (31, 13, 25) {real, imag} */,
  {32'hc4caf77c, 32'h00000000} /* (31, 13, 24) {real, imag} */,
  {32'hc48b7637, 32'h00000000} /* (31, 13, 23) {real, imag} */,
  {32'hc4a92ee2, 32'h00000000} /* (31, 13, 22) {real, imag} */,
  {32'hc406e075, 32'h00000000} /* (31, 13, 21) {real, imag} */,
  {32'h43c80490, 32'h00000000} /* (31, 13, 20) {real, imag} */,
  {32'h441b29b4, 32'h00000000} /* (31, 13, 19) {real, imag} */,
  {32'h442493fb, 32'h00000000} /* (31, 13, 18) {real, imag} */,
  {32'h445ffe57, 32'h00000000} /* (31, 13, 17) {real, imag} */,
  {32'h44556e80, 32'h00000000} /* (31, 13, 16) {real, imag} */,
  {32'h44b0e68a, 32'h00000000} /* (31, 13, 15) {real, imag} */,
  {32'h44569e71, 32'h00000000} /* (31, 13, 14) {real, imag} */,
  {32'h4443701b, 32'h00000000} /* (31, 13, 13) {real, imag} */,
  {32'h43943fc2, 32'h00000000} /* (31, 13, 12) {real, imag} */,
  {32'hc419698a, 32'h00000000} /* (31, 13, 11) {real, imag} */,
  {32'hc4088b1c, 32'h00000000} /* (31, 13, 10) {real, imag} */,
  {32'hc4d9a673, 32'h00000000} /* (31, 13, 9) {real, imag} */,
  {32'hc529fc4e, 32'h00000000} /* (31, 13, 8) {real, imag} */,
  {32'hc4ea6c75, 32'h00000000} /* (31, 13, 7) {real, imag} */,
  {32'hc4dfad7a, 32'h00000000} /* (31, 13, 6) {real, imag} */,
  {32'hc4e0b448, 32'h00000000} /* (31, 13, 5) {real, imag} */,
  {32'hc49eccb8, 32'h00000000} /* (31, 13, 4) {real, imag} */,
  {32'hc49b0f5d, 32'h00000000} /* (31, 13, 3) {real, imag} */,
  {32'hc4b7e23c, 32'h00000000} /* (31, 13, 2) {real, imag} */,
  {32'hc485e16c, 32'h00000000} /* (31, 13, 1) {real, imag} */,
  {32'hc46d40dc, 32'h00000000} /* (31, 13, 0) {real, imag} */,
  {32'hc47803f3, 32'h00000000} /* (31, 12, 31) {real, imag} */,
  {32'hc4ad53ff, 32'h00000000} /* (31, 12, 30) {real, imag} */,
  {32'hc430a6df, 32'h00000000} /* (31, 12, 29) {real, imag} */,
  {32'hc462ba86, 32'h00000000} /* (31, 12, 28) {real, imag} */,
  {32'hc4a190be, 32'h00000000} /* (31, 12, 27) {real, imag} */,
  {32'hc5039f3a, 32'h00000000} /* (31, 12, 26) {real, imag} */,
  {32'hc437aaf5, 32'h00000000} /* (31, 12, 25) {real, imag} */,
  {32'hc489b30c, 32'h00000000} /* (31, 12, 24) {real, imag} */,
  {32'hc4c2cb4e, 32'h00000000} /* (31, 12, 23) {real, imag} */,
  {32'hc4b87800, 32'h00000000} /* (31, 12, 22) {real, imag} */,
  {32'hc3fe1021, 32'h00000000} /* (31, 12, 21) {real, imag} */,
  {32'hc25d2e90, 32'h00000000} /* (31, 12, 20) {real, imag} */,
  {32'h43ce8667, 32'h00000000} /* (31, 12, 19) {real, imag} */,
  {32'h43e1066e, 32'h00000000} /* (31, 12, 18) {real, imag} */,
  {32'h444b513a, 32'h00000000} /* (31, 12, 17) {real, imag} */,
  {32'h44cd9363, 32'h00000000} /* (31, 12, 16) {real, imag} */,
  {32'h44250441, 32'h00000000} /* (31, 12, 15) {real, imag} */,
  {32'h44606fba, 32'h00000000} /* (31, 12, 14) {real, imag} */,
  {32'h43dfd166, 32'h00000000} /* (31, 12, 13) {real, imag} */,
  {32'h443a65a2, 32'h00000000} /* (31, 12, 12) {real, imag} */,
  {32'h43631c20, 32'h00000000} /* (31, 12, 11) {real, imag} */,
  {32'hc47d4576, 32'h00000000} /* (31, 12, 10) {real, imag} */,
  {32'hc4c80b72, 32'h00000000} /* (31, 12, 9) {real, imag} */,
  {32'hc517884c, 32'h00000000} /* (31, 12, 8) {real, imag} */,
  {32'hc49fb7f2, 32'h00000000} /* (31, 12, 7) {real, imag} */,
  {32'hc4dc2f72, 32'h00000000} /* (31, 12, 6) {real, imag} */,
  {32'hc4984590, 32'h00000000} /* (31, 12, 5) {real, imag} */,
  {32'hc48566d2, 32'h00000000} /* (31, 12, 4) {real, imag} */,
  {32'hc48dd923, 32'h00000000} /* (31, 12, 3) {real, imag} */,
  {32'hc446eb61, 32'h00000000} /* (31, 12, 2) {real, imag} */,
  {32'hc4cc6177, 32'h00000000} /* (31, 12, 1) {real, imag} */,
  {32'hc4914adf, 32'h00000000} /* (31, 12, 0) {real, imag} */,
  {32'hc38c4546, 32'h00000000} /* (31, 11, 31) {real, imag} */,
  {32'hc47cb954, 32'h00000000} /* (31, 11, 30) {real, imag} */,
  {32'hc40fb72c, 32'h00000000} /* (31, 11, 29) {real, imag} */,
  {32'hc423e852, 32'h00000000} /* (31, 11, 28) {real, imag} */,
  {32'hc4ac5547, 32'h00000000} /* (31, 11, 27) {real, imag} */,
  {32'hc3dd51ca, 32'h00000000} /* (31, 11, 26) {real, imag} */,
  {32'hc40e5c9a, 32'h00000000} /* (31, 11, 25) {real, imag} */,
  {32'hc43cfbfd, 32'h00000000} /* (31, 11, 24) {real, imag} */,
  {32'hc435ea86, 32'h00000000} /* (31, 11, 23) {real, imag} */,
  {32'hc495089c, 32'h00000000} /* (31, 11, 22) {real, imag} */,
  {32'hc402ad50, 32'h00000000} /* (31, 11, 21) {real, imag} */,
  {32'h43e5c4ec, 32'h00000000} /* (31, 11, 20) {real, imag} */,
  {32'h43200db4, 32'h00000000} /* (31, 11, 19) {real, imag} */,
  {32'h4419cb37, 32'h00000000} /* (31, 11, 18) {real, imag} */,
  {32'h44c69a0b, 32'h00000000} /* (31, 11, 17) {real, imag} */,
  {32'h44169943, 32'h00000000} /* (31, 11, 16) {real, imag} */,
  {32'h42f9e4fa, 32'h00000000} /* (31, 11, 15) {real, imag} */,
  {32'h44118d3a, 32'h00000000} /* (31, 11, 14) {real, imag} */,
  {32'hc38927fa, 32'h00000000} /* (31, 11, 13) {real, imag} */,
  {32'h43d7dd2c, 32'h00000000} /* (31, 11, 12) {real, imag} */,
  {32'h42b40fd0, 32'h00000000} /* (31, 11, 11) {real, imag} */,
  {32'hc463b11d, 32'h00000000} /* (31, 11, 10) {real, imag} */,
  {32'hc4644066, 32'h00000000} /* (31, 11, 9) {real, imag} */,
  {32'hc451c4ef, 32'h00000000} /* (31, 11, 8) {real, imag} */,
  {32'hc3e909d4, 32'h00000000} /* (31, 11, 7) {real, imag} */,
  {32'hc34b2d90, 32'h00000000} /* (31, 11, 6) {real, imag} */,
  {32'hc4a1e73c, 32'h00000000} /* (31, 11, 5) {real, imag} */,
  {32'hc3c57dc8, 32'h00000000} /* (31, 11, 4) {real, imag} */,
  {32'hc412c780, 32'h00000000} /* (31, 11, 3) {real, imag} */,
  {32'hc42a1a5f, 32'h00000000} /* (31, 11, 2) {real, imag} */,
  {32'hc3429aa8, 32'h00000000} /* (31, 11, 1) {real, imag} */,
  {32'hc311ceec, 32'h00000000} /* (31, 11, 0) {real, imag} */,
  {32'h44850ba4, 32'h00000000} /* (31, 10, 31) {real, imag} */,
  {32'h44663217, 32'h00000000} /* (31, 10, 30) {real, imag} */,
  {32'hc341cc62, 32'h00000000} /* (31, 10, 29) {real, imag} */,
  {32'hc1a26848, 32'h00000000} /* (31, 10, 28) {real, imag} */,
  {32'hc2fab624, 32'h00000000} /* (31, 10, 27) {real, imag} */,
  {32'hc2cc04bb, 32'h00000000} /* (31, 10, 26) {real, imag} */,
  {32'h441d2155, 32'h00000000} /* (31, 10, 25) {real, imag} */,
  {32'hc24ff358, 32'h00000000} /* (31, 10, 24) {real, imag} */,
  {32'h44429d5e, 32'h00000000} /* (31, 10, 23) {real, imag} */,
  {32'hc3e280f3, 32'h00000000} /* (31, 10, 22) {real, imag} */,
  {32'h40d365c0, 32'h00000000} /* (31, 10, 21) {real, imag} */,
  {32'hc3adb5df, 32'h00000000} /* (31, 10, 20) {real, imag} */,
  {32'hc4183b38, 32'h00000000} /* (31, 10, 19) {real, imag} */,
  {32'hc3828896, 32'h00000000} /* (31, 10, 18) {real, imag} */,
  {32'hc26896e0, 32'h00000000} /* (31, 10, 17) {real, imag} */,
  {32'hc387873c, 32'h00000000} /* (31, 10, 16) {real, imag} */,
  {32'hc522d34e, 32'h00000000} /* (31, 10, 15) {real, imag} */,
  {32'hc47bd719, 32'h00000000} /* (31, 10, 14) {real, imag} */,
  {32'hc48a27b6, 32'h00000000} /* (31, 10, 13) {real, imag} */,
  {32'hc3e4dcb4, 32'h00000000} /* (31, 10, 12) {real, imag} */,
  {32'hc3602b92, 32'h00000000} /* (31, 10, 11) {real, imag} */,
  {32'hc2a97513, 32'h00000000} /* (31, 10, 10) {real, imag} */,
  {32'h4409dc8d, 32'h00000000} /* (31, 10, 9) {real, imag} */,
  {32'h443cbcbe, 32'h00000000} /* (31, 10, 8) {real, imag} */,
  {32'h445d374c, 32'h00000000} /* (31, 10, 7) {real, imag} */,
  {32'h43e62925, 32'h00000000} /* (31, 10, 6) {real, imag} */,
  {32'h444d3eb6, 32'h00000000} /* (31, 10, 5) {real, imag} */,
  {32'h441ec150, 32'h00000000} /* (31, 10, 4) {real, imag} */,
  {32'h42734458, 32'h00000000} /* (31, 10, 3) {real, imag} */,
  {32'h4403d5ac, 32'h00000000} /* (31, 10, 2) {real, imag} */,
  {32'h4374f948, 32'h00000000} /* (31, 10, 1) {real, imag} */,
  {32'h42e087c6, 32'h00000000} /* (31, 10, 0) {real, imag} */,
  {32'h44c459ce, 32'h00000000} /* (31, 9, 31) {real, imag} */,
  {32'h449b5cb1, 32'h00000000} /* (31, 9, 30) {real, imag} */,
  {32'h43b73278, 32'h00000000} /* (31, 9, 29) {real, imag} */,
  {32'h43b90ae1, 32'h00000000} /* (31, 9, 28) {real, imag} */,
  {32'h43f21baa, 32'h00000000} /* (31, 9, 27) {real, imag} */,
  {32'h447750a3, 32'h00000000} /* (31, 9, 26) {real, imag} */,
  {32'h445a288a, 32'h00000000} /* (31, 9, 25) {real, imag} */,
  {32'h4480bc99, 32'h00000000} /* (31, 9, 24) {real, imag} */,
  {32'h43ac8244, 32'h00000000} /* (31, 9, 23) {real, imag} */,
  {32'h44aaee26, 32'h00000000} /* (31, 9, 22) {real, imag} */,
  {32'hc31047d4, 32'h00000000} /* (31, 9, 21) {real, imag} */,
  {32'hc38eed8c, 32'h00000000} /* (31, 9, 20) {real, imag} */,
  {32'hc4367ca6, 32'h00000000} /* (31, 9, 19) {real, imag} */,
  {32'hc49cf340, 32'h00000000} /* (31, 9, 18) {real, imag} */,
  {32'hc499e7c3, 32'h00000000} /* (31, 9, 17) {real, imag} */,
  {32'hc499bbe4, 32'h00000000} /* (31, 9, 16) {real, imag} */,
  {32'hc4d0a8a2, 32'h00000000} /* (31, 9, 15) {real, imag} */,
  {32'hc4b7b033, 32'h00000000} /* (31, 9, 14) {real, imag} */,
  {32'hc4aae096, 32'h00000000} /* (31, 9, 13) {real, imag} */,
  {32'hc48aa828, 32'h00000000} /* (31, 9, 12) {real, imag} */,
  {32'hc46b7de9, 32'h00000000} /* (31, 9, 11) {real, imag} */,
  {32'hc3546a2c, 32'h00000000} /* (31, 9, 10) {real, imag} */,
  {32'h445be53e, 32'h00000000} /* (31, 9, 9) {real, imag} */,
  {32'h44a57995, 32'h00000000} /* (31, 9, 8) {real, imag} */,
  {32'h44b4da77, 32'h00000000} /* (31, 9, 7) {real, imag} */,
  {32'h4468c078, 32'h00000000} /* (31, 9, 6) {real, imag} */,
  {32'h448ddba8, 32'h00000000} /* (31, 9, 5) {real, imag} */,
  {32'h44fda9ed, 32'h00000000} /* (31, 9, 4) {real, imag} */,
  {32'h448ebe72, 32'h00000000} /* (31, 9, 3) {real, imag} */,
  {32'h4466c6f9, 32'h00000000} /* (31, 9, 2) {real, imag} */,
  {32'h448af173, 32'h00000000} /* (31, 9, 1) {real, imag} */,
  {32'h4402b3fc, 32'h00000000} /* (31, 9, 0) {real, imag} */,
  {32'h4451f23e, 32'h00000000} /* (31, 8, 31) {real, imag} */,
  {32'h44748fea, 32'h00000000} /* (31, 8, 30) {real, imag} */,
  {32'h443449d3, 32'h00000000} /* (31, 8, 29) {real, imag} */,
  {32'h44420382, 32'h00000000} /* (31, 8, 28) {real, imag} */,
  {32'h4494e4c0, 32'h00000000} /* (31, 8, 27) {real, imag} */,
  {32'h44b1c330, 32'h00000000} /* (31, 8, 26) {real, imag} */,
  {32'h449a92fb, 32'h00000000} /* (31, 8, 25) {real, imag} */,
  {32'h44b8f8cc, 32'h00000000} /* (31, 8, 24) {real, imag} */,
  {32'h43fc0a53, 32'h00000000} /* (31, 8, 23) {real, imag} */,
  {32'h43856c10, 32'h00000000} /* (31, 8, 22) {real, imag} */,
  {32'hc2011878, 32'h00000000} /* (31, 8, 21) {real, imag} */,
  {32'hc4902770, 32'h00000000} /* (31, 8, 20) {real, imag} */,
  {32'hc46e0908, 32'h00000000} /* (31, 8, 19) {real, imag} */,
  {32'hc486ed2a, 32'h00000000} /* (31, 8, 18) {real, imag} */,
  {32'hc4c53860, 32'h00000000} /* (31, 8, 17) {real, imag} */,
  {32'hc48548a3, 32'h00000000} /* (31, 8, 16) {real, imag} */,
  {32'hc49db58d, 32'h00000000} /* (31, 8, 15) {real, imag} */,
  {32'hc498f5a7, 32'h00000000} /* (31, 8, 14) {real, imag} */,
  {32'hc4c03f1e, 32'h00000000} /* (31, 8, 13) {real, imag} */,
  {32'hc4f1f97f, 32'h00000000} /* (31, 8, 12) {real, imag} */,
  {32'hc4918df4, 32'h00000000} /* (31, 8, 11) {real, imag} */,
  {32'hc421db3f, 32'h00000000} /* (31, 8, 10) {real, imag} */,
  {32'h4461f14b, 32'h00000000} /* (31, 8, 9) {real, imag} */,
  {32'h4421ffb0, 32'h00000000} /* (31, 8, 8) {real, imag} */,
  {32'h44ae63df, 32'h00000000} /* (31, 8, 7) {real, imag} */,
  {32'h44b459cc, 32'h00000000} /* (31, 8, 6) {real, imag} */,
  {32'h445e127e, 32'h00000000} /* (31, 8, 5) {real, imag} */,
  {32'h44bcdd3e, 32'h00000000} /* (31, 8, 4) {real, imag} */,
  {32'h44a6e060, 32'h00000000} /* (31, 8, 3) {real, imag} */,
  {32'h44931ff0, 32'h00000000} /* (31, 8, 2) {real, imag} */,
  {32'h44ac4278, 32'h00000000} /* (31, 8, 1) {real, imag} */,
  {32'h448ed85f, 32'h00000000} /* (31, 8, 0) {real, imag} */,
  {32'h44bdde72, 32'h00000000} /* (31, 7, 31) {real, imag} */,
  {32'h44ad9146, 32'h00000000} /* (31, 7, 30) {real, imag} */,
  {32'h446e7298, 32'h00000000} /* (31, 7, 29) {real, imag} */,
  {32'h4441729e, 32'h00000000} /* (31, 7, 28) {real, imag} */,
  {32'h44428878, 32'h00000000} /* (31, 7, 27) {real, imag} */,
  {32'h43cd934b, 32'h00000000} /* (31, 7, 26) {real, imag} */,
  {32'h440ce764, 32'h00000000} /* (31, 7, 25) {real, imag} */,
  {32'h44010189, 32'h00000000} /* (31, 7, 24) {real, imag} */,
  {32'h443dd3c8, 32'h00000000} /* (31, 7, 23) {real, imag} */,
  {32'h43b63f54, 32'h00000000} /* (31, 7, 22) {real, imag} */,
  {32'hc4039fb9, 32'h00000000} /* (31, 7, 21) {real, imag} */,
  {32'hc4c6a8e4, 32'h00000000} /* (31, 7, 20) {real, imag} */,
  {32'hc3c59988, 32'h00000000} /* (31, 7, 19) {real, imag} */,
  {32'hc41c6aae, 32'h00000000} /* (31, 7, 18) {real, imag} */,
  {32'hc44e6664, 32'h00000000} /* (31, 7, 17) {real, imag} */,
  {32'hc47fdc3e, 32'h00000000} /* (31, 7, 16) {real, imag} */,
  {32'hc4d6c956, 32'h00000000} /* (31, 7, 15) {real, imag} */,
  {32'hc4d7acf6, 32'h00000000} /* (31, 7, 14) {real, imag} */,
  {32'hc4a89cee, 32'h00000000} /* (31, 7, 13) {real, imag} */,
  {32'hc4ccf20d, 32'h00000000} /* (31, 7, 12) {real, imag} */,
  {32'hc4fdf910, 32'h00000000} /* (31, 7, 11) {real, imag} */,
  {32'h42dfb784, 32'h00000000} /* (31, 7, 10) {real, imag} */,
  {32'h4402ba6c, 32'h00000000} /* (31, 7, 9) {real, imag} */,
  {32'h443c2a37, 32'h00000000} /* (31, 7, 8) {real, imag} */,
  {32'h4506b77c, 32'h00000000} /* (31, 7, 7) {real, imag} */,
  {32'h449d39af, 32'h00000000} /* (31, 7, 6) {real, imag} */,
  {32'h44b13cb6, 32'h00000000} /* (31, 7, 5) {real, imag} */,
  {32'h44b2100a, 32'h00000000} /* (31, 7, 4) {real, imag} */,
  {32'h44c1f214, 32'h00000000} /* (31, 7, 3) {real, imag} */,
  {32'h44c27559, 32'h00000000} /* (31, 7, 2) {real, imag} */,
  {32'h4480822f, 32'h00000000} /* (31, 7, 1) {real, imag} */,
  {32'h44815f65, 32'h00000000} /* (31, 7, 0) {real, imag} */,
  {32'h44bd2276, 32'h00000000} /* (31, 6, 31) {real, imag} */,
  {32'h442fe8a3, 32'h00000000} /* (31, 6, 30) {real, imag} */,
  {32'h4435494b, 32'h00000000} /* (31, 6, 29) {real, imag} */,
  {32'h4450a858, 32'h00000000} /* (31, 6, 28) {real, imag} */,
  {32'h434c46c8, 32'h00000000} /* (31, 6, 27) {real, imag} */,
  {32'h43663354, 32'h00000000} /* (31, 6, 26) {real, imag} */,
  {32'h43e53eb1, 32'h00000000} /* (31, 6, 25) {real, imag} */,
  {32'h444f4e60, 32'h00000000} /* (31, 6, 24) {real, imag} */,
  {32'h43f537c2, 32'h00000000} /* (31, 6, 23) {real, imag} */,
  {32'h44881239, 32'h00000000} /* (31, 6, 22) {real, imag} */,
  {32'h43aa3632, 32'h00000000} /* (31, 6, 21) {real, imag} */,
  {32'hc451ed68, 32'h00000000} /* (31, 6, 20) {real, imag} */,
  {32'hc3a2b8ea, 32'h00000000} /* (31, 6, 19) {real, imag} */,
  {32'hc48bc553, 32'h00000000} /* (31, 6, 18) {real, imag} */,
  {32'hc5022dde, 32'h00000000} /* (31, 6, 17) {real, imag} */,
  {32'hc48d34d8, 32'h00000000} /* (31, 6, 16) {real, imag} */,
  {32'hc4871cfa, 32'h00000000} /* (31, 6, 15) {real, imag} */,
  {32'hc4c81888, 32'h00000000} /* (31, 6, 14) {real, imag} */,
  {32'hc4ec1842, 32'h00000000} /* (31, 6, 13) {real, imag} */,
  {32'hc49d6a4a, 32'h00000000} /* (31, 6, 12) {real, imag} */,
  {32'hc4ce4079, 32'h00000000} /* (31, 6, 11) {real, imag} */,
  {32'hc4202418, 32'h00000000} /* (31, 6, 10) {real, imag} */,
  {32'hc24bdb30, 32'h00000000} /* (31, 6, 9) {real, imag} */,
  {32'h440a526c, 32'h00000000} /* (31, 6, 8) {real, imag} */,
  {32'h44e91798, 32'h00000000} /* (31, 6, 7) {real, imag} */,
  {32'h45032cb4, 32'h00000000} /* (31, 6, 6) {real, imag} */,
  {32'h44b94e38, 32'h00000000} /* (31, 6, 5) {real, imag} */,
  {32'h44bfb588, 32'h00000000} /* (31, 6, 4) {real, imag} */,
  {32'h44d187ae, 32'h00000000} /* (31, 6, 3) {real, imag} */,
  {32'h4498cf09, 32'h00000000} /* (31, 6, 2) {real, imag} */,
  {32'h44ddb0fd, 32'h00000000} /* (31, 6, 1) {real, imag} */,
  {32'h4452d3ae, 32'h00000000} /* (31, 6, 0) {real, imag} */,
  {32'h449a3906, 32'h00000000} /* (31, 5, 31) {real, imag} */,
  {32'h43e4b0fc, 32'h00000000} /* (31, 5, 30) {real, imag} */,
  {32'h449259e1, 32'h00000000} /* (31, 5, 29) {real, imag} */,
  {32'h44de6b42, 32'h00000000} /* (31, 5, 28) {real, imag} */,
  {32'h4327e310, 32'h00000000} /* (31, 5, 27) {real, imag} */,
  {32'h44493c35, 32'h00000000} /* (31, 5, 26) {real, imag} */,
  {32'h4386278e, 32'h00000000} /* (31, 5, 25) {real, imag} */,
  {32'h442c47c0, 32'h00000000} /* (31, 5, 24) {real, imag} */,
  {32'h449cda1b, 32'h00000000} /* (31, 5, 23) {real, imag} */,
  {32'h4461d77c, 32'h00000000} /* (31, 5, 22) {real, imag} */,
  {32'h448ad0d0, 32'h00000000} /* (31, 5, 21) {real, imag} */,
  {32'h438bb330, 32'h00000000} /* (31, 5, 20) {real, imag} */,
  {32'h435333b4, 32'h00000000} /* (31, 5, 19) {real, imag} */,
  {32'hc30f3e44, 32'h00000000} /* (31, 5, 18) {real, imag} */,
  {32'hc4898fb9, 32'h00000000} /* (31, 5, 17) {real, imag} */,
  {32'hc47dc41c, 32'h00000000} /* (31, 5, 16) {real, imag} */,
  {32'hc46104df, 32'h00000000} /* (31, 5, 15) {real, imag} */,
  {32'hc4be0a27, 32'h00000000} /* (31, 5, 14) {real, imag} */,
  {32'hc4e0d33f, 32'h00000000} /* (31, 5, 13) {real, imag} */,
  {32'hc4a4eff6, 32'h00000000} /* (31, 5, 12) {real, imag} */,
  {32'hc4bcfcab, 32'h00000000} /* (31, 5, 11) {real, imag} */,
  {32'hc4b54f12, 32'h00000000} /* (31, 5, 10) {real, imag} */,
  {32'hc469c899, 32'h00000000} /* (31, 5, 9) {real, imag} */,
  {32'hc3fb22cc, 32'h00000000} /* (31, 5, 8) {real, imag} */,
  {32'h43e3c6ff, 32'h00000000} /* (31, 5, 7) {real, imag} */,
  {32'h44872722, 32'h00000000} /* (31, 5, 6) {real, imag} */,
  {32'h44037358, 32'h00000000} /* (31, 5, 5) {real, imag} */,
  {32'h44d07248, 32'h00000000} /* (31, 5, 4) {real, imag} */,
  {32'h44ab9294, 32'h00000000} /* (31, 5, 3) {real, imag} */,
  {32'h445c70f3, 32'h00000000} /* (31, 5, 2) {real, imag} */,
  {32'h44a80493, 32'h00000000} /* (31, 5, 1) {real, imag} */,
  {32'h43903ae3, 32'h00000000} /* (31, 5, 0) {real, imag} */,
  {32'h43eb39a0, 32'h00000000} /* (31, 4, 31) {real, imag} */,
  {32'h42b2e818, 32'h00000000} /* (31, 4, 30) {real, imag} */,
  {32'hc129a780, 32'h00000000} /* (31, 4, 29) {real, imag} */,
  {32'h445e2e9e, 32'h00000000} /* (31, 4, 28) {real, imag} */,
  {32'h4440ca81, 32'h00000000} /* (31, 4, 27) {real, imag} */,
  {32'h445aa5d4, 32'h00000000} /* (31, 4, 26) {real, imag} */,
  {32'h43bcd4b8, 32'h00000000} /* (31, 4, 25) {real, imag} */,
  {32'h43b5fb6a, 32'h00000000} /* (31, 4, 24) {real, imag} */,
  {32'h43cf6ba4, 32'h00000000} /* (31, 4, 23) {real, imag} */,
  {32'h445c25a8, 32'h00000000} /* (31, 4, 22) {real, imag} */,
  {32'h443e97a4, 32'h00000000} /* (31, 4, 21) {real, imag} */,
  {32'h442e8a48, 32'h00000000} /* (31, 4, 20) {real, imag} */,
  {32'h4426bdb4, 32'h00000000} /* (31, 4, 19) {real, imag} */,
  {32'h42895b80, 32'h00000000} /* (31, 4, 18) {real, imag} */,
  {32'h43395a7e, 32'h00000000} /* (31, 4, 17) {real, imag} */,
  {32'hc41441ed, 32'h00000000} /* (31, 4, 16) {real, imag} */,
  {32'hc4a627c2, 32'h00000000} /* (31, 4, 15) {real, imag} */,
  {32'hc49b2666, 32'h00000000} /* (31, 4, 14) {real, imag} */,
  {32'hc4a78bf1, 32'h00000000} /* (31, 4, 13) {real, imag} */,
  {32'hc4a0f76f, 32'h00000000} /* (31, 4, 12) {real, imag} */,
  {32'hc5154570, 32'h00000000} /* (31, 4, 11) {real, imag} */,
  {32'hc4f682fe, 32'h00000000} /* (31, 4, 10) {real, imag} */,
  {32'hc4835729, 32'h00000000} /* (31, 4, 9) {real, imag} */,
  {32'hc4029a36, 32'h00000000} /* (31, 4, 8) {real, imag} */,
  {32'hc3cdeb28, 32'h00000000} /* (31, 4, 7) {real, imag} */,
  {32'hc3f9cbdb, 32'h00000000} /* (31, 4, 6) {real, imag} */,
  {32'h4443284c, 32'h00000000} /* (31, 4, 5) {real, imag} */,
  {32'h44673830, 32'h00000000} /* (31, 4, 4) {real, imag} */,
  {32'h443a67e6, 32'h00000000} /* (31, 4, 3) {real, imag} */,
  {32'h448d03c6, 32'h00000000} /* (31, 4, 2) {real, imag} */,
  {32'h448ee20f, 32'h00000000} /* (31, 4, 1) {real, imag} */,
  {32'h44669d1f, 32'h00000000} /* (31, 4, 0) {real, imag} */,
  {32'h4407ec94, 32'h00000000} /* (31, 3, 31) {real, imag} */,
  {32'h444cda68, 32'h00000000} /* (31, 3, 30) {real, imag} */,
  {32'h43d76e76, 32'h00000000} /* (31, 3, 29) {real, imag} */,
  {32'h44666533, 32'h00000000} /* (31, 3, 28) {real, imag} */,
  {32'h44347faa, 32'h00000000} /* (31, 3, 27) {real, imag} */,
  {32'h447394ed, 32'h00000000} /* (31, 3, 26) {real, imag} */,
  {32'h4480a4e4, 32'h00000000} /* (31, 3, 25) {real, imag} */,
  {32'h448b90a3, 32'h00000000} /* (31, 3, 24) {real, imag} */,
  {32'h44993c48, 32'h00000000} /* (31, 3, 23) {real, imag} */,
  {32'h448ef4ed, 32'h00000000} /* (31, 3, 22) {real, imag} */,
  {32'h445e2c1b, 32'h00000000} /* (31, 3, 21) {real, imag} */,
  {32'h445c5fc8, 32'h00000000} /* (31, 3, 20) {real, imag} */,
  {32'h4465835f, 32'h00000000} /* (31, 3, 19) {real, imag} */,
  {32'h4380cf94, 32'h00000000} /* (31, 3, 18) {real, imag} */,
  {32'h424cc6b0, 32'h00000000} /* (31, 3, 17) {real, imag} */,
  {32'hc4004bee, 32'h00000000} /* (31, 3, 16) {real, imag} */,
  {32'hc4812e14, 32'h00000000} /* (31, 3, 15) {real, imag} */,
  {32'hc4dc89a8, 32'h00000000} /* (31, 3, 14) {real, imag} */,
  {32'hc4f0b10e, 32'h00000000} /* (31, 3, 13) {real, imag} */,
  {32'hc4d16694, 32'h00000000} /* (31, 3, 12) {real, imag} */,
  {32'hc4ddc4a3, 32'h00000000} /* (31, 3, 11) {real, imag} */,
  {32'hc52ae747, 32'h00000000} /* (31, 3, 10) {real, imag} */,
  {32'hc48a4894, 32'h00000000} /* (31, 3, 9) {real, imag} */,
  {32'hc46918c2, 32'h00000000} /* (31, 3, 8) {real, imag} */,
  {32'hc4421e39, 32'h00000000} /* (31, 3, 7) {real, imag} */,
  {32'hc407762c, 32'h00000000} /* (31, 3, 6) {real, imag} */,
  {32'hc416166d, 32'h00000000} /* (31, 3, 5) {real, imag} */,
  {32'h44116c66, 32'h00000000} /* (31, 3, 4) {real, imag} */,
  {32'h4452d74d, 32'h00000000} /* (31, 3, 3) {real, imag} */,
  {32'h4483e624, 32'h00000000} /* (31, 3, 2) {real, imag} */,
  {32'h44b15c58, 32'h00000000} /* (31, 3, 1) {real, imag} */,
  {32'h43c6b6ea, 32'h00000000} /* (31, 3, 0) {real, imag} */,
  {32'h43c1fc14, 32'h00000000} /* (31, 2, 31) {real, imag} */,
  {32'h44414afd, 32'h00000000} /* (31, 2, 30) {real, imag} */,
  {32'h44654340, 32'h00000000} /* (31, 2, 29) {real, imag} */,
  {32'h43575bec, 32'h00000000} /* (31, 2, 28) {real, imag} */,
  {32'h4493ec1b, 32'h00000000} /* (31, 2, 27) {real, imag} */,
  {32'h44889a2a, 32'h00000000} /* (31, 2, 26) {real, imag} */,
  {32'h441c9ed8, 32'h00000000} /* (31, 2, 25) {real, imag} */,
  {32'h4439a3dc, 32'h00000000} /* (31, 2, 24) {real, imag} */,
  {32'h444cf2b7, 32'h00000000} /* (31, 2, 23) {real, imag} */,
  {32'h4469f3cf, 32'h00000000} /* (31, 2, 22) {real, imag} */,
  {32'h44717938, 32'h00000000} /* (31, 2, 21) {real, imag} */,
  {32'h4492cebe, 32'h00000000} /* (31, 2, 20) {real, imag} */,
  {32'h443386ca, 32'h00000000} /* (31, 2, 19) {real, imag} */,
  {32'h42920e70, 32'h00000000} /* (31, 2, 18) {real, imag} */,
  {32'hc38a4d60, 32'h00000000} /* (31, 2, 17) {real, imag} */,
  {32'hc3d292f2, 32'h00000000} /* (31, 2, 16) {real, imag} */,
  {32'hc4d0b4e9, 32'h00000000} /* (31, 2, 15) {real, imag} */,
  {32'hc48ef966, 32'h00000000} /* (31, 2, 14) {real, imag} */,
  {32'hc4bff4ee, 32'h00000000} /* (31, 2, 13) {real, imag} */,
  {32'hc4e05ebe, 32'h00000000} /* (31, 2, 12) {real, imag} */,
  {32'hc4ce89f3, 32'h00000000} /* (31, 2, 11) {real, imag} */,
  {32'hc4ae422e, 32'h00000000} /* (31, 2, 10) {real, imag} */,
  {32'hc4b3233a, 32'h00000000} /* (31, 2, 9) {real, imag} */,
  {32'hc46aaa40, 32'h00000000} /* (31, 2, 8) {real, imag} */,
  {32'hc4b15bca, 32'h00000000} /* (31, 2, 7) {real, imag} */,
  {32'hc4b638b4, 32'h00000000} /* (31, 2, 6) {real, imag} */,
  {32'hc40788fe, 32'h00000000} /* (31, 2, 5) {real, imag} */,
  {32'h4348e9cc, 32'h00000000} /* (31, 2, 4) {real, imag} */,
  {32'h448afcb9, 32'h00000000} /* (31, 2, 3) {real, imag} */,
  {32'h442ffad5, 32'h00000000} /* (31, 2, 2) {real, imag} */,
  {32'h43bb93ea, 32'h00000000} /* (31, 2, 1) {real, imag} */,
  {32'h43d11e4a, 32'h00000000} /* (31, 2, 0) {real, imag} */,
  {32'h435eba0e, 32'h00000000} /* (31, 1, 31) {real, imag} */,
  {32'h440dc1d7, 32'h00000000} /* (31, 1, 30) {real, imag} */,
  {32'h420bd4e4, 32'h00000000} /* (31, 1, 29) {real, imag} */,
  {32'h440fd1a7, 32'h00000000} /* (31, 1, 28) {real, imag} */,
  {32'h4498aea3, 32'h00000000} /* (31, 1, 27) {real, imag} */,
  {32'h444bd772, 32'h00000000} /* (31, 1, 26) {real, imag} */,
  {32'h44628ca4, 32'h00000000} /* (31, 1, 25) {real, imag} */,
  {32'h44da2da8, 32'h00000000} /* (31, 1, 24) {real, imag} */,
  {32'h4461cd20, 32'h00000000} /* (31, 1, 23) {real, imag} */,
  {32'h4471a1e0, 32'h00000000} /* (31, 1, 22) {real, imag} */,
  {32'h446fa238, 32'h00000000} /* (31, 1, 21) {real, imag} */,
  {32'h4479e401, 32'h00000000} /* (31, 1, 20) {real, imag} */,
  {32'h43fd8af4, 32'h00000000} /* (31, 1, 19) {real, imag} */,
  {32'h4340993e, 32'h00000000} /* (31, 1, 18) {real, imag} */,
  {32'hc2a5e062, 32'h00000000} /* (31, 1, 17) {real, imag} */,
  {32'hc3f3e15a, 32'h00000000} /* (31, 1, 16) {real, imag} */,
  {32'hc47c3b42, 32'h00000000} /* (31, 1, 15) {real, imag} */,
  {32'hc49d5258, 32'h00000000} /* (31, 1, 14) {real, imag} */,
  {32'hc3c353de, 32'h00000000} /* (31, 1, 13) {real, imag} */,
  {32'hc4774ded, 32'h00000000} /* (31, 1, 12) {real, imag} */,
  {32'hc4a162c7, 32'h00000000} /* (31, 1, 11) {real, imag} */,
  {32'hc4dccfdb, 32'h00000000} /* (31, 1, 10) {real, imag} */,
  {32'hc499ecb4, 32'h00000000} /* (31, 1, 9) {real, imag} */,
  {32'hc4733fcf, 32'h00000000} /* (31, 1, 8) {real, imag} */,
  {32'hc45906ea, 32'h00000000} /* (31, 1, 7) {real, imag} */,
  {32'hc49b94fe, 32'h00000000} /* (31, 1, 6) {real, imag} */,
  {32'h43407510, 32'h00000000} /* (31, 1, 5) {real, imag} */,
  {32'h43713c14, 32'h00000000} /* (31, 1, 4) {real, imag} */,
  {32'h44171ff2, 32'h00000000} /* (31, 1, 3) {real, imag} */,
  {32'h4424d18a, 32'h00000000} /* (31, 1, 2) {real, imag} */,
  {32'h42fbbb7a, 32'h00000000} /* (31, 1, 1) {real, imag} */,
  {32'h427b8df0, 32'h00000000} /* (31, 1, 0) {real, imag} */,
  {32'h43826886, 32'h00000000} /* (31, 0, 31) {real, imag} */,
  {32'h429ee038, 32'h00000000} /* (31, 0, 30) {real, imag} */,
  {32'h43146f3c, 32'h00000000} /* (31, 0, 29) {real, imag} */,
  {32'h433cd9bc, 32'h00000000} /* (31, 0, 28) {real, imag} */,
  {32'h43ac4e1f, 32'h00000000} /* (31, 0, 27) {real, imag} */,
  {32'h44390f20, 32'h00000000} /* (31, 0, 26) {real, imag} */,
  {32'h4489f6a6, 32'h00000000} /* (31, 0, 25) {real, imag} */,
  {32'h44645c6a, 32'h00000000} /* (31, 0, 24) {real, imag} */,
  {32'h4498670a, 32'h00000000} /* (31, 0, 23) {real, imag} */,
  {32'h4491fe7a, 32'h00000000} /* (31, 0, 22) {real, imag} */,
  {32'h4452ac94, 32'h00000000} /* (31, 0, 21) {real, imag} */,
  {32'h442b0909, 32'h00000000} /* (31, 0, 20) {real, imag} */,
  {32'h441d2260, 32'h00000000} /* (31, 0, 19) {real, imag} */,
  {32'h4011c880, 32'h00000000} /* (31, 0, 18) {real, imag} */,
  {32'hc33bb6a4, 32'h00000000} /* (31, 0, 17) {real, imag} */,
  {32'hc3da9bfa, 32'h00000000} /* (31, 0, 16) {real, imag} */,
  {32'hc4980614, 32'h00000000} /* (31, 0, 15) {real, imag} */,
  {32'hc4aff6f6, 32'h00000000} /* (31, 0, 14) {real, imag} */,
  {32'hc49d8aee, 32'h00000000} /* (31, 0, 13) {real, imag} */,
  {32'hc46f0635, 32'h00000000} /* (31, 0, 12) {real, imag} */,
  {32'hc42bed9e, 32'h00000000} /* (31, 0, 11) {real, imag} */,
  {32'hc49fa2a6, 32'h00000000} /* (31, 0, 10) {real, imag} */,
  {32'hc3d25915, 32'h00000000} /* (31, 0, 9) {real, imag} */,
  {32'hc40fb168, 32'h00000000} /* (31, 0, 8) {real, imag} */,
  {32'hc3824f1e, 32'h00000000} /* (31, 0, 7) {real, imag} */,
  {32'h421450f0, 32'h00000000} /* (31, 0, 6) {real, imag} */,
  {32'h420d2cf0, 32'h00000000} /* (31, 0, 5) {real, imag} */,
  {32'h4406c539, 32'h00000000} /* (31, 0, 4) {real, imag} */,
  {32'h4364194c, 32'h00000000} /* (31, 0, 3) {real, imag} */,
  {32'h4392824f, 32'h00000000} /* (31, 0, 2) {real, imag} */,
  {32'h43731c40, 32'h00000000} /* (31, 0, 1) {real, imag} */,
  {32'h42d346b8, 32'h00000000} /* (31, 0, 0) {real, imag} */,
  {32'h44851126, 32'h00000000} /* (30, 31, 31) {real, imag} */,
  {32'h448f0376, 32'h00000000} /* (30, 31, 30) {real, imag} */,
  {32'h44e3d04e, 32'h00000000} /* (30, 31, 29) {real, imag} */,
  {32'h44c1972a, 32'h00000000} /* (30, 31, 28) {real, imag} */,
  {32'h44d13684, 32'h00000000} /* (30, 31, 27) {real, imag} */,
  {32'h44ba9dac, 32'h00000000} /* (30, 31, 26) {real, imag} */,
  {32'h454aead1, 32'h00000000} /* (30, 31, 25) {real, imag} */,
  {32'h4518937e, 32'h00000000} /* (30, 31, 24) {real, imag} */,
  {32'h44e4daf4, 32'h00000000} /* (30, 31, 23) {real, imag} */,
  {32'h44da55f7, 32'h00000000} /* (30, 31, 22) {real, imag} */,
  {32'h44d3c24a, 32'h00000000} /* (30, 31, 21) {real, imag} */,
  {32'h43c5e5f2, 32'h00000000} /* (30, 31, 20) {real, imag} */,
  {32'hc3111ff8, 32'h00000000} /* (30, 31, 19) {real, imag} */,
  {32'hc3bbb2ea, 32'h00000000} /* (30, 31, 18) {real, imag} */,
  {32'hc481c874, 32'h00000000} /* (30, 31, 17) {real, imag} */,
  {32'hc5025021, 32'h00000000} /* (30, 31, 16) {real, imag} */,
  {32'hc501a774, 32'h00000000} /* (30, 31, 15) {real, imag} */,
  {32'hc527862f, 32'h00000000} /* (30, 31, 14) {real, imag} */,
  {32'hc54ad0df, 32'h00000000} /* (30, 31, 13) {real, imag} */,
  {32'hc5329fc1, 32'h00000000} /* (30, 31, 12) {real, imag} */,
  {32'hc5123603, 32'h00000000} /* (30, 31, 11) {real, imag} */,
  {32'hc47dc7b9, 32'h00000000} /* (30, 31, 10) {real, imag} */,
  {32'hc2d8d8e0, 32'h00000000} /* (30, 31, 9) {real, imag} */,
  {32'h4414a45e, 32'h00000000} /* (30, 31, 8) {real, imag} */,
  {32'h43d8b470, 32'h00000000} /* (30, 31, 7) {real, imag} */,
  {32'h44676292, 32'h00000000} /* (30, 31, 6) {real, imag} */,
  {32'h44ab0c0a, 32'h00000000} /* (30, 31, 5) {real, imag} */,
  {32'h44c2bba0, 32'h00000000} /* (30, 31, 4) {real, imag} */,
  {32'h44c9b22c, 32'h00000000} /* (30, 31, 3) {real, imag} */,
  {32'h44ee2154, 32'h00000000} /* (30, 31, 2) {real, imag} */,
  {32'h44cbf1a0, 32'h00000000} /* (30, 31, 1) {real, imag} */,
  {32'h44a249e8, 32'h00000000} /* (30, 31, 0) {real, imag} */,
  {32'h44c8be00, 32'h00000000} /* (30, 30, 31) {real, imag} */,
  {32'h450a5e08, 32'h00000000} /* (30, 30, 30) {real, imag} */,
  {32'h4510fffc, 32'h00000000} /* (30, 30, 29) {real, imag} */,
  {32'h44eed660, 32'h00000000} /* (30, 30, 28) {real, imag} */,
  {32'h4508cd56, 32'h00000000} /* (30, 30, 27) {real, imag} */,
  {32'h453ccfb8, 32'h00000000} /* (30, 30, 26) {real, imag} */,
  {32'h4572c051, 32'h00000000} /* (30, 30, 25) {real, imag} */,
  {32'h455f8bff, 32'h00000000} /* (30, 30, 24) {real, imag} */,
  {32'h454214e5, 32'h00000000} /* (30, 30, 23) {real, imag} */,
  {32'h45093b4c, 32'h00000000} /* (30, 30, 22) {real, imag} */,
  {32'h45127cb0, 32'h00000000} /* (30, 30, 21) {real, imag} */,
  {32'h43b3a8d0, 32'h00000000} /* (30, 30, 20) {real, imag} */,
  {32'hc45b86a9, 32'h00000000} /* (30, 30, 19) {real, imag} */,
  {32'hc4db5bf0, 32'h00000000} /* (30, 30, 18) {real, imag} */,
  {32'hc50454c1, 32'h00000000} /* (30, 30, 17) {real, imag} */,
  {32'hc5128734, 32'h00000000} /* (30, 30, 16) {real, imag} */,
  {32'hc5410b08, 32'h00000000} /* (30, 30, 15) {real, imag} */,
  {32'hc576d1b6, 32'h00000000} /* (30, 30, 14) {real, imag} */,
  {32'hc5a1ba11, 32'h00000000} /* (30, 30, 13) {real, imag} */,
  {32'hc5792cac, 32'h00000000} /* (30, 30, 12) {real, imag} */,
  {32'hc4fed974, 32'h00000000} /* (30, 30, 11) {real, imag} */,
  {32'hc3750208, 32'h00000000} /* (30, 30, 10) {real, imag} */,
  {32'h448b7f42, 32'h00000000} /* (30, 30, 9) {real, imag} */,
  {32'h44d5e57a, 32'h00000000} /* (30, 30, 8) {real, imag} */,
  {32'h44a762ea, 32'h00000000} /* (30, 30, 7) {real, imag} */,
  {32'h44edbaaf, 32'h00000000} /* (30, 30, 6) {real, imag} */,
  {32'h45142efe, 32'h00000000} /* (30, 30, 5) {real, imag} */,
  {32'h4547e5fc, 32'h00000000} /* (30, 30, 4) {real, imag} */,
  {32'h4520a4ad, 32'h00000000} /* (30, 30, 3) {real, imag} */,
  {32'h4502742b, 32'h00000000} /* (30, 30, 2) {real, imag} */,
  {32'h453dd3a3, 32'h00000000} /* (30, 30, 1) {real, imag} */,
  {32'h45126b42, 32'h00000000} /* (30, 30, 0) {real, imag} */,
  {32'h44af2aa0, 32'h00000000} /* (30, 29, 31) {real, imag} */,
  {32'h451beb62, 32'h00000000} /* (30, 29, 30) {real, imag} */,
  {32'h4522c75c, 32'h00000000} /* (30, 29, 29) {real, imag} */,
  {32'h4506af47, 32'h00000000} /* (30, 29, 28) {real, imag} */,
  {32'h450925c4, 32'h00000000} /* (30, 29, 27) {real, imag} */,
  {32'h450698fe, 32'h00000000} /* (30, 29, 26) {real, imag} */,
  {32'h453c1373, 32'h00000000} /* (30, 29, 25) {real, imag} */,
  {32'h4560f479, 32'h00000000} /* (30, 29, 24) {real, imag} */,
  {32'h452d8b16, 32'h00000000} /* (30, 29, 23) {real, imag} */,
  {32'h451b8c21, 32'h00000000} /* (30, 29, 22) {real, imag} */,
  {32'h445978fe, 32'h00000000} /* (30, 29, 21) {real, imag} */,
  {32'hc4953bcd, 32'h00000000} /* (30, 29, 20) {real, imag} */,
  {32'hc4bdbf60, 32'h00000000} /* (30, 29, 19) {real, imag} */,
  {32'hc4f9687a, 32'h00000000} /* (30, 29, 18) {real, imag} */,
  {32'hc528227f, 32'h00000000} /* (30, 29, 17) {real, imag} */,
  {32'hc5770157, 32'h00000000} /* (30, 29, 16) {real, imag} */,
  {32'hc559a464, 32'h00000000} /* (30, 29, 15) {real, imag} */,
  {32'hc57ee122, 32'h00000000} /* (30, 29, 14) {real, imag} */,
  {32'hc5730708, 32'h00000000} /* (30, 29, 13) {real, imag} */,
  {32'hc5467883, 32'h00000000} /* (30, 29, 12) {real, imag} */,
  {32'hc506d2fe, 32'h00000000} /* (30, 29, 11) {real, imag} */,
  {32'hc417da8a, 32'h00000000} /* (30, 29, 10) {real, imag} */,
  {32'h44eeebc2, 32'h00000000} /* (30, 29, 9) {real, imag} */,
  {32'h45014341, 32'h00000000} /* (30, 29, 8) {real, imag} */,
  {32'h44f10f9c, 32'h00000000} /* (30, 29, 7) {real, imag} */,
  {32'h4504c31b, 32'h00000000} /* (30, 29, 6) {real, imag} */,
  {32'h454324cc, 32'h00000000} /* (30, 29, 5) {real, imag} */,
  {32'h4522b1b2, 32'h00000000} /* (30, 29, 4) {real, imag} */,
  {32'h4559d5c8, 32'h00000000} /* (30, 29, 3) {real, imag} */,
  {32'h4509f43b, 32'h00000000} /* (30, 29, 2) {real, imag} */,
  {32'h44eba3a2, 32'h00000000} /* (30, 29, 1) {real, imag} */,
  {32'h44e755ca, 32'h00000000} /* (30, 29, 0) {real, imag} */,
  {32'h44ae7ec0, 32'h00000000} /* (30, 28, 31) {real, imag} */,
  {32'h45445f43, 32'h00000000} /* (30, 28, 30) {real, imag} */,
  {32'h457d1966, 32'h00000000} /* (30, 28, 29) {real, imag} */,
  {32'h450327a6, 32'h00000000} /* (30, 28, 28) {real, imag} */,
  {32'h4525e044, 32'h00000000} /* (30, 28, 27) {real, imag} */,
  {32'h45640194, 32'h00000000} /* (30, 28, 26) {real, imag} */,
  {32'h454f24c1, 32'h00000000} /* (30, 28, 25) {real, imag} */,
  {32'h4535e067, 32'h00000000} /* (30, 28, 24) {real, imag} */,
  {32'h44ffd43c, 32'h00000000} /* (30, 28, 23) {real, imag} */,
  {32'h44b4df22, 32'h00000000} /* (30, 28, 22) {real, imag} */,
  {32'h433e1dd8, 32'h00000000} /* (30, 28, 21) {real, imag} */,
  {32'hc4e43626, 32'h00000000} /* (30, 28, 20) {real, imag} */,
  {32'hc521aa28, 32'h00000000} /* (30, 28, 19) {real, imag} */,
  {32'hc51b39e8, 32'h00000000} /* (30, 28, 18) {real, imag} */,
  {32'hc52eed1b, 32'h00000000} /* (30, 28, 17) {real, imag} */,
  {32'hc539a0c4, 32'h00000000} /* (30, 28, 16) {real, imag} */,
  {32'hc5398d6e, 32'h00000000} /* (30, 28, 15) {real, imag} */,
  {32'hc5764bb1, 32'h00000000} /* (30, 28, 14) {real, imag} */,
  {32'hc554154e, 32'h00000000} /* (30, 28, 13) {real, imag} */,
  {32'hc5018d10, 32'h00000000} /* (30, 28, 12) {real, imag} */,
  {32'hc4c74d57, 32'h00000000} /* (30, 28, 11) {real, imag} */,
  {32'h43d93410, 32'h00000000} /* (30, 28, 10) {real, imag} */,
  {32'h44b8ecae, 32'h00000000} /* (30, 28, 9) {real, imag} */,
  {32'h453bbb69, 32'h00000000} /* (30, 28, 8) {real, imag} */,
  {32'h451842ca, 32'h00000000} /* (30, 28, 7) {real, imag} */,
  {32'h45515ee5, 32'h00000000} /* (30, 28, 6) {real, imag} */,
  {32'h4523a8fa, 32'h00000000} /* (30, 28, 5) {real, imag} */,
  {32'h45258ab7, 32'h00000000} /* (30, 28, 4) {real, imag} */,
  {32'h452e2b5c, 32'h00000000} /* (30, 28, 3) {real, imag} */,
  {32'h450c5ba8, 32'h00000000} /* (30, 28, 2) {real, imag} */,
  {32'h44e57f82, 32'h00000000} /* (30, 28, 1) {real, imag} */,
  {32'h44d2168f, 32'h00000000} /* (30, 28, 0) {real, imag} */,
  {32'h451b2c1a, 32'h00000000} /* (30, 27, 31) {real, imag} */,
  {32'h451e7986, 32'h00000000} /* (30, 27, 30) {real, imag} */,
  {32'h45284ff2, 32'h00000000} /* (30, 27, 29) {real, imag} */,
  {32'h4506f5e6, 32'h00000000} /* (30, 27, 28) {real, imag} */,
  {32'h45307cd0, 32'h00000000} /* (30, 27, 27) {real, imag} */,
  {32'h458f810f, 32'h00000000} /* (30, 27, 26) {real, imag} */,
  {32'h454e14bc, 32'h00000000} /* (30, 27, 25) {real, imag} */,
  {32'h45168889, 32'h00000000} /* (30, 27, 24) {real, imag} */,
  {32'h4504cbaf, 32'h00000000} /* (30, 27, 23) {real, imag} */,
  {32'h44ca1318, 32'h00000000} /* (30, 27, 22) {real, imag} */,
  {32'h4499db3a, 32'h00000000} /* (30, 27, 21) {real, imag} */,
  {32'hc424d224, 32'h00000000} /* (30, 27, 20) {real, imag} */,
  {32'hc4dc5065, 32'h00000000} /* (30, 27, 19) {real, imag} */,
  {32'hc52e21d2, 32'h00000000} /* (30, 27, 18) {real, imag} */,
  {32'hc529f1a2, 32'h00000000} /* (30, 27, 17) {real, imag} */,
  {32'hc539cec3, 32'h00000000} /* (30, 27, 16) {real, imag} */,
  {32'hc55f8d1a, 32'h00000000} /* (30, 27, 15) {real, imag} */,
  {32'hc57aa638, 32'h00000000} /* (30, 27, 14) {real, imag} */,
  {32'hc584425f, 32'h00000000} /* (30, 27, 13) {real, imag} */,
  {32'hc4b5f982, 32'h00000000} /* (30, 27, 12) {real, imag} */,
  {32'hc4b2fc33, 32'h00000000} /* (30, 27, 11) {real, imag} */,
  {32'h44a10483, 32'h00000000} /* (30, 27, 10) {real, imag} */,
  {32'h4553fbec, 32'h00000000} /* (30, 27, 9) {real, imag} */,
  {32'h45443977, 32'h00000000} /* (30, 27, 8) {real, imag} */,
  {32'h4566097d, 32'h00000000} /* (30, 27, 7) {real, imag} */,
  {32'h453c7966, 32'h00000000} /* (30, 27, 6) {real, imag} */,
  {32'h452e4f66, 32'h00000000} /* (30, 27, 5) {real, imag} */,
  {32'h454f6109, 32'h00000000} /* (30, 27, 4) {real, imag} */,
  {32'h451f482b, 32'h00000000} /* (30, 27, 3) {real, imag} */,
  {32'h4517a742, 32'h00000000} /* (30, 27, 2) {real, imag} */,
  {32'h44ff617b, 32'h00000000} /* (30, 27, 1) {real, imag} */,
  {32'h44bbb9ee, 32'h00000000} /* (30, 27, 0) {real, imag} */,
  {32'h44dbdb3c, 32'h00000000} /* (30, 26, 31) {real, imag} */,
  {32'h4518c796, 32'h00000000} /* (30, 26, 30) {real, imag} */,
  {32'h45208ac0, 32'h00000000} /* (30, 26, 29) {real, imag} */,
  {32'h450bdc81, 32'h00000000} /* (30, 26, 28) {real, imag} */,
  {32'h4547283b, 32'h00000000} /* (30, 26, 27) {real, imag} */,
  {32'h4532873e, 32'h00000000} /* (30, 26, 26) {real, imag} */,
  {32'h454afa21, 32'h00000000} /* (30, 26, 25) {real, imag} */,
  {32'h45436210, 32'h00000000} /* (30, 26, 24) {real, imag} */,
  {32'h44f845f6, 32'h00000000} /* (30, 26, 23) {real, imag} */,
  {32'h44d7b91e, 32'h00000000} /* (30, 26, 22) {real, imag} */,
  {32'h445544a4, 32'h00000000} /* (30, 26, 21) {real, imag} */,
  {32'hc47f4260, 32'h00000000} /* (30, 26, 20) {real, imag} */,
  {32'hc4f7e838, 32'h00000000} /* (30, 26, 19) {real, imag} */,
  {32'hc50093fe, 32'h00000000} /* (30, 26, 18) {real, imag} */,
  {32'hc51a60ca, 32'h00000000} /* (30, 26, 17) {real, imag} */,
  {32'hc53747e1, 32'h00000000} /* (30, 26, 16) {real, imag} */,
  {32'hc5815073, 32'h00000000} /* (30, 26, 15) {real, imag} */,
  {32'hc5661c38, 32'h00000000} /* (30, 26, 14) {real, imag} */,
  {32'hc54d57fc, 32'h00000000} /* (30, 26, 13) {real, imag} */,
  {32'hc52b5ded, 32'h00000000} /* (30, 26, 12) {real, imag} */,
  {32'hc4bb9562, 32'h00000000} /* (30, 26, 11) {real, imag} */,
  {32'h44089096, 32'h00000000} /* (30, 26, 10) {real, imag} */,
  {32'h451352bb, 32'h00000000} /* (30, 26, 9) {real, imag} */,
  {32'h454934be, 32'h00000000} /* (30, 26, 8) {real, imag} */,
  {32'h45698ee9, 32'h00000000} /* (30, 26, 7) {real, imag} */,
  {32'h457ca215, 32'h00000000} /* (30, 26, 6) {real, imag} */,
  {32'h454639e2, 32'h00000000} /* (30, 26, 5) {real, imag} */,
  {32'h4528c6fa, 32'h00000000} /* (30, 26, 4) {real, imag} */,
  {32'h45724650, 32'h00000000} /* (30, 26, 3) {real, imag} */,
  {32'h454870a2, 32'h00000000} /* (30, 26, 2) {real, imag} */,
  {32'h450ba1ec, 32'h00000000} /* (30, 26, 1) {real, imag} */,
  {32'h44f04792, 32'h00000000} /* (30, 26, 0) {real, imag} */,
  {32'h44d9f136, 32'h00000000} /* (30, 25, 31) {real, imag} */,
  {32'h4542a492, 32'h00000000} /* (30, 25, 30) {real, imag} */,
  {32'h4517298b, 32'h00000000} /* (30, 25, 29) {real, imag} */,
  {32'h450766eb, 32'h00000000} /* (30, 25, 28) {real, imag} */,
  {32'h45641b3a, 32'h00000000} /* (30, 25, 27) {real, imag} */,
  {32'h4556fce2, 32'h00000000} /* (30, 25, 26) {real, imag} */,
  {32'h455ceae6, 32'h00000000} /* (30, 25, 25) {real, imag} */,
  {32'h4537d7d6, 32'h00000000} /* (30, 25, 24) {real, imag} */,
  {32'h450aaa49, 32'h00000000} /* (30, 25, 23) {real, imag} */,
  {32'h44dcae77, 32'h00000000} /* (30, 25, 22) {real, imag} */,
  {32'h44950514, 32'h00000000} /* (30, 25, 21) {real, imag} */,
  {32'hc4c01550, 32'h00000000} /* (30, 25, 20) {real, imag} */,
  {32'hc519d151, 32'h00000000} /* (30, 25, 19) {real, imag} */,
  {32'hc50fb084, 32'h00000000} /* (30, 25, 18) {real, imag} */,
  {32'hc562a022, 32'h00000000} /* (30, 25, 17) {real, imag} */,
  {32'hc56b872c, 32'h00000000} /* (30, 25, 16) {real, imag} */,
  {32'hc5650d03, 32'h00000000} /* (30, 25, 15) {real, imag} */,
  {32'hc596dc2f, 32'h00000000} /* (30, 25, 14) {real, imag} */,
  {32'hc55f0a91, 32'h00000000} /* (30, 25, 13) {real, imag} */,
  {32'hc53003d3, 32'h00000000} /* (30, 25, 12) {real, imag} */,
  {32'hc48305a0, 32'h00000000} /* (30, 25, 11) {real, imag} */,
  {32'h449dd884, 32'h00000000} /* (30, 25, 10) {real, imag} */,
  {32'h44f6f683, 32'h00000000} /* (30, 25, 9) {real, imag} */,
  {32'h454db8e4, 32'h00000000} /* (30, 25, 8) {real, imag} */,
  {32'h4564784d, 32'h00000000} /* (30, 25, 7) {real, imag} */,
  {32'h45560538, 32'h00000000} /* (30, 25, 6) {real, imag} */,
  {32'h45853b42, 32'h00000000} /* (30, 25, 5) {real, imag} */,
  {32'h4570ae1a, 32'h00000000} /* (30, 25, 4) {real, imag} */,
  {32'h453c7b57, 32'h00000000} /* (30, 25, 3) {real, imag} */,
  {32'h451dc8fa, 32'h00000000} /* (30, 25, 2) {real, imag} */,
  {32'h44c86771, 32'h00000000} /* (30, 25, 1) {real, imag} */,
  {32'h44b32c84, 32'h00000000} /* (30, 25, 0) {real, imag} */,
  {32'h450d8696, 32'h00000000} /* (30, 24, 31) {real, imag} */,
  {32'h452ee3ee, 32'h00000000} /* (30, 24, 30) {real, imag} */,
  {32'h4545247f, 32'h00000000} /* (30, 24, 29) {real, imag} */,
  {32'h450fa7b1, 32'h00000000} /* (30, 24, 28) {real, imag} */,
  {32'h44a6752e, 32'h00000000} /* (30, 24, 27) {real, imag} */,
  {32'h4549f234, 32'h00000000} /* (30, 24, 26) {real, imag} */,
  {32'h451ccf1e, 32'h00000000} /* (30, 24, 25) {real, imag} */,
  {32'h4508d72c, 32'h00000000} /* (30, 24, 24) {real, imag} */,
  {32'h4515720f, 32'h00000000} /* (30, 24, 23) {real, imag} */,
  {32'h451b097e, 32'h00000000} /* (30, 24, 22) {real, imag} */,
  {32'h44972f03, 32'h00000000} /* (30, 24, 21) {real, imag} */,
  {32'hc4f5cede, 32'h00000000} /* (30, 24, 20) {real, imag} */,
  {32'hc4eb6e16, 32'h00000000} /* (30, 24, 19) {real, imag} */,
  {32'hc50cb0d5, 32'h00000000} /* (30, 24, 18) {real, imag} */,
  {32'hc54197b7, 32'h00000000} /* (30, 24, 17) {real, imag} */,
  {32'hc558d524, 32'h00000000} /* (30, 24, 16) {real, imag} */,
  {32'hc540cd44, 32'h00000000} /* (30, 24, 15) {real, imag} */,
  {32'hc55cb2a0, 32'h00000000} /* (30, 24, 14) {real, imag} */,
  {32'hc541667d, 32'h00000000} /* (30, 24, 13) {real, imag} */,
  {32'hc4bfdfe2, 32'h00000000} /* (30, 24, 12) {real, imag} */,
  {32'hc467beb3, 32'h00000000} /* (30, 24, 11) {real, imag} */,
  {32'h441e55fe, 32'h00000000} /* (30, 24, 10) {real, imag} */,
  {32'h45137e24, 32'h00000000} /* (30, 24, 9) {real, imag} */,
  {32'h4554083c, 32'h00000000} /* (30, 24, 8) {real, imag} */,
  {32'h45670f31, 32'h00000000} /* (30, 24, 7) {real, imag} */,
  {32'h455319b2, 32'h00000000} /* (30, 24, 6) {real, imag} */,
  {32'h45803a54, 32'h00000000} /* (30, 24, 5) {real, imag} */,
  {32'h45451a61, 32'h00000000} /* (30, 24, 4) {real, imag} */,
  {32'h456ff245, 32'h00000000} /* (30, 24, 3) {real, imag} */,
  {32'h4552f211, 32'h00000000} /* (30, 24, 2) {real, imag} */,
  {32'h44ebc1ca, 32'h00000000} /* (30, 24, 1) {real, imag} */,
  {32'h44b4e21f, 32'h00000000} /* (30, 24, 0) {real, imag} */,
  {32'h44cabffd, 32'h00000000} /* (30, 23, 31) {real, imag} */,
  {32'h45114e5e, 32'h00000000} /* (30, 23, 30) {real, imag} */,
  {32'h44d0628c, 32'h00000000} /* (30, 23, 29) {real, imag} */,
  {32'h44e85f31, 32'h00000000} /* (30, 23, 28) {real, imag} */,
  {32'h44a76401, 32'h00000000} /* (30, 23, 27) {real, imag} */,
  {32'h44b2f0fe, 32'h00000000} /* (30, 23, 26) {real, imag} */,
  {32'h45009e93, 32'h00000000} /* (30, 23, 25) {real, imag} */,
  {32'h44f5e36d, 32'h00000000} /* (30, 23, 24) {real, imag} */,
  {32'h452a2d4c, 32'h00000000} /* (30, 23, 23) {real, imag} */,
  {32'h451fe842, 32'h00000000} /* (30, 23, 22) {real, imag} */,
  {32'h449cd56a, 32'h00000000} /* (30, 23, 21) {real, imag} */,
  {32'hc45b0448, 32'h00000000} /* (30, 23, 20) {real, imag} */,
  {32'hc4d46a17, 32'h00000000} /* (30, 23, 19) {real, imag} */,
  {32'hc5020b05, 32'h00000000} /* (30, 23, 18) {real, imag} */,
  {32'hc5056cb7, 32'h00000000} /* (30, 23, 17) {real, imag} */,
  {32'hc52a7ac1, 32'h00000000} /* (30, 23, 16) {real, imag} */,
  {32'hc514de42, 32'h00000000} /* (30, 23, 15) {real, imag} */,
  {32'hc535cac8, 32'h00000000} /* (30, 23, 14) {real, imag} */,
  {32'hc506b9d0, 32'h00000000} /* (30, 23, 13) {real, imag} */,
  {32'hc403b43a, 32'h00000000} /* (30, 23, 12) {real, imag} */,
  {32'hc437cf12, 32'h00000000} /* (30, 23, 11) {real, imag} */,
  {32'h4402e413, 32'h00000000} /* (30, 23, 10) {real, imag} */,
  {32'h44f65aee, 32'h00000000} /* (30, 23, 9) {real, imag} */,
  {32'h453889ae, 32'h00000000} /* (30, 23, 8) {real, imag} */,
  {32'h45417f38, 32'h00000000} /* (30, 23, 7) {real, imag} */,
  {32'h4529defa, 32'h00000000} /* (30, 23, 6) {real, imag} */,
  {32'h4541e7db, 32'h00000000} /* (30, 23, 5) {real, imag} */,
  {32'h45455c4f, 32'h00000000} /* (30, 23, 4) {real, imag} */,
  {32'h454102ea, 32'h00000000} /* (30, 23, 3) {real, imag} */,
  {32'h4540604f, 32'h00000000} /* (30, 23, 2) {real, imag} */,
  {32'h45121b55, 32'h00000000} /* (30, 23, 1) {real, imag} */,
  {32'h4518dcb9, 32'h00000000} /* (30, 23, 0) {real, imag} */,
  {32'h4403fdf4, 32'h00000000} /* (30, 22, 31) {real, imag} */,
  {32'h44b3cf64, 32'h00000000} /* (30, 22, 30) {real, imag} */,
  {32'h44af5d32, 32'h00000000} /* (30, 22, 29) {real, imag} */,
  {32'h440ac741, 32'h00000000} /* (30, 22, 28) {real, imag} */,
  {32'h43fb5cf9, 32'h00000000} /* (30, 22, 27) {real, imag} */,
  {32'h43fa0878, 32'h00000000} /* (30, 22, 26) {real, imag} */,
  {32'h44a1c2e0, 32'h00000000} /* (30, 22, 25) {real, imag} */,
  {32'h44b0f878, 32'h00000000} /* (30, 22, 24) {real, imag} */,
  {32'h45113602, 32'h00000000} /* (30, 22, 23) {real, imag} */,
  {32'h4533bec2, 32'h00000000} /* (30, 22, 22) {real, imag} */,
  {32'h447a84a7, 32'h00000000} /* (30, 22, 21) {real, imag} */,
  {32'hc35626e8, 32'h00000000} /* (30, 22, 20) {real, imag} */,
  {32'hc49b43fd, 32'h00000000} /* (30, 22, 19) {real, imag} */,
  {32'hc4cd4420, 32'h00000000} /* (30, 22, 18) {real, imag} */,
  {32'hc5044c19, 32'h00000000} /* (30, 22, 17) {real, imag} */,
  {32'hc50ae992, 32'h00000000} /* (30, 22, 16) {real, imag} */,
  {32'hc51a2b52, 32'h00000000} /* (30, 22, 15) {real, imag} */,
  {32'hc4cd5d0c, 32'h00000000} /* (30, 22, 14) {real, imag} */,
  {32'hc49b268c, 32'h00000000} /* (30, 22, 13) {real, imag} */,
  {32'hc42e7ded, 32'h00000000} /* (30, 22, 12) {real, imag} */,
  {32'hc429bc96, 32'h00000000} /* (30, 22, 11) {real, imag} */,
  {32'h44986b7b, 32'h00000000} /* (30, 22, 10) {real, imag} */,
  {32'h44d15ab6, 32'h00000000} /* (30, 22, 9) {real, imag} */,
  {32'h44bccfc0, 32'h00000000} /* (30, 22, 8) {real, imag} */,
  {32'h45208202, 32'h00000000} /* (30, 22, 7) {real, imag} */,
  {32'h44e6b1ed, 32'h00000000} /* (30, 22, 6) {real, imag} */,
  {32'h4521feda, 32'h00000000} /* (30, 22, 5) {real, imag} */,
  {32'h45448f2e, 32'h00000000} /* (30, 22, 4) {real, imag} */,
  {32'h4514cdb0, 32'h00000000} /* (30, 22, 3) {real, imag} */,
  {32'h4506edcc, 32'h00000000} /* (30, 22, 2) {real, imag} */,
  {32'h44c29536, 32'h00000000} /* (30, 22, 1) {real, imag} */,
  {32'h447c076a, 32'h00000000} /* (30, 22, 0) {real, imag} */,
  {32'hc374fe10, 32'h00000000} /* (30, 21, 31) {real, imag} */,
  {32'h416dbf80, 32'h00000000} /* (30, 21, 30) {real, imag} */,
  {32'hc3dabc92, 32'h00000000} /* (30, 21, 29) {real, imag} */,
  {32'hc400c60c, 32'h00000000} /* (30, 21, 28) {real, imag} */,
  {32'hc3d075fa, 32'h00000000} /* (30, 21, 27) {real, imag} */,
  {32'h438a6b14, 32'h00000000} /* (30, 21, 26) {real, imag} */,
  {32'h41974680, 32'h00000000} /* (30, 21, 25) {real, imag} */,
  {32'h42d4bdae, 32'h00000000} /* (30, 21, 24) {real, imag} */,
  {32'h443d0d9b, 32'h00000000} /* (30, 21, 23) {real, imag} */,
  {32'hc34c2130, 32'h00000000} /* (30, 21, 22) {real, imag} */,
  {32'hc30e7a58, 32'h00000000} /* (30, 21, 21) {real, imag} */,
  {32'hc3871e68, 32'h00000000} /* (30, 21, 20) {real, imag} */,
  {32'hc3d01e74, 32'h00000000} /* (30, 21, 19) {real, imag} */,
  {32'hc39cd44c, 32'h00000000} /* (30, 21, 18) {real, imag} */,
  {32'hc49326de, 32'h00000000} /* (30, 21, 17) {real, imag} */,
  {32'hc494be2e, 32'h00000000} /* (30, 21, 16) {real, imag} */,
  {32'hc452a7e4, 32'h00000000} /* (30, 21, 15) {real, imag} */,
  {32'hc395a43e, 32'h00000000} /* (30, 21, 14) {real, imag} */,
  {32'hc32e2fe8, 32'h00000000} /* (30, 21, 13) {real, imag} */,
  {32'hc3bd2477, 32'h00000000} /* (30, 21, 12) {real, imag} */,
  {32'h4467064d, 32'h00000000} /* (30, 21, 11) {real, imag} */,
  {32'h441542e0, 32'h00000000} /* (30, 21, 10) {real, imag} */,
  {32'h44c1d79c, 32'h00000000} /* (30, 21, 9) {real, imag} */,
  {32'h439e41e0, 32'h00000000} /* (30, 21, 8) {real, imag} */,
  {32'h43b0b82a, 32'h00000000} /* (30, 21, 7) {real, imag} */,
  {32'h445d1684, 32'h00000000} /* (30, 21, 6) {real, imag} */,
  {32'h4384ddb8, 32'h00000000} /* (30, 21, 5) {real, imag} */,
  {32'h44af7aa6, 32'h00000000} /* (30, 21, 4) {real, imag} */,
  {32'h442ec410, 32'h00000000} /* (30, 21, 3) {real, imag} */,
  {32'h4437a3dc, 32'h00000000} /* (30, 21, 2) {real, imag} */,
  {32'h43d9ba88, 32'h00000000} /* (30, 21, 1) {real, imag} */,
  {32'hc3675bc8, 32'h00000000} /* (30, 21, 0) {real, imag} */,
  {32'hc4974786, 32'h00000000} /* (30, 20, 31) {real, imag} */,
  {32'hc49c84dc, 32'h00000000} /* (30, 20, 30) {real, imag} */,
  {32'hc503fc17, 32'h00000000} /* (30, 20, 29) {real, imag} */,
  {32'hc4db10a8, 32'h00000000} /* (30, 20, 28) {real, imag} */,
  {32'hc4f44b3e, 32'h00000000} /* (30, 20, 27) {real, imag} */,
  {32'hc50291c5, 32'h00000000} /* (30, 20, 26) {real, imag} */,
  {32'hc499a253, 32'h00000000} /* (30, 20, 25) {real, imag} */,
  {32'hc54ea90d, 32'h00000000} /* (30, 20, 24) {real, imag} */,
  {32'hc4cbb31d, 32'h00000000} /* (30, 20, 23) {real, imag} */,
  {32'hc4ab4203, 32'h00000000} /* (30, 20, 22) {real, imag} */,
  {32'hc4447360, 32'h00000000} /* (30, 20, 21) {real, imag} */,
  {32'h43e200a0, 32'h00000000} /* (30, 20, 20) {real, imag} */,
  {32'h43dec474, 32'h00000000} /* (30, 20, 19) {real, imag} */,
  {32'h441f603b, 32'h00000000} /* (30, 20, 18) {real, imag} */,
  {32'h44c0a8fc, 32'h00000000} /* (30, 20, 17) {real, imag} */,
  {32'h448086f3, 32'h00000000} /* (30, 20, 16) {real, imag} */,
  {32'h44c0fb62, 32'h00000000} /* (30, 20, 15) {real, imag} */,
  {32'h44d680e0, 32'h00000000} /* (30, 20, 14) {real, imag} */,
  {32'h451f6e61, 32'h00000000} /* (30, 20, 13) {real, imag} */,
  {32'h4509a538, 32'h00000000} /* (30, 20, 12) {real, imag} */,
  {32'h447e4c7c, 32'h00000000} /* (30, 20, 11) {real, imag} */,
  {32'h4397abb6, 32'h00000000} /* (30, 20, 10) {real, imag} */,
  {32'hc3e66b73, 32'h00000000} /* (30, 20, 9) {real, imag} */,
  {32'hc506bd4f, 32'h00000000} /* (30, 20, 8) {real, imag} */,
  {32'hc515eff3, 32'h00000000} /* (30, 20, 7) {real, imag} */,
  {32'hc51d05e6, 32'h00000000} /* (30, 20, 6) {real, imag} */,
  {32'hc4cb82d6, 32'h00000000} /* (30, 20, 5) {real, imag} */,
  {32'hc525c492, 32'h00000000} /* (30, 20, 4) {real, imag} */,
  {32'hc50f5330, 32'h00000000} /* (30, 20, 3) {real, imag} */,
  {32'hc49c404c, 32'h00000000} /* (30, 20, 2) {real, imag} */,
  {32'hc4d43b42, 32'h00000000} /* (30, 20, 1) {real, imag} */,
  {32'hc4e03cfd, 32'h00000000} /* (30, 20, 0) {real, imag} */,
  {32'hc4f55273, 32'h00000000} /* (30, 19, 31) {real, imag} */,
  {32'hc52cf16a, 32'h00000000} /* (30, 19, 30) {real, imag} */,
  {32'hc51e34b0, 32'h00000000} /* (30, 19, 29) {real, imag} */,
  {32'hc5290c44, 32'h00000000} /* (30, 19, 28) {real, imag} */,
  {32'hc523b4d0, 32'h00000000} /* (30, 19, 27) {real, imag} */,
  {32'hc52558a4, 32'h00000000} /* (30, 19, 26) {real, imag} */,
  {32'hc51d1bbc, 32'h00000000} /* (30, 19, 25) {real, imag} */,
  {32'hc53b4a3c, 32'h00000000} /* (30, 19, 24) {real, imag} */,
  {32'hc5126d7c, 32'h00000000} /* (30, 19, 23) {real, imag} */,
  {32'hc4c10b40, 32'h00000000} /* (30, 19, 22) {real, imag} */,
  {32'hc495c3a2, 32'h00000000} /* (30, 19, 21) {real, imag} */,
  {32'h444f2c52, 32'h00000000} /* (30, 19, 20) {real, imag} */,
  {32'h44b5a982, 32'h00000000} /* (30, 19, 19) {real, imag} */,
  {32'h45196dce, 32'h00000000} /* (30, 19, 18) {real, imag} */,
  {32'h450e5230, 32'h00000000} /* (30, 19, 17) {real, imag} */,
  {32'h44f77638, 32'h00000000} /* (30, 19, 16) {real, imag} */,
  {32'h453904cc, 32'h00000000} /* (30, 19, 15) {real, imag} */,
  {32'h45335d32, 32'h00000000} /* (30, 19, 14) {real, imag} */,
  {32'h45512158, 32'h00000000} /* (30, 19, 13) {real, imag} */,
  {32'h45380d1a, 32'h00000000} /* (30, 19, 12) {real, imag} */,
  {32'h450beda6, 32'h00000000} /* (30, 19, 11) {real, imag} */,
  {32'h42eb81f0, 32'h00000000} /* (30, 19, 10) {real, imag} */,
  {32'hc523b920, 32'h00000000} /* (30, 19, 9) {real, imag} */,
  {32'hc5445b6a, 32'h00000000} /* (30, 19, 8) {real, imag} */,
  {32'hc55bf6bc, 32'h00000000} /* (30, 19, 7) {real, imag} */,
  {32'hc5651810, 32'h00000000} /* (30, 19, 6) {real, imag} */,
  {32'hc50ccec3, 32'h00000000} /* (30, 19, 5) {real, imag} */,
  {32'hc55a0b70, 32'h00000000} /* (30, 19, 4) {real, imag} */,
  {32'hc551f8d9, 32'h00000000} /* (30, 19, 3) {real, imag} */,
  {32'hc522d706, 32'h00000000} /* (30, 19, 2) {real, imag} */,
  {32'hc54aa1a0, 32'h00000000} /* (30, 19, 1) {real, imag} */,
  {32'hc518fd0e, 32'h00000000} /* (30, 19, 0) {real, imag} */,
  {32'hc5620466, 32'h00000000} /* (30, 18, 31) {real, imag} */,
  {32'hc55ba463, 32'h00000000} /* (30, 18, 30) {real, imag} */,
  {32'hc534851e, 32'h00000000} /* (30, 18, 29) {real, imag} */,
  {32'hc535cbee, 32'h00000000} /* (30, 18, 28) {real, imag} */,
  {32'hc54c782a, 32'h00000000} /* (30, 18, 27) {real, imag} */,
  {32'hc52f1989, 32'h00000000} /* (30, 18, 26) {real, imag} */,
  {32'hc4f9aeaa, 32'h00000000} /* (30, 18, 25) {real, imag} */,
  {32'hc4ebc664, 32'h00000000} /* (30, 18, 24) {real, imag} */,
  {32'hc4d14f7c, 32'h00000000} /* (30, 18, 23) {real, imag} */,
  {32'hc4c687e2, 32'h00000000} /* (30, 18, 22) {real, imag} */,
  {32'hc4092e5c, 32'h00000000} /* (30, 18, 21) {real, imag} */,
  {32'h4466ce3e, 32'h00000000} /* (30, 18, 20) {real, imag} */,
  {32'h451fc519, 32'h00000000} /* (30, 18, 19) {real, imag} */,
  {32'h4526dc7a, 32'h00000000} /* (30, 18, 18) {real, imag} */,
  {32'h4539b9b8, 32'h00000000} /* (30, 18, 17) {real, imag} */,
  {32'h451d6e4b, 32'h00000000} /* (30, 18, 16) {real, imag} */,
  {32'h45235ab6, 32'h00000000} /* (30, 18, 15) {real, imag} */,
  {32'h4549ed65, 32'h00000000} /* (30, 18, 14) {real, imag} */,
  {32'h45417684, 32'h00000000} /* (30, 18, 13) {real, imag} */,
  {32'h454adec6, 32'h00000000} /* (30, 18, 12) {real, imag} */,
  {32'h4529285a, 32'h00000000} /* (30, 18, 11) {real, imag} */,
  {32'hc4a6cc6a, 32'h00000000} /* (30, 18, 10) {real, imag} */,
  {32'hc5493d83, 32'h00000000} /* (30, 18, 9) {real, imag} */,
  {32'hc554b9d2, 32'h00000000} /* (30, 18, 8) {real, imag} */,
  {32'hc589875b, 32'h00000000} /* (30, 18, 7) {real, imag} */,
  {32'hc5394e93, 32'h00000000} /* (30, 18, 6) {real, imag} */,
  {32'hc53c4e39, 32'h00000000} /* (30, 18, 5) {real, imag} */,
  {32'hc553b136, 32'h00000000} /* (30, 18, 4) {real, imag} */,
  {32'hc55dd891, 32'h00000000} /* (30, 18, 3) {real, imag} */,
  {32'hc547951e, 32'h00000000} /* (30, 18, 2) {real, imag} */,
  {32'hc5459658, 32'h00000000} /* (30, 18, 1) {real, imag} */,
  {32'hc5270675, 32'h00000000} /* (30, 18, 0) {real, imag} */,
  {32'hc5659244, 32'h00000000} /* (30, 17, 31) {real, imag} */,
  {32'hc581275f, 32'h00000000} /* (30, 17, 30) {real, imag} */,
  {32'hc55405dc, 32'h00000000} /* (30, 17, 29) {real, imag} */,
  {32'hc55e3520, 32'h00000000} /* (30, 17, 28) {real, imag} */,
  {32'hc565fd2f, 32'h00000000} /* (30, 17, 27) {real, imag} */,
  {32'hc5102152, 32'h00000000} /* (30, 17, 26) {real, imag} */,
  {32'hc51cdfc6, 32'h00000000} /* (30, 17, 25) {real, imag} */,
  {32'hc51527cf, 32'h00000000} /* (30, 17, 24) {real, imag} */,
  {32'hc4e5ab98, 32'h00000000} /* (30, 17, 23) {real, imag} */,
  {32'hc4df5207, 32'h00000000} /* (30, 17, 22) {real, imag} */,
  {32'hc4812f55, 32'h00000000} /* (30, 17, 21) {real, imag} */,
  {32'h44f80be3, 32'h00000000} /* (30, 17, 20) {real, imag} */,
  {32'h45059f02, 32'h00000000} /* (30, 17, 19) {real, imag} */,
  {32'h4529ecbe, 32'h00000000} /* (30, 17, 18) {real, imag} */,
  {32'h45594c5f, 32'h00000000} /* (30, 17, 17) {real, imag} */,
  {32'h45388c64, 32'h00000000} /* (30, 17, 16) {real, imag} */,
  {32'h4533a206, 32'h00000000} /* (30, 17, 15) {real, imag} */,
  {32'h455e9d9e, 32'h00000000} /* (30, 17, 14) {real, imag} */,
  {32'h45446f86, 32'h00000000} /* (30, 17, 13) {real, imag} */,
  {32'h451d3c9e, 32'h00000000} /* (30, 17, 12) {real, imag} */,
  {32'h4521c171, 32'h00000000} /* (30, 17, 11) {real, imag} */,
  {32'hc4a2c34e, 32'h00000000} /* (30, 17, 10) {real, imag} */,
  {32'hc523b59c, 32'h00000000} /* (30, 17, 9) {real, imag} */,
  {32'hc5492937, 32'h00000000} /* (30, 17, 8) {real, imag} */,
  {32'hc5426f40, 32'h00000000} /* (30, 17, 7) {real, imag} */,
  {32'hc56297f8, 32'h00000000} /* (30, 17, 6) {real, imag} */,
  {32'hc5585b44, 32'h00000000} /* (30, 17, 5) {real, imag} */,
  {32'hc5744d96, 32'h00000000} /* (30, 17, 4) {real, imag} */,
  {32'hc5630eee, 32'h00000000} /* (30, 17, 3) {real, imag} */,
  {32'hc55966fe, 32'h00000000} /* (30, 17, 2) {real, imag} */,
  {32'hc553989d, 32'h00000000} /* (30, 17, 1) {real, imag} */,
  {32'hc542048a, 32'h00000000} /* (30, 17, 0) {real, imag} */,
  {32'hc5461d16, 32'h00000000} /* (30, 16, 31) {real, imag} */,
  {32'hc5724746, 32'h00000000} /* (30, 16, 30) {real, imag} */,
  {32'hc58670ee, 32'h00000000} /* (30, 16, 29) {real, imag} */,
  {32'hc52f714d, 32'h00000000} /* (30, 16, 28) {real, imag} */,
  {32'hc532c23c, 32'h00000000} /* (30, 16, 27) {real, imag} */,
  {32'hc5413883, 32'h00000000} /* (30, 16, 26) {real, imag} */,
  {32'hc52efc5b, 32'h00000000} /* (30, 16, 25) {real, imag} */,
  {32'hc5946792, 32'h00000000} /* (30, 16, 24) {real, imag} */,
  {32'hc520f210, 32'h00000000} /* (30, 16, 23) {real, imag} */,
  {32'hc4d57060, 32'h00000000} /* (30, 16, 22) {real, imag} */,
  {32'h423c7040, 32'h00000000} /* (30, 16, 21) {real, imag} */,
  {32'h44ffaabd, 32'h00000000} /* (30, 16, 20) {real, imag} */,
  {32'h455315ea, 32'h00000000} /* (30, 16, 19) {real, imag} */,
  {32'h453290cd, 32'h00000000} /* (30, 16, 18) {real, imag} */,
  {32'h45498e4a, 32'h00000000} /* (30, 16, 17) {real, imag} */,
  {32'h454b70a7, 32'h00000000} /* (30, 16, 16) {real, imag} */,
  {32'h4562c84c, 32'h00000000} /* (30, 16, 15) {real, imag} */,
  {32'h453d6b8c, 32'h00000000} /* (30, 16, 14) {real, imag} */,
  {32'h452bec0e, 32'h00000000} /* (30, 16, 13) {real, imag} */,
  {32'h4527dbb7, 32'h00000000} /* (30, 16, 12) {real, imag} */,
  {32'h4439d51a, 32'h00000000} /* (30, 16, 11) {real, imag} */,
  {32'hc5079ce9, 32'h00000000} /* (30, 16, 10) {real, imag} */,
  {32'hc524158d, 32'h00000000} /* (30, 16, 9) {real, imag} */,
  {32'hc51333c7, 32'h00000000} /* (30, 16, 8) {real, imag} */,
  {32'hc54cd3d6, 32'h00000000} /* (30, 16, 7) {real, imag} */,
  {32'hc582352d, 32'h00000000} /* (30, 16, 6) {real, imag} */,
  {32'hc5815126, 32'h00000000} /* (30, 16, 5) {real, imag} */,
  {32'hc57ca65c, 32'h00000000} /* (30, 16, 4) {real, imag} */,
  {32'hc5793fda, 32'h00000000} /* (30, 16, 3) {real, imag} */,
  {32'hc576b655, 32'h00000000} /* (30, 16, 2) {real, imag} */,
  {32'hc55b2592, 32'h00000000} /* (30, 16, 1) {real, imag} */,
  {32'hc52db77f, 32'h00000000} /* (30, 16, 0) {real, imag} */,
  {32'hc52f048a, 32'h00000000} /* (30, 15, 31) {real, imag} */,
  {32'hc5605750, 32'h00000000} /* (30, 15, 30) {real, imag} */,
  {32'hc56ed273, 32'h00000000} /* (30, 15, 29) {real, imag} */,
  {32'hc56665ce, 32'h00000000} /* (30, 15, 28) {real, imag} */,
  {32'hc5402d28, 32'h00000000} /* (30, 15, 27) {real, imag} */,
  {32'hc5191c13, 32'h00000000} /* (30, 15, 26) {real, imag} */,
  {32'hc5474a7a, 32'h00000000} /* (30, 15, 25) {real, imag} */,
  {32'hc52dcde9, 32'h00000000} /* (30, 15, 24) {real, imag} */,
  {32'hc5056d49, 32'h00000000} /* (30, 15, 23) {real, imag} */,
  {32'hc4ea0127, 32'h00000000} /* (30, 15, 22) {real, imag} */,
  {32'hc38fe200, 32'h00000000} /* (30, 15, 21) {real, imag} */,
  {32'h441bb108, 32'h00000000} /* (30, 15, 20) {real, imag} */,
  {32'h452c7924, 32'h00000000} /* (30, 15, 19) {real, imag} */,
  {32'h453a14e6, 32'h00000000} /* (30, 15, 18) {real, imag} */,
  {32'h452b27b5, 32'h00000000} /* (30, 15, 17) {real, imag} */,
  {32'h454d7718, 32'h00000000} /* (30, 15, 16) {real, imag} */,
  {32'h455e0fa2, 32'h00000000} /* (30, 15, 15) {real, imag} */,
  {32'h45503c80, 32'h00000000} /* (30, 15, 14) {real, imag} */,
  {32'h452165df, 32'h00000000} /* (30, 15, 13) {real, imag} */,
  {32'h44c141d4, 32'h00000000} /* (30, 15, 12) {real, imag} */,
  {32'h43871e84, 32'h00000000} /* (30, 15, 11) {real, imag} */,
  {32'hc4e594e2, 32'h00000000} /* (30, 15, 10) {real, imag} */,
  {32'hc5398ca4, 32'h00000000} /* (30, 15, 9) {real, imag} */,
  {32'hc569fe2f, 32'h00000000} /* (30, 15, 8) {real, imag} */,
  {32'hc5634ceb, 32'h00000000} /* (30, 15, 7) {real, imag} */,
  {32'hc56789d4, 32'h00000000} /* (30, 15, 6) {real, imag} */,
  {32'hc59551a5, 32'h00000000} /* (30, 15, 5) {real, imag} */,
  {32'hc571042e, 32'h00000000} /* (30, 15, 4) {real, imag} */,
  {32'hc56d43cc, 32'h00000000} /* (30, 15, 3) {real, imag} */,
  {32'hc54c138e, 32'h00000000} /* (30, 15, 2) {real, imag} */,
  {32'hc5500abd, 32'h00000000} /* (30, 15, 1) {real, imag} */,
  {32'hc51ef5ec, 32'h00000000} /* (30, 15, 0) {real, imag} */,
  {32'hc5301ce9, 32'h00000000} /* (30, 14, 31) {real, imag} */,
  {32'hc5701c16, 32'h00000000} /* (30, 14, 30) {real, imag} */,
  {32'hc558986e, 32'h00000000} /* (30, 14, 29) {real, imag} */,
  {32'hc54b0212, 32'h00000000} /* (30, 14, 28) {real, imag} */,
  {32'hc520b631, 32'h00000000} /* (30, 14, 27) {real, imag} */,
  {32'hc5222886, 32'h00000000} /* (30, 14, 26) {real, imag} */,
  {32'hc553949a, 32'h00000000} /* (30, 14, 25) {real, imag} */,
  {32'hc53b03e0, 32'h00000000} /* (30, 14, 24) {real, imag} */,
  {32'hc516d9d0, 32'h00000000} /* (30, 14, 23) {real, imag} */,
  {32'hc5006514, 32'h00000000} /* (30, 14, 22) {real, imag} */,
  {32'hc4398a26, 32'h00000000} /* (30, 14, 21) {real, imag} */,
  {32'h44c277c4, 32'h00000000} /* (30, 14, 20) {real, imag} */,
  {32'h44b51b6e, 32'h00000000} /* (30, 14, 19) {real, imag} */,
  {32'h4528f367, 32'h00000000} /* (30, 14, 18) {real, imag} */,
  {32'h4502e96b, 32'h00000000} /* (30, 14, 17) {real, imag} */,
  {32'h4552620f, 32'h00000000} /* (30, 14, 16) {real, imag} */,
  {32'h455c2a0d, 32'h00000000} /* (30, 14, 15) {real, imag} */,
  {32'h452c28fa, 32'h00000000} /* (30, 14, 14) {real, imag} */,
  {32'h4516b5b4, 32'h00000000} /* (30, 14, 13) {real, imag} */,
  {32'h449fe780, 32'h00000000} /* (30, 14, 12) {real, imag} */,
  {32'h4455d08b, 32'h00000000} /* (30, 14, 11) {real, imag} */,
  {32'hc4a102dc, 32'h00000000} /* (30, 14, 10) {real, imag} */,
  {32'hc5461538, 32'h00000000} /* (30, 14, 9) {real, imag} */,
  {32'hc56dd7a6, 32'h00000000} /* (30, 14, 8) {real, imag} */,
  {32'hc55d4ea6, 32'h00000000} /* (30, 14, 7) {real, imag} */,
  {32'hc54eda7c, 32'h00000000} /* (30, 14, 6) {real, imag} */,
  {32'hc585071c, 32'h00000000} /* (30, 14, 5) {real, imag} */,
  {32'hc5594286, 32'h00000000} /* (30, 14, 4) {real, imag} */,
  {32'hc54ed697, 32'h00000000} /* (30, 14, 3) {real, imag} */,
  {32'hc5395a8b, 32'h00000000} /* (30, 14, 2) {real, imag} */,
  {32'hc4ff66ba, 32'h00000000} /* (30, 14, 1) {real, imag} */,
  {32'hc51346bf, 32'h00000000} /* (30, 14, 0) {real, imag} */,
  {32'hc5222940, 32'h00000000} /* (30, 13, 31) {real, imag} */,
  {32'hc54339b4, 32'h00000000} /* (30, 13, 30) {real, imag} */,
  {32'hc52badc9, 32'h00000000} /* (30, 13, 29) {real, imag} */,
  {32'hc537fd90, 32'h00000000} /* (30, 13, 28) {real, imag} */,
  {32'hc55626a4, 32'h00000000} /* (30, 13, 27) {real, imag} */,
  {32'hc533329a, 32'h00000000} /* (30, 13, 26) {real, imag} */,
  {32'hc535600c, 32'h00000000} /* (30, 13, 25) {real, imag} */,
  {32'hc57f3b46, 32'h00000000} /* (30, 13, 24) {real, imag} */,
  {32'hc55d5711, 32'h00000000} /* (30, 13, 23) {real, imag} */,
  {32'hc4ebf5f6, 32'h00000000} /* (30, 13, 22) {real, imag} */,
  {32'hc4a80ef9, 32'h00000000} /* (30, 13, 21) {real, imag} */,
  {32'h44a459d6, 32'h00000000} /* (30, 13, 20) {real, imag} */,
  {32'h44ecfbd9, 32'h00000000} /* (30, 13, 19) {real, imag} */,
  {32'h44c93394, 32'h00000000} /* (30, 13, 18) {real, imag} */,
  {32'h452cd1ea, 32'h00000000} /* (30, 13, 17) {real, imag} */,
  {32'h4530a433, 32'h00000000} /* (30, 13, 16) {real, imag} */,
  {32'h454ab808, 32'h00000000} /* (30, 13, 15) {real, imag} */,
  {32'h45188b5e, 32'h00000000} /* (30, 13, 14) {real, imag} */,
  {32'h44b0f04a, 32'h00000000} /* (30, 13, 13) {real, imag} */,
  {32'h449996d0, 32'h00000000} /* (30, 13, 12) {real, imag} */,
  {32'h444215da, 32'h00000000} /* (30, 13, 11) {real, imag} */,
  {32'hc4858ae4, 32'h00000000} /* (30, 13, 10) {real, imag} */,
  {32'hc5268088, 32'h00000000} /* (30, 13, 9) {real, imag} */,
  {32'hc55e5f60, 32'h00000000} /* (30, 13, 8) {real, imag} */,
  {32'hc5612755, 32'h00000000} /* (30, 13, 7) {real, imag} */,
  {32'hc56786b9, 32'h00000000} /* (30, 13, 6) {real, imag} */,
  {32'hc588bcd9, 32'h00000000} /* (30, 13, 5) {real, imag} */,
  {32'hc57a6167, 32'h00000000} /* (30, 13, 4) {real, imag} */,
  {32'hc56cb5ea, 32'h00000000} /* (30, 13, 3) {real, imag} */,
  {32'hc500ee82, 32'h00000000} /* (30, 13, 2) {real, imag} */,
  {32'hc51fc96c, 32'h00000000} /* (30, 13, 1) {real, imag} */,
  {32'hc51974b9, 32'h00000000} /* (30, 13, 0) {real, imag} */,
  {32'hc4f0e996, 32'h00000000} /* (30, 12, 31) {real, imag} */,
  {32'hc4ed20f2, 32'h00000000} /* (30, 12, 30) {real, imag} */,
  {32'hc50036bb, 32'h00000000} /* (30, 12, 29) {real, imag} */,
  {32'hc50084d9, 32'h00000000} /* (30, 12, 28) {real, imag} */,
  {32'hc548029e, 32'h00000000} /* (30, 12, 27) {real, imag} */,
  {32'hc5278546, 32'h00000000} /* (30, 12, 26) {real, imag} */,
  {32'hc52e52ad, 32'h00000000} /* (30, 12, 25) {real, imag} */,
  {32'hc52010b8, 32'h00000000} /* (30, 12, 24) {real, imag} */,
  {32'hc51131ff, 32'h00000000} /* (30, 12, 23) {real, imag} */,
  {32'hc521bdbc, 32'h00000000} /* (30, 12, 22) {real, imag} */,
  {32'hc4b1d233, 32'h00000000} /* (30, 12, 21) {real, imag} */,
  {32'h4394e0f4, 32'h00000000} /* (30, 12, 20) {real, imag} */,
  {32'h44ee0686, 32'h00000000} /* (30, 12, 19) {real, imag} */,
  {32'h450bdea5, 32'h00000000} /* (30, 12, 18) {real, imag} */,
  {32'h450d199b, 32'h00000000} /* (30, 12, 17) {real, imag} */,
  {32'h450f7d1b, 32'h00000000} /* (30, 12, 16) {real, imag} */,
  {32'h4506122b, 32'h00000000} /* (30, 12, 15) {real, imag} */,
  {32'h44d59e42, 32'h00000000} /* (30, 12, 14) {real, imag} */,
  {32'h44dc2f2c, 32'h00000000} /* (30, 12, 13) {real, imag} */,
  {32'h449e28ac, 32'h00000000} /* (30, 12, 12) {real, imag} */,
  {32'h4379dd38, 32'h00000000} /* (30, 12, 11) {real, imag} */,
  {32'hc47d3690, 32'h00000000} /* (30, 12, 10) {real, imag} */,
  {32'hc4f3251e, 32'h00000000} /* (30, 12, 9) {real, imag} */,
  {32'hc519463e, 32'h00000000} /* (30, 12, 8) {real, imag} */,
  {32'hc5301229, 32'h00000000} /* (30, 12, 7) {real, imag} */,
  {32'hc535b20a, 32'h00000000} /* (30, 12, 6) {real, imag} */,
  {32'hc52b4a96, 32'h00000000} /* (30, 12, 5) {real, imag} */,
  {32'hc5522db8, 32'h00000000} /* (30, 12, 4) {real, imag} */,
  {32'hc54efca5, 32'h00000000} /* (30, 12, 3) {real, imag} */,
  {32'hc51f6ea9, 32'h00000000} /* (30, 12, 2) {real, imag} */,
  {32'hc502e397, 32'h00000000} /* (30, 12, 1) {real, imag} */,
  {32'hc518b3ad, 32'h00000000} /* (30, 12, 0) {real, imag} */,
  {32'hc44fc1c6, 32'h00000000} /* (30, 11, 31) {real, imag} */,
  {32'hc44b63f1, 32'h00000000} /* (30, 11, 30) {real, imag} */,
  {32'hc4c548f9, 32'h00000000} /* (30, 11, 29) {real, imag} */,
  {32'hc4eb6fe7, 32'h00000000} /* (30, 11, 28) {real, imag} */,
  {32'hc4a23260, 32'h00000000} /* (30, 11, 27) {real, imag} */,
  {32'hc487bfa0, 32'h00000000} /* (30, 11, 26) {real, imag} */,
  {32'hc52a54cb, 32'h00000000} /* (30, 11, 25) {real, imag} */,
  {32'hc4974028, 32'h00000000} /* (30, 11, 24) {real, imag} */,
  {32'hc478848e, 32'h00000000} /* (30, 11, 23) {real, imag} */,
  {32'hc50f0802, 32'h00000000} /* (30, 11, 22) {real, imag} */,
  {32'hc4367cf3, 32'h00000000} /* (30, 11, 21) {real, imag} */,
  {32'h44006e28, 32'h00000000} /* (30, 11, 20) {real, imag} */,
  {32'h44b9b0fa, 32'h00000000} /* (30, 11, 19) {real, imag} */,
  {32'h445220de, 32'h00000000} /* (30, 11, 18) {real, imag} */,
  {32'h44e928fb, 32'h00000000} /* (30, 11, 17) {real, imag} */,
  {32'h45198ba4, 32'h00000000} /* (30, 11, 16) {real, imag} */,
  {32'h449494c3, 32'h00000000} /* (30, 11, 15) {real, imag} */,
  {32'h44d86278, 32'h00000000} /* (30, 11, 14) {real, imag} */,
  {32'h446d13fe, 32'h00000000} /* (30, 11, 13) {real, imag} */,
  {32'hc13cb780, 32'h00000000} /* (30, 11, 12) {real, imag} */,
  {32'h43e1be9a, 32'h00000000} /* (30, 11, 11) {real, imag} */,
  {32'hc4285478, 32'h00000000} /* (30, 11, 10) {real, imag} */,
  {32'hc51873df, 32'h00000000} /* (30, 11, 9) {real, imag} */,
  {32'hc4d0be9c, 32'h00000000} /* (30, 11, 8) {real, imag} */,
  {32'hc4394c2a, 32'h00000000} /* (30, 11, 7) {real, imag} */,
  {32'hc4a10b7b, 32'h00000000} /* (30, 11, 6) {real, imag} */,
  {32'hc4a94804, 32'h00000000} /* (30, 11, 5) {real, imag} */,
  {32'hc4707288, 32'h00000000} /* (30, 11, 4) {real, imag} */,
  {32'hc515075b, 32'h00000000} /* (30, 11, 3) {real, imag} */,
  {32'hc49a3771, 32'h00000000} /* (30, 11, 2) {real, imag} */,
  {32'hc4913197, 32'h00000000} /* (30, 11, 1) {real, imag} */,
  {32'hc495cbc4, 32'h00000000} /* (30, 11, 0) {real, imag} */,
  {32'h449050dc, 32'h00000000} /* (30, 10, 31) {real, imag} */,
  {32'h448394b6, 32'h00000000} /* (30, 10, 30) {real, imag} */,
  {32'h43063fe8, 32'h00000000} /* (30, 10, 29) {real, imag} */,
  {32'hc1975260, 32'h00000000} /* (30, 10, 28) {real, imag} */,
  {32'h43dd5fe3, 32'h00000000} /* (30, 10, 27) {real, imag} */,
  {32'h44144b8e, 32'h00000000} /* (30, 10, 26) {real, imag} */,
  {32'h4452b831, 32'h00000000} /* (30, 10, 25) {real, imag} */,
  {32'h434fd5cc, 32'h00000000} /* (30, 10, 24) {real, imag} */,
  {32'h442a3886, 32'h00000000} /* (30, 10, 23) {real, imag} */,
  {32'h43d2dbb2, 32'h00000000} /* (30, 10, 22) {real, imag} */,
  {32'hc43ab479, 32'h00000000} /* (30, 10, 21) {real, imag} */,
  {32'hc3be4102, 32'h00000000} /* (30, 10, 20) {real, imag} */,
  {32'hc3c68ee0, 32'h00000000} /* (30, 10, 19) {real, imag} */,
  {32'hc3acc98f, 32'h00000000} /* (30, 10, 18) {real, imag} */,
  {32'hc32e6092, 32'h00000000} /* (30, 10, 17) {real, imag} */,
  {32'hc429137c, 32'h00000000} /* (30, 10, 16) {real, imag} */,
  {32'hc48576d2, 32'h00000000} /* (30, 10, 15) {real, imag} */,
  {32'hc48db554, 32'h00000000} /* (30, 10, 14) {real, imag} */,
  {32'hc4da2797, 32'h00000000} /* (30, 10, 13) {real, imag} */,
  {32'hc4a70294, 32'h00000000} /* (30, 10, 12) {real, imag} */,
  {32'hc36c12ea, 32'h00000000} /* (30, 10, 11) {real, imag} */,
  {32'hc325b55a, 32'h00000000} /* (30, 10, 10) {real, imag} */,
  {32'hc31a63dc, 32'h00000000} /* (30, 10, 9) {real, imag} */,
  {32'h44409087, 32'h00000000} /* (30, 10, 8) {real, imag} */,
  {32'h44b775d3, 32'h00000000} /* (30, 10, 7) {real, imag} */,
  {32'h44ea1210, 32'h00000000} /* (30, 10, 6) {real, imag} */,
  {32'h4432bc85, 32'h00000000} /* (30, 10, 5) {real, imag} */,
  {32'h44da8f3e, 32'h00000000} /* (30, 10, 4) {real, imag} */,
  {32'h444cd738, 32'h00000000} /* (30, 10, 3) {real, imag} */,
  {32'h442eae7a, 32'h00000000} /* (30, 10, 2) {real, imag} */,
  {32'h442fbcda, 32'h00000000} /* (30, 10, 1) {real, imag} */,
  {32'h440e05b4, 32'h00000000} /* (30, 10, 0) {real, imag} */,
  {32'h44ba1168, 32'h00000000} /* (30, 9, 31) {real, imag} */,
  {32'h451cf285, 32'h00000000} /* (30, 9, 30) {real, imag} */,
  {32'h44cad46a, 32'h00000000} /* (30, 9, 29) {real, imag} */,
  {32'h44e7597b, 32'h00000000} /* (30, 9, 28) {real, imag} */,
  {32'h44e9798b, 32'h00000000} /* (30, 9, 27) {real, imag} */,
  {32'h44d5c43e, 32'h00000000} /* (30, 9, 26) {real, imag} */,
  {32'h4501ef44, 32'h00000000} /* (30, 9, 25) {real, imag} */,
  {32'h44cb3133, 32'h00000000} /* (30, 9, 24) {real, imag} */,
  {32'h4493c55f, 32'h00000000} /* (30, 9, 23) {real, imag} */,
  {32'h4447dc68, 32'h00000000} /* (30, 9, 22) {real, imag} */,
  {32'h44105c92, 32'h00000000} /* (30, 9, 21) {real, imag} */,
  {32'hc454eda8, 32'h00000000} /* (30, 9, 20) {real, imag} */,
  {32'hc4bcd35b, 32'h00000000} /* (30, 9, 19) {real, imag} */,
  {32'hc4a48c62, 32'h00000000} /* (30, 9, 18) {real, imag} */,
  {32'hc5073562, 32'h00000000} /* (30, 9, 17) {real, imag} */,
  {32'hc548a285, 32'h00000000} /* (30, 9, 16) {real, imag} */,
  {32'hc512a9f7, 32'h00000000} /* (30, 9, 15) {real, imag} */,
  {32'hc52d6385, 32'h00000000} /* (30, 9, 14) {real, imag} */,
  {32'hc509868f, 32'h00000000} /* (30, 9, 13) {real, imag} */,
  {32'hc4f4435d, 32'h00000000} /* (30, 9, 12) {real, imag} */,
  {32'hc4d30853, 32'h00000000} /* (30, 9, 11) {real, imag} */,
  {32'hc38a64b0, 32'h00000000} /* (30, 9, 10) {real, imag} */,
  {32'h4440b094, 32'h00000000} /* (30, 9, 9) {real, imag} */,
  {32'h4490078d, 32'h00000000} /* (30, 9, 8) {real, imag} */,
  {32'h44fca9f9, 32'h00000000} /* (30, 9, 7) {real, imag} */,
  {32'h44be6bb4, 32'h00000000} /* (30, 9, 6) {real, imag} */,
  {32'h454b234c, 32'h00000000} /* (30, 9, 5) {real, imag} */,
  {32'h450382f2, 32'h00000000} /* (30, 9, 4) {real, imag} */,
  {32'h45232346, 32'h00000000} /* (30, 9, 3) {real, imag} */,
  {32'h4515c69b, 32'h00000000} /* (30, 9, 2) {real, imag} */,
  {32'h452193c2, 32'h00000000} /* (30, 9, 1) {real, imag} */,
  {32'h44ebc8c2, 32'h00000000} /* (30, 9, 0) {real, imag} */,
  {32'h44f3fa77, 32'h00000000} /* (30, 8, 31) {real, imag} */,
  {32'h451f973e, 32'h00000000} /* (30, 8, 30) {real, imag} */,
  {32'h4525d573, 32'h00000000} /* (30, 8, 29) {real, imag} */,
  {32'h44f485f8, 32'h00000000} /* (30, 8, 28) {real, imag} */,
  {32'h4510ba28, 32'h00000000} /* (30, 8, 27) {real, imag} */,
  {32'h45313fbe, 32'h00000000} /* (30, 8, 26) {real, imag} */,
  {32'h45081c16, 32'h00000000} /* (30, 8, 25) {real, imag} */,
  {32'h4503502a, 32'h00000000} /* (30, 8, 24) {real, imag} */,
  {32'h44cb70aa, 32'h00000000} /* (30, 8, 23) {real, imag} */,
  {32'h44a23ffb, 32'h00000000} /* (30, 8, 22) {real, imag} */,
  {32'h44201bc1, 32'h00000000} /* (30, 8, 21) {real, imag} */,
  {32'hc4c10893, 32'h00000000} /* (30, 8, 20) {real, imag} */,
  {32'hc4e7cde1, 32'h00000000} /* (30, 8, 19) {real, imag} */,
  {32'hc5136cbf, 32'h00000000} /* (30, 8, 18) {real, imag} */,
  {32'hc53173de, 32'h00000000} /* (30, 8, 17) {real, imag} */,
  {32'hc53c641d, 32'h00000000} /* (30, 8, 16) {real, imag} */,
  {32'hc53e0fd0, 32'h00000000} /* (30, 8, 15) {real, imag} */,
  {32'hc58e1aeb, 32'h00000000} /* (30, 8, 14) {real, imag} */,
  {32'hc546ce71, 32'h00000000} /* (30, 8, 13) {real, imag} */,
  {32'hc58df0ec, 32'h00000000} /* (30, 8, 12) {real, imag} */,
  {32'hc515189a, 32'h00000000} /* (30, 8, 11) {real, imag} */,
  {32'hc413f59a, 32'h00000000} /* (30, 8, 10) {real, imag} */,
  {32'h44438843, 32'h00000000} /* (30, 8, 9) {real, imag} */,
  {32'h444e3f62, 32'h00000000} /* (30, 8, 8) {real, imag} */,
  {32'h44e9772c, 32'h00000000} /* (30, 8, 7) {real, imag} */,
  {32'h4518a548, 32'h00000000} /* (30, 8, 6) {real, imag} */,
  {32'h450c4ec2, 32'h00000000} /* (30, 8, 5) {real, imag} */,
  {32'h452b2f64, 32'h00000000} /* (30, 8, 4) {real, imag} */,
  {32'h45678a38, 32'h00000000} /* (30, 8, 3) {real, imag} */,
  {32'h4532e5f3, 32'h00000000} /* (30, 8, 2) {real, imag} */,
  {32'h45277200, 32'h00000000} /* (30, 8, 1) {real, imag} */,
  {32'h45108c6b, 32'h00000000} /* (30, 8, 0) {real, imag} */,
  {32'h45294bb8, 32'h00000000} /* (30, 7, 31) {real, imag} */,
  {32'h44f7cab2, 32'h00000000} /* (30, 7, 30) {real, imag} */,
  {32'h44faf2f5, 32'h00000000} /* (30, 7, 29) {real, imag} */,
  {32'h4532c572, 32'h00000000} /* (30, 7, 28) {real, imag} */,
  {32'h45001464, 32'h00000000} /* (30, 7, 27) {real, imag} */,
  {32'h4507158c, 32'h00000000} /* (30, 7, 26) {real, imag} */,
  {32'h4524ec6f, 32'h00000000} /* (30, 7, 25) {real, imag} */,
  {32'h450def5c, 32'h00000000} /* (30, 7, 24) {real, imag} */,
  {32'h45079682, 32'h00000000} /* (30, 7, 23) {real, imag} */,
  {32'h44f7d856, 32'h00000000} /* (30, 7, 22) {real, imag} */,
  {32'h42c7cbb0, 32'h00000000} /* (30, 7, 21) {real, imag} */,
  {32'hc4a514b6, 32'h00000000} /* (30, 7, 20) {real, imag} */,
  {32'hc4b59cdb, 32'h00000000} /* (30, 7, 19) {real, imag} */,
  {32'hc500601b, 32'h00000000} /* (30, 7, 18) {real, imag} */,
  {32'hc511e829, 32'h00000000} /* (30, 7, 17) {real, imag} */,
  {32'hc52a9a7c, 32'h00000000} /* (30, 7, 16) {real, imag} */,
  {32'hc52af4e8, 32'h00000000} /* (30, 7, 15) {real, imag} */,
  {32'hc5484959, 32'h00000000} /* (30, 7, 14) {real, imag} */,
  {32'hc5456d9c, 32'h00000000} /* (30, 7, 13) {real, imag} */,
  {32'hc5553718, 32'h00000000} /* (30, 7, 12) {real, imag} */,
  {32'hc5415f6e, 32'h00000000} /* (30, 7, 11) {real, imag} */,
  {32'hc3752e08, 32'h00000000} /* (30, 7, 10) {real, imag} */,
  {32'h444d6174, 32'h00000000} /* (30, 7, 9) {real, imag} */,
  {32'h44bef6ac, 32'h00000000} /* (30, 7, 8) {real, imag} */,
  {32'h45166736, 32'h00000000} /* (30, 7, 7) {real, imag} */,
  {32'h452e2d9d, 32'h00000000} /* (30, 7, 6) {real, imag} */,
  {32'h4560aed6, 32'h00000000} /* (30, 7, 5) {real, imag} */,
  {32'h4555931b, 32'h00000000} /* (30, 7, 4) {real, imag} */,
  {32'h457192da, 32'h00000000} /* (30, 7, 3) {real, imag} */,
  {32'h4578f94f, 32'h00000000} /* (30, 7, 2) {real, imag} */,
  {32'h45402bcb, 32'h00000000} /* (30, 7, 1) {real, imag} */,
  {32'h4512469c, 32'h00000000} /* (30, 7, 0) {real, imag} */,
  {32'h4500c00c, 32'h00000000} /* (30, 6, 31) {real, imag} */,
  {32'h4512c990, 32'h00000000} /* (30, 6, 30) {real, imag} */,
  {32'h45343e8c, 32'h00000000} /* (30, 6, 29) {real, imag} */,
  {32'h44f222be, 32'h00000000} /* (30, 6, 28) {real, imag} */,
  {32'h44e0953f, 32'h00000000} /* (30, 6, 27) {real, imag} */,
  {32'h44a80ffa, 32'h00000000} /* (30, 6, 26) {real, imag} */,
  {32'h4524b57e, 32'h00000000} /* (30, 6, 25) {real, imag} */,
  {32'h45414b7e, 32'h00000000} /* (30, 6, 24) {real, imag} */,
  {32'h451dbb65, 32'h00000000} /* (30, 6, 23) {real, imag} */,
  {32'h45037120, 32'h00000000} /* (30, 6, 22) {real, imag} */,
  {32'h44bea7a6, 32'h00000000} /* (30, 6, 21) {real, imag} */,
  {32'hc3ecc3a6, 32'h00000000} /* (30, 6, 20) {real, imag} */,
  {32'hc465bcd6, 32'h00000000} /* (30, 6, 19) {real, imag} */,
  {32'hc498fdca, 32'h00000000} /* (30, 6, 18) {real, imag} */,
  {32'hc5273ddc, 32'h00000000} /* (30, 6, 17) {real, imag} */,
  {32'hc51ec360, 32'h00000000} /* (30, 6, 16) {real, imag} */,
  {32'hc52235c2, 32'h00000000} /* (30, 6, 15) {real, imag} */,
  {32'hc57712a0, 32'h00000000} /* (30, 6, 14) {real, imag} */,
  {32'hc51a6224, 32'h00000000} /* (30, 6, 13) {real, imag} */,
  {32'hc5301483, 32'h00000000} /* (30, 6, 12) {real, imag} */,
  {32'hc55225cc, 32'h00000000} /* (30, 6, 11) {real, imag} */,
  {32'hc487f444, 32'h00000000} /* (30, 6, 10) {real, imag} */,
  {32'h449abcdd, 32'h00000000} /* (30, 6, 9) {real, imag} */,
  {32'h4453d0aa, 32'h00000000} /* (30, 6, 8) {real, imag} */,
  {32'h450ce793, 32'h00000000} /* (30, 6, 7) {real, imag} */,
  {32'h451b540c, 32'h00000000} /* (30, 6, 6) {real, imag} */,
  {32'h451fa97c, 32'h00000000} /* (30, 6, 5) {real, imag} */,
  {32'h45117465, 32'h00000000} /* (30, 6, 4) {real, imag} */,
  {32'h453d5130, 32'h00000000} /* (30, 6, 3) {real, imag} */,
  {32'h45650565, 32'h00000000} /* (30, 6, 2) {real, imag} */,
  {32'h452f8230, 32'h00000000} /* (30, 6, 1) {real, imag} */,
  {32'h450af82c, 32'h00000000} /* (30, 6, 0) {real, imag} */,
  {32'h44f06d7f, 32'h00000000} /* (30, 5, 31) {real, imag} */,
  {32'h450f4b75, 32'h00000000} /* (30, 5, 30) {real, imag} */,
  {32'h4528be3a, 32'h00000000} /* (30, 5, 29) {real, imag} */,
  {32'h453c61e0, 32'h00000000} /* (30, 5, 28) {real, imag} */,
  {32'h44c30c08, 32'h00000000} /* (30, 5, 27) {real, imag} */,
  {32'h4516e106, 32'h00000000} /* (30, 5, 26) {real, imag} */,
  {32'h4500765f, 32'h00000000} /* (30, 5, 25) {real, imag} */,
  {32'h45358efa, 32'h00000000} /* (30, 5, 24) {real, imag} */,
  {32'h451ba4f2, 32'h00000000} /* (30, 5, 23) {real, imag} */,
  {32'h450dd16b, 32'h00000000} /* (30, 5, 22) {real, imag} */,
  {32'h4505398a, 32'h00000000} /* (30, 5, 21) {real, imag} */,
  {32'h44ec4056, 32'h00000000} /* (30, 5, 20) {real, imag} */,
  {32'h4449bfd2, 32'h00000000} /* (30, 5, 19) {real, imag} */,
  {32'hc1092c80, 32'h00000000} /* (30, 5, 18) {real, imag} */,
  {32'hc463b9e8, 32'h00000000} /* (30, 5, 17) {real, imag} */,
  {32'hc48ea9e8, 32'h00000000} /* (30, 5, 16) {real, imag} */,
  {32'hc52f1080, 32'h00000000} /* (30, 5, 15) {real, imag} */,
  {32'hc540aa47, 32'h00000000} /* (30, 5, 14) {real, imag} */,
  {32'hc5404c2c, 32'h00000000} /* (30, 5, 13) {real, imag} */,
  {32'hc5590596, 32'h00000000} /* (30, 5, 12) {real, imag} */,
  {32'hc5497120, 32'h00000000} /* (30, 5, 11) {real, imag} */,
  {32'hc50b65c6, 32'h00000000} /* (30, 5, 10) {real, imag} */,
  {32'hc47301a4, 32'h00000000} /* (30, 5, 9) {real, imag} */,
  {32'hc4224888, 32'h00000000} /* (30, 5, 8) {real, imag} */,
  {32'hc3594f70, 32'h00000000} /* (30, 5, 7) {real, imag} */,
  {32'h443230d5, 32'h00000000} /* (30, 5, 6) {real, imag} */,
  {32'h4507fd5a, 32'h00000000} /* (30, 5, 5) {real, imag} */,
  {32'h453483f1, 32'h00000000} /* (30, 5, 4) {real, imag} */,
  {32'h4528cae0, 32'h00000000} /* (30, 5, 3) {real, imag} */,
  {32'h4548eae6, 32'h00000000} /* (30, 5, 2) {real, imag} */,
  {32'h4527ca08, 32'h00000000} /* (30, 5, 1) {real, imag} */,
  {32'h45048736, 32'h00000000} /* (30, 5, 0) {real, imag} */,
  {32'h44a706fe, 32'h00000000} /* (30, 4, 31) {real, imag} */,
  {32'h44cffc16, 32'h00000000} /* (30, 4, 30) {real, imag} */,
  {32'h44e1dd14, 32'h00000000} /* (30, 4, 29) {real, imag} */,
  {32'h45385b88, 32'h00000000} /* (30, 4, 28) {real, imag} */,
  {32'h451ac82d, 32'h00000000} /* (30, 4, 27) {real, imag} */,
  {32'h4513fa56, 32'h00000000} /* (30, 4, 26) {real, imag} */,
  {32'h450dc88f, 32'h00000000} /* (30, 4, 25) {real, imag} */,
  {32'h450581ff, 32'h00000000} /* (30, 4, 24) {real, imag} */,
  {32'h45173b72, 32'h00000000} /* (30, 4, 23) {real, imag} */,
  {32'h4520c906, 32'h00000000} /* (30, 4, 22) {real, imag} */,
  {32'h45296e48, 32'h00000000} /* (30, 4, 21) {real, imag} */,
  {32'h451fbb32, 32'h00000000} /* (30, 4, 20) {real, imag} */,
  {32'h4502420c, 32'h00000000} /* (30, 4, 19) {real, imag} */,
  {32'h4492b763, 32'h00000000} /* (30, 4, 18) {real, imag} */,
  {32'h43d2cd5c, 32'h00000000} /* (30, 4, 17) {real, imag} */,
  {32'hc2934e68, 32'h00000000} /* (30, 4, 16) {real, imag} */,
  {32'hc5116540, 32'h00000000} /* (30, 4, 15) {real, imag} */,
  {32'hc512f10f, 32'h00000000} /* (30, 4, 14) {real, imag} */,
  {32'hc542dedc, 32'h00000000} /* (30, 4, 13) {real, imag} */,
  {32'hc54cea68, 32'h00000000} /* (30, 4, 12) {real, imag} */,
  {32'hc56ce625, 32'h00000000} /* (30, 4, 11) {real, imag} */,
  {32'hc57360b2, 32'h00000000} /* (30, 4, 10) {real, imag} */,
  {32'hc532b219, 32'h00000000} /* (30, 4, 9) {real, imag} */,
  {32'hc4dfa6b0, 32'h00000000} /* (30, 4, 8) {real, imag} */,
  {32'hc42779d2, 32'h00000000} /* (30, 4, 7) {real, imag} */,
  {32'h426edc60, 32'h00000000} /* (30, 4, 6) {real, imag} */,
  {32'h44e1b7e4, 32'h00000000} /* (30, 4, 5) {real, imag} */,
  {32'h44f45494, 32'h00000000} /* (30, 4, 4) {real, imag} */,
  {32'h45431abc, 32'h00000000} /* (30, 4, 3) {real, imag} */,
  {32'h44f1f0a1, 32'h00000000} /* (30, 4, 2) {real, imag} */,
  {32'h44ff3ba9, 32'h00000000} /* (30, 4, 1) {real, imag} */,
  {32'h44e37a92, 32'h00000000} /* (30, 4, 0) {real, imag} */,
  {32'h44cd6d7a, 32'h00000000} /* (30, 3, 31) {real, imag} */,
  {32'h4501e645, 32'h00000000} /* (30, 3, 30) {real, imag} */,
  {32'h451fb243, 32'h00000000} /* (30, 3, 29) {real, imag} */,
  {32'h44c5a948, 32'h00000000} /* (30, 3, 28) {real, imag} */,
  {32'h4527b858, 32'h00000000} /* (30, 3, 27) {real, imag} */,
  {32'h45457120, 32'h00000000} /* (30, 3, 26) {real, imag} */,
  {32'h452c905c, 32'h00000000} /* (30, 3, 25) {real, imag} */,
  {32'h4516b435, 32'h00000000} /* (30, 3, 24) {real, imag} */,
  {32'h44fb0dc0, 32'h00000000} /* (30, 3, 23) {real, imag} */,
  {32'h4551e79c, 32'h00000000} /* (30, 3, 22) {real, imag} */,
  {32'h455ba2fd, 32'h00000000} /* (30, 3, 21) {real, imag} */,
  {32'h4526cbf8, 32'h00000000} /* (30, 3, 20) {real, imag} */,
  {32'h44c1750f, 32'h00000000} /* (30, 3, 19) {real, imag} */,
  {32'h4489f3ee, 32'h00000000} /* (30, 3, 18) {real, imag} */,
  {32'h448d08cc, 32'h00000000} /* (30, 3, 17) {real, imag} */,
  {32'hc3c2e820, 32'h00000000} /* (30, 3, 16) {real, imag} */,
  {32'hc5061923, 32'h00000000} /* (30, 3, 15) {real, imag} */,
  {32'hc527483f, 32'h00000000} /* (30, 3, 14) {real, imag} */,
  {32'hc51070c5, 32'h00000000} /* (30, 3, 13) {real, imag} */,
  {32'hc598ed05, 32'h00000000} /* (30, 3, 12) {real, imag} */,
  {32'hc57dfa7c, 32'h00000000} /* (30, 3, 11) {real, imag} */,
  {32'hc55f1002, 32'h00000000} /* (30, 3, 10) {real, imag} */,
  {32'hc5187810, 32'h00000000} /* (30, 3, 9) {real, imag} */,
  {32'hc50facd7, 32'h00000000} /* (30, 3, 8) {real, imag} */,
  {32'hc51aa3e2, 32'h00000000} /* (30, 3, 7) {real, imag} */,
  {32'hc49e4a39, 32'h00000000} /* (30, 3, 6) {real, imag} */,
  {32'h428178e0, 32'h00000000} /* (30, 3, 5) {real, imag} */,
  {32'h44ebc624, 32'h00000000} /* (30, 3, 4) {real, imag} */,
  {32'h44dcde79, 32'h00000000} /* (30, 3, 3) {real, imag} */,
  {32'h454a0c1d, 32'h00000000} /* (30, 3, 2) {real, imag} */,
  {32'h450109b5, 32'h00000000} /* (30, 3, 1) {real, imag} */,
  {32'h44b4fd32, 32'h00000000} /* (30, 3, 0) {real, imag} */,
  {32'h449a2c99, 32'h00000000} /* (30, 2, 31) {real, imag} */,
  {32'h450998e6, 32'h00000000} /* (30, 2, 30) {real, imag} */,
  {32'h4512a204, 32'h00000000} /* (30, 2, 29) {real, imag} */,
  {32'h45204163, 32'h00000000} /* (30, 2, 28) {real, imag} */,
  {32'h44e6cc7a, 32'h00000000} /* (30, 2, 27) {real, imag} */,
  {32'h45526bd2, 32'h00000000} /* (30, 2, 26) {real, imag} */,
  {32'h450319c8, 32'h00000000} /* (30, 2, 25) {real, imag} */,
  {32'h4522e250, 32'h00000000} /* (30, 2, 24) {real, imag} */,
  {32'h45055cde, 32'h00000000} /* (30, 2, 23) {real, imag} */,
  {32'h45058bed, 32'h00000000} /* (30, 2, 22) {real, imag} */,
  {32'h453e0056, 32'h00000000} /* (30, 2, 21) {real, imag} */,
  {32'h45198ced, 32'h00000000} /* (30, 2, 20) {real, imag} */,
  {32'h44f2bf7e, 32'h00000000} /* (30, 2, 19) {real, imag} */,
  {32'h447e5b00, 32'h00000000} /* (30, 2, 18) {real, imag} */,
  {32'h4449ae86, 32'h00000000} /* (30, 2, 17) {real, imag} */,
  {32'hc3dbb898, 32'h00000000} /* (30, 2, 16) {real, imag} */,
  {32'hc50f24ca, 32'h00000000} /* (30, 2, 15) {real, imag} */,
  {32'hc50da446, 32'h00000000} /* (30, 2, 14) {real, imag} */,
  {32'hc515ccf0, 32'h00000000} /* (30, 2, 13) {real, imag} */,
  {32'hc56731fb, 32'h00000000} /* (30, 2, 12) {real, imag} */,
  {32'hc5679875, 32'h00000000} /* (30, 2, 11) {real, imag} */,
  {32'hc55092f6, 32'h00000000} /* (30, 2, 10) {real, imag} */,
  {32'hc548fca0, 32'h00000000} /* (30, 2, 9) {real, imag} */,
  {32'hc50d16b8, 32'h00000000} /* (30, 2, 8) {real, imag} */,
  {32'hc53e4c0c, 32'h00000000} /* (30, 2, 7) {real, imag} */,
  {32'hc50f307b, 32'h00000000} /* (30, 2, 6) {real, imag} */,
  {32'hc3594798, 32'h00000000} /* (30, 2, 5) {real, imag} */,
  {32'h4490e31a, 32'h00000000} /* (30, 2, 4) {real, imag} */,
  {32'h44f64b72, 32'h00000000} /* (30, 2, 3) {real, imag} */,
  {32'h44d9c654, 32'h00000000} /* (30, 2, 2) {real, imag} */,
  {32'h44b9e9a1, 32'h00000000} /* (30, 2, 1) {real, imag} */,
  {32'h44888d5e, 32'h00000000} /* (30, 2, 0) {real, imag} */,
  {32'h4485c541, 32'h00000000} /* (30, 1, 31) {real, imag} */,
  {32'h44d014f1, 32'h00000000} /* (30, 1, 30) {real, imag} */,
  {32'h44e5e108, 32'h00000000} /* (30, 1, 29) {real, imag} */,
  {32'h44c6ef08, 32'h00000000} /* (30, 1, 28) {real, imag} */,
  {32'h44ff184b, 32'h00000000} /* (30, 1, 27) {real, imag} */,
  {32'h44f284e5, 32'h00000000} /* (30, 1, 26) {real, imag} */,
  {32'h4532cb61, 32'h00000000} /* (30, 1, 25) {real, imag} */,
  {32'h451bb02e, 32'h00000000} /* (30, 1, 24) {real, imag} */,
  {32'h44d50601, 32'h00000000} /* (30, 1, 23) {real, imag} */,
  {32'h452ff7cd, 32'h00000000} /* (30, 1, 22) {real, imag} */,
  {32'h451f373c, 32'h00000000} /* (30, 1, 21) {real, imag} */,
  {32'h44d32075, 32'h00000000} /* (30, 1, 20) {real, imag} */,
  {32'h4505e1a2, 32'h00000000} /* (30, 1, 19) {real, imag} */,
  {32'h44b156ab, 32'h00000000} /* (30, 1, 18) {real, imag} */,
  {32'h44e47102, 32'h00000000} /* (30, 1, 17) {real, imag} */,
  {32'hc3dfcc94, 32'h00000000} /* (30, 1, 16) {real, imag} */,
  {32'hc51734b8, 32'h00000000} /* (30, 1, 15) {real, imag} */,
  {32'hc502f63c, 32'h00000000} /* (30, 1, 14) {real, imag} */,
  {32'hc51b055c, 32'h00000000} /* (30, 1, 13) {real, imag} */,
  {32'hc520514c, 32'h00000000} /* (30, 1, 12) {real, imag} */,
  {32'hc56e05c0, 32'h00000000} /* (30, 1, 11) {real, imag} */,
  {32'hc53efac4, 32'h00000000} /* (30, 1, 10) {real, imag} */,
  {32'hc51e1cef, 32'h00000000} /* (30, 1, 9) {real, imag} */,
  {32'hc51a4d0a, 32'h00000000} /* (30, 1, 8) {real, imag} */,
  {32'hc4bfc38b, 32'h00000000} /* (30, 1, 7) {real, imag} */,
  {32'hc5027d2b, 32'h00000000} /* (30, 1, 6) {real, imag} */,
  {32'hc2e58530, 32'h00000000} /* (30, 1, 5) {real, imag} */,
  {32'h44c16187, 32'h00000000} /* (30, 1, 4) {real, imag} */,
  {32'h44f84bab, 32'h00000000} /* (30, 1, 3) {real, imag} */,
  {32'h44ddf1ff, 32'h00000000} /* (30, 1, 2) {real, imag} */,
  {32'h4483559e, 32'h00000000} /* (30, 1, 1) {real, imag} */,
  {32'h44700388, 32'h00000000} /* (30, 1, 0) {real, imag} */,
  {32'h449daf96, 32'h00000000} /* (30, 0, 31) {real, imag} */,
  {32'h4482a987, 32'h00000000} /* (30, 0, 30) {real, imag} */,
  {32'h4462cede, 32'h00000000} /* (30, 0, 29) {real, imag} */,
  {32'h44c97516, 32'h00000000} /* (30, 0, 28) {real, imag} */,
  {32'h44ca475e, 32'h00000000} /* (30, 0, 27) {real, imag} */,
  {32'h4508646a, 32'h00000000} /* (30, 0, 26) {real, imag} */,
  {32'h450f3644, 32'h00000000} /* (30, 0, 25) {real, imag} */,
  {32'h45066fd6, 32'h00000000} /* (30, 0, 24) {real, imag} */,
  {32'h44fcf396, 32'h00000000} /* (30, 0, 23) {real, imag} */,
  {32'h451e63fe, 32'h00000000} /* (30, 0, 22) {real, imag} */,
  {32'h450ab950, 32'h00000000} /* (30, 0, 21) {real, imag} */,
  {32'h44a20ddf, 32'h00000000} /* (30, 0, 20) {real, imag} */,
  {32'h44853e97, 32'h00000000} /* (30, 0, 19) {real, imag} */,
  {32'h445deed8, 32'h00000000} /* (30, 0, 18) {real, imag} */,
  {32'h4457754b, 32'h00000000} /* (30, 0, 17) {real, imag} */,
  {32'hc42de0a7, 32'h00000000} /* (30, 0, 16) {real, imag} */,
  {32'hc4e3bfea, 32'h00000000} /* (30, 0, 15) {real, imag} */,
  {32'hc53e70c2, 32'h00000000} /* (30, 0, 14) {real, imag} */,
  {32'hc546c1aa, 32'h00000000} /* (30, 0, 13) {real, imag} */,
  {32'hc513e33f, 32'h00000000} /* (30, 0, 12) {real, imag} */,
  {32'hc50fc58b, 32'h00000000} /* (30, 0, 11) {real, imag} */,
  {32'hc4d920cc, 32'h00000000} /* (30, 0, 10) {real, imag} */,
  {32'hc48c7bd9, 32'h00000000} /* (30, 0, 9) {real, imag} */,
  {32'hc4989c04, 32'h00000000} /* (30, 0, 8) {real, imag} */,
  {32'hc4ad702e, 32'h00000000} /* (30, 0, 7) {real, imag} */,
  {32'hc3a28fe4, 32'h00000000} /* (30, 0, 6) {real, imag} */,
  {32'h43f5e862, 32'h00000000} /* (30, 0, 5) {real, imag} */,
  {32'h44b6de05, 32'h00000000} /* (30, 0, 4) {real, imag} */,
  {32'h44ce3579, 32'h00000000} /* (30, 0, 3) {real, imag} */,
  {32'h44ad4e70, 32'h00000000} /* (30, 0, 2) {real, imag} */,
  {32'h4484aa22, 32'h00000000} /* (30, 0, 1) {real, imag} */,
  {32'h4441079b, 32'h00000000} /* (30, 0, 0) {real, imag} */,
  {32'h445a0551, 32'h00000000} /* (29, 31, 31) {real, imag} */,
  {32'h446c8d76, 32'h00000000} /* (29, 31, 30) {real, imag} */,
  {32'h44e9d98a, 32'h00000000} /* (29, 31, 29) {real, imag} */,
  {32'h44bc7210, 32'h00000000} /* (29, 31, 28) {real, imag} */,
  {32'h44d5f686, 32'h00000000} /* (29, 31, 27) {real, imag} */,
  {32'h450ac642, 32'h00000000} /* (29, 31, 26) {real, imag} */,
  {32'h44fe4bb3, 32'h00000000} /* (29, 31, 25) {real, imag} */,
  {32'h4532850e, 32'h00000000} /* (29, 31, 24) {real, imag} */,
  {32'h4509dee2, 32'h00000000} /* (29, 31, 23) {real, imag} */,
  {32'h450e8e51, 32'h00000000} /* (29, 31, 22) {real, imag} */,
  {32'h44998edf, 32'h00000000} /* (29, 31, 21) {real, imag} */,
  {32'h44256caf, 32'h00000000} /* (29, 31, 20) {real, imag} */,
  {32'h4372bee0, 32'h00000000} /* (29, 31, 19) {real, imag} */,
  {32'hc45431b6, 32'h00000000} /* (29, 31, 18) {real, imag} */,
  {32'hc487272e, 32'h00000000} /* (29, 31, 17) {real, imag} */,
  {32'hc4f3a866, 32'h00000000} /* (29, 31, 16) {real, imag} */,
  {32'hc516917a, 32'h00000000} /* (29, 31, 15) {real, imag} */,
  {32'hc54e262c, 32'h00000000} /* (29, 31, 14) {real, imag} */,
  {32'hc54c2a97, 32'h00000000} /* (29, 31, 13) {real, imag} */,
  {32'hc557ea66, 32'h00000000} /* (29, 31, 12) {real, imag} */,
  {32'hc5227095, 32'h00000000} /* (29, 31, 11) {real, imag} */,
  {32'hc489bca4, 32'h00000000} /* (29, 31, 10) {real, imag} */,
  {32'h43d82414, 32'h00000000} /* (29, 31, 9) {real, imag} */,
  {32'h4366f818, 32'h00000000} /* (29, 31, 8) {real, imag} */,
  {32'h4454f95a, 32'h00000000} /* (29, 31, 7) {real, imag} */,
  {32'h44a02b6c, 32'h00000000} /* (29, 31, 6) {real, imag} */,
  {32'h448f9775, 32'h00000000} /* (29, 31, 5) {real, imag} */,
  {32'h44ef390c, 32'h00000000} /* (29, 31, 4) {real, imag} */,
  {32'h4501a7ae, 32'h00000000} /* (29, 31, 3) {real, imag} */,
  {32'h44eb52f7, 32'h00000000} /* (29, 31, 2) {real, imag} */,
  {32'h44e0e29e, 32'h00000000} /* (29, 31, 1) {real, imag} */,
  {32'h449298be, 32'h00000000} /* (29, 31, 0) {real, imag} */,
  {32'h4436b054, 32'h00000000} /* (29, 30, 31) {real, imag} */,
  {32'h44d147d2, 32'h00000000} /* (29, 30, 30) {real, imag} */,
  {32'h45049846, 32'h00000000} /* (29, 30, 29) {real, imag} */,
  {32'h452818b7, 32'h00000000} /* (29, 30, 28) {real, imag} */,
  {32'h45358b1d, 32'h00000000} /* (29, 30, 27) {real, imag} */,
  {32'h4532234c, 32'h00000000} /* (29, 30, 26) {real, imag} */,
  {32'h457229c6, 32'h00000000} /* (29, 30, 25) {real, imag} */,
  {32'h453f562c, 32'h00000000} /* (29, 30, 24) {real, imag} */,
  {32'h453f9dc0, 32'h00000000} /* (29, 30, 23) {real, imag} */,
  {32'h450c3412, 32'h00000000} /* (29, 30, 22) {real, imag} */,
  {32'h44a9c2af, 32'h00000000} /* (29, 30, 21) {real, imag} */,
  {32'hc3b83800, 32'h00000000} /* (29, 30, 20) {real, imag} */,
  {32'hc489ef64, 32'h00000000} /* (29, 30, 19) {real, imag} */,
  {32'hc4f3e28f, 32'h00000000} /* (29, 30, 18) {real, imag} */,
  {32'hc5341e0b, 32'h00000000} /* (29, 30, 17) {real, imag} */,
  {32'hc53f7857, 32'h00000000} /* (29, 30, 16) {real, imag} */,
  {32'hc555bf49, 32'h00000000} /* (29, 30, 15) {real, imag} */,
  {32'hc58027f4, 32'h00000000} /* (29, 30, 14) {real, imag} */,
  {32'hc5826607, 32'h00000000} /* (29, 30, 13) {real, imag} */,
  {32'hc56b4ed1, 32'h00000000} /* (29, 30, 12) {real, imag} */,
  {32'hc52eed3b, 32'h00000000} /* (29, 30, 11) {real, imag} */,
  {32'hc448b830, 32'h00000000} /* (29, 30, 10) {real, imag} */,
  {32'h450b9a1a, 32'h00000000} /* (29, 30, 9) {real, imag} */,
  {32'h45087032, 32'h00000000} /* (29, 30, 8) {real, imag} */,
  {32'h44c1b2f8, 32'h00000000} /* (29, 30, 7) {real, imag} */,
  {32'h4532ded8, 32'h00000000} /* (29, 30, 6) {real, imag} */,
  {32'h450f9608, 32'h00000000} /* (29, 30, 5) {real, imag} */,
  {32'h452f5792, 32'h00000000} /* (29, 30, 4) {real, imag} */,
  {32'h456876a8, 32'h00000000} /* (29, 30, 3) {real, imag} */,
  {32'h4520f022, 32'h00000000} /* (29, 30, 2) {real, imag} */,
  {32'h4536f093, 32'h00000000} /* (29, 30, 1) {real, imag} */,
  {32'h4501cca5, 32'h00000000} /* (29, 30, 0) {real, imag} */,
  {32'h4529f65d, 32'h00000000} /* (29, 29, 31) {real, imag} */,
  {32'h452e3f24, 32'h00000000} /* (29, 29, 30) {real, imag} */,
  {32'h44dc77d6, 32'h00000000} /* (29, 29, 29) {real, imag} */,
  {32'h450f9b2e, 32'h00000000} /* (29, 29, 28) {real, imag} */,
  {32'h452c53bc, 32'h00000000} /* (29, 29, 27) {real, imag} */,
  {32'h4558dbe1, 32'h00000000} /* (29, 29, 26) {real, imag} */,
  {32'h455d96e6, 32'h00000000} /* (29, 29, 25) {real, imag} */,
  {32'h45622348, 32'h00000000} /* (29, 29, 24) {real, imag} */,
  {32'h456aa4d2, 32'h00000000} /* (29, 29, 23) {real, imag} */,
  {32'h44cb0bb8, 32'h00000000} /* (29, 29, 22) {real, imag} */,
  {32'h448280f8, 32'h00000000} /* (29, 29, 21) {real, imag} */,
  {32'hc523f388, 32'h00000000} /* (29, 29, 20) {real, imag} */,
  {32'hc4e49d24, 32'h00000000} /* (29, 29, 19) {real, imag} */,
  {32'hc53fefb2, 32'h00000000} /* (29, 29, 18) {real, imag} */,
  {32'hc589a69c, 32'h00000000} /* (29, 29, 17) {real, imag} */,
  {32'hc55c77e2, 32'h00000000} /* (29, 29, 16) {real, imag} */,
  {32'hc58117b8, 32'h00000000} /* (29, 29, 15) {real, imag} */,
  {32'hc5bee0be, 32'h00000000} /* (29, 29, 14) {real, imag} */,
  {32'hc5a12d6a, 32'h00000000} /* (29, 29, 13) {real, imag} */,
  {32'hc54c21ca, 32'h00000000} /* (29, 29, 12) {real, imag} */,
  {32'hc4c14f50, 32'h00000000} /* (29, 29, 11) {real, imag} */,
  {32'h43be6450, 32'h00000000} /* (29, 29, 10) {real, imag} */,
  {32'h4501b628, 32'h00000000} /* (29, 29, 9) {real, imag} */,
  {32'h4538940c, 32'h00000000} /* (29, 29, 8) {real, imag} */,
  {32'h451bc5aa, 32'h00000000} /* (29, 29, 7) {real, imag} */,
  {32'h454a274c, 32'h00000000} /* (29, 29, 6) {real, imag} */,
  {32'h45471162, 32'h00000000} /* (29, 29, 5) {real, imag} */,
  {32'h454a517a, 32'h00000000} /* (29, 29, 4) {real, imag} */,
  {32'h45519450, 32'h00000000} /* (29, 29, 3) {real, imag} */,
  {32'h4505d528, 32'h00000000} /* (29, 29, 2) {real, imag} */,
  {32'h44f37ca4, 32'h00000000} /* (29, 29, 1) {real, imag} */,
  {32'h44b3b29c, 32'h00000000} /* (29, 29, 0) {real, imag} */,
  {32'h44d10a61, 32'h00000000} /* (29, 28, 31) {real, imag} */,
  {32'h45335978, 32'h00000000} /* (29, 28, 30) {real, imag} */,
  {32'h453955f2, 32'h00000000} /* (29, 28, 29) {real, imag} */,
  {32'h4520d966, 32'h00000000} /* (29, 28, 28) {real, imag} */,
  {32'h45292bf4, 32'h00000000} /* (29, 28, 27) {real, imag} */,
  {32'h45519d6e, 32'h00000000} /* (29, 28, 26) {real, imag} */,
  {32'h45486e02, 32'h00000000} /* (29, 28, 25) {real, imag} */,
  {32'h45287b50, 32'h00000000} /* (29, 28, 24) {real, imag} */,
  {32'h4512dc10, 32'h00000000} /* (29, 28, 23) {real, imag} */,
  {32'h4508e5d4, 32'h00000000} /* (29, 28, 22) {real, imag} */,
  {32'h44bc884a, 32'h00000000} /* (29, 28, 21) {real, imag} */,
  {32'hc48fc2c8, 32'h00000000} /* (29, 28, 20) {real, imag} */,
  {32'hc51779fb, 32'h00000000} /* (29, 28, 19) {real, imag} */,
  {32'hc554f044, 32'h00000000} /* (29, 28, 18) {real, imag} */,
  {32'hc566330e, 32'h00000000} /* (29, 28, 17) {real, imag} */,
  {32'hc544bfa0, 32'h00000000} /* (29, 28, 16) {real, imag} */,
  {32'hc58cc3cf, 32'h00000000} /* (29, 28, 15) {real, imag} */,
  {32'hc58de20b, 32'h00000000} /* (29, 28, 14) {real, imag} */,
  {32'hc5941980, 32'h00000000} /* (29, 28, 13) {real, imag} */,
  {32'hc5473fca, 32'h00000000} /* (29, 28, 12) {real, imag} */,
  {32'hc4c75ad0, 32'h00000000} /* (29, 28, 11) {real, imag} */,
  {32'h448e43d5, 32'h00000000} /* (29, 28, 10) {real, imag} */,
  {32'h453632ca, 32'h00000000} /* (29, 28, 9) {real, imag} */,
  {32'h4570c9e0, 32'h00000000} /* (29, 28, 8) {real, imag} */,
  {32'h4592bba0, 32'h00000000} /* (29, 28, 7) {real, imag} */,
  {32'h45519820, 32'h00000000} /* (29, 28, 6) {real, imag} */,
  {32'h454bab73, 32'h00000000} /* (29, 28, 5) {real, imag} */,
  {32'h454b30b0, 32'h00000000} /* (29, 28, 4) {real, imag} */,
  {32'h452aea1d, 32'h00000000} /* (29, 28, 3) {real, imag} */,
  {32'h45113aca, 32'h00000000} /* (29, 28, 2) {real, imag} */,
  {32'h44d6f691, 32'h00000000} /* (29, 28, 1) {real, imag} */,
  {32'h450c090c, 32'h00000000} /* (29, 28, 0) {real, imag} */,
  {32'h44f167b9, 32'h00000000} /* (29, 27, 31) {real, imag} */,
  {32'h4519652e, 32'h00000000} /* (29, 27, 30) {real, imag} */,
  {32'h45150050, 32'h00000000} /* (29, 27, 29) {real, imag} */,
  {32'h4521b187, 32'h00000000} /* (29, 27, 28) {real, imag} */,
  {32'h456eaf36, 32'h00000000} /* (29, 27, 27) {real, imag} */,
  {32'h45601e20, 32'h00000000} /* (29, 27, 26) {real, imag} */,
  {32'h457dc2b8, 32'h00000000} /* (29, 27, 25) {real, imag} */,
  {32'h45489856, 32'h00000000} /* (29, 27, 24) {real, imag} */,
  {32'h4504bf9d, 32'h00000000} /* (29, 27, 23) {real, imag} */,
  {32'h45150da6, 32'h00000000} /* (29, 27, 22) {real, imag} */,
  {32'h44937c0f, 32'h00000000} /* (29, 27, 21) {real, imag} */,
  {32'hc4a78bb3, 32'h00000000} /* (29, 27, 20) {real, imag} */,
  {32'hc56197f6, 32'h00000000} /* (29, 27, 19) {real, imag} */,
  {32'hc563ed25, 32'h00000000} /* (29, 27, 18) {real, imag} */,
  {32'hc5559b32, 32'h00000000} /* (29, 27, 17) {real, imag} */,
  {32'hc5714870, 32'h00000000} /* (29, 27, 16) {real, imag} */,
  {32'hc57312f0, 32'h00000000} /* (29, 27, 15) {real, imag} */,
  {32'hc589594e, 32'h00000000} /* (29, 27, 14) {real, imag} */,
  {32'hc584cf67, 32'h00000000} /* (29, 27, 13) {real, imag} */,
  {32'hc5185027, 32'h00000000} /* (29, 27, 12) {real, imag} */,
  {32'hc487096b, 32'h00000000} /* (29, 27, 11) {real, imag} */,
  {32'h44b23641, 32'h00000000} /* (29, 27, 10) {real, imag} */,
  {32'h456ca590, 32'h00000000} /* (29, 27, 9) {real, imag} */,
  {32'h4591120e, 32'h00000000} /* (29, 27, 8) {real, imag} */,
  {32'h45936166, 32'h00000000} /* (29, 27, 7) {real, imag} */,
  {32'h4593ece3, 32'h00000000} /* (29, 27, 6) {real, imag} */,
  {32'h4572667c, 32'h00000000} /* (29, 27, 5) {real, imag} */,
  {32'h4546d770, 32'h00000000} /* (29, 27, 4) {real, imag} */,
  {32'h4581d3ab, 32'h00000000} /* (29, 27, 3) {real, imag} */,
  {32'h45114437, 32'h00000000} /* (29, 27, 2) {real, imag} */,
  {32'h44f283b5, 32'h00000000} /* (29, 27, 1) {real, imag} */,
  {32'h44d5ed6c, 32'h00000000} /* (29, 27, 0) {real, imag} */,
  {32'h44d12e6d, 32'h00000000} /* (29, 26, 31) {real, imag} */,
  {32'h44f792a2, 32'h00000000} /* (29, 26, 30) {real, imag} */,
  {32'h45492894, 32'h00000000} /* (29, 26, 29) {real, imag} */,
  {32'h453a8df1, 32'h00000000} /* (29, 26, 28) {real, imag} */,
  {32'h45598062, 32'h00000000} /* (29, 26, 27) {real, imag} */,
  {32'h456072e0, 32'h00000000} /* (29, 26, 26) {real, imag} */,
  {32'h453ac680, 32'h00000000} /* (29, 26, 25) {real, imag} */,
  {32'h4573e29c, 32'h00000000} /* (29, 26, 24) {real, imag} */,
  {32'h453117aa, 32'h00000000} /* (29, 26, 23) {real, imag} */,
  {32'h44c2dbd4, 32'h00000000} /* (29, 26, 22) {real, imag} */,
  {32'h440c3b14, 32'h00000000} /* (29, 26, 21) {real, imag} */,
  {32'hc4fc749e, 32'h00000000} /* (29, 26, 20) {real, imag} */,
  {32'hc53492f9, 32'h00000000} /* (29, 26, 19) {real, imag} */,
  {32'hc55e4fc8, 32'h00000000} /* (29, 26, 18) {real, imag} */,
  {32'hc569bf8c, 32'h00000000} /* (29, 26, 17) {real, imag} */,
  {32'hc58c093e, 32'h00000000} /* (29, 26, 16) {real, imag} */,
  {32'hc58e43e7, 32'h00000000} /* (29, 26, 15) {real, imag} */,
  {32'hc5824dfc, 32'h00000000} /* (29, 26, 14) {real, imag} */,
  {32'hc5630c60, 32'h00000000} /* (29, 26, 13) {real, imag} */,
  {32'hc53a9215, 32'h00000000} /* (29, 26, 12) {real, imag} */,
  {32'hc427d048, 32'h00000000} /* (29, 26, 11) {real, imag} */,
  {32'h4463035a, 32'h00000000} /* (29, 26, 10) {real, imag} */,
  {32'h452d1b28, 32'h00000000} /* (29, 26, 9) {real, imag} */,
  {32'h456e5018, 32'h00000000} /* (29, 26, 8) {real, imag} */,
  {32'h457c5c36, 32'h00000000} /* (29, 26, 7) {real, imag} */,
  {32'h456f5a78, 32'h00000000} /* (29, 26, 6) {real, imag} */,
  {32'h4577207b, 32'h00000000} /* (29, 26, 5) {real, imag} */,
  {32'h455e4d47, 32'h00000000} /* (29, 26, 4) {real, imag} */,
  {32'h45708851, 32'h00000000} /* (29, 26, 3) {real, imag} */,
  {32'h45155318, 32'h00000000} /* (29, 26, 2) {real, imag} */,
  {32'h44f50e21, 32'h00000000} /* (29, 26, 1) {real, imag} */,
  {32'h44fc585d, 32'h00000000} /* (29, 26, 0) {real, imag} */,
  {32'h4504b7b8, 32'h00000000} /* (29, 25, 31) {real, imag} */,
  {32'h450de79c, 32'h00000000} /* (29, 25, 30) {real, imag} */,
  {32'h453705f9, 32'h00000000} /* (29, 25, 29) {real, imag} */,
  {32'h4530db46, 32'h00000000} /* (29, 25, 28) {real, imag} */,
  {32'h454ca491, 32'h00000000} /* (29, 25, 27) {real, imag} */,
  {32'h45772382, 32'h00000000} /* (29, 25, 26) {real, imag} */,
  {32'h4563c792, 32'h00000000} /* (29, 25, 25) {real, imag} */,
  {32'h45469d72, 32'h00000000} /* (29, 25, 24) {real, imag} */,
  {32'h45344782, 32'h00000000} /* (29, 25, 23) {real, imag} */,
  {32'h45062259, 32'h00000000} /* (29, 25, 22) {real, imag} */,
  {32'h4407fd5c, 32'h00000000} /* (29, 25, 21) {real, imag} */,
  {32'hc4c07b1a, 32'h00000000} /* (29, 25, 20) {real, imag} */,
  {32'hc504d34d, 32'h00000000} /* (29, 25, 19) {real, imag} */,
  {32'hc561788c, 32'h00000000} /* (29, 25, 18) {real, imag} */,
  {32'hc54a317a, 32'h00000000} /* (29, 25, 17) {real, imag} */,
  {32'hc563d11e, 32'h00000000} /* (29, 25, 16) {real, imag} */,
  {32'hc59d05aa, 32'h00000000} /* (29, 25, 15) {real, imag} */,
  {32'hc5a5556e, 32'h00000000} /* (29, 25, 14) {real, imag} */,
  {32'hc584e47a, 32'h00000000} /* (29, 25, 13) {real, imag} */,
  {32'hc511aa92, 32'h00000000} /* (29, 25, 12) {real, imag} */,
  {32'hc4c35b26, 32'h00000000} /* (29, 25, 11) {real, imag} */,
  {32'h441558c8, 32'h00000000} /* (29, 25, 10) {real, imag} */,
  {32'h45523cac, 32'h00000000} /* (29, 25, 9) {real, imag} */,
  {32'h4576f12a, 32'h00000000} /* (29, 25, 8) {real, imag} */,
  {32'h457c5252, 32'h00000000} /* (29, 25, 7) {real, imag} */,
  {32'h45807269, 32'h00000000} /* (29, 25, 6) {real, imag} */,
  {32'h455ecf5f, 32'h00000000} /* (29, 25, 5) {real, imag} */,
  {32'h45889116, 32'h00000000} /* (29, 25, 4) {real, imag} */,
  {32'h4522e1ef, 32'h00000000} /* (29, 25, 3) {real, imag} */,
  {32'h450cd6b6, 32'h00000000} /* (29, 25, 2) {real, imag} */,
  {32'h44e77bb0, 32'h00000000} /* (29, 25, 1) {real, imag} */,
  {32'h44d5f9b5, 32'h00000000} /* (29, 25, 0) {real, imag} */,
  {32'h44e94e11, 32'h00000000} /* (29, 24, 31) {real, imag} */,
  {32'h451787c1, 32'h00000000} /* (29, 24, 30) {real, imag} */,
  {32'h44b8cec2, 32'h00000000} /* (29, 24, 29) {real, imag} */,
  {32'h450da6a8, 32'h00000000} /* (29, 24, 28) {real, imag} */,
  {32'h45345d4b, 32'h00000000} /* (29, 24, 27) {real, imag} */,
  {32'h455e9135, 32'h00000000} /* (29, 24, 26) {real, imag} */,
  {32'h459c5cf7, 32'h00000000} /* (29, 24, 25) {real, imag} */,
  {32'h4568b5e7, 32'h00000000} /* (29, 24, 24) {real, imag} */,
  {32'h453369ae, 32'h00000000} /* (29, 24, 23) {real, imag} */,
  {32'h45104c8c, 32'h00000000} /* (29, 24, 22) {real, imag} */,
  {32'h44a4b8e8, 32'h00000000} /* (29, 24, 21) {real, imag} */,
  {32'hc4e06162, 32'h00000000} /* (29, 24, 20) {real, imag} */,
  {32'hc52f52f9, 32'h00000000} /* (29, 24, 19) {real, imag} */,
  {32'hc5600546, 32'h00000000} /* (29, 24, 18) {real, imag} */,
  {32'hc56681db, 32'h00000000} /* (29, 24, 17) {real, imag} */,
  {32'hc57ce7ad, 32'h00000000} /* (29, 24, 16) {real, imag} */,
  {32'hc57759c2, 32'h00000000} /* (29, 24, 15) {real, imag} */,
  {32'hc592126a, 32'h00000000} /* (29, 24, 14) {real, imag} */,
  {32'hc5531d5f, 32'h00000000} /* (29, 24, 13) {real, imag} */,
  {32'hc4efadb4, 32'h00000000} /* (29, 24, 12) {real, imag} */,
  {32'hc49e4832, 32'h00000000} /* (29, 24, 11) {real, imag} */,
  {32'h4486fb06, 32'h00000000} /* (29, 24, 10) {real, imag} */,
  {32'h454b33b2, 32'h00000000} /* (29, 24, 9) {real, imag} */,
  {32'h458cfc4e, 32'h00000000} /* (29, 24, 8) {real, imag} */,
  {32'h459658eb, 32'h00000000} /* (29, 24, 7) {real, imag} */,
  {32'h459fa0d9, 32'h00000000} /* (29, 24, 6) {real, imag} */,
  {32'h4561e4d6, 32'h00000000} /* (29, 24, 5) {real, imag} */,
  {32'h4540469f, 32'h00000000} /* (29, 24, 4) {real, imag} */,
  {32'h455bacad, 32'h00000000} /* (29, 24, 3) {real, imag} */,
  {32'h454fd95a, 32'h00000000} /* (29, 24, 2) {real, imag} */,
  {32'h44f345da, 32'h00000000} /* (29, 24, 1) {real, imag} */,
  {32'h44be2f8a, 32'h00000000} /* (29, 24, 0) {real, imag} */,
  {32'h44f04c16, 32'h00000000} /* (29, 23, 31) {real, imag} */,
  {32'h44b8abaa, 32'h00000000} /* (29, 23, 30) {real, imag} */,
  {32'h44e137ac, 32'h00000000} /* (29, 23, 29) {real, imag} */,
  {32'h44cdfb5f, 32'h00000000} /* (29, 23, 28) {real, imag} */,
  {32'h44e8d642, 32'h00000000} /* (29, 23, 27) {real, imag} */,
  {32'h454f7efd, 32'h00000000} /* (29, 23, 26) {real, imag} */,
  {32'h45331eab, 32'h00000000} /* (29, 23, 25) {real, imag} */,
  {32'h45027220, 32'h00000000} /* (29, 23, 24) {real, imag} */,
  {32'h45112083, 32'h00000000} /* (29, 23, 23) {real, imag} */,
  {32'h45159a40, 32'h00000000} /* (29, 23, 22) {real, imag} */,
  {32'h446c9c5a, 32'h00000000} /* (29, 23, 21) {real, imag} */,
  {32'hc4507df6, 32'h00000000} /* (29, 23, 20) {real, imag} */,
  {32'hc516e737, 32'h00000000} /* (29, 23, 19) {real, imag} */,
  {32'hc5882274, 32'h00000000} /* (29, 23, 18) {real, imag} */,
  {32'hc534b77f, 32'h00000000} /* (29, 23, 17) {real, imag} */,
  {32'hc543c44c, 32'h00000000} /* (29, 23, 16) {real, imag} */,
  {32'hc52dd4bf, 32'h00000000} /* (29, 23, 15) {real, imag} */,
  {32'hc53797a1, 32'h00000000} /* (29, 23, 14) {real, imag} */,
  {32'hc50c50e8, 32'h00000000} /* (29, 23, 13) {real, imag} */,
  {32'hc4cded87, 32'h00000000} /* (29, 23, 12) {real, imag} */,
  {32'hc40df6b8, 32'h00000000} /* (29, 23, 11) {real, imag} */,
  {32'h441fc454, 32'h00000000} /* (29, 23, 10) {real, imag} */,
  {32'h44f878fb, 32'h00000000} /* (29, 23, 9) {real, imag} */,
  {32'h456ff5ba, 32'h00000000} /* (29, 23, 8) {real, imag} */,
  {32'h456d9c35, 32'h00000000} /* (29, 23, 7) {real, imag} */,
  {32'h4571e7ec, 32'h00000000} /* (29, 23, 6) {real, imag} */,
  {32'h455393e0, 32'h00000000} /* (29, 23, 5) {real, imag} */,
  {32'h454496b0, 32'h00000000} /* (29, 23, 4) {real, imag} */,
  {32'h45481cdf, 32'h00000000} /* (29, 23, 3) {real, imag} */,
  {32'h450defd9, 32'h00000000} /* (29, 23, 2) {real, imag} */,
  {32'h44eb0946, 32'h00000000} /* (29, 23, 1) {real, imag} */,
  {32'h448b8244, 32'h00000000} /* (29, 23, 0) {real, imag} */,
  {32'h44a51244, 32'h00000000} /* (29, 22, 31) {real, imag} */,
  {32'h44118901, 32'h00000000} /* (29, 22, 30) {real, imag} */,
  {32'h44955cdc, 32'h00000000} /* (29, 22, 29) {real, imag} */,
  {32'h449d3a43, 32'h00000000} /* (29, 22, 28) {real, imag} */,
  {32'h44491714, 32'h00000000} /* (29, 22, 27) {real, imag} */,
  {32'h44f1306a, 32'h00000000} /* (29, 22, 26) {real, imag} */,
  {32'h44c69233, 32'h00000000} /* (29, 22, 25) {real, imag} */,
  {32'h44e67ba1, 32'h00000000} /* (29, 22, 24) {real, imag} */,
  {32'h451a6e5a, 32'h00000000} /* (29, 22, 23) {real, imag} */,
  {32'h44de6495, 32'h00000000} /* (29, 22, 22) {real, imag} */,
  {32'h449cf5ba, 32'h00000000} /* (29, 22, 21) {real, imag} */,
  {32'hc4ba2be7, 32'h00000000} /* (29, 22, 20) {real, imag} */,
  {32'hc44588a8, 32'h00000000} /* (29, 22, 19) {real, imag} */,
  {32'hc4aa3aae, 32'h00000000} /* (29, 22, 18) {real, imag} */,
  {32'hc4d316f1, 32'h00000000} /* (29, 22, 17) {real, imag} */,
  {32'hc4d25b61, 32'h00000000} /* (29, 22, 16) {real, imag} */,
  {32'hc4d81026, 32'h00000000} /* (29, 22, 15) {real, imag} */,
  {32'hc4d132e8, 32'h00000000} /* (29, 22, 14) {real, imag} */,
  {32'hc4e26fb6, 32'h00000000} /* (29, 22, 13) {real, imag} */,
  {32'hc48c5507, 32'h00000000} /* (29, 22, 12) {real, imag} */,
  {32'hc439812c, 32'h00000000} /* (29, 22, 11) {real, imag} */,
  {32'h4422faed, 32'h00000000} /* (29, 22, 10) {real, imag} */,
  {32'h448a2825, 32'h00000000} /* (29, 22, 9) {real, imag} */,
  {32'h44fdb3f5, 32'h00000000} /* (29, 22, 8) {real, imag} */,
  {32'h4526b60a, 32'h00000000} /* (29, 22, 7) {real, imag} */,
  {32'h45184948, 32'h00000000} /* (29, 22, 6) {real, imag} */,
  {32'h45354db3, 32'h00000000} /* (29, 22, 5) {real, imag} */,
  {32'h451234f0, 32'h00000000} /* (29, 22, 4) {real, imag} */,
  {32'h450caffc, 32'h00000000} /* (29, 22, 3) {real, imag} */,
  {32'h453baea7, 32'h00000000} /* (29, 22, 2) {real, imag} */,
  {32'h45099444, 32'h00000000} /* (29, 22, 1) {real, imag} */,
  {32'h445d548e, 32'h00000000} /* (29, 22, 0) {real, imag} */,
  {32'hc2b30010, 32'h00000000} /* (29, 21, 31) {real, imag} */,
  {32'h436a53a2, 32'h00000000} /* (29, 21, 30) {real, imag} */,
  {32'h42f30f50, 32'h00000000} /* (29, 21, 29) {real, imag} */,
  {32'hc3fab5e0, 32'h00000000} /* (29, 21, 28) {real, imag} */,
  {32'hc4069919, 32'h00000000} /* (29, 21, 27) {real, imag} */,
  {32'hc455289e, 32'h00000000} /* (29, 21, 26) {real, imag} */,
  {32'hc3caa203, 32'h00000000} /* (29, 21, 25) {real, imag} */,
  {32'h444a7e3b, 32'h00000000} /* (29, 21, 24) {real, imag} */,
  {32'hc378eb88, 32'h00000000} /* (29, 21, 23) {real, imag} */,
  {32'h43eb6423, 32'h00000000} /* (29, 21, 22) {real, imag} */,
  {32'h43d317b0, 32'h00000000} /* (29, 21, 21) {real, imag} */,
  {32'hc3641061, 32'h00000000} /* (29, 21, 20) {real, imag} */,
  {32'hc3d59bfd, 32'h00000000} /* (29, 21, 19) {real, imag} */,
  {32'hc286dd50, 32'h00000000} /* (29, 21, 18) {real, imag} */,
  {32'hc3f26b22, 32'h00000000} /* (29, 21, 17) {real, imag} */,
  {32'hc401ad79, 32'h00000000} /* (29, 21, 16) {real, imag} */,
  {32'hc4992f9c, 32'h00000000} /* (29, 21, 15) {real, imag} */,
  {32'hc435a290, 32'h00000000} /* (29, 21, 14) {real, imag} */,
  {32'h42155188, 32'h00000000} /* (29, 21, 13) {real, imag} */,
  {32'h447e6036, 32'h00000000} /* (29, 21, 12) {real, imag} */,
  {32'h44411377, 32'h00000000} /* (29, 21, 11) {real, imag} */,
  {32'h448f295f, 32'h00000000} /* (29, 21, 10) {real, imag} */,
  {32'h446fe848, 32'h00000000} /* (29, 21, 9) {real, imag} */,
  {32'h4377f384, 32'h00000000} /* (29, 21, 8) {real, imag} */,
  {32'h44788050, 32'h00000000} /* (29, 21, 7) {real, imag} */,
  {32'hc38dfd95, 32'h00000000} /* (29, 21, 6) {real, imag} */,
  {32'hc36b2b9b, 32'h00000000} /* (29, 21, 5) {real, imag} */,
  {32'h427dc224, 32'h00000000} /* (29, 21, 4) {real, imag} */,
  {32'h4390e187, 32'h00000000} /* (29, 21, 3) {real, imag} */,
  {32'h43b6feae, 32'h00000000} /* (29, 21, 2) {real, imag} */,
  {32'h42964500, 32'h00000000} /* (29, 21, 1) {real, imag} */,
  {32'hc312ae43, 32'h00000000} /* (29, 21, 0) {real, imag} */,
  {32'hc4d5dd6e, 32'h00000000} /* (29, 20, 31) {real, imag} */,
  {32'hc4c26e67, 32'h00000000} /* (29, 20, 30) {real, imag} */,
  {32'hc50cf5a8, 32'h00000000} /* (29, 20, 29) {real, imag} */,
  {32'hc53b526a, 32'h00000000} /* (29, 20, 28) {real, imag} */,
  {32'hc5135447, 32'h00000000} /* (29, 20, 27) {real, imag} */,
  {32'hc517be4b, 32'h00000000} /* (29, 20, 26) {real, imag} */,
  {32'hc50f8a8c, 32'h00000000} /* (29, 20, 25) {real, imag} */,
  {32'hc51b1d1d, 32'h00000000} /* (29, 20, 24) {real, imag} */,
  {32'hc4d4b9fa, 32'h00000000} /* (29, 20, 23) {real, imag} */,
  {32'hc49342e0, 32'h00000000} /* (29, 20, 22) {real, imag} */,
  {32'hc3574288, 32'h00000000} /* (29, 20, 21) {real, imag} */,
  {32'h446b7e06, 32'h00000000} /* (29, 20, 20) {real, imag} */,
  {32'h44a7f333, 32'h00000000} /* (29, 20, 19) {real, imag} */,
  {32'h44fd4ff2, 32'h00000000} /* (29, 20, 18) {real, imag} */,
  {32'h44d82f3c, 32'h00000000} /* (29, 20, 17) {real, imag} */,
  {32'h44d532dd, 32'h00000000} /* (29, 20, 16) {real, imag} */,
  {32'h44e37fbe, 32'h00000000} /* (29, 20, 15) {real, imag} */,
  {32'h450af1ca, 32'h00000000} /* (29, 20, 14) {real, imag} */,
  {32'h451d6ae0, 32'h00000000} /* (29, 20, 13) {real, imag} */,
  {32'h44d84be4, 32'h00000000} /* (29, 20, 12) {real, imag} */,
  {32'h44983770, 32'h00000000} /* (29, 20, 11) {real, imag} */,
  {32'h420194c0, 32'h00000000} /* (29, 20, 10) {real, imag} */,
  {32'hc486b3cb, 32'h00000000} /* (29, 20, 9) {real, imag} */,
  {32'hc48cea96, 32'h00000000} /* (29, 20, 8) {real, imag} */,
  {32'hc4cfbdd2, 32'h00000000} /* (29, 20, 7) {real, imag} */,
  {32'hc5352a70, 32'h00000000} /* (29, 20, 6) {real, imag} */,
  {32'hc5338e80, 32'h00000000} /* (29, 20, 5) {real, imag} */,
  {32'hc508f9b4, 32'h00000000} /* (29, 20, 4) {real, imag} */,
  {32'hc560f400, 32'h00000000} /* (29, 20, 3) {real, imag} */,
  {32'hc53f7e8b, 32'h00000000} /* (29, 20, 2) {real, imag} */,
  {32'hc509fbbe, 32'h00000000} /* (29, 20, 1) {real, imag} */,
  {32'hc49b9001, 32'h00000000} /* (29, 20, 0) {real, imag} */,
  {32'hc55ef49c, 32'h00000000} /* (29, 19, 31) {real, imag} */,
  {32'hc53514d0, 32'h00000000} /* (29, 19, 30) {real, imag} */,
  {32'hc582ee92, 32'h00000000} /* (29, 19, 29) {real, imag} */,
  {32'hc557329a, 32'h00000000} /* (29, 19, 28) {real, imag} */,
  {32'hc5481d02, 32'h00000000} /* (29, 19, 27) {real, imag} */,
  {32'hc5211771, 32'h00000000} /* (29, 19, 26) {real, imag} */,
  {32'hc53d0ae4, 32'h00000000} /* (29, 19, 25) {real, imag} */,
  {32'hc50ee43e, 32'h00000000} /* (29, 19, 24) {real, imag} */,
  {32'hc5148840, 32'h00000000} /* (29, 19, 23) {real, imag} */,
  {32'hc541e8bf, 32'h00000000} /* (29, 19, 22) {real, imag} */,
  {32'hc2074400, 32'h00000000} /* (29, 19, 21) {real, imag} */,
  {32'h44d357ba, 32'h00000000} /* (29, 19, 20) {real, imag} */,
  {32'h4505c094, 32'h00000000} /* (29, 19, 19) {real, imag} */,
  {32'h450c881e, 32'h00000000} /* (29, 19, 18) {real, imag} */,
  {32'h4552060a, 32'h00000000} /* (29, 19, 17) {real, imag} */,
  {32'h45399cf8, 32'h00000000} /* (29, 19, 16) {real, imag} */,
  {32'h453091ac, 32'h00000000} /* (29, 19, 15) {real, imag} */,
  {32'h455e315a, 32'h00000000} /* (29, 19, 14) {real, imag} */,
  {32'h455f0858, 32'h00000000} /* (29, 19, 13) {real, imag} */,
  {32'h4544dbd4, 32'h00000000} /* (29, 19, 12) {real, imag} */,
  {32'h44fac5b9, 32'h00000000} /* (29, 19, 11) {real, imag} */,
  {32'hc3137750, 32'h00000000} /* (29, 19, 10) {real, imag} */,
  {32'hc4dde80b, 32'h00000000} /* (29, 19, 9) {real, imag} */,
  {32'hc554885c, 32'h00000000} /* (29, 19, 8) {real, imag} */,
  {32'hc56dc5a8, 32'h00000000} /* (29, 19, 7) {real, imag} */,
  {32'hc52a0661, 32'h00000000} /* (29, 19, 6) {real, imag} */,
  {32'hc5616e80, 32'h00000000} /* (29, 19, 5) {real, imag} */,
  {32'hc565a5a3, 32'h00000000} /* (29, 19, 4) {real, imag} */,
  {32'hc53260f8, 32'h00000000} /* (29, 19, 3) {real, imag} */,
  {32'hc57a81c2, 32'h00000000} /* (29, 19, 2) {real, imag} */,
  {32'hc561a034, 32'h00000000} /* (29, 19, 1) {real, imag} */,
  {32'hc52a6492, 32'h00000000} /* (29, 19, 0) {real, imag} */,
  {32'hc575c79f, 32'h00000000} /* (29, 18, 31) {real, imag} */,
  {32'hc56bf944, 32'h00000000} /* (29, 18, 30) {real, imag} */,
  {32'hc57ac56d, 32'h00000000} /* (29, 18, 29) {real, imag} */,
  {32'hc585be49, 32'h00000000} /* (29, 18, 28) {real, imag} */,
  {32'hc58d9767, 32'h00000000} /* (29, 18, 27) {real, imag} */,
  {32'hc581d586, 32'h00000000} /* (29, 18, 26) {real, imag} */,
  {32'hc5511aea, 32'h00000000} /* (29, 18, 25) {real, imag} */,
  {32'hc5457374, 32'h00000000} /* (29, 18, 24) {real, imag} */,
  {32'hc5754296, 32'h00000000} /* (29, 18, 23) {real, imag} */,
  {32'hc53f184a, 32'h00000000} /* (29, 18, 22) {real, imag} */,
  {32'hc4943c10, 32'h00000000} /* (29, 18, 21) {real, imag} */,
  {32'h44876cb3, 32'h00000000} /* (29, 18, 20) {real, imag} */,
  {32'h4521c72c, 32'h00000000} /* (29, 18, 19) {real, imag} */,
  {32'h4586ea5c, 32'h00000000} /* (29, 18, 18) {real, imag} */,
  {32'h4538c816, 32'h00000000} /* (29, 18, 17) {real, imag} */,
  {32'h456c8955, 32'h00000000} /* (29, 18, 16) {real, imag} */,
  {32'h45714df9, 32'h00000000} /* (29, 18, 15) {real, imag} */,
  {32'h45670b0e, 32'h00000000} /* (29, 18, 14) {real, imag} */,
  {32'h45528595, 32'h00000000} /* (29, 18, 13) {real, imag} */,
  {32'h4533a9da, 32'h00000000} /* (29, 18, 12) {real, imag} */,
  {32'h44df03b9, 32'h00000000} /* (29, 18, 11) {real, imag} */,
  {32'hc46226d8, 32'h00000000} /* (29, 18, 10) {real, imag} */,
  {32'hc550bc02, 32'h00000000} /* (29, 18, 9) {real, imag} */,
  {32'hc539e9b0, 32'h00000000} /* (29, 18, 8) {real, imag} */,
  {32'hc53e6524, 32'h00000000} /* (29, 18, 7) {real, imag} */,
  {32'hc565f6b2, 32'h00000000} /* (29, 18, 6) {real, imag} */,
  {32'hc567d210, 32'h00000000} /* (29, 18, 5) {real, imag} */,
  {32'hc58d4daf, 32'h00000000} /* (29, 18, 4) {real, imag} */,
  {32'hc591dc91, 32'h00000000} /* (29, 18, 3) {real, imag} */,
  {32'hc583d4dc, 32'h00000000} /* (29, 18, 2) {real, imag} */,
  {32'hc589c406, 32'h00000000} /* (29, 18, 1) {real, imag} */,
  {32'hc58af824, 32'h00000000} /* (29, 18, 0) {real, imag} */,
  {32'hc571df38, 32'h00000000} /* (29, 17, 31) {real, imag} */,
  {32'hc5a56b03, 32'h00000000} /* (29, 17, 30) {real, imag} */,
  {32'hc5896f22, 32'h00000000} /* (29, 17, 29) {real, imag} */,
  {32'hc5a9757d, 32'h00000000} /* (29, 17, 28) {real, imag} */,
  {32'hc5981c53, 32'h00000000} /* (29, 17, 27) {real, imag} */,
  {32'hc59da4db, 32'h00000000} /* (29, 17, 26) {real, imag} */,
  {32'hc56ef127, 32'h00000000} /* (29, 17, 25) {real, imag} */,
  {32'hc5728a19, 32'h00000000} /* (29, 17, 24) {real, imag} */,
  {32'hc576ae46, 32'h00000000} /* (29, 17, 23) {real, imag} */,
  {32'hc534729e, 32'h00000000} /* (29, 17, 22) {real, imag} */,
  {32'hc50f7e0e, 32'h00000000} /* (29, 17, 21) {real, imag} */,
  {32'h4360a6f0, 32'h00000000} /* (29, 17, 20) {real, imag} */,
  {32'h45152085, 32'h00000000} /* (29, 17, 19) {real, imag} */,
  {32'h4537970c, 32'h00000000} /* (29, 17, 18) {real, imag} */,
  {32'h459d4bb7, 32'h00000000} /* (29, 17, 17) {real, imag} */,
  {32'h45755eac, 32'h00000000} /* (29, 17, 16) {real, imag} */,
  {32'h45836a2f, 32'h00000000} /* (29, 17, 15) {real, imag} */,
  {32'h4591dfe3, 32'h00000000} /* (29, 17, 14) {real, imag} */,
  {32'h453884de, 32'h00000000} /* (29, 17, 13) {real, imag} */,
  {32'h45296160, 32'h00000000} /* (29, 17, 12) {real, imag} */,
  {32'h447968b8, 32'h00000000} /* (29, 17, 11) {real, imag} */,
  {32'hc420b0c8, 32'h00000000} /* (29, 17, 10) {real, imag} */,
  {32'hc5077759, 32'h00000000} /* (29, 17, 9) {real, imag} */,
  {32'hc56f4ddb, 32'h00000000} /* (29, 17, 8) {real, imag} */,
  {32'hc57d6026, 32'h00000000} /* (29, 17, 7) {real, imag} */,
  {32'hc580e07b, 32'h00000000} /* (29, 17, 6) {real, imag} */,
  {32'hc56d6ea8, 32'h00000000} /* (29, 17, 5) {real, imag} */,
  {32'hc58994fa, 32'h00000000} /* (29, 17, 4) {real, imag} */,
  {32'hc59395ea, 32'h00000000} /* (29, 17, 3) {real, imag} */,
  {32'hc58798d0, 32'h00000000} /* (29, 17, 2) {real, imag} */,
  {32'hc57520e6, 32'h00000000} /* (29, 17, 1) {real, imag} */,
  {32'hc552da6a, 32'h00000000} /* (29, 17, 0) {real, imag} */,
  {32'hc55a89c0, 32'h00000000} /* (29, 16, 31) {real, imag} */,
  {32'hc594057d, 32'h00000000} /* (29, 16, 30) {real, imag} */,
  {32'hc58787bd, 32'h00000000} /* (29, 16, 29) {real, imag} */,
  {32'hc58e917b, 32'h00000000} /* (29, 16, 28) {real, imag} */,
  {32'hc5ad24c2, 32'h00000000} /* (29, 16, 27) {real, imag} */,
  {32'hc56283a5, 32'h00000000} /* (29, 16, 26) {real, imag} */,
  {32'hc580d9b3, 32'h00000000} /* (29, 16, 25) {real, imag} */,
  {32'hc5910b99, 32'h00000000} /* (29, 16, 24) {real, imag} */,
  {32'hc55d1505, 32'h00000000} /* (29, 16, 23) {real, imag} */,
  {32'hc51f212b, 32'h00000000} /* (29, 16, 22) {real, imag} */,
  {32'hc4de8b54, 32'h00000000} /* (29, 16, 21) {real, imag} */,
  {32'h449b50e3, 32'h00000000} /* (29, 16, 20) {real, imag} */,
  {32'h4520c0ce, 32'h00000000} /* (29, 16, 19) {real, imag} */,
  {32'h4537e1b5, 32'h00000000} /* (29, 16, 18) {real, imag} */,
  {32'h456e460e, 32'h00000000} /* (29, 16, 17) {real, imag} */,
  {32'h45873dc5, 32'h00000000} /* (29, 16, 16) {real, imag} */,
  {32'h4596add8, 32'h00000000} /* (29, 16, 15) {real, imag} */,
  {32'h4579d54e, 32'h00000000} /* (29, 16, 14) {real, imag} */,
  {32'h454cb76a, 32'h00000000} /* (29, 16, 13) {real, imag} */,
  {32'h450068d8, 32'h00000000} /* (29, 16, 12) {real, imag} */,
  {32'h444b42ac, 32'h00000000} /* (29, 16, 11) {real, imag} */,
  {32'hc45eaf5c, 32'h00000000} /* (29, 16, 10) {real, imag} */,
  {32'hc5107169, 32'h00000000} /* (29, 16, 9) {real, imag} */,
  {32'hc58b941b, 32'h00000000} /* (29, 16, 8) {real, imag} */,
  {32'hc57e5c67, 32'h00000000} /* (29, 16, 7) {real, imag} */,
  {32'hc591c40a, 32'h00000000} /* (29, 16, 6) {real, imag} */,
  {32'hc586a7b3, 32'h00000000} /* (29, 16, 5) {real, imag} */,
  {32'hc58d3f89, 32'h00000000} /* (29, 16, 4) {real, imag} */,
  {32'hc598e15b, 32'h00000000} /* (29, 16, 3) {real, imag} */,
  {32'hc5831347, 32'h00000000} /* (29, 16, 2) {real, imag} */,
  {32'hc596a0df, 32'h00000000} /* (29, 16, 1) {real, imag} */,
  {32'hc5591296, 32'h00000000} /* (29, 16, 0) {real, imag} */,
  {32'hc55cab8d, 32'h00000000} /* (29, 15, 31) {real, imag} */,
  {32'hc5874f7c, 32'h00000000} /* (29, 15, 30) {real, imag} */,
  {32'hc57903ca, 32'h00000000} /* (29, 15, 29) {real, imag} */,
  {32'hc5712598, 32'h00000000} /* (29, 15, 28) {real, imag} */,
  {32'hc566f8b6, 32'h00000000} /* (29, 15, 27) {real, imag} */,
  {32'hc57633e6, 32'h00000000} /* (29, 15, 26) {real, imag} */,
  {32'hc58d8f4a, 32'h00000000} /* (29, 15, 25) {real, imag} */,
  {32'hc56e2b41, 32'h00000000} /* (29, 15, 24) {real, imag} */,
  {32'hc52c23f4, 32'h00000000} /* (29, 15, 23) {real, imag} */,
  {32'hc50341ad, 32'h00000000} /* (29, 15, 22) {real, imag} */,
  {32'hc40ae7bc, 32'h00000000} /* (29, 15, 21) {real, imag} */,
  {32'h44dae8a4, 32'h00000000} /* (29, 15, 20) {real, imag} */,
  {32'h44fa23fe, 32'h00000000} /* (29, 15, 19) {real, imag} */,
  {32'h4548433c, 32'h00000000} /* (29, 15, 18) {real, imag} */,
  {32'h453e41d2, 32'h00000000} /* (29, 15, 17) {real, imag} */,
  {32'h458ed82e, 32'h00000000} /* (29, 15, 16) {real, imag} */,
  {32'h45953b46, 32'h00000000} /* (29, 15, 15) {real, imag} */,
  {32'h458ae6e2, 32'h00000000} /* (29, 15, 14) {real, imag} */,
  {32'h455afcf6, 32'h00000000} /* (29, 15, 13) {real, imag} */,
  {32'h453d4b26, 32'h00000000} /* (29, 15, 12) {real, imag} */,
  {32'h444e5918, 32'h00000000} /* (29, 15, 11) {real, imag} */,
  {32'hc4e6c514, 32'h00000000} /* (29, 15, 10) {real, imag} */,
  {32'hc533eba5, 32'h00000000} /* (29, 15, 9) {real, imag} */,
  {32'hc578f50b, 32'h00000000} /* (29, 15, 8) {real, imag} */,
  {32'hc5bfedfa, 32'h00000000} /* (29, 15, 7) {real, imag} */,
  {32'hc58b698e, 32'h00000000} /* (29, 15, 6) {real, imag} */,
  {32'hc590c218, 32'h00000000} /* (29, 15, 5) {real, imag} */,
  {32'hc5803970, 32'h00000000} /* (29, 15, 4) {real, imag} */,
  {32'hc570ef17, 32'h00000000} /* (29, 15, 3) {real, imag} */,
  {32'hc57bd240, 32'h00000000} /* (29, 15, 2) {real, imag} */,
  {32'hc5646a0e, 32'h00000000} /* (29, 15, 1) {real, imag} */,
  {32'hc54a4c47, 32'h00000000} /* (29, 15, 0) {real, imag} */,
  {32'hc557c6d0, 32'h00000000} /* (29, 14, 31) {real, imag} */,
  {32'hc58ae58c, 32'h00000000} /* (29, 14, 30) {real, imag} */,
  {32'hc58fe40b, 32'h00000000} /* (29, 14, 29) {real, imag} */,
  {32'hc558332c, 32'h00000000} /* (29, 14, 28) {real, imag} */,
  {32'hc55e6afe, 32'h00000000} /* (29, 14, 27) {real, imag} */,
  {32'hc558dcc2, 32'h00000000} /* (29, 14, 26) {real, imag} */,
  {32'hc56abaee, 32'h00000000} /* (29, 14, 25) {real, imag} */,
  {32'hc5937768, 32'h00000000} /* (29, 14, 24) {real, imag} */,
  {32'hc568a988, 32'h00000000} /* (29, 14, 23) {real, imag} */,
  {32'hc54a0a22, 32'h00000000} /* (29, 14, 22) {real, imag} */,
  {32'hc4531b4c, 32'h00000000} /* (29, 14, 21) {real, imag} */,
  {32'h44c40df3, 32'h00000000} /* (29, 14, 20) {real, imag} */,
  {32'h45087bfb, 32'h00000000} /* (29, 14, 19) {real, imag} */,
  {32'h451e0df6, 32'h00000000} /* (29, 14, 18) {real, imag} */,
  {32'h45652d7a, 32'h00000000} /* (29, 14, 17) {real, imag} */,
  {32'h45842192, 32'h00000000} /* (29, 14, 16) {real, imag} */,
  {32'h457240f8, 32'h00000000} /* (29, 14, 15) {real, imag} */,
  {32'h458e4698, 32'h00000000} /* (29, 14, 14) {real, imag} */,
  {32'h452edfd9, 32'h00000000} /* (29, 14, 13) {real, imag} */,
  {32'h451cd262, 32'h00000000} /* (29, 14, 12) {real, imag} */,
  {32'h44d3e864, 32'h00000000} /* (29, 14, 11) {real, imag} */,
  {32'hc4728638, 32'h00000000} /* (29, 14, 10) {real, imag} */,
  {32'hc571bb2a, 32'h00000000} /* (29, 14, 9) {real, imag} */,
  {32'hc56bd60d, 32'h00000000} /* (29, 14, 8) {real, imag} */,
  {32'hc586b170, 32'h00000000} /* (29, 14, 7) {real, imag} */,
  {32'hc58444a7, 32'h00000000} /* (29, 14, 6) {real, imag} */,
  {32'hc5954218, 32'h00000000} /* (29, 14, 5) {real, imag} */,
  {32'hc55e1d96, 32'h00000000} /* (29, 14, 4) {real, imag} */,
  {32'hc591e04e, 32'h00000000} /* (29, 14, 3) {real, imag} */,
  {32'hc57fb2c4, 32'h00000000} /* (29, 14, 2) {real, imag} */,
  {32'hc53a1b92, 32'h00000000} /* (29, 14, 1) {real, imag} */,
  {32'hc55c1e33, 32'h00000000} /* (29, 14, 0) {real, imag} */,
  {32'hc55dfbb3, 32'h00000000} /* (29, 13, 31) {real, imag} */,
  {32'hc5644f3c, 32'h00000000} /* (29, 13, 30) {real, imag} */,
  {32'hc576181e, 32'h00000000} /* (29, 13, 29) {real, imag} */,
  {32'hc58cb54f, 32'h00000000} /* (29, 13, 28) {real, imag} */,
  {32'hc54c87fd, 32'h00000000} /* (29, 13, 27) {real, imag} */,
  {32'hc5561530, 32'h00000000} /* (29, 13, 26) {real, imag} */,
  {32'hc58b1fe2, 32'h00000000} /* (29, 13, 25) {real, imag} */,
  {32'hc5938d86, 32'h00000000} /* (29, 13, 24) {real, imag} */,
  {32'hc53b0e4c, 32'h00000000} /* (29, 13, 23) {real, imag} */,
  {32'hc54270d4, 32'h00000000} /* (29, 13, 22) {real, imag} */,
  {32'hc4aee69a, 32'h00000000} /* (29, 13, 21) {real, imag} */,
  {32'h44394a2a, 32'h00000000} /* (29, 13, 20) {real, imag} */,
  {32'h453cf044, 32'h00000000} /* (29, 13, 19) {real, imag} */,
  {32'h456222fa, 32'h00000000} /* (29, 13, 18) {real, imag} */,
  {32'h4543b37e, 32'h00000000} /* (29, 13, 17) {real, imag} */,
  {32'h456d6bf3, 32'h00000000} /* (29, 13, 16) {real, imag} */,
  {32'h45408761, 32'h00000000} /* (29, 13, 15) {real, imag} */,
  {32'h4523d990, 32'h00000000} /* (29, 13, 14) {real, imag} */,
  {32'h45317650, 32'h00000000} /* (29, 13, 13) {real, imag} */,
  {32'h45339ef0, 32'h00000000} /* (29, 13, 12) {real, imag} */,
  {32'h44ab2aba, 32'h00000000} /* (29, 13, 11) {real, imag} */,
  {32'hc4dc92d1, 32'h00000000} /* (29, 13, 10) {real, imag} */,
  {32'hc52d8fe9, 32'h00000000} /* (29, 13, 9) {real, imag} */,
  {32'hc58fc062, 32'h00000000} /* (29, 13, 8) {real, imag} */,
  {32'hc5578d72, 32'h00000000} /* (29, 13, 7) {real, imag} */,
  {32'hc551726e, 32'h00000000} /* (29, 13, 6) {real, imag} */,
  {32'hc5741ef5, 32'h00000000} /* (29, 13, 5) {real, imag} */,
  {32'hc57291d8, 32'h00000000} /* (29, 13, 4) {real, imag} */,
  {32'hc5916756, 32'h00000000} /* (29, 13, 3) {real, imag} */,
  {32'hc56e2c22, 32'h00000000} /* (29, 13, 2) {real, imag} */,
  {32'hc54d287c, 32'h00000000} /* (29, 13, 1) {real, imag} */,
  {32'hc53683db, 32'h00000000} /* (29, 13, 0) {real, imag} */,
  {32'hc50e68e4, 32'h00000000} /* (29, 12, 31) {real, imag} */,
  {32'hc516dce8, 32'h00000000} /* (29, 12, 30) {real, imag} */,
  {32'hc510c18a, 32'h00000000} /* (29, 12, 29) {real, imag} */,
  {32'hc56632a2, 32'h00000000} /* (29, 12, 28) {real, imag} */,
  {32'hc592a1ee, 32'h00000000} /* (29, 12, 27) {real, imag} */,
  {32'hc531bb0a, 32'h00000000} /* (29, 12, 26) {real, imag} */,
  {32'hc5496044, 32'h00000000} /* (29, 12, 25) {real, imag} */,
  {32'hc5530771, 32'h00000000} /* (29, 12, 24) {real, imag} */,
  {32'hc5035c20, 32'h00000000} /* (29, 12, 23) {real, imag} */,
  {32'hc4e4902c, 32'h00000000} /* (29, 12, 22) {real, imag} */,
  {32'hc4a9757e, 32'h00000000} /* (29, 12, 21) {real, imag} */,
  {32'h44806440, 32'h00000000} /* (29, 12, 20) {real, imag} */,
  {32'h45760250, 32'h00000000} /* (29, 12, 19) {real, imag} */,
  {32'h4546e493, 32'h00000000} /* (29, 12, 18) {real, imag} */,
  {32'h452bbbcc, 32'h00000000} /* (29, 12, 17) {real, imag} */,
  {32'h45431e8e, 32'h00000000} /* (29, 12, 16) {real, imag} */,
  {32'h45063f08, 32'h00000000} /* (29, 12, 15) {real, imag} */,
  {32'h451bc606, 32'h00000000} /* (29, 12, 14) {real, imag} */,
  {32'h45053fe8, 32'h00000000} /* (29, 12, 13) {real, imag} */,
  {32'h44ee3d61, 32'h00000000} /* (29, 12, 12) {real, imag} */,
  {32'h44bedc36, 32'h00000000} /* (29, 12, 11) {real, imag} */,
  {32'hc4255f56, 32'h00000000} /* (29, 12, 10) {real, imag} */,
  {32'hc511ad92, 32'h00000000} /* (29, 12, 9) {real, imag} */,
  {32'hc55fc2f9, 32'h00000000} /* (29, 12, 8) {real, imag} */,
  {32'hc5338be6, 32'h00000000} /* (29, 12, 7) {real, imag} */,
  {32'hc531d66e, 32'h00000000} /* (29, 12, 6) {real, imag} */,
  {32'hc54d0439, 32'h00000000} /* (29, 12, 5) {real, imag} */,
  {32'hc520489c, 32'h00000000} /* (29, 12, 4) {real, imag} */,
  {32'hc51fd3a8, 32'h00000000} /* (29, 12, 3) {real, imag} */,
  {32'hc586007c, 32'h00000000} /* (29, 12, 2) {real, imag} */,
  {32'hc59679d0, 32'h00000000} /* (29, 12, 1) {real, imag} */,
  {32'hc5236a2c, 32'h00000000} /* (29, 12, 0) {real, imag} */,
  {32'hc47885a7, 32'h00000000} /* (29, 11, 31) {real, imag} */,
  {32'hc4b155ca, 32'h00000000} /* (29, 11, 30) {real, imag} */,
  {32'hc4b281aa, 32'h00000000} /* (29, 11, 29) {real, imag} */,
  {32'hc50495c0, 32'h00000000} /* (29, 11, 28) {real, imag} */,
  {32'hc553eaaa, 32'h00000000} /* (29, 11, 27) {real, imag} */,
  {32'hc51492e2, 32'h00000000} /* (29, 11, 26) {real, imag} */,
  {32'hc4d020ae, 32'h00000000} /* (29, 11, 25) {real, imag} */,
  {32'hc4aea34c, 32'h00000000} /* (29, 11, 24) {real, imag} */,
  {32'hc4ac4a2b, 32'h00000000} /* (29, 11, 23) {real, imag} */,
  {32'hc46a9990, 32'h00000000} /* (29, 11, 22) {real, imag} */,
  {32'hc4d0cb9e, 32'h00000000} /* (29, 11, 21) {real, imag} */,
  {32'hc37808f2, 32'h00000000} /* (29, 11, 20) {real, imag} */,
  {32'h449ff040, 32'h00000000} /* (29, 11, 19) {real, imag} */,
  {32'h45170a9e, 32'h00000000} /* (29, 11, 18) {real, imag} */,
  {32'h450afb20, 32'h00000000} /* (29, 11, 17) {real, imag} */,
  {32'h44b9455a, 32'h00000000} /* (29, 11, 16) {real, imag} */,
  {32'h448ca766, 32'h00000000} /* (29, 11, 15) {real, imag} */,
  {32'h44583f10, 32'h00000000} /* (29, 11, 14) {real, imag} */,
  {32'h44c2f772, 32'h00000000} /* (29, 11, 13) {real, imag} */,
  {32'h43b84358, 32'h00000000} /* (29, 11, 12) {real, imag} */,
  {32'hc3071dd8, 32'h00000000} /* (29, 11, 11) {real, imag} */,
  {32'hc43932bf, 32'h00000000} /* (29, 11, 10) {real, imag} */,
  {32'hc4fb887e, 32'h00000000} /* (29, 11, 9) {real, imag} */,
  {32'hc485d880, 32'h00000000} /* (29, 11, 8) {real, imag} */,
  {32'hc511dee2, 32'h00000000} /* (29, 11, 7) {real, imag} */,
  {32'hc4f351bc, 32'h00000000} /* (29, 11, 6) {real, imag} */,
  {32'hc467a6bf, 32'h00000000} /* (29, 11, 5) {real, imag} */,
  {32'hc486b85c, 32'h00000000} /* (29, 11, 4) {real, imag} */,
  {32'hc52e3c28, 32'h00000000} /* (29, 11, 3) {real, imag} */,
  {32'hc53d5e16, 32'h00000000} /* (29, 11, 2) {real, imag} */,
  {32'hc525c03e, 32'h00000000} /* (29, 11, 1) {real, imag} */,
  {32'hc4fba130, 32'h00000000} /* (29, 11, 0) {real, imag} */,
  {32'h4434ea92, 32'h00000000} /* (29, 10, 31) {real, imag} */,
  {32'h446c5571, 32'h00000000} /* (29, 10, 30) {real, imag} */,
  {32'h44817d74, 32'h00000000} /* (29, 10, 29) {real, imag} */,
  {32'h44508bd5, 32'h00000000} /* (29, 10, 28) {real, imag} */,
  {32'h4506e308, 32'h00000000} /* (29, 10, 27) {real, imag} */,
  {32'hc1b5f4a0, 32'h00000000} /* (29, 10, 26) {real, imag} */,
  {32'h4457f45a, 32'h00000000} /* (29, 10, 25) {real, imag} */,
  {32'h44549e27, 32'h00000000} /* (29, 10, 24) {real, imag} */,
  {32'h4330f290, 32'h00000000} /* (29, 10, 23) {real, imag} */,
  {32'h432b1bae, 32'h00000000} /* (29, 10, 22) {real, imag} */,
  {32'hc41e1113, 32'h00000000} /* (29, 10, 21) {real, imag} */,
  {32'hc4e6fa09, 32'h00000000} /* (29, 10, 20) {real, imag} */,
  {32'hc46157bc, 32'h00000000} /* (29, 10, 19) {real, imag} */,
  {32'hc42b674d, 32'h00000000} /* (29, 10, 18) {real, imag} */,
  {32'hc4dd4597, 32'h00000000} /* (29, 10, 17) {real, imag} */,
  {32'hc3e61ca0, 32'h00000000} /* (29, 10, 16) {real, imag} */,
  {32'hc42cb59c, 32'h00000000} /* (29, 10, 15) {real, imag} */,
  {32'hc45d1bc7, 32'h00000000} /* (29, 10, 14) {real, imag} */,
  {32'hc4372697, 32'h00000000} /* (29, 10, 13) {real, imag} */,
  {32'hc4f3cfb0, 32'h00000000} /* (29, 10, 12) {real, imag} */,
  {32'hc42cef9a, 32'h00000000} /* (29, 10, 11) {real, imag} */,
  {32'hc40f284f, 32'h00000000} /* (29, 10, 10) {real, imag} */,
  {32'hc3f810e0, 32'h00000000} /* (29, 10, 9) {real, imag} */,
  {32'hc3c341ca, 32'h00000000} /* (29, 10, 8) {real, imag} */,
  {32'h42ca9074, 32'h00000000} /* (29, 10, 7) {real, imag} */,
  {32'h442a0ff2, 32'h00000000} /* (29, 10, 6) {real, imag} */,
  {32'h448ea03c, 32'h00000000} /* (29, 10, 5) {real, imag} */,
  {32'h44cb26a1, 32'h00000000} /* (29, 10, 4) {real, imag} */,
  {32'h440b8bd8, 32'h00000000} /* (29, 10, 3) {real, imag} */,
  {32'h448327c0, 32'h00000000} /* (29, 10, 2) {real, imag} */,
  {32'h4472000e, 32'h00000000} /* (29, 10, 1) {real, imag} */,
  {32'h44a19e8b, 32'h00000000} /* (29, 10, 0) {real, imag} */,
  {32'h44f7b4ec, 32'h00000000} /* (29, 9, 31) {real, imag} */,
  {32'h452e545e, 32'h00000000} /* (29, 9, 30) {real, imag} */,
  {32'h456adcc2, 32'h00000000} /* (29, 9, 29) {real, imag} */,
  {32'h45427540, 32'h00000000} /* (29, 9, 28) {real, imag} */,
  {32'h44fc7ec5, 32'h00000000} /* (29, 9, 27) {real, imag} */,
  {32'h44f1fb55, 32'h00000000} /* (29, 9, 26) {real, imag} */,
  {32'h44ddceba, 32'h00000000} /* (29, 9, 25) {real, imag} */,
  {32'h45050b7e, 32'h00000000} /* (29, 9, 24) {real, imag} */,
  {32'h4500ba8f, 32'h00000000} /* (29, 9, 23) {real, imag} */,
  {32'h44ca7fa4, 32'h00000000} /* (29, 9, 22) {real, imag} */,
  {32'hc4035e00, 32'h00000000} /* (29, 9, 21) {real, imag} */,
  {32'hc4d7c78e, 32'h00000000} /* (29, 9, 20) {real, imag} */,
  {32'hc4d126e8, 32'h00000000} /* (29, 9, 19) {real, imag} */,
  {32'hc507d4fd, 32'h00000000} /* (29, 9, 18) {real, imag} */,
  {32'hc51ac8b9, 32'h00000000} /* (29, 9, 17) {real, imag} */,
  {32'hc5286a84, 32'h00000000} /* (29, 9, 16) {real, imag} */,
  {32'hc5625df0, 32'h00000000} /* (29, 9, 15) {real, imag} */,
  {32'hc517ba32, 32'h00000000} /* (29, 9, 14) {real, imag} */,
  {32'hc518258a, 32'h00000000} /* (29, 9, 13) {real, imag} */,
  {32'hc56f6978, 32'h00000000} /* (29, 9, 12) {real, imag} */,
  {32'hc506c681, 32'h00000000} /* (29, 9, 11) {real, imag} */,
  {32'hc353a978, 32'h00000000} /* (29, 9, 10) {real, imag} */,
  {32'h43ad3c18, 32'h00000000} /* (29, 9, 9) {real, imag} */,
  {32'h442dfe76, 32'h00000000} /* (29, 9, 8) {real, imag} */,
  {32'h450b2b67, 32'h00000000} /* (29, 9, 7) {real, imag} */,
  {32'h44f140f2, 32'h00000000} /* (29, 9, 6) {real, imag} */,
  {32'h45159a60, 32'h00000000} /* (29, 9, 5) {real, imag} */,
  {32'h454982f9, 32'h00000000} /* (29, 9, 4) {real, imag} */,
  {32'h455c59a2, 32'h00000000} /* (29, 9, 3) {real, imag} */,
  {32'h4503e8d3, 32'h00000000} /* (29, 9, 2) {real, imag} */,
  {32'h4500ca57, 32'h00000000} /* (29, 9, 1) {real, imag} */,
  {32'h450ff780, 32'h00000000} /* (29, 9, 0) {real, imag} */,
  {32'h4527c8be, 32'h00000000} /* (29, 8, 31) {real, imag} */,
  {32'h45618529, 32'h00000000} /* (29, 8, 30) {real, imag} */,
  {32'h454ccd6c, 32'h00000000} /* (29, 8, 29) {real, imag} */,
  {32'h44e0d131, 32'h00000000} /* (29, 8, 28) {real, imag} */,
  {32'h4507c9f4, 32'h00000000} /* (29, 8, 27) {real, imag} */,
  {32'h4513315a, 32'h00000000} /* (29, 8, 26) {real, imag} */,
  {32'h44fa718a, 32'h00000000} /* (29, 8, 25) {real, imag} */,
  {32'h44e5ba68, 32'h00000000} /* (29, 8, 24) {real, imag} */,
  {32'h452db14e, 32'h00000000} /* (29, 8, 23) {real, imag} */,
  {32'h4511def0, 32'h00000000} /* (29, 8, 22) {real, imag} */,
  {32'h4469f6ad, 32'h00000000} /* (29, 8, 21) {real, imag} */,
  {32'hc4972a4b, 32'h00000000} /* (29, 8, 20) {real, imag} */,
  {32'hc514b40c, 32'h00000000} /* (29, 8, 19) {real, imag} */,
  {32'hc517209a, 32'h00000000} /* (29, 8, 18) {real, imag} */,
  {32'hc52157db, 32'h00000000} /* (29, 8, 17) {real, imag} */,
  {32'hc52487a8, 32'h00000000} /* (29, 8, 16) {real, imag} */,
  {32'hc53bdd9c, 32'h00000000} /* (29, 8, 15) {real, imag} */,
  {32'hc58e6cee, 32'h00000000} /* (29, 8, 14) {real, imag} */,
  {32'hc56829fe, 32'h00000000} /* (29, 8, 13) {real, imag} */,
  {32'hc53d2f34, 32'h00000000} /* (29, 8, 12) {real, imag} */,
  {32'hc52f2dbc, 32'h00000000} /* (29, 8, 11) {real, imag} */,
  {32'hc43996b4, 32'h00000000} /* (29, 8, 10) {real, imag} */,
  {32'h441f1a04, 32'h00000000} /* (29, 8, 9) {real, imag} */,
  {32'h44cffad8, 32'h00000000} /* (29, 8, 8) {real, imag} */,
  {32'h44ba0c18, 32'h00000000} /* (29, 8, 7) {real, imag} */,
  {32'h452c761a, 32'h00000000} /* (29, 8, 6) {real, imag} */,
  {32'h452ef7f3, 32'h00000000} /* (29, 8, 5) {real, imag} */,
  {32'h45851d29, 32'h00000000} /* (29, 8, 4) {real, imag} */,
  {32'h4573af86, 32'h00000000} /* (29, 8, 3) {real, imag} */,
  {32'h45579eca, 32'h00000000} /* (29, 8, 2) {real, imag} */,
  {32'h456516b7, 32'h00000000} /* (29, 8, 1) {real, imag} */,
  {32'h450fcd80, 32'h00000000} /* (29, 8, 0) {real, imag} */,
  {32'h4505b2b8, 32'h00000000} /* (29, 7, 31) {real, imag} */,
  {32'h45511598, 32'h00000000} /* (29, 7, 30) {real, imag} */,
  {32'h45257dba, 32'h00000000} /* (29, 7, 29) {real, imag} */,
  {32'h45002732, 32'h00000000} /* (29, 7, 28) {real, imag} */,
  {32'h45134c1a, 32'h00000000} /* (29, 7, 27) {real, imag} */,
  {32'h45375c12, 32'h00000000} /* (29, 7, 26) {real, imag} */,
  {32'h45313ff5, 32'h00000000} /* (29, 7, 25) {real, imag} */,
  {32'h452145da, 32'h00000000} /* (29, 7, 24) {real, imag} */,
  {32'h452a7c07, 32'h00000000} /* (29, 7, 23) {real, imag} */,
  {32'h44f01ea0, 32'h00000000} /* (29, 7, 22) {real, imag} */,
  {32'h44a9d734, 32'h00000000} /* (29, 7, 21) {real, imag} */,
  {32'hc2d330b0, 32'h00000000} /* (29, 7, 20) {real, imag} */,
  {32'hc53d18de, 32'h00000000} /* (29, 7, 19) {real, imag} */,
  {32'hc540d2ee, 32'h00000000} /* (29, 7, 18) {real, imag} */,
  {32'hc538651a, 32'h00000000} /* (29, 7, 17) {real, imag} */,
  {32'hc5508e87, 32'h00000000} /* (29, 7, 16) {real, imag} */,
  {32'hc527991c, 32'h00000000} /* (29, 7, 15) {real, imag} */,
  {32'hc582cf72, 32'h00000000} /* (29, 7, 14) {real, imag} */,
  {32'hc57ca0ee, 32'h00000000} /* (29, 7, 13) {real, imag} */,
  {32'hc52fda42, 32'h00000000} /* (29, 7, 12) {real, imag} */,
  {32'hc4fa7a9b, 32'h00000000} /* (29, 7, 11) {real, imag} */,
  {32'hc3e2a654, 32'h00000000} /* (29, 7, 10) {real, imag} */,
  {32'h443f7ff4, 32'h00000000} /* (29, 7, 9) {real, imag} */,
  {32'h45049c1c, 32'h00000000} /* (29, 7, 8) {real, imag} */,
  {32'h449f4abc, 32'h00000000} /* (29, 7, 7) {real, imag} */,
  {32'h45161d94, 32'h00000000} /* (29, 7, 6) {real, imag} */,
  {32'h455da198, 32'h00000000} /* (29, 7, 5) {real, imag} */,
  {32'h456ca3a4, 32'h00000000} /* (29, 7, 4) {real, imag} */,
  {32'h4584afa3, 32'h00000000} /* (29, 7, 3) {real, imag} */,
  {32'h45857702, 32'h00000000} /* (29, 7, 2) {real, imag} */,
  {32'h4538ef58, 32'h00000000} /* (29, 7, 1) {real, imag} */,
  {32'h45088d6f, 32'h00000000} /* (29, 7, 0) {real, imag} */,
  {32'h4524ff36, 32'h00000000} /* (29, 6, 31) {real, imag} */,
  {32'h45400566, 32'h00000000} /* (29, 6, 30) {real, imag} */,
  {32'h4545c5d0, 32'h00000000} /* (29, 6, 29) {real, imag} */,
  {32'h450c9f1c, 32'h00000000} /* (29, 6, 28) {real, imag} */,
  {32'h4518462b, 32'h00000000} /* (29, 6, 27) {real, imag} */,
  {32'h453114c0, 32'h00000000} /* (29, 6, 26) {real, imag} */,
  {32'h452fa0f7, 32'h00000000} /* (29, 6, 25) {real, imag} */,
  {32'h45348047, 32'h00000000} /* (29, 6, 24) {real, imag} */,
  {32'h453a52dc, 32'h00000000} /* (29, 6, 23) {real, imag} */,
  {32'h44fcc657, 32'h00000000} /* (29, 6, 22) {real, imag} */,
  {32'h44c97bec, 32'h00000000} /* (29, 6, 21) {real, imag} */,
  {32'h42945430, 32'h00000000} /* (29, 6, 20) {real, imag} */,
  {32'hc44081b0, 32'h00000000} /* (29, 6, 19) {real, imag} */,
  {32'hc4edfd4c, 32'h00000000} /* (29, 6, 18) {real, imag} */,
  {32'hc50a9c91, 32'h00000000} /* (29, 6, 17) {real, imag} */,
  {32'hc56a55ee, 32'h00000000} /* (29, 6, 16) {real, imag} */,
  {32'hc582939b, 32'h00000000} /* (29, 6, 15) {real, imag} */,
  {32'hc55d2d2a, 32'h00000000} /* (29, 6, 14) {real, imag} */,
  {32'hc569e4c2, 32'h00000000} /* (29, 6, 13) {real, imag} */,
  {32'hc567a938, 32'h00000000} /* (29, 6, 12) {real, imag} */,
  {32'hc54f6c15, 32'h00000000} /* (29, 6, 11) {real, imag} */,
  {32'hc483530c, 32'h00000000} /* (29, 6, 10) {real, imag} */,
  {32'h43cb9d68, 32'h00000000} /* (29, 6, 9) {real, imag} */,
  {32'h439227d0, 32'h00000000} /* (29, 6, 8) {real, imag} */,
  {32'h44a9e91c, 32'h00000000} /* (29, 6, 7) {real, imag} */,
  {32'h44ed171d, 32'h00000000} /* (29, 6, 6) {real, imag} */,
  {32'h45636d70, 32'h00000000} /* (29, 6, 5) {real, imag} */,
  {32'h456c5d38, 32'h00000000} /* (29, 6, 4) {real, imag} */,
  {32'h4545d6ec, 32'h00000000} /* (29, 6, 3) {real, imag} */,
  {32'h455b5716, 32'h00000000} /* (29, 6, 2) {real, imag} */,
  {32'h455187ed, 32'h00000000} /* (29, 6, 1) {real, imag} */,
  {32'h450c81ac, 32'h00000000} /* (29, 6, 0) {real, imag} */,
  {32'h450797c4, 32'h00000000} /* (29, 5, 31) {real, imag} */,
  {32'h45449dd4, 32'h00000000} /* (29, 5, 30) {real, imag} */,
  {32'h4557f324, 32'h00000000} /* (29, 5, 29) {real, imag} */,
  {32'h45254d50, 32'h00000000} /* (29, 5, 28) {real, imag} */,
  {32'h452059b0, 32'h00000000} /* (29, 5, 27) {real, imag} */,
  {32'h45360391, 32'h00000000} /* (29, 5, 26) {real, imag} */,
  {32'h453fe9fc, 32'h00000000} /* (29, 5, 25) {real, imag} */,
  {32'h453e9e5c, 32'h00000000} /* (29, 5, 24) {real, imag} */,
  {32'h453b3578, 32'h00000000} /* (29, 5, 23) {real, imag} */,
  {32'h4562b283, 32'h00000000} /* (29, 5, 22) {real, imag} */,
  {32'h457db4eb, 32'h00000000} /* (29, 5, 21) {real, imag} */,
  {32'h450d97e7, 32'h00000000} /* (29, 5, 20) {real, imag} */,
  {32'h44a0267f, 32'h00000000} /* (29, 5, 19) {real, imag} */,
  {32'hc38f3068, 32'h00000000} /* (29, 5, 18) {real, imag} */,
  {32'hc345de18, 32'h00000000} /* (29, 5, 17) {real, imag} */,
  {32'hc4a6a01b, 32'h00000000} /* (29, 5, 16) {real, imag} */,
  {32'hc54d1278, 32'h00000000} /* (29, 5, 15) {real, imag} */,
  {32'hc5504538, 32'h00000000} /* (29, 5, 14) {real, imag} */,
  {32'hc57fa7f8, 32'h00000000} /* (29, 5, 13) {real, imag} */,
  {32'hc581959f, 32'h00000000} /* (29, 5, 12) {real, imag} */,
  {32'hc59c1b50, 32'h00000000} /* (29, 5, 11) {real, imag} */,
  {32'hc5122e1b, 32'h00000000} /* (29, 5, 10) {real, imag} */,
  {32'hc4ed6638, 32'h00000000} /* (29, 5, 9) {real, imag} */,
  {32'hc4123056, 32'h00000000} /* (29, 5, 8) {real, imag} */,
  {32'h437f1468, 32'h00000000} /* (29, 5, 7) {real, imag} */,
  {32'h441972e4, 32'h00000000} /* (29, 5, 6) {real, imag} */,
  {32'h4507d3c9, 32'h00000000} /* (29, 5, 5) {real, imag} */,
  {32'h45802afc, 32'h00000000} /* (29, 5, 4) {real, imag} */,
  {32'h454fc448, 32'h00000000} /* (29, 5, 3) {real, imag} */,
  {32'h454812f3, 32'h00000000} /* (29, 5, 2) {real, imag} */,
  {32'h4559a81a, 32'h00000000} /* (29, 5, 1) {real, imag} */,
  {32'h45290c72, 32'h00000000} /* (29, 5, 0) {real, imag} */,
  {32'h44f87c01, 32'h00000000} /* (29, 4, 31) {real, imag} */,
  {32'h44eaef7c, 32'h00000000} /* (29, 4, 30) {real, imag} */,
  {32'h45245fa6, 32'h00000000} /* (29, 4, 29) {real, imag} */,
  {32'h453ca519, 32'h00000000} /* (29, 4, 28) {real, imag} */,
  {32'h45302fd6, 32'h00000000} /* (29, 4, 27) {real, imag} */,
  {32'h452a8998, 32'h00000000} /* (29, 4, 26) {real, imag} */,
  {32'h4526d2de, 32'h00000000} /* (29, 4, 25) {real, imag} */,
  {32'h451cf110, 32'h00000000} /* (29, 4, 24) {real, imag} */,
  {32'h453afee8, 32'h00000000} /* (29, 4, 23) {real, imag} */,
  {32'h4529c604, 32'h00000000} /* (29, 4, 22) {real, imag} */,
  {32'h456ff0cb, 32'h00000000} /* (29, 4, 21) {real, imag} */,
  {32'h4590bfa6, 32'h00000000} /* (29, 4, 20) {real, imag} */,
  {32'h451ce3bc, 32'h00000000} /* (29, 4, 19) {real, imag} */,
  {32'h45154640, 32'h00000000} /* (29, 4, 18) {real, imag} */,
  {32'h449f13f9, 32'h00000000} /* (29, 4, 17) {real, imag} */,
  {32'hc3cf14c8, 32'h00000000} /* (29, 4, 16) {real, imag} */,
  {32'hc52d62ea, 32'h00000000} /* (29, 4, 15) {real, imag} */,
  {32'hc55dda98, 32'h00000000} /* (29, 4, 14) {real, imag} */,
  {32'hc55fe63e, 32'h00000000} /* (29, 4, 13) {real, imag} */,
  {32'hc564f323, 32'h00000000} /* (29, 4, 12) {real, imag} */,
  {32'hc582a879, 32'h00000000} /* (29, 4, 11) {real, imag} */,
  {32'hc581ea3c, 32'h00000000} /* (29, 4, 10) {real, imag} */,
  {32'hc5191ca2, 32'h00000000} /* (29, 4, 9) {real, imag} */,
  {32'hc4da5f37, 32'h00000000} /* (29, 4, 8) {real, imag} */,
  {32'hc4d0362f, 32'h00000000} /* (29, 4, 7) {real, imag} */,
  {32'hc3ef5b84, 32'h00000000} /* (29, 4, 6) {real, imag} */,
  {32'h44ad83da, 32'h00000000} /* (29, 4, 5) {real, imag} */,
  {32'h454f7a63, 32'h00000000} /* (29, 4, 4) {real, imag} */,
  {32'h45310de4, 32'h00000000} /* (29, 4, 3) {real, imag} */,
  {32'h45596390, 32'h00000000} /* (29, 4, 2) {real, imag} */,
  {32'h45177cd8, 32'h00000000} /* (29, 4, 1) {real, imag} */,
  {32'h4500192f, 32'h00000000} /* (29, 4, 0) {real, imag} */,
  {32'h44a6a58c, 32'h00000000} /* (29, 3, 31) {real, imag} */,
  {32'h44fcc5ef, 32'h00000000} /* (29, 3, 30) {real, imag} */,
  {32'h4524d87b, 32'h00000000} /* (29, 3, 29) {real, imag} */,
  {32'h4503e013, 32'h00000000} /* (29, 3, 28) {real, imag} */,
  {32'h45271846, 32'h00000000} /* (29, 3, 27) {real, imag} */,
  {32'h45194cfa, 32'h00000000} /* (29, 3, 26) {real, imag} */,
  {32'h450231cb, 32'h00000000} /* (29, 3, 25) {real, imag} */,
  {32'h45196339, 32'h00000000} /* (29, 3, 24) {real, imag} */,
  {32'h45104b15, 32'h00000000} /* (29, 3, 23) {real, imag} */,
  {32'h451db402, 32'h00000000} /* (29, 3, 22) {real, imag} */,
  {32'h45392ffe, 32'h00000000} /* (29, 3, 21) {real, imag} */,
  {32'h4553c862, 32'h00000000} /* (29, 3, 20) {real, imag} */,
  {32'h45263ec6, 32'h00000000} /* (29, 3, 19) {real, imag} */,
  {32'h453e29aa, 32'h00000000} /* (29, 3, 18) {real, imag} */,
  {32'h4500453c, 32'h00000000} /* (29, 3, 17) {real, imag} */,
  {32'hc0f02a80, 32'h00000000} /* (29, 3, 16) {real, imag} */,
  {32'hc4b78690, 32'h00000000} /* (29, 3, 15) {real, imag} */,
  {32'hc5533b90, 32'h00000000} /* (29, 3, 14) {real, imag} */,
  {32'hc555d6ad, 32'h00000000} /* (29, 3, 13) {real, imag} */,
  {32'hc549b319, 32'h00000000} /* (29, 3, 12) {real, imag} */,
  {32'hc5847947, 32'h00000000} /* (29, 3, 11) {real, imag} */,
  {32'hc5752176, 32'h00000000} /* (29, 3, 10) {real, imag} */,
  {32'hc53e88df, 32'h00000000} /* (29, 3, 9) {real, imag} */,
  {32'hc52a211b, 32'h00000000} /* (29, 3, 8) {real, imag} */,
  {32'hc4fbb1e6, 32'h00000000} /* (29, 3, 7) {real, imag} */,
  {32'hc4c43478, 32'h00000000} /* (29, 3, 6) {real, imag} */,
  {32'hc1b43a00, 32'h00000000} /* (29, 3, 5) {real, imag} */,
  {32'h44d03f9b, 32'h00000000} /* (29, 3, 4) {real, imag} */,
  {32'h451159be, 32'h00000000} /* (29, 3, 3) {real, imag} */,
  {32'h450dea56, 32'h00000000} /* (29, 3, 2) {real, imag} */,
  {32'h44b43778, 32'h00000000} /* (29, 3, 1) {real, imag} */,
  {32'h44dc6704, 32'h00000000} /* (29, 3, 0) {real, imag} */,
  {32'h4509584e, 32'h00000000} /* (29, 2, 31) {real, imag} */,
  {32'h4548b3a7, 32'h00000000} /* (29, 2, 30) {real, imag} */,
  {32'h452b4bab, 32'h00000000} /* (29, 2, 29) {real, imag} */,
  {32'h4526c5e6, 32'h00000000} /* (29, 2, 28) {real, imag} */,
  {32'h4506a36a, 32'h00000000} /* (29, 2, 27) {real, imag} */,
  {32'h45105f6f, 32'h00000000} /* (29, 2, 26) {real, imag} */,
  {32'h4531d75c, 32'h00000000} /* (29, 2, 25) {real, imag} */,
  {32'h451bbc89, 32'h00000000} /* (29, 2, 24) {real, imag} */,
  {32'h4529c7c8, 32'h00000000} /* (29, 2, 23) {real, imag} */,
  {32'h45732368, 32'h00000000} /* (29, 2, 22) {real, imag} */,
  {32'h45644f0e, 32'h00000000} /* (29, 2, 21) {real, imag} */,
  {32'h453695c0, 32'h00000000} /* (29, 2, 20) {real, imag} */,
  {32'h4512c36c, 32'h00000000} /* (29, 2, 19) {real, imag} */,
  {32'h451a4d11, 32'h00000000} /* (29, 2, 18) {real, imag} */,
  {32'h45257c59, 32'h00000000} /* (29, 2, 17) {real, imag} */,
  {32'hc20a0740, 32'h00000000} /* (29, 2, 16) {real, imag} */,
  {32'hc48358fd, 32'h00000000} /* (29, 2, 15) {real, imag} */,
  {32'hc5214f11, 32'h00000000} /* (29, 2, 14) {real, imag} */,
  {32'hc5456d0d, 32'h00000000} /* (29, 2, 13) {real, imag} */,
  {32'hc54eb9be, 32'h00000000} /* (29, 2, 12) {real, imag} */,
  {32'hc56f483a, 32'h00000000} /* (29, 2, 11) {real, imag} */,
  {32'hc583dde3, 32'h00000000} /* (29, 2, 10) {real, imag} */,
  {32'hc565ab7c, 32'h00000000} /* (29, 2, 9) {real, imag} */,
  {32'hc52f818b, 32'h00000000} /* (29, 2, 8) {real, imag} */,
  {32'hc50fe256, 32'h00000000} /* (29, 2, 7) {real, imag} */,
  {32'hc513bbac, 32'h00000000} /* (29, 2, 6) {real, imag} */,
  {32'hc43c4c28, 32'h00000000} /* (29, 2, 5) {real, imag} */,
  {32'h44cc163c, 32'h00000000} /* (29, 2, 4) {real, imag} */,
  {32'h44ce2cc3, 32'h00000000} /* (29, 2, 3) {real, imag} */,
  {32'h448ec65a, 32'h00000000} /* (29, 2, 2) {real, imag} */,
  {32'h44d25fc9, 32'h00000000} /* (29, 2, 1) {real, imag} */,
  {32'h44c7823a, 32'h00000000} /* (29, 2, 0) {real, imag} */,
  {32'h44cd4cd0, 32'h00000000} /* (29, 1, 31) {real, imag} */,
  {32'h44d7f2b2, 32'h00000000} /* (29, 1, 30) {real, imag} */,
  {32'h44d5965e, 32'h00000000} /* (29, 1, 29) {real, imag} */,
  {32'h4529ed3c, 32'h00000000} /* (29, 1, 28) {real, imag} */,
  {32'h451233a6, 32'h00000000} /* (29, 1, 27) {real, imag} */,
  {32'h45246524, 32'h00000000} /* (29, 1, 26) {real, imag} */,
  {32'h452b932a, 32'h00000000} /* (29, 1, 25) {real, imag} */,
  {32'h4555bd22, 32'h00000000} /* (29, 1, 24) {real, imag} */,
  {32'h4554e1a4, 32'h00000000} /* (29, 1, 23) {real, imag} */,
  {32'h4554f04b, 32'h00000000} /* (29, 1, 22) {real, imag} */,
  {32'h455d6d07, 32'h00000000} /* (29, 1, 21) {real, imag} */,
  {32'h454ebf17, 32'h00000000} /* (29, 1, 20) {real, imag} */,
  {32'h4518df9b, 32'h00000000} /* (29, 1, 19) {real, imag} */,
  {32'h451d55e7, 32'h00000000} /* (29, 1, 18) {real, imag} */,
  {32'h450af91f, 32'h00000000} /* (29, 1, 17) {real, imag} */,
  {32'h4383b4c4, 32'h00000000} /* (29, 1, 16) {real, imag} */,
  {32'hc4d86bd4, 32'h00000000} /* (29, 1, 15) {real, imag} */,
  {32'hc54b0321, 32'h00000000} /* (29, 1, 14) {real, imag} */,
  {32'hc557b5a3, 32'h00000000} /* (29, 1, 13) {real, imag} */,
  {32'hc58dd0f4, 32'h00000000} /* (29, 1, 12) {real, imag} */,
  {32'hc5935216, 32'h00000000} /* (29, 1, 11) {real, imag} */,
  {32'hc53bbdac, 32'h00000000} /* (29, 1, 10) {real, imag} */,
  {32'hc53eedf2, 32'h00000000} /* (29, 1, 9) {real, imag} */,
  {32'hc51fb844, 32'h00000000} /* (29, 1, 8) {real, imag} */,
  {32'hc4fdd95b, 32'h00000000} /* (29, 1, 7) {real, imag} */,
  {32'hc4d0491e, 32'h00000000} /* (29, 1, 6) {real, imag} */,
  {32'hc33f6a70, 32'h00000000} /* (29, 1, 5) {real, imag} */,
  {32'h44c83c76, 32'h00000000} /* (29, 1, 4) {real, imag} */,
  {32'h4528f1f1, 32'h00000000} /* (29, 1, 3) {real, imag} */,
  {32'h4512a161, 32'h00000000} /* (29, 1, 2) {real, imag} */,
  {32'h44cd5124, 32'h00000000} /* (29, 1, 1) {real, imag} */,
  {32'h449b241b, 32'h00000000} /* (29, 1, 0) {real, imag} */,
  {32'h442ba2f6, 32'h00000000} /* (29, 0, 31) {real, imag} */,
  {32'h44af1eca, 32'h00000000} /* (29, 0, 30) {real, imag} */,
  {32'h44d93633, 32'h00000000} /* (29, 0, 29) {real, imag} */,
  {32'h44a08da2, 32'h00000000} /* (29, 0, 28) {real, imag} */,
  {32'h44c33f8b, 32'h00000000} /* (29, 0, 27) {real, imag} */,
  {32'h44cebeb7, 32'h00000000} /* (29, 0, 26) {real, imag} */,
  {32'h450773da, 32'h00000000} /* (29, 0, 25) {real, imag} */,
  {32'h45177ec4, 32'h00000000} /* (29, 0, 24) {real, imag} */,
  {32'h453277dc, 32'h00000000} /* (29, 0, 23) {real, imag} */,
  {32'h45107b53, 32'h00000000} /* (29, 0, 22) {real, imag} */,
  {32'h45127d07, 32'h00000000} /* (29, 0, 21) {real, imag} */,
  {32'h45099efb, 32'h00000000} /* (29, 0, 20) {real, imag} */,
  {32'h449e5d3f, 32'h00000000} /* (29, 0, 19) {real, imag} */,
  {32'h44c6fb5b, 32'h00000000} /* (29, 0, 18) {real, imag} */,
  {32'h4479d63c, 32'h00000000} /* (29, 0, 17) {real, imag} */,
  {32'hc3d7ffa4, 32'h00000000} /* (29, 0, 16) {real, imag} */,
  {32'hc4d3c41b, 32'h00000000} /* (29, 0, 15) {real, imag} */,
  {32'hc52ad8b5, 32'h00000000} /* (29, 0, 14) {real, imag} */,
  {32'hc581c47d, 32'h00000000} /* (29, 0, 13) {real, imag} */,
  {32'hc56bd273, 32'h00000000} /* (29, 0, 12) {real, imag} */,
  {32'hc5388ed2, 32'h00000000} /* (29, 0, 11) {real, imag} */,
  {32'hc5067ec4, 32'h00000000} /* (29, 0, 10) {real, imag} */,
  {32'hc50112b8, 32'h00000000} /* (29, 0, 9) {real, imag} */,
  {32'hc488e58e, 32'h00000000} /* (29, 0, 8) {real, imag} */,
  {32'hc486029b, 32'h00000000} /* (29, 0, 7) {real, imag} */,
  {32'hc4734368, 32'h00000000} /* (29, 0, 6) {real, imag} */,
  {32'h44a1e2bc, 32'h00000000} /* (29, 0, 5) {real, imag} */,
  {32'h44b40501, 32'h00000000} /* (29, 0, 4) {real, imag} */,
  {32'h4506b68e, 32'h00000000} /* (29, 0, 3) {real, imag} */,
  {32'h45196382, 32'h00000000} /* (29, 0, 2) {real, imag} */,
  {32'h44ae539e, 32'h00000000} /* (29, 0, 1) {real, imag} */,
  {32'h4481abf1, 32'h00000000} /* (29, 0, 0) {real, imag} */,
  {32'h423f9cc0, 32'h00000000} /* (28, 31, 31) {real, imag} */,
  {32'hc3901a00, 32'h00000000} /* (28, 31, 30) {real, imag} */,
  {32'h438bdab0, 32'h00000000} /* (28, 31, 29) {real, imag} */,
  {32'h447df510, 32'h00000000} /* (28, 31, 28) {real, imag} */,
  {32'h44bc9d92, 32'h00000000} /* (28, 31, 27) {real, imag} */,
  {32'h450f9755, 32'h00000000} /* (28, 31, 26) {real, imag} */,
  {32'h44da038b, 32'h00000000} /* (28, 31, 25) {real, imag} */,
  {32'h44bca465, 32'h00000000} /* (28, 31, 24) {real, imag} */,
  {32'h44d8b39d, 32'h00000000} /* (28, 31, 23) {real, imag} */,
  {32'h44ce92d6, 32'h00000000} /* (28, 31, 22) {real, imag} */,
  {32'h4485f3b4, 32'h00000000} /* (28, 31, 21) {real, imag} */,
  {32'h425d23d0, 32'h00000000} /* (28, 31, 20) {real, imag} */,
  {32'hc32af31c, 32'h00000000} /* (28, 31, 19) {real, imag} */,
  {32'hc3cc25ee, 32'h00000000} /* (28, 31, 18) {real, imag} */,
  {32'hc4aced4f, 32'h00000000} /* (28, 31, 17) {real, imag} */,
  {32'hc4c9280c, 32'h00000000} /* (28, 31, 16) {real, imag} */,
  {32'hc5191956, 32'h00000000} /* (28, 31, 15) {real, imag} */,
  {32'hc53f0460, 32'h00000000} /* (28, 31, 14) {real, imag} */,
  {32'hc55b97ee, 32'h00000000} /* (28, 31, 13) {real, imag} */,
  {32'hc54d6d50, 32'h00000000} /* (28, 31, 12) {real, imag} */,
  {32'hc4f8ca6c, 32'h00000000} /* (28, 31, 11) {real, imag} */,
  {32'hc4715cab, 32'h00000000} /* (28, 31, 10) {real, imag} */,
  {32'h42c34b10, 32'h00000000} /* (28, 31, 9) {real, imag} */,
  {32'h43fbf72b, 32'h00000000} /* (28, 31, 8) {real, imag} */,
  {32'h4445bf0a, 32'h00000000} /* (28, 31, 7) {real, imag} */,
  {32'h440c2efb, 32'h00000000} /* (28, 31, 6) {real, imag} */,
  {32'h448e3a60, 32'h00000000} /* (28, 31, 5) {real, imag} */,
  {32'h450102a3, 32'h00000000} /* (28, 31, 4) {real, imag} */,
  {32'h44c6fc64, 32'h00000000} /* (28, 31, 3) {real, imag} */,
  {32'h44edb766, 32'h00000000} /* (28, 31, 2) {real, imag} */,
  {32'h4495ce0b, 32'h00000000} /* (28, 31, 1) {real, imag} */,
  {32'h41e3a380, 32'h00000000} /* (28, 31, 0) {real, imag} */,
  {32'h443659f2, 32'h00000000} /* (28, 30, 31) {real, imag} */,
  {32'h430a8960, 32'h00000000} /* (28, 30, 30) {real, imag} */,
  {32'h44009266, 32'h00000000} /* (28, 30, 29) {real, imag} */,
  {32'h44c9bd0d, 32'h00000000} /* (28, 30, 28) {real, imag} */,
  {32'h45236abe, 32'h00000000} /* (28, 30, 27) {real, imag} */,
  {32'h452b5d1a, 32'h00000000} /* (28, 30, 26) {real, imag} */,
  {32'h452178e5, 32'h00000000} /* (28, 30, 25) {real, imag} */,
  {32'h45286d02, 32'h00000000} /* (28, 30, 24) {real, imag} */,
  {32'h451d938e, 32'h00000000} /* (28, 30, 23) {real, imag} */,
  {32'h44cc02dc, 32'h00000000} /* (28, 30, 22) {real, imag} */,
  {32'h44375230, 32'h00000000} /* (28, 30, 21) {real, imag} */,
  {32'hc443efd4, 32'h00000000} /* (28, 30, 20) {real, imag} */,
  {32'hc4a5dc5d, 32'h00000000} /* (28, 30, 19) {real, imag} */,
  {32'hc51c2d80, 32'h00000000} /* (28, 30, 18) {real, imag} */,
  {32'hc55e5296, 32'h00000000} /* (28, 30, 17) {real, imag} */,
  {32'hc5433138, 32'h00000000} /* (28, 30, 16) {real, imag} */,
  {32'hc557c922, 32'h00000000} /* (28, 30, 15) {real, imag} */,
  {32'hc585229d, 32'h00000000} /* (28, 30, 14) {real, imag} */,
  {32'hc56d2e64, 32'h00000000} /* (28, 30, 13) {real, imag} */,
  {32'hc56ec18e, 32'h00000000} /* (28, 30, 12) {real, imag} */,
  {32'hc51bd29a, 32'h00000000} /* (28, 30, 11) {real, imag} */,
  {32'hc390ef50, 32'h00000000} /* (28, 30, 10) {real, imag} */,
  {32'h4509b10f, 32'h00000000} /* (28, 30, 9) {real, imag} */,
  {32'h44dda147, 32'h00000000} /* (28, 30, 8) {real, imag} */,
  {32'h45252776, 32'h00000000} /* (28, 30, 7) {real, imag} */,
  {32'h44eb16b4, 32'h00000000} /* (28, 30, 6) {real, imag} */,
  {32'h4505e451, 32'h00000000} /* (28, 30, 5) {real, imag} */,
  {32'h454d6c5c, 32'h00000000} /* (28, 30, 4) {real, imag} */,
  {32'h452f4608, 32'h00000000} /* (28, 30, 3) {real, imag} */,
  {32'h44e5b6e9, 32'h00000000} /* (28, 30, 2) {real, imag} */,
  {32'h44728c02, 32'h00000000} /* (28, 30, 1) {real, imag} */,
  {32'h435e3278, 32'h00000000} /* (28, 30, 0) {real, imag} */,
  {32'h4474484c, 32'h00000000} /* (28, 29, 31) {real, imag} */,
  {32'h4492afbd, 32'h00000000} /* (28, 29, 30) {real, imag} */,
  {32'h44b22fd0, 32'h00000000} /* (28, 29, 29) {real, imag} */,
  {32'h45288836, 32'h00000000} /* (28, 29, 28) {real, imag} */,
  {32'h44f4c115, 32'h00000000} /* (28, 29, 27) {real, imag} */,
  {32'h45122da8, 32'h00000000} /* (28, 29, 26) {real, imag} */,
  {32'h455c5a66, 32'h00000000} /* (28, 29, 25) {real, imag} */,
  {32'h450f18ab, 32'h00000000} /* (28, 29, 24) {real, imag} */,
  {32'h44f12602, 32'h00000000} /* (28, 29, 23) {real, imag} */,
  {32'h44cb9b83, 32'h00000000} /* (28, 29, 22) {real, imag} */,
  {32'hc3181e80, 32'h00000000} /* (28, 29, 21) {real, imag} */,
  {32'hc50d1645, 32'h00000000} /* (28, 29, 20) {real, imag} */,
  {32'hc566d439, 32'h00000000} /* (28, 29, 19) {real, imag} */,
  {32'hc550d65a, 32'h00000000} /* (28, 29, 18) {real, imag} */,
  {32'hc55b60e4, 32'h00000000} /* (28, 29, 17) {real, imag} */,
  {32'hc584d0c7, 32'h00000000} /* (28, 29, 16) {real, imag} */,
  {32'hc5700c87, 32'h00000000} /* (28, 29, 15) {real, imag} */,
  {32'hc594b62c, 32'h00000000} /* (28, 29, 14) {real, imag} */,
  {32'hc5754f0c, 32'h00000000} /* (28, 29, 13) {real, imag} */,
  {32'hc554403a, 32'h00000000} /* (28, 29, 12) {real, imag} */,
  {32'hc4eb4d4b, 32'h00000000} /* (28, 29, 11) {real, imag} */,
  {32'h44097042, 32'h00000000} /* (28, 29, 10) {real, imag} */,
  {32'h44bfa15b, 32'h00000000} /* (28, 29, 9) {real, imag} */,
  {32'h4506822d, 32'h00000000} /* (28, 29, 8) {real, imag} */,
  {32'h453f2993, 32'h00000000} /* (28, 29, 7) {real, imag} */,
  {32'h45321d28, 32'h00000000} /* (28, 29, 6) {real, imag} */,
  {32'h452e415c, 32'h00000000} /* (28, 29, 5) {real, imag} */,
  {32'h4543a415, 32'h00000000} /* (28, 29, 4) {real, imag} */,
  {32'h452d5a05, 32'h00000000} /* (28, 29, 3) {real, imag} */,
  {32'h45059c54, 32'h00000000} /* (28, 29, 2) {real, imag} */,
  {32'h4457dcd2, 32'h00000000} /* (28, 29, 1) {real, imag} */,
  {32'h4407bf30, 32'h00000000} /* (28, 29, 0) {real, imag} */,
  {32'h4450936e, 32'h00000000} /* (28, 28, 31) {real, imag} */,
  {32'h448e4995, 32'h00000000} /* (28, 28, 30) {real, imag} */,
  {32'h44d37fe2, 32'h00000000} /* (28, 28, 29) {real, imag} */,
  {32'h452716e5, 32'h00000000} /* (28, 28, 28) {real, imag} */,
  {32'h44f1c0e9, 32'h00000000} /* (28, 28, 27) {real, imag} */,
  {32'h452b7d82, 32'h00000000} /* (28, 28, 26) {real, imag} */,
  {32'h45190e74, 32'h00000000} /* (28, 28, 25) {real, imag} */,
  {32'h45176734, 32'h00000000} /* (28, 28, 24) {real, imag} */,
  {32'h450e414c, 32'h00000000} /* (28, 28, 23) {real, imag} */,
  {32'h45133550, 32'h00000000} /* (28, 28, 22) {real, imag} */,
  {32'h4469c367, 32'h00000000} /* (28, 28, 21) {real, imag} */,
  {32'hc50644d6, 32'h00000000} /* (28, 28, 20) {real, imag} */,
  {32'hc58dcd92, 32'h00000000} /* (28, 28, 19) {real, imag} */,
  {32'hc555419c, 32'h00000000} /* (28, 28, 18) {real, imag} */,
  {32'hc5898698, 32'h00000000} /* (28, 28, 17) {real, imag} */,
  {32'hc5787e62, 32'h00000000} /* (28, 28, 16) {real, imag} */,
  {32'hc57a7976, 32'h00000000} /* (28, 28, 15) {real, imag} */,
  {32'hc593a9ae, 32'h00000000} /* (28, 28, 14) {real, imag} */,
  {32'hc56241a7, 32'h00000000} /* (28, 28, 13) {real, imag} */,
  {32'hc550a2a1, 32'h00000000} /* (28, 28, 12) {real, imag} */,
  {32'hc4da4baf, 32'h00000000} /* (28, 28, 11) {real, imag} */,
  {32'h44c529dc, 32'h00000000} /* (28, 28, 10) {real, imag} */,
  {32'h454ed22c, 32'h00000000} /* (28, 28, 9) {real, imag} */,
  {32'h45635a64, 32'h00000000} /* (28, 28, 8) {real, imag} */,
  {32'h4550f118, 32'h00000000} /* (28, 28, 7) {real, imag} */,
  {32'h4551fa2c, 32'h00000000} /* (28, 28, 6) {real, imag} */,
  {32'h4536a3c8, 32'h00000000} /* (28, 28, 5) {real, imag} */,
  {32'h45640524, 32'h00000000} /* (28, 28, 4) {real, imag} */,
  {32'h454341e4, 32'h00000000} /* (28, 28, 3) {real, imag} */,
  {32'h45162d46, 32'h00000000} /* (28, 28, 2) {real, imag} */,
  {32'h4463413c, 32'h00000000} /* (28, 28, 1) {real, imag} */,
  {32'h440cdba8, 32'h00000000} /* (28, 28, 0) {real, imag} */,
  {32'h44352206, 32'h00000000} /* (28, 27, 31) {real, imag} */,
  {32'h44bf0c21, 32'h00000000} /* (28, 27, 30) {real, imag} */,
  {32'h4525fe43, 32'h00000000} /* (28, 27, 29) {real, imag} */,
  {32'h4523f206, 32'h00000000} /* (28, 27, 28) {real, imag} */,
  {32'h44f614ef, 32'h00000000} /* (28, 27, 27) {real, imag} */,
  {32'h44ef62b1, 32'h00000000} /* (28, 27, 26) {real, imag} */,
  {32'h44ef1660, 32'h00000000} /* (28, 27, 25) {real, imag} */,
  {32'h4518df00, 32'h00000000} /* (28, 27, 24) {real, imag} */,
  {32'h44ae71cf, 32'h00000000} /* (28, 27, 23) {real, imag} */,
  {32'h450424ba, 32'h00000000} /* (28, 27, 22) {real, imag} */,
  {32'h44b09b50, 32'h00000000} /* (28, 27, 21) {real, imag} */,
  {32'hc4d2a3e0, 32'h00000000} /* (28, 27, 20) {real, imag} */,
  {32'hc52f60fc, 32'h00000000} /* (28, 27, 19) {real, imag} */,
  {32'hc571bcf8, 32'h00000000} /* (28, 27, 18) {real, imag} */,
  {32'hc55d0cfc, 32'h00000000} /* (28, 27, 17) {real, imag} */,
  {32'hc5909a7d, 32'h00000000} /* (28, 27, 16) {real, imag} */,
  {32'hc5717a92, 32'h00000000} /* (28, 27, 15) {real, imag} */,
  {32'hc56c787a, 32'h00000000} /* (28, 27, 14) {real, imag} */,
  {32'hc553f3a5, 32'h00000000} /* (28, 27, 13) {real, imag} */,
  {32'hc53a90e8, 32'h00000000} /* (28, 27, 12) {real, imag} */,
  {32'hc4bd5bcb, 32'h00000000} /* (28, 27, 11) {real, imag} */,
  {32'h44b37fcd, 32'h00000000} /* (28, 27, 10) {real, imag} */,
  {32'h456b40fa, 32'h00000000} /* (28, 27, 9) {real, imag} */,
  {32'h455da0a8, 32'h00000000} /* (28, 27, 8) {real, imag} */,
  {32'h45999306, 32'h00000000} /* (28, 27, 7) {real, imag} */,
  {32'h4548474a, 32'h00000000} /* (28, 27, 6) {real, imag} */,
  {32'h4583a94f, 32'h00000000} /* (28, 27, 5) {real, imag} */,
  {32'h454ca560, 32'h00000000} /* (28, 27, 4) {real, imag} */,
  {32'h45100fe2, 32'h00000000} /* (28, 27, 3) {real, imag} */,
  {32'h4523654e, 32'h00000000} /* (28, 27, 2) {real, imag} */,
  {32'h44a3d2b8, 32'h00000000} /* (28, 27, 1) {real, imag} */,
  {32'h44397d68, 32'h00000000} /* (28, 27, 0) {real, imag} */,
  {32'h446ca554, 32'h00000000} /* (28, 26, 31) {real, imag} */,
  {32'h449aed19, 32'h00000000} /* (28, 26, 30) {real, imag} */,
  {32'h448b74c6, 32'h00000000} /* (28, 26, 29) {real, imag} */,
  {32'h44c6064f, 32'h00000000} /* (28, 26, 28) {real, imag} */,
  {32'h45070edd, 32'h00000000} /* (28, 26, 27) {real, imag} */,
  {32'h452ca068, 32'h00000000} /* (28, 26, 26) {real, imag} */,
  {32'h44f80450, 32'h00000000} /* (28, 26, 25) {real, imag} */,
  {32'h45250af0, 32'h00000000} /* (28, 26, 24) {real, imag} */,
  {32'h4505035b, 32'h00000000} /* (28, 26, 23) {real, imag} */,
  {32'h44f195f8, 32'h00000000} /* (28, 26, 22) {real, imag} */,
  {32'h4476a1f4, 32'h00000000} /* (28, 26, 21) {real, imag} */,
  {32'hc4ff0f90, 32'h00000000} /* (28, 26, 20) {real, imag} */,
  {32'hc52c3e46, 32'h00000000} /* (28, 26, 19) {real, imag} */,
  {32'hc58a81af, 32'h00000000} /* (28, 26, 18) {real, imag} */,
  {32'hc57bf81b, 32'h00000000} /* (28, 26, 17) {real, imag} */,
  {32'hc59d619c, 32'h00000000} /* (28, 26, 16) {real, imag} */,
  {32'hc58079ac, 32'h00000000} /* (28, 26, 15) {real, imag} */,
  {32'hc55d7ad0, 32'h00000000} /* (28, 26, 14) {real, imag} */,
  {32'hc561a69b, 32'h00000000} /* (28, 26, 13) {real, imag} */,
  {32'hc50e60b0, 32'h00000000} /* (28, 26, 12) {real, imag} */,
  {32'hc4c52602, 32'h00000000} /* (28, 26, 11) {real, imag} */,
  {32'h43f5dae0, 32'h00000000} /* (28, 26, 10) {real, imag} */,
  {32'h453aafc4, 32'h00000000} /* (28, 26, 9) {real, imag} */,
  {32'h45966ef1, 32'h00000000} /* (28, 26, 8) {real, imag} */,
  {32'h4543bbb9, 32'h00000000} /* (28, 26, 7) {real, imag} */,
  {32'h4543fe84, 32'h00000000} /* (28, 26, 6) {real, imag} */,
  {32'h454cb2b3, 32'h00000000} /* (28, 26, 5) {real, imag} */,
  {32'h4520d18e, 32'h00000000} /* (28, 26, 4) {real, imag} */,
  {32'h450746cc, 32'h00000000} /* (28, 26, 3) {real, imag} */,
  {32'h44c074c8, 32'h00000000} /* (28, 26, 2) {real, imag} */,
  {32'h44dacf0e, 32'h00000000} /* (28, 26, 1) {real, imag} */,
  {32'h449b595a, 32'h00000000} /* (28, 26, 0) {real, imag} */,
  {32'h44d39acf, 32'h00000000} /* (28, 25, 31) {real, imag} */,
  {32'h44b88d1f, 32'h00000000} /* (28, 25, 30) {real, imag} */,
  {32'h44adad1c, 32'h00000000} /* (28, 25, 29) {real, imag} */,
  {32'h44db1bb2, 32'h00000000} /* (28, 25, 28) {real, imag} */,
  {32'h4506f343, 32'h00000000} /* (28, 25, 27) {real, imag} */,
  {32'h45162570, 32'h00000000} /* (28, 25, 26) {real, imag} */,
  {32'h4532d737, 32'h00000000} /* (28, 25, 25) {real, imag} */,
  {32'h45186a0e, 32'h00000000} /* (28, 25, 24) {real, imag} */,
  {32'h45384a86, 32'h00000000} /* (28, 25, 23) {real, imag} */,
  {32'h45373c89, 32'h00000000} /* (28, 25, 22) {real, imag} */,
  {32'h43fd7a44, 32'h00000000} /* (28, 25, 21) {real, imag} */,
  {32'hc4e7eb98, 32'h00000000} /* (28, 25, 20) {real, imag} */,
  {32'hc50ba9f9, 32'h00000000} /* (28, 25, 19) {real, imag} */,
  {32'hc54c4860, 32'h00000000} /* (28, 25, 18) {real, imag} */,
  {32'hc5571b74, 32'h00000000} /* (28, 25, 17) {real, imag} */,
  {32'hc55b9a15, 32'h00000000} /* (28, 25, 16) {real, imag} */,
  {32'hc56ffab6, 32'h00000000} /* (28, 25, 15) {real, imag} */,
  {32'hc5520548, 32'h00000000} /* (28, 25, 14) {real, imag} */,
  {32'hc53c6bd8, 32'h00000000} /* (28, 25, 13) {real, imag} */,
  {32'hc52850cb, 32'h00000000} /* (28, 25, 12) {real, imag} */,
  {32'hc47a2fcc, 32'h00000000} /* (28, 25, 11) {real, imag} */,
  {32'h44597255, 32'h00000000} /* (28, 25, 10) {real, imag} */,
  {32'h45142653, 32'h00000000} /* (28, 25, 9) {real, imag} */,
  {32'h457b3236, 32'h00000000} /* (28, 25, 8) {real, imag} */,
  {32'h4547fa02, 32'h00000000} /* (28, 25, 7) {real, imag} */,
  {32'h4536e4cb, 32'h00000000} /* (28, 25, 6) {real, imag} */,
  {32'h4579ee04, 32'h00000000} /* (28, 25, 5) {real, imag} */,
  {32'h4524a5aa, 32'h00000000} /* (28, 25, 4) {real, imag} */,
  {32'h44d5f96b, 32'h00000000} /* (28, 25, 3) {real, imag} */,
  {32'h44aa0b03, 32'h00000000} /* (28, 25, 2) {real, imag} */,
  {32'h4487cdf4, 32'h00000000} /* (28, 25, 1) {real, imag} */,
  {32'h44b293ca, 32'h00000000} /* (28, 25, 0) {real, imag} */,
  {32'h44203c8c, 32'h00000000} /* (28, 24, 31) {real, imag} */,
  {32'h44d79a09, 32'h00000000} /* (28, 24, 30) {real, imag} */,
  {32'h44b35360, 32'h00000000} /* (28, 24, 29) {real, imag} */,
  {32'h44b682f6, 32'h00000000} /* (28, 24, 28) {real, imag} */,
  {32'h45439b38, 32'h00000000} /* (28, 24, 27) {real, imag} */,
  {32'h4519b24a, 32'h00000000} /* (28, 24, 26) {real, imag} */,
  {32'h455bcc00, 32'h00000000} /* (28, 24, 25) {real, imag} */,
  {32'h4537979e, 32'h00000000} /* (28, 24, 24) {real, imag} */,
  {32'h4531e728, 32'h00000000} /* (28, 24, 23) {real, imag} */,
  {32'h45041a6b, 32'h00000000} /* (28, 24, 22) {real, imag} */,
  {32'h442475b8, 32'h00000000} /* (28, 24, 21) {real, imag} */,
  {32'hc42c1304, 32'h00000000} /* (28, 24, 20) {real, imag} */,
  {32'hc5043821, 32'h00000000} /* (28, 24, 19) {real, imag} */,
  {32'hc51b2415, 32'h00000000} /* (28, 24, 18) {real, imag} */,
  {32'hc52882a2, 32'h00000000} /* (28, 24, 17) {real, imag} */,
  {32'hc55654c6, 32'h00000000} /* (28, 24, 16) {real, imag} */,
  {32'hc58f1702, 32'h00000000} /* (28, 24, 15) {real, imag} */,
  {32'hc5a36159, 32'h00000000} /* (28, 24, 14) {real, imag} */,
  {32'hc54fc0d2, 32'h00000000} /* (28, 24, 13) {real, imag} */,
  {32'hc4e55e54, 32'h00000000} /* (28, 24, 12) {real, imag} */,
  {32'hc4aa0437, 32'h00000000} /* (28, 24, 11) {real, imag} */,
  {32'h4462022e, 32'h00000000} /* (28, 24, 10) {real, imag} */,
  {32'h4526c81c, 32'h00000000} /* (28, 24, 9) {real, imag} */,
  {32'h45914d9f, 32'h00000000} /* (28, 24, 8) {real, imag} */,
  {32'h4582da34, 32'h00000000} /* (28, 24, 7) {real, imag} */,
  {32'h4557b559, 32'h00000000} /* (28, 24, 6) {real, imag} */,
  {32'h45429080, 32'h00000000} /* (28, 24, 5) {real, imag} */,
  {32'h4524cfa6, 32'h00000000} /* (28, 24, 4) {real, imag} */,
  {32'h4503b62f, 32'h00000000} /* (28, 24, 3) {real, imag} */,
  {32'h44c9d6c2, 32'h00000000} /* (28, 24, 2) {real, imag} */,
  {32'h44bab0fd, 32'h00000000} /* (28, 24, 1) {real, imag} */,
  {32'h44537cf2, 32'h00000000} /* (28, 24, 0) {real, imag} */,
  {32'h44599170, 32'h00000000} /* (28, 23, 31) {real, imag} */,
  {32'h44c6d080, 32'h00000000} /* (28, 23, 30) {real, imag} */,
  {32'h44d1a6b0, 32'h00000000} /* (28, 23, 29) {real, imag} */,
  {32'h44f1aa85, 32'h00000000} /* (28, 23, 28) {real, imag} */,
  {32'h45342ebf, 32'h00000000} /* (28, 23, 27) {real, imag} */,
  {32'h45657742, 32'h00000000} /* (28, 23, 26) {real, imag} */,
  {32'h4505140b, 32'h00000000} /* (28, 23, 25) {real, imag} */,
  {32'h451943d4, 32'h00000000} /* (28, 23, 24) {real, imag} */,
  {32'h451a083b, 32'h00000000} /* (28, 23, 23) {real, imag} */,
  {32'h44cbd904, 32'h00000000} /* (28, 23, 22) {real, imag} */,
  {32'h4501c8ed, 32'h00000000} /* (28, 23, 21) {real, imag} */,
  {32'hc4037fbc, 32'h00000000} /* (28, 23, 20) {real, imag} */,
  {32'hc50af292, 32'h00000000} /* (28, 23, 19) {real, imag} */,
  {32'hc5292c9f, 32'h00000000} /* (28, 23, 18) {real, imag} */,
  {32'hc509127b, 32'h00000000} /* (28, 23, 17) {real, imag} */,
  {32'hc53ce5e6, 32'h00000000} /* (28, 23, 16) {real, imag} */,
  {32'hc5589760, 32'h00000000} /* (28, 23, 15) {real, imag} */,
  {32'hc544d99c, 32'h00000000} /* (28, 23, 14) {real, imag} */,
  {32'hc4cf2b26, 32'h00000000} /* (28, 23, 13) {real, imag} */,
  {32'hc4c4ed0b, 32'h00000000} /* (28, 23, 12) {real, imag} */,
  {32'hc48caed0, 32'h00000000} /* (28, 23, 11) {real, imag} */,
  {32'h43483ca0, 32'h00000000} /* (28, 23, 10) {real, imag} */,
  {32'h4536e2ef, 32'h00000000} /* (28, 23, 9) {real, imag} */,
  {32'h4545bc76, 32'h00000000} /* (28, 23, 8) {real, imag} */,
  {32'h456129cd, 32'h00000000} /* (28, 23, 7) {real, imag} */,
  {32'h452acb30, 32'h00000000} /* (28, 23, 6) {real, imag} */,
  {32'h451c6f4f, 32'h00000000} /* (28, 23, 5) {real, imag} */,
  {32'h44be2fa7, 32'h00000000} /* (28, 23, 4) {real, imag} */,
  {32'h44fed568, 32'h00000000} /* (28, 23, 3) {real, imag} */,
  {32'h44d02c02, 32'h00000000} /* (28, 23, 2) {real, imag} */,
  {32'h448fdfea, 32'h00000000} /* (28, 23, 1) {real, imag} */,
  {32'h442ef458, 32'h00000000} /* (28, 23, 0) {real, imag} */,
  {32'h44331ae1, 32'h00000000} /* (28, 22, 31) {real, imag} */,
  {32'h45210a0f, 32'h00000000} /* (28, 22, 30) {real, imag} */,
  {32'h44f3fd52, 32'h00000000} /* (28, 22, 29) {real, imag} */,
  {32'h449f9ba8, 32'h00000000} /* (28, 22, 28) {real, imag} */,
  {32'h44d542e3, 32'h00000000} /* (28, 22, 27) {real, imag} */,
  {32'h44cae093, 32'h00000000} /* (28, 22, 26) {real, imag} */,
  {32'h445c9742, 32'h00000000} /* (28, 22, 25) {real, imag} */,
  {32'h448b5492, 32'h00000000} /* (28, 22, 24) {real, imag} */,
  {32'h44bc7dc6, 32'h00000000} /* (28, 22, 23) {real, imag} */,
  {32'h44e23476, 32'h00000000} /* (28, 22, 22) {real, imag} */,
  {32'h44138ffc, 32'h00000000} /* (28, 22, 21) {real, imag} */,
  {32'hc3da78e6, 32'h00000000} /* (28, 22, 20) {real, imag} */,
  {32'hc48a588d, 32'h00000000} /* (28, 22, 19) {real, imag} */,
  {32'hc4a325f9, 32'h00000000} /* (28, 22, 18) {real, imag} */,
  {32'hc462d7ce, 32'h00000000} /* (28, 22, 17) {real, imag} */,
  {32'hc4e9c05c, 32'h00000000} /* (28, 22, 16) {real, imag} */,
  {32'hc4d50e2e, 32'h00000000} /* (28, 22, 15) {real, imag} */,
  {32'hc4a46b42, 32'h00000000} /* (28, 22, 14) {real, imag} */,
  {32'hc4814400, 32'h00000000} /* (28, 22, 13) {real, imag} */,
  {32'hc3878e5f, 32'h00000000} /* (28, 22, 12) {real, imag} */,
  {32'hc31d2e68, 32'h00000000} /* (28, 22, 11) {real, imag} */,
  {32'h43fc9dec, 32'h00000000} /* (28, 22, 10) {real, imag} */,
  {32'h44c55fa7, 32'h00000000} /* (28, 22, 9) {real, imag} */,
  {32'h450d5a65, 32'h00000000} /* (28, 22, 8) {real, imag} */,
  {32'h45002d41, 32'h00000000} /* (28, 22, 7) {real, imag} */,
  {32'h44c9b13e, 32'h00000000} /* (28, 22, 6) {real, imag} */,
  {32'h44990f74, 32'h00000000} /* (28, 22, 5) {real, imag} */,
  {32'h44f0299c, 32'h00000000} /* (28, 22, 4) {real, imag} */,
  {32'h44d6feb5, 32'h00000000} /* (28, 22, 3) {real, imag} */,
  {32'h4467ba1e, 32'h00000000} /* (28, 22, 2) {real, imag} */,
  {32'h44838a22, 32'h00000000} /* (28, 22, 1) {real, imag} */,
  {32'h440854b0, 32'h00000000} /* (28, 22, 0) {real, imag} */,
  {32'hc3c8581c, 32'h00000000} /* (28, 21, 31) {real, imag} */,
  {32'hc415202f, 32'h00000000} /* (28, 21, 30) {real, imag} */,
  {32'h4411054d, 32'h00000000} /* (28, 21, 29) {real, imag} */,
  {32'h424bda12, 32'h00000000} /* (28, 21, 28) {real, imag} */,
  {32'hc3d9a910, 32'h00000000} /* (28, 21, 27) {real, imag} */,
  {32'hc432679d, 32'h00000000} /* (28, 21, 26) {real, imag} */,
  {32'hc3d7e291, 32'h00000000} /* (28, 21, 25) {real, imag} */,
  {32'h440769fd, 32'h00000000} /* (28, 21, 24) {real, imag} */,
  {32'h42a45895, 32'h00000000} /* (28, 21, 23) {real, imag} */,
  {32'hc2ece03c, 32'h00000000} /* (28, 21, 22) {real, imag} */,
  {32'h43ab421e, 32'h00000000} /* (28, 21, 21) {real, imag} */,
  {32'h434873b1, 32'h00000000} /* (28, 21, 20) {real, imag} */,
  {32'h42fd7b60, 32'h00000000} /* (28, 21, 19) {real, imag} */,
  {32'h436e87b2, 32'h00000000} /* (28, 21, 18) {real, imag} */,
  {32'h4387f1bb, 32'h00000000} /* (28, 21, 17) {real, imag} */,
  {32'hc3048210, 32'h00000000} /* (28, 21, 16) {real, imag} */,
  {32'hc23a9fa0, 32'h00000000} /* (28, 21, 15) {real, imag} */,
  {32'hc3cfbb8a, 32'h00000000} /* (28, 21, 14) {real, imag} */,
  {32'h4444d743, 32'h00000000} /* (28, 21, 13) {real, imag} */,
  {32'h439384fa, 32'h00000000} /* (28, 21, 12) {real, imag} */,
  {32'hc39d666c, 32'h00000000} /* (28, 21, 11) {real, imag} */,
  {32'h44549e07, 32'h00000000} /* (28, 21, 10) {real, imag} */,
  {32'h432f739e, 32'h00000000} /* (28, 21, 9) {real, imag} */,
  {32'h41aeeca0, 32'h00000000} /* (28, 21, 8) {real, imag} */,
  {32'hc2f7c38f, 32'h00000000} /* (28, 21, 7) {real, imag} */,
  {32'h41de8680, 32'h00000000} /* (28, 21, 6) {real, imag} */,
  {32'hc3f93d46, 32'h00000000} /* (28, 21, 5) {real, imag} */,
  {32'h4422afe2, 32'h00000000} /* (28, 21, 4) {real, imag} */,
  {32'hc392f69c, 32'h00000000} /* (28, 21, 3) {real, imag} */,
  {32'hc4215166, 32'h00000000} /* (28, 21, 2) {real, imag} */,
  {32'h438182c7, 32'h00000000} /* (28, 21, 1) {real, imag} */,
  {32'hc3af52f5, 32'h00000000} /* (28, 21, 0) {real, imag} */,
  {32'hc4e47ee3, 32'h00000000} /* (28, 20, 31) {real, imag} */,
  {32'hc50790d8, 32'h00000000} /* (28, 20, 30) {real, imag} */,
  {32'hc4d3d338, 32'h00000000} /* (28, 20, 29) {real, imag} */,
  {32'hc50c1e70, 32'h00000000} /* (28, 20, 28) {real, imag} */,
  {32'hc51a23ae, 32'h00000000} /* (28, 20, 27) {real, imag} */,
  {32'hc50508ff, 32'h00000000} /* (28, 20, 26) {real, imag} */,
  {32'hc546a70c, 32'h00000000} /* (28, 20, 25) {real, imag} */,
  {32'hc52ad6fc, 32'h00000000} /* (28, 20, 24) {real, imag} */,
  {32'hc4d14e7e, 32'h00000000} /* (28, 20, 23) {real, imag} */,
  {32'hc4cdfe45, 32'h00000000} /* (28, 20, 22) {real, imag} */,
  {32'hc31ffde0, 32'h00000000} /* (28, 20, 21) {real, imag} */,
  {32'h44ae5964, 32'h00000000} /* (28, 20, 20) {real, imag} */,
  {32'h44f1766c, 32'h00000000} /* (28, 20, 19) {real, imag} */,
  {32'h44f7aaa1, 32'h00000000} /* (28, 20, 18) {real, imag} */,
  {32'h44c64c6f, 32'h00000000} /* (28, 20, 17) {real, imag} */,
  {32'h44f26900, 32'h00000000} /* (28, 20, 16) {real, imag} */,
  {32'h451465da, 32'h00000000} /* (28, 20, 15) {real, imag} */,
  {32'h4515af9a, 32'h00000000} /* (28, 20, 14) {real, imag} */,
  {32'h4522a7fc, 32'h00000000} /* (28, 20, 13) {real, imag} */,
  {32'h44f19a10, 32'h00000000} /* (28, 20, 12) {real, imag} */,
  {32'h44ea044c, 32'h00000000} /* (28, 20, 11) {real, imag} */,
  {32'h44197f4c, 32'h00000000} /* (28, 20, 10) {real, imag} */,
  {32'hc36c3920, 32'h00000000} /* (28, 20, 9) {real, imag} */,
  {32'hc5172e78, 32'h00000000} /* (28, 20, 8) {real, imag} */,
  {32'hc4d02338, 32'h00000000} /* (28, 20, 7) {real, imag} */,
  {32'hc4dcf253, 32'h00000000} /* (28, 20, 6) {real, imag} */,
  {32'hc53cb53c, 32'h00000000} /* (28, 20, 5) {real, imag} */,
  {32'hc51e82d1, 32'h00000000} /* (28, 20, 4) {real, imag} */,
  {32'hc4b14ef4, 32'h00000000} /* (28, 20, 3) {real, imag} */,
  {32'hc5477b7e, 32'h00000000} /* (28, 20, 2) {real, imag} */,
  {32'hc516b136, 32'h00000000} /* (28, 20, 1) {real, imag} */,
  {32'hc4570800, 32'h00000000} /* (28, 20, 0) {real, imag} */,
  {32'hc51b80a2, 32'h00000000} /* (28, 19, 31) {real, imag} */,
  {32'hc552f57a, 32'h00000000} /* (28, 19, 30) {real, imag} */,
  {32'hc520f2a8, 32'h00000000} /* (28, 19, 29) {real, imag} */,
  {32'hc54685ad, 32'h00000000} /* (28, 19, 28) {real, imag} */,
  {32'hc559b7d7, 32'h00000000} /* (28, 19, 27) {real, imag} */,
  {32'hc558fe5a, 32'h00000000} /* (28, 19, 26) {real, imag} */,
  {32'hc55184c6, 32'h00000000} /* (28, 19, 25) {real, imag} */,
  {32'hc55de348, 32'h00000000} /* (28, 19, 24) {real, imag} */,
  {32'hc53a8e00, 32'h00000000} /* (28, 19, 23) {real, imag} */,
  {32'hc4f3a649, 32'h00000000} /* (28, 19, 22) {real, imag} */,
  {32'hc44b7a4c, 32'h00000000} /* (28, 19, 21) {real, imag} */,
  {32'h44746698, 32'h00000000} /* (28, 19, 20) {real, imag} */,
  {32'h451fcd49, 32'h00000000} /* (28, 19, 19) {real, imag} */,
  {32'h4517c502, 32'h00000000} /* (28, 19, 18) {real, imag} */,
  {32'h45159d79, 32'h00000000} /* (28, 19, 17) {real, imag} */,
  {32'h4544f488, 32'h00000000} /* (28, 19, 16) {real, imag} */,
  {32'h455ad606, 32'h00000000} /* (28, 19, 15) {real, imag} */,
  {32'h4547665a, 32'h00000000} /* (28, 19, 14) {real, imag} */,
  {32'h453543f4, 32'h00000000} /* (28, 19, 13) {real, imag} */,
  {32'h44ee533a, 32'h00000000} /* (28, 19, 12) {real, imag} */,
  {32'h44a7373a, 32'h00000000} /* (28, 19, 11) {real, imag} */,
  {32'h4381b2bc, 32'h00000000} /* (28, 19, 10) {real, imag} */,
  {32'hc4a9ad74, 32'h00000000} /* (28, 19, 9) {real, imag} */,
  {32'hc4f81fc8, 32'h00000000} /* (28, 19, 8) {real, imag} */,
  {32'hc50eabd8, 32'h00000000} /* (28, 19, 7) {real, imag} */,
  {32'hc52e559e, 32'h00000000} /* (28, 19, 6) {real, imag} */,
  {32'hc585844e, 32'h00000000} /* (28, 19, 5) {real, imag} */,
  {32'hc5584318, 32'h00000000} /* (28, 19, 4) {real, imag} */,
  {32'hc53e3fbb, 32'h00000000} /* (28, 19, 3) {real, imag} */,
  {32'hc5658752, 32'h00000000} /* (28, 19, 2) {real, imag} */,
  {32'hc551216d, 32'h00000000} /* (28, 19, 1) {real, imag} */,
  {32'hc5611d90, 32'h00000000} /* (28, 19, 0) {real, imag} */,
  {32'hc530d183, 32'h00000000} /* (28, 18, 31) {real, imag} */,
  {32'hc57f450a, 32'h00000000} /* (28, 18, 30) {real, imag} */,
  {32'hc576b3c0, 32'h00000000} /* (28, 18, 29) {real, imag} */,
  {32'hc56b3679, 32'h00000000} /* (28, 18, 28) {real, imag} */,
  {32'hc583d330, 32'h00000000} /* (28, 18, 27) {real, imag} */,
  {32'hc582cad6, 32'h00000000} /* (28, 18, 26) {real, imag} */,
  {32'hc5706592, 32'h00000000} /* (28, 18, 25) {real, imag} */,
  {32'hc551abf8, 32'h00000000} /* (28, 18, 24) {real, imag} */,
  {32'hc5675b61, 32'h00000000} /* (28, 18, 23) {real, imag} */,
  {32'hc577f757, 32'h00000000} /* (28, 18, 22) {real, imag} */,
  {32'hc51f6df0, 32'h00000000} /* (28, 18, 21) {real, imag} */,
  {32'h443c5128, 32'h00000000} /* (28, 18, 20) {real, imag} */,
  {32'h4508fac0, 32'h00000000} /* (28, 18, 19) {real, imag} */,
  {32'h4558e672, 32'h00000000} /* (28, 18, 18) {real, imag} */,
  {32'h4532d2e8, 32'h00000000} /* (28, 18, 17) {real, imag} */,
  {32'h4573466c, 32'h00000000} /* (28, 18, 16) {real, imag} */,
  {32'h4565fb77, 32'h00000000} /* (28, 18, 15) {real, imag} */,
  {32'h456ddf06, 32'h00000000} /* (28, 18, 14) {real, imag} */,
  {32'h4580a621, 32'h00000000} /* (28, 18, 13) {real, imag} */,
  {32'h4511d5a9, 32'h00000000} /* (28, 18, 12) {real, imag} */,
  {32'h44b2c1af, 32'h00000000} /* (28, 18, 11) {real, imag} */,
  {32'hc0588000, 32'h00000000} /* (28, 18, 10) {real, imag} */,
  {32'hc4e313dd, 32'h00000000} /* (28, 18, 9) {real, imag} */,
  {32'hc53d691c, 32'h00000000} /* (28, 18, 8) {real, imag} */,
  {32'hc545ede7, 32'h00000000} /* (28, 18, 7) {real, imag} */,
  {32'hc55b9611, 32'h00000000} /* (28, 18, 6) {real, imag} */,
  {32'hc58bd71a, 32'h00000000} /* (28, 18, 5) {real, imag} */,
  {32'hc582d7af, 32'h00000000} /* (28, 18, 4) {real, imag} */,
  {32'hc55c708c, 32'h00000000} /* (28, 18, 3) {real, imag} */,
  {32'hc58333ea, 32'h00000000} /* (28, 18, 2) {real, imag} */,
  {32'hc5619d6e, 32'h00000000} /* (28, 18, 1) {real, imag} */,
  {32'hc562f8d8, 32'h00000000} /* (28, 18, 0) {real, imag} */,
  {32'hc5499008, 32'h00000000} /* (28, 17, 31) {real, imag} */,
  {32'hc58812d8, 32'h00000000} /* (28, 17, 30) {real, imag} */,
  {32'hc5a04cbc, 32'h00000000} /* (28, 17, 29) {real, imag} */,
  {32'hc5873912, 32'h00000000} /* (28, 17, 28) {real, imag} */,
  {32'hc597a702, 32'h00000000} /* (28, 17, 27) {real, imag} */,
  {32'hc5a58ec0, 32'h00000000} /* (28, 17, 26) {real, imag} */,
  {32'hc59f2840, 32'h00000000} /* (28, 17, 25) {real, imag} */,
  {32'hc57a994f, 32'h00000000} /* (28, 17, 24) {real, imag} */,
  {32'hc598fc70, 32'h00000000} /* (28, 17, 23) {real, imag} */,
  {32'hc53acdb5, 32'h00000000} /* (28, 17, 22) {real, imag} */,
  {32'hc4cf631d, 32'h00000000} /* (28, 17, 21) {real, imag} */,
  {32'h4439a33c, 32'h00000000} /* (28, 17, 20) {real, imag} */,
  {32'h4502a021, 32'h00000000} /* (28, 17, 19) {real, imag} */,
  {32'h455721a0, 32'h00000000} /* (28, 17, 18) {real, imag} */,
  {32'h4539bab6, 32'h00000000} /* (28, 17, 17) {real, imag} */,
  {32'h4550ff0d, 32'h00000000} /* (28, 17, 16) {real, imag} */,
  {32'h45598f6c, 32'h00000000} /* (28, 17, 15) {real, imag} */,
  {32'h4587f0dc, 32'h00000000} /* (28, 17, 14) {real, imag} */,
  {32'h453431d3, 32'h00000000} /* (28, 17, 13) {real, imag} */,
  {32'h452c7cf6, 32'h00000000} /* (28, 17, 12) {real, imag} */,
  {32'h44aca646, 32'h00000000} /* (28, 17, 11) {real, imag} */,
  {32'hc376f510, 32'h00000000} /* (28, 17, 10) {real, imag} */,
  {32'hc4ba9dff, 32'h00000000} /* (28, 17, 9) {real, imag} */,
  {32'hc52742cb, 32'h00000000} /* (28, 17, 8) {real, imag} */,
  {32'hc56d45c9, 32'h00000000} /* (28, 17, 7) {real, imag} */,
  {32'hc581c23c, 32'h00000000} /* (28, 17, 6) {real, imag} */,
  {32'hc55d0096, 32'h00000000} /* (28, 17, 5) {real, imag} */,
  {32'hc5853d08, 32'h00000000} /* (28, 17, 4) {real, imag} */,
  {32'hc5958ea0, 32'h00000000} /* (28, 17, 3) {real, imag} */,
  {32'hc56052c4, 32'h00000000} /* (28, 17, 2) {real, imag} */,
  {32'hc560f0da, 32'h00000000} /* (28, 17, 1) {real, imag} */,
  {32'hc53370fb, 32'h00000000} /* (28, 17, 0) {real, imag} */,
  {32'hc5422719, 32'h00000000} /* (28, 16, 31) {real, imag} */,
  {32'hc58f4b1a, 32'h00000000} /* (28, 16, 30) {real, imag} */,
  {32'hc57d06e3, 32'h00000000} /* (28, 16, 29) {real, imag} */,
  {32'hc5986064, 32'h00000000} /* (28, 16, 28) {real, imag} */,
  {32'hc584795a, 32'h00000000} /* (28, 16, 27) {real, imag} */,
  {32'hc58c7070, 32'h00000000} /* (28, 16, 26) {real, imag} */,
  {32'hc599b4a6, 32'h00000000} /* (28, 16, 25) {real, imag} */,
  {32'hc5865c76, 32'h00000000} /* (28, 16, 24) {real, imag} */,
  {32'hc57b9b18, 32'h00000000} /* (28, 16, 23) {real, imag} */,
  {32'hc50e7901, 32'h00000000} /* (28, 16, 22) {real, imag} */,
  {32'hc4ce7c53, 32'h00000000} /* (28, 16, 21) {real, imag} */,
  {32'h4476a0ac, 32'h00000000} /* (28, 16, 20) {real, imag} */,
  {32'h44da4db1, 32'h00000000} /* (28, 16, 19) {real, imag} */,
  {32'h452bf0c8, 32'h00000000} /* (28, 16, 18) {real, imag} */,
  {32'h4583fafd, 32'h00000000} /* (28, 16, 17) {real, imag} */,
  {32'h458768ee, 32'h00000000} /* (28, 16, 16) {real, imag} */,
  {32'h45655273, 32'h00000000} /* (28, 16, 15) {real, imag} */,
  {32'h454e4ebb, 32'h00000000} /* (28, 16, 14) {real, imag} */,
  {32'h4543964d, 32'h00000000} /* (28, 16, 13) {real, imag} */,
  {32'h450df45f, 32'h00000000} /* (28, 16, 12) {real, imag} */,
  {32'h44d249e7, 32'h00000000} /* (28, 16, 11) {real, imag} */,
  {32'h42bcb200, 32'h00000000} /* (28, 16, 10) {real, imag} */,
  {32'hc4fb4bf6, 32'h00000000} /* (28, 16, 9) {real, imag} */,
  {32'hc56a1f35, 32'h00000000} /* (28, 16, 8) {real, imag} */,
  {32'hc580d0f3, 32'h00000000} /* (28, 16, 7) {real, imag} */,
  {32'hc57eb827, 32'h00000000} /* (28, 16, 6) {real, imag} */,
  {32'hc5858394, 32'h00000000} /* (28, 16, 5) {real, imag} */,
  {32'hc5913df6, 32'h00000000} /* (28, 16, 4) {real, imag} */,
  {32'hc5505164, 32'h00000000} /* (28, 16, 3) {real, imag} */,
  {32'hc55c8772, 32'h00000000} /* (28, 16, 2) {real, imag} */,
  {32'hc56c7c44, 32'h00000000} /* (28, 16, 1) {real, imag} */,
  {32'hc53eca20, 32'h00000000} /* (28, 16, 0) {real, imag} */,
  {32'hc542e33c, 32'h00000000} /* (28, 15, 31) {real, imag} */,
  {32'hc590a18d, 32'h00000000} /* (28, 15, 30) {real, imag} */,
  {32'hc56679d2, 32'h00000000} /* (28, 15, 29) {real, imag} */,
  {32'hc56c5786, 32'h00000000} /* (28, 15, 28) {real, imag} */,
  {32'hc56b56c4, 32'h00000000} /* (28, 15, 27) {real, imag} */,
  {32'hc586c228, 32'h00000000} /* (28, 15, 26) {real, imag} */,
  {32'hc596eba0, 32'h00000000} /* (28, 15, 25) {real, imag} */,
  {32'hc5856cb8, 32'h00000000} /* (28, 15, 24) {real, imag} */,
  {32'hc57a34d2, 32'h00000000} /* (28, 15, 23) {real, imag} */,
  {32'hc53d223e, 32'h00000000} /* (28, 15, 22) {real, imag} */,
  {32'hc43fe538, 32'h00000000} /* (28, 15, 21) {real, imag} */,
  {32'h44b43b92, 32'h00000000} /* (28, 15, 20) {real, imag} */,
  {32'h45057471, 32'h00000000} /* (28, 15, 19) {real, imag} */,
  {32'h4536d3c2, 32'h00000000} /* (28, 15, 18) {real, imag} */,
  {32'h455fb89e, 32'h00000000} /* (28, 15, 17) {real, imag} */,
  {32'h457b0a8d, 32'h00000000} /* (28, 15, 16) {real, imag} */,
  {32'h458256c3, 32'h00000000} /* (28, 15, 15) {real, imag} */,
  {32'h452bc9a2, 32'h00000000} /* (28, 15, 14) {real, imag} */,
  {32'h454fe49a, 32'h00000000} /* (28, 15, 13) {real, imag} */,
  {32'h45496c4e, 32'h00000000} /* (28, 15, 12) {real, imag} */,
  {32'h44ef5768, 32'h00000000} /* (28, 15, 11) {real, imag} */,
  {32'hc4598e54, 32'h00000000} /* (28, 15, 10) {real, imag} */,
  {32'hc5127a38, 32'h00000000} /* (28, 15, 9) {real, imag} */,
  {32'hc579d650, 32'h00000000} /* (28, 15, 8) {real, imag} */,
  {32'hc589d1b7, 32'h00000000} /* (28, 15, 7) {real, imag} */,
  {32'hc58dbb27, 32'h00000000} /* (28, 15, 6) {real, imag} */,
  {32'hc588569f, 32'h00000000} /* (28, 15, 5) {real, imag} */,
  {32'hc57156d9, 32'h00000000} /* (28, 15, 4) {real, imag} */,
  {32'hc5788b77, 32'h00000000} /* (28, 15, 3) {real, imag} */,
  {32'hc54fe65c, 32'h00000000} /* (28, 15, 2) {real, imag} */,
  {32'hc567f37c, 32'h00000000} /* (28, 15, 1) {real, imag} */,
  {32'hc54269d9, 32'h00000000} /* (28, 15, 0) {real, imag} */,
  {32'hc53a42a9, 32'h00000000} /* (28, 14, 31) {real, imag} */,
  {32'hc5476d6d, 32'h00000000} /* (28, 14, 30) {real, imag} */,
  {32'hc56ed668, 32'h00000000} /* (28, 14, 29) {real, imag} */,
  {32'hc558cb79, 32'h00000000} /* (28, 14, 28) {real, imag} */,
  {32'hc54a9864, 32'h00000000} /* (28, 14, 27) {real, imag} */,
  {32'hc57d0180, 32'h00000000} /* (28, 14, 26) {real, imag} */,
  {32'hc5817df4, 32'h00000000} /* (28, 14, 25) {real, imag} */,
  {32'hc598edc7, 32'h00000000} /* (28, 14, 24) {real, imag} */,
  {32'hc58206ea, 32'h00000000} /* (28, 14, 23) {real, imag} */,
  {32'hc52a2e24, 32'h00000000} /* (28, 14, 22) {real, imag} */,
  {32'hc4385ace, 32'h00000000} /* (28, 14, 21) {real, imag} */,
  {32'h4489fa88, 32'h00000000} /* (28, 14, 20) {real, imag} */,
  {32'h451b7be6, 32'h00000000} /* (28, 14, 19) {real, imag} */,
  {32'h45447f50, 32'h00000000} /* (28, 14, 18) {real, imag} */,
  {32'h4549425a, 32'h00000000} /* (28, 14, 17) {real, imag} */,
  {32'h457a4081, 32'h00000000} /* (28, 14, 16) {real, imag} */,
  {32'h455fdccb, 32'h00000000} /* (28, 14, 15) {real, imag} */,
  {32'h453ccfc9, 32'h00000000} /* (28, 14, 14) {real, imag} */,
  {32'h456f7b4e, 32'h00000000} /* (28, 14, 13) {real, imag} */,
  {32'h45242d25, 32'h00000000} /* (28, 14, 12) {real, imag} */,
  {32'h447e50f2, 32'h00000000} /* (28, 14, 11) {real, imag} */,
  {32'hc3af8d94, 32'h00000000} /* (28, 14, 10) {real, imag} */,
  {32'hc51a5d5b, 32'h00000000} /* (28, 14, 9) {real, imag} */,
  {32'hc569a77b, 32'h00000000} /* (28, 14, 8) {real, imag} */,
  {32'hc5697566, 32'h00000000} /* (28, 14, 7) {real, imag} */,
  {32'hc553e080, 32'h00000000} /* (28, 14, 6) {real, imag} */,
  {32'hc545c2da, 32'h00000000} /* (28, 14, 5) {real, imag} */,
  {32'hc547f06c, 32'h00000000} /* (28, 14, 4) {real, imag} */,
  {32'hc57ccc48, 32'h00000000} /* (28, 14, 3) {real, imag} */,
  {32'hc56a71f6, 32'h00000000} /* (28, 14, 2) {real, imag} */,
  {32'hc57528d6, 32'h00000000} /* (28, 14, 1) {real, imag} */,
  {32'hc52c7543, 32'h00000000} /* (28, 14, 0) {real, imag} */,
  {32'hc53b00b8, 32'h00000000} /* (28, 13, 31) {real, imag} */,
  {32'hc5398001, 32'h00000000} /* (28, 13, 30) {real, imag} */,
  {32'hc566cdab, 32'h00000000} /* (28, 13, 29) {real, imag} */,
  {32'hc5468532, 32'h00000000} /* (28, 13, 28) {real, imag} */,
  {32'hc538cc79, 32'h00000000} /* (28, 13, 27) {real, imag} */,
  {32'hc5505d64, 32'h00000000} /* (28, 13, 26) {real, imag} */,
  {32'hc571f2e3, 32'h00000000} /* (28, 13, 25) {real, imag} */,
  {32'hc561c7d4, 32'h00000000} /* (28, 13, 24) {real, imag} */,
  {32'hc50c5332, 32'h00000000} /* (28, 13, 23) {real, imag} */,
  {32'hc4dac819, 32'h00000000} /* (28, 13, 22) {real, imag} */,
  {32'hc3df04c0, 32'h00000000} /* (28, 13, 21) {real, imag} */,
  {32'h44bb3008, 32'h00000000} /* (28, 13, 20) {real, imag} */,
  {32'h44f077f4, 32'h00000000} /* (28, 13, 19) {real, imag} */,
  {32'h4543f310, 32'h00000000} /* (28, 13, 18) {real, imag} */,
  {32'h454a518a, 32'h00000000} /* (28, 13, 17) {real, imag} */,
  {32'h4515825a, 32'h00000000} /* (28, 13, 16) {real, imag} */,
  {32'h455fae2c, 32'h00000000} /* (28, 13, 15) {real, imag} */,
  {32'h45427e73, 32'h00000000} /* (28, 13, 14) {real, imag} */,
  {32'h45210c87, 32'h00000000} /* (28, 13, 13) {real, imag} */,
  {32'h45095abe, 32'h00000000} /* (28, 13, 12) {real, imag} */,
  {32'h44395ff4, 32'h00000000} /* (28, 13, 11) {real, imag} */,
  {32'hc4ad6860, 32'h00000000} /* (28, 13, 10) {real, imag} */,
  {32'hc55f5231, 32'h00000000} /* (28, 13, 9) {real, imag} */,
  {32'hc542498c, 32'h00000000} /* (28, 13, 8) {real, imag} */,
  {32'hc52af616, 32'h00000000} /* (28, 13, 7) {real, imag} */,
  {32'hc525b198, 32'h00000000} /* (28, 13, 6) {real, imag} */,
  {32'hc51f6ba2, 32'h00000000} /* (28, 13, 5) {real, imag} */,
  {32'hc5274b52, 32'h00000000} /* (28, 13, 4) {real, imag} */,
  {32'hc541fa62, 32'h00000000} /* (28, 13, 3) {real, imag} */,
  {32'hc57a82e0, 32'h00000000} /* (28, 13, 2) {real, imag} */,
  {32'hc5542538, 32'h00000000} /* (28, 13, 1) {real, imag} */,
  {32'hc536c7ee, 32'h00000000} /* (28, 13, 0) {real, imag} */,
  {32'hc4de6989, 32'h00000000} /* (28, 12, 31) {real, imag} */,
  {32'hc562493e, 32'h00000000} /* (28, 12, 30) {real, imag} */,
  {32'hc53cc184, 32'h00000000} /* (28, 12, 29) {real, imag} */,
  {32'hc544f8bb, 32'h00000000} /* (28, 12, 28) {real, imag} */,
  {32'hc545c2ee, 32'h00000000} /* (28, 12, 27) {real, imag} */,
  {32'hc581b2e4, 32'h00000000} /* (28, 12, 26) {real, imag} */,
  {32'hc54843b9, 32'h00000000} /* (28, 12, 25) {real, imag} */,
  {32'hc5281782, 32'h00000000} /* (28, 12, 24) {real, imag} */,
  {32'hc50c6cbf, 32'h00000000} /* (28, 12, 23) {real, imag} */,
  {32'hc4da213b, 32'h00000000} /* (28, 12, 22) {real, imag} */,
  {32'hc44a0845, 32'h00000000} /* (28, 12, 21) {real, imag} */,
  {32'h44b9fd34, 32'h00000000} /* (28, 12, 20) {real, imag} */,
  {32'h44f647f9, 32'h00000000} /* (28, 12, 19) {real, imag} */,
  {32'h4536909a, 32'h00000000} /* (28, 12, 18) {real, imag} */,
  {32'h45181587, 32'h00000000} /* (28, 12, 17) {real, imag} */,
  {32'h450f61de, 32'h00000000} /* (28, 12, 16) {real, imag} */,
  {32'h44f201b3, 32'h00000000} /* (28, 12, 15) {real, imag} */,
  {32'h450cf6fe, 32'h00000000} /* (28, 12, 14) {real, imag} */,
  {32'h44f2701f, 32'h00000000} /* (28, 12, 13) {real, imag} */,
  {32'h44ae8ff6, 32'h00000000} /* (28, 12, 12) {real, imag} */,
  {32'h443c0c96, 32'h00000000} /* (28, 12, 11) {real, imag} */,
  {32'hc463e920, 32'h00000000} /* (28, 12, 10) {real, imag} */,
  {32'hc4faabde, 32'h00000000} /* (28, 12, 9) {real, imag} */,
  {32'hc52650d2, 32'h00000000} /* (28, 12, 8) {real, imag} */,
  {32'hc5173ad9, 32'h00000000} /* (28, 12, 7) {real, imag} */,
  {32'hc50f3720, 32'h00000000} /* (28, 12, 6) {real, imag} */,
  {32'hc51a32c6, 32'h00000000} /* (28, 12, 5) {real, imag} */,
  {32'hc52df86a, 32'h00000000} /* (28, 12, 4) {real, imag} */,
  {32'hc575ca02, 32'h00000000} /* (28, 12, 3) {real, imag} */,
  {32'hc5525a26, 32'h00000000} /* (28, 12, 2) {real, imag} */,
  {32'hc582d099, 32'h00000000} /* (28, 12, 1) {real, imag} */,
  {32'hc51f60ee, 32'h00000000} /* (28, 12, 0) {real, imag} */,
  {32'hc4b48a73, 32'h00000000} /* (28, 11, 31) {real, imag} */,
  {32'hc4a776a6, 32'h00000000} /* (28, 11, 30) {real, imag} */,
  {32'hc49e9f5a, 32'h00000000} /* (28, 11, 29) {real, imag} */,
  {32'hc4f2ae01, 32'h00000000} /* (28, 11, 28) {real, imag} */,
  {32'hc5227f09, 32'h00000000} /* (28, 11, 27) {real, imag} */,
  {32'hc5133981, 32'h00000000} /* (28, 11, 26) {real, imag} */,
  {32'hc4e510ef, 32'h00000000} /* (28, 11, 25) {real, imag} */,
  {32'hc50862fe, 32'h00000000} /* (28, 11, 24) {real, imag} */,
  {32'hc4d35394, 32'h00000000} /* (28, 11, 23) {real, imag} */,
  {32'hc4a04ee9, 32'h00000000} /* (28, 11, 22) {real, imag} */,
  {32'hc3e593a6, 32'h00000000} /* (28, 11, 21) {real, imag} */,
  {32'hc30ae120, 32'h00000000} /* (28, 11, 20) {real, imag} */,
  {32'h447da0b4, 32'h00000000} /* (28, 11, 19) {real, imag} */,
  {32'h444c2086, 32'h00000000} /* (28, 11, 18) {real, imag} */,
  {32'h44be8d60, 32'h00000000} /* (28, 11, 17) {real, imag} */,
  {32'h44965bbf, 32'h00000000} /* (28, 11, 16) {real, imag} */,
  {32'h4480687f, 32'h00000000} /* (28, 11, 15) {real, imag} */,
  {32'h44a0eef2, 32'h00000000} /* (28, 11, 14) {real, imag} */,
  {32'h44bea5c6, 32'h00000000} /* (28, 11, 13) {real, imag} */,
  {32'h43e6a8c4, 32'h00000000} /* (28, 11, 12) {real, imag} */,
  {32'h40e93200, 32'h00000000} /* (28, 11, 11) {real, imag} */,
  {32'hc4b9d714, 32'h00000000} /* (28, 11, 10) {real, imag} */,
  {32'hc46f6352, 32'h00000000} /* (28, 11, 9) {real, imag} */,
  {32'hc4a6017d, 32'h00000000} /* (28, 11, 8) {real, imag} */,
  {32'hc4f72d24, 32'h00000000} /* (28, 11, 7) {real, imag} */,
  {32'hc50caa78, 32'h00000000} /* (28, 11, 6) {real, imag} */,
  {32'hc50be1f9, 32'h00000000} /* (28, 11, 5) {real, imag} */,
  {32'hc4997a66, 32'h00000000} /* (28, 11, 4) {real, imag} */,
  {32'hc4bb465a, 32'h00000000} /* (28, 11, 3) {real, imag} */,
  {32'hc52c6a42, 32'h00000000} /* (28, 11, 2) {real, imag} */,
  {32'hc4ec1a22, 32'h00000000} /* (28, 11, 1) {real, imag} */,
  {32'hc4b6676d, 32'h00000000} /* (28, 11, 0) {real, imag} */,
  {32'h4422ef4a, 32'h00000000} /* (28, 10, 31) {real, imag} */,
  {32'h44046bb3, 32'h00000000} /* (28, 10, 30) {real, imag} */,
  {32'h42d39fa0, 32'h00000000} /* (28, 10, 29) {real, imag} */,
  {32'h42f85a30, 32'h00000000} /* (28, 10, 28) {real, imag} */,
  {32'h422ee790, 32'h00000000} /* (28, 10, 27) {real, imag} */,
  {32'hc369be7c, 32'h00000000} /* (28, 10, 26) {real, imag} */,
  {32'h44089b6a, 32'h00000000} /* (28, 10, 25) {real, imag} */,
  {32'h44e4917c, 32'h00000000} /* (28, 10, 24) {real, imag} */,
  {32'h448d32fa, 32'h00000000} /* (28, 10, 23) {real, imag} */,
  {32'h44b59c6d, 32'h00000000} /* (28, 10, 22) {real, imag} */,
  {32'h42957190, 32'h00000000} /* (28, 10, 21) {real, imag} */,
  {32'hc4e477dc, 32'h00000000} /* (28, 10, 20) {real, imag} */,
  {32'hc490dbe3, 32'h00000000} /* (28, 10, 19) {real, imag} */,
  {32'hc4837b91, 32'h00000000} /* (28, 10, 18) {real, imag} */,
  {32'hc4ebf506, 32'h00000000} /* (28, 10, 17) {real, imag} */,
  {32'hc43297df, 32'h00000000} /* (28, 10, 16) {real, imag} */,
  {32'hc4290856, 32'h00000000} /* (28, 10, 15) {real, imag} */,
  {32'hc4b4e9de, 32'h00000000} /* (28, 10, 14) {real, imag} */,
  {32'hc4198e12, 32'h00000000} /* (28, 10, 13) {real, imag} */,
  {32'hc4d7f260, 32'h00000000} /* (28, 10, 12) {real, imag} */,
  {32'hc4b9d666, 32'h00000000} /* (28, 10, 11) {real, imag} */,
  {32'hc34f2970, 32'h00000000} /* (28, 10, 10) {real, imag} */,
  {32'h43951d16, 32'h00000000} /* (28, 10, 9) {real, imag} */,
  {32'h440832c1, 32'h00000000} /* (28, 10, 8) {real, imag} */,
  {32'h43b1db72, 32'h00000000} /* (28, 10, 7) {real, imag} */,
  {32'h43b0ddac, 32'h00000000} /* (28, 10, 6) {real, imag} */,
  {32'h4487a854, 32'h00000000} /* (28, 10, 5) {real, imag} */,
  {32'h43d32f0e, 32'h00000000} /* (28, 10, 4) {real, imag} */,
  {32'h4310d966, 32'h00000000} /* (28, 10, 3) {real, imag} */,
  {32'h43563c22, 32'h00000000} /* (28, 10, 2) {real, imag} */,
  {32'h43787d60, 32'h00000000} /* (28, 10, 1) {real, imag} */,
  {32'h43aa388a, 32'h00000000} /* (28, 10, 0) {real, imag} */,
  {32'h45107109, 32'h00000000} /* (28, 9, 31) {real, imag} */,
  {32'h450be28d, 32'h00000000} /* (28, 9, 30) {real, imag} */,
  {32'h44db4980, 32'h00000000} /* (28, 9, 29) {real, imag} */,
  {32'h44b03a41, 32'h00000000} /* (28, 9, 28) {real, imag} */,
  {32'h44d48b9c, 32'h00000000} /* (28, 9, 27) {real, imag} */,
  {32'h4484c498, 32'h00000000} /* (28, 9, 26) {real, imag} */,
  {32'h451643a1, 32'h00000000} /* (28, 9, 25) {real, imag} */,
  {32'h452a84b2, 32'h00000000} /* (28, 9, 24) {real, imag} */,
  {32'h44f6636a, 32'h00000000} /* (28, 9, 23) {real, imag} */,
  {32'h45071ec0, 32'h00000000} /* (28, 9, 22) {real, imag} */,
  {32'h448352d8, 32'h00000000} /* (28, 9, 21) {real, imag} */,
  {32'hc4d69dee, 32'h00000000} /* (28, 9, 20) {real, imag} */,
  {32'hc5107411, 32'h00000000} /* (28, 9, 19) {real, imag} */,
  {32'hc50e5dba, 32'h00000000} /* (28, 9, 18) {real, imag} */,
  {32'hc56f537a, 32'h00000000} /* (28, 9, 17) {real, imag} */,
  {32'hc532386e, 32'h00000000} /* (28, 9, 16) {real, imag} */,
  {32'hc508e245, 32'h00000000} /* (28, 9, 15) {real, imag} */,
  {32'hc50845e7, 32'h00000000} /* (28, 9, 14) {real, imag} */,
  {32'hc4ed9c66, 32'h00000000} /* (28, 9, 13) {real, imag} */,
  {32'hc5145ada, 32'h00000000} /* (28, 9, 12) {real, imag} */,
  {32'hc4dea23a, 32'h00000000} /* (28, 9, 11) {real, imag} */,
  {32'h44049828, 32'h00000000} /* (28, 9, 10) {real, imag} */,
  {32'h4504508b, 32'h00000000} /* (28, 9, 9) {real, imag} */,
  {32'h44b20ea5, 32'h00000000} /* (28, 9, 8) {real, imag} */,
  {32'h44d20e2e, 32'h00000000} /* (28, 9, 7) {real, imag} */,
  {32'h44d25700, 32'h00000000} /* (28, 9, 6) {real, imag} */,
  {32'h44d5ea64, 32'h00000000} /* (28, 9, 5) {real, imag} */,
  {32'h452d4307, 32'h00000000} /* (28, 9, 4) {real, imag} */,
  {32'h45186beb, 32'h00000000} /* (28, 9, 3) {real, imag} */,
  {32'h44e564cc, 32'h00000000} /* (28, 9, 2) {real, imag} */,
  {32'h44b719f9, 32'h00000000} /* (28, 9, 1) {real, imag} */,
  {32'h44a7e00d, 32'h00000000} /* (28, 9, 0) {real, imag} */,
  {32'h4514eea6, 32'h00000000} /* (28, 8, 31) {real, imag} */,
  {32'h44ebbbbc, 32'h00000000} /* (28, 8, 30) {real, imag} */,
  {32'h45154eb3, 32'h00000000} /* (28, 8, 29) {real, imag} */,
  {32'h44b59c14, 32'h00000000} /* (28, 8, 28) {real, imag} */,
  {32'h44c44083, 32'h00000000} /* (28, 8, 27) {real, imag} */,
  {32'h452ce2f4, 32'h00000000} /* (28, 8, 26) {real, imag} */,
  {32'h44dd5634, 32'h00000000} /* (28, 8, 25) {real, imag} */,
  {32'h44fba33e, 32'h00000000} /* (28, 8, 24) {real, imag} */,
  {32'h4501e61f, 32'h00000000} /* (28, 8, 23) {real, imag} */,
  {32'h4504b56a, 32'h00000000} /* (28, 8, 22) {real, imag} */,
  {32'h44469f82, 32'h00000000} /* (28, 8, 21) {real, imag} */,
  {32'hc43637b1, 32'h00000000} /* (28, 8, 20) {real, imag} */,
  {32'hc4e567a6, 32'h00000000} /* (28, 8, 19) {real, imag} */,
  {32'hc57974f7, 32'h00000000} /* (28, 8, 18) {real, imag} */,
  {32'hc562bfd3, 32'h00000000} /* (28, 8, 17) {real, imag} */,
  {32'hc53da8e4, 32'h00000000} /* (28, 8, 16) {real, imag} */,
  {32'hc5238c42, 32'h00000000} /* (28, 8, 15) {real, imag} */,
  {32'hc5599482, 32'h00000000} /* (28, 8, 14) {real, imag} */,
  {32'hc55b03e1, 32'h00000000} /* (28, 8, 13) {real, imag} */,
  {32'hc51de3e6, 32'h00000000} /* (28, 8, 12) {real, imag} */,
  {32'hc51a5e74, 32'h00000000} /* (28, 8, 11) {real, imag} */,
  {32'h43c276c0, 32'h00000000} /* (28, 8, 10) {real, imag} */,
  {32'h44b4d77c, 32'h00000000} /* (28, 8, 9) {real, imag} */,
  {32'h44a7197c, 32'h00000000} /* (28, 8, 8) {real, imag} */,
  {32'h45026ea5, 32'h00000000} /* (28, 8, 7) {real, imag} */,
  {32'h44ff5bb1, 32'h00000000} /* (28, 8, 6) {real, imag} */,
  {32'h45095c5a, 32'h00000000} /* (28, 8, 5) {real, imag} */,
  {32'h45104f9d, 32'h00000000} /* (28, 8, 4) {real, imag} */,
  {32'h452b5c89, 32'h00000000} /* (28, 8, 3) {real, imag} */,
  {32'h45386477, 32'h00000000} /* (28, 8, 2) {real, imag} */,
  {32'h453dcb91, 32'h00000000} /* (28, 8, 1) {real, imag} */,
  {32'h44fd1a31, 32'h00000000} /* (28, 8, 0) {real, imag} */,
  {32'h44d950a2, 32'h00000000} /* (28, 7, 31) {real, imag} */,
  {32'h450a1510, 32'h00000000} /* (28, 7, 30) {real, imag} */,
  {32'h44d32900, 32'h00000000} /* (28, 7, 29) {real, imag} */,
  {32'h44aca5bc, 32'h00000000} /* (28, 7, 28) {real, imag} */,
  {32'h44e26927, 32'h00000000} /* (28, 7, 27) {real, imag} */,
  {32'h45165486, 32'h00000000} /* (28, 7, 26) {real, imag} */,
  {32'h45304c63, 32'h00000000} /* (28, 7, 25) {real, imag} */,
  {32'h456550aa, 32'h00000000} /* (28, 7, 24) {real, imag} */,
  {32'h45057bfa, 32'h00000000} /* (28, 7, 23) {real, imag} */,
  {32'h44d208a4, 32'h00000000} /* (28, 7, 22) {real, imag} */,
  {32'h44ad2664, 32'h00000000} /* (28, 7, 21) {real, imag} */,
  {32'hc4c1e240, 32'h00000000} /* (28, 7, 20) {real, imag} */,
  {32'hc53610de, 32'h00000000} /* (28, 7, 19) {real, imag} */,
  {32'hc50e29cc, 32'h00000000} /* (28, 7, 18) {real, imag} */,
  {32'hc562ee12, 32'h00000000} /* (28, 7, 17) {real, imag} */,
  {32'hc52d27a5, 32'h00000000} /* (28, 7, 16) {real, imag} */,
  {32'hc584315e, 32'h00000000} /* (28, 7, 15) {real, imag} */,
  {32'hc5576682, 32'h00000000} /* (28, 7, 14) {real, imag} */,
  {32'hc555ff36, 32'h00000000} /* (28, 7, 13) {real, imag} */,
  {32'hc54394d0, 32'h00000000} /* (28, 7, 12) {real, imag} */,
  {32'hc4fc591d, 32'h00000000} /* (28, 7, 11) {real, imag} */,
  {32'hc46a9a73, 32'h00000000} /* (28, 7, 10) {real, imag} */,
  {32'h44111460, 32'h00000000} /* (28, 7, 9) {real, imag} */,
  {32'h44eb24bd, 32'h00000000} /* (28, 7, 8) {real, imag} */,
  {32'h44ecc620, 32'h00000000} /* (28, 7, 7) {real, imag} */,
  {32'h44edeb7a, 32'h00000000} /* (28, 7, 6) {real, imag} */,
  {32'h4540e324, 32'h00000000} /* (28, 7, 5) {real, imag} */,
  {32'h454fc68e, 32'h00000000} /* (28, 7, 4) {real, imag} */,
  {32'h454a55b6, 32'h00000000} /* (28, 7, 3) {real, imag} */,
  {32'h455471f8, 32'h00000000} /* (28, 7, 2) {real, imag} */,
  {32'h451e4b82, 32'h00000000} /* (28, 7, 1) {real, imag} */,
  {32'h44d7d066, 32'h00000000} /* (28, 7, 0) {real, imag} */,
  {32'h44e8864c, 32'h00000000} /* (28, 6, 31) {real, imag} */,
  {32'h44c06b8e, 32'h00000000} /* (28, 6, 30) {real, imag} */,
  {32'h44fb4b1e, 32'h00000000} /* (28, 6, 29) {real, imag} */,
  {32'h44ebb278, 32'h00000000} /* (28, 6, 28) {real, imag} */,
  {32'h4514452c, 32'h00000000} /* (28, 6, 27) {real, imag} */,
  {32'h45468cb6, 32'h00000000} /* (28, 6, 26) {real, imag} */,
  {32'h4543d53c, 32'h00000000} /* (28, 6, 25) {real, imag} */,
  {32'h450192b3, 32'h00000000} /* (28, 6, 24) {real, imag} */,
  {32'h451ec7a8, 32'h00000000} /* (28, 6, 23) {real, imag} */,
  {32'h453dc027, 32'h00000000} /* (28, 6, 22) {real, imag} */,
  {32'h44e17ffb, 32'h00000000} /* (28, 6, 21) {real, imag} */,
  {32'hc3889368, 32'h00000000} /* (28, 6, 20) {real, imag} */,
  {32'hc4dc65c0, 32'h00000000} /* (28, 6, 19) {real, imag} */,
  {32'hc50c7122, 32'h00000000} /* (28, 6, 18) {real, imag} */,
  {32'hc505f786, 32'h00000000} /* (28, 6, 17) {real, imag} */,
  {32'hc52399c4, 32'h00000000} /* (28, 6, 16) {real, imag} */,
  {32'hc54b281e, 32'h00000000} /* (28, 6, 15) {real, imag} */,
  {32'hc5705c61, 32'h00000000} /* (28, 6, 14) {real, imag} */,
  {32'hc5741b2d, 32'h00000000} /* (28, 6, 13) {real, imag} */,
  {32'hc56151fa, 32'h00000000} /* (28, 6, 12) {real, imag} */,
  {32'hc50d05ae, 32'h00000000} /* (28, 6, 11) {real, imag} */,
  {32'hc4442dc2, 32'h00000000} /* (28, 6, 10) {real, imag} */,
  {32'h439d7560, 32'h00000000} /* (28, 6, 9) {real, imag} */,
  {32'h447e1264, 32'h00000000} /* (28, 6, 8) {real, imag} */,
  {32'h44aa79a8, 32'h00000000} /* (28, 6, 7) {real, imag} */,
  {32'h44e3a902, 32'h00000000} /* (28, 6, 6) {real, imag} */,
  {32'h4526d43a, 32'h00000000} /* (28, 6, 5) {real, imag} */,
  {32'h459502a8, 32'h00000000} /* (28, 6, 4) {real, imag} */,
  {32'h4558cbf4, 32'h00000000} /* (28, 6, 3) {real, imag} */,
  {32'h451423e2, 32'h00000000} /* (28, 6, 2) {real, imag} */,
  {32'h44e2e3b8, 32'h00000000} /* (28, 6, 1) {real, imag} */,
  {32'h44c264c8, 32'h00000000} /* (28, 6, 0) {real, imag} */,
  {32'h44b1888a, 32'h00000000} /* (28, 5, 31) {real, imag} */,
  {32'h44df3d92, 32'h00000000} /* (28, 5, 30) {real, imag} */,
  {32'h44fc75a9, 32'h00000000} /* (28, 5, 29) {real, imag} */,
  {32'h45058d5b, 32'h00000000} /* (28, 5, 28) {real, imag} */,
  {32'h453284ca, 32'h00000000} /* (28, 5, 27) {real, imag} */,
  {32'h452badee, 32'h00000000} /* (28, 5, 26) {real, imag} */,
  {32'h452e8468, 32'h00000000} /* (28, 5, 25) {real, imag} */,
  {32'h4541efea, 32'h00000000} /* (28, 5, 24) {real, imag} */,
  {32'h45422aa5, 32'h00000000} /* (28, 5, 23) {real, imag} */,
  {32'h452345d6, 32'h00000000} /* (28, 5, 22) {real, imag} */,
  {32'h4548527a, 32'h00000000} /* (28, 5, 21) {real, imag} */,
  {32'h450c8ce1, 32'h00000000} /* (28, 5, 20) {real, imag} */,
  {32'h445a742e, 32'h00000000} /* (28, 5, 19) {real, imag} */,
  {32'h438299d4, 32'h00000000} /* (28, 5, 18) {real, imag} */,
  {32'hc4157fd1, 32'h00000000} /* (28, 5, 17) {real, imag} */,
  {32'hc4b40600, 32'h00000000} /* (28, 5, 16) {real, imag} */,
  {32'hc4ec4142, 32'h00000000} /* (28, 5, 15) {real, imag} */,
  {32'hc545c209, 32'h00000000} /* (28, 5, 14) {real, imag} */,
  {32'hc57ba5fe, 32'h00000000} /* (28, 5, 13) {real, imag} */,
  {32'hc53f3413, 32'h00000000} /* (28, 5, 12) {real, imag} */,
  {32'hc568b310, 32'h00000000} /* (28, 5, 11) {real, imag} */,
  {32'hc52c1dde, 32'h00000000} /* (28, 5, 10) {real, imag} */,
  {32'hc48ddaca, 32'h00000000} /* (28, 5, 9) {real, imag} */,
  {32'hc401da96, 32'h00000000} /* (28, 5, 8) {real, imag} */,
  {32'hc3faa1d8, 32'h00000000} /* (28, 5, 7) {real, imag} */,
  {32'h43cf0150, 32'h00000000} /* (28, 5, 6) {real, imag} */,
  {32'h4528f4ae, 32'h00000000} /* (28, 5, 5) {real, imag} */,
  {32'h452c594b, 32'h00000000} /* (28, 5, 4) {real, imag} */,
  {32'h4545d9fc, 32'h00000000} /* (28, 5, 3) {real, imag} */,
  {32'h4511329c, 32'h00000000} /* (28, 5, 2) {real, imag} */,
  {32'h44fd88c8, 32'h00000000} /* (28, 5, 1) {real, imag} */,
  {32'h44d30dc2, 32'h00000000} /* (28, 5, 0) {real, imag} */,
  {32'h44a61d5a, 32'h00000000} /* (28, 4, 31) {real, imag} */,
  {32'h44e43c67, 32'h00000000} /* (28, 4, 30) {real, imag} */,
  {32'h4505393a, 32'h00000000} /* (28, 4, 29) {real, imag} */,
  {32'h44fedee7, 32'h00000000} /* (28, 4, 28) {real, imag} */,
  {32'h44cc0ed8, 32'h00000000} /* (28, 4, 27) {real, imag} */,
  {32'h4455d102, 32'h00000000} /* (28, 4, 26) {real, imag} */,
  {32'h4428df32, 32'h00000000} /* (28, 4, 25) {real, imag} */,
  {32'h45173be0, 32'h00000000} /* (28, 4, 24) {real, imag} */,
  {32'h451dc2ee, 32'h00000000} /* (28, 4, 23) {real, imag} */,
  {32'h450deb64, 32'h00000000} /* (28, 4, 22) {real, imag} */,
  {32'h453c38ce, 32'h00000000} /* (28, 4, 21) {real, imag} */,
  {32'h44efd665, 32'h00000000} /* (28, 4, 20) {real, imag} */,
  {32'h450538ea, 32'h00000000} /* (28, 4, 19) {real, imag} */,
  {32'h45098ef7, 32'h00000000} /* (28, 4, 18) {real, imag} */,
  {32'h44c894fe, 32'h00000000} /* (28, 4, 17) {real, imag} */,
  {32'h43284bf4, 32'h00000000} /* (28, 4, 16) {real, imag} */,
  {32'hc5039a00, 32'h00000000} /* (28, 4, 15) {real, imag} */,
  {32'hc52262ba, 32'h00000000} /* (28, 4, 14) {real, imag} */,
  {32'hc5576104, 32'h00000000} /* (28, 4, 13) {real, imag} */,
  {32'hc5325ca6, 32'h00000000} /* (28, 4, 12) {real, imag} */,
  {32'hc5505acc, 32'h00000000} /* (28, 4, 11) {real, imag} */,
  {32'hc55378fc, 32'h00000000} /* (28, 4, 10) {real, imag} */,
  {32'hc5037248, 32'h00000000} /* (28, 4, 9) {real, imag} */,
  {32'hc508cdae, 32'h00000000} /* (28, 4, 8) {real, imag} */,
  {32'hc4cdb031, 32'h00000000} /* (28, 4, 7) {real, imag} */,
  {32'hc4805b90, 32'h00000000} /* (28, 4, 6) {real, imag} */,
  {32'h4497727c, 32'h00000000} /* (28, 4, 5) {real, imag} */,
  {32'h44fd8411, 32'h00000000} /* (28, 4, 4) {real, imag} */,
  {32'h4514d904, 32'h00000000} /* (28, 4, 3) {real, imag} */,
  {32'h4534d005, 32'h00000000} /* (28, 4, 2) {real, imag} */,
  {32'h44aeb57c, 32'h00000000} /* (28, 4, 1) {real, imag} */,
  {32'h4483d14e, 32'h00000000} /* (28, 4, 0) {real, imag} */,
  {32'h448f9e32, 32'h00000000} /* (28, 3, 31) {real, imag} */,
  {32'h44cd607e, 32'h00000000} /* (28, 3, 30) {real, imag} */,
  {32'h45008199, 32'h00000000} /* (28, 3, 29) {real, imag} */,
  {32'h454393a0, 32'h00000000} /* (28, 3, 28) {real, imag} */,
  {32'h451cf182, 32'h00000000} /* (28, 3, 27) {real, imag} */,
  {32'h44cb27ef, 32'h00000000} /* (28, 3, 26) {real, imag} */,
  {32'h448a0030, 32'h00000000} /* (28, 3, 25) {real, imag} */,
  {32'h448ee032, 32'h00000000} /* (28, 3, 24) {real, imag} */,
  {32'h45013bc1, 32'h00000000} /* (28, 3, 23) {real, imag} */,
  {32'h45179dfd, 32'h00000000} /* (28, 3, 22) {real, imag} */,
  {32'h4516c6c1, 32'h00000000} /* (28, 3, 21) {real, imag} */,
  {32'h453f04ea, 32'h00000000} /* (28, 3, 20) {real, imag} */,
  {32'h4513aa5e, 32'h00000000} /* (28, 3, 19) {real, imag} */,
  {32'h451a2182, 32'h00000000} /* (28, 3, 18) {real, imag} */,
  {32'h450ba4ac, 32'h00000000} /* (28, 3, 17) {real, imag} */,
  {32'h44abf65c, 32'h00000000} /* (28, 3, 16) {real, imag} */,
  {32'hc4bf4706, 32'h00000000} /* (28, 3, 15) {real, imag} */,
  {32'hc5242d49, 32'h00000000} /* (28, 3, 14) {real, imag} */,
  {32'hc54de523, 32'h00000000} /* (28, 3, 13) {real, imag} */,
  {32'hc56b21e6, 32'h00000000} /* (28, 3, 12) {real, imag} */,
  {32'hc5350ee8, 32'h00000000} /* (28, 3, 11) {real, imag} */,
  {32'hc5494cbc, 32'h00000000} /* (28, 3, 10) {real, imag} */,
  {32'hc53eed62, 32'h00000000} /* (28, 3, 9) {real, imag} */,
  {32'hc51d7f2c, 32'h00000000} /* (28, 3, 8) {real, imag} */,
  {32'hc4ba61b3, 32'h00000000} /* (28, 3, 7) {real, imag} */,
  {32'hc50503d1, 32'h00000000} /* (28, 3, 6) {real, imag} */,
  {32'hc4253f45, 32'h00000000} /* (28, 3, 5) {real, imag} */,
  {32'h4480776f, 32'h00000000} /* (28, 3, 4) {real, imag} */,
  {32'h45100dfe, 32'h00000000} /* (28, 3, 3) {real, imag} */,
  {32'h4547a902, 32'h00000000} /* (28, 3, 2) {real, imag} */,
  {32'h4502f1f8, 32'h00000000} /* (28, 3, 1) {real, imag} */,
  {32'h4483deae, 32'h00000000} /* (28, 3, 0) {real, imag} */,
  {32'h4454c6e2, 32'h00000000} /* (28, 2, 31) {real, imag} */,
  {32'h44e41aba, 32'h00000000} /* (28, 2, 30) {real, imag} */,
  {32'h44b7da00, 32'h00000000} /* (28, 2, 29) {real, imag} */,
  {32'h44b07d57, 32'h00000000} /* (28, 2, 28) {real, imag} */,
  {32'h450658bc, 32'h00000000} /* (28, 2, 27) {real, imag} */,
  {32'h44cf4b60, 32'h00000000} /* (28, 2, 26) {real, imag} */,
  {32'h44df6c2a, 32'h00000000} /* (28, 2, 25) {real, imag} */,
  {32'h453d58e4, 32'h00000000} /* (28, 2, 24) {real, imag} */,
  {32'h452b0018, 32'h00000000} /* (28, 2, 23) {real, imag} */,
  {32'h45326738, 32'h00000000} /* (28, 2, 22) {real, imag} */,
  {32'h4523d0a2, 32'h00000000} /* (28, 2, 21) {real, imag} */,
  {32'h456e1916, 32'h00000000} /* (28, 2, 20) {real, imag} */,
  {32'h452f13c8, 32'h00000000} /* (28, 2, 19) {real, imag} */,
  {32'h44cba59c, 32'h00000000} /* (28, 2, 18) {real, imag} */,
  {32'h44adafe4, 32'h00000000} /* (28, 2, 17) {real, imag} */,
  {32'h447d0b54, 32'h00000000} /* (28, 2, 16) {real, imag} */,
  {32'hc50adf52, 32'h00000000} /* (28, 2, 15) {real, imag} */,
  {32'hc5318a3f, 32'h00000000} /* (28, 2, 14) {real, imag} */,
  {32'hc55b8516, 32'h00000000} /* (28, 2, 13) {real, imag} */,
  {32'hc54462d8, 32'h00000000} /* (28, 2, 12) {real, imag} */,
  {32'hc531650e, 32'h00000000} /* (28, 2, 11) {real, imag} */,
  {32'hc58eb077, 32'h00000000} /* (28, 2, 10) {real, imag} */,
  {32'hc5a188fa, 32'h00000000} /* (28, 2, 9) {real, imag} */,
  {32'hc536e768, 32'h00000000} /* (28, 2, 8) {real, imag} */,
  {32'hc50e256e, 32'h00000000} /* (28, 2, 7) {real, imag} */,
  {32'hc500e168, 32'h00000000} /* (28, 2, 6) {real, imag} */,
  {32'hc453c8b1, 32'h00000000} /* (28, 2, 5) {real, imag} */,
  {32'h4413a83a, 32'h00000000} /* (28, 2, 4) {real, imag} */,
  {32'h4507db1e, 32'h00000000} /* (28, 2, 3) {real, imag} */,
  {32'h44e37384, 32'h00000000} /* (28, 2, 2) {real, imag} */,
  {32'h44d75dc0, 32'h00000000} /* (28, 2, 1) {real, imag} */,
  {32'h449c0752, 32'h00000000} /* (28, 2, 0) {real, imag} */,
  {32'h4456c1cf, 32'h00000000} /* (28, 1, 31) {real, imag} */,
  {32'h44294db4, 32'h00000000} /* (28, 1, 30) {real, imag} */,
  {32'h44a46ccd, 32'h00000000} /* (28, 1, 29) {real, imag} */,
  {32'h442b46d2, 32'h00000000} /* (28, 1, 28) {real, imag} */,
  {32'h448cd924, 32'h00000000} /* (28, 1, 27) {real, imag} */,
  {32'h44802fe4, 32'h00000000} /* (28, 1, 26) {real, imag} */,
  {32'h4494aa75, 32'h00000000} /* (28, 1, 25) {real, imag} */,
  {32'h4520e8bb, 32'h00000000} /* (28, 1, 24) {real, imag} */,
  {32'h4563abf1, 32'h00000000} /* (28, 1, 23) {real, imag} */,
  {32'h454eeb4c, 32'h00000000} /* (28, 1, 22) {real, imag} */,
  {32'h454f90f2, 32'h00000000} /* (28, 1, 21) {real, imag} */,
  {32'h45060802, 32'h00000000} /* (28, 1, 20) {real, imag} */,
  {32'h4523c924, 32'h00000000} /* (28, 1, 19) {real, imag} */,
  {32'h453768c6, 32'h00000000} /* (28, 1, 18) {real, imag} */,
  {32'h4513a61f, 32'h00000000} /* (28, 1, 17) {real, imag} */,
  {32'h449f3341, 32'h00000000} /* (28, 1, 16) {real, imag} */,
  {32'hc4c591b8, 32'h00000000} /* (28, 1, 15) {real, imag} */,
  {32'hc51901f3, 32'h00000000} /* (28, 1, 14) {real, imag} */,
  {32'hc5713b3e, 32'h00000000} /* (28, 1, 13) {real, imag} */,
  {32'hc56e77ba, 32'h00000000} /* (28, 1, 12) {real, imag} */,
  {32'hc52fcc38, 32'h00000000} /* (28, 1, 11) {real, imag} */,
  {32'hc58a1a50, 32'h00000000} /* (28, 1, 10) {real, imag} */,
  {32'hc58923c2, 32'h00000000} /* (28, 1, 9) {real, imag} */,
  {32'hc50a5923, 32'h00000000} /* (28, 1, 8) {real, imag} */,
  {32'hc512f76d, 32'h00000000} /* (28, 1, 7) {real, imag} */,
  {32'hc4bc580b, 32'h00000000} /* (28, 1, 6) {real, imag} */,
  {32'hc40974b6, 32'h00000000} /* (28, 1, 5) {real, imag} */,
  {32'h446003bd, 32'h00000000} /* (28, 1, 4) {real, imag} */,
  {32'h44c1d708, 32'h00000000} /* (28, 1, 3) {real, imag} */,
  {32'h44c7b883, 32'h00000000} /* (28, 1, 2) {real, imag} */,
  {32'h448d4400, 32'h00000000} /* (28, 1, 1) {real, imag} */,
  {32'h4414b6e8, 32'h00000000} /* (28, 1, 0) {real, imag} */,
  {32'h42c39318, 32'h00000000} /* (28, 0, 31) {real, imag} */,
  {32'h43a1720c, 32'h00000000} /* (28, 0, 30) {real, imag} */,
  {32'h44073d8a, 32'h00000000} /* (28, 0, 29) {real, imag} */,
  {32'h4413304c, 32'h00000000} /* (28, 0, 28) {real, imag} */,
  {32'h440e435e, 32'h00000000} /* (28, 0, 27) {real, imag} */,
  {32'h440c260a, 32'h00000000} /* (28, 0, 26) {real, imag} */,
  {32'h44bc1110, 32'h00000000} /* (28, 0, 25) {real, imag} */,
  {32'h44e5f185, 32'h00000000} /* (28, 0, 24) {real, imag} */,
  {32'h44fdd86a, 32'h00000000} /* (28, 0, 23) {real, imag} */,
  {32'h44f5becc, 32'h00000000} /* (28, 0, 22) {real, imag} */,
  {32'h45061c12, 32'h00000000} /* (28, 0, 21) {real, imag} */,
  {32'h44dd34df, 32'h00000000} /* (28, 0, 20) {real, imag} */,
  {32'h44f168ec, 32'h00000000} /* (28, 0, 19) {real, imag} */,
  {32'h448d9009, 32'h00000000} /* (28, 0, 18) {real, imag} */,
  {32'h44418c67, 32'h00000000} /* (28, 0, 17) {real, imag} */,
  {32'h4246eb34, 32'h00000000} /* (28, 0, 16) {real, imag} */,
  {32'hc503f817, 32'h00000000} /* (28, 0, 15) {real, imag} */,
  {32'hc511dc8c, 32'h00000000} /* (28, 0, 14) {real, imag} */,
  {32'hc5301414, 32'h00000000} /* (28, 0, 13) {real, imag} */,
  {32'hc578ed35, 32'h00000000} /* (28, 0, 12) {real, imag} */,
  {32'hc54bba58, 32'h00000000} /* (28, 0, 11) {real, imag} */,
  {32'hc4d36a3f, 32'h00000000} /* (28, 0, 10) {real, imag} */,
  {32'hc4bc1584, 32'h00000000} /* (28, 0, 9) {real, imag} */,
  {32'hc49e34f9, 32'h00000000} /* (28, 0, 8) {real, imag} */,
  {32'hc4ab1d72, 32'h00000000} /* (28, 0, 7) {real, imag} */,
  {32'hc4660bb0, 32'h00000000} /* (28, 0, 6) {real, imag} */,
  {32'h42b2e110, 32'h00000000} /* (28, 0, 5) {real, imag} */,
  {32'h4464192a, 32'h00000000} /* (28, 0, 4) {real, imag} */,
  {32'h44770791, 32'h00000000} /* (28, 0, 3) {real, imag} */,
  {32'h448e280b, 32'h00000000} /* (28, 0, 2) {real, imag} */,
  {32'h442385f9, 32'h00000000} /* (28, 0, 1) {real, imag} */,
  {32'h43b37662, 32'h00000000} /* (28, 0, 0) {real, imag} */,
  {32'hc4caade2, 32'h00000000} /* (27, 31, 31) {real, imag} */,
  {32'hc4de8981, 32'h00000000} /* (27, 31, 30) {real, imag} */,
  {32'hc4dedc57, 32'h00000000} /* (27, 31, 29) {real, imag} */,
  {32'hc4425ca6, 32'h00000000} /* (27, 31, 28) {real, imag} */,
  {32'hc4048637, 32'h00000000} /* (27, 31, 27) {real, imag} */,
  {32'hc4025fd7, 32'h00000000} /* (27, 31, 26) {real, imag} */,
  {32'h441c6ae6, 32'h00000000} /* (27, 31, 25) {real, imag} */,
  {32'hc20b1d98, 32'h00000000} /* (27, 31, 24) {real, imag} */,
  {32'h42781ec8, 32'h00000000} /* (27, 31, 23) {real, imag} */,
  {32'hc2d772f0, 32'h00000000} /* (27, 31, 22) {real, imag} */,
  {32'hc35ae0c0, 32'h00000000} /* (27, 31, 21) {real, imag} */,
  {32'hc3d5bdb6, 32'h00000000} /* (27, 31, 20) {real, imag} */,
  {32'hc40138c4, 32'h00000000} /* (27, 31, 19) {real, imag} */,
  {32'hc3e511ac, 32'h00000000} /* (27, 31, 18) {real, imag} */,
  {32'hc3fd494c, 32'h00000000} /* (27, 31, 17) {real, imag} */,
  {32'hc43db676, 32'h00000000} /* (27, 31, 16) {real, imag} */,
  {32'hc494482e, 32'h00000000} /* (27, 31, 15) {real, imag} */,
  {32'hc50a470a, 32'h00000000} /* (27, 31, 14) {real, imag} */,
  {32'hc54a5edc, 32'h00000000} /* (27, 31, 13) {real, imag} */,
  {32'hc50c9ca4, 32'h00000000} /* (27, 31, 12) {real, imag} */,
  {32'hc4ed1782, 32'h00000000} /* (27, 31, 11) {real, imag} */,
  {32'hc431dc79, 32'h00000000} /* (27, 31, 10) {real, imag} */,
  {32'hc1e81760, 32'h00000000} /* (27, 31, 9) {real, imag} */,
  {32'h4390b49d, 32'h00000000} /* (27, 31, 8) {real, imag} */,
  {32'hc3ee52f1, 32'h00000000} /* (27, 31, 7) {real, imag} */,
  {32'h435c0628, 32'h00000000} /* (27, 31, 6) {real, imag} */,
  {32'h43ddeb58, 32'h00000000} /* (27, 31, 5) {real, imag} */,
  {32'h441d43eb, 32'h00000000} /* (27, 31, 4) {real, imag} */,
  {32'hc3d906b8, 32'h00000000} /* (27, 31, 3) {real, imag} */,
  {32'h441c0204, 32'h00000000} /* (27, 31, 2) {real, imag} */,
  {32'hc329cbd3, 32'h00000000} /* (27, 31, 1) {real, imag} */,
  {32'hc4bc1e4d, 32'h00000000} /* (27, 31, 0) {real, imag} */,
  {32'hc493d620, 32'h00000000} /* (27, 30, 31) {real, imag} */,
  {32'hc4b838db, 32'h00000000} /* (27, 30, 30) {real, imag} */,
  {32'hc4aca04c, 32'h00000000} /* (27, 30, 29) {real, imag} */,
  {32'h43e890c0, 32'h00000000} /* (27, 30, 28) {real, imag} */,
  {32'h43d7a69a, 32'h00000000} /* (27, 30, 27) {real, imag} */,
  {32'h42864248, 32'h00000000} /* (27, 30, 26) {real, imag} */,
  {32'h44b343c8, 32'h00000000} /* (27, 30, 25) {real, imag} */,
  {32'hc1639c20, 32'h00000000} /* (27, 30, 24) {real, imag} */,
  {32'h44b1b162, 32'h00000000} /* (27, 30, 23) {real, imag} */,
  {32'h4426a0a6, 32'h00000000} /* (27, 30, 22) {real, imag} */,
  {32'hc41e91a4, 32'h00000000} /* (27, 30, 21) {real, imag} */,
  {32'hc4aaed1a, 32'h00000000} /* (27, 30, 20) {real, imag} */,
  {32'hc503d15a, 32'h00000000} /* (27, 30, 19) {real, imag} */,
  {32'hc4c9b8e4, 32'h00000000} /* (27, 30, 18) {real, imag} */,
  {32'hc49584bc, 32'h00000000} /* (27, 30, 17) {real, imag} */,
  {32'hc513afc8, 32'h00000000} /* (27, 30, 16) {real, imag} */,
  {32'hc5112213, 32'h00000000} /* (27, 30, 15) {real, imag} */,
  {32'hc56857ca, 32'h00000000} /* (27, 30, 14) {real, imag} */,
  {32'hc5720eba, 32'h00000000} /* (27, 30, 13) {real, imag} */,
  {32'hc542f683, 32'h00000000} /* (27, 30, 12) {real, imag} */,
  {32'hc4f25d38, 32'h00000000} /* (27, 30, 11) {real, imag} */,
  {32'hc0478900, 32'h00000000} /* (27, 30, 10) {real, imag} */,
  {32'h44a2838c, 32'h00000000} /* (27, 30, 9) {real, imag} */,
  {32'h44467d3c, 32'h00000000} /* (27, 30, 8) {real, imag} */,
  {32'h4488f158, 32'h00000000} /* (27, 30, 7) {real, imag} */,
  {32'h43cfaf24, 32'h00000000} /* (27, 30, 6) {real, imag} */,
  {32'h449cedaa, 32'h00000000} /* (27, 30, 5) {real, imag} */,
  {32'h44abb014, 32'h00000000} /* (27, 30, 4) {real, imag} */,
  {32'h4460ec77, 32'h00000000} /* (27, 30, 3) {real, imag} */,
  {32'h442a5ec8, 32'h00000000} /* (27, 30, 2) {real, imag} */,
  {32'hc3f9739d, 32'h00000000} /* (27, 30, 1) {real, imag} */,
  {32'hc499073e, 32'h00000000} /* (27, 30, 0) {real, imag} */,
  {32'hc47e5b7d, 32'h00000000} /* (27, 29, 31) {real, imag} */,
  {32'hc426f8f6, 32'h00000000} /* (27, 29, 30) {real, imag} */,
  {32'hc3150ec8, 32'h00000000} /* (27, 29, 29) {real, imag} */,
  {32'h43dd5bc4, 32'h00000000} /* (27, 29, 28) {real, imag} */,
  {32'h443599bc, 32'h00000000} /* (27, 29, 27) {real, imag} */,
  {32'hc3ed027d, 32'h00000000} /* (27, 29, 26) {real, imag} */,
  {32'h443bc1f8, 32'h00000000} /* (27, 29, 25) {real, imag} */,
  {32'h447c8e46, 32'h00000000} /* (27, 29, 24) {real, imag} */,
  {32'h44349232, 32'h00000000} /* (27, 29, 23) {real, imag} */,
  {32'h43610d04, 32'h00000000} /* (27, 29, 22) {real, imag} */,
  {32'hc34599c0, 32'h00000000} /* (27, 29, 21) {real, imag} */,
  {32'hc4e44496, 32'h00000000} /* (27, 29, 20) {real, imag} */,
  {32'hc5224139, 32'h00000000} /* (27, 29, 19) {real, imag} */,
  {32'hc5487490, 32'h00000000} /* (27, 29, 18) {real, imag} */,
  {32'hc5137b08, 32'h00000000} /* (27, 29, 17) {real, imag} */,
  {32'hc533715c, 32'h00000000} /* (27, 29, 16) {real, imag} */,
  {32'hc537cbeb, 32'h00000000} /* (27, 29, 15) {real, imag} */,
  {32'hc555d9ae, 32'h00000000} /* (27, 29, 14) {real, imag} */,
  {32'hc519a33a, 32'h00000000} /* (27, 29, 13) {real, imag} */,
  {32'hc51ab450, 32'h00000000} /* (27, 29, 12) {real, imag} */,
  {32'hc4c4387e, 32'h00000000} /* (27, 29, 11) {real, imag} */,
  {32'h436ba2ca, 32'h00000000} /* (27, 29, 10) {real, imag} */,
  {32'h44ceba30, 32'h00000000} /* (27, 29, 9) {real, imag} */,
  {32'h44fc33b3, 32'h00000000} /* (27, 29, 8) {real, imag} */,
  {32'h44c4d95b, 32'h00000000} /* (27, 29, 7) {real, imag} */,
  {32'h4491ef5c, 32'h00000000} /* (27, 29, 6) {real, imag} */,
  {32'h44a8e46a, 32'h00000000} /* (27, 29, 5) {real, imag} */,
  {32'h450b1fd7, 32'h00000000} /* (27, 29, 4) {real, imag} */,
  {32'h45036587, 32'h00000000} /* (27, 29, 3) {real, imag} */,
  {32'hc1edc080, 32'h00000000} /* (27, 29, 2) {real, imag} */,
  {32'hc43a9e6a, 32'h00000000} /* (27, 29, 1) {real, imag} */,
  {32'hc48af712, 32'h00000000} /* (27, 29, 0) {real, imag} */,
  {32'hc43d9540, 32'h00000000} /* (27, 28, 31) {real, imag} */,
  {32'h43ca3fc4, 32'h00000000} /* (27, 28, 30) {real, imag} */,
  {32'hc35c0d50, 32'h00000000} /* (27, 28, 29) {real, imag} */,
  {32'hc3dcd3ba, 32'h00000000} /* (27, 28, 28) {real, imag} */,
  {32'h43f7888a, 32'h00000000} /* (27, 28, 27) {real, imag} */,
  {32'h440a6b23, 32'h00000000} /* (27, 28, 26) {real, imag} */,
  {32'hc3994a50, 32'h00000000} /* (27, 28, 25) {real, imag} */,
  {32'h448737bb, 32'h00000000} /* (27, 28, 24) {real, imag} */,
  {32'h444056ba, 32'h00000000} /* (27, 28, 23) {real, imag} */,
  {32'hc411e194, 32'h00000000} /* (27, 28, 22) {real, imag} */,
  {32'h43b60070, 32'h00000000} /* (27, 28, 21) {real, imag} */,
  {32'hc5123014, 32'h00000000} /* (27, 28, 20) {real, imag} */,
  {32'hc561243c, 32'h00000000} /* (27, 28, 19) {real, imag} */,
  {32'hc539fb18, 32'h00000000} /* (27, 28, 18) {real, imag} */,
  {32'hc52cbc04, 32'h00000000} /* (27, 28, 17) {real, imag} */,
  {32'hc54032de, 32'h00000000} /* (27, 28, 16) {real, imag} */,
  {32'hc5355924, 32'h00000000} /* (27, 28, 15) {real, imag} */,
  {32'hc530215a, 32'h00000000} /* (27, 28, 14) {real, imag} */,
  {32'hc5368ca5, 32'h00000000} /* (27, 28, 13) {real, imag} */,
  {32'hc5065c7f, 32'h00000000} /* (27, 28, 12) {real, imag} */,
  {32'hc48bab6c, 32'h00000000} /* (27, 28, 11) {real, imag} */,
  {32'h4466ae2d, 32'h00000000} /* (27, 28, 10) {real, imag} */,
  {32'h4541f4be, 32'h00000000} /* (27, 28, 9) {real, imag} */,
  {32'h45031d7f, 32'h00000000} /* (27, 28, 8) {real, imag} */,
  {32'h44ba7f2b, 32'h00000000} /* (27, 28, 7) {real, imag} */,
  {32'h44c61886, 32'h00000000} /* (27, 28, 6) {real, imag} */,
  {32'h4534adf8, 32'h00000000} /* (27, 28, 5) {real, imag} */,
  {32'h446d1fa6, 32'h00000000} /* (27, 28, 4) {real, imag} */,
  {32'h43df0d30, 32'h00000000} /* (27, 28, 3) {real, imag} */,
  {32'h448490dd, 32'h00000000} /* (27, 28, 2) {real, imag} */,
  {32'hc3a89374, 32'h00000000} /* (27, 28, 1) {real, imag} */,
  {32'hc41379a0, 32'h00000000} /* (27, 28, 0) {real, imag} */,
  {32'hc47e4b42, 32'h00000000} /* (27, 27, 31) {real, imag} */,
  {32'hc38b2b74, 32'h00000000} /* (27, 27, 30) {real, imag} */,
  {32'hc2b5a2c0, 32'h00000000} /* (27, 27, 29) {real, imag} */,
  {32'h44161200, 32'h00000000} /* (27, 27, 28) {real, imag} */,
  {32'h4435a17a, 32'h00000000} /* (27, 27, 27) {real, imag} */,
  {32'h4429efe8, 32'h00000000} /* (27, 27, 26) {real, imag} */,
  {32'h42263aa0, 32'h00000000} /* (27, 27, 25) {real, imag} */,
  {32'h42d0f5a0, 32'h00000000} /* (27, 27, 24) {real, imag} */,
  {32'h440b9424, 32'h00000000} /* (27, 27, 23) {real, imag} */,
  {32'h4403bea9, 32'h00000000} /* (27, 27, 22) {real, imag} */,
  {32'h4414290e, 32'h00000000} /* (27, 27, 21) {real, imag} */,
  {32'hc4c6eaad, 32'h00000000} /* (27, 27, 20) {real, imag} */,
  {32'hc5283690, 32'h00000000} /* (27, 27, 19) {real, imag} */,
  {32'hc557c98a, 32'h00000000} /* (27, 27, 18) {real, imag} */,
  {32'hc56850f4, 32'h00000000} /* (27, 27, 17) {real, imag} */,
  {32'hc555a2ba, 32'h00000000} /* (27, 27, 16) {real, imag} */,
  {32'hc53b5452, 32'h00000000} /* (27, 27, 15) {real, imag} */,
  {32'hc5118ee8, 32'h00000000} /* (27, 27, 14) {real, imag} */,
  {32'hc4f8965c, 32'h00000000} /* (27, 27, 13) {real, imag} */,
  {32'hc50d0078, 32'h00000000} /* (27, 27, 12) {real, imag} */,
  {32'hc4d4995f, 32'h00000000} /* (27, 27, 11) {real, imag} */,
  {32'h44268670, 32'h00000000} /* (27, 27, 10) {real, imag} */,
  {32'h450e6910, 32'h00000000} /* (27, 27, 9) {real, imag} */,
  {32'h45041853, 32'h00000000} /* (27, 27, 8) {real, imag} */,
  {32'h44e80ffe, 32'h00000000} /* (27, 27, 7) {real, imag} */,
  {32'h44f1c688, 32'h00000000} /* (27, 27, 6) {real, imag} */,
  {32'h44ef2079, 32'h00000000} /* (27, 27, 5) {real, imag} */,
  {32'h4491f425, 32'h00000000} /* (27, 27, 4) {real, imag} */,
  {32'h444dc696, 32'h00000000} /* (27, 27, 3) {real, imag} */,
  {32'h435e9be0, 32'h00000000} /* (27, 27, 2) {real, imag} */,
  {32'hc32b07c8, 32'h00000000} /* (27, 27, 1) {real, imag} */,
  {32'hc41aecf0, 32'h00000000} /* (27, 27, 0) {real, imag} */,
  {32'hc3f58af4, 32'h00000000} /* (27, 26, 31) {real, imag} */,
  {32'hc40b615c, 32'h00000000} /* (27, 26, 30) {real, imag} */,
  {32'hc3d44a00, 32'h00000000} /* (27, 26, 29) {real, imag} */,
  {32'hc37a9880, 32'h00000000} /* (27, 26, 28) {real, imag} */,
  {32'h42858e18, 32'h00000000} /* (27, 26, 27) {real, imag} */,
  {32'h44126d35, 32'h00000000} /* (27, 26, 26) {real, imag} */,
  {32'h443f5faa, 32'h00000000} /* (27, 26, 25) {real, imag} */,
  {32'h44225164, 32'h00000000} /* (27, 26, 24) {real, imag} */,
  {32'h4421ac3b, 32'h00000000} /* (27, 26, 23) {real, imag} */,
  {32'h447253a2, 32'h00000000} /* (27, 26, 22) {real, imag} */,
  {32'h428aabe0, 32'h00000000} /* (27, 26, 21) {real, imag} */,
  {32'hc4e2174e, 32'h00000000} /* (27, 26, 20) {real, imag} */,
  {32'hc501eaf7, 32'h00000000} /* (27, 26, 19) {real, imag} */,
  {32'hc568a716, 32'h00000000} /* (27, 26, 18) {real, imag} */,
  {32'hc5689880, 32'h00000000} /* (27, 26, 17) {real, imag} */,
  {32'hc52bd29e, 32'h00000000} /* (27, 26, 16) {real, imag} */,
  {32'hc57d27de, 32'h00000000} /* (27, 26, 15) {real, imag} */,
  {32'hc52208a4, 32'h00000000} /* (27, 26, 14) {real, imag} */,
  {32'hc52ceb24, 32'h00000000} /* (27, 26, 13) {real, imag} */,
  {32'hc51541c6, 32'h00000000} /* (27, 26, 12) {real, imag} */,
  {32'hc4e9baae, 32'h00000000} /* (27, 26, 11) {real, imag} */,
  {32'hc31242cc, 32'h00000000} /* (27, 26, 10) {real, imag} */,
  {32'h45009b52, 32'h00000000} /* (27, 26, 9) {real, imag} */,
  {32'h45041c12, 32'h00000000} /* (27, 26, 8) {real, imag} */,
  {32'h44d83e5c, 32'h00000000} /* (27, 26, 7) {real, imag} */,
  {32'h44c3d1f9, 32'h00000000} /* (27, 26, 6) {real, imag} */,
  {32'h44a2b6b2, 32'h00000000} /* (27, 26, 5) {real, imag} */,
  {32'h441fda43, 32'h00000000} /* (27, 26, 4) {real, imag} */,
  {32'h43d32ec8, 32'h00000000} /* (27, 26, 3) {real, imag} */,
  {32'h434348e0, 32'h00000000} /* (27, 26, 2) {real, imag} */,
  {32'h42cc5f40, 32'h00000000} /* (27, 26, 1) {real, imag} */,
  {32'hc462fccb, 32'h00000000} /* (27, 26, 0) {real, imag} */,
  {32'hc3eaf2b8, 32'h00000000} /* (27, 25, 31) {real, imag} */,
  {32'hc2b57460, 32'h00000000} /* (27, 25, 30) {real, imag} */,
  {32'hc3c1fa8a, 32'h00000000} /* (27, 25, 29) {real, imag} */,
  {32'hc42f8a49, 32'h00000000} /* (27, 25, 28) {real, imag} */,
  {32'h4399ca4e, 32'h00000000} /* (27, 25, 27) {real, imag} */,
  {32'h440c10a4, 32'h00000000} /* (27, 25, 26) {real, imag} */,
  {32'h43b0d36e, 32'h00000000} /* (27, 25, 25) {real, imag} */,
  {32'h44cb4b00, 32'h00000000} /* (27, 25, 24) {real, imag} */,
  {32'h4476c246, 32'h00000000} /* (27, 25, 23) {real, imag} */,
  {32'h444ba437, 32'h00000000} /* (27, 25, 22) {real, imag} */,
  {32'hc3cb7a78, 32'h00000000} /* (27, 25, 21) {real, imag} */,
  {32'hc4e32d18, 32'h00000000} /* (27, 25, 20) {real, imag} */,
  {32'hc4ca7873, 32'h00000000} /* (27, 25, 19) {real, imag} */,
  {32'hc50057b1, 32'h00000000} /* (27, 25, 18) {real, imag} */,
  {32'hc518f16a, 32'h00000000} /* (27, 25, 17) {real, imag} */,
  {32'hc4fcb212, 32'h00000000} /* (27, 25, 16) {real, imag} */,
  {32'hc53ce495, 32'h00000000} /* (27, 25, 15) {real, imag} */,
  {32'hc56144d0, 32'h00000000} /* (27, 25, 14) {real, imag} */,
  {32'hc4dd2b6e, 32'h00000000} /* (27, 25, 13) {real, imag} */,
  {32'hc511a81c, 32'h00000000} /* (27, 25, 12) {real, imag} */,
  {32'hc4b99548, 32'h00000000} /* (27, 25, 11) {real, imag} */,
  {32'hc2961540, 32'h00000000} /* (27, 25, 10) {real, imag} */,
  {32'h44aa6918, 32'h00000000} /* (27, 25, 9) {real, imag} */,
  {32'h4546428e, 32'h00000000} /* (27, 25, 8) {real, imag} */,
  {32'h45135de6, 32'h00000000} /* (27, 25, 7) {real, imag} */,
  {32'h44b25092, 32'h00000000} /* (27, 25, 6) {real, imag} */,
  {32'h4487b90a, 32'h00000000} /* (27, 25, 5) {real, imag} */,
  {32'h442a9440, 32'h00000000} /* (27, 25, 4) {real, imag} */,
  {32'hc2cb5410, 32'h00000000} /* (27, 25, 3) {real, imag} */,
  {32'h439945c8, 32'h00000000} /* (27, 25, 2) {real, imag} */,
  {32'hc44f3cf7, 32'h00000000} /* (27, 25, 1) {real, imag} */,
  {32'hc49cf19a, 32'h00000000} /* (27, 25, 0) {real, imag} */,
  {32'hc46758c6, 32'h00000000} /* (27, 24, 31) {real, imag} */,
  {32'h4307e1e8, 32'h00000000} /* (27, 24, 30) {real, imag} */,
  {32'h440474cf, 32'h00000000} /* (27, 24, 29) {real, imag} */,
  {32'h43ea123a, 32'h00000000} /* (27, 24, 28) {real, imag} */,
  {32'h449a4cba, 32'h00000000} /* (27, 24, 27) {real, imag} */,
  {32'h44c2d57f, 32'h00000000} /* (27, 24, 26) {real, imag} */,
  {32'h441bdb39, 32'h00000000} /* (27, 24, 25) {real, imag} */,
  {32'h446621b4, 32'h00000000} /* (27, 24, 24) {real, imag} */,
  {32'h4505cf33, 32'h00000000} /* (27, 24, 23) {real, imag} */,
  {32'h4469b08c, 32'h00000000} /* (27, 24, 22) {real, imag} */,
  {32'h44518f25, 32'h00000000} /* (27, 24, 21) {real, imag} */,
  {32'hc49f1d5e, 32'h00000000} /* (27, 24, 20) {real, imag} */,
  {32'hc506f626, 32'h00000000} /* (27, 24, 19) {real, imag} */,
  {32'hc506e8c1, 32'h00000000} /* (27, 24, 18) {real, imag} */,
  {32'hc4a4e3d8, 32'h00000000} /* (27, 24, 17) {real, imag} */,
  {32'hc507c51e, 32'h00000000} /* (27, 24, 16) {real, imag} */,
  {32'hc54f650c, 32'h00000000} /* (27, 24, 15) {real, imag} */,
  {32'hc534737e, 32'h00000000} /* (27, 24, 14) {real, imag} */,
  {32'hc4962590, 32'h00000000} /* (27, 24, 13) {real, imag} */,
  {32'hc50665ab, 32'h00000000} /* (27, 24, 12) {real, imag} */,
  {32'hc4f61e5c, 32'h00000000} /* (27, 24, 11) {real, imag} */,
  {32'h43134d88, 32'h00000000} /* (27, 24, 10) {real, imag} */,
  {32'h4505a136, 32'h00000000} /* (27, 24, 9) {real, imag} */,
  {32'h455d43bb, 32'h00000000} /* (27, 24, 8) {real, imag} */,
  {32'h44edd7a6, 32'h00000000} /* (27, 24, 7) {real, imag} */,
  {32'h45063d7d, 32'h00000000} /* (27, 24, 6) {real, imag} */,
  {32'h43ff9126, 32'h00000000} /* (27, 24, 5) {real, imag} */,
  {32'h43989bd6, 32'h00000000} /* (27, 24, 4) {real, imag} */,
  {32'h431ba10c, 32'h00000000} /* (27, 24, 3) {real, imag} */,
  {32'hc387dc68, 32'h00000000} /* (27, 24, 2) {real, imag} */,
  {32'h43447800, 32'h00000000} /* (27, 24, 1) {real, imag} */,
  {32'hc403909e, 32'h00000000} /* (27, 24, 0) {real, imag} */,
  {32'hc3c64a80, 32'h00000000} /* (27, 23, 31) {real, imag} */,
  {32'h441a7194, 32'h00000000} /* (27, 23, 30) {real, imag} */,
  {32'h44372461, 32'h00000000} /* (27, 23, 29) {real, imag} */,
  {32'h44505a22, 32'h00000000} /* (27, 23, 28) {real, imag} */,
  {32'h450da005, 32'h00000000} /* (27, 23, 27) {real, imag} */,
  {32'h4479ebf1, 32'h00000000} /* (27, 23, 26) {real, imag} */,
  {32'h4419c180, 32'h00000000} /* (27, 23, 25) {real, imag} */,
  {32'h449ad690, 32'h00000000} /* (27, 23, 24) {real, imag} */,
  {32'h450d1699, 32'h00000000} /* (27, 23, 23) {real, imag} */,
  {32'h44f3ff48, 32'h00000000} /* (27, 23, 22) {real, imag} */,
  {32'h440e70ff, 32'h00000000} /* (27, 23, 21) {real, imag} */,
  {32'hc43fc878, 32'h00000000} /* (27, 23, 20) {real, imag} */,
  {32'hc4d507f6, 32'h00000000} /* (27, 23, 19) {real, imag} */,
  {32'hc4e97540, 32'h00000000} /* (27, 23, 18) {real, imag} */,
  {32'hc4db5a8c, 32'h00000000} /* (27, 23, 17) {real, imag} */,
  {32'hc4bc21d1, 32'h00000000} /* (27, 23, 16) {real, imag} */,
  {32'hc4ff93e0, 32'h00000000} /* (27, 23, 15) {real, imag} */,
  {32'hc52669a4, 32'h00000000} /* (27, 23, 14) {real, imag} */,
  {32'hc49a7cc2, 32'h00000000} /* (27, 23, 13) {real, imag} */,
  {32'hc4ac26af, 32'h00000000} /* (27, 23, 12) {real, imag} */,
  {32'hc49334b4, 32'h00000000} /* (27, 23, 11) {real, imag} */,
  {32'h44bcbc74, 32'h00000000} /* (27, 23, 10) {real, imag} */,
  {32'h44fec88e, 32'h00000000} /* (27, 23, 9) {real, imag} */,
  {32'h4535835e, 32'h00000000} /* (27, 23, 8) {real, imag} */,
  {32'h450bcf71, 32'h00000000} /* (27, 23, 7) {real, imag} */,
  {32'h44c5c186, 32'h00000000} /* (27, 23, 6) {real, imag} */,
  {32'h4404ffa9, 32'h00000000} /* (27, 23, 5) {real, imag} */,
  {32'h440e7968, 32'h00000000} /* (27, 23, 4) {real, imag} */,
  {32'h4333b93c, 32'h00000000} /* (27, 23, 3) {real, imag} */,
  {32'h4401d9ef, 32'h00000000} /* (27, 23, 2) {real, imag} */,
  {32'hc358a8e8, 32'h00000000} /* (27, 23, 1) {real, imag} */,
  {32'hc24eabc0, 32'h00000000} /* (27, 23, 0) {real, imag} */,
  {32'hc36ad87c, 32'h00000000} /* (27, 22, 31) {real, imag} */,
  {32'h4410cc74, 32'h00000000} /* (27, 22, 30) {real, imag} */,
  {32'h4425d43a, 32'h00000000} /* (27, 22, 29) {real, imag} */,
  {32'h443eca86, 32'h00000000} /* (27, 22, 28) {real, imag} */,
  {32'h43fb3c8d, 32'h00000000} /* (27, 22, 27) {real, imag} */,
  {32'h4452ffe2, 32'h00000000} /* (27, 22, 26) {real, imag} */,
  {32'h431f1358, 32'h00000000} /* (27, 22, 25) {real, imag} */,
  {32'h438245ee, 32'h00000000} /* (27, 22, 24) {real, imag} */,
  {32'h43cfe118, 32'h00000000} /* (27, 22, 23) {real, imag} */,
  {32'h444bda7d, 32'h00000000} /* (27, 22, 22) {real, imag} */,
  {32'h41b09e20, 32'h00000000} /* (27, 22, 21) {real, imag} */,
  {32'hc49e3895, 32'h00000000} /* (27, 22, 20) {real, imag} */,
  {32'hc4688020, 32'h00000000} /* (27, 22, 19) {real, imag} */,
  {32'hc4a4f634, 32'h00000000} /* (27, 22, 18) {real, imag} */,
  {32'hc4a875dc, 32'h00000000} /* (27, 22, 17) {real, imag} */,
  {32'hc46a7442, 32'h00000000} /* (27, 22, 16) {real, imag} */,
  {32'hc432d383, 32'h00000000} /* (27, 22, 15) {real, imag} */,
  {32'hc420930a, 32'h00000000} /* (27, 22, 14) {real, imag} */,
  {32'hc4bb6aaf, 32'h00000000} /* (27, 22, 13) {real, imag} */,
  {32'hc401aaa6, 32'h00000000} /* (27, 22, 12) {real, imag} */,
  {32'h427243f8, 32'h00000000} /* (27, 22, 11) {real, imag} */,
  {32'h44855c74, 32'h00000000} /* (27, 22, 10) {real, imag} */,
  {32'h4478f646, 32'h00000000} /* (27, 22, 9) {real, imag} */,
  {32'h4491b42a, 32'h00000000} /* (27, 22, 8) {real, imag} */,
  {32'h44f04e12, 32'h00000000} /* (27, 22, 7) {real, imag} */,
  {32'h4481fdaa, 32'h00000000} /* (27, 22, 6) {real, imag} */,
  {32'h444eb93b, 32'h00000000} /* (27, 22, 5) {real, imag} */,
  {32'h43d49764, 32'h00000000} /* (27, 22, 4) {real, imag} */,
  {32'h448495a7, 32'h00000000} /* (27, 22, 3) {real, imag} */,
  {32'h43f21f16, 32'h00000000} /* (27, 22, 2) {real, imag} */,
  {32'h43bf7027, 32'h00000000} /* (27, 22, 1) {real, imag} */,
  {32'h441919e2, 32'h00000000} /* (27, 22, 0) {real, imag} */,
  {32'hc3b1977f, 32'h00000000} /* (27, 21, 31) {real, imag} */,
  {32'hc3f83491, 32'h00000000} /* (27, 21, 30) {real, imag} */,
  {32'hc419f432, 32'h00000000} /* (27, 21, 29) {real, imag} */,
  {32'hc402728a, 32'h00000000} /* (27, 21, 28) {real, imag} */,
  {32'h4269d038, 32'h00000000} /* (27, 21, 27) {real, imag} */,
  {32'hc2c56fa4, 32'h00000000} /* (27, 21, 26) {real, imag} */,
  {32'hc48a6e1e, 32'h00000000} /* (27, 21, 25) {real, imag} */,
  {32'hc47f43bf, 32'h00000000} /* (27, 21, 24) {real, imag} */,
  {32'hc43589b3, 32'h00000000} /* (27, 21, 23) {real, imag} */,
  {32'hc3a991d8, 32'h00000000} /* (27, 21, 22) {real, imag} */,
  {32'h41d95140, 32'h00000000} /* (27, 21, 21) {real, imag} */,
  {32'hc275ed18, 32'h00000000} /* (27, 21, 20) {real, imag} */,
  {32'h43f67630, 32'h00000000} /* (27, 21, 19) {real, imag} */,
  {32'h44164d27, 32'h00000000} /* (27, 21, 18) {real, imag} */,
  {32'h44603bce, 32'h00000000} /* (27, 21, 17) {real, imag} */,
  {32'hc409707d, 32'h00000000} /* (27, 21, 16) {real, imag} */,
  {32'hc21a1118, 32'h00000000} /* (27, 21, 15) {real, imag} */,
  {32'h442719f7, 32'h00000000} /* (27, 21, 14) {real, imag} */,
  {32'h4408e4ce, 32'h00000000} /* (27, 21, 13) {real, imag} */,
  {32'hc3790c73, 32'h00000000} /* (27, 21, 12) {real, imag} */,
  {32'h43a17d20, 32'h00000000} /* (27, 21, 11) {real, imag} */,
  {32'h446251e4, 32'h00000000} /* (27, 21, 10) {real, imag} */,
  {32'h44eb682e, 32'h00000000} /* (27, 21, 9) {real, imag} */,
  {32'h438245aa, 32'h00000000} /* (27, 21, 8) {real, imag} */,
  {32'hc24822a0, 32'h00000000} /* (27, 21, 7) {real, imag} */,
  {32'h441a3006, 32'h00000000} /* (27, 21, 6) {real, imag} */,
  {32'hc363443e, 32'h00000000} /* (27, 21, 5) {real, imag} */,
  {32'hc4424626, 32'h00000000} /* (27, 21, 4) {real, imag} */,
  {32'h44338a36, 32'h00000000} /* (27, 21, 3) {real, imag} */,
  {32'hc31e2cfb, 32'h00000000} /* (27, 21, 2) {real, imag} */,
  {32'hc3d9380c, 32'h00000000} /* (27, 21, 1) {real, imag} */,
  {32'hc3c3eb16, 32'h00000000} /* (27, 21, 0) {real, imag} */,
  {32'hc48c93d3, 32'h00000000} /* (27, 20, 31) {real, imag} */,
  {32'hc4983196, 32'h00000000} /* (27, 20, 30) {real, imag} */,
  {32'hc4d8613c, 32'h00000000} /* (27, 20, 29) {real, imag} */,
  {32'hc5383c70, 32'h00000000} /* (27, 20, 28) {real, imag} */,
  {32'hc4b585f0, 32'h00000000} /* (27, 20, 27) {real, imag} */,
  {32'hc4b15e22, 32'h00000000} /* (27, 20, 26) {real, imag} */,
  {32'hc538dd94, 32'h00000000} /* (27, 20, 25) {real, imag} */,
  {32'hc5085050, 32'h00000000} /* (27, 20, 24) {real, imag} */,
  {32'hc494e1fc, 32'h00000000} /* (27, 20, 23) {real, imag} */,
  {32'hc4bf0db8, 32'h00000000} /* (27, 20, 22) {real, imag} */,
  {32'hc3e8f368, 32'h00000000} /* (27, 20, 21) {real, imag} */,
  {32'h43c73028, 32'h00000000} /* (27, 20, 20) {real, imag} */,
  {32'h44768b69, 32'h00000000} /* (27, 20, 19) {real, imag} */,
  {32'h45314e62, 32'h00000000} /* (27, 20, 18) {real, imag} */,
  {32'h450bc0ae, 32'h00000000} /* (27, 20, 17) {real, imag} */,
  {32'h4519ee0b, 32'h00000000} /* (27, 20, 16) {real, imag} */,
  {32'h44d58bcf, 32'h00000000} /* (27, 20, 15) {real, imag} */,
  {32'h44f14620, 32'h00000000} /* (27, 20, 14) {real, imag} */,
  {32'h44d2fe6e, 32'h00000000} /* (27, 20, 13) {real, imag} */,
  {32'h449a4538, 32'h00000000} /* (27, 20, 12) {real, imag} */,
  {32'h4400901f, 32'h00000000} /* (27, 20, 11) {real, imag} */,
  {32'hc332f8d4, 32'h00000000} /* (27, 20, 10) {real, imag} */,
  {32'hc3bdd64c, 32'h00000000} /* (27, 20, 9) {real, imag} */,
  {32'hc4595209, 32'h00000000} /* (27, 20, 8) {real, imag} */,
  {32'hc4b9e398, 32'h00000000} /* (27, 20, 7) {real, imag} */,
  {32'hc4cdfce8, 32'h00000000} /* (27, 20, 6) {real, imag} */,
  {32'hc4dd5c52, 32'h00000000} /* (27, 20, 5) {real, imag} */,
  {32'hc4e3b034, 32'h00000000} /* (27, 20, 4) {real, imag} */,
  {32'hc50ee908, 32'h00000000} /* (27, 20, 3) {real, imag} */,
  {32'hc4f95c75, 32'h00000000} /* (27, 20, 2) {real, imag} */,
  {32'hc4e2ba42, 32'h00000000} /* (27, 20, 1) {real, imag} */,
  {32'hc4b00eb8, 32'h00000000} /* (27, 20, 0) {real, imag} */,
  {32'hc4f0530b, 32'h00000000} /* (27, 19, 31) {real, imag} */,
  {32'hc4cfe7dc, 32'h00000000} /* (27, 19, 30) {real, imag} */,
  {32'hc4e8b616, 32'h00000000} /* (27, 19, 29) {real, imag} */,
  {32'hc500448e, 32'h00000000} /* (27, 19, 28) {real, imag} */,
  {32'hc529f1c6, 32'h00000000} /* (27, 19, 27) {real, imag} */,
  {32'hc517610e, 32'h00000000} /* (27, 19, 26) {real, imag} */,
  {32'hc5036320, 32'h00000000} /* (27, 19, 25) {real, imag} */,
  {32'hc5373d94, 32'h00000000} /* (27, 19, 24) {real, imag} */,
  {32'hc527a327, 32'h00000000} /* (27, 19, 23) {real, imag} */,
  {32'hc4c75a84, 32'h00000000} /* (27, 19, 22) {real, imag} */,
  {32'hc4281342, 32'h00000000} /* (27, 19, 21) {real, imag} */,
  {32'h449a704e, 32'h00000000} /* (27, 19, 20) {real, imag} */,
  {32'h449aaa4b, 32'h00000000} /* (27, 19, 19) {real, imag} */,
  {32'h44ed24de, 32'h00000000} /* (27, 19, 18) {real, imag} */,
  {32'h451d27b9, 32'h00000000} /* (27, 19, 17) {real, imag} */,
  {32'h4515e452, 32'h00000000} /* (27, 19, 16) {real, imag} */,
  {32'h4559edbe, 32'h00000000} /* (27, 19, 15) {real, imag} */,
  {32'h452a430a, 32'h00000000} /* (27, 19, 14) {real, imag} */,
  {32'h4515d0cf, 32'h00000000} /* (27, 19, 13) {real, imag} */,
  {32'h44d50e5c, 32'h00000000} /* (27, 19, 12) {real, imag} */,
  {32'h44858ed4, 32'h00000000} /* (27, 19, 11) {real, imag} */,
  {32'h43669548, 32'h00000000} /* (27, 19, 10) {real, imag} */,
  {32'hc418989a, 32'h00000000} /* (27, 19, 9) {real, imag} */,
  {32'hc4c13ebf, 32'h00000000} /* (27, 19, 8) {real, imag} */,
  {32'hc4d33c69, 32'h00000000} /* (27, 19, 7) {real, imag} */,
  {32'hc4af5894, 32'h00000000} /* (27, 19, 6) {real, imag} */,
  {32'hc536a5c2, 32'h00000000} /* (27, 19, 5) {real, imag} */,
  {32'hc51e53a3, 32'h00000000} /* (27, 19, 4) {real, imag} */,
  {32'hc5208ef4, 32'h00000000} /* (27, 19, 3) {real, imag} */,
  {32'hc56606a5, 32'h00000000} /* (27, 19, 2) {real, imag} */,
  {32'hc4b53cd4, 32'h00000000} /* (27, 19, 1) {real, imag} */,
  {32'hc492ba3f, 32'h00000000} /* (27, 19, 0) {real, imag} */,
  {32'hc4f68367, 32'h00000000} /* (27, 18, 31) {real, imag} */,
  {32'hc512f073, 32'h00000000} /* (27, 18, 30) {real, imag} */,
  {32'hc5274ea1, 32'h00000000} /* (27, 18, 29) {real, imag} */,
  {32'hc5146f76, 32'h00000000} /* (27, 18, 28) {real, imag} */,
  {32'hc524ff94, 32'h00000000} /* (27, 18, 27) {real, imag} */,
  {32'hc53b03be, 32'h00000000} /* (27, 18, 26) {real, imag} */,
  {32'hc5348bdc, 32'h00000000} /* (27, 18, 25) {real, imag} */,
  {32'hc564134f, 32'h00000000} /* (27, 18, 24) {real, imag} */,
  {32'hc53392c7, 32'h00000000} /* (27, 18, 23) {real, imag} */,
  {32'hc51fe557, 32'h00000000} /* (27, 18, 22) {real, imag} */,
  {32'hc3f95170, 32'h00000000} /* (27, 18, 21) {real, imag} */,
  {32'hc1bd7300, 32'h00000000} /* (27, 18, 20) {real, imag} */,
  {32'h445d88bc, 32'h00000000} /* (27, 18, 19) {real, imag} */,
  {32'h45112766, 32'h00000000} /* (27, 18, 18) {real, imag} */,
  {32'h4513ed04, 32'h00000000} /* (27, 18, 17) {real, imag} */,
  {32'h4537e759, 32'h00000000} /* (27, 18, 16) {real, imag} */,
  {32'h4537680c, 32'h00000000} /* (27, 18, 15) {real, imag} */,
  {32'h451fa6a1, 32'h00000000} /* (27, 18, 14) {real, imag} */,
  {32'h455491a9, 32'h00000000} /* (27, 18, 13) {real, imag} */,
  {32'h45027fd6, 32'h00000000} /* (27, 18, 12) {real, imag} */,
  {32'h44c691bd, 32'h00000000} /* (27, 18, 11) {real, imag} */,
  {32'h424eece0, 32'h00000000} /* (27, 18, 10) {real, imag} */,
  {32'hc406d30e, 32'h00000000} /* (27, 18, 9) {real, imag} */,
  {32'hc4b5e87e, 32'h00000000} /* (27, 18, 8) {real, imag} */,
  {32'hc4f6ff0a, 32'h00000000} /* (27, 18, 7) {real, imag} */,
  {32'hc562a56b, 32'h00000000} /* (27, 18, 6) {real, imag} */,
  {32'hc56140f0, 32'h00000000} /* (27, 18, 5) {real, imag} */,
  {32'hc5240314, 32'h00000000} /* (27, 18, 4) {real, imag} */,
  {32'hc53c2332, 32'h00000000} /* (27, 18, 3) {real, imag} */,
  {32'hc4b8ad05, 32'h00000000} /* (27, 18, 2) {real, imag} */,
  {32'hc4e10343, 32'h00000000} /* (27, 18, 1) {real, imag} */,
  {32'hc4a313ca, 32'h00000000} /* (27, 18, 0) {real, imag} */,
  {32'hc4de2790, 32'h00000000} /* (27, 17, 31) {real, imag} */,
  {32'hc52ee9c1, 32'h00000000} /* (27, 17, 30) {real, imag} */,
  {32'hc5549000, 32'h00000000} /* (27, 17, 29) {real, imag} */,
  {32'hc53aa89f, 32'h00000000} /* (27, 17, 28) {real, imag} */,
  {32'hc53659a9, 32'h00000000} /* (27, 17, 27) {real, imag} */,
  {32'hc4fab4d0, 32'h00000000} /* (27, 17, 26) {real, imag} */,
  {32'hc5443297, 32'h00000000} /* (27, 17, 25) {real, imag} */,
  {32'hc569befc, 32'h00000000} /* (27, 17, 24) {real, imag} */,
  {32'hc552c16e, 32'h00000000} /* (27, 17, 23) {real, imag} */,
  {32'hc50700e6, 32'h00000000} /* (27, 17, 22) {real, imag} */,
  {32'hc4f16f03, 32'h00000000} /* (27, 17, 21) {real, imag} */,
  {32'h42d41720, 32'h00000000} /* (27, 17, 20) {real, imag} */,
  {32'h44c7739c, 32'h00000000} /* (27, 17, 19) {real, imag} */,
  {32'h451232b5, 32'h00000000} /* (27, 17, 18) {real, imag} */,
  {32'h457021e7, 32'h00000000} /* (27, 17, 17) {real, imag} */,
  {32'h452efd97, 32'h00000000} /* (27, 17, 16) {real, imag} */,
  {32'h4502c867, 32'h00000000} /* (27, 17, 15) {real, imag} */,
  {32'h45250291, 32'h00000000} /* (27, 17, 14) {real, imag} */,
  {32'h451373be, 32'h00000000} /* (27, 17, 13) {real, imag} */,
  {32'h44b8ade6, 32'h00000000} /* (27, 17, 12) {real, imag} */,
  {32'h44c6577e, 32'h00000000} /* (27, 17, 11) {real, imag} */,
  {32'hc0b15880, 32'h00000000} /* (27, 17, 10) {real, imag} */,
  {32'hc49a739e, 32'h00000000} /* (27, 17, 9) {real, imag} */,
  {32'hc4ca97b4, 32'h00000000} /* (27, 17, 8) {real, imag} */,
  {32'hc4fe095d, 32'h00000000} /* (27, 17, 7) {real, imag} */,
  {32'hc550370c, 32'h00000000} /* (27, 17, 6) {real, imag} */,
  {32'hc52974f8, 32'h00000000} /* (27, 17, 5) {real, imag} */,
  {32'hc5346591, 32'h00000000} /* (27, 17, 4) {real, imag} */,
  {32'hc52355e0, 32'h00000000} /* (27, 17, 3) {real, imag} */,
  {32'hc54e7cdb, 32'h00000000} /* (27, 17, 2) {real, imag} */,
  {32'hc4bd8d5e, 32'h00000000} /* (27, 17, 1) {real, imag} */,
  {32'hc471fba5, 32'h00000000} /* (27, 17, 0) {real, imag} */,
  {32'hc4be913b, 32'h00000000} /* (27, 16, 31) {real, imag} */,
  {32'hc534a272, 32'h00000000} /* (27, 16, 30) {real, imag} */,
  {32'hc5580512, 32'h00000000} /* (27, 16, 29) {real, imag} */,
  {32'hc52513f6, 32'h00000000} /* (27, 16, 28) {real, imag} */,
  {32'hc532abb1, 32'h00000000} /* (27, 16, 27) {real, imag} */,
  {32'hc52d997f, 32'h00000000} /* (27, 16, 26) {real, imag} */,
  {32'hc570c3cc, 32'h00000000} /* (27, 16, 25) {real, imag} */,
  {32'hc541b65c, 32'h00000000} /* (27, 16, 24) {real, imag} */,
  {32'hc5526651, 32'h00000000} /* (27, 16, 23) {real, imag} */,
  {32'hc503ee06, 32'h00000000} /* (27, 16, 22) {real, imag} */,
  {32'hc42500b4, 32'h00000000} /* (27, 16, 21) {real, imag} */,
  {32'h4461c132, 32'h00000000} /* (27, 16, 20) {real, imag} */,
  {32'h44e34473, 32'h00000000} /* (27, 16, 19) {real, imag} */,
  {32'h44fea8bc, 32'h00000000} /* (27, 16, 18) {real, imag} */,
  {32'h45195a29, 32'h00000000} /* (27, 16, 17) {real, imag} */,
  {32'h4501fcf6, 32'h00000000} /* (27, 16, 16) {real, imag} */,
  {32'h451ebeca, 32'h00000000} /* (27, 16, 15) {real, imag} */,
  {32'h44f7bd4f, 32'h00000000} /* (27, 16, 14) {real, imag} */,
  {32'h450a4cc2, 32'h00000000} /* (27, 16, 13) {real, imag} */,
  {32'h44f2975c, 32'h00000000} /* (27, 16, 12) {real, imag} */,
  {32'h44a08a36, 32'h00000000} /* (27, 16, 11) {real, imag} */,
  {32'hc4537b83, 32'h00000000} /* (27, 16, 10) {real, imag} */,
  {32'hc497c68d, 32'h00000000} /* (27, 16, 9) {real, imag} */,
  {32'hc4c99c85, 32'h00000000} /* (27, 16, 8) {real, imag} */,
  {32'hc5197edb, 32'h00000000} /* (27, 16, 7) {real, imag} */,
  {32'hc533e4ae, 32'h00000000} /* (27, 16, 6) {real, imag} */,
  {32'hc5168712, 32'h00000000} /* (27, 16, 5) {real, imag} */,
  {32'hc54305ca, 32'h00000000} /* (27, 16, 4) {real, imag} */,
  {32'hc5333a86, 32'h00000000} /* (27, 16, 3) {real, imag} */,
  {32'hc50cf176, 32'h00000000} /* (27, 16, 2) {real, imag} */,
  {32'hc5114a35, 32'h00000000} /* (27, 16, 1) {real, imag} */,
  {32'hc501dc0a, 32'h00000000} /* (27, 16, 0) {real, imag} */,
  {32'hc5116498, 32'h00000000} /* (27, 15, 31) {real, imag} */,
  {32'hc503925c, 32'h00000000} /* (27, 15, 30) {real, imag} */,
  {32'hc52bfff8, 32'h00000000} /* (27, 15, 29) {real, imag} */,
  {32'hc54c7dbc, 32'h00000000} /* (27, 15, 28) {real, imag} */,
  {32'hc530f754, 32'h00000000} /* (27, 15, 27) {real, imag} */,
  {32'hc56f87ec, 32'h00000000} /* (27, 15, 26) {real, imag} */,
  {32'hc55a8a1a, 32'h00000000} /* (27, 15, 25) {real, imag} */,
  {32'hc5463597, 32'h00000000} /* (27, 15, 24) {real, imag} */,
  {32'hc5135154, 32'h00000000} /* (27, 15, 23) {real, imag} */,
  {32'hc55cd22b, 32'h00000000} /* (27, 15, 22) {real, imag} */,
  {32'hc4c15922, 32'h00000000} /* (27, 15, 21) {real, imag} */,
  {32'h44404084, 32'h00000000} /* (27, 15, 20) {real, imag} */,
  {32'h44cdf26c, 32'h00000000} /* (27, 15, 19) {real, imag} */,
  {32'h44c8f170, 32'h00000000} /* (27, 15, 18) {real, imag} */,
  {32'h450365fc, 32'h00000000} /* (27, 15, 17) {real, imag} */,
  {32'h44f84247, 32'h00000000} /* (27, 15, 16) {real, imag} */,
  {32'h451080e4, 32'h00000000} /* (27, 15, 15) {real, imag} */,
  {32'h44cc2950, 32'h00000000} /* (27, 15, 14) {real, imag} */,
  {32'h44d5a19f, 32'h00000000} /* (27, 15, 13) {real, imag} */,
  {32'h443eacc0, 32'h00000000} /* (27, 15, 12) {real, imag} */,
  {32'h44c565e7, 32'h00000000} /* (27, 15, 11) {real, imag} */,
  {32'hc4511d9a, 32'h00000000} /* (27, 15, 10) {real, imag} */,
  {32'hc4fab535, 32'h00000000} /* (27, 15, 9) {real, imag} */,
  {32'hc500270d, 32'h00000000} /* (27, 15, 8) {real, imag} */,
  {32'hc51d528c, 32'h00000000} /* (27, 15, 7) {real, imag} */,
  {32'hc531b639, 32'h00000000} /* (27, 15, 6) {real, imag} */,
  {32'hc537a82b, 32'h00000000} /* (27, 15, 5) {real, imag} */,
  {32'hc5132a45, 32'h00000000} /* (27, 15, 4) {real, imag} */,
  {32'hc5137b56, 32'h00000000} /* (27, 15, 3) {real, imag} */,
  {32'hc4eda9a4, 32'h00000000} /* (27, 15, 2) {real, imag} */,
  {32'hc514035c, 32'h00000000} /* (27, 15, 1) {real, imag} */,
  {32'hc4dbf059, 32'h00000000} /* (27, 15, 0) {real, imag} */,
  {32'hc5016f1b, 32'h00000000} /* (27, 14, 31) {real, imag} */,
  {32'hc54f9d06, 32'h00000000} /* (27, 14, 30) {real, imag} */,
  {32'hc5140201, 32'h00000000} /* (27, 14, 29) {real, imag} */,
  {32'hc5485e8e, 32'h00000000} /* (27, 14, 28) {real, imag} */,
  {32'hc546e3c8, 32'h00000000} /* (27, 14, 27) {real, imag} */,
  {32'hc52f2d1f, 32'h00000000} /* (27, 14, 26) {real, imag} */,
  {32'hc54c8cea, 32'h00000000} /* (27, 14, 25) {real, imag} */,
  {32'hc5498fb2, 32'h00000000} /* (27, 14, 24) {real, imag} */,
  {32'hc546d1c8, 32'h00000000} /* (27, 14, 23) {real, imag} */,
  {32'hc53c4938, 32'h00000000} /* (27, 14, 22) {real, imag} */,
  {32'hc462f03c, 32'h00000000} /* (27, 14, 21) {real, imag} */,
  {32'h43b6cce6, 32'h00000000} /* (27, 14, 20) {real, imag} */,
  {32'h449f9313, 32'h00000000} /* (27, 14, 19) {real, imag} */,
  {32'h450cb815, 32'h00000000} /* (27, 14, 18) {real, imag} */,
  {32'h44b9684d, 32'h00000000} /* (27, 14, 17) {real, imag} */,
  {32'h44e11471, 32'h00000000} /* (27, 14, 16) {real, imag} */,
  {32'h45076e71, 32'h00000000} /* (27, 14, 15) {real, imag} */,
  {32'h44cd96d9, 32'h00000000} /* (27, 14, 14) {real, imag} */,
  {32'h44b48798, 32'h00000000} /* (27, 14, 13) {real, imag} */,
  {32'h44e5812c, 32'h00000000} /* (27, 14, 12) {real, imag} */,
  {32'h44735972, 32'h00000000} /* (27, 14, 11) {real, imag} */,
  {32'hc4371a5c, 32'h00000000} /* (27, 14, 10) {real, imag} */,
  {32'hc4f8dee5, 32'h00000000} /* (27, 14, 9) {real, imag} */,
  {32'hc515098a, 32'h00000000} /* (27, 14, 8) {real, imag} */,
  {32'hc53975fe, 32'h00000000} /* (27, 14, 7) {real, imag} */,
  {32'hc4de03f8, 32'h00000000} /* (27, 14, 6) {real, imag} */,
  {32'hc4dce20e, 32'h00000000} /* (27, 14, 5) {real, imag} */,
  {32'hc509aee4, 32'h00000000} /* (27, 14, 4) {real, imag} */,
  {32'hc4f3e6fd, 32'h00000000} /* (27, 14, 3) {real, imag} */,
  {32'hc501cd23, 32'h00000000} /* (27, 14, 2) {real, imag} */,
  {32'hc51e50ce, 32'h00000000} /* (27, 14, 1) {real, imag} */,
  {32'hc47c2cb6, 32'h00000000} /* (27, 14, 0) {real, imag} */,
  {32'hc509ee4f, 32'h00000000} /* (27, 13, 31) {real, imag} */,
  {32'hc531a8d0, 32'h00000000} /* (27, 13, 30) {real, imag} */,
  {32'hc5281215, 32'h00000000} /* (27, 13, 29) {real, imag} */,
  {32'hc5131085, 32'h00000000} /* (27, 13, 28) {real, imag} */,
  {32'hc520caca, 32'h00000000} /* (27, 13, 27) {real, imag} */,
  {32'hc4f57492, 32'h00000000} /* (27, 13, 26) {real, imag} */,
  {32'hc529af1e, 32'h00000000} /* (27, 13, 25) {real, imag} */,
  {32'hc52b22e8, 32'h00000000} /* (27, 13, 24) {real, imag} */,
  {32'hc524f782, 32'h00000000} /* (27, 13, 23) {real, imag} */,
  {32'hc4b941d8, 32'h00000000} /* (27, 13, 22) {real, imag} */,
  {32'hc4b8aaf4, 32'h00000000} /* (27, 13, 21) {real, imag} */,
  {32'hc30c31ac, 32'h00000000} /* (27, 13, 20) {real, imag} */,
  {32'h44323146, 32'h00000000} /* (27, 13, 19) {real, imag} */,
  {32'h44d4a97d, 32'h00000000} /* (27, 13, 18) {real, imag} */,
  {32'h44f9cbaf, 32'h00000000} /* (27, 13, 17) {real, imag} */,
  {32'h44ede642, 32'h00000000} /* (27, 13, 16) {real, imag} */,
  {32'h448c3c82, 32'h00000000} /* (27, 13, 15) {real, imag} */,
  {32'h44b55085, 32'h00000000} /* (27, 13, 14) {real, imag} */,
  {32'h44a75d5c, 32'h00000000} /* (27, 13, 13) {real, imag} */,
  {32'h44ad175a, 32'h00000000} /* (27, 13, 12) {real, imag} */,
  {32'h447faef4, 32'h00000000} /* (27, 13, 11) {real, imag} */,
  {32'hc457550c, 32'h00000000} /* (27, 13, 10) {real, imag} */,
  {32'hc50c1c5a, 32'h00000000} /* (27, 13, 9) {real, imag} */,
  {32'hc4ee0c20, 32'h00000000} /* (27, 13, 8) {real, imag} */,
  {32'hc545d208, 32'h00000000} /* (27, 13, 7) {real, imag} */,
  {32'hc4eb231a, 32'h00000000} /* (27, 13, 6) {real, imag} */,
  {32'hc491bd78, 32'h00000000} /* (27, 13, 5) {real, imag} */,
  {32'hc4dc670e, 32'h00000000} /* (27, 13, 4) {real, imag} */,
  {32'hc51fd4d0, 32'h00000000} /* (27, 13, 3) {real, imag} */,
  {32'hc503f0d4, 32'h00000000} /* (27, 13, 2) {real, imag} */,
  {32'hc4cc401f, 32'h00000000} /* (27, 13, 1) {real, imag} */,
  {32'hc4b0124c, 32'h00000000} /* (27, 13, 0) {real, imag} */,
  {32'hc4e6e43a, 32'h00000000} /* (27, 12, 31) {real, imag} */,
  {32'hc5039921, 32'h00000000} /* (27, 12, 30) {real, imag} */,
  {32'hc4d6c78c, 32'h00000000} /* (27, 12, 29) {real, imag} */,
  {32'hc51dae6f, 32'h00000000} /* (27, 12, 28) {real, imag} */,
  {32'hc5106786, 32'h00000000} /* (27, 12, 27) {real, imag} */,
  {32'hc5150c5c, 32'h00000000} /* (27, 12, 26) {real, imag} */,
  {32'hc5350734, 32'h00000000} /* (27, 12, 25) {real, imag} */,
  {32'hc4e4f0fe, 32'h00000000} /* (27, 12, 24) {real, imag} */,
  {32'hc4c4732d, 32'h00000000} /* (27, 12, 23) {real, imag} */,
  {32'hc51926ee, 32'h00000000} /* (27, 12, 22) {real, imag} */,
  {32'hc3d76346, 32'h00000000} /* (27, 12, 21) {real, imag} */,
  {32'hc3bdf9d1, 32'h00000000} /* (27, 12, 20) {real, imag} */,
  {32'h4387d3b0, 32'h00000000} /* (27, 12, 19) {real, imag} */,
  {32'h44a3621a, 32'h00000000} /* (27, 12, 18) {real, imag} */,
  {32'h44ededd8, 32'h00000000} /* (27, 12, 17) {real, imag} */,
  {32'h44882174, 32'h00000000} /* (27, 12, 16) {real, imag} */,
  {32'h44417093, 32'h00000000} /* (27, 12, 15) {real, imag} */,
  {32'h44bae588, 32'h00000000} /* (27, 12, 14) {real, imag} */,
  {32'h44aec51a, 32'h00000000} /* (27, 12, 13) {real, imag} */,
  {32'h41925780, 32'h00000000} /* (27, 12, 12) {real, imag} */,
  {32'h4471ae08, 32'h00000000} /* (27, 12, 11) {real, imag} */,
  {32'hc3eac318, 32'h00000000} /* (27, 12, 10) {real, imag} */,
  {32'hc4c43bfc, 32'h00000000} /* (27, 12, 9) {real, imag} */,
  {32'hc4566334, 32'h00000000} /* (27, 12, 8) {real, imag} */,
  {32'hc4c7c61f, 32'h00000000} /* (27, 12, 7) {real, imag} */,
  {32'hc50a8866, 32'h00000000} /* (27, 12, 6) {real, imag} */,
  {32'hc4c46f9a, 32'h00000000} /* (27, 12, 5) {real, imag} */,
  {32'hc4a5600b, 32'h00000000} /* (27, 12, 4) {real, imag} */,
  {32'hc4d195a8, 32'h00000000} /* (27, 12, 3) {real, imag} */,
  {32'hc4fd1a70, 32'h00000000} /* (27, 12, 2) {real, imag} */,
  {32'hc4be4b96, 32'h00000000} /* (27, 12, 1) {real, imag} */,
  {32'hc4b1d2b8, 32'h00000000} /* (27, 12, 0) {real, imag} */,
  {32'hc44d2972, 32'h00000000} /* (27, 11, 31) {real, imag} */,
  {32'hc452f533, 32'h00000000} /* (27, 11, 30) {real, imag} */,
  {32'hc4a5277e, 32'h00000000} /* (27, 11, 29) {real, imag} */,
  {32'hc50d7954, 32'h00000000} /* (27, 11, 28) {real, imag} */,
  {32'hc4b8800e, 32'h00000000} /* (27, 11, 27) {real, imag} */,
  {32'hc4d62132, 32'h00000000} /* (27, 11, 26) {real, imag} */,
  {32'hc510b070, 32'h00000000} /* (27, 11, 25) {real, imag} */,
  {32'hc4a5c518, 32'h00000000} /* (27, 11, 24) {real, imag} */,
  {32'hc41c76a2, 32'h00000000} /* (27, 11, 23) {real, imag} */,
  {32'hc4bd21d2, 32'h00000000} /* (27, 11, 22) {real, imag} */,
  {32'hc233e470, 32'h00000000} /* (27, 11, 21) {real, imag} */,
  {32'h44002f2c, 32'h00000000} /* (27, 11, 20) {real, imag} */,
  {32'hc3c27d58, 32'h00000000} /* (27, 11, 19) {real, imag} */,
  {32'h447a1501, 32'h00000000} /* (27, 11, 18) {real, imag} */,
  {32'h44dfe2fb, 32'h00000000} /* (27, 11, 17) {real, imag} */,
  {32'h42fd0014, 32'h00000000} /* (27, 11, 16) {real, imag} */,
  {32'h44526bb6, 32'h00000000} /* (27, 11, 15) {real, imag} */,
  {32'h44c4f484, 32'h00000000} /* (27, 11, 14) {real, imag} */,
  {32'h4450f4bc, 32'h00000000} /* (27, 11, 13) {real, imag} */,
  {32'h43825904, 32'h00000000} /* (27, 11, 12) {real, imag} */,
  {32'hc2216120, 32'h00000000} /* (27, 11, 11) {real, imag} */,
  {32'hc439c444, 32'h00000000} /* (27, 11, 10) {real, imag} */,
  {32'hc46b008a, 32'h00000000} /* (27, 11, 9) {real, imag} */,
  {32'hc48014f2, 32'h00000000} /* (27, 11, 8) {real, imag} */,
  {32'hc40044da, 32'h00000000} /* (27, 11, 7) {real, imag} */,
  {32'hc47caadc, 32'h00000000} /* (27, 11, 6) {real, imag} */,
  {32'hc3b0f71c, 32'h00000000} /* (27, 11, 5) {real, imag} */,
  {32'hc42d4286, 32'h00000000} /* (27, 11, 4) {real, imag} */,
  {32'hc4b5b397, 32'h00000000} /* (27, 11, 3) {real, imag} */,
  {32'hc4a5ffca, 32'h00000000} /* (27, 11, 2) {real, imag} */,
  {32'hc4bc5b6d, 32'h00000000} /* (27, 11, 1) {real, imag} */,
  {32'hc43fad2a, 32'h00000000} /* (27, 11, 0) {real, imag} */,
  {32'h4340d7d9, 32'h00000000} /* (27, 10, 31) {real, imag} */,
  {32'h42f8dc46, 32'h00000000} /* (27, 10, 30) {real, imag} */,
  {32'hc397d0e1, 32'h00000000} /* (27, 10, 29) {real, imag} */,
  {32'hc3b4b3dd, 32'h00000000} /* (27, 10, 28) {real, imag} */,
  {32'hc3d8a852, 32'h00000000} /* (27, 10, 27) {real, imag} */,
  {32'h426c6f08, 32'h00000000} /* (27, 10, 26) {real, imag} */,
  {32'hc393728a, 32'h00000000} /* (27, 10, 25) {real, imag} */,
  {32'hc1d70340, 32'h00000000} /* (27, 10, 24) {real, imag} */,
  {32'h440d83b3, 32'h00000000} /* (27, 10, 23) {real, imag} */,
  {32'h448bb860, 32'h00000000} /* (27, 10, 22) {real, imag} */,
  {32'h4323da24, 32'h00000000} /* (27, 10, 21) {real, imag} */,
  {32'hc45a4a5e, 32'h00000000} /* (27, 10, 20) {real, imag} */,
  {32'hc4daf7d9, 32'h00000000} /* (27, 10, 19) {real, imag} */,
  {32'hc492bf27, 32'h00000000} /* (27, 10, 18) {real, imag} */,
  {32'hc48e7da8, 32'h00000000} /* (27, 10, 17) {real, imag} */,
  {32'hc48cc1eb, 32'h00000000} /* (27, 10, 16) {real, imag} */,
  {32'hc3269cc1, 32'h00000000} /* (27, 10, 15) {real, imag} */,
  {32'hc2d1db96, 32'h00000000} /* (27, 10, 14) {real, imag} */,
  {32'hc4040264, 32'h00000000} /* (27, 10, 13) {real, imag} */,
  {32'hc4636536, 32'h00000000} /* (27, 10, 12) {real, imag} */,
  {32'hc5016216, 32'h00000000} /* (27, 10, 11) {real, imag} */,
  {32'hc3c5eccb, 32'h00000000} /* (27, 10, 10) {real, imag} */,
  {32'h43c37348, 32'h00000000} /* (27, 10, 9) {real, imag} */,
  {32'h449b6821, 32'h00000000} /* (27, 10, 8) {real, imag} */,
  {32'h44f70eb6, 32'h00000000} /* (27, 10, 7) {real, imag} */,
  {32'h44fc8248, 32'h00000000} /* (27, 10, 6) {real, imag} */,
  {32'h444d3d13, 32'h00000000} /* (27, 10, 5) {real, imag} */,
  {32'h446fadd0, 32'h00000000} /* (27, 10, 4) {real, imag} */,
  {32'hc33b4a38, 32'h00000000} /* (27, 10, 3) {real, imag} */,
  {32'hc3900d65, 32'h00000000} /* (27, 10, 2) {real, imag} */,
  {32'h43d671be, 32'h00000000} /* (27, 10, 1) {real, imag} */,
  {32'h43085e7a, 32'h00000000} /* (27, 10, 0) {real, imag} */,
  {32'h445c9962, 32'h00000000} /* (27, 9, 31) {real, imag} */,
  {32'h4468ad35, 32'h00000000} /* (27, 9, 30) {real, imag} */,
  {32'h4433443e, 32'h00000000} /* (27, 9, 29) {real, imag} */,
  {32'h4450640b, 32'h00000000} /* (27, 9, 28) {real, imag} */,
  {32'h420b98c8, 32'h00000000} /* (27, 9, 27) {real, imag} */,
  {32'h429baa40, 32'h00000000} /* (27, 9, 26) {real, imag} */,
  {32'h44166d6f, 32'h00000000} /* (27, 9, 25) {real, imag} */,
  {32'h4440dc5e, 32'h00000000} /* (27, 9, 24) {real, imag} */,
  {32'h449604aa, 32'h00000000} /* (27, 9, 23) {real, imag} */,
  {32'h44976f87, 32'h00000000} /* (27, 9, 22) {real, imag} */,
  {32'h4425d4f2, 32'h00000000} /* (27, 9, 21) {real, imag} */,
  {32'hc4b3db1d, 32'h00000000} /* (27, 9, 20) {real, imag} */,
  {32'hc5340c24, 32'h00000000} /* (27, 9, 19) {real, imag} */,
  {32'hc4f03719, 32'h00000000} /* (27, 9, 18) {real, imag} */,
  {32'hc51183bb, 32'h00000000} /* (27, 9, 17) {real, imag} */,
  {32'hc5083c66, 32'h00000000} /* (27, 9, 16) {real, imag} */,
  {32'hc507731c, 32'h00000000} /* (27, 9, 15) {real, imag} */,
  {32'hc4d24d66, 32'h00000000} /* (27, 9, 14) {real, imag} */,
  {32'hc5196c96, 32'h00000000} /* (27, 9, 13) {real, imag} */,
  {32'hc4c531d4, 32'h00000000} /* (27, 9, 12) {real, imag} */,
  {32'hc445278a, 32'h00000000} /* (27, 9, 11) {real, imag} */,
  {32'h4412d18c, 32'h00000000} /* (27, 9, 10) {real, imag} */,
  {32'h44e9f168, 32'h00000000} /* (27, 9, 9) {real, imag} */,
  {32'h44e363bd, 32'h00000000} /* (27, 9, 8) {real, imag} */,
  {32'h44bd8c12, 32'h00000000} /* (27, 9, 7) {real, imag} */,
  {32'h44ce08d1, 32'h00000000} /* (27, 9, 6) {real, imag} */,
  {32'h44afba23, 32'h00000000} /* (27, 9, 5) {real, imag} */,
  {32'h446ef7f3, 32'h00000000} /* (27, 9, 4) {real, imag} */,
  {32'h4473fb2a, 32'h00000000} /* (27, 9, 3) {real, imag} */,
  {32'h440926f6, 32'h00000000} /* (27, 9, 2) {real, imag} */,
  {32'h448a860e, 32'h00000000} /* (27, 9, 1) {real, imag} */,
  {32'h44523a85, 32'h00000000} /* (27, 9, 0) {real, imag} */,
  {32'h438d7480, 32'h00000000} /* (27, 8, 31) {real, imag} */,
  {32'h4399b47c, 32'h00000000} /* (27, 8, 30) {real, imag} */,
  {32'h44d6cce5, 32'h00000000} /* (27, 8, 29) {real, imag} */,
  {32'h43037108, 32'h00000000} /* (27, 8, 28) {real, imag} */,
  {32'h43e118cc, 32'h00000000} /* (27, 8, 27) {real, imag} */,
  {32'h443235c2, 32'h00000000} /* (27, 8, 26) {real, imag} */,
  {32'h44629614, 32'h00000000} /* (27, 8, 25) {real, imag} */,
  {32'h4471d393, 32'h00000000} /* (27, 8, 24) {real, imag} */,
  {32'h43bc3db8, 32'h00000000} /* (27, 8, 23) {real, imag} */,
  {32'h4525dce8, 32'h00000000} /* (27, 8, 22) {real, imag} */,
  {32'h43a567d4, 32'h00000000} /* (27, 8, 21) {real, imag} */,
  {32'hc495385a, 32'h00000000} /* (27, 8, 20) {real, imag} */,
  {32'hc50967f5, 32'h00000000} /* (27, 8, 19) {real, imag} */,
  {32'hc547dfb1, 32'h00000000} /* (27, 8, 18) {real, imag} */,
  {32'hc50d6cb5, 32'h00000000} /* (27, 8, 17) {real, imag} */,
  {32'hc548f628, 32'h00000000} /* (27, 8, 16) {real, imag} */,
  {32'hc55a1828, 32'h00000000} /* (27, 8, 15) {real, imag} */,
  {32'hc51111f2, 32'h00000000} /* (27, 8, 14) {real, imag} */,
  {32'hc50f1bd6, 32'h00000000} /* (27, 8, 13) {real, imag} */,
  {32'hc505e6a4, 32'h00000000} /* (27, 8, 12) {real, imag} */,
  {32'hc50dc72a, 32'h00000000} /* (27, 8, 11) {real, imag} */,
  {32'hc3141052, 32'h00000000} /* (27, 8, 10) {real, imag} */,
  {32'h44bfe45e, 32'h00000000} /* (27, 8, 9) {real, imag} */,
  {32'h44d2e89e, 32'h00000000} /* (27, 8, 8) {real, imag} */,
  {32'h44e9b252, 32'h00000000} /* (27, 8, 7) {real, imag} */,
  {32'h450e7108, 32'h00000000} /* (27, 8, 6) {real, imag} */,
  {32'h44d3d4b5, 32'h00000000} /* (27, 8, 5) {real, imag} */,
  {32'h44c1c7b4, 32'h00000000} /* (27, 8, 4) {real, imag} */,
  {32'h44cea428, 32'h00000000} /* (27, 8, 3) {real, imag} */,
  {32'h4414163c, 32'h00000000} /* (27, 8, 2) {real, imag} */,
  {32'h442084bb, 32'h00000000} /* (27, 8, 1) {real, imag} */,
  {32'h443d2260, 32'h00000000} /* (27, 8, 0) {real, imag} */,
  {32'h4363edb0, 32'h00000000} /* (27, 7, 31) {real, imag} */,
  {32'h431056e8, 32'h00000000} /* (27, 7, 30) {real, imag} */,
  {32'hc398acf0, 32'h00000000} /* (27, 7, 29) {real, imag} */,
  {32'h43c04900, 32'h00000000} /* (27, 7, 28) {real, imag} */,
  {32'h443f6fbb, 32'h00000000} /* (27, 7, 27) {real, imag} */,
  {32'h43b4ba81, 32'h00000000} /* (27, 7, 26) {real, imag} */,
  {32'h44b5a4fc, 32'h00000000} /* (27, 7, 25) {real, imag} */,
  {32'h44463ac1, 32'h00000000} /* (27, 7, 24) {real, imag} */,
  {32'h44a67fb9, 32'h00000000} /* (27, 7, 23) {real, imag} */,
  {32'h448e8c15, 32'h00000000} /* (27, 7, 22) {real, imag} */,
  {32'h43da13ac, 32'h00000000} /* (27, 7, 21) {real, imag} */,
  {32'hc45e1e8f, 32'h00000000} /* (27, 7, 20) {real, imag} */,
  {32'hc505ed73, 32'h00000000} /* (27, 7, 19) {real, imag} */,
  {32'hc50b2c0a, 32'h00000000} /* (27, 7, 18) {real, imag} */,
  {32'hc54e3f0b, 32'h00000000} /* (27, 7, 17) {real, imag} */,
  {32'hc523d03c, 32'h00000000} /* (27, 7, 16) {real, imag} */,
  {32'hc5134526, 32'h00000000} /* (27, 7, 15) {real, imag} */,
  {32'hc5359530, 32'h00000000} /* (27, 7, 14) {real, imag} */,
  {32'hc51a85a7, 32'h00000000} /* (27, 7, 13) {real, imag} */,
  {32'hc4bfef81, 32'h00000000} /* (27, 7, 12) {real, imag} */,
  {32'hc4bac7fc, 32'h00000000} /* (27, 7, 11) {real, imag} */,
  {32'hc45ecf70, 32'h00000000} /* (27, 7, 10) {real, imag} */,
  {32'h4455e660, 32'h00000000} /* (27, 7, 9) {real, imag} */,
  {32'h44b4830e, 32'h00000000} /* (27, 7, 8) {real, imag} */,
  {32'h44ebf9bd, 32'h00000000} /* (27, 7, 7) {real, imag} */,
  {32'h449ba5e7, 32'h00000000} /* (27, 7, 6) {real, imag} */,
  {32'h4526339a, 32'h00000000} /* (27, 7, 5) {real, imag} */,
  {32'h44f6164c, 32'h00000000} /* (27, 7, 4) {real, imag} */,
  {32'h448f9c38, 32'h00000000} /* (27, 7, 3) {real, imag} */,
  {32'h44c4aa84, 32'h00000000} /* (27, 7, 2) {real, imag} */,
  {32'h44516a94, 32'h00000000} /* (27, 7, 1) {real, imag} */,
  {32'h43af34ac, 32'h00000000} /* (27, 7, 0) {real, imag} */,
  {32'hc3877682, 32'h00000000} /* (27, 6, 31) {real, imag} */,
  {32'hc30dc0d0, 32'h00000000} /* (27, 6, 30) {real, imag} */,
  {32'hc3729468, 32'h00000000} /* (27, 6, 29) {real, imag} */,
  {32'hc35de438, 32'h00000000} /* (27, 6, 28) {real, imag} */,
  {32'h442ad5c7, 32'h00000000} /* (27, 6, 27) {real, imag} */,
  {32'h44624e0a, 32'h00000000} /* (27, 6, 26) {real, imag} */,
  {32'h44a8456d, 32'h00000000} /* (27, 6, 25) {real, imag} */,
  {32'h443f534f, 32'h00000000} /* (27, 6, 24) {real, imag} */,
  {32'h440e776f, 32'h00000000} /* (27, 6, 23) {real, imag} */,
  {32'h449bc98e, 32'h00000000} /* (27, 6, 22) {real, imag} */,
  {32'h44bba008, 32'h00000000} /* (27, 6, 21) {real, imag} */,
  {32'hc40ce24b, 32'h00000000} /* (27, 6, 20) {real, imag} */,
  {32'hc4bd285c, 32'h00000000} /* (27, 6, 19) {real, imag} */,
  {32'hc50b0420, 32'h00000000} /* (27, 6, 18) {real, imag} */,
  {32'hc4bd0296, 32'h00000000} /* (27, 6, 17) {real, imag} */,
  {32'hc4a99570, 32'h00000000} /* (27, 6, 16) {real, imag} */,
  {32'hc5004c15, 32'h00000000} /* (27, 6, 15) {real, imag} */,
  {32'hc522012f, 32'h00000000} /* (27, 6, 14) {real, imag} */,
  {32'hc55dfa7e, 32'h00000000} /* (27, 6, 13) {real, imag} */,
  {32'hc4e03950, 32'h00000000} /* (27, 6, 12) {real, imag} */,
  {32'hc4b7efea, 32'h00000000} /* (27, 6, 11) {real, imag} */,
  {32'h438d48ab, 32'h00000000} /* (27, 6, 10) {real, imag} */,
  {32'h44d5677b, 32'h00000000} /* (27, 6, 9) {real, imag} */,
  {32'h4439405f, 32'h00000000} /* (27, 6, 8) {real, imag} */,
  {32'h44c6b576, 32'h00000000} /* (27, 6, 7) {real, imag} */,
  {32'h44bc1fba, 32'h00000000} /* (27, 6, 6) {real, imag} */,
  {32'h450c10f3, 32'h00000000} /* (27, 6, 5) {real, imag} */,
  {32'h44eb9876, 32'h00000000} /* (27, 6, 4) {real, imag} */,
  {32'h44764f14, 32'h00000000} /* (27, 6, 3) {real, imag} */,
  {32'h44820d85, 32'h00000000} /* (27, 6, 2) {real, imag} */,
  {32'h44e19e9e, 32'h00000000} /* (27, 6, 1) {real, imag} */,
  {32'h4325c8b4, 32'h00000000} /* (27, 6, 0) {real, imag} */,
  {32'hc4163c2e, 32'h00000000} /* (27, 5, 31) {real, imag} */,
  {32'h41f66fc0, 32'h00000000} /* (27, 5, 30) {real, imag} */,
  {32'h42d97630, 32'h00000000} /* (27, 5, 29) {real, imag} */,
  {32'h42ec9890, 32'h00000000} /* (27, 5, 28) {real, imag} */,
  {32'h42807a98, 32'h00000000} /* (27, 5, 27) {real, imag} */,
  {32'h442c83ce, 32'h00000000} /* (27, 5, 26) {real, imag} */,
  {32'h44ce0f66, 32'h00000000} /* (27, 5, 25) {real, imag} */,
  {32'h4436b47f, 32'h00000000} /* (27, 5, 24) {real, imag} */,
  {32'h435ad988, 32'h00000000} /* (27, 5, 23) {real, imag} */,
  {32'h44dc3416, 32'h00000000} /* (27, 5, 22) {real, imag} */,
  {32'h44a2fe16, 32'h00000000} /* (27, 5, 21) {real, imag} */,
  {32'h4491c0d1, 32'h00000000} /* (27, 5, 20) {real, imag} */,
  {32'hc25a7c70, 32'h00000000} /* (27, 5, 19) {real, imag} */,
  {32'hc3e2732f, 32'h00000000} /* (27, 5, 18) {real, imag} */,
  {32'hc3e5e19a, 32'h00000000} /* (27, 5, 17) {real, imag} */,
  {32'hc4830281, 32'h00000000} /* (27, 5, 16) {real, imag} */,
  {32'hc4a39369, 32'h00000000} /* (27, 5, 15) {real, imag} */,
  {32'hc5364b3e, 32'h00000000} /* (27, 5, 14) {real, imag} */,
  {32'hc50dac14, 32'h00000000} /* (27, 5, 13) {real, imag} */,
  {32'hc4ed39f5, 32'h00000000} /* (27, 5, 12) {real, imag} */,
  {32'hc4d71b94, 32'h00000000} /* (27, 5, 11) {real, imag} */,
  {32'hc3dca4fd, 32'h00000000} /* (27, 5, 10) {real, imag} */,
  {32'h430a32c0, 32'h00000000} /* (27, 5, 9) {real, imag} */,
  {32'hc3f139d6, 32'h00000000} /* (27, 5, 8) {real, imag} */,
  {32'hc31b17a8, 32'h00000000} /* (27, 5, 7) {real, imag} */,
  {32'h43f4e4f0, 32'h00000000} /* (27, 5, 6) {real, imag} */,
  {32'h44583f94, 32'h00000000} /* (27, 5, 5) {real, imag} */,
  {32'h446cb362, 32'h00000000} /* (27, 5, 4) {real, imag} */,
  {32'h4482eaf2, 32'h00000000} /* (27, 5, 3) {real, imag} */,
  {32'h44980fc0, 32'h00000000} /* (27, 5, 2) {real, imag} */,
  {32'h44047ae8, 32'h00000000} /* (27, 5, 1) {real, imag} */,
  {32'h42849f80, 32'h00000000} /* (27, 5, 0) {real, imag} */,
  {32'hc42eb8ce, 32'h00000000} /* (27, 4, 31) {real, imag} */,
  {32'hc404c21a, 32'h00000000} /* (27, 4, 30) {real, imag} */,
  {32'hc3fd47f4, 32'h00000000} /* (27, 4, 29) {real, imag} */,
  {32'h436707b4, 32'h00000000} /* (27, 4, 28) {real, imag} */,
  {32'hc3b7a1b8, 32'h00000000} /* (27, 4, 27) {real, imag} */,
  {32'hc48d4e8f, 32'h00000000} /* (27, 4, 26) {real, imag} */,
  {32'hc452d40a, 32'h00000000} /* (27, 4, 25) {real, imag} */,
  {32'h434bc58c, 32'h00000000} /* (27, 4, 24) {real, imag} */,
  {32'h4483e172, 32'h00000000} /* (27, 4, 23) {real, imag} */,
  {32'h44b229aa, 32'h00000000} /* (27, 4, 22) {real, imag} */,
  {32'h448ddeec, 32'h00000000} /* (27, 4, 21) {real, imag} */,
  {32'h44f741cb, 32'h00000000} /* (27, 4, 20) {real, imag} */,
  {32'h4439b8e0, 32'h00000000} /* (27, 4, 19) {real, imag} */,
  {32'h44736b70, 32'h00000000} /* (27, 4, 18) {real, imag} */,
  {32'h44b016b0, 32'h00000000} /* (27, 4, 17) {real, imag} */,
  {32'h445f3b91, 32'h00000000} /* (27, 4, 16) {real, imag} */,
  {32'hc4586266, 32'h00000000} /* (27, 4, 15) {real, imag} */,
  {32'hc4df7393, 32'h00000000} /* (27, 4, 14) {real, imag} */,
  {32'hc5190a4e, 32'h00000000} /* (27, 4, 13) {real, imag} */,
  {32'hc4ecfb30, 32'h00000000} /* (27, 4, 12) {real, imag} */,
  {32'hc504a80f, 32'h00000000} /* (27, 4, 11) {real, imag} */,
  {32'hc4f63319, 32'h00000000} /* (27, 4, 10) {real, imag} */,
  {32'hc4a24447, 32'h00000000} /* (27, 4, 9) {real, imag} */,
  {32'hc4d990d8, 32'h00000000} /* (27, 4, 8) {real, imag} */,
  {32'hc46f2bde, 32'h00000000} /* (27, 4, 7) {real, imag} */,
  {32'hc452b0d8, 32'h00000000} /* (27, 4, 6) {real, imag} */,
  {32'h44c3fffc, 32'h00000000} /* (27, 4, 5) {real, imag} */,
  {32'h44b2c3c9, 32'h00000000} /* (27, 4, 4) {real, imag} */,
  {32'h44c142a8, 32'h00000000} /* (27, 4, 3) {real, imag} */,
  {32'h4459ba56, 32'h00000000} /* (27, 4, 2) {real, imag} */,
  {32'h420b3e00, 32'h00000000} /* (27, 4, 1) {real, imag} */,
  {32'hc3efb42e, 32'h00000000} /* (27, 4, 0) {real, imag} */,
  {32'hc47a2534, 32'h00000000} /* (27, 3, 31) {real, imag} */,
  {32'h438e2328, 32'h00000000} /* (27, 3, 30) {real, imag} */,
  {32'h4363eb80, 32'h00000000} /* (27, 3, 29) {real, imag} */,
  {32'h433fae98, 32'h00000000} /* (27, 3, 28) {real, imag} */,
  {32'h432dbd38, 32'h00000000} /* (27, 3, 27) {real, imag} */,
  {32'hc42c2167, 32'h00000000} /* (27, 3, 26) {real, imag} */,
  {32'hc3819c9e, 32'h00000000} /* (27, 3, 25) {real, imag} */,
  {32'h432153a0, 32'h00000000} /* (27, 3, 24) {real, imag} */,
  {32'h4453a268, 32'h00000000} /* (27, 3, 23) {real, imag} */,
  {32'h446bb628, 32'h00000000} /* (27, 3, 22) {real, imag} */,
  {32'h44fbb2d8, 32'h00000000} /* (27, 3, 21) {real, imag} */,
  {32'h44fba37e, 32'h00000000} /* (27, 3, 20) {real, imag} */,
  {32'h450d6752, 32'h00000000} /* (27, 3, 19) {real, imag} */,
  {32'h44d554bc, 32'h00000000} /* (27, 3, 18) {real, imag} */,
  {32'h44d9f714, 32'h00000000} /* (27, 3, 17) {real, imag} */,
  {32'h444cef37, 32'h00000000} /* (27, 3, 16) {real, imag} */,
  {32'hc42631f0, 32'h00000000} /* (27, 3, 15) {real, imag} */,
  {32'hc3f21f5c, 32'h00000000} /* (27, 3, 14) {real, imag} */,
  {32'hc52019e8, 32'h00000000} /* (27, 3, 13) {real, imag} */,
  {32'hc5068dec, 32'h00000000} /* (27, 3, 12) {real, imag} */,
  {32'hc50f0814, 32'h00000000} /* (27, 3, 11) {real, imag} */,
  {32'hc509637f, 32'h00000000} /* (27, 3, 10) {real, imag} */,
  {32'hc4eecbf4, 32'h00000000} /* (27, 3, 9) {real, imag} */,
  {32'hc4b54f8a, 32'h00000000} /* (27, 3, 8) {real, imag} */,
  {32'hc4d2e7ee, 32'h00000000} /* (27, 3, 7) {real, imag} */,
  {32'hc4983e32, 32'h00000000} /* (27, 3, 6) {real, imag} */,
  {32'h432e2ea0, 32'h00000000} /* (27, 3, 5) {real, imag} */,
  {32'h43e9f182, 32'h00000000} /* (27, 3, 4) {real, imag} */,
  {32'h4430178a, 32'h00000000} /* (27, 3, 3) {real, imag} */,
  {32'h4483ed92, 32'h00000000} /* (27, 3, 2) {real, imag} */,
  {32'h43ed8512, 32'h00000000} /* (27, 3, 1) {real, imag} */,
  {32'hc32f9c04, 32'h00000000} /* (27, 3, 0) {real, imag} */,
  {32'hc4840bd0, 32'h00000000} /* (27, 2, 31) {real, imag} */,
  {32'hc2a55be8, 32'h00000000} /* (27, 2, 30) {real, imag} */,
  {32'hc407de92, 32'h00000000} /* (27, 2, 29) {real, imag} */,
  {32'hc35847b8, 32'h00000000} /* (27, 2, 28) {real, imag} */,
  {32'hc37d2e90, 32'h00000000} /* (27, 2, 27) {real, imag} */,
  {32'hc3435730, 32'h00000000} /* (27, 2, 26) {real, imag} */,
  {32'hc3ddb054, 32'h00000000} /* (27, 2, 25) {real, imag} */,
  {32'h444f2425, 32'h00000000} /* (27, 2, 24) {real, imag} */,
  {32'h442b803b, 32'h00000000} /* (27, 2, 23) {real, imag} */,
  {32'h44893382, 32'h00000000} /* (27, 2, 22) {real, imag} */,
  {32'h4525c484, 32'h00000000} /* (27, 2, 21) {real, imag} */,
  {32'h4507b310, 32'h00000000} /* (27, 2, 20) {real, imag} */,
  {32'h4532fed3, 32'h00000000} /* (27, 2, 19) {real, imag} */,
  {32'h449b11d2, 32'h00000000} /* (27, 2, 18) {real, imag} */,
  {32'h450ab54a, 32'h00000000} /* (27, 2, 17) {real, imag} */,
  {32'h44cc27b4, 32'h00000000} /* (27, 2, 16) {real, imag} */,
  {32'hc4a09430, 32'h00000000} /* (27, 2, 15) {real, imag} */,
  {32'hc4a21fca, 32'h00000000} /* (27, 2, 14) {real, imag} */,
  {32'hc4d0b393, 32'h00000000} /* (27, 2, 13) {real, imag} */,
  {32'hc517bc32, 32'h00000000} /* (27, 2, 12) {real, imag} */,
  {32'hc52669f8, 32'h00000000} /* (27, 2, 11) {real, imag} */,
  {32'hc53ce4a7, 32'h00000000} /* (27, 2, 10) {real, imag} */,
  {32'hc52e4022, 32'h00000000} /* (27, 2, 9) {real, imag} */,
  {32'hc51acb0d, 32'h00000000} /* (27, 2, 8) {real, imag} */,
  {32'hc4c4f290, 32'h00000000} /* (27, 2, 7) {real, imag} */,
  {32'hc504f021, 32'h00000000} /* (27, 2, 6) {real, imag} */,
  {32'hc4663eca, 32'h00000000} /* (27, 2, 5) {real, imag} */,
  {32'hc2f34cb0, 32'h00000000} /* (27, 2, 4) {real, imag} */,
  {32'h43f9ffc0, 32'h00000000} /* (27, 2, 3) {real, imag} */,
  {32'h448ec576, 32'h00000000} /* (27, 2, 2) {real, imag} */,
  {32'h444c10b8, 32'h00000000} /* (27, 2, 1) {real, imag} */,
  {32'hc3bb7452, 32'h00000000} /* (27, 2, 0) {real, imag} */,
  {32'hc3ca552e, 32'h00000000} /* (27, 1, 31) {real, imag} */,
  {32'h43f065a4, 32'h00000000} /* (27, 1, 30) {real, imag} */,
  {32'hc3f54790, 32'h00000000} /* (27, 1, 29) {real, imag} */,
  {32'hc4895a54, 32'h00000000} /* (27, 1, 28) {real, imag} */,
  {32'hc1f5e500, 32'h00000000} /* (27, 1, 27) {real, imag} */,
  {32'hc4869d04, 32'h00000000} /* (27, 1, 26) {real, imag} */,
  {32'h44245092, 32'h00000000} /* (27, 1, 25) {real, imag} */,
  {32'h43961a7c, 32'h00000000} /* (27, 1, 24) {real, imag} */,
  {32'h4476bfb5, 32'h00000000} /* (27, 1, 23) {real, imag} */,
  {32'h45082d04, 32'h00000000} /* (27, 1, 22) {real, imag} */,
  {32'h44f3c297, 32'h00000000} /* (27, 1, 21) {real, imag} */,
  {32'h44af47a4, 32'h00000000} /* (27, 1, 20) {real, imag} */,
  {32'h4527afe6, 32'h00000000} /* (27, 1, 19) {real, imag} */,
  {32'h451c001a, 32'h00000000} /* (27, 1, 18) {real, imag} */,
  {32'h45058242, 32'h00000000} /* (27, 1, 17) {real, imag} */,
  {32'h44d69660, 32'h00000000} /* (27, 1, 16) {real, imag} */,
  {32'hc4531f47, 32'h00000000} /* (27, 1, 15) {real, imag} */,
  {32'hc4e2307d, 32'h00000000} /* (27, 1, 14) {real, imag} */,
  {32'hc4f8ec2c, 32'h00000000} /* (27, 1, 13) {real, imag} */,
  {32'hc539596e, 32'h00000000} /* (27, 1, 12) {real, imag} */,
  {32'hc53d37b4, 32'h00000000} /* (27, 1, 11) {real, imag} */,
  {32'hc51927c3, 32'h00000000} /* (27, 1, 10) {real, imag} */,
  {32'hc54fb36c, 32'h00000000} /* (27, 1, 9) {real, imag} */,
  {32'hc562a200, 32'h00000000} /* (27, 1, 8) {real, imag} */,
  {32'hc505ef7a, 32'h00000000} /* (27, 1, 7) {real, imag} */,
  {32'hc4f45cc8, 32'h00000000} /* (27, 1, 6) {real, imag} */,
  {32'hc4771d36, 32'h00000000} /* (27, 1, 5) {real, imag} */,
  {32'hc30a97c0, 32'h00000000} /* (27, 1, 4) {real, imag} */,
  {32'h42feefb0, 32'h00000000} /* (27, 1, 3) {real, imag} */,
  {32'h442d62e4, 32'h00000000} /* (27, 1, 2) {real, imag} */,
  {32'h443feb1a, 32'h00000000} /* (27, 1, 1) {real, imag} */,
  {32'h41db14e0, 32'h00000000} /* (27, 1, 0) {real, imag} */,
  {32'hc4adb52b, 32'h00000000} /* (27, 0, 31) {real, imag} */,
  {32'hc4935f4e, 32'h00000000} /* (27, 0, 30) {real, imag} */,
  {32'hc48ede01, 32'h00000000} /* (27, 0, 29) {real, imag} */,
  {32'hc4b144d2, 32'h00000000} /* (27, 0, 28) {real, imag} */,
  {32'hc4892967, 32'h00000000} /* (27, 0, 27) {real, imag} */,
  {32'hc453ba6b, 32'h00000000} /* (27, 0, 26) {real, imag} */,
  {32'hc3f45612, 32'h00000000} /* (27, 0, 25) {real, imag} */,
  {32'h41f4d840, 32'h00000000} /* (27, 0, 24) {real, imag} */,
  {32'h43a5ff78, 32'h00000000} /* (27, 0, 23) {real, imag} */,
  {32'h44966aa2, 32'h00000000} /* (27, 0, 22) {real, imag} */,
  {32'h441652e5, 32'h00000000} /* (27, 0, 21) {real, imag} */,
  {32'h43dc5f64, 32'h00000000} /* (27, 0, 20) {real, imag} */,
  {32'h449ce2bc, 32'h00000000} /* (27, 0, 19) {real, imag} */,
  {32'h45019bd8, 32'h00000000} /* (27, 0, 18) {real, imag} */,
  {32'h444041f0, 32'h00000000} /* (27, 0, 17) {real, imag} */,
  {32'hc358b704, 32'h00000000} /* (27, 0, 16) {real, imag} */,
  {32'hc46c71da, 32'h00000000} /* (27, 0, 15) {real, imag} */,
  {32'hc4ace716, 32'h00000000} /* (27, 0, 14) {real, imag} */,
  {32'hc4e532e1, 32'h00000000} /* (27, 0, 13) {real, imag} */,
  {32'hc500c17b, 32'h00000000} /* (27, 0, 12) {real, imag} */,
  {32'hc4d13643, 32'h00000000} /* (27, 0, 11) {real, imag} */,
  {32'hc4bc60c8, 32'h00000000} /* (27, 0, 10) {real, imag} */,
  {32'hc47da8a7, 32'h00000000} /* (27, 0, 9) {real, imag} */,
  {32'hc4d5784e, 32'h00000000} /* (27, 0, 8) {real, imag} */,
  {32'hc4c698ae, 32'h00000000} /* (27, 0, 7) {real, imag} */,
  {32'hc4cace24, 32'h00000000} /* (27, 0, 6) {real, imag} */,
  {32'hc4593951, 32'h00000000} /* (27, 0, 5) {real, imag} */,
  {32'hc3915024, 32'h00000000} /* (27, 0, 4) {real, imag} */,
  {32'h4349640c, 32'h00000000} /* (27, 0, 3) {real, imag} */,
  {32'hc3f2d204, 32'h00000000} /* (27, 0, 2) {real, imag} */,
  {32'hc4595688, 32'h00000000} /* (27, 0, 1) {real, imag} */,
  {32'hc48f5b96, 32'h00000000} /* (27, 0, 0) {real, imag} */,
  {32'hc5802176, 32'h00000000} /* (26, 31, 31) {real, imag} */,
  {32'hc5926f12, 32'h00000000} /* (26, 31, 30) {real, imag} */,
  {32'hc5830a2a, 32'h00000000} /* (26, 31, 29) {real, imag} */,
  {32'hc5809281, 32'h00000000} /* (26, 31, 28) {real, imag} */,
  {32'hc54e9560, 32'h00000000} /* (26, 31, 27) {real, imag} */,
  {32'hc558c4d6, 32'h00000000} /* (26, 31, 26) {real, imag} */,
  {32'hc5544017, 32'h00000000} /* (26, 31, 25) {real, imag} */,
  {32'hc525ed60, 32'h00000000} /* (26, 31, 24) {real, imag} */,
  {32'hc53d5201, 32'h00000000} /* (26, 31, 23) {real, imag} */,
  {32'hc51491e3, 32'h00000000} /* (26, 31, 22) {real, imag} */,
  {32'hc4e3db2b, 32'h00000000} /* (26, 31, 21) {real, imag} */,
  {32'hc51a9a75, 32'h00000000} /* (26, 31, 20) {real, imag} */,
  {32'hc3cf0f80, 32'h00000000} /* (26, 31, 19) {real, imag} */,
  {32'h42723360, 32'h00000000} /* (26, 31, 18) {real, imag} */,
  {32'h437f0230, 32'h00000000} /* (26, 31, 17) {real, imag} */,
  {32'h42729900, 32'h00000000} /* (26, 31, 16) {real, imag} */,
  {32'h4381ddb4, 32'h00000000} /* (26, 31, 15) {real, imag} */,
  {32'hc3c45370, 32'h00000000} /* (26, 31, 14) {real, imag} */,
  {32'hc3a25bc0, 32'h00000000} /* (26, 31, 13) {real, imag} */,
  {32'h438e0b80, 32'h00000000} /* (26, 31, 12) {real, imag} */,
  {32'hc373e6d0, 32'h00000000} /* (26, 31, 11) {real, imag} */,
  {32'hc3958f8c, 32'h00000000} /* (26, 31, 10) {real, imag} */,
  {32'hc42e8d3c, 32'h00000000} /* (26, 31, 9) {real, imag} */,
  {32'hc498cf76, 32'h00000000} /* (26, 31, 8) {real, imag} */,
  {32'hc481d0dc, 32'h00000000} /* (26, 31, 7) {real, imag} */,
  {32'hc4b6b1d6, 32'h00000000} /* (26, 31, 6) {real, imag} */,
  {32'hc4911fcd, 32'h00000000} /* (26, 31, 5) {real, imag} */,
  {32'hc523c061, 32'h00000000} /* (26, 31, 4) {real, imag} */,
  {32'hc5109e27, 32'h00000000} /* (26, 31, 3) {real, imag} */,
  {32'hc51f4226, 32'h00000000} /* (26, 31, 2) {real, imag} */,
  {32'hc537e965, 32'h00000000} /* (26, 31, 1) {real, imag} */,
  {32'hc52d12f9, 32'h00000000} /* (26, 31, 0) {real, imag} */,
  {32'hc56d8680, 32'h00000000} /* (26, 30, 31) {real, imag} */,
  {32'hc56da2c1, 32'h00000000} /* (26, 30, 30) {real, imag} */,
  {32'hc56f9ce2, 32'h00000000} /* (26, 30, 29) {real, imag} */,
  {32'hc5712a3c, 32'h00000000} /* (26, 30, 28) {real, imag} */,
  {32'hc529cdb4, 32'h00000000} /* (26, 30, 27) {real, imag} */,
  {32'hc55d5dcd, 32'h00000000} /* (26, 30, 26) {real, imag} */,
  {32'hc559d1f4, 32'h00000000} /* (26, 30, 25) {real, imag} */,
  {32'hc52c8f20, 32'h00000000} /* (26, 30, 24) {real, imag} */,
  {32'hc5005705, 32'h00000000} /* (26, 30, 23) {real, imag} */,
  {32'hc509001f, 32'h00000000} /* (26, 30, 22) {real, imag} */,
  {32'hc4c67416, 32'h00000000} /* (26, 30, 21) {real, imag} */,
  {32'hc49362dc, 32'h00000000} /* (26, 30, 20) {real, imag} */,
  {32'hc43ea947, 32'h00000000} /* (26, 30, 19) {real, imag} */,
  {32'h4422a3e0, 32'h00000000} /* (26, 30, 18) {real, imag} */,
  {32'hc413d256, 32'h00000000} /* (26, 30, 17) {real, imag} */,
  {32'h42c873a0, 32'h00000000} /* (26, 30, 16) {real, imag} */,
  {32'h4380de50, 32'h00000000} /* (26, 30, 15) {real, imag} */,
  {32'hc3e1ccd8, 32'h00000000} /* (26, 30, 14) {real, imag} */,
  {32'hc38ebf30, 32'h00000000} /* (26, 30, 13) {real, imag} */,
  {32'hc29379f0, 32'h00000000} /* (26, 30, 12) {real, imag} */,
  {32'hc3dda188, 32'h00000000} /* (26, 30, 11) {real, imag} */,
  {32'h4358bde0, 32'h00000000} /* (26, 30, 10) {real, imag} */,
  {32'hc4901f28, 32'h00000000} /* (26, 30, 9) {real, imag} */,
  {32'hc4cdaf77, 32'h00000000} /* (26, 30, 8) {real, imag} */,
  {32'hc48687ea, 32'h00000000} /* (26, 30, 7) {real, imag} */,
  {32'hc392cf9e, 32'h00000000} /* (26, 30, 6) {real, imag} */,
  {32'hc494abe2, 32'h00000000} /* (26, 30, 5) {real, imag} */,
  {32'hc4b1d9d0, 32'h00000000} /* (26, 30, 4) {real, imag} */,
  {32'hc516b389, 32'h00000000} /* (26, 30, 3) {real, imag} */,
  {32'hc525ee09, 32'h00000000} /* (26, 30, 2) {real, imag} */,
  {32'hc55f3f1e, 32'h00000000} /* (26, 30, 1) {real, imag} */,
  {32'hc55c913e, 32'h00000000} /* (26, 30, 0) {real, imag} */,
  {32'hc51e5155, 32'h00000000} /* (26, 29, 31) {real, imag} */,
  {32'hc53bbc16, 32'h00000000} /* (26, 29, 30) {real, imag} */,
  {32'hc5907a92, 32'h00000000} /* (26, 29, 29) {real, imag} */,
  {32'hc55ca87c, 32'h00000000} /* (26, 29, 28) {real, imag} */,
  {32'hc546aebf, 32'h00000000} /* (26, 29, 27) {real, imag} */,
  {32'hc56c5cc8, 32'h00000000} /* (26, 29, 26) {real, imag} */,
  {32'hc5721a1f, 32'h00000000} /* (26, 29, 25) {real, imag} */,
  {32'hc53356f7, 32'h00000000} /* (26, 29, 24) {real, imag} */,
  {32'hc509fec2, 32'h00000000} /* (26, 29, 23) {real, imag} */,
  {32'hc518ab18, 32'h00000000} /* (26, 29, 22) {real, imag} */,
  {32'hc4e64a28, 32'h00000000} /* (26, 29, 21) {real, imag} */,
  {32'hc447a9cd, 32'h00000000} /* (26, 29, 20) {real, imag} */,
  {32'hc3cea3dc, 32'h00000000} /* (26, 29, 19) {real, imag} */,
  {32'hc449443e, 32'h00000000} /* (26, 29, 18) {real, imag} */,
  {32'hc4237dd8, 32'h00000000} /* (26, 29, 17) {real, imag} */,
  {32'hc41681cc, 32'h00000000} /* (26, 29, 16) {real, imag} */,
  {32'hc3659d70, 32'h00000000} /* (26, 29, 15) {real, imag} */,
  {32'hc3178d78, 32'h00000000} /* (26, 29, 14) {real, imag} */,
  {32'hc4023df0, 32'h00000000} /* (26, 29, 13) {real, imag} */,
  {32'hc4890e37, 32'h00000000} /* (26, 29, 12) {real, imag} */,
  {32'hc4a9560a, 32'h00000000} /* (26, 29, 11) {real, imag} */,
  {32'h4354ad18, 32'h00000000} /* (26, 29, 10) {real, imag} */,
  {32'h44054944, 32'h00000000} /* (26, 29, 9) {real, imag} */,
  {32'hc44bef5c, 32'h00000000} /* (26, 29, 8) {real, imag} */,
  {32'hc49eded9, 32'h00000000} /* (26, 29, 7) {real, imag} */,
  {32'hc480436f, 32'h00000000} /* (26, 29, 6) {real, imag} */,
  {32'hc3cc17ae, 32'h00000000} /* (26, 29, 5) {real, imag} */,
  {32'hc4c4b6d8, 32'h00000000} /* (26, 29, 4) {real, imag} */,
  {32'hc52335c8, 32'h00000000} /* (26, 29, 3) {real, imag} */,
  {32'hc5339404, 32'h00000000} /* (26, 29, 2) {real, imag} */,
  {32'hc57d294a, 32'h00000000} /* (26, 29, 1) {real, imag} */,
  {32'hc56af197, 32'h00000000} /* (26, 29, 0) {real, imag} */,
  {32'hc5547a46, 32'h00000000} /* (26, 28, 31) {real, imag} */,
  {32'hc554bb7e, 32'h00000000} /* (26, 28, 30) {real, imag} */,
  {32'hc5940f5e, 32'h00000000} /* (26, 28, 29) {real, imag} */,
  {32'hc553511c, 32'h00000000} /* (26, 28, 28) {real, imag} */,
  {32'hc53891a2, 32'h00000000} /* (26, 28, 27) {real, imag} */,
  {32'hc589684e, 32'h00000000} /* (26, 28, 26) {real, imag} */,
  {32'hc587cfa5, 32'h00000000} /* (26, 28, 25) {real, imag} */,
  {32'hc51ce63f, 32'h00000000} /* (26, 28, 24) {real, imag} */,
  {32'hc507e0e4, 32'h00000000} /* (26, 28, 23) {real, imag} */,
  {32'hc506f898, 32'h00000000} /* (26, 28, 22) {real, imag} */,
  {32'hc4b0f5b8, 32'h00000000} /* (26, 28, 21) {real, imag} */,
  {32'hc4e56afb, 32'h00000000} /* (26, 28, 20) {real, imag} */,
  {32'hc4963413, 32'h00000000} /* (26, 28, 19) {real, imag} */,
  {32'hc4305b16, 32'h00000000} /* (26, 28, 18) {real, imag} */,
  {32'h43d2a818, 32'h00000000} /* (26, 28, 17) {real, imag} */,
  {32'hc49afcdc, 32'h00000000} /* (26, 28, 16) {real, imag} */,
  {32'hc5068ede, 32'h00000000} /* (26, 28, 15) {real, imag} */,
  {32'hc370d368, 32'h00000000} /* (26, 28, 14) {real, imag} */,
  {32'hc493043c, 32'h00000000} /* (26, 28, 13) {real, imag} */,
  {32'hc384f298, 32'h00000000} /* (26, 28, 12) {real, imag} */,
  {32'hc358af40, 32'h00000000} /* (26, 28, 11) {real, imag} */,
  {32'hc3bef890, 32'h00000000} /* (26, 28, 10) {real, imag} */,
  {32'hc31b4040, 32'h00000000} /* (26, 28, 9) {real, imag} */,
  {32'hc38e4a78, 32'h00000000} /* (26, 28, 8) {real, imag} */,
  {32'hc4481e1c, 32'h00000000} /* (26, 28, 7) {real, imag} */,
  {32'hc361edbc, 32'h00000000} /* (26, 28, 6) {real, imag} */,
  {32'hc4b74564, 32'h00000000} /* (26, 28, 5) {real, imag} */,
  {32'hc5123bbc, 32'h00000000} /* (26, 28, 4) {real, imag} */,
  {32'hc553c6b8, 32'h00000000} /* (26, 28, 3) {real, imag} */,
  {32'hc53e2d10, 32'h00000000} /* (26, 28, 2) {real, imag} */,
  {32'hc534f4a3, 32'h00000000} /* (26, 28, 1) {real, imag} */,
  {32'hc526722e, 32'h00000000} /* (26, 28, 0) {real, imag} */,
  {32'hc5591095, 32'h00000000} /* (26, 27, 31) {real, imag} */,
  {32'hc58be3e8, 32'h00000000} /* (26, 27, 30) {real, imag} */,
  {32'hc59ab8a2, 32'h00000000} /* (26, 27, 29) {real, imag} */,
  {32'hc541a992, 32'h00000000} /* (26, 27, 28) {real, imag} */,
  {32'hc51d57b7, 32'h00000000} /* (26, 27, 27) {real, imag} */,
  {32'hc56c50d8, 32'h00000000} /* (26, 27, 26) {real, imag} */,
  {32'hc56428fc, 32'h00000000} /* (26, 27, 25) {real, imag} */,
  {32'hc5355265, 32'h00000000} /* (26, 27, 24) {real, imag} */,
  {32'hc4ab97f3, 32'h00000000} /* (26, 27, 23) {real, imag} */,
  {32'hc4af7876, 32'h00000000} /* (26, 27, 22) {real, imag} */,
  {32'hc46bc4de, 32'h00000000} /* (26, 27, 21) {real, imag} */,
  {32'hc494d110, 32'h00000000} /* (26, 27, 20) {real, imag} */,
  {32'hc4563ee3, 32'h00000000} /* (26, 27, 19) {real, imag} */,
  {32'hc49610f4, 32'h00000000} /* (26, 27, 18) {real, imag} */,
  {32'hc4aaa83d, 32'h00000000} /* (26, 27, 17) {real, imag} */,
  {32'h43336940, 32'h00000000} /* (26, 27, 16) {real, imag} */,
  {32'hc4a92e3e, 32'h00000000} /* (26, 27, 15) {real, imag} */,
  {32'hc3af2ac8, 32'h00000000} /* (26, 27, 14) {real, imag} */,
  {32'hc38002e0, 32'h00000000} /* (26, 27, 13) {real, imag} */,
  {32'hc3afa69c, 32'h00000000} /* (26, 27, 12) {real, imag} */,
  {32'h43b34868, 32'h00000000} /* (26, 27, 11) {real, imag} */,
  {32'h43b6b3c4, 32'h00000000} /* (26, 27, 10) {real, imag} */,
  {32'hc4dae9e7, 32'h00000000} /* (26, 27, 9) {real, imag} */,
  {32'hc3908d88, 32'h00000000} /* (26, 27, 8) {real, imag} */,
  {32'hc41e2e6e, 32'h00000000} /* (26, 27, 7) {real, imag} */,
  {32'hc4609a33, 32'h00000000} /* (26, 27, 6) {real, imag} */,
  {32'hc4fba7f1, 32'h00000000} /* (26, 27, 5) {real, imag} */,
  {32'hc5292342, 32'h00000000} /* (26, 27, 4) {real, imag} */,
  {32'hc50cff1d, 32'h00000000} /* (26, 27, 3) {real, imag} */,
  {32'hc53c874e, 32'h00000000} /* (26, 27, 2) {real, imag} */,
  {32'hc533c6da, 32'h00000000} /* (26, 27, 1) {real, imag} */,
  {32'hc53a5d06, 32'h00000000} /* (26, 27, 0) {real, imag} */,
  {32'hc564671f, 32'h00000000} /* (26, 26, 31) {real, imag} */,
  {32'hc5775135, 32'h00000000} /* (26, 26, 30) {real, imag} */,
  {32'hc58fb776, 32'h00000000} /* (26, 26, 29) {real, imag} */,
  {32'hc586ddae, 32'h00000000} /* (26, 26, 28) {real, imag} */,
  {32'hc56a3156, 32'h00000000} /* (26, 26, 27) {real, imag} */,
  {32'hc54b1400, 32'h00000000} /* (26, 26, 26) {real, imag} */,
  {32'hc533fcf2, 32'h00000000} /* (26, 26, 25) {real, imag} */,
  {32'hc51021d6, 32'h00000000} /* (26, 26, 24) {real, imag} */,
  {32'hc4b58fb0, 32'h00000000} /* (26, 26, 23) {real, imag} */,
  {32'hc4bf8a4a, 32'h00000000} /* (26, 26, 22) {real, imag} */,
  {32'hc4e1027d, 32'h00000000} /* (26, 26, 21) {real, imag} */,
  {32'hc4a929b3, 32'h00000000} /* (26, 26, 20) {real, imag} */,
  {32'hc4826605, 32'h00000000} /* (26, 26, 19) {real, imag} */,
  {32'hc426951a, 32'h00000000} /* (26, 26, 18) {real, imag} */,
  {32'hc4793158, 32'h00000000} /* (26, 26, 17) {real, imag} */,
  {32'hc33e1000, 32'h00000000} /* (26, 26, 16) {real, imag} */,
  {32'hc3cb0200, 32'h00000000} /* (26, 26, 15) {real, imag} */,
  {32'hc49973aa, 32'h00000000} /* (26, 26, 14) {real, imag} */,
  {32'hc32e4170, 32'h00000000} /* (26, 26, 13) {real, imag} */,
  {32'hc46790a4, 32'h00000000} /* (26, 26, 12) {real, imag} */,
  {32'hc422f048, 32'h00000000} /* (26, 26, 11) {real, imag} */,
  {32'hc4b0bbfd, 32'h00000000} /* (26, 26, 10) {real, imag} */,
  {32'hc42a7ce6, 32'h00000000} /* (26, 26, 9) {real, imag} */,
  {32'hc49119fb, 32'h00000000} /* (26, 26, 8) {real, imag} */,
  {32'hc49dfe4e, 32'h00000000} /* (26, 26, 7) {real, imag} */,
  {32'hc4d8cb0a, 32'h00000000} /* (26, 26, 6) {real, imag} */,
  {32'hc49495d1, 32'h00000000} /* (26, 26, 5) {real, imag} */,
  {32'hc50a963e, 32'h00000000} /* (26, 26, 4) {real, imag} */,
  {32'hc52d93b6, 32'h00000000} /* (26, 26, 3) {real, imag} */,
  {32'hc529f96c, 32'h00000000} /* (26, 26, 2) {real, imag} */,
  {32'hc5897c4d, 32'h00000000} /* (26, 26, 1) {real, imag} */,
  {32'hc56d1022, 32'h00000000} /* (26, 26, 0) {real, imag} */,
  {32'hc5632917, 32'h00000000} /* (26, 25, 31) {real, imag} */,
  {32'hc589ee87, 32'h00000000} /* (26, 25, 30) {real, imag} */,
  {32'hc53e5366, 32'h00000000} /* (26, 25, 29) {real, imag} */,
  {32'hc54faf8b, 32'h00000000} /* (26, 25, 28) {real, imag} */,
  {32'hc54ed3c5, 32'h00000000} /* (26, 25, 27) {real, imag} */,
  {32'hc554b81b, 32'h00000000} /* (26, 25, 26) {real, imag} */,
  {32'hc5168dad, 32'h00000000} /* (26, 25, 25) {real, imag} */,
  {32'hc50ce41d, 32'h00000000} /* (26, 25, 24) {real, imag} */,
  {32'hc4b6d8e4, 32'h00000000} /* (26, 25, 23) {real, imag} */,
  {32'hc4866cf4, 32'h00000000} /* (26, 25, 22) {real, imag} */,
  {32'hc455110f, 32'h00000000} /* (26, 25, 21) {real, imag} */,
  {32'hc35f0bdc, 32'h00000000} /* (26, 25, 20) {real, imag} */,
  {32'h43778658, 32'h00000000} /* (26, 25, 19) {real, imag} */,
  {32'hc45d9716, 32'h00000000} /* (26, 25, 18) {real, imag} */,
  {32'hc42c350e, 32'h00000000} /* (26, 25, 17) {real, imag} */,
  {32'h43a23498, 32'h00000000} /* (26, 25, 16) {real, imag} */,
  {32'hc4443614, 32'h00000000} /* (26, 25, 15) {real, imag} */,
  {32'hc4097cb6, 32'h00000000} /* (26, 25, 14) {real, imag} */,
  {32'hc336ffa8, 32'h00000000} /* (26, 25, 13) {real, imag} */,
  {32'h42603b00, 32'h00000000} /* (26, 25, 12) {real, imag} */,
  {32'hc4ad50da, 32'h00000000} /* (26, 25, 11) {real, imag} */,
  {32'hc434d1ec, 32'h00000000} /* (26, 25, 10) {real, imag} */,
  {32'hc410def5, 32'h00000000} /* (26, 25, 9) {real, imag} */,
  {32'hc343a830, 32'h00000000} /* (26, 25, 8) {real, imag} */,
  {32'hc4252198, 32'h00000000} /* (26, 25, 7) {real, imag} */,
  {32'hc499e670, 32'h00000000} /* (26, 25, 6) {real, imag} */,
  {32'hc4a4b548, 32'h00000000} /* (26, 25, 5) {real, imag} */,
  {32'hc4cc12de, 32'h00000000} /* (26, 25, 4) {real, imag} */,
  {32'hc521d6e8, 32'h00000000} /* (26, 25, 3) {real, imag} */,
  {32'hc541afc4, 32'h00000000} /* (26, 25, 2) {real, imag} */,
  {32'hc54a351a, 32'h00000000} /* (26, 25, 1) {real, imag} */,
  {32'hc5435c13, 32'h00000000} /* (26, 25, 0) {real, imag} */,
  {32'hc531e59f, 32'h00000000} /* (26, 24, 31) {real, imag} */,
  {32'hc539e0c0, 32'h00000000} /* (26, 24, 30) {real, imag} */,
  {32'hc502a5ac, 32'h00000000} /* (26, 24, 29) {real, imag} */,
  {32'hc53d428f, 32'h00000000} /* (26, 24, 28) {real, imag} */,
  {32'hc4d70bb5, 32'h00000000} /* (26, 24, 27) {real, imag} */,
  {32'hc50e0b76, 32'h00000000} /* (26, 24, 26) {real, imag} */,
  {32'hc50a4d36, 32'h00000000} /* (26, 24, 25) {real, imag} */,
  {32'hc41b7dfb, 32'h00000000} /* (26, 24, 24) {real, imag} */,
  {32'hc4e71f07, 32'h00000000} /* (26, 24, 23) {real, imag} */,
  {32'hc464d11c, 32'h00000000} /* (26, 24, 22) {real, imag} */,
  {32'hc45c91f0, 32'h00000000} /* (26, 24, 21) {real, imag} */,
  {32'h431a65a0, 32'h00000000} /* (26, 24, 20) {real, imag} */,
  {32'hc1344380, 32'h00000000} /* (26, 24, 19) {real, imag} */,
  {32'h4373dc70, 32'h00000000} /* (26, 24, 18) {real, imag} */,
  {32'hc3e5e938, 32'h00000000} /* (26, 24, 17) {real, imag} */,
  {32'hc3448fe8, 32'h00000000} /* (26, 24, 16) {real, imag} */,
  {32'h42a64920, 32'h00000000} /* (26, 24, 15) {real, imag} */,
  {32'h43f3694c, 32'h00000000} /* (26, 24, 14) {real, imag} */,
  {32'h43e925bc, 32'h00000000} /* (26, 24, 13) {real, imag} */,
  {32'hc4d0553e, 32'h00000000} /* (26, 24, 12) {real, imag} */,
  {32'hc4786952, 32'h00000000} /* (26, 24, 11) {real, imag} */,
  {32'hc39eb65c, 32'h00000000} /* (26, 24, 10) {real, imag} */,
  {32'h43ee097c, 32'h00000000} /* (26, 24, 9) {real, imag} */,
  {32'hc2978f58, 32'h00000000} /* (26, 24, 8) {real, imag} */,
  {32'hc407f522, 32'h00000000} /* (26, 24, 7) {real, imag} */,
  {32'hc4ac3476, 32'h00000000} /* (26, 24, 6) {real, imag} */,
  {32'hc51273ed, 32'h00000000} /* (26, 24, 5) {real, imag} */,
  {32'hc541c9a2, 32'h00000000} /* (26, 24, 4) {real, imag} */,
  {32'hc511d7d4, 32'h00000000} /* (26, 24, 3) {real, imag} */,
  {32'hc51c9cc5, 32'h00000000} /* (26, 24, 2) {real, imag} */,
  {32'hc528e4ad, 32'h00000000} /* (26, 24, 1) {real, imag} */,
  {32'hc544b5fa, 32'h00000000} /* (26, 24, 0) {real, imag} */,
  {32'hc523f48c, 32'h00000000} /* (26, 23, 31) {real, imag} */,
  {32'hc511ac6e, 32'h00000000} /* (26, 23, 30) {real, imag} */,
  {32'hc5226974, 32'h00000000} /* (26, 23, 29) {real, imag} */,
  {32'hc51e7ab1, 32'h00000000} /* (26, 23, 28) {real, imag} */,
  {32'hc49f2692, 32'h00000000} /* (26, 23, 27) {real, imag} */,
  {32'hc4e837a0, 32'h00000000} /* (26, 23, 26) {real, imag} */,
  {32'hc516e92b, 32'h00000000} /* (26, 23, 25) {real, imag} */,
  {32'hc4c8877e, 32'h00000000} /* (26, 23, 24) {real, imag} */,
  {32'hc49fd904, 32'h00000000} /* (26, 23, 23) {real, imag} */,
  {32'hc3ea9864, 32'h00000000} /* (26, 23, 22) {real, imag} */,
  {32'hc3f915d8, 32'h00000000} /* (26, 23, 21) {real, imag} */,
  {32'hc2fc0d30, 32'h00000000} /* (26, 23, 20) {real, imag} */,
  {32'h43126880, 32'h00000000} /* (26, 23, 19) {real, imag} */,
  {32'hc3a3b94a, 32'h00000000} /* (26, 23, 18) {real, imag} */,
  {32'h42ffb300, 32'h00000000} /* (26, 23, 17) {real, imag} */,
  {32'hc29d2b00, 32'h00000000} /* (26, 23, 16) {real, imag} */,
  {32'h44e9192b, 32'h00000000} /* (26, 23, 15) {real, imag} */,
  {32'h440715e2, 32'h00000000} /* (26, 23, 14) {real, imag} */,
  {32'h43135b48, 32'h00000000} /* (26, 23, 13) {real, imag} */,
  {32'hc47242c1, 32'h00000000} /* (26, 23, 12) {real, imag} */,
  {32'hc4133511, 32'h00000000} /* (26, 23, 11) {real, imag} */,
  {32'h430940a4, 32'h00000000} /* (26, 23, 10) {real, imag} */,
  {32'hc3f1b678, 32'h00000000} /* (26, 23, 9) {real, imag} */,
  {32'hc0ff4180, 32'h00000000} /* (26, 23, 8) {real, imag} */,
  {32'hc3b2d95a, 32'h00000000} /* (26, 23, 7) {real, imag} */,
  {32'hc4d3093f, 32'h00000000} /* (26, 23, 6) {real, imag} */,
  {32'hc52ff225, 32'h00000000} /* (26, 23, 5) {real, imag} */,
  {32'hc528d99e, 32'h00000000} /* (26, 23, 4) {real, imag} */,
  {32'hc50d71e9, 32'h00000000} /* (26, 23, 3) {real, imag} */,
  {32'hc4c9647a, 32'h00000000} /* (26, 23, 2) {real, imag} */,
  {32'hc507113e, 32'h00000000} /* (26, 23, 1) {real, imag} */,
  {32'hc5314660, 32'h00000000} /* (26, 23, 0) {real, imag} */,
  {32'hc4a3544b, 32'h00000000} /* (26, 22, 31) {real, imag} */,
  {32'hc4baff5e, 32'h00000000} /* (26, 22, 30) {real, imag} */,
  {32'hc4d17d05, 32'h00000000} /* (26, 22, 29) {real, imag} */,
  {32'hc4be4906, 32'h00000000} /* (26, 22, 28) {real, imag} */,
  {32'hc4f6ff1d, 32'h00000000} /* (26, 22, 27) {real, imag} */,
  {32'hc4ae443a, 32'h00000000} /* (26, 22, 26) {real, imag} */,
  {32'hc48355ff, 32'h00000000} /* (26, 22, 25) {real, imag} */,
  {32'hc4ced5d3, 32'h00000000} /* (26, 22, 24) {real, imag} */,
  {32'hc3f28da6, 32'h00000000} /* (26, 22, 23) {real, imag} */,
  {32'hc246b610, 32'h00000000} /* (26, 22, 22) {real, imag} */,
  {32'hc3aa8b70, 32'h00000000} /* (26, 22, 21) {real, imag} */,
  {32'hc4684e2e, 32'h00000000} /* (26, 22, 20) {real, imag} */,
  {32'hc455b45b, 32'h00000000} /* (26, 22, 19) {real, imag} */,
  {32'h4434ef7a, 32'h00000000} /* (26, 22, 18) {real, imag} */,
  {32'h4423f71a, 32'h00000000} /* (26, 22, 17) {real, imag} */,
  {32'h4438a3b0, 32'h00000000} /* (26, 22, 16) {real, imag} */,
  {32'h44a5c571, 32'h00000000} /* (26, 22, 15) {real, imag} */,
  {32'h4459041c, 32'h00000000} /* (26, 22, 14) {real, imag} */,
  {32'h43c1343c, 32'h00000000} /* (26, 22, 13) {real, imag} */,
  {32'h44878c14, 32'h00000000} /* (26, 22, 12) {real, imag} */,
  {32'h44220b9a, 32'h00000000} /* (26, 22, 11) {real, imag} */,
  {32'h44214478, 32'h00000000} /* (26, 22, 10) {real, imag} */,
  {32'hc3e35b8c, 32'h00000000} /* (26, 22, 9) {real, imag} */,
  {32'h43e99484, 32'h00000000} /* (26, 22, 8) {real, imag} */,
  {32'h4306ee90, 32'h00000000} /* (26, 22, 7) {real, imag} */,
  {32'hc428dc91, 32'h00000000} /* (26, 22, 6) {real, imag} */,
  {32'hc4b7dcce, 32'h00000000} /* (26, 22, 5) {real, imag} */,
  {32'hc4bafcfb, 32'h00000000} /* (26, 22, 4) {real, imag} */,
  {32'hc44e775d, 32'h00000000} /* (26, 22, 3) {real, imag} */,
  {32'hc45bda0c, 32'h00000000} /* (26, 22, 2) {real, imag} */,
  {32'hc48913f5, 32'h00000000} /* (26, 22, 1) {real, imag} */,
  {32'hc4b03028, 32'h00000000} /* (26, 22, 0) {real, imag} */,
  {32'hc48427f0, 32'h00000000} /* (26, 21, 31) {real, imag} */,
  {32'hc447473d, 32'h00000000} /* (26, 21, 30) {real, imag} */,
  {32'hc49e06ae, 32'h00000000} /* (26, 21, 29) {real, imag} */,
  {32'hc4e82124, 32'h00000000} /* (26, 21, 28) {real, imag} */,
  {32'hc4e43109, 32'h00000000} /* (26, 21, 27) {real, imag} */,
  {32'hc4c89f93, 32'h00000000} /* (26, 21, 26) {real, imag} */,
  {32'hc4d24aee, 32'h00000000} /* (26, 21, 25) {real, imag} */,
  {32'hc497e02c, 32'h00000000} /* (26, 21, 24) {real, imag} */,
  {32'hc4b23bda, 32'h00000000} /* (26, 21, 23) {real, imag} */,
  {32'hc3625244, 32'h00000000} /* (26, 21, 22) {real, imag} */,
  {32'h437302e2, 32'h00000000} /* (26, 21, 21) {real, imag} */,
  {32'hc3b5a15b, 32'h00000000} /* (26, 21, 20) {real, imag} */,
  {32'hc32dc814, 32'h00000000} /* (26, 21, 19) {real, imag} */,
  {32'h44c17243, 32'h00000000} /* (26, 21, 18) {real, imag} */,
  {32'h43f377a0, 32'h00000000} /* (26, 21, 17) {real, imag} */,
  {32'h4467599e, 32'h00000000} /* (26, 21, 16) {real, imag} */,
  {32'h441011b1, 32'h00000000} /* (26, 21, 15) {real, imag} */,
  {32'h4441fceb, 32'h00000000} /* (26, 21, 14) {real, imag} */,
  {32'h4498c262, 32'h00000000} /* (26, 21, 13) {real, imag} */,
  {32'h4420f9c8, 32'h00000000} /* (26, 21, 12) {real, imag} */,
  {32'hc2ca04d0, 32'h00000000} /* (26, 21, 11) {real, imag} */,
  {32'h432c1c98, 32'h00000000} /* (26, 21, 10) {real, imag} */,
  {32'hc338bac0, 32'h00000000} /* (26, 21, 9) {real, imag} */,
  {32'hc4944580, 32'h00000000} /* (26, 21, 8) {real, imag} */,
  {32'hc357ecbc, 32'h00000000} /* (26, 21, 7) {real, imag} */,
  {32'h445a6547, 32'h00000000} /* (26, 21, 6) {real, imag} */,
  {32'hc336cd0a, 32'h00000000} /* (26, 21, 5) {real, imag} */,
  {32'hc42968f2, 32'h00000000} /* (26, 21, 4) {real, imag} */,
  {32'hc41db6fe, 32'h00000000} /* (26, 21, 3) {real, imag} */,
  {32'h40c01b00, 32'h00000000} /* (26, 21, 2) {real, imag} */,
  {32'hc426107c, 32'h00000000} /* (26, 21, 1) {real, imag} */,
  {32'hc40d6e06, 32'h00000000} /* (26, 21, 0) {real, imag} */,
  {32'hc34ba25a, 32'h00000000} /* (26, 20, 31) {real, imag} */,
  {32'hc3b22496, 32'h00000000} /* (26, 20, 30) {real, imag} */,
  {32'hc40fbac4, 32'h00000000} /* (26, 20, 29) {real, imag} */,
  {32'hc10d726e, 32'h00000000} /* (26, 20, 28) {real, imag} */,
  {32'hc48fbd30, 32'h00000000} /* (26, 20, 27) {real, imag} */,
  {32'hc4860242, 32'h00000000} /* (26, 20, 26) {real, imag} */,
  {32'hc4b2fb98, 32'h00000000} /* (26, 20, 25) {real, imag} */,
  {32'hc444464d, 32'h00000000} /* (26, 20, 24) {real, imag} */,
  {32'h42aa9758, 32'h00000000} /* (26, 20, 23) {real, imag} */,
  {32'hc2709010, 32'h00000000} /* (26, 20, 22) {real, imag} */,
  {32'h42e01eb0, 32'h00000000} /* (26, 20, 21) {real, imag} */,
  {32'h423b8490, 32'h00000000} /* (26, 20, 20) {real, imag} */,
  {32'h3f860200, 32'h00000000} /* (26, 20, 19) {real, imag} */,
  {32'h442f06ea, 32'h00000000} /* (26, 20, 18) {real, imag} */,
  {32'h44057e01, 32'h00000000} /* (26, 20, 17) {real, imag} */,
  {32'h44710e65, 32'h00000000} /* (26, 20, 16) {real, imag} */,
  {32'h44389608, 32'h00000000} /* (26, 20, 15) {real, imag} */,
  {32'h441160b4, 32'h00000000} /* (26, 20, 14) {real, imag} */,
  {32'h43e5f431, 32'h00000000} /* (26, 20, 13) {real, imag} */,
  {32'h4232497c, 32'h00000000} /* (26, 20, 12) {real, imag} */,
  {32'hc2ff4898, 32'h00000000} /* (26, 20, 11) {real, imag} */,
  {32'hc4676732, 32'h00000000} /* (26, 20, 10) {real, imag} */,
  {32'hc39d8d9e, 32'h00000000} /* (26, 20, 9) {real, imag} */,
  {32'h4385e592, 32'h00000000} /* (26, 20, 8) {real, imag} */,
  {32'hc3be4960, 32'h00000000} /* (26, 20, 7) {real, imag} */,
  {32'hc44e3764, 32'h00000000} /* (26, 20, 6) {real, imag} */,
  {32'hc4dbf471, 32'h00000000} /* (26, 20, 5) {real, imag} */,
  {32'hc44f2953, 32'h00000000} /* (26, 20, 4) {real, imag} */,
  {32'hc446c1d3, 32'h00000000} /* (26, 20, 3) {real, imag} */,
  {32'hc4390428, 32'h00000000} /* (26, 20, 2) {real, imag} */,
  {32'hc41a2fe5, 32'h00000000} /* (26, 20, 1) {real, imag} */,
  {32'hc40d65a3, 32'h00000000} /* (26, 20, 0) {real, imag} */,
  {32'h438648a9, 32'h00000000} /* (26, 19, 31) {real, imag} */,
  {32'h43e1c174, 32'h00000000} /* (26, 19, 30) {real, imag} */,
  {32'hc44280fc, 32'h00000000} /* (26, 19, 29) {real, imag} */,
  {32'hc252a51c, 32'h00000000} /* (26, 19, 28) {real, imag} */,
  {32'hc419c568, 32'h00000000} /* (26, 19, 27) {real, imag} */,
  {32'hc350c5b6, 32'h00000000} /* (26, 19, 26) {real, imag} */,
  {32'hc3d3de23, 32'h00000000} /* (26, 19, 25) {real, imag} */,
  {32'hc4024992, 32'h00000000} /* (26, 19, 24) {real, imag} */,
  {32'h42ca5d18, 32'h00000000} /* (26, 19, 23) {real, imag} */,
  {32'hc3bb8f1e, 32'h00000000} /* (26, 19, 22) {real, imag} */,
  {32'hc3511d76, 32'h00000000} /* (26, 19, 21) {real, imag} */,
  {32'hc34d1ed0, 32'h00000000} /* (26, 19, 20) {real, imag} */,
  {32'h4393f872, 32'h00000000} /* (26, 19, 19) {real, imag} */,
  {32'hc3088d44, 32'h00000000} /* (26, 19, 18) {real, imag} */,
  {32'hc3d20822, 32'h00000000} /* (26, 19, 17) {real, imag} */,
  {32'h44f95c82, 32'h00000000} /* (26, 19, 16) {real, imag} */,
  {32'h449f51dd, 32'h00000000} /* (26, 19, 15) {real, imag} */,
  {32'h441a7342, 32'h00000000} /* (26, 19, 14) {real, imag} */,
  {32'h44125be4, 32'h00000000} /* (26, 19, 13) {real, imag} */,
  {32'h43970d40, 32'h00000000} /* (26, 19, 12) {real, imag} */,
  {32'h443abe28, 32'h00000000} /* (26, 19, 11) {real, imag} */,
  {32'h4275a098, 32'h00000000} /* (26, 19, 10) {real, imag} */,
  {32'h4282fc0c, 32'h00000000} /* (26, 19, 9) {real, imag} */,
  {32'h43ef2024, 32'h00000000} /* (26, 19, 8) {real, imag} */,
  {32'hc387b5da, 32'h00000000} /* (26, 19, 7) {real, imag} */,
  {32'hc39b1624, 32'h00000000} /* (26, 19, 6) {real, imag} */,
  {32'hc473c416, 32'h00000000} /* (26, 19, 5) {real, imag} */,
  {32'hc4e23199, 32'h00000000} /* (26, 19, 4) {real, imag} */,
  {32'hc46f0c9f, 32'h00000000} /* (26, 19, 3) {real, imag} */,
  {32'hc4070027, 32'h00000000} /* (26, 19, 2) {real, imag} */,
  {32'hc2984ad8, 32'h00000000} /* (26, 19, 1) {real, imag} */,
  {32'hc18c9380, 32'h00000000} /* (26, 19, 0) {real, imag} */,
  {32'h44974634, 32'h00000000} /* (26, 18, 31) {real, imag} */,
  {32'h43cd448c, 32'h00000000} /* (26, 18, 30) {real, imag} */,
  {32'h434dedee, 32'h00000000} /* (26, 18, 29) {real, imag} */,
  {32'h428d9fe8, 32'h00000000} /* (26, 18, 28) {real, imag} */,
  {32'hc3d51288, 32'h00000000} /* (26, 18, 27) {real, imag} */,
  {32'h4285b3ac, 32'h00000000} /* (26, 18, 26) {real, imag} */,
  {32'hc32c9b10, 32'h00000000} /* (26, 18, 25) {real, imag} */,
  {32'hc4357c74, 32'h00000000} /* (26, 18, 24) {real, imag} */,
  {32'hc4ae167a, 32'h00000000} /* (26, 18, 23) {real, imag} */,
  {32'hc45c09a8, 32'h00000000} /* (26, 18, 22) {real, imag} */,
  {32'hc3b28f2c, 32'h00000000} /* (26, 18, 21) {real, imag} */,
  {32'hc3c9cc34, 32'h00000000} /* (26, 18, 20) {real, imag} */,
  {32'h42b15750, 32'h00000000} /* (26, 18, 19) {real, imag} */,
  {32'hc3d7ec95, 32'h00000000} /* (26, 18, 18) {real, imag} */,
  {32'h43fe6fbe, 32'h00000000} /* (26, 18, 17) {real, imag} */,
  {32'h442a4e76, 32'h00000000} /* (26, 18, 16) {real, imag} */,
  {32'h4483d834, 32'h00000000} /* (26, 18, 15) {real, imag} */,
  {32'h4414904a, 32'h00000000} /* (26, 18, 14) {real, imag} */,
  {32'hc3c6d52f, 32'h00000000} /* (26, 18, 13) {real, imag} */,
  {32'hc3ba6d5c, 32'h00000000} /* (26, 18, 12) {real, imag} */,
  {32'h44803bce, 32'h00000000} /* (26, 18, 11) {real, imag} */,
  {32'h445ca6ec, 32'h00000000} /* (26, 18, 10) {real, imag} */,
  {32'h42eb1ab0, 32'h00000000} /* (26, 18, 9) {real, imag} */,
  {32'h4375f71a, 32'h00000000} /* (26, 18, 8) {real, imag} */,
  {32'h4341be28, 32'h00000000} /* (26, 18, 7) {real, imag} */,
  {32'h40ed3300, 32'h00000000} /* (26, 18, 6) {real, imag} */,
  {32'h41aefe80, 32'h00000000} /* (26, 18, 5) {real, imag} */,
  {32'hc433aeb2, 32'h00000000} /* (26, 18, 4) {real, imag} */,
  {32'hc46a73d6, 32'h00000000} /* (26, 18, 3) {real, imag} */,
  {32'h43848c53, 32'h00000000} /* (26, 18, 2) {real, imag} */,
  {32'h44162949, 32'h00000000} /* (26, 18, 1) {real, imag} */,
  {32'h43069762, 32'h00000000} /* (26, 18, 0) {real, imag} */,
  {32'h442fff6e, 32'h00000000} /* (26, 17, 31) {real, imag} */,
  {32'h416eba00, 32'h00000000} /* (26, 17, 30) {real, imag} */,
  {32'h441acc78, 32'h00000000} /* (26, 17, 29) {real, imag} */,
  {32'hc3110ba7, 32'h00000000} /* (26, 17, 28) {real, imag} */,
  {32'hc329932f, 32'h00000000} /* (26, 17, 27) {real, imag} */,
  {32'h4475a0c8, 32'h00000000} /* (26, 17, 26) {real, imag} */,
  {32'hc4153bf2, 32'h00000000} /* (26, 17, 25) {real, imag} */,
  {32'hc4148bc6, 32'h00000000} /* (26, 17, 24) {real, imag} */,
  {32'hc454b3c9, 32'h00000000} /* (26, 17, 23) {real, imag} */,
  {32'hc40980bc, 32'h00000000} /* (26, 17, 22) {real, imag} */,
  {32'hc475c4f2, 32'h00000000} /* (26, 17, 21) {real, imag} */,
  {32'hc4613616, 32'h00000000} /* (26, 17, 20) {real, imag} */,
  {32'hc3bb0c22, 32'h00000000} /* (26, 17, 19) {real, imag} */,
  {32'h4322cd7a, 32'h00000000} /* (26, 17, 18) {real, imag} */,
  {32'h44317781, 32'h00000000} /* (26, 17, 17) {real, imag} */,
  {32'h43c3c5da, 32'h00000000} /* (26, 17, 16) {real, imag} */,
  {32'h440095aa, 32'h00000000} /* (26, 17, 15) {real, imag} */,
  {32'h4422c952, 32'h00000000} /* (26, 17, 14) {real, imag} */,
  {32'hc4232e82, 32'h00000000} /* (26, 17, 13) {real, imag} */,
  {32'hc395370c, 32'h00000000} /* (26, 17, 12) {real, imag} */,
  {32'h436c9e37, 32'h00000000} /* (26, 17, 11) {real, imag} */,
  {32'h43deeeb0, 32'h00000000} /* (26, 17, 10) {real, imag} */,
  {32'h44469456, 32'h00000000} /* (26, 17, 9) {real, imag} */,
  {32'h43b1e717, 32'h00000000} /* (26, 17, 8) {real, imag} */,
  {32'h448ead44, 32'h00000000} /* (26, 17, 7) {real, imag} */,
  {32'h448d8868, 32'h00000000} /* (26, 17, 6) {real, imag} */,
  {32'hc3685fa8, 32'h00000000} /* (26, 17, 5) {real, imag} */,
  {32'h438b686c, 32'h00000000} /* (26, 17, 4) {real, imag} */,
  {32'hc363f62c, 32'h00000000} /* (26, 17, 3) {real, imag} */,
  {32'hc4078f74, 32'h00000000} /* (26, 17, 2) {real, imag} */,
  {32'h43beefbe, 32'h00000000} /* (26, 17, 1) {real, imag} */,
  {32'h439d656a, 32'h00000000} /* (26, 17, 0) {real, imag} */,
  {32'h42eae377, 32'h00000000} /* (26, 16, 31) {real, imag} */,
  {32'h441876ba, 32'h00000000} /* (26, 16, 30) {real, imag} */,
  {32'h44342f85, 32'h00000000} /* (26, 16, 29) {real, imag} */,
  {32'h442ffefc, 32'h00000000} /* (26, 16, 28) {real, imag} */,
  {32'hc36ec18f, 32'h00000000} /* (26, 16, 27) {real, imag} */,
  {32'hc220f4b8, 32'h00000000} /* (26, 16, 26) {real, imag} */,
  {32'hc3d2e36d, 32'h00000000} /* (26, 16, 25) {real, imag} */,
  {32'hc32d50be, 32'h00000000} /* (26, 16, 24) {real, imag} */,
  {32'hc20d1970, 32'h00000000} /* (26, 16, 23) {real, imag} */,
  {32'hc4844d5e, 32'h00000000} /* (26, 16, 22) {real, imag} */,
  {32'hc40f8680, 32'h00000000} /* (26, 16, 21) {real, imag} */,
  {32'hc3e879dc, 32'h00000000} /* (26, 16, 20) {real, imag} */,
  {32'hc341e99e, 32'h00000000} /* (26, 16, 19) {real, imag} */,
  {32'h439d79e8, 32'h00000000} /* (26, 16, 18) {real, imag} */,
  {32'hc3c0a79c, 32'h00000000} /* (26, 16, 17) {real, imag} */,
  {32'hc1689ae0, 32'h00000000} /* (26, 16, 16) {real, imag} */,
  {32'h41a73424, 32'h00000000} /* (26, 16, 15) {real, imag} */,
  {32'hc2f0dc64, 32'h00000000} /* (26, 16, 14) {real, imag} */,
  {32'hc3fd96c2, 32'h00000000} /* (26, 16, 13) {real, imag} */,
  {32'h448156a5, 32'h00000000} /* (26, 16, 12) {real, imag} */,
  {32'hc3662fb5, 32'h00000000} /* (26, 16, 11) {real, imag} */,
  {32'h4444e2b4, 32'h00000000} /* (26, 16, 10) {real, imag} */,
  {32'h442aa272, 32'h00000000} /* (26, 16, 9) {real, imag} */,
  {32'h431126da, 32'h00000000} /* (26, 16, 8) {real, imag} */,
  {32'h44964938, 32'h00000000} /* (26, 16, 7) {real, imag} */,
  {32'h44ae3d7a, 32'h00000000} /* (26, 16, 6) {real, imag} */,
  {32'h440b0d48, 32'h00000000} /* (26, 16, 5) {real, imag} */,
  {32'h43921358, 32'h00000000} /* (26, 16, 4) {real, imag} */,
  {32'h430c9b86, 32'h00000000} /* (26, 16, 3) {real, imag} */,
  {32'hc3216a60, 32'h00000000} /* (26, 16, 2) {real, imag} */,
  {32'h43d146ec, 32'h00000000} /* (26, 16, 1) {real, imag} */,
  {32'h4481a9bc, 32'h00000000} /* (26, 16, 0) {real, imag} */,
  {32'h4390bb44, 32'h00000000} /* (26, 15, 31) {real, imag} */,
  {32'hc3d506dc, 32'h00000000} /* (26, 15, 30) {real, imag} */,
  {32'hc48096ee, 32'h00000000} /* (26, 15, 29) {real, imag} */,
  {32'h4468fc9c, 32'h00000000} /* (26, 15, 28) {real, imag} */,
  {32'hc353d298, 32'h00000000} /* (26, 15, 27) {real, imag} */,
  {32'hc34c6b53, 32'h00000000} /* (26, 15, 26) {real, imag} */,
  {32'hc48a9bf0, 32'h00000000} /* (26, 15, 25) {real, imag} */,
  {32'h43f96b88, 32'h00000000} /* (26, 15, 24) {real, imag} */,
  {32'h4324f212, 32'h00000000} /* (26, 15, 23) {real, imag} */,
  {32'hc4dc7cd7, 32'h00000000} /* (26, 15, 22) {real, imag} */,
  {32'hc4331a53, 32'h00000000} /* (26, 15, 21) {real, imag} */,
  {32'hc42f3074, 32'h00000000} /* (26, 15, 20) {real, imag} */,
  {32'hc4924e1a, 32'h00000000} /* (26, 15, 19) {real, imag} */,
  {32'hc497c4e6, 32'h00000000} /* (26, 15, 18) {real, imag} */,
  {32'hc4f41786, 32'h00000000} /* (26, 15, 17) {real, imag} */,
  {32'hc2ec247a, 32'h00000000} /* (26, 15, 16) {real, imag} */,
  {32'hc3c76798, 32'h00000000} /* (26, 15, 15) {real, imag} */,
  {32'hc42f5696, 32'h00000000} /* (26, 15, 14) {real, imag} */,
  {32'hc31b3722, 32'h00000000} /* (26, 15, 13) {real, imag} */,
  {32'h434b5d92, 32'h00000000} /* (26, 15, 12) {real, imag} */,
  {32'h432aed78, 32'h00000000} /* (26, 15, 11) {real, imag} */,
  {32'hc3ca1eba, 32'h00000000} /* (26, 15, 10) {real, imag} */,
  {32'hc2bd1748, 32'h00000000} /* (26, 15, 9) {real, imag} */,
  {32'hc3a97488, 32'h00000000} /* (26, 15, 8) {real, imag} */,
  {32'hc36e18ae, 32'h00000000} /* (26, 15, 7) {real, imag} */,
  {32'h4439b3be, 32'h00000000} /* (26, 15, 6) {real, imag} */,
  {32'h430aeb1c, 32'h00000000} /* (26, 15, 5) {real, imag} */,
  {32'h42f8470c, 32'h00000000} /* (26, 15, 4) {real, imag} */,
  {32'hc3c924f8, 32'h00000000} /* (26, 15, 3) {real, imag} */,
  {32'hc39241de, 32'h00000000} /* (26, 15, 2) {real, imag} */,
  {32'h440a40cd, 32'h00000000} /* (26, 15, 1) {real, imag} */,
  {32'h43c1aa10, 32'h00000000} /* (26, 15, 0) {real, imag} */,
  {32'h435ee43a, 32'h00000000} /* (26, 14, 31) {real, imag} */,
  {32'hc3fdcb85, 32'h00000000} /* (26, 14, 30) {real, imag} */,
  {32'hc4269aec, 32'h00000000} /* (26, 14, 29) {real, imag} */,
  {32'hc39821e9, 32'h00000000} /* (26, 14, 28) {real, imag} */,
  {32'hc414c376, 32'h00000000} /* (26, 14, 27) {real, imag} */,
  {32'hc3717dfc, 32'h00000000} /* (26, 14, 26) {real, imag} */,
  {32'hc4bf6d7f, 32'h00000000} /* (26, 14, 25) {real, imag} */,
  {32'hc3d433cd, 32'h00000000} /* (26, 14, 24) {real, imag} */,
  {32'hc452b288, 32'h00000000} /* (26, 14, 23) {real, imag} */,
  {32'hc4aebef4, 32'h00000000} /* (26, 14, 22) {real, imag} */,
  {32'hc484bbea, 32'h00000000} /* (26, 14, 21) {real, imag} */,
  {32'hc413ab55, 32'h00000000} /* (26, 14, 20) {real, imag} */,
  {32'hc36b41aa, 32'h00000000} /* (26, 14, 19) {real, imag} */,
  {32'hc435f516, 32'h00000000} /* (26, 14, 18) {real, imag} */,
  {32'hc44dd6f0, 32'h00000000} /* (26, 14, 17) {real, imag} */,
  {32'hc42ba794, 32'h00000000} /* (26, 14, 16) {real, imag} */,
  {32'hc3e1db4b, 32'h00000000} /* (26, 14, 15) {real, imag} */,
  {32'hc3dc0351, 32'h00000000} /* (26, 14, 14) {real, imag} */,
  {32'hc41ad552, 32'h00000000} /* (26, 14, 13) {real, imag} */,
  {32'hc3a7a577, 32'h00000000} /* (26, 14, 12) {real, imag} */,
  {32'hc2b5920c, 32'h00000000} /* (26, 14, 11) {real, imag} */,
  {32'hc3b0234a, 32'h00000000} /* (26, 14, 10) {real, imag} */,
  {32'hc3db12f4, 32'h00000000} /* (26, 14, 9) {real, imag} */,
  {32'h4205b678, 32'h00000000} /* (26, 14, 8) {real, imag} */,
  {32'h43cbf285, 32'h00000000} /* (26, 14, 7) {real, imag} */,
  {32'h439a83ac, 32'h00000000} /* (26, 14, 6) {real, imag} */,
  {32'hc28f0ee8, 32'h00000000} /* (26, 14, 5) {real, imag} */,
  {32'h445102d9, 32'h00000000} /* (26, 14, 4) {real, imag} */,
  {32'h446fc4b6, 32'h00000000} /* (26, 14, 3) {real, imag} */,
  {32'hc3d8219d, 32'h00000000} /* (26, 14, 2) {real, imag} */,
  {32'h43ce0d1d, 32'h00000000} /* (26, 14, 1) {real, imag} */,
  {32'h43abfda8, 32'h00000000} /* (26, 14, 0) {real, imag} */,
  {32'h43612380, 32'h00000000} /* (26, 13, 31) {real, imag} */,
  {32'hc3993422, 32'h00000000} /* (26, 13, 30) {real, imag} */,
  {32'hc40ae776, 32'h00000000} /* (26, 13, 29) {real, imag} */,
  {32'hc38cc8c8, 32'h00000000} /* (26, 13, 28) {real, imag} */,
  {32'h442c6373, 32'h00000000} /* (26, 13, 27) {real, imag} */,
  {32'hc3c4dd2c, 32'h00000000} /* (26, 13, 26) {real, imag} */,
  {32'hc427055b, 32'h00000000} /* (26, 13, 25) {real, imag} */,
  {32'hc48a5f92, 32'h00000000} /* (26, 13, 24) {real, imag} */,
  {32'hc3d5029a, 32'h00000000} /* (26, 13, 23) {real, imag} */,
  {32'hc49aab32, 32'h00000000} /* (26, 13, 22) {real, imag} */,
  {32'hc4a29b57, 32'h00000000} /* (26, 13, 21) {real, imag} */,
  {32'hc39859f0, 32'h00000000} /* (26, 13, 20) {real, imag} */,
  {32'hc41772be, 32'h00000000} /* (26, 13, 19) {real, imag} */,
  {32'h434a4ee8, 32'h00000000} /* (26, 13, 18) {real, imag} */,
  {32'hc42aab1c, 32'h00000000} /* (26, 13, 17) {real, imag} */,
  {32'hc493a830, 32'h00000000} /* (26, 13, 16) {real, imag} */,
  {32'hc49ccac2, 32'h00000000} /* (26, 13, 15) {real, imag} */,
  {32'hc492f1dc, 32'h00000000} /* (26, 13, 14) {real, imag} */,
  {32'hc4138c1e, 32'h00000000} /* (26, 13, 13) {real, imag} */,
  {32'hc2b5b0b1, 32'h00000000} /* (26, 13, 12) {real, imag} */,
  {32'h4305ddbc, 32'h00000000} /* (26, 13, 11) {real, imag} */,
  {32'h4317a948, 32'h00000000} /* (26, 13, 10) {real, imag} */,
  {32'h43bcec9a, 32'h00000000} /* (26, 13, 9) {real, imag} */,
  {32'h42fceb98, 32'h00000000} /* (26, 13, 8) {real, imag} */,
  {32'hc3d5831c, 32'h00000000} /* (26, 13, 7) {real, imag} */,
  {32'h429f7b58, 32'h00000000} /* (26, 13, 6) {real, imag} */,
  {32'h4438a87e, 32'h00000000} /* (26, 13, 5) {real, imag} */,
  {32'h4482085d, 32'h00000000} /* (26, 13, 4) {real, imag} */,
  {32'h4409f832, 32'h00000000} /* (26, 13, 3) {real, imag} */,
  {32'hc387d0c7, 32'h00000000} /* (26, 13, 2) {real, imag} */,
  {32'hc3408d49, 32'h00000000} /* (26, 13, 1) {real, imag} */,
  {32'h438de504, 32'h00000000} /* (26, 13, 0) {real, imag} */,
  {32'hc29da7f8, 32'h00000000} /* (26, 12, 31) {real, imag} */,
  {32'h42376480, 32'h00000000} /* (26, 12, 30) {real, imag} */,
  {32'h4231798a, 32'h00000000} /* (26, 12, 29) {real, imag} */,
  {32'h434bb10a, 32'h00000000} /* (26, 12, 28) {real, imag} */,
  {32'hc395d066, 32'h00000000} /* (26, 12, 27) {real, imag} */,
  {32'hc24d9354, 32'h00000000} /* (26, 12, 26) {real, imag} */,
  {32'hc457bd90, 32'h00000000} /* (26, 12, 25) {real, imag} */,
  {32'hc39f2d5c, 32'h00000000} /* (26, 12, 24) {real, imag} */,
  {32'hc23289f6, 32'h00000000} /* (26, 12, 23) {real, imag} */,
  {32'hc3abc3bd, 32'h00000000} /* (26, 12, 22) {real, imag} */,
  {32'hc3ac12a6, 32'h00000000} /* (26, 12, 21) {real, imag} */,
  {32'hc4362c33, 32'h00000000} /* (26, 12, 20) {real, imag} */,
  {32'hc45edcfe, 32'h00000000} /* (26, 12, 19) {real, imag} */,
  {32'hc3961758, 32'h00000000} /* (26, 12, 18) {real, imag} */,
  {32'hc3d65e7a, 32'h00000000} /* (26, 12, 17) {real, imag} */,
  {32'hc42c0f46, 32'h00000000} /* (26, 12, 16) {real, imag} */,
  {32'hc3fb381e, 32'h00000000} /* (26, 12, 15) {real, imag} */,
  {32'hc4232268, 32'h00000000} /* (26, 12, 14) {real, imag} */,
  {32'hc3036bac, 32'h00000000} /* (26, 12, 13) {real, imag} */,
  {32'hc3eff9e1, 32'h00000000} /* (26, 12, 12) {real, imag} */,
  {32'h4350c1a7, 32'h00000000} /* (26, 12, 11) {real, imag} */,
  {32'h4331e3fc, 32'h00000000} /* (26, 12, 10) {real, imag} */,
  {32'h43bd8fe1, 32'h00000000} /* (26, 12, 9) {real, imag} */,
  {32'hc3ecf0ec, 32'h00000000} /* (26, 12, 8) {real, imag} */,
  {32'hc2871cc1, 32'h00000000} /* (26, 12, 7) {real, imag} */,
  {32'h432c5742, 32'h00000000} /* (26, 12, 6) {real, imag} */,
  {32'h421b8a34, 32'h00000000} /* (26, 12, 5) {real, imag} */,
  {32'h4344c2b4, 32'h00000000} /* (26, 12, 4) {real, imag} */,
  {32'hc419815a, 32'h00000000} /* (26, 12, 3) {real, imag} */,
  {32'hc3a222be, 32'h00000000} /* (26, 12, 2) {real, imag} */,
  {32'hc4813a06, 32'h00000000} /* (26, 12, 1) {real, imag} */,
  {32'h440ab1fe, 32'h00000000} /* (26, 12, 0) {real, imag} */,
  {32'h43c271e9, 32'h00000000} /* (26, 11, 31) {real, imag} */,
  {32'h43aa2a80, 32'h00000000} /* (26, 11, 30) {real, imag} */,
  {32'hc40cf7c4, 32'h00000000} /* (26, 11, 29) {real, imag} */,
  {32'hc46be500, 32'h00000000} /* (26, 11, 28) {real, imag} */,
  {32'hc365c5ca, 32'h00000000} /* (26, 11, 27) {real, imag} */,
  {32'hc4690ee0, 32'h00000000} /* (26, 11, 26) {real, imag} */,
  {32'hc4140f77, 32'h00000000} /* (26, 11, 25) {real, imag} */,
  {32'h43a4ecf6, 32'h00000000} /* (26, 11, 24) {real, imag} */,
  {32'h426f1940, 32'h00000000} /* (26, 11, 23) {real, imag} */,
  {32'h43cdc2f0, 32'h00000000} /* (26, 11, 22) {real, imag} */,
  {32'h43bea196, 32'h00000000} /* (26, 11, 21) {real, imag} */,
  {32'h42e25f2e, 32'h00000000} /* (26, 11, 20) {real, imag} */,
  {32'hc48069ca, 32'h00000000} /* (26, 11, 19) {real, imag} */,
  {32'hc3f79590, 32'h00000000} /* (26, 11, 18) {real, imag} */,
  {32'h43a88622, 32'h00000000} /* (26, 11, 17) {real, imag} */,
  {32'hc3941ae5, 32'h00000000} /* (26, 11, 16) {real, imag} */,
  {32'h4311338a, 32'h00000000} /* (26, 11, 15) {real, imag} */,
  {32'hc405575f, 32'h00000000} /* (26, 11, 14) {real, imag} */,
  {32'hc45097e8, 32'h00000000} /* (26, 11, 13) {real, imag} */,
  {32'hc1ae9410, 32'h00000000} /* (26, 11, 12) {real, imag} */,
  {32'hc289d304, 32'h00000000} /* (26, 11, 11) {real, imag} */,
  {32'h441481ac, 32'h00000000} /* (26, 11, 10) {real, imag} */,
  {32'h443091f1, 32'h00000000} /* (26, 11, 9) {real, imag} */,
  {32'h448c19d6, 32'h00000000} /* (26, 11, 8) {real, imag} */,
  {32'h44ac7566, 32'h00000000} /* (26, 11, 7) {real, imag} */,
  {32'h439322f8, 32'h00000000} /* (26, 11, 6) {real, imag} */,
  {32'hc248d41c, 32'h00000000} /* (26, 11, 5) {real, imag} */,
  {32'h4418e8e2, 32'h00000000} /* (26, 11, 4) {real, imag} */,
  {32'hc458f968, 32'h00000000} /* (26, 11, 3) {real, imag} */,
  {32'hc4086088, 32'h00000000} /* (26, 11, 2) {real, imag} */,
  {32'hc402f19a, 32'h00000000} /* (26, 11, 1) {real, imag} */,
  {32'hc3aac9f3, 32'h00000000} /* (26, 11, 0) {real, imag} */,
  {32'hc41db0b6, 32'h00000000} /* (26, 10, 31) {real, imag} */,
  {32'h438d4656, 32'h00000000} /* (26, 10, 30) {real, imag} */,
  {32'hc492f074, 32'h00000000} /* (26, 10, 29) {real, imag} */,
  {32'hc4984444, 32'h00000000} /* (26, 10, 28) {real, imag} */,
  {32'hc3fe3712, 32'h00000000} /* (26, 10, 27) {real, imag} */,
  {32'hc4479c5e, 32'h00000000} /* (26, 10, 26) {real, imag} */,
  {32'hc4366b36, 32'h00000000} /* (26, 10, 25) {real, imag} */,
  {32'hc3ede142, 32'h00000000} /* (26, 10, 24) {real, imag} */,
  {32'h434543a8, 32'h00000000} /* (26, 10, 23) {real, imag} */,
  {32'hc40319c1, 32'h00000000} /* (26, 10, 22) {real, imag} */,
  {32'hc4906e21, 32'h00000000} /* (26, 10, 21) {real, imag} */,
  {32'h43b1c0e6, 32'h00000000} /* (26, 10, 20) {real, imag} */,
  {32'hc4649b6f, 32'h00000000} /* (26, 10, 19) {real, imag} */,
  {32'hc48e349c, 32'h00000000} /* (26, 10, 18) {real, imag} */,
  {32'hc4a139ae, 32'h00000000} /* (26, 10, 17) {real, imag} */,
  {32'h43990222, 32'h00000000} /* (26, 10, 16) {real, imag} */,
  {32'hc33b885e, 32'h00000000} /* (26, 10, 15) {real, imag} */,
  {32'hc4998664, 32'h00000000} /* (26, 10, 14) {real, imag} */,
  {32'hc38cca9a, 32'h00000000} /* (26, 10, 13) {real, imag} */,
  {32'hc3adb916, 32'h00000000} /* (26, 10, 12) {real, imag} */,
  {32'hc3e98ae2, 32'h00000000} /* (26, 10, 11) {real, imag} */,
  {32'h435ea644, 32'h00000000} /* (26, 10, 10) {real, imag} */,
  {32'h444a4146, 32'h00000000} /* (26, 10, 9) {real, imag} */,
  {32'h4452e9f7, 32'h00000000} /* (26, 10, 8) {real, imag} */,
  {32'h44959759, 32'h00000000} /* (26, 10, 7) {real, imag} */,
  {32'h448f7b04, 32'h00000000} /* (26, 10, 6) {real, imag} */,
  {32'h43bee8f9, 32'h00000000} /* (26, 10, 5) {real, imag} */,
  {32'h4404eb39, 32'h00000000} /* (26, 10, 4) {real, imag} */,
  {32'hc41eef67, 32'h00000000} /* (26, 10, 3) {real, imag} */,
  {32'hc44ede18, 32'h00000000} /* (26, 10, 2) {real, imag} */,
  {32'h43d6065a, 32'h00000000} /* (26, 10, 1) {real, imag} */,
  {32'h43da8ffe, 32'h00000000} /* (26, 10, 0) {real, imag} */,
  {32'hc42017fd, 32'h00000000} /* (26, 9, 31) {real, imag} */,
  {32'hc3fa2ce8, 32'h00000000} /* (26, 9, 30) {real, imag} */,
  {32'hc4755b86, 32'h00000000} /* (26, 9, 29) {real, imag} */,
  {32'hc4b9d6ff, 32'h00000000} /* (26, 9, 28) {real, imag} */,
  {32'hc4dbd1d4, 32'h00000000} /* (26, 9, 27) {real, imag} */,
  {32'hc44e0257, 32'h00000000} /* (26, 9, 26) {real, imag} */,
  {32'hc4b1e400, 32'h00000000} /* (26, 9, 25) {real, imag} */,
  {32'hc2f27f18, 32'h00000000} /* (26, 9, 24) {real, imag} */,
  {32'hc4847114, 32'h00000000} /* (26, 9, 23) {real, imag} */,
  {32'hc46988e4, 32'h00000000} /* (26, 9, 22) {real, imag} */,
  {32'hc3ba2ff4, 32'h00000000} /* (26, 9, 21) {real, imag} */,
  {32'hc3e8aa70, 32'h00000000} /* (26, 9, 20) {real, imag} */,
  {32'hc47ac8e9, 32'h00000000} /* (26, 9, 19) {real, imag} */,
  {32'hc4a74fd9, 32'h00000000} /* (26, 9, 18) {real, imag} */,
  {32'hc4642317, 32'h00000000} /* (26, 9, 17) {real, imag} */,
  {32'hc41deea4, 32'h00000000} /* (26, 9, 16) {real, imag} */,
  {32'hc47da7b1, 32'h00000000} /* (26, 9, 15) {real, imag} */,
  {32'hc3ee7b08, 32'h00000000} /* (26, 9, 14) {real, imag} */,
  {32'hc48b5c8d, 32'h00000000} /* (26, 9, 13) {real, imag} */,
  {32'hc43fda0e, 32'h00000000} /* (26, 9, 12) {real, imag} */,
  {32'h4325f7bc, 32'h00000000} /* (26, 9, 11) {real, imag} */,
  {32'h435fc75c, 32'h00000000} /* (26, 9, 10) {real, imag} */,
  {32'h4400e728, 32'h00000000} /* (26, 9, 9) {real, imag} */,
  {32'h4484fd5c, 32'h00000000} /* (26, 9, 8) {real, imag} */,
  {32'h44456ef8, 32'h00000000} /* (26, 9, 7) {real, imag} */,
  {32'h44769aae, 32'h00000000} /* (26, 9, 6) {real, imag} */,
  {32'hc213be40, 32'h00000000} /* (26, 9, 5) {real, imag} */,
  {32'h43020900, 32'h00000000} /* (26, 9, 4) {real, imag} */,
  {32'hc4261c75, 32'h00000000} /* (26, 9, 3) {real, imag} */,
  {32'hc40c14ca, 32'h00000000} /* (26, 9, 2) {real, imag} */,
  {32'hc38df4b2, 32'h00000000} /* (26, 9, 1) {real, imag} */,
  {32'hc47edcba, 32'h00000000} /* (26, 9, 0) {real, imag} */,
  {32'hc48bd49a, 32'h00000000} /* (26, 8, 31) {real, imag} */,
  {32'hc4b70161, 32'h00000000} /* (26, 8, 30) {real, imag} */,
  {32'hc51bdde2, 32'h00000000} /* (26, 8, 29) {real, imag} */,
  {32'hc50190e0, 32'h00000000} /* (26, 8, 28) {real, imag} */,
  {32'hc4f753f6, 32'h00000000} /* (26, 8, 27) {real, imag} */,
  {32'hc50fce7e, 32'h00000000} /* (26, 8, 26) {real, imag} */,
  {32'hc500e4a5, 32'h00000000} /* (26, 8, 25) {real, imag} */,
  {32'hc4ce80a6, 32'h00000000} /* (26, 8, 24) {real, imag} */,
  {32'hc48ffc7f, 32'h00000000} /* (26, 8, 23) {real, imag} */,
  {32'hc47f2123, 32'h00000000} /* (26, 8, 22) {real, imag} */,
  {32'hc48b1f0c, 32'h00000000} /* (26, 8, 21) {real, imag} */,
  {32'hc4851715, 32'h00000000} /* (26, 8, 20) {real, imag} */,
  {32'hc48e006a, 32'h00000000} /* (26, 8, 19) {real, imag} */,
  {32'hc4c384ca, 32'h00000000} /* (26, 8, 18) {real, imag} */,
  {32'hc496a14a, 32'h00000000} /* (26, 8, 17) {real, imag} */,
  {32'hc489917e, 32'h00000000} /* (26, 8, 16) {real, imag} */,
  {32'hc48e90b6, 32'h00000000} /* (26, 8, 15) {real, imag} */,
  {32'hc48fc5af, 32'h00000000} /* (26, 8, 14) {real, imag} */,
  {32'hc44ca95e, 32'h00000000} /* (26, 8, 13) {real, imag} */,
  {32'hc4438362, 32'h00000000} /* (26, 8, 12) {real, imag} */,
  {32'hc400ef80, 32'h00000000} /* (26, 8, 11) {real, imag} */,
  {32'h4379d438, 32'h00000000} /* (26, 8, 10) {real, imag} */,
  {32'h448f7962, 32'h00000000} /* (26, 8, 9) {real, imag} */,
  {32'h444f2e39, 32'h00000000} /* (26, 8, 8) {real, imag} */,
  {32'h444ad0cc, 32'h00000000} /* (26, 8, 7) {real, imag} */,
  {32'h442941a9, 32'h00000000} /* (26, 8, 6) {real, imag} */,
  {32'hc38a56fb, 32'h00000000} /* (26, 8, 5) {real, imag} */,
  {32'h4294571c, 32'h00000000} /* (26, 8, 4) {real, imag} */,
  {32'hc450c460, 32'h00000000} /* (26, 8, 3) {real, imag} */,
  {32'hc45fdc1c, 32'h00000000} /* (26, 8, 2) {real, imag} */,
  {32'hc481b87e, 32'h00000000} /* (26, 8, 1) {real, imag} */,
  {32'hc5092c51, 32'h00000000} /* (26, 8, 0) {real, imag} */,
  {32'hc51e171f, 32'h00000000} /* (26, 7, 31) {real, imag} */,
  {32'hc4ff2f72, 32'h00000000} /* (26, 7, 30) {real, imag} */,
  {32'hc5614b20, 32'h00000000} /* (26, 7, 29) {real, imag} */,
  {32'hc577e8ab, 32'h00000000} /* (26, 7, 28) {real, imag} */,
  {32'hc52c6289, 32'h00000000} /* (26, 7, 27) {real, imag} */,
  {32'hc4ff6ae3, 32'h00000000} /* (26, 7, 26) {real, imag} */,
  {32'hc51b8970, 32'h00000000} /* (26, 7, 25) {real, imag} */,
  {32'hc4e565bb, 32'h00000000} /* (26, 7, 24) {real, imag} */,
  {32'hc42f990d, 32'h00000000} /* (26, 7, 23) {real, imag} */,
  {32'hc446d8c6, 32'h00000000} /* (26, 7, 22) {real, imag} */,
  {32'hc4a66ebc, 32'h00000000} /* (26, 7, 21) {real, imag} */,
  {32'hc4792c9d, 32'h00000000} /* (26, 7, 20) {real, imag} */,
  {32'hc43f673a, 32'h00000000} /* (26, 7, 19) {real, imag} */,
  {32'hc4aad51b, 32'h00000000} /* (26, 7, 18) {real, imag} */,
  {32'hc4b59f1e, 32'h00000000} /* (26, 7, 17) {real, imag} */,
  {32'hc4a936ca, 32'h00000000} /* (26, 7, 16) {real, imag} */,
  {32'hc4043d8b, 32'h00000000} /* (26, 7, 15) {real, imag} */,
  {32'hc33818a0, 32'h00000000} /* (26, 7, 14) {real, imag} */,
  {32'hc3c42964, 32'h00000000} /* (26, 7, 13) {real, imag} */,
  {32'hc30cc610, 32'h00000000} /* (26, 7, 12) {real, imag} */,
  {32'hc46801a0, 32'h00000000} /* (26, 7, 11) {real, imag} */,
  {32'h43b89c14, 32'h00000000} /* (26, 7, 10) {real, imag} */,
  {32'h445d6d56, 32'h00000000} /* (26, 7, 9) {real, imag} */,
  {32'h42795760, 32'h00000000} /* (26, 7, 8) {real, imag} */,
  {32'h438ff81a, 32'h00000000} /* (26, 7, 7) {real, imag} */,
  {32'h437939be, 32'h00000000} /* (26, 7, 6) {real, imag} */,
  {32'hc3ef6c5a, 32'h00000000} /* (26, 7, 5) {real, imag} */,
  {32'hc15036c0, 32'h00000000} /* (26, 7, 4) {real, imag} */,
  {32'hc44f2ada, 32'h00000000} /* (26, 7, 3) {real, imag} */,
  {32'hc4e76b5f, 32'h00000000} /* (26, 7, 2) {real, imag} */,
  {32'hc4c72c90, 32'h00000000} /* (26, 7, 1) {real, imag} */,
  {32'hc4d168b2, 32'h00000000} /* (26, 7, 0) {real, imag} */,
  {32'hc51e63dc, 32'h00000000} /* (26, 6, 31) {real, imag} */,
  {32'hc5579f48, 32'h00000000} /* (26, 6, 30) {real, imag} */,
  {32'hc5395754, 32'h00000000} /* (26, 6, 29) {real, imag} */,
  {32'hc561cf0d, 32'h00000000} /* (26, 6, 28) {real, imag} */,
  {32'hc53042c0, 32'h00000000} /* (26, 6, 27) {real, imag} */,
  {32'hc4fb4eea, 32'h00000000} /* (26, 6, 26) {real, imag} */,
  {32'hc4ab6dd0, 32'h00000000} /* (26, 6, 25) {real, imag} */,
  {32'hc518c186, 32'h00000000} /* (26, 6, 24) {real, imag} */,
  {32'hc4a20bd6, 32'h00000000} /* (26, 6, 23) {real, imag} */,
  {32'hc45a6207, 32'h00000000} /* (26, 6, 22) {real, imag} */,
  {32'hc406ebfa, 32'h00000000} /* (26, 6, 21) {real, imag} */,
  {32'hc4a1c08b, 32'h00000000} /* (26, 6, 20) {real, imag} */,
  {32'hc479d8f4, 32'h00000000} /* (26, 6, 19) {real, imag} */,
  {32'hc4246500, 32'h00000000} /* (26, 6, 18) {real, imag} */,
  {32'hc49c0370, 32'h00000000} /* (26, 6, 17) {real, imag} */,
  {32'hc4257b13, 32'h00000000} /* (26, 6, 16) {real, imag} */,
  {32'hc2d45830, 32'h00000000} /* (26, 6, 15) {real, imag} */,
  {32'h40971d00, 32'h00000000} /* (26, 6, 14) {real, imag} */,
  {32'hc41874f6, 32'h00000000} /* (26, 6, 13) {real, imag} */,
  {32'h436dd8b0, 32'h00000000} /* (26, 6, 12) {real, imag} */,
  {32'hc397a2fc, 32'h00000000} /* (26, 6, 11) {real, imag} */,
  {32'h4449ca98, 32'h00000000} /* (26, 6, 10) {real, imag} */,
  {32'h4418cd87, 32'h00000000} /* (26, 6, 9) {real, imag} */,
  {32'h4472af08, 32'h00000000} /* (26, 6, 8) {real, imag} */,
  {32'hc24de380, 32'h00000000} /* (26, 6, 7) {real, imag} */,
  {32'hc448585b, 32'h00000000} /* (26, 6, 6) {real, imag} */,
  {32'hc44b69f2, 32'h00000000} /* (26, 6, 5) {real, imag} */,
  {32'hc4262472, 32'h00000000} /* (26, 6, 4) {real, imag} */,
  {32'hc4e03fa8, 32'h00000000} /* (26, 6, 3) {real, imag} */,
  {32'hc4d30176, 32'h00000000} /* (26, 6, 2) {real, imag} */,
  {32'hc5220096, 32'h00000000} /* (26, 6, 1) {real, imag} */,
  {32'hc5196e4f, 32'h00000000} /* (26, 6, 0) {real, imag} */,
  {32'hc5640451, 32'h00000000} /* (26, 5, 31) {real, imag} */,
  {32'hc5686a3a, 32'h00000000} /* (26, 5, 30) {real, imag} */,
  {32'hc53d4451, 32'h00000000} /* (26, 5, 29) {real, imag} */,
  {32'hc54281b0, 32'h00000000} /* (26, 5, 28) {real, imag} */,
  {32'hc5489a06, 32'h00000000} /* (26, 5, 27) {real, imag} */,
  {32'hc54128f5, 32'h00000000} /* (26, 5, 26) {real, imag} */,
  {32'hc555df09, 32'h00000000} /* (26, 5, 25) {real, imag} */,
  {32'hc51e5863, 32'h00000000} /* (26, 5, 24) {real, imag} */,
  {32'hc4f88927, 32'h00000000} /* (26, 5, 23) {real, imag} */,
  {32'hc4e26283, 32'h00000000} /* (26, 5, 22) {real, imag} */,
  {32'hc2f3feb8, 32'h00000000} /* (26, 5, 21) {real, imag} */,
  {32'hc44bd9de, 32'h00000000} /* (26, 5, 20) {real, imag} */,
  {32'hc4029862, 32'h00000000} /* (26, 5, 19) {real, imag} */,
  {32'hc4a37a39, 32'h00000000} /* (26, 5, 18) {real, imag} */,
  {32'h430921fc, 32'h00000000} /* (26, 5, 17) {real, imag} */,
  {32'hc4170a98, 32'h00000000} /* (26, 5, 16) {real, imag} */,
  {32'hc45dded4, 32'h00000000} /* (26, 5, 15) {real, imag} */,
  {32'hc320ee88, 32'h00000000} /* (26, 5, 14) {real, imag} */,
  {32'hc47ac135, 32'h00000000} /* (26, 5, 13) {real, imag} */,
  {32'h4262eee0, 32'h00000000} /* (26, 5, 12) {real, imag} */,
  {32'hc401231e, 32'h00000000} /* (26, 5, 11) {real, imag} */,
  {32'h43b50d30, 32'h00000000} /* (26, 5, 10) {real, imag} */,
  {32'h44899052, 32'h00000000} /* (26, 5, 9) {real, imag} */,
  {32'h44045529, 32'h00000000} /* (26, 5, 8) {real, imag} */,
  {32'hc3332da8, 32'h00000000} /* (26, 5, 7) {real, imag} */,
  {32'hc4e00135, 32'h00000000} /* (26, 5, 6) {real, imag} */,
  {32'hc4a78246, 32'h00000000} /* (26, 5, 5) {real, imag} */,
  {32'hc4ed3d5f, 32'h00000000} /* (26, 5, 4) {real, imag} */,
  {32'hc4d750bb, 32'h00000000} /* (26, 5, 3) {real, imag} */,
  {32'hc52246be, 32'h00000000} /* (26, 5, 2) {real, imag} */,
  {32'hc4bcf062, 32'h00000000} /* (26, 5, 1) {real, imag} */,
  {32'hc524378e, 32'h00000000} /* (26, 5, 0) {real, imag} */,
  {32'hc55eb312, 32'h00000000} /* (26, 4, 31) {real, imag} */,
  {32'hc56c42e2, 32'h00000000} /* (26, 4, 30) {real, imag} */,
  {32'hc5721c65, 32'h00000000} /* (26, 4, 29) {real, imag} */,
  {32'hc5839c2b, 32'h00000000} /* (26, 4, 28) {real, imag} */,
  {32'hc574e978, 32'h00000000} /* (26, 4, 27) {real, imag} */,
  {32'hc53d3fd7, 32'h00000000} /* (26, 4, 26) {real, imag} */,
  {32'hc5507166, 32'h00000000} /* (26, 4, 25) {real, imag} */,
  {32'hc54d3c8b, 32'h00000000} /* (26, 4, 24) {real, imag} */,
  {32'hc51f404e, 32'h00000000} /* (26, 4, 23) {real, imag} */,
  {32'hc4962a0e, 32'h00000000} /* (26, 4, 22) {real, imag} */,
  {32'h43932364, 32'h00000000} /* (26, 4, 21) {real, imag} */,
  {32'hc4116b03, 32'h00000000} /* (26, 4, 20) {real, imag} */,
  {32'hc486c3c1, 32'h00000000} /* (26, 4, 19) {real, imag} */,
  {32'hc3fc88bc, 32'h00000000} /* (26, 4, 18) {real, imag} */,
  {32'hc3ba8734, 32'h00000000} /* (26, 4, 17) {real, imag} */,
  {32'h43d7a4d4, 32'h00000000} /* (26, 4, 16) {real, imag} */,
  {32'h4402708a, 32'h00000000} /* (26, 4, 15) {real, imag} */,
  {32'hc413d7ba, 32'h00000000} /* (26, 4, 14) {real, imag} */,
  {32'h442cc8ac, 32'h00000000} /* (26, 4, 13) {real, imag} */,
  {32'h43ba28ac, 32'h00000000} /* (26, 4, 12) {real, imag} */,
  {32'h43df8f80, 32'h00000000} /* (26, 4, 11) {real, imag} */,
  {32'h439e9fd0, 32'h00000000} /* (26, 4, 10) {real, imag} */,
  {32'hc3c4e84c, 32'h00000000} /* (26, 4, 9) {real, imag} */,
  {32'h439bca68, 32'h00000000} /* (26, 4, 8) {real, imag} */,
  {32'hc3966b64, 32'h00000000} /* (26, 4, 7) {real, imag} */,
  {32'hc4a9fad0, 32'h00000000} /* (26, 4, 6) {real, imag} */,
  {32'h42fbe570, 32'h00000000} /* (26, 4, 5) {real, imag} */,
  {32'hc407c6b1, 32'h00000000} /* (26, 4, 4) {real, imag} */,
  {32'hc4fe5cc3, 32'h00000000} /* (26, 4, 3) {real, imag} */,
  {32'hc4caf6f7, 32'h00000000} /* (26, 4, 2) {real, imag} */,
  {32'hc51b678c, 32'h00000000} /* (26, 4, 1) {real, imag} */,
  {32'hc538b426, 32'h00000000} /* (26, 4, 0) {real, imag} */,
  {32'hc560f774, 32'h00000000} /* (26, 3, 31) {real, imag} */,
  {32'hc525c6de, 32'h00000000} /* (26, 3, 30) {real, imag} */,
  {32'hc5918f02, 32'h00000000} /* (26, 3, 29) {real, imag} */,
  {32'hc5732516, 32'h00000000} /* (26, 3, 28) {real, imag} */,
  {32'hc57ec86a, 32'h00000000} /* (26, 3, 27) {real, imag} */,
  {32'hc55eed02, 32'h00000000} /* (26, 3, 26) {real, imag} */,
  {32'hc54bdefa, 32'h00000000} /* (26, 3, 25) {real, imag} */,
  {32'hc5523d9f, 32'h00000000} /* (26, 3, 24) {real, imag} */,
  {32'hc53b5826, 32'h00000000} /* (26, 3, 23) {real, imag} */,
  {32'hc484a241, 32'h00000000} /* (26, 3, 22) {real, imag} */,
  {32'hc4a5d130, 32'h00000000} /* (26, 3, 21) {real, imag} */,
  {32'hc438de64, 32'h00000000} /* (26, 3, 20) {real, imag} */,
  {32'hc34b7418, 32'h00000000} /* (26, 3, 19) {real, imag} */,
  {32'h446aff4e, 32'h00000000} /* (26, 3, 18) {real, imag} */,
  {32'hc39f9ed0, 32'h00000000} /* (26, 3, 17) {real, imag} */,
  {32'h443720e0, 32'h00000000} /* (26, 3, 16) {real, imag} */,
  {32'h4452be56, 32'h00000000} /* (26, 3, 15) {real, imag} */,
  {32'h43a41e14, 32'h00000000} /* (26, 3, 14) {real, imag} */,
  {32'hc3277740, 32'h00000000} /* (26, 3, 13) {real, imag} */,
  {32'h44075950, 32'h00000000} /* (26, 3, 12) {real, imag} */,
  {32'h44a14655, 32'h00000000} /* (26, 3, 11) {real, imag} */,
  {32'hc3cfd42c, 32'h00000000} /* (26, 3, 10) {real, imag} */,
  {32'hc428403e, 32'h00000000} /* (26, 3, 9) {real, imag} */,
  {32'hc28f8f40, 32'h00000000} /* (26, 3, 8) {real, imag} */,
  {32'h440d4552, 32'h00000000} /* (26, 3, 7) {real, imag} */,
  {32'hc4913fdf, 32'h00000000} /* (26, 3, 6) {real, imag} */,
  {32'hc1b1cae0, 32'h00000000} /* (26, 3, 5) {real, imag} */,
  {32'hc4990639, 32'h00000000} /* (26, 3, 4) {real, imag} */,
  {32'hc4c248ef, 32'h00000000} /* (26, 3, 3) {real, imag} */,
  {32'hc48c5501, 32'h00000000} /* (26, 3, 2) {real, imag} */,
  {32'hc521490f, 32'h00000000} /* (26, 3, 1) {real, imag} */,
  {32'hc549d4b7, 32'h00000000} /* (26, 3, 0) {real, imag} */,
  {32'hc5453b1c, 32'h00000000} /* (26, 2, 31) {real, imag} */,
  {32'hc524093a, 32'h00000000} /* (26, 2, 30) {real, imag} */,
  {32'hc577d326, 32'h00000000} /* (26, 2, 29) {real, imag} */,
  {32'hc58ca2c9, 32'h00000000} /* (26, 2, 28) {real, imag} */,
  {32'hc584419a, 32'h00000000} /* (26, 2, 27) {real, imag} */,
  {32'hc56a4314, 32'h00000000} /* (26, 2, 26) {real, imag} */,
  {32'hc5460486, 32'h00000000} /* (26, 2, 25) {real, imag} */,
  {32'hc50a137a, 32'h00000000} /* (26, 2, 24) {real, imag} */,
  {32'hc50d2be6, 32'h00000000} /* (26, 2, 23) {real, imag} */,
  {32'hc4e883c5, 32'h00000000} /* (26, 2, 22) {real, imag} */,
  {32'hc428dbfa, 32'h00000000} /* (26, 2, 21) {real, imag} */,
  {32'hc44f5ad4, 32'h00000000} /* (26, 2, 20) {real, imag} */,
  {32'hc35a49ac, 32'h00000000} /* (26, 2, 19) {real, imag} */,
  {32'h431e9128, 32'h00000000} /* (26, 2, 18) {real, imag} */,
  {32'h44a56a0f, 32'h00000000} /* (26, 2, 17) {real, imag} */,
  {32'h44738640, 32'h00000000} /* (26, 2, 16) {real, imag} */,
  {32'h447453b0, 32'h00000000} /* (26, 2, 15) {real, imag} */,
  {32'h441f2672, 32'h00000000} /* (26, 2, 14) {real, imag} */,
  {32'h430b5df8, 32'h00000000} /* (26, 2, 13) {real, imag} */,
  {32'hc1ac4500, 32'h00000000} /* (26, 2, 12) {real, imag} */,
  {32'hc4161ee4, 32'h00000000} /* (26, 2, 11) {real, imag} */,
  {32'h41f90b00, 32'h00000000} /* (26, 2, 10) {real, imag} */,
  {32'hc29a4a50, 32'h00000000} /* (26, 2, 9) {real, imag} */,
  {32'hc48e9dc4, 32'h00000000} /* (26, 2, 8) {real, imag} */,
  {32'hc3db57dc, 32'h00000000} /* (26, 2, 7) {real, imag} */,
  {32'hc4be1483, 32'h00000000} /* (26, 2, 6) {real, imag} */,
  {32'hc5030ac4, 32'h00000000} /* (26, 2, 5) {real, imag} */,
  {32'hc4f6f40c, 32'h00000000} /* (26, 2, 4) {real, imag} */,
  {32'hc4d4716c, 32'h00000000} /* (26, 2, 3) {real, imag} */,
  {32'hc4eac845, 32'h00000000} /* (26, 2, 2) {real, imag} */,
  {32'hc52d7364, 32'h00000000} /* (26, 2, 1) {real, imag} */,
  {32'hc54500bc, 32'h00000000} /* (26, 2, 0) {real, imag} */,
  {32'hc56574d4, 32'h00000000} /* (26, 1, 31) {real, imag} */,
  {32'hc564a374, 32'h00000000} /* (26, 1, 30) {real, imag} */,
  {32'hc5840042, 32'h00000000} /* (26, 1, 29) {real, imag} */,
  {32'hc5916062, 32'h00000000} /* (26, 1, 28) {real, imag} */,
  {32'hc5609125, 32'h00000000} /* (26, 1, 27) {real, imag} */,
  {32'hc5561263, 32'h00000000} /* (26, 1, 26) {real, imag} */,
  {32'hc53a8d8a, 32'h00000000} /* (26, 1, 25) {real, imag} */,
  {32'hc4e2bd5a, 32'h00000000} /* (26, 1, 24) {real, imag} */,
  {32'hc51052e4, 32'h00000000} /* (26, 1, 23) {real, imag} */,
  {32'hc4f73748, 32'h00000000} /* (26, 1, 22) {real, imag} */,
  {32'hc4eb7bb0, 32'h00000000} /* (26, 1, 21) {real, imag} */,
  {32'hc2e1e68c, 32'h00000000} /* (26, 1, 20) {real, imag} */,
  {32'hc305468c, 32'h00000000} /* (26, 1, 19) {real, imag} */,
  {32'hc2ff08d0, 32'h00000000} /* (26, 1, 18) {real, imag} */,
  {32'h44bec048, 32'h00000000} /* (26, 1, 17) {real, imag} */,
  {32'h447bbd0c, 32'h00000000} /* (26, 1, 16) {real, imag} */,
  {32'hc399743c, 32'h00000000} /* (26, 1, 15) {real, imag} */,
  {32'hc3b5d680, 32'h00000000} /* (26, 1, 14) {real, imag} */,
  {32'h4384d278, 32'h00000000} /* (26, 1, 13) {real, imag} */,
  {32'h434722f0, 32'h00000000} /* (26, 1, 12) {real, imag} */,
  {32'h43a76850, 32'h00000000} /* (26, 1, 11) {real, imag} */,
  {32'hc44c081c, 32'h00000000} /* (26, 1, 10) {real, imag} */,
  {32'hc46a0de0, 32'h00000000} /* (26, 1, 9) {real, imag} */,
  {32'hc40c4a35, 32'h00000000} /* (26, 1, 8) {real, imag} */,
  {32'hc49b95be, 32'h00000000} /* (26, 1, 7) {real, imag} */,
  {32'hc52ba4c8, 32'h00000000} /* (26, 1, 6) {real, imag} */,
  {32'hc4fe9a9c, 32'h00000000} /* (26, 1, 5) {real, imag} */,
  {32'hc45e448c, 32'h00000000} /* (26, 1, 4) {real, imag} */,
  {32'hc4d7a884, 32'h00000000} /* (26, 1, 3) {real, imag} */,
  {32'hc51352a8, 32'h00000000} /* (26, 1, 2) {real, imag} */,
  {32'hc55092cc, 32'h00000000} /* (26, 1, 1) {real, imag} */,
  {32'hc559de1d, 32'h00000000} /* (26, 1, 0) {real, imag} */,
  {32'hc575f817, 32'h00000000} /* (26, 0, 31) {real, imag} */,
  {32'hc5633a7f, 32'h00000000} /* (26, 0, 30) {real, imag} */,
  {32'hc58214f6, 32'h00000000} /* (26, 0, 29) {real, imag} */,
  {32'hc586ff48, 32'h00000000} /* (26, 0, 28) {real, imag} */,
  {32'hc5841408, 32'h00000000} /* (26, 0, 27) {real, imag} */,
  {32'hc5651a43, 32'h00000000} /* (26, 0, 26) {real, imag} */,
  {32'hc554dcbf, 32'h00000000} /* (26, 0, 25) {real, imag} */,
  {32'hc53c6104, 32'h00000000} /* (26, 0, 24) {real, imag} */,
  {32'hc5052bb0, 32'h00000000} /* (26, 0, 23) {real, imag} */,
  {32'hc4f2b6c6, 32'h00000000} /* (26, 0, 22) {real, imag} */,
  {32'hc4c1e7e6, 32'h00000000} /* (26, 0, 21) {real, imag} */,
  {32'h43e9f8a8, 32'h00000000} /* (26, 0, 20) {real, imag} */,
  {32'h43c80da4, 32'h00000000} /* (26, 0, 19) {real, imag} */,
  {32'h4419c8ae, 32'h00000000} /* (26, 0, 18) {real, imag} */,
  {32'h447ed300, 32'h00000000} /* (26, 0, 17) {real, imag} */,
  {32'hc2c928c0, 32'h00000000} /* (26, 0, 16) {real, imag} */,
  {32'h41578200, 32'h00000000} /* (26, 0, 15) {real, imag} */,
  {32'h436ef130, 32'h00000000} /* (26, 0, 14) {real, imag} */,
  {32'hc2825760, 32'h00000000} /* (26, 0, 13) {real, imag} */,
  {32'hc350ea70, 32'h00000000} /* (26, 0, 12) {real, imag} */,
  {32'h42d779a0, 32'h00000000} /* (26, 0, 11) {real, imag} */,
  {32'hc44e87cc, 32'h00000000} /* (26, 0, 10) {real, imag} */,
  {32'hc441b55c, 32'h00000000} /* (26, 0, 9) {real, imag} */,
  {32'hc413bb10, 32'h00000000} /* (26, 0, 8) {real, imag} */,
  {32'hc512c852, 32'h00000000} /* (26, 0, 7) {real, imag} */,
  {32'hc510e9c3, 32'h00000000} /* (26, 0, 6) {real, imag} */,
  {32'hc4e1352e, 32'h00000000} /* (26, 0, 5) {real, imag} */,
  {32'hc4da11c8, 32'h00000000} /* (26, 0, 4) {real, imag} */,
  {32'hc51972e8, 32'h00000000} /* (26, 0, 3) {real, imag} */,
  {32'hc5424368, 32'h00000000} /* (26, 0, 2) {real, imag} */,
  {32'hc5547716, 32'h00000000} /* (26, 0, 1) {real, imag} */,
  {32'hc557b260, 32'h00000000} /* (26, 0, 0) {real, imag} */,
  {32'hc5d1a3dd, 32'h00000000} /* (25, 31, 31) {real, imag} */,
  {32'hc5ea9387, 32'h00000000} /* (25, 31, 30) {real, imag} */,
  {32'hc5ec4e4e, 32'h00000000} /* (25, 31, 29) {real, imag} */,
  {32'hc5f2c55a, 32'h00000000} /* (25, 31, 28) {real, imag} */,
  {32'hc5e5e296, 32'h00000000} /* (25, 31, 27) {real, imag} */,
  {32'hc5d97c24, 32'h00000000} /* (25, 31, 26) {real, imag} */,
  {32'hc5d82c9c, 32'h00000000} /* (25, 31, 25) {real, imag} */,
  {32'hc5bb4fd5, 32'h00000000} /* (25, 31, 24) {real, imag} */,
  {32'hc5b188b4, 32'h00000000} /* (25, 31, 23) {real, imag} */,
  {32'hc5887286, 32'h00000000} /* (25, 31, 22) {real, imag} */,
  {32'hc5461535, 32'h00000000} /* (25, 31, 21) {real, imag} */,
  {32'hc497ea61, 32'h00000000} /* (25, 31, 20) {real, imag} */,
  {32'hc09a8a00, 32'h00000000} /* (25, 31, 19) {real, imag} */,
  {32'h44774fc4, 32'h00000000} /* (25, 31, 18) {real, imag} */,
  {32'h4494befc, 32'h00000000} /* (25, 31, 17) {real, imag} */,
  {32'h449c4bda, 32'h00000000} /* (25, 31, 16) {real, imag} */,
  {32'h44f0392c, 32'h00000000} /* (25, 31, 15) {real, imag} */,
  {32'h4506036a, 32'h00000000} /* (25, 31, 14) {real, imag} */,
  {32'h452e0c05, 32'h00000000} /* (25, 31, 13) {real, imag} */,
  {32'h44ecedb0, 32'h00000000} /* (25, 31, 12) {real, imag} */,
  {32'h4491c496, 32'h00000000} /* (25, 31, 11) {real, imag} */,
  {32'h439da3e0, 32'h00000000} /* (25, 31, 10) {real, imag} */,
  {32'hc453e614, 32'h00000000} /* (25, 31, 9) {real, imag} */,
  {32'hc4c6c294, 32'h00000000} /* (25, 31, 8) {real, imag} */,
  {32'hc52dc631, 32'h00000000} /* (25, 31, 7) {real, imag} */,
  {32'hc53709d7, 32'h00000000} /* (25, 31, 6) {real, imag} */,
  {32'hc5860c3a, 32'h00000000} /* (25, 31, 5) {real, imag} */,
  {32'hc59422ba, 32'h00000000} /* (25, 31, 4) {real, imag} */,
  {32'hc5ac3c8e, 32'h00000000} /* (25, 31, 3) {real, imag} */,
  {32'hc5b192ce, 32'h00000000} /* (25, 31, 2) {real, imag} */,
  {32'hc5e27e49, 32'h00000000} /* (25, 31, 1) {real, imag} */,
  {32'hc5ccc3c4, 32'h00000000} /* (25, 31, 0) {real, imag} */,
  {32'hc5d2a7be, 32'h00000000} /* (25, 30, 31) {real, imag} */,
  {32'hc5e9319c, 32'h00000000} /* (25, 30, 30) {real, imag} */,
  {32'hc5f7fbab, 32'h00000000} /* (25, 30, 29) {real, imag} */,
  {32'hc5f9007e, 32'h00000000} /* (25, 30, 28) {real, imag} */,
  {32'hc5dd783c, 32'h00000000} /* (25, 30, 27) {real, imag} */,
  {32'hc5f02fa2, 32'h00000000} /* (25, 30, 26) {real, imag} */,
  {32'hc5ded9fd, 32'h00000000} /* (25, 30, 25) {real, imag} */,
  {32'hc5e46c1a, 32'h00000000} /* (25, 30, 24) {real, imag} */,
  {32'hc5c23d76, 32'h00000000} /* (25, 30, 23) {real, imag} */,
  {32'hc57e6b64, 32'h00000000} /* (25, 30, 22) {real, imag} */,
  {32'hc52732b0, 32'h00000000} /* (25, 30, 21) {real, imag} */,
  {32'hc3253f60, 32'h00000000} /* (25, 30, 20) {real, imag} */,
  {32'h43f89800, 32'h00000000} /* (25, 30, 19) {real, imag} */,
  {32'h44f59798, 32'h00000000} /* (25, 30, 18) {real, imag} */,
  {32'h45025d9f, 32'h00000000} /* (25, 30, 17) {real, imag} */,
  {32'h45389e44, 32'h00000000} /* (25, 30, 16) {real, imag} */,
  {32'h454da875, 32'h00000000} /* (25, 30, 15) {real, imag} */,
  {32'h452a98cc, 32'h00000000} /* (25, 30, 14) {real, imag} */,
  {32'h4553a4c2, 32'h00000000} /* (25, 30, 13) {real, imag} */,
  {32'h44f554c8, 32'h00000000} /* (25, 30, 12) {real, imag} */,
  {32'h449ec09a, 32'h00000000} /* (25, 30, 11) {real, imag} */,
  {32'hc39a01b8, 32'h00000000} /* (25, 30, 10) {real, imag} */,
  {32'hc4ce004c, 32'h00000000} /* (25, 30, 9) {real, imag} */,
  {32'hc51f1cbb, 32'h00000000} /* (25, 30, 8) {real, imag} */,
  {32'hc5668043, 32'h00000000} /* (25, 30, 7) {real, imag} */,
  {32'hc58a39a2, 32'h00000000} /* (25, 30, 6) {real, imag} */,
  {32'hc59490ea, 32'h00000000} /* (25, 30, 5) {real, imag} */,
  {32'hc5aca8ab, 32'h00000000} /* (25, 30, 4) {real, imag} */,
  {32'hc5baa229, 32'h00000000} /* (25, 30, 3) {real, imag} */,
  {32'hc5bd9be7, 32'h00000000} /* (25, 30, 2) {real, imag} */,
  {32'hc5e3802c, 32'h00000000} /* (25, 30, 1) {real, imag} */,
  {32'hc5d78580, 32'h00000000} /* (25, 30, 0) {real, imag} */,
  {32'hc5d79e96, 32'h00000000} /* (25, 29, 31) {real, imag} */,
  {32'hc5f220d4, 32'h00000000} /* (25, 29, 30) {real, imag} */,
  {32'hc5f3cef7, 32'h00000000} /* (25, 29, 29) {real, imag} */,
  {32'hc5eeaee5, 32'h00000000} /* (25, 29, 28) {real, imag} */,
  {32'hc605c500, 32'h00000000} /* (25, 29, 27) {real, imag} */,
  {32'hc609e38c, 32'h00000000} /* (25, 29, 26) {real, imag} */,
  {32'hc5f5d301, 32'h00000000} /* (25, 29, 25) {real, imag} */,
  {32'hc5d50211, 32'h00000000} /* (25, 29, 24) {real, imag} */,
  {32'hc5a3aef9, 32'h00000000} /* (25, 29, 23) {real, imag} */,
  {32'hc5909b29, 32'h00000000} /* (25, 29, 22) {real, imag} */,
  {32'hc5775046, 32'h00000000} /* (25, 29, 21) {real, imag} */,
  {32'hc22ec180, 32'h00000000} /* (25, 29, 20) {real, imag} */,
  {32'h441e1644, 32'h00000000} /* (25, 29, 19) {real, imag} */,
  {32'h44e8d550, 32'h00000000} /* (25, 29, 18) {real, imag} */,
  {32'h45154b4e, 32'h00000000} /* (25, 29, 17) {real, imag} */,
  {32'h45016092, 32'h00000000} /* (25, 29, 16) {real, imag} */,
  {32'h452ff4db, 32'h00000000} /* (25, 29, 15) {real, imag} */,
  {32'h4530a810, 32'h00000000} /* (25, 29, 14) {real, imag} */,
  {32'h44fa6e4c, 32'h00000000} /* (25, 29, 13) {real, imag} */,
  {32'h44eb7cac, 32'h00000000} /* (25, 29, 12) {real, imag} */,
  {32'h44b1af4a, 32'h00000000} /* (25, 29, 11) {real, imag} */,
  {32'hc48dbaf0, 32'h00000000} /* (25, 29, 10) {real, imag} */,
  {32'hc4de64e4, 32'h00000000} /* (25, 29, 9) {real, imag} */,
  {32'hc5555bb6, 32'h00000000} /* (25, 29, 8) {real, imag} */,
  {32'hc58b7c33, 32'h00000000} /* (25, 29, 7) {real, imag} */,
  {32'hc5781312, 32'h00000000} /* (25, 29, 6) {real, imag} */,
  {32'hc5787f22, 32'h00000000} /* (25, 29, 5) {real, imag} */,
  {32'hc59282c3, 32'h00000000} /* (25, 29, 4) {real, imag} */,
  {32'hc5c4f01c, 32'h00000000} /* (25, 29, 3) {real, imag} */,
  {32'hc5e3adea, 32'h00000000} /* (25, 29, 2) {real, imag} */,
  {32'hc5d31c09, 32'h00000000} /* (25, 29, 1) {real, imag} */,
  {32'hc5beea4d, 32'h00000000} /* (25, 29, 0) {real, imag} */,
  {32'hc5cfb982, 32'h00000000} /* (25, 28, 31) {real, imag} */,
  {32'hc6047e4a, 32'h00000000} /* (25, 28, 30) {real, imag} */,
  {32'hc5fcce2e, 32'h00000000} /* (25, 28, 29) {real, imag} */,
  {32'hc5f68970, 32'h00000000} /* (25, 28, 28) {real, imag} */,
  {32'hc60731d2, 32'h00000000} /* (25, 28, 27) {real, imag} */,
  {32'hc600a7e1, 32'h00000000} /* (25, 28, 26) {real, imag} */,
  {32'hc5fcc8bc, 32'h00000000} /* (25, 28, 25) {real, imag} */,
  {32'hc5ce54d0, 32'h00000000} /* (25, 28, 24) {real, imag} */,
  {32'hc5b82bcd, 32'h00000000} /* (25, 28, 23) {real, imag} */,
  {32'hc590802c, 32'h00000000} /* (25, 28, 22) {real, imag} */,
  {32'hc581f055, 32'h00000000} /* (25, 28, 21) {real, imag} */,
  {32'hc41bbb24, 32'h00000000} /* (25, 28, 20) {real, imag} */,
  {32'h444156a4, 32'h00000000} /* (25, 28, 19) {real, imag} */,
  {32'h45550e8e, 32'h00000000} /* (25, 28, 18) {real, imag} */,
  {32'h4530311a, 32'h00000000} /* (25, 28, 17) {real, imag} */,
  {32'h4514fe5e, 32'h00000000} /* (25, 28, 16) {real, imag} */,
  {32'h4517c3f4, 32'h00000000} /* (25, 28, 15) {real, imag} */,
  {32'h452c4cba, 32'h00000000} /* (25, 28, 14) {real, imag} */,
  {32'h44e78000, 32'h00000000} /* (25, 28, 13) {real, imag} */,
  {32'h451bceb1, 32'h00000000} /* (25, 28, 12) {real, imag} */,
  {32'h44a4ca04, 32'h00000000} /* (25, 28, 11) {real, imag} */,
  {32'hc481f786, 32'h00000000} /* (25, 28, 10) {real, imag} */,
  {32'hc50f3f28, 32'h00000000} /* (25, 28, 9) {real, imag} */,
  {32'hc5607328, 32'h00000000} /* (25, 28, 8) {real, imag} */,
  {32'hc5810045, 32'h00000000} /* (25, 28, 7) {real, imag} */,
  {32'hc588b0b2, 32'h00000000} /* (25, 28, 6) {real, imag} */,
  {32'hc5b94e0d, 32'h00000000} /* (25, 28, 5) {real, imag} */,
  {32'hc5b7afe8, 32'h00000000} /* (25, 28, 4) {real, imag} */,
  {32'hc5ccf95c, 32'h00000000} /* (25, 28, 3) {real, imag} */,
  {32'hc5da20cb, 32'h00000000} /* (25, 28, 2) {real, imag} */,
  {32'hc5f27931, 32'h00000000} /* (25, 28, 1) {real, imag} */,
  {32'hc5de3903, 32'h00000000} /* (25, 28, 0) {real, imag} */,
  {32'hc5c62cbb, 32'h00000000} /* (25, 27, 31) {real, imag} */,
  {32'hc5e07ebc, 32'h00000000} /* (25, 27, 30) {real, imag} */,
  {32'hc5e9656e, 32'h00000000} /* (25, 27, 29) {real, imag} */,
  {32'hc5fad791, 32'h00000000} /* (25, 27, 28) {real, imag} */,
  {32'hc608646d, 32'h00000000} /* (25, 27, 27) {real, imag} */,
  {32'hc60175e6, 32'h00000000} /* (25, 27, 26) {real, imag} */,
  {32'hc5f5f78e, 32'h00000000} /* (25, 27, 25) {real, imag} */,
  {32'hc5d9c33e, 32'h00000000} /* (25, 27, 24) {real, imag} */,
  {32'hc59b337a, 32'h00000000} /* (25, 27, 23) {real, imag} */,
  {32'hc58ddf13, 32'h00000000} /* (25, 27, 22) {real, imag} */,
  {32'hc54fc078, 32'h00000000} /* (25, 27, 21) {real, imag} */,
  {32'hc39f32a0, 32'h00000000} /* (25, 27, 20) {real, imag} */,
  {32'h44c308f0, 32'h00000000} /* (25, 27, 19) {real, imag} */,
  {32'h454214f2, 32'h00000000} /* (25, 27, 18) {real, imag} */,
  {32'h45385012, 32'h00000000} /* (25, 27, 17) {real, imag} */,
  {32'h45416825, 32'h00000000} /* (25, 27, 16) {real, imag} */,
  {32'h4544190e, 32'h00000000} /* (25, 27, 15) {real, imag} */,
  {32'h44f5162e, 32'h00000000} /* (25, 27, 14) {real, imag} */,
  {32'h45058d54, 32'h00000000} /* (25, 27, 13) {real, imag} */,
  {32'h44b533f4, 32'h00000000} /* (25, 27, 12) {real, imag} */,
  {32'h448f0428, 32'h00000000} /* (25, 27, 11) {real, imag} */,
  {32'hc48f83e0, 32'h00000000} /* (25, 27, 10) {real, imag} */,
  {32'hc587723c, 32'h00000000} /* (25, 27, 9) {real, imag} */,
  {32'hc567572b, 32'h00000000} /* (25, 27, 8) {real, imag} */,
  {32'hc5794e3c, 32'h00000000} /* (25, 27, 7) {real, imag} */,
  {32'hc59bdc3d, 32'h00000000} /* (25, 27, 6) {real, imag} */,
  {32'hc5b223ae, 32'h00000000} /* (25, 27, 5) {real, imag} */,
  {32'hc5dbe588, 32'h00000000} /* (25, 27, 4) {real, imag} */,
  {32'hc5f84230, 32'h00000000} /* (25, 27, 3) {real, imag} */,
  {32'hc5d34ae1, 32'h00000000} /* (25, 27, 2) {real, imag} */,
  {32'hc5dacf91, 32'h00000000} /* (25, 27, 1) {real, imag} */,
  {32'hc5d7d4dc, 32'h00000000} /* (25, 27, 0) {real, imag} */,
  {32'hc5c7e642, 32'h00000000} /* (25, 26, 31) {real, imag} */,
  {32'hc5e49582, 32'h00000000} /* (25, 26, 30) {real, imag} */,
  {32'hc60571ad, 32'h00000000} /* (25, 26, 29) {real, imag} */,
  {32'hc5fdc9bb, 32'h00000000} /* (25, 26, 28) {real, imag} */,
  {32'hc5e7fe98, 32'h00000000} /* (25, 26, 27) {real, imag} */,
  {32'hc5e13286, 32'h00000000} /* (25, 26, 26) {real, imag} */,
  {32'hc5e6b2cd, 32'h00000000} /* (25, 26, 25) {real, imag} */,
  {32'hc5afa3dd, 32'h00000000} /* (25, 26, 24) {real, imag} */,
  {32'hc58ba7cf, 32'h00000000} /* (25, 26, 23) {real, imag} */,
  {32'hc54fc83a, 32'h00000000} /* (25, 26, 22) {real, imag} */,
  {32'hc5293e14, 32'h00000000} /* (25, 26, 21) {real, imag} */,
  {32'hc3939670, 32'h00000000} /* (25, 26, 20) {real, imag} */,
  {32'h44d80c92, 32'h00000000} /* (25, 26, 19) {real, imag} */,
  {32'h452f710c, 32'h00000000} /* (25, 26, 18) {real, imag} */,
  {32'h451f33f6, 32'h00000000} /* (25, 26, 17) {real, imag} */,
  {32'h454766d4, 32'h00000000} /* (25, 26, 16) {real, imag} */,
  {32'h452ffac0, 32'h00000000} /* (25, 26, 15) {real, imag} */,
  {32'h4520c8c9, 32'h00000000} /* (25, 26, 14) {real, imag} */,
  {32'h44ec2eb6, 32'h00000000} /* (25, 26, 13) {real, imag} */,
  {32'h448d770c, 32'h00000000} /* (25, 26, 12) {real, imag} */,
  {32'h440fb094, 32'h00000000} /* (25, 26, 11) {real, imag} */,
  {32'hc4ab66de, 32'h00000000} /* (25, 26, 10) {real, imag} */,
  {32'hc56fdcde, 32'h00000000} /* (25, 26, 9) {real, imag} */,
  {32'hc571ca66, 32'h00000000} /* (25, 26, 8) {real, imag} */,
  {32'hc588ad0d, 32'h00000000} /* (25, 26, 7) {real, imag} */,
  {32'hc58b5dbc, 32'h00000000} /* (25, 26, 6) {real, imag} */,
  {32'hc5afc140, 32'h00000000} /* (25, 26, 5) {real, imag} */,
  {32'hc5aa591f, 32'h00000000} /* (25, 26, 4) {real, imag} */,
  {32'hc5baeb4a, 32'h00000000} /* (25, 26, 3) {real, imag} */,
  {32'hc5d171b6, 32'h00000000} /* (25, 26, 2) {real, imag} */,
  {32'hc5cb0381, 32'h00000000} /* (25, 26, 1) {real, imag} */,
  {32'hc5c71b88, 32'h00000000} /* (25, 26, 0) {real, imag} */,
  {32'hc5cf70e9, 32'h00000000} /* (25, 25, 31) {real, imag} */,
  {32'hc5e5daae, 32'h00000000} /* (25, 25, 30) {real, imag} */,
  {32'hc5ed9766, 32'h00000000} /* (25, 25, 29) {real, imag} */,
  {32'hc5d4b090, 32'h00000000} /* (25, 25, 28) {real, imag} */,
  {32'hc5e8525a, 32'h00000000} /* (25, 25, 27) {real, imag} */,
  {32'hc5cff561, 32'h00000000} /* (25, 25, 26) {real, imag} */,
  {32'hc5ae386e, 32'h00000000} /* (25, 25, 25) {real, imag} */,
  {32'hc5b440ca, 32'h00000000} /* (25, 25, 24) {real, imag} */,
  {32'hc586f453, 32'h00000000} /* (25, 25, 23) {real, imag} */,
  {32'hc5551bcf, 32'h00000000} /* (25, 25, 22) {real, imag} */,
  {32'hc4812b88, 32'h00000000} /* (25, 25, 21) {real, imag} */,
  {32'h44d522b8, 32'h00000000} /* (25, 25, 20) {real, imag} */,
  {32'h4466f9d8, 32'h00000000} /* (25, 25, 19) {real, imag} */,
  {32'h45282e2c, 32'h00000000} /* (25, 25, 18) {real, imag} */,
  {32'h45078ed2, 32'h00000000} /* (25, 25, 17) {real, imag} */,
  {32'h45494314, 32'h00000000} /* (25, 25, 16) {real, imag} */,
  {32'h452eed1e, 32'h00000000} /* (25, 25, 15) {real, imag} */,
  {32'h454bbe94, 32'h00000000} /* (25, 25, 14) {real, imag} */,
  {32'h45442b00, 32'h00000000} /* (25, 25, 13) {real, imag} */,
  {32'h44bdfb28, 32'h00000000} /* (25, 25, 12) {real, imag} */,
  {32'hc34b9b40, 32'h00000000} /* (25, 25, 11) {real, imag} */,
  {32'hc50b52ee, 32'h00000000} /* (25, 25, 10) {real, imag} */,
  {32'hc55222f0, 32'h00000000} /* (25, 25, 9) {real, imag} */,
  {32'hc58dd020, 32'h00000000} /* (25, 25, 8) {real, imag} */,
  {32'hc5775c06, 32'h00000000} /* (25, 25, 7) {real, imag} */,
  {32'hc591b252, 32'h00000000} /* (25, 25, 6) {real, imag} */,
  {32'hc59815ca, 32'h00000000} /* (25, 25, 5) {real, imag} */,
  {32'hc5a90558, 32'h00000000} /* (25, 25, 4) {real, imag} */,
  {32'hc5b8079f, 32'h00000000} /* (25, 25, 3) {real, imag} */,
  {32'hc5b4df00, 32'h00000000} /* (25, 25, 2) {real, imag} */,
  {32'hc5c32541, 32'h00000000} /* (25, 25, 1) {real, imag} */,
  {32'hc5c97478, 32'h00000000} /* (25, 25, 0) {real, imag} */,
  {32'hc5b3c6b0, 32'h00000000} /* (25, 24, 31) {real, imag} */,
  {32'hc5c541eb, 32'h00000000} /* (25, 24, 30) {real, imag} */,
  {32'hc5bc0591, 32'h00000000} /* (25, 24, 29) {real, imag} */,
  {32'hc5b58aee, 32'h00000000} /* (25, 24, 28) {real, imag} */,
  {32'hc5b0d6d6, 32'h00000000} /* (25, 24, 27) {real, imag} */,
  {32'hc5aa1bec, 32'h00000000} /* (25, 24, 26) {real, imag} */,
  {32'hc5bbd3aa, 32'h00000000} /* (25, 24, 25) {real, imag} */,
  {32'hc59b3481, 32'h00000000} /* (25, 24, 24) {real, imag} */,
  {32'hc567270a, 32'h00000000} /* (25, 24, 23) {real, imag} */,
  {32'hc553c40c, 32'h00000000} /* (25, 24, 22) {real, imag} */,
  {32'hc4949746, 32'h00000000} /* (25, 24, 21) {real, imag} */,
  {32'h442d3f0c, 32'h00000000} /* (25, 24, 20) {real, imag} */,
  {32'h44cab9be, 32'h00000000} /* (25, 24, 19) {real, imag} */,
  {32'h451c38fb, 32'h00000000} /* (25, 24, 18) {real, imag} */,
  {32'h4509f9ca, 32'h00000000} /* (25, 24, 17) {real, imag} */,
  {32'h45116308, 32'h00000000} /* (25, 24, 16) {real, imag} */,
  {32'h45424da0, 32'h00000000} /* (25, 24, 15) {real, imag} */,
  {32'h45626ba2, 32'h00000000} /* (25, 24, 14) {real, imag} */,
  {32'h4523b6de, 32'h00000000} /* (25, 24, 13) {real, imag} */,
  {32'h44a4093c, 32'h00000000} /* (25, 24, 12) {real, imag} */,
  {32'hc3d9c348, 32'h00000000} /* (25, 24, 11) {real, imag} */,
  {32'hc508584b, 32'h00000000} /* (25, 24, 10) {real, imag} */,
  {32'hc55ab678, 32'h00000000} /* (25, 24, 9) {real, imag} */,
  {32'hc54dfc0a, 32'h00000000} /* (25, 24, 8) {real, imag} */,
  {32'hc56620b6, 32'h00000000} /* (25, 24, 7) {real, imag} */,
  {32'hc58be57c, 32'h00000000} /* (25, 24, 6) {real, imag} */,
  {32'hc5882f42, 32'h00000000} /* (25, 24, 5) {real, imag} */,
  {32'hc5a1675a, 32'h00000000} /* (25, 24, 4) {real, imag} */,
  {32'hc5b27272, 32'h00000000} /* (25, 24, 3) {real, imag} */,
  {32'hc5ac54cc, 32'h00000000} /* (25, 24, 2) {real, imag} */,
  {32'hc5c6d70d, 32'h00000000} /* (25, 24, 1) {real, imag} */,
  {32'hc5b0227a, 32'h00000000} /* (25, 24, 0) {real, imag} */,
  {32'hc584a44a, 32'h00000000} /* (25, 23, 31) {real, imag} */,
  {32'hc58ceee2, 32'h00000000} /* (25, 23, 30) {real, imag} */,
  {32'hc5b8a76c, 32'h00000000} /* (25, 23, 29) {real, imag} */,
  {32'hc5a8b82e, 32'h00000000} /* (25, 23, 28) {real, imag} */,
  {32'hc59f5346, 32'h00000000} /* (25, 23, 27) {real, imag} */,
  {32'hc599b70e, 32'h00000000} /* (25, 23, 26) {real, imag} */,
  {32'hc5ae769c, 32'h00000000} /* (25, 23, 25) {real, imag} */,
  {32'hc560e50a, 32'h00000000} /* (25, 23, 24) {real, imag} */,
  {32'hc57fc932, 32'h00000000} /* (25, 23, 23) {real, imag} */,
  {32'hc5633cfe, 32'h00000000} /* (25, 23, 22) {real, imag} */,
  {32'hc42b7e64, 32'h00000000} /* (25, 23, 21) {real, imag} */,
  {32'h44b88f71, 32'h00000000} /* (25, 23, 20) {real, imag} */,
  {32'h44ca4bf1, 32'h00000000} /* (25, 23, 19) {real, imag} */,
  {32'h44feff26, 32'h00000000} /* (25, 23, 18) {real, imag} */,
  {32'h454dfb48, 32'h00000000} /* (25, 23, 17) {real, imag} */,
  {32'h452859b1, 32'h00000000} /* (25, 23, 16) {real, imag} */,
  {32'h456f2484, 32'h00000000} /* (25, 23, 15) {real, imag} */,
  {32'h4562f39f, 32'h00000000} /* (25, 23, 14) {real, imag} */,
  {32'h44dcfcb2, 32'h00000000} /* (25, 23, 13) {real, imag} */,
  {32'h44a68729, 32'h00000000} /* (25, 23, 12) {real, imag} */,
  {32'h42a1c3e0, 32'h00000000} /* (25, 23, 11) {real, imag} */,
  {32'hc4d3263f, 32'h00000000} /* (25, 23, 10) {real, imag} */,
  {32'hc512daf8, 32'h00000000} /* (25, 23, 9) {real, imag} */,
  {32'hc51b1402, 32'h00000000} /* (25, 23, 8) {real, imag} */,
  {32'hc528dee2, 32'h00000000} /* (25, 23, 7) {real, imag} */,
  {32'hc58a637b, 32'h00000000} /* (25, 23, 6) {real, imag} */,
  {32'hc59bb750, 32'h00000000} /* (25, 23, 5) {real, imag} */,
  {32'hc5a15444, 32'h00000000} /* (25, 23, 4) {real, imag} */,
  {32'hc584072e, 32'h00000000} /* (25, 23, 3) {real, imag} */,
  {32'hc5927b80, 32'h00000000} /* (25, 23, 2) {real, imag} */,
  {32'hc5b0a340, 32'h00000000} /* (25, 23, 1) {real, imag} */,
  {32'hc59b1ee0, 32'h00000000} /* (25, 23, 0) {real, imag} */,
  {32'hc5739b38, 32'h00000000} /* (25, 22, 31) {real, imag} */,
  {32'hc58113c7, 32'h00000000} /* (25, 22, 30) {real, imag} */,
  {32'hc5742457, 32'h00000000} /* (25, 22, 29) {real, imag} */,
  {32'hc58d09d7, 32'h00000000} /* (25, 22, 28) {real, imag} */,
  {32'hc555c158, 32'h00000000} /* (25, 22, 27) {real, imag} */,
  {32'hc56e05b2, 32'h00000000} /* (25, 22, 26) {real, imag} */,
  {32'hc54c42b6, 32'h00000000} /* (25, 22, 25) {real, imag} */,
  {32'hc55db48a, 32'h00000000} /* (25, 22, 24) {real, imag} */,
  {32'hc531cbc9, 32'h00000000} /* (25, 22, 23) {real, imag} */,
  {32'hc503de3e, 32'h00000000} /* (25, 22, 22) {real, imag} */,
  {32'hc455f93c, 32'h00000000} /* (25, 22, 21) {real, imag} */,
  {32'h447c6eda, 32'h00000000} /* (25, 22, 20) {real, imag} */,
  {32'h44c7c861, 32'h00000000} /* (25, 22, 19) {real, imag} */,
  {32'h45437f9a, 32'h00000000} /* (25, 22, 18) {real, imag} */,
  {32'h450c2588, 32'h00000000} /* (25, 22, 17) {real, imag} */,
  {32'h45136427, 32'h00000000} /* (25, 22, 16) {real, imag} */,
  {32'h4530bef2, 32'h00000000} /* (25, 22, 15) {real, imag} */,
  {32'h450dd80d, 32'h00000000} /* (25, 22, 14) {real, imag} */,
  {32'h45460723, 32'h00000000} /* (25, 22, 13) {real, imag} */,
  {32'h44e2cecf, 32'h00000000} /* (25, 22, 12) {real, imag} */,
  {32'h448d6d3f, 32'h00000000} /* (25, 22, 11) {real, imag} */,
  {32'hc47cb1e2, 32'h00000000} /* (25, 22, 10) {real, imag} */,
  {32'hc509d5d6, 32'h00000000} /* (25, 22, 9) {real, imag} */,
  {32'hc51feda4, 32'h00000000} /* (25, 22, 8) {real, imag} */,
  {32'hc55316f7, 32'h00000000} /* (25, 22, 7) {real, imag} */,
  {32'hc5544966, 32'h00000000} /* (25, 22, 6) {real, imag} */,
  {32'hc58dd53e, 32'h00000000} /* (25, 22, 5) {real, imag} */,
  {32'hc55d9d68, 32'h00000000} /* (25, 22, 4) {real, imag} */,
  {32'hc578f342, 32'h00000000} /* (25, 22, 3) {real, imag} */,
  {32'hc55cb5fc, 32'h00000000} /* (25, 22, 2) {real, imag} */,
  {32'hc537dcb4, 32'h00000000} /* (25, 22, 1) {real, imag} */,
  {32'hc5575f19, 32'h00000000} /* (25, 22, 0) {real, imag} */,
  {32'hc5116d40, 32'h00000000} /* (25, 21, 31) {real, imag} */,
  {32'hc5302a4f, 32'h00000000} /* (25, 21, 30) {real, imag} */,
  {32'hc4eb63d8, 32'h00000000} /* (25, 21, 29) {real, imag} */,
  {32'hc4ebd0e8, 32'h00000000} /* (25, 21, 28) {real, imag} */,
  {32'hc52f6873, 32'h00000000} /* (25, 21, 27) {real, imag} */,
  {32'hc4f0d0bd, 32'h00000000} /* (25, 21, 26) {real, imag} */,
  {32'hc4f1b396, 32'h00000000} /* (25, 21, 25) {real, imag} */,
  {32'hc4b9a5d6, 32'h00000000} /* (25, 21, 24) {real, imag} */,
  {32'hc4b0b45e, 32'h00000000} /* (25, 21, 23) {real, imag} */,
  {32'hc36ed088, 32'h00000000} /* (25, 21, 22) {real, imag} */,
  {32'h42217ee0, 32'h00000000} /* (25, 21, 21) {real, imag} */,
  {32'h43f7f6a8, 32'h00000000} /* (25, 21, 20) {real, imag} */,
  {32'h43538078, 32'h00000000} /* (25, 21, 19) {real, imag} */,
  {32'h442273cf, 32'h00000000} /* (25, 21, 18) {real, imag} */,
  {32'h44f5befa, 32'h00000000} /* (25, 21, 17) {real, imag} */,
  {32'h445ec162, 32'h00000000} /* (25, 21, 16) {real, imag} */,
  {32'h44bcf526, 32'h00000000} /* (25, 21, 15) {real, imag} */,
  {32'h44e74756, 32'h00000000} /* (25, 21, 14) {real, imag} */,
  {32'h44c58b5e, 32'h00000000} /* (25, 21, 13) {real, imag} */,
  {32'h44ea0cce, 32'h00000000} /* (25, 21, 12) {real, imag} */,
  {32'h4421953c, 32'h00000000} /* (25, 21, 11) {real, imag} */,
  {32'hc4922873, 32'h00000000} /* (25, 21, 10) {real, imag} */,
  {32'hc559a819, 32'h00000000} /* (25, 21, 9) {real, imag} */,
  {32'hc508a371, 32'h00000000} /* (25, 21, 8) {real, imag} */,
  {32'hc519efa0, 32'h00000000} /* (25, 21, 7) {real, imag} */,
  {32'hc48b590f, 32'h00000000} /* (25, 21, 6) {real, imag} */,
  {32'hc4d0b1ed, 32'h00000000} /* (25, 21, 5) {real, imag} */,
  {32'hc4c1c834, 32'h00000000} /* (25, 21, 4) {real, imag} */,
  {32'hc4c5b387, 32'h00000000} /* (25, 21, 3) {real, imag} */,
  {32'hc4937d18, 32'h00000000} /* (25, 21, 2) {real, imag} */,
  {32'hc4e3aa0c, 32'h00000000} /* (25, 21, 1) {real, imag} */,
  {32'hc486969d, 32'h00000000} /* (25, 21, 0) {real, imag} */,
  {32'h4386fe66, 32'h00000000} /* (25, 20, 31) {real, imag} */,
  {32'h42b7678c, 32'h00000000} /* (25, 20, 30) {real, imag} */,
  {32'h444d6ed0, 32'h00000000} /* (25, 20, 29) {real, imag} */,
  {32'h442dfec6, 32'h00000000} /* (25, 20, 28) {real, imag} */,
  {32'h4482a11d, 32'h00000000} /* (25, 20, 27) {real, imag} */,
  {32'h43f0554b, 32'h00000000} /* (25, 20, 26) {real, imag} */,
  {32'h428bcd94, 32'h00000000} /* (25, 20, 25) {real, imag} */,
  {32'h43d03b06, 32'h00000000} /* (25, 20, 24) {real, imag} */,
  {32'h44d103e8, 32'h00000000} /* (25, 20, 23) {real, imag} */,
  {32'h44bfb77c, 32'h00000000} /* (25, 20, 22) {real, imag} */,
  {32'h449d9ae8, 32'h00000000} /* (25, 20, 21) {real, imag} */,
  {32'hc35fefd4, 32'h00000000} /* (25, 20, 20) {real, imag} */,
  {32'hc484497c, 32'h00000000} /* (25, 20, 19) {real, imag} */,
  {32'hc45c43c2, 32'h00000000} /* (25, 20, 18) {real, imag} */,
  {32'hc385d8ea, 32'h00000000} /* (25, 20, 17) {real, imag} */,
  {32'hc4557a51, 32'h00000000} /* (25, 20, 16) {real, imag} */,
  {32'hc4b3788e, 32'h00000000} /* (25, 20, 15) {real, imag} */,
  {32'hc43dd8d6, 32'h00000000} /* (25, 20, 14) {real, imag} */,
  {32'hc2f5635c, 32'h00000000} /* (25, 20, 13) {real, imag} */,
  {32'hc2d7199c, 32'h00000000} /* (25, 20, 12) {real, imag} */,
  {32'hc462d8af, 32'h00000000} /* (25, 20, 11) {real, imag} */,
  {32'hc2e7c7a4, 32'h00000000} /* (25, 20, 10) {real, imag} */,
  {32'hc3cdd98d, 32'h00000000} /* (25, 20, 9) {real, imag} */,
  {32'h43f10a0a, 32'h00000000} /* (25, 20, 8) {real, imag} */,
  {32'h44114bd0, 32'h00000000} /* (25, 20, 7) {real, imag} */,
  {32'h44e13984, 32'h00000000} /* (25, 20, 6) {real, imag} */,
  {32'h43854f2a, 32'h00000000} /* (25, 20, 5) {real, imag} */,
  {32'h43d4b4d8, 32'h00000000} /* (25, 20, 4) {real, imag} */,
  {32'h43e42d10, 32'h00000000} /* (25, 20, 3) {real, imag} */,
  {32'h4306e1b6, 32'h00000000} /* (25, 20, 2) {real, imag} */,
  {32'h449d5514, 32'h00000000} /* (25, 20, 1) {real, imag} */,
  {32'h447cc1f1, 32'h00000000} /* (25, 20, 0) {real, imag} */,
  {32'h44ff42c8, 32'h00000000} /* (25, 19, 31) {real, imag} */,
  {32'h44fcb80e, 32'h00000000} /* (25, 19, 30) {real, imag} */,
  {32'h4505615e, 32'h00000000} /* (25, 19, 29) {real, imag} */,
  {32'h44fe480c, 32'h00000000} /* (25, 19, 28) {real, imag} */,
  {32'h452bb9f2, 32'h00000000} /* (25, 19, 27) {real, imag} */,
  {32'h450cdd50, 32'h00000000} /* (25, 19, 26) {real, imag} */,
  {32'h44d19120, 32'h00000000} /* (25, 19, 25) {real, imag} */,
  {32'h44a03fba, 32'h00000000} /* (25, 19, 24) {real, imag} */,
  {32'h44ec51dd, 32'h00000000} /* (25, 19, 23) {real, imag} */,
  {32'h45072f9a, 32'h00000000} /* (25, 19, 22) {real, imag} */,
  {32'h44449e5b, 32'h00000000} /* (25, 19, 21) {real, imag} */,
  {32'hc48b77d0, 32'h00000000} /* (25, 19, 20) {real, imag} */,
  {32'hc4827b34, 32'h00000000} /* (25, 19, 19) {real, imag} */,
  {32'hc4c10deb, 32'h00000000} /* (25, 19, 18) {real, imag} */,
  {32'hc4c8a816, 32'h00000000} /* (25, 19, 17) {real, imag} */,
  {32'hc4bce916, 32'h00000000} /* (25, 19, 16) {real, imag} */,
  {32'hc47ab1af, 32'h00000000} /* (25, 19, 15) {real, imag} */,
  {32'hc4a250bc, 32'h00000000} /* (25, 19, 14) {real, imag} */,
  {32'hc47978d6, 32'h00000000} /* (25, 19, 13) {real, imag} */,
  {32'hc4dde884, 32'h00000000} /* (25, 19, 12) {real, imag} */,
  {32'hc48195b5, 32'h00000000} /* (25, 19, 11) {real, imag} */,
  {32'h449e9a0a, 32'h00000000} /* (25, 19, 10) {real, imag} */,
  {32'h44c2dbe0, 32'h00000000} /* (25, 19, 9) {real, imag} */,
  {32'h44aaa7e6, 32'h00000000} /* (25, 19, 8) {real, imag} */,
  {32'h4515a49f, 32'h00000000} /* (25, 19, 7) {real, imag} */,
  {32'h44bb28f1, 32'h00000000} /* (25, 19, 6) {real, imag} */,
  {32'h44932336, 32'h00000000} /* (25, 19, 5) {real, imag} */,
  {32'h44bd0e08, 32'h00000000} /* (25, 19, 4) {real, imag} */,
  {32'h4496aa16, 32'h00000000} /* (25, 19, 3) {real, imag} */,
  {32'h448efdbd, 32'h00000000} /* (25, 19, 2) {real, imag} */,
  {32'h44d33938, 32'h00000000} /* (25, 19, 1) {real, imag} */,
  {32'h44dd1fea, 32'h00000000} /* (25, 19, 0) {real, imag} */,
  {32'h454c1698, 32'h00000000} /* (25, 18, 31) {real, imag} */,
  {32'h4540b322, 32'h00000000} /* (25, 18, 30) {real, imag} */,
  {32'h4500e725, 32'h00000000} /* (25, 18, 29) {real, imag} */,
  {32'h450bbf6b, 32'h00000000} /* (25, 18, 28) {real, imag} */,
  {32'h454f0f7e, 32'h00000000} /* (25, 18, 27) {real, imag} */,
  {32'h453292be, 32'h00000000} /* (25, 18, 26) {real, imag} */,
  {32'h4516049a, 32'h00000000} /* (25, 18, 25) {real, imag} */,
  {32'h452971f8, 32'h00000000} /* (25, 18, 24) {real, imag} */,
  {32'h44f98ae4, 32'h00000000} /* (25, 18, 23) {real, imag} */,
  {32'h44ad6070, 32'h00000000} /* (25, 18, 22) {real, imag} */,
  {32'hc212ab80, 32'h00000000} /* (25, 18, 21) {real, imag} */,
  {32'hc472bf30, 32'h00000000} /* (25, 18, 20) {real, imag} */,
  {32'hc4c64508, 32'h00000000} /* (25, 18, 19) {real, imag} */,
  {32'hc51350aa, 32'h00000000} /* (25, 18, 18) {real, imag} */,
  {32'hc52582c4, 32'h00000000} /* (25, 18, 17) {real, imag} */,
  {32'hc4eb7d76, 32'h00000000} /* (25, 18, 16) {real, imag} */,
  {32'hc50a3f28, 32'h00000000} /* (25, 18, 15) {real, imag} */,
  {32'hc4e687f5, 32'h00000000} /* (25, 18, 14) {real, imag} */,
  {32'hc504fa15, 32'h00000000} /* (25, 18, 13) {real, imag} */,
  {32'hc4c4e399, 32'h00000000} /* (25, 18, 12) {real, imag} */,
  {32'hc3fe5d30, 32'h00000000} /* (25, 18, 11) {real, imag} */,
  {32'hc290b630, 32'h00000000} /* (25, 18, 10) {real, imag} */,
  {32'h44f1989b, 32'h00000000} /* (25, 18, 9) {real, imag} */,
  {32'h450f3566, 32'h00000000} /* (25, 18, 8) {real, imag} */,
  {32'h4528ba28, 32'h00000000} /* (25, 18, 7) {real, imag} */,
  {32'h453f59c4, 32'h00000000} /* (25, 18, 6) {real, imag} */,
  {32'h4513ee0a, 32'h00000000} /* (25, 18, 5) {real, imag} */,
  {32'h45023e28, 32'h00000000} /* (25, 18, 4) {real, imag} */,
  {32'h44d64f5a, 32'h00000000} /* (25, 18, 3) {real, imag} */,
  {32'h455b8826, 32'h00000000} /* (25, 18, 2) {real, imag} */,
  {32'h45237da8, 32'h00000000} /* (25, 18, 1) {real, imag} */,
  {32'h450fe98f, 32'h00000000} /* (25, 18, 0) {real, imag} */,
  {32'h453e475f, 32'h00000000} /* (25, 17, 31) {real, imag} */,
  {32'h45409cbe, 32'h00000000} /* (25, 17, 30) {real, imag} */,
  {32'h455e74d0, 32'h00000000} /* (25, 17, 29) {real, imag} */,
  {32'h4559bc9a, 32'h00000000} /* (25, 17, 28) {real, imag} */,
  {32'h457f54b8, 32'h00000000} /* (25, 17, 27) {real, imag} */,
  {32'h4557ecb2, 32'h00000000} /* (25, 17, 26) {real, imag} */,
  {32'h4554aaaf, 32'h00000000} /* (25, 17, 25) {real, imag} */,
  {32'h456eaa2e, 32'h00000000} /* (25, 17, 24) {real, imag} */,
  {32'h4534c159, 32'h00000000} /* (25, 17, 23) {real, imag} */,
  {32'h44dbacae, 32'h00000000} /* (25, 17, 22) {real, imag} */,
  {32'h441385a6, 32'h00000000} /* (25, 17, 21) {real, imag} */,
  {32'hc4a1dfea, 32'h00000000} /* (25, 17, 20) {real, imag} */,
  {32'hc4e7a328, 32'h00000000} /* (25, 17, 19) {real, imag} */,
  {32'hc515b443, 32'h00000000} /* (25, 17, 18) {real, imag} */,
  {32'hc534db80, 32'h00000000} /* (25, 17, 17) {real, imag} */,
  {32'hc5293923, 32'h00000000} /* (25, 17, 16) {real, imag} */,
  {32'hc51f4dd7, 32'h00000000} /* (25, 17, 15) {real, imag} */,
  {32'hc53c0c0a, 32'h00000000} /* (25, 17, 14) {real, imag} */,
  {32'hc5300008, 32'h00000000} /* (25, 17, 13) {real, imag} */,
  {32'hc4e00e7c, 32'h00000000} /* (25, 17, 12) {real, imag} */,
  {32'hc4917c0c, 32'h00000000} /* (25, 17, 11) {real, imag} */,
  {32'h442a16ae, 32'h00000000} /* (25, 17, 10) {real, imag} */,
  {32'h44de58fa, 32'h00000000} /* (25, 17, 9) {real, imag} */,
  {32'h453eae8c, 32'h00000000} /* (25, 17, 8) {real, imag} */,
  {32'h4585f0ca, 32'h00000000} /* (25, 17, 7) {real, imag} */,
  {32'h455525b5, 32'h00000000} /* (25, 17, 6) {real, imag} */,
  {32'h45431fee, 32'h00000000} /* (25, 17, 5) {real, imag} */,
  {32'h451d89be, 32'h00000000} /* (25, 17, 4) {real, imag} */,
  {32'h45419dac, 32'h00000000} /* (25, 17, 3) {real, imag} */,
  {32'h45514899, 32'h00000000} /* (25, 17, 2) {real, imag} */,
  {32'h452846c8, 32'h00000000} /* (25, 17, 1) {real, imag} */,
  {32'h453c98d1, 32'h00000000} /* (25, 17, 0) {real, imag} */,
  {32'h455c4612, 32'h00000000} /* (25, 16, 31) {real, imag} */,
  {32'h456f40b4, 32'h00000000} /* (25, 16, 30) {real, imag} */,
  {32'h4564aff2, 32'h00000000} /* (25, 16, 29) {real, imag} */,
  {32'h458c3503, 32'h00000000} /* (25, 16, 28) {real, imag} */,
  {32'h4534ff3d, 32'h00000000} /* (25, 16, 27) {real, imag} */,
  {32'h453a4576, 32'h00000000} /* (25, 16, 26) {real, imag} */,
  {32'h456c73e0, 32'h00000000} /* (25, 16, 25) {real, imag} */,
  {32'h451e4830, 32'h00000000} /* (25, 16, 24) {real, imag} */,
  {32'h4525cac0, 32'h00000000} /* (25, 16, 23) {real, imag} */,
  {32'h44cd497c, 32'h00000000} /* (25, 16, 22) {real, imag} */,
  {32'hc23f9e80, 32'h00000000} /* (25, 16, 21) {real, imag} */,
  {32'hc495d399, 32'h00000000} /* (25, 16, 20) {real, imag} */,
  {32'hc5067e46, 32'h00000000} /* (25, 16, 19) {real, imag} */,
  {32'hc51dafe4, 32'h00000000} /* (25, 16, 18) {real, imag} */,
  {32'hc52ca6e0, 32'h00000000} /* (25, 16, 17) {real, imag} */,
  {32'hc557a3fc, 32'h00000000} /* (25, 16, 16) {real, imag} */,
  {32'hc529c7ee, 32'h00000000} /* (25, 16, 15) {real, imag} */,
  {32'hc54aac94, 32'h00000000} /* (25, 16, 14) {real, imag} */,
  {32'hc53f08fa, 32'h00000000} /* (25, 16, 13) {real, imag} */,
  {32'hc539a0fc, 32'h00000000} /* (25, 16, 12) {real, imag} */,
  {32'hc4f3a2f2, 32'h00000000} /* (25, 16, 11) {real, imag} */,
  {32'h43fd374c, 32'h00000000} /* (25, 16, 10) {real, imag} */,
  {32'h44a0d817, 32'h00000000} /* (25, 16, 9) {real, imag} */,
  {32'h4528a22c, 32'h00000000} /* (25, 16, 8) {real, imag} */,
  {32'h4583284c, 32'h00000000} /* (25, 16, 7) {real, imag} */,
  {32'h45c60925, 32'h00000000} /* (25, 16, 6) {real, imag} */,
  {32'h45649e0a, 32'h00000000} /* (25, 16, 5) {real, imag} */,
  {32'h4581a01c, 32'h00000000} /* (25, 16, 4) {real, imag} */,
  {32'h458ce651, 32'h00000000} /* (25, 16, 3) {real, imag} */,
  {32'h457620e2, 32'h00000000} /* (25, 16, 2) {real, imag} */,
  {32'h45605480, 32'h00000000} /* (25, 16, 1) {real, imag} */,
  {32'h45787474, 32'h00000000} /* (25, 16, 0) {real, imag} */,
  {32'h4562f148, 32'h00000000} /* (25, 15, 31) {real, imag} */,
  {32'h4570d850, 32'h00000000} /* (25, 15, 30) {real, imag} */,
  {32'h456795b6, 32'h00000000} /* (25, 15, 29) {real, imag} */,
  {32'h45827a28, 32'h00000000} /* (25, 15, 28) {real, imag} */,
  {32'h453ea7d6, 32'h00000000} /* (25, 15, 27) {real, imag} */,
  {32'h4522b6e5, 32'h00000000} /* (25, 15, 26) {real, imag} */,
  {32'h4507b92a, 32'h00000000} /* (25, 15, 25) {real, imag} */,
  {32'h45121086, 32'h00000000} /* (25, 15, 24) {real, imag} */,
  {32'h452f55f8, 32'h00000000} /* (25, 15, 23) {real, imag} */,
  {32'h44bd25e2, 32'h00000000} /* (25, 15, 22) {real, imag} */,
  {32'h4351c340, 32'h00000000} /* (25, 15, 21) {real, imag} */,
  {32'hc4adc80e, 32'h00000000} /* (25, 15, 20) {real, imag} */,
  {32'hc5281788, 32'h00000000} /* (25, 15, 19) {real, imag} */,
  {32'hc52a0fc4, 32'h00000000} /* (25, 15, 18) {real, imag} */,
  {32'hc5695707, 32'h00000000} /* (25, 15, 17) {real, imag} */,
  {32'hc565825c, 32'h00000000} /* (25, 15, 16) {real, imag} */,
  {32'hc55e6c14, 32'h00000000} /* (25, 15, 15) {real, imag} */,
  {32'hc55a0206, 32'h00000000} /* (25, 15, 14) {real, imag} */,
  {32'hc51e44ce, 32'h00000000} /* (25, 15, 13) {real, imag} */,
  {32'hc5012cd3, 32'h00000000} /* (25, 15, 12) {real, imag} */,
  {32'hc49050f3, 32'h00000000} /* (25, 15, 11) {real, imag} */,
  {32'h43eebb90, 32'h00000000} /* (25, 15, 10) {real, imag} */,
  {32'h44f11994, 32'h00000000} /* (25, 15, 9) {real, imag} */,
  {32'h451babd6, 32'h00000000} /* (25, 15, 8) {real, imag} */,
  {32'h454683ac, 32'h00000000} /* (25, 15, 7) {real, imag} */,
  {32'h455d1ddf, 32'h00000000} /* (25, 15, 6) {real, imag} */,
  {32'h457214b8, 32'h00000000} /* (25, 15, 5) {real, imag} */,
  {32'h458e545c, 32'h00000000} /* (25, 15, 4) {real, imag} */,
  {32'h4574c0ce, 32'h00000000} /* (25, 15, 3) {real, imag} */,
  {32'h455e6fe0, 32'h00000000} /* (25, 15, 2) {real, imag} */,
  {32'h454e44e1, 32'h00000000} /* (25, 15, 1) {real, imag} */,
  {32'h4554b0d6, 32'h00000000} /* (25, 15, 0) {real, imag} */,
  {32'h45406f8c, 32'h00000000} /* (25, 14, 31) {real, imag} */,
  {32'h4544113f, 32'h00000000} /* (25, 14, 30) {real, imag} */,
  {32'h455c65c1, 32'h00000000} /* (25, 14, 29) {real, imag} */,
  {32'h453e8160, 32'h00000000} /* (25, 14, 28) {real, imag} */,
  {32'h45611bf7, 32'h00000000} /* (25, 14, 27) {real, imag} */,
  {32'h45374de6, 32'h00000000} /* (25, 14, 26) {real, imag} */,
  {32'h45111ec5, 32'h00000000} /* (25, 14, 25) {real, imag} */,
  {32'h4509e91b, 32'h00000000} /* (25, 14, 24) {real, imag} */,
  {32'h4505b44e, 32'h00000000} /* (25, 14, 23) {real, imag} */,
  {32'h446fa596, 32'h00000000} /* (25, 14, 22) {real, imag} */,
  {32'h42d3f890, 32'h00000000} /* (25, 14, 21) {real, imag} */,
  {32'hc49b5281, 32'h00000000} /* (25, 14, 20) {real, imag} */,
  {32'hc52c475e, 32'h00000000} /* (25, 14, 19) {real, imag} */,
  {32'hc5540e32, 32'h00000000} /* (25, 14, 18) {real, imag} */,
  {32'hc55607be, 32'h00000000} /* (25, 14, 17) {real, imag} */,
  {32'hc584ceb2, 32'h00000000} /* (25, 14, 16) {real, imag} */,
  {32'hc55bc032, 32'h00000000} /* (25, 14, 15) {real, imag} */,
  {32'hc5426557, 32'h00000000} /* (25, 14, 14) {real, imag} */,
  {32'hc551f10f, 32'h00000000} /* (25, 14, 13) {real, imag} */,
  {32'hc5040b2e, 32'h00000000} /* (25, 14, 12) {real, imag} */,
  {32'hc49a258e, 32'h00000000} /* (25, 14, 11) {real, imag} */,
  {32'h43c71d34, 32'h00000000} /* (25, 14, 10) {real, imag} */,
  {32'h44db559e, 32'h00000000} /* (25, 14, 9) {real, imag} */,
  {32'h4523987b, 32'h00000000} /* (25, 14, 8) {real, imag} */,
  {32'h4554795a, 32'h00000000} /* (25, 14, 7) {real, imag} */,
  {32'h454cf57a, 32'h00000000} /* (25, 14, 6) {real, imag} */,
  {32'h45725a66, 32'h00000000} /* (25, 14, 5) {real, imag} */,
  {32'h45720bd8, 32'h00000000} /* (25, 14, 4) {real, imag} */,
  {32'h4558fece, 32'h00000000} /* (25, 14, 3) {real, imag} */,
  {32'h453de54a, 32'h00000000} /* (25, 14, 2) {real, imag} */,
  {32'h4558de8e, 32'h00000000} /* (25, 14, 1) {real, imag} */,
  {32'h452827da, 32'h00000000} /* (25, 14, 0) {real, imag} */,
  {32'h4518b4e5, 32'h00000000} /* (25, 13, 31) {real, imag} */,
  {32'h454ff4c2, 32'h00000000} /* (25, 13, 30) {real, imag} */,
  {32'h45319b63, 32'h00000000} /* (25, 13, 29) {real, imag} */,
  {32'h455ef79a, 32'h00000000} /* (25, 13, 28) {real, imag} */,
  {32'h455bd9a1, 32'h00000000} /* (25, 13, 27) {real, imag} */,
  {32'h45133e6a, 32'h00000000} /* (25, 13, 26) {real, imag} */,
  {32'h452a608b, 32'h00000000} /* (25, 13, 25) {real, imag} */,
  {32'h45214e90, 32'h00000000} /* (25, 13, 24) {real, imag} */,
  {32'h4514b354, 32'h00000000} /* (25, 13, 23) {real, imag} */,
  {32'h44df0036, 32'h00000000} /* (25, 13, 22) {real, imag} */,
  {32'h413d6e00, 32'h00000000} /* (25, 13, 21) {real, imag} */,
  {32'hc4d7b4cc, 32'h00000000} /* (25, 13, 20) {real, imag} */,
  {32'hc5055204, 32'h00000000} /* (25, 13, 19) {real, imag} */,
  {32'hc510efb7, 32'h00000000} /* (25, 13, 18) {real, imag} */,
  {32'hc5547923, 32'h00000000} /* (25, 13, 17) {real, imag} */,
  {32'hc58d042c, 32'h00000000} /* (25, 13, 16) {real, imag} */,
  {32'hc54fb365, 32'h00000000} /* (25, 13, 15) {real, imag} */,
  {32'hc528c968, 32'h00000000} /* (25, 13, 14) {real, imag} */,
  {32'hc5085ffd, 32'h00000000} /* (25, 13, 13) {real, imag} */,
  {32'hc4fd1dc8, 32'h00000000} /* (25, 13, 12) {real, imag} */,
  {32'hc48758fe, 32'h00000000} /* (25, 13, 11) {real, imag} */,
  {32'h44a36d0b, 32'h00000000} /* (25, 13, 10) {real, imag} */,
  {32'h44f9e0f2, 32'h00000000} /* (25, 13, 9) {real, imag} */,
  {32'h451c96b4, 32'h00000000} /* (25, 13, 8) {real, imag} */,
  {32'h455dddf2, 32'h00000000} /* (25, 13, 7) {real, imag} */,
  {32'h456ccc49, 32'h00000000} /* (25, 13, 6) {real, imag} */,
  {32'h4581a362, 32'h00000000} /* (25, 13, 5) {real, imag} */,
  {32'h458d22ad, 32'h00000000} /* (25, 13, 4) {real, imag} */,
  {32'h454f6dd4, 32'h00000000} /* (25, 13, 3) {real, imag} */,
  {32'h45318273, 32'h00000000} /* (25, 13, 2) {real, imag} */,
  {32'h4522d9af, 32'h00000000} /* (25, 13, 1) {real, imag} */,
  {32'h4522cfce, 32'h00000000} /* (25, 13, 0) {real, imag} */,
  {32'h4511367a, 32'h00000000} /* (25, 12, 31) {real, imag} */,
  {32'h453dd489, 32'h00000000} /* (25, 12, 30) {real, imag} */,
  {32'h44e41045, 32'h00000000} /* (25, 12, 29) {real, imag} */,
  {32'h451c3f3c, 32'h00000000} /* (25, 12, 28) {real, imag} */,
  {32'h450a225e, 32'h00000000} /* (25, 12, 27) {real, imag} */,
  {32'h44ba061a, 32'h00000000} /* (25, 12, 26) {real, imag} */,
  {32'h451437a3, 32'h00000000} /* (25, 12, 25) {real, imag} */,
  {32'h450ebb1d, 32'h00000000} /* (25, 12, 24) {real, imag} */,
  {32'h44d10009, 32'h00000000} /* (25, 12, 23) {real, imag} */,
  {32'h444f4ff8, 32'h00000000} /* (25, 12, 22) {real, imag} */,
  {32'h42f38f10, 32'h00000000} /* (25, 12, 21) {real, imag} */,
  {32'hc507b708, 32'h00000000} /* (25, 12, 20) {real, imag} */,
  {32'hc53e4cb2, 32'h00000000} /* (25, 12, 19) {real, imag} */,
  {32'hc558d718, 32'h00000000} /* (25, 12, 18) {real, imag} */,
  {32'hc5395428, 32'h00000000} /* (25, 12, 17) {real, imag} */,
  {32'hc53b91d8, 32'h00000000} /* (25, 12, 16) {real, imag} */,
  {32'hc53470c8, 32'h00000000} /* (25, 12, 15) {real, imag} */,
  {32'hc50f7335, 32'h00000000} /* (25, 12, 14) {real, imag} */,
  {32'hc4a39baf, 32'h00000000} /* (25, 12, 13) {real, imag} */,
  {32'hc4c12118, 32'h00000000} /* (25, 12, 12) {real, imag} */,
  {32'hc4b5aaed, 32'h00000000} /* (25, 12, 11) {real, imag} */,
  {32'h4510d3b3, 32'h00000000} /* (25, 12, 10) {real, imag} */,
  {32'h4516fa37, 32'h00000000} /* (25, 12, 9) {real, imag} */,
  {32'h450fadb3, 32'h00000000} /* (25, 12, 8) {real, imag} */,
  {32'h4546182e, 32'h00000000} /* (25, 12, 7) {real, imag} */,
  {32'h4560eeda, 32'h00000000} /* (25, 12, 6) {real, imag} */,
  {32'h454b8574, 32'h00000000} /* (25, 12, 5) {real, imag} */,
  {32'h452485ce, 32'h00000000} /* (25, 12, 4) {real, imag} */,
  {32'h44f55653, 32'h00000000} /* (25, 12, 3) {real, imag} */,
  {32'h451d2570, 32'h00000000} /* (25, 12, 2) {real, imag} */,
  {32'h4510d928, 32'h00000000} /* (25, 12, 1) {real, imag} */,
  {32'h44afe044, 32'h00000000} /* (25, 12, 0) {real, imag} */,
  {32'h44388350, 32'h00000000} /* (25, 11, 31) {real, imag} */,
  {32'h448e0f5a, 32'h00000000} /* (25, 11, 30) {real, imag} */,
  {32'h44282fe9, 32'h00000000} /* (25, 11, 29) {real, imag} */,
  {32'h4469fa43, 32'h00000000} /* (25, 11, 28) {real, imag} */,
  {32'h4402ed71, 32'h00000000} /* (25, 11, 27) {real, imag} */,
  {32'h43e56fb2, 32'h00000000} /* (25, 11, 26) {real, imag} */,
  {32'h446cd4b0, 32'h00000000} /* (25, 11, 25) {real, imag} */,
  {32'h44a93f04, 32'h00000000} /* (25, 11, 24) {real, imag} */,
  {32'h448478cc, 32'h00000000} /* (25, 11, 23) {real, imag} */,
  {32'h447fc82b, 32'h00000000} /* (25, 11, 22) {real, imag} */,
  {32'hc3a99574, 32'h00000000} /* (25, 11, 21) {real, imag} */,
  {32'hc4d257bd, 32'h00000000} /* (25, 11, 20) {real, imag} */,
  {32'hc4e64abc, 32'h00000000} /* (25, 11, 19) {real, imag} */,
  {32'hc5400968, 32'h00000000} /* (25, 11, 18) {real, imag} */,
  {32'hc53b8bbb, 32'h00000000} /* (25, 11, 17) {real, imag} */,
  {32'hc48991e6, 32'h00000000} /* (25, 11, 16) {real, imag} */,
  {32'hc48520de, 32'h00000000} /* (25, 11, 15) {real, imag} */,
  {32'hc46a45f4, 32'h00000000} /* (25, 11, 14) {real, imag} */,
  {32'hc45cb119, 32'h00000000} /* (25, 11, 13) {real, imag} */,
  {32'hc4741a19, 32'h00000000} /* (25, 11, 12) {real, imag} */,
  {32'hc4763ad7, 32'h00000000} /* (25, 11, 11) {real, imag} */,
  {32'h4428613b, 32'h00000000} /* (25, 11, 10) {real, imag} */,
  {32'h44f34ffc, 32'h00000000} /* (25, 11, 9) {real, imag} */,
  {32'h453aaa2e, 32'h00000000} /* (25, 11, 8) {real, imag} */,
  {32'h45636f72, 32'h00000000} /* (25, 11, 7) {real, imag} */,
  {32'h45227553, 32'h00000000} /* (25, 11, 6) {real, imag} */,
  {32'h44eed7d7, 32'h00000000} /* (25, 11, 5) {real, imag} */,
  {32'h44a44ac7, 32'h00000000} /* (25, 11, 4) {real, imag} */,
  {32'h44748605, 32'h00000000} /* (25, 11, 3) {real, imag} */,
  {32'h445fc648, 32'h00000000} /* (25, 11, 2) {real, imag} */,
  {32'h44c58616, 32'h00000000} /* (25, 11, 1) {real, imag} */,
  {32'h448df51a, 32'h00000000} /* (25, 11, 0) {real, imag} */,
  {32'hc4694b84, 32'h00000000} /* (25, 10, 31) {real, imag} */,
  {32'hc4ac0aac, 32'h00000000} /* (25, 10, 30) {real, imag} */,
  {32'hc5228902, 32'h00000000} /* (25, 10, 29) {real, imag} */,
  {32'hc503d949, 32'h00000000} /* (25, 10, 28) {real, imag} */,
  {32'hc5057cc2, 32'h00000000} /* (25, 10, 27) {real, imag} */,
  {32'hc50f1d16, 32'h00000000} /* (25, 10, 26) {real, imag} */,
  {32'hc519f066, 32'h00000000} /* (25, 10, 25) {real, imag} */,
  {32'hc478398c, 32'h00000000} /* (25, 10, 24) {real, imag} */,
  {32'hc4a4c295, 32'h00000000} /* (25, 10, 23) {real, imag} */,
  {32'hc49442ae, 32'h00000000} /* (25, 10, 22) {real, imag} */,
  {32'hc4aadaee, 32'h00000000} /* (25, 10, 21) {real, imag} */,
  {32'hc446e537, 32'h00000000} /* (25, 10, 20) {real, imag} */,
  {32'hc2313e90, 32'h00000000} /* (25, 10, 19) {real, imag} */,
  {32'hc3d42fc2, 32'h00000000} /* (25, 10, 18) {real, imag} */,
  {32'h4485315f, 32'h00000000} /* (25, 10, 17) {real, imag} */,
  {32'h44195d6e, 32'h00000000} /* (25, 10, 16) {real, imag} */,
  {32'h44471f68, 32'h00000000} /* (25, 10, 15) {real, imag} */,
  {32'h440c04c9, 32'h00000000} /* (25, 10, 14) {real, imag} */,
  {32'h42822380, 32'h00000000} /* (25, 10, 13) {real, imag} */,
  {32'h43840a38, 32'h00000000} /* (25, 10, 12) {real, imag} */,
  {32'h44c2c058, 32'h00000000} /* (25, 10, 11) {real, imag} */,
  {32'h4469a000, 32'h00000000} /* (25, 10, 10) {real, imag} */,
  {32'h43e3bc3c, 32'h00000000} /* (25, 10, 9) {real, imag} */,
  {32'h43764c18, 32'h00000000} /* (25, 10, 8) {real, imag} */,
  {32'h4500163d, 32'h00000000} /* (25, 10, 7) {real, imag} */,
  {32'h42a4d0a8, 32'h00000000} /* (25, 10, 6) {real, imag} */,
  {32'hc329d694, 32'h00000000} /* (25, 10, 5) {real, imag} */,
  {32'hc45471c1, 32'h00000000} /* (25, 10, 4) {real, imag} */,
  {32'hc4b31ec0, 32'h00000000} /* (25, 10, 3) {real, imag} */,
  {32'hc4874178, 32'h00000000} /* (25, 10, 2) {real, imag} */,
  {32'hc518616c, 32'h00000000} /* (25, 10, 1) {real, imag} */,
  {32'hc4db1d8b, 32'h00000000} /* (25, 10, 0) {real, imag} */,
  {32'hc534a540, 32'h00000000} /* (25, 9, 31) {real, imag} */,
  {32'hc55608f6, 32'h00000000} /* (25, 9, 30) {real, imag} */,
  {32'hc5612081, 32'h00000000} /* (25, 9, 29) {real, imag} */,
  {32'hc56c3fae, 32'h00000000} /* (25, 9, 28) {real, imag} */,
  {32'hc5907b9b, 32'h00000000} /* (25, 9, 27) {real, imag} */,
  {32'hc5860e86, 32'h00000000} /* (25, 9, 26) {real, imag} */,
  {32'hc552def1, 32'h00000000} /* (25, 9, 25) {real, imag} */,
  {32'hc553a1a2, 32'h00000000} /* (25, 9, 24) {real, imag} */,
  {32'hc513ecf2, 32'h00000000} /* (25, 9, 23) {real, imag} */,
  {32'hc51bc077, 32'h00000000} /* (25, 9, 22) {real, imag} */,
  {32'hc507083c, 32'h00000000} /* (25, 9, 21) {real, imag} */,
  {32'hc38575b0, 32'h00000000} /* (25, 9, 20) {real, imag} */,
  {32'h42f84ce0, 32'h00000000} /* (25, 9, 19) {real, imag} */,
  {32'h4445557a, 32'h00000000} /* (25, 9, 18) {real, imag} */,
  {32'h44788aa8, 32'h00000000} /* (25, 9, 17) {real, imag} */,
  {32'h4493c130, 32'h00000000} /* (25, 9, 16) {real, imag} */,
  {32'h44abcd93, 32'h00000000} /* (25, 9, 15) {real, imag} */,
  {32'h450e5dee, 32'h00000000} /* (25, 9, 14) {real, imag} */,
  {32'h44c70562, 32'h00000000} /* (25, 9, 13) {real, imag} */,
  {32'h44d21fd5, 32'h00000000} /* (25, 9, 12) {real, imag} */,
  {32'h44c191c4, 32'h00000000} /* (25, 9, 11) {real, imag} */,
  {32'h44163d6a, 32'h00000000} /* (25, 9, 10) {real, imag} */,
  {32'hc3112350, 32'h00000000} /* (25, 9, 9) {real, imag} */,
  {32'hc4776dc8, 32'h00000000} /* (25, 9, 8) {real, imag} */,
  {32'hc440a29c, 32'h00000000} /* (25, 9, 7) {real, imag} */,
  {32'hc47561f5, 32'h00000000} /* (25, 9, 6) {real, imag} */,
  {32'hc5037a3c, 32'h00000000} /* (25, 9, 5) {real, imag} */,
  {32'hc51ab479, 32'h00000000} /* (25, 9, 4) {real, imag} */,
  {32'hc52d7b9b, 32'h00000000} /* (25, 9, 3) {real, imag} */,
  {32'hc53c473e, 32'h00000000} /* (25, 9, 2) {real, imag} */,
  {32'hc5657924, 32'h00000000} /* (25, 9, 1) {real, imag} */,
  {32'hc545b346, 32'h00000000} /* (25, 9, 0) {real, imag} */,
  {32'hc567c95a, 32'h00000000} /* (25, 8, 31) {real, imag} */,
  {32'hc5772554, 32'h00000000} /* (25, 8, 30) {real, imag} */,
  {32'hc5ad2e15, 32'h00000000} /* (25, 8, 29) {real, imag} */,
  {32'hc5a82e1e, 32'h00000000} /* (25, 8, 28) {real, imag} */,
  {32'hc5936b5f, 32'h00000000} /* (25, 8, 27) {real, imag} */,
  {32'hc599901c, 32'h00000000} /* (25, 8, 26) {real, imag} */,
  {32'hc59f0e56, 32'h00000000} /* (25, 8, 25) {real, imag} */,
  {32'hc58bbf28, 32'h00000000} /* (25, 8, 24) {real, imag} */,
  {32'hc56447d6, 32'h00000000} /* (25, 8, 23) {real, imag} */,
  {32'hc554a7ac, 32'h00000000} /* (25, 8, 22) {real, imag} */,
  {32'hc5120406, 32'h00000000} /* (25, 8, 21) {real, imag} */,
  {32'hc3fd1048, 32'h00000000} /* (25, 8, 20) {real, imag} */,
  {32'h43a0d51c, 32'h00000000} /* (25, 8, 19) {real, imag} */,
  {32'h4468dd30, 32'h00000000} /* (25, 8, 18) {real, imag} */,
  {32'h448d3c7f, 32'h00000000} /* (25, 8, 17) {real, imag} */,
  {32'h44df4bea, 32'h00000000} /* (25, 8, 16) {real, imag} */,
  {32'h4510951a, 32'h00000000} /* (25, 8, 15) {real, imag} */,
  {32'h4515f98c, 32'h00000000} /* (25, 8, 14) {real, imag} */,
  {32'h4515308c, 32'h00000000} /* (25, 8, 13) {real, imag} */,
  {32'h44e9f0f7, 32'h00000000} /* (25, 8, 12) {real, imag} */,
  {32'h44dfddd0, 32'h00000000} /* (25, 8, 11) {real, imag} */,
  {32'h43c55908, 32'h00000000} /* (25, 8, 10) {real, imag} */,
  {32'hc3ac6be8, 32'h00000000} /* (25, 8, 9) {real, imag} */,
  {32'hc452c46a, 32'h00000000} /* (25, 8, 8) {real, imag} */,
  {32'hc4dcf911, 32'h00000000} /* (25, 8, 7) {real, imag} */,
  {32'hc51e0966, 32'h00000000} /* (25, 8, 6) {real, imag} */,
  {32'hc53d4f9e, 32'h00000000} /* (25, 8, 5) {real, imag} */,
  {32'hc5268d3a, 32'h00000000} /* (25, 8, 4) {real, imag} */,
  {32'hc5407988, 32'h00000000} /* (25, 8, 3) {real, imag} */,
  {32'hc56b3316, 32'h00000000} /* (25, 8, 2) {real, imag} */,
  {32'hc592b608, 32'h00000000} /* (25, 8, 1) {real, imag} */,
  {32'hc5933106, 32'h00000000} /* (25, 8, 0) {real, imag} */,
  {32'hc5867ffb, 32'h00000000} /* (25, 7, 31) {real, imag} */,
  {32'hc5ae0972, 32'h00000000} /* (25, 7, 30) {real, imag} */,
  {32'hc5e06eb2, 32'h00000000} /* (25, 7, 29) {real, imag} */,
  {32'hc5e87bc6, 32'h00000000} /* (25, 7, 28) {real, imag} */,
  {32'hc5bee1e6, 32'h00000000} /* (25, 7, 27) {real, imag} */,
  {32'hc5a439ba, 32'h00000000} /* (25, 7, 26) {real, imag} */,
  {32'hc5b6d7a3, 32'h00000000} /* (25, 7, 25) {real, imag} */,
  {32'hc5a05221, 32'h00000000} /* (25, 7, 24) {real, imag} */,
  {32'hc5a24ee6, 32'h00000000} /* (25, 7, 23) {real, imag} */,
  {32'hc587daf6, 32'h00000000} /* (25, 7, 22) {real, imag} */,
  {32'hc52c712f, 32'h00000000} /* (25, 7, 21) {real, imag} */,
  {32'hc3c556b4, 32'h00000000} /* (25, 7, 20) {real, imag} */,
  {32'h424c2500, 32'h00000000} /* (25, 7, 19) {real, imag} */,
  {32'h43c6cf00, 32'h00000000} /* (25, 7, 18) {real, imag} */,
  {32'h448826de, 32'h00000000} /* (25, 7, 17) {real, imag} */,
  {32'h449a0402, 32'h00000000} /* (25, 7, 16) {real, imag} */,
  {32'h44f85987, 32'h00000000} /* (25, 7, 15) {real, imag} */,
  {32'h450b3713, 32'h00000000} /* (25, 7, 14) {real, imag} */,
  {32'h4518738d, 32'h00000000} /* (25, 7, 13) {real, imag} */,
  {32'h44e61db2, 32'h00000000} /* (25, 7, 12) {real, imag} */,
  {32'h44c978ae, 32'h00000000} /* (25, 7, 11) {real, imag} */,
  {32'h43f54220, 32'h00000000} /* (25, 7, 10) {real, imag} */,
  {32'hc41bd5a0, 32'h00000000} /* (25, 7, 9) {real, imag} */,
  {32'hc4dff0bf, 32'h00000000} /* (25, 7, 8) {real, imag} */,
  {32'hc5070553, 32'h00000000} /* (25, 7, 7) {real, imag} */,
  {32'hc4fc6fba, 32'h00000000} /* (25, 7, 6) {real, imag} */,
  {32'hc566986b, 32'h00000000} /* (25, 7, 5) {real, imag} */,
  {32'hc584ddf8, 32'h00000000} /* (25, 7, 4) {real, imag} */,
  {32'hc5500622, 32'h00000000} /* (25, 7, 3) {real, imag} */,
  {32'hc5a62626, 32'h00000000} /* (25, 7, 2) {real, imag} */,
  {32'hc5be583c, 32'h00000000} /* (25, 7, 1) {real, imag} */,
  {32'hc591c338, 32'h00000000} /* (25, 7, 0) {real, imag} */,
  {32'hc5b9b636, 32'h00000000} /* (25, 6, 31) {real, imag} */,
  {32'hc5cd3e6c, 32'h00000000} /* (25, 6, 30) {real, imag} */,
  {32'hc5cf1070, 32'h00000000} /* (25, 6, 29) {real, imag} */,
  {32'hc5e81cdc, 32'h00000000} /* (25, 6, 28) {real, imag} */,
  {32'hc5ca6d33, 32'h00000000} /* (25, 6, 27) {real, imag} */,
  {32'hc5b5ba6b, 32'h00000000} /* (25, 6, 26) {real, imag} */,
  {32'hc5cbec16, 32'h00000000} /* (25, 6, 25) {real, imag} */,
  {32'hc5b8b527, 32'h00000000} /* (25, 6, 24) {real, imag} */,
  {32'hc59f2d81, 32'h00000000} /* (25, 6, 23) {real, imag} */,
  {32'hc578f2be, 32'h00000000} /* (25, 6, 22) {real, imag} */,
  {32'hc55917e2, 32'h00000000} /* (25, 6, 21) {real, imag} */,
  {32'hc4a6cf31, 32'h00000000} /* (25, 6, 20) {real, imag} */,
  {32'hc48f6da5, 32'h00000000} /* (25, 6, 19) {real, imag} */,
  {32'h42df9460, 32'h00000000} /* (25, 6, 18) {real, imag} */,
  {32'h44632190, 32'h00000000} /* (25, 6, 17) {real, imag} */,
  {32'h449d9946, 32'h00000000} /* (25, 6, 16) {real, imag} */,
  {32'h44f7b7e8, 32'h00000000} /* (25, 6, 15) {real, imag} */,
  {32'h45305521, 32'h00000000} /* (25, 6, 14) {real, imag} */,
  {32'h452901d4, 32'h00000000} /* (25, 6, 13) {real, imag} */,
  {32'h45402498, 32'h00000000} /* (25, 6, 12) {real, imag} */,
  {32'h45048d56, 32'h00000000} /* (25, 6, 11) {real, imag} */,
  {32'h43fdbdf0, 32'h00000000} /* (25, 6, 10) {real, imag} */,
  {32'hc2ff0020, 32'h00000000} /* (25, 6, 9) {real, imag} */,
  {32'hc3106540, 32'h00000000} /* (25, 6, 8) {real, imag} */,
  {32'hc4845154, 32'h00000000} /* (25, 6, 7) {real, imag} */,
  {32'hc5231cec, 32'h00000000} /* (25, 6, 6) {real, imag} */,
  {32'hc54c7232, 32'h00000000} /* (25, 6, 5) {real, imag} */,
  {32'hc5923364, 32'h00000000} /* (25, 6, 4) {real, imag} */,
  {32'hc5913245, 32'h00000000} /* (25, 6, 3) {real, imag} */,
  {32'hc5978f12, 32'h00000000} /* (25, 6, 2) {real, imag} */,
  {32'hc5aa04eb, 32'h00000000} /* (25, 6, 1) {real, imag} */,
  {32'hc59fd5ec, 32'h00000000} /* (25, 6, 0) {real, imag} */,
  {32'hc5cd7a5e, 32'h00000000} /* (25, 5, 31) {real, imag} */,
  {32'hc5f090c3, 32'h00000000} /* (25, 5, 30) {real, imag} */,
  {32'hc5e891f4, 32'h00000000} /* (25, 5, 29) {real, imag} */,
  {32'hc5ff8bcc, 32'h00000000} /* (25, 5, 28) {real, imag} */,
  {32'hc5d54030, 32'h00000000} /* (25, 5, 27) {real, imag} */,
  {32'hc5cdc63a, 32'h00000000} /* (25, 5, 26) {real, imag} */,
  {32'hc5dedbbe, 32'h00000000} /* (25, 5, 25) {real, imag} */,
  {32'hc5cb9d4e, 32'h00000000} /* (25, 5, 24) {real, imag} */,
  {32'hc5a25210, 32'h00000000} /* (25, 5, 23) {real, imag} */,
  {32'hc59956a2, 32'h00000000} /* (25, 5, 22) {real, imag} */,
  {32'hc581f29a, 32'h00000000} /* (25, 5, 21) {real, imag} */,
  {32'hc5381f8e, 32'h00000000} /* (25, 5, 20) {real, imag} */,
  {32'hc5044ff2, 32'h00000000} /* (25, 5, 19) {real, imag} */,
  {32'hc49b5e88, 32'h00000000} /* (25, 5, 18) {real, imag} */,
  {32'hc40b9f1c, 32'h00000000} /* (25, 5, 17) {real, imag} */,
  {32'h447b4b10, 32'h00000000} /* (25, 5, 16) {real, imag} */,
  {32'h450c2c83, 32'h00000000} /* (25, 5, 15) {real, imag} */,
  {32'h4507b326, 32'h00000000} /* (25, 5, 14) {real, imag} */,
  {32'h452e46f8, 32'h00000000} /* (25, 5, 13) {real, imag} */,
  {32'h4538dd2b, 32'h00000000} /* (25, 5, 12) {real, imag} */,
  {32'h451022d8, 32'h00000000} /* (25, 5, 11) {real, imag} */,
  {32'h44bb4cfe, 32'h00000000} /* (25, 5, 10) {real, imag} */,
  {32'h4480e57a, 32'h00000000} /* (25, 5, 9) {real, imag} */,
  {32'h44460038, 32'h00000000} /* (25, 5, 8) {real, imag} */,
  {32'h441923e8, 32'h00000000} /* (25, 5, 7) {real, imag} */,
  {32'hc49882d0, 32'h00000000} /* (25, 5, 6) {real, imag} */,
  {32'hc57c9c07, 32'h00000000} /* (25, 5, 5) {real, imag} */,
  {32'hc564b228, 32'h00000000} /* (25, 5, 4) {real, imag} */,
  {32'hc5a67f6f, 32'h00000000} /* (25, 5, 3) {real, imag} */,
  {32'hc5abfd62, 32'h00000000} /* (25, 5, 2) {real, imag} */,
  {32'hc5e0bb0a, 32'h00000000} /* (25, 5, 1) {real, imag} */,
  {32'hc5b62085, 32'h00000000} /* (25, 5, 0) {real, imag} */,
  {32'hc5cda57e, 32'h00000000} /* (25, 4, 31) {real, imag} */,
  {32'hc5eb1493, 32'h00000000} /* (25, 4, 30) {real, imag} */,
  {32'hc5fbef21, 32'h00000000} /* (25, 4, 29) {real, imag} */,
  {32'hc5f821f4, 32'h00000000} /* (25, 4, 28) {real, imag} */,
  {32'hc608525c, 32'h00000000} /* (25, 4, 27) {real, imag} */,
  {32'hc5da9042, 32'h00000000} /* (25, 4, 26) {real, imag} */,
  {32'hc5db6d08, 32'h00000000} /* (25, 4, 25) {real, imag} */,
  {32'hc5d8a6ed, 32'h00000000} /* (25, 4, 24) {real, imag} */,
  {32'hc5c80963, 32'h00000000} /* (25, 4, 23) {real, imag} */,
  {32'hc5988e49, 32'h00000000} /* (25, 4, 22) {real, imag} */,
  {32'hc584d148, 32'h00000000} /* (25, 4, 21) {real, imag} */,
  {32'hc5670f5a, 32'h00000000} /* (25, 4, 20) {real, imag} */,
  {32'hc5459bba, 32'h00000000} /* (25, 4, 19) {real, imag} */,
  {32'hc516404e, 32'h00000000} /* (25, 4, 18) {real, imag} */,
  {32'hc4bf07c5, 32'h00000000} /* (25, 4, 17) {real, imag} */,
  {32'hc42f9ee8, 32'h00000000} /* (25, 4, 16) {real, imag} */,
  {32'h44f8e072, 32'h00000000} /* (25, 4, 15) {real, imag} */,
  {32'h451b0002, 32'h00000000} /* (25, 4, 14) {real, imag} */,
  {32'h451613d2, 32'h00000000} /* (25, 4, 13) {real, imag} */,
  {32'h452fac05, 32'h00000000} /* (25, 4, 12) {real, imag} */,
  {32'h4542dd65, 32'h00000000} /* (25, 4, 11) {real, imag} */,
  {32'h450f743c, 32'h00000000} /* (25, 4, 10) {real, imag} */,
  {32'h44e2f25e, 32'h00000000} /* (25, 4, 9) {real, imag} */,
  {32'h4512ef66, 32'h00000000} /* (25, 4, 8) {real, imag} */,
  {32'h445585c0, 32'h00000000} /* (25, 4, 7) {real, imag} */,
  {32'h43703ee0, 32'h00000000} /* (25, 4, 6) {real, imag} */,
  {32'hc51a844f, 32'h00000000} /* (25, 4, 5) {real, imag} */,
  {32'hc58b3324, 32'h00000000} /* (25, 4, 4) {real, imag} */,
  {32'hc5825996, 32'h00000000} /* (25, 4, 3) {real, imag} */,
  {32'hc5abad49, 32'h00000000} /* (25, 4, 2) {real, imag} */,
  {32'hc5a9f482, 32'h00000000} /* (25, 4, 1) {real, imag} */,
  {32'hc5be58bf, 32'h00000000} /* (25, 4, 0) {real, imag} */,
  {32'hc5d02960, 32'h00000000} /* (25, 3, 31) {real, imag} */,
  {32'hc5e587f6, 32'h00000000} /* (25, 3, 30) {real, imag} */,
  {32'hc5fd4595, 32'h00000000} /* (25, 3, 29) {real, imag} */,
  {32'hc60b5dba, 32'h00000000} /* (25, 3, 28) {real, imag} */,
  {32'hc610f7d4, 32'h00000000} /* (25, 3, 27) {real, imag} */,
  {32'hc5f472f6, 32'h00000000} /* (25, 3, 26) {real, imag} */,
  {32'hc5decc24, 32'h00000000} /* (25, 3, 25) {real, imag} */,
  {32'hc5e03909, 32'h00000000} /* (25, 3, 24) {real, imag} */,
  {32'hc5c41796, 32'h00000000} /* (25, 3, 23) {real, imag} */,
  {32'hc5ab51dc, 32'h00000000} /* (25, 3, 22) {real, imag} */,
  {32'hc5901a11, 32'h00000000} /* (25, 3, 21) {real, imag} */,
  {32'hc58de7f5, 32'h00000000} /* (25, 3, 20) {real, imag} */,
  {32'hc556b1c3, 32'h00000000} /* (25, 3, 19) {real, imag} */,
  {32'hc4ba3338, 32'h00000000} /* (25, 3, 18) {real, imag} */,
  {32'hc4ba9122, 32'h00000000} /* (25, 3, 17) {real, imag} */,
  {32'hc49d10dc, 32'h00000000} /* (25, 3, 16) {real, imag} */,
  {32'h448366ae, 32'h00000000} /* (25, 3, 15) {real, imag} */,
  {32'h450d9b35, 32'h00000000} /* (25, 3, 14) {real, imag} */,
  {32'h457c18de, 32'h00000000} /* (25, 3, 13) {real, imag} */,
  {32'h452f28b8, 32'h00000000} /* (25, 3, 12) {real, imag} */,
  {32'h45702c39, 32'h00000000} /* (25, 3, 11) {real, imag} */,
  {32'h4541e999, 32'h00000000} /* (25, 3, 10) {real, imag} */,
  {32'h44eae310, 32'h00000000} /* (25, 3, 9) {real, imag} */,
  {32'h450d3f62, 32'h00000000} /* (25, 3, 8) {real, imag} */,
  {32'h45094550, 32'h00000000} /* (25, 3, 7) {real, imag} */,
  {32'h40ed0e00, 32'h00000000} /* (25, 3, 6) {real, imag} */,
  {32'hc515fa06, 32'h00000000} /* (25, 3, 5) {real, imag} */,
  {32'hc59befab, 32'h00000000} /* (25, 3, 4) {real, imag} */,
  {32'hc5a2216a, 32'h00000000} /* (25, 3, 3) {real, imag} */,
  {32'hc5aa873d, 32'h00000000} /* (25, 3, 2) {real, imag} */,
  {32'hc5ccb90e, 32'h00000000} /* (25, 3, 1) {real, imag} */,
  {32'hc5cffb69, 32'h00000000} /* (25, 3, 0) {real, imag} */,
  {32'hc5c9e5f5, 32'h00000000} /* (25, 2, 31) {real, imag} */,
  {32'hc5f0e860, 32'h00000000} /* (25, 2, 30) {real, imag} */,
  {32'hc5fede01, 32'h00000000} /* (25, 2, 29) {real, imag} */,
  {32'hc60f6583, 32'h00000000} /* (25, 2, 28) {real, imag} */,
  {32'hc60a16ab, 32'h00000000} /* (25, 2, 27) {real, imag} */,
  {32'hc5e9730e, 32'h00000000} /* (25, 2, 26) {real, imag} */,
  {32'hc5d02f70, 32'h00000000} /* (25, 2, 25) {real, imag} */,
  {32'hc5cd6602, 32'h00000000} /* (25, 2, 24) {real, imag} */,
  {32'hc5c2c584, 32'h00000000} /* (25, 2, 23) {real, imag} */,
  {32'hc5a0ac33, 32'h00000000} /* (25, 2, 22) {real, imag} */,
  {32'hc5926bd6, 32'h00000000} /* (25, 2, 21) {real, imag} */,
  {32'hc5936101, 32'h00000000} /* (25, 2, 20) {real, imag} */,
  {32'hc52fae8a, 32'h00000000} /* (25, 2, 19) {real, imag} */,
  {32'hc520fe4c, 32'h00000000} /* (25, 2, 18) {real, imag} */,
  {32'hc492b512, 32'h00000000} /* (25, 2, 17) {real, imag} */,
  {32'h43f62d80, 32'h00000000} /* (25, 2, 16) {real, imag} */,
  {32'h45003f5e, 32'h00000000} /* (25, 2, 15) {real, imag} */,
  {32'h4520d249, 32'h00000000} /* (25, 2, 14) {real, imag} */,
  {32'h4549ac52, 32'h00000000} /* (25, 2, 13) {real, imag} */,
  {32'h457c6669, 32'h00000000} /* (25, 2, 12) {real, imag} */,
  {32'h4547232c, 32'h00000000} /* (25, 2, 11) {real, imag} */,
  {32'h451671c3, 32'h00000000} /* (25, 2, 10) {real, imag} */,
  {32'h453b3363, 32'h00000000} /* (25, 2, 9) {real, imag} */,
  {32'h449147c8, 32'h00000000} /* (25, 2, 8) {real, imag} */,
  {32'h44a2d968, 32'h00000000} /* (25, 2, 7) {real, imag} */,
  {32'h44852c18, 32'h00000000} /* (25, 2, 6) {real, imag} */,
  {32'hc538a655, 32'h00000000} /* (25, 2, 5) {real, imag} */,
  {32'hc59fc0e7, 32'h00000000} /* (25, 2, 4) {real, imag} */,
  {32'hc5a82c3b, 32'h00000000} /* (25, 2, 3) {real, imag} */,
  {32'hc5b26a06, 32'h00000000} /* (25, 2, 2) {real, imag} */,
  {32'hc5c25d0c, 32'h00000000} /* (25, 2, 1) {real, imag} */,
  {32'hc5c57c16, 32'h00000000} /* (25, 2, 0) {real, imag} */,
  {32'hc5ca9236, 32'h00000000} /* (25, 1, 31) {real, imag} */,
  {32'hc5f935ed, 32'h00000000} /* (25, 1, 30) {real, imag} */,
  {32'hc5e88140, 32'h00000000} /* (25, 1, 29) {real, imag} */,
  {32'hc60e1f7e, 32'h00000000} /* (25, 1, 28) {real, imag} */,
  {32'hc60295e3, 32'h00000000} /* (25, 1, 27) {real, imag} */,
  {32'hc5f5e5ae, 32'h00000000} /* (25, 1, 26) {real, imag} */,
  {32'hc5d806eb, 32'h00000000} /* (25, 1, 25) {real, imag} */,
  {32'hc5c21321, 32'h00000000} /* (25, 1, 24) {real, imag} */,
  {32'hc5b34c52, 32'h00000000} /* (25, 1, 23) {real, imag} */,
  {32'hc58e4bb8, 32'h00000000} /* (25, 1, 22) {real, imag} */,
  {32'hc5a8695a, 32'h00000000} /* (25, 1, 21) {real, imag} */,
  {32'hc552833a, 32'h00000000} /* (25, 1, 20) {real, imag} */,
  {32'hc5303b54, 32'h00000000} /* (25, 1, 19) {real, imag} */,
  {32'hc4d0699c, 32'h00000000} /* (25, 1, 18) {real, imag} */,
  {32'hc4af2ad8, 32'h00000000} /* (25, 1, 17) {real, imag} */,
  {32'hc448f7d4, 32'h00000000} /* (25, 1, 16) {real, imag} */,
  {32'h44f3745a, 32'h00000000} /* (25, 1, 15) {real, imag} */,
  {32'h453787e6, 32'h00000000} /* (25, 1, 14) {real, imag} */,
  {32'h44d1de20, 32'h00000000} /* (25, 1, 13) {real, imag} */,
  {32'h4516f6be, 32'h00000000} /* (25, 1, 12) {real, imag} */,
  {32'h4532d274, 32'h00000000} /* (25, 1, 11) {real, imag} */,
  {32'h451b98bc, 32'h00000000} /* (25, 1, 10) {real, imag} */,
  {32'h44d81ffc, 32'h00000000} /* (25, 1, 9) {real, imag} */,
  {32'h44ba2fbc, 32'h00000000} /* (25, 1, 8) {real, imag} */,
  {32'hc3012e90, 32'h00000000} /* (25, 1, 7) {real, imag} */,
  {32'hc4afc6d6, 32'h00000000} /* (25, 1, 6) {real, imag} */,
  {32'hc52d906b, 32'h00000000} /* (25, 1, 5) {real, imag} */,
  {32'hc58d3c5d, 32'h00000000} /* (25, 1, 4) {real, imag} */,
  {32'hc5a28730, 32'h00000000} /* (25, 1, 3) {real, imag} */,
  {32'hc5b018b5, 32'h00000000} /* (25, 1, 2) {real, imag} */,
  {32'hc5b5a452, 32'h00000000} /* (25, 1, 1) {real, imag} */,
  {32'hc5c4dc52, 32'h00000000} /* (25, 1, 0) {real, imag} */,
  {32'hc5d066c0, 32'h00000000} /* (25, 0, 31) {real, imag} */,
  {32'hc5d4c487, 32'h00000000} /* (25, 0, 30) {real, imag} */,
  {32'hc5e6a1cc, 32'h00000000} /* (25, 0, 29) {real, imag} */,
  {32'hc5f4c345, 32'h00000000} /* (25, 0, 28) {real, imag} */,
  {32'hc5f2baa2, 32'h00000000} /* (25, 0, 27) {real, imag} */,
  {32'hc5f0dbaa, 32'h00000000} /* (25, 0, 26) {real, imag} */,
  {32'hc5c7b618, 32'h00000000} /* (25, 0, 25) {real, imag} */,
  {32'hc5b8201f, 32'h00000000} /* (25, 0, 24) {real, imag} */,
  {32'hc5a04321, 32'h00000000} /* (25, 0, 23) {real, imag} */,
  {32'hc59335fa, 32'h00000000} /* (25, 0, 22) {real, imag} */,
  {32'hc5679b3c, 32'h00000000} /* (25, 0, 21) {real, imag} */,
  {32'hc5177e66, 32'h00000000} /* (25, 0, 20) {real, imag} */,
  {32'hc4aa24bd, 32'h00000000} /* (25, 0, 19) {real, imag} */,
  {32'hc42a85d4, 32'h00000000} /* (25, 0, 18) {real, imag} */,
  {32'hc3d4c258, 32'h00000000} /* (25, 0, 17) {real, imag} */,
  {32'h44375234, 32'h00000000} /* (25, 0, 16) {real, imag} */,
  {32'h44a6c7ee, 32'h00000000} /* (25, 0, 15) {real, imag} */,
  {32'h44e12054, 32'h00000000} /* (25, 0, 14) {real, imag} */,
  {32'h45053fb1, 32'h00000000} /* (25, 0, 13) {real, imag} */,
  {32'h450be142, 32'h00000000} /* (25, 0, 12) {real, imag} */,
  {32'h44da3c26, 32'h00000000} /* (25, 0, 11) {real, imag} */,
  {32'h449e2618, 32'h00000000} /* (25, 0, 10) {real, imag} */,
  {32'h438ba6a8, 32'h00000000} /* (25, 0, 9) {real, imag} */,
  {32'hc32bb0e0, 32'h00000000} /* (25, 0, 8) {real, imag} */,
  {32'hc45117d8, 32'h00000000} /* (25, 0, 7) {real, imag} */,
  {32'hc4fe54f1, 32'h00000000} /* (25, 0, 6) {real, imag} */,
  {32'hc54ce9ca, 32'h00000000} /* (25, 0, 5) {real, imag} */,
  {32'hc588977b, 32'h00000000} /* (25, 0, 4) {real, imag} */,
  {32'hc5a09c34, 32'h00000000} /* (25, 0, 3) {real, imag} */,
  {32'hc5ca18fe, 32'h00000000} /* (25, 0, 2) {real, imag} */,
  {32'hc5ca8f0a, 32'h00000000} /* (25, 0, 1) {real, imag} */,
  {32'hc5b3229a, 32'h00000000} /* (25, 0, 0) {real, imag} */,
  {32'hc60fbc48, 32'h00000000} /* (24, 31, 31) {real, imag} */,
  {32'hc621eef0, 32'h00000000} /* (24, 31, 30) {real, imag} */,
  {32'hc626b856, 32'h00000000} /* (24, 31, 29) {real, imag} */,
  {32'hc625ea2f, 32'h00000000} /* (24, 31, 28) {real, imag} */,
  {32'hc632e088, 32'h00000000} /* (24, 31, 27) {real, imag} */,
  {32'hc61c13bc, 32'h00000000} /* (24, 31, 26) {real, imag} */,
  {32'hc611eff9, 32'h00000000} /* (24, 31, 25) {real, imag} */,
  {32'hc60c7b0a, 32'h00000000} /* (24, 31, 24) {real, imag} */,
  {32'hc5e8b32d, 32'h00000000} /* (24, 31, 23) {real, imag} */,
  {32'hc5cf7b33, 32'h00000000} /* (24, 31, 22) {real, imag} */,
  {32'hc58d7b8b, 32'h00000000} /* (24, 31, 21) {real, imag} */,
  {32'hc50a3c8b, 32'h00000000} /* (24, 31, 20) {real, imag} */,
  {32'h430f4850, 32'h00000000} /* (24, 31, 19) {real, imag} */,
  {32'h4413ee30, 32'h00000000} /* (24, 31, 18) {real, imag} */,
  {32'h44b3bc1c, 32'h00000000} /* (24, 31, 17) {real, imag} */,
  {32'h452e4aea, 32'h00000000} /* (24, 31, 16) {real, imag} */,
  {32'h4546d11d, 32'h00000000} /* (24, 31, 15) {real, imag} */,
  {32'h456adc80, 32'h00000000} /* (24, 31, 14) {real, imag} */,
  {32'h456b4680, 32'h00000000} /* (24, 31, 13) {real, imag} */,
  {32'h454f4863, 32'h00000000} /* (24, 31, 12) {real, imag} */,
  {32'h4515f0e6, 32'h00000000} /* (24, 31, 11) {real, imag} */,
  {32'hc330e280, 32'h00000000} /* (24, 31, 10) {real, imag} */,
  {32'hc429a090, 32'h00000000} /* (24, 31, 9) {real, imag} */,
  {32'hc51862d9, 32'h00000000} /* (24, 31, 8) {real, imag} */,
  {32'hc52a5b86, 32'h00000000} /* (24, 31, 7) {real, imag} */,
  {32'hc58e8425, 32'h00000000} /* (24, 31, 6) {real, imag} */,
  {32'hc5bc373d, 32'h00000000} /* (24, 31, 5) {real, imag} */,
  {32'hc5cee0cc, 32'h00000000} /* (24, 31, 4) {real, imag} */,
  {32'hc5e264a8, 32'h00000000} /* (24, 31, 3) {real, imag} */,
  {32'hc5ff6aaa, 32'h00000000} /* (24, 31, 2) {real, imag} */,
  {32'hc608d244, 32'h00000000} /* (24, 31, 1) {real, imag} */,
  {32'hc608962e, 32'h00000000} /* (24, 31, 0) {real, imag} */,
  {32'hc613a56a, 32'h00000000} /* (24, 30, 31) {real, imag} */,
  {32'hc6254504, 32'h00000000} /* (24, 30, 30) {real, imag} */,
  {32'hc62667f2, 32'h00000000} /* (24, 30, 29) {real, imag} */,
  {32'hc6293646, 32'h00000000} /* (24, 30, 28) {real, imag} */,
  {32'hc6302276, 32'h00000000} /* (24, 30, 27) {real, imag} */,
  {32'hc61d8a90, 32'h00000000} /* (24, 30, 26) {real, imag} */,
  {32'hc61f450b, 32'h00000000} /* (24, 30, 25) {real, imag} */,
  {32'hc6081a8e, 32'h00000000} /* (24, 30, 24) {real, imag} */,
  {32'hc5e5dd68, 32'h00000000} /* (24, 30, 23) {real, imag} */,
  {32'hc5e11ae0, 32'h00000000} /* (24, 30, 22) {real, imag} */,
  {32'hc57d3878, 32'h00000000} /* (24, 30, 21) {real, imag} */,
  {32'hc3b2cb88, 32'h00000000} /* (24, 30, 20) {real, imag} */,
  {32'h44282bfc, 32'h00000000} /* (24, 30, 19) {real, imag} */,
  {32'h45219f12, 32'h00000000} /* (24, 30, 18) {real, imag} */,
  {32'h45628227, 32'h00000000} /* (24, 30, 17) {real, imag} */,
  {32'h45820faf, 32'h00000000} /* (24, 30, 16) {real, imag} */,
  {32'h458011da, 32'h00000000} /* (24, 30, 15) {real, imag} */,
  {32'h4595327f, 32'h00000000} /* (24, 30, 14) {real, imag} */,
  {32'h4577d676, 32'h00000000} /* (24, 30, 13) {real, imag} */,
  {32'h45635bc9, 32'h00000000} /* (24, 30, 12) {real, imag} */,
  {32'h4543bd07, 32'h00000000} /* (24, 30, 11) {real, imag} */,
  {32'hc3c834e0, 32'h00000000} /* (24, 30, 10) {real, imag} */,
  {32'hc4fb1f78, 32'h00000000} /* (24, 30, 9) {real, imag} */,
  {32'hc578ec46, 32'h00000000} /* (24, 30, 8) {real, imag} */,
  {32'hc59294b6, 32'h00000000} /* (24, 30, 7) {real, imag} */,
  {32'hc5c24df8, 32'h00000000} /* (24, 30, 6) {real, imag} */,
  {32'hc5df68d2, 32'h00000000} /* (24, 30, 5) {real, imag} */,
  {32'hc5e6e2d6, 32'h00000000} /* (24, 30, 4) {real, imag} */,
  {32'hc606ba46, 32'h00000000} /* (24, 30, 3) {real, imag} */,
  {32'hc609cf3e, 32'h00000000} /* (24, 30, 2) {real, imag} */,
  {32'hc609c57b, 32'h00000000} /* (24, 30, 1) {real, imag} */,
  {32'hc60c09de, 32'h00000000} /* (24, 30, 0) {real, imag} */,
  {32'hc6171eaf, 32'h00000000} /* (24, 29, 31) {real, imag} */,
  {32'hc62f80e5, 32'h00000000} /* (24, 29, 30) {real, imag} */,
  {32'hc6304dd7, 32'h00000000} /* (24, 29, 29) {real, imag} */,
  {32'hc6270250, 32'h00000000} /* (24, 29, 28) {real, imag} */,
  {32'hc626af00, 32'h00000000} /* (24, 29, 27) {real, imag} */,
  {32'hc624d96a, 32'h00000000} /* (24, 29, 26) {real, imag} */,
  {32'hc627b898, 32'h00000000} /* (24, 29, 25) {real, imag} */,
  {32'hc60c5246, 32'h00000000} /* (24, 29, 24) {real, imag} */,
  {32'hc5e63689, 32'h00000000} /* (24, 29, 23) {real, imag} */,
  {32'hc5bd66f6, 32'h00000000} /* (24, 29, 22) {real, imag} */,
  {32'hc5513aea, 32'h00000000} /* (24, 29, 21) {real, imag} */,
  {32'hc389d540, 32'h00000000} /* (24, 29, 20) {real, imag} */,
  {32'h449928cc, 32'h00000000} /* (24, 29, 19) {real, imag} */,
  {32'h4544d4ba, 32'h00000000} /* (24, 29, 18) {real, imag} */,
  {32'h457da124, 32'h00000000} /* (24, 29, 17) {real, imag} */,
  {32'h458e5068, 32'h00000000} /* (24, 29, 16) {real, imag} */,
  {32'h4591975e, 32'h00000000} /* (24, 29, 15) {real, imag} */,
  {32'h4596708a, 32'h00000000} /* (24, 29, 14) {real, imag} */,
  {32'h45812bb0, 32'h00000000} /* (24, 29, 13) {real, imag} */,
  {32'h457fd503, 32'h00000000} /* (24, 29, 12) {real, imag} */,
  {32'h44e913e4, 32'h00000000} /* (24, 29, 11) {real, imag} */,
  {32'hc3532a60, 32'h00000000} /* (24, 29, 10) {real, imag} */,
  {32'hc5153036, 32'h00000000} /* (24, 29, 9) {real, imag} */,
  {32'hc595d048, 32'h00000000} /* (24, 29, 8) {real, imag} */,
  {32'hc5cf1d83, 32'h00000000} /* (24, 29, 7) {real, imag} */,
  {32'hc5be9b3e, 32'h00000000} /* (24, 29, 6) {real, imag} */,
  {32'hc5d5e943, 32'h00000000} /* (24, 29, 5) {real, imag} */,
  {32'hc5d2907d, 32'h00000000} /* (24, 29, 4) {real, imag} */,
  {32'hc61211b0, 32'h00000000} /* (24, 29, 3) {real, imag} */,
  {32'hc614d512, 32'h00000000} /* (24, 29, 2) {real, imag} */,
  {32'hc61215e7, 32'h00000000} /* (24, 29, 1) {real, imag} */,
  {32'hc61527b1, 32'h00000000} /* (24, 29, 0) {real, imag} */,
  {32'hc61b63a8, 32'h00000000} /* (24, 28, 31) {real, imag} */,
  {32'hc62fbb74, 32'h00000000} /* (24, 28, 30) {real, imag} */,
  {32'hc6340541, 32'h00000000} /* (24, 28, 29) {real, imag} */,
  {32'hc6267d5c, 32'h00000000} /* (24, 28, 28) {real, imag} */,
  {32'hc6283104, 32'h00000000} /* (24, 28, 27) {real, imag} */,
  {32'hc634859e, 32'h00000000} /* (24, 28, 26) {real, imag} */,
  {32'hc613e2d0, 32'h00000000} /* (24, 28, 25) {real, imag} */,
  {32'hc60d6c8a, 32'h00000000} /* (24, 28, 24) {real, imag} */,
  {32'hc5f81cf3, 32'h00000000} /* (24, 28, 23) {real, imag} */,
  {32'hc5c9d824, 32'h00000000} /* (24, 28, 22) {real, imag} */,
  {32'hc5893540, 32'h00000000} /* (24, 28, 21) {real, imag} */,
  {32'hc3b1a360, 32'h00000000} /* (24, 28, 20) {real, imag} */,
  {32'h4516ab4a, 32'h00000000} /* (24, 28, 19) {real, imag} */,
  {32'h45658c41, 32'h00000000} /* (24, 28, 18) {real, imag} */,
  {32'h4593e967, 32'h00000000} /* (24, 28, 17) {real, imag} */,
  {32'h45b68e57, 32'h00000000} /* (24, 28, 16) {real, imag} */,
  {32'h45b1b7f5, 32'h00000000} /* (24, 28, 15) {real, imag} */,
  {32'h458d0ac0, 32'h00000000} /* (24, 28, 14) {real, imag} */,
  {32'h4581dbca, 32'h00000000} /* (24, 28, 13) {real, imag} */,
  {32'h4553d363, 32'h00000000} /* (24, 28, 12) {real, imag} */,
  {32'h4523fd5e, 32'h00000000} /* (24, 28, 11) {real, imag} */,
  {32'hc4b1c254, 32'h00000000} /* (24, 28, 10) {real, imag} */,
  {32'hc57c3036, 32'h00000000} /* (24, 28, 9) {real, imag} */,
  {32'hc59dfada, 32'h00000000} /* (24, 28, 8) {real, imag} */,
  {32'hc5cf3483, 32'h00000000} /* (24, 28, 7) {real, imag} */,
  {32'hc5d3b91c, 32'h00000000} /* (24, 28, 6) {real, imag} */,
  {32'hc5ddf40c, 32'h00000000} /* (24, 28, 5) {real, imag} */,
  {32'hc6099a7a, 32'h00000000} /* (24, 28, 4) {real, imag} */,
  {32'hc618a94e, 32'h00000000} /* (24, 28, 3) {real, imag} */,
  {32'hc616a004, 32'h00000000} /* (24, 28, 2) {real, imag} */,
  {32'hc6229ba4, 32'h00000000} /* (24, 28, 1) {real, imag} */,
  {32'hc61fcdbc, 32'h00000000} /* (24, 28, 0) {real, imag} */,
  {32'hc6189455, 32'h00000000} /* (24, 27, 31) {real, imag} */,
  {32'hc61d48c4, 32'h00000000} /* (24, 27, 30) {real, imag} */,
  {32'hc624cb9b, 32'h00000000} /* (24, 27, 29) {real, imag} */,
  {32'hc61bb780, 32'h00000000} /* (24, 27, 28) {real, imag} */,
  {32'hc61d48d8, 32'h00000000} /* (24, 27, 27) {real, imag} */,
  {32'hc64097b4, 32'h00000000} /* (24, 27, 26) {real, imag} */,
  {32'hc624603e, 32'h00000000} /* (24, 27, 25) {real, imag} */,
  {32'hc60bfabb, 32'h00000000} /* (24, 27, 24) {real, imag} */,
  {32'hc5f3eb7f, 32'h00000000} /* (24, 27, 23) {real, imag} */,
  {32'hc5a8a436, 32'h00000000} /* (24, 27, 22) {real, imag} */,
  {32'hc55d703e, 32'h00000000} /* (24, 27, 21) {real, imag} */,
  {32'hc42abd38, 32'h00000000} /* (24, 27, 20) {real, imag} */,
  {32'h451791f2, 32'h00000000} /* (24, 27, 19) {real, imag} */,
  {32'h4594b904, 32'h00000000} /* (24, 27, 18) {real, imag} */,
  {32'h459c0956, 32'h00000000} /* (24, 27, 17) {real, imag} */,
  {32'h45a0fab8, 32'h00000000} /* (24, 27, 16) {real, imag} */,
  {32'h459bf4b8, 32'h00000000} /* (24, 27, 15) {real, imag} */,
  {32'h4584d582, 32'h00000000} /* (24, 27, 14) {real, imag} */,
  {32'h458c7e42, 32'h00000000} /* (24, 27, 13) {real, imag} */,
  {32'h45656d82, 32'h00000000} /* (24, 27, 12) {real, imag} */,
  {32'h451a1eea, 32'h00000000} /* (24, 27, 11) {real, imag} */,
  {32'hc4d4ca74, 32'h00000000} /* (24, 27, 10) {real, imag} */,
  {32'hc583c453, 32'h00000000} /* (24, 27, 9) {real, imag} */,
  {32'hc5a6f77e, 32'h00000000} /* (24, 27, 8) {real, imag} */,
  {32'hc5aa52af, 32'h00000000} /* (24, 27, 7) {real, imag} */,
  {32'hc5da58fc, 32'h00000000} /* (24, 27, 6) {real, imag} */,
  {32'hc5fadd85, 32'h00000000} /* (24, 27, 5) {real, imag} */,
  {32'hc612b672, 32'h00000000} /* (24, 27, 4) {real, imag} */,
  {32'hc619db34, 32'h00000000} /* (24, 27, 3) {real, imag} */,
  {32'hc619166b, 32'h00000000} /* (24, 27, 2) {real, imag} */,
  {32'hc618fc43, 32'h00000000} /* (24, 27, 1) {real, imag} */,
  {32'hc60f1174, 32'h00000000} /* (24, 27, 0) {real, imag} */,
  {32'hc60a2b62, 32'h00000000} /* (24, 26, 31) {real, imag} */,
  {32'hc61a1b44, 32'h00000000} /* (24, 26, 30) {real, imag} */,
  {32'hc61ae582, 32'h00000000} /* (24, 26, 29) {real, imag} */,
  {32'hc617e7da, 32'h00000000} /* (24, 26, 28) {real, imag} */,
  {32'hc6240dcf, 32'h00000000} /* (24, 26, 27) {real, imag} */,
  {32'hc630acf0, 32'h00000000} /* (24, 26, 26) {real, imag} */,
  {32'hc61b62e2, 32'h00000000} /* (24, 26, 25) {real, imag} */,
  {32'hc6027457, 32'h00000000} /* (24, 26, 24) {real, imag} */,
  {32'hc5d53ab4, 32'h00000000} /* (24, 26, 23) {real, imag} */,
  {32'hc593aa36, 32'h00000000} /* (24, 26, 22) {real, imag} */,
  {32'hc54fa756, 32'h00000000} /* (24, 26, 21) {real, imag} */,
  {32'h43321f20, 32'h00000000} /* (24, 26, 20) {real, imag} */,
  {32'h452cecbb, 32'h00000000} /* (24, 26, 19) {real, imag} */,
  {32'h4589db34, 32'h00000000} /* (24, 26, 18) {real, imag} */,
  {32'h45996392, 32'h00000000} /* (24, 26, 17) {real, imag} */,
  {32'h45aa4c9a, 32'h00000000} /* (24, 26, 16) {real, imag} */,
  {32'h459f2a4f, 32'h00000000} /* (24, 26, 15) {real, imag} */,
  {32'h459ccf09, 32'h00000000} /* (24, 26, 14) {real, imag} */,
  {32'h456ece80, 32'h00000000} /* (24, 26, 13) {real, imag} */,
  {32'h455429b0, 32'h00000000} /* (24, 26, 12) {real, imag} */,
  {32'h43db0160, 32'h00000000} /* (24, 26, 11) {real, imag} */,
  {32'hc51ddd0e, 32'h00000000} /* (24, 26, 10) {real, imag} */,
  {32'hc5834ddb, 32'h00000000} /* (24, 26, 9) {real, imag} */,
  {32'hc5950803, 32'h00000000} /* (24, 26, 8) {real, imag} */,
  {32'hc5c08a2e, 32'h00000000} /* (24, 26, 7) {real, imag} */,
  {32'hc5db217e, 32'h00000000} /* (24, 26, 6) {real, imag} */,
  {32'hc5f4993d, 32'h00000000} /* (24, 26, 5) {real, imag} */,
  {32'hc6031e7e, 32'h00000000} /* (24, 26, 4) {real, imag} */,
  {32'hc612c70b, 32'h00000000} /* (24, 26, 3) {real, imag} */,
  {32'hc60a5cc9, 32'h00000000} /* (24, 26, 2) {real, imag} */,
  {32'hc60586af, 32'h00000000} /* (24, 26, 1) {real, imag} */,
  {32'hc6079eb3, 32'h00000000} /* (24, 26, 0) {real, imag} */,
  {32'hc5fd9da6, 32'h00000000} /* (24, 25, 31) {real, imag} */,
  {32'hc615a392, 32'h00000000} /* (24, 25, 30) {real, imag} */,
  {32'hc6297fd7, 32'h00000000} /* (24, 25, 29) {real, imag} */,
  {32'hc6138e4c, 32'h00000000} /* (24, 25, 28) {real, imag} */,
  {32'hc6195fe4, 32'h00000000} /* (24, 25, 27) {real, imag} */,
  {32'hc60d579a, 32'h00000000} /* (24, 25, 26) {real, imag} */,
  {32'hc6109a9a, 32'h00000000} /* (24, 25, 25) {real, imag} */,
  {32'hc5e4c0f4, 32'h00000000} /* (24, 25, 24) {real, imag} */,
  {32'hc5b8a1c6, 32'h00000000} /* (24, 25, 23) {real, imag} */,
  {32'hc5858827, 32'h00000000} /* (24, 25, 22) {real, imag} */,
  {32'hc4da258e, 32'h00000000} /* (24, 25, 21) {real, imag} */,
  {32'h449827ea, 32'h00000000} /* (24, 25, 20) {real, imag} */,
  {32'h45476ae4, 32'h00000000} /* (24, 25, 19) {real, imag} */,
  {32'h457b4f16, 32'h00000000} /* (24, 25, 18) {real, imag} */,
  {32'h45b45ebf, 32'h00000000} /* (24, 25, 17) {real, imag} */,
  {32'h458cbd44, 32'h00000000} /* (24, 25, 16) {real, imag} */,
  {32'h45969414, 32'h00000000} /* (24, 25, 15) {real, imag} */,
  {32'h45aa3909, 32'h00000000} /* (24, 25, 14) {real, imag} */,
  {32'h4576da28, 32'h00000000} /* (24, 25, 13) {real, imag} */,
  {32'h45090fa1, 32'h00000000} /* (24, 25, 12) {real, imag} */,
  {32'hc3354620, 32'h00000000} /* (24, 25, 11) {real, imag} */,
  {32'hc50a0299, 32'h00000000} /* (24, 25, 10) {real, imag} */,
  {32'hc58b556e, 32'h00000000} /* (24, 25, 9) {real, imag} */,
  {32'hc5bbbb94, 32'h00000000} /* (24, 25, 8) {real, imag} */,
  {32'hc5cb4406, 32'h00000000} /* (24, 25, 7) {real, imag} */,
  {32'hc5c58ac3, 32'h00000000} /* (24, 25, 6) {real, imag} */,
  {32'hc5ec9c0e, 32'h00000000} /* (24, 25, 5) {real, imag} */,
  {32'hc60ec77a, 32'h00000000} /* (24, 25, 4) {real, imag} */,
  {32'hc605df84, 32'h00000000} /* (24, 25, 3) {real, imag} */,
  {32'hc5fa2cb7, 32'h00000000} /* (24, 25, 2) {real, imag} */,
  {32'hc60124fa, 32'h00000000} /* (24, 25, 1) {real, imag} */,
  {32'hc60aa5ce, 32'h00000000} /* (24, 25, 0) {real, imag} */,
  {32'hc5e14e58, 32'h00000000} /* (24, 24, 31) {real, imag} */,
  {32'hc5f7926b, 32'h00000000} /* (24, 24, 30) {real, imag} */,
  {32'hc5ff4bc0, 32'h00000000} /* (24, 24, 29) {real, imag} */,
  {32'hc606e804, 32'h00000000} /* (24, 24, 28) {real, imag} */,
  {32'hc5e56d9e, 32'h00000000} /* (24, 24, 27) {real, imag} */,
  {32'hc5f755c8, 32'h00000000} /* (24, 24, 26) {real, imag} */,
  {32'hc5f1ee12, 32'h00000000} /* (24, 24, 25) {real, imag} */,
  {32'hc5da34ae, 32'h00000000} /* (24, 24, 24) {real, imag} */,
  {32'hc5b4733e, 32'h00000000} /* (24, 24, 23) {real, imag} */,
  {32'hc55b9517, 32'h00000000} /* (24, 24, 22) {real, imag} */,
  {32'hc517007a, 32'h00000000} /* (24, 24, 21) {real, imag} */,
  {32'h444c5bfc, 32'h00000000} /* (24, 24, 20) {real, imag} */,
  {32'h4515f2da, 32'h00000000} /* (24, 24, 19) {real, imag} */,
  {32'h455815e6, 32'h00000000} /* (24, 24, 18) {real, imag} */,
  {32'h45928f12, 32'h00000000} /* (24, 24, 17) {real, imag} */,
  {32'h45a191c3, 32'h00000000} /* (24, 24, 16) {real, imag} */,
  {32'h459b3564, 32'h00000000} /* (24, 24, 15) {real, imag} */,
  {32'h459b2ad1, 32'h00000000} /* (24, 24, 14) {real, imag} */,
  {32'h456e6bbc, 32'h00000000} /* (24, 24, 13) {real, imag} */,
  {32'h44c2addc, 32'h00000000} /* (24, 24, 12) {real, imag} */,
  {32'h440a1480, 32'h00000000} /* (24, 24, 11) {real, imag} */,
  {32'hc50e96a5, 32'h00000000} /* (24, 24, 10) {real, imag} */,
  {32'hc57d0104, 32'h00000000} /* (24, 24, 9) {real, imag} */,
  {32'hc5b01b46, 32'h00000000} /* (24, 24, 8) {real, imag} */,
  {32'hc5b022ea, 32'h00000000} /* (24, 24, 7) {real, imag} */,
  {32'hc5b36a16, 32'h00000000} /* (24, 24, 6) {real, imag} */,
  {32'hc5c84e05, 32'h00000000} /* (24, 24, 5) {real, imag} */,
  {32'hc5d7a9e4, 32'h00000000} /* (24, 24, 4) {real, imag} */,
  {32'hc60649c8, 32'h00000000} /* (24, 24, 3) {real, imag} */,
  {32'hc5ef8105, 32'h00000000} /* (24, 24, 2) {real, imag} */,
  {32'hc5e48896, 32'h00000000} /* (24, 24, 1) {real, imag} */,
  {32'hc5ec664b, 32'h00000000} /* (24, 24, 0) {real, imag} */,
  {32'hc5b198e6, 32'h00000000} /* (24, 23, 31) {real, imag} */,
  {32'hc5c53f18, 32'h00000000} /* (24, 23, 30) {real, imag} */,
  {32'hc5d39988, 32'h00000000} /* (24, 23, 29) {real, imag} */,
  {32'hc5c563e4, 32'h00000000} /* (24, 23, 28) {real, imag} */,
  {32'hc5d6469e, 32'h00000000} /* (24, 23, 27) {real, imag} */,
  {32'hc5cd91d6, 32'h00000000} /* (24, 23, 26) {real, imag} */,
  {32'hc5ae73bc, 32'h00000000} /* (24, 23, 25) {real, imag} */,
  {32'hc5a9bb1f, 32'h00000000} /* (24, 23, 24) {real, imag} */,
  {32'hc59d918d, 32'h00000000} /* (24, 23, 23) {real, imag} */,
  {32'hc5870e4d, 32'h00000000} /* (24, 23, 22) {real, imag} */,
  {32'hc4ca8f90, 32'h00000000} /* (24, 23, 21) {real, imag} */,
  {32'h447dd61c, 32'h00000000} /* (24, 23, 20) {real, imag} */,
  {32'h450192a4, 32'h00000000} /* (24, 23, 19) {real, imag} */,
  {32'h456de716, 32'h00000000} /* (24, 23, 18) {real, imag} */,
  {32'h4581632c, 32'h00000000} /* (24, 23, 17) {real, imag} */,
  {32'h457800e6, 32'h00000000} /* (24, 23, 16) {real, imag} */,
  {32'h458cedba, 32'h00000000} /* (24, 23, 15) {real, imag} */,
  {32'h45a2596a, 32'h00000000} /* (24, 23, 14) {real, imag} */,
  {32'h4556ed07, 32'h00000000} /* (24, 23, 13) {real, imag} */,
  {32'h45124193, 32'h00000000} /* (24, 23, 12) {real, imag} */,
  {32'h44441804, 32'h00000000} /* (24, 23, 11) {real, imag} */,
  {32'hc4d71aba, 32'h00000000} /* (24, 23, 10) {real, imag} */,
  {32'hc53c9c01, 32'h00000000} /* (24, 23, 9) {real, imag} */,
  {32'hc58e422f, 32'h00000000} /* (24, 23, 8) {real, imag} */,
  {32'hc5a9bb97, 32'h00000000} /* (24, 23, 7) {real, imag} */,
  {32'hc5a1fdff, 32'h00000000} /* (24, 23, 6) {real, imag} */,
  {32'hc5cccbab, 32'h00000000} /* (24, 23, 5) {real, imag} */,
  {32'hc5b0efac, 32'h00000000} /* (24, 23, 4) {real, imag} */,
  {32'hc5a88a39, 32'h00000000} /* (24, 23, 3) {real, imag} */,
  {32'hc5d0823f, 32'h00000000} /* (24, 23, 2) {real, imag} */,
  {32'hc5e62eb2, 32'h00000000} /* (24, 23, 1) {real, imag} */,
  {32'hc5bf6c49, 32'h00000000} /* (24, 23, 0) {real, imag} */,
  {32'hc596f9be, 32'h00000000} /* (24, 22, 31) {real, imag} */,
  {32'hc59399e7, 32'h00000000} /* (24, 22, 30) {real, imag} */,
  {32'hc5b68eac, 32'h00000000} /* (24, 22, 29) {real, imag} */,
  {32'hc5a8b366, 32'h00000000} /* (24, 22, 28) {real, imag} */,
  {32'hc5a41e2c, 32'h00000000} /* (24, 22, 27) {real, imag} */,
  {32'hc599bdd8, 32'h00000000} /* (24, 22, 26) {real, imag} */,
  {32'hc572a7c8, 32'h00000000} /* (24, 22, 25) {real, imag} */,
  {32'hc57f2559, 32'h00000000} /* (24, 22, 24) {real, imag} */,
  {32'hc57524b0, 32'h00000000} /* (24, 22, 23) {real, imag} */,
  {32'hc5691e34, 32'h00000000} /* (24, 22, 22) {real, imag} */,
  {32'hc4345436, 32'h00000000} /* (24, 22, 21) {real, imag} */,
  {32'h44a4b74c, 32'h00000000} /* (24, 22, 20) {real, imag} */,
  {32'h45646fd2, 32'h00000000} /* (24, 22, 19) {real, imag} */,
  {32'h454eeca6, 32'h00000000} /* (24, 22, 18) {real, imag} */,
  {32'h45510d77, 32'h00000000} /* (24, 22, 17) {real, imag} */,
  {32'h4541b935, 32'h00000000} /* (24, 22, 16) {real, imag} */,
  {32'h45508031, 32'h00000000} /* (24, 22, 15) {real, imag} */,
  {32'h456f4c1a, 32'h00000000} /* (24, 22, 14) {real, imag} */,
  {32'h4569ad1c, 32'h00000000} /* (24, 22, 13) {real, imag} */,
  {32'h451c3468, 32'h00000000} /* (24, 22, 12) {real, imag} */,
  {32'h44670ca0, 32'h00000000} /* (24, 22, 11) {real, imag} */,
  {32'hc48cf7c7, 32'h00000000} /* (24, 22, 10) {real, imag} */,
  {32'hc53cfa96, 32'h00000000} /* (24, 22, 9) {real, imag} */,
  {32'hc55cd779, 32'h00000000} /* (24, 22, 8) {real, imag} */,
  {32'hc58c2466, 32'h00000000} /* (24, 22, 7) {real, imag} */,
  {32'hc5880c46, 32'h00000000} /* (24, 22, 6) {real, imag} */,
  {32'hc58d2ad7, 32'h00000000} /* (24, 22, 5) {real, imag} */,
  {32'hc5885757, 32'h00000000} /* (24, 22, 4) {real, imag} */,
  {32'hc588628f, 32'h00000000} /* (24, 22, 3) {real, imag} */,
  {32'hc58c7660, 32'h00000000} /* (24, 22, 2) {real, imag} */,
  {32'hc5996efa, 32'h00000000} /* (24, 22, 1) {real, imag} */,
  {32'hc597fb90, 32'h00000000} /* (24, 22, 0) {real, imag} */,
  {32'hc4d77892, 32'h00000000} /* (24, 21, 31) {real, imag} */,
  {32'hc4f5343b, 32'h00000000} /* (24, 21, 30) {real, imag} */,
  {32'hc542e068, 32'h00000000} /* (24, 21, 29) {real, imag} */,
  {32'hc50cf0bf, 32'h00000000} /* (24, 21, 28) {real, imag} */,
  {32'hc4d1d5af, 32'h00000000} /* (24, 21, 27) {real, imag} */,
  {32'hc4e9801e, 32'h00000000} /* (24, 21, 26) {real, imag} */,
  {32'hc4f34862, 32'h00000000} /* (24, 21, 25) {real, imag} */,
  {32'hc4e7e47c, 32'h00000000} /* (24, 21, 24) {real, imag} */,
  {32'hc4af5e9d, 32'h00000000} /* (24, 21, 23) {real, imag} */,
  {32'hc3f5cff0, 32'h00000000} /* (24, 21, 22) {real, imag} */,
  {32'hc40b3359, 32'h00000000} /* (24, 21, 21) {real, imag} */,
  {32'hc3b9366c, 32'h00000000} /* (24, 21, 20) {real, imag} */,
  {32'h448416a6, 32'h00000000} /* (24, 21, 19) {real, imag} */,
  {32'h44943d5e, 32'h00000000} /* (24, 21, 18) {real, imag} */,
  {32'h448b098d, 32'h00000000} /* (24, 21, 17) {real, imag} */,
  {32'h45095480, 32'h00000000} /* (24, 21, 16) {real, imag} */,
  {32'h448ded4a, 32'h00000000} /* (24, 21, 15) {real, imag} */,
  {32'h44d15419, 32'h00000000} /* (24, 21, 14) {real, imag} */,
  {32'h4512ee72, 32'h00000000} /* (24, 21, 13) {real, imag} */,
  {32'h44d032e8, 32'h00000000} /* (24, 21, 12) {real, imag} */,
  {32'hc3c24d4c, 32'h00000000} /* (24, 21, 11) {real, imag} */,
  {32'hc457ead4, 32'h00000000} /* (24, 21, 10) {real, imag} */,
  {32'hc4647dd8, 32'h00000000} /* (24, 21, 9) {real, imag} */,
  {32'hc49cda5a, 32'h00000000} /* (24, 21, 8) {real, imag} */,
  {32'hc4ca789f, 32'h00000000} /* (24, 21, 7) {real, imag} */,
  {32'hc4fe287a, 32'h00000000} /* (24, 21, 6) {real, imag} */,
  {32'hc4e4a194, 32'h00000000} /* (24, 21, 5) {real, imag} */,
  {32'hc5326ca0, 32'h00000000} /* (24, 21, 4) {real, imag} */,
  {32'hc529f019, 32'h00000000} /* (24, 21, 3) {real, imag} */,
  {32'hc4a450c6, 32'h00000000} /* (24, 21, 2) {real, imag} */,
  {32'hc48f590d, 32'h00000000} /* (24, 21, 1) {real, imag} */,
  {32'hc4d42fdb, 32'h00000000} /* (24, 21, 0) {real, imag} */,
  {32'h449ea2fd, 32'h00000000} /* (24, 20, 31) {real, imag} */,
  {32'h4496e580, 32'h00000000} /* (24, 20, 30) {real, imag} */,
  {32'h44881880, 32'h00000000} /* (24, 20, 29) {real, imag} */,
  {32'h44251251, 32'h00000000} /* (24, 20, 28) {real, imag} */,
  {32'h44a609b4, 32'h00000000} /* (24, 20, 27) {real, imag} */,
  {32'h451d5c30, 32'h00000000} /* (24, 20, 26) {real, imag} */,
  {32'h4486c28e, 32'h00000000} /* (24, 20, 25) {real, imag} */,
  {32'h4488898b, 32'h00000000} /* (24, 20, 24) {real, imag} */,
  {32'h451c9d90, 32'h00000000} /* (24, 20, 23) {real, imag} */,
  {32'h450dc2c7, 32'h00000000} /* (24, 20, 22) {real, imag} */,
  {32'h446bd429, 32'h00000000} /* (24, 20, 21) {real, imag} */,
  {32'hc4c9fbc2, 32'h00000000} /* (24, 20, 20) {real, imag} */,
  {32'hc4de7440, 32'h00000000} /* (24, 20, 19) {real, imag} */,
  {32'hc4a502ae, 32'h00000000} /* (24, 20, 18) {real, imag} */,
  {32'hc50d6723, 32'h00000000} /* (24, 20, 17) {real, imag} */,
  {32'hc4a4556f, 32'h00000000} /* (24, 20, 16) {real, imag} */,
  {32'hc4c0856b, 32'h00000000} /* (24, 20, 15) {real, imag} */,
  {32'hc49755a0, 32'h00000000} /* (24, 20, 14) {real, imag} */,
  {32'hc4a53f06, 32'h00000000} /* (24, 20, 13) {real, imag} */,
  {32'hc40ac21d, 32'h00000000} /* (24, 20, 12) {real, imag} */,
  {32'hc4b6a2aa, 32'h00000000} /* (24, 20, 11) {real, imag} */,
  {32'hc4489088, 32'h00000000} /* (24, 20, 10) {real, imag} */,
  {32'h44b5360c, 32'h00000000} /* (24, 20, 9) {real, imag} */,
  {32'h43f9a89c, 32'h00000000} /* (24, 20, 8) {real, imag} */,
  {32'h445bd98e, 32'h00000000} /* (24, 20, 7) {real, imag} */,
  {32'h44836da4, 32'h00000000} /* (24, 20, 6) {real, imag} */,
  {32'h447867b3, 32'h00000000} /* (24, 20, 5) {real, imag} */,
  {32'h44aa8d0e, 32'h00000000} /* (24, 20, 4) {real, imag} */,
  {32'h442d1375, 32'h00000000} /* (24, 20, 3) {real, imag} */,
  {32'h44989e8c, 32'h00000000} /* (24, 20, 2) {real, imag} */,
  {32'h44c1d40b, 32'h00000000} /* (24, 20, 1) {real, imag} */,
  {32'h449da7b3, 32'h00000000} /* (24, 20, 0) {real, imag} */,
  {32'h452ab8ce, 32'h00000000} /* (24, 19, 31) {real, imag} */,
  {32'h45532302, 32'h00000000} /* (24, 19, 30) {real, imag} */,
  {32'h454b5f89, 32'h00000000} /* (24, 19, 29) {real, imag} */,
  {32'h4527a7ba, 32'h00000000} /* (24, 19, 28) {real, imag} */,
  {32'h45488bd2, 32'h00000000} /* (24, 19, 27) {real, imag} */,
  {32'h45751662, 32'h00000000} /* (24, 19, 26) {real, imag} */,
  {32'h45329cc8, 32'h00000000} /* (24, 19, 25) {real, imag} */,
  {32'h453e5189, 32'h00000000} /* (24, 19, 24) {real, imag} */,
  {32'h454edf38, 32'h00000000} /* (24, 19, 23) {real, imag} */,
  {32'h451525aa, 32'h00000000} /* (24, 19, 22) {real, imag} */,
  {32'h44aa9e66, 32'h00000000} /* (24, 19, 21) {real, imag} */,
  {32'hc4d182e8, 32'h00000000} /* (24, 19, 20) {real, imag} */,
  {32'hc527e005, 32'h00000000} /* (24, 19, 19) {real, imag} */,
  {32'hc55b5466, 32'h00000000} /* (24, 19, 18) {real, imag} */,
  {32'hc54c2d3a, 32'h00000000} /* (24, 19, 17) {real, imag} */,
  {32'hc54f48dd, 32'h00000000} /* (24, 19, 16) {real, imag} */,
  {32'hc534cf2e, 32'h00000000} /* (24, 19, 15) {real, imag} */,
  {32'hc50e5cbe, 32'h00000000} /* (24, 19, 14) {real, imag} */,
  {32'hc5208165, 32'h00000000} /* (24, 19, 13) {real, imag} */,
  {32'hc526c38a, 32'h00000000} /* (24, 19, 12) {real, imag} */,
  {32'hc4c05aa5, 32'h00000000} /* (24, 19, 11) {real, imag} */,
  {32'h448b0a4c, 32'h00000000} /* (24, 19, 10) {real, imag} */,
  {32'h44feb28c, 32'h00000000} /* (24, 19, 9) {real, imag} */,
  {32'h45139f03, 32'h00000000} /* (24, 19, 8) {real, imag} */,
  {32'h45278444, 32'h00000000} /* (24, 19, 7) {real, imag} */,
  {32'h4563da1a, 32'h00000000} /* (24, 19, 6) {real, imag} */,
  {32'h454aa7f9, 32'h00000000} /* (24, 19, 5) {real, imag} */,
  {32'h453807ca, 32'h00000000} /* (24, 19, 4) {real, imag} */,
  {32'h4518b6b7, 32'h00000000} /* (24, 19, 3) {real, imag} */,
  {32'h45410952, 32'h00000000} /* (24, 19, 2) {real, imag} */,
  {32'h454e25ac, 32'h00000000} /* (24, 19, 1) {real, imag} */,
  {32'h4521fc61, 32'h00000000} /* (24, 19, 0) {real, imag} */,
  {32'h4599f38a, 32'h00000000} /* (24, 18, 31) {real, imag} */,
  {32'h45a345b9, 32'h00000000} /* (24, 18, 30) {real, imag} */,
  {32'h459d3808, 32'h00000000} /* (24, 18, 29) {real, imag} */,
  {32'h4590cac1, 32'h00000000} /* (24, 18, 28) {real, imag} */,
  {32'h456ee022, 32'h00000000} /* (24, 18, 27) {real, imag} */,
  {32'h456f6122, 32'h00000000} /* (24, 18, 26) {real, imag} */,
  {32'h45953e5f, 32'h00000000} /* (24, 18, 25) {real, imag} */,
  {32'h45819497, 32'h00000000} /* (24, 18, 24) {real, imag} */,
  {32'h45281d8b, 32'h00000000} /* (24, 18, 23) {real, imag} */,
  {32'h4539cb1c, 32'h00000000} /* (24, 18, 22) {real, imag} */,
  {32'h4509ca5a, 32'h00000000} /* (24, 18, 21) {real, imag} */,
  {32'hc50dab80, 32'h00000000} /* (24, 18, 20) {real, imag} */,
  {32'hc5577ad4, 32'h00000000} /* (24, 18, 19) {real, imag} */,
  {32'hc572d365, 32'h00000000} /* (24, 18, 18) {real, imag} */,
  {32'hc5980aee, 32'h00000000} /* (24, 18, 17) {real, imag} */,
  {32'hc53b09a6, 32'h00000000} /* (24, 18, 16) {real, imag} */,
  {32'hc560b7b0, 32'h00000000} /* (24, 18, 15) {real, imag} */,
  {32'hc57cd912, 32'h00000000} /* (24, 18, 14) {real, imag} */,
  {32'hc53bc9ec, 32'h00000000} /* (24, 18, 13) {real, imag} */,
  {32'hc5210f16, 32'h00000000} /* (24, 18, 12) {real, imag} */,
  {32'hc4dda4c1, 32'h00000000} /* (24, 18, 11) {real, imag} */,
  {32'h44c657e9, 32'h00000000} /* (24, 18, 10) {real, imag} */,
  {32'h451dc502, 32'h00000000} /* (24, 18, 9) {real, imag} */,
  {32'h4534562a, 32'h00000000} /* (24, 18, 8) {real, imag} */,
  {32'h45645cfd, 32'h00000000} /* (24, 18, 7) {real, imag} */,
  {32'h457a0688, 32'h00000000} /* (24, 18, 6) {real, imag} */,
  {32'h45849211, 32'h00000000} /* (24, 18, 5) {real, imag} */,
  {32'h455fb1f8, 32'h00000000} /* (24, 18, 4) {real, imag} */,
  {32'h45813712, 32'h00000000} /* (24, 18, 3) {real, imag} */,
  {32'h458082b6, 32'h00000000} /* (24, 18, 2) {real, imag} */,
  {32'h4598adf8, 32'h00000000} /* (24, 18, 1) {real, imag} */,
  {32'h458ee834, 32'h00000000} /* (24, 18, 0) {real, imag} */,
  {32'h45aa80de, 32'h00000000} /* (24, 17, 31) {real, imag} */,
  {32'h45b1b401, 32'h00000000} /* (24, 17, 30) {real, imag} */,
  {32'h45a7d3a4, 32'h00000000} /* (24, 17, 29) {real, imag} */,
  {32'h45a6bdbb, 32'h00000000} /* (24, 17, 28) {real, imag} */,
  {32'h45b3d889, 32'h00000000} /* (24, 17, 27) {real, imag} */,
  {32'h458d0dfd, 32'h00000000} /* (24, 17, 26) {real, imag} */,
  {32'h45980fd4, 32'h00000000} /* (24, 17, 25) {real, imag} */,
  {32'h4592be2a, 32'h00000000} /* (24, 17, 24) {real, imag} */,
  {32'h45882505, 32'h00000000} /* (24, 17, 23) {real, imag} */,
  {32'h451ab3c3, 32'h00000000} /* (24, 17, 22) {real, imag} */,
  {32'h4459d778, 32'h00000000} /* (24, 17, 21) {real, imag} */,
  {32'hc4e02446, 32'h00000000} /* (24, 17, 20) {real, imag} */,
  {32'hc56526b8, 32'h00000000} /* (24, 17, 19) {real, imag} */,
  {32'hc5746953, 32'h00000000} /* (24, 17, 18) {real, imag} */,
  {32'hc5971bc4, 32'h00000000} /* (24, 17, 17) {real, imag} */,
  {32'hc58b651c, 32'h00000000} /* (24, 17, 16) {real, imag} */,
  {32'hc59b40a6, 32'h00000000} /* (24, 17, 15) {real, imag} */,
  {32'hc59b409f, 32'h00000000} /* (24, 17, 14) {real, imag} */,
  {32'hc5843f76, 32'h00000000} /* (24, 17, 13) {real, imag} */,
  {32'hc54ef256, 32'h00000000} /* (24, 17, 12) {real, imag} */,
  {32'hc4f3df0c, 32'h00000000} /* (24, 17, 11) {real, imag} */,
  {32'h42918600, 32'h00000000} /* (24, 17, 10) {real, imag} */,
  {32'h45104f8f, 32'h00000000} /* (24, 17, 9) {real, imag} */,
  {32'h452b479e, 32'h00000000} /* (24, 17, 8) {real, imag} */,
  {32'h457ed1aa, 32'h00000000} /* (24, 17, 7) {real, imag} */,
  {32'h45932e9e, 32'h00000000} /* (24, 17, 6) {real, imag} */,
  {32'h4594d1f7, 32'h00000000} /* (24, 17, 5) {real, imag} */,
  {32'h45a2afbc, 32'h00000000} /* (24, 17, 4) {real, imag} */,
  {32'h45a84e92, 32'h00000000} /* (24, 17, 3) {real, imag} */,
  {32'h459fc418, 32'h00000000} /* (24, 17, 2) {real, imag} */,
  {32'h45bef92a, 32'h00000000} /* (24, 17, 1) {real, imag} */,
  {32'h45ce2fb6, 32'h00000000} /* (24, 17, 0) {real, imag} */,
  {32'h45b4537c, 32'h00000000} /* (24, 16, 31) {real, imag} */,
  {32'h45cd757a, 32'h00000000} /* (24, 16, 30) {real, imag} */,
  {32'h45bad576, 32'h00000000} /* (24, 16, 29) {real, imag} */,
  {32'h45a35d3a, 32'h00000000} /* (24, 16, 28) {real, imag} */,
  {32'h45a02b42, 32'h00000000} /* (24, 16, 27) {real, imag} */,
  {32'h4593a633, 32'h00000000} /* (24, 16, 26) {real, imag} */,
  {32'h459135a6, 32'h00000000} /* (24, 16, 25) {real, imag} */,
  {32'h45a450ae, 32'h00000000} /* (24, 16, 24) {real, imag} */,
  {32'h4586a27d, 32'h00000000} /* (24, 16, 23) {real, imag} */,
  {32'h4541110c, 32'h00000000} /* (24, 16, 22) {real, imag} */,
  {32'h4446bd5c, 32'h00000000} /* (24, 16, 21) {real, imag} */,
  {32'hc538bc05, 32'h00000000} /* (24, 16, 20) {real, imag} */,
  {32'hc58ecf6d, 32'h00000000} /* (24, 16, 19) {real, imag} */,
  {32'hc579bf1c, 32'h00000000} /* (24, 16, 18) {real, imag} */,
  {32'hc586e361, 32'h00000000} /* (24, 16, 17) {real, imag} */,
  {32'hc5a2fe94, 32'h00000000} /* (24, 16, 16) {real, imag} */,
  {32'hc5974b3c, 32'h00000000} /* (24, 16, 15) {real, imag} */,
  {32'hc59e64a4, 32'h00000000} /* (24, 16, 14) {real, imag} */,
  {32'hc597e892, 32'h00000000} /* (24, 16, 13) {real, imag} */,
  {32'hc59268bc, 32'h00000000} /* (24, 16, 12) {real, imag} */,
  {32'hc50ec9c1, 32'h00000000} /* (24, 16, 11) {real, imag} */,
  {32'h43e208d0, 32'h00000000} /* (24, 16, 10) {real, imag} */,
  {32'h45211554, 32'h00000000} /* (24, 16, 9) {real, imag} */,
  {32'h454f09e4, 32'h00000000} /* (24, 16, 8) {real, imag} */,
  {32'h459ef6d3, 32'h00000000} /* (24, 16, 7) {real, imag} */,
  {32'h45a86f7e, 32'h00000000} /* (24, 16, 6) {real, imag} */,
  {32'h45c78efe, 32'h00000000} /* (24, 16, 5) {real, imag} */,
  {32'h45cc2c4e, 32'h00000000} /* (24, 16, 4) {real, imag} */,
  {32'h45b7290f, 32'h00000000} /* (24, 16, 3) {real, imag} */,
  {32'h45c3f54c, 32'h00000000} /* (24, 16, 2) {real, imag} */,
  {32'h45cec649, 32'h00000000} /* (24, 16, 1) {real, imag} */,
  {32'h45c2e4bc, 32'h00000000} /* (24, 16, 0) {real, imag} */,
  {32'h45a8bc28, 32'h00000000} /* (24, 15, 31) {real, imag} */,
  {32'h45bdf3b3, 32'h00000000} /* (24, 15, 30) {real, imag} */,
  {32'h45b39d02, 32'h00000000} /* (24, 15, 29) {real, imag} */,
  {32'h45b6460e, 32'h00000000} /* (24, 15, 28) {real, imag} */,
  {32'h45aab668, 32'h00000000} /* (24, 15, 27) {real, imag} */,
  {32'h45998282, 32'h00000000} /* (24, 15, 26) {real, imag} */,
  {32'h458e7981, 32'h00000000} /* (24, 15, 25) {real, imag} */,
  {32'h4583aa6c, 32'h00000000} /* (24, 15, 24) {real, imag} */,
  {32'h457f83c9, 32'h00000000} /* (24, 15, 23) {real, imag} */,
  {32'h44f7603a, 32'h00000000} /* (24, 15, 22) {real, imag} */,
  {32'h4327fbb0, 32'h00000000} /* (24, 15, 21) {real, imag} */,
  {32'hc5037cbe, 32'h00000000} /* (24, 15, 20) {real, imag} */,
  {32'hc58569bf, 32'h00000000} /* (24, 15, 19) {real, imag} */,
  {32'hc57292b4, 32'h00000000} /* (24, 15, 18) {real, imag} */,
  {32'hc58b2804, 32'h00000000} /* (24, 15, 17) {real, imag} */,
  {32'hc5a41b12, 32'h00000000} /* (24, 15, 16) {real, imag} */,
  {32'hc595e61a, 32'h00000000} /* (24, 15, 15) {real, imag} */,
  {32'hc5aa6571, 32'h00000000} /* (24, 15, 14) {real, imag} */,
  {32'hc5893480, 32'h00000000} /* (24, 15, 13) {real, imag} */,
  {32'hc574c348, 32'h00000000} /* (24, 15, 12) {real, imag} */,
  {32'hc4f9012c, 32'h00000000} /* (24, 15, 11) {real, imag} */,
  {32'h4461a12e, 32'h00000000} /* (24, 15, 10) {real, imag} */,
  {32'h45059ad6, 32'h00000000} /* (24, 15, 9) {real, imag} */,
  {32'h45609d51, 32'h00000000} /* (24, 15, 8) {real, imag} */,
  {32'h4595da14, 32'h00000000} /* (24, 15, 7) {real, imag} */,
  {32'h45aaad4c, 32'h00000000} /* (24, 15, 6) {real, imag} */,
  {32'h45b9080a, 32'h00000000} /* (24, 15, 5) {real, imag} */,
  {32'h45b14bbd, 32'h00000000} /* (24, 15, 4) {real, imag} */,
  {32'h45cf683f, 32'h00000000} /* (24, 15, 3) {real, imag} */,
  {32'h45c8aca6, 32'h00000000} /* (24, 15, 2) {real, imag} */,
  {32'h45b86b5e, 32'h00000000} /* (24, 15, 1) {real, imag} */,
  {32'h45aca4bc, 32'h00000000} /* (24, 15, 0) {real, imag} */,
  {32'h45a31358, 32'h00000000} /* (24, 14, 31) {real, imag} */,
  {32'h45a2fd13, 32'h00000000} /* (24, 14, 30) {real, imag} */,
  {32'h459febec, 32'h00000000} /* (24, 14, 29) {real, imag} */,
  {32'h45aaad68, 32'h00000000} /* (24, 14, 28) {real, imag} */,
  {32'h45a2cb1d, 32'h00000000} /* (24, 14, 27) {real, imag} */,
  {32'h45a6e2ad, 32'h00000000} /* (24, 14, 26) {real, imag} */,
  {32'h458f9c55, 32'h00000000} /* (24, 14, 25) {real, imag} */,
  {32'h458a0fe1, 32'h00000000} /* (24, 14, 24) {real, imag} */,
  {32'h459b21dd, 32'h00000000} /* (24, 14, 23) {real, imag} */,
  {32'h45371ba2, 32'h00000000} /* (24, 14, 22) {real, imag} */,
  {32'h4310fd70, 32'h00000000} /* (24, 14, 21) {real, imag} */,
  {32'hc4ffc5be, 32'h00000000} /* (24, 14, 20) {real, imag} */,
  {32'hc585cb98, 32'h00000000} /* (24, 14, 19) {real, imag} */,
  {32'hc5872aa0, 32'h00000000} /* (24, 14, 18) {real, imag} */,
  {32'hc5a9af91, 32'h00000000} /* (24, 14, 17) {real, imag} */,
  {32'hc5adcca7, 32'h00000000} /* (24, 14, 16) {real, imag} */,
  {32'hc596a12c, 32'h00000000} /* (24, 14, 15) {real, imag} */,
  {32'hc589c76b, 32'h00000000} /* (24, 14, 14) {real, imag} */,
  {32'hc586ca0c, 32'h00000000} /* (24, 14, 13) {real, imag} */,
  {32'hc540d99f, 32'h00000000} /* (24, 14, 12) {real, imag} */,
  {32'hc4e3a5c8, 32'h00000000} /* (24, 14, 11) {real, imag} */,
  {32'h44021078, 32'h00000000} /* (24, 14, 10) {real, imag} */,
  {32'h4531ab4e, 32'h00000000} /* (24, 14, 9) {real, imag} */,
  {32'h45904e4b, 32'h00000000} /* (24, 14, 8) {real, imag} */,
  {32'h45959aa7, 32'h00000000} /* (24, 14, 7) {real, imag} */,
  {32'h45ab57f3, 32'h00000000} /* (24, 14, 6) {real, imag} */,
  {32'h45c9417a, 32'h00000000} /* (24, 14, 5) {real, imag} */,
  {32'h45c9e386, 32'h00000000} /* (24, 14, 4) {real, imag} */,
  {32'h45b6b08a, 32'h00000000} /* (24, 14, 3) {real, imag} */,
  {32'h45ab8f68, 32'h00000000} /* (24, 14, 2) {real, imag} */,
  {32'h45a24b1b, 32'h00000000} /* (24, 14, 1) {real, imag} */,
  {32'h459eb95b, 32'h00000000} /* (24, 14, 0) {real, imag} */,
  {32'h45871aa4, 32'h00000000} /* (24, 13, 31) {real, imag} */,
  {32'h458a1b34, 32'h00000000} /* (24, 13, 30) {real, imag} */,
  {32'h45900f40, 32'h00000000} /* (24, 13, 29) {real, imag} */,
  {32'h45abcd63, 32'h00000000} /* (24, 13, 28) {real, imag} */,
  {32'h459c7f24, 32'h00000000} /* (24, 13, 27) {real, imag} */,
  {32'h458b244c, 32'h00000000} /* (24, 13, 26) {real, imag} */,
  {32'h4565f94b, 32'h00000000} /* (24, 13, 25) {real, imag} */,
  {32'h45873296, 32'h00000000} /* (24, 13, 24) {real, imag} */,
  {32'h458f8316, 32'h00000000} /* (24, 13, 23) {real, imag} */,
  {32'h44dc22d8, 32'h00000000} /* (24, 13, 22) {real, imag} */,
  {32'h43890748, 32'h00000000} /* (24, 13, 21) {real, imag} */,
  {32'hc5051e08, 32'h00000000} /* (24, 13, 20) {real, imag} */,
  {32'hc580e278, 32'h00000000} /* (24, 13, 19) {real, imag} */,
  {32'hc5a1ca17, 32'h00000000} /* (24, 13, 18) {real, imag} */,
  {32'hc58e6b7e, 32'h00000000} /* (24, 13, 17) {real, imag} */,
  {32'hc57fe5ae, 32'h00000000} /* (24, 13, 16) {real, imag} */,
  {32'hc585c3d2, 32'h00000000} /* (24, 13, 15) {real, imag} */,
  {32'hc57df1cd, 32'h00000000} /* (24, 13, 14) {real, imag} */,
  {32'hc563b864, 32'h00000000} /* (24, 13, 13) {real, imag} */,
  {32'hc52acb7e, 32'h00000000} /* (24, 13, 12) {real, imag} */,
  {32'hc4ed04e6, 32'h00000000} /* (24, 13, 11) {real, imag} */,
  {32'h4485822e, 32'h00000000} /* (24, 13, 10) {real, imag} */,
  {32'h4532ed01, 32'h00000000} /* (24, 13, 9) {real, imag} */,
  {32'h458b7ab0, 32'h00000000} /* (24, 13, 8) {real, imag} */,
  {32'h459bd232, 32'h00000000} /* (24, 13, 7) {real, imag} */,
  {32'h45a7a0dc, 32'h00000000} /* (24, 13, 6) {real, imag} */,
  {32'h45cc9c5a, 32'h00000000} /* (24, 13, 5) {real, imag} */,
  {32'h45b47b54, 32'h00000000} /* (24, 13, 4) {real, imag} */,
  {32'h45a33ac8, 32'h00000000} /* (24, 13, 3) {real, imag} */,
  {32'h4581f501, 32'h00000000} /* (24, 13, 2) {real, imag} */,
  {32'h4580d2d4, 32'h00000000} /* (24, 13, 1) {real, imag} */,
  {32'h4580e179, 32'h00000000} /* (24, 13, 0) {real, imag} */,
  {32'h45220f3b, 32'h00000000} /* (24, 12, 31) {real, imag} */,
  {32'h45467e96, 32'h00000000} /* (24, 12, 30) {real, imag} */,
  {32'h453aa49a, 32'h00000000} /* (24, 12, 29) {real, imag} */,
  {32'h45660866, 32'h00000000} /* (24, 12, 28) {real, imag} */,
  {32'h4580b2e0, 32'h00000000} /* (24, 12, 27) {real, imag} */,
  {32'h455d1ac8, 32'h00000000} /* (24, 12, 26) {real, imag} */,
  {32'h45495477, 32'h00000000} /* (24, 12, 25) {real, imag} */,
  {32'h454ed2ee, 32'h00000000} /* (24, 12, 24) {real, imag} */,
  {32'h451e52b0, 32'h00000000} /* (24, 12, 23) {real, imag} */,
  {32'h4445c048, 32'h00000000} /* (24, 12, 22) {real, imag} */,
  {32'hc3ab7760, 32'h00000000} /* (24, 12, 21) {real, imag} */,
  {32'hc509418e, 32'h00000000} /* (24, 12, 20) {real, imag} */,
  {32'hc582dd76, 32'h00000000} /* (24, 12, 19) {real, imag} */,
  {32'hc5a0fc64, 32'h00000000} /* (24, 12, 18) {real, imag} */,
  {32'hc59107ac, 32'h00000000} /* (24, 12, 17) {real, imag} */,
  {32'hc57f0746, 32'h00000000} /* (24, 12, 16) {real, imag} */,
  {32'hc5868106, 32'h00000000} /* (24, 12, 15) {real, imag} */,
  {32'hc51f7ae6, 32'h00000000} /* (24, 12, 14) {real, imag} */,
  {32'hc5219d1a, 32'h00000000} /* (24, 12, 13) {real, imag} */,
  {32'hc509bf94, 32'h00000000} /* (24, 12, 12) {real, imag} */,
  {32'hc4ce1515, 32'h00000000} /* (24, 12, 11) {real, imag} */,
  {32'h45149a0c, 32'h00000000} /* (24, 12, 10) {real, imag} */,
  {32'h4535b765, 32'h00000000} /* (24, 12, 9) {real, imag} */,
  {32'h458e8fa3, 32'h00000000} /* (24, 12, 8) {real, imag} */,
  {32'h4568f43a, 32'h00000000} /* (24, 12, 7) {real, imag} */,
  {32'h45930789, 32'h00000000} /* (24, 12, 6) {real, imag} */,
  {32'h4590a088, 32'h00000000} /* (24, 12, 5) {real, imag} */,
  {32'h456bec48, 32'h00000000} /* (24, 12, 4) {real, imag} */,
  {32'h457df7e8, 32'h00000000} /* (24, 12, 3) {real, imag} */,
  {32'h454b6928, 32'h00000000} /* (24, 12, 2) {real, imag} */,
  {32'h4579f018, 32'h00000000} /* (24, 12, 1) {real, imag} */,
  {32'h454b3d36, 32'h00000000} /* (24, 12, 0) {real, imag} */,
  {32'h44624cfc, 32'h00000000} /* (24, 11, 31) {real, imag} */,
  {32'h4508bf10, 32'h00000000} /* (24, 11, 30) {real, imag} */,
  {32'h442e482a, 32'h00000000} /* (24, 11, 29) {real, imag} */,
  {32'h44335a08, 32'h00000000} /* (24, 11, 28) {real, imag} */,
  {32'h44934dbe, 32'h00000000} /* (24, 11, 27) {real, imag} */,
  {32'h450227ab, 32'h00000000} /* (24, 11, 26) {real, imag} */,
  {32'h44df76d3, 32'h00000000} /* (24, 11, 25) {real, imag} */,
  {32'h44f61b40, 32'h00000000} /* (24, 11, 24) {real, imag} */,
  {32'h44cb509e, 32'h00000000} /* (24, 11, 23) {real, imag} */,
  {32'h44ca8c64, 32'h00000000} /* (24, 11, 22) {real, imag} */,
  {32'hc474cff6, 32'h00000000} /* (24, 11, 21) {real, imag} */,
  {32'hc51d6997, 32'h00000000} /* (24, 11, 20) {real, imag} */,
  {32'hc54435e0, 32'h00000000} /* (24, 11, 19) {real, imag} */,
  {32'hc53fcdc2, 32'h00000000} /* (24, 11, 18) {real, imag} */,
  {32'hc53b1f24, 32'h00000000} /* (24, 11, 17) {real, imag} */,
  {32'hc4ec44cc, 32'h00000000} /* (24, 11, 16) {real, imag} */,
  {32'hc5141ef1, 32'h00000000} /* (24, 11, 15) {real, imag} */,
  {32'hc495a3c5, 32'h00000000} /* (24, 11, 14) {real, imag} */,
  {32'hc482b2f5, 32'h00000000} /* (24, 11, 13) {real, imag} */,
  {32'hc426234e, 32'h00000000} /* (24, 11, 12) {real, imag} */,
  {32'h42b81978, 32'h00000000} /* (24, 11, 11) {real, imag} */,
  {32'h440f5dfb, 32'h00000000} /* (24, 11, 10) {real, imag} */,
  {32'h452f9342, 32'h00000000} /* (24, 11, 9) {real, imag} */,
  {32'h453d8dfc, 32'h00000000} /* (24, 11, 8) {real, imag} */,
  {32'h45806d60, 32'h00000000} /* (24, 11, 7) {real, imag} */,
  {32'h457c4e4c, 32'h00000000} /* (24, 11, 6) {real, imag} */,
  {32'h45176640, 32'h00000000} /* (24, 11, 5) {real, imag} */,
  {32'h44a8b69a, 32'h00000000} /* (24, 11, 4) {real, imag} */,
  {32'h44a1d9d5, 32'h00000000} /* (24, 11, 3) {real, imag} */,
  {32'h44d68068, 32'h00000000} /* (24, 11, 2) {real, imag} */,
  {32'h44a5e943, 32'h00000000} /* (24, 11, 1) {real, imag} */,
  {32'h448f480a, 32'h00000000} /* (24, 11, 0) {real, imag} */,
  {32'hc4a0d1d8, 32'h00000000} /* (24, 10, 31) {real, imag} */,
  {32'hc52cec06, 32'h00000000} /* (24, 10, 30) {real, imag} */,
  {32'hc4f77bf1, 32'h00000000} /* (24, 10, 29) {real, imag} */,
  {32'hc5089fda, 32'h00000000} /* (24, 10, 28) {real, imag} */,
  {32'hc507ec27, 32'h00000000} /* (24, 10, 27) {real, imag} */,
  {32'hc4f5c587, 32'h00000000} /* (24, 10, 26) {real, imag} */,
  {32'hc4ea7257, 32'h00000000} /* (24, 10, 25) {real, imag} */,
  {32'hc4bda5f2, 32'h00000000} /* (24, 10, 24) {real, imag} */,
  {32'hc4b18eea, 32'h00000000} /* (24, 10, 23) {real, imag} */,
  {32'hc4e5e73e, 32'h00000000} /* (24, 10, 22) {real, imag} */,
  {32'hc5082f22, 32'h00000000} /* (24, 10, 21) {real, imag} */,
  {32'hc4860af0, 32'h00000000} /* (24, 10, 20) {real, imag} */,
  {32'hc3da2658, 32'h00000000} /* (24, 10, 19) {real, imag} */,
  {32'hc4230309, 32'h00000000} /* (24, 10, 18) {real, imag} */,
  {32'h43911698, 32'h00000000} /* (24, 10, 17) {real, imag} */,
  {32'h44524da1, 32'h00000000} /* (24, 10, 16) {real, imag} */,
  {32'h44e10960, 32'h00000000} /* (24, 10, 15) {real, imag} */,
  {32'h44b9f0a7, 32'h00000000} /* (24, 10, 14) {real, imag} */,
  {32'h4491593d, 32'h00000000} /* (24, 10, 13) {real, imag} */,
  {32'h44b08737, 32'h00000000} /* (24, 10, 12) {real, imag} */,
  {32'h4452821c, 32'h00000000} /* (24, 10, 11) {real, imag} */,
  {32'h441798da, 32'h00000000} /* (24, 10, 10) {real, imag} */,
  {32'h441f4d16, 32'h00000000} /* (24, 10, 9) {real, imag} */,
  {32'h4302eb6c, 32'h00000000} /* (24, 10, 8) {real, imag} */,
  {32'h447cc745, 32'h00000000} /* (24, 10, 7) {real, imag} */,
  {32'h433b9250, 32'h00000000} /* (24, 10, 6) {real, imag} */,
  {32'h43ab5d6c, 32'h00000000} /* (24, 10, 5) {real, imag} */,
  {32'hc4948416, 32'h00000000} /* (24, 10, 4) {real, imag} */,
  {32'hc536da69, 32'h00000000} /* (24, 10, 3) {real, imag} */,
  {32'hc4ad5ac8, 32'h00000000} /* (24, 10, 2) {real, imag} */,
  {32'hc4e45cf6, 32'h00000000} /* (24, 10, 1) {real, imag} */,
  {32'hc50507bc, 32'h00000000} /* (24, 10, 0) {real, imag} */,
  {32'hc585b9c3, 32'h00000000} /* (24, 9, 31) {real, imag} */,
  {32'hc596c07e, 32'h00000000} /* (24, 9, 30) {real, imag} */,
  {32'hc59b146e, 32'h00000000} /* (24, 9, 29) {real, imag} */,
  {32'hc59daaee, 32'h00000000} /* (24, 9, 28) {real, imag} */,
  {32'hc5b3dcd4, 32'h00000000} /* (24, 9, 27) {real, imag} */,
  {32'hc5b25ede, 32'h00000000} /* (24, 9, 26) {real, imag} */,
  {32'hc588322e, 32'h00000000} /* (24, 9, 25) {real, imag} */,
  {32'hc5a040df, 32'h00000000} /* (24, 9, 24) {real, imag} */,
  {32'hc58bf7aa, 32'h00000000} /* (24, 9, 23) {real, imag} */,
  {32'hc532a176, 32'h00000000} /* (24, 9, 22) {real, imag} */,
  {32'hc51f08fd, 32'h00000000} /* (24, 9, 21) {real, imag} */,
  {32'hc49e2602, 32'h00000000} /* (24, 9, 20) {real, imag} */,
  {32'h43c1ca98, 32'h00000000} /* (24, 9, 19) {real, imag} */,
  {32'h445b2ec4, 32'h00000000} /* (24, 9, 18) {real, imag} */,
  {32'h44d4e21c, 32'h00000000} /* (24, 9, 17) {real, imag} */,
  {32'h452f439e, 32'h00000000} /* (24, 9, 16) {real, imag} */,
  {32'h451c0697, 32'h00000000} /* (24, 9, 15) {real, imag} */,
  {32'h455c98d0, 32'h00000000} /* (24, 9, 14) {real, imag} */,
  {32'h4527b4aa, 32'h00000000} /* (24, 9, 13) {real, imag} */,
  {32'h45369fba, 32'h00000000} /* (24, 9, 12) {real, imag} */,
  {32'h44e859c7, 32'h00000000} /* (24, 9, 11) {real, imag} */,
  {32'h4416a730, 32'h00000000} /* (24, 9, 10) {real, imag} */,
  {32'hc3f952d8, 32'h00000000} /* (24, 9, 9) {real, imag} */,
  {32'hc4ab10cf, 32'h00000000} /* (24, 9, 8) {real, imag} */,
  {32'hc4ac2a10, 32'h00000000} /* (24, 9, 7) {real, imag} */,
  {32'hc51b5cf6, 32'h00000000} /* (24, 9, 6) {real, imag} */,
  {32'hc5168173, 32'h00000000} /* (24, 9, 5) {real, imag} */,
  {32'hc52f6b09, 32'h00000000} /* (24, 9, 4) {real, imag} */,
  {32'hc5958a9a, 32'h00000000} /* (24, 9, 3) {real, imag} */,
  {32'hc589723c, 32'h00000000} /* (24, 9, 2) {real, imag} */,
  {32'hc58a8fb9, 32'h00000000} /* (24, 9, 1) {real, imag} */,
  {32'hc56e5dfc, 32'h00000000} /* (24, 9, 0) {real, imag} */,
  {32'hc5b6a34e, 32'h00000000} /* (24, 8, 31) {real, imag} */,
  {32'hc5ae379c, 32'h00000000} /* (24, 8, 30) {real, imag} */,
  {32'hc5e6456c, 32'h00000000} /* (24, 8, 29) {real, imag} */,
  {32'hc5e9ff33, 32'h00000000} /* (24, 8, 28) {real, imag} */,
  {32'hc5d7073c, 32'h00000000} /* (24, 8, 27) {real, imag} */,
  {32'hc5d649e8, 32'h00000000} /* (24, 8, 26) {real, imag} */,
  {32'hc5e039cb, 32'h00000000} /* (24, 8, 25) {real, imag} */,
  {32'hc5c63aba, 32'h00000000} /* (24, 8, 24) {real, imag} */,
  {32'hc5a39498, 32'h00000000} /* (24, 8, 23) {real, imag} */,
  {32'hc593c471, 32'h00000000} /* (24, 8, 22) {real, imag} */,
  {32'hc54370c3, 32'h00000000} /* (24, 8, 21) {real, imag} */,
  {32'hc49782a8, 32'h00000000} /* (24, 8, 20) {real, imag} */,
  {32'h425875c0, 32'h00000000} /* (24, 8, 19) {real, imag} */,
  {32'h449557c0, 32'h00000000} /* (24, 8, 18) {real, imag} */,
  {32'h45026aa8, 32'h00000000} /* (24, 8, 17) {real, imag} */,
  {32'h4556eb14, 32'h00000000} /* (24, 8, 16) {real, imag} */,
  {32'h456527bb, 32'h00000000} /* (24, 8, 15) {real, imag} */,
  {32'h454e9085, 32'h00000000} /* (24, 8, 14) {real, imag} */,
  {32'h45887fa8, 32'h00000000} /* (24, 8, 13) {real, imag} */,
  {32'h4580ddbd, 32'h00000000} /* (24, 8, 12) {real, imag} */,
  {32'h453b195d, 32'h00000000} /* (24, 8, 11) {real, imag} */,
  {32'h44569420, 32'h00000000} /* (24, 8, 10) {real, imag} */,
  {32'hc2f5d2c0, 32'h00000000} /* (24, 8, 9) {real, imag} */,
  {32'hc50cdc28, 32'h00000000} /* (24, 8, 8) {real, imag} */,
  {32'hc580ac30, 32'h00000000} /* (24, 8, 7) {real, imag} */,
  {32'hc588705f, 32'h00000000} /* (24, 8, 6) {real, imag} */,
  {32'hc56dbd2f, 32'h00000000} /* (24, 8, 5) {real, imag} */,
  {32'hc57c99c0, 32'h00000000} /* (24, 8, 4) {real, imag} */,
  {32'hc58ecdfa, 32'h00000000} /* (24, 8, 3) {real, imag} */,
  {32'hc5c5c514, 32'h00000000} /* (24, 8, 2) {real, imag} */,
  {32'hc5c5fc1e, 32'h00000000} /* (24, 8, 1) {real, imag} */,
  {32'hc59a7f7c, 32'h00000000} /* (24, 8, 0) {real, imag} */,
  {32'hc5d6d77f, 32'h00000000} /* (24, 7, 31) {real, imag} */,
  {32'hc5fe3b74, 32'h00000000} /* (24, 7, 30) {real, imag} */,
  {32'hc5fd0e73, 32'h00000000} /* (24, 7, 29) {real, imag} */,
  {32'hc6038490, 32'h00000000} /* (24, 7, 28) {real, imag} */,
  {32'hc605642f, 32'h00000000} /* (24, 7, 27) {real, imag} */,
  {32'hc5f915f1, 32'h00000000} /* (24, 7, 26) {real, imag} */,
  {32'hc5f976ca, 32'h00000000} /* (24, 7, 25) {real, imag} */,
  {32'hc60312d8, 32'h00000000} /* (24, 7, 24) {real, imag} */,
  {32'hc5d348f3, 32'h00000000} /* (24, 7, 23) {real, imag} */,
  {32'hc5b28b1c, 32'h00000000} /* (24, 7, 22) {real, imag} */,
  {32'hc569de80, 32'h00000000} /* (24, 7, 21) {real, imag} */,
  {32'hc21e0000, 32'h00000000} /* (24, 7, 20) {real, imag} */,
  {32'hc2a30ae0, 32'h00000000} /* (24, 7, 19) {real, imag} */,
  {32'h4375de00, 32'h00000000} /* (24, 7, 18) {real, imag} */,
  {32'h4509c826, 32'h00000000} /* (24, 7, 17) {real, imag} */,
  {32'h4541c9b6, 32'h00000000} /* (24, 7, 16) {real, imag} */,
  {32'h454d528a, 32'h00000000} /* (24, 7, 15) {real, imag} */,
  {32'h455f383f, 32'h00000000} /* (24, 7, 14) {real, imag} */,
  {32'h45855db5, 32'h00000000} /* (24, 7, 13) {real, imag} */,
  {32'h458afdeb, 32'h00000000} /* (24, 7, 12) {real, imag} */,
  {32'h4530ec3d, 32'h00000000} /* (24, 7, 11) {real, imag} */,
  {32'h449a486c, 32'h00000000} /* (24, 7, 10) {real, imag} */,
  {32'hc48741a0, 32'h00000000} /* (24, 7, 9) {real, imag} */,
  {32'hc51416b2, 32'h00000000} /* (24, 7, 8) {real, imag} */,
  {32'hc51df3f2, 32'h00000000} /* (24, 7, 7) {real, imag} */,
  {32'hc5777490, 32'h00000000} /* (24, 7, 6) {real, imag} */,
  {32'hc5992ea4, 32'h00000000} /* (24, 7, 5) {real, imag} */,
  {32'hc5a1df7c, 32'h00000000} /* (24, 7, 4) {real, imag} */,
  {32'hc5bef564, 32'h00000000} /* (24, 7, 3) {real, imag} */,
  {32'hc5cee940, 32'h00000000} /* (24, 7, 2) {real, imag} */,
  {32'hc5e1cc6b, 32'h00000000} /* (24, 7, 1) {real, imag} */,
  {32'hc5da76a1, 32'h00000000} /* (24, 7, 0) {real, imag} */,
  {32'hc5ee306d, 32'h00000000} /* (24, 6, 31) {real, imag} */,
  {32'hc60000bc, 32'h00000000} /* (24, 6, 30) {real, imag} */,
  {32'hc6151e75, 32'h00000000} /* (24, 6, 29) {real, imag} */,
  {32'hc61af69a, 32'h00000000} /* (24, 6, 28) {real, imag} */,
  {32'hc60c660b, 32'h00000000} /* (24, 6, 27) {real, imag} */,
  {32'hc61282ec, 32'h00000000} /* (24, 6, 26) {real, imag} */,
  {32'hc6093aa3, 32'h00000000} /* (24, 6, 25) {real, imag} */,
  {32'hc60c1a16, 32'h00000000} /* (24, 6, 24) {real, imag} */,
  {32'hc6062462, 32'h00000000} /* (24, 6, 23) {real, imag} */,
  {32'hc5de1d74, 32'h00000000} /* (24, 6, 22) {real, imag} */,
  {32'hc59d0386, 32'h00000000} /* (24, 6, 21) {real, imag} */,
  {32'hc50b77e8, 32'h00000000} /* (24, 6, 20) {real, imag} */,
  {32'hc4654be4, 32'h00000000} /* (24, 6, 19) {real, imag} */,
  {32'h444cfb04, 32'h00000000} /* (24, 6, 18) {real, imag} */,
  {32'h44c76902, 32'h00000000} /* (24, 6, 17) {real, imag} */,
  {32'h45162964, 32'h00000000} /* (24, 6, 16) {real, imag} */,
  {32'h45546f06, 32'h00000000} /* (24, 6, 15) {real, imag} */,
  {32'h458c5492, 32'h00000000} /* (24, 6, 14) {real, imag} */,
  {32'h4594bb9e, 32'h00000000} /* (24, 6, 13) {real, imag} */,
  {32'h45873dac, 32'h00000000} /* (24, 6, 12) {real, imag} */,
  {32'h4528873c, 32'h00000000} /* (24, 6, 11) {real, imag} */,
  {32'h446cfb20, 32'h00000000} /* (24, 6, 10) {real, imag} */,
  {32'hc2a16b80, 32'h00000000} /* (24, 6, 9) {real, imag} */,
  {32'hc507f3f5, 32'h00000000} /* (24, 6, 8) {real, imag} */,
  {32'hc53bf45c, 32'h00000000} /* (24, 6, 7) {real, imag} */,
  {32'hc5699c0f, 32'h00000000} /* (24, 6, 6) {real, imag} */,
  {32'hc5888d80, 32'h00000000} /* (24, 6, 5) {real, imag} */,
  {32'hc5a1f70e, 32'h00000000} /* (24, 6, 4) {real, imag} */,
  {32'hc5d0d384, 32'h00000000} /* (24, 6, 3) {real, imag} */,
  {32'hc5f20b0c, 32'h00000000} /* (24, 6, 2) {real, imag} */,
  {32'hc6032b9c, 32'h00000000} /* (24, 6, 1) {real, imag} */,
  {32'hc5f82370, 32'h00000000} /* (24, 6, 0) {real, imag} */,
  {32'hc609bc5c, 32'h00000000} /* (24, 5, 31) {real, imag} */,
  {32'hc617376f, 32'h00000000} /* (24, 5, 30) {real, imag} */,
  {32'hc6256fe6, 32'h00000000} /* (24, 5, 29) {real, imag} */,
  {32'hc6263f17, 32'h00000000} /* (24, 5, 28) {real, imag} */,
  {32'hc61fd7a0, 32'h00000000} /* (24, 5, 27) {real, imag} */,
  {32'hc6192e6e, 32'h00000000} /* (24, 5, 26) {real, imag} */,
  {32'hc61a7ae4, 32'h00000000} /* (24, 5, 25) {real, imag} */,
  {32'hc60891bc, 32'h00000000} /* (24, 5, 24) {real, imag} */,
  {32'hc600f88d, 32'h00000000} /* (24, 5, 23) {real, imag} */,
  {32'hc5d873a0, 32'h00000000} /* (24, 5, 22) {real, imag} */,
  {32'hc5cf3870, 32'h00000000} /* (24, 5, 21) {real, imag} */,
  {32'hc585cef9, 32'h00000000} /* (24, 5, 20) {real, imag} */,
  {32'hc52b7205, 32'h00000000} /* (24, 5, 19) {real, imag} */,
  {32'hc4f3f20e, 32'h00000000} /* (24, 5, 18) {real, imag} */,
  {32'hc45e4e64, 32'h00000000} /* (24, 5, 17) {real, imag} */,
  {32'h44e6a6b0, 32'h00000000} /* (24, 5, 16) {real, imag} */,
  {32'h4580e1b0, 32'h00000000} /* (24, 5, 15) {real, imag} */,
  {32'h45881864, 32'h00000000} /* (24, 5, 14) {real, imag} */,
  {32'h4595f6b2, 32'h00000000} /* (24, 5, 13) {real, imag} */,
  {32'h458d3888, 32'h00000000} /* (24, 5, 12) {real, imag} */,
  {32'h45738610, 32'h00000000} /* (24, 5, 11) {real, imag} */,
  {32'h455512e6, 32'h00000000} /* (24, 5, 10) {real, imag} */,
  {32'h44b927b4, 32'h00000000} /* (24, 5, 9) {real, imag} */,
  {32'h43cb6630, 32'h00000000} /* (24, 5, 8) {real, imag} */,
  {32'hc4814bd8, 32'h00000000} /* (24, 5, 7) {real, imag} */,
  {32'hc50e4edc, 32'h00000000} /* (24, 5, 6) {real, imag} */,
  {32'hc574fc29, 32'h00000000} /* (24, 5, 5) {real, imag} */,
  {32'hc5a7e751, 32'h00000000} /* (24, 5, 4) {real, imag} */,
  {32'hc5e72542, 32'h00000000} /* (24, 5, 3) {real, imag} */,
  {32'hc5e2a114, 32'h00000000} /* (24, 5, 2) {real, imag} */,
  {32'hc5fe3cac, 32'h00000000} /* (24, 5, 1) {real, imag} */,
  {32'hc607985b, 32'h00000000} /* (24, 5, 0) {real, imag} */,
  {32'hc612e79c, 32'h00000000} /* (24, 4, 31) {real, imag} */,
  {32'hc6263c56, 32'h00000000} /* (24, 4, 30) {real, imag} */,
  {32'hc62546ee, 32'h00000000} /* (24, 4, 29) {real, imag} */,
  {32'hc6293af3, 32'h00000000} /* (24, 4, 28) {real, imag} */,
  {32'hc62329f6, 32'h00000000} /* (24, 4, 27) {real, imag} */,
  {32'hc6270b4c, 32'h00000000} /* (24, 4, 26) {real, imag} */,
  {32'hc61cbcd8, 32'h00000000} /* (24, 4, 25) {real, imag} */,
  {32'hc6164e6a, 32'h00000000} /* (24, 4, 24) {real, imag} */,
  {32'hc606c7cc, 32'h00000000} /* (24, 4, 23) {real, imag} */,
  {32'hc5fa39fa, 32'h00000000} /* (24, 4, 22) {real, imag} */,
  {32'hc5e5dc96, 32'h00000000} /* (24, 4, 21) {real, imag} */,
  {32'hc5c26f2c, 32'h00000000} /* (24, 4, 20) {real, imag} */,
  {32'hc5918896, 32'h00000000} /* (24, 4, 19) {real, imag} */,
  {32'hc56481f9, 32'h00000000} /* (24, 4, 18) {real, imag} */,
  {32'hc5069b0e, 32'h00000000} /* (24, 4, 17) {real, imag} */,
  {32'hc2cdbec0, 32'h00000000} /* (24, 4, 16) {real, imag} */,
  {32'h4557d3e0, 32'h00000000} /* (24, 4, 15) {real, imag} */,
  {32'h457eba7a, 32'h00000000} /* (24, 4, 14) {real, imag} */,
  {32'h458111af, 32'h00000000} /* (24, 4, 13) {real, imag} */,
  {32'h4599730e, 32'h00000000} /* (24, 4, 12) {real, imag} */,
  {32'h4575c015, 32'h00000000} /* (24, 4, 11) {real, imag} */,
  {32'h457e0786, 32'h00000000} /* (24, 4, 10) {real, imag} */,
  {32'h455877fb, 32'h00000000} /* (24, 4, 9) {real, imag} */,
  {32'h450a9f12, 32'h00000000} /* (24, 4, 8) {real, imag} */,
  {32'h44664298, 32'h00000000} /* (24, 4, 7) {real, imag} */,
  {32'hc42e3ab4, 32'h00000000} /* (24, 4, 6) {real, imag} */,
  {32'hc562c130, 32'h00000000} /* (24, 4, 5) {real, imag} */,
  {32'hc5acfaec, 32'h00000000} /* (24, 4, 4) {real, imag} */,
  {32'hc5e35bd2, 32'h00000000} /* (24, 4, 3) {real, imag} */,
  {32'hc5fbd476, 32'h00000000} /* (24, 4, 2) {real, imag} */,
  {32'hc6089520, 32'h00000000} /* (24, 4, 1) {real, imag} */,
  {32'hc60650ba, 32'h00000000} /* (24, 4, 0) {real, imag} */,
  {32'hc612eb28, 32'h00000000} /* (24, 3, 31) {real, imag} */,
  {32'hc61b6556, 32'h00000000} /* (24, 3, 30) {real, imag} */,
  {32'hc62ea7ae, 32'h00000000} /* (24, 3, 29) {real, imag} */,
  {32'hc63c39be, 32'h00000000} /* (24, 3, 28) {real, imag} */,
  {32'hc6345c72, 32'h00000000} /* (24, 3, 27) {real, imag} */,
  {32'hc62347f5, 32'h00000000} /* (24, 3, 26) {real, imag} */,
  {32'hc617a412, 32'h00000000} /* (24, 3, 25) {real, imag} */,
  {32'hc61c70b6, 32'h00000000} /* (24, 3, 24) {real, imag} */,
  {32'hc605c2fc, 32'h00000000} /* (24, 3, 23) {real, imag} */,
  {32'hc6029912, 32'h00000000} /* (24, 3, 22) {real, imag} */,
  {32'hc5e3c9e8, 32'h00000000} /* (24, 3, 21) {real, imag} */,
  {32'hc5bbfdef, 32'h00000000} /* (24, 3, 20) {real, imag} */,
  {32'hc5912be5, 32'h00000000} /* (24, 3, 19) {real, imag} */,
  {32'hc54e250d, 32'h00000000} /* (24, 3, 18) {real, imag} */,
  {32'hc50ace88, 32'h00000000} /* (24, 3, 17) {real, imag} */,
  {32'hc3e11370, 32'h00000000} /* (24, 3, 16) {real, imag} */,
  {32'h451efdef, 32'h00000000} /* (24, 3, 15) {real, imag} */,
  {32'h458654ce, 32'h00000000} /* (24, 3, 14) {real, imag} */,
  {32'h45c0cd0f, 32'h00000000} /* (24, 3, 13) {real, imag} */,
  {32'h45b8efb4, 32'h00000000} /* (24, 3, 12) {real, imag} */,
  {32'h4582be20, 32'h00000000} /* (24, 3, 11) {real, imag} */,
  {32'h457ee1c4, 32'h00000000} /* (24, 3, 10) {real, imag} */,
  {32'h45652d98, 32'h00000000} /* (24, 3, 9) {real, imag} */,
  {32'h452db0a4, 32'h00000000} /* (24, 3, 8) {real, imag} */,
  {32'h4497f09e, 32'h00000000} /* (24, 3, 7) {real, imag} */,
  {32'hc40481c8, 32'h00000000} /* (24, 3, 6) {real, imag} */,
  {32'hc5638d5f, 32'h00000000} /* (24, 3, 5) {real, imag} */,
  {32'hc5c98871, 32'h00000000} /* (24, 3, 4) {real, imag} */,
  {32'hc5cf7ea7, 32'h00000000} /* (24, 3, 3) {real, imag} */,
  {32'hc600dfa1, 32'h00000000} /* (24, 3, 2) {real, imag} */,
  {32'hc60f1c62, 32'h00000000} /* (24, 3, 1) {real, imag} */,
  {32'hc60a2230, 32'h00000000} /* (24, 3, 0) {real, imag} */,
  {32'hc60f56c5, 32'h00000000} /* (24, 2, 31) {real, imag} */,
  {32'hc62404c4, 32'h00000000} /* (24, 2, 30) {real, imag} */,
  {32'hc6252ed8, 32'h00000000} /* (24, 2, 29) {real, imag} */,
  {32'hc62b3f52, 32'h00000000} /* (24, 2, 28) {real, imag} */,
  {32'hc6372dc0, 32'h00000000} /* (24, 2, 27) {real, imag} */,
  {32'hc62abe92, 32'h00000000} /* (24, 2, 26) {real, imag} */,
  {32'hc620244a, 32'h00000000} /* (24, 2, 25) {real, imag} */,
  {32'hc6131c79, 32'h00000000} /* (24, 2, 24) {real, imag} */,
  {32'hc603abc4, 32'h00000000} /* (24, 2, 23) {real, imag} */,
  {32'hc5ecc50c, 32'h00000000} /* (24, 2, 22) {real, imag} */,
  {32'hc5de25a1, 32'h00000000} /* (24, 2, 21) {real, imag} */,
  {32'hc5ba07e6, 32'h00000000} /* (24, 2, 20) {real, imag} */,
  {32'hc5b69eb7, 32'h00000000} /* (24, 2, 19) {real, imag} */,
  {32'hc583e6cc, 32'h00000000} /* (24, 2, 18) {real, imag} */,
  {32'hc51a420a, 32'h00000000} /* (24, 2, 17) {real, imag} */,
  {32'hc3b8c8d0, 32'h00000000} /* (24, 2, 16) {real, imag} */,
  {32'h450d1c6f, 32'h00000000} /* (24, 2, 15) {real, imag} */,
  {32'h45551fa1, 32'h00000000} /* (24, 2, 14) {real, imag} */,
  {32'h45a25fa7, 32'h00000000} /* (24, 2, 13) {real, imag} */,
  {32'h45c493b8, 32'h00000000} /* (24, 2, 12) {real, imag} */,
  {32'h459183f0, 32'h00000000} /* (24, 2, 11) {real, imag} */,
  {32'h45986d9c, 32'h00000000} /* (24, 2, 10) {real, imag} */,
  {32'h456efe4e, 32'h00000000} /* (24, 2, 9) {real, imag} */,
  {32'h4513e46c, 32'h00000000} /* (24, 2, 8) {real, imag} */,
  {32'h44b44492, 32'h00000000} /* (24, 2, 7) {real, imag} */,
  {32'hc3a6e7b8, 32'h00000000} /* (24, 2, 6) {real, imag} */,
  {32'hc52762c6, 32'h00000000} /* (24, 2, 5) {real, imag} */,
  {32'hc5bdd042, 32'h00000000} /* (24, 2, 4) {real, imag} */,
  {32'hc5e797d1, 32'h00000000} /* (24, 2, 3) {real, imag} */,
  {32'hc600c87c, 32'h00000000} /* (24, 2, 2) {real, imag} */,
  {32'hc6078bac, 32'h00000000} /* (24, 2, 1) {real, imag} */,
  {32'hc607b5cc, 32'h00000000} /* (24, 2, 0) {real, imag} */,
  {32'hc60cc893, 32'h00000000} /* (24, 1, 31) {real, imag} */,
  {32'hc616ee0f, 32'h00000000} /* (24, 1, 30) {real, imag} */,
  {32'hc62a4f8a, 32'h00000000} /* (24, 1, 29) {real, imag} */,
  {32'hc62e8b20, 32'h00000000} /* (24, 1, 28) {real, imag} */,
  {32'hc637d9ee, 32'h00000000} /* (24, 1, 27) {real, imag} */,
  {32'hc62efb52, 32'h00000000} /* (24, 1, 26) {real, imag} */,
  {32'hc61dd0d2, 32'h00000000} /* (24, 1, 25) {real, imag} */,
  {32'hc60bdfe7, 32'h00000000} /* (24, 1, 24) {real, imag} */,
  {32'hc602b165, 32'h00000000} /* (24, 1, 23) {real, imag} */,
  {32'hc5e4316e, 32'h00000000} /* (24, 1, 22) {real, imag} */,
  {32'hc5d481a2, 32'h00000000} /* (24, 1, 21) {real, imag} */,
  {32'hc592781a, 32'h00000000} /* (24, 1, 20) {real, imag} */,
  {32'hc59ce2da, 32'h00000000} /* (24, 1, 19) {real, imag} */,
  {32'hc55f330c, 32'h00000000} /* (24, 1, 18) {real, imag} */,
  {32'hc4f016a8, 32'h00000000} /* (24, 1, 17) {real, imag} */,
  {32'h43e32048, 32'h00000000} /* (24, 1, 16) {real, imag} */,
  {32'h452d72af, 32'h00000000} /* (24, 1, 15) {real, imag} */,
  {32'h456fdb3b, 32'h00000000} /* (24, 1, 14) {real, imag} */,
  {32'h458d8c65, 32'h00000000} /* (24, 1, 13) {real, imag} */,
  {32'h4589454a, 32'h00000000} /* (24, 1, 12) {real, imag} */,
  {32'h45a84847, 32'h00000000} /* (24, 1, 11) {real, imag} */,
  {32'h456d4190, 32'h00000000} /* (24, 1, 10) {real, imag} */,
  {32'h4541071e, 32'h00000000} /* (24, 1, 9) {real, imag} */,
  {32'h44ead25a, 32'h00000000} /* (24, 1, 8) {real, imag} */,
  {32'h445af224, 32'h00000000} /* (24, 1, 7) {real, imag} */,
  {32'hc4a64638, 32'h00000000} /* (24, 1, 6) {real, imag} */,
  {32'hc57d9f93, 32'h00000000} /* (24, 1, 5) {real, imag} */,
  {32'hc5b7e9b6, 32'h00000000} /* (24, 1, 4) {real, imag} */,
  {32'hc5ecc174, 32'h00000000} /* (24, 1, 3) {real, imag} */,
  {32'hc602c4ab, 32'h00000000} /* (24, 1, 2) {real, imag} */,
  {32'hc6076c56, 32'h00000000} /* (24, 1, 1) {real, imag} */,
  {32'hc605f446, 32'h00000000} /* (24, 1, 0) {real, imag} */,
  {32'hc60ead88, 32'h00000000} /* (24, 0, 31) {real, imag} */,
  {32'hc61bd420, 32'h00000000} /* (24, 0, 30) {real, imag} */,
  {32'hc6298a96, 32'h00000000} /* (24, 0, 29) {real, imag} */,
  {32'hc62ba2da, 32'h00000000} /* (24, 0, 28) {real, imag} */,
  {32'hc62d15bb, 32'h00000000} /* (24, 0, 27) {real, imag} */,
  {32'hc62a4784, 32'h00000000} /* (24, 0, 26) {real, imag} */,
  {32'hc613d64e, 32'h00000000} /* (24, 0, 25) {real, imag} */,
  {32'hc6030012, 32'h00000000} /* (24, 0, 24) {real, imag} */,
  {32'hc5f38444, 32'h00000000} /* (24, 0, 23) {real, imag} */,
  {32'hc5c64d57, 32'h00000000} /* (24, 0, 22) {real, imag} */,
  {32'hc597d426, 32'h00000000} /* (24, 0, 21) {real, imag} */,
  {32'hc55da7d7, 32'h00000000} /* (24, 0, 20) {real, imag} */,
  {32'hc538abb1, 32'h00000000} /* (24, 0, 19) {real, imag} */,
  {32'hc485712e, 32'h00000000} /* (24, 0, 18) {real, imag} */,
  {32'h4286a940, 32'h00000000} /* (24, 0, 17) {real, imag} */,
  {32'h448ace7c, 32'h00000000} /* (24, 0, 16) {real, imag} */,
  {32'h451f785d, 32'h00000000} /* (24, 0, 15) {real, imag} */,
  {32'h4577f1fd, 32'h00000000} /* (24, 0, 14) {real, imag} */,
  {32'h45674dd8, 32'h00000000} /* (24, 0, 13) {real, imag} */,
  {32'h456305bd, 32'h00000000} /* (24, 0, 12) {real, imag} */,
  {32'h4548930b, 32'h00000000} /* (24, 0, 11) {real, imag} */,
  {32'h4504b678, 32'h00000000} /* (24, 0, 10) {real, imag} */,
  {32'h44898754, 32'h00000000} /* (24, 0, 9) {real, imag} */,
  {32'h445a1b98, 32'h00000000} /* (24, 0, 8) {real, imag} */,
  {32'hc48164e2, 32'h00000000} /* (24, 0, 7) {real, imag} */,
  {32'hc52981b2, 32'h00000000} /* (24, 0, 6) {real, imag} */,
  {32'hc58c334e, 32'h00000000} /* (24, 0, 5) {real, imag} */,
  {32'hc5c1ed34, 32'h00000000} /* (24, 0, 4) {real, imag} */,
  {32'hc5e22f1a, 32'h00000000} /* (24, 0, 3) {real, imag} */,
  {32'hc5fcf610, 32'h00000000} /* (24, 0, 2) {real, imag} */,
  {32'hc6033b94, 32'h00000000} /* (24, 0, 1) {real, imag} */,
  {32'hc60a65bc, 32'h00000000} /* (24, 0, 0) {real, imag} */,
  {32'hc62f4df8, 32'h00000000} /* (23, 31, 31) {real, imag} */,
  {32'hc63f57ad, 32'h00000000} /* (23, 31, 30) {real, imag} */,
  {32'hc63f450f, 32'h00000000} /* (23, 31, 29) {real, imag} */,
  {32'hc641a0fa, 32'h00000000} /* (23, 31, 28) {real, imag} */,
  {32'hc63b29aa, 32'h00000000} /* (23, 31, 27) {real, imag} */,
  {32'hc6475268, 32'h00000000} /* (23, 31, 26) {real, imag} */,
  {32'hc6370d49, 32'h00000000} /* (23, 31, 25) {real, imag} */,
  {32'hc62114c5, 32'h00000000} /* (23, 31, 24) {real, imag} */,
  {32'hc60d4464, 32'h00000000} /* (23, 31, 23) {real, imag} */,
  {32'hc600c474, 32'h00000000} /* (23, 31, 22) {real, imag} */,
  {32'hc5a2998a, 32'h00000000} /* (23, 31, 21) {real, imag} */,
  {32'hc4ef7802, 32'h00000000} /* (23, 31, 20) {real, imag} */,
  {32'hc495f8d2, 32'h00000000} /* (23, 31, 19) {real, imag} */,
  {32'h44246518, 32'h00000000} /* (23, 31, 18) {real, imag} */,
  {32'h4520a6c7, 32'h00000000} /* (23, 31, 17) {real, imag} */,
  {32'h4551059e, 32'h00000000} /* (23, 31, 16) {real, imag} */,
  {32'h458ee07a, 32'h00000000} /* (23, 31, 15) {real, imag} */,
  {32'h459e9cd6, 32'h00000000} /* (23, 31, 14) {real, imag} */,
  {32'h45a2a232, 32'h00000000} /* (23, 31, 13) {real, imag} */,
  {32'h458dfb08, 32'h00000000} /* (23, 31, 12) {real, imag} */,
  {32'h454f4d0a, 32'h00000000} /* (23, 31, 11) {real, imag} */,
  {32'h448b7664, 32'h00000000} /* (23, 31, 10) {real, imag} */,
  {32'hc43b7010, 32'h00000000} /* (23, 31, 9) {real, imag} */,
  {32'hc5297e59, 32'h00000000} /* (23, 31, 8) {real, imag} */,
  {32'hc544f4f4, 32'h00000000} /* (23, 31, 7) {real, imag} */,
  {32'hc5a089c0, 32'h00000000} /* (23, 31, 6) {real, imag} */,
  {32'hc5d19d1a, 32'h00000000} /* (23, 31, 5) {real, imag} */,
  {32'hc5f51bf4, 32'h00000000} /* (23, 31, 4) {real, imag} */,
  {32'hc60a8503, 32'h00000000} /* (23, 31, 3) {real, imag} */,
  {32'hc61313c4, 32'h00000000} /* (23, 31, 2) {real, imag} */,
  {32'hc61f28b8, 32'h00000000} /* (23, 31, 1) {real, imag} */,
  {32'hc625b1b0, 32'h00000000} /* (23, 31, 0) {real, imag} */,
  {32'hc62eb338, 32'h00000000} /* (23, 30, 31) {real, imag} */,
  {32'hc6438f85, 32'h00000000} /* (23, 30, 30) {real, imag} */,
  {32'hc64beef1, 32'h00000000} /* (23, 30, 29) {real, imag} */,
  {32'hc642989a, 32'h00000000} /* (23, 30, 28) {real, imag} */,
  {32'hc649673d, 32'h00000000} /* (23, 30, 27) {real, imag} */,
  {32'hc6444b26, 32'h00000000} /* (23, 30, 26) {real, imag} */,
  {32'hc636f3c6, 32'h00000000} /* (23, 30, 25) {real, imag} */,
  {32'hc63a6bba, 32'h00000000} /* (23, 30, 24) {real, imag} */,
  {32'hc619e326, 32'h00000000} /* (23, 30, 23) {real, imag} */,
  {32'hc5edf9e8, 32'h00000000} /* (23, 30, 22) {real, imag} */,
  {32'hc5a56a99, 32'h00000000} /* (23, 30, 21) {real, imag} */,
  {32'hc44be704, 32'h00000000} /* (23, 30, 20) {real, imag} */,
  {32'h43cf7470, 32'h00000000} /* (23, 30, 19) {real, imag} */,
  {32'h4526c9d8, 32'h00000000} /* (23, 30, 18) {real, imag} */,
  {32'h45764bce, 32'h00000000} /* (23, 30, 17) {real, imag} */,
  {32'h45b224f1, 32'h00000000} /* (23, 30, 16) {real, imag} */,
  {32'h45a40378, 32'h00000000} /* (23, 30, 15) {real, imag} */,
  {32'h45acc932, 32'h00000000} /* (23, 30, 14) {real, imag} */,
  {32'h45a21d4e, 32'h00000000} /* (23, 30, 13) {real, imag} */,
  {32'h45980b10, 32'h00000000} /* (23, 30, 12) {real, imag} */,
  {32'h4587c006, 32'h00000000} /* (23, 30, 11) {real, imag} */,
  {32'h4339f480, 32'h00000000} /* (23, 30, 10) {real, imag} */,
  {32'hc53ca800, 32'h00000000} /* (23, 30, 9) {real, imag} */,
  {32'hc58a1297, 32'h00000000} /* (23, 30, 8) {real, imag} */,
  {32'hc58fa339, 32'h00000000} /* (23, 30, 7) {real, imag} */,
  {32'hc5cca258, 32'h00000000} /* (23, 30, 6) {real, imag} */,
  {32'hc5f20cb7, 32'h00000000} /* (23, 30, 5) {real, imag} */,
  {32'hc60c9cdb, 32'h00000000} /* (23, 30, 4) {real, imag} */,
  {32'hc61fee90, 32'h00000000} /* (23, 30, 3) {real, imag} */,
  {32'hc61cf47a, 32'h00000000} /* (23, 30, 2) {real, imag} */,
  {32'hc6238228, 32'h00000000} /* (23, 30, 1) {real, imag} */,
  {32'hc62c65e4, 32'h00000000} /* (23, 30, 0) {real, imag} */,
  {32'hc635bc99, 32'h00000000} /* (23, 29, 31) {real, imag} */,
  {32'hc6438b04, 32'h00000000} /* (23, 29, 30) {real, imag} */,
  {32'hc6413562, 32'h00000000} /* (23, 29, 29) {real, imag} */,
  {32'hc64b0189, 32'h00000000} /* (23, 29, 28) {real, imag} */,
  {32'hc64829f7, 32'h00000000} /* (23, 29, 27) {real, imag} */,
  {32'hc6439232, 32'h00000000} /* (23, 29, 26) {real, imag} */,
  {32'hc64ba89c, 32'h00000000} /* (23, 29, 25) {real, imag} */,
  {32'hc632b7a8, 32'h00000000} /* (23, 29, 24) {real, imag} */,
  {32'hc616d9fa, 32'h00000000} /* (23, 29, 23) {real, imag} */,
  {32'hc5daa576, 32'h00000000} /* (23, 29, 22) {real, imag} */,
  {32'hc594379a, 32'h00000000} /* (23, 29, 21) {real, imag} */,
  {32'hc4ae34d6, 32'h00000000} /* (23, 29, 20) {real, imag} */,
  {32'h45039576, 32'h00000000} /* (23, 29, 19) {real, imag} */,
  {32'h4589bb8c, 32'h00000000} /* (23, 29, 18) {real, imag} */,
  {32'h45b1f987, 32'h00000000} /* (23, 29, 17) {real, imag} */,
  {32'h45bc8669, 32'h00000000} /* (23, 29, 16) {real, imag} */,
  {32'h45c06b46, 32'h00000000} /* (23, 29, 15) {real, imag} */,
  {32'h45b33773, 32'h00000000} /* (23, 29, 14) {real, imag} */,
  {32'h45a3b244, 32'h00000000} /* (23, 29, 13) {real, imag} */,
  {32'h458e61a6, 32'h00000000} /* (23, 29, 12) {real, imag} */,
  {32'h452dee3c, 32'h00000000} /* (23, 29, 11) {real, imag} */,
  {32'h4382ef80, 32'h00000000} /* (23, 29, 10) {real, imag} */,
  {32'hc5578bbe, 32'h00000000} /* (23, 29, 9) {real, imag} */,
  {32'hc5ada110, 32'h00000000} /* (23, 29, 8) {real, imag} */,
  {32'hc5dbb900, 32'h00000000} /* (23, 29, 7) {real, imag} */,
  {32'hc5eb58f0, 32'h00000000} /* (23, 29, 6) {real, imag} */,
  {32'hc605be6d, 32'h00000000} /* (23, 29, 5) {real, imag} */,
  {32'hc6126fbf, 32'h00000000} /* (23, 29, 4) {real, imag} */,
  {32'hc6160e22, 32'h00000000} /* (23, 29, 3) {real, imag} */,
  {32'hc62e644e, 32'h00000000} /* (23, 29, 2) {real, imag} */,
  {32'hc635e800, 32'h00000000} /* (23, 29, 1) {real, imag} */,
  {32'hc62f8a98, 32'h00000000} /* (23, 29, 0) {real, imag} */,
  {32'hc646658f, 32'h00000000} /* (23, 28, 31) {real, imag} */,
  {32'hc64327d7, 32'h00000000} /* (23, 28, 30) {real, imag} */,
  {32'hc644fc97, 32'h00000000} /* (23, 28, 29) {real, imag} */,
  {32'hc64333ae, 32'h00000000} /* (23, 28, 28) {real, imag} */,
  {32'hc644e848, 32'h00000000} /* (23, 28, 27) {real, imag} */,
  {32'hc63cc126, 32'h00000000} /* (23, 28, 26) {real, imag} */,
  {32'hc64582ca, 32'h00000000} /* (23, 28, 25) {real, imag} */,
  {32'hc62f72c3, 32'h00000000} /* (23, 28, 24) {real, imag} */,
  {32'hc60c9146, 32'h00000000} /* (23, 28, 23) {real, imag} */,
  {32'hc5d7dff5, 32'h00000000} /* (23, 28, 22) {real, imag} */,
  {32'hc581e6b4, 32'h00000000} /* (23, 28, 21) {real, imag} */,
  {32'hc307a340, 32'h00000000} /* (23, 28, 20) {real, imag} */,
  {32'h4533ca02, 32'h00000000} /* (23, 28, 19) {real, imag} */,
  {32'h458fc0e5, 32'h00000000} /* (23, 28, 18) {real, imag} */,
  {32'h45b9e23b, 32'h00000000} /* (23, 28, 17) {real, imag} */,
  {32'h45d9fec9, 32'h00000000} /* (23, 28, 16) {real, imag} */,
  {32'h45e878e2, 32'h00000000} /* (23, 28, 15) {real, imag} */,
  {32'h45d3b7b2, 32'h00000000} /* (23, 28, 14) {real, imag} */,
  {32'h45a7bac2, 32'h00000000} /* (23, 28, 13) {real, imag} */,
  {32'h45912ffd, 32'h00000000} /* (23, 28, 12) {real, imag} */,
  {32'h45117312, 32'h00000000} /* (23, 28, 11) {real, imag} */,
  {32'hc4764928, 32'h00000000} /* (23, 28, 10) {real, imag} */,
  {32'hc56f38f8, 32'h00000000} /* (23, 28, 9) {real, imag} */,
  {32'hc5e055ca, 32'h00000000} /* (23, 28, 8) {real, imag} */,
  {32'hc5fc0a28, 32'h00000000} /* (23, 28, 7) {real, imag} */,
  {32'hc608cebe, 32'h00000000} /* (23, 28, 6) {real, imag} */,
  {32'hc612c14a, 32'h00000000} /* (23, 28, 5) {real, imag} */,
  {32'hc61ae968, 32'h00000000} /* (23, 28, 4) {real, imag} */,
  {32'hc62faf6e, 32'h00000000} /* (23, 28, 3) {real, imag} */,
  {32'hc63c65a8, 32'h00000000} /* (23, 28, 2) {real, imag} */,
  {32'hc6361d1a, 32'h00000000} /* (23, 28, 1) {real, imag} */,
  {32'hc629eccc, 32'h00000000} /* (23, 28, 0) {real, imag} */,
  {32'hc62d0a20, 32'h00000000} /* (23, 27, 31) {real, imag} */,
  {32'hc64acf81, 32'h00000000} /* (23, 27, 30) {real, imag} */,
  {32'hc6415a1e, 32'h00000000} /* (23, 27, 29) {real, imag} */,
  {32'hc6448f4c, 32'h00000000} /* (23, 27, 28) {real, imag} */,
  {32'hc6541ab0, 32'h00000000} /* (23, 27, 27) {real, imag} */,
  {32'hc644f7ea, 32'h00000000} /* (23, 27, 26) {real, imag} */,
  {32'hc636b244, 32'h00000000} /* (23, 27, 25) {real, imag} */,
  {32'hc624a11c, 32'h00000000} /* (23, 27, 24) {real, imag} */,
  {32'hc603dad0, 32'h00000000} /* (23, 27, 23) {real, imag} */,
  {32'hc5c3d012, 32'h00000000} /* (23, 27, 22) {real, imag} */,
  {32'hc5636a15, 32'h00000000} /* (23, 27, 21) {real, imag} */,
  {32'hc3ae8580, 32'h00000000} /* (23, 27, 20) {real, imag} */,
  {32'h453a81a6, 32'h00000000} /* (23, 27, 19) {real, imag} */,
  {32'h45abc4d4, 32'h00000000} /* (23, 27, 18) {real, imag} */,
  {32'h45bd08fd, 32'h00000000} /* (23, 27, 17) {real, imag} */,
  {32'h45d5e986, 32'h00000000} /* (23, 27, 16) {real, imag} */,
  {32'h45ca0d19, 32'h00000000} /* (23, 27, 15) {real, imag} */,
  {32'h45c2fdd6, 32'h00000000} /* (23, 27, 14) {real, imag} */,
  {32'h45b78675, 32'h00000000} /* (23, 27, 13) {real, imag} */,
  {32'h457f2fc6, 32'h00000000} /* (23, 27, 12) {real, imag} */,
  {32'h45126fe8, 32'h00000000} /* (23, 27, 11) {real, imag} */,
  {32'hc4e3c43c, 32'h00000000} /* (23, 27, 10) {real, imag} */,
  {32'hc59f097f, 32'h00000000} /* (23, 27, 9) {real, imag} */,
  {32'hc5c92183, 32'h00000000} /* (23, 27, 8) {real, imag} */,
  {32'hc5fe9089, 32'h00000000} /* (23, 27, 7) {real, imag} */,
  {32'hc60d2f3f, 32'h00000000} /* (23, 27, 6) {real, imag} */,
  {32'hc61f2e9a, 32'h00000000} /* (23, 27, 5) {real, imag} */,
  {32'hc62aa51d, 32'h00000000} /* (23, 27, 4) {real, imag} */,
  {32'hc6420d96, 32'h00000000} /* (23, 27, 3) {real, imag} */,
  {32'hc63b73c6, 32'h00000000} /* (23, 27, 2) {real, imag} */,
  {32'hc623fb60, 32'h00000000} /* (23, 27, 1) {real, imag} */,
  {32'hc62b81f5, 32'h00000000} /* (23, 27, 0) {real, imag} */,
  {32'hc6280964, 32'h00000000} /* (23, 26, 31) {real, imag} */,
  {32'hc630fb8a, 32'h00000000} /* (23, 26, 30) {real, imag} */,
  {32'hc63cd6c0, 32'h00000000} /* (23, 26, 29) {real, imag} */,
  {32'hc644714f, 32'h00000000} /* (23, 26, 28) {real, imag} */,
  {32'hc6498613, 32'h00000000} /* (23, 26, 27) {real, imag} */,
  {32'hc64f1f8c, 32'h00000000} /* (23, 26, 26) {real, imag} */,
  {32'hc62f4a71, 32'h00000000} /* (23, 26, 25) {real, imag} */,
  {32'hc6195580, 32'h00000000} /* (23, 26, 24) {real, imag} */,
  {32'hc60b0f3c, 32'h00000000} /* (23, 26, 23) {real, imag} */,
  {32'hc5cbb816, 32'h00000000} /* (23, 26, 22) {real, imag} */,
  {32'hc51f460d, 32'h00000000} /* (23, 26, 21) {real, imag} */,
  {32'h431e6540, 32'h00000000} /* (23, 26, 20) {real, imag} */,
  {32'h4540696a, 32'h00000000} /* (23, 26, 19) {real, imag} */,
  {32'h45ab5642, 32'h00000000} /* (23, 26, 18) {real, imag} */,
  {32'h45cd439e, 32'h00000000} /* (23, 26, 17) {real, imag} */,
  {32'h45b5893a, 32'h00000000} /* (23, 26, 16) {real, imag} */,
  {32'h45d8ca0f, 32'h00000000} /* (23, 26, 15) {real, imag} */,
  {32'h45c08ab0, 32'h00000000} /* (23, 26, 14) {real, imag} */,
  {32'h45982f81, 32'h00000000} /* (23, 26, 13) {real, imag} */,
  {32'h455c3428, 32'h00000000} /* (23, 26, 12) {real, imag} */,
  {32'h44ab4608, 32'h00000000} /* (23, 26, 11) {real, imag} */,
  {32'hc4f3d5fc, 32'h00000000} /* (23, 26, 10) {real, imag} */,
  {32'hc5991c2a, 32'h00000000} /* (23, 26, 9) {real, imag} */,
  {32'hc5caaccf, 32'h00000000} /* (23, 26, 8) {real, imag} */,
  {32'hc5fcc9b8, 32'h00000000} /* (23, 26, 7) {real, imag} */,
  {32'hc6098b35, 32'h00000000} /* (23, 26, 6) {real, imag} */,
  {32'hc60d5ee2, 32'h00000000} /* (23, 26, 5) {real, imag} */,
  {32'hc62326a4, 32'h00000000} /* (23, 26, 4) {real, imag} */,
  {32'hc62615d6, 32'h00000000} /* (23, 26, 3) {real, imag} */,
  {32'hc62daa03, 32'h00000000} /* (23, 26, 2) {real, imag} */,
  {32'hc6268de9, 32'h00000000} /* (23, 26, 1) {real, imag} */,
  {32'hc6269469, 32'h00000000} /* (23, 26, 0) {real, imag} */,
  {32'hc62027a5, 32'h00000000} /* (23, 25, 31) {real, imag} */,
  {32'hc6348414, 32'h00000000} /* (23, 25, 30) {real, imag} */,
  {32'hc6309f6f, 32'h00000000} /* (23, 25, 29) {real, imag} */,
  {32'hc62fd1f7, 32'h00000000} /* (23, 25, 28) {real, imag} */,
  {32'hc62b7f7e, 32'h00000000} /* (23, 25, 27) {real, imag} */,
  {32'hc6292aa4, 32'h00000000} /* (23, 25, 26) {real, imag} */,
  {32'hc6283002, 32'h00000000} /* (23, 25, 25) {real, imag} */,
  {32'hc613b23c, 32'h00000000} /* (23, 25, 24) {real, imag} */,
  {32'hc5f833d2, 32'h00000000} /* (23, 25, 23) {real, imag} */,
  {32'hc5ae6915, 32'h00000000} /* (23, 25, 22) {real, imag} */,
  {32'hc53c5723, 32'h00000000} /* (23, 25, 21) {real, imag} */,
  {32'h4481db58, 32'h00000000} /* (23, 25, 20) {real, imag} */,
  {32'h4564b82e, 32'h00000000} /* (23, 25, 19) {real, imag} */,
  {32'h45a15d48, 32'h00000000} /* (23, 25, 18) {real, imag} */,
  {32'h45bc53c2, 32'h00000000} /* (23, 25, 17) {real, imag} */,
  {32'h45cc386e, 32'h00000000} /* (23, 25, 16) {real, imag} */,
  {32'h45d067ea, 32'h00000000} /* (23, 25, 15) {real, imag} */,
  {32'h45d11708, 32'h00000000} /* (23, 25, 14) {real, imag} */,
  {32'h45b7dffe, 32'h00000000} /* (23, 25, 13) {real, imag} */,
  {32'h45593bf5, 32'h00000000} /* (23, 25, 12) {real, imag} */,
  {32'h446d0f78, 32'h00000000} /* (23, 25, 11) {real, imag} */,
  {32'hc563b887, 32'h00000000} /* (23, 25, 10) {real, imag} */,
  {32'hc5a6925d, 32'h00000000} /* (23, 25, 9) {real, imag} */,
  {32'hc5c2530c, 32'h00000000} /* (23, 25, 8) {real, imag} */,
  {32'hc5f06db6, 32'h00000000} /* (23, 25, 7) {real, imag} */,
  {32'hc6089fa4, 32'h00000000} /* (23, 25, 6) {real, imag} */,
  {32'hc60afb27, 32'h00000000} /* (23, 25, 5) {real, imag} */,
  {32'hc61b7517, 32'h00000000} /* (23, 25, 4) {real, imag} */,
  {32'hc6250d04, 32'h00000000} /* (23, 25, 3) {real, imag} */,
  {32'hc6289f80, 32'h00000000} /* (23, 25, 2) {real, imag} */,
  {32'hc614a6e5, 32'h00000000} /* (23, 25, 1) {real, imag} */,
  {32'hc60bc807, 32'h00000000} /* (23, 25, 0) {real, imag} */,
  {32'hc607fd28, 32'h00000000} /* (23, 24, 31) {real, imag} */,
  {32'hc6136039, 32'h00000000} /* (23, 24, 30) {real, imag} */,
  {32'hc61b64c2, 32'h00000000} /* (23, 24, 29) {real, imag} */,
  {32'hc61ead9e, 32'h00000000} /* (23, 24, 28) {real, imag} */,
  {32'hc6247dc2, 32'h00000000} /* (23, 24, 27) {real, imag} */,
  {32'hc609be02, 32'h00000000} /* (23, 24, 26) {real, imag} */,
  {32'hc6040400, 32'h00000000} /* (23, 24, 25) {real, imag} */,
  {32'hc5ec5bb7, 32'h00000000} /* (23, 24, 24) {real, imag} */,
  {32'hc5d65da7, 32'h00000000} /* (23, 24, 23) {real, imag} */,
  {32'hc5af2756, 32'h00000000} /* (23, 24, 22) {real, imag} */,
  {32'hc520c8d7, 32'h00000000} /* (23, 24, 21) {real, imag} */,
  {32'h44388a9c, 32'h00000000} /* (23, 24, 20) {real, imag} */,
  {32'h45343103, 32'h00000000} /* (23, 24, 19) {real, imag} */,
  {32'h45988bc9, 32'h00000000} /* (23, 24, 18) {real, imag} */,
  {32'h45c987a9, 32'h00000000} /* (23, 24, 17) {real, imag} */,
  {32'h45d22dd6, 32'h00000000} /* (23, 24, 16) {real, imag} */,
  {32'h45b8e6e8, 32'h00000000} /* (23, 24, 15) {real, imag} */,
  {32'h45dfb092, 32'h00000000} /* (23, 24, 14) {real, imag} */,
  {32'h45992d2d, 32'h00000000} /* (23, 24, 13) {real, imag} */,
  {32'h4546aaaf, 32'h00000000} /* (23, 24, 12) {real, imag} */,
  {32'h43d48800, 32'h00000000} /* (23, 24, 11) {real, imag} */,
  {32'hc5127a16, 32'h00000000} /* (23, 24, 10) {real, imag} */,
  {32'hc595c60b, 32'h00000000} /* (23, 24, 9) {real, imag} */,
  {32'hc5c7b36f, 32'h00000000} /* (23, 24, 8) {real, imag} */,
  {32'hc5fbce65, 32'h00000000} /* (23, 24, 7) {real, imag} */,
  {32'hc5fb9662, 32'h00000000} /* (23, 24, 6) {real, imag} */,
  {32'hc6016579, 32'h00000000} /* (23, 24, 5) {real, imag} */,
  {32'hc603a2fe, 32'h00000000} /* (23, 24, 4) {real, imag} */,
  {32'hc616e6c9, 32'h00000000} /* (23, 24, 3) {real, imag} */,
  {32'hc614253a, 32'h00000000} /* (23, 24, 2) {real, imag} */,
  {32'hc60764b2, 32'h00000000} /* (23, 24, 1) {real, imag} */,
  {32'hc5fea286, 32'h00000000} /* (23, 24, 0) {real, imag} */,
  {32'hc5ed109c, 32'h00000000} /* (23, 23, 31) {real, imag} */,
  {32'hc5f29265, 32'h00000000} /* (23, 23, 30) {real, imag} */,
  {32'hc5ec064f, 32'h00000000} /* (23, 23, 29) {real, imag} */,
  {32'hc60695bc, 32'h00000000} /* (23, 23, 28) {real, imag} */,
  {32'hc603cb04, 32'h00000000} /* (23, 23, 27) {real, imag} */,
  {32'hc5e77276, 32'h00000000} /* (23, 23, 26) {real, imag} */,
  {32'hc5ea0742, 32'h00000000} /* (23, 23, 25) {real, imag} */,
  {32'hc5c31d85, 32'h00000000} /* (23, 23, 24) {real, imag} */,
  {32'hc5b93d0c, 32'h00000000} /* (23, 23, 23) {real, imag} */,
  {32'hc5843fad, 32'h00000000} /* (23, 23, 22) {real, imag} */,
  {32'hc4fef49c, 32'h00000000} /* (23, 23, 21) {real, imag} */,
  {32'h4468f4a8, 32'h00000000} /* (23, 23, 20) {real, imag} */,
  {32'h45536c7e, 32'h00000000} /* (23, 23, 19) {real, imag} */,
  {32'h458d7a7e, 32'h00000000} /* (23, 23, 18) {real, imag} */,
  {32'h45c4aa00, 32'h00000000} /* (23, 23, 17) {real, imag} */,
  {32'h45a6b1a4, 32'h00000000} /* (23, 23, 16) {real, imag} */,
  {32'h45af05d0, 32'h00000000} /* (23, 23, 15) {real, imag} */,
  {32'h45b5c01d, 32'h00000000} /* (23, 23, 14) {real, imag} */,
  {32'h457e5036, 32'h00000000} /* (23, 23, 13) {real, imag} */,
  {32'h4546ef04, 32'h00000000} /* (23, 23, 12) {real, imag} */,
  {32'h44409018, 32'h00000000} /* (23, 23, 11) {real, imag} */,
  {32'hc4f605f8, 32'h00000000} /* (23, 23, 10) {real, imag} */,
  {32'hc5577cc7, 32'h00000000} /* (23, 23, 9) {real, imag} */,
  {32'hc5a9b2ab, 32'h00000000} /* (23, 23, 8) {real, imag} */,
  {32'hc5ceaba0, 32'h00000000} /* (23, 23, 7) {real, imag} */,
  {32'hc5d0f5b5, 32'h00000000} /* (23, 23, 6) {real, imag} */,
  {32'hc5d6f85b, 32'h00000000} /* (23, 23, 5) {real, imag} */,
  {32'hc5f20645, 32'h00000000} /* (23, 23, 4) {real, imag} */,
  {32'hc5e5dd43, 32'h00000000} /* (23, 23, 3) {real, imag} */,
  {32'hc5d3e0d8, 32'h00000000} /* (23, 23, 2) {real, imag} */,
  {32'hc5d3aa94, 32'h00000000} /* (23, 23, 1) {real, imag} */,
  {32'hc5e618c4, 32'h00000000} /* (23, 23, 0) {real, imag} */,
  {32'hc59dc893, 32'h00000000} /* (23, 22, 31) {real, imag} */,
  {32'hc5a3a078, 32'h00000000} /* (23, 22, 30) {real, imag} */,
  {32'hc5afa9d4, 32'h00000000} /* (23, 22, 29) {real, imag} */,
  {32'hc5ac00b5, 32'h00000000} /* (23, 22, 28) {real, imag} */,
  {32'hc59b42a5, 32'h00000000} /* (23, 22, 27) {real, imag} */,
  {32'hc5990a47, 32'h00000000} /* (23, 22, 26) {real, imag} */,
  {32'hc590d7bc, 32'h00000000} /* (23, 22, 25) {real, imag} */,
  {32'hc590fdd3, 32'h00000000} /* (23, 22, 24) {real, imag} */,
  {32'hc571a3aa, 32'h00000000} /* (23, 22, 23) {real, imag} */,
  {32'hc54eb7df, 32'h00000000} /* (23, 22, 22) {real, imag} */,
  {32'hc4bdf069, 32'h00000000} /* (23, 22, 21) {real, imag} */,
  {32'h4496b01a, 32'h00000000} /* (23, 22, 20) {real, imag} */,
  {32'h454d1a39, 32'h00000000} /* (23, 22, 19) {real, imag} */,
  {32'h4579c06c, 32'h00000000} /* (23, 22, 18) {real, imag} */,
  {32'h45567e94, 32'h00000000} /* (23, 22, 17) {real, imag} */,
  {32'h458c044c, 32'h00000000} /* (23, 22, 16) {real, imag} */,
  {32'h456854fa, 32'h00000000} /* (23, 22, 15) {real, imag} */,
  {32'h455e29d1, 32'h00000000} /* (23, 22, 14) {real, imag} */,
  {32'h45484ac9, 32'h00000000} /* (23, 22, 13) {real, imag} */,
  {32'h4520df5c, 32'h00000000} /* (23, 22, 12) {real, imag} */,
  {32'h447b8ce8, 32'h00000000} /* (23, 22, 11) {real, imag} */,
  {32'hc49ddc93, 32'h00000000} /* (23, 22, 10) {real, imag} */,
  {32'hc532c664, 32'h00000000} /* (23, 22, 9) {real, imag} */,
  {32'hc574a0a3, 32'h00000000} /* (23, 22, 8) {real, imag} */,
  {32'hc584ce2d, 32'h00000000} /* (23, 22, 7) {real, imag} */,
  {32'hc58f484e, 32'h00000000} /* (23, 22, 6) {real, imag} */,
  {32'hc5a0ab4f, 32'h00000000} /* (23, 22, 5) {real, imag} */,
  {32'hc5a7ae0c, 32'h00000000} /* (23, 22, 4) {real, imag} */,
  {32'hc5a88c5a, 32'h00000000} /* (23, 22, 3) {real, imag} */,
  {32'hc590a062, 32'h00000000} /* (23, 22, 2) {real, imag} */,
  {32'hc59bccc8, 32'h00000000} /* (23, 22, 1) {real, imag} */,
  {32'hc5a0ed48, 32'h00000000} /* (23, 22, 0) {real, imag} */,
  {32'hc4eabe88, 32'h00000000} /* (23, 21, 31) {real, imag} */,
  {32'hc51d7910, 32'h00000000} /* (23, 21, 30) {real, imag} */,
  {32'hc54a47f7, 32'h00000000} /* (23, 21, 29) {real, imag} */,
  {32'hc548baac, 32'h00000000} /* (23, 21, 28) {real, imag} */,
  {32'hc5021ad5, 32'h00000000} /* (23, 21, 27) {real, imag} */,
  {32'hc4523bc0, 32'h00000000} /* (23, 21, 26) {real, imag} */,
  {32'hc4e1ef36, 32'h00000000} /* (23, 21, 25) {real, imag} */,
  {32'hc4df5cc2, 32'h00000000} /* (23, 21, 24) {real, imag} */,
  {32'hc46c9195, 32'h00000000} /* (23, 21, 23) {real, imag} */,
  {32'hc4f31a9e, 32'h00000000} /* (23, 21, 22) {real, imag} */,
  {32'hc4af0e90, 32'h00000000} /* (23, 21, 21) {real, imag} */,
  {32'hc38ba23c, 32'h00000000} /* (23, 21, 20) {real, imag} */,
  {32'h43af8008, 32'h00000000} /* (23, 21, 19) {real, imag} */,
  {32'h4508b504, 32'h00000000} /* (23, 21, 18) {real, imag} */,
  {32'h44c8b30d, 32'h00000000} /* (23, 21, 17) {real, imag} */,
  {32'h4487b181, 32'h00000000} /* (23, 21, 16) {real, imag} */,
  {32'h44429a6c, 32'h00000000} /* (23, 21, 15) {real, imag} */,
  {32'h451d0c2e, 32'h00000000} /* (23, 21, 14) {real, imag} */,
  {32'h44d09236, 32'h00000000} /* (23, 21, 13) {real, imag} */,
  {32'h44266244, 32'h00000000} /* (23, 21, 12) {real, imag} */,
  {32'h404b1000, 32'h00000000} /* (23, 21, 11) {real, imag} */,
  {32'hc4836fc1, 32'h00000000} /* (23, 21, 10) {real, imag} */,
  {32'hc4146ae8, 32'h00000000} /* (23, 21, 9) {real, imag} */,
  {32'hc50c9b05, 32'h00000000} /* (23, 21, 8) {real, imag} */,
  {32'hc50f4952, 32'h00000000} /* (23, 21, 7) {real, imag} */,
  {32'hc5114245, 32'h00000000} /* (23, 21, 6) {real, imag} */,
  {32'hc51b7a66, 32'h00000000} /* (23, 21, 5) {real, imag} */,
  {32'hc529659a, 32'h00000000} /* (23, 21, 4) {real, imag} */,
  {32'hc51d4464, 32'h00000000} /* (23, 21, 3) {real, imag} */,
  {32'hc5101400, 32'h00000000} /* (23, 21, 2) {real, imag} */,
  {32'hc5192323, 32'h00000000} /* (23, 21, 1) {real, imag} */,
  {32'hc522c4de, 32'h00000000} /* (23, 21, 0) {real, imag} */,
  {32'h44bbb24c, 32'h00000000} /* (23, 20, 31) {real, imag} */,
  {32'h451e1243, 32'h00000000} /* (23, 20, 30) {real, imag} */,
  {32'h44c04c6e, 32'h00000000} /* (23, 20, 29) {real, imag} */,
  {32'h44af2b3e, 32'h00000000} /* (23, 20, 28) {real, imag} */,
  {32'h44ce46fc, 32'h00000000} /* (23, 20, 27) {real, imag} */,
  {32'h452e05e0, 32'h00000000} /* (23, 20, 26) {real, imag} */,
  {32'h452ae903, 32'h00000000} /* (23, 20, 25) {real, imag} */,
  {32'h450556d1, 32'h00000000} /* (23, 20, 24) {real, imag} */,
  {32'h451239b4, 32'h00000000} /* (23, 20, 23) {real, imag} */,
  {32'h4432f7fa, 32'h00000000} /* (23, 20, 22) {real, imag} */,
  {32'h43a97cfc, 32'h00000000} /* (23, 20, 21) {real, imag} */,
  {32'hc4d7b508, 32'h00000000} /* (23, 20, 20) {real, imag} */,
  {32'hc5349c3c, 32'h00000000} /* (23, 20, 19) {real, imag} */,
  {32'hc4b5b1fe, 32'h00000000} /* (23, 20, 18) {real, imag} */,
  {32'hc52b0538, 32'h00000000} /* (23, 20, 17) {real, imag} */,
  {32'hc54cfcaa, 32'h00000000} /* (23, 20, 16) {real, imag} */,
  {32'hc4a174ba, 32'h00000000} /* (23, 20, 15) {real, imag} */,
  {32'hc40ee918, 32'h00000000} /* (23, 20, 14) {real, imag} */,
  {32'hc482136a, 32'h00000000} /* (23, 20, 13) {real, imag} */,
  {32'hc48aaf12, 32'h00000000} /* (23, 20, 12) {real, imag} */,
  {32'hc490afb8, 32'h00000000} /* (23, 20, 11) {real, imag} */,
  {32'hc169b880, 32'h00000000} /* (23, 20, 10) {real, imag} */,
  {32'h44ab16c2, 32'h00000000} /* (23, 20, 9) {real, imag} */,
  {32'h44b74fde, 32'h00000000} /* (23, 20, 8) {real, imag} */,
  {32'h448b8b39, 32'h00000000} /* (23, 20, 7) {real, imag} */,
  {32'h44d882a5, 32'h00000000} /* (23, 20, 6) {real, imag} */,
  {32'h448bb843, 32'h00000000} /* (23, 20, 5) {real, imag} */,
  {32'h44895f48, 32'h00000000} /* (23, 20, 4) {real, imag} */,
  {32'h44fd5a98, 32'h00000000} /* (23, 20, 3) {real, imag} */,
  {32'h44219be0, 32'h00000000} /* (23, 20, 2) {real, imag} */,
  {32'h44b5e210, 32'h00000000} /* (23, 20, 1) {real, imag} */,
  {32'h4461a4e8, 32'h00000000} /* (23, 20, 0) {real, imag} */,
  {32'h458c891b, 32'h00000000} /* (23, 19, 31) {real, imag} */,
  {32'h459e809f, 32'h00000000} /* (23, 19, 30) {real, imag} */,
  {32'h457658e8, 32'h00000000} /* (23, 19, 29) {real, imag} */,
  {32'h45801eaf, 32'h00000000} /* (23, 19, 28) {real, imag} */,
  {32'h457f4e6d, 32'h00000000} /* (23, 19, 27) {real, imag} */,
  {32'h45706f06, 32'h00000000} /* (23, 19, 26) {real, imag} */,
  {32'h457b9b1f, 32'h00000000} /* (23, 19, 25) {real, imag} */,
  {32'h45710692, 32'h00000000} /* (23, 19, 24) {real, imag} */,
  {32'h4573a3b6, 32'h00000000} /* (23, 19, 23) {real, imag} */,
  {32'h45451813, 32'h00000000} /* (23, 19, 22) {real, imag} */,
  {32'h43efe798, 32'h00000000} /* (23, 19, 21) {real, imag} */,
  {32'hc4b1a045, 32'h00000000} /* (23, 19, 20) {real, imag} */,
  {32'hc5386649, 32'h00000000} /* (23, 19, 19) {real, imag} */,
  {32'hc57655fa, 32'h00000000} /* (23, 19, 18) {real, imag} */,
  {32'hc576e601, 32'h00000000} /* (23, 19, 17) {real, imag} */,
  {32'hc58342cc, 32'h00000000} /* (23, 19, 16) {real, imag} */,
  {32'hc5481f92, 32'h00000000} /* (23, 19, 15) {real, imag} */,
  {32'hc559be92, 32'h00000000} /* (23, 19, 14) {real, imag} */,
  {32'hc5636214, 32'h00000000} /* (23, 19, 13) {real, imag} */,
  {32'hc520ed42, 32'h00000000} /* (23, 19, 12) {real, imag} */,
  {32'hc50b6557, 32'h00000000} /* (23, 19, 11) {real, imag} */,
  {32'hc470c238, 32'h00000000} /* (23, 19, 10) {real, imag} */,
  {32'h44d9412e, 32'h00000000} /* (23, 19, 9) {real, imag} */,
  {32'h4516455e, 32'h00000000} /* (23, 19, 8) {real, imag} */,
  {32'h4550bdde, 32'h00000000} /* (23, 19, 7) {real, imag} */,
  {32'h457904cd, 32'h00000000} /* (23, 19, 6) {real, imag} */,
  {32'h45908ad8, 32'h00000000} /* (23, 19, 5) {real, imag} */,
  {32'h45933416, 32'h00000000} /* (23, 19, 4) {real, imag} */,
  {32'h4560b221, 32'h00000000} /* (23, 19, 3) {real, imag} */,
  {32'h457db7de, 32'h00000000} /* (23, 19, 2) {real, imag} */,
  {32'h458834d0, 32'h00000000} /* (23, 19, 1) {real, imag} */,
  {32'h45693c2a, 32'h00000000} /* (23, 19, 0) {real, imag} */,
  {32'h45a55a88, 32'h00000000} /* (23, 18, 31) {real, imag} */,
  {32'h45cb366a, 32'h00000000} /* (23, 18, 30) {real, imag} */,
  {32'h45d4130b, 32'h00000000} /* (23, 18, 29) {real, imag} */,
  {32'h45ab5816, 32'h00000000} /* (23, 18, 28) {real, imag} */,
  {32'h45aa29c3, 32'h00000000} /* (23, 18, 27) {real, imag} */,
  {32'h45942505, 32'h00000000} /* (23, 18, 26) {real, imag} */,
  {32'h459ae79e, 32'h00000000} /* (23, 18, 25) {real, imag} */,
  {32'h45a145dc, 32'h00000000} /* (23, 18, 24) {real, imag} */,
  {32'h459188fb, 32'h00000000} /* (23, 18, 23) {real, imag} */,
  {32'h4539c8ba, 32'h00000000} /* (23, 18, 22) {real, imag} */,
  {32'h448d74fc, 32'h00000000} /* (23, 18, 21) {real, imag} */,
  {32'hc511fbb1, 32'h00000000} /* (23, 18, 20) {real, imag} */,
  {32'hc5a2b922, 32'h00000000} /* (23, 18, 19) {real, imag} */,
  {32'hc5ac174d, 32'h00000000} /* (23, 18, 18) {real, imag} */,
  {32'hc59282ce, 32'h00000000} /* (23, 18, 17) {real, imag} */,
  {32'hc5984782, 32'h00000000} /* (23, 18, 16) {real, imag} */,
  {32'hc59e0342, 32'h00000000} /* (23, 18, 15) {real, imag} */,
  {32'hc5af3a48, 32'h00000000} /* (23, 18, 14) {real, imag} */,
  {32'hc5a3ea2d, 32'h00000000} /* (23, 18, 13) {real, imag} */,
  {32'hc577cab9, 32'h00000000} /* (23, 18, 12) {real, imag} */,
  {32'hc527cdde, 32'h00000000} /* (23, 18, 11) {real, imag} */,
  {32'h443efd68, 32'h00000000} /* (23, 18, 10) {real, imag} */,
  {32'h451114a9, 32'h00000000} /* (23, 18, 9) {real, imag} */,
  {32'h457e1e0f, 32'h00000000} /* (23, 18, 8) {real, imag} */,
  {32'h45a0481d, 32'h00000000} /* (23, 18, 7) {real, imag} */,
  {32'h45a91703, 32'h00000000} /* (23, 18, 6) {real, imag} */,
  {32'h45bc71bb, 32'h00000000} /* (23, 18, 5) {real, imag} */,
  {32'h45bc137c, 32'h00000000} /* (23, 18, 4) {real, imag} */,
  {32'h45ae3bfc, 32'h00000000} /* (23, 18, 3) {real, imag} */,
  {32'h45b47ecb, 32'h00000000} /* (23, 18, 2) {real, imag} */,
  {32'h45d3c8e8, 32'h00000000} /* (23, 18, 1) {real, imag} */,
  {32'h45b316be, 32'h00000000} /* (23, 18, 0) {real, imag} */,
  {32'h45ee16e8, 32'h00000000} /* (23, 17, 31) {real, imag} */,
  {32'h45e5497b, 32'h00000000} /* (23, 17, 30) {real, imag} */,
  {32'h45d53306, 32'h00000000} /* (23, 17, 29) {real, imag} */,
  {32'h45ed3c4c, 32'h00000000} /* (23, 17, 28) {real, imag} */,
  {32'h45af4bb3, 32'h00000000} /* (23, 17, 27) {real, imag} */,
  {32'h45adf326, 32'h00000000} /* (23, 17, 26) {real, imag} */,
  {32'h45c28154, 32'h00000000} /* (23, 17, 25) {real, imag} */,
  {32'h45b9ff10, 32'h00000000} /* (23, 17, 24) {real, imag} */,
  {32'h45996c5a, 32'h00000000} /* (23, 17, 23) {real, imag} */,
  {32'h45440c81, 32'h00000000} /* (23, 17, 22) {real, imag} */,
  {32'h444e81e8, 32'h00000000} /* (23, 17, 21) {real, imag} */,
  {32'hc54ddac5, 32'h00000000} /* (23, 17, 20) {real, imag} */,
  {32'hc591e19c, 32'h00000000} /* (23, 17, 19) {real, imag} */,
  {32'hc5c04a4f, 32'h00000000} /* (23, 17, 18) {real, imag} */,
  {32'hc5cd6404, 32'h00000000} /* (23, 17, 17) {real, imag} */,
  {32'hc5be2b60, 32'h00000000} /* (23, 17, 16) {real, imag} */,
  {32'hc5d122c0, 32'h00000000} /* (23, 17, 15) {real, imag} */,
  {32'hc5ceaa7b, 32'h00000000} /* (23, 17, 14) {real, imag} */,
  {32'hc5acd4b8, 32'h00000000} /* (23, 17, 13) {real, imag} */,
  {32'hc59916ce, 32'h00000000} /* (23, 17, 12) {real, imag} */,
  {32'hc5641c2a, 32'h00000000} /* (23, 17, 11) {real, imag} */,
  {32'hc3f15fe8, 32'h00000000} /* (23, 17, 10) {real, imag} */,
  {32'h4543de00, 32'h00000000} /* (23, 17, 9) {real, imag} */,
  {32'h459d6220, 32'h00000000} /* (23, 17, 8) {real, imag} */,
  {32'h45ab43fc, 32'h00000000} /* (23, 17, 7) {real, imag} */,
  {32'h45cbbea0, 32'h00000000} /* (23, 17, 6) {real, imag} */,
  {32'h45cd1534, 32'h00000000} /* (23, 17, 5) {real, imag} */,
  {32'h45c7fafe, 32'h00000000} /* (23, 17, 4) {real, imag} */,
  {32'h45d87fd8, 32'h00000000} /* (23, 17, 3) {real, imag} */,
  {32'h45d8fb5f, 32'h00000000} /* (23, 17, 2) {real, imag} */,
  {32'h45e8a270, 32'h00000000} /* (23, 17, 1) {real, imag} */,
  {32'h45dbb75a, 32'h00000000} /* (23, 17, 0) {real, imag} */,
  {32'h45e441a9, 32'h00000000} /* (23, 16, 31) {real, imag} */,
  {32'h45f3cdd4, 32'h00000000} /* (23, 16, 30) {real, imag} */,
  {32'h45fd2ba4, 32'h00000000} /* (23, 16, 29) {real, imag} */,
  {32'h45d736ae, 32'h00000000} /* (23, 16, 28) {real, imag} */,
  {32'h45de1a06, 32'h00000000} /* (23, 16, 27) {real, imag} */,
  {32'h45ca8312, 32'h00000000} /* (23, 16, 26) {real, imag} */,
  {32'h45dfb682, 32'h00000000} /* (23, 16, 25) {real, imag} */,
  {32'h45c86294, 32'h00000000} /* (23, 16, 24) {real, imag} */,
  {32'h45b84164, 32'h00000000} /* (23, 16, 23) {real, imag} */,
  {32'h4577ddd0, 32'h00000000} /* (23, 16, 22) {real, imag} */,
  {32'h432935c0, 32'h00000000} /* (23, 16, 21) {real, imag} */,
  {32'hc53b6f32, 32'h00000000} /* (23, 16, 20) {real, imag} */,
  {32'hc58b6021, 32'h00000000} /* (23, 16, 19) {real, imag} */,
  {32'hc5b742ca, 32'h00000000} /* (23, 16, 18) {real, imag} */,
  {32'hc5cf1992, 32'h00000000} /* (23, 16, 17) {real, imag} */,
  {32'hc5d80016, 32'h00000000} /* (23, 16, 16) {real, imag} */,
  {32'hc5cb6c4f, 32'h00000000} /* (23, 16, 15) {real, imag} */,
  {32'hc5c4bde4, 32'h00000000} /* (23, 16, 14) {real, imag} */,
  {32'hc5b0e0e8, 32'h00000000} /* (23, 16, 13) {real, imag} */,
  {32'hc59fb18a, 32'h00000000} /* (23, 16, 12) {real, imag} */,
  {32'hc53dc2fc, 32'h00000000} /* (23, 16, 11) {real, imag} */,
  {32'hc29b4c60, 32'h00000000} /* (23, 16, 10) {real, imag} */,
  {32'h457a6a34, 32'h00000000} /* (23, 16, 9) {real, imag} */,
  {32'h459618a4, 32'h00000000} /* (23, 16, 8) {real, imag} */,
  {32'h45b492d0, 32'h00000000} /* (23, 16, 7) {real, imag} */,
  {32'h45be40ac, 32'h00000000} /* (23, 16, 6) {real, imag} */,
  {32'h45e3041c, 32'h00000000} /* (23, 16, 5) {real, imag} */,
  {32'h45f7a1dd, 32'h00000000} /* (23, 16, 4) {real, imag} */,
  {32'h45e3ba0f, 32'h00000000} /* (23, 16, 3) {real, imag} */,
  {32'h4604b9b3, 32'h00000000} /* (23, 16, 2) {real, imag} */,
  {32'h45fc64fe, 32'h00000000} /* (23, 16, 1) {real, imag} */,
  {32'h45dde128, 32'h00000000} /* (23, 16, 0) {real, imag} */,
  {32'h45e0bf6c, 32'h00000000} /* (23, 15, 31) {real, imag} */,
  {32'h45eda11f, 32'h00000000} /* (23, 15, 30) {real, imag} */,
  {32'h45ffcef2, 32'h00000000} /* (23, 15, 29) {real, imag} */,
  {32'h45db337e, 32'h00000000} /* (23, 15, 28) {real, imag} */,
  {32'h46000ed2, 32'h00000000} /* (23, 15, 27) {real, imag} */,
  {32'h45fbd2cf, 32'h00000000} /* (23, 15, 26) {real, imag} */,
  {32'h45c8b4df, 32'h00000000} /* (23, 15, 25) {real, imag} */,
  {32'h45bd4520, 32'h00000000} /* (23, 15, 24) {real, imag} */,
  {32'h45a8d6b0, 32'h00000000} /* (23, 15, 23) {real, imag} */,
  {32'h45438428, 32'h00000000} /* (23, 15, 22) {real, imag} */,
  {32'hc2edaba0, 32'h00000000} /* (23, 15, 21) {real, imag} */,
  {32'hc57cbeac, 32'h00000000} /* (23, 15, 20) {real, imag} */,
  {32'hc5885945, 32'h00000000} /* (23, 15, 19) {real, imag} */,
  {32'hc5c9ef39, 32'h00000000} /* (23, 15, 18) {real, imag} */,
  {32'hc5ce2660, 32'h00000000} /* (23, 15, 17) {real, imag} */,
  {32'hc5d0a91a, 32'h00000000} /* (23, 15, 16) {real, imag} */,
  {32'hc5c1de26, 32'h00000000} /* (23, 15, 15) {real, imag} */,
  {32'hc5a6ccd1, 32'h00000000} /* (23, 15, 14) {real, imag} */,
  {32'hc5c87bd6, 32'h00000000} /* (23, 15, 13) {real, imag} */,
  {32'hc5a66762, 32'h00000000} /* (23, 15, 12) {real, imag} */,
  {32'hc503c996, 32'h00000000} /* (23, 15, 11) {real, imag} */,
  {32'h43d32ff0, 32'h00000000} /* (23, 15, 10) {real, imag} */,
  {32'h45480656, 32'h00000000} /* (23, 15, 9) {real, imag} */,
  {32'h459f7704, 32'h00000000} /* (23, 15, 8) {real, imag} */,
  {32'h45c0c464, 32'h00000000} /* (23, 15, 7) {real, imag} */,
  {32'h45d97158, 32'h00000000} /* (23, 15, 6) {real, imag} */,
  {32'h45e9be3a, 32'h00000000} /* (23, 15, 5) {real, imag} */,
  {32'h45fa73ea, 32'h00000000} /* (23, 15, 4) {real, imag} */,
  {32'h460107b6, 32'h00000000} /* (23, 15, 3) {real, imag} */,
  {32'h45fc3795, 32'h00000000} /* (23, 15, 2) {real, imag} */,
  {32'h45e8cdf8, 32'h00000000} /* (23, 15, 1) {real, imag} */,
  {32'h45e64730, 32'h00000000} /* (23, 15, 0) {real, imag} */,
  {32'h45d26627, 32'h00000000} /* (23, 14, 31) {real, imag} */,
  {32'h45df279a, 32'h00000000} /* (23, 14, 30) {real, imag} */,
  {32'h45d8d58a, 32'h00000000} /* (23, 14, 29) {real, imag} */,
  {32'h45e1ab9e, 32'h00000000} /* (23, 14, 28) {real, imag} */,
  {32'h45d28541, 32'h00000000} /* (23, 14, 27) {real, imag} */,
  {32'h45c1b496, 32'h00000000} /* (23, 14, 26) {real, imag} */,
  {32'h45b64c34, 32'h00000000} /* (23, 14, 25) {real, imag} */,
  {32'h45d6ac08, 32'h00000000} /* (23, 14, 24) {real, imag} */,
  {32'h45aeeb55, 32'h00000000} /* (23, 14, 23) {real, imag} */,
  {32'h45398374, 32'h00000000} /* (23, 14, 22) {real, imag} */,
  {32'h41f78a80, 32'h00000000} /* (23, 14, 21) {real, imag} */,
  {32'hc5339e27, 32'h00000000} /* (23, 14, 20) {real, imag} */,
  {32'hc596e14c, 32'h00000000} /* (23, 14, 19) {real, imag} */,
  {32'hc5aedcdb, 32'h00000000} /* (23, 14, 18) {real, imag} */,
  {32'hc5c172c0, 32'h00000000} /* (23, 14, 17) {real, imag} */,
  {32'hc5b7cb90, 32'h00000000} /* (23, 14, 16) {real, imag} */,
  {32'hc5a93481, 32'h00000000} /* (23, 14, 15) {real, imag} */,
  {32'hc5b220fe, 32'h00000000} /* (23, 14, 14) {real, imag} */,
  {32'hc59226ac, 32'h00000000} /* (23, 14, 13) {real, imag} */,
  {32'hc57a5661, 32'h00000000} /* (23, 14, 12) {real, imag} */,
  {32'hc515d63e, 32'h00000000} /* (23, 14, 11) {real, imag} */,
  {32'h44a4dcce, 32'h00000000} /* (23, 14, 10) {real, imag} */,
  {32'h456e95ef, 32'h00000000} /* (23, 14, 9) {real, imag} */,
  {32'h45c79130, 32'h00000000} /* (23, 14, 8) {real, imag} */,
  {32'h45dd3b13, 32'h00000000} /* (23, 14, 7) {real, imag} */,
  {32'h45cf98f6, 32'h00000000} /* (23, 14, 6) {real, imag} */,
  {32'h45e6c580, 32'h00000000} /* (23, 14, 5) {real, imag} */,
  {32'h45f582e8, 32'h00000000} /* (23, 14, 4) {real, imag} */,
  {32'h45f21078, 32'h00000000} /* (23, 14, 3) {real, imag} */,
  {32'h45cdcdf5, 32'h00000000} /* (23, 14, 2) {real, imag} */,
  {32'h45d3879a, 32'h00000000} /* (23, 14, 1) {real, imag} */,
  {32'h45de609c, 32'h00000000} /* (23, 14, 0) {real, imag} */,
  {32'h45a92a26, 32'h00000000} /* (23, 13, 31) {real, imag} */,
  {32'h45a0c85e, 32'h00000000} /* (23, 13, 30) {real, imag} */,
  {32'h45c80204, 32'h00000000} /* (23, 13, 29) {real, imag} */,
  {32'h45c2371f, 32'h00000000} /* (23, 13, 28) {real, imag} */,
  {32'h45c29818, 32'h00000000} /* (23, 13, 27) {real, imag} */,
  {32'h45a17c24, 32'h00000000} /* (23, 13, 26) {real, imag} */,
  {32'h4597c414, 32'h00000000} /* (23, 13, 25) {real, imag} */,
  {32'h45ab98ff, 32'h00000000} /* (23, 13, 24) {real, imag} */,
  {32'h45a3b70c, 32'h00000000} /* (23, 13, 23) {real, imag} */,
  {32'h45530360, 32'h00000000} /* (23, 13, 22) {real, imag} */,
  {32'h44320920, 32'h00000000} /* (23, 13, 21) {real, imag} */,
  {32'hc533380e, 32'h00000000} /* (23, 13, 20) {real, imag} */,
  {32'hc59cb867, 32'h00000000} /* (23, 13, 19) {real, imag} */,
  {32'hc59f0372, 32'h00000000} /* (23, 13, 18) {real, imag} */,
  {32'hc5bca14e, 32'h00000000} /* (23, 13, 17) {real, imag} */,
  {32'hc5a07f19, 32'h00000000} /* (23, 13, 16) {real, imag} */,
  {32'hc58f9716, 32'h00000000} /* (23, 13, 15) {real, imag} */,
  {32'hc584bbd2, 32'h00000000} /* (23, 13, 14) {real, imag} */,
  {32'hc59a27a0, 32'h00000000} /* (23, 13, 13) {real, imag} */,
  {32'hc57a7986, 32'h00000000} /* (23, 13, 12) {real, imag} */,
  {32'hc4a8a886, 32'h00000000} /* (23, 13, 11) {real, imag} */,
  {32'h44a0d26c, 32'h00000000} /* (23, 13, 10) {real, imag} */,
  {32'h458cf7b4, 32'h00000000} /* (23, 13, 9) {real, imag} */,
  {32'h45a02199, 32'h00000000} /* (23, 13, 8) {real, imag} */,
  {32'h45c8c930, 32'h00000000} /* (23, 13, 7) {real, imag} */,
  {32'h45d710ae, 32'h00000000} /* (23, 13, 6) {real, imag} */,
  {32'h45cb6a24, 32'h00000000} /* (23, 13, 5) {real, imag} */,
  {32'h45cddd3d, 32'h00000000} /* (23, 13, 4) {real, imag} */,
  {32'h45b4ea47, 32'h00000000} /* (23, 13, 3) {real, imag} */,
  {32'h45916dd2, 32'h00000000} /* (23, 13, 2) {real, imag} */,
  {32'h45b1dc2e, 32'h00000000} /* (23, 13, 1) {real, imag} */,
  {32'h45b22b4f, 32'h00000000} /* (23, 13, 0) {real, imag} */,
  {32'h457b6285, 32'h00000000} /* (23, 12, 31) {real, imag} */,
  {32'h457db717, 32'h00000000} /* (23, 12, 30) {real, imag} */,
  {32'h4581c7d4, 32'h00000000} /* (23, 12, 29) {real, imag} */,
  {32'h4592c6cb, 32'h00000000} /* (23, 12, 28) {real, imag} */,
  {32'h457da625, 32'h00000000} /* (23, 12, 27) {real, imag} */,
  {32'h45980480, 32'h00000000} /* (23, 12, 26) {real, imag} */,
  {32'h4552fb5e, 32'h00000000} /* (23, 12, 25) {real, imag} */,
  {32'h4542648e, 32'h00000000} /* (23, 12, 24) {real, imag} */,
  {32'h4539d7a1, 32'h00000000} /* (23, 12, 23) {real, imag} */,
  {32'h453423f1, 32'h00000000} /* (23, 12, 22) {real, imag} */,
  {32'hc2dec040, 32'h00000000} /* (23, 12, 21) {real, imag} */,
  {32'hc536f038, 32'h00000000} /* (23, 12, 20) {real, imag} */,
  {32'hc5815d80, 32'h00000000} /* (23, 12, 19) {real, imag} */,
  {32'hc5a8c38b, 32'h00000000} /* (23, 12, 18) {real, imag} */,
  {32'hc5b6b2b2, 32'h00000000} /* (23, 12, 17) {real, imag} */,
  {32'hc592ce49, 32'h00000000} /* (23, 12, 16) {real, imag} */,
  {32'hc56895d1, 32'h00000000} /* (23, 12, 15) {real, imag} */,
  {32'hc53dea4f, 32'h00000000} /* (23, 12, 14) {real, imag} */,
  {32'hc56f5bc1, 32'h00000000} /* (23, 12, 13) {real, imag} */,
  {32'hc5457b15, 32'h00000000} /* (23, 12, 12) {real, imag} */,
  {32'hc506d4d5, 32'h00000000} /* (23, 12, 11) {real, imag} */,
  {32'h44c5dbd7, 32'h00000000} /* (23, 12, 10) {real, imag} */,
  {32'h457c3212, 32'h00000000} /* (23, 12, 9) {real, imag} */,
  {32'h45a4561f, 32'h00000000} /* (23, 12, 8) {real, imag} */,
  {32'h45a5981e, 32'h00000000} /* (23, 12, 7) {real, imag} */,
  {32'h45a75cba, 32'h00000000} /* (23, 12, 6) {real, imag} */,
  {32'h45aed305, 32'h00000000} /* (23, 12, 5) {real, imag} */,
  {32'h45918122, 32'h00000000} /* (23, 12, 4) {real, imag} */,
  {32'h45914b88, 32'h00000000} /* (23, 12, 3) {real, imag} */,
  {32'h45941387, 32'h00000000} /* (23, 12, 2) {real, imag} */,
  {32'h45864818, 32'h00000000} /* (23, 12, 1) {real, imag} */,
  {32'h45703252, 32'h00000000} /* (23, 12, 0) {real, imag} */,
  {32'h4499c836, 32'h00000000} /* (23, 11, 31) {real, imag} */,
  {32'h44ddabd6, 32'h00000000} /* (23, 11, 30) {real, imag} */,
  {32'h44df120d, 32'h00000000} /* (23, 11, 29) {real, imag} */,
  {32'h4535adb8, 32'h00000000} /* (23, 11, 28) {real, imag} */,
  {32'h45187a17, 32'h00000000} /* (23, 11, 27) {real, imag} */,
  {32'h44f17073, 32'h00000000} /* (23, 11, 26) {real, imag} */,
  {32'h44ee8070, 32'h00000000} /* (23, 11, 25) {real, imag} */,
  {32'h44e01698, 32'h00000000} /* (23, 11, 24) {real, imag} */,
  {32'h4499c37e, 32'h00000000} /* (23, 11, 23) {real, imag} */,
  {32'h43f23528, 32'h00000000} /* (23, 11, 22) {real, imag} */,
  {32'hc4855a71, 32'h00000000} /* (23, 11, 21) {real, imag} */,
  {32'hc51b3211, 32'h00000000} /* (23, 11, 20) {real, imag} */,
  {32'hc5584d95, 32'h00000000} /* (23, 11, 19) {real, imag} */,
  {32'hc51b3784, 32'h00000000} /* (23, 11, 18) {real, imag} */,
  {32'hc5430f9a, 32'h00000000} /* (23, 11, 17) {real, imag} */,
  {32'hc51ec09a, 32'h00000000} /* (23, 11, 16) {real, imag} */,
  {32'hc507bb3b, 32'h00000000} /* (23, 11, 15) {real, imag} */,
  {32'hc4e5f9b0, 32'h00000000} /* (23, 11, 14) {real, imag} */,
  {32'hc4d52f15, 32'h00000000} /* (23, 11, 13) {real, imag} */,
  {32'hc504fc80, 32'h00000000} /* (23, 11, 12) {real, imag} */,
  {32'hc445e3a8, 32'h00000000} /* (23, 11, 11) {real, imag} */,
  {32'h448fabad, 32'h00000000} /* (23, 11, 10) {real, imag} */,
  {32'h4524ecb8, 32'h00000000} /* (23, 11, 9) {real, imag} */,
  {32'h452f2520, 32'h00000000} /* (23, 11, 8) {real, imag} */,
  {32'h45413b57, 32'h00000000} /* (23, 11, 7) {real, imag} */,
  {32'h454a7ca5, 32'h00000000} /* (23, 11, 6) {real, imag} */,
  {32'h44fa130f, 32'h00000000} /* (23, 11, 5) {real, imag} */,
  {32'h452725a1, 32'h00000000} /* (23, 11, 4) {real, imag} */,
  {32'h44f5e5b2, 32'h00000000} /* (23, 11, 3) {real, imag} */,
  {32'h4502c0a6, 32'h00000000} /* (23, 11, 2) {real, imag} */,
  {32'h44a4d50c, 32'h00000000} /* (23, 11, 1) {real, imag} */,
  {32'h4457be5a, 32'h00000000} /* (23, 11, 0) {real, imag} */,
  {32'hc510baa9, 32'h00000000} /* (23, 10, 31) {real, imag} */,
  {32'hc50c9a15, 32'h00000000} /* (23, 10, 30) {real, imag} */,
  {32'hc50cd309, 32'h00000000} /* (23, 10, 29) {real, imag} */,
  {32'hc5015ff8, 32'h00000000} /* (23, 10, 28) {real, imag} */,
  {32'hc513d26a, 32'h00000000} /* (23, 10, 27) {real, imag} */,
  {32'hc4d4a0b5, 32'h00000000} /* (23, 10, 26) {real, imag} */,
  {32'hc442dd44, 32'h00000000} /* (23, 10, 25) {real, imag} */,
  {32'hc463fd26, 32'h00000000} /* (23, 10, 24) {real, imag} */,
  {32'hc55ebe6c, 32'h00000000} /* (23, 10, 23) {real, imag} */,
  {32'hc5281c90, 32'h00000000} /* (23, 10, 22) {real, imag} */,
  {32'hc514a55a, 32'h00000000} /* (23, 10, 21) {real, imag} */,
  {32'hc4e97ad7, 32'h00000000} /* (23, 10, 20) {real, imag} */,
  {32'hc4a0562a, 32'h00000000} /* (23, 10, 19) {real, imag} */,
  {32'hc0e5dd80, 32'h00000000} /* (23, 10, 18) {real, imag} */,
  {32'h4411daaa, 32'h00000000} /* (23, 10, 17) {real, imag} */,
  {32'h4498954b, 32'h00000000} /* (23, 10, 16) {real, imag} */,
  {32'h4479ea7b, 32'h00000000} /* (23, 10, 15) {real, imag} */,
  {32'h444367bb, 32'h00000000} /* (23, 10, 14) {real, imag} */,
  {32'h44936acc, 32'h00000000} /* (23, 10, 13) {real, imag} */,
  {32'h44a74535, 32'h00000000} /* (23, 10, 12) {real, imag} */,
  {32'h44988c14, 32'h00000000} /* (23, 10, 11) {real, imag} */,
  {32'h43c68dd4, 32'h00000000} /* (23, 10, 10) {real, imag} */,
  {32'h44713e1c, 32'h00000000} /* (23, 10, 9) {real, imag} */,
  {32'h44603ddc, 32'h00000000} /* (23, 10, 8) {real, imag} */,
  {32'h439417dc, 32'h00000000} /* (23, 10, 7) {real, imag} */,
  {32'hc44bb9da, 32'h00000000} /* (23, 10, 6) {real, imag} */,
  {32'hc428a6da, 32'h00000000} /* (23, 10, 5) {real, imag} */,
  {32'hc4ef269b, 32'h00000000} /* (23, 10, 4) {real, imag} */,
  {32'hc541fadd, 32'h00000000} /* (23, 10, 3) {real, imag} */,
  {32'hc4fc7440, 32'h00000000} /* (23, 10, 2) {real, imag} */,
  {32'hc509bfb4, 32'h00000000} /* (23, 10, 1) {real, imag} */,
  {32'hc4d2e20b, 32'h00000000} /* (23, 10, 0) {real, imag} */,
  {32'hc5997ee6, 32'h00000000} /* (23, 9, 31) {real, imag} */,
  {32'hc5b9804a, 32'h00000000} /* (23, 9, 30) {real, imag} */,
  {32'hc5cbca0b, 32'h00000000} /* (23, 9, 29) {real, imag} */,
  {32'hc5c08127, 32'h00000000} /* (23, 9, 28) {real, imag} */,
  {32'hc5b6ccb4, 32'h00000000} /* (23, 9, 27) {real, imag} */,
  {32'hc5a6716c, 32'h00000000} /* (23, 9, 26) {real, imag} */,
  {32'hc5b1f8da, 32'h00000000} /* (23, 9, 25) {real, imag} */,
  {32'hc5ad953f, 32'h00000000} /* (23, 9, 24) {real, imag} */,
  {32'hc59f1943, 32'h00000000} /* (23, 9, 23) {real, imag} */,
  {32'hc59bece3, 32'h00000000} /* (23, 9, 22) {real, imag} */,
  {32'hc5518b7e, 32'h00000000} /* (23, 9, 21) {real, imag} */,
  {32'hc4a60158, 32'h00000000} /* (23, 9, 20) {real, imag} */,
  {32'h42d83140, 32'h00000000} /* (23, 9, 19) {real, imag} */,
  {32'h449825d1, 32'h00000000} /* (23, 9, 18) {real, imag} */,
  {32'h451e0258, 32'h00000000} /* (23, 9, 17) {real, imag} */,
  {32'h451bd32c, 32'h00000000} /* (23, 9, 16) {real, imag} */,
  {32'h45664630, 32'h00000000} /* (23, 9, 15) {real, imag} */,
  {32'h4568d988, 32'h00000000} /* (23, 9, 14) {real, imag} */,
  {32'h455c0f1e, 32'h00000000} /* (23, 9, 13) {real, imag} */,
  {32'h454c59ea, 32'h00000000} /* (23, 9, 12) {real, imag} */,
  {32'h450a6426, 32'h00000000} /* (23, 9, 11) {real, imag} */,
  {32'hc3a1f5f0, 32'h00000000} /* (23, 9, 10) {real, imag} */,
  {32'hc447e584, 32'h00000000} /* (23, 9, 9) {real, imag} */,
  {32'hc4f2f87c, 32'h00000000} /* (23, 9, 8) {real, imag} */,
  {32'hc50b3756, 32'h00000000} /* (23, 9, 7) {real, imag} */,
  {32'hc5316be2, 32'h00000000} /* (23, 9, 6) {real, imag} */,
  {32'hc5691f32, 32'h00000000} /* (23, 9, 5) {real, imag} */,
  {32'hc55c1ac2, 32'h00000000} /* (23, 9, 4) {real, imag} */,
  {32'hc58b0513, 32'h00000000} /* (23, 9, 3) {real, imag} */,
  {32'hc5a26343, 32'h00000000} /* (23, 9, 2) {real, imag} */,
  {32'hc581df21, 32'h00000000} /* (23, 9, 1) {real, imag} */,
  {32'hc585a9fc, 32'h00000000} /* (23, 9, 0) {real, imag} */,
  {32'hc5d7268f, 32'h00000000} /* (23, 8, 31) {real, imag} */,
  {32'hc5f5dddd, 32'h00000000} /* (23, 8, 30) {real, imag} */,
  {32'hc606045c, 32'h00000000} /* (23, 8, 29) {real, imag} */,
  {32'hc60607c4, 32'h00000000} /* (23, 8, 28) {real, imag} */,
  {32'hc60b76f9, 32'h00000000} /* (23, 8, 27) {real, imag} */,
  {32'hc603e5c5, 32'h00000000} /* (23, 8, 26) {real, imag} */,
  {32'hc5ef0771, 32'h00000000} /* (23, 8, 25) {real, imag} */,
  {32'hc602a8e0, 32'h00000000} /* (23, 8, 24) {real, imag} */,
  {32'hc5d8cbcc, 32'h00000000} /* (23, 8, 23) {real, imag} */,
  {32'hc5bccba9, 32'h00000000} /* (23, 8, 22) {real, imag} */,
  {32'hc57e7eaa, 32'h00000000} /* (23, 8, 21) {real, imag} */,
  {32'hc47decf0, 32'h00000000} /* (23, 8, 20) {real, imag} */,
  {32'h41cac780, 32'h00000000} /* (23, 8, 19) {real, imag} */,
  {32'h44cecfac, 32'h00000000} /* (23, 8, 18) {real, imag} */,
  {32'h45126a60, 32'h00000000} /* (23, 8, 17) {real, imag} */,
  {32'h456618c5, 32'h00000000} /* (23, 8, 16) {real, imag} */,
  {32'h45a4656d, 32'h00000000} /* (23, 8, 15) {real, imag} */,
  {32'h456dd686, 32'h00000000} /* (23, 8, 14) {real, imag} */,
  {32'h45964054, 32'h00000000} /* (23, 8, 13) {real, imag} */,
  {32'h45b9649d, 32'h00000000} /* (23, 8, 12) {real, imag} */,
  {32'h4545378c, 32'h00000000} /* (23, 8, 11) {real, imag} */,
  {32'h449de1c8, 32'h00000000} /* (23, 8, 10) {real, imag} */,
  {32'hc41ba8f8, 32'h00000000} /* (23, 8, 9) {real, imag} */,
  {32'hc544485f, 32'h00000000} /* (23, 8, 8) {real, imag} */,
  {32'hc58651fe, 32'h00000000} /* (23, 8, 7) {real, imag} */,
  {32'hc57b00b2, 32'h00000000} /* (23, 8, 6) {real, imag} */,
  {32'hc59e1301, 32'h00000000} /* (23, 8, 5) {real, imag} */,
  {32'hc5b577c2, 32'h00000000} /* (23, 8, 4) {real, imag} */,
  {32'hc5db81a8, 32'h00000000} /* (23, 8, 3) {real, imag} */,
  {32'hc5c27887, 32'h00000000} /* (23, 8, 2) {real, imag} */,
  {32'hc5c78526, 32'h00000000} /* (23, 8, 1) {real, imag} */,
  {32'hc5cd54de, 32'h00000000} /* (23, 8, 0) {real, imag} */,
  {32'hc6038d44, 32'h00000000} /* (23, 7, 31) {real, imag} */,
  {32'hc608c6f0, 32'h00000000} /* (23, 7, 30) {real, imag} */,
  {32'hc6110132, 32'h00000000} /* (23, 7, 29) {real, imag} */,
  {32'hc6214ce8, 32'h00000000} /* (23, 7, 28) {real, imag} */,
  {32'hc6269774, 32'h00000000} /* (23, 7, 27) {real, imag} */,
  {32'hc6221bea, 32'h00000000} /* (23, 7, 26) {real, imag} */,
  {32'hc619535f, 32'h00000000} /* (23, 7, 25) {real, imag} */,
  {32'hc60b8922, 32'h00000000} /* (23, 7, 24) {real, imag} */,
  {32'hc60ff9a6, 32'h00000000} /* (23, 7, 23) {real, imag} */,
  {32'hc5d8efc8, 32'h00000000} /* (23, 7, 22) {real, imag} */,
  {32'hc577a0f5, 32'h00000000} /* (23, 7, 21) {real, imag} */,
  {32'hc4d0c344, 32'h00000000} /* (23, 7, 20) {real, imag} */,
  {32'h438e5cc8, 32'h00000000} /* (23, 7, 19) {real, imag} */,
  {32'h448d04ba, 32'h00000000} /* (23, 7, 18) {real, imag} */,
  {32'h4539471c, 32'h00000000} /* (23, 7, 17) {real, imag} */,
  {32'h458ba0eb, 32'h00000000} /* (23, 7, 16) {real, imag} */,
  {32'h458a8e84, 32'h00000000} /* (23, 7, 15) {real, imag} */,
  {32'h459e76db, 32'h00000000} /* (23, 7, 14) {real, imag} */,
  {32'h459d175f, 32'h00000000} /* (23, 7, 13) {real, imag} */,
  {32'h45851630, 32'h00000000} /* (23, 7, 12) {real, imag} */,
  {32'h456bc6ee, 32'h00000000} /* (23, 7, 11) {real, imag} */,
  {32'h44891b74, 32'h00000000} /* (23, 7, 10) {real, imag} */,
  {32'hc47df8d0, 32'h00000000} /* (23, 7, 9) {real, imag} */,
  {32'hc528794a, 32'h00000000} /* (23, 7, 8) {real, imag} */,
  {32'hc5433ca2, 32'h00000000} /* (23, 7, 7) {real, imag} */,
  {32'hc5a7b7bc, 32'h00000000} /* (23, 7, 6) {real, imag} */,
  {32'hc5ab1c72, 32'h00000000} /* (23, 7, 5) {real, imag} */,
  {32'hc5c953af, 32'h00000000} /* (23, 7, 4) {real, imag} */,
  {32'hc5e99180, 32'h00000000} /* (23, 7, 3) {real, imag} */,
  {32'hc605bec1, 32'h00000000} /* (23, 7, 2) {real, imag} */,
  {32'hc6014a86, 32'h00000000} /* (23, 7, 1) {real, imag} */,
  {32'hc5ec593d, 32'h00000000} /* (23, 7, 0) {real, imag} */,
  {32'hc612122a, 32'h00000000} /* (23, 6, 31) {real, imag} */,
  {32'hc61de586, 32'h00000000} /* (23, 6, 30) {real, imag} */,
  {32'hc62a0b2e, 32'h00000000} /* (23, 6, 29) {real, imag} */,
  {32'hc62d8d07, 32'h00000000} /* (23, 6, 28) {real, imag} */,
  {32'hc62d54af, 32'h00000000} /* (23, 6, 27) {real, imag} */,
  {32'hc62b13e8, 32'h00000000} /* (23, 6, 26) {real, imag} */,
  {32'hc6243b93, 32'h00000000} /* (23, 6, 25) {real, imag} */,
  {32'hc61b14a2, 32'h00000000} /* (23, 6, 24) {real, imag} */,
  {32'hc60fd103, 32'h00000000} /* (23, 6, 23) {real, imag} */,
  {32'hc5fca78b, 32'h00000000} /* (23, 6, 22) {real, imag} */,
  {32'hc5b4f032, 32'h00000000} /* (23, 6, 21) {real, imag} */,
  {32'hc543e557, 32'h00000000} /* (23, 6, 20) {real, imag} */,
  {32'hc489e1f0, 32'h00000000} /* (23, 6, 19) {real, imag} */,
  {32'h4420d1b0, 32'h00000000} /* (23, 6, 18) {real, imag} */,
  {32'h450b9105, 32'h00000000} /* (23, 6, 17) {real, imag} */,
  {32'h4579f750, 32'h00000000} /* (23, 6, 16) {real, imag} */,
  {32'h458ea8c8, 32'h00000000} /* (23, 6, 15) {real, imag} */,
  {32'h45b2fdd1, 32'h00000000} /* (23, 6, 14) {real, imag} */,
  {32'h45bbbc93, 32'h00000000} /* (23, 6, 13) {real, imag} */,
  {32'h45b0858a, 32'h00000000} /* (23, 6, 12) {real, imag} */,
  {32'h459c16ae, 32'h00000000} /* (23, 6, 11) {real, imag} */,
  {32'h44ee173c, 32'h00000000} /* (23, 6, 10) {real, imag} */,
  {32'hc3327640, 32'h00000000} /* (23, 6, 9) {real, imag} */,
  {32'hc4ba4eec, 32'h00000000} /* (23, 6, 8) {real, imag} */,
  {32'hc5322ff4, 32'h00000000} /* (23, 6, 7) {real, imag} */,
  {32'hc5990f4b, 32'h00000000} /* (23, 6, 6) {real, imag} */,
  {32'hc5ad0a24, 32'h00000000} /* (23, 6, 5) {real, imag} */,
  {32'hc5d1ec24, 32'h00000000} /* (23, 6, 4) {real, imag} */,
  {32'hc5f2aa9c, 32'h00000000} /* (23, 6, 3) {real, imag} */,
  {32'hc6039d12, 32'h00000000} /* (23, 6, 2) {real, imag} */,
  {32'hc60e5eba, 32'h00000000} /* (23, 6, 1) {real, imag} */,
  {32'hc616a55a, 32'h00000000} /* (23, 6, 0) {real, imag} */,
  {32'hc628c875, 32'h00000000} /* (23, 5, 31) {real, imag} */,
  {32'hc62f68af, 32'h00000000} /* (23, 5, 30) {real, imag} */,
  {32'hc6428d85, 32'h00000000} /* (23, 5, 29) {real, imag} */,
  {32'hc6422f5d, 32'h00000000} /* (23, 5, 28) {real, imag} */,
  {32'hc63dffaa, 32'h00000000} /* (23, 5, 27) {real, imag} */,
  {32'hc6403fbd, 32'h00000000} /* (23, 5, 26) {real, imag} */,
  {32'hc6311e2e, 32'h00000000} /* (23, 5, 25) {real, imag} */,
  {32'hc62e7fcb, 32'h00000000} /* (23, 5, 24) {real, imag} */,
  {32'hc61fdb96, 32'h00000000} /* (23, 5, 23) {real, imag} */,
  {32'hc60bdb60, 32'h00000000} /* (23, 5, 22) {real, imag} */,
  {32'hc5d6f0d2, 32'h00000000} /* (23, 5, 21) {real, imag} */,
  {32'hc5a74d35, 32'h00000000} /* (23, 5, 20) {real, imag} */,
  {32'hc5593709, 32'h00000000} /* (23, 5, 19) {real, imag} */,
  {32'hc4b13866, 32'h00000000} /* (23, 5, 18) {real, imag} */,
  {32'h43b4f3d0, 32'h00000000} /* (23, 5, 17) {real, imag} */,
  {32'h44a8c384, 32'h00000000} /* (23, 5, 16) {real, imag} */,
  {32'h456a0870, 32'h00000000} /* (23, 5, 15) {real, imag} */,
  {32'h45ae82a2, 32'h00000000} /* (23, 5, 14) {real, imag} */,
  {32'h45b20e26, 32'h00000000} /* (23, 5, 13) {real, imag} */,
  {32'h45a84ece, 32'h00000000} /* (23, 5, 12) {real, imag} */,
  {32'h45a6e014, 32'h00000000} /* (23, 5, 11) {real, imag} */,
  {32'h45616b88, 32'h00000000} /* (23, 5, 10) {real, imag} */,
  {32'h45207e2e, 32'h00000000} /* (23, 5, 9) {real, imag} */,
  {32'h44928880, 32'h00000000} /* (23, 5, 8) {real, imag} */,
  {32'hc4af713c, 32'h00000000} /* (23, 5, 7) {real, imag} */,
  {32'hc5123e40, 32'h00000000} /* (23, 5, 6) {real, imag} */,
  {32'hc59fd652, 32'h00000000} /* (23, 5, 5) {real, imag} */,
  {32'hc5d99097, 32'h00000000} /* (23, 5, 4) {real, imag} */,
  {32'hc6036a5c, 32'h00000000} /* (23, 5, 3) {real, imag} */,
  {32'hc60c1a76, 32'h00000000} /* (23, 5, 2) {real, imag} */,
  {32'hc61ae5e4, 32'h00000000} /* (23, 5, 1) {real, imag} */,
  {32'hc62128de, 32'h00000000} /* (23, 5, 0) {real, imag} */,
  {32'hc6302409, 32'h00000000} /* (23, 4, 31) {real, imag} */,
  {32'hc64cddb4, 32'h00000000} /* (23, 4, 30) {real, imag} */,
  {32'hc64c632c, 32'h00000000} /* (23, 4, 29) {real, imag} */,
  {32'hc64d0c03, 32'h00000000} /* (23, 4, 28) {real, imag} */,
  {32'hc64b9946, 32'h00000000} /* (23, 4, 27) {real, imag} */,
  {32'hc64dcb98, 32'h00000000} /* (23, 4, 26) {real, imag} */,
  {32'hc64f2d9e, 32'h00000000} /* (23, 4, 25) {real, imag} */,
  {32'hc644f5a6, 32'h00000000} /* (23, 4, 24) {real, imag} */,
  {32'hc627a868, 32'h00000000} /* (23, 4, 23) {real, imag} */,
  {32'hc613eb7e, 32'h00000000} /* (23, 4, 22) {real, imag} */,
  {32'hc5e7b5d6, 32'h00000000} /* (23, 4, 21) {real, imag} */,
  {32'hc5dea278, 32'h00000000} /* (23, 4, 20) {real, imag} */,
  {32'hc5a73730, 32'h00000000} /* (23, 4, 19) {real, imag} */,
  {32'hc51fab83, 32'h00000000} /* (23, 4, 18) {real, imag} */,
  {32'hc4b6e6e0, 32'h00000000} /* (23, 4, 17) {real, imag} */,
  {32'h441a65b8, 32'h00000000} /* (23, 4, 16) {real, imag} */,
  {32'h45476e6c, 32'h00000000} /* (23, 4, 15) {real, imag} */,
  {32'h458d1175, 32'h00000000} /* (23, 4, 14) {real, imag} */,
  {32'h45c06f88, 32'h00000000} /* (23, 4, 13) {real, imag} */,
  {32'h45ade4d6, 32'h00000000} /* (23, 4, 12) {real, imag} */,
  {32'h45995389, 32'h00000000} /* (23, 4, 11) {real, imag} */,
  {32'h459d2a61, 32'h00000000} /* (23, 4, 10) {real, imag} */,
  {32'h456eea18, 32'h00000000} /* (23, 4, 9) {real, imag} */,
  {32'h4515ee32, 32'h00000000} /* (23, 4, 8) {real, imag} */,
  {32'h449869d4, 32'h00000000} /* (23, 4, 7) {real, imag} */,
  {32'hc4047648, 32'h00000000} /* (23, 4, 6) {real, imag} */,
  {32'hc58bb272, 32'h00000000} /* (23, 4, 5) {real, imag} */,
  {32'hc5e3eee4, 32'h00000000} /* (23, 4, 4) {real, imag} */,
  {32'hc61045a3, 32'h00000000} /* (23, 4, 3) {real, imag} */,
  {32'hc614a6c0, 32'h00000000} /* (23, 4, 2) {real, imag} */,
  {32'hc61d3c90, 32'h00000000} /* (23, 4, 1) {real, imag} */,
  {32'hc61dd9d0, 32'h00000000} /* (23, 4, 0) {real, imag} */,
  {32'hc6374314, 32'h00000000} /* (23, 3, 31) {real, imag} */,
  {32'hc6582adc, 32'h00000000} /* (23, 3, 30) {real, imag} */,
  {32'hc64cb08d, 32'h00000000} /* (23, 3, 29) {real, imag} */,
  {32'hc650284f, 32'h00000000} /* (23, 3, 28) {real, imag} */,
  {32'hc64c17a0, 32'h00000000} /* (23, 3, 27) {real, imag} */,
  {32'hc64732a5, 32'h00000000} /* (23, 3, 26) {real, imag} */,
  {32'hc644d2f6, 32'h00000000} /* (23, 3, 25) {real, imag} */,
  {32'hc6384958, 32'h00000000} /* (23, 3, 24) {real, imag} */,
  {32'hc6273824, 32'h00000000} /* (23, 3, 23) {real, imag} */,
  {32'hc613cd54, 32'h00000000} /* (23, 3, 22) {real, imag} */,
  {32'hc5f4638c, 32'h00000000} /* (23, 3, 21) {real, imag} */,
  {32'hc5dccf02, 32'h00000000} /* (23, 3, 20) {real, imag} */,
  {32'hc5a6e327, 32'h00000000} /* (23, 3, 19) {real, imag} */,
  {32'hc59bc94e, 32'h00000000} /* (23, 3, 18) {real, imag} */,
  {32'hc5034f4e, 32'h00000000} /* (23, 3, 17) {real, imag} */,
  {32'hc3dadb30, 32'h00000000} /* (23, 3, 16) {real, imag} */,
  {32'h456218a0, 32'h00000000} /* (23, 3, 15) {real, imag} */,
  {32'h45b34725, 32'h00000000} /* (23, 3, 14) {real, imag} */,
  {32'h45b873fa, 32'h00000000} /* (23, 3, 13) {real, imag} */,
  {32'h45c806fe, 32'h00000000} /* (23, 3, 12) {real, imag} */,
  {32'h45c1e7d8, 32'h00000000} /* (23, 3, 11) {real, imag} */,
  {32'h45b13f6e, 32'h00000000} /* (23, 3, 10) {real, imag} */,
  {32'h45739852, 32'h00000000} /* (23, 3, 9) {real, imag} */,
  {32'h45252042, 32'h00000000} /* (23, 3, 8) {real, imag} */,
  {32'h44e0f56c, 32'h00000000} /* (23, 3, 7) {real, imag} */,
  {32'hc3c9e0f0, 32'h00000000} /* (23, 3, 6) {real, imag} */,
  {32'hc5639029, 32'h00000000} /* (23, 3, 5) {real, imag} */,
  {32'hc5ebf69a, 32'h00000000} /* (23, 3, 4) {real, imag} */,
  {32'hc611c766, 32'h00000000} /* (23, 3, 3) {real, imag} */,
  {32'hc62b82c7, 32'h00000000} /* (23, 3, 2) {real, imag} */,
  {32'hc6237614, 32'h00000000} /* (23, 3, 1) {real, imag} */,
  {32'hc632a74a, 32'h00000000} /* (23, 3, 0) {real, imag} */,
  {32'hc6357986, 32'h00000000} /* (23, 2, 31) {real, imag} */,
  {32'hc636f0d4, 32'h00000000} /* (23, 2, 30) {real, imag} */,
  {32'hc652a698, 32'h00000000} /* (23, 2, 29) {real, imag} */,
  {32'hc65b6b1c, 32'h00000000} /* (23, 2, 28) {real, imag} */,
  {32'hc650072c, 32'h00000000} /* (23, 2, 27) {real, imag} */,
  {32'hc6595f68, 32'h00000000} /* (23, 2, 26) {real, imag} */,
  {32'hc6464ecc, 32'h00000000} /* (23, 2, 25) {real, imag} */,
  {32'hc6378268, 32'h00000000} /* (23, 2, 24) {real, imag} */,
  {32'hc623546c, 32'h00000000} /* (23, 2, 23) {real, imag} */,
  {32'hc6262c93, 32'h00000000} /* (23, 2, 22) {real, imag} */,
  {32'hc6060fc2, 32'h00000000} /* (23, 2, 21) {real, imag} */,
  {32'hc5db3ae1, 32'h00000000} /* (23, 2, 20) {real, imag} */,
  {32'hc5bd8be0, 32'h00000000} /* (23, 2, 19) {real, imag} */,
  {32'hc58902c6, 32'h00000000} /* (23, 2, 18) {real, imag} */,
  {32'hc527fccf, 32'h00000000} /* (23, 2, 17) {real, imag} */,
  {32'hc4a665fc, 32'h00000000} /* (23, 2, 16) {real, imag} */,
  {32'h44ff9444, 32'h00000000} /* (23, 2, 15) {real, imag} */,
  {32'h45a9b8c9, 32'h00000000} /* (23, 2, 14) {real, imag} */,
  {32'h45ce9c48, 32'h00000000} /* (23, 2, 13) {real, imag} */,
  {32'h45b12c07, 32'h00000000} /* (23, 2, 12) {real, imag} */,
  {32'h45c16b8f, 32'h00000000} /* (23, 2, 11) {real, imag} */,
  {32'h45918ded, 32'h00000000} /* (23, 2, 10) {real, imag} */,
  {32'h456ac5f0, 32'h00000000} /* (23, 2, 9) {real, imag} */,
  {32'h450e59c4, 32'h00000000} /* (23, 2, 8) {real, imag} */,
  {32'h4425f268, 32'h00000000} /* (23, 2, 7) {real, imag} */,
  {32'h439b8b00, 32'h00000000} /* (23, 2, 6) {real, imag} */,
  {32'hc584c86c, 32'h00000000} /* (23, 2, 5) {real, imag} */,
  {32'hc5dee36d, 32'h00000000} /* (23, 2, 4) {real, imag} */,
  {32'hc60faec7, 32'h00000000} /* (23, 2, 3) {real, imag} */,
  {32'hc6283e0a, 32'h00000000} /* (23, 2, 2) {real, imag} */,
  {32'hc61f5438, 32'h00000000} /* (23, 2, 1) {real, imag} */,
  {32'hc62cbaba, 32'h00000000} /* (23, 2, 0) {real, imag} */,
  {32'hc6298b98, 32'h00000000} /* (23, 1, 31) {real, imag} */,
  {32'hc6383f72, 32'h00000000} /* (23, 1, 30) {real, imag} */,
  {32'hc64a030f, 32'h00000000} /* (23, 1, 29) {real, imag} */,
  {32'hc64ae64e, 32'h00000000} /* (23, 1, 28) {real, imag} */,
  {32'hc65cf8fe, 32'h00000000} /* (23, 1, 27) {real, imag} */,
  {32'hc6520041, 32'h00000000} /* (23, 1, 26) {real, imag} */,
  {32'hc63c36a8, 32'h00000000} /* (23, 1, 25) {real, imag} */,
  {32'hc62f9ce2, 32'h00000000} /* (23, 1, 24) {real, imag} */,
  {32'hc61d42cb, 32'h00000000} /* (23, 1, 23) {real, imag} */,
  {32'hc6091c01, 32'h00000000} /* (23, 1, 22) {real, imag} */,
  {32'hc5debc90, 32'h00000000} /* (23, 1, 21) {real, imag} */,
  {32'hc5bc6d33, 32'h00000000} /* (23, 1, 20) {real, imag} */,
  {32'hc594e576, 32'h00000000} /* (23, 1, 19) {real, imag} */,
  {32'hc5486db9, 32'h00000000} /* (23, 1, 18) {real, imag} */,
  {32'hc4edfc00, 32'h00000000} /* (23, 1, 17) {real, imag} */,
  {32'hc3dca380, 32'h00000000} /* (23, 1, 16) {real, imag} */,
  {32'h453598fa, 32'h00000000} /* (23, 1, 15) {real, imag} */,
  {32'h45990715, 32'h00000000} /* (23, 1, 14) {real, imag} */,
  {32'h45b4767a, 32'h00000000} /* (23, 1, 13) {real, imag} */,
  {32'h45cafe50, 32'h00000000} /* (23, 1, 12) {real, imag} */,
  {32'h45b0016b, 32'h00000000} /* (23, 1, 11) {real, imag} */,
  {32'h456535f4, 32'h00000000} /* (23, 1, 10) {real, imag} */,
  {32'h455c60c8, 32'h00000000} /* (23, 1, 9) {real, imag} */,
  {32'h4550db70, 32'h00000000} /* (23, 1, 8) {real, imag} */,
  {32'h4410ecb0, 32'h00000000} /* (23, 1, 7) {real, imag} */,
  {32'hc4680584, 32'h00000000} /* (23, 1, 6) {real, imag} */,
  {32'hc593d2e0, 32'h00000000} /* (23, 1, 5) {real, imag} */,
  {32'hc5d4b235, 32'h00000000} /* (23, 1, 4) {real, imag} */,
  {32'hc60a0b0e, 32'h00000000} /* (23, 1, 3) {real, imag} */,
  {32'hc61075f2, 32'h00000000} /* (23, 1, 2) {real, imag} */,
  {32'hc61f93cc, 32'h00000000} /* (23, 1, 1) {real, imag} */,
  {32'hc621de38, 32'h00000000} /* (23, 1, 0) {real, imag} */,
  {32'hc62a5a3e, 32'h00000000} /* (23, 0, 31) {real, imag} */,
  {32'hc638d1fd, 32'h00000000} /* (23, 0, 30) {real, imag} */,
  {32'hc641f37a, 32'h00000000} /* (23, 0, 29) {real, imag} */,
  {32'hc63ebab0, 32'h00000000} /* (23, 0, 28) {real, imag} */,
  {32'hc64e9d1b, 32'h00000000} /* (23, 0, 27) {real, imag} */,
  {32'hc6496d4c, 32'h00000000} /* (23, 0, 26) {real, imag} */,
  {32'hc63266c6, 32'h00000000} /* (23, 0, 25) {real, imag} */,
  {32'hc62ab3ce, 32'h00000000} /* (23, 0, 24) {real, imag} */,
  {32'hc617e8b9, 32'h00000000} /* (23, 0, 23) {real, imag} */,
  {32'hc5e42ff0, 32'h00000000} /* (23, 0, 22) {real, imag} */,
  {32'hc5bb1348, 32'h00000000} /* (23, 0, 21) {real, imag} */,
  {32'hc5a09eaa, 32'h00000000} /* (23, 0, 20) {real, imag} */,
  {32'hc53a324a, 32'h00000000} /* (23, 0, 19) {real, imag} */,
  {32'hc4e97580, 32'h00000000} /* (23, 0, 18) {real, imag} */,
  {32'hc3a80c40, 32'h00000000} /* (23, 0, 17) {real, imag} */,
  {32'h44efc9b8, 32'h00000000} /* (23, 0, 16) {real, imag} */,
  {32'h4573dc4e, 32'h00000000} /* (23, 0, 15) {real, imag} */,
  {32'h45982d9a, 32'h00000000} /* (23, 0, 14) {real, imag} */,
  {32'h459b2bb4, 32'h00000000} /* (23, 0, 13) {real, imag} */,
  {32'h4590d058, 32'h00000000} /* (23, 0, 12) {real, imag} */,
  {32'h4561c134, 32'h00000000} /* (23, 0, 11) {real, imag} */,
  {32'h453ae1ea, 32'h00000000} /* (23, 0, 10) {real, imag} */,
  {32'h44b6b990, 32'h00000000} /* (23, 0, 9) {real, imag} */,
  {32'h449b45ac, 32'h00000000} /* (23, 0, 8) {real, imag} */,
  {32'hc4b60b70, 32'h00000000} /* (23, 0, 7) {real, imag} */,
  {32'hc53f61e4, 32'h00000000} /* (23, 0, 6) {real, imag} */,
  {32'hc59b34c0, 32'h00000000} /* (23, 0, 5) {real, imag} */,
  {32'hc5d441e6, 32'h00000000} /* (23, 0, 4) {real, imag} */,
  {32'hc6052a4e, 32'h00000000} /* (23, 0, 3) {real, imag} */,
  {32'hc614726b, 32'h00000000} /* (23, 0, 2) {real, imag} */,
  {32'hc61c06ae, 32'h00000000} /* (23, 0, 1) {real, imag} */,
  {32'hc620307e, 32'h00000000} /* (23, 0, 0) {real, imag} */,
  {32'hc641a02f, 32'h00000000} /* (22, 31, 31) {real, imag} */,
  {32'hc64ac5ae, 32'h00000000} /* (22, 31, 30) {real, imag} */,
  {32'hc64dce54, 32'h00000000} /* (22, 31, 29) {real, imag} */,
  {32'hc651b2eb, 32'h00000000} /* (22, 31, 28) {real, imag} */,
  {32'hc6559e7a, 32'h00000000} /* (22, 31, 27) {real, imag} */,
  {32'hc649032a, 32'h00000000} /* (22, 31, 26) {real, imag} */,
  {32'hc6400e6a, 32'h00000000} /* (22, 31, 25) {real, imag} */,
  {32'hc63e357a, 32'h00000000} /* (22, 31, 24) {real, imag} */,
  {32'hc61cf330, 32'h00000000} /* (22, 31, 23) {real, imag} */,
  {32'hc600f97b, 32'h00000000} /* (22, 31, 22) {real, imag} */,
  {32'hc5bec5ab, 32'h00000000} /* (22, 31, 21) {real, imag} */,
  {32'hc546d3a3, 32'h00000000} /* (22, 31, 20) {real, imag} */,
  {32'hc4917048, 32'h00000000} /* (22, 31, 19) {real, imag} */,
  {32'h4465d450, 32'h00000000} /* (22, 31, 18) {real, imag} */,
  {32'h4501e474, 32'h00000000} /* (22, 31, 17) {real, imag} */,
  {32'h458115da, 32'h00000000} /* (22, 31, 16) {real, imag} */,
  {32'h45b00af6, 32'h00000000} /* (22, 31, 15) {real, imag} */,
  {32'h45a82e77, 32'h00000000} /* (22, 31, 14) {real, imag} */,
  {32'h45b585e4, 32'h00000000} /* (22, 31, 13) {real, imag} */,
  {32'h45ac8aca, 32'h00000000} /* (22, 31, 12) {real, imag} */,
  {32'h455dbca2, 32'h00000000} /* (22, 31, 11) {real, imag} */,
  {32'h44f35d3c, 32'h00000000} /* (22, 31, 10) {real, imag} */,
  {32'hc410aa98, 32'h00000000} /* (22, 31, 9) {real, imag} */,
  {32'hc5230da2, 32'h00000000} /* (22, 31, 8) {real, imag} */,
  {32'hc56547a8, 32'h00000000} /* (22, 31, 7) {real, imag} */,
  {32'hc5a6d61c, 32'h00000000} /* (22, 31, 6) {real, imag} */,
  {32'hc5d6cbd1, 32'h00000000} /* (22, 31, 5) {real, imag} */,
  {32'hc607339b, 32'h00000000} /* (22, 31, 4) {real, imag} */,
  {32'hc6110e04, 32'h00000000} /* (22, 31, 3) {real, imag} */,
  {32'hc62496ff, 32'h00000000} /* (22, 31, 2) {real, imag} */,
  {32'hc635fb45, 32'h00000000} /* (22, 31, 1) {real, imag} */,
  {32'hc633bcf1, 32'h00000000} /* (22, 31, 0) {real, imag} */,
  {32'hc647eae2, 32'h00000000} /* (22, 30, 31) {real, imag} */,
  {32'hc64efedc, 32'h00000000} /* (22, 30, 30) {real, imag} */,
  {32'hc659117b, 32'h00000000} /* (22, 30, 29) {real, imag} */,
  {32'hc65d3e0f, 32'h00000000} /* (22, 30, 28) {real, imag} */,
  {32'hc64980c9, 32'h00000000} /* (22, 30, 27) {real, imag} */,
  {32'hc64f2d7a, 32'h00000000} /* (22, 30, 26) {real, imag} */,
  {32'hc6519107, 32'h00000000} /* (22, 30, 25) {real, imag} */,
  {32'hc64ff00e, 32'h00000000} /* (22, 30, 24) {real, imag} */,
  {32'hc62690fa, 32'h00000000} /* (22, 30, 23) {real, imag} */,
  {32'hc6053f90, 32'h00000000} /* (22, 30, 22) {real, imag} */,
  {32'hc5b136d0, 32'h00000000} /* (22, 30, 21) {real, imag} */,
  {32'hc41cfb90, 32'h00000000} /* (22, 30, 20) {real, imag} */,
  {32'h4419f980, 32'h00000000} /* (22, 30, 19) {real, imag} */,
  {32'h452b01b6, 32'h00000000} /* (22, 30, 18) {real, imag} */,
  {32'h457dcb6a, 32'h00000000} /* (22, 30, 17) {real, imag} */,
  {32'h45b0cc6f, 32'h00000000} /* (22, 30, 16) {real, imag} */,
  {32'h45c78fb8, 32'h00000000} /* (22, 30, 15) {real, imag} */,
  {32'h45ca2d84, 32'h00000000} /* (22, 30, 14) {real, imag} */,
  {32'h45d9d306, 32'h00000000} /* (22, 30, 13) {real, imag} */,
  {32'h45bbd67e, 32'h00000000} /* (22, 30, 12) {real, imag} */,
  {32'h452f2a30, 32'h00000000} /* (22, 30, 11) {real, imag} */,
  {32'hc2c4cd40, 32'h00000000} /* (22, 30, 10) {real, imag} */,
  {32'hc5150478, 32'h00000000} /* (22, 30, 9) {real, imag} */,
  {32'hc58f61cd, 32'h00000000} /* (22, 30, 8) {real, imag} */,
  {32'hc5bade58, 32'h00000000} /* (22, 30, 7) {real, imag} */,
  {32'hc5cf85af, 32'h00000000} /* (22, 30, 6) {real, imag} */,
  {32'hc60d4a78, 32'h00000000} /* (22, 30, 5) {real, imag} */,
  {32'hc615d549, 32'h00000000} /* (22, 30, 4) {real, imag} */,
  {32'hc621803b, 32'h00000000} /* (22, 30, 3) {real, imag} */,
  {32'hc63183f6, 32'h00000000} /* (22, 30, 2) {real, imag} */,
  {32'hc6406702, 32'h00000000} /* (22, 30, 1) {real, imag} */,
  {32'hc64120f0, 32'h00000000} /* (22, 30, 0) {real, imag} */,
  {32'hc6424066, 32'h00000000} /* (22, 29, 31) {real, imag} */,
  {32'hc6503afb, 32'h00000000} /* (22, 29, 30) {real, imag} */,
  {32'hc6578bd4, 32'h00000000} /* (22, 29, 29) {real, imag} */,
  {32'hc65e0498, 32'h00000000} /* (22, 29, 28) {real, imag} */,
  {32'hc65d5924, 32'h00000000} /* (22, 29, 27) {real, imag} */,
  {32'hc64e57f9, 32'h00000000} /* (22, 29, 26) {real, imag} */,
  {32'hc64e2146, 32'h00000000} /* (22, 29, 25) {real, imag} */,
  {32'hc63adf44, 32'h00000000} /* (22, 29, 24) {real, imag} */,
  {32'hc6264036, 32'h00000000} /* (22, 29, 23) {real, imag} */,
  {32'hc6000ebd, 32'h00000000} /* (22, 29, 22) {real, imag} */,
  {32'hc5ae0860, 32'h00000000} /* (22, 29, 21) {real, imag} */,
  {32'hc4433768, 32'h00000000} /* (22, 29, 20) {real, imag} */,
  {32'h456b0039, 32'h00000000} /* (22, 29, 19) {real, imag} */,
  {32'h4585f002, 32'h00000000} /* (22, 29, 18) {real, imag} */,
  {32'h45c7ca86, 32'h00000000} /* (22, 29, 17) {real, imag} */,
  {32'h45e30978, 32'h00000000} /* (22, 29, 16) {real, imag} */,
  {32'h45e307bc, 32'h00000000} /* (22, 29, 15) {real, imag} */,
  {32'h45e3936a, 32'h00000000} /* (22, 29, 14) {real, imag} */,
  {32'h45d0628f, 32'h00000000} /* (22, 29, 13) {real, imag} */,
  {32'h45b94063, 32'h00000000} /* (22, 29, 12) {real, imag} */,
  {32'h45389de0, 32'h00000000} /* (22, 29, 11) {real, imag} */,
  {32'hc44abe90, 32'h00000000} /* (22, 29, 10) {real, imag} */,
  {32'hc56422d8, 32'h00000000} /* (22, 29, 9) {real, imag} */,
  {32'hc5c4def1, 32'h00000000} /* (22, 29, 8) {real, imag} */,
  {32'hc5e2d33c, 32'h00000000} /* (22, 29, 7) {real, imag} */,
  {32'hc60682d3, 32'h00000000} /* (22, 29, 6) {real, imag} */,
  {32'hc61bd849, 32'h00000000} /* (22, 29, 5) {real, imag} */,
  {32'hc623f7ba, 32'h00000000} /* (22, 29, 4) {real, imag} */,
  {32'hc6260b3f, 32'h00000000} /* (22, 29, 3) {real, imag} */,
  {32'hc6429915, 32'h00000000} /* (22, 29, 2) {real, imag} */,
  {32'hc65570d9, 32'h00000000} /* (22, 29, 1) {real, imag} */,
  {32'hc644a08c, 32'h00000000} /* (22, 29, 0) {real, imag} */,
  {32'hc647e07a, 32'h00000000} /* (22, 28, 31) {real, imag} */,
  {32'hc6510f10, 32'h00000000} /* (22, 28, 30) {real, imag} */,
  {32'hc65fa412, 32'h00000000} /* (22, 28, 29) {real, imag} */,
  {32'hc65ca0ce, 32'h00000000} /* (22, 28, 28) {real, imag} */,
  {32'hc65c4353, 32'h00000000} /* (22, 28, 27) {real, imag} */,
  {32'hc65136f1, 32'h00000000} /* (22, 28, 26) {real, imag} */,
  {32'hc654cc2e, 32'h00000000} /* (22, 28, 25) {real, imag} */,
  {32'hc6404657, 32'h00000000} /* (22, 28, 24) {real, imag} */,
  {32'hc623abe3, 32'h00000000} /* (22, 28, 23) {real, imag} */,
  {32'hc60ad23a, 32'h00000000} /* (22, 28, 22) {real, imag} */,
  {32'hc58feaa0, 32'h00000000} /* (22, 28, 21) {real, imag} */,
  {32'h42c896c0, 32'h00000000} /* (22, 28, 20) {real, imag} */,
  {32'h45819fbb, 32'h00000000} /* (22, 28, 19) {real, imag} */,
  {32'h45c5e770, 32'h00000000} /* (22, 28, 18) {real, imag} */,
  {32'h45c8994b, 32'h00000000} /* (22, 28, 17) {real, imag} */,
  {32'h45f46be3, 32'h00000000} /* (22, 28, 16) {real, imag} */,
  {32'h460b327c, 32'h00000000} /* (22, 28, 15) {real, imag} */,
  {32'h45e8d780, 32'h00000000} /* (22, 28, 14) {real, imag} */,
  {32'h45c604af, 32'h00000000} /* (22, 28, 13) {real, imag} */,
  {32'h45a8c00b, 32'h00000000} /* (22, 28, 12) {real, imag} */,
  {32'h45288b3c, 32'h00000000} /* (22, 28, 11) {real, imag} */,
  {32'hc4935078, 32'h00000000} /* (22, 28, 10) {real, imag} */,
  {32'hc59350fc, 32'h00000000} /* (22, 28, 9) {real, imag} */,
  {32'hc5e0016a, 32'h00000000} /* (22, 28, 8) {real, imag} */,
  {32'hc603cacd, 32'h00000000} /* (22, 28, 7) {real, imag} */,
  {32'hc61e5794, 32'h00000000} /* (22, 28, 6) {real, imag} */,
  {32'hc62ee53b, 32'h00000000} /* (22, 28, 5) {real, imag} */,
  {32'hc633834e, 32'h00000000} /* (22, 28, 4) {real, imag} */,
  {32'hc63b9ce8, 32'h00000000} /* (22, 28, 3) {real, imag} */,
  {32'hc64b0a8e, 32'h00000000} /* (22, 28, 2) {real, imag} */,
  {32'hc64852f0, 32'h00000000} /* (22, 28, 1) {real, imag} */,
  {32'hc641483e, 32'h00000000} /* (22, 28, 0) {real, imag} */,
  {32'hc63ea105, 32'h00000000} /* (22, 27, 31) {real, imag} */,
  {32'hc64999af, 32'h00000000} /* (22, 27, 30) {real, imag} */,
  {32'hc647db11, 32'h00000000} /* (22, 27, 29) {real, imag} */,
  {32'hc6575fa8, 32'h00000000} /* (22, 27, 28) {real, imag} */,
  {32'hc664cb86, 32'h00000000} /* (22, 27, 27) {real, imag} */,
  {32'hc64fc525, 32'h00000000} /* (22, 27, 26) {real, imag} */,
  {32'hc64589f8, 32'h00000000} /* (22, 27, 25) {real, imag} */,
  {32'hc636fd43, 32'h00000000} /* (22, 27, 24) {real, imag} */,
  {32'hc612a222, 32'h00000000} /* (22, 27, 23) {real, imag} */,
  {32'hc5dcfa58, 32'h00000000} /* (22, 27, 22) {real, imag} */,
  {32'hc5669ce0, 32'h00000000} /* (22, 27, 21) {real, imag} */,
  {32'h4438e890, 32'h00000000} /* (22, 27, 20) {real, imag} */,
  {32'h454f894c, 32'h00000000} /* (22, 27, 19) {real, imag} */,
  {32'h45b21d62, 32'h00000000} /* (22, 27, 18) {real, imag} */,
  {32'h45eb1bc2, 32'h00000000} /* (22, 27, 17) {real, imag} */,
  {32'h45f15513, 32'h00000000} /* (22, 27, 16) {real, imag} */,
  {32'h45fe5336, 32'h00000000} /* (22, 27, 15) {real, imag} */,
  {32'h45ec1c6e, 32'h00000000} /* (22, 27, 14) {real, imag} */,
  {32'h45dded56, 32'h00000000} /* (22, 27, 13) {real, imag} */,
  {32'h459bfc49, 32'h00000000} /* (22, 27, 12) {real, imag} */,
  {32'h4506aab6, 32'h00000000} /* (22, 27, 11) {real, imag} */,
  {32'hc4cd3538, 32'h00000000} /* (22, 27, 10) {real, imag} */,
  {32'hc5bcc6cc, 32'h00000000} /* (22, 27, 9) {real, imag} */,
  {32'hc606e4a1, 32'h00000000} /* (22, 27, 8) {real, imag} */,
  {32'hc61221fe, 32'h00000000} /* (22, 27, 7) {real, imag} */,
  {32'hc61aa0f2, 32'h00000000} /* (22, 27, 6) {real, imag} */,
  {32'hc640717c, 32'h00000000} /* (22, 27, 5) {real, imag} */,
  {32'hc646eb56, 32'h00000000} /* (22, 27, 4) {real, imag} */,
  {32'hc6466a00, 32'h00000000} /* (22, 27, 3) {real, imag} */,
  {32'hc64046c3, 32'h00000000} /* (22, 27, 2) {real, imag} */,
  {32'hc6494c31, 32'h00000000} /* (22, 27, 1) {real, imag} */,
  {32'hc6483508, 32'h00000000} /* (22, 27, 0) {real, imag} */,
  {32'hc6344aa6, 32'h00000000} /* (22, 26, 31) {real, imag} */,
  {32'hc63ac9d2, 32'h00000000} /* (22, 26, 30) {real, imag} */,
  {32'hc6452fce, 32'h00000000} /* (22, 26, 29) {real, imag} */,
  {32'hc64e2f9c, 32'h00000000} /* (22, 26, 28) {real, imag} */,
  {32'hc64a8b41, 32'h00000000} /* (22, 26, 27) {real, imag} */,
  {32'hc645eb70, 32'h00000000} /* (22, 26, 26) {real, imag} */,
  {32'hc63d974c, 32'h00000000} /* (22, 26, 25) {real, imag} */,
  {32'hc631967f, 32'h00000000} /* (22, 26, 24) {real, imag} */,
  {32'hc613affd, 32'h00000000} /* (22, 26, 23) {real, imag} */,
  {32'hc5eaf848, 32'h00000000} /* (22, 26, 22) {real, imag} */,
  {32'hc56496a4, 32'h00000000} /* (22, 26, 21) {real, imag} */,
  {32'h439b1010, 32'h00000000} /* (22, 26, 20) {real, imag} */,
  {32'h455f5aa4, 32'h00000000} /* (22, 26, 19) {real, imag} */,
  {32'h45aac134, 32'h00000000} /* (22, 26, 18) {real, imag} */,
  {32'h45e416d0, 32'h00000000} /* (22, 26, 17) {real, imag} */,
  {32'h45ea19a0, 32'h00000000} /* (22, 26, 16) {real, imag} */,
  {32'h45d7c7c8, 32'h00000000} /* (22, 26, 15) {real, imag} */,
  {32'h45e81b20, 32'h00000000} /* (22, 26, 14) {real, imag} */,
  {32'h45daa82d, 32'h00000000} /* (22, 26, 13) {real, imag} */,
  {32'h45978ae1, 32'h00000000} /* (22, 26, 12) {real, imag} */,
  {32'h450fcd1c, 32'h00000000} /* (22, 26, 11) {real, imag} */,
  {32'hc5097408, 32'h00000000} /* (22, 26, 10) {real, imag} */,
  {32'hc5d8ec91, 32'h00000000} /* (22, 26, 9) {real, imag} */,
  {32'hc5eb6c9e, 32'h00000000} /* (22, 26, 8) {real, imag} */,
  {32'hc608360f, 32'h00000000} /* (22, 26, 7) {real, imag} */,
  {32'hc621edc4, 32'h00000000} /* (22, 26, 6) {real, imag} */,
  {32'hc624935c, 32'h00000000} /* (22, 26, 5) {real, imag} */,
  {32'hc63b9072, 32'h00000000} /* (22, 26, 4) {real, imag} */,
  {32'hc641a179, 32'h00000000} /* (22, 26, 3) {real, imag} */,
  {32'hc64029da, 32'h00000000} /* (22, 26, 2) {real, imag} */,
  {32'hc64660e0, 32'h00000000} /* (22, 26, 1) {real, imag} */,
  {32'hc633fe0a, 32'h00000000} /* (22, 26, 0) {real, imag} */,
  {32'hc6285bf9, 32'h00000000} /* (22, 25, 31) {real, imag} */,
  {32'hc62eff9b, 32'h00000000} /* (22, 25, 30) {real, imag} */,
  {32'hc63b3ff4, 32'h00000000} /* (22, 25, 29) {real, imag} */,
  {32'hc6360a58, 32'h00000000} /* (22, 25, 28) {real, imag} */,
  {32'hc6328899, 32'h00000000} /* (22, 25, 27) {real, imag} */,
  {32'hc638bedb, 32'h00000000} /* (22, 25, 26) {real, imag} */,
  {32'hc6217871, 32'h00000000} /* (22, 25, 25) {real, imag} */,
  {32'hc6294e5e, 32'h00000000} /* (22, 25, 24) {real, imag} */,
  {32'hc6155551, 32'h00000000} /* (22, 25, 23) {real, imag} */,
  {32'hc5d6d539, 32'h00000000} /* (22, 25, 22) {real, imag} */,
  {32'hc555f0c4, 32'h00000000} /* (22, 25, 21) {real, imag} */,
  {32'h443f05d8, 32'h00000000} /* (22, 25, 20) {real, imag} */,
  {32'h45609fc1, 32'h00000000} /* (22, 25, 19) {real, imag} */,
  {32'h45b51280, 32'h00000000} /* (22, 25, 18) {real, imag} */,
  {32'h45dee356, 32'h00000000} /* (22, 25, 17) {real, imag} */,
  {32'h45f44b40, 32'h00000000} /* (22, 25, 16) {real, imag} */,
  {32'h45e247ee, 32'h00000000} /* (22, 25, 15) {real, imag} */,
  {32'h45de2832, 32'h00000000} /* (22, 25, 14) {real, imag} */,
  {32'h45b3a113, 32'h00000000} /* (22, 25, 13) {real, imag} */,
  {32'h45802037, 32'h00000000} /* (22, 25, 12) {real, imag} */,
  {32'h44b90da8, 32'h00000000} /* (22, 25, 11) {real, imag} */,
  {32'hc53bd2d4, 32'h00000000} /* (22, 25, 10) {real, imag} */,
  {32'hc5b4b8be, 32'h00000000} /* (22, 25, 9) {real, imag} */,
  {32'hc5f351c0, 32'h00000000} /* (22, 25, 8) {real, imag} */,
  {32'hc6005421, 32'h00000000} /* (22, 25, 7) {real, imag} */,
  {32'hc61d11a0, 32'h00000000} /* (22, 25, 6) {real, imag} */,
  {32'hc62385da, 32'h00000000} /* (22, 25, 5) {real, imag} */,
  {32'hc6291828, 32'h00000000} /* (22, 25, 4) {real, imag} */,
  {32'hc62b4588, 32'h00000000} /* (22, 25, 3) {real, imag} */,
  {32'hc63181ce, 32'h00000000} /* (22, 25, 2) {real, imag} */,
  {32'hc6353985, 32'h00000000} /* (22, 25, 1) {real, imag} */,
  {32'hc622ac90, 32'h00000000} /* (22, 25, 0) {real, imag} */,
  {32'hc60fecb2, 32'h00000000} /* (22, 24, 31) {real, imag} */,
  {32'hc6281b4f, 32'h00000000} /* (22, 24, 30) {real, imag} */,
  {32'hc6274924, 32'h00000000} /* (22, 24, 29) {real, imag} */,
  {32'hc6241178, 32'h00000000} /* (22, 24, 28) {real, imag} */,
  {32'hc62c45d6, 32'h00000000} /* (22, 24, 27) {real, imag} */,
  {32'hc6100f2a, 32'h00000000} /* (22, 24, 26) {real, imag} */,
  {32'hc618a5d0, 32'h00000000} /* (22, 24, 25) {real, imag} */,
  {32'hc603a62f, 32'h00000000} /* (22, 24, 24) {real, imag} */,
  {32'hc5dcd10a, 32'h00000000} /* (22, 24, 23) {real, imag} */,
  {32'hc5c6f250, 32'h00000000} /* (22, 24, 22) {real, imag} */,
  {32'hc535eeee, 32'h00000000} /* (22, 24, 21) {real, imag} */,
  {32'h4426c6f8, 32'h00000000} /* (22, 24, 20) {real, imag} */,
  {32'h45818fee, 32'h00000000} /* (22, 24, 19) {real, imag} */,
  {32'h45b79f1c, 32'h00000000} /* (22, 24, 18) {real, imag} */,
  {32'h45d770ec, 32'h00000000} /* (22, 24, 17) {real, imag} */,
  {32'h45ee6ea4, 32'h00000000} /* (22, 24, 16) {real, imag} */,
  {32'h45f8f7cf, 32'h00000000} /* (22, 24, 15) {real, imag} */,
  {32'h45c5c286, 32'h00000000} /* (22, 24, 14) {real, imag} */,
  {32'h45a28fc6, 32'h00000000} /* (22, 24, 13) {real, imag} */,
  {32'h45564d46, 32'h00000000} /* (22, 24, 12) {real, imag} */,
  {32'h447f0438, 32'h00000000} /* (22, 24, 11) {real, imag} */,
  {32'hc52e0ea4, 32'h00000000} /* (22, 24, 10) {real, imag} */,
  {32'hc588d341, 32'h00000000} /* (22, 24, 9) {real, imag} */,
  {32'hc5f421e2, 32'h00000000} /* (22, 24, 8) {real, imag} */,
  {32'hc600069e, 32'h00000000} /* (22, 24, 7) {real, imag} */,
  {32'hc6099478, 32'h00000000} /* (22, 24, 6) {real, imag} */,
  {32'hc60f84a4, 32'h00000000} /* (22, 24, 5) {real, imag} */,
  {32'hc611270e, 32'h00000000} /* (22, 24, 4) {real, imag} */,
  {32'hc619d021, 32'h00000000} /* (22, 24, 3) {real, imag} */,
  {32'hc618c7b6, 32'h00000000} /* (22, 24, 2) {real, imag} */,
  {32'hc60a41d9, 32'h00000000} /* (22, 24, 1) {real, imag} */,
  {32'hc60c2ed4, 32'h00000000} /* (22, 24, 0) {real, imag} */,
  {32'hc5e5836a, 32'h00000000} /* (22, 23, 31) {real, imag} */,
  {32'hc6034a46, 32'h00000000} /* (22, 23, 30) {real, imag} */,
  {32'hc60c1e4d, 32'h00000000} /* (22, 23, 29) {real, imag} */,
  {32'hc608e8cd, 32'h00000000} /* (22, 23, 28) {real, imag} */,
  {32'hc604d946, 32'h00000000} /* (22, 23, 27) {real, imag} */,
  {32'hc5f35d7d, 32'h00000000} /* (22, 23, 26) {real, imag} */,
  {32'hc5e8df92, 32'h00000000} /* (22, 23, 25) {real, imag} */,
  {32'hc5c8c321, 32'h00000000} /* (22, 23, 24) {real, imag} */,
  {32'hc5dc7a6d, 32'h00000000} /* (22, 23, 23) {real, imag} */,
  {32'hc5a3f76c, 32'h00000000} /* (22, 23, 22) {real, imag} */,
  {32'hc4d7dad4, 32'h00000000} /* (22, 23, 21) {real, imag} */,
  {32'h445ab9d4, 32'h00000000} /* (22, 23, 20) {real, imag} */,
  {32'h45594c6d, 32'h00000000} /* (22, 23, 19) {real, imag} */,
  {32'h45876ab0, 32'h00000000} /* (22, 23, 18) {real, imag} */,
  {32'h459d1f2e, 32'h00000000} /* (22, 23, 17) {real, imag} */,
  {32'h45aff597, 32'h00000000} /* (22, 23, 16) {real, imag} */,
  {32'h45a9ba9a, 32'h00000000} /* (22, 23, 15) {real, imag} */,
  {32'h45a7ade8, 32'h00000000} /* (22, 23, 14) {real, imag} */,
  {32'h45877c26, 32'h00000000} /* (22, 23, 13) {real, imag} */,
  {32'h45466f55, 32'h00000000} /* (22, 23, 12) {real, imag} */,
  {32'h443d0b44, 32'h00000000} /* (22, 23, 11) {real, imag} */,
  {32'hc4afae74, 32'h00000000} /* (22, 23, 10) {real, imag} */,
  {32'hc54f7bfd, 32'h00000000} /* (22, 23, 9) {real, imag} */,
  {32'hc5b2919b, 32'h00000000} /* (22, 23, 8) {real, imag} */,
  {32'hc5efbbfb, 32'h00000000} /* (22, 23, 7) {real, imag} */,
  {32'hc5e63cdc, 32'h00000000} /* (22, 23, 6) {real, imag} */,
  {32'hc5fcad13, 32'h00000000} /* (22, 23, 5) {real, imag} */,
  {32'hc602469a, 32'h00000000} /* (22, 23, 4) {real, imag} */,
  {32'hc60e12db, 32'h00000000} /* (22, 23, 3) {real, imag} */,
  {32'hc60225fd, 32'h00000000} /* (22, 23, 2) {real, imag} */,
  {32'hc5f34d32, 32'h00000000} /* (22, 23, 1) {real, imag} */,
  {32'hc5eb4f3b, 32'h00000000} /* (22, 23, 0) {real, imag} */,
  {32'hc5a0c780, 32'h00000000} /* (22, 22, 31) {real, imag} */,
  {32'hc5c6d228, 32'h00000000} /* (22, 22, 30) {real, imag} */,
  {32'hc5c035b4, 32'h00000000} /* (22, 22, 29) {real, imag} */,
  {32'hc5c9bd97, 32'h00000000} /* (22, 22, 28) {real, imag} */,
  {32'hc5b7b4ef, 32'h00000000} /* (22, 22, 27) {real, imag} */,
  {32'hc594f246, 32'h00000000} /* (22, 22, 26) {real, imag} */,
  {32'hc5957f21, 32'h00000000} /* (22, 22, 25) {real, imag} */,
  {32'hc58a6c24, 32'h00000000} /* (22, 22, 24) {real, imag} */,
  {32'hc59217e1, 32'h00000000} /* (22, 22, 23) {real, imag} */,
  {32'hc5610f4a, 32'h00000000} /* (22, 22, 22) {real, imag} */,
  {32'hc4d6e19a, 32'h00000000} /* (22, 22, 21) {real, imag} */,
  {32'h44990574, 32'h00000000} /* (22, 22, 20) {real, imag} */,
  {32'h44ededec, 32'h00000000} /* (22, 22, 19) {real, imag} */,
  {32'h4542cc50, 32'h00000000} /* (22, 22, 18) {real, imag} */,
  {32'h4551ee2d, 32'h00000000} /* (22, 22, 17) {real, imag} */,
  {32'h455f6ec3, 32'h00000000} /* (22, 22, 16) {real, imag} */,
  {32'h45605da8, 32'h00000000} /* (22, 22, 15) {real, imag} */,
  {32'h454fd840, 32'h00000000} /* (22, 22, 14) {real, imag} */,
  {32'h45464e50, 32'h00000000} /* (22, 22, 13) {real, imag} */,
  {32'h45209bfe, 32'h00000000} /* (22, 22, 12) {real, imag} */,
  {32'h44ae55fc, 32'h00000000} /* (22, 22, 11) {real, imag} */,
  {32'hc488a769, 32'h00000000} /* (22, 22, 10) {real, imag} */,
  {32'hc5529d8c, 32'h00000000} /* (22, 22, 9) {real, imag} */,
  {32'hc560b162, 32'h00000000} /* (22, 22, 8) {real, imag} */,
  {32'hc5977e57, 32'h00000000} /* (22, 22, 7) {real, imag} */,
  {32'hc5b7d383, 32'h00000000} /* (22, 22, 6) {real, imag} */,
  {32'hc5ac320e, 32'h00000000} /* (22, 22, 5) {real, imag} */,
  {32'hc5aa9aa6, 32'h00000000} /* (22, 22, 4) {real, imag} */,
  {32'hc5b45ed7, 32'h00000000} /* (22, 22, 3) {real, imag} */,
  {32'hc5a6c57c, 32'h00000000} /* (22, 22, 2) {real, imag} */,
  {32'hc5bf5380, 32'h00000000} /* (22, 22, 1) {real, imag} */,
  {32'hc5a86648, 32'h00000000} /* (22, 22, 0) {real, imag} */,
  {32'hc50e4d53, 32'h00000000} /* (22, 21, 31) {real, imag} */,
  {32'hc52bcbee, 32'h00000000} /* (22, 21, 30) {real, imag} */,
  {32'hc5295e76, 32'h00000000} /* (22, 21, 29) {real, imag} */,
  {32'hc524641d, 32'h00000000} /* (22, 21, 28) {real, imag} */,
  {32'hc4fc512d, 32'h00000000} /* (22, 21, 27) {real, imag} */,
  {32'hc4dfd4d8, 32'h00000000} /* (22, 21, 26) {real, imag} */,
  {32'hc4e9786f, 32'h00000000} /* (22, 21, 25) {real, imag} */,
  {32'hc4b5038b, 32'h00000000} /* (22, 21, 24) {real, imag} */,
  {32'hc4e56136, 32'h00000000} /* (22, 21, 23) {real, imag} */,
  {32'hc489ece7, 32'h00000000} /* (22, 21, 22) {real, imag} */,
  {32'hc4cf46c5, 32'h00000000} /* (22, 21, 21) {real, imag} */,
  {32'h432c27a0, 32'h00000000} /* (22, 21, 20) {real, imag} */,
  {32'h44812113, 32'h00000000} /* (22, 21, 19) {real, imag} */,
  {32'h4100a880, 32'h00000000} /* (22, 21, 18) {real, imag} */,
  {32'h445e28c8, 32'h00000000} /* (22, 21, 17) {real, imag} */,
  {32'h443b487c, 32'h00000000} /* (22, 21, 16) {real, imag} */,
  {32'h448a95b8, 32'h00000000} /* (22, 21, 15) {real, imag} */,
  {32'h446ad472, 32'h00000000} /* (22, 21, 14) {real, imag} */,
  {32'h44f1873d, 32'h00000000} /* (22, 21, 13) {real, imag} */,
  {32'h450dc2dd, 32'h00000000} /* (22, 21, 12) {real, imag} */,
  {32'h4424ea3e, 32'h00000000} /* (22, 21, 11) {real, imag} */,
  {32'hc4c92446, 32'h00000000} /* (22, 21, 10) {real, imag} */,
  {32'hc48e31c3, 32'h00000000} /* (22, 21, 9) {real, imag} */,
  {32'hc4d2d035, 32'h00000000} /* (22, 21, 8) {real, imag} */,
  {32'hc52482c1, 32'h00000000} /* (22, 21, 7) {real, imag} */,
  {32'hc514d332, 32'h00000000} /* (22, 21, 6) {real, imag} */,
  {32'hc518370e, 32'h00000000} /* (22, 21, 5) {real, imag} */,
  {32'hc518a680, 32'h00000000} /* (22, 21, 4) {real, imag} */,
  {32'hc4f99cbd, 32'h00000000} /* (22, 21, 3) {real, imag} */,
  {32'hc51cc1f0, 32'h00000000} /* (22, 21, 2) {real, imag} */,
  {32'hc53aad95, 32'h00000000} /* (22, 21, 1) {real, imag} */,
  {32'hc50a6a1d, 32'h00000000} /* (22, 21, 0) {real, imag} */,
  {32'h44d4a722, 32'h00000000} /* (22, 20, 31) {real, imag} */,
  {32'h452cdcea, 32'h00000000} /* (22, 20, 30) {real, imag} */,
  {32'h451f2344, 32'h00000000} /* (22, 20, 29) {real, imag} */,
  {32'h450be466, 32'h00000000} /* (22, 20, 28) {real, imag} */,
  {32'h4528ef64, 32'h00000000} /* (22, 20, 27) {real, imag} */,
  {32'h45140cfd, 32'h00000000} /* (22, 20, 26) {real, imag} */,
  {32'h4511f1e5, 32'h00000000} /* (22, 20, 25) {real, imag} */,
  {32'h45363196, 32'h00000000} /* (22, 20, 24) {real, imag} */,
  {32'h44b97cf4, 32'h00000000} /* (22, 20, 23) {real, imag} */,
  {32'h441ce226, 32'h00000000} /* (22, 20, 22) {real, imag} */,
  {32'hc2e74420, 32'h00000000} /* (22, 20, 21) {real, imag} */,
  {32'hc4ba54d4, 32'h00000000} /* (22, 20, 20) {real, imag} */,
  {32'hc5009b2a, 32'h00000000} /* (22, 20, 19) {real, imag} */,
  {32'hc53df774, 32'h00000000} /* (22, 20, 18) {real, imag} */,
  {32'hc5556c24, 32'h00000000} /* (22, 20, 17) {real, imag} */,
  {32'hc537ecd9, 32'h00000000} /* (22, 20, 16) {real, imag} */,
  {32'hc4ee59fc, 32'h00000000} /* (22, 20, 15) {real, imag} */,
  {32'hc4c0d281, 32'h00000000} /* (22, 20, 14) {real, imag} */,
  {32'hc5097b1e, 32'h00000000} /* (22, 20, 13) {real, imag} */,
  {32'hc4a67389, 32'h00000000} /* (22, 20, 12) {real, imag} */,
  {32'hc479db08, 32'h00000000} /* (22, 20, 11) {real, imag} */,
  {32'hc3548b30, 32'h00000000} /* (22, 20, 10) {real, imag} */,
  {32'h4493977e, 32'h00000000} /* (22, 20, 9) {real, imag} */,
  {32'h4428c850, 32'h00000000} /* (22, 20, 8) {real, imag} */,
  {32'h448a6248, 32'h00000000} /* (22, 20, 7) {real, imag} */,
  {32'h44d7881d, 32'h00000000} /* (22, 20, 6) {real, imag} */,
  {32'h4508d071, 32'h00000000} /* (22, 20, 5) {real, imag} */,
  {32'h4509f689, 32'h00000000} /* (22, 20, 4) {real, imag} */,
  {32'h44eb2c25, 32'h00000000} /* (22, 20, 3) {real, imag} */,
  {32'h44cbcfa4, 32'h00000000} /* (22, 20, 2) {real, imag} */,
  {32'h4483171c, 32'h00000000} /* (22, 20, 1) {real, imag} */,
  {32'h446723dc, 32'h00000000} /* (22, 20, 0) {real, imag} */,
  {32'h45848c32, 32'h00000000} /* (22, 19, 31) {real, imag} */,
  {32'h457bc2e0, 32'h00000000} /* (22, 19, 30) {real, imag} */,
  {32'h4589e3a6, 32'h00000000} /* (22, 19, 29) {real, imag} */,
  {32'h45940b2a, 32'h00000000} /* (22, 19, 28) {real, imag} */,
  {32'h45b7648a, 32'h00000000} /* (22, 19, 27) {real, imag} */,
  {32'h458eac5e, 32'h00000000} /* (22, 19, 26) {real, imag} */,
  {32'h4587c852, 32'h00000000} /* (22, 19, 25) {real, imag} */,
  {32'h45860ee2, 32'h00000000} /* (22, 19, 24) {real, imag} */,
  {32'h4569aced, 32'h00000000} /* (22, 19, 23) {real, imag} */,
  {32'h45299c3c, 32'h00000000} /* (22, 19, 22) {real, imag} */,
  {32'h434a6400, 32'h00000000} /* (22, 19, 21) {real, imag} */,
  {32'hc4f8558a, 32'h00000000} /* (22, 19, 20) {real, imag} */,
  {32'hc545ce76, 32'h00000000} /* (22, 19, 19) {real, imag} */,
  {32'hc586a37a, 32'h00000000} /* (22, 19, 18) {real, imag} */,
  {32'hc595ce34, 32'h00000000} /* (22, 19, 17) {real, imag} */,
  {32'hc5aa72c0, 32'h00000000} /* (22, 19, 16) {real, imag} */,
  {32'hc59633d4, 32'h00000000} /* (22, 19, 15) {real, imag} */,
  {32'hc58e5f6c, 32'h00000000} /* (22, 19, 14) {real, imag} */,
  {32'hc59c8704, 32'h00000000} /* (22, 19, 13) {real, imag} */,
  {32'hc5930db2, 32'h00000000} /* (22, 19, 12) {real, imag} */,
  {32'hc504d8d0, 32'h00000000} /* (22, 19, 11) {real, imag} */,
  {32'h42da7980, 32'h00000000} /* (22, 19, 10) {real, imag} */,
  {32'h44c762ef, 32'h00000000} /* (22, 19, 9) {real, imag} */,
  {32'h450e1c74, 32'h00000000} /* (22, 19, 8) {real, imag} */,
  {32'h4568c8d9, 32'h00000000} /* (22, 19, 7) {real, imag} */,
  {32'h458def64, 32'h00000000} /* (22, 19, 6) {real, imag} */,
  {32'h4596bb7b, 32'h00000000} /* (22, 19, 5) {real, imag} */,
  {32'h45a3d6f8, 32'h00000000} /* (22, 19, 4) {real, imag} */,
  {32'h45a102a7, 32'h00000000} /* (22, 19, 3) {real, imag} */,
  {32'h458810e8, 32'h00000000} /* (22, 19, 2) {real, imag} */,
  {32'h456cf394, 32'h00000000} /* (22, 19, 1) {real, imag} */,
  {32'h45764420, 32'h00000000} /* (22, 19, 0) {real, imag} */,
  {32'h45caf82b, 32'h00000000} /* (22, 18, 31) {real, imag} */,
  {32'h45d9df3a, 32'h00000000} /* (22, 18, 30) {real, imag} */,
  {32'h45c7a1d0, 32'h00000000} /* (22, 18, 29) {real, imag} */,
  {32'h45dccd8a, 32'h00000000} /* (22, 18, 28) {real, imag} */,
  {32'h45cd6b4c, 32'h00000000} /* (22, 18, 27) {real, imag} */,
  {32'h45cadfb8, 32'h00000000} /* (22, 18, 26) {real, imag} */,
  {32'h45c2702c, 32'h00000000} /* (22, 18, 25) {real, imag} */,
  {32'h45abb4fe, 32'h00000000} /* (22, 18, 24) {real, imag} */,
  {32'h45834584, 32'h00000000} /* (22, 18, 23) {real, imag} */,
  {32'h4520c544, 32'h00000000} /* (22, 18, 22) {real, imag} */,
  {32'h43e32780, 32'h00000000} /* (22, 18, 21) {real, imag} */,
  {32'hc504ad20, 32'h00000000} /* (22, 18, 20) {real, imag} */,
  {32'hc581dde8, 32'h00000000} /* (22, 18, 19) {real, imag} */,
  {32'hc5c19a8e, 32'h00000000} /* (22, 18, 18) {real, imag} */,
  {32'hc5beb3ba, 32'h00000000} /* (22, 18, 17) {real, imag} */,
  {32'hc5db44b4, 32'h00000000} /* (22, 18, 16) {real, imag} */,
  {32'hc5dce405, 32'h00000000} /* (22, 18, 15) {real, imag} */,
  {32'hc5cd93d8, 32'h00000000} /* (22, 18, 14) {real, imag} */,
  {32'hc5b40884, 32'h00000000} /* (22, 18, 13) {real, imag} */,
  {32'hc59b946c, 32'h00000000} /* (22, 18, 12) {real, imag} */,
  {32'hc562523b, 32'h00000000} /* (22, 18, 11) {real, imag} */,
  {32'hc45f0fb4, 32'h00000000} /* (22, 18, 10) {real, imag} */,
  {32'h452929fc, 32'h00000000} /* (22, 18, 9) {real, imag} */,
  {32'h45939af4, 32'h00000000} /* (22, 18, 8) {real, imag} */,
  {32'h45bcce22, 32'h00000000} /* (22, 18, 7) {real, imag} */,
  {32'h45c2cdf4, 32'h00000000} /* (22, 18, 6) {real, imag} */,
  {32'h45baead6, 32'h00000000} /* (22, 18, 5) {real, imag} */,
  {32'h45c4cf74, 32'h00000000} /* (22, 18, 4) {real, imag} */,
  {32'h45c00f60, 32'h00000000} /* (22, 18, 3) {real, imag} */,
  {32'h45d703bc, 32'h00000000} /* (22, 18, 2) {real, imag} */,
  {32'h45d92856, 32'h00000000} /* (22, 18, 1) {real, imag} */,
  {32'h45bb6e42, 32'h00000000} /* (22, 18, 0) {real, imag} */,
  {32'h45f63d08, 32'h00000000} /* (22, 17, 31) {real, imag} */,
  {32'h45f3f7e2, 32'h00000000} /* (22, 17, 30) {real, imag} */,
  {32'h46008d0e, 32'h00000000} /* (22, 17, 29) {real, imag} */,
  {32'h45fa26cd, 32'h00000000} /* (22, 17, 28) {real, imag} */,
  {32'h45d8d171, 32'h00000000} /* (22, 17, 27) {real, imag} */,
  {32'h45d9c976, 32'h00000000} /* (22, 17, 26) {real, imag} */,
  {32'h45ef8b86, 32'h00000000} /* (22, 17, 25) {real, imag} */,
  {32'h45e658f0, 32'h00000000} /* (22, 17, 24) {real, imag} */,
  {32'h45c32a19, 32'h00000000} /* (22, 17, 23) {real, imag} */,
  {32'h45538624, 32'h00000000} /* (22, 17, 22) {real, imag} */,
  {32'h433cc960, 32'h00000000} /* (22, 17, 21) {real, imag} */,
  {32'hc5103e06, 32'h00000000} /* (22, 17, 20) {real, imag} */,
  {32'hc5b96208, 32'h00000000} /* (22, 17, 19) {real, imag} */,
  {32'hc5ef6a9d, 32'h00000000} /* (22, 17, 18) {real, imag} */,
  {32'hc5dca374, 32'h00000000} /* (22, 17, 17) {real, imag} */,
  {32'hc5e30422, 32'h00000000} /* (22, 17, 16) {real, imag} */,
  {32'hc5e6c220, 32'h00000000} /* (22, 17, 15) {real, imag} */,
  {32'hc5e07512, 32'h00000000} /* (22, 17, 14) {real, imag} */,
  {32'hc5cc413a, 32'h00000000} /* (22, 17, 13) {real, imag} */,
  {32'hc5ce2969, 32'h00000000} /* (22, 17, 12) {real, imag} */,
  {32'hc54dcba2, 32'h00000000} /* (22, 17, 11) {real, imag} */,
  {32'hc259f600, 32'h00000000} /* (22, 17, 10) {real, imag} */,
  {32'h456e6f7b, 32'h00000000} /* (22, 17, 9) {real, imag} */,
  {32'h45b8f4c0, 32'h00000000} /* (22, 17, 8) {real, imag} */,
  {32'h45d100d1, 32'h00000000} /* (22, 17, 7) {real, imag} */,
  {32'h45e0811a, 32'h00000000} /* (22, 17, 6) {real, imag} */,
  {32'h45ec4d05, 32'h00000000} /* (22, 17, 5) {real, imag} */,
  {32'h46038f0a, 32'h00000000} /* (22, 17, 4) {real, imag} */,
  {32'h45ecba0e, 32'h00000000} /* (22, 17, 3) {real, imag} */,
  {32'h46051f9e, 32'h00000000} /* (22, 17, 2) {real, imag} */,
  {32'h46032537, 32'h00000000} /* (22, 17, 1) {real, imag} */,
  {32'h45f68aac, 32'h00000000} /* (22, 17, 0) {real, imag} */,
  {32'h46051bf8, 32'h00000000} /* (22, 16, 31) {real, imag} */,
  {32'h460b9e21, 32'h00000000} /* (22, 16, 30) {real, imag} */,
  {32'h460532ce, 32'h00000000} /* (22, 16, 29) {real, imag} */,
  {32'h45fc5512, 32'h00000000} /* (22, 16, 28) {real, imag} */,
  {32'h45f44cfa, 32'h00000000} /* (22, 16, 27) {real, imag} */,
  {32'h45fef1d5, 32'h00000000} /* (22, 16, 26) {real, imag} */,
  {32'h4605e82a, 32'h00000000} /* (22, 16, 25) {real, imag} */,
  {32'h45e4e1cd, 32'h00000000} /* (22, 16, 24) {real, imag} */,
  {32'h45d3b37e, 32'h00000000} /* (22, 16, 23) {real, imag} */,
  {32'h458a892a, 32'h00000000} /* (22, 16, 22) {real, imag} */,
  {32'hc31dc980, 32'h00000000} /* (22, 16, 21) {real, imag} */,
  {32'hc560492a, 32'h00000000} /* (22, 16, 20) {real, imag} */,
  {32'hc5ba1ac3, 32'h00000000} /* (22, 16, 19) {real, imag} */,
  {32'hc6012a5e, 32'h00000000} /* (22, 16, 18) {real, imag} */,
  {32'hc5e81db2, 32'h00000000} /* (22, 16, 17) {real, imag} */,
  {32'hc5eaf86e, 32'h00000000} /* (22, 16, 16) {real, imag} */,
  {32'hc5e93331, 32'h00000000} /* (22, 16, 15) {real, imag} */,
  {32'hc5c3d2e8, 32'h00000000} /* (22, 16, 14) {real, imag} */,
  {32'hc5d1cee9, 32'h00000000} /* (22, 16, 13) {real, imag} */,
  {32'hc5ac225e, 32'h00000000} /* (22, 16, 12) {real, imag} */,
  {32'hc56352d1, 32'h00000000} /* (22, 16, 11) {real, imag} */,
  {32'hc35a63e0, 32'h00000000} /* (22, 16, 10) {real, imag} */,
  {32'h457bef7e, 32'h00000000} /* (22, 16, 9) {real, imag} */,
  {32'h45a21833, 32'h00000000} /* (22, 16, 8) {real, imag} */,
  {32'h45cd9384, 32'h00000000} /* (22, 16, 7) {real, imag} */,
  {32'h45f776d2, 32'h00000000} /* (22, 16, 6) {real, imag} */,
  {32'h45fc85de, 32'h00000000} /* (22, 16, 5) {real, imag} */,
  {32'h460a8a28, 32'h00000000} /* (22, 16, 4) {real, imag} */,
  {32'h461097c0, 32'h00000000} /* (22, 16, 3) {real, imag} */,
  {32'h46001e12, 32'h00000000} /* (22, 16, 2) {real, imag} */,
  {32'h46081190, 32'h00000000} /* (22, 16, 1) {real, imag} */,
  {32'h45fe4ccc, 32'h00000000} /* (22, 16, 0) {real, imag} */,
  {32'h45fa0433, 32'h00000000} /* (22, 15, 31) {real, imag} */,
  {32'h460c0e98, 32'h00000000} /* (22, 15, 30) {real, imag} */,
  {32'h460bf5fb, 32'h00000000} /* (22, 15, 29) {real, imag} */,
  {32'h460cedb2, 32'h00000000} /* (22, 15, 28) {real, imag} */,
  {32'h46038252, 32'h00000000} /* (22, 15, 27) {real, imag} */,
  {32'h45f8df5c, 32'h00000000} /* (22, 15, 26) {real, imag} */,
  {32'h45efd753, 32'h00000000} /* (22, 15, 25) {real, imag} */,
  {32'h45e76184, 32'h00000000} /* (22, 15, 24) {real, imag} */,
  {32'h45b8fd0e, 32'h00000000} /* (22, 15, 23) {real, imag} */,
  {32'h45520ab8, 32'h00000000} /* (22, 15, 22) {real, imag} */,
  {32'hc1835a00, 32'h00000000} /* (22, 15, 21) {real, imag} */,
  {32'hc55ee370, 32'h00000000} /* (22, 15, 20) {real, imag} */,
  {32'hc5bc8652, 32'h00000000} /* (22, 15, 19) {real, imag} */,
  {32'hc5c7f948, 32'h00000000} /* (22, 15, 18) {real, imag} */,
  {32'hc5ee41b2, 32'h00000000} /* (22, 15, 17) {real, imag} */,
  {32'hc5f58278, 32'h00000000} /* (22, 15, 16) {real, imag} */,
  {32'hc5d1b1a7, 32'h00000000} /* (22, 15, 15) {real, imag} */,
  {32'hc5d22a6a, 32'h00000000} /* (22, 15, 14) {real, imag} */,
  {32'hc5b596ca, 32'h00000000} /* (22, 15, 13) {real, imag} */,
  {32'hc5af4e41, 32'h00000000} /* (22, 15, 12) {real, imag} */,
  {32'hc5896e19, 32'h00000000} /* (22, 15, 11) {real, imag} */,
  {32'hc2c20600, 32'h00000000} /* (22, 15, 10) {real, imag} */,
  {32'h455e558a, 32'h00000000} /* (22, 15, 9) {real, imag} */,
  {32'h45c0fcec, 32'h00000000} /* (22, 15, 8) {real, imag} */,
  {32'h45da67ac, 32'h00000000} /* (22, 15, 7) {real, imag} */,
  {32'h45ee19ac, 32'h00000000} /* (22, 15, 6) {real, imag} */,
  {32'h4600c1dd, 32'h00000000} /* (22, 15, 5) {real, imag} */,
  {32'h4612acff, 32'h00000000} /* (22, 15, 4) {real, imag} */,
  {32'h46171ffc, 32'h00000000} /* (22, 15, 3) {real, imag} */,
  {32'h460a0c6d, 32'h00000000} /* (22, 15, 2) {real, imag} */,
  {32'h4606c964, 32'h00000000} /* (22, 15, 1) {real, imag} */,
  {32'h45f329cc, 32'h00000000} /* (22, 15, 0) {real, imag} */,
  {32'h45e406e0, 32'h00000000} /* (22, 14, 31) {real, imag} */,
  {32'h4606ae68, 32'h00000000} /* (22, 14, 30) {real, imag} */,
  {32'h4602b7d1, 32'h00000000} /* (22, 14, 29) {real, imag} */,
  {32'h45f523e2, 32'h00000000} /* (22, 14, 28) {real, imag} */,
  {32'h45f117ec, 32'h00000000} /* (22, 14, 27) {real, imag} */,
  {32'h460403bb, 32'h00000000} /* (22, 14, 26) {real, imag} */,
  {32'h45f2de56, 32'h00000000} /* (22, 14, 25) {real, imag} */,
  {32'h45d29972, 32'h00000000} /* (22, 14, 24) {real, imag} */,
  {32'h45ccf952, 32'h00000000} /* (22, 14, 23) {real, imag} */,
  {32'h458727f6, 32'h00000000} /* (22, 14, 22) {real, imag} */,
  {32'hc2f95e80, 32'h00000000} /* (22, 14, 21) {real, imag} */,
  {32'hc553ac84, 32'h00000000} /* (22, 14, 20) {real, imag} */,
  {32'hc5896a9c, 32'h00000000} /* (22, 14, 19) {real, imag} */,
  {32'hc5c74f05, 32'h00000000} /* (22, 14, 18) {real, imag} */,
  {32'hc5cd0918, 32'h00000000} /* (22, 14, 17) {real, imag} */,
  {32'hc5d9001a, 32'h00000000} /* (22, 14, 16) {real, imag} */,
  {32'hc5e11b20, 32'h00000000} /* (22, 14, 15) {real, imag} */,
  {32'hc5b1ee80, 32'h00000000} /* (22, 14, 14) {real, imag} */,
  {32'hc5baa926, 32'h00000000} /* (22, 14, 13) {real, imag} */,
  {32'hc5a76636, 32'h00000000} /* (22, 14, 12) {real, imag} */,
  {32'hc5254e3c, 32'h00000000} /* (22, 14, 11) {real, imag} */,
  {32'h448f886e, 32'h00000000} /* (22, 14, 10) {real, imag} */,
  {32'h4581c3d6, 32'h00000000} /* (22, 14, 9) {real, imag} */,
  {32'h45bc3836, 32'h00000000} /* (22, 14, 8) {real, imag} */,
  {32'h45e8764e, 32'h00000000} /* (22, 14, 7) {real, imag} */,
  {32'h45e73e90, 32'h00000000} /* (22, 14, 6) {real, imag} */,
  {32'h45e95dac, 32'h00000000} /* (22, 14, 5) {real, imag} */,
  {32'h46054982, 32'h00000000} /* (22, 14, 4) {real, imag} */,
  {32'h460277b9, 32'h00000000} /* (22, 14, 3) {real, imag} */,
  {32'h45f4d135, 32'h00000000} /* (22, 14, 2) {real, imag} */,
  {32'h45fee2da, 32'h00000000} /* (22, 14, 1) {real, imag} */,
  {32'h4604a206, 32'h00000000} /* (22, 14, 0) {real, imag} */,
  {32'h45c1008d, 32'h00000000} /* (22, 13, 31) {real, imag} */,
  {32'h45deca2c, 32'h00000000} /* (22, 13, 30) {real, imag} */,
  {32'h45d8299d, 32'h00000000} /* (22, 13, 29) {real, imag} */,
  {32'h45d414eb, 32'h00000000} /* (22, 13, 28) {real, imag} */,
  {32'h45c14fce, 32'h00000000} /* (22, 13, 27) {real, imag} */,
  {32'h45d6fb22, 32'h00000000} /* (22, 13, 26) {real, imag} */,
  {32'h45c37268, 32'h00000000} /* (22, 13, 25) {real, imag} */,
  {32'h45998502, 32'h00000000} /* (22, 13, 24) {real, imag} */,
  {32'h45844460, 32'h00000000} /* (22, 13, 23) {real, imag} */,
  {32'h45760584, 32'h00000000} /* (22, 13, 22) {real, imag} */,
  {32'h44505c8c, 32'h00000000} /* (22, 13, 21) {real, imag} */,
  {32'hc5335edd, 32'h00000000} /* (22, 13, 20) {real, imag} */,
  {32'hc5a89f72, 32'h00000000} /* (22, 13, 19) {real, imag} */,
  {32'hc5b8ab62, 32'h00000000} /* (22, 13, 18) {real, imag} */,
  {32'hc5c161a8, 32'h00000000} /* (22, 13, 17) {real, imag} */,
  {32'hc5c9b66d, 32'h00000000} /* (22, 13, 16) {real, imag} */,
  {32'hc5a84159, 32'h00000000} /* (22, 13, 15) {real, imag} */,
  {32'hc598f726, 32'h00000000} /* (22, 13, 14) {real, imag} */,
  {32'hc58c3039, 32'h00000000} /* (22, 13, 13) {real, imag} */,
  {32'hc560a472, 32'h00000000} /* (22, 13, 12) {real, imag} */,
  {32'hc51d05ff, 32'h00000000} /* (22, 13, 11) {real, imag} */,
  {32'h44e56346, 32'h00000000} /* (22, 13, 10) {real, imag} */,
  {32'h45991108, 32'h00000000} /* (22, 13, 9) {real, imag} */,
  {32'h45ca6944, 32'h00000000} /* (22, 13, 8) {real, imag} */,
  {32'h45e118fe, 32'h00000000} /* (22, 13, 7) {real, imag} */,
  {32'h45d5af52, 32'h00000000} /* (22, 13, 6) {real, imag} */,
  {32'h45ea478a, 32'h00000000} /* (22, 13, 5) {real, imag} */,
  {32'h45db7c14, 32'h00000000} /* (22, 13, 4) {real, imag} */,
  {32'h45d526b8, 32'h00000000} /* (22, 13, 3) {real, imag} */,
  {32'h45ca0a34, 32'h00000000} /* (22, 13, 2) {real, imag} */,
  {32'h45d4cb08, 32'h00000000} /* (22, 13, 1) {real, imag} */,
  {32'h45d10dd7, 32'h00000000} /* (22, 13, 0) {real, imag} */,
  {32'h4589c1f5, 32'h00000000} /* (22, 12, 31) {real, imag} */,
  {32'h45787b31, 32'h00000000} /* (22, 12, 30) {real, imag} */,
  {32'h4585c85d, 32'h00000000} /* (22, 12, 29) {real, imag} */,
  {32'h45a9501a, 32'h00000000} /* (22, 12, 28) {real, imag} */,
  {32'h459df05e, 32'h00000000} /* (22, 12, 27) {real, imag} */,
  {32'h457a51a8, 32'h00000000} /* (22, 12, 26) {real, imag} */,
  {32'h456e9b99, 32'h00000000} /* (22, 12, 25) {real, imag} */,
  {32'h4570fed0, 32'h00000000} /* (22, 12, 24) {real, imag} */,
  {32'h458eee4a, 32'h00000000} /* (22, 12, 23) {real, imag} */,
  {32'h452c20c4, 32'h00000000} /* (22, 12, 22) {real, imag} */,
  {32'h42b2e0e0, 32'h00000000} /* (22, 12, 21) {real, imag} */,
  {32'hc5295088, 32'h00000000} /* (22, 12, 20) {real, imag} */,
  {32'hc5b1dfec, 32'h00000000} /* (22, 12, 19) {real, imag} */,
  {32'hc5a9ba08, 32'h00000000} /* (22, 12, 18) {real, imag} */,
  {32'hc596071a, 32'h00000000} /* (22, 12, 17) {real, imag} */,
  {32'hc5938295, 32'h00000000} /* (22, 12, 16) {real, imag} */,
  {32'hc567bacc, 32'h00000000} /* (22, 12, 15) {real, imag} */,
  {32'hc56a5d77, 32'h00000000} /* (22, 12, 14) {real, imag} */,
  {32'hc5414764, 32'h00000000} /* (22, 12, 13) {real, imag} */,
  {32'hc54cc4d4, 32'h00000000} /* (22, 12, 12) {real, imag} */,
  {32'hc483c558, 32'h00000000} /* (22, 12, 11) {real, imag} */,
  {32'h4519c9dc, 32'h00000000} /* (22, 12, 10) {real, imag} */,
  {32'h45460e53, 32'h00000000} /* (22, 12, 9) {real, imag} */,
  {32'h4596b9fc, 32'h00000000} /* (22, 12, 8) {real, imag} */,
  {32'h45b88a16, 32'h00000000} /* (22, 12, 7) {real, imag} */,
  {32'h45b89b96, 32'h00000000} /* (22, 12, 6) {real, imag} */,
  {32'h45c44b1e, 32'h00000000} /* (22, 12, 5) {real, imag} */,
  {32'h459aefae, 32'h00000000} /* (22, 12, 4) {real, imag} */,
  {32'h459820be, 32'h00000000} /* (22, 12, 3) {real, imag} */,
  {32'h45945140, 32'h00000000} /* (22, 12, 2) {real, imag} */,
  {32'h4592adf2, 32'h00000000} /* (22, 12, 1) {real, imag} */,
  {32'h45553f5c, 32'h00000000} /* (22, 12, 0) {real, imag} */,
  {32'h4494c1ce, 32'h00000000} /* (22, 11, 31) {real, imag} */,
  {32'h4485efb8, 32'h00000000} /* (22, 11, 30) {real, imag} */,
  {32'h449c9f0f, 32'h00000000} /* (22, 11, 29) {real, imag} */,
  {32'h44a5f240, 32'h00000000} /* (22, 11, 28) {real, imag} */,
  {32'h44d7fe38, 32'h00000000} /* (22, 11, 27) {real, imag} */,
  {32'h450d467e, 32'h00000000} /* (22, 11, 26) {real, imag} */,
  {32'h447b5db4, 32'h00000000} /* (22, 11, 25) {real, imag} */,
  {32'h44d7e531, 32'h00000000} /* (22, 11, 24) {real, imag} */,
  {32'h44c72a40, 32'h00000000} /* (22, 11, 23) {real, imag} */,
  {32'h4429d4b3, 32'h00000000} /* (22, 11, 22) {real, imag} */,
  {32'hc4964acd, 32'h00000000} /* (22, 11, 21) {real, imag} */,
  {32'hc54c7e23, 32'h00000000} /* (22, 11, 20) {real, imag} */,
  {32'hc54f2b6d, 32'h00000000} /* (22, 11, 19) {real, imag} */,
  {32'hc53b61c6, 32'h00000000} /* (22, 11, 18) {real, imag} */,
  {32'hc531136d, 32'h00000000} /* (22, 11, 17) {real, imag} */,
  {32'hc52595b4, 32'h00000000} /* (22, 11, 16) {real, imag} */,
  {32'hc50f4846, 32'h00000000} /* (22, 11, 15) {real, imag} */,
  {32'hc4ecc6cc, 32'h00000000} /* (22, 11, 14) {real, imag} */,
  {32'hc4cd4999, 32'h00000000} /* (22, 11, 13) {real, imag} */,
  {32'hc4ef3e18, 32'h00000000} /* (22, 11, 12) {real, imag} */,
  {32'hc3c0b076, 32'h00000000} /* (22, 11, 11) {real, imag} */,
  {32'h44fad274, 32'h00000000} /* (22, 11, 10) {real, imag} */,
  {32'h450ac40d, 32'h00000000} /* (22, 11, 9) {real, imag} */,
  {32'h459007c6, 32'h00000000} /* (22, 11, 8) {real, imag} */,
  {32'h45890da2, 32'h00000000} /* (22, 11, 7) {real, imag} */,
  {32'h45196bc3, 32'h00000000} /* (22, 11, 6) {real, imag} */,
  {32'h4539f252, 32'h00000000} /* (22, 11, 5) {real, imag} */,
  {32'h452b2d3f, 32'h00000000} /* (22, 11, 4) {real, imag} */,
  {32'h451671f7, 32'h00000000} /* (22, 11, 3) {real, imag} */,
  {32'h44d9c0c4, 32'h00000000} /* (22, 11, 2) {real, imag} */,
  {32'h44f58682, 32'h00000000} /* (22, 11, 1) {real, imag} */,
  {32'h44ca30ed, 32'h00000000} /* (22, 11, 0) {real, imag} */,
  {32'hc510872c, 32'h00000000} /* (22, 10, 31) {real, imag} */,
  {32'hc53c9090, 32'h00000000} /* (22, 10, 30) {real, imag} */,
  {32'hc5492c36, 32'h00000000} /* (22, 10, 29) {real, imag} */,
  {32'hc528eabc, 32'h00000000} /* (22, 10, 28) {real, imag} */,
  {32'hc5146139, 32'h00000000} /* (22, 10, 27) {real, imag} */,
  {32'hc504fdc0, 32'h00000000} /* (22, 10, 26) {real, imag} */,
  {32'hc523cdf6, 32'h00000000} /* (22, 10, 25) {real, imag} */,
  {32'hc5231cae, 32'h00000000} /* (22, 10, 24) {real, imag} */,
  {32'hc52ba19e, 32'h00000000} /* (22, 10, 23) {real, imag} */,
  {32'hc502c22c, 32'h00000000} /* (22, 10, 22) {real, imag} */,
  {32'hc550b799, 32'h00000000} /* (22, 10, 21) {real, imag} */,
  {32'hc4acdec4, 32'h00000000} /* (22, 10, 20) {real, imag} */,
  {32'h417b2cc0, 32'h00000000} /* (22, 10, 19) {real, imag} */,
  {32'hc4066ba0, 32'h00000000} /* (22, 10, 18) {real, imag} */,
  {32'h43bdac4b, 32'h00000000} /* (22, 10, 17) {real, imag} */,
  {32'h4421335f, 32'h00000000} /* (22, 10, 16) {real, imag} */,
  {32'h43f1053c, 32'h00000000} /* (22, 10, 15) {real, imag} */,
  {32'h44538e9a, 32'h00000000} /* (22, 10, 14) {real, imag} */,
  {32'h4484cd5c, 32'h00000000} /* (22, 10, 13) {real, imag} */,
  {32'h44b8e638, 32'h00000000} /* (22, 10, 12) {real, imag} */,
  {32'h44e17856, 32'h00000000} /* (22, 10, 11) {real, imag} */,
  {32'h44a99d62, 32'h00000000} /* (22, 10, 10) {real, imag} */,
  {32'h44165f68, 32'h00000000} /* (22, 10, 9) {real, imag} */,
  {32'h44a1e426, 32'h00000000} /* (22, 10, 8) {real, imag} */,
  {32'h44281ef8, 32'h00000000} /* (22, 10, 7) {real, imag} */,
  {32'hc387d37a, 32'h00000000} /* (22, 10, 6) {real, imag} */,
  {32'hc4435014, 32'h00000000} /* (22, 10, 5) {real, imag} */,
  {32'hc4cf4e38, 32'h00000000} /* (22, 10, 4) {real, imag} */,
  {32'hc4b44456, 32'h00000000} /* (22, 10, 3) {real, imag} */,
  {32'hc4f8d2b4, 32'h00000000} /* (22, 10, 2) {real, imag} */,
  {32'hc498dcef, 32'h00000000} /* (22, 10, 1) {real, imag} */,
  {32'hc4c17eb6, 32'h00000000} /* (22, 10, 0) {real, imag} */,
  {32'hc59cb822, 32'h00000000} /* (22, 9, 31) {real, imag} */,
  {32'hc5c60b4e, 32'h00000000} /* (22, 9, 30) {real, imag} */,
  {32'hc5c6c4c8, 32'h00000000} /* (22, 9, 29) {real, imag} */,
  {32'hc5c0894a, 32'h00000000} /* (22, 9, 28) {real, imag} */,
  {32'hc5c1a26e, 32'h00000000} /* (22, 9, 27) {real, imag} */,
  {32'hc5b831b0, 32'h00000000} /* (22, 9, 26) {real, imag} */,
  {32'hc5a3ad2c, 32'h00000000} /* (22, 9, 25) {real, imag} */,
  {32'hc5abf5b2, 32'h00000000} /* (22, 9, 24) {real, imag} */,
  {32'hc5a402f8, 32'h00000000} /* (22, 9, 23) {real, imag} */,
  {32'hc58c13ec, 32'h00000000} /* (22, 9, 22) {real, imag} */,
  {32'hc577791e, 32'h00000000} /* (22, 9, 21) {real, imag} */,
  {32'hc4b1b4d0, 32'h00000000} /* (22, 9, 20) {real, imag} */,
  {32'h424cbf40, 32'h00000000} /* (22, 9, 19) {real, imag} */,
  {32'h450b21ad, 32'h00000000} /* (22, 9, 18) {real, imag} */,
  {32'h4510a2a9, 32'h00000000} /* (22, 9, 17) {real, imag} */,
  {32'h4555e818, 32'h00000000} /* (22, 9, 16) {real, imag} */,
  {32'h455937f0, 32'h00000000} /* (22, 9, 15) {real, imag} */,
  {32'h453c26df, 32'h00000000} /* (22, 9, 14) {real, imag} */,
  {32'h457c0199, 32'h00000000} /* (22, 9, 13) {real, imag} */,
  {32'h4558d03f, 32'h00000000} /* (22, 9, 12) {real, imag} */,
  {32'h454336cf, 32'h00000000} /* (22, 9, 11) {real, imag} */,
  {32'h4497996a, 32'h00000000} /* (22, 9, 10) {real, imag} */,
  {32'hc3b7f8d8, 32'h00000000} /* (22, 9, 9) {real, imag} */,
  {32'hc4827566, 32'h00000000} /* (22, 9, 8) {real, imag} */,
  {32'hc5292434, 32'h00000000} /* (22, 9, 7) {real, imag} */,
  {32'hc54a220e, 32'h00000000} /* (22, 9, 6) {real, imag} */,
  {32'hc54f8ff8, 32'h00000000} /* (22, 9, 5) {real, imag} */,
  {32'hc5997d09, 32'h00000000} /* (22, 9, 4) {real, imag} */,
  {32'hc5bcb738, 32'h00000000} /* (22, 9, 3) {real, imag} */,
  {32'hc592ac40, 32'h00000000} /* (22, 9, 2) {real, imag} */,
  {32'hc5bb998a, 32'h00000000} /* (22, 9, 1) {real, imag} */,
  {32'hc5aaab58, 32'h00000000} /* (22, 9, 0) {real, imag} */,
  {32'hc5eac3bc, 32'h00000000} /* (22, 8, 31) {real, imag} */,
  {32'hc606693c, 32'h00000000} /* (22, 8, 30) {real, imag} */,
  {32'hc607e596, 32'h00000000} /* (22, 8, 29) {real, imag} */,
  {32'hc6066759, 32'h00000000} /* (22, 8, 28) {real, imag} */,
  {32'hc6064510, 32'h00000000} /* (22, 8, 27) {real, imag} */,
  {32'hc60c904b, 32'h00000000} /* (22, 8, 26) {real, imag} */,
  {32'hc6036e40, 32'h00000000} /* (22, 8, 25) {real, imag} */,
  {32'hc611bf1e, 32'h00000000} /* (22, 8, 24) {real, imag} */,
  {32'hc5fd3180, 32'h00000000} /* (22, 8, 23) {real, imag} */,
  {32'hc5b9deba, 32'h00000000} /* (22, 8, 22) {real, imag} */,
  {32'hc58b8f88, 32'h00000000} /* (22, 8, 21) {real, imag} */,
  {32'hc4ad4ce6, 32'h00000000} /* (22, 8, 20) {real, imag} */,
  {32'h4403a43c, 32'h00000000} /* (22, 8, 19) {real, imag} */,
  {32'h4529cf60, 32'h00000000} /* (22, 8, 18) {real, imag} */,
  {32'h4575c37c, 32'h00000000} /* (22, 8, 17) {real, imag} */,
  {32'h455894c7, 32'h00000000} /* (22, 8, 16) {real, imag} */,
  {32'h458e6d7c, 32'h00000000} /* (22, 8, 15) {real, imag} */,
  {32'h45bc564c, 32'h00000000} /* (22, 8, 14) {real, imag} */,
  {32'h459483fc, 32'h00000000} /* (22, 8, 13) {real, imag} */,
  {32'h458742c8, 32'h00000000} /* (22, 8, 12) {real, imag} */,
  {32'h454bdc69, 32'h00000000} /* (22, 8, 11) {real, imag} */,
  {32'h44a246a8, 32'h00000000} /* (22, 8, 10) {real, imag} */,
  {32'hc4a5faec, 32'h00000000} /* (22, 8, 9) {real, imag} */,
  {32'hc51a20f2, 32'h00000000} /* (22, 8, 8) {real, imag} */,
  {32'hc54d3121, 32'h00000000} /* (22, 8, 7) {real, imag} */,
  {32'hc58f7e3a, 32'h00000000} /* (22, 8, 6) {real, imag} */,
  {32'hc5a83fc0, 32'h00000000} /* (22, 8, 5) {real, imag} */,
  {32'hc5ceee88, 32'h00000000} /* (22, 8, 4) {real, imag} */,
  {32'hc5c95a46, 32'h00000000} /* (22, 8, 3) {real, imag} */,
  {32'hc5ec7c14, 32'h00000000} /* (22, 8, 2) {real, imag} */,
  {32'hc5ea6ab6, 32'h00000000} /* (22, 8, 1) {real, imag} */,
  {32'hc5c2a5ca, 32'h00000000} /* (22, 8, 0) {real, imag} */,
  {32'hc609c7ad, 32'h00000000} /* (22, 7, 31) {real, imag} */,
  {32'hc6250924, 32'h00000000} /* (22, 7, 30) {real, imag} */,
  {32'hc6258ded, 32'h00000000} /* (22, 7, 29) {real, imag} */,
  {32'hc629cfa1, 32'h00000000} /* (22, 7, 28) {real, imag} */,
  {32'hc62466a6, 32'h00000000} /* (22, 7, 27) {real, imag} */,
  {32'hc625aee0, 32'h00000000} /* (22, 7, 26) {real, imag} */,
  {32'hc636bf18, 32'h00000000} /* (22, 7, 25) {real, imag} */,
  {32'hc61c1818, 32'h00000000} /* (22, 7, 24) {real, imag} */,
  {32'hc60ea6b0, 32'h00000000} /* (22, 7, 23) {real, imag} */,
  {32'hc5f25c9a, 32'h00000000} /* (22, 7, 22) {real, imag} */,
  {32'hc5b002e0, 32'h00000000} /* (22, 7, 21) {real, imag} */,
  {32'hc502b3e8, 32'h00000000} /* (22, 7, 20) {real, imag} */,
  {32'h43e2a670, 32'h00000000} /* (22, 7, 19) {real, imag} */,
  {32'h44c7621c, 32'h00000000} /* (22, 7, 18) {real, imag} */,
  {32'h456f9ad9, 32'h00000000} /* (22, 7, 17) {real, imag} */,
  {32'h457bb9fc, 32'h00000000} /* (22, 7, 16) {real, imag} */,
  {32'h459c6238, 32'h00000000} /* (22, 7, 15) {real, imag} */,
  {32'h45bf97d5, 32'h00000000} /* (22, 7, 14) {real, imag} */,
  {32'h45c1f6c2, 32'h00000000} /* (22, 7, 13) {real, imag} */,
  {32'h45a4d82c, 32'h00000000} /* (22, 7, 12) {real, imag} */,
  {32'h457efa70, 32'h00000000} /* (22, 7, 11) {real, imag} */,
  {32'h44a9bce4, 32'h00000000} /* (22, 7, 10) {real, imag} */,
  {32'hc2c77ec0, 32'h00000000} /* (22, 7, 9) {real, imag} */,
  {32'hc503ab29, 32'h00000000} /* (22, 7, 8) {real, imag} */,
  {32'hc54e78e0, 32'h00000000} /* (22, 7, 7) {real, imag} */,
  {32'hc5941048, 32'h00000000} /* (22, 7, 6) {real, imag} */,
  {32'hc5ef3fcc, 32'h00000000} /* (22, 7, 5) {real, imag} */,
  {32'hc5d7ddb8, 32'h00000000} /* (22, 7, 4) {real, imag} */,
  {32'hc601a3d6, 32'h00000000} /* (22, 7, 3) {real, imag} */,
  {32'hc616db02, 32'h00000000} /* (22, 7, 2) {real, imag} */,
  {32'hc6048d0a, 32'h00000000} /* (22, 7, 1) {real, imag} */,
  {32'hc604aca1, 32'h00000000} /* (22, 7, 0) {real, imag} */,
  {32'hc6202633, 32'h00000000} /* (22, 6, 31) {real, imag} */,
  {32'hc628cfa1, 32'h00000000} /* (22, 6, 30) {real, imag} */,
  {32'hc6360aaf, 32'h00000000} /* (22, 6, 29) {real, imag} */,
  {32'hc6433b4b, 32'h00000000} /* (22, 6, 28) {real, imag} */,
  {32'hc641d98d, 32'h00000000} /* (22, 6, 27) {real, imag} */,
  {32'hc6421792, 32'h00000000} /* (22, 6, 26) {real, imag} */,
  {32'hc63b5709, 32'h00000000} /* (22, 6, 25) {real, imag} */,
  {32'hc6232a1a, 32'h00000000} /* (22, 6, 24) {real, imag} */,
  {32'hc6196bd6, 32'h00000000} /* (22, 6, 23) {real, imag} */,
  {32'hc607ebac, 32'h00000000} /* (22, 6, 22) {real, imag} */,
  {32'hc5c6d554, 32'h00000000} /* (22, 6, 21) {real, imag} */,
  {32'hc5327ec2, 32'h00000000} /* (22, 6, 20) {real, imag} */,
  {32'hc4a1effe, 32'h00000000} /* (22, 6, 19) {real, imag} */,
  {32'h44120438, 32'h00000000} /* (22, 6, 18) {real, imag} */,
  {32'h451f979c, 32'h00000000} /* (22, 6, 17) {real, imag} */,
  {32'h45767965, 32'h00000000} /* (22, 6, 16) {real, imag} */,
  {32'h45bf648c, 32'h00000000} /* (22, 6, 15) {real, imag} */,
  {32'h45ba6846, 32'h00000000} /* (22, 6, 14) {real, imag} */,
  {32'h45c9e3d2, 32'h00000000} /* (22, 6, 13) {real, imag} */,
  {32'h45c7756a, 32'h00000000} /* (22, 6, 12) {real, imag} */,
  {32'h45910fa2, 32'h00000000} /* (22, 6, 11) {real, imag} */,
  {32'h45197d0c, 32'h00000000} /* (22, 6, 10) {real, imag} */,
  {32'h4398b7a0, 32'h00000000} /* (22, 6, 9) {real, imag} */,
  {32'hc493b750, 32'h00000000} /* (22, 6, 8) {real, imag} */,
  {32'hc5067c52, 32'h00000000} /* (22, 6, 7) {real, imag} */,
  {32'hc5a24c58, 32'h00000000} /* (22, 6, 6) {real, imag} */,
  {32'hc5acf728, 32'h00000000} /* (22, 6, 5) {real, imag} */,
  {32'hc5eb37c3, 32'h00000000} /* (22, 6, 4) {real, imag} */,
  {32'hc60abe39, 32'h00000000} /* (22, 6, 3) {real, imag} */,
  {32'hc60ef0ba, 32'h00000000} /* (22, 6, 2) {real, imag} */,
  {32'hc61ca40b, 32'h00000000} /* (22, 6, 1) {real, imag} */,
  {32'hc61fae71, 32'h00000000} /* (22, 6, 0) {real, imag} */,
  {32'hc631de72, 32'h00000000} /* (22, 5, 31) {real, imag} */,
  {32'hc64f9ef7, 32'h00000000} /* (22, 5, 30) {real, imag} */,
  {32'hc648e54e, 32'h00000000} /* (22, 5, 29) {real, imag} */,
  {32'hc655ee54, 32'h00000000} /* (22, 5, 28) {real, imag} */,
  {32'hc657aaae, 32'h00000000} /* (22, 5, 27) {real, imag} */,
  {32'hc64e712f, 32'h00000000} /* (22, 5, 26) {real, imag} */,
  {32'hc64ea947, 32'h00000000} /* (22, 5, 25) {real, imag} */,
  {32'hc641b720, 32'h00000000} /* (22, 5, 24) {real, imag} */,
  {32'hc6255a56, 32'h00000000} /* (22, 5, 23) {real, imag} */,
  {32'hc6139a1a, 32'h00000000} /* (22, 5, 22) {real, imag} */,
  {32'hc5ef9451, 32'h00000000} /* (22, 5, 21) {real, imag} */,
  {32'hc5ac1189, 32'h00000000} /* (22, 5, 20) {real, imag} */,
  {32'hc5537185, 32'h00000000} /* (22, 5, 19) {real, imag} */,
  {32'hc4bd5e30, 32'h00000000} /* (22, 5, 18) {real, imag} */,
  {32'h4312c860, 32'h00000000} /* (22, 5, 17) {real, imag} */,
  {32'h44b13478, 32'h00000000} /* (22, 5, 16) {real, imag} */,
  {32'h458cd0a3, 32'h00000000} /* (22, 5, 15) {real, imag} */,
  {32'h45ce244e, 32'h00000000} /* (22, 5, 14) {real, imag} */,
  {32'h45cb782c, 32'h00000000} /* (22, 5, 13) {real, imag} */,
  {32'h45be4198, 32'h00000000} /* (22, 5, 12) {real, imag} */,
  {32'h45bef6d8, 32'h00000000} /* (22, 5, 11) {real, imag} */,
  {32'h45a73432, 32'h00000000} /* (22, 5, 10) {real, imag} */,
  {32'h44ed42b8, 32'h00000000} /* (22, 5, 9) {real, imag} */,
  {32'h44a5e42c, 32'h00000000} /* (22, 5, 8) {real, imag} */,
  {32'h431a2b40, 32'h00000000} /* (22, 5, 7) {real, imag} */,
  {32'hc4ef87d4, 32'h00000000} /* (22, 5, 6) {real, imag} */,
  {32'hc5ac110b, 32'h00000000} /* (22, 5, 5) {real, imag} */,
  {32'hc5e360fb, 32'h00000000} /* (22, 5, 4) {real, imag} */,
  {32'hc61dfca3, 32'h00000000} /* (22, 5, 3) {real, imag} */,
  {32'hc6276350, 32'h00000000} /* (22, 5, 2) {real, imag} */,
  {32'hc620168c, 32'h00000000} /* (22, 5, 1) {real, imag} */,
  {32'hc6295e0b, 32'h00000000} /* (22, 5, 0) {real, imag} */,
  {32'hc63ee352, 32'h00000000} /* (22, 4, 31) {real, imag} */,
  {32'hc65105a5, 32'h00000000} /* (22, 4, 30) {real, imag} */,
  {32'hc65da263, 32'h00000000} /* (22, 4, 29) {real, imag} */,
  {32'hc65d6ddb, 32'h00000000} /* (22, 4, 28) {real, imag} */,
  {32'hc66bad4e, 32'h00000000} /* (22, 4, 27) {real, imag} */,
  {32'hc65cff39, 32'h00000000} /* (22, 4, 26) {real, imag} */,
  {32'hc6522943, 32'h00000000} /* (22, 4, 25) {real, imag} */,
  {32'hc649c1eb, 32'h00000000} /* (22, 4, 24) {real, imag} */,
  {32'hc6303276, 32'h00000000} /* (22, 4, 23) {real, imag} */,
  {32'hc619995d, 32'h00000000} /* (22, 4, 22) {real, imag} */,
  {32'hc6035559, 32'h00000000} /* (22, 4, 21) {real, imag} */,
  {32'hc5dbb02c, 32'h00000000} /* (22, 4, 20) {real, imag} */,
  {32'hc5ab58d7, 32'h00000000} /* (22, 4, 19) {real, imag} */,
  {32'hc5421104, 32'h00000000} /* (22, 4, 18) {real, imag} */,
  {32'hc495d35c, 32'h00000000} /* (22, 4, 17) {real, imag} */,
  {32'h43b5d7b0, 32'h00000000} /* (22, 4, 16) {real, imag} */,
  {32'h45768436, 32'h00000000} /* (22, 4, 15) {real, imag} */,
  {32'h45be00ce, 32'h00000000} /* (22, 4, 14) {real, imag} */,
  {32'h45d0c972, 32'h00000000} /* (22, 4, 13) {real, imag} */,
  {32'h45cd2d72, 32'h00000000} /* (22, 4, 12) {real, imag} */,
  {32'h45d6955b, 32'h00000000} /* (22, 4, 11) {real, imag} */,
  {32'h45af5842, 32'h00000000} /* (22, 4, 10) {real, imag} */,
  {32'h45a65682, 32'h00000000} /* (22, 4, 9) {real, imag} */,
  {32'h4587a556, 32'h00000000} /* (22, 4, 8) {real, imag} */,
  {32'h449abb5c, 32'h00000000} /* (22, 4, 7) {real, imag} */,
  {32'hc44e28d0, 32'h00000000} /* (22, 4, 6) {real, imag} */,
  {32'hc59608ca, 32'h00000000} /* (22, 4, 5) {real, imag} */,
  {32'hc5f5e090, 32'h00000000} /* (22, 4, 4) {real, imag} */,
  {32'hc617a100, 32'h00000000} /* (22, 4, 3) {real, imag} */,
  {32'hc626724f, 32'h00000000} /* (22, 4, 2) {real, imag} */,
  {32'hc62d4266, 32'h00000000} /* (22, 4, 1) {real, imag} */,
  {32'hc6374ca6, 32'h00000000} /* (22, 4, 0) {real, imag} */,
  {32'hc63f5749, 32'h00000000} /* (22, 3, 31) {real, imag} */,
  {32'hc6554f1f, 32'h00000000} /* (22, 3, 30) {real, imag} */,
  {32'hc65c11e6, 32'h00000000} /* (22, 3, 29) {real, imag} */,
  {32'hc6681611, 32'h00000000} /* (22, 3, 28) {real, imag} */,
  {32'hc674c5a5, 32'h00000000} /* (22, 3, 27) {real, imag} */,
  {32'hc66061fa, 32'h00000000} /* (22, 3, 26) {real, imag} */,
  {32'hc6622f14, 32'h00000000} /* (22, 3, 25) {real, imag} */,
  {32'hc641b834, 32'h00000000} /* (22, 3, 24) {real, imag} */,
  {32'hc64b2d2e, 32'h00000000} /* (22, 3, 23) {real, imag} */,
  {32'hc625e892, 32'h00000000} /* (22, 3, 22) {real, imag} */,
  {32'hc611139e, 32'h00000000} /* (22, 3, 21) {real, imag} */,
  {32'hc5f40089, 32'h00000000} /* (22, 3, 20) {real, imag} */,
  {32'hc59a4b99, 32'h00000000} /* (22, 3, 19) {real, imag} */,
  {32'hc579e39a, 32'h00000000} /* (22, 3, 18) {real, imag} */,
  {32'hc52673da, 32'h00000000} /* (22, 3, 17) {real, imag} */,
  {32'h437dba00, 32'h00000000} /* (22, 3, 16) {real, imag} */,
  {32'h454d9708, 32'h00000000} /* (22, 3, 15) {real, imag} */,
  {32'h45c91e96, 32'h00000000} /* (22, 3, 14) {real, imag} */,
  {32'h45dc5fa1, 32'h00000000} /* (22, 3, 13) {real, imag} */,
  {32'h45d2ce06, 32'h00000000} /* (22, 3, 12) {real, imag} */,
  {32'h45d827f6, 32'h00000000} /* (22, 3, 11) {real, imag} */,
  {32'h45d26b41, 32'h00000000} /* (22, 3, 10) {real, imag} */,
  {32'h4597bc8c, 32'h00000000} /* (22, 3, 9) {real, imag} */,
  {32'h455aa5b0, 32'h00000000} /* (22, 3, 8) {real, imag} */,
  {32'h44f3ed8c, 32'h00000000} /* (22, 3, 7) {real, imag} */,
  {32'hc3a46490, 32'h00000000} /* (22, 3, 6) {real, imag} */,
  {32'hc59d5eba, 32'h00000000} /* (22, 3, 5) {real, imag} */,
  {32'hc605c94b, 32'h00000000} /* (22, 3, 4) {real, imag} */,
  {32'hc627d336, 32'h00000000} /* (22, 3, 3) {real, imag} */,
  {32'hc6435d5e, 32'h00000000} /* (22, 3, 2) {real, imag} */,
  {32'hc639c824, 32'h00000000} /* (22, 3, 1) {real, imag} */,
  {32'hc63ad7b2, 32'h00000000} /* (22, 3, 0) {real, imag} */,
  {32'hc6463336, 32'h00000000} /* (22, 2, 31) {real, imag} */,
  {32'hc66027b6, 32'h00000000} /* (22, 2, 30) {real, imag} */,
  {32'hc66bdab1, 32'h00000000} /* (22, 2, 29) {real, imag} */,
  {32'hc6605386, 32'h00000000} /* (22, 2, 28) {real, imag} */,
  {32'hc65eb511, 32'h00000000} /* (22, 2, 27) {real, imag} */,
  {32'hc6599a8c, 32'h00000000} /* (22, 2, 26) {real, imag} */,
  {32'hc6536b06, 32'h00000000} /* (22, 2, 25) {real, imag} */,
  {32'hc647b4f9, 32'h00000000} /* (22, 2, 24) {real, imag} */,
  {32'hc644f97b, 32'h00000000} /* (22, 2, 23) {real, imag} */,
  {32'hc61ec001, 32'h00000000} /* (22, 2, 22) {real, imag} */,
  {32'hc60a46b6, 32'h00000000} /* (22, 2, 21) {real, imag} */,
  {32'hc5e492ca, 32'h00000000} /* (22, 2, 20) {real, imag} */,
  {32'hc5b58d1d, 32'h00000000} /* (22, 2, 19) {real, imag} */,
  {32'hc57b8bd2, 32'h00000000} /* (22, 2, 18) {real, imag} */,
  {32'hc51196a6, 32'h00000000} /* (22, 2, 17) {real, imag} */,
  {32'h432ce240, 32'h00000000} /* (22, 2, 16) {real, imag} */,
  {32'h453ec1e2, 32'h00000000} /* (22, 2, 15) {real, imag} */,
  {32'h45c3ce4c, 32'h00000000} /* (22, 2, 14) {real, imag} */,
  {32'h45c5ae22, 32'h00000000} /* (22, 2, 13) {real, imag} */,
  {32'h45c81351, 32'h00000000} /* (22, 2, 12) {real, imag} */,
  {32'h45c5fcae, 32'h00000000} /* (22, 2, 11) {real, imag} */,
  {32'h459cf3f8, 32'h00000000} /* (22, 2, 10) {real, imag} */,
  {32'h459138fd, 32'h00000000} /* (22, 2, 9) {real, imag} */,
  {32'h4562f114, 32'h00000000} /* (22, 2, 8) {real, imag} */,
  {32'h44a8b468, 32'h00000000} /* (22, 2, 7) {real, imag} */,
  {32'hc4750d30, 32'h00000000} /* (22, 2, 6) {real, imag} */,
  {32'hc58c48bd, 32'h00000000} /* (22, 2, 5) {real, imag} */,
  {32'hc5eb047c, 32'h00000000} /* (22, 2, 4) {real, imag} */,
  {32'hc6183978, 32'h00000000} /* (22, 2, 3) {real, imag} */,
  {32'hc64170c4, 32'h00000000} /* (22, 2, 2) {real, imag} */,
  {32'hc64a16f0, 32'h00000000} /* (22, 2, 1) {real, imag} */,
  {32'hc6353e59, 32'h00000000} /* (22, 2, 0) {real, imag} */,
  {32'hc64018a4, 32'h00000000} /* (22, 1, 31) {real, imag} */,
  {32'hc64b5664, 32'h00000000} /* (22, 1, 30) {real, imag} */,
  {32'hc655c0f5, 32'h00000000} /* (22, 1, 29) {real, imag} */,
  {32'hc659dca4, 32'h00000000} /* (22, 1, 28) {real, imag} */,
  {32'hc6555a8e, 32'h00000000} /* (22, 1, 27) {real, imag} */,
  {32'hc6632045, 32'h00000000} /* (22, 1, 26) {real, imag} */,
  {32'hc65c8107, 32'h00000000} /* (22, 1, 25) {real, imag} */,
  {32'hc642b6a6, 32'h00000000} /* (22, 1, 24) {real, imag} */,
  {32'hc635353e, 32'h00000000} /* (22, 1, 23) {real, imag} */,
  {32'hc620d5f0, 32'h00000000} /* (22, 1, 22) {real, imag} */,
  {32'hc5fdb0a6, 32'h00000000} /* (22, 1, 21) {real, imag} */,
  {32'hc5d30317, 32'h00000000} /* (22, 1, 20) {real, imag} */,
  {32'hc5a3aae3, 32'h00000000} /* (22, 1, 19) {real, imag} */,
  {32'hc555696f, 32'h00000000} /* (22, 1, 18) {real, imag} */,
  {32'hc52f3b76, 32'h00000000} /* (22, 1, 17) {real, imag} */,
  {32'h438dda30, 32'h00000000} /* (22, 1, 16) {real, imag} */,
  {32'h455278b6, 32'h00000000} /* (22, 1, 15) {real, imag} */,
  {32'h45bc62a3, 32'h00000000} /* (22, 1, 14) {real, imag} */,
  {32'h45c9f22e, 32'h00000000} /* (22, 1, 13) {real, imag} */,
  {32'h45bceefb, 32'h00000000} /* (22, 1, 12) {real, imag} */,
  {32'h45a9afcc, 32'h00000000} /* (22, 1, 11) {real, imag} */,
  {32'h458e8ce6, 32'h00000000} /* (22, 1, 10) {real, imag} */,
  {32'h456ece24, 32'h00000000} /* (22, 1, 9) {real, imag} */,
  {32'h45396c2e, 32'h00000000} /* (22, 1, 8) {real, imag} */,
  {32'h44422b58, 32'h00000000} /* (22, 1, 7) {real, imag} */,
  {32'hc4e09cd8, 32'h00000000} /* (22, 1, 6) {real, imag} */,
  {32'hc58dc85e, 32'h00000000} /* (22, 1, 5) {real, imag} */,
  {32'hc5f41a27, 32'h00000000} /* (22, 1, 4) {real, imag} */,
  {32'hc61960f2, 32'h00000000} /* (22, 1, 3) {real, imag} */,
  {32'hc6332a04, 32'h00000000} /* (22, 1, 2) {real, imag} */,
  {32'hc6357a50, 32'h00000000} /* (22, 1, 1) {real, imag} */,
  {32'hc639095a, 32'h00000000} /* (22, 1, 0) {real, imag} */,
  {32'hc636bfa2, 32'h00000000} /* (22, 0, 31) {real, imag} */,
  {32'hc644a394, 32'h00000000} /* (22, 0, 30) {real, imag} */,
  {32'hc64d7204, 32'h00000000} /* (22, 0, 29) {real, imag} */,
  {32'hc64e555f, 32'h00000000} /* (22, 0, 28) {real, imag} */,
  {32'hc652d285, 32'h00000000} /* (22, 0, 27) {real, imag} */,
  {32'hc6698270, 32'h00000000} /* (22, 0, 26) {real, imag} */,
  {32'hc64b7124, 32'h00000000} /* (22, 0, 25) {real, imag} */,
  {32'hc62d4905, 32'h00000000} /* (22, 0, 24) {real, imag} */,
  {32'hc6219296, 32'h00000000} /* (22, 0, 23) {real, imag} */,
  {32'hc60eb806, 32'h00000000} /* (22, 0, 22) {real, imag} */,
  {32'hc5c90378, 32'h00000000} /* (22, 0, 21) {real, imag} */,
  {32'hc5b7d8fc, 32'h00000000} /* (22, 0, 20) {real, imag} */,
  {32'hc5486ca1, 32'h00000000} /* (22, 0, 19) {real, imag} */,
  {32'hc4c200b0, 32'h00000000} /* (22, 0, 18) {real, imag} */,
  {32'hc388bdd0, 32'h00000000} /* (22, 0, 17) {real, imag} */,
  {32'h44d00c6c, 32'h00000000} /* (22, 0, 16) {real, imag} */,
  {32'h4568e7c6, 32'h00000000} /* (22, 0, 15) {real, imag} */,
  {32'h45b900a5, 32'h00000000} /* (22, 0, 14) {real, imag} */,
  {32'h45ad5ea0, 32'h00000000} /* (22, 0, 13) {real, imag} */,
  {32'h45b06c86, 32'h00000000} /* (22, 0, 12) {real, imag} */,
  {32'h459edd1a, 32'h00000000} /* (22, 0, 11) {real, imag} */,
  {32'h4541c57e, 32'h00000000} /* (22, 0, 10) {real, imag} */,
  {32'h44edf870, 32'h00000000} /* (22, 0, 9) {real, imag} */,
  {32'h43935380, 32'h00000000} /* (22, 0, 8) {real, imag} */,
  {32'hc4bfa254, 32'h00000000} /* (22, 0, 7) {real, imag} */,
  {32'hc55d3042, 32'h00000000} /* (22, 0, 6) {real, imag} */,
  {32'hc5b59a4c, 32'h00000000} /* (22, 0, 5) {real, imag} */,
  {32'hc5ee1ff0, 32'h00000000} /* (22, 0, 4) {real, imag} */,
  {32'hc6112526, 32'h00000000} /* (22, 0, 3) {real, imag} */,
  {32'hc6238afd, 32'h00000000} /* (22, 0, 2) {real, imag} */,
  {32'hc6380a66, 32'h00000000} /* (22, 0, 1) {real, imag} */,
  {32'hc63d800e, 32'h00000000} /* (22, 0, 0) {real, imag} */,
  {32'hc645522a, 32'h00000000} /* (21, 31, 31) {real, imag} */,
  {32'hc652c6af, 32'h00000000} /* (21, 31, 30) {real, imag} */,
  {32'hc64e8453, 32'h00000000} /* (21, 31, 29) {real, imag} */,
  {32'hc6558b53, 32'h00000000} /* (21, 31, 28) {real, imag} */,
  {32'hc656b350, 32'h00000000} /* (21, 31, 27) {real, imag} */,
  {32'hc64d5753, 32'h00000000} /* (21, 31, 26) {real, imag} */,
  {32'hc649f920, 32'h00000000} /* (21, 31, 25) {real, imag} */,
  {32'hc638d7ff, 32'h00000000} /* (21, 31, 24) {real, imag} */,
  {32'hc61dd8f2, 32'h00000000} /* (21, 31, 23) {real, imag} */,
  {32'hc6029b10, 32'h00000000} /* (21, 31, 22) {real, imag} */,
  {32'hc5c49f7b, 32'h00000000} /* (21, 31, 21) {real, imag} */,
  {32'hc5567576, 32'h00000000} /* (21, 31, 20) {real, imag} */,
  {32'hc481b324, 32'h00000000} /* (21, 31, 19) {real, imag} */,
  {32'h44489298, 32'h00000000} /* (21, 31, 18) {real, imag} */,
  {32'h451f1e26, 32'h00000000} /* (21, 31, 17) {real, imag} */,
  {32'h4588107a, 32'h00000000} /* (21, 31, 16) {real, imag} */,
  {32'h45afad63, 32'h00000000} /* (21, 31, 15) {real, imag} */,
  {32'h45cb5f62, 32'h00000000} /* (21, 31, 14) {real, imag} */,
  {32'h45c74446, 32'h00000000} /* (21, 31, 13) {real, imag} */,
  {32'h45a1aece, 32'h00000000} /* (21, 31, 12) {real, imag} */,
  {32'h4576bf16, 32'h00000000} /* (21, 31, 11) {real, imag} */,
  {32'h44f1d030, 32'h00000000} /* (21, 31, 10) {real, imag} */,
  {32'hc41c48e8, 32'h00000000} /* (21, 31, 9) {real, imag} */,
  {32'hc4ff15e8, 32'h00000000} /* (21, 31, 8) {real, imag} */,
  {32'hc59ab507, 32'h00000000} /* (21, 31, 7) {real, imag} */,
  {32'hc5be303c, 32'h00000000} /* (21, 31, 6) {real, imag} */,
  {32'hc5de32b5, 32'h00000000} /* (21, 31, 5) {real, imag} */,
  {32'hc6052748, 32'h00000000} /* (21, 31, 4) {real, imag} */,
  {32'hc61e536a, 32'h00000000} /* (21, 31, 3) {real, imag} */,
  {32'hc62ef12c, 32'h00000000} /* (21, 31, 2) {real, imag} */,
  {32'hc636ec52, 32'h00000000} /* (21, 31, 1) {real, imag} */,
  {32'hc63aed9a, 32'h00000000} /* (21, 31, 0) {real, imag} */,
  {32'hc64eb626, 32'h00000000} /* (21, 30, 31) {real, imag} */,
  {32'hc6541e26, 32'h00000000} /* (21, 30, 30) {real, imag} */,
  {32'hc653fe2e, 32'h00000000} /* (21, 30, 29) {real, imag} */,
  {32'hc660f0c4, 32'h00000000} /* (21, 30, 28) {real, imag} */,
  {32'hc65ab14c, 32'h00000000} /* (21, 30, 27) {real, imag} */,
  {32'hc64efbaf, 32'h00000000} /* (21, 30, 26) {real, imag} */,
  {32'hc64c596a, 32'h00000000} /* (21, 30, 25) {real, imag} */,
  {32'hc635ff2e, 32'h00000000} /* (21, 30, 24) {real, imag} */,
  {32'hc6229dae, 32'h00000000} /* (21, 30, 23) {real, imag} */,
  {32'hc614a86e, 32'h00000000} /* (21, 30, 22) {real, imag} */,
  {32'hc59bbe5a, 32'h00000000} /* (21, 30, 21) {real, imag} */,
  {32'hc4e4ebde, 32'h00000000} /* (21, 30, 20) {real, imag} */,
  {32'h44e10724, 32'h00000000} /* (21, 30, 19) {real, imag} */,
  {32'h4539b7fa, 32'h00000000} /* (21, 30, 18) {real, imag} */,
  {32'h4567b47a, 32'h00000000} /* (21, 30, 17) {real, imag} */,
  {32'h45b2ddac, 32'h00000000} /* (21, 30, 16) {real, imag} */,
  {32'h45d656e4, 32'h00000000} /* (21, 30, 15) {real, imag} */,
  {32'h45fc2077, 32'h00000000} /* (21, 30, 14) {real, imag} */,
  {32'h45f04c73, 32'h00000000} /* (21, 30, 13) {real, imag} */,
  {32'h45b1372d, 32'h00000000} /* (21, 30, 12) {real, imag} */,
  {32'h457003b6, 32'h00000000} /* (21, 30, 11) {real, imag} */,
  {32'h447bbc90, 32'h00000000} /* (21, 30, 10) {real, imag} */,
  {32'hc50bf292, 32'h00000000} /* (21, 30, 9) {real, imag} */,
  {32'hc57c185e, 32'h00000000} /* (21, 30, 8) {real, imag} */,
  {32'hc5b46c01, 32'h00000000} /* (21, 30, 7) {real, imag} */,
  {32'hc5f60c2b, 32'h00000000} /* (21, 30, 6) {real, imag} */,
  {32'hc607d7a4, 32'h00000000} /* (21, 30, 5) {real, imag} */,
  {32'hc612d4c7, 32'h00000000} /* (21, 30, 4) {real, imag} */,
  {32'hc6249e2c, 32'h00000000} /* (21, 30, 3) {real, imag} */,
  {32'hc63e89dc, 32'h00000000} /* (21, 30, 2) {real, imag} */,
  {32'hc64fec12, 32'h00000000} /* (21, 30, 1) {real, imag} */,
  {32'hc6433e9c, 32'h00000000} /* (21, 30, 0) {real, imag} */,
  {32'hc65a0d24, 32'h00000000} /* (21, 29, 31) {real, imag} */,
  {32'hc66a8710, 32'h00000000} /* (21, 29, 30) {real, imag} */,
  {32'hc65665c3, 32'h00000000} /* (21, 29, 29) {real, imag} */,
  {32'hc65f0302, 32'h00000000} /* (21, 29, 28) {real, imag} */,
  {32'hc659efe2, 32'h00000000} /* (21, 29, 27) {real, imag} */,
  {32'hc65004dd, 32'h00000000} /* (21, 29, 26) {real, imag} */,
  {32'hc654db3a, 32'h00000000} /* (21, 29, 25) {real, imag} */,
  {32'hc63a8852, 32'h00000000} /* (21, 29, 24) {real, imag} */,
  {32'hc6253710, 32'h00000000} /* (21, 29, 23) {real, imag} */,
  {32'hc5fb93f6, 32'h00000000} /* (21, 29, 22) {real, imag} */,
  {32'hc57a7ee5, 32'h00000000} /* (21, 29, 21) {real, imag} */,
  {32'h440797d8, 32'h00000000} /* (21, 29, 20) {real, imag} */,
  {32'h4546d146, 32'h00000000} /* (21, 29, 19) {real, imag} */,
  {32'h45bc98df, 32'h00000000} /* (21, 29, 18) {real, imag} */,
  {32'h45c324b0, 32'h00000000} /* (21, 29, 17) {real, imag} */,
  {32'h45dedb0a, 32'h00000000} /* (21, 29, 16) {real, imag} */,
  {32'h45ef7f54, 32'h00000000} /* (21, 29, 15) {real, imag} */,
  {32'h45e80020, 32'h00000000} /* (21, 29, 14) {real, imag} */,
  {32'h45e54ece, 32'h00000000} /* (21, 29, 13) {real, imag} */,
  {32'h45c2e4d7, 32'h00000000} /* (21, 29, 12) {real, imag} */,
  {32'h454c2460, 32'h00000000} /* (21, 29, 11) {real, imag} */,
  {32'hc248c800, 32'h00000000} /* (21, 29, 10) {real, imag} */,
  {32'hc569cef8, 32'h00000000} /* (21, 29, 9) {real, imag} */,
  {32'hc5b6b19c, 32'h00000000} /* (21, 29, 8) {real, imag} */,
  {32'hc5e05838, 32'h00000000} /* (21, 29, 7) {real, imag} */,
  {32'hc60726db, 32'h00000000} /* (21, 29, 6) {real, imag} */,
  {32'hc619f7cf, 32'h00000000} /* (21, 29, 5) {real, imag} */,
  {32'hc62b5a50, 32'h00000000} /* (21, 29, 4) {real, imag} */,
  {32'hc636889a, 32'h00000000} /* (21, 29, 3) {real, imag} */,
  {32'hc644406c, 32'h00000000} /* (21, 29, 2) {real, imag} */,
  {32'hc651134c, 32'h00000000} /* (21, 29, 1) {real, imag} */,
  {32'hc642e85b, 32'h00000000} /* (21, 29, 0) {real, imag} */,
  {32'hc64af82c, 32'h00000000} /* (21, 28, 31) {real, imag} */,
  {32'hc65d952b, 32'h00000000} /* (21, 28, 30) {real, imag} */,
  {32'hc6557442, 32'h00000000} /* (21, 28, 29) {real, imag} */,
  {32'hc6631a50, 32'h00000000} /* (21, 28, 28) {real, imag} */,
  {32'hc6665428, 32'h00000000} /* (21, 28, 27) {real, imag} */,
  {32'hc64e644a, 32'h00000000} /* (21, 28, 26) {real, imag} */,
  {32'hc65721e3, 32'h00000000} /* (21, 28, 25) {real, imag} */,
  {32'hc6393e78, 32'h00000000} /* (21, 28, 24) {real, imag} */,
  {32'hc62ab6ac, 32'h00000000} /* (21, 28, 23) {real, imag} */,
  {32'hc6024d7e, 32'h00000000} /* (21, 28, 22) {real, imag} */,
  {32'hc597bca6, 32'h00000000} /* (21, 28, 21) {real, imag} */,
  {32'hc3771ee0, 32'h00000000} /* (21, 28, 20) {real, imag} */,
  {32'h4573e910, 32'h00000000} /* (21, 28, 19) {real, imag} */,
  {32'h45bbc83a, 32'h00000000} /* (21, 28, 18) {real, imag} */,
  {32'h45deef3e, 32'h00000000} /* (21, 28, 17) {real, imag} */,
  {32'h45fb77a6, 32'h00000000} /* (21, 28, 16) {real, imag} */,
  {32'h46015ff4, 32'h00000000} /* (21, 28, 15) {real, imag} */,
  {32'h46016d09, 32'h00000000} /* (21, 28, 14) {real, imag} */,
  {32'h45ce9300, 32'h00000000} /* (21, 28, 13) {real, imag} */,
  {32'h45c93c24, 32'h00000000} /* (21, 28, 12) {real, imag} */,
  {32'h455424f8, 32'h00000000} /* (21, 28, 11) {real, imag} */,
  {32'hc48ca54c, 32'h00000000} /* (21, 28, 10) {real, imag} */,
  {32'hc5b1330a, 32'h00000000} /* (21, 28, 9) {real, imag} */,
  {32'hc5dba4cd, 32'h00000000} /* (21, 28, 8) {real, imag} */,
  {32'hc610b960, 32'h00000000} /* (21, 28, 7) {real, imag} */,
  {32'hc6219514, 32'h00000000} /* (21, 28, 6) {real, imag} */,
  {32'hc62ede91, 32'h00000000} /* (21, 28, 5) {real, imag} */,
  {32'hc6418b04, 32'h00000000} /* (21, 28, 4) {real, imag} */,
  {32'hc6499bfc, 32'h00000000} /* (21, 28, 3) {real, imag} */,
  {32'hc6422bb5, 32'h00000000} /* (21, 28, 2) {real, imag} */,
  {32'hc64fb849, 32'h00000000} /* (21, 28, 1) {real, imag} */,
  {32'hc6590d07, 32'h00000000} /* (21, 28, 0) {real, imag} */,
  {32'hc64a8f92, 32'h00000000} /* (21, 27, 31) {real, imag} */,
  {32'hc64a6ae3, 32'h00000000} /* (21, 27, 30) {real, imag} */,
  {32'hc65992b8, 32'h00000000} /* (21, 27, 29) {real, imag} */,
  {32'hc665f15e, 32'h00000000} /* (21, 27, 28) {real, imag} */,
  {32'hc6613693, 32'h00000000} /* (21, 27, 27) {real, imag} */,
  {32'hc657b018, 32'h00000000} /* (21, 27, 26) {real, imag} */,
  {32'hc642bb1c, 32'h00000000} /* (21, 27, 25) {real, imag} */,
  {32'hc63e910a, 32'h00000000} /* (21, 27, 24) {real, imag} */,
  {32'hc628f8aa, 32'h00000000} /* (21, 27, 23) {real, imag} */,
  {32'hc6078f64, 32'h00000000} /* (21, 27, 22) {real, imag} */,
  {32'hc57d7874, 32'h00000000} /* (21, 27, 21) {real, imag} */,
  {32'hc26b4400, 32'h00000000} /* (21, 27, 20) {real, imag} */,
  {32'h453ac044, 32'h00000000} /* (21, 27, 19) {real, imag} */,
  {32'h45aeae18, 32'h00000000} /* (21, 27, 18) {real, imag} */,
  {32'h45d9dace, 32'h00000000} /* (21, 27, 17) {real, imag} */,
  {32'h45e70eec, 32'h00000000} /* (21, 27, 16) {real, imag} */,
  {32'h4609852e, 32'h00000000} /* (21, 27, 15) {real, imag} */,
  {32'h45ffd66a, 32'h00000000} /* (21, 27, 14) {real, imag} */,
  {32'h45d78bcf, 32'h00000000} /* (21, 27, 13) {real, imag} */,
  {32'h45a393ac, 32'h00000000} /* (21, 27, 12) {real, imag} */,
  {32'h452241a4, 32'h00000000} /* (21, 27, 11) {real, imag} */,
  {32'hc4f1c310, 32'h00000000} /* (21, 27, 10) {real, imag} */,
  {32'hc59dd764, 32'h00000000} /* (21, 27, 9) {real, imag} */,
  {32'hc6050946, 32'h00000000} /* (21, 27, 8) {real, imag} */,
  {32'hc6130982, 32'h00000000} /* (21, 27, 7) {real, imag} */,
  {32'hc633128c, 32'h00000000} /* (21, 27, 6) {real, imag} */,
  {32'hc63bd8fc, 32'h00000000} /* (21, 27, 5) {real, imag} */,
  {32'hc63f3da2, 32'h00000000} /* (21, 27, 4) {real, imag} */,
  {32'hc642d34d, 32'h00000000} /* (21, 27, 3) {real, imag} */,
  {32'hc65be5d0, 32'h00000000} /* (21, 27, 2) {real, imag} */,
  {32'hc653193b, 32'h00000000} /* (21, 27, 1) {real, imag} */,
  {32'hc6500cac, 32'h00000000} /* (21, 27, 0) {real, imag} */,
  {32'hc6379c23, 32'h00000000} /* (21, 26, 31) {real, imag} */,
  {32'hc655794e, 32'h00000000} /* (21, 26, 30) {real, imag} */,
  {32'hc64d3a10, 32'h00000000} /* (21, 26, 29) {real, imag} */,
  {32'hc646380a, 32'h00000000} /* (21, 26, 28) {real, imag} */,
  {32'hc6620ca9, 32'h00000000} /* (21, 26, 27) {real, imag} */,
  {32'hc64b78b8, 32'h00000000} /* (21, 26, 26) {real, imag} */,
  {32'hc63c7b52, 32'h00000000} /* (21, 26, 25) {real, imag} */,
  {32'hc64f6506, 32'h00000000} /* (21, 26, 24) {real, imag} */,
  {32'hc61e064d, 32'h00000000} /* (21, 26, 23) {real, imag} */,
  {32'hc5d087cf, 32'h00000000} /* (21, 26, 22) {real, imag} */,
  {32'hc5743b59, 32'h00000000} /* (21, 26, 21) {real, imag} */,
  {32'h4326dac0, 32'h00000000} /* (21, 26, 20) {real, imag} */,
  {32'h4581c352, 32'h00000000} /* (21, 26, 19) {real, imag} */,
  {32'h45b3ac01, 32'h00000000} /* (21, 26, 18) {real, imag} */,
  {32'h45e52e4c, 32'h00000000} /* (21, 26, 17) {real, imag} */,
  {32'h45fff3f5, 32'h00000000} /* (21, 26, 16) {real, imag} */,
  {32'h45f38942, 32'h00000000} /* (21, 26, 15) {real, imag} */,
  {32'h45f3cf1c, 32'h00000000} /* (21, 26, 14) {real, imag} */,
  {32'h45ec8684, 32'h00000000} /* (21, 26, 13) {real, imag} */,
  {32'h45ae6cf8, 32'h00000000} /* (21, 26, 12) {real, imag} */,
  {32'h4502314c, 32'h00000000} /* (21, 26, 11) {real, imag} */,
  {32'hc530b6fe, 32'h00000000} /* (21, 26, 10) {real, imag} */,
  {32'hc5ce3d01, 32'h00000000} /* (21, 26, 9) {real, imag} */,
  {32'hc5fc78eb, 32'h00000000} /* (21, 26, 8) {real, imag} */,
  {32'hc61bf6ff, 32'h00000000} /* (21, 26, 7) {real, imag} */,
  {32'hc62ae09a, 32'h00000000} /* (21, 26, 6) {real, imag} */,
  {32'hc62bfc1c, 32'h00000000} /* (21, 26, 5) {real, imag} */,
  {32'hc639a18b, 32'h00000000} /* (21, 26, 4) {real, imag} */,
  {32'hc6449ee5, 32'h00000000} /* (21, 26, 3) {real, imag} */,
  {32'hc645ab84, 32'h00000000} /* (21, 26, 2) {real, imag} */,
  {32'hc64d8fbc, 32'h00000000} /* (21, 26, 1) {real, imag} */,
  {32'hc63f1ffe, 32'h00000000} /* (21, 26, 0) {real, imag} */,
  {32'hc63068f8, 32'h00000000} /* (21, 25, 31) {real, imag} */,
  {32'hc631182f, 32'h00000000} /* (21, 25, 30) {real, imag} */,
  {32'hc63b4fae, 32'h00000000} /* (21, 25, 29) {real, imag} */,
  {32'hc6410920, 32'h00000000} /* (21, 25, 28) {real, imag} */,
  {32'hc64cec8e, 32'h00000000} /* (21, 25, 27) {real, imag} */,
  {32'hc643ffba, 32'h00000000} /* (21, 25, 26) {real, imag} */,
  {32'hc62eac0d, 32'h00000000} /* (21, 25, 25) {real, imag} */,
  {32'hc626b71a, 32'h00000000} /* (21, 25, 24) {real, imag} */,
  {32'hc6043172, 32'h00000000} /* (21, 25, 23) {real, imag} */,
  {32'hc5da383a, 32'h00000000} /* (21, 25, 22) {real, imag} */,
  {32'hc575bf92, 32'h00000000} /* (21, 25, 21) {real, imag} */,
  {32'h43b14a80, 32'h00000000} /* (21, 25, 20) {real, imag} */,
  {32'h4581f19a, 32'h00000000} /* (21, 25, 19) {real, imag} */,
  {32'h45c6d15e, 32'h00000000} /* (21, 25, 18) {real, imag} */,
  {32'h45de8554, 32'h00000000} /* (21, 25, 17) {real, imag} */,
  {32'h45f47d36, 32'h00000000} /* (21, 25, 16) {real, imag} */,
  {32'h460455b6, 32'h00000000} /* (21, 25, 15) {real, imag} */,
  {32'h46050713, 32'h00000000} /* (21, 25, 14) {real, imag} */,
  {32'h45cb125d, 32'h00000000} /* (21, 25, 13) {real, imag} */,
  {32'h459ea7a0, 32'h00000000} /* (21, 25, 12) {real, imag} */,
  {32'h44f78528, 32'h00000000} /* (21, 25, 11) {real, imag} */,
  {32'hc53aa5f8, 32'h00000000} /* (21, 25, 10) {real, imag} */,
  {32'hc5c85472, 32'h00000000} /* (21, 25, 9) {real, imag} */,
  {32'hc5f711e4, 32'h00000000} /* (21, 25, 8) {real, imag} */,
  {32'hc60e38fa, 32'h00000000} /* (21, 25, 7) {real, imag} */,
  {32'hc61609e5, 32'h00000000} /* (21, 25, 6) {real, imag} */,
  {32'hc62a1d2c, 32'h00000000} /* (21, 25, 5) {real, imag} */,
  {32'hc631b02a, 32'h00000000} /* (21, 25, 4) {real, imag} */,
  {32'hc6399ea8, 32'h00000000} /* (21, 25, 3) {real, imag} */,
  {32'hc6456da1, 32'h00000000} /* (21, 25, 2) {real, imag} */,
  {32'hc632e7c0, 32'h00000000} /* (21, 25, 1) {real, imag} */,
  {32'hc62fdf91, 32'h00000000} /* (21, 25, 0) {real, imag} */,
  {32'hc613672b, 32'h00000000} /* (21, 24, 31) {real, imag} */,
  {32'hc6159d08, 32'h00000000} /* (21, 24, 30) {real, imag} */,
  {32'hc6197119, 32'h00000000} /* (21, 24, 29) {real, imag} */,
  {32'hc61e146c, 32'h00000000} /* (21, 24, 28) {real, imag} */,
  {32'hc61bdf04, 32'h00000000} /* (21, 24, 27) {real, imag} */,
  {32'hc61eb4bc, 32'h00000000} /* (21, 24, 26) {real, imag} */,
  {32'hc604f602, 32'h00000000} /* (21, 24, 25) {real, imag} */,
  {32'hc60b8c63, 32'h00000000} /* (21, 24, 24) {real, imag} */,
  {32'hc5f10d70, 32'h00000000} /* (21, 24, 23) {real, imag} */,
  {32'hc5c03db9, 32'h00000000} /* (21, 24, 22) {real, imag} */,
  {32'hc54114f4, 32'h00000000} /* (21, 24, 21) {real, imag} */,
  {32'h446aed10, 32'h00000000} /* (21, 24, 20) {real, imag} */,
  {32'h458f63a8, 32'h00000000} /* (21, 24, 19) {real, imag} */,
  {32'h45d15da9, 32'h00000000} /* (21, 24, 18) {real, imag} */,
  {32'h45aece4d, 32'h00000000} /* (21, 24, 17) {real, imag} */,
  {32'h45f1071f, 32'h00000000} /* (21, 24, 16) {real, imag} */,
  {32'h45efc6e2, 32'h00000000} /* (21, 24, 15) {real, imag} */,
  {32'h45d68841, 32'h00000000} /* (21, 24, 14) {real, imag} */,
  {32'h45bbac48, 32'h00000000} /* (21, 24, 13) {real, imag} */,
  {32'h45908e6e, 32'h00000000} /* (21, 24, 12) {real, imag} */,
  {32'h45027002, 32'h00000000} /* (21, 24, 11) {real, imag} */,
  {32'hc4fbf178, 32'h00000000} /* (21, 24, 10) {real, imag} */,
  {32'hc5a51749, 32'h00000000} /* (21, 24, 9) {real, imag} */,
  {32'hc5d0310d, 32'h00000000} /* (21, 24, 8) {real, imag} */,
  {32'hc60392f6, 32'h00000000} /* (21, 24, 7) {real, imag} */,
  {32'hc6189812, 32'h00000000} /* (21, 24, 6) {real, imag} */,
  {32'hc61677fc, 32'h00000000} /* (21, 24, 5) {real, imag} */,
  {32'hc619fb49, 32'h00000000} /* (21, 24, 4) {real, imag} */,
  {32'hc6206b8f, 32'h00000000} /* (21, 24, 3) {real, imag} */,
  {32'hc62ba73c, 32'h00000000} /* (21, 24, 2) {real, imag} */,
  {32'hc6240cda, 32'h00000000} /* (21, 24, 1) {real, imag} */,
  {32'hc610b2e2, 32'h00000000} /* (21, 24, 0) {real, imag} */,
  {32'hc5e8af94, 32'h00000000} /* (21, 23, 31) {real, imag} */,
  {32'hc60631bc, 32'h00000000} /* (21, 23, 30) {real, imag} */,
  {32'hc60cc966, 32'h00000000} /* (21, 23, 29) {real, imag} */,
  {32'hc605b7aa, 32'h00000000} /* (21, 23, 28) {real, imag} */,
  {32'hc5f716b4, 32'h00000000} /* (21, 23, 27) {real, imag} */,
  {32'hc5fa7aaa, 32'h00000000} /* (21, 23, 26) {real, imag} */,
  {32'hc5e37b7d, 32'h00000000} /* (21, 23, 25) {real, imag} */,
  {32'hc5db1316, 32'h00000000} /* (21, 23, 24) {real, imag} */,
  {32'hc5ccf326, 32'h00000000} /* (21, 23, 23) {real, imag} */,
  {32'hc59c3c17, 32'h00000000} /* (21, 23, 22) {real, imag} */,
  {32'hc51c84cd, 32'h00000000} /* (21, 23, 21) {real, imag} */,
  {32'h44d3b734, 32'h00000000} /* (21, 23, 20) {real, imag} */,
  {32'h45252509, 32'h00000000} /* (21, 23, 19) {real, imag} */,
  {32'h45853ffb, 32'h00000000} /* (21, 23, 18) {real, imag} */,
  {32'h459f949c, 32'h00000000} /* (21, 23, 17) {real, imag} */,
  {32'h45c5c6b8, 32'h00000000} /* (21, 23, 16) {real, imag} */,
  {32'h45b6971e, 32'h00000000} /* (21, 23, 15) {real, imag} */,
  {32'h459dd2c0, 32'h00000000} /* (21, 23, 14) {real, imag} */,
  {32'h4597b971, 32'h00000000} /* (21, 23, 13) {real, imag} */,
  {32'h456b7ede, 32'h00000000} /* (21, 23, 12) {real, imag} */,
  {32'h44990a02, 32'h00000000} /* (21, 23, 11) {real, imag} */,
  {32'hc50e6c75, 32'h00000000} /* (21, 23, 10) {real, imag} */,
  {32'hc5828eef, 32'h00000000} /* (21, 23, 9) {real, imag} */,
  {32'hc5a85172, 32'h00000000} /* (21, 23, 8) {real, imag} */,
  {32'hc5e19bb6, 32'h00000000} /* (21, 23, 7) {real, imag} */,
  {32'hc5e7d1c1, 32'h00000000} /* (21, 23, 6) {real, imag} */,
  {32'hc608f0f4, 32'h00000000} /* (21, 23, 5) {real, imag} */,
  {32'hc60c0b42, 32'h00000000} /* (21, 23, 4) {real, imag} */,
  {32'hc60b64cf, 32'h00000000} /* (21, 23, 3) {real, imag} */,
  {32'hc6009c22, 32'h00000000} /* (21, 23, 2) {real, imag} */,
  {32'hc603ec43, 32'h00000000} /* (21, 23, 1) {real, imag} */,
  {32'hc5f711d6, 32'h00000000} /* (21, 23, 0) {real, imag} */,
  {32'hc5aa167b, 32'h00000000} /* (21, 22, 31) {real, imag} */,
  {32'hc5c34205, 32'h00000000} /* (21, 22, 30) {real, imag} */,
  {32'hc5ba52c4, 32'h00000000} /* (21, 22, 29) {real, imag} */,
  {32'hc5b5cd4c, 32'h00000000} /* (21, 22, 28) {real, imag} */,
  {32'hc5af7e4e, 32'h00000000} /* (21, 22, 27) {real, imag} */,
  {32'hc59887db, 32'h00000000} /* (21, 22, 26) {real, imag} */,
  {32'hc5882c66, 32'h00000000} /* (21, 22, 25) {real, imag} */,
  {32'hc5953bb1, 32'h00000000} /* (21, 22, 24) {real, imag} */,
  {32'hc5937ecd, 32'h00000000} /* (21, 22, 23) {real, imag} */,
  {32'hc5527ba0, 32'h00000000} /* (21, 22, 22) {real, imag} */,
  {32'hc4f540b4, 32'h00000000} /* (21, 22, 21) {real, imag} */,
  {32'h44ab1884, 32'h00000000} /* (21, 22, 20) {real, imag} */,
  {32'h4506c51c, 32'h00000000} /* (21, 22, 19) {real, imag} */,
  {32'h454b2dde, 32'h00000000} /* (21, 22, 18) {real, imag} */,
  {32'h4533bab8, 32'h00000000} /* (21, 22, 17) {real, imag} */,
  {32'h457a8fd8, 32'h00000000} /* (21, 22, 16) {real, imag} */,
  {32'h4585c4a3, 32'h00000000} /* (21, 22, 15) {real, imag} */,
  {32'h455c4ce6, 32'h00000000} /* (21, 22, 14) {real, imag} */,
  {32'h4580372a, 32'h00000000} /* (21, 22, 13) {real, imag} */,
  {32'h45327288, 32'h00000000} /* (21, 22, 12) {real, imag} */,
  {32'h441d1a64, 32'h00000000} /* (21, 22, 11) {real, imag} */,
  {32'hc4d0422b, 32'h00000000} /* (21, 22, 10) {real, imag} */,
  {32'hc515d7a8, 32'h00000000} /* (21, 22, 9) {real, imag} */,
  {32'hc589ea59, 32'h00000000} /* (21, 22, 8) {real, imag} */,
  {32'hc59fe0d9, 32'h00000000} /* (21, 22, 7) {real, imag} */,
  {32'hc5a9466e, 32'h00000000} /* (21, 22, 6) {real, imag} */,
  {32'hc5b98008, 32'h00000000} /* (21, 22, 5) {real, imag} */,
  {32'hc5d3612b, 32'h00000000} /* (21, 22, 4) {real, imag} */,
  {32'hc5e45672, 32'h00000000} /* (21, 22, 3) {real, imag} */,
  {32'hc5c12151, 32'h00000000} /* (21, 22, 2) {real, imag} */,
  {32'hc5d40d56, 32'h00000000} /* (21, 22, 1) {real, imag} */,
  {32'hc5b22ca0, 32'h00000000} /* (21, 22, 0) {real, imag} */,
  {32'hc50ed98c, 32'h00000000} /* (21, 21, 31) {real, imag} */,
  {32'hc4fe1ad0, 32'h00000000} /* (21, 21, 30) {real, imag} */,
  {32'hc4e743f2, 32'h00000000} /* (21, 21, 29) {real, imag} */,
  {32'hc4da67ef, 32'h00000000} /* (21, 21, 28) {real, imag} */,
  {32'hc4c22b60, 32'h00000000} /* (21, 21, 27) {real, imag} */,
  {32'hc4e8a488, 32'h00000000} /* (21, 21, 26) {real, imag} */,
  {32'hc4b32601, 32'h00000000} /* (21, 21, 25) {real, imag} */,
  {32'hc49a0bb8, 32'h00000000} /* (21, 21, 24) {real, imag} */,
  {32'hc4b05043, 32'h00000000} /* (21, 21, 23) {real, imag} */,
  {32'hc492980c, 32'h00000000} /* (21, 21, 22) {real, imag} */,
  {32'hc428922c, 32'h00000000} /* (21, 21, 21) {real, imag} */,
  {32'hc401ca0f, 32'h00000000} /* (21, 21, 20) {real, imag} */,
  {32'h43db8850, 32'h00000000} /* (21, 21, 19) {real, imag} */,
  {32'h43c93d1e, 32'h00000000} /* (21, 21, 18) {real, imag} */,
  {32'hc1d96b40, 32'h00000000} /* (21, 21, 17) {real, imag} */,
  {32'h43948208, 32'h00000000} /* (21, 21, 16) {real, imag} */,
  {32'h449ab1d5, 32'h00000000} /* (21, 21, 15) {real, imag} */,
  {32'h446100ac, 32'h00000000} /* (21, 21, 14) {real, imag} */,
  {32'h44b3a8c4, 32'h00000000} /* (21, 21, 13) {real, imag} */,
  {32'h446448aa, 32'h00000000} /* (21, 21, 12) {real, imag} */,
  {32'h43f790b0, 32'h00000000} /* (21, 21, 11) {real, imag} */,
  {32'hc495d19c, 32'h00000000} /* (21, 21, 10) {real, imag} */,
  {32'hc479d7de, 32'h00000000} /* (21, 21, 9) {real, imag} */,
  {32'hc4c1e438, 32'h00000000} /* (21, 21, 8) {real, imag} */,
  {32'hc4f13c1b, 32'h00000000} /* (21, 21, 7) {real, imag} */,
  {32'hc4e78e16, 32'h00000000} /* (21, 21, 6) {real, imag} */,
  {32'hc5029d3b, 32'h00000000} /* (21, 21, 5) {real, imag} */,
  {32'hc4fb6746, 32'h00000000} /* (21, 21, 4) {real, imag} */,
  {32'hc520ccea, 32'h00000000} /* (21, 21, 3) {real, imag} */,
  {32'hc506e944, 32'h00000000} /* (21, 21, 2) {real, imag} */,
  {32'hc563cd28, 32'h00000000} /* (21, 21, 1) {real, imag} */,
  {32'hc525fb45, 32'h00000000} /* (21, 21, 0) {real, imag} */,
  {32'h44908943, 32'h00000000} /* (21, 20, 31) {real, imag} */,
  {32'h44c8c630, 32'h00000000} /* (21, 20, 30) {real, imag} */,
  {32'h452180a6, 32'h00000000} /* (21, 20, 29) {real, imag} */,
  {32'h44f5307b, 32'h00000000} /* (21, 20, 28) {real, imag} */,
  {32'h453393bd, 32'h00000000} /* (21, 20, 27) {real, imag} */,
  {32'h44ea440e, 32'h00000000} /* (21, 20, 26) {real, imag} */,
  {32'h45199333, 32'h00000000} /* (21, 20, 25) {real, imag} */,
  {32'h45279267, 32'h00000000} /* (21, 20, 24) {real, imag} */,
  {32'h449d2a7a, 32'h00000000} /* (21, 20, 23) {real, imag} */,
  {32'h446836bd, 32'h00000000} /* (21, 20, 22) {real, imag} */,
  {32'hc34cac40, 32'h00000000} /* (21, 20, 21) {real, imag} */,
  {32'hc4a840b1, 32'h00000000} /* (21, 20, 20) {real, imag} */,
  {32'hc504b38d, 32'h00000000} /* (21, 20, 19) {real, imag} */,
  {32'hc529713c, 32'h00000000} /* (21, 20, 18) {real, imag} */,
  {32'hc59c2c70, 32'h00000000} /* (21, 20, 17) {real, imag} */,
  {32'hc54e3784, 32'h00000000} /* (21, 20, 16) {real, imag} */,
  {32'hc51cb836, 32'h00000000} /* (21, 20, 15) {real, imag} */,
  {32'hc516039c, 32'h00000000} /* (21, 20, 14) {real, imag} */,
  {32'hc52eac44, 32'h00000000} /* (21, 20, 13) {real, imag} */,
  {32'hc499436d, 32'h00000000} /* (21, 20, 12) {real, imag} */,
  {32'hc4f8222e, 32'h00000000} /* (21, 20, 11) {real, imag} */,
  {32'hc447bd3c, 32'h00000000} /* (21, 20, 10) {real, imag} */,
  {32'h449156a6, 32'h00000000} /* (21, 20, 9) {real, imag} */,
  {32'h4461407c, 32'h00000000} /* (21, 20, 8) {real, imag} */,
  {32'h4471e86b, 32'h00000000} /* (21, 20, 7) {real, imag} */,
  {32'h44e5f00e, 32'h00000000} /* (21, 20, 6) {real, imag} */,
  {32'h44fab8fa, 32'h00000000} /* (21, 20, 5) {real, imag} */,
  {32'h453d22b6, 32'h00000000} /* (21, 20, 4) {real, imag} */,
  {32'h4528dbe3, 32'h00000000} /* (21, 20, 3) {real, imag} */,
  {32'h44e505ff, 32'h00000000} /* (21, 20, 2) {real, imag} */,
  {32'h44804232, 32'h00000000} /* (21, 20, 1) {real, imag} */,
  {32'h446d1788, 32'h00000000} /* (21, 20, 0) {real, imag} */,
  {32'h4585b6c6, 32'h00000000} /* (21, 19, 31) {real, imag} */,
  {32'h45993137, 32'h00000000} /* (21, 19, 30) {real, imag} */,
  {32'h45b31e20, 32'h00000000} /* (21, 19, 29) {real, imag} */,
  {32'h45adbb36, 32'h00000000} /* (21, 19, 28) {real, imag} */,
  {32'h459affb4, 32'h00000000} /* (21, 19, 27) {real, imag} */,
  {32'h45a77988, 32'h00000000} /* (21, 19, 26) {real, imag} */,
  {32'h45937f49, 32'h00000000} /* (21, 19, 25) {real, imag} */,
  {32'h4595cfb5, 32'h00000000} /* (21, 19, 24) {real, imag} */,
  {32'h456f045e, 32'h00000000} /* (21, 19, 23) {real, imag} */,
  {32'h4505bf6a, 32'h00000000} /* (21, 19, 22) {real, imag} */,
  {32'h44212360, 32'h00000000} /* (21, 19, 21) {real, imag} */,
  {32'hc5193f8e, 32'h00000000} /* (21, 19, 20) {real, imag} */,
  {32'hc54f1841, 32'h00000000} /* (21, 19, 19) {real, imag} */,
  {32'hc59447e4, 32'h00000000} /* (21, 19, 18) {real, imag} */,
  {32'hc5c3ee03, 32'h00000000} /* (21, 19, 17) {real, imag} */,
  {32'hc5bbb44a, 32'h00000000} /* (21, 19, 16) {real, imag} */,
  {32'hc5b90270, 32'h00000000} /* (21, 19, 15) {real, imag} */,
  {32'hc5ab3e07, 32'h00000000} /* (21, 19, 14) {real, imag} */,
  {32'hc5a19b2c, 32'h00000000} /* (21, 19, 13) {real, imag} */,
  {32'hc587d416, 32'h00000000} /* (21, 19, 12) {real, imag} */,
  {32'hc5183208, 32'h00000000} /* (21, 19, 11) {real, imag} */,
  {32'hc2dd22a0, 32'h00000000} /* (21, 19, 10) {real, imag} */,
  {32'h44c2ecdc, 32'h00000000} /* (21, 19, 9) {real, imag} */,
  {32'h452187f6, 32'h00000000} /* (21, 19, 8) {real, imag} */,
  {32'h4537012e, 32'h00000000} /* (21, 19, 7) {real, imag} */,
  {32'h4591db02, 32'h00000000} /* (21, 19, 6) {real, imag} */,
  {32'h458ddc50, 32'h00000000} /* (21, 19, 5) {real, imag} */,
  {32'h457b2116, 32'h00000000} /* (21, 19, 4) {real, imag} */,
  {32'h459ec6df, 32'h00000000} /* (21, 19, 3) {real, imag} */,
  {32'h45bdfcd0, 32'h00000000} /* (21, 19, 2) {real, imag} */,
  {32'h45864ccf, 32'h00000000} /* (21, 19, 1) {real, imag} */,
  {32'h456ccb84, 32'h00000000} /* (21, 19, 0) {real, imag} */,
  {32'h45d3cc01, 32'h00000000} /* (21, 18, 31) {real, imag} */,
  {32'h45cce43c, 32'h00000000} /* (21, 18, 30) {real, imag} */,
  {32'h45f26268, 32'h00000000} /* (21, 18, 29) {real, imag} */,
  {32'h45f204ea, 32'h00000000} /* (21, 18, 28) {real, imag} */,
  {32'h45e4c89e, 32'h00000000} /* (21, 18, 27) {real, imag} */,
  {32'h45d8dd03, 32'h00000000} /* (21, 18, 26) {real, imag} */,
  {32'h45e34b2f, 32'h00000000} /* (21, 18, 25) {real, imag} */,
  {32'h45bfd9cc, 32'h00000000} /* (21, 18, 24) {real, imag} */,
  {32'h45b0d3c2, 32'h00000000} /* (21, 18, 23) {real, imag} */,
  {32'h454e4680, 32'h00000000} /* (21, 18, 22) {real, imag} */,
  {32'hc3f69c48, 32'h00000000} /* (21, 18, 21) {real, imag} */,
  {32'hc4c3325c, 32'h00000000} /* (21, 18, 20) {real, imag} */,
  {32'hc585cbf6, 32'h00000000} /* (21, 18, 19) {real, imag} */,
  {32'hc5db120a, 32'h00000000} /* (21, 18, 18) {real, imag} */,
  {32'hc5db70f3, 32'h00000000} /* (21, 18, 17) {real, imag} */,
  {32'hc5f31fd4, 32'h00000000} /* (21, 18, 16) {real, imag} */,
  {32'hc5f98469, 32'h00000000} /* (21, 18, 15) {real, imag} */,
  {32'hc5bc2a9c, 32'h00000000} /* (21, 18, 14) {real, imag} */,
  {32'hc5afda12, 32'h00000000} /* (21, 18, 13) {real, imag} */,
  {32'hc593eb4c, 32'h00000000} /* (21, 18, 12) {real, imag} */,
  {32'hc51071a4, 32'h00000000} /* (21, 18, 11) {real, imag} */,
  {32'hc373a080, 32'h00000000} /* (21, 18, 10) {real, imag} */,
  {32'h45078e96, 32'h00000000} /* (21, 18, 9) {real, imag} */,
  {32'h458d4f60, 32'h00000000} /* (21, 18, 8) {real, imag} */,
  {32'h45ae19f8, 32'h00000000} /* (21, 18, 7) {real, imag} */,
  {32'h45cb7114, 32'h00000000} /* (21, 18, 6) {real, imag} */,
  {32'h45dbf434, 32'h00000000} /* (21, 18, 5) {real, imag} */,
  {32'h45d3a57d, 32'h00000000} /* (21, 18, 4) {real, imag} */,
  {32'h45d61a28, 32'h00000000} /* (21, 18, 3) {real, imag} */,
  {32'h45ee6f26, 32'h00000000} /* (21, 18, 2) {real, imag} */,
  {32'h45ec6273, 32'h00000000} /* (21, 18, 1) {real, imag} */,
  {32'h45c39c04, 32'h00000000} /* (21, 18, 0) {real, imag} */,
  {32'h45e36a90, 32'h00000000} /* (21, 17, 31) {real, imag} */,
  {32'h45f68c9a, 32'h00000000} /* (21, 17, 30) {real, imag} */,
  {32'h4609043c, 32'h00000000} /* (21, 17, 29) {real, imag} */,
  {32'h460b3ad0, 32'h00000000} /* (21, 17, 28) {real, imag} */,
  {32'h4610ab3a, 32'h00000000} /* (21, 17, 27) {real, imag} */,
  {32'h45ff0fd6, 32'h00000000} /* (21, 17, 26) {real, imag} */,
  {32'h45ff9337, 32'h00000000} /* (21, 17, 25) {real, imag} */,
  {32'h45ec75f2, 32'h00000000} /* (21, 17, 24) {real, imag} */,
  {32'h45cc15ea, 32'h00000000} /* (21, 17, 23) {real, imag} */,
  {32'h4558cf98, 32'h00000000} /* (21, 17, 22) {real, imag} */,
  {32'h446ed30c, 32'h00000000} /* (21, 17, 21) {real, imag} */,
  {32'hc50eea10, 32'h00000000} /* (21, 17, 20) {real, imag} */,
  {32'hc5af446c, 32'h00000000} /* (21, 17, 19) {real, imag} */,
  {32'hc5f2436c, 32'h00000000} /* (21, 17, 18) {real, imag} */,
  {32'hc60d77c0, 32'h00000000} /* (21, 17, 17) {real, imag} */,
  {32'hc5fdeb8a, 32'h00000000} /* (21, 17, 16) {real, imag} */,
  {32'hc5eb4d56, 32'h00000000} /* (21, 17, 15) {real, imag} */,
  {32'hc5e29dee, 32'h00000000} /* (21, 17, 14) {real, imag} */,
  {32'hc5d123be, 32'h00000000} /* (21, 17, 13) {real, imag} */,
  {32'hc59afe36, 32'h00000000} /* (21, 17, 12) {real, imag} */,
  {32'hc54edf31, 32'h00000000} /* (21, 17, 11) {real, imag} */,
  {32'h4184de80, 32'h00000000} /* (21, 17, 10) {real, imag} */,
  {32'h45220aca, 32'h00000000} /* (21, 17, 9) {real, imag} */,
  {32'h4596699e, 32'h00000000} /* (21, 17, 8) {real, imag} */,
  {32'h45cab616, 32'h00000000} /* (21, 17, 7) {real, imag} */,
  {32'h45dc1f10, 32'h00000000} /* (21, 17, 6) {real, imag} */,
  {32'h460e5cd5, 32'h00000000} /* (21, 17, 5) {real, imag} */,
  {32'h4606b103, 32'h00000000} /* (21, 17, 4) {real, imag} */,
  {32'h4605d238, 32'h00000000} /* (21, 17, 3) {real, imag} */,
  {32'h4614e47e, 32'h00000000} /* (21, 17, 2) {real, imag} */,
  {32'h461c07a8, 32'h00000000} /* (21, 17, 1) {real, imag} */,
  {32'h45f9ae00, 32'h00000000} /* (21, 17, 0) {real, imag} */,
  {32'h46044780, 32'h00000000} /* (21, 16, 31) {real, imag} */,
  {32'h461275e2, 32'h00000000} /* (21, 16, 30) {real, imag} */,
  {32'h460dd01d, 32'h00000000} /* (21, 16, 29) {real, imag} */,
  {32'h461189cf, 32'h00000000} /* (21, 16, 28) {real, imag} */,
  {32'h4606c06a, 32'h00000000} /* (21, 16, 27) {real, imag} */,
  {32'h46118b7e, 32'h00000000} /* (21, 16, 26) {real, imag} */,
  {32'h45f6a16d, 32'h00000000} /* (21, 16, 25) {real, imag} */,
  {32'h45ede6fe, 32'h00000000} /* (21, 16, 24) {real, imag} */,
  {32'h45bc4e37, 32'h00000000} /* (21, 16, 23) {real, imag} */,
  {32'h456fb8fa, 32'h00000000} /* (21, 16, 22) {real, imag} */,
  {32'h4474db88, 32'h00000000} /* (21, 16, 21) {real, imag} */,
  {32'hc5738813, 32'h00000000} /* (21, 16, 20) {real, imag} */,
  {32'hc5c82b73, 32'h00000000} /* (21, 16, 19) {real, imag} */,
  {32'hc5db7cca, 32'h00000000} /* (21, 16, 18) {real, imag} */,
  {32'hc5eb390d, 32'h00000000} /* (21, 16, 17) {real, imag} */,
  {32'hc5da384c, 32'h00000000} /* (21, 16, 16) {real, imag} */,
  {32'hc5fba520, 32'h00000000} /* (21, 16, 15) {real, imag} */,
  {32'hc60667d8, 32'h00000000} /* (21, 16, 14) {real, imag} */,
  {32'hc5eb9016, 32'h00000000} /* (21, 16, 13) {real, imag} */,
  {32'hc5a5acaa, 32'h00000000} /* (21, 16, 12) {real, imag} */,
  {32'hc54af37e, 32'h00000000} /* (21, 16, 11) {real, imag} */,
  {32'h43f1ce00, 32'h00000000} /* (21, 16, 10) {real, imag} */,
  {32'h45687bd2, 32'h00000000} /* (21, 16, 9) {real, imag} */,
  {32'h45a855ae, 32'h00000000} /* (21, 16, 8) {real, imag} */,
  {32'h45cf8439, 32'h00000000} /* (21, 16, 7) {real, imag} */,
  {32'h45f8e8c5, 32'h00000000} /* (21, 16, 6) {real, imag} */,
  {32'h461586b2, 32'h00000000} /* (21, 16, 5) {real, imag} */,
  {32'h46100c2d, 32'h00000000} /* (21, 16, 4) {real, imag} */,
  {32'h46179654, 32'h00000000} /* (21, 16, 3) {real, imag} */,
  {32'h4619e2c3, 32'h00000000} /* (21, 16, 2) {real, imag} */,
  {32'h461a9d70, 32'h00000000} /* (21, 16, 1) {real, imag} */,
  {32'h4609e2ba, 32'h00000000} /* (21, 16, 0) {real, imag} */,
  {32'h4609046e, 32'h00000000} /* (21, 15, 31) {real, imag} */,
  {32'h46199bd4, 32'h00000000} /* (21, 15, 30) {real, imag} */,
  {32'h460d9d1a, 32'h00000000} /* (21, 15, 29) {real, imag} */,
  {32'h4612cadd, 32'h00000000} /* (21, 15, 28) {real, imag} */,
  {32'h4605ef00, 32'h00000000} /* (21, 15, 27) {real, imag} */,
  {32'h460d1dea, 32'h00000000} /* (21, 15, 26) {real, imag} */,
  {32'h4616d5fe, 32'h00000000} /* (21, 15, 25) {real, imag} */,
  {32'h45d2ca42, 32'h00000000} /* (21, 15, 24) {real, imag} */,
  {32'h45bf0f76, 32'h00000000} /* (21, 15, 23) {real, imag} */,
  {32'h4557dd66, 32'h00000000} /* (21, 15, 22) {real, imag} */,
  {32'h441ae034, 32'h00000000} /* (21, 15, 21) {real, imag} */,
  {32'hc5781cd2, 32'h00000000} /* (21, 15, 20) {real, imag} */,
  {32'hc59e59e5, 32'h00000000} /* (21, 15, 19) {real, imag} */,
  {32'hc5dd1b4c, 32'h00000000} /* (21, 15, 18) {real, imag} */,
  {32'hc5e1e166, 32'h00000000} /* (21, 15, 17) {real, imag} */,
  {32'hc5e8499e, 32'h00000000} /* (21, 15, 16) {real, imag} */,
  {32'hc5f88ce3, 32'h00000000} /* (21, 15, 15) {real, imag} */,
  {32'hc5eadb6c, 32'h00000000} /* (21, 15, 14) {real, imag} */,
  {32'hc5d74573, 32'h00000000} /* (21, 15, 13) {real, imag} */,
  {32'hc5b3ed6d, 32'h00000000} /* (21, 15, 12) {real, imag} */,
  {32'hc5525946, 32'h00000000} /* (21, 15, 11) {real, imag} */,
  {32'h44338c10, 32'h00000000} /* (21, 15, 10) {real, imag} */,
  {32'h457cbdf6, 32'h00000000} /* (21, 15, 9) {real, imag} */,
  {32'h45ad2656, 32'h00000000} /* (21, 15, 8) {real, imag} */,
  {32'h45d79d82, 32'h00000000} /* (21, 15, 7) {real, imag} */,
  {32'h45f26b15, 32'h00000000} /* (21, 15, 6) {real, imag} */,
  {32'h46080199, 32'h00000000} /* (21, 15, 5) {real, imag} */,
  {32'h4623463e, 32'h00000000} /* (21, 15, 4) {real, imag} */,
  {32'h461c3a2e, 32'h00000000} /* (21, 15, 3) {real, imag} */,
  {32'h460bb7df, 32'h00000000} /* (21, 15, 2) {real, imag} */,
  {32'h461bcc47, 32'h00000000} /* (21, 15, 1) {real, imag} */,
  {32'h4604301d, 32'h00000000} /* (21, 15, 0) {real, imag} */,
  {32'h45f10592, 32'h00000000} /* (21, 14, 31) {real, imag} */,
  {32'h460bb555, 32'h00000000} /* (21, 14, 30) {real, imag} */,
  {32'h4614b8cc, 32'h00000000} /* (21, 14, 29) {real, imag} */,
  {32'h460758e0, 32'h00000000} /* (21, 14, 28) {real, imag} */,
  {32'h46079afe, 32'h00000000} /* (21, 14, 27) {real, imag} */,
  {32'h46015682, 32'h00000000} /* (21, 14, 26) {real, imag} */,
  {32'h4600f63a, 32'h00000000} /* (21, 14, 25) {real, imag} */,
  {32'h45c88553, 32'h00000000} /* (21, 14, 24) {real, imag} */,
  {32'h459ab57a, 32'h00000000} /* (21, 14, 23) {real, imag} */,
  {32'h454f291b, 32'h00000000} /* (21, 14, 22) {real, imag} */,
  {32'h4465a80c, 32'h00000000} /* (21, 14, 21) {real, imag} */,
  {32'hc52d0678, 32'h00000000} /* (21, 14, 20) {real, imag} */,
  {32'hc595698f, 32'h00000000} /* (21, 14, 19) {real, imag} */,
  {32'hc5b73f28, 32'h00000000} /* (21, 14, 18) {real, imag} */,
  {32'hc5e83c60, 32'h00000000} /* (21, 14, 17) {real, imag} */,
  {32'hc5e4f5f8, 32'h00000000} /* (21, 14, 16) {real, imag} */,
  {32'hc5eeba4a, 32'h00000000} /* (21, 14, 15) {real, imag} */,
  {32'hc5d031ca, 32'h00000000} /* (21, 14, 14) {real, imag} */,
  {32'hc5c0b4fb, 32'h00000000} /* (21, 14, 13) {real, imag} */,
  {32'hc5a6d241, 32'h00000000} /* (21, 14, 12) {real, imag} */,
  {32'hc55e9986, 32'h00000000} /* (21, 14, 11) {real, imag} */,
  {32'h43fb7e98, 32'h00000000} /* (21, 14, 10) {real, imag} */,
  {32'h45660042, 32'h00000000} /* (21, 14, 9) {real, imag} */,
  {32'h45c53891, 32'h00000000} /* (21, 14, 8) {real, imag} */,
  {32'h45f0ed1c, 32'h00000000} /* (21, 14, 7) {real, imag} */,
  {32'h45efd41a, 32'h00000000} /* (21, 14, 6) {real, imag} */,
  {32'h460c9d71, 32'h00000000} /* (21, 14, 5) {real, imag} */,
  {32'h460f9747, 32'h00000000} /* (21, 14, 4) {real, imag} */,
  {32'h460131c7, 32'h00000000} /* (21, 14, 3) {real, imag} */,
  {32'h46102693, 32'h00000000} /* (21, 14, 2) {real, imag} */,
  {32'h4618b6f4, 32'h00000000} /* (21, 14, 1) {real, imag} */,
  {32'h45f593d8, 32'h00000000} /* (21, 14, 0) {real, imag} */,
  {32'h45c24f36, 32'h00000000} /* (21, 13, 31) {real, imag} */,
  {32'h45d6fefc, 32'h00000000} /* (21, 13, 30) {real, imag} */,
  {32'h45ea3410, 32'h00000000} /* (21, 13, 29) {real, imag} */,
  {32'h45db5a00, 32'h00000000} /* (21, 13, 28) {real, imag} */,
  {32'h45f795d3, 32'h00000000} /* (21, 13, 27) {real, imag} */,
  {32'h45e5425a, 32'h00000000} /* (21, 13, 26) {real, imag} */,
  {32'h45abf9a8, 32'h00000000} /* (21, 13, 25) {real, imag} */,
  {32'h45a8c112, 32'h00000000} /* (21, 13, 24) {real, imag} */,
  {32'h4588bc42, 32'h00000000} /* (21, 13, 23) {real, imag} */,
  {32'h458e20e5, 32'h00000000} /* (21, 13, 22) {real, imag} */,
  {32'h436be6f0, 32'h00000000} /* (21, 13, 21) {real, imag} */,
  {32'hc513a6a2, 32'h00000000} /* (21, 13, 20) {real, imag} */,
  {32'hc5a82423, 32'h00000000} /* (21, 13, 19) {real, imag} */,
  {32'hc5b907fd, 32'h00000000} /* (21, 13, 18) {real, imag} */,
  {32'hc5ab9aed, 32'h00000000} /* (21, 13, 17) {real, imag} */,
  {32'hc5c34a16, 32'h00000000} /* (21, 13, 16) {real, imag} */,
  {32'hc5bf4016, 32'h00000000} /* (21, 13, 15) {real, imag} */,
  {32'hc5b9eab4, 32'h00000000} /* (21, 13, 14) {real, imag} */,
  {32'hc5ad934a, 32'h00000000} /* (21, 13, 13) {real, imag} */,
  {32'hc57fcee8, 32'h00000000} /* (21, 13, 12) {real, imag} */,
  {32'hc538f8ce, 32'h00000000} /* (21, 13, 11) {real, imag} */,
  {32'h4458d480, 32'h00000000} /* (21, 13, 10) {real, imag} */,
  {32'h45716465, 32'h00000000} /* (21, 13, 9) {real, imag} */,
  {32'h45d1b0ae, 32'h00000000} /* (21, 13, 8) {real, imag} */,
  {32'h45deba7c, 32'h00000000} /* (21, 13, 7) {real, imag} */,
  {32'h45d2f203, 32'h00000000} /* (21, 13, 6) {real, imag} */,
  {32'h45f3345a, 32'h00000000} /* (21, 13, 5) {real, imag} */,
  {32'h45ef5d57, 32'h00000000} /* (21, 13, 4) {real, imag} */,
  {32'h45d61541, 32'h00000000} /* (21, 13, 3) {real, imag} */,
  {32'h45e240b7, 32'h00000000} /* (21, 13, 2) {real, imag} */,
  {32'h45fa070b, 32'h00000000} /* (21, 13, 1) {real, imag} */,
  {32'h45d5021a, 32'h00000000} /* (21, 13, 0) {real, imag} */,
  {32'h457f82c6, 32'h00000000} /* (21, 12, 31) {real, imag} */,
  {32'h45850c84, 32'h00000000} /* (21, 12, 30) {real, imag} */,
  {32'h4577fdf6, 32'h00000000} /* (21, 12, 29) {real, imag} */,
  {32'h458fea0a, 32'h00000000} /* (21, 12, 28) {real, imag} */,
  {32'h45a4d4e0, 32'h00000000} /* (21, 12, 27) {real, imag} */,
  {32'h4576de72, 32'h00000000} /* (21, 12, 26) {real, imag} */,
  {32'h456139a1, 32'h00000000} /* (21, 12, 25) {real, imag} */,
  {32'h4574a32c, 32'h00000000} /* (21, 12, 24) {real, imag} */,
  {32'h45717baa, 32'h00000000} /* (21, 12, 23) {real, imag} */,
  {32'h4558aeec, 32'h00000000} /* (21, 12, 22) {real, imag} */,
  {32'h433a8310, 32'h00000000} /* (21, 12, 21) {real, imag} */,
  {32'hc525f130, 32'h00000000} /* (21, 12, 20) {real, imag} */,
  {32'hc570639c, 32'h00000000} /* (21, 12, 19) {real, imag} */,
  {32'hc5a7b502, 32'h00000000} /* (21, 12, 18) {real, imag} */,
  {32'hc5a37b3a, 32'h00000000} /* (21, 12, 17) {real, imag} */,
  {32'hc58d4250, 32'h00000000} /* (21, 12, 16) {real, imag} */,
  {32'hc5810e4b, 32'h00000000} /* (21, 12, 15) {real, imag} */,
  {32'hc5a9ca1a, 32'h00000000} /* (21, 12, 14) {real, imag} */,
  {32'hc58185f7, 32'h00000000} /* (21, 12, 13) {real, imag} */,
  {32'hc510f956, 32'h00000000} /* (21, 12, 12) {real, imag} */,
  {32'hc4a0b7e6, 32'h00000000} /* (21, 12, 11) {real, imag} */,
  {32'h451bd404, 32'h00000000} /* (21, 12, 10) {real, imag} */,
  {32'h45807107, 32'h00000000} /* (21, 12, 9) {real, imag} */,
  {32'h459a3e16, 32'h00000000} /* (21, 12, 8) {real, imag} */,
  {32'h45a9bc2d, 32'h00000000} /* (21, 12, 7) {real, imag} */,
  {32'h45a26d76, 32'h00000000} /* (21, 12, 6) {real, imag} */,
  {32'h45a753ae, 32'h00000000} /* (21, 12, 5) {real, imag} */,
  {32'h45b1cd9e, 32'h00000000} /* (21, 12, 4) {real, imag} */,
  {32'h45872bcd, 32'h00000000} /* (21, 12, 3) {real, imag} */,
  {32'h4584a998, 32'h00000000} /* (21, 12, 2) {real, imag} */,
  {32'h459c6594, 32'h00000000} /* (21, 12, 1) {real, imag} */,
  {32'h45823af8, 32'h00000000} /* (21, 12, 0) {real, imag} */,
  {32'h44e39cd3, 32'h00000000} /* (21, 11, 31) {real, imag} */,
  {32'h4501b632, 32'h00000000} /* (21, 11, 30) {real, imag} */,
  {32'h44c9a65b, 32'h00000000} /* (21, 11, 29) {real, imag} */,
  {32'h44bf1684, 32'h00000000} /* (21, 11, 28) {real, imag} */,
  {32'h44aae569, 32'h00000000} /* (21, 11, 27) {real, imag} */,
  {32'h448b7a10, 32'h00000000} /* (21, 11, 26) {real, imag} */,
  {32'h44e87058, 32'h00000000} /* (21, 11, 25) {real, imag} */,
  {32'h44bf9068, 32'h00000000} /* (21, 11, 24) {real, imag} */,
  {32'h442a3a74, 32'h00000000} /* (21, 11, 23) {real, imag} */,
  {32'h44eb269b, 32'h00000000} /* (21, 11, 22) {real, imag} */,
  {32'hc4877e7b, 32'h00000000} /* (21, 11, 21) {real, imag} */,
  {32'hc50e9c9e, 32'h00000000} /* (21, 11, 20) {real, imag} */,
  {32'hc5152d3a, 32'h00000000} /* (21, 11, 19) {real, imag} */,
  {32'hc51c512e, 32'h00000000} /* (21, 11, 18) {real, imag} */,
  {32'hc5267fea, 32'h00000000} /* (21, 11, 17) {real, imag} */,
  {32'hc51d1a52, 32'h00000000} /* (21, 11, 16) {real, imag} */,
  {32'hc502ea64, 32'h00000000} /* (21, 11, 15) {real, imag} */,
  {32'hc4f90e5d, 32'h00000000} /* (21, 11, 14) {real, imag} */,
  {32'hc496346d, 32'h00000000} /* (21, 11, 13) {real, imag} */,
  {32'hc363e934, 32'h00000000} /* (21, 11, 12) {real, imag} */,
  {32'h42d18530, 32'h00000000} /* (21, 11, 11) {real, imag} */,
  {32'h452c1c0a, 32'h00000000} /* (21, 11, 10) {real, imag} */,
  {32'h45441850, 32'h00000000} /* (21, 11, 9) {real, imag} */,
  {32'h452cf09a, 32'h00000000} /* (21, 11, 8) {real, imag} */,
  {32'h457bfdad, 32'h00000000} /* (21, 11, 7) {real, imag} */,
  {32'h457e6582, 32'h00000000} /* (21, 11, 6) {real, imag} */,
  {32'h455701ac, 32'h00000000} /* (21, 11, 5) {real, imag} */,
  {32'h452e4dd0, 32'h00000000} /* (21, 11, 4) {real, imag} */,
  {32'h44cd2208, 32'h00000000} /* (21, 11, 3) {real, imag} */,
  {32'h450b89dc, 32'h00000000} /* (21, 11, 2) {real, imag} */,
  {32'h451d3910, 32'h00000000} /* (21, 11, 1) {real, imag} */,
  {32'h44e55e3c, 32'h00000000} /* (21, 11, 0) {real, imag} */,
  {32'hc4c57569, 32'h00000000} /* (21, 10, 31) {real, imag} */,
  {32'hc4e2b2e2, 32'h00000000} /* (21, 10, 30) {real, imag} */,
  {32'hc5231f98, 32'h00000000} /* (21, 10, 29) {real, imag} */,
  {32'hc525f4c2, 32'h00000000} /* (21, 10, 28) {real, imag} */,
  {32'hc56cea54, 32'h00000000} /* (21, 10, 27) {real, imag} */,
  {32'hc5298f81, 32'h00000000} /* (21, 10, 26) {real, imag} */,
  {32'hc51db8d0, 32'h00000000} /* (21, 10, 25) {real, imag} */,
  {32'hc5193844, 32'h00000000} /* (21, 10, 24) {real, imag} */,
  {32'hc504e9b9, 32'h00000000} /* (21, 10, 23) {real, imag} */,
  {32'hc548f65f, 32'h00000000} /* (21, 10, 22) {real, imag} */,
  {32'hc515bb5c, 32'h00000000} /* (21, 10, 21) {real, imag} */,
  {32'hc3e41f66, 32'h00000000} /* (21, 10, 20) {real, imag} */,
  {32'hc42c9772, 32'h00000000} /* (21, 10, 19) {real, imag} */,
  {32'hc404db04, 32'h00000000} /* (21, 10, 18) {real, imag} */,
  {32'h42c323a0, 32'h00000000} /* (21, 10, 17) {real, imag} */,
  {32'h44875eb4, 32'h00000000} /* (21, 10, 16) {real, imag} */,
  {32'h448ff1eb, 32'h00000000} /* (21, 10, 15) {real, imag} */,
  {32'h44c80dc2, 32'h00000000} /* (21, 10, 14) {real, imag} */,
  {32'h44a99567, 32'h00000000} /* (21, 10, 13) {real, imag} */,
  {32'h4505c71c, 32'h00000000} /* (21, 10, 12) {real, imag} */,
  {32'h44c4cf80, 32'h00000000} /* (21, 10, 11) {real, imag} */,
  {32'h44587cc0, 32'h00000000} /* (21, 10, 10) {real, imag} */,
  {32'h43409bc8, 32'h00000000} /* (21, 10, 9) {real, imag} */,
  {32'h442864ac, 32'h00000000} /* (21, 10, 8) {real, imag} */,
  {32'h443abc80, 32'h00000000} /* (21, 10, 7) {real, imag} */,
  {32'h43849a88, 32'h00000000} /* (21, 10, 6) {real, imag} */,
  {32'hc479a22b, 32'h00000000} /* (21, 10, 5) {real, imag} */,
  {32'hc4a53dce, 32'h00000000} /* (21, 10, 4) {real, imag} */,
  {32'hc4f39947, 32'h00000000} /* (21, 10, 3) {real, imag} */,
  {32'hc464a7d0, 32'h00000000} /* (21, 10, 2) {real, imag} */,
  {32'hc5008309, 32'h00000000} /* (21, 10, 1) {real, imag} */,
  {32'hc4fb04a6, 32'h00000000} /* (21, 10, 0) {real, imag} */,
  {32'hc5959fc9, 32'h00000000} /* (21, 9, 31) {real, imag} */,
  {32'hc5a504ec, 32'h00000000} /* (21, 9, 30) {real, imag} */,
  {32'hc5df45e1, 32'h00000000} /* (21, 9, 29) {real, imag} */,
  {32'hc5bfe084, 32'h00000000} /* (21, 9, 28) {real, imag} */,
  {32'hc5c8525c, 32'h00000000} /* (21, 9, 27) {real, imag} */,
  {32'hc5cc5bab, 32'h00000000} /* (21, 9, 26) {real, imag} */,
  {32'hc5bb0f7b, 32'h00000000} /* (21, 9, 25) {real, imag} */,
  {32'hc5ae1096, 32'h00000000} /* (21, 9, 24) {real, imag} */,
  {32'hc5b54862, 32'h00000000} /* (21, 9, 23) {real, imag} */,
  {32'hc591926d, 32'h00000000} /* (21, 9, 22) {real, imag} */,
  {32'hc56ca491, 32'h00000000} /* (21, 9, 21) {real, imag} */,
  {32'h42374500, 32'h00000000} /* (21, 9, 20) {real, imag} */,
  {32'h4431b28c, 32'h00000000} /* (21, 9, 19) {real, imag} */,
  {32'h447cfcb4, 32'h00000000} /* (21, 9, 18) {real, imag} */,
  {32'h450663d8, 32'h00000000} /* (21, 9, 17) {real, imag} */,
  {32'h4576368c, 32'h00000000} /* (21, 9, 16) {real, imag} */,
  {32'h456ced0e, 32'h00000000} /* (21, 9, 15) {real, imag} */,
  {32'h456afd30, 32'h00000000} /* (21, 9, 14) {real, imag} */,
  {32'h45621672, 32'h00000000} /* (21, 9, 13) {real, imag} */,
  {32'h453d7795, 32'h00000000} /* (21, 9, 12) {real, imag} */,
  {32'h4534eff9, 32'h00000000} /* (21, 9, 11) {real, imag} */,
  {32'h449ded6c, 32'h00000000} /* (21, 9, 10) {real, imag} */,
  {32'hc4983134, 32'h00000000} /* (21, 9, 9) {real, imag} */,
  {32'hc4ff9bb0, 32'h00000000} /* (21, 9, 8) {real, imag} */,
  {32'hc526b4a3, 32'h00000000} /* (21, 9, 7) {real, imag} */,
  {32'hc5824993, 32'h00000000} /* (21, 9, 6) {real, imag} */,
  {32'hc57b748f, 32'h00000000} /* (21, 9, 5) {real, imag} */,
  {32'hc5ad12d7, 32'h00000000} /* (21, 9, 4) {real, imag} */,
  {32'hc596b330, 32'h00000000} /* (21, 9, 3) {real, imag} */,
  {32'hc59d0d16, 32'h00000000} /* (21, 9, 2) {real, imag} */,
  {32'hc58d93c0, 32'h00000000} /* (21, 9, 1) {real, imag} */,
  {32'hc5972292, 32'h00000000} /* (21, 9, 0) {real, imag} */,
  {32'hc5eaf120, 32'h00000000} /* (21, 8, 31) {real, imag} */,
  {32'hc6052cb6, 32'h00000000} /* (21, 8, 30) {real, imag} */,
  {32'hc6136aa6, 32'h00000000} /* (21, 8, 29) {real, imag} */,
  {32'hc61644be, 32'h00000000} /* (21, 8, 28) {real, imag} */,
  {32'hc606f106, 32'h00000000} /* (21, 8, 27) {real, imag} */,
  {32'hc608947a, 32'h00000000} /* (21, 8, 26) {real, imag} */,
  {32'hc60c76f6, 32'h00000000} /* (21, 8, 25) {real, imag} */,
  {32'hc5f1fcb7, 32'h00000000} /* (21, 8, 24) {real, imag} */,
  {32'hc5ea54ce, 32'h00000000} /* (21, 8, 23) {real, imag} */,
  {32'hc5d1d514, 32'h00000000} /* (21, 8, 22) {real, imag} */,
  {32'hc59af022, 32'h00000000} /* (21, 8, 21) {real, imag} */,
  {32'hc49bf8e0, 32'h00000000} /* (21, 8, 20) {real, imag} */,
  {32'h449891ec, 32'h00000000} /* (21, 8, 19) {real, imag} */,
  {32'h4510a79a, 32'h00000000} /* (21, 8, 18) {real, imag} */,
  {32'h4579f80c, 32'h00000000} /* (21, 8, 17) {real, imag} */,
  {32'h4582caa6, 32'h00000000} /* (21, 8, 16) {real, imag} */,
  {32'h45ba2eea, 32'h00000000} /* (21, 8, 15) {real, imag} */,
  {32'h45b2070e, 32'h00000000} /* (21, 8, 14) {real, imag} */,
  {32'h459dfddf, 32'h00000000} /* (21, 8, 13) {real, imag} */,
  {32'h45819622, 32'h00000000} /* (21, 8, 12) {real, imag} */,
  {32'h458687d7, 32'h00000000} /* (21, 8, 11) {real, imag} */,
  {32'h44b9e5c4, 32'h00000000} /* (21, 8, 10) {real, imag} */,
  {32'hc44dee08, 32'h00000000} /* (21, 8, 9) {real, imag} */,
  {32'hc50ce9aa, 32'h00000000} /* (21, 8, 8) {real, imag} */,
  {32'hc53cc171, 32'h00000000} /* (21, 8, 7) {real, imag} */,
  {32'hc58f4636, 32'h00000000} /* (21, 8, 6) {real, imag} */,
  {32'hc5b32680, 32'h00000000} /* (21, 8, 5) {real, imag} */,
  {32'hc5b5bbbb, 32'h00000000} /* (21, 8, 4) {real, imag} */,
  {32'hc5d40d85, 32'h00000000} /* (21, 8, 3) {real, imag} */,
  {32'hc5ec1243, 32'h00000000} /* (21, 8, 2) {real, imag} */,
  {32'hc5e5331e, 32'h00000000} /* (21, 8, 1) {real, imag} */,
  {32'hc5c4721e, 32'h00000000} /* (21, 8, 0) {real, imag} */,
  {32'hc6188ff3, 32'h00000000} /* (21, 7, 31) {real, imag} */,
  {32'hc62c02c4, 32'h00000000} /* (21, 7, 30) {real, imag} */,
  {32'hc639b26a, 32'h00000000} /* (21, 7, 29) {real, imag} */,
  {32'hc62552aa, 32'h00000000} /* (21, 7, 28) {real, imag} */,
  {32'hc6290670, 32'h00000000} /* (21, 7, 27) {real, imag} */,
  {32'hc632eb44, 32'h00000000} /* (21, 7, 26) {real, imag} */,
  {32'hc62ef2f6, 32'h00000000} /* (21, 7, 25) {real, imag} */,
  {32'hc61e2f28, 32'h00000000} /* (21, 7, 24) {real, imag} */,
  {32'hc607f658, 32'h00000000} /* (21, 7, 23) {real, imag} */,
  {32'hc5f0c93e, 32'h00000000} /* (21, 7, 22) {real, imag} */,
  {32'hc5b138c2, 32'h00000000} /* (21, 7, 21) {real, imag} */,
  {32'hc5034dd0, 32'h00000000} /* (21, 7, 20) {real, imag} */,
  {32'h43963e80, 32'h00000000} /* (21, 7, 19) {real, imag} */,
  {32'h451a0a66, 32'h00000000} /* (21, 7, 18) {real, imag} */,
  {32'h4542081a, 32'h00000000} /* (21, 7, 17) {real, imag} */,
  {32'h45ac873c, 32'h00000000} /* (21, 7, 16) {real, imag} */,
  {32'h45c2d58c, 32'h00000000} /* (21, 7, 15) {real, imag} */,
  {32'h45d6e7dc, 32'h00000000} /* (21, 7, 14) {real, imag} */,
  {32'h45bf96b4, 32'h00000000} /* (21, 7, 13) {real, imag} */,
  {32'h45b4b6ed, 32'h00000000} /* (21, 7, 12) {real, imag} */,
  {32'h456be826, 32'h00000000} /* (21, 7, 11) {real, imag} */,
  {32'h4504155e, 32'h00000000} /* (21, 7, 10) {real, imag} */,
  {32'hc240ce80, 32'h00000000} /* (21, 7, 9) {real, imag} */,
  {32'hc4edf480, 32'h00000000} /* (21, 7, 8) {real, imag} */,
  {32'hc54f0550, 32'h00000000} /* (21, 7, 7) {real, imag} */,
  {32'hc59e9026, 32'h00000000} /* (21, 7, 6) {real, imag} */,
  {32'hc5d0f7f2, 32'h00000000} /* (21, 7, 5) {real, imag} */,
  {32'hc5f9f002, 32'h00000000} /* (21, 7, 4) {real, imag} */,
  {32'hc5fdf5c8, 32'h00000000} /* (21, 7, 3) {real, imag} */,
  {32'hc6119420, 32'h00000000} /* (21, 7, 2) {real, imag} */,
  {32'hc612c8a8, 32'h00000000} /* (21, 7, 1) {real, imag} */,
  {32'hc60943b1, 32'h00000000} /* (21, 7, 0) {real, imag} */,
  {32'hc6299a7a, 32'h00000000} /* (21, 6, 31) {real, imag} */,
  {32'hc62cdaeb, 32'h00000000} /* (21, 6, 30) {real, imag} */,
  {32'hc6314f6a, 32'h00000000} /* (21, 6, 29) {real, imag} */,
  {32'hc63ed4b4, 32'h00000000} /* (21, 6, 28) {real, imag} */,
  {32'hc645c6fa, 32'h00000000} /* (21, 6, 27) {real, imag} */,
  {32'hc63d169f, 32'h00000000} /* (21, 6, 26) {real, imag} */,
  {32'hc6430cb2, 32'h00000000} /* (21, 6, 25) {real, imag} */,
  {32'hc62db2d6, 32'h00000000} /* (21, 6, 24) {real, imag} */,
  {32'hc6160070, 32'h00000000} /* (21, 6, 23) {real, imag} */,
  {32'hc6037b63, 32'h00000000} /* (21, 6, 22) {real, imag} */,
  {32'hc5d09315, 32'h00000000} /* (21, 6, 21) {real, imag} */,
  {32'hc54b769a, 32'h00000000} /* (21, 6, 20) {real, imag} */,
  {32'hc4561338, 32'h00000000} /* (21, 6, 19) {real, imag} */,
  {32'h44e6b464, 32'h00000000} /* (21, 6, 18) {real, imag} */,
  {32'h4530d154, 32'h00000000} /* (21, 6, 17) {real, imag} */,
  {32'h458f5ed2, 32'h00000000} /* (21, 6, 16) {real, imag} */,
  {32'h45d29f98, 32'h00000000} /* (21, 6, 15) {real, imag} */,
  {32'h45e72916, 32'h00000000} /* (21, 6, 14) {real, imag} */,
  {32'h45fd51b4, 32'h00000000} /* (21, 6, 13) {real, imag} */,
  {32'h45b63709, 32'h00000000} /* (21, 6, 12) {real, imag} */,
  {32'h4587e309, 32'h00000000} /* (21, 6, 11) {real, imag} */,
  {32'h451e511c, 32'h00000000} /* (21, 6, 10) {real, imag} */,
  {32'h440ae2b8, 32'h00000000} /* (21, 6, 9) {real, imag} */,
  {32'hc4c01da4, 32'h00000000} /* (21, 6, 8) {real, imag} */,
  {32'hc4f81474, 32'h00000000} /* (21, 6, 7) {real, imag} */,
  {32'hc59a5af2, 32'h00000000} /* (21, 6, 6) {real, imag} */,
  {32'hc5d02a0b, 32'h00000000} /* (21, 6, 5) {real, imag} */,
  {32'hc5e7825d, 32'h00000000} /* (21, 6, 4) {real, imag} */,
  {32'hc61978c8, 32'h00000000} /* (21, 6, 3) {real, imag} */,
  {32'hc6274d28, 32'h00000000} /* (21, 6, 2) {real, imag} */,
  {32'hc61e9562, 32'h00000000} /* (21, 6, 1) {real, imag} */,
  {32'hc61d766a, 32'h00000000} /* (21, 6, 0) {real, imag} */,
  {32'hc633dae8, 32'h00000000} /* (21, 5, 31) {real, imag} */,
  {32'hc6455270, 32'h00000000} /* (21, 5, 30) {real, imag} */,
  {32'hc64dda1f, 32'h00000000} /* (21, 5, 29) {real, imag} */,
  {32'hc64d63ea, 32'h00000000} /* (21, 5, 28) {real, imag} */,
  {32'hc6560c41, 32'h00000000} /* (21, 5, 27) {real, imag} */,
  {32'hc6584831, 32'h00000000} /* (21, 5, 26) {real, imag} */,
  {32'hc64b6c78, 32'h00000000} /* (21, 5, 25) {real, imag} */,
  {32'hc6377a76, 32'h00000000} /* (21, 5, 24) {real, imag} */,
  {32'hc62448e5, 32'h00000000} /* (21, 5, 23) {real, imag} */,
  {32'hc61446a0, 32'h00000000} /* (21, 5, 22) {real, imag} */,
  {32'hc6074416, 32'h00000000} /* (21, 5, 21) {real, imag} */,
  {32'hc5b49c1e, 32'h00000000} /* (21, 5, 20) {real, imag} */,
  {32'hc5341db2, 32'h00000000} /* (21, 5, 19) {real, imag} */,
  {32'hc4175468, 32'h00000000} /* (21, 5, 18) {real, imag} */,
  {32'h44025260, 32'h00000000} /* (21, 5, 17) {real, imag} */,
  {32'h453df7f0, 32'h00000000} /* (21, 5, 16) {real, imag} */,
  {32'h45b66814, 32'h00000000} /* (21, 5, 15) {real, imag} */,
  {32'h45e19187, 32'h00000000} /* (21, 5, 14) {real, imag} */,
  {32'h45f2ac4e, 32'h00000000} /* (21, 5, 13) {real, imag} */,
  {32'h45cfcb69, 32'h00000000} /* (21, 5, 12) {real, imag} */,
  {32'h45bbda8e, 32'h00000000} /* (21, 5, 11) {real, imag} */,
  {32'h459dca16, 32'h00000000} /* (21, 5, 10) {real, imag} */,
  {32'h453a3996, 32'h00000000} /* (21, 5, 9) {real, imag} */,
  {32'h451af102, 32'h00000000} /* (21, 5, 8) {real, imag} */,
  {32'h443de0d0, 32'h00000000} /* (21, 5, 7) {real, imag} */,
  {32'hc5450afb, 32'h00000000} /* (21, 5, 6) {real, imag} */,
  {32'hc5b03370, 32'h00000000} /* (21, 5, 5) {real, imag} */,
  {32'hc60356c6, 32'h00000000} /* (21, 5, 4) {real, imag} */,
  {32'hc6212744, 32'h00000000} /* (21, 5, 3) {real, imag} */,
  {32'hc625bce8, 32'h00000000} /* (21, 5, 2) {real, imag} */,
  {32'hc62d51f5, 32'h00000000} /* (21, 5, 1) {real, imag} */,
  {32'hc6317104, 32'h00000000} /* (21, 5, 0) {real, imag} */,
  {32'hc6387873, 32'h00000000} /* (21, 4, 31) {real, imag} */,
  {32'hc642f74e, 32'h00000000} /* (21, 4, 30) {real, imag} */,
  {32'hc6509cf2, 32'h00000000} /* (21, 4, 29) {real, imag} */,
  {32'hc6529eaf, 32'h00000000} /* (21, 4, 28) {real, imag} */,
  {32'hc65dbf67, 32'h00000000} /* (21, 4, 27) {real, imag} */,
  {32'hc666eb56, 32'h00000000} /* (21, 4, 26) {real, imag} */,
  {32'hc658e0ce, 32'h00000000} /* (21, 4, 25) {real, imag} */,
  {32'hc65a1566, 32'h00000000} /* (21, 4, 24) {real, imag} */,
  {32'hc63b05ec, 32'h00000000} /* (21, 4, 23) {real, imag} */,
  {32'hc613e7b0, 32'h00000000} /* (21, 4, 22) {real, imag} */,
  {32'hc60ae809, 32'h00000000} /* (21, 4, 21) {real, imag} */,
  {32'hc5ff826a, 32'h00000000} /* (21, 4, 20) {real, imag} */,
  {32'hc5bc6b15, 32'h00000000} /* (21, 4, 19) {real, imag} */,
  {32'hc561acfe, 32'h00000000} /* (21, 4, 18) {real, imag} */,
  {32'hc474d3c0, 32'h00000000} /* (21, 4, 17) {real, imag} */,
  {32'h44611b00, 32'h00000000} /* (21, 4, 16) {real, imag} */,
  {32'h45773793, 32'h00000000} /* (21, 4, 15) {real, imag} */,
  {32'h45d76ec8, 32'h00000000} /* (21, 4, 14) {real, imag} */,
  {32'h45e5b7a4, 32'h00000000} /* (21, 4, 13) {real, imag} */,
  {32'h45d13eb2, 32'h00000000} /* (21, 4, 12) {real, imag} */,
  {32'h45c6867a, 32'h00000000} /* (21, 4, 11) {real, imag} */,
  {32'h45c903f3, 32'h00000000} /* (21, 4, 10) {real, imag} */,
  {32'h45923da9, 32'h00000000} /* (21, 4, 9) {real, imag} */,
  {32'h45265c2a, 32'h00000000} /* (21, 4, 8) {real, imag} */,
  {32'h44e407e0, 32'h00000000} /* (21, 4, 7) {real, imag} */,
  {32'hc42d9820, 32'h00000000} /* (21, 4, 6) {real, imag} */,
  {32'hc59a9242, 32'h00000000} /* (21, 4, 5) {real, imag} */,
  {32'hc5ed473e, 32'h00000000} /* (21, 4, 4) {real, imag} */,
  {32'hc625ccda, 32'h00000000} /* (21, 4, 3) {real, imag} */,
  {32'hc63c879c, 32'h00000000} /* (21, 4, 2) {real, imag} */,
  {32'hc6346755, 32'h00000000} /* (21, 4, 1) {real, imag} */,
  {32'hc63b2e47, 32'h00000000} /* (21, 4, 0) {real, imag} */,
  {32'hc64797b0, 32'h00000000} /* (21, 3, 31) {real, imag} */,
  {32'hc6630282, 32'h00000000} /* (21, 3, 30) {real, imag} */,
  {32'hc65a3d2e, 32'h00000000} /* (21, 3, 29) {real, imag} */,
  {32'hc665b822, 32'h00000000} /* (21, 3, 28) {real, imag} */,
  {32'hc6692019, 32'h00000000} /* (21, 3, 27) {real, imag} */,
  {32'hc65a5c57, 32'h00000000} /* (21, 3, 26) {real, imag} */,
  {32'hc654cd66, 32'h00000000} /* (21, 3, 25) {real, imag} */,
  {32'hc6574588, 32'h00000000} /* (21, 3, 24) {real, imag} */,
  {32'hc643e1e8, 32'h00000000} /* (21, 3, 23) {real, imag} */,
  {32'hc62ddb54, 32'h00000000} /* (21, 3, 22) {real, imag} */,
  {32'hc617cd19, 32'h00000000} /* (21, 3, 21) {real, imag} */,
  {32'hc5ee067f, 32'h00000000} /* (21, 3, 20) {real, imag} */,
  {32'hc5c694c1, 32'h00000000} /* (21, 3, 19) {real, imag} */,
  {32'hc5845d3c, 32'h00000000} /* (21, 3, 18) {real, imag} */,
  {32'hc5480f02, 32'h00000000} /* (21, 3, 17) {real, imag} */,
  {32'h432fdbe0, 32'h00000000} /* (21, 3, 16) {real, imag} */,
  {32'h4587b7f7, 32'h00000000} /* (21, 3, 15) {real, imag} */,
  {32'h45c934fc, 32'h00000000} /* (21, 3, 14) {real, imag} */,
  {32'h45dfa714, 32'h00000000} /* (21, 3, 13) {real, imag} */,
  {32'h45dbd67b, 32'h00000000} /* (21, 3, 12) {real, imag} */,
  {32'h45d2248e, 32'h00000000} /* (21, 3, 11) {real, imag} */,
  {32'h45aeb93a, 32'h00000000} /* (21, 3, 10) {real, imag} */,
  {32'h458f31f5, 32'h00000000} /* (21, 3, 9) {real, imag} */,
  {32'h455208ee, 32'h00000000} /* (21, 3, 8) {real, imag} */,
  {32'h453e74ec, 32'h00000000} /* (21, 3, 7) {real, imag} */,
  {32'hc3f117c0, 32'h00000000} /* (21, 3, 6) {real, imag} */,
  {32'hc5887c9a, 32'h00000000} /* (21, 3, 5) {real, imag} */,
  {32'hc5e443db, 32'h00000000} /* (21, 3, 4) {real, imag} */,
  {32'hc6281ee8, 32'h00000000} /* (21, 3, 3) {real, imag} */,
  {32'hc637637e, 32'h00000000} /* (21, 3, 2) {real, imag} */,
  {32'hc64cdae6, 32'h00000000} /* (21, 3, 1) {real, imag} */,
  {32'hc63b28ec, 32'h00000000} /* (21, 3, 0) {real, imag} */,
  {32'hc648bff5, 32'h00000000} /* (21, 2, 31) {real, imag} */,
  {32'hc65a3f2a, 32'h00000000} /* (21, 2, 30) {real, imag} */,
  {32'hc66120e1, 32'h00000000} /* (21, 2, 29) {real, imag} */,
  {32'hc662bfbe, 32'h00000000} /* (21, 2, 28) {real, imag} */,
  {32'hc65e8dae, 32'h00000000} /* (21, 2, 27) {real, imag} */,
  {32'hc65a1df0, 32'h00000000} /* (21, 2, 26) {real, imag} */,
  {32'hc65e1e32, 32'h00000000} /* (21, 2, 25) {real, imag} */,
  {32'hc64fbf05, 32'h00000000} /* (21, 2, 24) {real, imag} */,
  {32'hc63fd941, 32'h00000000} /* (21, 2, 23) {real, imag} */,
  {32'hc629ba48, 32'h00000000} /* (21, 2, 22) {real, imag} */,
  {32'hc61c6e07, 32'h00000000} /* (21, 2, 21) {real, imag} */,
  {32'hc5eb1832, 32'h00000000} /* (21, 2, 20) {real, imag} */,
  {32'hc5ba494f, 32'h00000000} /* (21, 2, 19) {real, imag} */,
  {32'hc575a3da, 32'h00000000} /* (21, 2, 18) {real, imag} */,
  {32'hc4d619cc, 32'h00000000} /* (21, 2, 17) {real, imag} */,
  {32'h43b75d40, 32'h00000000} /* (21, 2, 16) {real, imag} */,
  {32'h4558f998, 32'h00000000} /* (21, 2, 15) {real, imag} */,
  {32'h45b6b671, 32'h00000000} /* (21, 2, 14) {real, imag} */,
  {32'h45d43dd6, 32'h00000000} /* (21, 2, 13) {real, imag} */,
  {32'h45ce24d8, 32'h00000000} /* (21, 2, 12) {real, imag} */,
  {32'h45c44610, 32'h00000000} /* (21, 2, 11) {real, imag} */,
  {32'h45b0bd8f, 32'h00000000} /* (21, 2, 10) {real, imag} */,
  {32'h4598ad17, 32'h00000000} /* (21, 2, 9) {real, imag} */,
  {32'h4554eb04, 32'h00000000} /* (21, 2, 8) {real, imag} */,
  {32'h44da4700, 32'h00000000} /* (21, 2, 7) {real, imag} */,
  {32'hc42d20d8, 32'h00000000} /* (21, 2, 6) {real, imag} */,
  {32'hc5825652, 32'h00000000} /* (21, 2, 5) {real, imag} */,
  {32'hc6010cd5, 32'h00000000} /* (21, 2, 4) {real, imag} */,
  {32'hc617a6ea, 32'h00000000} /* (21, 2, 3) {real, imag} */,
  {32'hc63ecc22, 32'h00000000} /* (21, 2, 2) {real, imag} */,
  {32'hc6480f62, 32'h00000000} /* (21, 2, 1) {real, imag} */,
  {32'hc638e72e, 32'h00000000} /* (21, 2, 0) {real, imag} */,
  {32'hc6410171, 32'h00000000} /* (21, 1, 31) {real, imag} */,
  {32'hc64babc8, 32'h00000000} /* (21, 1, 30) {real, imag} */,
  {32'hc667e9f1, 32'h00000000} /* (21, 1, 29) {real, imag} */,
  {32'hc6672bc3, 32'h00000000} /* (21, 1, 28) {real, imag} */,
  {32'hc66a1215, 32'h00000000} /* (21, 1, 27) {real, imag} */,
  {32'hc662ea64, 32'h00000000} /* (21, 1, 26) {real, imag} */,
  {32'hc6587e52, 32'h00000000} /* (21, 1, 25) {real, imag} */,
  {32'hc6500dee, 32'h00000000} /* (21, 1, 24) {real, imag} */,
  {32'hc649a1a6, 32'h00000000} /* (21, 1, 23) {real, imag} */,
  {32'hc628d38c, 32'h00000000} /* (21, 1, 22) {real, imag} */,
  {32'hc610f064, 32'h00000000} /* (21, 1, 21) {real, imag} */,
  {32'hc5f07e08, 32'h00000000} /* (21, 1, 20) {real, imag} */,
  {32'hc5a3bc9c, 32'h00000000} /* (21, 1, 19) {real, imag} */,
  {32'hc55175ac, 32'h00000000} /* (21, 1, 18) {real, imag} */,
  {32'hc4791318, 32'h00000000} /* (21, 1, 17) {real, imag} */,
  {32'h43e1cc30, 32'h00000000} /* (21, 1, 16) {real, imag} */,
  {32'h456280ac, 32'h00000000} /* (21, 1, 15) {real, imag} */,
  {32'h45bc39f0, 32'h00000000} /* (21, 1, 14) {real, imag} */,
  {32'h45c988b6, 32'h00000000} /* (21, 1, 13) {real, imag} */,
  {32'h45db646a, 32'h00000000} /* (21, 1, 12) {real, imag} */,
  {32'h45b3b41a, 32'h00000000} /* (21, 1, 11) {real, imag} */,
  {32'h45b0474c, 32'h00000000} /* (21, 1, 10) {real, imag} */,
  {32'h45746828, 32'h00000000} /* (21, 1, 9) {real, imag} */,
  {32'h4506e742, 32'h00000000} /* (21, 1, 8) {real, imag} */,
  {32'hc38fa830, 32'h00000000} /* (21, 1, 7) {real, imag} */,
  {32'hc4a92850, 32'h00000000} /* (21, 1, 6) {real, imag} */,
  {32'hc59eaf0c, 32'h00000000} /* (21, 1, 5) {real, imag} */,
  {32'hc5fe8e88, 32'h00000000} /* (21, 1, 4) {real, imag} */,
  {32'hc624d6e8, 32'h00000000} /* (21, 1, 3) {real, imag} */,
  {32'hc64000f9, 32'h00000000} /* (21, 1, 2) {real, imag} */,
  {32'hc636b552, 32'h00000000} /* (21, 1, 1) {real, imag} */,
  {32'hc635b1de, 32'h00000000} /* (21, 1, 0) {real, imag} */,
  {32'hc640efb8, 32'h00000000} /* (21, 0, 31) {real, imag} */,
  {32'hc64ba30e, 32'h00000000} /* (21, 0, 30) {real, imag} */,
  {32'hc651ab75, 32'h00000000} /* (21, 0, 29) {real, imag} */,
  {32'hc657e54d, 32'h00000000} /* (21, 0, 28) {real, imag} */,
  {32'hc666ea9f, 32'h00000000} /* (21, 0, 27) {real, imag} */,
  {32'hc66249c7, 32'h00000000} /* (21, 0, 26) {real, imag} */,
  {32'hc6474bb0, 32'h00000000} /* (21, 0, 25) {real, imag} */,
  {32'hc63a4c6c, 32'h00000000} /* (21, 0, 24) {real, imag} */,
  {32'hc62f725a, 32'h00000000} /* (21, 0, 23) {real, imag} */,
  {32'hc6144aa6, 32'h00000000} /* (21, 0, 22) {real, imag} */,
  {32'hc5ddba97, 32'h00000000} /* (21, 0, 21) {real, imag} */,
  {32'hc5c3cc37, 32'h00000000} /* (21, 0, 20) {real, imag} */,
  {32'hc55cfa19, 32'h00000000} /* (21, 0, 19) {real, imag} */,
  {32'hc4bd44f8, 32'h00000000} /* (21, 0, 18) {real, imag} */,
  {32'hc4643548, 32'h00000000} /* (21, 0, 17) {real, imag} */,
  {32'h44edb084, 32'h00000000} /* (21, 0, 16) {real, imag} */,
  {32'h45902a28, 32'h00000000} /* (21, 0, 15) {real, imag} */,
  {32'h45a76829, 32'h00000000} /* (21, 0, 14) {real, imag} */,
  {32'h45d16332, 32'h00000000} /* (21, 0, 13) {real, imag} */,
  {32'h45c389d6, 32'h00000000} /* (21, 0, 12) {real, imag} */,
  {32'h45abd702, 32'h00000000} /* (21, 0, 11) {real, imag} */,
  {32'h457d4dac, 32'h00000000} /* (21, 0, 10) {real, imag} */,
  {32'h45121f06, 32'h00000000} /* (21, 0, 9) {real, imag} */,
  {32'hc279ae00, 32'h00000000} /* (21, 0, 8) {real, imag} */,
  {32'hc4cb3390, 32'h00000000} /* (21, 0, 7) {real, imag} */,
  {32'hc56fc5a2, 32'h00000000} /* (21, 0, 6) {real, imag} */,
  {32'hc5bbae11, 32'h00000000} /* (21, 0, 5) {real, imag} */,
  {32'hc606e94f, 32'h00000000} /* (21, 0, 4) {real, imag} */,
  {32'hc616b6f4, 32'h00000000} /* (21, 0, 3) {real, imag} */,
  {32'hc62760c9, 32'h00000000} /* (21, 0, 2) {real, imag} */,
  {32'hc639043c, 32'h00000000} /* (21, 0, 1) {real, imag} */,
  {32'hc639c326, 32'h00000000} /* (21, 0, 0) {real, imag} */,
  {32'hc63ff12e, 32'h00000000} /* (20, 31, 31) {real, imag} */,
  {32'hc6490776, 32'h00000000} /* (20, 31, 30) {real, imag} */,
  {32'hc649f40c, 32'h00000000} /* (20, 31, 29) {real, imag} */,
  {32'hc64e3ff2, 32'h00000000} /* (20, 31, 28) {real, imag} */,
  {32'hc6488553, 32'h00000000} /* (20, 31, 27) {real, imag} */,
  {32'hc6502876, 32'h00000000} /* (20, 31, 26) {real, imag} */,
  {32'hc645c88c, 32'h00000000} /* (20, 31, 25) {real, imag} */,
  {32'hc62f86bc, 32'h00000000} /* (20, 31, 24) {real, imag} */,
  {32'hc621fb96, 32'h00000000} /* (20, 31, 23) {real, imag} */,
  {32'hc6031936, 32'h00000000} /* (20, 31, 22) {real, imag} */,
  {32'hc5b770ba, 32'h00000000} /* (20, 31, 21) {real, imag} */,
  {32'hc54b290c, 32'h00000000} /* (20, 31, 20) {real, imag} */,
  {32'hc44a2d50, 32'h00000000} /* (20, 31, 19) {real, imag} */,
  {32'h448a75d8, 32'h00000000} /* (20, 31, 18) {real, imag} */,
  {32'h45232966, 32'h00000000} /* (20, 31, 17) {real, imag} */,
  {32'h458cf962, 32'h00000000} /* (20, 31, 16) {real, imag} */,
  {32'h45a48e53, 32'h00000000} /* (20, 31, 15) {real, imag} */,
  {32'h45bd7f3c, 32'h00000000} /* (20, 31, 14) {real, imag} */,
  {32'h45c69ee3, 32'h00000000} /* (20, 31, 13) {real, imag} */,
  {32'h45a2fabb, 32'h00000000} /* (20, 31, 12) {real, imag} */,
  {32'h45673084, 32'h00000000} /* (20, 31, 11) {real, imag} */,
  {32'h44fd6650, 32'h00000000} /* (20, 31, 10) {real, imag} */,
  {32'hc2958a40, 32'h00000000} /* (20, 31, 9) {real, imag} */,
  {32'hc526f466, 32'h00000000} /* (20, 31, 8) {real, imag} */,
  {32'hc58048bf, 32'h00000000} /* (20, 31, 7) {real, imag} */,
  {32'hc5b381c4, 32'h00000000} /* (20, 31, 6) {real, imag} */,
  {32'hc6007d34, 32'h00000000} /* (20, 31, 5) {real, imag} */,
  {32'hc60f59e8, 32'h00000000} /* (20, 31, 4) {real, imag} */,
  {32'hc61b6a1f, 32'h00000000} /* (20, 31, 3) {real, imag} */,
  {32'hc62aaa9b, 32'h00000000} /* (20, 31, 2) {real, imag} */,
  {32'hc63144a6, 32'h00000000} /* (20, 31, 1) {real, imag} */,
  {32'hc635f3b8, 32'h00000000} /* (20, 31, 0) {real, imag} */,
  {32'hc648b202, 32'h00000000} /* (20, 30, 31) {real, imag} */,
  {32'hc6548f4e, 32'h00000000} /* (20, 30, 30) {real, imag} */,
  {32'hc6587423, 32'h00000000} /* (20, 30, 29) {real, imag} */,
  {32'hc662daa6, 32'h00000000} /* (20, 30, 28) {real, imag} */,
  {32'hc65e31de, 32'h00000000} /* (20, 30, 27) {real, imag} */,
  {32'hc6470ce5, 32'h00000000} /* (20, 30, 26) {real, imag} */,
  {32'hc64b623a, 32'h00000000} /* (20, 30, 25) {real, imag} */,
  {32'hc6411353, 32'h00000000} /* (20, 30, 24) {real, imag} */,
  {32'hc62409b2, 32'h00000000} /* (20, 30, 23) {real, imag} */,
  {32'hc601d766, 32'h00000000} /* (20, 30, 22) {real, imag} */,
  {32'hc5a86a2a, 32'h00000000} /* (20, 30, 21) {real, imag} */,
  {32'hc4c14cc8, 32'h00000000} /* (20, 30, 20) {real, imag} */,
  {32'h44b6a044, 32'h00000000} /* (20, 30, 19) {real, imag} */,
  {32'h458ba64e, 32'h00000000} /* (20, 30, 18) {real, imag} */,
  {32'h45980345, 32'h00000000} /* (20, 30, 17) {real, imag} */,
  {32'h45e04026, 32'h00000000} /* (20, 30, 16) {real, imag} */,
  {32'h45e33ca4, 32'h00000000} /* (20, 30, 15) {real, imag} */,
  {32'h45f1b211, 32'h00000000} /* (20, 30, 14) {real, imag} */,
  {32'h45d4a026, 32'h00000000} /* (20, 30, 13) {real, imag} */,
  {32'h45a7b477, 32'h00000000} /* (20, 30, 12) {real, imag} */,
  {32'h45599c9a, 32'h00000000} /* (20, 30, 11) {real, imag} */,
  {32'h4351d940, 32'h00000000} /* (20, 30, 10) {real, imag} */,
  {32'hc4b4e09c, 32'h00000000} /* (20, 30, 9) {real, imag} */,
  {32'hc58ca3ea, 32'h00000000} /* (20, 30, 8) {real, imag} */,
  {32'hc5c5da2c, 32'h00000000} /* (20, 30, 7) {real, imag} */,
  {32'hc5fab0ae, 32'h00000000} /* (20, 30, 6) {real, imag} */,
  {32'hc616b21b, 32'h00000000} /* (20, 30, 5) {real, imag} */,
  {32'hc625cb78, 32'h00000000} /* (20, 30, 4) {real, imag} */,
  {32'hc633d6d6, 32'h00000000} /* (20, 30, 3) {real, imag} */,
  {32'hc631dd11, 32'h00000000} /* (20, 30, 2) {real, imag} */,
  {32'hc63a777a, 32'h00000000} /* (20, 30, 1) {real, imag} */,
  {32'hc63deca3, 32'h00000000} /* (20, 30, 0) {real, imag} */,
  {32'hc64c1110, 32'h00000000} /* (20, 29, 31) {real, imag} */,
  {32'hc654631a, 32'h00000000} /* (20, 29, 30) {real, imag} */,
  {32'hc653d4e4, 32'h00000000} /* (20, 29, 29) {real, imag} */,
  {32'hc6579556, 32'h00000000} /* (20, 29, 28) {real, imag} */,
  {32'hc658d911, 32'h00000000} /* (20, 29, 27) {real, imag} */,
  {32'hc65aeda1, 32'h00000000} /* (20, 29, 26) {real, imag} */,
  {32'hc6535d56, 32'h00000000} /* (20, 29, 25) {real, imag} */,
  {32'hc63e3e28, 32'h00000000} /* (20, 29, 24) {real, imag} */,
  {32'hc61ba390, 32'h00000000} /* (20, 29, 23) {real, imag} */,
  {32'hc6063164, 32'h00000000} /* (20, 29, 22) {real, imag} */,
  {32'hc580011e, 32'h00000000} /* (20, 29, 21) {real, imag} */,
  {32'h43809d80, 32'h00000000} /* (20, 29, 20) {real, imag} */,
  {32'h45236e26, 32'h00000000} /* (20, 29, 19) {real, imag} */,
  {32'h458ab3fe, 32'h00000000} /* (20, 29, 18) {real, imag} */,
  {32'h45cafade, 32'h00000000} /* (20, 29, 17) {real, imag} */,
  {32'h45d82824, 32'h00000000} /* (20, 29, 16) {real, imag} */,
  {32'h45ea5e48, 32'h00000000} /* (20, 29, 15) {real, imag} */,
  {32'h45f884af, 32'h00000000} /* (20, 29, 14) {real, imag} */,
  {32'h45e619a1, 32'h00000000} /* (20, 29, 13) {real, imag} */,
  {32'h45a43d64, 32'h00000000} /* (20, 29, 12) {real, imag} */,
  {32'h455b4f2c, 32'h00000000} /* (20, 29, 11) {real, imag} */,
  {32'h439f8ea0, 32'h00000000} /* (20, 29, 10) {real, imag} */,
  {32'hc53de948, 32'h00000000} /* (20, 29, 9) {real, imag} */,
  {32'hc5a955ab, 32'h00000000} /* (20, 29, 8) {real, imag} */,
  {32'hc5ed7e0b, 32'h00000000} /* (20, 29, 7) {real, imag} */,
  {32'hc60d934c, 32'h00000000} /* (20, 29, 6) {real, imag} */,
  {32'hc60e91d6, 32'h00000000} /* (20, 29, 5) {real, imag} */,
  {32'hc6258bc6, 32'h00000000} /* (20, 29, 4) {real, imag} */,
  {32'hc6308312, 32'h00000000} /* (20, 29, 3) {real, imag} */,
  {32'hc6382391, 32'h00000000} /* (20, 29, 2) {real, imag} */,
  {32'hc641355f, 32'h00000000} /* (20, 29, 1) {real, imag} */,
  {32'hc6487b46, 32'h00000000} /* (20, 29, 0) {real, imag} */,
  {32'hc6469d08, 32'h00000000} /* (20, 28, 31) {real, imag} */,
  {32'hc64ce2dc, 32'h00000000} /* (20, 28, 30) {real, imag} */,
  {32'hc64cdce7, 32'h00000000} /* (20, 28, 29) {real, imag} */,
  {32'hc65a76d8, 32'h00000000} /* (20, 28, 28) {real, imag} */,
  {32'hc6506fc9, 32'h00000000} /* (20, 28, 27) {real, imag} */,
  {32'hc6520e51, 32'h00000000} /* (20, 28, 26) {real, imag} */,
  {32'hc655b2f9, 32'h00000000} /* (20, 28, 25) {real, imag} */,
  {32'hc646b262, 32'h00000000} /* (20, 28, 24) {real, imag} */,
  {32'hc6276381, 32'h00000000} /* (20, 28, 23) {real, imag} */,
  {32'hc5ffa756, 32'h00000000} /* (20, 28, 22) {real, imag} */,
  {32'hc570f5ce, 32'h00000000} /* (20, 28, 21) {real, imag} */,
  {32'h42a71300, 32'h00000000} /* (20, 28, 20) {real, imag} */,
  {32'h452d84aa, 32'h00000000} /* (20, 28, 19) {real, imag} */,
  {32'h459c528f, 32'h00000000} /* (20, 28, 18) {real, imag} */,
  {32'h45d0e7fb, 32'h00000000} /* (20, 28, 17) {real, imag} */,
  {32'h45f2f5c5, 32'h00000000} /* (20, 28, 16) {real, imag} */,
  {32'h460933a6, 32'h00000000} /* (20, 28, 15) {real, imag} */,
  {32'h45f40a71, 32'h00000000} /* (20, 28, 14) {real, imag} */,
  {32'h45d375aa, 32'h00000000} /* (20, 28, 13) {real, imag} */,
  {32'h45bdaac4, 32'h00000000} /* (20, 28, 12) {real, imag} */,
  {32'h455ce4a4, 32'h00000000} /* (20, 28, 11) {real, imag} */,
  {32'hc2cbe500, 32'h00000000} /* (20, 28, 10) {real, imag} */,
  {32'hc5806abe, 32'h00000000} /* (20, 28, 9) {real, imag} */,
  {32'hc5eedfb4, 32'h00000000} /* (20, 28, 8) {real, imag} */,
  {32'hc605c86f, 32'h00000000} /* (20, 28, 7) {real, imag} */,
  {32'hc615ac49, 32'h00000000} /* (20, 28, 6) {real, imag} */,
  {32'hc628ee5c, 32'h00000000} /* (20, 28, 5) {real, imag} */,
  {32'hc63966d8, 32'h00000000} /* (20, 28, 4) {real, imag} */,
  {32'hc631f420, 32'h00000000} /* (20, 28, 3) {real, imag} */,
  {32'hc63cbd2a, 32'h00000000} /* (20, 28, 2) {real, imag} */,
  {32'hc64bd38c, 32'h00000000} /* (20, 28, 1) {real, imag} */,
  {32'hc64aee1a, 32'h00000000} /* (20, 28, 0) {real, imag} */,
  {32'hc6470780, 32'h00000000} /* (20, 27, 31) {real, imag} */,
  {32'hc64e81f4, 32'h00000000} /* (20, 27, 30) {real, imag} */,
  {32'hc6557146, 32'h00000000} /* (20, 27, 29) {real, imag} */,
  {32'hc66246b2, 32'h00000000} /* (20, 27, 28) {real, imag} */,
  {32'hc65528d7, 32'h00000000} /* (20, 27, 27) {real, imag} */,
  {32'hc64376ac, 32'h00000000} /* (20, 27, 26) {real, imag} */,
  {32'hc63a078e, 32'h00000000} /* (20, 27, 25) {real, imag} */,
  {32'hc64546ee, 32'h00000000} /* (20, 27, 24) {real, imag} */,
  {32'hc6289c0a, 32'h00000000} /* (20, 27, 23) {real, imag} */,
  {32'hc5cf92c8, 32'h00000000} /* (20, 27, 22) {real, imag} */,
  {32'hc5751c88, 32'h00000000} /* (20, 27, 21) {real, imag} */,
  {32'hc306ce00, 32'h00000000} /* (20, 27, 20) {real, imag} */,
  {32'h45415074, 32'h00000000} /* (20, 27, 19) {real, imag} */,
  {32'h45a28c0c, 32'h00000000} /* (20, 27, 18) {real, imag} */,
  {32'h45dd4e37, 32'h00000000} /* (20, 27, 17) {real, imag} */,
  {32'h45fd0de3, 32'h00000000} /* (20, 27, 16) {real, imag} */,
  {32'h4605e72c, 32'h00000000} /* (20, 27, 15) {real, imag} */,
  {32'h45fe2d90, 32'h00000000} /* (20, 27, 14) {real, imag} */,
  {32'h45e05e2c, 32'h00000000} /* (20, 27, 13) {real, imag} */,
  {32'h45ab8148, 32'h00000000} /* (20, 27, 12) {real, imag} */,
  {32'h452d9c04, 32'h00000000} /* (20, 27, 11) {real, imag} */,
  {32'hc49bc410, 32'h00000000} /* (20, 27, 10) {real, imag} */,
  {32'hc5a7062b, 32'h00000000} /* (20, 27, 9) {real, imag} */,
  {32'hc5e9d774, 32'h00000000} /* (20, 27, 8) {real, imag} */,
  {32'hc6114a9a, 32'h00000000} /* (20, 27, 7) {real, imag} */,
  {32'hc6283f02, 32'h00000000} /* (20, 27, 6) {real, imag} */,
  {32'hc63ee206, 32'h00000000} /* (20, 27, 5) {real, imag} */,
  {32'hc63b6f6c, 32'h00000000} /* (20, 27, 4) {real, imag} */,
  {32'hc63ffd37, 32'h00000000} /* (20, 27, 3) {real, imag} */,
  {32'hc64d0ae6, 32'h00000000} /* (20, 27, 2) {real, imag} */,
  {32'hc648c836, 32'h00000000} /* (20, 27, 1) {real, imag} */,
  {32'hc63ebad8, 32'h00000000} /* (20, 27, 0) {real, imag} */,
  {32'hc6367c01, 32'h00000000} /* (20, 26, 31) {real, imag} */,
  {32'hc63f59d6, 32'h00000000} /* (20, 26, 30) {real, imag} */,
  {32'hc64894b3, 32'h00000000} /* (20, 26, 29) {real, imag} */,
  {32'hc655bda1, 32'h00000000} /* (20, 26, 28) {real, imag} */,
  {32'hc641edca, 32'h00000000} /* (20, 26, 27) {real, imag} */,
  {32'hc63df2cb, 32'h00000000} /* (20, 26, 26) {real, imag} */,
  {32'hc638286c, 32'h00000000} /* (20, 26, 25) {real, imag} */,
  {32'hc62b6a52, 32'h00000000} /* (20, 26, 24) {real, imag} */,
  {32'hc61f328c, 32'h00000000} /* (20, 26, 23) {real, imag} */,
  {32'hc5e831b7, 32'h00000000} /* (20, 26, 22) {real, imag} */,
  {32'hc55679bb, 32'h00000000} /* (20, 26, 21) {real, imag} */,
  {32'h44540b28, 32'h00000000} /* (20, 26, 20) {real, imag} */,
  {32'h456d041e, 32'h00000000} /* (20, 26, 19) {real, imag} */,
  {32'h45bc9273, 32'h00000000} /* (20, 26, 18) {real, imag} */,
  {32'h45d86d6c, 32'h00000000} /* (20, 26, 17) {real, imag} */,
  {32'h45e48e60, 32'h00000000} /* (20, 26, 16) {real, imag} */,
  {32'h460dae57, 32'h00000000} /* (20, 26, 15) {real, imag} */,
  {32'h46065ebc, 32'h00000000} /* (20, 26, 14) {real, imag} */,
  {32'h45dc0572, 32'h00000000} /* (20, 26, 13) {real, imag} */,
  {32'h45ae1266, 32'h00000000} /* (20, 26, 12) {real, imag} */,
  {32'h451dd9bc, 32'h00000000} /* (20, 26, 11) {real, imag} */,
  {32'hc5297400, 32'h00000000} /* (20, 26, 10) {real, imag} */,
  {32'hc5a015e0, 32'h00000000} /* (20, 26, 9) {real, imag} */,
  {32'hc5f79e8f, 32'h00000000} /* (20, 26, 8) {real, imag} */,
  {32'hc6184bf6, 32'h00000000} /* (20, 26, 7) {real, imag} */,
  {32'hc6230402, 32'h00000000} /* (20, 26, 6) {real, imag} */,
  {32'hc627f6e7, 32'h00000000} /* (20, 26, 5) {real, imag} */,
  {32'hc6302db4, 32'h00000000} /* (20, 26, 4) {real, imag} */,
  {32'hc63c8658, 32'h00000000} /* (20, 26, 3) {real, imag} */,
  {32'hc6420f2a, 32'h00000000} /* (20, 26, 2) {real, imag} */,
  {32'hc640beb2, 32'h00000000} /* (20, 26, 1) {real, imag} */,
  {32'hc63f1382, 32'h00000000} /* (20, 26, 0) {real, imag} */,
  {32'hc62d1594, 32'h00000000} /* (20, 25, 31) {real, imag} */,
  {32'hc630e3ad, 32'h00000000} /* (20, 25, 30) {real, imag} */,
  {32'hc6353352, 32'h00000000} /* (20, 25, 29) {real, imag} */,
  {32'hc6423e94, 32'h00000000} /* (20, 25, 28) {real, imag} */,
  {32'hc63b3cf2, 32'h00000000} /* (20, 25, 27) {real, imag} */,
  {32'hc62c6cd8, 32'h00000000} /* (20, 25, 26) {real, imag} */,
  {32'hc62bc970, 32'h00000000} /* (20, 25, 25) {real, imag} */,
  {32'hc60ee01c, 32'h00000000} /* (20, 25, 24) {real, imag} */,
  {32'hc601383a, 32'h00000000} /* (20, 25, 23) {real, imag} */,
  {32'hc5e1aaea, 32'h00000000} /* (20, 25, 22) {real, imag} */,
  {32'hc5436fc8, 32'h00000000} /* (20, 25, 21) {real, imag} */,
  {32'h44ba0100, 32'h00000000} /* (20, 25, 20) {real, imag} */,
  {32'h4559572e, 32'h00000000} /* (20, 25, 19) {real, imag} */,
  {32'h45c71ce2, 32'h00000000} /* (20, 25, 18) {real, imag} */,
  {32'h45c81cc0, 32'h00000000} /* (20, 25, 17) {real, imag} */,
  {32'h45d78f8e, 32'h00000000} /* (20, 25, 16) {real, imag} */,
  {32'h45ecf41f, 32'h00000000} /* (20, 25, 15) {real, imag} */,
  {32'h460076b9, 32'h00000000} /* (20, 25, 14) {real, imag} */,
  {32'h45e1e273, 32'h00000000} /* (20, 25, 13) {real, imag} */,
  {32'h45a179ac, 32'h00000000} /* (20, 25, 12) {real, imag} */,
  {32'h45052322, 32'h00000000} /* (20, 25, 11) {real, imag} */,
  {32'hc51c4008, 32'h00000000} /* (20, 25, 10) {real, imag} */,
  {32'hc5ac2147, 32'h00000000} /* (20, 25, 9) {real, imag} */,
  {32'hc5fb04db, 32'h00000000} /* (20, 25, 8) {real, imag} */,
  {32'hc6167f76, 32'h00000000} /* (20, 25, 7) {real, imag} */,
  {32'hc626ac1f, 32'h00000000} /* (20, 25, 6) {real, imag} */,
  {32'hc61fd7f7, 32'h00000000} /* (20, 25, 5) {real, imag} */,
  {32'hc61dce97, 32'h00000000} /* (20, 25, 4) {real, imag} */,
  {32'hc6293f0e, 32'h00000000} /* (20, 25, 3) {real, imag} */,
  {32'hc638718f, 32'h00000000} /* (20, 25, 2) {real, imag} */,
  {32'hc62ed1a2, 32'h00000000} /* (20, 25, 1) {real, imag} */,
  {32'hc62acbc1, 32'h00000000} /* (20, 25, 0) {real, imag} */,
  {32'hc60b3bde, 32'h00000000} /* (20, 24, 31) {real, imag} */,
  {32'hc616d78b, 32'h00000000} /* (20, 24, 30) {real, imag} */,
  {32'hc616d86a, 32'h00000000} /* (20, 24, 29) {real, imag} */,
  {32'hc6174c15, 32'h00000000} /* (20, 24, 28) {real, imag} */,
  {32'hc61e674a, 32'h00000000} /* (20, 24, 27) {real, imag} */,
  {32'hc612e819, 32'h00000000} /* (20, 24, 26) {real, imag} */,
  {32'hc60fcb17, 32'h00000000} /* (20, 24, 25) {real, imag} */,
  {32'hc60a02dc, 32'h00000000} /* (20, 24, 24) {real, imag} */,
  {32'hc5f25252, 32'h00000000} /* (20, 24, 23) {real, imag} */,
  {32'hc5b2c44a, 32'h00000000} /* (20, 24, 22) {real, imag} */,
  {32'hc52dabf2, 32'h00000000} /* (20, 24, 21) {real, imag} */,
  {32'h44cc88e2, 32'h00000000} /* (20, 24, 20) {real, imag} */,
  {32'h45509e5a, 32'h00000000} /* (20, 24, 19) {real, imag} */,
  {32'h45948630, 32'h00000000} /* (20, 24, 18) {real, imag} */,
  {32'h45c9de31, 32'h00000000} /* (20, 24, 17) {real, imag} */,
  {32'h45ce2f74, 32'h00000000} /* (20, 24, 16) {real, imag} */,
  {32'h45dd503a, 32'h00000000} /* (20, 24, 15) {real, imag} */,
  {32'h45da1f3e, 32'h00000000} /* (20, 24, 14) {real, imag} */,
  {32'h45a7adaf, 32'h00000000} /* (20, 24, 13) {real, imag} */,
  {32'h4583c224, 32'h00000000} /* (20, 24, 12) {real, imag} */,
  {32'h4483b480, 32'h00000000} /* (20, 24, 11) {real, imag} */,
  {32'hc4f7d7da, 32'h00000000} /* (20, 24, 10) {real, imag} */,
  {32'hc5b52671, 32'h00000000} /* (20, 24, 9) {real, imag} */,
  {32'hc600c308, 32'h00000000} /* (20, 24, 8) {real, imag} */,
  {32'hc5fc8a6a, 32'h00000000} /* (20, 24, 7) {real, imag} */,
  {32'hc62214c7, 32'h00000000} /* (20, 24, 6) {real, imag} */,
  {32'hc60d0f72, 32'h00000000} /* (20, 24, 5) {real, imag} */,
  {32'hc6159606, 32'h00000000} /* (20, 24, 4) {real, imag} */,
  {32'hc62aec3e, 32'h00000000} /* (20, 24, 3) {real, imag} */,
  {32'hc629a1ed, 32'h00000000} /* (20, 24, 2) {real, imag} */,
  {32'hc619a56e, 32'h00000000} /* (20, 24, 1) {real, imag} */,
  {32'hc61a1e30, 32'h00000000} /* (20, 24, 0) {real, imag} */,
  {32'hc5de9229, 32'h00000000} /* (20, 23, 31) {real, imag} */,
  {32'hc5e3cc54, 32'h00000000} /* (20, 23, 30) {real, imag} */,
  {32'hc5edb3bf, 32'h00000000} /* (20, 23, 29) {real, imag} */,
  {32'hc600319e, 32'h00000000} /* (20, 23, 28) {real, imag} */,
  {32'hc601db3a, 32'h00000000} /* (20, 23, 27) {real, imag} */,
  {32'hc5e5283e, 32'h00000000} /* (20, 23, 26) {real, imag} */,
  {32'hc5e7d98e, 32'h00000000} /* (20, 23, 25) {real, imag} */,
  {32'hc5ee0bdd, 32'h00000000} /* (20, 23, 24) {real, imag} */,
  {32'hc5cd56a8, 32'h00000000} /* (20, 23, 23) {real, imag} */,
  {32'hc58e40b8, 32'h00000000} /* (20, 23, 22) {real, imag} */,
  {32'hc54e1bba, 32'h00000000} /* (20, 23, 21) {real, imag} */,
  {32'h44808700, 32'h00000000} /* (20, 23, 20) {real, imag} */,
  {32'h458303b6, 32'h00000000} /* (20, 23, 19) {real, imag} */,
  {32'h457a5384, 32'h00000000} /* (20, 23, 18) {real, imag} */,
  {32'h458cd37b, 32'h00000000} /* (20, 23, 17) {real, imag} */,
  {32'h45b5b864, 32'h00000000} /* (20, 23, 16) {real, imag} */,
  {32'h45b206c3, 32'h00000000} /* (20, 23, 15) {real, imag} */,
  {32'h45afceac, 32'h00000000} /* (20, 23, 14) {real, imag} */,
  {32'h45a0058f, 32'h00000000} /* (20, 23, 13) {real, imag} */,
  {32'h455059be, 32'h00000000} /* (20, 23, 12) {real, imag} */,
  {32'h444efc70, 32'h00000000} /* (20, 23, 11) {real, imag} */,
  {32'hc534098b, 32'h00000000} /* (20, 23, 10) {real, imag} */,
  {32'hc593c664, 32'h00000000} /* (20, 23, 9) {real, imag} */,
  {32'hc5c60483, 32'h00000000} /* (20, 23, 8) {real, imag} */,
  {32'hc5d51438, 32'h00000000} /* (20, 23, 7) {real, imag} */,
  {32'hc5f11c4c, 32'h00000000} /* (20, 23, 6) {real, imag} */,
  {32'hc5f70ca7, 32'h00000000} /* (20, 23, 5) {real, imag} */,
  {32'hc6034d87, 32'h00000000} /* (20, 23, 4) {real, imag} */,
  {32'hc60a5bab, 32'h00000000} /* (20, 23, 3) {real, imag} */,
  {32'hc6058908, 32'h00000000} /* (20, 23, 2) {real, imag} */,
  {32'hc60d2124, 32'h00000000} /* (20, 23, 1) {real, imag} */,
  {32'hc5ed1fca, 32'h00000000} /* (20, 23, 0) {real, imag} */,
  {32'hc5a12b98, 32'h00000000} /* (20, 22, 31) {real, imag} */,
  {32'hc5a10133, 32'h00000000} /* (20, 22, 30) {real, imag} */,
  {32'hc5b43f4c, 32'h00000000} /* (20, 22, 29) {real, imag} */,
  {32'hc5baeeac, 32'h00000000} /* (20, 22, 28) {real, imag} */,
  {32'hc5ad6c94, 32'h00000000} /* (20, 22, 27) {real, imag} */,
  {32'hc5a5d8aa, 32'h00000000} /* (20, 22, 26) {real, imag} */,
  {32'hc5acdfc2, 32'h00000000} /* (20, 22, 25) {real, imag} */,
  {32'hc5a43ab0, 32'h00000000} /* (20, 22, 24) {real, imag} */,
  {32'hc5852b64, 32'h00000000} /* (20, 22, 23) {real, imag} */,
  {32'hc551490e, 32'h00000000} /* (20, 22, 22) {real, imag} */,
  {32'hc4db7958, 32'h00000000} /* (20, 22, 21) {real, imag} */,
  {32'h4445e1e0, 32'h00000000} /* (20, 22, 20) {real, imag} */,
  {32'h4544a3d2, 32'h00000000} /* (20, 22, 19) {real, imag} */,
  {32'h454d95a8, 32'h00000000} /* (20, 22, 18) {real, imag} */,
  {32'h45404682, 32'h00000000} /* (20, 22, 17) {real, imag} */,
  {32'h455c98dc, 32'h00000000} /* (20, 22, 16) {real, imag} */,
  {32'h4570988f, 32'h00000000} /* (20, 22, 15) {real, imag} */,
  {32'h45850463, 32'h00000000} /* (20, 22, 14) {real, imag} */,
  {32'h4582eea2, 32'h00000000} /* (20, 22, 13) {real, imag} */,
  {32'h4558550c, 32'h00000000} /* (20, 22, 12) {real, imag} */,
  {32'h448b69ee, 32'h00000000} /* (20, 22, 11) {real, imag} */,
  {32'hc4f48a21, 32'h00000000} /* (20, 22, 10) {real, imag} */,
  {32'hc58adc24, 32'h00000000} /* (20, 22, 9) {real, imag} */,
  {32'hc591dd2a, 32'h00000000} /* (20, 22, 8) {real, imag} */,
  {32'hc5acbc80, 32'h00000000} /* (20, 22, 7) {real, imag} */,
  {32'hc5a7f647, 32'h00000000} /* (20, 22, 6) {real, imag} */,
  {32'hc5ab5c80, 32'h00000000} /* (20, 22, 5) {real, imag} */,
  {32'hc5bde08e, 32'h00000000} /* (20, 22, 4) {real, imag} */,
  {32'hc5c99793, 32'h00000000} /* (20, 22, 3) {real, imag} */,
  {32'hc5b620ac, 32'h00000000} /* (20, 22, 2) {real, imag} */,
  {32'hc5d9b1bb, 32'h00000000} /* (20, 22, 1) {real, imag} */,
  {32'hc5a8362c, 32'h00000000} /* (20, 22, 0) {real, imag} */,
  {32'hc5174d4a, 32'h00000000} /* (20, 21, 31) {real, imag} */,
  {32'hc5374609, 32'h00000000} /* (20, 21, 30) {real, imag} */,
  {32'hc532507d, 32'h00000000} /* (20, 21, 29) {real, imag} */,
  {32'hc52b73f1, 32'h00000000} /* (20, 21, 28) {real, imag} */,
  {32'hc4ee4480, 32'h00000000} /* (20, 21, 27) {real, imag} */,
  {32'hc4edf6df, 32'h00000000} /* (20, 21, 26) {real, imag} */,
  {32'hc4f6f146, 32'h00000000} /* (20, 21, 25) {real, imag} */,
  {32'hc4df53be, 32'h00000000} /* (20, 21, 24) {real, imag} */,
  {32'hc4c8e415, 32'h00000000} /* (20, 21, 23) {real, imag} */,
  {32'hc4d23bb6, 32'h00000000} /* (20, 21, 22) {real, imag} */,
  {32'h430b12a8, 32'h00000000} /* (20, 21, 21) {real, imag} */,
  {32'hc49ae354, 32'h00000000} /* (20, 21, 20) {real, imag} */,
  {32'h43668be0, 32'h00000000} /* (20, 21, 19) {real, imag} */,
  {32'h443146e2, 32'h00000000} /* (20, 21, 18) {real, imag} */,
  {32'h441daf0a, 32'h00000000} /* (20, 21, 17) {real, imag} */,
  {32'h4445643e, 32'h00000000} /* (20, 21, 16) {real, imag} */,
  {32'h44a1c51e, 32'h00000000} /* (20, 21, 15) {real, imag} */,
  {32'h45179889, 32'h00000000} /* (20, 21, 14) {real, imag} */,
  {32'h44952532, 32'h00000000} /* (20, 21, 13) {real, imag} */,
  {32'h442f0680, 32'h00000000} /* (20, 21, 12) {real, imag} */,
  {32'h44012620, 32'h00000000} /* (20, 21, 11) {real, imag} */,
  {32'hc4f64585, 32'h00000000} /* (20, 21, 10) {real, imag} */,
  {32'hc5113075, 32'h00000000} /* (20, 21, 9) {real, imag} */,
  {32'hc4b96962, 32'h00000000} /* (20, 21, 8) {real, imag} */,
  {32'hc523cc54, 32'h00000000} /* (20, 21, 7) {real, imag} */,
  {32'hc51bee73, 32'h00000000} /* (20, 21, 6) {real, imag} */,
  {32'hc4c2391f, 32'h00000000} /* (20, 21, 5) {real, imag} */,
  {32'hc53917fe, 32'h00000000} /* (20, 21, 4) {real, imag} */,
  {32'hc4d32880, 32'h00000000} /* (20, 21, 3) {real, imag} */,
  {32'hc5223e04, 32'h00000000} /* (20, 21, 2) {real, imag} */,
  {32'hc531e1ee, 32'h00000000} /* (20, 21, 1) {real, imag} */,
  {32'hc50f82da, 32'h00000000} /* (20, 21, 0) {real, imag} */,
  {32'h44f16a37, 32'h00000000} /* (20, 20, 31) {real, imag} */,
  {32'h453d7613, 32'h00000000} /* (20, 20, 30) {real, imag} */,
  {32'h4500424c, 32'h00000000} /* (20, 20, 29) {real, imag} */,
  {32'h44ea5895, 32'h00000000} /* (20, 20, 28) {real, imag} */,
  {32'h4529b5aa, 32'h00000000} /* (20, 20, 27) {real, imag} */,
  {32'h451977aa, 32'h00000000} /* (20, 20, 26) {real, imag} */,
  {32'h44fdec29, 32'h00000000} /* (20, 20, 25) {real, imag} */,
  {32'h44bc337e, 32'h00000000} /* (20, 20, 24) {real, imag} */,
  {32'h449e37c2, 32'h00000000} /* (20, 20, 23) {real, imag} */,
  {32'h44dfced4, 32'h00000000} /* (20, 20, 22) {real, imag} */,
  {32'h44921eef, 32'h00000000} /* (20, 20, 21) {real, imag} */,
  {32'hc4ac43c7, 32'h00000000} /* (20, 20, 20) {real, imag} */,
  {32'hc52a16ee, 32'h00000000} /* (20, 20, 19) {real, imag} */,
  {32'hc5141995, 32'h00000000} /* (20, 20, 18) {real, imag} */,
  {32'hc536c750, 32'h00000000} /* (20, 20, 17) {real, imag} */,
  {32'hc540098b, 32'h00000000} /* (20, 20, 16) {real, imag} */,
  {32'hc52bf835, 32'h00000000} /* (20, 20, 15) {real, imag} */,
  {32'hc50ce8b1, 32'h00000000} /* (20, 20, 14) {real, imag} */,
  {32'hc50d5b56, 32'h00000000} /* (20, 20, 13) {real, imag} */,
  {32'hc507742e, 32'h00000000} /* (20, 20, 12) {real, imag} */,
  {32'hc5165bfa, 32'h00000000} /* (20, 20, 11) {real, imag} */,
  {32'hc471bb5a, 32'h00000000} /* (20, 20, 10) {real, imag} */,
  {32'h43d55274, 32'h00000000} /* (20, 20, 9) {real, imag} */,
  {32'h43a55e1a, 32'h00000000} /* (20, 20, 8) {real, imag} */,
  {32'h442e9bb4, 32'h00000000} /* (20, 20, 7) {real, imag} */,
  {32'h450ec648, 32'h00000000} /* (20, 20, 6) {real, imag} */,
  {32'h450aedea, 32'h00000000} /* (20, 20, 5) {real, imag} */,
  {32'h4492ac63, 32'h00000000} /* (20, 20, 4) {real, imag} */,
  {32'h44d1d109, 32'h00000000} /* (20, 20, 3) {real, imag} */,
  {32'h44ebec06, 32'h00000000} /* (20, 20, 2) {real, imag} */,
  {32'h44b0e7b8, 32'h00000000} /* (20, 20, 1) {real, imag} */,
  {32'h44812692, 32'h00000000} /* (20, 20, 0) {real, imag} */,
  {32'h458de30d, 32'h00000000} /* (20, 19, 31) {real, imag} */,
  {32'h459bb0bc, 32'h00000000} /* (20, 19, 30) {real, imag} */,
  {32'h45b09162, 32'h00000000} /* (20, 19, 29) {real, imag} */,
  {32'h45b146d0, 32'h00000000} /* (20, 19, 28) {real, imag} */,
  {32'h45a3352e, 32'h00000000} /* (20, 19, 27) {real, imag} */,
  {32'h45947273, 32'h00000000} /* (20, 19, 26) {real, imag} */,
  {32'h459a9a90, 32'h00000000} /* (20, 19, 25) {real, imag} */,
  {32'h459b5f9b, 32'h00000000} /* (20, 19, 24) {real, imag} */,
  {32'h4597cb0b, 32'h00000000} /* (20, 19, 23) {real, imag} */,
  {32'h4535a354, 32'h00000000} /* (20, 19, 22) {real, imag} */,
  {32'h43e7fd7c, 32'h00000000} /* (20, 19, 21) {real, imag} */,
  {32'hc500516c, 32'h00000000} /* (20, 19, 20) {real, imag} */,
  {32'hc56712b5, 32'h00000000} /* (20, 19, 19) {real, imag} */,
  {32'hc5a1c31d, 32'h00000000} /* (20, 19, 18) {real, imag} */,
  {32'hc5afb593, 32'h00000000} /* (20, 19, 17) {real, imag} */,
  {32'hc5b9b5bc, 32'h00000000} /* (20, 19, 16) {real, imag} */,
  {32'hc5c28463, 32'h00000000} /* (20, 19, 15) {real, imag} */,
  {32'hc5aba5f0, 32'h00000000} /* (20, 19, 14) {real, imag} */,
  {32'hc59890bc, 32'h00000000} /* (20, 19, 13) {real, imag} */,
  {32'hc541fe20, 32'h00000000} /* (20, 19, 12) {real, imag} */,
  {32'hc53a61a0, 32'h00000000} /* (20, 19, 11) {real, imag} */,
  {32'hc3c089d0, 32'h00000000} /* (20, 19, 10) {real, imag} */,
  {32'h4517b154, 32'h00000000} /* (20, 19, 9) {real, imag} */,
  {32'h450bc822, 32'h00000000} /* (20, 19, 8) {real, imag} */,
  {32'h45336b02, 32'h00000000} /* (20, 19, 7) {real, imag} */,
  {32'h456a4ccc, 32'h00000000} /* (20, 19, 6) {real, imag} */,
  {32'h45755e18, 32'h00000000} /* (20, 19, 5) {real, imag} */,
  {32'h45971cad, 32'h00000000} /* (20, 19, 4) {real, imag} */,
  {32'h458e1595, 32'h00000000} /* (20, 19, 3) {real, imag} */,
  {32'h4597518f, 32'h00000000} /* (20, 19, 2) {real, imag} */,
  {32'h45b54a61, 32'h00000000} /* (20, 19, 1) {real, imag} */,
  {32'h4590897e, 32'h00000000} /* (20, 19, 0) {real, imag} */,
  {32'h45b4458a, 32'h00000000} /* (20, 18, 31) {real, imag} */,
  {32'h45dd2faa, 32'h00000000} /* (20, 18, 30) {real, imag} */,
  {32'h45ee661c, 32'h00000000} /* (20, 18, 29) {real, imag} */,
  {32'h45e55896, 32'h00000000} /* (20, 18, 28) {real, imag} */,
  {32'h45e998be, 32'h00000000} /* (20, 18, 27) {real, imag} */,
  {32'h45d44a34, 32'h00000000} /* (20, 18, 26) {real, imag} */,
  {32'h45c2d3ed, 32'h00000000} /* (20, 18, 25) {real, imag} */,
  {32'h45d63952, 32'h00000000} /* (20, 18, 24) {real, imag} */,
  {32'h45b9a938, 32'h00000000} /* (20, 18, 23) {real, imag} */,
  {32'h453eafce, 32'h00000000} /* (20, 18, 22) {real, imag} */,
  {32'h45047b12, 32'h00000000} /* (20, 18, 21) {real, imag} */,
  {32'hc50a5e4e, 32'h00000000} /* (20, 18, 20) {real, imag} */,
  {32'hc5909b58, 32'h00000000} /* (20, 18, 19) {real, imag} */,
  {32'hc5be783b, 32'h00000000} /* (20, 18, 18) {real, imag} */,
  {32'hc5ec0c18, 32'h00000000} /* (20, 18, 17) {real, imag} */,
  {32'hc60008eb, 32'h00000000} /* (20, 18, 16) {real, imag} */,
  {32'hc5e631f0, 32'h00000000} /* (20, 18, 15) {real, imag} */,
  {32'hc5ce8882, 32'h00000000} /* (20, 18, 14) {real, imag} */,
  {32'hc5a174c0, 32'h00000000} /* (20, 18, 13) {real, imag} */,
  {32'hc58c4ba2, 32'h00000000} /* (20, 18, 12) {real, imag} */,
  {32'hc5147c49, 32'h00000000} /* (20, 18, 11) {real, imag} */,
  {32'h44854848, 32'h00000000} /* (20, 18, 10) {real, imag} */,
  {32'h45126796, 32'h00000000} /* (20, 18, 9) {real, imag} */,
  {32'h458f21de, 32'h00000000} /* (20, 18, 8) {real, imag} */,
  {32'h459433da, 32'h00000000} /* (20, 18, 7) {real, imag} */,
  {32'h45b32079, 32'h00000000} /* (20, 18, 6) {real, imag} */,
  {32'h45e90a07, 32'h00000000} /* (20, 18, 5) {real, imag} */,
  {32'h45e1bf4b, 32'h00000000} /* (20, 18, 4) {real, imag} */,
  {32'h45e18afc, 32'h00000000} /* (20, 18, 3) {real, imag} */,
  {32'h45dd3f9d, 32'h00000000} /* (20, 18, 2) {real, imag} */,
  {32'h45fa08dc, 32'h00000000} /* (20, 18, 1) {real, imag} */,
  {32'h46040937, 32'h00000000} /* (20, 18, 0) {real, imag} */,
  {32'h45fb672b, 32'h00000000} /* (20, 17, 31) {real, imag} */,
  {32'h45ffae80, 32'h00000000} /* (20, 17, 30) {real, imag} */,
  {32'h46030032, 32'h00000000} /* (20, 17, 29) {real, imag} */,
  {32'h460cc5be, 32'h00000000} /* (20, 17, 28) {real, imag} */,
  {32'h46063506, 32'h00000000} /* (20, 17, 27) {real, imag} */,
  {32'h460dc230, 32'h00000000} /* (20, 17, 26) {real, imag} */,
  {32'h45faa76f, 32'h00000000} /* (20, 17, 25) {real, imag} */,
  {32'h45e9057d, 32'h00000000} /* (20, 17, 24) {real, imag} */,
  {32'h45adb01f, 32'h00000000} /* (20, 17, 23) {real, imag} */,
  {32'h45682b9e, 32'h00000000} /* (20, 17, 22) {real, imag} */,
  {32'h43e8e0f0, 32'h00000000} /* (20, 17, 21) {real, imag} */,
  {32'hc506c29f, 32'h00000000} /* (20, 17, 20) {real, imag} */,
  {32'hc5a61b3a, 32'h00000000} /* (20, 17, 19) {real, imag} */,
  {32'hc5db53a0, 32'h00000000} /* (20, 17, 18) {real, imag} */,
  {32'hc5d3c7f6, 32'h00000000} /* (20, 17, 17) {real, imag} */,
  {32'hc60c2a4a, 32'h00000000} /* (20, 17, 16) {real, imag} */,
  {32'hc605e284, 32'h00000000} /* (20, 17, 15) {real, imag} */,
  {32'hc5e40bdc, 32'h00000000} /* (20, 17, 14) {real, imag} */,
  {32'hc5b31b8b, 32'h00000000} /* (20, 17, 13) {real, imag} */,
  {32'hc588d4a4, 32'h00000000} /* (20, 17, 12) {real, imag} */,
  {32'hc52cf182, 32'h00000000} /* (20, 17, 11) {real, imag} */,
  {32'h43590e60, 32'h00000000} /* (20, 17, 10) {real, imag} */,
  {32'h456379ae, 32'h00000000} /* (20, 17, 9) {real, imag} */,
  {32'h45a70e7f, 32'h00000000} /* (20, 17, 8) {real, imag} */,
  {32'h45c37b19, 32'h00000000} /* (20, 17, 7) {real, imag} */,
  {32'h45e02d29, 32'h00000000} /* (20, 17, 6) {real, imag} */,
  {32'h46079224, 32'h00000000} /* (20, 17, 5) {real, imag} */,
  {32'h4611962b, 32'h00000000} /* (20, 17, 4) {real, imag} */,
  {32'h46050044, 32'h00000000} /* (20, 17, 3) {real, imag} */,
  {32'h460e988f, 32'h00000000} /* (20, 17, 2) {real, imag} */,
  {32'h461e9287, 32'h00000000} /* (20, 17, 1) {real, imag} */,
  {32'h45f8e480, 32'h00000000} /* (20, 17, 0) {real, imag} */,
  {32'h46078cd2, 32'h00000000} /* (20, 16, 31) {real, imag} */,
  {32'h460d15b3, 32'h00000000} /* (20, 16, 30) {real, imag} */,
  {32'h460d679b, 32'h00000000} /* (20, 16, 29) {real, imag} */,
  {32'h4613e49e, 32'h00000000} /* (20, 16, 28) {real, imag} */,
  {32'h4617a55b, 32'h00000000} /* (20, 16, 27) {real, imag} */,
  {32'h46090841, 32'h00000000} /* (20, 16, 26) {real, imag} */,
  {32'h460bb323, 32'h00000000} /* (20, 16, 25) {real, imag} */,
  {32'h45efe65a, 32'h00000000} /* (20, 16, 24) {real, imag} */,
  {32'h45b3ee36, 32'h00000000} /* (20, 16, 23) {real, imag} */,
  {32'h4552ca5c, 32'h00000000} /* (20, 16, 22) {real, imag} */,
  {32'h4340d6e0, 32'h00000000} /* (20, 16, 21) {real, imag} */,
  {32'hc53af5e1, 32'h00000000} /* (20, 16, 20) {real, imag} */,
  {32'hc5a17f39, 32'h00000000} /* (20, 16, 19) {real, imag} */,
  {32'hc5d2739c, 32'h00000000} /* (20, 16, 18) {real, imag} */,
  {32'hc5f604a7, 32'h00000000} /* (20, 16, 17) {real, imag} */,
  {32'hc6057672, 32'h00000000} /* (20, 16, 16) {real, imag} */,
  {32'hc5ec96fc, 32'h00000000} /* (20, 16, 15) {real, imag} */,
  {32'hc5f40066, 32'h00000000} /* (20, 16, 14) {real, imag} */,
  {32'hc5d83b25, 32'h00000000} /* (20, 16, 13) {real, imag} */,
  {32'hc5a9ca46, 32'h00000000} /* (20, 16, 12) {real, imag} */,
  {32'hc54b1a4c, 32'h00000000} /* (20, 16, 11) {real, imag} */,
  {32'h444ce0cc, 32'h00000000} /* (20, 16, 10) {real, imag} */,
  {32'h4586eb80, 32'h00000000} /* (20, 16, 9) {real, imag} */,
  {32'h45c83c12, 32'h00000000} /* (20, 16, 8) {real, imag} */,
  {32'h45cd901e, 32'h00000000} /* (20, 16, 7) {real, imag} */,
  {32'h45f84346, 32'h00000000} /* (20, 16, 6) {real, imag} */,
  {32'h460ed10c, 32'h00000000} /* (20, 16, 5) {real, imag} */,
  {32'h46133a1c, 32'h00000000} /* (20, 16, 4) {real, imag} */,
  {32'h46174348, 32'h00000000} /* (20, 16, 3) {real, imag} */,
  {32'h4616c6fe, 32'h00000000} /* (20, 16, 2) {real, imag} */,
  {32'h460bc0ca, 32'h00000000} /* (20, 16, 1) {real, imag} */,
  {32'h46105b0c, 32'h00000000} /* (20, 16, 0) {real, imag} */,
  {32'h46109c32, 32'h00000000} /* (20, 15, 31) {real, imag} */,
  {32'h4617f5fd, 32'h00000000} /* (20, 15, 30) {real, imag} */,
  {32'h461e91d6, 32'h00000000} /* (20, 15, 29) {real, imag} */,
  {32'h460b0aae, 32'h00000000} /* (20, 15, 28) {real, imag} */,
  {32'h4607f714, 32'h00000000} /* (20, 15, 27) {real, imag} */,
  {32'h460a8b81, 32'h00000000} /* (20, 15, 26) {real, imag} */,
  {32'h45f810e3, 32'h00000000} /* (20, 15, 25) {real, imag} */,
  {32'h45df4bf9, 32'h00000000} /* (20, 15, 24) {real, imag} */,
  {32'h45a6955e, 32'h00000000} /* (20, 15, 23) {real, imag} */,
  {32'h45701c40, 32'h00000000} /* (20, 15, 22) {real, imag} */,
  {32'h44bbb54c, 32'h00000000} /* (20, 15, 21) {real, imag} */,
  {32'hc534df28, 32'h00000000} /* (20, 15, 20) {real, imag} */,
  {32'hc5cbe282, 32'h00000000} /* (20, 15, 19) {real, imag} */,
  {32'hc5c616ea, 32'h00000000} /* (20, 15, 18) {real, imag} */,
  {32'hc5f6316a, 32'h00000000} /* (20, 15, 17) {real, imag} */,
  {32'hc600dc1c, 32'h00000000} /* (20, 15, 16) {real, imag} */,
  {32'hc6012bee, 32'h00000000} /* (20, 15, 15) {real, imag} */,
  {32'hc5e1d516, 32'h00000000} /* (20, 15, 14) {real, imag} */,
  {32'hc5e54bdc, 32'h00000000} /* (20, 15, 13) {real, imag} */,
  {32'hc5bd5ce3, 32'h00000000} /* (20, 15, 12) {real, imag} */,
  {32'hc5636da2, 32'h00000000} /* (20, 15, 11) {real, imag} */,
  {32'h43e449e0, 32'h00000000} /* (20, 15, 10) {real, imag} */,
  {32'h4576b1b2, 32'h00000000} /* (20, 15, 9) {real, imag} */,
  {32'h45b1087f, 32'h00000000} /* (20, 15, 8) {real, imag} */,
  {32'h45e8337e, 32'h00000000} /* (20, 15, 7) {real, imag} */,
  {32'h45faa8b4, 32'h00000000} /* (20, 15, 6) {real, imag} */,
  {32'h46156ae6, 32'h00000000} /* (20, 15, 5) {real, imag} */,
  {32'h46136e44, 32'h00000000} /* (20, 15, 4) {real, imag} */,
  {32'h462981fd, 32'h00000000} /* (20, 15, 3) {real, imag} */,
  {32'h461c8490, 32'h00000000} /* (20, 15, 2) {real, imag} */,
  {32'h46032d5f, 32'h00000000} /* (20, 15, 1) {real, imag} */,
  {32'h45fe9a84, 32'h00000000} /* (20, 15, 0) {real, imag} */,
  {32'h45f1f93d, 32'h00000000} /* (20, 14, 31) {real, imag} */,
  {32'h45fb1404, 32'h00000000} /* (20, 14, 30) {real, imag} */,
  {32'h46015735, 32'h00000000} /* (20, 14, 29) {real, imag} */,
  {32'h4608eb50, 32'h00000000} /* (20, 14, 28) {real, imag} */,
  {32'h45f3af2b, 32'h00000000} /* (20, 14, 27) {real, imag} */,
  {32'h45f9bf8f, 32'h00000000} /* (20, 14, 26) {real, imag} */,
  {32'h45e61343, 32'h00000000} /* (20, 14, 25) {real, imag} */,
  {32'h45d57132, 32'h00000000} /* (20, 14, 24) {real, imag} */,
  {32'h45b09832, 32'h00000000} /* (20, 14, 23) {real, imag} */,
  {32'h45745817, 32'h00000000} /* (20, 14, 22) {real, imag} */,
  {32'h44b49d9c, 32'h00000000} /* (20, 14, 21) {real, imag} */,
  {32'hc54f313d, 32'h00000000} /* (20, 14, 20) {real, imag} */,
  {32'hc5974681, 32'h00000000} /* (20, 14, 19) {real, imag} */,
  {32'hc5ba3cf6, 32'h00000000} /* (20, 14, 18) {real, imag} */,
  {32'hc5d9ee60, 32'h00000000} /* (20, 14, 17) {real, imag} */,
  {32'hc5e51fe3, 32'h00000000} /* (20, 14, 16) {real, imag} */,
  {32'hc5f49a47, 32'h00000000} /* (20, 14, 15) {real, imag} */,
  {32'hc5e55942, 32'h00000000} /* (20, 14, 14) {real, imag} */,
  {32'hc5c29e1e, 32'h00000000} /* (20, 14, 13) {real, imag} */,
  {32'hc5aac2c8, 32'h00000000} /* (20, 14, 12) {real, imag} */,
  {32'hc506b8b6, 32'h00000000} /* (20, 14, 11) {real, imag} */,
  {32'h44682f88, 32'h00000000} /* (20, 14, 10) {real, imag} */,
  {32'h45886159, 32'h00000000} /* (20, 14, 9) {real, imag} */,
  {32'h45d0fcb2, 32'h00000000} /* (20, 14, 8) {real, imag} */,
  {32'h45e5af96, 32'h00000000} /* (20, 14, 7) {real, imag} */,
  {32'h45f89ce0, 32'h00000000} /* (20, 14, 6) {real, imag} */,
  {32'h45fb91a5, 32'h00000000} /* (20, 14, 5) {real, imag} */,
  {32'h45fcce2a, 32'h00000000} /* (20, 14, 4) {real, imag} */,
  {32'h45fdb81f, 32'h00000000} /* (20, 14, 3) {real, imag} */,
  {32'h460006ed, 32'h00000000} /* (20, 14, 2) {real, imag} */,
  {32'h46056f8f, 32'h00000000} /* (20, 14, 1) {real, imag} */,
  {32'h45df4dcb, 32'h00000000} /* (20, 14, 0) {real, imag} */,
  {32'h45b6c588, 32'h00000000} /* (20, 13, 31) {real, imag} */,
  {32'h45c59cc1, 32'h00000000} /* (20, 13, 30) {real, imag} */,
  {32'h45daa441, 32'h00000000} /* (20, 13, 29) {real, imag} */,
  {32'h45d89808, 32'h00000000} /* (20, 13, 28) {real, imag} */,
  {32'h45e991a0, 32'h00000000} /* (20, 13, 27) {real, imag} */,
  {32'h45d0c156, 32'h00000000} /* (20, 13, 26) {real, imag} */,
  {32'h45a4d840, 32'h00000000} /* (20, 13, 25) {real, imag} */,
  {32'h45b02494, 32'h00000000} /* (20, 13, 24) {real, imag} */,
  {32'h459a816a, 32'h00000000} /* (20, 13, 23) {real, imag} */,
  {32'h4558e342, 32'h00000000} /* (20, 13, 22) {real, imag} */,
  {32'h448ee316, 32'h00000000} /* (20, 13, 21) {real, imag} */,
  {32'hc5078e86, 32'h00000000} /* (20, 13, 20) {real, imag} */,
  {32'hc57da880, 32'h00000000} /* (20, 13, 19) {real, imag} */,
  {32'hc59228c7, 32'h00000000} /* (20, 13, 18) {real, imag} */,
  {32'hc5bfea4a, 32'h00000000} /* (20, 13, 17) {real, imag} */,
  {32'hc5bf7dc8, 32'h00000000} /* (20, 13, 16) {real, imag} */,
  {32'hc5b86e08, 32'h00000000} /* (20, 13, 15) {real, imag} */,
  {32'hc5ccfa47, 32'h00000000} /* (20, 13, 14) {real, imag} */,
  {32'hc5bfbb31, 32'h00000000} /* (20, 13, 13) {real, imag} */,
  {32'hc58be30a, 32'h00000000} /* (20, 13, 12) {real, imag} */,
  {32'hc4de8180, 32'h00000000} /* (20, 13, 11) {real, imag} */,
  {32'h449424a6, 32'h00000000} /* (20, 13, 10) {real, imag} */,
  {32'h4592d480, 32'h00000000} /* (20, 13, 9) {real, imag} */,
  {32'h45ce4c68, 32'h00000000} /* (20, 13, 8) {real, imag} */,
  {32'h45bffa84, 32'h00000000} /* (20, 13, 7) {real, imag} */,
  {32'h45d3ba4d, 32'h00000000} /* (20, 13, 6) {real, imag} */,
  {32'h45de48a6, 32'h00000000} /* (20, 13, 5) {real, imag} */,
  {32'h45e6e081, 32'h00000000} /* (20, 13, 4) {real, imag} */,
  {32'h45cc6c2e, 32'h00000000} /* (20, 13, 3) {real, imag} */,
  {32'h45d4cd4f, 32'h00000000} /* (20, 13, 2) {real, imag} */,
  {32'h45de4cc2, 32'h00000000} /* (20, 13, 1) {real, imag} */,
  {32'h45c95c30, 32'h00000000} /* (20, 13, 0) {real, imag} */,
  {32'h4587a973, 32'h00000000} /* (20, 12, 31) {real, imag} */,
  {32'h4593c4b8, 32'h00000000} /* (20, 12, 30) {real, imag} */,
  {32'h457a8097, 32'h00000000} /* (20, 12, 29) {real, imag} */,
  {32'h4580b49e, 32'h00000000} /* (20, 12, 28) {real, imag} */,
  {32'h458be3d0, 32'h00000000} /* (20, 12, 27) {real, imag} */,
  {32'h458375d7, 32'h00000000} /* (20, 12, 26) {real, imag} */,
  {32'h454e3787, 32'h00000000} /* (20, 12, 25) {real, imag} */,
  {32'h452f117a, 32'h00000000} /* (20, 12, 24) {real, imag} */,
  {32'h4542a153, 32'h00000000} /* (20, 12, 23) {real, imag} */,
  {32'h452c7737, 32'h00000000} /* (20, 12, 22) {real, imag} */,
  {32'h449c5cc4, 32'h00000000} /* (20, 12, 21) {real, imag} */,
  {32'hc4f2d5e4, 32'h00000000} /* (20, 12, 20) {real, imag} */,
  {32'hc55a00f1, 32'h00000000} /* (20, 12, 19) {real, imag} */,
  {32'hc57a47a8, 32'h00000000} /* (20, 12, 18) {real, imag} */,
  {32'hc57fb815, 32'h00000000} /* (20, 12, 17) {real, imag} */,
  {32'hc58ab4fe, 32'h00000000} /* (20, 12, 16) {real, imag} */,
  {32'hc59c26e7, 32'h00000000} /* (20, 12, 15) {real, imag} */,
  {32'hc5a39992, 32'h00000000} /* (20, 12, 14) {real, imag} */,
  {32'hc5a37d98, 32'h00000000} /* (20, 12, 13) {real, imag} */,
  {32'hc5046ed2, 32'h00000000} /* (20, 12, 12) {real, imag} */,
  {32'hc429107c, 32'h00000000} /* (20, 12, 11) {real, imag} */,
  {32'h44f494b4, 32'h00000000} /* (20, 12, 10) {real, imag} */,
  {32'h458b6b11, 32'h00000000} /* (20, 12, 9) {real, imag} */,
  {32'h45a43f7d, 32'h00000000} /* (20, 12, 8) {real, imag} */,
  {32'h45b3111a, 32'h00000000} /* (20, 12, 7) {real, imag} */,
  {32'h45909995, 32'h00000000} /* (20, 12, 6) {real, imag} */,
  {32'h45963632, 32'h00000000} /* (20, 12, 5) {real, imag} */,
  {32'h45b55af2, 32'h00000000} /* (20, 12, 4) {real, imag} */,
  {32'h45af1996, 32'h00000000} /* (20, 12, 3) {real, imag} */,
  {32'h459ed8c6, 32'h00000000} /* (20, 12, 2) {real, imag} */,
  {32'h458e4584, 32'h00000000} /* (20, 12, 1) {real, imag} */,
  {32'h4574f574, 32'h00000000} /* (20, 12, 0) {real, imag} */,
  {32'h44b03379, 32'h00000000} /* (20, 11, 31) {real, imag} */,
  {32'h450c051c, 32'h00000000} /* (20, 11, 30) {real, imag} */,
  {32'h44cc3e56, 32'h00000000} /* (20, 11, 29) {real, imag} */,
  {32'h44fd3978, 32'h00000000} /* (20, 11, 28) {real, imag} */,
  {32'h4517f3da, 32'h00000000} /* (20, 11, 27) {real, imag} */,
  {32'h44baab4d, 32'h00000000} /* (20, 11, 26) {real, imag} */,
  {32'h43fbae14, 32'h00000000} /* (20, 11, 25) {real, imag} */,
  {32'h44929f6b, 32'h00000000} /* (20, 11, 24) {real, imag} */,
  {32'h44c08a15, 32'h00000000} /* (20, 11, 23) {real, imag} */,
  {32'h44331424, 32'h00000000} /* (20, 11, 22) {real, imag} */,
  {32'hc43aafaa, 32'h00000000} /* (20, 11, 21) {real, imag} */,
  {32'hc505c424, 32'h00000000} /* (20, 11, 20) {real, imag} */,
  {32'hc504b95d, 32'h00000000} /* (20, 11, 19) {real, imag} */,
  {32'hc53421f2, 32'h00000000} /* (20, 11, 18) {real, imag} */,
  {32'hc52ca658, 32'h00000000} /* (20, 11, 17) {real, imag} */,
  {32'hc4f3a91e, 32'h00000000} /* (20, 11, 16) {real, imag} */,
  {32'hc4fc308d, 32'h00000000} /* (20, 11, 15) {real, imag} */,
  {32'hc4c6d741, 32'h00000000} /* (20, 11, 14) {real, imag} */,
  {32'hc46f2944, 32'h00000000} /* (20, 11, 13) {real, imag} */,
  {32'hc4afb3f2, 32'h00000000} /* (20, 11, 12) {real, imag} */,
  {32'h440b221e, 32'h00000000} /* (20, 11, 11) {real, imag} */,
  {32'h451319d0, 32'h00000000} /* (20, 11, 10) {real, imag} */,
  {32'h455087ca, 32'h00000000} /* (20, 11, 9) {real, imag} */,
  {32'h4553d6c0, 32'h00000000} /* (20, 11, 8) {real, imag} */,
  {32'h454478ea, 32'h00000000} /* (20, 11, 7) {real, imag} */,
  {32'h455591b5, 32'h00000000} /* (20, 11, 6) {real, imag} */,
  {32'h450a9528, 32'h00000000} /* (20, 11, 5) {real, imag} */,
  {32'h44e54e81, 32'h00000000} /* (20, 11, 4) {real, imag} */,
  {32'h45212bf9, 32'h00000000} /* (20, 11, 3) {real, imag} */,
  {32'h45186aa2, 32'h00000000} /* (20, 11, 2) {real, imag} */,
  {32'h44d4e650, 32'h00000000} /* (20, 11, 1) {real, imag} */,
  {32'h448069fa, 32'h00000000} /* (20, 11, 0) {real, imag} */,
  {32'hc4e3f825, 32'h00000000} /* (20, 10, 31) {real, imag} */,
  {32'hc50b0e8f, 32'h00000000} /* (20, 10, 30) {real, imag} */,
  {32'hc50d0f9e, 32'h00000000} /* (20, 10, 29) {real, imag} */,
  {32'hc5188937, 32'h00000000} /* (20, 10, 28) {real, imag} */,
  {32'hc53d3bc3, 32'h00000000} /* (20, 10, 27) {real, imag} */,
  {32'hc54cc4fa, 32'h00000000} /* (20, 10, 26) {real, imag} */,
  {32'hc51dc334, 32'h00000000} /* (20, 10, 25) {real, imag} */,
  {32'hc515bd0d, 32'h00000000} /* (20, 10, 24) {real, imag} */,
  {32'hc51bb69c, 32'h00000000} /* (20, 10, 23) {real, imag} */,
  {32'hc5313909, 32'h00000000} /* (20, 10, 22) {real, imag} */,
  {32'hc4c84970, 32'h00000000} /* (20, 10, 21) {real, imag} */,
  {32'hc481d7ae, 32'h00000000} /* (20, 10, 20) {real, imag} */,
  {32'hc3bae3e0, 32'h00000000} /* (20, 10, 19) {real, imag} */,
  {32'h43337738, 32'h00000000} /* (20, 10, 18) {real, imag} */,
  {32'h43d2a6f2, 32'h00000000} /* (20, 10, 17) {real, imag} */,
  {32'h44f8da45, 32'h00000000} /* (20, 10, 16) {real, imag} */,
  {32'h4501d2da, 32'h00000000} /* (20, 10, 15) {real, imag} */,
  {32'h44aa61be, 32'h00000000} /* (20, 10, 14) {real, imag} */,
  {32'h44cdcb58, 32'h00000000} /* (20, 10, 13) {real, imag} */,
  {32'h44859b24, 32'h00000000} /* (20, 10, 12) {real, imag} */,
  {32'h44a08762, 32'h00000000} /* (20, 10, 11) {real, imag} */,
  {32'h44e367d5, 32'h00000000} /* (20, 10, 10) {real, imag} */,
  {32'h43100cf8, 32'h00000000} /* (20, 10, 9) {real, imag} */,
  {32'h436047c0, 32'h00000000} /* (20, 10, 8) {real, imag} */,
  {32'h4430a0eb, 32'h00000000} /* (20, 10, 7) {real, imag} */,
  {32'hc481a5ba, 32'h00000000} /* (20, 10, 6) {real, imag} */,
  {32'hc4a5d67c, 32'h00000000} /* (20, 10, 5) {real, imag} */,
  {32'hc4ab38d4, 32'h00000000} /* (20, 10, 4) {real, imag} */,
  {32'hc501ea90, 32'h00000000} /* (20, 10, 3) {real, imag} */,
  {32'hc54240fe, 32'h00000000} /* (20, 10, 2) {real, imag} */,
  {32'hc4c21ae4, 32'h00000000} /* (20, 10, 1) {real, imag} */,
  {32'hc4e3d37b, 32'h00000000} /* (20, 10, 0) {real, imag} */,
  {32'hc59c560e, 32'h00000000} /* (20, 9, 31) {real, imag} */,
  {32'hc5af70fa, 32'h00000000} /* (20, 9, 30) {real, imag} */,
  {32'hc5ac1399, 32'h00000000} /* (20, 9, 29) {real, imag} */,
  {32'hc5c91975, 32'h00000000} /* (20, 9, 28) {real, imag} */,
  {32'hc5d838cd, 32'h00000000} /* (20, 9, 27) {real, imag} */,
  {32'hc5ca04b2, 32'h00000000} /* (20, 9, 26) {real, imag} */,
  {32'hc5afea3f, 32'h00000000} /* (20, 9, 25) {real, imag} */,
  {32'hc5bcdb63, 32'h00000000} /* (20, 9, 24) {real, imag} */,
  {32'hc5a1400a, 32'h00000000} /* (20, 9, 23) {real, imag} */,
  {32'hc58c7c52, 32'h00000000} /* (20, 9, 22) {real, imag} */,
  {32'hc55cfa46, 32'h00000000} /* (20, 9, 21) {real, imag} */,
  {32'hc42bbc46, 32'h00000000} /* (20, 9, 20) {real, imag} */,
  {32'h4468dc3c, 32'h00000000} /* (20, 9, 19) {real, imag} */,
  {32'h451068ae, 32'h00000000} /* (20, 9, 18) {real, imag} */,
  {32'h4520d76f, 32'h00000000} /* (20, 9, 17) {real, imag} */,
  {32'h455b9790, 32'h00000000} /* (20, 9, 16) {real, imag} */,
  {32'h45883468, 32'h00000000} /* (20, 9, 15) {real, imag} */,
  {32'h45958842, 32'h00000000} /* (20, 9, 14) {real, imag} */,
  {32'h455905ae, 32'h00000000} /* (20, 9, 13) {real, imag} */,
  {32'h45663e42, 32'h00000000} /* (20, 9, 12) {real, imag} */,
  {32'h450ff77e, 32'h00000000} /* (20, 9, 11) {real, imag} */,
  {32'h4407a754, 32'h00000000} /* (20, 9, 10) {real, imag} */,
  {32'hc48c589c, 32'h00000000} /* (20, 9, 9) {real, imag} */,
  {32'hc5013faa, 32'h00000000} /* (20, 9, 8) {real, imag} */,
  {32'hc50b78f8, 32'h00000000} /* (20, 9, 7) {real, imag} */,
  {32'hc54f0f2d, 32'h00000000} /* (20, 9, 6) {real, imag} */,
  {32'hc579982e, 32'h00000000} /* (20, 9, 5) {real, imag} */,
  {32'hc57845c2, 32'h00000000} /* (20, 9, 4) {real, imag} */,
  {32'hc58dba4a, 32'h00000000} /* (20, 9, 3) {real, imag} */,
  {32'hc5915b54, 32'h00000000} /* (20, 9, 2) {real, imag} */,
  {32'hc59e20c6, 32'h00000000} /* (20, 9, 1) {real, imag} */,
  {32'hc5a3abce, 32'h00000000} /* (20, 9, 0) {real, imag} */,
  {32'hc5f14268, 32'h00000000} /* (20, 8, 31) {real, imag} */,
  {32'hc5f6da24, 32'h00000000} /* (20, 8, 30) {real, imag} */,
  {32'hc60a915e, 32'h00000000} /* (20, 8, 29) {real, imag} */,
  {32'hc60c862b, 32'h00000000} /* (20, 8, 28) {real, imag} */,
  {32'hc6071216, 32'h00000000} /* (20, 8, 27) {real, imag} */,
  {32'hc616019a, 32'h00000000} /* (20, 8, 26) {real, imag} */,
  {32'hc60cd764, 32'h00000000} /* (20, 8, 25) {real, imag} */,
  {32'hc5e9ce32, 32'h00000000} /* (20, 8, 24) {real, imag} */,
  {32'hc5eb260f, 32'h00000000} /* (20, 8, 23) {real, imag} */,
  {32'hc5e0ed9c, 32'h00000000} /* (20, 8, 22) {real, imag} */,
  {32'hc5a774ee, 32'h00000000} /* (20, 8, 21) {real, imag} */,
  {32'hc481de44, 32'h00000000} /* (20, 8, 20) {real, imag} */,
  {32'h449e54f8, 32'h00000000} /* (20, 8, 19) {real, imag} */,
  {32'h4501e3ab, 32'h00000000} /* (20, 8, 18) {real, imag} */,
  {32'h454790ec, 32'h00000000} /* (20, 8, 17) {real, imag} */,
  {32'h4596534b, 32'h00000000} /* (20, 8, 16) {real, imag} */,
  {32'h45d98a2e, 32'h00000000} /* (20, 8, 15) {real, imag} */,
  {32'h45cec44c, 32'h00000000} /* (20, 8, 14) {real, imag} */,
  {32'h45ac4318, 32'h00000000} /* (20, 8, 13) {real, imag} */,
  {32'h457d0e08, 32'h00000000} /* (20, 8, 12) {real, imag} */,
  {32'h454c2ed0, 32'h00000000} /* (20, 8, 11) {real, imag} */,
  {32'h44a9b2bc, 32'h00000000} /* (20, 8, 10) {real, imag} */,
  {32'hc4542db0, 32'h00000000} /* (20, 8, 9) {real, imag} */,
  {32'hc51da0e8, 32'h00000000} /* (20, 8, 8) {real, imag} */,
  {32'hc5477a46, 32'h00000000} /* (20, 8, 7) {real, imag} */,
  {32'hc5976adc, 32'h00000000} /* (20, 8, 6) {real, imag} */,
  {32'hc59dab22, 32'h00000000} /* (20, 8, 5) {real, imag} */,
  {32'hc5cdcabd, 32'h00000000} /* (20, 8, 4) {real, imag} */,
  {32'hc5d1cda6, 32'h00000000} /* (20, 8, 3) {real, imag} */,
  {32'hc5cb503a, 32'h00000000} /* (20, 8, 2) {real, imag} */,
  {32'hc5f399bc, 32'h00000000} /* (20, 8, 1) {real, imag} */,
  {32'hc5ec0019, 32'h00000000} /* (20, 8, 0) {real, imag} */,
  {32'hc60d2fba, 32'h00000000} /* (20, 7, 31) {real, imag} */,
  {32'hc61f6f46, 32'h00000000} /* (20, 7, 30) {real, imag} */,
  {32'hc62e378d, 32'h00000000} /* (20, 7, 29) {real, imag} */,
  {32'hc62a110a, 32'h00000000} /* (20, 7, 28) {real, imag} */,
  {32'hc6226030, 32'h00000000} /* (20, 7, 27) {real, imag} */,
  {32'hc62a0768, 32'h00000000} /* (20, 7, 26) {real, imag} */,
  {32'hc623704b, 32'h00000000} /* (20, 7, 25) {real, imag} */,
  {32'hc61ff58b, 32'h00000000} /* (20, 7, 24) {real, imag} */,
  {32'hc60cbdc8, 32'h00000000} /* (20, 7, 23) {real, imag} */,
  {32'hc5f5dbbe, 32'h00000000} /* (20, 7, 22) {real, imag} */,
  {32'hc5ad2f3b, 32'h00000000} /* (20, 7, 21) {real, imag} */,
  {32'hc4dba6e0, 32'h00000000} /* (20, 7, 20) {real, imag} */,
  {32'h44f605e0, 32'h00000000} /* (20, 7, 19) {real, imag} */,
  {32'h44ee26c6, 32'h00000000} /* (20, 7, 18) {real, imag} */,
  {32'h45722322, 32'h00000000} /* (20, 7, 17) {real, imag} */,
  {32'h45a59134, 32'h00000000} /* (20, 7, 16) {real, imag} */,
  {32'h45cc950d, 32'h00000000} /* (20, 7, 15) {real, imag} */,
  {32'h45d5d7f8, 32'h00000000} /* (20, 7, 14) {real, imag} */,
  {32'h45af5992, 32'h00000000} /* (20, 7, 13) {real, imag} */,
  {32'h45c28f08, 32'h00000000} /* (20, 7, 12) {real, imag} */,
  {32'h45767190, 32'h00000000} /* (20, 7, 11) {real, imag} */,
  {32'h44d1789c, 32'h00000000} /* (20, 7, 10) {real, imag} */,
  {32'hc352afc0, 32'h00000000} /* (20, 7, 9) {real, imag} */,
  {32'hc4d27110, 32'h00000000} /* (20, 7, 8) {real, imag} */,
  {32'hc55d5dda, 32'h00000000} /* (20, 7, 7) {real, imag} */,
  {32'hc5902cc6, 32'h00000000} /* (20, 7, 6) {real, imag} */,
  {32'hc5d10ab5, 32'h00000000} /* (20, 7, 5) {real, imag} */,
  {32'hc5f005dc, 32'h00000000} /* (20, 7, 4) {real, imag} */,
  {32'hc608331a, 32'h00000000} /* (20, 7, 3) {real, imag} */,
  {32'hc612511c, 32'h00000000} /* (20, 7, 2) {real, imag} */,
  {32'hc61008f6, 32'h00000000} /* (20, 7, 1) {real, imag} */,
  {32'hc608a359, 32'h00000000} /* (20, 7, 0) {real, imag} */,
  {32'hc62b45fa, 32'h00000000} /* (20, 6, 31) {real, imag} */,
  {32'hc62d5223, 32'h00000000} /* (20, 6, 30) {real, imag} */,
  {32'hc6383aca, 32'h00000000} /* (20, 6, 29) {real, imag} */,
  {32'hc6414050, 32'h00000000} /* (20, 6, 28) {real, imag} */,
  {32'hc63f556c, 32'h00000000} /* (20, 6, 27) {real, imag} */,
  {32'hc6291c32, 32'h00000000} /* (20, 6, 26) {real, imag} */,
  {32'hc62edeac, 32'h00000000} /* (20, 6, 25) {real, imag} */,
  {32'hc62af978, 32'h00000000} /* (20, 6, 24) {real, imag} */,
  {32'hc6193036, 32'h00000000} /* (20, 6, 23) {real, imag} */,
  {32'hc6039c5b, 32'h00000000} /* (20, 6, 22) {real, imag} */,
  {32'hc5b79711, 32'h00000000} /* (20, 6, 21) {real, imag} */,
  {32'hc548eb3d, 32'h00000000} /* (20, 6, 20) {real, imag} */,
  {32'hc363bc00, 32'h00000000} /* (20, 6, 19) {real, imag} */,
  {32'h445e9588, 32'h00000000} /* (20, 6, 18) {real, imag} */,
  {32'h451378bf, 32'h00000000} /* (20, 6, 17) {real, imag} */,
  {32'h4599f4bd, 32'h00000000} /* (20, 6, 16) {real, imag} */,
  {32'h45d3e0f3, 32'h00000000} /* (20, 6, 15) {real, imag} */,
  {32'h45da1b96, 32'h00000000} /* (20, 6, 14) {real, imag} */,
  {32'h45d9d077, 32'h00000000} /* (20, 6, 13) {real, imag} */,
  {32'h45e987f1, 32'h00000000} /* (20, 6, 12) {real, imag} */,
  {32'h459388e7, 32'h00000000} /* (20, 6, 11) {real, imag} */,
  {32'h4511b444, 32'h00000000} /* (20, 6, 10) {real, imag} */,
  {32'h440be908, 32'h00000000} /* (20, 6, 9) {real, imag} */,
  {32'hc48eff64, 32'h00000000} /* (20, 6, 8) {real, imag} */,
  {32'hc516784e, 32'h00000000} /* (20, 6, 7) {real, imag} */,
  {32'hc5852ff6, 32'h00000000} /* (20, 6, 6) {real, imag} */,
  {32'hc5bc0909, 32'h00000000} /* (20, 6, 5) {real, imag} */,
  {32'hc600fabe, 32'h00000000} /* (20, 6, 4) {real, imag} */,
  {32'hc60ca881, 32'h00000000} /* (20, 6, 3) {real, imag} */,
  {32'hc6114656, 32'h00000000} /* (20, 6, 2) {real, imag} */,
  {32'hc6176a9d, 32'h00000000} /* (20, 6, 1) {real, imag} */,
  {32'hc61aeba2, 32'h00000000} /* (20, 6, 0) {real, imag} */,
  {32'hc630235d, 32'h00000000} /* (20, 5, 31) {real, imag} */,
  {32'hc6407a2c, 32'h00000000} /* (20, 5, 30) {real, imag} */,
  {32'hc64ff786, 32'h00000000} /* (20, 5, 29) {real, imag} */,
  {32'hc63ee008, 32'h00000000} /* (20, 5, 28) {real, imag} */,
  {32'hc64da12a, 32'h00000000} /* (20, 5, 27) {real, imag} */,
  {32'hc64ef771, 32'h00000000} /* (20, 5, 26) {real, imag} */,
  {32'hc63e0ddc, 32'h00000000} /* (20, 5, 25) {real, imag} */,
  {32'hc638f7f0, 32'h00000000} /* (20, 5, 24) {real, imag} */,
  {32'hc6289be4, 32'h00000000} /* (20, 5, 23) {real, imag} */,
  {32'hc60b9119, 32'h00000000} /* (20, 5, 22) {real, imag} */,
  {32'hc5dde5c1, 32'h00000000} /* (20, 5, 21) {real, imag} */,
  {32'hc5a9f046, 32'h00000000} /* (20, 5, 20) {real, imag} */,
  {32'hc54a2bcf, 32'h00000000} /* (20, 5, 19) {real, imag} */,
  {32'hc4073580, 32'h00000000} /* (20, 5, 18) {real, imag} */,
  {32'h44156390, 32'h00000000} /* (20, 5, 17) {real, imag} */,
  {32'h45642e34, 32'h00000000} /* (20, 5, 16) {real, imag} */,
  {32'h45ac2d26, 32'h00000000} /* (20, 5, 15) {real, imag} */,
  {32'h45ca0c29, 32'h00000000} /* (20, 5, 14) {real, imag} */,
  {32'h45e17278, 32'h00000000} /* (20, 5, 13) {real, imag} */,
  {32'h45d4990d, 32'h00000000} /* (20, 5, 12) {real, imag} */,
  {32'h45d02d37, 32'h00000000} /* (20, 5, 11) {real, imag} */,
  {32'h457b91e4, 32'h00000000} /* (20, 5, 10) {real, imag} */,
  {32'h45221afa, 32'h00000000} /* (20, 5, 9) {real, imag} */,
  {32'h44a223b0, 32'h00000000} /* (20, 5, 8) {real, imag} */,
  {32'h436ad420, 32'h00000000} /* (20, 5, 7) {real, imag} */,
  {32'hc50dac1f, 32'h00000000} /* (20, 5, 6) {real, imag} */,
  {32'hc5a6aa57, 32'h00000000} /* (20, 5, 5) {real, imag} */,
  {32'hc5f86cc0, 32'h00000000} /* (20, 5, 4) {real, imag} */,
  {32'hc625d633, 32'h00000000} /* (20, 5, 3) {real, imag} */,
  {32'hc614c590, 32'h00000000} /* (20, 5, 2) {real, imag} */,
  {32'hc627a821, 32'h00000000} /* (20, 5, 1) {real, imag} */,
  {32'hc626f0c7, 32'h00000000} /* (20, 5, 0) {real, imag} */,
  {32'hc638fe0c, 32'h00000000} /* (20, 4, 31) {real, imag} */,
  {32'hc647d2d4, 32'h00000000} /* (20, 4, 30) {real, imag} */,
  {32'hc64f6f77, 32'h00000000} /* (20, 4, 29) {real, imag} */,
  {32'hc6530832, 32'h00000000} /* (20, 4, 28) {real, imag} */,
  {32'hc65219d6, 32'h00000000} /* (20, 4, 27) {real, imag} */,
  {32'hc64f33ae, 32'h00000000} /* (20, 4, 26) {real, imag} */,
  {32'hc6466f93, 32'h00000000} /* (20, 4, 25) {real, imag} */,
  {32'hc651a34e, 32'h00000000} /* (20, 4, 24) {real, imag} */,
  {32'hc633cf32, 32'h00000000} /* (20, 4, 23) {real, imag} */,
  {32'hc6207e18, 32'h00000000} /* (20, 4, 22) {real, imag} */,
  {32'hc6008af6, 32'h00000000} /* (20, 4, 21) {real, imag} */,
  {32'hc5d6803c, 32'h00000000} /* (20, 4, 20) {real, imag} */,
  {32'hc5a09e80, 32'h00000000} /* (20, 4, 19) {real, imag} */,
  {32'hc54c9f70, 32'h00000000} /* (20, 4, 18) {real, imag} */,
  {32'hc41ffeb0, 32'h00000000} /* (20, 4, 17) {real, imag} */,
  {32'h44dc5b14, 32'h00000000} /* (20, 4, 16) {real, imag} */,
  {32'h4573feb0, 32'h00000000} /* (20, 4, 15) {real, imag} */,
  {32'h45c61a8f, 32'h00000000} /* (20, 4, 14) {real, imag} */,
  {32'h45e5ab1a, 32'h00000000} /* (20, 4, 13) {real, imag} */,
  {32'h45d26c93, 32'h00000000} /* (20, 4, 12) {real, imag} */,
  {32'h45cf388c, 32'h00000000} /* (20, 4, 11) {real, imag} */,
  {32'h45bb8725, 32'h00000000} /* (20, 4, 10) {real, imag} */,
  {32'h4594b7ae, 32'h00000000} /* (20, 4, 9) {real, imag} */,
  {32'h459a2b1d, 32'h00000000} /* (20, 4, 8) {real, imag} */,
  {32'h450d2688, 32'h00000000} /* (20, 4, 7) {real, imag} */,
  {32'hc4406a18, 32'h00000000} /* (20, 4, 6) {real, imag} */,
  {32'hc59ca9e5, 32'h00000000} /* (20, 4, 5) {real, imag} */,
  {32'hc5ef7306, 32'h00000000} /* (20, 4, 4) {real, imag} */,
  {32'hc61a85e0, 32'h00000000} /* (20, 4, 3) {real, imag} */,
  {32'hc62a2087, 32'h00000000} /* (20, 4, 2) {real, imag} */,
  {32'hc6292cf7, 32'h00000000} /* (20, 4, 1) {real, imag} */,
  {32'hc6355ca6, 32'h00000000} /* (20, 4, 0) {real, imag} */,
  {32'hc640c90c, 32'h00000000} /* (20, 3, 31) {real, imag} */,
  {32'hc64b732a, 32'h00000000} /* (20, 3, 30) {real, imag} */,
  {32'hc6572f94, 32'h00000000} /* (20, 3, 29) {real, imag} */,
  {32'hc64cf890, 32'h00000000} /* (20, 3, 28) {real, imag} */,
  {32'hc64a5fca, 32'h00000000} /* (20, 3, 27) {real, imag} */,
  {32'hc64f908c, 32'h00000000} /* (20, 3, 26) {real, imag} */,
  {32'hc64dd8ea, 32'h00000000} /* (20, 3, 25) {real, imag} */,
  {32'hc650f21e, 32'h00000000} /* (20, 3, 24) {real, imag} */,
  {32'hc63a6f7e, 32'h00000000} /* (20, 3, 23) {real, imag} */,
  {32'hc6299010, 32'h00000000} /* (20, 3, 22) {real, imag} */,
  {32'hc618cd94, 32'h00000000} /* (20, 3, 21) {real, imag} */,
  {32'hc60bcb5f, 32'h00000000} /* (20, 3, 20) {real, imag} */,
  {32'hc5cc7d7c, 32'h00000000} /* (20, 3, 19) {real, imag} */,
  {32'hc587f11c, 32'h00000000} /* (20, 3, 18) {real, imag} */,
  {32'hc52a7a2e, 32'h00000000} /* (20, 3, 17) {real, imag} */,
  {32'h433e04c0, 32'h00000000} /* (20, 3, 16) {real, imag} */,
  {32'h45717e7e, 32'h00000000} /* (20, 3, 15) {real, imag} */,
  {32'h45b09434, 32'h00000000} /* (20, 3, 14) {real, imag} */,
  {32'h45d0bfe1, 32'h00000000} /* (20, 3, 13) {real, imag} */,
  {32'h45ee4fe5, 32'h00000000} /* (20, 3, 12) {real, imag} */,
  {32'h45d19254, 32'h00000000} /* (20, 3, 11) {real, imag} */,
  {32'h45beb4f0, 32'h00000000} /* (20, 3, 10) {real, imag} */,
  {32'h45c82484, 32'h00000000} /* (20, 3, 9) {real, imag} */,
  {32'h457d5186, 32'h00000000} /* (20, 3, 8) {real, imag} */,
  {32'h45411c9c, 32'h00000000} /* (20, 3, 7) {real, imag} */,
  {32'hc1c61c00, 32'h00000000} /* (20, 3, 6) {real, imag} */,
  {32'hc5a15441, 32'h00000000} /* (20, 3, 5) {real, imag} */,
  {32'hc5e85950, 32'h00000000} /* (20, 3, 4) {real, imag} */,
  {32'hc61b0d76, 32'h00000000} /* (20, 3, 3) {real, imag} */,
  {32'hc6334cd4, 32'h00000000} /* (20, 3, 2) {real, imag} */,
  {32'hc64353ec, 32'h00000000} /* (20, 3, 1) {real, imag} */,
  {32'hc633b07e, 32'h00000000} /* (20, 3, 0) {real, imag} */,
  {32'hc63ce5f7, 32'h00000000} /* (20, 2, 31) {real, imag} */,
  {32'hc653f431, 32'h00000000} /* (20, 2, 30) {real, imag} */,
  {32'hc6541458, 32'h00000000} /* (20, 2, 29) {real, imag} */,
  {32'hc659ec4a, 32'h00000000} /* (20, 2, 28) {real, imag} */,
  {32'hc65cf4cb, 32'h00000000} /* (20, 2, 27) {real, imag} */,
  {32'hc65339a8, 32'h00000000} /* (20, 2, 26) {real, imag} */,
  {32'hc64e1b1f, 32'h00000000} /* (20, 2, 25) {real, imag} */,
  {32'hc64ba5a2, 32'h00000000} /* (20, 2, 24) {real, imag} */,
  {32'hc6440f28, 32'h00000000} /* (20, 2, 23) {real, imag} */,
  {32'hc62e86aa, 32'h00000000} /* (20, 2, 22) {real, imag} */,
  {32'hc6109c24, 32'h00000000} /* (20, 2, 21) {real, imag} */,
  {32'hc5fde5f2, 32'h00000000} /* (20, 2, 20) {real, imag} */,
  {32'hc5c40b10, 32'h00000000} /* (20, 2, 19) {real, imag} */,
  {32'hc5867d38, 32'h00000000} /* (20, 2, 18) {real, imag} */,
  {32'hc505c802, 32'h00000000} /* (20, 2, 17) {real, imag} */,
  {32'hc28b3380, 32'h00000000} /* (20, 2, 16) {real, imag} */,
  {32'h45645c4c, 32'h00000000} /* (20, 2, 15) {real, imag} */,
  {32'h45abde7e, 32'h00000000} /* (20, 2, 14) {real, imag} */,
  {32'h45da27f4, 32'h00000000} /* (20, 2, 13) {real, imag} */,
  {32'h45e03318, 32'h00000000} /* (20, 2, 12) {real, imag} */,
  {32'h45c38fca, 32'h00000000} /* (20, 2, 11) {real, imag} */,
  {32'h45ba5467, 32'h00000000} /* (20, 2, 10) {real, imag} */,
  {32'h4583bca6, 32'h00000000} /* (20, 2, 9) {real, imag} */,
  {32'h453a2ef0, 32'h00000000} /* (20, 2, 8) {real, imag} */,
  {32'h44c0a500, 32'h00000000} /* (20, 2, 7) {real, imag} */,
  {32'hc43991c0, 32'h00000000} /* (20, 2, 6) {real, imag} */,
  {32'hc5746b40, 32'h00000000} /* (20, 2, 5) {real, imag} */,
  {32'hc5efbab6, 32'h00000000} /* (20, 2, 4) {real, imag} */,
  {32'hc625ad2e, 32'h00000000} /* (20, 2, 3) {real, imag} */,
  {32'hc62f872f, 32'h00000000} /* (20, 2, 2) {real, imag} */,
  {32'hc63a0822, 32'h00000000} /* (20, 2, 1) {real, imag} */,
  {32'hc637c301, 32'h00000000} /* (20, 2, 0) {real, imag} */,
  {32'hc6379337, 32'h00000000} /* (20, 1, 31) {real, imag} */,
  {32'hc6485bbb, 32'h00000000} /* (20, 1, 30) {real, imag} */,
  {32'hc650caf1, 32'h00000000} /* (20, 1, 29) {real, imag} */,
  {32'hc663555e, 32'h00000000} /* (20, 1, 28) {real, imag} */,
  {32'hc6600501, 32'h00000000} /* (20, 1, 27) {real, imag} */,
  {32'hc651abce, 32'h00000000} /* (20, 1, 26) {real, imag} */,
  {32'hc6415e54, 32'h00000000} /* (20, 1, 25) {real, imag} */,
  {32'hc646b664, 32'h00000000} /* (20, 1, 24) {real, imag} */,
  {32'hc63bde48, 32'h00000000} /* (20, 1, 23) {real, imag} */,
  {32'hc615411c, 32'h00000000} /* (20, 1, 22) {real, imag} */,
  {32'hc5fc58a6, 32'h00000000} /* (20, 1, 21) {real, imag} */,
  {32'hc5d71599, 32'h00000000} /* (20, 1, 20) {real, imag} */,
  {32'hc59f14d3, 32'h00000000} /* (20, 1, 19) {real, imag} */,
  {32'hc5751805, 32'h00000000} /* (20, 1, 18) {real, imag} */,
  {32'hc4d8f6d4, 32'h00000000} /* (20, 1, 17) {real, imag} */,
  {32'h44d16ea4, 32'h00000000} /* (20, 1, 16) {real, imag} */,
  {32'h458611dc, 32'h00000000} /* (20, 1, 15) {real, imag} */,
  {32'h45a9e9ea, 32'h00000000} /* (20, 1, 14) {real, imag} */,
  {32'h45bdb3e2, 32'h00000000} /* (20, 1, 13) {real, imag} */,
  {32'h45d76fe8, 32'h00000000} /* (20, 1, 12) {real, imag} */,
  {32'h45c226d6, 32'h00000000} /* (20, 1, 11) {real, imag} */,
  {32'h459bb13d, 32'h00000000} /* (20, 1, 10) {real, imag} */,
  {32'h458fcaec, 32'h00000000} /* (20, 1, 9) {real, imag} */,
  {32'h45140d84, 32'h00000000} /* (20, 1, 8) {real, imag} */,
  {32'h4320a380, 32'h00000000} /* (20, 1, 7) {real, imag} */,
  {32'hc42c6060, 32'h00000000} /* (20, 1, 6) {real, imag} */,
  {32'hc593390e, 32'h00000000} /* (20, 1, 5) {real, imag} */,
  {32'hc60ce59c, 32'h00000000} /* (20, 1, 4) {real, imag} */,
  {32'hc6220004, 32'h00000000} /* (20, 1, 3) {real, imag} */,
  {32'hc6265b50, 32'h00000000} /* (20, 1, 2) {real, imag} */,
  {32'hc634c30e, 32'h00000000} /* (20, 1, 1) {real, imag} */,
  {32'hc63811e0, 32'h00000000} /* (20, 1, 0) {real, imag} */,
  {32'hc634169e, 32'h00000000} /* (20, 0, 31) {real, imag} */,
  {32'hc6441e07, 32'h00000000} /* (20, 0, 30) {real, imag} */,
  {32'hc64974d3, 32'h00000000} /* (20, 0, 29) {real, imag} */,
  {32'hc656685c, 32'h00000000} /* (20, 0, 28) {real, imag} */,
  {32'hc656545c, 32'h00000000} /* (20, 0, 27) {real, imag} */,
  {32'hc648b80b, 32'h00000000} /* (20, 0, 26) {real, imag} */,
  {32'hc6422537, 32'h00000000} /* (20, 0, 25) {real, imag} */,
  {32'hc62ee433, 32'h00000000} /* (20, 0, 24) {real, imag} */,
  {32'hc61eb1c1, 32'h00000000} /* (20, 0, 23) {real, imag} */,
  {32'hc6053592, 32'h00000000} /* (20, 0, 22) {real, imag} */,
  {32'hc5da2010, 32'h00000000} /* (20, 0, 21) {real, imag} */,
  {32'hc59f886d, 32'h00000000} /* (20, 0, 20) {real, imag} */,
  {32'hc54cdc2c, 32'h00000000} /* (20, 0, 19) {real, imag} */,
  {32'hc4b92b4c, 32'h00000000} /* (20, 0, 18) {real, imag} */,
  {32'hc2f06900, 32'h00000000} /* (20, 0, 17) {real, imag} */,
  {32'h451c1136, 32'h00000000} /* (20, 0, 16) {real, imag} */,
  {32'h459c94a4, 32'h00000000} /* (20, 0, 15) {real, imag} */,
  {32'h45a6d862, 32'h00000000} /* (20, 0, 14) {real, imag} */,
  {32'h45b5349a, 32'h00000000} /* (20, 0, 13) {real, imag} */,
  {32'h45c16278, 32'h00000000} /* (20, 0, 12) {real, imag} */,
  {32'h45a9d737, 32'h00000000} /* (20, 0, 11) {real, imag} */,
  {32'h4565cab4, 32'h00000000} /* (20, 0, 10) {real, imag} */,
  {32'h4518d000, 32'h00000000} /* (20, 0, 9) {real, imag} */,
  {32'h443f9b60, 32'h00000000} /* (20, 0, 8) {real, imag} */,
  {32'hc4c97148, 32'h00000000} /* (20, 0, 7) {real, imag} */,
  {32'hc563e0b2, 32'h00000000} /* (20, 0, 6) {real, imag} */,
  {32'hc5ba82b0, 32'h00000000} /* (20, 0, 5) {real, imag} */,
  {32'hc5fb4233, 32'h00000000} /* (20, 0, 4) {real, imag} */,
  {32'hc615bbc6, 32'h00000000} /* (20, 0, 3) {real, imag} */,
  {32'hc6235e34, 32'h00000000} /* (20, 0, 2) {real, imag} */,
  {32'hc634b039, 32'h00000000} /* (20, 0, 1) {real, imag} */,
  {32'hc6445520, 32'h00000000} /* (20, 0, 0) {real, imag} */,
  {32'hc6320f18, 32'h00000000} /* (19, 31, 31) {real, imag} */,
  {32'hc6424258, 32'h00000000} /* (19, 31, 30) {real, imag} */,
  {32'hc638938c, 32'h00000000} /* (19, 31, 29) {real, imag} */,
  {32'hc63df1ca, 32'h00000000} /* (19, 31, 28) {real, imag} */,
  {32'hc6451140, 32'h00000000} /* (19, 31, 27) {real, imag} */,
  {32'hc63aebef, 32'h00000000} /* (19, 31, 26) {real, imag} */,
  {32'hc6264f68, 32'h00000000} /* (19, 31, 25) {real, imag} */,
  {32'hc61900b8, 32'h00000000} /* (19, 31, 24) {real, imag} */,
  {32'hc60ad893, 32'h00000000} /* (19, 31, 23) {real, imag} */,
  {32'hc5e660de, 32'h00000000} /* (19, 31, 22) {real, imag} */,
  {32'hc59f73f0, 32'h00000000} /* (19, 31, 21) {real, imag} */,
  {32'hc5409ef0, 32'h00000000} /* (19, 31, 20) {real, imag} */,
  {32'hc4204570, 32'h00000000} /* (19, 31, 19) {real, imag} */,
  {32'h44c8c55c, 32'h00000000} /* (19, 31, 18) {real, imag} */,
  {32'h45266602, 32'h00000000} /* (19, 31, 17) {real, imag} */,
  {32'h457a81f8, 32'h00000000} /* (19, 31, 16) {real, imag} */,
  {32'h45aa77d5, 32'h00000000} /* (19, 31, 15) {real, imag} */,
  {32'h45ad3d84, 32'h00000000} /* (19, 31, 14) {real, imag} */,
  {32'h45a8c82c, 32'h00000000} /* (19, 31, 13) {real, imag} */,
  {32'h45a9fc2d, 32'h00000000} /* (19, 31, 12) {real, imag} */,
  {32'h457a9808, 32'h00000000} /* (19, 31, 11) {real, imag} */,
  {32'h449ea430, 32'h00000000} /* (19, 31, 10) {real, imag} */,
  {32'hc38bd810, 32'h00000000} /* (19, 31, 9) {real, imag} */,
  {32'hc50a8190, 32'h00000000} /* (19, 31, 8) {real, imag} */,
  {32'hc5655398, 32'h00000000} /* (19, 31, 7) {real, imag} */,
  {32'hc5afc19e, 32'h00000000} /* (19, 31, 6) {real, imag} */,
  {32'hc5eb53cc, 32'h00000000} /* (19, 31, 5) {real, imag} */,
  {32'hc6030f9f, 32'h00000000} /* (19, 31, 4) {real, imag} */,
  {32'hc60f68a1, 32'h00000000} /* (19, 31, 3) {real, imag} */,
  {32'hc625dd3e, 32'h00000000} /* (19, 31, 2) {real, imag} */,
  {32'hc62c8f98, 32'h00000000} /* (19, 31, 1) {real, imag} */,
  {32'hc62bb8c4, 32'h00000000} /* (19, 31, 0) {real, imag} */,
  {32'hc6320db8, 32'h00000000} /* (19, 30, 31) {real, imag} */,
  {32'hc646632f, 32'h00000000} /* (19, 30, 30) {real, imag} */,
  {32'hc6436c36, 32'h00000000} /* (19, 30, 29) {real, imag} */,
  {32'hc63e4468, 32'h00000000} /* (19, 30, 28) {real, imag} */,
  {32'hc6477aa1, 32'h00000000} /* (19, 30, 27) {real, imag} */,
  {32'hc654c714, 32'h00000000} /* (19, 30, 26) {real, imag} */,
  {32'hc62e8332, 32'h00000000} /* (19, 30, 25) {real, imag} */,
  {32'hc621460c, 32'h00000000} /* (19, 30, 24) {real, imag} */,
  {32'hc6146b1e, 32'h00000000} /* (19, 30, 23) {real, imag} */,
  {32'hc5dbaebc, 32'h00000000} /* (19, 30, 22) {real, imag} */,
  {32'hc596b8f4, 32'h00000000} /* (19, 30, 21) {real, imag} */,
  {32'hc49bd970, 32'h00000000} /* (19, 30, 20) {real, imag} */,
  {32'h446de0a0, 32'h00000000} /* (19, 30, 19) {real, imag} */,
  {32'h4558a794, 32'h00000000} /* (19, 30, 18) {real, imag} */,
  {32'h45a10a92, 32'h00000000} /* (19, 30, 17) {real, imag} */,
  {32'h45cee1fa, 32'h00000000} /* (19, 30, 16) {real, imag} */,
  {32'h45d3ce65, 32'h00000000} /* (19, 30, 15) {real, imag} */,
  {32'h45e2c092, 32'h00000000} /* (19, 30, 14) {real, imag} */,
  {32'h45c90cd0, 32'h00000000} /* (19, 30, 13) {real, imag} */,
  {32'h4599233b, 32'h00000000} /* (19, 30, 12) {real, imag} */,
  {32'h455ea284, 32'h00000000} /* (19, 30, 11) {real, imag} */,
  {32'h44c2ad70, 32'h00000000} /* (19, 30, 10) {real, imag} */,
  {32'hc5066416, 32'h00000000} /* (19, 30, 9) {real, imag} */,
  {32'hc582ea6b, 32'h00000000} /* (19, 30, 8) {real, imag} */,
  {32'hc5c74e49, 32'h00000000} /* (19, 30, 7) {real, imag} */,
  {32'hc5ddca74, 32'h00000000} /* (19, 30, 6) {real, imag} */,
  {32'hc6063bc6, 32'h00000000} /* (19, 30, 5) {real, imag} */,
  {32'hc61a622b, 32'h00000000} /* (19, 30, 4) {real, imag} */,
  {32'hc624fe1e, 32'h00000000} /* (19, 30, 3) {real, imag} */,
  {32'hc62c2cf9, 32'h00000000} /* (19, 30, 2) {real, imag} */,
  {32'hc63043c7, 32'h00000000} /* (19, 30, 1) {real, imag} */,
  {32'hc62ae94f, 32'h00000000} /* (19, 30, 0) {real, imag} */,
  {32'hc63c1959, 32'h00000000} /* (19, 29, 31) {real, imag} */,
  {32'hc639fb82, 32'h00000000} /* (19, 29, 30) {real, imag} */,
  {32'hc63c6ab7, 32'h00000000} /* (19, 29, 29) {real, imag} */,
  {32'hc641480b, 32'h00000000} /* (19, 29, 28) {real, imag} */,
  {32'hc63cedfb, 32'h00000000} /* (19, 29, 27) {real, imag} */,
  {32'hc63b3094, 32'h00000000} /* (19, 29, 26) {real, imag} */,
  {32'hc6328208, 32'h00000000} /* (19, 29, 25) {real, imag} */,
  {32'hc62c6810, 32'h00000000} /* (19, 29, 24) {real, imag} */,
  {32'hc61f1dae, 32'h00000000} /* (19, 29, 23) {real, imag} */,
  {32'hc5dd7b6d, 32'h00000000} /* (19, 29, 22) {real, imag} */,
  {32'hc548710b, 32'h00000000} /* (19, 29, 21) {real, imag} */,
  {32'h449155c8, 32'h00000000} /* (19, 29, 20) {real, imag} */,
  {32'h45023af4, 32'h00000000} /* (19, 29, 19) {real, imag} */,
  {32'h45964ff4, 32'h00000000} /* (19, 29, 18) {real, imag} */,
  {32'h45cdeb04, 32'h00000000} /* (19, 29, 17) {real, imag} */,
  {32'h45d37aa4, 32'h00000000} /* (19, 29, 16) {real, imag} */,
  {32'h45de860a, 32'h00000000} /* (19, 29, 15) {real, imag} */,
  {32'h45f44fec, 32'h00000000} /* (19, 29, 14) {real, imag} */,
  {32'h45e47566, 32'h00000000} /* (19, 29, 13) {real, imag} */,
  {32'h45a8c406, 32'h00000000} /* (19, 29, 12) {real, imag} */,
  {32'h45386c04, 32'h00000000} /* (19, 29, 11) {real, imag} */,
  {32'h4374c160, 32'h00000000} /* (19, 29, 10) {real, imag} */,
  {32'hc539ae7e, 32'h00000000} /* (19, 29, 9) {real, imag} */,
  {32'hc5b64450, 32'h00000000} /* (19, 29, 8) {real, imag} */,
  {32'hc5ed1be4, 32'h00000000} /* (19, 29, 7) {real, imag} */,
  {32'hc602b65c, 32'h00000000} /* (19, 29, 6) {real, imag} */,
  {32'hc61890e7, 32'h00000000} /* (19, 29, 5) {real, imag} */,
  {32'hc61d4981, 32'h00000000} /* (19, 29, 4) {real, imag} */,
  {32'hc62ce92b, 32'h00000000} /* (19, 29, 3) {real, imag} */,
  {32'hc62eee61, 32'h00000000} /* (19, 29, 2) {real, imag} */,
  {32'hc63a6fb0, 32'h00000000} /* (19, 29, 1) {real, imag} */,
  {32'hc635eba6, 32'h00000000} /* (19, 29, 0) {real, imag} */,
  {32'hc635f538, 32'h00000000} /* (19, 28, 31) {real, imag} */,
  {32'hc63aa954, 32'h00000000} /* (19, 28, 30) {real, imag} */,
  {32'hc643c983, 32'h00000000} /* (19, 28, 29) {real, imag} */,
  {32'hc6563796, 32'h00000000} /* (19, 28, 28) {real, imag} */,
  {32'hc63cefcc, 32'h00000000} /* (19, 28, 27) {real, imag} */,
  {32'hc641c7af, 32'h00000000} /* (19, 28, 26) {real, imag} */,
  {32'hc63a5326, 32'h00000000} /* (19, 28, 25) {real, imag} */,
  {32'hc64716da, 32'h00000000} /* (19, 28, 24) {real, imag} */,
  {32'hc615a602, 32'h00000000} /* (19, 28, 23) {real, imag} */,
  {32'hc5d65474, 32'h00000000} /* (19, 28, 22) {real, imag} */,
  {32'hc548101f, 32'h00000000} /* (19, 28, 21) {real, imag} */,
  {32'h4501dae0, 32'h00000000} /* (19, 28, 20) {real, imag} */,
  {32'h454629b1, 32'h00000000} /* (19, 28, 19) {real, imag} */,
  {32'h45b14d44, 32'h00000000} /* (19, 28, 18) {real, imag} */,
  {32'h45ce5860, 32'h00000000} /* (19, 28, 17) {real, imag} */,
  {32'h45fd799b, 32'h00000000} /* (19, 28, 16) {real, imag} */,
  {32'h45ee1528, 32'h00000000} /* (19, 28, 15) {real, imag} */,
  {32'h45ecbacc, 32'h00000000} /* (19, 28, 14) {real, imag} */,
  {32'h45e09b1e, 32'h00000000} /* (19, 28, 13) {real, imag} */,
  {32'h459bc62f, 32'h00000000} /* (19, 28, 12) {real, imag} */,
  {32'h4529cd70, 32'h00000000} /* (19, 28, 11) {real, imag} */,
  {32'hc41536f0, 32'h00000000} /* (19, 28, 10) {real, imag} */,
  {32'hc5652ce6, 32'h00000000} /* (19, 28, 9) {real, imag} */,
  {32'hc5bcf3d4, 32'h00000000} /* (19, 28, 8) {real, imag} */,
  {32'hc5ea168b, 32'h00000000} /* (19, 28, 7) {real, imag} */,
  {32'hc6119f08, 32'h00000000} /* (19, 28, 6) {real, imag} */,
  {32'hc61aded0, 32'h00000000} /* (19, 28, 5) {real, imag} */,
  {32'hc625c09b, 32'h00000000} /* (19, 28, 4) {real, imag} */,
  {32'hc6314dbd, 32'h00000000} /* (19, 28, 3) {real, imag} */,
  {32'hc6371bf0, 32'h00000000} /* (19, 28, 2) {real, imag} */,
  {32'hc63f8e20, 32'h00000000} /* (19, 28, 1) {real, imag} */,
  {32'hc636d3e4, 32'h00000000} /* (19, 28, 0) {real, imag} */,
  {32'hc637b43a, 32'h00000000} /* (19, 27, 31) {real, imag} */,
  {32'hc63f394a, 32'h00000000} /* (19, 27, 30) {real, imag} */,
  {32'hc641059e, 32'h00000000} /* (19, 27, 29) {real, imag} */,
  {32'hc6330a98, 32'h00000000} /* (19, 27, 28) {real, imag} */,
  {32'hc633396e, 32'h00000000} /* (19, 27, 27) {real, imag} */,
  {32'hc63595d4, 32'h00000000} /* (19, 27, 26) {real, imag} */,
  {32'hc648988f, 32'h00000000} /* (19, 27, 25) {real, imag} */,
  {32'hc630b340, 32'h00000000} /* (19, 27, 24) {real, imag} */,
  {32'hc60fdf14, 32'h00000000} /* (19, 27, 23) {real, imag} */,
  {32'hc5b5ea9e, 32'h00000000} /* (19, 27, 22) {real, imag} */,
  {32'hc53e9c5a, 32'h00000000} /* (19, 27, 21) {real, imag} */,
  {32'h444bc668, 32'h00000000} /* (19, 27, 20) {real, imag} */,
  {32'h4556826f, 32'h00000000} /* (19, 27, 19) {real, imag} */,
  {32'h45917a59, 32'h00000000} /* (19, 27, 18) {real, imag} */,
  {32'h45d96305, 32'h00000000} /* (19, 27, 17) {real, imag} */,
  {32'h45f4c424, 32'h00000000} /* (19, 27, 16) {real, imag} */,
  {32'h46024274, 32'h00000000} /* (19, 27, 15) {real, imag} */,
  {32'h46009d88, 32'h00000000} /* (19, 27, 14) {real, imag} */,
  {32'h45c9d859, 32'h00000000} /* (19, 27, 13) {real, imag} */,
  {32'h45965180, 32'h00000000} /* (19, 27, 12) {real, imag} */,
  {32'h44e45514, 32'h00000000} /* (19, 27, 11) {real, imag} */,
  {32'hc4b7338c, 32'h00000000} /* (19, 27, 10) {real, imag} */,
  {32'hc5aae522, 32'h00000000} /* (19, 27, 9) {real, imag} */,
  {32'hc5d565a7, 32'h00000000} /* (19, 27, 8) {real, imag} */,
  {32'hc5ffb26c, 32'h00000000} /* (19, 27, 7) {real, imag} */,
  {32'hc61bad7d, 32'h00000000} /* (19, 27, 6) {real, imag} */,
  {32'hc6293b18, 32'h00000000} /* (19, 27, 5) {real, imag} */,
  {32'hc63128ae, 32'h00000000} /* (19, 27, 4) {real, imag} */,
  {32'hc62cf0f4, 32'h00000000} /* (19, 27, 3) {real, imag} */,
  {32'hc62f25e8, 32'h00000000} /* (19, 27, 2) {real, imag} */,
  {32'hc636157e, 32'h00000000} /* (19, 27, 1) {real, imag} */,
  {32'hc62f09de, 32'h00000000} /* (19, 27, 0) {real, imag} */,
  {32'hc62a38d7, 32'h00000000} /* (19, 26, 31) {real, imag} */,
  {32'hc62a607f, 32'h00000000} /* (19, 26, 30) {real, imag} */,
  {32'hc62ef102, 32'h00000000} /* (19, 26, 29) {real, imag} */,
  {32'hc63ea3ce, 32'h00000000} /* (19, 26, 28) {real, imag} */,
  {32'hc6314f74, 32'h00000000} /* (19, 26, 27) {real, imag} */,
  {32'hc629489a, 32'h00000000} /* (19, 26, 26) {real, imag} */,
  {32'hc62ede2f, 32'h00000000} /* (19, 26, 25) {real, imag} */,
  {32'hc619cdd3, 32'h00000000} /* (19, 26, 24) {real, imag} */,
  {32'hc60714e0, 32'h00000000} /* (19, 26, 23) {real, imag} */,
  {32'hc5bd5d5c, 32'h00000000} /* (19, 26, 22) {real, imag} */,
  {32'hc52df6e9, 32'h00000000} /* (19, 26, 21) {real, imag} */,
  {32'h438d9a70, 32'h00000000} /* (19, 26, 20) {real, imag} */,
  {32'h45433b2b, 32'h00000000} /* (19, 26, 19) {real, imag} */,
  {32'h459ac9e5, 32'h00000000} /* (19, 26, 18) {real, imag} */,
  {32'h45d1eff2, 32'h00000000} /* (19, 26, 17) {real, imag} */,
  {32'h45cb0081, 32'h00000000} /* (19, 26, 16) {real, imag} */,
  {32'h4600ac0d, 32'h00000000} /* (19, 26, 15) {real, imag} */,
  {32'h45fab77a, 32'h00000000} /* (19, 26, 14) {real, imag} */,
  {32'h45e09b24, 32'h00000000} /* (19, 26, 13) {real, imag} */,
  {32'h459edb30, 32'h00000000} /* (19, 26, 12) {real, imag} */,
  {32'h44b81450, 32'h00000000} /* (19, 26, 11) {real, imag} */,
  {32'hc4b3ca30, 32'h00000000} /* (19, 26, 10) {real, imag} */,
  {32'hc5a61312, 32'h00000000} /* (19, 26, 9) {real, imag} */,
  {32'hc60290dd, 32'h00000000} /* (19, 26, 8) {real, imag} */,
  {32'hc60a4808, 32'h00000000} /* (19, 26, 7) {real, imag} */,
  {32'hc613f614, 32'h00000000} /* (19, 26, 6) {real, imag} */,
  {32'hc6270848, 32'h00000000} /* (19, 26, 5) {real, imag} */,
  {32'hc62743e4, 32'h00000000} /* (19, 26, 4) {real, imag} */,
  {32'hc6274d72, 32'h00000000} /* (19, 26, 3) {real, imag} */,
  {32'hc62ec40a, 32'h00000000} /* (19, 26, 2) {real, imag} */,
  {32'hc6386683, 32'h00000000} /* (19, 26, 1) {real, imag} */,
  {32'hc631df56, 32'h00000000} /* (19, 26, 0) {real, imag} */,
  {32'hc61e019a, 32'h00000000} /* (19, 25, 31) {real, imag} */,
  {32'hc6286dd3, 32'h00000000} /* (19, 25, 30) {real, imag} */,
  {32'hc624d798, 32'h00000000} /* (19, 25, 29) {real, imag} */,
  {32'hc6245f56, 32'h00000000} /* (19, 25, 28) {real, imag} */,
  {32'hc62da435, 32'h00000000} /* (19, 25, 27) {real, imag} */,
  {32'hc6324ec4, 32'h00000000} /* (19, 25, 26) {real, imag} */,
  {32'hc61ff225, 32'h00000000} /* (19, 25, 25) {real, imag} */,
  {32'hc60a5b3c, 32'h00000000} /* (19, 25, 24) {real, imag} */,
  {32'hc5f9745a, 32'h00000000} /* (19, 25, 23) {real, imag} */,
  {32'hc5d77934, 32'h00000000} /* (19, 25, 22) {real, imag} */,
  {32'hc5612d9f, 32'h00000000} /* (19, 25, 21) {real, imag} */,
  {32'h449d4fc8, 32'h00000000} /* (19, 25, 20) {real, imag} */,
  {32'h4581a922, 32'h00000000} /* (19, 25, 19) {real, imag} */,
  {32'h45a2b670, 32'h00000000} /* (19, 25, 18) {real, imag} */,
  {32'h45c5d9fa, 32'h00000000} /* (19, 25, 17) {real, imag} */,
  {32'h45baee84, 32'h00000000} /* (19, 25, 16) {real, imag} */,
  {32'h45d86288, 32'h00000000} /* (19, 25, 15) {real, imag} */,
  {32'h45d0adba, 32'h00000000} /* (19, 25, 14) {real, imag} */,
  {32'h45ed2383, 32'h00000000} /* (19, 25, 13) {real, imag} */,
  {32'h457d91a6, 32'h00000000} /* (19, 25, 12) {real, imag} */,
  {32'h44a2e660, 32'h00000000} /* (19, 25, 11) {real, imag} */,
  {32'hc4e2ff4c, 32'h00000000} /* (19, 25, 10) {real, imag} */,
  {32'hc5ac3bba, 32'h00000000} /* (19, 25, 9) {real, imag} */,
  {32'hc5fd2d30, 32'h00000000} /* (19, 25, 8) {real, imag} */,
  {32'hc60aa845, 32'h00000000} /* (19, 25, 7) {real, imag} */,
  {32'hc60b1c4a, 32'h00000000} /* (19, 25, 6) {real, imag} */,
  {32'hc60c9bd9, 32'h00000000} /* (19, 25, 5) {real, imag} */,
  {32'hc61da218, 32'h00000000} /* (19, 25, 4) {real, imag} */,
  {32'hc61e884b, 32'h00000000} /* (19, 25, 3) {real, imag} */,
  {32'hc6313fe0, 32'h00000000} /* (19, 25, 2) {real, imag} */,
  {32'hc63c17f7, 32'h00000000} /* (19, 25, 1) {real, imag} */,
  {32'hc61f40a2, 32'h00000000} /* (19, 25, 0) {real, imag} */,
  {32'hc6058a22, 32'h00000000} /* (19, 24, 31) {real, imag} */,
  {32'hc6096a44, 32'h00000000} /* (19, 24, 30) {real, imag} */,
  {32'hc608705f, 32'h00000000} /* (19, 24, 29) {real, imag} */,
  {32'hc608e04a, 32'h00000000} /* (19, 24, 28) {real, imag} */,
  {32'hc617aac2, 32'h00000000} /* (19, 24, 27) {real, imag} */,
  {32'hc6087190, 32'h00000000} /* (19, 24, 26) {real, imag} */,
  {32'hc60ba91b, 32'h00000000} /* (19, 24, 25) {real, imag} */,
  {32'hc5f9cc5b, 32'h00000000} /* (19, 24, 24) {real, imag} */,
  {32'hc6094864, 32'h00000000} /* (19, 24, 23) {real, imag} */,
  {32'hc5aac069, 32'h00000000} /* (19, 24, 22) {real, imag} */,
  {32'hc50d56ed, 32'h00000000} /* (19, 24, 21) {real, imag} */,
  {32'h44d45370, 32'h00000000} /* (19, 24, 20) {real, imag} */,
  {32'h456af35f, 32'h00000000} /* (19, 24, 19) {real, imag} */,
  {32'h45a935c3, 32'h00000000} /* (19, 24, 18) {real, imag} */,
  {32'h45b3de7c, 32'h00000000} /* (19, 24, 17) {real, imag} */,
  {32'h45bbd9f7, 32'h00000000} /* (19, 24, 16) {real, imag} */,
  {32'h45d0bba1, 32'h00000000} /* (19, 24, 15) {real, imag} */,
  {32'h45d8d50c, 32'h00000000} /* (19, 24, 14) {real, imag} */,
  {32'h458db2fe, 32'h00000000} /* (19, 24, 13) {real, imag} */,
  {32'h455fbb0a, 32'h00000000} /* (19, 24, 12) {real, imag} */,
  {32'h44a299f4, 32'h00000000} /* (19, 24, 11) {real, imag} */,
  {32'hc528b6c0, 32'h00000000} /* (19, 24, 10) {real, imag} */,
  {32'hc5b6147a, 32'h00000000} /* (19, 24, 9) {real, imag} */,
  {32'hc5fff3d3, 32'h00000000} /* (19, 24, 8) {real, imag} */,
  {32'hc600bbd4, 32'h00000000} /* (19, 24, 7) {real, imag} */,
  {32'hc5f641bb, 32'h00000000} /* (19, 24, 6) {real, imag} */,
  {32'hc605a1cf, 32'h00000000} /* (19, 24, 5) {real, imag} */,
  {32'hc60af506, 32'h00000000} /* (19, 24, 4) {real, imag} */,
  {32'hc61143b9, 32'h00000000} /* (19, 24, 3) {real, imag} */,
  {32'hc61b3a46, 32'h00000000} /* (19, 24, 2) {real, imag} */,
  {32'hc616c244, 32'h00000000} /* (19, 24, 1) {real, imag} */,
  {32'hc60a8998, 32'h00000000} /* (19, 24, 0) {real, imag} */,
  {32'hc5e4c5b4, 32'h00000000} /* (19, 23, 31) {real, imag} */,
  {32'hc5e22428, 32'h00000000} /* (19, 23, 30) {real, imag} */,
  {32'hc5dd531c, 32'h00000000} /* (19, 23, 29) {real, imag} */,
  {32'hc5ef8d2c, 32'h00000000} /* (19, 23, 28) {real, imag} */,
  {32'hc5df66f5, 32'h00000000} /* (19, 23, 27) {real, imag} */,
  {32'hc5d95d1a, 32'h00000000} /* (19, 23, 26) {real, imag} */,
  {32'hc5dd488f, 32'h00000000} /* (19, 23, 25) {real, imag} */,
  {32'hc5f5bb77, 32'h00000000} /* (19, 23, 24) {real, imag} */,
  {32'hc5efa632, 32'h00000000} /* (19, 23, 23) {real, imag} */,
  {32'hc5b9f599, 32'h00000000} /* (19, 23, 22) {real, imag} */,
  {32'hc53d5367, 32'h00000000} /* (19, 23, 21) {real, imag} */,
  {32'h448f6fea, 32'h00000000} /* (19, 23, 20) {real, imag} */,
  {32'h45719664, 32'h00000000} /* (19, 23, 19) {real, imag} */,
  {32'h45b5a432, 32'h00000000} /* (19, 23, 18) {real, imag} */,
  {32'h458eb898, 32'h00000000} /* (19, 23, 17) {real, imag} */,
  {32'h45a7dd42, 32'h00000000} /* (19, 23, 16) {real, imag} */,
  {32'h45acb0f4, 32'h00000000} /* (19, 23, 15) {real, imag} */,
  {32'h45ac4a6e, 32'h00000000} /* (19, 23, 14) {real, imag} */,
  {32'h455d17f4, 32'h00000000} /* (19, 23, 13) {real, imag} */,
  {32'h454a3d67, 32'h00000000} /* (19, 23, 12) {real, imag} */,
  {32'h445f0118, 32'h00000000} /* (19, 23, 11) {real, imag} */,
  {32'hc53ef988, 32'h00000000} /* (19, 23, 10) {real, imag} */,
  {32'hc5882aad, 32'h00000000} /* (19, 23, 9) {real, imag} */,
  {32'hc5b5d015, 32'h00000000} /* (19, 23, 8) {real, imag} */,
  {32'hc5cce99a, 32'h00000000} /* (19, 23, 7) {real, imag} */,
  {32'hc5ed65af, 32'h00000000} /* (19, 23, 6) {real, imag} */,
  {32'hc600c7fe, 32'h00000000} /* (19, 23, 5) {real, imag} */,
  {32'hc5f3dd4c, 32'h00000000} /* (19, 23, 4) {real, imag} */,
  {32'hc5f54fce, 32'h00000000} /* (19, 23, 3) {real, imag} */,
  {32'hc5fb842e, 32'h00000000} /* (19, 23, 2) {real, imag} */,
  {32'hc5fa2e4c, 32'h00000000} /* (19, 23, 1) {real, imag} */,
  {32'hc5d83afa, 32'h00000000} /* (19, 23, 0) {real, imag} */,
  {32'hc5874a7f, 32'h00000000} /* (19, 22, 31) {real, imag} */,
  {32'hc5ba1a14, 32'h00000000} /* (19, 22, 30) {real, imag} */,
  {32'hc5be5598, 32'h00000000} /* (19, 22, 29) {real, imag} */,
  {32'hc5bc20a5, 32'h00000000} /* (19, 22, 28) {real, imag} */,
  {32'hc5bdb8ec, 32'h00000000} /* (19, 22, 27) {real, imag} */,
  {32'hc5b26197, 32'h00000000} /* (19, 22, 26) {real, imag} */,
  {32'hc590bbb8, 32'h00000000} /* (19, 22, 25) {real, imag} */,
  {32'hc592683d, 32'h00000000} /* (19, 22, 24) {real, imag} */,
  {32'hc5931f67, 32'h00000000} /* (19, 22, 23) {real, imag} */,
  {32'hc57e6fd0, 32'h00000000} /* (19, 22, 22) {real, imag} */,
  {32'hc5097384, 32'h00000000} /* (19, 22, 21) {real, imag} */,
  {32'h442ac3c4, 32'h00000000} /* (19, 22, 20) {real, imag} */,
  {32'h450e251c, 32'h00000000} /* (19, 22, 19) {real, imag} */,
  {32'h452a40db, 32'h00000000} /* (19, 22, 18) {real, imag} */,
  {32'h454e0b39, 32'h00000000} /* (19, 22, 17) {real, imag} */,
  {32'h45828064, 32'h00000000} /* (19, 22, 16) {real, imag} */,
  {32'h4549a1ae, 32'h00000000} /* (19, 22, 15) {real, imag} */,
  {32'h455b8f27, 32'h00000000} /* (19, 22, 14) {real, imag} */,
  {32'h4569d245, 32'h00000000} /* (19, 22, 13) {real, imag} */,
  {32'h449ee014, 32'h00000000} /* (19, 22, 12) {real, imag} */,
  {32'h43b03298, 32'h00000000} /* (19, 22, 11) {real, imag} */,
  {32'hc516f9ac, 32'h00000000} /* (19, 22, 10) {real, imag} */,
  {32'hc590d8f8, 32'h00000000} /* (19, 22, 9) {real, imag} */,
  {32'hc58e8fb7, 32'h00000000} /* (19, 22, 8) {real, imag} */,
  {32'hc5a41bef, 32'h00000000} /* (19, 22, 7) {real, imag} */,
  {32'hc59cd224, 32'h00000000} /* (19, 22, 6) {real, imag} */,
  {32'hc58bceed, 32'h00000000} /* (19, 22, 5) {real, imag} */,
  {32'hc5ac397e, 32'h00000000} /* (19, 22, 4) {real, imag} */,
  {32'hc5a0943e, 32'h00000000} /* (19, 22, 3) {real, imag} */,
  {32'hc5c4d644, 32'h00000000} /* (19, 22, 2) {real, imag} */,
  {32'hc5d201da, 32'h00000000} /* (19, 22, 1) {real, imag} */,
  {32'hc5b32a0a, 32'h00000000} /* (19, 22, 0) {real, imag} */,
  {32'hc5102ed6, 32'h00000000} /* (19, 21, 31) {real, imag} */,
  {32'hc516b8c8, 32'h00000000} /* (19, 21, 30) {real, imag} */,
  {32'hc5298e18, 32'h00000000} /* (19, 21, 29) {real, imag} */,
  {32'hc51b6df4, 32'h00000000} /* (19, 21, 28) {real, imag} */,
  {32'hc524f418, 32'h00000000} /* (19, 21, 27) {real, imag} */,
  {32'hc52a1083, 32'h00000000} /* (19, 21, 26) {real, imag} */,
  {32'hc50af0fc, 32'h00000000} /* (19, 21, 25) {real, imag} */,
  {32'hc4e84f14, 32'h00000000} /* (19, 21, 24) {real, imag} */,
  {32'hc4fe1720, 32'h00000000} /* (19, 21, 23) {real, imag} */,
  {32'hc4977a92, 32'h00000000} /* (19, 21, 22) {real, imag} */,
  {32'hc42d1c58, 32'h00000000} /* (19, 21, 21) {real, imag} */,
  {32'hc450013b, 32'h00000000} /* (19, 21, 20) {real, imag} */,
  {32'h42c22fb8, 32'h00000000} /* (19, 21, 19) {real, imag} */,
  {32'h43b77c3c, 32'h00000000} /* (19, 21, 18) {real, imag} */,
  {32'h443428a6, 32'h00000000} /* (19, 21, 17) {real, imag} */,
  {32'h44497272, 32'h00000000} /* (19, 21, 16) {real, imag} */,
  {32'h44997652, 32'h00000000} /* (19, 21, 15) {real, imag} */,
  {32'h44988154, 32'h00000000} /* (19, 21, 14) {real, imag} */,
  {32'h44949879, 32'h00000000} /* (19, 21, 13) {real, imag} */,
  {32'h43ef7194, 32'h00000000} /* (19, 21, 12) {real, imag} */,
  {32'hc3df0d2c, 32'h00000000} /* (19, 21, 11) {real, imag} */,
  {32'hc509c629, 32'h00000000} /* (19, 21, 10) {real, imag} */,
  {32'hc51d005a, 32'h00000000} /* (19, 21, 9) {real, imag} */,
  {32'hc51bd8fa, 32'h00000000} /* (19, 21, 8) {real, imag} */,
  {32'hc51d2748, 32'h00000000} /* (19, 21, 7) {real, imag} */,
  {32'hc4e2bf5a, 32'h00000000} /* (19, 21, 6) {real, imag} */,
  {32'hc4c6d994, 32'h00000000} /* (19, 21, 5) {real, imag} */,
  {32'hc49b2143, 32'h00000000} /* (19, 21, 4) {real, imag} */,
  {32'hc4e90336, 32'h00000000} /* (19, 21, 3) {real, imag} */,
  {32'hc5125aa0, 32'h00000000} /* (19, 21, 2) {real, imag} */,
  {32'hc507bf48, 32'h00000000} /* (19, 21, 1) {real, imag} */,
  {32'hc4e7ba7b, 32'h00000000} /* (19, 21, 0) {real, imag} */,
  {32'h44c11216, 32'h00000000} /* (19, 20, 31) {real, imag} */,
  {32'h44c4d97a, 32'h00000000} /* (19, 20, 30) {real, imag} */,
  {32'h448fbffb, 32'h00000000} /* (19, 20, 29) {real, imag} */,
  {32'h45148c4b, 32'h00000000} /* (19, 20, 28) {real, imag} */,
  {32'h452d4198, 32'h00000000} /* (19, 20, 27) {real, imag} */,
  {32'h44cf32f2, 32'h00000000} /* (19, 20, 26) {real, imag} */,
  {32'h448c4dd7, 32'h00000000} /* (19, 20, 25) {real, imag} */,
  {32'h44ef82cc, 32'h00000000} /* (19, 20, 24) {real, imag} */,
  {32'h44ec5f17, 32'h00000000} /* (19, 20, 23) {real, imag} */,
  {32'h44572b68, 32'h00000000} /* (19, 20, 22) {real, imag} */,
  {32'hc286d090, 32'h00000000} /* (19, 20, 21) {real, imag} */,
  {32'hc4ca3b93, 32'h00000000} /* (19, 20, 20) {real, imag} */,
  {32'hc4ee4f17, 32'h00000000} /* (19, 20, 19) {real, imag} */,
  {32'hc4de5300, 32'h00000000} /* (19, 20, 18) {real, imag} */,
  {32'hc518d678, 32'h00000000} /* (19, 20, 17) {real, imag} */,
  {32'hc4f0cb90, 32'h00000000} /* (19, 20, 16) {real, imag} */,
  {32'hc50fba23, 32'h00000000} /* (19, 20, 15) {real, imag} */,
  {32'hc4ffa174, 32'h00000000} /* (19, 20, 14) {real, imag} */,
  {32'hc532bdd8, 32'h00000000} /* (19, 20, 13) {real, imag} */,
  {32'hc54858bf, 32'h00000000} /* (19, 20, 12) {real, imag} */,
  {32'hc51bf750, 32'h00000000} /* (19, 20, 11) {real, imag} */,
  {32'h42419390, 32'h00000000} /* (19, 20, 10) {real, imag} */,
  {32'hc1be8780, 32'h00000000} /* (19, 20, 9) {real, imag} */,
  {32'h448239e6, 32'h00000000} /* (19, 20, 8) {real, imag} */,
  {32'h4472b212, 32'h00000000} /* (19, 20, 7) {real, imag} */,
  {32'h44dba5c8, 32'h00000000} /* (19, 20, 6) {real, imag} */,
  {32'h4500a264, 32'h00000000} /* (19, 20, 5) {real, imag} */,
  {32'h44870525, 32'h00000000} /* (19, 20, 4) {real, imag} */,
  {32'h450f6559, 32'h00000000} /* (19, 20, 3) {real, imag} */,
  {32'h4517d958, 32'h00000000} /* (19, 20, 2) {real, imag} */,
  {32'h44f9bcd0, 32'h00000000} /* (19, 20, 1) {real, imag} */,
  {32'h44c87bba, 32'h00000000} /* (19, 20, 0) {real, imag} */,
  {32'h457d97b2, 32'h00000000} /* (19, 19, 31) {real, imag} */,
  {32'h45867098, 32'h00000000} /* (19, 19, 30) {real, imag} */,
  {32'h4587b131, 32'h00000000} /* (19, 19, 29) {real, imag} */,
  {32'h45b7d732, 32'h00000000} /* (19, 19, 28) {real, imag} */,
  {32'h45afe5d4, 32'h00000000} /* (19, 19, 27) {real, imag} */,
  {32'h458c5334, 32'h00000000} /* (19, 19, 26) {real, imag} */,
  {32'h45852ef0, 32'h00000000} /* (19, 19, 25) {real, imag} */,
  {32'h45a78145, 32'h00000000} /* (19, 19, 24) {real, imag} */,
  {32'h45585371, 32'h00000000} /* (19, 19, 23) {real, imag} */,
  {32'h451b6500, 32'h00000000} /* (19, 19, 22) {real, imag} */,
  {32'h4421d72e, 32'h00000000} /* (19, 19, 21) {real, imag} */,
  {32'hc52405c8, 32'h00000000} /* (19, 19, 20) {real, imag} */,
  {32'hc58a8aa7, 32'h00000000} /* (19, 19, 19) {real, imag} */,
  {32'hc58c8f05, 32'h00000000} /* (19, 19, 18) {real, imag} */,
  {32'hc585efec, 32'h00000000} /* (19, 19, 17) {real, imag} */,
  {32'hc59a2d98, 32'h00000000} /* (19, 19, 16) {real, imag} */,
  {32'hc5a173df, 32'h00000000} /* (19, 19, 15) {real, imag} */,
  {32'hc578d6f8, 32'h00000000} /* (19, 19, 14) {real, imag} */,
  {32'hc56ae7e2, 32'h00000000} /* (19, 19, 13) {real, imag} */,
  {32'hc57daa0f, 32'h00000000} /* (19, 19, 12) {real, imag} */,
  {32'hc50c973e, 32'h00000000} /* (19, 19, 11) {real, imag} */,
  {32'hc405b64c, 32'h00000000} /* (19, 19, 10) {real, imag} */,
  {32'h44f48ce2, 32'h00000000} /* (19, 19, 9) {real, imag} */,
  {32'h454a6a5e, 32'h00000000} /* (19, 19, 8) {real, imag} */,
  {32'h4564fb6b, 32'h00000000} /* (19, 19, 7) {real, imag} */,
  {32'h4559c3bc, 32'h00000000} /* (19, 19, 6) {real, imag} */,
  {32'h4567467c, 32'h00000000} /* (19, 19, 5) {real, imag} */,
  {32'h4597d882, 32'h00000000} /* (19, 19, 4) {real, imag} */,
  {32'h458d8bb3, 32'h00000000} /* (19, 19, 3) {real, imag} */,
  {32'h45a105c1, 32'h00000000} /* (19, 19, 2) {real, imag} */,
  {32'h45a817c2, 32'h00000000} /* (19, 19, 1) {real, imag} */,
  {32'h459b7da4, 32'h00000000} /* (19, 19, 0) {real, imag} */,
  {32'h45c0c404, 32'h00000000} /* (19, 18, 31) {real, imag} */,
  {32'h45d6c909, 32'h00000000} /* (19, 18, 30) {real, imag} */,
  {32'h45b4b8de, 32'h00000000} /* (19, 18, 29) {real, imag} */,
  {32'h45bdf30e, 32'h00000000} /* (19, 18, 28) {real, imag} */,
  {32'h45b46e48, 32'h00000000} /* (19, 18, 27) {real, imag} */,
  {32'h45b85862, 32'h00000000} /* (19, 18, 26) {real, imag} */,
  {32'h45eccc68, 32'h00000000} /* (19, 18, 25) {real, imag} */,
  {32'h45d54510, 32'h00000000} /* (19, 18, 24) {real, imag} */,
  {32'h457c126e, 32'h00000000} /* (19, 18, 23) {real, imag} */,
  {32'h451b48cc, 32'h00000000} /* (19, 18, 22) {real, imag} */,
  {32'h44579bac, 32'h00000000} /* (19, 18, 21) {real, imag} */,
  {32'hc5212a5c, 32'h00000000} /* (19, 18, 20) {real, imag} */,
  {32'hc583e9ab, 32'h00000000} /* (19, 18, 19) {real, imag} */,
  {32'hc5b463ba, 32'h00000000} /* (19, 18, 18) {real, imag} */,
  {32'hc5d0157e, 32'h00000000} /* (19, 18, 17) {real, imag} */,
  {32'hc5d8eb6e, 32'h00000000} /* (19, 18, 16) {real, imag} */,
  {32'hc5d081ac, 32'h00000000} /* (19, 18, 15) {real, imag} */,
  {32'hc5b6a259, 32'h00000000} /* (19, 18, 14) {real, imag} */,
  {32'hc5978526, 32'h00000000} /* (19, 18, 13) {real, imag} */,
  {32'hc586bf34, 32'h00000000} /* (19, 18, 12) {real, imag} */,
  {32'hc526bfb8, 32'h00000000} /* (19, 18, 11) {real, imag} */,
  {32'h44a24c12, 32'h00000000} /* (19, 18, 10) {real, imag} */,
  {32'h4568759c, 32'h00000000} /* (19, 18, 9) {real, imag} */,
  {32'h456fd0b0, 32'h00000000} /* (19, 18, 8) {real, imag} */,
  {32'h45b25fb3, 32'h00000000} /* (19, 18, 7) {real, imag} */,
  {32'h45a5c142, 32'h00000000} /* (19, 18, 6) {real, imag} */,
  {32'h45baf5fe, 32'h00000000} /* (19, 18, 5) {real, imag} */,
  {32'h45e1821e, 32'h00000000} /* (19, 18, 4) {real, imag} */,
  {32'h45cc1f0d, 32'h00000000} /* (19, 18, 3) {real, imag} */,
  {32'h45c7a80c, 32'h00000000} /* (19, 18, 2) {real, imag} */,
  {32'h45d6f49c, 32'h00000000} /* (19, 18, 1) {real, imag} */,
  {32'h45e538ce, 32'h00000000} /* (19, 18, 0) {real, imag} */,
  {32'h45d7f6e5, 32'h00000000} /* (19, 17, 31) {real, imag} */,
  {32'h45e9c58f, 32'h00000000} /* (19, 17, 30) {real, imag} */,
  {32'h46001225, 32'h00000000} /* (19, 17, 29) {real, imag} */,
  {32'h45e5706d, 32'h00000000} /* (19, 17, 28) {real, imag} */,
  {32'h4601aa2b, 32'h00000000} /* (19, 17, 27) {real, imag} */,
  {32'h45edcc72, 32'h00000000} /* (19, 17, 26) {real, imag} */,
  {32'h45e2d677, 32'h00000000} /* (19, 17, 25) {real, imag} */,
  {32'h45c38ed6, 32'h00000000} /* (19, 17, 24) {real, imag} */,
  {32'h45a1f141, 32'h00000000} /* (19, 17, 23) {real, imag} */,
  {32'h45798c18, 32'h00000000} /* (19, 17, 22) {real, imag} */,
  {32'h43fff548, 32'h00000000} /* (19, 17, 21) {real, imag} */,
  {32'hc50228a2, 32'h00000000} /* (19, 17, 20) {real, imag} */,
  {32'hc591cbf3, 32'h00000000} /* (19, 17, 19) {real, imag} */,
  {32'hc5bba45e, 32'h00000000} /* (19, 17, 18) {real, imag} */,
  {32'hc5d33c40, 32'h00000000} /* (19, 17, 17) {real, imag} */,
  {32'hc602651a, 32'h00000000} /* (19, 17, 16) {real, imag} */,
  {32'hc5e49fb3, 32'h00000000} /* (19, 17, 15) {real, imag} */,
  {32'hc5be2d17, 32'h00000000} /* (19, 17, 14) {real, imag} */,
  {32'hc59fb9ec, 32'h00000000} /* (19, 17, 13) {real, imag} */,
  {32'hc592a267, 32'h00000000} /* (19, 17, 12) {real, imag} */,
  {32'hc523a538, 32'h00000000} /* (19, 17, 11) {real, imag} */,
  {32'h44c104c6, 32'h00000000} /* (19, 17, 10) {real, imag} */,
  {32'h45396f76, 32'h00000000} /* (19, 17, 9) {real, imag} */,
  {32'h45b7bfa0, 32'h00000000} /* (19, 17, 8) {real, imag} */,
  {32'h45c5f685, 32'h00000000} /* (19, 17, 7) {real, imag} */,
  {32'h45db9ce2, 32'h00000000} /* (19, 17, 6) {real, imag} */,
  {32'h45e50aaa, 32'h00000000} /* (19, 17, 5) {real, imag} */,
  {32'h46031da6, 32'h00000000} /* (19, 17, 4) {real, imag} */,
  {32'h45e39259, 32'h00000000} /* (19, 17, 3) {real, imag} */,
  {32'h45ff361e, 32'h00000000} /* (19, 17, 2) {real, imag} */,
  {32'h45ee0220, 32'h00000000} /* (19, 17, 1) {real, imag} */,
  {32'h45f463cb, 32'h00000000} /* (19, 17, 0) {real, imag} */,
  {32'h45fe776a, 32'h00000000} /* (19, 16, 31) {real, imag} */,
  {32'h45f4ec24, 32'h00000000} /* (19, 16, 30) {real, imag} */,
  {32'h460146ab, 32'h00000000} /* (19, 16, 29) {real, imag} */,
  {32'h460d0c51, 32'h00000000} /* (19, 16, 28) {real, imag} */,
  {32'h460f4bc5, 32'h00000000} /* (19, 16, 27) {real, imag} */,
  {32'h45fd6e2a, 32'h00000000} /* (19, 16, 26) {real, imag} */,
  {32'h45fdf875, 32'h00000000} /* (19, 16, 25) {real, imag} */,
  {32'h45e7e40c, 32'h00000000} /* (19, 16, 24) {real, imag} */,
  {32'h45a4b13e, 32'h00000000} /* (19, 16, 23) {real, imag} */,
  {32'h4555f4df, 32'h00000000} /* (19, 16, 22) {real, imag} */,
  {32'h443b5208, 32'h00000000} /* (19, 16, 21) {real, imag} */,
  {32'hc56425cf, 32'h00000000} /* (19, 16, 20) {real, imag} */,
  {32'hc59ec0cc, 32'h00000000} /* (19, 16, 19) {real, imag} */,
  {32'hc5cf2503, 32'h00000000} /* (19, 16, 18) {real, imag} */,
  {32'hc5e97808, 32'h00000000} /* (19, 16, 17) {real, imag} */,
  {32'hc5ea5732, 32'h00000000} /* (19, 16, 16) {real, imag} */,
  {32'hc5f811d2, 32'h00000000} /* (19, 16, 15) {real, imag} */,
  {32'hc5d916de, 32'h00000000} /* (19, 16, 14) {real, imag} */,
  {32'hc5ca672a, 32'h00000000} /* (19, 16, 13) {real, imag} */,
  {32'hc5898af0, 32'h00000000} /* (19, 16, 12) {real, imag} */,
  {32'hc542cf18, 32'h00000000} /* (19, 16, 11) {real, imag} */,
  {32'h4498ff7a, 32'h00000000} /* (19, 16, 10) {real, imag} */,
  {32'h4596f6cd, 32'h00000000} /* (19, 16, 9) {real, imag} */,
  {32'h45b4fe38, 32'h00000000} /* (19, 16, 8) {real, imag} */,
  {32'h45e73d80, 32'h00000000} /* (19, 16, 7) {real, imag} */,
  {32'h45edeb84, 32'h00000000} /* (19, 16, 6) {real, imag} */,
  {32'h45e31261, 32'h00000000} /* (19, 16, 5) {real, imag} */,
  {32'h45f677f0, 32'h00000000} /* (19, 16, 4) {real, imag} */,
  {32'h4600ae80, 32'h00000000} /* (19, 16, 3) {real, imag} */,
  {32'h45fe48b3, 32'h00000000} /* (19, 16, 2) {real, imag} */,
  {32'h45f2f1c8, 32'h00000000} /* (19, 16, 1) {real, imag} */,
  {32'h45d621aa, 32'h00000000} /* (19, 16, 0) {real, imag} */,
  {32'h45f3f286, 32'h00000000} /* (19, 15, 31) {real, imag} */,
  {32'h4604a3ce, 32'h00000000} /* (19, 15, 30) {real, imag} */,
  {32'h45fa1a83, 32'h00000000} /* (19, 15, 29) {real, imag} */,
  {32'h4609d213, 32'h00000000} /* (19, 15, 28) {real, imag} */,
  {32'h46024bf3, 32'h00000000} /* (19, 15, 27) {real, imag} */,
  {32'h460d4d38, 32'h00000000} /* (19, 15, 26) {real, imag} */,
  {32'h45fb73e1, 32'h00000000} /* (19, 15, 25) {real, imag} */,
  {32'h45ec2055, 32'h00000000} /* (19, 15, 24) {real, imag} */,
  {32'h45c971bf, 32'h00000000} /* (19, 15, 23) {real, imag} */,
  {32'h457333de, 32'h00000000} /* (19, 15, 22) {real, imag} */,
  {32'h4492812c, 32'h00000000} /* (19, 15, 21) {real, imag} */,
  {32'hc515e731, 32'h00000000} /* (19, 15, 20) {real, imag} */,
  {32'hc5b5d646, 32'h00000000} /* (19, 15, 19) {real, imag} */,
  {32'hc5d487d3, 32'h00000000} /* (19, 15, 18) {real, imag} */,
  {32'hc5db52fe, 32'h00000000} /* (19, 15, 17) {real, imag} */,
  {32'hc5dffc2e, 32'h00000000} /* (19, 15, 16) {real, imag} */,
  {32'hc5f7406e, 32'h00000000} /* (19, 15, 15) {real, imag} */,
  {32'hc5e9eb30, 32'h00000000} /* (19, 15, 14) {real, imag} */,
  {32'hc5c9a099, 32'h00000000} /* (19, 15, 13) {real, imag} */,
  {32'hc58176ae, 32'h00000000} /* (19, 15, 12) {real, imag} */,
  {32'hc545d418, 32'h00000000} /* (19, 15, 11) {real, imag} */,
  {32'h44e4fc40, 32'h00000000} /* (19, 15, 10) {real, imag} */,
  {32'h4596349b, 32'h00000000} /* (19, 15, 9) {real, imag} */,
  {32'h45deaaeb, 32'h00000000} /* (19, 15, 8) {real, imag} */,
  {32'h45fd7b39, 32'h00000000} /* (19, 15, 7) {real, imag} */,
  {32'h45ef3d11, 32'h00000000} /* (19, 15, 6) {real, imag} */,
  {32'h45fe3723, 32'h00000000} /* (19, 15, 5) {real, imag} */,
  {32'h45fb1960, 32'h00000000} /* (19, 15, 4) {real, imag} */,
  {32'h45fdbdae, 32'h00000000} /* (19, 15, 3) {real, imag} */,
  {32'h45f99e39, 32'h00000000} /* (19, 15, 2) {real, imag} */,
  {32'h45fa33a6, 32'h00000000} /* (19, 15, 1) {real, imag} */,
  {32'h45e2b570, 32'h00000000} /* (19, 15, 0) {real, imag} */,
  {32'h45cffa1a, 32'h00000000} /* (19, 14, 31) {real, imag} */,
  {32'h45de8470, 32'h00000000} /* (19, 14, 30) {real, imag} */,
  {32'h45eb1eab, 32'h00000000} /* (19, 14, 29) {real, imag} */,
  {32'h4604c080, 32'h00000000} /* (19, 14, 28) {real, imag} */,
  {32'h45e8abe1, 32'h00000000} /* (19, 14, 27) {real, imag} */,
  {32'h45ddeddd, 32'h00000000} /* (19, 14, 26) {real, imag} */,
  {32'h45da0ddb, 32'h00000000} /* (19, 14, 25) {real, imag} */,
  {32'h45dcf601, 32'h00000000} /* (19, 14, 24) {real, imag} */,
  {32'h45a329c6, 32'h00000000} /* (19, 14, 23) {real, imag} */,
  {32'h4584af61, 32'h00000000} /* (19, 14, 22) {real, imag} */,
  {32'h449abf0a, 32'h00000000} /* (19, 14, 21) {real, imag} */,
  {32'hc52fb348, 32'h00000000} /* (19, 14, 20) {real, imag} */,
  {32'hc5a1d350, 32'h00000000} /* (19, 14, 19) {real, imag} */,
  {32'hc5ada685, 32'h00000000} /* (19, 14, 18) {real, imag} */,
  {32'hc5d13900, 32'h00000000} /* (19, 14, 17) {real, imag} */,
  {32'hc5f40336, 32'h00000000} /* (19, 14, 16) {real, imag} */,
  {32'hc5f3cfc4, 32'h00000000} /* (19, 14, 15) {real, imag} */,
  {32'hc5e098da, 32'h00000000} /* (19, 14, 14) {real, imag} */,
  {32'hc5a8f533, 32'h00000000} /* (19, 14, 13) {real, imag} */,
  {32'hc578790a, 32'h00000000} /* (19, 14, 12) {real, imag} */,
  {32'hc4e5c744, 32'h00000000} /* (19, 14, 11) {real, imag} */,
  {32'h448fb574, 32'h00000000} /* (19, 14, 10) {real, imag} */,
  {32'h45849571, 32'h00000000} /* (19, 14, 9) {real, imag} */,
  {32'h45c4459f, 32'h00000000} /* (19, 14, 8) {real, imag} */,
  {32'h45d3da76, 32'h00000000} /* (19, 14, 7) {real, imag} */,
  {32'h45e61427, 32'h00000000} /* (19, 14, 6) {real, imag} */,
  {32'h45dec854, 32'h00000000} /* (19, 14, 5) {real, imag} */,
  {32'h45edc20c, 32'h00000000} /* (19, 14, 4) {real, imag} */,
  {32'h45f3d23c, 32'h00000000} /* (19, 14, 3) {real, imag} */,
  {32'h45e91035, 32'h00000000} /* (19, 14, 2) {real, imag} */,
  {32'h45df91f0, 32'h00000000} /* (19, 14, 1) {real, imag} */,
  {32'h45c9ac66, 32'h00000000} /* (19, 14, 0) {real, imag} */,
  {32'h45a8af74, 32'h00000000} /* (19, 13, 31) {real, imag} */,
  {32'h45d16e36, 32'h00000000} /* (19, 13, 30) {real, imag} */,
  {32'h45be59e5, 32'h00000000} /* (19, 13, 29) {real, imag} */,
  {32'h45e036f0, 32'h00000000} /* (19, 13, 28) {real, imag} */,
  {32'h45bbaa30, 32'h00000000} /* (19, 13, 27) {real, imag} */,
  {32'h45ab2749, 32'h00000000} /* (19, 13, 26) {real, imag} */,
  {32'h45ae5a4a, 32'h00000000} /* (19, 13, 25) {real, imag} */,
  {32'h4599017c, 32'h00000000} /* (19, 13, 24) {real, imag} */,
  {32'h45756fb6, 32'h00000000} /* (19, 13, 23) {real, imag} */,
  {32'h4525b326, 32'h00000000} /* (19, 13, 22) {real, imag} */,
  {32'h44da74da, 32'h00000000} /* (19, 13, 21) {real, imag} */,
  {32'hc540cf6d, 32'h00000000} /* (19, 13, 20) {real, imag} */,
  {32'hc57c3802, 32'h00000000} /* (19, 13, 19) {real, imag} */,
  {32'hc58c2650, 32'h00000000} /* (19, 13, 18) {real, imag} */,
  {32'hc5bda768, 32'h00000000} /* (19, 13, 17) {real, imag} */,
  {32'hc5bc8fe3, 32'h00000000} /* (19, 13, 16) {real, imag} */,
  {32'hc5d25e10, 32'h00000000} /* (19, 13, 15) {real, imag} */,
  {32'hc5cfa62a, 32'h00000000} /* (19, 13, 14) {real, imag} */,
  {32'hc5c3d8d3, 32'h00000000} /* (19, 13, 13) {real, imag} */,
  {32'hc5415261, 32'h00000000} /* (19, 13, 12) {real, imag} */,
  {32'hc484dc34, 32'h00000000} /* (19, 13, 11) {real, imag} */,
  {32'h44ebd0f1, 32'h00000000} /* (19, 13, 10) {real, imag} */,
  {32'h45737284, 32'h00000000} /* (19, 13, 9) {real, imag} */,
  {32'h45aec1e2, 32'h00000000} /* (19, 13, 8) {real, imag} */,
  {32'h45c47c99, 32'h00000000} /* (19, 13, 7) {real, imag} */,
  {32'h45c26035, 32'h00000000} /* (19, 13, 6) {real, imag} */,
  {32'h45ca3918, 32'h00000000} /* (19, 13, 5) {real, imag} */,
  {32'h45b68b16, 32'h00000000} /* (19, 13, 4) {real, imag} */,
  {32'h45babfc7, 32'h00000000} /* (19, 13, 3) {real, imag} */,
  {32'h45bcdff0, 32'h00000000} /* (19, 13, 2) {real, imag} */,
  {32'h45a9c714, 32'h00000000} /* (19, 13, 1) {real, imag} */,
  {32'h45b0223f, 32'h00000000} /* (19, 13, 0) {real, imag} */,
  {32'h454371b8, 32'h00000000} /* (19, 12, 31) {real, imag} */,
  {32'h4570e1c7, 32'h00000000} /* (19, 12, 30) {real, imag} */,
  {32'h45814c16, 32'h00000000} /* (19, 12, 29) {real, imag} */,
  {32'h45785e62, 32'h00000000} /* (19, 12, 28) {real, imag} */,
  {32'h457bd437, 32'h00000000} /* (19, 12, 27) {real, imag} */,
  {32'h4584029e, 32'h00000000} /* (19, 12, 26) {real, imag} */,
  {32'h455374fd, 32'h00000000} /* (19, 12, 25) {real, imag} */,
  {32'h45146244, 32'h00000000} /* (19, 12, 24) {real, imag} */,
  {32'h45590be0, 32'h00000000} /* (19, 12, 23) {real, imag} */,
  {32'h452b7a3d, 32'h00000000} /* (19, 12, 22) {real, imag} */,
  {32'h44c96086, 32'h00000000} /* (19, 12, 21) {real, imag} */,
  {32'hc4cff1a9, 32'h00000000} /* (19, 12, 20) {real, imag} */,
  {32'hc54c5f64, 32'h00000000} /* (19, 12, 19) {real, imag} */,
  {32'hc559a212, 32'h00000000} /* (19, 12, 18) {real, imag} */,
  {32'hc5ae8007, 32'h00000000} /* (19, 12, 17) {real, imag} */,
  {32'hc5937c4b, 32'h00000000} /* (19, 12, 16) {real, imag} */,
  {32'hc59686ce, 32'h00000000} /* (19, 12, 15) {real, imag} */,
  {32'hc5a4a62a, 32'h00000000} /* (19, 12, 14) {real, imag} */,
  {32'hc59236ac, 32'h00000000} /* (19, 12, 13) {real, imag} */,
  {32'hc5312924, 32'h00000000} /* (19, 12, 12) {real, imag} */,
  {32'hc31f03b0, 32'h00000000} /* (19, 12, 11) {real, imag} */,
  {32'h44f00c6e, 32'h00000000} /* (19, 12, 10) {real, imag} */,
  {32'h4560e1c7, 32'h00000000} /* (19, 12, 9) {real, imag} */,
  {32'h4599b7a2, 32'h00000000} /* (19, 12, 8) {real, imag} */,
  {32'h459d4ff6, 32'h00000000} /* (19, 12, 7) {real, imag} */,
  {32'h459b4f52, 32'h00000000} /* (19, 12, 6) {real, imag} */,
  {32'h4595a1c0, 32'h00000000} /* (19, 12, 5) {real, imag} */,
  {32'h457e07c4, 32'h00000000} /* (19, 12, 4) {real, imag} */,
  {32'h4591c896, 32'h00000000} /* (19, 12, 3) {real, imag} */,
  {32'h458594b4, 32'h00000000} /* (19, 12, 2) {real, imag} */,
  {32'h457c6302, 32'h00000000} /* (19, 12, 1) {real, imag} */,
  {32'h454daaae, 32'h00000000} /* (19, 12, 0) {real, imag} */,
  {32'h447b6c46, 32'h00000000} /* (19, 11, 31) {real, imag} */,
  {32'h44e977a2, 32'h00000000} /* (19, 11, 30) {real, imag} */,
  {32'h44977cd3, 32'h00000000} /* (19, 11, 29) {real, imag} */,
  {32'h44bc093e, 32'h00000000} /* (19, 11, 28) {real, imag} */,
  {32'h444404e7, 32'h00000000} /* (19, 11, 27) {real, imag} */,
  {32'h44450a7c, 32'h00000000} /* (19, 11, 26) {real, imag} */,
  {32'h44807a7d, 32'h00000000} /* (19, 11, 25) {real, imag} */,
  {32'h445a9160, 32'h00000000} /* (19, 11, 24) {real, imag} */,
  {32'h4404541c, 32'h00000000} /* (19, 11, 23) {real, imag} */,
  {32'h44b55e88, 32'h00000000} /* (19, 11, 22) {real, imag} */,
  {32'h43180de0, 32'h00000000} /* (19, 11, 21) {real, imag} */,
  {32'hc4b79722, 32'h00000000} /* (19, 11, 20) {real, imag} */,
  {32'hc51c827a, 32'h00000000} /* (19, 11, 19) {real, imag} */,
  {32'hc502db21, 32'h00000000} /* (19, 11, 18) {real, imag} */,
  {32'hc539220b, 32'h00000000} /* (19, 11, 17) {real, imag} */,
  {32'hc4c6b055, 32'h00000000} /* (19, 11, 16) {real, imag} */,
  {32'hc4fb9995, 32'h00000000} /* (19, 11, 15) {real, imag} */,
  {32'hc5319571, 32'h00000000} /* (19, 11, 14) {real, imag} */,
  {32'hc5130fe8, 32'h00000000} /* (19, 11, 13) {real, imag} */,
  {32'hc49d1fd4, 32'h00000000} /* (19, 11, 12) {real, imag} */,
  {32'h4496543e, 32'h00000000} /* (19, 11, 11) {real, imag} */,
  {32'h4505f19a, 32'h00000000} /* (19, 11, 10) {real, imag} */,
  {32'h45051d7c, 32'h00000000} /* (19, 11, 9) {real, imag} */,
  {32'h452aa2c9, 32'h00000000} /* (19, 11, 8) {real, imag} */,
  {32'h45237058, 32'h00000000} /* (19, 11, 7) {real, imag} */,
  {32'h453040c0, 32'h00000000} /* (19, 11, 6) {real, imag} */,
  {32'h45172f9f, 32'h00000000} /* (19, 11, 5) {real, imag} */,
  {32'h44ea3138, 32'h00000000} /* (19, 11, 4) {real, imag} */,
  {32'h4510e45a, 32'h00000000} /* (19, 11, 3) {real, imag} */,
  {32'h450eed3f, 32'h00000000} /* (19, 11, 2) {real, imag} */,
  {32'h44b7c5e2, 32'h00000000} /* (19, 11, 1) {real, imag} */,
  {32'h44a8d3a7, 32'h00000000} /* (19, 11, 0) {real, imag} */,
  {32'hc51dd336, 32'h00000000} /* (19, 10, 31) {real, imag} */,
  {32'hc50cc2ce, 32'h00000000} /* (19, 10, 30) {real, imag} */,
  {32'hc50e72e0, 32'h00000000} /* (19, 10, 29) {real, imag} */,
  {32'hc54757f4, 32'h00000000} /* (19, 10, 28) {real, imag} */,
  {32'hc5553be8, 32'h00000000} /* (19, 10, 27) {real, imag} */,
  {32'hc54e55e8, 32'h00000000} /* (19, 10, 26) {real, imag} */,
  {32'hc5444da2, 32'h00000000} /* (19, 10, 25) {real, imag} */,
  {32'hc57dae65, 32'h00000000} /* (19, 10, 24) {real, imag} */,
  {32'hc54b6771, 32'h00000000} /* (19, 10, 23) {real, imag} */,
  {32'hc512a720, 32'h00000000} /* (19, 10, 22) {real, imag} */,
  {32'hc4ba105e, 32'h00000000} /* (19, 10, 21) {real, imag} */,
  {32'hc42f4b28, 32'h00000000} /* (19, 10, 20) {real, imag} */,
  {32'h43ef083e, 32'h00000000} /* (19, 10, 19) {real, imag} */,
  {32'h43a66f40, 32'h00000000} /* (19, 10, 18) {real, imag} */,
  {32'h43898246, 32'h00000000} /* (19, 10, 17) {real, imag} */,
  {32'h44f5fcfd, 32'h00000000} /* (19, 10, 16) {real, imag} */,
  {32'h45231c88, 32'h00000000} /* (19, 10, 15) {real, imag} */,
  {32'h44d01b1c, 32'h00000000} /* (19, 10, 14) {real, imag} */,
  {32'h4426f598, 32'h00000000} /* (19, 10, 13) {real, imag} */,
  {32'h450685e6, 32'h00000000} /* (19, 10, 12) {real, imag} */,
  {32'h44c34f90, 32'h00000000} /* (19, 10, 11) {real, imag} */,
  {32'h44b30fa7, 32'h00000000} /* (19, 10, 10) {real, imag} */,
  {32'hc32d4080, 32'h00000000} /* (19, 10, 9) {real, imag} */,
  {32'hc3883278, 32'h00000000} /* (19, 10, 8) {real, imag} */,
  {32'h42918e20, 32'h00000000} /* (19, 10, 7) {real, imag} */,
  {32'hc4076f55, 32'h00000000} /* (19, 10, 6) {real, imag} */,
  {32'hc4a080f6, 32'h00000000} /* (19, 10, 5) {real, imag} */,
  {32'hc477bf1c, 32'h00000000} /* (19, 10, 4) {real, imag} */,
  {32'hc4bf2b42, 32'h00000000} /* (19, 10, 3) {real, imag} */,
  {32'hc4d6a008, 32'h00000000} /* (19, 10, 2) {real, imag} */,
  {32'hc4d3fa4e, 32'h00000000} /* (19, 10, 1) {real, imag} */,
  {32'hc4fa2325, 32'h00000000} /* (19, 10, 0) {real, imag} */,
  {32'hc5958a50, 32'h00000000} /* (19, 9, 31) {real, imag} */,
  {32'hc5b6dfb8, 32'h00000000} /* (19, 9, 30) {real, imag} */,
  {32'hc5aabf41, 32'h00000000} /* (19, 9, 29) {real, imag} */,
  {32'hc5e16527, 32'h00000000} /* (19, 9, 28) {real, imag} */,
  {32'hc5c02579, 32'h00000000} /* (19, 9, 27) {real, imag} */,
  {32'hc5c346f1, 32'h00000000} /* (19, 9, 26) {real, imag} */,
  {32'hc5c27450, 32'h00000000} /* (19, 9, 25) {real, imag} */,
  {32'hc5ac67da, 32'h00000000} /* (19, 9, 24) {real, imag} */,
  {32'hc5b4f23a, 32'h00000000} /* (19, 9, 23) {real, imag} */,
  {32'hc584252d, 32'h00000000} /* (19, 9, 22) {real, imag} */,
  {32'hc52af2a7, 32'h00000000} /* (19, 9, 21) {real, imag} */,
  {32'h42d06280, 32'h00000000} /* (19, 9, 20) {real, imag} */,
  {32'h4444ea5c, 32'h00000000} /* (19, 9, 19) {real, imag} */,
  {32'h45002716, 32'h00000000} /* (19, 9, 18) {real, imag} */,
  {32'h458288ce, 32'h00000000} /* (19, 9, 17) {real, imag} */,
  {32'h457f6c48, 32'h00000000} /* (19, 9, 16) {real, imag} */,
  {32'h45ca0b1c, 32'h00000000} /* (19, 9, 15) {real, imag} */,
  {32'h4597c2a0, 32'h00000000} /* (19, 9, 14) {real, imag} */,
  {32'h454142e6, 32'h00000000} /* (19, 9, 13) {real, imag} */,
  {32'h45653a0a, 32'h00000000} /* (19, 9, 12) {real, imag} */,
  {32'h4516a5ee, 32'h00000000} /* (19, 9, 11) {real, imag} */,
  {32'h42ba3b80, 32'h00000000} /* (19, 9, 10) {real, imag} */,
  {32'hc5012f37, 32'h00000000} /* (19, 9, 9) {real, imag} */,
  {32'hc4865c5e, 32'h00000000} /* (19, 9, 8) {real, imag} */,
  {32'hc4eec9eb, 32'h00000000} /* (19, 9, 7) {real, imag} */,
  {32'hc55a90c0, 32'h00000000} /* (19, 9, 6) {real, imag} */,
  {32'hc55e4161, 32'h00000000} /* (19, 9, 5) {real, imag} */,
  {32'hc58b7a33, 32'h00000000} /* (19, 9, 4) {real, imag} */,
  {32'hc581b68a, 32'h00000000} /* (19, 9, 3) {real, imag} */,
  {32'hc58a33da, 32'h00000000} /* (19, 9, 2) {real, imag} */,
  {32'hc599e468, 32'h00000000} /* (19, 9, 1) {real, imag} */,
  {32'hc59b238c, 32'h00000000} /* (19, 9, 0) {real, imag} */,
  {32'hc5da8f52, 32'h00000000} /* (19, 8, 31) {real, imag} */,
  {32'hc5feabd2, 32'h00000000} /* (19, 8, 30) {real, imag} */,
  {32'hc606f8de, 32'h00000000} /* (19, 8, 29) {real, imag} */,
  {32'hc5fbfde4, 32'h00000000} /* (19, 8, 28) {real, imag} */,
  {32'hc60a42ed, 32'h00000000} /* (19, 8, 27) {real, imag} */,
  {32'hc603b67d, 32'h00000000} /* (19, 8, 26) {real, imag} */,
  {32'hc5eba33e, 32'h00000000} /* (19, 8, 25) {real, imag} */,
  {32'hc5f25570, 32'h00000000} /* (19, 8, 24) {real, imag} */,
  {32'hc5dc9454, 32'h00000000} /* (19, 8, 23) {real, imag} */,
  {32'hc5b6f84a, 32'h00000000} /* (19, 8, 22) {real, imag} */,
  {32'hc555d9a0, 32'h00000000} /* (19, 8, 21) {real, imag} */,
  {32'hc3650090, 32'h00000000} /* (19, 8, 20) {real, imag} */,
  {32'h44b87a2e, 32'h00000000} /* (19, 8, 19) {real, imag} */,
  {32'h453e009c, 32'h00000000} /* (19, 8, 18) {real, imag} */,
  {32'h457ecbfc, 32'h00000000} /* (19, 8, 17) {real, imag} */,
  {32'h4588eace, 32'h00000000} /* (19, 8, 16) {real, imag} */,
  {32'h45b7cb3e, 32'h00000000} /* (19, 8, 15) {real, imag} */,
  {32'h45bafe52, 32'h00000000} /* (19, 8, 14) {real, imag} */,
  {32'h459cc5d6, 32'h00000000} /* (19, 8, 13) {real, imag} */,
  {32'h4581689e, 32'h00000000} /* (19, 8, 12) {real, imag} */,
  {32'h45724ee1, 32'h00000000} /* (19, 8, 11) {real, imag} */,
  {32'hc373f980, 32'h00000000} /* (19, 8, 10) {real, imag} */,
  {32'hc4ba4aca, 32'h00000000} /* (19, 8, 9) {real, imag} */,
  {32'hc4acf18e, 32'h00000000} /* (19, 8, 8) {real, imag} */,
  {32'hc5500cf8, 32'h00000000} /* (19, 8, 7) {real, imag} */,
  {32'hc593a858, 32'h00000000} /* (19, 8, 6) {real, imag} */,
  {32'hc590ed0c, 32'h00000000} /* (19, 8, 5) {real, imag} */,
  {32'hc5a1aa76, 32'h00000000} /* (19, 8, 4) {real, imag} */,
  {32'hc5d307fc, 32'h00000000} /* (19, 8, 3) {real, imag} */,
  {32'hc5c49ba2, 32'h00000000} /* (19, 8, 2) {real, imag} */,
  {32'hc5e2fe84, 32'h00000000} /* (19, 8, 1) {real, imag} */,
  {32'hc5e2f3c4, 32'h00000000} /* (19, 8, 0) {real, imag} */,
  {32'hc61580a3, 32'h00000000} /* (19, 7, 31) {real, imag} */,
  {32'hc614ab9a, 32'h00000000} /* (19, 7, 30) {real, imag} */,
  {32'hc61c9237, 32'h00000000} /* (19, 7, 29) {real, imag} */,
  {32'hc616b190, 32'h00000000} /* (19, 7, 28) {real, imag} */,
  {32'hc61c199c, 32'h00000000} /* (19, 7, 27) {real, imag} */,
  {32'hc6127fb4, 32'h00000000} /* (19, 7, 26) {real, imag} */,
  {32'hc61b5140, 32'h00000000} /* (19, 7, 25) {real, imag} */,
  {32'hc621dbec, 32'h00000000} /* (19, 7, 24) {real, imag} */,
  {32'hc5ef88fc, 32'h00000000} /* (19, 7, 23) {real, imag} */,
  {32'hc5e70222, 32'h00000000} /* (19, 7, 22) {real, imag} */,
  {32'hc5c7b534, 32'h00000000} /* (19, 7, 21) {real, imag} */,
  {32'hc4e4d228, 32'h00000000} /* (19, 7, 20) {real, imag} */,
  {32'h44822cea, 32'h00000000} /* (19, 7, 19) {real, imag} */,
  {32'h45237dea, 32'h00000000} /* (19, 7, 18) {real, imag} */,
  {32'h4589cc4e, 32'h00000000} /* (19, 7, 17) {real, imag} */,
  {32'h4597d6f9, 32'h00000000} /* (19, 7, 16) {real, imag} */,
  {32'h45c46120, 32'h00000000} /* (19, 7, 15) {real, imag} */,
  {32'h45cfe735, 32'h00000000} /* (19, 7, 14) {real, imag} */,
  {32'h45b6aeae, 32'h00000000} /* (19, 7, 13) {real, imag} */,
  {32'h459d7db2, 32'h00000000} /* (19, 7, 12) {real, imag} */,
  {32'h45892776, 32'h00000000} /* (19, 7, 11) {real, imag} */,
  {32'h448f6f14, 32'h00000000} /* (19, 7, 10) {real, imag} */,
  {32'hc3fb8780, 32'h00000000} /* (19, 7, 9) {real, imag} */,
  {32'hc5096778, 32'h00000000} /* (19, 7, 8) {real, imag} */,
  {32'hc5757247, 32'h00000000} /* (19, 7, 7) {real, imag} */,
  {32'hc591406c, 32'h00000000} /* (19, 7, 6) {real, imag} */,
  {32'hc5b5e6f4, 32'h00000000} /* (19, 7, 5) {real, imag} */,
  {32'hc5db1414, 32'h00000000} /* (19, 7, 4) {real, imag} */,
  {32'hc5dacf58, 32'h00000000} /* (19, 7, 3) {real, imag} */,
  {32'hc6021a4e, 32'h00000000} /* (19, 7, 2) {real, imag} */,
  {32'hc5f9db00, 32'h00000000} /* (19, 7, 1) {real, imag} */,
  {32'hc601c056, 32'h00000000} /* (19, 7, 0) {real, imag} */,
  {32'hc6114721, 32'h00000000} /* (19, 6, 31) {real, imag} */,
  {32'hc61e90af, 32'h00000000} /* (19, 6, 30) {real, imag} */,
  {32'hc628ee6d, 32'h00000000} /* (19, 6, 29) {real, imag} */,
  {32'hc624d1e3, 32'h00000000} /* (19, 6, 28) {real, imag} */,
  {32'hc614276a, 32'h00000000} /* (19, 6, 27) {real, imag} */,
  {32'hc62bbe1c, 32'h00000000} /* (19, 6, 26) {real, imag} */,
  {32'hc62c0b40, 32'h00000000} /* (19, 6, 25) {real, imag} */,
  {32'hc62023e2, 32'h00000000} /* (19, 6, 24) {real, imag} */,
  {32'hc6021cf8, 32'h00000000} /* (19, 6, 23) {real, imag} */,
  {32'hc5f7bbae, 32'h00000000} /* (19, 6, 22) {real, imag} */,
  {32'hc5c9a7c0, 32'h00000000} /* (19, 6, 21) {real, imag} */,
  {32'hc52cb9f4, 32'h00000000} /* (19, 6, 20) {real, imag} */,
  {32'hc42edfb8, 32'h00000000} /* (19, 6, 19) {real, imag} */,
  {32'h44e6d100, 32'h00000000} /* (19, 6, 18) {real, imag} */,
  {32'h454a6ed4, 32'h00000000} /* (19, 6, 17) {real, imag} */,
  {32'h459033f1, 32'h00000000} /* (19, 6, 16) {real, imag} */,
  {32'h45b2c436, 32'h00000000} /* (19, 6, 15) {real, imag} */,
  {32'h45e9fc4e, 32'h00000000} /* (19, 6, 14) {real, imag} */,
  {32'h45c06556, 32'h00000000} /* (19, 6, 13) {real, imag} */,
  {32'h45b29992, 32'h00000000} /* (19, 6, 12) {real, imag} */,
  {32'h458c4eab, 32'h00000000} /* (19, 6, 11) {real, imag} */,
  {32'h4517b042, 32'h00000000} /* (19, 6, 10) {real, imag} */,
  {32'h441e80d8, 32'h00000000} /* (19, 6, 9) {real, imag} */,
  {32'hc4bff234, 32'h00000000} /* (19, 6, 8) {real, imag} */,
  {32'hc50eef6e, 32'h00000000} /* (19, 6, 7) {real, imag} */,
  {32'hc59dd056, 32'h00000000} /* (19, 6, 6) {real, imag} */,
  {32'hc5bd70a4, 32'h00000000} /* (19, 6, 5) {real, imag} */,
  {32'hc5d91bc2, 32'h00000000} /* (19, 6, 4) {real, imag} */,
  {32'hc606873a, 32'h00000000} /* (19, 6, 3) {real, imag} */,
  {32'hc60de366, 32'h00000000} /* (19, 6, 2) {real, imag} */,
  {32'hc6179103, 32'h00000000} /* (19, 6, 1) {real, imag} */,
  {32'hc60d1e24, 32'h00000000} /* (19, 6, 0) {real, imag} */,
  {32'hc6236004, 32'h00000000} /* (19, 5, 31) {real, imag} */,
  {32'hc637a107, 32'h00000000} /* (19, 5, 30) {real, imag} */,
  {32'hc637f01e, 32'h00000000} /* (19, 5, 29) {real, imag} */,
  {32'hc62edfd6, 32'h00000000} /* (19, 5, 28) {real, imag} */,
  {32'hc62d688c, 32'h00000000} /* (19, 5, 27) {real, imag} */,
  {32'hc61ded84, 32'h00000000} /* (19, 5, 26) {real, imag} */,
  {32'hc6227f09, 32'h00000000} /* (19, 5, 25) {real, imag} */,
  {32'hc634691f, 32'h00000000} /* (19, 5, 24) {real, imag} */,
  {32'hc6195ec0, 32'h00000000} /* (19, 5, 23) {real, imag} */,
  {32'hc604bb16, 32'h00000000} /* (19, 5, 22) {real, imag} */,
  {32'hc5bdaa38, 32'h00000000} /* (19, 5, 21) {real, imag} */,
  {32'hc58206b3, 32'h00000000} /* (19, 5, 20) {real, imag} */,
  {32'hc508f520, 32'h00000000} /* (19, 5, 19) {real, imag} */,
  {32'hc4e920d0, 32'h00000000} /* (19, 5, 18) {real, imag} */,
  {32'h44239618, 32'h00000000} /* (19, 5, 17) {real, imag} */,
  {32'h454338ae, 32'h00000000} /* (19, 5, 16) {real, imag} */,
  {32'h458da0c7, 32'h00000000} /* (19, 5, 15) {real, imag} */,
  {32'h45c0438a, 32'h00000000} /* (19, 5, 14) {real, imag} */,
  {32'h45b48714, 32'h00000000} /* (19, 5, 13) {real, imag} */,
  {32'h45d3cf23, 32'h00000000} /* (19, 5, 12) {real, imag} */,
  {32'h45bd0959, 32'h00000000} /* (19, 5, 11) {real, imag} */,
  {32'h45a88a1b, 32'h00000000} /* (19, 5, 10) {real, imag} */,
  {32'h45318853, 32'h00000000} /* (19, 5, 9) {real, imag} */,
  {32'h44d40b88, 32'h00000000} /* (19, 5, 8) {real, imag} */,
  {32'hc4005500, 32'h00000000} /* (19, 5, 7) {real, imag} */,
  {32'hc4d7221e, 32'h00000000} /* (19, 5, 6) {real, imag} */,
  {32'hc5ae8e74, 32'h00000000} /* (19, 5, 5) {real, imag} */,
  {32'hc5f44883, 32'h00000000} /* (19, 5, 4) {real, imag} */,
  {32'hc6061ed0, 32'h00000000} /* (19, 5, 3) {real, imag} */,
  {32'hc621049a, 32'h00000000} /* (19, 5, 2) {real, imag} */,
  {32'hc6228894, 32'h00000000} /* (19, 5, 1) {real, imag} */,
  {32'hc61441fa, 32'h00000000} /* (19, 5, 0) {real, imag} */,
  {32'hc6347bd8, 32'h00000000} /* (19, 4, 31) {real, imag} */,
  {32'hc63b3b61, 32'h00000000} /* (19, 4, 30) {real, imag} */,
  {32'hc64223fa, 32'h00000000} /* (19, 4, 29) {real, imag} */,
  {32'hc639dca8, 32'h00000000} /* (19, 4, 28) {real, imag} */,
  {32'hc63abcbb, 32'h00000000} /* (19, 4, 27) {real, imag} */,
  {32'hc62b990e, 32'h00000000} /* (19, 4, 26) {real, imag} */,
  {32'hc6265c0e, 32'h00000000} /* (19, 4, 25) {real, imag} */,
  {32'hc63002a8, 32'h00000000} /* (19, 4, 24) {real, imag} */,
  {32'hc62aefb9, 32'h00000000} /* (19, 4, 23) {real, imag} */,
  {32'hc60cd964, 32'h00000000} /* (19, 4, 22) {real, imag} */,
  {32'hc60dc29f, 32'h00000000} /* (19, 4, 21) {real, imag} */,
  {32'hc5ccbc07, 32'h00000000} /* (19, 4, 20) {real, imag} */,
  {32'hc59f25c2, 32'h00000000} /* (19, 4, 19) {real, imag} */,
  {32'hc57eb291, 32'h00000000} /* (19, 4, 18) {real, imag} */,
  {32'hc4cbe1e4, 32'h00000000} /* (19, 4, 17) {real, imag} */,
  {32'h44056ee0, 32'h00000000} /* (19, 4, 16) {real, imag} */,
  {32'h45672ba3, 32'h00000000} /* (19, 4, 15) {real, imag} */,
  {32'h45c1eefe, 32'h00000000} /* (19, 4, 14) {real, imag} */,
  {32'h45c16edc, 32'h00000000} /* (19, 4, 13) {real, imag} */,
  {32'h45cfea58, 32'h00000000} /* (19, 4, 12) {real, imag} */,
  {32'h45d7007a, 32'h00000000} /* (19, 4, 11) {real, imag} */,
  {32'h45b57a89, 32'h00000000} /* (19, 4, 10) {real, imag} */,
  {32'h45a06fa8, 32'h00000000} /* (19, 4, 9) {real, imag} */,
  {32'h45786ff5, 32'h00000000} /* (19, 4, 8) {real, imag} */,
  {32'h448b0d80, 32'h00000000} /* (19, 4, 7) {real, imag} */,
  {32'hc3f02900, 32'h00000000} /* (19, 4, 6) {real, imag} */,
  {32'hc599b772, 32'h00000000} /* (19, 4, 5) {real, imag} */,
  {32'hc5f1a159, 32'h00000000} /* (19, 4, 4) {real, imag} */,
  {32'hc60a6f25, 32'h00000000} /* (19, 4, 3) {real, imag} */,
  {32'hc61706e7, 32'h00000000} /* (19, 4, 2) {real, imag} */,
  {32'hc62092ea, 32'h00000000} /* (19, 4, 1) {real, imag} */,
  {32'hc6193117, 32'h00000000} /* (19, 4, 0) {real, imag} */,
  {32'hc62752e1, 32'h00000000} /* (19, 3, 31) {real, imag} */,
  {32'hc63056fe, 32'h00000000} /* (19, 3, 30) {real, imag} */,
  {32'hc63a3568, 32'h00000000} /* (19, 3, 29) {real, imag} */,
  {32'hc633868b, 32'h00000000} /* (19, 3, 28) {real, imag} */,
  {32'hc63343c0, 32'h00000000} /* (19, 3, 27) {real, imag} */,
  {32'hc6392ea7, 32'h00000000} /* (19, 3, 26) {real, imag} */,
  {32'hc62e1c74, 32'h00000000} /* (19, 3, 25) {real, imag} */,
  {32'hc6366c30, 32'h00000000} /* (19, 3, 24) {real, imag} */,
  {32'hc635289c, 32'h00000000} /* (19, 3, 23) {real, imag} */,
  {32'hc62a5d2e, 32'h00000000} /* (19, 3, 22) {real, imag} */,
  {32'hc6071ad7, 32'h00000000} /* (19, 3, 21) {real, imag} */,
  {32'hc5f5c850, 32'h00000000} /* (19, 3, 20) {real, imag} */,
  {32'hc5def874, 32'h00000000} /* (19, 3, 19) {real, imag} */,
  {32'hc5748c69, 32'h00000000} /* (19, 3, 18) {real, imag} */,
  {32'hc5163d5a, 32'h00000000} /* (19, 3, 17) {real, imag} */,
  {32'h43da45c0, 32'h00000000} /* (19, 3, 16) {real, imag} */,
  {32'h453cdb67, 32'h00000000} /* (19, 3, 15) {real, imag} */,
  {32'h45a44508, 32'h00000000} /* (19, 3, 14) {real, imag} */,
  {32'h45d40198, 32'h00000000} /* (19, 3, 13) {real, imag} */,
  {32'h45d8c64e, 32'h00000000} /* (19, 3, 12) {real, imag} */,
  {32'h45d3641c, 32'h00000000} /* (19, 3, 11) {real, imag} */,
  {32'h45beeefa, 32'h00000000} /* (19, 3, 10) {real, imag} */,
  {32'h45b13898, 32'h00000000} /* (19, 3, 9) {real, imag} */,
  {32'h459b05ed, 32'h00000000} /* (19, 3, 8) {real, imag} */,
  {32'h453da326, 32'h00000000} /* (19, 3, 7) {real, imag} */,
  {32'hc3f9ac80, 32'h00000000} /* (19, 3, 6) {real, imag} */,
  {32'hc58b6686, 32'h00000000} /* (19, 3, 5) {real, imag} */,
  {32'hc5e7a504, 32'h00000000} /* (19, 3, 4) {real, imag} */,
  {32'hc607ce2e, 32'h00000000} /* (19, 3, 3) {real, imag} */,
  {32'hc61d8680, 32'h00000000} /* (19, 3, 2) {real, imag} */,
  {32'hc626c2b0, 32'h00000000} /* (19, 3, 1) {real, imag} */,
  {32'hc6218bef, 32'h00000000} /* (19, 3, 0) {real, imag} */,
  {32'hc62af0f5, 32'h00000000} /* (19, 2, 31) {real, imag} */,
  {32'hc6428bb6, 32'h00000000} /* (19, 2, 30) {real, imag} */,
  {32'hc630e5e3, 32'h00000000} /* (19, 2, 29) {real, imag} */,
  {32'hc630e6fe, 32'h00000000} /* (19, 2, 28) {real, imag} */,
  {32'hc639346c, 32'h00000000} /* (19, 2, 27) {real, imag} */,
  {32'hc62f60b0, 32'h00000000} /* (19, 2, 26) {real, imag} */,
  {32'hc632dc3c, 32'h00000000} /* (19, 2, 25) {real, imag} */,
  {32'hc62d65ec, 32'h00000000} /* (19, 2, 24) {real, imag} */,
  {32'hc63e278a, 32'h00000000} /* (19, 2, 23) {real, imag} */,
  {32'hc6250cc1, 32'h00000000} /* (19, 2, 22) {real, imag} */,
  {32'hc5e12afe, 32'h00000000} /* (19, 2, 21) {real, imag} */,
  {32'hc5dc16b9, 32'h00000000} /* (19, 2, 20) {real, imag} */,
  {32'hc5d1ac9c, 32'h00000000} /* (19, 2, 19) {real, imag} */,
  {32'hc5b0fe08, 32'h00000000} /* (19, 2, 18) {real, imag} */,
  {32'hc5343420, 32'h00000000} /* (19, 2, 17) {real, imag} */,
  {32'h43f38750, 32'h00000000} /* (19, 2, 16) {real, imag} */,
  {32'h451e7724, 32'h00000000} /* (19, 2, 15) {real, imag} */,
  {32'h45986734, 32'h00000000} /* (19, 2, 14) {real, imag} */,
  {32'h45c20a36, 32'h00000000} /* (19, 2, 13) {real, imag} */,
  {32'h45cbcf34, 32'h00000000} /* (19, 2, 12) {real, imag} */,
  {32'h45b539a8, 32'h00000000} /* (19, 2, 11) {real, imag} */,
  {32'h45a233c4, 32'h00000000} /* (19, 2, 10) {real, imag} */,
  {32'h45ada8df, 32'h00000000} /* (19, 2, 9) {real, imag} */,
  {32'h456ed736, 32'h00000000} /* (19, 2, 8) {real, imag} */,
  {32'h450a9d82, 32'h00000000} /* (19, 2, 7) {real, imag} */,
  {32'hc434ed50, 32'h00000000} /* (19, 2, 6) {real, imag} */,
  {32'hc57c89dc, 32'h00000000} /* (19, 2, 5) {real, imag} */,
  {32'hc5d86f4f, 32'h00000000} /* (19, 2, 4) {real, imag} */,
  {32'hc6173d90, 32'h00000000} /* (19, 2, 3) {real, imag} */,
  {32'hc62d4d4c, 32'h00000000} /* (19, 2, 2) {real, imag} */,
  {32'hc62d13c9, 32'h00000000} /* (19, 2, 1) {real, imag} */,
  {32'hc61d9cac, 32'h00000000} /* (19, 2, 0) {real, imag} */,
  {32'hc628ee66, 32'h00000000} /* (19, 1, 31) {real, imag} */,
  {32'hc63204f2, 32'h00000000} /* (19, 1, 30) {real, imag} */,
  {32'hc641fb1c, 32'h00000000} /* (19, 1, 29) {real, imag} */,
  {32'hc642b1f9, 32'h00000000} /* (19, 1, 28) {real, imag} */,
  {32'hc6396863, 32'h00000000} /* (19, 1, 27) {real, imag} */,
  {32'hc637c18e, 32'h00000000} /* (19, 1, 26) {real, imag} */,
  {32'hc62e38ae, 32'h00000000} /* (19, 1, 25) {real, imag} */,
  {32'hc627f495, 32'h00000000} /* (19, 1, 24) {real, imag} */,
  {32'hc62a3ef2, 32'h00000000} /* (19, 1, 23) {real, imag} */,
  {32'hc60ffa13, 32'h00000000} /* (19, 1, 22) {real, imag} */,
  {32'hc5ee2d9d, 32'h00000000} /* (19, 1, 21) {real, imag} */,
  {32'hc5bc7893, 32'h00000000} /* (19, 1, 20) {real, imag} */,
  {32'hc59c93a3, 32'h00000000} /* (19, 1, 19) {real, imag} */,
  {32'hc58b2a76, 32'h00000000} /* (19, 1, 18) {real, imag} */,
  {32'hc548a456, 32'h00000000} /* (19, 1, 17) {real, imag} */,
  {32'h445fe710, 32'h00000000} /* (19, 1, 16) {real, imag} */,
  {32'h4577d56d, 32'h00000000} /* (19, 1, 15) {real, imag} */,
  {32'h459b90ef, 32'h00000000} /* (19, 1, 14) {real, imag} */,
  {32'h45a88fbf, 32'h00000000} /* (19, 1, 13) {real, imag} */,
  {32'h45b3a8d6, 32'h00000000} /* (19, 1, 12) {real, imag} */,
  {32'h45b7f6f2, 32'h00000000} /* (19, 1, 11) {real, imag} */,
  {32'h45a0c658, 32'h00000000} /* (19, 1, 10) {real, imag} */,
  {32'h4570e082, 32'h00000000} /* (19, 1, 9) {real, imag} */,
  {32'h4513f648, 32'h00000000} /* (19, 1, 8) {real, imag} */,
  {32'h4459f870, 32'h00000000} /* (19, 1, 7) {real, imag} */,
  {32'hc4dc5576, 32'h00000000} /* (19, 1, 6) {real, imag} */,
  {32'hc564b572, 32'h00000000} /* (19, 1, 5) {real, imag} */,
  {32'hc5e63c81, 32'h00000000} /* (19, 1, 4) {real, imag} */,
  {32'hc622fa0e, 32'h00000000} /* (19, 1, 3) {real, imag} */,
  {32'hc6214857, 32'h00000000} /* (19, 1, 2) {real, imag} */,
  {32'hc62d6a4c, 32'h00000000} /* (19, 1, 1) {real, imag} */,
  {32'hc6272e1e, 32'h00000000} /* (19, 1, 0) {real, imag} */,
  {32'hc633775b, 32'h00000000} /* (19, 0, 31) {real, imag} */,
  {32'hc62e59d5, 32'h00000000} /* (19, 0, 30) {real, imag} */,
  {32'hc634ad59, 32'h00000000} /* (19, 0, 29) {real, imag} */,
  {32'hc63d445d, 32'h00000000} /* (19, 0, 28) {real, imag} */,
  {32'hc632dd2e, 32'h00000000} /* (19, 0, 27) {real, imag} */,
  {32'hc6323986, 32'h00000000} /* (19, 0, 26) {real, imag} */,
  {32'hc62e7e4b, 32'h00000000} /* (19, 0, 25) {real, imag} */,
  {32'hc62354d2, 32'h00000000} /* (19, 0, 24) {real, imag} */,
  {32'hc60dc64c, 32'h00000000} /* (19, 0, 23) {real, imag} */,
  {32'hc5f6ed80, 32'h00000000} /* (19, 0, 22) {real, imag} */,
  {32'hc5d0cf20, 32'h00000000} /* (19, 0, 21) {real, imag} */,
  {32'hc596a7ff, 32'h00000000} /* (19, 0, 20) {real, imag} */,
  {32'hc5537c54, 32'h00000000} /* (19, 0, 19) {real, imag} */,
  {32'hc4b27e60, 32'h00000000} /* (19, 0, 18) {real, imag} */,
  {32'hc1fb3400, 32'h00000000} /* (19, 0, 17) {real, imag} */,
  {32'h4503c2c0, 32'h00000000} /* (19, 0, 16) {real, imag} */,
  {32'h4581ec44, 32'h00000000} /* (19, 0, 15) {real, imag} */,
  {32'h4599b3f2, 32'h00000000} /* (19, 0, 14) {real, imag} */,
  {32'h45a81dca, 32'h00000000} /* (19, 0, 13) {real, imag} */,
  {32'h45a31dd2, 32'h00000000} /* (19, 0, 12) {real, imag} */,
  {32'h459b12d1, 32'h00000000} /* (19, 0, 11) {real, imag} */,
  {32'h456d3ee2, 32'h00000000} /* (19, 0, 10) {real, imag} */,
  {32'h450e5e3c, 32'h00000000} /* (19, 0, 9) {real, imag} */,
  {32'h43e7edd0, 32'h00000000} /* (19, 0, 8) {real, imag} */,
  {32'hc486ca40, 32'h00000000} /* (19, 0, 7) {real, imag} */,
  {32'hc52157ff, 32'h00000000} /* (19, 0, 6) {real, imag} */,
  {32'hc5b0f790, 32'h00000000} /* (19, 0, 5) {real, imag} */,
  {32'hc5ea1bf1, 32'h00000000} /* (19, 0, 4) {real, imag} */,
  {32'hc6107e36, 32'h00000000} /* (19, 0, 3) {real, imag} */,
  {32'hc613446a, 32'h00000000} /* (19, 0, 2) {real, imag} */,
  {32'hc628fbd2, 32'h00000000} /* (19, 0, 1) {real, imag} */,
  {32'hc6289581, 32'h00000000} /* (19, 0, 0) {real, imag} */,
  {32'hc60c2751, 32'h00000000} /* (18, 31, 31) {real, imag} */,
  {32'hc6167a68, 32'h00000000} /* (18, 31, 30) {real, imag} */,
  {32'hc61f7cb4, 32'h00000000} /* (18, 31, 29) {real, imag} */,
  {32'hc61f2f5d, 32'h00000000} /* (18, 31, 28) {real, imag} */,
  {32'hc6191e47, 32'h00000000} /* (18, 31, 27) {real, imag} */,
  {32'hc6169b04, 32'h00000000} /* (18, 31, 26) {real, imag} */,
  {32'hc613271a, 32'h00000000} /* (18, 31, 25) {real, imag} */,
  {32'hc5f5d806, 32'h00000000} /* (18, 31, 24) {real, imag} */,
  {32'hc5e00ab2, 32'h00000000} /* (18, 31, 23) {real, imag} */,
  {32'hc5b76c3c, 32'h00000000} /* (18, 31, 22) {real, imag} */,
  {32'hc5862302, 32'h00000000} /* (18, 31, 21) {real, imag} */,
  {32'hc522eb5c, 32'h00000000} /* (18, 31, 20) {real, imag} */,
  {32'hc492656c, 32'h00000000} /* (18, 31, 19) {real, imag} */,
  {32'h44673c70, 32'h00000000} /* (18, 31, 18) {real, imag} */,
  {32'h450a9363, 32'h00000000} /* (18, 31, 17) {real, imag} */,
  {32'h45410892, 32'h00000000} /* (18, 31, 16) {real, imag} */,
  {32'h458a0e22, 32'h00000000} /* (18, 31, 15) {real, imag} */,
  {32'h459b0c53, 32'h00000000} /* (18, 31, 14) {real, imag} */,
  {32'h459443e0, 32'h00000000} /* (18, 31, 13) {real, imag} */,
  {32'h457a7918, 32'h00000000} /* (18, 31, 12) {real, imag} */,
  {32'h4558ccf4, 32'h00000000} /* (18, 31, 11) {real, imag} */,
  {32'h44def88c, 32'h00000000} /* (18, 31, 10) {real, imag} */,
  {32'hc3f6e230, 32'h00000000} /* (18, 31, 9) {real, imag} */,
  {32'hc53d90e7, 32'h00000000} /* (18, 31, 8) {real, imag} */,
  {32'hc54d1281, 32'h00000000} /* (18, 31, 7) {real, imag} */,
  {32'hc58b704c, 32'h00000000} /* (18, 31, 6) {real, imag} */,
  {32'hc5cad28a, 32'h00000000} /* (18, 31, 5) {real, imag} */,
  {32'hc5c54940, 32'h00000000} /* (18, 31, 4) {real, imag} */,
  {32'hc6061198, 32'h00000000} /* (18, 31, 3) {real, imag} */,
  {32'hc6067fa7, 32'h00000000} /* (18, 31, 2) {real, imag} */,
  {32'hc6058f1b, 32'h00000000} /* (18, 31, 1) {real, imag} */,
  {32'hc60a5774, 32'h00000000} /* (18, 31, 0) {real, imag} */,
  {32'hc6219870, 32'h00000000} /* (18, 30, 31) {real, imag} */,
  {32'hc627852e, 32'h00000000} /* (18, 30, 30) {real, imag} */,
  {32'hc63be960, 32'h00000000} /* (18, 30, 29) {real, imag} */,
  {32'hc625fdb6, 32'h00000000} /* (18, 30, 28) {real, imag} */,
  {32'hc627fe14, 32'h00000000} /* (18, 30, 27) {real, imag} */,
  {32'hc62c06bf, 32'h00000000} /* (18, 30, 26) {real, imag} */,
  {32'hc60b60cf, 32'h00000000} /* (18, 30, 25) {real, imag} */,
  {32'hc606998c, 32'h00000000} /* (18, 30, 24) {real, imag} */,
  {32'hc5d33f9e, 32'h00000000} /* (18, 30, 23) {real, imag} */,
  {32'hc5c3e882, 32'h00000000} /* (18, 30, 22) {real, imag} */,
  {32'hc58191a2, 32'h00000000} /* (18, 30, 21) {real, imag} */,
  {32'hc4053cb0, 32'h00000000} /* (18, 30, 20) {real, imag} */,
  {32'h449c92cc, 32'h00000000} /* (18, 30, 19) {real, imag} */,
  {32'h4518ffd3, 32'h00000000} /* (18, 30, 18) {real, imag} */,
  {32'h4580f81f, 32'h00000000} /* (18, 30, 17) {real, imag} */,
  {32'h4593d2e2, 32'h00000000} /* (18, 30, 16) {real, imag} */,
  {32'h45be5fe8, 32'h00000000} /* (18, 30, 15) {real, imag} */,
  {32'h45d38223, 32'h00000000} /* (18, 30, 14) {real, imag} */,
  {32'h45c16571, 32'h00000000} /* (18, 30, 13) {real, imag} */,
  {32'h459b1c98, 32'h00000000} /* (18, 30, 12) {real, imag} */,
  {32'h4562aba6, 32'h00000000} /* (18, 30, 11) {real, imag} */,
  {32'h449d0a48, 32'h00000000} /* (18, 30, 10) {real, imag} */,
  {32'hc51f672b, 32'h00000000} /* (18, 30, 9) {real, imag} */,
  {32'hc5877a04, 32'h00000000} /* (18, 30, 8) {real, imag} */,
  {32'hc591d8a6, 32'h00000000} /* (18, 30, 7) {real, imag} */,
  {32'hc5d39e54, 32'h00000000} /* (18, 30, 6) {real, imag} */,
  {32'hc5cc7698, 32'h00000000} /* (18, 30, 5) {real, imag} */,
  {32'hc603f7d2, 32'h00000000} /* (18, 30, 4) {real, imag} */,
  {32'hc6093d80, 32'h00000000} /* (18, 30, 3) {real, imag} */,
  {32'hc6113e76, 32'h00000000} /* (18, 30, 2) {real, imag} */,
  {32'hc610499e, 32'h00000000} /* (18, 30, 1) {real, imag} */,
  {32'hc60ad306, 32'h00000000} /* (18, 30, 0) {real, imag} */,
  {32'hc61bba54, 32'h00000000} /* (18, 29, 31) {real, imag} */,
  {32'hc633afe8, 32'h00000000} /* (18, 29, 30) {real, imag} */,
  {32'hc62b01c3, 32'h00000000} /* (18, 29, 29) {real, imag} */,
  {32'hc6195b10, 32'h00000000} /* (18, 29, 28) {real, imag} */,
  {32'hc61ce3ab, 32'h00000000} /* (18, 29, 27) {real, imag} */,
  {32'hc61c9ff8, 32'h00000000} /* (18, 29, 26) {real, imag} */,
  {32'hc6194f32, 32'h00000000} /* (18, 29, 25) {real, imag} */,
  {32'hc6111b83, 32'h00000000} /* (18, 29, 24) {real, imag} */,
  {32'hc5ea9939, 32'h00000000} /* (18, 29, 23) {real, imag} */,
  {32'hc5a706ae, 32'h00000000} /* (18, 29, 22) {real, imag} */,
  {32'hc55774f0, 32'h00000000} /* (18, 29, 21) {real, imag} */,
  {32'h437d3ce0, 32'h00000000} /* (18, 29, 20) {real, imag} */,
  {32'h4501d3c0, 32'h00000000} /* (18, 29, 19) {real, imag} */,
  {32'h456115d0, 32'h00000000} /* (18, 29, 18) {real, imag} */,
  {32'h45a2fc1e, 32'h00000000} /* (18, 29, 17) {real, imag} */,
  {32'h45d69072, 32'h00000000} /* (18, 29, 16) {real, imag} */,
  {32'h45d4eba8, 32'h00000000} /* (18, 29, 15) {real, imag} */,
  {32'h45bf33dd, 32'h00000000} /* (18, 29, 14) {real, imag} */,
  {32'h45beceea, 32'h00000000} /* (18, 29, 13) {real, imag} */,
  {32'h45985c72, 32'h00000000} /* (18, 29, 12) {real, imag} */,
  {32'h45302c6d, 32'h00000000} /* (18, 29, 11) {real, imag} */,
  {32'h4367bde0, 32'h00000000} /* (18, 29, 10) {real, imag} */,
  {32'hc510a52d, 32'h00000000} /* (18, 29, 9) {real, imag} */,
  {32'hc5a48aef, 32'h00000000} /* (18, 29, 8) {real, imag} */,
  {32'hc5d254f3, 32'h00000000} /* (18, 29, 7) {real, imag} */,
  {32'hc5dcb798, 32'h00000000} /* (18, 29, 6) {real, imag} */,
  {32'hc5f4ae12, 32'h00000000} /* (18, 29, 5) {real, imag} */,
  {32'hc613a702, 32'h00000000} /* (18, 29, 4) {real, imag} */,
  {32'hc6215bc6, 32'h00000000} /* (18, 29, 3) {real, imag} */,
  {32'hc609b486, 32'h00000000} /* (18, 29, 2) {real, imag} */,
  {32'hc614fabc, 32'h00000000} /* (18, 29, 1) {real, imag} */,
  {32'hc61d767b, 32'h00000000} /* (18, 29, 0) {real, imag} */,
  {32'hc6144f3e, 32'h00000000} /* (18, 28, 31) {real, imag} */,
  {32'hc61d244f, 32'h00000000} /* (18, 28, 30) {real, imag} */,
  {32'hc6235656, 32'h00000000} /* (18, 28, 29) {real, imag} */,
  {32'hc6267565, 32'h00000000} /* (18, 28, 28) {real, imag} */,
  {32'hc61a4908, 32'h00000000} /* (18, 28, 27) {real, imag} */,
  {32'hc6160a08, 32'h00000000} /* (18, 28, 26) {real, imag} */,
  {32'hc625f180, 32'h00000000} /* (18, 28, 25) {real, imag} */,
  {32'hc620a79a, 32'h00000000} /* (18, 28, 24) {real, imag} */,
  {32'hc5f76423, 32'h00000000} /* (18, 28, 23) {real, imag} */,
  {32'hc5ac6167, 32'h00000000} /* (18, 28, 22) {real, imag} */,
  {32'hc53a4818, 32'h00000000} /* (18, 28, 21) {real, imag} */,
  {32'h424d8700, 32'h00000000} /* (18, 28, 20) {real, imag} */,
  {32'h45154f94, 32'h00000000} /* (18, 28, 19) {real, imag} */,
  {32'h45965833, 32'h00000000} /* (18, 28, 18) {real, imag} */,
  {32'h45be6ce6, 32'h00000000} /* (18, 28, 17) {real, imag} */,
  {32'h45d65b18, 32'h00000000} /* (18, 28, 16) {real, imag} */,
  {32'h45ddfa07, 32'h00000000} /* (18, 28, 15) {real, imag} */,
  {32'h45d5b0fe, 32'h00000000} /* (18, 28, 14) {real, imag} */,
  {32'h45acd507, 32'h00000000} /* (18, 28, 13) {real, imag} */,
  {32'h459ed852, 32'h00000000} /* (18, 28, 12) {real, imag} */,
  {32'h455bded2, 32'h00000000} /* (18, 28, 11) {real, imag} */,
  {32'hc46b5280, 32'h00000000} /* (18, 28, 10) {real, imag} */,
  {32'hc55e63a7, 32'h00000000} /* (18, 28, 9) {real, imag} */,
  {32'hc59c3644, 32'h00000000} /* (18, 28, 8) {real, imag} */,
  {32'hc5e9fc8f, 32'h00000000} /* (18, 28, 7) {real, imag} */,
  {32'hc6059a37, 32'h00000000} /* (18, 28, 6) {real, imag} */,
  {32'hc60b8c13, 32'h00000000} /* (18, 28, 5) {real, imag} */,
  {32'hc60ffb07, 32'h00000000} /* (18, 28, 4) {real, imag} */,
  {32'hc61a5972, 32'h00000000} /* (18, 28, 3) {real, imag} */,
  {32'hc61ce746, 32'h00000000} /* (18, 28, 2) {real, imag} */,
  {32'hc61d6469, 32'h00000000} /* (18, 28, 1) {real, imag} */,
  {32'hc61e96dc, 32'h00000000} /* (18, 28, 0) {real, imag} */,
  {32'hc614ca8f, 32'h00000000} /* (18, 27, 31) {real, imag} */,
  {32'hc6182230, 32'h00000000} /* (18, 27, 30) {real, imag} */,
  {32'hc61431f0, 32'h00000000} /* (18, 27, 29) {real, imag} */,
  {32'hc61814c5, 32'h00000000} /* (18, 27, 28) {real, imag} */,
  {32'hc6121c70, 32'h00000000} /* (18, 27, 27) {real, imag} */,
  {32'hc6237397, 32'h00000000} /* (18, 27, 26) {real, imag} */,
  {32'hc62091cc, 32'h00000000} /* (18, 27, 25) {real, imag} */,
  {32'hc608d922, 32'h00000000} /* (18, 27, 24) {real, imag} */,
  {32'hc5ddf1a6, 32'h00000000} /* (18, 27, 23) {real, imag} */,
  {32'hc59f56bc, 32'h00000000} /* (18, 27, 22) {real, imag} */,
  {32'hc5217bd6, 32'h00000000} /* (18, 27, 21) {real, imag} */,
  {32'h43cf2320, 32'h00000000} /* (18, 27, 20) {real, imag} */,
  {32'h45327d04, 32'h00000000} /* (18, 27, 19) {real, imag} */,
  {32'h4591f69a, 32'h00000000} /* (18, 27, 18) {real, imag} */,
  {32'h45bdd624, 32'h00000000} /* (18, 27, 17) {real, imag} */,
  {32'h45cd9476, 32'h00000000} /* (18, 27, 16) {real, imag} */,
  {32'h45ce3a94, 32'h00000000} /* (18, 27, 15) {real, imag} */,
  {32'h45f2804f, 32'h00000000} /* (18, 27, 14) {real, imag} */,
  {32'h45c24348, 32'h00000000} /* (18, 27, 13) {real, imag} */,
  {32'h4585b00e, 32'h00000000} /* (18, 27, 12) {real, imag} */,
  {32'h450dcec8, 32'h00000000} /* (18, 27, 11) {real, imag} */,
  {32'hc4c55ef8, 32'h00000000} /* (18, 27, 10) {real, imag} */,
  {32'hc588a2d4, 32'h00000000} /* (18, 27, 9) {real, imag} */,
  {32'hc5bc075f, 32'h00000000} /* (18, 27, 8) {real, imag} */,
  {32'hc5eb8d66, 32'h00000000} /* (18, 27, 7) {real, imag} */,
  {32'hc605a4ea, 32'h00000000} /* (18, 27, 6) {real, imag} */,
  {32'hc61bcc90, 32'h00000000} /* (18, 27, 5) {real, imag} */,
  {32'hc624faff, 32'h00000000} /* (18, 27, 4) {real, imag} */,
  {32'hc6182227, 32'h00000000} /* (18, 27, 3) {real, imag} */,
  {32'hc616b781, 32'h00000000} /* (18, 27, 2) {real, imag} */,
  {32'hc626359a, 32'h00000000} /* (18, 27, 1) {real, imag} */,
  {32'hc613b39b, 32'h00000000} /* (18, 27, 0) {real, imag} */,
  {32'hc6102642, 32'h00000000} /* (18, 26, 31) {real, imag} */,
  {32'hc61470c6, 32'h00000000} /* (18, 26, 30) {real, imag} */,
  {32'hc60c625c, 32'h00000000} /* (18, 26, 29) {real, imag} */,
  {32'hc60ada22, 32'h00000000} /* (18, 26, 28) {real, imag} */,
  {32'hc6081f32, 32'h00000000} /* (18, 26, 27) {real, imag} */,
  {32'hc6154d5a, 32'h00000000} /* (18, 26, 26) {real, imag} */,
  {32'hc618cd14, 32'h00000000} /* (18, 26, 25) {real, imag} */,
  {32'hc6041f47, 32'h00000000} /* (18, 26, 24) {real, imag} */,
  {32'hc5d33f94, 32'h00000000} /* (18, 26, 23) {real, imag} */,
  {32'hc59fe601, 32'h00000000} /* (18, 26, 22) {real, imag} */,
  {32'hc51f45ed, 32'h00000000} /* (18, 26, 21) {real, imag} */,
  {32'h439cb530, 32'h00000000} /* (18, 26, 20) {real, imag} */,
  {32'h452ff2b6, 32'h00000000} /* (18, 26, 19) {real, imag} */,
  {32'h458892cd, 32'h00000000} /* (18, 26, 18) {real, imag} */,
  {32'h45994d42, 32'h00000000} /* (18, 26, 17) {real, imag} */,
  {32'h45db3122, 32'h00000000} /* (18, 26, 16) {real, imag} */,
  {32'h45c0883a, 32'h00000000} /* (18, 26, 15) {real, imag} */,
  {32'h45d68f37, 32'h00000000} /* (18, 26, 14) {real, imag} */,
  {32'h45b71ff7, 32'h00000000} /* (18, 26, 13) {real, imag} */,
  {32'h458537c3, 32'h00000000} /* (18, 26, 12) {real, imag} */,
  {32'h44e562ac, 32'h00000000} /* (18, 26, 11) {real, imag} */,
  {32'hc4fa83a4, 32'h00000000} /* (18, 26, 10) {real, imag} */,
  {32'hc57e798a, 32'h00000000} /* (18, 26, 9) {real, imag} */,
  {32'hc5d5612e, 32'h00000000} /* (18, 26, 8) {real, imag} */,
  {32'hc5eebd4c, 32'h00000000} /* (18, 26, 7) {real, imag} */,
  {32'hc5fa6263, 32'h00000000} /* (18, 26, 6) {real, imag} */,
  {32'hc61912f7, 32'h00000000} /* (18, 26, 5) {real, imag} */,
  {32'hc61a41b6, 32'h00000000} /* (18, 26, 4) {real, imag} */,
  {32'hc619ecb0, 32'h00000000} /* (18, 26, 3) {real, imag} */,
  {32'hc6228694, 32'h00000000} /* (18, 26, 2) {real, imag} */,
  {32'hc6259118, 32'h00000000} /* (18, 26, 1) {real, imag} */,
  {32'hc611b41a, 32'h00000000} /* (18, 26, 0) {real, imag} */,
  {32'hc6036f98, 32'h00000000} /* (18, 25, 31) {real, imag} */,
  {32'hc5ff1196, 32'h00000000} /* (18, 25, 30) {real, imag} */,
  {32'hc60490cb, 32'h00000000} /* (18, 25, 29) {real, imag} */,
  {32'hc6025b37, 32'h00000000} /* (18, 25, 28) {real, imag} */,
  {32'hc61afe56, 32'h00000000} /* (18, 25, 27) {real, imag} */,
  {32'hc61d9047, 32'h00000000} /* (18, 25, 26) {real, imag} */,
  {32'hc5f8e102, 32'h00000000} /* (18, 25, 25) {real, imag} */,
  {32'hc5e4fe13, 32'h00000000} /* (18, 25, 24) {real, imag} */,
  {32'hc5d1bb9d, 32'h00000000} /* (18, 25, 23) {real, imag} */,
  {32'hc57c1e8e, 32'h00000000} /* (18, 25, 22) {real, imag} */,
  {32'hc548d7bf, 32'h00000000} /* (18, 25, 21) {real, imag} */,
  {32'h450ce116, 32'h00000000} /* (18, 25, 20) {real, imag} */,
  {32'h45ac6f3a, 32'h00000000} /* (18, 25, 19) {real, imag} */,
  {32'h45713be5, 32'h00000000} /* (18, 25, 18) {real, imag} */,
  {32'h458f504a, 32'h00000000} /* (18, 25, 17) {real, imag} */,
  {32'h45ae3412, 32'h00000000} /* (18, 25, 16) {real, imag} */,
  {32'h45b1ca67, 32'h00000000} /* (18, 25, 15) {real, imag} */,
  {32'h45b564aa, 32'h00000000} /* (18, 25, 14) {real, imag} */,
  {32'h45919596, 32'h00000000} /* (18, 25, 13) {real, imag} */,
  {32'h459b2478, 32'h00000000} /* (18, 25, 12) {real, imag} */,
  {32'h44c07430, 32'h00000000} /* (18, 25, 11) {real, imag} */,
  {32'hc5124cfd, 32'h00000000} /* (18, 25, 10) {real, imag} */,
  {32'hc58ea3fa, 32'h00000000} /* (18, 25, 9) {real, imag} */,
  {32'hc5da8ae1, 32'h00000000} /* (18, 25, 8) {real, imag} */,
  {32'hc5f13b39, 32'h00000000} /* (18, 25, 7) {real, imag} */,
  {32'hc5e3e37d, 32'h00000000} /* (18, 25, 6) {real, imag} */,
  {32'hc5f3f720, 32'h00000000} /* (18, 25, 5) {real, imag} */,
  {32'hc60561d2, 32'h00000000} /* (18, 25, 4) {real, imag} */,
  {32'hc60d214e, 32'h00000000} /* (18, 25, 3) {real, imag} */,
  {32'hc6139246, 32'h00000000} /* (18, 25, 2) {real, imag} */,
  {32'hc61a9d75, 32'h00000000} /* (18, 25, 1) {real, imag} */,
  {32'hc604b39d, 32'h00000000} /* (18, 25, 0) {real, imag} */,
  {32'hc5e8d14e, 32'h00000000} /* (18, 24, 31) {real, imag} */,
  {32'hc5dd2894, 32'h00000000} /* (18, 24, 30) {real, imag} */,
  {32'hc5e733e2, 32'h00000000} /* (18, 24, 29) {real, imag} */,
  {32'hc5fe8b14, 32'h00000000} /* (18, 24, 28) {real, imag} */,
  {32'hc5f502b8, 32'h00000000} /* (18, 24, 27) {real, imag} */,
  {32'hc601f851, 32'h00000000} /* (18, 24, 26) {real, imag} */,
  {32'hc5e1cb3f, 32'h00000000} /* (18, 24, 25) {real, imag} */,
  {32'hc5d7df3e, 32'h00000000} /* (18, 24, 24) {real, imag} */,
  {32'hc5b12a6e, 32'h00000000} /* (18, 24, 23) {real, imag} */,
  {32'hc593604b, 32'h00000000} /* (18, 24, 22) {real, imag} */,
  {32'hc4fbfa00, 32'h00000000} /* (18, 24, 21) {real, imag} */,
  {32'h4512ea22, 32'h00000000} /* (18, 24, 20) {real, imag} */,
  {32'h458bd012, 32'h00000000} /* (18, 24, 19) {real, imag} */,
  {32'h45709b86, 32'h00000000} /* (18, 24, 18) {real, imag} */,
  {32'h45929512, 32'h00000000} /* (18, 24, 17) {real, imag} */,
  {32'h4594b784, 32'h00000000} /* (18, 24, 16) {real, imag} */,
  {32'h4595615c, 32'h00000000} /* (18, 24, 15) {real, imag} */,
  {32'h45919432, 32'h00000000} /* (18, 24, 14) {real, imag} */,
  {32'h458dfbba, 32'h00000000} /* (18, 24, 13) {real, imag} */,
  {32'h45194e48, 32'h00000000} /* (18, 24, 12) {real, imag} */,
  {32'h44776ddc, 32'h00000000} /* (18, 24, 11) {real, imag} */,
  {32'hc5268a40, 32'h00000000} /* (18, 24, 10) {real, imag} */,
  {32'hc592786d, 32'h00000000} /* (18, 24, 9) {real, imag} */,
  {32'hc5b66c40, 32'h00000000} /* (18, 24, 8) {real, imag} */,
  {32'hc5e0d37a, 32'h00000000} /* (18, 24, 7) {real, imag} */,
  {32'hc5d6e4cd, 32'h00000000} /* (18, 24, 6) {real, imag} */,
  {32'hc5d0856c, 32'h00000000} /* (18, 24, 5) {real, imag} */,
  {32'hc5f6bbd1, 32'h00000000} /* (18, 24, 4) {real, imag} */,
  {32'hc5fd41c0, 32'h00000000} /* (18, 24, 3) {real, imag} */,
  {32'hc6024036, 32'h00000000} /* (18, 24, 2) {real, imag} */,
  {32'hc604d97f, 32'h00000000} /* (18, 24, 1) {real, imag} */,
  {32'hc5e37a42, 32'h00000000} /* (18, 24, 0) {real, imag} */,
  {32'hc5ad28a8, 32'h00000000} /* (18, 23, 31) {real, imag} */,
  {32'hc5b41d59, 32'h00000000} /* (18, 23, 30) {real, imag} */,
  {32'hc5c03deb, 32'h00000000} /* (18, 23, 29) {real, imag} */,
  {32'hc5db012e, 32'h00000000} /* (18, 23, 28) {real, imag} */,
  {32'hc5c4a3f5, 32'h00000000} /* (18, 23, 27) {real, imag} */,
  {32'hc5b9fc61, 32'h00000000} /* (18, 23, 26) {real, imag} */,
  {32'hc5b9a434, 32'h00000000} /* (18, 23, 25) {real, imag} */,
  {32'hc5c63c08, 32'h00000000} /* (18, 23, 24) {real, imag} */,
  {32'hc596b0ae, 32'h00000000} /* (18, 23, 23) {real, imag} */,
  {32'hc58438bf, 32'h00000000} /* (18, 23, 22) {real, imag} */,
  {32'hc4c19754, 32'h00000000} /* (18, 23, 21) {real, imag} */,
  {32'h44e49a70, 32'h00000000} /* (18, 23, 20) {real, imag} */,
  {32'h452ecc00, 32'h00000000} /* (18, 23, 19) {real, imag} */,
  {32'h454b13ba, 32'h00000000} /* (18, 23, 18) {real, imag} */,
  {32'h4598da74, 32'h00000000} /* (18, 23, 17) {real, imag} */,
  {32'h459bd8d5, 32'h00000000} /* (18, 23, 16) {real, imag} */,
  {32'h458bb8fe, 32'h00000000} /* (18, 23, 15) {real, imag} */,
  {32'h456f175a, 32'h00000000} /* (18, 23, 14) {real, imag} */,
  {32'h45554692, 32'h00000000} /* (18, 23, 13) {real, imag} */,
  {32'h452f467c, 32'h00000000} /* (18, 23, 12) {real, imag} */,
  {32'h43a7e9d0, 32'h00000000} /* (18, 23, 11) {real, imag} */,
  {32'hc52504b2, 32'h00000000} /* (18, 23, 10) {real, imag} */,
  {32'hc576faa9, 32'h00000000} /* (18, 23, 9) {real, imag} */,
  {32'hc595cb80, 32'h00000000} /* (18, 23, 8) {real, imag} */,
  {32'hc5b03922, 32'h00000000} /* (18, 23, 7) {real, imag} */,
  {32'hc5ac2b7b, 32'h00000000} /* (18, 23, 6) {real, imag} */,
  {32'hc5ad8c03, 32'h00000000} /* (18, 23, 5) {real, imag} */,
  {32'hc5ce90d2, 32'h00000000} /* (18, 23, 4) {real, imag} */,
  {32'hc5da9b9c, 32'h00000000} /* (18, 23, 3) {real, imag} */,
  {32'hc5f01939, 32'h00000000} /* (18, 23, 2) {real, imag} */,
  {32'hc5ce98f2, 32'h00000000} /* (18, 23, 1) {real, imag} */,
  {32'hc5b6bb5b, 32'h00000000} /* (18, 23, 0) {real, imag} */,
  {32'hc583244e, 32'h00000000} /* (18, 22, 31) {real, imag} */,
  {32'hc582dc0d, 32'h00000000} /* (18, 22, 30) {real, imag} */,
  {32'hc59234cc, 32'h00000000} /* (18, 22, 29) {real, imag} */,
  {32'hc5ba0721, 32'h00000000} /* (18, 22, 28) {real, imag} */,
  {32'hc5af7056, 32'h00000000} /* (18, 22, 27) {real, imag} */,
  {32'hc58f449a, 32'h00000000} /* (18, 22, 26) {real, imag} */,
  {32'hc54c5208, 32'h00000000} /* (18, 22, 25) {real, imag} */,
  {32'hc573d530, 32'h00000000} /* (18, 22, 24) {real, imag} */,
  {32'hc58a62fe, 32'h00000000} /* (18, 22, 23) {real, imag} */,
  {32'hc53fe034, 32'h00000000} /* (18, 22, 22) {real, imag} */,
  {32'hc4a06709, 32'h00000000} /* (18, 22, 21) {real, imag} */,
  {32'h43b49a90, 32'h00000000} /* (18, 22, 20) {real, imag} */,
  {32'h44dd3656, 32'h00000000} /* (18, 22, 19) {real, imag} */,
  {32'h4530c54a, 32'h00000000} /* (18, 22, 18) {real, imag} */,
  {32'h457caa24, 32'h00000000} /* (18, 22, 17) {real, imag} */,
  {32'h4579b04c, 32'h00000000} /* (18, 22, 16) {real, imag} */,
  {32'h45514c5a, 32'h00000000} /* (18, 22, 15) {real, imag} */,
  {32'h453d034e, 32'h00000000} /* (18, 22, 14) {real, imag} */,
  {32'h44f04a1e, 32'h00000000} /* (18, 22, 13) {real, imag} */,
  {32'h44e24c38, 32'h00000000} /* (18, 22, 12) {real, imag} */,
  {32'hc404853c, 32'h00000000} /* (18, 22, 11) {real, imag} */,
  {32'hc4f7012a, 32'h00000000} /* (18, 22, 10) {real, imag} */,
  {32'hc5377426, 32'h00000000} /* (18, 22, 9) {real, imag} */,
  {32'hc57f5920, 32'h00000000} /* (18, 22, 8) {real, imag} */,
  {32'hc5864a6a, 32'h00000000} /* (18, 22, 7) {real, imag} */,
  {32'hc57f0cec, 32'h00000000} /* (18, 22, 6) {real, imag} */,
  {32'hc58935b9, 32'h00000000} /* (18, 22, 5) {real, imag} */,
  {32'hc57e4f58, 32'h00000000} /* (18, 22, 4) {real, imag} */,
  {32'hc58e6690, 32'h00000000} /* (18, 22, 3) {real, imag} */,
  {32'hc58ddaa7, 32'h00000000} /* (18, 22, 2) {real, imag} */,
  {32'hc5a000a4, 32'h00000000} /* (18, 22, 1) {real, imag} */,
  {32'hc58f5964, 32'h00000000} /* (18, 22, 0) {real, imag} */,
  {32'hc50bd76d, 32'h00000000} /* (18, 21, 31) {real, imag} */,
  {32'hc54d7539, 32'h00000000} /* (18, 21, 30) {real, imag} */,
  {32'hc51d5da7, 32'h00000000} /* (18, 21, 29) {real, imag} */,
  {32'hc50db540, 32'h00000000} /* (18, 21, 28) {real, imag} */,
  {32'hc53fbcb1, 32'h00000000} /* (18, 21, 27) {real, imag} */,
  {32'hc52bd242, 32'h00000000} /* (18, 21, 26) {real, imag} */,
  {32'hc4fb2793, 32'h00000000} /* (18, 21, 25) {real, imag} */,
  {32'hc4c1c517, 32'h00000000} /* (18, 21, 24) {real, imag} */,
  {32'hc4cb60de, 32'h00000000} /* (18, 21, 23) {real, imag} */,
  {32'hc4bda8ec, 32'h00000000} /* (18, 21, 22) {real, imag} */,
  {32'hc4cbe1d5, 32'h00000000} /* (18, 21, 21) {real, imag} */,
  {32'hc32b0c5c, 32'h00000000} /* (18, 21, 20) {real, imag} */,
  {32'h4484862a, 32'h00000000} /* (18, 21, 19) {real, imag} */,
  {32'h447ed731, 32'h00000000} /* (18, 21, 18) {real, imag} */,
  {32'h4467dae8, 32'h00000000} /* (18, 21, 17) {real, imag} */,
  {32'h4473889a, 32'h00000000} /* (18, 21, 16) {real, imag} */,
  {32'h443b2548, 32'h00000000} /* (18, 21, 15) {real, imag} */,
  {32'h43f0ab40, 32'h00000000} /* (18, 21, 14) {real, imag} */,
  {32'h43ec7558, 32'h00000000} /* (18, 21, 13) {real, imag} */,
  {32'hc2ef5b50, 32'h00000000} /* (18, 21, 12) {real, imag} */,
  {32'hc39fd1b8, 32'h00000000} /* (18, 21, 11) {real, imag} */,
  {32'hc48afb40, 32'h00000000} /* (18, 21, 10) {real, imag} */,
  {32'hc4d3943b, 32'h00000000} /* (18, 21, 9) {real, imag} */,
  {32'hc4d211a9, 32'h00000000} /* (18, 21, 8) {real, imag} */,
  {32'hc4eefa84, 32'h00000000} /* (18, 21, 7) {real, imag} */,
  {32'hc4a5f8ea, 32'h00000000} /* (18, 21, 6) {real, imag} */,
  {32'hc4aecf33, 32'h00000000} /* (18, 21, 5) {real, imag} */,
  {32'hc4e77ed6, 32'h00000000} /* (18, 21, 4) {real, imag} */,
  {32'hc4a50900, 32'h00000000} /* (18, 21, 3) {real, imag} */,
  {32'hc500f697, 32'h00000000} /* (18, 21, 2) {real, imag} */,
  {32'hc523614b, 32'h00000000} /* (18, 21, 1) {real, imag} */,
  {32'hc4d5c0b7, 32'h00000000} /* (18, 21, 0) {real, imag} */,
  {32'h4473c082, 32'h00000000} /* (18, 20, 31) {real, imag} */,
  {32'h440b9487, 32'h00000000} /* (18, 20, 30) {real, imag} */,
  {32'h438d5fee, 32'h00000000} /* (18, 20, 29) {real, imag} */,
  {32'h4467090e, 32'h00000000} /* (18, 20, 28) {real, imag} */,
  {32'h446cdca2, 32'h00000000} /* (18, 20, 27) {real, imag} */,
  {32'h4413ae9c, 32'h00000000} /* (18, 20, 26) {real, imag} */,
  {32'h444b60fd, 32'h00000000} /* (18, 20, 25) {real, imag} */,
  {32'h4494860e, 32'h00000000} /* (18, 20, 24) {real, imag} */,
  {32'h44ff1d8f, 32'h00000000} /* (18, 20, 23) {real, imag} */,
  {32'h44491dc3, 32'h00000000} /* (18, 20, 22) {real, imag} */,
  {32'hc45e9321, 32'h00000000} /* (18, 20, 21) {real, imag} */,
  {32'hc4a60758, 32'h00000000} /* (18, 20, 20) {real, imag} */,
  {32'hc44e1640, 32'h00000000} /* (18, 20, 19) {real, imag} */,
  {32'hc4ca328a, 32'h00000000} /* (18, 20, 18) {real, imag} */,
  {32'hc4bbe548, 32'h00000000} /* (18, 20, 17) {real, imag} */,
  {32'hc516cabd, 32'h00000000} /* (18, 20, 16) {real, imag} */,
  {32'hc4f3eaa3, 32'h00000000} /* (18, 20, 15) {real, imag} */,
  {32'hc516c820, 32'h00000000} /* (18, 20, 14) {real, imag} */,
  {32'hc5082ad9, 32'h00000000} /* (18, 20, 13) {real, imag} */,
  {32'hc50c8be8, 32'h00000000} /* (18, 20, 12) {real, imag} */,
  {32'hc515faec, 32'h00000000} /* (18, 20, 11) {real, imag} */,
  {32'hc35f6462, 32'h00000000} /* (18, 20, 10) {real, imag} */,
  {32'h440ccc09, 32'h00000000} /* (18, 20, 9) {real, imag} */,
  {32'h44fbd066, 32'h00000000} /* (18, 20, 8) {real, imag} */,
  {32'h44fc3a7b, 32'h00000000} /* (18, 20, 7) {real, imag} */,
  {32'h4440185b, 32'h00000000} /* (18, 20, 6) {real, imag} */,
  {32'h449fe452, 32'h00000000} /* (18, 20, 5) {real, imag} */,
  {32'h44f421fa, 32'h00000000} /* (18, 20, 4) {real, imag} */,
  {32'h44ffa41a, 32'h00000000} /* (18, 20, 3) {real, imag} */,
  {32'h45043871, 32'h00000000} /* (18, 20, 2) {real, imag} */,
  {32'h44b1d324, 32'h00000000} /* (18, 20, 1) {real, imag} */,
  {32'h44c2dbea, 32'h00000000} /* (18, 20, 0) {real, imag} */,
  {32'h45573822, 32'h00000000} /* (18, 19, 31) {real, imag} */,
  {32'h45627462, 32'h00000000} /* (18, 19, 30) {real, imag} */,
  {32'h45531419, 32'h00000000} /* (18, 19, 29) {real, imag} */,
  {32'h45630eb7, 32'h00000000} /* (18, 19, 28) {real, imag} */,
  {32'h45469ac2, 32'h00000000} /* (18, 19, 27) {real, imag} */,
  {32'h454983a8, 32'h00000000} /* (18, 19, 26) {real, imag} */,
  {32'h455b4f9d, 32'h00000000} /* (18, 19, 25) {real, imag} */,
  {32'h458eba0c, 32'h00000000} /* (18, 19, 24) {real, imag} */,
  {32'h45366f33, 32'h00000000} /* (18, 19, 23) {real, imag} */,
  {32'h45031ded, 32'h00000000} /* (18, 19, 22) {real, imag} */,
  {32'h438d6b80, 32'h00000000} /* (18, 19, 21) {real, imag} */,
  {32'hc5338a69, 32'h00000000} /* (18, 19, 20) {real, imag} */,
  {32'hc524e79a, 32'h00000000} /* (18, 19, 19) {real, imag} */,
  {32'hc53247e8, 32'h00000000} /* (18, 19, 18) {real, imag} */,
  {32'hc581fa0f, 32'h00000000} /* (18, 19, 17) {real, imag} */,
  {32'hc55bdcc6, 32'h00000000} /* (18, 19, 16) {real, imag} */,
  {32'hc56e6344, 32'h00000000} /* (18, 19, 15) {real, imag} */,
  {32'hc5654a86, 32'h00000000} /* (18, 19, 14) {real, imag} */,
  {32'hc55908b5, 32'h00000000} /* (18, 19, 13) {real, imag} */,
  {32'hc5361879, 32'h00000000} /* (18, 19, 12) {real, imag} */,
  {32'hc521b88a, 32'h00000000} /* (18, 19, 11) {real, imag} */,
  {32'hc3c827f4, 32'h00000000} /* (18, 19, 10) {real, imag} */,
  {32'h451ce38f, 32'h00000000} /* (18, 19, 9) {real, imag} */,
  {32'h456f178b, 32'h00000000} /* (18, 19, 8) {real, imag} */,
  {32'h4587a92e, 32'h00000000} /* (18, 19, 7) {real, imag} */,
  {32'h45576111, 32'h00000000} /* (18, 19, 6) {real, imag} */,
  {32'h455c2370, 32'h00000000} /* (18, 19, 5) {real, imag} */,
  {32'h45814fe6, 32'h00000000} /* (18, 19, 4) {real, imag} */,
  {32'h45699270, 32'h00000000} /* (18, 19, 3) {real, imag} */,
  {32'h459b037c, 32'h00000000} /* (18, 19, 2) {real, imag} */,
  {32'h45958f65, 32'h00000000} /* (18, 19, 1) {real, imag} */,
  {32'h455045f2, 32'h00000000} /* (18, 19, 0) {real, imag} */,
  {32'h45b2df28, 32'h00000000} /* (18, 18, 31) {real, imag} */,
  {32'h45cf8cab, 32'h00000000} /* (18, 18, 30) {real, imag} */,
  {32'h45aacf16, 32'h00000000} /* (18, 18, 29) {real, imag} */,
  {32'h45a6dae0, 32'h00000000} /* (18, 18, 28) {real, imag} */,
  {32'h459ebd44, 32'h00000000} /* (18, 18, 27) {real, imag} */,
  {32'h45972984, 32'h00000000} /* (18, 18, 26) {real, imag} */,
  {32'h45a7a710, 32'h00000000} /* (18, 18, 25) {real, imag} */,
  {32'h459ea03b, 32'h00000000} /* (18, 18, 24) {real, imag} */,
  {32'h4582c1d6, 32'h00000000} /* (18, 18, 23) {real, imag} */,
  {32'h4528c88a, 32'h00000000} /* (18, 18, 22) {real, imag} */,
  {32'h439d3118, 32'h00000000} /* (18, 18, 21) {real, imag} */,
  {32'hc50516c6, 32'h00000000} /* (18, 18, 20) {real, imag} */,
  {32'hc55db0a8, 32'h00000000} /* (18, 18, 19) {real, imag} */,
  {32'hc592d6dc, 32'h00000000} /* (18, 18, 18) {real, imag} */,
  {32'hc5a32f44, 32'h00000000} /* (18, 18, 17) {real, imag} */,
  {32'hc5a3b31f, 32'h00000000} /* (18, 18, 16) {real, imag} */,
  {32'hc5a2ceca, 32'h00000000} /* (18, 18, 15) {real, imag} */,
  {32'hc59a0d01, 32'h00000000} /* (18, 18, 14) {real, imag} */,
  {32'hc598b746, 32'h00000000} /* (18, 18, 13) {real, imag} */,
  {32'hc5839126, 32'h00000000} /* (18, 18, 12) {real, imag} */,
  {32'hc501b338, 32'h00000000} /* (18, 18, 11) {real, imag} */,
  {32'h42da9720, 32'h00000000} /* (18, 18, 10) {real, imag} */,
  {32'h455a4ee9, 32'h00000000} /* (18, 18, 9) {real, imag} */,
  {32'h459c1b91, 32'h00000000} /* (18, 18, 8) {real, imag} */,
  {32'h45a1d2fe, 32'h00000000} /* (18, 18, 7) {real, imag} */,
  {32'h458de685, 32'h00000000} /* (18, 18, 6) {real, imag} */,
  {32'h45904ed6, 32'h00000000} /* (18, 18, 5) {real, imag} */,
  {32'h459e7e04, 32'h00000000} /* (18, 18, 4) {real, imag} */,
  {32'h459d9cde, 32'h00000000} /* (18, 18, 3) {real, imag} */,
  {32'h45a0308a, 32'h00000000} /* (18, 18, 2) {real, imag} */,
  {32'h45c4a53a, 32'h00000000} /* (18, 18, 1) {real, imag} */,
  {32'h45a3de4f, 32'h00000000} /* (18, 18, 0) {real, imag} */,
  {32'h45c96742, 32'h00000000} /* (18, 17, 31) {real, imag} */,
  {32'h45d8deed, 32'h00000000} /* (18, 17, 30) {real, imag} */,
  {32'h45c84c8b, 32'h00000000} /* (18, 17, 29) {real, imag} */,
  {32'h45d3826b, 32'h00000000} /* (18, 17, 28) {real, imag} */,
  {32'h45cf4c64, 32'h00000000} /* (18, 17, 27) {real, imag} */,
  {32'h45b12fed, 32'h00000000} /* (18, 17, 26) {real, imag} */,
  {32'h45b00ba0, 32'h00000000} /* (18, 17, 25) {real, imag} */,
  {32'h45a0645a, 32'h00000000} /* (18, 17, 24) {real, imag} */,
  {32'h45a28f6f, 32'h00000000} /* (18, 17, 23) {real, imag} */,
  {32'h452f428a, 32'h00000000} /* (18, 17, 22) {real, imag} */,
  {32'h43ff4570, 32'h00000000} /* (18, 17, 21) {real, imag} */,
  {32'hc52407fa, 32'h00000000} /* (18, 17, 20) {real, imag} */,
  {32'hc585579a, 32'h00000000} /* (18, 17, 19) {real, imag} */,
  {32'hc5930ec5, 32'h00000000} /* (18, 17, 18) {real, imag} */,
  {32'hc5b97e98, 32'h00000000} /* (18, 17, 17) {real, imag} */,
  {32'hc5b978b7, 32'h00000000} /* (18, 17, 16) {real, imag} */,
  {32'hc5bded84, 32'h00000000} /* (18, 17, 15) {real, imag} */,
  {32'hc5b6fcbf, 32'h00000000} /* (18, 17, 14) {real, imag} */,
  {32'hc59a4ac1, 32'h00000000} /* (18, 17, 13) {real, imag} */,
  {32'hc59f326b, 32'h00000000} /* (18, 17, 12) {real, imag} */,
  {32'hc50cbb80, 32'h00000000} /* (18, 17, 11) {real, imag} */,
  {32'h44bcbfbc, 32'h00000000} /* (18, 17, 10) {real, imag} */,
  {32'h458902c0, 32'h00000000} /* (18, 17, 9) {real, imag} */,
  {32'h4599dc12, 32'h00000000} /* (18, 17, 8) {real, imag} */,
  {32'h45a3eab1, 32'h00000000} /* (18, 17, 7) {real, imag} */,
  {32'h45b984ad, 32'h00000000} /* (18, 17, 6) {real, imag} */,
  {32'h45a857fd, 32'h00000000} /* (18, 17, 5) {real, imag} */,
  {32'h45b7fce9, 32'h00000000} /* (18, 17, 4) {real, imag} */,
  {32'h45caffea, 32'h00000000} /* (18, 17, 3) {real, imag} */,
  {32'h45d411e5, 32'h00000000} /* (18, 17, 2) {real, imag} */,
  {32'h45c14a74, 32'h00000000} /* (18, 17, 1) {real, imag} */,
  {32'h45d28bf3, 32'h00000000} /* (18, 17, 0) {real, imag} */,
  {32'h45c029f9, 32'h00000000} /* (18, 16, 31) {real, imag} */,
  {32'h45e693d5, 32'h00000000} /* (18, 16, 30) {real, imag} */,
  {32'h45f9d5c9, 32'h00000000} /* (18, 16, 29) {real, imag} */,
  {32'h45d6ef76, 32'h00000000} /* (18, 16, 28) {real, imag} */,
  {32'h45f13c77, 32'h00000000} /* (18, 16, 27) {real, imag} */,
  {32'h45e3fed8, 32'h00000000} /* (18, 16, 26) {real, imag} */,
  {32'h45c0533d, 32'h00000000} /* (18, 16, 25) {real, imag} */,
  {32'h45cbdd90, 32'h00000000} /* (18, 16, 24) {real, imag} */,
  {32'h45a9d106, 32'h00000000} /* (18, 16, 23) {real, imag} */,
  {32'h45451dd2, 32'h00000000} /* (18, 16, 22) {real, imag} */,
  {32'h449b1918, 32'h00000000} /* (18, 16, 21) {real, imag} */,
  {32'hc5603e4e, 32'h00000000} /* (18, 16, 20) {real, imag} */,
  {32'hc5931802, 32'h00000000} /* (18, 16, 19) {real, imag} */,
  {32'hc5aef3fa, 32'h00000000} /* (18, 16, 18) {real, imag} */,
  {32'hc5becdec, 32'h00000000} /* (18, 16, 17) {real, imag} */,
  {32'hc5d04fcc, 32'h00000000} /* (18, 16, 16) {real, imag} */,
  {32'hc5d5b851, 32'h00000000} /* (18, 16, 15) {real, imag} */,
  {32'hc5c6ca11, 32'h00000000} /* (18, 16, 14) {real, imag} */,
  {32'hc5a249b5, 32'h00000000} /* (18, 16, 13) {real, imag} */,
  {32'hc59397e2, 32'h00000000} /* (18, 16, 12) {real, imag} */,
  {32'hc48ab974, 32'h00000000} /* (18, 16, 11) {real, imag} */,
  {32'h4508f349, 32'h00000000} /* (18, 16, 10) {real, imag} */,
  {32'h45965267, 32'h00000000} /* (18, 16, 9) {real, imag} */,
  {32'h45cb9c4c, 32'h00000000} /* (18, 16, 8) {real, imag} */,
  {32'h45b96a7c, 32'h00000000} /* (18, 16, 7) {real, imag} */,
  {32'h45b5e9eb, 32'h00000000} /* (18, 16, 6) {real, imag} */,
  {32'h45c6c3aa, 32'h00000000} /* (18, 16, 5) {real, imag} */,
  {32'h45c5db33, 32'h00000000} /* (18, 16, 4) {real, imag} */,
  {32'h45d80042, 32'h00000000} /* (18, 16, 3) {real, imag} */,
  {32'h45dd3336, 32'h00000000} /* (18, 16, 2) {real, imag} */,
  {32'h45eaf3d6, 32'h00000000} /* (18, 16, 1) {real, imag} */,
  {32'h45c0fd88, 32'h00000000} /* (18, 16, 0) {real, imag} */,
  {32'h45b05dba, 32'h00000000} /* (18, 15, 31) {real, imag} */,
  {32'h45cf0a5a, 32'h00000000} /* (18, 15, 30) {real, imag} */,
  {32'h45df4104, 32'h00000000} /* (18, 15, 29) {real, imag} */,
  {32'h45d858c4, 32'h00000000} /* (18, 15, 28) {real, imag} */,
  {32'h45e8f1c0, 32'h00000000} /* (18, 15, 27) {real, imag} */,
  {32'h45e33832, 32'h00000000} /* (18, 15, 26) {real, imag} */,
  {32'h45b98d87, 32'h00000000} /* (18, 15, 25) {real, imag} */,
  {32'h45c41f91, 32'h00000000} /* (18, 15, 24) {real, imag} */,
  {32'h458f4642, 32'h00000000} /* (18, 15, 23) {real, imag} */,
  {32'h4570d044, 32'h00000000} /* (18, 15, 22) {real, imag} */,
  {32'h44df5440, 32'h00000000} /* (18, 15, 21) {real, imag} */,
  {32'hc4b009de, 32'h00000000} /* (18, 15, 20) {real, imag} */,
  {32'hc582d5ee, 32'h00000000} /* (18, 15, 19) {real, imag} */,
  {32'hc5b56dab, 32'h00000000} /* (18, 15, 18) {real, imag} */,
  {32'hc5d11e8c, 32'h00000000} /* (18, 15, 17) {real, imag} */,
  {32'hc5d688b8, 32'h00000000} /* (18, 15, 16) {real, imag} */,
  {32'hc5d644ee, 32'h00000000} /* (18, 15, 15) {real, imag} */,
  {32'hc5d46d36, 32'h00000000} /* (18, 15, 14) {real, imag} */,
  {32'hc5b3ac04, 32'h00000000} /* (18, 15, 13) {real, imag} */,
  {32'hc58b6e8a, 32'h00000000} /* (18, 15, 12) {real, imag} */,
  {32'hc50c3aa9, 32'h00000000} /* (18, 15, 11) {real, imag} */,
  {32'h44d66cd6, 32'h00000000} /* (18, 15, 10) {real, imag} */,
  {32'h457f0706, 32'h00000000} /* (18, 15, 9) {real, imag} */,
  {32'h45b4f4bf, 32'h00000000} /* (18, 15, 8) {real, imag} */,
  {32'h45e28826, 32'h00000000} /* (18, 15, 7) {real, imag} */,
  {32'h45bbe70e, 32'h00000000} /* (18, 15, 6) {real, imag} */,
  {32'h45ba2d5c, 32'h00000000} /* (18, 15, 5) {real, imag} */,
  {32'h45e39814, 32'h00000000} /* (18, 15, 4) {real, imag} */,
  {32'h45e634a6, 32'h00000000} /* (18, 15, 3) {real, imag} */,
  {32'h45c1d0bf, 32'h00000000} /* (18, 15, 2) {real, imag} */,
  {32'h45f2d14e, 32'h00000000} /* (18, 15, 1) {real, imag} */,
  {32'h45d7fdd2, 32'h00000000} /* (18, 15, 0) {real, imag} */,
  {32'h45b2f7fe, 32'h00000000} /* (18, 14, 31) {real, imag} */,
  {32'h45b3600c, 32'h00000000} /* (18, 14, 30) {real, imag} */,
  {32'h45c404a6, 32'h00000000} /* (18, 14, 29) {real, imag} */,
  {32'h45c0a670, 32'h00000000} /* (18, 14, 28) {real, imag} */,
  {32'h45b73f26, 32'h00000000} /* (18, 14, 27) {real, imag} */,
  {32'h45c53314, 32'h00000000} /* (18, 14, 26) {real, imag} */,
  {32'h45a639d0, 32'h00000000} /* (18, 14, 25) {real, imag} */,
  {32'h4594aa2f, 32'h00000000} /* (18, 14, 24) {real, imag} */,
  {32'h4582946d, 32'h00000000} /* (18, 14, 23) {real, imag} */,
  {32'h45909616, 32'h00000000} /* (18, 14, 22) {real, imag} */,
  {32'h450a442a, 32'h00000000} /* (18, 14, 21) {real, imag} */,
  {32'hc4ca33a4, 32'h00000000} /* (18, 14, 20) {real, imag} */,
  {32'hc566d725, 32'h00000000} /* (18, 14, 19) {real, imag} */,
  {32'hc5b39c00, 32'h00000000} /* (18, 14, 18) {real, imag} */,
  {32'hc5b37f27, 32'h00000000} /* (18, 14, 17) {real, imag} */,
  {32'hc5b5bfda, 32'h00000000} /* (18, 14, 16) {real, imag} */,
  {32'hc5c27eac, 32'h00000000} /* (18, 14, 15) {real, imag} */,
  {32'hc5dbc1da, 32'h00000000} /* (18, 14, 14) {real, imag} */,
  {32'hc5ac4702, 32'h00000000} /* (18, 14, 13) {real, imag} */,
  {32'hc54a46f4, 32'h00000000} /* (18, 14, 12) {real, imag} */,
  {32'hc4c0a564, 32'h00000000} /* (18, 14, 11) {real, imag} */,
  {32'h44e4f844, 32'h00000000} /* (18, 14, 10) {real, imag} */,
  {32'h4592d804, 32'h00000000} /* (18, 14, 9) {real, imag} */,
  {32'h45b19175, 32'h00000000} /* (18, 14, 8) {real, imag} */,
  {32'h45b8432f, 32'h00000000} /* (18, 14, 7) {real, imag} */,
  {32'h45c0a97a, 32'h00000000} /* (18, 14, 6) {real, imag} */,
  {32'h45b64f1e, 32'h00000000} /* (18, 14, 5) {real, imag} */,
  {32'h45bebe19, 32'h00000000} /* (18, 14, 4) {real, imag} */,
  {32'h45c23e92, 32'h00000000} /* (18, 14, 3) {real, imag} */,
  {32'h45df9b0e, 32'h00000000} /* (18, 14, 2) {real, imag} */,
  {32'h45d8334b, 32'h00000000} /* (18, 14, 1) {real, imag} */,
  {32'h45bc0c22, 32'h00000000} /* (18, 14, 0) {real, imag} */,
  {32'h45885a80, 32'h00000000} /* (18, 13, 31) {real, imag} */,
  {32'h45a206de, 32'h00000000} /* (18, 13, 30) {real, imag} */,
  {32'h45a0e95a, 32'h00000000} /* (18, 13, 29) {real, imag} */,
  {32'h45aa8f09, 32'h00000000} /* (18, 13, 28) {real, imag} */,
  {32'h4592214e, 32'h00000000} /* (18, 13, 27) {real, imag} */,
  {32'h45916de1, 32'h00000000} /* (18, 13, 26) {real, imag} */,
  {32'h458c8a6d, 32'h00000000} /* (18, 13, 25) {real, imag} */,
  {32'h457698c1, 32'h00000000} /* (18, 13, 24) {real, imag} */,
  {32'h455f5ee1, 32'h00000000} /* (18, 13, 23) {real, imag} */,
  {32'h45315fab, 32'h00000000} /* (18, 13, 22) {real, imag} */,
  {32'h4494e24a, 32'h00000000} /* (18, 13, 21) {real, imag} */,
  {32'hc4f3d26a, 32'h00000000} /* (18, 13, 20) {real, imag} */,
  {32'hc563b782, 32'h00000000} /* (18, 13, 19) {real, imag} */,
  {32'hc56a620c, 32'h00000000} /* (18, 13, 18) {real, imag} */,
  {32'hc5a714c2, 32'h00000000} /* (18, 13, 17) {real, imag} */,
  {32'hc5b859cd, 32'h00000000} /* (18, 13, 16) {real, imag} */,
  {32'hc5a432e8, 32'h00000000} /* (18, 13, 15) {real, imag} */,
  {32'hc5bc6fc8, 32'h00000000} /* (18, 13, 14) {real, imag} */,
  {32'hc5802432, 32'h00000000} /* (18, 13, 13) {real, imag} */,
  {32'hc51cb8be, 32'h00000000} /* (18, 13, 12) {real, imag} */,
  {32'h42116240, 32'h00000000} /* (18, 13, 11) {real, imag} */,
  {32'h4505eab2, 32'h00000000} /* (18, 13, 10) {real, imag} */,
  {32'h456350bf, 32'h00000000} /* (18, 13, 9) {real, imag} */,
  {32'h459fe4d0, 32'h00000000} /* (18, 13, 8) {real, imag} */,
  {32'h45ac6d80, 32'h00000000} /* (18, 13, 7) {real, imag} */,
  {32'h45a96922, 32'h00000000} /* (18, 13, 6) {real, imag} */,
  {32'h45b8d4ac, 32'h00000000} /* (18, 13, 5) {real, imag} */,
  {32'h459e22b6, 32'h00000000} /* (18, 13, 4) {real, imag} */,
  {32'h45c5f28b, 32'h00000000} /* (18, 13, 3) {real, imag} */,
  {32'h45b66a1c, 32'h00000000} /* (18, 13, 2) {real, imag} */,
  {32'h45b63828, 32'h00000000} /* (18, 13, 1) {real, imag} */,
  {32'h4599806d, 32'h00000000} /* (18, 13, 0) {real, imag} */,
  {32'h45440f77, 32'h00000000} /* (18, 12, 31) {real, imag} */,
  {32'h455418d6, 32'h00000000} /* (18, 12, 30) {real, imag} */,
  {32'h455392aa, 32'h00000000} /* (18, 12, 29) {real, imag} */,
  {32'h455d64d0, 32'h00000000} /* (18, 12, 28) {real, imag} */,
  {32'h4562f9fc, 32'h00000000} /* (18, 12, 27) {real, imag} */,
  {32'h454633f8, 32'h00000000} /* (18, 12, 26) {real, imag} */,
  {32'h45267b2a, 32'h00000000} /* (18, 12, 25) {real, imag} */,
  {32'h4502c754, 32'h00000000} /* (18, 12, 24) {real, imag} */,
  {32'h4527133e, 32'h00000000} /* (18, 12, 23) {real, imag} */,
  {32'h4505417e, 32'h00000000} /* (18, 12, 22) {real, imag} */,
  {32'h446c8260, 32'h00000000} /* (18, 12, 21) {real, imag} */,
  {32'hc4659bf6, 32'h00000000} /* (18, 12, 20) {real, imag} */,
  {32'hc5508d2c, 32'h00000000} /* (18, 12, 19) {real, imag} */,
  {32'hc5450c40, 32'h00000000} /* (18, 12, 18) {real, imag} */,
  {32'hc57bc760, 32'h00000000} /* (18, 12, 17) {real, imag} */,
  {32'hc591d88e, 32'h00000000} /* (18, 12, 16) {real, imag} */,
  {32'hc5886c6c, 32'h00000000} /* (18, 12, 15) {real, imag} */,
  {32'hc57e4c8e, 32'h00000000} /* (18, 12, 14) {real, imag} */,
  {32'hc5593a84, 32'h00000000} /* (18, 12, 13) {real, imag} */,
  {32'hc4fe0583, 32'h00000000} /* (18, 12, 12) {real, imag} */,
  {32'hc4782e0e, 32'h00000000} /* (18, 12, 11) {real, imag} */,
  {32'h44e6ecc8, 32'h00000000} /* (18, 12, 10) {real, imag} */,
  {32'h4548a6d2, 32'h00000000} /* (18, 12, 9) {real, imag} */,
  {32'h4581c163, 32'h00000000} /* (18, 12, 8) {real, imag} */,
  {32'h45a77594, 32'h00000000} /* (18, 12, 7) {real, imag} */,
  {32'h4593f6a3, 32'h00000000} /* (18, 12, 6) {real, imag} */,
  {32'h4592ac22, 32'h00000000} /* (18, 12, 5) {real, imag} */,
  {32'h4584c736, 32'h00000000} /* (18, 12, 4) {real, imag} */,
  {32'h45998338, 32'h00000000} /* (18, 12, 3) {real, imag} */,
  {32'h4555e246, 32'h00000000} /* (18, 12, 2) {real, imag} */,
  {32'h45708f70, 32'h00000000} /* (18, 12, 1) {real, imag} */,
  {32'h45743ac4, 32'h00000000} /* (18, 12, 0) {real, imag} */,
  {32'h4491960e, 32'h00000000} /* (18, 11, 31) {real, imag} */,
  {32'h44b5b34c, 32'h00000000} /* (18, 11, 30) {real, imag} */,
  {32'h443742c7, 32'h00000000} /* (18, 11, 29) {real, imag} */,
  {32'h44af28d6, 32'h00000000} /* (18, 11, 28) {real, imag} */,
  {32'h43ee8bba, 32'h00000000} /* (18, 11, 27) {real, imag} */,
  {32'h43f4f9f0, 32'h00000000} /* (18, 11, 26) {real, imag} */,
  {32'h4471a814, 32'h00000000} /* (18, 11, 25) {real, imag} */,
  {32'h442e3663, 32'h00000000} /* (18, 11, 24) {real, imag} */,
  {32'h449aa117, 32'h00000000} /* (18, 11, 23) {real, imag} */,
  {32'h44b7e4aa, 32'h00000000} /* (18, 11, 22) {real, imag} */,
  {32'h4416e988, 32'h00000000} /* (18, 11, 21) {real, imag} */,
  {32'hc4c460dc, 32'h00000000} /* (18, 11, 20) {real, imag} */,
  {32'hc4dc2656, 32'h00000000} /* (18, 11, 19) {real, imag} */,
  {32'hc4f28b7a, 32'h00000000} /* (18, 11, 18) {real, imag} */,
  {32'hc50e79d0, 32'h00000000} /* (18, 11, 17) {real, imag} */,
  {32'hc4fbc62d, 32'h00000000} /* (18, 11, 16) {real, imag} */,
  {32'hc4c4b348, 32'h00000000} /* (18, 11, 15) {real, imag} */,
  {32'hc53497f0, 32'h00000000} /* (18, 11, 14) {real, imag} */,
  {32'hc4c90114, 32'h00000000} /* (18, 11, 13) {real, imag} */,
  {32'h433388b4, 32'h00000000} /* (18, 11, 12) {real, imag} */,
  {32'h42b89b18, 32'h00000000} /* (18, 11, 11) {real, imag} */,
  {32'h45045afa, 32'h00000000} /* (18, 11, 10) {real, imag} */,
  {32'h450c8c79, 32'h00000000} /* (18, 11, 9) {real, imag} */,
  {32'h4514300c, 32'h00000000} /* (18, 11, 8) {real, imag} */,
  {32'h454aaba8, 32'h00000000} /* (18, 11, 7) {real, imag} */,
  {32'h454b64bd, 32'h00000000} /* (18, 11, 6) {real, imag} */,
  {32'h45245546, 32'h00000000} /* (18, 11, 5) {real, imag} */,
  {32'h45208452, 32'h00000000} /* (18, 11, 4) {real, imag} */,
  {32'h44d33f46, 32'h00000000} /* (18, 11, 3) {real, imag} */,
  {32'h45282b33, 32'h00000000} /* (18, 11, 2) {real, imag} */,
  {32'h451d0376, 32'h00000000} /* (18, 11, 1) {real, imag} */,
  {32'h4474c23e, 32'h00000000} /* (18, 11, 0) {real, imag} */,
  {32'hc4d8d3a2, 32'h00000000} /* (18, 10, 31) {real, imag} */,
  {32'hc508e724, 32'h00000000} /* (18, 10, 30) {real, imag} */,
  {32'hc50df346, 32'h00000000} /* (18, 10, 29) {real, imag} */,
  {32'hc518f7bc, 32'h00000000} /* (18, 10, 28) {real, imag} */,
  {32'hc55794c8, 32'h00000000} /* (18, 10, 27) {real, imag} */,
  {32'hc52d0be2, 32'h00000000} /* (18, 10, 26) {real, imag} */,
  {32'hc527a244, 32'h00000000} /* (18, 10, 25) {real, imag} */,
  {32'hc5263746, 32'h00000000} /* (18, 10, 24) {real, imag} */,
  {32'hc52add12, 32'h00000000} /* (18, 10, 23) {real, imag} */,
  {32'hc4d1693c, 32'h00000000} /* (18, 10, 22) {real, imag} */,
  {32'hc490181f, 32'h00000000} /* (18, 10, 21) {real, imag} */,
  {32'hc4157502, 32'h00000000} /* (18, 10, 20) {real, imag} */,
  {32'hc370c114, 32'h00000000} /* (18, 10, 19) {real, imag} */,
  {32'h4362ed7a, 32'h00000000} /* (18, 10, 18) {real, imag} */,
  {32'h4463a42c, 32'h00000000} /* (18, 10, 17) {real, imag} */,
  {32'h448e85e0, 32'h00000000} /* (18, 10, 16) {real, imag} */,
  {32'h44c95354, 32'h00000000} /* (18, 10, 15) {real, imag} */,
  {32'h44cbfd4a, 32'h00000000} /* (18, 10, 14) {real, imag} */,
  {32'h451e9ece, 32'h00000000} /* (18, 10, 13) {real, imag} */,
  {32'h44f3aefc, 32'h00000000} /* (18, 10, 12) {real, imag} */,
  {32'h45149006, 32'h00000000} /* (18, 10, 11) {real, imag} */,
  {32'hc13cc780, 32'h00000000} /* (18, 10, 10) {real, imag} */,
  {32'hc3af542c, 32'h00000000} /* (18, 10, 9) {real, imag} */,
  {32'h42ee46d0, 32'h00000000} /* (18, 10, 8) {real, imag} */,
  {32'hc45cb051, 32'h00000000} /* (18, 10, 7) {real, imag} */,
  {32'hc41ba9a8, 32'h00000000} /* (18, 10, 6) {real, imag} */,
  {32'hc47a82e2, 32'h00000000} /* (18, 10, 5) {real, imag} */,
  {32'hc4d86cf7, 32'h00000000} /* (18, 10, 4) {real, imag} */,
  {32'hc43bb575, 32'h00000000} /* (18, 10, 3) {real, imag} */,
  {32'hc36c23ba, 32'h00000000} /* (18, 10, 2) {real, imag} */,
  {32'hc4fa1256, 32'h00000000} /* (18, 10, 1) {real, imag} */,
  {32'hc4f48214, 32'h00000000} /* (18, 10, 0) {real, imag} */,
  {32'hc56aab42, 32'h00000000} /* (18, 9, 31) {real, imag} */,
  {32'hc5a2f6e0, 32'h00000000} /* (18, 9, 30) {real, imag} */,
  {32'hc5a05eb2, 32'h00000000} /* (18, 9, 29) {real, imag} */,
  {32'hc5aeeac8, 32'h00000000} /* (18, 9, 28) {real, imag} */,
  {32'hc5b14108, 32'h00000000} /* (18, 9, 27) {real, imag} */,
  {32'hc5ae7dea, 32'h00000000} /* (18, 9, 26) {real, imag} */,
  {32'hc5b09036, 32'h00000000} /* (18, 9, 25) {real, imag} */,
  {32'hc5b5b569, 32'h00000000} /* (18, 9, 24) {real, imag} */,
  {32'hc56b277a, 32'h00000000} /* (18, 9, 23) {real, imag} */,
  {32'hc55824aa, 32'h00000000} /* (18, 9, 22) {real, imag} */,
  {32'hc5027e52, 32'h00000000} /* (18, 9, 21) {real, imag} */,
  {32'hc3fa4c68, 32'h00000000} /* (18, 9, 20) {real, imag} */,
  {32'h4427c336, 32'h00000000} /* (18, 9, 19) {real, imag} */,
  {32'h453667a8, 32'h00000000} /* (18, 9, 18) {real, imag} */,
  {32'h45563764, 32'h00000000} /* (18, 9, 17) {real, imag} */,
  {32'h457be98b, 32'h00000000} /* (18, 9, 16) {real, imag} */,
  {32'h4589cb4f, 32'h00000000} /* (18, 9, 15) {real, imag} */,
  {32'h4585de4a, 32'h00000000} /* (18, 9, 14) {real, imag} */,
  {32'h4570ac18, 32'h00000000} /* (18, 9, 13) {real, imag} */,
  {32'h454361db, 32'h00000000} /* (18, 9, 12) {real, imag} */,
  {32'h451d9227, 32'h00000000} /* (18, 9, 11) {real, imag} */,
  {32'h428f7020, 32'h00000000} /* (18, 9, 10) {real, imag} */,
  {32'hc4f7681f, 32'h00000000} /* (18, 9, 9) {real, imag} */,
  {32'hc506e060, 32'h00000000} /* (18, 9, 8) {real, imag} */,
  {32'hc5124aa2, 32'h00000000} /* (18, 9, 7) {real, imag} */,
  {32'hc52a27e4, 32'h00000000} /* (18, 9, 6) {real, imag} */,
  {32'hc56b35be, 32'h00000000} /* (18, 9, 5) {real, imag} */,
  {32'hc59796ea, 32'h00000000} /* (18, 9, 4) {real, imag} */,
  {32'hc5554366, 32'h00000000} /* (18, 9, 3) {real, imag} */,
  {32'hc569d9f8, 32'h00000000} /* (18, 9, 2) {real, imag} */,
  {32'hc5a09736, 32'h00000000} /* (18, 9, 1) {real, imag} */,
  {32'hc58e9d1c, 32'h00000000} /* (18, 9, 0) {real, imag} */,
  {32'hc5bf411c, 32'h00000000} /* (18, 8, 31) {real, imag} */,
  {32'hc5dbb8a7, 32'h00000000} /* (18, 8, 30) {real, imag} */,
  {32'hc5f408f6, 32'h00000000} /* (18, 8, 29) {real, imag} */,
  {32'hc60808b1, 32'h00000000} /* (18, 8, 28) {real, imag} */,
  {32'hc5e89e4a, 32'h00000000} /* (18, 8, 27) {real, imag} */,
  {32'hc5e23d33, 32'h00000000} /* (18, 8, 26) {real, imag} */,
  {32'hc5dc150d, 32'h00000000} /* (18, 8, 25) {real, imag} */,
  {32'hc5ade58c, 32'h00000000} /* (18, 8, 24) {real, imag} */,
  {32'hc59f6c1e, 32'h00000000} /* (18, 8, 23) {real, imag} */,
  {32'hc58d02a0, 32'h00000000} /* (18, 8, 22) {real, imag} */,
  {32'hc5238e3d, 32'h00000000} /* (18, 8, 21) {real, imag} */,
  {32'hc3c30ba8, 32'h00000000} /* (18, 8, 20) {real, imag} */,
  {32'h443cf740, 32'h00000000} /* (18, 8, 19) {real, imag} */,
  {32'h452b5048, 32'h00000000} /* (18, 8, 18) {real, imag} */,
  {32'h4564d3a9, 32'h00000000} /* (18, 8, 17) {real, imag} */,
  {32'h458fe646, 32'h00000000} /* (18, 8, 16) {real, imag} */,
  {32'h459b3cee, 32'h00000000} /* (18, 8, 15) {real, imag} */,
  {32'h459b57f1, 32'h00000000} /* (18, 8, 14) {real, imag} */,
  {32'h4589c62e, 32'h00000000} /* (18, 8, 13) {real, imag} */,
  {32'h457b7407, 32'h00000000} /* (18, 8, 12) {real, imag} */,
  {32'h453bea0c, 32'h00000000} /* (18, 8, 11) {real, imag} */,
  {32'h4408b6c8, 32'h00000000} /* (18, 8, 10) {real, imag} */,
  {32'hc4ca6e6c, 32'h00000000} /* (18, 8, 9) {real, imag} */,
  {32'hc50bb7e9, 32'h00000000} /* (18, 8, 8) {real, imag} */,
  {32'hc521a78b, 32'h00000000} /* (18, 8, 7) {real, imag} */,
  {32'hc577c1a9, 32'h00000000} /* (18, 8, 6) {real, imag} */,
  {32'hc59d327c, 32'h00000000} /* (18, 8, 5) {real, imag} */,
  {32'hc59ee0ea, 32'h00000000} /* (18, 8, 4) {real, imag} */,
  {32'hc5b4b8b2, 32'h00000000} /* (18, 8, 3) {real, imag} */,
  {32'hc5c5ca50, 32'h00000000} /* (18, 8, 2) {real, imag} */,
  {32'hc5a795ec, 32'h00000000} /* (18, 8, 1) {real, imag} */,
  {32'hc5cc0f52, 32'h00000000} /* (18, 8, 0) {real, imag} */,
  {32'hc5eb3577, 32'h00000000} /* (18, 7, 31) {real, imag} */,
  {32'hc5fc045f, 32'h00000000} /* (18, 7, 30) {real, imag} */,
  {32'hc6013bfa, 32'h00000000} /* (18, 7, 29) {real, imag} */,
  {32'hc6061e79, 32'h00000000} /* (18, 7, 28) {real, imag} */,
  {32'hc6053d2e, 32'h00000000} /* (18, 7, 27) {real, imag} */,
  {32'hc6049823, 32'h00000000} /* (18, 7, 26) {real, imag} */,
  {32'hc614a47e, 32'h00000000} /* (18, 7, 25) {real, imag} */,
  {32'hc5f3f870, 32'h00000000} /* (18, 7, 24) {real, imag} */,
  {32'hc5ca1f18, 32'h00000000} /* (18, 7, 23) {real, imag} */,
  {32'hc5a126b6, 32'h00000000} /* (18, 7, 22) {real, imag} */,
  {32'hc5994685, 32'h00000000} /* (18, 7, 21) {real, imag} */,
  {32'hc482988a, 32'h00000000} /* (18, 7, 20) {real, imag} */,
  {32'h445c43bc, 32'h00000000} /* (18, 7, 19) {real, imag} */,
  {32'h454b0d27, 32'h00000000} /* (18, 7, 18) {real, imag} */,
  {32'h4576ee34, 32'h00000000} /* (18, 7, 17) {real, imag} */,
  {32'h45909fc5, 32'h00000000} /* (18, 7, 16) {real, imag} */,
  {32'h45bc94e7, 32'h00000000} /* (18, 7, 15) {real, imag} */,
  {32'h459a0641, 32'h00000000} /* (18, 7, 14) {real, imag} */,
  {32'h45999013, 32'h00000000} /* (18, 7, 13) {real, imag} */,
  {32'h4598d800, 32'h00000000} /* (18, 7, 12) {real, imag} */,
  {32'h4588c14d, 32'h00000000} /* (18, 7, 11) {real, imag} */,
  {32'h43f73be8, 32'h00000000} /* (18, 7, 10) {real, imag} */,
  {32'hc4ba9352, 32'h00000000} /* (18, 7, 9) {real, imag} */,
  {32'hc51012fc, 32'h00000000} /* (18, 7, 8) {real, imag} */,
  {32'hc528a310, 32'h00000000} /* (18, 7, 7) {real, imag} */,
  {32'hc59d849c, 32'h00000000} /* (18, 7, 6) {real, imag} */,
  {32'hc5ad0505, 32'h00000000} /* (18, 7, 5) {real, imag} */,
  {32'hc5b19906, 32'h00000000} /* (18, 7, 4) {real, imag} */,
  {32'hc5b70ce6, 32'h00000000} /* (18, 7, 3) {real, imag} */,
  {32'hc5c47f9c, 32'h00000000} /* (18, 7, 2) {real, imag} */,
  {32'hc5f134e2, 32'h00000000} /* (18, 7, 1) {real, imag} */,
  {32'hc5df9beb, 32'h00000000} /* (18, 7, 0) {real, imag} */,
  {32'hc5f54bb9, 32'h00000000} /* (18, 6, 31) {real, imag} */,
  {32'hc613eb45, 32'h00000000} /* (18, 6, 30) {real, imag} */,
  {32'hc6123eaa, 32'h00000000} /* (18, 6, 29) {real, imag} */,
  {32'hc5f5dd3e, 32'h00000000} /* (18, 6, 28) {real, imag} */,
  {32'hc5f92edb, 32'h00000000} /* (18, 6, 27) {real, imag} */,
  {32'hc60bf1c8, 32'h00000000} /* (18, 6, 26) {real, imag} */,
  {32'hc61ab6cc, 32'h00000000} /* (18, 6, 25) {real, imag} */,
  {32'hc6072024, 32'h00000000} /* (18, 6, 24) {real, imag} */,
  {32'hc5f59f1d, 32'h00000000} /* (18, 6, 23) {real, imag} */,
  {32'hc5d4d656, 32'h00000000} /* (18, 6, 22) {real, imag} */,
  {32'hc5bc6ed0, 32'h00000000} /* (18, 6, 21) {real, imag} */,
  {32'hc511ee1a, 32'h00000000} /* (18, 6, 20) {real, imag} */,
  {32'h43b5d390, 32'h00000000} /* (18, 6, 19) {real, imag} */,
  {32'h44e4d3e4, 32'h00000000} /* (18, 6, 18) {real, imag} */,
  {32'h45602682, 32'h00000000} /* (18, 6, 17) {real, imag} */,
  {32'h4569a048, 32'h00000000} /* (18, 6, 16) {real, imag} */,
  {32'h45ad750f, 32'h00000000} /* (18, 6, 15) {real, imag} */,
  {32'h45b1a7d1, 32'h00000000} /* (18, 6, 14) {real, imag} */,
  {32'h45acca18, 32'h00000000} /* (18, 6, 13) {real, imag} */,
  {32'h45b49780, 32'h00000000} /* (18, 6, 12) {real, imag} */,
  {32'h457c22fa, 32'h00000000} /* (18, 6, 11) {real, imag} */,
  {32'h4514566e, 32'h00000000} /* (18, 6, 10) {real, imag} */,
  {32'h442f3ac0, 32'h00000000} /* (18, 6, 9) {real, imag} */,
  {32'hc487b700, 32'h00000000} /* (18, 6, 8) {real, imag} */,
  {32'hc4fecaac, 32'h00000000} /* (18, 6, 7) {real, imag} */,
  {32'hc560e7c5, 32'h00000000} /* (18, 6, 6) {real, imag} */,
  {32'hc5ab207c, 32'h00000000} /* (18, 6, 5) {real, imag} */,
  {32'hc5c808f5, 32'h00000000} /* (18, 6, 4) {real, imag} */,
  {32'hc5f50771, 32'h00000000} /* (18, 6, 3) {real, imag} */,
  {32'hc60aef94, 32'h00000000} /* (18, 6, 2) {real, imag} */,
  {32'hc5f17aab, 32'h00000000} /* (18, 6, 1) {real, imag} */,
  {32'hc5f2b22c, 32'h00000000} /* (18, 6, 0) {real, imag} */,
  {32'hc605789e, 32'h00000000} /* (18, 5, 31) {real, imag} */,
  {32'hc608f057, 32'h00000000} /* (18, 5, 30) {real, imag} */,
  {32'hc61ec60d, 32'h00000000} /* (18, 5, 29) {real, imag} */,
  {32'hc6143ec4, 32'h00000000} /* (18, 5, 28) {real, imag} */,
  {32'hc6072bfa, 32'h00000000} /* (18, 5, 27) {real, imag} */,
  {32'hc60ca672, 32'h00000000} /* (18, 5, 26) {real, imag} */,
  {32'hc61559a2, 32'h00000000} /* (18, 5, 25) {real, imag} */,
  {32'hc603cb6c, 32'h00000000} /* (18, 5, 24) {real, imag} */,
  {32'hc60aba50, 32'h00000000} /* (18, 5, 23) {real, imag} */,
  {32'hc601bc5c, 32'h00000000} /* (18, 5, 22) {real, imag} */,
  {32'hc5a2d2ee, 32'h00000000} /* (18, 5, 21) {real, imag} */,
  {32'hc58c18e4, 32'h00000000} /* (18, 5, 20) {real, imag} */,
  {32'hc553cea2, 32'h00000000} /* (18, 5, 19) {real, imag} */,
  {32'hc4a7d230, 32'h00000000} /* (18, 5, 18) {real, imag} */,
  {32'h443a0b90, 32'h00000000} /* (18, 5, 17) {real, imag} */,
  {32'h45237ee8, 32'h00000000} /* (18, 5, 16) {real, imag} */,
  {32'h4576f1e8, 32'h00000000} /* (18, 5, 15) {real, imag} */,
  {32'h4590122a, 32'h00000000} /* (18, 5, 14) {real, imag} */,
  {32'h45b95a1a, 32'h00000000} /* (18, 5, 13) {real, imag} */,
  {32'h45a4ffc0, 32'h00000000} /* (18, 5, 12) {real, imag} */,
  {32'h458bfa72, 32'h00000000} /* (18, 5, 11) {real, imag} */,
  {32'h4584c393, 32'h00000000} /* (18, 5, 10) {real, imag} */,
  {32'h4506744a, 32'h00000000} /* (18, 5, 9) {real, imag} */,
  {32'h447b08d8, 32'h00000000} /* (18, 5, 8) {real, imag} */,
  {32'hc3a006a0, 32'h00000000} /* (18, 5, 7) {real, imag} */,
  {32'hc527af0a, 32'h00000000} /* (18, 5, 6) {real, imag} */,
  {32'hc5791368, 32'h00000000} /* (18, 5, 5) {real, imag} */,
  {32'hc5c30274, 32'h00000000} /* (18, 5, 4) {real, imag} */,
  {32'hc5f82a37, 32'h00000000} /* (18, 5, 3) {real, imag} */,
  {32'hc601e73f, 32'h00000000} /* (18, 5, 2) {real, imag} */,
  {32'hc6012212, 32'h00000000} /* (18, 5, 1) {real, imag} */,
  {32'hc5fb964a, 32'h00000000} /* (18, 5, 0) {real, imag} */,
  {32'hc6050060, 32'h00000000} /* (18, 4, 31) {real, imag} */,
  {32'hc619aab4, 32'h00000000} /* (18, 4, 30) {real, imag} */,
  {32'hc6264ede, 32'h00000000} /* (18, 4, 29) {real, imag} */,
  {32'hc615b5d8, 32'h00000000} /* (18, 4, 28) {real, imag} */,
  {32'hc609efd6, 32'h00000000} /* (18, 4, 27) {real, imag} */,
  {32'hc60bc2fe, 32'h00000000} /* (18, 4, 26) {real, imag} */,
  {32'hc607afe5, 32'h00000000} /* (18, 4, 25) {real, imag} */,
  {32'hc60c35ca, 32'h00000000} /* (18, 4, 24) {real, imag} */,
  {32'hc6115c3b, 32'h00000000} /* (18, 4, 23) {real, imag} */,
  {32'hc6018e3e, 32'h00000000} /* (18, 4, 22) {real, imag} */,
  {32'hc5f19ff0, 32'h00000000} /* (18, 4, 21) {real, imag} */,
  {32'hc5b9405c, 32'h00000000} /* (18, 4, 20) {real, imag} */,
  {32'hc5a47e13, 32'h00000000} /* (18, 4, 19) {real, imag} */,
  {32'hc5378b25, 32'h00000000} /* (18, 4, 18) {real, imag} */,
  {32'hc4c960bc, 32'h00000000} /* (18, 4, 17) {real, imag} */,
  {32'h44a821b6, 32'h00000000} /* (18, 4, 16) {real, imag} */,
  {32'h4551b42f, 32'h00000000} /* (18, 4, 15) {real, imag} */,
  {32'h4583afc6, 32'h00000000} /* (18, 4, 14) {real, imag} */,
  {32'h45a32309, 32'h00000000} /* (18, 4, 13) {real, imag} */,
  {32'h45b55e41, 32'h00000000} /* (18, 4, 12) {real, imag} */,
  {32'h45bd4761, 32'h00000000} /* (18, 4, 11) {real, imag} */,
  {32'h45a59240, 32'h00000000} /* (18, 4, 10) {real, imag} */,
  {32'h458caa5e, 32'h00000000} /* (18, 4, 9) {real, imag} */,
  {32'h451ea317, 32'h00000000} /* (18, 4, 8) {real, imag} */,
  {32'h44c612be, 32'h00000000} /* (18, 4, 7) {real, imag} */,
  {32'hc46127b8, 32'h00000000} /* (18, 4, 6) {real, imag} */,
  {32'hc5829e6e, 32'h00000000} /* (18, 4, 5) {real, imag} */,
  {32'hc5d4242c, 32'h00000000} /* (18, 4, 4) {real, imag} */,
  {32'hc5f31c17, 32'h00000000} /* (18, 4, 3) {real, imag} */,
  {32'hc5e81e76, 32'h00000000} /* (18, 4, 2) {real, imag} */,
  {32'hc60316cc, 32'h00000000} /* (18, 4, 1) {real, imag} */,
  {32'hc5f8653c, 32'h00000000} /* (18, 4, 0) {real, imag} */,
  {32'hc608f1a6, 32'h00000000} /* (18, 3, 31) {real, imag} */,
  {32'hc6162b73, 32'h00000000} /* (18, 3, 30) {real, imag} */,
  {32'hc6141361, 32'h00000000} /* (18, 3, 29) {real, imag} */,
  {32'hc60db355, 32'h00000000} /* (18, 3, 28) {real, imag} */,
  {32'hc60d2daa, 32'h00000000} /* (18, 3, 27) {real, imag} */,
  {32'hc607fb4f, 32'h00000000} /* (18, 3, 26) {real, imag} */,
  {32'hc60f8709, 32'h00000000} /* (18, 3, 25) {real, imag} */,
  {32'hc6067e67, 32'h00000000} /* (18, 3, 24) {real, imag} */,
  {32'hc60f0406, 32'h00000000} /* (18, 3, 23) {real, imag} */,
  {32'hc6122d0c, 32'h00000000} /* (18, 3, 22) {real, imag} */,
  {32'hc5ea30f4, 32'h00000000} /* (18, 3, 21) {real, imag} */,
  {32'hc5b80ad5, 32'h00000000} /* (18, 3, 20) {real, imag} */,
  {32'hc5a54c9c, 32'h00000000} /* (18, 3, 19) {real, imag} */,
  {32'hc57bac7d, 32'h00000000} /* (18, 3, 18) {real, imag} */,
  {32'hc51e28b8, 32'h00000000} /* (18, 3, 17) {real, imag} */,
  {32'h42858040, 32'h00000000} /* (18, 3, 16) {real, imag} */,
  {32'h453f8739, 32'h00000000} /* (18, 3, 15) {real, imag} */,
  {32'h4599293a, 32'h00000000} /* (18, 3, 14) {real, imag} */,
  {32'h45af678e, 32'h00000000} /* (18, 3, 13) {real, imag} */,
  {32'h45d1e7b6, 32'h00000000} /* (18, 3, 12) {real, imag} */,
  {32'h45b9b0a9, 32'h00000000} /* (18, 3, 11) {real, imag} */,
  {32'h459eb5a2, 32'h00000000} /* (18, 3, 10) {real, imag} */,
  {32'h45963004, 32'h00000000} /* (18, 3, 9) {real, imag} */,
  {32'h454ef044, 32'h00000000} /* (18, 3, 8) {real, imag} */,
  {32'h44c3820e, 32'h00000000} /* (18, 3, 7) {real, imag} */,
  {32'hc270b680, 32'h00000000} /* (18, 3, 6) {real, imag} */,
  {32'hc54762cf, 32'h00000000} /* (18, 3, 5) {real, imag} */,
  {32'hc5c69ee7, 32'h00000000} /* (18, 3, 4) {real, imag} */,
  {32'hc5e9093e, 32'h00000000} /* (18, 3, 3) {real, imag} */,
  {32'hc5ffc2be, 32'h00000000} /* (18, 3, 2) {real, imag} */,
  {32'hc60a619a, 32'h00000000} /* (18, 3, 1) {real, imag} */,
  {32'hc5ff9705, 32'h00000000} /* (18, 3, 0) {real, imag} */,
  {32'hc608d019, 32'h00000000} /* (18, 2, 31) {real, imag} */,
  {32'hc61aeca6, 32'h00000000} /* (18, 2, 30) {real, imag} */,
  {32'hc60df6c3, 32'h00000000} /* (18, 2, 29) {real, imag} */,
  {32'hc6131d4f, 32'h00000000} /* (18, 2, 28) {real, imag} */,
  {32'hc619de2b, 32'h00000000} /* (18, 2, 27) {real, imag} */,
  {32'hc61085ee, 32'h00000000} /* (18, 2, 26) {real, imag} */,
  {32'hc610af58, 32'h00000000} /* (18, 2, 25) {real, imag} */,
  {32'hc60866ea, 32'h00000000} /* (18, 2, 24) {real, imag} */,
  {32'hc60dd2d4, 32'h00000000} /* (18, 2, 23) {real, imag} */,
  {32'hc6007490, 32'h00000000} /* (18, 2, 22) {real, imag} */,
  {32'hc5da39aa, 32'h00000000} /* (18, 2, 21) {real, imag} */,
  {32'hc5bb0777, 32'h00000000} /* (18, 2, 20) {real, imag} */,
  {32'hc5c46748, 32'h00000000} /* (18, 2, 19) {real, imag} */,
  {32'hc598ebf8, 32'h00000000} /* (18, 2, 18) {real, imag} */,
  {32'hc51ac3be, 32'h00000000} /* (18, 2, 17) {real, imag} */,
  {32'hc4677314, 32'h00000000} /* (18, 2, 16) {real, imag} */,
  {32'h453dbe3c, 32'h00000000} /* (18, 2, 15) {real, imag} */,
  {32'h457ac011, 32'h00000000} /* (18, 2, 14) {real, imag} */,
  {32'h45b6c624, 32'h00000000} /* (18, 2, 13) {real, imag} */,
  {32'h45b568fe, 32'h00000000} /* (18, 2, 12) {real, imag} */,
  {32'h45a0c45c, 32'h00000000} /* (18, 2, 11) {real, imag} */,
  {32'h45a5ab44, 32'h00000000} /* (18, 2, 10) {real, imag} */,
  {32'h457a296a, 32'h00000000} /* (18, 2, 9) {real, imag} */,
  {32'h4561e8d6, 32'h00000000} /* (18, 2, 8) {real, imag} */,
  {32'h44dcb1f0, 32'h00000000} /* (18, 2, 7) {real, imag} */,
  {32'hc380cdb0, 32'h00000000} /* (18, 2, 6) {real, imag} */,
  {32'hc5805818, 32'h00000000} /* (18, 2, 5) {real, imag} */,
  {32'hc5c05c0d, 32'h00000000} /* (18, 2, 4) {real, imag} */,
  {32'hc5e171c2, 32'h00000000} /* (18, 2, 3) {real, imag} */,
  {32'hc6052598, 32'h00000000} /* (18, 2, 2) {real, imag} */,
  {32'hc60efc16, 32'h00000000} /* (18, 2, 1) {real, imag} */,
  {32'hc5ff4f92, 32'h00000000} /* (18, 2, 0) {real, imag} */,
  {32'hc60e540e, 32'h00000000} /* (18, 1, 31) {real, imag} */,
  {32'hc618d934, 32'h00000000} /* (18, 1, 30) {real, imag} */,
  {32'hc61f9c08, 32'h00000000} /* (18, 1, 29) {real, imag} */,
  {32'hc614b905, 32'h00000000} /* (18, 1, 28) {real, imag} */,
  {32'hc6146694, 32'h00000000} /* (18, 1, 27) {real, imag} */,
  {32'hc60f4e7d, 32'h00000000} /* (18, 1, 26) {real, imag} */,
  {32'hc613508e, 32'h00000000} /* (18, 1, 25) {real, imag} */,
  {32'hc60d817a, 32'h00000000} /* (18, 1, 24) {real, imag} */,
  {32'hc603c546, 32'h00000000} /* (18, 1, 23) {real, imag} */,
  {32'hc5e7a100, 32'h00000000} /* (18, 1, 22) {real, imag} */,
  {32'hc5c7d2e0, 32'h00000000} /* (18, 1, 21) {real, imag} */,
  {32'hc5ae6bac, 32'h00000000} /* (18, 1, 20) {real, imag} */,
  {32'hc5ab8b4e, 32'h00000000} /* (18, 1, 19) {real, imag} */,
  {32'hc596679e, 32'h00000000} /* (18, 1, 18) {real, imag} */,
  {32'hc5211dea, 32'h00000000} /* (18, 1, 17) {real, imag} */,
  {32'h436d3060, 32'h00000000} /* (18, 1, 16) {real, imag} */,
  {32'h453332ac, 32'h00000000} /* (18, 1, 15) {real, imag} */,
  {32'h4589f11b, 32'h00000000} /* (18, 1, 14) {real, imag} */,
  {32'h45af77e5, 32'h00000000} /* (18, 1, 13) {real, imag} */,
  {32'h45ad39ef, 32'h00000000} /* (18, 1, 12) {real, imag} */,
  {32'h45a9998c, 32'h00000000} /* (18, 1, 11) {real, imag} */,
  {32'h457e8e25, 32'h00000000} /* (18, 1, 10) {real, imag} */,
  {32'h4541b6a3, 32'h00000000} /* (18, 1, 9) {real, imag} */,
  {32'h45101954, 32'h00000000} /* (18, 1, 8) {real, imag} */,
  {32'h43cd46a0, 32'h00000000} /* (18, 1, 7) {real, imag} */,
  {32'hc4b03f7e, 32'h00000000} /* (18, 1, 6) {real, imag} */,
  {32'hc56a6f50, 32'h00000000} /* (18, 1, 5) {real, imag} */,
  {32'hc5b4e1de, 32'h00000000} /* (18, 1, 4) {real, imag} */,
  {32'hc5f39ca2, 32'h00000000} /* (18, 1, 3) {real, imag} */,
  {32'hc613687b, 32'h00000000} /* (18, 1, 2) {real, imag} */,
  {32'hc6076982, 32'h00000000} /* (18, 1, 1) {real, imag} */,
  {32'hc601bd32, 32'h00000000} /* (18, 1, 0) {real, imag} */,
  {32'hc60e3eab, 32'h00000000} /* (18, 0, 31) {real, imag} */,
  {32'hc6113fb6, 32'h00000000} /* (18, 0, 30) {real, imag} */,
  {32'hc614649e, 32'h00000000} /* (18, 0, 29) {real, imag} */,
  {32'hc613d590, 32'h00000000} /* (18, 0, 28) {real, imag} */,
  {32'hc6105b2b, 32'h00000000} /* (18, 0, 27) {real, imag} */,
  {32'hc6104d29, 32'h00000000} /* (18, 0, 26) {real, imag} */,
  {32'hc604a0f8, 32'h00000000} /* (18, 0, 25) {real, imag} */,
  {32'hc5fe694e, 32'h00000000} /* (18, 0, 24) {real, imag} */,
  {32'hc5e3295e, 32'h00000000} /* (18, 0, 23) {real, imag} */,
  {32'hc5ce6090, 32'h00000000} /* (18, 0, 22) {real, imag} */,
  {32'hc5b5702c, 32'h00000000} /* (18, 0, 21) {real, imag} */,
  {32'hc58b7e1e, 32'h00000000} /* (18, 0, 20) {real, imag} */,
  {32'hc51eb2f0, 32'h00000000} /* (18, 0, 19) {real, imag} */,
  {32'hc4e80d8e, 32'h00000000} /* (18, 0, 18) {real, imag} */,
  {32'hc420e818, 32'h00000000} /* (18, 0, 17) {real, imag} */,
  {32'h44d9c8d4, 32'h00000000} /* (18, 0, 16) {real, imag} */,
  {32'h45664893, 32'h00000000} /* (18, 0, 15) {real, imag} */,
  {32'h45872773, 32'h00000000} /* (18, 0, 14) {real, imag} */,
  {32'h459a6c90, 32'h00000000} /* (18, 0, 13) {real, imag} */,
  {32'h459e4f13, 32'h00000000} /* (18, 0, 12) {real, imag} */,
  {32'h45863e46, 32'h00000000} /* (18, 0, 11) {real, imag} */,
  {32'h453beca4, 32'h00000000} /* (18, 0, 10) {real, imag} */,
  {32'h44bfa258, 32'h00000000} /* (18, 0, 9) {real, imag} */,
  {32'h44545d60, 32'h00000000} /* (18, 0, 8) {real, imag} */,
  {32'hc43a6c7c, 32'h00000000} /* (18, 0, 7) {real, imag} */,
  {32'hc52ff0f1, 32'h00000000} /* (18, 0, 6) {real, imag} */,
  {32'hc5669247, 32'h00000000} /* (18, 0, 5) {real, imag} */,
  {32'hc5bcc46a, 32'h00000000} /* (18, 0, 4) {real, imag} */,
  {32'hc5e03fe2, 32'h00000000} /* (18, 0, 3) {real, imag} */,
  {32'hc6022d8c, 32'h00000000} /* (18, 0, 2) {real, imag} */,
  {32'hc610fd52, 32'h00000000} /* (18, 0, 1) {real, imag} */,
  {32'hc603d92e, 32'h00000000} /* (18, 0, 0) {real, imag} */,
  {32'hc5b7d743, 32'h00000000} /* (17, 31, 31) {real, imag} */,
  {32'hc5c5493a, 32'h00000000} /* (17, 31, 30) {real, imag} */,
  {32'hc5c7a22b, 32'h00000000} /* (17, 31, 29) {real, imag} */,
  {32'hc5cd7591, 32'h00000000} /* (17, 31, 28) {real, imag} */,
  {32'hc5c7399a, 32'h00000000} /* (17, 31, 27) {real, imag} */,
  {32'hc5b6b79e, 32'h00000000} /* (17, 31, 26) {real, imag} */,
  {32'hc5c46512, 32'h00000000} /* (17, 31, 25) {real, imag} */,
  {32'hc5b8c986, 32'h00000000} /* (17, 31, 24) {real, imag} */,
  {32'hc5999804, 32'h00000000} /* (17, 31, 23) {real, imag} */,
  {32'hc5839f1f, 32'h00000000} /* (17, 31, 22) {real, imag} */,
  {32'hc55e81e6, 32'h00000000} /* (17, 31, 21) {real, imag} */,
  {32'hc4e3f6de, 32'h00000000} /* (17, 31, 20) {real, imag} */,
  {32'hc40962f4, 32'h00000000} /* (17, 31, 19) {real, imag} */,
  {32'h439df550, 32'h00000000} /* (17, 31, 18) {real, imag} */,
  {32'h44f76750, 32'h00000000} /* (17, 31, 17) {real, imag} */,
  {32'h44f79276, 32'h00000000} /* (17, 31, 16) {real, imag} */,
  {32'h45591b6a, 32'h00000000} /* (17, 31, 15) {real, imag} */,
  {32'h455c37fc, 32'h00000000} /* (17, 31, 14) {real, imag} */,
  {32'h455c19ca, 32'h00000000} /* (17, 31, 13) {real, imag} */,
  {32'h454a030a, 32'h00000000} /* (17, 31, 12) {real, imag} */,
  {32'h452a6995, 32'h00000000} /* (17, 31, 11) {real, imag} */,
  {32'h44a5b3e2, 32'h00000000} /* (17, 31, 10) {real, imag} */,
  {32'hc409ec90, 32'h00000000} /* (17, 31, 9) {real, imag} */,
  {32'hc4b0d7a2, 32'h00000000} /* (17, 31, 8) {real, imag} */,
  {32'hc534cfe9, 32'h00000000} /* (17, 31, 7) {real, imag} */,
  {32'hc54bda42, 32'h00000000} /* (17, 31, 6) {real, imag} */,
  {32'hc5880bcf, 32'h00000000} /* (17, 31, 5) {real, imag} */,
  {32'hc5a10498, 32'h00000000} /* (17, 31, 4) {real, imag} */,
  {32'hc5aba4ac, 32'h00000000} /* (17, 31, 3) {real, imag} */,
  {32'hc5b6b11b, 32'h00000000} /* (17, 31, 2) {real, imag} */,
  {32'hc5b9b948, 32'h00000000} /* (17, 31, 1) {real, imag} */,
  {32'hc5b0500a, 32'h00000000} /* (17, 31, 0) {real, imag} */,
  {32'hc5c99c4a, 32'h00000000} /* (17, 30, 31) {real, imag} */,
  {32'hc5e1022d, 32'h00000000} /* (17, 30, 30) {real, imag} */,
  {32'hc5f79bfc, 32'h00000000} /* (17, 30, 29) {real, imag} */,
  {32'hc5ec1026, 32'h00000000} /* (17, 30, 28) {real, imag} */,
  {32'hc5c76440, 32'h00000000} /* (17, 30, 27) {real, imag} */,
  {32'hc5b6516e, 32'h00000000} /* (17, 30, 26) {real, imag} */,
  {32'hc5c6e41b, 32'h00000000} /* (17, 30, 25) {real, imag} */,
  {32'hc5c1bf1a, 32'h00000000} /* (17, 30, 24) {real, imag} */,
  {32'hc5a303c4, 32'h00000000} /* (17, 30, 23) {real, imag} */,
  {32'hc58778c4, 32'h00000000} /* (17, 30, 22) {real, imag} */,
  {32'hc54b58ef, 32'h00000000} /* (17, 30, 21) {real, imag} */,
  {32'h433749d0, 32'h00000000} /* (17, 30, 20) {real, imag} */,
  {32'h44e6e5d4, 32'h00000000} /* (17, 30, 19) {real, imag} */,
  {32'h4503a822, 32'h00000000} /* (17, 30, 18) {real, imag} */,
  {32'h45350826, 32'h00000000} /* (17, 30, 17) {real, imag} */,
  {32'h4570fa68, 32'h00000000} /* (17, 30, 16) {real, imag} */,
  {32'h4591a666, 32'h00000000} /* (17, 30, 15) {real, imag} */,
  {32'h458cd8ef, 32'h00000000} /* (17, 30, 14) {real, imag} */,
  {32'h458791f8, 32'h00000000} /* (17, 30, 13) {real, imag} */,
  {32'h45740b5c, 32'h00000000} /* (17, 30, 12) {real, imag} */,
  {32'h45174f60, 32'h00000000} /* (17, 30, 11) {real, imag} */,
  {32'hc3752290, 32'h00000000} /* (17, 30, 10) {real, imag} */,
  {32'hc4e7f984, 32'h00000000} /* (17, 30, 9) {real, imag} */,
  {32'hc542ce2c, 32'h00000000} /* (17, 30, 8) {real, imag} */,
  {32'hc58bd256, 32'h00000000} /* (17, 30, 7) {real, imag} */,
  {32'hc5a3c080, 32'h00000000} /* (17, 30, 6) {real, imag} */,
  {32'hc5b35588, 32'h00000000} /* (17, 30, 5) {real, imag} */,
  {32'hc5c0a414, 32'h00000000} /* (17, 30, 4) {real, imag} */,
  {32'hc5c9723f, 32'h00000000} /* (17, 30, 3) {real, imag} */,
  {32'hc5e79e65, 32'h00000000} /* (17, 30, 2) {real, imag} */,
  {32'hc5c92af1, 32'h00000000} /* (17, 30, 1) {real, imag} */,
  {32'hc5bc0e46, 32'h00000000} /* (17, 30, 0) {real, imag} */,
  {32'hc5d9372f, 32'h00000000} /* (17, 29, 31) {real, imag} */,
  {32'hc5f9309e, 32'h00000000} /* (17, 29, 30) {real, imag} */,
  {32'hc600168d, 32'h00000000} /* (17, 29, 29) {real, imag} */,
  {32'hc5ebc8f3, 32'h00000000} /* (17, 29, 28) {real, imag} */,
  {32'hc5d36a18, 32'h00000000} /* (17, 29, 27) {real, imag} */,
  {32'hc5cf56c5, 32'h00000000} /* (17, 29, 26) {real, imag} */,
  {32'hc5ca579e, 32'h00000000} /* (17, 29, 25) {real, imag} */,
  {32'hc5d87946, 32'h00000000} /* (17, 29, 24) {real, imag} */,
  {32'hc5ab2ae4, 32'h00000000} /* (17, 29, 23) {real, imag} */,
  {32'hc58c819c, 32'h00000000} /* (17, 29, 22) {real, imag} */,
  {32'hc5156958, 32'h00000000} /* (17, 29, 21) {real, imag} */,
  {32'h4485f3a0, 32'h00000000} /* (17, 29, 20) {real, imag} */,
  {32'h4504230c, 32'h00000000} /* (17, 29, 19) {real, imag} */,
  {32'h453575e3, 32'h00000000} /* (17, 29, 18) {real, imag} */,
  {32'h4595dcc1, 32'h00000000} /* (17, 29, 17) {real, imag} */,
  {32'h45ab8f14, 32'h00000000} /* (17, 29, 16) {real, imag} */,
  {32'h45a858c3, 32'h00000000} /* (17, 29, 15) {real, imag} */,
  {32'h4593ff2e, 32'h00000000} /* (17, 29, 14) {real, imag} */,
  {32'h45a9ae5a, 32'h00000000} /* (17, 29, 13) {real, imag} */,
  {32'h457dd33a, 32'h00000000} /* (17, 29, 12) {real, imag} */,
  {32'h44e33350, 32'h00000000} /* (17, 29, 11) {real, imag} */,
  {32'hc3ad58e0, 32'h00000000} /* (17, 29, 10) {real, imag} */,
  {32'hc51ea1bb, 32'h00000000} /* (17, 29, 9) {real, imag} */,
  {32'hc59e360e, 32'h00000000} /* (17, 29, 8) {real, imag} */,
  {32'hc59a94b4, 32'h00000000} /* (17, 29, 7) {real, imag} */,
  {32'hc5a9d2a8, 32'h00000000} /* (17, 29, 6) {real, imag} */,
  {32'hc5c1b8a4, 32'h00000000} /* (17, 29, 5) {real, imag} */,
  {32'hc5d4dac8, 32'h00000000} /* (17, 29, 4) {real, imag} */,
  {32'hc5d70a76, 32'h00000000} /* (17, 29, 3) {real, imag} */,
  {32'hc5e3ea06, 32'h00000000} /* (17, 29, 2) {real, imag} */,
  {32'hc5d5127d, 32'h00000000} /* (17, 29, 1) {real, imag} */,
  {32'hc5e6e0d0, 32'h00000000} /* (17, 29, 0) {real, imag} */,
  {32'hc5db7ac1, 32'h00000000} /* (17, 28, 31) {real, imag} */,
  {32'hc5f62795, 32'h00000000} /* (17, 28, 30) {real, imag} */,
  {32'hc5e7b200, 32'h00000000} /* (17, 28, 29) {real, imag} */,
  {32'hc5e07971, 32'h00000000} /* (17, 28, 28) {real, imag} */,
  {32'hc5e577f2, 32'h00000000} /* (17, 28, 27) {real, imag} */,
  {32'hc5c4d147, 32'h00000000} /* (17, 28, 26) {real, imag} */,
  {32'hc5dd2928, 32'h00000000} /* (17, 28, 25) {real, imag} */,
  {32'hc5d4536e, 32'h00000000} /* (17, 28, 24) {real, imag} */,
  {32'hc5ad7827, 32'h00000000} /* (17, 28, 23) {real, imag} */,
  {32'hc5705dd6, 32'h00000000} /* (17, 28, 22) {real, imag} */,
  {32'hc4b666e6, 32'h00000000} /* (17, 28, 21) {real, imag} */,
  {32'h43a058f0, 32'h00000000} /* (17, 28, 20) {real, imag} */,
  {32'h4511df56, 32'h00000000} /* (17, 28, 19) {real, imag} */,
  {32'h456305fd, 32'h00000000} /* (17, 28, 18) {real, imag} */,
  {32'h459c60a0, 32'h00000000} /* (17, 28, 17) {real, imag} */,
  {32'h45a2ab98, 32'h00000000} /* (17, 28, 16) {real, imag} */,
  {32'h45accced, 32'h00000000} /* (17, 28, 15) {real, imag} */,
  {32'h45a62071, 32'h00000000} /* (17, 28, 14) {real, imag} */,
  {32'h45949d1c, 32'h00000000} /* (17, 28, 13) {real, imag} */,
  {32'h4571571e, 32'h00000000} /* (17, 28, 12) {real, imag} */,
  {32'h45215e90, 32'h00000000} /* (17, 28, 11) {real, imag} */,
  {32'hc3983ec0, 32'h00000000} /* (17, 28, 10) {real, imag} */,
  {32'hc5358390, 32'h00000000} /* (17, 28, 9) {real, imag} */,
  {32'hc57d5a7c, 32'h00000000} /* (17, 28, 8) {real, imag} */,
  {32'hc5a821c3, 32'h00000000} /* (17, 28, 7) {real, imag} */,
  {32'hc5be06d9, 32'h00000000} /* (17, 28, 6) {real, imag} */,
  {32'hc5c9c20a, 32'h00000000} /* (17, 28, 5) {real, imag} */,
  {32'hc5e3a049, 32'h00000000} /* (17, 28, 4) {real, imag} */,
  {32'hc5ea188f, 32'h00000000} /* (17, 28, 3) {real, imag} */,
  {32'hc5f9f33c, 32'h00000000} /* (17, 28, 2) {real, imag} */,
  {32'hc5ed153e, 32'h00000000} /* (17, 28, 1) {real, imag} */,
  {32'hc5d3cab8, 32'h00000000} /* (17, 28, 0) {real, imag} */,
  {32'hc5ebb286, 32'h00000000} /* (17, 27, 31) {real, imag} */,
  {32'hc5f9247d, 32'h00000000} /* (17, 27, 30) {real, imag} */,
  {32'hc5d8eaa6, 32'h00000000} /* (17, 27, 29) {real, imag} */,
  {32'hc5c113d5, 32'h00000000} /* (17, 27, 28) {real, imag} */,
  {32'hc5c7abff, 32'h00000000} /* (17, 27, 27) {real, imag} */,
  {32'hc5cb5fab, 32'h00000000} /* (17, 27, 26) {real, imag} */,
  {32'hc5cec972, 32'h00000000} /* (17, 27, 25) {real, imag} */,
  {32'hc5c40ee9, 32'h00000000} /* (17, 27, 24) {real, imag} */,
  {32'hc5c8dcac, 32'h00000000} /* (17, 27, 23) {real, imag} */,
  {32'hc583a34b, 32'h00000000} /* (17, 27, 22) {real, imag} */,
  {32'hc50d8b8c, 32'h00000000} /* (17, 27, 21) {real, imag} */,
  {32'h44669118, 32'h00000000} /* (17, 27, 20) {real, imag} */,
  {32'h4516a496, 32'h00000000} /* (17, 27, 19) {real, imag} */,
  {32'h45872d8d, 32'h00000000} /* (17, 27, 18) {real, imag} */,
  {32'h45a9e577, 32'h00000000} /* (17, 27, 17) {real, imag} */,
  {32'h459e00ea, 32'h00000000} /* (17, 27, 16) {real, imag} */,
  {32'h459eec3e, 32'h00000000} /* (17, 27, 15) {real, imag} */,
  {32'h459651bf, 32'h00000000} /* (17, 27, 14) {real, imag} */,
  {32'h459432f6, 32'h00000000} /* (17, 27, 13) {real, imag} */,
  {32'h455c8bd6, 32'h00000000} /* (17, 27, 12) {real, imag} */,
  {32'h452c91e6, 32'h00000000} /* (17, 27, 11) {real, imag} */,
  {32'hc487aa74, 32'h00000000} /* (17, 27, 10) {real, imag} */,
  {32'hc552ed0d, 32'h00000000} /* (17, 27, 9) {real, imag} */,
  {32'hc58de79b, 32'h00000000} /* (17, 27, 8) {real, imag} */,
  {32'hc5c37e00, 32'h00000000} /* (17, 27, 7) {real, imag} */,
  {32'hc5d0c78b, 32'h00000000} /* (17, 27, 6) {real, imag} */,
  {32'hc5e265de, 32'h00000000} /* (17, 27, 5) {real, imag} */,
  {32'hc5f81329, 32'h00000000} /* (17, 27, 4) {real, imag} */,
  {32'hc5e3fd4b, 32'h00000000} /* (17, 27, 3) {real, imag} */,
  {32'hc5fe95d9, 32'h00000000} /* (17, 27, 2) {real, imag} */,
  {32'hc5f594a1, 32'h00000000} /* (17, 27, 1) {real, imag} */,
  {32'hc5c77c96, 32'h00000000} /* (17, 27, 0) {real, imag} */,
  {32'hc5c551c4, 32'h00000000} /* (17, 26, 31) {real, imag} */,
  {32'hc5d00ea2, 32'h00000000} /* (17, 26, 30) {real, imag} */,
  {32'hc5be2e72, 32'h00000000} /* (17, 26, 29) {real, imag} */,
  {32'hc5b81cf8, 32'h00000000} /* (17, 26, 28) {real, imag} */,
  {32'hc5bb6f2a, 32'h00000000} /* (17, 26, 27) {real, imag} */,
  {32'hc5d59f4a, 32'h00000000} /* (17, 26, 26) {real, imag} */,
  {32'hc5c38622, 32'h00000000} /* (17, 26, 25) {real, imag} */,
  {32'hc5a9092d, 32'h00000000} /* (17, 26, 24) {real, imag} */,
  {32'hc59de882, 32'h00000000} /* (17, 26, 23) {real, imag} */,
  {32'hc56c9fdc, 32'h00000000} /* (17, 26, 22) {real, imag} */,
  {32'hc4b29ace, 32'h00000000} /* (17, 26, 21) {real, imag} */,
  {32'h448621f0, 32'h00000000} /* (17, 26, 20) {real, imag} */,
  {32'h451d2843, 32'h00000000} /* (17, 26, 19) {real, imag} */,
  {32'h452df02e, 32'h00000000} /* (17, 26, 18) {real, imag} */,
  {32'h457a5975, 32'h00000000} /* (17, 26, 17) {real, imag} */,
  {32'h459100a8, 32'h00000000} /* (17, 26, 16) {real, imag} */,
  {32'h458a4602, 32'h00000000} /* (17, 26, 15) {real, imag} */,
  {32'h45a536be, 32'h00000000} /* (17, 26, 14) {real, imag} */,
  {32'h458f405e, 32'h00000000} /* (17, 26, 13) {real, imag} */,
  {32'h453431d4, 32'h00000000} /* (17, 26, 12) {real, imag} */,
  {32'h44d1fa62, 32'h00000000} /* (17, 26, 11) {real, imag} */,
  {32'hc50629b5, 32'h00000000} /* (17, 26, 10) {real, imag} */,
  {32'hc55e9e5c, 32'h00000000} /* (17, 26, 9) {real, imag} */,
  {32'hc5ac05df, 32'h00000000} /* (17, 26, 8) {real, imag} */,
  {32'hc5b38a2a, 32'h00000000} /* (17, 26, 7) {real, imag} */,
  {32'hc5c1460a, 32'h00000000} /* (17, 26, 6) {real, imag} */,
  {32'hc5d74c6a, 32'h00000000} /* (17, 26, 5) {real, imag} */,
  {32'hc5e23696, 32'h00000000} /* (17, 26, 4) {real, imag} */,
  {32'hc5e5ee24, 32'h00000000} /* (17, 26, 3) {real, imag} */,
  {32'hc5ea1115, 32'h00000000} /* (17, 26, 2) {real, imag} */,
  {32'hc5e4f8aa, 32'h00000000} /* (17, 26, 1) {real, imag} */,
  {32'hc5d8a684, 32'h00000000} /* (17, 26, 0) {real, imag} */,
  {32'hc5afd1f6, 32'h00000000} /* (17, 25, 31) {real, imag} */,
  {32'hc5cfd9ea, 32'h00000000} /* (17, 25, 30) {real, imag} */,
  {32'hc5bd14de, 32'h00000000} /* (17, 25, 29) {real, imag} */,
  {32'hc5b6283b, 32'h00000000} /* (17, 25, 28) {real, imag} */,
  {32'hc5b70516, 32'h00000000} /* (17, 25, 27) {real, imag} */,
  {32'hc5b99d41, 32'h00000000} /* (17, 25, 26) {real, imag} */,
  {32'hc5b1980e, 32'h00000000} /* (17, 25, 25) {real, imag} */,
  {32'hc5a2da8f, 32'h00000000} /* (17, 25, 24) {real, imag} */,
  {32'hc58b96c7, 32'h00000000} /* (17, 25, 23) {real, imag} */,
  {32'hc5516276, 32'h00000000} /* (17, 25, 22) {real, imag} */,
  {32'hc45445a8, 32'h00000000} /* (17, 25, 21) {real, imag} */,
  {32'h44e2d7f2, 32'h00000000} /* (17, 25, 20) {real, imag} */,
  {32'h45304a52, 32'h00000000} /* (17, 25, 19) {real, imag} */,
  {32'h452e4426, 32'h00000000} /* (17, 25, 18) {real, imag} */,
  {32'h454161e6, 32'h00000000} /* (17, 25, 17) {real, imag} */,
  {32'h458d6cae, 32'h00000000} /* (17, 25, 16) {real, imag} */,
  {32'h458dc528, 32'h00000000} /* (17, 25, 15) {real, imag} */,
  {32'h45706fdc, 32'h00000000} /* (17, 25, 14) {real, imag} */,
  {32'h455d3a08, 32'h00000000} /* (17, 25, 13) {real, imag} */,
  {32'h454c1ac6, 32'h00000000} /* (17, 25, 12) {real, imag} */,
  {32'h44fa14a6, 32'h00000000} /* (17, 25, 11) {real, imag} */,
  {32'hc50f6f1a, 32'h00000000} /* (17, 25, 10) {real, imag} */,
  {32'hc575e6dc, 32'h00000000} /* (17, 25, 9) {real, imag} */,
  {32'hc58b403d, 32'h00000000} /* (17, 25, 8) {real, imag} */,
  {32'hc59bfd5d, 32'h00000000} /* (17, 25, 7) {real, imag} */,
  {32'hc5b4308b, 32'h00000000} /* (17, 25, 6) {real, imag} */,
  {32'hc5c0cbc9, 32'h00000000} /* (17, 25, 5) {real, imag} */,
  {32'hc5bbc402, 32'h00000000} /* (17, 25, 4) {real, imag} */,
  {32'hc5ddd0f3, 32'h00000000} /* (17, 25, 3) {real, imag} */,
  {32'hc5e6ae83, 32'h00000000} /* (17, 25, 2) {real, imag} */,
  {32'hc5eb4537, 32'h00000000} /* (17, 25, 1) {real, imag} */,
  {32'hc5c51046, 32'h00000000} /* (17, 25, 0) {real, imag} */,
  {32'hc59f1aa1, 32'h00000000} /* (17, 24, 31) {real, imag} */,
  {32'hc5bce946, 32'h00000000} /* (17, 24, 30) {real, imag} */,
  {32'hc5a2ef33, 32'h00000000} /* (17, 24, 29) {real, imag} */,
  {32'hc5b911db, 32'h00000000} /* (17, 24, 28) {real, imag} */,
  {32'hc5b9a8b6, 32'h00000000} /* (17, 24, 27) {real, imag} */,
  {32'hc5c6fb30, 32'h00000000} /* (17, 24, 26) {real, imag} */,
  {32'hc59e221e, 32'h00000000} /* (17, 24, 25) {real, imag} */,
  {32'hc593fcfe, 32'h00000000} /* (17, 24, 24) {real, imag} */,
  {32'hc584ac43, 32'h00000000} /* (17, 24, 23) {real, imag} */,
  {32'hc58006bd, 32'h00000000} /* (17, 24, 22) {real, imag} */,
  {32'hc4beb5ec, 32'h00000000} /* (17, 24, 21) {real, imag} */,
  {32'h453244bc, 32'h00000000} /* (17, 24, 20) {real, imag} */,
  {32'h453cf8fa, 32'h00000000} /* (17, 24, 19) {real, imag} */,
  {32'h451de098, 32'h00000000} /* (17, 24, 18) {real, imag} */,
  {32'h45807868, 32'h00000000} /* (17, 24, 17) {real, imag} */,
  {32'h4552735c, 32'h00000000} /* (17, 24, 16) {real, imag} */,
  {32'h45562736, 32'h00000000} /* (17, 24, 15) {real, imag} */,
  {32'h45387b98, 32'h00000000} /* (17, 24, 14) {real, imag} */,
  {32'h456ac28e, 32'h00000000} /* (17, 24, 13) {real, imag} */,
  {32'h4527d7ca, 32'h00000000} /* (17, 24, 12) {real, imag} */,
  {32'h442ad860, 32'h00000000} /* (17, 24, 11) {real, imag} */,
  {32'hc53b3218, 32'h00000000} /* (17, 24, 10) {real, imag} */,
  {32'hc570a244, 32'h00000000} /* (17, 24, 9) {real, imag} */,
  {32'hc5919f14, 32'h00000000} /* (17, 24, 8) {real, imag} */,
  {32'hc59e45af, 32'h00000000} /* (17, 24, 7) {real, imag} */,
  {32'hc5a71bd3, 32'h00000000} /* (17, 24, 6) {real, imag} */,
  {32'hc598ba8e, 32'h00000000} /* (17, 24, 5) {real, imag} */,
  {32'hc59f08e9, 32'h00000000} /* (17, 24, 4) {real, imag} */,
  {32'hc5cafcfb, 32'h00000000} /* (17, 24, 3) {real, imag} */,
  {32'hc5d00cc6, 32'h00000000} /* (17, 24, 2) {real, imag} */,
  {32'hc5da2fc2, 32'h00000000} /* (17, 24, 1) {real, imag} */,
  {32'hc5aec9cc, 32'h00000000} /* (17, 24, 0) {real, imag} */,
  {32'hc57c426f, 32'h00000000} /* (17, 23, 31) {real, imag} */,
  {32'hc577eac2, 32'h00000000} /* (17, 23, 30) {real, imag} */,
  {32'hc5a664ed, 32'h00000000} /* (17, 23, 29) {real, imag} */,
  {32'hc5b40052, 32'h00000000} /* (17, 23, 28) {real, imag} */,
  {32'hc5a48afb, 32'h00000000} /* (17, 23, 27) {real, imag} */,
  {32'hc5a00660, 32'h00000000} /* (17, 23, 26) {real, imag} */,
  {32'hc5988f73, 32'h00000000} /* (17, 23, 25) {real, imag} */,
  {32'hc54b4642, 32'h00000000} /* (17, 23, 24) {real, imag} */,
  {32'hc56e9d93, 32'h00000000} /* (17, 23, 23) {real, imag} */,
  {32'hc52b7e1e, 32'h00000000} /* (17, 23, 22) {real, imag} */,
  {32'hc41d2a50, 32'h00000000} /* (17, 23, 21) {real, imag} */,
  {32'h44bbeb08, 32'h00000000} /* (17, 23, 20) {real, imag} */,
  {32'h450f35ac, 32'h00000000} /* (17, 23, 19) {real, imag} */,
  {32'h4528ce69, 32'h00000000} /* (17, 23, 18) {real, imag} */,
  {32'h45339226, 32'h00000000} /* (17, 23, 17) {real, imag} */,
  {32'h45368a48, 32'h00000000} /* (17, 23, 16) {real, imag} */,
  {32'h45536ff5, 32'h00000000} /* (17, 23, 15) {real, imag} */,
  {32'h45333b06, 32'h00000000} /* (17, 23, 14) {real, imag} */,
  {32'h454f2b02, 32'h00000000} /* (17, 23, 13) {real, imag} */,
  {32'h44e0cad2, 32'h00000000} /* (17, 23, 12) {real, imag} */,
  {32'h418abf00, 32'h00000000} /* (17, 23, 11) {real, imag} */,
  {32'hc4c7c574, 32'h00000000} /* (17, 23, 10) {real, imag} */,
  {32'hc55cbb32, 32'h00000000} /* (17, 23, 9) {real, imag} */,
  {32'hc5866cbc, 32'h00000000} /* (17, 23, 8) {real, imag} */,
  {32'hc584ad9f, 32'h00000000} /* (17, 23, 7) {real, imag} */,
  {32'hc5916367, 32'h00000000} /* (17, 23, 6) {real, imag} */,
  {32'hc5975e16, 32'h00000000} /* (17, 23, 5) {real, imag} */,
  {32'hc58de41d, 32'h00000000} /* (17, 23, 4) {real, imag} */,
  {32'hc5a27d29, 32'h00000000} /* (17, 23, 3) {real, imag} */,
  {32'hc5b0a790, 32'h00000000} /* (17, 23, 2) {real, imag} */,
  {32'hc59a290e, 32'h00000000} /* (17, 23, 1) {real, imag} */,
  {32'hc5858dab, 32'h00000000} /* (17, 23, 0) {real, imag} */,
  {32'hc553f53c, 32'h00000000} /* (17, 22, 31) {real, imag} */,
  {32'hc54e1f32, 32'h00000000} /* (17, 22, 30) {real, imag} */,
  {32'hc53b898a, 32'h00000000} /* (17, 22, 29) {real, imag} */,
  {32'hc570b770, 32'h00000000} /* (17, 22, 28) {real, imag} */,
  {32'hc559a201, 32'h00000000} /* (17, 22, 27) {real, imag} */,
  {32'hc5528dc7, 32'h00000000} /* (17, 22, 26) {real, imag} */,
  {32'hc55af6b7, 32'h00000000} /* (17, 22, 25) {real, imag} */,
  {32'hc52b849f, 32'h00000000} /* (17, 22, 24) {real, imag} */,
  {32'hc52b6b51, 32'h00000000} /* (17, 22, 23) {real, imag} */,
  {32'hc526f6c8, 32'h00000000} /* (17, 22, 22) {real, imag} */,
  {32'hc4a5f3f6, 32'h00000000} /* (17, 22, 21) {real, imag} */,
  {32'h4423b55c, 32'h00000000} /* (17, 22, 20) {real, imag} */,
  {32'h44954d06, 32'h00000000} /* (17, 22, 19) {real, imag} */,
  {32'h4504f517, 32'h00000000} /* (17, 22, 18) {real, imag} */,
  {32'h4523eb84, 32'h00000000} /* (17, 22, 17) {real, imag} */,
  {32'h44f8aec1, 32'h00000000} /* (17, 22, 16) {real, imag} */,
  {32'h451c38e4, 32'h00000000} /* (17, 22, 15) {real, imag} */,
  {32'h450f6c56, 32'h00000000} /* (17, 22, 14) {real, imag} */,
  {32'h44cae6af, 32'h00000000} /* (17, 22, 13) {real, imag} */,
  {32'h449e4728, 32'h00000000} /* (17, 22, 12) {real, imag} */,
  {32'h446901f4, 32'h00000000} /* (17, 22, 11) {real, imag} */,
  {32'hc4c71e02, 32'h00000000} /* (17, 22, 10) {real, imag} */,
  {32'hc51aa385, 32'h00000000} /* (17, 22, 9) {real, imag} */,
  {32'hc5433955, 32'h00000000} /* (17, 22, 8) {real, imag} */,
  {32'hc53a5cd7, 32'h00000000} /* (17, 22, 7) {real, imag} */,
  {32'hc53ded58, 32'h00000000} /* (17, 22, 6) {real, imag} */,
  {32'hc55bfd81, 32'h00000000} /* (17, 22, 5) {real, imag} */,
  {32'hc5623539, 32'h00000000} /* (17, 22, 4) {real, imag} */,
  {32'hc541fe3d, 32'h00000000} /* (17, 22, 3) {real, imag} */,
  {32'hc57796e5, 32'h00000000} /* (17, 22, 2) {real, imag} */,
  {32'hc563ef18, 32'h00000000} /* (17, 22, 1) {real, imag} */,
  {32'hc54b4e00, 32'h00000000} /* (17, 22, 0) {real, imag} */,
  {32'hc49c6966, 32'h00000000} /* (17, 21, 31) {real, imag} */,
  {32'hc51a809e, 32'h00000000} /* (17, 21, 30) {real, imag} */,
  {32'hc4fcfd6e, 32'h00000000} /* (17, 21, 29) {real, imag} */,
  {32'hc4e8cf98, 32'h00000000} /* (17, 21, 28) {real, imag} */,
  {32'hc531a4be, 32'h00000000} /* (17, 21, 27) {real, imag} */,
  {32'hc515c24c, 32'h00000000} /* (17, 21, 26) {real, imag} */,
  {32'hc49487a5, 32'h00000000} /* (17, 21, 25) {real, imag} */,
  {32'hc4bcb86c, 32'h00000000} /* (17, 21, 24) {real, imag} */,
  {32'hc4aabc40, 32'h00000000} /* (17, 21, 23) {real, imag} */,
  {32'hc49cae96, 32'h00000000} /* (17, 21, 22) {real, imag} */,
  {32'hc46605a6, 32'h00000000} /* (17, 21, 21) {real, imag} */,
  {32'h43da21ee, 32'h00000000} /* (17, 21, 20) {real, imag} */,
  {32'h4454f66b, 32'h00000000} /* (17, 21, 19) {real, imag} */,
  {32'h44221818, 32'h00000000} /* (17, 21, 18) {real, imag} */,
  {32'h4430f628, 32'h00000000} /* (17, 21, 17) {real, imag} */,
  {32'h44058fcf, 32'h00000000} /* (17, 21, 16) {real, imag} */,
  {32'h44850b22, 32'h00000000} /* (17, 21, 15) {real, imag} */,
  {32'h443f15be, 32'h00000000} /* (17, 21, 14) {real, imag} */,
  {32'h43792f8c, 32'h00000000} /* (17, 21, 13) {real, imag} */,
  {32'h40cee680, 32'h00000000} /* (17, 21, 12) {real, imag} */,
  {32'h41bb0f40, 32'h00000000} /* (17, 21, 11) {real, imag} */,
  {32'hc43bd55a, 32'h00000000} /* (17, 21, 10) {real, imag} */,
  {32'hc4948a09, 32'h00000000} /* (17, 21, 9) {real, imag} */,
  {32'hc4929e18, 32'h00000000} /* (17, 21, 8) {real, imag} */,
  {32'hc47c0b89, 32'h00000000} /* (17, 21, 7) {real, imag} */,
  {32'hc4803218, 32'h00000000} /* (17, 21, 6) {real, imag} */,
  {32'hc35495c0, 32'h00000000} /* (17, 21, 5) {real, imag} */,
  {32'hc4946e10, 32'h00000000} /* (17, 21, 4) {real, imag} */,
  {32'hc4a03d86, 32'h00000000} /* (17, 21, 3) {real, imag} */,
  {32'hc48b3d22, 32'h00000000} /* (17, 21, 2) {real, imag} */,
  {32'hc4c16382, 32'h00000000} /* (17, 21, 1) {real, imag} */,
  {32'hc4b7d706, 32'h00000000} /* (17, 21, 0) {real, imag} */,
  {32'h4483b318, 32'h00000000} /* (17, 20, 31) {real, imag} */,
  {32'h44b40342, 32'h00000000} /* (17, 20, 30) {real, imag} */,
  {32'hc3bc6904, 32'h00000000} /* (17, 20, 29) {real, imag} */,
  {32'h437d0818, 32'h00000000} /* (17, 20, 28) {real, imag} */,
  {32'hc2b3bb38, 32'h00000000} /* (17, 20, 27) {real, imag} */,
  {32'h40e5ce00, 32'h00000000} /* (17, 20, 26) {real, imag} */,
  {32'h43ed9630, 32'h00000000} /* (17, 20, 25) {real, imag} */,
  {32'h4496f940, 32'h00000000} /* (17, 20, 24) {real, imag} */,
  {32'h43ac131a, 32'h00000000} /* (17, 20, 23) {real, imag} */,
  {32'h44615748, 32'h00000000} /* (17, 20, 22) {real, imag} */,
  {32'h43cd448a, 32'h00000000} /* (17, 20, 21) {real, imag} */,
  {32'hc4929dd1, 32'h00000000} /* (17, 20, 20) {real, imag} */,
  {32'hc22d8cb8, 32'h00000000} /* (17, 20, 19) {real, imag} */,
  {32'hc4222591, 32'h00000000} /* (17, 20, 18) {real, imag} */,
  {32'hc4790827, 32'h00000000} /* (17, 20, 17) {real, imag} */,
  {32'hc4b0f2ba, 32'h00000000} /* (17, 20, 16) {real, imag} */,
  {32'hc4712f51, 32'h00000000} /* (17, 20, 15) {real, imag} */,
  {32'hc4ea3d3c, 32'h00000000} /* (17, 20, 14) {real, imag} */,
  {32'hc4ea2c41, 32'h00000000} /* (17, 20, 13) {real, imag} */,
  {32'hc4d1b49d, 32'h00000000} /* (17, 20, 12) {real, imag} */,
  {32'hc48ce822, 32'h00000000} /* (17, 20, 11) {real, imag} */,
  {32'h43c84f7d, 32'h00000000} /* (17, 20, 10) {real, imag} */,
  {32'h44a708f5, 32'h00000000} /* (17, 20, 9) {real, imag} */,
  {32'h448719e4, 32'h00000000} /* (17, 20, 8) {real, imag} */,
  {32'h448e84a4, 32'h00000000} /* (17, 20, 7) {real, imag} */,
  {32'h44feb010, 32'h00000000} /* (17, 20, 6) {real, imag} */,
  {32'h44e833e4, 32'h00000000} /* (17, 20, 5) {real, imag} */,
  {32'h44701122, 32'h00000000} /* (17, 20, 4) {real, imag} */,
  {32'h4467f2b2, 32'h00000000} /* (17, 20, 3) {real, imag} */,
  {32'h445f431b, 32'h00000000} /* (17, 20, 2) {real, imag} */,
  {32'h449e5436, 32'h00000000} /* (17, 20, 1) {real, imag} */,
  {32'h443b765d, 32'h00000000} /* (17, 20, 0) {real, imag} */,
  {32'h44f71df0, 32'h00000000} /* (17, 19, 31) {real, imag} */,
  {32'h451e8356, 32'h00000000} /* (17, 19, 30) {real, imag} */,
  {32'h451f0021, 32'h00000000} /* (17, 19, 29) {real, imag} */,
  {32'h44b82e46, 32'h00000000} /* (17, 19, 28) {real, imag} */,
  {32'h4505c09a, 32'h00000000} /* (17, 19, 27) {real, imag} */,
  {32'h44f9d9d2, 32'h00000000} /* (17, 19, 26) {real, imag} */,
  {32'h452db08d, 32'h00000000} /* (17, 19, 25) {real, imag} */,
  {32'h45309d31, 32'h00000000} /* (17, 19, 24) {real, imag} */,
  {32'h4549bae4, 32'h00000000} /* (17, 19, 23) {real, imag} */,
  {32'h44d0c73c, 32'h00000000} /* (17, 19, 22) {real, imag} */,
  {32'h441afc26, 32'h00000000} /* (17, 19, 21) {real, imag} */,
  {32'hc44b9188, 32'h00000000} /* (17, 19, 20) {real, imag} */,
  {32'hc4fd6b2c, 32'h00000000} /* (17, 19, 19) {real, imag} */,
  {32'hc513fdc6, 32'h00000000} /* (17, 19, 18) {real, imag} */,
  {32'hc50f896c, 32'h00000000} /* (17, 19, 17) {real, imag} */,
  {32'hc532eadf, 32'h00000000} /* (17, 19, 16) {real, imag} */,
  {32'hc55886ce, 32'h00000000} /* (17, 19, 15) {real, imag} */,
  {32'hc5420f4c, 32'h00000000} /* (17, 19, 14) {real, imag} */,
  {32'hc5057e67, 32'h00000000} /* (17, 19, 13) {real, imag} */,
  {32'hc50ca839, 32'h00000000} /* (17, 19, 12) {real, imag} */,
  {32'hc4d5b574, 32'h00000000} /* (17, 19, 11) {real, imag} */,
  {32'hc32e5270, 32'h00000000} /* (17, 19, 10) {real, imag} */,
  {32'h44bba6c6, 32'h00000000} /* (17, 19, 9) {real, imag} */,
  {32'h451fa9ab, 32'h00000000} /* (17, 19, 8) {real, imag} */,
  {32'h44fd239c, 32'h00000000} /* (17, 19, 7) {real, imag} */,
  {32'h44fa2b0c, 32'h00000000} /* (17, 19, 6) {real, imag} */,
  {32'h452b1354, 32'h00000000} /* (17, 19, 5) {real, imag} */,
  {32'h453f25ac, 32'h00000000} /* (17, 19, 4) {real, imag} */,
  {32'h453f011e, 32'h00000000} /* (17, 19, 3) {real, imag} */,
  {32'h45457048, 32'h00000000} /* (17, 19, 2) {real, imag} */,
  {32'h455a9bbc, 32'h00000000} /* (17, 19, 1) {real, imag} */,
  {32'h454567e7, 32'h00000000} /* (17, 19, 0) {real, imag} */,
  {32'h455825ef, 32'h00000000} /* (17, 18, 31) {real, imag} */,
  {32'h455acbba, 32'h00000000} /* (17, 18, 30) {real, imag} */,
  {32'h4591a169, 32'h00000000} /* (17, 18, 29) {real, imag} */,
  {32'h4570f179, 32'h00000000} /* (17, 18, 28) {real, imag} */,
  {32'h455c55a8, 32'h00000000} /* (17, 18, 27) {real, imag} */,
  {32'h4538766d, 32'h00000000} /* (17, 18, 26) {real, imag} */,
  {32'h4565230a, 32'h00000000} /* (17, 18, 25) {real, imag} */,
  {32'h455f76f7, 32'h00000000} /* (17, 18, 24) {real, imag} */,
  {32'h45625245, 32'h00000000} /* (17, 18, 23) {real, imag} */,
  {32'h4509400c, 32'h00000000} /* (17, 18, 22) {real, imag} */,
  {32'h4403ec7a, 32'h00000000} /* (17, 18, 21) {real, imag} */,
  {32'hc4a9e8f2, 32'h00000000} /* (17, 18, 20) {real, imag} */,
  {32'hc558d9e7, 32'h00000000} /* (17, 18, 19) {real, imag} */,
  {32'hc5483b63, 32'h00000000} /* (17, 18, 18) {real, imag} */,
  {32'hc55f9958, 32'h00000000} /* (17, 18, 17) {real, imag} */,
  {32'hc55bc38e, 32'h00000000} /* (17, 18, 16) {real, imag} */,
  {32'hc5702387, 32'h00000000} /* (17, 18, 15) {real, imag} */,
  {32'hc54d90c2, 32'h00000000} /* (17, 18, 14) {real, imag} */,
  {32'hc5351db6, 32'h00000000} /* (17, 18, 13) {real, imag} */,
  {32'hc4d95d26, 32'h00000000} /* (17, 18, 12) {real, imag} */,
  {32'hc5135120, 32'h00000000} /* (17, 18, 11) {real, imag} */,
  {32'h449292b6, 32'h00000000} /* (17, 18, 10) {real, imag} */,
  {32'h457d234a, 32'h00000000} /* (17, 18, 9) {real, imag} */,
  {32'h45665769, 32'h00000000} /* (17, 18, 8) {real, imag} */,
  {32'h453de6cb, 32'h00000000} /* (17, 18, 7) {real, imag} */,
  {32'h45571ad4, 32'h00000000} /* (17, 18, 6) {real, imag} */,
  {32'h4544552c, 32'h00000000} /* (17, 18, 5) {real, imag} */,
  {32'h45827dc6, 32'h00000000} /* (17, 18, 4) {real, imag} */,
  {32'h4583d956, 32'h00000000} /* (17, 18, 3) {real, imag} */,
  {32'h45a24c9e, 32'h00000000} /* (17, 18, 2) {real, imag} */,
  {32'h45963c60, 32'h00000000} /* (17, 18, 1) {real, imag} */,
  {32'h457cb552, 32'h00000000} /* (17, 18, 0) {real, imag} */,
  {32'h45822a2a, 32'h00000000} /* (17, 17, 31) {real, imag} */,
  {32'h459e7acf, 32'h00000000} /* (17, 17, 30) {real, imag} */,
  {32'h4598a935, 32'h00000000} /* (17, 17, 29) {real, imag} */,
  {32'h45907188, 32'h00000000} /* (17, 17, 28) {real, imag} */,
  {32'h457a599c, 32'h00000000} /* (17, 17, 27) {real, imag} */,
  {32'h4582da48, 32'h00000000} /* (17, 17, 26) {real, imag} */,
  {32'h45763d86, 32'h00000000} /* (17, 17, 25) {real, imag} */,
  {32'h45910fd5, 32'h00000000} /* (17, 17, 24) {real, imag} */,
  {32'h45826bda, 32'h00000000} /* (17, 17, 23) {real, imag} */,
  {32'h4524b65a, 32'h00000000} /* (17, 17, 22) {real, imag} */,
  {32'h442c0460, 32'h00000000} /* (17, 17, 21) {real, imag} */,
  {32'hc4ab3c9c, 32'h00000000} /* (17, 17, 20) {real, imag} */,
  {32'hc5447f42, 32'h00000000} /* (17, 17, 19) {real, imag} */,
  {32'hc5713f00, 32'h00000000} /* (17, 17, 18) {real, imag} */,
  {32'hc58afb1a, 32'h00000000} /* (17, 17, 17) {real, imag} */,
  {32'hc599765e, 32'h00000000} /* (17, 17, 16) {real, imag} */,
  {32'hc571a9fd, 32'h00000000} /* (17, 17, 15) {real, imag} */,
  {32'hc572911e, 32'h00000000} /* (17, 17, 14) {real, imag} */,
  {32'hc54e7e88, 32'h00000000} /* (17, 17, 13) {real, imag} */,
  {32'hc528016a, 32'h00000000} /* (17, 17, 12) {real, imag} */,
  {32'hc49f41a7, 32'h00000000} /* (17, 17, 11) {real, imag} */,
  {32'h45521b5c, 32'h00000000} /* (17, 17, 10) {real, imag} */,
  {32'h457830b8, 32'h00000000} /* (17, 17, 9) {real, imag} */,
  {32'h45a07bc3, 32'h00000000} /* (17, 17, 8) {real, imag} */,
  {32'h458c73a8, 32'h00000000} /* (17, 17, 7) {real, imag} */,
  {32'h45442aa2, 32'h00000000} /* (17, 17, 6) {real, imag} */,
  {32'h458a18b6, 32'h00000000} /* (17, 17, 5) {real, imag} */,
  {32'h45896a6a, 32'h00000000} /* (17, 17, 4) {real, imag} */,
  {32'h458fbded, 32'h00000000} /* (17, 17, 3) {real, imag} */,
  {32'h459c7cb6, 32'h00000000} /* (17, 17, 2) {real, imag} */,
  {32'h4590cf56, 32'h00000000} /* (17, 17, 1) {real, imag} */,
  {32'h4586f78a, 32'h00000000} /* (17, 17, 0) {real, imag} */,
  {32'h4580136a, 32'h00000000} /* (17, 16, 31) {real, imag} */,
  {32'h4590abda, 32'h00000000} /* (17, 16, 30) {real, imag} */,
  {32'h459d5b57, 32'h00000000} /* (17, 16, 29) {real, imag} */,
  {32'h45987eea, 32'h00000000} /* (17, 16, 28) {real, imag} */,
  {32'h4590237d, 32'h00000000} /* (17, 16, 27) {real, imag} */,
  {32'h458c1b68, 32'h00000000} /* (17, 16, 26) {real, imag} */,
  {32'h4586fe5e, 32'h00000000} /* (17, 16, 25) {real, imag} */,
  {32'h457f3f71, 32'h00000000} /* (17, 16, 24) {real, imag} */,
  {32'h45769390, 32'h00000000} /* (17, 16, 23) {real, imag} */,
  {32'h45236465, 32'h00000000} /* (17, 16, 22) {real, imag} */,
  {32'h4454723e, 32'h00000000} /* (17, 16, 21) {real, imag} */,
  {32'hc4782d54, 32'h00000000} /* (17, 16, 20) {real, imag} */,
  {32'hc58174ae, 32'h00000000} /* (17, 16, 19) {real, imag} */,
  {32'hc57a618a, 32'h00000000} /* (17, 16, 18) {real, imag} */,
  {32'hc593f0e0, 32'h00000000} /* (17, 16, 17) {real, imag} */,
  {32'hc592112f, 32'h00000000} /* (17, 16, 16) {real, imag} */,
  {32'hc59ea3fa, 32'h00000000} /* (17, 16, 15) {real, imag} */,
  {32'hc579804f, 32'h00000000} /* (17, 16, 14) {real, imag} */,
  {32'hc5b0101b, 32'h00000000} /* (17, 16, 13) {real, imag} */,
  {32'hc56b584d, 32'h00000000} /* (17, 16, 12) {real, imag} */,
  {32'hc47365d8, 32'h00000000} /* (17, 16, 11) {real, imag} */,
  {32'h44eb5e04, 32'h00000000} /* (17, 16, 10) {real, imag} */,
  {32'h458b3426, 32'h00000000} /* (17, 16, 9) {real, imag} */,
  {32'h458cf9b7, 32'h00000000} /* (17, 16, 8) {real, imag} */,
  {32'h458e92d8, 32'h00000000} /* (17, 16, 7) {real, imag} */,
  {32'h45745557, 32'h00000000} /* (17, 16, 6) {real, imag} */,
  {32'h45851e97, 32'h00000000} /* (17, 16, 5) {real, imag} */,
  {32'h458725fe, 32'h00000000} /* (17, 16, 4) {real, imag} */,
  {32'h458f7502, 32'h00000000} /* (17, 16, 3) {real, imag} */,
  {32'h458a5f6f, 32'h00000000} /* (17, 16, 2) {real, imag} */,
  {32'h459b78ba, 32'h00000000} /* (17, 16, 1) {real, imag} */,
  {32'h458eb885, 32'h00000000} /* (17, 16, 0) {real, imag} */,
  {32'h457002f8, 32'h00000000} /* (17, 15, 31) {real, imag} */,
  {32'h459183ec, 32'h00000000} /* (17, 15, 30) {real, imag} */,
  {32'h4597d105, 32'h00000000} /* (17, 15, 29) {real, imag} */,
  {32'h4571b044, 32'h00000000} /* (17, 15, 28) {real, imag} */,
  {32'h4598bde6, 32'h00000000} /* (17, 15, 27) {real, imag} */,
  {32'h4591573a, 32'h00000000} /* (17, 15, 26) {real, imag} */,
  {32'h456fce06, 32'h00000000} /* (17, 15, 25) {real, imag} */,
  {32'h455d288c, 32'h00000000} /* (17, 15, 24) {real, imag} */,
  {32'h4550ae44, 32'h00000000} /* (17, 15, 23) {real, imag} */,
  {32'h45167b03, 32'h00000000} /* (17, 15, 22) {real, imag} */,
  {32'h44b6cbf1, 32'h00000000} /* (17, 15, 21) {real, imag} */,
  {32'hc4b3b1e0, 32'h00000000} /* (17, 15, 20) {real, imag} */,
  {32'hc5253d7a, 32'h00000000} /* (17, 15, 19) {real, imag} */,
  {32'hc57c751f, 32'h00000000} /* (17, 15, 18) {real, imag} */,
  {32'hc59883fa, 32'h00000000} /* (17, 15, 17) {real, imag} */,
  {32'hc586796c, 32'h00000000} /* (17, 15, 16) {real, imag} */,
  {32'hc5836615, 32'h00000000} /* (17, 15, 15) {real, imag} */,
  {32'hc5717eeb, 32'h00000000} /* (17, 15, 14) {real, imag} */,
  {32'hc579e73a, 32'h00000000} /* (17, 15, 13) {real, imag} */,
  {32'hc5658f96, 32'h00000000} /* (17, 15, 12) {real, imag} */,
  {32'hc502c693, 32'h00000000} /* (17, 15, 11) {real, imag} */,
  {32'h4540a126, 32'h00000000} /* (17, 15, 10) {real, imag} */,
  {32'h459fcca5, 32'h00000000} /* (17, 15, 9) {real, imag} */,
  {32'h4590a8ee, 32'h00000000} /* (17, 15, 8) {real, imag} */,
  {32'h457283c6, 32'h00000000} /* (17, 15, 7) {real, imag} */,
  {32'h458b4fd8, 32'h00000000} /* (17, 15, 6) {real, imag} */,
  {32'h458a2df2, 32'h00000000} /* (17, 15, 5) {real, imag} */,
  {32'h459cbcce, 32'h00000000} /* (17, 15, 4) {real, imag} */,
  {32'h45abce7f, 32'h00000000} /* (17, 15, 3) {real, imag} */,
  {32'h45ac38ce, 32'h00000000} /* (17, 15, 2) {real, imag} */,
  {32'h458b5c2a, 32'h00000000} /* (17, 15, 1) {real, imag} */,
  {32'h45832ca6, 32'h00000000} /* (17, 15, 0) {real, imag} */,
  {32'h4550b540, 32'h00000000} /* (17, 14, 31) {real, imag} */,
  {32'h4566622c, 32'h00000000} /* (17, 14, 30) {real, imag} */,
  {32'h45a68535, 32'h00000000} /* (17, 14, 29) {real, imag} */,
  {32'h458eed17, 32'h00000000} /* (17, 14, 28) {real, imag} */,
  {32'h45898e8e, 32'h00000000} /* (17, 14, 27) {real, imag} */,
  {32'h4569dc14, 32'h00000000} /* (17, 14, 26) {real, imag} */,
  {32'h455563c3, 32'h00000000} /* (17, 14, 25) {real, imag} */,
  {32'h453533bc, 32'h00000000} /* (17, 14, 24) {real, imag} */,
  {32'h4532a471, 32'h00000000} /* (17, 14, 23) {real, imag} */,
  {32'h4536918c, 32'h00000000} /* (17, 14, 22) {real, imag} */,
  {32'h448e1358, 32'h00000000} /* (17, 14, 21) {real, imag} */,
  {32'hc488358a, 32'h00000000} /* (17, 14, 20) {real, imag} */,
  {32'hc5866e86, 32'h00000000} /* (17, 14, 19) {real, imag} */,
  {32'hc576cfce, 32'h00000000} /* (17, 14, 18) {real, imag} */,
  {32'hc5510a5a, 32'h00000000} /* (17, 14, 17) {real, imag} */,
  {32'hc577f9a6, 32'h00000000} /* (17, 14, 16) {real, imag} */,
  {32'hc56cb338, 32'h00000000} /* (17, 14, 15) {real, imag} */,
  {32'hc5910818, 32'h00000000} /* (17, 14, 14) {real, imag} */,
  {32'hc54e49de, 32'h00000000} /* (17, 14, 13) {real, imag} */,
  {32'hc531e91f, 32'h00000000} /* (17, 14, 12) {real, imag} */,
  {32'hc321a090, 32'h00000000} /* (17, 14, 11) {real, imag} */,
  {32'h4512ca04, 32'h00000000} /* (17, 14, 10) {real, imag} */,
  {32'h4569b4b1, 32'h00000000} /* (17, 14, 9) {real, imag} */,
  {32'h4568839a, 32'h00000000} /* (17, 14, 8) {real, imag} */,
  {32'h45864233, 32'h00000000} /* (17, 14, 7) {real, imag} */,
  {32'h4577ab38, 32'h00000000} /* (17, 14, 6) {real, imag} */,
  {32'h455507a4, 32'h00000000} /* (17, 14, 5) {real, imag} */,
  {32'h459af650, 32'h00000000} /* (17, 14, 4) {real, imag} */,
  {32'h45a2dac8, 32'h00000000} /* (17, 14, 3) {real, imag} */,
  {32'h45aa52a1, 32'h00000000} /* (17, 14, 2) {real, imag} */,
  {32'h45980831, 32'h00000000} /* (17, 14, 1) {real, imag} */,
  {32'h4566ece8, 32'h00000000} /* (17, 14, 0) {real, imag} */,
  {32'h45349cf9, 32'h00000000} /* (17, 13, 31) {real, imag} */,
  {32'h4542de31, 32'h00000000} /* (17, 13, 30) {real, imag} */,
  {32'h457e5efb, 32'h00000000} /* (17, 13, 29) {real, imag} */,
  {32'h457f0252, 32'h00000000} /* (17, 13, 28) {real, imag} */,
  {32'h453897f7, 32'h00000000} /* (17, 13, 27) {real, imag} */,
  {32'h454b0301, 32'h00000000} /* (17, 13, 26) {real, imag} */,
  {32'h454994ec, 32'h00000000} /* (17, 13, 25) {real, imag} */,
  {32'h451845aa, 32'h00000000} /* (17, 13, 24) {real, imag} */,
  {32'h4505f30b, 32'h00000000} /* (17, 13, 23) {real, imag} */,
  {32'h4527a129, 32'h00000000} /* (17, 13, 22) {real, imag} */,
  {32'h44a81aa6, 32'h00000000} /* (17, 13, 21) {real, imag} */,
  {32'h42bdc100, 32'h00000000} /* (17, 13, 20) {real, imag} */,
  {32'hc522eff3, 32'h00000000} /* (17, 13, 19) {real, imag} */,
  {32'hc54b50ef, 32'h00000000} /* (17, 13, 18) {real, imag} */,
  {32'hc556cd44, 32'h00000000} /* (17, 13, 17) {real, imag} */,
  {32'hc5587f2c, 32'h00000000} /* (17, 13, 16) {real, imag} */,
  {32'hc56451bb, 32'h00000000} /* (17, 13, 15) {real, imag} */,
  {32'hc56aaa3f, 32'h00000000} /* (17, 13, 14) {real, imag} */,
  {32'hc52bae9d, 32'h00000000} /* (17, 13, 13) {real, imag} */,
  {32'hc48c93bb, 32'h00000000} /* (17, 13, 12) {real, imag} */,
  {32'h435ec9f0, 32'h00000000} /* (17, 13, 11) {real, imag} */,
  {32'h451cba49, 32'h00000000} /* (17, 13, 10) {real, imag} */,
  {32'h4571e164, 32'h00000000} /* (17, 13, 9) {real, imag} */,
  {32'h459dba17, 32'h00000000} /* (17, 13, 8) {real, imag} */,
  {32'h4585cfc6, 32'h00000000} /* (17, 13, 7) {real, imag} */,
  {32'h45667111, 32'h00000000} /* (17, 13, 6) {real, imag} */,
  {32'h4562cbc9, 32'h00000000} /* (17, 13, 5) {real, imag} */,
  {32'h458ba4e6, 32'h00000000} /* (17, 13, 4) {real, imag} */,
  {32'h458b3436, 32'h00000000} /* (17, 13, 3) {real, imag} */,
  {32'h4599786a, 32'h00000000} /* (17, 13, 2) {real, imag} */,
  {32'h4568b008, 32'h00000000} /* (17, 13, 1) {real, imag} */,
  {32'h4561afa0, 32'h00000000} /* (17, 13, 0) {real, imag} */,
  {32'h453dd6c2, 32'h00000000} /* (17, 12, 31) {real, imag} */,
  {32'h453b6aed, 32'h00000000} /* (17, 12, 30) {real, imag} */,
  {32'h4538f325, 32'h00000000} /* (17, 12, 29) {real, imag} */,
  {32'h4510491d, 32'h00000000} /* (17, 12, 28) {real, imag} */,
  {32'h44f392b8, 32'h00000000} /* (17, 12, 27) {real, imag} */,
  {32'h4523024b, 32'h00000000} /* (17, 12, 26) {real, imag} */,
  {32'h454366a0, 32'h00000000} /* (17, 12, 25) {real, imag} */,
  {32'h4530a098, 32'h00000000} /* (17, 12, 24) {real, imag} */,
  {32'h44fe0930, 32'h00000000} /* (17, 12, 23) {real, imag} */,
  {32'h454472d0, 32'h00000000} /* (17, 12, 22) {real, imag} */,
  {32'h447e2152, 32'h00000000} /* (17, 12, 21) {real, imag} */,
  {32'hc4812e5b, 32'h00000000} /* (17, 12, 20) {real, imag} */,
  {32'hc5251808, 32'h00000000} /* (17, 12, 19) {real, imag} */,
  {32'hc4f27e01, 32'h00000000} /* (17, 12, 18) {real, imag} */,
  {32'hc510d996, 32'h00000000} /* (17, 12, 17) {real, imag} */,
  {32'hc55a8c8e, 32'h00000000} /* (17, 12, 16) {real, imag} */,
  {32'hc5632886, 32'h00000000} /* (17, 12, 15) {real, imag} */,
  {32'hc52a0b8f, 32'h00000000} /* (17, 12, 14) {real, imag} */,
  {32'hc4a0177a, 32'h00000000} /* (17, 12, 13) {real, imag} */,
  {32'hc4737328, 32'h00000000} /* (17, 12, 12) {real, imag} */,
  {32'h43698970, 32'h00000000} /* (17, 12, 11) {real, imag} */,
  {32'h450b735d, 32'h00000000} /* (17, 12, 10) {real, imag} */,
  {32'h454e85a4, 32'h00000000} /* (17, 12, 9) {real, imag} */,
  {32'h45702840, 32'h00000000} /* (17, 12, 8) {real, imag} */,
  {32'h456f5054, 32'h00000000} /* (17, 12, 7) {real, imag} */,
  {32'h454db800, 32'h00000000} /* (17, 12, 6) {real, imag} */,
  {32'h4544c828, 32'h00000000} /* (17, 12, 5) {real, imag} */,
  {32'h4552ec72, 32'h00000000} /* (17, 12, 4) {real, imag} */,
  {32'h4589aea9, 32'h00000000} /* (17, 12, 3) {real, imag} */,
  {32'h45765012, 32'h00000000} /* (17, 12, 2) {real, imag} */,
  {32'h45578f70, 32'h00000000} /* (17, 12, 1) {real, imag} */,
  {32'h451b530e, 32'h00000000} /* (17, 12, 0) {real, imag} */,
  {32'h4449ef73, 32'h00000000} /* (17, 11, 31) {real, imag} */,
  {32'h44a05162, 32'h00000000} /* (17, 11, 30) {real, imag} */,
  {32'h44e6649f, 32'h00000000} /* (17, 11, 29) {real, imag} */,
  {32'h442d87f4, 32'h00000000} /* (17, 11, 28) {real, imag} */,
  {32'h43b38530, 32'h00000000} /* (17, 11, 27) {real, imag} */,
  {32'h43fdd3d8, 32'h00000000} /* (17, 11, 26) {real, imag} */,
  {32'h44bac2dc, 32'h00000000} /* (17, 11, 25) {real, imag} */,
  {32'h43e45228, 32'h00000000} /* (17, 11, 24) {real, imag} */,
  {32'h44a69146, 32'h00000000} /* (17, 11, 23) {real, imag} */,
  {32'h444ba8c1, 32'h00000000} /* (17, 11, 22) {real, imag} */,
  {32'h44b6f470, 32'h00000000} /* (17, 11, 21) {real, imag} */,
  {32'hc3acd618, 32'h00000000} /* (17, 11, 20) {real, imag} */,
  {32'hc4d53ba4, 32'h00000000} /* (17, 11, 19) {real, imag} */,
  {32'hc4cf2fe2, 32'h00000000} /* (17, 11, 18) {real, imag} */,
  {32'hc491665c, 32'h00000000} /* (17, 11, 17) {real, imag} */,
  {32'hc52105d4, 32'h00000000} /* (17, 11, 16) {real, imag} */,
  {32'hc504e0ee, 32'h00000000} /* (17, 11, 15) {real, imag} */,
  {32'hc35df464, 32'h00000000} /* (17, 11, 14) {real, imag} */,
  {32'hc3f41c84, 32'h00000000} /* (17, 11, 13) {real, imag} */,
  {32'hc4411f90, 32'h00000000} /* (17, 11, 12) {real, imag} */,
  {32'h43353a40, 32'h00000000} /* (17, 11, 11) {real, imag} */,
  {32'h449b4d6d, 32'h00000000} /* (17, 11, 10) {real, imag} */,
  {32'h453395da, 32'h00000000} /* (17, 11, 9) {real, imag} */,
  {32'h452294a7, 32'h00000000} /* (17, 11, 8) {real, imag} */,
  {32'h451071ad, 32'h00000000} /* (17, 11, 7) {real, imag} */,
  {32'h45011186, 32'h00000000} /* (17, 11, 6) {real, imag} */,
  {32'h45570710, 32'h00000000} /* (17, 11, 5) {real, imag} */,
  {32'h45069dd1, 32'h00000000} /* (17, 11, 4) {real, imag} */,
  {32'h45060c57, 32'h00000000} /* (17, 11, 3) {real, imag} */,
  {32'h45102d6d, 32'h00000000} /* (17, 11, 2) {real, imag} */,
  {32'h45354c30, 32'h00000000} /* (17, 11, 1) {real, imag} */,
  {32'h44c58a78, 32'h00000000} /* (17, 11, 0) {real, imag} */,
  {32'hc4b7e36a, 32'h00000000} /* (17, 10, 31) {real, imag} */,
  {32'hc4dffebe, 32'h00000000} /* (17, 10, 30) {real, imag} */,
  {32'hc523f725, 32'h00000000} /* (17, 10, 29) {real, imag} */,
  {32'hc4bc5921, 32'h00000000} /* (17, 10, 28) {real, imag} */,
  {32'hc4dcb44a, 32'h00000000} /* (17, 10, 27) {real, imag} */,
  {32'hc515d941, 32'h00000000} /* (17, 10, 26) {real, imag} */,
  {32'hc4ee62a8, 32'h00000000} /* (17, 10, 25) {real, imag} */,
  {32'hc4a086ee, 32'h00000000} /* (17, 10, 24) {real, imag} */,
  {32'hc450886e, 32'h00000000} /* (17, 10, 23) {real, imag} */,
  {32'hc437bad1, 32'h00000000} /* (17, 10, 22) {real, imag} */,
  {32'hc3f3ac2f, 32'h00000000} /* (17, 10, 21) {real, imag} */,
  {32'h4430da6d, 32'h00000000} /* (17, 10, 20) {real, imag} */,
  {32'hc29c88dc, 32'h00000000} /* (17, 10, 19) {real, imag} */,
  {32'hc2ff1830, 32'h00000000} /* (17, 10, 18) {real, imag} */,
  {32'h4407139b, 32'h00000000} /* (17, 10, 17) {real, imag} */,
  {32'h4459aad6, 32'h00000000} /* (17, 10, 16) {real, imag} */,
  {32'h44e95432, 32'h00000000} /* (17, 10, 15) {real, imag} */,
  {32'h44a3e70a, 32'h00000000} /* (17, 10, 14) {real, imag} */,
  {32'h45042741, 32'h00000000} /* (17, 10, 13) {real, imag} */,
  {32'h451f34e6, 32'h00000000} /* (17, 10, 12) {real, imag} */,
  {32'h44af6256, 32'h00000000} /* (17, 10, 11) {real, imag} */,
  {32'h447ba4db, 32'h00000000} /* (17, 10, 10) {real, imag} */,
  {32'h43d2ea6a, 32'h00000000} /* (17, 10, 9) {real, imag} */,
  {32'h43b80d4b, 32'h00000000} /* (17, 10, 8) {real, imag} */,
  {32'hc230c8e8, 32'h00000000} /* (17, 10, 7) {real, imag} */,
  {32'hc342dcd0, 32'h00000000} /* (17, 10, 6) {real, imag} */,
  {32'h422781e8, 32'h00000000} /* (17, 10, 5) {real, imag} */,
  {32'hc348e0b8, 32'h00000000} /* (17, 10, 4) {real, imag} */,
  {32'hc3c5b4df, 32'h00000000} /* (17, 10, 3) {real, imag} */,
  {32'hc4f57e09, 32'h00000000} /* (17, 10, 2) {real, imag} */,
  {32'hc41df249, 32'h00000000} /* (17, 10, 1) {real, imag} */,
  {32'hc4b1edd9, 32'h00000000} /* (17, 10, 0) {real, imag} */,
  {32'hc5502a65, 32'h00000000} /* (17, 9, 31) {real, imag} */,
  {32'hc577c95c, 32'h00000000} /* (17, 9, 30) {real, imag} */,
  {32'hc54ce1f4, 32'h00000000} /* (17, 9, 29) {real, imag} */,
  {32'hc55cc421, 32'h00000000} /* (17, 9, 28) {real, imag} */,
  {32'hc576ac2f, 32'h00000000} /* (17, 9, 27) {real, imag} */,
  {32'hc56ebd01, 32'h00000000} /* (17, 9, 26) {real, imag} */,
  {32'hc5340252, 32'h00000000} /* (17, 9, 25) {real, imag} */,
  {32'hc5401837, 32'h00000000} /* (17, 9, 24) {real, imag} */,
  {32'hc4e7eb0a, 32'h00000000} /* (17, 9, 23) {real, imag} */,
  {32'hc52d8850, 32'h00000000} /* (17, 9, 22) {real, imag} */,
  {32'hc5004a10, 32'h00000000} /* (17, 9, 21) {real, imag} */,
  {32'h442b1153, 32'h00000000} /* (17, 9, 20) {real, imag} */,
  {32'h4486445a, 32'h00000000} /* (17, 9, 19) {real, imag} */,
  {32'h44d1e212, 32'h00000000} /* (17, 9, 18) {real, imag} */,
  {32'h45264ef3, 32'h00000000} /* (17, 9, 17) {real, imag} */,
  {32'h454873fc, 32'h00000000} /* (17, 9, 16) {real, imag} */,
  {32'h4578058b, 32'h00000000} /* (17, 9, 15) {real, imag} */,
  {32'h456f7f50, 32'h00000000} /* (17, 9, 14) {real, imag} */,
  {32'h45429f36, 32'h00000000} /* (17, 9, 13) {real, imag} */,
  {32'h450cc73d, 32'h00000000} /* (17, 9, 12) {real, imag} */,
  {32'h44c33d32, 32'h00000000} /* (17, 9, 11) {real, imag} */,
  {32'h439f2158, 32'h00000000} /* (17, 9, 10) {real, imag} */,
  {32'hc40707e4, 32'h00000000} /* (17, 9, 9) {real, imag} */,
  {32'hc438c7fc, 32'h00000000} /* (17, 9, 8) {real, imag} */,
  {32'hc4da1186, 32'h00000000} /* (17, 9, 7) {real, imag} */,
  {32'hc4c32554, 32'h00000000} /* (17, 9, 6) {real, imag} */,
  {32'hc532e594, 32'h00000000} /* (17, 9, 5) {real, imag} */,
  {32'hc50feded, 32'h00000000} /* (17, 9, 4) {real, imag} */,
  {32'hc50ac536, 32'h00000000} /* (17, 9, 3) {real, imag} */,
  {32'hc51410a1, 32'h00000000} /* (17, 9, 2) {real, imag} */,
  {32'hc54a9b1d, 32'h00000000} /* (17, 9, 1) {real, imag} */,
  {32'hc5459b5c, 32'h00000000} /* (17, 9, 0) {real, imag} */,
  {32'hc599a797, 32'h00000000} /* (17, 8, 31) {real, imag} */,
  {32'hc5a19d95, 32'h00000000} /* (17, 8, 30) {real, imag} */,
  {32'hc585cf52, 32'h00000000} /* (17, 8, 29) {real, imag} */,
  {32'hc5a110b3, 32'h00000000} /* (17, 8, 28) {real, imag} */,
  {32'hc5a67600, 32'h00000000} /* (17, 8, 27) {real, imag} */,
  {32'hc5a38130, 32'h00000000} /* (17, 8, 26) {real, imag} */,
  {32'hc591d58d, 32'h00000000} /* (17, 8, 25) {real, imag} */,
  {32'hc56ac091, 32'h00000000} /* (17, 8, 24) {real, imag} */,
  {32'hc56c1d03, 32'h00000000} /* (17, 8, 23) {real, imag} */,
  {32'hc536c798, 32'h00000000} /* (17, 8, 22) {real, imag} */,
  {32'hc4dd9f5f, 32'h00000000} /* (17, 8, 21) {real, imag} */,
  {32'hc40ca788, 32'h00000000} /* (17, 8, 20) {real, imag} */,
  {32'h4478e586, 32'h00000000} /* (17, 8, 19) {real, imag} */,
  {32'h44e79ecc, 32'h00000000} /* (17, 8, 18) {real, imag} */,
  {32'h451dd6ea, 32'h00000000} /* (17, 8, 17) {real, imag} */,
  {32'h45a5792c, 32'h00000000} /* (17, 8, 16) {real, imag} */,
  {32'h45875199, 32'h00000000} /* (17, 8, 15) {real, imag} */,
  {32'h457b3ee6, 32'h00000000} /* (17, 8, 14) {real, imag} */,
  {32'h456e1177, 32'h00000000} /* (17, 8, 13) {real, imag} */,
  {32'h456fd592, 32'h00000000} /* (17, 8, 12) {real, imag} */,
  {32'h44a6fb0b, 32'h00000000} /* (17, 8, 11) {real, imag} */,
  {32'h42b90da0, 32'h00000000} /* (17, 8, 10) {real, imag} */,
  {32'hc484f544, 32'h00000000} /* (17, 8, 9) {real, imag} */,
  {32'hc4ee7a06, 32'h00000000} /* (17, 8, 8) {real, imag} */,
  {32'hc4cffab2, 32'h00000000} /* (17, 8, 7) {real, imag} */,
  {32'hc4fd3619, 32'h00000000} /* (17, 8, 6) {real, imag} */,
  {32'hc5839f5d, 32'h00000000} /* (17, 8, 5) {real, imag} */,
  {32'hc59026c8, 32'h00000000} /* (17, 8, 4) {real, imag} */,
  {32'hc55c5f9a, 32'h00000000} /* (17, 8, 3) {real, imag} */,
  {32'hc5873933, 32'h00000000} /* (17, 8, 2) {real, imag} */,
  {32'hc58bd0b4, 32'h00000000} /* (17, 8, 1) {real, imag} */,
  {32'hc5879c62, 32'h00000000} /* (17, 8, 0) {real, imag} */,
  {32'hc5c1e04a, 32'h00000000} /* (17, 7, 31) {real, imag} */,
  {32'hc5ce169c, 32'h00000000} /* (17, 7, 30) {real, imag} */,
  {32'hc5c7516c, 32'h00000000} /* (17, 7, 29) {real, imag} */,
  {32'hc5ac2bb8, 32'h00000000} /* (17, 7, 28) {real, imag} */,
  {32'hc5b85e46, 32'h00000000} /* (17, 7, 27) {real, imag} */,
  {32'hc5bc7ce6, 32'h00000000} /* (17, 7, 26) {real, imag} */,
  {32'hc5a91364, 32'h00000000} /* (17, 7, 25) {real, imag} */,
  {32'hc593b334, 32'h00000000} /* (17, 7, 24) {real, imag} */,
  {32'hc5ba7af9, 32'h00000000} /* (17, 7, 23) {real, imag} */,
  {32'hc5753d1e, 32'h00000000} /* (17, 7, 22) {real, imag} */,
  {32'hc52c0fbe, 32'h00000000} /* (17, 7, 21) {real, imag} */,
  {32'hc49909d5, 32'h00000000} /* (17, 7, 20) {real, imag} */,
  {32'h442d9cd0, 32'h00000000} /* (17, 7, 19) {real, imag} */,
  {32'h4531103a, 32'h00000000} /* (17, 7, 18) {real, imag} */,
  {32'h453b89cc, 32'h00000000} /* (17, 7, 17) {real, imag} */,
  {32'h455a92ec, 32'h00000000} /* (17, 7, 16) {real, imag} */,
  {32'h455ff1d1, 32'h00000000} /* (17, 7, 15) {real, imag} */,
  {32'h45815d4c, 32'h00000000} /* (17, 7, 14) {real, imag} */,
  {32'h457e4bc5, 32'h00000000} /* (17, 7, 13) {real, imag} */,
  {32'h45940482, 32'h00000000} /* (17, 7, 12) {real, imag} */,
  {32'h454a8851, 32'h00000000} /* (17, 7, 11) {real, imag} */,
  {32'h43351080, 32'h00000000} /* (17, 7, 10) {real, imag} */,
  {32'hc49e2350, 32'h00000000} /* (17, 7, 9) {real, imag} */,
  {32'hc4f8e656, 32'h00000000} /* (17, 7, 8) {real, imag} */,
  {32'hc4df7178, 32'h00000000} /* (17, 7, 7) {real, imag} */,
  {32'hc559f928, 32'h00000000} /* (17, 7, 6) {real, imag} */,
  {32'hc581f6de, 32'h00000000} /* (17, 7, 5) {real, imag} */,
  {32'hc58f19c4, 32'h00000000} /* (17, 7, 4) {real, imag} */,
  {32'hc5a2bb19, 32'h00000000} /* (17, 7, 3) {real, imag} */,
  {32'hc5a40a4c, 32'h00000000} /* (17, 7, 2) {real, imag} */,
  {32'hc5a554ac, 32'h00000000} /* (17, 7, 1) {real, imag} */,
  {32'hc5930442, 32'h00000000} /* (17, 7, 0) {real, imag} */,
  {32'hc5b6f08d, 32'h00000000} /* (17, 6, 31) {real, imag} */,
  {32'hc5e096ae, 32'h00000000} /* (17, 6, 30) {real, imag} */,
  {32'hc5df76dc, 32'h00000000} /* (17, 6, 29) {real, imag} */,
  {32'hc5c70023, 32'h00000000} /* (17, 6, 28) {real, imag} */,
  {32'hc5b31b72, 32'h00000000} /* (17, 6, 27) {real, imag} */,
  {32'hc5b835fa, 32'h00000000} /* (17, 6, 26) {real, imag} */,
  {32'hc5c9e14e, 32'h00000000} /* (17, 6, 25) {real, imag} */,
  {32'hc5d6db82, 32'h00000000} /* (17, 6, 24) {real, imag} */,
  {32'hc5a3b3d6, 32'h00000000} /* (17, 6, 23) {real, imag} */,
  {32'hc58fddfc, 32'h00000000} /* (17, 6, 22) {real, imag} */,
  {32'hc581a83e, 32'h00000000} /* (17, 6, 21) {real, imag} */,
  {32'hc44526d4, 32'h00000000} /* (17, 6, 20) {real, imag} */,
  {32'h43ab9bf0, 32'h00000000} /* (17, 6, 19) {real, imag} */,
  {32'h449c2bfe, 32'h00000000} /* (17, 6, 18) {real, imag} */,
  {32'h4518cf66, 32'h00000000} /* (17, 6, 17) {real, imag} */,
  {32'h45531b92, 32'h00000000} /* (17, 6, 16) {real, imag} */,
  {32'h457dea56, 32'h00000000} /* (17, 6, 15) {real, imag} */,
  {32'h4585452c, 32'h00000000} /* (17, 6, 14) {real, imag} */,
  {32'h45830cba, 32'h00000000} /* (17, 6, 13) {real, imag} */,
  {32'h45812075, 32'h00000000} /* (17, 6, 12) {real, imag} */,
  {32'h45482591, 32'h00000000} /* (17, 6, 11) {real, imag} */,
  {32'h4496ec78, 32'h00000000} /* (17, 6, 10) {real, imag} */,
  {32'hc4cbfdde, 32'h00000000} /* (17, 6, 9) {real, imag} */,
  {32'hc479e0e0, 32'h00000000} /* (17, 6, 8) {real, imag} */,
  {32'hc4baf752, 32'h00000000} /* (17, 6, 7) {real, imag} */,
  {32'hc5406758, 32'h00000000} /* (17, 6, 6) {real, imag} */,
  {32'hc54bffc6, 32'h00000000} /* (17, 6, 5) {real, imag} */,
  {32'hc5a36460, 32'h00000000} /* (17, 6, 4) {real, imag} */,
  {32'hc5acc01e, 32'h00000000} /* (17, 6, 3) {real, imag} */,
  {32'hc5ab11f2, 32'h00000000} /* (17, 6, 2) {real, imag} */,
  {32'hc5b3c09d, 32'h00000000} /* (17, 6, 1) {real, imag} */,
  {32'hc5a51243, 32'h00000000} /* (17, 6, 0) {real, imag} */,
  {32'hc5bf39f9, 32'h00000000} /* (17, 5, 31) {real, imag} */,
  {32'hc5d1dd38, 32'h00000000} /* (17, 5, 30) {real, imag} */,
  {32'hc5eb0662, 32'h00000000} /* (17, 5, 29) {real, imag} */,
  {32'hc5d4d2fa, 32'h00000000} /* (17, 5, 28) {real, imag} */,
  {32'hc5c287cc, 32'h00000000} /* (17, 5, 27) {real, imag} */,
  {32'hc5ab32fc, 32'h00000000} /* (17, 5, 26) {real, imag} */,
  {32'hc5d4d73f, 32'h00000000} /* (17, 5, 25) {real, imag} */,
  {32'hc5c4ae23, 32'h00000000} /* (17, 5, 24) {real, imag} */,
  {32'hc598d3fe, 32'h00000000} /* (17, 5, 23) {real, imag} */,
  {32'hc5a12fe2, 32'h00000000} /* (17, 5, 22) {real, imag} */,
  {32'hc59a443c, 32'h00000000} /* (17, 5, 21) {real, imag} */,
  {32'hc56a0656, 32'h00000000} /* (17, 5, 20) {real, imag} */,
  {32'hc51d5b46, 32'h00000000} /* (17, 5, 19) {real, imag} */,
  {32'hc44020c0, 32'h00000000} /* (17, 5, 18) {real, imag} */,
  {32'h447702ec, 32'h00000000} /* (17, 5, 17) {real, imag} */,
  {32'h44cd7692, 32'h00000000} /* (17, 5, 16) {real, imag} */,
  {32'h453c12fa, 32'h00000000} /* (17, 5, 15) {real, imag} */,
  {32'h457706ff, 32'h00000000} /* (17, 5, 14) {real, imag} */,
  {32'h457e7b8b, 32'h00000000} /* (17, 5, 13) {real, imag} */,
  {32'h4558bc97, 32'h00000000} /* (17, 5, 12) {real, imag} */,
  {32'h45734f31, 32'h00000000} /* (17, 5, 11) {real, imag} */,
  {32'h451d44b3, 32'h00000000} /* (17, 5, 10) {real, imag} */,
  {32'h44ab07bc, 32'h00000000} /* (17, 5, 9) {real, imag} */,
  {32'h44745208, 32'h00000000} /* (17, 5, 8) {real, imag} */,
  {32'h40f7ce00, 32'h00000000} /* (17, 5, 7) {real, imag} */,
  {32'hc4b10195, 32'h00000000} /* (17, 5, 6) {real, imag} */,
  {32'hc5526be1, 32'h00000000} /* (17, 5, 5) {real, imag} */,
  {32'hc5a07fa9, 32'h00000000} /* (17, 5, 4) {real, imag} */,
  {32'hc59d064c, 32'h00000000} /* (17, 5, 3) {real, imag} */,
  {32'hc5ba0bb2, 32'h00000000} /* (17, 5, 2) {real, imag} */,
  {32'hc5aa7b54, 32'h00000000} /* (17, 5, 1) {real, imag} */,
  {32'hc5b4d5dc, 32'h00000000} /* (17, 5, 0) {real, imag} */,
  {32'hc5baba9c, 32'h00000000} /* (17, 4, 31) {real, imag} */,
  {32'hc5dad458, 32'h00000000} /* (17, 4, 30) {real, imag} */,
  {32'hc5e116a2, 32'h00000000} /* (17, 4, 29) {real, imag} */,
  {32'hc5d184da, 32'h00000000} /* (17, 4, 28) {real, imag} */,
  {32'hc5c3df05, 32'h00000000} /* (17, 4, 27) {real, imag} */,
  {32'hc5b470de, 32'h00000000} /* (17, 4, 26) {real, imag} */,
  {32'hc5b4f872, 32'h00000000} /* (17, 4, 25) {real, imag} */,
  {32'hc5a704fd, 32'h00000000} /* (17, 4, 24) {real, imag} */,
  {32'hc5b89bd4, 32'h00000000} /* (17, 4, 23) {real, imag} */,
  {32'hc5a56e28, 32'h00000000} /* (17, 4, 22) {real, imag} */,
  {32'hc5a423aa, 32'h00000000} /* (17, 4, 21) {real, imag} */,
  {32'hc58fbc6c, 32'h00000000} /* (17, 4, 20) {real, imag} */,
  {32'hc54e2e02, 32'h00000000} /* (17, 4, 19) {real, imag} */,
  {32'hc4cf5830, 32'h00000000} /* (17, 4, 18) {real, imag} */,
  {32'hc5047eeb, 32'h00000000} /* (17, 4, 17) {real, imag} */,
  {32'h43cb3d28, 32'h00000000} /* (17, 4, 16) {real, imag} */,
  {32'h4512eceb, 32'h00000000} /* (17, 4, 15) {real, imag} */,
  {32'h45862154, 32'h00000000} /* (17, 4, 14) {real, imag} */,
  {32'h4581d6dc, 32'h00000000} /* (17, 4, 13) {real, imag} */,
  {32'h455e81dc, 32'h00000000} /* (17, 4, 12) {real, imag} */,
  {32'h45807199, 32'h00000000} /* (17, 4, 11) {real, imag} */,
  {32'h455a95a5, 32'h00000000} /* (17, 4, 10) {real, imag} */,
  {32'h455180c1, 32'h00000000} /* (17, 4, 9) {real, imag} */,
  {32'h455fd0bd, 32'h00000000} /* (17, 4, 8) {real, imag} */,
  {32'h44e7da5c, 32'h00000000} /* (17, 4, 7) {real, imag} */,
  {32'hc3b54e00, 32'h00000000} /* (17, 4, 6) {real, imag} */,
  {32'hc5248db2, 32'h00000000} /* (17, 4, 5) {real, imag} */,
  {32'hc5a85de6, 32'h00000000} /* (17, 4, 4) {real, imag} */,
  {32'hc5989c8f, 32'h00000000} /* (17, 4, 3) {real, imag} */,
  {32'hc59eae51, 32'h00000000} /* (17, 4, 2) {real, imag} */,
  {32'hc5ae8188, 32'h00000000} /* (17, 4, 1) {real, imag} */,
  {32'hc5af57aa, 32'h00000000} /* (17, 4, 0) {real, imag} */,
  {32'hc5a96b96, 32'h00000000} /* (17, 3, 31) {real, imag} */,
  {32'hc5f57a56, 32'h00000000} /* (17, 3, 30) {real, imag} */,
  {32'hc5f00516, 32'h00000000} /* (17, 3, 29) {real, imag} */,
  {32'hc5c87a7c, 32'h00000000} /* (17, 3, 28) {real, imag} */,
  {32'hc5d49e49, 32'h00000000} /* (17, 3, 27) {real, imag} */,
  {32'hc5c1f187, 32'h00000000} /* (17, 3, 26) {real, imag} */,
  {32'hc5becf1e, 32'h00000000} /* (17, 3, 25) {real, imag} */,
  {32'hc5c0264c, 32'h00000000} /* (17, 3, 24) {real, imag} */,
  {32'hc5b2dfec, 32'h00000000} /* (17, 3, 23) {real, imag} */,
  {32'hc5b057be, 32'h00000000} /* (17, 3, 22) {real, imag} */,
  {32'hc5a3fe1e, 32'h00000000} /* (17, 3, 21) {real, imag} */,
  {32'hc5898c8d, 32'h00000000} /* (17, 3, 20) {real, imag} */,
  {32'hc576820f, 32'h00000000} /* (17, 3, 19) {real, imag} */,
  {32'hc59908b6, 32'h00000000} /* (17, 3, 18) {real, imag} */,
  {32'hc50315ef, 32'h00000000} /* (17, 3, 17) {real, imag} */,
  {32'hc018ac00, 32'h00000000} /* (17, 3, 16) {real, imag} */,
  {32'h45639667, 32'h00000000} /* (17, 3, 15) {real, imag} */,
  {32'h4591462e, 32'h00000000} /* (17, 3, 14) {real, imag} */,
  {32'h45a10392, 32'h00000000} /* (17, 3, 13) {real, imag} */,
  {32'h459c878a, 32'h00000000} /* (17, 3, 12) {real, imag} */,
  {32'h45abf28f, 32'h00000000} /* (17, 3, 11) {real, imag} */,
  {32'h45907099, 32'h00000000} /* (17, 3, 10) {real, imag} */,
  {32'h457e65d5, 32'h00000000} /* (17, 3, 9) {real, imag} */,
  {32'h457a4098, 32'h00000000} /* (17, 3, 8) {real, imag} */,
  {32'h44b354a2, 32'h00000000} /* (17, 3, 7) {real, imag} */,
  {32'hc3463a90, 32'h00000000} /* (17, 3, 6) {real, imag} */,
  {32'hc535412d, 32'h00000000} /* (17, 3, 5) {real, imag} */,
  {32'hc596e94d, 32'h00000000} /* (17, 3, 4) {real, imag} */,
  {32'hc5999716, 32'h00000000} /* (17, 3, 3) {real, imag} */,
  {32'hc59ff4ec, 32'h00000000} /* (17, 3, 2) {real, imag} */,
  {32'hc5ac5fba, 32'h00000000} /* (17, 3, 1) {real, imag} */,
  {32'hc5ad7f58, 32'h00000000} /* (17, 3, 0) {real, imag} */,
  {32'hc5b01f7a, 32'h00000000} /* (17, 2, 31) {real, imag} */,
  {32'hc5cba343, 32'h00000000} /* (17, 2, 30) {real, imag} */,
  {32'hc5dbaee1, 32'h00000000} /* (17, 2, 29) {real, imag} */,
  {32'hc5c07622, 32'h00000000} /* (17, 2, 28) {real, imag} */,
  {32'hc5c61c18, 32'h00000000} /* (17, 2, 27) {real, imag} */,
  {32'hc5e2ecd1, 32'h00000000} /* (17, 2, 26) {real, imag} */,
  {32'hc5c2ffe6, 32'h00000000} /* (17, 2, 25) {real, imag} */,
  {32'hc5b3bb6c, 32'h00000000} /* (17, 2, 24) {real, imag} */,
  {32'hc5a701f4, 32'h00000000} /* (17, 2, 23) {real, imag} */,
  {32'hc59c1a4f, 32'h00000000} /* (17, 2, 22) {real, imag} */,
  {32'hc59034d8, 32'h00000000} /* (17, 2, 21) {real, imag} */,
  {32'hc57a163e, 32'h00000000} /* (17, 2, 20) {real, imag} */,
  {32'hc578ec8d, 32'h00000000} /* (17, 2, 19) {real, imag} */,
  {32'hc5c22af2, 32'h00000000} /* (17, 2, 18) {real, imag} */,
  {32'hc5600a53, 32'h00000000} /* (17, 2, 17) {real, imag} */,
  {32'h432acb20, 32'h00000000} /* (17, 2, 16) {real, imag} */,
  {32'h45386eb1, 32'h00000000} /* (17, 2, 15) {real, imag} */,
  {32'h457f5cc2, 32'h00000000} /* (17, 2, 14) {real, imag} */,
  {32'h45aecfcb, 32'h00000000} /* (17, 2, 13) {real, imag} */,
  {32'h458b5e2e, 32'h00000000} /* (17, 2, 12) {real, imag} */,
  {32'h45b2f674, 32'h00000000} /* (17, 2, 11) {real, imag} */,
  {32'h45768d3a, 32'h00000000} /* (17, 2, 10) {real, imag} */,
  {32'h4540b1e4, 32'h00000000} /* (17, 2, 9) {real, imag} */,
  {32'h451f2ad4, 32'h00000000} /* (17, 2, 8) {real, imag} */,
  {32'h44828a94, 32'h00000000} /* (17, 2, 7) {real, imag} */,
  {32'hc3bf08b0, 32'h00000000} /* (17, 2, 6) {real, imag} */,
  {32'hc526db19, 32'h00000000} /* (17, 2, 5) {real, imag} */,
  {32'hc58d6139, 32'h00000000} /* (17, 2, 4) {real, imag} */,
  {32'hc59854be, 32'h00000000} /* (17, 2, 3) {real, imag} */,
  {32'hc5ae432a, 32'h00000000} /* (17, 2, 2) {real, imag} */,
  {32'hc5b8a928, 32'h00000000} /* (17, 2, 1) {real, imag} */,
  {32'hc5b12097, 32'h00000000} /* (17, 2, 0) {real, imag} */,
  {32'hc5b47070, 32'h00000000} /* (17, 1, 31) {real, imag} */,
  {32'hc5c15e5e, 32'h00000000} /* (17, 1, 30) {real, imag} */,
  {32'hc5d691ef, 32'h00000000} /* (17, 1, 29) {real, imag} */,
  {32'hc5c74d56, 32'h00000000} /* (17, 1, 28) {real, imag} */,
  {32'hc5d1a4bc, 32'h00000000} /* (17, 1, 27) {real, imag} */,
  {32'hc5d65eda, 32'h00000000} /* (17, 1, 26) {real, imag} */,
  {32'hc5d40025, 32'h00000000} /* (17, 1, 25) {real, imag} */,
  {32'hc5ae5a01, 32'h00000000} /* (17, 1, 24) {real, imag} */,
  {32'hc5b300ea, 32'h00000000} /* (17, 1, 23) {real, imag} */,
  {32'hc5a8eb9c, 32'h00000000} /* (17, 1, 22) {real, imag} */,
  {32'hc58458da, 32'h00000000} /* (17, 1, 21) {real, imag} */,
  {32'hc58aebec, 32'h00000000} /* (17, 1, 20) {real, imag} */,
  {32'hc57a32a4, 32'h00000000} /* (17, 1, 19) {real, imag} */,
  {32'hc59c9c52, 32'h00000000} /* (17, 1, 18) {real, imag} */,
  {32'hc544e142, 32'h00000000} /* (17, 1, 17) {real, imag} */,
  {32'hc39b67e0, 32'h00000000} /* (17, 1, 16) {real, imag} */,
  {32'h452077f0, 32'h00000000} /* (17, 1, 15) {real, imag} */,
  {32'h459a7506, 32'h00000000} /* (17, 1, 14) {real, imag} */,
  {32'h4593255b, 32'h00000000} /* (17, 1, 13) {real, imag} */,
  {32'h458ba89e, 32'h00000000} /* (17, 1, 12) {real, imag} */,
  {32'h45729790, 32'h00000000} /* (17, 1, 11) {real, imag} */,
  {32'h4547a441, 32'h00000000} /* (17, 1, 10) {real, imag} */,
  {32'h45004d2e, 32'h00000000} /* (17, 1, 9) {real, imag} */,
  {32'h44e54384, 32'h00000000} /* (17, 1, 8) {real, imag} */,
  {32'h44134cf0, 32'h00000000} /* (17, 1, 7) {real, imag} */,
  {32'hc447ade0, 32'h00000000} /* (17, 1, 6) {real, imag} */,
  {32'hc54c8d4b, 32'h00000000} /* (17, 1, 5) {real, imag} */,
  {32'hc59f7546, 32'h00000000} /* (17, 1, 4) {real, imag} */,
  {32'hc5923052, 32'h00000000} /* (17, 1, 3) {real, imag} */,
  {32'hc5adda72, 32'h00000000} /* (17, 1, 2) {real, imag} */,
  {32'hc5c27081, 32'h00000000} /* (17, 1, 1) {real, imag} */,
  {32'hc5adba2c, 32'h00000000} /* (17, 1, 0) {real, imag} */,
  {32'hc5c0a854, 32'h00000000} /* (17, 0, 31) {real, imag} */,
  {32'hc5ba0034, 32'h00000000} /* (17, 0, 30) {real, imag} */,
  {32'hc5cc3603, 32'h00000000} /* (17, 0, 29) {real, imag} */,
  {32'hc5c81a40, 32'h00000000} /* (17, 0, 28) {real, imag} */,
  {32'hc5c8338a, 32'h00000000} /* (17, 0, 27) {real, imag} */,
  {32'hc5cad03b, 32'h00000000} /* (17, 0, 26) {real, imag} */,
  {32'hc5b69b3b, 32'h00000000} /* (17, 0, 25) {real, imag} */,
  {32'hc5a5d0a8, 32'h00000000} /* (17, 0, 24) {real, imag} */,
  {32'hc5a6f2d4, 32'h00000000} /* (17, 0, 23) {real, imag} */,
  {32'hc59a476e, 32'h00000000} /* (17, 0, 22) {real, imag} */,
  {32'hc57c36b3, 32'h00000000} /* (17, 0, 21) {real, imag} */,
  {32'hc55a59a0, 32'h00000000} /* (17, 0, 20) {real, imag} */,
  {32'hc5236220, 32'h00000000} /* (17, 0, 19) {real, imag} */,
  {32'hc4e2d3a8, 32'h00000000} /* (17, 0, 18) {real, imag} */,
  {32'hc43d7974, 32'h00000000} /* (17, 0, 17) {real, imag} */,
  {32'h44880504, 32'h00000000} /* (17, 0, 16) {real, imag} */,
  {32'h450b3bdb, 32'h00000000} /* (17, 0, 15) {real, imag} */,
  {32'h4557a514, 32'h00000000} /* (17, 0, 14) {real, imag} */,
  {32'h4563a206, 32'h00000000} /* (17, 0, 13) {real, imag} */,
  {32'h456d52bc, 32'h00000000} /* (17, 0, 12) {real, imag} */,
  {32'h4560613f, 32'h00000000} /* (17, 0, 11) {real, imag} */,
  {32'h451332c2, 32'h00000000} /* (17, 0, 10) {real, imag} */,
  {32'h447acfa8, 32'h00000000} /* (17, 0, 9) {real, imag} */,
  {32'h439f1ca0, 32'h00000000} /* (17, 0, 8) {real, imag} */,
  {32'hc4440adc, 32'h00000000} /* (17, 0, 7) {real, imag} */,
  {32'hc4e0a352, 32'h00000000} /* (17, 0, 6) {real, imag} */,
  {32'hc53711f5, 32'h00000000} /* (17, 0, 5) {real, imag} */,
  {32'hc584280c, 32'h00000000} /* (17, 0, 4) {real, imag} */,
  {32'hc59a6153, 32'h00000000} /* (17, 0, 3) {real, imag} */,
  {32'hc5b23f98, 32'h00000000} /* (17, 0, 2) {real, imag} */,
  {32'hc5a3d114, 32'h00000000} /* (17, 0, 1) {real, imag} */,
  {32'hc5adca1d, 32'h00000000} /* (17, 0, 0) {real, imag} */,
  {32'hc51848bb, 32'h00000000} /* (16, 31, 31) {real, imag} */,
  {32'hc5264072, 32'h00000000} /* (16, 31, 30) {real, imag} */,
  {32'hc51abc39, 32'h00000000} /* (16, 31, 29) {real, imag} */,
  {32'hc51fd146, 32'h00000000} /* (16, 31, 28) {real, imag} */,
  {32'hc5120795, 32'h00000000} /* (16, 31, 27) {real, imag} */,
  {32'hc4d771e2, 32'h00000000} /* (16, 31, 26) {real, imag} */,
  {32'hc4ff082e, 32'h00000000} /* (16, 31, 25) {real, imag} */,
  {32'hc4f0750c, 32'h00000000} /* (16, 31, 24) {real, imag} */,
  {32'hc5144f67, 32'h00000000} /* (16, 31, 23) {real, imag} */,
  {32'hc4fce94a, 32'h00000000} /* (16, 31, 22) {real, imag} */,
  {32'hc462765a, 32'h00000000} /* (16, 31, 21) {real, imag} */,
  {32'hc44446da, 32'h00000000} /* (16, 31, 20) {real, imag} */,
  {32'hc3bea488, 32'h00000000} /* (16, 31, 19) {real, imag} */,
  {32'h42234860, 32'h00000000} /* (16, 31, 18) {real, imag} */,
  {32'h42c20fa0, 32'h00000000} /* (16, 31, 17) {real, imag} */,
  {32'h444f77c6, 32'h00000000} /* (16, 31, 16) {real, imag} */,
  {32'h43a62808, 32'h00000000} /* (16, 31, 15) {real, imag} */,
  {32'h44b07017, 32'h00000000} /* (16, 31, 14) {real, imag} */,
  {32'h44b0e6f6, 32'h00000000} /* (16, 31, 13) {real, imag} */,
  {32'h44c423ac, 32'h00000000} /* (16, 31, 12) {real, imag} */,
  {32'h44759163, 32'h00000000} /* (16, 31, 11) {real, imag} */,
  {32'hc23339d0, 32'h00000000} /* (16, 31, 10) {real, imag} */,
  {32'hc34e1d60, 32'h00000000} /* (16, 31, 9) {real, imag} */,
  {32'hc4c3d0f0, 32'h00000000} /* (16, 31, 8) {real, imag} */,
  {32'hc4e32bde, 32'h00000000} /* (16, 31, 7) {real, imag} */,
  {32'hc4b71310, 32'h00000000} /* (16, 31, 6) {real, imag} */,
  {32'hc5158f26, 32'h00000000} /* (16, 31, 5) {real, imag} */,
  {32'hc4e285b3, 32'h00000000} /* (16, 31, 4) {real, imag} */,
  {32'hc53943e7, 32'h00000000} /* (16, 31, 3) {real, imag} */,
  {32'hc502c0b2, 32'h00000000} /* (16, 31, 2) {real, imag} */,
  {32'hc50e8512, 32'h00000000} /* (16, 31, 1) {real, imag} */,
  {32'hc50bd258, 32'h00000000} /* (16, 31, 0) {real, imag} */,
  {32'hc509bb1f, 32'h00000000} /* (16, 30, 31) {real, imag} */,
  {32'hc538bbbd, 32'h00000000} /* (16, 30, 30) {real, imag} */,
  {32'hc561dc32, 32'h00000000} /* (16, 30, 29) {real, imag} */,
  {32'hc54888fc, 32'h00000000} /* (16, 30, 28) {real, imag} */,
  {32'hc54fb773, 32'h00000000} /* (16, 30, 27) {real, imag} */,
  {32'hc5052864, 32'h00000000} /* (16, 30, 26) {real, imag} */,
  {32'hc4dc0ec7, 32'h00000000} /* (16, 30, 25) {real, imag} */,
  {32'hc4d08c56, 32'h00000000} /* (16, 30, 24) {real, imag} */,
  {32'hc4e421bd, 32'h00000000} /* (16, 30, 23) {real, imag} */,
  {32'hc4e26ea2, 32'h00000000} /* (16, 30, 22) {real, imag} */,
  {32'hc3fc59d0, 32'h00000000} /* (16, 30, 21) {real, imag} */,
  {32'h43c0dcb8, 32'h00000000} /* (16, 30, 20) {real, imag} */,
  {32'h448497ca, 32'h00000000} /* (16, 30, 19) {real, imag} */,
  {32'h446b0a74, 32'h00000000} /* (16, 30, 18) {real, imag} */,
  {32'h4485a32a, 32'h00000000} /* (16, 30, 17) {real, imag} */,
  {32'h4493431e, 32'h00000000} /* (16, 30, 16) {real, imag} */,
  {32'h4503525d, 32'h00000000} /* (16, 30, 15) {real, imag} */,
  {32'h45034e69, 32'h00000000} /* (16, 30, 14) {real, imag} */,
  {32'h44c448cb, 32'h00000000} /* (16, 30, 13) {real, imag} */,
  {32'h44ce41c3, 32'h00000000} /* (16, 30, 12) {real, imag} */,
  {32'h4489829e, 32'h00000000} /* (16, 30, 11) {real, imag} */,
  {32'h438c284e, 32'h00000000} /* (16, 30, 10) {real, imag} */,
  {32'hc4b7bb41, 32'h00000000} /* (16, 30, 9) {real, imag} */,
  {32'hc50c568a, 32'h00000000} /* (16, 30, 8) {real, imag} */,
  {32'hc53b1ef4, 32'h00000000} /* (16, 30, 7) {real, imag} */,
  {32'hc4e1ac6a, 32'h00000000} /* (16, 30, 6) {real, imag} */,
  {32'hc5095909, 32'h00000000} /* (16, 30, 5) {real, imag} */,
  {32'hc5576f4e, 32'h00000000} /* (16, 30, 4) {real, imag} */,
  {32'hc53c1a79, 32'h00000000} /* (16, 30, 3) {real, imag} */,
  {32'hc55e9cc1, 32'h00000000} /* (16, 30, 2) {real, imag} */,
  {32'hc50b516e, 32'h00000000} /* (16, 30, 1) {real, imag} */,
  {32'hc51a9478, 32'h00000000} /* (16, 30, 0) {real, imag} */,
  {32'hc50cb5b6, 32'h00000000} /* (16, 29, 31) {real, imag} */,
  {32'hc53ae7c9, 32'h00000000} /* (16, 29, 30) {real, imag} */,
  {32'hc559f73f, 32'h00000000} /* (16, 29, 29) {real, imag} */,
  {32'hc550915f, 32'h00000000} /* (16, 29, 28) {real, imag} */,
  {32'hc54084e3, 32'h00000000} /* (16, 29, 27) {real, imag} */,
  {32'hc4eabe32, 32'h00000000} /* (16, 29, 26) {real, imag} */,
  {32'hc4ea2bea, 32'h00000000} /* (16, 29, 25) {real, imag} */,
  {32'hc51a6aa8, 32'h00000000} /* (16, 29, 24) {real, imag} */,
  {32'hc5272940, 32'h00000000} /* (16, 29, 23) {real, imag} */,
  {32'hc4260d70, 32'h00000000} /* (16, 29, 22) {real, imag} */,
  {32'h439d8dc4, 32'h00000000} /* (16, 29, 21) {real, imag} */,
  {32'h44d410e1, 32'h00000000} /* (16, 29, 20) {real, imag} */,
  {32'h44d29d9a, 32'h00000000} /* (16, 29, 19) {real, imag} */,
  {32'h44cdff82, 32'h00000000} /* (16, 29, 18) {real, imag} */,
  {32'h45397862, 32'h00000000} /* (16, 29, 17) {real, imag} */,
  {32'h450e6e8a, 32'h00000000} /* (16, 29, 16) {real, imag} */,
  {32'h453a4284, 32'h00000000} /* (16, 29, 15) {real, imag} */,
  {32'h454022f5, 32'h00000000} /* (16, 29, 14) {real, imag} */,
  {32'h451e9fbf, 32'h00000000} /* (16, 29, 13) {real, imag} */,
  {32'h451cb237, 32'h00000000} /* (16, 29, 12) {real, imag} */,
  {32'h45026873, 32'h00000000} /* (16, 29, 11) {real, imag} */,
  {32'h4465df48, 32'h00000000} /* (16, 29, 10) {real, imag} */,
  {32'hc4c6cdbc, 32'h00000000} /* (16, 29, 9) {real, imag} */,
  {32'hc51d8ac0, 32'h00000000} /* (16, 29, 8) {real, imag} */,
  {32'hc519f44c, 32'h00000000} /* (16, 29, 7) {real, imag} */,
  {32'hc5435016, 32'h00000000} /* (16, 29, 6) {real, imag} */,
  {32'hc51a3cd4, 32'h00000000} /* (16, 29, 5) {real, imag} */,
  {32'hc53ee6da, 32'h00000000} /* (16, 29, 4) {real, imag} */,
  {32'hc562e539, 32'h00000000} /* (16, 29, 3) {real, imag} */,
  {32'hc58b9b24, 32'h00000000} /* (16, 29, 2) {real, imag} */,
  {32'hc5685a42, 32'h00000000} /* (16, 29, 1) {real, imag} */,
  {32'hc5381076, 32'h00000000} /* (16, 29, 0) {real, imag} */,
  {32'hc55b2396, 32'h00000000} /* (16, 28, 31) {real, imag} */,
  {32'hc55e2167, 32'h00000000} /* (16, 28, 30) {real, imag} */,
  {32'hc51cbeb5, 32'h00000000} /* (16, 28, 29) {real, imag} */,
  {32'hc5202c5c, 32'h00000000} /* (16, 28, 28) {real, imag} */,
  {32'hc53934d6, 32'h00000000} /* (16, 28, 27) {real, imag} */,
  {32'hc51e11ae, 32'h00000000} /* (16, 28, 26) {real, imag} */,
  {32'hc538bc3a, 32'h00000000} /* (16, 28, 25) {real, imag} */,
  {32'hc53dc102, 32'h00000000} /* (16, 28, 24) {real, imag} */,
  {32'hc5380702, 32'h00000000} /* (16, 28, 23) {real, imag} */,
  {32'hc3df8c34, 32'h00000000} /* (16, 28, 22) {real, imag} */,
  {32'h43f790f4, 32'h00000000} /* (16, 28, 21) {real, imag} */,
  {32'h43f75cdc, 32'h00000000} /* (16, 28, 20) {real, imag} */,
  {32'h43bc0810, 32'h00000000} /* (16, 28, 19) {real, imag} */,
  {32'h453c42a0, 32'h00000000} /* (16, 28, 18) {real, imag} */,
  {32'h44f8029e, 32'h00000000} /* (16, 28, 17) {real, imag} */,
  {32'h45098ac8, 32'h00000000} /* (16, 28, 16) {real, imag} */,
  {32'h453a397c, 32'h00000000} /* (16, 28, 15) {real, imag} */,
  {32'h45488cb3, 32'h00000000} /* (16, 28, 14) {real, imag} */,
  {32'h4554be67, 32'h00000000} /* (16, 28, 13) {real, imag} */,
  {32'h451b7752, 32'h00000000} /* (16, 28, 12) {real, imag} */,
  {32'h44c5f27f, 32'h00000000} /* (16, 28, 11) {real, imag} */,
  {32'h439c8e04, 32'h00000000} /* (16, 28, 10) {real, imag} */,
  {32'hc4ef4284, 32'h00000000} /* (16, 28, 9) {real, imag} */,
  {32'hc4fdfe8d, 32'h00000000} /* (16, 28, 8) {real, imag} */,
  {32'hc5004f06, 32'h00000000} /* (16, 28, 7) {real, imag} */,
  {32'hc53d808e, 32'h00000000} /* (16, 28, 6) {real, imag} */,
  {32'hc525ed10, 32'h00000000} /* (16, 28, 5) {real, imag} */,
  {32'hc53d53ec, 32'h00000000} /* (16, 28, 4) {real, imag} */,
  {32'hc591ee8d, 32'h00000000} /* (16, 28, 3) {real, imag} */,
  {32'hc57914ce, 32'h00000000} /* (16, 28, 2) {real, imag} */,
  {32'hc5859ab4, 32'h00000000} /* (16, 28, 1) {real, imag} */,
  {32'hc532053a, 32'h00000000} /* (16, 28, 0) {real, imag} */,
  {32'hc5310ea2, 32'h00000000} /* (16, 27, 31) {real, imag} */,
  {32'hc5325b06, 32'h00000000} /* (16, 27, 30) {real, imag} */,
  {32'hc53178be, 32'h00000000} /* (16, 27, 29) {real, imag} */,
  {32'hc52a5f7e, 32'h00000000} /* (16, 27, 28) {real, imag} */,
  {32'hc521087c, 32'h00000000} /* (16, 27, 27) {real, imag} */,
  {32'hc51033ed, 32'h00000000} /* (16, 27, 26) {real, imag} */,
  {32'hc50305d2, 32'h00000000} /* (16, 27, 25) {real, imag} */,
  {32'hc5406864, 32'h00000000} /* (16, 27, 24) {real, imag} */,
  {32'hc4f0d56f, 32'h00000000} /* (16, 27, 23) {real, imag} */,
  {32'hc477bf5e, 32'h00000000} /* (16, 27, 22) {real, imag} */,
  {32'h43b03af4, 32'h00000000} /* (16, 27, 21) {real, imag} */,
  {32'h448f5862, 32'h00000000} /* (16, 27, 20) {real, imag} */,
  {32'h44b33065, 32'h00000000} /* (16, 27, 19) {real, imag} */,
  {32'h44cd547f, 32'h00000000} /* (16, 27, 18) {real, imag} */,
  {32'h448f24c4, 32'h00000000} /* (16, 27, 17) {real, imag} */,
  {32'h44d1e972, 32'h00000000} /* (16, 27, 16) {real, imag} */,
  {32'h45375294, 32'h00000000} /* (16, 27, 15) {real, imag} */,
  {32'h451d8718, 32'h00000000} /* (16, 27, 14) {real, imag} */,
  {32'h4500f754, 32'h00000000} /* (16, 27, 13) {real, imag} */,
  {32'h44e4ffb0, 32'h00000000} /* (16, 27, 12) {real, imag} */,
  {32'h4497639b, 32'h00000000} /* (16, 27, 11) {real, imag} */,
  {32'hc2f720c0, 32'h00000000} /* (16, 27, 10) {real, imag} */,
  {32'hc4e90cd0, 32'h00000000} /* (16, 27, 9) {real, imag} */,
  {32'hc4f200b5, 32'h00000000} /* (16, 27, 8) {real, imag} */,
  {32'hc52dc120, 32'h00000000} /* (16, 27, 7) {real, imag} */,
  {32'hc526f956, 32'h00000000} /* (16, 27, 6) {real, imag} */,
  {32'hc51ff71c, 32'h00000000} /* (16, 27, 5) {real, imag} */,
  {32'hc557d4cb, 32'h00000000} /* (16, 27, 4) {real, imag} */,
  {32'hc5653542, 32'h00000000} /* (16, 27, 3) {real, imag} */,
  {32'hc560b184, 32'h00000000} /* (16, 27, 2) {real, imag} */,
  {32'hc56b83f6, 32'h00000000} /* (16, 27, 1) {real, imag} */,
  {32'hc553ec8f, 32'h00000000} /* (16, 27, 0) {real, imag} */,
  {32'hc52be629, 32'h00000000} /* (16, 26, 31) {real, imag} */,
  {32'hc5494020, 32'h00000000} /* (16, 26, 30) {real, imag} */,
  {32'hc507ed6d, 32'h00000000} /* (16, 26, 29) {real, imag} */,
  {32'hc515f594, 32'h00000000} /* (16, 26, 28) {real, imag} */,
  {32'hc54173f2, 32'h00000000} /* (16, 26, 27) {real, imag} */,
  {32'hc5130d64, 32'h00000000} /* (16, 26, 26) {real, imag} */,
  {32'hc50e917e, 32'h00000000} /* (16, 26, 25) {real, imag} */,
  {32'hc53c9a61, 32'h00000000} /* (16, 26, 24) {real, imag} */,
  {32'hc4bfdf23, 32'h00000000} /* (16, 26, 23) {real, imag} */,
  {32'hc441e8f8, 32'h00000000} /* (16, 26, 22) {real, imag} */,
  {32'hc33d1628, 32'h00000000} /* (16, 26, 21) {real, imag} */,
  {32'h44bb13fc, 32'h00000000} /* (16, 26, 20) {real, imag} */,
  {32'h4462e6f4, 32'h00000000} /* (16, 26, 19) {real, imag} */,
  {32'h4477b2aa, 32'h00000000} /* (16, 26, 18) {real, imag} */,
  {32'h44e23a5c, 32'h00000000} /* (16, 26, 17) {real, imag} */,
  {32'h44ac92fe, 32'h00000000} /* (16, 26, 16) {real, imag} */,
  {32'h44c013ae, 32'h00000000} /* (16, 26, 15) {real, imag} */,
  {32'h44dcd710, 32'h00000000} /* (16, 26, 14) {real, imag} */,
  {32'h44b3dfd4, 32'h00000000} /* (16, 26, 13) {real, imag} */,
  {32'h44aa7702, 32'h00000000} /* (16, 26, 12) {real, imag} */,
  {32'h44249650, 32'h00000000} /* (16, 26, 11) {real, imag} */,
  {32'hc36938f8, 32'h00000000} /* (16, 26, 10) {real, imag} */,
  {32'hc4f4b2ad, 32'h00000000} /* (16, 26, 9) {real, imag} */,
  {32'hc50a8bdd, 32'h00000000} /* (16, 26, 8) {real, imag} */,
  {32'hc5262c68, 32'h00000000} /* (16, 26, 7) {real, imag} */,
  {32'hc5359bf8, 32'h00000000} /* (16, 26, 6) {real, imag} */,
  {32'hc52b4706, 32'h00000000} /* (16, 26, 5) {real, imag} */,
  {32'hc533b70e, 32'h00000000} /* (16, 26, 4) {real, imag} */,
  {32'hc5363863, 32'h00000000} /* (16, 26, 3) {real, imag} */,
  {32'hc58a22b5, 32'h00000000} /* (16, 26, 2) {real, imag} */,
  {32'hc573d046, 32'h00000000} /* (16, 26, 1) {real, imag} */,
  {32'hc5488a87, 32'h00000000} /* (16, 26, 0) {real, imag} */,
  {32'hc52b8ba8, 32'h00000000} /* (16, 25, 31) {real, imag} */,
  {32'hc533f1ca, 32'h00000000} /* (16, 25, 30) {real, imag} */,
  {32'hc53952bc, 32'h00000000} /* (16, 25, 29) {real, imag} */,
  {32'hc51486d6, 32'h00000000} /* (16, 25, 28) {real, imag} */,
  {32'hc50e5702, 32'h00000000} /* (16, 25, 27) {real, imag} */,
  {32'hc51a25d2, 32'h00000000} /* (16, 25, 26) {real, imag} */,
  {32'hc5243584, 32'h00000000} /* (16, 25, 25) {real, imag} */,
  {32'hc51a2de5, 32'h00000000} /* (16, 25, 24) {real, imag} */,
  {32'hc510efb0, 32'h00000000} /* (16, 25, 23) {real, imag} */,
  {32'hc4c98824, 32'h00000000} /* (16, 25, 22) {real, imag} */,
  {32'hc2c3fd90, 32'h00000000} /* (16, 25, 21) {real, imag} */,
  {32'h44b58add, 32'h00000000} /* (16, 25, 20) {real, imag} */,
  {32'h44b09939, 32'h00000000} /* (16, 25, 19) {real, imag} */,
  {32'h446cd118, 32'h00000000} /* (16, 25, 18) {real, imag} */,
  {32'h44a798fe, 32'h00000000} /* (16, 25, 17) {real, imag} */,
  {32'h44bc5dfc, 32'h00000000} /* (16, 25, 16) {real, imag} */,
  {32'h44f8ad40, 32'h00000000} /* (16, 25, 15) {real, imag} */,
  {32'h44807164, 32'h00000000} /* (16, 25, 14) {real, imag} */,
  {32'h4508392c, 32'h00000000} /* (16, 25, 13) {real, imag} */,
  {32'h447ef386, 32'h00000000} /* (16, 25, 12) {real, imag} */,
  {32'h445bb15a, 32'h00000000} /* (16, 25, 11) {real, imag} */,
  {32'hc430aa96, 32'h00000000} /* (16, 25, 10) {real, imag} */,
  {32'hc5079aba, 32'h00000000} /* (16, 25, 9) {real, imag} */,
  {32'hc4cca02a, 32'h00000000} /* (16, 25, 8) {real, imag} */,
  {32'hc4d65478, 32'h00000000} /* (16, 25, 7) {real, imag} */,
  {32'hc51bb694, 32'h00000000} /* (16, 25, 6) {real, imag} */,
  {32'hc5141c0e, 32'h00000000} /* (16, 25, 5) {real, imag} */,
  {32'hc53d6fda, 32'h00000000} /* (16, 25, 4) {real, imag} */,
  {32'hc56218a2, 32'h00000000} /* (16, 25, 3) {real, imag} */,
  {32'hc55ff0e8, 32'h00000000} /* (16, 25, 2) {real, imag} */,
  {32'hc57d7a29, 32'h00000000} /* (16, 25, 1) {real, imag} */,
  {32'hc52f0d74, 32'h00000000} /* (16, 25, 0) {real, imag} */,
  {32'hc52e9745, 32'h00000000} /* (16, 24, 31) {real, imag} */,
  {32'hc4fb9ad7, 32'h00000000} /* (16, 24, 30) {real, imag} */,
  {32'hc4d2a824, 32'h00000000} /* (16, 24, 29) {real, imag} */,
  {32'hc4dc8d9a, 32'h00000000} /* (16, 24, 28) {real, imag} */,
  {32'hc5277d42, 32'h00000000} /* (16, 24, 27) {real, imag} */,
  {32'hc52045d2, 32'h00000000} /* (16, 24, 26) {real, imag} */,
  {32'hc51f332d, 32'h00000000} /* (16, 24, 25) {real, imag} */,
  {32'hc54d2455, 32'h00000000} /* (16, 24, 24) {real, imag} */,
  {32'hc521d7c6, 32'h00000000} /* (16, 24, 23) {real, imag} */,
  {32'hc4e9ee26, 32'h00000000} /* (16, 24, 22) {real, imag} */,
  {32'hc361ef28, 32'h00000000} /* (16, 24, 21) {real, imag} */,
  {32'h4389407c, 32'h00000000} /* (16, 24, 20) {real, imag} */,
  {32'h44d39344, 32'h00000000} /* (16, 24, 19) {real, imag} */,
  {32'h448bf424, 32'h00000000} /* (16, 24, 18) {real, imag} */,
  {32'h44ddd114, 32'h00000000} /* (16, 24, 17) {real, imag} */,
  {32'h44e2f6eb, 32'h00000000} /* (16, 24, 16) {real, imag} */,
  {32'h4454b235, 32'h00000000} /* (16, 24, 15) {real, imag} */,
  {32'h44d4657d, 32'h00000000} /* (16, 24, 14) {real, imag} */,
  {32'h44939fd0, 32'h00000000} /* (16, 24, 13) {real, imag} */,
  {32'h45080074, 32'h00000000} /* (16, 24, 12) {real, imag} */,
  {32'h448032b0, 32'h00000000} /* (16, 24, 11) {real, imag} */,
  {32'hc4a0cb88, 32'h00000000} /* (16, 24, 10) {real, imag} */,
  {32'hc520191d, 32'h00000000} /* (16, 24, 9) {real, imag} */,
  {32'hc4f8eb3e, 32'h00000000} /* (16, 24, 8) {real, imag} */,
  {32'hc4f0cc64, 32'h00000000} /* (16, 24, 7) {real, imag} */,
  {32'hc4f1fbf4, 32'h00000000} /* (16, 24, 6) {real, imag} */,
  {32'hc52f62e8, 32'h00000000} /* (16, 24, 5) {real, imag} */,
  {32'hc51794be, 32'h00000000} /* (16, 24, 4) {real, imag} */,
  {32'hc558aa8c, 32'h00000000} /* (16, 24, 3) {real, imag} */,
  {32'hc5840039, 32'h00000000} /* (16, 24, 2) {real, imag} */,
  {32'hc5597068, 32'h00000000} /* (16, 24, 1) {real, imag} */,
  {32'hc50d27ca, 32'h00000000} /* (16, 24, 0) {real, imag} */,
  {32'hc4e99b25, 32'h00000000} /* (16, 23, 31) {real, imag} */,
  {32'hc4c4552a, 32'h00000000} /* (16, 23, 30) {real, imag} */,
  {32'hc496bb17, 32'h00000000} /* (16, 23, 29) {real, imag} */,
  {32'hc4f09c78, 32'h00000000} /* (16, 23, 28) {real, imag} */,
  {32'hc52fea8a, 32'h00000000} /* (16, 23, 27) {real, imag} */,
  {32'hc55bb656, 32'h00000000} /* (16, 23, 26) {real, imag} */,
  {32'hc50ac4e8, 32'h00000000} /* (16, 23, 25) {real, imag} */,
  {32'hc50bca80, 32'h00000000} /* (16, 23, 24) {real, imag} */,
  {32'hc543bfb6, 32'h00000000} /* (16, 23, 23) {real, imag} */,
  {32'hc4c9b162, 32'h00000000} /* (16, 23, 22) {real, imag} */,
  {32'hc481fcac, 32'h00000000} /* (16, 23, 21) {real, imag} */,
  {32'h44a5fd0c, 32'h00000000} /* (16, 23, 20) {real, imag} */,
  {32'h4437fa20, 32'h00000000} /* (16, 23, 19) {real, imag} */,
  {32'h4497cfd1, 32'h00000000} /* (16, 23, 18) {real, imag} */,
  {32'h445a03e2, 32'h00000000} /* (16, 23, 17) {real, imag} */,
  {32'h44a4aabd, 32'h00000000} /* (16, 23, 16) {real, imag} */,
  {32'h44c9139f, 32'h00000000} /* (16, 23, 15) {real, imag} */,
  {32'h448646be, 32'h00000000} /* (16, 23, 14) {real, imag} */,
  {32'h4487df1d, 32'h00000000} /* (16, 23, 13) {real, imag} */,
  {32'h449023f8, 32'h00000000} /* (16, 23, 12) {real, imag} */,
  {32'hc37dd7d8, 32'h00000000} /* (16, 23, 11) {real, imag} */,
  {32'hc4e9de7c, 32'h00000000} /* (16, 23, 10) {real, imag} */,
  {32'hc4d467f2, 32'h00000000} /* (16, 23, 9) {real, imag} */,
  {32'hc5084204, 32'h00000000} /* (16, 23, 8) {real, imag} */,
  {32'hc4a8f77d, 32'h00000000} /* (16, 23, 7) {real, imag} */,
  {32'hc4bc75fa, 32'h00000000} /* (16, 23, 6) {real, imag} */,
  {32'hc5397b75, 32'h00000000} /* (16, 23, 5) {real, imag} */,
  {32'hc4aad60e, 32'h00000000} /* (16, 23, 4) {real, imag} */,
  {32'hc4afa842, 32'h00000000} /* (16, 23, 3) {real, imag} */,
  {32'hc53bda52, 32'h00000000} /* (16, 23, 2) {real, imag} */,
  {32'hc5346fb0, 32'h00000000} /* (16, 23, 1) {real, imag} */,
  {32'hc501c422, 32'h00000000} /* (16, 23, 0) {real, imag} */,
  {32'hc4f5049c, 32'h00000000} /* (16, 22, 31) {real, imag} */,
  {32'hc4baa078, 32'h00000000} /* (16, 22, 30) {real, imag} */,
  {32'hc4d0486c, 32'h00000000} /* (16, 22, 29) {real, imag} */,
  {32'hc4dba952, 32'h00000000} /* (16, 22, 28) {real, imag} */,
  {32'hc4e38ee9, 32'h00000000} /* (16, 22, 27) {real, imag} */,
  {32'hc5085ab2, 32'h00000000} /* (16, 22, 26) {real, imag} */,
  {32'hc516a43c, 32'h00000000} /* (16, 22, 25) {real, imag} */,
  {32'hc50b937a, 32'h00000000} /* (16, 22, 24) {real, imag} */,
  {32'hc4e1254e, 32'h00000000} /* (16, 22, 23) {real, imag} */,
  {32'hc4dc89cb, 32'h00000000} /* (16, 22, 22) {real, imag} */,
  {32'hc4766d59, 32'h00000000} /* (16, 22, 21) {real, imag} */,
  {32'h448ef299, 32'h00000000} /* (16, 22, 20) {real, imag} */,
  {32'h4469f6ee, 32'h00000000} /* (16, 22, 19) {real, imag} */,
  {32'h44129a5c, 32'h00000000} /* (16, 22, 18) {real, imag} */,
  {32'h443a2c18, 32'h00000000} /* (16, 22, 17) {real, imag} */,
  {32'h449222c0, 32'h00000000} /* (16, 22, 16) {real, imag} */,
  {32'h44791528, 32'h00000000} /* (16, 22, 15) {real, imag} */,
  {32'h449204aa, 32'h00000000} /* (16, 22, 14) {real, imag} */,
  {32'h44c7b8e8, 32'h00000000} /* (16, 22, 13) {real, imag} */,
  {32'hc3485250, 32'h00000000} /* (16, 22, 12) {real, imag} */,
  {32'h423200a0, 32'h00000000} /* (16, 22, 11) {real, imag} */,
  {32'hc450d82c, 32'h00000000} /* (16, 22, 10) {real, imag} */,
  {32'hc4dee784, 32'h00000000} /* (16, 22, 9) {real, imag} */,
  {32'hc4fd266b, 32'h00000000} /* (16, 22, 8) {real, imag} */,
  {32'hc4d4fc7a, 32'h00000000} /* (16, 22, 7) {real, imag} */,
  {32'hc4e21e3b, 32'h00000000} /* (16, 22, 6) {real, imag} */,
  {32'hc48154a8, 32'h00000000} /* (16, 22, 5) {real, imag} */,
  {32'hc4d052c5, 32'h00000000} /* (16, 22, 4) {real, imag} */,
  {32'hc4f02d7d, 32'h00000000} /* (16, 22, 3) {real, imag} */,
  {32'hc4e75018, 32'h00000000} /* (16, 22, 2) {real, imag} */,
  {32'hc52794ec, 32'h00000000} /* (16, 22, 1) {real, imag} */,
  {32'hc4b2d98e, 32'h00000000} /* (16, 22, 0) {real, imag} */,
  {32'hc41bec78, 32'h00000000} /* (16, 21, 31) {real, imag} */,
  {32'hc4480621, 32'h00000000} /* (16, 21, 30) {real, imag} */,
  {32'hc4af6ad1, 32'h00000000} /* (16, 21, 29) {real, imag} */,
  {32'hc4b25108, 32'h00000000} /* (16, 21, 28) {real, imag} */,
  {32'hc4d3b721, 32'h00000000} /* (16, 21, 27) {real, imag} */,
  {32'hc4f34963, 32'h00000000} /* (16, 21, 26) {real, imag} */,
  {32'hc4d3034a, 32'h00000000} /* (16, 21, 25) {real, imag} */,
  {32'hc4ab8c2c, 32'h00000000} /* (16, 21, 24) {real, imag} */,
  {32'hc3a89a0a, 32'h00000000} /* (16, 21, 23) {real, imag} */,
  {32'hc3ed6ea4, 32'h00000000} /* (16, 21, 22) {real, imag} */,
  {32'hc4025e05, 32'h00000000} /* (16, 21, 21) {real, imag} */,
  {32'hc3cf68cd, 32'h00000000} /* (16, 21, 20) {real, imag} */,
  {32'h44330ec8, 32'h00000000} /* (16, 21, 19) {real, imag} */,
  {32'hc2b0bde8, 32'h00000000} /* (16, 21, 18) {real, imag} */,
  {32'h433662e2, 32'h00000000} /* (16, 21, 17) {real, imag} */,
  {32'h438b9d34, 32'h00000000} /* (16, 21, 16) {real, imag} */,
  {32'h443bc640, 32'h00000000} /* (16, 21, 15) {real, imag} */,
  {32'h4429a603, 32'h00000000} /* (16, 21, 14) {real, imag} */,
  {32'hc3ef126f, 32'h00000000} /* (16, 21, 13) {real, imag} */,
  {32'hc3c6001e, 32'h00000000} /* (16, 21, 12) {real, imag} */,
  {32'hc441fb92, 32'h00000000} /* (16, 21, 11) {real, imag} */,
  {32'hc38953cc, 32'h00000000} /* (16, 21, 10) {real, imag} */,
  {32'hc47c0a6f, 32'h00000000} /* (16, 21, 9) {real, imag} */,
  {32'hc4b3d764, 32'h00000000} /* (16, 21, 8) {real, imag} */,
  {32'hc43175f7, 32'h00000000} /* (16, 21, 7) {real, imag} */,
  {32'hc4ae1aba, 32'h00000000} /* (16, 21, 6) {real, imag} */,
  {32'hc48fa7d4, 32'h00000000} /* (16, 21, 5) {real, imag} */,
  {32'hc32af58e, 32'h00000000} /* (16, 21, 4) {real, imag} */,
  {32'hc4d846e2, 32'h00000000} /* (16, 21, 3) {real, imag} */,
  {32'hc49073b2, 32'h00000000} /* (16, 21, 2) {real, imag} */,
  {32'hc3eeae59, 32'h00000000} /* (16, 21, 1) {real, imag} */,
  {32'hc427f804, 32'h00000000} /* (16, 21, 0) {real, imag} */,
  {32'h44019c36, 32'h00000000} /* (16, 20, 31) {real, imag} */,
  {32'h44708f46, 32'h00000000} /* (16, 20, 30) {real, imag} */,
  {32'hc1f59f90, 32'h00000000} /* (16, 20, 29) {real, imag} */,
  {32'hc450562d, 32'h00000000} /* (16, 20, 28) {real, imag} */,
  {32'hc4a9c655, 32'h00000000} /* (16, 20, 27) {real, imag} */,
  {32'hc3cf56f9, 32'h00000000} /* (16, 20, 26) {real, imag} */,
  {32'h41be6950, 32'h00000000} /* (16, 20, 25) {real, imag} */,
  {32'h44886f2f, 32'h00000000} /* (16, 20, 24) {real, imag} */,
  {32'h4457d15c, 32'h00000000} /* (16, 20, 23) {real, imag} */,
  {32'h43110cda, 32'h00000000} /* (16, 20, 22) {real, imag} */,
  {32'hc2748efc, 32'h00000000} /* (16, 20, 21) {real, imag} */,
  {32'hc43610fe, 32'h00000000} /* (16, 20, 20) {real, imag} */,
  {32'hc426ba9c, 32'h00000000} /* (16, 20, 19) {real, imag} */,
  {32'hc36c0024, 32'h00000000} /* (16, 20, 18) {real, imag} */,
  {32'hc42a46b2, 32'h00000000} /* (16, 20, 17) {real, imag} */,
  {32'hc47c0770, 32'h00000000} /* (16, 20, 16) {real, imag} */,
  {32'h4369dcde, 32'h00000000} /* (16, 20, 15) {real, imag} */,
  {32'h44000222, 32'h00000000} /* (16, 20, 14) {real, imag} */,
  {32'hc4498132, 32'h00000000} /* (16, 20, 13) {real, imag} */,
  {32'hc4ee40ec, 32'h00000000} /* (16, 20, 12) {real, imag} */,
  {32'hc4792616, 32'h00000000} /* (16, 20, 11) {real, imag} */,
  {32'hc460f2f0, 32'h00000000} /* (16, 20, 10) {real, imag} */,
  {32'h443f4602, 32'h00000000} /* (16, 20, 9) {real, imag} */,
  {32'h441474fa, 32'h00000000} /* (16, 20, 8) {real, imag} */,
  {32'hc042bf80, 32'h00000000} /* (16, 20, 7) {real, imag} */,
  {32'h43a6d14d, 32'h00000000} /* (16, 20, 6) {real, imag} */,
  {32'h43f54b8a, 32'h00000000} /* (16, 20, 5) {real, imag} */,
  {32'h44015562, 32'h00000000} /* (16, 20, 4) {real, imag} */,
  {32'h449a1ba8, 32'h00000000} /* (16, 20, 3) {real, imag} */,
  {32'h44b01f90, 32'h00000000} /* (16, 20, 2) {real, imag} */,
  {32'h4353f36e, 32'h00000000} /* (16, 20, 1) {real, imag} */,
  {32'h43dafe2d, 32'h00000000} /* (16, 20, 0) {real, imag} */,
  {32'h44473271, 32'h00000000} /* (16, 19, 31) {real, imag} */,
  {32'h4422dc19, 32'h00000000} /* (16, 19, 30) {real, imag} */,
  {32'h43b41009, 32'h00000000} /* (16, 19, 29) {real, imag} */,
  {32'h4394980d, 32'h00000000} /* (16, 19, 28) {real, imag} */,
  {32'hc266cbc0, 32'h00000000} /* (16, 19, 27) {real, imag} */,
  {32'h43f45174, 32'h00000000} /* (16, 19, 26) {real, imag} */,
  {32'h43df3162, 32'h00000000} /* (16, 19, 25) {real, imag} */,
  {32'h443821b1, 32'h00000000} /* (16, 19, 24) {real, imag} */,
  {32'h44cfffab, 32'h00000000} /* (16, 19, 23) {real, imag} */,
  {32'h45140952, 32'h00000000} /* (16, 19, 22) {real, imag} */,
  {32'h4442ac34, 32'h00000000} /* (16, 19, 21) {real, imag} */,
  {32'hc418a7b6, 32'h00000000} /* (16, 19, 20) {real, imag} */,
  {32'hc4c4a5f2, 32'h00000000} /* (16, 19, 19) {real, imag} */,
  {32'hc3c6a9f6, 32'h00000000} /* (16, 19, 18) {real, imag} */,
  {32'hc375bf00, 32'h00000000} /* (16, 19, 17) {real, imag} */,
  {32'hc4c306d8, 32'h00000000} /* (16, 19, 16) {real, imag} */,
  {32'hc4b0a502, 32'h00000000} /* (16, 19, 15) {real, imag} */,
  {32'hc48bf2cc, 32'h00000000} /* (16, 19, 14) {real, imag} */,
  {32'hc48dd073, 32'h00000000} /* (16, 19, 13) {real, imag} */,
  {32'hc43d46f0, 32'h00000000} /* (16, 19, 12) {real, imag} */,
  {32'hc49bd0fd, 32'h00000000} /* (16, 19, 11) {real, imag} */,
  {32'h44219ba0, 32'h00000000} /* (16, 19, 10) {real, imag} */,
  {32'h44bd51e6, 32'h00000000} /* (16, 19, 9) {real, imag} */,
  {32'h44449c45, 32'h00000000} /* (16, 19, 8) {real, imag} */,
  {32'h4403d40a, 32'h00000000} /* (16, 19, 7) {real, imag} */,
  {32'h44431446, 32'h00000000} /* (16, 19, 6) {real, imag} */,
  {32'h44bf9516, 32'h00000000} /* (16, 19, 5) {real, imag} */,
  {32'h44b0cc1b, 32'h00000000} /* (16, 19, 4) {real, imag} */,
  {32'h44b180d8, 32'h00000000} /* (16, 19, 3) {real, imag} */,
  {32'h44d9149a, 32'h00000000} /* (16, 19, 2) {real, imag} */,
  {32'h45176398, 32'h00000000} /* (16, 19, 1) {real, imag} */,
  {32'h449beb6e, 32'h00000000} /* (16, 19, 0) {real, imag} */,
  {32'h44dece78, 32'h00000000} /* (16, 18, 31) {real, imag} */,
  {32'h44b1a24c, 32'h00000000} /* (16, 18, 30) {real, imag} */,
  {32'h444a50e8, 32'h00000000} /* (16, 18, 29) {real, imag} */,
  {32'h44482e4f, 32'h00000000} /* (16, 18, 28) {real, imag} */,
  {32'h44c2faf8, 32'h00000000} /* (16, 18, 27) {real, imag} */,
  {32'h4500ecfa, 32'h00000000} /* (16, 18, 26) {real, imag} */,
  {32'h448a0225, 32'h00000000} /* (16, 18, 25) {real, imag} */,
  {32'h4524de5e, 32'h00000000} /* (16, 18, 24) {real, imag} */,
  {32'h452b00e7, 32'h00000000} /* (16, 18, 23) {real, imag} */,
  {32'h44635772, 32'h00000000} /* (16, 18, 22) {real, imag} */,
  {32'h447abac8, 32'h00000000} /* (16, 18, 21) {real, imag} */,
  {32'hc381d560, 32'h00000000} /* (16, 18, 20) {real, imag} */,
  {32'hc48988d7, 32'h00000000} /* (16, 18, 19) {real, imag} */,
  {32'hc4ef998c, 32'h00000000} /* (16, 18, 18) {real, imag} */,
  {32'hc513d640, 32'h00000000} /* (16, 18, 17) {real, imag} */,
  {32'hc4e6f153, 32'h00000000} /* (16, 18, 16) {real, imag} */,
  {32'hc4e5b4bc, 32'h00000000} /* (16, 18, 15) {real, imag} */,
  {32'hc48cfa04, 32'h00000000} /* (16, 18, 14) {real, imag} */,
  {32'hc4d905a4, 32'h00000000} /* (16, 18, 13) {real, imag} */,
  {32'hc3dc7cc6, 32'h00000000} /* (16, 18, 12) {real, imag} */,
  {32'hc329b50c, 32'h00000000} /* (16, 18, 11) {real, imag} */,
  {32'h449cae50, 32'h00000000} /* (16, 18, 10) {real, imag} */,
  {32'h44fe9bf3, 32'h00000000} /* (16, 18, 9) {real, imag} */,
  {32'h44a14d4a, 32'h00000000} /* (16, 18, 8) {real, imag} */,
  {32'h44905dda, 32'h00000000} /* (16, 18, 7) {real, imag} */,
  {32'h4496f0f5, 32'h00000000} /* (16, 18, 6) {real, imag} */,
  {32'h449160c0, 32'h00000000} /* (16, 18, 5) {real, imag} */,
  {32'h450ba759, 32'h00000000} /* (16, 18, 4) {real, imag} */,
  {32'h44a31011, 32'h00000000} /* (16, 18, 3) {real, imag} */,
  {32'h44e90e06, 32'h00000000} /* (16, 18, 2) {real, imag} */,
  {32'h452dedb0, 32'h00000000} /* (16, 18, 1) {real, imag} */,
  {32'h44ed8e79, 32'h00000000} /* (16, 18, 0) {real, imag} */,
  {32'h4507cf38, 32'h00000000} /* (16, 17, 31) {real, imag} */,
  {32'h44ef9e42, 32'h00000000} /* (16, 17, 30) {real, imag} */,
  {32'h44a130a2, 32'h00000000} /* (16, 17, 29) {real, imag} */,
  {32'h44f211c0, 32'h00000000} /* (16, 17, 28) {real, imag} */,
  {32'h44be6c26, 32'h00000000} /* (16, 17, 27) {real, imag} */,
  {32'h44afbaa6, 32'h00000000} /* (16, 17, 26) {real, imag} */,
  {32'h451af26b, 32'h00000000} /* (16, 17, 25) {real, imag} */,
  {32'h4541b83a, 32'h00000000} /* (16, 17, 24) {real, imag} */,
  {32'h4475055b, 32'h00000000} /* (16, 17, 23) {real, imag} */,
  {32'h44e9093e, 32'h00000000} /* (16, 17, 22) {real, imag} */,
  {32'h44da4b9b, 32'h00000000} /* (16, 17, 21) {real, imag} */,
  {32'hc485e4de, 32'h00000000} /* (16, 17, 20) {real, imag} */,
  {32'hc463ff47, 32'h00000000} /* (16, 17, 19) {real, imag} */,
  {32'hc4d95710, 32'h00000000} /* (16, 17, 18) {real, imag} */,
  {32'hc50e5162, 32'h00000000} /* (16, 17, 17) {real, imag} */,
  {32'hc50788ec, 32'h00000000} /* (16, 17, 16) {real, imag} */,
  {32'hc51f650a, 32'h00000000} /* (16, 17, 15) {real, imag} */,
  {32'hc52ee4ef, 32'h00000000} /* (16, 17, 14) {real, imag} */,
  {32'hc5001185, 32'h00000000} /* (16, 17, 13) {real, imag} */,
  {32'hc456a61d, 32'h00000000} /* (16, 17, 12) {real, imag} */,
  {32'hc3b6419c, 32'h00000000} /* (16, 17, 11) {real, imag} */,
  {32'h44b04ca8, 32'h00000000} /* (16, 17, 10) {real, imag} */,
  {32'h453ac949, 32'h00000000} /* (16, 17, 9) {real, imag} */,
  {32'h4519b70e, 32'h00000000} /* (16, 17, 8) {real, imag} */,
  {32'h44af6e8f, 32'h00000000} /* (16, 17, 7) {real, imag} */,
  {32'h44881a2e, 32'h00000000} /* (16, 17, 6) {real, imag} */,
  {32'h4449e06a, 32'h00000000} /* (16, 17, 5) {real, imag} */,
  {32'h4503e0f5, 32'h00000000} /* (16, 17, 4) {real, imag} */,
  {32'h44f270ce, 32'h00000000} /* (16, 17, 3) {real, imag} */,
  {32'h448647b2, 32'h00000000} /* (16, 17, 2) {real, imag} */,
  {32'h44f98183, 32'h00000000} /* (16, 17, 1) {real, imag} */,
  {32'h45182dce, 32'h00000000} /* (16, 17, 0) {real, imag} */,
  {32'h44d18218, 32'h00000000} /* (16, 16, 31) {real, imag} */,
  {32'h448960ee, 32'h00000000} /* (16, 16, 30) {real, imag} */,
  {32'h44ed80db, 32'h00000000} /* (16, 16, 29) {real, imag} */,
  {32'h4508e19f, 32'h00000000} /* (16, 16, 28) {real, imag} */,
  {32'h44f90640, 32'h00000000} /* (16, 16, 27) {real, imag} */,
  {32'h449eb7f8, 32'h00000000} /* (16, 16, 26) {real, imag} */,
  {32'h4485d9e4, 32'h00000000} /* (16, 16, 25) {real, imag} */,
  {32'h44ea7982, 32'h00000000} /* (16, 16, 24) {real, imag} */,
  {32'h44a10b58, 32'h00000000} /* (16, 16, 23) {real, imag} */,
  {32'h44acbdf8, 32'h00000000} /* (16, 16, 22) {real, imag} */,
  {32'h43fd9374, 32'h00000000} /* (16, 16, 21) {real, imag} */,
  {32'hc4841a34, 32'h00000000} /* (16, 16, 20) {real, imag} */,
  {32'hc4ce71aa, 32'h00000000} /* (16, 16, 19) {real, imag} */,
  {32'hc4c69551, 32'h00000000} /* (16, 16, 18) {real, imag} */,
  {32'hc5124c0c, 32'h00000000} /* (16, 16, 17) {real, imag} */,
  {32'hc5202118, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'hc4e725a2, 32'h00000000} /* (16, 16, 15) {real, imag} */,
  {32'hc53c3279, 32'h00000000} /* (16, 16, 14) {real, imag} */,
  {32'hc4b151e1, 32'h00000000} /* (16, 16, 13) {real, imag} */,
  {32'hc509aeaf, 32'h00000000} /* (16, 16, 12) {real, imag} */,
  {32'hc45b6ad9, 32'h00000000} /* (16, 16, 11) {real, imag} */,
  {32'h44ce488a, 32'h00000000} /* (16, 16, 10) {real, imag} */,
  {32'h44c606ae, 32'h00000000} /* (16, 16, 9) {real, imag} */,
  {32'h4521459b, 32'h00000000} /* (16, 16, 8) {real, imag} */,
  {32'h44debf14, 32'h00000000} /* (16, 16, 7) {real, imag} */,
  {32'h442e66f9, 32'h00000000} /* (16, 16, 6) {real, imag} */,
  {32'h44b74ae1, 32'h00000000} /* (16, 16, 5) {real, imag} */,
  {32'h44bf6858, 32'h00000000} /* (16, 16, 4) {real, imag} */,
  {32'h4507a432, 32'h00000000} /* (16, 16, 3) {real, imag} */,
  {32'h451e2df4, 32'h00000000} /* (16, 16, 2) {real, imag} */,
  {32'h44e48195, 32'h00000000} /* (16, 16, 1) {real, imag} */,
  {32'h44b4b8b5, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'h4474d972, 32'h00000000} /* (16, 15, 31) {real, imag} */,
  {32'h44870c03, 32'h00000000} /* (16, 15, 30) {real, imag} */,
  {32'h44b75ea0, 32'h00000000} /* (16, 15, 29) {real, imag} */,
  {32'h450f2220, 32'h00000000} /* (16, 15, 28) {real, imag} */,
  {32'h44d07baa, 32'h00000000} /* (16, 15, 27) {real, imag} */,
  {32'h44a5b490, 32'h00000000} /* (16, 15, 26) {real, imag} */,
  {32'h443debab, 32'h00000000} /* (16, 15, 25) {real, imag} */,
  {32'h43b9e418, 32'h00000000} /* (16, 15, 24) {real, imag} */,
  {32'h445c3938, 32'h00000000} /* (16, 15, 23) {real, imag} */,
  {32'h44b309cc, 32'h00000000} /* (16, 15, 22) {real, imag} */,
  {32'h43c82c4c, 32'h00000000} /* (16, 15, 21) {real, imag} */,
  {32'hc44205e4, 32'h00000000} /* (16, 15, 20) {real, imag} */,
  {32'hc4aba937, 32'h00000000} /* (16, 15, 19) {real, imag} */,
  {32'hc4b074d4, 32'h00000000} /* (16, 15, 18) {real, imag} */,
  {32'hc4dc61a9, 32'h00000000} /* (16, 15, 17) {real, imag} */,
  {32'hc4ec26cc, 32'h00000000} /* (16, 15, 16) {real, imag} */,
  {32'hc5059c2e, 32'h00000000} /* (16, 15, 15) {real, imag} */,
  {32'hc508aa6a, 32'h00000000} /* (16, 15, 14) {real, imag} */,
  {32'hc498ef70, 32'h00000000} /* (16, 15, 13) {real, imag} */,
  {32'hc39e9da4, 32'h00000000} /* (16, 15, 12) {real, imag} */,
  {32'h43f5ed50, 32'h00000000} /* (16, 15, 11) {real, imag} */,
  {32'h44c1b938, 32'h00000000} /* (16, 15, 10) {real, imag} */,
  {32'h452675b4, 32'h00000000} /* (16, 15, 9) {real, imag} */,
  {32'h44e15526, 32'h00000000} /* (16, 15, 8) {real, imag} */,
  {32'h4507370f, 32'h00000000} /* (16, 15, 7) {real, imag} */,
  {32'h44adb808, 32'h00000000} /* (16, 15, 6) {real, imag} */,
  {32'h449c43ba, 32'h00000000} /* (16, 15, 5) {real, imag} */,
  {32'h4501f8aa, 32'h00000000} /* (16, 15, 4) {real, imag} */,
  {32'h4519b7ce, 32'h00000000} /* (16, 15, 3) {real, imag} */,
  {32'h4510406d, 32'h00000000} /* (16, 15, 2) {real, imag} */,
  {32'h44e93ac3, 32'h00000000} /* (16, 15, 1) {real, imag} */,
  {32'h44975ea8, 32'h00000000} /* (16, 15, 0) {real, imag} */,
  {32'h44899915, 32'h00000000} /* (16, 14, 31) {real, imag} */,
  {32'h44783784, 32'h00000000} /* (16, 14, 30) {real, imag} */,
  {32'h44bfb22c, 32'h00000000} /* (16, 14, 29) {real, imag} */,
  {32'h440bff8d, 32'h00000000} /* (16, 14, 28) {real, imag} */,
  {32'h44ad7050, 32'h00000000} /* (16, 14, 27) {real, imag} */,
  {32'h446c1023, 32'h00000000} /* (16, 14, 26) {real, imag} */,
  {32'h4407308a, 32'h00000000} /* (16, 14, 25) {real, imag} */,
  {32'h4431bc32, 32'h00000000} /* (16, 14, 24) {real, imag} */,
  {32'h44902907, 32'h00000000} /* (16, 14, 23) {real, imag} */,
  {32'h44c61f64, 32'h00000000} /* (16, 14, 22) {real, imag} */,
  {32'h43e570dc, 32'h00000000} /* (16, 14, 21) {real, imag} */,
  {32'hc481a892, 32'h00000000} /* (16, 14, 20) {real, imag} */,
  {32'hc506e148, 32'h00000000} /* (16, 14, 19) {real, imag} */,
  {32'hc48bb260, 32'h00000000} /* (16, 14, 18) {real, imag} */,
  {32'hc42333d9, 32'h00000000} /* (16, 14, 17) {real, imag} */,
  {32'hc49c89f4, 32'h00000000} /* (16, 14, 16) {real, imag} */,
  {32'hc49c1c7f, 32'h00000000} /* (16, 14, 15) {real, imag} */,
  {32'hc4a2c4c2, 32'h00000000} /* (16, 14, 14) {real, imag} */,
  {32'hc4a77e5c, 32'h00000000} /* (16, 14, 13) {real, imag} */,
  {32'hc3e4bb8e, 32'h00000000} /* (16, 14, 12) {real, imag} */,
  {32'h42fc1640, 32'h00000000} /* (16, 14, 11) {real, imag} */,
  {32'h44c76626, 32'h00000000} /* (16, 14, 10) {real, imag} */,
  {32'h4504b184, 32'h00000000} /* (16, 14, 9) {real, imag} */,
  {32'h44f0b0f7, 32'h00000000} /* (16, 14, 8) {real, imag} */,
  {32'h44b75489, 32'h00000000} /* (16, 14, 7) {real, imag} */,
  {32'h44b8818c, 32'h00000000} /* (16, 14, 6) {real, imag} */,
  {32'h44cb1159, 32'h00000000} /* (16, 14, 5) {real, imag} */,
  {32'h44fb1446, 32'h00000000} /* (16, 14, 4) {real, imag} */,
  {32'h45132df4, 32'h00000000} /* (16, 14, 3) {real, imag} */,
  {32'h44cca680, 32'h00000000} /* (16, 14, 2) {real, imag} */,
  {32'h44a905aa, 32'h00000000} /* (16, 14, 1) {real, imag} */,
  {32'h4484b31e, 32'h00000000} /* (16, 14, 0) {real, imag} */,
  {32'h448907ea, 32'h00000000} /* (16, 13, 31) {real, imag} */,
  {32'h44b0078b, 32'h00000000} /* (16, 13, 30) {real, imag} */,
  {32'h44cdde27, 32'h00000000} /* (16, 13, 29) {real, imag} */,
  {32'h44479dba, 32'h00000000} /* (16, 13, 28) {real, imag} */,
  {32'h448b9f8a, 32'h00000000} /* (16, 13, 27) {real, imag} */,
  {32'h44d5fdb6, 32'h00000000} /* (16, 13, 26) {real, imag} */,
  {32'h44a8fea9, 32'h00000000} /* (16, 13, 25) {real, imag} */,
  {32'h44964edd, 32'h00000000} /* (16, 13, 24) {real, imag} */,
  {32'h445d9ad3, 32'h00000000} /* (16, 13, 23) {real, imag} */,
  {32'h442cf734, 32'h00000000} /* (16, 13, 22) {real, imag} */,
  {32'h42a0bd48, 32'h00000000} /* (16, 13, 21) {real, imag} */,
  {32'hc4af8c9c, 32'h00000000} /* (16, 13, 20) {real, imag} */,
  {32'hc4806eb8, 32'h00000000} /* (16, 13, 19) {real, imag} */,
  {32'hc45ead9c, 32'h00000000} /* (16, 13, 18) {real, imag} */,
  {32'hc44547fc, 32'h00000000} /* (16, 13, 17) {real, imag} */,
  {32'hc410f795, 32'h00000000} /* (16, 13, 16) {real, imag} */,
  {32'hc4517517, 32'h00000000} /* (16, 13, 15) {real, imag} */,
  {32'hc48b4e57, 32'h00000000} /* (16, 13, 14) {real, imag} */,
  {32'hc472e1a6, 32'h00000000} /* (16, 13, 13) {real, imag} */,
  {32'hc3a47358, 32'h00000000} /* (16, 13, 12) {real, imag} */,
  {32'hc323c224, 32'h00000000} /* (16, 13, 11) {real, imag} */,
  {32'h44b8899a, 32'h00000000} /* (16, 13, 10) {real, imag} */,
  {32'h44d5894b, 32'h00000000} /* (16, 13, 9) {real, imag} */,
  {32'h4511c66c, 32'h00000000} /* (16, 13, 8) {real, imag} */,
  {32'h450502a7, 32'h00000000} /* (16, 13, 7) {real, imag} */,
  {32'h44af586a, 32'h00000000} /* (16, 13, 6) {real, imag} */,
  {32'h44c9a6d0, 32'h00000000} /* (16, 13, 5) {real, imag} */,
  {32'h4505dc7c, 32'h00000000} /* (16, 13, 4) {real, imag} */,
  {32'h4553a228, 32'h00000000} /* (16, 13, 3) {real, imag} */,
  {32'h450178fd, 32'h00000000} /* (16, 13, 2) {real, imag} */,
  {32'h44ca22ce, 32'h00000000} /* (16, 13, 1) {real, imag} */,
  {32'h444db43b, 32'h00000000} /* (16, 13, 0) {real, imag} */,
  {32'h444cb864, 32'h00000000} /* (16, 12, 31) {real, imag} */,
  {32'h4433bd88, 32'h00000000} /* (16, 12, 30) {real, imag} */,
  {32'h44cbe5a2, 32'h00000000} /* (16, 12, 29) {real, imag} */,
  {32'h4475f2b5, 32'h00000000} /* (16, 12, 28) {real, imag} */,
  {32'h44c4550e, 32'h00000000} /* (16, 12, 27) {real, imag} */,
  {32'h44c15a28, 32'h00000000} /* (16, 12, 26) {real, imag} */,
  {32'h44cd900c, 32'h00000000} /* (16, 12, 25) {real, imag} */,
  {32'h44a63188, 32'h00000000} /* (16, 12, 24) {real, imag} */,
  {32'h4485c0b5, 32'h00000000} /* (16, 12, 23) {real, imag} */,
  {32'h445d42e8, 32'h00000000} /* (16, 12, 22) {real, imag} */,
  {32'h44c0bbf5, 32'h00000000} /* (16, 12, 21) {real, imag} */,
  {32'hc2ae7e20, 32'h00000000} /* (16, 12, 20) {real, imag} */,
  {32'hc493d905, 32'h00000000} /* (16, 12, 19) {real, imag} */,
  {32'hc48a37af, 32'h00000000} /* (16, 12, 18) {real, imag} */,
  {32'hc3c24abc, 32'h00000000} /* (16, 12, 17) {real, imag} */,
  {32'hc45ea319, 32'h00000000} /* (16, 12, 16) {real, imag} */,
  {32'hc4abacf4, 32'h00000000} /* (16, 12, 15) {real, imag} */,
  {32'hc48c8547, 32'h00000000} /* (16, 12, 14) {real, imag} */,
  {32'h42da8798, 32'h00000000} /* (16, 12, 13) {real, imag} */,
  {32'hc325cb54, 32'h00000000} /* (16, 12, 12) {real, imag} */,
  {32'h4458f8df, 32'h00000000} /* (16, 12, 11) {real, imag} */,
  {32'h44d868ce, 32'h00000000} /* (16, 12, 10) {real, imag} */,
  {32'h44f4b738, 32'h00000000} /* (16, 12, 9) {real, imag} */,
  {32'h44cfabd4, 32'h00000000} /* (16, 12, 8) {real, imag} */,
  {32'h44ee8e57, 32'h00000000} /* (16, 12, 7) {real, imag} */,
  {32'h451270d0, 32'h00000000} /* (16, 12, 6) {real, imag} */,
  {32'h44bc6aff, 32'h00000000} /* (16, 12, 5) {real, imag} */,
  {32'h450e9c97, 32'h00000000} /* (16, 12, 4) {real, imag} */,
  {32'h44f2ad19, 32'h00000000} /* (16, 12, 3) {real, imag} */,
  {32'h4532b0a0, 32'h00000000} /* (16, 12, 2) {real, imag} */,
  {32'h45019546, 32'h00000000} /* (16, 12, 1) {real, imag} */,
  {32'h44a7bd2e, 32'h00000000} /* (16, 12, 0) {real, imag} */,
  {32'h440ecc52, 32'h00000000} /* (16, 11, 31) {real, imag} */,
  {32'h44b33ea6, 32'h00000000} /* (16, 11, 30) {real, imag} */,
  {32'h440d2506, 32'h00000000} /* (16, 11, 29) {real, imag} */,
  {32'h446b4f74, 32'h00000000} /* (16, 11, 28) {real, imag} */,
  {32'h44813f0c, 32'h00000000} /* (16, 11, 27) {real, imag} */,
  {32'h42a9ae5c, 32'h00000000} /* (16, 11, 26) {real, imag} */,
  {32'hc3a3f4ce, 32'h00000000} /* (16, 11, 25) {real, imag} */,
  {32'h441d31bc, 32'h00000000} /* (16, 11, 24) {real, imag} */,
  {32'h4426295f, 32'h00000000} /* (16, 11, 23) {real, imag} */,
  {32'h4469099f, 32'h00000000} /* (16, 11, 22) {real, imag} */,
  {32'h44f0f30a, 32'h00000000} /* (16, 11, 21) {real, imag} */,
  {32'hc000f000, 32'h00000000} /* (16, 11, 20) {real, imag} */,
  {32'hc4763582, 32'h00000000} /* (16, 11, 19) {real, imag} */,
  {32'hc37bacd0, 32'h00000000} /* (16, 11, 18) {real, imag} */,
  {32'h43cbaa20, 32'h00000000} /* (16, 11, 17) {real, imag} */,
  {32'hc3123064, 32'h00000000} /* (16, 11, 16) {real, imag} */,
  {32'hc45f9e90, 32'h00000000} /* (16, 11, 15) {real, imag} */,
  {32'h432db3b4, 32'h00000000} /* (16, 11, 14) {real, imag} */,
  {32'h440b4c48, 32'h00000000} /* (16, 11, 13) {real, imag} */,
  {32'h4408ead4, 32'h00000000} /* (16, 11, 12) {real, imag} */,
  {32'h44803d26, 32'h00000000} /* (16, 11, 11) {real, imag} */,
  {32'h44791d22, 32'h00000000} /* (16, 11, 10) {real, imag} */,
  {32'h44d4bdaa, 32'h00000000} /* (16, 11, 9) {real, imag} */,
  {32'h453ae48e, 32'h00000000} /* (16, 11, 8) {real, imag} */,
  {32'h44a44ab0, 32'h00000000} /* (16, 11, 7) {real, imag} */,
  {32'h4524c00e, 32'h00000000} /* (16, 11, 6) {real, imag} */,
  {32'h452a8361, 32'h00000000} /* (16, 11, 5) {real, imag} */,
  {32'h44e80dc0, 32'h00000000} /* (16, 11, 4) {real, imag} */,
  {32'h44a98297, 32'h00000000} /* (16, 11, 3) {real, imag} */,
  {32'h449e0d29, 32'h00000000} /* (16, 11, 2) {real, imag} */,
  {32'h44981b16, 32'h00000000} /* (16, 11, 1) {real, imag} */,
  {32'h44aa8d7a, 32'h00000000} /* (16, 11, 0) {real, imag} */,
  {32'hc450ce74, 32'h00000000} /* (16, 10, 31) {real, imag} */,
  {32'hc397a236, 32'h00000000} /* (16, 10, 30) {real, imag} */,
  {32'h41788940, 32'h00000000} /* (16, 10, 29) {real, imag} */,
  {32'hc3fd5ca2, 32'h00000000} /* (16, 10, 28) {real, imag} */,
  {32'hc4a279fe, 32'h00000000} /* (16, 10, 27) {real, imag} */,
  {32'hc4c1e994, 32'h00000000} /* (16, 10, 26) {real, imag} */,
  {32'hc44a4402, 32'h00000000} /* (16, 10, 25) {real, imag} */,
  {32'hc47e331e, 32'h00000000} /* (16, 10, 24) {real, imag} */,
  {32'hc4136c13, 32'h00000000} /* (16, 10, 23) {real, imag} */,
  {32'hc35c7fac, 32'h00000000} /* (16, 10, 22) {real, imag} */,
  {32'hc3cdd881, 32'h00000000} /* (16, 10, 21) {real, imag} */,
  {32'h43e63bc4, 32'h00000000} /* (16, 10, 20) {real, imag} */,
  {32'h447189b4, 32'h00000000} /* (16, 10, 19) {real, imag} */,
  {32'h44b68776, 32'h00000000} /* (16, 10, 18) {real, imag} */,
  {32'h447efaf6, 32'h00000000} /* (16, 10, 17) {real, imag} */,
  {32'h44ad6759, 32'h00000000} /* (16, 10, 16) {real, imag} */,
  {32'h450f78c8, 32'h00000000} /* (16, 10, 15) {real, imag} */,
  {32'h4466c4a5, 32'h00000000} /* (16, 10, 14) {real, imag} */,
  {32'h449c1d8e, 32'h00000000} /* (16, 10, 13) {real, imag} */,
  {32'h449128f8, 32'h00000000} /* (16, 10, 12) {real, imag} */,
  {32'h4432a070, 32'h00000000} /* (16, 10, 11) {real, imag} */,
  {32'h4431fd55, 32'h00000000} /* (16, 10, 10) {real, imag} */,
  {32'h4357c512, 32'h00000000} /* (16, 10, 9) {real, imag} */,
  {32'h445639b6, 32'h00000000} /* (16, 10, 8) {real, imag} */,
  {32'h43185e28, 32'h00000000} /* (16, 10, 7) {real, imag} */,
  {32'h44a07a00, 32'h00000000} /* (16, 10, 6) {real, imag} */,
  {32'h445f6a68, 32'h00000000} /* (16, 10, 5) {real, imag} */,
  {32'h4337d078, 32'h00000000} /* (16, 10, 4) {real, imag} */,
  {32'h43b2e3b7, 32'h00000000} /* (16, 10, 3) {real, imag} */,
  {32'h4385f26a, 32'h00000000} /* (16, 10, 2) {real, imag} */,
  {32'hc33afe6a, 32'h00000000} /* (16, 10, 1) {real, imag} */,
  {32'h42acb6b0, 32'h00000000} /* (16, 10, 0) {real, imag} */,
  {32'hc49aa6e0, 32'h00000000} /* (16, 9, 31) {real, imag} */,
  {32'hc5030eb8, 32'h00000000} /* (16, 9, 30) {real, imag} */,
  {32'hc4b1da8d, 32'h00000000} /* (16, 9, 29) {real, imag} */,
  {32'hc49c0d6e, 32'h00000000} /* (16, 9, 28) {real, imag} */,
  {32'hc51b53cd, 32'h00000000} /* (16, 9, 27) {real, imag} */,
  {32'hc493c75b, 32'h00000000} /* (16, 9, 26) {real, imag} */,
  {32'hc4ab9dca, 32'h00000000} /* (16, 9, 25) {real, imag} */,
  {32'hc4873b03, 32'h00000000} /* (16, 9, 24) {real, imag} */,
  {32'hc4c120f5, 32'h00000000} /* (16, 9, 23) {real, imag} */,
  {32'hc4dbf3ba, 32'h00000000} /* (16, 9, 22) {real, imag} */,
  {32'hc35214f8, 32'h00000000} /* (16, 9, 21) {real, imag} */,
  {32'h44272177, 32'h00000000} /* (16, 9, 20) {real, imag} */,
  {32'h449e930e, 32'h00000000} /* (16, 9, 19) {real, imag} */,
  {32'h44bc4a26, 32'h00000000} /* (16, 9, 18) {real, imag} */,
  {32'h4516bad8, 32'h00000000} /* (16, 9, 17) {real, imag} */,
  {32'h451fa1ea, 32'h00000000} /* (16, 9, 16) {real, imag} */,
  {32'h454986ba, 32'h00000000} /* (16, 9, 15) {real, imag} */,
  {32'h450b65d2, 32'h00000000} /* (16, 9, 14) {real, imag} */,
  {32'h44bfbc21, 32'h00000000} /* (16, 9, 13) {real, imag} */,
  {32'h44bbf426, 32'h00000000} /* (16, 9, 12) {real, imag} */,
  {32'h44a230b0, 32'h00000000} /* (16, 9, 11) {real, imag} */,
  {32'h43083b40, 32'h00000000} /* (16, 9, 10) {real, imag} */,
  {32'hc3fc194a, 32'h00000000} /* (16, 9, 9) {real, imag} */,
  {32'hc482a38d, 32'h00000000} /* (16, 9, 8) {real, imag} */,
  {32'hc387a13c, 32'h00000000} /* (16, 9, 7) {real, imag} */,
  {32'h42cefe88, 32'h00000000} /* (16, 9, 6) {real, imag} */,
  {32'hc4a014d7, 32'h00000000} /* (16, 9, 5) {real, imag} */,
  {32'hc42ba6bd, 32'h00000000} /* (16, 9, 4) {real, imag} */,
  {32'hc3ecf775, 32'h00000000} /* (16, 9, 3) {real, imag} */,
  {32'hc46bc750, 32'h00000000} /* (16, 9, 2) {real, imag} */,
  {32'hc43fbe6c, 32'h00000000} /* (16, 9, 1) {real, imag} */,
  {32'hc49a3b4a, 32'h00000000} /* (16, 9, 0) {real, imag} */,
  {32'hc4c6eb1b, 32'h00000000} /* (16, 8, 31) {real, imag} */,
  {32'hc4e95e3c, 32'h00000000} /* (16, 8, 30) {real, imag} */,
  {32'hc5080e93, 32'h00000000} /* (16, 8, 29) {real, imag} */,
  {32'hc499c6ba, 32'h00000000} /* (16, 8, 28) {real, imag} */,
  {32'hc4aba6a7, 32'h00000000} /* (16, 8, 27) {real, imag} */,
  {32'hc4f9a8df, 32'h00000000} /* (16, 8, 26) {real, imag} */,
  {32'hc4e7c6c0, 32'h00000000} /* (16, 8, 25) {real, imag} */,
  {32'hc4a1cc70, 32'h00000000} /* (16, 8, 24) {real, imag} */,
  {32'hc4ef4100, 32'h00000000} /* (16, 8, 23) {real, imag} */,
  {32'hc4acb21e, 32'h00000000} /* (16, 8, 22) {real, imag} */,
  {32'hc430b8fb, 32'h00000000} /* (16, 8, 21) {real, imag} */,
  {32'hc38848f6, 32'h00000000} /* (16, 8, 20) {real, imag} */,
  {32'h44e70551, 32'h00000000} /* (16, 8, 19) {real, imag} */,
  {32'h44bfea12, 32'h00000000} /* (16, 8, 18) {real, imag} */,
  {32'h4518c0d6, 32'h00000000} /* (16, 8, 17) {real, imag} */,
  {32'h455209c8, 32'h00000000} /* (16, 8, 16) {real, imag} */,
  {32'h450904ae, 32'h00000000} /* (16, 8, 15) {real, imag} */,
  {32'h452fe8ec, 32'h00000000} /* (16, 8, 14) {real, imag} */,
  {32'h45198d9b, 32'h00000000} /* (16, 8, 13) {real, imag} */,
  {32'h44eaa424, 32'h00000000} /* (16, 8, 12) {real, imag} */,
  {32'h448a04cb, 32'h00000000} /* (16, 8, 11) {real, imag} */,
  {32'hc1f5c9c0, 32'h00000000} /* (16, 8, 10) {real, imag} */,
  {32'hc404d379, 32'h00000000} /* (16, 8, 9) {real, imag} */,
  {32'h42f2d6e0, 32'h00000000} /* (16, 8, 8) {real, imag} */,
  {32'hc3b9e060, 32'h00000000} /* (16, 8, 7) {real, imag} */,
  {32'hc41d3c82, 32'h00000000} /* (16, 8, 6) {real, imag} */,
  {32'hc4e2a82a, 32'h00000000} /* (16, 8, 5) {real, imag} */,
  {32'hc48f439e, 32'h00000000} /* (16, 8, 4) {real, imag} */,
  {32'hc4460742, 32'h00000000} /* (16, 8, 3) {real, imag} */,
  {32'hc4bdaef2, 32'h00000000} /* (16, 8, 2) {real, imag} */,
  {32'hc52e1760, 32'h00000000} /* (16, 8, 1) {real, imag} */,
  {32'hc544b508, 32'h00000000} /* (16, 8, 0) {real, imag} */,
  {32'hc5265164, 32'h00000000} /* (16, 7, 31) {real, imag} */,
  {32'hc53139dc, 32'h00000000} /* (16, 7, 30) {real, imag} */,
  {32'hc5030e5e, 32'h00000000} /* (16, 7, 29) {real, imag} */,
  {32'hc50b41eb, 32'h00000000} /* (16, 7, 28) {real, imag} */,
  {32'hc5094f63, 32'h00000000} /* (16, 7, 27) {real, imag} */,
  {32'hc50bed86, 32'h00000000} /* (16, 7, 26) {real, imag} */,
  {32'hc52fbc3c, 32'h00000000} /* (16, 7, 25) {real, imag} */,
  {32'hc507c21a, 32'h00000000} /* (16, 7, 24) {real, imag} */,
  {32'hc4c8e6c3, 32'h00000000} /* (16, 7, 23) {real, imag} */,
  {32'hc4e8454e, 32'h00000000} /* (16, 7, 22) {real, imag} */,
  {32'hc49c5ef8, 32'h00000000} /* (16, 7, 21) {real, imag} */,
  {32'hc3b8dff4, 32'h00000000} /* (16, 7, 20) {real, imag} */,
  {32'h440713aa, 32'h00000000} /* (16, 7, 19) {real, imag} */,
  {32'h44432fa4, 32'h00000000} /* (16, 7, 18) {real, imag} */,
  {32'h451267fc, 32'h00000000} /* (16, 7, 17) {real, imag} */,
  {32'h44d34c11, 32'h00000000} /* (16, 7, 16) {real, imag} */,
  {32'h449ae503, 32'h00000000} /* (16, 7, 15) {real, imag} */,
  {32'h45358f4a, 32'h00000000} /* (16, 7, 14) {real, imag} */,
  {32'h45412c76, 32'h00000000} /* (16, 7, 13) {real, imag} */,
  {32'h44c83b72, 32'h00000000} /* (16, 7, 12) {real, imag} */,
  {32'h45246fb5, 32'h00000000} /* (16, 7, 11) {real, imag} */,
  {32'hc2b72360, 32'h00000000} /* (16, 7, 10) {real, imag} */,
  {32'hc43a6fce, 32'h00000000} /* (16, 7, 9) {real, imag} */,
  {32'hc3d725a2, 32'h00000000} /* (16, 7, 8) {real, imag} */,
  {32'hc3033a18, 32'h00000000} /* (16, 7, 7) {real, imag} */,
  {32'hc4aa4f82, 32'h00000000} /* (16, 7, 6) {real, imag} */,
  {32'hc48d38cc, 32'h00000000} /* (16, 7, 5) {real, imag} */,
  {32'hc51c87c2, 32'h00000000} /* (16, 7, 4) {real, imag} */,
  {32'hc4d1182b, 32'h00000000} /* (16, 7, 3) {real, imag} */,
  {32'hc512598d, 32'h00000000} /* (16, 7, 2) {real, imag} */,
  {32'hc523329c, 32'h00000000} /* (16, 7, 1) {real, imag} */,
  {32'hc50cc592, 32'h00000000} /* (16, 7, 0) {real, imag} */,
  {32'hc51555e4, 32'h00000000} /* (16, 6, 31) {real, imag} */,
  {32'hc513440b, 32'h00000000} /* (16, 6, 30) {real, imag} */,
  {32'hc5403009, 32'h00000000} /* (16, 6, 29) {real, imag} */,
  {32'hc535ace8, 32'h00000000} /* (16, 6, 28) {real, imag} */,
  {32'hc4f9e2c2, 32'h00000000} /* (16, 6, 27) {real, imag} */,
  {32'hc527a431, 32'h00000000} /* (16, 6, 26) {real, imag} */,
  {32'hc527e730, 32'h00000000} /* (16, 6, 25) {real, imag} */,
  {32'hc4f91d96, 32'h00000000} /* (16, 6, 24) {real, imag} */,
  {32'hc4e870c2, 32'h00000000} /* (16, 6, 23) {real, imag} */,
  {32'hc4efcc24, 32'h00000000} /* (16, 6, 22) {real, imag} */,
  {32'hc4c70780, 32'h00000000} /* (16, 6, 21) {real, imag} */,
  {32'hc296b718, 32'h00000000} /* (16, 6, 20) {real, imag} */,
  {32'h44333851, 32'h00000000} /* (16, 6, 19) {real, imag} */,
  {32'h448422d2, 32'h00000000} /* (16, 6, 18) {real, imag} */,
  {32'h44af805b, 32'h00000000} /* (16, 6, 17) {real, imag} */,
  {32'h44ff8d78, 32'h00000000} /* (16, 6, 16) {real, imag} */,
  {32'h450cd1be, 32'h00000000} /* (16, 6, 15) {real, imag} */,
  {32'h44fc2eae, 32'h00000000} /* (16, 6, 14) {real, imag} */,
  {32'h45278473, 32'h00000000} /* (16, 6, 13) {real, imag} */,
  {32'h44b0851c, 32'h00000000} /* (16, 6, 12) {real, imag} */,
  {32'h450bb2e7, 32'h00000000} /* (16, 6, 11) {real, imag} */,
  {32'h447c85a3, 32'h00000000} /* (16, 6, 10) {real, imag} */,
  {32'hc4514914, 32'h00000000} /* (16, 6, 9) {real, imag} */,
  {32'hc222d710, 32'h00000000} /* (16, 6, 8) {real, imag} */,
  {32'hc3850998, 32'h00000000} /* (16, 6, 7) {real, imag} */,
  {32'hc49194f8, 32'h00000000} /* (16, 6, 6) {real, imag} */,
  {32'hc4456710, 32'h00000000} /* (16, 6, 5) {real, imag} */,
  {32'hc4bb775e, 32'h00000000} /* (16, 6, 4) {real, imag} */,
  {32'hc50ed698, 32'h00000000} /* (16, 6, 3) {real, imag} */,
  {32'hc52a7f5f, 32'h00000000} /* (16, 6, 2) {real, imag} */,
  {32'hc54fc3de, 32'h00000000} /* (16, 6, 1) {real, imag} */,
  {32'hc50a79fc, 32'h00000000} /* (16, 6, 0) {real, imag} */,
  {32'hc5043320, 32'h00000000} /* (16, 5, 31) {real, imag} */,
  {32'hc559cc85, 32'h00000000} /* (16, 5, 30) {real, imag} */,
  {32'hc54059e0, 32'h00000000} /* (16, 5, 29) {real, imag} */,
  {32'hc53a7316, 32'h00000000} /* (16, 5, 28) {real, imag} */,
  {32'hc51015ac, 32'h00000000} /* (16, 5, 27) {real, imag} */,
  {32'hc540c815, 32'h00000000} /* (16, 5, 26) {real, imag} */,
  {32'hc4de495a, 32'h00000000} /* (16, 5, 25) {real, imag} */,
  {32'hc4ddc17b, 32'h00000000} /* (16, 5, 24) {real, imag} */,
  {32'hc5131196, 32'h00000000} /* (16, 5, 23) {real, imag} */,
  {32'hc4e1d87c, 32'h00000000} /* (16, 5, 22) {real, imag} */,
  {32'hc50dfd20, 32'h00000000} /* (16, 5, 21) {real, imag} */,
  {32'hc48436a6, 32'h00000000} /* (16, 5, 20) {real, imag} */,
  {32'h43baee58, 32'h00000000} /* (16, 5, 19) {real, imag} */,
  {32'hc2e21b50, 32'h00000000} /* (16, 5, 18) {real, imag} */,
  {32'h438eeae8, 32'h00000000} /* (16, 5, 17) {real, imag} */,
  {32'h4489a33e, 32'h00000000} /* (16, 5, 16) {real, imag} */,
  {32'h44dcf76f, 32'h00000000} /* (16, 5, 15) {real, imag} */,
  {32'h4520fcd7, 32'h00000000} /* (16, 5, 14) {real, imag} */,
  {32'h450bd77a, 32'h00000000} /* (16, 5, 13) {real, imag} */,
  {32'h45024b9a, 32'h00000000} /* (16, 5, 12) {real, imag} */,
  {32'h448ef4a2, 32'h00000000} /* (16, 5, 11) {real, imag} */,
  {32'h44d52b96, 32'h00000000} /* (16, 5, 10) {real, imag} */,
  {32'h44c1176e, 32'h00000000} /* (16, 5, 9) {real, imag} */,
  {32'h44ab5c07, 32'h00000000} /* (16, 5, 8) {real, imag} */,
  {32'h4454063e, 32'h00000000} /* (16, 5, 7) {real, imag} */,
  {32'h43306ac4, 32'h00000000} /* (16, 5, 6) {real, imag} */,
  {32'hc452abe8, 32'h00000000} /* (16, 5, 5) {real, imag} */,
  {32'hc4c6e2b2, 32'h00000000} /* (16, 5, 4) {real, imag} */,
  {32'hc535f951, 32'h00000000} /* (16, 5, 3) {real, imag} */,
  {32'hc5629254, 32'h00000000} /* (16, 5, 2) {real, imag} */,
  {32'hc54042b3, 32'h00000000} /* (16, 5, 1) {real, imag} */,
  {32'hc5117912, 32'h00000000} /* (16, 5, 0) {real, imag} */,
  {32'hc4f78a73, 32'h00000000} /* (16, 4, 31) {real, imag} */,
  {32'hc52a8b24, 32'h00000000} /* (16, 4, 30) {real, imag} */,
  {32'hc560002c, 32'h00000000} /* (16, 4, 29) {real, imag} */,
  {32'hc5253f38, 32'h00000000} /* (16, 4, 28) {real, imag} */,
  {32'hc5039c5f, 32'h00000000} /* (16, 4, 27) {real, imag} */,
  {32'hc4f929ce, 32'h00000000} /* (16, 4, 26) {real, imag} */,
  {32'hc4ee4ddb, 32'h00000000} /* (16, 4, 25) {real, imag} */,
  {32'hc4e55dda, 32'h00000000} /* (16, 4, 24) {real, imag} */,
  {32'hc4a056e6, 32'h00000000} /* (16, 4, 23) {real, imag} */,
  {32'hc4928063, 32'h00000000} /* (16, 4, 22) {real, imag} */,
  {32'hc4dc1085, 32'h00000000} /* (16, 4, 21) {real, imag} */,
  {32'hc54a7e15, 32'h00000000} /* (16, 4, 20) {real, imag} */,
  {32'hc4c96eea, 32'h00000000} /* (16, 4, 19) {real, imag} */,
  {32'hc43635ac, 32'h00000000} /* (16, 4, 18) {real, imag} */,
  {32'hc43330b6, 32'h00000000} /* (16, 4, 17) {real, imag} */,
  {32'hc47d0aa3, 32'h00000000} /* (16, 4, 16) {real, imag} */,
  {32'h43f5488c, 32'h00000000} /* (16, 4, 15) {real, imag} */,
  {32'h451b628e, 32'h00000000} /* (16, 4, 14) {real, imag} */,
  {32'h4510c940, 32'h00000000} /* (16, 4, 13) {real, imag} */,
  {32'h4502b2f2, 32'h00000000} /* (16, 4, 12) {real, imag} */,
  {32'h451ecda7, 32'h00000000} /* (16, 4, 11) {real, imag} */,
  {32'h44bb5814, 32'h00000000} /* (16, 4, 10) {real, imag} */,
  {32'h450d2508, 32'h00000000} /* (16, 4, 9) {real, imag} */,
  {32'h45122b03, 32'h00000000} /* (16, 4, 8) {real, imag} */,
  {32'h4488f516, 32'h00000000} /* (16, 4, 7) {real, imag} */,
  {32'h44b81071, 32'h00000000} /* (16, 4, 6) {real, imag} */,
  {32'h43a35864, 32'h00000000} /* (16, 4, 5) {real, imag} */,
  {32'hc505c61d, 32'h00000000} /* (16, 4, 4) {real, imag} */,
  {32'hc52c85ab, 32'h00000000} /* (16, 4, 3) {real, imag} */,
  {32'hc53abfad, 32'h00000000} /* (16, 4, 2) {real, imag} */,
  {32'hc509d3fc, 32'h00000000} /* (16, 4, 1) {real, imag} */,
  {32'hc524b905, 32'h00000000} /* (16, 4, 0) {real, imag} */,
  {32'hc5073714, 32'h00000000} /* (16, 3, 31) {real, imag} */,
  {32'hc54622c0, 32'h00000000} /* (16, 3, 30) {real, imag} */,
  {32'hc54c2cbd, 32'h00000000} /* (16, 3, 29) {real, imag} */,
  {32'hc4fa2690, 32'h00000000} /* (16, 3, 28) {real, imag} */,
  {32'hc512144c, 32'h00000000} /* (16, 3, 27) {real, imag} */,
  {32'hc50755bf, 32'h00000000} /* (16, 3, 26) {real, imag} */,
  {32'hc4f965c2, 32'h00000000} /* (16, 3, 25) {real, imag} */,
  {32'hc50e4e0d, 32'h00000000} /* (16, 3, 24) {real, imag} */,
  {32'hc4e3918e, 32'h00000000} /* (16, 3, 23) {real, imag} */,
  {32'hc5095318, 32'h00000000} /* (16, 3, 22) {real, imag} */,
  {32'hc50256be, 32'h00000000} /* (16, 3, 21) {real, imag} */,
  {32'hc500d75b, 32'h00000000} /* (16, 3, 20) {real, imag} */,
  {32'hc4967901, 32'h00000000} /* (16, 3, 19) {real, imag} */,
  {32'hc50f0760, 32'h00000000} /* (16, 3, 18) {real, imag} */,
  {32'hc4995c0c, 32'h00000000} /* (16, 3, 17) {real, imag} */,
  {32'hc3b535a4, 32'h00000000} /* (16, 3, 16) {real, imag} */,
  {32'h4483dfa1, 32'h00000000} /* (16, 3, 15) {real, imag} */,
  {32'h451435ce, 32'h00000000} /* (16, 3, 14) {real, imag} */,
  {32'h44e36256, 32'h00000000} /* (16, 3, 13) {real, imag} */,
  {32'h44fadce2, 32'h00000000} /* (16, 3, 12) {real, imag} */,
  {32'h4519d900, 32'h00000000} /* (16, 3, 11) {real, imag} */,
  {32'h44fff42e, 32'h00000000} /* (16, 3, 10) {real, imag} */,
  {32'h44ddcd96, 32'h00000000} /* (16, 3, 9) {real, imag} */,
  {32'h44f616ae, 32'h00000000} /* (16, 3, 8) {real, imag} */,
  {32'h445b737c, 32'h00000000} /* (16, 3, 7) {real, imag} */,
  {32'h44904bc6, 32'h00000000} /* (16, 3, 6) {real, imag} */,
  {32'hc422cd92, 32'h00000000} /* (16, 3, 5) {real, imag} */,
  {32'hc4acecba, 32'h00000000} /* (16, 3, 4) {real, imag} */,
  {32'hc4980827, 32'h00000000} /* (16, 3, 3) {real, imag} */,
  {32'hc4e08d21, 32'h00000000} /* (16, 3, 2) {real, imag} */,
  {32'hc4e851a4, 32'h00000000} /* (16, 3, 1) {real, imag} */,
  {32'hc4ed2c79, 32'h00000000} /* (16, 3, 0) {real, imag} */,
  {32'hc501cde9, 32'h00000000} /* (16, 2, 31) {real, imag} */,
  {32'hc50620dc, 32'h00000000} /* (16, 2, 30) {real, imag} */,
  {32'hc5053f77, 32'h00000000} /* (16, 2, 29) {real, imag} */,
  {32'hc5206a72, 32'h00000000} /* (16, 2, 28) {real, imag} */,
  {32'hc512b055, 32'h00000000} /* (16, 2, 27) {real, imag} */,
  {32'hc5411a35, 32'h00000000} /* (16, 2, 26) {real, imag} */,
  {32'hc5372eba, 32'h00000000} /* (16, 2, 25) {real, imag} */,
  {32'hc50b7cbf, 32'h00000000} /* (16, 2, 24) {real, imag} */,
  {32'hc4ea8615, 32'h00000000} /* (16, 2, 23) {real, imag} */,
  {32'hc4e0ae66, 32'h00000000} /* (16, 2, 22) {real, imag} */,
  {32'hc514234f, 32'h00000000} /* (16, 2, 21) {real, imag} */,
  {32'hc4aeb9f8, 32'h00000000} /* (16, 2, 20) {real, imag} */,
  {32'hc4f543f5, 32'h00000000} /* (16, 2, 19) {real, imag} */,
  {32'hc5216626, 32'h00000000} /* (16, 2, 18) {real, imag} */,
  {32'hc4fe3b9a, 32'h00000000} /* (16, 2, 17) {real, imag} */,
  {32'h44014ff9, 32'h00000000} /* (16, 2, 16) {real, imag} */,
  {32'h44aa39c6, 32'h00000000} /* (16, 2, 15) {real, imag} */,
  {32'h44f4c0b0, 32'h00000000} /* (16, 2, 14) {real, imag} */,
  {32'h452d7f67, 32'h00000000} /* (16, 2, 13) {real, imag} */,
  {32'h451d8cea, 32'h00000000} /* (16, 2, 12) {real, imag} */,
  {32'h44eb1d56, 32'h00000000} /* (16, 2, 11) {real, imag} */,
  {32'h450011e1, 32'h00000000} /* (16, 2, 10) {real, imag} */,
  {32'h450d6d86, 32'h00000000} /* (16, 2, 9) {real, imag} */,
  {32'h44b47f8a, 32'h00000000} /* (16, 2, 8) {real, imag} */,
  {32'h44688d5e, 32'h00000000} /* (16, 2, 7) {real, imag} */,
  {32'hc392d55a, 32'h00000000} /* (16, 2, 6) {real, imag} */,
  {32'hc445d6a5, 32'h00000000} /* (16, 2, 5) {real, imag} */,
  {32'hc4a66f52, 32'h00000000} /* (16, 2, 4) {real, imag} */,
  {32'hc4ea8dcf, 32'h00000000} /* (16, 2, 3) {real, imag} */,
  {32'hc523b610, 32'h00000000} /* (16, 2, 2) {real, imag} */,
  {32'hc50416df, 32'h00000000} /* (16, 2, 1) {real, imag} */,
  {32'hc4f2ce40, 32'h00000000} /* (16, 2, 0) {real, imag} */,
  {32'hc4c7ff46, 32'h00000000} /* (16, 1, 31) {real, imag} */,
  {32'hc515ff10, 32'h00000000} /* (16, 1, 30) {real, imag} */,
  {32'hc506668e, 32'h00000000} /* (16, 1, 29) {real, imag} */,
  {32'hc5578c6a, 32'h00000000} /* (16, 1, 28) {real, imag} */,
  {32'hc503c76f, 32'h00000000} /* (16, 1, 27) {real, imag} */,
  {32'hc5091627, 32'h00000000} /* (16, 1, 26) {real, imag} */,
  {32'hc50f958e, 32'h00000000} /* (16, 1, 25) {real, imag} */,
  {32'hc52bec66, 32'h00000000} /* (16, 1, 24) {real, imag} */,
  {32'hc4bdfcfc, 32'h00000000} /* (16, 1, 23) {real, imag} */,
  {32'hc51a231f, 32'h00000000} /* (16, 1, 22) {real, imag} */,
  {32'hc4f03bd8, 32'h00000000} /* (16, 1, 21) {real, imag} */,
  {32'hc4ad7fd5, 32'h00000000} /* (16, 1, 20) {real, imag} */,
  {32'hc4ecac34, 32'h00000000} /* (16, 1, 19) {real, imag} */,
  {32'hc4e4dd26, 32'h00000000} /* (16, 1, 18) {real, imag} */,
  {32'hc47977f1, 32'h00000000} /* (16, 1, 17) {real, imag} */,
  {32'h437a7e20, 32'h00000000} /* (16, 1, 16) {real, imag} */,
  {32'h44b00f26, 32'h00000000} /* (16, 1, 15) {real, imag} */,
  {32'h44f203e8, 32'h00000000} /* (16, 1, 14) {real, imag} */,
  {32'h4512a516, 32'h00000000} /* (16, 1, 13) {real, imag} */,
  {32'h453987bc, 32'h00000000} /* (16, 1, 12) {real, imag} */,
  {32'h44c6a284, 32'h00000000} /* (16, 1, 11) {real, imag} */,
  {32'h44c7a032, 32'h00000000} /* (16, 1, 10) {real, imag} */,
  {32'h4455c081, 32'h00000000} /* (16, 1, 9) {real, imag} */,
  {32'h448e4d7e, 32'h00000000} /* (16, 1, 8) {real, imag} */,
  {32'hc3964248, 32'h00000000} /* (16, 1, 7) {real, imag} */,
  {32'hc41e0653, 32'h00000000} /* (16, 1, 6) {real, imag} */,
  {32'hc454bc7d, 32'h00000000} /* (16, 1, 5) {real, imag} */,
  {32'hc4fdec89, 32'h00000000} /* (16, 1, 4) {real, imag} */,
  {32'hc508322c, 32'h00000000} /* (16, 1, 3) {real, imag} */,
  {32'hc5033449, 32'h00000000} /* (16, 1, 2) {real, imag} */,
  {32'hc5086ea2, 32'h00000000} /* (16, 1, 1) {real, imag} */,
  {32'hc525478d, 32'h00000000} /* (16, 1, 0) {real, imag} */,
  {32'hc4efc8de, 32'h00000000} /* (16, 0, 31) {real, imag} */,
  {32'hc5104d7d, 32'h00000000} /* (16, 0, 30) {real, imag} */,
  {32'hc5164f2f, 32'h00000000} /* (16, 0, 29) {real, imag} */,
  {32'hc50802a0, 32'h00000000} /* (16, 0, 28) {real, imag} */,
  {32'hc504353a, 32'h00000000} /* (16, 0, 27) {real, imag} */,
  {32'hc5100b69, 32'h00000000} /* (16, 0, 26) {real, imag} */,
  {32'hc50a4b1a, 32'h00000000} /* (16, 0, 25) {real, imag} */,
  {32'hc527a698, 32'h00000000} /* (16, 0, 24) {real, imag} */,
  {32'hc4ec1934, 32'h00000000} /* (16, 0, 23) {real, imag} */,
  {32'hc5161f25, 32'h00000000} /* (16, 0, 22) {real, imag} */,
  {32'hc4de73dc, 32'h00000000} /* (16, 0, 21) {real, imag} */,
  {32'hc49ef082, 32'h00000000} /* (16, 0, 20) {real, imag} */,
  {32'hc4760eaf, 32'h00000000} /* (16, 0, 19) {real, imag} */,
  {32'hc47fbae5, 32'h00000000} /* (16, 0, 18) {real, imag} */,
  {32'hc2894410, 32'h00000000} /* (16, 0, 17) {real, imag} */,
  {32'h43446c50, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h449347a6, 32'h00000000} /* (16, 0, 15) {real, imag} */,
  {32'h44da624a, 32'h00000000} /* (16, 0, 14) {real, imag} */,
  {32'h44bc3c0e, 32'h00000000} /* (16, 0, 13) {real, imag} */,
  {32'h44cb71d0, 32'h00000000} /* (16, 0, 12) {real, imag} */,
  {32'h450a239a, 32'h00000000} /* (16, 0, 11) {real, imag} */,
  {32'h447e6d48, 32'h00000000} /* (16, 0, 10) {real, imag} */,
  {32'h43888a9c, 32'h00000000} /* (16, 0, 9) {real, imag} */,
  {32'hc3a9d3a0, 32'h00000000} /* (16, 0, 8) {real, imag} */,
  {32'hc3bc08d0, 32'h00000000} /* (16, 0, 7) {real, imag} */,
  {32'hc41e4bd3, 32'h00000000} /* (16, 0, 6) {real, imag} */,
  {32'hc4bfedcc, 32'h00000000} /* (16, 0, 5) {real, imag} */,
  {32'hc503ae5d, 32'h00000000} /* (16, 0, 4) {real, imag} */,
  {32'hc4e64e36, 32'h00000000} /* (16, 0, 3) {real, imag} */,
  {32'hc4f10270, 32'h00000000} /* (16, 0, 2) {real, imag} */,
  {32'hc4fc3ed3, 32'h00000000} /* (16, 0, 1) {real, imag} */,
  {32'hc515ab47, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h44dcbbc6, 32'h00000000} /* (15, 31, 31) {real, imag} */,
  {32'h451ee499, 32'h00000000} /* (15, 31, 30) {real, imag} */,
  {32'h4526d64a, 32'h00000000} /* (15, 31, 29) {real, imag} */,
  {32'h450f1c83, 32'h00000000} /* (15, 31, 28) {real, imag} */,
  {32'h4520fbff, 32'h00000000} /* (15, 31, 27) {real, imag} */,
  {32'h450f8bc6, 32'h00000000} /* (15, 31, 26) {real, imag} */,
  {32'h450cc173, 32'h00000000} /* (15, 31, 25) {real, imag} */,
  {32'h4501069a, 32'h00000000} /* (15, 31, 24) {real, imag} */,
  {32'h451bb670, 32'h00000000} /* (15, 31, 23) {real, imag} */,
  {32'h45023189, 32'h00000000} /* (15, 31, 22) {real, imag} */,
  {32'h44861d9e, 32'h00000000} /* (15, 31, 21) {real, imag} */,
  {32'h42e22b30, 32'h00000000} /* (15, 31, 20) {real, imag} */,
  {32'h417ef4c0, 32'h00000000} /* (15, 31, 19) {real, imag} */,
  {32'hc12c8d80, 32'h00000000} /* (15, 31, 18) {real, imag} */,
  {32'hc4b75234, 32'h00000000} /* (15, 31, 17) {real, imag} */,
  {32'hc46ab414, 32'h00000000} /* (15, 31, 16) {real, imag} */,
  {32'hc4c31092, 32'h00000000} /* (15, 31, 15) {real, imag} */,
  {32'hc4b5e62e, 32'h00000000} /* (15, 31, 14) {real, imag} */,
  {32'hc4cf815c, 32'h00000000} /* (15, 31, 13) {real, imag} */,
  {32'hc4d829fc, 32'h00000000} /* (15, 31, 12) {real, imag} */,
  {32'hc49da52a, 32'h00000000} /* (15, 31, 11) {real, imag} */,
  {32'hc42cd2b0, 32'h00000000} /* (15, 31, 10) {real, imag} */,
  {32'hc3068cf0, 32'h00000000} /* (15, 31, 9) {real, imag} */,
  {32'h42c7f010, 32'h00000000} /* (15, 31, 8) {real, imag} */,
  {32'h43335098, 32'h00000000} /* (15, 31, 7) {real, imag} */,
  {32'h44d897ca, 32'h00000000} /* (15, 31, 6) {real, imag} */,
  {32'h44adef3a, 32'h00000000} /* (15, 31, 5) {real, imag} */,
  {32'h4497562c, 32'h00000000} /* (15, 31, 4) {real, imag} */,
  {32'h44ddb426, 32'h00000000} /* (15, 31, 3) {real, imag} */,
  {32'h4500ffcc, 32'h00000000} /* (15, 31, 2) {real, imag} */,
  {32'h450698f2, 32'h00000000} /* (15, 31, 1) {real, imag} */,
  {32'h44cae17e, 32'h00000000} /* (15, 31, 0) {real, imag} */,
  {32'h44cc994a, 32'h00000000} /* (15, 30, 31) {real, imag} */,
  {32'h4508e6e2, 32'h00000000} /* (15, 30, 30) {real, imag} */,
  {32'h44d01e63, 32'h00000000} /* (15, 30, 29) {real, imag} */,
  {32'h45115e96, 32'h00000000} /* (15, 30, 28) {real, imag} */,
  {32'h451ba5f2, 32'h00000000} /* (15, 30, 27) {real, imag} */,
  {32'h44fbbd72, 32'h00000000} /* (15, 30, 26) {real, imag} */,
  {32'h45347132, 32'h00000000} /* (15, 30, 25) {real, imag} */,
  {32'h451cc18c, 32'h00000000} /* (15, 30, 24) {real, imag} */,
  {32'h452fe9cc, 32'h00000000} /* (15, 30, 23) {real, imag} */,
  {32'h45279d24, 32'h00000000} /* (15, 30, 22) {real, imag} */,
  {32'h4494e8d6, 32'h00000000} /* (15, 30, 21) {real, imag} */,
  {32'h438a1a54, 32'h00000000} /* (15, 30, 20) {real, imag} */,
  {32'h4213ac70, 32'h00000000} /* (15, 30, 19) {real, imag} */,
  {32'hc43b19ce, 32'h00000000} /* (15, 30, 18) {real, imag} */,
  {32'hc4dfee89, 32'h00000000} /* (15, 30, 17) {real, imag} */,
  {32'hc4d86cec, 32'h00000000} /* (15, 30, 16) {real, imag} */,
  {32'hc4420a6b, 32'h00000000} /* (15, 30, 15) {real, imag} */,
  {32'hc468d993, 32'h00000000} /* (15, 30, 14) {real, imag} */,
  {32'hc4acb135, 32'h00000000} /* (15, 30, 13) {real, imag} */,
  {32'hc50fbbea, 32'h00000000} /* (15, 30, 12) {real, imag} */,
  {32'hc3cbfdd0, 32'h00000000} /* (15, 30, 11) {real, imag} */,
  {32'h40842180, 32'h00000000} /* (15, 30, 10) {real, imag} */,
  {32'h433d0378, 32'h00000000} /* (15, 30, 9) {real, imag} */,
  {32'h448afaf8, 32'h00000000} /* (15, 30, 8) {real, imag} */,
  {32'h43b395fc, 32'h00000000} /* (15, 30, 7) {real, imag} */,
  {32'h44dfa1ed, 32'h00000000} /* (15, 30, 6) {real, imag} */,
  {32'h4533891a, 32'h00000000} /* (15, 30, 5) {real, imag} */,
  {32'h4460f106, 32'h00000000} /* (15, 30, 4) {real, imag} */,
  {32'h44a2daa0, 32'h00000000} /* (15, 30, 3) {real, imag} */,
  {32'h44d35e25, 32'h00000000} /* (15, 30, 2) {real, imag} */,
  {32'h45454c60, 32'h00000000} /* (15, 30, 1) {real, imag} */,
  {32'h4521cc3a, 32'h00000000} /* (15, 30, 0) {real, imag} */,
  {32'h44bfb591, 32'h00000000} /* (15, 29, 31) {real, imag} */,
  {32'h44eb92bb, 32'h00000000} /* (15, 29, 30) {real, imag} */,
  {32'h448eebe6, 32'h00000000} /* (15, 29, 29) {real, imag} */,
  {32'h45315f53, 32'h00000000} /* (15, 29, 28) {real, imag} */,
  {32'h45474970, 32'h00000000} /* (15, 29, 27) {real, imag} */,
  {32'h450096e5, 32'h00000000} /* (15, 29, 26) {real, imag} */,
  {32'h451aca9e, 32'h00000000} /* (15, 29, 25) {real, imag} */,
  {32'h4530a2d8, 32'h00000000} /* (15, 29, 24) {real, imag} */,
  {32'h450bb0a6, 32'h00000000} /* (15, 29, 23) {real, imag} */,
  {32'h45205964, 32'h00000000} /* (15, 29, 22) {real, imag} */,
  {32'h450a119b, 32'h00000000} /* (15, 29, 21) {real, imag} */,
  {32'h44417d06, 32'h00000000} /* (15, 29, 20) {real, imag} */,
  {32'hc236c2a0, 32'h00000000} /* (15, 29, 19) {real, imag} */,
  {32'hc413e97f, 32'h00000000} /* (15, 29, 18) {real, imag} */,
  {32'hc4444c7a, 32'h00000000} /* (15, 29, 17) {real, imag} */,
  {32'hc4e5e1bf, 32'h00000000} /* (15, 29, 16) {real, imag} */,
  {32'hc49d2bdb, 32'h00000000} /* (15, 29, 15) {real, imag} */,
  {32'hc4a01d8f, 32'h00000000} /* (15, 29, 14) {real, imag} */,
  {32'hc403b573, 32'h00000000} /* (15, 29, 13) {real, imag} */,
  {32'hc382fbb8, 32'h00000000} /* (15, 29, 12) {real, imag} */,
  {32'hc37318e8, 32'h00000000} /* (15, 29, 11) {real, imag} */,
  {32'h43a7f6ca, 32'h00000000} /* (15, 29, 10) {real, imag} */,
  {32'h44688a14, 32'h00000000} /* (15, 29, 9) {real, imag} */,
  {32'h440a67f6, 32'h00000000} /* (15, 29, 8) {real, imag} */,
  {32'h44a9ba12, 32'h00000000} /* (15, 29, 7) {real, imag} */,
  {32'h44999540, 32'h00000000} /* (15, 29, 6) {real, imag} */,
  {32'h4527b73b, 32'h00000000} /* (15, 29, 5) {real, imag} */,
  {32'h44e15ae1, 32'h00000000} /* (15, 29, 4) {real, imag} */,
  {32'h4428666c, 32'h00000000} /* (15, 29, 3) {real, imag} */,
  {32'h446ada29, 32'h00000000} /* (15, 29, 2) {real, imag} */,
  {32'h44c28347, 32'h00000000} /* (15, 29, 1) {real, imag} */,
  {32'h45047f9c, 32'h00000000} /* (15, 29, 0) {real, imag} */,
  {32'h44c352cd, 32'h00000000} /* (15, 28, 31) {real, imag} */,
  {32'h44e8b5c0, 32'h00000000} /* (15, 28, 30) {real, imag} */,
  {32'h44f5eb52, 32'h00000000} /* (15, 28, 29) {real, imag} */,
  {32'h452fd3c2, 32'h00000000} /* (15, 28, 28) {real, imag} */,
  {32'h452d3300, 32'h00000000} /* (15, 28, 27) {real, imag} */,
  {32'h452ea2b2, 32'h00000000} /* (15, 28, 26) {real, imag} */,
  {32'h450eed1c, 32'h00000000} /* (15, 28, 25) {real, imag} */,
  {32'h45047d4b, 32'h00000000} /* (15, 28, 24) {real, imag} */,
  {32'h453f89a7, 32'h00000000} /* (15, 28, 23) {real, imag} */,
  {32'h454e18f9, 32'h00000000} /* (15, 28, 22) {real, imag} */,
  {32'h44ea3e62, 32'h00000000} /* (15, 28, 21) {real, imag} */,
  {32'h42f49ff8, 32'h00000000} /* (15, 28, 20) {real, imag} */,
  {32'hc404dab2, 32'h00000000} /* (15, 28, 19) {real, imag} */,
  {32'hc39e4596, 32'h00000000} /* (15, 28, 18) {real, imag} */,
  {32'hc4494d93, 32'h00000000} /* (15, 28, 17) {real, imag} */,
  {32'hc47a849b, 32'h00000000} /* (15, 28, 16) {real, imag} */,
  {32'hc3ebcd1c, 32'h00000000} /* (15, 28, 15) {real, imag} */,
  {32'hc4034b6f, 32'h00000000} /* (15, 28, 14) {real, imag} */,
  {32'hc3318640, 32'h00000000} /* (15, 28, 13) {real, imag} */,
  {32'hc350dd48, 32'h00000000} /* (15, 28, 12) {real, imag} */,
  {32'h438c0d14, 32'h00000000} /* (15, 28, 11) {real, imag} */,
  {32'h449ebd9c, 32'h00000000} /* (15, 28, 10) {real, imag} */,
  {32'h443e987e, 32'h00000000} /* (15, 28, 9) {real, imag} */,
  {32'h450065f3, 32'h00000000} /* (15, 28, 8) {real, imag} */,
  {32'h4487a452, 32'h00000000} /* (15, 28, 7) {real, imag} */,
  {32'h44a4670e, 32'h00000000} /* (15, 28, 6) {real, imag} */,
  {32'h44c34c5c, 32'h00000000} /* (15, 28, 5) {real, imag} */,
  {32'h4491d13e, 32'h00000000} /* (15, 28, 4) {real, imag} */,
  {32'h44930e2d, 32'h00000000} /* (15, 28, 3) {real, imag} */,
  {32'h429edf4a, 32'h00000000} /* (15, 28, 2) {real, imag} */,
  {32'h448266ba, 32'h00000000} /* (15, 28, 1) {real, imag} */,
  {32'h44d2fdb0, 32'h00000000} /* (15, 28, 0) {real, imag} */,
  {32'h44c2f3a7, 32'h00000000} /* (15, 27, 31) {real, imag} */,
  {32'h451581f4, 32'h00000000} /* (15, 27, 30) {real, imag} */,
  {32'h44f90d82, 32'h00000000} /* (15, 27, 29) {real, imag} */,
  {32'h45021888, 32'h00000000} /* (15, 27, 28) {real, imag} */,
  {32'h44ea0b20, 32'h00000000} /* (15, 27, 27) {real, imag} */,
  {32'h4529446a, 32'h00000000} /* (15, 27, 26) {real, imag} */,
  {32'h45517a86, 32'h00000000} /* (15, 27, 25) {real, imag} */,
  {32'h4504509b, 32'h00000000} /* (15, 27, 24) {real, imag} */,
  {32'h44ec6604, 32'h00000000} /* (15, 27, 23) {real, imag} */,
  {32'h44fc2eb1, 32'h00000000} /* (15, 27, 22) {real, imag} */,
  {32'h453fb9c2, 32'h00000000} /* (15, 27, 21) {real, imag} */,
  {32'hc3889483, 32'h00000000} /* (15, 27, 20) {real, imag} */,
  {32'hc47abcf2, 32'h00000000} /* (15, 27, 19) {real, imag} */,
  {32'hc44b6872, 32'h00000000} /* (15, 27, 18) {real, imag} */,
  {32'hc4c71924, 32'h00000000} /* (15, 27, 17) {real, imag} */,
  {32'hc4ee3d20, 32'h00000000} /* (15, 27, 16) {real, imag} */,
  {32'hc5033c9c, 32'h00000000} /* (15, 27, 15) {real, imag} */,
  {32'hc40f46e6, 32'h00000000} /* (15, 27, 14) {real, imag} */,
  {32'hc441b9ac, 32'h00000000} /* (15, 27, 13) {real, imag} */,
  {32'hc3dae15c, 32'h00000000} /* (15, 27, 12) {real, imag} */,
  {32'h42759310, 32'h00000000} /* (15, 27, 11) {real, imag} */,
  {32'h449e9fa0, 32'h00000000} /* (15, 27, 10) {real, imag} */,
  {32'h44b02e5c, 32'h00000000} /* (15, 27, 9) {real, imag} */,
  {32'h449bd2de, 32'h00000000} /* (15, 27, 8) {real, imag} */,
  {32'h449aee72, 32'h00000000} /* (15, 27, 7) {real, imag} */,
  {32'h44e820bb, 32'h00000000} /* (15, 27, 6) {real, imag} */,
  {32'h451fefd8, 32'h00000000} /* (15, 27, 5) {real, imag} */,
  {32'h44926ea8, 32'h00000000} /* (15, 27, 4) {real, imag} */,
  {32'h445841d4, 32'h00000000} /* (15, 27, 3) {real, imag} */,
  {32'h44805c1e, 32'h00000000} /* (15, 27, 2) {real, imag} */,
  {32'h4480f1dc, 32'h00000000} /* (15, 27, 1) {real, imag} */,
  {32'h449e1b00, 32'h00000000} /* (15, 27, 0) {real, imag} */,
  {32'h4486cdab, 32'h00000000} /* (15, 26, 31) {real, imag} */,
  {32'h44fe0c33, 32'h00000000} /* (15, 26, 30) {real, imag} */,
  {32'h450e1da5, 32'h00000000} /* (15, 26, 29) {real, imag} */,
  {32'h45220552, 32'h00000000} /* (15, 26, 28) {real, imag} */,
  {32'h450f70c8, 32'h00000000} /* (15, 26, 27) {real, imag} */,
  {32'h450bd482, 32'h00000000} /* (15, 26, 26) {real, imag} */,
  {32'h450ee919, 32'h00000000} /* (15, 26, 25) {real, imag} */,
  {32'h4484e965, 32'h00000000} /* (15, 26, 24) {real, imag} */,
  {32'h44beef7c, 32'h00000000} /* (15, 26, 23) {real, imag} */,
  {32'h44cfe704, 32'h00000000} /* (15, 26, 22) {real, imag} */,
  {32'h44efa739, 32'h00000000} /* (15, 26, 21) {real, imag} */,
  {32'hc3ebd332, 32'h00000000} /* (15, 26, 20) {real, imag} */,
  {32'hc464fcd6, 32'h00000000} /* (15, 26, 19) {real, imag} */,
  {32'hc4bceb58, 32'h00000000} /* (15, 26, 18) {real, imag} */,
  {32'hc5468de2, 32'h00000000} /* (15, 26, 17) {real, imag} */,
  {32'hc51fe566, 32'h00000000} /* (15, 26, 16) {real, imag} */,
  {32'hc4906a77, 32'h00000000} /* (15, 26, 15) {real, imag} */,
  {32'hc4a1c3c9, 32'h00000000} /* (15, 26, 14) {real, imag} */,
  {32'hc4a54b78, 32'h00000000} /* (15, 26, 13) {real, imag} */,
  {32'hc47cb45e, 32'h00000000} /* (15, 26, 12) {real, imag} */,
  {32'hc465993c, 32'h00000000} /* (15, 26, 11) {real, imag} */,
  {32'h446c845a, 32'h00000000} /* (15, 26, 10) {real, imag} */,
  {32'h44937f5c, 32'h00000000} /* (15, 26, 9) {real, imag} */,
  {32'h44156d57, 32'h00000000} /* (15, 26, 8) {real, imag} */,
  {32'h45037e3e, 32'h00000000} /* (15, 26, 7) {real, imag} */,
  {32'h44f454b6, 32'h00000000} /* (15, 26, 6) {real, imag} */,
  {32'h44c2f947, 32'h00000000} /* (15, 26, 5) {real, imag} */,
  {32'h44b0eba4, 32'h00000000} /* (15, 26, 4) {real, imag} */,
  {32'h450fd178, 32'h00000000} /* (15, 26, 3) {real, imag} */,
  {32'h44f1d9f6, 32'h00000000} /* (15, 26, 2) {real, imag} */,
  {32'h4443d9d2, 32'h00000000} /* (15, 26, 1) {real, imag} */,
  {32'h44ac3418, 32'h00000000} /* (15, 26, 0) {real, imag} */,
  {32'h44a5342b, 32'h00000000} /* (15, 25, 31) {real, imag} */,
  {32'h44bc410d, 32'h00000000} /* (15, 25, 30) {real, imag} */,
  {32'h45025371, 32'h00000000} /* (15, 25, 29) {real, imag} */,
  {32'h4520a0e9, 32'h00000000} /* (15, 25, 28) {real, imag} */,
  {32'h4505f5fc, 32'h00000000} /* (15, 25, 27) {real, imag} */,
  {32'h450ac548, 32'h00000000} /* (15, 25, 26) {real, imag} */,
  {32'h44c230ba, 32'h00000000} /* (15, 25, 25) {real, imag} */,
  {32'h44bbc4ee, 32'h00000000} /* (15, 25, 24) {real, imag} */,
  {32'h44d95b1f, 32'h00000000} /* (15, 25, 23) {real, imag} */,
  {32'h44c6be3e, 32'h00000000} /* (15, 25, 22) {real, imag} */,
  {32'h44983ffd, 32'h00000000} /* (15, 25, 21) {real, imag} */,
  {32'h415722c0, 32'h00000000} /* (15, 25, 20) {real, imag} */,
  {32'hc45a8bbd, 32'h00000000} /* (15, 25, 19) {real, imag} */,
  {32'hc4ea7fc2, 32'h00000000} /* (15, 25, 18) {real, imag} */,
  {32'hc4e44d5e, 32'h00000000} /* (15, 25, 17) {real, imag} */,
  {32'hc518fbc5, 32'h00000000} /* (15, 25, 16) {real, imag} */,
  {32'hc501562e, 32'h00000000} /* (15, 25, 15) {real, imag} */,
  {32'hc4b2db0f, 32'h00000000} /* (15, 25, 14) {real, imag} */,
  {32'hc514732f, 32'h00000000} /* (15, 25, 13) {real, imag} */,
  {32'hc4bd45fe, 32'h00000000} /* (15, 25, 12) {real, imag} */,
  {32'hc13b2c00, 32'h00000000} /* (15, 25, 11) {real, imag} */,
  {32'h44273999, 32'h00000000} /* (15, 25, 10) {real, imag} */,
  {32'h446266a4, 32'h00000000} /* (15, 25, 9) {real, imag} */,
  {32'h45008caf, 32'h00000000} /* (15, 25, 8) {real, imag} */,
  {32'h44ddf8f9, 32'h00000000} /* (15, 25, 7) {real, imag} */,
  {32'h44ee15f8, 32'h00000000} /* (15, 25, 6) {real, imag} */,
  {32'h44e5d143, 32'h00000000} /* (15, 25, 5) {real, imag} */,
  {32'h44dd42e8, 32'h00000000} /* (15, 25, 4) {real, imag} */,
  {32'h44c3c878, 32'h00000000} /* (15, 25, 3) {real, imag} */,
  {32'h449cd94e, 32'h00000000} /* (15, 25, 2) {real, imag} */,
  {32'h451d7f4b, 32'h00000000} /* (15, 25, 1) {real, imag} */,
  {32'h44d403da, 32'h00000000} /* (15, 25, 0) {real, imag} */,
  {32'h44b1e162, 32'h00000000} /* (15, 24, 31) {real, imag} */,
  {32'h45045bfc, 32'h00000000} /* (15, 24, 30) {real, imag} */,
  {32'h450e8756, 32'h00000000} /* (15, 24, 29) {real, imag} */,
  {32'h451f74d6, 32'h00000000} /* (15, 24, 28) {real, imag} */,
  {32'h44de5d58, 32'h00000000} /* (15, 24, 27) {real, imag} */,
  {32'h4467a317, 32'h00000000} /* (15, 24, 26) {real, imag} */,
  {32'h4466999b, 32'h00000000} /* (15, 24, 25) {real, imag} */,
  {32'h44d54db8, 32'h00000000} /* (15, 24, 24) {real, imag} */,
  {32'h45069784, 32'h00000000} /* (15, 24, 23) {real, imag} */,
  {32'h44cba839, 32'h00000000} /* (15, 24, 22) {real, imag} */,
  {32'h4440fa5f, 32'h00000000} /* (15, 24, 21) {real, imag} */,
  {32'hc2c190e0, 32'h00000000} /* (15, 24, 20) {real, imag} */,
  {32'hc4719004, 32'h00000000} /* (15, 24, 19) {real, imag} */,
  {32'hc46ead4a, 32'h00000000} /* (15, 24, 18) {real, imag} */,
  {32'hc4c21d11, 32'h00000000} /* (15, 24, 17) {real, imag} */,
  {32'hc51264d4, 32'h00000000} /* (15, 24, 16) {real, imag} */,
  {32'hc50cb5c2, 32'h00000000} /* (15, 24, 15) {real, imag} */,
  {32'hc5149e22, 32'h00000000} /* (15, 24, 14) {real, imag} */,
  {32'hc4d0d523, 32'h00000000} /* (15, 24, 13) {real, imag} */,
  {32'hc40272ea, 32'h00000000} /* (15, 24, 12) {real, imag} */,
  {32'hc4da33c8, 32'h00000000} /* (15, 24, 11) {real, imag} */,
  {32'hc2e3a758, 32'h00000000} /* (15, 24, 10) {real, imag} */,
  {32'h448517f8, 32'h00000000} /* (15, 24, 9) {real, imag} */,
  {32'h44d896ec, 32'h00000000} /* (15, 24, 8) {real, imag} */,
  {32'h44c54de7, 32'h00000000} /* (15, 24, 7) {real, imag} */,
  {32'h44f2f05f, 32'h00000000} /* (15, 24, 6) {real, imag} */,
  {32'h44d7ab28, 32'h00000000} /* (15, 24, 5) {real, imag} */,
  {32'h44a12362, 32'h00000000} /* (15, 24, 4) {real, imag} */,
  {32'h44ae1002, 32'h00000000} /* (15, 24, 3) {real, imag} */,
  {32'h44a4eb45, 32'h00000000} /* (15, 24, 2) {real, imag} */,
  {32'h44b79ba5, 32'h00000000} /* (15, 24, 1) {real, imag} */,
  {32'h44ab419c, 32'h00000000} /* (15, 24, 0) {real, imag} */,
  {32'h4493ca60, 32'h00000000} /* (15, 23, 31) {real, imag} */,
  {32'h4504adbc, 32'h00000000} /* (15, 23, 30) {real, imag} */,
  {32'h4546c6af, 32'h00000000} /* (15, 23, 29) {real, imag} */,
  {32'h44ed2732, 32'h00000000} /* (15, 23, 28) {real, imag} */,
  {32'h447952cf, 32'h00000000} /* (15, 23, 27) {real, imag} */,
  {32'h44447792, 32'h00000000} /* (15, 23, 26) {real, imag} */,
  {32'h44028b6e, 32'h00000000} /* (15, 23, 25) {real, imag} */,
  {32'h4491799b, 32'h00000000} /* (15, 23, 24) {real, imag} */,
  {32'h44765748, 32'h00000000} /* (15, 23, 23) {real, imag} */,
  {32'h4426a848, 32'h00000000} /* (15, 23, 22) {real, imag} */,
  {32'h44667934, 32'h00000000} /* (15, 23, 21) {real, imag} */,
  {32'hc393b010, 32'h00000000} /* (15, 23, 20) {real, imag} */,
  {32'hc452a392, 32'h00000000} /* (15, 23, 19) {real, imag} */,
  {32'hc486857d, 32'h00000000} /* (15, 23, 18) {real, imag} */,
  {32'hc4f15cc0, 32'h00000000} /* (15, 23, 17) {real, imag} */,
  {32'hc50fb979, 32'h00000000} /* (15, 23, 16) {real, imag} */,
  {32'hc4f7509a, 32'h00000000} /* (15, 23, 15) {real, imag} */,
  {32'hc4aaed46, 32'h00000000} /* (15, 23, 14) {real, imag} */,
  {32'hc4b83b3e, 32'h00000000} /* (15, 23, 13) {real, imag} */,
  {32'hc50c0533, 32'h00000000} /* (15, 23, 12) {real, imag} */,
  {32'hc49bb0ca, 32'h00000000} /* (15, 23, 11) {real, imag} */,
  {32'hc33b9086, 32'h00000000} /* (15, 23, 10) {real, imag} */,
  {32'h44a733c6, 32'h00000000} /* (15, 23, 9) {real, imag} */,
  {32'h44593d28, 32'h00000000} /* (15, 23, 8) {real, imag} */,
  {32'h450c3eae, 32'h00000000} /* (15, 23, 7) {real, imag} */,
  {32'h448b3402, 32'h00000000} /* (15, 23, 6) {real, imag} */,
  {32'h45278f23, 32'h00000000} /* (15, 23, 5) {real, imag} */,
  {32'h44cda4b3, 32'h00000000} /* (15, 23, 4) {real, imag} */,
  {32'h446e842a, 32'h00000000} /* (15, 23, 3) {real, imag} */,
  {32'h439ba197, 32'h00000000} /* (15, 23, 2) {real, imag} */,
  {32'h434e1e64, 32'h00000000} /* (15, 23, 1) {real, imag} */,
  {32'h43e46e06, 32'h00000000} /* (15, 23, 0) {real, imag} */,
  {32'h44ded202, 32'h00000000} /* (15, 22, 31) {real, imag} */,
  {32'h44f52769, 32'h00000000} /* (15, 22, 30) {real, imag} */,
  {32'h44e5f840, 32'h00000000} /* (15, 22, 29) {real, imag} */,
  {32'h44e20de5, 32'h00000000} /* (15, 22, 28) {real, imag} */,
  {32'h4420ddd1, 32'h00000000} /* (15, 22, 27) {real, imag} */,
  {32'h42a96c68, 32'h00000000} /* (15, 22, 26) {real, imag} */,
  {32'h436b94a2, 32'h00000000} /* (15, 22, 25) {real, imag} */,
  {32'h444e8c4c, 32'h00000000} /* (15, 22, 24) {real, imag} */,
  {32'h4450be1d, 32'h00000000} /* (15, 22, 23) {real, imag} */,
  {32'h43f11cfb, 32'h00000000} /* (15, 22, 22) {real, imag} */,
  {32'h43780240, 32'h00000000} /* (15, 22, 21) {real, imag} */,
  {32'h42b520d8, 32'h00000000} /* (15, 22, 20) {real, imag} */,
  {32'hc405bf34, 32'h00000000} /* (15, 22, 19) {real, imag} */,
  {32'hc44edfd7, 32'h00000000} /* (15, 22, 18) {real, imag} */,
  {32'hc4d74e40, 32'h00000000} /* (15, 22, 17) {real, imag} */,
  {32'hc5230df2, 32'h00000000} /* (15, 22, 16) {real, imag} */,
  {32'hc4b86a38, 32'h00000000} /* (15, 22, 15) {real, imag} */,
  {32'hc483a1cb, 32'h00000000} /* (15, 22, 14) {real, imag} */,
  {32'hc4993824, 32'h00000000} /* (15, 22, 13) {real, imag} */,
  {32'hc4ba2259, 32'h00000000} /* (15, 22, 12) {real, imag} */,
  {32'hc4bec4a6, 32'h00000000} /* (15, 22, 11) {real, imag} */,
  {32'h424f5790, 32'h00000000} /* (15, 22, 10) {real, imag} */,
  {32'h43f855d3, 32'h00000000} /* (15, 22, 9) {real, imag} */,
  {32'h44ded85e, 32'h00000000} /* (15, 22, 8) {real, imag} */,
  {32'h44256907, 32'h00000000} /* (15, 22, 7) {real, imag} */,
  {32'h44731d06, 32'h00000000} /* (15, 22, 6) {real, imag} */,
  {32'h44c2a496, 32'h00000000} /* (15, 22, 5) {real, imag} */,
  {32'h44c1c070, 32'h00000000} /* (15, 22, 4) {real, imag} */,
  {32'h440b94e0, 32'h00000000} /* (15, 22, 3) {real, imag} */,
  {32'h444edb07, 32'h00000000} /* (15, 22, 2) {real, imag} */,
  {32'h441f32db, 32'h00000000} /* (15, 22, 1) {real, imag} */,
  {32'h43960024, 32'h00000000} /* (15, 22, 0) {real, imag} */,
  {32'h437cc676, 32'h00000000} /* (15, 21, 31) {real, imag} */,
  {32'h4499de22, 32'h00000000} /* (15, 21, 30) {real, imag} */,
  {32'h432e19f0, 32'h00000000} /* (15, 21, 29) {real, imag} */,
  {32'h43118c90, 32'h00000000} /* (15, 21, 28) {real, imag} */,
  {32'h4303c892, 32'h00000000} /* (15, 21, 27) {real, imag} */,
  {32'hc3e6c528, 32'h00000000} /* (15, 21, 26) {real, imag} */,
  {32'hc42e9f5e, 32'h00000000} /* (15, 21, 25) {real, imag} */,
  {32'h439891a7, 32'h00000000} /* (15, 21, 24) {real, imag} */,
  {32'h43e49bff, 32'h00000000} /* (15, 21, 23) {real, imag} */,
  {32'h44514a6c, 32'h00000000} /* (15, 21, 22) {real, imag} */,
  {32'h443c1a05, 32'h00000000} /* (15, 21, 21) {real, imag} */,
  {32'hc32ebe16, 32'h00000000} /* (15, 21, 20) {real, imag} */,
  {32'hc10d3718, 32'h00000000} /* (15, 21, 19) {real, imag} */,
  {32'hc3e4ec69, 32'h00000000} /* (15, 21, 18) {real, imag} */,
  {32'hc3de947c, 32'h00000000} /* (15, 21, 17) {real, imag} */,
  {32'hc46b99f6, 32'h00000000} /* (15, 21, 16) {real, imag} */,
  {32'hc2cf2044, 32'h00000000} /* (15, 21, 15) {real, imag} */,
  {32'hc42d52fc, 32'h00000000} /* (15, 21, 14) {real, imag} */,
  {32'hc46959a4, 32'h00000000} /* (15, 21, 13) {real, imag} */,
  {32'hc484368e, 32'h00000000} /* (15, 21, 12) {real, imag} */,
  {32'hc427beae, 32'h00000000} /* (15, 21, 11) {real, imag} */,
  {32'hc3299621, 32'h00000000} /* (15, 21, 10) {real, imag} */,
  {32'h43ee0c6c, 32'h00000000} /* (15, 21, 9) {real, imag} */,
  {32'hc3bfea4d, 32'h00000000} /* (15, 21, 8) {real, imag} */,
  {32'h43d31403, 32'h00000000} /* (15, 21, 7) {real, imag} */,
  {32'h44608484, 32'h00000000} /* (15, 21, 6) {real, imag} */,
  {32'h4208f210, 32'h00000000} /* (15, 21, 5) {real, imag} */,
  {32'h4406ee2e, 32'h00000000} /* (15, 21, 4) {real, imag} */,
  {32'h4337fa54, 32'h00000000} /* (15, 21, 3) {real, imag} */,
  {32'hc408638e, 32'h00000000} /* (15, 21, 2) {real, imag} */,
  {32'h41d14cb8, 32'h00000000} /* (15, 21, 1) {real, imag} */,
  {32'h440f54c4, 32'h00000000} /* (15, 21, 0) {real, imag} */,
  {32'h41d857e0, 32'h00000000} /* (15, 20, 31) {real, imag} */,
  {32'hc433533f, 32'h00000000} /* (15, 20, 30) {real, imag} */,
  {32'hc4aac688, 32'h00000000} /* (15, 20, 29) {real, imag} */,
  {32'hc4c73a4b, 32'h00000000} /* (15, 20, 28) {real, imag} */,
  {32'hc4fc2d52, 32'h00000000} /* (15, 20, 27) {real, imag} */,
  {32'hc4cf4614, 32'h00000000} /* (15, 20, 26) {real, imag} */,
  {32'hc4a71ea7, 32'h00000000} /* (15, 20, 25) {real, imag} */,
  {32'hc4a1165a, 32'h00000000} /* (15, 20, 24) {real, imag} */,
  {32'hc4903937, 32'h00000000} /* (15, 20, 23) {real, imag} */,
  {32'hc3c4b25e, 32'h00000000} /* (15, 20, 22) {real, imag} */,
  {32'hc2c782d8, 32'h00000000} /* (15, 20, 21) {real, imag} */,
  {32'h44323621, 32'h00000000} /* (15, 20, 20) {real, imag} */,
  {32'h44514595, 32'h00000000} /* (15, 20, 19) {real, imag} */,
  {32'h4223c930, 32'h00000000} /* (15, 20, 18) {real, imag} */,
  {32'h43f72d3d, 32'h00000000} /* (15, 20, 17) {real, imag} */,
  {32'h44a49b94, 32'h00000000} /* (15, 20, 16) {real, imag} */,
  {32'h44a95b4a, 32'h00000000} /* (15, 20, 15) {real, imag} */,
  {32'h446c50cb, 32'h00000000} /* (15, 20, 14) {real, imag} */,
  {32'h44027fd3, 32'h00000000} /* (15, 20, 13) {real, imag} */,
  {32'h4491c131, 32'h00000000} /* (15, 20, 12) {real, imag} */,
  {32'h44755d60, 32'h00000000} /* (15, 20, 11) {real, imag} */,
  {32'hc3b06732, 32'h00000000} /* (15, 20, 10) {real, imag} */,
  {32'hc3f77364, 32'h00000000} /* (15, 20, 9) {real, imag} */,
  {32'hc374e4c4, 32'h00000000} /* (15, 20, 8) {real, imag} */,
  {32'hc32722fe, 32'h00000000} /* (15, 20, 7) {real, imag} */,
  {32'hc4840088, 32'h00000000} /* (15, 20, 6) {real, imag} */,
  {32'hc4e064b4, 32'h00000000} /* (15, 20, 5) {real, imag} */,
  {32'hc3eb4966, 32'h00000000} /* (15, 20, 4) {real, imag} */,
  {32'hc4392aa3, 32'h00000000} /* (15, 20, 3) {real, imag} */,
  {32'hc44ae18b, 32'h00000000} /* (15, 20, 2) {real, imag} */,
  {32'hc486c6a3, 32'h00000000} /* (15, 20, 1) {real, imag} */,
  {32'hc442e9ac, 32'h00000000} /* (15, 20, 0) {real, imag} */,
  {32'hc41fab30, 32'h00000000} /* (15, 19, 31) {real, imag} */,
  {32'hc47e0714, 32'h00000000} /* (15, 19, 30) {real, imag} */,
  {32'hc4dbfc5c, 32'h00000000} /* (15, 19, 29) {real, imag} */,
  {32'hc4ed3306, 32'h00000000} /* (15, 19, 28) {real, imag} */,
  {32'hc53d50a1, 32'h00000000} /* (15, 19, 27) {real, imag} */,
  {32'hc4e6ff82, 32'h00000000} /* (15, 19, 26) {real, imag} */,
  {32'hc5077099, 32'h00000000} /* (15, 19, 25) {real, imag} */,
  {32'hc4958ae3, 32'h00000000} /* (15, 19, 24) {real, imag} */,
  {32'hc4485bb0, 32'h00000000} /* (15, 19, 23) {real, imag} */,
  {32'hc4487178, 32'h00000000} /* (15, 19, 22) {real, imag} */,
  {32'h428443b4, 32'h00000000} /* (15, 19, 21) {real, imag} */,
  {32'h44499fe3, 32'h00000000} /* (15, 19, 20) {real, imag} */,
  {32'h44a39f86, 32'h00000000} /* (15, 19, 19) {real, imag} */,
  {32'h441c6712, 32'h00000000} /* (15, 19, 18) {real, imag} */,
  {32'h44489d5f, 32'h00000000} /* (15, 19, 17) {real, imag} */,
  {32'h44f55a1c, 32'h00000000} /* (15, 19, 16) {real, imag} */,
  {32'h4501729e, 32'h00000000} /* (15, 19, 15) {real, imag} */,
  {32'h44dbdd02, 32'h00000000} /* (15, 19, 14) {real, imag} */,
  {32'h45043c88, 32'h00000000} /* (15, 19, 13) {real, imag} */,
  {32'h44c79650, 32'h00000000} /* (15, 19, 12) {real, imag} */,
  {32'h441d2fd4, 32'h00000000} /* (15, 19, 11) {real, imag} */,
  {32'hc3acccc8, 32'h00000000} /* (15, 19, 10) {real, imag} */,
  {32'hc3fb61da, 32'h00000000} /* (15, 19, 9) {real, imag} */,
  {32'hc36cb1d0, 32'h00000000} /* (15, 19, 8) {real, imag} */,
  {32'hc472a334, 32'h00000000} /* (15, 19, 7) {real, imag} */,
  {32'hc4b7372c, 32'h00000000} /* (15, 19, 6) {real, imag} */,
  {32'hc48238ff, 32'h00000000} /* (15, 19, 5) {real, imag} */,
  {32'hc52226f7, 32'h00000000} /* (15, 19, 4) {real, imag} */,
  {32'hc48ba698, 32'h00000000} /* (15, 19, 3) {real, imag} */,
  {32'hc42c4848, 32'h00000000} /* (15, 19, 2) {real, imag} */,
  {32'hc49bdf14, 32'h00000000} /* (15, 19, 1) {real, imag} */,
  {32'hc485637a, 32'h00000000} /* (15, 19, 0) {real, imag} */,
  {32'hc48bf031, 32'h00000000} /* (15, 18, 31) {real, imag} */,
  {32'hc4f3f3e2, 32'h00000000} /* (15, 18, 30) {real, imag} */,
  {32'hc4c6daa7, 32'h00000000} /* (15, 18, 29) {real, imag} */,
  {32'hc50f1da2, 32'h00000000} /* (15, 18, 28) {real, imag} */,
  {32'hc4d4eabc, 32'h00000000} /* (15, 18, 27) {real, imag} */,
  {32'hc4d94538, 32'h00000000} /* (15, 18, 26) {real, imag} */,
  {32'hc4c09210, 32'h00000000} /* (15, 18, 25) {real, imag} */,
  {32'hc3ba6c66, 32'h00000000} /* (15, 18, 24) {real, imag} */,
  {32'hc4d0e870, 32'h00000000} /* (15, 18, 23) {real, imag} */,
  {32'hc4b3b0de, 32'h00000000} /* (15, 18, 22) {real, imag} */,
  {32'h440f16fa, 32'h00000000} /* (15, 18, 21) {real, imag} */,
  {32'h44520b57, 32'h00000000} /* (15, 18, 20) {real, imag} */,
  {32'h44aa4e1e, 32'h00000000} /* (15, 18, 19) {real, imag} */,
  {32'h450d77b9, 32'h00000000} /* (15, 18, 18) {real, imag} */,
  {32'h44d7f283, 32'h00000000} /* (15, 18, 17) {real, imag} */,
  {32'h44ace962, 32'h00000000} /* (15, 18, 16) {real, imag} */,
  {32'h44711636, 32'h00000000} /* (15, 18, 15) {real, imag} */,
  {32'h4483f474, 32'h00000000} /* (15, 18, 14) {real, imag} */,
  {32'h44f68c11, 32'h00000000} /* (15, 18, 13) {real, imag} */,
  {32'h44d1d552, 32'h00000000} /* (15, 18, 12) {real, imag} */,
  {32'h44923a08, 32'h00000000} /* (15, 18, 11) {real, imag} */,
  {32'hc271aba0, 32'h00000000} /* (15, 18, 10) {real, imag} */,
  {32'hc4576d38, 32'h00000000} /* (15, 18, 9) {real, imag} */,
  {32'hc4b51f9a, 32'h00000000} /* (15, 18, 8) {real, imag} */,
  {32'hc523ca1c, 32'h00000000} /* (15, 18, 7) {real, imag} */,
  {32'hc516468a, 32'h00000000} /* (15, 18, 6) {real, imag} */,
  {32'hc4e4a8d9, 32'h00000000} /* (15, 18, 5) {real, imag} */,
  {32'hc44acaa7, 32'h00000000} /* (15, 18, 4) {real, imag} */,
  {32'hc4c69960, 32'h00000000} /* (15, 18, 3) {real, imag} */,
  {32'hc4bca792, 32'h00000000} /* (15, 18, 2) {real, imag} */,
  {32'hc43b8db2, 32'h00000000} /* (15, 18, 1) {real, imag} */,
  {32'hc4b0f930, 32'h00000000} /* (15, 18, 0) {real, imag} */,
  {32'hc4a235cf, 32'h00000000} /* (15, 17, 31) {real, imag} */,
  {32'hc50add90, 32'h00000000} /* (15, 17, 30) {real, imag} */,
  {32'hc4fba8fe, 32'h00000000} /* (15, 17, 29) {real, imag} */,
  {32'hc4ef84f6, 32'h00000000} /* (15, 17, 28) {real, imag} */,
  {32'hc527e296, 32'h00000000} /* (15, 17, 27) {real, imag} */,
  {32'hc50b09b2, 32'h00000000} /* (15, 17, 26) {real, imag} */,
  {32'hc5012209, 32'h00000000} /* (15, 17, 25) {real, imag} */,
  {32'hc4a934a5, 32'h00000000} /* (15, 17, 24) {real, imag} */,
  {32'hc4a3495e, 32'h00000000} /* (15, 17, 23) {real, imag} */,
  {32'hc4d6f0ba, 32'h00000000} /* (15, 17, 22) {real, imag} */,
  {32'hc3bb4788, 32'h00000000} /* (15, 17, 21) {real, imag} */,
  {32'h44758168, 32'h00000000} /* (15, 17, 20) {real, imag} */,
  {32'h44b16d8c, 32'h00000000} /* (15, 17, 19) {real, imag} */,
  {32'h44fcb8ae, 32'h00000000} /* (15, 17, 18) {real, imag} */,
  {32'h4516f0e9, 32'h00000000} /* (15, 17, 17) {real, imag} */,
  {32'h44c599f8, 32'h00000000} /* (15, 17, 16) {real, imag} */,
  {32'h44bf35db, 32'h00000000} /* (15, 17, 15) {real, imag} */,
  {32'h443917a2, 32'h00000000} /* (15, 17, 14) {real, imag} */,
  {32'h44278577, 32'h00000000} /* (15, 17, 13) {real, imag} */,
  {32'h44bff420, 32'h00000000} /* (15, 17, 12) {real, imag} */,
  {32'h4468ea92, 32'h00000000} /* (15, 17, 11) {real, imag} */,
  {32'hc4834e86, 32'h00000000} /* (15, 17, 10) {real, imag} */,
  {32'hc4a0d809, 32'h00000000} /* (15, 17, 9) {real, imag} */,
  {32'hc498b807, 32'h00000000} /* (15, 17, 8) {real, imag} */,
  {32'hc4d092fe, 32'h00000000} /* (15, 17, 7) {real, imag} */,
  {32'hc548d133, 32'h00000000} /* (15, 17, 6) {real, imag} */,
  {32'hc5284a2d, 32'h00000000} /* (15, 17, 5) {real, imag} */,
  {32'hc503cf23, 32'h00000000} /* (15, 17, 4) {real, imag} */,
  {32'hc4c61d58, 32'h00000000} /* (15, 17, 3) {real, imag} */,
  {32'hc49228b8, 32'h00000000} /* (15, 17, 2) {real, imag} */,
  {32'hc4d3ad06, 32'h00000000} /* (15, 17, 1) {real, imag} */,
  {32'hc4f93d14, 32'h00000000} /* (15, 17, 0) {real, imag} */,
  {32'hc4de2056, 32'h00000000} /* (15, 16, 31) {real, imag} */,
  {32'hc51a5c27, 32'h00000000} /* (15, 16, 30) {real, imag} */,
  {32'hc5158c55, 32'h00000000} /* (15, 16, 29) {real, imag} */,
  {32'hc4d63a8f, 32'h00000000} /* (15, 16, 28) {real, imag} */,
  {32'hc548ba92, 32'h00000000} /* (15, 16, 27) {real, imag} */,
  {32'hc5462fd6, 32'h00000000} /* (15, 16, 26) {real, imag} */,
  {32'hc540178d, 32'h00000000} /* (15, 16, 25) {real, imag} */,
  {32'hc526eac6, 32'h00000000} /* (15, 16, 24) {real, imag} */,
  {32'hc4bd86a2, 32'h00000000} /* (15, 16, 23) {real, imag} */,
  {32'hc4f9def0, 32'h00000000} /* (15, 16, 22) {real, imag} */,
  {32'hc3e8b280, 32'h00000000} /* (15, 16, 21) {real, imag} */,
  {32'h4476ff5a, 32'h00000000} /* (15, 16, 20) {real, imag} */,
  {32'h44f31586, 32'h00000000} /* (15, 16, 19) {real, imag} */,
  {32'h451fd005, 32'h00000000} /* (15, 16, 18) {real, imag} */,
  {32'h44ff3842, 32'h00000000} /* (15, 16, 17) {real, imag} */,
  {32'h449a2826, 32'h00000000} /* (15, 16, 16) {real, imag} */,
  {32'h4492ece0, 32'h00000000} /* (15, 16, 15) {real, imag} */,
  {32'h449e2822, 32'h00000000} /* (15, 16, 14) {real, imag} */,
  {32'h44b5db7e, 32'h00000000} /* (15, 16, 13) {real, imag} */,
  {32'h449c77e7, 32'h00000000} /* (15, 16, 12) {real, imag} */,
  {32'h44604aa8, 32'h00000000} /* (15, 16, 11) {real, imag} */,
  {32'h43c25ea4, 32'h00000000} /* (15, 16, 10) {real, imag} */,
  {32'hc40ba5d4, 32'h00000000} /* (15, 16, 9) {real, imag} */,
  {32'hc4c05adb, 32'h00000000} /* (15, 16, 8) {real, imag} */,
  {32'hc51dc520, 32'h00000000} /* (15, 16, 7) {real, imag} */,
  {32'hc5356556, 32'h00000000} /* (15, 16, 6) {real, imag} */,
  {32'hc525c18a, 32'h00000000} /* (15, 16, 5) {real, imag} */,
  {32'hc4e6dfc7, 32'h00000000} /* (15, 16, 4) {real, imag} */,
  {32'hc4b51c1e, 32'h00000000} /* (15, 16, 3) {real, imag} */,
  {32'hc4d41c26, 32'h00000000} /* (15, 16, 2) {real, imag} */,
  {32'hc4f29340, 32'h00000000} /* (15, 16, 1) {real, imag} */,
  {32'hc4aabb44, 32'h00000000} /* (15, 16, 0) {real, imag} */,
  {32'hc5058161, 32'h00000000} /* (15, 15, 31) {real, imag} */,
  {32'hc51e1594, 32'h00000000} /* (15, 15, 30) {real, imag} */,
  {32'hc4fc05f6, 32'h00000000} /* (15, 15, 29) {real, imag} */,
  {32'hc5079621, 32'h00000000} /* (15, 15, 28) {real, imag} */,
  {32'hc52b267a, 32'h00000000} /* (15, 15, 27) {real, imag} */,
  {32'hc5636870, 32'h00000000} /* (15, 15, 26) {real, imag} */,
  {32'hc55d113a, 32'h00000000} /* (15, 15, 25) {real, imag} */,
  {32'hc51ae1ca, 32'h00000000} /* (15, 15, 24) {real, imag} */,
  {32'hc4c11d47, 32'h00000000} /* (15, 15, 23) {real, imag} */,
  {32'hc4b7b9fd, 32'h00000000} /* (15, 15, 22) {real, imag} */,
  {32'h43cbce1c, 32'h00000000} /* (15, 15, 21) {real, imag} */,
  {32'h43e8dc66, 32'h00000000} /* (15, 15, 20) {real, imag} */,
  {32'h44cb1e1b, 32'h00000000} /* (15, 15, 19) {real, imag} */,
  {32'h454d32d3, 32'h00000000} /* (15, 15, 18) {real, imag} */,
  {32'h45020558, 32'h00000000} /* (15, 15, 17) {real, imag} */,
  {32'h452b828a, 32'h00000000} /* (15, 15, 16) {real, imag} */,
  {32'h44c23c16, 32'h00000000} /* (15, 15, 15) {real, imag} */,
  {32'h44e41ae8, 32'h00000000} /* (15, 15, 14) {real, imag} */,
  {32'h45079c5f, 32'h00000000} /* (15, 15, 13) {real, imag} */,
  {32'h44c73bac, 32'h00000000} /* (15, 15, 12) {real, imag} */,
  {32'h44b8ced1, 32'h00000000} /* (15, 15, 11) {real, imag} */,
  {32'h431bd678, 32'h00000000} /* (15, 15, 10) {real, imag} */,
  {32'hc463973e, 32'h00000000} /* (15, 15, 9) {real, imag} */,
  {32'hc4807ce4, 32'h00000000} /* (15, 15, 8) {real, imag} */,
  {32'hc4e29e03, 32'h00000000} /* (15, 15, 7) {real, imag} */,
  {32'hc512f6ed, 32'h00000000} /* (15, 15, 6) {real, imag} */,
  {32'hc528ac62, 32'h00000000} /* (15, 15, 5) {real, imag} */,
  {32'hc4e1a4a8, 32'h00000000} /* (15, 15, 4) {real, imag} */,
  {32'hc4c1a553, 32'h00000000} /* (15, 15, 3) {real, imag} */,
  {32'hc4eeb2e6, 32'h00000000} /* (15, 15, 2) {real, imag} */,
  {32'hc4ed5be8, 32'h00000000} /* (15, 15, 1) {real, imag} */,
  {32'hc4e3979c, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hc501fa40, 32'h00000000} /* (15, 14, 31) {real, imag} */,
  {32'hc504d9d6, 32'h00000000} /* (15, 14, 30) {real, imag} */,
  {32'hc57e4104, 32'h00000000} /* (15, 14, 29) {real, imag} */,
  {32'hc5819b1a, 32'h00000000} /* (15, 14, 28) {real, imag} */,
  {32'hc5394545, 32'h00000000} /* (15, 14, 27) {real, imag} */,
  {32'hc53d2b69, 32'h00000000} /* (15, 14, 26) {real, imag} */,
  {32'hc577af09, 32'h00000000} /* (15, 14, 25) {real, imag} */,
  {32'hc50be0f3, 32'h00000000} /* (15, 14, 24) {real, imag} */,
  {32'hc4d1b8d8, 32'h00000000} /* (15, 14, 23) {real, imag} */,
  {32'hc48c5912, 32'h00000000} /* (15, 14, 22) {real, imag} */,
  {32'hc43ed14c, 32'h00000000} /* (15, 14, 21) {real, imag} */,
  {32'h4497d7ce, 32'h00000000} /* (15, 14, 20) {real, imag} */,
  {32'h44df9181, 32'h00000000} /* (15, 14, 19) {real, imag} */,
  {32'h4532567f, 32'h00000000} /* (15, 14, 18) {real, imag} */,
  {32'h453d86af, 32'h00000000} /* (15, 14, 17) {real, imag} */,
  {32'h4504993f, 32'h00000000} /* (15, 14, 16) {real, imag} */,
  {32'h452184a4, 32'h00000000} /* (15, 14, 15) {real, imag} */,
  {32'h44dd9e80, 32'h00000000} /* (15, 14, 14) {real, imag} */,
  {32'h450598a4, 32'h00000000} /* (15, 14, 13) {real, imag} */,
  {32'h44dd3afe, 32'h00000000} /* (15, 14, 12) {real, imag} */,
  {32'h450b2b27, 32'h00000000} /* (15, 14, 11) {real, imag} */,
  {32'h447b0ddb, 32'h00000000} /* (15, 14, 10) {real, imag} */,
  {32'hc3dfb9f8, 32'h00000000} /* (15, 14, 9) {real, imag} */,
  {32'hc43bbb34, 32'h00000000} /* (15, 14, 8) {real, imag} */,
  {32'hc4d44308, 32'h00000000} /* (15, 14, 7) {real, imag} */,
  {32'hc511f815, 32'h00000000} /* (15, 14, 6) {real, imag} */,
  {32'hc4e5eeda, 32'h00000000} /* (15, 14, 5) {real, imag} */,
  {32'hc4bfbdb2, 32'h00000000} /* (15, 14, 4) {real, imag} */,
  {32'hc4a16713, 32'h00000000} /* (15, 14, 3) {real, imag} */,
  {32'hc4f194f2, 32'h00000000} /* (15, 14, 2) {real, imag} */,
  {32'hc50f9e0b, 32'h00000000} /* (15, 14, 1) {real, imag} */,
  {32'hc4df4160, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'hc49eddf9, 32'h00000000} /* (15, 13, 31) {real, imag} */,
  {32'hc5068f06, 32'h00000000} /* (15, 13, 30) {real, imag} */,
  {32'hc52746a3, 32'h00000000} /* (15, 13, 29) {real, imag} */,
  {32'hc50a6e7b, 32'h00000000} /* (15, 13, 28) {real, imag} */,
  {32'hc5034f01, 32'h00000000} /* (15, 13, 27) {real, imag} */,
  {32'hc508a367, 32'h00000000} /* (15, 13, 26) {real, imag} */,
  {32'hc503dcfc, 32'h00000000} /* (15, 13, 25) {real, imag} */,
  {32'hc513178d, 32'h00000000} /* (15, 13, 24) {real, imag} */,
  {32'hc5075f45, 32'h00000000} /* (15, 13, 23) {real, imag} */,
  {32'hc4b522fa, 32'h00000000} /* (15, 13, 22) {real, imag} */,
  {32'hc4596ebc, 32'h00000000} /* (15, 13, 21) {real, imag} */,
  {32'h4363dba8, 32'h00000000} /* (15, 13, 20) {real, imag} */,
  {32'h44dc6cb9, 32'h00000000} /* (15, 13, 19) {real, imag} */,
  {32'h45179a3a, 32'h00000000} /* (15, 13, 18) {real, imag} */,
  {32'h44cafe39, 32'h00000000} /* (15, 13, 17) {real, imag} */,
  {32'h44f3b63e, 32'h00000000} /* (15, 13, 16) {real, imag} */,
  {32'h44ea917b, 32'h00000000} /* (15, 13, 15) {real, imag} */,
  {32'h4519dfd0, 32'h00000000} /* (15, 13, 14) {real, imag} */,
  {32'h44e22382, 32'h00000000} /* (15, 13, 13) {real, imag} */,
  {32'h44f007aa, 32'h00000000} /* (15, 13, 12) {real, imag} */,
  {32'h44b24fbf, 32'h00000000} /* (15, 13, 11) {real, imag} */,
  {32'h43eac7c6, 32'h00000000} /* (15, 13, 10) {real, imag} */,
  {32'h43a8b44c, 32'h00000000} /* (15, 13, 9) {real, imag} */,
  {32'hc3225eb0, 32'h00000000} /* (15, 13, 8) {real, imag} */,
  {32'hc4e1b0dc, 32'h00000000} /* (15, 13, 7) {real, imag} */,
  {32'hc5159b6f, 32'h00000000} /* (15, 13, 6) {real, imag} */,
  {32'hc46f506a, 32'h00000000} /* (15, 13, 5) {real, imag} */,
  {32'hc4b2b79b, 32'h00000000} /* (15, 13, 4) {real, imag} */,
  {32'hc4999633, 32'h00000000} /* (15, 13, 3) {real, imag} */,
  {32'hc497145a, 32'h00000000} /* (15, 13, 2) {real, imag} */,
  {32'hc48a5f0f, 32'h00000000} /* (15, 13, 1) {real, imag} */,
  {32'hc50327bf, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'hc49d1693, 32'h00000000} /* (15, 12, 31) {real, imag} */,
  {32'hc4dd848e, 32'h00000000} /* (15, 12, 30) {real, imag} */,
  {32'hc4da14fd, 32'h00000000} /* (15, 12, 29) {real, imag} */,
  {32'hc44a6d1e, 32'h00000000} /* (15, 12, 28) {real, imag} */,
  {32'hc4bdadff, 32'h00000000} /* (15, 12, 27) {real, imag} */,
  {32'hc4987f7e, 32'h00000000} /* (15, 12, 26) {real, imag} */,
  {32'hc4d729ca, 32'h00000000} /* (15, 12, 25) {real, imag} */,
  {32'hc4c4ce20, 32'h00000000} /* (15, 12, 24) {real, imag} */,
  {32'hc44ace51, 32'h00000000} /* (15, 12, 23) {real, imag} */,
  {32'hc45211aa, 32'h00000000} /* (15, 12, 22) {real, imag} */,
  {32'h43ce3380, 32'h00000000} /* (15, 12, 21) {real, imag} */,
  {32'h44ab1f6c, 32'h00000000} /* (15, 12, 20) {real, imag} */,
  {32'h44d560d0, 32'h00000000} /* (15, 12, 19) {real, imag} */,
  {32'h44dbf4e2, 32'h00000000} /* (15, 12, 18) {real, imag} */,
  {32'h45264ed5, 32'h00000000} /* (15, 12, 17) {real, imag} */,
  {32'h452d3a12, 32'h00000000} /* (15, 12, 16) {real, imag} */,
  {32'h44760c7e, 32'h00000000} /* (15, 12, 15) {real, imag} */,
  {32'h44922540, 32'h00000000} /* (15, 12, 14) {real, imag} */,
  {32'h44f0a083, 32'h00000000} /* (15, 12, 13) {real, imag} */,
  {32'h45467734, 32'h00000000} /* (15, 12, 12) {real, imag} */,
  {32'h450e1d34, 32'h00000000} /* (15, 12, 11) {real, imag} */,
  {32'h437effd4, 32'h00000000} /* (15, 12, 10) {real, imag} */,
  {32'h4139e400, 32'h00000000} /* (15, 12, 9) {real, imag} */,
  {32'hc4b5b918, 32'h00000000} /* (15, 12, 8) {real, imag} */,
  {32'hc3ee5eda, 32'h00000000} /* (15, 12, 7) {real, imag} */,
  {32'hc3dc8dfc, 32'h00000000} /* (15, 12, 6) {real, imag} */,
  {32'hc41f33ec, 32'h00000000} /* (15, 12, 5) {real, imag} */,
  {32'hc424f226, 32'h00000000} /* (15, 12, 4) {real, imag} */,
  {32'hc47c95c9, 32'h00000000} /* (15, 12, 3) {real, imag} */,
  {32'hc3df24a2, 32'h00000000} /* (15, 12, 2) {real, imag} */,
  {32'hc419dd64, 32'h00000000} /* (15, 12, 1) {real, imag} */,
  {32'hc47acbc1, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'h436f0b70, 32'h00000000} /* (15, 11, 31) {real, imag} */,
  {32'hc3289ed0, 32'h00000000} /* (15, 11, 30) {real, imag} */,
  {32'hc48257e4, 32'h00000000} /* (15, 11, 29) {real, imag} */,
  {32'hc478c9fa, 32'h00000000} /* (15, 11, 28) {real, imag} */,
  {32'hc4237007, 32'h00000000} /* (15, 11, 27) {real, imag} */,
  {32'hc41f5eb0, 32'h00000000} /* (15, 11, 26) {real, imag} */,
  {32'hc4415917, 32'h00000000} /* (15, 11, 25) {real, imag} */,
  {32'h429fe634, 32'h00000000} /* (15, 11, 24) {real, imag} */,
  {32'hc5041904, 32'h00000000} /* (15, 11, 23) {real, imag} */,
  {32'hc34fa09e, 32'h00000000} /* (15, 11, 22) {real, imag} */,
  {32'h44a123b8, 32'h00000000} /* (15, 11, 21) {real, imag} */,
  {32'h44d432fa, 32'h00000000} /* (15, 11, 20) {real, imag} */,
  {32'h44f4ee67, 32'h00000000} /* (15, 11, 19) {real, imag} */,
  {32'h450ced28, 32'h00000000} /* (15, 11, 18) {real, imag} */,
  {32'h44f805ba, 32'h00000000} /* (15, 11, 17) {real, imag} */,
  {32'h450733c1, 32'h00000000} /* (15, 11, 16) {real, imag} */,
  {32'h44cb9f58, 32'h00000000} /* (15, 11, 15) {real, imag} */,
  {32'h44d2802c, 32'h00000000} /* (15, 11, 14) {real, imag} */,
  {32'h44bcfa8c, 32'h00000000} /* (15, 11, 13) {real, imag} */,
  {32'h449e6f95, 32'h00000000} /* (15, 11, 12) {real, imag} */,
  {32'h451cc1ef, 32'h00000000} /* (15, 11, 11) {real, imag} */,
  {32'h438aa6df, 32'h00000000} /* (15, 11, 10) {real, imag} */,
  {32'hc283a018, 32'h00000000} /* (15, 11, 9) {real, imag} */,
  {32'hc439da2e, 32'h00000000} /* (15, 11, 8) {real, imag} */,
  {32'hc396c43c, 32'h00000000} /* (15, 11, 7) {real, imag} */,
  {32'h4395665d, 32'h00000000} /* (15, 11, 6) {real, imag} */,
  {32'hc38237c6, 32'h00000000} /* (15, 11, 5) {real, imag} */,
  {32'h41af18e0, 32'h00000000} /* (15, 11, 4) {real, imag} */,
  {32'h43b69a04, 32'h00000000} /* (15, 11, 3) {real, imag} */,
  {32'h436ccbdc, 32'h00000000} /* (15, 11, 2) {real, imag} */,
  {32'hc358fdb4, 32'h00000000} /* (15, 11, 1) {real, imag} */,
  {32'hc3947278, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h43f2647e, 32'h00000000} /* (15, 10, 31) {real, imag} */,
  {32'h44ae305d, 32'h00000000} /* (15, 10, 30) {real, imag} */,
  {32'h44b4211b, 32'h00000000} /* (15, 10, 29) {real, imag} */,
  {32'h4427f95e, 32'h00000000} /* (15, 10, 28) {real, imag} */,
  {32'h43e40687, 32'h00000000} /* (15, 10, 27) {real, imag} */,
  {32'h441af90a, 32'h00000000} /* (15, 10, 26) {real, imag} */,
  {32'h439e1e99, 32'h00000000} /* (15, 10, 25) {real, imag} */,
  {32'hc2c4e350, 32'h00000000} /* (15, 10, 24) {real, imag} */,
  {32'hc48cc90f, 32'h00000000} /* (15, 10, 23) {real, imag} */,
  {32'h44efb254, 32'h00000000} /* (15, 10, 22) {real, imag} */,
  {32'h4469ae43, 32'h00000000} /* (15, 10, 21) {real, imag} */,
  {32'h44486043, 32'h00000000} /* (15, 10, 20) {real, imag} */,
  {32'hc1a8f740, 32'h00000000} /* (15, 10, 19) {real, imag} */,
  {32'h44989240, 32'h00000000} /* (15, 10, 18) {real, imag} */,
  {32'h44a91848, 32'h00000000} /* (15, 10, 17) {real, imag} */,
  {32'h440b4737, 32'h00000000} /* (15, 10, 16) {real, imag} */,
  {32'h42c724c6, 32'h00000000} /* (15, 10, 15) {real, imag} */,
  {32'h447059b6, 32'h00000000} /* (15, 10, 14) {real, imag} */,
  {32'h43d66479, 32'h00000000} /* (15, 10, 13) {real, imag} */,
  {32'h4302da26, 32'h00000000} /* (15, 10, 12) {real, imag} */,
  {32'h43babcd9, 32'h00000000} /* (15, 10, 11) {real, imag} */,
  {32'h43a107e4, 32'h00000000} /* (15, 10, 10) {real, imag} */,
  {32'h44502bd6, 32'h00000000} /* (15, 10, 9) {real, imag} */,
  {32'h445aa204, 32'h00000000} /* (15, 10, 8) {real, imag} */,
  {32'h449a1203, 32'h00000000} /* (15, 10, 7) {real, imag} */,
  {32'h443a6128, 32'h00000000} /* (15, 10, 6) {real, imag} */,
  {32'h4508088d, 32'h00000000} /* (15, 10, 5) {real, imag} */,
  {32'h4425a4c5, 32'h00000000} /* (15, 10, 4) {real, imag} */,
  {32'h44b3c109, 32'h00000000} /* (15, 10, 3) {real, imag} */,
  {32'h44fbbb9a, 32'h00000000} /* (15, 10, 2) {real, imag} */,
  {32'h44806734, 32'h00000000} /* (15, 10, 1) {real, imag} */,
  {32'h44861318, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'h4495758c, 32'h00000000} /* (15, 9, 31) {real, imag} */,
  {32'h44631de8, 32'h00000000} /* (15, 9, 30) {real, imag} */,
  {32'h44a8c5d6, 32'h00000000} /* (15, 9, 29) {real, imag} */,
  {32'h4514d472, 32'h00000000} /* (15, 9, 28) {real, imag} */,
  {32'h449d7fd0, 32'h00000000} /* (15, 9, 27) {real, imag} */,
  {32'h44c3c5ee, 32'h00000000} /* (15, 9, 26) {real, imag} */,
  {32'h446c9921, 32'h00000000} /* (15, 9, 25) {real, imag} */,
  {32'h444d4de9, 32'h00000000} /* (15, 9, 24) {real, imag} */,
  {32'h44be89c2, 32'h00000000} /* (15, 9, 23) {real, imag} */,
  {32'h45048e26, 32'h00000000} /* (15, 9, 22) {real, imag} */,
  {32'h4428addb, 32'h00000000} /* (15, 9, 21) {real, imag} */,
  {32'h41b2ae00, 32'h00000000} /* (15, 9, 20) {real, imag} */,
  {32'h435e4ab8, 32'h00000000} /* (15, 9, 19) {real, imag} */,
  {32'h43c074a0, 32'h00000000} /* (15, 9, 18) {real, imag} */,
  {32'h43c387b8, 32'h00000000} /* (15, 9, 17) {real, imag} */,
  {32'h44a79742, 32'h00000000} /* (15, 9, 16) {real, imag} */,
  {32'hc48bd7e4, 32'h00000000} /* (15, 9, 15) {real, imag} */,
  {32'hc27fbe20, 32'h00000000} /* (15, 9, 14) {real, imag} */,
  {32'hc2cc2180, 32'h00000000} /* (15, 9, 13) {real, imag} */,
  {32'h43b4c04e, 32'h00000000} /* (15, 9, 12) {real, imag} */,
  {32'hc215fd10, 32'h00000000} /* (15, 9, 11) {real, imag} */,
  {32'hc275e350, 32'h00000000} /* (15, 9, 10) {real, imag} */,
  {32'h4482415a, 32'h00000000} /* (15, 9, 9) {real, imag} */,
  {32'h4430f87f, 32'h00000000} /* (15, 9, 8) {real, imag} */,
  {32'h4451e7db, 32'h00000000} /* (15, 9, 7) {real, imag} */,
  {32'h45114a56, 32'h00000000} /* (15, 9, 6) {real, imag} */,
  {32'h4504ab9c, 32'h00000000} /* (15, 9, 5) {real, imag} */,
  {32'h45066540, 32'h00000000} /* (15, 9, 4) {real, imag} */,
  {32'h45108b32, 32'h00000000} /* (15, 9, 3) {real, imag} */,
  {32'h44dc1120, 32'h00000000} /* (15, 9, 2) {real, imag} */,
  {32'h44d25648, 32'h00000000} /* (15, 9, 1) {real, imag} */,
  {32'h4483d542, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'h4381c05d, 32'h00000000} /* (15, 8, 31) {real, imag} */,
  {32'h44ee5109, 32'h00000000} /* (15, 8, 30) {real, imag} */,
  {32'h44e5cc25, 32'h00000000} /* (15, 8, 29) {real, imag} */,
  {32'h44b0b6c9, 32'h00000000} /* (15, 8, 28) {real, imag} */,
  {32'h450b82a0, 32'h00000000} /* (15, 8, 27) {real, imag} */,
  {32'h450ff0c8, 32'h00000000} /* (15, 8, 26) {real, imag} */,
  {32'h44a7d27a, 32'h00000000} /* (15, 8, 25) {real, imag} */,
  {32'h44d3e225, 32'h00000000} /* (15, 8, 24) {real, imag} */,
  {32'h44c9c850, 32'h00000000} /* (15, 8, 23) {real, imag} */,
  {32'h44d9fa90, 32'h00000000} /* (15, 8, 22) {real, imag} */,
  {32'h4520145e, 32'h00000000} /* (15, 8, 21) {real, imag} */,
  {32'h4393c50c, 32'h00000000} /* (15, 8, 20) {real, imag} */,
  {32'h435908b8, 32'h00000000} /* (15, 8, 19) {real, imag} */,
  {32'hc3eaf2d9, 32'h00000000} /* (15, 8, 18) {real, imag} */,
  {32'h437c6c94, 32'h00000000} /* (15, 8, 17) {real, imag} */,
  {32'h43edb83c, 32'h00000000} /* (15, 8, 16) {real, imag} */,
  {32'hc3ffc94d, 32'h00000000} /* (15, 8, 15) {real, imag} */,
  {32'hc3a88234, 32'h00000000} /* (15, 8, 14) {real, imag} */,
  {32'hc3b26f24, 32'h00000000} /* (15, 8, 13) {real, imag} */,
  {32'hc492e009, 32'h00000000} /* (15, 8, 12) {real, imag} */,
  {32'hc439b5b9, 32'h00000000} /* (15, 8, 11) {real, imag} */,
  {32'h43eaffa4, 32'h00000000} /* (15, 8, 10) {real, imag} */,
  {32'h448b66fc, 32'h00000000} /* (15, 8, 9) {real, imag} */,
  {32'h448a624f, 32'h00000000} /* (15, 8, 8) {real, imag} */,
  {32'h447f7538, 32'h00000000} /* (15, 8, 7) {real, imag} */,
  {32'h455671be, 32'h00000000} /* (15, 8, 6) {real, imag} */,
  {32'h44cf651f, 32'h00000000} /* (15, 8, 5) {real, imag} */,
  {32'h45067006, 32'h00000000} /* (15, 8, 4) {real, imag} */,
  {32'h450229fe, 32'h00000000} /* (15, 8, 3) {real, imag} */,
  {32'h44a49c17, 32'h00000000} /* (15, 8, 2) {real, imag} */,
  {32'h4486ebfe, 32'h00000000} /* (15, 8, 1) {real, imag} */,
  {32'h449c1391, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h44d004ae, 32'h00000000} /* (15, 7, 31) {real, imag} */,
  {32'h44fe4fb0, 32'h00000000} /* (15, 7, 30) {real, imag} */,
  {32'h4518225e, 32'h00000000} /* (15, 7, 29) {real, imag} */,
  {32'h44e52ca8, 32'h00000000} /* (15, 7, 28) {real, imag} */,
  {32'h44d01310, 32'h00000000} /* (15, 7, 27) {real, imag} */,
  {32'h44e1fe1a, 32'h00000000} /* (15, 7, 26) {real, imag} */,
  {32'h44f399de, 32'h00000000} /* (15, 7, 25) {real, imag} */,
  {32'h44d2c3da, 32'h00000000} /* (15, 7, 24) {real, imag} */,
  {32'h44fbe5c1, 32'h00000000} /* (15, 7, 23) {real, imag} */,
  {32'h4516ef12, 32'h00000000} /* (15, 7, 22) {real, imag} */,
  {32'h44c8e505, 32'h00000000} /* (15, 7, 21) {real, imag} */,
  {32'h4368cfa8, 32'h00000000} /* (15, 7, 20) {real, imag} */,
  {32'hc38509c2, 32'h00000000} /* (15, 7, 19) {real, imag} */,
  {32'hc3b1b986, 32'h00000000} /* (15, 7, 18) {real, imag} */,
  {32'h43e0d12a, 32'h00000000} /* (15, 7, 17) {real, imag} */,
  {32'hc3d9e7b4, 32'h00000000} /* (15, 7, 16) {real, imag} */,
  {32'hc3d8b4a2, 32'h00000000} /* (15, 7, 15) {real, imag} */,
  {32'hc40d4450, 32'h00000000} /* (15, 7, 14) {real, imag} */,
  {32'hc4572591, 32'h00000000} /* (15, 7, 13) {real, imag} */,
  {32'hc4786208, 32'h00000000} /* (15, 7, 12) {real, imag} */,
  {32'hc211e7f0, 32'h00000000} /* (15, 7, 11) {real, imag} */,
  {32'h44926dfa, 32'h00000000} /* (15, 7, 10) {real, imag} */,
  {32'h4405ee8f, 32'h00000000} /* (15, 7, 9) {real, imag} */,
  {32'h45002142, 32'h00000000} /* (15, 7, 8) {real, imag} */,
  {32'h4505d0b5, 32'h00000000} /* (15, 7, 7) {real, imag} */,
  {32'h44e1238b, 32'h00000000} /* (15, 7, 6) {real, imag} */,
  {32'h452c37a2, 32'h00000000} /* (15, 7, 5) {real, imag} */,
  {32'h450c4902, 32'h00000000} /* (15, 7, 4) {real, imag} */,
  {32'h44fff660, 32'h00000000} /* (15, 7, 3) {real, imag} */,
  {32'h4497bf14, 32'h00000000} /* (15, 7, 2) {real, imag} */,
  {32'h44ce3814, 32'h00000000} /* (15, 7, 1) {real, imag} */,
  {32'h44ac8e03, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'h44b36be9, 32'h00000000} /* (15, 6, 31) {real, imag} */,
  {32'h44e0c2f8, 32'h00000000} /* (15, 6, 30) {real, imag} */,
  {32'h4487ab99, 32'h00000000} /* (15, 6, 29) {real, imag} */,
  {32'h44ce1af0, 32'h00000000} /* (15, 6, 28) {real, imag} */,
  {32'h44c907da, 32'h00000000} /* (15, 6, 27) {real, imag} */,
  {32'h45256e9e, 32'h00000000} /* (15, 6, 26) {real, imag} */,
  {32'h44f3ade6, 32'h00000000} /* (15, 6, 25) {real, imag} */,
  {32'h4519fa55, 32'h00000000} /* (15, 6, 24) {real, imag} */,
  {32'h451ff2ba, 32'h00000000} /* (15, 6, 23) {real, imag} */,
  {32'h450de46b, 32'h00000000} /* (15, 6, 22) {real, imag} */,
  {32'h4508e4a1, 32'h00000000} /* (15, 6, 21) {real, imag} */,
  {32'h44052ef2, 32'h00000000} /* (15, 6, 20) {real, imag} */,
  {32'h4117ef00, 32'h00000000} /* (15, 6, 19) {real, imag} */,
  {32'hc395d38c, 32'h00000000} /* (15, 6, 18) {real, imag} */,
  {32'hc42b2664, 32'h00000000} /* (15, 6, 17) {real, imag} */,
  {32'hc3f08f3a, 32'h00000000} /* (15, 6, 16) {real, imag} */,
  {32'hc36a0308, 32'h00000000} /* (15, 6, 15) {real, imag} */,
  {32'hc40bb823, 32'h00000000} /* (15, 6, 14) {real, imag} */,
  {32'hc3cecf7c, 32'h00000000} /* (15, 6, 13) {real, imag} */,
  {32'hc433d2d7, 32'h00000000} /* (15, 6, 12) {real, imag} */,
  {32'hc312b878, 32'h00000000} /* (15, 6, 11) {real, imag} */,
  {32'h441fcadd, 32'h00000000} /* (15, 6, 10) {real, imag} */,
  {32'h44067ff8, 32'h00000000} /* (15, 6, 9) {real, imag} */,
  {32'h44b34842, 32'h00000000} /* (15, 6, 8) {real, imag} */,
  {32'h448f9048, 32'h00000000} /* (15, 6, 7) {real, imag} */,
  {32'h44c6bb2a, 32'h00000000} /* (15, 6, 6) {real, imag} */,
  {32'h451cc6b7, 32'h00000000} /* (15, 6, 5) {real, imag} */,
  {32'h4513021e, 32'h00000000} /* (15, 6, 4) {real, imag} */,
  {32'h44e54e63, 32'h00000000} /* (15, 6, 3) {real, imag} */,
  {32'h44d4a981, 32'h00000000} /* (15, 6, 2) {real, imag} */,
  {32'h44cce4a8, 32'h00000000} /* (15, 6, 1) {real, imag} */,
  {32'h44a8c388, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h44bf4c00, 32'h00000000} /* (15, 5, 31) {real, imag} */,
  {32'h4521c590, 32'h00000000} /* (15, 5, 30) {real, imag} */,
  {32'h44d3097d, 32'h00000000} /* (15, 5, 29) {real, imag} */,
  {32'h45399ea0, 32'h00000000} /* (15, 5, 28) {real, imag} */,
  {32'h4530fa13, 32'h00000000} /* (15, 5, 27) {real, imag} */,
  {32'h45192597, 32'h00000000} /* (15, 5, 26) {real, imag} */,
  {32'h45081360, 32'h00000000} /* (15, 5, 25) {real, imag} */,
  {32'h45519de0, 32'h00000000} /* (15, 5, 24) {real, imag} */,
  {32'h4526756a, 32'h00000000} /* (15, 5, 23) {real, imag} */,
  {32'h4504f9fe, 32'h00000000} /* (15, 5, 22) {real, imag} */,
  {32'h44c6bc38, 32'h00000000} /* (15, 5, 21) {real, imag} */,
  {32'h44da34ca, 32'h00000000} /* (15, 5, 20) {real, imag} */,
  {32'h43a9f6fe, 32'h00000000} /* (15, 5, 19) {real, imag} */,
  {32'h43383720, 32'h00000000} /* (15, 5, 18) {real, imag} */,
  {32'hc40cc782, 32'h00000000} /* (15, 5, 17) {real, imag} */,
  {32'hc22391a0, 32'h00000000} /* (15, 5, 16) {real, imag} */,
  {32'hc3eeadd0, 32'h00000000} /* (15, 5, 15) {real, imag} */,
  {32'hc4833c9c, 32'h00000000} /* (15, 5, 14) {real, imag} */,
  {32'hc371f8b8, 32'h00000000} /* (15, 5, 13) {real, imag} */,
  {32'hc4d5ac4d, 32'h00000000} /* (15, 5, 12) {real, imag} */,
  {32'hc4adb556, 32'h00000000} /* (15, 5, 11) {real, imag} */,
  {32'hc4cebf86, 32'h00000000} /* (15, 5, 10) {real, imag} */,
  {32'h435f8374, 32'h00000000} /* (15, 5, 9) {real, imag} */,
  {32'h42ea5950, 32'h00000000} /* (15, 5, 8) {real, imag} */,
  {32'hc39ff048, 32'h00000000} /* (15, 5, 7) {real, imag} */,
  {32'h44c4e45f, 32'h00000000} /* (15, 5, 6) {real, imag} */,
  {32'h44df592a, 32'h00000000} /* (15, 5, 5) {real, imag} */,
  {32'h4555f1b7, 32'h00000000} /* (15, 5, 4) {real, imag} */,
  {32'h44d7b31e, 32'h00000000} /* (15, 5, 3) {real, imag} */,
  {32'h44c58ccd, 32'h00000000} /* (15, 5, 2) {real, imag} */,
  {32'h44d99a8d, 32'h00000000} /* (15, 5, 1) {real, imag} */,
  {32'h44a52f6b, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'h44cd0bae, 32'h00000000} /* (15, 4, 31) {real, imag} */,
  {32'h4509421e, 32'h00000000} /* (15, 4, 30) {real, imag} */,
  {32'h451e84d9, 32'h00000000} /* (15, 4, 29) {real, imag} */,
  {32'h45332bca, 32'h00000000} /* (15, 4, 28) {real, imag} */,
  {32'h453f433e, 32'h00000000} /* (15, 4, 27) {real, imag} */,
  {32'h4529da74, 32'h00000000} /* (15, 4, 26) {real, imag} */,
  {32'h4520ff6f, 32'h00000000} /* (15, 4, 25) {real, imag} */,
  {32'h455cf6bc, 32'h00000000} /* (15, 4, 24) {real, imag} */,
  {32'h452b08e6, 32'h00000000} /* (15, 4, 23) {real, imag} */,
  {32'h452f9160, 32'h00000000} /* (15, 4, 22) {real, imag} */,
  {32'h452398bb, 32'h00000000} /* (15, 4, 21) {real, imag} */,
  {32'h45010249, 32'h00000000} /* (15, 4, 20) {real, imag} */,
  {32'h4482cd14, 32'h00000000} /* (15, 4, 19) {real, imag} */,
  {32'h44429766, 32'h00000000} /* (15, 4, 18) {real, imag} */,
  {32'h4446c110, 32'h00000000} /* (15, 4, 17) {real, imag} */,
  {32'h43840258, 32'h00000000} /* (15, 4, 16) {real, imag} */,
  {32'hc45b34d4, 32'h00000000} /* (15, 4, 15) {real, imag} */,
  {32'hc41446d8, 32'h00000000} /* (15, 4, 14) {real, imag} */,
  {32'hc4a70ad6, 32'h00000000} /* (15, 4, 13) {real, imag} */,
  {32'hc40f79a0, 32'h00000000} /* (15, 4, 12) {real, imag} */,
  {32'hc502cf42, 32'h00000000} /* (15, 4, 11) {real, imag} */,
  {32'hc4128210, 32'h00000000} /* (15, 4, 10) {real, imag} */,
  {32'hc42e50cd, 32'h00000000} /* (15, 4, 9) {real, imag} */,
  {32'hc4a33f39, 32'h00000000} /* (15, 4, 8) {real, imag} */,
  {32'hc3cdd538, 32'h00000000} /* (15, 4, 7) {real, imag} */,
  {32'h438e930c, 32'h00000000} /* (15, 4, 6) {real, imag} */,
  {32'h449837c2, 32'h00000000} /* (15, 4, 5) {real, imag} */,
  {32'h4505714d, 32'h00000000} /* (15, 4, 4) {real, imag} */,
  {32'h45274c23, 32'h00000000} /* (15, 4, 3) {real, imag} */,
  {32'h44ff12d9, 32'h00000000} /* (15, 4, 2) {real, imag} */,
  {32'h44f1edec, 32'h00000000} /* (15, 4, 1) {real, imag} */,
  {32'h44fa03ec, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'h4513e36e, 32'h00000000} /* (15, 3, 31) {real, imag} */,
  {32'h451613a0, 32'h00000000} /* (15, 3, 30) {real, imag} */,
  {32'h45215fc3, 32'h00000000} /* (15, 3, 29) {real, imag} */,
  {32'h453544a0, 32'h00000000} /* (15, 3, 28) {real, imag} */,
  {32'h4526e3d4, 32'h00000000} /* (15, 3, 27) {real, imag} */,
  {32'h4556ceb6, 32'h00000000} /* (15, 3, 26) {real, imag} */,
  {32'h451ff65f, 32'h00000000} /* (15, 3, 25) {real, imag} */,
  {32'h452f9636, 32'h00000000} /* (15, 3, 24) {real, imag} */,
  {32'h452aba90, 32'h00000000} /* (15, 3, 23) {real, imag} */,
  {32'h454c8792, 32'h00000000} /* (15, 3, 22) {real, imag} */,
  {32'h4512e768, 32'h00000000} /* (15, 3, 21) {real, imag} */,
  {32'h44f7fdf2, 32'h00000000} /* (15, 3, 20) {real, imag} */,
  {32'h44a7303f, 32'h00000000} /* (15, 3, 19) {real, imag} */,
  {32'h44c15dc2, 32'h00000000} /* (15, 3, 18) {real, imag} */,
  {32'h43e8cd14, 32'h00000000} /* (15, 3, 17) {real, imag} */,
  {32'h43d86220, 32'h00000000} /* (15, 3, 16) {real, imag} */,
  {32'hc4bca346, 32'h00000000} /* (15, 3, 15) {real, imag} */,
  {32'hc4af5c96, 32'h00000000} /* (15, 3, 14) {real, imag} */,
  {32'hc48960aa, 32'h00000000} /* (15, 3, 13) {real, imag} */,
  {32'hc49e3e6b, 32'h00000000} /* (15, 3, 12) {real, imag} */,
  {32'hc4506837, 32'h00000000} /* (15, 3, 11) {real, imag} */,
  {32'hc42ced16, 32'h00000000} /* (15, 3, 10) {real, imag} */,
  {32'hc490906a, 32'h00000000} /* (15, 3, 9) {real, imag} */,
  {32'hc40c0e7e, 32'h00000000} /* (15, 3, 8) {real, imag} */,
  {32'hc336ad40, 32'h00000000} /* (15, 3, 7) {real, imag} */,
  {32'h43b78290, 32'h00000000} /* (15, 3, 6) {real, imag} */,
  {32'h45002664, 32'h00000000} /* (15, 3, 5) {real, imag} */,
  {32'h4543969b, 32'h00000000} /* (15, 3, 4) {real, imag} */,
  {32'h4552c2f4, 32'h00000000} /* (15, 3, 3) {real, imag} */,
  {32'h44ced104, 32'h00000000} /* (15, 3, 2) {real, imag} */,
  {32'h44f50ea3, 32'h00000000} /* (15, 3, 1) {real, imag} */,
  {32'h450c4931, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'h44ff3713, 32'h00000000} /* (15, 2, 31) {real, imag} */,
  {32'h4555be75, 32'h00000000} /* (15, 2, 30) {real, imag} */,
  {32'h451b49da, 32'h00000000} /* (15, 2, 29) {real, imag} */,
  {32'h454314f7, 32'h00000000} /* (15, 2, 28) {real, imag} */,
  {32'h452c3182, 32'h00000000} /* (15, 2, 27) {real, imag} */,
  {32'h45325dbe, 32'h00000000} /* (15, 2, 26) {real, imag} */,
  {32'h4514fb6d, 32'h00000000} /* (15, 2, 25) {real, imag} */,
  {32'h453754aa, 32'h00000000} /* (15, 2, 24) {real, imag} */,
  {32'h4532b0b8, 32'h00000000} /* (15, 2, 23) {real, imag} */,
  {32'h4505dc86, 32'h00000000} /* (15, 2, 22) {real, imag} */,
  {32'h44f97b80, 32'h00000000} /* (15, 2, 21) {real, imag} */,
  {32'h44b0f931, 32'h00000000} /* (15, 2, 20) {real, imag} */,
  {32'h44de82bf, 32'h00000000} /* (15, 2, 19) {real, imag} */,
  {32'h447f398b, 32'h00000000} /* (15, 2, 18) {real, imag} */,
  {32'h4483e940, 32'h00000000} /* (15, 2, 17) {real, imag} */,
  {32'h44bb8388, 32'h00000000} /* (15, 2, 16) {real, imag} */,
  {32'hc43698da, 32'h00000000} /* (15, 2, 15) {real, imag} */,
  {32'hc4b56a4e, 32'h00000000} /* (15, 2, 14) {real, imag} */,
  {32'hc4b0d7d9, 32'h00000000} /* (15, 2, 13) {real, imag} */,
  {32'hc49d87aa, 32'h00000000} /* (15, 2, 12) {real, imag} */,
  {32'hc4d9089c, 32'h00000000} /* (15, 2, 11) {real, imag} */,
  {32'hc4826a70, 32'h00000000} /* (15, 2, 10) {real, imag} */,
  {32'hc475b383, 32'h00000000} /* (15, 2, 9) {real, imag} */,
  {32'hc3c88ca4, 32'h00000000} /* (15, 2, 8) {real, imag} */,
  {32'hc378dde8, 32'h00000000} /* (15, 2, 7) {real, imag} */,
  {32'h42e52618, 32'h00000000} /* (15, 2, 6) {real, imag} */,
  {32'h44f9b43e, 32'h00000000} /* (15, 2, 5) {real, imag} */,
  {32'h450e680c, 32'h00000000} /* (15, 2, 4) {real, imag} */,
  {32'h4514be00, 32'h00000000} /* (15, 2, 3) {real, imag} */,
  {32'h45233a2b, 32'h00000000} /* (15, 2, 2) {real, imag} */,
  {32'h44eb2b90, 32'h00000000} /* (15, 2, 1) {real, imag} */,
  {32'h45012899, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'h44e4350c, 32'h00000000} /* (15, 1, 31) {real, imag} */,
  {32'h451a78bc, 32'h00000000} /* (15, 1, 30) {real, imag} */,
  {32'h4514d45e, 32'h00000000} /* (15, 1, 29) {real, imag} */,
  {32'h4529c25a, 32'h00000000} /* (15, 1, 28) {real, imag} */,
  {32'h453a38d4, 32'h00000000} /* (15, 1, 27) {real, imag} */,
  {32'h451010be, 32'h00000000} /* (15, 1, 26) {real, imag} */,
  {32'h451f1af8, 32'h00000000} /* (15, 1, 25) {real, imag} */,
  {32'h450bf724, 32'h00000000} /* (15, 1, 24) {real, imag} */,
  {32'h45231e9a, 32'h00000000} /* (15, 1, 23) {real, imag} */,
  {32'h45314afa, 32'h00000000} /* (15, 1, 22) {real, imag} */,
  {32'h44da124a, 32'h00000000} /* (15, 1, 21) {real, imag} */,
  {32'h44e3e6db, 32'h00000000} /* (15, 1, 20) {real, imag} */,
  {32'h44c0f07c, 32'h00000000} /* (15, 1, 19) {real, imag} */,
  {32'h43695ccc, 32'h00000000} /* (15, 1, 18) {real, imag} */,
  {32'h446cd448, 32'h00000000} /* (15, 1, 17) {real, imag} */,
  {32'h4359c574, 32'h00000000} /* (15, 1, 16) {real, imag} */,
  {32'hc48f2e7c, 32'h00000000} /* (15, 1, 15) {real, imag} */,
  {32'hc4cf83f7, 32'h00000000} /* (15, 1, 14) {real, imag} */,
  {32'hc474f997, 32'h00000000} /* (15, 1, 13) {real, imag} */,
  {32'hc4a91e34, 32'h00000000} /* (15, 1, 12) {real, imag} */,
  {32'hc4adc37b, 32'h00000000} /* (15, 1, 11) {real, imag} */,
  {32'hc4e774e5, 32'h00000000} /* (15, 1, 10) {real, imag} */,
  {32'hc4bd5772, 32'h00000000} /* (15, 1, 9) {real, imag} */,
  {32'hc4a03c6a, 32'h00000000} /* (15, 1, 8) {real, imag} */,
  {32'hc41d6af6, 32'h00000000} /* (15, 1, 7) {real, imag} */,
  {32'hc4871889, 32'h00000000} /* (15, 1, 6) {real, imag} */,
  {32'hc3efd576, 32'h00000000} /* (15, 1, 5) {real, imag} */,
  {32'h449110a9, 32'h00000000} /* (15, 1, 4) {real, imag} */,
  {32'h44c711c2, 32'h00000000} /* (15, 1, 3) {real, imag} */,
  {32'h450bec64, 32'h00000000} /* (15, 1, 2) {real, imag} */,
  {32'h450346f6, 32'h00000000} /* (15, 1, 1) {real, imag} */,
  {32'h44a5517c, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'h44dbbbf5, 32'h00000000} /* (15, 0, 31) {real, imag} */,
  {32'h44e3ae33, 32'h00000000} /* (15, 0, 30) {real, imag} */,
  {32'h44f51e4a, 32'h00000000} /* (15, 0, 29) {real, imag} */,
  {32'h451f8dd4, 32'h00000000} /* (15, 0, 28) {real, imag} */,
  {32'h45080a74, 32'h00000000} /* (15, 0, 27) {real, imag} */,
  {32'h4513157a, 32'h00000000} /* (15, 0, 26) {real, imag} */,
  {32'h450c8388, 32'h00000000} /* (15, 0, 25) {real, imag} */,
  {32'h44fde2c7, 32'h00000000} /* (15, 0, 24) {real, imag} */,
  {32'h451fb5e6, 32'h00000000} /* (15, 0, 23) {real, imag} */,
  {32'h44ef3847, 32'h00000000} /* (15, 0, 22) {real, imag} */,
  {32'h44a1beb8, 32'h00000000} /* (15, 0, 21) {real, imag} */,
  {32'h446572eb, 32'h00000000} /* (15, 0, 20) {real, imag} */,
  {32'h44053adb, 32'h00000000} /* (15, 0, 19) {real, imag} */,
  {32'hc1b768c0, 32'h00000000} /* (15, 0, 18) {real, imag} */,
  {32'h431d65ec, 32'h00000000} /* (15, 0, 17) {real, imag} */,
  {32'hc22cfb40, 32'h00000000} /* (15, 0, 16) {real, imag} */,
  {32'hc46fbb6e, 32'h00000000} /* (15, 0, 15) {real, imag} */,
  {32'hc4c8bd31, 32'h00000000} /* (15, 0, 14) {real, imag} */,
  {32'hc4d01366, 32'h00000000} /* (15, 0, 13) {real, imag} */,
  {32'hc42d64a0, 32'h00000000} /* (15, 0, 12) {real, imag} */,
  {32'hc48e48db, 32'h00000000} /* (15, 0, 11) {real, imag} */,
  {32'hc49ecc0f, 32'h00000000} /* (15, 0, 10) {real, imag} */,
  {32'hc48a3b5a, 32'h00000000} /* (15, 0, 9) {real, imag} */,
  {32'hc430c8b6, 32'h00000000} /* (15, 0, 8) {real, imag} */,
  {32'hc3d8e550, 32'h00000000} /* (15, 0, 7) {real, imag} */,
  {32'hc39cbf64, 32'h00000000} /* (15, 0, 6) {real, imag} */,
  {32'h4412f785, 32'h00000000} /* (15, 0, 5) {real, imag} */,
  {32'h447d396d, 32'h00000000} /* (15, 0, 4) {real, imag} */,
  {32'h44d4c1e6, 32'h00000000} /* (15, 0, 3) {real, imag} */,
  {32'h4515f448, 32'h00000000} /* (15, 0, 2) {real, imag} */,
  {32'h44b9f838, 32'h00000000} /* (15, 0, 1) {real, imag} */,
  {32'h44a750b6, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h45afe6c3, 32'h00000000} /* (14, 31, 31) {real, imag} */,
  {32'h45b1b5b8, 32'h00000000} /* (14, 31, 30) {real, imag} */,
  {32'h45c4b0fb, 32'h00000000} /* (14, 31, 29) {real, imag} */,
  {32'h45c9b0ca, 32'h00000000} /* (14, 31, 28) {real, imag} */,
  {32'h45c71b43, 32'h00000000} /* (14, 31, 27) {real, imag} */,
  {32'h45ce142a, 32'h00000000} /* (14, 31, 26) {real, imag} */,
  {32'h45c5d998, 32'h00000000} /* (14, 31, 25) {real, imag} */,
  {32'h45d45eab, 32'h00000000} /* (14, 31, 24) {real, imag} */,
  {32'h459fc5ee, 32'h00000000} /* (14, 31, 23) {real, imag} */,
  {32'h4599bdce, 32'h00000000} /* (14, 31, 22) {real, imag} */,
  {32'h453f335a, 32'h00000000} /* (14, 31, 21) {real, imag} */,
  {32'h44da0819, 32'h00000000} /* (14, 31, 20) {real, imag} */,
  {32'h444d480c, 32'h00000000} /* (14, 31, 19) {real, imag} */,
  {32'hc4254dcc, 32'h00000000} /* (14, 31, 18) {real, imag} */,
  {32'hc4d812a6, 32'h00000000} /* (14, 31, 17) {real, imag} */,
  {32'hc4fe864b, 32'h00000000} /* (14, 31, 16) {real, imag} */,
  {32'hc5222732, 32'h00000000} /* (14, 31, 15) {real, imag} */,
  {32'hc540cef4, 32'h00000000} /* (14, 31, 14) {real, imag} */,
  {32'hc53949da, 32'h00000000} /* (14, 31, 13) {real, imag} */,
  {32'hc5182b03, 32'h00000000} /* (14, 31, 12) {real, imag} */,
  {32'hc5146a2a, 32'h00000000} /* (14, 31, 11) {real, imag} */,
  {32'hc4a07014, 32'h00000000} /* (14, 31, 10) {real, imag} */,
  {32'hc390dda8, 32'h00000000} /* (14, 31, 9) {real, imag} */,
  {32'h443f0218, 32'h00000000} /* (14, 31, 8) {real, imag} */,
  {32'h44cc6108, 32'h00000000} /* (14, 31, 7) {real, imag} */,
  {32'h4521f610, 32'h00000000} /* (14, 31, 6) {real, imag} */,
  {32'h455e1b2a, 32'h00000000} /* (14, 31, 5) {real, imag} */,
  {32'h45752402, 32'h00000000} /* (14, 31, 4) {real, imag} */,
  {32'h45889b02, 32'h00000000} /* (14, 31, 3) {real, imag} */,
  {32'h45a487cc, 32'h00000000} /* (14, 31, 2) {real, imag} */,
  {32'h45a82300, 32'h00000000} /* (14, 31, 1) {real, imag} */,
  {32'h45a355f9, 32'h00000000} /* (14, 31, 0) {real, imag} */,
  {32'h45accbb2, 32'h00000000} /* (14, 30, 31) {real, imag} */,
  {32'h45c5d202, 32'h00000000} /* (14, 30, 30) {real, imag} */,
  {32'h45c97a84, 32'h00000000} /* (14, 30, 29) {real, imag} */,
  {32'h45c89ff8, 32'h00000000} /* (14, 30, 28) {real, imag} */,
  {32'h45cede52, 32'h00000000} /* (14, 30, 27) {real, imag} */,
  {32'h46007d2c, 32'h00000000} /* (14, 30, 26) {real, imag} */,
  {32'h45e96046, 32'h00000000} /* (14, 30, 25) {real, imag} */,
  {32'h45f381f2, 32'h00000000} /* (14, 30, 24) {real, imag} */,
  {32'h45be4665, 32'h00000000} /* (14, 30, 23) {real, imag} */,
  {32'h4588ff7c, 32'h00000000} /* (14, 30, 22) {real, imag} */,
  {32'h4533f416, 32'h00000000} /* (14, 30, 21) {real, imag} */,
  {32'h446e4546, 32'h00000000} /* (14, 30, 20) {real, imag} */,
  {32'hc42a81f4, 32'h00000000} /* (14, 30, 19) {real, imag} */,
  {32'hc5419248, 32'h00000000} /* (14, 30, 18) {real, imag} */,
  {32'hc55c5908, 32'h00000000} /* (14, 30, 17) {real, imag} */,
  {32'hc5339908, 32'h00000000} /* (14, 30, 16) {real, imag} */,
  {32'hc5886e52, 32'h00000000} /* (14, 30, 15) {real, imag} */,
  {32'hc586a0fe, 32'h00000000} /* (14, 30, 14) {real, imag} */,
  {32'hc55df650, 32'h00000000} /* (14, 30, 13) {real, imag} */,
  {32'hc55337ff, 32'h00000000} /* (14, 30, 12) {real, imag} */,
  {32'hc5092c71, 32'h00000000} /* (14, 30, 11) {real, imag} */,
  {32'h424aa480, 32'h00000000} /* (14, 30, 10) {real, imag} */,
  {32'h44cd3f3e, 32'h00000000} /* (14, 30, 9) {real, imag} */,
  {32'h44cfe336, 32'h00000000} /* (14, 30, 8) {real, imag} */,
  {32'h4526f282, 32'h00000000} /* (14, 30, 7) {real, imag} */,
  {32'h455f9c5b, 32'h00000000} /* (14, 30, 6) {real, imag} */,
  {32'h45803d55, 32'h00000000} /* (14, 30, 5) {real, imag} */,
  {32'h458da4d8, 32'h00000000} /* (14, 30, 4) {real, imag} */,
  {32'h45963508, 32'h00000000} /* (14, 30, 3) {real, imag} */,
  {32'h4597fb26, 32'h00000000} /* (14, 30, 2) {real, imag} */,
  {32'h45b8d992, 32'h00000000} /* (14, 30, 1) {real, imag} */,
  {32'h45c4bf92, 32'h00000000} /* (14, 30, 0) {real, imag} */,
  {32'h45ae90aa, 32'h00000000} /* (14, 29, 31) {real, imag} */,
  {32'h45ca1c7e, 32'h00000000} /* (14, 29, 30) {real, imag} */,
  {32'h45c07866, 32'h00000000} /* (14, 29, 29) {real, imag} */,
  {32'h45cfbdb4, 32'h00000000} /* (14, 29, 28) {real, imag} */,
  {32'h45de207c, 32'h00000000} /* (14, 29, 27) {real, imag} */,
  {32'h45cdc2cb, 32'h00000000} /* (14, 29, 26) {real, imag} */,
  {32'h45c894d7, 32'h00000000} /* (14, 29, 25) {real, imag} */,
  {32'h45ba09b8, 32'h00000000} /* (14, 29, 24) {real, imag} */,
  {32'h45b7b58f, 32'h00000000} /* (14, 29, 23) {real, imag} */,
  {32'h455c54fb, 32'h00000000} /* (14, 29, 22) {real, imag} */,
  {32'h450ac01e, 32'h00000000} /* (14, 29, 21) {real, imag} */,
  {32'h4269c140, 32'h00000000} /* (14, 29, 20) {real, imag} */,
  {32'hc49f562e, 32'h00000000} /* (14, 29, 19) {real, imag} */,
  {32'hc5337cb6, 32'h00000000} /* (14, 29, 18) {real, imag} */,
  {32'hc552d6d6, 32'h00000000} /* (14, 29, 17) {real, imag} */,
  {32'hc581e3b7, 32'h00000000} /* (14, 29, 16) {real, imag} */,
  {32'hc5837712, 32'h00000000} /* (14, 29, 15) {real, imag} */,
  {32'hc56f4475, 32'h00000000} /* (14, 29, 14) {real, imag} */,
  {32'hc53a14f7, 32'h00000000} /* (14, 29, 13) {real, imag} */,
  {32'hc526d94b, 32'h00000000} /* (14, 29, 12) {real, imag} */,
  {32'hc4af30a8, 32'h00000000} /* (14, 29, 11) {real, imag} */,
  {32'h447594f8, 32'h00000000} /* (14, 29, 10) {real, imag} */,
  {32'h44d74d6c, 32'h00000000} /* (14, 29, 9) {real, imag} */,
  {32'h452b95d4, 32'h00000000} /* (14, 29, 8) {real, imag} */,
  {32'h454c2f2a, 32'h00000000} /* (14, 29, 7) {real, imag} */,
  {32'h4582ed74, 32'h00000000} /* (14, 29, 6) {real, imag} */,
  {32'h45b2611e, 32'h00000000} /* (14, 29, 5) {real, imag} */,
  {32'h45a3690a, 32'h00000000} /* (14, 29, 4) {real, imag} */,
  {32'h459b1062, 32'h00000000} /* (14, 29, 3) {real, imag} */,
  {32'h4594bdfa, 32'h00000000} /* (14, 29, 2) {real, imag} */,
  {32'h45d915cd, 32'h00000000} /* (14, 29, 1) {real, imag} */,
  {32'h45c25ecd, 32'h00000000} /* (14, 29, 0) {real, imag} */,
  {32'h45ad9c71, 32'h00000000} /* (14, 28, 31) {real, imag} */,
  {32'h45be8110, 32'h00000000} /* (14, 28, 30) {real, imag} */,
  {32'h45c501c4, 32'h00000000} /* (14, 28, 29) {real, imag} */,
  {32'h45dc54f0, 32'h00000000} /* (14, 28, 28) {real, imag} */,
  {32'h45dad48a, 32'h00000000} /* (14, 28, 27) {real, imag} */,
  {32'h45c7be7b, 32'h00000000} /* (14, 28, 26) {real, imag} */,
  {32'h45b39190, 32'h00000000} /* (14, 28, 25) {real, imag} */,
  {32'h45ae1244, 32'h00000000} /* (14, 28, 24) {real, imag} */,
  {32'h459bd35e, 32'h00000000} /* (14, 28, 23) {real, imag} */,
  {32'h45827aee, 32'h00000000} /* (14, 28, 22) {real, imag} */,
  {32'h4524399c, 32'h00000000} /* (14, 28, 21) {real, imag} */,
  {32'h4389f2a0, 32'h00000000} /* (14, 28, 20) {real, imag} */,
  {32'hc49f536c, 32'h00000000} /* (14, 28, 19) {real, imag} */,
  {32'hc549878b, 32'h00000000} /* (14, 28, 18) {real, imag} */,
  {32'hc584807e, 32'h00000000} /* (14, 28, 17) {real, imag} */,
  {32'hc598b53e, 32'h00000000} /* (14, 28, 16) {real, imag} */,
  {32'hc56e0eea, 32'h00000000} /* (14, 28, 15) {real, imag} */,
  {32'hc56b0adf, 32'h00000000} /* (14, 28, 14) {real, imag} */,
  {32'hc537f97b, 32'h00000000} /* (14, 28, 13) {real, imag} */,
  {32'hc4d29122, 32'h00000000} /* (14, 28, 12) {real, imag} */,
  {32'hc4b4f710, 32'h00000000} /* (14, 28, 11) {real, imag} */,
  {32'h44377d20, 32'h00000000} /* (14, 28, 10) {real, imag} */,
  {32'h455e0813, 32'h00000000} /* (14, 28, 9) {real, imag} */,
  {32'h456dc91c, 32'h00000000} /* (14, 28, 8) {real, imag} */,
  {32'h4573d2fc, 32'h00000000} /* (14, 28, 7) {real, imag} */,
  {32'h459f81ee, 32'h00000000} /* (14, 28, 6) {real, imag} */,
  {32'h45aeb4d6, 32'h00000000} /* (14, 28, 5) {real, imag} */,
  {32'h459ff3a5, 32'h00000000} /* (14, 28, 4) {real, imag} */,
  {32'h45a0d065, 32'h00000000} /* (14, 28, 3) {real, imag} */,
  {32'h45a41344, 32'h00000000} /* (14, 28, 2) {real, imag} */,
  {32'h45acee1a, 32'h00000000} /* (14, 28, 1) {real, imag} */,
  {32'h45ae51e2, 32'h00000000} /* (14, 28, 0) {real, imag} */,
  {32'h45a55db4, 32'h00000000} /* (14, 27, 31) {real, imag} */,
  {32'h45dab152, 32'h00000000} /* (14, 27, 30) {real, imag} */,
  {32'h45e41fec, 32'h00000000} /* (14, 27, 29) {real, imag} */,
  {32'h45d4900f, 32'h00000000} /* (14, 27, 28) {real, imag} */,
  {32'h45c30150, 32'h00000000} /* (14, 27, 27) {real, imag} */,
  {32'h45c8faec, 32'h00000000} /* (14, 27, 26) {real, imag} */,
  {32'h45b1934c, 32'h00000000} /* (14, 27, 25) {real, imag} */,
  {32'h45b983d7, 32'h00000000} /* (14, 27, 24) {real, imag} */,
  {32'h4595f644, 32'h00000000} /* (14, 27, 23) {real, imag} */,
  {32'h4599262c, 32'h00000000} /* (14, 27, 22) {real, imag} */,
  {32'h45537f3e, 32'h00000000} /* (14, 27, 21) {real, imag} */,
  {32'h42739ac0, 32'h00000000} /* (14, 27, 20) {real, imag} */,
  {32'hc4e43ca2, 32'h00000000} /* (14, 27, 19) {real, imag} */,
  {32'hc5496ff0, 32'h00000000} /* (14, 27, 18) {real, imag} */,
  {32'hc5726fba, 32'h00000000} /* (14, 27, 17) {real, imag} */,
  {32'hc5896ffe, 32'h00000000} /* (14, 27, 16) {real, imag} */,
  {32'hc55d296c, 32'h00000000} /* (14, 27, 15) {real, imag} */,
  {32'hc58322ac, 32'h00000000} /* (14, 27, 14) {real, imag} */,
  {32'hc53814a8, 32'h00000000} /* (14, 27, 13) {real, imag} */,
  {32'hc4fe2b54, 32'h00000000} /* (14, 27, 12) {real, imag} */,
  {32'hc556663b, 32'h00000000} /* (14, 27, 11) {real, imag} */,
  {32'h44196abc, 32'h00000000} /* (14, 27, 10) {real, imag} */,
  {32'h454a4ad1, 32'h00000000} /* (14, 27, 9) {real, imag} */,
  {32'h45860f81, 32'h00000000} /* (14, 27, 8) {real, imag} */,
  {32'h45928ec6, 32'h00000000} /* (14, 27, 7) {real, imag} */,
  {32'h45bc128e, 32'h00000000} /* (14, 27, 6) {real, imag} */,
  {32'h45b05739, 32'h00000000} /* (14, 27, 5) {real, imag} */,
  {32'h45a0f93c, 32'h00000000} /* (14, 27, 4) {real, imag} */,
  {32'h459a902e, 32'h00000000} /* (14, 27, 3) {real, imag} */,
  {32'h45af3484, 32'h00000000} /* (14, 27, 2) {real, imag} */,
  {32'h4599e141, 32'h00000000} /* (14, 27, 1) {real, imag} */,
  {32'h45963b72, 32'h00000000} /* (14, 27, 0) {real, imag} */,
  {32'h459310fa, 32'h00000000} /* (14, 26, 31) {real, imag} */,
  {32'h45ab4500, 32'h00000000} /* (14, 26, 30) {real, imag} */,
  {32'h45cd6cc0, 32'h00000000} /* (14, 26, 29) {real, imag} */,
  {32'h45e42fc8, 32'h00000000} /* (14, 26, 28) {real, imag} */,
  {32'h45cb6598, 32'h00000000} /* (14, 26, 27) {real, imag} */,
  {32'h45b4b00a, 32'h00000000} /* (14, 26, 26) {real, imag} */,
  {32'h45c93639, 32'h00000000} /* (14, 26, 25) {real, imag} */,
  {32'h45a9d935, 32'h00000000} /* (14, 26, 24) {real, imag} */,
  {32'h457ddaec, 32'h00000000} /* (14, 26, 23) {real, imag} */,
  {32'h4565c258, 32'h00000000} /* (14, 26, 22) {real, imag} */,
  {32'h450b7b46, 32'h00000000} /* (14, 26, 21) {real, imag} */,
  {32'hc4145424, 32'h00000000} /* (14, 26, 20) {real, imag} */,
  {32'hc4fd748e, 32'h00000000} /* (14, 26, 19) {real, imag} */,
  {32'hc55fb147, 32'h00000000} /* (14, 26, 18) {real, imag} */,
  {32'hc575674c, 32'h00000000} /* (14, 26, 17) {real, imag} */,
  {32'hc5ace0d4, 32'h00000000} /* (14, 26, 16) {real, imag} */,
  {32'hc581c55e, 32'h00000000} /* (14, 26, 15) {real, imag} */,
  {32'hc58798d8, 32'h00000000} /* (14, 26, 14) {real, imag} */,
  {32'hc5770210, 32'h00000000} /* (14, 26, 13) {real, imag} */,
  {32'hc52f00ab, 32'h00000000} /* (14, 26, 12) {real, imag} */,
  {32'hc5009ff7, 32'h00000000} /* (14, 26, 11) {real, imag} */,
  {32'h444d19bc, 32'h00000000} /* (14, 26, 10) {real, imag} */,
  {32'h44f4303c, 32'h00000000} /* (14, 26, 9) {real, imag} */,
  {32'h458474e9, 32'h00000000} /* (14, 26, 8) {real, imag} */,
  {32'h45b67aee, 32'h00000000} /* (14, 26, 7) {real, imag} */,
  {32'h45c69d90, 32'h00000000} /* (14, 26, 6) {real, imag} */,
  {32'h45acb3fb, 32'h00000000} /* (14, 26, 5) {real, imag} */,
  {32'h45a62746, 32'h00000000} /* (14, 26, 4) {real, imag} */,
  {32'h45b0be42, 32'h00000000} /* (14, 26, 3) {real, imag} */,
  {32'h45b3ad4e, 32'h00000000} /* (14, 26, 2) {real, imag} */,
  {32'h45a391ec, 32'h00000000} /* (14, 26, 1) {real, imag} */,
  {32'h45a18842, 32'h00000000} /* (14, 26, 0) {real, imag} */,
  {32'h45941e8c, 32'h00000000} /* (14, 25, 31) {real, imag} */,
  {32'h45bc960f, 32'h00000000} /* (14, 25, 30) {real, imag} */,
  {32'h45b59138, 32'h00000000} /* (14, 25, 29) {real, imag} */,
  {32'h45cdbb40, 32'h00000000} /* (14, 25, 28) {real, imag} */,
  {32'h45caa4a4, 32'h00000000} /* (14, 25, 27) {real, imag} */,
  {32'h45a6f77e, 32'h00000000} /* (14, 25, 26) {real, imag} */,
  {32'h45b99f13, 32'h00000000} /* (14, 25, 25) {real, imag} */,
  {32'h45add0a0, 32'h00000000} /* (14, 25, 24) {real, imag} */,
  {32'h458a445e, 32'h00000000} /* (14, 25, 23) {real, imag} */,
  {32'h45768e54, 32'h00000000} /* (14, 25, 22) {real, imag} */,
  {32'h450e3680, 32'h00000000} /* (14, 25, 21) {real, imag} */,
  {32'hc476665c, 32'h00000000} /* (14, 25, 20) {real, imag} */,
  {32'hc550f738, 32'h00000000} /* (14, 25, 19) {real, imag} */,
  {32'hc56cd009, 32'h00000000} /* (14, 25, 18) {real, imag} */,
  {32'hc597e141, 32'h00000000} /* (14, 25, 17) {real, imag} */,
  {32'hc5aaa538, 32'h00000000} /* (14, 25, 16) {real, imag} */,
  {32'hc596936e, 32'h00000000} /* (14, 25, 15) {real, imag} */,
  {32'hc58f541d, 32'h00000000} /* (14, 25, 14) {real, imag} */,
  {32'hc5955128, 32'h00000000} /* (14, 25, 13) {real, imag} */,
  {32'hc5810c76, 32'h00000000} /* (14, 25, 12) {real, imag} */,
  {32'hc4744ea0, 32'h00000000} /* (14, 25, 11) {real, imag} */,
  {32'h4484b4ce, 32'h00000000} /* (14, 25, 10) {real, imag} */,
  {32'h45368536, 32'h00000000} /* (14, 25, 9) {real, imag} */,
  {32'h455f9317, 32'h00000000} /* (14, 25, 8) {real, imag} */,
  {32'h4592e34a, 32'h00000000} /* (14, 25, 7) {real, imag} */,
  {32'h45a4bc66, 32'h00000000} /* (14, 25, 6) {real, imag} */,
  {32'h45b38f09, 32'h00000000} /* (14, 25, 5) {real, imag} */,
  {32'h45a08f04, 32'h00000000} /* (14, 25, 4) {real, imag} */,
  {32'h45ab1264, 32'h00000000} /* (14, 25, 3) {real, imag} */,
  {32'h45a2180a, 32'h00000000} /* (14, 25, 2) {real, imag} */,
  {32'h45b10eab, 32'h00000000} /* (14, 25, 1) {real, imag} */,
  {32'h458e8a1e, 32'h00000000} /* (14, 25, 0) {real, imag} */,
  {32'h45ab583b, 32'h00000000} /* (14, 24, 31) {real, imag} */,
  {32'h45964c28, 32'h00000000} /* (14, 24, 30) {real, imag} */,
  {32'h45a8c2db, 32'h00000000} /* (14, 24, 29) {real, imag} */,
  {32'h45c4efa9, 32'h00000000} /* (14, 24, 28) {real, imag} */,
  {32'h45a0eff7, 32'h00000000} /* (14, 24, 27) {real, imag} */,
  {32'h45815861, 32'h00000000} /* (14, 24, 26) {real, imag} */,
  {32'h4580b7c7, 32'h00000000} /* (14, 24, 25) {real, imag} */,
  {32'h459fde19, 32'h00000000} /* (14, 24, 24) {real, imag} */,
  {32'h4583342d, 32'h00000000} /* (14, 24, 23) {real, imag} */,
  {32'h457f93bc, 32'h00000000} /* (14, 24, 22) {real, imag} */,
  {32'h44afdb97, 32'h00000000} /* (14, 24, 21) {real, imag} */,
  {32'hc437a240, 32'h00000000} /* (14, 24, 20) {real, imag} */,
  {32'hc51a1ea6, 32'h00000000} /* (14, 24, 19) {real, imag} */,
  {32'hc54db524, 32'h00000000} /* (14, 24, 18) {real, imag} */,
  {32'hc58ec822, 32'h00000000} /* (14, 24, 17) {real, imag} */,
  {32'hc5a339c7, 32'h00000000} /* (14, 24, 16) {real, imag} */,
  {32'hc5946791, 32'h00000000} /* (14, 24, 15) {real, imag} */,
  {32'hc58d7814, 32'h00000000} /* (14, 24, 14) {real, imag} */,
  {32'hc592c763, 32'h00000000} /* (14, 24, 13) {real, imag} */,
  {32'hc57f9a7a, 32'h00000000} /* (14, 24, 12) {real, imag} */,
  {32'hc52c8e86, 32'h00000000} /* (14, 24, 11) {real, imag} */,
  {32'h4246fa60, 32'h00000000} /* (14, 24, 10) {real, imag} */,
  {32'h454456ea, 32'h00000000} /* (14, 24, 9) {real, imag} */,
  {32'h45932f65, 32'h00000000} /* (14, 24, 8) {real, imag} */,
  {32'h4594487d, 32'h00000000} /* (14, 24, 7) {real, imag} */,
  {32'h458b147e, 32'h00000000} /* (14, 24, 6) {real, imag} */,
  {32'h45905c62, 32'h00000000} /* (14, 24, 5) {real, imag} */,
  {32'h45a70ff1, 32'h00000000} /* (14, 24, 4) {real, imag} */,
  {32'h45abd3eb, 32'h00000000} /* (14, 24, 3) {real, imag} */,
  {32'h45817d52, 32'h00000000} /* (14, 24, 2) {real, imag} */,
  {32'h459bc6b2, 32'h00000000} /* (14, 24, 1) {real, imag} */,
  {32'h45694a32, 32'h00000000} /* (14, 24, 0) {real, imag} */,
  {32'h456121ae, 32'h00000000} /* (14, 23, 31) {real, imag} */,
  {32'h458b7bef, 32'h00000000} /* (14, 23, 30) {real, imag} */,
  {32'h4587b16e, 32'h00000000} /* (14, 23, 29) {real, imag} */,
  {32'h4594c14b, 32'h00000000} /* (14, 23, 28) {real, imag} */,
  {32'h4567ac18, 32'h00000000} /* (14, 23, 27) {real, imag} */,
  {32'h45664360, 32'h00000000} /* (14, 23, 26) {real, imag} */,
  {32'h4553842a, 32'h00000000} /* (14, 23, 25) {real, imag} */,
  {32'h455196a1, 32'h00000000} /* (14, 23, 24) {real, imag} */,
  {32'h455e9ea6, 32'h00000000} /* (14, 23, 23) {real, imag} */,
  {32'h453aedae, 32'h00000000} /* (14, 23, 22) {real, imag} */,
  {32'h447410ce, 32'h00000000} /* (14, 23, 21) {real, imag} */,
  {32'hc4a48863, 32'h00000000} /* (14, 23, 20) {real, imag} */,
  {32'hc4f25e1e, 32'h00000000} /* (14, 23, 19) {real, imag} */,
  {32'hc5449836, 32'h00000000} /* (14, 23, 18) {real, imag} */,
  {32'hc583b212, 32'h00000000} /* (14, 23, 17) {real, imag} */,
  {32'hc58ff1db, 32'h00000000} /* (14, 23, 16) {real, imag} */,
  {32'hc567a826, 32'h00000000} /* (14, 23, 15) {real, imag} */,
  {32'hc58077ef, 32'h00000000} /* (14, 23, 14) {real, imag} */,
  {32'hc585b662, 32'h00000000} /* (14, 23, 13) {real, imag} */,
  {32'hc5471fe0, 32'h00000000} /* (14, 23, 12) {real, imag} */,
  {32'hc4bcd310, 32'h00000000} /* (14, 23, 11) {real, imag} */,
  {32'h42bf2d70, 32'h00000000} /* (14, 23, 10) {real, imag} */,
  {32'h4528c022, 32'h00000000} /* (14, 23, 9) {real, imag} */,
  {32'h456a0c2b, 32'h00000000} /* (14, 23, 8) {real, imag} */,
  {32'h45454c5e, 32'h00000000} /* (14, 23, 7) {real, imag} */,
  {32'h4575af2e, 32'h00000000} /* (14, 23, 6) {real, imag} */,
  {32'h4595780c, 32'h00000000} /* (14, 23, 5) {real, imag} */,
  {32'h455b7f2c, 32'h00000000} /* (14, 23, 4) {real, imag} */,
  {32'h456ecb15, 32'h00000000} /* (14, 23, 3) {real, imag} */,
  {32'h455646a8, 32'h00000000} /* (14, 23, 2) {real, imag} */,
  {32'h455fd624, 32'h00000000} /* (14, 23, 1) {real, imag} */,
  {32'h4577bd72, 32'h00000000} /* (14, 23, 0) {real, imag} */,
  {32'h452f8d9f, 32'h00000000} /* (14, 22, 31) {real, imag} */,
  {32'h456171fe, 32'h00000000} /* (14, 22, 30) {real, imag} */,
  {32'h4584763f, 32'h00000000} /* (14, 22, 29) {real, imag} */,
  {32'h4553df35, 32'h00000000} /* (14, 22, 28) {real, imag} */,
  {32'h45352757, 32'h00000000} /* (14, 22, 27) {real, imag} */,
  {32'h451ae45d, 32'h00000000} /* (14, 22, 26) {real, imag} */,
  {32'h4504cbb4, 32'h00000000} /* (14, 22, 25) {real, imag} */,
  {32'h4515b4b4, 32'h00000000} /* (14, 22, 24) {real, imag} */,
  {32'h4550b02a, 32'h00000000} /* (14, 22, 23) {real, imag} */,
  {32'h452266a0, 32'h00000000} /* (14, 22, 22) {real, imag} */,
  {32'h443fa278, 32'h00000000} /* (14, 22, 21) {real, imag} */,
  {32'hc4826100, 32'h00000000} /* (14, 22, 20) {real, imag} */,
  {32'hc4832430, 32'h00000000} /* (14, 22, 19) {real, imag} */,
  {32'hc50e6ed4, 32'h00000000} /* (14, 22, 18) {real, imag} */,
  {32'hc527ecce, 32'h00000000} /* (14, 22, 17) {real, imag} */,
  {32'hc511dabe, 32'h00000000} /* (14, 22, 16) {real, imag} */,
  {32'hc52c17c3, 32'h00000000} /* (14, 22, 15) {real, imag} */,
  {32'hc5115d00, 32'h00000000} /* (14, 22, 14) {real, imag} */,
  {32'hc515d044, 32'h00000000} /* (14, 22, 13) {real, imag} */,
  {32'hc50b7a6b, 32'h00000000} /* (14, 22, 12) {real, imag} */,
  {32'hc4ef317e, 32'h00000000} /* (14, 22, 11) {real, imag} */,
  {32'h44564ec0, 32'h00000000} /* (14, 22, 10) {real, imag} */,
  {32'h44b94659, 32'h00000000} /* (14, 22, 9) {real, imag} */,
  {32'h457d8adc, 32'h00000000} /* (14, 22, 8) {real, imag} */,
  {32'h452955e0, 32'h00000000} /* (14, 22, 7) {real, imag} */,
  {32'h452df192, 32'h00000000} /* (14, 22, 6) {real, imag} */,
  {32'h4579baa6, 32'h00000000} /* (14, 22, 5) {real, imag} */,
  {32'h45396a31, 32'h00000000} /* (14, 22, 4) {real, imag} */,
  {32'h44d89d14, 32'h00000000} /* (14, 22, 3) {real, imag} */,
  {32'h45474d14, 32'h00000000} /* (14, 22, 2) {real, imag} */,
  {32'h454572fa, 32'h00000000} /* (14, 22, 1) {real, imag} */,
  {32'h4516013c, 32'h00000000} /* (14, 22, 0) {real, imag} */,
  {32'h44aeb54c, 32'h00000000} /* (14, 21, 31) {real, imag} */,
  {32'h44a0e64c, 32'h00000000} /* (14, 21, 30) {real, imag} */,
  {32'h448b6410, 32'h00000000} /* (14, 21, 29) {real, imag} */,
  {32'h441cc87d, 32'h00000000} /* (14, 21, 28) {real, imag} */,
  {32'h441abd19, 32'h00000000} /* (14, 21, 27) {real, imag} */,
  {32'hc3c1108a, 32'h00000000} /* (14, 21, 26) {real, imag} */,
  {32'h43d68c2e, 32'h00000000} /* (14, 21, 25) {real, imag} */,
  {32'h44404c12, 32'h00000000} /* (14, 21, 24) {real, imag} */,
  {32'h44598577, 32'h00000000} /* (14, 21, 23) {real, imag} */,
  {32'h44fd53aa, 32'h00000000} /* (14, 21, 22) {real, imag} */,
  {32'h43bd20e9, 32'h00000000} /* (14, 21, 21) {real, imag} */,
  {32'h4383bf94, 32'h00000000} /* (14, 21, 20) {real, imag} */,
  {32'hc26a2780, 32'h00000000} /* (14, 21, 19) {real, imag} */,
  {32'hc42fda2d, 32'h00000000} /* (14, 21, 18) {real, imag} */,
  {32'hc39e6618, 32'h00000000} /* (14, 21, 17) {real, imag} */,
  {32'hc4085ab9, 32'h00000000} /* (14, 21, 16) {real, imag} */,
  {32'hc3ad2d76, 32'h00000000} /* (14, 21, 15) {real, imag} */,
  {32'hc4277c57, 32'h00000000} /* (14, 21, 14) {real, imag} */,
  {32'hc4163f1c, 32'h00000000} /* (14, 21, 13) {real, imag} */,
  {32'hc3bdb312, 32'h00000000} /* (14, 21, 12) {real, imag} */,
  {32'hc38aa702, 32'h00000000} /* (14, 21, 11) {real, imag} */,
  {32'hc2cfaebe, 32'h00000000} /* (14, 21, 10) {real, imag} */,
  {32'h44e6aa3c, 32'h00000000} /* (14, 21, 9) {real, imag} */,
  {32'h451f0366, 32'h00000000} /* (14, 21, 8) {real, imag} */,
  {32'h44c1429a, 32'h00000000} /* (14, 21, 7) {real, imag} */,
  {32'h448a66c2, 32'h00000000} /* (14, 21, 6) {real, imag} */,
  {32'h441da994, 32'h00000000} /* (14, 21, 5) {real, imag} */,
  {32'h44a9270b, 32'h00000000} /* (14, 21, 4) {real, imag} */,
  {32'h44d9c0e1, 32'h00000000} /* (14, 21, 3) {real, imag} */,
  {32'h442e4f21, 32'h00000000} /* (14, 21, 2) {real, imag} */,
  {32'h449ed30c, 32'h00000000} /* (14, 21, 1) {real, imag} */,
  {32'h446fbaff, 32'h00000000} /* (14, 21, 0) {real, imag} */,
  {32'hc48b583a, 32'h00000000} /* (14, 20, 31) {real, imag} */,
  {32'hc470993f, 32'h00000000} /* (14, 20, 30) {real, imag} */,
  {32'hc51b9030, 32'h00000000} /* (14, 20, 29) {real, imag} */,
  {32'hc5602a20, 32'h00000000} /* (14, 20, 28) {real, imag} */,
  {32'hc504871e, 32'h00000000} /* (14, 20, 27) {real, imag} */,
  {32'hc520c9c8, 32'h00000000} /* (14, 20, 26) {real, imag} */,
  {32'hc528e07d, 32'h00000000} /* (14, 20, 25) {real, imag} */,
  {32'hc4b509a3, 32'h00000000} /* (14, 20, 24) {real, imag} */,
  {32'hc4881a0c, 32'h00000000} /* (14, 20, 23) {real, imag} */,
  {32'hc4a3270b, 32'h00000000} /* (14, 20, 22) {real, imag} */,
  {32'hc2a06b20, 32'h00000000} /* (14, 20, 21) {real, imag} */,
  {32'h44a39625, 32'h00000000} /* (14, 20, 20) {real, imag} */,
  {32'h445382c7, 32'h00000000} /* (14, 20, 19) {real, imag} */,
  {32'h44e3e5cc, 32'h00000000} /* (14, 20, 18) {real, imag} */,
  {32'h44c68154, 32'h00000000} /* (14, 20, 17) {real, imag} */,
  {32'h451044c8, 32'h00000000} /* (14, 20, 16) {real, imag} */,
  {32'h44e82174, 32'h00000000} /* (14, 20, 15) {real, imag} */,
  {32'h44ef9686, 32'h00000000} /* (14, 20, 14) {real, imag} */,
  {32'h44cb27b4, 32'h00000000} /* (14, 20, 13) {real, imag} */,
  {32'h4450bb96, 32'h00000000} /* (14, 20, 12) {real, imag} */,
  {32'h44f43cac, 32'h00000000} /* (14, 20, 11) {real, imag} */,
  {32'hc42511a3, 32'h00000000} /* (14, 20, 10) {real, imag} */,
  {32'hc304e510, 32'h00000000} /* (14, 20, 9) {real, imag} */,
  {32'hc48b1833, 32'h00000000} /* (14, 20, 8) {real, imag} */,
  {32'hc4f42784, 32'h00000000} /* (14, 20, 7) {real, imag} */,
  {32'hc4c215b5, 32'h00000000} /* (14, 20, 6) {real, imag} */,
  {32'hc4c2e494, 32'h00000000} /* (14, 20, 5) {real, imag} */,
  {32'hc4a05ddb, 32'h00000000} /* (14, 20, 4) {real, imag} */,
  {32'hc4c338e0, 32'h00000000} /* (14, 20, 3) {real, imag} */,
  {32'hc50f9952, 32'h00000000} /* (14, 20, 2) {real, imag} */,
  {32'hc4d93c78, 32'h00000000} /* (14, 20, 1) {real, imag} */,
  {32'hc4ac0a6b, 32'h00000000} /* (14, 20, 0) {real, imag} */,
  {32'hc50e180a, 32'h00000000} /* (14, 19, 31) {real, imag} */,
  {32'hc52cef70, 32'h00000000} /* (14, 19, 30) {real, imag} */,
  {32'hc5436af4, 32'h00000000} /* (14, 19, 29) {real, imag} */,
  {32'hc54c36e0, 32'h00000000} /* (14, 19, 28) {real, imag} */,
  {32'hc58f5508, 32'h00000000} /* (14, 19, 27) {real, imag} */,
  {32'hc5825ad3, 32'h00000000} /* (14, 19, 26) {real, imag} */,
  {32'hc53cea1b, 32'h00000000} /* (14, 19, 25) {real, imag} */,
  {32'hc52eeac7, 32'h00000000} /* (14, 19, 24) {real, imag} */,
  {32'hc50fed2d, 32'h00000000} /* (14, 19, 23) {real, imag} */,
  {32'hc516fe57, 32'h00000000} /* (14, 19, 22) {real, imag} */,
  {32'hc2975230, 32'h00000000} /* (14, 19, 21) {real, imag} */,
  {32'h44bb9e68, 32'h00000000} /* (14, 19, 20) {real, imag} */,
  {32'h45215237, 32'h00000000} /* (14, 19, 19) {real, imag} */,
  {32'h45391eb6, 32'h00000000} /* (14, 19, 18) {real, imag} */,
  {32'h4525cf63, 32'h00000000} /* (14, 19, 17) {real, imag} */,
  {32'h452cfbc2, 32'h00000000} /* (14, 19, 16) {real, imag} */,
  {32'h45391bb0, 32'h00000000} /* (14, 19, 15) {real, imag} */,
  {32'h453b09ac, 32'h00000000} /* (14, 19, 14) {real, imag} */,
  {32'h453a2c44, 32'h00000000} /* (14, 19, 13) {real, imag} */,
  {32'h453930e2, 32'h00000000} /* (14, 19, 12) {real, imag} */,
  {32'h44f656a4, 32'h00000000} /* (14, 19, 11) {real, imag} */,
  {32'hc328c568, 32'h00000000} /* (14, 19, 10) {real, imag} */,
  {32'hc4b264fa, 32'h00000000} /* (14, 19, 9) {real, imag} */,
  {32'hc4d54ab2, 32'h00000000} /* (14, 19, 8) {real, imag} */,
  {32'hc5780f83, 32'h00000000} /* (14, 19, 7) {real, imag} */,
  {32'hc54ea9e9, 32'h00000000} /* (14, 19, 6) {real, imag} */,
  {32'hc5281ff4, 32'h00000000} /* (14, 19, 5) {real, imag} */,
  {32'hc54973f2, 32'h00000000} /* (14, 19, 4) {real, imag} */,
  {32'hc53eccf5, 32'h00000000} /* (14, 19, 3) {real, imag} */,
  {32'hc5219a64, 32'h00000000} /* (14, 19, 2) {real, imag} */,
  {32'hc51603fb, 32'h00000000} /* (14, 19, 1) {real, imag} */,
  {32'hc51940c6, 32'h00000000} /* (14, 19, 0) {real, imag} */,
  {32'hc5599d92, 32'h00000000} /* (14, 18, 31) {real, imag} */,
  {32'hc55ab64a, 32'h00000000} /* (14, 18, 30) {real, imag} */,
  {32'hc569e5bc, 32'h00000000} /* (14, 18, 29) {real, imag} */,
  {32'hc57268db, 32'h00000000} /* (14, 18, 28) {real, imag} */,
  {32'hc5862d76, 32'h00000000} /* (14, 18, 27) {real, imag} */,
  {32'hc58fe8be, 32'h00000000} /* (14, 18, 26) {real, imag} */,
  {32'hc563f928, 32'h00000000} /* (14, 18, 25) {real, imag} */,
  {32'hc56e3613, 32'h00000000} /* (14, 18, 24) {real, imag} */,
  {32'hc55b11c2, 32'h00000000} /* (14, 18, 23) {real, imag} */,
  {32'hc5154cfd, 32'h00000000} /* (14, 18, 22) {real, imag} */,
  {32'hc41aed48, 32'h00000000} /* (14, 18, 21) {real, imag} */,
  {32'h44b17554, 32'h00000000} /* (14, 18, 20) {real, imag} */,
  {32'h45341143, 32'h00000000} /* (14, 18, 19) {real, imag} */,
  {32'h45350496, 32'h00000000} /* (14, 18, 18) {real, imag} */,
  {32'h45460332, 32'h00000000} /* (14, 18, 17) {real, imag} */,
  {32'h45827c28, 32'h00000000} /* (14, 18, 16) {real, imag} */,
  {32'h45676cb0, 32'h00000000} /* (14, 18, 15) {real, imag} */,
  {32'h454ae8f6, 32'h00000000} /* (14, 18, 14) {real, imag} */,
  {32'h4570cdca, 32'h00000000} /* (14, 18, 13) {real, imag} */,
  {32'h452491e5, 32'h00000000} /* (14, 18, 12) {real, imag} */,
  {32'h4505755b, 32'h00000000} /* (14, 18, 11) {real, imag} */,
  {32'h42458ac0, 32'h00000000} /* (14, 18, 10) {real, imag} */,
  {32'hc4a70bd9, 32'h00000000} /* (14, 18, 9) {real, imag} */,
  {32'hc52174b1, 32'h00000000} /* (14, 18, 8) {real, imag} */,
  {32'hc54ae19e, 32'h00000000} /* (14, 18, 7) {real, imag} */,
  {32'hc58f378a, 32'h00000000} /* (14, 18, 6) {real, imag} */,
  {32'hc58da065, 32'h00000000} /* (14, 18, 5) {real, imag} */,
  {32'hc583e877, 32'h00000000} /* (14, 18, 4) {real, imag} */,
  {32'hc5868a9d, 32'h00000000} /* (14, 18, 3) {real, imag} */,
  {32'hc520a5a8, 32'h00000000} /* (14, 18, 2) {real, imag} */,
  {32'hc58ce793, 32'h00000000} /* (14, 18, 1) {real, imag} */,
  {32'hc55af12c, 32'h00000000} /* (14, 18, 0) {real, imag} */,
  {32'hc564acae, 32'h00000000} /* (14, 17, 31) {real, imag} */,
  {32'hc58b4ee6, 32'h00000000} /* (14, 17, 30) {real, imag} */,
  {32'hc58451f3, 32'h00000000} /* (14, 17, 29) {real, imag} */,
  {32'hc58efea4, 32'h00000000} /* (14, 17, 28) {real, imag} */,
  {32'hc5ac1034, 32'h00000000} /* (14, 17, 27) {real, imag} */,
  {32'hc595e541, 32'h00000000} /* (14, 17, 26) {real, imag} */,
  {32'hc5ab29bd, 32'h00000000} /* (14, 17, 25) {real, imag} */,
  {32'hc5827719, 32'h00000000} /* (14, 17, 24) {real, imag} */,
  {32'hc586d85e, 32'h00000000} /* (14, 17, 23) {real, imag} */,
  {32'hc542b97c, 32'h00000000} /* (14, 17, 22) {real, imag} */,
  {32'hc4702164, 32'h00000000} /* (14, 17, 21) {real, imag} */,
  {32'h44df00c3, 32'h00000000} /* (14, 17, 20) {real, imag} */,
  {32'h455e69e3, 32'h00000000} /* (14, 17, 19) {real, imag} */,
  {32'h4575276c, 32'h00000000} /* (14, 17, 18) {real, imag} */,
  {32'h455b9549, 32'h00000000} /* (14, 17, 17) {real, imag} */,
  {32'h457db64e, 32'h00000000} /* (14, 17, 16) {real, imag} */,
  {32'h456594ca, 32'h00000000} /* (14, 17, 15) {real, imag} */,
  {32'h455e92c9, 32'h00000000} /* (14, 17, 14) {real, imag} */,
  {32'h45609c58, 32'h00000000} /* (14, 17, 13) {real, imag} */,
  {32'h452b561c, 32'h00000000} /* (14, 17, 12) {real, imag} */,
  {32'h4482292a, 32'h00000000} /* (14, 17, 11) {real, imag} */,
  {32'hc495eb50, 32'h00000000} /* (14, 17, 10) {real, imag} */,
  {32'hc4f378c9, 32'h00000000} /* (14, 17, 9) {real, imag} */,
  {32'hc5386ade, 32'h00000000} /* (14, 17, 8) {real, imag} */,
  {32'hc5779fc4, 32'h00000000} /* (14, 17, 7) {real, imag} */,
  {32'hc5af4ac0, 32'h00000000} /* (14, 17, 6) {real, imag} */,
  {32'hc5c67c14, 32'h00000000} /* (14, 17, 5) {real, imag} */,
  {32'hc5a49805, 32'h00000000} /* (14, 17, 4) {real, imag} */,
  {32'hc57ec30f, 32'h00000000} /* (14, 17, 3) {real, imag} */,
  {32'hc5889368, 32'h00000000} /* (14, 17, 2) {real, imag} */,
  {32'hc59917f6, 32'h00000000} /* (14, 17, 1) {real, imag} */,
  {32'hc583cf85, 32'h00000000} /* (14, 17, 0) {real, imag} */,
  {32'hc5885c04, 32'h00000000} /* (14, 16, 31) {real, imag} */,
  {32'hc5995e00, 32'h00000000} /* (14, 16, 30) {real, imag} */,
  {32'hc5a4175c, 32'h00000000} /* (14, 16, 29) {real, imag} */,
  {32'hc5923c72, 32'h00000000} /* (14, 16, 28) {real, imag} */,
  {32'hc5b59c26, 32'h00000000} /* (14, 16, 27) {real, imag} */,
  {32'hc59e7338, 32'h00000000} /* (14, 16, 26) {real, imag} */,
  {32'hc58d50ea, 32'h00000000} /* (14, 16, 25) {real, imag} */,
  {32'hc5a9cc03, 32'h00000000} /* (14, 16, 24) {real, imag} */,
  {32'hc59f55f6, 32'h00000000} /* (14, 16, 23) {real, imag} */,
  {32'hc56eb400, 32'h00000000} /* (14, 16, 22) {real, imag} */,
  {32'hc453f244, 32'h00000000} /* (14, 16, 21) {real, imag} */,
  {32'h44edcb4b, 32'h00000000} /* (14, 16, 20) {real, imag} */,
  {32'h454fc2d7, 32'h00000000} /* (14, 16, 19) {real, imag} */,
  {32'h458dbad1, 32'h00000000} /* (14, 16, 18) {real, imag} */,
  {32'h45a4c06a, 32'h00000000} /* (14, 16, 17) {real, imag} */,
  {32'h459a6389, 32'h00000000} /* (14, 16, 16) {real, imag} */,
  {32'h45843ca0, 32'h00000000} /* (14, 16, 15) {real, imag} */,
  {32'h4587b306, 32'h00000000} /* (14, 16, 14) {real, imag} */,
  {32'h4564da81, 32'h00000000} /* (14, 16, 13) {real, imag} */,
  {32'h4546af0e, 32'h00000000} /* (14, 16, 12) {real, imag} */,
  {32'h452486a5, 32'h00000000} /* (14, 16, 11) {real, imag} */,
  {32'hc399e200, 32'h00000000} /* (14, 16, 10) {real, imag} */,
  {32'hc4abe6b6, 32'h00000000} /* (14, 16, 9) {real, imag} */,
  {32'hc545e30a, 32'h00000000} /* (14, 16, 8) {real, imag} */,
  {32'hc5a1b3e2, 32'h00000000} /* (14, 16, 7) {real, imag} */,
  {32'hc5941628, 32'h00000000} /* (14, 16, 6) {real, imag} */,
  {32'hc5a944a8, 32'h00000000} /* (14, 16, 5) {real, imag} */,
  {32'hc5b0c825, 32'h00000000} /* (14, 16, 4) {real, imag} */,
  {32'hc5929406, 32'h00000000} /* (14, 16, 3) {real, imag} */,
  {32'hc5a46777, 32'h00000000} /* (14, 16, 2) {real, imag} */,
  {32'hc58bbe2c, 32'h00000000} /* (14, 16, 1) {real, imag} */,
  {32'hc58276dd, 32'h00000000} /* (14, 16, 0) {real, imag} */,
  {32'hc586873e, 32'h00000000} /* (14, 15, 31) {real, imag} */,
  {32'hc5b8454a, 32'h00000000} /* (14, 15, 30) {real, imag} */,
  {32'hc5b86f0e, 32'h00000000} /* (14, 15, 29) {real, imag} */,
  {32'hc5b37518, 32'h00000000} /* (14, 15, 28) {real, imag} */,
  {32'hc5b53c30, 32'h00000000} /* (14, 15, 27) {real, imag} */,
  {32'hc5b9f63f, 32'h00000000} /* (14, 15, 26) {real, imag} */,
  {32'hc59af356, 32'h00000000} /* (14, 15, 25) {real, imag} */,
  {32'hc582a8a4, 32'h00000000} /* (14, 15, 24) {real, imag} */,
  {32'hc5c5d94f, 32'h00000000} /* (14, 15, 23) {real, imag} */,
  {32'hc57db52a, 32'h00000000} /* (14, 15, 22) {real, imag} */,
  {32'hc3964558, 32'h00000000} /* (14, 15, 21) {real, imag} */,
  {32'h44c1cc61, 32'h00000000} /* (14, 15, 20) {real, imag} */,
  {32'h4569ac1f, 32'h00000000} /* (14, 15, 19) {real, imag} */,
  {32'h4572858f, 32'h00000000} /* (14, 15, 18) {real, imag} */,
  {32'h45892464, 32'h00000000} /* (14, 15, 17) {real, imag} */,
  {32'h45b007fb, 32'h00000000} /* (14, 15, 16) {real, imag} */,
  {32'h459d744e, 32'h00000000} /* (14, 15, 15) {real, imag} */,
  {32'h45924308, 32'h00000000} /* (14, 15, 14) {real, imag} */,
  {32'h45505228, 32'h00000000} /* (14, 15, 13) {real, imag} */,
  {32'h453df22c, 32'h00000000} /* (14, 15, 12) {real, imag} */,
  {32'h452cd927, 32'h00000000} /* (14, 15, 11) {real, imag} */,
  {32'h43b3b700, 32'h00000000} /* (14, 15, 10) {real, imag} */,
  {32'hc487571c, 32'h00000000} /* (14, 15, 9) {real, imag} */,
  {32'hc54bfd71, 32'h00000000} /* (14, 15, 8) {real, imag} */,
  {32'hc59225a9, 32'h00000000} /* (14, 15, 7) {real, imag} */,
  {32'hc5b7bb17, 32'h00000000} /* (14, 15, 6) {real, imag} */,
  {32'hc5b6ec0e, 32'h00000000} /* (14, 15, 5) {real, imag} */,
  {32'hc58316c9, 32'h00000000} /* (14, 15, 4) {real, imag} */,
  {32'hc5977e22, 32'h00000000} /* (14, 15, 3) {real, imag} */,
  {32'hc5b5e5e4, 32'h00000000} /* (14, 15, 2) {real, imag} */,
  {32'hc59bdd66, 32'h00000000} /* (14, 15, 1) {real, imag} */,
  {32'hc59e9f1f, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'hc5952bf7, 32'h00000000} /* (14, 14, 31) {real, imag} */,
  {32'hc5a9a166, 32'h00000000} /* (14, 14, 30) {real, imag} */,
  {32'hc5c1bec9, 32'h00000000} /* (14, 14, 29) {real, imag} */,
  {32'hc5aff56a, 32'h00000000} /* (14, 14, 28) {real, imag} */,
  {32'hc5bcc336, 32'h00000000} /* (14, 14, 27) {real, imag} */,
  {32'hc58d15e8, 32'h00000000} /* (14, 14, 26) {real, imag} */,
  {32'hc574ab2e, 32'h00000000} /* (14, 14, 25) {real, imag} */,
  {32'hc56f3402, 32'h00000000} /* (14, 14, 24) {real, imag} */,
  {32'hc56fc7aa, 32'h00000000} /* (14, 14, 23) {real, imag} */,
  {32'hc52fbaa6, 32'h00000000} /* (14, 14, 22) {real, imag} */,
  {32'hc4193b08, 32'h00000000} /* (14, 14, 21) {real, imag} */,
  {32'h44f92d16, 32'h00000000} /* (14, 14, 20) {real, imag} */,
  {32'h4531e73f, 32'h00000000} /* (14, 14, 19) {real, imag} */,
  {32'h456b0e83, 32'h00000000} /* (14, 14, 18) {real, imag} */,
  {32'h459922e2, 32'h00000000} /* (14, 14, 17) {real, imag} */,
  {32'h45a2a1b6, 32'h00000000} /* (14, 14, 16) {real, imag} */,
  {32'h459796cb, 32'h00000000} /* (14, 14, 15) {real, imag} */,
  {32'h4580524a, 32'h00000000} /* (14, 14, 14) {real, imag} */,
  {32'h458524d9, 32'h00000000} /* (14, 14, 13) {real, imag} */,
  {32'h4546b96d, 32'h00000000} /* (14, 14, 12) {real, imag} */,
  {32'h452610eb, 32'h00000000} /* (14, 14, 11) {real, imag} */,
  {32'h4201e540, 32'h00000000} /* (14, 14, 10) {real, imag} */,
  {32'hc4b8469b, 32'h00000000} /* (14, 14, 9) {real, imag} */,
  {32'hc5135342, 32'h00000000} /* (14, 14, 8) {real, imag} */,
  {32'hc571c3ee, 32'h00000000} /* (14, 14, 7) {real, imag} */,
  {32'hc59cc05c, 32'h00000000} /* (14, 14, 6) {real, imag} */,
  {32'hc59065e2, 32'h00000000} /* (14, 14, 5) {real, imag} */,
  {32'hc59a93aa, 32'h00000000} /* (14, 14, 4) {real, imag} */,
  {32'hc5a0ac7c, 32'h00000000} /* (14, 14, 3) {real, imag} */,
  {32'hc59a7b44, 32'h00000000} /* (14, 14, 2) {real, imag} */,
  {32'hc59fdcea, 32'h00000000} /* (14, 14, 1) {real, imag} */,
  {32'hc5884782, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'hc5670afc, 32'h00000000} /* (14, 13, 31) {real, imag} */,
  {32'hc5a26783, 32'h00000000} /* (14, 13, 30) {real, imag} */,
  {32'hc5850ba1, 32'h00000000} /* (14, 13, 29) {real, imag} */,
  {32'hc59aca7a, 32'h00000000} /* (14, 13, 28) {real, imag} */,
  {32'hc59cf362, 32'h00000000} /* (14, 13, 27) {real, imag} */,
  {32'hc54c519a, 32'h00000000} /* (14, 13, 26) {real, imag} */,
  {32'hc546e295, 32'h00000000} /* (14, 13, 25) {real, imag} */,
  {32'hc551420e, 32'h00000000} /* (14, 13, 24) {real, imag} */,
  {32'hc50dbc4d, 32'h00000000} /* (14, 13, 23) {real, imag} */,
  {32'hc4ac5a62, 32'h00000000} /* (14, 13, 22) {real, imag} */,
  {32'hc407921c, 32'h00000000} /* (14, 13, 21) {real, imag} */,
  {32'h452c202b, 32'h00000000} /* (14, 13, 20) {real, imag} */,
  {32'h4549155e, 32'h00000000} /* (14, 13, 19) {real, imag} */,
  {32'h45759021, 32'h00000000} /* (14, 13, 18) {real, imag} */,
  {32'h458cbdb6, 32'h00000000} /* (14, 13, 17) {real, imag} */,
  {32'h45856974, 32'h00000000} /* (14, 13, 16) {real, imag} */,
  {32'h4580aef2, 32'h00000000} /* (14, 13, 15) {real, imag} */,
  {32'h4559eea7, 32'h00000000} /* (14, 13, 14) {real, imag} */,
  {32'h455f51fc, 32'h00000000} /* (14, 13, 13) {real, imag} */,
  {32'h4554aeb4, 32'h00000000} /* (14, 13, 12) {real, imag} */,
  {32'h45148286, 32'h00000000} /* (14, 13, 11) {real, imag} */,
  {32'h43e9a9b4, 32'h00000000} /* (14, 13, 10) {real, imag} */,
  {32'hc4a421fe, 32'h00000000} /* (14, 13, 9) {real, imag} */,
  {32'hc51c3f6e, 32'h00000000} /* (14, 13, 8) {real, imag} */,
  {32'hc5815dd8, 32'h00000000} /* (14, 13, 7) {real, imag} */,
  {32'hc585119e, 32'h00000000} /* (14, 13, 6) {real, imag} */,
  {32'hc55ef621, 32'h00000000} /* (14, 13, 5) {real, imag} */,
  {32'hc5630645, 32'h00000000} /* (14, 13, 4) {real, imag} */,
  {32'hc58e3089, 32'h00000000} /* (14, 13, 3) {real, imag} */,
  {32'hc56e7d8d, 32'h00000000} /* (14, 13, 2) {real, imag} */,
  {32'hc585c01e, 32'h00000000} /* (14, 13, 1) {real, imag} */,
  {32'hc5694c3d, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'hc52549e1, 32'h00000000} /* (14, 12, 31) {real, imag} */,
  {32'hc57f81e2, 32'h00000000} /* (14, 12, 30) {real, imag} */,
  {32'hc5714c22, 32'h00000000} /* (14, 12, 29) {real, imag} */,
  {32'hc55cbc1c, 32'h00000000} /* (14, 12, 28) {real, imag} */,
  {32'hc5397e47, 32'h00000000} /* (14, 12, 27) {real, imag} */,
  {32'hc5270180, 32'h00000000} /* (14, 12, 26) {real, imag} */,
  {32'hc506885a, 32'h00000000} /* (14, 12, 25) {real, imag} */,
  {32'hc5394daf, 32'h00000000} /* (14, 12, 24) {real, imag} */,
  {32'hc4c76111, 32'h00000000} /* (14, 12, 23) {real, imag} */,
  {32'hc4ca4968, 32'h00000000} /* (14, 12, 22) {real, imag} */,
  {32'h43284a5c, 32'h00000000} /* (14, 12, 21) {real, imag} */,
  {32'h45017d47, 32'h00000000} /* (14, 12, 20) {real, imag} */,
  {32'h45658e86, 32'h00000000} /* (14, 12, 19) {real, imag} */,
  {32'h45881505, 32'h00000000} /* (14, 12, 18) {real, imag} */,
  {32'h4585668d, 32'h00000000} /* (14, 12, 17) {real, imag} */,
  {32'h45438b2c, 32'h00000000} /* (14, 12, 16) {real, imag} */,
  {32'h4549f4a9, 32'h00000000} /* (14, 12, 15) {real, imag} */,
  {32'h45337666, 32'h00000000} /* (14, 12, 14) {real, imag} */,
  {32'h455b2a0a, 32'h00000000} /* (14, 12, 13) {real, imag} */,
  {32'h455b5f5a, 32'h00000000} /* (14, 12, 12) {real, imag} */,
  {32'h45001151, 32'h00000000} /* (14, 12, 11) {real, imag} */,
  {32'h43a06c0c, 32'h00000000} /* (14, 12, 10) {real, imag} */,
  {32'hc4739e3a, 32'h00000000} /* (14, 12, 9) {real, imag} */,
  {32'hc4de263a, 32'h00000000} /* (14, 12, 8) {real, imag} */,
  {32'hc52c7d38, 32'h00000000} /* (14, 12, 7) {real, imag} */,
  {32'hc52dff38, 32'h00000000} /* (14, 12, 6) {real, imag} */,
  {32'hc4eef974, 32'h00000000} /* (14, 12, 5) {real, imag} */,
  {32'hc51f070b, 32'h00000000} /* (14, 12, 4) {real, imag} */,
  {32'hc532f332, 32'h00000000} /* (14, 12, 3) {real, imag} */,
  {32'hc5412d1b, 32'h00000000} /* (14, 12, 2) {real, imag} */,
  {32'hc54bfcae, 32'h00000000} /* (14, 12, 1) {real, imag} */,
  {32'hc50463be, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'hc415abc8, 32'h00000000} /* (14, 11, 31) {real, imag} */,
  {32'hc3a68df6, 32'h00000000} /* (14, 11, 30) {real, imag} */,
  {32'hc5426ef1, 32'h00000000} /* (14, 11, 29) {real, imag} */,
  {32'hc4f4165b, 32'h00000000} /* (14, 11, 28) {real, imag} */,
  {32'hc46bbdf1, 32'h00000000} /* (14, 11, 27) {real, imag} */,
  {32'hc51c750d, 32'h00000000} /* (14, 11, 26) {real, imag} */,
  {32'hc46ba868, 32'h00000000} /* (14, 11, 25) {real, imag} */,
  {32'hc49ca259, 32'h00000000} /* (14, 11, 24) {real, imag} */,
  {32'hc49a8cd6, 32'h00000000} /* (14, 11, 23) {real, imag} */,
  {32'hc332be76, 32'h00000000} /* (14, 11, 22) {real, imag} */,
  {32'h4381d7ba, 32'h00000000} /* (14, 11, 21) {real, imag} */,
  {32'h44cc5f5c, 32'h00000000} /* (14, 11, 20) {real, imag} */,
  {32'h450bb6a1, 32'h00000000} /* (14, 11, 19) {real, imag} */,
  {32'h45063a86, 32'h00000000} /* (14, 11, 18) {real, imag} */,
  {32'h456c930c, 32'h00000000} /* (14, 11, 17) {real, imag} */,
  {32'h4537e054, 32'h00000000} /* (14, 11, 16) {real, imag} */,
  {32'h44ef411c, 32'h00000000} /* (14, 11, 15) {real, imag} */,
  {32'h44e77974, 32'h00000000} /* (14, 11, 14) {real, imag} */,
  {32'h450ca503, 32'h00000000} /* (14, 11, 13) {real, imag} */,
  {32'h45156b1c, 32'h00000000} /* (14, 11, 12) {real, imag} */,
  {32'h44bebe70, 32'h00000000} /* (14, 11, 11) {real, imag} */,
  {32'hc3993648, 32'h00000000} /* (14, 11, 10) {real, imag} */,
  {32'hc448767e, 32'h00000000} /* (14, 11, 9) {real, imag} */,
  {32'hc4a413c1, 32'h00000000} /* (14, 11, 8) {real, imag} */,
  {32'hc4c164ca, 32'h00000000} /* (14, 11, 7) {real, imag} */,
  {32'hc4902e44, 32'h00000000} /* (14, 11, 6) {real, imag} */,
  {32'hc41e5b15, 32'h00000000} /* (14, 11, 5) {real, imag} */,
  {32'hc498916c, 32'h00000000} /* (14, 11, 4) {real, imag} */,
  {32'hc4234451, 32'h00000000} /* (14, 11, 3) {real, imag} */,
  {32'hc3e42baa, 32'h00000000} /* (14, 11, 2) {real, imag} */,
  {32'hc489c60c, 32'h00000000} /* (14, 11, 1) {real, imag} */,
  {32'hc41c9444, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h44f4bace, 32'h00000000} /* (14, 10, 31) {real, imag} */,
  {32'h44989789, 32'h00000000} /* (14, 10, 30) {real, imag} */,
  {32'h456817d9, 32'h00000000} /* (14, 10, 29) {real, imag} */,
  {32'h44d2711a, 32'h00000000} /* (14, 10, 28) {real, imag} */,
  {32'h44a55efe, 32'h00000000} /* (14, 10, 27) {real, imag} */,
  {32'h44ba1103, 32'h00000000} /* (14, 10, 26) {real, imag} */,
  {32'h4475d782, 32'h00000000} /* (14, 10, 25) {real, imag} */,
  {32'h44bdd066, 32'h00000000} /* (14, 10, 24) {real, imag} */,
  {32'h449abbcf, 32'h00000000} /* (14, 10, 23) {real, imag} */,
  {32'h4500ece4, 32'h00000000} /* (14, 10, 22) {real, imag} */,
  {32'h448c5454, 32'h00000000} /* (14, 10, 21) {real, imag} */,
  {32'h44002077, 32'h00000000} /* (14, 10, 20) {real, imag} */,
  {32'h441bd5e0, 32'h00000000} /* (14, 10, 19) {real, imag} */,
  {32'hc346ddc8, 32'h00000000} /* (14, 10, 18) {real, imag} */,
  {32'h4353ff98, 32'h00000000} /* (14, 10, 17) {real, imag} */,
  {32'h4411b147, 32'h00000000} /* (14, 10, 16) {real, imag} */,
  {32'h3f88b600, 32'h00000000} /* (14, 10, 15) {real, imag} */,
  {32'hc35cbb08, 32'h00000000} /* (14, 10, 14) {real, imag} */,
  {32'hc44ece7c, 32'h00000000} /* (14, 10, 13) {real, imag} */,
  {32'h4291c528, 32'h00000000} /* (14, 10, 12) {real, imag} */,
  {32'hc2384810, 32'h00000000} /* (14, 10, 11) {real, imag} */,
  {32'hc21993a0, 32'h00000000} /* (14, 10, 10) {real, imag} */,
  {32'hc328e146, 32'h00000000} /* (14, 10, 9) {real, imag} */,
  {32'h4457ba58, 32'h00000000} /* (14, 10, 8) {real, imag} */,
  {32'h43591050, 32'h00000000} /* (14, 10, 7) {real, imag} */,
  {32'h43e2b40c, 32'h00000000} /* (14, 10, 6) {real, imag} */,
  {32'h44914458, 32'h00000000} /* (14, 10, 5) {real, imag} */,
  {32'h44dd8730, 32'h00000000} /* (14, 10, 4) {real, imag} */,
  {32'h450da7ae, 32'h00000000} /* (14, 10, 3) {real, imag} */,
  {32'h4527f90c, 32'h00000000} /* (14, 10, 2) {real, imag} */,
  {32'h451d6c02, 32'h00000000} /* (14, 10, 1) {real, imag} */,
  {32'h449e7182, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'h44eb6e35, 32'h00000000} /* (14, 9, 31) {real, imag} */,
  {32'h4548c85f, 32'h00000000} /* (14, 9, 30) {real, imag} */,
  {32'h457c08de, 32'h00000000} /* (14, 9, 29) {real, imag} */,
  {32'h4568c44c, 32'h00000000} /* (14, 9, 28) {real, imag} */,
  {32'h457eedf2, 32'h00000000} /* (14, 9, 27) {real, imag} */,
  {32'h458f32a4, 32'h00000000} /* (14, 9, 26) {real, imag} */,
  {32'h45518486, 32'h00000000} /* (14, 9, 25) {real, imag} */,
  {32'h45687928, 32'h00000000} /* (14, 9, 24) {real, imag} */,
  {32'h4531facc, 32'h00000000} /* (14, 9, 23) {real, imag} */,
  {32'h452d6d5b, 32'h00000000} /* (14, 9, 22) {real, imag} */,
  {32'h455e6f94, 32'h00000000} /* (14, 9, 21) {real, imag} */,
  {32'h43cbe580, 32'h00000000} /* (14, 9, 20) {real, imag} */,
  {32'hc3ea4170, 32'h00000000} /* (14, 9, 19) {real, imag} */,
  {32'hc507b8a1, 32'h00000000} /* (14, 9, 18) {real, imag} */,
  {32'hc4b4d6dd, 32'h00000000} /* (14, 9, 17) {real, imag} */,
  {32'hc4444368, 32'h00000000} /* (14, 9, 16) {real, imag} */,
  {32'hc4afc0cb, 32'h00000000} /* (14, 9, 15) {real, imag} */,
  {32'hc4cdab42, 32'h00000000} /* (14, 9, 14) {real, imag} */,
  {32'hc4aface0, 32'h00000000} /* (14, 9, 13) {real, imag} */,
  {32'hc49e04f5, 32'h00000000} /* (14, 9, 12) {real, imag} */,
  {32'hc46639a8, 32'h00000000} /* (14, 9, 11) {real, imag} */,
  {32'h4439c258, 32'h00000000} /* (14, 9, 10) {real, imag} */,
  {32'h446a31d0, 32'h00000000} /* (14, 9, 9) {real, imag} */,
  {32'h44f36783, 32'h00000000} /* (14, 9, 8) {real, imag} */,
  {32'h45033558, 32'h00000000} /* (14, 9, 7) {real, imag} */,
  {32'h450d0dcf, 32'h00000000} /* (14, 9, 6) {real, imag} */,
  {32'h45307f7e, 32'h00000000} /* (14, 9, 5) {real, imag} */,
  {32'h4569d558, 32'h00000000} /* (14, 9, 4) {real, imag} */,
  {32'h4570d9e2, 32'h00000000} /* (14, 9, 3) {real, imag} */,
  {32'h45839b40, 32'h00000000} /* (14, 9, 2) {real, imag} */,
  {32'h456c8e00, 32'h00000000} /* (14, 9, 1) {real, imag} */,
  {32'h454137f2, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'h4566f46e, 32'h00000000} /* (14, 8, 31) {real, imag} */,
  {32'h456c66cb, 32'h00000000} /* (14, 8, 30) {real, imag} */,
  {32'h456c5812, 32'h00000000} /* (14, 8, 29) {real, imag} */,
  {32'h458cb990, 32'h00000000} /* (14, 8, 28) {real, imag} */,
  {32'h45747224, 32'h00000000} /* (14, 8, 27) {real, imag} */,
  {32'h458676a2, 32'h00000000} /* (14, 8, 26) {real, imag} */,
  {32'h45999070, 32'h00000000} /* (14, 8, 25) {real, imag} */,
  {32'h45abef8c, 32'h00000000} /* (14, 8, 24) {real, imag} */,
  {32'h45801187, 32'h00000000} /* (14, 8, 23) {real, imag} */,
  {32'h4586c1f3, 32'h00000000} /* (14, 8, 22) {real, imag} */,
  {32'h4502f2bd, 32'h00000000} /* (14, 8, 21) {real, imag} */,
  {32'h4462150a, 32'h00000000} /* (14, 8, 20) {real, imag} */,
  {32'hc4201036, 32'h00000000} /* (14, 8, 19) {real, imag} */,
  {32'hc48d804e, 32'h00000000} /* (14, 8, 18) {real, imag} */,
  {32'hc48baf80, 32'h00000000} /* (14, 8, 17) {real, imag} */,
  {32'hc4e9f294, 32'h00000000} /* (14, 8, 16) {real, imag} */,
  {32'hc50e628e, 32'h00000000} /* (14, 8, 15) {real, imag} */,
  {32'hc513a639, 32'h00000000} /* (14, 8, 14) {real, imag} */,
  {32'hc51ebbc6, 32'h00000000} /* (14, 8, 13) {real, imag} */,
  {32'hc4bcc353, 32'h00000000} /* (14, 8, 12) {real, imag} */,
  {32'hc4aedd75, 32'h00000000} /* (14, 8, 11) {real, imag} */,
  {32'h43b98c58, 32'h00000000} /* (14, 8, 10) {real, imag} */,
  {32'h44b3eca6, 32'h00000000} /* (14, 8, 9) {real, imag} */,
  {32'h44ddd0d4, 32'h00000000} /* (14, 8, 8) {real, imag} */,
  {32'h454f5395, 32'h00000000} /* (14, 8, 7) {real, imag} */,
  {32'h457a370a, 32'h00000000} /* (14, 8, 6) {real, imag} */,
  {32'h459b4370, 32'h00000000} /* (14, 8, 5) {real, imag} */,
  {32'h453dafba, 32'h00000000} /* (14, 8, 4) {real, imag} */,
  {32'h4584ba1f, 32'h00000000} /* (14, 8, 3) {real, imag} */,
  {32'h459807f2, 32'h00000000} /* (14, 8, 2) {real, imag} */,
  {32'h45951853, 32'h00000000} /* (14, 8, 1) {real, imag} */,
  {32'h453bafe0, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'h457fbb7f, 32'h00000000} /* (14, 7, 31) {real, imag} */,
  {32'h4590141e, 32'h00000000} /* (14, 7, 30) {real, imag} */,
  {32'h458d9d74, 32'h00000000} /* (14, 7, 29) {real, imag} */,
  {32'h459c330d, 32'h00000000} /* (14, 7, 28) {real, imag} */,
  {32'h4594c77e, 32'h00000000} /* (14, 7, 27) {real, imag} */,
  {32'h45b07d14, 32'h00000000} /* (14, 7, 26) {real, imag} */,
  {32'h45a13d7e, 32'h00000000} /* (14, 7, 25) {real, imag} */,
  {32'h45ac94e5, 32'h00000000} /* (14, 7, 24) {real, imag} */,
  {32'h4596cd83, 32'h00000000} /* (14, 7, 23) {real, imag} */,
  {32'h45a39486, 32'h00000000} /* (14, 7, 22) {real, imag} */,
  {32'h45257961, 32'h00000000} /* (14, 7, 21) {real, imag} */,
  {32'h42dc6150, 32'h00000000} /* (14, 7, 20) {real, imag} */,
  {32'h428ec700, 32'h00000000} /* (14, 7, 19) {real, imag} */,
  {32'hc487f58c, 32'h00000000} /* (14, 7, 18) {real, imag} */,
  {32'hc4f47e61, 32'h00000000} /* (14, 7, 17) {real, imag} */,
  {32'hc4dc392e, 32'h00000000} /* (14, 7, 16) {real, imag} */,
  {32'hc5115e2b, 32'h00000000} /* (14, 7, 15) {real, imag} */,
  {32'hc543c535, 32'h00000000} /* (14, 7, 14) {real, imag} */,
  {32'hc54c2101, 32'h00000000} /* (14, 7, 13) {real, imag} */,
  {32'hc4f13677, 32'h00000000} /* (14, 7, 12) {real, imag} */,
  {32'hc4cd50d8, 32'h00000000} /* (14, 7, 11) {real, imag} */,
  {32'h43d5b1f8, 32'h00000000} /* (14, 7, 10) {real, imag} */,
  {32'h448f5546, 32'h00000000} /* (14, 7, 9) {real, imag} */,
  {32'h450ed1bc, 32'h00000000} /* (14, 7, 8) {real, imag} */,
  {32'h45731032, 32'h00000000} /* (14, 7, 7) {real, imag} */,
  {32'h4583880a, 32'h00000000} /* (14, 7, 6) {real, imag} */,
  {32'h459196d4, 32'h00000000} /* (14, 7, 5) {real, imag} */,
  {32'h45792a4e, 32'h00000000} /* (14, 7, 4) {real, imag} */,
  {32'h458b71ca, 32'h00000000} /* (14, 7, 3) {real, imag} */,
  {32'h45a46506, 32'h00000000} /* (14, 7, 2) {real, imag} */,
  {32'h4586aac4, 32'h00000000} /* (14, 7, 1) {real, imag} */,
  {32'h4580ff3c, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'h458cfeb0, 32'h00000000} /* (14, 6, 31) {real, imag} */,
  {32'h458be6fd, 32'h00000000} /* (14, 6, 30) {real, imag} */,
  {32'h45a7164b, 32'h00000000} /* (14, 6, 29) {real, imag} */,
  {32'h45a0f02a, 32'h00000000} /* (14, 6, 28) {real, imag} */,
  {32'h45d2d238, 32'h00000000} /* (14, 6, 27) {real, imag} */,
  {32'h45cab1e8, 32'h00000000} /* (14, 6, 26) {real, imag} */,
  {32'h45b806f4, 32'h00000000} /* (14, 6, 25) {real, imag} */,
  {32'h45a44586, 32'h00000000} /* (14, 6, 24) {real, imag} */,
  {32'h45b484fc, 32'h00000000} /* (14, 6, 23) {real, imag} */,
  {32'h45a83f96, 32'h00000000} /* (14, 6, 22) {real, imag} */,
  {32'h45703420, 32'h00000000} /* (14, 6, 21) {real, imag} */,
  {32'h448a0dba, 32'h00000000} /* (14, 6, 20) {real, imag} */,
  {32'h436cad50, 32'h00000000} /* (14, 6, 19) {real, imag} */,
  {32'hc4533a94, 32'h00000000} /* (14, 6, 18) {real, imag} */,
  {32'hc4c2bab8, 32'h00000000} /* (14, 6, 17) {real, imag} */,
  {32'hc4a46bd7, 32'h00000000} /* (14, 6, 16) {real, imag} */,
  {32'hc51d5017, 32'h00000000} /* (14, 6, 15) {real, imag} */,
  {32'hc55467ba, 32'h00000000} /* (14, 6, 14) {real, imag} */,
  {32'hc54b48b6, 32'h00000000} /* (14, 6, 13) {real, imag} */,
  {32'hc5473790, 32'h00000000} /* (14, 6, 12) {real, imag} */,
  {32'hc51bf97f, 32'h00000000} /* (14, 6, 11) {real, imag} */,
  {32'hc468703c, 32'h00000000} /* (14, 6, 10) {real, imag} */,
  {32'h4469ed04, 32'h00000000} /* (14, 6, 9) {real, imag} */,
  {32'h4511528f, 32'h00000000} /* (14, 6, 8) {real, imag} */,
  {32'h452267a7, 32'h00000000} /* (14, 6, 7) {real, imag} */,
  {32'h455e7bcc, 32'h00000000} /* (14, 6, 6) {real, imag} */,
  {32'h45617118, 32'h00000000} /* (14, 6, 5) {real, imag} */,
  {32'h45b3bfb4, 32'h00000000} /* (14, 6, 4) {real, imag} */,
  {32'h45aeaaf0, 32'h00000000} /* (14, 6, 3) {real, imag} */,
  {32'h458dc422, 32'h00000000} /* (14, 6, 2) {real, imag} */,
  {32'h45bbb395, 32'h00000000} /* (14, 6, 1) {real, imag} */,
  {32'h4592a758, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h45991d56, 32'h00000000} /* (14, 5, 31) {real, imag} */,
  {32'h45b160bc, 32'h00000000} /* (14, 5, 30) {real, imag} */,
  {32'h45b787b5, 32'h00000000} /* (14, 5, 29) {real, imag} */,
  {32'h45d5d43f, 32'h00000000} /* (14, 5, 28) {real, imag} */,
  {32'h45d5308f, 32'h00000000} /* (14, 5, 27) {real, imag} */,
  {32'h45c3a032, 32'h00000000} /* (14, 5, 26) {real, imag} */,
  {32'h45b10952, 32'h00000000} /* (14, 5, 25) {real, imag} */,
  {32'h45cbe0e4, 32'h00000000} /* (14, 5, 24) {real, imag} */,
  {32'h45b41f92, 32'h00000000} /* (14, 5, 23) {real, imag} */,
  {32'h45c21635, 32'h00000000} /* (14, 5, 22) {real, imag} */,
  {32'h45a00315, 32'h00000000} /* (14, 5, 21) {real, imag} */,
  {32'h454e6249, 32'h00000000} /* (14, 5, 20) {real, imag} */,
  {32'h44ccc972, 32'h00000000} /* (14, 5, 19) {real, imag} */,
  {32'h4400aab8, 32'h00000000} /* (14, 5, 18) {real, imag} */,
  {32'hc2966360, 32'h00000000} /* (14, 5, 17) {real, imag} */,
  {32'hc3d7ca08, 32'h00000000} /* (14, 5, 16) {real, imag} */,
  {32'hc50ef5c9, 32'h00000000} /* (14, 5, 15) {real, imag} */,
  {32'hc5784c37, 32'h00000000} /* (14, 5, 14) {real, imag} */,
  {32'hc55af2f2, 32'h00000000} /* (14, 5, 13) {real, imag} */,
  {32'hc543b0c6, 32'h00000000} /* (14, 5, 12) {real, imag} */,
  {32'hc53e3d7e, 32'h00000000} /* (14, 5, 11) {real, imag} */,
  {32'hc5363ef4, 32'h00000000} /* (14, 5, 10) {real, imag} */,
  {32'hc505cdac, 32'h00000000} /* (14, 5, 9) {real, imag} */,
  {32'hc46ea0cc, 32'h00000000} /* (14, 5, 8) {real, imag} */,
  {32'h43c9e4b0, 32'h00000000} /* (14, 5, 7) {real, imag} */,
  {32'h44f1d508, 32'h00000000} /* (14, 5, 6) {real, imag} */,
  {32'h455e8c16, 32'h00000000} /* (14, 5, 5) {real, imag} */,
  {32'h45846117, 32'h00000000} /* (14, 5, 4) {real, imag} */,
  {32'h45b4e5de, 32'h00000000} /* (14, 5, 3) {real, imag} */,
  {32'h45b592b1, 32'h00000000} /* (14, 5, 2) {real, imag} */,
  {32'h459e3e1e, 32'h00000000} /* (14, 5, 1) {real, imag} */,
  {32'h459ca0b6, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'h45a9319e, 32'h00000000} /* (14, 4, 31) {real, imag} */,
  {32'h45c612e7, 32'h00000000} /* (14, 4, 30) {real, imag} */,
  {32'h45d3ada4, 32'h00000000} /* (14, 4, 29) {real, imag} */,
  {32'h45e4f475, 32'h00000000} /* (14, 4, 28) {real, imag} */,
  {32'h45e1f066, 32'h00000000} /* (14, 4, 27) {real, imag} */,
  {32'h45d91a3e, 32'h00000000} /* (14, 4, 26) {real, imag} */,
  {32'h45d2545f, 32'h00000000} /* (14, 4, 25) {real, imag} */,
  {32'h45d79503, 32'h00000000} /* (14, 4, 24) {real, imag} */,
  {32'h45d38c58, 32'h00000000} /* (14, 4, 23) {real, imag} */,
  {32'h45de60e9, 32'h00000000} /* (14, 4, 22) {real, imag} */,
  {32'h45c9d04f, 32'h00000000} /* (14, 4, 21) {real, imag} */,
  {32'h459ab89b, 32'h00000000} /* (14, 4, 20) {real, imag} */,
  {32'h453b3896, 32'h00000000} /* (14, 4, 19) {real, imag} */,
  {32'h44e62d74, 32'h00000000} /* (14, 4, 18) {real, imag} */,
  {32'h44b6bb00, 32'h00000000} /* (14, 4, 17) {real, imag} */,
  {32'h43d52b50, 32'h00000000} /* (14, 4, 16) {real, imag} */,
  {32'hc4aa2512, 32'h00000000} /* (14, 4, 15) {real, imag} */,
  {32'hc52e0526, 32'h00000000} /* (14, 4, 14) {real, imag} */,
  {32'hc55734d7, 32'h00000000} /* (14, 4, 13) {real, imag} */,
  {32'hc5453c5e, 32'h00000000} /* (14, 4, 12) {real, imag} */,
  {32'hc5428304, 32'h00000000} /* (14, 4, 11) {real, imag} */,
  {32'hc547524c, 32'h00000000} /* (14, 4, 10) {real, imag} */,
  {32'hc5732ff2, 32'h00000000} /* (14, 4, 9) {real, imag} */,
  {32'hc4fca434, 32'h00000000} /* (14, 4, 8) {real, imag} */,
  {32'hc4156464, 32'h00000000} /* (14, 4, 7) {real, imag} */,
  {32'h4472fcd8, 32'h00000000} /* (14, 4, 6) {real, imag} */,
  {32'h45318b92, 32'h00000000} /* (14, 4, 5) {real, imag} */,
  {32'h458749e3, 32'h00000000} /* (14, 4, 4) {real, imag} */,
  {32'h45afa927, 32'h00000000} /* (14, 4, 3) {real, imag} */,
  {32'h45c52e8f, 32'h00000000} /* (14, 4, 2) {real, imag} */,
  {32'h45abfa3e, 32'h00000000} /* (14, 4, 1) {real, imag} */,
  {32'h45a129b5, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'h45d427cb, 32'h00000000} /* (14, 3, 31) {real, imag} */,
  {32'h45c044ec, 32'h00000000} /* (14, 3, 30) {real, imag} */,
  {32'h45c8c79a, 32'h00000000} /* (14, 3, 29) {real, imag} */,
  {32'h45dc9476, 32'h00000000} /* (14, 3, 28) {real, imag} */,
  {32'h46055b64, 32'h00000000} /* (14, 3, 27) {real, imag} */,
  {32'h45ddf748, 32'h00000000} /* (14, 3, 26) {real, imag} */,
  {32'h45d98c31, 32'h00000000} /* (14, 3, 25) {real, imag} */,
  {32'h45e33f60, 32'h00000000} /* (14, 3, 24) {real, imag} */,
  {32'h45d55964, 32'h00000000} /* (14, 3, 23) {real, imag} */,
  {32'h45de0c17, 32'h00000000} /* (14, 3, 22) {real, imag} */,
  {32'h45b9aa54, 32'h00000000} /* (14, 3, 21) {real, imag} */,
  {32'h45a43f4e, 32'h00000000} /* (14, 3, 20) {real, imag} */,
  {32'h455503f9, 32'h00000000} /* (14, 3, 19) {real, imag} */,
  {32'h4579cb55, 32'h00000000} /* (14, 3, 18) {real, imag} */,
  {32'h44d330b8, 32'h00000000} /* (14, 3, 17) {real, imag} */,
  {32'h4446de88, 32'h00000000} /* (14, 3, 16) {real, imag} */,
  {32'hc4bd89e4, 32'h00000000} /* (14, 3, 15) {real, imag} */,
  {32'hc51eb58f, 32'h00000000} /* (14, 3, 14) {real, imag} */,
  {32'hc552a1ec, 32'h00000000} /* (14, 3, 13) {real, imag} */,
  {32'hc56531ec, 32'h00000000} /* (14, 3, 12) {real, imag} */,
  {32'hc5617276, 32'h00000000} /* (14, 3, 11) {real, imag} */,
  {32'hc5512ac5, 32'h00000000} /* (14, 3, 10) {real, imag} */,
  {32'hc51cbfe6, 32'h00000000} /* (14, 3, 9) {real, imag} */,
  {32'hc507a774, 32'h00000000} /* (14, 3, 8) {real, imag} */,
  {32'hc3eaa6c0, 32'h00000000} /* (14, 3, 7) {real, imag} */,
  {32'h44215e20, 32'h00000000} /* (14, 3, 6) {real, imag} */,
  {32'h4554b9ad, 32'h00000000} /* (14, 3, 5) {real, imag} */,
  {32'h45986e2a, 32'h00000000} /* (14, 3, 4) {real, imag} */,
  {32'h45ab5524, 32'h00000000} /* (14, 3, 3) {real, imag} */,
  {32'h45a9ea26, 32'h00000000} /* (14, 3, 2) {real, imag} */,
  {32'h45a61276, 32'h00000000} /* (14, 3, 1) {real, imag} */,
  {32'h45aef315, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h45c6ca84, 32'h00000000} /* (14, 2, 31) {real, imag} */,
  {32'h45def0da, 32'h00000000} /* (14, 2, 30) {real, imag} */,
  {32'h45bf45d6, 32'h00000000} /* (14, 2, 29) {real, imag} */,
  {32'h45de2fa0, 32'h00000000} /* (14, 2, 28) {real, imag} */,
  {32'h45ddfe0a, 32'h00000000} /* (14, 2, 27) {real, imag} */,
  {32'h45d4f6ef, 32'h00000000} /* (14, 2, 26) {real, imag} */,
  {32'h45d34e1c, 32'h00000000} /* (14, 2, 25) {real, imag} */,
  {32'h45da2252, 32'h00000000} /* (14, 2, 24) {real, imag} */,
  {32'h45d32f1d, 32'h00000000} /* (14, 2, 23) {real, imag} */,
  {32'h45b5879a, 32'h00000000} /* (14, 2, 22) {real, imag} */,
  {32'h45b3236f, 32'h00000000} /* (14, 2, 21) {real, imag} */,
  {32'h458044ff, 32'h00000000} /* (14, 2, 20) {real, imag} */,
  {32'h455e8638, 32'h00000000} /* (14, 2, 19) {real, imag} */,
  {32'h4524bd58, 32'h00000000} /* (14, 2, 18) {real, imag} */,
  {32'h4503c80a, 32'h00000000} /* (14, 2, 17) {real, imag} */,
  {32'h441c0cd0, 32'h00000000} /* (14, 2, 16) {real, imag} */,
  {32'hc5058944, 32'h00000000} /* (14, 2, 15) {real, imag} */,
  {32'hc4f9e146, 32'h00000000} /* (14, 2, 14) {real, imag} */,
  {32'hc55bb63c, 32'h00000000} /* (14, 2, 13) {real, imag} */,
  {32'hc57f4718, 32'h00000000} /* (14, 2, 12) {real, imag} */,
  {32'hc548109d, 32'h00000000} /* (14, 2, 11) {real, imag} */,
  {32'hc52eb2de, 32'h00000000} /* (14, 2, 10) {real, imag} */,
  {32'hc5472fdc, 32'h00000000} /* (14, 2, 9) {real, imag} */,
  {32'hc4d10050, 32'h00000000} /* (14, 2, 8) {real, imag} */,
  {32'hc48543e4, 32'h00000000} /* (14, 2, 7) {real, imag} */,
  {32'h431dea90, 32'h00000000} /* (14, 2, 6) {real, imag} */,
  {32'h44f7acdd, 32'h00000000} /* (14, 2, 5) {real, imag} */,
  {32'h45899dad, 32'h00000000} /* (14, 2, 4) {real, imag} */,
  {32'h45cb61cc, 32'h00000000} /* (14, 2, 3) {real, imag} */,
  {32'h45b85464, 32'h00000000} /* (14, 2, 2) {real, imag} */,
  {32'h45a768af, 32'h00000000} /* (14, 2, 1) {real, imag} */,
  {32'h45a11058, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h45a87b34, 32'h00000000} /* (14, 1, 31) {real, imag} */,
  {32'h45ce7fef, 32'h00000000} /* (14, 1, 30) {real, imag} */,
  {32'h45dae557, 32'h00000000} /* (14, 1, 29) {real, imag} */,
  {32'h45ecaf1b, 32'h00000000} /* (14, 1, 28) {real, imag} */,
  {32'h45ddbe9c, 32'h00000000} /* (14, 1, 27) {real, imag} */,
  {32'h45d16b1f, 32'h00000000} /* (14, 1, 26) {real, imag} */,
  {32'h45d9d6d0, 32'h00000000} /* (14, 1, 25) {real, imag} */,
  {32'h45e66032, 32'h00000000} /* (14, 1, 24) {real, imag} */,
  {32'h45a51428, 32'h00000000} /* (14, 1, 23) {real, imag} */,
  {32'h45b45af3, 32'h00000000} /* (14, 1, 22) {real, imag} */,
  {32'h4594bcdc, 32'h00000000} /* (14, 1, 21) {real, imag} */,
  {32'h4565447d, 32'h00000000} /* (14, 1, 20) {real, imag} */,
  {32'h455824d0, 32'h00000000} /* (14, 1, 19) {real, imag} */,
  {32'h44f8519b, 32'h00000000} /* (14, 1, 18) {real, imag} */,
  {32'h449882fe, 32'h00000000} /* (14, 1, 17) {real, imag} */,
  {32'h42540980, 32'h00000000} /* (14, 1, 16) {real, imag} */,
  {32'hc4b804da, 32'h00000000} /* (14, 1, 15) {real, imag} */,
  {32'hc52579ce, 32'h00000000} /* (14, 1, 14) {real, imag} */,
  {32'hc5789dea, 32'h00000000} /* (14, 1, 13) {real, imag} */,
  {32'hc56001ca, 32'h00000000} /* (14, 1, 12) {real, imag} */,
  {32'hc54a12b0, 32'h00000000} /* (14, 1, 11) {real, imag} */,
  {32'hc56c219a, 32'h00000000} /* (14, 1, 10) {real, imag} */,
  {32'hc5354617, 32'h00000000} /* (14, 1, 9) {real, imag} */,
  {32'hc514532c, 32'h00000000} /* (14, 1, 8) {real, imag} */,
  {32'hc4680564, 32'h00000000} /* (14, 1, 7) {real, imag} */,
  {32'h43b3ac30, 32'h00000000} /* (14, 1, 6) {real, imag} */,
  {32'h4528ffb4, 32'h00000000} /* (14, 1, 5) {real, imag} */,
  {32'h456af7ef, 32'h00000000} /* (14, 1, 4) {real, imag} */,
  {32'h45996cba, 32'h00000000} /* (14, 1, 3) {real, imag} */,
  {32'h45b4eb85, 32'h00000000} /* (14, 1, 2) {real, imag} */,
  {32'h4597e494, 32'h00000000} /* (14, 1, 1) {real, imag} */,
  {32'h459a8bf9, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h45a3d16b, 32'h00000000} /* (14, 0, 31) {real, imag} */,
  {32'h45b7114a, 32'h00000000} /* (14, 0, 30) {real, imag} */,
  {32'h45c75188, 32'h00000000} /* (14, 0, 29) {real, imag} */,
  {32'h45cdac92, 32'h00000000} /* (14, 0, 28) {real, imag} */,
  {32'h45e9250e, 32'h00000000} /* (14, 0, 27) {real, imag} */,
  {32'h45cf0e0a, 32'h00000000} /* (14, 0, 26) {real, imag} */,
  {32'h45c3ba0e, 32'h00000000} /* (14, 0, 25) {real, imag} */,
  {32'h45afda04, 32'h00000000} /* (14, 0, 24) {real, imag} */,
  {32'h45ad8390, 32'h00000000} /* (14, 0, 23) {real, imag} */,
  {32'h4590fb8d, 32'h00000000} /* (14, 0, 22) {real, imag} */,
  {32'h4560f2e9, 32'h00000000} /* (14, 0, 21) {real, imag} */,
  {32'h453f70e1, 32'h00000000} /* (14, 0, 20) {real, imag} */,
  {32'h44e7df82, 32'h00000000} /* (14, 0, 19) {real, imag} */,
  {32'h44ba042b, 32'h00000000} /* (14, 0, 18) {real, imag} */,
  {32'hc36b2410, 32'h00000000} /* (14, 0, 17) {real, imag} */,
  {32'hc44d3192, 32'h00000000} /* (14, 0, 16) {real, imag} */,
  {32'hc4faad8f, 32'h00000000} /* (14, 0, 15) {real, imag} */,
  {32'hc551df38, 32'h00000000} /* (14, 0, 14) {real, imag} */,
  {32'hc55f7de0, 32'h00000000} /* (14, 0, 13) {real, imag} */,
  {32'hc5489437, 32'h00000000} /* (14, 0, 12) {real, imag} */,
  {32'hc528b111, 32'h00000000} /* (14, 0, 11) {real, imag} */,
  {32'hc511f1a4, 32'h00000000} /* (14, 0, 10) {real, imag} */,
  {32'hc49ac036, 32'h00000000} /* (14, 0, 9) {real, imag} */,
  {32'hc4b46574, 32'h00000000} /* (14, 0, 8) {real, imag} */,
  {32'hc3c45518, 32'h00000000} /* (14, 0, 7) {real, imag} */,
  {32'h44936f6d, 32'h00000000} /* (14, 0, 6) {real, imag} */,
  {32'h4520dd83, 32'h00000000} /* (14, 0, 5) {real, imag} */,
  {32'h45666b51, 32'h00000000} /* (14, 0, 4) {real, imag} */,
  {32'h4591c224, 32'h00000000} /* (14, 0, 3) {real, imag} */,
  {32'h458e0c23, 32'h00000000} /* (14, 0, 2) {real, imag} */,
  {32'h458fa91a, 32'h00000000} /* (14, 0, 1) {real, imag} */,
  {32'h4595f487, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h4602f99e, 32'h00000000} /* (13, 31, 31) {real, imag} */,
  {32'h462018d0, 32'h00000000} /* (13, 31, 30) {real, imag} */,
  {32'h46182a7c, 32'h00000000} /* (13, 31, 29) {real, imag} */,
  {32'h46140f86, 32'h00000000} /* (13, 31, 28) {real, imag} */,
  {32'h4616175c, 32'h00000000} /* (13, 31, 27) {real, imag} */,
  {32'h4625b9d9, 32'h00000000} /* (13, 31, 26) {real, imag} */,
  {32'h46110fee, 32'h00000000} /* (13, 31, 25) {real, imag} */,
  {32'h4609d1f6, 32'h00000000} /* (13, 31, 24) {real, imag} */,
  {32'h45f85342, 32'h00000000} /* (13, 31, 23) {real, imag} */,
  {32'h45c0c942, 32'h00000000} /* (13, 31, 22) {real, imag} */,
  {32'h458c6310, 32'h00000000} /* (13, 31, 21) {real, imag} */,
  {32'h45188bdd, 32'h00000000} /* (13, 31, 20) {real, imag} */,
  {32'h446c9a84, 32'h00000000} /* (13, 31, 19) {real, imag} */,
  {32'hc4507d40, 32'h00000000} /* (13, 31, 18) {real, imag} */,
  {32'hc513692b, 32'h00000000} /* (13, 31, 17) {real, imag} */,
  {32'hc52e8c69, 32'h00000000} /* (13, 31, 16) {real, imag} */,
  {32'hc573e4ca, 32'h00000000} /* (13, 31, 15) {real, imag} */,
  {32'hc59008a1, 32'h00000000} /* (13, 31, 14) {real, imag} */,
  {32'hc597115c, 32'h00000000} /* (13, 31, 13) {real, imag} */,
  {32'hc564c952, 32'h00000000} /* (13, 31, 12) {real, imag} */,
  {32'hc5184a58, 32'h00000000} /* (13, 31, 11) {real, imag} */,
  {32'hc45de2b0, 32'h00000000} /* (13, 31, 10) {real, imag} */,
  {32'h43df1c10, 32'h00000000} /* (13, 31, 9) {real, imag} */,
  {32'h445e0c64, 32'h00000000} /* (13, 31, 8) {real, imag} */,
  {32'h4523f678, 32'h00000000} /* (13, 31, 7) {real, imag} */,
  {32'h458a9cea, 32'h00000000} /* (13, 31, 6) {real, imag} */,
  {32'h45c88cc0, 32'h00000000} /* (13, 31, 5) {real, imag} */,
  {32'h45d9a7dc, 32'h00000000} /* (13, 31, 4) {real, imag} */,
  {32'h45d34ba2, 32'h00000000} /* (13, 31, 3) {real, imag} */,
  {32'h45e3f494, 32'h00000000} /* (13, 31, 2) {real, imag} */,
  {32'h45f1678a, 32'h00000000} /* (13, 31, 1) {real, imag} */,
  {32'h45f2874e, 32'h00000000} /* (13, 31, 0) {real, imag} */,
  {32'h460e2d46, 32'h00000000} /* (13, 30, 31) {real, imag} */,
  {32'h4612a30d, 32'h00000000} /* (13, 30, 30) {real, imag} */,
  {32'h46179db2, 32'h00000000} /* (13, 30, 29) {real, imag} */,
  {32'h4616c9b4, 32'h00000000} /* (13, 30, 28) {real, imag} */,
  {32'h461704ce, 32'h00000000} /* (13, 30, 27) {real, imag} */,
  {32'h46168b56, 32'h00000000} /* (13, 30, 26) {real, imag} */,
  {32'h46256b52, 32'h00000000} /* (13, 30, 25) {real, imag} */,
  {32'h4613de9e, 32'h00000000} /* (13, 30, 24) {real, imag} */,
  {32'h46007250, 32'h00000000} /* (13, 30, 23) {real, imag} */,
  {32'h45e92de6, 32'h00000000} /* (13, 30, 22) {real, imag} */,
  {32'h455ed31d, 32'h00000000} /* (13, 30, 21) {real, imag} */,
  {32'h43c8f0f8, 32'h00000000} /* (13, 30, 20) {real, imag} */,
  {32'hc4589af8, 32'h00000000} /* (13, 30, 19) {real, imag} */,
  {32'hc53a316b, 32'h00000000} /* (13, 30, 18) {real, imag} */,
  {32'hc55b9378, 32'h00000000} /* (13, 30, 17) {real, imag} */,
  {32'hc5846a8c, 32'h00000000} /* (13, 30, 16) {real, imag} */,
  {32'hc5a8c985, 32'h00000000} /* (13, 30, 15) {real, imag} */,
  {32'hc5a9db0e, 32'h00000000} /* (13, 30, 14) {real, imag} */,
  {32'hc5a1d365, 32'h00000000} /* (13, 30, 13) {real, imag} */,
  {32'hc5590109, 32'h00000000} /* (13, 30, 12) {real, imag} */,
  {32'hc50f402a, 32'h00000000} /* (13, 30, 11) {real, imag} */,
  {32'hc3315460, 32'h00000000} /* (13, 30, 10) {real, imag} */,
  {32'h453af010, 32'h00000000} /* (13, 30, 9) {real, imag} */,
  {32'h453f421e, 32'h00000000} /* (13, 30, 8) {real, imag} */,
  {32'h457bf12a, 32'h00000000} /* (13, 30, 7) {real, imag} */,
  {32'h45e058d6, 32'h00000000} /* (13, 30, 6) {real, imag} */,
  {32'h45d51538, 32'h00000000} /* (13, 30, 5) {real, imag} */,
  {32'h45f3468e, 32'h00000000} /* (13, 30, 4) {real, imag} */,
  {32'h45fb0faf, 32'h00000000} /* (13, 30, 3) {real, imag} */,
  {32'h45f6a982, 32'h00000000} /* (13, 30, 2) {real, imag} */,
  {32'h45fab324, 32'h00000000} /* (13, 30, 1) {real, imag} */,
  {32'h45ff6576, 32'h00000000} /* (13, 30, 0) {real, imag} */,
  {32'h46119cfc, 32'h00000000} /* (13, 29, 31) {real, imag} */,
  {32'h461c899e, 32'h00000000} /* (13, 29, 30) {real, imag} */,
  {32'h461f8848, 32'h00000000} /* (13, 29, 29) {real, imag} */,
  {32'h4608336a, 32'h00000000} /* (13, 29, 28) {real, imag} */,
  {32'h460eb11b, 32'h00000000} /* (13, 29, 27) {real, imag} */,
  {32'h461fd03e, 32'h00000000} /* (13, 29, 26) {real, imag} */,
  {32'h461b7c1e, 32'h00000000} /* (13, 29, 25) {real, imag} */,
  {32'h45fe86f8, 32'h00000000} /* (13, 29, 24) {real, imag} */,
  {32'h45fbd43a, 32'h00000000} /* (13, 29, 23) {real, imag} */,
  {32'h45d53556, 32'h00000000} /* (13, 29, 22) {real, imag} */,
  {32'h45597bb4, 32'h00000000} /* (13, 29, 21) {real, imag} */,
  {32'h42b1b240, 32'h00000000} /* (13, 29, 20) {real, imag} */,
  {32'hc50dd03c, 32'h00000000} /* (13, 29, 19) {real, imag} */,
  {32'hc5547c1e, 32'h00000000} /* (13, 29, 18) {real, imag} */,
  {32'hc5a6cf39, 32'h00000000} /* (13, 29, 17) {real, imag} */,
  {32'hc5af0a08, 32'h00000000} /* (13, 29, 16) {real, imag} */,
  {32'hc5c2b4c3, 32'h00000000} /* (13, 29, 15) {real, imag} */,
  {32'hc5abde1f, 32'h00000000} /* (13, 29, 14) {real, imag} */,
  {32'hc5931658, 32'h00000000} /* (13, 29, 13) {real, imag} */,
  {32'hc557f423, 32'h00000000} /* (13, 29, 12) {real, imag} */,
  {32'hc4d1da08, 32'h00000000} /* (13, 29, 11) {real, imag} */,
  {32'h446f2998, 32'h00000000} /* (13, 29, 10) {real, imag} */,
  {32'h457512e4, 32'h00000000} /* (13, 29, 9) {real, imag} */,
  {32'h458202b4, 32'h00000000} /* (13, 29, 8) {real, imag} */,
  {32'h45a6cc50, 32'h00000000} /* (13, 29, 7) {real, imag} */,
  {32'h45df0d62, 32'h00000000} /* (13, 29, 6) {real, imag} */,
  {32'h45f4a6e6, 32'h00000000} /* (13, 29, 5) {real, imag} */,
  {32'h46020108, 32'h00000000} /* (13, 29, 4) {real, imag} */,
  {32'h46003cca, 32'h00000000} /* (13, 29, 3) {real, imag} */,
  {32'h460f6ba2, 32'h00000000} /* (13, 29, 2) {real, imag} */,
  {32'h461b8f6e, 32'h00000000} /* (13, 29, 1) {real, imag} */,
  {32'h4600ce7d, 32'h00000000} /* (13, 29, 0) {real, imag} */,
  {32'h4608f380, 32'h00000000} /* (13, 28, 31) {real, imag} */,
  {32'h461b0062, 32'h00000000} /* (13, 28, 30) {real, imag} */,
  {32'h461a381d, 32'h00000000} /* (13, 28, 29) {real, imag} */,
  {32'h461b7ae8, 32'h00000000} /* (13, 28, 28) {real, imag} */,
  {32'h46202307, 32'h00000000} /* (13, 28, 27) {real, imag} */,
  {32'h4617b3b0, 32'h00000000} /* (13, 28, 26) {real, imag} */,
  {32'h460b35c1, 32'h00000000} /* (13, 28, 25) {real, imag} */,
  {32'h4606eba2, 32'h00000000} /* (13, 28, 24) {real, imag} */,
  {32'h45e76c36, 32'h00000000} /* (13, 28, 23) {real, imag} */,
  {32'h45a2abfa, 32'h00000000} /* (13, 28, 22) {real, imag} */,
  {32'h455c5f11, 32'h00000000} /* (13, 28, 21) {real, imag} */,
  {32'h4306a9f0, 32'h00000000} /* (13, 28, 20) {real, imag} */,
  {32'hc5218baa, 32'h00000000} /* (13, 28, 19) {real, imag} */,
  {32'hc58f24cb, 32'h00000000} /* (13, 28, 18) {real, imag} */,
  {32'hc5ab2990, 32'h00000000} /* (13, 28, 17) {real, imag} */,
  {32'hc5c8432a, 32'h00000000} /* (13, 28, 16) {real, imag} */,
  {32'hc5c1603c, 32'h00000000} /* (13, 28, 15) {real, imag} */,
  {32'hc5b6e152, 32'h00000000} /* (13, 28, 14) {real, imag} */,
  {32'hc5901ed6, 32'h00000000} /* (13, 28, 13) {real, imag} */,
  {32'hc561a664, 32'h00000000} /* (13, 28, 12) {real, imag} */,
  {32'hc4fd8d20, 32'h00000000} /* (13, 28, 11) {real, imag} */,
  {32'h4446e888, 32'h00000000} /* (13, 28, 10) {real, imag} */,
  {32'h454a13bc, 32'h00000000} /* (13, 28, 9) {real, imag} */,
  {32'h459dca92, 32'h00000000} /* (13, 28, 8) {real, imag} */,
  {32'h45cc005e, 32'h00000000} /* (13, 28, 7) {real, imag} */,
  {32'h45e43b46, 32'h00000000} /* (13, 28, 6) {real, imag} */,
  {32'h46142fd2, 32'h00000000} /* (13, 28, 5) {real, imag} */,
  {32'h45f69eec, 32'h00000000} /* (13, 28, 4) {real, imag} */,
  {32'h45ed4c39, 32'h00000000} /* (13, 28, 3) {real, imag} */,
  {32'h4609cd78, 32'h00000000} /* (13, 28, 2) {real, imag} */,
  {32'h4607ca17, 32'h00000000} /* (13, 28, 1) {real, imag} */,
  {32'h4607a95f, 32'h00000000} /* (13, 28, 0) {real, imag} */,
  {32'h4606b404, 32'h00000000} /* (13, 27, 31) {real, imag} */,
  {32'h46175ec6, 32'h00000000} /* (13, 27, 30) {real, imag} */,
  {32'h4621313e, 32'h00000000} /* (13, 27, 29) {real, imag} */,
  {32'h4629623c, 32'h00000000} /* (13, 27, 28) {real, imag} */,
  {32'h462a150c, 32'h00000000} /* (13, 27, 27) {real, imag} */,
  {32'h460ac4a8, 32'h00000000} /* (13, 27, 26) {real, imag} */,
  {32'h4610cd14, 32'h00000000} /* (13, 27, 25) {real, imag} */,
  {32'h460461fc, 32'h00000000} /* (13, 27, 24) {real, imag} */,
  {32'h45d5c614, 32'h00000000} /* (13, 27, 23) {real, imag} */,
  {32'h45c5db37, 32'h00000000} /* (13, 27, 22) {real, imag} */,
  {32'h453943ba, 32'h00000000} /* (13, 27, 21) {real, imag} */,
  {32'h428884c0, 32'h00000000} /* (13, 27, 20) {real, imag} */,
  {32'hc51190d6, 32'h00000000} /* (13, 27, 19) {real, imag} */,
  {32'hc598bde2, 32'h00000000} /* (13, 27, 18) {real, imag} */,
  {32'hc5bea64e, 32'h00000000} /* (13, 27, 17) {real, imag} */,
  {32'hc5baa474, 32'h00000000} /* (13, 27, 16) {real, imag} */,
  {32'hc5e96d50, 32'h00000000} /* (13, 27, 15) {real, imag} */,
  {32'hc5a98e3d, 32'h00000000} /* (13, 27, 14) {real, imag} */,
  {32'hc593b2eb, 32'h00000000} /* (13, 27, 13) {real, imag} */,
  {32'hc57549f8, 32'h00000000} /* (13, 27, 12) {real, imag} */,
  {32'hc50c454a, 32'h00000000} /* (13, 27, 11) {real, imag} */,
  {32'h44968302, 32'h00000000} /* (13, 27, 10) {real, imag} */,
  {32'h45809217, 32'h00000000} /* (13, 27, 9) {real, imag} */,
  {32'h45b22918, 32'h00000000} /* (13, 27, 8) {real, imag} */,
  {32'h45de970c, 32'h00000000} /* (13, 27, 7) {real, imag} */,
  {32'h45f55cdd, 32'h00000000} /* (13, 27, 6) {real, imag} */,
  {32'h45f4befd, 32'h00000000} /* (13, 27, 5) {real, imag} */,
  {32'h45f9bfcb, 32'h00000000} /* (13, 27, 4) {real, imag} */,
  {32'h460935ee, 32'h00000000} /* (13, 27, 3) {real, imag} */,
  {32'h45f5cf34, 32'h00000000} /* (13, 27, 2) {real, imag} */,
  {32'h4603dbea, 32'h00000000} /* (13, 27, 1) {real, imag} */,
  {32'h460c0d34, 32'h00000000} /* (13, 27, 0) {real, imag} */,
  {32'h46066207, 32'h00000000} /* (13, 26, 31) {real, imag} */,
  {32'h461470e4, 32'h00000000} /* (13, 26, 30) {real, imag} */,
  {32'h461d9048, 32'h00000000} /* (13, 26, 29) {real, imag} */,
  {32'h4618d9f2, 32'h00000000} /* (13, 26, 28) {real, imag} */,
  {32'h460c6816, 32'h00000000} /* (13, 26, 27) {real, imag} */,
  {32'h4620d043, 32'h00000000} /* (13, 26, 26) {real, imag} */,
  {32'h461ba937, 32'h00000000} /* (13, 26, 25) {real, imag} */,
  {32'h45dce2be, 32'h00000000} /* (13, 26, 24) {real, imag} */,
  {32'h45dad520, 32'h00000000} /* (13, 26, 23) {real, imag} */,
  {32'h45ae6344, 32'h00000000} /* (13, 26, 22) {real, imag} */,
  {32'h44e73ce4, 32'h00000000} /* (13, 26, 21) {real, imag} */,
  {32'hc4132e48, 32'h00000000} /* (13, 26, 20) {real, imag} */,
  {32'hc539caba, 32'h00000000} /* (13, 26, 19) {real, imag} */,
  {32'hc5ab7a16, 32'h00000000} /* (13, 26, 18) {real, imag} */,
  {32'hc5b5f7d6, 32'h00000000} /* (13, 26, 17) {real, imag} */,
  {32'hc5d9ce1d, 32'h00000000} /* (13, 26, 16) {real, imag} */,
  {32'hc5d77380, 32'h00000000} /* (13, 26, 15) {real, imag} */,
  {32'hc5a6472c, 32'h00000000} /* (13, 26, 14) {real, imag} */,
  {32'hc58ef6fb, 32'h00000000} /* (13, 26, 13) {real, imag} */,
  {32'hc592a800, 32'h00000000} /* (13, 26, 12) {real, imag} */,
  {32'hc4be9ecc, 32'h00000000} /* (13, 26, 11) {real, imag} */,
  {32'h447fdaf0, 32'h00000000} /* (13, 26, 10) {real, imag} */,
  {32'h45717a7b, 32'h00000000} /* (13, 26, 9) {real, imag} */,
  {32'h45c280c0, 32'h00000000} /* (13, 26, 8) {real, imag} */,
  {32'h45f4cc82, 32'h00000000} /* (13, 26, 7) {real, imag} */,
  {32'h45f3d2d0, 32'h00000000} /* (13, 26, 6) {real, imag} */,
  {32'h46045584, 32'h00000000} /* (13, 26, 5) {real, imag} */,
  {32'h45fd600b, 32'h00000000} /* (13, 26, 4) {real, imag} */,
  {32'h45f8d159, 32'h00000000} /* (13, 26, 3) {real, imag} */,
  {32'h4603cef1, 32'h00000000} /* (13, 26, 2) {real, imag} */,
  {32'h45f86592, 32'h00000000} /* (13, 26, 1) {real, imag} */,
  {32'h45ecb879, 32'h00000000} /* (13, 26, 0) {real, imag} */,
  {32'h45fb9bc1, 32'h00000000} /* (13, 25, 31) {real, imag} */,
  {32'h460531f8, 32'h00000000} /* (13, 25, 30) {real, imag} */,
  {32'h461897be, 32'h00000000} /* (13, 25, 29) {real, imag} */,
  {32'h46085cc5, 32'h00000000} /* (13, 25, 28) {real, imag} */,
  {32'h460b12f2, 32'h00000000} /* (13, 25, 27) {real, imag} */,
  {32'h4609d72a, 32'h00000000} /* (13, 25, 26) {real, imag} */,
  {32'h4610d523, 32'h00000000} /* (13, 25, 25) {real, imag} */,
  {32'h45f2e18e, 32'h00000000} /* (13, 25, 24) {real, imag} */,
  {32'h45c5fe96, 32'h00000000} /* (13, 25, 23) {real, imag} */,
  {32'h4591d3d1, 32'h00000000} /* (13, 25, 22) {real, imag} */,
  {32'h45290c70, 32'h00000000} /* (13, 25, 21) {real, imag} */,
  {32'hc495ceac, 32'h00000000} /* (13, 25, 20) {real, imag} */,
  {32'hc563275a, 32'h00000000} /* (13, 25, 19) {real, imag} */,
  {32'hc599d7a7, 32'h00000000} /* (13, 25, 18) {real, imag} */,
  {32'hc5b685ff, 32'h00000000} /* (13, 25, 17) {real, imag} */,
  {32'hc5d51dba, 32'h00000000} /* (13, 25, 16) {real, imag} */,
  {32'hc5c07ed5, 32'h00000000} /* (13, 25, 15) {real, imag} */,
  {32'hc5b71a54, 32'h00000000} /* (13, 25, 14) {real, imag} */,
  {32'hc5d0c520, 32'h00000000} /* (13, 25, 13) {real, imag} */,
  {32'hc581416a, 32'h00000000} /* (13, 25, 12) {real, imag} */,
  {32'hc5088df4, 32'h00000000} /* (13, 25, 11) {real, imag} */,
  {32'h4483f6b8, 32'h00000000} /* (13, 25, 10) {real, imag} */,
  {32'h45897fd0, 32'h00000000} /* (13, 25, 9) {real, imag} */,
  {32'h45cced72, 32'h00000000} /* (13, 25, 8) {real, imag} */,
  {32'h45c970d2, 32'h00000000} /* (13, 25, 7) {real, imag} */,
  {32'h45d7cf9f, 32'h00000000} /* (13, 25, 6) {real, imag} */,
  {32'h46031ab8, 32'h00000000} /* (13, 25, 5) {real, imag} */,
  {32'h45f4748f, 32'h00000000} /* (13, 25, 4) {real, imag} */,
  {32'h45f47e33, 32'h00000000} /* (13, 25, 3) {real, imag} */,
  {32'h45e7a199, 32'h00000000} /* (13, 25, 2) {real, imag} */,
  {32'h45f0e89f, 32'h00000000} /* (13, 25, 1) {real, imag} */,
  {32'h45eef876, 32'h00000000} /* (13, 25, 0) {real, imag} */,
  {32'h45d47808, 32'h00000000} /* (13, 24, 31) {real, imag} */,
  {32'h45db457c, 32'h00000000} /* (13, 24, 30) {real, imag} */,
  {32'h46004936, 32'h00000000} /* (13, 24, 29) {real, imag} */,
  {32'h45f7c7ec, 32'h00000000} /* (13, 24, 28) {real, imag} */,
  {32'h45e41d0e, 32'h00000000} /* (13, 24, 27) {real, imag} */,
  {32'h45ebe121, 32'h00000000} /* (13, 24, 26) {real, imag} */,
  {32'h45ed512e, 32'h00000000} /* (13, 24, 25) {real, imag} */,
  {32'h45ec1550, 32'h00000000} /* (13, 24, 24) {real, imag} */,
  {32'h459d5832, 32'h00000000} /* (13, 24, 23) {real, imag} */,
  {32'h458588b0, 32'h00000000} /* (13, 24, 22) {real, imag} */,
  {32'h451c9dc8, 32'h00000000} /* (13, 24, 21) {real, imag} */,
  {32'hc41ca1ec, 32'h00000000} /* (13, 24, 20) {real, imag} */,
  {32'hc53eb227, 32'h00000000} /* (13, 24, 19) {real, imag} */,
  {32'hc59c575b, 32'h00000000} /* (13, 24, 18) {real, imag} */,
  {32'hc5ba6694, 32'h00000000} /* (13, 24, 17) {real, imag} */,
  {32'hc5dd0227, 32'h00000000} /* (13, 24, 16) {real, imag} */,
  {32'hc5b812e8, 32'h00000000} /* (13, 24, 15) {real, imag} */,
  {32'hc5bb328c, 32'h00000000} /* (13, 24, 14) {real, imag} */,
  {32'hc5ebb057, 32'h00000000} /* (13, 24, 13) {real, imag} */,
  {32'hc5a5b2f0, 32'h00000000} /* (13, 24, 12) {real, imag} */,
  {32'hc5327617, 32'h00000000} /* (13, 24, 11) {real, imag} */,
  {32'h44717168, 32'h00000000} /* (13, 24, 10) {real, imag} */,
  {32'h4585eb34, 32'h00000000} /* (13, 24, 9) {real, imag} */,
  {32'h45abf83e, 32'h00000000} /* (13, 24, 8) {real, imag} */,
  {32'h45becd92, 32'h00000000} /* (13, 24, 7) {real, imag} */,
  {32'h45b6d754, 32'h00000000} /* (13, 24, 6) {real, imag} */,
  {32'h45cab154, 32'h00000000} /* (13, 24, 5) {real, imag} */,
  {32'h45e141ae, 32'h00000000} /* (13, 24, 4) {real, imag} */,
  {32'h45cf1128, 32'h00000000} /* (13, 24, 3) {real, imag} */,
  {32'h45c4329f, 32'h00000000} /* (13, 24, 2) {real, imag} */,
  {32'h45caf61a, 32'h00000000} /* (13, 24, 1) {real, imag} */,
  {32'h45d82679, 32'h00000000} /* (13, 24, 0) {real, imag} */,
  {32'h45aaab2c, 32'h00000000} /* (13, 23, 31) {real, imag} */,
  {32'h45d2577b, 32'h00000000} /* (13, 23, 30) {real, imag} */,
  {32'h45bbd9dc, 32'h00000000} /* (13, 23, 29) {real, imag} */,
  {32'h45c61c24, 32'h00000000} /* (13, 23, 28) {real, imag} */,
  {32'h45b0f7dc, 32'h00000000} /* (13, 23, 27) {real, imag} */,
  {32'h45b83427, 32'h00000000} /* (13, 23, 26) {real, imag} */,
  {32'h45aaa4f8, 32'h00000000} /* (13, 23, 25) {real, imag} */,
  {32'h45a68897, 32'h00000000} /* (13, 23, 24) {real, imag} */,
  {32'h45919492, 32'h00000000} /* (13, 23, 23) {real, imag} */,
  {32'h4550cf5c, 32'h00000000} /* (13, 23, 22) {real, imag} */,
  {32'h44cf5084, 32'h00000000} /* (13, 23, 21) {real, imag} */,
  {32'hc4e150aa, 32'h00000000} /* (13, 23, 20) {real, imag} */,
  {32'hc5207082, 32'h00000000} /* (13, 23, 19) {real, imag} */,
  {32'hc57215c5, 32'h00000000} /* (13, 23, 18) {real, imag} */,
  {32'hc58f2417, 32'h00000000} /* (13, 23, 17) {real, imag} */,
  {32'hc5a59d46, 32'h00000000} /* (13, 23, 16) {real, imag} */,
  {32'hc5ae344e, 32'h00000000} /* (13, 23, 15) {real, imag} */,
  {32'hc5a282d3, 32'h00000000} /* (13, 23, 14) {real, imag} */,
  {32'hc5a7afc8, 32'h00000000} /* (13, 23, 13) {real, imag} */,
  {32'hc5912d6a, 32'h00000000} /* (13, 23, 12) {real, imag} */,
  {32'hc527d358, 32'h00000000} /* (13, 23, 11) {real, imag} */,
  {32'h42c40900, 32'h00000000} /* (13, 23, 10) {real, imag} */,
  {32'h4517b6dd, 32'h00000000} /* (13, 23, 9) {real, imag} */,
  {32'h45a20759, 32'h00000000} /* (13, 23, 8) {real, imag} */,
  {32'h45a88206, 32'h00000000} /* (13, 23, 7) {real, imag} */,
  {32'h45aa2af8, 32'h00000000} /* (13, 23, 6) {real, imag} */,
  {32'h45b138de, 32'h00000000} /* (13, 23, 5) {real, imag} */,
  {32'h45b504d4, 32'h00000000} /* (13, 23, 4) {real, imag} */,
  {32'h45b16dfb, 32'h00000000} /* (13, 23, 3) {real, imag} */,
  {32'h45ac7e7e, 32'h00000000} /* (13, 23, 2) {real, imag} */,
  {32'h45ac735f, 32'h00000000} /* (13, 23, 1) {real, imag} */,
  {32'h45a6dfa2, 32'h00000000} /* (13, 23, 0) {real, imag} */,
  {32'h4589768e, 32'h00000000} /* (13, 22, 31) {real, imag} */,
  {32'h4599d120, 32'h00000000} /* (13, 22, 30) {real, imag} */,
  {32'h4596b4c0, 32'h00000000} /* (13, 22, 29) {real, imag} */,
  {32'h459b4772, 32'h00000000} /* (13, 22, 28) {real, imag} */,
  {32'h4567393d, 32'h00000000} /* (13, 22, 27) {real, imag} */,
  {32'h45754eed, 32'h00000000} /* (13, 22, 26) {real, imag} */,
  {32'h4550b9ee, 32'h00000000} /* (13, 22, 25) {real, imag} */,
  {32'h455915e1, 32'h00000000} /* (13, 22, 24) {real, imag} */,
  {32'h454d1cf6, 32'h00000000} /* (13, 22, 23) {real, imag} */,
  {32'h4527a481, 32'h00000000} /* (13, 22, 22) {real, imag} */,
  {32'h4421f3c8, 32'h00000000} /* (13, 22, 21) {real, imag} */,
  {32'hc4e8e4f6, 32'h00000000} /* (13, 22, 20) {real, imag} */,
  {32'hc50fd68e, 32'h00000000} /* (13, 22, 19) {real, imag} */,
  {32'hc5398712, 32'h00000000} /* (13, 22, 18) {real, imag} */,
  {32'hc5406d38, 32'h00000000} /* (13, 22, 17) {real, imag} */,
  {32'hc53185d0, 32'h00000000} /* (13, 22, 16) {real, imag} */,
  {32'hc5347ce3, 32'h00000000} /* (13, 22, 15) {real, imag} */,
  {32'hc53ac0bf, 32'h00000000} /* (13, 22, 14) {real, imag} */,
  {32'hc5525d83, 32'h00000000} /* (13, 22, 13) {real, imag} */,
  {32'hc5405ecc, 32'h00000000} /* (13, 22, 12) {real, imag} */,
  {32'hc5091eab, 32'h00000000} /* (13, 22, 11) {real, imag} */,
  {32'hc3c4aef8, 32'h00000000} /* (13, 22, 10) {real, imag} */,
  {32'h451e8888, 32'h00000000} /* (13, 22, 9) {real, imag} */,
  {32'h45385193, 32'h00000000} /* (13, 22, 8) {real, imag} */,
  {32'h458dff81, 32'h00000000} /* (13, 22, 7) {real, imag} */,
  {32'h457602a7, 32'h00000000} /* (13, 22, 6) {real, imag} */,
  {32'h45781c0e, 32'h00000000} /* (13, 22, 5) {real, imag} */,
  {32'h456fdd53, 32'h00000000} /* (13, 22, 4) {real, imag} */,
  {32'h45603504, 32'h00000000} /* (13, 22, 3) {real, imag} */,
  {32'h458b1c55, 32'h00000000} /* (13, 22, 2) {real, imag} */,
  {32'h4568a1f6, 32'h00000000} /* (13, 22, 1) {real, imag} */,
  {32'h454c3684, 32'h00000000} /* (13, 22, 0) {real, imag} */,
  {32'h4499f7e0, 32'h00000000} /* (13, 21, 31) {real, imag} */,
  {32'h44a8209d, 32'h00000000} /* (13, 21, 30) {real, imag} */,
  {32'h44d29e91, 32'h00000000} /* (13, 21, 29) {real, imag} */,
  {32'h447fd638, 32'h00000000} /* (13, 21, 28) {real, imag} */,
  {32'h4483469e, 32'h00000000} /* (13, 21, 27) {real, imag} */,
  {32'h441dc180, 32'h00000000} /* (13, 21, 26) {real, imag} */,
  {32'hc3267460, 32'h00000000} /* (13, 21, 25) {real, imag} */,
  {32'h44de94d3, 32'h00000000} /* (13, 21, 24) {real, imag} */,
  {32'h4475aa8d, 32'h00000000} /* (13, 21, 23) {real, imag} */,
  {32'h447b040a, 32'h00000000} /* (13, 21, 22) {real, imag} */,
  {32'h4355337c, 32'h00000000} /* (13, 21, 21) {real, imag} */,
  {32'h4417baf6, 32'h00000000} /* (13, 21, 20) {real, imag} */,
  {32'hc44a1674, 32'h00000000} /* (13, 21, 19) {real, imag} */,
  {32'hc465b52d, 32'h00000000} /* (13, 21, 18) {real, imag} */,
  {32'hc48914b7, 32'h00000000} /* (13, 21, 17) {real, imag} */,
  {32'hc3e6daa4, 32'h00000000} /* (13, 21, 16) {real, imag} */,
  {32'hc3cf057e, 32'h00000000} /* (13, 21, 15) {real, imag} */,
  {32'hc409b4c4, 32'h00000000} /* (13, 21, 14) {real, imag} */,
  {32'hc3a1c414, 32'h00000000} /* (13, 21, 13) {real, imag} */,
  {32'hc3ab5d07, 32'h00000000} /* (13, 21, 12) {real, imag} */,
  {32'hc483542a, 32'h00000000} /* (13, 21, 11) {real, imag} */,
  {32'hc39e995f, 32'h00000000} /* (13, 21, 10) {real, imag} */,
  {32'h44fca984, 32'h00000000} /* (13, 21, 9) {real, imag} */,
  {32'h4513dd28, 32'h00000000} /* (13, 21, 8) {real, imag} */,
  {32'h44f22a3a, 32'h00000000} /* (13, 21, 7) {real, imag} */,
  {32'h4303656e, 32'h00000000} /* (13, 21, 6) {real, imag} */,
  {32'h44b6a09a, 32'h00000000} /* (13, 21, 5) {real, imag} */,
  {32'h44c2475b, 32'h00000000} /* (13, 21, 4) {real, imag} */,
  {32'h44841913, 32'h00000000} /* (13, 21, 3) {real, imag} */,
  {32'h44ad7384, 32'h00000000} /* (13, 21, 2) {real, imag} */,
  {32'h4499f895, 32'h00000000} /* (13, 21, 1) {real, imag} */,
  {32'h44daaee5, 32'h00000000} /* (13, 21, 0) {real, imag} */,
  {32'hc4c41192, 32'h00000000} /* (13, 20, 31) {real, imag} */,
  {32'hc4f8fdb4, 32'h00000000} /* (13, 20, 30) {real, imag} */,
  {32'hc5088433, 32'h00000000} /* (13, 20, 29) {real, imag} */,
  {32'hc5427a32, 32'h00000000} /* (13, 20, 28) {real, imag} */,
  {32'hc53571d0, 32'h00000000} /* (13, 20, 27) {real, imag} */,
  {32'hc512b75c, 32'h00000000} /* (13, 20, 26) {real, imag} */,
  {32'hc511e03c, 32'h00000000} /* (13, 20, 25) {real, imag} */,
  {32'hc4bb454d, 32'h00000000} /* (13, 20, 24) {real, imag} */,
  {32'hc4c55019, 32'h00000000} /* (13, 20, 23) {real, imag} */,
  {32'hc4c2898d, 32'h00000000} /* (13, 20, 22) {real, imag} */,
  {32'hc4015302, 32'h00000000} /* (13, 20, 21) {real, imag} */,
  {32'h44595ee1, 32'h00000000} /* (13, 20, 20) {real, imag} */,
  {32'h44cfdc12, 32'h00000000} /* (13, 20, 19) {real, imag} */,
  {32'h451e4248, 32'h00000000} /* (13, 20, 18) {real, imag} */,
  {32'h451b3f25, 32'h00000000} /* (13, 20, 17) {real, imag} */,
  {32'h45057da3, 32'h00000000} /* (13, 20, 16) {real, imag} */,
  {32'h4502218a, 32'h00000000} /* (13, 20, 15) {real, imag} */,
  {32'h45298938, 32'h00000000} /* (13, 20, 14) {real, imag} */,
  {32'h44df1966, 32'h00000000} /* (13, 20, 13) {real, imag} */,
  {32'h44eadca0, 32'h00000000} /* (13, 20, 12) {real, imag} */,
  {32'h44880073, 32'h00000000} /* (13, 20, 11) {real, imag} */,
  {32'hc4766dc3, 32'h00000000} /* (13, 20, 10) {real, imag} */,
  {32'hc391dbec, 32'h00000000} /* (13, 20, 9) {real, imag} */,
  {32'hc49030c3, 32'h00000000} /* (13, 20, 8) {real, imag} */,
  {32'hc4e02217, 32'h00000000} /* (13, 20, 7) {real, imag} */,
  {32'hc516f9c5, 32'h00000000} /* (13, 20, 6) {real, imag} */,
  {32'hc513d9cc, 32'h00000000} /* (13, 20, 5) {real, imag} */,
  {32'hc51cce9e, 32'h00000000} /* (13, 20, 4) {real, imag} */,
  {32'hc5018a0b, 32'h00000000} /* (13, 20, 3) {real, imag} */,
  {32'hc545bef4, 32'h00000000} /* (13, 20, 2) {real, imag} */,
  {32'hc507ac67, 32'h00000000} /* (13, 20, 1) {real, imag} */,
  {32'hc4da6c8c, 32'h00000000} /* (13, 20, 0) {real, imag} */,
  {32'hc5527718, 32'h00000000} /* (13, 19, 31) {real, imag} */,
  {32'hc57337f6, 32'h00000000} /* (13, 19, 30) {real, imag} */,
  {32'hc5a53449, 32'h00000000} /* (13, 19, 29) {real, imag} */,
  {32'hc596cb66, 32'h00000000} /* (13, 19, 28) {real, imag} */,
  {32'hc5a03ce4, 32'h00000000} /* (13, 19, 27) {real, imag} */,
  {32'hc57a0311, 32'h00000000} /* (13, 19, 26) {real, imag} */,
  {32'hc56b31a2, 32'h00000000} /* (13, 19, 25) {real, imag} */,
  {32'hc5687667, 32'h00000000} /* (13, 19, 24) {real, imag} */,
  {32'hc56f737a, 32'h00000000} /* (13, 19, 23) {real, imag} */,
  {32'hc525909c, 32'h00000000} /* (13, 19, 22) {real, imag} */,
  {32'hc4917eed, 32'h00000000} /* (13, 19, 21) {real, imag} */,
  {32'h44aaf581, 32'h00000000} /* (13, 19, 20) {real, imag} */,
  {32'h455bd612, 32'h00000000} /* (13, 19, 19) {real, imag} */,
  {32'h4582dd77, 32'h00000000} /* (13, 19, 18) {real, imag} */,
  {32'h456a321a, 32'h00000000} /* (13, 19, 17) {real, imag} */,
  {32'h4580c01b, 32'h00000000} /* (13, 19, 16) {real, imag} */,
  {32'h458ff503, 32'h00000000} /* (13, 19, 15) {real, imag} */,
  {32'h457e6eb2, 32'h00000000} /* (13, 19, 14) {real, imag} */,
  {32'h452969a2, 32'h00000000} /* (13, 19, 13) {real, imag} */,
  {32'h454e2e52, 32'h00000000} /* (13, 19, 12) {real, imag} */,
  {32'h44eaba1e, 32'h00000000} /* (13, 19, 11) {real, imag} */,
  {32'hc4406cac, 32'h00000000} /* (13, 19, 10) {real, imag} */,
  {32'hc4ea795c, 32'h00000000} /* (13, 19, 9) {real, imag} */,
  {32'hc52bb465, 32'h00000000} /* (13, 19, 8) {real, imag} */,
  {32'hc58f9131, 32'h00000000} /* (13, 19, 7) {real, imag} */,
  {32'hc56d6784, 32'h00000000} /* (13, 19, 6) {real, imag} */,
  {32'hc5848bbb, 32'h00000000} /* (13, 19, 5) {real, imag} */,
  {32'hc570b652, 32'h00000000} /* (13, 19, 4) {real, imag} */,
  {32'hc589a73f, 32'h00000000} /* (13, 19, 3) {real, imag} */,
  {32'hc58f2c99, 32'h00000000} /* (13, 19, 2) {real, imag} */,
  {32'hc57239aa, 32'h00000000} /* (13, 19, 1) {real, imag} */,
  {32'hc55672aa, 32'h00000000} /* (13, 19, 0) {real, imag} */,
  {32'hc58d636c, 32'h00000000} /* (13, 18, 31) {real, imag} */,
  {32'hc5b81eb7, 32'h00000000} /* (13, 18, 30) {real, imag} */,
  {32'hc5b1203e, 32'h00000000} /* (13, 18, 29) {real, imag} */,
  {32'hc5b5ba4e, 32'h00000000} /* (13, 18, 28) {real, imag} */,
  {32'hc5b69964, 32'h00000000} /* (13, 18, 27) {real, imag} */,
  {32'hc5b3883a, 32'h00000000} /* (13, 18, 26) {real, imag} */,
  {32'hc5a0e74b, 32'h00000000} /* (13, 18, 25) {real, imag} */,
  {32'hc5b29f8d, 32'h00000000} /* (13, 18, 24) {real, imag} */,
  {32'hc5a564b4, 32'h00000000} /* (13, 18, 23) {real, imag} */,
  {32'hc5525beb, 32'h00000000} /* (13, 18, 22) {real, imag} */,
  {32'hc4c1ee54, 32'h00000000} /* (13, 18, 21) {real, imag} */,
  {32'h44ae9eaa, 32'h00000000} /* (13, 18, 20) {real, imag} */,
  {32'h4571da73, 32'h00000000} /* (13, 18, 19) {real, imag} */,
  {32'h4573ba43, 32'h00000000} /* (13, 18, 18) {real, imag} */,
  {32'h458e1c0e, 32'h00000000} /* (13, 18, 17) {real, imag} */,
  {32'h45a43f88, 32'h00000000} /* (13, 18, 16) {real, imag} */,
  {32'h45926922, 32'h00000000} /* (13, 18, 15) {real, imag} */,
  {32'h459b66cf, 32'h00000000} /* (13, 18, 14) {real, imag} */,
  {32'h458faf88, 32'h00000000} /* (13, 18, 13) {real, imag} */,
  {32'h45487c77, 32'h00000000} /* (13, 18, 12) {real, imag} */,
  {32'h4524bfe9, 32'h00000000} /* (13, 18, 11) {real, imag} */,
  {32'hc43c6ca4, 32'h00000000} /* (13, 18, 10) {real, imag} */,
  {32'hc5176400, 32'h00000000} /* (13, 18, 9) {real, imag} */,
  {32'hc58701b9, 32'h00000000} /* (13, 18, 8) {real, imag} */,
  {32'hc58e7b0c, 32'h00000000} /* (13, 18, 7) {real, imag} */,
  {32'hc5b2c8f4, 32'h00000000} /* (13, 18, 6) {real, imag} */,
  {32'hc5cbf85e, 32'h00000000} /* (13, 18, 5) {real, imag} */,
  {32'hc5c00b96, 32'h00000000} /* (13, 18, 4) {real, imag} */,
  {32'hc5b4b8a3, 32'h00000000} /* (13, 18, 3) {real, imag} */,
  {32'hc5b3f110, 32'h00000000} /* (13, 18, 2) {real, imag} */,
  {32'hc59f99ac, 32'h00000000} /* (13, 18, 1) {real, imag} */,
  {32'hc59536fc, 32'h00000000} /* (13, 18, 0) {real, imag} */,
  {32'hc5ae6095, 32'h00000000} /* (13, 17, 31) {real, imag} */,
  {32'hc5c6baa6, 32'h00000000} /* (13, 17, 30) {real, imag} */,
  {32'hc5f8037b, 32'h00000000} /* (13, 17, 29) {real, imag} */,
  {32'hc5cba277, 32'h00000000} /* (13, 17, 28) {real, imag} */,
  {32'hc5ddd382, 32'h00000000} /* (13, 17, 27) {real, imag} */,
  {32'hc5d81bb6, 32'h00000000} /* (13, 17, 26) {real, imag} */,
  {32'hc5b585e4, 32'h00000000} /* (13, 17, 25) {real, imag} */,
  {32'hc5d3fba0, 32'h00000000} /* (13, 17, 24) {real, imag} */,
  {32'hc5bc2082, 32'h00000000} /* (13, 17, 23) {real, imag} */,
  {32'hc59dee01, 32'h00000000} /* (13, 17, 22) {real, imag} */,
  {32'hc432e088, 32'h00000000} /* (13, 17, 21) {real, imag} */,
  {32'h44bbc9b0, 32'h00000000} /* (13, 17, 20) {real, imag} */,
  {32'h4571f250, 32'h00000000} /* (13, 17, 19) {real, imag} */,
  {32'h45898134, 32'h00000000} /* (13, 17, 18) {real, imag} */,
  {32'h45a6c68b, 32'h00000000} /* (13, 17, 17) {real, imag} */,
  {32'h45b367fa, 32'h00000000} /* (13, 17, 16) {real, imag} */,
  {32'h45b6578d, 32'h00000000} /* (13, 17, 15) {real, imag} */,
  {32'h45a0dae6, 32'h00000000} /* (13, 17, 14) {real, imag} */,
  {32'h45855335, 32'h00000000} /* (13, 17, 13) {real, imag} */,
  {32'h457b2182, 32'h00000000} /* (13, 17, 12) {real, imag} */,
  {32'h450a10f4, 32'h00000000} /* (13, 17, 11) {real, imag} */,
  {32'hc404d790, 32'h00000000} /* (13, 17, 10) {real, imag} */,
  {32'hc540bf05, 32'h00000000} /* (13, 17, 9) {real, imag} */,
  {32'hc59cfdb0, 32'h00000000} /* (13, 17, 8) {real, imag} */,
  {32'hc5acdd34, 32'h00000000} /* (13, 17, 7) {real, imag} */,
  {32'hc5ebad0b, 32'h00000000} /* (13, 17, 6) {real, imag} */,
  {32'hc5d539f9, 32'h00000000} /* (13, 17, 5) {real, imag} */,
  {32'hc5e81efa, 32'h00000000} /* (13, 17, 4) {real, imag} */,
  {32'hc5da57f2, 32'h00000000} /* (13, 17, 3) {real, imag} */,
  {32'hc5b82340, 32'h00000000} /* (13, 17, 2) {real, imag} */,
  {32'hc5cd8875, 32'h00000000} /* (13, 17, 1) {real, imag} */,
  {32'hc5af52b6, 32'h00000000} /* (13, 17, 0) {real, imag} */,
  {32'hc5c33f59, 32'h00000000} /* (13, 16, 31) {real, imag} */,
  {32'hc5d48c0c, 32'h00000000} /* (13, 16, 30) {real, imag} */,
  {32'hc5e6f25e, 32'h00000000} /* (13, 16, 29) {real, imag} */,
  {32'hc5eb3718, 32'h00000000} /* (13, 16, 28) {real, imag} */,
  {32'hc5f66959, 32'h00000000} /* (13, 16, 27) {real, imag} */,
  {32'hc5e76c3a, 32'h00000000} /* (13, 16, 26) {real, imag} */,
  {32'hc5db8e8f, 32'h00000000} /* (13, 16, 25) {real, imag} */,
  {32'hc5d3a122, 32'h00000000} /* (13, 16, 24) {real, imag} */,
  {32'hc5b1c260, 32'h00000000} /* (13, 16, 23) {real, imag} */,
  {32'hc59d8a2f, 32'h00000000} /* (13, 16, 22) {real, imag} */,
  {32'hc4502418, 32'h00000000} /* (13, 16, 21) {real, imag} */,
  {32'h452a2a6a, 32'h00000000} /* (13, 16, 20) {real, imag} */,
  {32'h4569ae84, 32'h00000000} /* (13, 16, 19) {real, imag} */,
  {32'h45a0a490, 32'h00000000} /* (13, 16, 18) {real, imag} */,
  {32'h45d60fa4, 32'h00000000} /* (13, 16, 17) {real, imag} */,
  {32'h45ce160a, 32'h00000000} /* (13, 16, 16) {real, imag} */,
  {32'h45d83c7f, 32'h00000000} /* (13, 16, 15) {real, imag} */,
  {32'h45a84cac, 32'h00000000} /* (13, 16, 14) {real, imag} */,
  {32'h459623c4, 32'h00000000} /* (13, 16, 13) {real, imag} */,
  {32'h45a11eb0, 32'h00000000} /* (13, 16, 12) {real, imag} */,
  {32'h4521c796, 32'h00000000} /* (13, 16, 11) {real, imag} */,
  {32'h43463b20, 32'h00000000} /* (13, 16, 10) {real, imag} */,
  {32'hc534f612, 32'h00000000} /* (13, 16, 9) {real, imag} */,
  {32'hc58107f0, 32'h00000000} /* (13, 16, 8) {real, imag} */,
  {32'hc5ae0fde, 32'h00000000} /* (13, 16, 7) {real, imag} */,
  {32'hc5cce33b, 32'h00000000} /* (13, 16, 6) {real, imag} */,
  {32'hc5e444bc, 32'h00000000} /* (13, 16, 5) {real, imag} */,
  {32'hc5d2eeed, 32'h00000000} /* (13, 16, 4) {real, imag} */,
  {32'hc5d88e58, 32'h00000000} /* (13, 16, 3) {real, imag} */,
  {32'hc5d34714, 32'h00000000} /* (13, 16, 2) {real, imag} */,
  {32'hc5dd9116, 32'h00000000} /* (13, 16, 1) {real, imag} */,
  {32'hc5c59ad8, 32'h00000000} /* (13, 16, 0) {real, imag} */,
  {32'hc5dca29e, 32'h00000000} /* (13, 15, 31) {real, imag} */,
  {32'hc5dabc4c, 32'h00000000} /* (13, 15, 30) {real, imag} */,
  {32'hc600cb21, 32'h00000000} /* (13, 15, 29) {real, imag} */,
  {32'hc6032aaf, 32'h00000000} /* (13, 15, 28) {real, imag} */,
  {32'hc5f25549, 32'h00000000} /* (13, 15, 27) {real, imag} */,
  {32'hc5df274a, 32'h00000000} /* (13, 15, 26) {real, imag} */,
  {32'hc5ce67bd, 32'h00000000} /* (13, 15, 25) {real, imag} */,
  {32'hc5a86202, 32'h00000000} /* (13, 15, 24) {real, imag} */,
  {32'hc5b2d5c9, 32'h00000000} /* (13, 15, 23) {real, imag} */,
  {32'hc56e506e, 32'h00000000} /* (13, 15, 22) {real, imag} */,
  {32'hc4c03d68, 32'h00000000} /* (13, 15, 21) {real, imag} */,
  {32'h450e97cf, 32'h00000000} /* (13, 15, 20) {real, imag} */,
  {32'h4584084b, 32'h00000000} /* (13, 15, 19) {real, imag} */,
  {32'h45ac2d92, 32'h00000000} /* (13, 15, 18) {real, imag} */,
  {32'h45d35a49, 32'h00000000} /* (13, 15, 17) {real, imag} */,
  {32'h45c5abdc, 32'h00000000} /* (13, 15, 16) {real, imag} */,
  {32'h45c987fc, 32'h00000000} /* (13, 15, 15) {real, imag} */,
  {32'h45b3094a, 32'h00000000} /* (13, 15, 14) {real, imag} */,
  {32'h45a0aa02, 32'h00000000} /* (13, 15, 13) {real, imag} */,
  {32'h458fde04, 32'h00000000} /* (13, 15, 12) {real, imag} */,
  {32'h453d4e2e, 32'h00000000} /* (13, 15, 11) {real, imag} */,
  {32'h4329d150, 32'h00000000} /* (13, 15, 10) {real, imag} */,
  {32'hc53417d2, 32'h00000000} /* (13, 15, 9) {real, imag} */,
  {32'hc58c67b6, 32'h00000000} /* (13, 15, 8) {real, imag} */,
  {32'hc5c29a7b, 32'h00000000} /* (13, 15, 7) {real, imag} */,
  {32'hc5dd51c9, 32'h00000000} /* (13, 15, 6) {real, imag} */,
  {32'hc5c4e186, 32'h00000000} /* (13, 15, 5) {real, imag} */,
  {32'hc5d82afe, 32'h00000000} /* (13, 15, 4) {real, imag} */,
  {32'hc5d07c23, 32'h00000000} /* (13, 15, 3) {real, imag} */,
  {32'hc5e1592e, 32'h00000000} /* (13, 15, 2) {real, imag} */,
  {32'hc602d522, 32'h00000000} /* (13, 15, 1) {real, imag} */,
  {32'hc5e6e0c4, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'hc5b92eab, 32'h00000000} /* (13, 14, 31) {real, imag} */,
  {32'hc5c6c863, 32'h00000000} /* (13, 14, 30) {real, imag} */,
  {32'hc5e1ef16, 32'h00000000} /* (13, 14, 29) {real, imag} */,
  {32'hc5eec738, 32'h00000000} /* (13, 14, 28) {real, imag} */,
  {32'hc5d59f12, 32'h00000000} /* (13, 14, 27) {real, imag} */,
  {32'hc5bb78ff, 32'h00000000} /* (13, 14, 26) {real, imag} */,
  {32'hc5aa2553, 32'h00000000} /* (13, 14, 25) {real, imag} */,
  {32'hc5967316, 32'h00000000} /* (13, 14, 24) {real, imag} */,
  {32'hc5977adc, 32'h00000000} /* (13, 14, 23) {real, imag} */,
  {32'hc51d9195, 32'h00000000} /* (13, 14, 22) {real, imag} */,
  {32'h44009d94, 32'h00000000} /* (13, 14, 21) {real, imag} */,
  {32'h44e73a1a, 32'h00000000} /* (13, 14, 20) {real, imag} */,
  {32'h4586a40a, 32'h00000000} /* (13, 14, 19) {real, imag} */,
  {32'h459d861a, 32'h00000000} /* (13, 14, 18) {real, imag} */,
  {32'h45a6e936, 32'h00000000} /* (13, 14, 17) {real, imag} */,
  {32'h45d27f62, 32'h00000000} /* (13, 14, 16) {real, imag} */,
  {32'h45bc4b65, 32'h00000000} /* (13, 14, 15) {real, imag} */,
  {32'h45a62905, 32'h00000000} /* (13, 14, 14) {real, imag} */,
  {32'h459ab132, 32'h00000000} /* (13, 14, 13) {real, imag} */,
  {32'h455c6c01, 32'h00000000} /* (13, 14, 12) {real, imag} */,
  {32'h4509f6c4, 32'h00000000} /* (13, 14, 11) {real, imag} */,
  {32'hc412ea40, 32'h00000000} /* (13, 14, 10) {real, imag} */,
  {32'hc5185930, 32'h00000000} /* (13, 14, 9) {real, imag} */,
  {32'hc57ba8e7, 32'h00000000} /* (13, 14, 8) {real, imag} */,
  {32'hc5af038a, 32'h00000000} /* (13, 14, 7) {real, imag} */,
  {32'hc5ccc354, 32'h00000000} /* (13, 14, 6) {real, imag} */,
  {32'hc5c10902, 32'h00000000} /* (13, 14, 5) {real, imag} */,
  {32'hc5d17c1a, 32'h00000000} /* (13, 14, 4) {real, imag} */,
  {32'hc5d3365e, 32'h00000000} /* (13, 14, 3) {real, imag} */,
  {32'hc5e0300a, 32'h00000000} /* (13, 14, 2) {real, imag} */,
  {32'hc5f1db28, 32'h00000000} /* (13, 14, 1) {real, imag} */,
  {32'hc5ef45da, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'hc5a07434, 32'h00000000} /* (13, 13, 31) {real, imag} */,
  {32'hc5bb1d4d, 32'h00000000} /* (13, 13, 30) {real, imag} */,
  {32'hc5c08dd5, 32'h00000000} /* (13, 13, 29) {real, imag} */,
  {32'hc5b9ae06, 32'h00000000} /* (13, 13, 28) {real, imag} */,
  {32'hc5c1ec7d, 32'h00000000} /* (13, 13, 27) {real, imag} */,
  {32'hc595b8e6, 32'h00000000} /* (13, 13, 26) {real, imag} */,
  {32'hc589b9bf, 32'h00000000} /* (13, 13, 25) {real, imag} */,
  {32'hc5939f46, 32'h00000000} /* (13, 13, 24) {real, imag} */,
  {32'hc5443a41, 32'h00000000} /* (13, 13, 23) {real, imag} */,
  {32'hc4d69de2, 32'h00000000} /* (13, 13, 22) {real, imag} */,
  {32'hc2e94700, 32'h00000000} /* (13, 13, 21) {real, imag} */,
  {32'h44e8c973, 32'h00000000} /* (13, 13, 20) {real, imag} */,
  {32'h457b3786, 32'h00000000} /* (13, 13, 19) {real, imag} */,
  {32'h4596aa02, 32'h00000000} /* (13, 13, 18) {real, imag} */,
  {32'h45a780ba, 32'h00000000} /* (13, 13, 17) {real, imag} */,
  {32'h459942b7, 32'h00000000} /* (13, 13, 16) {real, imag} */,
  {32'h45b4b20c, 32'h00000000} /* (13, 13, 15) {real, imag} */,
  {32'h45a92fb5, 32'h00000000} /* (13, 13, 14) {real, imag} */,
  {32'h457a1aca, 32'h00000000} /* (13, 13, 13) {real, imag} */,
  {32'h45478f30, 32'h00000000} /* (13, 13, 12) {real, imag} */,
  {32'h450c9a1a, 32'h00000000} /* (13, 13, 11) {real, imag} */,
  {32'hc384a360, 32'h00000000} /* (13, 13, 10) {real, imag} */,
  {32'hc5119b74, 32'h00000000} /* (13, 13, 9) {real, imag} */,
  {32'hc5618ad4, 32'h00000000} /* (13, 13, 8) {real, imag} */,
  {32'hc5b5e848, 32'h00000000} /* (13, 13, 7) {real, imag} */,
  {32'hc5aa9946, 32'h00000000} /* (13, 13, 6) {real, imag} */,
  {32'hc5a5ad6a, 32'h00000000} /* (13, 13, 5) {real, imag} */,
  {32'hc5afc80b, 32'h00000000} /* (13, 13, 4) {real, imag} */,
  {32'hc5abdc69, 32'h00000000} /* (13, 13, 3) {real, imag} */,
  {32'hc5ad883a, 32'h00000000} /* (13, 13, 2) {real, imag} */,
  {32'hc5b389de, 32'h00000000} /* (13, 13, 1) {real, imag} */,
  {32'hc5ae9419, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'hc569f598, 32'h00000000} /* (13, 12, 31) {real, imag} */,
  {32'hc58f5948, 32'h00000000} /* (13, 12, 30) {real, imag} */,
  {32'hc5b4f62b, 32'h00000000} /* (13, 12, 29) {real, imag} */,
  {32'hc5a28b0b, 32'h00000000} /* (13, 12, 28) {real, imag} */,
  {32'hc55b924f, 32'h00000000} /* (13, 12, 27) {real, imag} */,
  {32'hc53f416c, 32'h00000000} /* (13, 12, 26) {real, imag} */,
  {32'hc552f8ba, 32'h00000000} /* (13, 12, 25) {real, imag} */,
  {32'hc5318c00, 32'h00000000} /* (13, 12, 24) {real, imag} */,
  {32'hc5133233, 32'h00000000} /* (13, 12, 23) {real, imag} */,
  {32'hc4b0e158, 32'h00000000} /* (13, 12, 22) {real, imag} */,
  {32'h43b84240, 32'h00000000} /* (13, 12, 21) {real, imag} */,
  {32'h45315860, 32'h00000000} /* (13, 12, 20) {real, imag} */,
  {32'h45ab42f3, 32'h00000000} /* (13, 12, 19) {real, imag} */,
  {32'h4586d409, 32'h00000000} /* (13, 12, 18) {real, imag} */,
  {32'h458198ae, 32'h00000000} /* (13, 12, 17) {real, imag} */,
  {32'h458db2e3, 32'h00000000} /* (13, 12, 16) {real, imag} */,
  {32'h4593dba8, 32'h00000000} /* (13, 12, 15) {real, imag} */,
  {32'h4559a190, 32'h00000000} /* (13, 12, 14) {real, imag} */,
  {32'h452d639e, 32'h00000000} /* (13, 12, 13) {real, imag} */,
  {32'h455c8896, 32'h00000000} /* (13, 12, 12) {real, imag} */,
  {32'h4535d64d, 32'h00000000} /* (13, 12, 11) {real, imag} */,
  {32'hc3a34cec, 32'h00000000} /* (13, 12, 10) {real, imag} */,
  {32'hc50457ca, 32'h00000000} /* (13, 12, 9) {real, imag} */,
  {32'hc5365928, 32'h00000000} /* (13, 12, 8) {real, imag} */,
  {32'hc5884832, 32'h00000000} /* (13, 12, 7) {real, imag} */,
  {32'hc575739c, 32'h00000000} /* (13, 12, 6) {real, imag} */,
  {32'hc5901468, 32'h00000000} /* (13, 12, 5) {real, imag} */,
  {32'hc55cea5e, 32'h00000000} /* (13, 12, 4) {real, imag} */,
  {32'hc58221ef, 32'h00000000} /* (13, 12, 3) {real, imag} */,
  {32'hc5870ae1, 32'h00000000} /* (13, 12, 2) {real, imag} */,
  {32'hc56bc302, 32'h00000000} /* (13, 12, 1) {real, imag} */,
  {32'hc559ccaa, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'hc4b79dc2, 32'h00000000} /* (13, 11, 31) {real, imag} */,
  {32'hc4e812dc, 32'h00000000} /* (13, 11, 30) {real, imag} */,
  {32'hc4bed3d4, 32'h00000000} /* (13, 11, 29) {real, imag} */,
  {32'hc52a61c8, 32'h00000000} /* (13, 11, 28) {real, imag} */,
  {32'hc49d30c4, 32'h00000000} /* (13, 11, 27) {real, imag} */,
  {32'hc4af3f94, 32'h00000000} /* (13, 11, 26) {real, imag} */,
  {32'hc433a1aa, 32'h00000000} /* (13, 11, 25) {real, imag} */,
  {32'hc47e093e, 32'h00000000} /* (13, 11, 24) {real, imag} */,
  {32'hc45067dd, 32'h00000000} /* (13, 11, 23) {real, imag} */,
  {32'h44022f60, 32'h00000000} /* (13, 11, 22) {real, imag} */,
  {32'h44727cf0, 32'h00000000} /* (13, 11, 21) {real, imag} */,
  {32'h44f84aea, 32'h00000000} /* (13, 11, 20) {real, imag} */,
  {32'h451a70f0, 32'h00000000} /* (13, 11, 19) {real, imag} */,
  {32'h454abb55, 32'h00000000} /* (13, 11, 18) {real, imag} */,
  {32'h457d6f54, 32'h00000000} /* (13, 11, 17) {real, imag} */,
  {32'h45530fdd, 32'h00000000} /* (13, 11, 16) {real, imag} */,
  {32'h4505a4cf, 32'h00000000} /* (13, 11, 15) {real, imag} */,
  {32'h44fa7970, 32'h00000000} /* (13, 11, 14) {real, imag} */,
  {32'h45115393, 32'h00000000} /* (13, 11, 13) {real, imag} */,
  {32'h45104a8a, 32'h00000000} /* (13, 11, 12) {real, imag} */,
  {32'h44f998d4, 32'h00000000} /* (13, 11, 11) {real, imag} */,
  {32'hc41f5fd1, 32'h00000000} /* (13, 11, 10) {real, imag} */,
  {32'hc4e78261, 32'h00000000} /* (13, 11, 9) {real, imag} */,
  {32'hc4e3e325, 32'h00000000} /* (13, 11, 8) {real, imag} */,
  {32'hc50c2ea7, 32'h00000000} /* (13, 11, 7) {real, imag} */,
  {32'hc5742618, 32'h00000000} /* (13, 11, 6) {real, imag} */,
  {32'hc4f20e08, 32'h00000000} /* (13, 11, 5) {real, imag} */,
  {32'hc4d2e73e, 32'h00000000} /* (13, 11, 4) {real, imag} */,
  {32'hc5124556, 32'h00000000} /* (13, 11, 3) {real, imag} */,
  {32'hc4cb0022, 32'h00000000} /* (13, 11, 2) {real, imag} */,
  {32'hc4c337f5, 32'h00000000} /* (13, 11, 1) {real, imag} */,
  {32'hc4cf4db6, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'h4529cecb, 32'h00000000} /* (13, 10, 31) {real, imag} */,
  {32'h452cbc1e, 32'h00000000} /* (13, 10, 30) {real, imag} */,
  {32'h450a9c16, 32'h00000000} /* (13, 10, 29) {real, imag} */,
  {32'h4555d839, 32'h00000000} /* (13, 10, 28) {real, imag} */,
  {32'h44eaf214, 32'h00000000} /* (13, 10, 27) {real, imag} */,
  {32'h44f155a6, 32'h00000000} /* (13, 10, 26) {real, imag} */,
  {32'h44e33434, 32'h00000000} /* (13, 10, 25) {real, imag} */,
  {32'h450d6044, 32'h00000000} /* (13, 10, 24) {real, imag} */,
  {32'h44c0a4e6, 32'h00000000} /* (13, 10, 23) {real, imag} */,
  {32'h44fbaea2, 32'h00000000} /* (13, 10, 22) {real, imag} */,
  {32'h4437e8bc, 32'h00000000} /* (13, 10, 21) {real, imag} */,
  {32'h440f9f36, 32'h00000000} /* (13, 10, 20) {real, imag} */,
  {32'h43e7da8c, 32'h00000000} /* (13, 10, 19) {real, imag} */,
  {32'h431859c8, 32'h00000000} /* (13, 10, 18) {real, imag} */,
  {32'h44f0bc65, 32'h00000000} /* (13, 10, 17) {real, imag} */,
  {32'h421bd240, 32'h00000000} /* (13, 10, 16) {real, imag} */,
  {32'hc3a15fd0, 32'h00000000} /* (13, 10, 15) {real, imag} */,
  {32'h42d77850, 32'h00000000} /* (13, 10, 14) {real, imag} */,
  {32'h43fd98ac, 32'h00000000} /* (13, 10, 13) {real, imag} */,
  {32'hc446df64, 32'h00000000} /* (13, 10, 12) {real, imag} */,
  {32'hc492c0f8, 32'h00000000} /* (13, 10, 11) {real, imag} */,
  {32'hc3166350, 32'h00000000} /* (13, 10, 10) {real, imag} */,
  {32'hc152e440, 32'h00000000} /* (13, 10, 9) {real, imag} */,
  {32'hc2558720, 32'h00000000} /* (13, 10, 8) {real, imag} */,
  {32'h441fcbf9, 32'h00000000} /* (13, 10, 7) {real, imag} */,
  {32'h441208a4, 32'h00000000} /* (13, 10, 6) {real, imag} */,
  {32'h4452b630, 32'h00000000} /* (13, 10, 5) {real, imag} */,
  {32'h448ef124, 32'h00000000} /* (13, 10, 4) {real, imag} */,
  {32'h44dafe75, 32'h00000000} /* (13, 10, 3) {real, imag} */,
  {32'h44bf5597, 32'h00000000} /* (13, 10, 2) {real, imag} */,
  {32'h44bc16ab, 32'h00000000} /* (13, 10, 1) {real, imag} */,
  {32'h449887bf, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h455178d8, 32'h00000000} /* (13, 9, 31) {real, imag} */,
  {32'h456e049b, 32'h00000000} /* (13, 9, 30) {real, imag} */,
  {32'h4583b7fb, 32'h00000000} /* (13, 9, 29) {real, imag} */,
  {32'h45a2fd79, 32'h00000000} /* (13, 9, 28) {real, imag} */,
  {32'h45a6b74c, 32'h00000000} /* (13, 9, 27) {real, imag} */,
  {32'h4593471f, 32'h00000000} /* (13, 9, 26) {real, imag} */,
  {32'h4597c5b2, 32'h00000000} /* (13, 9, 25) {real, imag} */,
  {32'h45add2f5, 32'h00000000} /* (13, 9, 24) {real, imag} */,
  {32'h45691cf4, 32'h00000000} /* (13, 9, 23) {real, imag} */,
  {32'h45576300, 32'h00000000} /* (13, 9, 22) {real, imag} */,
  {32'h4520c4f9, 32'h00000000} /* (13, 9, 21) {real, imag} */,
  {32'h43a45870, 32'h00000000} /* (13, 9, 20) {real, imag} */,
  {32'h43c10bb8, 32'h00000000} /* (13, 9, 19) {real, imag} */,
  {32'hc4acbcce, 32'h00000000} /* (13, 9, 18) {real, imag} */,
  {32'hc4dbc59e, 32'h00000000} /* (13, 9, 17) {real, imag} */,
  {32'hc52ba9a6, 32'h00000000} /* (13, 9, 16) {real, imag} */,
  {32'hc4d50b9c, 32'h00000000} /* (13, 9, 15) {real, imag} */,
  {32'hc569bebf, 32'h00000000} /* (13, 9, 14) {real, imag} */,
  {32'hc50a3522, 32'h00000000} /* (13, 9, 13) {real, imag} */,
  {32'hc5034524, 32'h00000000} /* (13, 9, 12) {real, imag} */,
  {32'hc4ee6021, 32'h00000000} /* (13, 9, 11) {real, imag} */,
  {32'h4441cfa0, 32'h00000000} /* (13, 9, 10) {real, imag} */,
  {32'h448db45e, 32'h00000000} /* (13, 9, 9) {real, imag} */,
  {32'h44f68025, 32'h00000000} /* (13, 9, 8) {real, imag} */,
  {32'h4541a96e, 32'h00000000} /* (13, 9, 7) {real, imag} */,
  {32'h451accf6, 32'h00000000} /* (13, 9, 6) {real, imag} */,
  {32'h4588e001, 32'h00000000} /* (13, 9, 5) {real, imag} */,
  {32'h45792d4c, 32'h00000000} /* (13, 9, 4) {real, imag} */,
  {32'h456d7eab, 32'h00000000} /* (13, 9, 3) {real, imag} */,
  {32'h4572e49f, 32'h00000000} /* (13, 9, 2) {real, imag} */,
  {32'h4571ffbd, 32'h00000000} /* (13, 9, 1) {real, imag} */,
  {32'h456fe7f4, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'h45a2001d, 32'h00000000} /* (13, 8, 31) {real, imag} */,
  {32'h45ac8934, 32'h00000000} /* (13, 8, 30) {real, imag} */,
  {32'h459ea2a6, 32'h00000000} /* (13, 8, 29) {real, imag} */,
  {32'h45bdcacf, 32'h00000000} /* (13, 8, 28) {real, imag} */,
  {32'h45d45988, 32'h00000000} /* (13, 8, 27) {real, imag} */,
  {32'h45c46156, 32'h00000000} /* (13, 8, 26) {real, imag} */,
  {32'h45bf622c, 32'h00000000} /* (13, 8, 25) {real, imag} */,
  {32'h45cb1952, 32'h00000000} /* (13, 8, 24) {real, imag} */,
  {32'h45a9ecfd, 32'h00000000} /* (13, 8, 23) {real, imag} */,
  {32'h458468da, 32'h00000000} /* (13, 8, 22) {real, imag} */,
  {32'h4548304e, 32'h00000000} /* (13, 8, 21) {real, imag} */,
  {32'h448b995b, 32'h00000000} /* (13, 8, 20) {real, imag} */,
  {32'hc4883d6a, 32'h00000000} /* (13, 8, 19) {real, imag} */,
  {32'hc48f7ba0, 32'h00000000} /* (13, 8, 18) {real, imag} */,
  {32'hc4ed25ae, 32'h00000000} /* (13, 8, 17) {real, imag} */,
  {32'hc541d778, 32'h00000000} /* (13, 8, 16) {real, imag} */,
  {32'hc57299ba, 32'h00000000} /* (13, 8, 15) {real, imag} */,
  {32'hc57ab673, 32'h00000000} /* (13, 8, 14) {real, imag} */,
  {32'hc54e0304, 32'h00000000} /* (13, 8, 13) {real, imag} */,
  {32'hc5339a42, 32'h00000000} /* (13, 8, 12) {real, imag} */,
  {32'hc521adff, 32'h00000000} /* (13, 8, 11) {real, imag} */,
  {32'hc3ab5d70, 32'h00000000} /* (13, 8, 10) {real, imag} */,
  {32'h44f83248, 32'h00000000} /* (13, 8, 9) {real, imag} */,
  {32'h45337c48, 32'h00000000} /* (13, 8, 8) {real, imag} */,
  {32'h457d307e, 32'h00000000} /* (13, 8, 7) {real, imag} */,
  {32'h45866f62, 32'h00000000} /* (13, 8, 6) {real, imag} */,
  {32'h459e55e3, 32'h00000000} /* (13, 8, 5) {real, imag} */,
  {32'h45a1994f, 32'h00000000} /* (13, 8, 4) {real, imag} */,
  {32'h45a9d09a, 32'h00000000} /* (13, 8, 3) {real, imag} */,
  {32'h45c68121, 32'h00000000} /* (13, 8, 2) {real, imag} */,
  {32'h45a3a1ac, 32'h00000000} /* (13, 8, 1) {real, imag} */,
  {32'h4597bd52, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'h45b953ba, 32'h00000000} /* (13, 7, 31) {real, imag} */,
  {32'h45cbac04, 32'h00000000} /* (13, 7, 30) {real, imag} */,
  {32'h45cbaed6, 32'h00000000} /* (13, 7, 29) {real, imag} */,
  {32'h45ddf4d0, 32'h00000000} /* (13, 7, 28) {real, imag} */,
  {32'h45e8c39e, 32'h00000000} /* (13, 7, 27) {real, imag} */,
  {32'h45f10bd8, 32'h00000000} /* (13, 7, 26) {real, imag} */,
  {32'h45d30301, 32'h00000000} /* (13, 7, 25) {real, imag} */,
  {32'h45f3b48c, 32'h00000000} /* (13, 7, 24) {real, imag} */,
  {32'h45e404b6, 32'h00000000} /* (13, 7, 23) {real, imag} */,
  {32'h45da5f0d, 32'h00000000} /* (13, 7, 22) {real, imag} */,
  {32'h456e4245, 32'h00000000} /* (13, 7, 21) {real, imag} */,
  {32'h42fb4a60, 32'h00000000} /* (13, 7, 20) {real, imag} */,
  {32'hc41123a4, 32'h00000000} /* (13, 7, 19) {real, imag} */,
  {32'hc492d4d6, 32'h00000000} /* (13, 7, 18) {real, imag} */,
  {32'hc52751ee, 32'h00000000} /* (13, 7, 17) {real, imag} */,
  {32'hc5315e5a, 32'h00000000} /* (13, 7, 16) {real, imag} */,
  {32'hc57133a7, 32'h00000000} /* (13, 7, 15) {real, imag} */,
  {32'hc589550c, 32'h00000000} /* (13, 7, 14) {real, imag} */,
  {32'hc56e412b, 32'h00000000} /* (13, 7, 13) {real, imag} */,
  {32'hc5809c2a, 32'h00000000} /* (13, 7, 12) {real, imag} */,
  {32'hc57869f3, 32'h00000000} /* (13, 7, 11) {real, imag} */,
  {32'hc458c994, 32'h00000000} /* (13, 7, 10) {real, imag} */,
  {32'h449655ec, 32'h00000000} /* (13, 7, 9) {real, imag} */,
  {32'h45089737, 32'h00000000} /* (13, 7, 8) {real, imag} */,
  {32'h45a1b1d2, 32'h00000000} /* (13, 7, 7) {real, imag} */,
  {32'h4598a757, 32'h00000000} /* (13, 7, 6) {real, imag} */,
  {32'h45a55426, 32'h00000000} /* (13, 7, 5) {real, imag} */,
  {32'h45cbc87e, 32'h00000000} /* (13, 7, 4) {real, imag} */,
  {32'h45cebc9e, 32'h00000000} /* (13, 7, 3) {real, imag} */,
  {32'h45d56012, 32'h00000000} /* (13, 7, 2) {real, imag} */,
  {32'h45d08c2d, 32'h00000000} /* (13, 7, 1) {real, imag} */,
  {32'h45b230a3, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'h45d9073e, 32'h00000000} /* (13, 6, 31) {real, imag} */,
  {32'h45dcda84, 32'h00000000} /* (13, 6, 30) {real, imag} */,
  {32'h45ecb61a, 32'h00000000} /* (13, 6, 29) {real, imag} */,
  {32'h4608c172, 32'h00000000} /* (13, 6, 28) {real, imag} */,
  {32'h460c78ec, 32'h00000000} /* (13, 6, 27) {real, imag} */,
  {32'h45f9168f, 32'h00000000} /* (13, 6, 26) {real, imag} */,
  {32'h460abb6a, 32'h00000000} /* (13, 6, 25) {real, imag} */,
  {32'h45fe4d76, 32'h00000000} /* (13, 6, 24) {real, imag} */,
  {32'h45efe1d6, 32'h00000000} /* (13, 6, 23) {real, imag} */,
  {32'h45f136c5, 32'h00000000} /* (13, 6, 22) {real, imag} */,
  {32'h45b53ce0, 32'h00000000} /* (13, 6, 21) {real, imag} */,
  {32'h451a7d37, 32'h00000000} /* (13, 6, 20) {real, imag} */,
  {32'h44299f84, 32'h00000000} /* (13, 6, 19) {real, imag} */,
  {32'hc451ee88, 32'h00000000} /* (13, 6, 18) {real, imag} */,
  {32'hc4eabfbe, 32'h00000000} /* (13, 6, 17) {real, imag} */,
  {32'hc5221488, 32'h00000000} /* (13, 6, 16) {real, imag} */,
  {32'hc55605f8, 32'h00000000} /* (13, 6, 15) {real, imag} */,
  {32'hc57325c3, 32'h00000000} /* (13, 6, 14) {real, imag} */,
  {32'hc5992e0a, 32'h00000000} /* (13, 6, 13) {real, imag} */,
  {32'hc58f5e4f, 32'h00000000} /* (13, 6, 12) {real, imag} */,
  {32'hc55fbfda, 32'h00000000} /* (13, 6, 11) {real, imag} */,
  {32'hc4d26d64, 32'h00000000} /* (13, 6, 10) {real, imag} */,
  {32'h42163880, 32'h00000000} /* (13, 6, 9) {real, imag} */,
  {32'h44ced9f0, 32'h00000000} /* (13, 6, 8) {real, imag} */,
  {32'h454f60cd, 32'h00000000} /* (13, 6, 7) {real, imag} */,
  {32'h45944de7, 32'h00000000} /* (13, 6, 6) {real, imag} */,
  {32'h459b46d4, 32'h00000000} /* (13, 6, 5) {real, imag} */,
  {32'h45d4cc4a, 32'h00000000} /* (13, 6, 4) {real, imag} */,
  {32'h45cd6cdc, 32'h00000000} /* (13, 6, 3) {real, imag} */,
  {32'h45dbbed9, 32'h00000000} /* (13, 6, 2) {real, imag} */,
  {32'h45d9d41a, 32'h00000000} /* (13, 6, 1) {real, imag} */,
  {32'h45d2c902, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'h45f621fb, 32'h00000000} /* (13, 5, 31) {real, imag} */,
  {32'h4606873d, 32'h00000000} /* (13, 5, 30) {real, imag} */,
  {32'h460febfc, 32'h00000000} /* (13, 5, 29) {real, imag} */,
  {32'h460cb144, 32'h00000000} /* (13, 5, 28) {real, imag} */,
  {32'h461e2a26, 32'h00000000} /* (13, 5, 27) {real, imag} */,
  {32'h46120a26, 32'h00000000} /* (13, 5, 26) {real, imag} */,
  {32'h460c34bd, 32'h00000000} /* (13, 5, 25) {real, imag} */,
  {32'h4604014e, 32'h00000000} /* (13, 5, 24) {real, imag} */,
  {32'h45fabc86, 32'h00000000} /* (13, 5, 23) {real, imag} */,
  {32'h45f3b723, 32'h00000000} /* (13, 5, 22) {real, imag} */,
  {32'h45e87020, 32'h00000000} /* (13, 5, 21) {real, imag} */,
  {32'h4592ffa3, 32'h00000000} /* (13, 5, 20) {real, imag} */,
  {32'h45380c77, 32'h00000000} /* (13, 5, 19) {real, imag} */,
  {32'h44a19f68, 32'h00000000} /* (13, 5, 18) {real, imag} */,
  {32'h44c0f04a, 32'h00000000} /* (13, 5, 17) {real, imag} */,
  {32'hc47b183c, 32'h00000000} /* (13, 5, 16) {real, imag} */,
  {32'hc5437ada, 32'h00000000} /* (13, 5, 15) {real, imag} */,
  {32'hc594a771, 32'h00000000} /* (13, 5, 14) {real, imag} */,
  {32'hc58c50ed, 32'h00000000} /* (13, 5, 13) {real, imag} */,
  {32'hc5966c36, 32'h00000000} /* (13, 5, 12) {real, imag} */,
  {32'hc586641d, 32'h00000000} /* (13, 5, 11) {real, imag} */,
  {32'hc545aeae, 32'h00000000} /* (13, 5, 10) {real, imag} */,
  {32'hc4f87da2, 32'h00000000} /* (13, 5, 9) {real, imag} */,
  {32'hc482f3ce, 32'h00000000} /* (13, 5, 8) {real, imag} */,
  {32'h42a2a880, 32'h00000000} /* (13, 5, 7) {real, imag} */,
  {32'h45242636, 32'h00000000} /* (13, 5, 6) {real, imag} */,
  {32'h45a37b96, 32'h00000000} /* (13, 5, 5) {real, imag} */,
  {32'h45c241b1, 32'h00000000} /* (13, 5, 4) {real, imag} */,
  {32'h45e61448, 32'h00000000} /* (13, 5, 3) {real, imag} */,
  {32'h45e9dcf6, 32'h00000000} /* (13, 5, 2) {real, imag} */,
  {32'h45f58aac, 32'h00000000} /* (13, 5, 1) {real, imag} */,
  {32'h45e8eaa4, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h46053978, 32'h00000000} /* (13, 4, 31) {real, imag} */,
  {32'h460e1b86, 32'h00000000} /* (13, 4, 30) {real, imag} */,
  {32'h461c159a, 32'h00000000} /* (13, 4, 29) {real, imag} */,
  {32'h4617961a, 32'h00000000} /* (13, 4, 28) {real, imag} */,
  {32'h4619dd32, 32'h00000000} /* (13, 4, 27) {real, imag} */,
  {32'h461777a8, 32'h00000000} /* (13, 4, 26) {real, imag} */,
  {32'h46166272, 32'h00000000} /* (13, 4, 25) {real, imag} */,
  {32'h4613c392, 32'h00000000} /* (13, 4, 24) {real, imag} */,
  {32'h461be70c, 32'h00000000} /* (13, 4, 23) {real, imag} */,
  {32'h4618ac5a, 32'h00000000} /* (13, 4, 22) {real, imag} */,
  {32'h460e9fea, 32'h00000000} /* (13, 4, 21) {real, imag} */,
  {32'h45d833d8, 32'h00000000} /* (13, 4, 20) {real, imag} */,
  {32'h4592893a, 32'h00000000} /* (13, 4, 19) {real, imag} */,
  {32'h45773021, 32'h00000000} /* (13, 4, 18) {real, imag} */,
  {32'h451b958a, 32'h00000000} /* (13, 4, 17) {real, imag} */,
  {32'h447a7a4c, 32'h00000000} /* (13, 4, 16) {real, imag} */,
  {32'hc52625b2, 32'h00000000} /* (13, 4, 15) {real, imag} */,
  {32'hc591f352, 32'h00000000} /* (13, 4, 14) {real, imag} */,
  {32'hc58f5843, 32'h00000000} /* (13, 4, 13) {real, imag} */,
  {32'hc5a6b2b4, 32'h00000000} /* (13, 4, 12) {real, imag} */,
  {32'hc58873f9, 32'h00000000} /* (13, 4, 11) {real, imag} */,
  {32'hc59b9cad, 32'h00000000} /* (13, 4, 10) {real, imag} */,
  {32'hc575810c, 32'h00000000} /* (13, 4, 9) {real, imag} */,
  {32'hc52361b2, 32'h00000000} /* (13, 4, 8) {real, imag} */,
  {32'hc47bacb8, 32'h00000000} /* (13, 4, 7) {real, imag} */,
  {32'h44879140, 32'h00000000} /* (13, 4, 6) {real, imag} */,
  {32'h458a44b7, 32'h00000000} /* (13, 4, 5) {real, imag} */,
  {32'h45c08330, 32'h00000000} /* (13, 4, 4) {real, imag} */,
  {32'h45e988f2, 32'h00000000} /* (13, 4, 3) {real, imag} */,
  {32'h46021f4a, 32'h00000000} /* (13, 4, 2) {real, imag} */,
  {32'h45fe8a33, 32'h00000000} /* (13, 4, 1) {real, imag} */,
  {32'h45f90dc6, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'h4606ec77, 32'h00000000} /* (13, 3, 31) {real, imag} */,
  {32'h460fc454, 32'h00000000} /* (13, 3, 30) {real, imag} */,
  {32'h4610ae85, 32'h00000000} /* (13, 3, 29) {real, imag} */,
  {32'h46270376, 32'h00000000} /* (13, 3, 28) {real, imag} */,
  {32'h4628ba69, 32'h00000000} /* (13, 3, 27) {real, imag} */,
  {32'h462255c6, 32'h00000000} /* (13, 3, 26) {real, imag} */,
  {32'h461f3f03, 32'h00000000} /* (13, 3, 25) {real, imag} */,
  {32'h4632ca74, 32'h00000000} /* (13, 3, 24) {real, imag} */,
  {32'h46183756, 32'h00000000} /* (13, 3, 23) {real, imag} */,
  {32'h461007c7, 32'h00000000} /* (13, 3, 22) {real, imag} */,
  {32'h46046240, 32'h00000000} /* (13, 3, 21) {real, imag} */,
  {32'h45ca9c05, 32'h00000000} /* (13, 3, 20) {real, imag} */,
  {32'h45982cf4, 32'h00000000} /* (13, 3, 19) {real, imag} */,
  {32'h457277c8, 32'h00000000} /* (13, 3, 18) {real, imag} */,
  {32'h452fa2ae, 32'h00000000} /* (13, 3, 17) {real, imag} */,
  {32'hc2b0c4c0, 32'h00000000} /* (13, 3, 16) {real, imag} */,
  {32'hc508a179, 32'h00000000} /* (13, 3, 15) {real, imag} */,
  {32'hc5817a8d, 32'h00000000} /* (13, 3, 14) {real, imag} */,
  {32'hc5aa6746, 32'h00000000} /* (13, 3, 13) {real, imag} */,
  {32'hc5a34972, 32'h00000000} /* (13, 3, 12) {real, imag} */,
  {32'hc5d7a702, 32'h00000000} /* (13, 3, 11) {real, imag} */,
  {32'hc58f33a1, 32'h00000000} /* (13, 3, 10) {real, imag} */,
  {32'hc5942dee, 32'h00000000} /* (13, 3, 9) {real, imag} */,
  {32'hc5267544, 32'h00000000} /* (13, 3, 8) {real, imag} */,
  {32'hc4480c48, 32'h00000000} /* (13, 3, 7) {real, imag} */,
  {32'h4489b4d8, 32'h00000000} /* (13, 3, 6) {real, imag} */,
  {32'h4569bea0, 32'h00000000} /* (13, 3, 5) {real, imag} */,
  {32'h45dd084f, 32'h00000000} /* (13, 3, 4) {real, imag} */,
  {32'h45e9d28c, 32'h00000000} /* (13, 3, 3) {real, imag} */,
  {32'h45ecd3c6, 32'h00000000} /* (13, 3, 2) {real, imag} */,
  {32'h45fbc001, 32'h00000000} /* (13, 3, 1) {real, imag} */,
  {32'h4607baa8, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h4604c31b, 32'h00000000} /* (13, 2, 31) {real, imag} */,
  {32'h46122838, 32'h00000000} /* (13, 2, 30) {real, imag} */,
  {32'h462d27b2, 32'h00000000} /* (13, 2, 29) {real, imag} */,
  {32'h462b2e99, 32'h00000000} /* (13, 2, 28) {real, imag} */,
  {32'h462b6299, 32'h00000000} /* (13, 2, 27) {real, imag} */,
  {32'h4635c7fc, 32'h00000000} /* (13, 2, 26) {real, imag} */,
  {32'h4620243d, 32'h00000000} /* (13, 2, 25) {real, imag} */,
  {32'h4632a95e, 32'h00000000} /* (13, 2, 24) {real, imag} */,
  {32'h46109f45, 32'h00000000} /* (13, 2, 23) {real, imag} */,
  {32'h4601e75a, 32'h00000000} /* (13, 2, 22) {real, imag} */,
  {32'h45f000e7, 32'h00000000} /* (13, 2, 21) {real, imag} */,
  {32'h45be1ea9, 32'h00000000} /* (13, 2, 20) {real, imag} */,
  {32'h45aa7c1b, 32'h00000000} /* (13, 2, 19) {real, imag} */,
  {32'h456081f1, 32'h00000000} /* (13, 2, 18) {real, imag} */,
  {32'h44e9ffac, 32'h00000000} /* (13, 2, 17) {real, imag} */,
  {32'h444d73d0, 32'h00000000} /* (13, 2, 16) {real, imag} */,
  {32'hc507305b, 32'h00000000} /* (13, 2, 15) {real, imag} */,
  {32'hc59f02d0, 32'h00000000} /* (13, 2, 14) {real, imag} */,
  {32'hc5909b03, 32'h00000000} /* (13, 2, 13) {real, imag} */,
  {32'hc59eb01a, 32'h00000000} /* (13, 2, 12) {real, imag} */,
  {32'hc59fc996, 32'h00000000} /* (13, 2, 11) {real, imag} */,
  {32'hc592e069, 32'h00000000} /* (13, 2, 10) {real, imag} */,
  {32'hc57941e7, 32'h00000000} /* (13, 2, 9) {real, imag} */,
  {32'hc53bfc3e, 32'h00000000} /* (13, 2, 8) {real, imag} */,
  {32'hc4c61216, 32'h00000000} /* (13, 2, 7) {real, imag} */,
  {32'h4466ce24, 32'h00000000} /* (13, 2, 6) {real, imag} */,
  {32'h459394c3, 32'h00000000} /* (13, 2, 5) {real, imag} */,
  {32'h45d3d317, 32'h00000000} /* (13, 2, 4) {real, imag} */,
  {32'h45d33fc1, 32'h00000000} /* (13, 2, 3) {real, imag} */,
  {32'h4608a155, 32'h00000000} /* (13, 2, 2) {real, imag} */,
  {32'h460072ce, 32'h00000000} /* (13, 2, 1) {real, imag} */,
  {32'h460137b5, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h460246ea, 32'h00000000} /* (13, 1, 31) {real, imag} */,
  {32'h460da136, 32'h00000000} /* (13, 1, 30) {real, imag} */,
  {32'h46202c4f, 32'h00000000} /* (13, 1, 29) {real, imag} */,
  {32'h461efc9e, 32'h00000000} /* (13, 1, 28) {real, imag} */,
  {32'h46255cde, 32'h00000000} /* (13, 1, 27) {real, imag} */,
  {32'h4620f187, 32'h00000000} /* (13, 1, 26) {real, imag} */,
  {32'h46179c38, 32'h00000000} /* (13, 1, 25) {real, imag} */,
  {32'h460e8704, 32'h00000000} /* (13, 1, 24) {real, imag} */,
  {32'h4615906f, 32'h00000000} /* (13, 1, 23) {real, imag} */,
  {32'h45f014c2, 32'h00000000} /* (13, 1, 22) {real, imag} */,
  {32'h45d0e3aa, 32'h00000000} /* (13, 1, 21) {real, imag} */,
  {32'h45c6b68c, 32'h00000000} /* (13, 1, 20) {real, imag} */,
  {32'h4593d555, 32'h00000000} /* (13, 1, 19) {real, imag} */,
  {32'h452642be, 32'h00000000} /* (13, 1, 18) {real, imag} */,
  {32'h44de3d9c, 32'h00000000} /* (13, 1, 17) {real, imag} */,
  {32'h441910e0, 32'h00000000} /* (13, 1, 16) {real, imag} */,
  {32'hc51c6c51, 32'h00000000} /* (13, 1, 15) {real, imag} */,
  {32'hc57421e0, 32'h00000000} /* (13, 1, 14) {real, imag} */,
  {32'hc5a27a66, 32'h00000000} /* (13, 1, 13) {real, imag} */,
  {32'hc5a3382d, 32'h00000000} /* (13, 1, 12) {real, imag} */,
  {32'hc587909d, 32'h00000000} /* (13, 1, 11) {real, imag} */,
  {32'hc5861d7c, 32'h00000000} /* (13, 1, 10) {real, imag} */,
  {32'hc551505a, 32'h00000000} /* (13, 1, 9) {real, imag} */,
  {32'hc501c0ff, 32'h00000000} /* (13, 1, 8) {real, imag} */,
  {32'hc4b3f80a, 32'h00000000} /* (13, 1, 7) {real, imag} */,
  {32'hc36bb600, 32'h00000000} /* (13, 1, 6) {real, imag} */,
  {32'h4598dfe6, 32'h00000000} /* (13, 1, 5) {real, imag} */,
  {32'h45b2d840, 32'h00000000} /* (13, 1, 4) {real, imag} */,
  {32'h45d15e61, 32'h00000000} /* (13, 1, 3) {real, imag} */,
  {32'h45ff1b37, 32'h00000000} /* (13, 1, 2) {real, imag} */,
  {32'h4605f1de, 32'h00000000} /* (13, 1, 1) {real, imag} */,
  {32'h45ffe828, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h45ff2fbd, 32'h00000000} /* (13, 0, 31) {real, imag} */,
  {32'h4605be78, 32'h00000000} /* (13, 0, 30) {real, imag} */,
  {32'h460c2169, 32'h00000000} /* (13, 0, 29) {real, imag} */,
  {32'h461831cc, 32'h00000000} /* (13, 0, 28) {real, imag} */,
  {32'h461ef84f, 32'h00000000} /* (13, 0, 27) {real, imag} */,
  {32'h461bfc4b, 32'h00000000} /* (13, 0, 26) {real, imag} */,
  {32'h460d6f62, 32'h00000000} /* (13, 0, 25) {real, imag} */,
  {32'h460b44d8, 32'h00000000} /* (13, 0, 24) {real, imag} */,
  {32'h46000346, 32'h00000000} /* (13, 0, 23) {real, imag} */,
  {32'h45d6019c, 32'h00000000} /* (13, 0, 22) {real, imag} */,
  {32'h45b8a117, 32'h00000000} /* (13, 0, 21) {real, imag} */,
  {32'h45a48b27, 32'h00000000} /* (13, 0, 20) {real, imag} */,
  {32'h45510002, 32'h00000000} /* (13, 0, 19) {real, imag} */,
  {32'h44fe4680, 32'h00000000} /* (13, 0, 18) {real, imag} */,
  {32'h4499d73c, 32'h00000000} /* (13, 0, 17) {real, imag} */,
  {32'hc4ef500c, 32'h00000000} /* (13, 0, 16) {real, imag} */,
  {32'hc548bfee, 32'h00000000} /* (13, 0, 15) {real, imag} */,
  {32'hc56d7f13, 32'h00000000} /* (13, 0, 14) {real, imag} */,
  {32'hc588a08e, 32'h00000000} /* (13, 0, 13) {real, imag} */,
  {32'hc58114c0, 32'h00000000} /* (13, 0, 12) {real, imag} */,
  {32'hc56997ab, 32'h00000000} /* (13, 0, 11) {real, imag} */,
  {32'hc55e6374, 32'h00000000} /* (13, 0, 10) {real, imag} */,
  {32'hc4cd1794, 32'h00000000} /* (13, 0, 9) {real, imag} */,
  {32'hc3aa9690, 32'h00000000} /* (13, 0, 8) {real, imag} */,
  {32'h4404d6bc, 32'h00000000} /* (13, 0, 7) {real, imag} */,
  {32'h44d17d50, 32'h00000000} /* (13, 0, 6) {real, imag} */,
  {32'h457a8dc2, 32'h00000000} /* (13, 0, 5) {real, imag} */,
  {32'h45b1c995, 32'h00000000} /* (13, 0, 4) {real, imag} */,
  {32'h45e161ff, 32'h00000000} /* (13, 0, 3) {real, imag} */,
  {32'h45ddf54e, 32'h00000000} /* (13, 0, 2) {real, imag} */,
  {32'h45f9d6f1, 32'h00000000} /* (13, 0, 1) {real, imag} */,
  {32'h4608acf4, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h4628b9fa, 32'h00000000} /* (12, 31, 31) {real, imag} */,
  {32'h462e0a93, 32'h00000000} /* (12, 31, 30) {real, imag} */,
  {32'h46339af6, 32'h00000000} /* (12, 31, 29) {real, imag} */,
  {32'h46385f4a, 32'h00000000} /* (12, 31, 28) {real, imag} */,
  {32'h46395667, 32'h00000000} /* (12, 31, 27) {real, imag} */,
  {32'h46429c84, 32'h00000000} /* (12, 31, 26) {real, imag} */,
  {32'h462f04e0, 32'h00000000} /* (12, 31, 25) {real, imag} */,
  {32'h46229552, 32'h00000000} /* (12, 31, 24) {real, imag} */,
  {32'h4610b313, 32'h00000000} /* (12, 31, 23) {real, imag} */,
  {32'h45f9f654, 32'h00000000} /* (12, 31, 22) {real, imag} */,
  {32'h45a7d5a6, 32'h00000000} /* (12, 31, 21) {real, imag} */,
  {32'h453c2d92, 32'h00000000} /* (12, 31, 20) {real, imag} */,
  {32'h4442b3c8, 32'h00000000} /* (12, 31, 19) {real, imag} */,
  {32'hc3f695a0, 32'h00000000} /* (12, 31, 18) {real, imag} */,
  {32'hc4e0c37a, 32'h00000000} /* (12, 31, 17) {real, imag} */,
  {32'hc54e7ecc, 32'h00000000} /* (12, 31, 16) {real, imag} */,
  {32'hc589ea08, 32'h00000000} /* (12, 31, 15) {real, imag} */,
  {32'hc5aba896, 32'h00000000} /* (12, 31, 14) {real, imag} */,
  {32'hc5af28ed, 32'h00000000} /* (12, 31, 13) {real, imag} */,
  {32'hc58ccc6a, 32'h00000000} /* (12, 31, 12) {real, imag} */,
  {32'hc54ca408, 32'h00000000} /* (12, 31, 11) {real, imag} */,
  {32'hc4625b88, 32'h00000000} /* (12, 31, 10) {real, imag} */,
  {32'h446b0508, 32'h00000000} /* (12, 31, 9) {real, imag} */,
  {32'h44e8bb44, 32'h00000000} /* (12, 31, 8) {real, imag} */,
  {32'h4564791c, 32'h00000000} /* (12, 31, 7) {real, imag} */,
  {32'h45b75c74, 32'h00000000} /* (12, 31, 6) {real, imag} */,
  {32'h45da71c0, 32'h00000000} /* (12, 31, 5) {real, imag} */,
  {32'h4603f654, 32'h00000000} /* (12, 31, 4) {real, imag} */,
  {32'h460f2b46, 32'h00000000} /* (12, 31, 3) {real, imag} */,
  {32'h4623e05a, 32'h00000000} /* (12, 31, 2) {real, imag} */,
  {32'h461a0475, 32'h00000000} /* (12, 31, 1) {real, imag} */,
  {32'h461ade47, 32'h00000000} /* (12, 31, 0) {real, imag} */,
  {32'h462ca885, 32'h00000000} /* (12, 30, 31) {real, imag} */,
  {32'h4641b90d, 32'h00000000} /* (12, 30, 30) {real, imag} */,
  {32'h46332e75, 32'h00000000} /* (12, 30, 29) {real, imag} */,
  {32'h46358236, 32'h00000000} /* (12, 30, 28) {real, imag} */,
  {32'h463f7b92, 32'h00000000} /* (12, 30, 27) {real, imag} */,
  {32'h46375f0e, 32'h00000000} /* (12, 30, 26) {real, imag} */,
  {32'h46312a6a, 32'h00000000} /* (12, 30, 25) {real, imag} */,
  {32'h4625a43b, 32'h00000000} /* (12, 30, 24) {real, imag} */,
  {32'h4617ae6b, 32'h00000000} /* (12, 30, 23) {real, imag} */,
  {32'h46092a9c, 32'h00000000} /* (12, 30, 22) {real, imag} */,
  {32'h45973252, 32'h00000000} /* (12, 30, 21) {real, imag} */,
  {32'h44ec1450, 32'h00000000} /* (12, 30, 20) {real, imag} */,
  {32'hc49ec160, 32'h00000000} /* (12, 30, 19) {real, imag} */,
  {32'hc529a742, 32'h00000000} /* (12, 30, 18) {real, imag} */,
  {32'hc5707dd6, 32'h00000000} /* (12, 30, 17) {real, imag} */,
  {32'hc59702af, 32'h00000000} /* (12, 30, 16) {real, imag} */,
  {32'hc5b85b06, 32'h00000000} /* (12, 30, 15) {real, imag} */,
  {32'hc5b90b9a, 32'h00000000} /* (12, 30, 14) {real, imag} */,
  {32'hc5a42276, 32'h00000000} /* (12, 30, 13) {real, imag} */,
  {32'hc58ec0fe, 32'h00000000} /* (12, 30, 12) {real, imag} */,
  {32'hc504b252, 32'h00000000} /* (12, 30, 11) {real, imag} */,
  {32'h449e9df8, 32'h00000000} /* (12, 30, 10) {real, imag} */,
  {32'h4532f68a, 32'h00000000} /* (12, 30, 9) {real, imag} */,
  {32'h458c37b2, 32'h00000000} /* (12, 30, 8) {real, imag} */,
  {32'h45b80e02, 32'h00000000} /* (12, 30, 7) {real, imag} */,
  {32'h45e7e4a0, 32'h00000000} /* (12, 30, 6) {real, imag} */,
  {32'h460ca7ff, 32'h00000000} /* (12, 30, 5) {real, imag} */,
  {32'h46227ecb, 32'h00000000} /* (12, 30, 4) {real, imag} */,
  {32'h4626e5fc, 32'h00000000} /* (12, 30, 3) {real, imag} */,
  {32'h462d169c, 32'h00000000} /* (12, 30, 2) {real, imag} */,
  {32'h461fc62a, 32'h00000000} /* (12, 30, 1) {real, imag} */,
  {32'h46215684, 32'h00000000} /* (12, 30, 0) {real, imag} */,
  {32'h462e09ca, 32'h00000000} /* (12, 29, 31) {real, imag} */,
  {32'h464a65f8, 32'h00000000} /* (12, 29, 30) {real, imag} */,
  {32'h46392d3c, 32'h00000000} /* (12, 29, 29) {real, imag} */,
  {32'h463c8473, 32'h00000000} /* (12, 29, 28) {real, imag} */,
  {32'h463b3a70, 32'h00000000} /* (12, 29, 27) {real, imag} */,
  {32'h463542ba, 32'h00000000} /* (12, 29, 26) {real, imag} */,
  {32'h4639316d, 32'h00000000} /* (12, 29, 25) {real, imag} */,
  {32'h4623814a, 32'h00000000} /* (12, 29, 24) {real, imag} */,
  {32'h46213797, 32'h00000000} /* (12, 29, 23) {real, imag} */,
  {32'h45fadcdd, 32'h00000000} /* (12, 29, 22) {real, imag} */,
  {32'h458df027, 32'h00000000} /* (12, 29, 21) {real, imag} */,
  {32'h442fddf0, 32'h00000000} /* (12, 29, 20) {real, imag} */,
  {32'hc525f3b0, 32'h00000000} /* (12, 29, 19) {real, imag} */,
  {32'hc5835155, 32'h00000000} /* (12, 29, 18) {real, imag} */,
  {32'hc59d747e, 32'h00000000} /* (12, 29, 17) {real, imag} */,
  {32'hc5d08c9e, 32'h00000000} /* (12, 29, 16) {real, imag} */,
  {32'hc5ca8337, 32'h00000000} /* (12, 29, 15) {real, imag} */,
  {32'hc5ce8de3, 32'h00000000} /* (12, 29, 14) {real, imag} */,
  {32'hc5cce575, 32'h00000000} /* (12, 29, 13) {real, imag} */,
  {32'hc57acef4, 32'h00000000} /* (12, 29, 12) {real, imag} */,
  {32'hc4eb4974, 32'h00000000} /* (12, 29, 11) {real, imag} */,
  {32'h442e6d40, 32'h00000000} /* (12, 29, 10) {real, imag} */,
  {32'h454e07b4, 32'h00000000} /* (12, 29, 9) {real, imag} */,
  {32'h45a6f3ed, 32'h00000000} /* (12, 29, 8) {real, imag} */,
  {32'h45f22942, 32'h00000000} /* (12, 29, 7) {real, imag} */,
  {32'h461122be, 32'h00000000} /* (12, 29, 6) {real, imag} */,
  {32'h461de248, 32'h00000000} /* (12, 29, 5) {real, imag} */,
  {32'h461f4ddb, 32'h00000000} /* (12, 29, 4) {real, imag} */,
  {32'h463851aa, 32'h00000000} /* (12, 29, 3) {real, imag} */,
  {32'h46296724, 32'h00000000} /* (12, 29, 2) {real, imag} */,
  {32'h462d5c39, 32'h00000000} /* (12, 29, 1) {real, imag} */,
  {32'h4626e39b, 32'h00000000} /* (12, 29, 0) {real, imag} */,
  {32'h462cbe48, 32'h00000000} /* (12, 28, 31) {real, imag} */,
  {32'h464d0d98, 32'h00000000} /* (12, 28, 30) {real, imag} */,
  {32'h4650ece8, 32'h00000000} /* (12, 28, 29) {real, imag} */,
  {32'h463ec02b, 32'h00000000} /* (12, 28, 28) {real, imag} */,
  {32'h463da6ee, 32'h00000000} /* (12, 28, 27) {real, imag} */,
  {32'h4646e254, 32'h00000000} /* (12, 28, 26) {real, imag} */,
  {32'h46306e2c, 32'h00000000} /* (12, 28, 25) {real, imag} */,
  {32'h462093c0, 32'h00000000} /* (12, 28, 24) {real, imag} */,
  {32'h461ca2f5, 32'h00000000} /* (12, 28, 23) {real, imag} */,
  {32'h45c7f0e2, 32'h00000000} /* (12, 28, 22) {real, imag} */,
  {32'h45639ab2, 32'h00000000} /* (12, 28, 21) {real, imag} */,
  {32'hc4251e48, 32'h00000000} /* (12, 28, 20) {real, imag} */,
  {32'hc556c74e, 32'h00000000} /* (12, 28, 19) {real, imag} */,
  {32'hc5afeca0, 32'h00000000} /* (12, 28, 18) {real, imag} */,
  {32'hc5d9b670, 32'h00000000} /* (12, 28, 17) {real, imag} */,
  {32'hc5e80b38, 32'h00000000} /* (12, 28, 16) {real, imag} */,
  {32'hc5de7c61, 32'h00000000} /* (12, 28, 15) {real, imag} */,
  {32'hc5c7fcd8, 32'h00000000} /* (12, 28, 14) {real, imag} */,
  {32'hc5cd6653, 32'h00000000} /* (12, 28, 13) {real, imag} */,
  {32'hc59dff0e, 32'h00000000} /* (12, 28, 12) {real, imag} */,
  {32'hc4dc645c, 32'h00000000} /* (12, 28, 11) {real, imag} */,
  {32'h444cd268, 32'h00000000} /* (12, 28, 10) {real, imag} */,
  {32'h45735656, 32'h00000000} /* (12, 28, 9) {real, imag} */,
  {32'h45bb3854, 32'h00000000} /* (12, 28, 8) {real, imag} */,
  {32'h45f6fa06, 32'h00000000} /* (12, 28, 7) {real, imag} */,
  {32'h461a7477, 32'h00000000} /* (12, 28, 6) {real, imag} */,
  {32'h461b1306, 32'h00000000} /* (12, 28, 5) {real, imag} */,
  {32'h46374ec4, 32'h00000000} /* (12, 28, 4) {real, imag} */,
  {32'h46221de2, 32'h00000000} /* (12, 28, 3) {real, imag} */,
  {32'h462f096a, 32'h00000000} /* (12, 28, 2) {real, imag} */,
  {32'h4633a5f4, 32'h00000000} /* (12, 28, 1) {real, imag} */,
  {32'h462b62a6, 32'h00000000} /* (12, 28, 0) {real, imag} */,
  {32'h462cb7a2, 32'h00000000} /* (12, 27, 31) {real, imag} */,
  {32'h46538e14, 32'h00000000} /* (12, 27, 30) {real, imag} */,
  {32'h4650b774, 32'h00000000} /* (12, 27, 29) {real, imag} */,
  {32'h464dcdbc, 32'h00000000} /* (12, 27, 28) {real, imag} */,
  {32'h46482235, 32'h00000000} /* (12, 27, 27) {real, imag} */,
  {32'h4635ff18, 32'h00000000} /* (12, 27, 26) {real, imag} */,
  {32'h462714ac, 32'h00000000} /* (12, 27, 25) {real, imag} */,
  {32'h461b46fb, 32'h00000000} /* (12, 27, 24) {real, imag} */,
  {32'h46038db8, 32'h00000000} /* (12, 27, 23) {real, imag} */,
  {32'h45c4a7eb, 32'h00000000} /* (12, 27, 22) {real, imag} */,
  {32'h454099e2, 32'h00000000} /* (12, 27, 21) {real, imag} */,
  {32'hc440fa28, 32'h00000000} /* (12, 27, 20) {real, imag} */,
  {32'hc583aa28, 32'h00000000} /* (12, 27, 19) {real, imag} */,
  {32'hc5d3178f, 32'h00000000} /* (12, 27, 18) {real, imag} */,
  {32'hc5df89b4, 32'h00000000} /* (12, 27, 17) {real, imag} */,
  {32'hc5f42c72, 32'h00000000} /* (12, 27, 16) {real, imag} */,
  {32'hc609b532, 32'h00000000} /* (12, 27, 15) {real, imag} */,
  {32'hc5e7d218, 32'h00000000} /* (12, 27, 14) {real, imag} */,
  {32'hc5976340, 32'h00000000} /* (12, 27, 13) {real, imag} */,
  {32'hc59b4275, 32'h00000000} /* (12, 27, 12) {real, imag} */,
  {32'hc4f87358, 32'h00000000} /* (12, 27, 11) {real, imag} */,
  {32'h44845e58, 32'h00000000} /* (12, 27, 10) {real, imag} */,
  {32'h45832c8c, 32'h00000000} /* (12, 27, 9) {real, imag} */,
  {32'h45dc944a, 32'h00000000} /* (12, 27, 8) {real, imag} */,
  {32'h45f4f34b, 32'h00000000} /* (12, 27, 7) {real, imag} */,
  {32'h46216046, 32'h00000000} /* (12, 27, 6) {real, imag} */,
  {32'h4626b0e8, 32'h00000000} /* (12, 27, 5) {real, imag} */,
  {32'h461cf07e, 32'h00000000} /* (12, 27, 4) {real, imag} */,
  {32'h4626e4cc, 32'h00000000} /* (12, 27, 3) {real, imag} */,
  {32'h4626869c, 32'h00000000} /* (12, 27, 2) {real, imag} */,
  {32'h4632c7b4, 32'h00000000} /* (12, 27, 1) {real, imag} */,
  {32'h46320f81, 32'h00000000} /* (12, 27, 0) {real, imag} */,
  {32'h4626cd6f, 32'h00000000} /* (12, 26, 31) {real, imag} */,
  {32'h463622c2, 32'h00000000} /* (12, 26, 30) {real, imag} */,
  {32'h463c1432, 32'h00000000} /* (12, 26, 29) {real, imag} */,
  {32'h4639e13a, 32'h00000000} /* (12, 26, 28) {real, imag} */,
  {32'h463a9c5a, 32'h00000000} /* (12, 26, 27) {real, imag} */,
  {32'h4630ca66, 32'h00000000} /* (12, 26, 26) {real, imag} */,
  {32'h463395d7, 32'h00000000} /* (12, 26, 25) {real, imag} */,
  {32'h4611af16, 32'h00000000} /* (12, 26, 24) {real, imag} */,
  {32'h45f371d9, 32'h00000000} /* (12, 26, 23) {real, imag} */,
  {32'h45c209b8, 32'h00000000} /* (12, 26, 22) {real, imag} */,
  {32'h4527dbf2, 32'h00000000} /* (12, 26, 21) {real, imag} */,
  {32'hc45652f8, 32'h00000000} /* (12, 26, 20) {real, imag} */,
  {32'hc57f5962, 32'h00000000} /* (12, 26, 19) {real, imag} */,
  {32'hc5b296c0, 32'h00000000} /* (12, 26, 18) {real, imag} */,
  {32'hc5d71ee5, 32'h00000000} /* (12, 26, 17) {real, imag} */,
  {32'hc5fea058, 32'h00000000} /* (12, 26, 16) {real, imag} */,
  {32'hc5ff870a, 32'h00000000} /* (12, 26, 15) {real, imag} */,
  {32'hc5f0e064, 32'h00000000} /* (12, 26, 14) {real, imag} */,
  {32'hc5b3e9e0, 32'h00000000} /* (12, 26, 13) {real, imag} */,
  {32'hc5771932, 32'h00000000} /* (12, 26, 12) {real, imag} */,
  {32'hc5177876, 32'h00000000} /* (12, 26, 11) {real, imag} */,
  {32'h44ab5f80, 32'h00000000} /* (12, 26, 10) {real, imag} */,
  {32'h45b2676a, 32'h00000000} /* (12, 26, 9) {real, imag} */,
  {32'h45f4f178, 32'h00000000} /* (12, 26, 8) {real, imag} */,
  {32'h45f5a763, 32'h00000000} /* (12, 26, 7) {real, imag} */,
  {32'h460b1d68, 32'h00000000} /* (12, 26, 6) {real, imag} */,
  {32'h460f8fd0, 32'h00000000} /* (12, 26, 5) {real, imag} */,
  {32'h461afbae, 32'h00000000} /* (12, 26, 4) {real, imag} */,
  {32'h4625c878, 32'h00000000} /* (12, 26, 3) {real, imag} */,
  {32'h4621248e, 32'h00000000} /* (12, 26, 2) {real, imag} */,
  {32'h462bce6e, 32'h00000000} /* (12, 26, 1) {real, imag} */,
  {32'h462494fe, 32'h00000000} /* (12, 26, 0) {real, imag} */,
  {32'h4615f49a, 32'h00000000} /* (12, 25, 31) {real, imag} */,
  {32'h46277620, 32'h00000000} /* (12, 25, 30) {real, imag} */,
  {32'h46251e8b, 32'h00000000} /* (12, 25, 29) {real, imag} */,
  {32'h46327d63, 32'h00000000} /* (12, 25, 28) {real, imag} */,
  {32'h462a4d0a, 32'h00000000} /* (12, 25, 27) {real, imag} */,
  {32'h461ad10d, 32'h00000000} /* (12, 25, 26) {real, imag} */,
  {32'h462d0df2, 32'h00000000} /* (12, 25, 25) {real, imag} */,
  {32'h46128f2e, 32'h00000000} /* (12, 25, 24) {real, imag} */,
  {32'h45cb9830, 32'h00000000} /* (12, 25, 23) {real, imag} */,
  {32'h45a72df6, 32'h00000000} /* (12, 25, 22) {real, imag} */,
  {32'h4518f0d6, 32'h00000000} /* (12, 25, 21) {real, imag} */,
  {32'hc4ee46f4, 32'h00000000} /* (12, 25, 20) {real, imag} */,
  {32'hc567f000, 32'h00000000} /* (12, 25, 19) {real, imag} */,
  {32'hc5bca617, 32'h00000000} /* (12, 25, 18) {real, imag} */,
  {32'hc5f248a6, 32'h00000000} /* (12, 25, 17) {real, imag} */,
  {32'hc6067ec2, 32'h00000000} /* (12, 25, 16) {real, imag} */,
  {32'hc5e5d32f, 32'h00000000} /* (12, 25, 15) {real, imag} */,
  {32'hc5b73017, 32'h00000000} /* (12, 25, 14) {real, imag} */,
  {32'hc5baa1e2, 32'h00000000} /* (12, 25, 13) {real, imag} */,
  {32'hc584e888, 32'h00000000} /* (12, 25, 12) {real, imag} */,
  {32'hc51e75c6, 32'h00000000} /* (12, 25, 11) {real, imag} */,
  {32'h44b343e8, 32'h00000000} /* (12, 25, 10) {real, imag} */,
  {32'h45a0dd1c, 32'h00000000} /* (12, 25, 9) {real, imag} */,
  {32'h45de4e1b, 32'h00000000} /* (12, 25, 8) {real, imag} */,
  {32'h45e6a706, 32'h00000000} /* (12, 25, 7) {real, imag} */,
  {32'h46055710, 32'h00000000} /* (12, 25, 6) {real, imag} */,
  {32'h460609ba, 32'h00000000} /* (12, 25, 5) {real, imag} */,
  {32'h46130b5a, 32'h00000000} /* (12, 25, 4) {real, imag} */,
  {32'h4613ba06, 32'h00000000} /* (12, 25, 3) {real, imag} */,
  {32'h4625ea28, 32'h00000000} /* (12, 25, 2) {real, imag} */,
  {32'h461c3c59, 32'h00000000} /* (12, 25, 1) {real, imag} */,
  {32'h4610ff0a, 32'h00000000} /* (12, 25, 0) {real, imag} */,
  {32'h45ffe039, 32'h00000000} /* (12, 24, 31) {real, imag} */,
  {32'h46069ca5, 32'h00000000} /* (12, 24, 30) {real, imag} */,
  {32'h461a6e0c, 32'h00000000} /* (12, 24, 29) {real, imag} */,
  {32'h461785fa, 32'h00000000} /* (12, 24, 28) {real, imag} */,
  {32'h460dcfda, 32'h00000000} /* (12, 24, 27) {real, imag} */,
  {32'h461240a6, 32'h00000000} /* (12, 24, 26) {real, imag} */,
  {32'h4612aa6e, 32'h00000000} /* (12, 24, 25) {real, imag} */,
  {32'h45f8bc26, 32'h00000000} /* (12, 24, 24) {real, imag} */,
  {32'h45a1204c, 32'h00000000} /* (12, 24, 23) {real, imag} */,
  {32'h458f2e79, 32'h00000000} /* (12, 24, 22) {real, imag} */,
  {32'h44ecde6e, 32'h00000000} /* (12, 24, 21) {real, imag} */,
  {32'hc513f089, 32'h00000000} /* (12, 24, 20) {real, imag} */,
  {32'hc56d615f, 32'h00000000} /* (12, 24, 19) {real, imag} */,
  {32'hc598417e, 32'h00000000} /* (12, 24, 18) {real, imag} */,
  {32'hc5dfc1ae, 32'h00000000} /* (12, 24, 17) {real, imag} */,
  {32'hc5e9766a, 32'h00000000} /* (12, 24, 16) {real, imag} */,
  {32'hc5d2f9f3, 32'h00000000} /* (12, 24, 15) {real, imag} */,
  {32'hc5bd5212, 32'h00000000} /* (12, 24, 14) {real, imag} */,
  {32'hc5a2bff9, 32'h00000000} /* (12, 24, 13) {real, imag} */,
  {32'hc58b8c90, 32'h00000000} /* (12, 24, 12) {real, imag} */,
  {32'hc53c9721, 32'h00000000} /* (12, 24, 11) {real, imag} */,
  {32'h4442aab8, 32'h00000000} /* (12, 24, 10) {real, imag} */,
  {32'h45a484ba, 32'h00000000} /* (12, 24, 9) {real, imag} */,
  {32'h45c2d8d4, 32'h00000000} /* (12, 24, 8) {real, imag} */,
  {32'h45e6ea4a, 32'h00000000} /* (12, 24, 7) {real, imag} */,
  {32'h45eea157, 32'h00000000} /* (12, 24, 6) {real, imag} */,
  {32'h46017155, 32'h00000000} /* (12, 24, 5) {real, imag} */,
  {32'h46053f11, 32'h00000000} /* (12, 24, 4) {real, imag} */,
  {32'h46016052, 32'h00000000} /* (12, 24, 3) {real, imag} */,
  {32'h460a9123, 32'h00000000} /* (12, 24, 2) {real, imag} */,
  {32'h46054044, 32'h00000000} /* (12, 24, 1) {real, imag} */,
  {32'h4603be7a, 32'h00000000} /* (12, 24, 0) {real, imag} */,
  {32'h45c5b406, 32'h00000000} /* (12, 23, 31) {real, imag} */,
  {32'h45fab8d0, 32'h00000000} /* (12, 23, 30) {real, imag} */,
  {32'h4603d3c5, 32'h00000000} /* (12, 23, 29) {real, imag} */,
  {32'h45e6d383, 32'h00000000} /* (12, 23, 28) {real, imag} */,
  {32'h45f2505c, 32'h00000000} /* (12, 23, 27) {real, imag} */,
  {32'h45df451c, 32'h00000000} /* (12, 23, 26) {real, imag} */,
  {32'h45d3207b, 32'h00000000} /* (12, 23, 25) {real, imag} */,
  {32'h45b8707a, 32'h00000000} /* (12, 23, 24) {real, imag} */,
  {32'h45b6f797, 32'h00000000} /* (12, 23, 23) {real, imag} */,
  {32'h455d9ae4, 32'h00000000} /* (12, 23, 22) {real, imag} */,
  {32'h446b5e3c, 32'h00000000} /* (12, 23, 21) {real, imag} */,
  {32'hc4b1c530, 32'h00000000} /* (12, 23, 20) {real, imag} */,
  {32'hc56785c8, 32'h00000000} /* (12, 23, 19) {real, imag} */,
  {32'hc5a07dab, 32'h00000000} /* (12, 23, 18) {real, imag} */,
  {32'hc598aaba, 32'h00000000} /* (12, 23, 17) {real, imag} */,
  {32'hc5ad191e, 32'h00000000} /* (12, 23, 16) {real, imag} */,
  {32'hc5a3a3e8, 32'h00000000} /* (12, 23, 15) {real, imag} */,
  {32'hc5adbd1a, 32'h00000000} /* (12, 23, 14) {real, imag} */,
  {32'hc59b3f34, 32'h00000000} /* (12, 23, 13) {real, imag} */,
  {32'hc559b65e, 32'h00000000} /* (12, 23, 12) {real, imag} */,
  {32'hc51dfeb0, 32'h00000000} /* (12, 23, 11) {real, imag} */,
  {32'h43c3c200, 32'h00000000} /* (12, 23, 10) {real, imag} */,
  {32'h4545162a, 32'h00000000} /* (12, 23, 9) {real, imag} */,
  {32'h4593a032, 32'h00000000} /* (12, 23, 8) {real, imag} */,
  {32'h45aeb5d1, 32'h00000000} /* (12, 23, 7) {real, imag} */,
  {32'h45c767f2, 32'h00000000} /* (12, 23, 6) {real, imag} */,
  {32'h45cc9e7a, 32'h00000000} /* (12, 23, 5) {real, imag} */,
  {32'h45e0c82a, 32'h00000000} /* (12, 23, 4) {real, imag} */,
  {32'h45d62386, 32'h00000000} /* (12, 23, 3) {real, imag} */,
  {32'h45cd2771, 32'h00000000} /* (12, 23, 2) {real, imag} */,
  {32'h45d4c4be, 32'h00000000} /* (12, 23, 1) {real, imag} */,
  {32'h45c5ec5c, 32'h00000000} /* (12, 23, 0) {real, imag} */,
  {32'h459157ea, 32'h00000000} /* (12, 22, 31) {real, imag} */,
  {32'h45bc5b54, 32'h00000000} /* (12, 22, 30) {real, imag} */,
  {32'h45a85b7d, 32'h00000000} /* (12, 22, 29) {real, imag} */,
  {32'h45a010bc, 32'h00000000} /* (12, 22, 28) {real, imag} */,
  {32'h4598009a, 32'h00000000} /* (12, 22, 27) {real, imag} */,
  {32'h459076c7, 32'h00000000} /* (12, 22, 26) {real, imag} */,
  {32'h458b0111, 32'h00000000} /* (12, 22, 25) {real, imag} */,
  {32'h456ca7d2, 32'h00000000} /* (12, 22, 24) {real, imag} */,
  {32'h4595762b, 32'h00000000} /* (12, 22, 23) {real, imag} */,
  {32'h4551f799, 32'h00000000} /* (12, 22, 22) {real, imag} */,
  {32'h429e2980, 32'h00000000} /* (12, 22, 21) {real, imag} */,
  {32'hc4f7870c, 32'h00000000} /* (12, 22, 20) {real, imag} */,
  {32'hc50541d5, 32'h00000000} /* (12, 22, 19) {real, imag} */,
  {32'hc579421b, 32'h00000000} /* (12, 22, 18) {real, imag} */,
  {32'hc5839fc6, 32'h00000000} /* (12, 22, 17) {real, imag} */,
  {32'hc5743c8a, 32'h00000000} /* (12, 22, 16) {real, imag} */,
  {32'hc53308e1, 32'h00000000} /* (12, 22, 15) {real, imag} */,
  {32'hc55d2958, 32'h00000000} /* (12, 22, 14) {real, imag} */,
  {32'hc55165fa, 32'h00000000} /* (12, 22, 13) {real, imag} */,
  {32'hc5910398, 32'h00000000} /* (12, 22, 12) {real, imag} */,
  {32'hc52ed3a8, 32'h00000000} /* (12, 22, 11) {real, imag} */,
  {32'h4315d1a0, 32'h00000000} /* (12, 22, 10) {real, imag} */,
  {32'h45602190, 32'h00000000} /* (12, 22, 9) {real, imag} */,
  {32'h456aebde, 32'h00000000} /* (12, 22, 8) {real, imag} */,
  {32'h458ca8a1, 32'h00000000} /* (12, 22, 7) {real, imag} */,
  {32'h457be1a7, 32'h00000000} /* (12, 22, 6) {real, imag} */,
  {32'h45889776, 32'h00000000} /* (12, 22, 5) {real, imag} */,
  {32'h4599536a, 32'h00000000} /* (12, 22, 4) {real, imag} */,
  {32'h459cbf3a, 32'h00000000} /* (12, 22, 3) {real, imag} */,
  {32'h45aa76dd, 32'h00000000} /* (12, 22, 2) {real, imag} */,
  {32'h45a8e0e8, 32'h00000000} /* (12, 22, 1) {real, imag} */,
  {32'h458d21bf, 32'h00000000} /* (12, 22, 0) {real, imag} */,
  {32'h44e58640, 32'h00000000} /* (12, 21, 31) {real, imag} */,
  {32'h44e322ba, 32'h00000000} /* (12, 21, 30) {real, imag} */,
  {32'h44bb16fe, 32'h00000000} /* (12, 21, 29) {real, imag} */,
  {32'h451386f8, 32'h00000000} /* (12, 21, 28) {real, imag} */,
  {32'h448efe26, 32'h00000000} /* (12, 21, 27) {real, imag} */,
  {32'h44b11fa4, 32'h00000000} /* (12, 21, 26) {real, imag} */,
  {32'h44bb4bef, 32'h00000000} /* (12, 21, 25) {real, imag} */,
  {32'h44abdb9d, 32'h00000000} /* (12, 21, 24) {real, imag} */,
  {32'h4462d756, 32'h00000000} /* (12, 21, 23) {real, imag} */,
  {32'h449fe140, 32'h00000000} /* (12, 21, 22) {real, imag} */,
  {32'hc285a3d8, 32'h00000000} /* (12, 21, 21) {real, imag} */,
  {32'hc4ad92ab, 32'h00000000} /* (12, 21, 20) {real, imag} */,
  {32'hc4b11364, 32'h00000000} /* (12, 21, 19) {real, imag} */,
  {32'hc3a5d79c, 32'h00000000} /* (12, 21, 18) {real, imag} */,
  {32'hc4b71c65, 32'h00000000} /* (12, 21, 17) {real, imag} */,
  {32'hc444cc9d, 32'h00000000} /* (12, 21, 16) {real, imag} */,
  {32'hc40d0300, 32'h00000000} /* (12, 21, 15) {real, imag} */,
  {32'hc41bcf1c, 32'h00000000} /* (12, 21, 14) {real, imag} */,
  {32'hc498e8ac, 32'h00000000} /* (12, 21, 13) {real, imag} */,
  {32'hc49856ca, 32'h00000000} /* (12, 21, 12) {real, imag} */,
  {32'hc48197dc, 32'h00000000} /* (12, 21, 11) {real, imag} */,
  {32'h446e77d8, 32'h00000000} /* (12, 21, 10) {real, imag} */,
  {32'h44a7932b, 32'h00000000} /* (12, 21, 9) {real, imag} */,
  {32'h44ef8dc3, 32'h00000000} /* (12, 21, 8) {real, imag} */,
  {32'h44e496ab, 32'h00000000} /* (12, 21, 7) {real, imag} */,
  {32'h449fce84, 32'h00000000} /* (12, 21, 6) {real, imag} */,
  {32'h4492f798, 32'h00000000} /* (12, 21, 5) {real, imag} */,
  {32'h44c3453f, 32'h00000000} /* (12, 21, 4) {real, imag} */,
  {32'h44dc1294, 32'h00000000} /* (12, 21, 3) {real, imag} */,
  {32'h4518e6f4, 32'h00000000} /* (12, 21, 2) {real, imag} */,
  {32'h44e1ca37, 32'h00000000} /* (12, 21, 1) {real, imag} */,
  {32'h44904a60, 32'h00000000} /* (12, 21, 0) {real, imag} */,
  {32'hc500ff60, 32'h00000000} /* (12, 20, 31) {real, imag} */,
  {32'hc54aef48, 32'h00000000} /* (12, 20, 30) {real, imag} */,
  {32'hc52065b3, 32'h00000000} /* (12, 20, 29) {real, imag} */,
  {32'hc52e1c4a, 32'h00000000} /* (12, 20, 28) {real, imag} */,
  {32'hc4feaf00, 32'h00000000} /* (12, 20, 27) {real, imag} */,
  {32'hc4e0d863, 32'h00000000} /* (12, 20, 26) {real, imag} */,
  {32'hc512db39, 32'h00000000} /* (12, 20, 25) {real, imag} */,
  {32'hc5048040, 32'h00000000} /* (12, 20, 24) {real, imag} */,
  {32'hc5297608, 32'h00000000} /* (12, 20, 23) {real, imag} */,
  {32'hc54b5a21, 32'h00000000} /* (12, 20, 22) {real, imag} */,
  {32'hc40931f2, 32'h00000000} /* (12, 20, 21) {real, imag} */,
  {32'h440c9c6d, 32'h00000000} /* (12, 20, 20) {real, imag} */,
  {32'h44b07e4d, 32'h00000000} /* (12, 20, 19) {real, imag} */,
  {32'h45022a61, 32'h00000000} /* (12, 20, 18) {real, imag} */,
  {32'h45573380, 32'h00000000} /* (12, 20, 17) {real, imag} */,
  {32'h44fb2c09, 32'h00000000} /* (12, 20, 16) {real, imag} */,
  {32'h452e3200, 32'h00000000} /* (12, 20, 15) {real, imag} */,
  {32'h451074d4, 32'h00000000} /* (12, 20, 14) {real, imag} */,
  {32'h44dcc7ea, 32'h00000000} /* (12, 20, 13) {real, imag} */,
  {32'h4508292c, 32'h00000000} /* (12, 20, 12) {real, imag} */,
  {32'h445d1a20, 32'h00000000} /* (12, 20, 11) {real, imag} */,
  {32'hc3bd4634, 32'h00000000} /* (12, 20, 10) {real, imag} */,
  {32'hc507cd1b, 32'h00000000} /* (12, 20, 9) {real, imag} */,
  {32'hc4a93390, 32'h00000000} /* (12, 20, 8) {real, imag} */,
  {32'hc4f93fc1, 32'h00000000} /* (12, 20, 7) {real, imag} */,
  {32'hc50e4837, 32'h00000000} /* (12, 20, 6) {real, imag} */,
  {32'hc522ca72, 32'h00000000} /* (12, 20, 5) {real, imag} */,
  {32'hc507d5f7, 32'h00000000} /* (12, 20, 4) {real, imag} */,
  {32'hc521115e, 32'h00000000} /* (12, 20, 3) {real, imag} */,
  {32'hc4fe67f6, 32'h00000000} /* (12, 20, 2) {real, imag} */,
  {32'hc5054e4a, 32'h00000000} /* (12, 20, 1) {real, imag} */,
  {32'hc4e088a9, 32'h00000000} /* (12, 20, 0) {real, imag} */,
  {32'hc56ee0b2, 32'h00000000} /* (12, 19, 31) {real, imag} */,
  {32'hc5b10fe4, 32'h00000000} /* (12, 19, 30) {real, imag} */,
  {32'hc5928878, 32'h00000000} /* (12, 19, 29) {real, imag} */,
  {32'hc5993f53, 32'h00000000} /* (12, 19, 28) {real, imag} */,
  {32'hc591dc9c, 32'h00000000} /* (12, 19, 27) {real, imag} */,
  {32'hc59f6429, 32'h00000000} /* (12, 19, 26) {real, imag} */,
  {32'hc591785c, 32'h00000000} /* (12, 19, 25) {real, imag} */,
  {32'hc5785a85, 32'h00000000} /* (12, 19, 24) {real, imag} */,
  {32'hc5880020, 32'h00000000} /* (12, 19, 23) {real, imag} */,
  {32'hc546559b, 32'h00000000} /* (12, 19, 22) {real, imag} */,
  {32'hc4c41d21, 32'h00000000} /* (12, 19, 21) {real, imag} */,
  {32'h44dee493, 32'h00000000} /* (12, 19, 20) {real, imag} */,
  {32'h453b9737, 32'h00000000} /* (12, 19, 19) {real, imag} */,
  {32'h45684359, 32'h00000000} /* (12, 19, 18) {real, imag} */,
  {32'h45710aa0, 32'h00000000} /* (12, 19, 17) {real, imag} */,
  {32'h4596fa64, 32'h00000000} /* (12, 19, 16) {real, imag} */,
  {32'h45b19b51, 32'h00000000} /* (12, 19, 15) {real, imag} */,
  {32'h458e6b14, 32'h00000000} /* (12, 19, 14) {real, imag} */,
  {32'h4565f8b0, 32'h00000000} /* (12, 19, 13) {real, imag} */,
  {32'h452b9754, 32'h00000000} /* (12, 19, 12) {real, imag} */,
  {32'h44c63942, 32'h00000000} /* (12, 19, 11) {real, imag} */,
  {32'hc4c4e78d, 32'h00000000} /* (12, 19, 10) {real, imag} */,
  {32'hc54475f3, 32'h00000000} /* (12, 19, 9) {real, imag} */,
  {32'hc52e09e9, 32'h00000000} /* (12, 19, 8) {real, imag} */,
  {32'hc58bc028, 32'h00000000} /* (12, 19, 7) {real, imag} */,
  {32'hc5801198, 32'h00000000} /* (12, 19, 6) {real, imag} */,
  {32'hc5ad24da, 32'h00000000} /* (12, 19, 5) {real, imag} */,
  {32'hc5af1b37, 32'h00000000} /* (12, 19, 4) {real, imag} */,
  {32'hc5812678, 32'h00000000} /* (12, 19, 3) {real, imag} */,
  {32'hc5951e58, 32'h00000000} /* (12, 19, 2) {real, imag} */,
  {32'hc5a2191a, 32'h00000000} /* (12, 19, 1) {real, imag} */,
  {32'hc590efcc, 32'h00000000} /* (12, 19, 0) {real, imag} */,
  {32'hc5c0deb0, 32'h00000000} /* (12, 18, 31) {real, imag} */,
  {32'hc5d0bdae, 32'h00000000} /* (12, 18, 30) {real, imag} */,
  {32'hc5fab1e2, 32'h00000000} /* (12, 18, 29) {real, imag} */,
  {32'hc5e8c6aa, 32'h00000000} /* (12, 18, 28) {real, imag} */,
  {32'hc5dfeed7, 32'h00000000} /* (12, 18, 27) {real, imag} */,
  {32'hc5db0060, 32'h00000000} /* (12, 18, 26) {real, imag} */,
  {32'hc5b4c741, 32'h00000000} /* (12, 18, 25) {real, imag} */,
  {32'hc5bf4d95, 32'h00000000} /* (12, 18, 24) {real, imag} */,
  {32'hc5a8e454, 32'h00000000} /* (12, 18, 23) {real, imag} */,
  {32'hc56e7c1e, 32'h00000000} /* (12, 18, 22) {real, imag} */,
  {32'hc52880ea, 32'h00000000} /* (12, 18, 21) {real, imag} */,
  {32'h44e08cae, 32'h00000000} /* (12, 18, 20) {real, imag} */,
  {32'h454be414, 32'h00000000} /* (12, 18, 19) {real, imag} */,
  {32'h45bbedfe, 32'h00000000} /* (12, 18, 18) {real, imag} */,
  {32'h45af56d8, 32'h00000000} /* (12, 18, 17) {real, imag} */,
  {32'h45a83eb0, 32'h00000000} /* (12, 18, 16) {real, imag} */,
  {32'h45b18930, 32'h00000000} /* (12, 18, 15) {real, imag} */,
  {32'h45becf50, 32'h00000000} /* (12, 18, 14) {real, imag} */,
  {32'h45a4dde8, 32'h00000000} /* (12, 18, 13) {real, imag} */,
  {32'h455a42bf, 32'h00000000} /* (12, 18, 12) {real, imag} */,
  {32'h452030fe, 32'h00000000} /* (12, 18, 11) {real, imag} */,
  {32'hc4ad086a, 32'h00000000} /* (12, 18, 10) {real, imag} */,
  {32'hc57be706, 32'h00000000} /* (12, 18, 9) {real, imag} */,
  {32'hc5780776, 32'h00000000} /* (12, 18, 8) {real, imag} */,
  {32'hc5a198fc, 32'h00000000} /* (12, 18, 7) {real, imag} */,
  {32'hc5c5ca3b, 32'h00000000} /* (12, 18, 6) {real, imag} */,
  {32'hc5d5f135, 32'h00000000} /* (12, 18, 5) {real, imag} */,
  {32'hc5d04768, 32'h00000000} /* (12, 18, 4) {real, imag} */,
  {32'hc5db0712, 32'h00000000} /* (12, 18, 3) {real, imag} */,
  {32'hc5e11fac, 32'h00000000} /* (12, 18, 2) {real, imag} */,
  {32'hc5c103f8, 32'h00000000} /* (12, 18, 1) {real, imag} */,
  {32'hc5b8ae80, 32'h00000000} /* (12, 18, 0) {real, imag} */,
  {32'hc5cfb8f6, 32'h00000000} /* (12, 17, 31) {real, imag} */,
  {32'hc5f55292, 32'h00000000} /* (12, 17, 30) {real, imag} */,
  {32'hc6050a7c, 32'h00000000} /* (12, 17, 29) {real, imag} */,
  {32'hc6219c61, 32'h00000000} /* (12, 17, 28) {real, imag} */,
  {32'hc60b0b1c, 32'h00000000} /* (12, 17, 27) {real, imag} */,
  {32'hc5ec225a, 32'h00000000} /* (12, 17, 26) {real, imag} */,
  {32'hc5dde8da, 32'h00000000} /* (12, 17, 25) {real, imag} */,
  {32'hc5cfcc22, 32'h00000000} /* (12, 17, 24) {real, imag} */,
  {32'hc5c1bd06, 32'h00000000} /* (12, 17, 23) {real, imag} */,
  {32'hc5795fa8, 32'h00000000} /* (12, 17, 22) {real, imag} */,
  {32'hc4c3d858, 32'h00000000} /* (12, 17, 21) {real, imag} */,
  {32'h450f592c, 32'h00000000} /* (12, 17, 20) {real, imag} */,
  {32'h457ec6dc, 32'h00000000} /* (12, 17, 19) {real, imag} */,
  {32'h45b1fd1a, 32'h00000000} /* (12, 17, 18) {real, imag} */,
  {32'h45cc4666, 32'h00000000} /* (12, 17, 17) {real, imag} */,
  {32'h45d588a6, 32'h00000000} /* (12, 17, 16) {real, imag} */,
  {32'h45ee825c, 32'h00000000} /* (12, 17, 15) {real, imag} */,
  {32'h45c677c6, 32'h00000000} /* (12, 17, 14) {real, imag} */,
  {32'h45adaeb8, 32'h00000000} /* (12, 17, 13) {real, imag} */,
  {32'h459724f0, 32'h00000000} /* (12, 17, 12) {real, imag} */,
  {32'h44f09b94, 32'h00000000} /* (12, 17, 11) {real, imag} */,
  {32'hc4bdea28, 32'h00000000} /* (12, 17, 10) {real, imag} */,
  {32'hc53ea1c4, 32'h00000000} /* (12, 17, 9) {real, imag} */,
  {32'hc59e8eba, 32'h00000000} /* (12, 17, 8) {real, imag} */,
  {32'hc5c461d8, 32'h00000000} /* (12, 17, 7) {real, imag} */,
  {32'hc5dd63f8, 32'h00000000} /* (12, 17, 6) {real, imag} */,
  {32'hc5f0573e, 32'h00000000} /* (12, 17, 5) {real, imag} */,
  {32'hc60555a8, 32'h00000000} /* (12, 17, 4) {real, imag} */,
  {32'hc60ab21a, 32'h00000000} /* (12, 17, 3) {real, imag} */,
  {32'hc5f0016c, 32'h00000000} /* (12, 17, 2) {real, imag} */,
  {32'hc5d4a152, 32'h00000000} /* (12, 17, 1) {real, imag} */,
  {32'hc5dc3586, 32'h00000000} /* (12, 17, 0) {real, imag} */,
  {32'hc5f57d44, 32'h00000000} /* (12, 16, 31) {real, imag} */,
  {32'hc60997c1, 32'h00000000} /* (12, 16, 30) {real, imag} */,
  {32'hc60cd070, 32'h00000000} /* (12, 16, 29) {real, imag} */,
  {32'hc6084830, 32'h00000000} /* (12, 16, 28) {real, imag} */,
  {32'hc608eddc, 32'h00000000} /* (12, 16, 27) {real, imag} */,
  {32'hc60ae8ec, 32'h00000000} /* (12, 16, 26) {real, imag} */,
  {32'hc5fd77c2, 32'h00000000} /* (12, 16, 25) {real, imag} */,
  {32'hc5ef79fc, 32'h00000000} /* (12, 16, 24) {real, imag} */,
  {32'hc5cc7d04, 32'h00000000} /* (12, 16, 23) {real, imag} */,
  {32'hc5920383, 32'h00000000} /* (12, 16, 22) {real, imag} */,
  {32'hc3e6bae0, 32'h00000000} /* (12, 16, 21) {real, imag} */,
  {32'h45453c81, 32'h00000000} /* (12, 16, 20) {real, imag} */,
  {32'h459a9fb6, 32'h00000000} /* (12, 16, 19) {real, imag} */,
  {32'h45c6ecfe, 32'h00000000} /* (12, 16, 18) {real, imag} */,
  {32'h45d1f53e, 32'h00000000} /* (12, 16, 17) {real, imag} */,
  {32'h45f5da51, 32'h00000000} /* (12, 16, 16) {real, imag} */,
  {32'h45d5e7d8, 32'h00000000} /* (12, 16, 15) {real, imag} */,
  {32'h45e2be86, 32'h00000000} /* (12, 16, 14) {real, imag} */,
  {32'h45d24aad, 32'h00000000} /* (12, 16, 13) {real, imag} */,
  {32'h45973622, 32'h00000000} /* (12, 16, 12) {real, imag} */,
  {32'h44e074cc, 32'h00000000} /* (12, 16, 11) {real, imag} */,
  {32'hc49e846e, 32'h00000000} /* (12, 16, 10) {real, imag} */,
  {32'hc55b6975, 32'h00000000} /* (12, 16, 9) {real, imag} */,
  {32'hc58c9e16, 32'h00000000} /* (12, 16, 8) {real, imag} */,
  {32'hc5d5d01c, 32'h00000000} /* (12, 16, 7) {real, imag} */,
  {32'hc5f299c1, 32'h00000000} /* (12, 16, 6) {real, imag} */,
  {32'hc5fa4198, 32'h00000000} /* (12, 16, 5) {real, imag} */,
  {32'hc609a23d, 32'h00000000} /* (12, 16, 4) {real, imag} */,
  {32'hc60cd0ce, 32'h00000000} /* (12, 16, 3) {real, imag} */,
  {32'hc5e7ae1a, 32'h00000000} /* (12, 16, 2) {real, imag} */,
  {32'hc60597c0, 32'h00000000} /* (12, 16, 1) {real, imag} */,
  {32'hc60194d4, 32'h00000000} /* (12, 16, 0) {real, imag} */,
  {32'hc5faa28d, 32'h00000000} /* (12, 15, 31) {real, imag} */,
  {32'hc6037618, 32'h00000000} /* (12, 15, 30) {real, imag} */,
  {32'hc604ca89, 32'h00000000} /* (12, 15, 29) {real, imag} */,
  {32'hc61cbfca, 32'h00000000} /* (12, 15, 28) {real, imag} */,
  {32'hc60a9fc8, 32'h00000000} /* (12, 15, 27) {real, imag} */,
  {32'hc602fa66, 32'h00000000} /* (12, 15, 26) {real, imag} */,
  {32'hc601ea08, 32'h00000000} /* (12, 15, 25) {real, imag} */,
  {32'hc5ecbd53, 32'h00000000} /* (12, 15, 24) {real, imag} */,
  {32'hc5b25e51, 32'h00000000} /* (12, 15, 23) {real, imag} */,
  {32'hc567aaa2, 32'h00000000} /* (12, 15, 22) {real, imag} */,
  {32'hc41140e8, 32'h00000000} /* (12, 15, 21) {real, imag} */,
  {32'h4519924f, 32'h00000000} /* (12, 15, 20) {real, imag} */,
  {32'h4592f201, 32'h00000000} /* (12, 15, 19) {real, imag} */,
  {32'h45c5c8dd, 32'h00000000} /* (12, 15, 18) {real, imag} */,
  {32'h45dd955e, 32'h00000000} /* (12, 15, 17) {real, imag} */,
  {32'h45dd6c1a, 32'h00000000} /* (12, 15, 16) {real, imag} */,
  {32'h45dbaff3, 32'h00000000} /* (12, 15, 15) {real, imag} */,
  {32'h45d45bd8, 32'h00000000} /* (12, 15, 14) {real, imag} */,
  {32'h45bb9245, 32'h00000000} /* (12, 15, 13) {real, imag} */,
  {32'h458f9c6e, 32'h00000000} /* (12, 15, 12) {real, imag} */,
  {32'h44e2b320, 32'h00000000} /* (12, 15, 11) {real, imag} */,
  {32'hc48918ac, 32'h00000000} /* (12, 15, 10) {real, imag} */,
  {32'hc545574a, 32'h00000000} /* (12, 15, 9) {real, imag} */,
  {32'hc5a90571, 32'h00000000} /* (12, 15, 8) {real, imag} */,
  {32'hc5d75055, 32'h00000000} /* (12, 15, 7) {real, imag} */,
  {32'hc6039506, 32'h00000000} /* (12, 15, 6) {real, imag} */,
  {32'hc5f6612b, 32'h00000000} /* (12, 15, 5) {real, imag} */,
  {32'hc6016bef, 32'h00000000} /* (12, 15, 4) {real, imag} */,
  {32'hc60646e6, 32'h00000000} /* (12, 15, 3) {real, imag} */,
  {32'hc600faf6, 32'h00000000} /* (12, 15, 2) {real, imag} */,
  {32'hc60a7d34, 32'h00000000} /* (12, 15, 1) {real, imag} */,
  {32'hc6127a7d, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'hc5fa3548, 32'h00000000} /* (12, 14, 31) {real, imag} */,
  {32'hc600f9bc, 32'h00000000} /* (12, 14, 30) {real, imag} */,
  {32'hc5fcdc8d, 32'h00000000} /* (12, 14, 29) {real, imag} */,
  {32'hc604c331, 32'h00000000} /* (12, 14, 28) {real, imag} */,
  {32'hc609cc20, 32'h00000000} /* (12, 14, 27) {real, imag} */,
  {32'hc5fb9143, 32'h00000000} /* (12, 14, 26) {real, imag} */,
  {32'hc5d65b3e, 32'h00000000} /* (12, 14, 25) {real, imag} */,
  {32'hc5c2ad16, 32'h00000000} /* (12, 14, 24) {real, imag} */,
  {32'hc5a661cd, 32'h00000000} /* (12, 14, 23) {real, imag} */,
  {32'hc54e42aa, 32'h00000000} /* (12, 14, 22) {real, imag} */,
  {32'hc48ec52a, 32'h00000000} /* (12, 14, 21) {real, imag} */,
  {32'h4529399b, 32'h00000000} /* (12, 14, 20) {real, imag} */,
  {32'h457f5866, 32'h00000000} /* (12, 14, 19) {real, imag} */,
  {32'h45b41806, 32'h00000000} /* (12, 14, 18) {real, imag} */,
  {32'h45d86cae, 32'h00000000} /* (12, 14, 17) {real, imag} */,
  {32'h45d68426, 32'h00000000} /* (12, 14, 16) {real, imag} */,
  {32'h45ed6b72, 32'h00000000} /* (12, 14, 15) {real, imag} */,
  {32'h45d08a2d, 32'h00000000} /* (12, 14, 14) {real, imag} */,
  {32'h45a6e9b7, 32'h00000000} /* (12, 14, 13) {real, imag} */,
  {32'h4583c7e6, 32'h00000000} /* (12, 14, 12) {real, imag} */,
  {32'h452d18ae, 32'h00000000} /* (12, 14, 11) {real, imag} */,
  {32'hc3799620, 32'h00000000} /* (12, 14, 10) {real, imag} */,
  {32'hc54234dc, 32'h00000000} /* (12, 14, 9) {real, imag} */,
  {32'hc5a2d0de, 32'h00000000} /* (12, 14, 8) {real, imag} */,
  {32'hc6000307, 32'h00000000} /* (12, 14, 7) {real, imag} */,
  {32'hc6029f06, 32'h00000000} /* (12, 14, 6) {real, imag} */,
  {32'hc5e17794, 32'h00000000} /* (12, 14, 5) {real, imag} */,
  {32'hc5e9a060, 32'h00000000} /* (12, 14, 4) {real, imag} */,
  {32'hc5e73fdd, 32'h00000000} /* (12, 14, 3) {real, imag} */,
  {32'hc5f42f50, 32'h00000000} /* (12, 14, 2) {real, imag} */,
  {32'hc613b8c9, 32'h00000000} /* (12, 14, 1) {real, imag} */,
  {32'hc60bc362, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'hc5d39d36, 32'h00000000} /* (12, 13, 31) {real, imag} */,
  {32'hc5ffa745, 32'h00000000} /* (12, 13, 30) {real, imag} */,
  {32'hc5ebb2de, 32'h00000000} /* (12, 13, 29) {real, imag} */,
  {32'hc5ef819d, 32'h00000000} /* (12, 13, 28) {real, imag} */,
  {32'hc5d0bc14, 32'h00000000} /* (12, 13, 27) {real, imag} */,
  {32'hc5a17c2e, 32'h00000000} /* (12, 13, 26) {real, imag} */,
  {32'hc5adedfe, 32'h00000000} /* (12, 13, 25) {real, imag} */,
  {32'hc5b620d3, 32'h00000000} /* (12, 13, 24) {real, imag} */,
  {32'hc58d3a32, 32'h00000000} /* (12, 13, 23) {real, imag} */,
  {32'hc572341b, 32'h00000000} /* (12, 13, 22) {real, imag} */,
  {32'hc4222318, 32'h00000000} /* (12, 13, 21) {real, imag} */,
  {32'h451e5e5e, 32'h00000000} /* (12, 13, 20) {real, imag} */,
  {32'h4580be58, 32'h00000000} /* (12, 13, 19) {real, imag} */,
  {32'h45c28762, 32'h00000000} /* (12, 13, 18) {real, imag} */,
  {32'h45c48a57, 32'h00000000} /* (12, 13, 17) {real, imag} */,
  {32'h45bec772, 32'h00000000} /* (12, 13, 16) {real, imag} */,
  {32'h45be6ed0, 32'h00000000} /* (12, 13, 15) {real, imag} */,
  {32'h45ce3c6d, 32'h00000000} /* (12, 13, 14) {real, imag} */,
  {32'h4592744e, 32'h00000000} /* (12, 13, 13) {real, imag} */,
  {32'h4568cc82, 32'h00000000} /* (12, 13, 12) {real, imag} */,
  {32'h451ec449, 32'h00000000} /* (12, 13, 11) {real, imag} */,
  {32'hc4530c10, 32'h00000000} /* (12, 13, 10) {real, imag} */,
  {32'hc53d0750, 32'h00000000} /* (12, 13, 9) {real, imag} */,
  {32'hc5871985, 32'h00000000} /* (12, 13, 8) {real, imag} */,
  {32'hc5c5981e, 32'h00000000} /* (12, 13, 7) {real, imag} */,
  {32'hc5bbfc1c, 32'h00000000} /* (12, 13, 6) {real, imag} */,
  {32'hc5c1ff0c, 32'h00000000} /* (12, 13, 5) {real, imag} */,
  {32'hc5da6707, 32'h00000000} /* (12, 13, 4) {real, imag} */,
  {32'hc5ca5066, 32'h00000000} /* (12, 13, 3) {real, imag} */,
  {32'hc5ebea94, 32'h00000000} /* (12, 13, 2) {real, imag} */,
  {32'hc5f367f7, 32'h00000000} /* (12, 13, 1) {real, imag} */,
  {32'hc5d5a98a, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'hc5ab0d9c, 32'h00000000} /* (12, 12, 31) {real, imag} */,
  {32'hc5b58336, 32'h00000000} /* (12, 12, 30) {real, imag} */,
  {32'hc5aa2b6f, 32'h00000000} /* (12, 12, 29) {real, imag} */,
  {32'hc5ac16e1, 32'h00000000} /* (12, 12, 28) {real, imag} */,
  {32'hc5959129, 32'h00000000} /* (12, 12, 27) {real, imag} */,
  {32'hc55e66cc, 32'h00000000} /* (12, 12, 26) {real, imag} */,
  {32'hc56a69b1, 32'h00000000} /* (12, 12, 25) {real, imag} */,
  {32'hc58506f2, 32'h00000000} /* (12, 12, 24) {real, imag} */,
  {32'hc530d0d9, 32'h00000000} /* (12, 12, 23) {real, imag} */,
  {32'hc4be77da, 32'h00000000} /* (12, 12, 22) {real, imag} */,
  {32'hc25aeb00, 32'h00000000} /* (12, 12, 21) {real, imag} */,
  {32'h450d1674, 32'h00000000} /* (12, 12, 20) {real, imag} */,
  {32'h457da0ba, 32'h00000000} /* (12, 12, 19) {real, imag} */,
  {32'h45acdefa, 32'h00000000} /* (12, 12, 18) {real, imag} */,
  {32'h45b7aa63, 32'h00000000} /* (12, 12, 17) {real, imag} */,
  {32'h45be33e0, 32'h00000000} /* (12, 12, 16) {real, imag} */,
  {32'h459d3bea, 32'h00000000} /* (12, 12, 15) {real, imag} */,
  {32'h4591117e, 32'h00000000} /* (12, 12, 14) {real, imag} */,
  {32'h456f4026, 32'h00000000} /* (12, 12, 13) {real, imag} */,
  {32'h452c8412, 32'h00000000} /* (12, 12, 12) {real, imag} */,
  {32'h44c8016f, 32'h00000000} /* (12, 12, 11) {real, imag} */,
  {32'hc4918cb8, 32'h00000000} /* (12, 12, 10) {real, imag} */,
  {32'hc549f1db, 32'h00000000} /* (12, 12, 9) {real, imag} */,
  {32'hc55f8816, 32'h00000000} /* (12, 12, 8) {real, imag} */,
  {32'hc59325fc, 32'h00000000} /* (12, 12, 7) {real, imag} */,
  {32'hc5bd9100, 32'h00000000} /* (12, 12, 6) {real, imag} */,
  {32'hc5ba5070, 32'h00000000} /* (12, 12, 5) {real, imag} */,
  {32'hc596028b, 32'h00000000} /* (12, 12, 4) {real, imag} */,
  {32'hc5b1b6ff, 32'h00000000} /* (12, 12, 3) {real, imag} */,
  {32'hc5a2789e, 32'h00000000} /* (12, 12, 2) {real, imag} */,
  {32'hc5988c9f, 32'h00000000} /* (12, 12, 1) {real, imag} */,
  {32'hc580445c, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'hc4afb494, 32'h00000000} /* (12, 11, 31) {real, imag} */,
  {32'hc50e961e, 32'h00000000} /* (12, 11, 30) {real, imag} */,
  {32'hc4769728, 32'h00000000} /* (12, 11, 29) {real, imag} */,
  {32'hc4ce5c43, 32'h00000000} /* (12, 11, 28) {real, imag} */,
  {32'hc4b5860f, 32'h00000000} /* (12, 11, 27) {real, imag} */,
  {32'hc46ac4f0, 32'h00000000} /* (12, 11, 26) {real, imag} */,
  {32'hc407a1d8, 32'h00000000} /* (12, 11, 25) {real, imag} */,
  {32'hc4b27bc2, 32'h00000000} /* (12, 11, 24) {real, imag} */,
  {32'hc4b208a0, 32'h00000000} /* (12, 11, 23) {real, imag} */,
  {32'hc2930a60, 32'h00000000} /* (12, 11, 22) {real, imag} */,
  {32'h4481b788, 32'h00000000} /* (12, 11, 21) {real, imag} */,
  {32'h451cbde4, 32'h00000000} /* (12, 11, 20) {real, imag} */,
  {32'h453f42f4, 32'h00000000} /* (12, 11, 19) {real, imag} */,
  {32'h45562ad2, 32'h00000000} /* (12, 11, 18) {real, imag} */,
  {32'h455d970d, 32'h00000000} /* (12, 11, 17) {real, imag} */,
  {32'h453785fd, 32'h00000000} /* (12, 11, 16) {real, imag} */,
  {32'h452e4696, 32'h00000000} /* (12, 11, 15) {real, imag} */,
  {32'h45428eca, 32'h00000000} /* (12, 11, 14) {real, imag} */,
  {32'h452317d4, 32'h00000000} /* (12, 11, 13) {real, imag} */,
  {32'h44acabd5, 32'h00000000} /* (12, 11, 12) {real, imag} */,
  {32'h4483ed19, 32'h00000000} /* (12, 11, 11) {real, imag} */,
  {32'hc491843a, 32'h00000000} /* (12, 11, 10) {real, imag} */,
  {32'hc53cc332, 32'h00000000} /* (12, 11, 9) {real, imag} */,
  {32'hc50f9805, 32'h00000000} /* (12, 11, 8) {real, imag} */,
  {32'hc53130a4, 32'h00000000} /* (12, 11, 7) {real, imag} */,
  {32'hc5525007, 32'h00000000} /* (12, 11, 6) {real, imag} */,
  {32'hc545f7c4, 32'h00000000} /* (12, 11, 5) {real, imag} */,
  {32'hc53635c0, 32'h00000000} /* (12, 11, 4) {real, imag} */,
  {32'hc4f361f9, 32'h00000000} /* (12, 11, 3) {real, imag} */,
  {32'hc50006b2, 32'h00000000} /* (12, 11, 2) {real, imag} */,
  {32'hc51f85b5, 32'h00000000} /* (12, 11, 1) {real, imag} */,
  {32'hc501ce13, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'h44ae7beb, 32'h00000000} /* (12, 10, 31) {real, imag} */,
  {32'h450a5408, 32'h00000000} /* (12, 10, 30) {real, imag} */,
  {32'h450a4f54, 32'h00000000} /* (12, 10, 29) {real, imag} */,
  {32'h45402750, 32'h00000000} /* (12, 10, 28) {real, imag} */,
  {32'h4569c79d, 32'h00000000} /* (12, 10, 27) {real, imag} */,
  {32'h4519cc9c, 32'h00000000} /* (12, 10, 26) {real, imag} */,
  {32'h45271f9a, 32'h00000000} /* (12, 10, 25) {real, imag} */,
  {32'h452b2fe1, 32'h00000000} /* (12, 10, 24) {real, imag} */,
  {32'h44edb083, 32'h00000000} /* (12, 10, 23) {real, imag} */,
  {32'h44e9f960, 32'h00000000} /* (12, 10, 22) {real, imag} */,
  {32'h44c75b6b, 32'h00000000} /* (12, 10, 21) {real, imag} */,
  {32'h447f95e6, 32'h00000000} /* (12, 10, 20) {real, imag} */,
  {32'h448828d6, 32'h00000000} /* (12, 10, 19) {real, imag} */,
  {32'h43d6df0f, 32'h00000000} /* (12, 10, 18) {real, imag} */,
  {32'h446d9268, 32'h00000000} /* (12, 10, 17) {real, imag} */,
  {32'hc2889768, 32'h00000000} /* (12, 10, 16) {real, imag} */,
  {32'hc3ad5ad8, 32'h00000000} /* (12, 10, 15) {real, imag} */,
  {32'h438e8280, 32'h00000000} /* (12, 10, 14) {real, imag} */,
  {32'hc454b511, 32'h00000000} /* (12, 10, 13) {real, imag} */,
  {32'hc34cca90, 32'h00000000} /* (12, 10, 12) {real, imag} */,
  {32'hc4898d5a, 32'h00000000} /* (12, 10, 11) {real, imag} */,
  {32'hc423b33d, 32'h00000000} /* (12, 10, 10) {real, imag} */,
  {32'hc3b7cc4c, 32'h00000000} /* (12, 10, 9) {real, imag} */,
  {32'h43dbb4a0, 32'h00000000} /* (12, 10, 8) {real, imag} */,
  {32'h443b298a, 32'h00000000} /* (12, 10, 7) {real, imag} */,
  {32'h44055161, 32'h00000000} /* (12, 10, 6) {real, imag} */,
  {32'h451a963e, 32'h00000000} /* (12, 10, 5) {real, imag} */,
  {32'h44bc29cf, 32'h00000000} /* (12, 10, 4) {real, imag} */,
  {32'h4479d99c, 32'h00000000} /* (12, 10, 3) {real, imag} */,
  {32'h44a28e09, 32'h00000000} /* (12, 10, 2) {real, imag} */,
  {32'h4503dca1, 32'h00000000} /* (12, 10, 1) {real, imag} */,
  {32'h44f14114, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h458ce497, 32'h00000000} /* (12, 9, 31) {real, imag} */,
  {32'h458f97bf, 32'h00000000} /* (12, 9, 30) {real, imag} */,
  {32'h4598f00e, 32'h00000000} /* (12, 9, 29) {real, imag} */,
  {32'h45c6d007, 32'h00000000} /* (12, 9, 28) {real, imag} */,
  {32'h45bad61a, 32'h00000000} /* (12, 9, 27) {real, imag} */,
  {32'h45bd1333, 32'h00000000} /* (12, 9, 26) {real, imag} */,
  {32'h45babc82, 32'h00000000} /* (12, 9, 25) {real, imag} */,
  {32'h45b9471e, 32'h00000000} /* (12, 9, 24) {real, imag} */,
  {32'h459bb4a7, 32'h00000000} /* (12, 9, 23) {real, imag} */,
  {32'h45811831, 32'h00000000} /* (12, 9, 22) {real, imag} */,
  {32'h4547d238, 32'h00000000} /* (12, 9, 21) {real, imag} */,
  {32'h44b3d9e3, 32'h00000000} /* (12, 9, 20) {real, imag} */,
  {32'hc2897f00, 32'h00000000} /* (12, 9, 19) {real, imag} */,
  {32'hc45fa424, 32'h00000000} /* (12, 9, 18) {real, imag} */,
  {32'hc4d302a4, 32'h00000000} /* (12, 9, 17) {real, imag} */,
  {32'hc51d2e38, 32'h00000000} /* (12, 9, 16) {real, imag} */,
  {32'hc51695b8, 32'h00000000} /* (12, 9, 15) {real, imag} */,
  {32'hc53bdf0c, 32'h00000000} /* (12, 9, 14) {real, imag} */,
  {32'hc5435f3c, 32'h00000000} /* (12, 9, 13) {real, imag} */,
  {32'hc5165e26, 32'h00000000} /* (12, 9, 12) {real, imag} */,
  {32'hc4e0b9f2, 32'h00000000} /* (12, 9, 11) {real, imag} */,
  {32'hc306aa60, 32'h00000000} /* (12, 9, 10) {real, imag} */,
  {32'h44a9c426, 32'h00000000} /* (12, 9, 9) {real, imag} */,
  {32'h452f429d, 32'h00000000} /* (12, 9, 8) {real, imag} */,
  {32'h4527da50, 32'h00000000} /* (12, 9, 7) {real, imag} */,
  {32'h455198a0, 32'h00000000} /* (12, 9, 6) {real, imag} */,
  {32'h4576ebf0, 32'h00000000} /* (12, 9, 5) {real, imag} */,
  {32'h4554ad56, 32'h00000000} /* (12, 9, 4) {real, imag} */,
  {32'h456d8727, 32'h00000000} /* (12, 9, 3) {real, imag} */,
  {32'h456568fd, 32'h00000000} /* (12, 9, 2) {real, imag} */,
  {32'h4591c3b9, 32'h00000000} /* (12, 9, 1) {real, imag} */,
  {32'h456a8328, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'h45c00370, 32'h00000000} /* (12, 8, 31) {real, imag} */,
  {32'h45c727cd, 32'h00000000} /* (12, 8, 30) {real, imag} */,
  {32'h45dc4879, 32'h00000000} /* (12, 8, 29) {real, imag} */,
  {32'h46040637, 32'h00000000} /* (12, 8, 28) {real, imag} */,
  {32'h45f6994e, 32'h00000000} /* (12, 8, 27) {real, imag} */,
  {32'h4607a53e, 32'h00000000} /* (12, 8, 26) {real, imag} */,
  {32'h45e5ca08, 32'h00000000} /* (12, 8, 25) {real, imag} */,
  {32'h46138477, 32'h00000000} /* (12, 8, 24) {real, imag} */,
  {32'h45ea2b4e, 32'h00000000} /* (12, 8, 23) {real, imag} */,
  {32'h45a72a76, 32'h00000000} /* (12, 8, 22) {real, imag} */,
  {32'h459bca42, 32'h00000000} /* (12, 8, 21) {real, imag} */,
  {32'h44a103b4, 32'h00000000} /* (12, 8, 20) {real, imag} */,
  {32'h438afd90, 32'h00000000} /* (12, 8, 19) {real, imag} */,
  {32'hc49c0c9e, 32'h00000000} /* (12, 8, 18) {real, imag} */,
  {32'hc5223b6d, 32'h00000000} /* (12, 8, 17) {real, imag} */,
  {32'hc556ee61, 32'h00000000} /* (12, 8, 16) {real, imag} */,
  {32'hc5a03ff2, 32'h00000000} /* (12, 8, 15) {real, imag} */,
  {32'hc58b14cf, 32'h00000000} /* (12, 8, 14) {real, imag} */,
  {32'hc559c4de, 32'h00000000} /* (12, 8, 13) {real, imag} */,
  {32'hc54cf4db, 32'h00000000} /* (12, 8, 12) {real, imag} */,
  {32'hc5089db0, 32'h00000000} /* (12, 8, 11) {real, imag} */,
  {32'h43323280, 32'h00000000} /* (12, 8, 10) {real, imag} */,
  {32'h44c3253e, 32'h00000000} /* (12, 8, 9) {real, imag} */,
  {32'h452e398c, 32'h00000000} /* (12, 8, 8) {real, imag} */,
  {32'h457cd7c4, 32'h00000000} /* (12, 8, 7) {real, imag} */,
  {32'h458953ec, 32'h00000000} /* (12, 8, 6) {real, imag} */,
  {32'h459f0c8c, 32'h00000000} /* (12, 8, 5) {real, imag} */,
  {32'h45af8fc8, 32'h00000000} /* (12, 8, 4) {real, imag} */,
  {32'h45ab512f, 32'h00000000} /* (12, 8, 3) {real, imag} */,
  {32'h45a51bc4, 32'h00000000} /* (12, 8, 2) {real, imag} */,
  {32'h45b9e114, 32'h00000000} /* (12, 8, 1) {real, imag} */,
  {32'h45b60402, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'h45e3e9d4, 32'h00000000} /* (12, 7, 31) {real, imag} */,
  {32'h46018147, 32'h00000000} /* (12, 7, 30) {real, imag} */,
  {32'h4603c716, 32'h00000000} /* (12, 7, 29) {real, imag} */,
  {32'h460ad02c, 32'h00000000} /* (12, 7, 28) {real, imag} */,
  {32'h46169efa, 32'h00000000} /* (12, 7, 27) {real, imag} */,
  {32'h460e7bb6, 32'h00000000} /* (12, 7, 26) {real, imag} */,
  {32'h460a74e6, 32'h00000000} /* (12, 7, 25) {real, imag} */,
  {32'h46080b2a, 32'h00000000} /* (12, 7, 24) {real, imag} */,
  {32'h45fa7739, 32'h00000000} /* (12, 7, 23) {real, imag} */,
  {32'h45dda19b, 32'h00000000} /* (12, 7, 22) {real, imag} */,
  {32'h45b18889, 32'h00000000} /* (12, 7, 21) {real, imag} */,
  {32'h451046f1, 32'h00000000} /* (12, 7, 20) {real, imag} */,
  {32'hc38fa2b0, 32'h00000000} /* (12, 7, 19) {real, imag} */,
  {32'hc4bf8a80, 32'h00000000} /* (12, 7, 18) {real, imag} */,
  {32'hc50b956c, 32'h00000000} /* (12, 7, 17) {real, imag} */,
  {32'hc573c953, 32'h00000000} /* (12, 7, 16) {real, imag} */,
  {32'hc5b6afee, 32'h00000000} /* (12, 7, 15) {real, imag} */,
  {32'hc59ea8a0, 32'h00000000} /* (12, 7, 14) {real, imag} */,
  {32'hc58f2040, 32'h00000000} /* (12, 7, 13) {real, imag} */,
  {32'hc5aa5ed4, 32'h00000000} /* (12, 7, 12) {real, imag} */,
  {32'hc563d1fa, 32'h00000000} /* (12, 7, 11) {real, imag} */,
  {32'hc3ad24a0, 32'h00000000} /* (12, 7, 10) {real, imag} */,
  {32'h44247d18, 32'h00000000} /* (12, 7, 9) {real, imag} */,
  {32'h455adf47, 32'h00000000} /* (12, 7, 8) {real, imag} */,
  {32'h457b5ab2, 32'h00000000} /* (12, 7, 7) {real, imag} */,
  {32'h459a430d, 32'h00000000} /* (12, 7, 6) {real, imag} */,
  {32'h45b572ab, 32'h00000000} /* (12, 7, 5) {real, imag} */,
  {32'h4604412c, 32'h00000000} /* (12, 7, 4) {real, imag} */,
  {32'h45e86e9f, 32'h00000000} /* (12, 7, 3) {real, imag} */,
  {32'h45ebf5d8, 32'h00000000} /* (12, 7, 2) {real, imag} */,
  {32'h45f6294c, 32'h00000000} /* (12, 7, 1) {real, imag} */,
  {32'h45de3432, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'h4603c949, 32'h00000000} /* (12, 6, 31) {real, imag} */,
  {32'h46085232, 32'h00000000} /* (12, 6, 30) {real, imag} */,
  {32'h4613ba43, 32'h00000000} /* (12, 6, 29) {real, imag} */,
  {32'h461e72a6, 32'h00000000} /* (12, 6, 28) {real, imag} */,
  {32'h46227560, 32'h00000000} /* (12, 6, 27) {real, imag} */,
  {32'h46293797, 32'h00000000} /* (12, 6, 26) {real, imag} */,
  {32'h4625284d, 32'h00000000} /* (12, 6, 25) {real, imag} */,
  {32'h4616a9a2, 32'h00000000} /* (12, 6, 24) {real, imag} */,
  {32'h460c5323, 32'h00000000} /* (12, 6, 23) {real, imag} */,
  {32'h4604fb35, 32'h00000000} /* (12, 6, 22) {real, imag} */,
  {32'h45d9aa50, 32'h00000000} /* (12, 6, 21) {real, imag} */,
  {32'h4576f55e, 32'h00000000} /* (12, 6, 20) {real, imag} */,
  {32'h44c76fe4, 32'h00000000} /* (12, 6, 19) {real, imag} */,
  {32'hc3d24620, 32'h00000000} /* (12, 6, 18) {real, imag} */,
  {32'hc4e38d40, 32'h00000000} /* (12, 6, 17) {real, imag} */,
  {32'hc58c8f2e, 32'h00000000} /* (12, 6, 16) {real, imag} */,
  {32'hc56df763, 32'h00000000} /* (12, 6, 15) {real, imag} */,
  {32'hc5bc4400, 32'h00000000} /* (12, 6, 14) {real, imag} */,
  {32'hc5b8bb76, 32'h00000000} /* (12, 6, 13) {real, imag} */,
  {32'hc5a1c5eb, 32'h00000000} /* (12, 6, 12) {real, imag} */,
  {32'hc586bff0, 32'h00000000} /* (12, 6, 11) {real, imag} */,
  {32'hc5262f4b, 32'h00000000} /* (12, 6, 10) {real, imag} */,
  {32'hc38aac00, 32'h00000000} /* (12, 6, 9) {real, imag} */,
  {32'h45271ea7, 32'h00000000} /* (12, 6, 8) {real, imag} */,
  {32'h45612cc4, 32'h00000000} /* (12, 6, 7) {real, imag} */,
  {32'h458b79f6, 32'h00000000} /* (12, 6, 6) {real, imag} */,
  {32'h45c2cf08, 32'h00000000} /* (12, 6, 5) {real, imag} */,
  {32'h45e4d049, 32'h00000000} /* (12, 6, 4) {real, imag} */,
  {32'h4607649a, 32'h00000000} /* (12, 6, 3) {real, imag} */,
  {32'h461382ed, 32'h00000000} /* (12, 6, 2) {real, imag} */,
  {32'h460e1db3, 32'h00000000} /* (12, 6, 1) {real, imag} */,
  {32'h46003d86, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'h461306dc, 32'h00000000} /* (12, 5, 31) {real, imag} */,
  {32'h461d8a14, 32'h00000000} /* (12, 5, 30) {real, imag} */,
  {32'h46323366, 32'h00000000} /* (12, 5, 29) {real, imag} */,
  {32'h463aaf54, 32'h00000000} /* (12, 5, 28) {real, imag} */,
  {32'h4638cad6, 32'h00000000} /* (12, 5, 27) {real, imag} */,
  {32'h46359814, 32'h00000000} /* (12, 5, 26) {real, imag} */,
  {32'h46304099, 32'h00000000} /* (12, 5, 25) {real, imag} */,
  {32'h462a1db0, 32'h00000000} /* (12, 5, 24) {real, imag} */,
  {32'h462dc22e, 32'h00000000} /* (12, 5, 23) {real, imag} */,
  {32'h460a73ae, 32'h00000000} /* (12, 5, 22) {real, imag} */,
  {32'h45f886f7, 32'h00000000} /* (12, 5, 21) {real, imag} */,
  {32'h45c1126b, 32'h00000000} /* (12, 5, 20) {real, imag} */,
  {32'h45734015, 32'h00000000} /* (12, 5, 19) {real, imag} */,
  {32'h453470c0, 32'h00000000} /* (12, 5, 18) {real, imag} */,
  {32'h44ad4314, 32'h00000000} /* (12, 5, 17) {real, imag} */,
  {32'hc4c5d522, 32'h00000000} /* (12, 5, 16) {real, imag} */,
  {32'hc585bd21, 32'h00000000} /* (12, 5, 15) {real, imag} */,
  {32'hc5998e13, 32'h00000000} /* (12, 5, 14) {real, imag} */,
  {32'hc5a9ffdb, 32'h00000000} /* (12, 5, 13) {real, imag} */,
  {32'hc5b40734, 32'h00000000} /* (12, 5, 12) {real, imag} */,
  {32'hc5b168b3, 32'h00000000} /* (12, 5, 11) {real, imag} */,
  {32'hc558e02a, 32'h00000000} /* (12, 5, 10) {real, imag} */,
  {32'hc4fa2aa0, 32'h00000000} /* (12, 5, 9) {real, imag} */,
  {32'hc2b223c0, 32'h00000000} /* (12, 5, 8) {real, imag} */,
  {32'h44861b50, 32'h00000000} /* (12, 5, 7) {real, imag} */,
  {32'h4543fb0e, 32'h00000000} /* (12, 5, 6) {real, imag} */,
  {32'h45a7767f, 32'h00000000} /* (12, 5, 5) {real, imag} */,
  {32'h45dd145d, 32'h00000000} /* (12, 5, 4) {real, imag} */,
  {32'h460eacbe, 32'h00000000} /* (12, 5, 3) {real, imag} */,
  {32'h46177257, 32'h00000000} /* (12, 5, 2) {real, imag} */,
  {32'h4617a288, 32'h00000000} /* (12, 5, 1) {real, imag} */,
  {32'h4611c17a, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'h461eca52, 32'h00000000} /* (12, 4, 31) {real, imag} */,
  {32'h463ab5a9, 32'h00000000} /* (12, 4, 30) {real, imag} */,
  {32'h463bdd66, 32'h00000000} /* (12, 4, 29) {real, imag} */,
  {32'h4637657a, 32'h00000000} /* (12, 4, 28) {real, imag} */,
  {32'h464bdb25, 32'h00000000} /* (12, 4, 27) {real, imag} */,
  {32'h4641f71a, 32'h00000000} /* (12, 4, 26) {real, imag} */,
  {32'h4639da04, 32'h00000000} /* (12, 4, 25) {real, imag} */,
  {32'h462a1c75, 32'h00000000} /* (12, 4, 24) {real, imag} */,
  {32'h46301806, 32'h00000000} /* (12, 4, 23) {real, imag} */,
  {32'h46207d0d, 32'h00000000} /* (12, 4, 22) {real, imag} */,
  {32'h461b8d50, 32'h00000000} /* (12, 4, 21) {real, imag} */,
  {32'h45fd886e, 32'h00000000} /* (12, 4, 20) {real, imag} */,
  {32'h45b33626, 32'h00000000} /* (12, 4, 19) {real, imag} */,
  {32'h45a2c598, 32'h00000000} /* (12, 4, 18) {real, imag} */,
  {32'h4527ba36, 32'h00000000} /* (12, 4, 17) {real, imag} */,
  {32'hc3106400, 32'h00000000} /* (12, 4, 16) {real, imag} */,
  {32'hc5516e68, 32'h00000000} /* (12, 4, 15) {real, imag} */,
  {32'hc5a188d2, 32'h00000000} /* (12, 4, 14) {real, imag} */,
  {32'hc5b71d1c, 32'h00000000} /* (12, 4, 13) {real, imag} */,
  {32'hc5c03dc0, 32'h00000000} /* (12, 4, 12) {real, imag} */,
  {32'hc5b16986, 32'h00000000} /* (12, 4, 11) {real, imag} */,
  {32'hc5a56afb, 32'h00000000} /* (12, 4, 10) {real, imag} */,
  {32'hc5642b28, 32'h00000000} /* (12, 4, 9) {real, imag} */,
  {32'hc50233f4, 32'h00000000} /* (12, 4, 8) {real, imag} */,
  {32'hc3db2c10, 32'h00000000} /* (12, 4, 7) {real, imag} */,
  {32'h44c5c0c8, 32'h00000000} /* (12, 4, 6) {real, imag} */,
  {32'h4581e010, 32'h00000000} /* (12, 4, 5) {real, imag} */,
  {32'h45e694f2, 32'h00000000} /* (12, 4, 4) {real, imag} */,
  {32'h4606367d, 32'h00000000} /* (12, 4, 3) {real, imag} */,
  {32'h461ab00d, 32'h00000000} /* (12, 4, 2) {real, imag} */,
  {32'h46201c78, 32'h00000000} /* (12, 4, 1) {real, imag} */,
  {32'h46181e82, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'h4626ccb5, 32'h00000000} /* (12, 3, 31) {real, imag} */,
  {32'h463c948e, 32'h00000000} /* (12, 3, 30) {real, imag} */,
  {32'h464fd232, 32'h00000000} /* (12, 3, 29) {real, imag} */,
  {32'h463e0466, 32'h00000000} /* (12, 3, 28) {real, imag} */,
  {32'h463c9510, 32'h00000000} /* (12, 3, 27) {real, imag} */,
  {32'h4638fbd9, 32'h00000000} /* (12, 3, 26) {real, imag} */,
  {32'h463fa024, 32'h00000000} /* (12, 3, 25) {real, imag} */,
  {32'h463ab39a, 32'h00000000} /* (12, 3, 24) {real, imag} */,
  {32'h4637cbe5, 32'h00000000} /* (12, 3, 23) {real, imag} */,
  {32'h4635889c, 32'h00000000} /* (12, 3, 22) {real, imag} */,
  {32'h4614aebc, 32'h00000000} /* (12, 3, 21) {real, imag} */,
  {32'h45fba591, 32'h00000000} /* (12, 3, 20) {real, imag} */,
  {32'h45c8bfce, 32'h00000000} /* (12, 3, 19) {real, imag} */,
  {32'h459b855a, 32'h00000000} /* (12, 3, 18) {real, imag} */,
  {32'h453950cc, 32'h00000000} /* (12, 3, 17) {real, imag} */,
  {32'h43bfb170, 32'h00000000} /* (12, 3, 16) {real, imag} */,
  {32'hc54e06b8, 32'h00000000} /* (12, 3, 15) {real, imag} */,
  {32'hc59e40bc, 32'h00000000} /* (12, 3, 14) {real, imag} */,
  {32'hc59c5815, 32'h00000000} /* (12, 3, 13) {real, imag} */,
  {32'hc5badf71, 32'h00000000} /* (12, 3, 12) {real, imag} */,
  {32'hc5b80de5, 32'h00000000} /* (12, 3, 11) {real, imag} */,
  {32'hc5aa188a, 32'h00000000} /* (12, 3, 10) {real, imag} */,
  {32'hc588fcf5, 32'h00000000} /* (12, 3, 9) {real, imag} */,
  {32'hc54cc096, 32'h00000000} /* (12, 3, 8) {real, imag} */,
  {32'hc49d7a70, 32'h00000000} /* (12, 3, 7) {real, imag} */,
  {32'hc377da80, 32'h00000000} /* (12, 3, 6) {real, imag} */,
  {32'h459af126, 32'h00000000} /* (12, 3, 5) {real, imag} */,
  {32'h45f953ad, 32'h00000000} /* (12, 3, 4) {real, imag} */,
  {32'h45f9d3e4, 32'h00000000} /* (12, 3, 3) {real, imag} */,
  {32'h46199819, 32'h00000000} /* (12, 3, 2) {real, imag} */,
  {32'h461be9ea, 32'h00000000} /* (12, 3, 1) {real, imag} */,
  {32'h4618a858, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'h462e62c2, 32'h00000000} /* (12, 2, 31) {real, imag} */,
  {32'h463baa1e, 32'h00000000} /* (12, 2, 30) {real, imag} */,
  {32'h463ff43a, 32'h00000000} /* (12, 2, 29) {real, imag} */,
  {32'h464acce0, 32'h00000000} /* (12, 2, 28) {real, imag} */,
  {32'h464507fc, 32'h00000000} /* (12, 2, 27) {real, imag} */,
  {32'h463d9fb0, 32'h00000000} /* (12, 2, 26) {real, imag} */,
  {32'h46570121, 32'h00000000} /* (12, 2, 25) {real, imag} */,
  {32'h464a4225, 32'h00000000} /* (12, 2, 24) {real, imag} */,
  {32'h463f91a0, 32'h00000000} /* (12, 2, 23) {real, imag} */,
  {32'h461df6c9, 32'h00000000} /* (12, 2, 22) {real, imag} */,
  {32'h45f57aec, 32'h00000000} /* (12, 2, 21) {real, imag} */,
  {32'h460333f7, 32'h00000000} /* (12, 2, 20) {real, imag} */,
  {32'h45ccb7d8, 32'h00000000} /* (12, 2, 19) {real, imag} */,
  {32'h45a3c362, 32'h00000000} /* (12, 2, 18) {real, imag} */,
  {32'h450ccf6c, 32'h00000000} /* (12, 2, 17) {real, imag} */,
  {32'h442c0fb0, 32'h00000000} /* (12, 2, 16) {real, imag} */,
  {32'hc5127616, 32'h00000000} /* (12, 2, 15) {real, imag} */,
  {32'hc58b1098, 32'h00000000} /* (12, 2, 14) {real, imag} */,
  {32'hc5ca28c4, 32'h00000000} /* (12, 2, 13) {real, imag} */,
  {32'hc5cf90a7, 32'h00000000} /* (12, 2, 12) {real, imag} */,
  {32'hc5afa59f, 32'h00000000} /* (12, 2, 11) {real, imag} */,
  {32'hc59e06b7, 32'h00000000} /* (12, 2, 10) {real, imag} */,
  {32'hc5747a34, 32'h00000000} /* (12, 2, 9) {real, imag} */,
  {32'hc55a6da4, 32'h00000000} /* (12, 2, 8) {real, imag} */,
  {32'hc4ad0750, 32'h00000000} /* (12, 2, 7) {real, imag} */,
  {32'h44203850, 32'h00000000} /* (12, 2, 6) {real, imag} */,
  {32'h458917b8, 32'h00000000} /* (12, 2, 5) {real, imag} */,
  {32'h460538f5, 32'h00000000} /* (12, 2, 4) {real, imag} */,
  {32'h46062ed1, 32'h00000000} /* (12, 2, 3) {real, imag} */,
  {32'h4619fdb2, 32'h00000000} /* (12, 2, 2) {real, imag} */,
  {32'h462869cb, 32'h00000000} /* (12, 2, 1) {real, imag} */,
  {32'h462102a9, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'h4630f56e, 32'h00000000} /* (12, 1, 31) {real, imag} */,
  {32'h463a4544, 32'h00000000} /* (12, 1, 30) {real, imag} */,
  {32'h4636f69a, 32'h00000000} /* (12, 1, 29) {real, imag} */,
  {32'h463b6a0c, 32'h00000000} /* (12, 1, 28) {real, imag} */,
  {32'h4648d02a, 32'h00000000} /* (12, 1, 27) {real, imag} */,
  {32'h46408714, 32'h00000000} /* (12, 1, 26) {real, imag} */,
  {32'h4641d8cc, 32'h00000000} /* (12, 1, 25) {real, imag} */,
  {32'h46426414, 32'h00000000} /* (12, 1, 24) {real, imag} */,
  {32'h46317212, 32'h00000000} /* (12, 1, 23) {real, imag} */,
  {32'h460b66f9, 32'h00000000} /* (12, 1, 22) {real, imag} */,
  {32'h4602a6b7, 32'h00000000} /* (12, 1, 21) {real, imag} */,
  {32'h45f1ac03, 32'h00000000} /* (12, 1, 20) {real, imag} */,
  {32'h45abe6d2, 32'h00000000} /* (12, 1, 19) {real, imag} */,
  {32'h45979c4c, 32'h00000000} /* (12, 1, 18) {real, imag} */,
  {32'h45013600, 32'h00000000} /* (12, 1, 17) {real, imag} */,
  {32'h41a93e00, 32'h00000000} /* (12, 1, 16) {real, imag} */,
  {32'hc5610b38, 32'h00000000} /* (12, 1, 15) {real, imag} */,
  {32'hc5c08430, 32'h00000000} /* (12, 1, 14) {real, imag} */,
  {32'hc5c1cf5d, 32'h00000000} /* (12, 1, 13) {real, imag} */,
  {32'hc5b85dcd, 32'h00000000} /* (12, 1, 12) {real, imag} */,
  {32'hc58adb9d, 32'h00000000} /* (12, 1, 11) {real, imag} */,
  {32'hc5893169, 32'h00000000} /* (12, 1, 10) {real, imag} */,
  {32'hc54f9ab2, 32'h00000000} /* (12, 1, 9) {real, imag} */,
  {32'hc52c94ae, 32'h00000000} /* (12, 1, 8) {real, imag} */,
  {32'hc49c9dc0, 32'h00000000} /* (12, 1, 7) {real, imag} */,
  {32'h44969a28, 32'h00000000} /* (12, 1, 6) {real, imag} */,
  {32'h4584524c, 32'h00000000} /* (12, 1, 5) {real, imag} */,
  {32'h45f1fdc3, 32'h00000000} /* (12, 1, 4) {real, imag} */,
  {32'h46099566, 32'h00000000} /* (12, 1, 3) {real, imag} */,
  {32'h461456d5, 32'h00000000} /* (12, 1, 2) {real, imag} */,
  {32'h462c17a5, 32'h00000000} /* (12, 1, 1) {real, imag} */,
  {32'h4629aa9d, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'h46237b7b, 32'h00000000} /* (12, 0, 31) {real, imag} */,
  {32'h4631a44a, 32'h00000000} /* (12, 0, 30) {real, imag} */,
  {32'h463281a4, 32'h00000000} /* (12, 0, 29) {real, imag} */,
  {32'h463a2521, 32'h00000000} /* (12, 0, 28) {real, imag} */,
  {32'h463a2f5c, 32'h00000000} /* (12, 0, 27) {real, imag} */,
  {32'h463c46d0, 32'h00000000} /* (12, 0, 26) {real, imag} */,
  {32'h4632142e, 32'h00000000} /* (12, 0, 25) {real, imag} */,
  {32'h462c9b29, 32'h00000000} /* (12, 0, 24) {real, imag} */,
  {32'h462a135b, 32'h00000000} /* (12, 0, 23) {real, imag} */,
  {32'h46083a50, 32'h00000000} /* (12, 0, 22) {real, imag} */,
  {32'h45e56c2e, 32'h00000000} /* (12, 0, 21) {real, imag} */,
  {32'h45b07a05, 32'h00000000} /* (12, 0, 20) {real, imag} */,
  {32'h457e91d6, 32'h00000000} /* (12, 0, 19) {real, imag} */,
  {32'h4506aa68, 32'h00000000} /* (12, 0, 18) {real, imag} */,
  {32'h43a66020, 32'h00000000} /* (12, 0, 17) {real, imag} */,
  {32'hc4d0e5b0, 32'h00000000} /* (12, 0, 16) {real, imag} */,
  {32'hc57a3bd5, 32'h00000000} /* (12, 0, 15) {real, imag} */,
  {32'hc5b5b4ac, 32'h00000000} /* (12, 0, 14) {real, imag} */,
  {32'hc59d850f, 32'h00000000} /* (12, 0, 13) {real, imag} */,
  {32'hc5982f4a, 32'h00000000} /* (12, 0, 12) {real, imag} */,
  {32'hc578ecda, 32'h00000000} /* (12, 0, 11) {real, imag} */,
  {32'hc5402b46, 32'h00000000} /* (12, 0, 10) {real, imag} */,
  {32'hc4c71d6c, 32'h00000000} /* (12, 0, 9) {real, imag} */,
  {32'hc3401c40, 32'h00000000} /* (12, 0, 8) {real, imag} */,
  {32'h44910258, 32'h00000000} /* (12, 0, 7) {real, imag} */,
  {32'h4539a2b9, 32'h00000000} /* (12, 0, 6) {real, imag} */,
  {32'h45b1a484, 32'h00000000} /* (12, 0, 5) {real, imag} */,
  {32'h45ecc8b3, 32'h00000000} /* (12, 0, 4) {real, imag} */,
  {32'h46101236, 32'h00000000} /* (12, 0, 3) {real, imag} */,
  {32'h460ddd5a, 32'h00000000} /* (12, 0, 2) {real, imag} */,
  {32'h46143e0c, 32'h00000000} /* (12, 0, 1) {real, imag} */,
  {32'h4620edb2, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h46358279, 32'h00000000} /* (11, 31, 31) {real, imag} */,
  {32'h4643b177, 32'h00000000} /* (11, 31, 30) {real, imag} */,
  {32'h4649b95c, 32'h00000000} /* (11, 31, 29) {real, imag} */,
  {32'h46474ab5, 32'h00000000} /* (11, 31, 28) {real, imag} */,
  {32'h4651b511, 32'h00000000} /* (11, 31, 27) {real, imag} */,
  {32'h4650b51a, 32'h00000000} /* (11, 31, 26) {real, imag} */,
  {32'h46433809, 32'h00000000} /* (11, 31, 25) {real, imag} */,
  {32'h4638069c, 32'h00000000} /* (11, 31, 24) {real, imag} */,
  {32'h46289f9b, 32'h00000000} /* (11, 31, 23) {real, imag} */,
  {32'h460d7300, 32'h00000000} /* (11, 31, 22) {real, imag} */,
  {32'h45cf0ce7, 32'h00000000} /* (11, 31, 21) {real, imag} */,
  {32'h455b927b, 32'h00000000} /* (11, 31, 20) {real, imag} */,
  {32'h44b9ed44, 32'h00000000} /* (11, 31, 19) {real, imag} */,
  {32'hc3954410, 32'h00000000} /* (11, 31, 18) {real, imag} */,
  {32'hc506f9c4, 32'h00000000} /* (11, 31, 17) {real, imag} */,
  {32'hc58b30d1, 32'h00000000} /* (11, 31, 16) {real, imag} */,
  {32'hc5b3f612, 32'h00000000} /* (11, 31, 15) {real, imag} */,
  {32'hc5b0695e, 32'h00000000} /* (11, 31, 14) {real, imag} */,
  {32'hc5c89d88, 32'h00000000} /* (11, 31, 13) {real, imag} */,
  {32'hc5a613b6, 32'h00000000} /* (11, 31, 12) {real, imag} */,
  {32'hc597aede, 32'h00000000} /* (11, 31, 11) {real, imag} */,
  {32'hc430a578, 32'h00000000} /* (11, 31, 10) {real, imag} */,
  {32'h444ba930, 32'h00000000} /* (11, 31, 9) {real, imag} */,
  {32'h45210bfc, 32'h00000000} /* (11, 31, 8) {real, imag} */,
  {32'h4582a45e, 32'h00000000} /* (11, 31, 7) {real, imag} */,
  {32'h45c06c60, 32'h00000000} /* (11, 31, 6) {real, imag} */,
  {32'h45fd7491, 32'h00000000} /* (11, 31, 5) {real, imag} */,
  {32'h46173a19, 32'h00000000} /* (11, 31, 4) {real, imag} */,
  {32'h46258844, 32'h00000000} /* (11, 31, 3) {real, imag} */,
  {32'h46395eee, 32'h00000000} /* (11, 31, 2) {real, imag} */,
  {32'h462b3581, 32'h00000000} /* (11, 31, 1) {real, imag} */,
  {32'h464154bc, 32'h00000000} /* (11, 31, 0) {real, imag} */,
  {32'h4645cebd, 32'h00000000} /* (11, 30, 31) {real, imag} */,
  {32'h46419ad6, 32'h00000000} /* (11, 30, 30) {real, imag} */,
  {32'h4642da7c, 32'h00000000} /* (11, 30, 29) {real, imag} */,
  {32'h464c760c, 32'h00000000} /* (11, 30, 28) {real, imag} */,
  {32'h464d871d, 32'h00000000} /* (11, 30, 27) {real, imag} */,
  {32'h46518eac, 32'h00000000} /* (11, 30, 26) {real, imag} */,
  {32'h464c65e6, 32'h00000000} /* (11, 30, 25) {real, imag} */,
  {32'h4645b416, 32'h00000000} /* (11, 30, 24) {real, imag} */,
  {32'h46263051, 32'h00000000} /* (11, 30, 23) {real, imag} */,
  {32'h45f68bde, 32'h00000000} /* (11, 30, 22) {real, imag} */,
  {32'h45afba34, 32'h00000000} /* (11, 30, 21) {real, imag} */,
  {32'h451d13d2, 32'h00000000} /* (11, 30, 20) {real, imag} */,
  {32'hc2d39a00, 32'h00000000} /* (11, 30, 19) {real, imag} */,
  {32'hc519313e, 32'h00000000} /* (11, 30, 18) {real, imag} */,
  {32'hc599f9fa, 32'h00000000} /* (11, 30, 17) {real, imag} */,
  {32'hc5adbd31, 32'h00000000} /* (11, 30, 16) {real, imag} */,
  {32'hc5d1b16a, 32'h00000000} /* (11, 30, 15) {real, imag} */,
  {32'hc5e96020, 32'h00000000} /* (11, 30, 14) {real, imag} */,
  {32'hc5c94ca1, 32'h00000000} /* (11, 30, 13) {real, imag} */,
  {32'hc5a8255d, 32'h00000000} /* (11, 30, 12) {real, imag} */,
  {32'hc5472694, 32'h00000000} /* (11, 30, 11) {real, imag} */,
  {32'h44a4b204, 32'h00000000} /* (11, 30, 10) {real, imag} */,
  {32'h453bf2ce, 32'h00000000} /* (11, 30, 9) {real, imag} */,
  {32'h457ebbaa, 32'h00000000} /* (11, 30, 8) {real, imag} */,
  {32'h45cdbefe, 32'h00000000} /* (11, 30, 7) {real, imag} */,
  {32'h460300ab, 32'h00000000} /* (11, 30, 6) {real, imag} */,
  {32'h46215761, 32'h00000000} /* (11, 30, 5) {real, imag} */,
  {32'h463b1c80, 32'h00000000} /* (11, 30, 4) {real, imag} */,
  {32'h463591b0, 32'h00000000} /* (11, 30, 3) {real, imag} */,
  {32'h46416a72, 32'h00000000} /* (11, 30, 2) {real, imag} */,
  {32'h4632f2e1, 32'h00000000} /* (11, 30, 1) {real, imag} */,
  {32'h46388d16, 32'h00000000} /* (11, 30, 0) {real, imag} */,
  {32'h464821f7, 32'h00000000} /* (11, 29, 31) {real, imag} */,
  {32'h4652ed56, 32'h00000000} /* (11, 29, 30) {real, imag} */,
  {32'h4651b4d0, 32'h00000000} /* (11, 29, 29) {real, imag} */,
  {32'h4652d8be, 32'h00000000} /* (11, 29, 28) {real, imag} */,
  {32'h4643b536, 32'h00000000} /* (11, 29, 27) {real, imag} */,
  {32'h464958ac, 32'h00000000} /* (11, 29, 26) {real, imag} */,
  {32'h4642e181, 32'h00000000} /* (11, 29, 25) {real, imag} */,
  {32'h4638b9c9, 32'h00000000} /* (11, 29, 24) {real, imag} */,
  {32'h4623f76a, 32'h00000000} /* (11, 29, 23) {real, imag} */,
  {32'h45fa4c10, 32'h00000000} /* (11, 29, 22) {real, imag} */,
  {32'h458f898a, 32'h00000000} /* (11, 29, 21) {real, imag} */,
  {32'h44afe108, 32'h00000000} /* (11, 29, 20) {real, imag} */,
  {32'hc4d3ede0, 32'h00000000} /* (11, 29, 19) {real, imag} */,
  {32'hc5848048, 32'h00000000} /* (11, 29, 18) {real, imag} */,
  {32'hc5aa8fde, 32'h00000000} /* (11, 29, 17) {real, imag} */,
  {32'hc5bda4f6, 32'h00000000} /* (11, 29, 16) {real, imag} */,
  {32'hc5df6ec2, 32'h00000000} /* (11, 29, 15) {real, imag} */,
  {32'hc5e84aab, 32'h00000000} /* (11, 29, 14) {real, imag} */,
  {32'hc5cfd38d, 32'h00000000} /* (11, 29, 13) {real, imag} */,
  {32'hc5ab09bc, 32'h00000000} /* (11, 29, 12) {real, imag} */,
  {32'hc504e8b0, 32'h00000000} /* (11, 29, 11) {real, imag} */,
  {32'h44aa9dcc, 32'h00000000} /* (11, 29, 10) {real, imag} */,
  {32'h456f47e4, 32'h00000000} /* (11, 29, 9) {real, imag} */,
  {32'h45b8620a, 32'h00000000} /* (11, 29, 8) {real, imag} */,
  {32'h45e82cbc, 32'h00000000} /* (11, 29, 7) {real, imag} */,
  {32'h4617041c, 32'h00000000} /* (11, 29, 6) {real, imag} */,
  {32'h46239c08, 32'h00000000} /* (11, 29, 5) {real, imag} */,
  {32'h4635a6f3, 32'h00000000} /* (11, 29, 4) {real, imag} */,
  {32'h463c49f8, 32'h00000000} /* (11, 29, 3) {real, imag} */,
  {32'h463dc70a, 32'h00000000} /* (11, 29, 2) {real, imag} */,
  {32'h4644002b, 32'h00000000} /* (11, 29, 1) {real, imag} */,
  {32'h463e1629, 32'h00000000} /* (11, 29, 0) {real, imag} */,
  {32'h4644db73, 32'h00000000} /* (11, 28, 31) {real, imag} */,
  {32'h46552c2e, 32'h00000000} /* (11, 28, 30) {real, imag} */,
  {32'h465913c5, 32'h00000000} /* (11, 28, 29) {real, imag} */,
  {32'h464f3f80, 32'h00000000} /* (11, 28, 28) {real, imag} */,
  {32'h46579ae8, 32'h00000000} /* (11, 28, 27) {real, imag} */,
  {32'h46513541, 32'h00000000} /* (11, 28, 26) {real, imag} */,
  {32'h4643fec7, 32'h00000000} /* (11, 28, 25) {real, imag} */,
  {32'h4629cfc8, 32'h00000000} /* (11, 28, 24) {real, imag} */,
  {32'h462176df, 32'h00000000} /* (11, 28, 23) {real, imag} */,
  {32'h45fbd628, 32'h00000000} /* (11, 28, 22) {real, imag} */,
  {32'h458b3e34, 32'h00000000} /* (11, 28, 21) {real, imag} */,
  {32'hc46b1210, 32'h00000000} /* (11, 28, 20) {real, imag} */,
  {32'hc53c50d6, 32'h00000000} /* (11, 28, 19) {real, imag} */,
  {32'hc5ac94ec, 32'h00000000} /* (11, 28, 18) {real, imag} */,
  {32'hc5e3e9b3, 32'h00000000} /* (11, 28, 17) {real, imag} */,
  {32'hc5f72ca0, 32'h00000000} /* (11, 28, 16) {real, imag} */,
  {32'hc604138d, 32'h00000000} /* (11, 28, 15) {real, imag} */,
  {32'hc5e6fedb, 32'h00000000} /* (11, 28, 14) {real, imag} */,
  {32'hc5cd2b6a, 32'h00000000} /* (11, 28, 13) {real, imag} */,
  {32'hc596d098, 32'h00000000} /* (11, 28, 12) {real, imag} */,
  {32'hc4d38efc, 32'h00000000} /* (11, 28, 11) {real, imag} */,
  {32'h4444e8b0, 32'h00000000} /* (11, 28, 10) {real, imag} */,
  {32'h45843362, 32'h00000000} /* (11, 28, 9) {real, imag} */,
  {32'h45d83ddd, 32'h00000000} /* (11, 28, 8) {real, imag} */,
  {32'h45f62d26, 32'h00000000} /* (11, 28, 7) {real, imag} */,
  {32'h461f3eb4, 32'h00000000} /* (11, 28, 6) {real, imag} */,
  {32'h462e5f6e, 32'h00000000} /* (11, 28, 5) {real, imag} */,
  {32'h463beb79, 32'h00000000} /* (11, 28, 4) {real, imag} */,
  {32'h4641bb70, 32'h00000000} /* (11, 28, 3) {real, imag} */,
  {32'h464ced90, 32'h00000000} /* (11, 28, 2) {real, imag} */,
  {32'h464949ce, 32'h00000000} /* (11, 28, 1) {real, imag} */,
  {32'h463f8a1e, 32'h00000000} /* (11, 28, 0) {real, imag} */,
  {32'h46490483, 32'h00000000} /* (11, 27, 31) {real, imag} */,
  {32'h464fbc2e, 32'h00000000} /* (11, 27, 30) {real, imag} */,
  {32'h465f7fe9, 32'h00000000} /* (11, 27, 29) {real, imag} */,
  {32'h46534540, 32'h00000000} /* (11, 27, 28) {real, imag} */,
  {32'h4645b9d0, 32'h00000000} /* (11, 27, 27) {real, imag} */,
  {32'h465ad26d, 32'h00000000} /* (11, 27, 26) {real, imag} */,
  {32'h46465299, 32'h00000000} /* (11, 27, 25) {real, imag} */,
  {32'h4624cf1e, 32'h00000000} /* (11, 27, 24) {real, imag} */,
  {32'h46289185, 32'h00000000} /* (11, 27, 23) {real, imag} */,
  {32'h45ec6358, 32'h00000000} /* (11, 27, 22) {real, imag} */,
  {32'h4538e34a, 32'h00000000} /* (11, 27, 21) {real, imag} */,
  {32'hc48178bc, 32'h00000000} /* (11, 27, 20) {real, imag} */,
  {32'hc58e88d8, 32'h00000000} /* (11, 27, 19) {real, imag} */,
  {32'hc5cded56, 32'h00000000} /* (11, 27, 18) {real, imag} */,
  {32'hc5eb71fd, 32'h00000000} /* (11, 27, 17) {real, imag} */,
  {32'hc607f47a, 32'h00000000} /* (11, 27, 16) {real, imag} */,
  {32'hc602b0ad, 32'h00000000} /* (11, 27, 15) {real, imag} */,
  {32'hc60005ba, 32'h00000000} /* (11, 27, 14) {real, imag} */,
  {32'hc5b86d32, 32'h00000000} /* (11, 27, 13) {real, imag} */,
  {32'hc5848469, 32'h00000000} /* (11, 27, 12) {real, imag} */,
  {32'hc51e6770, 32'h00000000} /* (11, 27, 11) {real, imag} */,
  {32'h449545c8, 32'h00000000} /* (11, 27, 10) {real, imag} */,
  {32'h458beb8e, 32'h00000000} /* (11, 27, 9) {real, imag} */,
  {32'h45e52acc, 32'h00000000} /* (11, 27, 8) {real, imag} */,
  {32'h4615af73, 32'h00000000} /* (11, 27, 7) {real, imag} */,
  {32'h462e73da, 32'h00000000} /* (11, 27, 6) {real, imag} */,
  {32'h4628f9b6, 32'h00000000} /* (11, 27, 5) {real, imag} */,
  {32'h464b2084, 32'h00000000} /* (11, 27, 4) {real, imag} */,
  {32'h463e1246, 32'h00000000} /* (11, 27, 3) {real, imag} */,
  {32'h463d79c7, 32'h00000000} /* (11, 27, 2) {real, imag} */,
  {32'h46422adc, 32'h00000000} /* (11, 27, 1) {real, imag} */,
  {32'h463e3a70, 32'h00000000} /* (11, 27, 0) {real, imag} */,
  {32'h4635b3f4, 32'h00000000} /* (11, 26, 31) {real, imag} */,
  {32'h46518b92, 32'h00000000} /* (11, 26, 30) {real, imag} */,
  {32'h465586a2, 32'h00000000} /* (11, 26, 29) {real, imag} */,
  {32'h464a9fc8, 32'h00000000} /* (11, 26, 28) {real, imag} */,
  {32'h464d3db5, 32'h00000000} /* (11, 26, 27) {real, imag} */,
  {32'h463fb20f, 32'h00000000} /* (11, 26, 26) {real, imag} */,
  {32'h46381bf4, 32'h00000000} /* (11, 26, 25) {real, imag} */,
  {32'h46297754, 32'h00000000} /* (11, 26, 24) {real, imag} */,
  {32'h460d4de3, 32'h00000000} /* (11, 26, 23) {real, imag} */,
  {32'h45c0d9cb, 32'h00000000} /* (11, 26, 22) {real, imag} */,
  {32'h451c573a, 32'h00000000} /* (11, 26, 21) {real, imag} */,
  {32'hc48a7138, 32'h00000000} /* (11, 26, 20) {real, imag} */,
  {32'hc5844fe0, 32'h00000000} /* (11, 26, 19) {real, imag} */,
  {32'hc5bbd874, 32'h00000000} /* (11, 26, 18) {real, imag} */,
  {32'hc5ed9357, 32'h00000000} /* (11, 26, 17) {real, imag} */,
  {32'hc60893ce, 32'h00000000} /* (11, 26, 16) {real, imag} */,
  {32'hc60c8c7e, 32'h00000000} /* (11, 26, 15) {real, imag} */,
  {32'hc5feb628, 32'h00000000} /* (11, 26, 14) {real, imag} */,
  {32'hc5c4ed28, 32'h00000000} /* (11, 26, 13) {real, imag} */,
  {32'hc5811140, 32'h00000000} /* (11, 26, 12) {real, imag} */,
  {32'hc4e7ee08, 32'h00000000} /* (11, 26, 11) {real, imag} */,
  {32'h44d91b68, 32'h00000000} /* (11, 26, 10) {real, imag} */,
  {32'h45a0924f, 32'h00000000} /* (11, 26, 9) {real, imag} */,
  {32'h45f341c0, 32'h00000000} /* (11, 26, 8) {real, imag} */,
  {32'h46132a2b, 32'h00000000} /* (11, 26, 7) {real, imag} */,
  {32'h461a8ea8, 32'h00000000} /* (11, 26, 6) {real, imag} */,
  {32'h462cc6b2, 32'h00000000} /* (11, 26, 5) {real, imag} */,
  {32'h4634e6b9, 32'h00000000} /* (11, 26, 4) {real, imag} */,
  {32'h46396dd4, 32'h00000000} /* (11, 26, 3) {real, imag} */,
  {32'h4635e89a, 32'h00000000} /* (11, 26, 2) {real, imag} */,
  {32'h463ae046, 32'h00000000} /* (11, 26, 1) {real, imag} */,
  {32'h464085f6, 32'h00000000} /* (11, 26, 0) {real, imag} */,
  {32'h46218e10, 32'h00000000} /* (11, 25, 31) {real, imag} */,
  {32'h462f3b79, 32'h00000000} /* (11, 25, 30) {real, imag} */,
  {32'h463c364b, 32'h00000000} /* (11, 25, 29) {real, imag} */,
  {32'h4641b82b, 32'h00000000} /* (11, 25, 28) {real, imag} */,
  {32'h4635c281, 32'h00000000} /* (11, 25, 27) {real, imag} */,
  {32'h462adf83, 32'h00000000} /* (11, 25, 26) {real, imag} */,
  {32'h4638fc7c, 32'h00000000} /* (11, 25, 25) {real, imag} */,
  {32'h4616df37, 32'h00000000} /* (11, 25, 24) {real, imag} */,
  {32'h45e4e658, 32'h00000000} /* (11, 25, 23) {real, imag} */,
  {32'h45abd0fa, 32'h00000000} /* (11, 25, 22) {real, imag} */,
  {32'h44eb1e04, 32'h00000000} /* (11, 25, 21) {real, imag} */,
  {32'hc496f504, 32'h00000000} /* (11, 25, 20) {real, imag} */,
  {32'hc57ad8f7, 32'h00000000} /* (11, 25, 19) {real, imag} */,
  {32'hc5cb860b, 32'h00000000} /* (11, 25, 18) {real, imag} */,
  {32'hc609e9d2, 32'h00000000} /* (11, 25, 17) {real, imag} */,
  {32'hc6114698, 32'h00000000} /* (11, 25, 16) {real, imag} */,
  {32'hc5e4b920, 32'h00000000} /* (11, 25, 15) {real, imag} */,
  {32'hc5c62fb6, 32'h00000000} /* (11, 25, 14) {real, imag} */,
  {32'hc5a9cb36, 32'h00000000} /* (11, 25, 13) {real, imag} */,
  {32'hc59e4d3a, 32'h00000000} /* (11, 25, 12) {real, imag} */,
  {32'hc4f2b2b8, 32'h00000000} /* (11, 25, 11) {real, imag} */,
  {32'h44d3cc30, 32'h00000000} /* (11, 25, 10) {real, imag} */,
  {32'h45b38898, 32'h00000000} /* (11, 25, 9) {real, imag} */,
  {32'h45fede22, 32'h00000000} /* (11, 25, 8) {real, imag} */,
  {32'h461180f2, 32'h00000000} /* (11, 25, 7) {real, imag} */,
  {32'h4613152d, 32'h00000000} /* (11, 25, 6) {real, imag} */,
  {32'h462be290, 32'h00000000} /* (11, 25, 5) {real, imag} */,
  {32'h4637b352, 32'h00000000} /* (11, 25, 4) {real, imag} */,
  {32'h46325d81, 32'h00000000} /* (11, 25, 3) {real, imag} */,
  {32'h463212a4, 32'h00000000} /* (11, 25, 2) {real, imag} */,
  {32'h4625cbf6, 32'h00000000} /* (11, 25, 1) {real, imag} */,
  {32'h4621281a, 32'h00000000} /* (11, 25, 0) {real, imag} */,
  {32'h460d62df, 32'h00000000} /* (11, 24, 31) {real, imag} */,
  {32'h4619e802, 32'h00000000} /* (11, 24, 30) {real, imag} */,
  {32'h461b3e8b, 32'h00000000} /* (11, 24, 29) {real, imag} */,
  {32'h462549c4, 32'h00000000} /* (11, 24, 28) {real, imag} */,
  {32'h462879b2, 32'h00000000} /* (11, 24, 27) {real, imag} */,
  {32'h460ff0a8, 32'h00000000} /* (11, 24, 26) {real, imag} */,
  {32'h46145144, 32'h00000000} /* (11, 24, 25) {real, imag} */,
  {32'h4603cb86, 32'h00000000} /* (11, 24, 24) {real, imag} */,
  {32'h45c17b54, 32'h00000000} /* (11, 24, 23) {real, imag} */,
  {32'h4587a507, 32'h00000000} /* (11, 24, 22) {real, imag} */,
  {32'h447cb9d8, 32'h00000000} /* (11, 24, 21) {real, imag} */,
  {32'hc5371046, 32'h00000000} /* (11, 24, 20) {real, imag} */,
  {32'hc5929c67, 32'h00000000} /* (11, 24, 19) {real, imag} */,
  {32'hc5d69aa8, 32'h00000000} /* (11, 24, 18) {real, imag} */,
  {32'hc60481c6, 32'h00000000} /* (11, 24, 17) {real, imag} */,
  {32'hc5d1375c, 32'h00000000} /* (11, 24, 16) {real, imag} */,
  {32'hc5cfc16c, 32'h00000000} /* (11, 24, 15) {real, imag} */,
  {32'hc5a4ccf4, 32'h00000000} /* (11, 24, 14) {real, imag} */,
  {32'hc5a3d8f6, 32'h00000000} /* (11, 24, 13) {real, imag} */,
  {32'hc58500b7, 32'h00000000} /* (11, 24, 12) {real, imag} */,
  {32'hc446efb8, 32'h00000000} /* (11, 24, 11) {real, imag} */,
  {32'h450f9ab2, 32'h00000000} /* (11, 24, 10) {real, imag} */,
  {32'h45bd0090, 32'h00000000} /* (11, 24, 9) {real, imag} */,
  {32'h45e2996d, 32'h00000000} /* (11, 24, 8) {real, imag} */,
  {32'h460c7448, 32'h00000000} /* (11, 24, 7) {real, imag} */,
  {32'h46139bb6, 32'h00000000} /* (11, 24, 6) {real, imag} */,
  {32'h461393be, 32'h00000000} /* (11, 24, 5) {real, imag} */,
  {32'h461d6e98, 32'h00000000} /* (11, 24, 4) {real, imag} */,
  {32'h462d3bcc, 32'h00000000} /* (11, 24, 3) {real, imag} */,
  {32'h461d9e26, 32'h00000000} /* (11, 24, 2) {real, imag} */,
  {32'h460de706, 32'h00000000} /* (11, 24, 1) {real, imag} */,
  {32'h46031e07, 32'h00000000} /* (11, 24, 0) {real, imag} */,
  {32'h45ebd7f9, 32'h00000000} /* (11, 23, 31) {real, imag} */,
  {32'h4601ad63, 32'h00000000} /* (11, 23, 30) {real, imag} */,
  {32'h45ffdc9a, 32'h00000000} /* (11, 23, 29) {real, imag} */,
  {32'h46003af0, 32'h00000000} /* (11, 23, 28) {real, imag} */,
  {32'h46009a68, 32'h00000000} /* (11, 23, 27) {real, imag} */,
  {32'h45f688d8, 32'h00000000} /* (11, 23, 26) {real, imag} */,
  {32'h45d2e132, 32'h00000000} /* (11, 23, 25) {real, imag} */,
  {32'h45c522cd, 32'h00000000} /* (11, 23, 24) {real, imag} */,
  {32'h459cc9f6, 32'h00000000} /* (11, 23, 23) {real, imag} */,
  {32'h453cf668, 32'h00000000} /* (11, 23, 22) {real, imag} */,
  {32'h44896a60, 32'h00000000} /* (11, 23, 21) {real, imag} */,
  {32'hc524237e, 32'h00000000} /* (11, 23, 20) {real, imag} */,
  {32'hc598152d, 32'h00000000} /* (11, 23, 19) {real, imag} */,
  {32'hc5ae0304, 32'h00000000} /* (11, 23, 18) {real, imag} */,
  {32'hc5c46129, 32'h00000000} /* (11, 23, 17) {real, imag} */,
  {32'hc5b05af4, 32'h00000000} /* (11, 23, 16) {real, imag} */,
  {32'hc5a1ec4d, 32'h00000000} /* (11, 23, 15) {real, imag} */,
  {32'hc596c1b8, 32'h00000000} /* (11, 23, 14) {real, imag} */,
  {32'hc583e912, 32'h00000000} /* (11, 23, 13) {real, imag} */,
  {32'hc54790b6, 32'h00000000} /* (11, 23, 12) {real, imag} */,
  {32'hc4ac3b10, 32'h00000000} /* (11, 23, 11) {real, imag} */,
  {32'h44bec340, 32'h00000000} /* (11, 23, 10) {real, imag} */,
  {32'h459cc72e, 32'h00000000} /* (11, 23, 9) {real, imag} */,
  {32'h45b4e4df, 32'h00000000} /* (11, 23, 8) {real, imag} */,
  {32'h45d93b84, 32'h00000000} /* (11, 23, 7) {real, imag} */,
  {32'h45e8d45c, 32'h00000000} /* (11, 23, 6) {real, imag} */,
  {32'h45ef44ac, 32'h00000000} /* (11, 23, 5) {real, imag} */,
  {32'h4600838c, 32'h00000000} /* (11, 23, 4) {real, imag} */,
  {32'h460626eb, 32'h00000000} /* (11, 23, 3) {real, imag} */,
  {32'h45f37634, 32'h00000000} /* (11, 23, 2) {real, imag} */,
  {32'h45fd1369, 32'h00000000} /* (11, 23, 1) {real, imag} */,
  {32'h45e7b840, 32'h00000000} /* (11, 23, 0) {real, imag} */,
  {32'h458f2f11, 32'h00000000} /* (11, 22, 31) {real, imag} */,
  {32'h45b77d89, 32'h00000000} /* (11, 22, 30) {real, imag} */,
  {32'h45bb36f0, 32'h00000000} /* (11, 22, 29) {real, imag} */,
  {32'h45b0d8c2, 32'h00000000} /* (11, 22, 28) {real, imag} */,
  {32'h45a45d7f, 32'h00000000} /* (11, 22, 27) {real, imag} */,
  {32'h459bf0fc, 32'h00000000} /* (11, 22, 26) {real, imag} */,
  {32'h45899ecf, 32'h00000000} /* (11, 22, 25) {real, imag} */,
  {32'h4581631a, 32'h00000000} /* (11, 22, 24) {real, imag} */,
  {32'h45818849, 32'h00000000} /* (11, 22, 23) {real, imag} */,
  {32'h452db2f9, 32'h00000000} /* (11, 22, 22) {real, imag} */,
  {32'h4445e070, 32'h00000000} /* (11, 22, 21) {real, imag} */,
  {32'hc505eb4c, 32'h00000000} /* (11, 22, 20) {real, imag} */,
  {32'hc579a65a, 32'h00000000} /* (11, 22, 19) {real, imag} */,
  {32'hc5622507, 32'h00000000} /* (11, 22, 18) {real, imag} */,
  {32'hc5598514, 32'h00000000} /* (11, 22, 17) {real, imag} */,
  {32'hc58da699, 32'h00000000} /* (11, 22, 16) {real, imag} */,
  {32'hc5509454, 32'h00000000} /* (11, 22, 15) {real, imag} */,
  {32'hc540b52a, 32'h00000000} /* (11, 22, 14) {real, imag} */,
  {32'hc53abdcb, 32'h00000000} /* (11, 22, 13) {real, imag} */,
  {32'hc52ae858, 32'h00000000} /* (11, 22, 12) {real, imag} */,
  {32'hc50acf3e, 32'h00000000} /* (11, 22, 11) {real, imag} */,
  {32'h447988ac, 32'h00000000} /* (11, 22, 10) {real, imag} */,
  {32'h454ec302, 32'h00000000} /* (11, 22, 9) {real, imag} */,
  {32'h458da52e, 32'h00000000} /* (11, 22, 8) {real, imag} */,
  {32'h4589b6b1, 32'h00000000} /* (11, 22, 7) {real, imag} */,
  {32'h459bc316, 32'h00000000} /* (11, 22, 6) {real, imag} */,
  {32'h458bc443, 32'h00000000} /* (11, 22, 5) {real, imag} */,
  {32'h45979461, 32'h00000000} /* (11, 22, 4) {real, imag} */,
  {32'h459b8d79, 32'h00000000} /* (11, 22, 3) {real, imag} */,
  {32'h45a96dc4, 32'h00000000} /* (11, 22, 2) {real, imag} */,
  {32'h45c894b2, 32'h00000000} /* (11, 22, 1) {real, imag} */,
  {32'h45ac2a77, 32'h00000000} /* (11, 22, 0) {real, imag} */,
  {32'h44da69fc, 32'h00000000} /* (11, 21, 31) {real, imag} */,
  {32'h44e752fc, 32'h00000000} /* (11, 21, 30) {real, imag} */,
  {32'h452428c2, 32'h00000000} /* (11, 21, 29) {real, imag} */,
  {32'h455ac92b, 32'h00000000} /* (11, 21, 28) {real, imag} */,
  {32'h44ff666f, 32'h00000000} /* (11, 21, 27) {real, imag} */,
  {32'h44b2212c, 32'h00000000} /* (11, 21, 26) {real, imag} */,
  {32'h44db78fe, 32'h00000000} /* (11, 21, 25) {real, imag} */,
  {32'h44e992b8, 32'h00000000} /* (11, 21, 24) {real, imag} */,
  {32'h43b0da8c, 32'h00000000} /* (11, 21, 23) {real, imag} */,
  {32'h438b5896, 32'h00000000} /* (11, 21, 22) {real, imag} */,
  {32'h44045d5d, 32'h00000000} /* (11, 21, 21) {real, imag} */,
  {32'hc43bdd45, 32'h00000000} /* (11, 21, 20) {real, imag} */,
  {32'hc4979178, 32'h00000000} /* (11, 21, 19) {real, imag} */,
  {32'hc4cdbf34, 32'h00000000} /* (11, 21, 18) {real, imag} */,
  {32'hc47f5b5e, 32'h00000000} /* (11, 21, 17) {real, imag} */,
  {32'hc454025a, 32'h00000000} /* (11, 21, 16) {real, imag} */,
  {32'hc39b8628, 32'h00000000} /* (11, 21, 15) {real, imag} */,
  {32'hc4552974, 32'h00000000} /* (11, 21, 14) {real, imag} */,
  {32'hc4a4b8da, 32'h00000000} /* (11, 21, 13) {real, imag} */,
  {32'hc35b5570, 32'h00000000} /* (11, 21, 12) {real, imag} */,
  {32'hc34829c8, 32'h00000000} /* (11, 21, 11) {real, imag} */,
  {32'h4386246c, 32'h00000000} /* (11, 21, 10) {real, imag} */,
  {32'h443edcec, 32'h00000000} /* (11, 21, 9) {real, imag} */,
  {32'h444d68c5, 32'h00000000} /* (11, 21, 8) {real, imag} */,
  {32'h448040a3, 32'h00000000} /* (11, 21, 7) {real, imag} */,
  {32'h44ef7ea2, 32'h00000000} /* (11, 21, 6) {real, imag} */,
  {32'h44e79e02, 32'h00000000} /* (11, 21, 5) {real, imag} */,
  {32'h44fcea96, 32'h00000000} /* (11, 21, 4) {real, imag} */,
  {32'h450c7d59, 32'h00000000} /* (11, 21, 3) {real, imag} */,
  {32'h44eedb38, 32'h00000000} /* (11, 21, 2) {real, imag} */,
  {32'h452b2516, 32'h00000000} /* (11, 21, 1) {real, imag} */,
  {32'h44cbad43, 32'h00000000} /* (11, 21, 0) {real, imag} */,
  {32'hc4cf3a50, 32'h00000000} /* (11, 20, 31) {real, imag} */,
  {32'hc52e2ba7, 32'h00000000} /* (11, 20, 30) {real, imag} */,
  {32'hc510907d, 32'h00000000} /* (11, 20, 29) {real, imag} */,
  {32'hc4d19f45, 32'h00000000} /* (11, 20, 28) {real, imag} */,
  {32'hc4bdb592, 32'h00000000} /* (11, 20, 27) {real, imag} */,
  {32'hc48aeef5, 32'h00000000} /* (11, 20, 26) {real, imag} */,
  {32'hc5115cf9, 32'h00000000} /* (11, 20, 25) {real, imag} */,
  {32'hc527802b, 32'h00000000} /* (11, 20, 24) {real, imag} */,
  {32'hc4c03c6d, 32'h00000000} /* (11, 20, 23) {real, imag} */,
  {32'hc4fcc538, 32'h00000000} /* (11, 20, 22) {real, imag} */,
  {32'hc463afbe, 32'h00000000} /* (11, 20, 21) {real, imag} */,
  {32'h43579188, 32'h00000000} /* (11, 20, 20) {real, imag} */,
  {32'h44aaa99f, 32'h00000000} /* (11, 20, 19) {real, imag} */,
  {32'h45199b01, 32'h00000000} /* (11, 20, 18) {real, imag} */,
  {32'h4523fe2e, 32'h00000000} /* (11, 20, 17) {real, imag} */,
  {32'h45615a2d, 32'h00000000} /* (11, 20, 16) {real, imag} */,
  {32'h45518636, 32'h00000000} /* (11, 20, 15) {real, imag} */,
  {32'h451eeec5, 32'h00000000} /* (11, 20, 14) {real, imag} */,
  {32'h4501d5cb, 32'h00000000} /* (11, 20, 13) {real, imag} */,
  {32'h45118469, 32'h00000000} /* (11, 20, 12) {real, imag} */,
  {32'h44b17142, 32'h00000000} /* (11, 20, 11) {real, imag} */,
  {32'hc4952207, 32'h00000000} /* (11, 20, 10) {real, imag} */,
  {32'hc4a44bde, 32'h00000000} /* (11, 20, 9) {real, imag} */,
  {32'hc4d1dfd6, 32'h00000000} /* (11, 20, 8) {real, imag} */,
  {32'hc4f44c77, 32'h00000000} /* (11, 20, 7) {real, imag} */,
  {32'hc51264ca, 32'h00000000} /* (11, 20, 6) {real, imag} */,
  {32'hc53b56ca, 32'h00000000} /* (11, 20, 5) {real, imag} */,
  {32'hc503238a, 32'h00000000} /* (11, 20, 4) {real, imag} */,
  {32'hc4d2b411, 32'h00000000} /* (11, 20, 3) {real, imag} */,
  {32'hc5241ca1, 32'h00000000} /* (11, 20, 2) {real, imag} */,
  {32'hc532a656, 32'h00000000} /* (11, 20, 1) {real, imag} */,
  {32'hc4c3e24a, 32'h00000000} /* (11, 20, 0) {real, imag} */,
  {32'hc58999d1, 32'h00000000} /* (11, 19, 31) {real, imag} */,
  {32'hc5b34464, 32'h00000000} /* (11, 19, 30) {real, imag} */,
  {32'hc5c3fcff, 32'h00000000} /* (11, 19, 29) {real, imag} */,
  {32'hc59f6820, 32'h00000000} /* (11, 19, 28) {real, imag} */,
  {32'hc592d639, 32'h00000000} /* (11, 19, 27) {real, imag} */,
  {32'hc5a6756b, 32'h00000000} /* (11, 19, 26) {real, imag} */,
  {32'hc5a1de10, 32'h00000000} /* (11, 19, 25) {real, imag} */,
  {32'hc5a59ea4, 32'h00000000} /* (11, 19, 24) {real, imag} */,
  {32'hc5436a46, 32'h00000000} /* (11, 19, 23) {real, imag} */,
  {32'hc5331de9, 32'h00000000} /* (11, 19, 22) {real, imag} */,
  {32'hc4aa2ca0, 32'h00000000} /* (11, 19, 21) {real, imag} */,
  {32'h44f9a1b9, 32'h00000000} /* (11, 19, 20) {real, imag} */,
  {32'h45146e1a, 32'h00000000} /* (11, 19, 19) {real, imag} */,
  {32'h455de67c, 32'h00000000} /* (11, 19, 18) {real, imag} */,
  {32'h4594f7cc, 32'h00000000} /* (11, 19, 17) {real, imag} */,
  {32'h45af324c, 32'h00000000} /* (11, 19, 16) {real, imag} */,
  {32'h45d60e01, 32'h00000000} /* (11, 19, 15) {real, imag} */,
  {32'h4596ab9e, 32'h00000000} /* (11, 19, 14) {real, imag} */,
  {32'h4583b331, 32'h00000000} /* (11, 19, 13) {real, imag} */,
  {32'h454b0d58, 32'h00000000} /* (11, 19, 12) {real, imag} */,
  {32'h44b73430, 32'h00000000} /* (11, 19, 11) {real, imag} */,
  {32'hc4aa21e3, 32'h00000000} /* (11, 19, 10) {real, imag} */,
  {32'hc5329348, 32'h00000000} /* (11, 19, 9) {real, imag} */,
  {32'hc543768b, 32'h00000000} /* (11, 19, 8) {real, imag} */,
  {32'hc581a24b, 32'h00000000} /* (11, 19, 7) {real, imag} */,
  {32'hc591ba64, 32'h00000000} /* (11, 19, 6) {real, imag} */,
  {32'hc5a02846, 32'h00000000} /* (11, 19, 5) {real, imag} */,
  {32'hc5b7ab12, 32'h00000000} /* (11, 19, 4) {real, imag} */,
  {32'hc5b28f64, 32'h00000000} /* (11, 19, 3) {real, imag} */,
  {32'hc5a181cc, 32'h00000000} /* (11, 19, 2) {real, imag} */,
  {32'hc596415a, 32'h00000000} /* (11, 19, 1) {real, imag} */,
  {32'hc594c1aa, 32'h00000000} /* (11, 19, 0) {real, imag} */,
  {32'hc5dc6f0c, 32'h00000000} /* (11, 18, 31) {real, imag} */,
  {32'hc5fc2886, 32'h00000000} /* (11, 18, 30) {real, imag} */,
  {32'hc60086b2, 32'h00000000} /* (11, 18, 29) {real, imag} */,
  {32'hc6018aee, 32'h00000000} /* (11, 18, 28) {real, imag} */,
  {32'hc5ec1104, 32'h00000000} /* (11, 18, 27) {real, imag} */,
  {32'hc5e5bef2, 32'h00000000} /* (11, 18, 26) {real, imag} */,
  {32'hc5d893bf, 32'h00000000} /* (11, 18, 25) {real, imag} */,
  {32'hc5b56191, 32'h00000000} /* (11, 18, 24) {real, imag} */,
  {32'hc5ac3e64, 32'h00000000} /* (11, 18, 23) {real, imag} */,
  {32'hc580bb83, 32'h00000000} /* (11, 18, 22) {real, imag} */,
  {32'hc4857680, 32'h00000000} /* (11, 18, 21) {real, imag} */,
  {32'h44ea319c, 32'h00000000} /* (11, 18, 20) {real, imag} */,
  {32'h45872bea, 32'h00000000} /* (11, 18, 19) {real, imag} */,
  {32'h458cf584, 32'h00000000} /* (11, 18, 18) {real, imag} */,
  {32'h45ae8266, 32'h00000000} /* (11, 18, 17) {real, imag} */,
  {32'h45bec5a4, 32'h00000000} /* (11, 18, 16) {real, imag} */,
  {32'h45dc8e0e, 32'h00000000} /* (11, 18, 15) {real, imag} */,
  {32'h45abd93a, 32'h00000000} /* (11, 18, 14) {real, imag} */,
  {32'h45af708e, 32'h00000000} /* (11, 18, 13) {real, imag} */,
  {32'h45698560, 32'h00000000} /* (11, 18, 12) {real, imag} */,
  {32'h44b033b8, 32'h00000000} /* (11, 18, 11) {real, imag} */,
  {32'hc49a8118, 32'h00000000} /* (11, 18, 10) {real, imag} */,
  {32'hc530d1c2, 32'h00000000} /* (11, 18, 9) {real, imag} */,
  {32'hc58a134b, 32'h00000000} /* (11, 18, 8) {real, imag} */,
  {32'hc5def230, 32'h00000000} /* (11, 18, 7) {real, imag} */,
  {32'hc5da0635, 32'h00000000} /* (11, 18, 6) {real, imag} */,
  {32'hc5e94ae2, 32'h00000000} /* (11, 18, 5) {real, imag} */,
  {32'hc5e492ff, 32'h00000000} /* (11, 18, 4) {real, imag} */,
  {32'hc5d68be0, 32'h00000000} /* (11, 18, 3) {real, imag} */,
  {32'hc5eb7212, 32'h00000000} /* (11, 18, 2) {real, imag} */,
  {32'hc5d83986, 32'h00000000} /* (11, 18, 1) {real, imag} */,
  {32'hc5c344a0, 32'h00000000} /* (11, 18, 0) {real, imag} */,
  {32'hc5e92a10, 32'h00000000} /* (11, 17, 31) {real, imag} */,
  {32'hc5ff23ec, 32'h00000000} /* (11, 17, 30) {real, imag} */,
  {32'hc60a2844, 32'h00000000} /* (11, 17, 29) {real, imag} */,
  {32'hc60fa1c0, 32'h00000000} /* (11, 17, 28) {real, imag} */,
  {32'hc609c190, 32'h00000000} /* (11, 17, 27) {real, imag} */,
  {32'hc602a568, 32'h00000000} /* (11, 17, 26) {real, imag} */,
  {32'hc5edc562, 32'h00000000} /* (11, 17, 25) {real, imag} */,
  {32'hc5d42e80, 32'h00000000} /* (11, 17, 24) {real, imag} */,
  {32'hc5d80757, 32'h00000000} /* (11, 17, 23) {real, imag} */,
  {32'hc57ec442, 32'h00000000} /* (11, 17, 22) {real, imag} */,
  {32'hc4c08ee8, 32'h00000000} /* (11, 17, 21) {real, imag} */,
  {32'h450aa3a0, 32'h00000000} /* (11, 17, 20) {real, imag} */,
  {32'h459f0844, 32'h00000000} /* (11, 17, 19) {real, imag} */,
  {32'h45ddffe2, 32'h00000000} /* (11, 17, 18) {real, imag} */,
  {32'h45d3b5b7, 32'h00000000} /* (11, 17, 17) {real, imag} */,
  {32'h45d982c4, 32'h00000000} /* (11, 17, 16) {real, imag} */,
  {32'h45e73604, 32'h00000000} /* (11, 17, 15) {real, imag} */,
  {32'h45f28b6e, 32'h00000000} /* (11, 17, 14) {real, imag} */,
  {32'h45c7ae8f, 32'h00000000} /* (11, 17, 13) {real, imag} */,
  {32'h4592965f, 32'h00000000} /* (11, 17, 12) {real, imag} */,
  {32'h44eacf0c, 32'h00000000} /* (11, 17, 11) {real, imag} */,
  {32'hc4b2266c, 32'h00000000} /* (11, 17, 10) {real, imag} */,
  {32'hc548fc04, 32'h00000000} /* (11, 17, 9) {real, imag} */,
  {32'hc5a40fa2, 32'h00000000} /* (11, 17, 8) {real, imag} */,
  {32'hc5e2e5b1, 32'h00000000} /* (11, 17, 7) {real, imag} */,
  {32'hc61013a2, 32'h00000000} /* (11, 17, 6) {real, imag} */,
  {32'hc6061823, 32'h00000000} /* (11, 17, 5) {real, imag} */,
  {32'hc615165c, 32'h00000000} /* (11, 17, 4) {real, imag} */,
  {32'hc627ba64, 32'h00000000} /* (11, 17, 3) {real, imag} */,
  {32'hc612db17, 32'h00000000} /* (11, 17, 2) {real, imag} */,
  {32'hc5ff211b, 32'h00000000} /* (11, 17, 1) {real, imag} */,
  {32'hc5ee9f5a, 32'h00000000} /* (11, 17, 0) {real, imag} */,
  {32'hc609ce2e, 32'h00000000} /* (11, 16, 31) {real, imag} */,
  {32'hc614aa3e, 32'h00000000} /* (11, 16, 30) {real, imag} */,
  {32'hc60e772e, 32'h00000000} /* (11, 16, 29) {real, imag} */,
  {32'hc6202853, 32'h00000000} /* (11, 16, 28) {real, imag} */,
  {32'hc618dccd, 32'h00000000} /* (11, 16, 27) {real, imag} */,
  {32'hc60bde69, 32'h00000000} /* (11, 16, 26) {real, imag} */,
  {32'hc60157ee, 32'h00000000} /* (11, 16, 25) {real, imag} */,
  {32'hc5f7cfae, 32'h00000000} /* (11, 16, 24) {real, imag} */,
  {32'hc5c0d4d8, 32'h00000000} /* (11, 16, 23) {real, imag} */,
  {32'hc551966e, 32'h00000000} /* (11, 16, 22) {real, imag} */,
  {32'hc4ae751e, 32'h00000000} /* (11, 16, 21) {real, imag} */,
  {32'h451dbc09, 32'h00000000} /* (11, 16, 20) {real, imag} */,
  {32'h45a2168c, 32'h00000000} /* (11, 16, 19) {real, imag} */,
  {32'h45ca6404, 32'h00000000} /* (11, 16, 18) {real, imag} */,
  {32'h45e84b34, 32'h00000000} /* (11, 16, 17) {real, imag} */,
  {32'h460069a6, 32'h00000000} /* (11, 16, 16) {real, imag} */,
  {32'h45f4d7bc, 32'h00000000} /* (11, 16, 15) {real, imag} */,
  {32'h45f2d3d1, 32'h00000000} /* (11, 16, 14) {real, imag} */,
  {32'h45daf79d, 32'h00000000} /* (11, 16, 13) {real, imag} */,
  {32'h459b3f72, 32'h00000000} /* (11, 16, 12) {real, imag} */,
  {32'h45049168, 32'h00000000} /* (11, 16, 11) {real, imag} */,
  {32'hc505beab, 32'h00000000} /* (11, 16, 10) {real, imag} */,
  {32'hc5961311, 32'h00000000} /* (11, 16, 9) {real, imag} */,
  {32'hc5d668f4, 32'h00000000} /* (11, 16, 8) {real, imag} */,
  {32'hc5f68f00, 32'h00000000} /* (11, 16, 7) {real, imag} */,
  {32'hc5f1d7b3, 32'h00000000} /* (11, 16, 6) {real, imag} */,
  {32'hc60ebee0, 32'h00000000} /* (11, 16, 5) {real, imag} */,
  {32'hc6138134, 32'h00000000} /* (11, 16, 4) {real, imag} */,
  {32'hc62ea553, 32'h00000000} /* (11, 16, 3) {real, imag} */,
  {32'hc61db2f2, 32'h00000000} /* (11, 16, 2) {real, imag} */,
  {32'hc60edc9c, 32'h00000000} /* (11, 16, 1) {real, imag} */,
  {32'hc606a61c, 32'h00000000} /* (11, 16, 0) {real, imag} */,
  {32'hc606598c, 32'h00000000} /* (11, 15, 31) {real, imag} */,
  {32'hc61d3438, 32'h00000000} /* (11, 15, 30) {real, imag} */,
  {32'hc61e7494, 32'h00000000} /* (11, 15, 29) {real, imag} */,
  {32'hc616c099, 32'h00000000} /* (11, 15, 28) {real, imag} */,
  {32'hc6140d2a, 32'h00000000} /* (11, 15, 27) {real, imag} */,
  {32'hc6121bcf, 32'h00000000} /* (11, 15, 26) {real, imag} */,
  {32'hc60218c4, 32'h00000000} /* (11, 15, 25) {real, imag} */,
  {32'hc5e66d44, 32'h00000000} /* (11, 15, 24) {real, imag} */,
  {32'hc5be8d16, 32'h00000000} /* (11, 15, 23) {real, imag} */,
  {32'hc5465728, 32'h00000000} /* (11, 15, 22) {real, imag} */,
  {32'h449083a8, 32'h00000000} /* (11, 15, 21) {real, imag} */,
  {32'h4536a959, 32'h00000000} /* (11, 15, 20) {real, imag} */,
  {32'h458f2d00, 32'h00000000} /* (11, 15, 19) {real, imag} */,
  {32'h45c5dc84, 32'h00000000} /* (11, 15, 18) {real, imag} */,
  {32'h45e579e0, 32'h00000000} /* (11, 15, 17) {real, imag} */,
  {32'h45fd7928, 32'h00000000} /* (11, 15, 16) {real, imag} */,
  {32'h460415a8, 32'h00000000} /* (11, 15, 15) {real, imag} */,
  {32'h45dd9ca8, 32'h00000000} /* (11, 15, 14) {real, imag} */,
  {32'h45c5b121, 32'h00000000} /* (11, 15, 13) {real, imag} */,
  {32'h458a217c, 32'h00000000} /* (11, 15, 12) {real, imag} */,
  {32'h4510604f, 32'h00000000} /* (11, 15, 11) {real, imag} */,
  {32'hc4dca088, 32'h00000000} /* (11, 15, 10) {real, imag} */,
  {32'hc5a0ed30, 32'h00000000} /* (11, 15, 9) {real, imag} */,
  {32'hc5d617fc, 32'h00000000} /* (11, 15, 8) {real, imag} */,
  {32'hc6057320, 32'h00000000} /* (11, 15, 7) {real, imag} */,
  {32'hc60506ce, 32'h00000000} /* (11, 15, 6) {real, imag} */,
  {32'hc60c3bba, 32'h00000000} /* (11, 15, 5) {real, imag} */,
  {32'hc6177ceb, 32'h00000000} /* (11, 15, 4) {real, imag} */,
  {32'hc61a3623, 32'h00000000} /* (11, 15, 3) {real, imag} */,
  {32'hc61942aa, 32'h00000000} /* (11, 15, 2) {real, imag} */,
  {32'hc6157608, 32'h00000000} /* (11, 15, 1) {real, imag} */,
  {32'hc60fe714, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'hc6005368, 32'h00000000} /* (11, 14, 31) {real, imag} */,
  {32'hc61c7093, 32'h00000000} /* (11, 14, 30) {real, imag} */,
  {32'hc61d7d16, 32'h00000000} /* (11, 14, 29) {real, imag} */,
  {32'hc60638a5, 32'h00000000} /* (11, 14, 28) {real, imag} */,
  {32'hc6032c9a, 32'h00000000} /* (11, 14, 27) {real, imag} */,
  {32'hc606df72, 32'h00000000} /* (11, 14, 26) {real, imag} */,
  {32'hc5e2d340, 32'h00000000} /* (11, 14, 25) {real, imag} */,
  {32'hc5d24a46, 32'h00000000} /* (11, 14, 24) {real, imag} */,
  {32'hc5af013d, 32'h00000000} /* (11, 14, 23) {real, imag} */,
  {32'hc5591faf, 32'h00000000} /* (11, 14, 22) {real, imag} */,
  {32'hc4d9b6d4, 32'h00000000} /* (11, 14, 21) {real, imag} */,
  {32'h45383e27, 32'h00000000} /* (11, 14, 20) {real, imag} */,
  {32'h459d1c47, 32'h00000000} /* (11, 14, 19) {real, imag} */,
  {32'h45cbfa28, 32'h00000000} /* (11, 14, 18) {real, imag} */,
  {32'h45dacaa0, 32'h00000000} /* (11, 14, 17) {real, imag} */,
  {32'h45db3a5c, 32'h00000000} /* (11, 14, 16) {real, imag} */,
  {32'h45f3423d, 32'h00000000} /* (11, 14, 15) {real, imag} */,
  {32'h45ed9aea, 32'h00000000} /* (11, 14, 14) {real, imag} */,
  {32'h45ba3448, 32'h00000000} /* (11, 14, 13) {real, imag} */,
  {32'h45b92f3e, 32'h00000000} /* (11, 14, 12) {real, imag} */,
  {32'h45122d24, 32'h00000000} /* (11, 14, 11) {real, imag} */,
  {32'hc463d648, 32'h00000000} /* (11, 14, 10) {real, imag} */,
  {32'hc5786d10, 32'h00000000} /* (11, 14, 9) {real, imag} */,
  {32'hc5bf38a2, 32'h00000000} /* (11, 14, 8) {real, imag} */,
  {32'hc5efcea5, 32'h00000000} /* (11, 14, 7) {real, imag} */,
  {32'hc5fc8d72, 32'h00000000} /* (11, 14, 6) {real, imag} */,
  {32'hc5f3a61f, 32'h00000000} /* (11, 14, 5) {real, imag} */,
  {32'hc60986a6, 32'h00000000} /* (11, 14, 4) {real, imag} */,
  {32'hc60f37c6, 32'h00000000} /* (11, 14, 3) {real, imag} */,
  {32'hc60fb8f8, 32'h00000000} /* (11, 14, 2) {real, imag} */,
  {32'hc6122691, 32'h00000000} /* (11, 14, 1) {real, imag} */,
  {32'hc60ba29a, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'hc5ef961a, 32'h00000000} /* (11, 13, 31) {real, imag} */,
  {32'hc60d92c7, 32'h00000000} /* (11, 13, 30) {real, imag} */,
  {32'hc5e12ff0, 32'h00000000} /* (11, 13, 29) {real, imag} */,
  {32'hc5f8b030, 32'h00000000} /* (11, 13, 28) {real, imag} */,
  {32'hc5d25502, 32'h00000000} /* (11, 13, 27) {real, imag} */,
  {32'hc5cb6c7e, 32'h00000000} /* (11, 13, 26) {real, imag} */,
  {32'hc5df9174, 32'h00000000} /* (11, 13, 25) {real, imag} */,
  {32'hc5a51490, 32'h00000000} /* (11, 13, 24) {real, imag} */,
  {32'hc595b9a4, 32'h00000000} /* (11, 13, 23) {real, imag} */,
  {32'hc5438a62, 32'h00000000} /* (11, 13, 22) {real, imag} */,
  {32'hc487102a, 32'h00000000} /* (11, 13, 21) {real, imag} */,
  {32'h451052c5, 32'h00000000} /* (11, 13, 20) {real, imag} */,
  {32'h45a754f4, 32'h00000000} /* (11, 13, 19) {real, imag} */,
  {32'h45c27f8b, 32'h00000000} /* (11, 13, 18) {real, imag} */,
  {32'h45da878b, 32'h00000000} /* (11, 13, 17) {real, imag} */,
  {32'h45de21f4, 32'h00000000} /* (11, 13, 16) {real, imag} */,
  {32'h45df85d4, 32'h00000000} /* (11, 13, 15) {real, imag} */,
  {32'h45b7954e, 32'h00000000} /* (11, 13, 14) {real, imag} */,
  {32'h459fddd0, 32'h00000000} /* (11, 13, 13) {real, imag} */,
  {32'h457ee460, 32'h00000000} /* (11, 13, 12) {real, imag} */,
  {32'h45054311, 32'h00000000} /* (11, 13, 11) {real, imag} */,
  {32'hc48941e8, 32'h00000000} /* (11, 13, 10) {real, imag} */,
  {32'hc54f9eac, 32'h00000000} /* (11, 13, 9) {real, imag} */,
  {32'hc5a0f870, 32'h00000000} /* (11, 13, 8) {real, imag} */,
  {32'hc5b002c4, 32'h00000000} /* (11, 13, 7) {real, imag} */,
  {32'hc5f57cdb, 32'h00000000} /* (11, 13, 6) {real, imag} */,
  {32'hc5d517a2, 32'h00000000} /* (11, 13, 5) {real, imag} */,
  {32'hc5ccdd02, 32'h00000000} /* (11, 13, 4) {real, imag} */,
  {32'hc5e2f09a, 32'h00000000} /* (11, 13, 3) {real, imag} */,
  {32'hc5d993c1, 32'h00000000} /* (11, 13, 2) {real, imag} */,
  {32'hc5e5c7b7, 32'h00000000} /* (11, 13, 1) {real, imag} */,
  {32'hc5df0018, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'hc59da233, 32'h00000000} /* (11, 12, 31) {real, imag} */,
  {32'hc59db63d, 32'h00000000} /* (11, 12, 30) {real, imag} */,
  {32'hc59d7f24, 32'h00000000} /* (11, 12, 29) {real, imag} */,
  {32'hc59ad2fa, 32'h00000000} /* (11, 12, 28) {real, imag} */,
  {32'hc586419c, 32'h00000000} /* (11, 12, 27) {real, imag} */,
  {32'hc5717235, 32'h00000000} /* (11, 12, 26) {real, imag} */,
  {32'hc565f2be, 32'h00000000} /* (11, 12, 25) {real, imag} */,
  {32'hc5730e82, 32'h00000000} /* (11, 12, 24) {real, imag} */,
  {32'hc55e76b0, 32'h00000000} /* (11, 12, 23) {real, imag} */,
  {32'hc4ec3ca8, 32'h00000000} /* (11, 12, 22) {real, imag} */,
  {32'hc3d23240, 32'h00000000} /* (11, 12, 21) {real, imag} */,
  {32'h451276c2, 32'h00000000} /* (11, 12, 20) {real, imag} */,
  {32'h457d083d, 32'h00000000} /* (11, 12, 19) {real, imag} */,
  {32'h45b53e48, 32'h00000000} /* (11, 12, 18) {real, imag} */,
  {32'h45bd9f92, 32'h00000000} /* (11, 12, 17) {real, imag} */,
  {32'h45c1d76a, 32'h00000000} /* (11, 12, 16) {real, imag} */,
  {32'h45ae4f95, 32'h00000000} /* (11, 12, 15) {real, imag} */,
  {32'h45a0594f, 32'h00000000} /* (11, 12, 14) {real, imag} */,
  {32'h4577b844, 32'h00000000} /* (11, 12, 13) {real, imag} */,
  {32'h453b7270, 32'h00000000} /* (11, 12, 12) {real, imag} */,
  {32'h441f89d4, 32'h00000000} /* (11, 12, 11) {real, imag} */,
  {32'hc4ce8c16, 32'h00000000} /* (11, 12, 10) {real, imag} */,
  {32'hc5277ac6, 32'h00000000} /* (11, 12, 9) {real, imag} */,
  {32'hc5766278, 32'h00000000} /* (11, 12, 8) {real, imag} */,
  {32'hc5897c1e, 32'h00000000} /* (11, 12, 7) {real, imag} */,
  {32'hc5ad5758, 32'h00000000} /* (11, 12, 6) {real, imag} */,
  {32'hc5af0b0e, 32'h00000000} /* (11, 12, 5) {real, imag} */,
  {32'hc5afe23d, 32'h00000000} /* (11, 12, 4) {real, imag} */,
  {32'hc59abf8e, 32'h00000000} /* (11, 12, 3) {real, imag} */,
  {32'hc5a3ed4e, 32'h00000000} /* (11, 12, 2) {real, imag} */,
  {32'hc5a81d58, 32'h00000000} /* (11, 12, 1) {real, imag} */,
  {32'hc58e27ea, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'hc50a0a2a, 32'h00000000} /* (11, 11, 31) {real, imag} */,
  {32'hc514b917, 32'h00000000} /* (11, 11, 30) {real, imag} */,
  {32'hc4ed67c0, 32'h00000000} /* (11, 11, 29) {real, imag} */,
  {32'hc4965bfe, 32'h00000000} /* (11, 11, 28) {real, imag} */,
  {32'hc4a8b2b4, 32'h00000000} /* (11, 11, 27) {real, imag} */,
  {32'hc46fb04f, 32'h00000000} /* (11, 11, 26) {real, imag} */,
  {32'hc4c30edf, 32'h00000000} /* (11, 11, 25) {real, imag} */,
  {32'hc5186a4c, 32'h00000000} /* (11, 11, 24) {real, imag} */,
  {32'hc48759a5, 32'h00000000} /* (11, 11, 23) {real, imag} */,
  {32'hc1333600, 32'h00000000} /* (11, 11, 22) {real, imag} */,
  {32'h44772542, 32'h00000000} /* (11, 11, 21) {real, imag} */,
  {32'h450cf002, 32'h00000000} /* (11, 11, 20) {real, imag} */,
  {32'h45571908, 32'h00000000} /* (11, 11, 19) {real, imag} */,
  {32'h4548b2b4, 32'h00000000} /* (11, 11, 18) {real, imag} */,
  {32'h455ab4de, 32'h00000000} /* (11, 11, 17) {real, imag} */,
  {32'h45a49fc7, 32'h00000000} /* (11, 11, 16) {real, imag} */,
  {32'h4549c360, 32'h00000000} /* (11, 11, 15) {real, imag} */,
  {32'h452b0e55, 32'h00000000} /* (11, 11, 14) {real, imag} */,
  {32'h45251538, 32'h00000000} /* (11, 11, 13) {real, imag} */,
  {32'h4518f4a3, 32'h00000000} /* (11, 11, 12) {real, imag} */,
  {32'h43bbfc34, 32'h00000000} /* (11, 11, 11) {real, imag} */,
  {32'hc412c1c1, 32'h00000000} /* (11, 11, 10) {real, imag} */,
  {32'hc4a4305f, 32'h00000000} /* (11, 11, 9) {real, imag} */,
  {32'hc5217c88, 32'h00000000} /* (11, 11, 8) {real, imag} */,
  {32'hc53f4e46, 32'h00000000} /* (11, 11, 7) {real, imag} */,
  {32'hc522cec3, 32'h00000000} /* (11, 11, 6) {real, imag} */,
  {32'hc5077db6, 32'h00000000} /* (11, 11, 5) {real, imag} */,
  {32'hc544eef6, 32'h00000000} /* (11, 11, 4) {real, imag} */,
  {32'hc55c6514, 32'h00000000} /* (11, 11, 3) {real, imag} */,
  {32'hc513d5bc, 32'h00000000} /* (11, 11, 2) {real, imag} */,
  {32'hc506bf98, 32'h00000000} /* (11, 11, 1) {real, imag} */,
  {32'hc4c77184, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'h44da6bc0, 32'h00000000} /* (11, 10, 31) {real, imag} */,
  {32'h451bddac, 32'h00000000} /* (11, 10, 30) {real, imag} */,
  {32'h451c9a7c, 32'h00000000} /* (11, 10, 29) {real, imag} */,
  {32'h4541dc1c, 32'h00000000} /* (11, 10, 28) {real, imag} */,
  {32'h45507892, 32'h00000000} /* (11, 10, 27) {real, imag} */,
  {32'h4515524e, 32'h00000000} /* (11, 10, 26) {real, imag} */,
  {32'h453c418f, 32'h00000000} /* (11, 10, 25) {real, imag} */,
  {32'h4520dad0, 32'h00000000} /* (11, 10, 24) {real, imag} */,
  {32'h4535523a, 32'h00000000} /* (11, 10, 23) {real, imag} */,
  {32'h45737125, 32'h00000000} /* (11, 10, 22) {real, imag} */,
  {32'h457d2824, 32'h00000000} /* (11, 10, 21) {real, imag} */,
  {32'h4514463e, 32'h00000000} /* (11, 10, 20) {real, imag} */,
  {32'h446a2f82, 32'h00000000} /* (11, 10, 19) {real, imag} */,
  {32'h42f0a4ec, 32'h00000000} /* (11, 10, 18) {real, imag} */,
  {32'hc3820388, 32'h00000000} /* (11, 10, 17) {real, imag} */,
  {32'h43c1f070, 32'h00000000} /* (11, 10, 16) {real, imag} */,
  {32'h43071cd4, 32'h00000000} /* (11, 10, 15) {real, imag} */,
  {32'hc2a63c40, 32'h00000000} /* (11, 10, 14) {real, imag} */,
  {32'hc40f2f76, 32'h00000000} /* (11, 10, 13) {real, imag} */,
  {32'hc453edda, 32'h00000000} /* (11, 10, 12) {real, imag} */,
  {32'hc41012da, 32'h00000000} /* (11, 10, 11) {real, imag} */,
  {32'hc40a14d6, 32'h00000000} /* (11, 10, 10) {real, imag} */,
  {32'h4434dbfc, 32'h00000000} /* (11, 10, 9) {real, imag} */,
  {32'h42d17180, 32'h00000000} /* (11, 10, 8) {real, imag} */,
  {32'h44ccf674, 32'h00000000} /* (11, 10, 7) {real, imag} */,
  {32'h44cec7e6, 32'h00000000} /* (11, 10, 6) {real, imag} */,
  {32'h44abc2e8, 32'h00000000} /* (11, 10, 5) {real, imag} */,
  {32'h44c9f77e, 32'h00000000} /* (11, 10, 4) {real, imag} */,
  {32'h44153a12, 32'h00000000} /* (11, 10, 3) {real, imag} */,
  {32'h4420041c, 32'h00000000} /* (11, 10, 2) {real, imag} */,
  {32'h4502d4ab, 32'h00000000} /* (11, 10, 1) {real, imag} */,
  {32'h44d2dd98, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h45895dab, 32'h00000000} /* (11, 9, 31) {real, imag} */,
  {32'h45a7479c, 32'h00000000} /* (11, 9, 30) {real, imag} */,
  {32'h45d38281, 32'h00000000} /* (11, 9, 29) {real, imag} */,
  {32'h45d86aca, 32'h00000000} /* (11, 9, 28) {real, imag} */,
  {32'h45d411b6, 32'h00000000} /* (11, 9, 27) {real, imag} */,
  {32'h45ca6272, 32'h00000000} /* (11, 9, 26) {real, imag} */,
  {32'h45bf3e02, 32'h00000000} /* (11, 9, 25) {real, imag} */,
  {32'h45a7e85b, 32'h00000000} /* (11, 9, 24) {real, imag} */,
  {32'h45c38c58, 32'h00000000} /* (11, 9, 23) {real, imag} */,
  {32'h459b0f03, 32'h00000000} /* (11, 9, 22) {real, imag} */,
  {32'h45762e8a, 32'h00000000} /* (11, 9, 21) {real, imag} */,
  {32'h45043853, 32'h00000000} /* (11, 9, 20) {real, imag} */,
  {32'h43eb434c, 32'h00000000} /* (11, 9, 19) {real, imag} */,
  {32'hc3d8b748, 32'h00000000} /* (11, 9, 18) {real, imag} */,
  {32'hc4ad3a1c, 32'h00000000} /* (11, 9, 17) {real, imag} */,
  {32'hc52c0e66, 32'h00000000} /* (11, 9, 16) {real, imag} */,
  {32'hc5379bca, 32'h00000000} /* (11, 9, 15) {real, imag} */,
  {32'hc521da44, 32'h00000000} /* (11, 9, 14) {real, imag} */,
  {32'hc53a5442, 32'h00000000} /* (11, 9, 13) {real, imag} */,
  {32'hc53441d4, 32'h00000000} /* (11, 9, 12) {real, imag} */,
  {32'hc501b424, 32'h00000000} /* (11, 9, 11) {real, imag} */,
  {32'h41bed680, 32'h00000000} /* (11, 9, 10) {real, imag} */,
  {32'h44be3bf4, 32'h00000000} /* (11, 9, 9) {real, imag} */,
  {32'h4521e1fe, 32'h00000000} /* (11, 9, 8) {real, imag} */,
  {32'h45867b9a, 32'h00000000} /* (11, 9, 7) {real, imag} */,
  {32'h45789fc6, 32'h00000000} /* (11, 9, 6) {real, imag} */,
  {32'h454ed19e, 32'h00000000} /* (11, 9, 5) {real, imag} */,
  {32'h4585e5e0, 32'h00000000} /* (11, 9, 4) {real, imag} */,
  {32'h458bf383, 32'h00000000} /* (11, 9, 3) {real, imag} */,
  {32'h4581c3e0, 32'h00000000} /* (11, 9, 2) {real, imag} */,
  {32'h458862d0, 32'h00000000} /* (11, 9, 1) {real, imag} */,
  {32'h4590887b, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h45bc6cd6, 32'h00000000} /* (11, 8, 31) {real, imag} */,
  {32'h45e9e363, 32'h00000000} /* (11, 8, 30) {real, imag} */,
  {32'h45fffa6a, 32'h00000000} /* (11, 8, 29) {real, imag} */,
  {32'h460eccb6, 32'h00000000} /* (11, 8, 28) {real, imag} */,
  {32'h46187657, 32'h00000000} /* (11, 8, 27) {real, imag} */,
  {32'h46171ee6, 32'h00000000} /* (11, 8, 26) {real, imag} */,
  {32'h4604a276, 32'h00000000} /* (11, 8, 25) {real, imag} */,
  {32'h45eefa2b, 32'h00000000} /* (11, 8, 24) {real, imag} */,
  {32'h45fb81aa, 32'h00000000} /* (11, 8, 23) {real, imag} */,
  {32'h45d10338, 32'h00000000} /* (11, 8, 22) {real, imag} */,
  {32'h45829734, 32'h00000000} /* (11, 8, 21) {real, imag} */,
  {32'h45223ede, 32'h00000000} /* (11, 8, 20) {real, imag} */,
  {32'h44461184, 32'h00000000} /* (11, 8, 19) {real, imag} */,
  {32'hc4acdab4, 32'h00000000} /* (11, 8, 18) {real, imag} */,
  {32'hc536e0f6, 32'h00000000} /* (11, 8, 17) {real, imag} */,
  {32'hc55ba975, 32'h00000000} /* (11, 8, 16) {real, imag} */,
  {32'hc5979c44, 32'h00000000} /* (11, 8, 15) {real, imag} */,
  {32'hc584ccd7, 32'h00000000} /* (11, 8, 14) {real, imag} */,
  {32'hc5568584, 32'h00000000} /* (11, 8, 13) {real, imag} */,
  {32'hc56323a6, 32'h00000000} /* (11, 8, 12) {real, imag} */,
  {32'hc51ba5d9, 32'h00000000} /* (11, 8, 11) {real, imag} */,
  {32'hc3a9e090, 32'h00000000} /* (11, 8, 10) {real, imag} */,
  {32'h444881e0, 32'h00000000} /* (11, 8, 9) {real, imag} */,
  {32'h4573600a, 32'h00000000} /* (11, 8, 8) {real, imag} */,
  {32'h455b740c, 32'h00000000} /* (11, 8, 7) {real, imag} */,
  {32'h45913286, 32'h00000000} /* (11, 8, 6) {real, imag} */,
  {32'h45c01eb8, 32'h00000000} /* (11, 8, 5) {real, imag} */,
  {32'h45b4b1dd, 32'h00000000} /* (11, 8, 4) {real, imag} */,
  {32'h45c602c6, 32'h00000000} /* (11, 8, 3) {real, imag} */,
  {32'h45cff8e9, 32'h00000000} /* (11, 8, 2) {real, imag} */,
  {32'h45e17b6b, 32'h00000000} /* (11, 8, 1) {real, imag} */,
  {32'h45d3ac76, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h4609d990, 32'h00000000} /* (11, 7, 31) {real, imag} */,
  {32'h46094180, 32'h00000000} /* (11, 7, 30) {real, imag} */,
  {32'h4614f4c0, 32'h00000000} /* (11, 7, 29) {real, imag} */,
  {32'h461a9c14, 32'h00000000} /* (11, 7, 28) {real, imag} */,
  {32'h463094f6, 32'h00000000} /* (11, 7, 27) {real, imag} */,
  {32'h462c4a4c, 32'h00000000} /* (11, 7, 26) {real, imag} */,
  {32'h4621db82, 32'h00000000} /* (11, 7, 25) {real, imag} */,
  {32'h461a416e, 32'h00000000} /* (11, 7, 24) {real, imag} */,
  {32'h4607f676, 32'h00000000} /* (11, 7, 23) {real, imag} */,
  {32'h46000680, 32'h00000000} /* (11, 7, 22) {real, imag} */,
  {32'h45d4f98b, 32'h00000000} /* (11, 7, 21) {real, imag} */,
  {32'h45643ca4, 32'h00000000} /* (11, 7, 20) {real, imag} */,
  {32'h444f35d0, 32'h00000000} /* (11, 7, 19) {real, imag} */,
  {32'hc4b906d8, 32'h00000000} /* (11, 7, 18) {real, imag} */,
  {32'hc5174334, 32'h00000000} /* (11, 7, 17) {real, imag} */,
  {32'hc5841bea, 32'h00000000} /* (11, 7, 16) {real, imag} */,
  {32'hc596cc48, 32'h00000000} /* (11, 7, 15) {real, imag} */,
  {32'hc5a85bdc, 32'h00000000} /* (11, 7, 14) {real, imag} */,
  {32'hc5a0e982, 32'h00000000} /* (11, 7, 13) {real, imag} */,
  {32'hc59b295b, 32'h00000000} /* (11, 7, 12) {real, imag} */,
  {32'hc55a5968, 32'h00000000} /* (11, 7, 11) {real, imag} */,
  {32'hc4aebbb0, 32'h00000000} /* (11, 7, 10) {real, imag} */,
  {32'h44aae50c, 32'h00000000} /* (11, 7, 9) {real, imag} */,
  {32'h452dead0, 32'h00000000} /* (11, 7, 8) {real, imag} */,
  {32'h45ad446c, 32'h00000000} /* (11, 7, 7) {real, imag} */,
  {32'h45c66151, 32'h00000000} /* (11, 7, 6) {real, imag} */,
  {32'h45e0e37b, 32'h00000000} /* (11, 7, 5) {real, imag} */,
  {32'h45f06004, 32'h00000000} /* (11, 7, 4) {real, imag} */,
  {32'h460cda87, 32'h00000000} /* (11, 7, 3) {real, imag} */,
  {32'h460e08c3, 32'h00000000} /* (11, 7, 2) {real, imag} */,
  {32'h45f17e7e, 32'h00000000} /* (11, 7, 1) {real, imag} */,
  {32'h45f610d6, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'h46197056, 32'h00000000} /* (11, 6, 31) {real, imag} */,
  {32'h46226030, 32'h00000000} /* (11, 6, 30) {real, imag} */,
  {32'h4623d2b4, 32'h00000000} /* (11, 6, 29) {real, imag} */,
  {32'h46387c50, 32'h00000000} /* (11, 6, 28) {real, imag} */,
  {32'h463d3ba8, 32'h00000000} /* (11, 6, 27) {real, imag} */,
  {32'h4645c250, 32'h00000000} /* (11, 6, 26) {real, imag} */,
  {32'h462def8a, 32'h00000000} /* (11, 6, 25) {real, imag} */,
  {32'h462a884a, 32'h00000000} /* (11, 6, 24) {real, imag} */,
  {32'h4619434e, 32'h00000000} /* (11, 6, 23) {real, imag} */,
  {32'h4602662f, 32'h00000000} /* (11, 6, 22) {real, imag} */,
  {32'h45f4bdf6, 32'h00000000} /* (11, 6, 21) {real, imag} */,
  {32'h45831609, 32'h00000000} /* (11, 6, 20) {real, imag} */,
  {32'h45184bad, 32'h00000000} /* (11, 6, 19) {real, imag} */,
  {32'hc4cc1aec, 32'h00000000} /* (11, 6, 18) {real, imag} */,
  {32'hc5149175, 32'h00000000} /* (11, 6, 17) {real, imag} */,
  {32'hc575f5a2, 32'h00000000} /* (11, 6, 16) {real, imag} */,
  {32'hc5968282, 32'h00000000} /* (11, 6, 15) {real, imag} */,
  {32'hc5b8d724, 32'h00000000} /* (11, 6, 14) {real, imag} */,
  {32'hc5c3cab8, 32'h00000000} /* (11, 6, 13) {real, imag} */,
  {32'hc5d2db74, 32'h00000000} /* (11, 6, 12) {real, imag} */,
  {32'hc59dee95, 32'h00000000} /* (11, 6, 11) {real, imag} */,
  {32'hc51a6908, 32'h00000000} /* (11, 6, 10) {real, imag} */,
  {32'hc3530000, 32'h00000000} /* (11, 6, 9) {real, imag} */,
  {32'h456c63b2, 32'h00000000} /* (11, 6, 8) {real, imag} */,
  {32'h45a0e139, 32'h00000000} /* (11, 6, 7) {real, imag} */,
  {32'h45b427aa, 32'h00000000} /* (11, 6, 6) {real, imag} */,
  {32'h45c15442, 32'h00000000} /* (11, 6, 5) {real, imag} */,
  {32'h460800f0, 32'h00000000} /* (11, 6, 4) {real, imag} */,
  {32'h460d2d80, 32'h00000000} /* (11, 6, 3) {real, imag} */,
  {32'h4616dff6, 32'h00000000} /* (11, 6, 2) {real, imag} */,
  {32'h4623ae2f, 32'h00000000} /* (11, 6, 1) {real, imag} */,
  {32'h461a6c28, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'h4624fe68, 32'h00000000} /* (11, 5, 31) {real, imag} */,
  {32'h463230de, 32'h00000000} /* (11, 5, 30) {real, imag} */,
  {32'h46410ca8, 32'h00000000} /* (11, 5, 29) {real, imag} */,
  {32'h463f9c91, 32'h00000000} /* (11, 5, 28) {real, imag} */,
  {32'h465e64b5, 32'h00000000} /* (11, 5, 27) {real, imag} */,
  {32'h4650b9b2, 32'h00000000} /* (11, 5, 26) {real, imag} */,
  {32'h463bd93d, 32'h00000000} /* (11, 5, 25) {real, imag} */,
  {32'h46363bc2, 32'h00000000} /* (11, 5, 24) {real, imag} */,
  {32'h46361b1a, 32'h00000000} /* (11, 5, 23) {real, imag} */,
  {32'h462577fe, 32'h00000000} /* (11, 5, 22) {real, imag} */,
  {32'h45fb8aa4, 32'h00000000} /* (11, 5, 21) {real, imag} */,
  {32'h45bd6a05, 32'h00000000} /* (11, 5, 20) {real, imag} */,
  {32'h45a09224, 32'h00000000} /* (11, 5, 19) {real, imag} */,
  {32'h4545b6b8, 32'h00000000} /* (11, 5, 18) {real, imag} */,
  {32'hc31f9720, 32'h00000000} /* (11, 5, 17) {real, imag} */,
  {32'hc517e772, 32'h00000000} /* (11, 5, 16) {real, imag} */,
  {32'hc580ac82, 32'h00000000} /* (11, 5, 15) {real, imag} */,
  {32'hc5d33fab, 32'h00000000} /* (11, 5, 14) {real, imag} */,
  {32'hc5b8e830, 32'h00000000} /* (11, 5, 13) {real, imag} */,
  {32'hc5bf73ea, 32'h00000000} /* (11, 5, 12) {real, imag} */,
  {32'hc5cc3e06, 32'h00000000} /* (11, 5, 11) {real, imag} */,
  {32'hc565a25a, 32'h00000000} /* (11, 5, 10) {real, imag} */,
  {32'hc4ed7608, 32'h00000000} /* (11, 5, 9) {real, imag} */,
  {32'h442ce6a8, 32'h00000000} /* (11, 5, 8) {real, imag} */,
  {32'h44dd7640, 32'h00000000} /* (11, 5, 7) {real, imag} */,
  {32'h45269adc, 32'h00000000} /* (11, 5, 6) {real, imag} */,
  {32'h45a6b34c, 32'h00000000} /* (11, 5, 5) {real, imag} */,
  {32'h45f4b443, 32'h00000000} /* (11, 5, 4) {real, imag} */,
  {32'h461f550e, 32'h00000000} /* (11, 5, 3) {real, imag} */,
  {32'h462acf3d, 32'h00000000} /* (11, 5, 2) {real, imag} */,
  {32'h4636ac64, 32'h00000000} /* (11, 5, 1) {real, imag} */,
  {32'h46240ee4, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h462dbbed, 32'h00000000} /* (11, 4, 31) {real, imag} */,
  {32'h46434241, 32'h00000000} /* (11, 4, 30) {real, imag} */,
  {32'h464c521b, 32'h00000000} /* (11, 4, 29) {real, imag} */,
  {32'h464b9877, 32'h00000000} /* (11, 4, 28) {real, imag} */,
  {32'h46498a97, 32'h00000000} /* (11, 4, 27) {real, imag} */,
  {32'h46486719, 32'h00000000} /* (11, 4, 26) {real, imag} */,
  {32'h4657ca2c, 32'h00000000} /* (11, 4, 25) {real, imag} */,
  {32'h463d2b36, 32'h00000000} /* (11, 4, 24) {real, imag} */,
  {32'h464267f8, 32'h00000000} /* (11, 4, 23) {real, imag} */,
  {32'h463f982c, 32'h00000000} /* (11, 4, 22) {real, imag} */,
  {32'h4623ce8d, 32'h00000000} /* (11, 4, 21) {real, imag} */,
  {32'h460f1d1a, 32'h00000000} /* (11, 4, 20) {real, imag} */,
  {32'h45de1b8e, 32'h00000000} /* (11, 4, 19) {real, imag} */,
  {32'h459f893e, 32'h00000000} /* (11, 4, 18) {real, imag} */,
  {32'h45672314, 32'h00000000} /* (11, 4, 17) {real, imag} */,
  {32'h445232d0, 32'h00000000} /* (11, 4, 16) {real, imag} */,
  {32'hc5744cf1, 32'h00000000} /* (11, 4, 15) {real, imag} */,
  {32'hc5a2b82e, 32'h00000000} /* (11, 4, 14) {real, imag} */,
  {32'hc5bdef8a, 32'h00000000} /* (11, 4, 13) {real, imag} */,
  {32'hc5c04042, 32'h00000000} /* (11, 4, 12) {real, imag} */,
  {32'hc5d262ca, 32'h00000000} /* (11, 4, 11) {real, imag} */,
  {32'hc590b72e, 32'h00000000} /* (11, 4, 10) {real, imag} */,
  {32'hc56be1c0, 32'h00000000} /* (11, 4, 9) {real, imag} */,
  {32'hc55148ca, 32'h00000000} /* (11, 4, 8) {real, imag} */,
  {32'hc407c548, 32'h00000000} /* (11, 4, 7) {real, imag} */,
  {32'h450a58aa, 32'h00000000} /* (11, 4, 6) {real, imag} */,
  {32'h45a54926, 32'h00000000} /* (11, 4, 5) {real, imag} */,
  {32'h45f11478, 32'h00000000} /* (11, 4, 4) {real, imag} */,
  {32'h461fe9b3, 32'h00000000} /* (11, 4, 3) {real, imag} */,
  {32'h46291e5f, 32'h00000000} /* (11, 4, 2) {real, imag} */,
  {32'h462f3949, 32'h00000000} /* (11, 4, 1) {real, imag} */,
  {32'h462bb083, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h46385cd9, 32'h00000000} /* (11, 3, 31) {real, imag} */,
  {32'h4649e2ae, 32'h00000000} /* (11, 3, 30) {real, imag} */,
  {32'h4667d460, 32'h00000000} /* (11, 3, 29) {real, imag} */,
  {32'h465ee080, 32'h00000000} /* (11, 3, 28) {real, imag} */,
  {32'h4655d828, 32'h00000000} /* (11, 3, 27) {real, imag} */,
  {32'h46527077, 32'h00000000} /* (11, 3, 26) {real, imag} */,
  {32'h465592a4, 32'h00000000} /* (11, 3, 25) {real, imag} */,
  {32'h464b07a5, 32'h00000000} /* (11, 3, 24) {real, imag} */,
  {32'h463f7f7a, 32'h00000000} /* (11, 3, 23) {real, imag} */,
  {32'h4639f0b2, 32'h00000000} /* (11, 3, 22) {real, imag} */,
  {32'h462154b2, 32'h00000000} /* (11, 3, 21) {real, imag} */,
  {32'h46075114, 32'h00000000} /* (11, 3, 20) {real, imag} */,
  {32'h45ebca17, 32'h00000000} /* (11, 3, 19) {real, imag} */,
  {32'h45a448f8, 32'h00000000} /* (11, 3, 18) {real, imag} */,
  {32'h453f5372, 32'h00000000} /* (11, 3, 17) {real, imag} */,
  {32'h440afb30, 32'h00000000} /* (11, 3, 16) {real, imag} */,
  {32'hc5769c0b, 32'h00000000} /* (11, 3, 15) {real, imag} */,
  {32'hc59ed60b, 32'h00000000} /* (11, 3, 14) {real, imag} */,
  {32'hc5d81ad5, 32'h00000000} /* (11, 3, 13) {real, imag} */,
  {32'hc5d7027c, 32'h00000000} /* (11, 3, 12) {real, imag} */,
  {32'hc5c530a4, 32'h00000000} /* (11, 3, 11) {real, imag} */,
  {32'hc5bbb172, 32'h00000000} /* (11, 3, 10) {real, imag} */,
  {32'hc589246b, 32'h00000000} /* (11, 3, 9) {real, imag} */,
  {32'hc569f7ac, 32'h00000000} /* (11, 3, 8) {real, imag} */,
  {32'hc47caab8, 32'h00000000} /* (11, 3, 7) {real, imag} */,
  {32'h44186808, 32'h00000000} /* (11, 3, 6) {real, imag} */,
  {32'h45872839, 32'h00000000} /* (11, 3, 5) {real, imag} */,
  {32'h45f75a3b, 32'h00000000} /* (11, 3, 4) {real, imag} */,
  {32'h460be04e, 32'h00000000} /* (11, 3, 3) {real, imag} */,
  {32'h462b2afe, 32'h00000000} /* (11, 3, 2) {real, imag} */,
  {32'h4631bac4, 32'h00000000} /* (11, 3, 1) {real, imag} */,
  {32'h46300993, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'h464025d2, 32'h00000000} /* (11, 2, 31) {real, imag} */,
  {32'h464b076c, 32'h00000000} /* (11, 2, 30) {real, imag} */,
  {32'h465b5b5d, 32'h00000000} /* (11, 2, 29) {real, imag} */,
  {32'h4669953f, 32'h00000000} /* (11, 2, 28) {real, imag} */,
  {32'h4657fceb, 32'h00000000} /* (11, 2, 27) {real, imag} */,
  {32'h4651bb1b, 32'h00000000} /* (11, 2, 26) {real, imag} */,
  {32'h46506d99, 32'h00000000} /* (11, 2, 25) {real, imag} */,
  {32'h464d0326, 32'h00000000} /* (11, 2, 24) {real, imag} */,
  {32'h46496865, 32'h00000000} /* (11, 2, 23) {real, imag} */,
  {32'h4622d612, 32'h00000000} /* (11, 2, 22) {real, imag} */,
  {32'h461dbc03, 32'h00000000} /* (11, 2, 21) {real, imag} */,
  {32'h460e6253, 32'h00000000} /* (11, 2, 20) {real, imag} */,
  {32'h45e33ca7, 32'h00000000} /* (11, 2, 19) {real, imag} */,
  {32'h459a7424, 32'h00000000} /* (11, 2, 18) {real, imag} */,
  {32'h453a97e8, 32'h00000000} /* (11, 2, 17) {real, imag} */,
  {32'hc40fc010, 32'h00000000} /* (11, 2, 16) {real, imag} */,
  {32'hc5715aaa, 32'h00000000} /* (11, 2, 15) {real, imag} */,
  {32'hc5aebad4, 32'h00000000} /* (11, 2, 14) {real, imag} */,
  {32'hc5dbca1a, 32'h00000000} /* (11, 2, 13) {real, imag} */,
  {32'hc5d498b6, 32'h00000000} /* (11, 2, 12) {real, imag} */,
  {32'hc5c8512a, 32'h00000000} /* (11, 2, 11) {real, imag} */,
  {32'hc5b82cde, 32'h00000000} /* (11, 2, 10) {real, imag} */,
  {32'hc5892996, 32'h00000000} /* (11, 2, 9) {real, imag} */,
  {32'hc549b864, 32'h00000000} /* (11, 2, 8) {real, imag} */,
  {32'hc4af36d8, 32'h00000000} /* (11, 2, 7) {real, imag} */,
  {32'hc2f53640, 32'h00000000} /* (11, 2, 6) {real, imag} */,
  {32'h457e4b13, 32'h00000000} /* (11, 2, 5) {real, imag} */,
  {32'h460480c1, 32'h00000000} /* (11, 2, 4) {real, imag} */,
  {32'h4616ee44, 32'h00000000} /* (11, 2, 3) {real, imag} */,
  {32'h46331758, 32'h00000000} /* (11, 2, 2) {real, imag} */,
  {32'h46354080, 32'h00000000} /* (11, 2, 1) {real, imag} */,
  {32'h462fb550, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'h463a797f, 32'h00000000} /* (11, 1, 31) {real, imag} */,
  {32'h46515d8f, 32'h00000000} /* (11, 1, 30) {real, imag} */,
  {32'h465f4afa, 32'h00000000} /* (11, 1, 29) {real, imag} */,
  {32'h4666f005, 32'h00000000} /* (11, 1, 28) {real, imag} */,
  {32'h466883b5, 32'h00000000} /* (11, 1, 27) {real, imag} */,
  {32'h4659e048, 32'h00000000} /* (11, 1, 26) {real, imag} */,
  {32'h464bb670, 32'h00000000} /* (11, 1, 25) {real, imag} */,
  {32'h46500db5, 32'h00000000} /* (11, 1, 24) {real, imag} */,
  {32'h464218b5, 32'h00000000} /* (11, 1, 23) {real, imag} */,
  {32'h461ba59f, 32'h00000000} /* (11, 1, 22) {real, imag} */,
  {32'h460d0116, 32'h00000000} /* (11, 1, 21) {real, imag} */,
  {32'h4600f96a, 32'h00000000} /* (11, 1, 20) {real, imag} */,
  {32'h45bebc54, 32'h00000000} /* (11, 1, 19) {real, imag} */,
  {32'h4590fc99, 32'h00000000} /* (11, 1, 18) {real, imag} */,
  {32'h44ad69e8, 32'h00000000} /* (11, 1, 17) {real, imag} */,
  {32'hc42e66e0, 32'h00000000} /* (11, 1, 16) {real, imag} */,
  {32'hc57d262d, 32'h00000000} /* (11, 1, 15) {real, imag} */,
  {32'hc5a9f492, 32'h00000000} /* (11, 1, 14) {real, imag} */,
  {32'hc5c26955, 32'h00000000} /* (11, 1, 13) {real, imag} */,
  {32'hc5d7ccd6, 32'h00000000} /* (11, 1, 12) {real, imag} */,
  {32'hc5aca126, 32'h00000000} /* (11, 1, 11) {real, imag} */,
  {32'hc5938321, 32'h00000000} /* (11, 1, 10) {real, imag} */,
  {32'hc54c97be, 32'h00000000} /* (11, 1, 9) {real, imag} */,
  {32'hc4f58538, 32'h00000000} /* (11, 1, 8) {real, imag} */,
  {32'hc48179e8, 32'h00000000} /* (11, 1, 7) {real, imag} */,
  {32'h44e39fda, 32'h00000000} /* (11, 1, 6) {real, imag} */,
  {32'h45a90b5a, 32'h00000000} /* (11, 1, 5) {real, imag} */,
  {32'h45f8ed3b, 32'h00000000} /* (11, 1, 4) {real, imag} */,
  {32'h461429b4, 32'h00000000} /* (11, 1, 3) {real, imag} */,
  {32'h46218250, 32'h00000000} /* (11, 1, 2) {real, imag} */,
  {32'h46377665, 32'h00000000} /* (11, 1, 1) {real, imag} */,
  {32'h4639507a, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h4639222b, 32'h00000000} /* (11, 0, 31) {real, imag} */,
  {32'h46432ecb, 32'h00000000} /* (11, 0, 30) {real, imag} */,
  {32'h464f42c5, 32'h00000000} /* (11, 0, 29) {real, imag} */,
  {32'h465a04a4, 32'h00000000} /* (11, 0, 28) {real, imag} */,
  {32'h46607c24, 32'h00000000} /* (11, 0, 27) {real, imag} */,
  {32'h464d1426, 32'h00000000} /* (11, 0, 26) {real, imag} */,
  {32'h46484ad2, 32'h00000000} /* (11, 0, 25) {real, imag} */,
  {32'h463fd360, 32'h00000000} /* (11, 0, 24) {real, imag} */,
  {32'h462e6024, 32'h00000000} /* (11, 0, 23) {real, imag} */,
  {32'h461300dd, 32'h00000000} /* (11, 0, 22) {real, imag} */,
  {32'h45e8a0d2, 32'h00000000} /* (11, 0, 21) {real, imag} */,
  {32'h45a9339e, 32'h00000000} /* (11, 0, 20) {real, imag} */,
  {32'h45926cbe, 32'h00000000} /* (11, 0, 19) {real, imag} */,
  {32'h4521672e, 32'h00000000} /* (11, 0, 18) {real, imag} */,
  {32'h438ccb30, 32'h00000000} /* (11, 0, 17) {real, imag} */,
  {32'hc4c19e48, 32'h00000000} /* (11, 0, 16) {real, imag} */,
  {32'hc579ad60, 32'h00000000} /* (11, 0, 15) {real, imag} */,
  {32'hc5b35322, 32'h00000000} /* (11, 0, 14) {real, imag} */,
  {32'hc5b14072, 32'h00000000} /* (11, 0, 13) {real, imag} */,
  {32'hc5abb938, 32'h00000000} /* (11, 0, 12) {real, imag} */,
  {32'hc585553c, 32'h00000000} /* (11, 0, 11) {real, imag} */,
  {32'hc54029aa, 32'h00000000} /* (11, 0, 10) {real, imag} */,
  {32'hc4a6009c, 32'h00000000} /* (11, 0, 9) {real, imag} */,
  {32'hc3e7c250, 32'h00000000} /* (11, 0, 8) {real, imag} */,
  {32'h448e22d8, 32'h00000000} /* (11, 0, 7) {real, imag} */,
  {32'h455a13fd, 32'h00000000} /* (11, 0, 6) {real, imag} */,
  {32'h45c3cd66, 32'h00000000} /* (11, 0, 5) {real, imag} */,
  {32'h45f9a58a, 32'h00000000} /* (11, 0, 4) {real, imag} */,
  {32'h461867a1, 32'h00000000} /* (11, 0, 3) {real, imag} */,
  {32'h462952ac, 32'h00000000} /* (11, 0, 2) {real, imag} */,
  {32'h46370858, 32'h00000000} /* (11, 0, 1) {real, imag} */,
  {32'h46357e28, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h463cabe1, 32'h00000000} /* (10, 31, 31) {real, imag} */,
  {32'h4649481b, 32'h00000000} /* (10, 31, 30) {real, imag} */,
  {32'h4650a9b4, 32'h00000000} /* (10, 31, 29) {real, imag} */,
  {32'h46535b94, 32'h00000000} /* (10, 31, 28) {real, imag} */,
  {32'h4655098e, 32'h00000000} /* (10, 31, 27) {real, imag} */,
  {32'h4646d42e, 32'h00000000} /* (10, 31, 26) {real, imag} */,
  {32'h464c61e6, 32'h00000000} /* (10, 31, 25) {real, imag} */,
  {32'h4642e756, 32'h00000000} /* (10, 31, 24) {real, imag} */,
  {32'h4630d567, 32'h00000000} /* (10, 31, 23) {real, imag} */,
  {32'h461b2848, 32'h00000000} /* (10, 31, 22) {real, imag} */,
  {32'h45e08430, 32'h00000000} /* (10, 31, 21) {real, imag} */,
  {32'h45708f80, 32'h00000000} /* (10, 31, 20) {real, imag} */,
  {32'h44f1efd0, 32'h00000000} /* (10, 31, 19) {real, imag} */,
  {32'h43034ba0, 32'h00000000} /* (10, 31, 18) {real, imag} */,
  {32'hc4a1bb98, 32'h00000000} /* (10, 31, 17) {real, imag} */,
  {32'hc57bf1e8, 32'h00000000} /* (10, 31, 16) {real, imag} */,
  {32'hc5b765c2, 32'h00000000} /* (10, 31, 15) {real, imag} */,
  {32'hc5ba5b3a, 32'h00000000} /* (10, 31, 14) {real, imag} */,
  {32'hc5d2ca7c, 32'h00000000} /* (10, 31, 13) {real, imag} */,
  {32'hc5b1e778, 32'h00000000} /* (10, 31, 12) {real, imag} */,
  {32'hc560a126, 32'h00000000} /* (10, 31, 11) {real, imag} */,
  {32'hc4d96674, 32'h00000000} /* (10, 31, 10) {real, imag} */,
  {32'h44314b70, 32'h00000000} /* (10, 31, 9) {real, imag} */,
  {32'h452af38e, 32'h00000000} /* (10, 31, 8) {real, imag} */,
  {32'h458d02da, 32'h00000000} /* (10, 31, 7) {real, imag} */,
  {32'h45dcfffc, 32'h00000000} /* (10, 31, 6) {real, imag} */,
  {32'h45f1bddc, 32'h00000000} /* (10, 31, 5) {real, imag} */,
  {32'h4613c7e8, 32'h00000000} /* (10, 31, 4) {real, imag} */,
  {32'h46250841, 32'h00000000} /* (10, 31, 3) {real, imag} */,
  {32'h462caca2, 32'h00000000} /* (10, 31, 2) {real, imag} */,
  {32'h4644cf86, 32'h00000000} /* (10, 31, 1) {real, imag} */,
  {32'h4642461c, 32'h00000000} /* (10, 31, 0) {real, imag} */,
  {32'h464d5442, 32'h00000000} /* (10, 30, 31) {real, imag} */,
  {32'h465cd559, 32'h00000000} /* (10, 30, 30) {real, imag} */,
  {32'h46557a89, 32'h00000000} /* (10, 30, 29) {real, imag} */,
  {32'h4663151e, 32'h00000000} /* (10, 30, 28) {real, imag} */,
  {32'h4652a012, 32'h00000000} /* (10, 30, 27) {real, imag} */,
  {32'h464b5118, 32'h00000000} /* (10, 30, 26) {real, imag} */,
  {32'h464a513c, 32'h00000000} /* (10, 30, 25) {real, imag} */,
  {32'h4640b09c, 32'h00000000} /* (10, 30, 24) {real, imag} */,
  {32'h46250a33, 32'h00000000} /* (10, 30, 23) {real, imag} */,
  {32'h460d100f, 32'h00000000} /* (10, 30, 22) {real, imag} */,
  {32'h45b8500d, 32'h00000000} /* (10, 30, 21) {real, imag} */,
  {32'h4521e110, 32'h00000000} /* (10, 30, 20) {real, imag} */,
  {32'h42396a80, 32'h00000000} /* (10, 30, 19) {real, imag} */,
  {32'hc507f2fc, 32'h00000000} /* (10, 30, 18) {real, imag} */,
  {32'hc54828fa, 32'h00000000} /* (10, 30, 17) {real, imag} */,
  {32'hc5b5920b, 32'h00000000} /* (10, 30, 16) {real, imag} */,
  {32'hc5caffa9, 32'h00000000} /* (10, 30, 15) {real, imag} */,
  {32'hc5dd5386, 32'h00000000} /* (10, 30, 14) {real, imag} */,
  {32'hc5e2c65a, 32'h00000000} /* (10, 30, 13) {real, imag} */,
  {32'hc5bef4eb, 32'h00000000} /* (10, 30, 12) {real, imag} */,
  {32'hc534d300, 32'h00000000} /* (10, 30, 11) {real, imag} */,
  {32'hc373a000, 32'h00000000} /* (10, 30, 10) {real, imag} */,
  {32'h45263a98, 32'h00000000} /* (10, 30, 9) {real, imag} */,
  {32'h45bdb418, 32'h00000000} /* (10, 30, 8) {real, imag} */,
  {32'h45d2c52b, 32'h00000000} /* (10, 30, 7) {real, imag} */,
  {32'h45faee0a, 32'h00000000} /* (10, 30, 6) {real, imag} */,
  {32'h4619fd6e, 32'h00000000} /* (10, 30, 5) {real, imag} */,
  {32'h462e8727, 32'h00000000} /* (10, 30, 4) {real, imag} */,
  {32'h4634606e, 32'h00000000} /* (10, 30, 3) {real, imag} */,
  {32'h4644afa1, 32'h00000000} /* (10, 30, 2) {real, imag} */,
  {32'h464d6454, 32'h00000000} /* (10, 30, 1) {real, imag} */,
  {32'h463fde8c, 32'h00000000} /* (10, 30, 0) {real, imag} */,
  {32'h4652b0a6, 32'h00000000} /* (10, 29, 31) {real, imag} */,
  {32'h465e644a, 32'h00000000} /* (10, 29, 30) {real, imag} */,
  {32'h4656fca3, 32'h00000000} /* (10, 29, 29) {real, imag} */,
  {32'h46539aeb, 32'h00000000} /* (10, 29, 28) {real, imag} */,
  {32'h46573edd, 32'h00000000} /* (10, 29, 27) {real, imag} */,
  {32'h465bf123, 32'h00000000} /* (10, 29, 26) {real, imag} */,
  {32'h46453827, 32'h00000000} /* (10, 29, 25) {real, imag} */,
  {32'h4634747e, 32'h00000000} /* (10, 29, 24) {real, imag} */,
  {32'h461e172a, 32'h00000000} /* (10, 29, 23) {real, imag} */,
  {32'h45f3ce34, 32'h00000000} /* (10, 29, 22) {real, imag} */,
  {32'h459fea0d, 32'h00000000} /* (10, 29, 21) {real, imag} */,
  {32'h446af208, 32'h00000000} /* (10, 29, 20) {real, imag} */,
  {32'hc4cd3b28, 32'h00000000} /* (10, 29, 19) {real, imag} */,
  {32'hc580730e, 32'h00000000} /* (10, 29, 18) {real, imag} */,
  {32'hc59ec090, 32'h00000000} /* (10, 29, 17) {real, imag} */,
  {32'hc5bb81b7, 32'h00000000} /* (10, 29, 16) {real, imag} */,
  {32'hc5eb7a37, 32'h00000000} /* (10, 29, 15) {real, imag} */,
  {32'hc5d8997b, 32'h00000000} /* (10, 29, 14) {real, imag} */,
  {32'hc5c3ad46, 32'h00000000} /* (10, 29, 13) {real, imag} */,
  {32'hc59e209e, 32'h00000000} /* (10, 29, 12) {real, imag} */,
  {32'hc5453b74, 32'h00000000} /* (10, 29, 11) {real, imag} */,
  {32'h44b39b78, 32'h00000000} /* (10, 29, 10) {real, imag} */,
  {32'h456c9684, 32'h00000000} /* (10, 29, 9) {real, imag} */,
  {32'h45cb0053, 32'h00000000} /* (10, 29, 8) {real, imag} */,
  {32'h460496ce, 32'h00000000} /* (10, 29, 7) {real, imag} */,
  {32'h460def46, 32'h00000000} /* (10, 29, 6) {real, imag} */,
  {32'h4625f44e, 32'h00000000} /* (10, 29, 5) {real, imag} */,
  {32'h463d1ff4, 32'h00000000} /* (10, 29, 4) {real, imag} */,
  {32'h464a72b3, 32'h00000000} /* (10, 29, 3) {real, imag} */,
  {32'h46447e61, 32'h00000000} /* (10, 29, 2) {real, imag} */,
  {32'h464d5ad4, 32'h00000000} /* (10, 29, 1) {real, imag} */,
  {32'h464d3354, 32'h00000000} /* (10, 29, 0) {real, imag} */,
  {32'h4650a966, 32'h00000000} /* (10, 28, 31) {real, imag} */,
  {32'h46561250, 32'h00000000} /* (10, 28, 30) {real, imag} */,
  {32'h46516c0a, 32'h00000000} /* (10, 28, 29) {real, imag} */,
  {32'h4656f3fe, 32'h00000000} /* (10, 28, 28) {real, imag} */,
  {32'h46586c87, 32'h00000000} /* (10, 28, 27) {real, imag} */,
  {32'h46545e32, 32'h00000000} /* (10, 28, 26) {real, imag} */,
  {32'h46435cb2, 32'h00000000} /* (10, 28, 25) {real, imag} */,
  {32'h46441a77, 32'h00000000} /* (10, 28, 24) {real, imag} */,
  {32'h461e23cc, 32'h00000000} /* (10, 28, 23) {real, imag} */,
  {32'h45f5350c, 32'h00000000} /* (10, 28, 22) {real, imag} */,
  {32'h456ebaf8, 32'h00000000} /* (10, 28, 21) {real, imag} */,
  {32'h4396aa90, 32'h00000000} /* (10, 28, 20) {real, imag} */,
  {32'hc539fbbe, 32'h00000000} /* (10, 28, 19) {real, imag} */,
  {32'hc5a5454b, 32'h00000000} /* (10, 28, 18) {real, imag} */,
  {32'hc5bd595e, 32'h00000000} /* (10, 28, 17) {real, imag} */,
  {32'hc5ed2d50, 32'h00000000} /* (10, 28, 16) {real, imag} */,
  {32'hc60682a4, 32'h00000000} /* (10, 28, 15) {real, imag} */,
  {32'hc5ed3911, 32'h00000000} /* (10, 28, 14) {real, imag} */,
  {32'hc5c318c9, 32'h00000000} /* (10, 28, 13) {real, imag} */,
  {32'hc5a71200, 32'h00000000} /* (10, 28, 12) {real, imag} */,
  {32'hc4f864c8, 32'h00000000} /* (10, 28, 11) {real, imag} */,
  {32'h44a4672c, 32'h00000000} /* (10, 28, 10) {real, imag} */,
  {32'h458e406b, 32'h00000000} /* (10, 28, 9) {real, imag} */,
  {32'h45bea9b6, 32'h00000000} /* (10, 28, 8) {real, imag} */,
  {32'h460d51f6, 32'h00000000} /* (10, 28, 7) {real, imag} */,
  {32'h46289292, 32'h00000000} /* (10, 28, 6) {real, imag} */,
  {32'h463576ed, 32'h00000000} /* (10, 28, 5) {real, imag} */,
  {32'h46516016, 32'h00000000} /* (10, 28, 4) {real, imag} */,
  {32'h464aff92, 32'h00000000} /* (10, 28, 3) {real, imag} */,
  {32'h4644c6ba, 32'h00000000} /* (10, 28, 2) {real, imag} */,
  {32'h4659377b, 32'h00000000} /* (10, 28, 1) {real, imag} */,
  {32'h464cf8ea, 32'h00000000} /* (10, 28, 0) {real, imag} */,
  {32'h464b8c3d, 32'h00000000} /* (10, 27, 31) {real, imag} */,
  {32'h4653c28a, 32'h00000000} /* (10, 27, 30) {real, imag} */,
  {32'h4668e3e8, 32'h00000000} /* (10, 27, 29) {real, imag} */,
  {32'h46527b3e, 32'h00000000} /* (10, 27, 28) {real, imag} */,
  {32'h466a48ee, 32'h00000000} /* (10, 27, 27) {real, imag} */,
  {32'h4662019c, 32'h00000000} /* (10, 27, 26) {real, imag} */,
  {32'h4642a012, 32'h00000000} /* (10, 27, 25) {real, imag} */,
  {32'h4640e1f1, 32'h00000000} /* (10, 27, 24) {real, imag} */,
  {32'h46234c97, 32'h00000000} /* (10, 27, 23) {real, imag} */,
  {32'h45eed403, 32'h00000000} /* (10, 27, 22) {real, imag} */,
  {32'h45376c48, 32'h00000000} /* (10, 27, 21) {real, imag} */,
  {32'hc474d790, 32'h00000000} /* (10, 27, 20) {real, imag} */,
  {32'hc584015a, 32'h00000000} /* (10, 27, 19) {real, imag} */,
  {32'hc5b8171e, 32'h00000000} /* (10, 27, 18) {real, imag} */,
  {32'hc5fcbef3, 32'h00000000} /* (10, 27, 17) {real, imag} */,
  {32'hc60cb4ce, 32'h00000000} /* (10, 27, 16) {real, imag} */,
  {32'hc60897ff, 32'h00000000} /* (10, 27, 15) {real, imag} */,
  {32'hc6019b46, 32'h00000000} /* (10, 27, 14) {real, imag} */,
  {32'hc5cd6741, 32'h00000000} /* (10, 27, 13) {real, imag} */,
  {32'hc5828137, 32'h00000000} /* (10, 27, 12) {real, imag} */,
  {32'hc51be8c8, 32'h00000000} /* (10, 27, 11) {real, imag} */,
  {32'h44a12f60, 32'h00000000} /* (10, 27, 10) {real, imag} */,
  {32'h45aa97cc, 32'h00000000} /* (10, 27, 9) {real, imag} */,
  {32'h45d8e926, 32'h00000000} /* (10, 27, 8) {real, imag} */,
  {32'h460e99f1, 32'h00000000} /* (10, 27, 7) {real, imag} */,
  {32'h46243526, 32'h00000000} /* (10, 27, 6) {real, imag} */,
  {32'h4645bef3, 32'h00000000} /* (10, 27, 5) {real, imag} */,
  {32'h46558bc2, 32'h00000000} /* (10, 27, 4) {real, imag} */,
  {32'h464578af, 32'h00000000} /* (10, 27, 3) {real, imag} */,
  {32'h4648e853, 32'h00000000} /* (10, 27, 2) {real, imag} */,
  {32'h464ce1ca, 32'h00000000} /* (10, 27, 1) {real, imag} */,
  {32'h46520310, 32'h00000000} /* (10, 27, 0) {real, imag} */,
  {32'h463b3a6a, 32'h00000000} /* (10, 26, 31) {real, imag} */,
  {32'h46470cdf, 32'h00000000} /* (10, 26, 30) {real, imag} */,
  {32'h46600031, 32'h00000000} /* (10, 26, 29) {real, imag} */,
  {32'h4643919e, 32'h00000000} /* (10, 26, 28) {real, imag} */,
  {32'h464e33e7, 32'h00000000} /* (10, 26, 27) {real, imag} */,
  {32'h4642d4c0, 32'h00000000} /* (10, 26, 26) {real, imag} */,
  {32'h464b074e, 32'h00000000} /* (10, 26, 25) {real, imag} */,
  {32'h46327bb1, 32'h00000000} /* (10, 26, 24) {real, imag} */,
  {32'h45fa8389, 32'h00000000} /* (10, 26, 23) {real, imag} */,
  {32'h45cd7c42, 32'h00000000} /* (10, 26, 22) {real, imag} */,
  {32'h45171f06, 32'h00000000} /* (10, 26, 21) {real, imag} */,
  {32'hc4dbfd0c, 32'h00000000} /* (10, 26, 20) {real, imag} */,
  {32'hc58b0bd7, 32'h00000000} /* (10, 26, 19) {real, imag} */,
  {32'hc5c2b9fe, 32'h00000000} /* (10, 26, 18) {real, imag} */,
  {32'hc603070f, 32'h00000000} /* (10, 26, 17) {real, imag} */,
  {32'hc6112f39, 32'h00000000} /* (10, 26, 16) {real, imag} */,
  {32'hc5fc5800, 32'h00000000} /* (10, 26, 15) {real, imag} */,
  {32'hc5d562fa, 32'h00000000} /* (10, 26, 14) {real, imag} */,
  {32'hc5c794ea, 32'h00000000} /* (10, 26, 13) {real, imag} */,
  {32'hc596c417, 32'h00000000} /* (10, 26, 12) {real, imag} */,
  {32'hc4b335f0, 32'h00000000} /* (10, 26, 11) {real, imag} */,
  {32'h4500c5ae, 32'h00000000} /* (10, 26, 10) {real, imag} */,
  {32'h45cb65b4, 32'h00000000} /* (10, 26, 9) {real, imag} */,
  {32'h45fe35aa, 32'h00000000} /* (10, 26, 8) {real, imag} */,
  {32'h46206296, 32'h00000000} /* (10, 26, 7) {real, imag} */,
  {32'h4623bf15, 32'h00000000} /* (10, 26, 6) {real, imag} */,
  {32'h46384ab2, 32'h00000000} /* (10, 26, 5) {real, imag} */,
  {32'h463b3016, 32'h00000000} /* (10, 26, 4) {real, imag} */,
  {32'h46431526, 32'h00000000} /* (10, 26, 3) {real, imag} */,
  {32'h4651c197, 32'h00000000} /* (10, 26, 2) {real, imag} */,
  {32'h463f26cf, 32'h00000000} /* (10, 26, 1) {real, imag} */,
  {32'h4641d7bf, 32'h00000000} /* (10, 26, 0) {real, imag} */,
  {32'h4630a237, 32'h00000000} /* (10, 25, 31) {real, imag} */,
  {32'h462badc4, 32'h00000000} /* (10, 25, 30) {real, imag} */,
  {32'h463d72b2, 32'h00000000} /* (10, 25, 29) {real, imag} */,
  {32'h463d7084, 32'h00000000} /* (10, 25, 28) {real, imag} */,
  {32'h462d5995, 32'h00000000} /* (10, 25, 27) {real, imag} */,
  {32'h462b6b3a, 32'h00000000} /* (10, 25, 26) {real, imag} */,
  {32'h46354d02, 32'h00000000} /* (10, 25, 25) {real, imag} */,
  {32'h4616932a, 32'h00000000} /* (10, 25, 24) {real, imag} */,
  {32'h45e11ec4, 32'h00000000} /* (10, 25, 23) {real, imag} */,
  {32'h45a8a723, 32'h00000000} /* (10, 25, 22) {real, imag} */,
  {32'h4509a3ea, 32'h00000000} /* (10, 25, 21) {real, imag} */,
  {32'hc4714988, 32'h00000000} /* (10, 25, 20) {real, imag} */,
  {32'hc58adeec, 32'h00000000} /* (10, 25, 19) {real, imag} */,
  {32'hc5bcfd8b, 32'h00000000} /* (10, 25, 18) {real, imag} */,
  {32'hc60285ee, 32'h00000000} /* (10, 25, 17) {real, imag} */,
  {32'hc60269c3, 32'h00000000} /* (10, 25, 16) {real, imag} */,
  {32'hc5e8c3c2, 32'h00000000} /* (10, 25, 15) {real, imag} */,
  {32'hc5e13481, 32'h00000000} /* (10, 25, 14) {real, imag} */,
  {32'hc5b1bcd7, 32'h00000000} /* (10, 25, 13) {real, imag} */,
  {32'hc57c711e, 32'h00000000} /* (10, 25, 12) {real, imag} */,
  {32'hc4799c40, 32'h00000000} /* (10, 25, 11) {real, imag} */,
  {32'h4519cb86, 32'h00000000} /* (10, 25, 10) {real, imag} */,
  {32'h45b63418, 32'h00000000} /* (10, 25, 9) {real, imag} */,
  {32'h46037aee, 32'h00000000} /* (10, 25, 8) {real, imag} */,
  {32'h4615c29c, 32'h00000000} /* (10, 25, 7) {real, imag} */,
  {32'h4628b1a4, 32'h00000000} /* (10, 25, 6) {real, imag} */,
  {32'h46390166, 32'h00000000} /* (10, 25, 5) {real, imag} */,
  {32'h463b344a, 32'h00000000} /* (10, 25, 4) {real, imag} */,
  {32'h46327eb0, 32'h00000000} /* (10, 25, 3) {real, imag} */,
  {32'h463380da, 32'h00000000} /* (10, 25, 2) {real, imag} */,
  {32'h46327928, 32'h00000000} /* (10, 25, 1) {real, imag} */,
  {32'h4625f0a5, 32'h00000000} /* (10, 25, 0) {real, imag} */,
  {32'h460c2b5f, 32'h00000000} /* (10, 24, 31) {real, imag} */,
  {32'h46176f4f, 32'h00000000} /* (10, 24, 30) {real, imag} */,
  {32'h46248bc4, 32'h00000000} /* (10, 24, 29) {real, imag} */,
  {32'h4629f066, 32'h00000000} /* (10, 24, 28) {real, imag} */,
  {32'h46278da2, 32'h00000000} /* (10, 24, 27) {real, imag} */,
  {32'h4617855c, 32'h00000000} /* (10, 24, 26) {real, imag} */,
  {32'h461082ff, 32'h00000000} /* (10, 24, 25) {real, imag} */,
  {32'h45f58d0a, 32'h00000000} /* (10, 24, 24) {real, imag} */,
  {32'h45c770d2, 32'h00000000} /* (10, 24, 23) {real, imag} */,
  {32'h458492ab, 32'h00000000} /* (10, 24, 22) {real, imag} */,
  {32'h44af9bc4, 32'h00000000} /* (10, 24, 21) {real, imag} */,
  {32'hc53ba192, 32'h00000000} /* (10, 24, 20) {real, imag} */,
  {32'hc584c538, 32'h00000000} /* (10, 24, 19) {real, imag} */,
  {32'hc5a51d53, 32'h00000000} /* (10, 24, 18) {real, imag} */,
  {32'hc5d1f5b5, 32'h00000000} /* (10, 24, 17) {real, imag} */,
  {32'hc5cfac0e, 32'h00000000} /* (10, 24, 16) {real, imag} */,
  {32'hc5ca10e8, 32'h00000000} /* (10, 24, 15) {real, imag} */,
  {32'hc5bc7120, 32'h00000000} /* (10, 24, 14) {real, imag} */,
  {32'hc5944263, 32'h00000000} /* (10, 24, 13) {real, imag} */,
  {32'hc5875936, 32'h00000000} /* (10, 24, 12) {real, imag} */,
  {32'hc5035ef8, 32'h00000000} /* (10, 24, 11) {real, imag} */,
  {32'h452cf24a, 32'h00000000} /* (10, 24, 10) {real, imag} */,
  {32'h45a7ec3c, 32'h00000000} /* (10, 24, 9) {real, imag} */,
  {32'h45ed226e, 32'h00000000} /* (10, 24, 8) {real, imag} */,
  {32'h4612d3df, 32'h00000000} /* (10, 24, 7) {real, imag} */,
  {32'h46182552, 32'h00000000} /* (10, 24, 6) {real, imag} */,
  {32'h4616c9be, 32'h00000000} /* (10, 24, 5) {real, imag} */,
  {32'h461d2c34, 32'h00000000} /* (10, 24, 4) {real, imag} */,
  {32'h4621ed0e, 32'h00000000} /* (10, 24, 3) {real, imag} */,
  {32'h4634d2cc, 32'h00000000} /* (10, 24, 2) {real, imag} */,
  {32'h46160b1c, 32'h00000000} /* (10, 24, 1) {real, imag} */,
  {32'h461e0099, 32'h00000000} /* (10, 24, 0) {real, imag} */,
  {32'h45d81136, 32'h00000000} /* (10, 23, 31) {real, imag} */,
  {32'h45e85d38, 32'h00000000} /* (10, 23, 30) {real, imag} */,
  {32'h46011c58, 32'h00000000} /* (10, 23, 29) {real, imag} */,
  {32'h4601d513, 32'h00000000} /* (10, 23, 28) {real, imag} */,
  {32'h45f9a6f2, 32'h00000000} /* (10, 23, 27) {real, imag} */,
  {32'h45f9b426, 32'h00000000} /* (10, 23, 26) {real, imag} */,
  {32'h45e4f504, 32'h00000000} /* (10, 23, 25) {real, imag} */,
  {32'h45d1ddb6, 32'h00000000} /* (10, 23, 24) {real, imag} */,
  {32'h4583f906, 32'h00000000} /* (10, 23, 23) {real, imag} */,
  {32'h4564c360, 32'h00000000} /* (10, 23, 22) {real, imag} */,
  {32'h44b52544, 32'h00000000} /* (10, 23, 21) {real, imag} */,
  {32'hc54d9b76, 32'h00000000} /* (10, 23, 20) {real, imag} */,
  {32'hc58faef0, 32'h00000000} /* (10, 23, 19) {real, imag} */,
  {32'hc5b0e6c4, 32'h00000000} /* (10, 23, 18) {real, imag} */,
  {32'hc5b602bb, 32'h00000000} /* (10, 23, 17) {real, imag} */,
  {32'hc595a394, 32'h00000000} /* (10, 23, 16) {real, imag} */,
  {32'hc58cc084, 32'h00000000} /* (10, 23, 15) {real, imag} */,
  {32'hc57c72c3, 32'h00000000} /* (10, 23, 14) {real, imag} */,
  {32'hc5756122, 32'h00000000} /* (10, 23, 13) {real, imag} */,
  {32'hc561a618, 32'h00000000} /* (10, 23, 12) {real, imag} */,
  {32'hc502d7cb, 32'h00000000} /* (10, 23, 11) {real, imag} */,
  {32'h44e65a50, 32'h00000000} /* (10, 23, 10) {real, imag} */,
  {32'h45ab2bda, 32'h00000000} /* (10, 23, 9) {real, imag} */,
  {32'h45c24d16, 32'h00000000} /* (10, 23, 8) {real, imag} */,
  {32'h45f1e8de, 32'h00000000} /* (10, 23, 7) {real, imag} */,
  {32'h4606b02e, 32'h00000000} /* (10, 23, 6) {real, imag} */,
  {32'h45eda0f3, 32'h00000000} /* (10, 23, 5) {real, imag} */,
  {32'h46026714, 32'h00000000} /* (10, 23, 4) {real, imag} */,
  {32'h460b5392, 32'h00000000} /* (10, 23, 3) {real, imag} */,
  {32'h46018cd4, 32'h00000000} /* (10, 23, 2) {real, imag} */,
  {32'h46067ad8, 32'h00000000} /* (10, 23, 1) {real, imag} */,
  {32'h45eb20f2, 32'h00000000} /* (10, 23, 0) {real, imag} */,
  {32'h45975daa, 32'h00000000} /* (10, 22, 31) {real, imag} */,
  {32'h45b1e8f7, 32'h00000000} /* (10, 22, 30) {real, imag} */,
  {32'h45a2dcad, 32'h00000000} /* (10, 22, 29) {real, imag} */,
  {32'h45b72082, 32'h00000000} /* (10, 22, 28) {real, imag} */,
  {32'h459f0b38, 32'h00000000} /* (10, 22, 27) {real, imag} */,
  {32'h45b31b11, 32'h00000000} /* (10, 22, 26) {real, imag} */,
  {32'h45ab4640, 32'h00000000} /* (10, 22, 25) {real, imag} */,
  {32'h4583a076, 32'h00000000} /* (10, 22, 24) {real, imag} */,
  {32'h45552b11, 32'h00000000} /* (10, 22, 23) {real, imag} */,
  {32'h4513aae7, 32'h00000000} /* (10, 22, 22) {real, imag} */,
  {32'h447d3e74, 32'h00000000} /* (10, 22, 21) {real, imag} */,
  {32'hc4fcec44, 32'h00000000} /* (10, 22, 20) {real, imag} */,
  {32'hc57a274b, 32'h00000000} /* (10, 22, 19) {real, imag} */,
  {32'hc56691fe, 32'h00000000} /* (10, 22, 18) {real, imag} */,
  {32'hc55764ce, 32'h00000000} /* (10, 22, 17) {real, imag} */,
  {32'hc542691e, 32'h00000000} /* (10, 22, 16) {real, imag} */,
  {32'hc53fc254, 32'h00000000} /* (10, 22, 15) {real, imag} */,
  {32'hc577db86, 32'h00000000} /* (10, 22, 14) {real, imag} */,
  {32'hc56ed522, 32'h00000000} /* (10, 22, 13) {real, imag} */,
  {32'hc4c35562, 32'h00000000} /* (10, 22, 12) {real, imag} */,
  {32'hc458a388, 32'h00000000} /* (10, 22, 11) {real, imag} */,
  {32'h448c0704, 32'h00000000} /* (10, 22, 10) {real, imag} */,
  {32'h451bbe1d, 32'h00000000} /* (10, 22, 9) {real, imag} */,
  {32'h455c1960, 32'h00000000} /* (10, 22, 8) {real, imag} */,
  {32'h45958da4, 32'h00000000} /* (10, 22, 7) {real, imag} */,
  {32'h45a87dd6, 32'h00000000} /* (10, 22, 6) {real, imag} */,
  {32'h45b03a40, 32'h00000000} /* (10, 22, 5) {real, imag} */,
  {32'h45a7ad75, 32'h00000000} /* (10, 22, 4) {real, imag} */,
  {32'h45bd4ff4, 32'h00000000} /* (10, 22, 3) {real, imag} */,
  {32'h45d9c58b, 32'h00000000} /* (10, 22, 2) {real, imag} */,
  {32'h45a77493, 32'h00000000} /* (10, 22, 1) {real, imag} */,
  {32'h459fac17, 32'h00000000} /* (10, 22, 0) {real, imag} */,
  {32'h44a96038, 32'h00000000} /* (10, 21, 31) {real, imag} */,
  {32'h4525b8c4, 32'h00000000} /* (10, 21, 30) {real, imag} */,
  {32'h45004cad, 32'h00000000} /* (10, 21, 29) {real, imag} */,
  {32'h44c587a3, 32'h00000000} /* (10, 21, 28) {real, imag} */,
  {32'h450c92a4, 32'h00000000} /* (10, 21, 27) {real, imag} */,
  {32'h45012a3c, 32'h00000000} /* (10, 21, 26) {real, imag} */,
  {32'h44ab8202, 32'h00000000} /* (10, 21, 25) {real, imag} */,
  {32'h44ae82a6, 32'h00000000} /* (10, 21, 24) {real, imag} */,
  {32'h44c90966, 32'h00000000} /* (10, 21, 23) {real, imag} */,
  {32'h44cd7aaa, 32'h00000000} /* (10, 21, 22) {real, imag} */,
  {32'h4496095a, 32'h00000000} /* (10, 21, 21) {real, imag} */,
  {32'hc46452e0, 32'h00000000} /* (10, 21, 20) {real, imag} */,
  {32'hc4bdec5c, 32'h00000000} /* (10, 21, 19) {real, imag} */,
  {32'hc424db4e, 32'h00000000} /* (10, 21, 18) {real, imag} */,
  {32'hc41f7753, 32'h00000000} /* (10, 21, 17) {real, imag} */,
  {32'hc2748b30, 32'h00000000} /* (10, 21, 16) {real, imag} */,
  {32'h43242abc, 32'h00000000} /* (10, 21, 15) {real, imag} */,
  {32'hc4909480, 32'h00000000} /* (10, 21, 14) {real, imag} */,
  {32'hc408ba5c, 32'h00000000} /* (10, 21, 13) {real, imag} */,
  {32'hc3db67f8, 32'h00000000} /* (10, 21, 12) {real, imag} */,
  {32'h42889cc0, 32'h00000000} /* (10, 21, 11) {real, imag} */,
  {32'h43d7cdcc, 32'h00000000} /* (10, 21, 10) {real, imag} */,
  {32'h44962efa, 32'h00000000} /* (10, 21, 9) {real, imag} */,
  {32'h449466ea, 32'h00000000} /* (10, 21, 8) {real, imag} */,
  {32'h447d0804, 32'h00000000} /* (10, 21, 7) {real, imag} */,
  {32'h44abde9e, 32'h00000000} /* (10, 21, 6) {real, imag} */,
  {32'h450812e3, 32'h00000000} /* (10, 21, 5) {real, imag} */,
  {32'h44d1a714, 32'h00000000} /* (10, 21, 4) {real, imag} */,
  {32'h44eddc92, 32'h00000000} /* (10, 21, 3) {real, imag} */,
  {32'h450df27a, 32'h00000000} /* (10, 21, 2) {real, imag} */,
  {32'h44e41162, 32'h00000000} /* (10, 21, 1) {real, imag} */,
  {32'h4502d719, 32'h00000000} /* (10, 21, 0) {real, imag} */,
  {32'hc4cd39a8, 32'h00000000} /* (10, 20, 31) {real, imag} */,
  {32'hc513200f, 32'h00000000} /* (10, 20, 30) {real, imag} */,
  {32'hc4df8a36, 32'h00000000} /* (10, 20, 29) {real, imag} */,
  {32'hc4dd5600, 32'h00000000} /* (10, 20, 28) {real, imag} */,
  {32'hc4cf9c02, 32'h00000000} /* (10, 20, 27) {real, imag} */,
  {32'hc4dee636, 32'h00000000} /* (10, 20, 26) {real, imag} */,
  {32'hc51898c4, 32'h00000000} /* (10, 20, 25) {real, imag} */,
  {32'hc527e416, 32'h00000000} /* (10, 20, 24) {real, imag} */,
  {32'hc50743cf, 32'h00000000} /* (10, 20, 23) {real, imag} */,
  {32'hc4c0f3bb, 32'h00000000} /* (10, 20, 22) {real, imag} */,
  {32'h42e41f20, 32'h00000000} /* (10, 20, 21) {real, imag} */,
  {32'h44a6d2d6, 32'h00000000} /* (10, 20, 20) {real, imag} */,
  {32'h450b04ac, 32'h00000000} /* (10, 20, 19) {real, imag} */,
  {32'h44c62fce, 32'h00000000} /* (10, 20, 18) {real, imag} */,
  {32'h44f6ae1a, 32'h00000000} /* (10, 20, 17) {real, imag} */,
  {32'h456239ef, 32'h00000000} /* (10, 20, 16) {real, imag} */,
  {32'h45682f46, 32'h00000000} /* (10, 20, 15) {real, imag} */,
  {32'h455fee9f, 32'h00000000} /* (10, 20, 14) {real, imag} */,
  {32'h4541933f, 32'h00000000} /* (10, 20, 13) {real, imag} */,
  {32'h44fc7228, 32'h00000000} /* (10, 20, 12) {real, imag} */,
  {32'h44b394b4, 32'h00000000} /* (10, 20, 11) {real, imag} */,
  {32'hc3f5bac0, 32'h00000000} /* (10, 20, 10) {real, imag} */,
  {32'hc402b912, 32'h00000000} /* (10, 20, 9) {real, imag} */,
  {32'hc503c4ac, 32'h00000000} /* (10, 20, 8) {real, imag} */,
  {32'hc5292dcb, 32'h00000000} /* (10, 20, 7) {real, imag} */,
  {32'hc5126d30, 32'h00000000} /* (10, 20, 6) {real, imag} */,
  {32'hc52250d3, 32'h00000000} /* (10, 20, 5) {real, imag} */,
  {32'hc4ef58be, 32'h00000000} /* (10, 20, 4) {real, imag} */,
  {32'hc5463188, 32'h00000000} /* (10, 20, 3) {real, imag} */,
  {32'hc50d16f2, 32'h00000000} /* (10, 20, 2) {real, imag} */,
  {32'hc53561e9, 32'h00000000} /* (10, 20, 1) {real, imag} */,
  {32'hc515e73d, 32'h00000000} /* (10, 20, 0) {real, imag} */,
  {32'hc5a5beb7, 32'h00000000} /* (10, 19, 31) {real, imag} */,
  {32'hc5bed5fd, 32'h00000000} /* (10, 19, 30) {real, imag} */,
  {32'hc5b92b93, 32'h00000000} /* (10, 19, 29) {real, imag} */,
  {32'hc5aae034, 32'h00000000} /* (10, 19, 28) {real, imag} */,
  {32'hc59e26e9, 32'h00000000} /* (10, 19, 27) {real, imag} */,
  {32'hc599a7be, 32'h00000000} /* (10, 19, 26) {real, imag} */,
  {32'hc5960b8e, 32'h00000000} /* (10, 19, 25) {real, imag} */,
  {32'hc592b6ae, 32'h00000000} /* (10, 19, 24) {real, imag} */,
  {32'hc580e3bb, 32'h00000000} /* (10, 19, 23) {real, imag} */,
  {32'hc55ee3f2, 32'h00000000} /* (10, 19, 22) {real, imag} */,
  {32'hc45cf1b4, 32'h00000000} /* (10, 19, 21) {real, imag} */,
  {32'h448f9a26, 32'h00000000} /* (10, 19, 20) {real, imag} */,
  {32'h452ea7ea, 32'h00000000} /* (10, 19, 19) {real, imag} */,
  {32'h4558dd79, 32'h00000000} /* (10, 19, 18) {real, imag} */,
  {32'h459c3472, 32'h00000000} /* (10, 19, 17) {real, imag} */,
  {32'h45ba9c46, 32'h00000000} /* (10, 19, 16) {real, imag} */,
  {32'h45b4457b, 32'h00000000} /* (10, 19, 15) {real, imag} */,
  {32'h45b35025, 32'h00000000} /* (10, 19, 14) {real, imag} */,
  {32'h45876521, 32'h00000000} /* (10, 19, 13) {real, imag} */,
  {32'h456ad093, 32'h00000000} /* (10, 19, 12) {real, imag} */,
  {32'h44c120d1, 32'h00000000} /* (10, 19, 11) {real, imag} */,
  {32'hc3860d38, 32'h00000000} /* (10, 19, 10) {real, imag} */,
  {32'hc50a58b4, 32'h00000000} /* (10, 19, 9) {real, imag} */,
  {32'hc5559602, 32'h00000000} /* (10, 19, 8) {real, imag} */,
  {32'hc5919667, 32'h00000000} /* (10, 19, 7) {real, imag} */,
  {32'hc58fc64f, 32'h00000000} /* (10, 19, 6) {real, imag} */,
  {32'hc5b1698e, 32'h00000000} /* (10, 19, 5) {real, imag} */,
  {32'hc5b5e81c, 32'h00000000} /* (10, 19, 4) {real, imag} */,
  {32'hc5995c54, 32'h00000000} /* (10, 19, 3) {real, imag} */,
  {32'hc5b6c9b2, 32'h00000000} /* (10, 19, 2) {real, imag} */,
  {32'hc5b5ac62, 32'h00000000} /* (10, 19, 1) {real, imag} */,
  {32'hc5a62eac, 32'h00000000} /* (10, 19, 0) {real, imag} */,
  {32'hc5da1e0b, 32'h00000000} /* (10, 18, 31) {real, imag} */,
  {32'hc606ab4e, 32'h00000000} /* (10, 18, 30) {real, imag} */,
  {32'hc5df7dc0, 32'h00000000} /* (10, 18, 29) {real, imag} */,
  {32'hc6090d05, 32'h00000000} /* (10, 18, 28) {real, imag} */,
  {32'hc5f9deed, 32'h00000000} /* (10, 18, 27) {real, imag} */,
  {32'hc5db4aec, 32'h00000000} /* (10, 18, 26) {real, imag} */,
  {32'hc5c8e549, 32'h00000000} /* (10, 18, 25) {real, imag} */,
  {32'hc5d2c786, 32'h00000000} /* (10, 18, 24) {real, imag} */,
  {32'hc593f716, 32'h00000000} /* (10, 18, 23) {real, imag} */,
  {32'hc54a5ede, 32'h00000000} /* (10, 18, 22) {real, imag} */,
  {32'hc4aa3728, 32'h00000000} /* (10, 18, 21) {real, imag} */,
  {32'h44edb390, 32'h00000000} /* (10, 18, 20) {real, imag} */,
  {32'h454cc8c8, 32'h00000000} /* (10, 18, 19) {real, imag} */,
  {32'h459131d1, 32'h00000000} /* (10, 18, 18) {real, imag} */,
  {32'h45b5621e, 32'h00000000} /* (10, 18, 17) {real, imag} */,
  {32'h45d74ffa, 32'h00000000} /* (10, 18, 16) {real, imag} */,
  {32'h45f27d6f, 32'h00000000} /* (10, 18, 15) {real, imag} */,
  {32'h45c92f3c, 32'h00000000} /* (10, 18, 14) {real, imag} */,
  {32'h45b7ab04, 32'h00000000} /* (10, 18, 13) {real, imag} */,
  {32'h459fe543, 32'h00000000} /* (10, 18, 12) {real, imag} */,
  {32'h452612fa, 32'h00000000} /* (10, 18, 11) {real, imag} */,
  {32'hc4bdc470, 32'h00000000} /* (10, 18, 10) {real, imag} */,
  {32'hc54a8ede, 32'h00000000} /* (10, 18, 9) {real, imag} */,
  {32'hc5c0d01a, 32'h00000000} /* (10, 18, 8) {real, imag} */,
  {32'hc5f17986, 32'h00000000} /* (10, 18, 7) {real, imag} */,
  {32'hc5e305b9, 32'h00000000} /* (10, 18, 6) {real, imag} */,
  {32'hc5f68fe0, 32'h00000000} /* (10, 18, 5) {real, imag} */,
  {32'hc5f953b2, 32'h00000000} /* (10, 18, 4) {real, imag} */,
  {32'hc60367aa, 32'h00000000} /* (10, 18, 3) {real, imag} */,
  {32'hc5ed32ff, 32'h00000000} /* (10, 18, 2) {real, imag} */,
  {32'hc5eb19f8, 32'h00000000} /* (10, 18, 1) {real, imag} */,
  {32'hc5e42216, 32'h00000000} /* (10, 18, 0) {real, imag} */,
  {32'hc5fbb9dd, 32'h00000000} /* (10, 17, 31) {real, imag} */,
  {32'hc6057771, 32'h00000000} /* (10, 17, 30) {real, imag} */,
  {32'hc6118476, 32'h00000000} /* (10, 17, 29) {real, imag} */,
  {32'hc6103c5c, 32'h00000000} /* (10, 17, 28) {real, imag} */,
  {32'hc6157e48, 32'h00000000} /* (10, 17, 27) {real, imag} */,
  {32'hc60b6288, 32'h00000000} /* (10, 17, 26) {real, imag} */,
  {32'hc601ee9a, 32'h00000000} /* (10, 17, 25) {real, imag} */,
  {32'hc5f39d30, 32'h00000000} /* (10, 17, 24) {real, imag} */,
  {32'hc5b21238, 32'h00000000} /* (10, 17, 23) {real, imag} */,
  {32'hc58ef7fe, 32'h00000000} /* (10, 17, 22) {real, imag} */,
  {32'hc501fbd9, 32'h00000000} /* (10, 17, 21) {real, imag} */,
  {32'h450ba110, 32'h00000000} /* (10, 17, 20) {real, imag} */,
  {32'h458be1a0, 32'h00000000} /* (10, 17, 19) {real, imag} */,
  {32'h45d84078, 32'h00000000} /* (10, 17, 18) {real, imag} */,
  {32'h45e19f6e, 32'h00000000} /* (10, 17, 17) {real, imag} */,
  {32'h45e673c7, 32'h00000000} /* (10, 17, 16) {real, imag} */,
  {32'h45f629ed, 32'h00000000} /* (10, 17, 15) {real, imag} */,
  {32'h45f9c71e, 32'h00000000} /* (10, 17, 14) {real, imag} */,
  {32'h45c813c9, 32'h00000000} /* (10, 17, 13) {real, imag} */,
  {32'h45a663c8, 32'h00000000} /* (10, 17, 12) {real, imag} */,
  {32'h451ecf3f, 32'h00000000} /* (10, 17, 11) {real, imag} */,
  {32'hc51eb8be, 32'h00000000} /* (10, 17, 10) {real, imag} */,
  {32'hc59937f0, 32'h00000000} /* (10, 17, 9) {real, imag} */,
  {32'hc5cfd406, 32'h00000000} /* (10, 17, 8) {real, imag} */,
  {32'hc5f4a12e, 32'h00000000} /* (10, 17, 7) {real, imag} */,
  {32'hc6152b0f, 32'h00000000} /* (10, 17, 6) {real, imag} */,
  {32'hc60636d0, 32'h00000000} /* (10, 17, 5) {real, imag} */,
  {32'hc609751a, 32'h00000000} /* (10, 17, 4) {real, imag} */,
  {32'hc617e503, 32'h00000000} /* (10, 17, 3) {real, imag} */,
  {32'hc61ddbac, 32'h00000000} /* (10, 17, 2) {real, imag} */,
  {32'hc60c0994, 32'h00000000} /* (10, 17, 1) {real, imag} */,
  {32'hc604ca7e, 32'h00000000} /* (10, 17, 0) {real, imag} */,
  {32'hc607a61e, 32'h00000000} /* (10, 16, 31) {real, imag} */,
  {32'hc6173cdb, 32'h00000000} /* (10, 16, 30) {real, imag} */,
  {32'hc61a6153, 32'h00000000} /* (10, 16, 29) {real, imag} */,
  {32'hc61dce46, 32'h00000000} /* (10, 16, 28) {real, imag} */,
  {32'hc6274184, 32'h00000000} /* (10, 16, 27) {real, imag} */,
  {32'hc60e8e07, 32'h00000000} /* (10, 16, 26) {real, imag} */,
  {32'hc60651c3, 32'h00000000} /* (10, 16, 25) {real, imag} */,
  {32'hc5ef168b, 32'h00000000} /* (10, 16, 24) {real, imag} */,
  {32'hc5c695c9, 32'h00000000} /* (10, 16, 23) {real, imag} */,
  {32'hc57f83b0, 32'h00000000} /* (10, 16, 22) {real, imag} */,
  {32'hc3af50f0, 32'h00000000} /* (10, 16, 21) {real, imag} */,
  {32'h45176371, 32'h00000000} /* (10, 16, 20) {real, imag} */,
  {32'h45ad8486, 32'h00000000} /* (10, 16, 19) {real, imag} */,
  {32'h45dc7c44, 32'h00000000} /* (10, 16, 18) {real, imag} */,
  {32'h45ef64bd, 32'h00000000} /* (10, 16, 17) {real, imag} */,
  {32'h4606c386, 32'h00000000} /* (10, 16, 16) {real, imag} */,
  {32'h45f425a8, 32'h00000000} /* (10, 16, 15) {real, imag} */,
  {32'h45fff882, 32'h00000000} /* (10, 16, 14) {real, imag} */,
  {32'h45e79086, 32'h00000000} /* (10, 16, 13) {real, imag} */,
  {32'h4589cad8, 32'h00000000} /* (10, 16, 12) {real, imag} */,
  {32'h4501210a, 32'h00000000} /* (10, 16, 11) {real, imag} */,
  {32'hc505e231, 32'h00000000} /* (10, 16, 10) {real, imag} */,
  {32'hc59738e0, 32'h00000000} /* (10, 16, 9) {real, imag} */,
  {32'hc5d08aff, 32'h00000000} /* (10, 16, 8) {real, imag} */,
  {32'hc5eede47, 32'h00000000} /* (10, 16, 7) {real, imag} */,
  {32'hc6071954, 32'h00000000} /* (10, 16, 6) {real, imag} */,
  {32'hc603003a, 32'h00000000} /* (10, 16, 5) {real, imag} */,
  {32'hc60f8b3f, 32'h00000000} /* (10, 16, 4) {real, imag} */,
  {32'hc6172fd3, 32'h00000000} /* (10, 16, 3) {real, imag} */,
  {32'hc6296b30, 32'h00000000} /* (10, 16, 2) {real, imag} */,
  {32'hc616c43c, 32'h00000000} /* (10, 16, 1) {real, imag} */,
  {32'hc606d66e, 32'h00000000} /* (10, 16, 0) {real, imag} */,
  {32'hc60fcb34, 32'h00000000} /* (10, 15, 31) {real, imag} */,
  {32'hc61beba4, 32'h00000000} /* (10, 15, 30) {real, imag} */,
  {32'hc6196852, 32'h00000000} /* (10, 15, 29) {real, imag} */,
  {32'hc619fac0, 32'h00000000} /* (10, 15, 28) {real, imag} */,
  {32'hc614225e, 32'h00000000} /* (10, 15, 27) {real, imag} */,
  {32'hc61675b0, 32'h00000000} /* (10, 15, 26) {real, imag} */,
  {32'hc6001835, 32'h00000000} /* (10, 15, 25) {real, imag} */,
  {32'hc5f1559a, 32'h00000000} /* (10, 15, 24) {real, imag} */,
  {32'hc5bad77c, 32'h00000000} /* (10, 15, 23) {real, imag} */,
  {32'hc55274ac, 32'h00000000} /* (10, 15, 22) {real, imag} */,
  {32'h44165f58, 32'h00000000} /* (10, 15, 21) {real, imag} */,
  {32'h45619cf8, 32'h00000000} /* (10, 15, 20) {real, imag} */,
  {32'h4593d2fe, 32'h00000000} /* (10, 15, 19) {real, imag} */,
  {32'h45e35734, 32'h00000000} /* (10, 15, 18) {real, imag} */,
  {32'h45ef611f, 32'h00000000} /* (10, 15, 17) {real, imag} */,
  {32'h45ffec57, 32'h00000000} /* (10, 15, 16) {real, imag} */,
  {32'h45f68663, 32'h00000000} /* (10, 15, 15) {real, imag} */,
  {32'h45e70dd8, 32'h00000000} /* (10, 15, 14) {real, imag} */,
  {32'h45c6b3a4, 32'h00000000} /* (10, 15, 13) {real, imag} */,
  {32'h459f678c, 32'h00000000} /* (10, 15, 12) {real, imag} */,
  {32'h44f4a480, 32'h00000000} /* (10, 15, 11) {real, imag} */,
  {32'hc4e04980, 32'h00000000} /* (10, 15, 10) {real, imag} */,
  {32'hc599be93, 32'h00000000} /* (10, 15, 9) {real, imag} */,
  {32'hc5eed1de, 32'h00000000} /* (10, 15, 8) {real, imag} */,
  {32'hc60169b1, 32'h00000000} /* (10, 15, 7) {real, imag} */,
  {32'hc5fee0d6, 32'h00000000} /* (10, 15, 6) {real, imag} */,
  {32'hc609a1f8, 32'h00000000} /* (10, 15, 5) {real, imag} */,
  {32'hc61d7bf5, 32'h00000000} /* (10, 15, 4) {real, imag} */,
  {32'hc61a8b13, 32'h00000000} /* (10, 15, 3) {real, imag} */,
  {32'hc621bdfe, 32'h00000000} /* (10, 15, 2) {real, imag} */,
  {32'hc6201cdc, 32'h00000000} /* (10, 15, 1) {real, imag} */,
  {32'hc60b5394, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'hc5ff2e80, 32'h00000000} /* (10, 14, 31) {real, imag} */,
  {32'hc60a035e, 32'h00000000} /* (10, 14, 30) {real, imag} */,
  {32'hc60a2955, 32'h00000000} /* (10, 14, 29) {real, imag} */,
  {32'hc6105341, 32'h00000000} /* (10, 14, 28) {real, imag} */,
  {32'hc60029da, 32'h00000000} /* (10, 14, 27) {real, imag} */,
  {32'hc5fef206, 32'h00000000} /* (10, 14, 26) {real, imag} */,
  {32'hc6006523, 32'h00000000} /* (10, 14, 25) {real, imag} */,
  {32'hc5cf96f7, 32'h00000000} /* (10, 14, 24) {real, imag} */,
  {32'hc595d434, 32'h00000000} /* (10, 14, 23) {real, imag} */,
  {32'hc519a910, 32'h00000000} /* (10, 14, 22) {real, imag} */,
  {32'hc4167e48, 32'h00000000} /* (10, 14, 21) {real, imag} */,
  {32'h45213904, 32'h00000000} /* (10, 14, 20) {real, imag} */,
  {32'h459cc538, 32'h00000000} /* (10, 14, 19) {real, imag} */,
  {32'h45c8e5a9, 32'h00000000} /* (10, 14, 18) {real, imag} */,
  {32'h45ed14cb, 32'h00000000} /* (10, 14, 17) {real, imag} */,
  {32'h45ec22a0, 32'h00000000} /* (10, 14, 16) {real, imag} */,
  {32'h45ded652, 32'h00000000} /* (10, 14, 15) {real, imag} */,
  {32'h45de5fdc, 32'h00000000} /* (10, 14, 14) {real, imag} */,
  {32'h45bcc390, 32'h00000000} /* (10, 14, 13) {real, imag} */,
  {32'h45759188, 32'h00000000} /* (10, 14, 12) {real, imag} */,
  {32'h45223139, 32'h00000000} /* (10, 14, 11) {real, imag} */,
  {32'hc48c8dc6, 32'h00000000} /* (10, 14, 10) {real, imag} */,
  {32'hc5995e22, 32'h00000000} /* (10, 14, 9) {real, imag} */,
  {32'hc5c4140d, 32'h00000000} /* (10, 14, 8) {real, imag} */,
  {32'hc5dba57c, 32'h00000000} /* (10, 14, 7) {real, imag} */,
  {32'hc60145d2, 32'h00000000} /* (10, 14, 6) {real, imag} */,
  {32'hc60ad4ce, 32'h00000000} /* (10, 14, 5) {real, imag} */,
  {32'hc60c5f68, 32'h00000000} /* (10, 14, 4) {real, imag} */,
  {32'hc60bc54b, 32'h00000000} /* (10, 14, 3) {real, imag} */,
  {32'hc604b402, 32'h00000000} /* (10, 14, 2) {real, imag} */,
  {32'hc6164944, 32'h00000000} /* (10, 14, 1) {real, imag} */,
  {32'hc6148fcc, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'hc5d25a73, 32'h00000000} /* (10, 13, 31) {real, imag} */,
  {32'hc5d8987e, 32'h00000000} /* (10, 13, 30) {real, imag} */,
  {32'hc5e26268, 32'h00000000} /* (10, 13, 29) {real, imag} */,
  {32'hc5e6b0a6, 32'h00000000} /* (10, 13, 28) {real, imag} */,
  {32'hc5ea4010, 32'h00000000} /* (10, 13, 27) {real, imag} */,
  {32'hc5cebe4b, 32'h00000000} /* (10, 13, 26) {real, imag} */,
  {32'hc5c97d6c, 32'h00000000} /* (10, 13, 25) {real, imag} */,
  {32'hc5b2a204, 32'h00000000} /* (10, 13, 24) {real, imag} */,
  {32'hc58357ac, 32'h00000000} /* (10, 13, 23) {real, imag} */,
  {32'hc52d4a19, 32'h00000000} /* (10, 13, 22) {real, imag} */,
  {32'h43cf8cd8, 32'h00000000} /* (10, 13, 21) {real, imag} */,
  {32'h4517e5f4, 32'h00000000} /* (10, 13, 20) {real, imag} */,
  {32'h4592ea9b, 32'h00000000} /* (10, 13, 19) {real, imag} */,
  {32'h45bfb16b, 32'h00000000} /* (10, 13, 18) {real, imag} */,
  {32'h45bc842a, 32'h00000000} /* (10, 13, 17) {real, imag} */,
  {32'h45c6f238, 32'h00000000} /* (10, 13, 16) {real, imag} */,
  {32'h45c9ac07, 32'h00000000} /* (10, 13, 15) {real, imag} */,
  {32'h45ab7756, 32'h00000000} /* (10, 13, 14) {real, imag} */,
  {32'h459f43fe, 32'h00000000} /* (10, 13, 13) {real, imag} */,
  {32'h4578b63c, 32'h00000000} /* (10, 13, 12) {real, imag} */,
  {32'h45162200, 32'h00000000} /* (10, 13, 11) {real, imag} */,
  {32'hc45b5f28, 32'h00000000} /* (10, 13, 10) {real, imag} */,
  {32'hc5706799, 32'h00000000} /* (10, 13, 9) {real, imag} */,
  {32'hc5b18d92, 32'h00000000} /* (10, 13, 8) {real, imag} */,
  {32'hc5d90bb6, 32'h00000000} /* (10, 13, 7) {real, imag} */,
  {32'hc5e73584, 32'h00000000} /* (10, 13, 6) {real, imag} */,
  {32'hc5ea419e, 32'h00000000} /* (10, 13, 5) {real, imag} */,
  {32'hc5dd3ac8, 32'h00000000} /* (10, 13, 4) {real, imag} */,
  {32'hc5f9d031, 32'h00000000} /* (10, 13, 3) {real, imag} */,
  {32'hc5d744df, 32'h00000000} /* (10, 13, 2) {real, imag} */,
  {32'hc5f8d9c4, 32'h00000000} /* (10, 13, 1) {real, imag} */,
  {32'hc5e9adf2, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'hc597c72a, 32'h00000000} /* (10, 12, 31) {real, imag} */,
  {32'hc5b44e9e, 32'h00000000} /* (10, 12, 30) {real, imag} */,
  {32'hc5a35a8d, 32'h00000000} /* (10, 12, 29) {real, imag} */,
  {32'hc58be364, 32'h00000000} /* (10, 12, 28) {real, imag} */,
  {32'hc587f506, 32'h00000000} /* (10, 12, 27) {real, imag} */,
  {32'hc59b2720, 32'h00000000} /* (10, 12, 26) {real, imag} */,
  {32'hc56e50b7, 32'h00000000} /* (10, 12, 25) {real, imag} */,
  {32'hc58dae6b, 32'h00000000} /* (10, 12, 24) {real, imag} */,
  {32'hc56334f2, 32'h00000000} /* (10, 12, 23) {real, imag} */,
  {32'hc4c627e9, 32'h00000000} /* (10, 12, 22) {real, imag} */,
  {32'hc28ef4a0, 32'h00000000} /* (10, 12, 21) {real, imag} */,
  {32'h4529d717, 32'h00000000} /* (10, 12, 20) {real, imag} */,
  {32'h4592983c, 32'h00000000} /* (10, 12, 19) {real, imag} */,
  {32'h4585ff9a, 32'h00000000} /* (10, 12, 18) {real, imag} */,
  {32'h45ac7a4a, 32'h00000000} /* (10, 12, 17) {real, imag} */,
  {32'h45b9190e, 32'h00000000} /* (10, 12, 16) {real, imag} */,
  {32'h45962582, 32'h00000000} /* (10, 12, 15) {real, imag} */,
  {32'h45867814, 32'h00000000} /* (10, 12, 14) {real, imag} */,
  {32'h456d72e2, 32'h00000000} /* (10, 12, 13) {real, imag} */,
  {32'h452df2ef, 32'h00000000} /* (10, 12, 12) {real, imag} */,
  {32'h44698d4c, 32'h00000000} /* (10, 12, 11) {real, imag} */,
  {32'hc4c252d0, 32'h00000000} /* (10, 12, 10) {real, imag} */,
  {32'hc550b715, 32'h00000000} /* (10, 12, 9) {real, imag} */,
  {32'hc5890221, 32'h00000000} /* (10, 12, 8) {real, imag} */,
  {32'hc5afbfbf, 32'h00000000} /* (10, 12, 7) {real, imag} */,
  {32'hc5a9e9a7, 32'h00000000} /* (10, 12, 6) {real, imag} */,
  {32'hc5b3afa0, 32'h00000000} /* (10, 12, 5) {real, imag} */,
  {32'hc5b10a00, 32'h00000000} /* (10, 12, 4) {real, imag} */,
  {32'hc59ce864, 32'h00000000} /* (10, 12, 3) {real, imag} */,
  {32'hc594259a, 32'h00000000} /* (10, 12, 2) {real, imag} */,
  {32'hc5a4d4d4, 32'h00000000} /* (10, 12, 1) {real, imag} */,
  {32'hc59e8a2a, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hc4f42490, 32'h00000000} /* (10, 11, 31) {real, imag} */,
  {32'hc497c213, 32'h00000000} /* (10, 11, 30) {real, imag} */,
  {32'hc4a9bcb4, 32'h00000000} /* (10, 11, 29) {real, imag} */,
  {32'hc4fcd667, 32'h00000000} /* (10, 11, 28) {real, imag} */,
  {32'hc4d32a8c, 32'h00000000} /* (10, 11, 27) {real, imag} */,
  {32'hc4dadd4a, 32'h00000000} /* (10, 11, 26) {real, imag} */,
  {32'hc497e385, 32'h00000000} /* (10, 11, 25) {real, imag} */,
  {32'hc434f2a6, 32'h00000000} /* (10, 11, 24) {real, imag} */,
  {32'hc3c61c54, 32'h00000000} /* (10, 11, 23) {real, imag} */,
  {32'h439b7c04, 32'h00000000} /* (10, 11, 22) {real, imag} */,
  {32'h446553b0, 32'h00000000} /* (10, 11, 21) {real, imag} */,
  {32'h450b661a, 32'h00000000} /* (10, 11, 20) {real, imag} */,
  {32'h456975de, 32'h00000000} /* (10, 11, 19) {real, imag} */,
  {32'h45817bfd, 32'h00000000} /* (10, 11, 18) {real, imag} */,
  {32'h4549a0b3, 32'h00000000} /* (10, 11, 17) {real, imag} */,
  {32'h45806287, 32'h00000000} /* (10, 11, 16) {real, imag} */,
  {32'h457a6f2a, 32'h00000000} /* (10, 11, 15) {real, imag} */,
  {32'h453ba140, 32'h00000000} /* (10, 11, 14) {real, imag} */,
  {32'h45081faa, 32'h00000000} /* (10, 11, 13) {real, imag} */,
  {32'h44b7695b, 32'h00000000} /* (10, 11, 12) {real, imag} */,
  {32'h44875cc4, 32'h00000000} /* (10, 11, 11) {real, imag} */,
  {32'hc486cd40, 32'h00000000} /* (10, 11, 10) {real, imag} */,
  {32'hc4b5eeb7, 32'h00000000} /* (10, 11, 9) {real, imag} */,
  {32'hc4e747bf, 32'h00000000} /* (10, 11, 8) {real, imag} */,
  {32'hc50c0c18, 32'h00000000} /* (10, 11, 7) {real, imag} */,
  {32'hc52e3e1c, 32'h00000000} /* (10, 11, 6) {real, imag} */,
  {32'hc50189bf, 32'h00000000} /* (10, 11, 5) {real, imag} */,
  {32'hc51a9048, 32'h00000000} /* (10, 11, 4) {real, imag} */,
  {32'hc51cb90e, 32'h00000000} /* (10, 11, 3) {real, imag} */,
  {32'hc53a6952, 32'h00000000} /* (10, 11, 2) {real, imag} */,
  {32'hc506003f, 32'h00000000} /* (10, 11, 1) {real, imag} */,
  {32'hc4d43e25, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h44d5d1c2, 32'h00000000} /* (10, 10, 31) {real, imag} */,
  {32'h4528d565, 32'h00000000} /* (10, 10, 30) {real, imag} */,
  {32'h456ef72a, 32'h00000000} /* (10, 10, 29) {real, imag} */,
  {32'h451483c2, 32'h00000000} /* (10, 10, 28) {real, imag} */,
  {32'h450639da, 32'h00000000} /* (10, 10, 27) {real, imag} */,
  {32'h4555b119, 32'h00000000} /* (10, 10, 26) {real, imag} */,
  {32'h45304cf9, 32'h00000000} /* (10, 10, 25) {real, imag} */,
  {32'h453e2628, 32'h00000000} /* (10, 10, 24) {real, imag} */,
  {32'h4560e307, 32'h00000000} /* (10, 10, 23) {real, imag} */,
  {32'h452d99ae, 32'h00000000} /* (10, 10, 22) {real, imag} */,
  {32'h454cddc0, 32'h00000000} /* (10, 10, 21) {real, imag} */,
  {32'h4515cc19, 32'h00000000} /* (10, 10, 20) {real, imag} */,
  {32'h44036e99, 32'h00000000} /* (10, 10, 19) {real, imag} */,
  {32'h4465babe, 32'h00000000} /* (10, 10, 18) {real, imag} */,
  {32'h44663b74, 32'h00000000} /* (10, 10, 17) {real, imag} */,
  {32'hc33a9214, 32'h00000000} /* (10, 10, 16) {real, imag} */,
  {32'hc355ef44, 32'h00000000} /* (10, 10, 15) {real, imag} */,
  {32'hc3de9fd0, 32'h00000000} /* (10, 10, 14) {real, imag} */,
  {32'hc43999aa, 32'h00000000} /* (10, 10, 13) {real, imag} */,
  {32'hc4b94c1d, 32'h00000000} /* (10, 10, 12) {real, imag} */,
  {32'hc48df5b5, 32'h00000000} /* (10, 10, 11) {real, imag} */,
  {32'hc423ac20, 32'h00000000} /* (10, 10, 10) {real, imag} */,
  {32'hc2092440, 32'h00000000} /* (10, 10, 9) {real, imag} */,
  {32'h43d75754, 32'h00000000} /* (10, 10, 8) {real, imag} */,
  {32'h45014195, 32'h00000000} /* (10, 10, 7) {real, imag} */,
  {32'h450a799e, 32'h00000000} /* (10, 10, 6) {real, imag} */,
  {32'h4512a020, 32'h00000000} /* (10, 10, 5) {real, imag} */,
  {32'h451d0bdf, 32'h00000000} /* (10, 10, 4) {real, imag} */,
  {32'h4469f5af, 32'h00000000} /* (10, 10, 3) {real, imag} */,
  {32'h446bf85e, 32'h00000000} /* (10, 10, 2) {real, imag} */,
  {32'h44be8bc6, 32'h00000000} /* (10, 10, 1) {real, imag} */,
  {32'h44d57f64, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h45a53551, 32'h00000000} /* (10, 9, 31) {real, imag} */,
  {32'h45a3874e, 32'h00000000} /* (10, 9, 30) {real, imag} */,
  {32'h45c55e7c, 32'h00000000} /* (10, 9, 29) {real, imag} */,
  {32'h45faa747, 32'h00000000} /* (10, 9, 28) {real, imag} */,
  {32'h45d5e574, 32'h00000000} /* (10, 9, 27) {real, imag} */,
  {32'h45c7259e, 32'h00000000} /* (10, 9, 26) {real, imag} */,
  {32'h45c5aa34, 32'h00000000} /* (10, 9, 25) {real, imag} */,
  {32'h45ca879c, 32'h00000000} /* (10, 9, 24) {real, imag} */,
  {32'h45b1a8d0, 32'h00000000} /* (10, 9, 23) {real, imag} */,
  {32'h45b22211, 32'h00000000} /* (10, 9, 22) {real, imag} */,
  {32'h456a017c, 32'h00000000} /* (10, 9, 21) {real, imag} */,
  {32'h4516c11c, 32'h00000000} /* (10, 9, 20) {real, imag} */,
  {32'hc4095360, 32'h00000000} /* (10, 9, 19) {real, imag} */,
  {32'hc4b7ff2e, 32'h00000000} /* (10, 9, 18) {real, imag} */,
  {32'hc4bb8d04, 32'h00000000} /* (10, 9, 17) {real, imag} */,
  {32'hc55d1af9, 32'h00000000} /* (10, 9, 16) {real, imag} */,
  {32'hc55b219a, 32'h00000000} /* (10, 9, 15) {real, imag} */,
  {32'hc52e5f6d, 32'h00000000} /* (10, 9, 14) {real, imag} */,
  {32'hc519565b, 32'h00000000} /* (10, 9, 13) {real, imag} */,
  {32'hc536679a, 32'h00000000} /* (10, 9, 12) {real, imag} */,
  {32'hc5289aff, 32'h00000000} /* (10, 9, 11) {real, imag} */,
  {32'hc3f10248, 32'h00000000} /* (10, 9, 10) {real, imag} */,
  {32'h44d83208, 32'h00000000} /* (10, 9, 9) {real, imag} */,
  {32'h453520d4, 32'h00000000} /* (10, 9, 8) {real, imag} */,
  {32'h45737944, 32'h00000000} /* (10, 9, 7) {real, imag} */,
  {32'h457f050a, 32'h00000000} /* (10, 9, 6) {real, imag} */,
  {32'h4587bc95, 32'h00000000} /* (10, 9, 5) {real, imag} */,
  {32'h45901784, 32'h00000000} /* (10, 9, 4) {real, imag} */,
  {32'h45b2e1ed, 32'h00000000} /* (10, 9, 3) {real, imag} */,
  {32'h4581f38c, 32'h00000000} /* (10, 9, 2) {real, imag} */,
  {32'h458cefad, 32'h00000000} /* (10, 9, 1) {real, imag} */,
  {32'h458a1eb2, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'h45c9bf51, 32'h00000000} /* (10, 8, 31) {real, imag} */,
  {32'h45e5c75b, 32'h00000000} /* (10, 8, 30) {real, imag} */,
  {32'h460a8cb6, 32'h00000000} /* (10, 8, 29) {real, imag} */,
  {32'h4606d14e, 32'h00000000} /* (10, 8, 28) {real, imag} */,
  {32'h46210348, 32'h00000000} /* (10, 8, 27) {real, imag} */,
  {32'h46132818, 32'h00000000} /* (10, 8, 26) {real, imag} */,
  {32'h46079600, 32'h00000000} /* (10, 8, 25) {real, imag} */,
  {32'h45fe3e40, 32'h00000000} /* (10, 8, 24) {real, imag} */,
  {32'h45fd1a51, 32'h00000000} /* (10, 8, 23) {real, imag} */,
  {32'h45d41713, 32'h00000000} /* (10, 8, 22) {real, imag} */,
  {32'h45952260, 32'h00000000} /* (10, 8, 21) {real, imag} */,
  {32'h4521082c, 32'h00000000} /* (10, 8, 20) {real, imag} */,
  {32'h43501dc0, 32'h00000000} /* (10, 8, 19) {real, imag} */,
  {32'hc4dff264, 32'h00000000} /* (10, 8, 18) {real, imag} */,
  {32'hc538a149, 32'h00000000} /* (10, 8, 17) {real, imag} */,
  {32'hc56a91f8, 32'h00000000} /* (10, 8, 16) {real, imag} */,
  {32'hc5845f13, 32'h00000000} /* (10, 8, 15) {real, imag} */,
  {32'hc595cb23, 32'h00000000} /* (10, 8, 14) {real, imag} */,
  {32'hc59242e4, 32'h00000000} /* (10, 8, 13) {real, imag} */,
  {32'hc5808d25, 32'h00000000} /* (10, 8, 12) {real, imag} */,
  {32'hc5812661, 32'h00000000} /* (10, 8, 11) {real, imag} */,
  {32'hc48ba12c, 32'h00000000} /* (10, 8, 10) {real, imag} */,
  {32'h4529374a, 32'h00000000} /* (10, 8, 9) {real, imag} */,
  {32'h45533d0c, 32'h00000000} /* (10, 8, 8) {real, imag} */,
  {32'h45ac42b5, 32'h00000000} /* (10, 8, 7) {real, imag} */,
  {32'h45b6e907, 32'h00000000} /* (10, 8, 6) {real, imag} */,
  {32'h45b883ac, 32'h00000000} /* (10, 8, 5) {real, imag} */,
  {32'h45db10fe, 32'h00000000} /* (10, 8, 4) {real, imag} */,
  {32'h45db4d78, 32'h00000000} /* (10, 8, 3) {real, imag} */,
  {32'h45f041ab, 32'h00000000} /* (10, 8, 2) {real, imag} */,
  {32'h45e6b1fe, 32'h00000000} /* (10, 8, 1) {real, imag} */,
  {32'h45e16f3a, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h460d889e, 32'h00000000} /* (10, 7, 31) {real, imag} */,
  {32'h4612be18, 32'h00000000} /* (10, 7, 30) {real, imag} */,
  {32'h4634b021, 32'h00000000} /* (10, 7, 29) {real, imag} */,
  {32'h4627617e, 32'h00000000} /* (10, 7, 28) {real, imag} */,
  {32'h462f5bcf, 32'h00000000} /* (10, 7, 27) {real, imag} */,
  {32'h462d641e, 32'h00000000} /* (10, 7, 26) {real, imag} */,
  {32'h461e8886, 32'h00000000} /* (10, 7, 25) {real, imag} */,
  {32'h461edf12, 32'h00000000} /* (10, 7, 24) {real, imag} */,
  {32'h4615a881, 32'h00000000} /* (10, 7, 23) {real, imag} */,
  {32'h460a11d4, 32'h00000000} /* (10, 7, 22) {real, imag} */,
  {32'h45bfc064, 32'h00000000} /* (10, 7, 21) {real, imag} */,
  {32'h455ae567, 32'h00000000} /* (10, 7, 20) {real, imag} */,
  {32'h44c4184a, 32'h00000000} /* (10, 7, 19) {real, imag} */,
  {32'hc4bf6ae4, 32'h00000000} /* (10, 7, 18) {real, imag} */,
  {32'hc52af071, 32'h00000000} /* (10, 7, 17) {real, imag} */,
  {32'hc58a8304, 32'h00000000} /* (10, 7, 16) {real, imag} */,
  {32'hc5a6c846, 32'h00000000} /* (10, 7, 15) {real, imag} */,
  {32'hc5b479a7, 32'h00000000} /* (10, 7, 14) {real, imag} */,
  {32'hc5a9bf2a, 32'h00000000} /* (10, 7, 13) {real, imag} */,
  {32'hc5b15a8c, 32'h00000000} /* (10, 7, 12) {real, imag} */,
  {32'hc58e2a3a, 32'h00000000} /* (10, 7, 11) {real, imag} */,
  {32'hc4b2139c, 32'h00000000} /* (10, 7, 10) {real, imag} */,
  {32'h44199058, 32'h00000000} /* (10, 7, 9) {real, imag} */,
  {32'h45672789, 32'h00000000} /* (10, 7, 8) {real, imag} */,
  {32'h45c01f9d, 32'h00000000} /* (10, 7, 7) {real, imag} */,
  {32'h45d11d4f, 32'h00000000} /* (10, 7, 6) {real, imag} */,
  {32'h45d572b8, 32'h00000000} /* (10, 7, 5) {real, imag} */,
  {32'h46046f54, 32'h00000000} /* (10, 7, 4) {real, imag} */,
  {32'h461544cf, 32'h00000000} /* (10, 7, 3) {real, imag} */,
  {32'h46069ba6, 32'h00000000} /* (10, 7, 2) {real, imag} */,
  {32'h4617cc5a, 32'h00000000} /* (10, 7, 1) {real, imag} */,
  {32'h4605f05b, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h46297092, 32'h00000000} /* (10, 6, 31) {real, imag} */,
  {32'h46263adc, 32'h00000000} /* (10, 6, 30) {real, imag} */,
  {32'h4630af67, 32'h00000000} /* (10, 6, 29) {real, imag} */,
  {32'h4642fa22, 32'h00000000} /* (10, 6, 28) {real, imag} */,
  {32'h464223e3, 32'h00000000} /* (10, 6, 27) {real, imag} */,
  {32'h46422f26, 32'h00000000} /* (10, 6, 26) {real, imag} */,
  {32'h4637b650, 32'h00000000} /* (10, 6, 25) {real, imag} */,
  {32'h46390750, 32'h00000000} /* (10, 6, 24) {real, imag} */,
  {32'h46276a19, 32'h00000000} /* (10, 6, 23) {real, imag} */,
  {32'h461738b1, 32'h00000000} /* (10, 6, 22) {real, imag} */,
  {32'h46024691, 32'h00000000} /* (10, 6, 21) {real, imag} */,
  {32'h459dc003, 32'h00000000} /* (10, 6, 20) {real, imag} */,
  {32'h452c57eb, 32'h00000000} /* (10, 6, 19) {real, imag} */,
  {32'h430e1de0, 32'h00000000} /* (10, 6, 18) {real, imag} */,
  {32'hc4d392fc, 32'h00000000} /* (10, 6, 17) {real, imag} */,
  {32'hc57c6ffd, 32'h00000000} /* (10, 6, 16) {real, imag} */,
  {32'hc599d156, 32'h00000000} /* (10, 6, 15) {real, imag} */,
  {32'hc5c52cb0, 32'h00000000} /* (10, 6, 14) {real, imag} */,
  {32'hc5c1da42, 32'h00000000} /* (10, 6, 13) {real, imag} */,
  {32'hc5bfcc2d, 32'h00000000} /* (10, 6, 12) {real, imag} */,
  {32'hc596daee, 32'h00000000} /* (10, 6, 11) {real, imag} */,
  {32'hc4dc94d4, 32'h00000000} /* (10, 6, 10) {real, imag} */,
  {32'hc3a30a70, 32'h00000000} /* (10, 6, 9) {real, imag} */,
  {32'h44c3535c, 32'h00000000} /* (10, 6, 8) {real, imag} */,
  {32'h45809ea6, 32'h00000000} /* (10, 6, 7) {real, imag} */,
  {32'h45b5eaee, 32'h00000000} /* (10, 6, 6) {real, imag} */,
  {32'h45e78196, 32'h00000000} /* (10, 6, 5) {real, imag} */,
  {32'h460d72fe, 32'h00000000} /* (10, 6, 4) {real, imag} */,
  {32'h4624c717, 32'h00000000} /* (10, 6, 3) {real, imag} */,
  {32'h461ef9ae, 32'h00000000} /* (10, 6, 2) {real, imag} */,
  {32'h462ac870, 32'h00000000} /* (10, 6, 1) {real, imag} */,
  {32'h462700ee, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'h462930be, 32'h00000000} /* (10, 5, 31) {real, imag} */,
  {32'h46375582, 32'h00000000} /* (10, 5, 30) {real, imag} */,
  {32'h46412d00, 32'h00000000} /* (10, 5, 29) {real, imag} */,
  {32'h46498a40, 32'h00000000} /* (10, 5, 28) {real, imag} */,
  {32'h465ee984, 32'h00000000} /* (10, 5, 27) {real, imag} */,
  {32'h4657edc2, 32'h00000000} /* (10, 5, 26) {real, imag} */,
  {32'h4654b7d4, 32'h00000000} /* (10, 5, 25) {real, imag} */,
  {32'h46381d46, 32'h00000000} /* (10, 5, 24) {real, imag} */,
  {32'h463c023e, 32'h00000000} /* (10, 5, 23) {real, imag} */,
  {32'h4629bcc6, 32'h00000000} /* (10, 5, 22) {real, imag} */,
  {32'h461a6c03, 32'h00000000} /* (10, 5, 21) {real, imag} */,
  {32'h45edec52, 32'h00000000} /* (10, 5, 20) {real, imag} */,
  {32'h459d0091, 32'h00000000} /* (10, 5, 19) {real, imag} */,
  {32'h4514d214, 32'h00000000} /* (10, 5, 18) {real, imag} */,
  {32'h445472f0, 32'h00000000} /* (10, 5, 17) {real, imag} */,
  {32'hc4c033d0, 32'h00000000} /* (10, 5, 16) {real, imag} */,
  {32'hc58c12bc, 32'h00000000} /* (10, 5, 15) {real, imag} */,
  {32'hc5b23f0f, 32'h00000000} /* (10, 5, 14) {real, imag} */,
  {32'hc5c4422d, 32'h00000000} /* (10, 5, 13) {real, imag} */,
  {32'hc5e3d6b3, 32'h00000000} /* (10, 5, 12) {real, imag} */,
  {32'hc5ce2ce8, 32'h00000000} /* (10, 5, 11) {real, imag} */,
  {32'hc54500b0, 32'h00000000} /* (10, 5, 10) {real, imag} */,
  {32'hc4bafefc, 32'h00000000} /* (10, 5, 9) {real, imag} */,
  {32'h43284800, 32'h00000000} /* (10, 5, 8) {real, imag} */,
  {32'h44f59bb0, 32'h00000000} /* (10, 5, 7) {real, imag} */,
  {32'h456caa56, 32'h00000000} /* (10, 5, 6) {real, imag} */,
  {32'h45cf4aba, 32'h00000000} /* (10, 5, 5) {real, imag} */,
  {32'h460197ac, 32'h00000000} /* (10, 5, 4) {real, imag} */,
  {32'h46157c18, 32'h00000000} /* (10, 5, 3) {real, imag} */,
  {32'h46356877, 32'h00000000} /* (10, 5, 2) {real, imag} */,
  {32'h4639b6b6, 32'h00000000} /* (10, 5, 1) {real, imag} */,
  {32'h4628fc88, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h46394a78, 32'h00000000} /* (10, 4, 31) {real, imag} */,
  {32'h46475b54, 32'h00000000} /* (10, 4, 30) {real, imag} */,
  {32'h4650547b, 32'h00000000} /* (10, 4, 29) {real, imag} */,
  {32'h465c759a, 32'h00000000} /* (10, 4, 28) {real, imag} */,
  {32'h4664786f, 32'h00000000} /* (10, 4, 27) {real, imag} */,
  {32'h4661c8f4, 32'h00000000} /* (10, 4, 26) {real, imag} */,
  {32'h465720a9, 32'h00000000} /* (10, 4, 25) {real, imag} */,
  {32'h46457839, 32'h00000000} /* (10, 4, 24) {real, imag} */,
  {32'h463d456c, 32'h00000000} /* (10, 4, 23) {real, imag} */,
  {32'h463a6aff, 32'h00000000} /* (10, 4, 22) {real, imag} */,
  {32'h4625a597, 32'h00000000} /* (10, 4, 21) {real, imag} */,
  {32'h46065b1e, 32'h00000000} /* (10, 4, 20) {real, imag} */,
  {32'h45be280d, 32'h00000000} /* (10, 4, 19) {real, imag} */,
  {32'h45861d09, 32'h00000000} /* (10, 4, 18) {real, imag} */,
  {32'h45414166, 32'h00000000} /* (10, 4, 17) {real, imag} */,
  {32'hc40fcbe0, 32'h00000000} /* (10, 4, 16) {real, imag} */,
  {32'hc58f2fc3, 32'h00000000} /* (10, 4, 15) {real, imag} */,
  {32'hc58f0c2d, 32'h00000000} /* (10, 4, 14) {real, imag} */,
  {32'hc5c004ba, 32'h00000000} /* (10, 4, 13) {real, imag} */,
  {32'hc5dc0d28, 32'h00000000} /* (10, 4, 12) {real, imag} */,
  {32'hc5cf9116, 32'h00000000} /* (10, 4, 11) {real, imag} */,
  {32'hc591de53, 32'h00000000} /* (10, 4, 10) {real, imag} */,
  {32'hc5374124, 32'h00000000} /* (10, 4, 9) {real, imag} */,
  {32'hc4f464c8, 32'h00000000} /* (10, 4, 8) {real, imag} */,
  {32'h430dc620, 32'h00000000} /* (10, 4, 7) {real, imag} */,
  {32'h45252ee8, 32'h00000000} /* (10, 4, 6) {real, imag} */,
  {32'h45b21fb2, 32'h00000000} /* (10, 4, 5) {real, imag} */,
  {32'h45f7b37f, 32'h00000000} /* (10, 4, 4) {real, imag} */,
  {32'h461b0306, 32'h00000000} /* (10, 4, 3) {real, imag} */,
  {32'h4632f59a, 32'h00000000} /* (10, 4, 2) {real, imag} */,
  {32'h4643cf24, 32'h00000000} /* (10, 4, 1) {real, imag} */,
  {32'h4639e642, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'h463e3029, 32'h00000000} /* (10, 3, 31) {real, imag} */,
  {32'h46503fc5, 32'h00000000} /* (10, 3, 30) {real, imag} */,
  {32'h46559aca, 32'h00000000} /* (10, 3, 29) {real, imag} */,
  {32'h466eae4c, 32'h00000000} /* (10, 3, 28) {real, imag} */,
  {32'h4657e89e, 32'h00000000} /* (10, 3, 27) {real, imag} */,
  {32'h46591661, 32'h00000000} /* (10, 3, 26) {real, imag} */,
  {32'h4654c72e, 32'h00000000} /* (10, 3, 25) {real, imag} */,
  {32'h4668b703, 32'h00000000} /* (10, 3, 24) {real, imag} */,
  {32'h4645d6ce, 32'h00000000} /* (10, 3, 23) {real, imag} */,
  {32'h4632105c, 32'h00000000} /* (10, 3, 22) {real, imag} */,
  {32'h4630bd2a, 32'h00000000} /* (10, 3, 21) {real, imag} */,
  {32'h4610dc4b, 32'h00000000} /* (10, 3, 20) {real, imag} */,
  {32'h45e1e1d8, 32'h00000000} /* (10, 3, 19) {real, imag} */,
  {32'h459a871b, 32'h00000000} /* (10, 3, 18) {real, imag} */,
  {32'h454ac1a2, 32'h00000000} /* (10, 3, 17) {real, imag} */,
  {32'hc3a80270, 32'h00000000} /* (10, 3, 16) {real, imag} */,
  {32'hc56d5248, 32'h00000000} /* (10, 3, 15) {real, imag} */,
  {32'hc5ab934e, 32'h00000000} /* (10, 3, 14) {real, imag} */,
  {32'hc5c9c6e0, 32'h00000000} /* (10, 3, 13) {real, imag} */,
  {32'hc5c3fdec, 32'h00000000} /* (10, 3, 12) {real, imag} */,
  {32'hc5ded268, 32'h00000000} /* (10, 3, 11) {real, imag} */,
  {32'hc5ad8f3e, 32'h00000000} /* (10, 3, 10) {real, imag} */,
  {32'hc5827505, 32'h00000000} /* (10, 3, 9) {real, imag} */,
  {32'hc569c664, 32'h00000000} /* (10, 3, 8) {real, imag} */,
  {32'hc4cb7a38, 32'h00000000} /* (10, 3, 7) {real, imag} */,
  {32'h44c6765c, 32'h00000000} /* (10, 3, 6) {real, imag} */,
  {32'h4590b0b3, 32'h00000000} /* (10, 3, 5) {real, imag} */,
  {32'h46070ded, 32'h00000000} /* (10, 3, 4) {real, imag} */,
  {32'h461f2ec8, 32'h00000000} /* (10, 3, 3) {real, imag} */,
  {32'h463efb5e, 32'h00000000} /* (10, 3, 2) {real, imag} */,
  {32'h4642483a, 32'h00000000} /* (10, 3, 1) {real, imag} */,
  {32'h46428400, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'h463cffda, 32'h00000000} /* (10, 2, 31) {real, imag} */,
  {32'h464cd155, 32'h00000000} /* (10, 2, 30) {real, imag} */,
  {32'h465e2171, 32'h00000000} /* (10, 2, 29) {real, imag} */,
  {32'h4663a652, 32'h00000000} /* (10, 2, 28) {real, imag} */,
  {32'h46623f5c, 32'h00000000} /* (10, 2, 27) {real, imag} */,
  {32'h46578ebc, 32'h00000000} /* (10, 2, 26) {real, imag} */,
  {32'h465e6ab5, 32'h00000000} /* (10, 2, 25) {real, imag} */,
  {32'h464e6f84, 32'h00000000} /* (10, 2, 24) {real, imag} */,
  {32'h464907f1, 32'h00000000} /* (10, 2, 23) {real, imag} */,
  {32'h462f13ff, 32'h00000000} /* (10, 2, 22) {real, imag} */,
  {32'h461baea0, 32'h00000000} /* (10, 2, 21) {real, imag} */,
  {32'h4609ea6e, 32'h00000000} /* (10, 2, 20) {real, imag} */,
  {32'h45fa0aa8, 32'h00000000} /* (10, 2, 19) {real, imag} */,
  {32'h45aba438, 32'h00000000} /* (10, 2, 18) {real, imag} */,
  {32'h454c3b6c, 32'h00000000} /* (10, 2, 17) {real, imag} */,
  {32'hc22ad580, 32'h00000000} /* (10, 2, 16) {real, imag} */,
  {32'hc56e844c, 32'h00000000} /* (10, 2, 15) {real, imag} */,
  {32'hc5d30afa, 32'h00000000} /* (10, 2, 14) {real, imag} */,
  {32'hc5bfbcfe, 32'h00000000} /* (10, 2, 13) {real, imag} */,
  {32'hc5dce9dc, 32'h00000000} /* (10, 2, 12) {real, imag} */,
  {32'hc5debaf1, 32'h00000000} /* (10, 2, 11) {real, imag} */,
  {32'hc5bbea67, 32'h00000000} /* (10, 2, 10) {real, imag} */,
  {32'hc58ce916, 32'h00000000} /* (10, 2, 9) {real, imag} */,
  {32'hc571c008, 32'h00000000} /* (10, 2, 8) {real, imag} */,
  {32'hc4eb7df0, 32'h00000000} /* (10, 2, 7) {real, imag} */,
  {32'h44c83678, 32'h00000000} /* (10, 2, 6) {real, imag} */,
  {32'h45925934, 32'h00000000} /* (10, 2, 5) {real, imag} */,
  {32'h45ee827c, 32'h00000000} /* (10, 2, 4) {real, imag} */,
  {32'h4620aea4, 32'h00000000} /* (10, 2, 3) {real, imag} */,
  {32'h4631e4e4, 32'h00000000} /* (10, 2, 2) {real, imag} */,
  {32'h463a80fb, 32'h00000000} /* (10, 2, 1) {real, imag} */,
  {32'h463f8d44, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'h463fb5f4, 32'h00000000} /* (10, 1, 31) {real, imag} */,
  {32'h464cfc28, 32'h00000000} /* (10, 1, 30) {real, imag} */,
  {32'h46635db0, 32'h00000000} /* (10, 1, 29) {real, imag} */,
  {32'h466c4fb5, 32'h00000000} /* (10, 1, 28) {real, imag} */,
  {32'h4667a144, 32'h00000000} /* (10, 1, 27) {real, imag} */,
  {32'h465f741f, 32'h00000000} /* (10, 1, 26) {real, imag} */,
  {32'h465510f0, 32'h00000000} /* (10, 1, 25) {real, imag} */,
  {32'h465076ba, 32'h00000000} /* (10, 1, 24) {real, imag} */,
  {32'h4639b24e, 32'h00000000} /* (10, 1, 23) {real, imag} */,
  {32'h46215f78, 32'h00000000} /* (10, 1, 22) {real, imag} */,
  {32'h460e5928, 32'h00000000} /* (10, 1, 21) {real, imag} */,
  {32'h45f2bc2e, 32'h00000000} /* (10, 1, 20) {real, imag} */,
  {32'h45cefdbd, 32'h00000000} /* (10, 1, 19) {real, imag} */,
  {32'h459e3b25, 32'h00000000} /* (10, 1, 18) {real, imag} */,
  {32'h45191cdc, 32'h00000000} /* (10, 1, 17) {real, imag} */,
  {32'hc4331978, 32'h00000000} /* (10, 1, 16) {real, imag} */,
  {32'hc580c75f, 32'h00000000} /* (10, 1, 15) {real, imag} */,
  {32'hc5b85434, 32'h00000000} /* (10, 1, 14) {real, imag} */,
  {32'hc5f6c1f5, 32'h00000000} /* (10, 1, 13) {real, imag} */,
  {32'hc5df65ee, 32'h00000000} /* (10, 1, 12) {real, imag} */,
  {32'hc5bb66b4, 32'h00000000} /* (10, 1, 11) {real, imag} */,
  {32'hc5b22022, 32'h00000000} /* (10, 1, 10) {real, imag} */,
  {32'hc54858f2, 32'h00000000} /* (10, 1, 9) {real, imag} */,
  {32'hc4d58604, 32'h00000000} /* (10, 1, 8) {real, imag} */,
  {32'hc3c628b0, 32'h00000000} /* (10, 1, 7) {real, imag} */,
  {32'h44f2cb0c, 32'h00000000} /* (10, 1, 6) {real, imag} */,
  {32'h45a11f91, 32'h00000000} /* (10, 1, 5) {real, imag} */,
  {32'h45fba82a, 32'h00000000} /* (10, 1, 4) {real, imag} */,
  {32'h461d0a56, 32'h00000000} /* (10, 1, 3) {real, imag} */,
  {32'h462ce1a0, 32'h00000000} /* (10, 1, 2) {real, imag} */,
  {32'h4639faa4, 32'h00000000} /* (10, 1, 1) {real, imag} */,
  {32'h4636e57c, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h464108d5, 32'h00000000} /* (10, 0, 31) {real, imag} */,
  {32'h464bf7e1, 32'h00000000} /* (10, 0, 30) {real, imag} */,
  {32'h4657a7b0, 32'h00000000} /* (10, 0, 29) {real, imag} */,
  {32'h46610ea7, 32'h00000000} /* (10, 0, 28) {real, imag} */,
  {32'h4665685b, 32'h00000000} /* (10, 0, 27) {real, imag} */,
  {32'h4655942c, 32'h00000000} /* (10, 0, 26) {real, imag} */,
  {32'h4647d43a, 32'h00000000} /* (10, 0, 25) {real, imag} */,
  {32'h4640e946, 32'h00000000} /* (10, 0, 24) {real, imag} */,
  {32'h462ac504, 32'h00000000} /* (10, 0, 23) {real, imag} */,
  {32'h46134545, 32'h00000000} /* (10, 0, 22) {real, imag} */,
  {32'h45f18fd4, 32'h00000000} /* (10, 0, 21) {real, imag} */,
  {32'h45b6a5d6, 32'h00000000} /* (10, 0, 20) {real, imag} */,
  {32'h457d4dff, 32'h00000000} /* (10, 0, 19) {real, imag} */,
  {32'h4536cdb1, 32'h00000000} /* (10, 0, 18) {real, imag} */,
  {32'h441f7ec8, 32'h00000000} /* (10, 0, 17) {real, imag} */,
  {32'hc4eeeb60, 32'h00000000} /* (10, 0, 16) {real, imag} */,
  {32'hc562ea9c, 32'h00000000} /* (10, 0, 15) {real, imag} */,
  {32'hc5a775a6, 32'h00000000} /* (10, 0, 14) {real, imag} */,
  {32'hc5cc937f, 32'h00000000} /* (10, 0, 13) {real, imag} */,
  {32'hc5adfd3e, 32'h00000000} /* (10, 0, 12) {real, imag} */,
  {32'hc5960776, 32'h00000000} /* (10, 0, 11) {real, imag} */,
  {32'hc5353c02, 32'h00000000} /* (10, 0, 10) {real, imag} */,
  {32'hc4c0cbb8, 32'h00000000} /* (10, 0, 9) {real, imag} */,
  {32'hc1b7f700, 32'h00000000} /* (10, 0, 8) {real, imag} */,
  {32'h44c5e360, 32'h00000000} /* (10, 0, 7) {real, imag} */,
  {32'h455696f4, 32'h00000000} /* (10, 0, 6) {real, imag} */,
  {32'h45c8384e, 32'h00000000} /* (10, 0, 5) {real, imag} */,
  {32'h4605ebc1, 32'h00000000} /* (10, 0, 4) {real, imag} */,
  {32'h462245a6, 32'h00000000} /* (10, 0, 3) {real, imag} */,
  {32'h462d8789, 32'h00000000} /* (10, 0, 2) {real, imag} */,
  {32'h4634b6b2, 32'h00000000} /* (10, 0, 1) {real, imag} */,
  {32'h4638e936, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h463b2aff, 32'h00000000} /* (9, 31, 31) {real, imag} */,
  {32'h463f221b, 32'h00000000} /* (9, 31, 30) {real, imag} */,
  {32'h4651f1f5, 32'h00000000} /* (9, 31, 29) {real, imag} */,
  {32'h464b8bce, 32'h00000000} /* (9, 31, 28) {real, imag} */,
  {32'h464c57ea, 32'h00000000} /* (9, 31, 27) {real, imag} */,
  {32'h464f2640, 32'h00000000} /* (9, 31, 26) {real, imag} */,
  {32'h4642e657, 32'h00000000} /* (9, 31, 25) {real, imag} */,
  {32'h463dbb11, 32'h00000000} /* (9, 31, 24) {real, imag} */,
  {32'h4625da46, 32'h00000000} /* (9, 31, 23) {real, imag} */,
  {32'h4610ce6f, 32'h00000000} /* (9, 31, 22) {real, imag} */,
  {32'h45da73c1, 32'h00000000} /* (9, 31, 21) {real, imag} */,
  {32'h457eb26c, 32'h00000000} /* (9, 31, 20) {real, imag} */,
  {32'h44f5edc0, 32'h00000000} /* (9, 31, 19) {real, imag} */,
  {32'h43a73470, 32'h00000000} /* (9, 31, 18) {real, imag} */,
  {32'hc4b1fc20, 32'h00000000} /* (9, 31, 17) {real, imag} */,
  {32'hc55ad174, 32'h00000000} /* (9, 31, 16) {real, imag} */,
  {32'hc59767ea, 32'h00000000} /* (9, 31, 15) {real, imag} */,
  {32'hc5c385a6, 32'h00000000} /* (9, 31, 14) {real, imag} */,
  {32'hc5cd6e4a, 32'h00000000} /* (9, 31, 13) {real, imag} */,
  {32'hc5af303b, 32'h00000000} /* (9, 31, 12) {real, imag} */,
  {32'hc53f309e, 32'h00000000} /* (9, 31, 11) {real, imag} */,
  {32'hc45b3a38, 32'h00000000} /* (9, 31, 10) {real, imag} */,
  {32'h4437c2d0, 32'h00000000} /* (9, 31, 9) {real, imag} */,
  {32'h4546c77c, 32'h00000000} /* (9, 31, 8) {real, imag} */,
  {32'h4594f7f8, 32'h00000000} /* (9, 31, 7) {real, imag} */,
  {32'h45c52bae, 32'h00000000} /* (9, 31, 6) {real, imag} */,
  {32'h45f665cf, 32'h00000000} /* (9, 31, 5) {real, imag} */,
  {32'h460d9ddc, 32'h00000000} /* (9, 31, 4) {real, imag} */,
  {32'h4622dd42, 32'h00000000} /* (9, 31, 3) {real, imag} */,
  {32'h462ef38e, 32'h00000000} /* (9, 31, 2) {real, imag} */,
  {32'h46315618, 32'h00000000} /* (9, 31, 1) {real, imag} */,
  {32'h4637b3e1, 32'h00000000} /* (9, 31, 0) {real, imag} */,
  {32'h463c6b18, 32'h00000000} /* (9, 30, 31) {real, imag} */,
  {32'h464c616c, 32'h00000000} /* (9, 30, 30) {real, imag} */,
  {32'h466151a0, 32'h00000000} /* (9, 30, 29) {real, imag} */,
  {32'h464bcdfc, 32'h00000000} /* (9, 30, 28) {real, imag} */,
  {32'h465b51f9, 32'h00000000} /* (9, 30, 27) {real, imag} */,
  {32'h464e6464, 32'h00000000} /* (9, 30, 26) {real, imag} */,
  {32'h463ee77a, 32'h00000000} /* (9, 30, 25) {real, imag} */,
  {32'h4643732e, 32'h00000000} /* (9, 30, 24) {real, imag} */,
  {32'h46205384, 32'h00000000} /* (9, 30, 23) {real, imag} */,
  {32'h4605b691, 32'h00000000} /* (9, 30, 22) {real, imag} */,
  {32'h45bb0102, 32'h00000000} /* (9, 30, 21) {real, imag} */,
  {32'h450a1cb4, 32'h00000000} /* (9, 30, 20) {real, imag} */,
  {32'h439b0c00, 32'h00000000} /* (9, 30, 19) {real, imag} */,
  {32'hc4fd8720, 32'h00000000} /* (9, 30, 18) {real, imag} */,
  {32'hc5604cd4, 32'h00000000} /* (9, 30, 17) {real, imag} */,
  {32'hc59f77c4, 32'h00000000} /* (9, 30, 16) {real, imag} */,
  {32'hc5c2fb68, 32'h00000000} /* (9, 30, 15) {real, imag} */,
  {32'hc5cb2994, 32'h00000000} /* (9, 30, 14) {real, imag} */,
  {32'hc5de7817, 32'h00000000} /* (9, 30, 13) {real, imag} */,
  {32'hc5b6dabb, 32'h00000000} /* (9, 30, 12) {real, imag} */,
  {32'hc5348014, 32'h00000000} /* (9, 30, 11) {real, imag} */,
  {32'h448398e4, 32'h00000000} /* (9, 30, 10) {real, imag} */,
  {32'h451ad984, 32'h00000000} /* (9, 30, 9) {real, imag} */,
  {32'h458acd29, 32'h00000000} /* (9, 30, 8) {real, imag} */,
  {32'h45e2b9ac, 32'h00000000} /* (9, 30, 7) {real, imag} */,
  {32'h45edeed2, 32'h00000000} /* (9, 30, 6) {real, imag} */,
  {32'h46174178, 32'h00000000} /* (9, 30, 5) {real, imag} */,
  {32'h462c0386, 32'h00000000} /* (9, 30, 4) {real, imag} */,
  {32'h463583fa, 32'h00000000} /* (9, 30, 3) {real, imag} */,
  {32'h4636fd27, 32'h00000000} /* (9, 30, 2) {real, imag} */,
  {32'h463e3a50, 32'h00000000} /* (9, 30, 1) {real, imag} */,
  {32'h464c344e, 32'h00000000} /* (9, 30, 0) {real, imag} */,
  {32'h464f476e, 32'h00000000} /* (9, 29, 31) {real, imag} */,
  {32'h465c83f2, 32'h00000000} /* (9, 29, 30) {real, imag} */,
  {32'h46514da4, 32'h00000000} /* (9, 29, 29) {real, imag} */,
  {32'h46548458, 32'h00000000} /* (9, 29, 28) {real, imag} */,
  {32'h464e4696, 32'h00000000} /* (9, 29, 27) {real, imag} */,
  {32'h46488e78, 32'h00000000} /* (9, 29, 26) {real, imag} */,
  {32'h4646af2c, 32'h00000000} /* (9, 29, 25) {real, imag} */,
  {32'h46365fc2, 32'h00000000} /* (9, 29, 24) {real, imag} */,
  {32'h461a9be0, 32'h00000000} /* (9, 29, 23) {real, imag} */,
  {32'h45fa7af4, 32'h00000000} /* (9, 29, 22) {real, imag} */,
  {32'h45a7fd32, 32'h00000000} /* (9, 29, 21) {real, imag} */,
  {32'h44c22320, 32'h00000000} /* (9, 29, 20) {real, imag} */,
  {32'hc4809ebc, 32'h00000000} /* (9, 29, 19) {real, imag} */,
  {32'hc54dd0ae, 32'h00000000} /* (9, 29, 18) {real, imag} */,
  {32'hc588f412, 32'h00000000} /* (9, 29, 17) {real, imag} */,
  {32'hc5caf094, 32'h00000000} /* (9, 29, 16) {real, imag} */,
  {32'hc6050252, 32'h00000000} /* (9, 29, 15) {real, imag} */,
  {32'hc5e7caac, 32'h00000000} /* (9, 29, 14) {real, imag} */,
  {32'hc5cd8df8, 32'h00000000} /* (9, 29, 13) {real, imag} */,
  {32'hc5a33347, 32'h00000000} /* (9, 29, 12) {real, imag} */,
  {32'hc5095644, 32'h00000000} /* (9, 29, 11) {real, imag} */,
  {32'h43c75570, 32'h00000000} /* (9, 29, 10) {real, imag} */,
  {32'h454aceb8, 32'h00000000} /* (9, 29, 9) {real, imag} */,
  {32'h45b84458, 32'h00000000} /* (9, 29, 8) {real, imag} */,
  {32'h45ed050c, 32'h00000000} /* (9, 29, 7) {real, imag} */,
  {32'h460d5ad6, 32'h00000000} /* (9, 29, 6) {real, imag} */,
  {32'h461b4fed, 32'h00000000} /* (9, 29, 5) {real, imag} */,
  {32'h463dc75f, 32'h00000000} /* (9, 29, 4) {real, imag} */,
  {32'h46499228, 32'h00000000} /* (9, 29, 3) {real, imag} */,
  {32'h463ec3ec, 32'h00000000} /* (9, 29, 2) {real, imag} */,
  {32'h46441a99, 32'h00000000} /* (9, 29, 1) {real, imag} */,
  {32'h46382194, 32'h00000000} /* (9, 29, 0) {real, imag} */,
  {32'h4656844b, 32'h00000000} /* (9, 28, 31) {real, imag} */,
  {32'h465b7602, 32'h00000000} /* (9, 28, 30) {real, imag} */,
  {32'h4648a666, 32'h00000000} /* (9, 28, 29) {real, imag} */,
  {32'h46489222, 32'h00000000} /* (9, 28, 28) {real, imag} */,
  {32'h464d0a08, 32'h00000000} /* (9, 28, 27) {real, imag} */,
  {32'h463d0334, 32'h00000000} /* (9, 28, 26) {real, imag} */,
  {32'h46387b0d, 32'h00000000} /* (9, 28, 25) {real, imag} */,
  {32'h46409615, 32'h00000000} /* (9, 28, 24) {real, imag} */,
  {32'h461dedc8, 32'h00000000} /* (9, 28, 23) {real, imag} */,
  {32'h460331dc, 32'h00000000} /* (9, 28, 22) {real, imag} */,
  {32'h456a8972, 32'h00000000} /* (9, 28, 21) {real, imag} */,
  {32'h441905a0, 32'h00000000} /* (9, 28, 20) {real, imag} */,
  {32'hc52e2fb2, 32'h00000000} /* (9, 28, 19) {real, imag} */,
  {32'hc58c5bb4, 32'h00000000} /* (9, 28, 18) {real, imag} */,
  {32'hc5c39a04, 32'h00000000} /* (9, 28, 17) {real, imag} */,
  {32'hc5e5e66c, 32'h00000000} /* (9, 28, 16) {real, imag} */,
  {32'hc60b3a7d, 32'h00000000} /* (9, 28, 15) {real, imag} */,
  {32'hc5f449a0, 32'h00000000} /* (9, 28, 14) {real, imag} */,
  {32'hc5c63030, 32'h00000000} /* (9, 28, 13) {real, imag} */,
  {32'hc591bf91, 32'h00000000} /* (9, 28, 12) {real, imag} */,
  {32'hc53c5122, 32'h00000000} /* (9, 28, 11) {real, imag} */,
  {32'h450a971a, 32'h00000000} /* (9, 28, 10) {real, imag} */,
  {32'h459a61b2, 32'h00000000} /* (9, 28, 9) {real, imag} */,
  {32'h45e1f70e, 32'h00000000} /* (9, 28, 8) {real, imag} */,
  {32'h4603aca4, 32'h00000000} /* (9, 28, 7) {real, imag} */,
  {32'h46151dc6, 32'h00000000} /* (9, 28, 6) {real, imag} */,
  {32'h4633c83c, 32'h00000000} /* (9, 28, 5) {real, imag} */,
  {32'h46403beb, 32'h00000000} /* (9, 28, 4) {real, imag} */,
  {32'h465484cc, 32'h00000000} /* (9, 28, 3) {real, imag} */,
  {32'h46414e90, 32'h00000000} /* (9, 28, 2) {real, imag} */,
  {32'h46473dd6, 32'h00000000} /* (9, 28, 1) {real, imag} */,
  {32'h46415f80, 32'h00000000} /* (9, 28, 0) {real, imag} */,
  {32'h46415c7c, 32'h00000000} /* (9, 27, 31) {real, imag} */,
  {32'h4649e438, 32'h00000000} /* (9, 27, 30) {real, imag} */,
  {32'h464ccb9d, 32'h00000000} /* (9, 27, 29) {real, imag} */,
  {32'h46430178, 32'h00000000} /* (9, 27, 28) {real, imag} */,
  {32'h464a25fa, 32'h00000000} /* (9, 27, 27) {real, imag} */,
  {32'h4642a20e, 32'h00000000} /* (9, 27, 26) {real, imag} */,
  {32'h4658b600, 32'h00000000} /* (9, 27, 25) {real, imag} */,
  {32'h4630deb2, 32'h00000000} /* (9, 27, 24) {real, imag} */,
  {32'h46148c53, 32'h00000000} /* (9, 27, 23) {real, imag} */,
  {32'h45d0892c, 32'h00000000} /* (9, 27, 22) {real, imag} */,
  {32'h45228f68, 32'h00000000} /* (9, 27, 21) {real, imag} */,
  {32'hc4b7164c, 32'h00000000} /* (9, 27, 20) {real, imag} */,
  {32'hc545b23c, 32'h00000000} /* (9, 27, 19) {real, imag} */,
  {32'hc5a38b31, 32'h00000000} /* (9, 27, 18) {real, imag} */,
  {32'hc5cc3708, 32'h00000000} /* (9, 27, 17) {real, imag} */,
  {32'hc5ff2f0c, 32'h00000000} /* (9, 27, 16) {real, imag} */,
  {32'hc60189fe, 32'h00000000} /* (9, 27, 15) {real, imag} */,
  {32'hc5da6287, 32'h00000000} /* (9, 27, 14) {real, imag} */,
  {32'hc5cf0736, 32'h00000000} /* (9, 27, 13) {real, imag} */,
  {32'hc59012b4, 32'h00000000} /* (9, 27, 12) {real, imag} */,
  {32'hc524e176, 32'h00000000} /* (9, 27, 11) {real, imag} */,
  {32'h44edd564, 32'h00000000} /* (9, 27, 10) {real, imag} */,
  {32'h459f74e3, 32'h00000000} /* (9, 27, 9) {real, imag} */,
  {32'h45effc6d, 32'h00000000} /* (9, 27, 8) {real, imag} */,
  {32'h4620dd63, 32'h00000000} /* (9, 27, 7) {real, imag} */,
  {32'h4627a25a, 32'h00000000} /* (9, 27, 6) {real, imag} */,
  {32'h46413f50, 32'h00000000} /* (9, 27, 5) {real, imag} */,
  {32'h46444a98, 32'h00000000} /* (9, 27, 4) {real, imag} */,
  {32'h4647a0da, 32'h00000000} /* (9, 27, 3) {real, imag} */,
  {32'h464489f2, 32'h00000000} /* (9, 27, 2) {real, imag} */,
  {32'h4649c452, 32'h00000000} /* (9, 27, 1) {real, imag} */,
  {32'h46434732, 32'h00000000} /* (9, 27, 0) {real, imag} */,
  {32'h46388b23, 32'h00000000} /* (9, 26, 31) {real, imag} */,
  {32'h46412f4a, 32'h00000000} /* (9, 26, 30) {real, imag} */,
  {32'h4652400a, 32'h00000000} /* (9, 26, 29) {real, imag} */,
  {32'h464bd55b, 32'h00000000} /* (9, 26, 28) {real, imag} */,
  {32'h4636f278, 32'h00000000} /* (9, 26, 27) {real, imag} */,
  {32'h4642f11f, 32'h00000000} /* (9, 26, 26) {real, imag} */,
  {32'h463cff99, 32'h00000000} /* (9, 26, 25) {real, imag} */,
  {32'h46300e03, 32'h00000000} /* (9, 26, 24) {real, imag} */,
  {32'h45fc48df, 32'h00000000} /* (9, 26, 23) {real, imag} */,
  {32'h45b78674, 32'h00000000} /* (9, 26, 22) {real, imag} */,
  {32'h4552f324, 32'h00000000} /* (9, 26, 21) {real, imag} */,
  {32'hc4bc5fa0, 32'h00000000} /* (9, 26, 20) {real, imag} */,
  {32'hc592a858, 32'h00000000} /* (9, 26, 19) {real, imag} */,
  {32'hc5af8b4c, 32'h00000000} /* (9, 26, 18) {real, imag} */,
  {32'hc5d4819e, 32'h00000000} /* (9, 26, 17) {real, imag} */,
  {32'hc5fb4a3c, 32'h00000000} /* (9, 26, 16) {real, imag} */,
  {32'hc5f4655a, 32'h00000000} /* (9, 26, 15) {real, imag} */,
  {32'hc5d839c8, 32'h00000000} /* (9, 26, 14) {real, imag} */,
  {32'hc5b87d31, 32'h00000000} /* (9, 26, 13) {real, imag} */,
  {32'hc578ba54, 32'h00000000} /* (9, 26, 12) {real, imag} */,
  {32'hc4695f48, 32'h00000000} /* (9, 26, 11) {real, imag} */,
  {32'h44f8b148, 32'h00000000} /* (9, 26, 10) {real, imag} */,
  {32'h45b84f6a, 32'h00000000} /* (9, 26, 9) {real, imag} */,
  {32'h45fca8c1, 32'h00000000} /* (9, 26, 8) {real, imag} */,
  {32'h46114edf, 32'h00000000} /* (9, 26, 7) {real, imag} */,
  {32'h462c3cb0, 32'h00000000} /* (9, 26, 6) {real, imag} */,
  {32'h4633058a, 32'h00000000} /* (9, 26, 5) {real, imag} */,
  {32'h463f69f6, 32'h00000000} /* (9, 26, 4) {real, imag} */,
  {32'h463f1a58, 32'h00000000} /* (9, 26, 3) {real, imag} */,
  {32'h464135f2, 32'h00000000} /* (9, 26, 2) {real, imag} */,
  {32'h46435639, 32'h00000000} /* (9, 26, 1) {real, imag} */,
  {32'h4639baae, 32'h00000000} /* (9, 26, 0) {real, imag} */,
  {32'h462b2b9c, 32'h00000000} /* (9, 25, 31) {real, imag} */,
  {32'h463353b8, 32'h00000000} /* (9, 25, 30) {real, imag} */,
  {32'h463d1c11, 32'h00000000} /* (9, 25, 29) {real, imag} */,
  {32'h464e6351, 32'h00000000} /* (9, 25, 28) {real, imag} */,
  {32'h4626fce8, 32'h00000000} /* (9, 25, 27) {real, imag} */,
  {32'h462762bc, 32'h00000000} /* (9, 25, 26) {real, imag} */,
  {32'h4624e99a, 32'h00000000} /* (9, 25, 25) {real, imag} */,
  {32'h46132b3e, 32'h00000000} /* (9, 25, 24) {real, imag} */,
  {32'h45e5ec47, 32'h00000000} /* (9, 25, 23) {real, imag} */,
  {32'h45936d69, 32'h00000000} /* (9, 25, 22) {real, imag} */,
  {32'h451bf826, 32'h00000000} /* (9, 25, 21) {real, imag} */,
  {32'hc4c511b8, 32'h00000000} /* (9, 25, 20) {real, imag} */,
  {32'hc56b5afe, 32'h00000000} /* (9, 25, 19) {real, imag} */,
  {32'hc5baaa3c, 32'h00000000} /* (9, 25, 18) {real, imag} */,
  {32'hc5e56943, 32'h00000000} /* (9, 25, 17) {real, imag} */,
  {32'hc5dfbf39, 32'h00000000} /* (9, 25, 16) {real, imag} */,
  {32'hc5db2690, 32'h00000000} /* (9, 25, 15) {real, imag} */,
  {32'hc5cb9ca8, 32'h00000000} /* (9, 25, 14) {real, imag} */,
  {32'hc5b57092, 32'h00000000} /* (9, 25, 13) {real, imag} */,
  {32'hc53f39e4, 32'h00000000} /* (9, 25, 12) {real, imag} */,
  {32'hc4c64aa8, 32'h00000000} /* (9, 25, 11) {real, imag} */,
  {32'h45181328, 32'h00000000} /* (9, 25, 10) {real, imag} */,
  {32'h45cfb5a4, 32'h00000000} /* (9, 25, 9) {real, imag} */,
  {32'h45e55254, 32'h00000000} /* (9, 25, 8) {real, imag} */,
  {32'h460b1a9c, 32'h00000000} /* (9, 25, 7) {real, imag} */,
  {32'h462bbf14, 32'h00000000} /* (9, 25, 6) {real, imag} */,
  {32'h46382132, 32'h00000000} /* (9, 25, 5) {real, imag} */,
  {32'h46395a87, 32'h00000000} /* (9, 25, 4) {real, imag} */,
  {32'h463ca324, 32'h00000000} /* (9, 25, 3) {real, imag} */,
  {32'h463169d4, 32'h00000000} /* (9, 25, 2) {real, imag} */,
  {32'h46357f4c, 32'h00000000} /* (9, 25, 1) {real, imag} */,
  {32'h462d58bc, 32'h00000000} /* (9, 25, 0) {real, imag} */,
  {32'h46116f54, 32'h00000000} /* (9, 24, 31) {real, imag} */,
  {32'h462d204f, 32'h00000000} /* (9, 24, 30) {real, imag} */,
  {32'h4615f47e, 32'h00000000} /* (9, 24, 29) {real, imag} */,
  {32'h4612df20, 32'h00000000} /* (9, 24, 28) {real, imag} */,
  {32'h4614124f, 32'h00000000} /* (9, 24, 27) {real, imag} */,
  {32'h4613a858, 32'h00000000} /* (9, 24, 26) {real, imag} */,
  {32'h460a8e60, 32'h00000000} /* (9, 24, 25) {real, imag} */,
  {32'h45ee8efd, 32'h00000000} /* (9, 24, 24) {real, imag} */,
  {32'h45bc6db9, 32'h00000000} /* (9, 24, 23) {real, imag} */,
  {32'h45606c82, 32'h00000000} /* (9, 24, 22) {real, imag} */,
  {32'h44ac695c, 32'h00000000} /* (9, 24, 21) {real, imag} */,
  {32'hc5067756, 32'h00000000} /* (9, 24, 20) {real, imag} */,
  {32'hc56f1012, 32'h00000000} /* (9, 24, 19) {real, imag} */,
  {32'hc589a999, 32'h00000000} /* (9, 24, 18) {real, imag} */,
  {32'hc589bcc2, 32'h00000000} /* (9, 24, 17) {real, imag} */,
  {32'hc5b8b3d4, 32'h00000000} /* (9, 24, 16) {real, imag} */,
  {32'hc5d9e233, 32'h00000000} /* (9, 24, 15) {real, imag} */,
  {32'hc5ac005a, 32'h00000000} /* (9, 24, 14) {real, imag} */,
  {32'hc5933c27, 32'h00000000} /* (9, 24, 13) {real, imag} */,
  {32'hc58d902c, 32'h00000000} /* (9, 24, 12) {real, imag} */,
  {32'hc50538c8, 32'h00000000} /* (9, 24, 11) {real, imag} */,
  {32'h456ae8a2, 32'h00000000} /* (9, 24, 10) {real, imag} */,
  {32'h45b5a390, 32'h00000000} /* (9, 24, 9) {real, imag} */,
  {32'h45e2aad9, 32'h00000000} /* (9, 24, 8) {real, imag} */,
  {32'h460a351c, 32'h00000000} /* (9, 24, 7) {real, imag} */,
  {32'h46124174, 32'h00000000} /* (9, 24, 6) {real, imag} */,
  {32'h462200a4, 32'h00000000} /* (9, 24, 5) {real, imag} */,
  {32'h462046f8, 32'h00000000} /* (9, 24, 4) {real, imag} */,
  {32'h46214788, 32'h00000000} /* (9, 24, 3) {real, imag} */,
  {32'h461fdcda, 32'h00000000} /* (9, 24, 2) {real, imag} */,
  {32'h46143b67, 32'h00000000} /* (9, 24, 1) {real, imag} */,
  {32'h460d37f7, 32'h00000000} /* (9, 24, 0) {real, imag} */,
  {32'h45e477dc, 32'h00000000} /* (9, 23, 31) {real, imag} */,
  {32'h45ef11d4, 32'h00000000} /* (9, 23, 30) {real, imag} */,
  {32'h45f717e4, 32'h00000000} /* (9, 23, 29) {real, imag} */,
  {32'h45fa4d68, 32'h00000000} /* (9, 23, 28) {real, imag} */,
  {32'h45fb17b8, 32'h00000000} /* (9, 23, 27) {real, imag} */,
  {32'h45e4a36c, 32'h00000000} /* (9, 23, 26) {real, imag} */,
  {32'h45c7a7e9, 32'h00000000} /* (9, 23, 25) {real, imag} */,
  {32'h45c633b8, 32'h00000000} /* (9, 23, 24) {real, imag} */,
  {32'h45c5996a, 32'h00000000} /* (9, 23, 23) {real, imag} */,
  {32'h455749b1, 32'h00000000} /* (9, 23, 22) {real, imag} */,
  {32'h449a06fc, 32'h00000000} /* (9, 23, 21) {real, imag} */,
  {32'hc4aa8d0a, 32'h00000000} /* (9, 23, 20) {real, imag} */,
  {32'hc5672607, 32'h00000000} /* (9, 23, 19) {real, imag} */,
  {32'hc57fb1b3, 32'h00000000} /* (9, 23, 18) {real, imag} */,
  {32'hc58cac12, 32'h00000000} /* (9, 23, 17) {real, imag} */,
  {32'hc58fe289, 32'h00000000} /* (9, 23, 16) {real, imag} */,
  {32'hc5954c7a, 32'h00000000} /* (9, 23, 15) {real, imag} */,
  {32'hc592470c, 32'h00000000} /* (9, 23, 14) {real, imag} */,
  {32'hc57e1cbf, 32'h00000000} /* (9, 23, 13) {real, imag} */,
  {32'hc533bcdf, 32'h00000000} /* (9, 23, 12) {real, imag} */,
  {32'hc4f1aea2, 32'h00000000} /* (9, 23, 11) {real, imag} */,
  {32'h4516a738, 32'h00000000} /* (9, 23, 10) {real, imag} */,
  {32'h4585513f, 32'h00000000} /* (9, 23, 9) {real, imag} */,
  {32'h45ce73bc, 32'h00000000} /* (9, 23, 8) {real, imag} */,
  {32'h45de9b86, 32'h00000000} /* (9, 23, 7) {real, imag} */,
  {32'h45ef77c4, 32'h00000000} /* (9, 23, 6) {real, imag} */,
  {32'h45eb243d, 32'h00000000} /* (9, 23, 5) {real, imag} */,
  {32'h46027d3c, 32'h00000000} /* (9, 23, 4) {real, imag} */,
  {32'h45fddd30, 32'h00000000} /* (9, 23, 3) {real, imag} */,
  {32'h45f4427e, 32'h00000000} /* (9, 23, 2) {real, imag} */,
  {32'h45f7f410, 32'h00000000} /* (9, 23, 1) {real, imag} */,
  {32'h45dd2587, 32'h00000000} /* (9, 23, 0) {real, imag} */,
  {32'h45900f65, 32'h00000000} /* (9, 22, 31) {real, imag} */,
  {32'h45b188ef, 32'h00000000} /* (9, 22, 30) {real, imag} */,
  {32'h45ce8d47, 32'h00000000} /* (9, 22, 29) {real, imag} */,
  {32'h45c37ade, 32'h00000000} /* (9, 22, 28) {real, imag} */,
  {32'h459bfb56, 32'h00000000} /* (9, 22, 27) {real, imag} */,
  {32'h45a81aef, 32'h00000000} /* (9, 22, 26) {real, imag} */,
  {32'h45a50a93, 32'h00000000} /* (9, 22, 25) {real, imag} */,
  {32'h458edbd7, 32'h00000000} /* (9, 22, 24) {real, imag} */,
  {32'h4598678d, 32'h00000000} /* (9, 22, 23) {real, imag} */,
  {32'h4530ab6e, 32'h00000000} /* (9, 22, 22) {real, imag} */,
  {32'h44a4fffe, 32'h00000000} /* (9, 22, 21) {real, imag} */,
  {32'hc4a5d0fc, 32'h00000000} /* (9, 22, 20) {real, imag} */,
  {32'hc500caa0, 32'h00000000} /* (9, 22, 19) {real, imag} */,
  {32'hc57e0e46, 32'h00000000} /* (9, 22, 18) {real, imag} */,
  {32'hc54bad7d, 32'h00000000} /* (9, 22, 17) {real, imag} */,
  {32'hc52ba6b1, 32'h00000000} /* (9, 22, 16) {real, imag} */,
  {32'hc5234c02, 32'h00000000} /* (9, 22, 15) {real, imag} */,
  {32'hc545bbd2, 32'h00000000} /* (9, 22, 14) {real, imag} */,
  {32'hc520517e, 32'h00000000} /* (9, 22, 13) {real, imag} */,
  {32'hc4d65f5c, 32'h00000000} /* (9, 22, 12) {real, imag} */,
  {32'hc219a040, 32'h00000000} /* (9, 22, 11) {real, imag} */,
  {32'h44be3623, 32'h00000000} /* (9, 22, 10) {real, imag} */,
  {32'h453a3472, 32'h00000000} /* (9, 22, 9) {real, imag} */,
  {32'h4568906a, 32'h00000000} /* (9, 22, 8) {real, imag} */,
  {32'h45817cad, 32'h00000000} /* (9, 22, 7) {real, imag} */,
  {32'h459d66cd, 32'h00000000} /* (9, 22, 6) {real, imag} */,
  {32'h45af0844, 32'h00000000} /* (9, 22, 5) {real, imag} */,
  {32'h45aeb740, 32'h00000000} /* (9, 22, 4) {real, imag} */,
  {32'h45c3d3f4, 32'h00000000} /* (9, 22, 3) {real, imag} */,
  {32'h45c5f821, 32'h00000000} /* (9, 22, 2) {real, imag} */,
  {32'h45a18786, 32'h00000000} /* (9, 22, 1) {real, imag} */,
  {32'h458c296e, 32'h00000000} /* (9, 22, 0) {real, imag} */,
  {32'h44e90226, 32'h00000000} /* (9, 21, 31) {real, imag} */,
  {32'h44f8584c, 32'h00000000} /* (9, 21, 30) {real, imag} */,
  {32'h44eeb9be, 32'h00000000} /* (9, 21, 29) {real, imag} */,
  {32'h44e2c395, 32'h00000000} /* (9, 21, 28) {real, imag} */,
  {32'h44d3fd7c, 32'h00000000} /* (9, 21, 27) {real, imag} */,
  {32'h451629c8, 32'h00000000} /* (9, 21, 26) {real, imag} */,
  {32'h451cbabe, 32'h00000000} /* (9, 21, 25) {real, imag} */,
  {32'h44f21ea6, 32'h00000000} /* (9, 21, 24) {real, imag} */,
  {32'h44b4ad4e, 32'h00000000} /* (9, 21, 23) {real, imag} */,
  {32'h4492404d, 32'h00000000} /* (9, 21, 22) {real, imag} */,
  {32'h45058848, 32'h00000000} /* (9, 21, 21) {real, imag} */,
  {32'hc4abceb6, 32'h00000000} /* (9, 21, 20) {real, imag} */,
  {32'hc4b5c1ba, 32'h00000000} /* (9, 21, 19) {real, imag} */,
  {32'hc421e818, 32'h00000000} /* (9, 21, 18) {real, imag} */,
  {32'hc42c00e7, 32'h00000000} /* (9, 21, 17) {real, imag} */,
  {32'h441354d9, 32'h00000000} /* (9, 21, 16) {real, imag} */,
  {32'hc426295c, 32'h00000000} /* (9, 21, 15) {real, imag} */,
  {32'hc27e50c0, 32'h00000000} /* (9, 21, 14) {real, imag} */,
  {32'h41ec8880, 32'h00000000} /* (9, 21, 13) {real, imag} */,
  {32'h4390aa14, 32'h00000000} /* (9, 21, 12) {real, imag} */,
  {32'hc354e464, 32'h00000000} /* (9, 21, 11) {real, imag} */,
  {32'h44a528d4, 32'h00000000} /* (9, 21, 10) {real, imag} */,
  {32'h449c78d3, 32'h00000000} /* (9, 21, 9) {real, imag} */,
  {32'h448c7cc6, 32'h00000000} /* (9, 21, 8) {real, imag} */,
  {32'h44b60cda, 32'h00000000} /* (9, 21, 7) {real, imag} */,
  {32'h44a53fe5, 32'h00000000} /* (9, 21, 6) {real, imag} */,
  {32'h4501902e, 32'h00000000} /* (9, 21, 5) {real, imag} */,
  {32'h4501b1ad, 32'h00000000} /* (9, 21, 4) {real, imag} */,
  {32'h44df7ca8, 32'h00000000} /* (9, 21, 3) {real, imag} */,
  {32'h4553bffc, 32'h00000000} /* (9, 21, 2) {real, imag} */,
  {32'h44d618e8, 32'h00000000} /* (9, 21, 1) {real, imag} */,
  {32'h44afd0b8, 32'h00000000} /* (9, 21, 0) {real, imag} */,
  {32'hc4f9f147, 32'h00000000} /* (9, 20, 31) {real, imag} */,
  {32'hc50bd9ac, 32'h00000000} /* (9, 20, 30) {real, imag} */,
  {32'hc52137b6, 32'h00000000} /* (9, 20, 29) {real, imag} */,
  {32'hc50a5517, 32'h00000000} /* (9, 20, 28) {real, imag} */,
  {32'hc4ce13a2, 32'h00000000} /* (9, 20, 27) {real, imag} */,
  {32'hc4e0647c, 32'h00000000} /* (9, 20, 26) {real, imag} */,
  {32'hc50abf5d, 32'h00000000} /* (9, 20, 25) {real, imag} */,
  {32'hc4f6cabc, 32'h00000000} /* (9, 20, 24) {real, imag} */,
  {32'hc4b09d96, 32'h00000000} /* (9, 20, 23) {real, imag} */,
  {32'hc3e97f8e, 32'h00000000} /* (9, 20, 22) {real, imag} */,
  {32'hc3ab7680, 32'h00000000} /* (9, 20, 21) {real, imag} */,
  {32'h44daaea0, 32'h00000000} /* (9, 20, 20) {real, imag} */,
  {32'h44645f87, 32'h00000000} /* (9, 20, 19) {real, imag} */,
  {32'h44af07c8, 32'h00000000} /* (9, 20, 18) {real, imag} */,
  {32'h4516e082, 32'h00000000} /* (9, 20, 17) {real, imag} */,
  {32'h453780cb, 32'h00000000} /* (9, 20, 16) {real, imag} */,
  {32'h453dbef8, 32'h00000000} /* (9, 20, 15) {real, imag} */,
  {32'h453b1976, 32'h00000000} /* (9, 20, 14) {real, imag} */,
  {32'h45465420, 32'h00000000} /* (9, 20, 13) {real, imag} */,
  {32'h45352bfb, 32'h00000000} /* (9, 20, 12) {real, imag} */,
  {32'h44cb3642, 32'h00000000} /* (9, 20, 11) {real, imag} */,
  {32'h426d08d0, 32'h00000000} /* (9, 20, 10) {real, imag} */,
  {32'hc4be4a72, 32'h00000000} /* (9, 20, 9) {real, imag} */,
  {32'hc4ee52ac, 32'h00000000} /* (9, 20, 8) {real, imag} */,
  {32'hc51a365c, 32'h00000000} /* (9, 20, 7) {real, imag} */,
  {32'hc51a732e, 32'h00000000} /* (9, 20, 6) {real, imag} */,
  {32'hc4cfa74c, 32'h00000000} /* (9, 20, 5) {real, imag} */,
  {32'hc5122a56, 32'h00000000} /* (9, 20, 4) {real, imag} */,
  {32'hc52aeac0, 32'h00000000} /* (9, 20, 3) {real, imag} */,
  {32'hc506254a, 32'h00000000} /* (9, 20, 2) {real, imag} */,
  {32'hc5397bac, 32'h00000000} /* (9, 20, 1) {real, imag} */,
  {32'hc4ec1826, 32'h00000000} /* (9, 20, 0) {real, imag} */,
  {32'hc5a29a89, 32'h00000000} /* (9, 19, 31) {real, imag} */,
  {32'hc5b282ea, 32'h00000000} /* (9, 19, 30) {real, imag} */,
  {32'hc59fe4fb, 32'h00000000} /* (9, 19, 29) {real, imag} */,
  {32'hc5900bbe, 32'h00000000} /* (9, 19, 28) {real, imag} */,
  {32'hc59cad9b, 32'h00000000} /* (9, 19, 27) {real, imag} */,
  {32'hc59fb164, 32'h00000000} /* (9, 19, 26) {real, imag} */,
  {32'hc5763a4a, 32'h00000000} /* (9, 19, 25) {real, imag} */,
  {32'hc592989a, 32'h00000000} /* (9, 19, 24) {real, imag} */,
  {32'hc57520c1, 32'h00000000} /* (9, 19, 23) {real, imag} */,
  {32'hc543bf4b, 32'h00000000} /* (9, 19, 22) {real, imag} */,
  {32'hc43027d8, 32'h00000000} /* (9, 19, 21) {real, imag} */,
  {32'h44ea20fc, 32'h00000000} /* (9, 19, 20) {real, imag} */,
  {32'h453219c6, 32'h00000000} /* (9, 19, 19) {real, imag} */,
  {32'h455a5ebe, 32'h00000000} /* (9, 19, 18) {real, imag} */,
  {32'h457d43b6, 32'h00000000} /* (9, 19, 17) {real, imag} */,
  {32'h45b99de0, 32'h00000000} /* (9, 19, 16) {real, imag} */,
  {32'h45b8b0f9, 32'h00000000} /* (9, 19, 15) {real, imag} */,
  {32'h45c6509c, 32'h00000000} /* (9, 19, 14) {real, imag} */,
  {32'h45914df1, 32'h00000000} /* (9, 19, 13) {real, imag} */,
  {32'h454b387b, 32'h00000000} /* (9, 19, 12) {real, imag} */,
  {32'h45197b7e, 32'h00000000} /* (9, 19, 11) {real, imag} */,
  {32'hc48174c0, 32'h00000000} /* (9, 19, 10) {real, imag} */,
  {32'hc529a36a, 32'h00000000} /* (9, 19, 9) {real, imag} */,
  {32'hc59641ec, 32'h00000000} /* (9, 19, 8) {real, imag} */,
  {32'hc5a802d6, 32'h00000000} /* (9, 19, 7) {real, imag} */,
  {32'hc5aae50a, 32'h00000000} /* (9, 19, 6) {real, imag} */,
  {32'hc5aebdc9, 32'h00000000} /* (9, 19, 5) {real, imag} */,
  {32'hc5a7764f, 32'h00000000} /* (9, 19, 4) {real, imag} */,
  {32'hc5afa957, 32'h00000000} /* (9, 19, 3) {real, imag} */,
  {32'hc5a9dab7, 32'h00000000} /* (9, 19, 2) {real, imag} */,
  {32'hc5a756a9, 32'h00000000} /* (9, 19, 1) {real, imag} */,
  {32'hc58adc7e, 32'h00000000} /* (9, 19, 0) {real, imag} */,
  {32'hc5ee7e01, 32'h00000000} /* (9, 18, 31) {real, imag} */,
  {32'hc5eccf8e, 32'h00000000} /* (9, 18, 30) {real, imag} */,
  {32'hc5f1d8e8, 32'h00000000} /* (9, 18, 29) {real, imag} */,
  {32'hc5e4b738, 32'h00000000} /* (9, 18, 28) {real, imag} */,
  {32'hc5dbed1c, 32'h00000000} /* (9, 18, 27) {real, imag} */,
  {32'hc5cb4134, 32'h00000000} /* (9, 18, 26) {real, imag} */,
  {32'hc5caecc4, 32'h00000000} /* (9, 18, 25) {real, imag} */,
  {32'hc5cfd390, 32'h00000000} /* (9, 18, 24) {real, imag} */,
  {32'hc5ae2e5e, 32'h00000000} /* (9, 18, 23) {real, imag} */,
  {32'hc533a865, 32'h00000000} /* (9, 18, 22) {real, imag} */,
  {32'hc480aecc, 32'h00000000} /* (9, 18, 21) {real, imag} */,
  {32'h453a9228, 32'h00000000} /* (9, 18, 20) {real, imag} */,
  {32'h4580ac3a, 32'h00000000} /* (9, 18, 19) {real, imag} */,
  {32'h458ce080, 32'h00000000} /* (9, 18, 18) {real, imag} */,
  {32'h45b289a4, 32'h00000000} /* (9, 18, 17) {real, imag} */,
  {32'h45fab7ce, 32'h00000000} /* (9, 18, 16) {real, imag} */,
  {32'h45e27187, 32'h00000000} /* (9, 18, 15) {real, imag} */,
  {32'h45d63cb2, 32'h00000000} /* (9, 18, 14) {real, imag} */,
  {32'h45cdabd6, 32'h00000000} /* (9, 18, 13) {real, imag} */,
  {32'h45962408, 32'h00000000} /* (9, 18, 12) {real, imag} */,
  {32'h45083465, 32'h00000000} /* (9, 18, 11) {real, imag} */,
  {32'hc491a6ea, 32'h00000000} /* (9, 18, 10) {real, imag} */,
  {32'hc5789ee8, 32'h00000000} /* (9, 18, 9) {real, imag} */,
  {32'hc59d7cbc, 32'h00000000} /* (9, 18, 8) {real, imag} */,
  {32'hc5b75ec8, 32'h00000000} /* (9, 18, 7) {real, imag} */,
  {32'hc5d27c1e, 32'h00000000} /* (9, 18, 6) {real, imag} */,
  {32'hc5e02eb9, 32'h00000000} /* (9, 18, 5) {real, imag} */,
  {32'hc5f331dc, 32'h00000000} /* (9, 18, 4) {real, imag} */,
  {32'hc5fded88, 32'h00000000} /* (9, 18, 3) {real, imag} */,
  {32'hc5e67e02, 32'h00000000} /* (9, 18, 2) {real, imag} */,
  {32'hc5f1ce80, 32'h00000000} /* (9, 18, 1) {real, imag} */,
  {32'hc5e15734, 32'h00000000} /* (9, 18, 0) {real, imag} */,
  {32'hc609a6dd, 32'h00000000} /* (9, 17, 31) {real, imag} */,
  {32'hc61576c5, 32'h00000000} /* (9, 17, 30) {real, imag} */,
  {32'hc615d612, 32'h00000000} /* (9, 17, 29) {real, imag} */,
  {32'hc616d588, 32'h00000000} /* (9, 17, 28) {real, imag} */,
  {32'hc60eff52, 32'h00000000} /* (9, 17, 27) {real, imag} */,
  {32'hc603c070, 32'h00000000} /* (9, 17, 26) {real, imag} */,
  {32'hc5ed2931, 32'h00000000} /* (9, 17, 25) {real, imag} */,
  {32'hc5fd3466, 32'h00000000} /* (9, 17, 24) {real, imag} */,
  {32'hc5c7f6d8, 32'h00000000} /* (9, 17, 23) {real, imag} */,
  {32'hc552d7df, 32'h00000000} /* (9, 17, 22) {real, imag} */,
  {32'hc40d5998, 32'h00000000} /* (9, 17, 21) {real, imag} */,
  {32'h455f861d, 32'h00000000} /* (9, 17, 20) {real, imag} */,
  {32'h4599d91f, 32'h00000000} /* (9, 17, 19) {real, imag} */,
  {32'h45a4dc05, 32'h00000000} /* (9, 17, 18) {real, imag} */,
  {32'h45e95a92, 32'h00000000} /* (9, 17, 17) {real, imag} */,
  {32'h45e1fcac, 32'h00000000} /* (9, 17, 16) {real, imag} */,
  {32'h45e6ed84, 32'h00000000} /* (9, 17, 15) {real, imag} */,
  {32'h45d17c6e, 32'h00000000} /* (9, 17, 14) {real, imag} */,
  {32'h45c70e82, 32'h00000000} /* (9, 17, 13) {real, imag} */,
  {32'h45873440, 32'h00000000} /* (9, 17, 12) {real, imag} */,
  {32'h44ee0728, 32'h00000000} /* (9, 17, 11) {real, imag} */,
  {32'hc4b294c6, 32'h00000000} /* (9, 17, 10) {real, imag} */,
  {32'hc59307d5, 32'h00000000} /* (9, 17, 9) {real, imag} */,
  {32'hc5cc4f7e, 32'h00000000} /* (9, 17, 8) {real, imag} */,
  {32'hc5cd1832, 32'h00000000} /* (9, 17, 7) {real, imag} */,
  {32'hc5f2a6d0, 32'h00000000} /* (9, 17, 6) {real, imag} */,
  {32'hc6092b14, 32'h00000000} /* (9, 17, 5) {real, imag} */,
  {32'hc60705ee, 32'h00000000} /* (9, 17, 4) {real, imag} */,
  {32'hc613637e, 32'h00000000} /* (9, 17, 3) {real, imag} */,
  {32'hc61a8684, 32'h00000000} /* (9, 17, 2) {real, imag} */,
  {32'hc6064077, 32'h00000000} /* (9, 17, 1) {real, imag} */,
  {32'hc5fbd460, 32'h00000000} /* (9, 17, 0) {real, imag} */,
  {32'hc60bbb68, 32'h00000000} /* (9, 16, 31) {real, imag} */,
  {32'hc623cc65, 32'h00000000} /* (9, 16, 30) {real, imag} */,
  {32'hc617680f, 32'h00000000} /* (9, 16, 29) {real, imag} */,
  {32'hc622f57a, 32'h00000000} /* (9, 16, 28) {real, imag} */,
  {32'hc614fac6, 32'h00000000} /* (9, 16, 27) {real, imag} */,
  {32'hc60853fc, 32'h00000000} /* (9, 16, 26) {real, imag} */,
  {32'hc602c113, 32'h00000000} /* (9, 16, 25) {real, imag} */,
  {32'hc5e11b26, 32'h00000000} /* (9, 16, 24) {real, imag} */,
  {32'hc5c2e2c7, 32'h00000000} /* (9, 16, 23) {real, imag} */,
  {32'hc57f4227, 32'h00000000} /* (9, 16, 22) {real, imag} */,
  {32'hc3e1cb80, 32'h00000000} /* (9, 16, 21) {real, imag} */,
  {32'h451d261e, 32'h00000000} /* (9, 16, 20) {real, imag} */,
  {32'h458da052, 32'h00000000} /* (9, 16, 19) {real, imag} */,
  {32'h45d24dd8, 32'h00000000} /* (9, 16, 18) {real, imag} */,
  {32'h45eea070, 32'h00000000} /* (9, 16, 17) {real, imag} */,
  {32'h46023706, 32'h00000000} /* (9, 16, 16) {real, imag} */,
  {32'h4600113a, 32'h00000000} /* (9, 16, 15) {real, imag} */,
  {32'h45e409ba, 32'h00000000} /* (9, 16, 14) {real, imag} */,
  {32'h45b6eca6, 32'h00000000} /* (9, 16, 13) {real, imag} */,
  {32'h458b8037, 32'h00000000} /* (9, 16, 12) {real, imag} */,
  {32'h44b9a2b0, 32'h00000000} /* (9, 16, 11) {real, imag} */,
  {32'hc4f3cc10, 32'h00000000} /* (9, 16, 10) {real, imag} */,
  {32'hc586f3b3, 32'h00000000} /* (9, 16, 9) {real, imag} */,
  {32'hc5cf3526, 32'h00000000} /* (9, 16, 8) {real, imag} */,
  {32'hc5e754b9, 32'h00000000} /* (9, 16, 7) {real, imag} */,
  {32'hc5f77ea2, 32'h00000000} /* (9, 16, 6) {real, imag} */,
  {32'hc60a5923, 32'h00000000} /* (9, 16, 5) {real, imag} */,
  {32'hc60d2ade, 32'h00000000} /* (9, 16, 4) {real, imag} */,
  {32'hc620763e, 32'h00000000} /* (9, 16, 3) {real, imag} */,
  {32'hc618700c, 32'h00000000} /* (9, 16, 2) {real, imag} */,
  {32'hc60dbc6a, 32'h00000000} /* (9, 16, 1) {real, imag} */,
  {32'hc601316e, 32'h00000000} /* (9, 16, 0) {real, imag} */,
  {32'hc60557fd, 32'h00000000} /* (9, 15, 31) {real, imag} */,
  {32'hc618f91b, 32'h00000000} /* (9, 15, 30) {real, imag} */,
  {32'hc612f77e, 32'h00000000} /* (9, 15, 29) {real, imag} */,
  {32'hc60f97fd, 32'h00000000} /* (9, 15, 28) {real, imag} */,
  {32'hc614bb4a, 32'h00000000} /* (9, 15, 27) {real, imag} */,
  {32'hc608a25e, 32'h00000000} /* (9, 15, 26) {real, imag} */,
  {32'hc60297e3, 32'h00000000} /* (9, 15, 25) {real, imag} */,
  {32'hc5e8c1bd, 32'h00000000} /* (9, 15, 24) {real, imag} */,
  {32'hc5b393ba, 32'h00000000} /* (9, 15, 23) {real, imag} */,
  {32'hc5685b42, 32'h00000000} /* (9, 15, 22) {real, imag} */,
  {32'hc3944038, 32'h00000000} /* (9, 15, 21) {real, imag} */,
  {32'h45302fce, 32'h00000000} /* (9, 15, 20) {real, imag} */,
  {32'h45949a43, 32'h00000000} /* (9, 15, 19) {real, imag} */,
  {32'h45d4bfc6, 32'h00000000} /* (9, 15, 18) {real, imag} */,
  {32'h45ebf5fc, 32'h00000000} /* (9, 15, 17) {real, imag} */,
  {32'h4602807c, 32'h00000000} /* (9, 15, 16) {real, imag} */,
  {32'h45f372da, 32'h00000000} /* (9, 15, 15) {real, imag} */,
  {32'h45d3cf52, 32'h00000000} /* (9, 15, 14) {real, imag} */,
  {32'h45c4c507, 32'h00000000} /* (9, 15, 13) {real, imag} */,
  {32'h459dcfdc, 32'h00000000} /* (9, 15, 12) {real, imag} */,
  {32'h4501c37a, 32'h00000000} /* (9, 15, 11) {real, imag} */,
  {32'hc4e751de, 32'h00000000} /* (9, 15, 10) {real, imag} */,
  {32'hc581008e, 32'h00000000} /* (9, 15, 9) {real, imag} */,
  {32'hc5ccea85, 32'h00000000} /* (9, 15, 8) {real, imag} */,
  {32'hc5ee6f1a, 32'h00000000} /* (9, 15, 7) {real, imag} */,
  {32'hc602e800, 32'h00000000} /* (9, 15, 6) {real, imag} */,
  {32'hc60297f5, 32'h00000000} /* (9, 15, 5) {real, imag} */,
  {32'hc60fae36, 32'h00000000} /* (9, 15, 4) {real, imag} */,
  {32'hc617ba94, 32'h00000000} /* (9, 15, 3) {real, imag} */,
  {32'hc617be65, 32'h00000000} /* (9, 15, 2) {real, imag} */,
  {32'hc60f3014, 32'h00000000} /* (9, 15, 1) {real, imag} */,
  {32'hc60de194, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'hc60189c2, 32'h00000000} /* (9, 14, 31) {real, imag} */,
  {32'hc60c3870, 32'h00000000} /* (9, 14, 30) {real, imag} */,
  {32'hc5fadee6, 32'h00000000} /* (9, 14, 29) {real, imag} */,
  {32'hc600224c, 32'h00000000} /* (9, 14, 28) {real, imag} */,
  {32'hc61c513c, 32'h00000000} /* (9, 14, 27) {real, imag} */,
  {32'hc6022970, 32'h00000000} /* (9, 14, 26) {real, imag} */,
  {32'hc5fb63db, 32'h00000000} /* (9, 14, 25) {real, imag} */,
  {32'hc5c72028, 32'h00000000} /* (9, 14, 24) {real, imag} */,
  {32'hc59d3be9, 32'h00000000} /* (9, 14, 23) {real, imag} */,
  {32'hc54bb9b4, 32'h00000000} /* (9, 14, 22) {real, imag} */,
  {32'hc417e8a4, 32'h00000000} /* (9, 14, 21) {real, imag} */,
  {32'h45301372, 32'h00000000} /* (9, 14, 20) {real, imag} */,
  {32'h457c67f7, 32'h00000000} /* (9, 14, 19) {real, imag} */,
  {32'h45acec16, 32'h00000000} /* (9, 14, 18) {real, imag} */,
  {32'h45cea910, 32'h00000000} /* (9, 14, 17) {real, imag} */,
  {32'h45db62ee, 32'h00000000} /* (9, 14, 16) {real, imag} */,
  {32'h45d3b642, 32'h00000000} /* (9, 14, 15) {real, imag} */,
  {32'h45d9e8f4, 32'h00000000} /* (9, 14, 14) {real, imag} */,
  {32'h45d7a41c, 32'h00000000} /* (9, 14, 13) {real, imag} */,
  {32'h4592b619, 32'h00000000} /* (9, 14, 12) {real, imag} */,
  {32'h44fa39ea, 32'h00000000} /* (9, 14, 11) {real, imag} */,
  {32'hc4998f40, 32'h00000000} /* (9, 14, 10) {real, imag} */,
  {32'hc5909065, 32'h00000000} /* (9, 14, 9) {real, imag} */,
  {32'hc5c326ac, 32'h00000000} /* (9, 14, 8) {real, imag} */,
  {32'hc5d8d10b, 32'h00000000} /* (9, 14, 7) {real, imag} */,
  {32'hc5e84994, 32'h00000000} /* (9, 14, 6) {real, imag} */,
  {32'hc5f8497c, 32'h00000000} /* (9, 14, 5) {real, imag} */,
  {32'hc5f837b9, 32'h00000000} /* (9, 14, 4) {real, imag} */,
  {32'hc5fc337e, 32'h00000000} /* (9, 14, 3) {real, imag} */,
  {32'hc6082a7c, 32'h00000000} /* (9, 14, 2) {real, imag} */,
  {32'hc603209a, 32'h00000000} /* (9, 14, 1) {real, imag} */,
  {32'hc5eb1a10, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hc5cbcbfc, 32'h00000000} /* (9, 13, 31) {real, imag} */,
  {32'hc5d16727, 32'h00000000} /* (9, 13, 30) {real, imag} */,
  {32'hc5da2c08, 32'h00000000} /* (9, 13, 29) {real, imag} */,
  {32'hc5ed5a96, 32'h00000000} /* (9, 13, 28) {real, imag} */,
  {32'hc5c51f5c, 32'h00000000} /* (9, 13, 27) {real, imag} */,
  {32'hc5ce7dbe, 32'h00000000} /* (9, 13, 26) {real, imag} */,
  {32'hc5bf4842, 32'h00000000} /* (9, 13, 25) {real, imag} */,
  {32'hc5a6ba1a, 32'h00000000} /* (9, 13, 24) {real, imag} */,
  {32'hc58b7ae0, 32'h00000000} /* (9, 13, 23) {real, imag} */,
  {32'hc513b496, 32'h00000000} /* (9, 13, 22) {real, imag} */,
  {32'hc2c6b360, 32'h00000000} /* (9, 13, 21) {real, imag} */,
  {32'h4544012e, 32'h00000000} /* (9, 13, 20) {real, imag} */,
  {32'h45689b33, 32'h00000000} /* (9, 13, 19) {real, imag} */,
  {32'h45b2cdb5, 32'h00000000} /* (9, 13, 18) {real, imag} */,
  {32'h45b66fc8, 32'h00000000} /* (9, 13, 17) {real, imag} */,
  {32'h45ab54c2, 32'h00000000} /* (9, 13, 16) {real, imag} */,
  {32'h45af3d34, 32'h00000000} /* (9, 13, 15) {real, imag} */,
  {32'h45a5ac29, 32'h00000000} /* (9, 13, 14) {real, imag} */,
  {32'h45b3061c, 32'h00000000} /* (9, 13, 13) {real, imag} */,
  {32'h455e6bf4, 32'h00000000} /* (9, 13, 12) {real, imag} */,
  {32'h44d8dd2e, 32'h00000000} /* (9, 13, 11) {real, imag} */,
  {32'hc4f33c22, 32'h00000000} /* (9, 13, 10) {real, imag} */,
  {32'hc5943cb2, 32'h00000000} /* (9, 13, 9) {real, imag} */,
  {32'hc5ab1a42, 32'h00000000} /* (9, 13, 8) {real, imag} */,
  {32'hc5d86370, 32'h00000000} /* (9, 13, 7) {real, imag} */,
  {32'hc5c13669, 32'h00000000} /* (9, 13, 6) {real, imag} */,
  {32'hc5d7bc74, 32'h00000000} /* (9, 13, 5) {real, imag} */,
  {32'hc5dc3073, 32'h00000000} /* (9, 13, 4) {real, imag} */,
  {32'hc5eade10, 32'h00000000} /* (9, 13, 3) {real, imag} */,
  {32'hc5ce02a1, 32'h00000000} /* (9, 13, 2) {real, imag} */,
  {32'hc5d7fd20, 32'h00000000} /* (9, 13, 1) {real, imag} */,
  {32'hc5e01e52, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'hc588db62, 32'h00000000} /* (9, 12, 31) {real, imag} */,
  {32'hc5a4e773, 32'h00000000} /* (9, 12, 30) {real, imag} */,
  {32'hc59e9588, 32'h00000000} /* (9, 12, 29) {real, imag} */,
  {32'hc599b46c, 32'h00000000} /* (9, 12, 28) {real, imag} */,
  {32'hc5994d1a, 32'h00000000} /* (9, 12, 27) {real, imag} */,
  {32'hc58c35ac, 32'h00000000} /* (9, 12, 26) {real, imag} */,
  {32'hc57eb774, 32'h00000000} /* (9, 12, 25) {real, imag} */,
  {32'hc563368d, 32'h00000000} /* (9, 12, 24) {real, imag} */,
  {32'hc51d640d, 32'h00000000} /* (9, 12, 23) {real, imag} */,
  {32'hc4b4164a, 32'h00000000} /* (9, 12, 22) {real, imag} */,
  {32'h445cafe4, 32'h00000000} /* (9, 12, 21) {real, imag} */,
  {32'h45281482, 32'h00000000} /* (9, 12, 20) {real, imag} */,
  {32'h4582a053, 32'h00000000} /* (9, 12, 19) {real, imag} */,
  {32'h456ee25e, 32'h00000000} /* (9, 12, 18) {real, imag} */,
  {32'h458b948c, 32'h00000000} /* (9, 12, 17) {real, imag} */,
  {32'h459da4b2, 32'h00000000} /* (9, 12, 16) {real, imag} */,
  {32'h458bfb7e, 32'h00000000} /* (9, 12, 15) {real, imag} */,
  {32'h458d6e59, 32'h00000000} /* (9, 12, 14) {real, imag} */,
  {32'h453ad519, 32'h00000000} /* (9, 12, 13) {real, imag} */,
  {32'h453a6ccc, 32'h00000000} /* (9, 12, 12) {real, imag} */,
  {32'h4433b49c, 32'h00000000} /* (9, 12, 11) {real, imag} */,
  {32'hc4ef79da, 32'h00000000} /* (9, 12, 10) {real, imag} */,
  {32'hc582e39a, 32'h00000000} /* (9, 12, 9) {real, imag} */,
  {32'hc57211d3, 32'h00000000} /* (9, 12, 8) {real, imag} */,
  {32'hc59e12a8, 32'h00000000} /* (9, 12, 7) {real, imag} */,
  {32'hc5b25b16, 32'h00000000} /* (9, 12, 6) {real, imag} */,
  {32'hc59bdd6c, 32'h00000000} /* (9, 12, 5) {real, imag} */,
  {32'hc5a0f7c8, 32'h00000000} /* (9, 12, 4) {real, imag} */,
  {32'hc5a11b27, 32'h00000000} /* (9, 12, 3) {real, imag} */,
  {32'hc5966093, 32'h00000000} /* (9, 12, 2) {real, imag} */,
  {32'hc5900758, 32'h00000000} /* (9, 12, 1) {real, imag} */,
  {32'hc5926964, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'hc48c56d2, 32'h00000000} /* (9, 11, 31) {real, imag} */,
  {32'hc4b8c2da, 32'h00000000} /* (9, 11, 30) {real, imag} */,
  {32'hc4b12fef, 32'h00000000} /* (9, 11, 29) {real, imag} */,
  {32'hc4a2ea58, 32'h00000000} /* (9, 11, 28) {real, imag} */,
  {32'hc50d04f6, 32'h00000000} /* (9, 11, 27) {real, imag} */,
  {32'hc49b5962, 32'h00000000} /* (9, 11, 26) {real, imag} */,
  {32'hc4a11a6c, 32'h00000000} /* (9, 11, 25) {real, imag} */,
  {32'hc4af2617, 32'h00000000} /* (9, 11, 24) {real, imag} */,
  {32'hc38af2f4, 32'h00000000} /* (9, 11, 23) {real, imag} */,
  {32'h4418d374, 32'h00000000} /* (9, 11, 22) {real, imag} */,
  {32'h4443428a, 32'h00000000} /* (9, 11, 21) {real, imag} */,
  {32'h4524a7fd, 32'h00000000} /* (9, 11, 20) {real, imag} */,
  {32'h451aa5a9, 32'h00000000} /* (9, 11, 19) {real, imag} */,
  {32'h45085626, 32'h00000000} /* (9, 11, 18) {real, imag} */,
  {32'h451f1618, 32'h00000000} /* (9, 11, 17) {real, imag} */,
  {32'h4529c012, 32'h00000000} /* (9, 11, 16) {real, imag} */,
  {32'h451be9a8, 32'h00000000} /* (9, 11, 15) {real, imag} */,
  {32'h452bbac5, 32'h00000000} /* (9, 11, 14) {real, imag} */,
  {32'h44f65eaf, 32'h00000000} /* (9, 11, 13) {real, imag} */,
  {32'h44a32b5c, 32'h00000000} /* (9, 11, 12) {real, imag} */,
  {32'hc3e3676c, 32'h00000000} /* (9, 11, 11) {real, imag} */,
  {32'hc4c6d480, 32'h00000000} /* (9, 11, 10) {real, imag} */,
  {32'hc4bba698, 32'h00000000} /* (9, 11, 9) {real, imag} */,
  {32'hc50f217b, 32'h00000000} /* (9, 11, 8) {real, imag} */,
  {32'hc52984b2, 32'h00000000} /* (9, 11, 7) {real, imag} */,
  {32'hc50d10f9, 32'h00000000} /* (9, 11, 6) {real, imag} */,
  {32'hc4d4bc7d, 32'h00000000} /* (9, 11, 5) {real, imag} */,
  {32'hc50766c5, 32'h00000000} /* (9, 11, 4) {real, imag} */,
  {32'hc4ddad8e, 32'h00000000} /* (9, 11, 3) {real, imag} */,
  {32'hc50ef45c, 32'h00000000} /* (9, 11, 2) {real, imag} */,
  {32'hc5229aa2, 32'h00000000} /* (9, 11, 1) {real, imag} */,
  {32'hc4972f9e, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h4508a910, 32'h00000000} /* (9, 10, 31) {real, imag} */,
  {32'h4508ee3f, 32'h00000000} /* (9, 10, 30) {real, imag} */,
  {32'h455e2724, 32'h00000000} /* (9, 10, 29) {real, imag} */,
  {32'h452c9946, 32'h00000000} /* (9, 10, 28) {real, imag} */,
  {32'h4540e8eb, 32'h00000000} /* (9, 10, 27) {real, imag} */,
  {32'h45155b11, 32'h00000000} /* (9, 10, 26) {real, imag} */,
  {32'h452308ea, 32'h00000000} /* (9, 10, 25) {real, imag} */,
  {32'h45230e5c, 32'h00000000} /* (9, 10, 24) {real, imag} */,
  {32'h4528fc75, 32'h00000000} /* (9, 10, 23) {real, imag} */,
  {32'h458284ed, 32'h00000000} /* (9, 10, 22) {real, imag} */,
  {32'h451bf0e8, 32'h00000000} /* (9, 10, 21) {real, imag} */,
  {32'h44c8e5aa, 32'h00000000} /* (9, 10, 20) {real, imag} */,
  {32'h442fa84e, 32'h00000000} /* (9, 10, 19) {real, imag} */,
  {32'hc43ac0e6, 32'h00000000} /* (9, 10, 18) {real, imag} */,
  {32'h43b9a83e, 32'h00000000} /* (9, 10, 17) {real, imag} */,
  {32'hc458a7a9, 32'h00000000} /* (9, 10, 16) {real, imag} */,
  {32'hc42e2865, 32'h00000000} /* (9, 10, 15) {real, imag} */,
  {32'hc499dfaa, 32'h00000000} /* (9, 10, 14) {real, imag} */,
  {32'hc47023f8, 32'h00000000} /* (9, 10, 13) {real, imag} */,
  {32'hc4cc0fcb, 32'h00000000} /* (9, 10, 12) {real, imag} */,
  {32'hc488456e, 32'h00000000} /* (9, 10, 11) {real, imag} */,
  {32'hc46cdb9c, 32'h00000000} /* (9, 10, 10) {real, imag} */,
  {32'hc31d9858, 32'h00000000} /* (9, 10, 9) {real, imag} */,
  {32'hc38c21c0, 32'h00000000} /* (9, 10, 8) {real, imag} */,
  {32'h446259bd, 32'h00000000} /* (9, 10, 7) {real, imag} */,
  {32'h44beb5b1, 32'h00000000} /* (9, 10, 6) {real, imag} */,
  {32'h450ef98e, 32'h00000000} /* (9, 10, 5) {real, imag} */,
  {32'h44e2fa64, 32'h00000000} /* (9, 10, 4) {real, imag} */,
  {32'h44a2996d, 32'h00000000} /* (9, 10, 3) {real, imag} */,
  {32'h4476cca2, 32'h00000000} /* (9, 10, 2) {real, imag} */,
  {32'h448b03c2, 32'h00000000} /* (9, 10, 1) {real, imag} */,
  {32'h4503725a, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'h45964cea, 32'h00000000} /* (9, 9, 31) {real, imag} */,
  {32'h45b497da, 32'h00000000} /* (9, 9, 30) {real, imag} */,
  {32'h45c80832, 32'h00000000} /* (9, 9, 29) {real, imag} */,
  {32'h45cc1460, 32'h00000000} /* (9, 9, 28) {real, imag} */,
  {32'h45d455cf, 32'h00000000} /* (9, 9, 27) {real, imag} */,
  {32'h45b709e4, 32'h00000000} /* (9, 9, 26) {real, imag} */,
  {32'h45b4dcee, 32'h00000000} /* (9, 9, 25) {real, imag} */,
  {32'h45bf2876, 32'h00000000} /* (9, 9, 24) {real, imag} */,
  {32'h45bb9ca4, 32'h00000000} /* (9, 9, 23) {real, imag} */,
  {32'h459694e0, 32'h00000000} /* (9, 9, 22) {real, imag} */,
  {32'h45805d23, 32'h00000000} /* (9, 9, 21) {real, imag} */,
  {32'h44ef7172, 32'h00000000} /* (9, 9, 20) {real, imag} */,
  {32'h43b02e70, 32'h00000000} /* (9, 9, 19) {real, imag} */,
  {32'hc509a79b, 32'h00000000} /* (9, 9, 18) {real, imag} */,
  {32'hc52fbc88, 32'h00000000} /* (9, 9, 17) {real, imag} */,
  {32'hc5350ed6, 32'h00000000} /* (9, 9, 16) {real, imag} */,
  {32'hc550ccc4, 32'h00000000} /* (9, 9, 15) {real, imag} */,
  {32'hc55ef514, 32'h00000000} /* (9, 9, 14) {real, imag} */,
  {32'hc57a9fdc, 32'h00000000} /* (9, 9, 13) {real, imag} */,
  {32'hc56dc950, 32'h00000000} /* (9, 9, 12) {real, imag} */,
  {32'hc51801ba, 32'h00000000} /* (9, 9, 11) {real, imag} */,
  {32'hc4192b7c, 32'h00000000} /* (9, 9, 10) {real, imag} */,
  {32'h438066d8, 32'h00000000} /* (9, 9, 9) {real, imag} */,
  {32'h449f7bfe, 32'h00000000} /* (9, 9, 8) {real, imag} */,
  {32'h4519e0ed, 32'h00000000} /* (9, 9, 7) {real, imag} */,
  {32'h4565cd48, 32'h00000000} /* (9, 9, 6) {real, imag} */,
  {32'h45910ef1, 32'h00000000} /* (9, 9, 5) {real, imag} */,
  {32'h45816a6e, 32'h00000000} /* (9, 9, 4) {real, imag} */,
  {32'h458f2b85, 32'h00000000} /* (9, 9, 3) {real, imag} */,
  {32'h458956b8, 32'h00000000} /* (9, 9, 2) {real, imag} */,
  {32'h45816708, 32'h00000000} /* (9, 9, 1) {real, imag} */,
  {32'h4587fae6, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h45e3f7c3, 32'h00000000} /* (9, 8, 31) {real, imag} */,
  {32'h45ee0a5a, 32'h00000000} /* (9, 8, 30) {real, imag} */,
  {32'h460fd818, 32'h00000000} /* (9, 8, 29) {real, imag} */,
  {32'h460aee74, 32'h00000000} /* (9, 8, 28) {real, imag} */,
  {32'h460f8b0d, 32'h00000000} /* (9, 8, 27) {real, imag} */,
  {32'h4606689a, 32'h00000000} /* (9, 8, 26) {real, imag} */,
  {32'h46014182, 32'h00000000} /* (9, 8, 25) {real, imag} */,
  {32'h46061896, 32'h00000000} /* (9, 8, 24) {real, imag} */,
  {32'h4600ee49, 32'h00000000} /* (9, 8, 23) {real, imag} */,
  {32'h45d84078, 32'h00000000} /* (9, 8, 22) {real, imag} */,
  {32'h4591b520, 32'h00000000} /* (9, 8, 21) {real, imag} */,
  {32'h44f41b02, 32'h00000000} /* (9, 8, 20) {real, imag} */,
  {32'h444579a4, 32'h00000000} /* (9, 8, 19) {real, imag} */,
  {32'hc4cc8e8c, 32'h00000000} /* (9, 8, 18) {real, imag} */,
  {32'hc54f5059, 32'h00000000} /* (9, 8, 17) {real, imag} */,
  {32'hc586bca4, 32'h00000000} /* (9, 8, 16) {real, imag} */,
  {32'hc598d2c1, 32'h00000000} /* (9, 8, 15) {real, imag} */,
  {32'hc59dea70, 32'h00000000} /* (9, 8, 14) {real, imag} */,
  {32'hc59c4f42, 32'h00000000} /* (9, 8, 13) {real, imag} */,
  {32'hc58e6515, 32'h00000000} /* (9, 8, 12) {real, imag} */,
  {32'hc5433431, 32'h00000000} /* (9, 8, 11) {real, imag} */,
  {32'hc3ec6ef0, 32'h00000000} /* (9, 8, 10) {real, imag} */,
  {32'h44830434, 32'h00000000} /* (9, 8, 9) {real, imag} */,
  {32'h454af21a, 32'h00000000} /* (9, 8, 8) {real, imag} */,
  {32'h459c14b9, 32'h00000000} /* (9, 8, 7) {real, imag} */,
  {32'h45b7b9c8, 32'h00000000} /* (9, 8, 6) {real, imag} */,
  {32'h45b416bc, 32'h00000000} /* (9, 8, 5) {real, imag} */,
  {32'h45cf7aa2, 32'h00000000} /* (9, 8, 4) {real, imag} */,
  {32'h45caa574, 32'h00000000} /* (9, 8, 3) {real, imag} */,
  {32'h45d07083, 32'h00000000} /* (9, 8, 2) {real, imag} */,
  {32'h45d30498, 32'h00000000} /* (9, 8, 1) {real, imag} */,
  {32'h45c592bc, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h460561ce, 32'h00000000} /* (9, 7, 31) {real, imag} */,
  {32'h460d0c2d, 32'h00000000} /* (9, 7, 30) {real, imag} */,
  {32'h462140c8, 32'h00000000} /* (9, 7, 29) {real, imag} */,
  {32'h462a86e4, 32'h00000000} /* (9, 7, 28) {real, imag} */,
  {32'h4620246e, 32'h00000000} /* (9, 7, 27) {real, imag} */,
  {32'h4622254e, 32'h00000000} /* (9, 7, 26) {real, imag} */,
  {32'h461a75cd, 32'h00000000} /* (9, 7, 25) {real, imag} */,
  {32'h46158bf8, 32'h00000000} /* (9, 7, 24) {real, imag} */,
  {32'h46142b06, 32'h00000000} /* (9, 7, 23) {real, imag} */,
  {32'h46059e42, 32'h00000000} /* (9, 7, 22) {real, imag} */,
  {32'h45bd742e, 32'h00000000} /* (9, 7, 21) {real, imag} */,
  {32'h4548c656, 32'h00000000} /* (9, 7, 20) {real, imag} */,
  {32'h443d6534, 32'h00000000} /* (9, 7, 19) {real, imag} */,
  {32'hc484d340, 32'h00000000} /* (9, 7, 18) {real, imag} */,
  {32'hc5614ff6, 32'h00000000} /* (9, 7, 17) {real, imag} */,
  {32'hc57a1cce, 32'h00000000} /* (9, 7, 16) {real, imag} */,
  {32'hc5a6ba29, 32'h00000000} /* (9, 7, 15) {real, imag} */,
  {32'hc5bb653a, 32'h00000000} /* (9, 7, 14) {real, imag} */,
  {32'hc5c1ffec, 32'h00000000} /* (9, 7, 13) {real, imag} */,
  {32'hc5bd7f64, 32'h00000000} /* (9, 7, 12) {real, imag} */,
  {32'hc58147a8, 32'h00000000} /* (9, 7, 11) {real, imag} */,
  {32'hc4858220, 32'h00000000} /* (9, 7, 10) {real, imag} */,
  {32'h44ed74b0, 32'h00000000} /* (9, 7, 9) {real, imag} */,
  {32'h454f1e34, 32'h00000000} /* (9, 7, 8) {real, imag} */,
  {32'h459ba173, 32'h00000000} /* (9, 7, 7) {real, imag} */,
  {32'h45b829f9, 32'h00000000} /* (9, 7, 6) {real, imag} */,
  {32'h45d86b16, 32'h00000000} /* (9, 7, 5) {real, imag} */,
  {32'h46043618, 32'h00000000} /* (9, 7, 4) {real, imag} */,
  {32'h45f84d52, 32'h00000000} /* (9, 7, 3) {real, imag} */,
  {32'h460a7338, 32'h00000000} /* (9, 7, 2) {real, imag} */,
  {32'h460e2912, 32'h00000000} /* (9, 7, 1) {real, imag} */,
  {32'h4607464e, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h4619d6c7, 32'h00000000} /* (9, 6, 31) {real, imag} */,
  {32'h461d0773, 32'h00000000} /* (9, 6, 30) {real, imag} */,
  {32'h4633a488, 32'h00000000} /* (9, 6, 29) {real, imag} */,
  {32'h463b5eb7, 32'h00000000} /* (9, 6, 28) {real, imag} */,
  {32'h46337664, 32'h00000000} /* (9, 6, 27) {real, imag} */,
  {32'h462db054, 32'h00000000} /* (9, 6, 26) {real, imag} */,
  {32'h462bc328, 32'h00000000} /* (9, 6, 25) {real, imag} */,
  {32'h4634b776, 32'h00000000} /* (9, 6, 24) {real, imag} */,
  {32'h46356ca6, 32'h00000000} /* (9, 6, 23) {real, imag} */,
  {32'h4614346b, 32'h00000000} /* (9, 6, 22) {real, imag} */,
  {32'h45eb4729, 32'h00000000} /* (9, 6, 21) {real, imag} */,
  {32'h4594f560, 32'h00000000} /* (9, 6, 20) {real, imag} */,
  {32'h450ad5b7, 32'h00000000} /* (9, 6, 19) {real, imag} */,
  {32'hc3ca92d0, 32'h00000000} /* (9, 6, 18) {real, imag} */,
  {32'hc4f16e28, 32'h00000000} /* (9, 6, 17) {real, imag} */,
  {32'hc56cb8a4, 32'h00000000} /* (9, 6, 16) {real, imag} */,
  {32'hc5b44ca4, 32'h00000000} /* (9, 6, 15) {real, imag} */,
  {32'hc5bc401e, 32'h00000000} /* (9, 6, 14) {real, imag} */,
  {32'hc5db13b0, 32'h00000000} /* (9, 6, 13) {real, imag} */,
  {32'hc5c5435a, 32'h00000000} /* (9, 6, 12) {real, imag} */,
  {32'hc5987348, 32'h00000000} /* (9, 6, 11) {real, imag} */,
  {32'hc5096a1c, 32'h00000000} /* (9, 6, 10) {real, imag} */,
  {32'h434a98a0, 32'h00000000} /* (9, 6, 9) {real, imag} */,
  {32'h44c78044, 32'h00000000} /* (9, 6, 8) {real, imag} */,
  {32'h458299f8, 32'h00000000} /* (9, 6, 7) {real, imag} */,
  {32'h45aa083a, 32'h00000000} /* (9, 6, 6) {real, imag} */,
  {32'h46096ea6, 32'h00000000} /* (9, 6, 5) {real, imag} */,
  {32'h4600bcbc, 32'h00000000} /* (9, 6, 4) {real, imag} */,
  {32'h460ce3ca, 32'h00000000} /* (9, 6, 3) {real, imag} */,
  {32'h4617e206, 32'h00000000} /* (9, 6, 2) {real, imag} */,
  {32'h4624ab68, 32'h00000000} /* (9, 6, 1) {real, imag} */,
  {32'h461dac75, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'h462c383e, 32'h00000000} /* (9, 5, 31) {real, imag} */,
  {32'h46320b94, 32'h00000000} /* (9, 5, 30) {real, imag} */,
  {32'h463887e0, 32'h00000000} /* (9, 5, 29) {real, imag} */,
  {32'h464c219e, 32'h00000000} /* (9, 5, 28) {real, imag} */,
  {32'h46426d4f, 32'h00000000} /* (9, 5, 27) {real, imag} */,
  {32'h46523226, 32'h00000000} /* (9, 5, 26) {real, imag} */,
  {32'h463e5e84, 32'h00000000} /* (9, 5, 25) {real, imag} */,
  {32'h463841ce, 32'h00000000} /* (9, 5, 24) {real, imag} */,
  {32'h463d4af8, 32'h00000000} /* (9, 5, 23) {real, imag} */,
  {32'h462c0ed8, 32'h00000000} /* (9, 5, 22) {real, imag} */,
  {32'h460cc92a, 32'h00000000} /* (9, 5, 21) {real, imag} */,
  {32'h45ee8521, 32'h00000000} /* (9, 5, 20) {real, imag} */,
  {32'h458bb724, 32'h00000000} /* (9, 5, 19) {real, imag} */,
  {32'h44e77494, 32'h00000000} /* (9, 5, 18) {real, imag} */,
  {32'h44a98d14, 32'h00000000} /* (9, 5, 17) {real, imag} */,
  {32'hc4f3c95c, 32'h00000000} /* (9, 5, 16) {real, imag} */,
  {32'hc58fdb30, 32'h00000000} /* (9, 5, 15) {real, imag} */,
  {32'hc5b80825, 32'h00000000} /* (9, 5, 14) {real, imag} */,
  {32'hc5bf6f78, 32'h00000000} /* (9, 5, 13) {real, imag} */,
  {32'hc5d46333, 32'h00000000} /* (9, 5, 12) {real, imag} */,
  {32'hc5cc4982, 32'h00000000} /* (9, 5, 11) {real, imag} */,
  {32'hc5606ade, 32'h00000000} /* (9, 5, 10) {real, imag} */,
  {32'hc5124e82, 32'h00000000} /* (9, 5, 9) {real, imag} */,
  {32'hc28fe140, 32'h00000000} /* (9, 5, 8) {real, imag} */,
  {32'h44db224c, 32'h00000000} /* (9, 5, 7) {real, imag} */,
  {32'h45a402c6, 32'h00000000} /* (9, 5, 6) {real, imag} */,
  {32'h45e8363c, 32'h00000000} /* (9, 5, 5) {real, imag} */,
  {32'h45f02fb1, 32'h00000000} /* (9, 5, 4) {real, imag} */,
  {32'h4621ab70, 32'h00000000} /* (9, 5, 3) {real, imag} */,
  {32'h462513f6, 32'h00000000} /* (9, 5, 2) {real, imag} */,
  {32'h463843a6, 32'h00000000} /* (9, 5, 1) {real, imag} */,
  {32'h4637f1ae, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'h463f6dee, 32'h00000000} /* (9, 4, 31) {real, imag} */,
  {32'h46401d6f, 32'h00000000} /* (9, 4, 30) {real, imag} */,
  {32'h465031e5, 32'h00000000} /* (9, 4, 29) {real, imag} */,
  {32'h46507606, 32'h00000000} /* (9, 4, 28) {real, imag} */,
  {32'h466886b4, 32'h00000000} /* (9, 4, 27) {real, imag} */,
  {32'h465d4320, 32'h00000000} /* (9, 4, 26) {real, imag} */,
  {32'h46484b6e, 32'h00000000} /* (9, 4, 25) {real, imag} */,
  {32'h4644fdf7, 32'h00000000} /* (9, 4, 24) {real, imag} */,
  {32'h463c5382, 32'h00000000} /* (9, 4, 23) {real, imag} */,
  {32'h46350262, 32'h00000000} /* (9, 4, 22) {real, imag} */,
  {32'h46136484, 32'h00000000} /* (9, 4, 21) {real, imag} */,
  {32'h4608737e, 32'h00000000} /* (9, 4, 20) {real, imag} */,
  {32'h45cd7157, 32'h00000000} /* (9, 4, 19) {real, imag} */,
  {32'h457ac211, 32'h00000000} /* (9, 4, 18) {real, imag} */,
  {32'h44ebabc0, 32'h00000000} /* (9, 4, 17) {real, imag} */,
  {32'hc484ab60, 32'h00000000} /* (9, 4, 16) {real, imag} */,
  {32'hc57ac13a, 32'h00000000} /* (9, 4, 15) {real, imag} */,
  {32'hc59f8482, 32'h00000000} /* (9, 4, 14) {real, imag} */,
  {32'hc5c693de, 32'h00000000} /* (9, 4, 13) {real, imag} */,
  {32'hc5f806af, 32'h00000000} /* (9, 4, 12) {real, imag} */,
  {32'hc5d183a9, 32'h00000000} /* (9, 4, 11) {real, imag} */,
  {32'hc5968273, 32'h00000000} /* (9, 4, 10) {real, imag} */,
  {32'hc5353e0e, 32'h00000000} /* (9, 4, 9) {real, imag} */,
  {32'hc4c1b520, 32'h00000000} /* (9, 4, 8) {real, imag} */,
  {32'h43d24840, 32'h00000000} /* (9, 4, 7) {real, imag} */,
  {32'h44c96d20, 32'h00000000} /* (9, 4, 6) {real, imag} */,
  {32'h45a8a998, 32'h00000000} /* (9, 4, 5) {real, imag} */,
  {32'h4604caee, 32'h00000000} /* (9, 4, 4) {real, imag} */,
  {32'h4619b698, 32'h00000000} /* (9, 4, 3) {real, imag} */,
  {32'h462fd45d, 32'h00000000} /* (9, 4, 2) {real, imag} */,
  {32'h463475a7, 32'h00000000} /* (9, 4, 1) {real, imag} */,
  {32'h463f2aeb, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'h46376e36, 32'h00000000} /* (9, 3, 31) {real, imag} */,
  {32'h464f161a, 32'h00000000} /* (9, 3, 30) {real, imag} */,
  {32'h4658d7e8, 32'h00000000} /* (9, 3, 29) {real, imag} */,
  {32'h4654fb74, 32'h00000000} /* (9, 3, 28) {real, imag} */,
  {32'h4661488e, 32'h00000000} /* (9, 3, 27) {real, imag} */,
  {32'h465cacb6, 32'h00000000} /* (9, 3, 26) {real, imag} */,
  {32'h465c0808, 32'h00000000} /* (9, 3, 25) {real, imag} */,
  {32'h464e1750, 32'h00000000} /* (9, 3, 24) {real, imag} */,
  {32'h464346f2, 32'h00000000} /* (9, 3, 23) {real, imag} */,
  {32'h462e14b6, 32'h00000000} /* (9, 3, 22) {real, imag} */,
  {32'h461eaa0b, 32'h00000000} /* (9, 3, 21) {real, imag} */,
  {32'h460e487a, 32'h00000000} /* (9, 3, 20) {real, imag} */,
  {32'h45dd84df, 32'h00000000} /* (9, 3, 19) {real, imag} */,
  {32'h45a34059, 32'h00000000} /* (9, 3, 18) {real, imag} */,
  {32'h4522921a, 32'h00000000} /* (9, 3, 17) {real, imag} */,
  {32'h43562de0, 32'h00000000} /* (9, 3, 16) {real, imag} */,
  {32'hc551bb6c, 32'h00000000} /* (9, 3, 15) {real, imag} */,
  {32'hc5904c2b, 32'h00000000} /* (9, 3, 14) {real, imag} */,
  {32'hc5b8ecb9, 32'h00000000} /* (9, 3, 13) {real, imag} */,
  {32'hc5e3d33f, 32'h00000000} /* (9, 3, 12) {real, imag} */,
  {32'hc5f634f4, 32'h00000000} /* (9, 3, 11) {real, imag} */,
  {32'hc5aa1077, 32'h00000000} /* (9, 3, 10) {real, imag} */,
  {32'hc58736e9, 32'h00000000} /* (9, 3, 9) {real, imag} */,
  {32'hc542d1fe, 32'h00000000} /* (9, 3, 8) {real, imag} */,
  {32'hc4ee7af4, 32'h00000000} /* (9, 3, 7) {real, imag} */,
  {32'h4492a0d4, 32'h00000000} /* (9, 3, 6) {real, imag} */,
  {32'h459bc618, 32'h00000000} /* (9, 3, 5) {real, imag} */,
  {32'h45f61c6b, 32'h00000000} /* (9, 3, 4) {real, imag} */,
  {32'h461d3f76, 32'h00000000} /* (9, 3, 3) {real, imag} */,
  {32'h462bc7a2, 32'h00000000} /* (9, 3, 2) {real, imag} */,
  {32'h464b84dc, 32'h00000000} /* (9, 3, 1) {real, imag} */,
  {32'h4645d1a2, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'h4643e502, 32'h00000000} /* (9, 2, 31) {real, imag} */,
  {32'h46500e06, 32'h00000000} /* (9, 2, 30) {real, imag} */,
  {32'h4652a451, 32'h00000000} /* (9, 2, 29) {real, imag} */,
  {32'h4657ea24, 32'h00000000} /* (9, 2, 28) {real, imag} */,
  {32'h46583a0e, 32'h00000000} /* (9, 2, 27) {real, imag} */,
  {32'h4659e6c1, 32'h00000000} /* (9, 2, 26) {real, imag} */,
  {32'h46656280, 32'h00000000} /* (9, 2, 25) {real, imag} */,
  {32'h46656480, 32'h00000000} /* (9, 2, 24) {real, imag} */,
  {32'h463a91a4, 32'h00000000} /* (9, 2, 23) {real, imag} */,
  {32'h462c7986, 32'h00000000} /* (9, 2, 22) {real, imag} */,
  {32'h46121757, 32'h00000000} /* (9, 2, 21) {real, imag} */,
  {32'h46046e61, 32'h00000000} /* (9, 2, 20) {real, imag} */,
  {32'h45eef07d, 32'h00000000} /* (9, 2, 19) {real, imag} */,
  {32'h45abad4e, 32'h00000000} /* (9, 2, 18) {real, imag} */,
  {32'h4584e478, 32'h00000000} /* (9, 2, 17) {real, imag} */,
  {32'h444e8a88, 32'h00000000} /* (9, 2, 16) {real, imag} */,
  {32'hc5398ec2, 32'h00000000} /* (9, 2, 15) {real, imag} */,
  {32'hc57d01f2, 32'h00000000} /* (9, 2, 14) {real, imag} */,
  {32'hc5b451d6, 32'h00000000} /* (9, 2, 13) {real, imag} */,
  {32'hc5ca2af4, 32'h00000000} /* (9, 2, 12) {real, imag} */,
  {32'hc5c66781, 32'h00000000} /* (9, 2, 11) {real, imag} */,
  {32'hc5ba65c6, 32'h00000000} /* (9, 2, 10) {real, imag} */,
  {32'hc59c5985, 32'h00000000} /* (9, 2, 9) {real, imag} */,
  {32'hc539f20a, 32'h00000000} /* (9, 2, 8) {real, imag} */,
  {32'hc4ccd858, 32'h00000000} /* (9, 2, 7) {real, imag} */,
  {32'h43dbcc90, 32'h00000000} /* (9, 2, 6) {real, imag} */,
  {32'h45a94c76, 32'h00000000} /* (9, 2, 5) {real, imag} */,
  {32'h45fd092a, 32'h00000000} /* (9, 2, 4) {real, imag} */,
  {32'h46132246, 32'h00000000} /* (9, 2, 3) {real, imag} */,
  {32'h4631b033, 32'h00000000} /* (9, 2, 2) {real, imag} */,
  {32'h46377d93, 32'h00000000} /* (9, 2, 1) {real, imag} */,
  {32'h4638999e, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'h46409042, 32'h00000000} /* (9, 1, 31) {real, imag} */,
  {32'h464b82b2, 32'h00000000} /* (9, 1, 30) {real, imag} */,
  {32'h46583012, 32'h00000000} /* (9, 1, 29) {real, imag} */,
  {32'h465d455a, 32'h00000000} /* (9, 1, 28) {real, imag} */,
  {32'h4663c563, 32'h00000000} /* (9, 1, 27) {real, imag} */,
  {32'h4650897e, 32'h00000000} /* (9, 1, 26) {real, imag} */,
  {32'h465de495, 32'h00000000} /* (9, 1, 25) {real, imag} */,
  {32'h4656f428, 32'h00000000} /* (9, 1, 24) {real, imag} */,
  {32'h462e3eee, 32'h00000000} /* (9, 1, 23) {real, imag} */,
  {32'h4621b1c8, 32'h00000000} /* (9, 1, 22) {real, imag} */,
  {32'h4606ee88, 32'h00000000} /* (9, 1, 21) {real, imag} */,
  {32'h45df5b38, 32'h00000000} /* (9, 1, 20) {real, imag} */,
  {32'h45d1d67a, 32'h00000000} /* (9, 1, 19) {real, imag} */,
  {32'h4598ee14, 32'h00000000} /* (9, 1, 18) {real, imag} */,
  {32'h457da27a, 32'h00000000} /* (9, 1, 17) {real, imag} */,
  {32'h43a0e870, 32'h00000000} /* (9, 1, 16) {real, imag} */,
  {32'hc5302df8, 32'h00000000} /* (9, 1, 15) {real, imag} */,
  {32'hc5965ca1, 32'h00000000} /* (9, 1, 14) {real, imag} */,
  {32'hc5d0eb09, 32'h00000000} /* (9, 1, 13) {real, imag} */,
  {32'hc5c87ccc, 32'h00000000} /* (9, 1, 12) {real, imag} */,
  {32'hc5c20c56, 32'h00000000} /* (9, 1, 11) {real, imag} */,
  {32'hc59f4d3c, 32'h00000000} /* (9, 1, 10) {real, imag} */,
  {32'hc583104e, 32'h00000000} /* (9, 1, 9) {real, imag} */,
  {32'hc51be4be, 32'h00000000} /* (9, 1, 8) {real, imag} */,
  {32'hc40a57a8, 32'h00000000} /* (9, 1, 7) {real, imag} */,
  {32'h44de5838, 32'h00000000} /* (9, 1, 6) {real, imag} */,
  {32'h45ad829f, 32'h00000000} /* (9, 1, 5) {real, imag} */,
  {32'h4600e810, 32'h00000000} /* (9, 1, 4) {real, imag} */,
  {32'h4619cf67, 32'h00000000} /* (9, 1, 3) {real, imag} */,
  {32'h462ee4d2, 32'h00000000} /* (9, 1, 2) {real, imag} */,
  {32'h4638c7cc, 32'h00000000} /* (9, 1, 1) {real, imag} */,
  {32'h463b5e78, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'h463fcf9a, 32'h00000000} /* (9, 0, 31) {real, imag} */,
  {32'h46470c62, 32'h00000000} /* (9, 0, 30) {real, imag} */,
  {32'h463e4f9f, 32'h00000000} /* (9, 0, 29) {real, imag} */,
  {32'h465098ed, 32'h00000000} /* (9, 0, 28) {real, imag} */,
  {32'h464ff53d, 32'h00000000} /* (9, 0, 27) {real, imag} */,
  {32'h464a0187, 32'h00000000} /* (9, 0, 26) {real, imag} */,
  {32'h46489606, 32'h00000000} /* (9, 0, 25) {real, imag} */,
  {32'h463f0042, 32'h00000000} /* (9, 0, 24) {real, imag} */,
  {32'h462a92e5, 32'h00000000} /* (9, 0, 23) {real, imag} */,
  {32'h460ccae3, 32'h00000000} /* (9, 0, 22) {real, imag} */,
  {32'h45ed376a, 32'h00000000} /* (9, 0, 21) {real, imag} */,
  {32'h45b0f128, 32'h00000000} /* (9, 0, 20) {real, imag} */,
  {32'h45719829, 32'h00000000} /* (9, 0, 19) {real, imag} */,
  {32'h4530565d, 32'h00000000} /* (9, 0, 18) {real, imag} */,
  {32'h44123968, 32'h00000000} /* (9, 0, 17) {real, imag} */,
  {32'hc48ee420, 32'h00000000} /* (9, 0, 16) {real, imag} */,
  {32'hc557f3c6, 32'h00000000} /* (9, 0, 15) {real, imag} */,
  {32'hc598ab6c, 32'h00000000} /* (9, 0, 14) {real, imag} */,
  {32'hc5c5083e, 32'h00000000} /* (9, 0, 13) {real, imag} */,
  {32'hc5b8c45a, 32'h00000000} /* (9, 0, 12) {real, imag} */,
  {32'hc59fe906, 32'h00000000} /* (9, 0, 11) {real, imag} */,
  {32'hc558fb74, 32'h00000000} /* (9, 0, 10) {real, imag} */,
  {32'hc50fdffe, 32'h00000000} /* (9, 0, 9) {real, imag} */,
  {32'hc4089c78, 32'h00000000} /* (9, 0, 8) {real, imag} */,
  {32'h44a47d20, 32'h00000000} /* (9, 0, 7) {real, imag} */,
  {32'h457dd6b4, 32'h00000000} /* (9, 0, 6) {real, imag} */,
  {32'h45bef22e, 32'h00000000} /* (9, 0, 5) {real, imag} */,
  {32'h4606a30c, 32'h00000000} /* (9, 0, 4) {real, imag} */,
  {32'h461ad8ee, 32'h00000000} /* (9, 0, 3) {real, imag} */,
  {32'h4625cae7, 32'h00000000} /* (9, 0, 2) {real, imag} */,
  {32'h46329c22, 32'h00000000} /* (9, 0, 1) {real, imag} */,
  {32'h46343ae5, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h462c36ad, 32'h00000000} /* (8, 31, 31) {real, imag} */,
  {32'h463166a6, 32'h00000000} /* (8, 31, 30) {real, imag} */,
  {32'h463f6150, 32'h00000000} /* (8, 31, 29) {real, imag} */,
  {32'h463f1b06, 32'h00000000} /* (8, 31, 28) {real, imag} */,
  {32'h463ed4b6, 32'h00000000} /* (8, 31, 27) {real, imag} */,
  {32'h463c9a91, 32'h00000000} /* (8, 31, 26) {real, imag} */,
  {32'h46341c12, 32'h00000000} /* (8, 31, 25) {real, imag} */,
  {32'h46229b78, 32'h00000000} /* (8, 31, 24) {real, imag} */,
  {32'h4612ad54, 32'h00000000} /* (8, 31, 23) {real, imag} */,
  {32'h46021eaa, 32'h00000000} /* (8, 31, 22) {real, imag} */,
  {32'h45b89d7c, 32'h00000000} /* (8, 31, 21) {real, imag} */,
  {32'h454e01e2, 32'h00000000} /* (8, 31, 20) {real, imag} */,
  {32'h44ec6d10, 32'h00000000} /* (8, 31, 19) {real, imag} */,
  {32'h438794d0, 32'h00000000} /* (8, 31, 18) {real, imag} */,
  {32'hc4ca0530, 32'h00000000} /* (8, 31, 17) {real, imag} */,
  {32'hc558aa1b, 32'h00000000} /* (8, 31, 16) {real, imag} */,
  {32'hc5890af0, 32'h00000000} /* (8, 31, 15) {real, imag} */,
  {32'hc59a6f5c, 32'h00000000} /* (8, 31, 14) {real, imag} */,
  {32'hc59f432f, 32'h00000000} /* (8, 31, 13) {real, imag} */,
  {32'hc582844c, 32'h00000000} /* (8, 31, 12) {real, imag} */,
  {32'hc559c510, 32'h00000000} /* (8, 31, 11) {real, imag} */,
  {32'h43dcaea0, 32'h00000000} /* (8, 31, 10) {real, imag} */,
  {32'h44682998, 32'h00000000} /* (8, 31, 9) {real, imag} */,
  {32'h450f1856, 32'h00000000} /* (8, 31, 8) {real, imag} */,
  {32'h458cc0f4, 32'h00000000} /* (8, 31, 7) {real, imag} */,
  {32'h45b7f8a0, 32'h00000000} /* (8, 31, 6) {real, imag} */,
  {32'h45dc72a6, 32'h00000000} /* (8, 31, 5) {real, imag} */,
  {32'h460d2b14, 32'h00000000} /* (8, 31, 4) {real, imag} */,
  {32'h4617c1aa, 32'h00000000} /* (8, 31, 3) {real, imag} */,
  {32'h461ee9b6, 32'h00000000} /* (8, 31, 2) {real, imag} */,
  {32'h46265921, 32'h00000000} /* (8, 31, 1) {real, imag} */,
  {32'h46288e78, 32'h00000000} /* (8, 31, 0) {real, imag} */,
  {32'h4634884d, 32'h00000000} /* (8, 30, 31) {real, imag} */,
  {32'h463c41b4, 32'h00000000} /* (8, 30, 30) {real, imag} */,
  {32'h46399050, 32'h00000000} /* (8, 30, 29) {real, imag} */,
  {32'h464af106, 32'h00000000} /* (8, 30, 28) {real, imag} */,
  {32'h464882bc, 32'h00000000} /* (8, 30, 27) {real, imag} */,
  {32'h46379292, 32'h00000000} /* (8, 30, 26) {real, imag} */,
  {32'h4638b216, 32'h00000000} /* (8, 30, 25) {real, imag} */,
  {32'h4627a533, 32'h00000000} /* (8, 30, 24) {real, imag} */,
  {32'h4609941f, 32'h00000000} /* (8, 30, 23) {real, imag} */,
  {32'h460385ec, 32'h00000000} /* (8, 30, 22) {real, imag} */,
  {32'h45bb0f12, 32'h00000000} /* (8, 30, 21) {real, imag} */,
  {32'h44e55e48, 32'h00000000} /* (8, 30, 20) {real, imag} */,
  {32'hc43c2378, 32'h00000000} /* (8, 30, 19) {real, imag} */,
  {32'hc4f77234, 32'h00000000} /* (8, 30, 18) {real, imag} */,
  {32'hc53eab90, 32'h00000000} /* (8, 30, 17) {real, imag} */,
  {32'hc5a600e7, 32'h00000000} /* (8, 30, 16) {real, imag} */,
  {32'hc5ae8726, 32'h00000000} /* (8, 30, 15) {real, imag} */,
  {32'hc5ad74e0, 32'h00000000} /* (8, 30, 14) {real, imag} */,
  {32'hc5a70080, 32'h00000000} /* (8, 30, 13) {real, imag} */,
  {32'hc5874a74, 32'h00000000} /* (8, 30, 12) {real, imag} */,
  {32'hc52a6d36, 32'h00000000} /* (8, 30, 11) {real, imag} */,
  {32'h449f48b0, 32'h00000000} /* (8, 30, 10) {real, imag} */,
  {32'h4512aee8, 32'h00000000} /* (8, 30, 9) {real, imag} */,
  {32'h458762f6, 32'h00000000} /* (8, 30, 8) {real, imag} */,
  {32'h45c085c6, 32'h00000000} /* (8, 30, 7) {real, imag} */,
  {32'h45df0758, 32'h00000000} /* (8, 30, 6) {real, imag} */,
  {32'h461a6071, 32'h00000000} /* (8, 30, 5) {real, imag} */,
  {32'h461ff33d, 32'h00000000} /* (8, 30, 4) {real, imag} */,
  {32'h46213d1c, 32'h00000000} /* (8, 30, 3) {real, imag} */,
  {32'h463029a6, 32'h00000000} /* (8, 30, 2) {real, imag} */,
  {32'h4640ea1a, 32'h00000000} /* (8, 30, 1) {real, imag} */,
  {32'h462aff30, 32'h00000000} /* (8, 30, 0) {real, imag} */,
  {32'h463fa60c, 32'h00000000} /* (8, 29, 31) {real, imag} */,
  {32'h4646b05e, 32'h00000000} /* (8, 29, 30) {real, imag} */,
  {32'h46370870, 32'h00000000} /* (8, 29, 29) {real, imag} */,
  {32'h463926f1, 32'h00000000} /* (8, 29, 28) {real, imag} */,
  {32'h463745b9, 32'h00000000} /* (8, 29, 27) {real, imag} */,
  {32'h463129e6, 32'h00000000} /* (8, 29, 26) {real, imag} */,
  {32'h4628aefb, 32'h00000000} /* (8, 29, 25) {real, imag} */,
  {32'h461bd695, 32'h00000000} /* (8, 29, 24) {real, imag} */,
  {32'h4609504d, 32'h00000000} /* (8, 29, 23) {real, imag} */,
  {32'h45ee6b2c, 32'h00000000} /* (8, 29, 22) {real, imag} */,
  {32'h45953f30, 32'h00000000} /* (8, 29, 21) {real, imag} */,
  {32'hc2abc9c0, 32'h00000000} /* (8, 29, 20) {real, imag} */,
  {32'hc4d1b6f0, 32'h00000000} /* (8, 29, 19) {real, imag} */,
  {32'hc56f0426, 32'h00000000} /* (8, 29, 18) {real, imag} */,
  {32'hc591a7fa, 32'h00000000} /* (8, 29, 17) {real, imag} */,
  {32'hc5ad0bea, 32'h00000000} /* (8, 29, 16) {real, imag} */,
  {32'hc5c7afbf, 32'h00000000} /* (8, 29, 15) {real, imag} */,
  {32'hc5bf8e73, 32'h00000000} /* (8, 29, 14) {real, imag} */,
  {32'hc5b62650, 32'h00000000} /* (8, 29, 13) {real, imag} */,
  {32'hc58701d2, 32'h00000000} /* (8, 29, 12) {real, imag} */,
  {32'hc5295bdc, 32'h00000000} /* (8, 29, 11) {real, imag} */,
  {32'h449856e0, 32'h00000000} /* (8, 29, 10) {real, imag} */,
  {32'h455a2034, 32'h00000000} /* (8, 29, 9) {real, imag} */,
  {32'h45ace47a, 32'h00000000} /* (8, 29, 8) {real, imag} */,
  {32'h45d89903, 32'h00000000} /* (8, 29, 7) {real, imag} */,
  {32'h45f6ffba, 32'h00000000} /* (8, 29, 6) {real, imag} */,
  {32'h461a80d2, 32'h00000000} /* (8, 29, 5) {real, imag} */,
  {32'h4627f0fa, 32'h00000000} /* (8, 29, 4) {real, imag} */,
  {32'h46326da0, 32'h00000000} /* (8, 29, 3) {real, imag} */,
  {32'h463fdb30, 32'h00000000} /* (8, 29, 2) {real, imag} */,
  {32'h46465f93, 32'h00000000} /* (8, 29, 1) {real, imag} */,
  {32'h463134b5, 32'h00000000} /* (8, 29, 0) {real, imag} */,
  {32'h46323b55, 32'h00000000} /* (8, 28, 31) {real, imag} */,
  {32'h4643b872, 32'h00000000} /* (8, 28, 30) {real, imag} */,
  {32'h46372a34, 32'h00000000} /* (8, 28, 29) {real, imag} */,
  {32'h462cdf11, 32'h00000000} /* (8, 28, 28) {real, imag} */,
  {32'h462e1775, 32'h00000000} /* (8, 28, 27) {real, imag} */,
  {32'h463550e4, 32'h00000000} /* (8, 28, 26) {real, imag} */,
  {32'h462ecb9a, 32'h00000000} /* (8, 28, 25) {real, imag} */,
  {32'h46175238, 32'h00000000} /* (8, 28, 24) {real, imag} */,
  {32'h4609d3fa, 32'h00000000} /* (8, 28, 23) {real, imag} */,
  {32'h45ce35b1, 32'h00000000} /* (8, 28, 22) {real, imag} */,
  {32'h457d3a4d, 32'h00000000} /* (8, 28, 21) {real, imag} */,
  {32'h43096180, 32'h00000000} /* (8, 28, 20) {real, imag} */,
  {32'hc50706fa, 32'h00000000} /* (8, 28, 19) {real, imag} */,
  {32'hc5816d8b, 32'h00000000} /* (8, 28, 18) {real, imag} */,
  {32'hc5909fb5, 32'h00000000} /* (8, 28, 17) {real, imag} */,
  {32'hc5c6ce65, 32'h00000000} /* (8, 28, 16) {real, imag} */,
  {32'hc5cc99a2, 32'h00000000} /* (8, 28, 15) {real, imag} */,
  {32'hc5ea10b4, 32'h00000000} /* (8, 28, 14) {real, imag} */,
  {32'hc5ca4dcd, 32'h00000000} /* (8, 28, 13) {real, imag} */,
  {32'hc5814782, 32'h00000000} /* (8, 28, 12) {real, imag} */,
  {32'hc52cfa70, 32'h00000000} /* (8, 28, 11) {real, imag} */,
  {32'h44956f88, 32'h00000000} /* (8, 28, 10) {real, imag} */,
  {32'h45815fdd, 32'h00000000} /* (8, 28, 9) {real, imag} */,
  {32'h45db4bb8, 32'h00000000} /* (8, 28, 8) {real, imag} */,
  {32'h45e29f97, 32'h00000000} /* (8, 28, 7) {real, imag} */,
  {32'h460cd542, 32'h00000000} /* (8, 28, 6) {real, imag} */,
  {32'h461cae10, 32'h00000000} /* (8, 28, 5) {real, imag} */,
  {32'h4634a30a, 32'h00000000} /* (8, 28, 4) {real, imag} */,
  {32'h46327b10, 32'h00000000} /* (8, 28, 3) {real, imag} */,
  {32'h4642d036, 32'h00000000} /* (8, 28, 2) {real, imag} */,
  {32'h462f9d96, 32'h00000000} /* (8, 28, 1) {real, imag} */,
  {32'h462e07fe, 32'h00000000} /* (8, 28, 0) {real, imag} */,
  {32'h4633e354, 32'h00000000} /* (8, 27, 31) {real, imag} */,
  {32'h463a7b98, 32'h00000000} /* (8, 27, 30) {real, imag} */,
  {32'h462f825d, 32'h00000000} /* (8, 27, 29) {real, imag} */,
  {32'h463a4610, 32'h00000000} /* (8, 27, 28) {real, imag} */,
  {32'h462ac47c, 32'h00000000} /* (8, 27, 27) {real, imag} */,
  {32'h4637ff52, 32'h00000000} /* (8, 27, 26) {real, imag} */,
  {32'h46277900, 32'h00000000} /* (8, 27, 25) {real, imag} */,
  {32'h461a2ac7, 32'h00000000} /* (8, 27, 24) {real, imag} */,
  {32'h46156c96, 32'h00000000} /* (8, 27, 23) {real, imag} */,
  {32'h45afa7a4, 32'h00000000} /* (8, 27, 22) {real, imag} */,
  {32'h456f1dca, 32'h00000000} /* (8, 27, 21) {real, imag} */,
  {32'h43c9c450, 32'h00000000} /* (8, 27, 20) {real, imag} */,
  {32'hc53ee288, 32'h00000000} /* (8, 27, 19) {real, imag} */,
  {32'hc58cc883, 32'h00000000} /* (8, 27, 18) {real, imag} */,
  {32'hc5d3181f, 32'h00000000} /* (8, 27, 17) {real, imag} */,
  {32'hc5de2a0c, 32'h00000000} /* (8, 27, 16) {real, imag} */,
  {32'hc5e75d73, 32'h00000000} /* (8, 27, 15) {real, imag} */,
  {32'hc5e1b63c, 32'h00000000} /* (8, 27, 14) {real, imag} */,
  {32'hc5b22d96, 32'h00000000} /* (8, 27, 13) {real, imag} */,
  {32'hc582800c, 32'h00000000} /* (8, 27, 12) {real, imag} */,
  {32'hc4beede4, 32'h00000000} /* (8, 27, 11) {real, imag} */,
  {32'h44ef372c, 32'h00000000} /* (8, 27, 10) {real, imag} */,
  {32'h45a96c62, 32'h00000000} /* (8, 27, 9) {real, imag} */,
  {32'h45e52891, 32'h00000000} /* (8, 27, 8) {real, imag} */,
  {32'h4609c842, 32'h00000000} /* (8, 27, 7) {real, imag} */,
  {32'h460ab8da, 32'h00000000} /* (8, 27, 6) {real, imag} */,
  {32'h4622dfa6, 32'h00000000} /* (8, 27, 5) {real, imag} */,
  {32'h464637fa, 32'h00000000} /* (8, 27, 4) {real, imag} */,
  {32'h46300022, 32'h00000000} /* (8, 27, 3) {real, imag} */,
  {32'h462cc824, 32'h00000000} /* (8, 27, 2) {real, imag} */,
  {32'h463516c8, 32'h00000000} /* (8, 27, 1) {real, imag} */,
  {32'h4635a188, 32'h00000000} /* (8, 27, 0) {real, imag} */,
  {32'h462f9412, 32'h00000000} /* (8, 26, 31) {real, imag} */,
  {32'h462880e5, 32'h00000000} /* (8, 26, 30) {real, imag} */,
  {32'h462e051a, 32'h00000000} /* (8, 26, 29) {real, imag} */,
  {32'h463565e9, 32'h00000000} /* (8, 26, 28) {real, imag} */,
  {32'h4626e89b, 32'h00000000} /* (8, 26, 27) {real, imag} */,
  {32'h4631378c, 32'h00000000} /* (8, 26, 26) {real, imag} */,
  {32'h462a8932, 32'h00000000} /* (8, 26, 25) {real, imag} */,
  {32'h460dcb62, 32'h00000000} /* (8, 26, 24) {real, imag} */,
  {32'h45fcb52e, 32'h00000000} /* (8, 26, 23) {real, imag} */,
  {32'h45af1c8c, 32'h00000000} /* (8, 26, 22) {real, imag} */,
  {32'h45131e2e, 32'h00000000} /* (8, 26, 21) {real, imag} */,
  {32'hc467e4d0, 32'h00000000} /* (8, 26, 20) {real, imag} */,
  {32'hc553944a, 32'h00000000} /* (8, 26, 19) {real, imag} */,
  {32'hc59e75bf, 32'h00000000} /* (8, 26, 18) {real, imag} */,
  {32'hc5c31f9c, 32'h00000000} /* (8, 26, 17) {real, imag} */,
  {32'hc5d456e6, 32'h00000000} /* (8, 26, 16) {real, imag} */,
  {32'hc5df84bf, 32'h00000000} /* (8, 26, 15) {real, imag} */,
  {32'hc5e1bac2, 32'h00000000} /* (8, 26, 14) {real, imag} */,
  {32'hc5b86243, 32'h00000000} /* (8, 26, 13) {real, imag} */,
  {32'hc5496398, 32'h00000000} /* (8, 26, 12) {real, imag} */,
  {32'hc4da3340, 32'h00000000} /* (8, 26, 11) {real, imag} */,
  {32'h45146fa6, 32'h00000000} /* (8, 26, 10) {real, imag} */,
  {32'h45b1f2f3, 32'h00000000} /* (8, 26, 9) {real, imag} */,
  {32'h45f3fd3d, 32'h00000000} /* (8, 26, 8) {real, imag} */,
  {32'h460e171d, 32'h00000000} /* (8, 26, 7) {real, imag} */,
  {32'h460bc9d4, 32'h00000000} /* (8, 26, 6) {real, imag} */,
  {32'h4619e526, 32'h00000000} /* (8, 26, 5) {real, imag} */,
  {32'h4637f85c, 32'h00000000} /* (8, 26, 4) {real, imag} */,
  {32'h4625fffe, 32'h00000000} /* (8, 26, 3) {real, imag} */,
  {32'h462b7018, 32'h00000000} /* (8, 26, 2) {real, imag} */,
  {32'h462cf540, 32'h00000000} /* (8, 26, 1) {real, imag} */,
  {32'h46231115, 32'h00000000} /* (8, 26, 0) {real, imag} */,
  {32'h4617938d, 32'h00000000} /* (8, 25, 31) {real, imag} */,
  {32'h4624af82, 32'h00000000} /* (8, 25, 30) {real, imag} */,
  {32'h4622c0ba, 32'h00000000} /* (8, 25, 29) {real, imag} */,
  {32'h462785a5, 32'h00000000} /* (8, 25, 28) {real, imag} */,
  {32'h4622be8c, 32'h00000000} /* (8, 25, 27) {real, imag} */,
  {32'h4618f580, 32'h00000000} /* (8, 25, 26) {real, imag} */,
  {32'h4618438a, 32'h00000000} /* (8, 25, 25) {real, imag} */,
  {32'h4603be64, 32'h00000000} /* (8, 25, 24) {real, imag} */,
  {32'h45d7c22a, 32'h00000000} /* (8, 25, 23) {real, imag} */,
  {32'h459d7534, 32'h00000000} /* (8, 25, 22) {real, imag} */,
  {32'h450751f4, 32'h00000000} /* (8, 25, 21) {real, imag} */,
  {32'hc4a5e42c, 32'h00000000} /* (8, 25, 20) {real, imag} */,
  {32'hc56d2914, 32'h00000000} /* (8, 25, 19) {real, imag} */,
  {32'hc5955123, 32'h00000000} /* (8, 25, 18) {real, imag} */,
  {32'hc5a4fbb8, 32'h00000000} /* (8, 25, 17) {real, imag} */,
  {32'hc5b6897f, 32'h00000000} /* (8, 25, 16) {real, imag} */,
  {32'hc5ccdaf0, 32'h00000000} /* (8, 25, 15) {real, imag} */,
  {32'hc5d84da0, 32'h00000000} /* (8, 25, 14) {real, imag} */,
  {32'hc5b12ca2, 32'h00000000} /* (8, 25, 13) {real, imag} */,
  {32'hc53b662f, 32'h00000000} /* (8, 25, 12) {real, imag} */,
  {32'hc4883404, 32'h00000000} /* (8, 25, 11) {real, imag} */,
  {32'h450ac770, 32'h00000000} /* (8, 25, 10) {real, imag} */,
  {32'h45a54e9b, 32'h00000000} /* (8, 25, 9) {real, imag} */,
  {32'h45d82329, 32'h00000000} /* (8, 25, 8) {real, imag} */,
  {32'h4607ec83, 32'h00000000} /* (8, 25, 7) {real, imag} */,
  {32'h460123be, 32'h00000000} /* (8, 25, 6) {real, imag} */,
  {32'h461868b9, 32'h00000000} /* (8, 25, 5) {real, imag} */,
  {32'h46263c5e, 32'h00000000} /* (8, 25, 4) {real, imag} */,
  {32'h461994fd, 32'h00000000} /* (8, 25, 3) {real, imag} */,
  {32'h461817ec, 32'h00000000} /* (8, 25, 2) {real, imag} */,
  {32'h461c43e4, 32'h00000000} /* (8, 25, 1) {real, imag} */,
  {32'h46193156, 32'h00000000} /* (8, 25, 0) {real, imag} */,
  {32'h460656be, 32'h00000000} /* (8, 24, 31) {real, imag} */,
  {32'h460f910e, 32'h00000000} /* (8, 24, 30) {real, imag} */,
  {32'h46093eb6, 32'h00000000} /* (8, 24, 29) {real, imag} */,
  {32'h4625f59a, 32'h00000000} /* (8, 24, 28) {real, imag} */,
  {32'h461b4b6d, 32'h00000000} /* (8, 24, 27) {real, imag} */,
  {32'h4617d785, 32'h00000000} /* (8, 24, 26) {real, imag} */,
  {32'h46091b28, 32'h00000000} /* (8, 24, 25) {real, imag} */,
  {32'h45e67fb1, 32'h00000000} /* (8, 24, 24) {real, imag} */,
  {32'h45b311d6, 32'h00000000} /* (8, 24, 23) {real, imag} */,
  {32'h459786a0, 32'h00000000} /* (8, 24, 22) {real, imag} */,
  {32'h4508930d, 32'h00000000} /* (8, 24, 21) {real, imag} */,
  {32'hc434b4c0, 32'h00000000} /* (8, 24, 20) {real, imag} */,
  {32'hc5840d4e, 32'h00000000} /* (8, 24, 19) {real, imag} */,
  {32'hc58b4de3, 32'h00000000} /* (8, 24, 18) {real, imag} */,
  {32'hc5965a16, 32'h00000000} /* (8, 24, 17) {real, imag} */,
  {32'hc598ea56, 32'h00000000} /* (8, 24, 16) {real, imag} */,
  {32'hc5cd3d0c, 32'h00000000} /* (8, 24, 15) {real, imag} */,
  {32'hc5b1b341, 32'h00000000} /* (8, 24, 14) {real, imag} */,
  {32'hc599181d, 32'h00000000} /* (8, 24, 13) {real, imag} */,
  {32'hc54d00ae, 32'h00000000} /* (8, 24, 12) {real, imag} */,
  {32'hc3f121a0, 32'h00000000} /* (8, 24, 11) {real, imag} */,
  {32'h453c14b5, 32'h00000000} /* (8, 24, 10) {real, imag} */,
  {32'h45a227f9, 32'h00000000} /* (8, 24, 9) {real, imag} */,
  {32'h45c4d455, 32'h00000000} /* (8, 24, 8) {real, imag} */,
  {32'h45ef2eda, 32'h00000000} /* (8, 24, 7) {real, imag} */,
  {32'h46082253, 32'h00000000} /* (8, 24, 6) {real, imag} */,
  {32'h46034ab3, 32'h00000000} /* (8, 24, 5) {real, imag} */,
  {32'h4611bd3d, 32'h00000000} /* (8, 24, 4) {real, imag} */,
  {32'h460f9dde, 32'h00000000} /* (8, 24, 3) {real, imag} */,
  {32'h4607ac54, 32'h00000000} /* (8, 24, 2) {real, imag} */,
  {32'h46147b03, 32'h00000000} /* (8, 24, 1) {real, imag} */,
  {32'h45fdac8c, 32'h00000000} /* (8, 24, 0) {real, imag} */,
  {32'h45d12abe, 32'h00000000} /* (8, 23, 31) {real, imag} */,
  {32'h460279d8, 32'h00000000} /* (8, 23, 30) {real, imag} */,
  {32'h45f54489, 32'h00000000} /* (8, 23, 29) {real, imag} */,
  {32'h46067442, 32'h00000000} /* (8, 23, 28) {real, imag} */,
  {32'h45f6aa08, 32'h00000000} /* (8, 23, 27) {real, imag} */,
  {32'h45e5a7ff, 32'h00000000} /* (8, 23, 26) {real, imag} */,
  {32'h45d0f3bb, 32'h00000000} /* (8, 23, 25) {real, imag} */,
  {32'h45b8850d, 32'h00000000} /* (8, 23, 24) {real, imag} */,
  {32'h45a218a4, 32'h00000000} /* (8, 23, 23) {real, imag} */,
  {32'h4571d05c, 32'h00000000} /* (8, 23, 22) {real, imag} */,
  {32'h4501dff6, 32'h00000000} /* (8, 23, 21) {real, imag} */,
  {32'hc48bd114, 32'h00000000} /* (8, 23, 20) {real, imag} */,
  {32'hc53afb58, 32'h00000000} /* (8, 23, 19) {real, imag} */,
  {32'hc5451f3b, 32'h00000000} /* (8, 23, 18) {real, imag} */,
  {32'hc5532d89, 32'h00000000} /* (8, 23, 17) {real, imag} */,
  {32'hc58228c8, 32'h00000000} /* (8, 23, 16) {real, imag} */,
  {32'hc5886a62, 32'h00000000} /* (8, 23, 15) {real, imag} */,
  {32'hc58ef5d2, 32'h00000000} /* (8, 23, 14) {real, imag} */,
  {32'hc595fa0b, 32'h00000000} /* (8, 23, 13) {real, imag} */,
  {32'hc5520146, 32'h00000000} /* (8, 23, 12) {real, imag} */,
  {32'hc4420b20, 32'h00000000} /* (8, 23, 11) {real, imag} */,
  {32'h44daf364, 32'h00000000} /* (8, 23, 10) {real, imag} */,
  {32'h45a4eb0d, 32'h00000000} /* (8, 23, 9) {real, imag} */,
  {32'h45a26f73, 32'h00000000} /* (8, 23, 8) {real, imag} */,
  {32'h45e5bf1c, 32'h00000000} /* (8, 23, 7) {real, imag} */,
  {32'h45d19668, 32'h00000000} /* (8, 23, 6) {real, imag} */,
  {32'h45e73ffb, 32'h00000000} /* (8, 23, 5) {real, imag} */,
  {32'h45eb0ef9, 32'h00000000} /* (8, 23, 4) {real, imag} */,
  {32'h45ee3684, 32'h00000000} /* (8, 23, 3) {real, imag} */,
  {32'h45ec61e4, 32'h00000000} /* (8, 23, 2) {real, imag} */,
  {32'h45c6f99a, 32'h00000000} /* (8, 23, 1) {real, imag} */,
  {32'h45bca778, 32'h00000000} /* (8, 23, 0) {real, imag} */,
  {32'h4583e7ac, 32'h00000000} /* (8, 22, 31) {real, imag} */,
  {32'h459e300f, 32'h00000000} /* (8, 22, 30) {real, imag} */,
  {32'h45cd1c59, 32'h00000000} /* (8, 22, 29) {real, imag} */,
  {32'h459323fe, 32'h00000000} /* (8, 22, 28) {real, imag} */,
  {32'h45a5feb8, 32'h00000000} /* (8, 22, 27) {real, imag} */,
  {32'h45a8b6f7, 32'h00000000} /* (8, 22, 26) {real, imag} */,
  {32'h458f002e, 32'h00000000} /* (8, 22, 25) {real, imag} */,
  {32'h4594a9a6, 32'h00000000} /* (8, 22, 24) {real, imag} */,
  {32'h458ae6c7, 32'h00000000} /* (8, 22, 23) {real, imag} */,
  {32'h4544c642, 32'h00000000} /* (8, 22, 22) {real, imag} */,
  {32'h45055b00, 32'h00000000} /* (8, 22, 21) {real, imag} */,
  {32'hc2c7fd00, 32'h00000000} /* (8, 22, 20) {real, imag} */,
  {32'hc4e97fb2, 32'h00000000} /* (8, 22, 19) {real, imag} */,
  {32'hc50a29e4, 32'h00000000} /* (8, 22, 18) {real, imag} */,
  {32'hc51d13d6, 32'h00000000} /* (8, 22, 17) {real, imag} */,
  {32'hc5126f2a, 32'h00000000} /* (8, 22, 16) {real, imag} */,
  {32'hc512a663, 32'h00000000} /* (8, 22, 15) {real, imag} */,
  {32'hc54cdfa2, 32'h00000000} /* (8, 22, 14) {real, imag} */,
  {32'hc51cda9e, 32'h00000000} /* (8, 22, 13) {real, imag} */,
  {32'hc4d80426, 32'h00000000} /* (8, 22, 12) {real, imag} */,
  {32'hc434930c, 32'h00000000} /* (8, 22, 11) {real, imag} */,
  {32'h45260296, 32'h00000000} /* (8, 22, 10) {real, imag} */,
  {32'h45400b74, 32'h00000000} /* (8, 22, 9) {real, imag} */,
  {32'h45552184, 32'h00000000} /* (8, 22, 8) {real, imag} */,
  {32'h459bd741, 32'h00000000} /* (8, 22, 7) {real, imag} */,
  {32'h458c6927, 32'h00000000} /* (8, 22, 6) {real, imag} */,
  {32'h459e6d50, 32'h00000000} /* (8, 22, 5) {real, imag} */,
  {32'h458cf3e5, 32'h00000000} /* (8, 22, 4) {real, imag} */,
  {32'h45ab020e, 32'h00000000} /* (8, 22, 3) {real, imag} */,
  {32'h459792f6, 32'h00000000} /* (8, 22, 2) {real, imag} */,
  {32'h458942e6, 32'h00000000} /* (8, 22, 1) {real, imag} */,
  {32'h45790b0a, 32'h00000000} /* (8, 22, 0) {real, imag} */,
  {32'h44d6c092, 32'h00000000} /* (8, 21, 31) {real, imag} */,
  {32'h450941ce, 32'h00000000} /* (8, 21, 30) {real, imag} */,
  {32'h45077653, 32'h00000000} /* (8, 21, 29) {real, imag} */,
  {32'h45044758, 32'h00000000} /* (8, 21, 28) {real, imag} */,
  {32'h45054126, 32'h00000000} /* (8, 21, 27) {real, imag} */,
  {32'h44d57f1c, 32'h00000000} /* (8, 21, 26) {real, imag} */,
  {32'h44f224dd, 32'h00000000} /* (8, 21, 25) {real, imag} */,
  {32'h44b62f27, 32'h00000000} /* (8, 21, 24) {real, imag} */,
  {32'h449e8e73, 32'h00000000} /* (8, 21, 23) {real, imag} */,
  {32'h447b775c, 32'h00000000} /* (8, 21, 22) {real, imag} */,
  {32'h448dc0fc, 32'h00000000} /* (8, 21, 21) {real, imag} */,
  {32'h43f771ae, 32'h00000000} /* (8, 21, 20) {real, imag} */,
  {32'hc493021e, 32'h00000000} /* (8, 21, 19) {real, imag} */,
  {32'hc402d326, 32'h00000000} /* (8, 21, 18) {real, imag} */,
  {32'hc3dc1172, 32'h00000000} /* (8, 21, 17) {real, imag} */,
  {32'hc40f7a4a, 32'h00000000} /* (8, 21, 16) {real, imag} */,
  {32'h43197d74, 32'h00000000} /* (8, 21, 15) {real, imag} */,
  {32'hc466cc28, 32'h00000000} /* (8, 21, 14) {real, imag} */,
  {32'h41f9ac80, 32'h00000000} /* (8, 21, 13) {real, imag} */,
  {32'h441a48e6, 32'h00000000} /* (8, 21, 12) {real, imag} */,
  {32'h436b2414, 32'h00000000} /* (8, 21, 11) {real, imag} */,
  {32'h44c063f2, 32'h00000000} /* (8, 21, 10) {real, imag} */,
  {32'h44ab570f, 32'h00000000} /* (8, 21, 9) {real, imag} */,
  {32'h449e0db9, 32'h00000000} /* (8, 21, 8) {real, imag} */,
  {32'h449ad971, 32'h00000000} /* (8, 21, 7) {real, imag} */,
  {32'h44b5daba, 32'h00000000} /* (8, 21, 6) {real, imag} */,
  {32'h44b5bd60, 32'h00000000} /* (8, 21, 5) {real, imag} */,
  {32'h4487f554, 32'h00000000} /* (8, 21, 4) {real, imag} */,
  {32'h4510b425, 32'h00000000} /* (8, 21, 3) {real, imag} */,
  {32'h449aa079, 32'h00000000} /* (8, 21, 2) {real, imag} */,
  {32'h44c1f24c, 32'h00000000} /* (8, 21, 1) {real, imag} */,
  {32'h4452d028, 32'h00000000} /* (8, 21, 0) {real, imag} */,
  {32'hc4ba04f1, 32'h00000000} /* (8, 20, 31) {real, imag} */,
  {32'hc530b061, 32'h00000000} /* (8, 20, 30) {real, imag} */,
  {32'hc4c7d171, 32'h00000000} /* (8, 20, 29) {real, imag} */,
  {32'hc491519b, 32'h00000000} /* (8, 20, 28) {real, imag} */,
  {32'hc50ce315, 32'h00000000} /* (8, 20, 27) {real, imag} */,
  {32'hc4f299d4, 32'h00000000} /* (8, 20, 26) {real, imag} */,
  {32'hc4b211fe, 32'h00000000} /* (8, 20, 25) {real, imag} */,
  {32'hc4cc59c2, 32'h00000000} /* (8, 20, 24) {real, imag} */,
  {32'hc4d8f36f, 32'h00000000} /* (8, 20, 23) {real, imag} */,
  {32'hc47707f8, 32'h00000000} /* (8, 20, 22) {real, imag} */,
  {32'hc28c68d0, 32'h00000000} /* (8, 20, 21) {real, imag} */,
  {32'h4453503e, 32'h00000000} /* (8, 20, 20) {real, imag} */,
  {32'h44cdc44a, 32'h00000000} /* (8, 20, 19) {real, imag} */,
  {32'h450cf7ba, 32'h00000000} /* (8, 20, 18) {real, imag} */,
  {32'h454c0cb6, 32'h00000000} /* (8, 20, 17) {real, imag} */,
  {32'h4534be13, 32'h00000000} /* (8, 20, 16) {real, imag} */,
  {32'h453a48ba, 32'h00000000} /* (8, 20, 15) {real, imag} */,
  {32'h45222847, 32'h00000000} /* (8, 20, 14) {real, imag} */,
  {32'h4545c930, 32'h00000000} /* (8, 20, 13) {real, imag} */,
  {32'h451cc5a0, 32'h00000000} /* (8, 20, 12) {real, imag} */,
  {32'h44b98f2a, 32'h00000000} /* (8, 20, 11) {real, imag} */,
  {32'hc3373224, 32'h00000000} /* (8, 20, 10) {real, imag} */,
  {32'hc458d33c, 32'h00000000} /* (8, 20, 9) {real, imag} */,
  {32'hc50710e1, 32'h00000000} /* (8, 20, 8) {real, imag} */,
  {32'hc5261c0c, 32'h00000000} /* (8, 20, 7) {real, imag} */,
  {32'hc502d30a, 32'h00000000} /* (8, 20, 6) {real, imag} */,
  {32'hc531fe9a, 32'h00000000} /* (8, 20, 5) {real, imag} */,
  {32'hc551c91a, 32'h00000000} /* (8, 20, 4) {real, imag} */,
  {32'hc4fe93e2, 32'h00000000} /* (8, 20, 3) {real, imag} */,
  {32'hc5203986, 32'h00000000} /* (8, 20, 2) {real, imag} */,
  {32'hc5217af8, 32'h00000000} /* (8, 20, 1) {real, imag} */,
  {32'hc4d9562e, 32'h00000000} /* (8, 20, 0) {real, imag} */,
  {32'hc57d6dc0, 32'h00000000} /* (8, 19, 31) {real, imag} */,
  {32'hc57fb628, 32'h00000000} /* (8, 19, 30) {real, imag} */,
  {32'hc58e6e4c, 32'h00000000} /* (8, 19, 29) {real, imag} */,
  {32'hc5977ab6, 32'h00000000} /* (8, 19, 28) {real, imag} */,
  {32'hc57b88ab, 32'h00000000} /* (8, 19, 27) {real, imag} */,
  {32'hc5952929, 32'h00000000} /* (8, 19, 26) {real, imag} */,
  {32'hc58e3346, 32'h00000000} /* (8, 19, 25) {real, imag} */,
  {32'hc55d20d5, 32'h00000000} /* (8, 19, 24) {real, imag} */,
  {32'hc53ac08e, 32'h00000000} /* (8, 19, 23) {real, imag} */,
  {32'hc4dd51cd, 32'h00000000} /* (8, 19, 22) {real, imag} */,
  {32'hc4116c42, 32'h00000000} /* (8, 19, 21) {real, imag} */,
  {32'h4539a4d5, 32'h00000000} /* (8, 19, 20) {real, imag} */,
  {32'h45768832, 32'h00000000} /* (8, 19, 19) {real, imag} */,
  {32'h45596b3c, 32'h00000000} /* (8, 19, 18) {real, imag} */,
  {32'h4597998c, 32'h00000000} /* (8, 19, 17) {real, imag} */,
  {32'h45995cb8, 32'h00000000} /* (8, 19, 16) {real, imag} */,
  {32'h45a72dd6, 32'h00000000} /* (8, 19, 15) {real, imag} */,
  {32'h45a1ae24, 32'h00000000} /* (8, 19, 14) {real, imag} */,
  {32'h45b1447c, 32'h00000000} /* (8, 19, 13) {real, imag} */,
  {32'h452d0d72, 32'h00000000} /* (8, 19, 12) {real, imag} */,
  {32'h44bbc6b6, 32'h00000000} /* (8, 19, 11) {real, imag} */,
  {32'h42e73040, 32'h00000000} /* (8, 19, 10) {real, imag} */,
  {32'hc580ad3a, 32'h00000000} /* (8, 19, 9) {real, imag} */,
  {32'hc58eea72, 32'h00000000} /* (8, 19, 8) {real, imag} */,
  {32'hc58cb8f1, 32'h00000000} /* (8, 19, 7) {real, imag} */,
  {32'hc587f00f, 32'h00000000} /* (8, 19, 6) {real, imag} */,
  {32'hc589c67d, 32'h00000000} /* (8, 19, 5) {real, imag} */,
  {32'hc59fcfea, 32'h00000000} /* (8, 19, 4) {real, imag} */,
  {32'hc5c4fd15, 32'h00000000} /* (8, 19, 3) {real, imag} */,
  {32'hc5b4cf4e, 32'h00000000} /* (8, 19, 2) {real, imag} */,
  {32'hc5907cf0, 32'h00000000} /* (8, 19, 1) {real, imag} */,
  {32'hc583b73a, 32'h00000000} /* (8, 19, 0) {real, imag} */,
  {32'hc5d501d0, 32'h00000000} /* (8, 18, 31) {real, imag} */,
  {32'hc5e3923a, 32'h00000000} /* (8, 18, 30) {real, imag} */,
  {32'hc5c5e3cd, 32'h00000000} /* (8, 18, 29) {real, imag} */,
  {32'hc5ba7238, 32'h00000000} /* (8, 18, 28) {real, imag} */,
  {32'hc5c3e1ac, 32'h00000000} /* (8, 18, 27) {real, imag} */,
  {32'hc5c9c712, 32'h00000000} /* (8, 18, 26) {real, imag} */,
  {32'hc5bfc501, 32'h00000000} /* (8, 18, 25) {real, imag} */,
  {32'hc5bd9420, 32'h00000000} /* (8, 18, 24) {real, imag} */,
  {32'hc5b24c52, 32'h00000000} /* (8, 18, 23) {real, imag} */,
  {32'hc55258f2, 32'h00000000} /* (8, 18, 22) {real, imag} */,
  {32'hc180ad80, 32'h00000000} /* (8, 18, 21) {real, imag} */,
  {32'h455523a3, 32'h00000000} /* (8, 18, 20) {real, imag} */,
  {32'h4592b041, 32'h00000000} /* (8, 18, 19) {real, imag} */,
  {32'h459a3f9f, 32'h00000000} /* (8, 18, 18) {real, imag} */,
  {32'h45b2d35f, 32'h00000000} /* (8, 18, 17) {real, imag} */,
  {32'h45d066e0, 32'h00000000} /* (8, 18, 16) {real, imag} */,
  {32'h45db341c, 32'h00000000} /* (8, 18, 15) {real, imag} */,
  {32'h45d8ca9a, 32'h00000000} /* (8, 18, 14) {real, imag} */,
  {32'h45a57f93, 32'h00000000} /* (8, 18, 13) {real, imag} */,
  {32'h458cbbd0, 32'h00000000} /* (8, 18, 12) {real, imag} */,
  {32'h44c40c32, 32'h00000000} /* (8, 18, 11) {real, imag} */,
  {32'hc4fb53d0, 32'h00000000} /* (8, 18, 10) {real, imag} */,
  {32'hc51fb9ea, 32'h00000000} /* (8, 18, 9) {real, imag} */,
  {32'hc594de3c, 32'h00000000} /* (8, 18, 8) {real, imag} */,
  {32'hc5b04ab8, 32'h00000000} /* (8, 18, 7) {real, imag} */,
  {32'hc5b92941, 32'h00000000} /* (8, 18, 6) {real, imag} */,
  {32'hc5b52dcc, 32'h00000000} /* (8, 18, 5) {real, imag} */,
  {32'hc5d264ca, 32'h00000000} /* (8, 18, 4) {real, imag} */,
  {32'hc5fea3bb, 32'h00000000} /* (8, 18, 3) {real, imag} */,
  {32'hc5ece3a7, 32'h00000000} /* (8, 18, 2) {real, imag} */,
  {32'hc5e7b55d, 32'h00000000} /* (8, 18, 1) {real, imag} */,
  {32'hc5d1959c, 32'h00000000} /* (8, 18, 0) {real, imag} */,
  {32'hc5fb09e2, 32'h00000000} /* (8, 17, 31) {real, imag} */,
  {32'hc61a34d0, 32'h00000000} /* (8, 17, 30) {real, imag} */,
  {32'hc60a820a, 32'h00000000} /* (8, 17, 29) {real, imag} */,
  {32'hc5fe6192, 32'h00000000} /* (8, 17, 28) {real, imag} */,
  {32'hc5f77fbd, 32'h00000000} /* (8, 17, 27) {real, imag} */,
  {32'hc5dac325, 32'h00000000} /* (8, 17, 26) {real, imag} */,
  {32'hc5d50a15, 32'h00000000} /* (8, 17, 25) {real, imag} */,
  {32'hc5d96097, 32'h00000000} /* (8, 17, 24) {real, imag} */,
  {32'hc5d06348, 32'h00000000} /* (8, 17, 23) {real, imag} */,
  {32'hc55371b2, 32'h00000000} /* (8, 17, 22) {real, imag} */,
  {32'h43d1e200, 32'h00000000} /* (8, 17, 21) {real, imag} */,
  {32'h45226f39, 32'h00000000} /* (8, 17, 20) {real, imag} */,
  {32'h4566f7da, 32'h00000000} /* (8, 17, 19) {real, imag} */,
  {32'h45a40304, 32'h00000000} /* (8, 17, 18) {real, imag} */,
  {32'h45bfb6e1, 32'h00000000} /* (8, 17, 17) {real, imag} */,
  {32'h45e4a8f4, 32'h00000000} /* (8, 17, 16) {real, imag} */,
  {32'h45cf2e8a, 32'h00000000} /* (8, 17, 15) {real, imag} */,
  {32'h45c63f60, 32'h00000000} /* (8, 17, 14) {real, imag} */,
  {32'h45a1b71e, 32'h00000000} /* (8, 17, 13) {real, imag} */,
  {32'h45585ca1, 32'h00000000} /* (8, 17, 12) {real, imag} */,
  {32'h448a183c, 32'h00000000} /* (8, 17, 11) {real, imag} */,
  {32'hc4a239fc, 32'h00000000} /* (8, 17, 10) {real, imag} */,
  {32'hc550f12e, 32'h00000000} /* (8, 17, 9) {real, imag} */,
  {32'hc5b2f7f9, 32'h00000000} /* (8, 17, 8) {real, imag} */,
  {32'hc5bf39c0, 32'h00000000} /* (8, 17, 7) {real, imag} */,
  {32'hc5e84da3, 32'h00000000} /* (8, 17, 6) {real, imag} */,
  {32'hc5ee90f3, 32'h00000000} /* (8, 17, 5) {real, imag} */,
  {32'hc6057605, 32'h00000000} /* (8, 17, 4) {real, imag} */,
  {32'hc616bc9e, 32'h00000000} /* (8, 17, 3) {real, imag} */,
  {32'hc606742e, 32'h00000000} /* (8, 17, 2) {real, imag} */,
  {32'hc6004860, 32'h00000000} /* (8, 17, 1) {real, imag} */,
  {32'hc5e7864e, 32'h00000000} /* (8, 17, 0) {real, imag} */,
  {32'hc600919d, 32'h00000000} /* (8, 16, 31) {real, imag} */,
  {32'hc61997ab, 32'h00000000} /* (8, 16, 30) {real, imag} */,
  {32'hc6061361, 32'h00000000} /* (8, 16, 29) {real, imag} */,
  {32'hc6081918, 32'h00000000} /* (8, 16, 28) {real, imag} */,
  {32'hc60739b9, 32'h00000000} /* (8, 16, 27) {real, imag} */,
  {32'hc5e45422, 32'h00000000} /* (8, 16, 26) {real, imag} */,
  {32'hc5e23e82, 32'h00000000} /* (8, 16, 25) {real, imag} */,
  {32'hc5cdee78, 32'h00000000} /* (8, 16, 24) {real, imag} */,
  {32'hc5b15c0a, 32'h00000000} /* (8, 16, 23) {real, imag} */,
  {32'hc55a02d6, 32'h00000000} /* (8, 16, 22) {real, imag} */,
  {32'hc3ca3558, 32'h00000000} /* (8, 16, 21) {real, imag} */,
  {32'h452abf90, 32'h00000000} /* (8, 16, 20) {real, imag} */,
  {32'h458c59d8, 32'h00000000} /* (8, 16, 19) {real, imag} */,
  {32'h45c011ca, 32'h00000000} /* (8, 16, 18) {real, imag} */,
  {32'h45e15bdd, 32'h00000000} /* (8, 16, 17) {real, imag} */,
  {32'h45db1168, 32'h00000000} /* (8, 16, 16) {real, imag} */,
  {32'h45f9af4a, 32'h00000000} /* (8, 16, 15) {real, imag} */,
  {32'h45d29433, 32'h00000000} /* (8, 16, 14) {real, imag} */,
  {32'h45c09a75, 32'h00000000} /* (8, 16, 13) {real, imag} */,
  {32'h457dd3a4, 32'h00000000} /* (8, 16, 12) {real, imag} */,
  {32'h44aeecd2, 32'h00000000} /* (8, 16, 11) {real, imag} */,
  {32'hc48d149e, 32'h00000000} /* (8, 16, 10) {real, imag} */,
  {32'hc5814942, 32'h00000000} /* (8, 16, 9) {real, imag} */,
  {32'hc5b7575c, 32'h00000000} /* (8, 16, 8) {real, imag} */,
  {32'hc5c1a266, 32'h00000000} /* (8, 16, 7) {real, imag} */,
  {32'hc5eaacb9, 32'h00000000} /* (8, 16, 6) {real, imag} */,
  {32'hc5fa5256, 32'h00000000} /* (8, 16, 5) {real, imag} */,
  {32'hc60d7ffc, 32'h00000000} /* (8, 16, 4) {real, imag} */,
  {32'hc6149522, 32'h00000000} /* (8, 16, 3) {real, imag} */,
  {32'hc613ec77, 32'h00000000} /* (8, 16, 2) {real, imag} */,
  {32'hc60ebcbc, 32'h00000000} /* (8, 16, 1) {real, imag} */,
  {32'hc5f50914, 32'h00000000} /* (8, 16, 0) {real, imag} */,
  {32'hc6066564, 32'h00000000} /* (8, 15, 31) {real, imag} */,
  {32'hc6122302, 32'h00000000} /* (8, 15, 30) {real, imag} */,
  {32'hc6119e1a, 32'h00000000} /* (8, 15, 29) {real, imag} */,
  {32'hc601d6f2, 32'h00000000} /* (8, 15, 28) {real, imag} */,
  {32'hc5ecae45, 32'h00000000} /* (8, 15, 27) {real, imag} */,
  {32'hc5f852e3, 32'h00000000} /* (8, 15, 26) {real, imag} */,
  {32'hc5e18704, 32'h00000000} /* (8, 15, 25) {real, imag} */,
  {32'hc5e2b291, 32'h00000000} /* (8, 15, 24) {real, imag} */,
  {32'hc5a3d58b, 32'h00000000} /* (8, 15, 23) {real, imag} */,
  {32'hc53292c2, 32'h00000000} /* (8, 15, 22) {real, imag} */,
  {32'hc2e52ba0, 32'h00000000} /* (8, 15, 21) {real, imag} */,
  {32'h453ebc50, 32'h00000000} /* (8, 15, 20) {real, imag} */,
  {32'h4576ff9a, 32'h00000000} /* (8, 15, 19) {real, imag} */,
  {32'h45c455e9, 32'h00000000} /* (8, 15, 18) {real, imag} */,
  {32'h45eb8f04, 32'h00000000} /* (8, 15, 17) {real, imag} */,
  {32'h45ebe688, 32'h00000000} /* (8, 15, 16) {real, imag} */,
  {32'h45e0c91a, 32'h00000000} /* (8, 15, 15) {real, imag} */,
  {32'h45dee3f4, 32'h00000000} /* (8, 15, 14) {real, imag} */,
  {32'h45c0284f, 32'h00000000} /* (8, 15, 13) {real, imag} */,
  {32'h458b44b8, 32'h00000000} /* (8, 15, 12) {real, imag} */,
  {32'h44f3bc2c, 32'h00000000} /* (8, 15, 11) {real, imag} */,
  {32'hc4d05b94, 32'h00000000} /* (8, 15, 10) {real, imag} */,
  {32'hc5645409, 32'h00000000} /* (8, 15, 9) {real, imag} */,
  {32'hc5b52307, 32'h00000000} /* (8, 15, 8) {real, imag} */,
  {32'hc5fb5a91, 32'h00000000} /* (8, 15, 7) {real, imag} */,
  {32'hc5f359d7, 32'h00000000} /* (8, 15, 6) {real, imag} */,
  {32'hc5e9c274, 32'h00000000} /* (8, 15, 5) {real, imag} */,
  {32'hc60249c4, 32'h00000000} /* (8, 15, 4) {real, imag} */,
  {32'hc60a4258, 32'h00000000} /* (8, 15, 3) {real, imag} */,
  {32'hc60dbb22, 32'h00000000} /* (8, 15, 2) {real, imag} */,
  {32'hc602bd13, 32'h00000000} /* (8, 15, 1) {real, imag} */,
  {32'hc5f38fa6, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'hc5d2b620, 32'h00000000} /* (8, 14, 31) {real, imag} */,
  {32'hc5eaa245, 32'h00000000} /* (8, 14, 30) {real, imag} */,
  {32'hc5e6703c, 32'h00000000} /* (8, 14, 29) {real, imag} */,
  {32'hc5fb6434, 32'h00000000} /* (8, 14, 28) {real, imag} */,
  {32'hc5f2cb6c, 32'h00000000} /* (8, 14, 27) {real, imag} */,
  {32'hc5ef9e76, 32'h00000000} /* (8, 14, 26) {real, imag} */,
  {32'hc5ee444e, 32'h00000000} /* (8, 14, 25) {real, imag} */,
  {32'hc5af6bd6, 32'h00000000} /* (8, 14, 24) {real, imag} */,
  {32'hc59a2eaa, 32'h00000000} /* (8, 14, 23) {real, imag} */,
  {32'hc57483bb, 32'h00000000} /* (8, 14, 22) {real, imag} */,
  {32'hc43f3f48, 32'h00000000} /* (8, 14, 21) {real, imag} */,
  {32'h4508849a, 32'h00000000} /* (8, 14, 20) {real, imag} */,
  {32'h4563cde4, 32'h00000000} /* (8, 14, 19) {real, imag} */,
  {32'h45a15b8d, 32'h00000000} /* (8, 14, 18) {real, imag} */,
  {32'h45c3ffea, 32'h00000000} /* (8, 14, 17) {real, imag} */,
  {32'h45bb82c7, 32'h00000000} /* (8, 14, 16) {real, imag} */,
  {32'h45b90f7a, 32'h00000000} /* (8, 14, 15) {real, imag} */,
  {32'h45b14893, 32'h00000000} /* (8, 14, 14) {real, imag} */,
  {32'h45a2e8d4, 32'h00000000} /* (8, 14, 13) {real, imag} */,
  {32'h4556c19c, 32'h00000000} /* (8, 14, 12) {real, imag} */,
  {32'h44fe8cc8, 32'h00000000} /* (8, 14, 11) {real, imag} */,
  {32'hc4439aa4, 32'h00000000} /* (8, 14, 10) {real, imag} */,
  {32'hc58ec3c2, 32'h00000000} /* (8, 14, 9) {real, imag} */,
  {32'hc5c82004, 32'h00000000} /* (8, 14, 8) {real, imag} */,
  {32'hc5ed7c16, 32'h00000000} /* (8, 14, 7) {real, imag} */,
  {32'hc5e08394, 32'h00000000} /* (8, 14, 6) {real, imag} */,
  {32'hc5daca57, 32'h00000000} /* (8, 14, 5) {real, imag} */,
  {32'hc5ecb769, 32'h00000000} /* (8, 14, 4) {real, imag} */,
  {32'hc5f55bee, 32'h00000000} /* (8, 14, 3) {real, imag} */,
  {32'hc5f6a21b, 32'h00000000} /* (8, 14, 2) {real, imag} */,
  {32'hc5fb8136, 32'h00000000} /* (8, 14, 1) {real, imag} */,
  {32'hc5f0ceef, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'hc5b081f4, 32'h00000000} /* (8, 13, 31) {real, imag} */,
  {32'hc5c379c4, 32'h00000000} /* (8, 13, 30) {real, imag} */,
  {32'hc5b39a06, 32'h00000000} /* (8, 13, 29) {real, imag} */,
  {32'hc5be7f88, 32'h00000000} /* (8, 13, 28) {real, imag} */,
  {32'hc5d036d0, 32'h00000000} /* (8, 13, 27) {real, imag} */,
  {32'hc5c38716, 32'h00000000} /* (8, 13, 26) {real, imag} */,
  {32'hc5a87e29, 32'h00000000} /* (8, 13, 25) {real, imag} */,
  {32'hc59f23d6, 32'h00000000} /* (8, 13, 24) {real, imag} */,
  {32'hc56cb4b9, 32'h00000000} /* (8, 13, 23) {real, imag} */,
  {32'hc55f2e93, 32'h00000000} /* (8, 13, 22) {real, imag} */,
  {32'hc4477d8c, 32'h00000000} /* (8, 13, 21) {real, imag} */,
  {32'h4526ba3c, 32'h00000000} /* (8, 13, 20) {real, imag} */,
  {32'h455837f2, 32'h00000000} /* (8, 13, 19) {real, imag} */,
  {32'h4583e976, 32'h00000000} /* (8, 13, 18) {real, imag} */,
  {32'h45a257e9, 32'h00000000} /* (8, 13, 17) {real, imag} */,
  {32'h45b6336a, 32'h00000000} /* (8, 13, 16) {real, imag} */,
  {32'h45b8d882, 32'h00000000} /* (8, 13, 15) {real, imag} */,
  {32'h4597dedc, 32'h00000000} /* (8, 13, 14) {real, imag} */,
  {32'h458b122c, 32'h00000000} /* (8, 13, 13) {real, imag} */,
  {32'h457e7751, 32'h00000000} /* (8, 13, 12) {real, imag} */,
  {32'h450d74f9, 32'h00000000} /* (8, 13, 11) {real, imag} */,
  {32'hc4c9db6e, 32'h00000000} /* (8, 13, 10) {real, imag} */,
  {32'hc5738749, 32'h00000000} /* (8, 13, 9) {real, imag} */,
  {32'hc5a29f36, 32'h00000000} /* (8, 13, 8) {real, imag} */,
  {32'hc5ac859c, 32'h00000000} /* (8, 13, 7) {real, imag} */,
  {32'hc5d53746, 32'h00000000} /* (8, 13, 6) {real, imag} */,
  {32'hc5e9107a, 32'h00000000} /* (8, 13, 5) {real, imag} */,
  {32'hc5cbed36, 32'h00000000} /* (8, 13, 4) {real, imag} */,
  {32'hc5bf6c55, 32'h00000000} /* (8, 13, 3) {real, imag} */,
  {32'hc5d6c524, 32'h00000000} /* (8, 13, 2) {real, imag} */,
  {32'hc5d5294d, 32'h00000000} /* (8, 13, 1) {real, imag} */,
  {32'hc5b32ddc, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'hc5427b92, 32'h00000000} /* (8, 12, 31) {real, imag} */,
  {32'hc55bf1e0, 32'h00000000} /* (8, 12, 30) {real, imag} */,
  {32'hc581966c, 32'h00000000} /* (8, 12, 29) {real, imag} */,
  {32'hc5ab4670, 32'h00000000} /* (8, 12, 28) {real, imag} */,
  {32'hc59eceb1, 32'h00000000} /* (8, 12, 27) {real, imag} */,
  {32'hc596752a, 32'h00000000} /* (8, 12, 26) {real, imag} */,
  {32'hc58ca4f7, 32'h00000000} /* (8, 12, 25) {real, imag} */,
  {32'hc55a84cd, 32'h00000000} /* (8, 12, 24) {real, imag} */,
  {32'hc5145904, 32'h00000000} /* (8, 12, 23) {real, imag} */,
  {32'hc464ab90, 32'h00000000} /* (8, 12, 22) {real, imag} */,
  {32'h43f5dcd0, 32'h00000000} /* (8, 12, 21) {real, imag} */,
  {32'h454038b4, 32'h00000000} /* (8, 12, 20) {real, imag} */,
  {32'h45397800, 32'h00000000} /* (8, 12, 19) {real, imag} */,
  {32'h453f0f3d, 32'h00000000} /* (8, 12, 18) {real, imag} */,
  {32'h4582a01a, 32'h00000000} /* (8, 12, 17) {real, imag} */,
  {32'h4586f6bf, 32'h00000000} /* (8, 12, 16) {real, imag} */,
  {32'h459857ae, 32'h00000000} /* (8, 12, 15) {real, imag} */,
  {32'h45671836, 32'h00000000} /* (8, 12, 14) {real, imag} */,
  {32'h453c436c, 32'h00000000} /* (8, 12, 13) {real, imag} */,
  {32'h450a805f, 32'h00000000} /* (8, 12, 12) {real, imag} */,
  {32'h44842758, 32'h00000000} /* (8, 12, 11) {real, imag} */,
  {32'hc4a6792a, 32'h00000000} /* (8, 12, 10) {real, imag} */,
  {32'hc5766782, 32'h00000000} /* (8, 12, 9) {real, imag} */,
  {32'hc56cdc37, 32'h00000000} /* (8, 12, 8) {real, imag} */,
  {32'hc588329e, 32'h00000000} /* (8, 12, 7) {real, imag} */,
  {32'hc59a5440, 32'h00000000} /* (8, 12, 6) {real, imag} */,
  {32'hc599c41f, 32'h00000000} /* (8, 12, 5) {real, imag} */,
  {32'hc59cb2e5, 32'h00000000} /* (8, 12, 4) {real, imag} */,
  {32'hc5a7b284, 32'h00000000} /* (8, 12, 3) {real, imag} */,
  {32'hc5872828, 32'h00000000} /* (8, 12, 2) {real, imag} */,
  {32'hc56a92c6, 32'h00000000} /* (8, 12, 1) {real, imag} */,
  {32'hc561fe52, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'hc418bbd6, 32'h00000000} /* (8, 11, 31) {real, imag} */,
  {32'hc46860b9, 32'h00000000} /* (8, 11, 30) {real, imag} */,
  {32'hc4b2609c, 32'h00000000} /* (8, 11, 29) {real, imag} */,
  {32'hc526fc82, 32'h00000000} /* (8, 11, 28) {real, imag} */,
  {32'hc5215b82, 32'h00000000} /* (8, 11, 27) {real, imag} */,
  {32'hc4c5be50, 32'h00000000} /* (8, 11, 26) {real, imag} */,
  {32'hc4b62540, 32'h00000000} /* (8, 11, 25) {real, imag} */,
  {32'hc5005910, 32'h00000000} /* (8, 11, 24) {real, imag} */,
  {32'hc30bd3c0, 32'h00000000} /* (8, 11, 23) {real, imag} */,
  {32'h444828c0, 32'h00000000} /* (8, 11, 22) {real, imag} */,
  {32'h44d50e54, 32'h00000000} /* (8, 11, 21) {real, imag} */,
  {32'h44d1893d, 32'h00000000} /* (8, 11, 20) {real, imag} */,
  {32'h44e30d29, 32'h00000000} /* (8, 11, 19) {real, imag} */,
  {32'h44cc67b2, 32'h00000000} /* (8, 11, 18) {real, imag} */,
  {32'h44bd9399, 32'h00000000} /* (8, 11, 17) {real, imag} */,
  {32'h450dea04, 32'h00000000} /* (8, 11, 16) {real, imag} */,
  {32'h4506914c, 32'h00000000} /* (8, 11, 15) {real, imag} */,
  {32'h44cbca56, 32'h00000000} /* (8, 11, 14) {real, imag} */,
  {32'h44fa0760, 32'h00000000} /* (8, 11, 13) {real, imag} */,
  {32'h446811d8, 32'h00000000} /* (8, 11, 12) {real, imag} */,
  {32'h444c3050, 32'h00000000} /* (8, 11, 11) {real, imag} */,
  {32'hc4a633a8, 32'h00000000} /* (8, 11, 10) {real, imag} */,
  {32'hc52344b3, 32'h00000000} /* (8, 11, 9) {real, imag} */,
  {32'hc5304838, 32'h00000000} /* (8, 11, 8) {real, imag} */,
  {32'hc50a903c, 32'h00000000} /* (8, 11, 7) {real, imag} */,
  {32'hc5465862, 32'h00000000} /* (8, 11, 6) {real, imag} */,
  {32'hc54bf2c6, 32'h00000000} /* (8, 11, 5) {real, imag} */,
  {32'hc4cc54c1, 32'h00000000} /* (8, 11, 4) {real, imag} */,
  {32'hc4c923ab, 32'h00000000} /* (8, 11, 3) {real, imag} */,
  {32'hc520117f, 32'h00000000} /* (8, 11, 2) {real, imag} */,
  {32'hc5296d20, 32'h00000000} /* (8, 11, 1) {real, imag} */,
  {32'hc4baac0f, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h44d96f84, 32'h00000000} /* (8, 10, 31) {real, imag} */,
  {32'h4513776e, 32'h00000000} /* (8, 10, 30) {real, imag} */,
  {32'h44dc1ed0, 32'h00000000} /* (8, 10, 29) {real, imag} */,
  {32'h451e7d6a, 32'h00000000} /* (8, 10, 28) {real, imag} */,
  {32'h453b6c79, 32'h00000000} /* (8, 10, 27) {real, imag} */,
  {32'h4500e0cc, 32'h00000000} /* (8, 10, 26) {real, imag} */,
  {32'h450f7b26, 32'h00000000} /* (8, 10, 25) {real, imag} */,
  {32'h44ee840e, 32'h00000000} /* (8, 10, 24) {real, imag} */,
  {32'h457cddd6, 32'h00000000} /* (8, 10, 23) {real, imag} */,
  {32'h45439a72, 32'h00000000} /* (8, 10, 22) {real, imag} */,
  {32'h452ec898, 32'h00000000} /* (8, 10, 21) {real, imag} */,
  {32'h4500e749, 32'h00000000} /* (8, 10, 20) {real, imag} */,
  {32'h43dcd430, 32'h00000000} /* (8, 10, 19) {real, imag} */,
  {32'hc42f8860, 32'h00000000} /* (8, 10, 18) {real, imag} */,
  {32'hc45f9cc0, 32'h00000000} /* (8, 10, 17) {real, imag} */,
  {32'hc3e6abdc, 32'h00000000} /* (8, 10, 16) {real, imag} */,
  {32'hc46e9cfc, 32'h00000000} /* (8, 10, 15) {real, imag} */,
  {32'hc463ca2e, 32'h00000000} /* (8, 10, 14) {real, imag} */,
  {32'hc46348e7, 32'h00000000} /* (8, 10, 13) {real, imag} */,
  {32'hc457853c, 32'h00000000} /* (8, 10, 12) {real, imag} */,
  {32'hc4b50d6a, 32'h00000000} /* (8, 10, 11) {real, imag} */,
  {32'hc44adbe8, 32'h00000000} /* (8, 10, 10) {real, imag} */,
  {32'hc37d5370, 32'h00000000} /* (8, 10, 9) {real, imag} */,
  {32'h44110b70, 32'h00000000} /* (8, 10, 8) {real, imag} */,
  {32'h441c4e36, 32'h00000000} /* (8, 10, 7) {real, imag} */,
  {32'h43951698, 32'h00000000} /* (8, 10, 6) {real, imag} */,
  {32'h432234b8, 32'h00000000} /* (8, 10, 5) {real, imag} */,
  {32'h44d60404, 32'h00000000} /* (8, 10, 4) {real, imag} */,
  {32'h44ffd046, 32'h00000000} /* (8, 10, 3) {real, imag} */,
  {32'h4459a564, 32'h00000000} /* (8, 10, 2) {real, imag} */,
  {32'h4494c06e, 32'h00000000} /* (8, 10, 1) {real, imag} */,
  {32'h44d20045, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'h458d7547, 32'h00000000} /* (8, 9, 31) {real, imag} */,
  {32'h459b44b0, 32'h00000000} /* (8, 9, 30) {real, imag} */,
  {32'h45b84e68, 32'h00000000} /* (8, 9, 29) {real, imag} */,
  {32'h45b1c9fe, 32'h00000000} /* (8, 9, 28) {real, imag} */,
  {32'h45adc19c, 32'h00000000} /* (8, 9, 27) {real, imag} */,
  {32'h459c55a6, 32'h00000000} /* (8, 9, 26) {real, imag} */,
  {32'h45b69bae, 32'h00000000} /* (8, 9, 25) {real, imag} */,
  {32'h45aae31e, 32'h00000000} /* (8, 9, 24) {real, imag} */,
  {32'h45ab39ec, 32'h00000000} /* (8, 9, 23) {real, imag} */,
  {32'h459403ac, 32'h00000000} /* (8, 9, 22) {real, imag} */,
  {32'h455ad7f5, 32'h00000000} /* (8, 9, 21) {real, imag} */,
  {32'h450a0699, 32'h00000000} /* (8, 9, 20) {real, imag} */,
  {32'hc4065034, 32'h00000000} /* (8, 9, 19) {real, imag} */,
  {32'hc4eb83ba, 32'h00000000} /* (8, 9, 18) {real, imag} */,
  {32'hc4e11255, 32'h00000000} /* (8, 9, 17) {real, imag} */,
  {32'hc528db2c, 32'h00000000} /* (8, 9, 16) {real, imag} */,
  {32'hc5610096, 32'h00000000} /* (8, 9, 15) {real, imag} */,
  {32'hc55eee3b, 32'h00000000} /* (8, 9, 14) {real, imag} */,
  {32'hc5a45f56, 32'h00000000} /* (8, 9, 13) {real, imag} */,
  {32'hc5528387, 32'h00000000} /* (8, 9, 12) {real, imag} */,
  {32'hc4cd486a, 32'h00000000} /* (8, 9, 11) {real, imag} */,
  {32'hc465a84c, 32'h00000000} /* (8, 9, 10) {real, imag} */,
  {32'h44886a22, 32'h00000000} /* (8, 9, 9) {real, imag} */,
  {32'h451d9d47, 32'h00000000} /* (8, 9, 8) {real, imag} */,
  {32'h45524860, 32'h00000000} /* (8, 9, 7) {real, imag} */,
  {32'h4537d916, 32'h00000000} /* (8, 9, 6) {real, imag} */,
  {32'h457aebb9, 32'h00000000} /* (8, 9, 5) {real, imag} */,
  {32'h457b9245, 32'h00000000} /* (8, 9, 4) {real, imag} */,
  {32'h4572e1f9, 32'h00000000} /* (8, 9, 3) {real, imag} */,
  {32'h4583e00c, 32'h00000000} /* (8, 9, 2) {real, imag} */,
  {32'h458c93c7, 32'h00000000} /* (8, 9, 1) {real, imag} */,
  {32'h45968f87, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'h45ec09a5, 32'h00000000} /* (8, 8, 31) {real, imag} */,
  {32'h45dc055f, 32'h00000000} /* (8, 8, 30) {real, imag} */,
  {32'h45fced3a, 32'h00000000} /* (8, 8, 29) {real, imag} */,
  {32'h45eb3ae4, 32'h00000000} /* (8, 8, 28) {real, imag} */,
  {32'h45e9d0e2, 32'h00000000} /* (8, 8, 27) {real, imag} */,
  {32'h4605b0ce, 32'h00000000} /* (8, 8, 26) {real, imag} */,
  {32'h45e82179, 32'h00000000} /* (8, 8, 25) {real, imag} */,
  {32'h4605e336, 32'h00000000} /* (8, 8, 24) {real, imag} */,
  {32'h45eb3c4e, 32'h00000000} /* (8, 8, 23) {real, imag} */,
  {32'h45cd4118, 32'h00000000} /* (8, 8, 22) {real, imag} */,
  {32'h4585abf1, 32'h00000000} /* (8, 8, 21) {real, imag} */,
  {32'h44ed4098, 32'h00000000} /* (8, 8, 20) {real, imag} */,
  {32'hc3b31930, 32'h00000000} /* (8, 8, 19) {real, imag} */,
  {32'hc503b44f, 32'h00000000} /* (8, 8, 18) {real, imag} */,
  {32'hc552193e, 32'h00000000} /* (8, 8, 17) {real, imag} */,
  {32'hc571e0c3, 32'h00000000} /* (8, 8, 16) {real, imag} */,
  {32'hc5a0fc69, 32'h00000000} /* (8, 8, 15) {real, imag} */,
  {32'hc5b2d73d, 32'h00000000} /* (8, 8, 14) {real, imag} */,
  {32'hc59f591e, 32'h00000000} /* (8, 8, 13) {real, imag} */,
  {32'hc57c56c8, 32'h00000000} /* (8, 8, 12) {real, imag} */,
  {32'hc5367569, 32'h00000000} /* (8, 8, 11) {real, imag} */,
  {32'hc1485000, 32'h00000000} /* (8, 8, 10) {real, imag} */,
  {32'h44b3d12c, 32'h00000000} /* (8, 8, 9) {real, imag} */,
  {32'h452a5d20, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'h4546fe44, 32'h00000000} /* (8, 8, 7) {real, imag} */,
  {32'h45a8781e, 32'h00000000} /* (8, 8, 6) {real, imag} */,
  {32'h45a08bc7, 32'h00000000} /* (8, 8, 5) {real, imag} */,
  {32'h45be87c6, 32'h00000000} /* (8, 8, 4) {real, imag} */,
  {32'h45bdd172, 32'h00000000} /* (8, 8, 3) {real, imag} */,
  {32'h45bed928, 32'h00000000} /* (8, 8, 2) {real, imag} */,
  {32'h45c77987, 32'h00000000} /* (8, 8, 1) {real, imag} */,
  {32'h45cc6cb6, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h45f17b1c, 32'h00000000} /* (8, 7, 31) {real, imag} */,
  {32'h46078a09, 32'h00000000} /* (8, 7, 30) {real, imag} */,
  {32'h46228e00, 32'h00000000} /* (8, 7, 29) {real, imag} */,
  {32'h46117b1e, 32'h00000000} /* (8, 7, 28) {real, imag} */,
  {32'h46166108, 32'h00000000} /* (8, 7, 27) {real, imag} */,
  {32'h460640bc, 32'h00000000} /* (8, 7, 26) {real, imag} */,
  {32'h460bb9cc, 32'h00000000} /* (8, 7, 25) {real, imag} */,
  {32'h461401d0, 32'h00000000} /* (8, 7, 24) {real, imag} */,
  {32'h460893b6, 32'h00000000} /* (8, 7, 23) {real, imag} */,
  {32'h45fd3ab5, 32'h00000000} /* (8, 7, 22) {real, imag} */,
  {32'h45a98cc0, 32'h00000000} /* (8, 7, 21) {real, imag} */,
  {32'h450525b6, 32'h00000000} /* (8, 7, 20) {real, imag} */,
  {32'hc3715b90, 32'h00000000} /* (8, 7, 19) {real, imag} */,
  {32'hc50c4bf6, 32'h00000000} /* (8, 7, 18) {real, imag} */,
  {32'hc559e6b5, 32'h00000000} /* (8, 7, 17) {real, imag} */,
  {32'hc5961aa4, 32'h00000000} /* (8, 7, 16) {real, imag} */,
  {32'hc5bba932, 32'h00000000} /* (8, 7, 15) {real, imag} */,
  {32'hc5b1ef3e, 32'h00000000} /* (8, 7, 14) {real, imag} */,
  {32'hc5b74647, 32'h00000000} /* (8, 7, 13) {real, imag} */,
  {32'hc594e416, 32'h00000000} /* (8, 7, 12) {real, imag} */,
  {32'hc585b3e0, 32'h00000000} /* (8, 7, 11) {real, imag} */,
  {32'hc44c8978, 32'h00000000} /* (8, 7, 10) {real, imag} */,
  {32'h44ec895e, 32'h00000000} /* (8, 7, 9) {real, imag} */,
  {32'h458a62ac, 32'h00000000} /* (8, 7, 8) {real, imag} */,
  {32'h4589d1d4, 32'h00000000} /* (8, 7, 7) {real, imag} */,
  {32'h4593a313, 32'h00000000} /* (8, 7, 6) {real, imag} */,
  {32'h45c60d04, 32'h00000000} /* (8, 7, 5) {real, imag} */,
  {32'h45deb26b, 32'h00000000} /* (8, 7, 4) {real, imag} */,
  {32'h45fb1acc, 32'h00000000} /* (8, 7, 3) {real, imag} */,
  {32'h45f207df, 32'h00000000} /* (8, 7, 2) {real, imag} */,
  {32'h4603547f, 32'h00000000} /* (8, 7, 1) {real, imag} */,
  {32'h460777de, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h460f6e64, 32'h00000000} /* (8, 6, 31) {real, imag} */,
  {32'h461907a2, 32'h00000000} /* (8, 6, 30) {real, imag} */,
  {32'h461ef6da, 32'h00000000} /* (8, 6, 29) {real, imag} */,
  {32'h462708f8, 32'h00000000} /* (8, 6, 28) {real, imag} */,
  {32'h4624d71e, 32'h00000000} /* (8, 6, 27) {real, imag} */,
  {32'h4629d91e, 32'h00000000} /* (8, 6, 26) {real, imag} */,
  {32'h461f5438, 32'h00000000} /* (8, 6, 25) {real, imag} */,
  {32'h461ebe86, 32'h00000000} /* (8, 6, 24) {real, imag} */,
  {32'h46178c78, 32'h00000000} /* (8, 6, 23) {real, imag} */,
  {32'h460322c6, 32'h00000000} /* (8, 6, 22) {real, imag} */,
  {32'h45d2a1f9, 32'h00000000} /* (8, 6, 21) {real, imag} */,
  {32'h455a08ec, 32'h00000000} /* (8, 6, 20) {real, imag} */,
  {32'h43d165c8, 32'h00000000} /* (8, 6, 19) {real, imag} */,
  {32'hc41f6458, 32'h00000000} /* (8, 6, 18) {real, imag} */,
  {32'hc512ecfb, 32'h00000000} /* (8, 6, 17) {real, imag} */,
  {32'hc5886bae, 32'h00000000} /* (8, 6, 16) {real, imag} */,
  {32'hc5ab709f, 32'h00000000} /* (8, 6, 15) {real, imag} */,
  {32'hc5c9a892, 32'h00000000} /* (8, 6, 14) {real, imag} */,
  {32'hc5d1de1c, 32'h00000000} /* (8, 6, 13) {real, imag} */,
  {32'hc5c1a0d3, 32'h00000000} /* (8, 6, 12) {real, imag} */,
  {32'hc58893c0, 32'h00000000} /* (8, 6, 11) {real, imag} */,
  {32'hc4f17514, 32'h00000000} /* (8, 6, 10) {real, imag} */,
  {32'h43b5c2b0, 32'h00000000} /* (8, 6, 9) {real, imag} */,
  {32'h4524f5fa, 32'h00000000} /* (8, 6, 8) {real, imag} */,
  {32'h45555983, 32'h00000000} /* (8, 6, 7) {real, imag} */,
  {32'h45ac493c, 32'h00000000} /* (8, 6, 6) {real, imag} */,
  {32'h45c69473, 32'h00000000} /* (8, 6, 5) {real, imag} */,
  {32'h45ec8e68, 32'h00000000} /* (8, 6, 4) {real, imag} */,
  {32'h4605f1f0, 32'h00000000} /* (8, 6, 3) {real, imag} */,
  {32'h461c8e80, 32'h00000000} /* (8, 6, 2) {real, imag} */,
  {32'h460a2f43, 32'h00000000} /* (8, 6, 1) {real, imag} */,
  {32'h460dca32, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'h4624015e, 32'h00000000} /* (8, 5, 31) {real, imag} */,
  {32'h4620db3b, 32'h00000000} /* (8, 5, 30) {real, imag} */,
  {32'h463453fc, 32'h00000000} /* (8, 5, 29) {real, imag} */,
  {32'h463a56f6, 32'h00000000} /* (8, 5, 28) {real, imag} */,
  {32'h463cca6e, 32'h00000000} /* (8, 5, 27) {real, imag} */,
  {32'h463bf334, 32'h00000000} /* (8, 5, 26) {real, imag} */,
  {32'h463680df, 32'h00000000} /* (8, 5, 25) {real, imag} */,
  {32'h462d178d, 32'h00000000} /* (8, 5, 24) {real, imag} */,
  {32'h4625d9f6, 32'h00000000} /* (8, 5, 23) {real, imag} */,
  {32'h46251df9, 32'h00000000} /* (8, 5, 22) {real, imag} */,
  {32'h45f5cdee, 32'h00000000} /* (8, 5, 21) {real, imag} */,
  {32'h45cb9528, 32'h00000000} /* (8, 5, 20) {real, imag} */,
  {32'h45931f44, 32'h00000000} /* (8, 5, 19) {real, imag} */,
  {32'h45058509, 32'h00000000} /* (8, 5, 18) {real, imag} */,
  {32'h43920400, 32'h00000000} /* (8, 5, 17) {real, imag} */,
  {32'hc50eeac4, 32'h00000000} /* (8, 5, 16) {real, imag} */,
  {32'hc5925029, 32'h00000000} /* (8, 5, 15) {real, imag} */,
  {32'hc5c846ea, 32'h00000000} /* (8, 5, 14) {real, imag} */,
  {32'hc5cac77c, 32'h00000000} /* (8, 5, 13) {real, imag} */,
  {32'hc5b52898, 32'h00000000} /* (8, 5, 12) {real, imag} */,
  {32'hc59cb624, 32'h00000000} /* (8, 5, 11) {real, imag} */,
  {32'hc55bb13e, 32'h00000000} /* (8, 5, 10) {real, imag} */,
  {32'hc4c42868, 32'h00000000} /* (8, 5, 9) {real, imag} */,
  {32'hc3bd70c0, 32'h00000000} /* (8, 5, 8) {real, imag} */,
  {32'h451a8cda, 32'h00000000} /* (8, 5, 7) {real, imag} */,
  {32'h451677c5, 32'h00000000} /* (8, 5, 6) {real, imag} */,
  {32'h45c7184e, 32'h00000000} /* (8, 5, 5) {real, imag} */,
  {32'h45f23c80, 32'h00000000} /* (8, 5, 4) {real, imag} */,
  {32'h460226e4, 32'h00000000} /* (8, 5, 3) {real, imag} */,
  {32'h461b0b62, 32'h00000000} /* (8, 5, 2) {real, imag} */,
  {32'h46319a12, 32'h00000000} /* (8, 5, 1) {real, imag} */,
  {32'h462d97dc, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'h46283d82, 32'h00000000} /* (8, 4, 31) {real, imag} */,
  {32'h4631217e, 32'h00000000} /* (8, 4, 30) {real, imag} */,
  {32'h462b552e, 32'h00000000} /* (8, 4, 29) {real, imag} */,
  {32'h4640e90e, 32'h00000000} /* (8, 4, 28) {real, imag} */,
  {32'h465515f6, 32'h00000000} /* (8, 4, 27) {real, imag} */,
  {32'h46387268, 32'h00000000} /* (8, 4, 26) {real, imag} */,
  {32'h4634663e, 32'h00000000} /* (8, 4, 25) {real, imag} */,
  {32'h46323d3c, 32'h00000000} /* (8, 4, 24) {real, imag} */,
  {32'h462bc792, 32'h00000000} /* (8, 4, 23) {real, imag} */,
  {32'h462d3fc6, 32'h00000000} /* (8, 4, 22) {real, imag} */,
  {32'h4614014c, 32'h00000000} /* (8, 4, 21) {real, imag} */,
  {32'h45f96a53, 32'h00000000} /* (8, 4, 20) {real, imag} */,
  {32'h45b1d074, 32'h00000000} /* (8, 4, 19) {real, imag} */,
  {32'h4579e878, 32'h00000000} /* (8, 4, 18) {real, imag} */,
  {32'h4519768c, 32'h00000000} /* (8, 4, 17) {real, imag} */,
  {32'hc2da3a00, 32'h00000000} /* (8, 4, 16) {real, imag} */,
  {32'hc570676c, 32'h00000000} /* (8, 4, 15) {real, imag} */,
  {32'hc592260e, 32'h00000000} /* (8, 4, 14) {real, imag} */,
  {32'hc5a247b7, 32'h00000000} /* (8, 4, 13) {real, imag} */,
  {32'hc5c9a419, 32'h00000000} /* (8, 4, 12) {real, imag} */,
  {32'hc5b81d51, 32'h00000000} /* (8, 4, 11) {real, imag} */,
  {32'hc580d9d5, 32'h00000000} /* (8, 4, 10) {real, imag} */,
  {32'hc550cd76, 32'h00000000} /* (8, 4, 9) {real, imag} */,
  {32'hc4da42ac, 32'h00000000} /* (8, 4, 8) {real, imag} */,
  {32'h43e82e70, 32'h00000000} /* (8, 4, 7) {real, imag} */,
  {32'h44f8be24, 32'h00000000} /* (8, 4, 6) {real, imag} */,
  {32'h45a476cb, 32'h00000000} /* (8, 4, 5) {real, imag} */,
  {32'h45e947d7, 32'h00000000} /* (8, 4, 4) {real, imag} */,
  {32'h46143dcd, 32'h00000000} /* (8, 4, 3) {real, imag} */,
  {32'h4623bc1f, 32'h00000000} /* (8, 4, 2) {real, imag} */,
  {32'h462ee290, 32'h00000000} /* (8, 4, 1) {real, imag} */,
  {32'h4629da23, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'h463037a9, 32'h00000000} /* (8, 3, 31) {real, imag} */,
  {32'h4638b458, 32'h00000000} /* (8, 3, 30) {real, imag} */,
  {32'h4643680d, 32'h00000000} /* (8, 3, 29) {real, imag} */,
  {32'h463d6693, 32'h00000000} /* (8, 3, 28) {real, imag} */,
  {32'h46429bca, 32'h00000000} /* (8, 3, 27) {real, imag} */,
  {32'h464ac746, 32'h00000000} /* (8, 3, 26) {real, imag} */,
  {32'h4648d2ac, 32'h00000000} /* (8, 3, 25) {real, imag} */,
  {32'h4649a7d4, 32'h00000000} /* (8, 3, 24) {real, imag} */,
  {32'h462c4098, 32'h00000000} /* (8, 3, 23) {real, imag} */,
  {32'h461bfa20, 32'h00000000} /* (8, 3, 22) {real, imag} */,
  {32'h46187bc2, 32'h00000000} /* (8, 3, 21) {real, imag} */,
  {32'h45f24b8b, 32'h00000000} /* (8, 3, 20) {real, imag} */,
  {32'h45e21f5d, 32'h00000000} /* (8, 3, 19) {real, imag} */,
  {32'h459c1cf0, 32'h00000000} /* (8, 3, 18) {real, imag} */,
  {32'h45131ab6, 32'h00000000} /* (8, 3, 17) {real, imag} */,
  {32'h42fb34c0, 32'h00000000} /* (8, 3, 16) {real, imag} */,
  {32'hc5223068, 32'h00000000} /* (8, 3, 15) {real, imag} */,
  {32'hc5772787, 32'h00000000} /* (8, 3, 14) {real, imag} */,
  {32'hc5b71d0a, 32'h00000000} /* (8, 3, 13) {real, imag} */,
  {32'hc5ebbf8a, 32'h00000000} /* (8, 3, 12) {real, imag} */,
  {32'hc5a57664, 32'h00000000} /* (8, 3, 11) {real, imag} */,
  {32'hc58cc8f7, 32'h00000000} /* (8, 3, 10) {real, imag} */,
  {32'hc5845e0b, 32'h00000000} /* (8, 3, 9) {real, imag} */,
  {32'hc51a3682, 32'h00000000} /* (8, 3, 8) {real, imag} */,
  {32'hc4b9a98c, 32'h00000000} /* (8, 3, 7) {real, imag} */,
  {32'h44192138, 32'h00000000} /* (8, 3, 6) {real, imag} */,
  {32'h4588f579, 32'h00000000} /* (8, 3, 5) {real, imag} */,
  {32'h45e6d195, 32'h00000000} /* (8, 3, 4) {real, imag} */,
  {32'h46164090, 32'h00000000} /* (8, 3, 3) {real, imag} */,
  {32'h461b9623, 32'h00000000} /* (8, 3, 2) {real, imag} */,
  {32'h4630af82, 32'h00000000} /* (8, 3, 1) {real, imag} */,
  {32'h462793fe, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'h46325050, 32'h00000000} /* (8, 2, 31) {real, imag} */,
  {32'h463cff34, 32'h00000000} /* (8, 2, 30) {real, imag} */,
  {32'h4646f81f, 32'h00000000} /* (8, 2, 29) {real, imag} */,
  {32'h46483b46, 32'h00000000} /* (8, 2, 28) {real, imag} */,
  {32'h46443cde, 32'h00000000} /* (8, 2, 27) {real, imag} */,
  {32'h464ed7b5, 32'h00000000} /* (8, 2, 26) {real, imag} */,
  {32'h464a2800, 32'h00000000} /* (8, 2, 25) {real, imag} */,
  {32'h46496042, 32'h00000000} /* (8, 2, 24) {real, imag} */,
  {32'h463c1c58, 32'h00000000} /* (8, 2, 23) {real, imag} */,
  {32'h461d30e5, 32'h00000000} /* (8, 2, 22) {real, imag} */,
  {32'h4608ba26, 32'h00000000} /* (8, 2, 21) {real, imag} */,
  {32'h45f7c116, 32'h00000000} /* (8, 2, 20) {real, imag} */,
  {32'h45e70b3d, 32'h00000000} /* (8, 2, 19) {real, imag} */,
  {32'h45920adc, 32'h00000000} /* (8, 2, 18) {real, imag} */,
  {32'h4556f390, 32'h00000000} /* (8, 2, 17) {real, imag} */,
  {32'h447e7400, 32'h00000000} /* (8, 2, 16) {real, imag} */,
  {32'hc50498e8, 32'h00000000} /* (8, 2, 15) {real, imag} */,
  {32'hc5842de7, 32'h00000000} /* (8, 2, 14) {real, imag} */,
  {32'hc5b6f7e6, 32'h00000000} /* (8, 2, 13) {real, imag} */,
  {32'hc5b8fbb0, 32'h00000000} /* (8, 2, 12) {real, imag} */,
  {32'hc5b39de9, 32'h00000000} /* (8, 2, 11) {real, imag} */,
  {32'hc5b22ae6, 32'h00000000} /* (8, 2, 10) {real, imag} */,
  {32'hc5a2c908, 32'h00000000} /* (8, 2, 9) {real, imag} */,
  {32'hc55121cc, 32'h00000000} /* (8, 2, 8) {real, imag} */,
  {32'hc49f0654, 32'h00000000} /* (8, 2, 7) {real, imag} */,
  {32'hc2f92c00, 32'h00000000} /* (8, 2, 6) {real, imag} */,
  {32'h45c1da70, 32'h00000000} /* (8, 2, 5) {real, imag} */,
  {32'h4601bef9, 32'h00000000} /* (8, 2, 4) {real, imag} */,
  {32'h4614afce, 32'h00000000} /* (8, 2, 3) {real, imag} */,
  {32'h462f59e6, 32'h00000000} /* (8, 2, 2) {real, imag} */,
  {32'h463859ce, 32'h00000000} /* (8, 2, 1) {real, imag} */,
  {32'h462db16b, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'h462f103a, 32'h00000000} /* (8, 1, 31) {real, imag} */,
  {32'h463647b3, 32'h00000000} /* (8, 1, 30) {real, imag} */,
  {32'h464229dc, 32'h00000000} /* (8, 1, 29) {real, imag} */,
  {32'h46442ad4, 32'h00000000} /* (8, 1, 28) {real, imag} */,
  {32'h464f047c, 32'h00000000} /* (8, 1, 27) {real, imag} */,
  {32'h464d06ef, 32'h00000000} /* (8, 1, 26) {real, imag} */,
  {32'h464dab4c, 32'h00000000} /* (8, 1, 25) {real, imag} */,
  {32'h464319cb, 32'h00000000} /* (8, 1, 24) {real, imag} */,
  {32'h462c7408, 32'h00000000} /* (8, 1, 23) {real, imag} */,
  {32'h4607179a, 32'h00000000} /* (8, 1, 22) {real, imag} */,
  {32'h45fe70c0, 32'h00000000} /* (8, 1, 21) {real, imag} */,
  {32'h45e9071c, 32'h00000000} /* (8, 1, 20) {real, imag} */,
  {32'h45b2adf6, 32'h00000000} /* (8, 1, 19) {real, imag} */,
  {32'h4584a9aa, 32'h00000000} /* (8, 1, 18) {real, imag} */,
  {32'h450f5818, 32'h00000000} /* (8, 1, 17) {real, imag} */,
  {32'h445bb4a8, 32'h00000000} /* (8, 1, 16) {real, imag} */,
  {32'hc50365fe, 32'h00000000} /* (8, 1, 15) {real, imag} */,
  {32'hc59502da, 32'h00000000} /* (8, 1, 14) {real, imag} */,
  {32'hc59a34e9, 32'h00000000} /* (8, 1, 13) {real, imag} */,
  {32'hc5b9ccfc, 32'h00000000} /* (8, 1, 12) {real, imag} */,
  {32'hc59a8ec9, 32'h00000000} /* (8, 1, 11) {real, imag} */,
  {32'hc5707ab4, 32'h00000000} /* (8, 1, 10) {real, imag} */,
  {32'hc5919a90, 32'h00000000} /* (8, 1, 9) {real, imag} */,
  {32'hc50db61c, 32'h00000000} /* (8, 1, 8) {real, imag} */,
  {32'hc3f4f820, 32'h00000000} /* (8, 1, 7) {real, imag} */,
  {32'h44cbe38c, 32'h00000000} /* (8, 1, 6) {real, imag} */,
  {32'h45a095d2, 32'h00000000} /* (8, 1, 5) {real, imag} */,
  {32'h45f0e3d4, 32'h00000000} /* (8, 1, 4) {real, imag} */,
  {32'h461855e4, 32'h00000000} /* (8, 1, 3) {real, imag} */,
  {32'h4626451b, 32'h00000000} /* (8, 1, 2) {real, imag} */,
  {32'h462ae7ae, 32'h00000000} /* (8, 1, 1) {real, imag} */,
  {32'h462c58b0, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'h462752ec, 32'h00000000} /* (8, 0, 31) {real, imag} */,
  {32'h46326e3d, 32'h00000000} /* (8, 0, 30) {real, imag} */,
  {32'h463fe1d4, 32'h00000000} /* (8, 0, 29) {real, imag} */,
  {32'h4638459f, 32'h00000000} /* (8, 0, 28) {real, imag} */,
  {32'h46454342, 32'h00000000} /* (8, 0, 27) {real, imag} */,
  {32'h46421727, 32'h00000000} /* (8, 0, 26) {real, imag} */,
  {32'h463a9d36, 32'h00000000} /* (8, 0, 25) {real, imag} */,
  {32'h463ac910, 32'h00000000} /* (8, 0, 24) {real, imag} */,
  {32'h46129aa6, 32'h00000000} /* (8, 0, 23) {real, imag} */,
  {32'h46017dac, 32'h00000000} /* (8, 0, 22) {real, imag} */,
  {32'h45db33a6, 32'h00000000} /* (8, 0, 21) {real, imag} */,
  {32'h459fb36e, 32'h00000000} /* (8, 0, 20) {real, imag} */,
  {32'h45850ffe, 32'h00000000} /* (8, 0, 19) {real, imag} */,
  {32'h45425cf1, 32'h00000000} /* (8, 0, 18) {real, imag} */,
  {32'h449627f0, 32'h00000000} /* (8, 0, 17) {real, imag} */,
  {32'hc4300a88, 32'h00000000} /* (8, 0, 16) {real, imag} */,
  {32'hc528cbb6, 32'h00000000} /* (8, 0, 15) {real, imag} */,
  {32'hc59b5842, 32'h00000000} /* (8, 0, 14) {real, imag} */,
  {32'hc599d9d8, 32'h00000000} /* (8, 0, 13) {real, imag} */,
  {32'hc59be84a, 32'h00000000} /* (8, 0, 12) {real, imag} */,
  {32'hc5721be8, 32'h00000000} /* (8, 0, 11) {real, imag} */,
  {32'hc566d9ec, 32'h00000000} /* (8, 0, 10) {real, imag} */,
  {32'hc4f84510, 32'h00000000} /* (8, 0, 9) {real, imag} */,
  {32'hc4048680, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'h448910b0, 32'h00000000} /* (8, 0, 7) {real, imag} */,
  {32'h45599487, 32'h00000000} /* (8, 0, 6) {real, imag} */,
  {32'h45b130be, 32'h00000000} /* (8, 0, 5) {real, imag} */,
  {32'h45ea3f2e, 32'h00000000} /* (8, 0, 4) {real, imag} */,
  {32'h4616abaf, 32'h00000000} /* (8, 0, 3) {real, imag} */,
  {32'h4620137e, 32'h00000000} /* (8, 0, 2) {real, imag} */,
  {32'h4623a924, 32'h00000000} /* (8, 0, 1) {real, imag} */,
  {32'h4627e9b8, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h4614ee4e, 32'h00000000} /* (7, 31, 31) {real, imag} */,
  {32'h461e1c72, 32'h00000000} /* (7, 31, 30) {real, imag} */,
  {32'h46247ee5, 32'h00000000} /* (7, 31, 29) {real, imag} */,
  {32'h46220bb0, 32'h00000000} /* (7, 31, 28) {real, imag} */,
  {32'h46200cd7, 32'h00000000} /* (7, 31, 27) {real, imag} */,
  {32'h461c9892, 32'h00000000} /* (7, 31, 26) {real, imag} */,
  {32'h46189ea2, 32'h00000000} /* (7, 31, 25) {real, imag} */,
  {32'h46081b68, 32'h00000000} /* (7, 31, 24) {real, imag} */,
  {32'h45f775ae, 32'h00000000} /* (7, 31, 23) {real, imag} */,
  {32'h45cb75c6, 32'h00000000} /* (7, 31, 22) {real, imag} */,
  {32'h4593ef35, 32'h00000000} /* (7, 31, 21) {real, imag} */,
  {32'h450f0589, 32'h00000000} /* (7, 31, 20) {real, imag} */,
  {32'h44965b80, 32'h00000000} /* (7, 31, 19) {real, imag} */,
  {32'h41abf000, 32'h00000000} /* (7, 31, 18) {real, imag} */,
  {32'hc46cc988, 32'h00000000} /* (7, 31, 17) {real, imag} */,
  {32'hc4fbc90a, 32'h00000000} /* (7, 31, 16) {real, imag} */,
  {32'hc54071e0, 32'h00000000} /* (7, 31, 15) {real, imag} */,
  {32'hc559e8d6, 32'h00000000} /* (7, 31, 14) {real, imag} */,
  {32'hc560542c, 32'h00000000} /* (7, 31, 13) {real, imag} */,
  {32'hc57b6b9a, 32'h00000000} /* (7, 31, 12) {real, imag} */,
  {32'hc52b67b9, 32'h00000000} /* (7, 31, 11) {real, imag} */,
  {32'h430e3d00, 32'h00000000} /* (7, 31, 10) {real, imag} */,
  {32'h44628a80, 32'h00000000} /* (7, 31, 9) {real, imag} */,
  {32'h44bf00d4, 32'h00000000} /* (7, 31, 8) {real, imag} */,
  {32'h45907a4e, 32'h00000000} /* (7, 31, 7) {real, imag} */,
  {32'h45963c20, 32'h00000000} /* (7, 31, 6) {real, imag} */,
  {32'h45bc4167, 32'h00000000} /* (7, 31, 5) {real, imag} */,
  {32'h45dc4058, 32'h00000000} /* (7, 31, 4) {real, imag} */,
  {32'h46005648, 32'h00000000} /* (7, 31, 3) {real, imag} */,
  {32'h460a2f32, 32'h00000000} /* (7, 31, 2) {real, imag} */,
  {32'h4619f4ca, 32'h00000000} /* (7, 31, 1) {real, imag} */,
  {32'h46122ecf, 32'h00000000} /* (7, 31, 0) {real, imag} */,
  {32'h461ac09b, 32'h00000000} /* (7, 30, 31) {real, imag} */,
  {32'h462251b3, 32'h00000000} /* (7, 30, 30) {real, imag} */,
  {32'h462b4ca6, 32'h00000000} /* (7, 30, 29) {real, imag} */,
  {32'h462a55d0, 32'h00000000} /* (7, 30, 28) {real, imag} */,
  {32'h461fbc54, 32'h00000000} /* (7, 30, 27) {real, imag} */,
  {32'h4613923c, 32'h00000000} /* (7, 30, 26) {real, imag} */,
  {32'h460eb112, 32'h00000000} /* (7, 30, 25) {real, imag} */,
  {32'h46048e66, 32'h00000000} /* (7, 30, 24) {real, imag} */,
  {32'h4608b6a1, 32'h00000000} /* (7, 30, 23) {real, imag} */,
  {32'h45e00efa, 32'h00000000} /* (7, 30, 22) {real, imag} */,
  {32'h456cb8e1, 32'h00000000} /* (7, 30, 21) {real, imag} */,
  {32'h422b1780, 32'h00000000} /* (7, 30, 20) {real, imag} */,
  {32'hc4859d48, 32'h00000000} /* (7, 30, 19) {real, imag} */,
  {32'hc505f4f8, 32'h00000000} /* (7, 30, 18) {real, imag} */,
  {32'hc53b917c, 32'h00000000} /* (7, 30, 17) {real, imag} */,
  {32'hc5890b7e, 32'h00000000} /* (7, 30, 16) {real, imag} */,
  {32'hc5897652, 32'h00000000} /* (7, 30, 15) {real, imag} */,
  {32'hc595319e, 32'h00000000} /* (7, 30, 14) {real, imag} */,
  {32'hc589cc74, 32'h00000000} /* (7, 30, 13) {real, imag} */,
  {32'hc578de3e, 32'h00000000} /* (7, 30, 12) {real, imag} */,
  {32'hc52afef2, 32'h00000000} /* (7, 30, 11) {real, imag} */,
  {32'h432c6380, 32'h00000000} /* (7, 30, 10) {real, imag} */,
  {32'h44f74a24, 32'h00000000} /* (7, 30, 9) {real, imag} */,
  {32'h45828404, 32'h00000000} /* (7, 30, 8) {real, imag} */,
  {32'h45a6217b, 32'h00000000} /* (7, 30, 7) {real, imag} */,
  {32'h45d4bb42, 32'h00000000} /* (7, 30, 6) {real, imag} */,
  {32'h45ea5518, 32'h00000000} /* (7, 30, 5) {real, imag} */,
  {32'h460e9eae, 32'h00000000} /* (7, 30, 4) {real, imag} */,
  {32'h4608adee, 32'h00000000} /* (7, 30, 3) {real, imag} */,
  {32'h4625cf5e, 32'h00000000} /* (7, 30, 2) {real, imag} */,
  {32'h4622d595, 32'h00000000} /* (7, 30, 1) {real, imag} */,
  {32'h4613dabd, 32'h00000000} /* (7, 30, 0) {real, imag} */,
  {32'h46171c34, 32'h00000000} /* (7, 29, 31) {real, imag} */,
  {32'h461f6534, 32'h00000000} /* (7, 29, 30) {real, imag} */,
  {32'h46213ad2, 32'h00000000} /* (7, 29, 29) {real, imag} */,
  {32'h46209960, 32'h00000000} /* (7, 29, 28) {real, imag} */,
  {32'h46184020, 32'h00000000} /* (7, 29, 27) {real, imag} */,
  {32'h461213f0, 32'h00000000} /* (7, 29, 26) {real, imag} */,
  {32'h460c91c0, 32'h00000000} /* (7, 29, 25) {real, imag} */,
  {32'h45f72e18, 32'h00000000} /* (7, 29, 24) {real, imag} */,
  {32'h45dca524, 32'h00000000} /* (7, 29, 23) {real, imag} */,
  {32'h45b3035e, 32'h00000000} /* (7, 29, 22) {real, imag} */,
  {32'h4580943c, 32'h00000000} /* (7, 29, 21) {real, imag} */,
  {32'hc4a2cf58, 32'h00000000} /* (7, 29, 20) {real, imag} */,
  {32'hc4ed2c14, 32'h00000000} /* (7, 29, 19) {real, imag} */,
  {32'hc52977a2, 32'h00000000} /* (7, 29, 18) {real, imag} */,
  {32'hc571c75e, 32'h00000000} /* (7, 29, 17) {real, imag} */,
  {32'hc589935c, 32'h00000000} /* (7, 29, 16) {real, imag} */,
  {32'hc5a23cdc, 32'h00000000} /* (7, 29, 15) {real, imag} */,
  {32'hc5a52bdf, 32'h00000000} /* (7, 29, 14) {real, imag} */,
  {32'hc592dcf4, 32'h00000000} /* (7, 29, 13) {real, imag} */,
  {32'hc56a3356, 32'h00000000} /* (7, 29, 12) {real, imag} */,
  {32'hc504cf42, 32'h00000000} /* (7, 29, 11) {real, imag} */,
  {32'h449016fc, 32'h00000000} /* (7, 29, 10) {real, imag} */,
  {32'h4565e7a5, 32'h00000000} /* (7, 29, 9) {real, imag} */,
  {32'h45aa03d4, 32'h00000000} /* (7, 29, 8) {real, imag} */,
  {32'h45bdc150, 32'h00000000} /* (7, 29, 7) {real, imag} */,
  {32'h45edd248, 32'h00000000} /* (7, 29, 6) {real, imag} */,
  {32'h4612a400, 32'h00000000} /* (7, 29, 5) {real, imag} */,
  {32'h46143b09, 32'h00000000} /* (7, 29, 4) {real, imag} */,
  {32'h4621a490, 32'h00000000} /* (7, 29, 3) {real, imag} */,
  {32'h462d0be4, 32'h00000000} /* (7, 29, 2) {real, imag} */,
  {32'h461f99b4, 32'h00000000} /* (7, 29, 1) {real, imag} */,
  {32'h461cf984, 32'h00000000} /* (7, 29, 0) {real, imag} */,
  {32'h461a315f, 32'h00000000} /* (7, 28, 31) {real, imag} */,
  {32'h461a17ab, 32'h00000000} /* (7, 28, 30) {real, imag} */,
  {32'h4622ad66, 32'h00000000} /* (7, 28, 29) {real, imag} */,
  {32'h462a038e, 32'h00000000} /* (7, 28, 28) {real, imag} */,
  {32'h460b4bdf, 32'h00000000} /* (7, 28, 27) {real, imag} */,
  {32'h460a93ce, 32'h00000000} /* (7, 28, 26) {real, imag} */,
  {32'h46053789, 32'h00000000} /* (7, 28, 25) {real, imag} */,
  {32'h45f8af0c, 32'h00000000} /* (7, 28, 24) {real, imag} */,
  {32'h45da0d0d, 32'h00000000} /* (7, 28, 23) {real, imag} */,
  {32'h45a97771, 32'h00000000} /* (7, 28, 22) {real, imag} */,
  {32'h454cfb46, 32'h00000000} /* (7, 28, 21) {real, imag} */,
  {32'h441eb108, 32'h00000000} /* (7, 28, 20) {real, imag} */,
  {32'hc4abfb80, 32'h00000000} /* (7, 28, 19) {real, imag} */,
  {32'hc54aeda9, 32'h00000000} /* (7, 28, 18) {real, imag} */,
  {32'hc58537b2, 32'h00000000} /* (7, 28, 17) {real, imag} */,
  {32'hc58171a0, 32'h00000000} /* (7, 28, 16) {real, imag} */,
  {32'hc5a1f196, 32'h00000000} /* (7, 28, 15) {real, imag} */,
  {32'hc5a0a174, 32'h00000000} /* (7, 28, 14) {real, imag} */,
  {32'hc58d8461, 32'h00000000} /* (7, 28, 13) {real, imag} */,
  {32'hc539e141, 32'h00000000} /* (7, 28, 12) {real, imag} */,
  {32'hc496a01e, 32'h00000000} /* (7, 28, 11) {real, imag} */,
  {32'h446ced88, 32'h00000000} /* (7, 28, 10) {real, imag} */,
  {32'h4583422e, 32'h00000000} /* (7, 28, 9) {real, imag} */,
  {32'h45a2bd9c, 32'h00000000} /* (7, 28, 8) {real, imag} */,
  {32'h45f9e36b, 32'h00000000} /* (7, 28, 7) {real, imag} */,
  {32'h45efd4af, 32'h00000000} /* (7, 28, 6) {real, imag} */,
  {32'h460a9edc, 32'h00000000} /* (7, 28, 5) {real, imag} */,
  {32'h4613ff8e, 32'h00000000} /* (7, 28, 4) {real, imag} */,
  {32'h461f79ec, 32'h00000000} /* (7, 28, 3) {real, imag} */,
  {32'h4617d3ce, 32'h00000000} /* (7, 28, 2) {real, imag} */,
  {32'h46117827, 32'h00000000} /* (7, 28, 1) {real, imag} */,
  {32'h461368dc, 32'h00000000} /* (7, 28, 0) {real, imag} */,
  {32'h461a3d9f, 32'h00000000} /* (7, 27, 31) {real, imag} */,
  {32'h4614070c, 32'h00000000} /* (7, 27, 30) {real, imag} */,
  {32'h4614ccb3, 32'h00000000} /* (7, 27, 29) {real, imag} */,
  {32'h461c6b2a, 32'h00000000} /* (7, 27, 28) {real, imag} */,
  {32'h46129f98, 32'h00000000} /* (7, 27, 27) {real, imag} */,
  {32'h460dcf1a, 32'h00000000} /* (7, 27, 26) {real, imag} */,
  {32'h45f5f0d0, 32'h00000000} /* (7, 27, 25) {real, imag} */,
  {32'h4605683f, 32'h00000000} /* (7, 27, 24) {real, imag} */,
  {32'h45df9f8b, 32'h00000000} /* (7, 27, 23) {real, imag} */,
  {32'h45a70c16, 32'h00000000} /* (7, 27, 22) {real, imag} */,
  {32'h45456a14, 32'h00000000} /* (7, 27, 21) {real, imag} */,
  {32'hc414b960, 32'h00000000} /* (7, 27, 20) {real, imag} */,
  {32'hc5095435, 32'h00000000} /* (7, 27, 19) {real, imag} */,
  {32'hc563ad1c, 32'h00000000} /* (7, 27, 18) {real, imag} */,
  {32'hc593f697, 32'h00000000} /* (7, 27, 17) {real, imag} */,
  {32'hc5a997ca, 32'h00000000} /* (7, 27, 16) {real, imag} */,
  {32'hc5a872c6, 32'h00000000} /* (7, 27, 15) {real, imag} */,
  {32'hc59cb2a0, 32'h00000000} /* (7, 27, 14) {real, imag} */,
  {32'hc58d4a1a, 32'h00000000} /* (7, 27, 13) {real, imag} */,
  {32'hc556aa9a, 32'h00000000} /* (7, 27, 12) {real, imag} */,
  {32'hc4f728f6, 32'h00000000} /* (7, 27, 11) {real, imag} */,
  {32'h44d94c00, 32'h00000000} /* (7, 27, 10) {real, imag} */,
  {32'h458c65ac, 32'h00000000} /* (7, 27, 9) {real, imag} */,
  {32'h45b5ab6e, 32'h00000000} /* (7, 27, 8) {real, imag} */,
  {32'h45ecb4d1, 32'h00000000} /* (7, 27, 7) {real, imag} */,
  {32'h45ef6f16, 32'h00000000} /* (7, 27, 6) {real, imag} */,
  {32'h460a9c15, 32'h00000000} /* (7, 27, 5) {real, imag} */,
  {32'h4615f905, 32'h00000000} /* (7, 27, 4) {real, imag} */,
  {32'h461575fa, 32'h00000000} /* (7, 27, 3) {real, imag} */,
  {32'h460daf2b, 32'h00000000} /* (7, 27, 2) {real, imag} */,
  {32'h460f8e2e, 32'h00000000} /* (7, 27, 1) {real, imag} */,
  {32'h460fd4ed, 32'h00000000} /* (7, 27, 0) {real, imag} */,
  {32'h46029111, 32'h00000000} /* (7, 26, 31) {real, imag} */,
  {32'h46090cc6, 32'h00000000} /* (7, 26, 30) {real, imag} */,
  {32'h461b906b, 32'h00000000} /* (7, 26, 29) {real, imag} */,
  {32'h4619f84c, 32'h00000000} /* (7, 26, 28) {real, imag} */,
  {32'h46168799, 32'h00000000} /* (7, 26, 27) {real, imag} */,
  {32'h460f474f, 32'h00000000} /* (7, 26, 26) {real, imag} */,
  {32'h4609801c, 32'h00000000} /* (7, 26, 25) {real, imag} */,
  {32'h45f5014f, 32'h00000000} /* (7, 26, 24) {real, imag} */,
  {32'h45cc9a32, 32'h00000000} /* (7, 26, 23) {real, imag} */,
  {32'h45a52470, 32'h00000000} /* (7, 26, 22) {real, imag} */,
  {32'h4543a236, 32'h00000000} /* (7, 26, 21) {real, imag} */,
  {32'hc3c37070, 32'h00000000} /* (7, 26, 20) {real, imag} */,
  {32'hc51c1264, 32'h00000000} /* (7, 26, 19) {real, imag} */,
  {32'hc556c76b, 32'h00000000} /* (7, 26, 18) {real, imag} */,
  {32'hc58b8b28, 32'h00000000} /* (7, 26, 17) {real, imag} */,
  {32'hc5baafe3, 32'h00000000} /* (7, 26, 16) {real, imag} */,
  {32'hc5aee452, 32'h00000000} /* (7, 26, 15) {real, imag} */,
  {32'hc5aedd6f, 32'h00000000} /* (7, 26, 14) {real, imag} */,
  {32'hc599028c, 32'h00000000} /* (7, 26, 13) {real, imag} */,
  {32'hc5374366, 32'h00000000} /* (7, 26, 12) {real, imag} */,
  {32'hc40ffb50, 32'h00000000} /* (7, 26, 11) {real, imag} */,
  {32'h4507b164, 32'h00000000} /* (7, 26, 10) {real, imag} */,
  {32'h459a949c, 32'h00000000} /* (7, 26, 9) {real, imag} */,
  {32'h45b6a5af, 32'h00000000} /* (7, 26, 8) {real, imag} */,
  {32'h45d167fe, 32'h00000000} /* (7, 26, 7) {real, imag} */,
  {32'h45def472, 32'h00000000} /* (7, 26, 6) {real, imag} */,
  {32'h4600c49a, 32'h00000000} /* (7, 26, 5) {real, imag} */,
  {32'h4608576a, 32'h00000000} /* (7, 26, 4) {real, imag} */,
  {32'h460b5051, 32'h00000000} /* (7, 26, 3) {real, imag} */,
  {32'h4601eff1, 32'h00000000} /* (7, 26, 2) {real, imag} */,
  {32'h460c4b50, 32'h00000000} /* (7, 26, 1) {real, imag} */,
  {32'h4613417e, 32'h00000000} /* (7, 26, 0) {real, imag} */,
  {32'h4605c5c7, 32'h00000000} /* (7, 25, 31) {real, imag} */,
  {32'h460217e2, 32'h00000000} /* (7, 25, 30) {real, imag} */,
  {32'h46099710, 32'h00000000} /* (7, 25, 29) {real, imag} */,
  {32'h4609e237, 32'h00000000} /* (7, 25, 28) {real, imag} */,
  {32'h461098a2, 32'h00000000} /* (7, 25, 27) {real, imag} */,
  {32'h4610115e, 32'h00000000} /* (7, 25, 26) {real, imag} */,
  {32'h45f52b0e, 32'h00000000} /* (7, 25, 25) {real, imag} */,
  {32'h45e51782, 32'h00000000} /* (7, 25, 24) {real, imag} */,
  {32'h45ccfa4e, 32'h00000000} /* (7, 25, 23) {real, imag} */,
  {32'h4599e232, 32'h00000000} /* (7, 25, 22) {real, imag} */,
  {32'h452104c0, 32'h00000000} /* (7, 25, 21) {real, imag} */,
  {32'h43522e70, 32'h00000000} /* (7, 25, 20) {real, imag} */,
  {32'hc54daab2, 32'h00000000} /* (7, 25, 19) {real, imag} */,
  {32'hc54f6f05, 32'h00000000} /* (7, 25, 18) {real, imag} */,
  {32'hc58661b2, 32'h00000000} /* (7, 25, 17) {real, imag} */,
  {32'hc59d1b1a, 32'h00000000} /* (7, 25, 16) {real, imag} */,
  {32'hc59771b2, 32'h00000000} /* (7, 25, 15) {real, imag} */,
  {32'hc5c1981d, 32'h00000000} /* (7, 25, 14) {real, imag} */,
  {32'hc560ab0c, 32'h00000000} /* (7, 25, 13) {real, imag} */,
  {32'hc5578474, 32'h00000000} /* (7, 25, 12) {real, imag} */,
  {32'hc4ac9dbc, 32'h00000000} /* (7, 25, 11) {real, imag} */,
  {32'h451fb6aa, 32'h00000000} /* (7, 25, 10) {real, imag} */,
  {32'h45872790, 32'h00000000} /* (7, 25, 9) {real, imag} */,
  {32'h45d0617e, 32'h00000000} /* (7, 25, 8) {real, imag} */,
  {32'h45d3fb42, 32'h00000000} /* (7, 25, 7) {real, imag} */,
  {32'h45dbbc9c, 32'h00000000} /* (7, 25, 6) {real, imag} */,
  {32'h45eb23e0, 32'h00000000} /* (7, 25, 5) {real, imag} */,
  {32'h45f8b176, 32'h00000000} /* (7, 25, 4) {real, imag} */,
  {32'h45fd705f, 32'h00000000} /* (7, 25, 3) {real, imag} */,
  {32'h45f92a02, 32'h00000000} /* (7, 25, 2) {real, imag} */,
  {32'h45f2f512, 32'h00000000} /* (7, 25, 1) {real, imag} */,
  {32'h45e90b56, 32'h00000000} /* (7, 25, 0) {real, imag} */,
  {32'h45e2c66f, 32'h00000000} /* (7, 24, 31) {real, imag} */,
  {32'h45f72210, 32'h00000000} /* (7, 24, 30) {real, imag} */,
  {32'h45e641de, 32'h00000000} /* (7, 24, 29) {real, imag} */,
  {32'h45fedab7, 32'h00000000} /* (7, 24, 28) {real, imag} */,
  {32'h46038705, 32'h00000000} /* (7, 24, 27) {real, imag} */,
  {32'h45ecf34f, 32'h00000000} /* (7, 24, 26) {real, imag} */,
  {32'h45fc0014, 32'h00000000} /* (7, 24, 25) {real, imag} */,
  {32'h45da443f, 32'h00000000} /* (7, 24, 24) {real, imag} */,
  {32'h45be1371, 32'h00000000} /* (7, 24, 23) {real, imag} */,
  {32'h45a66f94, 32'h00000000} /* (7, 24, 22) {real, imag} */,
  {32'h45261986, 32'h00000000} /* (7, 24, 21) {real, imag} */,
  {32'hc472c840, 32'h00000000} /* (7, 24, 20) {real, imag} */,
  {32'hc4b33f6e, 32'h00000000} /* (7, 24, 19) {real, imag} */,
  {32'hc549ae18, 32'h00000000} /* (7, 24, 18) {real, imag} */,
  {32'hc57b588a, 32'h00000000} /* (7, 24, 17) {real, imag} */,
  {32'hc58f21b0, 32'h00000000} /* (7, 24, 16) {real, imag} */,
  {32'hc5a28d63, 32'h00000000} /* (7, 24, 15) {real, imag} */,
  {32'hc582b370, 32'h00000000} /* (7, 24, 14) {real, imag} */,
  {32'hc5a92724, 32'h00000000} /* (7, 24, 13) {real, imag} */,
  {32'hc539bdda, 32'h00000000} /* (7, 24, 12) {real, imag} */,
  {32'hc42a589c, 32'h00000000} /* (7, 24, 11) {real, imag} */,
  {32'h44a042f4, 32'h00000000} /* (7, 24, 10) {real, imag} */,
  {32'h45a4f040, 32'h00000000} /* (7, 24, 9) {real, imag} */,
  {32'h45acc5db, 32'h00000000} /* (7, 24, 8) {real, imag} */,
  {32'h45bfac47, 32'h00000000} /* (7, 24, 7) {real, imag} */,
  {32'h45d1c894, 32'h00000000} /* (7, 24, 6) {real, imag} */,
  {32'h45cd9103, 32'h00000000} /* (7, 24, 5) {real, imag} */,
  {32'h45dbe75c, 32'h00000000} /* (7, 24, 4) {real, imag} */,
  {32'h45eed818, 32'h00000000} /* (7, 24, 3) {real, imag} */,
  {32'h45f201d4, 32'h00000000} /* (7, 24, 2) {real, imag} */,
  {32'h45cf51e9, 32'h00000000} /* (7, 24, 1) {real, imag} */,
  {32'h45ca30cc, 32'h00000000} /* (7, 24, 0) {real, imag} */,
  {32'h45a70ac0, 32'h00000000} /* (7, 23, 31) {real, imag} */,
  {32'h45c5411b, 32'h00000000} /* (7, 23, 30) {real, imag} */,
  {32'h45cd4eff, 32'h00000000} /* (7, 23, 29) {real, imag} */,
  {32'h45cfc958, 32'h00000000} /* (7, 23, 28) {real, imag} */,
  {32'h45f01217, 32'h00000000} /* (7, 23, 27) {real, imag} */,
  {32'h45e04358, 32'h00000000} /* (7, 23, 26) {real, imag} */,
  {32'h45c20e6b, 32'h00000000} /* (7, 23, 25) {real, imag} */,
  {32'h45a66c2c, 32'h00000000} /* (7, 23, 24) {real, imag} */,
  {32'h45a29766, 32'h00000000} /* (7, 23, 23) {real, imag} */,
  {32'h45783c94, 32'h00000000} /* (7, 23, 22) {real, imag} */,
  {32'h450be6fe, 32'h00000000} /* (7, 23, 21) {real, imag} */,
  {32'hc0fde600, 32'h00000000} /* (7, 23, 20) {real, imag} */,
  {32'hc494d514, 32'h00000000} /* (7, 23, 19) {real, imag} */,
  {32'hc50c8dbe, 32'h00000000} /* (7, 23, 18) {real, imag} */,
  {32'hc536404e, 32'h00000000} /* (7, 23, 17) {real, imag} */,
  {32'hc540b97c, 32'h00000000} /* (7, 23, 16) {real, imag} */,
  {32'hc551bea4, 32'h00000000} /* (7, 23, 15) {real, imag} */,
  {32'hc568fbf2, 32'h00000000} /* (7, 23, 14) {real, imag} */,
  {32'hc582d759, 32'h00000000} /* (7, 23, 13) {real, imag} */,
  {32'hc505b1eb, 32'h00000000} /* (7, 23, 12) {real, imag} */,
  {32'hc3d94130, 32'h00000000} /* (7, 23, 11) {real, imag} */,
  {32'h44a80b38, 32'h00000000} /* (7, 23, 10) {real, imag} */,
  {32'h45625692, 32'h00000000} /* (7, 23, 9) {real, imag} */,
  {32'h4598b024, 32'h00000000} /* (7, 23, 8) {real, imag} */,
  {32'h45aa6f5a, 32'h00000000} /* (7, 23, 7) {real, imag} */,
  {32'h45ccd592, 32'h00000000} /* (7, 23, 6) {real, imag} */,
  {32'h45c78f53, 32'h00000000} /* (7, 23, 5) {real, imag} */,
  {32'h45b09bae, 32'h00000000} /* (7, 23, 4) {real, imag} */,
  {32'h45b183af, 32'h00000000} /* (7, 23, 3) {real, imag} */,
  {32'h45af4ad0, 32'h00000000} /* (7, 23, 2) {real, imag} */,
  {32'h45a585bf, 32'h00000000} /* (7, 23, 1) {real, imag} */,
  {32'h45a1b522, 32'h00000000} /* (7, 23, 0) {real, imag} */,
  {32'h45593c90, 32'h00000000} /* (7, 22, 31) {real, imag} */,
  {32'h456c5638, 32'h00000000} /* (7, 22, 30) {real, imag} */,
  {32'h459241d7, 32'h00000000} /* (7, 22, 29) {real, imag} */,
  {32'h45a6a10d, 32'h00000000} /* (7, 22, 28) {real, imag} */,
  {32'h45bcce95, 32'h00000000} /* (7, 22, 27) {real, imag} */,
  {32'h4596d39c, 32'h00000000} /* (7, 22, 26) {real, imag} */,
  {32'h45965966, 32'h00000000} /* (7, 22, 25) {real, imag} */,
  {32'h45799516, 32'h00000000} /* (7, 22, 24) {real, imag} */,
  {32'h456e998e, 32'h00000000} /* (7, 22, 23) {real, imag} */,
  {32'h457768d6, 32'h00000000} /* (7, 22, 22) {real, imag} */,
  {32'h44caeed6, 32'h00000000} /* (7, 22, 21) {real, imag} */,
  {32'h437bffc8, 32'h00000000} /* (7, 22, 20) {real, imag} */,
  {32'hc4a48b30, 32'h00000000} /* (7, 22, 19) {real, imag} */,
  {32'hc40ce128, 32'h00000000} /* (7, 22, 18) {real, imag} */,
  {32'hc4a1771f, 32'h00000000} /* (7, 22, 17) {real, imag} */,
  {32'hc530c490, 32'h00000000} /* (7, 22, 16) {real, imag} */,
  {32'hc4d7239f, 32'h00000000} /* (7, 22, 15) {real, imag} */,
  {32'hc51d05cc, 32'h00000000} /* (7, 22, 14) {real, imag} */,
  {32'hc50de308, 32'h00000000} /* (7, 22, 13) {real, imag} */,
  {32'hc50f5a22, 32'h00000000} /* (7, 22, 12) {real, imag} */,
  {32'hc4239f18, 32'h00000000} /* (7, 22, 11) {real, imag} */,
  {32'h44e1de10, 32'h00000000} /* (7, 22, 10) {real, imag} */,
  {32'h4531d7e3, 32'h00000000} /* (7, 22, 9) {real, imag} */,
  {32'h459c842b, 32'h00000000} /* (7, 22, 8) {real, imag} */,
  {32'h45953ff7, 32'h00000000} /* (7, 22, 7) {real, imag} */,
  {32'h45887b31, 32'h00000000} /* (7, 22, 6) {real, imag} */,
  {32'h4596d9de, 32'h00000000} /* (7, 22, 5) {real, imag} */,
  {32'h45640c66, 32'h00000000} /* (7, 22, 4) {real, imag} */,
  {32'h4563dd60, 32'h00000000} /* (7, 22, 3) {real, imag} */,
  {32'h45828037, 32'h00000000} /* (7, 22, 2) {real, imag} */,
  {32'h4538364c, 32'h00000000} /* (7, 22, 1) {real, imag} */,
  {32'h454252a0, 32'h00000000} /* (7, 22, 0) {real, imag} */,
  {32'h44a98b2e, 32'h00000000} /* (7, 21, 31) {real, imag} */,
  {32'h451bba06, 32'h00000000} /* (7, 21, 30) {real, imag} */,
  {32'h45096ed1, 32'h00000000} /* (7, 21, 29) {real, imag} */,
  {32'h45265862, 32'h00000000} /* (7, 21, 28) {real, imag} */,
  {32'h45743e21, 32'h00000000} /* (7, 21, 27) {real, imag} */,
  {32'h451f5ae0, 32'h00000000} /* (7, 21, 26) {real, imag} */,
  {32'h450d3383, 32'h00000000} /* (7, 21, 25) {real, imag} */,
  {32'h44a20253, 32'h00000000} /* (7, 21, 24) {real, imag} */,
  {32'h450cdce9, 32'h00000000} /* (7, 21, 23) {real, imag} */,
  {32'h44bf90f4, 32'h00000000} /* (7, 21, 22) {real, imag} */,
  {32'h44503464, 32'h00000000} /* (7, 21, 21) {real, imag} */,
  {32'hc3cd828f, 32'h00000000} /* (7, 21, 20) {real, imag} */,
  {32'h43860358, 32'h00000000} /* (7, 21, 19) {real, imag} */,
  {32'h4389e7b8, 32'h00000000} /* (7, 21, 18) {real, imag} */,
  {32'h43005308, 32'h00000000} /* (7, 21, 17) {real, imag} */,
  {32'h442ec4d3, 32'h00000000} /* (7, 21, 16) {real, imag} */,
  {32'hc30ee094, 32'h00000000} /* (7, 21, 15) {real, imag} */,
  {32'hc36b8900, 32'h00000000} /* (7, 21, 14) {real, imag} */,
  {32'h43a1d2e8, 32'h00000000} /* (7, 21, 13) {real, imag} */,
  {32'hc418410a, 32'h00000000} /* (7, 21, 12) {real, imag} */,
  {32'h43f85a48, 32'h00000000} /* (7, 21, 11) {real, imag} */,
  {32'h44a2f030, 32'h00000000} /* (7, 21, 10) {real, imag} */,
  {32'h4505a31d, 32'h00000000} /* (7, 21, 9) {real, imag} */,
  {32'h44fdbeb7, 32'h00000000} /* (7, 21, 8) {real, imag} */,
  {32'h45103cc9, 32'h00000000} /* (7, 21, 7) {real, imag} */,
  {32'h4487bc7c, 32'h00000000} /* (7, 21, 6) {real, imag} */,
  {32'h44209234, 32'h00000000} /* (7, 21, 5) {real, imag} */,
  {32'h44909ed7, 32'h00000000} /* (7, 21, 4) {real, imag} */,
  {32'h449e77c6, 32'h00000000} /* (7, 21, 3) {real, imag} */,
  {32'h44ad3d57, 32'h00000000} /* (7, 21, 2) {real, imag} */,
  {32'h449965d9, 32'h00000000} /* (7, 21, 1) {real, imag} */,
  {32'h4499437c, 32'h00000000} /* (7, 21, 0) {real, imag} */,
  {32'hc475918e, 32'h00000000} /* (7, 20, 31) {real, imag} */,
  {32'hc451c016, 32'h00000000} /* (7, 20, 30) {real, imag} */,
  {32'hc4d6e6a7, 32'h00000000} /* (7, 20, 29) {real, imag} */,
  {32'hc412ffb6, 32'h00000000} /* (7, 20, 28) {real, imag} */,
  {32'hc39de19d, 32'h00000000} /* (7, 20, 27) {real, imag} */,
  {32'hc463803d, 32'h00000000} /* (7, 20, 26) {real, imag} */,
  {32'hc4731e3a, 32'h00000000} /* (7, 20, 25) {real, imag} */,
  {32'hc4bab4b9, 32'h00000000} /* (7, 20, 24) {real, imag} */,
  {32'hc4f9f580, 32'h00000000} /* (7, 20, 23) {real, imag} */,
  {32'hc4f9ab88, 32'h00000000} /* (7, 20, 22) {real, imag} */,
  {32'hc32417dc, 32'h00000000} /* (7, 20, 21) {real, imag} */,
  {32'h444221a0, 32'h00000000} /* (7, 20, 20) {real, imag} */,
  {32'h44e67870, 32'h00000000} /* (7, 20, 19) {real, imag} */,
  {32'h45360bb3, 32'h00000000} /* (7, 20, 18) {real, imag} */,
  {32'h45273779, 32'h00000000} /* (7, 20, 17) {real, imag} */,
  {32'h451503c0, 32'h00000000} /* (7, 20, 16) {real, imag} */,
  {32'h450ac2b2, 32'h00000000} /* (7, 20, 15) {real, imag} */,
  {32'h45416fc6, 32'h00000000} /* (7, 20, 14) {real, imag} */,
  {32'h45028b35, 32'h00000000} /* (7, 20, 13) {real, imag} */,
  {32'h44f53d61, 32'h00000000} /* (7, 20, 12) {real, imag} */,
  {32'h44a4b0c3, 32'h00000000} /* (7, 20, 11) {real, imag} */,
  {32'h4298b9b0, 32'h00000000} /* (7, 20, 10) {real, imag} */,
  {32'hc484506d, 32'h00000000} /* (7, 20, 9) {real, imag} */,
  {32'hc4be50c3, 32'h00000000} /* (7, 20, 8) {real, imag} */,
  {32'hc4b5206e, 32'h00000000} /* (7, 20, 7) {real, imag} */,
  {32'hc50ccb82, 32'h00000000} /* (7, 20, 6) {real, imag} */,
  {32'hc4c42f34, 32'h00000000} /* (7, 20, 5) {real, imag} */,
  {32'hc4f5ebd8, 32'h00000000} /* (7, 20, 4) {real, imag} */,
  {32'hc53b66a0, 32'h00000000} /* (7, 20, 3) {real, imag} */,
  {32'hc509e649, 32'h00000000} /* (7, 20, 2) {real, imag} */,
  {32'hc517d2d1, 32'h00000000} /* (7, 20, 1) {real, imag} */,
  {32'hc4c0bf67, 32'h00000000} /* (7, 20, 0) {real, imag} */,
  {32'hc54848a1, 32'h00000000} /* (7, 19, 31) {real, imag} */,
  {32'hc53c9f1c, 32'h00000000} /* (7, 19, 30) {real, imag} */,
  {32'hc533fdb7, 32'h00000000} /* (7, 19, 29) {real, imag} */,
  {32'hc5559317, 32'h00000000} /* (7, 19, 28) {real, imag} */,
  {32'hc5359ac2, 32'h00000000} /* (7, 19, 27) {real, imag} */,
  {32'hc5628022, 32'h00000000} /* (7, 19, 26) {real, imag} */,
  {32'hc55abce0, 32'h00000000} /* (7, 19, 25) {real, imag} */,
  {32'hc5423bde, 32'h00000000} /* (7, 19, 24) {real, imag} */,
  {32'hc55f624d, 32'h00000000} /* (7, 19, 23) {real, imag} */,
  {32'hc531e1d9, 32'h00000000} /* (7, 19, 22) {real, imag} */,
  {32'hc2e6d680, 32'h00000000} /* (7, 19, 21) {real, imag} */,
  {32'h44d14cf0, 32'h00000000} /* (7, 19, 20) {real, imag} */,
  {32'h453d5de4, 32'h00000000} /* (7, 19, 19) {real, imag} */,
  {32'h4588139d, 32'h00000000} /* (7, 19, 18) {real, imag} */,
  {32'h459d9ffa, 32'h00000000} /* (7, 19, 17) {real, imag} */,
  {32'h459dee10, 32'h00000000} /* (7, 19, 16) {real, imag} */,
  {32'h459e113e, 32'h00000000} /* (7, 19, 15) {real, imag} */,
  {32'h459b6e91, 32'h00000000} /* (7, 19, 14) {real, imag} */,
  {32'h457f6bc9, 32'h00000000} /* (7, 19, 13) {real, imag} */,
  {32'h453599b1, 32'h00000000} /* (7, 19, 12) {real, imag} */,
  {32'h44bec544, 32'h00000000} /* (7, 19, 11) {real, imag} */,
  {32'hc4a1efbd, 32'h00000000} /* (7, 19, 10) {real, imag} */,
  {32'hc4c8f701, 32'h00000000} /* (7, 19, 9) {real, imag} */,
  {32'hc57b4400, 32'h00000000} /* (7, 19, 8) {real, imag} */,
  {32'hc5347875, 32'h00000000} /* (7, 19, 7) {real, imag} */,
  {32'hc52a5f7b, 32'h00000000} /* (7, 19, 6) {real, imag} */,
  {32'hc5532d82, 32'h00000000} /* (7, 19, 5) {real, imag} */,
  {32'hc5872b77, 32'h00000000} /* (7, 19, 4) {real, imag} */,
  {32'hc58a8be0, 32'h00000000} /* (7, 19, 3) {real, imag} */,
  {32'hc58f7671, 32'h00000000} /* (7, 19, 2) {real, imag} */,
  {32'hc58a4142, 32'h00000000} /* (7, 19, 1) {real, imag} */,
  {32'hc55892e1, 32'h00000000} /* (7, 19, 0) {real, imag} */,
  {32'hc5969668, 32'h00000000} /* (7, 18, 31) {real, imag} */,
  {32'hc5b8aebf, 32'h00000000} /* (7, 18, 30) {real, imag} */,
  {32'hc59fbece, 32'h00000000} /* (7, 18, 29) {real, imag} */,
  {32'hc5944010, 32'h00000000} /* (7, 18, 28) {real, imag} */,
  {32'hc5a4dfb4, 32'h00000000} /* (7, 18, 27) {real, imag} */,
  {32'hc59a10a3, 32'h00000000} /* (7, 18, 26) {real, imag} */,
  {32'hc594ca43, 32'h00000000} /* (7, 18, 25) {real, imag} */,
  {32'hc5a52063, 32'h00000000} /* (7, 18, 24) {real, imag} */,
  {32'hc57f9663, 32'h00000000} /* (7, 18, 23) {real, imag} */,
  {32'hc520c8de, 32'h00000000} /* (7, 18, 22) {real, imag} */,
  {32'hc3b81508, 32'h00000000} /* (7, 18, 21) {real, imag} */,
  {32'h4504b62a, 32'h00000000} /* (7, 18, 20) {real, imag} */,
  {32'h4540766e, 32'h00000000} /* (7, 18, 19) {real, imag} */,
  {32'h456befaf, 32'h00000000} /* (7, 18, 18) {real, imag} */,
  {32'h45da5c20, 32'h00000000} /* (7, 18, 17) {real, imag} */,
  {32'h45d47d1a, 32'h00000000} /* (7, 18, 16) {real, imag} */,
  {32'h45b2d7ae, 32'h00000000} /* (7, 18, 15) {real, imag} */,
  {32'h45c7f843, 32'h00000000} /* (7, 18, 14) {real, imag} */,
  {32'h459f9486, 32'h00000000} /* (7, 18, 13) {real, imag} */,
  {32'h45386d84, 32'h00000000} /* (7, 18, 12) {real, imag} */,
  {32'h4501963c, 32'h00000000} /* (7, 18, 11) {real, imag} */,
  {32'hc3c39140, 32'h00000000} /* (7, 18, 10) {real, imag} */,
  {32'hc536cfe7, 32'h00000000} /* (7, 18, 9) {real, imag} */,
  {32'hc57988fa, 32'h00000000} /* (7, 18, 8) {real, imag} */,
  {32'hc57af85d, 32'h00000000} /* (7, 18, 7) {real, imag} */,
  {32'hc595265d, 32'h00000000} /* (7, 18, 6) {real, imag} */,
  {32'hc59e5db6, 32'h00000000} /* (7, 18, 5) {real, imag} */,
  {32'hc5aefb13, 32'h00000000} /* (7, 18, 4) {real, imag} */,
  {32'hc5c320f7, 32'h00000000} /* (7, 18, 3) {real, imag} */,
  {32'hc5b2da57, 32'h00000000} /* (7, 18, 2) {real, imag} */,
  {32'hc5b50956, 32'h00000000} /* (7, 18, 1) {real, imag} */,
  {32'hc5a0f43c, 32'h00000000} /* (7, 18, 0) {real, imag} */,
  {32'hc5c73eab, 32'h00000000} /* (7, 17, 31) {real, imag} */,
  {32'hc5e9906e, 32'h00000000} /* (7, 17, 30) {real, imag} */,
  {32'hc5c72366, 32'h00000000} /* (7, 17, 29) {real, imag} */,
  {32'hc5afe08c, 32'h00000000} /* (7, 17, 28) {real, imag} */,
  {32'hc5cbc6dc, 32'h00000000} /* (7, 17, 27) {real, imag} */,
  {32'hc5afca84, 32'h00000000} /* (7, 17, 26) {real, imag} */,
  {32'hc5bf0ea9, 32'h00000000} /* (7, 17, 25) {real, imag} */,
  {32'hc5c908e8, 32'h00000000} /* (7, 17, 24) {real, imag} */,
  {32'hc58166ca, 32'h00000000} /* (7, 17, 23) {real, imag} */,
  {32'hc521b9cc, 32'h00000000} /* (7, 17, 22) {real, imag} */,
  {32'hc42a7dac, 32'h00000000} /* (7, 17, 21) {real, imag} */,
  {32'h44e7c2b8, 32'h00000000} /* (7, 17, 20) {real, imag} */,
  {32'h457090e7, 32'h00000000} /* (7, 17, 19) {real, imag} */,
  {32'h45945daa, 32'h00000000} /* (7, 17, 18) {real, imag} */,
  {32'h45b00493, 32'h00000000} /* (7, 17, 17) {real, imag} */,
  {32'h45a75934, 32'h00000000} /* (7, 17, 16) {real, imag} */,
  {32'h45d9fbd9, 32'h00000000} /* (7, 17, 15) {real, imag} */,
  {32'h45c9d276, 32'h00000000} /* (7, 17, 14) {real, imag} */,
  {32'h45915696, 32'h00000000} /* (7, 17, 13) {real, imag} */,
  {32'h4583b6e6, 32'h00000000} /* (7, 17, 12) {real, imag} */,
  {32'h44d712d2, 32'h00000000} /* (7, 17, 11) {real, imag} */,
  {32'hc49e663c, 32'h00000000} /* (7, 17, 10) {real, imag} */,
  {32'hc5354f26, 32'h00000000} /* (7, 17, 9) {real, imag} */,
  {32'hc5833968, 32'h00000000} /* (7, 17, 8) {real, imag} */,
  {32'hc5951848, 32'h00000000} /* (7, 17, 7) {real, imag} */,
  {32'hc5b986a2, 32'h00000000} /* (7, 17, 6) {real, imag} */,
  {32'hc5c1ba36, 32'h00000000} /* (7, 17, 5) {real, imag} */,
  {32'hc5d5619e, 32'h00000000} /* (7, 17, 4) {real, imag} */,
  {32'hc5f4a478, 32'h00000000} /* (7, 17, 3) {real, imag} */,
  {32'hc5dfc0cc, 32'h00000000} /* (7, 17, 2) {real, imag} */,
  {32'hc5c8a33b, 32'h00000000} /* (7, 17, 1) {real, imag} */,
  {32'hc5b742ba, 32'h00000000} /* (7, 17, 0) {real, imag} */,
  {32'hc5c0d453, 32'h00000000} /* (7, 16, 31) {real, imag} */,
  {32'hc5eab12d, 32'h00000000} /* (7, 16, 30) {real, imag} */,
  {32'hc5d59cc1, 32'h00000000} /* (7, 16, 29) {real, imag} */,
  {32'hc5dc9d54, 32'h00000000} /* (7, 16, 28) {real, imag} */,
  {32'hc5d34490, 32'h00000000} /* (7, 16, 27) {real, imag} */,
  {32'hc5badf70, 32'h00000000} /* (7, 16, 26) {real, imag} */,
  {32'hc5e11140, 32'h00000000} /* (7, 16, 25) {real, imag} */,
  {32'hc5c000e2, 32'h00000000} /* (7, 16, 24) {real, imag} */,
  {32'hc58802dd, 32'h00000000} /* (7, 16, 23) {real, imag} */,
  {32'hc55f0fea, 32'h00000000} /* (7, 16, 22) {real, imag} */,
  {32'hc30f3d40, 32'h00000000} /* (7, 16, 21) {real, imag} */,
  {32'h44fc4666, 32'h00000000} /* (7, 16, 20) {real, imag} */,
  {32'h45828a5c, 32'h00000000} /* (7, 16, 19) {real, imag} */,
  {32'h45b3b7c4, 32'h00000000} /* (7, 16, 18) {real, imag} */,
  {32'h45bed193, 32'h00000000} /* (7, 16, 17) {real, imag} */,
  {32'h45bed292, 32'h00000000} /* (7, 16, 16) {real, imag} */,
  {32'h45be2877, 32'h00000000} /* (7, 16, 15) {real, imag} */,
  {32'h45b70d35, 32'h00000000} /* (7, 16, 14) {real, imag} */,
  {32'h458b8469, 32'h00000000} /* (7, 16, 13) {real, imag} */,
  {32'h4532b2c1, 32'h00000000} /* (7, 16, 12) {real, imag} */,
  {32'h44ce5990, 32'h00000000} /* (7, 16, 11) {real, imag} */,
  {32'hc49e8aaa, 32'h00000000} /* (7, 16, 10) {real, imag} */,
  {32'hc52fa0e1, 32'h00000000} /* (7, 16, 9) {real, imag} */,
  {32'hc581d7ce, 32'h00000000} /* (7, 16, 8) {real, imag} */,
  {32'hc5a99ec1, 32'h00000000} /* (7, 16, 7) {real, imag} */,
  {32'hc5d415bd, 32'h00000000} /* (7, 16, 6) {real, imag} */,
  {32'hc5c525ee, 32'h00000000} /* (7, 16, 5) {real, imag} */,
  {32'hc5c64c82, 32'h00000000} /* (7, 16, 4) {real, imag} */,
  {32'hc5da49ee, 32'h00000000} /* (7, 16, 3) {real, imag} */,
  {32'hc5fa311c, 32'h00000000} /* (7, 16, 2) {real, imag} */,
  {32'hc5e89663, 32'h00000000} /* (7, 16, 1) {real, imag} */,
  {32'hc5c7da82, 32'h00000000} /* (7, 16, 0) {real, imag} */,
  {32'hc5c17bdc, 32'h00000000} /* (7, 15, 31) {real, imag} */,
  {32'hc5c74e7b, 32'h00000000} /* (7, 15, 30) {real, imag} */,
  {32'hc5e9353c, 32'h00000000} /* (7, 15, 29) {real, imag} */,
  {32'hc5f62d69, 32'h00000000} /* (7, 15, 28) {real, imag} */,
  {32'hc5f1df52, 32'h00000000} /* (7, 15, 27) {real, imag} */,
  {32'hc5f012ce, 32'h00000000} /* (7, 15, 26) {real, imag} */,
  {32'hc5ded1d6, 32'h00000000} /* (7, 15, 25) {real, imag} */,
  {32'hc5b64a0a, 32'h00000000} /* (7, 15, 24) {real, imag} */,
  {32'hc58dabb5, 32'h00000000} /* (7, 15, 23) {real, imag} */,
  {32'hc577025f, 32'h00000000} /* (7, 15, 22) {real, imag} */,
  {32'h42e16320, 32'h00000000} /* (7, 15, 21) {real, imag} */,
  {32'h4517bdf2, 32'h00000000} /* (7, 15, 20) {real, imag} */,
  {32'h456035bd, 32'h00000000} /* (7, 15, 19) {real, imag} */,
  {32'h45931d78, 32'h00000000} /* (7, 15, 18) {real, imag} */,
  {32'h45be4b6c, 32'h00000000} /* (7, 15, 17) {real, imag} */,
  {32'h45d0c202, 32'h00000000} /* (7, 15, 16) {real, imag} */,
  {32'h45bb5298, 32'h00000000} /* (7, 15, 15) {real, imag} */,
  {32'h45a35085, 32'h00000000} /* (7, 15, 14) {real, imag} */,
  {32'h459ddeac, 32'h00000000} /* (7, 15, 13) {real, imag} */,
  {32'h455836c2, 32'h00000000} /* (7, 15, 12) {real, imag} */,
  {32'h44788a6c, 32'h00000000} /* (7, 15, 11) {real, imag} */,
  {32'hc47da634, 32'h00000000} /* (7, 15, 10) {real, imag} */,
  {32'hc5775ae3, 32'h00000000} /* (7, 15, 9) {real, imag} */,
  {32'hc590a04e, 32'h00000000} /* (7, 15, 8) {real, imag} */,
  {32'hc5af7553, 32'h00000000} /* (7, 15, 7) {real, imag} */,
  {32'hc5c18dd4, 32'h00000000} /* (7, 15, 6) {real, imag} */,
  {32'hc5c0e3b2, 32'h00000000} /* (7, 15, 5) {real, imag} */,
  {32'hc5d84799, 32'h00000000} /* (7, 15, 4) {real, imag} */,
  {32'hc5e14cbc, 32'h00000000} /* (7, 15, 3) {real, imag} */,
  {32'hc5f742d0, 32'h00000000} /* (7, 15, 2) {real, imag} */,
  {32'hc6065737, 32'h00000000} /* (7, 15, 1) {real, imag} */,
  {32'hc5cb6382, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'hc5b066f2, 32'h00000000} /* (7, 14, 31) {real, imag} */,
  {32'hc5b5d72a, 32'h00000000} /* (7, 14, 30) {real, imag} */,
  {32'hc5bb251d, 32'h00000000} /* (7, 14, 29) {real, imag} */,
  {32'hc5d1f91a, 32'h00000000} /* (7, 14, 28) {real, imag} */,
  {32'hc5d928c9, 32'h00000000} /* (7, 14, 27) {real, imag} */,
  {32'hc5ba53ec, 32'h00000000} /* (7, 14, 26) {real, imag} */,
  {32'hc5d2245c, 32'h00000000} /* (7, 14, 25) {real, imag} */,
  {32'hc5a59805, 32'h00000000} /* (7, 14, 24) {real, imag} */,
  {32'hc58c05d7, 32'h00000000} /* (7, 14, 23) {real, imag} */,
  {32'hc51f83ec, 32'h00000000} /* (7, 14, 22) {real, imag} */,
  {32'hc4388138, 32'h00000000} /* (7, 14, 21) {real, imag} */,
  {32'h450182b6, 32'h00000000} /* (7, 14, 20) {real, imag} */,
  {32'h454188ef, 32'h00000000} /* (7, 14, 19) {real, imag} */,
  {32'h457a684c, 32'h00000000} /* (7, 14, 18) {real, imag} */,
  {32'h4590c09e, 32'h00000000} /* (7, 14, 17) {real, imag} */,
  {32'h45ab55fc, 32'h00000000} /* (7, 14, 16) {real, imag} */,
  {32'h45b95a6a, 32'h00000000} /* (7, 14, 15) {real, imag} */,
  {32'h45905a62, 32'h00000000} /* (7, 14, 14) {real, imag} */,
  {32'h45969b17, 32'h00000000} /* (7, 14, 13) {real, imag} */,
  {32'h4549027c, 32'h00000000} /* (7, 14, 12) {real, imag} */,
  {32'h444c6bf0, 32'h00000000} /* (7, 14, 11) {real, imag} */,
  {32'hc4b87f5a, 32'h00000000} /* (7, 14, 10) {real, imag} */,
  {32'hc57c1fd1, 32'h00000000} /* (7, 14, 9) {real, imag} */,
  {32'hc5ab6c13, 32'h00000000} /* (7, 14, 8) {real, imag} */,
  {32'hc5ce54f1, 32'h00000000} /* (7, 14, 7) {real, imag} */,
  {32'hc5b71172, 32'h00000000} /* (7, 14, 6) {real, imag} */,
  {32'hc5c60aad, 32'h00000000} /* (7, 14, 5) {real, imag} */,
  {32'hc5dd0c2b, 32'h00000000} /* (7, 14, 4) {real, imag} */,
  {32'hc5dca290, 32'h00000000} /* (7, 14, 3) {real, imag} */,
  {32'hc5ce2a10, 32'h00000000} /* (7, 14, 2) {real, imag} */,
  {32'hc5e44214, 32'h00000000} /* (7, 14, 1) {real, imag} */,
  {32'hc5ae0c94, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hc59026e0, 32'h00000000} /* (7, 13, 31) {real, imag} */,
  {32'hc59ff916, 32'h00000000} /* (7, 13, 30) {real, imag} */,
  {32'hc5aaafbd, 32'h00000000} /* (7, 13, 29) {real, imag} */,
  {32'hc5aa1dc8, 32'h00000000} /* (7, 13, 28) {real, imag} */,
  {32'hc5aad110, 32'h00000000} /* (7, 13, 27) {real, imag} */,
  {32'hc5a74d9e, 32'h00000000} /* (7, 13, 26) {real, imag} */,
  {32'hc59adb68, 32'h00000000} /* (7, 13, 25) {real, imag} */,
  {32'hc58dc076, 32'h00000000} /* (7, 13, 24) {real, imag} */,
  {32'hc578ccc4, 32'h00000000} /* (7, 13, 23) {real, imag} */,
  {32'hc5322c36, 32'h00000000} /* (7, 13, 22) {real, imag} */,
  {32'hc1a58d00, 32'h00000000} /* (7, 13, 21) {real, imag} */,
  {32'h44e16d32, 32'h00000000} /* (7, 13, 20) {real, imag} */,
  {32'h4558825a, 32'h00000000} /* (7, 13, 19) {real, imag} */,
  {32'h457a546e, 32'h00000000} /* (7, 13, 18) {real, imag} */,
  {32'h4576eb11, 32'h00000000} /* (7, 13, 17) {real, imag} */,
  {32'h45995297, 32'h00000000} /* (7, 13, 16) {real, imag} */,
  {32'h4591251c, 32'h00000000} /* (7, 13, 15) {real, imag} */,
  {32'h45816524, 32'h00000000} /* (7, 13, 14) {real, imag} */,
  {32'h4536c6d6, 32'h00000000} /* (7, 13, 13) {real, imag} */,
  {32'h45135957, 32'h00000000} /* (7, 13, 12) {real, imag} */,
  {32'h4489623a, 32'h00000000} /* (7, 13, 11) {real, imag} */,
  {32'hc493f28e, 32'h00000000} /* (7, 13, 10) {real, imag} */,
  {32'hc59d87c0, 32'h00000000} /* (7, 13, 9) {real, imag} */,
  {32'hc594eb68, 32'h00000000} /* (7, 13, 8) {real, imag} */,
  {32'hc586d1b2, 32'h00000000} /* (7, 13, 7) {real, imag} */,
  {32'hc5a46bde, 32'h00000000} /* (7, 13, 6) {real, imag} */,
  {32'hc5cacc23, 32'h00000000} /* (7, 13, 5) {real, imag} */,
  {32'hc5b7f212, 32'h00000000} /* (7, 13, 4) {real, imag} */,
  {32'hc5c2b13f, 32'h00000000} /* (7, 13, 3) {real, imag} */,
  {32'hc5adaee9, 32'h00000000} /* (7, 13, 2) {real, imag} */,
  {32'hc5aa0c32, 32'h00000000} /* (7, 13, 1) {real, imag} */,
  {32'hc58eb1e5, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'hc5155836, 32'h00000000} /* (7, 12, 31) {real, imag} */,
  {32'hc539378c, 32'h00000000} /* (7, 12, 30) {real, imag} */,
  {32'hc57a673a, 32'h00000000} /* (7, 12, 29) {real, imag} */,
  {32'hc59fe736, 32'h00000000} /* (7, 12, 28) {real, imag} */,
  {32'hc5894724, 32'h00000000} /* (7, 12, 27) {real, imag} */,
  {32'hc5706513, 32'h00000000} /* (7, 12, 26) {real, imag} */,
  {32'hc5944434, 32'h00000000} /* (7, 12, 25) {real, imag} */,
  {32'hc5807ea5, 32'h00000000} /* (7, 12, 24) {real, imag} */,
  {32'hc50c2311, 32'h00000000} /* (7, 12, 23) {real, imag} */,
  {32'hc437de34, 32'h00000000} /* (7, 12, 22) {real, imag} */,
  {32'h43ac8b48, 32'h00000000} /* (7, 12, 21) {real, imag} */,
  {32'h44eb9a92, 32'h00000000} /* (7, 12, 20) {real, imag} */,
  {32'h44e4fd4e, 32'h00000000} /* (7, 12, 19) {real, imag} */,
  {32'h451ef7ba, 32'h00000000} /* (7, 12, 18) {real, imag} */,
  {32'h45427af8, 32'h00000000} /* (7, 12, 17) {real, imag} */,
  {32'h4538f942, 32'h00000000} /* (7, 12, 16) {real, imag} */,
  {32'h4563770c, 32'h00000000} /* (7, 12, 15) {real, imag} */,
  {32'h4535a50c, 32'h00000000} /* (7, 12, 14) {real, imag} */,
  {32'h45282174, 32'h00000000} /* (7, 12, 13) {real, imag} */,
  {32'h4509216a, 32'h00000000} /* (7, 12, 12) {real, imag} */,
  {32'h4482f6f2, 32'h00000000} /* (7, 12, 11) {real, imag} */,
  {32'hc48cb372, 32'h00000000} /* (7, 12, 10) {real, imag} */,
  {32'hc559056f, 32'h00000000} /* (7, 12, 9) {real, imag} */,
  {32'hc54dc941, 32'h00000000} /* (7, 12, 8) {real, imag} */,
  {32'hc57dde33, 32'h00000000} /* (7, 12, 7) {real, imag} */,
  {32'hc5a9a7c8, 32'h00000000} /* (7, 12, 6) {real, imag} */,
  {32'hc5906ac8, 32'h00000000} /* (7, 12, 5) {real, imag} */,
  {32'hc5828116, 32'h00000000} /* (7, 12, 4) {real, imag} */,
  {32'hc549eabb, 32'h00000000} /* (7, 12, 3) {real, imag} */,
  {32'hc5570658, 32'h00000000} /* (7, 12, 2) {real, imag} */,
  {32'hc55edf02, 32'h00000000} /* (7, 12, 1) {real, imag} */,
  {32'hc53692ea, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'hc3c27740, 32'h00000000} /* (7, 11, 31) {real, imag} */,
  {32'hc49846d4, 32'h00000000} /* (7, 11, 30) {real, imag} */,
  {32'hc489a931, 32'h00000000} /* (7, 11, 29) {real, imag} */,
  {32'hc4903d7f, 32'h00000000} /* (7, 11, 28) {real, imag} */,
  {32'hc4ef77a3, 32'h00000000} /* (7, 11, 27) {real, imag} */,
  {32'hc4c058f7, 32'h00000000} /* (7, 11, 26) {real, imag} */,
  {32'hc50de300, 32'h00000000} /* (7, 11, 25) {real, imag} */,
  {32'hc42bcf9a, 32'h00000000} /* (7, 11, 24) {real, imag} */,
  {32'h42222ec0, 32'h00000000} /* (7, 11, 23) {real, imag} */,
  {32'h420740c0, 32'h00000000} /* (7, 11, 22) {real, imag} */,
  {32'h4423b1b2, 32'h00000000} /* (7, 11, 21) {real, imag} */,
  {32'h44ed67f8, 32'h00000000} /* (7, 11, 20) {real, imag} */,
  {32'h44d1db94, 32'h00000000} /* (7, 11, 19) {real, imag} */,
  {32'h44c223d2, 32'h00000000} /* (7, 11, 18) {real, imag} */,
  {32'h449954e8, 32'h00000000} /* (7, 11, 17) {real, imag} */,
  {32'h44f7528f, 32'h00000000} /* (7, 11, 16) {real, imag} */,
  {32'h44e8ae62, 32'h00000000} /* (7, 11, 15) {real, imag} */,
  {32'h44ef80b8, 32'h00000000} /* (7, 11, 14) {real, imag} */,
  {32'h44c4437f, 32'h00000000} /* (7, 11, 13) {real, imag} */,
  {32'h44dd6113, 32'h00000000} /* (7, 11, 12) {real, imag} */,
  {32'h44729b32, 32'h00000000} /* (7, 11, 11) {real, imag} */,
  {32'hc4eebdd9, 32'h00000000} /* (7, 11, 10) {real, imag} */,
  {32'hc4f61054, 32'h00000000} /* (7, 11, 9) {real, imag} */,
  {32'hc50a30fa, 32'h00000000} /* (7, 11, 8) {real, imag} */,
  {32'hc510b2df, 32'h00000000} /* (7, 11, 7) {real, imag} */,
  {32'hc534dfaf, 32'h00000000} /* (7, 11, 6) {real, imag} */,
  {32'hc540fc04, 32'h00000000} /* (7, 11, 5) {real, imag} */,
  {32'hc4c021f0, 32'h00000000} /* (7, 11, 4) {real, imag} */,
  {32'hc4daac58, 32'h00000000} /* (7, 11, 3) {real, imag} */,
  {32'hc4bca118, 32'h00000000} /* (7, 11, 2) {real, imag} */,
  {32'hc500ea0a, 32'h00000000} /* (7, 11, 1) {real, imag} */,
  {32'hc4b0bae7, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'h44f2f6de, 32'h00000000} /* (7, 10, 31) {real, imag} */,
  {32'h44e77e91, 32'h00000000} /* (7, 10, 30) {real, imag} */,
  {32'h44d136d3, 32'h00000000} /* (7, 10, 29) {real, imag} */,
  {32'h450892fb, 32'h00000000} /* (7, 10, 28) {real, imag} */,
  {32'h4502fa0f, 32'h00000000} /* (7, 10, 27) {real, imag} */,
  {32'h44c10b93, 32'h00000000} /* (7, 10, 26) {real, imag} */,
  {32'h44db7419, 32'h00000000} /* (7, 10, 25) {real, imag} */,
  {32'h4521732c, 32'h00000000} /* (7, 10, 24) {real, imag} */,
  {32'h45278bd8, 32'h00000000} /* (7, 10, 23) {real, imag} */,
  {32'h44f72952, 32'h00000000} /* (7, 10, 22) {real, imag} */,
  {32'h4501974f, 32'h00000000} /* (7, 10, 21) {real, imag} */,
  {32'h449b14cd, 32'h00000000} /* (7, 10, 20) {real, imag} */,
  {32'h43bafa88, 32'h00000000} /* (7, 10, 19) {real, imag} */,
  {32'h42ae1a00, 32'h00000000} /* (7, 10, 18) {real, imag} */,
  {32'hc4712b32, 32'h00000000} /* (7, 10, 17) {real, imag} */,
  {32'hc51d246d, 32'h00000000} /* (7, 10, 16) {real, imag} */,
  {32'hc49ba3dc, 32'h00000000} /* (7, 10, 15) {real, imag} */,
  {32'hc4708036, 32'h00000000} /* (7, 10, 14) {real, imag} */,
  {32'hc42b4916, 32'h00000000} /* (7, 10, 13) {real, imag} */,
  {32'hc4b86e5c, 32'h00000000} /* (7, 10, 12) {real, imag} */,
  {32'hc5057917, 32'h00000000} /* (7, 10, 11) {real, imag} */,
  {32'hc37007e8, 32'h00000000} /* (7, 10, 10) {real, imag} */,
  {32'hc372f2b8, 32'h00000000} /* (7, 10, 9) {real, imag} */,
  {32'hc20a42a0, 32'h00000000} /* (7, 10, 8) {real, imag} */,
  {32'h44568acc, 32'h00000000} /* (7, 10, 7) {real, imag} */,
  {32'h4405811c, 32'h00000000} /* (7, 10, 6) {real, imag} */,
  {32'h4472fbdd, 32'h00000000} /* (7, 10, 5) {real, imag} */,
  {32'h4419ea04, 32'h00000000} /* (7, 10, 4) {real, imag} */,
  {32'h445b9da8, 32'h00000000} /* (7, 10, 3) {real, imag} */,
  {32'h44b48cf4, 32'h00000000} /* (7, 10, 2) {real, imag} */,
  {32'h44b1a26f, 32'h00000000} /* (7, 10, 1) {real, imag} */,
  {32'h44fa94c5, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'h4595a4fd, 32'h00000000} /* (7, 9, 31) {real, imag} */,
  {32'h459a4d68, 32'h00000000} /* (7, 9, 30) {real, imag} */,
  {32'h4584fee6, 32'h00000000} /* (7, 9, 29) {real, imag} */,
  {32'h458c831a, 32'h00000000} /* (7, 9, 28) {real, imag} */,
  {32'h45895cfe, 32'h00000000} /* (7, 9, 27) {real, imag} */,
  {32'h45819167, 32'h00000000} /* (7, 9, 26) {real, imag} */,
  {32'h45ae443e, 32'h00000000} /* (7, 9, 25) {real, imag} */,
  {32'h45b25892, 32'h00000000} /* (7, 9, 24) {real, imag} */,
  {32'h45970ccb, 32'h00000000} /* (7, 9, 23) {real, imag} */,
  {32'h45a37fa4, 32'h00000000} /* (7, 9, 22) {real, imag} */,
  {32'h4584762e, 32'h00000000} /* (7, 9, 21) {real, imag} */,
  {32'h44ba6df2, 32'h00000000} /* (7, 9, 20) {real, imag} */,
  {32'h4238f500, 32'h00000000} /* (7, 9, 19) {real, imag} */,
  {32'hc4cf222e, 32'h00000000} /* (7, 9, 18) {real, imag} */,
  {32'hc533a63f, 32'h00000000} /* (7, 9, 17) {real, imag} */,
  {32'hc5525b1a, 32'h00000000} /* (7, 9, 16) {real, imag} */,
  {32'hc5329aa4, 32'h00000000} /* (7, 9, 15) {real, imag} */,
  {32'hc4fbe37a, 32'h00000000} /* (7, 9, 14) {real, imag} */,
  {32'hc5489015, 32'h00000000} /* (7, 9, 13) {real, imag} */,
  {32'hc51d0648, 32'h00000000} /* (7, 9, 12) {real, imag} */,
  {32'hc4e33122, 32'h00000000} /* (7, 9, 11) {real, imag} */,
  {32'hc414c690, 32'h00000000} /* (7, 9, 10) {real, imag} */,
  {32'h43969370, 32'h00000000} /* (7, 9, 9) {real, imag} */,
  {32'h450d9ee5, 32'h00000000} /* (7, 9, 8) {real, imag} */,
  {32'h453dd4a0, 32'h00000000} /* (7, 9, 7) {real, imag} */,
  {32'h451d696f, 32'h00000000} /* (7, 9, 6) {real, imag} */,
  {32'h4526c534, 32'h00000000} /* (7, 9, 5) {real, imag} */,
  {32'h45355693, 32'h00000000} /* (7, 9, 4) {real, imag} */,
  {32'h4578d85e, 32'h00000000} /* (7, 9, 3) {real, imag} */,
  {32'h4587691e, 32'h00000000} /* (7, 9, 2) {real, imag} */,
  {32'h45a28b10, 32'h00000000} /* (7, 9, 1) {real, imag} */,
  {32'h4587d427, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'h45b10caa, 32'h00000000} /* (7, 8, 31) {real, imag} */,
  {32'h45c670ab, 32'h00000000} /* (7, 8, 30) {real, imag} */,
  {32'h45b7e2b8, 32'h00000000} /* (7, 8, 29) {real, imag} */,
  {32'h45c90ddc, 32'h00000000} /* (7, 8, 28) {real, imag} */,
  {32'h45b46607, 32'h00000000} /* (7, 8, 27) {real, imag} */,
  {32'h45c498ae, 32'h00000000} /* (7, 8, 26) {real, imag} */,
  {32'h45c8284a, 32'h00000000} /* (7, 8, 25) {real, imag} */,
  {32'h45bbb6f9, 32'h00000000} /* (7, 8, 24) {real, imag} */,
  {32'h45da3dba, 32'h00000000} /* (7, 8, 23) {real, imag} */,
  {32'h45d6018c, 32'h00000000} /* (7, 8, 22) {real, imag} */,
  {32'h453fdbd0, 32'h00000000} /* (7, 8, 21) {real, imag} */,
  {32'h44874cd6, 32'h00000000} /* (7, 8, 20) {real, imag} */,
  {32'hc3200cd0, 32'h00000000} /* (7, 8, 19) {real, imag} */,
  {32'hc51ae02a, 32'h00000000} /* (7, 8, 18) {real, imag} */,
  {32'hc5484044, 32'h00000000} /* (7, 8, 17) {real, imag} */,
  {32'hc535c91d, 32'h00000000} /* (7, 8, 16) {real, imag} */,
  {32'hc55c8a5b, 32'h00000000} /* (7, 8, 15) {real, imag} */,
  {32'hc5687886, 32'h00000000} /* (7, 8, 14) {real, imag} */,
  {32'hc56ab960, 32'h00000000} /* (7, 8, 13) {real, imag} */,
  {32'hc53d7634, 32'h00000000} /* (7, 8, 12) {real, imag} */,
  {32'hc50846d6, 32'h00000000} /* (7, 8, 11) {real, imag} */,
  {32'hc42f5cf0, 32'h00000000} /* (7, 8, 10) {real, imag} */,
  {32'h44813116, 32'h00000000} /* (7, 8, 9) {real, imag} */,
  {32'h45167f96, 32'h00000000} /* (7, 8, 8) {real, imag} */,
  {32'h456d67cb, 32'h00000000} /* (7, 8, 7) {real, imag} */,
  {32'h453b0abc, 32'h00000000} /* (7, 8, 6) {real, imag} */,
  {32'h45818950, 32'h00000000} /* (7, 8, 5) {real, imag} */,
  {32'h45a26464, 32'h00000000} /* (7, 8, 4) {real, imag} */,
  {32'h45a2f606, 32'h00000000} /* (7, 8, 3) {real, imag} */,
  {32'h45c61c23, 32'h00000000} /* (7, 8, 2) {real, imag} */,
  {32'h45c6d9c2, 32'h00000000} /* (7, 8, 1) {real, imag} */,
  {32'h45b90198, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'h45ea96b5, 32'h00000000} /* (7, 7, 31) {real, imag} */,
  {32'h46063670, 32'h00000000} /* (7, 7, 30) {real, imag} */,
  {32'h45e6481c, 32'h00000000} /* (7, 7, 29) {real, imag} */,
  {32'h45db9014, 32'h00000000} /* (7, 7, 28) {real, imag} */,
  {32'h45ed583f, 32'h00000000} /* (7, 7, 27) {real, imag} */,
  {32'h45d6e424, 32'h00000000} /* (7, 7, 26) {real, imag} */,
  {32'h45d48e91, 32'h00000000} /* (7, 7, 25) {real, imag} */,
  {32'h460197e2, 32'h00000000} /* (7, 7, 24) {real, imag} */,
  {32'h45e9f556, 32'h00000000} /* (7, 7, 23) {real, imag} */,
  {32'h45de1538, 32'h00000000} /* (7, 7, 22) {real, imag} */,
  {32'h458a4eb1, 32'h00000000} /* (7, 7, 21) {real, imag} */,
  {32'h44ecfd7e, 32'h00000000} /* (7, 7, 20) {real, imag} */,
  {32'hc39cb320, 32'h00000000} /* (7, 7, 19) {real, imag} */,
  {32'hc4f360b2, 32'h00000000} /* (7, 7, 18) {real, imag} */,
  {32'hc5195b8a, 32'h00000000} /* (7, 7, 17) {real, imag} */,
  {32'hc58140d6, 32'h00000000} /* (7, 7, 16) {real, imag} */,
  {32'hc58e3cc7, 32'h00000000} /* (7, 7, 15) {real, imag} */,
  {32'hc5a39e37, 32'h00000000} /* (7, 7, 14) {real, imag} */,
  {32'hc58ba618, 32'h00000000} /* (7, 7, 13) {real, imag} */,
  {32'hc57f4638, 32'h00000000} /* (7, 7, 12) {real, imag} */,
  {32'hc553bb42, 32'h00000000} /* (7, 7, 11) {real, imag} */,
  {32'hc2551940, 32'h00000000} /* (7, 7, 10) {real, imag} */,
  {32'h4495951c, 32'h00000000} /* (7, 7, 9) {real, imag} */,
  {32'h45533549, 32'h00000000} /* (7, 7, 8) {real, imag} */,
  {32'h4561f341, 32'h00000000} /* (7, 7, 7) {real, imag} */,
  {32'h45800202, 32'h00000000} /* (7, 7, 6) {real, imag} */,
  {32'h4590b973, 32'h00000000} /* (7, 7, 5) {real, imag} */,
  {32'h45c3dac8, 32'h00000000} /* (7, 7, 4) {real, imag} */,
  {32'h45e5e220, 32'h00000000} /* (7, 7, 3) {real, imag} */,
  {32'h45c7a644, 32'h00000000} /* (7, 7, 2) {real, imag} */,
  {32'h45d8a72d, 32'h00000000} /* (7, 7, 1) {real, imag} */,
  {32'h45cddfc8, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'h45fa6156, 32'h00000000} /* (7, 6, 31) {real, imag} */,
  {32'h46131b88, 32'h00000000} /* (7, 6, 30) {real, imag} */,
  {32'h460a36c2, 32'h00000000} /* (7, 6, 29) {real, imag} */,
  {32'h46071179, 32'h00000000} /* (7, 6, 28) {real, imag} */,
  {32'h46108ab4, 32'h00000000} /* (7, 6, 27) {real, imag} */,
  {32'h46102587, 32'h00000000} /* (7, 6, 26) {real, imag} */,
  {32'h460797aa, 32'h00000000} /* (7, 6, 25) {real, imag} */,
  {32'h46086ebb, 32'h00000000} /* (7, 6, 24) {real, imag} */,
  {32'h45f08920, 32'h00000000} /* (7, 6, 23) {real, imag} */,
  {32'h45f96f42, 32'h00000000} /* (7, 6, 22) {real, imag} */,
  {32'h45b5ea02, 32'h00000000} /* (7, 6, 21) {real, imag} */,
  {32'h44d8f7a0, 32'h00000000} /* (7, 6, 20) {real, imag} */,
  {32'h445b13d8, 32'h00000000} /* (7, 6, 19) {real, imag} */,
  {32'h42b328c0, 32'h00000000} /* (7, 6, 18) {real, imag} */,
  {32'hc509287e, 32'h00000000} /* (7, 6, 17) {real, imag} */,
  {32'hc55c0c27, 32'h00000000} /* (7, 6, 16) {real, imag} */,
  {32'hc583ae26, 32'h00000000} /* (7, 6, 15) {real, imag} */,
  {32'hc5930169, 32'h00000000} /* (7, 6, 14) {real, imag} */,
  {32'hc59aadb2, 32'h00000000} /* (7, 6, 13) {real, imag} */,
  {32'hc58399ce, 32'h00000000} /* (7, 6, 12) {real, imag} */,
  {32'hc58a3dfc, 32'h00000000} /* (7, 6, 11) {real, imag} */,
  {32'hc4b67946, 32'h00000000} /* (7, 6, 10) {real, imag} */,
  {32'h43b90030, 32'h00000000} /* (7, 6, 9) {real, imag} */,
  {32'h4554f8e4, 32'h00000000} /* (7, 6, 8) {real, imag} */,
  {32'h45101138, 32'h00000000} /* (7, 6, 7) {real, imag} */,
  {32'h456ff2c7, 32'h00000000} /* (7, 6, 6) {real, imag} */,
  {32'h45c0c5ae, 32'h00000000} /* (7, 6, 5) {real, imag} */,
  {32'h45cfa74c, 32'h00000000} /* (7, 6, 4) {real, imag} */,
  {32'h45e7e7b1, 32'h00000000} /* (7, 6, 3) {real, imag} */,
  {32'h46051bf6, 32'h00000000} /* (7, 6, 2) {real, imag} */,
  {32'h46105796, 32'h00000000} /* (7, 6, 1) {real, imag} */,
  {32'h45fb0c52, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'h460bcf24, 32'h00000000} /* (7, 5, 31) {real, imag} */,
  {32'h46013be2, 32'h00000000} /* (7, 5, 30) {real, imag} */,
  {32'h4610e8f2, 32'h00000000} /* (7, 5, 29) {real, imag} */,
  {32'h461c4cd6, 32'h00000000} /* (7, 5, 28) {real, imag} */,
  {32'h46223376, 32'h00000000} /* (7, 5, 27) {real, imag} */,
  {32'h46112d74, 32'h00000000} /* (7, 5, 26) {real, imag} */,
  {32'h4616faee, 32'h00000000} /* (7, 5, 25) {real, imag} */,
  {32'h460c3f32, 32'h00000000} /* (7, 5, 24) {real, imag} */,
  {32'h460ad1aa, 32'h00000000} /* (7, 5, 23) {real, imag} */,
  {32'h4603a72e, 32'h00000000} /* (7, 5, 22) {real, imag} */,
  {32'h45ca3008, 32'h00000000} /* (7, 5, 21) {real, imag} */,
  {32'h4585053b, 32'h00000000} /* (7, 5, 20) {real, imag} */,
  {32'h454e32c1, 32'h00000000} /* (7, 5, 19) {real, imag} */,
  {32'h44d3f4be, 32'h00000000} /* (7, 5, 18) {real, imag} */,
  {32'h43652040, 32'h00000000} /* (7, 5, 17) {real, imag} */,
  {32'hc4c7d106, 32'h00000000} /* (7, 5, 16) {real, imag} */,
  {32'hc5846c9b, 32'h00000000} /* (7, 5, 15) {real, imag} */,
  {32'hc5afe79c, 32'h00000000} /* (7, 5, 14) {real, imag} */,
  {32'hc59ff009, 32'h00000000} /* (7, 5, 13) {real, imag} */,
  {32'hc5afe55d, 32'h00000000} /* (7, 5, 12) {real, imag} */,
  {32'hc57f0284, 32'h00000000} /* (7, 5, 11) {real, imag} */,
  {32'hc513369f, 32'h00000000} /* (7, 5, 10) {real, imag} */,
  {32'hc48eb134, 32'h00000000} /* (7, 5, 9) {real, imag} */,
  {32'h43cc33f0, 32'h00000000} /* (7, 5, 8) {real, imag} */,
  {32'h443263d0, 32'h00000000} /* (7, 5, 7) {real, imag} */,
  {32'h452f3a36, 32'h00000000} /* (7, 5, 6) {real, imag} */,
  {32'h45ac7728, 32'h00000000} /* (7, 5, 5) {real, imag} */,
  {32'h45e69eb9, 32'h00000000} /* (7, 5, 4) {real, imag} */,
  {32'h45dc0b72, 32'h00000000} /* (7, 5, 3) {real, imag} */,
  {32'h460fbea3, 32'h00000000} /* (7, 5, 2) {real, imag} */,
  {32'h461ec715, 32'h00000000} /* (7, 5, 1) {real, imag} */,
  {32'h46019c25, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'h460e66a8, 32'h00000000} /* (7, 4, 31) {real, imag} */,
  {32'h4620842a, 32'h00000000} /* (7, 4, 30) {real, imag} */,
  {32'h460e9ca2, 32'h00000000} /* (7, 4, 29) {real, imag} */,
  {32'h461a4aa0, 32'h00000000} /* (7, 4, 28) {real, imag} */,
  {32'h462242b2, 32'h00000000} /* (7, 4, 27) {real, imag} */,
  {32'h461ad0c0, 32'h00000000} /* (7, 4, 26) {real, imag} */,
  {32'h46187d0b, 32'h00000000} /* (7, 4, 25) {real, imag} */,
  {32'h46106dc4, 32'h00000000} /* (7, 4, 24) {real, imag} */,
  {32'h461cd391, 32'h00000000} /* (7, 4, 23) {real, imag} */,
  {32'h46066c45, 32'h00000000} /* (7, 4, 22) {real, imag} */,
  {32'h45fa914a, 32'h00000000} /* (7, 4, 21) {real, imag} */,
  {32'h45bcbcf3, 32'h00000000} /* (7, 4, 20) {real, imag} */,
  {32'h45997bc4, 32'h00000000} /* (7, 4, 19) {real, imag} */,
  {32'h4584ae47, 32'h00000000} /* (7, 4, 18) {real, imag} */,
  {32'h45145afc, 32'h00000000} /* (7, 4, 17) {real, imag} */,
  {32'hc36a3480, 32'h00000000} /* (7, 4, 16) {real, imag} */,
  {32'hc565d2f3, 32'h00000000} /* (7, 4, 15) {real, imag} */,
  {32'hc583de77, 32'h00000000} /* (7, 4, 14) {real, imag} */,
  {32'hc5913487, 32'h00000000} /* (7, 4, 13) {real, imag} */,
  {32'hc59fd62c, 32'h00000000} /* (7, 4, 12) {real, imag} */,
  {32'hc596e7d8, 32'h00000000} /* (7, 4, 11) {real, imag} */,
  {32'hc54e23ea, 32'h00000000} /* (7, 4, 10) {real, imag} */,
  {32'hc50369dc, 32'h00000000} /* (7, 4, 9) {real, imag} */,
  {32'hc4c06838, 32'h00000000} /* (7, 4, 8) {real, imag} */,
  {32'h443f0f30, 32'h00000000} /* (7, 4, 7) {real, imag} */,
  {32'h44d82980, 32'h00000000} /* (7, 4, 6) {real, imag} */,
  {32'h455ee603, 32'h00000000} /* (7, 4, 5) {real, imag} */,
  {32'h45b556e5, 32'h00000000} /* (7, 4, 4) {real, imag} */,
  {32'h4601c350, 32'h00000000} /* (7, 4, 3) {real, imag} */,
  {32'h46044058, 32'h00000000} /* (7, 4, 2) {real, imag} */,
  {32'h461806b7, 32'h00000000} /* (7, 4, 1) {real, imag} */,
  {32'h46119ec3, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'h4613034a, 32'h00000000} /* (7, 3, 31) {real, imag} */,
  {32'h4621bc36, 32'h00000000} /* (7, 3, 30) {real, imag} */,
  {32'h4618785a, 32'h00000000} /* (7, 3, 29) {real, imag} */,
  {32'h461adfd4, 32'h00000000} /* (7, 3, 28) {real, imag} */,
  {32'h46247d3a, 32'h00000000} /* (7, 3, 27) {real, imag} */,
  {32'h46282c16, 32'h00000000} /* (7, 3, 26) {real, imag} */,
  {32'h461a9b91, 32'h00000000} /* (7, 3, 25) {real, imag} */,
  {32'h4626528e, 32'h00000000} /* (7, 3, 24) {real, imag} */,
  {32'h4615ed50, 32'h00000000} /* (7, 3, 23) {real, imag} */,
  {32'h4603f07c, 32'h00000000} /* (7, 3, 22) {real, imag} */,
  {32'h460257bd, 32'h00000000} /* (7, 3, 21) {real, imag} */,
  {32'h45c753e0, 32'h00000000} /* (7, 3, 20) {real, imag} */,
  {32'h459f5edf, 32'h00000000} /* (7, 3, 19) {real, imag} */,
  {32'h4598e924, 32'h00000000} /* (7, 3, 18) {real, imag} */,
  {32'h451f2382, 32'h00000000} /* (7, 3, 17) {real, imag} */,
  {32'h43d54640, 32'h00000000} /* (7, 3, 16) {real, imag} */,
  {32'hc511815e, 32'h00000000} /* (7, 3, 15) {real, imag} */,
  {32'hc561df0d, 32'h00000000} /* (7, 3, 14) {real, imag} */,
  {32'hc5946494, 32'h00000000} /* (7, 3, 13) {real, imag} */,
  {32'hc5890963, 32'h00000000} /* (7, 3, 12) {real, imag} */,
  {32'hc588d96f, 32'h00000000} /* (7, 3, 11) {real, imag} */,
  {32'hc5667e6e, 32'h00000000} /* (7, 3, 10) {real, imag} */,
  {32'hc532e931, 32'h00000000} /* (7, 3, 9) {real, imag} */,
  {32'hc503cade, 32'h00000000} /* (7, 3, 8) {real, imag} */,
  {32'hc508b5a2, 32'h00000000} /* (7, 3, 7) {real, imag} */,
  {32'h43aa0450, 32'h00000000} /* (7, 3, 6) {real, imag} */,
  {32'h4578bddd, 32'h00000000} /* (7, 3, 5) {real, imag} */,
  {32'h45b88f80, 32'h00000000} /* (7, 3, 4) {real, imag} */,
  {32'h460d5740, 32'h00000000} /* (7, 3, 3) {real, imag} */,
  {32'h461a579b, 32'h00000000} /* (7, 3, 2) {real, imag} */,
  {32'h460fb464, 32'h00000000} /* (7, 3, 1) {real, imag} */,
  {32'h4613a0e6, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'h4613cc1c, 32'h00000000} /* (7, 2, 31) {real, imag} */,
  {32'h461e7cad, 32'h00000000} /* (7, 2, 30) {real, imag} */,
  {32'h462ae2a6, 32'h00000000} /* (7, 2, 29) {real, imag} */,
  {32'h4624ed18, 32'h00000000} /* (7, 2, 28) {real, imag} */,
  {32'h4623c0b3, 32'h00000000} /* (7, 2, 27) {real, imag} */,
  {32'h462d7308, 32'h00000000} /* (7, 2, 26) {real, imag} */,
  {32'h4626cc3b, 32'h00000000} /* (7, 2, 25) {real, imag} */,
  {32'h4619885a, 32'h00000000} /* (7, 2, 24) {real, imag} */,
  {32'h460fba68, 32'h00000000} /* (7, 2, 23) {real, imag} */,
  {32'h460c5c4e, 32'h00000000} /* (7, 2, 22) {real, imag} */,
  {32'h460a4c32, 32'h00000000} /* (7, 2, 21) {real, imag} */,
  {32'h45e02c12, 32'h00000000} /* (7, 2, 20) {real, imag} */,
  {32'h45b8d226, 32'h00000000} /* (7, 2, 19) {real, imag} */,
  {32'h4597ac27, 32'h00000000} /* (7, 2, 18) {real, imag} */,
  {32'h453fb12a, 32'h00000000} /* (7, 2, 17) {real, imag} */,
  {32'h446b4768, 32'h00000000} /* (7, 2, 16) {real, imag} */,
  {32'hc4b3efe6, 32'h00000000} /* (7, 2, 15) {real, imag} */,
  {32'hc54c6033, 32'h00000000} /* (7, 2, 14) {real, imag} */,
  {32'hc57b506f, 32'h00000000} /* (7, 2, 13) {real, imag} */,
  {32'hc5864d0a, 32'h00000000} /* (7, 2, 12) {real, imag} */,
  {32'hc587e6ae, 32'h00000000} /* (7, 2, 11) {real, imag} */,
  {32'hc556d6ee, 32'h00000000} /* (7, 2, 10) {real, imag} */,
  {32'hc54ec4fc, 32'h00000000} /* (7, 2, 9) {real, imag} */,
  {32'hc5145506, 32'h00000000} /* (7, 2, 8) {real, imag} */,
  {32'hc4cd41be, 32'h00000000} /* (7, 2, 7) {real, imag} */,
  {32'h43c98c20, 32'h00000000} /* (7, 2, 6) {real, imag} */,
  {32'h45506372, 32'h00000000} /* (7, 2, 5) {real, imag} */,
  {32'h45da37ce, 32'h00000000} /* (7, 2, 4) {real, imag} */,
  {32'h45fa6042, 32'h00000000} /* (7, 2, 3) {real, imag} */,
  {32'h460ec3e4, 32'h00000000} /* (7, 2, 2) {real, imag} */,
  {32'h461b5072, 32'h00000000} /* (7, 2, 1) {real, imag} */,
  {32'h461b3488, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'h460fc7cc, 32'h00000000} /* (7, 1, 31) {real, imag} */,
  {32'h461fc973, 32'h00000000} /* (7, 1, 30) {real, imag} */,
  {32'h4625935b, 32'h00000000} /* (7, 1, 29) {real, imag} */,
  {32'h462f8e6b, 32'h00000000} /* (7, 1, 28) {real, imag} */,
  {32'h4626df39, 32'h00000000} /* (7, 1, 27) {real, imag} */,
  {32'h461ff92a, 32'h00000000} /* (7, 1, 26) {real, imag} */,
  {32'h462445fc, 32'h00000000} /* (7, 1, 25) {real, imag} */,
  {32'h46148a20, 32'h00000000} /* (7, 1, 24) {real, imag} */,
  {32'h460c4a40, 32'h00000000} /* (7, 1, 23) {real, imag} */,
  {32'h45e9e7c6, 32'h00000000} /* (7, 1, 22) {real, imag} */,
  {32'h45f656b8, 32'h00000000} /* (7, 1, 21) {real, imag} */,
  {32'h45cebc0a, 32'h00000000} /* (7, 1, 20) {real, imag} */,
  {32'h459abb92, 32'h00000000} /* (7, 1, 19) {real, imag} */,
  {32'h45991c9e, 32'h00000000} /* (7, 1, 18) {real, imag} */,
  {32'h453498e5, 32'h00000000} /* (7, 1, 17) {real, imag} */,
  {32'h4454c440, 32'h00000000} /* (7, 1, 16) {real, imag} */,
  {32'hc4cf4b72, 32'h00000000} /* (7, 1, 15) {real, imag} */,
  {32'hc51c8dab, 32'h00000000} /* (7, 1, 14) {real, imag} */,
  {32'hc54befc4, 32'h00000000} /* (7, 1, 13) {real, imag} */,
  {32'hc57611b1, 32'h00000000} /* (7, 1, 12) {real, imag} */,
  {32'hc5990866, 32'h00000000} /* (7, 1, 11) {real, imag} */,
  {32'hc582071b, 32'h00000000} /* (7, 1, 10) {real, imag} */,
  {32'hc5230cab, 32'h00000000} /* (7, 1, 9) {real, imag} */,
  {32'hc50b1556, 32'h00000000} /* (7, 1, 8) {real, imag} */,
  {32'h42ae7dc0, 32'h00000000} /* (7, 1, 7) {real, imag} */,
  {32'h44e6ec7e, 32'h00000000} /* (7, 1, 6) {real, imag} */,
  {32'h453a92f8, 32'h00000000} /* (7, 1, 5) {real, imag} */,
  {32'h45cdfc1e, 32'h00000000} /* (7, 1, 4) {real, imag} */,
  {32'h46082969, 32'h00000000} /* (7, 1, 3) {real, imag} */,
  {32'h4603cf09, 32'h00000000} /* (7, 1, 2) {real, imag} */,
  {32'h4615bfe1, 32'h00000000} /* (7, 1, 1) {real, imag} */,
  {32'h46157eef, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'h4619853f, 32'h00000000} /* (7, 0, 31) {real, imag} */,
  {32'h4619a700, 32'h00000000} /* (7, 0, 30) {real, imag} */,
  {32'h46177ee2, 32'h00000000} /* (7, 0, 29) {real, imag} */,
  {32'h461a5603, 32'h00000000} /* (7, 0, 28) {real, imag} */,
  {32'h461fee8a, 32'h00000000} /* (7, 0, 27) {real, imag} */,
  {32'h46214c64, 32'h00000000} /* (7, 0, 26) {real, imag} */,
  {32'h46131fbb, 32'h00000000} /* (7, 0, 25) {real, imag} */,
  {32'h4600df8c, 32'h00000000} /* (7, 0, 24) {real, imag} */,
  {32'h45ed2574, 32'h00000000} /* (7, 0, 23) {real, imag} */,
  {32'h45d56fdc, 32'h00000000} /* (7, 0, 22) {real, imag} */,
  {32'h45ae5573, 32'h00000000} /* (7, 0, 21) {real, imag} */,
  {32'h459dd903, 32'h00000000} /* (7, 0, 20) {real, imag} */,
  {32'h456944e3, 32'h00000000} /* (7, 0, 19) {real, imag} */,
  {32'h4523d116, 32'h00000000} /* (7, 0, 18) {real, imag} */,
  {32'h44a6edfc, 32'h00000000} /* (7, 0, 17) {real, imag} */,
  {32'hc41406f8, 32'h00000000} /* (7, 0, 16) {real, imag} */,
  {32'hc4e8b200, 32'h00000000} /* (7, 0, 15) {real, imag} */,
  {32'hc565cef8, 32'h00000000} /* (7, 0, 14) {real, imag} */,
  {32'hc5601dd3, 32'h00000000} /* (7, 0, 13) {real, imag} */,
  {32'hc5852a6a, 32'h00000000} /* (7, 0, 12) {real, imag} */,
  {32'hc559b93a, 32'h00000000} /* (7, 0, 11) {real, imag} */,
  {32'hc4fac084, 32'h00000000} /* (7, 0, 10) {real, imag} */,
  {32'hc4cee548, 32'h00000000} /* (7, 0, 9) {real, imag} */,
  {32'h4397f2b8, 32'h00000000} /* (7, 0, 8) {real, imag} */,
  {32'h449e0cca, 32'h00000000} /* (7, 0, 7) {real, imag} */,
  {32'h4566c43f, 32'h00000000} /* (7, 0, 6) {real, imag} */,
  {32'h458e042b, 32'h00000000} /* (7, 0, 5) {real, imag} */,
  {32'h45b24b71, 32'h00000000} /* (7, 0, 4) {real, imag} */,
  {32'h46010931, 32'h00000000} /* (7, 0, 3) {real, imag} */,
  {32'h4601ede0, 32'h00000000} /* (7, 0, 2) {real, imag} */,
  {32'h46079f0a, 32'h00000000} /* (7, 0, 1) {real, imag} */,
  {32'h460db81e, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h45e04974, 32'h00000000} /* (6, 31, 31) {real, imag} */,
  {32'h45f880e2, 32'h00000000} /* (6, 31, 30) {real, imag} */,
  {32'h45e95f36, 32'h00000000} /* (6, 31, 29) {real, imag} */,
  {32'h45ff7760, 32'h00000000} /* (6, 31, 28) {real, imag} */,
  {32'h45e035b8, 32'h00000000} /* (6, 31, 27) {real, imag} */,
  {32'h45e3419e, 32'h00000000} /* (6, 31, 26) {real, imag} */,
  {32'h45e25624, 32'h00000000} /* (6, 31, 25) {real, imag} */,
  {32'h45ca27f7, 32'h00000000} /* (6, 31, 24) {real, imag} */,
  {32'h45b09dad, 32'h00000000} /* (6, 31, 23) {real, imag} */,
  {32'h458c1782, 32'h00000000} /* (6, 31, 22) {real, imag} */,
  {32'h45595e2e, 32'h00000000} /* (6, 31, 21) {real, imag} */,
  {32'h44fc0996, 32'h00000000} /* (6, 31, 20) {real, imag} */,
  {32'h445aa078, 32'h00000000} /* (6, 31, 19) {real, imag} */,
  {32'h438545a0, 32'h00000000} /* (6, 31, 18) {real, imag} */,
  {32'hc3fa7168, 32'h00000000} /* (6, 31, 17) {real, imag} */,
  {32'hc4bd3512, 32'h00000000} /* (6, 31, 16) {real, imag} */,
  {32'hc4c3cb88, 32'h00000000} /* (6, 31, 15) {real, imag} */,
  {32'hc50bae1c, 32'h00000000} /* (6, 31, 14) {real, imag} */,
  {32'hc4fa57d2, 32'h00000000} /* (6, 31, 13) {real, imag} */,
  {32'hc4d17b92, 32'h00000000} /* (6, 31, 12) {real, imag} */,
  {32'hc4ad2410, 32'h00000000} /* (6, 31, 11) {real, imag} */,
  {32'h43c50188, 32'h00000000} /* (6, 31, 10) {real, imag} */,
  {32'h446d8ee0, 32'h00000000} /* (6, 31, 9) {real, imag} */,
  {32'h44fe0e54, 32'h00000000} /* (6, 31, 8) {real, imag} */,
  {32'h450c0eca, 32'h00000000} /* (6, 31, 7) {real, imag} */,
  {32'h45566c64, 32'h00000000} /* (6, 31, 6) {real, imag} */,
  {32'h4585b910, 32'h00000000} /* (6, 31, 5) {real, imag} */,
  {32'h459699f8, 32'h00000000} /* (6, 31, 4) {real, imag} */,
  {32'h45c1ee25, 32'h00000000} /* (6, 31, 3) {real, imag} */,
  {32'h45c1fd24, 32'h00000000} /* (6, 31, 2) {real, imag} */,
  {32'h45e08c5a, 32'h00000000} /* (6, 31, 1) {real, imag} */,
  {32'h45eff0de, 32'h00000000} /* (6, 31, 0) {real, imag} */,
  {32'h45f78729, 32'h00000000} /* (6, 30, 31) {real, imag} */,
  {32'h460d2843, 32'h00000000} /* (6, 30, 30) {real, imag} */,
  {32'h460904a4, 32'h00000000} /* (6, 30, 29) {real, imag} */,
  {32'h4602a7f3, 32'h00000000} /* (6, 30, 28) {real, imag} */,
  {32'h45ed83f3, 32'h00000000} /* (6, 30, 27) {real, imag} */,
  {32'h45eab71d, 32'h00000000} /* (6, 30, 26) {real, imag} */,
  {32'h45d96318, 32'h00000000} /* (6, 30, 25) {real, imag} */,
  {32'h45cad0d2, 32'h00000000} /* (6, 30, 24) {real, imag} */,
  {32'h45abd164, 32'h00000000} /* (6, 30, 23) {real, imag} */,
  {32'h45add88a, 32'h00000000} /* (6, 30, 22) {real, imag} */,
  {32'h45363ce2, 32'h00000000} /* (6, 30, 21) {real, imag} */,
  {32'hc3190330, 32'h00000000} /* (6, 30, 20) {real, imag} */,
  {32'hc3bdea50, 32'h00000000} /* (6, 30, 19) {real, imag} */,
  {32'hc4725604, 32'h00000000} /* (6, 30, 18) {real, imag} */,
  {32'hc507a88f, 32'h00000000} /* (6, 30, 17) {real, imag} */,
  {32'hc505c035, 32'h00000000} /* (6, 30, 16) {real, imag} */,
  {32'hc5277c72, 32'h00000000} /* (6, 30, 15) {real, imag} */,
  {32'hc59347ba, 32'h00000000} /* (6, 30, 14) {real, imag} */,
  {32'hc527b392, 32'h00000000} /* (6, 30, 13) {real, imag} */,
  {32'hc4db2a60, 32'h00000000} /* (6, 30, 12) {real, imag} */,
  {32'hc4ab9144, 32'h00000000} /* (6, 30, 11) {real, imag} */,
  {32'h4471bad8, 32'h00000000} /* (6, 30, 10) {real, imag} */,
  {32'h44a9a590, 32'h00000000} /* (6, 30, 9) {real, imag} */,
  {32'h4513fa73, 32'h00000000} /* (6, 30, 8) {real, imag} */,
  {32'h456bd4dd, 32'h00000000} /* (6, 30, 7) {real, imag} */,
  {32'h458104ca, 32'h00000000} /* (6, 30, 6) {real, imag} */,
  {32'h45a0af87, 32'h00000000} /* (6, 30, 5) {real, imag} */,
  {32'h45b44902, 32'h00000000} /* (6, 30, 4) {real, imag} */,
  {32'h45de3741, 32'h00000000} /* (6, 30, 3) {real, imag} */,
  {32'h45ec3b28, 32'h00000000} /* (6, 30, 2) {real, imag} */,
  {32'h45fba9a6, 32'h00000000} /* (6, 30, 1) {real, imag} */,
  {32'h45ebe05a, 32'h00000000} /* (6, 30, 0) {real, imag} */,
  {32'h45f57db4, 32'h00000000} /* (6, 29, 31) {real, imag} */,
  {32'h4601e5de, 32'h00000000} /* (6, 29, 30) {real, imag} */,
  {32'h45fb5884, 32'h00000000} /* (6, 29, 29) {real, imag} */,
  {32'h45f26e30, 32'h00000000} /* (6, 29, 28) {real, imag} */,
  {32'h45ded0f6, 32'h00000000} /* (6, 29, 27) {real, imag} */,
  {32'h45d8bbfe, 32'h00000000} /* (6, 29, 26) {real, imag} */,
  {32'h45ab0b08, 32'h00000000} /* (6, 29, 25) {real, imag} */,
  {32'h45bfcb59, 32'h00000000} /* (6, 29, 24) {real, imag} */,
  {32'h45af9b5b, 32'h00000000} /* (6, 29, 23) {real, imag} */,
  {32'h4596f8b3, 32'h00000000} /* (6, 29, 22) {real, imag} */,
  {32'h45543097, 32'h00000000} /* (6, 29, 21) {real, imag} */,
  {32'h441f0e54, 32'h00000000} /* (6, 29, 20) {real, imag} */,
  {32'hc399d600, 32'h00000000} /* (6, 29, 19) {real, imag} */,
  {32'hc4c63706, 32'h00000000} /* (6, 29, 18) {real, imag} */,
  {32'hc4f25f74, 32'h00000000} /* (6, 29, 17) {real, imag} */,
  {32'hc50ac5f2, 32'h00000000} /* (6, 29, 16) {real, imag} */,
  {32'hc51d1a78, 32'h00000000} /* (6, 29, 15) {real, imag} */,
  {32'hc543b1ca, 32'h00000000} /* (6, 29, 14) {real, imag} */,
  {32'hc53c4dd9, 32'h00000000} /* (6, 29, 13) {real, imag} */,
  {32'hc4c2d5ee, 32'h00000000} /* (6, 29, 12) {real, imag} */,
  {32'hc44899c0, 32'h00000000} /* (6, 29, 11) {real, imag} */,
  {32'h4499ddb2, 32'h00000000} /* (6, 29, 10) {real, imag} */,
  {32'h454bbde1, 32'h00000000} /* (6, 29, 9) {real, imag} */,
  {32'h458f83c5, 32'h00000000} /* (6, 29, 8) {real, imag} */,
  {32'h45982d6f, 32'h00000000} /* (6, 29, 7) {real, imag} */,
  {32'h45afc35f, 32'h00000000} /* (6, 29, 6) {real, imag} */,
  {32'h45b664a0, 32'h00000000} /* (6, 29, 5) {real, imag} */,
  {32'h45d492fe, 32'h00000000} /* (6, 29, 4) {real, imag} */,
  {32'h45be05bc, 32'h00000000} /* (6, 29, 3) {real, imag} */,
  {32'h45c9ea60, 32'h00000000} /* (6, 29, 2) {real, imag} */,
  {32'h45f262ef, 32'h00000000} /* (6, 29, 1) {real, imag} */,
  {32'h45e49381, 32'h00000000} /* (6, 29, 0) {real, imag} */,
  {32'h45d8e7ae, 32'h00000000} /* (6, 28, 31) {real, imag} */,
  {32'h45ed8096, 32'h00000000} /* (6, 28, 30) {real, imag} */,
  {32'h45e6141a, 32'h00000000} /* (6, 28, 29) {real, imag} */,
  {32'h45de9b85, 32'h00000000} /* (6, 28, 28) {real, imag} */,
  {32'h45d8c814, 32'h00000000} /* (6, 28, 27) {real, imag} */,
  {32'h45badc58, 32'h00000000} /* (6, 28, 26) {real, imag} */,
  {32'h45ad5341, 32'h00000000} /* (6, 28, 25) {real, imag} */,
  {32'h45bbcb95, 32'h00000000} /* (6, 28, 24) {real, imag} */,
  {32'h45ad7994, 32'h00000000} /* (6, 28, 23) {real, imag} */,
  {32'h458d8f47, 32'h00000000} /* (6, 28, 22) {real, imag} */,
  {32'h45559c33, 32'h00000000} /* (6, 28, 21) {real, imag} */,
  {32'hc29a8120, 32'h00000000} /* (6, 28, 20) {real, imag} */,
  {32'hc448319c, 32'h00000000} /* (6, 28, 19) {real, imag} */,
  {32'hc4f56e54, 32'h00000000} /* (6, 28, 18) {real, imag} */,
  {32'hc5238894, 32'h00000000} /* (6, 28, 17) {real, imag} */,
  {32'hc510865c, 32'h00000000} /* (6, 28, 16) {real, imag} */,
  {32'hc5338ec0, 32'h00000000} /* (6, 28, 15) {real, imag} */,
  {32'hc553a571, 32'h00000000} /* (6, 28, 14) {real, imag} */,
  {32'hc51fba75, 32'h00000000} /* (6, 28, 13) {real, imag} */,
  {32'hc4c6098c, 32'h00000000} /* (6, 28, 12) {real, imag} */,
  {32'hc44c6c74, 32'h00000000} /* (6, 28, 11) {real, imag} */,
  {32'h45216cec, 32'h00000000} /* (6, 28, 10) {real, imag} */,
  {32'h4582ba25, 32'h00000000} /* (6, 28, 9) {real, imag} */,
  {32'h45972a65, 32'h00000000} /* (6, 28, 8) {real, imag} */,
  {32'h45a24ca0, 32'h00000000} /* (6, 28, 7) {real, imag} */,
  {32'h45af8461, 32'h00000000} /* (6, 28, 6) {real, imag} */,
  {32'h45d25a96, 32'h00000000} /* (6, 28, 5) {real, imag} */,
  {32'h45d83970, 32'h00000000} /* (6, 28, 4) {real, imag} */,
  {32'h45f6b388, 32'h00000000} /* (6, 28, 3) {real, imag} */,
  {32'h45e76b03, 32'h00000000} /* (6, 28, 2) {real, imag} */,
  {32'h45cf0820, 32'h00000000} /* (6, 28, 1) {real, imag} */,
  {32'h45d4355e, 32'h00000000} /* (6, 28, 0) {real, imag} */,
  {32'h45d4959c, 32'h00000000} /* (6, 27, 31) {real, imag} */,
  {32'h45dae40c, 32'h00000000} /* (6, 27, 30) {real, imag} */,
  {32'h45d49150, 32'h00000000} /* (6, 27, 29) {real, imag} */,
  {32'h45d72fb6, 32'h00000000} /* (6, 27, 28) {real, imag} */,
  {32'h45cd712d, 32'h00000000} /* (6, 27, 27) {real, imag} */,
  {32'h45c4b48e, 32'h00000000} /* (6, 27, 26) {real, imag} */,
  {32'h45ad08c4, 32'h00000000} /* (6, 27, 25) {real, imag} */,
  {32'h45c96497, 32'h00000000} /* (6, 27, 24) {real, imag} */,
  {32'h45b1341c, 32'h00000000} /* (6, 27, 23) {real, imag} */,
  {32'h45a0b63d, 32'h00000000} /* (6, 27, 22) {real, imag} */,
  {32'h4548014e, 32'h00000000} /* (6, 27, 21) {real, imag} */,
  {32'hc2e04980, 32'h00000000} /* (6, 27, 20) {real, imag} */,
  {32'hc4944f12, 32'h00000000} /* (6, 27, 19) {real, imag} */,
  {32'hc5291a01, 32'h00000000} /* (6, 27, 18) {real, imag} */,
  {32'hc5188d83, 32'h00000000} /* (6, 27, 17) {real, imag} */,
  {32'hc539b470, 32'h00000000} /* (6, 27, 16) {real, imag} */,
  {32'hc534e0f8, 32'h00000000} /* (6, 27, 15) {real, imag} */,
  {32'hc52f0ebc, 32'h00000000} /* (6, 27, 14) {real, imag} */,
  {32'hc54b1654, 32'h00000000} /* (6, 27, 13) {real, imag} */,
  {32'hc4ec1140, 32'h00000000} /* (6, 27, 12) {real, imag} */,
  {32'hc3ce8b70, 32'h00000000} /* (6, 27, 11) {real, imag} */,
  {32'h450aa72b, 32'h00000000} /* (6, 27, 10) {real, imag} */,
  {32'h4514929f, 32'h00000000} /* (6, 27, 9) {real, imag} */,
  {32'h458fc0c9, 32'h00000000} /* (6, 27, 8) {real, imag} */,
  {32'h45a745e0, 32'h00000000} /* (6, 27, 7) {real, imag} */,
  {32'h45b90eb7, 32'h00000000} /* (6, 27, 6) {real, imag} */,
  {32'h45cded9b, 32'h00000000} /* (6, 27, 5) {real, imag} */,
  {32'h45c4f712, 32'h00000000} /* (6, 27, 4) {real, imag} */,
  {32'h45d8c282, 32'h00000000} /* (6, 27, 3) {real, imag} */,
  {32'h45d0ceb4, 32'h00000000} /* (6, 27, 2) {real, imag} */,
  {32'h45d78b8e, 32'h00000000} /* (6, 27, 1) {real, imag} */,
  {32'h45d3bc26, 32'h00000000} /* (6, 27, 0) {real, imag} */,
  {32'h45c54f09, 32'h00000000} /* (6, 26, 31) {real, imag} */,
  {32'h45bf93bc, 32'h00000000} /* (6, 26, 30) {real, imag} */,
  {32'h45dfe8bf, 32'h00000000} /* (6, 26, 29) {real, imag} */,
  {32'h45d242d4, 32'h00000000} /* (6, 26, 28) {real, imag} */,
  {32'h45c8c6aa, 32'h00000000} /* (6, 26, 27) {real, imag} */,
  {32'h45c74499, 32'h00000000} /* (6, 26, 26) {real, imag} */,
  {32'h45a6bdb3, 32'h00000000} /* (6, 26, 25) {real, imag} */,
  {32'h459d4970, 32'h00000000} /* (6, 26, 24) {real, imag} */,
  {32'h45879715, 32'h00000000} /* (6, 26, 23) {real, imag} */,
  {32'h45791627, 32'h00000000} /* (6, 26, 22) {real, imag} */,
  {32'h45243412, 32'h00000000} /* (6, 26, 21) {real, imag} */,
  {32'hc11dad00, 32'h00000000} /* (6, 26, 20) {real, imag} */,
  {32'hc4a1e946, 32'h00000000} /* (6, 26, 19) {real, imag} */,
  {32'hc523927c, 32'h00000000} /* (6, 26, 18) {real, imag} */,
  {32'hc531447d, 32'h00000000} /* (6, 26, 17) {real, imag} */,
  {32'hc51c69f1, 32'h00000000} /* (6, 26, 16) {real, imag} */,
  {32'hc51cbb72, 32'h00000000} /* (6, 26, 15) {real, imag} */,
  {32'hc53a31f9, 32'h00000000} /* (6, 26, 14) {real, imag} */,
  {32'hc553faf2, 32'h00000000} /* (6, 26, 13) {real, imag} */,
  {32'hc4ab0542, 32'h00000000} /* (6, 26, 12) {real, imag} */,
  {32'hc4196570, 32'h00000000} /* (6, 26, 11) {real, imag} */,
  {32'h4509298e, 32'h00000000} /* (6, 26, 10) {real, imag} */,
  {32'h458143c1, 32'h00000000} /* (6, 26, 9) {real, imag} */,
  {32'h458ef2ec, 32'h00000000} /* (6, 26, 8) {real, imag} */,
  {32'h45a4013f, 32'h00000000} /* (6, 26, 7) {real, imag} */,
  {32'h45b1eff4, 32'h00000000} /* (6, 26, 6) {real, imag} */,
  {32'h45c4e9bd, 32'h00000000} /* (6, 26, 5) {real, imag} */,
  {32'h45bfea5c, 32'h00000000} /* (6, 26, 4) {real, imag} */,
  {32'h45ac4152, 32'h00000000} /* (6, 26, 3) {real, imag} */,
  {32'h45b0d0be, 32'h00000000} /* (6, 26, 2) {real, imag} */,
  {32'h45c92e28, 32'h00000000} /* (6, 26, 1) {real, imag} */,
  {32'h45b67866, 32'h00000000} /* (6, 26, 0) {real, imag} */,
  {32'h45b5ec05, 32'h00000000} /* (6, 25, 31) {real, imag} */,
  {32'h45d03a84, 32'h00000000} /* (6, 25, 30) {real, imag} */,
  {32'h45b764c0, 32'h00000000} /* (6, 25, 29) {real, imag} */,
  {32'h45b59cf8, 32'h00000000} /* (6, 25, 28) {real, imag} */,
  {32'h45b3a0b2, 32'h00000000} /* (6, 25, 27) {real, imag} */,
  {32'h45cf2e30, 32'h00000000} /* (6, 25, 26) {real, imag} */,
  {32'h45a6ce43, 32'h00000000} /* (6, 25, 25) {real, imag} */,
  {32'h45926ca7, 32'h00000000} /* (6, 25, 24) {real, imag} */,
  {32'h45734743, 32'h00000000} /* (6, 25, 23) {real, imag} */,
  {32'h45564808, 32'h00000000} /* (6, 25, 22) {real, imag} */,
  {32'h4519856f, 32'h00000000} /* (6, 25, 21) {real, imag} */,
  {32'h4384c1f0, 32'h00000000} /* (6, 25, 20) {real, imag} */,
  {32'hc41f1e7c, 32'h00000000} /* (6, 25, 19) {real, imag} */,
  {32'hc5017f30, 32'h00000000} /* (6, 25, 18) {real, imag} */,
  {32'hc5533242, 32'h00000000} /* (6, 25, 17) {real, imag} */,
  {32'hc51a5600, 32'h00000000} /* (6, 25, 16) {real, imag} */,
  {32'hc53e0016, 32'h00000000} /* (6, 25, 15) {real, imag} */,
  {32'hc5202cb4, 32'h00000000} /* (6, 25, 14) {real, imag} */,
  {32'hc50aabd7, 32'h00000000} /* (6, 25, 13) {real, imag} */,
  {32'hc5027b07, 32'h00000000} /* (6, 25, 12) {real, imag} */,
  {32'h3f385000, 32'h00000000} /* (6, 25, 11) {real, imag} */,
  {32'h4514c674, 32'h00000000} /* (6, 25, 10) {real, imag} */,
  {32'h4579f336, 32'h00000000} /* (6, 25, 9) {real, imag} */,
  {32'h4567c1f1, 32'h00000000} /* (6, 25, 8) {real, imag} */,
  {32'h4593bcac, 32'h00000000} /* (6, 25, 7) {real, imag} */,
  {32'h45a02b68, 32'h00000000} /* (6, 25, 6) {real, imag} */,
  {32'h45b8e71c, 32'h00000000} /* (6, 25, 5) {real, imag} */,
  {32'h45a3a7b9, 32'h00000000} /* (6, 25, 4) {real, imag} */,
  {32'h45a902f8, 32'h00000000} /* (6, 25, 3) {real, imag} */,
  {32'h45b5f794, 32'h00000000} /* (6, 25, 2) {real, imag} */,
  {32'h45bcf067, 32'h00000000} /* (6, 25, 1) {real, imag} */,
  {32'h459ed288, 32'h00000000} /* (6, 25, 0) {real, imag} */,
  {32'h4592707c, 32'h00000000} /* (6, 24, 31) {real, imag} */,
  {32'h45b129bd, 32'h00000000} /* (6, 24, 30) {real, imag} */,
  {32'h45a55328, 32'h00000000} /* (6, 24, 29) {real, imag} */,
  {32'h45b182d9, 32'h00000000} /* (6, 24, 28) {real, imag} */,
  {32'h45b5c53c, 32'h00000000} /* (6, 24, 27) {real, imag} */,
  {32'h45a445ef, 32'h00000000} /* (6, 24, 26) {real, imag} */,
  {32'h45959568, 32'h00000000} /* (6, 24, 25) {real, imag} */,
  {32'h45945909, 32'h00000000} /* (6, 24, 24) {real, imag} */,
  {32'h4585fc3a, 32'h00000000} /* (6, 24, 23) {real, imag} */,
  {32'h453cccb2, 32'h00000000} /* (6, 24, 22) {real, imag} */,
  {32'h45239753, 32'h00000000} /* (6, 24, 21) {real, imag} */,
  {32'h43dcea58, 32'h00000000} /* (6, 24, 20) {real, imag} */,
  {32'hc48b1fee, 32'h00000000} /* (6, 24, 19) {real, imag} */,
  {32'hc4428c70, 32'h00000000} /* (6, 24, 18) {real, imag} */,
  {32'hc51e47fe, 32'h00000000} /* (6, 24, 17) {real, imag} */,
  {32'hc5394a4c, 32'h00000000} /* (6, 24, 16) {real, imag} */,
  {32'hc505a53c, 32'h00000000} /* (6, 24, 15) {real, imag} */,
  {32'hc513d160, 32'h00000000} /* (6, 24, 14) {real, imag} */,
  {32'hc4adcab6, 32'h00000000} /* (6, 24, 13) {real, imag} */,
  {32'hc49f7018, 32'h00000000} /* (6, 24, 12) {real, imag} */,
  {32'hc3bd8750, 32'h00000000} /* (6, 24, 11) {real, imag} */,
  {32'h4523b1a2, 32'h00000000} /* (6, 24, 10) {real, imag} */,
  {32'h452be630, 32'h00000000} /* (6, 24, 9) {real, imag} */,
  {32'h4572276f, 32'h00000000} /* (6, 24, 8) {real, imag} */,
  {32'h457aff88, 32'h00000000} /* (6, 24, 7) {real, imag} */,
  {32'h45824f37, 32'h00000000} /* (6, 24, 6) {real, imag} */,
  {32'h45b71ffe, 32'h00000000} /* (6, 24, 5) {real, imag} */,
  {32'h4596ab18, 32'h00000000} /* (6, 24, 4) {real, imag} */,
  {32'h45991704, 32'h00000000} /* (6, 24, 3) {real, imag} */,
  {32'h45a96c14, 32'h00000000} /* (6, 24, 2) {real, imag} */,
  {32'h45917b32, 32'h00000000} /* (6, 24, 1) {real, imag} */,
  {32'h45975a12, 32'h00000000} /* (6, 24, 0) {real, imag} */,
  {32'h4588d0fc, 32'h00000000} /* (6, 23, 31) {real, imag} */,
  {32'h459fcc0b, 32'h00000000} /* (6, 23, 30) {real, imag} */,
  {32'h45911f84, 32'h00000000} /* (6, 23, 29) {real, imag} */,
  {32'h45814032, 32'h00000000} /* (6, 23, 28) {real, imag} */,
  {32'h4599d6a0, 32'h00000000} /* (6, 23, 27) {real, imag} */,
  {32'h45989ce6, 32'h00000000} /* (6, 23, 26) {real, imag} */,
  {32'h458de049, 32'h00000000} /* (6, 23, 25) {real, imag} */,
  {32'h457f3a86, 32'h00000000} /* (6, 23, 24) {real, imag} */,
  {32'h4564a8f3, 32'h00000000} /* (6, 23, 23) {real, imag} */,
  {32'h45523d48, 32'h00000000} /* (6, 23, 22) {real, imag} */,
  {32'h450db30a, 32'h00000000} /* (6, 23, 21) {real, imag} */,
  {32'h445c1d14, 32'h00000000} /* (6, 23, 20) {real, imag} */,
  {32'hc290e350, 32'h00000000} /* (6, 23, 19) {real, imag} */,
  {32'hc3c2920c, 32'h00000000} /* (6, 23, 18) {real, imag} */,
  {32'hc4c8b3e6, 32'h00000000} /* (6, 23, 17) {real, imag} */,
  {32'hc507b008, 32'h00000000} /* (6, 23, 16) {real, imag} */,
  {32'hc48be75a, 32'h00000000} /* (6, 23, 15) {real, imag} */,
  {32'hc4fe80c5, 32'h00000000} /* (6, 23, 14) {real, imag} */,
  {32'hc4bb6276, 32'h00000000} /* (6, 23, 13) {real, imag} */,
  {32'hc4641f68, 32'h00000000} /* (6, 23, 12) {real, imag} */,
  {32'h43cc9740, 32'h00000000} /* (6, 23, 11) {real, imag} */,
  {32'h44d1305c, 32'h00000000} /* (6, 23, 10) {real, imag} */,
  {32'h45039220, 32'h00000000} /* (6, 23, 9) {real, imag} */,
  {32'h45648772, 32'h00000000} /* (6, 23, 8) {real, imag} */,
  {32'h454e3e4d, 32'h00000000} /* (6, 23, 7) {real, imag} */,
  {32'h45561ac8, 32'h00000000} /* (6, 23, 6) {real, imag} */,
  {32'h45535630, 32'h00000000} /* (6, 23, 5) {real, imag} */,
  {32'h457bc56d, 32'h00000000} /* (6, 23, 4) {real, imag} */,
  {32'h455a476e, 32'h00000000} /* (6, 23, 3) {real, imag} */,
  {32'h455ef16c, 32'h00000000} /* (6, 23, 2) {real, imag} */,
  {32'h45596271, 32'h00000000} /* (6, 23, 1) {real, imag} */,
  {32'h455c542e, 32'h00000000} /* (6, 23, 0) {real, imag} */,
  {32'h452d3f31, 32'h00000000} /* (6, 22, 31) {real, imag} */,
  {32'h45337060, 32'h00000000} /* (6, 22, 30) {real, imag} */,
  {32'h453af758, 32'h00000000} /* (6, 22, 29) {real, imag} */,
  {32'h4575b192, 32'h00000000} /* (6, 22, 28) {real, imag} */,
  {32'h4587f6a5, 32'h00000000} /* (6, 22, 27) {real, imag} */,
  {32'h458cfdf5, 32'h00000000} /* (6, 22, 26) {real, imag} */,
  {32'h455d27d4, 32'h00000000} /* (6, 22, 25) {real, imag} */,
  {32'h453cfc34, 32'h00000000} /* (6, 22, 24) {real, imag} */,
  {32'h45807478, 32'h00000000} /* (6, 22, 23) {real, imag} */,
  {32'h453ba361, 32'h00000000} /* (6, 22, 22) {real, imag} */,
  {32'h44fcde82, 32'h00000000} /* (6, 22, 21) {real, imag} */,
  {32'h43f2ba86, 32'h00000000} /* (6, 22, 20) {real, imag} */,
  {32'h439fd114, 32'h00000000} /* (6, 22, 19) {real, imag} */,
  {32'hc398a148, 32'h00000000} /* (6, 22, 18) {real, imag} */,
  {32'hc4882e31, 32'h00000000} /* (6, 22, 17) {real, imag} */,
  {32'hc40dc7ae, 32'h00000000} /* (6, 22, 16) {real, imag} */,
  {32'hc4b000ee, 32'h00000000} /* (6, 22, 15) {real, imag} */,
  {32'hc4af2dab, 32'h00000000} /* (6, 22, 14) {real, imag} */,
  {32'hc45b21da, 32'h00000000} /* (6, 22, 13) {real, imag} */,
  {32'hc491ff60, 32'h00000000} /* (6, 22, 12) {real, imag} */,
  {32'hc401dd3a, 32'h00000000} /* (6, 22, 11) {real, imag} */,
  {32'h44c107dc, 32'h00000000} /* (6, 22, 10) {real, imag} */,
  {32'h4545c7b8, 32'h00000000} /* (6, 22, 9) {real, imag} */,
  {32'h454a9014, 32'h00000000} /* (6, 22, 8) {real, imag} */,
  {32'h453addb5, 32'h00000000} /* (6, 22, 7) {real, imag} */,
  {32'h455f7767, 32'h00000000} /* (6, 22, 6) {real, imag} */,
  {32'h4537ee27, 32'h00000000} /* (6, 22, 5) {real, imag} */,
  {32'h44f30726, 32'h00000000} /* (6, 22, 4) {real, imag} */,
  {32'h4514db22, 32'h00000000} /* (6, 22, 3) {real, imag} */,
  {32'h45030e81, 32'h00000000} /* (6, 22, 2) {real, imag} */,
  {32'h4518f5d2, 32'h00000000} /* (6, 22, 1) {real, imag} */,
  {32'h450f9968, 32'h00000000} /* (6, 22, 0) {real, imag} */,
  {32'h440f0186, 32'h00000000} /* (6, 21, 31) {real, imag} */,
  {32'h44c22f92, 32'h00000000} /* (6, 21, 30) {real, imag} */,
  {32'h450ade89, 32'h00000000} /* (6, 21, 29) {real, imag} */,
  {32'h454e1bfa, 32'h00000000} /* (6, 21, 28) {real, imag} */,
  {32'h455b10a8, 32'h00000000} /* (6, 21, 27) {real, imag} */,
  {32'h45012a4a, 32'h00000000} /* (6, 21, 26) {real, imag} */,
  {32'h4535d3e2, 32'h00000000} /* (6, 21, 25) {real, imag} */,
  {32'h44ec925c, 32'h00000000} /* (6, 21, 24) {real, imag} */,
  {32'h44ab2677, 32'h00000000} /* (6, 21, 23) {real, imag} */,
  {32'h449cea4e, 32'h00000000} /* (6, 21, 22) {real, imag} */,
  {32'h44677389, 32'h00000000} /* (6, 21, 21) {real, imag} */,
  {32'h43cebce8, 32'h00000000} /* (6, 21, 20) {real, imag} */,
  {32'h44935b08, 32'h00000000} /* (6, 21, 19) {real, imag} */,
  {32'h4497364a, 32'h00000000} /* (6, 21, 18) {real, imag} */,
  {32'h43472eb4, 32'h00000000} /* (6, 21, 17) {real, imag} */,
  {32'hc28911a0, 32'h00000000} /* (6, 21, 16) {real, imag} */,
  {32'h41526da0, 32'h00000000} /* (6, 21, 15) {real, imag} */,
  {32'h43e43252, 32'h00000000} /* (6, 21, 14) {real, imag} */,
  {32'h426504c0, 32'h00000000} /* (6, 21, 13) {real, imag} */,
  {32'h43f502bc, 32'h00000000} /* (6, 21, 12) {real, imag} */,
  {32'h43a3c264, 32'h00000000} /* (6, 21, 11) {real, imag} */,
  {32'h44d63cfc, 32'h00000000} /* (6, 21, 10) {real, imag} */,
  {32'h44920a9d, 32'h00000000} /* (6, 21, 9) {real, imag} */,
  {32'h451b58b4, 32'h00000000} /* (6, 21, 8) {real, imag} */,
  {32'h44d095ab, 32'h00000000} /* (6, 21, 7) {real, imag} */,
  {32'h4522671c, 32'h00000000} /* (6, 21, 6) {real, imag} */,
  {32'h44a8ad34, 32'h00000000} /* (6, 21, 5) {real, imag} */,
  {32'h442faf90, 32'h00000000} /* (6, 21, 4) {real, imag} */,
  {32'h440c8dcb, 32'h00000000} /* (6, 21, 3) {real, imag} */,
  {32'h44514d65, 32'h00000000} /* (6, 21, 2) {real, imag} */,
  {32'h4495ccc0, 32'h00000000} /* (6, 21, 1) {real, imag} */,
  {32'h4451b772, 32'h00000000} /* (6, 21, 0) {real, imag} */,
  {32'hc442ba52, 32'h00000000} /* (6, 20, 31) {real, imag} */,
  {32'hc2ca0ec0, 32'h00000000} /* (6, 20, 30) {real, imag} */,
  {32'hc2670f80, 32'h00000000} /* (6, 20, 29) {real, imag} */,
  {32'h43e46760, 32'h00000000} /* (6, 20, 28) {real, imag} */,
  {32'h43219f78, 32'h00000000} /* (6, 20, 27) {real, imag} */,
  {32'h42f5d854, 32'h00000000} /* (6, 20, 26) {real, imag} */,
  {32'hc491fa4c, 32'h00000000} /* (6, 20, 25) {real, imag} */,
  {32'hc3a7e6a3, 32'h00000000} /* (6, 20, 24) {real, imag} */,
  {32'hc447ecb6, 32'h00000000} /* (6, 20, 23) {real, imag} */,
  {32'hc391af04, 32'h00000000} /* (6, 20, 22) {real, imag} */,
  {32'h43d00a63, 32'h00000000} /* (6, 20, 21) {real, imag} */,
  {32'h44c518ee, 32'h00000000} /* (6, 20, 20) {real, imag} */,
  {32'h4505c7f1, 32'h00000000} /* (6, 20, 19) {real, imag} */,
  {32'h451e3c46, 32'h00000000} /* (6, 20, 18) {real, imag} */,
  {32'h4519460e, 32'h00000000} /* (6, 20, 17) {real, imag} */,
  {32'h450da9b0, 32'h00000000} /* (6, 20, 16) {real, imag} */,
  {32'h4511830a, 32'h00000000} /* (6, 20, 15) {real, imag} */,
  {32'h4519a20a, 32'h00000000} /* (6, 20, 14) {real, imag} */,
  {32'h44f1d44e, 32'h00000000} /* (6, 20, 13) {real, imag} */,
  {32'h44c33295, 32'h00000000} /* (6, 20, 12) {real, imag} */,
  {32'h44727922, 32'h00000000} /* (6, 20, 11) {real, imag} */,
  {32'hc46674ba, 32'h00000000} /* (6, 20, 10) {real, imag} */,
  {32'hc3fb951a, 32'h00000000} /* (6, 20, 9) {real, imag} */,
  {32'hc3c63b3b, 32'h00000000} /* (6, 20, 8) {real, imag} */,
  {32'hc482c647, 32'h00000000} /* (6, 20, 7) {real, imag} */,
  {32'hc441898a, 32'h00000000} /* (6, 20, 6) {real, imag} */,
  {32'hc410bb2a, 32'h00000000} /* (6, 20, 5) {real, imag} */,
  {32'hc4ad8570, 32'h00000000} /* (6, 20, 4) {real, imag} */,
  {32'hc4febb2f, 32'h00000000} /* (6, 20, 3) {real, imag} */,
  {32'hc48e7e7d, 32'h00000000} /* (6, 20, 2) {real, imag} */,
  {32'hc4d27a73, 32'h00000000} /* (6, 20, 1) {real, imag} */,
  {32'hc458da26, 32'h00000000} /* (6, 20, 0) {real, imag} */,
  {32'hc4dd9638, 32'h00000000} /* (6, 19, 31) {real, imag} */,
  {32'hc4d06a88, 32'h00000000} /* (6, 19, 30) {real, imag} */,
  {32'hc4fcb124, 32'h00000000} /* (6, 19, 29) {real, imag} */,
  {32'hc4c31e62, 32'h00000000} /* (6, 19, 28) {real, imag} */,
  {32'hc4e95b7f, 32'h00000000} /* (6, 19, 27) {real, imag} */,
  {32'hc50cbcbc, 32'h00000000} /* (6, 19, 26) {real, imag} */,
  {32'hc53a933a, 32'h00000000} /* (6, 19, 25) {real, imag} */,
  {32'hc53aa898, 32'h00000000} /* (6, 19, 24) {real, imag} */,
  {32'hc5164d14, 32'h00000000} /* (6, 19, 23) {real, imag} */,
  {32'hc4d60c64, 32'h00000000} /* (6, 19, 22) {real, imag} */,
  {32'h42151760, 32'h00000000} /* (6, 19, 21) {real, imag} */,
  {32'h44df8bf4, 32'h00000000} /* (6, 19, 20) {real, imag} */,
  {32'h4528608e, 32'h00000000} /* (6, 19, 19) {real, imag} */,
  {32'h455ac0f6, 32'h00000000} /* (6, 19, 18) {real, imag} */,
  {32'h457fa20d, 32'h00000000} /* (6, 19, 17) {real, imag} */,
  {32'h4554a48e, 32'h00000000} /* (6, 19, 16) {real, imag} */,
  {32'h454cff4e, 32'h00000000} /* (6, 19, 15) {real, imag} */,
  {32'h45419400, 32'h00000000} /* (6, 19, 14) {real, imag} */,
  {32'h451c414c, 32'h00000000} /* (6, 19, 13) {real, imag} */,
  {32'h4522bc21, 32'h00000000} /* (6, 19, 12) {real, imag} */,
  {32'h43882d24, 32'h00000000} /* (6, 19, 11) {real, imag} */,
  {32'hc4539969, 32'h00000000} /* (6, 19, 10) {real, imag} */,
  {32'hc20a0400, 32'h00000000} /* (6, 19, 9) {real, imag} */,
  {32'hc464bf2a, 32'h00000000} /* (6, 19, 8) {real, imag} */,
  {32'hc48b23d1, 32'h00000000} /* (6, 19, 7) {real, imag} */,
  {32'hc44dd699, 32'h00000000} /* (6, 19, 6) {real, imag} */,
  {32'hc50b7868, 32'h00000000} /* (6, 19, 5) {real, imag} */,
  {32'hc51c4238, 32'h00000000} /* (6, 19, 4) {real, imag} */,
  {32'hc515608a, 32'h00000000} /* (6, 19, 3) {real, imag} */,
  {32'hc532c918, 32'h00000000} /* (6, 19, 2) {real, imag} */,
  {32'hc54d6901, 32'h00000000} /* (6, 19, 1) {real, imag} */,
  {32'hc51935a2, 32'h00000000} /* (6, 19, 0) {real, imag} */,
  {32'hc545d692, 32'h00000000} /* (6, 18, 31) {real, imag} */,
  {32'hc53f0720, 32'h00000000} /* (6, 18, 30) {real, imag} */,
  {32'hc53abac2, 32'h00000000} /* (6, 18, 29) {real, imag} */,
  {32'hc5359248, 32'h00000000} /* (6, 18, 28) {real, imag} */,
  {32'hc54a6de3, 32'h00000000} /* (6, 18, 27) {real, imag} */,
  {32'hc541690c, 32'h00000000} /* (6, 18, 26) {real, imag} */,
  {32'hc539bf1b, 32'h00000000} /* (6, 18, 25) {real, imag} */,
  {32'hc58b505a, 32'h00000000} /* (6, 18, 24) {real, imag} */,
  {32'hc5176dd2, 32'h00000000} /* (6, 18, 23) {real, imag} */,
  {32'hc457cf78, 32'h00000000} /* (6, 18, 22) {real, imag} */,
  {32'hc17f7780, 32'h00000000} /* (6, 18, 21) {real, imag} */,
  {32'h4513e0f3, 32'h00000000} /* (6, 18, 20) {real, imag} */,
  {32'h455b44c5, 32'h00000000} /* (6, 18, 19) {real, imag} */,
  {32'h456b77de, 32'h00000000} /* (6, 18, 18) {real, imag} */,
  {32'h458beef2, 32'h00000000} /* (6, 18, 17) {real, imag} */,
  {32'h4584450e, 32'h00000000} /* (6, 18, 16) {real, imag} */,
  {32'h457e723a, 32'h00000000} /* (6, 18, 15) {real, imag} */,
  {32'h45751a26, 32'h00000000} /* (6, 18, 14) {real, imag} */,
  {32'h45621036, 32'h00000000} /* (6, 18, 13) {real, imag} */,
  {32'h44f3dcac, 32'h00000000} /* (6, 18, 12) {real, imag} */,
  {32'h442addec, 32'h00000000} /* (6, 18, 11) {real, imag} */,
  {32'hc3ab197c, 32'h00000000} /* (6, 18, 10) {real, imag} */,
  {32'hc4a7b31a, 32'h00000000} /* (6, 18, 9) {real, imag} */,
  {32'hc52afd44, 32'h00000000} /* (6, 18, 8) {real, imag} */,
  {32'hc4f409ec, 32'h00000000} /* (6, 18, 7) {real, imag} */,
  {32'hc4fa552a, 32'h00000000} /* (6, 18, 6) {real, imag} */,
  {32'hc50ba172, 32'h00000000} /* (6, 18, 5) {real, imag} */,
  {32'hc556df1b, 32'h00000000} /* (6, 18, 4) {real, imag} */,
  {32'hc57052b5, 32'h00000000} /* (6, 18, 3) {real, imag} */,
  {32'hc55900a4, 32'h00000000} /* (6, 18, 2) {real, imag} */,
  {32'hc54c842c, 32'h00000000} /* (6, 18, 1) {real, imag} */,
  {32'hc547414c, 32'h00000000} /* (6, 18, 0) {real, imag} */,
  {32'hc566605a, 32'h00000000} /* (6, 17, 31) {real, imag} */,
  {32'hc57fd9bb, 32'h00000000} /* (6, 17, 30) {real, imag} */,
  {32'hc57a8169, 32'h00000000} /* (6, 17, 29) {real, imag} */,
  {32'hc569d33a, 32'h00000000} /* (6, 17, 28) {real, imag} */,
  {32'hc55e69e8, 32'h00000000} /* (6, 17, 27) {real, imag} */,
  {32'hc56b12c9, 32'h00000000} /* (6, 17, 26) {real, imag} */,
  {32'hc58ea239, 32'h00000000} /* (6, 17, 25) {real, imag} */,
  {32'hc56eedbe, 32'h00000000} /* (6, 17, 24) {real, imag} */,
  {32'hc5092988, 32'h00000000} /* (6, 17, 23) {real, imag} */,
  {32'hc4b192f6, 32'h00000000} /* (6, 17, 22) {real, imag} */,
  {32'h41f4b680, 32'h00000000} /* (6, 17, 21) {real, imag} */,
  {32'h4501ed58, 32'h00000000} /* (6, 17, 20) {real, imag} */,
  {32'h4531814c, 32'h00000000} /* (6, 17, 19) {real, imag} */,
  {32'h455ba022, 32'h00000000} /* (6, 17, 18) {real, imag} */,
  {32'h45963e2e, 32'h00000000} /* (6, 17, 17) {real, imag} */,
  {32'h458be4dd, 32'h00000000} /* (6, 17, 16) {real, imag} */,
  {32'h459023ff, 32'h00000000} /* (6, 17, 15) {real, imag} */,
  {32'h4583b290, 32'h00000000} /* (6, 17, 14) {real, imag} */,
  {32'h45617769, 32'h00000000} /* (6, 17, 13) {real, imag} */,
  {32'h45431cbc, 32'h00000000} /* (6, 17, 12) {real, imag} */,
  {32'h4413df08, 32'h00000000} /* (6, 17, 11) {real, imag} */,
  {32'hc499e8fe, 32'h00000000} /* (6, 17, 10) {real, imag} */,
  {32'hc529d34e, 32'h00000000} /* (6, 17, 9) {real, imag} */,
  {32'hc4cc61ed, 32'h00000000} /* (6, 17, 8) {real, imag} */,
  {32'hc5466948, 32'h00000000} /* (6, 17, 7) {real, imag} */,
  {32'hc57ef44b, 32'h00000000} /* (6, 17, 6) {real, imag} */,
  {32'hc564a1ab, 32'h00000000} /* (6, 17, 5) {real, imag} */,
  {32'hc57b9f6c, 32'h00000000} /* (6, 17, 4) {real, imag} */,
  {32'hc58291f1, 32'h00000000} /* (6, 17, 3) {real, imag} */,
  {32'hc5743f5a, 32'h00000000} /* (6, 17, 2) {real, imag} */,
  {32'hc56fe26c, 32'h00000000} /* (6, 17, 1) {real, imag} */,
  {32'hc562a23a, 32'h00000000} /* (6, 17, 0) {real, imag} */,
  {32'hc568f52d, 32'h00000000} /* (6, 16, 31) {real, imag} */,
  {32'hc58af931, 32'h00000000} /* (6, 16, 30) {real, imag} */,
  {32'hc59c8e4a, 32'h00000000} /* (6, 16, 29) {real, imag} */,
  {32'hc5795ebe, 32'h00000000} /* (6, 16, 28) {real, imag} */,
  {32'hc58bdaee, 32'h00000000} /* (6, 16, 27) {real, imag} */,
  {32'hc58a2a24, 32'h00000000} /* (6, 16, 26) {real, imag} */,
  {32'hc56d1d5e, 32'h00000000} /* (6, 16, 25) {real, imag} */,
  {32'hc561b851, 32'h00000000} /* (6, 16, 24) {real, imag} */,
  {32'hc50c22a2, 32'h00000000} /* (6, 16, 23) {real, imag} */,
  {32'hc50c253a, 32'h00000000} /* (6, 16, 22) {real, imag} */,
  {32'hc3cb2b00, 32'h00000000} /* (6, 16, 21) {real, imag} */,
  {32'h44e6eb3e, 32'h00000000} /* (6, 16, 20) {real, imag} */,
  {32'h4529643e, 32'h00000000} /* (6, 16, 19) {real, imag} */,
  {32'h4552ddc8, 32'h00000000} /* (6, 16, 18) {real, imag} */,
  {32'h45624d5c, 32'h00000000} /* (6, 16, 17) {real, imag} */,
  {32'h458673d9, 32'h00000000} /* (6, 16, 16) {real, imag} */,
  {32'h45a982a4, 32'h00000000} /* (6, 16, 15) {real, imag} */,
  {32'h457eeb62, 32'h00000000} /* (6, 16, 14) {real, imag} */,
  {32'h454e50c4, 32'h00000000} /* (6, 16, 13) {real, imag} */,
  {32'h4509b9e6, 32'h00000000} /* (6, 16, 12) {real, imag} */,
  {32'h43a97260, 32'h00000000} /* (6, 16, 11) {real, imag} */,
  {32'hc46662f2, 32'h00000000} /* (6, 16, 10) {real, imag} */,
  {32'hc509e9ae, 32'h00000000} /* (6, 16, 9) {real, imag} */,
  {32'hc54fbe5b, 32'h00000000} /* (6, 16, 8) {real, imag} */,
  {32'hc5906802, 32'h00000000} /* (6, 16, 7) {real, imag} */,
  {32'hc569944a, 32'h00000000} /* (6, 16, 6) {real, imag} */,
  {32'hc586b42c, 32'h00000000} /* (6, 16, 5) {real, imag} */,
  {32'hc5a2385e, 32'h00000000} /* (6, 16, 4) {real, imag} */,
  {32'hc5a344f1, 32'h00000000} /* (6, 16, 3) {real, imag} */,
  {32'hc5ae1606, 32'h00000000} /* (6, 16, 2) {real, imag} */,
  {32'hc5c6fa3e, 32'h00000000} /* (6, 16, 1) {real, imag} */,
  {32'hc58adc2b, 32'h00000000} /* (6, 16, 0) {real, imag} */,
  {32'hc5598693, 32'h00000000} /* (6, 15, 31) {real, imag} */,
  {32'hc584dc81, 32'h00000000} /* (6, 15, 30) {real, imag} */,
  {32'hc57f1fdb, 32'h00000000} /* (6, 15, 29) {real, imag} */,
  {32'hc58ce1f2, 32'h00000000} /* (6, 15, 28) {real, imag} */,
  {32'hc59fdc52, 32'h00000000} /* (6, 15, 27) {real, imag} */,
  {32'hc56f8d2e, 32'h00000000} /* (6, 15, 26) {real, imag} */,
  {32'hc59a781c, 32'h00000000} /* (6, 15, 25) {real, imag} */,
  {32'hc562fa11, 32'h00000000} /* (6, 15, 24) {real, imag} */,
  {32'hc52effa2, 32'h00000000} /* (6, 15, 23) {real, imag} */,
  {32'hc4beee49, 32'h00000000} /* (6, 15, 22) {real, imag} */,
  {32'hc23e5d00, 32'h00000000} /* (6, 15, 21) {real, imag} */,
  {32'h450e2432, 32'h00000000} /* (6, 15, 20) {real, imag} */,
  {32'h45428bf8, 32'h00000000} /* (6, 15, 19) {real, imag} */,
  {32'h4531a37c, 32'h00000000} /* (6, 15, 18) {real, imag} */,
  {32'h453bb734, 32'h00000000} /* (6, 15, 17) {real, imag} */,
  {32'h45938e7a, 32'h00000000} /* (6, 15, 16) {real, imag} */,
  {32'h458191da, 32'h00000000} /* (6, 15, 15) {real, imag} */,
  {32'h45634e1a, 32'h00000000} /* (6, 15, 14) {real, imag} */,
  {32'h4537cd1f, 32'h00000000} /* (6, 15, 13) {real, imag} */,
  {32'h44b18d2f, 32'h00000000} /* (6, 15, 12) {real, imag} */,
  {32'h43a36e08, 32'h00000000} /* (6, 15, 11) {real, imag} */,
  {32'hc43640da, 32'h00000000} /* (6, 15, 10) {real, imag} */,
  {32'hc51d3d67, 32'h00000000} /* (6, 15, 9) {real, imag} */,
  {32'hc568a9c5, 32'h00000000} /* (6, 15, 8) {real, imag} */,
  {32'hc58c960f, 32'h00000000} /* (6, 15, 7) {real, imag} */,
  {32'hc5843da1, 32'h00000000} /* (6, 15, 6) {real, imag} */,
  {32'hc569d3c8, 32'h00000000} /* (6, 15, 5) {real, imag} */,
  {32'hc58fff01, 32'h00000000} /* (6, 15, 4) {real, imag} */,
  {32'hc5bc18bc, 32'h00000000} /* (6, 15, 3) {real, imag} */,
  {32'hc5ce41e0, 32'h00000000} /* (6, 15, 2) {real, imag} */,
  {32'hc5be2384, 32'h00000000} /* (6, 15, 1) {real, imag} */,
  {32'hc58a059c, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'hc555dc43, 32'h00000000} /* (6, 14, 31) {real, imag} */,
  {32'hc56b7316, 32'h00000000} /* (6, 14, 30) {real, imag} */,
  {32'hc578e5e0, 32'h00000000} /* (6, 14, 29) {real, imag} */,
  {32'hc58d3434, 32'h00000000} /* (6, 14, 28) {real, imag} */,
  {32'hc5751890, 32'h00000000} /* (6, 14, 27) {real, imag} */,
  {32'hc59405be, 32'h00000000} /* (6, 14, 26) {real, imag} */,
  {32'hc597d164, 32'h00000000} /* (6, 14, 25) {real, imag} */,
  {32'hc56d9fda, 32'h00000000} /* (6, 14, 24) {real, imag} */,
  {32'hc5787920, 32'h00000000} /* (6, 14, 23) {real, imag} */,
  {32'hc4f31fd4, 32'h00000000} /* (6, 14, 22) {real, imag} */,
  {32'h4241e300, 32'h00000000} /* (6, 14, 21) {real, imag} */,
  {32'h450837f8, 32'h00000000} /* (6, 14, 20) {real, imag} */,
  {32'h44d5e434, 32'h00000000} /* (6, 14, 19) {real, imag} */,
  {32'h450d8738, 32'h00000000} /* (6, 14, 18) {real, imag} */,
  {32'h453233fb, 32'h00000000} /* (6, 14, 17) {real, imag} */,
  {32'h456a1885, 32'h00000000} /* (6, 14, 16) {real, imag} */,
  {32'h454b479f, 32'h00000000} /* (6, 14, 15) {real, imag} */,
  {32'h456ad2c8, 32'h00000000} /* (6, 14, 14) {real, imag} */,
  {32'h453942cc, 32'h00000000} /* (6, 14, 13) {real, imag} */,
  {32'h44acb315, 32'h00000000} /* (6, 14, 12) {real, imag} */,
  {32'h443fc298, 32'h00000000} /* (6, 14, 11) {real, imag} */,
  {32'hc5319b3b, 32'h00000000} /* (6, 14, 10) {real, imag} */,
  {32'hc544a651, 32'h00000000} /* (6, 14, 9) {real, imag} */,
  {32'hc531b584, 32'h00000000} /* (6, 14, 8) {real, imag} */,
  {32'hc5826a6c, 32'h00000000} /* (6, 14, 7) {real, imag} */,
  {32'hc591dbbc, 32'h00000000} /* (6, 14, 6) {real, imag} */,
  {32'hc587a262, 32'h00000000} /* (6, 14, 5) {real, imag} */,
  {32'hc58773b9, 32'h00000000} /* (6, 14, 4) {real, imag} */,
  {32'hc591b3a2, 32'h00000000} /* (6, 14, 3) {real, imag} */,
  {32'hc5ad0034, 32'h00000000} /* (6, 14, 2) {real, imag} */,
  {32'hc57b934f, 32'h00000000} /* (6, 14, 1) {real, imag} */,
  {32'hc55191b3, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hc52e5b20, 32'h00000000} /* (6, 13, 31) {real, imag} */,
  {32'hc5542d76, 32'h00000000} /* (6, 13, 30) {real, imag} */,
  {32'hc55b13cf, 32'h00000000} /* (6, 13, 29) {real, imag} */,
  {32'hc566ddfd, 32'h00000000} /* (6, 13, 28) {real, imag} */,
  {32'hc5739697, 32'h00000000} /* (6, 13, 27) {real, imag} */,
  {32'hc54adf1f, 32'h00000000} /* (6, 13, 26) {real, imag} */,
  {32'hc571aee2, 32'h00000000} /* (6, 13, 25) {real, imag} */,
  {32'hc5919cd4, 32'h00000000} /* (6, 13, 24) {real, imag} */,
  {32'hc51f2e74, 32'h00000000} /* (6, 13, 23) {real, imag} */,
  {32'hc4e5c302, 32'h00000000} /* (6, 13, 22) {real, imag} */,
  {32'hc4420ed8, 32'h00000000} /* (6, 13, 21) {real, imag} */,
  {32'h44f170bc, 32'h00000000} /* (6, 13, 20) {real, imag} */,
  {32'h449bd45e, 32'h00000000} /* (6, 13, 19) {real, imag} */,
  {32'h450865f8, 32'h00000000} /* (6, 13, 18) {real, imag} */,
  {32'h452e4027, 32'h00000000} /* (6, 13, 17) {real, imag} */,
  {32'h452bbba5, 32'h00000000} /* (6, 13, 16) {real, imag} */,
  {32'h4552aeea, 32'h00000000} /* (6, 13, 15) {real, imag} */,
  {32'h4502a2ec, 32'h00000000} /* (6, 13, 14) {real, imag} */,
  {32'h454480b5, 32'h00000000} /* (6, 13, 13) {real, imag} */,
  {32'h44bb964e, 32'h00000000} /* (6, 13, 12) {real, imag} */,
  {32'h4460f35c, 32'h00000000} /* (6, 13, 11) {real, imag} */,
  {32'hc5303e89, 32'h00000000} /* (6, 13, 10) {real, imag} */,
  {32'hc590fb53, 32'h00000000} /* (6, 13, 9) {real, imag} */,
  {32'hc50ed93a, 32'h00000000} /* (6, 13, 8) {real, imag} */,
  {32'hc593fafb, 32'h00000000} /* (6, 13, 7) {real, imag} */,
  {32'hc59022bc, 32'h00000000} /* (6, 13, 6) {real, imag} */,
  {32'hc554e794, 32'h00000000} /* (6, 13, 5) {real, imag} */,
  {32'hc580da04, 32'h00000000} /* (6, 13, 4) {real, imag} */,
  {32'hc59e14c0, 32'h00000000} /* (6, 13, 3) {real, imag} */,
  {32'hc563dbe4, 32'h00000000} /* (6, 13, 2) {real, imag} */,
  {32'hc52f5801, 32'h00000000} /* (6, 13, 1) {real, imag} */,
  {32'hc50ae2d3, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'hc4d9e008, 32'h00000000} /* (6, 12, 31) {real, imag} */,
  {32'hc516f286, 32'h00000000} /* (6, 12, 30) {real, imag} */,
  {32'hc5010bdc, 32'h00000000} /* (6, 12, 29) {real, imag} */,
  {32'hc4f7f9d1, 32'h00000000} /* (6, 12, 28) {real, imag} */,
  {32'hc517acb4, 32'h00000000} /* (6, 12, 27) {real, imag} */,
  {32'hc53aed7f, 32'h00000000} /* (6, 12, 26) {real, imag} */,
  {32'hc531b3ab, 32'h00000000} /* (6, 12, 25) {real, imag} */,
  {32'hc532a53e, 32'h00000000} /* (6, 12, 24) {real, imag} */,
  {32'hc50a124d, 32'h00000000} /* (6, 12, 23) {real, imag} */,
  {32'hc3986004, 32'h00000000} /* (6, 12, 22) {real, imag} */,
  {32'hc42edc08, 32'h00000000} /* (6, 12, 21) {real, imag} */,
  {32'h4486013a, 32'h00000000} /* (6, 12, 20) {real, imag} */,
  {32'h44b84129, 32'h00000000} /* (6, 12, 19) {real, imag} */,
  {32'h449685bb, 32'h00000000} /* (6, 12, 18) {real, imag} */,
  {32'h4520a43a, 32'h00000000} /* (6, 12, 17) {real, imag} */,
  {32'h4514c42c, 32'h00000000} /* (6, 12, 16) {real, imag} */,
  {32'h44f085a0, 32'h00000000} /* (6, 12, 15) {real, imag} */,
  {32'h450048bc, 32'h00000000} /* (6, 12, 14) {real, imag} */,
  {32'h4513e13e, 32'h00000000} /* (6, 12, 13) {real, imag} */,
  {32'h45586538, 32'h00000000} /* (6, 12, 12) {real, imag} */,
  {32'hc2524be0, 32'h00000000} /* (6, 12, 11) {real, imag} */,
  {32'hc49d7312, 32'h00000000} /* (6, 12, 10) {real, imag} */,
  {32'hc4ed3db9, 32'h00000000} /* (6, 12, 9) {real, imag} */,
  {32'hc55f66cc, 32'h00000000} /* (6, 12, 8) {real, imag} */,
  {32'hc5249ab1, 32'h00000000} /* (6, 12, 7) {real, imag} */,
  {32'hc552f066, 32'h00000000} /* (6, 12, 6) {real, imag} */,
  {32'hc549cfe4, 32'h00000000} /* (6, 12, 5) {real, imag} */,
  {32'hc538c4d8, 32'h00000000} /* (6, 12, 4) {real, imag} */,
  {32'hc5283358, 32'h00000000} /* (6, 12, 3) {real, imag} */,
  {32'hc5299e6e, 32'h00000000} /* (6, 12, 2) {real, imag} */,
  {32'hc505d3b2, 32'h00000000} /* (6, 12, 1) {real, imag} */,
  {32'hc4bdb3e5, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'hc1aa0e00, 32'h00000000} /* (6, 11, 31) {real, imag} */,
  {32'hc13b3c40, 32'h00000000} /* (6, 11, 30) {real, imag} */,
  {32'hc4b10509, 32'h00000000} /* (6, 11, 29) {real, imag} */,
  {32'hc49ecaeb, 32'h00000000} /* (6, 11, 28) {real, imag} */,
  {32'hc4b4542d, 32'h00000000} /* (6, 11, 27) {real, imag} */,
  {32'hc4bbeb4a, 32'h00000000} /* (6, 11, 26) {real, imag} */,
  {32'hc4adda77, 32'h00000000} /* (6, 11, 25) {real, imag} */,
  {32'hc43f8b50, 32'h00000000} /* (6, 11, 24) {real, imag} */,
  {32'hc33cde58, 32'h00000000} /* (6, 11, 23) {real, imag} */,
  {32'h430eb158, 32'h00000000} /* (6, 11, 22) {real, imag} */,
  {32'h434b5b50, 32'h00000000} /* (6, 11, 21) {real, imag} */,
  {32'h44669400, 32'h00000000} /* (6, 11, 20) {real, imag} */,
  {32'h4431d268, 32'h00000000} /* (6, 11, 19) {real, imag} */,
  {32'h4470aa86, 32'h00000000} /* (6, 11, 18) {real, imag} */,
  {32'h44c98f41, 32'h00000000} /* (6, 11, 17) {real, imag} */,
  {32'h44aac48e, 32'h00000000} /* (6, 11, 16) {real, imag} */,
  {32'h4431dcd5, 32'h00000000} /* (6, 11, 15) {real, imag} */,
  {32'h44c79c4c, 32'h00000000} /* (6, 11, 14) {real, imag} */,
  {32'h44bd9dc5, 32'h00000000} /* (6, 11, 13) {real, imag} */,
  {32'h443d25fc, 32'h00000000} /* (6, 11, 12) {real, imag} */,
  {32'h435f1a80, 32'h00000000} /* (6, 11, 11) {real, imag} */,
  {32'hc4779efc, 32'h00000000} /* (6, 11, 10) {real, imag} */,
  {32'hc515a292, 32'h00000000} /* (6, 11, 9) {real, imag} */,
  {32'hc50ee7d4, 32'h00000000} /* (6, 11, 8) {real, imag} */,
  {32'hc4f5a4ab, 32'h00000000} /* (6, 11, 7) {real, imag} */,
  {32'hc51b4936, 32'h00000000} /* (6, 11, 6) {real, imag} */,
  {32'hc531ae13, 32'h00000000} /* (6, 11, 5) {real, imag} */,
  {32'hc521899b, 32'h00000000} /* (6, 11, 4) {real, imag} */,
  {32'hc481b180, 32'h00000000} /* (6, 11, 3) {real, imag} */,
  {32'hc4d5a5dd, 32'h00000000} /* (6, 11, 2) {real, imag} */,
  {32'hc48fcc6b, 32'h00000000} /* (6, 11, 1) {real, imag} */,
  {32'hc2e7f2b8, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h44d364d9, 32'h00000000} /* (6, 10, 31) {real, imag} */,
  {32'h44d5f81d, 32'h00000000} /* (6, 10, 30) {real, imag} */,
  {32'h44c925f3, 32'h00000000} /* (6, 10, 29) {real, imag} */,
  {32'h451d568d, 32'h00000000} /* (6, 10, 28) {real, imag} */,
  {32'h44e84850, 32'h00000000} /* (6, 10, 27) {real, imag} */,
  {32'h4470fb96, 32'h00000000} /* (6, 10, 26) {real, imag} */,
  {32'h44f1fd24, 32'h00000000} /* (6, 10, 25) {real, imag} */,
  {32'h45111775, 32'h00000000} /* (6, 10, 24) {real, imag} */,
  {32'h45048c07, 32'h00000000} /* (6, 10, 23) {real, imag} */,
  {32'h451122ec, 32'h00000000} /* (6, 10, 22) {real, imag} */,
  {32'h44ee6693, 32'h00000000} /* (6, 10, 21) {real, imag} */,
  {32'h441bb10a, 32'h00000000} /* (6, 10, 20) {real, imag} */,
  {32'hc436a49f, 32'h00000000} /* (6, 10, 19) {real, imag} */,
  {32'h435014b0, 32'h00000000} /* (6, 10, 18) {real, imag} */,
  {32'hc44cffb4, 32'h00000000} /* (6, 10, 17) {real, imag} */,
  {32'hc41d544d, 32'h00000000} /* (6, 10, 16) {real, imag} */,
  {32'hc2eeaf90, 32'h00000000} /* (6, 10, 15) {real, imag} */,
  {32'hc344f9d8, 32'h00000000} /* (6, 10, 14) {real, imag} */,
  {32'hc3ecee34, 32'h00000000} /* (6, 10, 13) {real, imag} */,
  {32'hc46f6160, 32'h00000000} /* (6, 10, 12) {real, imag} */,
  {32'hc489a9d6, 32'h00000000} /* (6, 10, 11) {real, imag} */,
  {32'hc4879dd9, 32'h00000000} /* (6, 10, 10) {real, imag} */,
  {32'hc2781f90, 32'h00000000} /* (6, 10, 9) {real, imag} */,
  {32'hc3e979b2, 32'h00000000} /* (6, 10, 8) {real, imag} */,
  {32'h4416facd, 32'h00000000} /* (6, 10, 7) {real, imag} */,
  {32'h43cf751c, 32'h00000000} /* (6, 10, 6) {real, imag} */,
  {32'h439838c4, 32'h00000000} /* (6, 10, 5) {real, imag} */,
  {32'h443cb566, 32'h00000000} /* (6, 10, 4) {real, imag} */,
  {32'h43f15ca2, 32'h00000000} /* (6, 10, 3) {real, imag} */,
  {32'h43f6f488, 32'h00000000} /* (6, 10, 2) {real, imag} */,
  {32'h44d72e80, 32'h00000000} /* (6, 10, 1) {real, imag} */,
  {32'h44fdb36c, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'h454e5927, 32'h00000000} /* (6, 9, 31) {real, imag} */,
  {32'h45894af8, 32'h00000000} /* (6, 9, 30) {real, imag} */,
  {32'h455c5483, 32'h00000000} /* (6, 9, 29) {real, imag} */,
  {32'h453a36fd, 32'h00000000} /* (6, 9, 28) {real, imag} */,
  {32'h4592b004, 32'h00000000} /* (6, 9, 27) {real, imag} */,
  {32'h4556cec0, 32'h00000000} /* (6, 9, 26) {real, imag} */,
  {32'h455a5620, 32'h00000000} /* (6, 9, 25) {real, imag} */,
  {32'h454bbe74, 32'h00000000} /* (6, 9, 24) {real, imag} */,
  {32'h4593491a, 32'h00000000} /* (6, 9, 23) {real, imag} */,
  {32'h458e0f1a, 32'h00000000} /* (6, 9, 22) {real, imag} */,
  {32'h45527925, 32'h00000000} /* (6, 9, 21) {real, imag} */,
  {32'hc3955986, 32'h00000000} /* (6, 9, 20) {real, imag} */,
  {32'hc31c7990, 32'h00000000} /* (6, 9, 19) {real, imag} */,
  {32'hc3918ebc, 32'h00000000} /* (6, 9, 18) {real, imag} */,
  {32'hc50ba432, 32'h00000000} /* (6, 9, 17) {real, imag} */,
  {32'hc4d022fa, 32'h00000000} /* (6, 9, 16) {real, imag} */,
  {32'hc490f972, 32'h00000000} /* (6, 9, 15) {real, imag} */,
  {32'hc4d0fcf0, 32'h00000000} /* (6, 9, 14) {real, imag} */,
  {32'hc4b1e52a, 32'h00000000} /* (6, 9, 13) {real, imag} */,
  {32'hc499c6e6, 32'h00000000} /* (6, 9, 12) {real, imag} */,
  {32'hc5070fd9, 32'h00000000} /* (6, 9, 11) {real, imag} */,
  {32'hc4631ca8, 32'h00000000} /* (6, 9, 10) {real, imag} */,
  {32'h432e6c40, 32'h00000000} /* (6, 9, 9) {real, imag} */,
  {32'h44c79d53, 32'h00000000} /* (6, 9, 8) {real, imag} */,
  {32'h453c2b22, 32'h00000000} /* (6, 9, 7) {real, imag} */,
  {32'h44ba2046, 32'h00000000} /* (6, 9, 6) {real, imag} */,
  {32'h44d56fb2, 32'h00000000} /* (6, 9, 5) {real, imag} */,
  {32'h450d2cf7, 32'h00000000} /* (6, 9, 4) {real, imag} */,
  {32'h452dfbb3, 32'h00000000} /* (6, 9, 3) {real, imag} */,
  {32'h4558073c, 32'h00000000} /* (6, 9, 2) {real, imag} */,
  {32'h453e27f6, 32'h00000000} /* (6, 9, 1) {real, imag} */,
  {32'h4532f0d7, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'h4575a438, 32'h00000000} /* (6, 8, 31) {real, imag} */,
  {32'h45abb67b, 32'h00000000} /* (6, 8, 30) {real, imag} */,
  {32'h458cdeec, 32'h00000000} /* (6, 8, 29) {real, imag} */,
  {32'h45614308, 32'h00000000} /* (6, 8, 28) {real, imag} */,
  {32'h4582172c, 32'h00000000} /* (6, 8, 27) {real, imag} */,
  {32'h458406ad, 32'h00000000} /* (6, 8, 26) {real, imag} */,
  {32'h455c351a, 32'h00000000} /* (6, 8, 25) {real, imag} */,
  {32'h458048d5, 32'h00000000} /* (6, 8, 24) {real, imag} */,
  {32'h459670b6, 32'h00000000} /* (6, 8, 23) {real, imag} */,
  {32'h4592b924, 32'h00000000} /* (6, 8, 22) {real, imag} */,
  {32'h4546b130, 32'h00000000} /* (6, 8, 21) {real, imag} */,
  {32'h448d7ba6, 32'h00000000} /* (6, 8, 20) {real, imag} */,
  {32'h43694300, 32'h00000000} /* (6, 8, 19) {real, imag} */,
  {32'hc3a943bc, 32'h00000000} /* (6, 8, 18) {real, imag} */,
  {32'hc4b68255, 32'h00000000} /* (6, 8, 17) {real, imag} */,
  {32'hc523ae9b, 32'h00000000} /* (6, 8, 16) {real, imag} */,
  {32'hc503435e, 32'h00000000} /* (6, 8, 15) {real, imag} */,
  {32'hc527de34, 32'h00000000} /* (6, 8, 14) {real, imag} */,
  {32'hc526a4ba, 32'h00000000} /* (6, 8, 13) {real, imag} */,
  {32'hc4e2e210, 32'h00000000} /* (6, 8, 12) {real, imag} */,
  {32'hc4cac508, 32'h00000000} /* (6, 8, 11) {real, imag} */,
  {32'hc35f03b8, 32'h00000000} /* (6, 8, 10) {real, imag} */,
  {32'h43a3a444, 32'h00000000} /* (6, 8, 9) {real, imag} */,
  {32'h44fb6ec7, 32'h00000000} /* (6, 8, 8) {real, imag} */,
  {32'h452d33b9, 32'h00000000} /* (6, 8, 7) {real, imag} */,
  {32'h4523fb45, 32'h00000000} /* (6, 8, 6) {real, imag} */,
  {32'h450422c6, 32'h00000000} /* (6, 8, 5) {real, imag} */,
  {32'h4547473d, 32'h00000000} /* (6, 8, 4) {real, imag} */,
  {32'h459498dd, 32'h00000000} /* (6, 8, 3) {real, imag} */,
  {32'h45873654, 32'h00000000} /* (6, 8, 2) {real, imag} */,
  {32'h45875ac6, 32'h00000000} /* (6, 8, 1) {real, imag} */,
  {32'h458ea0c0, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h45b10b5b, 32'h00000000} /* (6, 7, 31) {real, imag} */,
  {32'h45a6a151, 32'h00000000} /* (6, 7, 30) {real, imag} */,
  {32'h45906598, 32'h00000000} /* (6, 7, 29) {real, imag} */,
  {32'h4594a638, 32'h00000000} /* (6, 7, 28) {real, imag} */,
  {32'h458e258c, 32'h00000000} /* (6, 7, 27) {real, imag} */,
  {32'h459b42e9, 32'h00000000} /* (6, 7, 26) {real, imag} */,
  {32'h458eec0d, 32'h00000000} /* (6, 7, 25) {real, imag} */,
  {32'h45a2d918, 32'h00000000} /* (6, 7, 24) {real, imag} */,
  {32'h45a9356c, 32'h00000000} /* (6, 7, 23) {real, imag} */,
  {32'h45a62252, 32'h00000000} /* (6, 7, 22) {real, imag} */,
  {32'h458154d6, 32'h00000000} /* (6, 7, 21) {real, imag} */,
  {32'h44f0c93b, 32'h00000000} /* (6, 7, 20) {real, imag} */,
  {32'h4426ef48, 32'h00000000} /* (6, 7, 19) {real, imag} */,
  {32'hc33764d0, 32'h00000000} /* (6, 7, 18) {real, imag} */,
  {32'hc4a9e74c, 32'h00000000} /* (6, 7, 17) {real, imag} */,
  {32'hc521f56c, 32'h00000000} /* (6, 7, 16) {real, imag} */,
  {32'hc554977e, 32'h00000000} /* (6, 7, 15) {real, imag} */,
  {32'hc55774e2, 32'h00000000} /* (6, 7, 14) {real, imag} */,
  {32'hc57ad65f, 32'h00000000} /* (6, 7, 13) {real, imag} */,
  {32'hc534aba8, 32'h00000000} /* (6, 7, 12) {real, imag} */,
  {32'hc4bb2a10, 32'h00000000} /* (6, 7, 11) {real, imag} */,
  {32'hc3f75fd0, 32'h00000000} /* (6, 7, 10) {real, imag} */,
  {32'h444de782, 32'h00000000} /* (6, 7, 9) {real, imag} */,
  {32'h45042a58, 32'h00000000} /* (6, 7, 8) {real, imag} */,
  {32'h44ce9886, 32'h00000000} /* (6, 7, 7) {real, imag} */,
  {32'h45336c04, 32'h00000000} /* (6, 7, 6) {real, imag} */,
  {32'h456ce6b2, 32'h00000000} /* (6, 7, 5) {real, imag} */,
  {32'h45854525, 32'h00000000} /* (6, 7, 4) {real, imag} */,
  {32'h459f1d8d, 32'h00000000} /* (6, 7, 3) {real, imag} */,
  {32'h45b6a52a, 32'h00000000} /* (6, 7, 2) {real, imag} */,
  {32'h459e0d36, 32'h00000000} /* (6, 7, 1) {real, imag} */,
  {32'h459c8696, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'h45b1e27c, 32'h00000000} /* (6, 6, 31) {real, imag} */,
  {32'h45c3c679, 32'h00000000} /* (6, 6, 30) {real, imag} */,
  {32'h45c49f3d, 32'h00000000} /* (6, 6, 29) {real, imag} */,
  {32'h45a4fb2f, 32'h00000000} /* (6, 6, 28) {real, imag} */,
  {32'h45c43f87, 32'h00000000} /* (6, 6, 27) {real, imag} */,
  {32'h45b75438, 32'h00000000} /* (6, 6, 26) {real, imag} */,
  {32'h45a5f398, 32'h00000000} /* (6, 6, 25) {real, imag} */,
  {32'h45c0fe2c, 32'h00000000} /* (6, 6, 24) {real, imag} */,
  {32'h45b0418d, 32'h00000000} /* (6, 6, 23) {real, imag} */,
  {32'h45ab127e, 32'h00000000} /* (6, 6, 22) {real, imag} */,
  {32'h4585d73f, 32'h00000000} /* (6, 6, 21) {real, imag} */,
  {32'h44be9a38, 32'h00000000} /* (6, 6, 20) {real, imag} */,
  {32'h447f5f06, 32'h00000000} /* (6, 6, 19) {real, imag} */,
  {32'hc3bfd970, 32'h00000000} /* (6, 6, 18) {real, imag} */,
  {32'hc49668b0, 32'h00000000} /* (6, 6, 17) {real, imag} */,
  {32'hc4d7d688, 32'h00000000} /* (6, 6, 16) {real, imag} */,
  {32'hc5330558, 32'h00000000} /* (6, 6, 15) {real, imag} */,
  {32'hc537a716, 32'h00000000} /* (6, 6, 14) {real, imag} */,
  {32'hc5293ee2, 32'h00000000} /* (6, 6, 13) {real, imag} */,
  {32'hc5638f7a, 32'h00000000} /* (6, 6, 12) {real, imag} */,
  {32'hc50187e2, 32'h00000000} /* (6, 6, 11) {real, imag} */,
  {32'h4396e200, 32'h00000000} /* (6, 6, 10) {real, imag} */,
  {32'h445bbdd0, 32'h00000000} /* (6, 6, 9) {real, imag} */,
  {32'h450171a8, 32'h00000000} /* (6, 6, 8) {real, imag} */,
  {32'h45259e06, 32'h00000000} /* (6, 6, 7) {real, imag} */,
  {32'h457c7d64, 32'h00000000} /* (6, 6, 6) {real, imag} */,
  {32'h45b5a86b, 32'h00000000} /* (6, 6, 5) {real, imag} */,
  {32'h45b57374, 32'h00000000} /* (6, 6, 4) {real, imag} */,
  {32'h4599da15, 32'h00000000} /* (6, 6, 3) {real, imag} */,
  {32'h45b97dcd, 32'h00000000} /* (6, 6, 2) {real, imag} */,
  {32'h45bff4d8, 32'h00000000} /* (6, 6, 1) {real, imag} */,
  {32'h45b5b9e3, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'h45e94a98, 32'h00000000} /* (6, 5, 31) {real, imag} */,
  {32'h45c8935e, 32'h00000000} /* (6, 5, 30) {real, imag} */,
  {32'h45bd804c, 32'h00000000} /* (6, 5, 29) {real, imag} */,
  {32'h45d13e12, 32'h00000000} /* (6, 5, 28) {real, imag} */,
  {32'h45cfce64, 32'h00000000} /* (6, 5, 27) {real, imag} */,
  {32'h45c5ec1a, 32'h00000000} /* (6, 5, 26) {real, imag} */,
  {32'h45cc2b4d, 32'h00000000} /* (6, 5, 25) {real, imag} */,
  {32'h45c43651, 32'h00000000} /* (6, 5, 24) {real, imag} */,
  {32'h45d678ce, 32'h00000000} /* (6, 5, 23) {real, imag} */,
  {32'h45b82874, 32'h00000000} /* (6, 5, 22) {real, imag} */,
  {32'h458e98ec, 32'h00000000} /* (6, 5, 21) {real, imag} */,
  {32'h4544537e, 32'h00000000} /* (6, 5, 20) {real, imag} */,
  {32'h451dfd68, 32'h00000000} /* (6, 5, 19) {real, imag} */,
  {32'h44617924, 32'h00000000} /* (6, 5, 18) {real, imag} */,
  {32'h439c35e8, 32'h00000000} /* (6, 5, 17) {real, imag} */,
  {32'hc3e0bde8, 32'h00000000} /* (6, 5, 16) {real, imag} */,
  {32'hc51d5af5, 32'h00000000} /* (6, 5, 15) {real, imag} */,
  {32'hc55b9ad4, 32'h00000000} /* (6, 5, 14) {real, imag} */,
  {32'hc53587ef, 32'h00000000} /* (6, 5, 13) {real, imag} */,
  {32'hc5329164, 32'h00000000} /* (6, 5, 12) {real, imag} */,
  {32'hc562d2c8, 32'h00000000} /* (6, 5, 11) {real, imag} */,
  {32'hc497df0c, 32'h00000000} /* (6, 5, 10) {real, imag} */,
  {32'hc3b6e1f0, 32'h00000000} /* (6, 5, 9) {real, imag} */,
  {32'hc46e6c78, 32'h00000000} /* (6, 5, 8) {real, imag} */,
  {32'h449279ba, 32'h00000000} /* (6, 5, 7) {real, imag} */,
  {32'h452dd418, 32'h00000000} /* (6, 5, 6) {real, imag} */,
  {32'h455961aa, 32'h00000000} /* (6, 5, 5) {real, imag} */,
  {32'h45a7146d, 32'h00000000} /* (6, 5, 4) {real, imag} */,
  {32'h45b53152, 32'h00000000} /* (6, 5, 3) {real, imag} */,
  {32'h45b724ac, 32'h00000000} /* (6, 5, 2) {real, imag} */,
  {32'h45bfecf6, 32'h00000000} /* (6, 5, 1) {real, imag} */,
  {32'h45bea12c, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'h45db3501, 32'h00000000} /* (6, 4, 31) {real, imag} */,
  {32'h45c447a7, 32'h00000000} /* (6, 4, 30) {real, imag} */,
  {32'h45c291ea, 32'h00000000} /* (6, 4, 29) {real, imag} */,
  {32'h45d5a4cf, 32'h00000000} /* (6, 4, 28) {real, imag} */,
  {32'h45d22a58, 32'h00000000} /* (6, 4, 27) {real, imag} */,
  {32'h45e1abb0, 32'h00000000} /* (6, 4, 26) {real, imag} */,
  {32'h45c83c7a, 32'h00000000} /* (6, 4, 25) {real, imag} */,
  {32'h45c80b21, 32'h00000000} /* (6, 4, 24) {real, imag} */,
  {32'h45c6d7a4, 32'h00000000} /* (6, 4, 23) {real, imag} */,
  {32'h45c05cf8, 32'h00000000} /* (6, 4, 22) {real, imag} */,
  {32'h4597b209, 32'h00000000} /* (6, 4, 21) {real, imag} */,
  {32'h45a04c6d, 32'h00000000} /* (6, 4, 20) {real, imag} */,
  {32'h4556ad37, 32'h00000000} /* (6, 4, 19) {real, imag} */,
  {32'h4545fc53, 32'h00000000} /* (6, 4, 18) {real, imag} */,
  {32'h44c91554, 32'h00000000} /* (6, 4, 17) {real, imag} */,
  {32'hc233b380, 32'h00000000} /* (6, 4, 16) {real, imag} */,
  {32'hc56b1c52, 32'h00000000} /* (6, 4, 15) {real, imag} */,
  {32'hc57efd0e, 32'h00000000} /* (6, 4, 14) {real, imag} */,
  {32'hc53680e1, 32'h00000000} /* (6, 4, 13) {real, imag} */,
  {32'hc56a213a, 32'h00000000} /* (6, 4, 12) {real, imag} */,
  {32'hc538d4cf, 32'h00000000} /* (6, 4, 11) {real, imag} */,
  {32'hc516c33c, 32'h00000000} /* (6, 4, 10) {real, imag} */,
  {32'hc4b06e60, 32'h00000000} /* (6, 4, 9) {real, imag} */,
  {32'hc4d6df58, 32'h00000000} /* (6, 4, 8) {real, imag} */,
  {32'hc4446bf4, 32'h00000000} /* (6, 4, 7) {real, imag} */,
  {32'h442704cc, 32'h00000000} /* (6, 4, 6) {real, imag} */,
  {32'h45320800, 32'h00000000} /* (6, 4, 5) {real, imag} */,
  {32'h45a37d89, 32'h00000000} /* (6, 4, 4) {real, imag} */,
  {32'h45b9bc54, 32'h00000000} /* (6, 4, 3) {real, imag} */,
  {32'h45bb4042, 32'h00000000} /* (6, 4, 2) {real, imag} */,
  {32'h45fa8087, 32'h00000000} /* (6, 4, 1) {real, imag} */,
  {32'h45da1a04, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'h45d902ab, 32'h00000000} /* (6, 3, 31) {real, imag} */,
  {32'h45e36010, 32'h00000000} /* (6, 3, 30) {real, imag} */,
  {32'h45d5f1bc, 32'h00000000} /* (6, 3, 29) {real, imag} */,
  {32'h45f06951, 32'h00000000} /* (6, 3, 28) {real, imag} */,
  {32'h45e89b8c, 32'h00000000} /* (6, 3, 27) {real, imag} */,
  {32'h45d95510, 32'h00000000} /* (6, 3, 26) {real, imag} */,
  {32'h45eff3df, 32'h00000000} /* (6, 3, 25) {real, imag} */,
  {32'h45eee7c6, 32'h00000000} /* (6, 3, 24) {real, imag} */,
  {32'h45c8820e, 32'h00000000} /* (6, 3, 23) {real, imag} */,
  {32'h45c4c844, 32'h00000000} /* (6, 3, 22) {real, imag} */,
  {32'h45aa354b, 32'h00000000} /* (6, 3, 21) {real, imag} */,
  {32'h458c026f, 32'h00000000} /* (6, 3, 20) {real, imag} */,
  {32'h4573b6df, 32'h00000000} /* (6, 3, 19) {real, imag} */,
  {32'h454b0d98, 32'h00000000} /* (6, 3, 18) {real, imag} */,
  {32'h44f5c806, 32'h00000000} /* (6, 3, 17) {real, imag} */,
  {32'h439f2ab0, 32'h00000000} /* (6, 3, 16) {real, imag} */,
  {32'hc4a330e4, 32'h00000000} /* (6, 3, 15) {real, imag} */,
  {32'hc55d5ff5, 32'h00000000} /* (6, 3, 14) {real, imag} */,
  {32'hc5291c78, 32'h00000000} /* (6, 3, 13) {real, imag} */,
  {32'hc556534a, 32'h00000000} /* (6, 3, 12) {real, imag} */,
  {32'hc54827b8, 32'h00000000} /* (6, 3, 11) {real, imag} */,
  {32'hc5077330, 32'h00000000} /* (6, 3, 10) {real, imag} */,
  {32'hc5188806, 32'h00000000} /* (6, 3, 9) {real, imag} */,
  {32'hc4a34260, 32'h00000000} /* (6, 3, 8) {real, imag} */,
  {32'hc38c14a8, 32'h00000000} /* (6, 3, 7) {real, imag} */,
  {32'h4355f310, 32'h00000000} /* (6, 3, 6) {real, imag} */,
  {32'h4510b8ea, 32'h00000000} /* (6, 3, 5) {real, imag} */,
  {32'h45939649, 32'h00000000} /* (6, 3, 4) {real, imag} */,
  {32'h45af5b5e, 32'h00000000} /* (6, 3, 3) {real, imag} */,
  {32'h45af8bf6, 32'h00000000} /* (6, 3, 2) {real, imag} */,
  {32'h45e19fa6, 32'h00000000} /* (6, 3, 1) {real, imag} */,
  {32'h45e4fddf, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'h45dad18e, 32'h00000000} /* (6, 2, 31) {real, imag} */,
  {32'h45f9445c, 32'h00000000} /* (6, 2, 30) {real, imag} */,
  {32'h45e3ff02, 32'h00000000} /* (6, 2, 29) {real, imag} */,
  {32'h45fda5f0, 32'h00000000} /* (6, 2, 28) {real, imag} */,
  {32'h45fb848c, 32'h00000000} /* (6, 2, 27) {real, imag} */,
  {32'h45d36033, 32'h00000000} /* (6, 2, 26) {real, imag} */,
  {32'h45fd03c1, 32'h00000000} /* (6, 2, 25) {real, imag} */,
  {32'h45f7710b, 32'h00000000} /* (6, 2, 24) {real, imag} */,
  {32'h45c90e20, 32'h00000000} /* (6, 2, 23) {real, imag} */,
  {32'h45f71893, 32'h00000000} /* (6, 2, 22) {real, imag} */,
  {32'h45c28b5f, 32'h00000000} /* (6, 2, 21) {real, imag} */,
  {32'h45a2cb60, 32'h00000000} /* (6, 2, 20) {real, imag} */,
  {32'h4583950f, 32'h00000000} /* (6, 2, 19) {real, imag} */,
  {32'h454ed874, 32'h00000000} /* (6, 2, 18) {real, imag} */,
  {32'h453b791b, 32'h00000000} /* (6, 2, 17) {real, imag} */,
  {32'h44b76e48, 32'h00000000} /* (6, 2, 16) {real, imag} */,
  {32'hc44489ac, 32'h00000000} /* (6, 2, 15) {real, imag} */,
  {32'hc5009c43, 32'h00000000} /* (6, 2, 14) {real, imag} */,
  {32'hc4fc6270, 32'h00000000} /* (6, 2, 13) {real, imag} */,
  {32'hc521d218, 32'h00000000} /* (6, 2, 12) {real, imag} */,
  {32'hc52d0390, 32'h00000000} /* (6, 2, 11) {real, imag} */,
  {32'hc5200f7a, 32'h00000000} /* (6, 2, 10) {real, imag} */,
  {32'hc47257d8, 32'h00000000} /* (6, 2, 9) {real, imag} */,
  {32'hc49102cc, 32'h00000000} /* (6, 2, 8) {real, imag} */,
  {32'hc3c55080, 32'h00000000} /* (6, 2, 7) {real, imag} */,
  {32'h448a0f24, 32'h00000000} /* (6, 2, 6) {real, imag} */,
  {32'h4536fb2a, 32'h00000000} /* (6, 2, 5) {real, imag} */,
  {32'h456d4181, 32'h00000000} /* (6, 2, 4) {real, imag} */,
  {32'h45b2a42d, 32'h00000000} /* (6, 2, 3) {real, imag} */,
  {32'h45dc1376, 32'h00000000} /* (6, 2, 2) {real, imag} */,
  {32'h45cd0310, 32'h00000000} /* (6, 2, 1) {real, imag} */,
  {32'h45e7f916, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'h45dbaa5a, 32'h00000000} /* (6, 1, 31) {real, imag} */,
  {32'h45e5733e, 32'h00000000} /* (6, 1, 30) {real, imag} */,
  {32'h45ef9b52, 32'h00000000} /* (6, 1, 29) {real, imag} */,
  {32'h45f5b5b0, 32'h00000000} /* (6, 1, 28) {real, imag} */,
  {32'h45f7d115, 32'h00000000} /* (6, 1, 27) {real, imag} */,
  {32'h45e0fb60, 32'h00000000} /* (6, 1, 26) {real, imag} */,
  {32'h45e69641, 32'h00000000} /* (6, 1, 25) {real, imag} */,
  {32'h45d2cd00, 32'h00000000} /* (6, 1, 24) {real, imag} */,
  {32'h45c2bd46, 32'h00000000} /* (6, 1, 23) {real, imag} */,
  {32'h45b64798, 32'h00000000} /* (6, 1, 22) {real, imag} */,
  {32'h45a5e135, 32'h00000000} /* (6, 1, 21) {real, imag} */,
  {32'h458234f2, 32'h00000000} /* (6, 1, 20) {real, imag} */,
  {32'h452d7fd8, 32'h00000000} /* (6, 1, 19) {real, imag} */,
  {32'h453e2100, 32'h00000000} /* (6, 1, 18) {real, imag} */,
  {32'h4504ea33, 32'h00000000} /* (6, 1, 17) {real, imag} */,
  {32'h44194fd0, 32'h00000000} /* (6, 1, 16) {real, imag} */,
  {32'hc3ff4040, 32'h00000000} /* (6, 1, 15) {real, imag} */,
  {32'hc4341358, 32'h00000000} /* (6, 1, 14) {real, imag} */,
  {32'hc509a3c5, 32'h00000000} /* (6, 1, 13) {real, imag} */,
  {32'hc514e473, 32'h00000000} /* (6, 1, 12) {real, imag} */,
  {32'hc52d8aa6, 32'h00000000} /* (6, 1, 11) {real, imag} */,
  {32'hc4eea398, 32'h00000000} /* (6, 1, 10) {real, imag} */,
  {32'hc48ce66c, 32'h00000000} /* (6, 1, 9) {real, imag} */,
  {32'hc41795a8, 32'h00000000} /* (6, 1, 8) {real, imag} */,
  {32'h4350fc80, 32'h00000000} /* (6, 1, 7) {real, imag} */,
  {32'h448dde0e, 32'h00000000} /* (6, 1, 6) {real, imag} */,
  {32'h454e58e2, 32'h00000000} /* (6, 1, 5) {real, imag} */,
  {32'h4581bdbe, 32'h00000000} /* (6, 1, 4) {real, imag} */,
  {32'h45b10886, 32'h00000000} /* (6, 1, 3) {real, imag} */,
  {32'h45b65cac, 32'h00000000} /* (6, 1, 2) {real, imag} */,
  {32'h45d11746, 32'h00000000} /* (6, 1, 1) {real, imag} */,
  {32'h45d054a1, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'h45e8a6b6, 32'h00000000} /* (6, 0, 31) {real, imag} */,
  {32'h45e9d082, 32'h00000000} /* (6, 0, 30) {real, imag} */,
  {32'h45e62778, 32'h00000000} /* (6, 0, 29) {real, imag} */,
  {32'h45e0f491, 32'h00000000} /* (6, 0, 28) {real, imag} */,
  {32'h460c82a7, 32'h00000000} /* (6, 0, 27) {real, imag} */,
  {32'h45da2cc3, 32'h00000000} /* (6, 0, 26) {real, imag} */,
  {32'h45dbe484, 32'h00000000} /* (6, 0, 25) {real, imag} */,
  {32'h45c48ef2, 32'h00000000} /* (6, 0, 24) {real, imag} */,
  {32'h45ae670c, 32'h00000000} /* (6, 0, 23) {real, imag} */,
  {32'h4593e9c3, 32'h00000000} /* (6, 0, 22) {real, imag} */,
  {32'h45928ed7, 32'h00000000} /* (6, 0, 21) {real, imag} */,
  {32'h45610d18, 32'h00000000} /* (6, 0, 20) {real, imag} */,
  {32'h45090a40, 32'h00000000} /* (6, 0, 19) {real, imag} */,
  {32'h44c976de, 32'h00000000} /* (6, 0, 18) {real, imag} */,
  {32'h443dc9f4, 32'h00000000} /* (6, 0, 17) {real, imag} */,
  {32'hc31ba3b0, 32'h00000000} /* (6, 0, 16) {real, imag} */,
  {32'hc494c9b8, 32'h00000000} /* (6, 0, 15) {real, imag} */,
  {32'hc49235ae, 32'h00000000} /* (6, 0, 14) {real, imag} */,
  {32'hc5021ef7, 32'h00000000} /* (6, 0, 13) {real, imag} */,
  {32'hc51b3a32, 32'h00000000} /* (6, 0, 12) {real, imag} */,
  {32'hc4c5cf40, 32'h00000000} /* (6, 0, 11) {real, imag} */,
  {32'hc45b0058, 32'h00000000} /* (6, 0, 10) {real, imag} */,
  {32'hc3b2d5f0, 32'h00000000} /* (6, 0, 9) {real, imag} */,
  {32'h43db7158, 32'h00000000} /* (6, 0, 8) {real, imag} */,
  {32'h4487cfba, 32'h00000000} /* (6, 0, 7) {real, imag} */,
  {32'h44f521f7, 32'h00000000} /* (6, 0, 6) {real, imag} */,
  {32'h456d26f2, 32'h00000000} /* (6, 0, 5) {real, imag} */,
  {32'h459f46a8, 32'h00000000} /* (6, 0, 4) {real, imag} */,
  {32'h45afe808, 32'h00000000} /* (6, 0, 3) {real, imag} */,
  {32'h45bdfb80, 32'h00000000} /* (6, 0, 2) {real, imag} */,
  {32'h45c62e9e, 32'h00000000} /* (6, 0, 1) {real, imag} */,
  {32'h45d228aa, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'h45848ef2, 32'h00000000} /* (5, 31, 31) {real, imag} */,
  {32'h458db585, 32'h00000000} /* (5, 31, 30) {real, imag} */,
  {32'h4588616c, 32'h00000000} /* (5, 31, 29) {real, imag} */,
  {32'h45853928, 32'h00000000} /* (5, 31, 28) {real, imag} */,
  {32'h4575bf8e, 32'h00000000} /* (5, 31, 27) {real, imag} */,
  {32'h454f53ec, 32'h00000000} /* (5, 31, 26) {real, imag} */,
  {32'h455c4ec9, 32'h00000000} /* (5, 31, 25) {real, imag} */,
  {32'h45315df8, 32'h00000000} /* (5, 31, 24) {real, imag} */,
  {32'h451d88a8, 32'h00000000} /* (5, 31, 23) {real, imag} */,
  {32'h4510f020, 32'h00000000} /* (5, 31, 22) {real, imag} */,
  {32'h450f152e, 32'h00000000} /* (5, 31, 21) {real, imag} */,
  {32'h4498d052, 32'h00000000} /* (5, 31, 20) {real, imag} */,
  {32'h448e924a, 32'h00000000} /* (5, 31, 19) {real, imag} */,
  {32'h44921b34, 32'h00000000} /* (5, 31, 18) {real, imag} */,
  {32'h433dabb0, 32'h00000000} /* (5, 31, 17) {real, imag} */,
  {32'h4372d1c8, 32'h00000000} /* (5, 31, 16) {real, imag} */,
  {32'h43986710, 32'h00000000} /* (5, 31, 15) {real, imag} */,
  {32'hc416b4b6, 32'h00000000} /* (5, 31, 14) {real, imag} */,
  {32'h4388ff00, 32'h00000000} /* (5, 31, 13) {real, imag} */,
  {32'h43424c90, 32'h00000000} /* (5, 31, 12) {real, imag} */,
  {32'h43d31410, 32'h00000000} /* (5, 31, 11) {real, imag} */,
  {32'h446c7446, 32'h00000000} /* (5, 31, 10) {real, imag} */,
  {32'h442114bc, 32'h00000000} /* (5, 31, 9) {real, imag} */,
  {32'h4468278c, 32'h00000000} /* (5, 31, 8) {real, imag} */,
  {32'h44c2100c, 32'h00000000} /* (5, 31, 7) {real, imag} */,
  {32'h44d61b5b, 32'h00000000} /* (5, 31, 6) {real, imag} */,
  {32'h44f90c6c, 32'h00000000} /* (5, 31, 5) {real, imag} */,
  {32'h4500c7ee, 32'h00000000} /* (5, 31, 4) {real, imag} */,
  {32'h44f86de0, 32'h00000000} /* (5, 31, 3) {real, imag} */,
  {32'h452e0928, 32'h00000000} /* (5, 31, 2) {real, imag} */,
  {32'h457a8101, 32'h00000000} /* (5, 31, 1) {real, imag} */,
  {32'h4587268a, 32'h00000000} /* (5, 31, 0) {real, imag} */,
  {32'h4584e8b4, 32'h00000000} /* (5, 30, 31) {real, imag} */,
  {32'h4599b7a0, 32'h00000000} /* (5, 30, 30) {real, imag} */,
  {32'h4592c6ec, 32'h00000000} /* (5, 30, 29) {real, imag} */,
  {32'h45738dd6, 32'h00000000} /* (5, 30, 28) {real, imag} */,
  {32'h457b6667, 32'h00000000} /* (5, 30, 27) {real, imag} */,
  {32'h45326c6c, 32'h00000000} /* (5, 30, 26) {real, imag} */,
  {32'h451e126a, 32'h00000000} /* (5, 30, 25) {real, imag} */,
  {32'h453946a3, 32'h00000000} /* (5, 30, 24) {real, imag} */,
  {32'h452bab89, 32'h00000000} /* (5, 30, 23) {real, imag} */,
  {32'h449ec8b6, 32'h00000000} /* (5, 30, 22) {real, imag} */,
  {32'h4525aac9, 32'h00000000} /* (5, 30, 21) {real, imag} */,
  {32'h4509c5a6, 32'h00000000} /* (5, 30, 20) {real, imag} */,
  {32'h4449e460, 32'h00000000} /* (5, 30, 19) {real, imag} */,
  {32'h444b51ac, 32'h00000000} /* (5, 30, 18) {real, imag} */,
  {32'h4498160c, 32'h00000000} /* (5, 30, 17) {real, imag} */,
  {32'h440561ac, 32'h00000000} /* (5, 30, 16) {real, imag} */,
  {32'h43c8fa2c, 32'h00000000} /* (5, 30, 15) {real, imag} */,
  {32'hc2f24b00, 32'h00000000} /* (5, 30, 14) {real, imag} */,
  {32'hc2f03380, 32'h00000000} /* (5, 30, 13) {real, imag} */,
  {32'h43eafa90, 32'h00000000} /* (5, 30, 12) {real, imag} */,
  {32'h441b277c, 32'h00000000} /* (5, 30, 11) {real, imag} */,
  {32'h4409c40c, 32'h00000000} /* (5, 30, 10) {real, imag} */,
  {32'h43fb844c, 32'h00000000} /* (5, 30, 9) {real, imag} */,
  {32'h44ad56f6, 32'h00000000} /* (5, 30, 8) {real, imag} */,
  {32'h450d8c59, 32'h00000000} /* (5, 30, 7) {real, imag} */,
  {32'h4419c7cb, 32'h00000000} /* (5, 30, 6) {real, imag} */,
  {32'h44565943, 32'h00000000} /* (5, 30, 5) {real, imag} */,
  {32'h44f95014, 32'h00000000} /* (5, 30, 4) {real, imag} */,
  {32'h453ffbd2, 32'h00000000} /* (5, 30, 3) {real, imag} */,
  {32'h456f30d5, 32'h00000000} /* (5, 30, 2) {real, imag} */,
  {32'h4587b15f, 32'h00000000} /* (5, 30, 1) {real, imag} */,
  {32'h458eb610, 32'h00000000} /* (5, 30, 0) {real, imag} */,
  {32'h458f578a, 32'h00000000} /* (5, 29, 31) {real, imag} */,
  {32'h458058a3, 32'h00000000} /* (5, 29, 30) {real, imag} */,
  {32'h45188298, 32'h00000000} /* (5, 29, 29) {real, imag} */,
  {32'h4576be89, 32'h00000000} /* (5, 29, 28) {real, imag} */,
  {32'h454783a7, 32'h00000000} /* (5, 29, 27) {real, imag} */,
  {32'h44f86326, 32'h00000000} /* (5, 29, 26) {real, imag} */,
  {32'h44aeb021, 32'h00000000} /* (5, 29, 25) {real, imag} */,
  {32'h4529449a, 32'h00000000} /* (5, 29, 24) {real, imag} */,
  {32'h44e2fd0e, 32'h00000000} /* (5, 29, 23) {real, imag} */,
  {32'h44ebb7e2, 32'h00000000} /* (5, 29, 22) {real, imag} */,
  {32'h4510ebd6, 32'h00000000} /* (5, 29, 21) {real, imag} */,
  {32'h44969a17, 32'h00000000} /* (5, 29, 20) {real, imag} */,
  {32'h442f8e90, 32'h00000000} /* (5, 29, 19) {real, imag} */,
  {32'h43567b80, 32'h00000000} /* (5, 29, 18) {real, imag} */,
  {32'h4449ce2a, 32'h00000000} /* (5, 29, 17) {real, imag} */,
  {32'h4401f680, 32'h00000000} /* (5, 29, 16) {real, imag} */,
  {32'h43bfedc0, 32'h00000000} /* (5, 29, 15) {real, imag} */,
  {32'h43ab70f0, 32'h00000000} /* (5, 29, 14) {real, imag} */,
  {32'h4350bf60, 32'h00000000} /* (5, 29, 13) {real, imag} */,
  {32'h440d24ac, 32'h00000000} /* (5, 29, 12) {real, imag} */,
  {32'h430efb60, 32'h00000000} /* (5, 29, 11) {real, imag} */,
  {32'h430bc550, 32'h00000000} /* (5, 29, 10) {real, imag} */,
  {32'h438f6f24, 32'h00000000} /* (5, 29, 9) {real, imag} */,
  {32'h45124b8e, 32'h00000000} /* (5, 29, 8) {real, imag} */,
  {32'h4511f235, 32'h00000000} /* (5, 29, 7) {real, imag} */,
  {32'h44132a5c, 32'h00000000} /* (5, 29, 6) {real, imag} */,
  {32'h44da7cfc, 32'h00000000} /* (5, 29, 5) {real, imag} */,
  {32'h44e58a8b, 32'h00000000} /* (5, 29, 4) {real, imag} */,
  {32'h455f4c5c, 32'h00000000} /* (5, 29, 3) {real, imag} */,
  {32'h4564dfd4, 32'h00000000} /* (5, 29, 2) {real, imag} */,
  {32'h4583492f, 32'h00000000} /* (5, 29, 1) {real, imag} */,
  {32'h458418bc, 32'h00000000} /* (5, 29, 0) {real, imag} */,
  {32'h45850086, 32'h00000000} /* (5, 28, 31) {real, imag} */,
  {32'h4529d6ba, 32'h00000000} /* (5, 28, 30) {real, imag} */,
  {32'h452f5266, 32'h00000000} /* (5, 28, 29) {real, imag} */,
  {32'h455879ca, 32'h00000000} /* (5, 28, 28) {real, imag} */,
  {32'h4538d23a, 32'h00000000} /* (5, 28, 27) {real, imag} */,
  {32'h44c9c314, 32'h00000000} /* (5, 28, 26) {real, imag} */,
  {32'h44d8d93e, 32'h00000000} /* (5, 28, 25) {real, imag} */,
  {32'h452bf30d, 32'h00000000} /* (5, 28, 24) {real, imag} */,
  {32'h44cbfb36, 32'h00000000} /* (5, 28, 23) {real, imag} */,
  {32'h44ffd1e8, 32'h00000000} /* (5, 28, 22) {real, imag} */,
  {32'h451d7d70, 32'h00000000} /* (5, 28, 21) {real, imag} */,
  {32'h449594d1, 32'h00000000} /* (5, 28, 20) {real, imag} */,
  {32'h441238ec, 32'h00000000} /* (5, 28, 19) {real, imag} */,
  {32'h442af718, 32'h00000000} /* (5, 28, 18) {real, imag} */,
  {32'h43d273a8, 32'h00000000} /* (5, 28, 17) {real, imag} */,
  {32'h43ba023c, 32'h00000000} /* (5, 28, 16) {real, imag} */,
  {32'h438e6428, 32'h00000000} /* (5, 28, 15) {real, imag} */,
  {32'hc2a2b360, 32'h00000000} /* (5, 28, 14) {real, imag} */,
  {32'h43d9360c, 32'h00000000} /* (5, 28, 13) {real, imag} */,
  {32'h44ad8ba7, 32'h00000000} /* (5, 28, 12) {real, imag} */,
  {32'h44809406, 32'h00000000} /* (5, 28, 11) {real, imag} */,
  {32'h4522e35a, 32'h00000000} /* (5, 28, 10) {real, imag} */,
  {32'h448f5e56, 32'h00000000} /* (5, 28, 9) {real, imag} */,
  {32'h445c32e0, 32'h00000000} /* (5, 28, 8) {real, imag} */,
  {32'h44903bd8, 32'h00000000} /* (5, 28, 7) {real, imag} */,
  {32'h44dfc956, 32'h00000000} /* (5, 28, 6) {real, imag} */,
  {32'h4504dfe8, 32'h00000000} /* (5, 28, 5) {real, imag} */,
  {32'h4547cfee, 32'h00000000} /* (5, 28, 4) {real, imag} */,
  {32'h4529cfc6, 32'h00000000} /* (5, 28, 3) {real, imag} */,
  {32'h45460bf8, 32'h00000000} /* (5, 28, 2) {real, imag} */,
  {32'h4559f0b7, 32'h00000000} /* (5, 28, 1) {real, imag} */,
  {32'h455e2cf8, 32'h00000000} /* (5, 28, 0) {real, imag} */,
  {32'h455ba7c4, 32'h00000000} /* (5, 27, 31) {real, imag} */,
  {32'h4528e284, 32'h00000000} /* (5, 27, 30) {real, imag} */,
  {32'h4554d7b3, 32'h00000000} /* (5, 27, 29) {real, imag} */,
  {32'h451e975e, 32'h00000000} /* (5, 27, 28) {real, imag} */,
  {32'h44c8bc2e, 32'h00000000} /* (5, 27, 27) {real, imag} */,
  {32'h451a8f2b, 32'h00000000} /* (5, 27, 26) {real, imag} */,
  {32'h44ccf30c, 32'h00000000} /* (5, 27, 25) {real, imag} */,
  {32'h43099a34, 32'h00000000} /* (5, 27, 24) {real, imag} */,
  {32'h44a69f1c, 32'h00000000} /* (5, 27, 23) {real, imag} */,
  {32'h44dd234c, 32'h00000000} /* (5, 27, 22) {real, imag} */,
  {32'h450cd8b7, 32'h00000000} /* (5, 27, 21) {real, imag} */,
  {32'h44e752a9, 32'h00000000} /* (5, 27, 20) {real, imag} */,
  {32'h44995827, 32'h00000000} /* (5, 27, 19) {real, imag} */,
  {32'h440074a8, 32'h00000000} /* (5, 27, 18) {real, imag} */,
  {32'h43e5c934, 32'h00000000} /* (5, 27, 17) {real, imag} */,
  {32'h43dce928, 32'h00000000} /* (5, 27, 16) {real, imag} */,
  {32'h44106788, 32'h00000000} /* (5, 27, 15) {real, imag} */,
  {32'hc3409108, 32'h00000000} /* (5, 27, 14) {real, imag} */,
  {32'h4450379c, 32'h00000000} /* (5, 27, 13) {real, imag} */,
  {32'h444f52f5, 32'h00000000} /* (5, 27, 12) {real, imag} */,
  {32'h45045e9a, 32'h00000000} /* (5, 27, 11) {real, imag} */,
  {32'h44cf93b2, 32'h00000000} /* (5, 27, 10) {real, imag} */,
  {32'h44e0ac3e, 32'h00000000} /* (5, 27, 9) {real, imag} */,
  {32'h44efe77a, 32'h00000000} /* (5, 27, 8) {real, imag} */,
  {32'h45036b2a, 32'h00000000} /* (5, 27, 7) {real, imag} */,
  {32'h4519958a, 32'h00000000} /* (5, 27, 6) {real, imag} */,
  {32'h4519080b, 32'h00000000} /* (5, 27, 5) {real, imag} */,
  {32'h45215853, 32'h00000000} /* (5, 27, 4) {real, imag} */,
  {32'h4513b352, 32'h00000000} /* (5, 27, 3) {real, imag} */,
  {32'h45316dff, 32'h00000000} /* (5, 27, 2) {real, imag} */,
  {32'h4543cdfc, 32'h00000000} /* (5, 27, 1) {real, imag} */,
  {32'h4520e2d1, 32'h00000000} /* (5, 27, 0) {real, imag} */,
  {32'h453ae44c, 32'h00000000} /* (5, 26, 31) {real, imag} */,
  {32'h4549b81e, 32'h00000000} /* (5, 26, 30) {real, imag} */,
  {32'h451ea4ca, 32'h00000000} /* (5, 26, 29) {real, imag} */,
  {32'h45172ddd, 32'h00000000} /* (5, 26, 28) {real, imag} */,
  {32'h4527e898, 32'h00000000} /* (5, 26, 27) {real, imag} */,
  {32'h452c7064, 32'h00000000} /* (5, 26, 26) {real, imag} */,
  {32'h44bc0248, 32'h00000000} /* (5, 26, 25) {real, imag} */,
  {32'h441c2754, 32'h00000000} /* (5, 26, 24) {real, imag} */,
  {32'h449571a6, 32'h00000000} /* (5, 26, 23) {real, imag} */,
  {32'h44b53eec, 32'h00000000} /* (5, 26, 22) {real, imag} */,
  {32'h448e1c86, 32'h00000000} /* (5, 26, 21) {real, imag} */,
  {32'h44c5b01f, 32'h00000000} /* (5, 26, 20) {real, imag} */,
  {32'h449869e1, 32'h00000000} /* (5, 26, 19) {real, imag} */,
  {32'h44c9d32a, 32'h00000000} /* (5, 26, 18) {real, imag} */,
  {32'h438bf0e0, 32'h00000000} /* (5, 26, 17) {real, imag} */,
  {32'h431dcd28, 32'h00000000} /* (5, 26, 16) {real, imag} */,
  {32'h448b6208, 32'h00000000} /* (5, 26, 15) {real, imag} */,
  {32'h444287a2, 32'h00000000} /* (5, 26, 14) {real, imag} */,
  {32'h423199a0, 32'h00000000} /* (5, 26, 13) {real, imag} */,
  {32'h448b198e, 32'h00000000} /* (5, 26, 12) {real, imag} */,
  {32'h4436117c, 32'h00000000} /* (5, 26, 11) {real, imag} */,
  {32'h44095e70, 32'h00000000} /* (5, 26, 10) {real, imag} */,
  {32'h44d38bd0, 32'h00000000} /* (5, 26, 9) {real, imag} */,
  {32'h4515f68a, 32'h00000000} /* (5, 26, 8) {real, imag} */,
  {32'h4512c6df, 32'h00000000} /* (5, 26, 7) {real, imag} */,
  {32'h451ee5cb, 32'h00000000} /* (5, 26, 6) {real, imag} */,
  {32'h450f0551, 32'h00000000} /* (5, 26, 5) {real, imag} */,
  {32'h4527b5b4, 32'h00000000} /* (5, 26, 4) {real, imag} */,
  {32'h451523ae, 32'h00000000} /* (5, 26, 3) {real, imag} */,
  {32'h45363cbf, 32'h00000000} /* (5, 26, 2) {real, imag} */,
  {32'h454414e4, 32'h00000000} /* (5, 26, 1) {real, imag} */,
  {32'h4516c022, 32'h00000000} /* (5, 26, 0) {real, imag} */,
  {32'h4521d28c, 32'h00000000} /* (5, 25, 31) {real, imag} */,
  {32'h44ccf7c6, 32'h00000000} /* (5, 25, 30) {real, imag} */,
  {32'h44f86e9a, 32'h00000000} /* (5, 25, 29) {real, imag} */,
  {32'h45064ad0, 32'h00000000} /* (5, 25, 28) {real, imag} */,
  {32'h45180e8d, 32'h00000000} /* (5, 25, 27) {real, imag} */,
  {32'h44df8c5f, 32'h00000000} /* (5, 25, 26) {real, imag} */,
  {32'h44af50be, 32'h00000000} /* (5, 25, 25) {real, imag} */,
  {32'h4408ffa6, 32'h00000000} /* (5, 25, 24) {real, imag} */,
  {32'h448d4199, 32'h00000000} /* (5, 25, 23) {real, imag} */,
  {32'h4478f8b5, 32'h00000000} /* (5, 25, 22) {real, imag} */,
  {32'h442f59d0, 32'h00000000} /* (5, 25, 21) {real, imag} */,
  {32'h450c676b, 32'h00000000} /* (5, 25, 20) {real, imag} */,
  {32'h44e120a0, 32'h00000000} /* (5, 25, 19) {real, imag} */,
  {32'h4489f9b0, 32'h00000000} /* (5, 25, 18) {real, imag} */,
  {32'h44d52f1e, 32'h00000000} /* (5, 25, 17) {real, imag} */,
  {32'h44124a01, 32'h00000000} /* (5, 25, 16) {real, imag} */,
  {32'h44984c30, 32'h00000000} /* (5, 25, 15) {real, imag} */,
  {32'h44987f52, 32'h00000000} /* (5, 25, 14) {real, imag} */,
  {32'hc2062af0, 32'h00000000} /* (5, 25, 13) {real, imag} */,
  {32'h44945e3d, 32'h00000000} /* (5, 25, 12) {real, imag} */,
  {32'h449bf4c4, 32'h00000000} /* (5, 25, 11) {real, imag} */,
  {32'h44730576, 32'h00000000} /* (5, 25, 10) {real, imag} */,
  {32'h44a8fe0a, 32'h00000000} /* (5, 25, 9) {real, imag} */,
  {32'h44347a78, 32'h00000000} /* (5, 25, 8) {real, imag} */,
  {32'h44c74b0b, 32'h00000000} /* (5, 25, 7) {real, imag} */,
  {32'h4516117b, 32'h00000000} /* (5, 25, 6) {real, imag} */,
  {32'h45326038, 32'h00000000} /* (5, 25, 5) {real, imag} */,
  {32'h45119131, 32'h00000000} /* (5, 25, 4) {real, imag} */,
  {32'h44b94eb6, 32'h00000000} /* (5, 25, 3) {real, imag} */,
  {32'h44a4ad7e, 32'h00000000} /* (5, 25, 2) {real, imag} */,
  {32'h4521628f, 32'h00000000} /* (5, 25, 1) {real, imag} */,
  {32'h4509e744, 32'h00000000} /* (5, 25, 0) {real, imag} */,
  {32'h44f3806c, 32'h00000000} /* (5, 24, 31) {real, imag} */,
  {32'h451ba292, 32'h00000000} /* (5, 24, 30) {real, imag} */,
  {32'h44b0ba6a, 32'h00000000} /* (5, 24, 29) {real, imag} */,
  {32'h44e1f140, 32'h00000000} /* (5, 24, 28) {real, imag} */,
  {32'h4466841f, 32'h00000000} /* (5, 24, 27) {real, imag} */,
  {32'h44abeef2, 32'h00000000} /* (5, 24, 26) {real, imag} */,
  {32'h44b7b1d8, 32'h00000000} /* (5, 24, 25) {real, imag} */,
  {32'h449e220c, 32'h00000000} /* (5, 24, 24) {real, imag} */,
  {32'h44a357ad, 32'h00000000} /* (5, 24, 23) {real, imag} */,
  {32'h447f9cd0, 32'h00000000} /* (5, 24, 22) {real, imag} */,
  {32'h44e18655, 32'h00000000} /* (5, 24, 21) {real, imag} */,
  {32'h450fb5ac, 32'h00000000} /* (5, 24, 20) {real, imag} */,
  {32'h450479ea, 32'h00000000} /* (5, 24, 19) {real, imag} */,
  {32'h44a53ce1, 32'h00000000} /* (5, 24, 18) {real, imag} */,
  {32'h44627bda, 32'h00000000} /* (5, 24, 17) {real, imag} */,
  {32'h447d4564, 32'h00000000} /* (5, 24, 16) {real, imag} */,
  {32'h441672ef, 32'h00000000} /* (5, 24, 15) {real, imag} */,
  {32'hc2a367d0, 32'h00000000} /* (5, 24, 14) {real, imag} */,
  {32'h4455ceaf, 32'h00000000} /* (5, 24, 13) {real, imag} */,
  {32'h43bea30e, 32'h00000000} /* (5, 24, 12) {real, imag} */,
  {32'h44edb5f6, 32'h00000000} /* (5, 24, 11) {real, imag} */,
  {32'h44cf2bae, 32'h00000000} /* (5, 24, 10) {real, imag} */,
  {32'h4407ac19, 32'h00000000} /* (5, 24, 9) {real, imag} */,
  {32'h443b2153, 32'h00000000} /* (5, 24, 8) {real, imag} */,
  {32'h44ad5673, 32'h00000000} /* (5, 24, 7) {real, imag} */,
  {32'h44f4e27c, 32'h00000000} /* (5, 24, 6) {real, imag} */,
  {32'h44e7b8c1, 32'h00000000} /* (5, 24, 5) {real, imag} */,
  {32'h44e6f508, 32'h00000000} /* (5, 24, 4) {real, imag} */,
  {32'h44e80742, 32'h00000000} /* (5, 24, 3) {real, imag} */,
  {32'h4401d2d6, 32'h00000000} /* (5, 24, 2) {real, imag} */,
  {32'h451b25e4, 32'h00000000} /* (5, 24, 1) {real, imag} */,
  {32'h44e8420c, 32'h00000000} /* (5, 24, 0) {real, imag} */,
  {32'h44a9f394, 32'h00000000} /* (5, 23, 31) {real, imag} */,
  {32'h450d2173, 32'h00000000} /* (5, 23, 30) {real, imag} */,
  {32'h44a23772, 32'h00000000} /* (5, 23, 29) {real, imag} */,
  {32'h44b57a95, 32'h00000000} /* (5, 23, 28) {real, imag} */,
  {32'h4485e9b6, 32'h00000000} /* (5, 23, 27) {real, imag} */,
  {32'h449c47b3, 32'h00000000} /* (5, 23, 26) {real, imag} */,
  {32'h44cd60eb, 32'h00000000} /* (5, 23, 25) {real, imag} */,
  {32'h44e8aa61, 32'h00000000} /* (5, 23, 24) {real, imag} */,
  {32'h447d67f6, 32'h00000000} /* (5, 23, 23) {real, imag} */,
  {32'h441ed6f6, 32'h00000000} /* (5, 23, 22) {real, imag} */,
  {32'h4501b107, 32'h00000000} /* (5, 23, 21) {real, imag} */,
  {32'h44cd692a, 32'h00000000} /* (5, 23, 20) {real, imag} */,
  {32'h44efed49, 32'h00000000} /* (5, 23, 19) {real, imag} */,
  {32'h45029d0f, 32'h00000000} /* (5, 23, 18) {real, imag} */,
  {32'h44e28bb6, 32'h00000000} /* (5, 23, 17) {real, imag} */,
  {32'h44784fb6, 32'h00000000} /* (5, 23, 16) {real, imag} */,
  {32'h449922f6, 32'h00000000} /* (5, 23, 15) {real, imag} */,
  {32'h446f0f39, 32'h00000000} /* (5, 23, 14) {real, imag} */,
  {32'h441212ae, 32'h00000000} /* (5, 23, 13) {real, imag} */,
  {32'h4464b36a, 32'h00000000} /* (5, 23, 12) {real, imag} */,
  {32'h4419ebdf, 32'h00000000} /* (5, 23, 11) {real, imag} */,
  {32'h4446f52e, 32'h00000000} /* (5, 23, 10) {real, imag} */,
  {32'h43c9d598, 32'h00000000} /* (5, 23, 9) {real, imag} */,
  {32'h442f0c96, 32'h00000000} /* (5, 23, 8) {real, imag} */,
  {32'h4440f128, 32'h00000000} /* (5, 23, 7) {real, imag} */,
  {32'h445a3236, 32'h00000000} /* (5, 23, 6) {real, imag} */,
  {32'h44627b7b, 32'h00000000} /* (5, 23, 5) {real, imag} */,
  {32'h44a0197c, 32'h00000000} /* (5, 23, 4) {real, imag} */,
  {32'h4442dee2, 32'h00000000} /* (5, 23, 3) {real, imag} */,
  {32'h43993b80, 32'h00000000} /* (5, 23, 2) {real, imag} */,
  {32'h445f16dd, 32'h00000000} /* (5, 23, 1) {real, imag} */,
  {32'h448b2529, 32'h00000000} /* (5, 23, 0) {real, imag} */,
  {32'h4430c1bc, 32'h00000000} /* (5, 22, 31) {real, imag} */,
  {32'h4477d4ac, 32'h00000000} /* (5, 22, 30) {real, imag} */,
  {32'h44661968, 32'h00000000} /* (5, 22, 29) {real, imag} */,
  {32'h44322939, 32'h00000000} /* (5, 22, 28) {real, imag} */,
  {32'h44cd2e51, 32'h00000000} /* (5, 22, 27) {real, imag} */,
  {32'h44ad918f, 32'h00000000} /* (5, 22, 26) {real, imag} */,
  {32'h449e1a45, 32'h00000000} /* (5, 22, 25) {real, imag} */,
  {32'h43d9e176, 32'h00000000} /* (5, 22, 24) {real, imag} */,
  {32'h44869344, 32'h00000000} /* (5, 22, 23) {real, imag} */,
  {32'h447a87f4, 32'h00000000} /* (5, 22, 22) {real, imag} */,
  {32'h4470af74, 32'h00000000} /* (5, 22, 21) {real, imag} */,
  {32'h44f28d09, 32'h00000000} /* (5, 22, 20) {real, imag} */,
  {32'h4529f7fa, 32'h00000000} /* (5, 22, 19) {real, imag} */,
  {32'h45189706, 32'h00000000} /* (5, 22, 18) {real, imag} */,
  {32'h4481abae, 32'h00000000} /* (5, 22, 17) {real, imag} */,
  {32'h448c5cdc, 32'h00000000} /* (5, 22, 16) {real, imag} */,
  {32'h4421e962, 32'h00000000} /* (5, 22, 15) {real, imag} */,
  {32'h43731c52, 32'h00000000} /* (5, 22, 14) {real, imag} */,
  {32'h4430368a, 32'h00000000} /* (5, 22, 13) {real, imag} */,
  {32'h435ebcc1, 32'h00000000} /* (5, 22, 12) {real, imag} */,
  {32'h443a750e, 32'h00000000} /* (5, 22, 11) {real, imag} */,
  {32'h4400e8c4, 32'h00000000} /* (5, 22, 10) {real, imag} */,
  {32'h44042ca4, 32'h00000000} /* (5, 22, 9) {real, imag} */,
  {32'h42a37c48, 32'h00000000} /* (5, 22, 8) {real, imag} */,
  {32'h4457d2d3, 32'h00000000} /* (5, 22, 7) {real, imag} */,
  {32'h43ac8c91, 32'h00000000} /* (5, 22, 6) {real, imag} */,
  {32'h445870b6, 32'h00000000} /* (5, 22, 5) {real, imag} */,
  {32'h443d2422, 32'h00000000} /* (5, 22, 4) {real, imag} */,
  {32'h421537e0, 32'h00000000} /* (5, 22, 3) {real, imag} */,
  {32'hc34dad48, 32'h00000000} /* (5, 22, 2) {real, imag} */,
  {32'h43f05e56, 32'h00000000} /* (5, 22, 1) {real, imag} */,
  {32'h43f81151, 32'h00000000} /* (5, 22, 0) {real, imag} */,
  {32'h43e70b97, 32'h00000000} /* (5, 21, 31) {real, imag} */,
  {32'h4441181b, 32'h00000000} /* (5, 21, 30) {real, imag} */,
  {32'h446de988, 32'h00000000} /* (5, 21, 29) {real, imag} */,
  {32'h44aa3c59, 32'h00000000} /* (5, 21, 28) {real, imag} */,
  {32'h441b5ad2, 32'h00000000} /* (5, 21, 27) {real, imag} */,
  {32'h4466017c, 32'h00000000} /* (5, 21, 26) {real, imag} */,
  {32'h434ebd1c, 32'h00000000} /* (5, 21, 25) {real, imag} */,
  {32'h4491738a, 32'h00000000} /* (5, 21, 24) {real, imag} */,
  {32'h449e4f81, 32'h00000000} /* (5, 21, 23) {real, imag} */,
  {32'h44873a83, 32'h00000000} /* (5, 21, 22) {real, imag} */,
  {32'h43d3f14c, 32'h00000000} /* (5, 21, 21) {real, imag} */,
  {32'h44cfb370, 32'h00000000} /* (5, 21, 20) {real, imag} */,
  {32'h4523f410, 32'h00000000} /* (5, 21, 19) {real, imag} */,
  {32'h44a9e99e, 32'h00000000} /* (5, 21, 18) {real, imag} */,
  {32'h43f6e106, 32'h00000000} /* (5, 21, 17) {real, imag} */,
  {32'h42e390f8, 32'h00000000} /* (5, 21, 16) {real, imag} */,
  {32'h441797e0, 32'h00000000} /* (5, 21, 15) {real, imag} */,
  {32'h4498fb0e, 32'h00000000} /* (5, 21, 14) {real, imag} */,
  {32'h439e9c65, 32'h00000000} /* (5, 21, 13) {real, imag} */,
  {32'h438142a4, 32'h00000000} /* (5, 21, 12) {real, imag} */,
  {32'h44990c5b, 32'h00000000} /* (5, 21, 11) {real, imag} */,
  {32'h4484ad7a, 32'h00000000} /* (5, 21, 10) {real, imag} */,
  {32'h443e1d1f, 32'h00000000} /* (5, 21, 9) {real, imag} */,
  {32'h44550a87, 32'h00000000} /* (5, 21, 8) {real, imag} */,
  {32'h443bb596, 32'h00000000} /* (5, 21, 7) {real, imag} */,
  {32'h433f36e2, 32'h00000000} /* (5, 21, 6) {real, imag} */,
  {32'h444079d4, 32'h00000000} /* (5, 21, 5) {real, imag} */,
  {32'h4342235c, 32'h00000000} /* (5, 21, 4) {real, imag} */,
  {32'h4402a9e0, 32'h00000000} /* (5, 21, 3) {real, imag} */,
  {32'h438bde50, 32'h00000000} /* (5, 21, 2) {real, imag} */,
  {32'hbea60e00, 32'h00000000} /* (5, 21, 1) {real, imag} */,
  {32'h42df1588, 32'h00000000} /* (5, 21, 0) {real, imag} */,
  {32'h43aa5f81, 32'h00000000} /* (5, 20, 31) {real, imag} */,
  {32'h44d0b148, 32'h00000000} /* (5, 20, 30) {real, imag} */,
  {32'h44872c05, 32'h00000000} /* (5, 20, 29) {real, imag} */,
  {32'h4488651e, 32'h00000000} /* (5, 20, 28) {real, imag} */,
  {32'h44893550, 32'h00000000} /* (5, 20, 27) {real, imag} */,
  {32'hc3bacebc, 32'h00000000} /* (5, 20, 26) {real, imag} */,
  {32'h4433eecf, 32'h00000000} /* (5, 20, 25) {real, imag} */,
  {32'h449a737c, 32'h00000000} /* (5, 20, 24) {real, imag} */,
  {32'h445502cb, 32'h00000000} /* (5, 20, 23) {real, imag} */,
  {32'h447c3a97, 32'h00000000} /* (5, 20, 22) {real, imag} */,
  {32'h44a79ee6, 32'h00000000} /* (5, 20, 21) {real, imag} */,
  {32'h449529a7, 32'h00000000} /* (5, 20, 20) {real, imag} */,
  {32'h448473d6, 32'h00000000} /* (5, 20, 19) {real, imag} */,
  {32'h449ee416, 32'h00000000} /* (5, 20, 18) {real, imag} */,
  {32'h43f6ad1a, 32'h00000000} /* (5, 20, 17) {real, imag} */,
  {32'h4312bbaf, 32'h00000000} /* (5, 20, 16) {real, imag} */,
  {32'h449831f4, 32'h00000000} /* (5, 20, 15) {real, imag} */,
  {32'h4425fb51, 32'h00000000} /* (5, 20, 14) {real, imag} */,
  {32'h41d65180, 32'h00000000} /* (5, 20, 13) {real, imag} */,
  {32'h440d43c0, 32'h00000000} /* (5, 20, 12) {real, imag} */,
  {32'h442c94e1, 32'h00000000} /* (5, 20, 11) {real, imag} */,
  {32'h45023d78, 32'h00000000} /* (5, 20, 10) {real, imag} */,
  {32'h44734f95, 32'h00000000} /* (5, 20, 9) {real, imag} */,
  {32'h433d6814, 32'h00000000} /* (5, 20, 8) {real, imag} */,
  {32'h445bc531, 32'h00000000} /* (5, 20, 7) {real, imag} */,
  {32'h448d7130, 32'h00000000} /* (5, 20, 6) {real, imag} */,
  {32'h44d5727a, 32'h00000000} /* (5, 20, 5) {real, imag} */,
  {32'hc0b55d00, 32'h00000000} /* (5, 20, 4) {real, imag} */,
  {32'h414e0a00, 32'h00000000} /* (5, 20, 3) {real, imag} */,
  {32'h43b3a83a, 32'h00000000} /* (5, 20, 2) {real, imag} */,
  {32'h44223b0f, 32'h00000000} /* (5, 20, 1) {real, imag} */,
  {32'hc194e0f8, 32'h00000000} /* (5, 20, 0) {real, imag} */,
  {32'h42e9ff02, 32'h00000000} /* (5, 19, 31) {real, imag} */,
  {32'h44457e1a, 32'h00000000} /* (5, 19, 30) {real, imag} */,
  {32'hc20d4f20, 32'h00000000} /* (5, 19, 29) {real, imag} */,
  {32'h44680044, 32'h00000000} /* (5, 19, 28) {real, imag} */,
  {32'h440d9821, 32'h00000000} /* (5, 19, 27) {real, imag} */,
  {32'h4217f1a8, 32'h00000000} /* (5, 19, 26) {real, imag} */,
  {32'hc3ed62ec, 32'h00000000} /* (5, 19, 25) {real, imag} */,
  {32'h42b6c60e, 32'h00000000} /* (5, 19, 24) {real, imag} */,
  {32'h440d967e, 32'h00000000} /* (5, 19, 23) {real, imag} */,
  {32'h445e2812, 32'h00000000} /* (5, 19, 22) {real, imag} */,
  {32'h43ebc781, 32'h00000000} /* (5, 19, 21) {real, imag} */,
  {32'h43a47296, 32'h00000000} /* (5, 19, 20) {real, imag} */,
  {32'h4461509c, 32'h00000000} /* (5, 19, 19) {real, imag} */,
  {32'h446bafd0, 32'h00000000} /* (5, 19, 18) {real, imag} */,
  {32'h44197cb5, 32'h00000000} /* (5, 19, 17) {real, imag} */,
  {32'h4385f1e6, 32'h00000000} /* (5, 19, 16) {real, imag} */,
  {32'h437ed99f, 32'h00000000} /* (5, 19, 15) {real, imag} */,
  {32'h43c5536b, 32'h00000000} /* (5, 19, 14) {real, imag} */,
  {32'h44106b10, 32'h00000000} /* (5, 19, 13) {real, imag} */,
  {32'h43b86f78, 32'h00000000} /* (5, 19, 12) {real, imag} */,
  {32'h43974a36, 32'h00000000} /* (5, 19, 11) {real, imag} */,
  {32'h44753d8e, 32'h00000000} /* (5, 19, 10) {real, imag} */,
  {32'h448e15e4, 32'h00000000} /* (5, 19, 9) {real, imag} */,
  {32'hc3783ca5, 32'h00000000} /* (5, 19, 8) {real, imag} */,
  {32'h43b1773c, 32'h00000000} /* (5, 19, 7) {real, imag} */,
  {32'h44034a66, 32'h00000000} /* (5, 19, 6) {real, imag} */,
  {32'h440f3a52, 32'h00000000} /* (5, 19, 5) {real, imag} */,
  {32'h4337daa0, 32'h00000000} /* (5, 19, 4) {real, imag} */,
  {32'hc48b9424, 32'h00000000} /* (5, 19, 3) {real, imag} */,
  {32'hc4021c26, 32'h00000000} /* (5, 19, 2) {real, imag} */,
  {32'hc33ff98c, 32'h00000000} /* (5, 19, 1) {real, imag} */,
  {32'hc4995f90, 32'h00000000} /* (5, 19, 0) {real, imag} */,
  {32'hc3be7f23, 32'h00000000} /* (5, 18, 31) {real, imag} */,
  {32'hc43bf0ce, 32'h00000000} /* (5, 18, 30) {real, imag} */,
  {32'h422e9460, 32'h00000000} /* (5, 18, 29) {real, imag} */,
  {32'h43ad8e9d, 32'h00000000} /* (5, 18, 28) {real, imag} */,
  {32'hc45de714, 32'h00000000} /* (5, 18, 27) {real, imag} */,
  {32'hc0cd6360, 32'h00000000} /* (5, 18, 26) {real, imag} */,
  {32'hc3e7e23e, 32'h00000000} /* (5, 18, 25) {real, imag} */,
  {32'hc424d928, 32'h00000000} /* (5, 18, 24) {real, imag} */,
  {32'hc369025e, 32'h00000000} /* (5, 18, 23) {real, imag} */,
  {32'h43d8a8ea, 32'h00000000} /* (5, 18, 22) {real, imag} */,
  {32'h4401c08f, 32'h00000000} /* (5, 18, 21) {real, imag} */,
  {32'h44923086, 32'h00000000} /* (5, 18, 20) {real, imag} */,
  {32'h443ce5c2, 32'h00000000} /* (5, 18, 19) {real, imag} */,
  {32'h447d9bda, 32'h00000000} /* (5, 18, 18) {real, imag} */,
  {32'h444b4eb8, 32'h00000000} /* (5, 18, 17) {real, imag} */,
  {32'hc3d95cc6, 32'h00000000} /* (5, 18, 16) {real, imag} */,
  {32'h44492466, 32'h00000000} /* (5, 18, 15) {real, imag} */,
  {32'h42cefcd4, 32'h00000000} /* (5, 18, 14) {real, imag} */,
  {32'h4413891e, 32'h00000000} /* (5, 18, 13) {real, imag} */,
  {32'h43a866d1, 32'h00000000} /* (5, 18, 12) {real, imag} */,
  {32'h42355458, 32'h00000000} /* (5, 18, 11) {real, imag} */,
  {32'hc3038f0f, 32'h00000000} /* (5, 18, 10) {real, imag} */,
  {32'hc2bcb552, 32'h00000000} /* (5, 18, 9) {real, imag} */,
  {32'h4325a632, 32'h00000000} /* (5, 18, 8) {real, imag} */,
  {32'h43771ae6, 32'h00000000} /* (5, 18, 7) {real, imag} */,
  {32'h4403cf68, 32'h00000000} /* (5, 18, 6) {real, imag} */,
  {32'h44313ae5, 32'h00000000} /* (5, 18, 5) {real, imag} */,
  {32'hc22dcfa0, 32'h00000000} /* (5, 18, 4) {real, imag} */,
  {32'hc3f2c71c, 32'h00000000} /* (5, 18, 3) {real, imag} */,
  {32'hc4ccff1f, 32'h00000000} /* (5, 18, 2) {real, imag} */,
  {32'hc16ebdc0, 32'h00000000} /* (5, 18, 1) {real, imag} */,
  {32'hc498975c, 32'h00000000} /* (5, 18, 0) {real, imag} */,
  {32'hc491a5b4, 32'h00000000} /* (5, 17, 31) {real, imag} */,
  {32'hc44c0106, 32'h00000000} /* (5, 17, 30) {real, imag} */,
  {32'hc4950a3f, 32'h00000000} /* (5, 17, 29) {real, imag} */,
  {32'hc4b45e29, 32'h00000000} /* (5, 17, 28) {real, imag} */,
  {32'hc468eaf6, 32'h00000000} /* (5, 17, 27) {real, imag} */,
  {32'hc4110eb4, 32'h00000000} /* (5, 17, 26) {real, imag} */,
  {32'h430b3c39, 32'h00000000} /* (5, 17, 25) {real, imag} */,
  {32'hc375be53, 32'h00000000} /* (5, 17, 24) {real, imag} */,
  {32'hc1ee77b0, 32'h00000000} /* (5, 17, 23) {real, imag} */,
  {32'h43f253e8, 32'h00000000} /* (5, 17, 22) {real, imag} */,
  {32'h44220d46, 32'h00000000} /* (5, 17, 21) {real, imag} */,
  {32'h44a6a9f4, 32'h00000000} /* (5, 17, 20) {real, imag} */,
  {32'h444abd6f, 32'h00000000} /* (5, 17, 19) {real, imag} */,
  {32'h43cbf068, 32'h00000000} /* (5, 17, 18) {real, imag} */,
  {32'h439eddb4, 32'h00000000} /* (5, 17, 17) {real, imag} */,
  {32'h44b7e15a, 32'h00000000} /* (5, 17, 16) {real, imag} */,
  {32'h445552a8, 32'h00000000} /* (5, 17, 15) {real, imag} */,
  {32'h44643052, 32'h00000000} /* (5, 17, 14) {real, imag} */,
  {32'h43b68e40, 32'h00000000} /* (5, 17, 13) {real, imag} */,
  {32'h42cc2fd0, 32'h00000000} /* (5, 17, 12) {real, imag} */,
  {32'hc30f8122, 32'h00000000} /* (5, 17, 11) {real, imag} */,
  {32'h43411823, 32'h00000000} /* (5, 17, 10) {real, imag} */,
  {32'hc26dad6c, 32'h00000000} /* (5, 17, 9) {real, imag} */,
  {32'h4399690c, 32'h00000000} /* (5, 17, 8) {real, imag} */,
  {32'hc3c9c595, 32'h00000000} /* (5, 17, 7) {real, imag} */,
  {32'hc3868ffc, 32'h00000000} /* (5, 17, 6) {real, imag} */,
  {32'hc3dd2e2c, 32'h00000000} /* (5, 17, 5) {real, imag} */,
  {32'hc4140940, 32'h00000000} /* (5, 17, 4) {real, imag} */,
  {32'hc3fdf9ca, 32'h00000000} /* (5, 17, 3) {real, imag} */,
  {32'hc3f6793c, 32'h00000000} /* (5, 17, 2) {real, imag} */,
  {32'hc38bf7c2, 32'h00000000} /* (5, 17, 1) {real, imag} */,
  {32'hc45c4ff9, 32'h00000000} /* (5, 17, 0) {real, imag} */,
  {32'hc4704053, 32'h00000000} /* (5, 16, 31) {real, imag} */,
  {32'hc49e76a8, 32'h00000000} /* (5, 16, 30) {real, imag} */,
  {32'hc4c564cd, 32'h00000000} /* (5, 16, 29) {real, imag} */,
  {32'hc40880f8, 32'h00000000} /* (5, 16, 28) {real, imag} */,
  {32'hc44dbf90, 32'h00000000} /* (5, 16, 27) {real, imag} */,
  {32'hc41f266a, 32'h00000000} /* (5, 16, 26) {real, imag} */,
  {32'hc20625c4, 32'h00000000} /* (5, 16, 25) {real, imag} */,
  {32'hc34bddfe, 32'h00000000} /* (5, 16, 24) {real, imag} */,
  {32'h4477f089, 32'h00000000} /* (5, 16, 23) {real, imag} */,
  {32'h444be54d, 32'h00000000} /* (5, 16, 22) {real, imag} */,
  {32'h445f9592, 32'h00000000} /* (5, 16, 21) {real, imag} */,
  {32'h448cb008, 32'h00000000} /* (5, 16, 20) {real, imag} */,
  {32'h447ffdfc, 32'h00000000} /* (5, 16, 19) {real, imag} */,
  {32'h445b3cd0, 32'h00000000} /* (5, 16, 18) {real, imag} */,
  {32'h44700540, 32'h00000000} /* (5, 16, 17) {real, imag} */,
  {32'hc406cb5e, 32'h00000000} /* (5, 16, 16) {real, imag} */,
  {32'h434ba04c, 32'h00000000} /* (5, 16, 15) {real, imag} */,
  {32'h44a66da2, 32'h00000000} /* (5, 16, 14) {real, imag} */,
  {32'h44922f93, 32'h00000000} /* (5, 16, 13) {real, imag} */,
  {32'hc3badeb4, 32'h00000000} /* (5, 16, 12) {real, imag} */,
  {32'hc3a1925f, 32'h00000000} /* (5, 16, 11) {real, imag} */,
  {32'h438d3ea8, 32'h00000000} /* (5, 16, 10) {real, imag} */,
  {32'hc396ccb6, 32'h00000000} /* (5, 16, 9) {real, imag} */,
  {32'h4351d7ae, 32'h00000000} /* (5, 16, 8) {real, imag} */,
  {32'hc3283e6c, 32'h00000000} /* (5, 16, 7) {real, imag} */,
  {32'hc3e6b5f2, 32'h00000000} /* (5, 16, 6) {real, imag} */,
  {32'hc3da5d00, 32'h00000000} /* (5, 16, 5) {real, imag} */,
  {32'hc425e44a, 32'h00000000} /* (5, 16, 4) {real, imag} */,
  {32'hc4e6efc4, 32'h00000000} /* (5, 16, 3) {real, imag} */,
  {32'hc4b78786, 32'h00000000} /* (5, 16, 2) {real, imag} */,
  {32'hc473f6e4, 32'h00000000} /* (5, 16, 1) {real, imag} */,
  {32'hc450413e, 32'h00000000} /* (5, 16, 0) {real, imag} */,
  {32'hc3d907ba, 32'h00000000} /* (5, 15, 31) {real, imag} */,
  {32'hc48acf20, 32'h00000000} /* (5, 15, 30) {real, imag} */,
  {32'hc4333977, 32'h00000000} /* (5, 15, 29) {real, imag} */,
  {32'hc4521a29, 32'h00000000} /* (5, 15, 28) {real, imag} */,
  {32'hc42eb11c, 32'h00000000} /* (5, 15, 27) {real, imag} */,
  {32'hc3e9a92e, 32'h00000000} /* (5, 15, 26) {real, imag} */,
  {32'hc49b26f7, 32'h00000000} /* (5, 15, 25) {real, imag} */,
  {32'hc3c0f7f6, 32'h00000000} /* (5, 15, 24) {real, imag} */,
  {32'h43cf301b, 32'h00000000} /* (5, 15, 23) {real, imag} */,
  {32'h43c273c3, 32'h00000000} /* (5, 15, 22) {real, imag} */,
  {32'h43b97b5b, 32'h00000000} /* (5, 15, 21) {real, imag} */,
  {32'h44a740cb, 32'h00000000} /* (5, 15, 20) {real, imag} */,
  {32'h448aa428, 32'h00000000} /* (5, 15, 19) {real, imag} */,
  {32'h4411eabd, 32'h00000000} /* (5, 15, 18) {real, imag} */,
  {32'h4436b247, 32'h00000000} /* (5, 15, 17) {real, imag} */,
  {32'h4458d697, 32'h00000000} /* (5, 15, 16) {real, imag} */,
  {32'hc3fa59c8, 32'h00000000} /* (5, 15, 15) {real, imag} */,
  {32'h4397419b, 32'h00000000} /* (5, 15, 14) {real, imag} */,
  {32'hc497c653, 32'h00000000} /* (5, 15, 13) {real, imag} */,
  {32'hc4a477fe, 32'h00000000} /* (5, 15, 12) {real, imag} */,
  {32'hc34625da, 32'h00000000} /* (5, 15, 11) {real, imag} */,
  {32'hc45c83df, 32'h00000000} /* (5, 15, 10) {real, imag} */,
  {32'h43f680b0, 32'h00000000} /* (5, 15, 9) {real, imag} */,
  {32'hc448250f, 32'h00000000} /* (5, 15, 8) {real, imag} */,
  {32'hc47371c2, 32'h00000000} /* (5, 15, 7) {real, imag} */,
  {32'hc434d230, 32'h00000000} /* (5, 15, 6) {real, imag} */,
  {32'hc4857433, 32'h00000000} /* (5, 15, 5) {real, imag} */,
  {32'hc4b6e891, 32'h00000000} /* (5, 15, 4) {real, imag} */,
  {32'hc5056511, 32'h00000000} /* (5, 15, 3) {real, imag} */,
  {32'hc5057dd8, 32'h00000000} /* (5, 15, 2) {real, imag} */,
  {32'hc41f9dbb, 32'h00000000} /* (5, 15, 1) {real, imag} */,
  {32'hc4aec78e, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'hc45854ef, 32'h00000000} /* (5, 14, 31) {real, imag} */,
  {32'hc3f213c7, 32'h00000000} /* (5, 14, 30) {real, imag} */,
  {32'hc3ee25e5, 32'h00000000} /* (5, 14, 29) {real, imag} */,
  {32'hc450075a, 32'h00000000} /* (5, 14, 28) {real, imag} */,
  {32'hc3c17040, 32'h00000000} /* (5, 14, 27) {real, imag} */,
  {32'hc4640b15, 32'h00000000} /* (5, 14, 26) {real, imag} */,
  {32'hc4bbd0bc, 32'h00000000} /* (5, 14, 25) {real, imag} */,
  {32'hc4a6c2ca, 32'h00000000} /* (5, 14, 24) {real, imag} */,
  {32'hc3542fde, 32'h00000000} /* (5, 14, 23) {real, imag} */,
  {32'h42b7d258, 32'h00000000} /* (5, 14, 22) {real, imag} */,
  {32'h43a50ede, 32'h00000000} /* (5, 14, 21) {real, imag} */,
  {32'hc3c53550, 32'h00000000} /* (5, 14, 20) {real, imag} */,
  {32'hc376f958, 32'h00000000} /* (5, 14, 19) {real, imag} */,
  {32'h44097928, 32'h00000000} /* (5, 14, 18) {real, imag} */,
  {32'hc470c590, 32'h00000000} /* (5, 14, 17) {real, imag} */,
  {32'h43ae67c3, 32'h00000000} /* (5, 14, 16) {real, imag} */,
  {32'h43934b52, 32'h00000000} /* (5, 14, 15) {real, imag} */,
  {32'h434e5b5e, 32'h00000000} /* (5, 14, 14) {real, imag} */,
  {32'hc43c6044, 32'h00000000} /* (5, 14, 13) {real, imag} */,
  {32'h4336ed60, 32'h00000000} /* (5, 14, 12) {real, imag} */,
  {32'hc3cac5da, 32'h00000000} /* (5, 14, 11) {real, imag} */,
  {32'hc441fdeb, 32'h00000000} /* (5, 14, 10) {real, imag} */,
  {32'hc29dd4e8, 32'h00000000} /* (5, 14, 9) {real, imag} */,
  {32'hc37e8bc0, 32'h00000000} /* (5, 14, 8) {real, imag} */,
  {32'hc48c9b7f, 32'h00000000} /* (5, 14, 7) {real, imag} */,
  {32'hc48ed938, 32'h00000000} /* (5, 14, 6) {real, imag} */,
  {32'hc4d92458, 32'h00000000} /* (5, 14, 5) {real, imag} */,
  {32'hc4dcf08c, 32'h00000000} /* (5, 14, 4) {real, imag} */,
  {32'hc4d2d345, 32'h00000000} /* (5, 14, 3) {real, imag} */,
  {32'hc503c1b2, 32'h00000000} /* (5, 14, 2) {real, imag} */,
  {32'hc4ca160e, 32'h00000000} /* (5, 14, 1) {real, imag} */,
  {32'hc42362ea, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hc3718e5c, 32'h00000000} /* (5, 13, 31) {real, imag} */,
  {32'hc420842a, 32'h00000000} /* (5, 13, 30) {real, imag} */,
  {32'h438a715e, 32'h00000000} /* (5, 13, 29) {real, imag} */,
  {32'h4481ae0e, 32'h00000000} /* (5, 13, 28) {real, imag} */,
  {32'h43cd6578, 32'h00000000} /* (5, 13, 27) {real, imag} */,
  {32'h4349981e, 32'h00000000} /* (5, 13, 26) {real, imag} */,
  {32'hc489120c, 32'h00000000} /* (5, 13, 25) {real, imag} */,
  {32'hc4956309, 32'h00000000} /* (5, 13, 24) {real, imag} */,
  {32'hc3d5c4ca, 32'h00000000} /* (5, 13, 23) {real, imag} */,
  {32'h44c19a36, 32'h00000000} /* (5, 13, 22) {real, imag} */,
  {32'h44a0df53, 32'h00000000} /* (5, 13, 21) {real, imag} */,
  {32'hc4d6fa26, 32'h00000000} /* (5, 13, 20) {real, imag} */,
  {32'hc3cc0f00, 32'h00000000} /* (5, 13, 19) {real, imag} */,
  {32'hc49fc3c2, 32'h00000000} /* (5, 13, 18) {real, imag} */,
  {32'hc46c318d, 32'h00000000} /* (5, 13, 17) {real, imag} */,
  {32'hc3aa3c37, 32'h00000000} /* (5, 13, 16) {real, imag} */,
  {32'hc14f93b8, 32'h00000000} /* (5, 13, 15) {real, imag} */,
  {32'hc1309500, 32'h00000000} /* (5, 13, 14) {real, imag} */,
  {32'hc39828a2, 32'h00000000} /* (5, 13, 13) {real, imag} */,
  {32'hc30d0944, 32'h00000000} /* (5, 13, 12) {real, imag} */,
  {32'hc39b76ac, 32'h00000000} /* (5, 13, 11) {real, imag} */,
  {32'hc3e0095d, 32'h00000000} /* (5, 13, 10) {real, imag} */,
  {32'hc42e44b2, 32'h00000000} /* (5, 13, 9) {real, imag} */,
  {32'hc4535a62, 32'h00000000} /* (5, 13, 8) {real, imag} */,
  {32'hc4870d96, 32'h00000000} /* (5, 13, 7) {real, imag} */,
  {32'hc478717f, 32'h00000000} /* (5, 13, 6) {real, imag} */,
  {32'hc4aae351, 32'h00000000} /* (5, 13, 5) {real, imag} */,
  {32'hc4cb7650, 32'h00000000} /* (5, 13, 4) {real, imag} */,
  {32'hc4f5dc40, 32'h00000000} /* (5, 13, 3) {real, imag} */,
  {32'hc47b4875, 32'h00000000} /* (5, 13, 2) {real, imag} */,
  {32'hc41d40e1, 32'h00000000} /* (5, 13, 1) {real, imag} */,
  {32'hc3f199f3, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'h43403706, 32'h00000000} /* (5, 12, 31) {real, imag} */,
  {32'hc359da64, 32'h00000000} /* (5, 12, 30) {real, imag} */,
  {32'h444bb2bf, 32'h00000000} /* (5, 12, 29) {real, imag} */,
  {32'h4465afcd, 32'h00000000} /* (5, 12, 28) {real, imag} */,
  {32'h43bf0897, 32'h00000000} /* (5, 12, 27) {real, imag} */,
  {32'hc43e73a2, 32'h00000000} /* (5, 12, 26) {real, imag} */,
  {32'hc3119280, 32'h00000000} /* (5, 12, 25) {real, imag} */,
  {32'hc46c63b1, 32'h00000000} /* (5, 12, 24) {real, imag} */,
  {32'h423de8c0, 32'h00000000} /* (5, 12, 23) {real, imag} */,
  {32'h4380482e, 32'h00000000} /* (5, 12, 22) {real, imag} */,
  {32'h448bdd6f, 32'h00000000} /* (5, 12, 21) {real, imag} */,
  {32'hc39fd8c9, 32'h00000000} /* (5, 12, 20) {real, imag} */,
  {32'hc4b62a76, 32'h00000000} /* (5, 12, 19) {real, imag} */,
  {32'hc409ed7c, 32'h00000000} /* (5, 12, 18) {real, imag} */,
  {32'hc3367b42, 32'h00000000} /* (5, 12, 17) {real, imag} */,
  {32'h41428538, 32'h00000000} /* (5, 12, 16) {real, imag} */,
  {32'h43be188d, 32'h00000000} /* (5, 12, 15) {real, imag} */,
  {32'hc43371eb, 32'h00000000} /* (5, 12, 14) {real, imag} */,
  {32'h4323e1b4, 32'h00000000} /* (5, 12, 13) {real, imag} */,
  {32'h43d50ede, 32'h00000000} /* (5, 12, 12) {real, imag} */,
  {32'h43198fa2, 32'h00000000} /* (5, 12, 11) {real, imag} */,
  {32'hc318a2ea, 32'h00000000} /* (5, 12, 10) {real, imag} */,
  {32'hc481db1c, 32'h00000000} /* (5, 12, 9) {real, imag} */,
  {32'hc4143cf7, 32'h00000000} /* (5, 12, 8) {real, imag} */,
  {32'hc47877e4, 32'h00000000} /* (5, 12, 7) {real, imag} */,
  {32'hc4876422, 32'h00000000} /* (5, 12, 6) {real, imag} */,
  {32'hc43b6b9a, 32'h00000000} /* (5, 12, 5) {real, imag} */,
  {32'hc4457624, 32'h00000000} /* (5, 12, 4) {real, imag} */,
  {32'hc38608ca, 32'h00000000} /* (5, 12, 3) {real, imag} */,
  {32'h441880b4, 32'h00000000} /* (5, 12, 2) {real, imag} */,
  {32'h4424ff82, 32'h00000000} /* (5, 12, 1) {real, imag} */,
  {32'h4318c6e4, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h441a8118, 32'h00000000} /* (5, 11, 31) {real, imag} */,
  {32'h4499bc49, 32'h00000000} /* (5, 11, 30) {real, imag} */,
  {32'h43ac4f3a, 32'h00000000} /* (5, 11, 29) {real, imag} */,
  {32'h448470a4, 32'h00000000} /* (5, 11, 28) {real, imag} */,
  {32'h44328a27, 32'h00000000} /* (5, 11, 27) {real, imag} */,
  {32'h427996fd, 32'h00000000} /* (5, 11, 26) {real, imag} */,
  {32'h448211cf, 32'h00000000} /* (5, 11, 25) {real, imag} */,
  {32'h4369b0cc, 32'h00000000} /* (5, 11, 24) {real, imag} */,
  {32'h43ab4f41, 32'h00000000} /* (5, 11, 23) {real, imag} */,
  {32'h44e91592, 32'h00000000} /* (5, 11, 22) {real, imag} */,
  {32'h447f4f26, 32'h00000000} /* (5, 11, 21) {real, imag} */,
  {32'h4451a211, 32'h00000000} /* (5, 11, 20) {real, imag} */,
  {32'hc46829ea, 32'h00000000} /* (5, 11, 19) {real, imag} */,
  {32'h42ad4050, 32'h00000000} /* (5, 11, 18) {real, imag} */,
  {32'hc41a9977, 32'h00000000} /* (5, 11, 17) {real, imag} */,
  {32'h420b9920, 32'h00000000} /* (5, 11, 16) {real, imag} */,
  {32'h433a9f56, 32'h00000000} /* (5, 11, 15) {real, imag} */,
  {32'h43695e18, 32'h00000000} /* (5, 11, 14) {real, imag} */,
  {32'hc46cd35d, 32'h00000000} /* (5, 11, 13) {real, imag} */,
  {32'hc30a3f3c, 32'h00000000} /* (5, 11, 12) {real, imag} */,
  {32'hc289b1a8, 32'h00000000} /* (5, 11, 11) {real, imag} */,
  {32'hbf3c6340, 32'h00000000} /* (5, 11, 10) {real, imag} */,
  {32'hc40c2b4c, 32'h00000000} /* (5, 11, 9) {real, imag} */,
  {32'hc44a8e69, 32'h00000000} /* (5, 11, 8) {real, imag} */,
  {32'hc31afdf2, 32'h00000000} /* (5, 11, 7) {real, imag} */,
  {32'hc4821ab6, 32'h00000000} /* (5, 11, 6) {real, imag} */,
  {32'hc447ebce, 32'h00000000} /* (5, 11, 5) {real, imag} */,
  {32'h42cdf468, 32'h00000000} /* (5, 11, 4) {real, imag} */,
  {32'hc4242428, 32'h00000000} /* (5, 11, 3) {real, imag} */,
  {32'hc36ba1a4, 32'h00000000} /* (5, 11, 2) {real, imag} */,
  {32'h44ff08cc, 32'h00000000} /* (5, 11, 1) {real, imag} */,
  {32'h449e86ca, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'h44862128, 32'h00000000} /* (5, 10, 31) {real, imag} */,
  {32'h44d39284, 32'h00000000} /* (5, 10, 30) {real, imag} */,
  {32'h44969a3f, 32'h00000000} /* (5, 10, 29) {real, imag} */,
  {32'h43ee17c9, 32'h00000000} /* (5, 10, 28) {real, imag} */,
  {32'h445c7002, 32'h00000000} /* (5, 10, 27) {real, imag} */,
  {32'h4498f7d0, 32'h00000000} /* (5, 10, 26) {real, imag} */,
  {32'h433969ac, 32'h00000000} /* (5, 10, 25) {real, imag} */,
  {32'h43e0037d, 32'h00000000} /* (5, 10, 24) {real, imag} */,
  {32'h44e6dc88, 32'h00000000} /* (5, 10, 23) {real, imag} */,
  {32'h44c81c6c, 32'h00000000} /* (5, 10, 22) {real, imag} */,
  {32'hc3defaf9, 32'h00000000} /* (5, 10, 21) {real, imag} */,
  {32'h442bd004, 32'h00000000} /* (5, 10, 20) {real, imag} */,
  {32'h44e6ba8b, 32'h00000000} /* (5, 10, 19) {real, imag} */,
  {32'hc3e1694d, 32'h00000000} /* (5, 10, 18) {real, imag} */,
  {32'hc2e92604, 32'h00000000} /* (5, 10, 17) {real, imag} */,
  {32'h44109e22, 32'h00000000} /* (5, 10, 16) {real, imag} */,
  {32'h4410ddde, 32'h00000000} /* (5, 10, 15) {real, imag} */,
  {32'h4357fc1c, 32'h00000000} /* (5, 10, 14) {real, imag} */,
  {32'hc3c6531d, 32'h00000000} /* (5, 10, 13) {real, imag} */,
  {32'hc402714a, 32'h00000000} /* (5, 10, 12) {real, imag} */,
  {32'h4380e07c, 32'h00000000} /* (5, 10, 11) {real, imag} */,
  {32'hc44b77a5, 32'h00000000} /* (5, 10, 10) {real, imag} */,
  {32'hc4ad6712, 32'h00000000} /* (5, 10, 9) {real, imag} */,
  {32'h438c9527, 32'h00000000} /* (5, 10, 8) {real, imag} */,
  {32'hc263ac10, 32'h00000000} /* (5, 10, 7) {real, imag} */,
  {32'hc4aca4f0, 32'h00000000} /* (5, 10, 6) {real, imag} */,
  {32'hc38706a1, 32'h00000000} /* (5, 10, 5) {real, imag} */,
  {32'hc3e5b2ed, 32'h00000000} /* (5, 10, 4) {real, imag} */,
  {32'h43f529dc, 32'h00000000} /* (5, 10, 3) {real, imag} */,
  {32'hc393f0db, 32'h00000000} /* (5, 10, 2) {real, imag} */,
  {32'h44153bea, 32'h00000000} /* (5, 10, 1) {real, imag} */,
  {32'h44816b72, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'h44a7cf8b, 32'h00000000} /* (5, 9, 31) {real, imag} */,
  {32'h4458e278, 32'h00000000} /* (5, 9, 30) {real, imag} */,
  {32'h4483bd4d, 32'h00000000} /* (5, 9, 29) {real, imag} */,
  {32'h44a785b2, 32'h00000000} /* (5, 9, 28) {real, imag} */,
  {32'h442dd824, 32'h00000000} /* (5, 9, 27) {real, imag} */,
  {32'h449e6664, 32'h00000000} /* (5, 9, 26) {real, imag} */,
  {32'h449b6fae, 32'h00000000} /* (5, 9, 25) {real, imag} */,
  {32'h44042f56, 32'h00000000} /* (5, 9, 24) {real, imag} */,
  {32'h44fabe48, 32'h00000000} /* (5, 9, 23) {real, imag} */,
  {32'h44bcb3b3, 32'h00000000} /* (5, 9, 22) {real, imag} */,
  {32'h446f2b6a, 32'h00000000} /* (5, 9, 21) {real, imag} */,
  {32'h4499d73c, 32'h00000000} /* (5, 9, 20) {real, imag} */,
  {32'h443cf9ce, 32'h00000000} /* (5, 9, 19) {real, imag} */,
  {32'h444a8d6b, 32'h00000000} /* (5, 9, 18) {real, imag} */,
  {32'h440aedfd, 32'h00000000} /* (5, 9, 17) {real, imag} */,
  {32'h449569a5, 32'h00000000} /* (5, 9, 16) {real, imag} */,
  {32'h449584dd, 32'h00000000} /* (5, 9, 15) {real, imag} */,
  {32'hc41d1aec, 32'h00000000} /* (5, 9, 14) {real, imag} */,
  {32'h4107b480, 32'h00000000} /* (5, 9, 13) {real, imag} */,
  {32'h431355bc, 32'h00000000} /* (5, 9, 12) {real, imag} */,
  {32'h44351862, 32'h00000000} /* (5, 9, 11) {real, imag} */,
  {32'hc3b35d1c, 32'h00000000} /* (5, 9, 10) {real, imag} */,
  {32'hc23088f0, 32'h00000000} /* (5, 9, 9) {real, imag} */,
  {32'hc45eae3e, 32'h00000000} /* (5, 9, 8) {real, imag} */,
  {32'h438d9670, 32'h00000000} /* (5, 9, 7) {real, imag} */,
  {32'h436a04b8, 32'h00000000} /* (5, 9, 6) {real, imag} */,
  {32'hc310b8b0, 32'h00000000} /* (5, 9, 5) {real, imag} */,
  {32'h43eb384b, 32'h00000000} /* (5, 9, 4) {real, imag} */,
  {32'h43f6eee9, 32'h00000000} /* (5, 9, 3) {real, imag} */,
  {32'h43d83e86, 32'h00000000} /* (5, 9, 2) {real, imag} */,
  {32'h44956c68, 32'h00000000} /* (5, 9, 1) {real, imag} */,
  {32'h44c12cb3, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'h4503804f, 32'h00000000} /* (5, 8, 31) {real, imag} */,
  {32'h4499dc92, 32'h00000000} /* (5, 8, 30) {real, imag} */,
  {32'h44c5c4cf, 32'h00000000} /* (5, 8, 29) {real, imag} */,
  {32'h44098c45, 32'h00000000} /* (5, 8, 28) {real, imag} */,
  {32'h446e1ba6, 32'h00000000} /* (5, 8, 27) {real, imag} */,
  {32'h445eea79, 32'h00000000} /* (5, 8, 26) {real, imag} */,
  {32'h414e1b40, 32'h00000000} /* (5, 8, 25) {real, imag} */,
  {32'h44dad77a, 32'h00000000} /* (5, 8, 24) {real, imag} */,
  {32'h450a2028, 32'h00000000} /* (5, 8, 23) {real, imag} */,
  {32'h44b24a7c, 32'h00000000} /* (5, 8, 22) {real, imag} */,
  {32'h450d63cc, 32'h00000000} /* (5, 8, 21) {real, imag} */,
  {32'h4505c6c4, 32'h00000000} /* (5, 8, 20) {real, imag} */,
  {32'h44dc0f9c, 32'h00000000} /* (5, 8, 19) {real, imag} */,
  {32'h44c0a027, 32'h00000000} /* (5, 8, 18) {real, imag} */,
  {32'h44abe251, 32'h00000000} /* (5, 8, 17) {real, imag} */,
  {32'h43bf4f8e, 32'h00000000} /* (5, 8, 16) {real, imag} */,
  {32'h441ff3ab, 32'h00000000} /* (5, 8, 15) {real, imag} */,
  {32'hc3ebf782, 32'h00000000} /* (5, 8, 14) {real, imag} */,
  {32'hc4b943fd, 32'h00000000} /* (5, 8, 13) {real, imag} */,
  {32'hc4205f85, 32'h00000000} /* (5, 8, 12) {real, imag} */,
  {32'h44278bd2, 32'h00000000} /* (5, 8, 11) {real, imag} */,
  {32'hbef98800, 32'h00000000} /* (5, 8, 10) {real, imag} */,
  {32'hc408025d, 32'h00000000} /* (5, 8, 9) {real, imag} */,
  {32'h434ebc4c, 32'h00000000} /* (5, 8, 8) {real, imag} */,
  {32'h433e5028, 32'h00000000} /* (5, 8, 7) {real, imag} */,
  {32'hc1a3cfe0, 32'h00000000} /* (5, 8, 6) {real, imag} */,
  {32'hc28a53a0, 32'h00000000} /* (5, 8, 5) {real, imag} */,
  {32'h44101fd7, 32'h00000000} /* (5, 8, 4) {real, imag} */,
  {32'h44a511b8, 32'h00000000} /* (5, 8, 3) {real, imag} */,
  {32'h44b9682f, 32'h00000000} /* (5, 8, 2) {real, imag} */,
  {32'h45045388, 32'h00000000} /* (5, 8, 1) {real, imag} */,
  {32'h44e0420c, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'h452d71ce, 32'h00000000} /* (5, 7, 31) {real, imag} */,
  {32'h44de7a6a, 32'h00000000} /* (5, 7, 30) {real, imag} */,
  {32'h44c7208c, 32'h00000000} /* (5, 7, 29) {real, imag} */,
  {32'h44a9c050, 32'h00000000} /* (5, 7, 28) {real, imag} */,
  {32'h4471f3a2, 32'h00000000} /* (5, 7, 27) {real, imag} */,
  {32'h44ddc2dc, 32'h00000000} /* (5, 7, 26) {real, imag} */,
  {32'h42639900, 32'h00000000} /* (5, 7, 25) {real, imag} */,
  {32'h4399d461, 32'h00000000} /* (5, 7, 24) {real, imag} */,
  {32'h4539f6f5, 32'h00000000} /* (5, 7, 23) {real, imag} */,
  {32'h45250e7e, 32'h00000000} /* (5, 7, 22) {real, imag} */,
  {32'h44b81740, 32'h00000000} /* (5, 7, 21) {real, imag} */,
  {32'h453cfc82, 32'h00000000} /* (5, 7, 20) {real, imag} */,
  {32'h44e43928, 32'h00000000} /* (5, 7, 19) {real, imag} */,
  {32'h44dab80f, 32'h00000000} /* (5, 7, 18) {real, imag} */,
  {32'h44b7a814, 32'h00000000} /* (5, 7, 17) {real, imag} */,
  {32'h4485f960, 32'h00000000} /* (5, 7, 16) {real, imag} */,
  {32'hc2995b00, 32'h00000000} /* (5, 7, 15) {real, imag} */,
  {32'hc4dd8fba, 32'h00000000} /* (5, 7, 14) {real, imag} */,
  {32'hc4aa9d52, 32'h00000000} /* (5, 7, 13) {real, imag} */,
  {32'h411072c0, 32'h00000000} /* (5, 7, 12) {real, imag} */,
  {32'h43e3c620, 32'h00000000} /* (5, 7, 11) {real, imag} */,
  {32'hc41c5f21, 32'h00000000} /* (5, 7, 10) {real, imag} */,
  {32'hc3d42930, 32'h00000000} /* (5, 7, 9) {real, imag} */,
  {32'h4463e22c, 32'h00000000} /* (5, 7, 8) {real, imag} */,
  {32'h4487a0d6, 32'h00000000} /* (5, 7, 7) {real, imag} */,
  {32'hc3c48894, 32'h00000000} /* (5, 7, 6) {real, imag} */,
  {32'h4406127a, 32'h00000000} /* (5, 7, 5) {real, imag} */,
  {32'h4454aa26, 32'h00000000} /* (5, 7, 4) {real, imag} */,
  {32'h44d752d4, 32'h00000000} /* (5, 7, 3) {real, imag} */,
  {32'h4554a81e, 32'h00000000} /* (5, 7, 2) {real, imag} */,
  {32'h4504f5f4, 32'h00000000} /* (5, 7, 1) {real, imag} */,
  {32'h450280db, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'h45188ab6, 32'h00000000} /* (5, 6, 31) {real, imag} */,
  {32'h453ac8e8, 32'h00000000} /* (5, 6, 30) {real, imag} */,
  {32'h44767d8a, 32'h00000000} /* (5, 6, 29) {real, imag} */,
  {32'h44c35c1e, 32'h00000000} /* (5, 6, 28) {real, imag} */,
  {32'h44f74fd6, 32'h00000000} /* (5, 6, 27) {real, imag} */,
  {32'h44c975ce, 32'h00000000} /* (5, 6, 26) {real, imag} */,
  {32'h4514e3e1, 32'h00000000} /* (5, 6, 25) {real, imag} */,
  {32'h44f25a0a, 32'h00000000} /* (5, 6, 24) {real, imag} */,
  {32'h452e7d18, 32'h00000000} /* (5, 6, 23) {real, imag} */,
  {32'h454f078e, 32'h00000000} /* (5, 6, 22) {real, imag} */,
  {32'h450ba4ee, 32'h00000000} /* (5, 6, 21) {real, imag} */,
  {32'h44cac787, 32'h00000000} /* (5, 6, 20) {real, imag} */,
  {32'h44abf7ba, 32'h00000000} /* (5, 6, 19) {real, imag} */,
  {32'h4485e3d7, 32'h00000000} /* (5, 6, 18) {real, imag} */,
  {32'h43ddfab8, 32'h00000000} /* (5, 6, 17) {real, imag} */,
  {32'h43ba7098, 32'h00000000} /* (5, 6, 16) {real, imag} */,
  {32'hc438b392, 32'h00000000} /* (5, 6, 15) {real, imag} */,
  {32'h42befc90, 32'h00000000} /* (5, 6, 14) {real, imag} */,
  {32'hc3aab674, 32'h00000000} /* (5, 6, 13) {real, imag} */,
  {32'hc407f34b, 32'h00000000} /* (5, 6, 12) {real, imag} */,
  {32'h44214860, 32'h00000000} /* (5, 6, 11) {real, imag} */,
  {32'h43917750, 32'h00000000} /* (5, 6, 10) {real, imag} */,
  {32'h444df3fd, 32'h00000000} /* (5, 6, 9) {real, imag} */,
  {32'h448398ea, 32'h00000000} /* (5, 6, 8) {real, imag} */,
  {32'h4426ee8a, 32'h00000000} /* (5, 6, 7) {real, imag} */,
  {32'h448b966c, 32'h00000000} /* (5, 6, 6) {real, imag} */,
  {32'h44e8f3f4, 32'h00000000} /* (5, 6, 5) {real, imag} */,
  {32'h44d86909, 32'h00000000} /* (5, 6, 4) {real, imag} */,
  {32'h45000f5c, 32'h00000000} /* (5, 6, 3) {real, imag} */,
  {32'h452624ae, 32'h00000000} /* (5, 6, 2) {real, imag} */,
  {32'h451825dd, 32'h00000000} /* (5, 6, 1) {real, imag} */,
  {32'h452bef1b, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'h455b71f6, 32'h00000000} /* (5, 5, 31) {real, imag} */,
  {32'h4544563a, 32'h00000000} /* (5, 5, 30) {real, imag} */,
  {32'h45163561, 32'h00000000} /* (5, 5, 29) {real, imag} */,
  {32'h44b1de38, 32'h00000000} /* (5, 5, 28) {real, imag} */,
  {32'h4526b48e, 32'h00000000} /* (5, 5, 27) {real, imag} */,
  {32'h452e58e4, 32'h00000000} /* (5, 5, 26) {real, imag} */,
  {32'h44dab882, 32'h00000000} /* (5, 5, 25) {real, imag} */,
  {32'h451fd4b2, 32'h00000000} /* (5, 5, 24) {real, imag} */,
  {32'h452ac0f6, 32'h00000000} /* (5, 5, 23) {real, imag} */,
  {32'h4521807c, 32'h00000000} /* (5, 5, 22) {real, imag} */,
  {32'h4514e968, 32'h00000000} /* (5, 5, 21) {real, imag} */,
  {32'h4423bd0f, 32'h00000000} /* (5, 5, 20) {real, imag} */,
  {32'h43f38c30, 32'h00000000} /* (5, 5, 19) {real, imag} */,
  {32'h44447001, 32'h00000000} /* (5, 5, 18) {real, imag} */,
  {32'hc410c872, 32'h00000000} /* (5, 5, 17) {real, imag} */,
  {32'hc38660a8, 32'h00000000} /* (5, 5, 16) {real, imag} */,
  {32'hc37f8ea8, 32'h00000000} /* (5, 5, 15) {real, imag} */,
  {32'h42e0b7c0, 32'h00000000} /* (5, 5, 14) {real, imag} */,
  {32'hc4470f58, 32'h00000000} /* (5, 5, 13) {real, imag} */,
  {32'h43665844, 32'h00000000} /* (5, 5, 12) {real, imag} */,
  {32'hc428ea30, 32'h00000000} /* (5, 5, 11) {real, imag} */,
  {32'h43d8f154, 32'h00000000} /* (5, 5, 10) {real, imag} */,
  {32'h42b71e88, 32'h00000000} /* (5, 5, 9) {real, imag} */,
  {32'h444f4e2a, 32'h00000000} /* (5, 5, 8) {real, imag} */,
  {32'h4498ba80, 32'h00000000} /* (5, 5, 7) {real, imag} */,
  {32'h448a1080, 32'h00000000} /* (5, 5, 6) {real, imag} */,
  {32'h45388b74, 32'h00000000} /* (5, 5, 5) {real, imag} */,
  {32'h4519d834, 32'h00000000} /* (5, 5, 4) {real, imag} */,
  {32'h452d5b62, 32'h00000000} /* (5, 5, 3) {real, imag} */,
  {32'h451e44c2, 32'h00000000} /* (5, 5, 2) {real, imag} */,
  {32'h452f0bf6, 32'h00000000} /* (5, 5, 1) {real, imag} */,
  {32'h453b839d, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'h4546d699, 32'h00000000} /* (5, 4, 31) {real, imag} */,
  {32'h453b2eaa, 32'h00000000} /* (5, 4, 30) {real, imag} */,
  {32'h45166a40, 32'h00000000} /* (5, 4, 29) {real, imag} */,
  {32'h4510048e, 32'h00000000} /* (5, 4, 28) {real, imag} */,
  {32'h4526c3ee, 32'h00000000} /* (5, 4, 27) {real, imag} */,
  {32'h4523f504, 32'h00000000} /* (5, 4, 26) {real, imag} */,
  {32'h4518a2ee, 32'h00000000} /* (5, 4, 25) {real, imag} */,
  {32'h45058f8d, 32'h00000000} /* (5, 4, 24) {real, imag} */,
  {32'h453da3c5, 32'h00000000} /* (5, 4, 23) {real, imag} */,
  {32'h4528b3a8, 32'h00000000} /* (5, 4, 22) {real, imag} */,
  {32'h44c776e2, 32'h00000000} /* (5, 4, 21) {real, imag} */,
  {32'h44d72f98, 32'h00000000} /* (5, 4, 20) {real, imag} */,
  {32'h43ed2f34, 32'h00000000} /* (5, 4, 19) {real, imag} */,
  {32'hc238a120, 32'h00000000} /* (5, 4, 18) {real, imag} */,
  {32'h43325c58, 32'h00000000} /* (5, 4, 17) {real, imag} */,
  {32'hc357d978, 32'h00000000} /* (5, 4, 16) {real, imag} */,
  {32'hc499733a, 32'h00000000} /* (5, 4, 15) {real, imag} */,
  {32'hc4057b24, 32'h00000000} /* (5, 4, 14) {real, imag} */,
  {32'hc41d15aa, 32'h00000000} /* (5, 4, 13) {real, imag} */,
  {32'hc3c6f016, 32'h00000000} /* (5, 4, 12) {real, imag} */,
  {32'hc405f520, 32'h00000000} /* (5, 4, 11) {real, imag} */,
  {32'h412b2200, 32'h00000000} /* (5, 4, 10) {real, imag} */,
  {32'h440db87e, 32'h00000000} /* (5, 4, 9) {real, imag} */,
  {32'h43beaa20, 32'h00000000} /* (5, 4, 8) {real, imag} */,
  {32'h44a1b336, 32'h00000000} /* (5, 4, 7) {real, imag} */,
  {32'h45052bf0, 32'h00000000} /* (5, 4, 6) {real, imag} */,
  {32'h4501edf9, 32'h00000000} /* (5, 4, 5) {real, imag} */,
  {32'h4510a424, 32'h00000000} /* (5, 4, 4) {real, imag} */,
  {32'h44fb6b77, 32'h00000000} /* (5, 4, 3) {real, imag} */,
  {32'h452b0862, 32'h00000000} /* (5, 4, 2) {real, imag} */,
  {32'h4555d6aa, 32'h00000000} /* (5, 4, 1) {real, imag} */,
  {32'h456e440e, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'h453d0740, 32'h00000000} /* (5, 3, 31) {real, imag} */,
  {32'h4552755c, 32'h00000000} /* (5, 3, 30) {real, imag} */,
  {32'h453b1051, 32'h00000000} /* (5, 3, 29) {real, imag} */,
  {32'h451bc8f5, 32'h00000000} /* (5, 3, 28) {real, imag} */,
  {32'h4543907a, 32'h00000000} /* (5, 3, 27) {real, imag} */,
  {32'h453fb370, 32'h00000000} /* (5, 3, 26) {real, imag} */,
  {32'h45729b92, 32'h00000000} /* (5, 3, 25) {real, imag} */,
  {32'h45199f49, 32'h00000000} /* (5, 3, 24) {real, imag} */,
  {32'h45145b2c, 32'h00000000} /* (5, 3, 23) {real, imag} */,
  {32'h452680c5, 32'h00000000} /* (5, 3, 22) {real, imag} */,
  {32'h44fceb89, 32'h00000000} /* (5, 3, 21) {real, imag} */,
  {32'h450847ee, 32'h00000000} /* (5, 3, 20) {real, imag} */,
  {32'h44983c0a, 32'h00000000} /* (5, 3, 19) {real, imag} */,
  {32'h43a44e7c, 32'h00000000} /* (5, 3, 18) {real, imag} */,
  {32'h4400528a, 32'h00000000} /* (5, 3, 17) {real, imag} */,
  {32'hc456d02c, 32'h00000000} /* (5, 3, 16) {real, imag} */,
  {32'hc3f10af4, 32'h00000000} /* (5, 3, 15) {real, imag} */,
  {32'hc2dced90, 32'h00000000} /* (5, 3, 14) {real, imag} */,
  {32'hc3e25518, 32'h00000000} /* (5, 3, 13) {real, imag} */,
  {32'hc3baf3a8, 32'h00000000} /* (5, 3, 12) {real, imag} */,
  {32'hc298d000, 32'h00000000} /* (5, 3, 11) {real, imag} */,
  {32'h42020fe0, 32'h00000000} /* (5, 3, 10) {real, imag} */,
  {32'h43cfdb5c, 32'h00000000} /* (5, 3, 9) {real, imag} */,
  {32'h43bbec38, 32'h00000000} /* (5, 3, 8) {real, imag} */,
  {32'h44a1a0a1, 32'h00000000} /* (5, 3, 7) {real, imag} */,
  {32'h446e4a50, 32'h00000000} /* (5, 3, 6) {real, imag} */,
  {32'h44a3222b, 32'h00000000} /* (5, 3, 5) {real, imag} */,
  {32'h4529c08e, 32'h00000000} /* (5, 3, 4) {real, imag} */,
  {32'h44e3debe, 32'h00000000} /* (5, 3, 3) {real, imag} */,
  {32'h450497da, 32'h00000000} /* (5, 3, 2) {real, imag} */,
  {32'h45582f3a, 32'h00000000} /* (5, 3, 1) {real, imag} */,
  {32'h457f41cf, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'h4582da80, 32'h00000000} /* (5, 2, 31) {real, imag} */,
  {32'h458881cb, 32'h00000000} /* (5, 2, 30) {real, imag} */,
  {32'h455228da, 32'h00000000} /* (5, 2, 29) {real, imag} */,
  {32'h45224af4, 32'h00000000} /* (5, 2, 28) {real, imag} */,
  {32'h454d9fee, 32'h00000000} /* (5, 2, 27) {real, imag} */,
  {32'h45654320, 32'h00000000} /* (5, 2, 26) {real, imag} */,
  {32'h45405c2b, 32'h00000000} /* (5, 2, 25) {real, imag} */,
  {32'h454f876c, 32'h00000000} /* (5, 2, 24) {real, imag} */,
  {32'h45080893, 32'h00000000} /* (5, 2, 23) {real, imag} */,
  {32'h452d800b, 32'h00000000} /* (5, 2, 22) {real, imag} */,
  {32'h451a6a48, 32'h00000000} /* (5, 2, 21) {real, imag} */,
  {32'h44be654f, 32'h00000000} /* (5, 2, 20) {real, imag} */,
  {32'h4460a8ae, 32'h00000000} /* (5, 2, 19) {real, imag} */,
  {32'h441e7bfe, 32'h00000000} /* (5, 2, 18) {real, imag} */,
  {32'hc2933fe0, 32'h00000000} /* (5, 2, 17) {real, imag} */,
  {32'h4393d874, 32'h00000000} /* (5, 2, 16) {real, imag} */,
  {32'h442f8f3c, 32'h00000000} /* (5, 2, 15) {real, imag} */,
  {32'hc3856360, 32'h00000000} /* (5, 2, 14) {real, imag} */,
  {32'h43b8e6e4, 32'h00000000} /* (5, 2, 13) {real, imag} */,
  {32'h442ab5bd, 32'h00000000} /* (5, 2, 12) {real, imag} */,
  {32'h440d2e66, 32'h00000000} /* (5, 2, 11) {real, imag} */,
  {32'hc3e3024c, 32'h00000000} /* (5, 2, 10) {real, imag} */,
  {32'h442df3e0, 32'h00000000} /* (5, 2, 9) {real, imag} */,
  {32'h444532e8, 32'h00000000} /* (5, 2, 8) {real, imag} */,
  {32'h44a3b5f4, 32'h00000000} /* (5, 2, 7) {real, imag} */,
  {32'h44b3201e, 32'h00000000} /* (5, 2, 6) {real, imag} */,
  {32'h44b74656, 32'h00000000} /* (5, 2, 5) {real, imag} */,
  {32'h44cd9ae7, 32'h00000000} /* (5, 2, 4) {real, imag} */,
  {32'h45134970, 32'h00000000} /* (5, 2, 3) {real, imag} */,
  {32'h45425b70, 32'h00000000} /* (5, 2, 2) {real, imag} */,
  {32'h453e011a, 32'h00000000} /* (5, 2, 1) {real, imag} */,
  {32'h4539f7ac, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'h457b1027, 32'h00000000} /* (5, 1, 31) {real, imag} */,
  {32'h45814596, 32'h00000000} /* (5, 1, 30) {real, imag} */,
  {32'h458b80a8, 32'h00000000} /* (5, 1, 29) {real, imag} */,
  {32'h457fad22, 32'h00000000} /* (5, 1, 28) {real, imag} */,
  {32'h45549468, 32'h00000000} /* (5, 1, 27) {real, imag} */,
  {32'h4517a39d, 32'h00000000} /* (5, 1, 26) {real, imag} */,
  {32'h452a5471, 32'h00000000} /* (5, 1, 25) {real, imag} */,
  {32'h456c75b1, 32'h00000000} /* (5, 1, 24) {real, imag} */,
  {32'h454c41ac, 32'h00000000} /* (5, 1, 23) {real, imag} */,
  {32'h44c8e1e5, 32'h00000000} /* (5, 1, 22) {real, imag} */,
  {32'h44dbf1ec, 32'h00000000} /* (5, 1, 21) {real, imag} */,
  {32'h44a83700, 32'h00000000} /* (5, 1, 20) {real, imag} */,
  {32'h4484050f, 32'h00000000} /* (5, 1, 19) {real, imag} */,
  {32'hc3ff1368, 32'h00000000} /* (5, 1, 18) {real, imag} */,
  {32'hc40aac6c, 32'h00000000} /* (5, 1, 17) {real, imag} */,
  {32'h4486189c, 32'h00000000} /* (5, 1, 16) {real, imag} */,
  {32'h44211d6c, 32'h00000000} /* (5, 1, 15) {real, imag} */,
  {32'h442320a0, 32'h00000000} /* (5, 1, 14) {real, imag} */,
  {32'hc29aa5e0, 32'h00000000} /* (5, 1, 13) {real, imag} */,
  {32'h42fbc8d0, 32'h00000000} /* (5, 1, 12) {real, imag} */,
  {32'h4493a4b4, 32'h00000000} /* (5, 1, 11) {real, imag} */,
  {32'h445fd124, 32'h00000000} /* (5, 1, 10) {real, imag} */,
  {32'h4488113e, 32'h00000000} /* (5, 1, 9) {real, imag} */,
  {32'h44b40a2e, 32'h00000000} /* (5, 1, 8) {real, imag} */,
  {32'h44cc7a7b, 32'h00000000} /* (5, 1, 7) {real, imag} */,
  {32'h44d977a9, 32'h00000000} /* (5, 1, 6) {real, imag} */,
  {32'h448ebc32, 32'h00000000} /* (5, 1, 5) {real, imag} */,
  {32'h44ff2a0a, 32'h00000000} /* (5, 1, 4) {real, imag} */,
  {32'h450b8532, 32'h00000000} /* (5, 1, 3) {real, imag} */,
  {32'h4534ecc9, 32'h00000000} /* (5, 1, 2) {real, imag} */,
  {32'h4550c4db, 32'h00000000} /* (5, 1, 1) {real, imag} */,
  {32'h455e9e16, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'h4583ceaa, 32'h00000000} /* (5, 0, 31) {real, imag} */,
  {32'h45924180, 32'h00000000} /* (5, 0, 30) {real, imag} */,
  {32'h458e4fad, 32'h00000000} /* (5, 0, 29) {real, imag} */,
  {32'h458acb1a, 32'h00000000} /* (5, 0, 28) {real, imag} */,
  {32'h456bd21e, 32'h00000000} /* (5, 0, 27) {real, imag} */,
  {32'h4549e036, 32'h00000000} /* (5, 0, 26) {real, imag} */,
  {32'h454fdbeb, 32'h00000000} /* (5, 0, 25) {real, imag} */,
  {32'h456f325a, 32'h00000000} /* (5, 0, 24) {real, imag} */,
  {32'h453e4e4d, 32'h00000000} /* (5, 0, 23) {real, imag} */,
  {32'h451add7e, 32'h00000000} /* (5, 0, 22) {real, imag} */,
  {32'h4501c89a, 32'h00000000} /* (5, 0, 21) {real, imag} */,
  {32'h44d30077, 32'h00000000} /* (5, 0, 20) {real, imag} */,
  {32'h44904b1a, 32'h00000000} /* (5, 0, 19) {real, imag} */,
  {32'h433130e0, 32'h00000000} /* (5, 0, 18) {real, imag} */,
  {32'h43fb1f58, 32'h00000000} /* (5, 0, 17) {real, imag} */,
  {32'h43e24d2c, 32'h00000000} /* (5, 0, 16) {real, imag} */,
  {32'hc1055b00, 32'h00000000} /* (5, 0, 15) {real, imag} */,
  {32'h441235a8, 32'h00000000} /* (5, 0, 14) {real, imag} */,
  {32'h430527e0, 32'h00000000} /* (5, 0, 13) {real, imag} */,
  {32'h444479fa, 32'h00000000} /* (5, 0, 12) {real, imag} */,
  {32'h43aa6cd0, 32'h00000000} /* (5, 0, 11) {real, imag} */,
  {32'h441571f2, 32'h00000000} /* (5, 0, 10) {real, imag} */,
  {32'h437234f0, 32'h00000000} /* (5, 0, 9) {real, imag} */,
  {32'h447137b0, 32'h00000000} /* (5, 0, 8) {real, imag} */,
  {32'h445b43dc, 32'h00000000} /* (5, 0, 7) {real, imag} */,
  {32'h448af1d0, 32'h00000000} /* (5, 0, 6) {real, imag} */,
  {32'h44df6044, 32'h00000000} /* (5, 0, 5) {real, imag} */,
  {32'h44edf055, 32'h00000000} /* (5, 0, 4) {real, imag} */,
  {32'h4540f02f, 32'h00000000} /* (5, 0, 3) {real, imag} */,
  {32'h45512cd3, 32'h00000000} /* (5, 0, 2) {real, imag} */,
  {32'h4563f35f, 32'h00000000} /* (5, 0, 1) {real, imag} */,
  {32'h456d748c, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'h44bb8a80, 32'h00000000} /* (4, 31, 31) {real, imag} */,
  {32'h44cbdfab, 32'h00000000} /* (4, 31, 30) {real, imag} */,
  {32'h44c10338, 32'h00000000} /* (4, 31, 29) {real, imag} */,
  {32'h444ef230, 32'h00000000} /* (4, 31, 28) {real, imag} */,
  {32'h430b63d8, 32'h00000000} /* (4, 31, 27) {real, imag} */,
  {32'hc4074366, 32'h00000000} /* (4, 31, 26) {real, imag} */,
  {32'hc34b57c1, 32'h00000000} /* (4, 31, 25) {real, imag} */,
  {32'hc437d18d, 32'h00000000} /* (4, 31, 24) {real, imag} */,
  {32'h43f7101e, 32'h00000000} /* (4, 31, 23) {real, imag} */,
  {32'h440b5571, 32'h00000000} /* (4, 31, 22) {real, imag} */,
  {32'h442a80b1, 32'h00000000} /* (4, 31, 21) {real, imag} */,
  {32'h44ba903a, 32'h00000000} /* (4, 31, 20) {real, imag} */,
  {32'h44e40cd3, 32'h00000000} /* (4, 31, 19) {real, imag} */,
  {32'h44a0cbcc, 32'h00000000} /* (4, 31, 18) {real, imag} */,
  {32'h44d41244, 32'h00000000} /* (4, 31, 17) {real, imag} */,
  {32'h44a710cf, 32'h00000000} /* (4, 31, 16) {real, imag} */,
  {32'h44c2902c, 32'h00000000} /* (4, 31, 15) {real, imag} */,
  {32'h44c2ad0d, 32'h00000000} /* (4, 31, 14) {real, imag} */,
  {32'h452caf2c, 32'h00000000} /* (4, 31, 13) {real, imag} */,
  {32'h4506dbe0, 32'h00000000} /* (4, 31, 12) {real, imag} */,
  {32'h44bc3693, 32'h00000000} /* (4, 31, 11) {real, imag} */,
  {32'h43d213eb, 32'h00000000} /* (4, 31, 10) {real, imag} */,
  {32'h43658359, 32'h00000000} /* (4, 31, 9) {real, imag} */,
  {32'h43bd131e, 32'h00000000} /* (4, 31, 8) {real, imag} */,
  {32'h43572b25, 32'h00000000} /* (4, 31, 7) {real, imag} */,
  {32'hc35eea24, 32'h00000000} /* (4, 31, 6) {real, imag} */,
  {32'h42899958, 32'h00000000} /* (4, 31, 5) {real, imag} */,
  {32'h43d18c5a, 32'h00000000} /* (4, 31, 4) {real, imag} */,
  {32'h43bb8e8c, 32'h00000000} /* (4, 31, 3) {real, imag} */,
  {32'h446aba50, 32'h00000000} /* (4, 31, 2) {real, imag} */,
  {32'h44ac858c, 32'h00000000} /* (4, 31, 1) {real, imag} */,
  {32'h44b39405, 32'h00000000} /* (4, 31, 0) {real, imag} */,
  {32'h4488e3f8, 32'h00000000} /* (4, 30, 31) {real, imag} */,
  {32'h43d80196, 32'h00000000} /* (4, 30, 30) {real, imag} */,
  {32'h44833cac, 32'h00000000} /* (4, 30, 29) {real, imag} */,
  {32'h437becc8, 32'h00000000} /* (4, 30, 28) {real, imag} */,
  {32'hc39a1e18, 32'h00000000} /* (4, 30, 27) {real, imag} */,
  {32'hc4a7f438, 32'h00000000} /* (4, 30, 26) {real, imag} */,
  {32'hc4608ebc, 32'h00000000} /* (4, 30, 25) {real, imag} */,
  {32'hc449cb4d, 32'h00000000} /* (4, 30, 24) {real, imag} */,
  {32'hc3fe1d18, 32'h00000000} /* (4, 30, 23) {real, imag} */,
  {32'h4305cc1c, 32'h00000000} /* (4, 30, 22) {real, imag} */,
  {32'h4443558e, 32'h00000000} /* (4, 30, 21) {real, imag} */,
  {32'h44d3fb0d, 32'h00000000} /* (4, 30, 20) {real, imag} */,
  {32'h451e2816, 32'h00000000} /* (4, 30, 19) {real, imag} */,
  {32'h4511ba92, 32'h00000000} /* (4, 30, 18) {real, imag} */,
  {32'h451b6c29, 32'h00000000} /* (4, 30, 17) {real, imag} */,
  {32'h4502165c, 32'h00000000} /* (4, 30, 16) {real, imag} */,
  {32'h451fcfa9, 32'h00000000} /* (4, 30, 15) {real, imag} */,
  {32'h4504952f, 32'h00000000} /* (4, 30, 14) {real, imag} */,
  {32'h453af6c0, 32'h00000000} /* (4, 30, 13) {real, imag} */,
  {32'h4520dec6, 32'h00000000} /* (4, 30, 12) {real, imag} */,
  {32'h44fe3b48, 32'h00000000} /* (4, 30, 11) {real, imag} */,
  {32'h4366cdf0, 32'h00000000} /* (4, 30, 10) {real, imag} */,
  {32'hc3ccb870, 32'h00000000} /* (4, 30, 9) {real, imag} */,
  {32'hc3a54afe, 32'h00000000} /* (4, 30, 8) {real, imag} */,
  {32'hc486badc, 32'h00000000} /* (4, 30, 7) {real, imag} */,
  {32'hc473caed, 32'h00000000} /* (4, 30, 6) {real, imag} */,
  {32'hc46ea526, 32'h00000000} /* (4, 30, 5) {real, imag} */,
  {32'hc3b0e9b4, 32'h00000000} /* (4, 30, 4) {real, imag} */,
  {32'h41c6fe40, 32'h00000000} /* (4, 30, 3) {real, imag} */,
  {32'h443619da, 32'h00000000} /* (4, 30, 2) {real, imag} */,
  {32'h4404a080, 32'h00000000} /* (4, 30, 1) {real, imag} */,
  {32'h449bce3a, 32'h00000000} /* (4, 30, 0) {real, imag} */,
  {32'h446cd837, 32'h00000000} /* (4, 29, 31) {real, imag} */,
  {32'hc315b9e0, 32'h00000000} /* (4, 29, 30) {real, imag} */,
  {32'hc2757ce0, 32'h00000000} /* (4, 29, 29) {real, imag} */,
  {32'h4370a548, 32'h00000000} /* (4, 29, 28) {real, imag} */,
  {32'h42da9878, 32'h00000000} /* (4, 29, 27) {real, imag} */,
  {32'hc4797d14, 32'h00000000} /* (4, 29, 26) {real, imag} */,
  {32'hc4927c45, 32'h00000000} /* (4, 29, 25) {real, imag} */,
  {32'hc47d7540, 32'h00000000} /* (4, 29, 24) {real, imag} */,
  {32'hc49dda43, 32'h00000000} /* (4, 29, 23) {real, imag} */,
  {32'hc37d855e, 32'h00000000} /* (4, 29, 22) {real, imag} */,
  {32'h44373886, 32'h00000000} /* (4, 29, 21) {real, imag} */,
  {32'h4500a3cf, 32'h00000000} /* (4, 29, 20) {real, imag} */,
  {32'h453ad6e8, 32'h00000000} /* (4, 29, 19) {real, imag} */,
  {32'h4509cc6c, 32'h00000000} /* (4, 29, 18) {real, imag} */,
  {32'h456479b4, 32'h00000000} /* (4, 29, 17) {real, imag} */,
  {32'h45674b30, 32'h00000000} /* (4, 29, 16) {real, imag} */,
  {32'h453b07ec, 32'h00000000} /* (4, 29, 15) {real, imag} */,
  {32'h450a6b62, 32'h00000000} /* (4, 29, 14) {real, imag} */,
  {32'h44ffa12f, 32'h00000000} /* (4, 29, 13) {real, imag} */,
  {32'h452370c6, 32'h00000000} /* (4, 29, 12) {real, imag} */,
  {32'h45041c77, 32'h00000000} /* (4, 29, 11) {real, imag} */,
  {32'hc44bf0cc, 32'h00000000} /* (4, 29, 10) {real, imag} */,
  {32'hc45f5a12, 32'h00000000} /* (4, 29, 9) {real, imag} */,
  {32'hc450bf12, 32'h00000000} /* (4, 29, 8) {real, imag} */,
  {32'hc4b12c29, 32'h00000000} /* (4, 29, 7) {real, imag} */,
  {32'hc41a28c6, 32'h00000000} /* (4, 29, 6) {real, imag} */,
  {32'hc47611b8, 32'h00000000} /* (4, 29, 5) {real, imag} */,
  {32'hc46e4288, 32'h00000000} /* (4, 29, 4) {real, imag} */,
  {32'h43a20f6c, 32'h00000000} /* (4, 29, 3) {real, imag} */,
  {32'h444f393a, 32'h00000000} /* (4, 29, 2) {real, imag} */,
  {32'h4357d478, 32'h00000000} /* (4, 29, 1) {real, imag} */,
  {32'h43f6ee40, 32'h00000000} /* (4, 29, 0) {real, imag} */,
  {32'h44925559, 32'h00000000} /* (4, 28, 31) {real, imag} */,
  {32'h4399d040, 32'h00000000} /* (4, 28, 30) {real, imag} */,
  {32'hc4730df9, 32'h00000000} /* (4, 28, 29) {real, imag} */,
  {32'h41ed8540, 32'h00000000} /* (4, 28, 28) {real, imag} */,
  {32'hc3ff0c8c, 32'h00000000} /* (4, 28, 27) {real, imag} */,
  {32'hc4827a2a, 32'h00000000} /* (4, 28, 26) {real, imag} */,
  {32'hc4827a28, 32'h00000000} /* (4, 28, 25) {real, imag} */,
  {32'hc4a59e17, 32'h00000000} /* (4, 28, 24) {real, imag} */,
  {32'hc4481b2a, 32'h00000000} /* (4, 28, 23) {real, imag} */,
  {32'h42841258, 32'h00000000} /* (4, 28, 22) {real, imag} */,
  {32'h44fc9d46, 32'h00000000} /* (4, 28, 21) {real, imag} */,
  {32'h453ad114, 32'h00000000} /* (4, 28, 20) {real, imag} */,
  {32'h453c53d1, 32'h00000000} /* (4, 28, 19) {real, imag} */,
  {32'h4514361e, 32'h00000000} /* (4, 28, 18) {real, imag} */,
  {32'h452afb8e, 32'h00000000} /* (4, 28, 17) {real, imag} */,
  {32'h453343a7, 32'h00000000} /* (4, 28, 16) {real, imag} */,
  {32'h45040ac6, 32'h00000000} /* (4, 28, 15) {real, imag} */,
  {32'h44f35d40, 32'h00000000} /* (4, 28, 14) {real, imag} */,
  {32'h4523f810, 32'h00000000} /* (4, 28, 13) {real, imag} */,
  {32'h450b3ff4, 32'h00000000} /* (4, 28, 12) {real, imag} */,
  {32'h452b5ea2, 32'h00000000} /* (4, 28, 11) {real, imag} */,
  {32'h4463206b, 32'h00000000} /* (4, 28, 10) {real, imag} */,
  {32'hc4a9ffc0, 32'h00000000} /* (4, 28, 9) {real, imag} */,
  {32'hc4c07669, 32'h00000000} /* (4, 28, 8) {real, imag} */,
  {32'hc4032b46, 32'h00000000} /* (4, 28, 7) {real, imag} */,
  {32'hc43c1c91, 32'h00000000} /* (4, 28, 6) {real, imag} */,
  {32'hc3fc8eee, 32'h00000000} /* (4, 28, 5) {real, imag} */,
  {32'hc44c1e86, 32'h00000000} /* (4, 28, 4) {real, imag} */,
  {32'hc428ba4c, 32'h00000000} /* (4, 28, 3) {real, imag} */,
  {32'hc2f09e70, 32'h00000000} /* (4, 28, 2) {real, imag} */,
  {32'h4398c964, 32'h00000000} /* (4, 28, 1) {real, imag} */,
  {32'h443a36e4, 32'h00000000} /* (4, 28, 0) {real, imag} */,
  {32'h4436cfea, 32'h00000000} /* (4, 27, 31) {real, imag} */,
  {32'hc3371e08, 32'h00000000} /* (4, 27, 30) {real, imag} */,
  {32'h43535190, 32'h00000000} /* (4, 27, 29) {real, imag} */,
  {32'hc48682e4, 32'h00000000} /* (4, 27, 28) {real, imag} */,
  {32'hc47cce05, 32'h00000000} /* (4, 27, 27) {real, imag} */,
  {32'hc472608f, 32'h00000000} /* (4, 27, 26) {real, imag} */,
  {32'hc4c2e596, 32'h00000000} /* (4, 27, 25) {real, imag} */,
  {32'hc4feac20, 32'h00000000} /* (4, 27, 24) {real, imag} */,
  {32'hc4003bb0, 32'h00000000} /* (4, 27, 23) {real, imag} */,
  {32'hc420705e, 32'h00000000} /* (4, 27, 22) {real, imag} */,
  {32'h443cd09b, 32'h00000000} /* (4, 27, 21) {real, imag} */,
  {32'h4560275a, 32'h00000000} /* (4, 27, 20) {real, imag} */,
  {32'h4546ece6, 32'h00000000} /* (4, 27, 19) {real, imag} */,
  {32'h4579cefa, 32'h00000000} /* (4, 27, 18) {real, imag} */,
  {32'h45331b90, 32'h00000000} /* (4, 27, 17) {real, imag} */,
  {32'h4511c170, 32'h00000000} /* (4, 27, 16) {real, imag} */,
  {32'h4577ddca, 32'h00000000} /* (4, 27, 15) {real, imag} */,
  {32'h451b5a36, 32'h00000000} /* (4, 27, 14) {real, imag} */,
  {32'h451fe635, 32'h00000000} /* (4, 27, 13) {real, imag} */,
  {32'h4542bc46, 32'h00000000} /* (4, 27, 12) {real, imag} */,
  {32'h453945db, 32'h00000000} /* (4, 27, 11) {real, imag} */,
  {32'h4311d4e4, 32'h00000000} /* (4, 27, 10) {real, imag} */,
  {32'hc429f778, 32'h00000000} /* (4, 27, 9) {real, imag} */,
  {32'hc46325a4, 32'h00000000} /* (4, 27, 8) {real, imag} */,
  {32'hc3d95f47, 32'h00000000} /* (4, 27, 7) {real, imag} */,
  {32'hc48f9c24, 32'h00000000} /* (4, 27, 6) {real, imag} */,
  {32'hc3f85c76, 32'h00000000} /* (4, 27, 5) {real, imag} */,
  {32'h42b31600, 32'h00000000} /* (4, 27, 4) {real, imag} */,
  {32'hc43129c8, 32'h00000000} /* (4, 27, 3) {real, imag} */,
  {32'hc383ec70, 32'h00000000} /* (4, 27, 2) {real, imag} */,
  {32'hc3b62f6c, 32'h00000000} /* (4, 27, 1) {real, imag} */,
  {32'hc1a3ea40, 32'h00000000} /* (4, 27, 0) {real, imag} */,
  {32'h43beaafc, 32'h00000000} /* (4, 26, 31) {real, imag} */,
  {32'hc3c41df0, 32'h00000000} /* (4, 26, 30) {real, imag} */,
  {32'hc402d1aa, 32'h00000000} /* (4, 26, 29) {real, imag} */,
  {32'hc4261c72, 32'h00000000} /* (4, 26, 28) {real, imag} */,
  {32'hc40eef30, 32'h00000000} /* (4, 26, 27) {real, imag} */,
  {32'hc4d09cb7, 32'h00000000} /* (4, 26, 26) {real, imag} */,
  {32'hc4cc9806, 32'h00000000} /* (4, 26, 25) {real, imag} */,
  {32'hc5167aa2, 32'h00000000} /* (4, 26, 24) {real, imag} */,
  {32'hc4f10fea, 32'h00000000} /* (4, 26, 23) {real, imag} */,
  {32'hc3a68256, 32'h00000000} /* (4, 26, 22) {real, imag} */,
  {32'h444d81c0, 32'h00000000} /* (4, 26, 21) {real, imag} */,
  {32'h4505cad5, 32'h00000000} /* (4, 26, 20) {real, imag} */,
  {32'h453823e4, 32'h00000000} /* (4, 26, 19) {real, imag} */,
  {32'h45458d4c, 32'h00000000} /* (4, 26, 18) {real, imag} */,
  {32'h455c3494, 32'h00000000} /* (4, 26, 17) {real, imag} */,
  {32'h45316a67, 32'h00000000} /* (4, 26, 16) {real, imag} */,
  {32'h45630476, 32'h00000000} /* (4, 26, 15) {real, imag} */,
  {32'h456a3af4, 32'h00000000} /* (4, 26, 14) {real, imag} */,
  {32'h452357a6, 32'h00000000} /* (4, 26, 13) {real, imag} */,
  {32'h453c2ed6, 32'h00000000} /* (4, 26, 12) {real, imag} */,
  {32'h44d0434c, 32'h00000000} /* (4, 26, 11) {real, imag} */,
  {32'h439963f4, 32'h00000000} /* (4, 26, 10) {real, imag} */,
  {32'hc42089f7, 32'h00000000} /* (4, 26, 9) {real, imag} */,
  {32'hc3f69b10, 32'h00000000} /* (4, 26, 8) {real, imag} */,
  {32'hc3a2e7c2, 32'h00000000} /* (4, 26, 7) {real, imag} */,
  {32'hc3b6d4aa, 32'h00000000} /* (4, 26, 6) {real, imag} */,
  {32'hc3f29739, 32'h00000000} /* (4, 26, 5) {real, imag} */,
  {32'hc43f0fdf, 32'h00000000} /* (4, 26, 4) {real, imag} */,
  {32'hc31afa78, 32'h00000000} /* (4, 26, 3) {real, imag} */,
  {32'hc41108e6, 32'h00000000} /* (4, 26, 2) {real, imag} */,
  {32'hc38a9eec, 32'h00000000} /* (4, 26, 1) {real, imag} */,
  {32'h43e040b8, 32'h00000000} /* (4, 26, 0) {real, imag} */,
  {32'hc3dd468c, 32'h00000000} /* (4, 25, 31) {real, imag} */,
  {32'hc46d78e6, 32'h00000000} /* (4, 25, 30) {real, imag} */,
  {32'hc4795d0e, 32'h00000000} /* (4, 25, 29) {real, imag} */,
  {32'hc4b4202c, 32'h00000000} /* (4, 25, 28) {real, imag} */,
  {32'hc4dbeadd, 32'h00000000} /* (4, 25, 27) {real, imag} */,
  {32'hc4eac974, 32'h00000000} /* (4, 25, 26) {real, imag} */,
  {32'hc52d9b68, 32'h00000000} /* (4, 25, 25) {real, imag} */,
  {32'hc4df8b95, 32'h00000000} /* (4, 25, 24) {real, imag} */,
  {32'hc4eba8d0, 32'h00000000} /* (4, 25, 23) {real, imag} */,
  {32'hc4a31380, 32'h00000000} /* (4, 25, 22) {real, imag} */,
  {32'h42941480, 32'h00000000} /* (4, 25, 21) {real, imag} */,
  {32'h454d36c6, 32'h00000000} /* (4, 25, 20) {real, imag} */,
  {32'h4553f45e, 32'h00000000} /* (4, 25, 19) {real, imag} */,
  {32'h453f71ac, 32'h00000000} /* (4, 25, 18) {real, imag} */,
  {32'h45450d58, 32'h00000000} /* (4, 25, 17) {real, imag} */,
  {32'h4541d296, 32'h00000000} /* (4, 25, 16) {real, imag} */,
  {32'h454bb62c, 32'h00000000} /* (4, 25, 15) {real, imag} */,
  {32'h451d93f0, 32'h00000000} /* (4, 25, 14) {real, imag} */,
  {32'h453f4dda, 32'h00000000} /* (4, 25, 13) {real, imag} */,
  {32'h44e43f50, 32'h00000000} /* (4, 25, 12) {real, imag} */,
  {32'h4511ef2b, 32'h00000000} /* (4, 25, 11) {real, imag} */,
  {32'h4357aa94, 32'h00000000} /* (4, 25, 10) {real, imag} */,
  {32'hc3dd9184, 32'h00000000} /* (4, 25, 9) {real, imag} */,
  {32'hc4f86135, 32'h00000000} /* (4, 25, 8) {real, imag} */,
  {32'hc48052e2, 32'h00000000} /* (4, 25, 7) {real, imag} */,
  {32'hc41ca819, 32'h00000000} /* (4, 25, 6) {real, imag} */,
  {32'hc5090147, 32'h00000000} /* (4, 25, 5) {real, imag} */,
  {32'hc4c28000, 32'h00000000} /* (4, 25, 4) {real, imag} */,
  {32'hc448d670, 32'h00000000} /* (4, 25, 3) {real, imag} */,
  {32'hc4b95aa4, 32'h00000000} /* (4, 25, 2) {real, imag} */,
  {32'hc40e93ce, 32'h00000000} /* (4, 25, 1) {real, imag} */,
  {32'hc330d098, 32'h00000000} /* (4, 25, 0) {real, imag} */,
  {32'hc3a677b8, 32'h00000000} /* (4, 24, 31) {real, imag} */,
  {32'hc49be776, 32'h00000000} /* (4, 24, 30) {real, imag} */,
  {32'hc4fef988, 32'h00000000} /* (4, 24, 29) {real, imag} */,
  {32'hc4ec0ccb, 32'h00000000} /* (4, 24, 28) {real, imag} */,
  {32'hc4ba11ff, 32'h00000000} /* (4, 24, 27) {real, imag} */,
  {32'hc510159c, 32'h00000000} /* (4, 24, 26) {real, imag} */,
  {32'hc4def374, 32'h00000000} /* (4, 24, 25) {real, imag} */,
  {32'hc4a61c44, 32'h00000000} /* (4, 24, 24) {real, imag} */,
  {32'hc4864d12, 32'h00000000} /* (4, 24, 23) {real, imag} */,
  {32'hc3b6bec1, 32'h00000000} /* (4, 24, 22) {real, imag} */,
  {32'h44102eb0, 32'h00000000} /* (4, 24, 21) {real, imag} */,
  {32'h455ab170, 32'h00000000} /* (4, 24, 20) {real, imag} */,
  {32'h4578b3b1, 32'h00000000} /* (4, 24, 19) {real, imag} */,
  {32'h45821f8e, 32'h00000000} /* (4, 24, 18) {real, imag} */,
  {32'h454e37b3, 32'h00000000} /* (4, 24, 17) {real, imag} */,
  {32'h4566c206, 32'h00000000} /* (4, 24, 16) {real, imag} */,
  {32'h4581d0cc, 32'h00000000} /* (4, 24, 15) {real, imag} */,
  {32'h4544e7d7, 32'h00000000} /* (4, 24, 14) {real, imag} */,
  {32'h452ea178, 32'h00000000} /* (4, 24, 13) {real, imag} */,
  {32'h4508002a, 32'h00000000} /* (4, 24, 12) {real, imag} */,
  {32'h44f3fddf, 32'h00000000} /* (4, 24, 11) {real, imag} */,
  {32'hc396f864, 32'h00000000} /* (4, 24, 10) {real, imag} */,
  {32'hc4576620, 32'h00000000} /* (4, 24, 9) {real, imag} */,
  {32'hc4b48db4, 32'h00000000} /* (4, 24, 8) {real, imag} */,
  {32'hc444783b, 32'h00000000} /* (4, 24, 7) {real, imag} */,
  {32'hc4949ba3, 32'h00000000} /* (4, 24, 6) {real, imag} */,
  {32'hc48505eb, 32'h00000000} /* (4, 24, 5) {real, imag} */,
  {32'hc449b330, 32'h00000000} /* (4, 24, 4) {real, imag} */,
  {32'hc40b2f24, 32'h00000000} /* (4, 24, 3) {real, imag} */,
  {32'hc4efdcbb, 32'h00000000} /* (4, 24, 2) {real, imag} */,
  {32'hc50771ef, 32'h00000000} /* (4, 24, 1) {real, imag} */,
  {32'hc47fdf70, 32'h00000000} /* (4, 24, 0) {real, imag} */,
  {32'hc4925d0d, 32'h00000000} /* (4, 23, 31) {real, imag} */,
  {32'hc4cd5dd5, 32'h00000000} /* (4, 23, 30) {real, imag} */,
  {32'hc4b68eb6, 32'h00000000} /* (4, 23, 29) {real, imag} */,
  {32'hc4fd2674, 32'h00000000} /* (4, 23, 28) {real, imag} */,
  {32'hc5091f77, 32'h00000000} /* (4, 23, 27) {real, imag} */,
  {32'hc4a4831c, 32'h00000000} /* (4, 23, 26) {real, imag} */,
  {32'hc4b74eca, 32'h00000000} /* (4, 23, 25) {real, imag} */,
  {32'hc4c13c9e, 32'h00000000} /* (4, 23, 24) {real, imag} */,
  {32'hc42746b0, 32'h00000000} /* (4, 23, 23) {real, imag} */,
  {32'hc2cbcca8, 32'h00000000} /* (4, 23, 22) {real, imag} */,
  {32'h449b38b4, 32'h00000000} /* (4, 23, 21) {real, imag} */,
  {32'h454f8caf, 32'h00000000} /* (4, 23, 20) {real, imag} */,
  {32'h4555bf92, 32'h00000000} /* (4, 23, 19) {real, imag} */,
  {32'h45864252, 32'h00000000} /* (4, 23, 18) {real, imag} */,
  {32'h45825dde, 32'h00000000} /* (4, 23, 17) {real, imag} */,
  {32'h454bc241, 32'h00000000} /* (4, 23, 16) {real, imag} */,
  {32'h453f27ba, 32'h00000000} /* (4, 23, 15) {real, imag} */,
  {32'h45533906, 32'h00000000} /* (4, 23, 14) {real, imag} */,
  {32'h45173047, 32'h00000000} /* (4, 23, 13) {real, imag} */,
  {32'h44bd20e0, 32'h00000000} /* (4, 23, 12) {real, imag} */,
  {32'h44f7111e, 32'h00000000} /* (4, 23, 11) {real, imag} */,
  {32'hc2c5e658, 32'h00000000} /* (4, 23, 10) {real, imag} */,
  {32'hc4db5726, 32'h00000000} /* (4, 23, 9) {real, imag} */,
  {32'hc5054edf, 32'h00000000} /* (4, 23, 8) {real, imag} */,
  {32'hc4bcf57c, 32'h00000000} /* (4, 23, 7) {real, imag} */,
  {32'hc4801c5a, 32'h00000000} /* (4, 23, 6) {real, imag} */,
  {32'hc44714a6, 32'h00000000} /* (4, 23, 5) {real, imag} */,
  {32'hc4269d7c, 32'h00000000} /* (4, 23, 4) {real, imag} */,
  {32'hc4c44438, 32'h00000000} /* (4, 23, 3) {real, imag} */,
  {32'hc48151ca, 32'h00000000} /* (4, 23, 2) {real, imag} */,
  {32'hc4ea8194, 32'h00000000} /* (4, 23, 1) {real, imag} */,
  {32'hc495a292, 32'h00000000} /* (4, 23, 0) {real, imag} */,
  {32'hc3dc273c, 32'h00000000} /* (4, 22, 31) {real, imag} */,
  {32'hc4ed9e09, 32'h00000000} /* (4, 22, 30) {real, imag} */,
  {32'hc4887b84, 32'h00000000} /* (4, 22, 29) {real, imag} */,
  {32'hc49cd8ee, 32'h00000000} /* (4, 22, 28) {real, imag} */,
  {32'hc4acee0c, 32'h00000000} /* (4, 22, 27) {real, imag} */,
  {32'hc405a2ec, 32'h00000000} /* (4, 22, 26) {real, imag} */,
  {32'hc4ab1860, 32'h00000000} /* (4, 22, 25) {real, imag} */,
  {32'hc49789ce, 32'h00000000} /* (4, 22, 24) {real, imag} */,
  {32'hc4a83a8d, 32'h00000000} /* (4, 22, 23) {real, imag} */,
  {32'h438a8d9e, 32'h00000000} /* (4, 22, 22) {real, imag} */,
  {32'h441d1892, 32'h00000000} /* (4, 22, 21) {real, imag} */,
  {32'h45437b1b, 32'h00000000} /* (4, 22, 20) {real, imag} */,
  {32'h454bc641, 32'h00000000} /* (4, 22, 19) {real, imag} */,
  {32'h4551e2ec, 32'h00000000} /* (4, 22, 18) {real, imag} */,
  {32'h455c76ba, 32'h00000000} /* (4, 22, 17) {real, imag} */,
  {32'h44f2640b, 32'h00000000} /* (4, 22, 16) {real, imag} */,
  {32'h450d2aa6, 32'h00000000} /* (4, 22, 15) {real, imag} */,
  {32'h452e638f, 32'h00000000} /* (4, 22, 14) {real, imag} */,
  {32'h44e78f86, 32'h00000000} /* (4, 22, 13) {real, imag} */,
  {32'h44bc9566, 32'h00000000} /* (4, 22, 12) {real, imag} */,
  {32'h449391aa, 32'h00000000} /* (4, 22, 11) {real, imag} */,
  {32'hc4438b6c, 32'h00000000} /* (4, 22, 10) {real, imag} */,
  {32'hc4bc0704, 32'h00000000} /* (4, 22, 9) {real, imag} */,
  {32'hc4a7af4e, 32'h00000000} /* (4, 22, 8) {real, imag} */,
  {32'hc4390fba, 32'h00000000} /* (4, 22, 7) {real, imag} */,
  {32'hc4af0c76, 32'h00000000} /* (4, 22, 6) {real, imag} */,
  {32'hc497b161, 32'h00000000} /* (4, 22, 5) {real, imag} */,
  {32'hc48e2d06, 32'h00000000} /* (4, 22, 4) {real, imag} */,
  {32'hc4a012ee, 32'h00000000} /* (4, 22, 3) {real, imag} */,
  {32'hc42e653a, 32'h00000000} /* (4, 22, 2) {real, imag} */,
  {32'hc4eb26bc, 32'h00000000} /* (4, 22, 1) {real, imag} */,
  {32'hc47fb38e, 32'h00000000} /* (4, 22, 0) {real, imag} */,
  {32'h42e1db48, 32'h00000000} /* (4, 21, 31) {real, imag} */,
  {32'h44020553, 32'h00000000} /* (4, 21, 30) {real, imag} */,
  {32'hc409d0ff, 32'h00000000} /* (4, 21, 29) {real, imag} */,
  {32'hc21ba7ac, 32'h00000000} /* (4, 21, 28) {real, imag} */,
  {32'h441dab6a, 32'h00000000} /* (4, 21, 27) {real, imag} */,
  {32'hc49d6aa8, 32'h00000000} /* (4, 21, 26) {real, imag} */,
  {32'h448dad59, 32'h00000000} /* (4, 21, 25) {real, imag} */,
  {32'h443d2b72, 32'h00000000} /* (4, 21, 24) {real, imag} */,
  {32'h42aba6d0, 32'h00000000} /* (4, 21, 23) {real, imag} */,
  {32'h443bc1fd, 32'h00000000} /* (4, 21, 22) {real, imag} */,
  {32'h447234ce, 32'h00000000} /* (4, 21, 21) {real, imag} */,
  {32'h44b486fb, 32'h00000000} /* (4, 21, 20) {real, imag} */,
  {32'h450fb3d6, 32'h00000000} /* (4, 21, 19) {real, imag} */,
  {32'h44d6dc89, 32'h00000000} /* (4, 21, 18) {real, imag} */,
  {32'h44e5313c, 32'h00000000} /* (4, 21, 17) {real, imag} */,
  {32'h442f9d04, 32'h00000000} /* (4, 21, 16) {real, imag} */,
  {32'h44881bcc, 32'h00000000} /* (4, 21, 15) {real, imag} */,
  {32'h44e984c6, 32'h00000000} /* (4, 21, 14) {real, imag} */,
  {32'h44ab6f36, 32'h00000000} /* (4, 21, 13) {real, imag} */,
  {32'h4405cbbb, 32'h00000000} /* (4, 21, 12) {real, imag} */,
  {32'h4454bf82, 32'h00000000} /* (4, 21, 11) {real, imag} */,
  {32'h442285f7, 32'h00000000} /* (4, 21, 10) {real, imag} */,
  {32'h43157932, 32'h00000000} /* (4, 21, 9) {real, imag} */,
  {32'h4359396a, 32'h00000000} /* (4, 21, 8) {real, imag} */,
  {32'hc38c3bf4, 32'h00000000} /* (4, 21, 7) {real, imag} */,
  {32'hc3f89dca, 32'h00000000} /* (4, 21, 6) {real, imag} */,
  {32'h43498280, 32'h00000000} /* (4, 21, 5) {real, imag} */,
  {32'hc2d727d0, 32'h00000000} /* (4, 21, 4) {real, imag} */,
  {32'hc47cce3e, 32'h00000000} /* (4, 21, 3) {real, imag} */,
  {32'h43024d20, 32'h00000000} /* (4, 21, 2) {real, imag} */,
  {32'hc41050d7, 32'h00000000} /* (4, 21, 1) {real, imag} */,
  {32'hc3bb7599, 32'h00000000} /* (4, 21, 0) {real, imag} */,
  {32'h44f57e4e, 32'h00000000} /* (4, 20, 31) {real, imag} */,
  {32'h45342fe2, 32'h00000000} /* (4, 20, 30) {real, imag} */,
  {32'h4501167e, 32'h00000000} /* (4, 20, 29) {real, imag} */,
  {32'h4539950e, 32'h00000000} /* (4, 20, 28) {real, imag} */,
  {32'h450b9aca, 32'h00000000} /* (4, 20, 27) {real, imag} */,
  {32'h44e289bf, 32'h00000000} /* (4, 20, 26) {real, imag} */,
  {32'h4533aaca, 32'h00000000} /* (4, 20, 25) {real, imag} */,
  {32'h452c8290, 32'h00000000} /* (4, 20, 24) {real, imag} */,
  {32'h45453c4f, 32'h00000000} /* (4, 20, 23) {real, imag} */,
  {32'h4492d1d8, 32'h00000000} /* (4, 20, 22) {real, imag} */,
  {32'h4493e602, 32'h00000000} /* (4, 20, 21) {real, imag} */,
  {32'hc0f8d800, 32'h00000000} /* (4, 20, 20) {real, imag} */,
  {32'h43e0bf89, 32'h00000000} /* (4, 20, 19) {real, imag} */,
  {32'hc15ae0c0, 32'h00000000} /* (4, 20, 18) {real, imag} */,
  {32'hc4091e25, 32'h00000000} /* (4, 20, 17) {real, imag} */,
  {32'hc412162a, 32'h00000000} /* (4, 20, 16) {real, imag} */,
  {32'hc3a34762, 32'h00000000} /* (4, 20, 15) {real, imag} */,
  {32'hc3e8f58c, 32'h00000000} /* (4, 20, 14) {real, imag} */,
  {32'hc4391c0e, 32'h00000000} /* (4, 20, 13) {real, imag} */,
  {32'hc471bc43, 32'h00000000} /* (4, 20, 12) {real, imag} */,
  {32'h43cd26f6, 32'h00000000} /* (4, 20, 11) {real, imag} */,
  {32'h44dd90f7, 32'h00000000} /* (4, 20, 10) {real, imag} */,
  {32'h44a1d32f, 32'h00000000} /* (4, 20, 9) {real, imag} */,
  {32'h449e9655, 32'h00000000} /* (4, 20, 8) {real, imag} */,
  {32'h447ae08c, 32'h00000000} /* (4, 20, 7) {real, imag} */,
  {32'h44e3f8ae, 32'h00000000} /* (4, 20, 6) {real, imag} */,
  {32'h44f3beb0, 32'h00000000} /* (4, 20, 5) {real, imag} */,
  {32'h448bc3a9, 32'h00000000} /* (4, 20, 4) {real, imag} */,
  {32'h439bd1ad, 32'h00000000} /* (4, 20, 3) {real, imag} */,
  {32'h44a08c1c, 32'h00000000} /* (4, 20, 2) {real, imag} */,
  {32'h4474d41d, 32'h00000000} /* (4, 20, 1) {real, imag} */,
  {32'h43772bd8, 32'h00000000} /* (4, 20, 0) {real, imag} */,
  {32'h4497dec5, 32'h00000000} /* (4, 19, 31) {real, imag} */,
  {32'h45311185, 32'h00000000} /* (4, 19, 30) {real, imag} */,
  {32'h44f1e3eb, 32'h00000000} /* (4, 19, 29) {real, imag} */,
  {32'h452652e9, 32'h00000000} /* (4, 19, 28) {real, imag} */,
  {32'h44f438f0, 32'h00000000} /* (4, 19, 27) {real, imag} */,
  {32'h450644d1, 32'h00000000} /* (4, 19, 26) {real, imag} */,
  {32'h452096e6, 32'h00000000} /* (4, 19, 25) {real, imag} */,
  {32'h4523773d, 32'h00000000} /* (4, 19, 24) {real, imag} */,
  {32'h44f61fdc, 32'h00000000} /* (4, 19, 23) {real, imag} */,
  {32'h44dad5e9, 32'h00000000} /* (4, 19, 22) {real, imag} */,
  {32'h4448a6e3, 32'h00000000} /* (4, 19, 21) {real, imag} */,
  {32'hc3fea794, 32'h00000000} /* (4, 19, 20) {real, imag} */,
  {32'hc4a0fa57, 32'h00000000} /* (4, 19, 19) {real, imag} */,
  {32'hc47852fd, 32'h00000000} /* (4, 19, 18) {real, imag} */,
  {32'hc5182796, 32'h00000000} /* (4, 19, 17) {real, imag} */,
  {32'hc4a3b833, 32'h00000000} /* (4, 19, 16) {real, imag} */,
  {32'hc4b234f1, 32'h00000000} /* (4, 19, 15) {real, imag} */,
  {32'hc4922242, 32'h00000000} /* (4, 19, 14) {real, imag} */,
  {32'hc49074a7, 32'h00000000} /* (4, 19, 13) {real, imag} */,
  {32'hc498969e, 32'h00000000} /* (4, 19, 12) {real, imag} */,
  {32'hc436f97c, 32'h00000000} /* (4, 19, 11) {real, imag} */,
  {32'h444a493c, 32'h00000000} /* (4, 19, 10) {real, imag} */,
  {32'h44b7040d, 32'h00000000} /* (4, 19, 9) {real, imag} */,
  {32'h44ac4838, 32'h00000000} /* (4, 19, 8) {real, imag} */,
  {32'h450ea128, 32'h00000000} /* (4, 19, 7) {real, imag} */,
  {32'h44e1a83f, 32'h00000000} /* (4, 19, 6) {real, imag} */,
  {32'h4519245d, 32'h00000000} /* (4, 19, 5) {real, imag} */,
  {32'h450cc134, 32'h00000000} /* (4, 19, 4) {real, imag} */,
  {32'h44f445d5, 32'h00000000} /* (4, 19, 3) {real, imag} */,
  {32'h43d52cf6, 32'h00000000} /* (4, 19, 2) {real, imag} */,
  {32'h4464f246, 32'h00000000} /* (4, 19, 1) {real, imag} */,
  {32'h44b74171, 32'h00000000} /* (4, 19, 0) {real, imag} */,
  {32'h44be1306, 32'h00000000} /* (4, 18, 31) {real, imag} */,
  {32'h450ebe20, 32'h00000000} /* (4, 18, 30) {real, imag} */,
  {32'h45000a4c, 32'h00000000} /* (4, 18, 29) {real, imag} */,
  {32'h45088eda, 32'h00000000} /* (4, 18, 28) {real, imag} */,
  {32'h44ec1d3f, 32'h00000000} /* (4, 18, 27) {real, imag} */,
  {32'h44c26e86, 32'h00000000} /* (4, 18, 26) {real, imag} */,
  {32'h44fb00a4, 32'h00000000} /* (4, 18, 25) {real, imag} */,
  {32'h4510bf80, 32'h00000000} /* (4, 18, 24) {real, imag} */,
  {32'h450155ff, 32'h00000000} /* (4, 18, 23) {real, imag} */,
  {32'h44d284fb, 32'h00000000} /* (4, 18, 22) {real, imag} */,
  {32'h44c72db6, 32'h00000000} /* (4, 18, 21) {real, imag} */,
  {32'hc442f772, 32'h00000000} /* (4, 18, 20) {real, imag} */,
  {32'hc4aaee04, 32'h00000000} /* (4, 18, 19) {real, imag} */,
  {32'hc434ddfa, 32'h00000000} /* (4, 18, 18) {real, imag} */,
  {32'hc4ac91ba, 32'h00000000} /* (4, 18, 17) {real, imag} */,
  {32'hc4b3cb71, 32'h00000000} /* (4, 18, 16) {real, imag} */,
  {32'hc4e44cfa, 32'h00000000} /* (4, 18, 15) {real, imag} */,
  {32'hc4d67756, 32'h00000000} /* (4, 18, 14) {real, imag} */,
  {32'hc50a7b94, 32'h00000000} /* (4, 18, 13) {real, imag} */,
  {32'hc48e4d67, 32'h00000000} /* (4, 18, 12) {real, imag} */,
  {32'hc4ad3529, 32'h00000000} /* (4, 18, 11) {real, imag} */,
  {32'h439ca860, 32'h00000000} /* (4, 18, 10) {real, imag} */,
  {32'h44fd467c, 32'h00000000} /* (4, 18, 9) {real, imag} */,
  {32'h44ce07c4, 32'h00000000} /* (4, 18, 8) {real, imag} */,
  {32'h44f9531e, 32'h00000000} /* (4, 18, 7) {real, imag} */,
  {32'h453d7032, 32'h00000000} /* (4, 18, 6) {real, imag} */,
  {32'h452f31b5, 32'h00000000} /* (4, 18, 5) {real, imag} */,
  {32'h4530f1f8, 32'h00000000} /* (4, 18, 4) {real, imag} */,
  {32'h44bdcdae, 32'h00000000} /* (4, 18, 3) {real, imag} */,
  {32'h44a20f5f, 32'h00000000} /* (4, 18, 2) {real, imag} */,
  {32'h44cd9ab6, 32'h00000000} /* (4, 18, 1) {real, imag} */,
  {32'h44902bf9, 32'h00000000} /* (4, 18, 0) {real, imag} */,
  {32'h44c2d668, 32'h00000000} /* (4, 17, 31) {real, imag} */,
  {32'h450d52ee, 32'h00000000} /* (4, 17, 30) {real, imag} */,
  {32'h44e642d4, 32'h00000000} /* (4, 17, 29) {real, imag} */,
  {32'h44fc4ecb, 32'h00000000} /* (4, 17, 28) {real, imag} */,
  {32'h450e3218, 32'h00000000} /* (4, 17, 27) {real, imag} */,
  {32'h45180f91, 32'h00000000} /* (4, 17, 26) {real, imag} */,
  {32'h44e09a3f, 32'h00000000} /* (4, 17, 25) {real, imag} */,
  {32'h44ec8a3c, 32'h00000000} /* (4, 17, 24) {real, imag} */,
  {32'h450c4eca, 32'h00000000} /* (4, 17, 23) {real, imag} */,
  {32'h44d7e58e, 32'h00000000} /* (4, 17, 22) {real, imag} */,
  {32'h446651a2, 32'h00000000} /* (4, 17, 21) {real, imag} */,
  {32'hc45090ee, 32'h00000000} /* (4, 17, 20) {real, imag} */,
  {32'hc4d4567c, 32'h00000000} /* (4, 17, 19) {real, imag} */,
  {32'hc471c853, 32'h00000000} /* (4, 17, 18) {real, imag} */,
  {32'hc4c746bb, 32'h00000000} /* (4, 17, 17) {real, imag} */,
  {32'hc515989f, 32'h00000000} /* (4, 17, 16) {real, imag} */,
  {32'hc5118fd4, 32'h00000000} /* (4, 17, 15) {real, imag} */,
  {32'hc4d70ef6, 32'h00000000} /* (4, 17, 14) {real, imag} */,
  {32'hc4e6a58c, 32'h00000000} /* (4, 17, 13) {real, imag} */,
  {32'hc4dce115, 32'h00000000} /* (4, 17, 12) {real, imag} */,
  {32'hc4d6a6e3, 32'h00000000} /* (4, 17, 11) {real, imag} */,
  {32'h449d51a2, 32'h00000000} /* (4, 17, 10) {real, imag} */,
  {32'h44ba1f3b, 32'h00000000} /* (4, 17, 9) {real, imag} */,
  {32'h44c5cd90, 32'h00000000} /* (4, 17, 8) {real, imag} */,
  {32'h44f804a1, 32'h00000000} /* (4, 17, 7) {real, imag} */,
  {32'h450753c7, 32'h00000000} /* (4, 17, 6) {real, imag} */,
  {32'h4567d266, 32'h00000000} /* (4, 17, 5) {real, imag} */,
  {32'h45276b9e, 32'h00000000} /* (4, 17, 4) {real, imag} */,
  {32'h451bb102, 32'h00000000} /* (4, 17, 3) {real, imag} */,
  {32'h450a98ee, 32'h00000000} /* (4, 17, 2) {real, imag} */,
  {32'h44d51599, 32'h00000000} /* (4, 17, 1) {real, imag} */,
  {32'h443b92c5, 32'h00000000} /* (4, 17, 0) {real, imag} */,
  {32'h44a2aa10, 32'h00000000} /* (4, 16, 31) {real, imag} */,
  {32'h44cf11d4, 32'h00000000} /* (4, 16, 30) {real, imag} */,
  {32'h4516fb94, 32'h00000000} /* (4, 16, 29) {real, imag} */,
  {32'h44ae36e5, 32'h00000000} /* (4, 16, 28) {real, imag} */,
  {32'h45079693, 32'h00000000} /* (4, 16, 27) {real, imag} */,
  {32'h4526fe0e, 32'h00000000} /* (4, 16, 26) {real, imag} */,
  {32'h451c4639, 32'h00000000} /* (4, 16, 25) {real, imag} */,
  {32'h44d6b033, 32'h00000000} /* (4, 16, 24) {real, imag} */,
  {32'h4510a141, 32'h00000000} /* (4, 16, 23) {real, imag} */,
  {32'h44f8f1b4, 32'h00000000} /* (4, 16, 22) {real, imag} */,
  {32'h44adf964, 32'h00000000} /* (4, 16, 21) {real, imag} */,
  {32'hc406083a, 32'h00000000} /* (4, 16, 20) {real, imag} */,
  {32'hc5011dbe, 32'h00000000} /* (4, 16, 19) {real, imag} */,
  {32'hc4fb16ae, 32'h00000000} /* (4, 16, 18) {real, imag} */,
  {32'hc4e2e778, 32'h00000000} /* (4, 16, 17) {real, imag} */,
  {32'hc52630fc, 32'h00000000} /* (4, 16, 16) {real, imag} */,
  {32'hc52e2baa, 32'h00000000} /* (4, 16, 15) {real, imag} */,
  {32'hc4cd7614, 32'h00000000} /* (4, 16, 14) {real, imag} */,
  {32'hc4e6dbdc, 32'h00000000} /* (4, 16, 13) {real, imag} */,
  {32'hc519d232, 32'h00000000} /* (4, 16, 12) {real, imag} */,
  {32'hc4f36a42, 32'h00000000} /* (4, 16, 11) {real, imag} */,
  {32'h4253a400, 32'h00000000} /* (4, 16, 10) {real, imag} */,
  {32'h44955922, 32'h00000000} /* (4, 16, 9) {real, imag} */,
  {32'h4510c1f0, 32'h00000000} /* (4, 16, 8) {real, imag} */,
  {32'h451a939f, 32'h00000000} /* (4, 16, 7) {real, imag} */,
  {32'h44d54dcc, 32'h00000000} /* (4, 16, 6) {real, imag} */,
  {32'h450aebdc, 32'h00000000} /* (4, 16, 5) {real, imag} */,
  {32'h44f50d29, 32'h00000000} /* (4, 16, 4) {real, imag} */,
  {32'h44fdbe8a, 32'h00000000} /* (4, 16, 3) {real, imag} */,
  {32'h44fe3902, 32'h00000000} /* (4, 16, 2) {real, imag} */,
  {32'h44a72228, 32'h00000000} /* (4, 16, 1) {real, imag} */,
  {32'h44e33c4c, 32'h00000000} /* (4, 16, 0) {real, imag} */,
  {32'h4476bc33, 32'h00000000} /* (4, 15, 31) {real, imag} */,
  {32'h452661cd, 32'h00000000} /* (4, 15, 30) {real, imag} */,
  {32'h452ce830, 32'h00000000} /* (4, 15, 29) {real, imag} */,
  {32'h4529c86d, 32'h00000000} /* (4, 15, 28) {real, imag} */,
  {32'h451c541d, 32'h00000000} /* (4, 15, 27) {real, imag} */,
  {32'h450a0788, 32'h00000000} /* (4, 15, 26) {real, imag} */,
  {32'h451529f5, 32'h00000000} /* (4, 15, 25) {real, imag} */,
  {32'h4501807d, 32'h00000000} /* (4, 15, 24) {real, imag} */,
  {32'h454125b1, 32'h00000000} /* (4, 15, 23) {real, imag} */,
  {32'h4521b2b8, 32'h00000000} /* (4, 15, 22) {real, imag} */,
  {32'h44c77abd, 32'h00000000} /* (4, 15, 21) {real, imag} */,
  {32'hc4824392, 32'h00000000} /* (4, 15, 20) {real, imag} */,
  {32'hc4aa4a83, 32'h00000000} /* (4, 15, 19) {real, imag} */,
  {32'hc4e6e562, 32'h00000000} /* (4, 15, 18) {real, imag} */,
  {32'hc4ecf602, 32'h00000000} /* (4, 15, 17) {real, imag} */,
  {32'hc4dad015, 32'h00000000} /* (4, 15, 16) {real, imag} */,
  {32'hc518e256, 32'h00000000} /* (4, 15, 15) {real, imag} */,
  {32'hc50c703b, 32'h00000000} /* (4, 15, 14) {real, imag} */,
  {32'hc55a13c6, 32'h00000000} /* (4, 15, 13) {real, imag} */,
  {32'hc50aa5b3, 32'h00000000} /* (4, 15, 12) {real, imag} */,
  {32'hc4aae9d2, 32'h00000000} /* (4, 15, 11) {real, imag} */,
  {32'h4439d986, 32'h00000000} /* (4, 15, 10) {real, imag} */,
  {32'h44b6874a, 32'h00000000} /* (4, 15, 9) {real, imag} */,
  {32'h44f7679d, 32'h00000000} /* (4, 15, 8) {real, imag} */,
  {32'h44bf6d12, 32'h00000000} /* (4, 15, 7) {real, imag} */,
  {32'h44a6b7d4, 32'h00000000} /* (4, 15, 6) {real, imag} */,
  {32'h4454940a, 32'h00000000} /* (4, 15, 5) {real, imag} */,
  {32'h44a3d5da, 32'h00000000} /* (4, 15, 4) {real, imag} */,
  {32'h44a0bb21, 32'h00000000} /* (4, 15, 3) {real, imag} */,
  {32'h44a98696, 32'h00000000} /* (4, 15, 2) {real, imag} */,
  {32'h45069edb, 32'h00000000} /* (4, 15, 1) {real, imag} */,
  {32'h44eb1f3b, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'h4520bb48, 32'h00000000} /* (4, 14, 31) {real, imag} */,
  {32'h44fa8cdc, 32'h00000000} /* (4, 14, 30) {real, imag} */,
  {32'h4519e758, 32'h00000000} /* (4, 14, 29) {real, imag} */,
  {32'h45603404, 32'h00000000} /* (4, 14, 28) {real, imag} */,
  {32'h4516ff6e, 32'h00000000} /* (4, 14, 27) {real, imag} */,
  {32'h4504efca, 32'h00000000} /* (4, 14, 26) {real, imag} */,
  {32'h44f0a84d, 32'h00000000} /* (4, 14, 25) {real, imag} */,
  {32'h44c1ac7e, 32'h00000000} /* (4, 14, 24) {real, imag} */,
  {32'h44f30e0a, 32'h00000000} /* (4, 14, 23) {real, imag} */,
  {32'h45185896, 32'h00000000} /* (4, 14, 22) {real, imag} */,
  {32'h44883c3c, 32'h00000000} /* (4, 14, 21) {real, imag} */,
  {32'hc452438a, 32'h00000000} /* (4, 14, 20) {real, imag} */,
  {32'hc48a10fd, 32'h00000000} /* (4, 14, 19) {real, imag} */,
  {32'hc4cbbf0f, 32'h00000000} /* (4, 14, 18) {real, imag} */,
  {32'hc5220306, 32'h00000000} /* (4, 14, 17) {real, imag} */,
  {32'hc4efacd4, 32'h00000000} /* (4, 14, 16) {real, imag} */,
  {32'hc52e3570, 32'h00000000} /* (4, 14, 15) {real, imag} */,
  {32'hc501e6d0, 32'h00000000} /* (4, 14, 14) {real, imag} */,
  {32'hc4fd6bc9, 32'h00000000} /* (4, 14, 13) {real, imag} */,
  {32'hc4de9c11, 32'h00000000} /* (4, 14, 12) {real, imag} */,
  {32'hc436a73e, 32'h00000000} /* (4, 14, 11) {real, imag} */,
  {32'h440b53ee, 32'h00000000} /* (4, 14, 10) {real, imag} */,
  {32'h44c4df6f, 32'h00000000} /* (4, 14, 9) {real, imag} */,
  {32'h44dc9a42, 32'h00000000} /* (4, 14, 8) {real, imag} */,
  {32'h45232bbf, 32'h00000000} /* (4, 14, 7) {real, imag} */,
  {32'h44c0982b, 32'h00000000} /* (4, 14, 6) {real, imag} */,
  {32'h44afb8a8, 32'h00000000} /* (4, 14, 5) {real, imag} */,
  {32'h448e1712, 32'h00000000} /* (4, 14, 4) {real, imag} */,
  {32'h4447c396, 32'h00000000} /* (4, 14, 3) {real, imag} */,
  {32'h44222446, 32'h00000000} /* (4, 14, 2) {real, imag} */,
  {32'h452881bc, 32'h00000000} /* (4, 14, 1) {real, imag} */,
  {32'h44dd2f74, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'h44d14602, 32'h00000000} /* (4, 13, 31) {real, imag} */,
  {32'h44d820fb, 32'h00000000} /* (4, 13, 30) {real, imag} */,
  {32'h45158bfc, 32'h00000000} /* (4, 13, 29) {real, imag} */,
  {32'h4514aa18, 32'h00000000} /* (4, 13, 28) {real, imag} */,
  {32'h45459cbb, 32'h00000000} /* (4, 13, 27) {real, imag} */,
  {32'h45183e68, 32'h00000000} /* (4, 13, 26) {real, imag} */,
  {32'h44b9a094, 32'h00000000} /* (4, 13, 25) {real, imag} */,
  {32'h44ce578b, 32'h00000000} /* (4, 13, 24) {real, imag} */,
  {32'h44b0dfb1, 32'h00000000} /* (4, 13, 23) {real, imag} */,
  {32'h450d0861, 32'h00000000} /* (4, 13, 22) {real, imag} */,
  {32'h44f1df5a, 32'h00000000} /* (4, 13, 21) {real, imag} */,
  {32'hc4b45684, 32'h00000000} /* (4, 13, 20) {real, imag} */,
  {32'hc51da5c3, 32'h00000000} /* (4, 13, 19) {real, imag} */,
  {32'hc50970d2, 32'h00000000} /* (4, 13, 18) {real, imag} */,
  {32'hc52ee14d, 32'h00000000} /* (4, 13, 17) {real, imag} */,
  {32'hc4fd040c, 32'h00000000} /* (4, 13, 16) {real, imag} */,
  {32'hc4cd27c2, 32'h00000000} /* (4, 13, 15) {real, imag} */,
  {32'hc4eb985f, 32'h00000000} /* (4, 13, 14) {real, imag} */,
  {32'hc4fffa58, 32'h00000000} /* (4, 13, 13) {real, imag} */,
  {32'hc48ea8c7, 32'h00000000} /* (4, 13, 12) {real, imag} */,
  {32'hc4338cdc, 32'h00000000} /* (4, 13, 11) {real, imag} */,
  {32'h44236a1f, 32'h00000000} /* (4, 13, 10) {real, imag} */,
  {32'h44683ab8, 32'h00000000} /* (4, 13, 9) {real, imag} */,
  {32'h4481eee9, 32'h00000000} /* (4, 13, 8) {real, imag} */,
  {32'h44bb1773, 32'h00000000} /* (4, 13, 7) {real, imag} */,
  {32'h44acc766, 32'h00000000} /* (4, 13, 6) {real, imag} */,
  {32'h447ca9b7, 32'h00000000} /* (4, 13, 5) {real, imag} */,
  {32'h443e7db0, 32'h00000000} /* (4, 13, 4) {real, imag} */,
  {32'h449d388a, 32'h00000000} /* (4, 13, 3) {real, imag} */,
  {32'h4515c82c, 32'h00000000} /* (4, 13, 2) {real, imag} */,
  {32'h4517504d, 32'h00000000} /* (4, 13, 1) {real, imag} */,
  {32'h452c8778, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'h449a1de1, 32'h00000000} /* (4, 12, 31) {real, imag} */,
  {32'h44f29952, 32'h00000000} /* (4, 12, 30) {real, imag} */,
  {32'h451eb1e3, 32'h00000000} /* (4, 12, 29) {real, imag} */,
  {32'h4512a7fc, 32'h00000000} /* (4, 12, 28) {real, imag} */,
  {32'h450a9f84, 32'h00000000} /* (4, 12, 27) {real, imag} */,
  {32'h44ddfb9a, 32'h00000000} /* (4, 12, 26) {real, imag} */,
  {32'h44c16fa6, 32'h00000000} /* (4, 12, 25) {real, imag} */,
  {32'h451777d2, 32'h00000000} /* (4, 12, 24) {real, imag} */,
  {32'h44f8aa7e, 32'h00000000} /* (4, 12, 23) {real, imag} */,
  {32'h4524edca, 32'h00000000} /* (4, 12, 22) {real, imag} */,
  {32'h448ebe6a, 32'h00000000} /* (4, 12, 21) {real, imag} */,
  {32'hc4653ee5, 32'h00000000} /* (4, 12, 20) {real, imag} */,
  {32'hc5144918, 32'h00000000} /* (4, 12, 19) {real, imag} */,
  {32'hc4c764d1, 32'h00000000} /* (4, 12, 18) {real, imag} */,
  {32'hc5003d94, 32'h00000000} /* (4, 12, 17) {real, imag} */,
  {32'hc4cf05d9, 32'h00000000} /* (4, 12, 16) {real, imag} */,
  {32'hc4c5bd01, 32'h00000000} /* (4, 12, 15) {real, imag} */,
  {32'hc4dd881e, 32'h00000000} /* (4, 12, 14) {real, imag} */,
  {32'hc4bb3dcc, 32'h00000000} /* (4, 12, 13) {real, imag} */,
  {32'hc489868e, 32'h00000000} /* (4, 12, 12) {real, imag} */,
  {32'hc3525330, 32'h00000000} /* (4, 12, 11) {real, imag} */,
  {32'h449dd22e, 32'h00000000} /* (4, 12, 10) {real, imag} */,
  {32'h4494f21c, 32'h00000000} /* (4, 12, 9) {real, imag} */,
  {32'h442d6506, 32'h00000000} /* (4, 12, 8) {real, imag} */,
  {32'h44a0f542, 32'h00000000} /* (4, 12, 7) {real, imag} */,
  {32'h44944158, 32'h00000000} /* (4, 12, 6) {real, imag} */,
  {32'h4464e049, 32'h00000000} /* (4, 12, 5) {real, imag} */,
  {32'h44e21906, 32'h00000000} /* (4, 12, 4) {real, imag} */,
  {32'h449765f3, 32'h00000000} /* (4, 12, 3) {real, imag} */,
  {32'h4509c770, 32'h00000000} /* (4, 12, 2) {real, imag} */,
  {32'h45057c5c, 32'h00000000} /* (4, 12, 1) {real, imag} */,
  {32'h44fca23f, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'h449c5ce6, 32'h00000000} /* (4, 11, 31) {real, imag} */,
  {32'h44e6a684, 32'h00000000} /* (4, 11, 30) {real, imag} */,
  {32'h44c998a4, 32'h00000000} /* (4, 11, 29) {real, imag} */,
  {32'h4525dc2a, 32'h00000000} /* (4, 11, 28) {real, imag} */,
  {32'h44dfbad7, 32'h00000000} /* (4, 11, 27) {real, imag} */,
  {32'h44c8507a, 32'h00000000} /* (4, 11, 26) {real, imag} */,
  {32'h44a197a3, 32'h00000000} /* (4, 11, 25) {real, imag} */,
  {32'h447d160f, 32'h00000000} /* (4, 11, 24) {real, imag} */,
  {32'h450dc966, 32'h00000000} /* (4, 11, 23) {real, imag} */,
  {32'h450545bc, 32'h00000000} /* (4, 11, 22) {real, imag} */,
  {32'h447c72a1, 32'h00000000} /* (4, 11, 21) {real, imag} */,
  {32'hc38ab563, 32'h00000000} /* (4, 11, 20) {real, imag} */,
  {32'hc487ba25, 32'h00000000} /* (4, 11, 19) {real, imag} */,
  {32'hc4f224b3, 32'h00000000} /* (4, 11, 18) {real, imag} */,
  {32'hc4b6f84e, 32'h00000000} /* (4, 11, 17) {real, imag} */,
  {32'hc42f7fbd, 32'h00000000} /* (4, 11, 16) {real, imag} */,
  {32'hc4c639e8, 32'h00000000} /* (4, 11, 15) {real, imag} */,
  {32'hc4d5c18c, 32'h00000000} /* (4, 11, 14) {real, imag} */,
  {32'hc4b78666, 32'h00000000} /* (4, 11, 13) {real, imag} */,
  {32'hc4595fae, 32'h00000000} /* (4, 11, 12) {real, imag} */,
  {32'hc4185666, 32'h00000000} /* (4, 11, 11) {real, imag} */,
  {32'h44e9f6d6, 32'h00000000} /* (4, 11, 10) {real, imag} */,
  {32'h4479d38b, 32'h00000000} /* (4, 11, 9) {real, imag} */,
  {32'h439a5736, 32'h00000000} /* (4, 11, 8) {real, imag} */,
  {32'h445fd448, 32'h00000000} /* (4, 11, 7) {real, imag} */,
  {32'h448b64d0, 32'h00000000} /* (4, 11, 6) {real, imag} */,
  {32'h448ae840, 32'h00000000} /* (4, 11, 5) {real, imag} */,
  {32'h442b933c, 32'h00000000} /* (4, 11, 4) {real, imag} */,
  {32'h449ba3eb, 32'h00000000} /* (4, 11, 3) {real, imag} */,
  {32'h447fba96, 32'h00000000} /* (4, 11, 2) {real, imag} */,
  {32'h4501f47a, 32'h00000000} /* (4, 11, 1) {real, imag} */,
  {32'h44ccddfe, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'h4424bc3b, 32'h00000000} /* (4, 10, 31) {real, imag} */,
  {32'h44347bc1, 32'h00000000} /* (4, 10, 30) {real, imag} */,
  {32'h43762da4, 32'h00000000} /* (4, 10, 29) {real, imag} */,
  {32'hc2ea2c5c, 32'h00000000} /* (4, 10, 28) {real, imag} */,
  {32'hc3dcf08d, 32'h00000000} /* (4, 10, 27) {real, imag} */,
  {32'hc2fe4824, 32'h00000000} /* (4, 10, 26) {real, imag} */,
  {32'hc3c06c72, 32'h00000000} /* (4, 10, 25) {real, imag} */,
  {32'hc1d3e800, 32'h00000000} /* (4, 10, 24) {real, imag} */,
  {32'hc419f7b8, 32'h00000000} /* (4, 10, 23) {real, imag} */,
  {32'h4396bfbb, 32'h00000000} /* (4, 10, 22) {real, imag} */,
  {32'hc331738a, 32'h00000000} /* (4, 10, 21) {real, imag} */,
  {32'h4446fb66, 32'h00000000} /* (4, 10, 20) {real, imag} */,
  {32'h44a0ba6b, 32'h00000000} /* (4, 10, 19) {real, imag} */,
  {32'hc45a4dae, 32'h00000000} /* (4, 10, 18) {real, imag} */,
  {32'h4321c04a, 32'h00000000} /* (4, 10, 17) {real, imag} */,
  {32'h442d07b6, 32'h00000000} /* (4, 10, 16) {real, imag} */,
  {32'h440e01a9, 32'h00000000} /* (4, 10, 15) {real, imag} */,
  {32'hc330ce78, 32'h00000000} /* (4, 10, 14) {real, imag} */,
  {32'hc3611cae, 32'h00000000} /* (4, 10, 13) {real, imag} */,
  {32'h442b5b22, 32'h00000000} /* (4, 10, 12) {real, imag} */,
  {32'h44a2c1bd, 32'h00000000} /* (4, 10, 11) {real, imag} */,
  {32'hc3fa6f67, 32'h00000000} /* (4, 10, 10) {real, imag} */,
  {32'hc45b55d1, 32'h00000000} /* (4, 10, 9) {real, imag} */,
  {32'hc485db1c, 32'h00000000} /* (4, 10, 8) {real, imag} */,
  {32'hc4aab16a, 32'h00000000} /* (4, 10, 7) {real, imag} */,
  {32'hc4019f0e, 32'h00000000} /* (4, 10, 6) {real, imag} */,
  {32'hc36a01a2, 32'h00000000} /* (4, 10, 5) {real, imag} */,
  {32'hc468a21c, 32'h00000000} /* (4, 10, 4) {real, imag} */,
  {32'hc45d840e, 32'h00000000} /* (4, 10, 3) {real, imag} */,
  {32'hc36d2690, 32'h00000000} /* (4, 10, 2) {real, imag} */,
  {32'h43cdd21b, 32'h00000000} /* (4, 10, 1) {real, imag} */,
  {32'h43467d6e, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'h42ef0c48, 32'h00000000} /* (4, 9, 31) {real, imag} */,
  {32'hc4012152, 32'h00000000} /* (4, 9, 30) {real, imag} */,
  {32'hc490834a, 32'h00000000} /* (4, 9, 29) {real, imag} */,
  {32'hc49e5896, 32'h00000000} /* (4, 9, 28) {real, imag} */,
  {32'hc46c6ee2, 32'h00000000} /* (4, 9, 27) {real, imag} */,
  {32'hc47b22fe, 32'h00000000} /* (4, 9, 26) {real, imag} */,
  {32'hc418ab88, 32'h00000000} /* (4, 9, 25) {real, imag} */,
  {32'hc45132a8, 32'h00000000} /* (4, 9, 24) {real, imag} */,
  {32'hc49d833b, 32'h00000000} /* (4, 9, 23) {real, imag} */,
  {32'hc30f09c2, 32'h00000000} /* (4, 9, 22) {real, imag} */,
  {32'hc3a76d1c, 32'h00000000} /* (4, 9, 21) {real, imag} */,
  {32'h450d3438, 32'h00000000} /* (4, 9, 20) {real, imag} */,
  {32'h44d6fd50, 32'h00000000} /* (4, 9, 19) {real, imag} */,
  {32'h44fb2862, 32'h00000000} /* (4, 9, 18) {real, imag} */,
  {32'h44c21133, 32'h00000000} /* (4, 9, 17) {real, imag} */,
  {32'h44d5b228, 32'h00000000} /* (4, 9, 16) {real, imag} */,
  {32'h44ad26f6, 32'h00000000} /* (4, 9, 15) {real, imag} */,
  {32'h4485752f, 32'h00000000} /* (4, 9, 14) {real, imag} */,
  {32'h4467ab65, 32'h00000000} /* (4, 9, 13) {real, imag} */,
  {32'h44b9c256, 32'h00000000} /* (4, 9, 12) {real, imag} */,
  {32'h44a5951d, 32'h00000000} /* (4, 9, 11) {real, imag} */,
  {32'hc3185dfe, 32'h00000000} /* (4, 9, 10) {real, imag} */,
  {32'hc4eee732, 32'h00000000} /* (4, 9, 9) {real, imag} */,
  {32'hc4ceb25e, 32'h00000000} /* (4, 9, 8) {real, imag} */,
  {32'hc4b5d289, 32'h00000000} /* (4, 9, 7) {real, imag} */,
  {32'hc4470c7e, 32'h00000000} /* (4, 9, 6) {real, imag} */,
  {32'hc48a462d, 32'h00000000} /* (4, 9, 5) {real, imag} */,
  {32'hc48e1492, 32'h00000000} /* (4, 9, 4) {real, imag} */,
  {32'hc4734b40, 32'h00000000} /* (4, 9, 3) {real, imag} */,
  {32'hc4e208b0, 32'h00000000} /* (4, 9, 2) {real, imag} */,
  {32'hc39b1ae4, 32'h00000000} /* (4, 9, 1) {real, imag} */,
  {32'hc2397b40, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'h430520f0, 32'h00000000} /* (4, 8, 31) {real, imag} */,
  {32'hc3fed945, 32'h00000000} /* (4, 8, 30) {real, imag} */,
  {32'hc49feb0f, 32'h00000000} /* (4, 8, 29) {real, imag} */,
  {32'hc4cd382e, 32'h00000000} /* (4, 8, 28) {real, imag} */,
  {32'hc4b3d9b4, 32'h00000000} /* (4, 8, 27) {real, imag} */,
  {32'hc4dc9f0e, 32'h00000000} /* (4, 8, 26) {real, imag} */,
  {32'hc4b1d911, 32'h00000000} /* (4, 8, 25) {real, imag} */,
  {32'hc4225589, 32'h00000000} /* (4, 8, 24) {real, imag} */,
  {32'hc34f65f7, 32'h00000000} /* (4, 8, 23) {real, imag} */,
  {32'hc354870c, 32'h00000000} /* (4, 8, 22) {real, imag} */,
  {32'h444fd4b8, 32'h00000000} /* (4, 8, 21) {real, imag} */,
  {32'h44fa25a2, 32'h00000000} /* (4, 8, 20) {real, imag} */,
  {32'h4514de55, 32'h00000000} /* (4, 8, 19) {real, imag} */,
  {32'h4532d74f, 32'h00000000} /* (4, 8, 18) {real, imag} */,
  {32'h450c5cb2, 32'h00000000} /* (4, 8, 17) {real, imag} */,
  {32'h45120d1a, 32'h00000000} /* (4, 8, 16) {real, imag} */,
  {32'h45273363, 32'h00000000} /* (4, 8, 15) {real, imag} */,
  {32'h44319c5c, 32'h00000000} /* (4, 8, 14) {real, imag} */,
  {32'h4479cf63, 32'h00000000} /* (4, 8, 13) {real, imag} */,
  {32'h4505166a, 32'h00000000} /* (4, 8, 12) {real, imag} */,
  {32'h440c6412, 32'h00000000} /* (4, 8, 11) {real, imag} */,
  {32'hc3b4ca66, 32'h00000000} /* (4, 8, 10) {real, imag} */,
  {32'hc49807f5, 32'h00000000} /* (4, 8, 9) {real, imag} */,
  {32'hc4f929fa, 32'h00000000} /* (4, 8, 8) {real, imag} */,
  {32'hc42462cf, 32'h00000000} /* (4, 8, 7) {real, imag} */,
  {32'hc4abae1e, 32'h00000000} /* (4, 8, 6) {real, imag} */,
  {32'hc4d054d6, 32'h00000000} /* (4, 8, 5) {real, imag} */,
  {32'hc4eb6242, 32'h00000000} /* (4, 8, 4) {real, imag} */,
  {32'hc497b406, 32'h00000000} /* (4, 8, 3) {real, imag} */,
  {32'hc417a594, 32'h00000000} /* (4, 8, 2) {real, imag} */,
  {32'hc44cfa70, 32'h00000000} /* (4, 8, 1) {real, imag} */,
  {32'hc22e40c0, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'h43b34e90, 32'h00000000} /* (4, 7, 31) {real, imag} */,
  {32'hc3843230, 32'h00000000} /* (4, 7, 30) {real, imag} */,
  {32'hc3e0bbcd, 32'h00000000} /* (4, 7, 29) {real, imag} */,
  {32'hc490b9e7, 32'h00000000} /* (4, 7, 28) {real, imag} */,
  {32'hc4e2d4ea, 32'h00000000} /* (4, 7, 27) {real, imag} */,
  {32'hc5288204, 32'h00000000} /* (4, 7, 26) {real, imag} */,
  {32'hc4d01447, 32'h00000000} /* (4, 7, 25) {real, imag} */,
  {32'hc4b492db, 32'h00000000} /* (4, 7, 24) {real, imag} */,
  {32'hc28b28be, 32'h00000000} /* (4, 7, 23) {real, imag} */,
  {32'h435eeb82, 32'h00000000} /* (4, 7, 22) {real, imag} */,
  {32'h448f6469, 32'h00000000} /* (4, 7, 21) {real, imag} */,
  {32'h44eca48f, 32'h00000000} /* (4, 7, 20) {real, imag} */,
  {32'h4510c8f0, 32'h00000000} /* (4, 7, 19) {real, imag} */,
  {32'h45280fd0, 32'h00000000} /* (4, 7, 18) {real, imag} */,
  {32'h4547da82, 32'h00000000} /* (4, 7, 17) {real, imag} */,
  {32'h451ac866, 32'h00000000} /* (4, 7, 16) {real, imag} */,
  {32'h45395a40, 32'h00000000} /* (4, 7, 15) {real, imag} */,
  {32'h4528bf36, 32'h00000000} /* (4, 7, 14) {real, imag} */,
  {32'h44b712ad, 32'h00000000} /* (4, 7, 13) {real, imag} */,
  {32'h44e03ba5, 32'h00000000} /* (4, 7, 12) {real, imag} */,
  {32'h44ea7346, 32'h00000000} /* (4, 7, 11) {real, imag} */,
  {32'hc38800a4, 32'h00000000} /* (4, 7, 10) {real, imag} */,
  {32'h43ace10c, 32'h00000000} /* (4, 7, 9) {real, imag} */,
  {32'hc436c282, 32'h00000000} /* (4, 7, 8) {real, imag} */,
  {32'hc4064e12, 32'h00000000} /* (4, 7, 7) {real, imag} */,
  {32'hc497d904, 32'h00000000} /* (4, 7, 6) {real, imag} */,
  {32'hc4bd1553, 32'h00000000} /* (4, 7, 5) {real, imag} */,
  {32'hc5010f67, 32'h00000000} /* (4, 7, 4) {real, imag} */,
  {32'hc4327393, 32'h00000000} /* (4, 7, 3) {real, imag} */,
  {32'hc3a6c0c4, 32'h00000000} /* (4, 7, 2) {real, imag} */,
  {32'h43dea794, 32'h00000000} /* (4, 7, 1) {real, imag} */,
  {32'h43b4a010, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'h43a81b74, 32'h00000000} /* (4, 6, 31) {real, imag} */,
  {32'h43de1996, 32'h00000000} /* (4, 6, 30) {real, imag} */,
  {32'hc50aa6dc, 32'h00000000} /* (4, 6, 29) {real, imag} */,
  {32'hc49c06ba, 32'h00000000} /* (4, 6, 28) {real, imag} */,
  {32'hc44835a3, 32'h00000000} /* (4, 6, 27) {real, imag} */,
  {32'hc4c80aa6, 32'h00000000} /* (4, 6, 26) {real, imag} */,
  {32'hc4a16e13, 32'h00000000} /* (4, 6, 25) {real, imag} */,
  {32'hc4776696, 32'h00000000} /* (4, 6, 24) {real, imag} */,
  {32'h440a67e8, 32'h00000000} /* (4, 6, 23) {real, imag} */,
  {32'h4430683b, 32'h00000000} /* (4, 6, 22) {real, imag} */,
  {32'h4429027b, 32'h00000000} /* (4, 6, 21) {real, imag} */,
  {32'h443e4c70, 32'h00000000} /* (4, 6, 20) {real, imag} */,
  {32'h44a4f4b4, 32'h00000000} /* (4, 6, 19) {real, imag} */,
  {32'h44f3b599, 32'h00000000} /* (4, 6, 18) {real, imag} */,
  {32'h4529f25a, 32'h00000000} /* (4, 6, 17) {real, imag} */,
  {32'h4506acc7, 32'h00000000} /* (4, 6, 16) {real, imag} */,
  {32'h44e2e2dd, 32'h00000000} /* (4, 6, 15) {real, imag} */,
  {32'h450fd463, 32'h00000000} /* (4, 6, 14) {real, imag} */,
  {32'h45107606, 32'h00000000} /* (4, 6, 13) {real, imag} */,
  {32'h44dca19a, 32'h00000000} /* (4, 6, 12) {real, imag} */,
  {32'h447fd245, 32'h00000000} /* (4, 6, 11) {real, imag} */,
  {32'h44420280, 32'h00000000} /* (4, 6, 10) {real, imag} */,
  {32'h417cf000, 32'h00000000} /* (4, 6, 9) {real, imag} */,
  {32'hc3d088f4, 32'h00000000} /* (4, 6, 8) {real, imag} */,
  {32'hc3f5cf18, 32'h00000000} /* (4, 6, 7) {real, imag} */,
  {32'hc4b41f60, 32'h00000000} /* (4, 6, 6) {real, imag} */,
  {32'hc340059c, 32'h00000000} /* (4, 6, 5) {real, imag} */,
  {32'hc45c8374, 32'h00000000} /* (4, 6, 4) {real, imag} */,
  {32'hc42d8246, 32'h00000000} /* (4, 6, 3) {real, imag} */,
  {32'hc38d95dc, 32'h00000000} /* (4, 6, 2) {real, imag} */,
  {32'h431ac2c8, 32'h00000000} /* (4, 6, 1) {real, imag} */,
  {32'h43af4998, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'h443514ac, 32'h00000000} /* (4, 5, 31) {real, imag} */,
  {32'h42dbc040, 32'h00000000} /* (4, 5, 30) {real, imag} */,
  {32'hc4c54d09, 32'h00000000} /* (4, 5, 29) {real, imag} */,
  {32'hc458f232, 32'h00000000} /* (4, 5, 28) {real, imag} */,
  {32'hc50a39f9, 32'h00000000} /* (4, 5, 27) {real, imag} */,
  {32'hc5245978, 32'h00000000} /* (4, 5, 26) {real, imag} */,
  {32'hc514ce91, 32'h00000000} /* (4, 5, 25) {real, imag} */,
  {32'hc4be992c, 32'h00000000} /* (4, 5, 24) {real, imag} */,
  {32'hc42d7473, 32'h00000000} /* (4, 5, 23) {real, imag} */,
  {32'h42007a20, 32'h00000000} /* (4, 5, 22) {real, imag} */,
  {32'hc34023e0, 32'h00000000} /* (4, 5, 21) {real, imag} */,
  {32'hc3fd5b2a, 32'h00000000} /* (4, 5, 20) {real, imag} */,
  {32'h42c0509e, 32'h00000000} /* (4, 5, 19) {real, imag} */,
  {32'h443f8ef4, 32'h00000000} /* (4, 5, 18) {real, imag} */,
  {32'hc351bf61, 32'h00000000} /* (4, 5, 17) {real, imag} */,
  {32'h43c30200, 32'h00000000} /* (4, 5, 16) {real, imag} */,
  {32'h4455cfee, 32'h00000000} /* (4, 5, 15) {real, imag} */,
  {32'h44fa47c6, 32'h00000000} /* (4, 5, 14) {real, imag} */,
  {32'h44e09e73, 32'h00000000} /* (4, 5, 13) {real, imag} */,
  {32'h452cbb58, 32'h00000000} /* (4, 5, 12) {real, imag} */,
  {32'h44c094c2, 32'h00000000} /* (4, 5, 11) {real, imag} */,
  {32'h44810489, 32'h00000000} /* (4, 5, 10) {real, imag} */,
  {32'h44b8a382, 32'h00000000} /* (4, 5, 9) {real, imag} */,
  {32'h448302f0, 32'h00000000} /* (4, 5, 8) {real, imag} */,
  {32'h450e3f80, 32'h00000000} /* (4, 5, 7) {real, imag} */,
  {32'h44a5aef1, 32'h00000000} /* (4, 5, 6) {real, imag} */,
  {32'h43bec8d0, 32'h00000000} /* (4, 5, 5) {real, imag} */,
  {32'h4195e180, 32'h00000000} /* (4, 5, 4) {real, imag} */,
  {32'hc39e2664, 32'h00000000} /* (4, 5, 3) {real, imag} */,
  {32'h436f272a, 32'h00000000} /* (4, 5, 2) {real, imag} */,
  {32'hc1e1f148, 32'h00000000} /* (4, 5, 1) {real, imag} */,
  {32'h43e9b4cc, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'h44662ca4, 32'h00000000} /* (4, 4, 31) {real, imag} */,
  {32'h42f89c30, 32'h00000000} /* (4, 4, 30) {real, imag} */,
  {32'hc4b3ea0b, 32'h00000000} /* (4, 4, 29) {real, imag} */,
  {32'hc51f4c12, 32'h00000000} /* (4, 4, 28) {real, imag} */,
  {32'hc49a15ff, 32'h00000000} /* (4, 4, 27) {real, imag} */,
  {32'hc42ca639, 32'h00000000} /* (4, 4, 26) {real, imag} */,
  {32'hc493e676, 32'h00000000} /* (4, 4, 25) {real, imag} */,
  {32'hc50b5030, 32'h00000000} /* (4, 4, 24) {real, imag} */,
  {32'hc4ca9bf3, 32'h00000000} /* (4, 4, 23) {real, imag} */,
  {32'h434cbc60, 32'h00000000} /* (4, 4, 22) {real, imag} */,
  {32'hc44b0639, 32'h00000000} /* (4, 4, 21) {real, imag} */,
  {32'hc3fef51c, 32'h00000000} /* (4, 4, 20) {real, imag} */,
  {32'hc4583b89, 32'h00000000} /* (4, 4, 19) {real, imag} */,
  {32'hc45668ce, 32'h00000000} /* (4, 4, 18) {real, imag} */,
  {32'hc43b73ca, 32'h00000000} /* (4, 4, 17) {real, imag} */,
  {32'hc42048ad, 32'h00000000} /* (4, 4, 16) {real, imag} */,
  {32'h4497d7ee, 32'h00000000} /* (4, 4, 15) {real, imag} */,
  {32'h45004868, 32'h00000000} /* (4, 4, 14) {real, imag} */,
  {32'h452cfe0e, 32'h00000000} /* (4, 4, 13) {real, imag} */,
  {32'h45079eaa, 32'h00000000} /* (4, 4, 12) {real, imag} */,
  {32'h4517da5c, 32'h00000000} /* (4, 4, 11) {real, imag} */,
  {32'h44e7b098, 32'h00000000} /* (4, 4, 10) {real, imag} */,
  {32'h44e26fee, 32'h00000000} /* (4, 4, 9) {real, imag} */,
  {32'h452f05d4, 32'h00000000} /* (4, 4, 8) {real, imag} */,
  {32'h45068ac3, 32'h00000000} /* (4, 4, 7) {real, imag} */,
  {32'h45221b7f, 32'h00000000} /* (4, 4, 6) {real, imag} */,
  {32'h44a7af90, 32'h00000000} /* (4, 4, 5) {real, imag} */,
  {32'hc41a5862, 32'h00000000} /* (4, 4, 4) {real, imag} */,
  {32'hc42f77f7, 32'h00000000} /* (4, 4, 3) {real, imag} */,
  {32'hc3dacabf, 32'h00000000} /* (4, 4, 2) {real, imag} */,
  {32'hc3bd4813, 32'h00000000} /* (4, 4, 1) {real, imag} */,
  {32'h42db2e08, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'h43dc5771, 32'h00000000} /* (4, 3, 31) {real, imag} */,
  {32'hc235b3a0, 32'h00000000} /* (4, 3, 30) {real, imag} */,
  {32'hc4714384, 32'h00000000} /* (4, 3, 29) {real, imag} */,
  {32'hc4c95d0d, 32'h00000000} /* (4, 3, 28) {real, imag} */,
  {32'hc3034230, 32'h00000000} /* (4, 3, 27) {real, imag} */,
  {32'h43384608, 32'h00000000} /* (4, 3, 26) {real, imag} */,
  {32'hc398fff8, 32'h00000000} /* (4, 3, 25) {real, imag} */,
  {32'hc433a1c8, 32'h00000000} /* (4, 3, 24) {real, imag} */,
  {32'hc3fda854, 32'h00000000} /* (4, 3, 23) {real, imag} */,
  {32'hc42f6320, 32'h00000000} /* (4, 3, 22) {real, imag} */,
  {32'hc2c767a0, 32'h00000000} /* (4, 3, 21) {real, imag} */,
  {32'hc3f1cf11, 32'h00000000} /* (4, 3, 20) {real, imag} */,
  {32'hc4ac589c, 32'h00000000} /* (4, 3, 19) {real, imag} */,
  {32'hc4eb7987, 32'h00000000} /* (4, 3, 18) {real, imag} */,
  {32'hc4c71e8e, 32'h00000000} /* (4, 3, 17) {real, imag} */,
  {32'hc46a4058, 32'h00000000} /* (4, 3, 16) {real, imag} */,
  {32'h446a9054, 32'h00000000} /* (4, 3, 15) {real, imag} */,
  {32'h4526e83e, 32'h00000000} /* (4, 3, 14) {real, imag} */,
  {32'h45476af7, 32'h00000000} /* (4, 3, 13) {real, imag} */,
  {32'h44ea1b53, 32'h00000000} /* (4, 3, 12) {real, imag} */,
  {32'h45090533, 32'h00000000} /* (4, 3, 11) {real, imag} */,
  {32'h4535f4f6, 32'h00000000} /* (4, 3, 10) {real, imag} */,
  {32'h45146425, 32'h00000000} /* (4, 3, 9) {real, imag} */,
  {32'h4510cb59, 32'h00000000} /* (4, 3, 8) {real, imag} */,
  {32'h4524471c, 32'h00000000} /* (4, 3, 7) {real, imag} */,
  {32'h4540c5ff, 32'h00000000} /* (4, 3, 6) {real, imag} */,
  {32'h4506d87f, 32'h00000000} /* (4, 3, 5) {real, imag} */,
  {32'h435a089a, 32'h00000000} /* (4, 3, 4) {real, imag} */,
  {32'hc4a25320, 32'h00000000} /* (4, 3, 3) {real, imag} */,
  {32'hc407d3d2, 32'h00000000} /* (4, 3, 2) {real, imag} */,
  {32'hc26abe30, 32'h00000000} /* (4, 3, 1) {real, imag} */,
  {32'h4450f476, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'h4426ae70, 32'h00000000} /* (4, 2, 31) {real, imag} */,
  {32'h43075d34, 32'h00000000} /* (4, 2, 30) {real, imag} */,
  {32'h43a7f870, 32'h00000000} /* (4, 2, 29) {real, imag} */,
  {32'hc44258c8, 32'h00000000} /* (4, 2, 28) {real, imag} */,
  {32'hc3de6b9e, 32'h00000000} /* (4, 2, 27) {real, imag} */,
  {32'hc4826592, 32'h00000000} /* (4, 2, 26) {real, imag} */,
  {32'h42109800, 32'h00000000} /* (4, 2, 25) {real, imag} */,
  {32'h443a3f8c, 32'h00000000} /* (4, 2, 24) {real, imag} */,
  {32'h428727a0, 32'h00000000} /* (4, 2, 23) {real, imag} */,
  {32'h4399e178, 32'h00000000} /* (4, 2, 22) {real, imag} */,
  {32'hc42db8f2, 32'h00000000} /* (4, 2, 21) {real, imag} */,
  {32'hc4dd2e2c, 32'h00000000} /* (4, 2, 20) {real, imag} */,
  {32'hc4d2444f, 32'h00000000} /* (4, 2, 19) {real, imag} */,
  {32'hc4ac3830, 32'h00000000} /* (4, 2, 18) {real, imag} */,
  {32'hc46c2dcd, 32'h00000000} /* (4, 2, 17) {real, imag} */,
  {32'hc3b21d66, 32'h00000000} /* (4, 2, 16) {real, imag} */,
  {32'h4500c8f5, 32'h00000000} /* (4, 2, 15) {real, imag} */,
  {32'h44e54532, 32'h00000000} /* (4, 2, 14) {real, imag} */,
  {32'h44d68f8a, 32'h00000000} /* (4, 2, 13) {real, imag} */,
  {32'h456e23f8, 32'h00000000} /* (4, 2, 12) {real, imag} */,
  {32'h450ce166, 32'h00000000} /* (4, 2, 11) {real, imag} */,
  {32'h45143d2f, 32'h00000000} /* (4, 2, 10) {real, imag} */,
  {32'h451e22ed, 32'h00000000} /* (4, 2, 9) {real, imag} */,
  {32'h454180f5, 32'h00000000} /* (4, 2, 8) {real, imag} */,
  {32'h4531f96e, 32'h00000000} /* (4, 2, 7) {real, imag} */,
  {32'h45234a1b, 32'h00000000} /* (4, 2, 6) {real, imag} */,
  {32'h44dc5fd9, 32'h00000000} /* (4, 2, 5) {real, imag} */,
  {32'hc0c07f80, 32'h00000000} /* (4, 2, 4) {real, imag} */,
  {32'hc46c038a, 32'h00000000} /* (4, 2, 3) {real, imag} */,
  {32'hc3935bc6, 32'h00000000} /* (4, 2, 2) {real, imag} */,
  {32'hc3810ed6, 32'h00000000} /* (4, 2, 1) {real, imag} */,
  {32'h444413c1, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'h44adc2ee, 32'h00000000} /* (4, 1, 31) {real, imag} */,
  {32'h4451f8fa, 32'h00000000} /* (4, 1, 30) {real, imag} */,
  {32'hc1bac3c0, 32'h00000000} /* (4, 1, 29) {real, imag} */,
  {32'h433cfae8, 32'h00000000} /* (4, 1, 28) {real, imag} */,
  {32'hc35644e8, 32'h00000000} /* (4, 1, 27) {real, imag} */,
  {32'h43c0aad8, 32'h00000000} /* (4, 1, 26) {real, imag} */,
  {32'h4303bca8, 32'h00000000} /* (4, 1, 25) {real, imag} */,
  {32'h4318daa8, 32'h00000000} /* (4, 1, 24) {real, imag} */,
  {32'hc42e4798, 32'h00000000} /* (4, 1, 23) {real, imag} */,
  {32'hc1b22400, 32'h00000000} /* (4, 1, 22) {real, imag} */,
  {32'hc456c458, 32'h00000000} /* (4, 1, 21) {real, imag} */,
  {32'hc4452c9b, 32'h00000000} /* (4, 1, 20) {real, imag} */,
  {32'hc42d92e9, 32'h00000000} /* (4, 1, 19) {real, imag} */,
  {32'hc4a129ca, 32'h00000000} /* (4, 1, 18) {real, imag} */,
  {32'hc426222f, 32'h00000000} /* (4, 1, 17) {real, imag} */,
  {32'h42cc7168, 32'h00000000} /* (4, 1, 16) {real, imag} */,
  {32'h44a9d2a0, 32'h00000000} /* (4, 1, 15) {real, imag} */,
  {32'h45122c02, 32'h00000000} /* (4, 1, 14) {real, imag} */,
  {32'h454d3710, 32'h00000000} /* (4, 1, 13) {real, imag} */,
  {32'h450d5cba, 32'h00000000} /* (4, 1, 12) {real, imag} */,
  {32'h44e30a9f, 32'h00000000} /* (4, 1, 11) {real, imag} */,
  {32'h453441e1, 32'h00000000} /* (4, 1, 10) {real, imag} */,
  {32'h454c02e6, 32'h00000000} /* (4, 1, 9) {real, imag} */,
  {32'h451315c0, 32'h00000000} /* (4, 1, 8) {real, imag} */,
  {32'h45422953, 32'h00000000} /* (4, 1, 7) {real, imag} */,
  {32'h4540b233, 32'h00000000} /* (4, 1, 6) {real, imag} */,
  {32'h43c37178, 32'h00000000} /* (4, 1, 5) {real, imag} */,
  {32'hc4782767, 32'h00000000} /* (4, 1, 4) {real, imag} */,
  {32'hc3b5e076, 32'h00000000} /* (4, 1, 3) {real, imag} */,
  {32'h441eb08f, 32'h00000000} /* (4, 1, 2) {real, imag} */,
  {32'h442c7c13, 32'h00000000} /* (4, 1, 1) {real, imag} */,
  {32'h44870448, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'h44ddc9ab, 32'h00000000} /* (4, 0, 31) {real, imag} */,
  {32'h44ca0270, 32'h00000000} /* (4, 0, 30) {real, imag} */,
  {32'h437e1e88, 32'h00000000} /* (4, 0, 29) {real, imag} */,
  {32'h4416dfc4, 32'h00000000} /* (4, 0, 28) {real, imag} */,
  {32'h447ab4e7, 32'h00000000} /* (4, 0, 27) {real, imag} */,
  {32'h440622cf, 32'h00000000} /* (4, 0, 26) {real, imag} */,
  {32'h4387ce14, 32'h00000000} /* (4, 0, 25) {real, imag} */,
  {32'h43cbd27a, 32'h00000000} /* (4, 0, 24) {real, imag} */,
  {32'hc42aa80a, 32'h00000000} /* (4, 0, 23) {real, imag} */,
  {32'hc2513200, 32'h00000000} /* (4, 0, 22) {real, imag} */,
  {32'h43ab6c8a, 32'h00000000} /* (4, 0, 21) {real, imag} */,
  {32'h40ba9be0, 32'h00000000} /* (4, 0, 20) {real, imag} */,
  {32'h42a7cc38, 32'h00000000} /* (4, 0, 19) {real, imag} */,
  {32'h438296ce, 32'h00000000} /* (4, 0, 18) {real, imag} */,
  {32'hc1ec04d0, 32'h00000000} /* (4, 0, 17) {real, imag} */,
  {32'h446099ad, 32'h00000000} /* (4, 0, 16) {real, imag} */,
  {32'h44ae0d57, 32'h00000000} /* (4, 0, 15) {real, imag} */,
  {32'h450a01b8, 32'h00000000} /* (4, 0, 14) {real, imag} */,
  {32'h453f6c48, 32'h00000000} /* (4, 0, 13) {real, imag} */,
  {32'h44f037fc, 32'h00000000} /* (4, 0, 12) {real, imag} */,
  {32'h44d1b470, 32'h00000000} /* (4, 0, 11) {real, imag} */,
  {32'h44d1f600, 32'h00000000} /* (4, 0, 10) {real, imag} */,
  {32'h44e88c6d, 32'h00000000} /* (4, 0, 9) {real, imag} */,
  {32'h44b2d104, 32'h00000000} /* (4, 0, 8) {real, imag} */,
  {32'h4508969a, 32'h00000000} /* (4, 0, 7) {real, imag} */,
  {32'h450eae48, 32'h00000000} /* (4, 0, 6) {real, imag} */,
  {32'h43ba0632, 32'h00000000} /* (4, 0, 5) {real, imag} */,
  {32'hc3a96198, 32'h00000000} /* (4, 0, 4) {real, imag} */,
  {32'h426cebb0, 32'h00000000} /* (4, 0, 3) {real, imag} */,
  {32'h44319fc8, 32'h00000000} /* (4, 0, 2) {real, imag} */,
  {32'h4443b734, 32'h00000000} /* (4, 0, 1) {real, imag} */,
  {32'h44807796, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hc2395f80, 32'h00000000} /* (3, 31, 31) {real, imag} */,
  {32'hc3b1a968, 32'h00000000} /* (3, 31, 30) {real, imag} */,
  {32'hc490a89e, 32'h00000000} /* (3, 31, 29) {real, imag} */,
  {32'hc4d039fc, 32'h00000000} /* (3, 31, 28) {real, imag} */,
  {32'hc50dac03, 32'h00000000} /* (3, 31, 27) {real, imag} */,
  {32'hc4cbe736, 32'h00000000} /* (3, 31, 26) {real, imag} */,
  {32'hc4fc6adc, 32'h00000000} /* (3, 31, 25) {real, imag} */,
  {32'hc4dc8eda, 32'h00000000} /* (3, 31, 24) {real, imag} */,
  {32'hc4db2699, 32'h00000000} /* (3, 31, 23) {real, imag} */,
  {32'hc4922b81, 32'h00000000} /* (3, 31, 22) {real, imag} */,
  {32'hc20f1018, 32'h00000000} /* (3, 31, 21) {real, imag} */,
  {32'h440a0b3a, 32'h00000000} /* (3, 31, 20) {real, imag} */,
  {32'h44dab800, 32'h00000000} /* (3, 31, 19) {real, imag} */,
  {32'h44c096b5, 32'h00000000} /* (3, 31, 18) {real, imag} */,
  {32'h44cb8f74, 32'h00000000} /* (3, 31, 17) {real, imag} */,
  {32'h44f73c40, 32'h00000000} /* (3, 31, 16) {real, imag} */,
  {32'h4508c6a3, 32'h00000000} /* (3, 31, 15) {real, imag} */,
  {32'h457c111d, 32'h00000000} /* (3, 31, 14) {real, imag} */,
  {32'h4552471b, 32'h00000000} /* (3, 31, 13) {real, imag} */,
  {32'h451ede96, 32'h00000000} /* (3, 31, 12) {real, imag} */,
  {32'h45218717, 32'h00000000} /* (3, 31, 11) {real, imag} */,
  {32'h44821dfe, 32'h00000000} /* (3, 31, 10) {real, imag} */,
  {32'h40532100, 32'h00000000} /* (3, 31, 9) {real, imag} */,
  {32'hc4372774, 32'h00000000} /* (3, 31, 8) {real, imag} */,
  {32'hc36356e8, 32'h00000000} /* (3, 31, 7) {real, imag} */,
  {32'hc4078d68, 32'h00000000} /* (3, 31, 6) {real, imag} */,
  {32'hc45641b8, 32'h00000000} /* (3, 31, 5) {real, imag} */,
  {32'hc4651414, 32'h00000000} /* (3, 31, 4) {real, imag} */,
  {32'hc4bb96fc, 32'h00000000} /* (3, 31, 3) {real, imag} */,
  {32'hc4d1349b, 32'h00000000} /* (3, 31, 2) {real, imag} */,
  {32'hc4a21400, 32'h00000000} /* (3, 31, 1) {real, imag} */,
  {32'hc436b61f, 32'h00000000} /* (3, 31, 0) {real, imag} */,
  {32'hc41a887c, 32'h00000000} /* (3, 30, 31) {real, imag} */,
  {32'hc41fc224, 32'h00000000} /* (3, 30, 30) {real, imag} */,
  {32'hc497aa4b, 32'h00000000} /* (3, 30, 29) {real, imag} */,
  {32'hc50bc1a4, 32'h00000000} /* (3, 30, 28) {real, imag} */,
  {32'hc53ec1d4, 32'h00000000} /* (3, 30, 27) {real, imag} */,
  {32'hc539480c, 32'h00000000} /* (3, 30, 26) {real, imag} */,
  {32'hc503c31d, 32'h00000000} /* (3, 30, 25) {real, imag} */,
  {32'hc519a700, 32'h00000000} /* (3, 30, 24) {real, imag} */,
  {32'hc5049961, 32'h00000000} /* (3, 30, 23) {real, imag} */,
  {32'hc48f657b, 32'h00000000} /* (3, 30, 22) {real, imag} */,
  {32'hc3f66c90, 32'h00000000} /* (3, 30, 21) {real, imag} */,
  {32'h44c575d2, 32'h00000000} /* (3, 30, 20) {real, imag} */,
  {32'h453b38f2, 32'h00000000} /* (3, 30, 19) {real, imag} */,
  {32'h453b1db2, 32'h00000000} /* (3, 30, 18) {real, imag} */,
  {32'h45287038, 32'h00000000} /* (3, 30, 17) {real, imag} */,
  {32'h453cca23, 32'h00000000} /* (3, 30, 16) {real, imag} */,
  {32'h4551b135, 32'h00000000} /* (3, 30, 15) {real, imag} */,
  {32'h4552696a, 32'h00000000} /* (3, 30, 14) {real, imag} */,
  {32'h4564eef0, 32'h00000000} /* (3, 30, 13) {real, imag} */,
  {32'h455f3b50, 32'h00000000} /* (3, 30, 12) {real, imag} */,
  {32'h453445aa, 32'h00000000} /* (3, 30, 11) {real, imag} */,
  {32'h40d80000, 32'h00000000} /* (3, 30, 10) {real, imag} */,
  {32'hc4df0710, 32'h00000000} /* (3, 30, 9) {real, imag} */,
  {32'hc4b68a00, 32'h00000000} /* (3, 30, 8) {real, imag} */,
  {32'hc4e91731, 32'h00000000} /* (3, 30, 7) {real, imag} */,
  {32'hc5156cbe, 32'h00000000} /* (3, 30, 6) {real, imag} */,
  {32'hc480e035, 32'h00000000} /* (3, 30, 5) {real, imag} */,
  {32'hc502665f, 32'h00000000} /* (3, 30, 4) {real, imag} */,
  {32'hc508be6a, 32'h00000000} /* (3, 30, 3) {real, imag} */,
  {32'hc506e1d0, 32'h00000000} /* (3, 30, 2) {real, imag} */,
  {32'hc4638466, 32'h00000000} /* (3, 30, 1) {real, imag} */,
  {32'h43626f30, 32'h00000000} /* (3, 30, 0) {real, imag} */,
  {32'hc4901aba, 32'h00000000} /* (3, 29, 31) {real, imag} */,
  {32'hc4ef25ab, 32'h00000000} /* (3, 29, 30) {real, imag} */,
  {32'hc4c86a76, 32'h00000000} /* (3, 29, 29) {real, imag} */,
  {32'hc50f2656, 32'h00000000} /* (3, 29, 28) {real, imag} */,
  {32'hc5449ab6, 32'h00000000} /* (3, 29, 27) {real, imag} */,
  {32'hc51c9823, 32'h00000000} /* (3, 29, 26) {real, imag} */,
  {32'hc55e52e2, 32'h00000000} /* (3, 29, 25) {real, imag} */,
  {32'hc52c85d4, 32'h00000000} /* (3, 29, 24) {real, imag} */,
  {32'hc4f3f24b, 32'h00000000} /* (3, 29, 23) {real, imag} */,
  {32'hc49717e6, 32'h00000000} /* (3, 29, 22) {real, imag} */,
  {32'h438ae00a, 32'h00000000} /* (3, 29, 21) {real, imag} */,
  {32'h45271238, 32'h00000000} /* (3, 29, 20) {real, imag} */,
  {32'h45988884, 32'h00000000} /* (3, 29, 19) {real, imag} */,
  {32'h457d4768, 32'h00000000} /* (3, 29, 18) {real, imag} */,
  {32'h4585258e, 32'h00000000} /* (3, 29, 17) {real, imag} */,
  {32'h45732020, 32'h00000000} /* (3, 29, 16) {real, imag} */,
  {32'h4569c1a9, 32'h00000000} /* (3, 29, 15) {real, imag} */,
  {32'h4537db08, 32'h00000000} /* (3, 29, 14) {real, imag} */,
  {32'h45294937, 32'h00000000} /* (3, 29, 13) {real, imag} */,
  {32'h459b33ca, 32'h00000000} /* (3, 29, 12) {real, imag} */,
  {32'h45471cea, 32'h00000000} /* (3, 29, 11) {real, imag} */,
  {32'hc34e2ea0, 32'h00000000} /* (3, 29, 10) {real, imag} */,
  {32'hc4d53093, 32'h00000000} /* (3, 29, 9) {real, imag} */,
  {32'hc4c50a23, 32'h00000000} /* (3, 29, 8) {real, imag} */,
  {32'hc511b7ed, 32'h00000000} /* (3, 29, 7) {real, imag} */,
  {32'hc4f37c3c, 32'h00000000} /* (3, 29, 6) {real, imag} */,
  {32'hc4d1c0f0, 32'h00000000} /* (3, 29, 5) {real, imag} */,
  {32'hc53b74b0, 32'h00000000} /* (3, 29, 4) {real, imag} */,
  {32'hc520a7a2, 32'h00000000} /* (3, 29, 3) {real, imag} */,
  {32'hc484c263, 32'h00000000} /* (3, 29, 2) {real, imag} */,
  {32'hc46f7e4c, 32'h00000000} /* (3, 29, 1) {real, imag} */,
  {32'hc37151c0, 32'h00000000} /* (3, 29, 0) {real, imag} */,
  {32'hc43a0fce, 32'h00000000} /* (3, 28, 31) {real, imag} */,
  {32'hc4ce1f14, 32'h00000000} /* (3, 28, 30) {real, imag} */,
  {32'hc4fe597e, 32'h00000000} /* (3, 28, 29) {real, imag} */,
  {32'hc53ceb66, 32'h00000000} /* (3, 28, 28) {real, imag} */,
  {32'hc579f6fc, 32'h00000000} /* (3, 28, 27) {real, imag} */,
  {32'hc50b7db0, 32'h00000000} /* (3, 28, 26) {real, imag} */,
  {32'hc5224222, 32'h00000000} /* (3, 28, 25) {real, imag} */,
  {32'hc525512e, 32'h00000000} /* (3, 28, 24) {real, imag} */,
  {32'hc4e30009, 32'h00000000} /* (3, 28, 23) {real, imag} */,
  {32'hc4db1038, 32'h00000000} /* (3, 28, 22) {real, imag} */,
  {32'h43293808, 32'h00000000} /* (3, 28, 21) {real, imag} */,
  {32'h453b084b, 32'h00000000} /* (3, 28, 20) {real, imag} */,
  {32'h4584eeea, 32'h00000000} /* (3, 28, 19) {real, imag} */,
  {32'h455b5f24, 32'h00000000} /* (3, 28, 18) {real, imag} */,
  {32'h45878de0, 32'h00000000} /* (3, 28, 17) {real, imag} */,
  {32'h45949e0c, 32'h00000000} /* (3, 28, 16) {real, imag} */,
  {32'h456e967e, 32'h00000000} /* (3, 28, 15) {real, imag} */,
  {32'h456dedc0, 32'h00000000} /* (3, 28, 14) {real, imag} */,
  {32'h4537d0cd, 32'h00000000} /* (3, 28, 13) {real, imag} */,
  {32'h4582af68, 32'h00000000} /* (3, 28, 12) {real, imag} */,
  {32'h45086142, 32'h00000000} /* (3, 28, 11) {real, imag} */,
  {32'h42e96890, 32'h00000000} /* (3, 28, 10) {real, imag} */,
  {32'hc4a0da9a, 32'h00000000} /* (3, 28, 9) {real, imag} */,
  {32'hc50045d0, 32'h00000000} /* (3, 28, 8) {real, imag} */,
  {32'hc5164384, 32'h00000000} /* (3, 28, 7) {real, imag} */,
  {32'hc4c55710, 32'h00000000} /* (3, 28, 6) {real, imag} */,
  {32'hc5130f02, 32'h00000000} /* (3, 28, 5) {real, imag} */,
  {32'hc513646d, 32'h00000000} /* (3, 28, 4) {real, imag} */,
  {32'hc5244b86, 32'h00000000} /* (3, 28, 3) {real, imag} */,
  {32'hc4f9e90c, 32'h00000000} /* (3, 28, 2) {real, imag} */,
  {32'hc49f9f99, 32'h00000000} /* (3, 28, 1) {real, imag} */,
  {32'hc483ea0e, 32'h00000000} /* (3, 28, 0) {real, imag} */,
  {32'hc4a8fd90, 32'h00000000} /* (3, 27, 31) {real, imag} */,
  {32'hc4b787d8, 32'h00000000} /* (3, 27, 30) {real, imag} */,
  {32'hc508db52, 32'h00000000} /* (3, 27, 29) {real, imag} */,
  {32'hc50d38a0, 32'h00000000} /* (3, 27, 28) {real, imag} */,
  {32'hc528b52a, 32'h00000000} /* (3, 27, 27) {real, imag} */,
  {32'hc5498716, 32'h00000000} /* (3, 27, 26) {real, imag} */,
  {32'hc539c9b4, 32'h00000000} /* (3, 27, 25) {real, imag} */,
  {32'hc51bc031, 32'h00000000} /* (3, 27, 24) {real, imag} */,
  {32'hc53c62b5, 32'h00000000} /* (3, 27, 23) {real, imag} */,
  {32'hc4ecb3b0, 32'h00000000} /* (3, 27, 22) {real, imag} */,
  {32'h443a2772, 32'h00000000} /* (3, 27, 21) {real, imag} */,
  {32'h451ffcd2, 32'h00000000} /* (3, 27, 20) {real, imag} */,
  {32'h458d11c4, 32'h00000000} /* (3, 27, 19) {real, imag} */,
  {32'h457edb20, 32'h00000000} /* (3, 27, 18) {real, imag} */,
  {32'h457f511a, 32'h00000000} /* (3, 27, 17) {real, imag} */,
  {32'h45544078, 32'h00000000} /* (3, 27, 16) {real, imag} */,
  {32'h4569cab6, 32'h00000000} /* (3, 27, 15) {real, imag} */,
  {32'h45654f82, 32'h00000000} /* (3, 27, 14) {real, imag} */,
  {32'h458c6372, 32'h00000000} /* (3, 27, 13) {real, imag} */,
  {32'h455ffdc0, 32'h00000000} /* (3, 27, 12) {real, imag} */,
  {32'h451bc4f8, 32'h00000000} /* (3, 27, 11) {real, imag} */,
  {32'hc436426a, 32'h00000000} /* (3, 27, 10) {real, imag} */,
  {32'hc482867f, 32'h00000000} /* (3, 27, 9) {real, imag} */,
  {32'hc4c4d98a, 32'h00000000} /* (3, 27, 8) {real, imag} */,
  {32'hc4e55126, 32'h00000000} /* (3, 27, 7) {real, imag} */,
  {32'hc51db6da, 32'h00000000} /* (3, 27, 6) {real, imag} */,
  {32'hc5116bb0, 32'h00000000} /* (3, 27, 5) {real, imag} */,
  {32'hc529a094, 32'h00000000} /* (3, 27, 4) {real, imag} */,
  {32'hc532799c, 32'h00000000} /* (3, 27, 3) {real, imag} */,
  {32'hc502bf40, 32'h00000000} /* (3, 27, 2) {real, imag} */,
  {32'hc52336f4, 32'h00000000} /* (3, 27, 1) {real, imag} */,
  {32'hc4442df0, 32'h00000000} /* (3, 27, 0) {real, imag} */,
  {32'hc4a13810, 32'h00000000} /* (3, 26, 31) {real, imag} */,
  {32'hc4d316f9, 32'h00000000} /* (3, 26, 30) {real, imag} */,
  {32'hc5278ae0, 32'h00000000} /* (3, 26, 29) {real, imag} */,
  {32'hc5007c40, 32'h00000000} /* (3, 26, 28) {real, imag} */,
  {32'hc52f8935, 32'h00000000} /* (3, 26, 27) {real, imag} */,
  {32'hc53ad3d2, 32'h00000000} /* (3, 26, 26) {real, imag} */,
  {32'hc5510c09, 32'h00000000} /* (3, 26, 25) {real, imag} */,
  {32'hc5614bce, 32'h00000000} /* (3, 26, 24) {real, imag} */,
  {32'hc53d323b, 32'h00000000} /* (3, 26, 23) {real, imag} */,
  {32'hc4b799c0, 32'h00000000} /* (3, 26, 22) {real, imag} */,
  {32'h4489fb7c, 32'h00000000} /* (3, 26, 21) {real, imag} */,
  {32'h4574d1aa, 32'h00000000} /* (3, 26, 20) {real, imag} */,
  {32'h457bd35c, 32'h00000000} /* (3, 26, 19) {real, imag} */,
  {32'h458d036c, 32'h00000000} /* (3, 26, 18) {real, imag} */,
  {32'h458e55a0, 32'h00000000} /* (3, 26, 17) {real, imag} */,
  {32'h456657d8, 32'h00000000} /* (3, 26, 16) {real, imag} */,
  {32'h4599ad34, 32'h00000000} /* (3, 26, 15) {real, imag} */,
  {32'h45812350, 32'h00000000} /* (3, 26, 14) {real, imag} */,
  {32'h4568c68c, 32'h00000000} /* (3, 26, 13) {real, imag} */,
  {32'h455a3dac, 32'h00000000} /* (3, 26, 12) {real, imag} */,
  {32'h450b2b35, 32'h00000000} /* (3, 26, 11) {real, imag} */,
  {32'h4419191e, 32'h00000000} /* (3, 26, 10) {real, imag} */,
  {32'hc4a059b6, 32'h00000000} /* (3, 26, 9) {real, imag} */,
  {32'hc50eb6a2, 32'h00000000} /* (3, 26, 8) {real, imag} */,
  {32'hc5013339, 32'h00000000} /* (3, 26, 7) {real, imag} */,
  {32'hc4f86c1e, 32'h00000000} /* (3, 26, 6) {real, imag} */,
  {32'hc541736c, 32'h00000000} /* (3, 26, 5) {real, imag} */,
  {32'hc5003ca4, 32'h00000000} /* (3, 26, 4) {real, imag} */,
  {32'hc4ee0d44, 32'h00000000} /* (3, 26, 3) {real, imag} */,
  {32'hc5350b19, 32'h00000000} /* (3, 26, 2) {real, imag} */,
  {32'hc50266fe, 32'h00000000} /* (3, 26, 1) {real, imag} */,
  {32'hc4be7748, 32'h00000000} /* (3, 26, 0) {real, imag} */,
  {32'hc4cc1e6c, 32'h00000000} /* (3, 25, 31) {real, imag} */,
  {32'hc4ee8c16, 32'h00000000} /* (3, 25, 30) {real, imag} */,
  {32'hc52c4a8e, 32'h00000000} /* (3, 25, 29) {real, imag} */,
  {32'hc558de99, 32'h00000000} /* (3, 25, 28) {real, imag} */,
  {32'hc56afe19, 32'h00000000} /* (3, 25, 27) {real, imag} */,
  {32'hc57ad04e, 32'h00000000} /* (3, 25, 26) {real, imag} */,
  {32'hc52bb6ac, 32'h00000000} /* (3, 25, 25) {real, imag} */,
  {32'hc548cb8f, 32'h00000000} /* (3, 25, 24) {real, imag} */,
  {32'hc517ec20, 32'h00000000} /* (3, 25, 23) {real, imag} */,
  {32'hc4c378f2, 32'h00000000} /* (3, 25, 22) {real, imag} */,
  {32'h44807216, 32'h00000000} /* (3, 25, 21) {real, imag} */,
  {32'h4556f784, 32'h00000000} /* (3, 25, 20) {real, imag} */,
  {32'h458a4df9, 32'h00000000} /* (3, 25, 19) {real, imag} */,
  {32'h4597ef05, 32'h00000000} /* (3, 25, 18) {real, imag} */,
  {32'h459cd21e, 32'h00000000} /* (3, 25, 17) {real, imag} */,
  {32'h458c6fa8, 32'h00000000} /* (3, 25, 16) {real, imag} */,
  {32'h459888d1, 32'h00000000} /* (3, 25, 15) {real, imag} */,
  {32'h458b52e0, 32'h00000000} /* (3, 25, 14) {real, imag} */,
  {32'h4540a066, 32'h00000000} /* (3, 25, 13) {real, imag} */,
  {32'h456a5dc5, 32'h00000000} /* (3, 25, 12) {real, imag} */,
  {32'h4509332d, 32'h00000000} /* (3, 25, 11) {real, imag} */,
  {32'h43f4f244, 32'h00000000} /* (3, 25, 10) {real, imag} */,
  {32'hc4f1d6dc, 32'h00000000} /* (3, 25, 9) {real, imag} */,
  {32'hc513261b, 32'h00000000} /* (3, 25, 8) {real, imag} */,
  {32'hc52315cc, 32'h00000000} /* (3, 25, 7) {real, imag} */,
  {32'hc519dc89, 32'h00000000} /* (3, 25, 6) {real, imag} */,
  {32'hc52ca71c, 32'h00000000} /* (3, 25, 5) {real, imag} */,
  {32'hc52f069c, 32'h00000000} /* (3, 25, 4) {real, imag} */,
  {32'hc50105ac, 32'h00000000} /* (3, 25, 3) {real, imag} */,
  {32'hc53a448a, 32'h00000000} /* (3, 25, 2) {real, imag} */,
  {32'hc52aeb30, 32'h00000000} /* (3, 25, 1) {real, imag} */,
  {32'hc4e70202, 32'h00000000} /* (3, 25, 0) {real, imag} */,
  {32'hc4de0a0c, 32'h00000000} /* (3, 24, 31) {real, imag} */,
  {32'hc54e94d0, 32'h00000000} /* (3, 24, 30) {real, imag} */,
  {32'hc51c39d8, 32'h00000000} /* (3, 24, 29) {real, imag} */,
  {32'hc58ad91a, 32'h00000000} /* (3, 24, 28) {real, imag} */,
  {32'hc535732c, 32'h00000000} /* (3, 24, 27) {real, imag} */,
  {32'hc52ef4c2, 32'h00000000} /* (3, 24, 26) {real, imag} */,
  {32'hc57f637b, 32'h00000000} /* (3, 24, 25) {real, imag} */,
  {32'hc51cbb55, 32'h00000000} /* (3, 24, 24) {real, imag} */,
  {32'hc52a23af, 32'h00000000} /* (3, 24, 23) {real, imag} */,
  {32'hc48f239c, 32'h00000000} /* (3, 24, 22) {real, imag} */,
  {32'h4488520e, 32'h00000000} /* (3, 24, 21) {real, imag} */,
  {32'h45388117, 32'h00000000} /* (3, 24, 20) {real, imag} */,
  {32'h45703168, 32'h00000000} /* (3, 24, 19) {real, imag} */,
  {32'h458d5fd6, 32'h00000000} /* (3, 24, 18) {real, imag} */,
  {32'h45908ae8, 32'h00000000} /* (3, 24, 17) {real, imag} */,
  {32'h45834b91, 32'h00000000} /* (3, 24, 16) {real, imag} */,
  {32'h4584bf05, 32'h00000000} /* (3, 24, 15) {real, imag} */,
  {32'h45a221bc, 32'h00000000} /* (3, 24, 14) {real, imag} */,
  {32'h453a207e, 32'h00000000} /* (3, 24, 13) {real, imag} */,
  {32'h456ee08c, 32'h00000000} /* (3, 24, 12) {real, imag} */,
  {32'h450dda9e, 32'h00000000} /* (3, 24, 11) {real, imag} */,
  {32'hc2f65840, 32'h00000000} /* (3, 24, 10) {real, imag} */,
  {32'hc4ec917a, 32'h00000000} /* (3, 24, 9) {real, imag} */,
  {32'hc52b76df, 32'h00000000} /* (3, 24, 8) {real, imag} */,
  {32'hc505bfb7, 32'h00000000} /* (3, 24, 7) {real, imag} */,
  {32'hc527c7a0, 32'h00000000} /* (3, 24, 6) {real, imag} */,
  {32'hc5150a1d, 32'h00000000} /* (3, 24, 5) {real, imag} */,
  {32'hc50777f9, 32'h00000000} /* (3, 24, 4) {real, imag} */,
  {32'hc52d70f8, 32'h00000000} /* (3, 24, 3) {real, imag} */,
  {32'hc535bccf, 32'h00000000} /* (3, 24, 2) {real, imag} */,
  {32'hc528bed4, 32'h00000000} /* (3, 24, 1) {real, imag} */,
  {32'hc521b0a4, 32'h00000000} /* (3, 24, 0) {real, imag} */,
  {32'hc50af076, 32'h00000000} /* (3, 23, 31) {real, imag} */,
  {32'hc513759b, 32'h00000000} /* (3, 23, 30) {real, imag} */,
  {32'hc5290bcc, 32'h00000000} /* (3, 23, 29) {real, imag} */,
  {32'hc5453d8a, 32'h00000000} /* (3, 23, 28) {real, imag} */,
  {32'hc55f757a, 32'h00000000} /* (3, 23, 27) {real, imag} */,
  {32'hc52af946, 32'h00000000} /* (3, 23, 26) {real, imag} */,
  {32'hc51fabfa, 32'h00000000} /* (3, 23, 25) {real, imag} */,
  {32'hc5054f24, 32'h00000000} /* (3, 23, 24) {real, imag} */,
  {32'hc47341c7, 32'h00000000} /* (3, 23, 23) {real, imag} */,
  {32'hc4a19a94, 32'h00000000} /* (3, 23, 22) {real, imag} */,
  {32'h446c14ae, 32'h00000000} /* (3, 23, 21) {real, imag} */,
  {32'h45314712, 32'h00000000} /* (3, 23, 20) {real, imag} */,
  {32'h45502578, 32'h00000000} /* (3, 23, 19) {real, imag} */,
  {32'h456961b0, 32'h00000000} /* (3, 23, 18) {real, imag} */,
  {32'h45611db0, 32'h00000000} /* (3, 23, 17) {real, imag} */,
  {32'h4557d36a, 32'h00000000} /* (3, 23, 16) {real, imag} */,
  {32'h455694a4, 32'h00000000} /* (3, 23, 15) {real, imag} */,
  {32'h4582d140, 32'h00000000} /* (3, 23, 14) {real, imag} */,
  {32'h456f1760, 32'h00000000} /* (3, 23, 13) {real, imag} */,
  {32'h454f2654, 32'h00000000} /* (3, 23, 12) {real, imag} */,
  {32'h451789d2, 32'h00000000} /* (3, 23, 11) {real, imag} */,
  {32'hc3ece84c, 32'h00000000} /* (3, 23, 10) {real, imag} */,
  {32'hc4bb778e, 32'h00000000} /* (3, 23, 9) {real, imag} */,
  {32'hc505192c, 32'h00000000} /* (3, 23, 8) {real, imag} */,
  {32'hc508d531, 32'h00000000} /* (3, 23, 7) {real, imag} */,
  {32'hc4f78ec4, 32'h00000000} /* (3, 23, 6) {real, imag} */,
  {32'hc518e564, 32'h00000000} /* (3, 23, 5) {real, imag} */,
  {32'hc4d7b000, 32'h00000000} /* (3, 23, 4) {real, imag} */,
  {32'hc570bdf8, 32'h00000000} /* (3, 23, 3) {real, imag} */,
  {32'hc540e03c, 32'h00000000} /* (3, 23, 2) {real, imag} */,
  {32'hc50b80fa, 32'h00000000} /* (3, 23, 1) {real, imag} */,
  {32'hc5023704, 32'h00000000} /* (3, 23, 0) {real, imag} */,
  {32'hc4b1d918, 32'h00000000} /* (3, 22, 31) {real, imag} */,
  {32'hc52206da, 32'h00000000} /* (3, 22, 30) {real, imag} */,
  {32'hc52b6a6c, 32'h00000000} /* (3, 22, 29) {real, imag} */,
  {32'hc51b7d8b, 32'h00000000} /* (3, 22, 28) {real, imag} */,
  {32'hc5384bbb, 32'h00000000} /* (3, 22, 27) {real, imag} */,
  {32'hc52c0666, 32'h00000000} /* (3, 22, 26) {real, imag} */,
  {32'hc47ba698, 32'h00000000} /* (3, 22, 25) {real, imag} */,
  {32'hc49d29c8, 32'h00000000} /* (3, 22, 24) {real, imag} */,
  {32'hc43b0770, 32'h00000000} /* (3, 22, 23) {real, imag} */,
  {32'h43842fea, 32'h00000000} /* (3, 22, 22) {real, imag} */,
  {32'h4474e3d1, 32'h00000000} /* (3, 22, 21) {real, imag} */,
  {32'h44fa397d, 32'h00000000} /* (3, 22, 20) {real, imag} */,
  {32'h45152ff5, 32'h00000000} /* (3, 22, 19) {real, imag} */,
  {32'h4528cfee, 32'h00000000} /* (3, 22, 18) {real, imag} */,
  {32'h45547ca4, 32'h00000000} /* (3, 22, 17) {real, imag} */,
  {32'h450c5dc4, 32'h00000000} /* (3, 22, 16) {real, imag} */,
  {32'h4506b980, 32'h00000000} /* (3, 22, 15) {real, imag} */,
  {32'h454363b6, 32'h00000000} /* (3, 22, 14) {real, imag} */,
  {32'h455a2e96, 32'h00000000} /* (3, 22, 13) {real, imag} */,
  {32'h44f4faa2, 32'h00000000} /* (3, 22, 12) {real, imag} */,
  {32'h447ab80c, 32'h00000000} /* (3, 22, 11) {real, imag} */,
  {32'hc20fdc60, 32'h00000000} /* (3, 22, 10) {real, imag} */,
  {32'hc4d0b78c, 32'h00000000} /* (3, 22, 9) {real, imag} */,
  {32'hc4ae8664, 32'h00000000} /* (3, 22, 8) {real, imag} */,
  {32'hc51d7e1e, 32'h00000000} /* (3, 22, 7) {real, imag} */,
  {32'hc4aada80, 32'h00000000} /* (3, 22, 6) {real, imag} */,
  {32'hc513dabb, 32'h00000000} /* (3, 22, 5) {real, imag} */,
  {32'hc4dc0ddf, 32'h00000000} /* (3, 22, 4) {real, imag} */,
  {32'hc4eaafd6, 32'h00000000} /* (3, 22, 3) {real, imag} */,
  {32'hc53243fc, 32'h00000000} /* (3, 22, 2) {real, imag} */,
  {32'hc5115caa, 32'h00000000} /* (3, 22, 1) {real, imag} */,
  {32'hc4a130d5, 32'h00000000} /* (3, 22, 0) {real, imag} */,
  {32'hc2c90cd4, 32'h00000000} /* (3, 21, 31) {real, imag} */,
  {32'hc2843ef0, 32'h00000000} /* (3, 21, 30) {real, imag} */,
  {32'h443a0570, 32'h00000000} /* (3, 21, 29) {real, imag} */,
  {32'hc305bb30, 32'h00000000} /* (3, 21, 28) {real, imag} */,
  {32'hc4658f06, 32'h00000000} /* (3, 21, 27) {real, imag} */,
  {32'hc37cdb42, 32'h00000000} /* (3, 21, 26) {real, imag} */,
  {32'h44238b95, 32'h00000000} /* (3, 21, 25) {real, imag} */,
  {32'h446bd36a, 32'h00000000} /* (3, 21, 24) {real, imag} */,
  {32'hc2981c98, 32'h00000000} /* (3, 21, 23) {real, imag} */,
  {32'h4411f246, 32'h00000000} /* (3, 21, 22) {real, imag} */,
  {32'h44267260, 32'h00000000} /* (3, 21, 21) {real, imag} */,
  {32'h442e3aa5, 32'h00000000} /* (3, 21, 20) {real, imag} */,
  {32'h44a0ab10, 32'h00000000} /* (3, 21, 19) {real, imag} */,
  {32'h44bbc4af, 32'h00000000} /* (3, 21, 18) {real, imag} */,
  {32'h44d27d18, 32'h00000000} /* (3, 21, 17) {real, imag} */,
  {32'h44f08758, 32'h00000000} /* (3, 21, 16) {real, imag} */,
  {32'h444eff60, 32'h00000000} /* (3, 21, 15) {real, imag} */,
  {32'h4498df14, 32'h00000000} /* (3, 21, 14) {real, imag} */,
  {32'h4499a497, 32'h00000000} /* (3, 21, 13) {real, imag} */,
  {32'h43f0f914, 32'h00000000} /* (3, 21, 12) {real, imag} */,
  {32'h43ad4554, 32'h00000000} /* (3, 21, 11) {real, imag} */,
  {32'h424e3948, 32'h00000000} /* (3, 21, 10) {real, imag} */,
  {32'hc4829210, 32'h00000000} /* (3, 21, 9) {real, imag} */,
  {32'hc439d616, 32'h00000000} /* (3, 21, 8) {real, imag} */,
  {32'h43e5cc74, 32'h00000000} /* (3, 21, 7) {real, imag} */,
  {32'hc29a8f66, 32'h00000000} /* (3, 21, 6) {real, imag} */,
  {32'hc413950a, 32'h00000000} /* (3, 21, 5) {real, imag} */,
  {32'hc43a0ea1, 32'h00000000} /* (3, 21, 4) {real, imag} */,
  {32'hc4a43e50, 32'h00000000} /* (3, 21, 3) {real, imag} */,
  {32'hc467534e, 32'h00000000} /* (3, 21, 2) {real, imag} */,
  {32'hc3ead342, 32'h00000000} /* (3, 21, 1) {real, imag} */,
  {32'hc3ac33d0, 32'h00000000} /* (3, 21, 0) {real, imag} */,
  {32'h44c952b0, 32'h00000000} /* (3, 20, 31) {real, imag} */,
  {32'h44ea03c2, 32'h00000000} /* (3, 20, 30) {real, imag} */,
  {32'h45242160, 32'h00000000} /* (3, 20, 29) {real, imag} */,
  {32'h451a25b9, 32'h00000000} /* (3, 20, 28) {real, imag} */,
  {32'h451a376c, 32'h00000000} /* (3, 20, 27) {real, imag} */,
  {32'h450b2ded, 32'h00000000} /* (3, 20, 26) {real, imag} */,
  {32'h45684d4c, 32'h00000000} /* (3, 20, 25) {real, imag} */,
  {32'h45503b52, 32'h00000000} /* (3, 20, 24) {real, imag} */,
  {32'h4526c3d4, 32'h00000000} /* (3, 20, 23) {real, imag} */,
  {32'h44a9b234, 32'h00000000} /* (3, 20, 22) {real, imag} */,
  {32'h441dad33, 32'h00000000} /* (3, 20, 21) {real, imag} */,
  {32'hc483f1ec, 32'h00000000} /* (3, 20, 20) {real, imag} */,
  {32'hc3d2790e, 32'h00000000} /* (3, 20, 19) {real, imag} */,
  {32'hc4077394, 32'h00000000} /* (3, 20, 18) {real, imag} */,
  {32'hc38c96ee, 32'h00000000} /* (3, 20, 17) {real, imag} */,
  {32'hc3b5ae46, 32'h00000000} /* (3, 20, 16) {real, imag} */,
  {32'hc4389b2c, 32'h00000000} /* (3, 20, 15) {real, imag} */,
  {32'hc4817f64, 32'h00000000} /* (3, 20, 14) {real, imag} */,
  {32'hc470058a, 32'h00000000} /* (3, 20, 13) {real, imag} */,
  {32'hc4ee1e26, 32'h00000000} /* (3, 20, 12) {real, imag} */,
  {32'hc387fb4c, 32'h00000000} /* (3, 20, 11) {real, imag} */,
  {32'h4496040e, 32'h00000000} /* (3, 20, 10) {real, imag} */,
  {32'h43e3a3f4, 32'h00000000} /* (3, 20, 9) {real, imag} */,
  {32'h43c642f0, 32'h00000000} /* (3, 20, 8) {real, imag} */,
  {32'h45233efc, 32'h00000000} /* (3, 20, 7) {real, imag} */,
  {32'h44cf58e8, 32'h00000000} /* (3, 20, 6) {real, imag} */,
  {32'h4519614c, 32'h00000000} /* (3, 20, 5) {real, imag} */,
  {32'h44bb45aa, 32'h00000000} /* (3, 20, 4) {real, imag} */,
  {32'h44540d39, 32'h00000000} /* (3, 20, 3) {real, imag} */,
  {32'h44951b6a, 32'h00000000} /* (3, 20, 2) {real, imag} */,
  {32'h4444c2a5, 32'h00000000} /* (3, 20, 1) {real, imag} */,
  {32'h441633ed, 32'h00000000} /* (3, 20, 0) {real, imag} */,
  {32'h4501a14b, 32'h00000000} /* (3, 19, 31) {real, imag} */,
  {32'h4516ab52, 32'h00000000} /* (3, 19, 30) {real, imag} */,
  {32'h45303f84, 32'h00000000} /* (3, 19, 29) {real, imag} */,
  {32'h454c38dd, 32'h00000000} /* (3, 19, 28) {real, imag} */,
  {32'h455d17ac, 32'h00000000} /* (3, 19, 27) {real, imag} */,
  {32'h453173a2, 32'h00000000} /* (3, 19, 26) {real, imag} */,
  {32'h459143fb, 32'h00000000} /* (3, 19, 25) {real, imag} */,
  {32'h456f9986, 32'h00000000} /* (3, 19, 24) {real, imag} */,
  {32'h45258628, 32'h00000000} /* (3, 19, 23) {real, imag} */,
  {32'h45000f7c, 32'h00000000} /* (3, 19, 22) {real, imag} */,
  {32'h43295180, 32'h00000000} /* (3, 19, 21) {real, imag} */,
  {32'hc4f02a24, 32'h00000000} /* (3, 19, 20) {real, imag} */,
  {32'hc4b97f5a, 32'h00000000} /* (3, 19, 19) {real, imag} */,
  {32'hc4e43528, 32'h00000000} /* (3, 19, 18) {real, imag} */,
  {32'hc508a9e9, 32'h00000000} /* (3, 19, 17) {real, imag} */,
  {32'hc4dbe28d, 32'h00000000} /* (3, 19, 16) {real, imag} */,
  {32'hc50a6ac3, 32'h00000000} /* (3, 19, 15) {real, imag} */,
  {32'hc4f45e59, 32'h00000000} /* (3, 19, 14) {real, imag} */,
  {32'hc4ff0454, 32'h00000000} /* (3, 19, 13) {real, imag} */,
  {32'hc531b68b, 32'h00000000} /* (3, 19, 12) {real, imag} */,
  {32'hc4da3cb5, 32'h00000000} /* (3, 19, 11) {real, imag} */,
  {32'h44a2de5d, 32'h00000000} /* (3, 19, 10) {real, imag} */,
  {32'h44df0e04, 32'h00000000} /* (3, 19, 9) {real, imag} */,
  {32'h4503a99a, 32'h00000000} /* (3, 19, 8) {real, imag} */,
  {32'h4540aa6c, 32'h00000000} /* (3, 19, 7) {real, imag} */,
  {32'h44eb1116, 32'h00000000} /* (3, 19, 6) {real, imag} */,
  {32'h45301320, 32'h00000000} /* (3, 19, 5) {real, imag} */,
  {32'h4537ef96, 32'h00000000} /* (3, 19, 4) {real, imag} */,
  {32'h44fd30fa, 32'h00000000} /* (3, 19, 3) {real, imag} */,
  {32'h44d60c0e, 32'h00000000} /* (3, 19, 2) {real, imag} */,
  {32'h4514ad97, 32'h00000000} /* (3, 19, 1) {real, imag} */,
  {32'h44df156d, 32'h00000000} /* (3, 19, 0) {real, imag} */,
  {32'h4502f490, 32'h00000000} /* (3, 18, 31) {real, imag} */,
  {32'h4528215e, 32'h00000000} /* (3, 18, 30) {real, imag} */,
  {32'h45400dd1, 32'h00000000} /* (3, 18, 29) {real, imag} */,
  {32'h45724b2f, 32'h00000000} /* (3, 18, 28) {real, imag} */,
  {32'h452bcebb, 32'h00000000} /* (3, 18, 27) {real, imag} */,
  {32'h4588edd4, 32'h00000000} /* (3, 18, 26) {real, imag} */,
  {32'h45512452, 32'h00000000} /* (3, 18, 25) {real, imag} */,
  {32'h458f37d9, 32'h00000000} /* (3, 18, 24) {real, imag} */,
  {32'h453630a1, 32'h00000000} /* (3, 18, 23) {real, imag} */,
  {32'h45009ba0, 32'h00000000} /* (3, 18, 22) {real, imag} */,
  {32'h449e6aaa, 32'h00000000} /* (3, 18, 21) {real, imag} */,
  {32'hc51b19cf, 32'h00000000} /* (3, 18, 20) {real, imag} */,
  {32'hc4a7cf11, 32'h00000000} /* (3, 18, 19) {real, imag} */,
  {32'hc53fd2c5, 32'h00000000} /* (3, 18, 18) {real, imag} */,
  {32'hc572f800, 32'h00000000} /* (3, 18, 17) {real, imag} */,
  {32'hc4e6b550, 32'h00000000} /* (3, 18, 16) {real, imag} */,
  {32'hc54ff3a4, 32'h00000000} /* (3, 18, 15) {real, imag} */,
  {32'hc54e17b2, 32'h00000000} /* (3, 18, 14) {real, imag} */,
  {32'hc54dc1a9, 32'h00000000} /* (3, 18, 13) {real, imag} */,
  {32'hc55b71f5, 32'h00000000} /* (3, 18, 12) {real, imag} */,
  {32'hc52ee02d, 32'h00000000} /* (3, 18, 11) {real, imag} */,
  {32'h426d8200, 32'h00000000} /* (3, 18, 10) {real, imag} */,
  {32'h44f27ea4, 32'h00000000} /* (3, 18, 9) {real, imag} */,
  {32'h45641e0e, 32'h00000000} /* (3, 18, 8) {real, imag} */,
  {32'h455698c7, 32'h00000000} /* (3, 18, 7) {real, imag} */,
  {32'h452c7380, 32'h00000000} /* (3, 18, 6) {real, imag} */,
  {32'h45488769, 32'h00000000} /* (3, 18, 5) {real, imag} */,
  {32'h45391abd, 32'h00000000} /* (3, 18, 4) {real, imag} */,
  {32'h453cda9c, 32'h00000000} /* (3, 18, 3) {real, imag} */,
  {32'h451ae391, 32'h00000000} /* (3, 18, 2) {real, imag} */,
  {32'h45137a3c, 32'h00000000} /* (3, 18, 1) {real, imag} */,
  {32'h44f93d20, 32'h00000000} /* (3, 18, 0) {real, imag} */,
  {32'h4532e206, 32'h00000000} /* (3, 17, 31) {real, imag} */,
  {32'h4544ffa2, 32'h00000000} /* (3, 17, 30) {real, imag} */,
  {32'h454a3b96, 32'h00000000} /* (3, 17, 29) {real, imag} */,
  {32'h4565297f, 32'h00000000} /* (3, 17, 28) {real, imag} */,
  {32'h45620186, 32'h00000000} /* (3, 17, 27) {real, imag} */,
  {32'h458a255c, 32'h00000000} /* (3, 17, 26) {real, imag} */,
  {32'h4568c7f5, 32'h00000000} /* (3, 17, 25) {real, imag} */,
  {32'h454713c4, 32'h00000000} /* (3, 17, 24) {real, imag} */,
  {32'h45410a98, 32'h00000000} /* (3, 17, 23) {real, imag} */,
  {32'h45143407, 32'h00000000} /* (3, 17, 22) {real, imag} */,
  {32'h44140cde, 32'h00000000} /* (3, 17, 21) {real, imag} */,
  {32'hc5031da5, 32'h00000000} /* (3, 17, 20) {real, imag} */,
  {32'hc508c8f4, 32'h00000000} /* (3, 17, 19) {real, imag} */,
  {32'hc5418e12, 32'h00000000} /* (3, 17, 18) {real, imag} */,
  {32'hc54ebb8d, 32'h00000000} /* (3, 17, 17) {real, imag} */,
  {32'hc56e093a, 32'h00000000} /* (3, 17, 16) {real, imag} */,
  {32'hc556a6c0, 32'h00000000} /* (3, 17, 15) {real, imag} */,
  {32'hc5533d56, 32'h00000000} /* (3, 17, 14) {real, imag} */,
  {32'hc532f204, 32'h00000000} /* (3, 17, 13) {real, imag} */,
  {32'hc4fa8c9e, 32'h00000000} /* (3, 17, 12) {real, imag} */,
  {32'hc500f6c8, 32'h00000000} /* (3, 17, 11) {real, imag} */,
  {32'h43d220c8, 32'h00000000} /* (3, 17, 10) {real, imag} */,
  {32'h44f703ae, 32'h00000000} /* (3, 17, 9) {real, imag} */,
  {32'h45161002, 32'h00000000} /* (3, 17, 8) {real, imag} */,
  {32'h453a2748, 32'h00000000} /* (3, 17, 7) {real, imag} */,
  {32'h4544cc6d, 32'h00000000} /* (3, 17, 6) {real, imag} */,
  {32'h454c61b8, 32'h00000000} /* (3, 17, 5) {real, imag} */,
  {32'h4580afff, 32'h00000000} /* (3, 17, 4) {real, imag} */,
  {32'h45392a08, 32'h00000000} /* (3, 17, 3) {real, imag} */,
  {32'h4513a820, 32'h00000000} /* (3, 17, 2) {real, imag} */,
  {32'h45081bc9, 32'h00000000} /* (3, 17, 1) {real, imag} */,
  {32'h451bbd0a, 32'h00000000} /* (3, 17, 0) {real, imag} */,
  {32'h4533b01e, 32'h00000000} /* (3, 16, 31) {real, imag} */,
  {32'h4585fbc7, 32'h00000000} /* (3, 16, 30) {real, imag} */,
  {32'h4557bb1c, 32'h00000000} /* (3, 16, 29) {real, imag} */,
  {32'h454490a7, 32'h00000000} /* (3, 16, 28) {real, imag} */,
  {32'h4547e14c, 32'h00000000} /* (3, 16, 27) {real, imag} */,
  {32'h4540251a, 32'h00000000} /* (3, 16, 26) {real, imag} */,
  {32'h456d7d37, 32'h00000000} /* (3, 16, 25) {real, imag} */,
  {32'h454a54b1, 32'h00000000} /* (3, 16, 24) {real, imag} */,
  {32'h452da77e, 32'h00000000} /* (3, 16, 23) {real, imag} */,
  {32'h450f56a8, 32'h00000000} /* (3, 16, 22) {real, imag} */,
  {32'h446f5164, 32'h00000000} /* (3, 16, 21) {real, imag} */,
  {32'hc4f2c0c3, 32'h00000000} /* (3, 16, 20) {real, imag} */,
  {32'hc530c043, 32'h00000000} /* (3, 16, 19) {real, imag} */,
  {32'hc54d0e9c, 32'h00000000} /* (3, 16, 18) {real, imag} */,
  {32'hc57ba7ff, 32'h00000000} /* (3, 16, 17) {real, imag} */,
  {32'hc58aea6b, 32'h00000000} /* (3, 16, 16) {real, imag} */,
  {32'hc5886bf6, 32'h00000000} /* (3, 16, 15) {real, imag} */,
  {32'hc5399f40, 32'h00000000} /* (3, 16, 14) {real, imag} */,
  {32'hc57f0e98, 32'h00000000} /* (3, 16, 13) {real, imag} */,
  {32'hc523b5fb, 32'h00000000} /* (3, 16, 12) {real, imag} */,
  {32'hc4e0c920, 32'h00000000} /* (3, 16, 11) {real, imag} */,
  {32'h43d08ec4, 32'h00000000} /* (3, 16, 10) {real, imag} */,
  {32'h452282d5, 32'h00000000} /* (3, 16, 9) {real, imag} */,
  {32'h45238417, 32'h00000000} /* (3, 16, 8) {real, imag} */,
  {32'h45451afa, 32'h00000000} /* (3, 16, 7) {real, imag} */,
  {32'h45307dc2, 32'h00000000} /* (3, 16, 6) {real, imag} */,
  {32'h45403dc2, 32'h00000000} /* (3, 16, 5) {real, imag} */,
  {32'h454f49e6, 32'h00000000} /* (3, 16, 4) {real, imag} */,
  {32'h455abaa5, 32'h00000000} /* (3, 16, 3) {real, imag} */,
  {32'h4557bc7e, 32'h00000000} /* (3, 16, 2) {real, imag} */,
  {32'h45574b97, 32'h00000000} /* (3, 16, 1) {real, imag} */,
  {32'h45505582, 32'h00000000} /* (3, 16, 0) {real, imag} */,
  {32'h45446c07, 32'h00000000} /* (3, 15, 31) {real, imag} */,
  {32'h4565294a, 32'h00000000} /* (3, 15, 30) {real, imag} */,
  {32'h454e96a4, 32'h00000000} /* (3, 15, 29) {real, imag} */,
  {32'h453be63a, 32'h00000000} /* (3, 15, 28) {real, imag} */,
  {32'h45773a66, 32'h00000000} /* (3, 15, 27) {real, imag} */,
  {32'h455d9862, 32'h00000000} /* (3, 15, 26) {real, imag} */,
  {32'h455dacc5, 32'h00000000} /* (3, 15, 25) {real, imag} */,
  {32'h45537f79, 32'h00000000} /* (3, 15, 24) {real, imag} */,
  {32'h45609618, 32'h00000000} /* (3, 15, 23) {real, imag} */,
  {32'h455a0470, 32'h00000000} /* (3, 15, 22) {real, imag} */,
  {32'h449e4927, 32'h00000000} /* (3, 15, 21) {real, imag} */,
  {32'hc4ad0ca1, 32'h00000000} /* (3, 15, 20) {real, imag} */,
  {32'hc50c7bce, 32'h00000000} /* (3, 15, 19) {real, imag} */,
  {32'hc5295302, 32'h00000000} /* (3, 15, 18) {real, imag} */,
  {32'hc5530c99, 32'h00000000} /* (3, 15, 17) {real, imag} */,
  {32'hc53fb71f, 32'h00000000} /* (3, 15, 16) {real, imag} */,
  {32'hc555eb91, 32'h00000000} /* (3, 15, 15) {real, imag} */,
  {32'hc5592ace, 32'h00000000} /* (3, 15, 14) {real, imag} */,
  {32'hc53833ec, 32'h00000000} /* (3, 15, 13) {real, imag} */,
  {32'hc544f888, 32'h00000000} /* (3, 15, 12) {real, imag} */,
  {32'hc4be60f7, 32'h00000000} /* (3, 15, 11) {real, imag} */,
  {32'h44368860, 32'h00000000} /* (3, 15, 10) {real, imag} */,
  {32'h45145de9, 32'h00000000} /* (3, 15, 9) {real, imag} */,
  {32'h450a96a3, 32'h00000000} /* (3, 15, 8) {real, imag} */,
  {32'h454d3fec, 32'h00000000} /* (3, 15, 7) {real, imag} */,
  {32'h452621a4, 32'h00000000} /* (3, 15, 6) {real, imag} */,
  {32'h4563d254, 32'h00000000} /* (3, 15, 5) {real, imag} */,
  {32'h452cade6, 32'h00000000} /* (3, 15, 4) {real, imag} */,
  {32'h455bb496, 32'h00000000} /* (3, 15, 3) {real, imag} */,
  {32'h456c4bf0, 32'h00000000} /* (3, 15, 2) {real, imag} */,
  {32'h453f8395, 32'h00000000} /* (3, 15, 1) {real, imag} */,
  {32'h455026ef, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'h4531e2a8, 32'h00000000} /* (3, 14, 31) {real, imag} */,
  {32'h4559b8fa, 32'h00000000} /* (3, 14, 30) {real, imag} */,
  {32'h45529fd4, 32'h00000000} /* (3, 14, 29) {real, imag} */,
  {32'h456c82c7, 32'h00000000} /* (3, 14, 28) {real, imag} */,
  {32'h457ede55, 32'h00000000} /* (3, 14, 27) {real, imag} */,
  {32'h4565f57c, 32'h00000000} /* (3, 14, 26) {real, imag} */,
  {32'h4520dd58, 32'h00000000} /* (3, 14, 25) {real, imag} */,
  {32'h45403d22, 32'h00000000} /* (3, 14, 24) {real, imag} */,
  {32'h455c6614, 32'h00000000} /* (3, 14, 23) {real, imag} */,
  {32'h456d6e37, 32'h00000000} /* (3, 14, 22) {real, imag} */,
  {32'h45146531, 32'h00000000} /* (3, 14, 21) {real, imag} */,
  {32'hc4b11228, 32'h00000000} /* (3, 14, 20) {real, imag} */,
  {32'hc51f888a, 32'h00000000} /* (3, 14, 19) {real, imag} */,
  {32'hc568bbb5, 32'h00000000} /* (3, 14, 18) {real, imag} */,
  {32'hc5377389, 32'h00000000} /* (3, 14, 17) {real, imag} */,
  {32'hc57e3da2, 32'h00000000} /* (3, 14, 16) {real, imag} */,
  {32'hc55b0322, 32'h00000000} /* (3, 14, 15) {real, imag} */,
  {32'hc5094edc, 32'h00000000} /* (3, 14, 14) {real, imag} */,
  {32'hc53018f0, 32'h00000000} /* (3, 14, 13) {real, imag} */,
  {32'hc514fcf7, 32'h00000000} /* (3, 14, 12) {real, imag} */,
  {32'hc497d066, 32'h00000000} /* (3, 14, 11) {real, imag} */,
  {32'h4445aa6e, 32'h00000000} /* (3, 14, 10) {real, imag} */,
  {32'h4514a180, 32'h00000000} /* (3, 14, 9) {real, imag} */,
  {32'h454da1fe, 32'h00000000} /* (3, 14, 8) {real, imag} */,
  {32'h45202c28, 32'h00000000} /* (3, 14, 7) {real, imag} */,
  {32'h453e9f23, 32'h00000000} /* (3, 14, 6) {real, imag} */,
  {32'h453b22af, 32'h00000000} /* (3, 14, 5) {real, imag} */,
  {32'h452ed91c, 32'h00000000} /* (3, 14, 4) {real, imag} */,
  {32'h4545122a, 32'h00000000} /* (3, 14, 3) {real, imag} */,
  {32'h4555a715, 32'h00000000} /* (3, 14, 2) {real, imag} */,
  {32'h455c7c01, 32'h00000000} /* (3, 14, 1) {real, imag} */,
  {32'h45605954, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'h453e4630, 32'h00000000} /* (3, 13, 31) {real, imag} */,
  {32'h4572ce12, 32'h00000000} /* (3, 13, 30) {real, imag} */,
  {32'h45840d69, 32'h00000000} /* (3, 13, 29) {real, imag} */,
  {32'h458f840e, 32'h00000000} /* (3, 13, 28) {real, imag} */,
  {32'h4526da26, 32'h00000000} /* (3, 13, 27) {real, imag} */,
  {32'h4550169a, 32'h00000000} /* (3, 13, 26) {real, imag} */,
  {32'h455f535c, 32'h00000000} /* (3, 13, 25) {real, imag} */,
  {32'h453d4457, 32'h00000000} /* (3, 13, 24) {real, imag} */,
  {32'h455878f0, 32'h00000000} /* (3, 13, 23) {real, imag} */,
  {32'h45398251, 32'h00000000} /* (3, 13, 22) {real, imag} */,
  {32'h44acd66e, 32'h00000000} /* (3, 13, 21) {real, imag} */,
  {32'hc494e620, 32'h00000000} /* (3, 13, 20) {real, imag} */,
  {32'hc548a583, 32'h00000000} /* (3, 13, 19) {real, imag} */,
  {32'hc4fd6b26, 32'h00000000} /* (3, 13, 18) {real, imag} */,
  {32'hc57a7368, 32'h00000000} /* (3, 13, 17) {real, imag} */,
  {32'hc56b21dd, 32'h00000000} /* (3, 13, 16) {real, imag} */,
  {32'hc5213614, 32'h00000000} /* (3, 13, 15) {real, imag} */,
  {32'hc53da8a0, 32'h00000000} /* (3, 13, 14) {real, imag} */,
  {32'hc523308e, 32'h00000000} /* (3, 13, 13) {real, imag} */,
  {32'hc50fe6cb, 32'h00000000} /* (3, 13, 12) {real, imag} */,
  {32'hc4a3d52b, 32'h00000000} /* (3, 13, 11) {real, imag} */,
  {32'h4417080e, 32'h00000000} /* (3, 13, 10) {real, imag} */,
  {32'h44cb65c0, 32'h00000000} /* (3, 13, 9) {real, imag} */,
  {32'h451237a5, 32'h00000000} /* (3, 13, 8) {real, imag} */,
  {32'h453ff8f8, 32'h00000000} /* (3, 13, 7) {real, imag} */,
  {32'h450f2e71, 32'h00000000} /* (3, 13, 6) {real, imag} */,
  {32'h45273869, 32'h00000000} /* (3, 13, 5) {real, imag} */,
  {32'h45084040, 32'h00000000} /* (3, 13, 4) {real, imag} */,
  {32'h4525f57f, 32'h00000000} /* (3, 13, 3) {real, imag} */,
  {32'h4556d135, 32'h00000000} /* (3, 13, 2) {real, imag} */,
  {32'h4592336c, 32'h00000000} /* (3, 13, 1) {real, imag} */,
  {32'h453b90d9, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'h4509d7e8, 32'h00000000} /* (3, 12, 31) {real, imag} */,
  {32'h454e7a7a, 32'h00000000} /* (3, 12, 30) {real, imag} */,
  {32'h456f1bf5, 32'h00000000} /* (3, 12, 29) {real, imag} */,
  {32'h455b04e7, 32'h00000000} /* (3, 12, 28) {real, imag} */,
  {32'h4533da41, 32'h00000000} /* (3, 12, 27) {real, imag} */,
  {32'h4508f014, 32'h00000000} /* (3, 12, 26) {real, imag} */,
  {32'h45305695, 32'h00000000} /* (3, 12, 25) {real, imag} */,
  {32'h455ac882, 32'h00000000} /* (3, 12, 24) {real, imag} */,
  {32'h450ff832, 32'h00000000} /* (3, 12, 23) {real, imag} */,
  {32'h45193054, 32'h00000000} /* (3, 12, 22) {real, imag} */,
  {32'h440f05f1, 32'h00000000} /* (3, 12, 21) {real, imag} */,
  {32'hc4b56412, 32'h00000000} /* (3, 12, 20) {real, imag} */,
  {32'hc4a6e701, 32'h00000000} /* (3, 12, 19) {real, imag} */,
  {32'hc521ad35, 32'h00000000} /* (3, 12, 18) {real, imag} */,
  {32'hc524e4a1, 32'h00000000} /* (3, 12, 17) {real, imag} */,
  {32'hc54dfa2c, 32'h00000000} /* (3, 12, 16) {real, imag} */,
  {32'hc52af1f4, 32'h00000000} /* (3, 12, 15) {real, imag} */,
  {32'hc52c94e6, 32'h00000000} /* (3, 12, 14) {real, imag} */,
  {32'hc517da73, 32'h00000000} /* (3, 12, 13) {real, imag} */,
  {32'hc4942236, 32'h00000000} /* (3, 12, 12) {real, imag} */,
  {32'hc4574788, 32'h00000000} /* (3, 12, 11) {real, imag} */,
  {32'h4401b500, 32'h00000000} /* (3, 12, 10) {real, imag} */,
  {32'h44a69216, 32'h00000000} /* (3, 12, 9) {real, imag} */,
  {32'h44e44dcb, 32'h00000000} /* (3, 12, 8) {real, imag} */,
  {32'h452968ba, 32'h00000000} /* (3, 12, 7) {real, imag} */,
  {32'h45353bb8, 32'h00000000} /* (3, 12, 6) {real, imag} */,
  {32'h44eb2e1c, 32'h00000000} /* (3, 12, 5) {real, imag} */,
  {32'h44e29652, 32'h00000000} /* (3, 12, 4) {real, imag} */,
  {32'h45221cba, 32'h00000000} /* (3, 12, 3) {real, imag} */,
  {32'h450c99c9, 32'h00000000} /* (3, 12, 2) {real, imag} */,
  {32'h4590ecef, 32'h00000000} /* (3, 12, 1) {real, imag} */,
  {32'h453313e0, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'h44c401c2, 32'h00000000} /* (3, 11, 31) {real, imag} */,
  {32'h45179a9f, 32'h00000000} /* (3, 11, 30) {real, imag} */,
  {32'h451bbeac, 32'h00000000} /* (3, 11, 29) {real, imag} */,
  {32'h44eb25b6, 32'h00000000} /* (3, 11, 28) {real, imag} */,
  {32'h4514a600, 32'h00000000} /* (3, 11, 27) {real, imag} */,
  {32'h44bb24f4, 32'h00000000} /* (3, 11, 26) {real, imag} */,
  {32'h4481aecc, 32'h00000000} /* (3, 11, 25) {real, imag} */,
  {32'h44fef7a5, 32'h00000000} /* (3, 11, 24) {real, imag} */,
  {32'h44a64c96, 32'h00000000} /* (3, 11, 23) {real, imag} */,
  {32'h4489ea76, 32'h00000000} /* (3, 11, 22) {real, imag} */,
  {32'h44600f87, 32'h00000000} /* (3, 11, 21) {real, imag} */,
  {32'hc4651f0e, 32'h00000000} /* (3, 11, 20) {real, imag} */,
  {32'hc528c201, 32'h00000000} /* (3, 11, 19) {real, imag} */,
  {32'hc505d6a4, 32'h00000000} /* (3, 11, 18) {real, imag} */,
  {32'hc4b46d98, 32'h00000000} /* (3, 11, 17) {real, imag} */,
  {32'hc4ecd555, 32'h00000000} /* (3, 11, 16) {real, imag} */,
  {32'hc503cc73, 32'h00000000} /* (3, 11, 15) {real, imag} */,
  {32'hc4bbd002, 32'h00000000} /* (3, 11, 14) {real, imag} */,
  {32'hc4b0fb01, 32'h00000000} /* (3, 11, 13) {real, imag} */,
  {32'hc4adf8e0, 32'h00000000} /* (3, 11, 12) {real, imag} */,
  {32'hc451f3e7, 32'h00000000} /* (3, 11, 11) {real, imag} */,
  {32'h445324a7, 32'h00000000} /* (3, 11, 10) {real, imag} */,
  {32'h45015772, 32'h00000000} /* (3, 11, 9) {real, imag} */,
  {32'h44e3b223, 32'h00000000} /* (3, 11, 8) {real, imag} */,
  {32'h44fc44be, 32'h00000000} /* (3, 11, 7) {real, imag} */,
  {32'h44c8e91e, 32'h00000000} /* (3, 11, 6) {real, imag} */,
  {32'h44a4b726, 32'h00000000} /* (3, 11, 5) {real, imag} */,
  {32'h44d3afe5, 32'h00000000} /* (3, 11, 4) {real, imag} */,
  {32'h44eb1e0e, 32'h00000000} /* (3, 11, 3) {real, imag} */,
  {32'h44c58e97, 32'h00000000} /* (3, 11, 2) {real, imag} */,
  {32'h44ca444c, 32'h00000000} /* (3, 11, 1) {real, imag} */,
  {32'h44cb3d51, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'h4335702b, 32'h00000000} /* (3, 10, 31) {real, imag} */,
  {32'hc2e727ab, 32'h00000000} /* (3, 10, 30) {real, imag} */,
  {32'h435feb1a, 32'h00000000} /* (3, 10, 29) {real, imag} */,
  {32'h430475e7, 32'h00000000} /* (3, 10, 28) {real, imag} */,
  {32'hc2de7388, 32'h00000000} /* (3, 10, 27) {real, imag} */,
  {32'hc479b26d, 32'h00000000} /* (3, 10, 26) {real, imag} */,
  {32'h4178a9b0, 32'h00000000} /* (3, 10, 25) {real, imag} */,
  {32'hc4b8e0e2, 32'h00000000} /* (3, 10, 24) {real, imag} */,
  {32'hc3dc2938, 32'h00000000} /* (3, 10, 23) {real, imag} */,
  {32'hc41d7368, 32'h00000000} /* (3, 10, 22) {real, imag} */,
  {32'hc2b2a1ac, 32'h00000000} /* (3, 10, 21) {real, imag} */,
  {32'h43842743, 32'h00000000} /* (3, 10, 20) {real, imag} */,
  {32'hc305bbbc, 32'h00000000} /* (3, 10, 19) {real, imag} */,
  {32'h44311c55, 32'h00000000} /* (3, 10, 18) {real, imag} */,
  {32'h43a07b87, 32'h00000000} /* (3, 10, 17) {real, imag} */,
  {32'h44931df6, 32'h00000000} /* (3, 10, 16) {real, imag} */,
  {32'hc382e160, 32'h00000000} /* (3, 10, 15) {real, imag} */,
  {32'h42c094cb, 32'h00000000} /* (3, 10, 14) {real, imag} */,
  {32'hc2b50a74, 32'h00000000} /* (3, 10, 13) {real, imag} */,
  {32'h437d6709, 32'h00000000} /* (3, 10, 12) {real, imag} */,
  {32'h4470b81f, 32'h00000000} /* (3, 10, 11) {real, imag} */,
  {32'h4412c54f, 32'h00000000} /* (3, 10, 10) {real, imag} */,
  {32'h43654dd5, 32'h00000000} /* (3, 10, 9) {real, imag} */,
  {32'hc36cac84, 32'h00000000} /* (3, 10, 8) {real, imag} */,
  {32'h428adb2e, 32'h00000000} /* (3, 10, 7) {real, imag} */,
  {32'hc3a81645, 32'h00000000} /* (3, 10, 6) {real, imag} */,
  {32'hc40fbbc4, 32'h00000000} /* (3, 10, 5) {real, imag} */,
  {32'hc3f6924b, 32'h00000000} /* (3, 10, 4) {real, imag} */,
  {32'hc48d050e, 32'h00000000} /* (3, 10, 3) {real, imag} */,
  {32'hc4329bc1, 32'h00000000} /* (3, 10, 2) {real, imag} */,
  {32'hc1bc97f0, 32'h00000000} /* (3, 10, 1) {real, imag} */,
  {32'hc407c001, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'hc47b53e9, 32'h00000000} /* (3, 9, 31) {real, imag} */,
  {32'hc4ffac48, 32'h00000000} /* (3, 9, 30) {real, imag} */,
  {32'hc4a3cbf0, 32'h00000000} /* (3, 9, 29) {real, imag} */,
  {32'hc4cd2ea8, 32'h00000000} /* (3, 9, 28) {real, imag} */,
  {32'hc4c73a23, 32'h00000000} /* (3, 9, 27) {real, imag} */,
  {32'hc4e59f54, 32'h00000000} /* (3, 9, 26) {real, imag} */,
  {32'hc492919a, 32'h00000000} /* (3, 9, 25) {real, imag} */,
  {32'hc4921ed3, 32'h00000000} /* (3, 9, 24) {real, imag} */,
  {32'hc4d7f119, 32'h00000000} /* (3, 9, 23) {real, imag} */,
  {32'hc4d535e0, 32'h00000000} /* (3, 9, 22) {real, imag} */,
  {32'hc38e7b12, 32'h00000000} /* (3, 9, 21) {real, imag} */,
  {32'h4408ca1f, 32'h00000000} /* (3, 9, 20) {real, imag} */,
  {32'h44e90f72, 32'h00000000} /* (3, 9, 19) {real, imag} */,
  {32'h44dc8316, 32'h00000000} /* (3, 9, 18) {real, imag} */,
  {32'h4522aefa, 32'h00000000} /* (3, 9, 17) {real, imag} */,
  {32'h450d9516, 32'h00000000} /* (3, 9, 16) {real, imag} */,
  {32'h44ce4f48, 32'h00000000} /* (3, 9, 15) {real, imag} */,
  {32'h44ff766a, 32'h00000000} /* (3, 9, 14) {real, imag} */,
  {32'h44830bbc, 32'h00000000} /* (3, 9, 13) {real, imag} */,
  {32'h455023ee, 32'h00000000} /* (3, 9, 12) {real, imag} */,
  {32'h44d6ecd1, 32'h00000000} /* (3, 9, 11) {real, imag} */,
  {32'hc34a69ac, 32'h00000000} /* (3, 9, 10) {real, imag} */,
  {32'hc4a3ea50, 32'h00000000} /* (3, 9, 9) {real, imag} */,
  {32'hc4c8f197, 32'h00000000} /* (3, 9, 8) {real, imag} */,
  {32'hc453f64e, 32'h00000000} /* (3, 9, 7) {real, imag} */,
  {32'hc5016f98, 32'h00000000} /* (3, 9, 6) {real, imag} */,
  {32'hc4dcbb0c, 32'h00000000} /* (3, 9, 5) {real, imag} */,
  {32'hc50ec59c, 32'h00000000} /* (3, 9, 4) {real, imag} */,
  {32'hc52632dd, 32'h00000000} /* (3, 9, 3) {real, imag} */,
  {32'hc4d4e806, 32'h00000000} /* (3, 9, 2) {real, imag} */,
  {32'hc4e1ac1b, 32'h00000000} /* (3, 9, 1) {real, imag} */,
  {32'hc44d6e4e, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'hc491fed6, 32'h00000000} /* (3, 8, 31) {real, imag} */,
  {32'hc4d84536, 32'h00000000} /* (3, 8, 30) {real, imag} */,
  {32'hc502ab19, 32'h00000000} /* (3, 8, 29) {real, imag} */,
  {32'hc51ef64a, 32'h00000000} /* (3, 8, 28) {real, imag} */,
  {32'hc53bcd98, 32'h00000000} /* (3, 8, 27) {real, imag} */,
  {32'hc5456dff, 32'h00000000} /* (3, 8, 26) {real, imag} */,
  {32'hc5107b58, 32'h00000000} /* (3, 8, 25) {real, imag} */,
  {32'hc4fc751c, 32'h00000000} /* (3, 8, 24) {real, imag} */,
  {32'hc4fea843, 32'h00000000} /* (3, 8, 23) {real, imag} */,
  {32'hc4606fd4, 32'h00000000} /* (3, 8, 22) {real, imag} */,
  {32'h4378bcf0, 32'h00000000} /* (3, 8, 21) {real, imag} */,
  {32'h4498c3d8, 32'h00000000} /* (3, 8, 20) {real, imag} */,
  {32'h45256311, 32'h00000000} /* (3, 8, 19) {real, imag} */,
  {32'h454b85ec, 32'h00000000} /* (3, 8, 18) {real, imag} */,
  {32'h45099f93, 32'h00000000} /* (3, 8, 17) {real, imag} */,
  {32'h44ead742, 32'h00000000} /* (3, 8, 16) {real, imag} */,
  {32'h4547b847, 32'h00000000} /* (3, 8, 15) {real, imag} */,
  {32'h45059b62, 32'h00000000} /* (3, 8, 14) {real, imag} */,
  {32'h44be1128, 32'h00000000} /* (3, 8, 13) {real, imag} */,
  {32'h453ee89e, 32'h00000000} /* (3, 8, 12) {real, imag} */,
  {32'h448fa283, 32'h00000000} /* (3, 8, 11) {real, imag} */,
  {32'hc4eaa092, 32'h00000000} /* (3, 8, 10) {real, imag} */,
  {32'hc50225e2, 32'h00000000} /* (3, 8, 9) {real, imag} */,
  {32'hc526ad80, 32'h00000000} /* (3, 8, 8) {real, imag} */,
  {32'hc4de6fc5, 32'h00000000} /* (3, 8, 7) {real, imag} */,
  {32'hc5102adc, 32'h00000000} /* (3, 8, 6) {real, imag} */,
  {32'hc50df412, 32'h00000000} /* (3, 8, 5) {real, imag} */,
  {32'hc5141abf, 32'h00000000} /* (3, 8, 4) {real, imag} */,
  {32'hc53e2d07, 32'h00000000} /* (3, 8, 3) {real, imag} */,
  {32'hc4f8fe97, 32'h00000000} /* (3, 8, 2) {real, imag} */,
  {32'hc506e111, 32'h00000000} /* (3, 8, 1) {real, imag} */,
  {32'hc4b347d2, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'hc4c1e8d4, 32'h00000000} /* (3, 7, 31) {real, imag} */,
  {32'hc4c4cd74, 32'h00000000} /* (3, 7, 30) {real, imag} */,
  {32'hc52aa326, 32'h00000000} /* (3, 7, 29) {real, imag} */,
  {32'hc5879a4a, 32'h00000000} /* (3, 7, 28) {real, imag} */,
  {32'hc5654d80, 32'h00000000} /* (3, 7, 27) {real, imag} */,
  {32'hc591a6b8, 32'h00000000} /* (3, 7, 26) {real, imag} */,
  {32'hc52f5c3b, 32'h00000000} /* (3, 7, 25) {real, imag} */,
  {32'hc51b5ca0, 32'h00000000} /* (3, 7, 24) {real, imag} */,
  {32'hc500c773, 32'h00000000} /* (3, 7, 23) {real, imag} */,
  {32'hc467c71f, 32'h00000000} /* (3, 7, 22) {real, imag} */,
  {32'hc32b1818, 32'h00000000} /* (3, 7, 21) {real, imag} */,
  {32'h44d4c240, 32'h00000000} /* (3, 7, 20) {real, imag} */,
  {32'h450ce84b, 32'h00000000} /* (3, 7, 19) {real, imag} */,
  {32'h45145c48, 32'h00000000} /* (3, 7, 18) {real, imag} */,
  {32'h4572f1c9, 32'h00000000} /* (3, 7, 17) {real, imag} */,
  {32'h45445960, 32'h00000000} /* (3, 7, 16) {real, imag} */,
  {32'h450ebe6a, 32'h00000000} /* (3, 7, 15) {real, imag} */,
  {32'h4544b72a, 32'h00000000} /* (3, 7, 14) {real, imag} */,
  {32'h450927e8, 32'h00000000} /* (3, 7, 13) {real, imag} */,
  {32'h4517590e, 32'h00000000} /* (3, 7, 12) {real, imag} */,
  {32'h449d161b, 32'h00000000} /* (3, 7, 11) {real, imag} */,
  {32'hc4689364, 32'h00000000} /* (3, 7, 10) {real, imag} */,
  {32'hc5077bf3, 32'h00000000} /* (3, 7, 9) {real, imag} */,
  {32'hc4a32e82, 32'h00000000} /* (3, 7, 8) {real, imag} */,
  {32'hc4f6fade, 32'h00000000} /* (3, 7, 7) {real, imag} */,
  {32'hc4a7bb18, 32'h00000000} /* (3, 7, 6) {real, imag} */,
  {32'hc51833be, 32'h00000000} /* (3, 7, 5) {real, imag} */,
  {32'hc523d8da, 32'h00000000} /* (3, 7, 4) {real, imag} */,
  {32'hc5684da9, 32'h00000000} /* (3, 7, 3) {real, imag} */,
  {32'hc5029eee, 32'h00000000} /* (3, 7, 2) {real, imag} */,
  {32'hc4cb4b06, 32'h00000000} /* (3, 7, 1) {real, imag} */,
  {32'hc4a77477, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'hc48d618f, 32'h00000000} /* (3, 6, 31) {real, imag} */,
  {32'hc5130aec, 32'h00000000} /* (3, 6, 30) {real, imag} */,
  {32'hc531d158, 32'h00000000} /* (3, 6, 29) {real, imag} */,
  {32'hc54f3713, 32'h00000000} /* (3, 6, 28) {real, imag} */,
  {32'hc5802f74, 32'h00000000} /* (3, 6, 27) {real, imag} */,
  {32'hc561dc02, 32'h00000000} /* (3, 6, 26) {real, imag} */,
  {32'hc5638f10, 32'h00000000} /* (3, 6, 25) {real, imag} */,
  {32'hc5301a8f, 32'h00000000} /* (3, 6, 24) {real, imag} */,
  {32'hc50210fe, 32'h00000000} /* (3, 6, 23) {real, imag} */,
  {32'hc49c2e40, 32'h00000000} /* (3, 6, 22) {real, imag} */,
  {32'hc3003e3c, 32'h00000000} /* (3, 6, 21) {real, imag} */,
  {32'h446dc9ee, 32'h00000000} /* (3, 6, 20) {real, imag} */,
  {32'h44ac3611, 32'h00000000} /* (3, 6, 19) {real, imag} */,
  {32'h44b3a924, 32'h00000000} /* (3, 6, 18) {real, imag} */,
  {32'h4505c552, 32'h00000000} /* (3, 6, 17) {real, imag} */,
  {32'h450f1c1a, 32'h00000000} /* (3, 6, 16) {real, imag} */,
  {32'h4532645a, 32'h00000000} /* (3, 6, 15) {real, imag} */,
  {32'h45525836, 32'h00000000} /* (3, 6, 14) {real, imag} */,
  {32'h451ede58, 32'h00000000} /* (3, 6, 13) {real, imag} */,
  {32'h4503ab0f, 32'h00000000} /* (3, 6, 12) {real, imag} */,
  {32'h45211347, 32'h00000000} /* (3, 6, 11) {real, imag} */,
  {32'hc2e2b580, 32'h00000000} /* (3, 6, 10) {real, imag} */,
  {32'hc3d02518, 32'h00000000} /* (3, 6, 9) {real, imag} */,
  {32'hc3947158, 32'h00000000} /* (3, 6, 8) {real, imag} */,
  {32'hc43124e8, 32'h00000000} /* (3, 6, 7) {real, imag} */,
  {32'hc5049e93, 32'h00000000} /* (3, 6, 6) {real, imag} */,
  {32'hc4ee2f86, 32'h00000000} /* (3, 6, 5) {real, imag} */,
  {32'hc4c190cf, 32'h00000000} /* (3, 6, 4) {real, imag} */,
  {32'hc50167fe, 32'h00000000} /* (3, 6, 3) {real, imag} */,
  {32'hc53dd474, 32'h00000000} /* (3, 6, 2) {real, imag} */,
  {32'hc517499e, 32'h00000000} /* (3, 6, 1) {real, imag} */,
  {32'hc4c09ac2, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hc4b8e679, 32'h00000000} /* (3, 5, 31) {real, imag} */,
  {32'hc50f6c94, 32'h00000000} /* (3, 5, 30) {real, imag} */,
  {32'hc539edbc, 32'h00000000} /* (3, 5, 29) {real, imag} */,
  {32'hc54a9e8c, 32'h00000000} /* (3, 5, 28) {real, imag} */,
  {32'hc558a5bc, 32'h00000000} /* (3, 5, 27) {real, imag} */,
  {32'hc56783b1, 32'h00000000} /* (3, 5, 26) {real, imag} */,
  {32'hc56769fc, 32'h00000000} /* (3, 5, 25) {real, imag} */,
  {32'hc575a242, 32'h00000000} /* (3, 5, 24) {real, imag} */,
  {32'hc4fe65a6, 32'h00000000} /* (3, 5, 23) {real, imag} */,
  {32'hc483cf92, 32'h00000000} /* (3, 5, 22) {real, imag} */,
  {32'hc414d7f2, 32'h00000000} /* (3, 5, 21) {real, imag} */,
  {32'hc46b35be, 32'h00000000} /* (3, 5, 20) {real, imag} */,
  {32'h42dfff80, 32'h00000000} /* (3, 5, 19) {real, imag} */,
  {32'h4357a4e8, 32'h00000000} /* (3, 5, 18) {real, imag} */,
  {32'hc229e580, 32'h00000000} /* (3, 5, 17) {real, imag} */,
  {32'h4475f0ba, 32'h00000000} /* (3, 5, 16) {real, imag} */,
  {32'h44de0def, 32'h00000000} /* (3, 5, 15) {real, imag} */,
  {32'h452b2e32, 32'h00000000} /* (3, 5, 14) {real, imag} */,
  {32'h45477b4c, 32'h00000000} /* (3, 5, 13) {real, imag} */,
  {32'h455788e4, 32'h00000000} /* (3, 5, 12) {real, imag} */,
  {32'h45249b9c, 32'h00000000} /* (3, 5, 11) {real, imag} */,
  {32'h4548ff79, 32'h00000000} /* (3, 5, 10) {real, imag} */,
  {32'h44872165, 32'h00000000} /* (3, 5, 9) {real, imag} */,
  {32'h445bd4f6, 32'h00000000} /* (3, 5, 8) {real, imag} */,
  {32'h4468a078, 32'h00000000} /* (3, 5, 7) {real, imag} */,
  {32'hc311f634, 32'h00000000} /* (3, 5, 6) {real, imag} */,
  {32'hc40a020a, 32'h00000000} /* (3, 5, 5) {real, imag} */,
  {32'hc4a2a475, 32'h00000000} /* (3, 5, 4) {real, imag} */,
  {32'hc4ca12e6, 32'h00000000} /* (3, 5, 3) {real, imag} */,
  {32'hc5015350, 32'h00000000} /* (3, 5, 2) {real, imag} */,
  {32'hc4d0f1fa, 32'h00000000} /* (3, 5, 1) {real, imag} */,
  {32'hc4bffee7, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hc502d5f7, 32'h00000000} /* (3, 4, 31) {real, imag} */,
  {32'hc52c57d9, 32'h00000000} /* (3, 4, 30) {real, imag} */,
  {32'hc5524ec3, 32'h00000000} /* (3, 4, 29) {real, imag} */,
  {32'hc56dbb25, 32'h00000000} /* (3, 4, 28) {real, imag} */,
  {32'hc5793d86, 32'h00000000} /* (3, 4, 27) {real, imag} */,
  {32'hc56cf9b6, 32'h00000000} /* (3, 4, 26) {real, imag} */,
  {32'hc53f233d, 32'h00000000} /* (3, 4, 25) {real, imag} */,
  {32'hc5257cee, 32'h00000000} /* (3, 4, 24) {real, imag} */,
  {32'hc535a9db, 32'h00000000} /* (3, 4, 23) {real, imag} */,
  {32'hc4fe2507, 32'h00000000} /* (3, 4, 22) {real, imag} */,
  {32'hc4699e07, 32'h00000000} /* (3, 4, 21) {real, imag} */,
  {32'hc4abb4f8, 32'h00000000} /* (3, 4, 20) {real, imag} */,
  {32'hc4f77106, 32'h00000000} /* (3, 4, 19) {real, imag} */,
  {32'hc487bc99, 32'h00000000} /* (3, 4, 18) {real, imag} */,
  {32'hc4716fd8, 32'h00000000} /* (3, 4, 17) {real, imag} */,
  {32'h44038cf8, 32'h00000000} /* (3, 4, 16) {real, imag} */,
  {32'h4504eae9, 32'h00000000} /* (3, 4, 15) {real, imag} */,
  {32'h452b089f, 32'h00000000} /* (3, 4, 14) {real, imag} */,
  {32'h45743329, 32'h00000000} /* (3, 4, 13) {real, imag} */,
  {32'h4575d807, 32'h00000000} /* (3, 4, 12) {real, imag} */,
  {32'h454e9252, 32'h00000000} /* (3, 4, 11) {real, imag} */,
  {32'h4563b3a6, 32'h00000000} /* (3, 4, 10) {real, imag} */,
  {32'h45342e6d, 32'h00000000} /* (3, 4, 9) {real, imag} */,
  {32'h45394a0e, 32'h00000000} /* (3, 4, 8) {real, imag} */,
  {32'h4514fa8f, 32'h00000000} /* (3, 4, 7) {real, imag} */,
  {32'h450e900b, 32'h00000000} /* (3, 4, 6) {real, imag} */,
  {32'h440bf109, 32'h00000000} /* (3, 4, 5) {real, imag} */,
  {32'hc426920b, 32'h00000000} /* (3, 4, 4) {real, imag} */,
  {32'hc4a4798e, 32'h00000000} /* (3, 4, 3) {real, imag} */,
  {32'hc4c1063f, 32'h00000000} /* (3, 4, 2) {real, imag} */,
  {32'hc4ce5048, 32'h00000000} /* (3, 4, 1) {real, imag} */,
  {32'hc4856456, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hc4ac4d6c, 32'h00000000} /* (3, 3, 31) {real, imag} */,
  {32'hc5376400, 32'h00000000} /* (3, 3, 30) {real, imag} */,
  {32'hc5771ec4, 32'h00000000} /* (3, 3, 29) {real, imag} */,
  {32'hc53f74a4, 32'h00000000} /* (3, 3, 28) {real, imag} */,
  {32'hc54b2f03, 32'h00000000} /* (3, 3, 27) {real, imag} */,
  {32'hc53e27d4, 32'h00000000} /* (3, 3, 26) {real, imag} */,
  {32'hc53bbc52, 32'h00000000} /* (3, 3, 25) {real, imag} */,
  {32'hc53d8c19, 32'h00000000} /* (3, 3, 24) {real, imag} */,
  {32'hc5197c02, 32'h00000000} /* (3, 3, 23) {real, imag} */,
  {32'hc50d878e, 32'h00000000} /* (3, 3, 22) {real, imag} */,
  {32'hc500fc24, 32'h00000000} /* (3, 3, 21) {real, imag} */,
  {32'hc51131d4, 32'h00000000} /* (3, 3, 20) {real, imag} */,
  {32'hc502586b, 32'h00000000} /* (3, 3, 19) {real, imag} */,
  {32'hc5115cd8, 32'h00000000} /* (3, 3, 18) {real, imag} */,
  {32'hc4a65471, 32'h00000000} /* (3, 3, 17) {real, imag} */,
  {32'hc485cd7c, 32'h00000000} /* (3, 3, 16) {real, imag} */,
  {32'h44cc4920, 32'h00000000} /* (3, 3, 15) {real, imag} */,
  {32'h45296db2, 32'h00000000} /* (3, 3, 14) {real, imag} */,
  {32'h457521de, 32'h00000000} /* (3, 3, 13) {real, imag} */,
  {32'h4586ef8c, 32'h00000000} /* (3, 3, 12) {real, imag} */,
  {32'h4568de15, 32'h00000000} /* (3, 3, 11) {real, imag} */,
  {32'h45820162, 32'h00000000} /* (3, 3, 10) {real, imag} */,
  {32'h4542a3c2, 32'h00000000} /* (3, 3, 9) {real, imag} */,
  {32'h455182a9, 32'h00000000} /* (3, 3, 8) {real, imag} */,
  {32'h451a6c6c, 32'h00000000} /* (3, 3, 7) {real, imag} */,
  {32'h4514289a, 32'h00000000} /* (3, 3, 6) {real, imag} */,
  {32'h43dceaa0, 32'h00000000} /* (3, 3, 5) {real, imag} */,
  {32'hc45b02d3, 32'h00000000} /* (3, 3, 4) {real, imag} */,
  {32'hc4fe4ae6, 32'h00000000} /* (3, 3, 3) {real, imag} */,
  {32'hc4e04248, 32'h00000000} /* (3, 3, 2) {real, imag} */,
  {32'hc5179a8e, 32'h00000000} /* (3, 3, 1) {real, imag} */,
  {32'hc4a44618, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hc4ae580d, 32'h00000000} /* (3, 2, 31) {real, imag} */,
  {32'hc513185c, 32'h00000000} /* (3, 2, 30) {real, imag} */,
  {32'hc5341439, 32'h00000000} /* (3, 2, 29) {real, imag} */,
  {32'hc51a9496, 32'h00000000} /* (3, 2, 28) {real, imag} */,
  {32'hc523a65a, 32'h00000000} /* (3, 2, 27) {real, imag} */,
  {32'hc50ae792, 32'h00000000} /* (3, 2, 26) {real, imag} */,
  {32'hc52e526f, 32'h00000000} /* (3, 2, 25) {real, imag} */,
  {32'hc4f2af55, 32'h00000000} /* (3, 2, 24) {real, imag} */,
  {32'hc4cd4968, 32'h00000000} /* (3, 2, 23) {real, imag} */,
  {32'hc4ecad9e, 32'h00000000} /* (3, 2, 22) {real, imag} */,
  {32'hc4f8c4cc, 32'h00000000} /* (3, 2, 21) {real, imag} */,
  {32'hc53d24c9, 32'h00000000} /* (3, 2, 20) {real, imag} */,
  {32'hc52171e0, 32'h00000000} /* (3, 2, 19) {real, imag} */,
  {32'hc506852e, 32'h00000000} /* (3, 2, 18) {real, imag} */,
  {32'hc4c9a92c, 32'h00000000} /* (3, 2, 17) {real, imag} */,
  {32'hc2903360, 32'h00000000} /* (3, 2, 16) {real, imag} */,
  {32'h44d936db, 32'h00000000} /* (3, 2, 15) {real, imag} */,
  {32'h455eb0c2, 32'h00000000} /* (3, 2, 14) {real, imag} */,
  {32'h453c4369, 32'h00000000} /* (3, 2, 13) {real, imag} */,
  {32'h455c8dfe, 32'h00000000} /* (3, 2, 12) {real, imag} */,
  {32'h457bcbb6, 32'h00000000} /* (3, 2, 11) {real, imag} */,
  {32'h457a3e9c, 32'h00000000} /* (3, 2, 10) {real, imag} */,
  {32'h45803a48, 32'h00000000} /* (3, 2, 9) {real, imag} */,
  {32'h45223844, 32'h00000000} /* (3, 2, 8) {real, imag} */,
  {32'h452f9622, 32'h00000000} /* (3, 2, 7) {real, imag} */,
  {32'h453315f9, 32'h00000000} /* (3, 2, 6) {real, imag} */,
  {32'h439cc1a2, 32'h00000000} /* (3, 2, 5) {real, imag} */,
  {32'hc4a66546, 32'h00000000} /* (3, 2, 4) {real, imag} */,
  {32'hc48e066b, 32'h00000000} /* (3, 2, 3) {real, imag} */,
  {32'hc4f263b4, 32'h00000000} /* (3, 2, 2) {real, imag} */,
  {32'hc4a60fc8, 32'h00000000} /* (3, 2, 1) {real, imag} */,
  {32'hc48d7768, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hc433f5fc, 32'h00000000} /* (3, 1, 31) {real, imag} */,
  {32'hc4bfcb68, 32'h00000000} /* (3, 1, 30) {real, imag} */,
  {32'hc4f61656, 32'h00000000} /* (3, 1, 29) {real, imag} */,
  {32'hc4d2c383, 32'h00000000} /* (3, 1, 28) {real, imag} */,
  {32'hc51111be, 32'h00000000} /* (3, 1, 27) {real, imag} */,
  {32'hc508f8e0, 32'h00000000} /* (3, 1, 26) {real, imag} */,
  {32'hc5059286, 32'h00000000} /* (3, 1, 25) {real, imag} */,
  {32'hc4c850bd, 32'h00000000} /* (3, 1, 24) {real, imag} */,
  {32'hc48c8b97, 32'h00000000} /* (3, 1, 23) {real, imag} */,
  {32'hc4bede0a, 32'h00000000} /* (3, 1, 22) {real, imag} */,
  {32'hc52076d2, 32'h00000000} /* (3, 1, 21) {real, imag} */,
  {32'hc4f1cee2, 32'h00000000} /* (3, 1, 20) {real, imag} */,
  {32'hc4da9767, 32'h00000000} /* (3, 1, 19) {real, imag} */,
  {32'hc49e3cf6, 32'h00000000} /* (3, 1, 18) {real, imag} */,
  {32'hc427ba94, 32'h00000000} /* (3, 1, 17) {real, imag} */,
  {32'hc2988b20, 32'h00000000} /* (3, 1, 16) {real, imag} */,
  {32'h44e845d8, 32'h00000000} /* (3, 1, 15) {real, imag} */,
  {32'h452060bc, 32'h00000000} /* (3, 1, 14) {real, imag} */,
  {32'h455509c5, 32'h00000000} /* (3, 1, 13) {real, imag} */,
  {32'h45630ba6, 32'h00000000} /* (3, 1, 12) {real, imag} */,
  {32'h456b638e, 32'h00000000} /* (3, 1, 11) {real, imag} */,
  {32'h458351d6, 32'h00000000} /* (3, 1, 10) {real, imag} */,
  {32'h45385472, 32'h00000000} /* (3, 1, 9) {real, imag} */,
  {32'h452ef812, 32'h00000000} /* (3, 1, 8) {real, imag} */,
  {32'h4566e14a, 32'h00000000} /* (3, 1, 7) {real, imag} */,
  {32'h4545af93, 32'h00000000} /* (3, 1, 6) {real, imag} */,
  {32'h4413f96e, 32'h00000000} /* (3, 1, 5) {real, imag} */,
  {32'hc465a6d8, 32'h00000000} /* (3, 1, 4) {real, imag} */,
  {32'hc4b5e7f7, 32'h00000000} /* (3, 1, 3) {real, imag} */,
  {32'hc4ccbb3e, 32'h00000000} /* (3, 1, 2) {real, imag} */,
  {32'hc510a0a8, 32'h00000000} /* (3, 1, 1) {real, imag} */,
  {32'hc46f1960, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'hc4048657, 32'h00000000} /* (3, 0, 31) {real, imag} */,
  {32'hc4512919, 32'h00000000} /* (3, 0, 30) {real, imag} */,
  {32'hc4bf02bd, 32'h00000000} /* (3, 0, 29) {real, imag} */,
  {32'hc4b0ca60, 32'h00000000} /* (3, 0, 28) {real, imag} */,
  {32'hc463b0f7, 32'h00000000} /* (3, 0, 27) {real, imag} */,
  {32'hc4bcaa79, 32'h00000000} /* (3, 0, 26) {real, imag} */,
  {32'hc4b57c2a, 32'h00000000} /* (3, 0, 25) {real, imag} */,
  {32'hc4b2034c, 32'h00000000} /* (3, 0, 24) {real, imag} */,
  {32'hc478f18f, 32'h00000000} /* (3, 0, 23) {real, imag} */,
  {32'hc46032e9, 32'h00000000} /* (3, 0, 22) {real, imag} */,
  {32'hc46eab5a, 32'h00000000} /* (3, 0, 21) {real, imag} */,
  {32'hc41cc741, 32'h00000000} /* (3, 0, 20) {real, imag} */,
  {32'hc4016be3, 32'h00000000} /* (3, 0, 19) {real, imag} */,
  {32'hc401f9ab, 32'h00000000} /* (3, 0, 18) {real, imag} */,
  {32'h40e00cc0, 32'h00000000} /* (3, 0, 17) {real, imag} */,
  {32'h44444a69, 32'h00000000} /* (3, 0, 16) {real, imag} */,
  {32'h44ecf3b0, 32'h00000000} /* (3, 0, 15) {real, imag} */,
  {32'h451e9ae8, 32'h00000000} /* (3, 0, 14) {real, imag} */,
  {32'h455f539c, 32'h00000000} /* (3, 0, 13) {real, imag} */,
  {32'h453939d4, 32'h00000000} /* (3, 0, 12) {real, imag} */,
  {32'h452780f8, 32'h00000000} /* (3, 0, 11) {real, imag} */,
  {32'h450a42f8, 32'h00000000} /* (3, 0, 10) {real, imag} */,
  {32'h45274a29, 32'h00000000} /* (3, 0, 9) {real, imag} */,
  {32'h450c5ebf, 32'h00000000} /* (3, 0, 8) {real, imag} */,
  {32'h44fb05e8, 32'h00000000} /* (3, 0, 7) {real, imag} */,
  {32'h4500b281, 32'h00000000} /* (3, 0, 6) {real, imag} */,
  {32'h438b7874, 32'h00000000} /* (3, 0, 5) {real, imag} */,
  {32'hc4077b11, 32'h00000000} /* (3, 0, 4) {real, imag} */,
  {32'hc4ebc19a, 32'h00000000} /* (3, 0, 3) {real, imag} */,
  {32'hc496eacc, 32'h00000000} /* (3, 0, 2) {real, imag} */,
  {32'hc4601cda, 32'h00000000} /* (3, 0, 1) {real, imag} */,
  {32'hc42ac80b, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc4958656, 32'h00000000} /* (2, 31, 31) {real, imag} */,
  {32'hc4cad067, 32'h00000000} /* (2, 31, 30) {real, imag} */,
  {32'hc4e6b186, 32'h00000000} /* (2, 31, 29) {real, imag} */,
  {32'hc50164ac, 32'h00000000} /* (2, 31, 28) {real, imag} */,
  {32'hc52f5152, 32'h00000000} /* (2, 31, 27) {real, imag} */,
  {32'hc50d3318, 32'h00000000} /* (2, 31, 26) {real, imag} */,
  {32'hc4f39402, 32'h00000000} /* (2, 31, 25) {real, imag} */,
  {32'hc502663c, 32'h00000000} /* (2, 31, 24) {real, imag} */,
  {32'hc4df7c4a, 32'h00000000} /* (2, 31, 23) {real, imag} */,
  {32'hc499c7c6, 32'h00000000} /* (2, 31, 22) {real, imag} */,
  {32'hc4a30fcc, 32'h00000000} /* (2, 31, 21) {real, imag} */,
  {32'h444231fa, 32'h00000000} /* (2, 31, 20) {real, imag} */,
  {32'h44950d10, 32'h00000000} /* (2, 31, 19) {real, imag} */,
  {32'h4470e738, 32'h00000000} /* (2, 31, 18) {real, imag} */,
  {32'h44d2b9aa, 32'h00000000} /* (2, 31, 17) {real, imag} */,
  {32'h45065e0a, 32'h00000000} /* (2, 31, 16) {real, imag} */,
  {32'h453fdba7, 32'h00000000} /* (2, 31, 15) {real, imag} */,
  {32'h454f9822, 32'h00000000} /* (2, 31, 14) {real, imag} */,
  {32'h45543367, 32'h00000000} /* (2, 31, 13) {real, imag} */,
  {32'h45170500, 32'h00000000} /* (2, 31, 12) {real, imag} */,
  {32'h45017286, 32'h00000000} /* (2, 31, 11) {real, imag} */,
  {32'h4458257e, 32'h00000000} /* (2, 31, 10) {real, imag} */,
  {32'hc4153ad8, 32'h00000000} /* (2, 31, 9) {real, imag} */,
  {32'hc39c779e, 32'h00000000} /* (2, 31, 8) {real, imag} */,
  {32'hc4a5b8b2, 32'h00000000} /* (2, 31, 7) {real, imag} */,
  {32'hc4e66860, 32'h00000000} /* (2, 31, 6) {real, imag} */,
  {32'hc4c93f64, 32'h00000000} /* (2, 31, 5) {real, imag} */,
  {32'hc4b5dc35, 32'h00000000} /* (2, 31, 4) {real, imag} */,
  {32'hc503a61e, 32'h00000000} /* (2, 31, 3) {real, imag} */,
  {32'hc51cd9eb, 32'h00000000} /* (2, 31, 2) {real, imag} */,
  {32'hc52394af, 32'h00000000} /* (2, 31, 1) {real, imag} */,
  {32'hc47c3cde, 32'h00000000} /* (2, 31, 0) {real, imag} */,
  {32'hc4a9b46c, 32'h00000000} /* (2, 30, 31) {real, imag} */,
  {32'hc50e37d5, 32'h00000000} /* (2, 30, 30) {real, imag} */,
  {32'hc4e2ed7e, 32'h00000000} /* (2, 30, 29) {real, imag} */,
  {32'hc557d3ad, 32'h00000000} /* (2, 30, 28) {real, imag} */,
  {32'hc53a3e72, 32'h00000000} /* (2, 30, 27) {real, imag} */,
  {32'hc5269333, 32'h00000000} /* (2, 30, 26) {real, imag} */,
  {32'hc53ebad8, 32'h00000000} /* (2, 30, 25) {real, imag} */,
  {32'hc501e1cb, 32'h00000000} /* (2, 30, 24) {real, imag} */,
  {32'hc4e17a2e, 32'h00000000} /* (2, 30, 23) {real, imag} */,
  {32'hc50ec8d4, 32'h00000000} /* (2, 30, 22) {real, imag} */,
  {32'hc40a8032, 32'h00000000} /* (2, 30, 21) {real, imag} */,
  {32'h4505033c, 32'h00000000} /* (2, 30, 20) {real, imag} */,
  {32'h4542c51f, 32'h00000000} /* (2, 30, 19) {real, imag} */,
  {32'h450129bf, 32'h00000000} /* (2, 30, 18) {real, imag} */,
  {32'h4549307c, 32'h00000000} /* (2, 30, 17) {real, imag} */,
  {32'h454c58c4, 32'h00000000} /* (2, 30, 16) {real, imag} */,
  {32'h4564e2e0, 32'h00000000} /* (2, 30, 15) {real, imag} */,
  {32'h4579c60d, 32'h00000000} /* (2, 30, 14) {real, imag} */,
  {32'h4556987f, 32'h00000000} /* (2, 30, 13) {real, imag} */,
  {32'h45395e3d, 32'h00000000} /* (2, 30, 12) {real, imag} */,
  {32'h44f8bc60, 32'h00000000} /* (2, 30, 11) {real, imag} */,
  {32'hc38cfc18, 32'h00000000} /* (2, 30, 10) {real, imag} */,
  {32'hc4a06110, 32'h00000000} /* (2, 30, 9) {real, imag} */,
  {32'hc4a8dc75, 32'h00000000} /* (2, 30, 8) {real, imag} */,
  {32'hc51008a9, 32'h00000000} /* (2, 30, 7) {real, imag} */,
  {32'hc51281ba, 32'h00000000} /* (2, 30, 6) {real, imag} */,
  {32'hc5189808, 32'h00000000} /* (2, 30, 5) {real, imag} */,
  {32'hc547b4c0, 32'h00000000} /* (2, 30, 4) {real, imag} */,
  {32'hc4ec07fe, 32'h00000000} /* (2, 30, 3) {real, imag} */,
  {32'hc5768889, 32'h00000000} /* (2, 30, 2) {real, imag} */,
  {32'hc4ec6fab, 32'h00000000} /* (2, 30, 1) {real, imag} */,
  {32'hc485f664, 32'h00000000} /* (2, 30, 0) {real, imag} */,
  {32'hc4cd9a6b, 32'h00000000} /* (2, 29, 31) {real, imag} */,
  {32'hc503c03e, 32'h00000000} /* (2, 29, 30) {real, imag} */,
  {32'hc5470d2e, 32'h00000000} /* (2, 29, 29) {real, imag} */,
  {32'hc544b4aa, 32'h00000000} /* (2, 29, 28) {real, imag} */,
  {32'hc5609a5a, 32'h00000000} /* (2, 29, 27) {real, imag} */,
  {32'hc5813d9c, 32'h00000000} /* (2, 29, 26) {real, imag} */,
  {32'hc54acd34, 32'h00000000} /* (2, 29, 25) {real, imag} */,
  {32'hc580970b, 32'h00000000} /* (2, 29, 24) {real, imag} */,
  {32'hc502e10d, 32'h00000000} /* (2, 29, 23) {real, imag} */,
  {32'hc5073ad2, 32'h00000000} /* (2, 29, 22) {real, imag} */,
  {32'hc3565560, 32'h00000000} /* (2, 29, 21) {real, imag} */,
  {32'h45276321, 32'h00000000} /* (2, 29, 20) {real, imag} */,
  {32'h458baa06, 32'h00000000} /* (2, 29, 19) {real, imag} */,
  {32'h458c649a, 32'h00000000} /* (2, 29, 18) {real, imag} */,
  {32'h45644d33, 32'h00000000} /* (2, 29, 17) {real, imag} */,
  {32'h458782b6, 32'h00000000} /* (2, 29, 16) {real, imag} */,
  {32'h4560a152, 32'h00000000} /* (2, 29, 15) {real, imag} */,
  {32'h454eed62, 32'h00000000} /* (2, 29, 14) {real, imag} */,
  {32'h455dab04, 32'h00000000} /* (2, 29, 13) {real, imag} */,
  {32'h4531e2e6, 32'h00000000} /* (2, 29, 12) {real, imag} */,
  {32'h44e39643, 32'h00000000} /* (2, 29, 11) {real, imag} */,
  {32'hc4264234, 32'h00000000} /* (2, 29, 10) {real, imag} */,
  {32'hc4c3b4e3, 32'h00000000} /* (2, 29, 9) {real, imag} */,
  {32'hc4c0b1fc, 32'h00000000} /* (2, 29, 8) {real, imag} */,
  {32'hc5000dc3, 32'h00000000} /* (2, 29, 7) {real, imag} */,
  {32'hc5317306, 32'h00000000} /* (2, 29, 6) {real, imag} */,
  {32'hc51aab2e, 32'h00000000} /* (2, 29, 5) {real, imag} */,
  {32'hc54a2033, 32'h00000000} /* (2, 29, 4) {real, imag} */,
  {32'hc53e9e7c, 32'h00000000} /* (2, 29, 3) {real, imag} */,
  {32'hc56055fb, 32'h00000000} /* (2, 29, 2) {real, imag} */,
  {32'hc4db0fb6, 32'h00000000} /* (2, 29, 1) {real, imag} */,
  {32'hc492f808, 32'h00000000} /* (2, 29, 0) {real, imag} */,
  {32'hc5126674, 32'h00000000} /* (2, 28, 31) {real, imag} */,
  {32'hc5294757, 32'h00000000} /* (2, 28, 30) {real, imag} */,
  {32'hc5435a24, 32'h00000000} /* (2, 28, 29) {real, imag} */,
  {32'hc5776da7, 32'h00000000} /* (2, 28, 28) {real, imag} */,
  {32'hc57088c3, 32'h00000000} /* (2, 28, 27) {real, imag} */,
  {32'hc57e219e, 32'h00000000} /* (2, 28, 26) {real, imag} */,
  {32'hc5404a4e, 32'h00000000} /* (2, 28, 25) {real, imag} */,
  {32'hc5334fd5, 32'h00000000} /* (2, 28, 24) {real, imag} */,
  {32'hc53bed2f, 32'h00000000} /* (2, 28, 23) {real, imag} */,
  {32'hc537886a, 32'h00000000} /* (2, 28, 22) {real, imag} */,
  {32'h42ef09a0, 32'h00000000} /* (2, 28, 21) {real, imag} */,
  {32'h455cfa58, 32'h00000000} /* (2, 28, 20) {real, imag} */,
  {32'h458fd0c4, 32'h00000000} /* (2, 28, 19) {real, imag} */,
  {32'h4599f173, 32'h00000000} /* (2, 28, 18) {real, imag} */,
  {32'h45954e84, 32'h00000000} /* (2, 28, 17) {real, imag} */,
  {32'h459c9e0b, 32'h00000000} /* (2, 28, 16) {real, imag} */,
  {32'h4564008e, 32'h00000000} /* (2, 28, 15) {real, imag} */,
  {32'h4573dbf9, 32'h00000000} /* (2, 28, 14) {real, imag} */,
  {32'h455279d6, 32'h00000000} /* (2, 28, 13) {real, imag} */,
  {32'h453c9b6b, 32'h00000000} /* (2, 28, 12) {real, imag} */,
  {32'h44bbde3a, 32'h00000000} /* (2, 28, 11) {real, imag} */,
  {32'hc3abe010, 32'h00000000} /* (2, 28, 10) {real, imag} */,
  {32'hc51f6a82, 32'h00000000} /* (2, 28, 9) {real, imag} */,
  {32'hc537dacd, 32'h00000000} /* (2, 28, 8) {real, imag} */,
  {32'hc56b45d9, 32'h00000000} /* (2, 28, 7) {real, imag} */,
  {32'hc5107588, 32'h00000000} /* (2, 28, 6) {real, imag} */,
  {32'hc5292a0b, 32'h00000000} /* (2, 28, 5) {real, imag} */,
  {32'hc5800f27, 32'h00000000} /* (2, 28, 4) {real, imag} */,
  {32'hc5557d00, 32'h00000000} /* (2, 28, 3) {real, imag} */,
  {32'hc528e45a, 32'h00000000} /* (2, 28, 2) {real, imag} */,
  {32'hc501d98d, 32'h00000000} /* (2, 28, 1) {real, imag} */,
  {32'hc4bec628, 32'h00000000} /* (2, 28, 0) {real, imag} */,
  {32'hc4e300f7, 32'h00000000} /* (2, 27, 31) {real, imag} */,
  {32'hc537cf5c, 32'h00000000} /* (2, 27, 30) {real, imag} */,
  {32'hc5267ade, 32'h00000000} /* (2, 27, 29) {real, imag} */,
  {32'hc5404270, 32'h00000000} /* (2, 27, 28) {real, imag} */,
  {32'hc57e3048, 32'h00000000} /* (2, 27, 27) {real, imag} */,
  {32'hc5742b4d, 32'h00000000} /* (2, 27, 26) {real, imag} */,
  {32'hc5517ad1, 32'h00000000} /* (2, 27, 25) {real, imag} */,
  {32'hc537f969, 32'h00000000} /* (2, 27, 24) {real, imag} */,
  {32'hc51f9675, 32'h00000000} /* (2, 27, 23) {real, imag} */,
  {32'hc4d122fc, 32'h00000000} /* (2, 27, 22) {real, imag} */,
  {32'h4322e4c8, 32'h00000000} /* (2, 27, 21) {real, imag} */,
  {32'h45396fd0, 32'h00000000} /* (2, 27, 20) {real, imag} */,
  {32'h45986daa, 32'h00000000} /* (2, 27, 19) {real, imag} */,
  {32'h4585e2e1, 32'h00000000} /* (2, 27, 18) {real, imag} */,
  {32'h4592d64e, 32'h00000000} /* (2, 27, 17) {real, imag} */,
  {32'h458fc77c, 32'h00000000} /* (2, 27, 16) {real, imag} */,
  {32'h457b9534, 32'h00000000} /* (2, 27, 15) {real, imag} */,
  {32'h4567e3bc, 32'h00000000} /* (2, 27, 14) {real, imag} */,
  {32'h458494e5, 32'h00000000} /* (2, 27, 13) {real, imag} */,
  {32'h454924c4, 32'h00000000} /* (2, 27, 12) {real, imag} */,
  {32'h451a7134, 32'h00000000} /* (2, 27, 11) {real, imag} */,
  {32'hc415575c, 32'h00000000} /* (2, 27, 10) {real, imag} */,
  {32'hc4cf238e, 32'h00000000} /* (2, 27, 9) {real, imag} */,
  {32'hc505ac81, 32'h00000000} /* (2, 27, 8) {real, imag} */,
  {32'hc555faef, 32'h00000000} /* (2, 27, 7) {real, imag} */,
  {32'hc53f97e8, 32'h00000000} /* (2, 27, 6) {real, imag} */,
  {32'hc5650ad2, 32'h00000000} /* (2, 27, 5) {real, imag} */,
  {32'hc53e85cc, 32'h00000000} /* (2, 27, 4) {real, imag} */,
  {32'hc550e8b3, 32'h00000000} /* (2, 27, 3) {real, imag} */,
  {32'hc591127d, 32'h00000000} /* (2, 27, 2) {real, imag} */,
  {32'hc51061c0, 32'h00000000} /* (2, 27, 1) {real, imag} */,
  {32'hc504308e, 32'h00000000} /* (2, 27, 0) {real, imag} */,
  {32'hc51e0944, 32'h00000000} /* (2, 26, 31) {real, imag} */,
  {32'hc53a1a19, 32'h00000000} /* (2, 26, 30) {real, imag} */,
  {32'hc52bbb5a, 32'h00000000} /* (2, 26, 29) {real, imag} */,
  {32'hc57dd9b0, 32'h00000000} /* (2, 26, 28) {real, imag} */,
  {32'hc55fc3b6, 32'h00000000} /* (2, 26, 27) {real, imag} */,
  {32'hc53040da, 32'h00000000} /* (2, 26, 26) {real, imag} */,
  {32'hc55b4ff6, 32'h00000000} /* (2, 26, 25) {real, imag} */,
  {32'hc5368989, 32'h00000000} /* (2, 26, 24) {real, imag} */,
  {32'hc52e0c45, 32'h00000000} /* (2, 26, 23) {real, imag} */,
  {32'hc4908601, 32'h00000000} /* (2, 26, 22) {real, imag} */,
  {32'h44383469, 32'h00000000} /* (2, 26, 21) {real, imag} */,
  {32'h4571e5c7, 32'h00000000} /* (2, 26, 20) {real, imag} */,
  {32'h4582240e, 32'h00000000} /* (2, 26, 19) {real, imag} */,
  {32'h456d7581, 32'h00000000} /* (2, 26, 18) {real, imag} */,
  {32'h459840d4, 32'h00000000} /* (2, 26, 17) {real, imag} */,
  {32'h45883bcf, 32'h00000000} /* (2, 26, 16) {real, imag} */,
  {32'h4562204a, 32'h00000000} /* (2, 26, 15) {real, imag} */,
  {32'h458d5786, 32'h00000000} /* (2, 26, 14) {real, imag} */,
  {32'h45735c74, 32'h00000000} /* (2, 26, 13) {real, imag} */,
  {32'h458acd7c, 32'h00000000} /* (2, 26, 12) {real, imag} */,
  {32'h44fd69cc, 32'h00000000} /* (2, 26, 11) {real, imag} */,
  {32'h43d691c4, 32'h00000000} /* (2, 26, 10) {real, imag} */,
  {32'hc4b6cb1f, 32'h00000000} /* (2, 26, 9) {real, imag} */,
  {32'hc4f617b6, 32'h00000000} /* (2, 26, 8) {real, imag} */,
  {32'hc51888dd, 32'h00000000} /* (2, 26, 7) {real, imag} */,
  {32'hc55516b2, 32'h00000000} /* (2, 26, 6) {real, imag} */,
  {32'hc51bc29a, 32'h00000000} /* (2, 26, 5) {real, imag} */,
  {32'hc518c28f, 32'h00000000} /* (2, 26, 4) {real, imag} */,
  {32'hc54bf0e7, 32'h00000000} /* (2, 26, 3) {real, imag} */,
  {32'hc5628d91, 32'h00000000} /* (2, 26, 2) {real, imag} */,
  {32'hc54b3f0a, 32'h00000000} /* (2, 26, 1) {real, imag} */,
  {32'hc502c3fa, 32'h00000000} /* (2, 26, 0) {real, imag} */,
  {32'hc5196d89, 32'h00000000} /* (2, 25, 31) {real, imag} */,
  {32'hc55a90d9, 32'h00000000} /* (2, 25, 30) {real, imag} */,
  {32'hc535731e, 32'h00000000} /* (2, 25, 29) {real, imag} */,
  {32'hc543be88, 32'h00000000} /* (2, 25, 28) {real, imag} */,
  {32'hc567b227, 32'h00000000} /* (2, 25, 27) {real, imag} */,
  {32'hc5496fb2, 32'h00000000} /* (2, 25, 26) {real, imag} */,
  {32'hc5755c3c, 32'h00000000} /* (2, 25, 25) {real, imag} */,
  {32'hc5618654, 32'h00000000} /* (2, 25, 24) {real, imag} */,
  {32'hc50ff869, 32'h00000000} /* (2, 25, 23) {real, imag} */,
  {32'hc4ddc7a0, 32'h00000000} /* (2, 25, 22) {real, imag} */,
  {32'h4484c669, 32'h00000000} /* (2, 25, 21) {real, imag} */,
  {32'h4562290e, 32'h00000000} /* (2, 25, 20) {real, imag} */,
  {32'h4578500b, 32'h00000000} /* (2, 25, 19) {real, imag} */,
  {32'h459318f3, 32'h00000000} /* (2, 25, 18) {real, imag} */,
  {32'h45887cbd, 32'h00000000} /* (2, 25, 17) {real, imag} */,
  {32'h457efb40, 32'h00000000} /* (2, 25, 16) {real, imag} */,
  {32'h458d0aec, 32'h00000000} /* (2, 25, 15) {real, imag} */,
  {32'h459634a5, 32'h00000000} /* (2, 25, 14) {real, imag} */,
  {32'h4551ed84, 32'h00000000} /* (2, 25, 13) {real, imag} */,
  {32'h453622bc, 32'h00000000} /* (2, 25, 12) {real, imag} */,
  {32'h454926e3, 32'h00000000} /* (2, 25, 11) {real, imag} */,
  {32'h43eb23c4, 32'h00000000} /* (2, 25, 10) {real, imag} */,
  {32'hc4ea1cb8, 32'h00000000} /* (2, 25, 9) {real, imag} */,
  {32'hc52aa440, 32'h00000000} /* (2, 25, 8) {real, imag} */,
  {32'hc5334685, 32'h00000000} /* (2, 25, 7) {real, imag} */,
  {32'hc559d7f8, 32'h00000000} /* (2, 25, 6) {real, imag} */,
  {32'hc54d2414, 32'h00000000} /* (2, 25, 5) {real, imag} */,
  {32'hc520ea48, 32'h00000000} /* (2, 25, 4) {real, imag} */,
  {32'hc5457153, 32'h00000000} /* (2, 25, 3) {real, imag} */,
  {32'hc5661fb6, 32'h00000000} /* (2, 25, 2) {real, imag} */,
  {32'hc53b038a, 32'h00000000} /* (2, 25, 1) {real, imag} */,
  {32'hc558d7c0, 32'h00000000} /* (2, 25, 0) {real, imag} */,
  {32'hc53e39bb, 32'h00000000} /* (2, 24, 31) {real, imag} */,
  {32'hc548aea8, 32'h00000000} /* (2, 24, 30) {real, imag} */,
  {32'hc53277e4, 32'h00000000} /* (2, 24, 29) {real, imag} */,
  {32'hc53a4fc8, 32'h00000000} /* (2, 24, 28) {real, imag} */,
  {32'hc560bcc2, 32'h00000000} /* (2, 24, 27) {real, imag} */,
  {32'hc5809ab0, 32'h00000000} /* (2, 24, 26) {real, imag} */,
  {32'hc561c28d, 32'h00000000} /* (2, 24, 25) {real, imag} */,
  {32'hc52bc70d, 32'h00000000} /* (2, 24, 24) {real, imag} */,
  {32'hc4f37231, 32'h00000000} /* (2, 24, 23) {real, imag} */,
  {32'hc4ce23e6, 32'h00000000} /* (2, 24, 22) {real, imag} */,
  {32'h4499ffe8, 32'h00000000} /* (2, 24, 21) {real, imag} */,
  {32'h4543e784, 32'h00000000} /* (2, 24, 20) {real, imag} */,
  {32'h4570ae3c, 32'h00000000} /* (2, 24, 19) {real, imag} */,
  {32'h45989188, 32'h00000000} /* (2, 24, 18) {real, imag} */,
  {32'h458ada74, 32'h00000000} /* (2, 24, 17) {real, imag} */,
  {32'h45838330, 32'h00000000} /* (2, 24, 16) {real, imag} */,
  {32'h4577100f, 32'h00000000} /* (2, 24, 15) {real, imag} */,
  {32'h453e68ba, 32'h00000000} /* (2, 24, 14) {real, imag} */,
  {32'h454de298, 32'h00000000} /* (2, 24, 13) {real, imag} */,
  {32'h453bbbc2, 32'h00000000} /* (2, 24, 12) {real, imag} */,
  {32'h44f18994, 32'h00000000} /* (2, 24, 11) {real, imag} */,
  {32'hc4a97062, 32'h00000000} /* (2, 24, 10) {real, imag} */,
  {32'hc51451a1, 32'h00000000} /* (2, 24, 9) {real, imag} */,
  {32'hc4baac12, 32'h00000000} /* (2, 24, 8) {real, imag} */,
  {32'hc549a1de, 32'h00000000} /* (2, 24, 7) {real, imag} */,
  {32'hc53a7f55, 32'h00000000} /* (2, 24, 6) {real, imag} */,
  {32'hc551038c, 32'h00000000} /* (2, 24, 5) {real, imag} */,
  {32'hc536d47e, 32'h00000000} /* (2, 24, 4) {real, imag} */,
  {32'hc55e811c, 32'h00000000} /* (2, 24, 3) {real, imag} */,
  {32'hc5661218, 32'h00000000} /* (2, 24, 2) {real, imag} */,
  {32'hc57a5301, 32'h00000000} /* (2, 24, 1) {real, imag} */,
  {32'hc53c9451, 32'h00000000} /* (2, 24, 0) {real, imag} */,
  {32'hc51c0e17, 32'h00000000} /* (2, 23, 31) {real, imag} */,
  {32'hc51be6c1, 32'h00000000} /* (2, 23, 30) {real, imag} */,
  {32'hc55b85ea, 32'h00000000} /* (2, 23, 29) {real, imag} */,
  {32'hc523309a, 32'h00000000} /* (2, 23, 28) {real, imag} */,
  {32'hc5416e38, 32'h00000000} /* (2, 23, 27) {real, imag} */,
  {32'hc53f3f1a, 32'h00000000} /* (2, 23, 26) {real, imag} */,
  {32'hc52c6ff2, 32'h00000000} /* (2, 23, 25) {real, imag} */,
  {32'hc4e29acc, 32'h00000000} /* (2, 23, 24) {real, imag} */,
  {32'hc4b8b906, 32'h00000000} /* (2, 23, 23) {real, imag} */,
  {32'hc48c1668, 32'h00000000} /* (2, 23, 22) {real, imag} */,
  {32'h4403a0be, 32'h00000000} /* (2, 23, 21) {real, imag} */,
  {32'h45327d22, 32'h00000000} /* (2, 23, 20) {real, imag} */,
  {32'h456c6a9e, 32'h00000000} /* (2, 23, 19) {real, imag} */,
  {32'h456ec928, 32'h00000000} /* (2, 23, 18) {real, imag} */,
  {32'h45a12cf8, 32'h00000000} /* (2, 23, 17) {real, imag} */,
  {32'h4554fbea, 32'h00000000} /* (2, 23, 16) {real, imag} */,
  {32'h453dfbf7, 32'h00000000} /* (2, 23, 15) {real, imag} */,
  {32'h45524919, 32'h00000000} /* (2, 23, 14) {real, imag} */,
  {32'h453dd3fe, 32'h00000000} /* (2, 23, 13) {real, imag} */,
  {32'h450724c0, 32'h00000000} /* (2, 23, 12) {real, imag} */,
  {32'h450024e8, 32'h00000000} /* (2, 23, 11) {real, imag} */,
  {32'hc343c8c8, 32'h00000000} /* (2, 23, 10) {real, imag} */,
  {32'hc513c872, 32'h00000000} /* (2, 23, 9) {real, imag} */,
  {32'hc4f0045c, 32'h00000000} /* (2, 23, 8) {real, imag} */,
  {32'hc51b1f61, 32'h00000000} /* (2, 23, 7) {real, imag} */,
  {32'hc500b6e8, 32'h00000000} /* (2, 23, 6) {real, imag} */,
  {32'hc50dfadc, 32'h00000000} /* (2, 23, 5) {real, imag} */,
  {32'hc528cbb8, 32'h00000000} /* (2, 23, 4) {real, imag} */,
  {32'hc51267e6, 32'h00000000} /* (2, 23, 3) {real, imag} */,
  {32'hc54d9276, 32'h00000000} /* (2, 23, 2) {real, imag} */,
  {32'hc592b522, 32'h00000000} /* (2, 23, 1) {real, imag} */,
  {32'hc5193176, 32'h00000000} /* (2, 23, 0) {real, imag} */,
  {32'hc4dc8bc6, 32'h00000000} /* (2, 22, 31) {real, imag} */,
  {32'hc5027da0, 32'h00000000} /* (2, 22, 30) {real, imag} */,
  {32'hc525b2c7, 32'h00000000} /* (2, 22, 29) {real, imag} */,
  {32'hc4f139d3, 32'h00000000} /* (2, 22, 28) {real, imag} */,
  {32'hc520c7c7, 32'h00000000} /* (2, 22, 27) {real, imag} */,
  {32'hc4e0469c, 32'h00000000} /* (2, 22, 26) {real, imag} */,
  {32'hc498b789, 32'h00000000} /* (2, 22, 25) {real, imag} */,
  {32'hc4d2fae5, 32'h00000000} /* (2, 22, 24) {real, imag} */,
  {32'hc4407df8, 32'h00000000} /* (2, 22, 23) {real, imag} */,
  {32'h418deba0, 32'h00000000} /* (2, 22, 22) {real, imag} */,
  {32'hc45aa608, 32'h00000000} /* (2, 22, 21) {real, imag} */,
  {32'h44d8a783, 32'h00000000} /* (2, 22, 20) {real, imag} */,
  {32'h454ec1c9, 32'h00000000} /* (2, 22, 19) {real, imag} */,
  {32'h454363e8, 32'h00000000} /* (2, 22, 18) {real, imag} */,
  {32'h452270d0, 32'h00000000} /* (2, 22, 17) {real, imag} */,
  {32'h45334736, 32'h00000000} /* (2, 22, 16) {real, imag} */,
  {32'h45222bad, 32'h00000000} /* (2, 22, 15) {real, imag} */,
  {32'h45661638, 32'h00000000} /* (2, 22, 14) {real, imag} */,
  {32'h454531c1, 32'h00000000} /* (2, 22, 13) {real, imag} */,
  {32'h45183914, 32'h00000000} /* (2, 22, 12) {real, imag} */,
  {32'h4497293c, 32'h00000000} /* (2, 22, 11) {real, imag} */,
  {32'hc4614979, 32'h00000000} /* (2, 22, 10) {real, imag} */,
  {32'hc4cfe779, 32'h00000000} /* (2, 22, 9) {real, imag} */,
  {32'hc53fd93e, 32'h00000000} /* (2, 22, 8) {real, imag} */,
  {32'hc4e6cd74, 32'h00000000} /* (2, 22, 7) {real, imag} */,
  {32'hc4cc8c58, 32'h00000000} /* (2, 22, 6) {real, imag} */,
  {32'hc4f58714, 32'h00000000} /* (2, 22, 5) {real, imag} */,
  {32'hc4b586e1, 32'h00000000} /* (2, 22, 4) {real, imag} */,
  {32'hc50c0991, 32'h00000000} /* (2, 22, 3) {real, imag} */,
  {32'hc518f92a, 32'h00000000} /* (2, 22, 2) {real, imag} */,
  {32'hc4fc3e6b, 32'h00000000} /* (2, 22, 1) {real, imag} */,
  {32'hc52b80aa, 32'h00000000} /* (2, 22, 0) {real, imag} */,
  {32'hc481f552, 32'h00000000} /* (2, 21, 31) {real, imag} */,
  {32'hc438db32, 32'h00000000} /* (2, 21, 30) {real, imag} */,
  {32'hc3349754, 32'h00000000} /* (2, 21, 29) {real, imag} */,
  {32'hc42e3530, 32'h00000000} /* (2, 21, 28) {real, imag} */,
  {32'hc48022dc, 32'h00000000} /* (2, 21, 27) {real, imag} */,
  {32'h428de0fa, 32'h00000000} /* (2, 21, 26) {real, imag} */,
  {32'h43e5dbda, 32'h00000000} /* (2, 21, 25) {real, imag} */,
  {32'h4344f570, 32'h00000000} /* (2, 21, 24) {real, imag} */,
  {32'h443cf982, 32'h00000000} /* (2, 21, 23) {real, imag} */,
  {32'h419c9114, 32'h00000000} /* (2, 21, 22) {real, imag} */,
  {32'hc3dde6cf, 32'h00000000} /* (2, 21, 21) {real, imag} */,
  {32'h4498fe93, 32'h00000000} /* (2, 21, 20) {real, imag} */,
  {32'h44b31d60, 32'h00000000} /* (2, 21, 19) {real, imag} */,
  {32'h44ae3e8f, 32'h00000000} /* (2, 21, 18) {real, imag} */,
  {32'h44d39064, 32'h00000000} /* (2, 21, 17) {real, imag} */,
  {32'h450a429d, 32'h00000000} /* (2, 21, 16) {real, imag} */,
  {32'h4414e758, 32'h00000000} /* (2, 21, 15) {real, imag} */,
  {32'h449331f5, 32'h00000000} /* (2, 21, 14) {real, imag} */,
  {32'h449c4840, 32'h00000000} /* (2, 21, 13) {real, imag} */,
  {32'h43e41ac4, 32'h00000000} /* (2, 21, 12) {real, imag} */,
  {32'h448d656e, 32'h00000000} /* (2, 21, 11) {real, imag} */,
  {32'h43d00594, 32'h00000000} /* (2, 21, 10) {real, imag} */,
  {32'hc400ce26, 32'h00000000} /* (2, 21, 9) {real, imag} */,
  {32'hc483a2de, 32'h00000000} /* (2, 21, 8) {real, imag} */,
  {32'hc44a3d86, 32'h00000000} /* (2, 21, 7) {real, imag} */,
  {32'hc187288c, 32'h00000000} /* (2, 21, 6) {real, imag} */,
  {32'hc38394d3, 32'h00000000} /* (2, 21, 5) {real, imag} */,
  {32'hc463a392, 32'h00000000} /* (2, 21, 4) {real, imag} */,
  {32'hc47716b0, 32'h00000000} /* (2, 21, 3) {real, imag} */,
  {32'hc498d355, 32'h00000000} /* (2, 21, 2) {real, imag} */,
  {32'hc4af5924, 32'h00000000} /* (2, 21, 1) {real, imag} */,
  {32'hc46fb81c, 32'h00000000} /* (2, 21, 0) {real, imag} */,
  {32'h43d1057e, 32'h00000000} /* (2, 20, 31) {real, imag} */,
  {32'h44e07c6b, 32'h00000000} /* (2, 20, 30) {real, imag} */,
  {32'h44fffa23, 32'h00000000} /* (2, 20, 29) {real, imag} */,
  {32'h453a6439, 32'h00000000} /* (2, 20, 28) {real, imag} */,
  {32'h451bcedd, 32'h00000000} /* (2, 20, 27) {real, imag} */,
  {32'h44c6a40e, 32'h00000000} /* (2, 20, 26) {real, imag} */,
  {32'h45593517, 32'h00000000} /* (2, 20, 25) {real, imag} */,
  {32'h452f3cc2, 32'h00000000} /* (2, 20, 24) {real, imag} */,
  {32'h44f677de, 32'h00000000} /* (2, 20, 23) {real, imag} */,
  {32'h44eeadae, 32'h00000000} /* (2, 20, 22) {real, imag} */,
  {32'h443d334e, 32'h00000000} /* (2, 20, 21) {real, imag} */,
  {32'hc4093a3f, 32'h00000000} /* (2, 20, 20) {real, imag} */,
  {32'hc4395dfc, 32'h00000000} /* (2, 20, 19) {real, imag} */,
  {32'hc35f6d60, 32'h00000000} /* (2, 20, 18) {real, imag} */,
  {32'hc490180c, 32'h00000000} /* (2, 20, 17) {real, imag} */,
  {32'hc4376415, 32'h00000000} /* (2, 20, 16) {real, imag} */,
  {32'hc463b355, 32'h00000000} /* (2, 20, 15) {real, imag} */,
  {32'hc5144edc, 32'h00000000} /* (2, 20, 14) {real, imag} */,
  {32'hc4af5de5, 32'h00000000} /* (2, 20, 13) {real, imag} */,
  {32'hc47070f3, 32'h00000000} /* (2, 20, 12) {real, imag} */,
  {32'hc4516928, 32'h00000000} /* (2, 20, 11) {real, imag} */,
  {32'hc2ad19d8, 32'h00000000} /* (2, 20, 10) {real, imag} */,
  {32'h44a498b2, 32'h00000000} /* (2, 20, 9) {real, imag} */,
  {32'h443d7d50, 32'h00000000} /* (2, 20, 8) {real, imag} */,
  {32'h4485b8c6, 32'h00000000} /* (2, 20, 7) {real, imag} */,
  {32'h45147c9d, 32'h00000000} /* (2, 20, 6) {real, imag} */,
  {32'h450a7158, 32'h00000000} /* (2, 20, 5) {real, imag} */,
  {32'h44bb8542, 32'h00000000} /* (2, 20, 4) {real, imag} */,
  {32'h448a2c95, 32'h00000000} /* (2, 20, 3) {real, imag} */,
  {32'h44a612dc, 32'h00000000} /* (2, 20, 2) {real, imag} */,
  {32'h44471787, 32'h00000000} /* (2, 20, 1) {real, imag} */,
  {32'h442518fb, 32'h00000000} /* (2, 20, 0) {real, imag} */,
  {32'h451724e6, 32'h00000000} /* (2, 19, 31) {real, imag} */,
  {32'h451c1a28, 32'h00000000} /* (2, 19, 30) {real, imag} */,
  {32'h4520e599, 32'h00000000} /* (2, 19, 29) {real, imag} */,
  {32'h45825186, 32'h00000000} /* (2, 19, 28) {real, imag} */,
  {32'h456da58d, 32'h00000000} /* (2, 19, 27) {real, imag} */,
  {32'h45485dad, 32'h00000000} /* (2, 19, 26) {real, imag} */,
  {32'h45685ee3, 32'h00000000} /* (2, 19, 25) {real, imag} */,
  {32'h45990404, 32'h00000000} /* (2, 19, 24) {real, imag} */,
  {32'h453ea0ce, 32'h00000000} /* (2, 19, 23) {real, imag} */,
  {32'h4528e2ae, 32'h00000000} /* (2, 19, 22) {real, imag} */,
  {32'h443a27f6, 32'h00000000} /* (2, 19, 21) {real, imag} */,
  {32'hc4a9a6e8, 32'h00000000} /* (2, 19, 20) {real, imag} */,
  {32'hc4c9f334, 32'h00000000} /* (2, 19, 19) {real, imag} */,
  {32'hc53b5e79, 32'h00000000} /* (2, 19, 18) {real, imag} */,
  {32'hc51151ce, 32'h00000000} /* (2, 19, 17) {real, imag} */,
  {32'hc4ef15bc, 32'h00000000} /* (2, 19, 16) {real, imag} */,
  {32'hc51c9a4c, 32'h00000000} /* (2, 19, 15) {real, imag} */,
  {32'hc4f7ef7b, 32'h00000000} /* (2, 19, 14) {real, imag} */,
  {32'hc509b321, 32'h00000000} /* (2, 19, 13) {real, imag} */,
  {32'hc4e87bac, 32'h00000000} /* (2, 19, 12) {real, imag} */,
  {32'hc4a1bbae, 32'h00000000} /* (2, 19, 11) {real, imag} */,
  {32'h447571cc, 32'h00000000} /* (2, 19, 10) {real, imag} */,
  {32'h44b2a5ea, 32'h00000000} /* (2, 19, 9) {real, imag} */,
  {32'h44f26aa2, 32'h00000000} /* (2, 19, 8) {real, imag} */,
  {32'h4527489e, 32'h00000000} /* (2, 19, 7) {real, imag} */,
  {32'h4518ff26, 32'h00000000} /* (2, 19, 6) {real, imag} */,
  {32'h451f370e, 32'h00000000} /* (2, 19, 5) {real, imag} */,
  {32'h45102ee4, 32'h00000000} /* (2, 19, 4) {real, imag} */,
  {32'h451f1f16, 32'h00000000} /* (2, 19, 3) {real, imag} */,
  {32'h4533b78b, 32'h00000000} /* (2, 19, 2) {real, imag} */,
  {32'h450680c2, 32'h00000000} /* (2, 19, 1) {real, imag} */,
  {32'h44ad8224, 32'h00000000} /* (2, 19, 0) {real, imag} */,
  {32'h45128682, 32'h00000000} /* (2, 18, 31) {real, imag} */,
  {32'h455166e4, 32'h00000000} /* (2, 18, 30) {real, imag} */,
  {32'h45487b57, 32'h00000000} /* (2, 18, 29) {real, imag} */,
  {32'h457bbe12, 32'h00000000} /* (2, 18, 28) {real, imag} */,
  {32'h457c9c05, 32'h00000000} /* (2, 18, 27) {real, imag} */,
  {32'h4586ce2d, 32'h00000000} /* (2, 18, 26) {real, imag} */,
  {32'h458eb0bc, 32'h00000000} /* (2, 18, 25) {real, imag} */,
  {32'h45552159, 32'h00000000} /* (2, 18, 24) {real, imag} */,
  {32'h4537f236, 32'h00000000} /* (2, 18, 23) {real, imag} */,
  {32'h4505f7ed, 32'h00000000} /* (2, 18, 22) {real, imag} */,
  {32'h440c74e2, 32'h00000000} /* (2, 18, 21) {real, imag} */,
  {32'hc4e0190c, 32'h00000000} /* (2, 18, 20) {real, imag} */,
  {32'hc524f8cc, 32'h00000000} /* (2, 18, 19) {real, imag} */,
  {32'hc560390a, 32'h00000000} /* (2, 18, 18) {real, imag} */,
  {32'hc5395cb3, 32'h00000000} /* (2, 18, 17) {real, imag} */,
  {32'hc531005b, 32'h00000000} /* (2, 18, 16) {real, imag} */,
  {32'hc52e504e, 32'h00000000} /* (2, 18, 15) {real, imag} */,
  {32'hc5183448, 32'h00000000} /* (2, 18, 14) {real, imag} */,
  {32'hc516aaaf, 32'h00000000} /* (2, 18, 13) {real, imag} */,
  {32'hc525a4a0, 32'h00000000} /* (2, 18, 12) {real, imag} */,
  {32'hc509461d, 32'h00000000} /* (2, 18, 11) {real, imag} */,
  {32'h443ce0e8, 32'h00000000} /* (2, 18, 10) {real, imag} */,
  {32'h44eea174, 32'h00000000} /* (2, 18, 9) {real, imag} */,
  {32'h45304285, 32'h00000000} /* (2, 18, 8) {real, imag} */,
  {32'h45687cee, 32'h00000000} /* (2, 18, 7) {real, imag} */,
  {32'h4514314d, 32'h00000000} /* (2, 18, 6) {real, imag} */,
  {32'h45385590, 32'h00000000} /* (2, 18, 5) {real, imag} */,
  {32'h454252de, 32'h00000000} /* (2, 18, 4) {real, imag} */,
  {32'h45107566, 32'h00000000} /* (2, 18, 3) {real, imag} */,
  {32'h454a57c0, 32'h00000000} /* (2, 18, 2) {real, imag} */,
  {32'h452eab79, 32'h00000000} /* (2, 18, 1) {real, imag} */,
  {32'h44fd0a6a, 32'h00000000} /* (2, 18, 0) {real, imag} */,
  {32'h452344ea, 32'h00000000} /* (2, 17, 31) {real, imag} */,
  {32'h45436abe, 32'h00000000} /* (2, 17, 30) {real, imag} */,
  {32'h45815ae6, 32'h00000000} /* (2, 17, 29) {real, imag} */,
  {32'h454eca58, 32'h00000000} /* (2, 17, 28) {real, imag} */,
  {32'h45798cff, 32'h00000000} /* (2, 17, 27) {real, imag} */,
  {32'h4568ab98, 32'h00000000} /* (2, 17, 26) {real, imag} */,
  {32'h4560ed8d, 32'h00000000} /* (2, 17, 25) {real, imag} */,
  {32'h453cc7ab, 32'h00000000} /* (2, 17, 24) {real, imag} */,
  {32'h4556b061, 32'h00000000} /* (2, 17, 23) {real, imag} */,
  {32'h45319938, 32'h00000000} /* (2, 17, 22) {real, imag} */,
  {32'h442d6880, 32'h00000000} /* (2, 17, 21) {real, imag} */,
  {32'hc46a45cc, 32'h00000000} /* (2, 17, 20) {real, imag} */,
  {32'hc5184098, 32'h00000000} /* (2, 17, 19) {real, imag} */,
  {32'hc54ac2e9, 32'h00000000} /* (2, 17, 18) {real, imag} */,
  {32'hc5a1533a, 32'h00000000} /* (2, 17, 17) {real, imag} */,
  {32'hc57177a0, 32'h00000000} /* (2, 17, 16) {real, imag} */,
  {32'hc530e846, 32'h00000000} /* (2, 17, 15) {real, imag} */,
  {32'hc553581a, 32'h00000000} /* (2, 17, 14) {real, imag} */,
  {32'hc54dfc9d, 32'h00000000} /* (2, 17, 13) {real, imag} */,
  {32'hc50661c8, 32'h00000000} /* (2, 17, 12) {real, imag} */,
  {32'hc49f128a, 32'h00000000} /* (2, 17, 11) {real, imag} */,
  {32'hc0cafc00, 32'h00000000} /* (2, 17, 10) {real, imag} */,
  {32'h450e54ed, 32'h00000000} /* (2, 17, 9) {real, imag} */,
  {32'h452936b5, 32'h00000000} /* (2, 17, 8) {real, imag} */,
  {32'h455cf08f, 32'h00000000} /* (2, 17, 7) {real, imag} */,
  {32'h458d32fc, 32'h00000000} /* (2, 17, 6) {real, imag} */,
  {32'h4548141a, 32'h00000000} /* (2, 17, 5) {real, imag} */,
  {32'h453bc85b, 32'h00000000} /* (2, 17, 4) {real, imag} */,
  {32'h453a76a4, 32'h00000000} /* (2, 17, 3) {real, imag} */,
  {32'h452d19fd, 32'h00000000} /* (2, 17, 2) {real, imag} */,
  {32'h4521aaf1, 32'h00000000} /* (2, 17, 1) {real, imag} */,
  {32'h453d0036, 32'h00000000} /* (2, 17, 0) {real, imag} */,
  {32'h45631a45, 32'h00000000} /* (2, 16, 31) {real, imag} */,
  {32'h4567061e, 32'h00000000} /* (2, 16, 30) {real, imag} */,
  {32'h454748b2, 32'h00000000} /* (2, 16, 29) {real, imag} */,
  {32'h4561f9f7, 32'h00000000} /* (2, 16, 28) {real, imag} */,
  {32'h454b5027, 32'h00000000} /* (2, 16, 27) {real, imag} */,
  {32'h457b5559, 32'h00000000} /* (2, 16, 26) {real, imag} */,
  {32'h4560eaa8, 32'h00000000} /* (2, 16, 25) {real, imag} */,
  {32'h455e8e56, 32'h00000000} /* (2, 16, 24) {real, imag} */,
  {32'h45621c32, 32'h00000000} /* (2, 16, 23) {real, imag} */,
  {32'h45433ffb, 32'h00000000} /* (2, 16, 22) {real, imag} */,
  {32'h44a5c2de, 32'h00000000} /* (2, 16, 21) {real, imag} */,
  {32'hc4f418c8, 32'h00000000} /* (2, 16, 20) {real, imag} */,
  {32'hc534af62, 32'h00000000} /* (2, 16, 19) {real, imag} */,
  {32'hc54892b0, 32'h00000000} /* (2, 16, 18) {real, imag} */,
  {32'hc555d1ae, 32'h00000000} /* (2, 16, 17) {real, imag} */,
  {32'hc56bdc78, 32'h00000000} /* (2, 16, 16) {real, imag} */,
  {32'hc5707c37, 32'h00000000} /* (2, 16, 15) {real, imag} */,
  {32'hc5496030, 32'h00000000} /* (2, 16, 14) {real, imag} */,
  {32'hc525d806, 32'h00000000} /* (2, 16, 13) {real, imag} */,
  {32'hc51b94f5, 32'h00000000} /* (2, 16, 12) {real, imag} */,
  {32'hc4cd32fa, 32'h00000000} /* (2, 16, 11) {real, imag} */,
  {32'h448a65d6, 32'h00000000} /* (2, 16, 10) {real, imag} */,
  {32'h44f99329, 32'h00000000} /* (2, 16, 9) {real, imag} */,
  {32'h4542be7e, 32'h00000000} /* (2, 16, 8) {real, imag} */,
  {32'h4558a304, 32'h00000000} /* (2, 16, 7) {real, imag} */,
  {32'h456f1f8d, 32'h00000000} /* (2, 16, 6) {real, imag} */,
  {32'h455e53a1, 32'h00000000} /* (2, 16, 5) {real, imag} */,
  {32'h4520c344, 32'h00000000} /* (2, 16, 4) {real, imag} */,
  {32'h4585bdbb, 32'h00000000} /* (2, 16, 3) {real, imag} */,
  {32'h45795fbc, 32'h00000000} /* (2, 16, 2) {real, imag} */,
  {32'h45335466, 32'h00000000} /* (2, 16, 1) {real, imag} */,
  {32'h4553be84, 32'h00000000} /* (2, 16, 0) {real, imag} */,
  {32'h4571b3e4, 32'h00000000} /* (2, 15, 31) {real, imag} */,
  {32'h4570c213, 32'h00000000} /* (2, 15, 30) {real, imag} */,
  {32'h4561c436, 32'h00000000} /* (2, 15, 29) {real, imag} */,
  {32'h458a6e5c, 32'h00000000} /* (2, 15, 28) {real, imag} */,
  {32'h45596069, 32'h00000000} /* (2, 15, 27) {real, imag} */,
  {32'h455fe699, 32'h00000000} /* (2, 15, 26) {real, imag} */,
  {32'h45500d5b, 32'h00000000} /* (2, 15, 25) {real, imag} */,
  {32'h456aa87c, 32'h00000000} /* (2, 15, 24) {real, imag} */,
  {32'h45364b7d, 32'h00000000} /* (2, 15, 23) {real, imag} */,
  {32'h452876fa, 32'h00000000} /* (2, 15, 22) {real, imag} */,
  {32'h448e378a, 32'h00000000} /* (2, 15, 21) {real, imag} */,
  {32'hc4acab38, 32'h00000000} /* (2, 15, 20) {real, imag} */,
  {32'hc50f3d2f, 32'h00000000} /* (2, 15, 19) {real, imag} */,
  {32'hc53050f1, 32'h00000000} /* (2, 15, 18) {real, imag} */,
  {32'hc57884f3, 32'h00000000} /* (2, 15, 17) {real, imag} */,
  {32'hc55c5dc5, 32'h00000000} /* (2, 15, 16) {real, imag} */,
  {32'hc54a1304, 32'h00000000} /* (2, 15, 15) {real, imag} */,
  {32'hc554759f, 32'h00000000} /* (2, 15, 14) {real, imag} */,
  {32'hc535f140, 32'h00000000} /* (2, 15, 13) {real, imag} */,
  {32'hc524e74e, 32'h00000000} /* (2, 15, 12) {real, imag} */,
  {32'hc4d06db6, 32'h00000000} /* (2, 15, 11) {real, imag} */,
  {32'h440e64f4, 32'h00000000} /* (2, 15, 10) {real, imag} */,
  {32'h44eafa4a, 32'h00000000} /* (2, 15, 9) {real, imag} */,
  {32'h4555c07c, 32'h00000000} /* (2, 15, 8) {real, imag} */,
  {32'h45775d37, 32'h00000000} /* (2, 15, 7) {real, imag} */,
  {32'h451df54e, 32'h00000000} /* (2, 15, 6) {real, imag} */,
  {32'h45326c19, 32'h00000000} /* (2, 15, 5) {real, imag} */,
  {32'h4565c404, 32'h00000000} /* (2, 15, 4) {real, imag} */,
  {32'h455ae629, 32'h00000000} /* (2, 15, 3) {real, imag} */,
  {32'h457568c7, 32'h00000000} /* (2, 15, 2) {real, imag} */,
  {32'h455acb53, 32'h00000000} /* (2, 15, 1) {real, imag} */,
  {32'h452f5295, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'h45734b2e, 32'h00000000} /* (2, 14, 31) {real, imag} */,
  {32'h4576256f, 32'h00000000} /* (2, 14, 30) {real, imag} */,
  {32'h458cf09e, 32'h00000000} /* (2, 14, 29) {real, imag} */,
  {32'h4581c9ae, 32'h00000000} /* (2, 14, 28) {real, imag} */,
  {32'h457e5e48, 32'h00000000} /* (2, 14, 27) {real, imag} */,
  {32'h45744fad, 32'h00000000} /* (2, 14, 26) {real, imag} */,
  {32'h455c0fc9, 32'h00000000} /* (2, 14, 25) {real, imag} */,
  {32'h453dfc6b, 32'h00000000} /* (2, 14, 24) {real, imag} */,
  {32'h4541d3f1, 32'h00000000} /* (2, 14, 23) {real, imag} */,
  {32'h45204eaf, 32'h00000000} /* (2, 14, 22) {real, imag} */,
  {32'h4499821b, 32'h00000000} /* (2, 14, 21) {real, imag} */,
  {32'hc484974c, 32'h00000000} /* (2, 14, 20) {real, imag} */,
  {32'hc539fec3, 32'h00000000} /* (2, 14, 19) {real, imag} */,
  {32'hc53b96cb, 32'h00000000} /* (2, 14, 18) {real, imag} */,
  {32'hc5690640, 32'h00000000} /* (2, 14, 17) {real, imag} */,
  {32'hc5861fe2, 32'h00000000} /* (2, 14, 16) {real, imag} */,
  {32'hc538efd6, 32'h00000000} /* (2, 14, 15) {real, imag} */,
  {32'hc57ddb4b, 32'h00000000} /* (2, 14, 14) {real, imag} */,
  {32'hc55813e6, 32'h00000000} /* (2, 14, 13) {real, imag} */,
  {32'hc51a76e1, 32'h00000000} /* (2, 14, 12) {real, imag} */,
  {32'hc4d7ba6c, 32'h00000000} /* (2, 14, 11) {real, imag} */,
  {32'h44a59be2, 32'h00000000} /* (2, 14, 10) {real, imag} */,
  {32'h4524d98b, 32'h00000000} /* (2, 14, 9) {real, imag} */,
  {32'h45669bd1, 32'h00000000} /* (2, 14, 8) {real, imag} */,
  {32'h4554a8eb, 32'h00000000} /* (2, 14, 7) {real, imag} */,
  {32'h453cb8d1, 32'h00000000} /* (2, 14, 6) {real, imag} */,
  {32'h4547f6c6, 32'h00000000} /* (2, 14, 5) {real, imag} */,
  {32'h453ecb0e, 32'h00000000} /* (2, 14, 4) {real, imag} */,
  {32'h45863f69, 32'h00000000} /* (2, 14, 3) {real, imag} */,
  {32'h4599bc36, 32'h00000000} /* (2, 14, 2) {real, imag} */,
  {32'h45716784, 32'h00000000} /* (2, 14, 1) {real, imag} */,
  {32'h453cf90a, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h4549736a, 32'h00000000} /* (2, 13, 31) {real, imag} */,
  {32'h4590a05f, 32'h00000000} /* (2, 13, 30) {real, imag} */,
  {32'h45aa26cf, 32'h00000000} /* (2, 13, 29) {real, imag} */,
  {32'h45a5361c, 32'h00000000} /* (2, 13, 28) {real, imag} */,
  {32'h45671386, 32'h00000000} /* (2, 13, 27) {real, imag} */,
  {32'h4589ba70, 32'h00000000} /* (2, 13, 26) {real, imag} */,
  {32'h455f871c, 32'h00000000} /* (2, 13, 25) {real, imag} */,
  {32'h456b5178, 32'h00000000} /* (2, 13, 24) {real, imag} */,
  {32'h45633240, 32'h00000000} /* (2, 13, 23) {real, imag} */,
  {32'h4556f62e, 32'h00000000} /* (2, 13, 22) {real, imag} */,
  {32'h443c034a, 32'h00000000} /* (2, 13, 21) {real, imag} */,
  {32'hc4cb4d06, 32'h00000000} /* (2, 13, 20) {real, imag} */,
  {32'hc50c461a, 32'h00000000} /* (2, 13, 19) {real, imag} */,
  {32'hc54300fa, 32'h00000000} /* (2, 13, 18) {real, imag} */,
  {32'hc551e574, 32'h00000000} /* (2, 13, 17) {real, imag} */,
  {32'hc5785074, 32'h00000000} /* (2, 13, 16) {real, imag} */,
  {32'hc549154c, 32'h00000000} /* (2, 13, 15) {real, imag} */,
  {32'hc56e5d3e, 32'h00000000} /* (2, 13, 14) {real, imag} */,
  {32'hc5559f1a, 32'h00000000} /* (2, 13, 13) {real, imag} */,
  {32'hc4f68a72, 32'h00000000} /* (2, 13, 12) {real, imag} */,
  {32'hc4cc4df7, 32'h00000000} /* (2, 13, 11) {real, imag} */,
  {32'h44828b06, 32'h00000000} /* (2, 13, 10) {real, imag} */,
  {32'h44e813a0, 32'h00000000} /* (2, 13, 9) {real, imag} */,
  {32'h45261360, 32'h00000000} /* (2, 13, 8) {real, imag} */,
  {32'h4534298e, 32'h00000000} /* (2, 13, 7) {real, imag} */,
  {32'h4548fd70, 32'h00000000} /* (2, 13, 6) {real, imag} */,
  {32'h454d9138, 32'h00000000} /* (2, 13, 5) {real, imag} */,
  {32'h4525a591, 32'h00000000} /* (2, 13, 4) {real, imag} */,
  {32'h453d8ede, 32'h00000000} /* (2, 13, 3) {real, imag} */,
  {32'h454696f8, 32'h00000000} /* (2, 13, 2) {real, imag} */,
  {32'h45634d5c, 32'h00000000} /* (2, 13, 1) {real, imag} */,
  {32'h4552085e, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'h4515e5ae, 32'h00000000} /* (2, 12, 31) {real, imag} */,
  {32'h454b2884, 32'h00000000} /* (2, 12, 30) {real, imag} */,
  {32'h45763c84, 32'h00000000} /* (2, 12, 29) {real, imag} */,
  {32'h4587b94e, 32'h00000000} /* (2, 12, 28) {real, imag} */,
  {32'h4558e70e, 32'h00000000} /* (2, 12, 27) {real, imag} */,
  {32'h451a78aa, 32'h00000000} /* (2, 12, 26) {real, imag} */,
  {32'h456248e9, 32'h00000000} /* (2, 12, 25) {real, imag} */,
  {32'h4562167e, 32'h00000000} /* (2, 12, 24) {real, imag} */,
  {32'h4559da73, 32'h00000000} /* (2, 12, 23) {real, imag} */,
  {32'h45018d6f, 32'h00000000} /* (2, 12, 22) {real, imag} */,
  {32'h4390d0b8, 32'h00000000} /* (2, 12, 21) {real, imag} */,
  {32'hc4b53e04, 32'h00000000} /* (2, 12, 20) {real, imag} */,
  {32'hc50b2c9a, 32'h00000000} /* (2, 12, 19) {real, imag} */,
  {32'hc528b07b, 32'h00000000} /* (2, 12, 18) {real, imag} */,
  {32'hc5403893, 32'h00000000} /* (2, 12, 17) {real, imag} */,
  {32'hc5366a58, 32'h00000000} /* (2, 12, 16) {real, imag} */,
  {32'hc557b9cc, 32'h00000000} /* (2, 12, 15) {real, imag} */,
  {32'hc547aad4, 32'h00000000} /* (2, 12, 14) {real, imag} */,
  {32'hc4f14c03, 32'h00000000} /* (2, 12, 13) {real, imag} */,
  {32'hc531a112, 32'h00000000} /* (2, 12, 12) {real, imag} */,
  {32'hc4bd71a3, 32'h00000000} /* (2, 12, 11) {real, imag} */,
  {32'h3fac7c00, 32'h00000000} /* (2, 12, 10) {real, imag} */,
  {32'h448aac32, 32'h00000000} /* (2, 12, 9) {real, imag} */,
  {32'h4510e812, 32'h00000000} /* (2, 12, 8) {real, imag} */,
  {32'h452a5829, 32'h00000000} /* (2, 12, 7) {real, imag} */,
  {32'h452c88d9, 32'h00000000} /* (2, 12, 6) {real, imag} */,
  {32'h452928cc, 32'h00000000} /* (2, 12, 5) {real, imag} */,
  {32'h45194c1c, 32'h00000000} /* (2, 12, 4) {real, imag} */,
  {32'h4549a7e8, 32'h00000000} /* (2, 12, 3) {real, imag} */,
  {32'h456562d1, 32'h00000000} /* (2, 12, 2) {real, imag} */,
  {32'h45558323, 32'h00000000} /* (2, 12, 1) {real, imag} */,
  {32'h45339fda, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h44e18e39, 32'h00000000} /* (2, 11, 31) {real, imag} */,
  {32'h45094f88, 32'h00000000} /* (2, 11, 30) {real, imag} */,
  {32'h452135e7, 32'h00000000} /* (2, 11, 29) {real, imag} */,
  {32'h45271903, 32'h00000000} /* (2, 11, 28) {real, imag} */,
  {32'h44cb145c, 32'h00000000} /* (2, 11, 27) {real, imag} */,
  {32'h449d1510, 32'h00000000} /* (2, 11, 26) {real, imag} */,
  {32'h4500a33b, 32'h00000000} /* (2, 11, 25) {real, imag} */,
  {32'h44dd8b29, 32'h00000000} /* (2, 11, 24) {real, imag} */,
  {32'h44a998b6, 32'h00000000} /* (2, 11, 23) {real, imag} */,
  {32'h4488881f, 32'h00000000} /* (2, 11, 22) {real, imag} */,
  {32'h43d6ccb0, 32'h00000000} /* (2, 11, 21) {real, imag} */,
  {32'hc4838d6a, 32'h00000000} /* (2, 11, 20) {real, imag} */,
  {32'hc4bc026c, 32'h00000000} /* (2, 11, 19) {real, imag} */,
  {32'hc4ece956, 32'h00000000} /* (2, 11, 18) {real, imag} */,
  {32'hc4e27fb8, 32'h00000000} /* (2, 11, 17) {real, imag} */,
  {32'hc51c3d93, 32'h00000000} /* (2, 11, 16) {real, imag} */,
  {32'hc5138504, 32'h00000000} /* (2, 11, 15) {real, imag} */,
  {32'hc514b980, 32'h00000000} /* (2, 11, 14) {real, imag} */,
  {32'hc51171cd, 32'h00000000} /* (2, 11, 13) {real, imag} */,
  {32'hc4fa2432, 32'h00000000} /* (2, 11, 12) {real, imag} */,
  {32'hc50f6b83, 32'h00000000} /* (2, 11, 11) {real, imag} */,
  {32'hc2a1e878, 32'h00000000} /* (2, 11, 10) {real, imag} */,
  {32'h44e94f96, 32'h00000000} /* (2, 11, 9) {real, imag} */,
  {32'h45167e22, 32'h00000000} /* (2, 11, 8) {real, imag} */,
  {32'h4525ce68, 32'h00000000} /* (2, 11, 7) {real, imag} */,
  {32'h451c832c, 32'h00000000} /* (2, 11, 6) {real, imag} */,
  {32'h44b65aea, 32'h00000000} /* (2, 11, 5) {real, imag} */,
  {32'h451f5d70, 32'h00000000} /* (2, 11, 4) {real, imag} */,
  {32'h4503314e, 32'h00000000} /* (2, 11, 3) {real, imag} */,
  {32'h44829cb2, 32'h00000000} /* (2, 11, 2) {real, imag} */,
  {32'h4500c23c, 32'h00000000} /* (2, 11, 1) {real, imag} */,
  {32'h44f834de, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'hc2e83c88, 32'h00000000} /* (2, 10, 31) {real, imag} */,
  {32'h42fd47be, 32'h00000000} /* (2, 10, 30) {real, imag} */,
  {32'h43d41f31, 32'h00000000} /* (2, 10, 29) {real, imag} */,
  {32'hc327de0e, 32'h00000000} /* (2, 10, 28) {real, imag} */,
  {32'h43b9021d, 32'h00000000} /* (2, 10, 27) {real, imag} */,
  {32'hc4bd87dc, 32'h00000000} /* (2, 10, 26) {real, imag} */,
  {32'hc470719b, 32'h00000000} /* (2, 10, 25) {real, imag} */,
  {32'hc3697a72, 32'h00000000} /* (2, 10, 24) {real, imag} */,
  {32'hc3e338ce, 32'h00000000} /* (2, 10, 23) {real, imag} */,
  {32'hc39e7516, 32'h00000000} /* (2, 10, 22) {real, imag} */,
  {32'hc211d3d0, 32'h00000000} /* (2, 10, 21) {real, imag} */,
  {32'h43ea2b2d, 32'h00000000} /* (2, 10, 20) {real, imag} */,
  {32'hc2894b20, 32'h00000000} /* (2, 10, 19) {real, imag} */,
  {32'h43c484e5, 32'h00000000} /* (2, 10, 18) {real, imag} */,
  {32'h4480c0e6, 32'h00000000} /* (2, 10, 17) {real, imag} */,
  {32'hc22d3e30, 32'h00000000} /* (2, 10, 16) {real, imag} */,
  {32'h43ec3060, 32'h00000000} /* (2, 10, 15) {real, imag} */,
  {32'h43900f72, 32'h00000000} /* (2, 10, 14) {real, imag} */,
  {32'h43ddb0bd, 32'h00000000} /* (2, 10, 13) {real, imag} */,
  {32'h42d44397, 32'h00000000} /* (2, 10, 12) {real, imag} */,
  {32'h43db5129, 32'h00000000} /* (2, 10, 11) {real, imag} */,
  {32'h4302ba68, 32'h00000000} /* (2, 10, 10) {real, imag} */,
  {32'h4377fbcc, 32'h00000000} /* (2, 10, 9) {real, imag} */,
  {32'hc41ccddc, 32'h00000000} /* (2, 10, 8) {real, imag} */,
  {32'h413c6900, 32'h00000000} /* (2, 10, 7) {real, imag} */,
  {32'hc281d35c, 32'h00000000} /* (2, 10, 6) {real, imag} */,
  {32'hc31c79a0, 32'h00000000} /* (2, 10, 5) {real, imag} */,
  {32'hc4193f7e, 32'h00000000} /* (2, 10, 4) {real, imag} */,
  {32'hc4b3bc96, 32'h00000000} /* (2, 10, 3) {real, imag} */,
  {32'hc4a702ef, 32'h00000000} /* (2, 10, 2) {real, imag} */,
  {32'hc522df3b, 32'h00000000} /* (2, 10, 1) {real, imag} */,
  {32'hc4546d78, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'hc50fd2b3, 32'h00000000} /* (2, 9, 31) {real, imag} */,
  {32'hc4f3ba53, 32'h00000000} /* (2, 9, 30) {real, imag} */,
  {32'hc48ee6cd, 32'h00000000} /* (2, 9, 29) {real, imag} */,
  {32'hc4d679ec, 32'h00000000} /* (2, 9, 28) {real, imag} */,
  {32'hc4e1cf5e, 32'h00000000} /* (2, 9, 27) {real, imag} */,
  {32'hc527cabd, 32'h00000000} /* (2, 9, 26) {real, imag} */,
  {32'hc5312a59, 32'h00000000} /* (2, 9, 25) {real, imag} */,
  {32'hc50c948a, 32'h00000000} /* (2, 9, 24) {real, imag} */,
  {32'hc4b1cf64, 32'h00000000} /* (2, 9, 23) {real, imag} */,
  {32'hc501496d, 32'h00000000} /* (2, 9, 22) {real, imag} */,
  {32'hc4811188, 32'h00000000} /* (2, 9, 21) {real, imag} */,
  {32'h44423e58, 32'h00000000} /* (2, 9, 20) {real, imag} */,
  {32'h44dbe522, 32'h00000000} /* (2, 9, 19) {real, imag} */,
  {32'h4489f88c, 32'h00000000} /* (2, 9, 18) {real, imag} */,
  {32'h448fbf0c, 32'h00000000} /* (2, 9, 17) {real, imag} */,
  {32'h44d0fd82, 32'h00000000} /* (2, 9, 16) {real, imag} */,
  {32'h4521d11f, 32'h00000000} /* (2, 9, 15) {real, imag} */,
  {32'h449aea77, 32'h00000000} /* (2, 9, 14) {real, imag} */,
  {32'h44ee00a7, 32'h00000000} /* (2, 9, 13) {real, imag} */,
  {32'h44d0441c, 32'h00000000} /* (2, 9, 12) {real, imag} */,
  {32'h44c00bcc, 32'h00000000} /* (2, 9, 11) {real, imag} */,
  {32'hc350f230, 32'h00000000} /* (2, 9, 10) {real, imag} */,
  {32'hc404012c, 32'h00000000} /* (2, 9, 9) {real, imag} */,
  {32'hc487b3cd, 32'h00000000} /* (2, 9, 8) {real, imag} */,
  {32'hc4865a94, 32'h00000000} /* (2, 9, 7) {real, imag} */,
  {32'hc4d6c3fe, 32'h00000000} /* (2, 9, 6) {real, imag} */,
  {32'hc503c97d, 32'h00000000} /* (2, 9, 5) {real, imag} */,
  {32'hc520a01e, 32'h00000000} /* (2, 9, 4) {real, imag} */,
  {32'hc557529f, 32'h00000000} /* (2, 9, 3) {real, imag} */,
  {32'hc54efd04, 32'h00000000} /* (2, 9, 2) {real, imag} */,
  {32'hc5049c5a, 32'h00000000} /* (2, 9, 1) {real, imag} */,
  {32'hc4befcfa, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'hc5344fa6, 32'h00000000} /* (2, 8, 31) {real, imag} */,
  {32'hc56b1e88, 32'h00000000} /* (2, 8, 30) {real, imag} */,
  {32'hc50fdd0a, 32'h00000000} /* (2, 8, 29) {real, imag} */,
  {32'hc53358ce, 32'h00000000} /* (2, 8, 28) {real, imag} */,
  {32'hc542539d, 32'h00000000} /* (2, 8, 27) {real, imag} */,
  {32'hc54e0d82, 32'h00000000} /* (2, 8, 26) {real, imag} */,
  {32'hc5476e28, 32'h00000000} /* (2, 8, 25) {real, imag} */,
  {32'hc52ca2da, 32'h00000000} /* (2, 8, 24) {real, imag} */,
  {32'hc536ac24, 32'h00000000} /* (2, 8, 23) {real, imag} */,
  {32'hc50af6d4, 32'h00000000} /* (2, 8, 22) {real, imag} */,
  {32'hc455558e, 32'h00000000} /* (2, 8, 21) {real, imag} */,
  {32'h441c35c6, 32'h00000000} /* (2, 8, 20) {real, imag} */,
  {32'h45339ffb, 32'h00000000} /* (2, 8, 19) {real, imag} */,
  {32'h45164fbf, 32'h00000000} /* (2, 8, 18) {real, imag} */,
  {32'h4516c00c, 32'h00000000} /* (2, 8, 17) {real, imag} */,
  {32'h4551effd, 32'h00000000} /* (2, 8, 16) {real, imag} */,
  {32'h450eb6c4, 32'h00000000} /* (2, 8, 15) {real, imag} */,
  {32'h4520a49c, 32'h00000000} /* (2, 8, 14) {real, imag} */,
  {32'h44e0933d, 32'h00000000} /* (2, 8, 13) {real, imag} */,
  {32'h44d7133b, 32'h00000000} /* (2, 8, 12) {real, imag} */,
  {32'h448fc446, 32'h00000000} /* (2, 8, 11) {real, imag} */,
  {32'hc42963fa, 32'h00000000} /* (2, 8, 10) {real, imag} */,
  {32'hc528d8e4, 32'h00000000} /* (2, 8, 9) {real, imag} */,
  {32'hc5141de0, 32'h00000000} /* (2, 8, 8) {real, imag} */,
  {32'hc507b598, 32'h00000000} /* (2, 8, 7) {real, imag} */,
  {32'hc510d442, 32'h00000000} /* (2, 8, 6) {real, imag} */,
  {32'hc518047c, 32'h00000000} /* (2, 8, 5) {real, imag} */,
  {32'hc53cf750, 32'h00000000} /* (2, 8, 4) {real, imag} */,
  {32'hc56fa2fd, 32'h00000000} /* (2, 8, 3) {real, imag} */,
  {32'hc534c3f1, 32'h00000000} /* (2, 8, 2) {real, imag} */,
  {32'hc4fa3aa9, 32'h00000000} /* (2, 8, 1) {real, imag} */,
  {32'hc4e2eb0e, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'hc4f74a9e, 32'h00000000} /* (2, 7, 31) {real, imag} */,
  {32'hc526fee4, 32'h00000000} /* (2, 7, 30) {real, imag} */,
  {32'hc58d8efd, 32'h00000000} /* (2, 7, 29) {real, imag} */,
  {32'hc571ab82, 32'h00000000} /* (2, 7, 28) {real, imag} */,
  {32'hc57bf252, 32'h00000000} /* (2, 7, 27) {real, imag} */,
  {32'hc591f5d8, 32'h00000000} /* (2, 7, 26) {real, imag} */,
  {32'hc583cc97, 32'h00000000} /* (2, 7, 25) {real, imag} */,
  {32'hc59e0168, 32'h00000000} /* (2, 7, 24) {real, imag} */,
  {32'hc53d35fe, 32'h00000000} /* (2, 7, 23) {real, imag} */,
  {32'hc4e8a097, 32'h00000000} /* (2, 7, 22) {real, imag} */,
  {32'hc4805fe6, 32'h00000000} /* (2, 7, 21) {real, imag} */,
  {32'h451aa899, 32'h00000000} /* (2, 7, 20) {real, imag} */,
  {32'h448423d7, 32'h00000000} /* (2, 7, 19) {real, imag} */,
  {32'h44ef369c, 32'h00000000} /* (2, 7, 18) {real, imag} */,
  {32'h4536282c, 32'h00000000} /* (2, 7, 17) {real, imag} */,
  {32'h45319618, 32'h00000000} /* (2, 7, 16) {real, imag} */,
  {32'h4574a379, 32'h00000000} /* (2, 7, 15) {real, imag} */,
  {32'h454ab5bc, 32'h00000000} /* (2, 7, 14) {real, imag} */,
  {32'h45172156, 32'h00000000} /* (2, 7, 13) {real, imag} */,
  {32'h44fccb5f, 32'h00000000} /* (2, 7, 12) {real, imag} */,
  {32'h444ad8a2, 32'h00000000} /* (2, 7, 11) {real, imag} */,
  {32'hc4384ae8, 32'h00000000} /* (2, 7, 10) {real, imag} */,
  {32'hc509774a, 32'h00000000} /* (2, 7, 9) {real, imag} */,
  {32'hc4bdfe68, 32'h00000000} /* (2, 7, 8) {real, imag} */,
  {32'hc51abf38, 32'h00000000} /* (2, 7, 7) {real, imag} */,
  {32'hc532f26c, 32'h00000000} /* (2, 7, 6) {real, imag} */,
  {32'hc52702fc, 32'h00000000} /* (2, 7, 5) {real, imag} */,
  {32'hc55059a9, 32'h00000000} /* (2, 7, 4) {real, imag} */,
  {32'hc575b88e, 32'h00000000} /* (2, 7, 3) {real, imag} */,
  {32'hc537f21e, 32'h00000000} /* (2, 7, 2) {real, imag} */,
  {32'hc56d4b38, 32'h00000000} /* (2, 7, 1) {real, imag} */,
  {32'hc51c6846, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'hc50c92d6, 32'h00000000} /* (2, 6, 31) {real, imag} */,
  {32'hc54ed665, 32'h00000000} /* (2, 6, 30) {real, imag} */,
  {32'hc57200ca, 32'h00000000} /* (2, 6, 29) {real, imag} */,
  {32'hc58ec36a, 32'h00000000} /* (2, 6, 28) {real, imag} */,
  {32'hc5a5e440, 32'h00000000} /* (2, 6, 27) {real, imag} */,
  {32'hc59beb6a, 32'h00000000} /* (2, 6, 26) {real, imag} */,
  {32'hc58d9e22, 32'h00000000} /* (2, 6, 25) {real, imag} */,
  {32'hc588b5de, 32'h00000000} /* (2, 6, 24) {real, imag} */,
  {32'hc538bcc0, 32'h00000000} /* (2, 6, 23) {real, imag} */,
  {32'hc4d54b7b, 32'h00000000} /* (2, 6, 22) {real, imag} */,
  {32'hc4840a5a, 32'h00000000} /* (2, 6, 21) {real, imag} */,
  {32'h44246ce4, 32'h00000000} /* (2, 6, 20) {real, imag} */,
  {32'h448ae35c, 32'h00000000} /* (2, 6, 19) {real, imag} */,
  {32'h446c98c8, 32'h00000000} /* (2, 6, 18) {real, imag} */,
  {32'h44da454a, 32'h00000000} /* (2, 6, 17) {real, imag} */,
  {32'h4539c436, 32'h00000000} /* (2, 6, 16) {real, imag} */,
  {32'h45192404, 32'h00000000} /* (2, 6, 15) {real, imag} */,
  {32'h4553739b, 32'h00000000} /* (2, 6, 14) {real, imag} */,
  {32'h4539904e, 32'h00000000} /* (2, 6, 13) {real, imag} */,
  {32'h4580d3fa, 32'h00000000} /* (2, 6, 12) {real, imag} */,
  {32'h451c6aff, 32'h00000000} /* (2, 6, 11) {real, imag} */,
  {32'h441bb080, 32'h00000000} /* (2, 6, 10) {real, imag} */,
  {32'hc40bd63c, 32'h00000000} /* (2, 6, 9) {real, imag} */,
  {32'hc4bc3812, 32'h00000000} /* (2, 6, 8) {real, imag} */,
  {32'hc4ba80b7, 32'h00000000} /* (2, 6, 7) {real, imag} */,
  {32'hc4c95345, 32'h00000000} /* (2, 6, 6) {real, imag} */,
  {32'hc50b2944, 32'h00000000} /* (2, 6, 5) {real, imag} */,
  {32'hc50e56a8, 32'h00000000} /* (2, 6, 4) {real, imag} */,
  {32'hc52deadc, 32'h00000000} /* (2, 6, 3) {real, imag} */,
  {32'hc5584936, 32'h00000000} /* (2, 6, 2) {real, imag} */,
  {32'hc5143057, 32'h00000000} /* (2, 6, 1) {real, imag} */,
  {32'hc4f9bcec, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hc552eb26, 32'h00000000} /* (2, 5, 31) {real, imag} */,
  {32'hc54012f6, 32'h00000000} /* (2, 5, 30) {real, imag} */,
  {32'hc5554260, 32'h00000000} /* (2, 5, 29) {real, imag} */,
  {32'hc5788827, 32'h00000000} /* (2, 5, 28) {real, imag} */,
  {32'hc59b8183, 32'h00000000} /* (2, 5, 27) {real, imag} */,
  {32'hc58951a6, 32'h00000000} /* (2, 5, 26) {real, imag} */,
  {32'hc5981a5a, 32'h00000000} /* (2, 5, 25) {real, imag} */,
  {32'hc574717e, 32'h00000000} /* (2, 5, 24) {real, imag} */,
  {32'hc54c3cf1, 32'h00000000} /* (2, 5, 23) {real, imag} */,
  {32'hc5171ead, 32'h00000000} /* (2, 5, 22) {real, imag} */,
  {32'hc484ee62, 32'h00000000} /* (2, 5, 21) {real, imag} */,
  {32'hc43f0dc3, 32'h00000000} /* (2, 5, 20) {real, imag} */,
  {32'hc3ab43d4, 32'h00000000} /* (2, 5, 19) {real, imag} */,
  {32'hc3d8b326, 32'h00000000} /* (2, 5, 18) {real, imag} */,
  {32'h43b332c4, 32'h00000000} /* (2, 5, 17) {real, imag} */,
  {32'hc3158a18, 32'h00000000} /* (2, 5, 16) {real, imag} */,
  {32'h44efeb18, 32'h00000000} /* (2, 5, 15) {real, imag} */,
  {32'h44f478ab, 32'h00000000} /* (2, 5, 14) {real, imag} */,
  {32'h45621892, 32'h00000000} /* (2, 5, 13) {real, imag} */,
  {32'h458f7b08, 32'h00000000} /* (2, 5, 12) {real, imag} */,
  {32'h455e02ce, 32'h00000000} /* (2, 5, 11) {real, imag} */,
  {32'h44e7096f, 32'h00000000} /* (2, 5, 10) {real, imag} */,
  {32'h44a2b21b, 32'h00000000} /* (2, 5, 9) {real, imag} */,
  {32'h4482ec95, 32'h00000000} /* (2, 5, 8) {real, imag} */,
  {32'h42b99320, 32'h00000000} /* (2, 5, 7) {real, imag} */,
  {32'hc3c00ba2, 32'h00000000} /* (2, 5, 6) {real, imag} */,
  {32'hc46fbf04, 32'h00000000} /* (2, 5, 5) {real, imag} */,
  {32'hc52492c5, 32'h00000000} /* (2, 5, 4) {real, imag} */,
  {32'hc51c69a2, 32'h00000000} /* (2, 5, 3) {real, imag} */,
  {32'hc50f9540, 32'h00000000} /* (2, 5, 2) {real, imag} */,
  {32'hc50f8934, 32'h00000000} /* (2, 5, 1) {real, imag} */,
  {32'hc5258a54, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hc5569172, 32'h00000000} /* (2, 4, 31) {real, imag} */,
  {32'hc59d3f2d, 32'h00000000} /* (2, 4, 30) {real, imag} */,
  {32'hc591073c, 32'h00000000} /* (2, 4, 29) {real, imag} */,
  {32'hc56105ce, 32'h00000000} /* (2, 4, 28) {real, imag} */,
  {32'hc597c86b, 32'h00000000} /* (2, 4, 27) {real, imag} */,
  {32'hc5af9e1c, 32'h00000000} /* (2, 4, 26) {real, imag} */,
  {32'hc595c3be, 32'h00000000} /* (2, 4, 25) {real, imag} */,
  {32'hc58915ce, 32'h00000000} /* (2, 4, 24) {real, imag} */,
  {32'hc54a9a0c, 32'h00000000} /* (2, 4, 23) {real, imag} */,
  {32'hc529ceab, 32'h00000000} /* (2, 4, 22) {real, imag} */,
  {32'hc5315194, 32'h00000000} /* (2, 4, 21) {real, imag} */,
  {32'hc5374afc, 32'h00000000} /* (2, 4, 20) {real, imag} */,
  {32'hc4b7332a, 32'h00000000} /* (2, 4, 19) {real, imag} */,
  {32'hc4cf09e6, 32'h00000000} /* (2, 4, 18) {real, imag} */,
  {32'hc4a081bf, 32'h00000000} /* (2, 4, 17) {real, imag} */,
  {32'hc4bbd3fe, 32'h00000000} /* (2, 4, 16) {real, imag} */,
  {32'h44ff3cd5, 32'h00000000} /* (2, 4, 15) {real, imag} */,
  {32'h451454a0, 32'h00000000} /* (2, 4, 14) {real, imag} */,
  {32'h453f28c5, 32'h00000000} /* (2, 4, 13) {real, imag} */,
  {32'h457280aa, 32'h00000000} /* (2, 4, 12) {real, imag} */,
  {32'h4565763e, 32'h00000000} /* (2, 4, 11) {real, imag} */,
  {32'h4580a202, 32'h00000000} /* (2, 4, 10) {real, imag} */,
  {32'h454fdd5b, 32'h00000000} /* (2, 4, 9) {real, imag} */,
  {32'h45300104, 32'h00000000} /* (2, 4, 8) {real, imag} */,
  {32'h45177156, 32'h00000000} /* (2, 4, 7) {real, imag} */,
  {32'h44c1fd22, 32'h00000000} /* (2, 4, 6) {real, imag} */,
  {32'h432bb718, 32'h00000000} /* (2, 4, 5) {real, imag} */,
  {32'hc4a226e5, 32'h00000000} /* (2, 4, 4) {real, imag} */,
  {32'hc507ddc9, 32'h00000000} /* (2, 4, 3) {real, imag} */,
  {32'hc51563bd, 32'h00000000} /* (2, 4, 2) {real, imag} */,
  {32'hc536b1c6, 32'h00000000} /* (2, 4, 1) {real, imag} */,
  {32'hc527c3af, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hc53944a6, 32'h00000000} /* (2, 3, 31) {real, imag} */,
  {32'hc58f3c68, 32'h00000000} /* (2, 3, 30) {real, imag} */,
  {32'hc5707c31, 32'h00000000} /* (2, 3, 29) {real, imag} */,
  {32'hc561173a, 32'h00000000} /* (2, 3, 28) {real, imag} */,
  {32'hc5884c91, 32'h00000000} /* (2, 3, 27) {real, imag} */,
  {32'hc5865a33, 32'h00000000} /* (2, 3, 26) {real, imag} */,
  {32'hc5775f8f, 32'h00000000} /* (2, 3, 25) {real, imag} */,
  {32'hc560f3e1, 32'h00000000} /* (2, 3, 24) {real, imag} */,
  {32'hc5488336, 32'h00000000} /* (2, 3, 23) {real, imag} */,
  {32'hc5312cb8, 32'h00000000} /* (2, 3, 22) {real, imag} */,
  {32'hc51ccf2d, 32'h00000000} /* (2, 3, 21) {real, imag} */,
  {32'hc529f3a9, 32'h00000000} /* (2, 3, 20) {real, imag} */,
  {32'hc5416957, 32'h00000000} /* (2, 3, 19) {real, imag} */,
  {32'hc4c1dbbe, 32'h00000000} /* (2, 3, 18) {real, imag} */,
  {32'hc50333ef, 32'h00000000} /* (2, 3, 17) {real, imag} */,
  {32'hc4ab3bb3, 32'h00000000} /* (2, 3, 16) {real, imag} */,
  {32'h44895f20, 32'h00000000} /* (2, 3, 15) {real, imag} */,
  {32'h453bbea6, 32'h00000000} /* (2, 3, 14) {real, imag} */,
  {32'h455ad853, 32'h00000000} /* (2, 3, 13) {real, imag} */,
  {32'h457480d6, 32'h00000000} /* (2, 3, 12) {real, imag} */,
  {32'h45960667, 32'h00000000} /* (2, 3, 11) {real, imag} */,
  {32'h45811747, 32'h00000000} /* (2, 3, 10) {real, imag} */,
  {32'h454b38c7, 32'h00000000} /* (2, 3, 9) {real, imag} */,
  {32'h45469d29, 32'h00000000} /* (2, 3, 8) {real, imag} */,
  {32'h453a7b08, 32'h00000000} /* (2, 3, 7) {real, imag} */,
  {32'h450be784, 32'h00000000} /* (2, 3, 6) {real, imag} */,
  {32'hc413d7e4, 32'h00000000} /* (2, 3, 5) {real, imag} */,
  {32'hc4a9f5c6, 32'h00000000} /* (2, 3, 4) {real, imag} */,
  {32'hc523a55d, 32'h00000000} /* (2, 3, 3) {real, imag} */,
  {32'hc52c0cb9, 32'h00000000} /* (2, 3, 2) {real, imag} */,
  {32'hc5282e49, 32'h00000000} /* (2, 3, 1) {real, imag} */,
  {32'hc50ad300, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hc50d2dff, 32'h00000000} /* (2, 2, 31) {real, imag} */,
  {32'hc53b0b14, 32'h00000000} /* (2, 2, 30) {real, imag} */,
  {32'hc565ffd6, 32'h00000000} /* (2, 2, 29) {real, imag} */,
  {32'hc55d1f56, 32'h00000000} /* (2, 2, 28) {real, imag} */,
  {32'hc55b51fc, 32'h00000000} /* (2, 2, 27) {real, imag} */,
  {32'hc5560733, 32'h00000000} /* (2, 2, 26) {real, imag} */,
  {32'hc5747e10, 32'h00000000} /* (2, 2, 25) {real, imag} */,
  {32'hc53ea21c, 32'h00000000} /* (2, 2, 24) {real, imag} */,
  {32'hc515dd53, 32'h00000000} /* (2, 2, 23) {real, imag} */,
  {32'hc519dabb, 32'h00000000} /* (2, 2, 22) {real, imag} */,
  {32'hc553c1a8, 32'h00000000} /* (2, 2, 21) {real, imag} */,
  {32'hc57b48fb, 32'h00000000} /* (2, 2, 20) {real, imag} */,
  {32'hc564bd5c, 32'h00000000} /* (2, 2, 19) {real, imag} */,
  {32'hc5342ea6, 32'h00000000} /* (2, 2, 18) {real, imag} */,
  {32'hc51c8aec, 32'h00000000} /* (2, 2, 17) {real, imag} */,
  {32'hc3af3120, 32'h00000000} /* (2, 2, 16) {real, imag} */,
  {32'h45015785, 32'h00000000} /* (2, 2, 15) {real, imag} */,
  {32'h4540decc, 32'h00000000} /* (2, 2, 14) {real, imag} */,
  {32'h4584ebb5, 32'h00000000} /* (2, 2, 13) {real, imag} */,
  {32'h4576b252, 32'h00000000} /* (2, 2, 12) {real, imag} */,
  {32'h459f4a7a, 32'h00000000} /* (2, 2, 11) {real, imag} */,
  {32'h45605355, 32'h00000000} /* (2, 2, 10) {real, imag} */,
  {32'h45855f1e, 32'h00000000} /* (2, 2, 9) {real, imag} */,
  {32'h454f2d90, 32'h00000000} /* (2, 2, 8) {real, imag} */,
  {32'h452bee09, 32'h00000000} /* (2, 2, 7) {real, imag} */,
  {32'h44d19a9a, 32'h00000000} /* (2, 2, 6) {real, imag} */,
  {32'hc465c660, 32'h00000000} /* (2, 2, 5) {real, imag} */,
  {32'hc5064eb3, 32'h00000000} /* (2, 2, 4) {real, imag} */,
  {32'hc5695394, 32'h00000000} /* (2, 2, 3) {real, imag} */,
  {32'hc527b27c, 32'h00000000} /* (2, 2, 2) {real, imag} */,
  {32'hc5648eba, 32'h00000000} /* (2, 2, 1) {real, imag} */,
  {32'hc510bcf4, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hc5126efc, 32'h00000000} /* (2, 1, 31) {real, imag} */,
  {32'hc522f07c, 32'h00000000} /* (2, 1, 30) {real, imag} */,
  {32'hc50bca10, 32'h00000000} /* (2, 1, 29) {real, imag} */,
  {32'hc527a7b6, 32'h00000000} /* (2, 1, 28) {real, imag} */,
  {32'hc52a62e2, 32'h00000000} /* (2, 1, 27) {real, imag} */,
  {32'hc550f52b, 32'h00000000} /* (2, 1, 26) {real, imag} */,
  {32'hc53be200, 32'h00000000} /* (2, 1, 25) {real, imag} */,
  {32'hc51c3b9d, 32'h00000000} /* (2, 1, 24) {real, imag} */,
  {32'hc50929b4, 32'h00000000} /* (2, 1, 23) {real, imag} */,
  {32'hc516a187, 32'h00000000} /* (2, 1, 22) {real, imag} */,
  {32'hc4e02049, 32'h00000000} /* (2, 1, 21) {real, imag} */,
  {32'hc50fdc58, 32'h00000000} /* (2, 1, 20) {real, imag} */,
  {32'hc5119833, 32'h00000000} /* (2, 1, 19) {real, imag} */,
  {32'hc5156ad0, 32'h00000000} /* (2, 1, 18) {real, imag} */,
  {32'hc445e3ce, 32'h00000000} /* (2, 1, 17) {real, imag} */,
  {32'h43c5e7a0, 32'h00000000} /* (2, 1, 16) {real, imag} */,
  {32'h451554ec, 32'h00000000} /* (2, 1, 15) {real, imag} */,
  {32'h4554ce24, 32'h00000000} /* (2, 1, 14) {real, imag} */,
  {32'h45813692, 32'h00000000} /* (2, 1, 13) {real, imag} */,
  {32'h458ebe64, 32'h00000000} /* (2, 1, 12) {real, imag} */,
  {32'h4581de41, 32'h00000000} /* (2, 1, 11) {real, imag} */,
  {32'h4568b7af, 32'h00000000} /* (2, 1, 10) {real, imag} */,
  {32'h457fda58, 32'h00000000} /* (2, 1, 9) {real, imag} */,
  {32'h4534d429, 32'h00000000} /* (2, 1, 8) {real, imag} */,
  {32'h450c5172, 32'h00000000} /* (2, 1, 7) {real, imag} */,
  {32'h452f1b43, 32'h00000000} /* (2, 1, 6) {real, imag} */,
  {32'hc3240c08, 32'h00000000} /* (2, 1, 5) {real, imag} */,
  {32'hc5392aca, 32'h00000000} /* (2, 1, 4) {real, imag} */,
  {32'hc50bfdc1, 32'h00000000} /* (2, 1, 3) {real, imag} */,
  {32'hc50daa9e, 32'h00000000} /* (2, 1, 2) {real, imag} */,
  {32'hc546a186, 32'h00000000} /* (2, 1, 1) {real, imag} */,
  {32'hc51c5017, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hc4d594c2, 32'h00000000} /* (2, 0, 31) {real, imag} */,
  {32'hc4ede7ff, 32'h00000000} /* (2, 0, 30) {real, imag} */,
  {32'hc4dad4f0, 32'h00000000} /* (2, 0, 29) {real, imag} */,
  {32'hc50b2c94, 32'h00000000} /* (2, 0, 28) {real, imag} */,
  {32'hc50901c0, 32'h00000000} /* (2, 0, 27) {real, imag} */,
  {32'hc507330f, 32'h00000000} /* (2, 0, 26) {real, imag} */,
  {32'hc500c56e, 32'h00000000} /* (2, 0, 25) {real, imag} */,
  {32'hc5091859, 32'h00000000} /* (2, 0, 24) {real, imag} */,
  {32'hc52e0a0a, 32'h00000000} /* (2, 0, 23) {real, imag} */,
  {32'hc4ed629e, 32'h00000000} /* (2, 0, 22) {real, imag} */,
  {32'hc44551c5, 32'h00000000} /* (2, 0, 21) {real, imag} */,
  {32'hc4851d6e, 32'h00000000} /* (2, 0, 20) {real, imag} */,
  {32'hc429cb14, 32'h00000000} /* (2, 0, 19) {real, imag} */,
  {32'hc430a016, 32'h00000000} /* (2, 0, 18) {real, imag} */,
  {32'h423e54a0, 32'h00000000} /* (2, 0, 17) {real, imag} */,
  {32'h449530ad, 32'h00000000} /* (2, 0, 16) {real, imag} */,
  {32'h44fad60c, 32'h00000000} /* (2, 0, 15) {real, imag} */,
  {32'h451a3060, 32'h00000000} /* (2, 0, 14) {real, imag} */,
  {32'h4556a3be, 32'h00000000} /* (2, 0, 13) {real, imag} */,
  {32'h45621a8e, 32'h00000000} /* (2, 0, 12) {real, imag} */,
  {32'h4523b15c, 32'h00000000} /* (2, 0, 11) {real, imag} */,
  {32'h45297d0b, 32'h00000000} /* (2, 0, 10) {real, imag} */,
  {32'h4505bf90, 32'h00000000} /* (2, 0, 9) {real, imag} */,
  {32'h4494b6a0, 32'h00000000} /* (2, 0, 8) {real, imag} */,
  {32'h44a85eb7, 32'h00000000} /* (2, 0, 7) {real, imag} */,
  {32'h45180371, 32'h00000000} /* (2, 0, 6) {real, imag} */,
  {32'hc42e55e1, 32'h00000000} /* (2, 0, 5) {real, imag} */,
  {32'hc50c7bcc, 32'h00000000} /* (2, 0, 4) {real, imag} */,
  {32'hc4e21904, 32'h00000000} /* (2, 0, 3) {real, imag} */,
  {32'hc517ba26, 32'h00000000} /* (2, 0, 2) {real, imag} */,
  {32'hc50c5fac, 32'h00000000} /* (2, 0, 1) {real, imag} */,
  {32'hc505ccc4, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc4a517f9, 32'h00000000} /* (1, 31, 31) {real, imag} */,
  {32'hc4f75d18, 32'h00000000} /* (1, 31, 30) {real, imag} */,
  {32'hc4fb43f6, 32'h00000000} /* (1, 31, 29) {real, imag} */,
  {32'hc5378e8e, 32'h00000000} /* (1, 31, 28) {real, imag} */,
  {32'hc510c6e1, 32'h00000000} /* (1, 31, 27) {real, imag} */,
  {32'hc4d801c0, 32'h00000000} /* (1, 31, 26) {real, imag} */,
  {32'hc4d1476b, 32'h00000000} /* (1, 31, 25) {real, imag} */,
  {32'hc50a8985, 32'h00000000} /* (1, 31, 24) {real, imag} */,
  {32'hc4dcdd64, 32'h00000000} /* (1, 31, 23) {real, imag} */,
  {32'hc4e14056, 32'h00000000} /* (1, 31, 22) {real, imag} */,
  {32'hc4a0b25d, 32'h00000000} /* (1, 31, 21) {real, imag} */,
  {32'h430ff718, 32'h00000000} /* (1, 31, 20) {real, imag} */,
  {32'h44784a07, 32'h00000000} /* (1, 31, 19) {real, imag} */,
  {32'h44a5053d, 32'h00000000} /* (1, 31, 18) {real, imag} */,
  {32'h441c4f2e, 32'h00000000} /* (1, 31, 17) {real, imag} */,
  {32'h44c0e8ba, 32'h00000000} /* (1, 31, 16) {real, imag} */,
  {32'h450a8b8a, 32'h00000000} /* (1, 31, 15) {real, imag} */,
  {32'h45261834, 32'h00000000} /* (1, 31, 14) {real, imag} */,
  {32'h450c7213, 32'h00000000} /* (1, 31, 13) {real, imag} */,
  {32'h4500c502, 32'h00000000} /* (1, 31, 12) {real, imag} */,
  {32'h44f6423e, 32'h00000000} /* (1, 31, 11) {real, imag} */,
  {32'h44053b57, 32'h00000000} /* (1, 31, 10) {real, imag} */,
  {32'h425d6960, 32'h00000000} /* (1, 31, 9) {real, imag} */,
  {32'hc372a410, 32'h00000000} /* (1, 31, 8) {real, imag} */,
  {32'hc46258c8, 32'h00000000} /* (1, 31, 7) {real, imag} */,
  {32'hc4374433, 32'h00000000} /* (1, 31, 6) {real, imag} */,
  {32'hc4e904db, 32'h00000000} /* (1, 31, 5) {real, imag} */,
  {32'hc4f9d133, 32'h00000000} /* (1, 31, 4) {real, imag} */,
  {32'hc4b79d40, 32'h00000000} /* (1, 31, 3) {real, imag} */,
  {32'hc4e79fe5, 32'h00000000} /* (1, 31, 2) {real, imag} */,
  {32'hc4e344f1, 32'h00000000} /* (1, 31, 1) {real, imag} */,
  {32'hc48fff5a, 32'h00000000} /* (1, 31, 0) {real, imag} */,
  {32'hc499a0b4, 32'h00000000} /* (1, 30, 31) {real, imag} */,
  {32'hc4964fa0, 32'h00000000} /* (1, 30, 30) {real, imag} */,
  {32'hc50183f4, 32'h00000000} /* (1, 30, 29) {real, imag} */,
  {32'hc56c39a6, 32'h00000000} /* (1, 30, 28) {real, imag} */,
  {32'hc524f954, 32'h00000000} /* (1, 30, 27) {real, imag} */,
  {32'hc4febc00, 32'h00000000} /* (1, 30, 26) {real, imag} */,
  {32'hc501fbe0, 32'h00000000} /* (1, 30, 25) {real, imag} */,
  {32'hc4dfd902, 32'h00000000} /* (1, 30, 24) {real, imag} */,
  {32'hc4e6521e, 32'h00000000} /* (1, 30, 23) {real, imag} */,
  {32'hc5011a06, 32'h00000000} /* (1, 30, 22) {real, imag} */,
  {32'hc489385e, 32'h00000000} /* (1, 30, 21) {real, imag} */,
  {32'h44cba70e, 32'h00000000} /* (1, 30, 20) {real, imag} */,
  {32'h449a5d98, 32'h00000000} /* (1, 30, 19) {real, imag} */,
  {32'h44e88850, 32'h00000000} /* (1, 30, 18) {real, imag} */,
  {32'h44fe3412, 32'h00000000} /* (1, 30, 17) {real, imag} */,
  {32'h4542d77e, 32'h00000000} /* (1, 30, 16) {real, imag} */,
  {32'h4532c3be, 32'h00000000} /* (1, 30, 15) {real, imag} */,
  {32'h4517aa84, 32'h00000000} /* (1, 30, 14) {real, imag} */,
  {32'h44f77a8f, 32'h00000000} /* (1, 30, 13) {real, imag} */,
  {32'h44e2e830, 32'h00000000} /* (1, 30, 12) {real, imag} */,
  {32'h44f98fe7, 32'h00000000} /* (1, 30, 11) {real, imag} */,
  {32'h43cea880, 32'h00000000} /* (1, 30, 10) {real, imag} */,
  {32'hc4a597c0, 32'h00000000} /* (1, 30, 9) {real, imag} */,
  {32'hc4a637fc, 32'h00000000} /* (1, 30, 8) {real, imag} */,
  {32'hc5002403, 32'h00000000} /* (1, 30, 7) {real, imag} */,
  {32'hc52410ec, 32'h00000000} /* (1, 30, 6) {real, imag} */,
  {32'hc5128e5f, 32'h00000000} /* (1, 30, 5) {real, imag} */,
  {32'hc51b97c1, 32'h00000000} /* (1, 30, 4) {real, imag} */,
  {32'hc537886e, 32'h00000000} /* (1, 30, 3) {real, imag} */,
  {32'hc50c8734, 32'h00000000} /* (1, 30, 2) {real, imag} */,
  {32'hc4a6610a, 32'h00000000} /* (1, 30, 1) {real, imag} */,
  {32'hc4da3f9b, 32'h00000000} /* (1, 30, 0) {real, imag} */,
  {32'hc4de571a, 32'h00000000} /* (1, 29, 31) {real, imag} */,
  {32'hc4ff565a, 32'h00000000} /* (1, 29, 30) {real, imag} */,
  {32'hc53951dc, 32'h00000000} /* (1, 29, 29) {real, imag} */,
  {32'hc5354b62, 32'h00000000} /* (1, 29, 28) {real, imag} */,
  {32'hc511a9e0, 32'h00000000} /* (1, 29, 27) {real, imag} */,
  {32'hc5184c7c, 32'h00000000} /* (1, 29, 26) {real, imag} */,
  {32'hc50ea5e6, 32'h00000000} /* (1, 29, 25) {real, imag} */,
  {32'hc4f06c27, 32'h00000000} /* (1, 29, 24) {real, imag} */,
  {32'hc51cc06e, 32'h00000000} /* (1, 29, 23) {real, imag} */,
  {32'hc519fa6e, 32'h00000000} /* (1, 29, 22) {real, imag} */,
  {32'hc3883ce0, 32'h00000000} /* (1, 29, 21) {real, imag} */,
  {32'h44edaf6e, 32'h00000000} /* (1, 29, 20) {real, imag} */,
  {32'h45102550, 32'h00000000} /* (1, 29, 19) {real, imag} */,
  {32'h45226132, 32'h00000000} /* (1, 29, 18) {real, imag} */,
  {32'h454b181d, 32'h00000000} /* (1, 29, 17) {real, imag} */,
  {32'h454481c6, 32'h00000000} /* (1, 29, 16) {real, imag} */,
  {32'h453fe781, 32'h00000000} /* (1, 29, 15) {real, imag} */,
  {32'h4553246b, 32'h00000000} /* (1, 29, 14) {real, imag} */,
  {32'h451fbb6c, 32'h00000000} /* (1, 29, 13) {real, imag} */,
  {32'h4501a0bc, 32'h00000000} /* (1, 29, 12) {real, imag} */,
  {32'h44ae4469, 32'h00000000} /* (1, 29, 11) {real, imag} */,
  {32'hc4426549, 32'h00000000} /* (1, 29, 10) {real, imag} */,
  {32'hc50447bc, 32'h00000000} /* (1, 29, 9) {real, imag} */,
  {32'hc51714e9, 32'h00000000} /* (1, 29, 8) {real, imag} */,
  {32'hc507aec6, 32'h00000000} /* (1, 29, 7) {real, imag} */,
  {32'hc51f0e30, 32'h00000000} /* (1, 29, 6) {real, imag} */,
  {32'hc55cfb3d, 32'h00000000} /* (1, 29, 5) {real, imag} */,
  {32'hc587d03e, 32'h00000000} /* (1, 29, 4) {real, imag} */,
  {32'hc551ef90, 32'h00000000} /* (1, 29, 3) {real, imag} */,
  {32'hc5263dea, 32'h00000000} /* (1, 29, 2) {real, imag} */,
  {32'hc4ffe572, 32'h00000000} /* (1, 29, 1) {real, imag} */,
  {32'hc4ccbc3f, 32'h00000000} /* (1, 29, 0) {real, imag} */,
  {32'hc50856c2, 32'h00000000} /* (1, 28, 31) {real, imag} */,
  {32'hc5420114, 32'h00000000} /* (1, 28, 30) {real, imag} */,
  {32'hc567c42e, 32'h00000000} /* (1, 28, 29) {real, imag} */,
  {32'hc5197ed1, 32'h00000000} /* (1, 28, 28) {real, imag} */,
  {32'hc526042c, 32'h00000000} /* (1, 28, 27) {real, imag} */,
  {32'hc5573ad4, 32'h00000000} /* (1, 28, 26) {real, imag} */,
  {32'hc52eb319, 32'h00000000} /* (1, 28, 25) {real, imag} */,
  {32'hc51f7fc7, 32'h00000000} /* (1, 28, 24) {real, imag} */,
  {32'hc5164886, 32'h00000000} /* (1, 28, 23) {real, imag} */,
  {32'hc4f4837c, 32'h00000000} /* (1, 28, 22) {real, imag} */,
  {32'hc406ca90, 32'h00000000} /* (1, 28, 21) {real, imag} */,
  {32'h4505d297, 32'h00000000} /* (1, 28, 20) {real, imag} */,
  {32'h456ae308, 32'h00000000} /* (1, 28, 19) {real, imag} */,
  {32'h454893a8, 32'h00000000} /* (1, 28, 18) {real, imag} */,
  {32'h4547d10c, 32'h00000000} /* (1, 28, 17) {real, imag} */,
  {32'h454b26cd, 32'h00000000} /* (1, 28, 16) {real, imag} */,
  {32'h4538ce4c, 32'h00000000} /* (1, 28, 15) {real, imag} */,
  {32'h452c3854, 32'h00000000} /* (1, 28, 14) {real, imag} */,
  {32'h452ce30c, 32'h00000000} /* (1, 28, 13) {real, imag} */,
  {32'h452e42c7, 32'h00000000} /* (1, 28, 12) {real, imag} */,
  {32'h44c1d03f, 32'h00000000} /* (1, 28, 11) {real, imag} */,
  {32'hc4685b62, 32'h00000000} /* (1, 28, 10) {real, imag} */,
  {32'hc4c95342, 32'h00000000} /* (1, 28, 9) {real, imag} */,
  {32'hc4f55e06, 32'h00000000} /* (1, 28, 8) {real, imag} */,
  {32'hc53e4d8e, 32'h00000000} /* (1, 28, 7) {real, imag} */,
  {32'hc516405e, 32'h00000000} /* (1, 28, 6) {real, imag} */,
  {32'hc52de692, 32'h00000000} /* (1, 28, 5) {real, imag} */,
  {32'hc5423935, 32'h00000000} /* (1, 28, 4) {real, imag} */,
  {32'hc53083ae, 32'h00000000} /* (1, 28, 3) {real, imag} */,
  {32'hc514a10e, 32'h00000000} /* (1, 28, 2) {real, imag} */,
  {32'hc516ede0, 32'h00000000} /* (1, 28, 1) {real, imag} */,
  {32'hc51a42d5, 32'h00000000} /* (1, 28, 0) {real, imag} */,
  {32'hc4f2137e, 32'h00000000} /* (1, 27, 31) {real, imag} */,
  {32'hc5503fa8, 32'h00000000} /* (1, 27, 30) {real, imag} */,
  {32'hc58b5f89, 32'h00000000} /* (1, 27, 29) {real, imag} */,
  {32'hc562eb52, 32'h00000000} /* (1, 27, 28) {real, imag} */,
  {32'hc5188977, 32'h00000000} /* (1, 27, 27) {real, imag} */,
  {32'hc500cd71, 32'h00000000} /* (1, 27, 26) {real, imag} */,
  {32'hc5360d6f, 32'h00000000} /* (1, 27, 25) {real, imag} */,
  {32'hc4ff94dc, 32'h00000000} /* (1, 27, 24) {real, imag} */,
  {32'hc52d73e6, 32'h00000000} /* (1, 27, 23) {real, imag} */,
  {32'hc49708dc, 32'h00000000} /* (1, 27, 22) {real, imag} */,
  {32'h433227a8, 32'h00000000} /* (1, 27, 21) {real, imag} */,
  {32'h454c07c3, 32'h00000000} /* (1, 27, 20) {real, imag} */,
  {32'h457d99a8, 32'h00000000} /* (1, 27, 19) {real, imag} */,
  {32'h4574b494, 32'h00000000} /* (1, 27, 18) {real, imag} */,
  {32'h455faeaa, 32'h00000000} /* (1, 27, 17) {real, imag} */,
  {32'h454d513c, 32'h00000000} /* (1, 27, 16) {real, imag} */,
  {32'h454a090f, 32'h00000000} /* (1, 27, 15) {real, imag} */,
  {32'h4542cac8, 32'h00000000} /* (1, 27, 14) {real, imag} */,
  {32'h45304691, 32'h00000000} /* (1, 27, 13) {real, imag} */,
  {32'h4522b7c4, 32'h00000000} /* (1, 27, 12) {real, imag} */,
  {32'h44e1fea1, 32'h00000000} /* (1, 27, 11) {real, imag} */,
  {32'hc25ed5c0, 32'h00000000} /* (1, 27, 10) {real, imag} */,
  {32'hc47bcfd7, 32'h00000000} /* (1, 27, 9) {real, imag} */,
  {32'hc50806ee, 32'h00000000} /* (1, 27, 8) {real, imag} */,
  {32'hc516404c, 32'h00000000} /* (1, 27, 7) {real, imag} */,
  {32'hc502b35a, 32'h00000000} /* (1, 27, 6) {real, imag} */,
  {32'hc53805de, 32'h00000000} /* (1, 27, 5) {real, imag} */,
  {32'hc51e3d3f, 32'h00000000} /* (1, 27, 4) {real, imag} */,
  {32'hc53180b0, 32'h00000000} /* (1, 27, 3) {real, imag} */,
  {32'hc54c6c84, 32'h00000000} /* (1, 27, 2) {real, imag} */,
  {32'hc516605a, 32'h00000000} /* (1, 27, 1) {real, imag} */,
  {32'hc4fa1a79, 32'h00000000} /* (1, 27, 0) {real, imag} */,
  {32'hc50ffd48, 32'h00000000} /* (1, 26, 31) {real, imag} */,
  {32'hc559403f, 32'h00000000} /* (1, 26, 30) {real, imag} */,
  {32'hc56c9cf1, 32'h00000000} /* (1, 26, 29) {real, imag} */,
  {32'hc52fc45e, 32'h00000000} /* (1, 26, 28) {real, imag} */,
  {32'hc518d37f, 32'h00000000} /* (1, 26, 27) {real, imag} */,
  {32'hc524120d, 32'h00000000} /* (1, 26, 26) {real, imag} */,
  {32'hc519ceb0, 32'h00000000} /* (1, 26, 25) {real, imag} */,
  {32'hc51152ed, 32'h00000000} /* (1, 26, 24) {real, imag} */,
  {32'hc4fa12d0, 32'h00000000} /* (1, 26, 23) {real, imag} */,
  {32'hc4b1d6e8, 32'h00000000} /* (1, 26, 22) {real, imag} */,
  {32'h43c49172, 32'h00000000} /* (1, 26, 21) {real, imag} */,
  {32'h44f0dc0b, 32'h00000000} /* (1, 26, 20) {real, imag} */,
  {32'h454eb691, 32'h00000000} /* (1, 26, 19) {real, imag} */,
  {32'h4546670c, 32'h00000000} /* (1, 26, 18) {real, imag} */,
  {32'h456c9b62, 32'h00000000} /* (1, 26, 17) {real, imag} */,
  {32'h45616df4, 32'h00000000} /* (1, 26, 16) {real, imag} */,
  {32'h4524412a, 32'h00000000} /* (1, 26, 15) {real, imag} */,
  {32'h452ae5e3, 32'h00000000} /* (1, 26, 14) {real, imag} */,
  {32'h45156b35, 32'h00000000} /* (1, 26, 13) {real, imag} */,
  {32'h4506ae3a, 32'h00000000} /* (1, 26, 12) {real, imag} */,
  {32'h44f0847e, 32'h00000000} /* (1, 26, 11) {real, imag} */,
  {32'h43396980, 32'h00000000} /* (1, 26, 10) {real, imag} */,
  {32'hc50ea2d0, 32'h00000000} /* (1, 26, 9) {real, imag} */,
  {32'hc5078ef5, 32'h00000000} /* (1, 26, 8) {real, imag} */,
  {32'hc4ae9cce, 32'h00000000} /* (1, 26, 7) {real, imag} */,
  {32'hc50cddd2, 32'h00000000} /* (1, 26, 6) {real, imag} */,
  {32'hc511dffc, 32'h00000000} /* (1, 26, 5) {real, imag} */,
  {32'hc5371ec0, 32'h00000000} /* (1, 26, 4) {real, imag} */,
  {32'hc54a6e5f, 32'h00000000} /* (1, 26, 3) {real, imag} */,
  {32'hc56bb262, 32'h00000000} /* (1, 26, 2) {real, imag} */,
  {32'hc54b295c, 32'h00000000} /* (1, 26, 1) {real, imag} */,
  {32'hc5206246, 32'h00000000} /* (1, 26, 0) {real, imag} */,
  {32'hc530386c, 32'h00000000} /* (1, 25, 31) {real, imag} */,
  {32'hc55544d0, 32'h00000000} /* (1, 25, 30) {real, imag} */,
  {32'hc55387d1, 32'h00000000} /* (1, 25, 29) {real, imag} */,
  {32'hc5272e46, 32'h00000000} /* (1, 25, 28) {real, imag} */,
  {32'hc536792f, 32'h00000000} /* (1, 25, 27) {real, imag} */,
  {32'hc5385f00, 32'h00000000} /* (1, 25, 26) {real, imag} */,
  {32'hc5364302, 32'h00000000} /* (1, 25, 25) {real, imag} */,
  {32'hc50c0a24, 32'h00000000} /* (1, 25, 24) {real, imag} */,
  {32'hc4d8a7a0, 32'h00000000} /* (1, 25, 23) {real, imag} */,
  {32'hc4718a2c, 32'h00000000} /* (1, 25, 22) {real, imag} */,
  {32'h443b096b, 32'h00000000} /* (1, 25, 21) {real, imag} */,
  {32'h4558eeb5, 32'h00000000} /* (1, 25, 20) {real, imag} */,
  {32'h457deb22, 32'h00000000} /* (1, 25, 19) {real, imag} */,
  {32'h45633a92, 32'h00000000} /* (1, 25, 18) {real, imag} */,
  {32'h45374d79, 32'h00000000} /* (1, 25, 17) {real, imag} */,
  {32'h454da442, 32'h00000000} /* (1, 25, 16) {real, imag} */,
  {32'h45619cc8, 32'h00000000} /* (1, 25, 15) {real, imag} */,
  {32'h452ebecc, 32'h00000000} /* (1, 25, 14) {real, imag} */,
  {32'h4503cd6f, 32'h00000000} /* (1, 25, 13) {real, imag} */,
  {32'h45073348, 32'h00000000} /* (1, 25, 12) {real, imag} */,
  {32'h44d68fbe, 32'h00000000} /* (1, 25, 11) {real, imag} */,
  {32'h4392e010, 32'h00000000} /* (1, 25, 10) {real, imag} */,
  {32'hc533abec, 32'h00000000} /* (1, 25, 9) {real, imag} */,
  {32'hc5260c14, 32'h00000000} /* (1, 25, 8) {real, imag} */,
  {32'hc517fd82, 32'h00000000} /* (1, 25, 7) {real, imag} */,
  {32'hc5109969, 32'h00000000} /* (1, 25, 6) {real, imag} */,
  {32'hc4e6202c, 32'h00000000} /* (1, 25, 5) {real, imag} */,
  {32'hc5490f8b, 32'h00000000} /* (1, 25, 4) {real, imag} */,
  {32'hc53795b4, 32'h00000000} /* (1, 25, 3) {real, imag} */,
  {32'hc50989ea, 32'h00000000} /* (1, 25, 2) {real, imag} */,
  {32'hc57b5fff, 32'h00000000} /* (1, 25, 1) {real, imag} */,
  {32'hc53df45c, 32'h00000000} /* (1, 25, 0) {real, imag} */,
  {32'hc528975a, 32'h00000000} /* (1, 24, 31) {real, imag} */,
  {32'hc52dc10d, 32'h00000000} /* (1, 24, 30) {real, imag} */,
  {32'hc5155a2e, 32'h00000000} /* (1, 24, 29) {real, imag} */,
  {32'hc50ff145, 32'h00000000} /* (1, 24, 28) {real, imag} */,
  {32'hc51d00be, 32'h00000000} /* (1, 24, 27) {real, imag} */,
  {32'hc54282b6, 32'h00000000} /* (1, 24, 26) {real, imag} */,
  {32'hc512e4ce, 32'h00000000} /* (1, 24, 25) {real, imag} */,
  {32'hc522044c, 32'h00000000} /* (1, 24, 24) {real, imag} */,
  {32'hc4cbe75f, 32'h00000000} /* (1, 24, 23) {real, imag} */,
  {32'hc43bc2f7, 32'h00000000} /* (1, 24, 22) {real, imag} */,
  {32'h445ea5b2, 32'h00000000} /* (1, 24, 21) {real, imag} */,
  {32'h4585c773, 32'h00000000} /* (1, 24, 20) {real, imag} */,
  {32'h45665c06, 32'h00000000} /* (1, 24, 19) {real, imag} */,
  {32'h4573326e, 32'h00000000} /* (1, 24, 18) {real, imag} */,
  {32'h45633824, 32'h00000000} /* (1, 24, 17) {real, imag} */,
  {32'h452776b4, 32'h00000000} /* (1, 24, 16) {real, imag} */,
  {32'h454824a6, 32'h00000000} /* (1, 24, 15) {real, imag} */,
  {32'h456880ff, 32'h00000000} /* (1, 24, 14) {real, imag} */,
  {32'h4521ef6a, 32'h00000000} /* (1, 24, 13) {real, imag} */,
  {32'h44ecdab2, 32'h00000000} /* (1, 24, 12) {real, imag} */,
  {32'h44b393a2, 32'h00000000} /* (1, 24, 11) {real, imag} */,
  {32'hc4b6497b, 32'h00000000} /* (1, 24, 10) {real, imag} */,
  {32'hc517c418, 32'h00000000} /* (1, 24, 9) {real, imag} */,
  {32'hc523a0c0, 32'h00000000} /* (1, 24, 8) {real, imag} */,
  {32'hc509a5ad, 32'h00000000} /* (1, 24, 7) {real, imag} */,
  {32'hc4f33724, 32'h00000000} /* (1, 24, 6) {real, imag} */,
  {32'hc5205ae2, 32'h00000000} /* (1, 24, 5) {real, imag} */,
  {32'hc50bee67, 32'h00000000} /* (1, 24, 4) {real, imag} */,
  {32'hc5191f40, 32'h00000000} /* (1, 24, 3) {real, imag} */,
  {32'hc52ae28c, 32'h00000000} /* (1, 24, 2) {real, imag} */,
  {32'hc50fd938, 32'h00000000} /* (1, 24, 1) {real, imag} */,
  {32'hc523b6fc, 32'h00000000} /* (1, 24, 0) {real, imag} */,
  {32'hc5128138, 32'h00000000} /* (1, 23, 31) {real, imag} */,
  {32'hc51aab54, 32'h00000000} /* (1, 23, 30) {real, imag} */,
  {32'hc5183605, 32'h00000000} /* (1, 23, 29) {real, imag} */,
  {32'hc5004e51, 32'h00000000} /* (1, 23, 28) {real, imag} */,
  {32'hc51c9cb8, 32'h00000000} /* (1, 23, 27) {real, imag} */,
  {32'hc525d278, 32'h00000000} /* (1, 23, 26) {real, imag} */,
  {32'hc506c1dc, 32'h00000000} /* (1, 23, 25) {real, imag} */,
  {32'hc4b62862, 32'h00000000} /* (1, 23, 24) {real, imag} */,
  {32'hc459611d, 32'h00000000} /* (1, 23, 23) {real, imag} */,
  {32'h43afa1a8, 32'h00000000} /* (1, 23, 22) {real, imag} */,
  {32'h443a4861, 32'h00000000} /* (1, 23, 21) {real, imag} */,
  {32'h45288a47, 32'h00000000} /* (1, 23, 20) {real, imag} */,
  {32'h4532aa4d, 32'h00000000} /* (1, 23, 19) {real, imag} */,
  {32'h4541b742, 32'h00000000} /* (1, 23, 18) {real, imag} */,
  {32'h453389be, 32'h00000000} /* (1, 23, 17) {real, imag} */,
  {32'h452a94ab, 32'h00000000} /* (1, 23, 16) {real, imag} */,
  {32'h45244c10, 32'h00000000} /* (1, 23, 15) {real, imag} */,
  {32'h45175f3e, 32'h00000000} /* (1, 23, 14) {real, imag} */,
  {32'h452dab05, 32'h00000000} /* (1, 23, 13) {real, imag} */,
  {32'h44fa7be1, 32'h00000000} /* (1, 23, 12) {real, imag} */,
  {32'h451f1b14, 32'h00000000} /* (1, 23, 11) {real, imag} */,
  {32'hc398838c, 32'h00000000} /* (1, 23, 10) {real, imag} */,
  {32'hc48476a1, 32'h00000000} /* (1, 23, 9) {real, imag} */,
  {32'hc510759d, 32'h00000000} /* (1, 23, 8) {real, imag} */,
  {32'hc500a206, 32'h00000000} /* (1, 23, 7) {real, imag} */,
  {32'hc4979234, 32'h00000000} /* (1, 23, 6) {real, imag} */,
  {32'hc4dfa970, 32'h00000000} /* (1, 23, 5) {real, imag} */,
  {32'hc4fe9fbe, 32'h00000000} /* (1, 23, 4) {real, imag} */,
  {32'hc4d301b6, 32'h00000000} /* (1, 23, 3) {real, imag} */,
  {32'hc4ef5233, 32'h00000000} /* (1, 23, 2) {real, imag} */,
  {32'hc52bb37a, 32'h00000000} /* (1, 23, 1) {real, imag} */,
  {32'hc4e9c8a6, 32'h00000000} /* (1, 23, 0) {real, imag} */,
  {32'hc4e41c28, 32'h00000000} /* (1, 22, 31) {real, imag} */,
  {32'hc486e158, 32'h00000000} /* (1, 22, 30) {real, imag} */,
  {32'hc4a773d4, 32'h00000000} /* (1, 22, 29) {real, imag} */,
  {32'hc5337d12, 32'h00000000} /* (1, 22, 28) {real, imag} */,
  {32'hc53416da, 32'h00000000} /* (1, 22, 27) {real, imag} */,
  {32'hc4f76a1e, 32'h00000000} /* (1, 22, 26) {real, imag} */,
  {32'hc4db878a, 32'h00000000} /* (1, 22, 25) {real, imag} */,
  {32'hc45b373d, 32'h00000000} /* (1, 22, 24) {real, imag} */,
  {32'hc37606b0, 32'h00000000} /* (1, 22, 23) {real, imag} */,
  {32'hc2ebcdd4, 32'h00000000} /* (1, 22, 22) {real, imag} */,
  {32'h4252cb70, 32'h00000000} /* (1, 22, 21) {real, imag} */,
  {32'h451e98fd, 32'h00000000} /* (1, 22, 20) {real, imag} */,
  {32'h450ecb97, 32'h00000000} /* (1, 22, 19) {real, imag} */,
  {32'h44ccc1b8, 32'h00000000} /* (1, 22, 18) {real, imag} */,
  {32'h45119ff6, 32'h00000000} /* (1, 22, 17) {real, imag} */,
  {32'h453c9b77, 32'h00000000} /* (1, 22, 16) {real, imag} */,
  {32'h44e8a2dc, 32'h00000000} /* (1, 22, 15) {real, imag} */,
  {32'h4511a02a, 32'h00000000} /* (1, 22, 14) {real, imag} */,
  {32'h4515ed77, 32'h00000000} /* (1, 22, 13) {real, imag} */,
  {32'h450f6430, 32'h00000000} /* (1, 22, 12) {real, imag} */,
  {32'h44c70efb, 32'h00000000} /* (1, 22, 11) {real, imag} */,
  {32'hc2912788, 32'h00000000} /* (1, 22, 10) {real, imag} */,
  {32'hc4c68808, 32'h00000000} /* (1, 22, 9) {real, imag} */,
  {32'hc4c9b8f4, 32'h00000000} /* (1, 22, 8) {real, imag} */,
  {32'hc496f45a, 32'h00000000} /* (1, 22, 7) {real, imag} */,
  {32'hc48be82f, 32'h00000000} /* (1, 22, 6) {real, imag} */,
  {32'hc4aff420, 32'h00000000} /* (1, 22, 5) {real, imag} */,
  {32'hc49dc344, 32'h00000000} /* (1, 22, 4) {real, imag} */,
  {32'hc4ae7e7a, 32'h00000000} /* (1, 22, 3) {real, imag} */,
  {32'hc4d095d6, 32'h00000000} /* (1, 22, 2) {real, imag} */,
  {32'hc4d9dca3, 32'h00000000} /* (1, 22, 1) {real, imag} */,
  {32'hc4b5e0ea, 32'h00000000} /* (1, 22, 0) {real, imag} */,
  {32'hc4bbd3d7, 32'h00000000} /* (1, 21, 31) {real, imag} */,
  {32'hc44d969b, 32'h00000000} /* (1, 21, 30) {real, imag} */,
  {32'h4172acc0, 32'h00000000} /* (1, 21, 29) {real, imag} */,
  {32'hc4ccd4c8, 32'h00000000} /* (1, 21, 28) {real, imag} */,
  {32'hc4184858, 32'h00000000} /* (1, 21, 27) {real, imag} */,
  {32'hc313c7de, 32'h00000000} /* (1, 21, 26) {real, imag} */,
  {32'hc3482d96, 32'h00000000} /* (1, 21, 25) {real, imag} */,
  {32'hc39164ac, 32'h00000000} /* (1, 21, 24) {real, imag} */,
  {32'h3e603800, 32'h00000000} /* (1, 21, 23) {real, imag} */,
  {32'hc262e2dc, 32'h00000000} /* (1, 21, 22) {real, imag} */,
  {32'h43440398, 32'h00000000} /* (1, 21, 21) {real, imag} */,
  {32'h43e38859, 32'h00000000} /* (1, 21, 20) {real, imag} */,
  {32'h44714d84, 32'h00000000} /* (1, 21, 19) {real, imag} */,
  {32'h44c3a7bb, 32'h00000000} /* (1, 21, 18) {real, imag} */,
  {32'h43ae4b5e, 32'h00000000} /* (1, 21, 17) {real, imag} */,
  {32'h44135814, 32'h00000000} /* (1, 21, 16) {real, imag} */,
  {32'h44c6cee5, 32'h00000000} /* (1, 21, 15) {real, imag} */,
  {32'h4476f705, 32'h00000000} /* (1, 21, 14) {real, imag} */,
  {32'h44962a34, 32'h00000000} /* (1, 21, 13) {real, imag} */,
  {32'h448602ec, 32'h00000000} /* (1, 21, 12) {real, imag} */,
  {32'h4443253c, 32'h00000000} /* (1, 21, 11) {real, imag} */,
  {32'h4332c31e, 32'h00000000} /* (1, 21, 10) {real, imag} */,
  {32'hc4427b2a, 32'h00000000} /* (1, 21, 9) {real, imag} */,
  {32'hc46d98e6, 32'h00000000} /* (1, 21, 8) {real, imag} */,
  {32'hc3c38bfd, 32'h00000000} /* (1, 21, 7) {real, imag} */,
  {32'hc3d38d58, 32'h00000000} /* (1, 21, 6) {real, imag} */,
  {32'hc3df9a9a, 32'h00000000} /* (1, 21, 5) {real, imag} */,
  {32'hc3ea91a5, 32'h00000000} /* (1, 21, 4) {real, imag} */,
  {32'hc1d21ea0, 32'h00000000} /* (1, 21, 3) {real, imag} */,
  {32'hc426016e, 32'h00000000} /* (1, 21, 2) {real, imag} */,
  {32'hc4287f4c, 32'h00000000} /* (1, 21, 1) {real, imag} */,
  {32'hc429b634, 32'h00000000} /* (1, 21, 0) {real, imag} */,
  {32'h44457de4, 32'h00000000} /* (1, 20, 31) {real, imag} */,
  {32'h448ce8dd, 32'h00000000} /* (1, 20, 30) {real, imag} */,
  {32'h44f0a9aa, 32'h00000000} /* (1, 20, 29) {real, imag} */,
  {32'h44d6843a, 32'h00000000} /* (1, 20, 28) {real, imag} */,
  {32'h44a8be24, 32'h00000000} /* (1, 20, 27) {real, imag} */,
  {32'h44831464, 32'h00000000} /* (1, 20, 26) {real, imag} */,
  {32'h4526a292, 32'h00000000} /* (1, 20, 25) {real, imag} */,
  {32'h451396ce, 32'h00000000} /* (1, 20, 24) {real, imag} */,
  {32'h44c77cbe, 32'h00000000} /* (1, 20, 23) {real, imag} */,
  {32'h45075418, 32'h00000000} /* (1, 20, 22) {real, imag} */,
  {32'h446f17a7, 32'h00000000} /* (1, 20, 21) {real, imag} */,
  {32'hc02ac700, 32'h00000000} /* (1, 20, 20) {real, imag} */,
  {32'hc485b11b, 32'h00000000} /* (1, 20, 19) {real, imag} */,
  {32'hc4abafd3, 32'h00000000} /* (1, 20, 18) {real, imag} */,
  {32'hc4670380, 32'h00000000} /* (1, 20, 17) {real, imag} */,
  {32'hc4a245b8, 32'h00000000} /* (1, 20, 16) {real, imag} */,
  {32'hc4eb12e2, 32'h00000000} /* (1, 20, 15) {real, imag} */,
  {32'hc4167dce, 32'h00000000} /* (1, 20, 14) {real, imag} */,
  {32'hc4267fcc, 32'h00000000} /* (1, 20, 13) {real, imag} */,
  {32'hc40c2508, 32'h00000000} /* (1, 20, 12) {real, imag} */,
  {32'hc3e3aa0c, 32'h00000000} /* (1, 20, 11) {real, imag} */,
  {32'h41e1bde0, 32'h00000000} /* (1, 20, 10) {real, imag} */,
  {32'h442a5cad, 32'h00000000} /* (1, 20, 9) {real, imag} */,
  {32'h442a61d8, 32'h00000000} /* (1, 20, 8) {real, imag} */,
  {32'h445fe2d9, 32'h00000000} /* (1, 20, 7) {real, imag} */,
  {32'h448ed306, 32'h00000000} /* (1, 20, 6) {real, imag} */,
  {32'h447087a5, 32'h00000000} /* (1, 20, 5) {real, imag} */,
  {32'h44851e8c, 32'h00000000} /* (1, 20, 4) {real, imag} */,
  {32'h44a5ecf1, 32'h00000000} /* (1, 20, 3) {real, imag} */,
  {32'h4506bb00, 32'h00000000} /* (1, 20, 2) {real, imag} */,
  {32'h44378bd8, 32'h00000000} /* (1, 20, 1) {real, imag} */,
  {32'h41c38f20, 32'h00000000} /* (1, 20, 0) {real, imag} */,
  {32'h44f9c0f4, 32'h00000000} /* (1, 19, 31) {real, imag} */,
  {32'h4505be4c, 32'h00000000} /* (1, 19, 30) {real, imag} */,
  {32'h4510c4a2, 32'h00000000} /* (1, 19, 29) {real, imag} */,
  {32'h44ecc32f, 32'h00000000} /* (1, 19, 28) {real, imag} */,
  {32'h451714c6, 32'h00000000} /* (1, 19, 27) {real, imag} */,
  {32'h450a1082, 32'h00000000} /* (1, 19, 26) {real, imag} */,
  {32'h4541c212, 32'h00000000} /* (1, 19, 25) {real, imag} */,
  {32'h45281a92, 32'h00000000} /* (1, 19, 24) {real, imag} */,
  {32'h454f2fde, 32'h00000000} /* (1, 19, 23) {real, imag} */,
  {32'h452973fe, 32'h00000000} /* (1, 19, 22) {real, imag} */,
  {32'h44b62cb0, 32'h00000000} /* (1, 19, 21) {real, imag} */,
  {32'hc41734b6, 32'h00000000} /* (1, 19, 20) {real, imag} */,
  {32'hc47f9022, 32'h00000000} /* (1, 19, 19) {real, imag} */,
  {32'hc4ebfe03, 32'h00000000} /* (1, 19, 18) {real, imag} */,
  {32'hc4f3c562, 32'h00000000} /* (1, 19, 17) {real, imag} */,
  {32'hc4f8266c, 32'h00000000} /* (1, 19, 16) {real, imag} */,
  {32'hc4e0d348, 32'h00000000} /* (1, 19, 15) {real, imag} */,
  {32'hc4d2f036, 32'h00000000} /* (1, 19, 14) {real, imag} */,
  {32'hc4d65381, 32'h00000000} /* (1, 19, 13) {real, imag} */,
  {32'hc4fe34fb, 32'h00000000} /* (1, 19, 12) {real, imag} */,
  {32'hc49ee524, 32'h00000000} /* (1, 19, 11) {real, imag} */,
  {32'hc34fdde8, 32'h00000000} /* (1, 19, 10) {real, imag} */,
  {32'h4462b998, 32'h00000000} /* (1, 19, 9) {real, imag} */,
  {32'h44d673fc, 32'h00000000} /* (1, 19, 8) {real, imag} */,
  {32'h45060244, 32'h00000000} /* (1, 19, 7) {real, imag} */,
  {32'h45015fd2, 32'h00000000} /* (1, 19, 6) {real, imag} */,
  {32'h4509c038, 32'h00000000} /* (1, 19, 5) {real, imag} */,
  {32'h45248f0c, 32'h00000000} /* (1, 19, 4) {real, imag} */,
  {32'h4550bd42, 32'h00000000} /* (1, 19, 3) {real, imag} */,
  {32'h44cef083, 32'h00000000} /* (1, 19, 2) {real, imag} */,
  {32'h4510ce93, 32'h00000000} /* (1, 19, 1) {real, imag} */,
  {32'h44c1f866, 32'h00000000} /* (1, 19, 0) {real, imag} */,
  {32'h44d49553, 32'h00000000} /* (1, 18, 31) {real, imag} */,
  {32'h451addca, 32'h00000000} /* (1, 18, 30) {real, imag} */,
  {32'h44efafb2, 32'h00000000} /* (1, 18, 29) {real, imag} */,
  {32'h44ffdae3, 32'h00000000} /* (1, 18, 28) {real, imag} */,
  {32'h45554013, 32'h00000000} /* (1, 18, 27) {real, imag} */,
  {32'h455ffc6f, 32'h00000000} /* (1, 18, 26) {real, imag} */,
  {32'h45348bc3, 32'h00000000} /* (1, 18, 25) {real, imag} */,
  {32'h4542a3ca, 32'h00000000} /* (1, 18, 24) {real, imag} */,
  {32'h45264d18, 32'h00000000} /* (1, 18, 23) {real, imag} */,
  {32'h4515472c, 32'h00000000} /* (1, 18, 22) {real, imag} */,
  {32'h43a31b40, 32'h00000000} /* (1, 18, 21) {real, imag} */,
  {32'hc42a4980, 32'h00000000} /* (1, 18, 20) {real, imag} */,
  {32'hc4abcd86, 32'h00000000} /* (1, 18, 19) {real, imag} */,
  {32'hc4df2728, 32'h00000000} /* (1, 18, 18) {real, imag} */,
  {32'hc5064b4a, 32'h00000000} /* (1, 18, 17) {real, imag} */,
  {32'hc4f8dcfa, 32'h00000000} /* (1, 18, 16) {real, imag} */,
  {32'hc4e88559, 32'h00000000} /* (1, 18, 15) {real, imag} */,
  {32'hc51e7d1e, 32'h00000000} /* (1, 18, 14) {real, imag} */,
  {32'hc52d772f, 32'h00000000} /* (1, 18, 13) {real, imag} */,
  {32'hc4b09fc7, 32'h00000000} /* (1, 18, 12) {real, imag} */,
  {32'hc43732b4, 32'h00000000} /* (1, 18, 11) {real, imag} */,
  {32'h44726abc, 32'h00000000} /* (1, 18, 10) {real, imag} */,
  {32'h44cd273e, 32'h00000000} /* (1, 18, 9) {real, imag} */,
  {32'h44e78409, 32'h00000000} /* (1, 18, 8) {real, imag} */,
  {32'h45666c00, 32'h00000000} /* (1, 18, 7) {real, imag} */,
  {32'h45047f70, 32'h00000000} /* (1, 18, 6) {real, imag} */,
  {32'h451a0914, 32'h00000000} /* (1, 18, 5) {real, imag} */,
  {32'h450c54a8, 32'h00000000} /* (1, 18, 4) {real, imag} */,
  {32'h4521fe67, 32'h00000000} /* (1, 18, 3) {real, imag} */,
  {32'h452956c6, 32'h00000000} /* (1, 18, 2) {real, imag} */,
  {32'h44b6f5ee, 32'h00000000} /* (1, 18, 1) {real, imag} */,
  {32'h451ad1a1, 32'h00000000} /* (1, 18, 0) {real, imag} */,
  {32'h452e9926, 32'h00000000} /* (1, 17, 31) {real, imag} */,
  {32'h45413776, 32'h00000000} /* (1, 17, 30) {real, imag} */,
  {32'h451d5862, 32'h00000000} /* (1, 17, 29) {real, imag} */,
  {32'h4555ee2c, 32'h00000000} /* (1, 17, 28) {real, imag} */,
  {32'h4558f71e, 32'h00000000} /* (1, 17, 27) {real, imag} */,
  {32'h4558eb1b, 32'h00000000} /* (1, 17, 26) {real, imag} */,
  {32'h456fea82, 32'h00000000} /* (1, 17, 25) {real, imag} */,
  {32'h4525442d, 32'h00000000} /* (1, 17, 24) {real, imag} */,
  {32'h455c581f, 32'h00000000} /* (1, 17, 23) {real, imag} */,
  {32'h453b55cb, 32'h00000000} /* (1, 17, 22) {real, imag} */,
  {32'h430ed150, 32'h00000000} /* (1, 17, 21) {real, imag} */,
  {32'hc406ca98, 32'h00000000} /* (1, 17, 20) {real, imag} */,
  {32'hc4d66bbc, 32'h00000000} /* (1, 17, 19) {real, imag} */,
  {32'hc511504a, 32'h00000000} /* (1, 17, 18) {real, imag} */,
  {32'hc51ea37c, 32'h00000000} /* (1, 17, 17) {real, imag} */,
  {32'hc534f20f, 32'h00000000} /* (1, 17, 16) {real, imag} */,
  {32'hc5196d6e, 32'h00000000} /* (1, 17, 15) {real, imag} */,
  {32'hc4f5b6a7, 32'h00000000} /* (1, 17, 14) {real, imag} */,
  {32'hc52180aa, 32'h00000000} /* (1, 17, 13) {real, imag} */,
  {32'hc5096c10, 32'h00000000} /* (1, 17, 12) {real, imag} */,
  {32'hc48e876d, 32'h00000000} /* (1, 17, 11) {real, imag} */,
  {32'h449e166a, 32'h00000000} /* (1, 17, 10) {real, imag} */,
  {32'h450ef5e6, 32'h00000000} /* (1, 17, 9) {real, imag} */,
  {32'h45362a95, 32'h00000000} /* (1, 17, 8) {real, imag} */,
  {32'h450c117d, 32'h00000000} /* (1, 17, 7) {real, imag} */,
  {32'h4581b04c, 32'h00000000} /* (1, 17, 6) {real, imag} */,
  {32'h4533b7f5, 32'h00000000} /* (1, 17, 5) {real, imag} */,
  {32'h450510bf, 32'h00000000} /* (1, 17, 4) {real, imag} */,
  {32'h45015014, 32'h00000000} /* (1, 17, 3) {real, imag} */,
  {32'h4502e608, 32'h00000000} /* (1, 17, 2) {real, imag} */,
  {32'h450bbda0, 32'h00000000} /* (1, 17, 1) {real, imag} */,
  {32'h44ec18a2, 32'h00000000} /* (1, 17, 0) {real, imag} */,
  {32'h44f2f5ca, 32'h00000000} /* (1, 16, 31) {real, imag} */,
  {32'h4522afce, 32'h00000000} /* (1, 16, 30) {real, imag} */,
  {32'h454cc5c3, 32'h00000000} /* (1, 16, 29) {real, imag} */,
  {32'h454d5d7f, 32'h00000000} /* (1, 16, 28) {real, imag} */,
  {32'h4554559f, 32'h00000000} /* (1, 16, 27) {real, imag} */,
  {32'h45403460, 32'h00000000} /* (1, 16, 26) {real, imag} */,
  {32'h454acf64, 32'h00000000} /* (1, 16, 25) {real, imag} */,
  {32'h45071c20, 32'h00000000} /* (1, 16, 24) {real, imag} */,
  {32'h453477e3, 32'h00000000} /* (1, 16, 23) {real, imag} */,
  {32'h454a3952, 32'h00000000} /* (1, 16, 22) {real, imag} */,
  {32'h44c7b88e, 32'h00000000} /* (1, 16, 21) {real, imag} */,
  {32'hc43a9f46, 32'h00000000} /* (1, 16, 20) {real, imag} */,
  {32'hc4e94b02, 32'h00000000} /* (1, 16, 19) {real, imag} */,
  {32'hc51445d6, 32'h00000000} /* (1, 16, 18) {real, imag} */,
  {32'hc5402bce, 32'h00000000} /* (1, 16, 17) {real, imag} */,
  {32'hc533be96, 32'h00000000} /* (1, 16, 16) {real, imag} */,
  {32'hc5360871, 32'h00000000} /* (1, 16, 15) {real, imag} */,
  {32'hc53506e4, 32'h00000000} /* (1, 16, 14) {real, imag} */,
  {32'hc50d11dd, 32'h00000000} /* (1, 16, 13) {real, imag} */,
  {32'hc501eca9, 32'h00000000} /* (1, 16, 12) {real, imag} */,
  {32'hc4ac99b2, 32'h00000000} /* (1, 16, 11) {real, imag} */,
  {32'h4411c00e, 32'h00000000} /* (1, 16, 10) {real, imag} */,
  {32'h453c2d1c, 32'h00000000} /* (1, 16, 9) {real, imag} */,
  {32'h452eed2c, 32'h00000000} /* (1, 16, 8) {real, imag} */,
  {32'h45412079, 32'h00000000} /* (1, 16, 7) {real, imag} */,
  {32'h45648068, 32'h00000000} /* (1, 16, 6) {real, imag} */,
  {32'h451bf1e1, 32'h00000000} /* (1, 16, 5) {real, imag} */,
  {32'h45094dae, 32'h00000000} /* (1, 16, 4) {real, imag} */,
  {32'h4500aa69, 32'h00000000} /* (1, 16, 3) {real, imag} */,
  {32'h44fb04b9, 32'h00000000} /* (1, 16, 2) {real, imag} */,
  {32'h453fcbf6, 32'h00000000} /* (1, 16, 1) {real, imag} */,
  {32'h4525c63e, 32'h00000000} /* (1, 16, 0) {real, imag} */,
  {32'h4511979d, 32'h00000000} /* (1, 15, 31) {real, imag} */,
  {32'h453bcf0e, 32'h00000000} /* (1, 15, 30) {real, imag} */,
  {32'h45806980, 32'h00000000} /* (1, 15, 29) {real, imag} */,
  {32'h4558917a, 32'h00000000} /* (1, 15, 28) {real, imag} */,
  {32'h4552e967, 32'h00000000} /* (1, 15, 27) {real, imag} */,
  {32'h4550a94e, 32'h00000000} /* (1, 15, 26) {real, imag} */,
  {32'h452e2ada, 32'h00000000} /* (1, 15, 25) {real, imag} */,
  {32'h452ca672, 32'h00000000} /* (1, 15, 24) {real, imag} */,
  {32'h44fee8b7, 32'h00000000} /* (1, 15, 23) {real, imag} */,
  {32'h450b3231, 32'h00000000} /* (1, 15, 22) {real, imag} */,
  {32'h44bd0f02, 32'h00000000} /* (1, 15, 21) {real, imag} */,
  {32'hc4b5d4ab, 32'h00000000} /* (1, 15, 20) {real, imag} */,
  {32'hc50fccb5, 32'h00000000} /* (1, 15, 19) {real, imag} */,
  {32'hc504fe5a, 32'h00000000} /* (1, 15, 18) {real, imag} */,
  {32'hc50e6acf, 32'h00000000} /* (1, 15, 17) {real, imag} */,
  {32'hc546962c, 32'h00000000} /* (1, 15, 16) {real, imag} */,
  {32'hc522ad0f, 32'h00000000} /* (1, 15, 15) {real, imag} */,
  {32'hc522e3fc, 32'h00000000} /* (1, 15, 14) {real, imag} */,
  {32'hc54365fa, 32'h00000000} /* (1, 15, 13) {real, imag} */,
  {32'hc52e2d26, 32'h00000000} /* (1, 15, 12) {real, imag} */,
  {32'hc4ba00e6, 32'h00000000} /* (1, 15, 11) {real, imag} */,
  {32'h4335e088, 32'h00000000} /* (1, 15, 10) {real, imag} */,
  {32'h4502f1a4, 32'h00000000} /* (1, 15, 9) {real, imag} */,
  {32'h45157476, 32'h00000000} /* (1, 15, 8) {real, imag} */,
  {32'h454062cc, 32'h00000000} /* (1, 15, 7) {real, imag} */,
  {32'h4550e9f7, 32'h00000000} /* (1, 15, 6) {real, imag} */,
  {32'h453456d7, 32'h00000000} /* (1, 15, 5) {real, imag} */,
  {32'h4554e734, 32'h00000000} /* (1, 15, 4) {real, imag} */,
  {32'h4523d7cb, 32'h00000000} /* (1, 15, 3) {real, imag} */,
  {32'h4542b8c4, 32'h00000000} /* (1, 15, 2) {real, imag} */,
  {32'h456da98b, 32'h00000000} /* (1, 15, 1) {real, imag} */,
  {32'h451bd0c8, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'h452f84a3, 32'h00000000} /* (1, 14, 31) {real, imag} */,
  {32'h457fb6f5, 32'h00000000} /* (1, 14, 30) {real, imag} */,
  {32'h45672af4, 32'h00000000} /* (1, 14, 29) {real, imag} */,
  {32'h45516986, 32'h00000000} /* (1, 14, 28) {real, imag} */,
  {32'h456fbc28, 32'h00000000} /* (1, 14, 27) {real, imag} */,
  {32'h456190fe, 32'h00000000} /* (1, 14, 26) {real, imag} */,
  {32'h453f04bd, 32'h00000000} /* (1, 14, 25) {real, imag} */,
  {32'h452607dd, 32'h00000000} /* (1, 14, 24) {real, imag} */,
  {32'h450aa5d1, 32'h00000000} /* (1, 14, 23) {real, imag} */,
  {32'h450ac7cc, 32'h00000000} /* (1, 14, 22) {real, imag} */,
  {32'h43e724d4, 32'h00000000} /* (1, 14, 21) {real, imag} */,
  {32'hc48b611e, 32'h00000000} /* (1, 14, 20) {real, imag} */,
  {32'hc518f307, 32'h00000000} /* (1, 14, 19) {real, imag} */,
  {32'hc54efafd, 32'h00000000} /* (1, 14, 18) {real, imag} */,
  {32'hc571d8dd, 32'h00000000} /* (1, 14, 17) {real, imag} */,
  {32'hc505b2fa, 32'h00000000} /* (1, 14, 16) {real, imag} */,
  {32'hc547d1f5, 32'h00000000} /* (1, 14, 15) {real, imag} */,
  {32'hc54e62b5, 32'h00000000} /* (1, 14, 14) {real, imag} */,
  {32'hc56e1c1a, 32'h00000000} /* (1, 14, 13) {real, imag} */,
  {32'hc52a2038, 32'h00000000} /* (1, 14, 12) {real, imag} */,
  {32'hc4af8d40, 32'h00000000} /* (1, 14, 11) {real, imag} */,
  {32'h440ed7c6, 32'h00000000} /* (1, 14, 10) {real, imag} */,
  {32'h44ca4462, 32'h00000000} /* (1, 14, 9) {real, imag} */,
  {32'h451826f3, 32'h00000000} /* (1, 14, 8) {real, imag} */,
  {32'h451367bd, 32'h00000000} /* (1, 14, 7) {real, imag} */,
  {32'h452df120, 32'h00000000} /* (1, 14, 6) {real, imag} */,
  {32'h45351324, 32'h00000000} /* (1, 14, 5) {real, imag} */,
  {32'h453349d3, 32'h00000000} /* (1, 14, 4) {real, imag} */,
  {32'h45474561, 32'h00000000} /* (1, 14, 3) {real, imag} */,
  {32'h4547fc17, 32'h00000000} /* (1, 14, 2) {real, imag} */,
  {32'h4530e4df, 32'h00000000} /* (1, 14, 1) {real, imag} */,
  {32'h45021e8c, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'h4508e36e, 32'h00000000} /* (1, 13, 31) {real, imag} */,
  {32'h452f3849, 32'h00000000} /* (1, 13, 30) {real, imag} */,
  {32'h45878032, 32'h00000000} /* (1, 13, 29) {real, imag} */,
  {32'h45573d90, 32'h00000000} /* (1, 13, 28) {real, imag} */,
  {32'h457551df, 32'h00000000} /* (1, 13, 27) {real, imag} */,
  {32'h45787d88, 32'h00000000} /* (1, 13, 26) {real, imag} */,
  {32'h45565da5, 32'h00000000} /* (1, 13, 25) {real, imag} */,
  {32'h451404e4, 32'h00000000} /* (1, 13, 24) {real, imag} */,
  {32'h44f400b2, 32'h00000000} /* (1, 13, 23) {real, imag} */,
  {32'h45003503, 32'h00000000} /* (1, 13, 22) {real, imag} */,
  {32'h43e9d518, 32'h00000000} /* (1, 13, 21) {real, imag} */,
  {32'hc4a9ea72, 32'h00000000} /* (1, 13, 20) {real, imag} */,
  {32'hc549ece3, 32'h00000000} /* (1, 13, 19) {real, imag} */,
  {32'hc5460487, 32'h00000000} /* (1, 13, 18) {real, imag} */,
  {32'hc56a1033, 32'h00000000} /* (1, 13, 17) {real, imag} */,
  {32'hc58b1ead, 32'h00000000} /* (1, 13, 16) {real, imag} */,
  {32'hc51ca294, 32'h00000000} /* (1, 13, 15) {real, imag} */,
  {32'hc5234ae5, 32'h00000000} /* (1, 13, 14) {real, imag} */,
  {32'hc515ca4f, 32'h00000000} /* (1, 13, 13) {real, imag} */,
  {32'hc522e9ce, 32'h00000000} /* (1, 13, 12) {real, imag} */,
  {32'hc50bc14d, 32'h00000000} /* (1, 13, 11) {real, imag} */,
  {32'h41d4b3c0, 32'h00000000} /* (1, 13, 10) {real, imag} */,
  {32'h44bf3216, 32'h00000000} /* (1, 13, 9) {real, imag} */,
  {32'h45375e5c, 32'h00000000} /* (1, 13, 8) {real, imag} */,
  {32'h4529c097, 32'h00000000} /* (1, 13, 7) {real, imag} */,
  {32'h44c66ac2, 32'h00000000} /* (1, 13, 6) {real, imag} */,
  {32'h452e48a7, 32'h00000000} /* (1, 13, 5) {real, imag} */,
  {32'h450bea7e, 32'h00000000} /* (1, 13, 4) {real, imag} */,
  {32'h452f8ea9, 32'h00000000} /* (1, 13, 3) {real, imag} */,
  {32'h456302bb, 32'h00000000} /* (1, 13, 2) {real, imag} */,
  {32'h45194955, 32'h00000000} /* (1, 13, 1) {real, imag} */,
  {32'h4528d222, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'h44cc5af9, 32'h00000000} /* (1, 12, 31) {real, imag} */,
  {32'h450d36d0, 32'h00000000} /* (1, 12, 30) {real, imag} */,
  {32'h45305ea5, 32'h00000000} /* (1, 12, 29) {real, imag} */,
  {32'h45452dd8, 32'h00000000} /* (1, 12, 28) {real, imag} */,
  {32'h452b2b85, 32'h00000000} /* (1, 12, 27) {real, imag} */,
  {32'h452933c5, 32'h00000000} /* (1, 12, 26) {real, imag} */,
  {32'h450991cc, 32'h00000000} /* (1, 12, 25) {real, imag} */,
  {32'h454218f7, 32'h00000000} /* (1, 12, 24) {real, imag} */,
  {32'h4564511a, 32'h00000000} /* (1, 12, 23) {real, imag} */,
  {32'h451897f8, 32'h00000000} /* (1, 12, 22) {real, imag} */,
  {32'h4481ec36, 32'h00000000} /* (1, 12, 21) {real, imag} */,
  {32'hc4b318cc, 32'h00000000} /* (1, 12, 20) {real, imag} */,
  {32'hc536e66c, 32'h00000000} /* (1, 12, 19) {real, imag} */,
  {32'hc5085457, 32'h00000000} /* (1, 12, 18) {real, imag} */,
  {32'hc55dfad6, 32'h00000000} /* (1, 12, 17) {real, imag} */,
  {32'hc5563243, 32'h00000000} /* (1, 12, 16) {real, imag} */,
  {32'hc4ec9ea3, 32'h00000000} /* (1, 12, 15) {real, imag} */,
  {32'hc4ffa63d, 32'h00000000} /* (1, 12, 14) {real, imag} */,
  {32'hc4e84ede, 32'h00000000} /* (1, 12, 13) {real, imag} */,
  {32'hc4e36a18, 32'h00000000} /* (1, 12, 12) {real, imag} */,
  {32'hc504cd6f, 32'h00000000} /* (1, 12, 11) {real, imag} */,
  {32'h43a9f1f8, 32'h00000000} /* (1, 12, 10) {real, imag} */,
  {32'h44b53ed0, 32'h00000000} /* (1, 12, 9) {real, imag} */,
  {32'h44c27b2e, 32'h00000000} /* (1, 12, 8) {real, imag} */,
  {32'h45101eae, 32'h00000000} /* (1, 12, 7) {real, imag} */,
  {32'h4518f7ac, 32'h00000000} /* (1, 12, 6) {real, imag} */,
  {32'h4522c22f, 32'h00000000} /* (1, 12, 5) {real, imag} */,
  {32'h451336fd, 32'h00000000} /* (1, 12, 4) {real, imag} */,
  {32'h45281b26, 32'h00000000} /* (1, 12, 3) {real, imag} */,
  {32'h4509b1e1, 32'h00000000} /* (1, 12, 2) {real, imag} */,
  {32'h45213888, 32'h00000000} /* (1, 12, 1) {real, imag} */,
  {32'h451588d9, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'h44a79c6f, 32'h00000000} /* (1, 11, 31) {real, imag} */,
  {32'h44bf7878, 32'h00000000} /* (1, 11, 30) {real, imag} */,
  {32'h44c20d8a, 32'h00000000} /* (1, 11, 29) {real, imag} */,
  {32'h44c8adac, 32'h00000000} /* (1, 11, 28) {real, imag} */,
  {32'h44f75ddf, 32'h00000000} /* (1, 11, 27) {real, imag} */,
  {32'h44b05708, 32'h00000000} /* (1, 11, 26) {real, imag} */,
  {32'h447a8534, 32'h00000000} /* (1, 11, 25) {real, imag} */,
  {32'h4504ce19, 32'h00000000} /* (1, 11, 24) {real, imag} */,
  {32'h4513c3b7, 32'h00000000} /* (1, 11, 23) {real, imag} */,
  {32'h447e91df, 32'h00000000} /* (1, 11, 22) {real, imag} */,
  {32'h442f01c6, 32'h00000000} /* (1, 11, 21) {real, imag} */,
  {32'hc47f1122, 32'h00000000} /* (1, 11, 20) {real, imag} */,
  {32'hc4687262, 32'h00000000} /* (1, 11, 19) {real, imag} */,
  {32'hc4c735b5, 32'h00000000} /* (1, 11, 18) {real, imag} */,
  {32'hc515d7d8, 32'h00000000} /* (1, 11, 17) {real, imag} */,
  {32'hc4afaea0, 32'h00000000} /* (1, 11, 16) {real, imag} */,
  {32'hc50b0fb4, 32'h00000000} /* (1, 11, 15) {real, imag} */,
  {32'hc4fac9d6, 32'h00000000} /* (1, 11, 14) {real, imag} */,
  {32'hc4a38ee6, 32'h00000000} /* (1, 11, 13) {real, imag} */,
  {32'hc51277bc, 32'h00000000} /* (1, 11, 12) {real, imag} */,
  {32'hc4a79915, 32'h00000000} /* (1, 11, 11) {real, imag} */,
  {32'hc328278c, 32'h00000000} /* (1, 11, 10) {real, imag} */,
  {32'h436e1252, 32'h00000000} /* (1, 11, 9) {real, imag} */,
  {32'h44907d1e, 32'h00000000} /* (1, 11, 8) {real, imag} */,
  {32'h44d291f0, 32'h00000000} /* (1, 11, 7) {real, imag} */,
  {32'h450e627d, 32'h00000000} /* (1, 11, 6) {real, imag} */,
  {32'h44e7f409, 32'h00000000} /* (1, 11, 5) {real, imag} */,
  {32'h44a8fdeb, 32'h00000000} /* (1, 11, 4) {real, imag} */,
  {32'h445af9ca, 32'h00000000} /* (1, 11, 3) {real, imag} */,
  {32'h44815d63, 32'h00000000} /* (1, 11, 2) {real, imag} */,
  {32'h44847ab0, 32'h00000000} /* (1, 11, 1) {real, imag} */,
  {32'h447a9328, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'h427c2ff8, 32'h00000000} /* (1, 10, 31) {real, imag} */,
  {32'h42780c12, 32'h00000000} /* (1, 10, 30) {real, imag} */,
  {32'h43822fba, 32'h00000000} /* (1, 10, 29) {real, imag} */,
  {32'hc274177c, 32'h00000000} /* (1, 10, 28) {real, imag} */,
  {32'hc4993854, 32'h00000000} /* (1, 10, 27) {real, imag} */,
  {32'hc454be95, 32'h00000000} /* (1, 10, 26) {real, imag} */,
  {32'hc3a4aa51, 32'h00000000} /* (1, 10, 25) {real, imag} */,
  {32'hc3351d31, 32'h00000000} /* (1, 10, 24) {real, imag} */,
  {32'h42609884, 32'h00000000} /* (1, 10, 23) {real, imag} */,
  {32'hc3b2779b, 32'h00000000} /* (1, 10, 22) {real, imag} */,
  {32'hc428d970, 32'h00000000} /* (1, 10, 21) {real, imag} */,
  {32'h43bf846f, 32'h00000000} /* (1, 10, 20) {real, imag} */,
  {32'h4411d1de, 32'h00000000} /* (1, 10, 19) {real, imag} */,
  {32'h4395ecd4, 32'h00000000} /* (1, 10, 18) {real, imag} */,
  {32'hc40b0e48, 32'h00000000} /* (1, 10, 17) {real, imag} */,
  {32'h4285dc48, 32'h00000000} /* (1, 10, 16) {real, imag} */,
  {32'hc44d58c4, 32'h00000000} /* (1, 10, 15) {real, imag} */,
  {32'hc39a8e70, 32'h00000000} /* (1, 10, 14) {real, imag} */,
  {32'h43df284a, 32'h00000000} /* (1, 10, 13) {real, imag} */,
  {32'hc3f7df14, 32'h00000000} /* (1, 10, 12) {real, imag} */,
  {32'hc3c9d78c, 32'h00000000} /* (1, 10, 11) {real, imag} */,
  {32'hc303f46c, 32'h00000000} /* (1, 10, 10) {real, imag} */,
  {32'hc488ff96, 32'h00000000} /* (1, 10, 9) {real, imag} */,
  {32'hc31e9137, 32'h00000000} /* (1, 10, 8) {real, imag} */,
  {32'hc3510763, 32'h00000000} /* (1, 10, 7) {real, imag} */,
  {32'h43bf6f1f, 32'h00000000} /* (1, 10, 6) {real, imag} */,
  {32'h4317dcda, 32'h00000000} /* (1, 10, 5) {real, imag} */,
  {32'h41e0d300, 32'h00000000} /* (1, 10, 4) {real, imag} */,
  {32'hc34962b2, 32'h00000000} /* (1, 10, 3) {real, imag} */,
  {32'hc470e0a2, 32'h00000000} /* (1, 10, 2) {real, imag} */,
  {32'hc423dcec, 32'h00000000} /* (1, 10, 1) {real, imag} */,
  {32'hc3542cf8, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'hc4a64c1e, 32'h00000000} /* (1, 9, 31) {real, imag} */,
  {32'hc4ddc6b3, 32'h00000000} /* (1, 9, 30) {real, imag} */,
  {32'hc481ec12, 32'h00000000} /* (1, 9, 29) {real, imag} */,
  {32'hc4d2b3a4, 32'h00000000} /* (1, 9, 28) {real, imag} */,
  {32'hc4db7866, 32'h00000000} /* (1, 9, 27) {real, imag} */,
  {32'hc511de8e, 32'h00000000} /* (1, 9, 26) {real, imag} */,
  {32'hc4fae56c, 32'h00000000} /* (1, 9, 25) {real, imag} */,
  {32'hc4ef92d6, 32'h00000000} /* (1, 9, 24) {real, imag} */,
  {32'hc5091859, 32'h00000000} /* (1, 9, 23) {real, imag} */,
  {32'hc4db3f65, 32'h00000000} /* (1, 9, 22) {real, imag} */,
  {32'hc4bcbb74, 32'h00000000} /* (1, 9, 21) {real, imag} */,
  {32'h441a341c, 32'h00000000} /* (1, 9, 20) {real, imag} */,
  {32'h44eafa9c, 32'h00000000} /* (1, 9, 19) {real, imag} */,
  {32'h4433e644, 32'h00000000} /* (1, 9, 18) {real, imag} */,
  {32'h4424988f, 32'h00000000} /* (1, 9, 17) {real, imag} */,
  {32'h44481c0a, 32'h00000000} /* (1, 9, 16) {real, imag} */,
  {32'h450a4728, 32'h00000000} /* (1, 9, 15) {real, imag} */,
  {32'h449749bd, 32'h00000000} /* (1, 9, 14) {real, imag} */,
  {32'h442d9d9f, 32'h00000000} /* (1, 9, 13) {real, imag} */,
  {32'h44b06f38, 32'h00000000} /* (1, 9, 12) {real, imag} */,
  {32'h449c2a22, 32'h00000000} /* (1, 9, 11) {real, imag} */,
  {32'hc40ee122, 32'h00000000} /* (1, 9, 10) {real, imag} */,
  {32'hc4c3646c, 32'h00000000} /* (1, 9, 9) {real, imag} */,
  {32'hc49a4db4, 32'h00000000} /* (1, 9, 8) {real, imag} */,
  {32'hc4d88986, 32'h00000000} /* (1, 9, 7) {real, imag} */,
  {32'hc40f877e, 32'h00000000} /* (1, 9, 6) {real, imag} */,
  {32'hc4ded5de, 32'h00000000} /* (1, 9, 5) {real, imag} */,
  {32'hc4a8bc84, 32'h00000000} /* (1, 9, 4) {real, imag} */,
  {32'hc4e9b73c, 32'h00000000} /* (1, 9, 3) {real, imag} */,
  {32'hc537e8b2, 32'h00000000} /* (1, 9, 2) {real, imag} */,
  {32'hc4d41a7c, 32'h00000000} /* (1, 9, 1) {real, imag} */,
  {32'hc4a9bd9b, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'hc4dd101f, 32'h00000000} /* (1, 8, 31) {real, imag} */,
  {32'hc4be42d0, 32'h00000000} /* (1, 8, 30) {real, imag} */,
  {32'hc50ffc11, 32'h00000000} /* (1, 8, 29) {real, imag} */,
  {32'hc4f1d06b, 32'h00000000} /* (1, 8, 28) {real, imag} */,
  {32'hc5025c81, 32'h00000000} /* (1, 8, 27) {real, imag} */,
  {32'hc5035aec, 32'h00000000} /* (1, 8, 26) {real, imag} */,
  {32'hc532b4d4, 32'h00000000} /* (1, 8, 25) {real, imag} */,
  {32'hc5501426, 32'h00000000} /* (1, 8, 24) {real, imag} */,
  {32'hc53157be, 32'h00000000} /* (1, 8, 23) {real, imag} */,
  {32'hc521d523, 32'h00000000} /* (1, 8, 22) {real, imag} */,
  {32'hc479da4b, 32'h00000000} /* (1, 8, 21) {real, imag} */,
  {32'h44457626, 32'h00000000} /* (1, 8, 20) {real, imag} */,
  {32'h44b5feb0, 32'h00000000} /* (1, 8, 19) {real, imag} */,
  {32'h444968ec, 32'h00000000} /* (1, 8, 18) {real, imag} */,
  {32'h44e6ed5f, 32'h00000000} /* (1, 8, 17) {real, imag} */,
  {32'h450bf8a6, 32'h00000000} /* (1, 8, 16) {real, imag} */,
  {32'h44e84129, 32'h00000000} /* (1, 8, 15) {real, imag} */,
  {32'h4511baad, 32'h00000000} /* (1, 8, 14) {real, imag} */,
  {32'h44c1c8c6, 32'h00000000} /* (1, 8, 13) {real, imag} */,
  {32'h44a4c97d, 32'h00000000} /* (1, 8, 12) {real, imag} */,
  {32'h4492408a, 32'h00000000} /* (1, 8, 11) {real, imag} */,
  {32'hc4a40898, 32'h00000000} /* (1, 8, 10) {real, imag} */,
  {32'hc4906bbe, 32'h00000000} /* (1, 8, 9) {real, imag} */,
  {32'hc484afb5, 32'h00000000} /* (1, 8, 8) {real, imag} */,
  {32'hc4d9d3dc, 32'h00000000} /* (1, 8, 7) {real, imag} */,
  {32'hc491fcf2, 32'h00000000} /* (1, 8, 6) {real, imag} */,
  {32'hc5001cd1, 32'h00000000} /* (1, 8, 5) {real, imag} */,
  {32'hc521ae06, 32'h00000000} /* (1, 8, 4) {real, imag} */,
  {32'hc4da603e, 32'h00000000} /* (1, 8, 3) {real, imag} */,
  {32'hc54fd3b3, 32'h00000000} /* (1, 8, 2) {real, imag} */,
  {32'hc50a67b0, 32'h00000000} /* (1, 8, 1) {real, imag} */,
  {32'hc48f2c38, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'hc4fcc2a4, 32'h00000000} /* (1, 7, 31) {real, imag} */,
  {32'hc5229e62, 32'h00000000} /* (1, 7, 30) {real, imag} */,
  {32'hc50f084e, 32'h00000000} /* (1, 7, 29) {real, imag} */,
  {32'hc54552b2, 32'h00000000} /* (1, 7, 28) {real, imag} */,
  {32'hc54e8007, 32'h00000000} /* (1, 7, 27) {real, imag} */,
  {32'hc56a1d9a, 32'h00000000} /* (1, 7, 26) {real, imag} */,
  {32'hc57eca1f, 32'h00000000} /* (1, 7, 25) {real, imag} */,
  {32'hc556843e, 32'h00000000} /* (1, 7, 24) {real, imag} */,
  {32'hc53ec36c, 32'h00000000} /* (1, 7, 23) {real, imag} */,
  {32'hc527ac40, 32'h00000000} /* (1, 7, 22) {real, imag} */,
  {32'hc38bd8dc, 32'h00000000} /* (1, 7, 21) {real, imag} */,
  {32'h4493459f, 32'h00000000} /* (1, 7, 20) {real, imag} */,
  {32'h448a4fca, 32'h00000000} /* (1, 7, 19) {real, imag} */,
  {32'h44d76541, 32'h00000000} /* (1, 7, 18) {real, imag} */,
  {32'h450ebafc, 32'h00000000} /* (1, 7, 17) {real, imag} */,
  {32'h4517efe4, 32'h00000000} /* (1, 7, 16) {real, imag} */,
  {32'h453fd37a, 32'h00000000} /* (1, 7, 15) {real, imag} */,
  {32'h453f5c8e, 32'h00000000} /* (1, 7, 14) {real, imag} */,
  {32'h45214320, 32'h00000000} /* (1, 7, 13) {real, imag} */,
  {32'h44eb78bc, 32'h00000000} /* (1, 7, 12) {real, imag} */,
  {32'h428a2260, 32'h00000000} /* (1, 7, 11) {real, imag} */,
  {32'hc45bbbca, 32'h00000000} /* (1, 7, 10) {real, imag} */,
  {32'hc4b5f092, 32'h00000000} /* (1, 7, 9) {real, imag} */,
  {32'hc495568c, 32'h00000000} /* (1, 7, 8) {real, imag} */,
  {32'hc4c0d1db, 32'h00000000} /* (1, 7, 7) {real, imag} */,
  {32'hc5006a1c, 32'h00000000} /* (1, 7, 6) {real, imag} */,
  {32'hc520b332, 32'h00000000} /* (1, 7, 5) {real, imag} */,
  {32'hc5540272, 32'h00000000} /* (1, 7, 4) {real, imag} */,
  {32'hc50a6b15, 32'h00000000} /* (1, 7, 3) {real, imag} */,
  {32'hc56e5d72, 32'h00000000} /* (1, 7, 2) {real, imag} */,
  {32'hc532c4e6, 32'h00000000} /* (1, 7, 1) {real, imag} */,
  {32'hc49cc47a, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'hc4e4daa1, 32'h00000000} /* (1, 6, 31) {real, imag} */,
  {32'hc5051662, 32'h00000000} /* (1, 6, 30) {real, imag} */,
  {32'hc534ae0c, 32'h00000000} /* (1, 6, 29) {real, imag} */,
  {32'hc54b11f7, 32'h00000000} /* (1, 6, 28) {real, imag} */,
  {32'hc5405c7c, 32'h00000000} /* (1, 6, 27) {real, imag} */,
  {32'hc58e4dfa, 32'h00000000} /* (1, 6, 26) {real, imag} */,
  {32'hc589cfa1, 32'h00000000} /* (1, 6, 25) {real, imag} */,
  {32'hc5562cbd, 32'h00000000} /* (1, 6, 24) {real, imag} */,
  {32'hc512187e, 32'h00000000} /* (1, 6, 23) {real, imag} */,
  {32'hc50a5a58, 32'h00000000} /* (1, 6, 22) {real, imag} */,
  {32'hc51b39c4, 32'h00000000} /* (1, 6, 21) {real, imag} */,
  {32'h44e4c868, 32'h00000000} /* (1, 6, 20) {real, imag} */,
  {32'h4433122a, 32'h00000000} /* (1, 6, 19) {real, imag} */,
  {32'h440d50f9, 32'h00000000} /* (1, 6, 18) {real, imag} */,
  {32'h44c63311, 32'h00000000} /* (1, 6, 17) {real, imag} */,
  {32'h451144e5, 32'h00000000} /* (1, 6, 16) {real, imag} */,
  {32'h45352832, 32'h00000000} /* (1, 6, 15) {real, imag} */,
  {32'h4518456c, 32'h00000000} /* (1, 6, 14) {real, imag} */,
  {32'h452d8f64, 32'h00000000} /* (1, 6, 13) {real, imag} */,
  {32'h451c80a1, 32'h00000000} /* (1, 6, 12) {real, imag} */,
  {32'h448a836d, 32'h00000000} /* (1, 6, 11) {real, imag} */,
  {32'h43418db0, 32'h00000000} /* (1, 6, 10) {real, imag} */,
  {32'hc507fc30, 32'h00000000} /* (1, 6, 9) {real, imag} */,
  {32'hc4ab3fba, 32'h00000000} /* (1, 6, 8) {real, imag} */,
  {32'hc48f2f8a, 32'h00000000} /* (1, 6, 7) {real, imag} */,
  {32'hc4b3e7d8, 32'h00000000} /* (1, 6, 6) {real, imag} */,
  {32'hc5022cc2, 32'h00000000} /* (1, 6, 5) {real, imag} */,
  {32'hc50a67bd, 32'h00000000} /* (1, 6, 4) {real, imag} */,
  {32'hc5254634, 32'h00000000} /* (1, 6, 3) {real, imag} */,
  {32'hc4f378b8, 32'h00000000} /* (1, 6, 2) {real, imag} */,
  {32'hc4d90ef1, 32'h00000000} /* (1, 6, 1) {real, imag} */,
  {32'hc4f3753a, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'hc5222772, 32'h00000000} /* (1, 5, 31) {real, imag} */,
  {32'hc552e7b8, 32'h00000000} /* (1, 5, 30) {real, imag} */,
  {32'hc550dfe6, 32'h00000000} /* (1, 5, 29) {real, imag} */,
  {32'hc56455da, 32'h00000000} /* (1, 5, 28) {real, imag} */,
  {32'hc542a0ee, 32'h00000000} /* (1, 5, 27) {real, imag} */,
  {32'hc597b74d, 32'h00000000} /* (1, 5, 26) {real, imag} */,
  {32'hc5615cf9, 32'h00000000} /* (1, 5, 25) {real, imag} */,
  {32'hc535f562, 32'h00000000} /* (1, 5, 24) {real, imag} */,
  {32'hc55512e2, 32'h00000000} /* (1, 5, 23) {real, imag} */,
  {32'hc556c2c8, 32'h00000000} /* (1, 5, 22) {real, imag} */,
  {32'hc510cd74, 32'h00000000} /* (1, 5, 21) {real, imag} */,
  {32'hc2d65450, 32'h00000000} /* (1, 5, 20) {real, imag} */,
  {32'hc40d022a, 32'h00000000} /* (1, 5, 19) {real, imag} */,
  {32'hc420bcb4, 32'h00000000} /* (1, 5, 18) {real, imag} */,
  {32'hc4661a78, 32'h00000000} /* (1, 5, 17) {real, imag} */,
  {32'h433309d4, 32'h00000000} /* (1, 5, 16) {real, imag} */,
  {32'h44650062, 32'h00000000} /* (1, 5, 15) {real, imag} */,
  {32'h449e2aab, 32'h00000000} /* (1, 5, 14) {real, imag} */,
  {32'h4517edc2, 32'h00000000} /* (1, 5, 13) {real, imag} */,
  {32'h453159ea, 32'h00000000} /* (1, 5, 12) {real, imag} */,
  {32'h45288092, 32'h00000000} /* (1, 5, 11) {real, imag} */,
  {32'h448abbcc, 32'h00000000} /* (1, 5, 10) {real, imag} */,
  {32'h4478f4ec, 32'h00000000} /* (1, 5, 9) {real, imag} */,
  {32'h433d60c0, 32'h00000000} /* (1, 5, 8) {real, imag} */,
  {32'h420621a0, 32'h00000000} /* (1, 5, 7) {real, imag} */,
  {32'hc3c936a4, 32'h00000000} /* (1, 5, 6) {real, imag} */,
  {32'hc43ec4f6, 32'h00000000} /* (1, 5, 5) {real, imag} */,
  {32'hc4f0eced, 32'h00000000} /* (1, 5, 4) {real, imag} */,
  {32'hc503ddaa, 32'h00000000} /* (1, 5, 3) {real, imag} */,
  {32'hc51d288f, 32'h00000000} /* (1, 5, 2) {real, imag} */,
  {32'hc519a10e, 32'h00000000} /* (1, 5, 1) {real, imag} */,
  {32'hc4f2fe0a, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'hc52e0498, 32'h00000000} /* (1, 4, 31) {real, imag} */,
  {32'hc5429e86, 32'h00000000} /* (1, 4, 30) {real, imag} */,
  {32'hc55e86d0, 32'h00000000} /* (1, 4, 29) {real, imag} */,
  {32'hc564f9b2, 32'h00000000} /* (1, 4, 28) {real, imag} */,
  {32'hc58401ba, 32'h00000000} /* (1, 4, 27) {real, imag} */,
  {32'hc580a25f, 32'h00000000} /* (1, 4, 26) {real, imag} */,
  {32'hc5889318, 32'h00000000} /* (1, 4, 25) {real, imag} */,
  {32'hc56664b7, 32'h00000000} /* (1, 4, 24) {real, imag} */,
  {32'hc53f9931, 32'h00000000} /* (1, 4, 23) {real, imag} */,
  {32'hc5149fa7, 32'h00000000} /* (1, 4, 22) {real, imag} */,
  {32'hc4c0b6e9, 32'h00000000} /* (1, 4, 21) {real, imag} */,
  {32'hc51c8cd9, 32'h00000000} /* (1, 4, 20) {real, imag} */,
  {32'hc5038fc4, 32'h00000000} /* (1, 4, 19) {real, imag} */,
  {32'hc497cc10, 32'h00000000} /* (1, 4, 18) {real, imag} */,
  {32'hc4f20fc5, 32'h00000000} /* (1, 4, 17) {real, imag} */,
  {32'hc4942869, 32'h00000000} /* (1, 4, 16) {real, imag} */,
  {32'h43eb5770, 32'h00000000} /* (1, 4, 15) {real, imag} */,
  {32'h44cd8751, 32'h00000000} /* (1, 4, 14) {real, imag} */,
  {32'h44e150f8, 32'h00000000} /* (1, 4, 13) {real, imag} */,
  {32'h4514d302, 32'h00000000} /* (1, 4, 12) {real, imag} */,
  {32'h451e4b98, 32'h00000000} /* (1, 4, 11) {real, imag} */,
  {32'h45126af8, 32'h00000000} /* (1, 4, 10) {real, imag} */,
  {32'h452c4ab8, 32'h00000000} /* (1, 4, 9) {real, imag} */,
  {32'h44d613ee, 32'h00000000} /* (1, 4, 8) {real, imag} */,
  {32'h44e40e5a, 32'h00000000} /* (1, 4, 7) {real, imag} */,
  {32'h446572a8, 32'h00000000} /* (1, 4, 6) {real, imag} */,
  {32'hc3fa1394, 32'h00000000} /* (1, 4, 5) {real, imag} */,
  {32'hc4cd5777, 32'h00000000} /* (1, 4, 4) {real, imag} */,
  {32'hc52f458a, 32'h00000000} /* (1, 4, 3) {real, imag} */,
  {32'hc54a20a4, 32'h00000000} /* (1, 4, 2) {real, imag} */,
  {32'hc5508752, 32'h00000000} /* (1, 4, 1) {real, imag} */,
  {32'hc508fcfc, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hc516c025, 32'h00000000} /* (1, 3, 31) {real, imag} */,
  {32'hc53e2986, 32'h00000000} /* (1, 3, 30) {real, imag} */,
  {32'hc55c7ad0, 32'h00000000} /* (1, 3, 29) {real, imag} */,
  {32'hc54b43de, 32'h00000000} /* (1, 3, 28) {real, imag} */,
  {32'hc56ee9ba, 32'h00000000} /* (1, 3, 27) {real, imag} */,
  {32'hc5676668, 32'h00000000} /* (1, 3, 26) {real, imag} */,
  {32'hc55525c2, 32'h00000000} /* (1, 3, 25) {real, imag} */,
  {32'hc57d6174, 32'h00000000} /* (1, 3, 24) {real, imag} */,
  {32'hc565e69b, 32'h00000000} /* (1, 3, 23) {real, imag} */,
  {32'hc51c6e52, 32'h00000000} /* (1, 3, 22) {real, imag} */,
  {32'hc51532e6, 32'h00000000} /* (1, 3, 21) {real, imag} */,
  {32'hc50880e9, 32'h00000000} /* (1, 3, 20) {real, imag} */,
  {32'hc5581399, 32'h00000000} /* (1, 3, 19) {real, imag} */,
  {32'hc54573ce, 32'h00000000} /* (1, 3, 18) {real, imag} */,
  {32'hc4e9d872, 32'h00000000} /* (1, 3, 17) {real, imag} */,
  {32'hc43ac8b4, 32'h00000000} /* (1, 3, 16) {real, imag} */,
  {32'h4448f0f7, 32'h00000000} /* (1, 3, 15) {real, imag} */,
  {32'h44f7a27f, 32'h00000000} /* (1, 3, 14) {real, imag} */,
  {32'h452a6750, 32'h00000000} /* (1, 3, 13) {real, imag} */,
  {32'h4522882e, 32'h00000000} /* (1, 3, 12) {real, imag} */,
  {32'h45390030, 32'h00000000} /* (1, 3, 11) {real, imag} */,
  {32'h456f942c, 32'h00000000} /* (1, 3, 10) {real, imag} */,
  {32'h4527bbbc, 32'h00000000} /* (1, 3, 9) {real, imag} */,
  {32'h44fedf99, 32'h00000000} /* (1, 3, 8) {real, imag} */,
  {32'h44fd0606, 32'h00000000} /* (1, 3, 7) {real, imag} */,
  {32'h4442a29a, 32'h00000000} /* (1, 3, 6) {real, imag} */,
  {32'hc4c08633, 32'h00000000} /* (1, 3, 5) {real, imag} */,
  {32'hc49debd1, 32'h00000000} /* (1, 3, 4) {real, imag} */,
  {32'hc525ce85, 32'h00000000} /* (1, 3, 3) {real, imag} */,
  {32'hc51e7bb8, 32'h00000000} /* (1, 3, 2) {real, imag} */,
  {32'hc4f69cd2, 32'h00000000} /* (1, 3, 1) {real, imag} */,
  {32'hc50efb86, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hc51930b6, 32'h00000000} /* (1, 2, 31) {real, imag} */,
  {32'hc552ca68, 32'h00000000} /* (1, 2, 30) {real, imag} */,
  {32'hc53d7e87, 32'h00000000} /* (1, 2, 29) {real, imag} */,
  {32'hc5896781, 32'h00000000} /* (1, 2, 28) {real, imag} */,
  {32'hc547526c, 32'h00000000} /* (1, 2, 27) {real, imag} */,
  {32'hc52daed5, 32'h00000000} /* (1, 2, 26) {real, imag} */,
  {32'hc55c5546, 32'h00000000} /* (1, 2, 25) {real, imag} */,
  {32'hc522bb27, 32'h00000000} /* (1, 2, 24) {real, imag} */,
  {32'hc5189c8c, 32'h00000000} /* (1, 2, 23) {real, imag} */,
  {32'hc5157436, 32'h00000000} /* (1, 2, 22) {real, imag} */,
  {32'hc4f6024a, 32'h00000000} /* (1, 2, 21) {real, imag} */,
  {32'hc4d0af62, 32'h00000000} /* (1, 2, 20) {real, imag} */,
  {32'hc5166e65, 32'h00000000} /* (1, 2, 19) {real, imag} */,
  {32'hc52d9a2a, 32'h00000000} /* (1, 2, 18) {real, imag} */,
  {32'hc50ec3c8, 32'h00000000} /* (1, 2, 17) {real, imag} */,
  {32'hc439e1f2, 32'h00000000} /* (1, 2, 16) {real, imag} */,
  {32'h447fd4f0, 32'h00000000} /* (1, 2, 15) {real, imag} */,
  {32'h45028d4c, 32'h00000000} /* (1, 2, 14) {real, imag} */,
  {32'h458cb77c, 32'h00000000} /* (1, 2, 13) {real, imag} */,
  {32'h4555e466, 32'h00000000} /* (1, 2, 12) {real, imag} */,
  {32'h4553abe0, 32'h00000000} /* (1, 2, 11) {real, imag} */,
  {32'h45613ecd, 32'h00000000} /* (1, 2, 10) {real, imag} */,
  {32'h4555b348, 32'h00000000} /* (1, 2, 9) {real, imag} */,
  {32'h451f8091, 32'h00000000} /* (1, 2, 8) {real, imag} */,
  {32'h44a6329f, 32'h00000000} /* (1, 2, 7) {real, imag} */,
  {32'h45051e04, 32'h00000000} /* (1, 2, 6) {real, imag} */,
  {32'hc443b804, 32'h00000000} /* (1, 2, 5) {real, imag} */,
  {32'hc5393c43, 32'h00000000} /* (1, 2, 4) {real, imag} */,
  {32'hc52fddab, 32'h00000000} /* (1, 2, 3) {real, imag} */,
  {32'hc51fbcde, 32'h00000000} /* (1, 2, 2) {real, imag} */,
  {32'hc5726856, 32'h00000000} /* (1, 2, 1) {real, imag} */,
  {32'hc5399d24, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hc500f771, 32'h00000000} /* (1, 1, 31) {real, imag} */,
  {32'hc526aa48, 32'h00000000} /* (1, 1, 30) {real, imag} */,
  {32'hc523095d, 32'h00000000} /* (1, 1, 29) {real, imag} */,
  {32'hc51fbc3e, 32'h00000000} /* (1, 1, 28) {real, imag} */,
  {32'hc509aea3, 32'h00000000} /* (1, 1, 27) {real, imag} */,
  {32'hc51b95de, 32'h00000000} /* (1, 1, 26) {real, imag} */,
  {32'hc51b0a28, 32'h00000000} /* (1, 1, 25) {real, imag} */,
  {32'hc51c2dbf, 32'h00000000} /* (1, 1, 24) {real, imag} */,
  {32'hc51e9efc, 32'h00000000} /* (1, 1, 23) {real, imag} */,
  {32'hc4df5bf6, 32'h00000000} /* (1, 1, 22) {real, imag} */,
  {32'hc49fcc4e, 32'h00000000} /* (1, 1, 21) {real, imag} */,
  {32'hc4b965c5, 32'h00000000} /* (1, 1, 20) {real, imag} */,
  {32'hc4d967e3, 32'h00000000} /* (1, 1, 19) {real, imag} */,
  {32'hc511a7b0, 32'h00000000} /* (1, 1, 18) {real, imag} */,
  {32'hc4a3a250, 32'h00000000} /* (1, 1, 17) {real, imag} */,
  {32'hc39c455c, 32'h00000000} /* (1, 1, 16) {real, imag} */,
  {32'h4483f032, 32'h00000000} /* (1, 1, 15) {real, imag} */,
  {32'h453285b6, 32'h00000000} /* (1, 1, 14) {real, imag} */,
  {32'h45862d6c, 32'h00000000} /* (1, 1, 13) {real, imag} */,
  {32'h45637fb6, 32'h00000000} /* (1, 1, 12) {real, imag} */,
  {32'h45657ee5, 32'h00000000} /* (1, 1, 11) {real, imag} */,
  {32'h452acd28, 32'h00000000} /* (1, 1, 10) {real, imag} */,
  {32'h4530b602, 32'h00000000} /* (1, 1, 9) {real, imag} */,
  {32'h451db5b9, 32'h00000000} /* (1, 1, 8) {real, imag} */,
  {32'h4508a5ac, 32'h00000000} /* (1, 1, 7) {real, imag} */,
  {32'h44a84d72, 32'h00000000} /* (1, 1, 6) {real, imag} */,
  {32'hc43276ac, 32'h00000000} /* (1, 1, 5) {real, imag} */,
  {32'hc576bcf2, 32'h00000000} /* (1, 1, 4) {real, imag} */,
  {32'hc53a389c, 32'h00000000} /* (1, 1, 3) {real, imag} */,
  {32'hc516f822, 32'h00000000} /* (1, 1, 2) {real, imag} */,
  {32'hc518277e, 32'h00000000} /* (1, 1, 1) {real, imag} */,
  {32'hc507d150, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hc4e73418, 32'h00000000} /* (1, 0, 31) {real, imag} */,
  {32'hc4d83004, 32'h00000000} /* (1, 0, 30) {real, imag} */,
  {32'hc4e21e35, 32'h00000000} /* (1, 0, 29) {real, imag} */,
  {32'hc4dd9686, 32'h00000000} /* (1, 0, 28) {real, imag} */,
  {32'hc4ec6542, 32'h00000000} /* (1, 0, 27) {real, imag} */,
  {32'hc5046ecd, 32'h00000000} /* (1, 0, 26) {real, imag} */,
  {32'hc4c5db91, 32'h00000000} /* (1, 0, 25) {real, imag} */,
  {32'hc4903f94, 32'h00000000} /* (1, 0, 24) {real, imag} */,
  {32'hc52d797a, 32'h00000000} /* (1, 0, 23) {real, imag} */,
  {32'hc4f948ac, 32'h00000000} /* (1, 0, 22) {real, imag} */,
  {32'hc42b8f8e, 32'h00000000} /* (1, 0, 21) {real, imag} */,
  {32'hc430650a, 32'h00000000} /* (1, 0, 20) {real, imag} */,
  {32'hc48042b2, 32'h00000000} /* (1, 0, 19) {real, imag} */,
  {32'hc46dd936, 32'h00000000} /* (1, 0, 18) {real, imag} */,
  {32'h431d6ca8, 32'h00000000} /* (1, 0, 17) {real, imag} */,
  {32'h43a96d38, 32'h00000000} /* (1, 0, 16) {real, imag} */,
  {32'h4496c812, 32'h00000000} /* (1, 0, 15) {real, imag} */,
  {32'h451cda52, 32'h00000000} /* (1, 0, 14) {real, imag} */,
  {32'h451c0103, 32'h00000000} /* (1, 0, 13) {real, imag} */,
  {32'h4507774a, 32'h00000000} /* (1, 0, 12) {real, imag} */,
  {32'h451765e9, 32'h00000000} /* (1, 0, 11) {real, imag} */,
  {32'h45197cf3, 32'h00000000} /* (1, 0, 10) {real, imag} */,
  {32'h44badc1d, 32'h00000000} /* (1, 0, 9) {real, imag} */,
  {32'h44802622, 32'h00000000} /* (1, 0, 8) {real, imag} */,
  {32'h44b3070f, 32'h00000000} /* (1, 0, 7) {real, imag} */,
  {32'h4384746e, 32'h00000000} /* (1, 0, 6) {real, imag} */,
  {32'hc48a1a5d, 32'h00000000} /* (1, 0, 5) {real, imag} */,
  {32'hc4abcc25, 32'h00000000} /* (1, 0, 4) {real, imag} */,
  {32'hc51010af, 32'h00000000} /* (1, 0, 3) {real, imag} */,
  {32'hc51648c0, 32'h00000000} /* (1, 0, 2) {real, imag} */,
  {32'hc4fdebc3, 32'h00000000} /* (1, 0, 1) {real, imag} */,
  {32'hc4e6d2e0, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hc419ef60, 32'h00000000} /* (0, 31, 31) {real, imag} */,
  {32'hc429c344, 32'h00000000} /* (0, 31, 30) {real, imag} */,
  {32'hc4e86658, 32'h00000000} /* (0, 31, 29) {real, imag} */,
  {32'hc50abf84, 32'h00000000} /* (0, 31, 28) {real, imag} */,
  {32'hc44caf0a, 32'h00000000} /* (0, 31, 27) {real, imag} */,
  {32'hc412a5f9, 32'h00000000} /* (0, 31, 26) {real, imag} */,
  {32'hc3f09df0, 32'h00000000} /* (0, 31, 25) {real, imag} */,
  {32'hc38a8780, 32'h00000000} /* (0, 31, 24) {real, imag} */,
  {32'hc40598ff, 32'h00000000} /* (0, 31, 23) {real, imag} */,
  {32'hc3bebe27, 32'h00000000} /* (0, 31, 22) {real, imag} */,
  {32'hc225c078, 32'h00000000} /* (0, 31, 21) {real, imag} */,
  {32'h4357e800, 32'h00000000} /* (0, 31, 20) {real, imag} */,
  {32'h439ce662, 32'h00000000} /* (0, 31, 19) {real, imag} */,
  {32'hc090f700, 32'h00000000} /* (0, 31, 18) {real, imag} */,
  {32'h42ea0880, 32'h00000000} /* (0, 31, 17) {real, imag} */,
  {32'h433f8c96, 32'h00000000} /* (0, 31, 16) {real, imag} */,
  {32'h43bdb315, 32'h00000000} /* (0, 31, 15) {real, imag} */,
  {32'h447de2bc, 32'h00000000} /* (0, 31, 14) {real, imag} */,
  {32'h4418f71c, 32'h00000000} /* (0, 31, 13) {real, imag} */,
  {32'h43eee2be, 32'h00000000} /* (0, 31, 12) {real, imag} */,
  {32'h446e6c8a, 32'h00000000} /* (0, 31, 11) {real, imag} */,
  {32'h43e2a896, 32'h00000000} /* (0, 31, 10) {real, imag} */,
  {32'h432fdb21, 32'h00000000} /* (0, 31, 9) {real, imag} */,
  {32'hc32e618f, 32'h00000000} /* (0, 31, 8) {real, imag} */,
  {32'hc2d9843e, 32'h00000000} /* (0, 31, 7) {real, imag} */,
  {32'hc3b35cf1, 32'h00000000} /* (0, 31, 6) {real, imag} */,
  {32'hc462b74c, 32'h00000000} /* (0, 31, 5) {real, imag} */,
  {32'hc47eae56, 32'h00000000} /* (0, 31, 4) {real, imag} */,
  {32'hc4798633, 32'h00000000} /* (0, 31, 3) {real, imag} */,
  {32'hc42de936, 32'h00000000} /* (0, 31, 2) {real, imag} */,
  {32'hc4318f78, 32'h00000000} /* (0, 31, 1) {real, imag} */,
  {32'hc43c5580, 32'h00000000} /* (0, 31, 0) {real, imag} */,
  {32'hc4a25a02, 32'h00000000} /* (0, 30, 31) {real, imag} */,
  {32'hc4135638, 32'h00000000} /* (0, 30, 30) {real, imag} */,
  {32'hc4c4c1c8, 32'h00000000} /* (0, 30, 29) {real, imag} */,
  {32'hc4f68a91, 32'h00000000} /* (0, 30, 28) {real, imag} */,
  {32'hc4a306be, 32'h00000000} /* (0, 30, 27) {real, imag} */,
  {32'hc419a5da, 32'h00000000} /* (0, 30, 26) {real, imag} */,
  {32'hc4357aa0, 32'h00000000} /* (0, 30, 25) {real, imag} */,
  {32'hc4907e2b, 32'h00000000} /* (0, 30, 24) {real, imag} */,
  {32'hc43bda44, 32'h00000000} /* (0, 30, 23) {real, imag} */,
  {32'hc36b4e32, 32'h00000000} /* (0, 30, 22) {real, imag} */,
  {32'hc1fd37e0, 32'h00000000} /* (0, 30, 21) {real, imag} */,
  {32'h442d7e9a, 32'h00000000} /* (0, 30, 20) {real, imag} */,
  {32'h443c63b5, 32'h00000000} /* (0, 30, 19) {real, imag} */,
  {32'h43986398, 32'h00000000} /* (0, 30, 18) {real, imag} */,
  {32'h443b1ba0, 32'h00000000} /* (0, 30, 17) {real, imag} */,
  {32'h44961366, 32'h00000000} /* (0, 30, 16) {real, imag} */,
  {32'h44263aaa, 32'h00000000} /* (0, 30, 15) {real, imag} */,
  {32'h4464f26a, 32'h00000000} /* (0, 30, 14) {real, imag} */,
  {32'h43f3042a, 32'h00000000} /* (0, 30, 13) {real, imag} */,
  {32'h43d15884, 32'h00000000} /* (0, 30, 12) {real, imag} */,
  {32'h43d738be, 32'h00000000} /* (0, 30, 11) {real, imag} */,
  {32'hc32f5a9e, 32'h00000000} /* (0, 30, 10) {real, imag} */,
  {32'hc1652c60, 32'h00000000} /* (0, 30, 9) {real, imag} */,
  {32'hc42ecec4, 32'h00000000} /* (0, 30, 8) {real, imag} */,
  {32'hc4355e60, 32'h00000000} /* (0, 30, 7) {real, imag} */,
  {32'hc4248728, 32'h00000000} /* (0, 30, 6) {real, imag} */,
  {32'hc4d324da, 32'h00000000} /* (0, 30, 5) {real, imag} */,
  {32'hc4cb6bbd, 32'h00000000} /* (0, 30, 4) {real, imag} */,
  {32'hc4aa96c8, 32'h00000000} /* (0, 30, 3) {real, imag} */,
  {32'hc4a7e5a2, 32'h00000000} /* (0, 30, 2) {real, imag} */,
  {32'hc38916f5, 32'h00000000} /* (0, 30, 1) {real, imag} */,
  {32'hc3dbabba, 32'h00000000} /* (0, 30, 0) {real, imag} */,
  {32'hc4b26de2, 32'h00000000} /* (0, 29, 31) {real, imag} */,
  {32'hc46957b4, 32'h00000000} /* (0, 29, 30) {real, imag} */,
  {32'hc4cdfcdf, 32'h00000000} /* (0, 29, 29) {real, imag} */,
  {32'hc4c5dfb2, 32'h00000000} /* (0, 29, 28) {real, imag} */,
  {32'hc46202f6, 32'h00000000} /* (0, 29, 27) {real, imag} */,
  {32'hc482fcbc, 32'h00000000} /* (0, 29, 26) {real, imag} */,
  {32'hc48a574a, 32'h00000000} /* (0, 29, 25) {real, imag} */,
  {32'hc49ded23, 32'h00000000} /* (0, 29, 24) {real, imag} */,
  {32'hc45ab0b3, 32'h00000000} /* (0, 29, 23) {real, imag} */,
  {32'hc39e7db7, 32'h00000000} /* (0, 29, 22) {real, imag} */,
  {32'hc28ce878, 32'h00000000} /* (0, 29, 21) {real, imag} */,
  {32'h442f55d0, 32'h00000000} /* (0, 29, 20) {real, imag} */,
  {32'h441b5f9c, 32'h00000000} /* (0, 29, 19) {real, imag} */,
  {32'h4473196d, 32'h00000000} /* (0, 29, 18) {real, imag} */,
  {32'h44b3bde2, 32'h00000000} /* (0, 29, 17) {real, imag} */,
  {32'h44c896ec, 32'h00000000} /* (0, 29, 16) {real, imag} */,
  {32'h444d3bfc, 32'h00000000} /* (0, 29, 15) {real, imag} */,
  {32'h44afed7a, 32'h00000000} /* (0, 29, 14) {real, imag} */,
  {32'h4488f2af, 32'h00000000} /* (0, 29, 13) {real, imag} */,
  {32'h444267ec, 32'h00000000} /* (0, 29, 12) {real, imag} */,
  {32'h4460b306, 32'h00000000} /* (0, 29, 11) {real, imag} */,
  {32'hc3ad04dd, 32'h00000000} /* (0, 29, 10) {real, imag} */,
  {32'hc4860822, 32'h00000000} /* (0, 29, 9) {real, imag} */,
  {32'hc44bbc2e, 32'h00000000} /* (0, 29, 8) {real, imag} */,
  {32'hc499dfc6, 32'h00000000} /* (0, 29, 7) {real, imag} */,
  {32'hc4952afc, 32'h00000000} /* (0, 29, 6) {real, imag} */,
  {32'hc4bc34dc, 32'h00000000} /* (0, 29, 5) {real, imag} */,
  {32'hc49cd45a, 32'h00000000} /* (0, 29, 4) {real, imag} */,
  {32'hc4937b60, 32'h00000000} /* (0, 29, 3) {real, imag} */,
  {32'hc4a4be44, 32'h00000000} /* (0, 29, 2) {real, imag} */,
  {32'hc4316229, 32'h00000000} /* (0, 29, 1) {real, imag} */,
  {32'hc46aec74, 32'h00000000} /* (0, 29, 0) {real, imag} */,
  {32'hc48f38bf, 32'h00000000} /* (0, 28, 31) {real, imag} */,
  {32'hc4cdf25f, 32'h00000000} /* (0, 28, 30) {real, imag} */,
  {32'hc4ea83cd, 32'h00000000} /* (0, 28, 29) {real, imag} */,
  {32'hc4d03246, 32'h00000000} /* (0, 28, 28) {real, imag} */,
  {32'hc3dd7e1c, 32'h00000000} /* (0, 28, 27) {real, imag} */,
  {32'hc46ca761, 32'h00000000} /* (0, 28, 26) {real, imag} */,
  {32'hc43e57c8, 32'h00000000} /* (0, 28, 25) {real, imag} */,
  {32'hc3c8931b, 32'h00000000} /* (0, 28, 24) {real, imag} */,
  {32'hc4550537, 32'h00000000} /* (0, 28, 23) {real, imag} */,
  {32'hc4055a73, 32'h00000000} /* (0, 28, 22) {real, imag} */,
  {32'hc1aad680, 32'h00000000} /* (0, 28, 21) {real, imag} */,
  {32'h447500f3, 32'h00000000} /* (0, 28, 20) {real, imag} */,
  {32'h44e4eab8, 32'h00000000} /* (0, 28, 19) {real, imag} */,
  {32'h44e18812, 32'h00000000} /* (0, 28, 18) {real, imag} */,
  {32'h44a20e8b, 32'h00000000} /* (0, 28, 17) {real, imag} */,
  {32'h44a5969c, 32'h00000000} /* (0, 28, 16) {real, imag} */,
  {32'h447931ca, 32'h00000000} /* (0, 28, 15) {real, imag} */,
  {32'h4473c41e, 32'h00000000} /* (0, 28, 14) {real, imag} */,
  {32'h44801c85, 32'h00000000} /* (0, 28, 13) {real, imag} */,
  {32'h44a4a686, 32'h00000000} /* (0, 28, 12) {real, imag} */,
  {32'h4468975a, 32'h00000000} /* (0, 28, 11) {real, imag} */,
  {32'hc3d59bb2, 32'h00000000} /* (0, 28, 10) {real, imag} */,
  {32'hc449b2cc, 32'h00000000} /* (0, 28, 9) {real, imag} */,
  {32'hc47c2376, 32'h00000000} /* (0, 28, 8) {real, imag} */,
  {32'hc4158379, 32'h00000000} /* (0, 28, 7) {real, imag} */,
  {32'hc467757d, 32'h00000000} /* (0, 28, 6) {real, imag} */,
  {32'hc4e08774, 32'h00000000} /* (0, 28, 5) {real, imag} */,
  {32'hc4809cb0, 32'h00000000} /* (0, 28, 4) {real, imag} */,
  {32'hc4b420e8, 32'h00000000} /* (0, 28, 3) {real, imag} */,
  {32'hc49a257a, 32'h00000000} /* (0, 28, 2) {real, imag} */,
  {32'hc486525b, 32'h00000000} /* (0, 28, 1) {real, imag} */,
  {32'hc48f8a6c, 32'h00000000} /* (0, 28, 0) {real, imag} */,
  {32'hc486e01a, 32'h00000000} /* (0, 27, 31) {real, imag} */,
  {32'hc4d5f17c, 32'h00000000} /* (0, 27, 30) {real, imag} */,
  {32'hc4c7c71a, 32'h00000000} /* (0, 27, 29) {real, imag} */,
  {32'hc4ce5088, 32'h00000000} /* (0, 27, 28) {real, imag} */,
  {32'hc4738ec6, 32'h00000000} /* (0, 27, 27) {real, imag} */,
  {32'hc48b4746, 32'h00000000} /* (0, 27, 26) {real, imag} */,
  {32'hc452467c, 32'h00000000} /* (0, 27, 25) {real, imag} */,
  {32'hc429e613, 32'h00000000} /* (0, 27, 24) {real, imag} */,
  {32'hc48293de, 32'h00000000} /* (0, 27, 23) {real, imag} */,
  {32'hc42b8dc8, 32'h00000000} /* (0, 27, 22) {real, imag} */,
  {32'h43b3d17e, 32'h00000000} /* (0, 27, 21) {real, imag} */,
  {32'h44960b80, 32'h00000000} /* (0, 27, 20) {real, imag} */,
  {32'h44843cf4, 32'h00000000} /* (0, 27, 19) {real, imag} */,
  {32'h44d993c4, 32'h00000000} /* (0, 27, 18) {real, imag} */,
  {32'h4502b2d4, 32'h00000000} /* (0, 27, 17) {real, imag} */,
  {32'h4469d739, 32'h00000000} /* (0, 27, 16) {real, imag} */,
  {32'h44781840, 32'h00000000} /* (0, 27, 15) {real, imag} */,
  {32'h444e9809, 32'h00000000} /* (0, 27, 14) {real, imag} */,
  {32'h445cc421, 32'h00000000} /* (0, 27, 13) {real, imag} */,
  {32'h4441de58, 32'h00000000} /* (0, 27, 12) {real, imag} */,
  {32'h444f9d0a, 32'h00000000} /* (0, 27, 11) {real, imag} */,
  {32'hc21f8cd0, 32'h00000000} /* (0, 27, 10) {real, imag} */,
  {32'hc20b71f8, 32'h00000000} /* (0, 27, 9) {real, imag} */,
  {32'hc44678c3, 32'h00000000} /* (0, 27, 8) {real, imag} */,
  {32'hc3e2e1af, 32'h00000000} /* (0, 27, 7) {real, imag} */,
  {32'hc448f48a, 32'h00000000} /* (0, 27, 6) {real, imag} */,
  {32'hc48924e0, 32'h00000000} /* (0, 27, 5) {real, imag} */,
  {32'hc4b71956, 32'h00000000} /* (0, 27, 4) {real, imag} */,
  {32'hc4720588, 32'h00000000} /* (0, 27, 3) {real, imag} */,
  {32'hc4680630, 32'h00000000} /* (0, 27, 2) {real, imag} */,
  {32'hc498bbe8, 32'h00000000} /* (0, 27, 1) {real, imag} */,
  {32'hc49f0630, 32'h00000000} /* (0, 27, 0) {real, imag} */,
  {32'hc4b569dc, 32'h00000000} /* (0, 26, 31) {real, imag} */,
  {32'hc51557f2, 32'h00000000} /* (0, 26, 30) {real, imag} */,
  {32'hc4fe908b, 32'h00000000} /* (0, 26, 29) {real, imag} */,
  {32'hc4911c7d, 32'h00000000} /* (0, 26, 28) {real, imag} */,
  {32'hc480c5fa, 32'h00000000} /* (0, 26, 27) {real, imag} */,
  {32'hc4a651e4, 32'h00000000} /* (0, 26, 26) {real, imag} */,
  {32'hc475153e, 32'h00000000} /* (0, 26, 25) {real, imag} */,
  {32'hc42ca317, 32'h00000000} /* (0, 26, 24) {real, imag} */,
  {32'hc4902f91, 32'h00000000} /* (0, 26, 23) {real, imag} */,
  {32'hc41c8e45, 32'h00000000} /* (0, 26, 22) {real, imag} */,
  {32'h4398da44, 32'h00000000} /* (0, 26, 21) {real, imag} */,
  {32'h44a779c5, 32'h00000000} /* (0, 26, 20) {real, imag} */,
  {32'h45094e99, 32'h00000000} /* (0, 26, 19) {real, imag} */,
  {32'h44fd9206, 32'h00000000} /* (0, 26, 18) {real, imag} */,
  {32'h44b2d656, 32'h00000000} /* (0, 26, 17) {real, imag} */,
  {32'h448b2af5, 32'h00000000} /* (0, 26, 16) {real, imag} */,
  {32'h44a9c208, 32'h00000000} /* (0, 26, 15) {real, imag} */,
  {32'h44b350e6, 32'h00000000} /* (0, 26, 14) {real, imag} */,
  {32'h4451b2ba, 32'h00000000} /* (0, 26, 13) {real, imag} */,
  {32'h4449eb03, 32'h00000000} /* (0, 26, 12) {real, imag} */,
  {32'h44a57b36, 32'h00000000} /* (0, 26, 11) {real, imag} */,
  {32'h421d80f0, 32'h00000000} /* (0, 26, 10) {real, imag} */,
  {32'hc47b2a5a, 32'h00000000} /* (0, 26, 9) {real, imag} */,
  {32'hc42579d1, 32'h00000000} /* (0, 26, 8) {real, imag} */,
  {32'hc40b70aa, 32'h00000000} /* (0, 26, 7) {real, imag} */,
  {32'hc47ceaad, 32'h00000000} /* (0, 26, 6) {real, imag} */,
  {32'hc4452d2a, 32'h00000000} /* (0, 26, 5) {real, imag} */,
  {32'hc468f07e, 32'h00000000} /* (0, 26, 4) {real, imag} */,
  {32'hc4b5151d, 32'h00000000} /* (0, 26, 3) {real, imag} */,
  {32'hc4ac4716, 32'h00000000} /* (0, 26, 2) {real, imag} */,
  {32'hc4cba0e4, 32'h00000000} /* (0, 26, 1) {real, imag} */,
  {32'hc4a7e665, 32'h00000000} /* (0, 26, 0) {real, imag} */,
  {32'hc4855598, 32'h00000000} /* (0, 25, 31) {real, imag} */,
  {32'hc50851ad, 32'h00000000} /* (0, 25, 30) {real, imag} */,
  {32'hc51ad650, 32'h00000000} /* (0, 25, 29) {real, imag} */,
  {32'hc4c10422, 32'h00000000} /* (0, 25, 28) {real, imag} */,
  {32'hc43bafde, 32'h00000000} /* (0, 25, 27) {real, imag} */,
  {32'hc469a366, 32'h00000000} /* (0, 25, 26) {real, imag} */,
  {32'hc43e93eb, 32'h00000000} /* (0, 25, 25) {real, imag} */,
  {32'hc368ab08, 32'h00000000} /* (0, 25, 24) {real, imag} */,
  {32'hc33115c0, 32'h00000000} /* (0, 25, 23) {real, imag} */,
  {32'hc318daea, 32'h00000000} /* (0, 25, 22) {real, imag} */,
  {32'h44217e7c, 32'h00000000} /* (0, 25, 21) {real, imag} */,
  {32'h45013c28, 32'h00000000} /* (0, 25, 20) {real, imag} */,
  {32'h45467b02, 32'h00000000} /* (0, 25, 19) {real, imag} */,
  {32'h450e628b, 32'h00000000} /* (0, 25, 18) {real, imag} */,
  {32'h44af0f22, 32'h00000000} /* (0, 25, 17) {real, imag} */,
  {32'h45144529, 32'h00000000} /* (0, 25, 16) {real, imag} */,
  {32'h44d2a6ba, 32'h00000000} /* (0, 25, 15) {real, imag} */,
  {32'h44718648, 32'h00000000} /* (0, 25, 14) {real, imag} */,
  {32'h4455bd6a, 32'h00000000} /* (0, 25, 13) {real, imag} */,
  {32'h44834222, 32'h00000000} /* (0, 25, 12) {real, imag} */,
  {32'h433a203a, 32'h00000000} /* (0, 25, 11) {real, imag} */,
  {32'hc368203a, 32'h00000000} /* (0, 25, 10) {real, imag} */,
  {32'hc50c5679, 32'h00000000} /* (0, 25, 9) {real, imag} */,
  {32'hc50ae132, 32'h00000000} /* (0, 25, 8) {real, imag} */,
  {32'hc4a693a2, 32'h00000000} /* (0, 25, 7) {real, imag} */,
  {32'hc39cbd59, 32'h00000000} /* (0, 25, 6) {real, imag} */,
  {32'hc44b6ade, 32'h00000000} /* (0, 25, 5) {real, imag} */,
  {32'hc4a84c58, 32'h00000000} /* (0, 25, 4) {real, imag} */,
  {32'hc4dc0028, 32'h00000000} /* (0, 25, 3) {real, imag} */,
  {32'hc4d8aa74, 32'h00000000} /* (0, 25, 2) {real, imag} */,
  {32'hc4fbb3f0, 32'h00000000} /* (0, 25, 1) {real, imag} */,
  {32'hc4d0e97f, 32'h00000000} /* (0, 25, 0) {real, imag} */,
  {32'hc474fde1, 32'h00000000} /* (0, 24, 31) {real, imag} */,
  {32'hc4899550, 32'h00000000} /* (0, 24, 30) {real, imag} */,
  {32'hc48516d2, 32'h00000000} /* (0, 24, 29) {real, imag} */,
  {32'hc4624cad, 32'h00000000} /* (0, 24, 28) {real, imag} */,
  {32'hc48016ca, 32'h00000000} /* (0, 24, 27) {real, imag} */,
  {32'hc4534d2d, 32'h00000000} /* (0, 24, 26) {real, imag} */,
  {32'hc3f1437a, 32'h00000000} /* (0, 24, 25) {real, imag} */,
  {32'hc3e0606c, 32'h00000000} /* (0, 24, 24) {real, imag} */,
  {32'h422829ac, 32'h00000000} /* (0, 24, 23) {real, imag} */,
  {32'h42e3364a, 32'h00000000} /* (0, 24, 22) {real, imag} */,
  {32'h43db58e2, 32'h00000000} /* (0, 24, 21) {real, imag} */,
  {32'h44e43351, 32'h00000000} /* (0, 24, 20) {real, imag} */,
  {32'h44da6bd8, 32'h00000000} /* (0, 24, 19) {real, imag} */,
  {32'h44ded263, 32'h00000000} /* (0, 24, 18) {real, imag} */,
  {32'h44a4ddc0, 32'h00000000} /* (0, 24, 17) {real, imag} */,
  {32'h44b8b0d1, 32'h00000000} /* (0, 24, 16) {real, imag} */,
  {32'h443b9abf, 32'h00000000} /* (0, 24, 15) {real, imag} */,
  {32'h44c2d204, 32'h00000000} /* (0, 24, 14) {real, imag} */,
  {32'h44ea4d66, 32'h00000000} /* (0, 24, 13) {real, imag} */,
  {32'h4425f90d, 32'h00000000} /* (0, 24, 12) {real, imag} */,
  {32'h442d7104, 32'h00000000} /* (0, 24, 11) {real, imag} */,
  {32'hc293cc38, 32'h00000000} /* (0, 24, 10) {real, imag} */,
  {32'hc457353f, 32'h00000000} /* (0, 24, 9) {real, imag} */,
  {32'hc4c71d45, 32'h00000000} /* (0, 24, 8) {real, imag} */,
  {32'hc3b5bba0, 32'h00000000} /* (0, 24, 7) {real, imag} */,
  {32'hc3c5aa94, 32'h00000000} /* (0, 24, 6) {real, imag} */,
  {32'hc4201e33, 32'h00000000} /* (0, 24, 5) {real, imag} */,
  {32'hc3c66404, 32'h00000000} /* (0, 24, 4) {real, imag} */,
  {32'hc44fe9f8, 32'h00000000} /* (0, 24, 3) {real, imag} */,
  {32'hc4a13147, 32'h00000000} /* (0, 24, 2) {real, imag} */,
  {32'hc492d9d2, 32'h00000000} /* (0, 24, 1) {real, imag} */,
  {32'hc4ad20c1, 32'h00000000} /* (0, 24, 0) {real, imag} */,
  {32'hc449cc6d, 32'h00000000} /* (0, 23, 31) {real, imag} */,
  {32'hc4a6b2f4, 32'h00000000} /* (0, 23, 30) {real, imag} */,
  {32'hc463a5f7, 32'h00000000} /* (0, 23, 29) {real, imag} */,
  {32'hc4c6b632, 32'h00000000} /* (0, 23, 28) {real, imag} */,
  {32'hc4994310, 32'h00000000} /* (0, 23, 27) {real, imag} */,
  {32'hc4b01c19, 32'h00000000} /* (0, 23, 26) {real, imag} */,
  {32'hc31b3a77, 32'h00000000} /* (0, 23, 25) {real, imag} */,
  {32'h41a6d3b8, 32'h00000000} /* (0, 23, 24) {real, imag} */,
  {32'h4279adc8, 32'h00000000} /* (0, 23, 23) {real, imag} */,
  {32'hc2d6eb2e, 32'h00000000} /* (0, 23, 22) {real, imag} */,
  {32'h4463be5a, 32'h00000000} /* (0, 23, 21) {real, imag} */,
  {32'h44decc04, 32'h00000000} /* (0, 23, 20) {real, imag} */,
  {32'h44a8d35e, 32'h00000000} /* (0, 23, 19) {real, imag} */,
  {32'h449d5a60, 32'h00000000} /* (0, 23, 18) {real, imag} */,
  {32'h44598da5, 32'h00000000} /* (0, 23, 17) {real, imag} */,
  {32'h4480ab38, 32'h00000000} /* (0, 23, 16) {real, imag} */,
  {32'h444fddff, 32'h00000000} /* (0, 23, 15) {real, imag} */,
  {32'h448799e6, 32'h00000000} /* (0, 23, 14) {real, imag} */,
  {32'h44866485, 32'h00000000} /* (0, 23, 13) {real, imag} */,
  {32'h44b5be8c, 32'h00000000} /* (0, 23, 12) {real, imag} */,
  {32'h4472387b, 32'h00000000} /* (0, 23, 11) {real, imag} */,
  {32'hc26451a0, 32'h00000000} /* (0, 23, 10) {real, imag} */,
  {32'hc3084271, 32'h00000000} /* (0, 23, 9) {real, imag} */,
  {32'hc3892de2, 32'h00000000} /* (0, 23, 8) {real, imag} */,
  {32'hc3e8f6f3, 32'h00000000} /* (0, 23, 7) {real, imag} */,
  {32'hc3373e9b, 32'h00000000} /* (0, 23, 6) {real, imag} */,
  {32'hc3a2e9a9, 32'h00000000} /* (0, 23, 5) {real, imag} */,
  {32'hc4609974, 32'h00000000} /* (0, 23, 4) {real, imag} */,
  {32'hc40cf38d, 32'h00000000} /* (0, 23, 3) {real, imag} */,
  {32'hc43850f2, 32'h00000000} /* (0, 23, 2) {real, imag} */,
  {32'hc45c78b7, 32'h00000000} /* (0, 23, 1) {real, imag} */,
  {32'hc4377faa, 32'h00000000} /* (0, 23, 0) {real, imag} */,
  {32'hc41b2308, 32'h00000000} /* (0, 22, 31) {real, imag} */,
  {32'hc41683e3, 32'h00000000} /* (0, 22, 30) {real, imag} */,
  {32'hc47c936a, 32'h00000000} /* (0, 22, 29) {real, imag} */,
  {32'hc4acb460, 32'h00000000} /* (0, 22, 28) {real, imag} */,
  {32'hc4cd5e50, 32'h00000000} /* (0, 22, 27) {real, imag} */,
  {32'hc4778f6a, 32'h00000000} /* (0, 22, 26) {real, imag} */,
  {32'hc40a7aca, 32'h00000000} /* (0, 22, 25) {real, imag} */,
  {32'hc394061f, 32'h00000000} /* (0, 22, 24) {real, imag} */,
  {32'hc397257e, 32'h00000000} /* (0, 22, 23) {real, imag} */,
  {32'hc1dff8c8, 32'h00000000} /* (0, 22, 22) {real, imag} */,
  {32'h442efa56, 32'h00000000} /* (0, 22, 21) {real, imag} */,
  {32'h44820e01, 32'h00000000} /* (0, 22, 20) {real, imag} */,
  {32'h44904079, 32'h00000000} /* (0, 22, 19) {real, imag} */,
  {32'h441448ce, 32'h00000000} /* (0, 22, 18) {real, imag} */,
  {32'h43f345d7, 32'h00000000} /* (0, 22, 17) {real, imag} */,
  {32'h445a0e58, 32'h00000000} /* (0, 22, 16) {real, imag} */,
  {32'h44621e92, 32'h00000000} /* (0, 22, 15) {real, imag} */,
  {32'h43e9d2ba, 32'h00000000} /* (0, 22, 14) {real, imag} */,
  {32'h44f3d87b, 32'h00000000} /* (0, 22, 13) {real, imag} */,
  {32'h44d67876, 32'h00000000} /* (0, 22, 12) {real, imag} */,
  {32'h4496b550, 32'h00000000} /* (0, 22, 11) {real, imag} */,
  {32'h43b08c4d, 32'h00000000} /* (0, 22, 10) {real, imag} */,
  {32'hc40aaccc, 32'h00000000} /* (0, 22, 9) {real, imag} */,
  {32'hc2c4743c, 32'h00000000} /* (0, 22, 8) {real, imag} */,
  {32'hc397c2aa, 32'h00000000} /* (0, 22, 7) {real, imag} */,
  {32'hc39cce18, 32'h00000000} /* (0, 22, 6) {real, imag} */,
  {32'hc36568be, 32'h00000000} /* (0, 22, 5) {real, imag} */,
  {32'hc427da1a, 32'h00000000} /* (0, 22, 4) {real, imag} */,
  {32'h4197b300, 32'h00000000} /* (0, 22, 3) {real, imag} */,
  {32'hc45b2f32, 32'h00000000} /* (0, 22, 2) {real, imag} */,
  {32'hc3e57d2f, 32'h00000000} /* (0, 22, 1) {real, imag} */,
  {32'hc429a466, 32'h00000000} /* (0, 22, 0) {real, imag} */,
  {32'hc3ea89b1, 32'h00000000} /* (0, 21, 31) {real, imag} */,
  {32'hc3fc696c, 32'h00000000} /* (0, 21, 30) {real, imag} */,
  {32'hc37cbe30, 32'h00000000} /* (0, 21, 29) {real, imag} */,
  {32'hc4c545d5, 32'h00000000} /* (0, 21, 28) {real, imag} */,
  {32'hc42e30b9, 32'h00000000} /* (0, 21, 27) {real, imag} */,
  {32'h429280b4, 32'h00000000} /* (0, 21, 26) {real, imag} */,
  {32'hc391ca28, 32'h00000000} /* (0, 21, 25) {real, imag} */,
  {32'hc3d6759a, 32'h00000000} /* (0, 21, 24) {real, imag} */,
  {32'h43a9f378, 32'h00000000} /* (0, 21, 23) {real, imag} */,
  {32'h43f2732c, 32'h00000000} /* (0, 21, 22) {real, imag} */,
  {32'h430f2078, 32'h00000000} /* (0, 21, 21) {real, imag} */,
  {32'h4345aba9, 32'h00000000} /* (0, 21, 20) {real, imag} */,
  {32'h4343bd84, 32'h00000000} /* (0, 21, 19) {real, imag} */,
  {32'h44272522, 32'h00000000} /* (0, 21, 18) {real, imag} */,
  {32'h43e05ec0, 32'h00000000} /* (0, 21, 17) {real, imag} */,
  {32'h430e6882, 32'h00000000} /* (0, 21, 16) {real, imag} */,
  {32'h43522876, 32'h00000000} /* (0, 21, 15) {real, imag} */,
  {32'h43d71b5a, 32'h00000000} /* (0, 21, 14) {real, imag} */,
  {32'h44b6a8d0, 32'h00000000} /* (0, 21, 13) {real, imag} */,
  {32'h445aa866, 32'h00000000} /* (0, 21, 12) {real, imag} */,
  {32'h447eeeaf, 32'h00000000} /* (0, 21, 11) {real, imag} */,
  {32'hc29807fc, 32'h00000000} /* (0, 21, 10) {real, imag} */,
  {32'hc38e504c, 32'h00000000} /* (0, 21, 9) {real, imag} */,
  {32'h441bfa15, 32'h00000000} /* (0, 21, 8) {real, imag} */,
  {32'hc3c1a9ba, 32'h00000000} /* (0, 21, 7) {real, imag} */,
  {32'hc397301c, 32'h00000000} /* (0, 21, 6) {real, imag} */,
  {32'hc12d5640, 32'h00000000} /* (0, 21, 5) {real, imag} */,
  {32'h430da5cf, 32'h00000000} /* (0, 21, 4) {real, imag} */,
  {32'hc23cd960, 32'h00000000} /* (0, 21, 3) {real, imag} */,
  {32'hc2caf84c, 32'h00000000} /* (0, 21, 2) {real, imag} */,
  {32'hc4249ef4, 32'h00000000} /* (0, 21, 1) {real, imag} */,
  {32'hc40e2d22, 32'h00000000} /* (0, 21, 0) {real, imag} */,
  {32'hbff3f600, 32'h00000000} /* (0, 20, 31) {real, imag} */,
  {32'h43145868, 32'h00000000} /* (0, 20, 30) {real, imag} */,
  {32'h4404ccfa, 32'h00000000} /* (0, 20, 29) {real, imag} */,
  {32'h4326a834, 32'h00000000} /* (0, 20, 28) {real, imag} */,
  {32'h43ec5ba7, 32'h00000000} /* (0, 20, 27) {real, imag} */,
  {32'h440f0d3f, 32'h00000000} /* (0, 20, 26) {real, imag} */,
  {32'h44bb98a0, 32'h00000000} /* (0, 20, 25) {real, imag} */,
  {32'h44cabb44, 32'h00000000} /* (0, 20, 24) {real, imag} */,
  {32'h4481ce0c, 32'h00000000} /* (0, 20, 23) {real, imag} */,
  {32'h4433c368, 32'h00000000} /* (0, 20, 22) {real, imag} */,
  {32'h4440a2a4, 32'h00000000} /* (0, 20, 21) {real, imag} */,
  {32'hc3d1a984, 32'h00000000} /* (0, 20, 20) {real, imag} */,
  {32'hc4269a4e, 32'h00000000} /* (0, 20, 19) {real, imag} */,
  {32'h42e678c2, 32'h00000000} /* (0, 20, 18) {real, imag} */,
  {32'hc3a36526, 32'h00000000} /* (0, 20, 17) {real, imag} */,
  {32'h439be89f, 32'h00000000} /* (0, 20, 16) {real, imag} */,
  {32'hc42784d6, 32'h00000000} /* (0, 20, 15) {real, imag} */,
  {32'hc399938e, 32'h00000000} /* (0, 20, 14) {real, imag} */,
  {32'hc3046bc9, 32'h00000000} /* (0, 20, 13) {real, imag} */,
  {32'h43cfd4da, 32'h00000000} /* (0, 20, 12) {real, imag} */,
  {32'h4401976a, 32'h00000000} /* (0, 20, 11) {real, imag} */,
  {32'hc3c451e2, 32'h00000000} /* (0, 20, 10) {real, imag} */,
  {32'h438533de, 32'h00000000} /* (0, 20, 9) {real, imag} */,
  {32'h4412e6eb, 32'h00000000} /* (0, 20, 8) {real, imag} */,
  {32'h43de7251, 32'h00000000} /* (0, 20, 7) {real, imag} */,
  {32'h44547e20, 32'h00000000} /* (0, 20, 6) {real, imag} */,
  {32'h43e4b3bc, 32'h00000000} /* (0, 20, 5) {real, imag} */,
  {32'h44264f1e, 32'h00000000} /* (0, 20, 4) {real, imag} */,
  {32'h43fe641c, 32'h00000000} /* (0, 20, 3) {real, imag} */,
  {32'h438ec48e, 32'h00000000} /* (0, 20, 2) {real, imag} */,
  {32'hc304776f, 32'h00000000} /* (0, 20, 1) {real, imag} */,
  {32'hc2e45fe4, 32'h00000000} /* (0, 20, 0) {real, imag} */,
  {32'h43ada329, 32'h00000000} /* (0, 19, 31) {real, imag} */,
  {32'h44bff794, 32'h00000000} /* (0, 19, 30) {real, imag} */,
  {32'h4487ca6c, 32'h00000000} /* (0, 19, 29) {real, imag} */,
  {32'h441d907c, 32'h00000000} /* (0, 19, 28) {real, imag} */,
  {32'h4489ca3a, 32'h00000000} /* (0, 19, 27) {real, imag} */,
  {32'h44973a87, 32'h00000000} /* (0, 19, 26) {real, imag} */,
  {32'h44c89ded, 32'h00000000} /* (0, 19, 25) {real, imag} */,
  {32'h44a67e7b, 32'h00000000} /* (0, 19, 24) {real, imag} */,
  {32'h444d2f8e, 32'h00000000} /* (0, 19, 23) {real, imag} */,
  {32'h4425b66a, 32'h00000000} /* (0, 19, 22) {real, imag} */,
  {32'h44302744, 32'h00000000} /* (0, 19, 21) {real, imag} */,
  {32'h4387b408, 32'h00000000} /* (0, 19, 20) {real, imag} */,
  {32'hc3573246, 32'h00000000} /* (0, 19, 19) {real, imag} */,
  {32'hc3ddae52, 32'h00000000} /* (0, 19, 18) {real, imag} */,
  {32'hc3f8e016, 32'h00000000} /* (0, 19, 17) {real, imag} */,
  {32'hc3c67dab, 32'h00000000} /* (0, 19, 16) {real, imag} */,
  {32'hc3b12317, 32'h00000000} /* (0, 19, 15) {real, imag} */,
  {32'hc3c596c8, 32'h00000000} /* (0, 19, 14) {real, imag} */,
  {32'h435e6584, 32'h00000000} /* (0, 19, 13) {real, imag} */,
  {32'h42ac7550, 32'h00000000} /* (0, 19, 12) {real, imag} */,
  {32'hc42e7dbc, 32'h00000000} /* (0, 19, 11) {real, imag} */,
  {32'h42808790, 32'h00000000} /* (0, 19, 10) {real, imag} */,
  {32'h444c67be, 32'h00000000} /* (0, 19, 9) {real, imag} */,
  {32'h43f29c1c, 32'h00000000} /* (0, 19, 8) {real, imag} */,
  {32'h448acd57, 32'h00000000} /* (0, 19, 7) {real, imag} */,
  {32'h4432cbb6, 32'h00000000} /* (0, 19, 6) {real, imag} */,
  {32'h4451430a, 32'h00000000} /* (0, 19, 5) {real, imag} */,
  {32'h44b55e55, 32'h00000000} /* (0, 19, 4) {real, imag} */,
  {32'h442d54e8, 32'h00000000} /* (0, 19, 3) {real, imag} */,
  {32'h43baa6d2, 32'h00000000} /* (0, 19, 2) {real, imag} */,
  {32'h441bac8b, 32'h00000000} /* (0, 19, 1) {real, imag} */,
  {32'h437c572a, 32'h00000000} /* (0, 19, 0) {real, imag} */,
  {32'h44207978, 32'h00000000} /* (0, 18, 31) {real, imag} */,
  {32'h4481df48, 32'h00000000} /* (0, 18, 30) {real, imag} */,
  {32'h4485f72c, 32'h00000000} /* (0, 18, 29) {real, imag} */,
  {32'h44232e1f, 32'h00000000} /* (0, 18, 28) {real, imag} */,
  {32'h445c02ee, 32'h00000000} /* (0, 18, 27) {real, imag} */,
  {32'h44c46261, 32'h00000000} /* (0, 18, 26) {real, imag} */,
  {32'h44991d68, 32'h00000000} /* (0, 18, 25) {real, imag} */,
  {32'h4500098f, 32'h00000000} /* (0, 18, 24) {real, imag} */,
  {32'h44b1cb0d, 32'h00000000} /* (0, 18, 23) {real, imag} */,
  {32'h44274442, 32'h00000000} /* (0, 18, 22) {real, imag} */,
  {32'h442900c4, 32'h00000000} /* (0, 18, 21) {real, imag} */,
  {32'h419ac550, 32'h00000000} /* (0, 18, 20) {real, imag} */,
  {32'hc3cb568c, 32'h00000000} /* (0, 18, 19) {real, imag} */,
  {32'hc475aaca, 32'h00000000} /* (0, 18, 18) {real, imag} */,
  {32'hc485bb26, 32'h00000000} /* (0, 18, 17) {real, imag} */,
  {32'hc39245f0, 32'h00000000} /* (0, 18, 16) {real, imag} */,
  {32'hc38dab25, 32'h00000000} /* (0, 18, 15) {real, imag} */,
  {32'hc40ad2ef, 32'h00000000} /* (0, 18, 14) {real, imag} */,
  {32'hc4a1105a, 32'h00000000} /* (0, 18, 13) {real, imag} */,
  {32'hc49f9102, 32'h00000000} /* (0, 18, 12) {real, imag} */,
  {32'hc42e7852, 32'h00000000} /* (0, 18, 11) {real, imag} */,
  {32'h4301c7f8, 32'h00000000} /* (0, 18, 10) {real, imag} */,
  {32'h42443f00, 32'h00000000} /* (0, 18, 9) {real, imag} */,
  {32'h441c67fd, 32'h00000000} /* (0, 18, 8) {real, imag} */,
  {32'h448be55f, 32'h00000000} /* (0, 18, 7) {real, imag} */,
  {32'h449b0dc5, 32'h00000000} /* (0, 18, 6) {real, imag} */,
  {32'h44ab6e69, 32'h00000000} /* (0, 18, 5) {real, imag} */,
  {32'h4471b52e, 32'h00000000} /* (0, 18, 4) {real, imag} */,
  {32'h4473dae8, 32'h00000000} /* (0, 18, 3) {real, imag} */,
  {32'h4446d7c6, 32'h00000000} /* (0, 18, 2) {real, imag} */,
  {32'h446d9e54, 32'h00000000} /* (0, 18, 1) {real, imag} */,
  {32'h41caa440, 32'h00000000} /* (0, 18, 0) {real, imag} */,
  {32'h4425ffd3, 32'h00000000} /* (0, 17, 31) {real, imag} */,
  {32'h4448ab2f, 32'h00000000} /* (0, 17, 30) {real, imag} */,
  {32'h44599c50, 32'h00000000} /* (0, 17, 29) {real, imag} */,
  {32'h44d226ae, 32'h00000000} /* (0, 17, 28) {real, imag} */,
  {32'h44a8997e, 32'h00000000} /* (0, 17, 27) {real, imag} */,
  {32'h44ccf7b0, 32'h00000000} /* (0, 17, 26) {real, imag} */,
  {32'h44ce8030, 32'h00000000} /* (0, 17, 25) {real, imag} */,
  {32'h44cfa580, 32'h00000000} /* (0, 17, 24) {real, imag} */,
  {32'h4478f102, 32'h00000000} /* (0, 17, 23) {real, imag} */,
  {32'h4482e6bb, 32'h00000000} /* (0, 17, 22) {real, imag} */,
  {32'h441f0dec, 32'h00000000} /* (0, 17, 21) {real, imag} */,
  {32'hc2a0480a, 32'h00000000} /* (0, 17, 20) {real, imag} */,
  {32'hbfc07600, 32'h00000000} /* (0, 17, 19) {real, imag} */,
  {32'hc4845123, 32'h00000000} /* (0, 17, 18) {real, imag} */,
  {32'hc4b51b8b, 32'h00000000} /* (0, 17, 17) {real, imag} */,
  {32'hc40da9d9, 32'h00000000} /* (0, 17, 16) {real, imag} */,
  {32'hc4823788, 32'h00000000} /* (0, 17, 15) {real, imag} */,
  {32'hc44158b9, 32'h00000000} /* (0, 17, 14) {real, imag} */,
  {32'hc42a7cc0, 32'h00000000} /* (0, 17, 13) {real, imag} */,
  {32'hc46c899d, 32'h00000000} /* (0, 17, 12) {real, imag} */,
  {32'hc406d12c, 32'h00000000} /* (0, 17, 11) {real, imag} */,
  {32'h4439e2e0, 32'h00000000} /* (0, 17, 10) {real, imag} */,
  {32'h442af347, 32'h00000000} /* (0, 17, 9) {real, imag} */,
  {32'h44113780, 32'h00000000} /* (0, 17, 8) {real, imag} */,
  {32'h44887353, 32'h00000000} /* (0, 17, 7) {real, imag} */,
  {32'h448410ad, 32'h00000000} /* (0, 17, 6) {real, imag} */,
  {32'h442268e8, 32'h00000000} /* (0, 17, 5) {real, imag} */,
  {32'h440eb50e, 32'h00000000} /* (0, 17, 4) {real, imag} */,
  {32'h43e660e4, 32'h00000000} /* (0, 17, 3) {real, imag} */,
  {32'h43a93a2d, 32'h00000000} /* (0, 17, 2) {real, imag} */,
  {32'h442bc9ee, 32'h00000000} /* (0, 17, 1) {real, imag} */,
  {32'h441b1bb1, 32'h00000000} /* (0, 17, 0) {real, imag} */,
  {32'h43b84c52, 32'h00000000} /* (0, 16, 31) {real, imag} */,
  {32'h44a0a804, 32'h00000000} /* (0, 16, 30) {real, imag} */,
  {32'h44d475ff, 32'h00000000} /* (0, 16, 29) {real, imag} */,
  {32'h44e55fae, 32'h00000000} /* (0, 16, 28) {real, imag} */,
  {32'h4505b6cc, 32'h00000000} /* (0, 16, 27) {real, imag} */,
  {32'h44b3e490, 32'h00000000} /* (0, 16, 26) {real, imag} */,
  {32'h44d98b20, 32'h00000000} /* (0, 16, 25) {real, imag} */,
  {32'h44a0f1bc, 32'h00000000} /* (0, 16, 24) {real, imag} */,
  {32'h447a5fd2, 32'h00000000} /* (0, 16, 23) {real, imag} */,
  {32'h44bb9c56, 32'h00000000} /* (0, 16, 22) {real, imag} */,
  {32'h4402f8e6, 32'h00000000} /* (0, 16, 21) {real, imag} */,
  {32'h42d319ae, 32'h00000000} /* (0, 16, 20) {real, imag} */,
  {32'hc3aa41e3, 32'h00000000} /* (0, 16, 19) {real, imag} */,
  {32'hc2f07358, 32'h00000000} /* (0, 16, 18) {real, imag} */,
  {32'hc4a68a34, 32'h00000000} /* (0, 16, 17) {real, imag} */,
  {32'hc49ce7e8, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hc48fc186, 32'h00000000} /* (0, 16, 15) {real, imag} */,
  {32'hc48269cc, 32'h00000000} /* (0, 16, 14) {real, imag} */,
  {32'hc4c5f6e1, 32'h00000000} /* (0, 16, 13) {real, imag} */,
  {32'hc4bb0752, 32'h00000000} /* (0, 16, 12) {real, imag} */,
  {32'hc4025ec8, 32'h00000000} /* (0, 16, 11) {real, imag} */,
  {32'h43852128, 32'h00000000} /* (0, 16, 10) {real, imag} */,
  {32'h450ce082, 32'h00000000} /* (0, 16, 9) {real, imag} */,
  {32'h44da05be, 32'h00000000} /* (0, 16, 8) {real, imag} */,
  {32'h44afb47f, 32'h00000000} /* (0, 16, 7) {real, imag} */,
  {32'h44aff816, 32'h00000000} /* (0, 16, 6) {real, imag} */,
  {32'h44473bd6, 32'h00000000} /* (0, 16, 5) {real, imag} */,
  {32'h43f0310c, 32'h00000000} /* (0, 16, 4) {real, imag} */,
  {32'h4401346e, 32'h00000000} /* (0, 16, 3) {real, imag} */,
  {32'h43f02500, 32'h00000000} /* (0, 16, 2) {real, imag} */,
  {32'h442e1779, 32'h00000000} /* (0, 16, 1) {real, imag} */,
  {32'h444fe01c, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h448f92af, 32'h00000000} /* (0, 15, 31) {real, imag} */,
  {32'h448b7ca2, 32'h00000000} /* (0, 15, 30) {real, imag} */,
  {32'h44dc2735, 32'h00000000} /* (0, 15, 29) {real, imag} */,
  {32'h44c32c6e, 32'h00000000} /* (0, 15, 28) {real, imag} */,
  {32'h44c4b1ee, 32'h00000000} /* (0, 15, 27) {real, imag} */,
  {32'h44a6cf33, 32'h00000000} /* (0, 15, 26) {real, imag} */,
  {32'h4476e0c0, 32'h00000000} /* (0, 15, 25) {real, imag} */,
  {32'h4440e306, 32'h00000000} /* (0, 15, 24) {real, imag} */,
  {32'h44897c54, 32'h00000000} /* (0, 15, 23) {real, imag} */,
  {32'h4406e278, 32'h00000000} /* (0, 15, 22) {real, imag} */,
  {32'h43ca5100, 32'h00000000} /* (0, 15, 21) {real, imag} */,
  {32'h422cdd60, 32'h00000000} /* (0, 15, 20) {real, imag} */,
  {32'hc4050cee, 32'h00000000} /* (0, 15, 19) {real, imag} */,
  {32'hc4438938, 32'h00000000} /* (0, 15, 18) {real, imag} */,
  {32'hc4510511, 32'h00000000} /* (0, 15, 17) {real, imag} */,
  {32'hc463127d, 32'h00000000} /* (0, 15, 16) {real, imag} */,
  {32'hc4d53cf1, 32'h00000000} /* (0, 15, 15) {real, imag} */,
  {32'hc4d76dca, 32'h00000000} /* (0, 15, 14) {real, imag} */,
  {32'hc4ffb22d, 32'h00000000} /* (0, 15, 13) {real, imag} */,
  {32'hc533ef05, 32'h00000000} /* (0, 15, 12) {real, imag} */,
  {32'hc4c227d4, 32'h00000000} /* (0, 15, 11) {real, imag} */,
  {32'hc3c12cdf, 32'h00000000} /* (0, 15, 10) {real, imag} */,
  {32'h44337826, 32'h00000000} /* (0, 15, 9) {real, imag} */,
  {32'h434bdb20, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'h4423e6cc, 32'h00000000} /* (0, 15, 7) {real, imag} */,
  {32'h44c94840, 32'h00000000} /* (0, 15, 6) {real, imag} */,
  {32'h44a238d2, 32'h00000000} /* (0, 15, 5) {real, imag} */,
  {32'h44c436d9, 32'h00000000} /* (0, 15, 4) {real, imag} */,
  {32'h445f6f2e, 32'h00000000} /* (0, 15, 3) {real, imag} */,
  {32'h44d966fa, 32'h00000000} /* (0, 15, 2) {real, imag} */,
  {32'h44a5fe72, 32'h00000000} /* (0, 15, 1) {real, imag} */,
  {32'h43ed3ece, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h443beb52, 32'h00000000} /* (0, 14, 31) {real, imag} */,
  {32'h447b319e, 32'h00000000} /* (0, 14, 30) {real, imag} */,
  {32'h44a36bba, 32'h00000000} /* (0, 14, 29) {real, imag} */,
  {32'h44c29233, 32'h00000000} /* (0, 14, 28) {real, imag} */,
  {32'h44ad261c, 32'h00000000} /* (0, 14, 27) {real, imag} */,
  {32'h44bd7170, 32'h00000000} /* (0, 14, 26) {real, imag} */,
  {32'h448ab3a7, 32'h00000000} /* (0, 14, 25) {real, imag} */,
  {32'h443b7ab8, 32'h00000000} /* (0, 14, 24) {real, imag} */,
  {32'h44802618, 32'h00000000} /* (0, 14, 23) {real, imag} */,
  {32'h44149b15, 32'h00000000} /* (0, 14, 22) {real, imag} */,
  {32'h432a5168, 32'h00000000} /* (0, 14, 21) {real, imag} */,
  {32'hc43b435a, 32'h00000000} /* (0, 14, 20) {real, imag} */,
  {32'hc4624c26, 32'h00000000} /* (0, 14, 19) {real, imag} */,
  {32'hc49e510c, 32'h00000000} /* (0, 14, 18) {real, imag} */,
  {32'hc4f2871c, 32'h00000000} /* (0, 14, 17) {real, imag} */,
  {32'hc47f9ee8, 32'h00000000} /* (0, 14, 16) {real, imag} */,
  {32'hc48ff896, 32'h00000000} /* (0, 14, 15) {real, imag} */,
  {32'hc48ac3b5, 32'h00000000} /* (0, 14, 14) {real, imag} */,
  {32'hc494ea38, 32'h00000000} /* (0, 14, 13) {real, imag} */,
  {32'hc4b674e1, 32'h00000000} /* (0, 14, 12) {real, imag} */,
  {32'hc4736c00, 32'h00000000} /* (0, 14, 11) {real, imag} */,
  {32'hc3d559ea, 32'h00000000} /* (0, 14, 10) {real, imag} */,
  {32'hc3100b78, 32'h00000000} /* (0, 14, 9) {real, imag} */,
  {32'h43af9121, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'h44016dfe, 32'h00000000} /* (0, 14, 7) {real, imag} */,
  {32'h4416a73b, 32'h00000000} /* (0, 14, 6) {real, imag} */,
  {32'h44be973c, 32'h00000000} /* (0, 14, 5) {real, imag} */,
  {32'h44c1f441, 32'h00000000} /* (0, 14, 4) {real, imag} */,
  {32'h44bf8ca5, 32'h00000000} /* (0, 14, 3) {real, imag} */,
  {32'h44a856d8, 32'h00000000} /* (0, 14, 2) {real, imag} */,
  {32'h448d8faa, 32'h00000000} /* (0, 14, 1) {real, imag} */,
  {32'h4462937c, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h44244e88, 32'h00000000} /* (0, 13, 31) {real, imag} */,
  {32'h44888a68, 32'h00000000} /* (0, 13, 30) {real, imag} */,
  {32'h44bd743c, 32'h00000000} /* (0, 13, 29) {real, imag} */,
  {32'h44a0e401, 32'h00000000} /* (0, 13, 28) {real, imag} */,
  {32'h44b5ad39, 32'h00000000} /* (0, 13, 27) {real, imag} */,
  {32'h44ab2043, 32'h00000000} /* (0, 13, 26) {real, imag} */,
  {32'h44adeb02, 32'h00000000} /* (0, 13, 25) {real, imag} */,
  {32'h44512309, 32'h00000000} /* (0, 13, 24) {real, imag} */,
  {32'h44300d96, 32'h00000000} /* (0, 13, 23) {real, imag} */,
  {32'h448969c0, 32'h00000000} /* (0, 13, 22) {real, imag} */,
  {32'hc3b50e8b, 32'h00000000} /* (0, 13, 21) {real, imag} */,
  {32'hc4a59eee, 32'h00000000} /* (0, 13, 20) {real, imag} */,
  {32'hc49e0cfc, 32'h00000000} /* (0, 13, 19) {real, imag} */,
  {32'hc4db49f1, 32'h00000000} /* (0, 13, 18) {real, imag} */,
  {32'hc4c6918a, 32'h00000000} /* (0, 13, 17) {real, imag} */,
  {32'hc4b0ce66, 32'h00000000} /* (0, 13, 16) {real, imag} */,
  {32'hc480bf11, 32'h00000000} /* (0, 13, 15) {real, imag} */,
  {32'hc444bac0, 32'h00000000} /* (0, 13, 14) {real, imag} */,
  {32'hc48a18bc, 32'h00000000} /* (0, 13, 13) {real, imag} */,
  {32'hc49fcf9f, 32'h00000000} /* (0, 13, 12) {real, imag} */,
  {32'hc47f46ee, 32'h00000000} /* (0, 13, 11) {real, imag} */,
  {32'hc45b681e, 32'h00000000} /* (0, 13, 10) {real, imag} */,
  {32'h41c40340, 32'h00000000} /* (0, 13, 9) {real, imag} */,
  {32'h43ccdc26, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'h44b32e1d, 32'h00000000} /* (0, 13, 7) {real, imag} */,
  {32'h444e42b1, 32'h00000000} /* (0, 13, 6) {real, imag} */,
  {32'h4445bf32, 32'h00000000} /* (0, 13, 5) {real, imag} */,
  {32'h44658ba7, 32'h00000000} /* (0, 13, 4) {real, imag} */,
  {32'h44836d04, 32'h00000000} /* (0, 13, 3) {real, imag} */,
  {32'h448ec92d, 32'h00000000} /* (0, 13, 2) {real, imag} */,
  {32'h44aee210, 32'h00000000} /* (0, 13, 1) {real, imag} */,
  {32'h4445b578, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'h4446f2d0, 32'h00000000} /* (0, 12, 31) {real, imag} */,
  {32'h448f95db, 32'h00000000} /* (0, 12, 30) {real, imag} */,
  {32'h44186f19, 32'h00000000} /* (0, 12, 29) {real, imag} */,
  {32'h44aabeca, 32'h00000000} /* (0, 12, 28) {real, imag} */,
  {32'h44822eba, 32'h00000000} /* (0, 12, 27) {real, imag} */,
  {32'h447edc31, 32'h00000000} /* (0, 12, 26) {real, imag} */,
  {32'h448944b6, 32'h00000000} /* (0, 12, 25) {real, imag} */,
  {32'h444b7b00, 32'h00000000} /* (0, 12, 24) {real, imag} */,
  {32'h4424f0ee, 32'h00000000} /* (0, 12, 23) {real, imag} */,
  {32'h4424341e, 32'h00000000} /* (0, 12, 22) {real, imag} */,
  {32'h44146cca, 32'h00000000} /* (0, 12, 21) {real, imag} */,
  {32'hc3bdb4db, 32'h00000000} /* (0, 12, 20) {real, imag} */,
  {32'hc483c3be, 32'h00000000} /* (0, 12, 19) {real, imag} */,
  {32'hc4845b30, 32'h00000000} /* (0, 12, 18) {real, imag} */,
  {32'hc46257a4, 32'h00000000} /* (0, 12, 17) {real, imag} */,
  {32'hc4dabdbb, 32'h00000000} /* (0, 12, 16) {real, imag} */,
  {32'hc41696c6, 32'h00000000} /* (0, 12, 15) {real, imag} */,
  {32'hc4822c09, 32'h00000000} /* (0, 12, 14) {real, imag} */,
  {32'hc4822b36, 32'h00000000} /* (0, 12, 13) {real, imag} */,
  {32'hc44f72cc, 32'h00000000} /* (0, 12, 12) {real, imag} */,
  {32'hc4528f69, 32'h00000000} /* (0, 12, 11) {real, imag} */,
  {32'hc3f72b6a, 32'h00000000} /* (0, 12, 10) {real, imag} */,
  {32'hc38ab7b6, 32'h00000000} /* (0, 12, 9) {real, imag} */,
  {32'h43e608ef, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'h44971dad, 32'h00000000} /* (0, 12, 7) {real, imag} */,
  {32'h446a647e, 32'h00000000} /* (0, 12, 6) {real, imag} */,
  {32'h448c8365, 32'h00000000} /* (0, 12, 5) {real, imag} */,
  {32'h447d92a2, 32'h00000000} /* (0, 12, 4) {real, imag} */,
  {32'h43c360f6, 32'h00000000} /* (0, 12, 3) {real, imag} */,
  {32'h4442b2bd, 32'h00000000} /* (0, 12, 2) {real, imag} */,
  {32'h44a8a066, 32'h00000000} /* (0, 12, 1) {real, imag} */,
  {32'h440bf576, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h43d654e1, 32'h00000000} /* (0, 11, 31) {real, imag} */,
  {32'h441bd21c, 32'h00000000} /* (0, 11, 30) {real, imag} */,
  {32'h443c81f8, 32'h00000000} /* (0, 11, 29) {real, imag} */,
  {32'h441ec5ee, 32'h00000000} /* (0, 11, 28) {real, imag} */,
  {32'h44228034, 32'h00000000} /* (0, 11, 27) {real, imag} */,
  {32'hc1855ed8, 32'h00000000} /* (0, 11, 26) {real, imag} */,
  {32'h43ffd667, 32'h00000000} /* (0, 11, 25) {real, imag} */,
  {32'h4471d495, 32'h00000000} /* (0, 11, 24) {real, imag} */,
  {32'h42a172e4, 32'h00000000} /* (0, 11, 23) {real, imag} */,
  {32'h441fdf8a, 32'h00000000} /* (0, 11, 22) {real, imag} */,
  {32'h44333d86, 32'h00000000} /* (0, 11, 21) {real, imag} */,
  {32'hc4309d9b, 32'h00000000} /* (0, 11, 20) {real, imag} */,
  {32'hc4046f22, 32'h00000000} /* (0, 11, 19) {real, imag} */,
  {32'hc4389c80, 32'h00000000} /* (0, 11, 18) {real, imag} */,
  {32'hc4f54306, 32'h00000000} /* (0, 11, 17) {real, imag} */,
  {32'hc4804234, 32'h00000000} /* (0, 11, 16) {real, imag} */,
  {32'hc42c6b5a, 32'h00000000} /* (0, 11, 15) {real, imag} */,
  {32'hc4938643, 32'h00000000} /* (0, 11, 14) {real, imag} */,
  {32'hc4538f0c, 32'h00000000} /* (0, 11, 13) {real, imag} */,
  {32'hc42950a8, 32'h00000000} /* (0, 11, 12) {real, imag} */,
  {32'hc43f45a0, 32'h00000000} /* (0, 11, 11) {real, imag} */,
  {32'hc3dda666, 32'h00000000} /* (0, 11, 10) {real, imag} */,
  {32'hc29fd124, 32'h00000000} /* (0, 11, 9) {real, imag} */,
  {32'h4387d8b6, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'h4466f90c, 32'h00000000} /* (0, 11, 7) {real, imag} */,
  {32'h442959d6, 32'h00000000} /* (0, 11, 6) {real, imag} */,
  {32'h44ab4923, 32'h00000000} /* (0, 11, 5) {real, imag} */,
  {32'h4426b06b, 32'h00000000} /* (0, 11, 4) {real, imag} */,
  {32'h43569b01, 32'h00000000} /* (0, 11, 3) {real, imag} */,
  {32'h43a3b760, 32'h00000000} /* (0, 11, 2) {real, imag} */,
  {32'h4369b500, 32'h00000000} /* (0, 11, 1) {real, imag} */,
  {32'h437c4fe6, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h42960cec, 32'h00000000} /* (0, 10, 31) {real, imag} */,
  {32'hc40b919a, 32'h00000000} /* (0, 10, 30) {real, imag} */,
  {32'h43b3fb32, 32'h00000000} /* (0, 10, 29) {real, imag} */,
  {32'hc1770d50, 32'h00000000} /* (0, 10, 28) {real, imag} */,
  {32'hc48b335a, 32'h00000000} /* (0, 10, 27) {real, imag} */,
  {32'hc418255a, 32'h00000000} /* (0, 10, 26) {real, imag} */,
  {32'hc3ba6947, 32'h00000000} /* (0, 10, 25) {real, imag} */,
  {32'hc323fe17, 32'h00000000} /* (0, 10, 24) {real, imag} */,
  {32'hc4836341, 32'h00000000} /* (0, 10, 23) {real, imag} */,
  {32'hc4181d72, 32'h00000000} /* (0, 10, 22) {real, imag} */,
  {32'hc4a4e026, 32'h00000000} /* (0, 10, 21) {real, imag} */,
  {32'h44019e40, 32'h00000000} /* (0, 10, 20) {real, imag} */,
  {32'h43c7bc62, 32'h00000000} /* (0, 10, 19) {real, imag} */,
  {32'hc3d9786d, 32'h00000000} /* (0, 10, 18) {real, imag} */,
  {32'hc21190ce, 32'h00000000} /* (0, 10, 17) {real, imag} */,
  {32'hc2997686, 32'h00000000} /* (0, 10, 16) {real, imag} */,
  {32'hc3d958dd, 32'h00000000} /* (0, 10, 15) {real, imag} */,
  {32'hc3db6ca9, 32'h00000000} /* (0, 10, 14) {real, imag} */,
  {32'hc3eb131a, 32'h00000000} /* (0, 10, 13) {real, imag} */,
  {32'hc3e0797c, 32'h00000000} /* (0, 10, 12) {real, imag} */,
  {32'hc417b41e, 32'h00000000} /* (0, 10, 11) {real, imag} */,
  {32'hc411afa8, 32'h00000000} /* (0, 10, 10) {real, imag} */,
  {32'hc46edf56, 32'h00000000} /* (0, 10, 9) {real, imag} */,
  {32'hc3a7eb5c, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'hc3b3da3c, 32'h00000000} /* (0, 10, 7) {real, imag} */,
  {32'h43f9cda0, 32'h00000000} /* (0, 10, 6) {real, imag} */,
  {32'hc3a3ed88, 32'h00000000} /* (0, 10, 5) {real, imag} */,
  {32'h43d08725, 32'h00000000} /* (0, 10, 4) {real, imag} */,
  {32'h42d24a48, 32'h00000000} /* (0, 10, 3) {real, imag} */,
  {32'hc40d65fd, 32'h00000000} /* (0, 10, 2) {real, imag} */,
  {32'hc37371d4, 32'h00000000} /* (0, 10, 1) {real, imag} */,
  {32'h431f2044, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'hc397a8e4, 32'h00000000} /* (0, 9, 31) {real, imag} */,
  {32'hc426728a, 32'h00000000} /* (0, 9, 30) {real, imag} */,
  {32'hc407fa31, 32'h00000000} /* (0, 9, 29) {real, imag} */,
  {32'hc46637af, 32'h00000000} /* (0, 9, 28) {real, imag} */,
  {32'hc4813db6, 32'h00000000} /* (0, 9, 27) {real, imag} */,
  {32'hc46c8d37, 32'h00000000} /* (0, 9, 26) {real, imag} */,
  {32'hc4407adc, 32'h00000000} /* (0, 9, 25) {real, imag} */,
  {32'hc433ebd5, 32'h00000000} /* (0, 9, 24) {real, imag} */,
  {32'hc417d487, 32'h00000000} /* (0, 9, 23) {real, imag} */,
  {32'hc4c5ae1a, 32'h00000000} /* (0, 9, 22) {real, imag} */,
  {32'hc42a9c67, 32'h00000000} /* (0, 9, 21) {real, imag} */,
  {32'hc388b260, 32'h00000000} /* (0, 9, 20) {real, imag} */,
  {32'h42264596, 32'h00000000} /* (0, 9, 19) {real, imag} */,
  {32'h43d39a7f, 32'h00000000} /* (0, 9, 18) {real, imag} */,
  {32'h438b258b, 32'h00000000} /* (0, 9, 17) {real, imag} */,
  {32'h4381ed28, 32'h00000000} /* (0, 9, 16) {real, imag} */,
  {32'hc38afd5c, 32'h00000000} /* (0, 9, 15) {real, imag} */,
  {32'h4389b38f, 32'h00000000} /* (0, 9, 14) {real, imag} */,
  {32'hc316273c, 32'h00000000} /* (0, 9, 13) {real, imag} */,
  {32'h442e7a71, 32'h00000000} /* (0, 9, 12) {real, imag} */,
  {32'h444c3cf0, 32'h00000000} /* (0, 9, 11) {real, imag} */,
  {32'hc4091c07, 32'h00000000} /* (0, 9, 10) {real, imag} */,
  {32'hc3e4111f, 32'h00000000} /* (0, 9, 9) {real, imag} */,
  {32'hc3d90f82, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'hc44294b1, 32'h00000000} /* (0, 9, 7) {real, imag} */,
  {32'hc31555dc, 32'h00000000} /* (0, 9, 6) {real, imag} */,
  {32'hc3db5632, 32'h00000000} /* (0, 9, 5) {real, imag} */,
  {32'hc3e75bb6, 32'h00000000} /* (0, 9, 4) {real, imag} */,
  {32'hc3120946, 32'h00000000} /* (0, 9, 3) {real, imag} */,
  {32'hc3a762a7, 32'h00000000} /* (0, 9, 2) {real, imag} */,
  {32'hc4527f9e, 32'h00000000} /* (0, 9, 1) {real, imag} */,
  {32'hc3cb628c, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'hc3b87906, 32'h00000000} /* (0, 8, 31) {real, imag} */,
  {32'hc3ad64d8, 32'h00000000} /* (0, 8, 30) {real, imag} */,
  {32'hc45ded70, 32'h00000000} /* (0, 8, 29) {real, imag} */,
  {32'hc493705a, 32'h00000000} /* (0, 8, 28) {real, imag} */,
  {32'hc473678e, 32'h00000000} /* (0, 8, 27) {real, imag} */,
  {32'hc4ba307e, 32'h00000000} /* (0, 8, 26) {real, imag} */,
  {32'hc49852ea, 32'h00000000} /* (0, 8, 25) {real, imag} */,
  {32'hc4a6c207, 32'h00000000} /* (0, 8, 24) {real, imag} */,
  {32'hc4a154c6, 32'h00000000} /* (0, 8, 23) {real, imag} */,
  {32'hc4aa697c, 32'h00000000} /* (0, 8, 22) {real, imag} */,
  {32'hc3f2585a, 32'h00000000} /* (0, 8, 21) {real, imag} */,
  {32'h431dccf2, 32'h00000000} /* (0, 8, 20) {real, imag} */,
  {32'h439a3b91, 32'h00000000} /* (0, 8, 19) {real, imag} */,
  {32'h43cedca1, 32'h00000000} /* (0, 8, 18) {real, imag} */,
  {32'h43987636, 32'h00000000} /* (0, 8, 17) {real, imag} */,
  {32'h4407062c, 32'h00000000} /* (0, 8, 16) {real, imag} */,
  {32'h4483fa58, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'h442354ac, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'h43bc7bd9, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'h44123093, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'h42b325ec, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'hc301bf20, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hc400395e, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'hc30e42d8, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hc35cde3c, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hc3b72c5a, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'hc370a390, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'hc398774a, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'hc40a0464, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'hc4513592, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'hc470ab55, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'hc4336910, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'hc45f5106, 32'h00000000} /* (0, 7, 31) {real, imag} */,
  {32'hc47430c4, 32'h00000000} /* (0, 7, 30) {real, imag} */,
  {32'hc47a051c, 32'h00000000} /* (0, 7, 29) {real, imag} */,
  {32'hc4b85ace, 32'h00000000} /* (0, 7, 28) {real, imag} */,
  {32'hc4afe19e, 32'h00000000} /* (0, 7, 27) {real, imag} */,
  {32'hc4cfd6c3, 32'h00000000} /* (0, 7, 26) {real, imag} */,
  {32'hc4c7f91a, 32'h00000000} /* (0, 7, 25) {real, imag} */,
  {32'hc4b02c66, 32'h00000000} /* (0, 7, 24) {real, imag} */,
  {32'hc4c57f3f, 32'h00000000} /* (0, 7, 23) {real, imag} */,
  {32'hc40949e5, 32'h00000000} /* (0, 7, 22) {real, imag} */,
  {32'hc3a8a6be, 32'h00000000} /* (0, 7, 21) {real, imag} */,
  {32'h43a85e16, 32'h00000000} /* (0, 7, 20) {real, imag} */,
  {32'h44321500, 32'h00000000} /* (0, 7, 19) {real, imag} */,
  {32'h436709f0, 32'h00000000} /* (0, 7, 18) {real, imag} */,
  {32'h43acb5f1, 32'h00000000} /* (0, 7, 17) {real, imag} */,
  {32'h43d1d305, 32'h00000000} /* (0, 7, 16) {real, imag} */,
  {32'h445bda4a, 32'h00000000} /* (0, 7, 15) {real, imag} */,
  {32'h44c86a96, 32'h00000000} /* (0, 7, 14) {real, imag} */,
  {32'h44476b36, 32'h00000000} /* (0, 7, 13) {real, imag} */,
  {32'h4420a495, 32'h00000000} /* (0, 7, 12) {real, imag} */,
  {32'hc271a8f0, 32'h00000000} /* (0, 7, 11) {real, imag} */,
  {32'hc4848ab9, 32'h00000000} /* (0, 7, 10) {real, imag} */,
  {32'hc3bf6a28, 32'h00000000} /* (0, 7, 9) {real, imag} */,
  {32'hc318ad94, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'hc3ab537c, 32'h00000000} /* (0, 7, 7) {real, imag} */,
  {32'hc4600abb, 32'h00000000} /* (0, 7, 6) {real, imag} */,
  {32'hc4550d3d, 32'h00000000} /* (0, 7, 5) {real, imag} */,
  {32'hc3f60be8, 32'h00000000} /* (0, 7, 4) {real, imag} */,
  {32'hc40acba8, 32'h00000000} /* (0, 7, 3) {real, imag} */,
  {32'hc4a177d2, 32'h00000000} /* (0, 7, 2) {real, imag} */,
  {32'hc4a7b884, 32'h00000000} /* (0, 7, 1) {real, imag} */,
  {32'hc38d2371, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'hc455fba6, 32'h00000000} /* (0, 6, 31) {real, imag} */,
  {32'hc4370190, 32'h00000000} /* (0, 6, 30) {real, imag} */,
  {32'hc4a048e2, 32'h00000000} /* (0, 6, 29) {real, imag} */,
  {32'hc4ffc31a, 32'h00000000} /* (0, 6, 28) {real, imag} */,
  {32'hc4d4ea65, 32'h00000000} /* (0, 6, 27) {real, imag} */,
  {32'hc5082070, 32'h00000000} /* (0, 6, 26) {real, imag} */,
  {32'hc4ed220f, 32'h00000000} /* (0, 6, 25) {real, imag} */,
  {32'hc512792e, 32'h00000000} /* (0, 6, 24) {real, imag} */,
  {32'hc484b6c4, 32'h00000000} /* (0, 6, 23) {real, imag} */,
  {32'hc4cb6e63, 32'h00000000} /* (0, 6, 22) {real, imag} */,
  {32'hc414c418, 32'h00000000} /* (0, 6, 21) {real, imag} */,
  {32'h44862c60, 32'h00000000} /* (0, 6, 20) {real, imag} */,
  {32'h43bbf3e4, 32'h00000000} /* (0, 6, 19) {real, imag} */,
  {32'h43ea6168, 32'h00000000} /* (0, 6, 18) {real, imag} */,
  {32'h441dc7e4, 32'h00000000} /* (0, 6, 17) {real, imag} */,
  {32'h430c9f28, 32'h00000000} /* (0, 6, 16) {real, imag} */,
  {32'h441cff24, 32'h00000000} /* (0, 6, 15) {real, imag} */,
  {32'h449d0dea, 32'h00000000} /* (0, 6, 14) {real, imag} */,
  {32'h43970a9a, 32'h00000000} /* (0, 6, 13) {real, imag} */,
  {32'h43e55f68, 32'h00000000} /* (0, 6, 12) {real, imag} */,
  {32'h439bff9c, 32'h00000000} /* (0, 6, 11) {real, imag} */,
  {32'hc38ed88c, 32'h00000000} /* (0, 6, 10) {real, imag} */,
  {32'hc473d8ca, 32'h00000000} /* (0, 6, 9) {real, imag} */,
  {32'hc45fbfc3, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'hc3ba95c5, 32'h00000000} /* (0, 6, 7) {real, imag} */,
  {32'hc44e1d5e, 32'h00000000} /* (0, 6, 6) {real, imag} */,
  {32'hc44b8a04, 32'h00000000} /* (0, 6, 5) {real, imag} */,
  {32'hc4157fa0, 32'h00000000} /* (0, 6, 4) {real, imag} */,
  {32'hc3aa0b5e, 32'h00000000} /* (0, 6, 3) {real, imag} */,
  {32'hc42b5dd4, 32'h00000000} /* (0, 6, 2) {real, imag} */,
  {32'hc3af5274, 32'h00000000} /* (0, 6, 1) {real, imag} */,
  {32'hc3f3d78c, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hc4ad85cb, 32'h00000000} /* (0, 5, 31) {real, imag} */,
  {32'hc4d69c4c, 32'h00000000} /* (0, 5, 30) {real, imag} */,
  {32'hc4e86475, 32'h00000000} /* (0, 5, 29) {real, imag} */,
  {32'hc529ec26, 32'h00000000} /* (0, 5, 28) {real, imag} */,
  {32'hc5331266, 32'h00000000} /* (0, 5, 27) {real, imag} */,
  {32'hc4d148c0, 32'h00000000} /* (0, 5, 26) {real, imag} */,
  {32'hc4ea4b4a, 32'h00000000} /* (0, 5, 25) {real, imag} */,
  {32'hc50494e2, 32'h00000000} /* (0, 5, 24) {real, imag} */,
  {32'hc4ff30ae, 32'h00000000} /* (0, 5, 23) {real, imag} */,
  {32'hc4a09444, 32'h00000000} /* (0, 5, 22) {real, imag} */,
  {32'hc445504e, 32'h00000000} /* (0, 5, 21) {real, imag} */,
  {32'hc44744ee, 32'h00000000} /* (0, 5, 20) {real, imag} */,
  {32'hc3849ea7, 32'h00000000} /* (0, 5, 19) {real, imag} */,
  {32'hc3a35ab0, 32'h00000000} /* (0, 5, 18) {real, imag} */,
  {32'hc498d107, 32'h00000000} /* (0, 5, 17) {real, imag} */,
  {32'hc417b03d, 32'h00000000} /* (0, 5, 16) {real, imag} */,
  {32'hc3b3655c, 32'h00000000} /* (0, 5, 15) {real, imag} */,
  {32'h43f1a9e8, 32'h00000000} /* (0, 5, 14) {real, imag} */,
  {32'h438fadac, 32'h00000000} /* (0, 5, 13) {real, imag} */,
  {32'h436b3600, 32'h00000000} /* (0, 5, 12) {real, imag} */,
  {32'h42d9b9f0, 32'h00000000} /* (0, 5, 11) {real, imag} */,
  {32'h434e3b30, 32'h00000000} /* (0, 5, 10) {real, imag} */,
  {32'h409ce180, 32'h00000000} /* (0, 5, 9) {real, imag} */,
  {32'h43d7ad04, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'hc2adcf88, 32'h00000000} /* (0, 5, 7) {real, imag} */,
  {32'hc426f289, 32'h00000000} /* (0, 5, 6) {real, imag} */,
  {32'hc28f2dc8, 32'h00000000} /* (0, 5, 5) {real, imag} */,
  {32'hc3e81f48, 32'h00000000} /* (0, 5, 4) {real, imag} */,
  {32'hc438a53a, 32'h00000000} /* (0, 5, 3) {real, imag} */,
  {32'hc4399770, 32'h00000000} /* (0, 5, 2) {real, imag} */,
  {32'hc49d2e67, 32'h00000000} /* (0, 5, 1) {real, imag} */,
  {32'hc416e823, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hc4c0c9fc, 32'h00000000} /* (0, 4, 31) {real, imag} */,
  {32'hc4d5969a, 32'h00000000} /* (0, 4, 30) {real, imag} */,
  {32'hc4eb1e4e, 32'h00000000} /* (0, 4, 29) {real, imag} */,
  {32'hc53bb586, 32'h00000000} /* (0, 4, 28) {real, imag} */,
  {32'hc4ffa3b3, 32'h00000000} /* (0, 4, 27) {real, imag} */,
  {32'hc4f9b5ac, 32'h00000000} /* (0, 4, 26) {real, imag} */,
  {32'hc4bc2ff2, 32'h00000000} /* (0, 4, 25) {real, imag} */,
  {32'hc4f87529, 32'h00000000} /* (0, 4, 24) {real, imag} */,
  {32'hc4bdc201, 32'h00000000} /* (0, 4, 23) {real, imag} */,
  {32'hc4acc367, 32'h00000000} /* (0, 4, 22) {real, imag} */,
  {32'hc433d83c, 32'h00000000} /* (0, 4, 21) {real, imag} */,
  {32'hc46ff544, 32'h00000000} /* (0, 4, 20) {real, imag} */,
  {32'hc4da1565, 32'h00000000} /* (0, 4, 19) {real, imag} */,
  {32'hc4391788, 32'h00000000} /* (0, 4, 18) {real, imag} */,
  {32'hc498f03f, 32'h00000000} /* (0, 4, 17) {real, imag} */,
  {32'hc4a06d57, 32'h00000000} /* (0, 4, 16) {real, imag} */,
  {32'h43c5a2c0, 32'h00000000} /* (0, 4, 15) {real, imag} */,
  {32'h449c9ed6, 32'h00000000} /* (0, 4, 14) {real, imag} */,
  {32'h44018344, 32'h00000000} /* (0, 4, 13) {real, imag} */,
  {32'h43a27f34, 32'h00000000} /* (0, 4, 12) {real, imag} */,
  {32'h443c342a, 32'h00000000} /* (0, 4, 11) {real, imag} */,
  {32'h44024c19, 32'h00000000} /* (0, 4, 10) {real, imag} */,
  {32'h44872796, 32'h00000000} /* (0, 4, 9) {real, imag} */,
  {32'h4411a05a, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'h4447005e, 32'h00000000} /* (0, 4, 7) {real, imag} */,
  {32'h441b92e6, 32'h00000000} /* (0, 4, 6) {real, imag} */,
  {32'hc41600e8, 32'h00000000} /* (0, 4, 5) {real, imag} */,
  {32'hc402110e, 32'h00000000} /* (0, 4, 4) {real, imag} */,
  {32'hc4494d8e, 32'h00000000} /* (0, 4, 3) {real, imag} */,
  {32'hc4851735, 32'h00000000} /* (0, 4, 2) {real, imag} */,
  {32'hc4a669f7, 32'h00000000} /* (0, 4, 1) {real, imag} */,
  {32'hc4678276, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hc4a2af5b, 32'h00000000} /* (0, 3, 31) {real, imag} */,
  {32'hc4bb190c, 32'h00000000} /* (0, 3, 30) {real, imag} */,
  {32'hc4a53da7, 32'h00000000} /* (0, 3, 29) {real, imag} */,
  {32'hc4e95e66, 32'h00000000} /* (0, 3, 28) {real, imag} */,
  {32'hc4ce6cac, 32'h00000000} /* (0, 3, 27) {real, imag} */,
  {32'hc4d3dac6, 32'h00000000} /* (0, 3, 26) {real, imag} */,
  {32'hc50da333, 32'h00000000} /* (0, 3, 25) {real, imag} */,
  {32'hc5197652, 32'h00000000} /* (0, 3, 24) {real, imag} */,
  {32'hc4d34646, 32'h00000000} /* (0, 3, 23) {real, imag} */,
  {32'hc4bba893, 32'h00000000} /* (0, 3, 22) {real, imag} */,
  {32'hc46caab2, 32'h00000000} /* (0, 3, 21) {real, imag} */,
  {32'hc4839b64, 32'h00000000} /* (0, 3, 20) {real, imag} */,
  {32'hc4ab2f53, 32'h00000000} /* (0, 3, 19) {real, imag} */,
  {32'hc5022d2b, 32'h00000000} /* (0, 3, 18) {real, imag} */,
  {32'hc4b33496, 32'h00000000} /* (0, 3, 17) {real, imag} */,
  {32'hc45b9b9b, 32'h00000000} /* (0, 3, 16) {real, imag} */,
  {32'h421b6b20, 32'h00000000} /* (0, 3, 15) {real, imag} */,
  {32'h44710f68, 32'h00000000} /* (0, 3, 14) {real, imag} */,
  {32'h446ff822, 32'h00000000} /* (0, 3, 13) {real, imag} */,
  {32'h44adeb58, 32'h00000000} /* (0, 3, 12) {real, imag} */,
  {32'h4483525a, 32'h00000000} /* (0, 3, 11) {real, imag} */,
  {32'h4441ff01, 32'h00000000} /* (0, 3, 10) {real, imag} */,
  {32'h43e8f980, 32'h00000000} /* (0, 3, 9) {real, imag} */,
  {32'h4420d705, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h441a37ac, 32'h00000000} /* (0, 3, 7) {real, imag} */,
  {32'h432694e8, 32'h00000000} /* (0, 3, 6) {real, imag} */,
  {32'hc26de888, 32'h00000000} /* (0, 3, 5) {real, imag} */,
  {32'hc4535496, 32'h00000000} /* (0, 3, 4) {real, imag} */,
  {32'hc4809771, 32'h00000000} /* (0, 3, 3) {real, imag} */,
  {32'hc48e048e, 32'h00000000} /* (0, 3, 2) {real, imag} */,
  {32'hc4abe468, 32'h00000000} /* (0, 3, 1) {real, imag} */,
  {32'hc45e1e3b, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hc4b7f144, 32'h00000000} /* (0, 2, 31) {real, imag} */,
  {32'hc49e8b25, 32'h00000000} /* (0, 2, 30) {real, imag} */,
  {32'hc4a5936c, 32'h00000000} /* (0, 2, 29) {real, imag} */,
  {32'hc4845c2c, 32'h00000000} /* (0, 2, 28) {real, imag} */,
  {32'hc4dec616, 32'h00000000} /* (0, 2, 27) {real, imag} */,
  {32'hc4cfb2d2, 32'h00000000} /* (0, 2, 26) {real, imag} */,
  {32'hc4b26736, 32'h00000000} /* (0, 2, 25) {real, imag} */,
  {32'hc48e1de7, 32'h00000000} /* (0, 2, 24) {real, imag} */,
  {32'hc496a273, 32'h00000000} /* (0, 2, 23) {real, imag} */,
  {32'hc48fd00e, 32'h00000000} /* (0, 2, 22) {real, imag} */,
  {32'hc38385b5, 32'h00000000} /* (0, 2, 21) {real, imag} */,
  {32'hc40689aa, 32'h00000000} /* (0, 2, 20) {real, imag} */,
  {32'hc46baaea, 32'h00000000} /* (0, 2, 19) {real, imag} */,
  {32'hc4c6aace, 32'h00000000} /* (0, 2, 18) {real, imag} */,
  {32'hc4a22f33, 32'h00000000} /* (0, 2, 17) {real, imag} */,
  {32'hc459db03, 32'h00000000} /* (0, 2, 16) {real, imag} */,
  {32'h41f24680, 32'h00000000} /* (0, 2, 15) {real, imag} */,
  {32'h4449d8fe, 32'h00000000} /* (0, 2, 14) {real, imag} */,
  {32'h44a899fc, 32'h00000000} /* (0, 2, 13) {real, imag} */,
  {32'h448ed5ca, 32'h00000000} /* (0, 2, 12) {real, imag} */,
  {32'h44ec1b12, 32'h00000000} /* (0, 2, 11) {real, imag} */,
  {32'h44b163de, 32'h00000000} /* (0, 2, 10) {real, imag} */,
  {32'h444c7709, 32'h00000000} /* (0, 2, 9) {real, imag} */,
  {32'h444d0d22, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'h440faf44, 32'h00000000} /* (0, 2, 7) {real, imag} */,
  {32'h440536b2, 32'h00000000} /* (0, 2, 6) {real, imag} */,
  {32'hc3a85139, 32'h00000000} /* (0, 2, 5) {real, imag} */,
  {32'hc4819f95, 32'h00000000} /* (0, 2, 4) {real, imag} */,
  {32'hc4511a7a, 32'h00000000} /* (0, 2, 3) {real, imag} */,
  {32'hc47098e4, 32'h00000000} /* (0, 2, 2) {real, imag} */,
  {32'hc438b0c0, 32'h00000000} /* (0, 2, 1) {real, imag} */,
  {32'hc4a14194, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hc484bd02, 32'h00000000} /* (0, 1, 31) {real, imag} */,
  {32'hc4a43b0a, 32'h00000000} /* (0, 1, 30) {real, imag} */,
  {32'hc4a52c39, 32'h00000000} /* (0, 1, 29) {real, imag} */,
  {32'hc4acd73f, 32'h00000000} /* (0, 1, 28) {real, imag} */,
  {32'hc4ac7c6a, 32'h00000000} /* (0, 1, 27) {real, imag} */,
  {32'hc4934890, 32'h00000000} /* (0, 1, 26) {real, imag} */,
  {32'hc490da67, 32'h00000000} /* (0, 1, 25) {real, imag} */,
  {32'hc422bbf5, 32'h00000000} /* (0, 1, 24) {real, imag} */,
  {32'hc416fbde, 32'h00000000} /* (0, 1, 23) {real, imag} */,
  {32'hc453f4b4, 32'h00000000} /* (0, 1, 22) {real, imag} */,
  {32'hc3fa1d16, 32'h00000000} /* (0, 1, 21) {real, imag} */,
  {32'hc351e070, 32'h00000000} /* (0, 1, 20) {real, imag} */,
  {32'hc4108f13, 32'h00000000} /* (0, 1, 19) {real, imag} */,
  {32'hc48bd5f9, 32'h00000000} /* (0, 1, 18) {real, imag} */,
  {32'hc46f6729, 32'h00000000} /* (0, 1, 17) {real, imag} */,
  {32'hc4661022, 32'h00000000} /* (0, 1, 16) {real, imag} */,
  {32'h439a6f66, 32'h00000000} /* (0, 1, 15) {real, imag} */,
  {32'h44820e1a, 32'h00000000} /* (0, 1, 14) {real, imag} */,
  {32'h4457ba76, 32'h00000000} /* (0, 1, 13) {real, imag} */,
  {32'h44ab2c9d, 32'h00000000} /* (0, 1, 12) {real, imag} */,
  {32'h44f669a2, 32'h00000000} /* (0, 1, 11) {real, imag} */,
  {32'h449aedd2, 32'h00000000} /* (0, 1, 10) {real, imag} */,
  {32'h44a46ebf, 32'h00000000} /* (0, 1, 9) {real, imag} */,
  {32'h44e2eb16, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'h44b80723, 32'h00000000} /* (0, 1, 7) {real, imag} */,
  {32'h44b83a14, 32'h00000000} /* (0, 1, 6) {real, imag} */,
  {32'hc476bc29, 32'h00000000} /* (0, 1, 5) {real, imag} */,
  {32'hc447d146, 32'h00000000} /* (0, 1, 4) {real, imag} */,
  {32'hc4c27d16, 32'h00000000} /* (0, 1, 3) {real, imag} */,
  {32'hc4939deb, 32'h00000000} /* (0, 1, 2) {real, imag} */,
  {32'hc4692b17, 32'h00000000} /* (0, 1, 1) {real, imag} */,
  {32'hc4837fb6, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hc486fdb0, 32'h00000000} /* (0, 0, 31) {real, imag} */,
  {32'hc4a1a8da, 32'h00000000} /* (0, 0, 30) {real, imag} */,
  {32'hc4e606f7, 32'h00000000} /* (0, 0, 29) {real, imag} */,
  {32'hc482bcdd, 32'h00000000} /* (0, 0, 28) {real, imag} */,
  {32'hc4a60c0b, 32'h00000000} /* (0, 0, 27) {real, imag} */,
  {32'hc48ef37c, 32'h00000000} /* (0, 0, 26) {real, imag} */,
  {32'hc3e87071, 32'h00000000} /* (0, 0, 25) {real, imag} */,
  {32'hc3f44ec6, 32'h00000000} /* (0, 0, 24) {real, imag} */,
  {32'hc3f09116, 32'h00000000} /* (0, 0, 23) {real, imag} */,
  {32'hc3cc47a7, 32'h00000000} /* (0, 0, 22) {real, imag} */,
  {32'hc39e2d11, 32'h00000000} /* (0, 0, 21) {real, imag} */,
  {32'hc30b9946, 32'h00000000} /* (0, 0, 20) {real, imag} */,
  {32'hc38f908e, 32'h00000000} /* (0, 0, 19) {real, imag} */,
  {32'hc3199e96, 32'h00000000} /* (0, 0, 18) {real, imag} */,
  {32'hc333b1d8, 32'h00000000} /* (0, 0, 17) {real, imag} */,
  {32'hc4097c09, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'h441a0f1f, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'h448c4a2e, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'h446ee6fa, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h4483c453, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'h4450a90a, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'h442678cd, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'h43d94211, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'h44868972, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h4420b475, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'h43b1ad7f, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'h421f7d58, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'hc460176e, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'hc460b4a9, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'hc490e786, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'hc437a788, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'hc42ae10d, 32'h00000000} /* (0, 0, 0) {real, imag} */};
