-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
O2oShzPUNdaj2K6fhET5SnDaNKEgHDNst4TmzIjPCYOdgAKpJ8ft3d0U22Z4BsBY
GU6e8jj2zXxb2waH4WSKPnuTcWQcuknL+ztIHAMdkbEr2+n9pAwOl1hgbY0a1Jz7
mPEDwbL6y9t0AplpLfNst5J/JONkL4Gd5Whnda8qSCr9C62FAuuL2g==
--pragma protect end_key_block
--pragma protect digest_block
AG+DD7VlnqbSOEB0AA269XxuJ4E=
--pragma protect end_digest_block
--pragma protect data_block
q4Ysub4FIiEGhpZIWTOeEytJ4gacJUw9BZKcaiaDvf/8zuw7+d84216HtfvQBXgD
8g8yqBGcezVSI9deLudhf6+yWrNpbeY2vuwzLwehTo5M0iPceNTx4qs7W7uaMxcc
aiuYx3BqFnZN8h8Jrj8L0H41aV8WVG1FPh2fQOFW+iHjBL3Dt4aKoR3TOi6nsUlF
w/NbOjh+0H0pWbEPqKZZ2MpIPhftnjvsUunRdkAL1THSuZb9M5KDjaz/T41H4Lko
JthbpdVsjBrlFI0CuviTw7OCHxwvOnP37/zpDnseNv9v+MTTV6DEFRN8jdQVnN83
P0okXY0kQrampEzJXQtk+yyREnidTVIjr30FW9Q10DVRtVWKr1xthZSuwur7hz7l
C2+V39xqSn1bsyQ3hDSIAOkOLAWGSUSj+pkkfLY1JQcEpbgzOiC8GY5L9HVf2RDy
CKj1hS6f47XlCicoW8YSRmw36Inqed2CGV/ydMfhqOet2vSP8ceN7LZbNSWlw8lp
/0aXxNuQ8BJiWPY1wwRJ8BrrgSmdEXw2aAm5R4ZLcHqylk0AjZL+SEFMSPGy/6HL
uqaiMvbYig0LEtxW3ZJ6zEP/iY2Cnr/lTuBsm9Ep1cKKWlhcW/56LpoWc2pX10cL
X6d/NqEumbyhkRt4kmOTxDJb/nO3F142yRU/Fh0C/qArhdUWALStQfloMsuUaIHB
jrNi+tFCLMHBLSiTRJwQvRXfVt7SD+gKbgroXZOAl0QIdAa3edlAYNj2rCbKUJWl
O6DP1xyxjJpr9wER3RWMMLvdb505RO22jSRzihridWCPrz8tquGFLin3Leo+gdOQ
1jbOMg+zbUm4P8hMKDomfh2fnc0/0kKUyaIpOYvrnzrOq7JSz0qhGJS2Ns3bBjG9
9zlCrAiuooVZniLn1bzqqr+5cAAplYSg3h7LFsm0HWHpeZXxGbhYFrEPNE6CfKtu
IOhNo46Sm3tV6I23emPLQxe/te5/sZPv4D3BCD3RNaJO01CcXAv4O8vsAkesMbcZ
7MWv3A4td06kBy6Ea9kxtKlowUHSA/FOWcTmZjO4LY1vbjBHu7lUSvqzLzv9PyxE
C61HZwyHkZfi4tJAlsJPPG3iUWk1dt1pcTkABkXfzAx1nzB/o8gm65ZtNGfP3H4c
wnHIkL9hbNS67AQp88CL+AcLPXb72Kb+SWuIFrpsF/gt7HNCTSBaW9lVFuH8Drng
uWyur5ygZh35Yap/FDYT08Id5YMWQzTuEEybWkdE4FjhoLGHMLYRr0PnHj6Q3DHk
YE60gyWTaXgCFreFFKa42XhuCh/E+48GzWILRszRTtKirlbpOR8FLQw+E4VHCr5L
fvsi+LPcqmDla4KPRQOl5FOAPo+lBwdeuGi37ZFE1tRRyC4nYIupmvssdv/zQUoh
/HxI1+dTeS3Ior+iDQFl8Qb/843QaMMJoegDg/FVf0zTrQJS0D7Wb3xGbRvzpjWH
XsqMexifoKpQwghMql/cghfxt8BDneRW0r4t4l1FuOaX0aG2xsld14cxcsxJ4AXf
JcHCbmgBZ6RbrqY+9GdNdDUzPZYF/8wHgqKxWu2dOzm/GWQycJNNyirYb6WyYaQG
nLu5p8GZHb/tjAkpl1fobFJomsQZHqcdtFzDY+AJLihYxupaaQS8YRT2TsCfAX48
B7u41/7SpQc6AQTZycKIiJFkHqwbk6AQhWak4H+HupxzxPwvyNjfcgftFJnjgxD5
isCDb9b5H/nS/qgD6Uuj/KlGBPbfIPn57tc4vT12hHSlHqdhYzIB31rf0nbkmr6f
zW2eEwPZYsudknEnWOzoa3Gt31g/A9M5RSH2PjkBTTTA+wYl3dSckih36XzGzcby
cu0QhnVuQ8oBJiRHkDWBjZmh3dzfCw8/JXFdG/r3RwH3MQcNplYQcet3RjB+Yefn
RWD+K/E7dbEsoE5uiBfFgLG2H2mnZ9FZuwvK/xTbqFat5D8FC2JPX5rKQKeUS5FB
05YaOoRCT0hL9up8MsgPtTKo3qPjAqxzVKWiZYM4VjBATCNsfijFMZJhIMrG5Gg/
7RaFfbw56dC1zwIhX5LD0AMIslCwb7yYUlIbyGGqfKr4huBALtn7CHLBSDy8oh+B
HwWq+ZblCXJ+Bj2ggqYa5ulvZlnbtkTIfhaZK9E6BAHAlN5CQicu9tKyHX5VYuHp
kWN2OMnH4X01n2yElHP38BB3pMD9tKgqGj7x0/8auVJ7Rdh4o4KIgI6wXVEF+007
s/kaCFEwIJAMVCnkmf5Uy8VP25on8ZF9Bjc7jVhrCgP58nw310VRClUY9jEmSSMX
710ClnEcVcsyOV8bcITynW6NkTeQ0o3uy7VnuYcieKcgIsF+15w+MAEUh7GcxUb+
UMpeR8I2mf4L1x0XC34x3fnMS/CfMj7X724cgIvWMjIz3t93YUf6sIC9+rtugwJz
eTcHuCekOR0ddIi3pLtTP1Sez7jXEOGHYxt2tMJX2Nqh6EfYx5UB8kGO/uMBtpcT
Hc4V2gDW22OYbLml9G9MBGAzYEhRuWSh0IvI9G57Qf5NHh6dVBNld+MFdqQQiyoo
WgKk8FyEO0CUWdvjWZMTYzYdlUHJohffxJLm2VCwcjBV/DcAu9vbMn6b+E2GGO3O
zLWd3OreI3u6EIxviHVzq8d+KIbkKPxp+k/GgtUbbwOeiIkHVyNPDP6CoeW10k02
npeiA8p4COYH8LZFccrxjqnTXyfBHO/pfG63R7iPdqKqlbhLyehwH3wnPXfPhntW
Fo7U9RyWHCNlaOzyqbpakn7X4BV1D5C/QXUwhtKyA4jHp3uP+7cWoGAaTQYNox4r
p1hK+orJ6RC8VcQAgzGKTZbOmJvqNkT6E4MSBQcP2vIAa8tqclwScGV6BvEIGwL8
jS1orTv3waCdqEkm6cw5KQmxw9Klbf1YkMvkX+MglSXzwPKoOjdIK1iBEOzB4O/N
oNMm20USuJsw6RhLy6hPc7cPPvNSDi48b7xhLWRtiPXtLJ3k47rtmEvY7wpAnNyS
VZH/WDqM44Cr5v1f/rZ3TQxDOjRR7Hx0yKx2824myATAvCkqTnnN5vGdL4lkWJVs
yDJ6/zUD3wL8AflTYGNowtz4mQf+DUpYAKnpcJs8OuhS8bHAzBVN2WtNpm8ryrkA
B6nl3OgnDT480SiX3AX/0iWSnvXmSVgJn5I41xY3jTCiSlYQRdU2AkEKEXI9k5Hi
6eH34QpVtPpFVvoo78lzhyOZ7FPVJU73iItJiw2TTXlJb+BKCxrrYaoiMdc26+GI
wriPAoZTaBt+ddIN76FZrpuHEMZA05xJyrdd4BybXHxvnXjv1z8FDA/JyxfYRlOu
K7uQYAPEPrV82NWgVtwIiambr+50cEba856jZvIqQ60W19laVLZMe1qzt+QfHBsi
XHKYN2YwS+IWL7pbh5xYD3GW8RxWBrSsSKFmdgGc1UCmDYbbAR1tzEiZecUvXYb7
XgTA3Ruth5LCqrX/HJd6pkWpPFM46roJ27cI4feZm1yAjAp2sXVTWhUd3f06mLa6
TeTDutBfdGMKfGGgkGhRBZkXUqZ0dNC3OD9fddIVsll3dimMYXP9r+DNJYbgZQ0W
3QZtLFbhDZ+wU3FE23S/2eBb/0eVkEl6nLqFeWwi744UO8sfytY8+Td1JMmpe6DO
TRXsLE+1gSwpTXsKQW9z0poOwiBhLd+9aENf3aIEO7uGJqMaEEgmP86ehNWCb46O
TkbUQr7ZkbSHl6oMfJVL9ZgoqM1N71M1DiK2hw4VcbE3ZaidkXcFpOe8Fgm6rwqN
4Fx3jSWaYkZ7KB9iAaNZqS370q3gU+DDvxKqLA4zXRcKTvXA8h0dXy1BYycfXdeC
cfLgEmRuuYA+/vcFvqqjzn7th0NX8uGDFiKz05Y5ankIDWePEShIDHJgdPr9vzGH
pTrw7sBBanvqWJ/R2NyaKhM+LrA80aq1apdxGf6aJqru920W7oOfXER9fCH1DwBx
yYnAMHhPxWQMn+sEjwyyfdyNNW80DsHbGrXB+3A3pjg3wEQ8QdxBJyTqQpgdOrKX
UrlRTkI21fNCoEl9m2BlDv+Y4rSEHmOp//jHw1syzjXDiC1Mboob+ebHndw49O6F
LEIMMtwZHdPa3j/VknyHXKp3OAuPdEP93ty04hx1RQ89+WbKpB1ofuXfnYmNF6Sk
C1XuZZYHKCJDexH24SFmNs48XOuE2UVqsQ4SW36v83278XTnqpjeJSd1eYHzj+vr
+j+m5JeIhTeUGV7hJT+qANHrGyBJRn14cBk0lgTw7lsYRIBUQX9UlTMj2TjUSdgy
jY2/Bt4btNREDSYZ0Z3YdWi7b5/MvkXjecIF6y5Po7n4ZzJ6M78wd/WhVmSmHxjF
b3QijnCIrkrnJmhNoEHlpP0MMTbzyAwpCwjXh0XplRB9tUcJh2C4RdhE2XityG1O
XBULkhryd2/mhCcpJ0UZPolxHLee8+JT2WBraFyWE89EF4VQfZG6EQNl9+FNtLrf
hLidUcExcR+GFJoVlIPvVcifKGv3qZg9+hN+sswnlVgkcmFaFfRtgb1JFUkHmigV
imekrd9KDpb1ij7b/eSXCP92TnW7FZdaHqoMG7obdVI00dUbJ7Qqr8VVAjbD8jQz
vYdpO7l/zfMZV0qpWwvyR7d4mqo0OaL2GVKdGNO0EyMenNdooEkaf3mayNctIUhk
u/StLSpnghFHCetCnxCgU3XQfjnD/NABPGZutjr48qx9YM6N7vqEaF1LPwu4Evbx
A8SkWxvW6iPALQv/iMRpknMEh+6r1Iv/J+KEWCeqQQ5N2OaL0j5O1d5WINwbf20f
5tl/XumdlfFm6E0UtfogBM7XOwqXBO/QFraNdqNAGg6xadpyMHUuWYU27Wxy25vg
22URmqoJGwBqBEXqzFhMk1h9Ht004cM33IF3eSUt3Lo1hT39liH9YieFR6M9rS55
mMuLXs4gzqG06rGajWCKjqB2X7nnLtuBpuM1Wp5C7S545j7dywnok/vNI9dmo/X3
NGfRmLuq3nH+E59rsVojDeFuN0KHQibaDh/4v/Pv3d+55a2kodj40E6HcXmLcLaq
WXid1HHoLk9PFgJJZsd8YBh4hApB2xt6A/jB3EtGIt+FS2/X/wKKVqZkbDDVP4qh
5C+TSUy4O9qaa4MRzp9PdVIuh8p75N+D6xi0XLUv0MXTHf6YWZH7YKIq9LppOzqK
HrMs941+Pl2scj+K0ITE1KjU/EDfXA3BwPJpctaMU2ymCabDj8qVVHmyUQBTWkDM
JwtE5TewIfbyKs5G6vKSqUo6sowCFz68X3zHS0WaMsU/E13TbjtpuV51IbLXlyUz
gDzH/+3wPHQ4HetA1BW1TjTutLprM4HweI++isMSGVRKcwSoPfCiMtCAyXwgOrmG
kCY+skHYD11XWz/fVtImQ/hwm7pLLinN5kNFHsLOGnDo67WeMNh4tZjKFO4IP+hJ
jN8J8UEIUsCpYizWAGSrA5dBqg/03pw0RuDlRmiQGEAW20dHjFVbvRUK70yLkzzz
ENYtlmC9ZvsF4MHRsEy+j/Sziax8GZ/zAps0MYnnRgsMHIm/eYIIotf0tDA931zY
iZ+aAsq249+OejDav8CbU04onbFQ7UlngZn8erQe9P2LLUvaYzwhvUM8rR58UTp+
o7i3EeO92OVZDkioEN84aaWHxUP8LRMKU7Lx+2UQjAlR9DrLacDVkmws6ogfR560
Lztmq75y1832cBEOsxNtgwI1ahz56n7lw6QIeGqtlrqPEQqEczo+jmlUvy11ks6s
++qaOWR2BTeFMQg95WDaAh80mCDBi3BWAFYVqCSs1IER2jItyWFfEWtegNzg0eyi
x/kWUsAfFU5yQLs7IDoJhsB/LUSLxctPDVN+wu7Y7M9fw7lBxcOogKXQ317ZSyAX
ddS/vKMhqvH0rviWBQDdVqdqqeKELynVlmK/qin0LsgegWQfBKRUYfdZwLFMH9Ur
j2jWpytGC+il/mbKagc+TeUHB+TO2CrHNuegiRES1rlZXFzmpZHNb39f5qkH1XJ6
7L1BW5TWvD6Zm8mNJ0uc/BIikgY5dzsSr3vWLPKl++COi8SG3X6dvDOVsvoOmNcQ
D9dgpP4K1W5QGnZRAoeciUxUcFErF3LE104wwmvDiQE0hg2SXXMBB8YIjPD/RGSZ
MRUMiRHA1WPSesjjmBkxlzShxTr2sks5nzSEHj6CAFguNqFGKtI/x0yRiZ4L44EJ
+ui+OZuXDf977YpTvhlJKlrrpf19E3HADPdy3KW1j6asPoC2438J1GSnOd4AiKAE
fvLYX0kUv3/tDN/phpXbnfP/EOLMtU+3/vavDN2PVOvISYdBBAhJBjMVu3vSwQ1D
KxzFnTBhdF3dWsRG7br85uj70MKHIyHLXRHwFSIUWbs=
--pragma protect end_data_block
--pragma protect digest_block
3xhUkSQwHWkBK+WhFRlwBO3H/Tw=
--pragma protect end_digest_block
--pragma protect end_protected
