-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
r/Q2piqO2yvgdnMc46AAuKceOG0o5wkKpWnbBxui4Ss42UDq9aGi+SjRqMSBwXF7
fEhQ5qOnI2iXys8X+lkdHThb78njwVlBfoXf6nto1ccuXKKnH/BxzRPJCkCWYAHg
81nG2Ae9T4TyDjxV5dNIxW4Zfu8YYhpUx1pJJNzTX/Ej4RGXukToMw==
--pragma protect end_key_block
--pragma protect digest_block
OrY3hwdfI1dOv62nAOxSVzhbuZw=
--pragma protect end_digest_block
--pragma protect data_block
mWNyGddehGYmUrDrgnJ7wwys7QXTua9yj3ksO2rWmbdAl5kiRy6zeYSjk5n+dqWd
MwqBgxJVtONu4dG62Tl3jP/yp6wvTwy+WJW8qh9k9YLguT0WbQWOD0KYNdW4x/pj
EqzLnIZOAgOJoszMggeoYO4z8aRoPRodeOqoT8xV0UVVtl+nmJ3rvkHo+fS40aZY
a6foFk3BLtoh2oltrhxvsZGkfaHTj0d6sjrof9i0UT/1PcXvjUj5SzgsO9j6jzL/
grr4y9txHKbPv/uQRyHNaRz197c9+kVKCk4AnItW+m9/31f8tFDRM/1C0Z950BCg
fL+VkGdVlvBu3XT6L/L14aG02OrexZVZ/+aTt8RdtC6+DLC7WLBHvzip8uiqaU5m
xgcvMD0u2vbT/ICg/v7W+6+nlx3dgcjaqNa5n3ldTDZ/rlnhE021IFIzoTaz93Fv
gZrxzz/EHQcQaOdbwlD+5+ORh/oUvbcUJYS7MKOmR01G1aZj117j8vcDcZwk1eU1
ctulMBWh2Fq9eJIr++Yb4WaJrP27X3ZUDPaHPFGlX2s2KRRS7V7qaBMSPi+ruU9o
lIH5+xiK/hYu6bc0/oC6Z4fUjx3fxxdKeHTE8UOkryyItg2fsTNwHKAx5iU2qcG0
Kw538EuBaQ6v2BsHHPIGjcT4tRiiOP3FM0+WNCxK0G8j7JqSS63IZOvoMY3WOXO9
SVMhrXkYe8JeXe2oy8LW3EwDFiei+OOF5m/aLYJaYSsqPdUMhAPM2jJos3GSLPrn
vQGllWg9Y7DU4zNkeK2O59aLQVWBlU2Icj+vQv9kMtnRD+CmiODDbptqGbuYHOTo
ggDzMSkrEJr49XIqF4BTG0A39TncnLuTdBgjRIs+iVQckFrdaqITMGuUhWt+MV8x
uj0banhV/JF9cDPY9wpiu0Exw8Z3Rq5vgGjKlCoNfO50c2aG3ohqal2/MhB4i1gy
sGP5L/nsa8FWTTmu30xwNZfgYKIcbT/ZepUCcLiEaM6qRwsSLyXYtciMXt62sDKG
Rp7u7tDW30Mz/8Cyzmc/ubMgFEH/i+YFvbcjWvUp4Nx5oV9lfP+Ulqcii4BWV4bh
YLVkhLqSOduW+3Jglhk8qhcHjG4IgCsjKMnKQqaFbIw1BrF5AE3wsQi39HulOVZd
T64ysBHXV8d6oKHpCzkfKJYlFmUsv3QWW7Vq96ubXtZ116hvRwv3e59huZgvU/su
2W9YCTAjenWoT1p64cqDvI9eb/8C8EJetiHIG651mRaahM9sc+oRDs2a33D6DCsf
k33K2wVyjD3FlVW1KX227600kCniQW6WUDrUX862emdqGE7tF1EdyaN2a17Lwedm
1+6rwPzZ4vn2WeMFLbRGmrulrG2fCdlHm0mV4m4PdZ7eVTVd2VpTWGBoaOFb/a16
uhn0/JXnAQrFq0kvxX3pjCK9eppCQ4PLusfagrP+mftwMD7ST/+snvYXrrHKZjCs
S6jUXAUVFEcmit0vJPwrhbZ/0UKz5ADCdfQO8NIEc9Sf8bBqX4HsYxpuF0jR6L+h
xtndba6bZtQg/BVtsozHCu1VoXhFB2z/H5lpfA+9aNkK9TrJ/8ZsgsCRMk3pSLN9
xCbJpBc+V95R6WQN7d9cZHjIi3aeq0zYxxy0SRoh3GGdeDIdDHK+wyVihAYF4aY9
VLoy+iWO9KEWxHAdd9Kvqdqff5moBOLPAa3+kJSoa+l88hB++ERV+M3nxYnJIjnr
CGRd/JhOGjaMAb0nzx/Ys4JgiFw97aC8phfNQK5RWsR3A+p7MJBwG3zC4FzF1GUA
j8wKaURSxqHuLNO36uEhq7auqBwpA+yqu+gDfQscoqIyNZPjnJpztXkse9MkKQFS
Sme1pba3e2Hvdopzo0rX3hqWmfGTDgYsZCovg6IAXSSZeDWb9V5Z0Kd6a0x+ZHTF
2HMGYAbOSGDvYEiXfV6zpH0mkGxEoilT5RXDyu4zXhvqrKb4wjUonfHZSp8CacEb
8l7VTHF7ztT3LUu9vquyv3OvGFXOeiJu8mdBVSgwUQbTy3p1rzvUtCC4U5UbB1wM
qIjwFDrXMDQh8RFK7iJY6v8Zj4+N/OzFq9y3clym9nPm8CcatSRkk+8wEm4/MFoM
5llC5U3QjMG/ZfoEQPoVp0UBDwlrmH0jmNF9NfwjZg/BME6iplEsoW7jF8Ljtw+j
1xsUGtwL9rps5PkUftVL4TM3B9YhSSiw9e6y909IGWac7w2vdfr61PBJsEtvjAO+
9ypYbq7LEzlpuMSIpmiN7aQv2P5jOnYtQD5dMq+csk+RigH7X53Q5sbRAlb/HDuq
qn3VegOKXuLhtr6B6hQyoJaGpCEoVYZHC6Mf+pqTrWlpJmuj++EWNL9HUlU1NIh3
lOTIZJeRWFNGj0spYMBYzEM2nBMSte9neNG2V38Urvd1nRDv5RanTdoCjd00O86x
boXFdE4wUsAIyczMxXV6nqPx+Xc48MxjHa3YnXXDrR2hg5VBDYTBNwy1UCA0Ot5J
uNUBvUhNQrqGN1CtZCWn+qQoBkEhvT92xAHbb7dRs+NXWjdzAjgLVd5bjqQPj1VI
11jOa8MO8vFNuBCiqrDR3H2lw+aYnNnVTx1+4p4EXjsFDOhO5r/bfxvjy16giK+g
CZJE6H1yl/PpoHqzmQPpjUnV2GbYJxjZDM/yc6rOSX+Z1zBU2VfhygdCqY4WQ2XO
xYuAYcXVpIRtySKUV4HqYZd2iMrv8tXTvO4ye3EMQdBcZCTfONGr3fAdG0ooE9Kg
5/DjRMrbUsHULKzyNgZWpHGTt3Z3P3MfbHHsmPdZJmqrMFTW7Z4Oq7i3ZrnSsgC3
YJdXXxjrAtnaqMGoRLJ1+vpYrQ4PKEAXDOhvrydpOQlBmdaCZkuMyN1K+1+EwpAy
tYUw+d9wIVJrSBtdYaw+I4dseayy9ItqoqZxWq19rWGycbVqF84FJi/i38GebWpk
Ix3VRG4bHk1uwDP7qh/7aeyn2dwIw3LxoJrx78lhiLylgi5iU3KPq7NysiSS2N19
zlDyHhclBzTTr8oTURBbU44v9poWFmJZiRYilDdKs9YYiT7JTELMfr11Vk7rvRJm
DhlOfxe9wqqA6y21qwiQyu05P+F1ZanpSehEPjR6HIpTwoKO3klBkXkGy18c3bYs
T5ZnCyYgF1VzGcuxwseQI7jtwaP74R3O7c6XxwEz5JerM12J5gbDDrH0ovZaNIVG
D9NeTnfGgULI3Qz817+mf2TlBnxF/cHQ552hlQKcW0lfiD9MBxOR3CH+YLHiC0wl
0wsGHJ07GZ+6r3iSFDIZXU9ZxbkuimJHtNt1uFlAgnmDVjt4Sq6ae3dyB5KjU6xm
q6VGMGYaIaLjQVFVKK77+F9HTZYUlWLUYSEasGkyANEwwoPtak1TbzvkBZmUUxZs
eFC1CHkUEvX4pihFLnefZRvwLt03vAHYxF9Y4trdtBYbQaSkfnk4oVVKmE+DXK8m
Jc4vxlPHlRBRNKRbQ+qvyRHPIxHK8mb9+067wa9k0jPWh4sqtki0kOGL9fuUes/b
e94v2NMcZddostGAMEB0638yhbeEpSmWL+/y6PbSjlv5zmJr1EHu2R1DOA3Qh2Zp
oJDzNHVufXhQC5zHZQXO5FaMR48ROTiTsbW9/mHLU555P2ZbOepAO4tUcxOLowkt
YQQUIK/LII/fbAoL/Ky5WqpB3gtboPIeJrqN8c/DIEHiHAkkhUK89HccnCnDh8jV
F2DCEGokjeQZg1vAhfNbKjPNckP3kLnoepHiH+FhNiUD+WLhtTmehmvm5tz6qkzw
Otppq0kSSkLbIdRmczVAx7DbdZwAjesL6NZUQCqlPWmwCgSapkzD0XeZedxauY6A
csYR6KJrxap/h3sxLSOu4vPZ+fFLyJWpbNESsE5gO51QlqD6bo/yxTMJRgKp+zZX
Bpqsv2AFN6tO2/VG7biTSxqF62sde7BbCY+kfoli0KBMdBQSh8V8O6qctGbLuT6V
Sa15a+EYY8wyG5PCHz07hZ9lgdteE/eBtToOLdY/MyWLUCtKhFxKR5/Jt6PJz7tH
1TPgioLlWUh58ZHZuZHkl9R9wKsa2NmnZxpv6TTNB1a4EaPY/vs3zxYyl4OzhSTa
sY98I1De/xdovnRMovADPyZ5F0xrLS2fGlKNB5n9we2r9jq1ym99Yi3QsbDlIBUx
+hYUoHDgG6JuuvHDJttfBWTP8htG5B6IkyA9s/ya8b1bd8ntTGTBZR4ulgMlZciA
Ab82x36/wNOAkX2WMu/IssiFz02YzwpWhvc7ZZeVEJ5APBvX7aiW6fGz0mhKwZz0
lDNXjZ0XkAObH9Wtnz8XhepNsI1y1q9snjvEGrw17uFw06KltGL2kO5yA/pttrBF
ov9YhB7ICaTvQMm+sWbZIUOtK+ZSawzAEXf5nczgPX7c9IAmoOfjOHjEcLsz48Af
5c179ETaT4xJLjPyx+W085r1rMl5aH1KpZfc+2VP9JfIx+ulNiFjZzeQm9j20TT8
3Ks7tgipycCcd7LBsowCkq78bpZ3XYR7l1Gr0YHoOfOww6mf68vfnzAcRrhhDw/b
Bq07iaBUNpsBVZhAud4U822fi/+/eDpuTRBYNwJMGnxo57hjsTkNF8IowCaTL0X2
noJ/aw52aX20DrHDpkYLNDy4NVLgHo4YOx0Q4fNMK+PolGYDBq5j6lgrbYggzrOa
59673CpnwG4j1IjQl2yNwxgwMOhnJ/8uNvaeUF25q03OEpiXH9/NhfzWzhObRpyC
Ft5tbmMjSkBSbojFazKoey1lQbnCNILhEzE9aUNI+NeC3qcxrXQnvyTYNeTrFDJ6
fsc2hlWT2Rr5spm/RSP2QmAC78s3RK9TIkIupLiD9K6wFIvof9ehOAoPRnq507Zh
Nrig2oClNBX+2jNDKR+ljs5nhH3MY4lVd8F00yrPYDmctipgdq4ReXnSv9sGpiKk
CUdIYvlDh6eUreP9YGnYqeRGMrJ5c7DBuxcqpEw3uDr4YFCJjE96mk2yAPQCAFh5
KFawkgftCesqUJRfFfNeF1uYDWgRr02ELih1kE6mTO7neexPg8qllj7zDtem7HrI
/ig3nAcemp/J9PmK2/MChY3mxm8HXD4x3pfmC494brKosMVy+L1rXe20wZ4CCXPV
RblsucG+gfbfPBC0+yWmQiEbC7ii0hW+mVVYorcZKHgaa3df9sNrfII70V/Ktfib
XE7cLCaeInqGB89AMs34spLw6u7Ee7Jte84JNy10pwsZKnRGXprkPwvB3saAV82O
2Pt0KYYUTmZFIPEnMlcav/jy9jGv5n5BxPxPUmvalx4Oe4bge35GDzrNGJQtp4Dl
iziuhh/C/zZItkKqB837D45nR6oluZQZ7EfUmAI5ewy14/7xR8qFYw4bximOrH5S
uywdjor86EQmTpQojwADHEXFzjDHhxbBKpIfIqryI1SJuOzgTbtkUL29RWgCK8aV
AvLoWkx9++AFs3+5QnjUOc1eYtg4kSTsTsGE1Avp+uP0irGgxq1xxwHMlGM/Ydhj
5q3Q1bD7UL9jOLlM72OjCeViYWm9VtBw2Jg4Ss6ip/WzW8wnmNv/hbaeGBKkWFMH
9SDsjxX+wYSzvQ/UZvfRi/g6Fs2Gxn2wuzORtwl19Vbujfb5qSoDbNV4w/O5f8TX
D+93pioCXLgPxOhfy59KaBiwE6jnvoi+92Arg/MTx7TNZiDzSgjNQtRixHWC+94D
68MSCH+1Chp2kFa7v9Ih8vkmVoeDAZfBqiu+bDoJgRHa8tsYCbJLIq5rhzeeXZIx
eHjvqa72iYwbotdLECNM97oEaq8ERwsn/pId5+/F98e+edY/qBWWyGinAV45xJrF
QmUx2jzRk8blzchmWoFOWmCxh3b/k7odSqd2ITwgBry6ropAsP9WgHJS+3ntlM1E
XHceZq4MEp28ybHCghynAzFrPSGNvvC2Y3cfnW0Jho2/dD8d0p6dvx3VTppY3XOx
tEC63/kUNnuYhC7OqqQ3lIO/f/5mxcp2MN7+63BC41+s2DkrGv/3zxWe57fE+xjk
iRxlXBCzajHEWIUbPYRGvwkHrbochtbYaCATJH9cjX/ZBuNSe9fQ8juxE6M3jBJY
PCvX31CIRIMXvAYX4ni+wRRkhbtYQyi8+XaM3SYwaPRXzV00RwzM6t4bxMzr2DNm
2IKg80DZRjwZSPcr4PYanS1tAReKcPvunF58aU+qPv+pqwciu+OhajE/A/wXt2HM
+rx6wcT0PQVcG0cM1f6lNvTOHkcXyadRgy4tgLKQfZssnE7HRomP8tYh8cUZRm+n
v6+mGhVgyGvmJHuGbhgkBEnBcs4GwwWQvEblVITSXw0nmVljnbguIFOQ5n2tYcMn
v1CbEvo8GvHGMaX9R8oz6fvk4ggR5BEAHKGl2PiOWk2q3cQJuj173Tb7RCs0NJFb
RImUjopmM2/zrvOWj9Dga62IGM8J+ccEiaUukD2HawoR7BkF8t4K2n7nGQ2xxnvl
REXssvRJgVNAUj3eVlQjsvzbBuH2vCt+MuAKN1ObL3I3MmBVARUNSG7wmCVNZ7PD
rJs1HQk+T/FeW0U5Zur0KL59uei46gOmAEYsHVBwLsn3vaerhtPKg+OLsKqPdtFu
CNoYKfeqX9S4+Q0lndlN5nv7b2BZBnOp2LE6lOINiWN+4ZRjtyOkesn1+1YFbxL8
E5/bjSanl/H2X36598Tj5PEpHw7Tiv1yJJIMdxkYx1qeUgcNxmC37UDm8u+biA89
JwrKK1UV1exmdOKGMq2hlxtBHwoN+209O2pDmZMjiQEWcUzGuLBXDlUgZt+UrG/g
b/hXk/1our1nEzmT49u8Pvkn45ITOXKx9xh27BXye9Ip7DP9LJ3hj5kVYrcObXYg
DAdo/RzE7HpxRKHK5d+MvfsV1EydjHRf6i1f7u8LPBwy2vrSHiDHIRnbKYoEg14S
kLPpD89DhNgoj5lHtwQD0m/CSaYleR3ojS4OCCf99+ATl8J9+L3hxsYORnmQq13C
9Yn78uoBHOXMN9DKo/+4uDI1WUQIro2rpu8LMWAv6F2Uq5eU5W9c1ylWycX4V1Z1
IagZTJoh9htiGa2KpUOJYjKbUFgWo6rjZmJEv8FT923H+eMfoifrkv+txnhm581S
bfygwE/PjsXKgtVXAHoTUzo9uGuMQiPsoFDlPEOCpByBxq+i2h+5vZx6X+w8FU05
H7OPWw3FI0Dh8N0ZTUrt7ewFGaZWCt+p3N5NBlFO5yuiSE3165KCMIDR2Gij8geb
fEDAs41CgtnRcrRYo1cphltzXiExlIatBI7rI0rm8Wz/a3KLLZZbSbugTf6jS3D1
hkAeSjQxk3NWfQDhGNIIAfe8jw/vA97R0QmVARDXCyzL5AyizuGDvyJGjIzt8VMt
HMLZK14/ScVgIB3XtkOGr8PH7brhwdRFbI+nUBiaV3jXPcujHeBNvmqVXCqCmvI3
vtp/ZKmaHDR0qFr7Tgq0oy4Gux92JxUiSnd8iktlpm555Xgwm9m2m5pUOYt8Nq27
BQlw6z3wxpeT08gMzeZ8TdGiXojIy9IKdVTDr4ReXaQrbvd5qGe3XAkX+bIQHrkN
VD1cOPYZCojvMqryEWvoSjjcjM5qlWu+QB5BNI1QNUlGhhnlCgYMkux0ej5Scb9E
AVYty4pnKMBzu+1JcbSZDLpO1isLZboUwqY1doFiBBdPi+BN84FF1Zw5GwRwHwnG
mNAd6FKwfUzPDe4VWscqv0fCgs7sZkh1TWos34WzumgImENAFMiC9cw3LWX5M9QX
Gfba+MY5tHvbQaqFpDgkJXfOI/5OZmH19dwFtaUILpNiQaJpRSfG4/TUkf9XBB+7
Xn3kevfr5abPvtxLxyTM9d01TXEwnNA++5+xADPwDmQSZSty58gfWEzVXmhewZ4J
l31BGJJbPfTMFVyeKAzdvsej48u4Edcr6JgxwJY9Zh6YSn7P7nMMhz+w9JcCBL+X
5M698HHWpPZnGeAmJ2hViRchaj0UGPDLGbwXNm7SryGYlaUwpeRnjlUogTozsWV+
M5S8Gt6FMi0+Q0jAzOAe35zLD5+LqFZIiWLlWh4wXH/S5ZXAPnvCZBObSP5ruGMy
1T8UtNwyHMFC78eroM60+8VknpagsZVhxoYV2XpPqbg76KCy6mUCy/PGJ0YVfGf6
cL2xfKql3HICtbFg1kqHLtyRyygwTz8eyjvCsi8BbXuPs0L+x19rFCZo0LG4TeYw
1y0ddl2IvyN1BGcVnNz2Tk8FgI6q77hFwk6YXojDq+7uD13XAPJBB5BbdTt1AU9a
gnm6KSwXzOc1oLgTXBF5hnRaSviBGFjUtEhcfB03Q/IkSKaidMhIvBclM7kUJCkz
NTG2oD8wyuIspB1Gy44Sfcr/+9xG95QmMd6g+CBt3wLGWV2dXSdBfkoU8CMngnoy
JUl7iNY3H7X2cwNf6Pz7nqpy+k9eTo4vtXU/DszAXmCogby2jB8vZEGNtumaXco9
coRntwqhjATv2q1uBdpkRqN2Hh9Q2NkfttctKEGMiKCaGPx5UObDexrxoOdRGXlO
Te9Udj8Q5vcd5hYV/jiP5He3YtaP33HyBrinK66yKPj5ddhNFhgiLbZQFyTeeW2V
WHYpFvHBV7QYXyr23MAGdVjvwGtAdHux8mjQ+mZ7qgVoA07wx/DJtoSPZsKdagPx
q/TpuiSnFZ51avTYgWqAXhvnFzqgs/UZWm22UB/CYFdN0dkO1BfQAWASD1MjRZMO
VJUQAnq2fH3v19aR0XkalJslvrq+0T6Z436tj3NzthRwJ3uVmmLbm5r5nU8LVM7a
yqVmfitjw0IqZR2NkgCAE65o7SUK6XIGpDO6IktD+hb3XDy3HDzMJJYBw9LNALdS
o+ZHbWo3DI64bDStBLmQm6vZSAu/QejVlS7rqlln2c1KTrQ606va1fpp2O+0b98p
XE/CIP8m/qgps/Z1e3JB6lnEDVgLZDovznKvX4ZrWkiMeMT3uhufLJotHMif+PaQ
ZscSenN0uovrsZn0ETXH7UeAnUzAkf37wnoO2gWlbbhg0jdsO9NFFHA5K6XOkK9/
n838T9OmpcgJgoamYQ5zTMhw0o3O1kB+vjeTeXHra8oTuolXn9PLdikrjKZ3chWY
pf9oc5NDEgRdOBwZCm1PGMkh8KuPzpblLQxutMaWqzJwnLC3gDXeRB1TiIkiV5Ar
L02Wq3nmFcGUo0nUOdHIAMATZOeeeT1XbZtoswaKkEkTfnG2Duf38bFnXMm4SxN6
9tYswWhlmnHXSfcvXG2odLz2PRhz3+FD/SGCJ5CTyTwfkcyARfJXkMIqITZahau9
H2d85Owg2uvAYD6dCudWuNB21rWGy2oyGucXzqyOkULrPJq7k9Qpg4IOU5AI0TNR
9YPBu+xReccbehSYYXNUo11ToI4nutBH1hd07okG0cb4w1DWIzIPRQevqE2wyiYf
yXevQ3NIyHOWwCZwbGI1u6awIzcGVfCxV+xBtj3W6SGGbXxoy+ANXXQCU8pg7eEC
ysl8T6okVVzYO3nWZMMCsyFb9V9BpU0AHTypdTpkHLy/URr7gXGwOlrrSntLET5d
RQHP3mqTRIYoj4ju9JMK0DEDPz2PSPUKOe0aabLgxIICCbN355oOnCkbrJZsy5uE
fmnc2KEAHHeebHSjr3T2aYrzTFYroOwy1O4nLYs0KpAHvzS8opyIYqJfD5jH8KGY
VD2hXFfWic2O6FdrMluuHLYDJcWjh8zEf2RqoPiulFblLi815d33waCcq53L/fN4
RxdXoTl2J4qBh1xTJLwwZ/rc/NhlebnC933jUs1iCAMCfm6Q05FA4dzEoJ7PjUdi
2dkAd1Eqkyr6Jv2TIDu4QGHnwx/lOiQ76OSZ0iqH8mPaEhRzJLLHqCWmooi4D4hH
itMZ2YFrDNcWQpMctSR1oYS3wzQkXMwMj2Df7+udnVfd3CcBcx7RI/FYYaK7LK+l
ltA/KryO95YRCjf2ZlDtrJDKLL3pypmE13aQTtTUz50zLgw9uUK+U9yzW32PJ09h
2Nrs3lHBa27ue4q/iCKjmSZ4MqfFjGzPQEBShuxHBNUla/pYP+g31IIO4Q+e3ubN
Z+DVj8HBHfyYogeRBkTNoIHkxw31Tkn0JIJaVyGnk3OvzqUEdnOibxETvwyfg9tw
1dXyQpFUbfG+zWsQw02aDQqaptjubyRlfITNTUEduhqRzZ4y9hoU4mmnznLcm6iq
ptrl5V4rMb4/tLe1EP8y5diCKsYi2lakupzHuRrjXO5zX2nq69KyEUxa9QEvMg2C
IpaYuDYp5XWR7Fp0qe2puL09A/9UEahwtyWsIHlw/xJNDrfk5m0KEBwHA5it3mQA
26tTSfJW7dvN7QulR1M4F6L1r6nhgl/JJHgnejBq9tTc8T2JS4xti1XEScBBm4Qv
k9V3IFKqk3x0eBJT3PaZ4Im9Cfymzuoi5o/LbC9pPZQdANukfWiM8RkxPY45iFz/
YrsuWWQubWsO9uM2SNoHCcPeuBFHtCP9LUGs6xVby5iYZdLKZOLhhMSjzE+9S6Hb
TU42K1UwAYZXQYW8dtVvANXxHnVDn69dgUy3INFaNKhRv8YCCDiC5Ftc0hU/yApV
sckFCOWj2SaWrsUTRY6VTrHg2mm929Adm5jgEnP8qKUtiqUnjflOiGzBL0QoNgeG
+bEgCWebEmtB3W7c8s5gM3mCrOj3EPIkJW+cbzQzQEzCqGeBJd7NVUBWf8E3bcyg
V591LO53HjN/iHYblwzCKn3PVF096Wra1dFjPM4Qx5/5otauXACk8MAUjJdGzPg/
p0VcN/Wsv+vZ2+NQ3bYLeJUKnhUd3ofAdAfLAOadT7Disi83+dy3+vbudZqRbtuO
LtiBvOaacYYew3aecYpjJX8iklykMeJetQc/3+Nk/UFRwwlNbYS5F1g3W5rJdVGv
SRSdqpTKyzxIta5Mz7ZrxkhDph5CcC6Omz6pPt5JVnbTtfGAIuEHp4fOgpqTC1iF
GqMGNBcmSGgBaykByhoD+LH0+txA6P/jL7Wf+HHYsKqAVAVCl4syy/f2CGU9oA2z
P0Vme/AzyORgzPzNYv/cQ/kYLiPzYtz4F2vBOXmiHm4HAyB/WEFmh0IRPksnSQPw
0ZsDuBmZseVempod9QM+kxcYXeu7OYxh8qKXidZU7+03b8D9qAgfPQmrf65+RlJ+
nI3wm2vwo0UT+o4m0JcReTwV1jTOIJAxqBavOibAcC3tbYQo22JuD/aNB2gQ/4HR
t9E5BVNZ9LFAzB5zEIwiuMJLO3TqO9uE9McbDF+ghU1Njsr1elOfXqor8BV9AoDi
zBHYvEQ0k+FcRhaPzfkZ8c8YyzvRN9utPvwCoHLbE5yI+Of8+Gkz1UizARbThNzA
IqZJb/Nc/0EZH4bZwMNvcLqHxRmhe0PYKMDzs5r+FkPsuIVO5l6PTAMb81llItae
hY3u2ZZdjHjYJQihpJk85H1kVcU0eNY5U4EebbDW9UITZ/fHZlwEJcH8rCakUExg
FoqFuCKzS8wD44DHN7iz0QVVaQ1maLByi7Db+onPto5NhISRKDXP0zLF+3Vfn3fC
4E/GdHSjndTUf6HNL64DLsnCDv2TXLQTS2Oajp46Izq2ZWKhz9VCZPyBgNenPDJr
+UdxWdjRp71HSfxI52DUw359mkBK0PP3eGJe7xuH7M03cLf5GTT/a9XG6kxuemMk
RVwdUdqxtLnMbSQKV8xuSDcc3+etZWh639t5Hd0peCgjWh0tXASSNJ1HuJfr3Y5B
uDYtX2div2zwbAgIf8vqhv76YMU59TRriL9/H78I5bKMnbBXOJv4KCU9SuNND85z
Y2QlAVcu1vVq0KiwPUFFNE7uoeIaWieDyZ93ExCyPcTpubo0P7PWiZ7Hd+fbi7Uh
aFcTQzUc5YCm6EeyDmD8xRULPi4K120M5zl4gQJYuTazVuYu0jvSq6SvvcoLVwV5
g0IeZDoW+9MpIjimdqBKqRRpnsNZHf0LJgT+jvJIdFvMYgtGSLzl6H53siz7WMVs
X20QImbG0G2a3WWWTCp9vPCzhcYfRM6wMLgmRxxlSYlnVIl/X9RmFBL2G16+guSm
M5hABK78L5TMi8hMpAC5v44U5Y8cwNAL0zWiXfjTL5pIZodbD8nfZQk7FHCcRCxf
RvvuHDeN9XzYR94KkJGzb2mqbLRuDTcS/t5hVwcdKTTT8TuFrGND0MxdQFEK8C9q
Zho8569WENIAgizssNkeegnunH6a+bbBlbpjlNQJqu//01yHcM2ZO8zawuZbIBaS
ov2KWwg27N6LARp/10X458kVKC9iAVvY4QbdeRAbm22k2nX2bkkhV61XeTfzXFr/
XBEF/nQLkmb35PBQtxg2imw3NbyK+FDmrE50FaxFGLIaMSvpnldiSsn99TSNuRKz
J5kG/s8y8PG8N36qRN6AuVuj4DowbS8y3Nm1L3LXw9cMyeCUPnsU4L3jw6MpS5cB
GkycUrbxJ3nuIRwRewNb2kkpmnRDpt7KTvH18bbqaG9I4qKl/DHJddkHNxQuqMyw
+Ugc+GrEBx+PacoBeMdrusleQxbJRO/XwzcLu/4qQzDTHGwXbVR8T3cszvpyc8TS
eA6f9X1LVN7hwNciCqZQVFJGofSjyLR3Lg0X5KrUUdUb9NkzBViq//Jsfos0DL+S
YOGrMmW2PyZOpE+E71UoEnjYeDwYL+BmWk0wb0iiSRHu/2o0EX1NIlwcYLVM60s2
0x9LKTgxGbu8befHquQmR4DARvrsxOYQNK1xG0M0Wnb9Z8X3/CTl4W+fU7NtSsFf
0dD4Pvg6CH+2TVVQ6JWFSpV/7JXyf4EHtLE14f6xEcyM1iGlV3QG6bROoHnCDbXo
K19e6hleURgLo8XFiP/1jKTLHMR7SlDSmgMxZ7oAyHLh0wxfLZikf7/1pZVu5Oek
cZCwKGtgqeqxIX/K9o50f3TsJlWt18utJf8XEBgSk5HxsTyBSnsXzPF/psmb8xBY
837wpxGq4V0260DkA6V8XNiRoizJmkNg7+yPm+E7f/6ftvK5BdiPtvXnhQeV0Qyg
0PVaV+33PBKY0QeQ7gNjHo0Ab2SMlUjjAsHw6phzBv4iO3ieVeeHg2MWBhJaxa2A
83iz3WAydXCrjZ0O8NC9UXkFxUexagA1mpTVQLQDSBhGMNbBkAGwXEahkREKDJ6u
njRRDjKLrn2mBwCC/P+a7lBLXURXfQ07TogWG/nJto1UqECNkBDVG71MEZYb+QMZ
qemjO6TCHhstrLvrB85w5HmbXJQ7evMUnb/56VXG5HPOd1+0yDjTU4Iy9RY7bTz1
/HAgaPXAjkF0AMvMJui9Stl4KtyhVYitpfk2/J1m9IoeTDuXYoPt1qJu37YHx0t5
gCCq1NbU9zNgZ/t/vnmTbwrOIXquIv2u50agkOg9e3vw41puY/lOxAkGQVBrbLBH
fdVokDIeu4sMl5n9F4RM24KjpLO1QsRgpMBEVQuDkB8RnGoHAHrpVeCeYrPhA1uI
B4XQG/HIJ7JYW9LqSCdWM47SdX08trh7H/vSvXBM+8xyx47VatHwCe2vupG6+xSa
eQZXaE/4iyQh7PuKHdep8wSdaKCIKy41s4uppkzBdazMpk1KAldvnT+9IBitKRo7
9kPd14agZfz6QJUhqgFiPvovhXaS9VPZWJ5U5N3x33khZSnEwXInW7DCEMAmLFO2
wSwgnamCRATOKZFOOtMz1pGpmmJX1x1lBuynhwHj8h+ef5etk1i1QsT5hwnvKbg9
ekYnee6jIpXVWxymmkPqjip15o8bIaTnJC6XOnEl+j/zcOxzBoxxjQuHa2l9i2yS
Na0Af961+jDhwO9XQMCotqVW7QwtB2hZjlCZkHYubIljtGP2Ma8hCMPT5ADljbG2
jq6d4TrpP6QA7LGNJ8z4vGY84ZPwJWVUpVB6NU0PRyu3ExrNBZMRGpTxEeT8PP2F
IbHGDm+hMpv6mrC6cc4l0Wkn0MkkAKSgNlG10JG46DXyE02elvT91pPmEnB1bjK2
6oaph1TxC+ZRgHcbHMoSOzsz0ujCG5UAaqwFglgx60Bd9H0Y9+snR1ygwU/dOrWv
bb9Q+r3fvyswEdCAyU70o+lAmWIny9Z9zu+hYO9pTXHYE0zgvRrCknjQgJjbO+4S
xQtdCp2QFhO2ASMwVj6nxxmk9uWygdSTtSnmtYlusCjt69bJMFJvx2mR+5fSCPjx
evQwlIPbLmuTblVjw1N5DEgmxCxtzetOle18typTa7Va33iWx2XRqhSJbJLfocYd
QwlG5r+mW9CxS3AMB/QEUYXOblP/lE8kXJXg5Zx53L2bHBZbMiP8uGHAYAW0mrFH
9KW7vqL8BZOO3O6lXJLm25URsJ2uOFutM18E/2j/1p7XmAAgS7CHX2DjzD85gIHB
kXYNdgwIkfc3JXSauftV1Nwv+WGbyhJYsSoy2WYZbscyyPE5nhNKpHrAt5LazMuV
/vLW+BUgEgARtBhfIABJpovDpx7I6oCHh4NirwKCglukQNDN6ZRgKIsIoE8XXCaP
010H+xd4CArr9aZaOyYDJIOvA7LqqIbxulLR3kdeBVYdictouASKjtF8rAN21Kfm
d5RsEUnksdA8NfnuAyMsV1u1HRUfokmQewRAcN6lbbkWYHedh7fp7WlOsjROfcQ1
1LQrQpgsgdoG8rlIRvg/mo3/3g8MNTiJI4+NlRUjwSBm/exx1WUEjcDQpicbO667
W5LikRZ8oDgDv5+xgMxosU18Toe1pc9fUM3Z9Ch1wOh4HuZmgSl9ISKfJ16BtMYt
UJE9wZf4huizKINnHEcEftBTIviZlLx/xwHmoKBYF+hF13Bwy6rNKM8z0iZgm8lq
OS1LC3nHp+jF1XC4vhKoU1Bn+ZoAsBzbVJN0CpwFD/dJwMvG/7DvQEe6087Lylx0
WRiBM+tPBX3E2GLWAQ9N0NOg7tFjRJOYWglqw+lUpZQOP+jvOAkDtegeA2pWdKdp
dGxm6Ub6S9s9cOJbr0v4REhxjSMkVr1XXRExcF5NCBecp4Xk+v7LGYCG+8/SogfA
WkOEVA87ZJNq6gr+b3hfBFtGCs/gqzRoLMpkBE0fxmoiMGnc9IaQBPmV7ya+ndvl
jGMEnZCEBXBSMbEt2zw0y0v+eexibFrdhL9p6Q0nVKjzzsEsWaY+RBEUMhjEViyx
a7nYScjRhqSAmlN21kLCQXsKKcEVJ2U351C3vVgGeqNv926hSWwiMDL8aL5a6Vly
SOq7hiL8bVpTr/4u0/fMQ7BjqKv6q1STu4krZGa955wxaCCEZmpttEGpp+m3QuT1
MACVN7xxNUBtGDps1EpEyIn13ie/yCHLgSEIqcROtHxr5z0iFSs6VOnY0l2ENPMl
HtVGDlef8tmA0IArGLCxAoYvfvnP1p0kg/k45cSxyCsi7IRN78a/znEMwbWpzrcO
9MLf9gEQiFHDv7EVnAyIP29e2PlxHzKXaoYXF215cB/rIqE3ZWtGgtkDOgPWGLdc
Yc25AvsRvDUACQsblIIn46TMHvYcgtROcSpdleOffmP+6uRkKzWDgSYwR89GuikT
E+HFuoGflMUOaRkQ9ENPnHkfDP/3KEjX90vapFMXoy5APP+de+LlaKQgR9OWlUx5
4wiyajqimr32UZI8XePEnK+DODmz8iIGG/6hR170k362+DifUQYJ6rIm3vuBzW8L
oef/iwbcA+QbOLZ/zDgRh/KjhHs4zDc2ma+L0vDyNVOF0B4LQIcC+BP48myJRbQx
QDW5/vWFhHalIIKMswVYWnrAfozvl1XqhTTXKrYUn8kCf2HKLnnmNWoPtrztc7go
zpjzbSekQNDhc9vxg9V870cweVzfJaYCawc8dS+ZRBSmHTZYqjwoolCmzz4Dn/2Z
tozju6tgQkz5o8yvMKJHiUI2kZah99LMKp7hWpWnHgHEpXVkVl12C/dkDDVizh9r
CjSwmnJfoDoWO1xPVO2d3RZa+ZS2qMDI8YuaoJPkrAsTsLWymZ6gVh+eGrnkJLEh
pjXYpVOL8bAIQcG8FDfEOG/AX2RgzLhjrbemiiiKuDvZj0Sf3Qicm0+Tu/lRuK6O
mLAWxKAZoNYad7XIk/D0ERYEq3msn5LCP8o3a+W5uxi6vvbnCkG4Z4KSzNmXKG8K
1x9XuI6A8AMK7b9yPujnzhCmNbimMk8uOVZ0SPAJWGWNR4OsgAAJH1KZdkYLodrY
zLWSfFeAkSahBBLVrwxAE/71FXkJctvCzYoBHqufW79PtgVjFpTVRH3+Hh6Fb+b4
CjWeDNfSqvcCUjKymKneY3TrTNawyr04pMtN1zF/K5IhX1BbWhO7/Yji0Nam+h/E
fVx+hWFLm7BbucDX0fGVuLRSONMxU4FYp5CMHVJNNh3ZFjA/xC9MdsPmey3C2KZ/
kzzE3hAaD7tHGt1nP1iHlkPLTblvFYTIRLQr8zMBMWce9X9K6bTWfx9BIqXMD9Xl
8DCfWN6v5aCoHDU80wHyjE8w1FljOrCmEq06XP28mp+3losnTADpzIsN19LIMg3h
AhmwqpqH2/c0fmyCkPvde5QDUMmca0gygf7XuWb7+eAOLnFKccUhP9z/xrM3v8lf
v7iC2KgBb1b0ng5Wx9xbfUq3RIsTyZvqfyTU80VhEtMsJclxpNhXz0HwJrt0neg1
PBgigXaJOWOp2PvKBWhnMbUdO9uF5oAKKkcwCBvADXXZprAlfDgJxw9MpX4xD+qX
XbUtiLrP+w+Zk1+kFOB+erqFm0mRJ11gr8w81FuA972LoJP5a5o0ep4t8iTiFaXn
llWFOCyJY4rkM7/AmA9IXnsq5sN0WcU/OxaGeEWqFxC+szTKfvJqhn0+fBp1r0us
Y3IweTg5P++qLHEwFAu1ihLZ6SHiFpUw5j7akKaLveufX5JjFm2cpUNOXgSA8ULh
0ai3/BarJVAkg9/d89aSrkmuxOyK3lBasmhwr3C6t6PAV1Cfv+l16JW3oFxam5Wb
ej47JOZxQ/uPR+RHzJKs5IAEgZDYTckbG/IN7iMP2B0L/3mtwODVo033rx+rzqQO
fB51+iZpdYNuC487FtA3pnlPxklFQ3zs7WVv9luuMDL27kiFQXw+p+mK0nlYbvnC
7p5RD1MVX1+AgMhSeeFZMrbd2rBPiugwGQlYRUyaTNlsbpaXg3DAi2C/ZGmAKy8n
u66+jXxgonGIUHQ4PxX6qyzZCRO25zqK9AikcMYprV+iXcKwuvksJdqf5y8QwaBT
Gyerp3KuiSGRD9cZZg/NATt2wH1uDote8i9AGGLGkbFIPdSL7sEVrU2Tvdk3OOUy
yM1rwQ/pOCiWle62/5zJWGuWC6ej6KjQOyjLJ1rSt/IlQTvgddK1egQxRf+wgc4l
CIucTKZZ354mZUZSQ0+UnvCY6GWIGwwurqqYY5AgkUv6Ei5FuNsXE1YDq2J3ohSa
MzxHXtpy7keVurDFmDQCmfm+f4Pf9oLuHS6u95ZizIbYMCPleVavxwCL03arNTlZ
xOrmoBT3Nd9CWSpj+Wqgjkk+NGiiY6G8DoRuTsZAfO1l2a2TGuoD9KXnK1tPahGG
UB7yAtLgqDtkK4kKvxiFg8ensEQ3EaoLhGm86p93su+0V/NGXgBzLr8QEcVGXPuO
gvC292khkH0oSmsyA/3vYlI/ZWI6l+UnWudY6wVborzAcH60sPvWseqiD2nfT50d
8N20Ikg5HdSgzHj8EpUTu5AIILWgVq6cGPY4T+xnR9TvfdDyyfCjY+bdHWkCkU0V
0expll1Bhog+ZaflpZZI4t+nS3fiT0kVBRB4dGsvNvjruujfOFWn3YJP/z2oe8dT
8Xds5rabYGjVWIrM482HJi41FRA72n5yxmAa9Fp+GOAC5zW3ZYAi1k8Z7NYM+QWE
FyPvE0Fd4Vat11pwzj6k6siKhPJei/z6fQRNHZzqxKr6BifMpDsbZbE6KnCqI9R/
fp4aM/qpzoUl4jHNwVAIDw9MdbMHr7M5B02htfaymxw0XKiKjE2n1XH0pQo6l4y5
AP6DfNQUPGFlKaBFCiB5l8Kuax3IPOqPoBZVbgV5yuEQ0R6YkpeM4c1sI2Sfk2Qc
ff5CtzuRnT4Bs+s5DDpI9eT/ABVKf9REHoFD+Dl2fjHUMknCY02y6ymMHsh0sO/7
jD9879DwQXasI2oxV8Wpqgx06Q8y1D6C9sMtXhHBHaHQsPLsZfIKzs6PnoQk1/hL
wyRRDhT0eGM2DTgSVfP6zztQRRcIwbxVReiCoQrdgwS4uNiTb4+YSzDxDdOwt8UN
O2jVv+mWKbrLN36hx3pdduVcfFIYxmvDf7s23hBlHTCTBiF/Iok8TGF6vK2BdwAl
BYGeLq15c44G2NymVuGiBemFptM8Vit8r8diwrTEjkcJuskMBszjdbbf2vFMoE57
qywGBPQh29l34VoTR02ucax7f71+CteTme2EgZLQNkDfyjNBuDsMyh7/D9yqZoJU
bXCGHOS61SdzeTxbnv8Ih0Va3HiROnMeqFlgBp+rznyVTDiRQF2BCAgWXOaF8pg8
/5l24fSvosfp7V836cYHP8uLEwWQT7DSOPFdZt1LFayh3DfA1tzPViwQ95HRulTS
ZsQ/o5Vf+bU4qODNtjK6lcKVc7DK8Biev8ocG7u7cMgCh6MPDekaJSKYH70MmUtk
Iu22Wz4DKmcR6NTM+YFd274Nqb9yh0lQxblQo6lsxoDnXK+I43vjDay6M1mVeDiI
SGL6NRNPfzgQPSDyhedA/gJxLO7q62ubCvDA82GWpgPRES86Hru0/626eZFf9/Fu
hwwgPr4hrc2sdiR3oUwzgXnPkXeNUZ6UkoIHDTTmpvUDi04nyRX1QQbjC4Ejq7Eb
SPdOGuI2pYIEw22y+Yu62O+qzura6Z87fmrrouHGr8y5StlaqUnYZMrnjvU9NMXo
TIVGRgIMFMDGoBa7BTFdzzU7olTg6aJBfK1qZT0Wsm2A3hYT9GbNRwr/mZVMCGyw
reSE870g+h/WPQWfYgUa5D/lZBglQIm8kT+roKsvBDoT2bHPVWjSNkyhlD8aF05M
JJ4IbAJX8r7ExuS8hJVq/q5eP9smiyjM1wCyRSsukWgrRt1mVXHB8sC/AJbgtT/U
fUjIoD/1HpjEQZtAe7KWUHWp8NquOCLqAFbvXeB/MGSSjzuMgg5zDaP8cqr3pyC4
jwwh64QNu6OkZj6AfMUYH8VBJOqvwxXq5Yhm8MDGKKRJs5DHsb0DECjNrd1RbUF2
i7YmtlBjXgFohi8nriAKqCyeiLnEBk8eKJLgqXorI2Rlpw6FTNDInbnZPxzDQhXN
MLVcXjU5El1BS1jbCx2SYu5k03x7yWJFcMs2Nq4kZpEO8f+DSOP8PmKheor2qNuc
MTyo+Vf9SVpih1p7fxryyAPItHx9MzAJjLcDBGl7hNkS4tAeFZEptPV5Lf0jyh4G
ixn4Z8qFyWsp8TJoXnopezEijHWiAOQ/naAiC2nfEqVYDci0DCRVhVmUGKhLX2W7
Fs9YVCzrizUorhs9ZfEHYBoCpMwrt9BC9gWtBfbw1BmoXNGUKgTONy1lTjGfySMl
Zeh1OvldUmjYrZVyLTgUgqU7kkIWnyFBwru4BpxbNfJ8pZlaPKx/d/ptBKjDyqXq
wddDcqq80GZsXfTuo679bkkXbjXy7B84QMZ3WfSx6JN3vM14LlYzozPxmEZanVp3
KRBuxqiEUeW25QwyrXgWci/mUTctX1tW1oAukgiSkkbnHe3jXUOeHsm1ScM4IrQV
hKaQI3L1CgWJ1DMfE+3WbMsj3L0MpsMvKZH/ahAFoaykOB+xnlLWBCo5OJ7m5wdG
Y2wnxxtdDnub5R4tBJ1lZ8ym5SuS+9y4Y+m9on5uKKeR1Jzsw+9P10CNXzFFAeEG
g+7w1ploxRE4A87WrhsmxWtQQguLyyQ/7q1yUyuak6D3ZSncc16M9zqR+PaWuVo4
1BMSYjmv10YGb/OSMjYYEz5LeRxRLeqQSjBwkiq9syo0Oc4V1BLDQ9sGlREKNMNK
ALD0JKBCKJqJP9DoY/fpKq96GCmCoIXX5DngCRDNDke8kfxiFuXhWG4j76g8w1Ov
uUr2KgBuF/5Fyh2CJ6yYLV2+GUTNmFkDTAttLIY13Gf35bi1ionJXBbTqQ7pooCs
QElhZu0JcJy4ZmWP/+2zH91oPrxEEMTiA/bhcVJQt3jJ9JHGLbiSwkATnujbUp3b
SGs3o1VYv4jvl2ippmx4nbXRd0z2x0/SUVPZZJMOIrlSMM9Ts2kIJtMMgrCi1zrR
Wz7yNs4jv2YJw0PRwNzbnzPYZQr9tuhgE9fFDwlJhHk1qkyaLn+sL622VZRGm2l6
/NXda2Xrb/UBoMHjyoAvjfKkOAtbyyAVKsKztLcs7fg9wJTlqYZXQPBwYtOpxjYb
bymI2/8lYSp7XOzr8Pnv6B9KzbF+iUsM4QWaFv/U5uNpfCRZKrlGF5yAQ4wjlUIh
ZVxElXtMnRIyI/yWYul6osjUILpzwUb+yYUp3rVaLF7o4Ep5HviHOGxRcvoC630u
YqEdVV9T9uBKCrHoEkI1bJ5h/0VaL+XKhOHYXu+pHdrEot9dVtMZE8o47Vcw/fgi
06RM3HSoeh4zQHAgeNhTEctyaNkHEEaNT4zL3NXq5hW9isq9JtBIn7vbwg9yvzFD
nAyGvHDo2uHA7pMAgKef8Yv9CGFTo4GHILy/TOxABM4xYO9aVlYbPOJYKmFFgs+4
Ikg4WnMFIagbxYxc+lKMNGW+FNafdniVUSmxVfHGcCCq7WeTZAeFAs5Yir3aKnWI
581uxmMsi+NVqZkBoKnXO6Pqo65638CmmxmHR6D+SkOu9IEDgVlMdLP7OflSNYto
3AnbkZoqOas2T8+xSFyWgzFY9S4LA+1hnmxcQnEdgNDSwPwqWhbj9wMBmlW8tUNS
rLFQToJ5edTynM2G2uC1gcGKXF7C0zGqEXcW2IpDuv+EbC3w+RojFfNIYRah7pkb
3HkchCUO84cduNy6/rEdTkJR72L1u+GjBE5u/XfQbXk7zND48nEeN9y+nt7pGIzd
5Vf3wNbT+O03OoXtQ48jgSFCoeT6v3qmsR7iMei/QIw+BzpO4cetJ/0Om5cW9AMJ
QNc9XHUK5knXPOlBfPD/HJlqyh9XPd6osw7gnP8oPL7kjUQboppCgf0llfFx74XG
Wd+ICjS1dCrHEyYfOhgUCCmnNrmypcb/hH7hn6UeT6VrZIbP42nAq7zcTi6RebC0
U6l6lJQnPZXeToJkPHDleBCT/Sz+GCs8aNm6+33877WH6Sry3VsQIXyQaCZpS1Lv
2SS4UmVZSNLChbIUUie0MF2UiKC8unR7aZ6uOTEFiidhAC7VE2jKjuvXo66RpYYs
Clo+oQWR4lDMbNPOWMLTgrMAYAiObHc8/SkzamXhdmgVo/cW0bgRfbqvQcHIML0I
InXgNXRYdCu79rgDYp89Ze+zsaCPlMaXGLy6eHowN+TvPFFECI5SJLB1co5dxO47
/dBD/Y2hBYyq8xn+zP3WUhRhOz/S7pm/iKdIqfdP97DraToUY9tMXGdRzAMFtznx
TCea/d/pLpUzC24HZ6AfwPS3T9h5la5MNY7s0KT6NOi4YL7gHjXEkRk9nxyRhQQH
LrpttgR1dBfGCvn+MkKYSXODxXvsnKoH/DZ0pu2MRgcdevlZ7/+OjVrfLF0C73jY
R+2bNFp3+TIamKq85oO3R9/Toi3takD+EFJXxl6A7s/AmyMUEhj45w+Bhpy6L8J1
JmTJTLZWrX0R6Qd+CGYlvEKv4u0EWForhRs6FBPvHWqCaMxVdKf4bvboP86sR4IT
X8aJwa0WM1PspkkGF/Fa9PjcIo11Myu+woCu5gvdpoW1lLGHp+rmI9aQ0nxPvs5F
EUwz2bMTbwSeDYQlvRexiRnc8PXXZCTdbFxwDMhDJOgWaBPvaYUvYPqQPbscjRbW
esTtlv6+l45bF2e7K75/zoTDCpFvqPlnSgYn+Xl+q7Kj1uxEQ67IfeVyjv67AgL4
QZxOTl42woEBUqwe8lUI1C+C1e2AvcGEJ8Dcgbvy7f/WbgRAtx0Y/zv5m5aNH+pQ
N1DdTW5/9+YqNr3ccyxr10iI1nL5eO8x1FinmwYe90gd0h622CA7jzLkemE6aOMw
vFHbab9yMeQ+OkUZAzex8y9LERmo/BSmPj4V5s+ZF76l0G7vFnYb2QM5mBVpnUyw
n+k1Tja68uVJkD1XHb351kS1p0uouheUWQknl2U/rz+1FzY8B9tp5EL4P/JpN2mD
NPyeoLLywbPo0jZ/5inetmqalYQ+cAgdrqFWdB2wCJ288Gr88UUGbDxhNnYRX+ey
lFpUITdZ9F9ZWCY4llUPfZYmgNrrVFygXUAbSnpbKKuDAM14PwZR6WOmHssAnsUB
SdL8i5/vCz9yyApxyXYwH1O5mmhHtLr2IZtOkSzQSgFuMgL4QdvKeFSE0W5AM4rP
PjME0JjFz8+0yz3+7hj50zVkchd9K6HIr5J0d+ZaupOF/qL7h0rIIQ5TW1KQnZ2a
RS4JJBE2+y7Oo3B01/0sqZSm8gfwNxdjMHWjdRTRyqdIQGM+X9CeowrB6r+2iJaP
qtSwZipF6KYpEuSRfCTua+hZCdWRg7iKCPeG3Pfse1XQeMJgKK80DeFtQnOTgM4t
C9fTrVrU7h3MUf71ZjnCrnIb2BGKh/tBvY6mgjb+mjjl3xn7hk5J5BZAGgfj76R2
wqDz96tKOhxmVol9jMFIr3mIygJfYENOjNISuO21QDpo5ukEPaDgObi7fXYrm3sh
IDf8Pmm3aSlnWOO02l8UL1zlup9S1ghTrrVfAxjil49xRisT//fds22+42VSE2K/
AYCVUDlWtIgQHiJSSfS6Quxe79bFObBmwWQKPpUCMiLH7bTCVTUdkRYrzBzeNDBA
9c2LYy3B32kolsh2koqVQ5JIjappPMOTOGg3E635FjiNTogHLZ+2k9o/7+SB8tJb
I8W9gkWXdIVUijj61taaDoUgzNwwBgi4EMGWZjmWKuCNex128KbR7NyN+5FQssMt
YOwSEPd8DufElO/0bRHIoyRLEu8MVbfH/nPfqdNqtbIDQdeYkFWTmoE9755gM0W8
3F5AegbSBh4msO1Lb2HXVx/9jRUf40L+komVNEJ46PRT1jakJdnYJzhvfTbyPUJO
DGLo+A8W8X5HlLNi4NXoAYrzC0RyoXVWNlyGXI9QBeH5V82L8jV+wQgmrrDXa/wg
BcZ7/pV+zsSAmC/mPjK2kbJ4plAa3zTr8RMJdrZIXA77QztZY1pGLZ1B4kvbdAGf
uYDCgQ1YES0Ms5J/+o4iPiwSJmWUiiTu22ylHCFcBhQgj/G75x7BoHFUqHm8idAd
cmeiR/Ayk0Ke0dr5bZ3kfWncVs1pqdg11OPb5OMvj9KXxOsBZcnRcWUX2fItNw/2
vVr+byp8grcTPJuabSZKAYAlC2r4D/a+eNCjfxqb+GAab1CN38SBzTGgWCMPxrAZ
tpvgR0KrRiVYFBQK3BVk4LR5PCKFHpG4bd5d73aSsOGuky7puQHpRXePV+HVR/cw
jzEu+hOJDfa5I6K+SkCSwnulqrMZUV8S+Es2C7ugJM9+zcUpgM8fUSwKnTV2mO6V
wKsMtOrfEcFQmwwD8Perfzmn4dSYrFjeQWdPV887qOushq8cselSGdw63Xt+Z5qr
1/edeNEmkf5XjqfX4C7h/EFuuCEE3P67sEPrIBAEcgOamFA3aZ424WB24FavC+Jw
TfZmHFypGvKXAXPJ9TkBLRHxRzTVfosy/rEa80AH1l2SpRAclq0Ak0lmJTzivg3o
z+f/uUXGfFn03Mv1PafPiNsoORXTOVj4MBvfiOMnWl18F/B5l3dMbGLs32srPzWH
knd0LzhXoZbO4iXxxJf+wI5UudDctWEqtcFGryz7z6SJhvLUu1kRRW+J/vBCK3KL
7wAiJp2Z+V4lIvepbflAZKsTSZ5VDlcQw3LXzmUJ51a+jhAmVIW9DIvIEsJSpreg
Xhq5DATk/U6zLAo5QfgmSGAhm8oLL2t4ZRAVGIz2SR4jXzb79i+WogbjhhNylhWR
ZKrjCTqjH6USDx5ASENRLR+cA8rdRqVRbvf3wCmyqz+yIPjsgkhrxj+ui5PKqJ5t
tb3bnZEV35aQbXzRclEU0MjDbf9G0CwaY/PBCRDJB/oZY9+M21Sz0p4uSymOxqjT
v9v0GsOyRuPrwMRnE32J5mqFEIwjijWIAt/vvWyrQ/v3a+/OGLqInhQEzepxxb4n
NQ9WpW6PFaNfDVjTUfowlVl1zWimHNhHwGbUKc9U3tC+/N8TyAccaUFIR9yWwqb2
szbpzqSNy58LqiMVXvFrftDaLHkx0ke5GN+uVhRspaNeH7EC9MlSRFlnNhUvX5hb
FkbTsKDfdl3SiHsmfVT9PNU+sIaeLgvkxDxLZGAKReq2cavznrleMu3SyAjUmOSR
gTQnM53AJiCjI+cV5MyKxzeLHkmyJVPEtLtsxrrY5mLXDlZ521T5djD/5UdWxLFl
Zah6B+h+TNPo1jKx+U0MCe36sO35mrA8t1WlWwvYP9InwEUf37z5RtF9hIfm7o7N
S1LbQ4do0qCbCIJJAErWDGXoowGpg5INt12SPQhK+A+X7zPhfmPZP7dWnVHxEKsm
SNiI9zWBIvazhONljnRvOga6CvcLbEhtK6Ojrq9MdSYpbgbAnA4DaFfOmf3Yazgl
Ios72P5ZQAW0HmihYcZySrYlVMHaXc1tNbthEW0spAu+CT9fx4dLmAhOizQbw9sN
wGuz3391fc99wf4aGqLFU9fjrco7cGbwQ6XbXX2nBbi0zd72Ut2fzD9+s6B/GOPb
npZS6VVJc1BRnuyP59jk+NJ3f1bf9Zrw8/JM0+q720Tf0hBYo9wqHy8zUr1sOmdX
QNW9OVm9AZxN8VRB1p7SD5iLM9GWKFWC/o35S4ODOXqh2RJPfgdYl01egzxgcZBN
1b6YiA/ufU7pQGNU5vrGuvYpHrEMAmGcpTJvMRYUYSim+mx6W67zmH6Yh0gId15H
WfJBFIYPN21v+Er0n+genQvfkx8xH0ip9EzOVRFE+31aonNo2GOnf7JSX8kiRVZl
HdUjHPT8AQIDF8aZO6GuF3pXi/Hzk6sEeB9ud7lrdNhht2EcUs/ZhYwbIr8hoUmT
0vxerNk3SqB5YDYU1NO2xbzGFn1fuI6tXdtSQEHBpD2pw49lq/pOJUG4VF+2tMEg
QTCdhJrDWGpQ+BCsxudo1F9PL2vb3eWTw1lrYCzcpockMD8MhETbPZTMsIGPEhtY
V6qc38Mi7UrS3wXuTO1q4zDA4TyndQUtuY3o2oNiLLMV4uaPfU88w3Ls5xx9i6Dz
tIl9Dl/spZOffwUoNqrEMlG0+3rrRaMrsid4YnzkrU8IKbuWbTgsNC1VEN0i1AyI
6upD5KRTNgieEkWzNn1ZaHqul3UM77LjuijmVPihZuafrd8pM6jkOIoPge6AH2U8
j8uoXY6HazxgU/+42gxgKI6kIqhsSwwq6B/CIhg09SkH7IJEtMMNguCR+/cJuggX
eyyDz+OkneIuMm+rHPj2FoBd0OUiGQNVUhHTpESfKoTWusoooF/FEtPSfsv+istn
2KklSf5BxWoTV6onwc2tkB+IFhxoPYgMp8c+g/P3prMxELTo0lwG3VMBSLorhWWA
3CQ8/JHbU/1hgXuG1hCDN5EkMx5vF/L64ly6VFaWgEVZfrg/piahPlb4qOZ1ELo2
rKdSSoU+KOq5vijmS4uq6CFjjP9LImVtZUrsMnohS+JL3g9uv0ZGU7gnBRvGWgjq
S00/EXe5MohpZopAmjAAQ+OToUIGkHbRlGJrPDStL4C+HX1tIpVYCvO33hejrtrs
1P1iVm3gwAAILUyMkAA1V4J+yx8JQj/61DApauc4c7uffvRsXr+sweKj0gvB98ap
IqTnBgTiHIRRVDnbVlvjgg48uh7VhnyvTxwz0RjgwGO3MWjL2P/lp1uQdSfEso2e
gmjIZqdxuVICxt7LxN5VBvsoL8sqWda67e7pJBWvJt2D8x21HlDbTfVd1YctVGhE
yOZtUop2c4b5DnY1fS9DlCS9hitDqZ5fhFzOvPyAqQpGRvcrStYa0awH24bIS9MF
USeAghdVcUAIbIxAihKAC1c15RVg6SXT7ehvMqKgZkVI7V8ljpXNzRRzu9AzNqQP
Ral65mrmiZG+x/K3az6op4jeNQG7LFVWaJDEyCvbpBYur4qIOX+HYq/y6Wodk4AZ
roTlWCSXSACBIuA9sVsma4Qgq03ia9PrQKfdutrOhjbnqSQ6laghDsmegbus5ket
L3DMtuyc2iilnark/k8Z5vceB3UiSoN4KLi8V8tO06m0kTgIvDL2NkIOa/XHHqk8
d/tBNrDKbf8ho7vm+GnQ0bCAziT2jDm2drZIBUu8EiSMaUT539t4kjGAfZ17TrwW
AAQINKIGa/Bq8GGFUUNb6vmae1WMilWDVDGXgV5D6/AEbFqvl+wbUHNygYBvZNVK
jdcuZIwH57xJhTaXchjk1izLIUQuG86K2YVQEij4Wz352ggAGRRzfaTgj8mgKUZi
2FyKpzpTfJRopf+LSfjt7zQma69Wa1LVDA4sY02R1sSdCOVyo2ZabvYGwIipkrSj
dNXqtyJu8f/rsEf8I7o76VIpFj1GYjPHZx2SUhgpCTBgdmGS7bO47VeVecIrgzFI
Uv5y684+rtbW4oagMxAkoZJlxo2L5QllAp3Zar3UFJhoBaQPf+/uEfiUYA8d8/e4
kbFPaA7oR9oER6vLxIlAHcbuNRza7ILPpd0qdOpOY3jAN/bJoyrmK/qxhSDfIy1J
pBQosd92l623zmznSbmiP5tYe0WX6jCKPEuX+oP2ZxAp74ElF7lKUc1pNbEgMihA
bGQLO7DN7aWkhlwCe2vBlz0PIVZLlu5PUjKwIbR8xBtJxA1xCkZEmggPgNfYC3v+
3MWWKsFoEXSbi9xnRTA4VM2XXQ8JD0dyNKye1oUmRiVwo7MxUSzH/BPw/tBwKap6
vl5c0UwsFEYj/oJK5Q/PCx23GkGFfPpy9QD9JfhkYrogG572Tq2a2EqEwpwUhaPG
InTXYKXwFSri+N4GJoLCuY92+ri2E/P0p64BDMILx6mmxZYqR8IaE8s7BBWzjIww
VBTZ3Kyovo6PKl3lMrq+dMSklW91lefdJuxakEFbMEeux3Y+mHa0teje6m4NqXHD
GxfNg/ZkXKd8N2k8iBKMfC/4VljUfO5cSXWLK9MQJ0KHnU6GHB0HP4FFqn46hOxy
pLoRCCWnb1kCwZ8crN9f74W0giacTqKlCO+LqUiYpA6mg6YV+jzSkOoOKJINnsWk
MCdjh/zi3tGqgnuYeWy0nwTUyG5TDdc+6nt0kQjMLdnu+PWsABCj7y9hvwsgkHMf
wcGa4pcm+Rrlqb6OK0JZP4PlKe2ylyzL9nWhY1eNBx92lQWmruDwD/vRjQicP9ft
+r/KiXvYrvQMIWxtej85rgkH0uLrhIgHTbL+4BU7dZCUPjJ8Jw/RiY5L2ekr4I0/
xaGz5E7Kf23LywSZoPxoUlnpPvYY/uxjWFBjiXUZ5shI0UgNT1Z2jpnI0W5cWGVh
c3NgcPK7G+7qLJPnHr3avFDkFhoXbtuD1YW15d0sdUjxUEnQwgd6K15+Qt35pyAk
QTwrT0Lk+QWTXz7aaxl6WDd2qADf+f5Z9Tj2NUue1sOvIBkTzSxAIZBft2Tr92LA
jsupeWszhBavH9cQmCvyjaPvebsAeQKMhcOQ9VrVnIpPPjKgzAW0hRPxU010Ch+G
qpTUIcIe0pHThahU3ERXa5ESamUbxATx1OWPUNt0XYcDjQ98ujVAQnjQL4G6Yiti
uDz9NmOsvR4ktF4UOiSyu8OkkdIUp7VbDL21/R98SduSti9O/BMwpbT9MrW16B/4
8/iVzTI6urx4YcKh4Z1eTYZ7q/VAYnbGvHjS8RmNrXHQteL2O6ySqtHqUN50Deu1
A6AKN/APf3IFKy892vvyV44qWphpSPJ42qoBEcn/CqhUkRrgECDWZX9Ly4HhtsIT
11747622khPP9rNj29icvt39z0YVnshYZjZUCprFRro/9Y3mXHKXNNtp7MsnILma
P3v4oajUfb2lVyBamlEABBNPP2XdgBXV880uPbaj8BarRy+dDneosJP6kgqweCWq
ALXvo+bmL8190QFm8QjyZToi2thL/s4rtqKnniolb96z7M5gbRN+V4d3VORagHra
TsZlhwUn6NP6AvBpDRPKLC0htvQ6HpUp8TH9jIbCKDfBElTzNicdouLDhuPI6Nju
KQj1ZTdOLVLrZf5+rdOtTnkI0x1QVKBurGAPGu++8kEOUoVgYsQwsSpPiTm/YhGk
kkqyrFXC7L7T/WZC0WJKuGnikDcmJzGsFOpmzHsYCM+A6x68sofL0fu9dzrOM4tq
wL5T+am9kty0Ap400Xrw5LhBW8pHS/dKg0KeKs2Hj5LL8cdAWd7igb5gvyHiV2Lz
HyJNobKVDa4hJZiRU+vxvnVyjPIHtUO+EYje8M3VvARwnn63m2fUt/eTJYVoJG3y
DaYf5+4ONHCww4Puf9dW594BOIrAMl2sWAvB/QHB+a+44ISMeYppKTeNSxc+2nxt
4lpqC0Lza9Pl5YrXhX59Wh8hIzPZVRhsSPNDt1vYrpFAOpIOaKlz61CQmycy2/Nn
sBy/l2OxdnUcktnlCsxkdEmDZ/gAvXmfSuTSsADn+aVHKfXXKkktoCIejlrpm16c
IHIe3rDWvXDZAiGgyD8Ht/XT3IIabeZJmDzGPSiQohpvSWTL8/2Dk9RzlwTdHxyR
lwTblqdFLht8dL75JOUYTSvJM7Q05izOXLylxdQd7Iz8RT2asGGC9F/IrcZ4zZ8e
0miRm50cGooAWkixpZZtI5S6UXGAX7cNO8SE+lpH7601aclSFdeAnRniiYCxS5T/
aiz0KpWDYndHIt9uX8U8wHNHuCHOsY+3u9hsK0v/9J4=
--pragma protect end_data_block
--pragma protect digest_block
0VGn3PYPF4TJOQ0KFFMSD1sA13w=
--pragma protect end_digest_block
--pragma protect end_protected
