-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
JODtHgykZIhpPV5lXQ7rKZb6ev1L+M/rhs9oEIhCHllsXPtZcrdhnw7GbHioqH0S
MrZKferIXtIAa7Mf1jhhkil8i/FfYxnKjjQirEFWixutkWAhKE8rJdhXnbUNti1i
4aio+OiE9L72AS5AkLJaYnd5Q38iv7SB9zUO+acuqTU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1680)
`protect data_block
bwF9PlXrnUSorpipSZQZvmQy966IiBshEV3ShLv8GPSyt9ysIIxlBAo3p8DL+Hum
rOWEWm8PBYbyCcmGe+6Ux/sk72AXTXDM1cu2jq9nd01ZMxzL9o2q+da79sN+Bvat
Sg7jBK28YwbYzJNplQdqSr3cg7v0YnH/B4OAQY+lhn2IQr8CDpPl1I/K2JpjkLBm
sM0DbzgpkvhlmgLblCBTtzDsT/w3M8h2Ilgdj/qOy0hr4Bv4dODvQaTQUoWWX0+e
Q4orz63rQTPxMqpz6RA9Mflcos5TBnJcJdFAHnYGMIMUhKPkKquBj+L6IlcqTSD7
5XxmwYZapmSk8E8birpTn/UBLKqj8/1AhOUAO6XEN2i0+lqNXwHsVcvdGi5rnJEL
iBsMg6Vc069K3PtnUUjDUH8bExK/7Wu/LgBs0SJQ8ByJaAui7wtCm9MmVFzSIkMp
dbqBWCNsG00oBwZksg+QSOZ54yqxVpdZf1UMVg9TS6ySPbPEtRX7aoqNa/s8mKLg
WCkm0ETxS08iY+Xe7yg4rHT5RJ9TMbmwPeRMwQEAhRGnZrOsynUps+m6iKC6t/Zu
VkELr8AoEBPBIOLO3YPKyd00ayMtAdEb4MAUPeYiharN/XV7jdQFu09kjcpSUsJQ
PDoj30fEltFl+rzi76KSfDqgG3JUXOU0lKdclcOUwsysE513/jmiGyyqYlUgLXar
NdZU3WEp+5lPDYbHy+3GfjeBZeQ3bOdCH43jh8VAAcT35vWqB/aQJ99CLwW5Z5OR
UX0TbN4XZouXuWRDiBCHdYp0SG+cjfpZ91vwa8s1SMNuEFrEVhqon4IqiyLVpcrE
XfAJQxCTUttv5A+OwbfaI0tF4HaSVARKzjOQ6Kv1CxSRVMaB5IsNKsvjX4bM++xD
FBYCtVHNyj84VK1yDfSPsXnoHZ4c7MSYr4uAF7UtRTq2OdGciedu6cB7alH2kplp
fKV0Lcy+n6H9ORhDgsT10yBXCHoDvYyu9D6XLjmTDIzRsH6TTRzyJ3PPUgnPvzY2
Cjc7RpxK/7+PQJNJeyKyrwZvAhbg50nFqd7pRb/pt5ORmshSntXgRxKgdYnW28WN
tYPYTH67qFgjfzcaGNfPDVtkeCOXO+jP9p2edyIDvc8raRCCMpR7kw1US1Am8MXv
zpcweIWv5gxQ0dhaN8S1JZ/2UAMxDhMQDkxwShKTBv9GtpYazmCOKUy+af+icTBM
dsJoe8oe8aLwBohgnxuvXxkFOtxsebSWc0uSXRrh+eIcCHzRVlrE18lLotP/TFE7
y9LkC78GTyZYnB4crBiqGhywC5KkNJmflKIp7UubNsh4Kx/kBA/qpHuD6VEj9XT9
tMPR97sq8s9e4oSU8yxhxQioyPXXPLsbnB6RYT9d0hUaRacIVJaFCn32CuKmEz5u
OtTgbjfKCc8cVT5yyjUMhvO0DSCQ1N1B4Xvuf1Vxiii5Y+0InQqpRjbjUpbau5Df
3s2VNxcNkb82DqUHJq8QmmGThgz0gbaq0VCCSEJziK3O/cm+aqWLq3bMPcrOUzDb
d55s7fh6lwymFPe0I4SADLxX/gvGTdkrd0ZiGBtjD24QLEpv6h/5O1v8Jf0kKvgk
+YUV43zTaUs2Uawm7a9cuZ4JyPDlD/e910oXvlLPfMIae25vfimYI/pu95fFK8OS
efYHVPpxt3laZczXAFD/7/cIwxxtPripgdcxODa+oV2HaJO4nNOYSsqYJfgRaDLr
ewX3cMw77w0i/Z9Ss8Q/VjQjU54jqtyCB/umE57LIqpJFCYuIIYq0jYdM7AYtgSo
WzTVlq8c1DlYPVzefAy6Yc83lJHXnFX4Xn/cZm/xH4XLg7RKyITmEr8WwlYRKnrN
cQUAwKt2itNWxXnoTpDxy3G9E8HvH2iaS7c9A/rvRMi1MCj5hNvwpFcqrdfpkZM1
0t19EnDgou/owalDuZ7fVP7IWlSWee9l7mOWDw8X+HwY4fjdMkWaF8YrLGqyw1VX
NPvNdkOhCS7Ot895ZcqYPclmL1qSe/ctLFAADfRT2fcMNotdZFvtGOKdre5tKTam
PJ3em88yoWUgzBkJnFZjYtU+0NkGHpMpueDt7IK6JZQ3cM6Eu1sR4J9lok0LqlPq
xZNrsB8WCGPDW15iW+tgxGGoN24zLLA5IPvoABgdDqq31oRAf1hO4LRY0o4wJiAo
4Ube3C/qTC4wHJbfmgFjOFLnCOGAS6crllyPPs/9nrid3qM2AARNeead0CYnxJT1
`protect end_protected
