-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EDAgESiXRqjVHH6HFQjKoP3dNA/pvr7TzeG4QcsqL9WoM7M3wx9P7vEF7CX4zISqjtqlI5WyQLBI
mY1Sr1lWKLkDdNHpGVXbhHRIEUNqsPy8CsghO0WubTlR6qnij574czzH7lAXnv/RDn2Kq02+ppYb
xppJf1jEZYBDE90JtobvmUD+1Ngu6ByvQlFztbAf6mRsfgJWyooini31eqHtP4HGkWcuXi1ItTXT
LwNVXCP3eMUNJCg5sfpE6RsUqTpfhsN7wVrK8FAzBfxtc0RLGqw8lI4QEDQOPSYvPyAGEUNNd9Gm
jniUYm1uNszeXVOzbRGDFxU/ke+JiYt1FUVBig==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13664)
`protect data_block
q/qgjG75JzXeR8Yu8/nLtwDXJS42wkDSwnXftdAaMa5DD+1YGnmgNTpdfWcG3bC7YRPER2tXbSm1
qoy1J0X0tBG0nLL5FJ8rxTrVE72lOmnf9/A3kJkZB2xYlRUg0unKGpLwC6txecZk0C9WAAR/I2yx
hfX112DKeR0pd3UzhCpPb7rwzOFEQ+LYJsi2KDUfp7hE5zNc/iTl0SYgg9YxVNQkKvGU41h1tUZi
jTmu/Wr6enqgjdF/sMSi40vwmxMuWYHU4Ns/i3pxBcwHD1EE8DLQqgrcux0TqkDnUcUC/5s3RRVG
35WB2PD/qPF7pLjJr4y2ev8BjaeOjOursK/ujrz2fRl+/OwPj/agNIlpldNazGeOxwQw+0RXRGpZ
gyu093+/z4aBbkpbjLPQrKuekXQHt6ok6wJvk+W8tPZPgd0a1lv7rRdGhzK+EiE4prvyexaeO9Yf
Ktss2S2dTPVyYyPe98qK1Gc5NpVwjNBoUz3njjIBQwaX8MkWdZYhRGROJL6suOEmQedt7AacUZtq
MzrbM5K/7erl+l/qKHJ3GhZHZCK6yFcCpxpwGnGnA8as/iK21GcS3txICWagm3OgwVCT2Bhvx+Ic
Ru16yI7wttiirmGqUD5QrusKcpgpaZG+19XXrn+qkdjS5CQUzHPQzgqUP4UBqQUk4c1/swp7Zvfh
v97/vLVPMfpLzTiN9p3jQw9Ue7d08CkMpDcPZEZhJKrfSf1dMOHMIe8NpVE2u30SSt4TSAT6XYNi
XvGbj4kfTH4VVVivYQSAP2z1WZWTOLmuYcqJt1ax2jNGr+FoZda65HeHafu19eL/ql6QCvMfnKps
Yxm0ZYjVpMf9Rzl6oPNlkRShl/iI3Th38fDHB4XGFlxnLdS86bs26eON8W8VZjHFiP3CuWdxShJo
faEIeg4WnCoHSUT1e07oTeyfMWkqit9BN4xlAAEUOBxTgewgL+8L1OL9L9v+vOa+OXHfhK2u7Wfp
joxzPrURLnj8iiiV5hYDAtzQasbnme3KD+jAH+CWs9Gk1NFhr5gK8VBr2K8RS2RZeukiQccHZzx0
HbTs9ZdoAKjQKeQBLl9YT4VUH2m27OGsMQUvt9JAbV78wIOrowQeIEEjTJaGphjQ0OMASwOZEBLN
spjVi+HomiiqIxv4wyNJxRVabzy0kPf9UN41ERwLffZTvbbuEVudK9RkZJx2OZns7yVLQFCeNFrh
Uq4WBwmghWnfnEDHfF1gQIrexVrRyRj8PIJM/tjzWFhqHchyXPJ5HRMzWxZ6NdGaWznvXXh7gDN5
2X74jAOTdLP5owhSM0ZLNyYdBz0P+1yTvlXLh6jUIF9jP3jlnUHkidPKaWmZVGH5huNxAeP79iGd
caWyAE8aB7hveBZ1qBYwA2mFqCcrTtLzTV1A5S4iM/dye+ynimRoYRtE16IVJm0KCNOYrkH10SsS
zYUNctx5JZdoHD9a5Xk34EVRkCd1Fev/lbXNb0v8Tg3c6E9vfPj716vQWv8/gaEHkV4UKEVHI8qC
Tr7P46h6vTfoe6XYsYbVPLO5mSS3faAupQIsRnsi5tvMPXaNtFH2OwakJyPGGOvBej/Hqb4jDd8/
6bQ0EAj/tp9f/ppFkdRchJb+5oHRFoX35tw4QlTK1vdMSeinmDMLUfjdH2OlcMu9X6xmie0qgHBj
6z7cPJMRw0sKb6bV81FRPDDdRg7Jlo9mufwN/AVxoqBnSawJ6T+fvbszzVyi6d+u2FkJcvPAeyzZ
RtGQGWTm4ZCqJwFzwyrIVzJC+4erfvKicgQxN2f0xy2btHbrtvfpzTlx099wWoFgkW8vM2L4+SxC
CsQkys4cCo7ClYNg+4B54exstYVHG9Tw5YJdjPE2m52PCOWFwLjXSJEgZstpsj2E3kfehaix8n2G
Yr57WzXfyV6ZreSC6bTdn1Gwurg3JEh1eFlacul66L1brHxdPFRv3lrjqOczZCV2DK0XzLS/C5bf
4W/LDSwKxtEDnCbhBcqRV4LDwOFIEhSpo4EAKTVRrpNDt2CAzbr6b3/nkhu4HcBpPkkkcOw9UooI
QERv/ah4oR4dEY/9i+INcEFSBgXUGq5c8YEGgiK1x0y13sP8kYJRnCCJvXBEg/WnKNi9r+mmPn6K
HN02Q5lUxXfioCWZ3li+2BXJxUf8C4qdlRtEmuMFv0nXwgRcJ5y00yzoYPH03pok5gerBNem3geE
fGMdnYj2U7H0VkRyxX5k8/cERXIMNGAF/u+S6WYUoMHAqDhpC6xBWB+aEQiznkLFs6bO865iCedt
cNua8FcIEYLEpLGAPV/FIQMKo5aHW4IMkayPwgk7W+/SlAMNNd1sY5fLAeny09uzN6HEI/S68/kI
DGla+y3lYY4JvTiFbIHg+XyP2oAHiv2DoCDh60x9acwlYcjJHmjQL91NGOe17JHhjXWNrBa5TBWC
obuJq0giviPagyHadqsN807B4v8Y5ocywuLkgbokKDV68NBjjoHiHYo6jyJHVVC66zQOrEIff4ix
Vt5Q5v533BewxThR3hyrRczybfffuf6YGKxkw3Bd9GTonmzDCBgeXVt2l7C1Vl0PtPDYinE6Unz+
DOHvhOdOS9+fPFCmTQrByd9/M0UY/rS4uJVz1qMzGXqvKO2G3YNcv2MT0TE5G3anZFt/50wJZnq9
LbKbYmiTYfp5PwhWs9k6KGTlO96z3cjlIx0BDODzZoAKSfr31hRBxfl0Pnd8FIysUxr7dPvYCYJl
P6FN/8Y1E+OMMNHmUCjSSnWjSsBnJj0+mnl39/baVT3YLkbkSvBm3jN1gaSKZFjSk9XuqVcGaX3C
KUcug/cK4VcQshbczdVdVpC+Yeo0XtokGncMKT0QGJajIEKHUroxlTk5X+79LBfQ6eu7ZzThoAJU
GgU/7vrQmgGSh642FZCa4IX86Qs+uiI2jD3QHgLSsT/QDxtqKATm+MB+HSqZC3UYkP75d3SMfg8E
JLrT5+Rz1xK+JC2Sbwbtm730zJrZqOozq3k+YafgWkocOHMHsL9e3VeSQERE96iRdwXakwfOYk6O
FswreNUkUwQYu55RqRoyZyHodbncRaTGA699Ufg+zng3bha8MoXqw5cc5cLI2hllFN8m/amTZehj
kOtzDIfhqb64Y7Z8qPcupTmh4EBvoMkaqLIfjJLtZQq3ugIoJjKRLxJxU31axwGy7uFehNU6AB1e
tyx5hTEs8DLnXJTHSYxo+AM8E69g3EoFJFuNKyfplq/ZV3d0u9Fp1r+fX93KMa8nVG+NLb+0dCl7
+E72xG98X3FB5JfCk6k737+GsYsO2mZ0vMhaXpRVnS/VWhmcCUyby49D4KecZ0DLHTz3lS3T3IKr
AOP6scsdIy14Ttr2l4iqu9b8vAIlD68G80a5y9/GzpjN6O1f5Px57wgspJ+9+mXq0dPWkI0srKfA
MKrYElbs5vkwNumKC2TfJhXgfQbOt2dAmQN6wW7aV/OslTL9d2T4Q1DcX0wdpPrxulbR2Vh6q0Zm
bu2huYdiS6d8i+dTg4kJciLyLA7dyzQGtv0gmSuJHTO6Apq+DRyjZaYiZLlv0SYzHNp3V9Om/FsW
wh8WbcWZXqjL+IgqVhxtyB68lwLIrcvicCAqPygMJN4bbFC6VBBBAlUh3MPT8eJR1UP+Af4J17Xv
z6R7j51yOSWvp38lcJkh9vL/ICbGQ1k6y2nvSnLVU6ItwYrCOMQ8GSppBGMtZF0FXj1HA5ch3735
feP6/4ClrFW5tZ/cyi7ZZF74ruu14Qwp25QVFPrUIB7MA/mtgJNI4O+37wVIDDsdCB55kreJqrNN
rf6rGaNyxmbfM8bW5Cnna281mxMpqh/R1S8bm6HFSm3RvDnyOu9cJQ4O/cy35ZemQYLSh5qSzWkh
+Ewd+gQsQSoMdpdGppBU0hm/GWvlTleG/hj+Ub9xglM857o9JW+IEAJNrF47cwgNSeZ0k91FMB/r
ycut7UgkfCC5YHBmGfj3auDqPS6nAdaK4qJrZ9UiBeofeKTG9DAQOjW9siA3k9gO2m8NFKo/J1RL
YYLOXS01LV4QLhfEva+J8+o0TYjkLmNYx3CzOtltZAKY5LMPts5HFP5S7CbKz+bOMFGObmx9nW8h
rZHBtHt0MFGmDaBpIO6HF69JDO9zdhrsEuDJRpGH/7lFaW2n0JvPyBjzyl0r7T5Vu7Csvmu9htmf
oPoQIevYMqnGKxj5NsaxVyjs+t+Owp7lHo0zgnRAo0UwbmTY1EEVPfLmFSg8wRCXvXBn1FE1a2Xi
7sSLxijq2T+jG/6VDxf04A094qfd1+wfL/yI+VuvDthdIulzbknxGD9hTzgx5KadBT76E/3onU+2
+zXgyQCrwIZIYasP/1J6vaKto/zMAVH0f/xqBDnDjZKXTyv57LbL8Ptxsk+cTaHf7EiqgN82vCdQ
96WRBWjUhtH4M9o42DrWxV6824NMBP0OFcY+gitQBGKAB0XrTVIGwIWFBzIE269JrzH0gKzkEx07
7/Pv7gZmHYVfqpLt2pNTwSViYKf6JajU8GqrsUQByrrgEOLB+/74Az3fHAPAJZyuh70ENmY2llf/
Nu39qbkR268+pjxHIyZe2KVZGkYL9KeFPxrTyPecnzLqGB8PvMlgLqA5tFBvaw+2OgpEcs3GVzJ7
17DtcChLmD1+2bEMXUTyqHPvZpSQjdEMjWDVTJK/IkV+UlGAP9/jAw6HJMd040II0I0/pnEl3lOp
Z6YzwmBCGWbV16mlv0ja7v/QB8QsKBA97MEhYhf14jsGnu77i3v55IvYMP0On35Q/kjkF5G71MDi
Z1kBZ9z+YKTXZ6bIYOF8+ja0Uj+td13qc/T2zQTd+POFVtJepN/NQfSFUCrsMsbx6BTwhWq+30vf
Uqo/VJq/mNfMsAgxd3wfQ80qpjLONH3n0kXSe8ZUbsLmup8u12QgX8OrutxDSjUjHEWsvrQbshIc
eyWM1tRiLPCyjewZ0tk6ZXliMOpoGnRYY7yAqsaJ2CZeG7NHxTAQW9J0+JGP6E2ZaMwoHkNADDz1
VBLsn9hM3K8D1x7qrhig5THpw9o7kdcMcuciJI51+Sh+yljhxKACNVewdta3bbD2xLG8NyeqRWyd
aqI/Ld/wBRlXKkX5wXSxW9OgfdTEEr50eoCeJSXav5uJQ+V6kJj/rqI1IuxwF1KjDvtee6iC2Ocy
OiBu8FKFrsbaCbaVnSnpQNXzRsObqNnzWAQezM+lNidKcMMc7FWq9sEYcOV+jmvpGhEly/83n+Ci
2FIuoZ1RLzZIxDIKvbNqUonaXhB2XNIcwdSFok79YEtS1sqqCvcStvaGMBi0wpDE6zN1P0WsMPOe
l1SujAkiN6rx6vGuzh2j+DdtutTDtBFJ6m3J00qzpmT9ZkjvSmr+6G+J38LEJOy5zDjNFpo8V6sq
snUZRgoe9YQIJj6C9i6s5/ouuz8wWiNSLQSGtglkNkLrHrFNd024yP+4sFqH05ozqqGfUy6lcVZ0
lFfYLGtWbiriDJu9lpCKJ2ij90AemqjnTXKo/VfhafKSIIGKJjRSHlAjN+VTlNrR8sYIHR1lPIFt
ynj52rRNICABAI+AfIalKcMcoU3wedw9Nu7Mt+T6s377lroks9QoyOqPZNPaOQHs5QOL0YUrl1ou
7Ns2rEO7ZkDXySYnh/LIzYGPGHosA9j1MoLjjPqe+B8FxPd3VaQOKF+xmiDgJrsYJIwkGP02Y7pe
69ovGr+8ZfTyPoq6AV8NIMBvSlu9nZuB9Ob/dF0+eoi4Anmmes155/ngDuXvQEGOrCUlcVfAiNDm
kqwhQ+qAvRDY7ZEyYnF5d9fhZkm6Rjf3CPF4CtXBQ0eegD/9ZqLPp1J/SKMwPW4yIMJns2HVnZqU
5P9+eLz8vMwMKgI2Ohroe45/3njWad0z3JUAsOPI3n5YqxNke+JP+duIiEKHTHgGwYmyOXbScENG
xNrr3/slEiUosNqW6jplb1Qwx8V8/r7I1kJ+uZeHgSskW6qT5P6OPXK4MmG9ARqmH5PjRmJ/xv+7
R2oW7+KnBpyzI3y0O9JAzUfwlxYyC1bNPf4dIg4Y+l0kihfFzL7q2N1gy2/ktY052Yz6NZ6JpQYq
cgTkpWpSElRFsqD/VW3nEhMhfGvBsZYrwtBfcceLkiMxJ9Xj+V6MjHd4SVFpSV+ZXUs0KAqieQpi
a8M9H6v4aKi7KSRvRiALSOW+O0uFuGiJb7WJ9TEn3zHO34p+yFsWu02+V4yXeM9G6vqzUuD27U6a
OE1LFgGQzhXp3jU/R2utbWWPisbxqh1EByrMRrJq4JUOJKqyAb5udhVlIlRp9Hmt0zcr2VF78vLc
U3Wprm/PK4oIZeyDD5eu+6mKZpjlTqrX9opiJYwqXMIU5vYI0kMk/hBBZoMP6Azr3byBDZu9xpRa
BDpVnyaJQ9ypZoPfCBCST6u2J/JKtkEhHauc5S/52A0gF4rpuZ4vx77BsL8/QHPq07Y3PbW+zf6H
EQShiLWcXaQaMM8j8rJrK6tXhmGj6nHKvu5JppqLIClLSkZR6bDtBKdER3TsZjmcPe/z1Ynwo4jT
5C2pvAvTS+2+QwgdNaqZClGqnZrdSn1DAI6jNB85cyuDmXBZeWHb6l7zWtbcEpW7+LxbChHsHzOc
BsdSi8iFTlHM8BofLDmajoRhXAEPq1uoWuq6GA61ulAgHdDdGmR+A5sGM8dSS1sfeUa2pdDT8bsi
GRpwt14DUe3P+NOyjLi9QCYmX9yj+dJCK9kXrwRbTUu7At2usq2gqAHQyOOCLiQtknVIBqOmEBFE
9csOCoIQUiyXSFqPX5RXNvFK5VqfaXl1OjVFqtKKipSum3QFlYzIHWHYza8jKZi+zpD3jRtDpyaR
jSC0bMDwskwIDP2R39zrM+qon/sa1OznOnmlb8Lx5sPXdaXB+8I6t0iVstnVc4TjzgJx1wwo2SFr
YW+QspBkjuMNM8pgf8sQ/WsOb8RvoR5q3QaeFoFSwlqWdDWm+ijOTSaazfXHTWVJS8N9/keXPoIS
eGq1nFW9TvoWYttPc2jEqSriP9bCTMrmSIbyysjbi/j9mDfl+9+aWvA+IPusj7A+rA+TzjMoRvve
jW+UNe16DylnpS0ypD1IWUxBSaAQ8Llg89C+GyVzqSef/sXhspzbmeMpxvrUvUmalXGAupQxSlpI
Q9288WW9nyYMpK6qHWaw3BSTtnzaSnptIjAgtQA1BrIFpFXE9rnZ6XqVIo2nIabQALx1qB0Ogmj2
wmP6BQQnpDhqj/2cBBPpc6OMM8yypobmGqb/BfcGAlve4rKidDhFeTAlPqMGW/R1XB21fgPNnOC9
e4ZP5tdkv1oogiU3m89W1atARdsAcfboKJ+jnLR/7od4Ws3DXSUSdt8x2wmmFLA7ANEB97aHs/h4
2C3du9TH3j+d8if83H3T1a+fORzMHUObKXwHnKA8BFu93LJSp+kiv/1YK+RrlOqVdd/2dUnmSVLW
gvEzN7ItRx4vkWDPSDu0BMQxGWgIL+Onb/qlA6wQK3YYBK/Df0mN5FORXV1QSeGv80nlZSZX4dLC
CoEa0WSaqbV5X3+tYKEQCs6+KPkmDJ6DTaj1Lq50eGzCdh6HG9pJAWxMyOeeMYfqkTX6fcJ3hd3w
lqSx+yWLCQ/TXFkcv9+thVRAyFeNer6As/G547CXBSh+jQrurkUdSRA1wwlpcuvVAh4NM2CKvbKR
6uWlZZFxy12VQClmcYYOz0P0ck2U+d2ofj24U17f22Cd3gkr+3aBenSRWy0UrHvRELWufXdmZo7M
0k9S8Xni6RDUHN+JI0JgBG3QxLZ3Om8jxCdBzalCW5LiAP+bbpJ0iIZBJr7X2t+b42S866MT9+AY
aII6JN+LR0ZCvmRP0OafwjGY3mSpXdTlxEfzq642u4NmEU4WAf/9AlqPwaZQF8GhBX1j96Jaol1n
hznRgqeyphoLrRRM9qW5fMNRBgiDOJx6y3c2/9SKZjVeAaFFjtPCe+OIvYYQvaiT/tdySB+NqKpr
xUWU9gR6Mbbx0ib4x7OBSk0GhkH8bC5WkgaW1cuu24gorQRdrFhTW6hPo4s0zHdqMxgsd4fmo9Yk
kzhwuDvuwRlZz+Jjm9EXWcP8r07rBVt6lMUyVQRvECQtPx+7cpHqhnI9vGaNLaC3ZYjnB4/sCQn3
VxhEsU5wTVJRzz3rlPr0UF9VzeK+YO0wxuBzhSxZG7lMSIqiDO7wO0MFNGUhRmF64q9Zi//xES9m
8nuwi8Cu5GCTC0IiUE5ZMkCmDC4iE3W+5hGY/UH16joLmcVXjnm7gkOmf7lm0pKcdFUmPmBpMDRa
azdzv+ZfMRXk1ZBMY2EU2lA0cVAFDrcLhtU6fJdWV6mTS7VRdptqgyvQT3vrSUtXYwD0jHKSt0aF
vOmrwqi6BdwBIqxMuQnD51jQ/1gn7pSb/+kkkRtKfOmLGDNv/nuB+wwdvvR4tjed+laj2NY6hCGN
dlyK/G29USRgNsg6NPgH6KgVrAuMJE08g8ytieBl45eYAHDLZV5JHgV7g9IlFGTez+WeJQePVGyB
pu0QMGIsd39p3R5DjEKd9JagVeqIVNnHh8gI3w72iIx2sx98/dGZ+m4G7yMZaJxaaIjgI9qm+0ZV
k002exS0eOTuQwAtKhleBZBbDU5ggKOjePCmHjmIkiQN7dB6u4KwnN7u6TscSWulyy9nDUuJVOHe
q7UFZqyM2ER0P0R9TPwpvAzj6O9KdIvqal36tMGlZO9vl05Gf8LtckDYxqWOdkZIyrv9bo2FlGfA
6uGtUMdTyWNfny8ppy45bUmysBi1rYfLIvG1pnFk8WKuOPXRMV+/RFnc8scqqSl9FoDfytpny+WX
6vHmma6aBdLWjmKdsx01XMJx4cZDYLJEcVWcGm4RuGJQA4yJqfCWDAIfs+gdGuXWJekwlaks+ngl
cvxIgZB801UaY2p0QVmsCNo9cvkMibGlS3pN3/onMdRZhyVuLas+sfpnRAmlD2ISqsyIbnEMz3+1
UlaXNkAAVG7IohHDNJ0GkYB/zP23fMrhidQCvp7RfMxafm7Happ9Z/NShCVTAoPyMz2A/ogGccVR
8bHLIpJG7sLTJmWQEmU8nT5ndrNoSs53e3CgSwz4e05tUlpGlnAm4zB8+OgkjcA1ExFRXlY/LEif
FAlPyyR8xibJUXcrXOr//MPulXQF1LFCOwIHUsYy1TM8hffLuVqBqArJT8nZTlKIG8PiM0fKEc4h
yNfVgDIo361Uiz8YT169zTZchWlewZf+Y7HL46Qaiu6jITIgKR7n4d8ESQPve2auzWvpoiVNlzqf
b1DpixfuXXpeHrkNCSgXWHrsHUzDop6QZx8BVuZmhbBJ2jHOC7CWZDl76XgX0L3vU6e0YpPgCaMx
RAwwMvFz85v41ndmcVRFmzScYzIrKdxnveWha6Cux56VDdMmVYNEPN/OEmcdjPqDrcyB5BaVa/Sf
ZrVfUXCzWzOgh7AVDG4DiKM2eLeYmIw22xBCnJarcScRWJLfX/Msp+BXxX1m2dCZHJ6OJO6nRfTc
d5Y8znzqE0dy2Zf+5h/vTQxhQbS+DzkzBIe1zRVwOhmkPVrsRJQA1E165eA9VZfVf7c2Sn7lKiNL
b1geUFoV49uZGrPBr0jItSLAVJGpVdlLAS5/9m6OYZLaW48/J/xW1ubhlmuYyU5Z46Y6OAKvWvm0
+dUgAMxcl4o9xObt6WuNzfzUeMEaOKWXDv8wJUTUSmPUSI1DXnSSZ6iaHIYtqpSBkIwtRnPrsnVR
BiJ209UkRqY67OhNu+mqz2o02D5Q6UyqkbfcFtPVKD/r6pXOH6E90CCAlmSaMPs3kCA5pjLhei2N
aSEkgmaCHdmCq2WQoR7Uy8V2wehExnKpNsAp3XjNdw/yTfetnPKyaJxd05zb/FA43CgnZMP/ocms
JueDHXSYDt9mxM6PIHZ9LlJ4KXjIQv10ff9KWkmd4Q0Hvv6Dz5L7mnryTml1FRk5xXSQvb7evm6S
fiN5puiO3LPoy1tw8p2AigLLYDDBors2pmuEErOE3fa/z4XhCA5YgbSHEtfe++rUUthAgaBXIWKA
LKVmjKvnKfZ4Z8Bcyxi+MntsKQx60ZqNZbwmZxgYZTpT9TiMJ3ADDWUOfbgWaR2wX2zwKM6iSYWb
w36NjIel2462FX9kgzKSNsyQnPjGBPGNVGaNyMgTN/Slj3g2mG9jsMGEmzD34D9pME3XId/LD8lg
txGmnk1FVtb+C1l3okL4ueLxhMkdnaeK9CniRQIQdjzWB4xlbZat0l6gzR0O508PF3kTspzUESjJ
Bo9A8NcMunrjTeIyAsMBVbTqO11IGnuHAZUtgp+S2hj8bBTVWuQfvDDZxfT7i0VZqm9Zoj8mxXo6
dbj3SKfh7TwGtzXW896KUpu4bPC/XeWVj3f4/4n7+BqAFNtincaCPxOcDbCTU7u3Pna9ibkRdc2V
XstmUAfqZ621b2Agc4a03/aqkLF9MY6u7e1M7MJM/KXRUvKD/COaAdaTxWcG01WtbISRs+l8AdUm
qMqRJ9XnnbAtgl7j3uWpMAjPmip1JAeNcBtcrz3ADGWAvx71Bb7QKi5Rigw0vyUwsmJdkJws4i+A
ucvfhMiayQUEdPgIAxCxVbrvG/xUGd7frdrbkPBcDTxU6GyDdEj/w/sDLXUjR8RxBpH8nsSQ1Obv
WmULIOaNM8RxUYR9BEb1oypApz69bV7TBsGAy2kLMbBU1FRHItzZQC8y4pVE3KU/PHokDkXEki0o
yoOxkuRGTOSYRxh9etmrUaT+1CqSbOw5OxF4VfpSAZHjqQuf2Rt0Iqssgh1xSMotI2Rkud79dgnE
WzTYlz1bazU98BWa9nN+Wc6/r56fa6xTfGCBX6lFWf3Rd8CPTKGBE3hMqwPJvTZ4MKIgThl732Rc
klZ0z8yMKeq+rQbkbVO0WzvFcRMNSxID1VMOdJVtDR8rxpAx9K3zKZmywKq+/RgSFDjtX5x0zb3a
kpaTZXhxhAvP5IqeWkh5WOkfSo/iBpa7jOhBZ7BfZeFWcZOOKr4jEk8QeqVkfqXx8Yo7tXXoXMih
N015woepqZStU1H77oPQCjtHg1/7sYp1a+JyDf5DZmQy2j9WKXycMbBKByvOlwjygf6Jej40DDMD
qAlrnQ+DvdlDoUTYh7VHYDx01ZJyiup1Ke5+fbCK+U2RPV/bug7tPvCj1vteu9pCQQfRLfiM7eKs
0ixig9yEkzFx6hVssfWB3BX4EHi5EcYT+zq5cuRXAVGw3UyN0f5D1u0D2h7Yw5BFoqg8BDYRoEsN
Rwp0NHzloesNe8ikiGMC/oPv1OKqaKkdxLkKMskKx+GBEag4BlqhjHHvIF5lJ50YuX9IcjQtPg32
/5vBxWdIAGykXReCstliRYgQCUKccAJOvLSARR3wIFDStODKwAcDtLV1lUvDKwAaWHGhXoY2Py0A
MNFTz4IyLodijTbQj48jvBL86TJXXY70aqgmmUwtby2eUiqDNWdVHRCNRzhWdp2Oh17ZIBNbqW52
kiYAOSXlsTC/Lztp8zddAsUm6qGkwfJL4H6zno/V0q75y133NK6OOx0vsKexaqbfcVMwWBxo1Ztk
+g1d7pVq+tQjLmqfRBH6oIhkHhTCxTJocJGPFEYGhyeG8Y8XY9dwWBTXv3LTYIl0gaoNcHPNeeED
52iAo5Ra/QFUVvgCqsKpJZnG7uAZ5lTLoR1967QCAfHkQuhcxAM3f38uUKUxyC+FOrAC7Ce6R0SZ
9JAZIzvv/9/IC5wxq7qrbf5tITjGF9hihd0PLU9Ju1AE0DpBR+5gVXp0BwAUFqqjFHPevFIiplG5
VV+i0Xe+rp2ZmSmVwGKBHbACUKTCNpoiwRJhPJTXLhE2vrr9ytGE0+UNomJtKWeATB54hl6M0TWg
T0zwKSZ6EKtNVkxxcW8v9v/3jCLsyz8OwcdZ8m1DJd2pjmsRuVcmbzV10YDkScsqh/n2Kb1esRZQ
zAH12rRFDGV7ol7VEDG06buMxP2axHHDudbQOKJndJVGi9otqfWAzATTSkd0DnnfP6eTOeVQ+wlK
4dlY8uemX3gjPrPjzTSBCFxy+i+Uf29czY8X8YB2svqldtuclqgjacr5g0DhRDHOJEFzbxZ3bRnT
KIWGbiTotk0oaMuzlaoxWk73zbLOf2IAcSWubKuuueNakPhdryrqZsn4X3sZ2xU1WZzmS0qRAbq2
moR+M8M3DM1vfa668PJP3W4yqL+3rpMURXZhLDTC3qdIjP95IK//yrBi0Uzx/e/XI9XD1Je34bT5
ZFGCoWloIimq199lSLrCLtxhKUDPcPKPu2uqJNQJVrWvCWlKRPdJ5YognjmrG2jnFkuWPKisBGsX
7O3mxrF5NMDAqjOt6vDTg7koL8Gh7cpKqelfOuW9U0KYvKR9Q+nhYiMV2xiyhPmI68eJm2/n39rX
eNxXCFj/tg3n56MCGdXwvOmI56cmJUk0gr4tbmR0UzCBCqGBEPzw8QZeaE1nYVVdO1FvHMQgmzwQ
F8PA6sO3gFWSXOBEZusIypM6QgDc2nGEgqJG3bLTQ5OStuo6fYceJiFpYMV2VmyPdPUcgF13HPEc
f4xNRzznynJJs7I0HLHFb78ryR5GsL6sVOnBmTlvOat/rNR5hc8jdWbrRivlMUNQxfpofSXvQKDj
roFNATVGlrGtOxcF4u97U1Jno6vuC3XFkfWa3mWo5fPSeByY/1+P+jA23+KBp9BV2C7MoagoUUvJ
UOXmX28Uz8WuKytff/mnVp8UbMtUVGj62sUarsnYprQHLtLNiEUBj81UYaw49XyHVbARsIWCoTw7
pR1DdVbKsujoy8HQMsJkGUc0GqxPGAEIdqJOnyiTzST0fqk5lWt4hbbrc7SXFg2ObUC1sY0A+OGh
H8+kdb2wMaA6KCNucIBUPrhRWX8g43HbD6KEuF5bY3+DvCmcSiPo29nvLF+SQo5yhNKMUJ6wMX6e
LpH4sV0p5aqNy/xfpDRPQRXfXjbUd3NKwA/ZIejbpnwp5UUiRHIQUdtsLsI7zUEqDGQf8C3Tna3z
0A70IFqxc2RxItBCarlh0cMKcCfCK64xnDpjvQzJt0duBI1GNzsBE+UOK+Sdy9XNrVHIvAxEEAQD
kjfR0BG/i3k2R5sTTzAKP1x7gfJ6qEHg+bsi0V8CIrW/FFSAzHx31cQcBDd/2gQ1qPxoyubLWnwn
WbIBK0AQ/1RDL+GCN3G1Du7sWam2doq4CCPjbyH+6mXAMf6hsEhkOcbMqxVDzGg+Pf7a1XGLQjMv
OwLxM+v6Y7BZD+zyhu5CBLcAvCIEkvapkOE8eM1qlWaz2PWLKeDW/PUjIdoT/kBmVHXBlZWQu0ML
ZtPp2Nf1f9DQ+pxNRaLJ4JgH+E1zub/tzeTiHrXqJsS4YE4L3sJeKrQvUkLqnUyEpfNtvzWrTLCX
l3IpQOeBAdm/vXmwqpXeINc2NdveGcw2UpJH7of3AKuS7d7SqpaUnwrXdXVf1blQylsyDs4uP7AD
1Lr/jXe37aJTrqjmOdQHUngnRHbNO6Y6t5LU7CpwRgcx5Sp8A0QF5wSU8/RTd01NrHPDGzRz5bq1
oVI2Q8AyTC/70kVEpweajPlnlPB3Rf7mzCOZ57EaazdH/fdYm4g7rqwQBCfb2U0MVSox2Fk5Ont+
dcuOz5rDqGEN/RCkQyewqOGBDbBTsQlrhxh6qBL2mZgPwU99JlQhVEDVTzISjuExgR7YHU2Do2bM
SI++xb8g9ME4p9+uGffIlU26z4B0/7xqs9ew5XiBbn9gcI+2BIRYNipWBnzk9IXHJQ0ccAJlJm3C
aax8bqey5m8TvIS/gsFwoS8ebRN3wx5ip8Gn0UulWoEhlwCZyD6AsoL3hZ8dnIs35hGncKqj/RgX
d28qJhpFHodt9T25AfddEJknAlAvA1FjXGUtIO0AbXXWD1Xja10CBS4cLDtOA+7f8dEoc1bRNqLo
nJ2v2KaAcMMAHuUfeR9tsBXFpByyFE/PYmoecGzG36YS+UUgGYTihUapVFc4mnboeJ7Zfcgmg8Kf
x8J0w/InxpjQGKdr3YRNBUu2u0ceh8LxtoaVl2wyidLkCEcTmCz3FCE7tAWiQH44KuhMGjfT2E2R
yTQFV6tNSHG+Jt9kFLAWER8C+sNNHxiLp3/lFz8YLFWyduPuydK56yWoe7yumAmsSqXhkp6fvQEp
5f43BmucMXKjWO9B7Wo98hb5bzMUlkwC8pa7WGXDdBSw6invAZ9C4faIMNVAA+szl5/TQoSxcKbV
Y0lSq7152T+x7bciZfZeDfcUR+PI3QTMGgWV20YrCjYTqmte/zzTOIldDfZFQm2XNHnQQ2hXgraQ
CB7bm0Wza6ALK/ItPvKxmzZ9OExs2q+64fiOIcpnFafMyBcMiXnAW2d+gHOe5/KfuwQGoZEI4zlY
x/n29ms6okSrXAC2yV+nAXi2R4uMZFYzjYhuGJ+tf+Wutqgu1wgtajbPlN5kBbrcraS37TPYbdaC
4rqSXXyrXhqE1zBDcrIZ0o4zcuUQze/VSwWkFdVh5lLp+RlauzoH7bVeGkIFZU6D8TXJoSVAR5kU
izhUQVcWexqurgRAwpvSDlCA5EvdZjkOI0i77x8Ne5DiE2XFeJzsGhsiPSwYzzqUCoNACZK9IxbY
iZdEYygU58iey56nDDUwzu5PL5ycYDKl/DiPH8GtT9BCiattUxUyryiFy9acLfkKgjBeMq/z/Z+T
g5gYWGHGMHL+a1rXRwfRLFnUcQaXhpEFC06Wwdfw/RRhgkPsUpUMQQj2vnFb/kR5IkeM9C2WHlpP
oR0LyVuQe68kg3im6FcECgZWIfb4Mc0fjxh2esYhG90iYFSQ3gIwl0DynSZWIJePbh4BHUbUQABg
tT/XDQ6HcWz5uHzhEwi5RkbCeC/DM0vIWHZL33MZR19c9L2gv06wKnZWHH7HNTH0gAgslg7hGC94
DSV7qBsLzD9cBUJU0oj7HXDJovsk+FEbi63yzp+YRbDkfpckfhuR18Xt+PmOaNWI9QqkL32PyrCi
o1sTeIadaK90Z81bkG+QrFFsi5QXvN8a8mR04wq4rZ3CiYF1noNWI408uCjvHy4viXrvSKlTQNXf
iHWc6isux69jAQAGmoUkEGyS82x+78LdjZ76XIPTHXO9l50tMQOM9gwL7emi6O3Vz22BfPzueATJ
Uqu1PGJXW1FKHcYsUtrjm+Aq/NReTDNCZpLxE5m2//WC9B3ZulHIttaMBwp2qCP3H+DnL0nDRxdV
L8A0W6wjpjlVTt9qhC8Lp24JMxXY0PryMvTg4qiuErcq9pmRroAuHGJZdlKp4nbuEeOZYUz6ZoMY
0LtdQV3d8xTHJ3MHNCv9eGvsYkm782WnPcMXMBWGiCzM5s6x2Ra3O5YuubU//BoltU/z1cfkhTiL
68hJnYCG/2Xe89JmfhKGQ+K41e+o1kYnH2x/IKHIbgm4YDy9Nm8Z6myssNFp/iz8TQJ/C7PKVuux
hrqSNTb2uM0Zh0aZg2D0TcSdW2ObNjfuTGsXdc8YB+J1VAwX8LUh+DNsdm7VAgLYbgD1IiNhh5hl
cWyxnnN27jTiMGCMgW/T4JDq7iec8si/pOSRPOtcQMor3M0pZ0M/2O1yBisfXrBAbma+E4F/PNzP
Qp9YT6TNBf6xvjcSG51T54ouXahqipGO+o1WPghN75Z+1F5llXfzBLH8KbOqNcZVaEupccQ6k493
J7DRuMX2VlrkGKiH5e8OTW+jiOsWpCsZu91V/fPSp1NI68hsQEMmReCNg65WaWKJsrYQgoPTsCiV
VRunvCdLfHSG/aTMWjZqQoEBTYBYO/+mH8B7+0mr6CkhOmkhEM7Gbqw9dgN2GOdmRn9esPn6A43x
oKGc5ig8dFJ37NVaW8ywxfXSrn2E0s7usf7RhKeOJaDzyTeDu9aQVS6csAPEO/Kmci0T9PCBBksr
MKNcsDfMK8Iwjf19FMN7S2yWqYanRrOwWpGAkZ2M2VNuUeRRMFkfgJBOggoia/HRBw0NIiYhQ7v7
dBNebIMwa02hBuptQZaQ0cwxm00vBn24LHM3Upyk3wOwjpEGctQ1QK8C86aqZoOTuNKXyPnvuuQT
Ws3oMP102Y9U3bweClP9uDZz9WfMxqvdh3BQNu2XRkvh6UIzjYd32mmkjTAyhClUGFbpPGlPu53v
be+APfg8XbUxPlfDq3HqxbFNS354Or2WzK1cDB5eroQ3h4GKN/owpb9xxuGjOBxjPi/MzVIGVF2+
k+pVcS7HSnr28Y6d0aD3XSFUC0tEt5xbiYJAG3Mf0HGnTNtGVZwzBS+qRlcQx9D+qIMy0lGj+o6+
hWxHRHEXYksMqNBOyxfJgxnR/bzfH8w+Blj3VBalJUC1pEJADDiq2ABy2zlDHXxfvpOpxQwiDyqT
k9xF+TAYnf537Y2MBcvZKatoClVNtf5xuzxpltUHyGI3IpPVmc3LdIjX+1zPKIQYd9TyTScmDcdJ
9TLQ/0/Hli0/dedO3gjH6Iu+j/IqJFQi29TXVEHVH3ZrRap2UMJr8H7fqFbx/6scjySHZxYLh8LI
TEa8DFVLLrPMHh56cIpsTVig/R3bIkmp3/fGIYE3tBgn2QDXLSIwsSBb1k3w1clYdOzCrQAvml2w
kw7bD6akhj0ZsKP9q/PtgYucRTFdwd3/G/leETn7EjFt+3qYc380wwabLiBcLWcVT/ZBfyySh6iw
4F1TsAnxvmxql8tXgkLmRugZhlJZiOcMBEd7YjUrL//84l1gAjX/mrZV5UsZoZ7E2a+NDDtuc1iV
n7ocMiqumFKYRzfvn1P82OY/e94grqLDSz2DQj/IVVYld3DobZVizE9vrji25IZNGiRzQQWrVPcQ
U2hghVbx5x5Kq5iYblTzG0OVWh7C1ha3jL50WGnLiW40xs0Ca8n811zHrdjoPspnoc0k8KSZ7fNp
iDa5tlRykqqBEt24NwUlmWSYLUG98hs5RSmFQmjoh1P8OG9f45qP+0KcYyxZDaFaAOBeSD9hxMUN
/Wb20a8y/2bOlFQ5gMMaJ2z/X0XRRnXsqtUzI50GB9Q/WOPyLW3ZIh2r8+NCe7h83tsUeYMMSBl0
ziHmoBYGFbfeE8xUNpKjKmTA6mJ6jJkvoFFVwzBXPQoMTQLuReln6LViXYdqX76qXEXQFw1qQ3Gj
CmGTp71Z1ltGhFc000eaFiBkMJDyegSTzKJ3vFBdbc7xzE0/FeRsPt+t2PoGbEazUwEbt8UiyfVN
ikYTU4qHHrFMMxQrxqRvW04DQUIr+/Upjvr6Bb2HgOtobJ9QQi8aCQOF6SGcU4YoN5hqRRWm3zat
iCEoqZlaRSL9ZpaSf71AZO0rgAyZheUhztUGEG3jZJi6Vq9V2eThNu+Izp/d4/pIlrlRnxAnNxh3
p4Xm7/dUbcy3B5rjBqwYEzp7e4awgsyc3CnZrIPjO4f9cpoAeWGP886eUqHOYFb5060TrrLKbXsP
Z6dO86VnWXqsovwdvrM7kbSULUllhAmeylqdyaQ4mDghOtl3QKpelDbqdt5rf/BjUpzmo8zJthMa
VaErjMQw4p806r7Vt9WHS/u3wF0iKNCfsCIr9SYZ0t+W8aUrWCMxCHvO5jEEcVx5AU7hyoU+WbbN
EhciR1AYHBvfsjVYSH4d+KFf7IPYvKdwhYMTwK4ESKrjDhrq5aXNwtPJPApRlscc7I8U1dHFPsx0
aoWaAyZgffj6S5a+arVjtJEZzyR2TLcGCjSnnCwNDsXz0GqKz4CfDvGHekQWjkQdH0A2QyHnh4r2
kLpm48CV37KcinxYSe75nXa7O2FOVxXw7WUFROcDAw9wV9Df+ZJViDUn8WQ/grRCnlUE22ZwES3G
PmpOuw5PmpDs4FbN0z51QPhMtX3UE5GjtVM4BECl84X0z/tbVQhpYZUby6Q61V0XT2cZCSv3Qz6P
F9X3l0My8727ciLbDNl5kCr/rtaA5VwiLFnz0hCerqqo337L9RWrchwNAd3PeivU7fmhFWVpPyaN
lgh9gSW9fFx0/dYronvE4DhPkL9I7DOuV7dVFKYaqrTn4eT5Fx4Bp9H5+YJFVOUYmal5oXnyR99/
KVDrP3qvTr0LRPUqMVlfq9Z+lvkjKK+i0kiAo3b2ZbdoU9uN8Xk5XIHxMlzDyNvRbbtg6TkVwrFv
2hqkSkzxxcANsC7M/u2TiP1Oh47uk4GzReBLG/zX7PXP9kHzcHsndti2RKLAPv2nJvyAEIbviI01
IrGkrDCLySut4pZjaUyMRpTwxl3pAZEMbbIfFU8V2OhPkk793l7ctPk=
`protect end_protected
