-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WLFa7YGthChyih2g6gb7N/ceb63VCGNcP7XkBswXr6UGY/YF1wVKgk5xTBWLzhJvCm7LGAwLmIKX
YFbn4ACwfJqAeKMtbzHcJ9aE50UNkU9bFWxPEN7OSY1Q+K6MdLiXMxNOxEwYulvTgE+aimnEOn7+
2IRKcBRiN/ajVR1U8k4MB9sKPqRYTeNPRfo54ec/lpQWSfegL91s6LhwKivZ3BmC/hZqAP6X6XCP
PiTUFztvu1gPN/4HRlr3/vHQmBJEFwgubgs9JzRnqaLv6ijm1ZCfmZ2Ltfk1S2DKhM6JxchJVxLh
9grl3ow61LWPyPZJCg7Aa8/39JR+2xCBddc7Ng==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13568)
`protect data_block
e+FGZP2xsJAr14/p9oupt1SAMS55lLcIWUw4WoNHTt1ZqdUpLGYGyPeBGYT6G4c6oNVKB1wuO/dK
iIPWEmA2xQrcZpfMHwBdYC8cn8ft6WzldhxU+gpOPlKgh3bpKvSkZkrhmIxfANU4gFzjpZ8jk+rA
L67MSbXmdXYNg6ZP1iAneXRNL74lBlZdqArNvvoYXV+mhRluSoL5FauawyoRbTLmQUP6VTuB3m/Z
l8AT4cFsNoxu+9Y3ugOQcelmSwm9/WSeDwpCenJtmAGxRlgJYh3mp49dPhIaKZehww4xXgZCutlc
1Rv1VveY3bhww+iDiaFPe8XwUHyOgOgEisK5EWy5dvMOnThLk9f7s38xGDtGYDyRpj2j9l68YOJp
k33lSUa0TGZBd4ZpO1OfFzjLGLjHudaD5+iUTXwcsnHC6NmpKZ2IgxWfx3sKFZpffBrFhUo0qB/n
MU4FTcgUqS/Fd06PtGs0twOea+QhkrP0tRQB5P4qiUeg5ZsFhqCifYfHDwGWT1n7MjzDWMKcre7C
3WA5rHj4mn1WmGtWv/b4rDrAOM1Oxpi8mSKksH2eU9REl9gZ7QZtcGru7FSkMnWbvt/tpdiolpFI
wvVdtlDZaE0fbLiZbT2P0comeDxRFU5aF11flLEcx57hDF5VY26SFQMuILd2QQUCmbETJKoMh/W0
5wOtW8AJ+93YyIkx0UBirIQxIgSu4sK9BdIjX3PXwmNfz/2N4TsofNsJZq3l9dPIpawFXiAe9VEN
K+SRNp867iXLTnHk240/8HDM4Yuv+did/aX++Ht24jXW/r5NL/xSNOaFgt3D65e9eryYsb7tYJJk
C6DeB7VID3S8MG2cGaiwQoinP/OnNvmg7JeUXsmpymB752nM181SZjAx2iZgMRRXnE41n3AZCEI2
UPCbvh8NvQwjSYjXPOMupHwwIkZlcg5aDmzvOsoeo6CESsIeu1oDOu+fxtOBQdfWtAhNYrPXAkcE
UfBYjXhFBrTMQIGPshDSGYilB9XBRRt/l4R5J5qmdRdCteTR7kA+xdcW/wzWTeAoa+GiSG6QTxlR
WERthAQJSWbwdnae9JxWRkM9w+eS5iH8c+R5w4zNbHei2DqUE7ZKiOCynsRxIPmTUTKiVQ1OFspg
hK1SKMo9ajwBoCEVr7+0diRsvaH9WX4puHD4XvyzdHa8JMMrYtY2sCc+/EMAPf1IdAtomjUPajj3
oyHMcz18VrN86+M8XhncqAN3aGnyTbwRDH2X/utdbzrYbCsf6tE2YqsNL0mfktj092IZarYjI9Gt
un3IHz7dnSjc+G0CjpWM+R47nk3GcqRMMAOC1enB1NPpPfbm7mn4aEao0xGjnlQlWKM1K/P1gqPi
9bhVdSrgCCbKJWfuLWmpcl9d3IsOedJ3gpgMlAT3PGMYv4Z6lIyxbuKAcuUywN+mGADnZETmNrPj
r8+q22lkwetUaY02dDHBq23T4T90hIfSg2WkKBP517Z43dqcPWrARyTeTICy4c5Rc6DilPj0BUe6
wpPZUxCVrvWvg0rrudYLSm5x9N9ERaUmxlQUR7DJ5qr/TCbTyKbSbTm9OVbuH/3KCcWVMegwBRyy
7rnIs546fzwuW8lOw7LTgPJXo/DK1lFUVLXmnPdz6hLb4Ff4hbiLTw8+9l6IT1uuL+3mTi6GddQ5
C0ePbgKnpaW9QYXFQXeoV7eny+pV/WHcCsvnU9LW7qNvntLbAV2RmTWqTLU57mT2mvHeYm9n6u3B
R08CRGCMKJTP9fDT9U0XSSxT7Q12ESDuE6Psu0KgZAUUMaFp9TfcndJ39l+ZMTQR1MFhYS6jW2bm
iKW1Cw8DjFl5LyIPbPhGedkFsDHnDpJOP0YTp48tpmrk7DcBsjFOeKUqo+Vlpzd1uYQH9BvXdN31
lF3KddcDbfKSsLHisFMgk1axKsIjMiOabHG4Zi4DqJkJT2GMQmsOz+LzIbgilkRWeg3lBSl5xBAK
9kFMqvmshIKoIkvcJJqBpoLLverWOMDxPyQ6Z8WkP2kbpKywrtHioWJdxF4lNpm0vOR0zLPjbUNa
eap8TRo+NJV57U2msnB2RhDZQyjjs84ddPhreKpW/ZjPnGaJLkMC5hTbQxelasnJCq0AQNiVhX4G
qHrPrzI/OEzlXPiJsCa188yIlTvWu0QUVrO8RgdLkqadLotdj06FFhCQBEy8fzVjUSN5ff5Z4Ep+
+0N6iwas8H+4tcxZdGlftPdeJLoklDC0resFzHW8CiraObbHNKIxgQcJNaiwqq2a1rb69DnGVN37
0yOjQ7SYPeloTtsDKosH7YbZl/BVCnURVjw03qdH8oGU95JFByQP1C2m5yYhVI0PfbUEddQpdLjB
8KrTVQMpo6YZIoC2OiaqRZF7DgPEnZNS6ZqeV/xHdPsGGAJ5ieQUEn01SJgjB7DP6M7fDoNCCNus
xwv8f/ADsTK14UldJ/c0hA9arIf2+XIaUoKpWdVUGF7ZG5a1VPjfvWNcoTGvsb0ai1RYbJxBdzfH
ix5w4IsOoVFwrT3J3ulo0opMu5g/Td0i2Zlj6IJs3ilCb2y1gV0ULx4sN35fxk6hzduLoy/1uV77
mv38mXvdMGzP/p9nsySOfJfOHDXIvkZn7E+jpq4851QphXLI7hL1N6I7ZKhn4AM/dJe3Dij0nJEj
xEKH+nz57/6T6FDDVrC+4yCe1ezMsDECxnxgUKZM+6WDIiP/XVrKi4okszaaB6xLyYk9HgBvSlRa
65UFUXM3rvPYfbApBrlX9ra9nMBogURAJ+HQfwzJtOEKxY74BA2L9FHp8OPuAmlSqXyCR6bOFpZn
uoSDNc2IlmZEX2aRRId7lJ9GvhM1Qzm4AhiF+mqZlDL/XKxqxOcjQh4WXI9Sk3Zs2EdaAsZ0DVIr
ctX2pfH5DYgWt8o/FRVJ+As5+GWAPT6epzKYY38r0C7nj90k+hlbzVmnrdkT1XE+r1a0eNQ66sxP
rjex8FTiZh2aQjUWF/ilLO7X4IHAX2hVPbiA6A3uaC8wpSIKrj6J7XW4jc5Bzh1Qe9QSI5rdHaic
MA71qqMABxmBLt3n4I+o9bldPAy5nKwwiUdhNhnbTljRglVRqijl62B3r2ZIbmmT/FVd3D9zGa6A
vdECE7R4f9rwW19J/Od2VBCrIuA8D8LKthvURAvfOGslCMcxwTCYD2F8O9KSkqAJY5HFD5Fz2G5E
r5hrIhkgCnEqZrBatYrLTERPGzeUtUGxIwxc+cUBwnlaxZVWxa6Czm+gwD53G+MbEyxZLzePUDDM
P7z3c/gVNEv/0dS5eiWc2oiW8hVonUWU8lVbYL/BaT0yL43EsawT2IRkMiTvx69BkXWHzxo3Tq4M
173vJl1pCULDqumLEej3uf2mD6QnDE0jEjGjvreaJT5rCuS0RycCNVeY9r5gcbh3LWU71YHLjOg+
sb+5FKhnviJ/4PjCyRnUJOrvaJJWMO01LW/ePLeBDnc4HbA5sAZBgy7/271InFOnxr7CPGAcRBkG
3I8T2yMRRQKm9MtOry1LUHx3iGGbqAaMdC9dkMZza19Ju8Q/seUKX2XZ3AP6+/wObVhOXDmEBH2Y
S5X8FslW2p8uayFLkVkq68iRIwtZBCoNj47BmV/H3qkQElxH2gM1ghQbiKKGH1ulctHAY/DaWiiZ
+9AI09RKkkjZUULWmUDCdtUtldhYmPmh1PRs1Wll+FOn2/ugJR1wxGUjrufUrYajKS+BW/QMPtja
jB/dFf2Dnk0SyYZAVfzx9mYza8OrHe2A5I3FTI+9OhELco9BjPhklXBDHuyEApm9mujdHDaWWCYe
t2rfCnFgTG07fWpICkeyXIYnDpeN4+ny+qjpCjP+eSDJg3jExOMgZNSAw+h8fh+dnyN20uRTW8Cq
yFlaihALkGOUdIy3OvECMS6spwamjPScw79+JEoE8to29tkF2hJZSNJxgNLi3YKgRE3+qcdzRaz0
618ZMC169Dwonbz7RZuBRRw9IubDr94ZoP7ipFn7TMA0mx3CJyIjRfYhJE6AhvJ+gEEGKUHMHY60
RSS/1T3maYdAkhqIExXQBCrAn5wMixt0t3/3eG7q17pWHBS4fxH4wC0DP9T2F9DQdXA39F2GjrWE
d5fSXr3e2PguLOe6MXROi6FSN5abQHrw8YIULhDfEOj8neQX/69IOSXH8AbVsKLdJccV9lj/M52T
wUoulhvYE56GQL9w//N/1h8DfQffWaRt/nIZqGrK/PWuOzXGtCw0iYKAbDMwRXV6/f1yhMZKCLgu
Q5K6yIOaB0fnRRmGDsKcczQDS9rB7ldR2JZzGyIKIz5CZ4f3qrLBMwdxDgva15jIV0tBJyVkTDCZ
VhUnUyiczmTBBl7W6loTQ0LaXFvFbEBFcROaOOg9gqnON6JpDltMaJFFcRoTs52jZPzl17a+3euF
SvE3d3bYFcMrvhq/vdQStkPgpn+c/uSRRrhkr7lF6T4TxEG9mWicP4a2psWYmRRskVyczQN+UmOU
LfYwYJJnFY1ld8XOEvE4McAi9LQIynr+NJkCzOnh/43LtbPv0fu6oJ8KcaUn3dp3pHAU83krGxfz
aqoG1dgqwm04yK+Q6+VKV0ltSwfXoJ5ePsCu+KgCcST/ZZ4t62fBMyed/0PsGTANyt9bBQspQhM0
W5iCwy7GfvkXQ8mml2MrrY3F/TlApogOmmRxh11tsrccfJplOfpTjsfkKtOEhFg47k2yxBYq3P3i
1mDFd/ioaXhiZmTKXap+H90xouUP+/UA3jSSXkykJBsQiy22K6DCf/tbuRMJ4YmE/tRiizOjxx8P
uK5rpAvnCnwlZlvlL41PP237XmKzSm3hVY9V+d+8kQblFI8BCBbOqGh3VxAuhxr/PtbO0KUe+1ne
/52IO6cevXLzjONJ5p3ozjlM47vXRY4dqTyIrsxgM6Rj56dkrISs7n1d0hohhApcSakdtXHXir2P
ItdlsXeLIperpGRrDxILA7oPybrSEenzYANGOvLhW/6X88T5YzCEQ6QW2D0U4C52q5xmI8PDIi/T
hKirNR5bElRQZvxxU2lD+xxwQ+kW2B1RGpMew+yEZbbs3Z4viR98OCriWYVRT2XDGPsihGC+Em7I
6nB3RxwG0L2RxguiKvDvvMSs4H7CYIAqumRilQGfWAIdrHiSN/TeQuCkMWXGTpw23mWaTv6nrvCC
KV2gqIOIAWrEjU8Dvg71yTkpgDZjWlnUP3rouIFWtsjccYek1Qau24lTJwS9CatnjUE+9I+cSmAh
egaQkZZuSB9POwLcuDrGDxKBr4WvJg9Ef580znfcHbnvWSjgVyeRASmt/G/5NipvPGmn2GFSH7DQ
PB+SrdWiyT9Ll49RMJDYg5Qk79nFKbVBT3VIPF9FrOwFh/5So0hI1A6+tEXjSyXJJn+T++LoDrk1
JNIuJUrrndcS0fDDYaY89X1T4yGGaJ7D7imnW87rsIelPHCvSy+dmBkC6rt4edqte/bvSNadN8LR
xF/cyDpN9YmbObdlMiNYWkf5ltNRRp2Os9U2j8Rvjl/bVICFz2zWXApcyNJp2A3ubSNX1BEQ4RlF
tFbIi7lIe2/mJO/p4yVIq2KM1HuLwAM2WNK6yo57Gbkdhd8HDoaPSgDqNp5IdpUVbipcHjXn78ez
WZUopL/hF9B/nFmAUwtZIUjZjx6kr/0zNVlHbPFpZycFVQDhuZ/o3y708O7ObtyOqLAIhMrm+RFP
G06h2EWBfFt9P+2f1pvbF2BTnvlLhRz1hs4KEN4ODgKi+KovL6lmounjE0SZ+ZLCs30dw+upPhYd
XSqMn0wFSHdNnp0azizEvxfYKDlsJRzEqxkCJ74pafVRINcFlEe1o+xDjgz5Ja7vrUru2hsHeeS4
RseuGm20DKsSD8yC37IETbL/RxKtk3sMtU+w7QIs+v6PsU+1ygcbGSfwMm1MTLZo28tlrUsgLqX0
nZtSpXjUNJ3fJzrLa86W9Av3onSE7XGAyXgCrDg/F6qLxlhiO/IJCeNDC3d/2Asm5xEEOQtzGX17
eDcWJX4EiRoUSqS/sm1RBAKIE24SeWFoElXNhTWxbYIlJOGVPkQNKUv1GYKqJvbVNPPYp634l6YS
Y+u/qu3L++CXEHC6svocAdQsaxpUMuNog3aDii0+ID6wWESMeNws7J9/LXEeV/6FymzBkGdiIncW
kxmaGCjmNNcEZZ9GR7wNJo69dfW5P49ou6xMLu/YZsAPuRIT00CNbYFEK00W2nJ2gvjYa5XomStQ
FEzXBAdII9JB+xMQIVZhNV6vzdyh9bzD/R/vHH7n30nNmCnmbW+90hy90ScdS6OZqOb8v6YY8ZD6
nZ21OdMq3/4AVqn92z/uCQfc+R0lfLoEubSfkHhPFn5t3NsdbtQVfejTzduAMZDWdmqrEswYZ7hJ
lhmrv1trCM3Q84/Pf/9CxceVyAtfc2v92/rv/DJh9jet6E2B0XiEKbDAERcaLWFOdz2agO/rr01P
Q/MRGXSfk6P0hnmFnl+d/Qdo9+p4eutJBKpZhAW5vgsubkUTuu6nEZxj4/LuhXc5De3Iqv1VXmOF
3dcRUNgLJGXUlz5RIPXF8KGKVpdz89DtLReP564xuf20FmxDN1hs9STUimzwSwLj1J4+dm6wIXwu
6zO5DarBNNACsA3IQt3EQ1rZlFHfn+YrRmoQci1lUsHqQgNCcxE8iWldRipI2CUk+NL1KGzloS2E
vhypp8ZK/Bcp8QrprPNtc45HHQgLiVoJFxrc9mmkax+hAehJuM9LUlNH2ExEmeUZrQJP68gxlsfZ
6QKQ4EWdz82T1Px3LZSs9Kx2OSaIwBjzZDxnCyaSMz5Zl2blf1s5SKmQFx1vqycaNzYGX4V0glLA
GB4CLwoSz6i4C6ohpEQl25YrGqd695B/eETeFxLSJbcgEi/qUrwJIx8G27NAJPFG9RfLUU1fAvjc
kPLEOF3B3TDnj50p4dup6BXPhMKeoZnzoeKlZ+zI21jYW+huCqimwaqq3mUHgpoqAQxe2UbzYNPc
xNC+H/bYskzMR6qfzQ8Rvp6mxR35Kr6SPHFfQ8YCTWrmXy6hst6k2Gzv2ShQSXdK74ba3xeuJ2Eb
bI+b7i3GTW4lGXa8Uvz6hrkHZ2ll/EXo1imD2GVZXVWpgYKTANUY2x2m3caRReBOfimogIM/pCFA
bZ+5Bq0Qp0BBl/Gdw0NVw+5kYyPBa2REjms1ovDbHns1pKgbmzM0vV3FFadWjfl7nBJ8Pzn7hAhg
51EiMgbZDDSaJJcT7nwIUOG49IvFK33WbhDoVrHNml0x1VZH26ABAIR33/wrp3FQUrRhFD1G+RD0
fcjvcISZXnC9uZFrdQgpWx11VVjhI3yMl32fM7TPgX3XHMLe5DmtaXc3feNdY6h69MF25uX69w7K
QBWg8j3W5o+BT3ZCP+3IxFAGguF+RJzreI7tpmDXsKdwmHXShrO8PY32f693jshunnPB6FH0rFbu
o22d9hnyGwuulSDTKaTAgYzf7IF5z14qa/oRm7JRzOotfCHjx/7FNAmefxybM3kx+wh051ipEMed
giPC7zMm61Rsz7RdRQVaFr2M/ha+v7gIj9Kq/XXEkQ0VxufWTpz33ViQ3Al9K3YYBi1l0pWIcblq
dHB+/T393o4WIBtbKdRJJIdYd6aSz1u/9VmspI3HaIjh3zj7Rm/lcRam0MSjwj77p6jkgS9UEweO
3VKHjV3+Pg98tGB3TOTovF2X+4KmFmC8AHO9OU8Bm7Zv1nL5Xiroxq3r67NTAh/PVvLVPWSudUCf
EWM3PW7EZh9JqtlTuT2mMRnrnigwUm9oMDI97rqIW6iJjmk4FfyskFtj39pyiimk6qfwCRU//Z5s
lvRp4j2/C6Zj2wlztkZtzEq5mRXvZWbGVLrOtkz/0gxdNf/eDgpBoTxKWBiJzIyliv3JhiumHyQB
1u2PLP8ctYkgeKN0qhcBKMdRLTdz3ryVOqCU7HL5ZCDMpN/V4Cd5ZaQO0YJsY2iQVmdPpaLonorw
2QTJMzkiYsJ5QRfLI6B+LfkqcdLhk+5HvYYiVGxngE7Dq5jeRFA6U1P0E4PmZcOvV5+Qe0srVx0b
MG8j6bgGKTlPgkSqDnK950uFegdZ2aUDi8hcURZV+fW+t5H3bpHWiwcDwMZGlKX4Igdf/dEbTl3k
KSz5OVvh44ARAfrOA3qBOJzxj42lPTksZtpFIbcQxRlwKhlIwRc6h03Y0m/Ch+lRvbcvkp+KIMFJ
7Wji6oJKwpORxa2ls8mvnl7jzPh/u2xhss3FK6aJrWpyFGMJncEcP5AhD+qKkdnmdZDiFt5vEs4T
gx15qU9bc16KZGlOiBP+crSibuo3yanJXlGuLJX5KiCygb3mrsBfpu+EVFlxxH2WeI4EdNUHdT8l
6DHDPoTGU0FqmzpuFXbmprz+kl/V6Uogwz/GHPWKWhuKdQwy+sXWSHb1/u6AROgKNXrQ6TJ7QaYj
oWO36xIgbkUhqFwvi7+e72vBwVA22+92imcrSaq08ACD9jomchPJLH4Mc2QyrnOfjzuLfH4/Tmyw
yMmxgwjzMNbwfBM2RaVRVt6FRLyvVZJJlhtt5SO94Rjcq/OU+daJATDUYNYK1PSEslo5O7sjT/qf
PRA7pViM8jPaORUEC4uE41RBhS9MJydJJfYkXVffMyJleT0TL5b+TndmcpH1a5iSYPjmDp/NLrnV
TOOJd3JWp6J9niNw0vxubQChA8Juy3w0qfWxZChbKk4D5YEDjNSP90z8eyngagRrLXnDtBUU8y1v
aSB9xmmNC6wQciMc2xz7xIEV/hZNo1VWLH2j9+72zZgbrhelL6R9BR8MI6kfM1hajMxpvqEekh2K
R/zL6yFN9gsWIekFPYiWWlOGmDMwu9ihZAJAGShgzPZaeMaW6oxOo0tkZNHHDiqarCGlJHbhxx5Z
kGX5spTlLB8u+ABMHikpizSsd9LpbEIS/5TOoaG+Req9MrZFwj94iojC/9brHR/iOeeX6Wsxp8RJ
00vCEgLSON9v1CdTF3pZCSuHl9pMcTMkoMlCxEgL9bSvB2lq3FtjNDGmX/QJSmkUiweAXRJyoNPu
XHi+lLp6nD7p33wZaQq0Y448uwTwhTs7VlmHmQ1CGdbQyjn/2rlDeGYoelJ0emrYxfX2623FCI5v
rhbu4fh9Etkvo0YGr0b35XAmMq7amvKZqH5GVFbeq+tF1kXOd4HV+zWmB30RlyBLcOpazA2eu6qS
P7shAzaJs8OM+fF1PrnbiGhPeBom9LTzVfHY8wmZ32t7t2YnK+bvG4NjM/J7DB7ibJ6H5k/RowR0
EL4WkInaNnAfBB8rtJetPRKN7wz9tJSygxgs9qVPBlCnzOalO4nVm7jvxt9bk+Rhyh4vkVXa2iM9
cUzlbKuhjt+SqvG+7lGkOePQU10WlQYDhWZxFlbsKQPBHAFC0AzIO/vG8to61z5s363q9/qiR+qE
x06z3zRETyimRMvgDETQk6iOu5M3KW93K+Bs2cS4o2N8vNdp4RM9V3W+m885vaWrC+oZTqjkUFaj
7MxUtknzA2otHZLp/45VmIyyzkq4JEZ30I8sMRLXcn9H/ZRiMFmg8Xb+nMok5fhSufQVHqG2Dpyl
upbpTwvw1oz7e7POC/u/xQ1aatiIokuSNnpAJ4BbsWklEUspPHq86X1X9n8Q4Lnbgd9h5LiU6yCx
mjbHqyA2AQr3RwN/Z1kAeq4zclzs+HHX23YcOYmyPuTkSJ10CXCE1emA2Hg+73VYVQW35iALW3eg
xvxArvuVmRMprVmfcddhNusyyGQz6kR4/vUqIyQet8iDlfklMaBrWbhQFuljYn54Fwx/B8EaVuQ8
a9NCccoNWMEUrt8gaQ8z6p2wPVtxKTonsvM1blYp5Lw2edMuTvUIVkzSLDm1ZZeA6MvcIEPX/QYc
Cby+2tnAAbhQcVvvgsEVVwah9OxNKdHJHGNSGJyFDUD8JDLvrSjWjusDH3EcYyKR8NOxQXc8BsoA
ebERLiEj+IyrilAWveTrEtRPApDonoD2hrPAMYYTMuiVbQs7DTdSYzPiLsYr4GCrAz32SEa6NpQe
PQ/96A/4O6Fy16/rIt4lEvvXkGiI8jbdZ2s2Z8NEvyIxsBr8SIdD1jqaDHUQCEF6jQp8YslJKgUM
ayrO+/Mh03RUhA/V+iVOeuG6Dq/xIyO45udLi/INoWhhgTl2N2FCn3jifut7PXJ4H3BpARiImC4z
2Os1R+GbAlhGdJcpA9CcavgPDMgjJZcElXJK8nGmc5OKFWb1qXTimaZB2w9+9K8QVd9m7NW/mo8m
UyHOy8lVZ2qbAHde9nfVrpF00MLZm6hWYifW/zLFRjF2STjqm7DoDX6FCq14lpzqEDKrmClx+4jG
f7MaZo1T9OYWDgPtDWlQygQkPUL2k4wYCw/LAnAtzjW+jAD/SWMKju/64lEKGifiDKciyQGJDa2W
YGn0QqeTHW3QUBjBKIvyJXaTwdoszDX8bluHyRos9s58y+zTnQ6RNI8OYMK7qnXnXqonYUaOVJTZ
egZeZpG+8T5g9zA2PkIUBOt3ozE6A4hCguHLchRwZI5adcLpDfjvEeFhwVaE4SxpJwDn39bnAzXT
xe3JoLzxl22MOvgo8BupTPpoOPqeGRz4VI4PN0QBrwkXIVOEHRE/11ga4hdHqOYS9eWMji9rw2mz
SAKaeRA1nGzr3XZr3CuTFGF5IDd00PrEwhDxiyj3CMTvIPsoug7iLQcTOjajYhVh7BgDB7kwHys0
fLtvt9wuGBG64GwGzn4n+98cExY6bWxIX4mJ+ZvcpAgkWNzt7dFB6PRzhc+TKqkuQFQy74ALeDQv
K/NA16oukeSTX2+qcHbHl65oTm6ke5JRHK8Jm/PLqhYV2L8af9JpzEROWwbI1HrBFSSEzFhZdjwX
qOegaT8tN/cKFrujs7saEozRUB2qoMgCTFg3OwVipieckRwKIyj3VP3t0fGS82xcdopOitYUfRar
h1yik/9V+ton1TF+SWU0jM4ASYt3F3GKWOmvoCOk7MbEeId8HoRAMP7oDV2D9tlyDW81uQxUO27E
VwuFkoWHxwEtIwLOKs68pwyJRZ4IGYn3y2h2MR7TsFoEOcIjPTI74LK7chbIPDA3YM3xT0FXfOnU
ig8GgULZlfVd6bcrxDxDlFW61lItqvPE50w3n02Riv7ZHHRMzSjD40Wlp5To1px5ZEnfgtbTcGJT
jgzmlJKFSBBJwL9P1pO5NlCmPBVFJaEt0aG5as2v2JwehTdmNbHJUs6oV7OB94qwhU1o9sj4QZUo
NG3+gOHNwquzUfvo+P+EVLYxN/JUkkC5D3TSX4Ds3vWkX2dSO1gQH3SVIOQLokBiOdResp7z0KUg
x3kFuSeUNA28QjCyCAk5hq3QS/SRdMKUCVKFgwSYsuEXGL8GloZAtGxWcOs2YAhphko3nmZMQtFZ
WDddVlmsRLHfq1jWCndGUCNHvn3yOJV9DVys5rWYRsHiybfUI6CxrI/CiAtEZvAj+/6MWSA4bonS
Vs5CEd+Xbe+2N2eKrdWSgDs/CrxiQUajSpD6iLODFluB4vNmDtLoI61aXVjtk9axfCZljjPv+PHp
yNW+S1DeL/lJNUrZhRRVYrUOwLpQCJMQyxBXxv6HUovGbPFrPXzvWUgpJwkxUZ1BTr+4jj28zqZ8
gTDBLqaYhIZaNsWqC92SafvQFqvFFn9PPbs6H5hPzhKTS0gC43ST2c53qdQ6jP7MVTRazIYc/dDL
qnSh3Qs+EorSCaEKX5ASd4VAzy2O0BR9h5kFPqRs8g90UTH2nKV2pf+XLqbyGOyQYrGtPakcOAfQ
U5n3lyQSn6hv6V+96JCW92ezkwpmHMpyik4PA/A5v8I0jgWCaNHbj/T+blJZemKnIinSag87rW47
F6imLb+0rWNjZzOKJMw9bzmUQiKG4y66+NmpAQeuEifJjdmCklhjf90ska0siIrkpRJDsTMSiAm0
2fYco4L4KNHXh6IC6LGe9Pj7mhcrmsn0rre6AwYqMiDvJCxGE8lVs8ocuMi54ux7ZeU2CWvOKhKy
tzm/HDDz/shZ+i++R6nc0Ym+LWm9CEIOXtqMedSc+JgO9hNwVZqdHcrEbBol4y7bvm2JgqhIhDK6
IwKxdbam/HsDwFvJExLr7xBI1Xvs/hmcAy+B4VX6UQ9lWX49N0Lh2g09/NSS/va3TZI+j/itCxrt
SvTQisDAJTt1I4tTc2EsR4jeCGehOPnN9Y8IHaJaoB1mJc9/ftEiDj3q1ViLhNkGGe/BRqjKn7+n
ZXIHrSIGZL74/7gls0D0i4DkHsAQSU7jqPAluFCSu7ddk0jlBlzrEo1SvpwHzf7DIHaIbUzSgPD0
dj3o7XUDEYv4yEh/q6alugcaqDAQoPwMfkDkfGZP0h80VtmRyDISQUvjkbzCRas0Z0wcQe0j9OYu
JeDZuCRtOV2u/dBiFdhvXWxYr4qe+xpW6T4bst6CdT6eG5ujI+HLrSrpprpo7auLZ+roQmgJT7Mu
48pbGgcSdn0AiJ6GABmla8MowbPw6MFi8Iybm3b5jswJ0bc3utQu1oVlDxoxTJd6EBxBq2U5V+Kg
FxQFvQQwt9TlyZj/Wgl4WkRfBENr/JEYLj5SUur4Gjck5sUPha/UyTFA+fZCS27fjA9F9kinQwQZ
Abo88fhVu2OeZPfI1gq2CSgCcCoOveXGFa5Vuglsjo+4MPYk5pFVFUf18BP2JSYCnR8e3IA+DMX9
o+c6pes7SKeih6n9Lu9XwDFOULff1rKFQ6uiBhlDEQi1J3VK2yV6G79nHP/MYt672MqoieQM1gR6
6xSRYCprf9pEhLXytnZjDkNS0+9kmPGHuyWytIRLLxaqfRZrnmbS6ZfFsbk43wS5R7XrcOaEcHBD
AAGFTiKFyWgtL9TKtzKybOTi6GD3/nAc4qNwbU0A56z/ANQzvmDNyciINDNoGZKrbWX71iLbVF+x
FG1UI4NAU7OiY8ZcoGbEdHwsdlef2OjOLtXWVp9CK0HGuEniRoOAH1rtfw66MaO0fy7/Qh9uwHHg
zam2PeYCg+fAMRynwnT7NyZdOVpYCrtfaE+2UqEan/emx2ZO8e/GG6BRGbHvSjS8/xf3yv/mwJif
3wvZj/KyctxplVpdYTQoa2yTOe5F65C91S7T25JoRFRrgBFxnx5XlONWm11Bi+ULR2OOzW5D9s3Z
chWuIAmr72k0VEZkLlHZI+MekpyJZZj5xOEDlcbOUTR3ox9mhIdCtMK7oi7jkDLFMi4fM6uus3zp
qeQiqLNr6GZjmhKyioQEPUOrSmHLxyc3GjdVvVopfFNYmTuTTUnyQLi0eKVioWDtdBLRA6Aos6An
xq9WNvWw9Ne8QzscbhMxMsWtic7bi44xH/GWbaMkpKpHg1FwpT1HDciyZcwBjKF2MpgHnRG4esQA
nqtKAGjQleKRTOQ8P2fmdDo/eUhHNymtGpMl7Nrdow7Pu7BKSLon9ATxht1n9u2MbvRm7k7BLJ+E
me5rtxQ2i9rSIrKQOia/s9YhY0eVdYq3YPJz1i4yFNKik04VdSBsKaaqxVdyL9MPqqEbwK8OLxjH
DGPJg7az3eolBUx34kxQOU/kaczstNFbVmJ9MaQndl3lCmEH3kpoSS6+7FZZr9XmkFBOuw2QYrR+
5+hMRo8b97QgkHmY459gc1Xh9kRO5CnexCeNWCb1+RG5s06ycoGkj1u6gYsF+EctxjoRaWj7DSry
zuSqzJtjbtXqaLsBMPTn27PiAnH3mHw60DQqySHEvZxHm+mID9IXIk+tVJJVvWB8g49BeGcw5xQU
e+9ICZMiOQte5DAjYrYqKsfyIGHAChP88gj93XeHvvitFcohkony439N/Say0aEQcTuOR8iZ8Pmd
VpSritZd//iydobtPwgoforTSh310Q2KedqW2IJ4r1RssT5eifAWNhA+LJztbNnvBvXjdxTmirjb
YzBrUB0X/7YUV+AUXLXSn247JIKpJymi3t8oZeU6JXRCMO4se3XlCHST9aRnOKXy1vcLn4uZsa8l
Zoa6XvMMtzgcuDtzKbfIVLY5a9UV9OSs8h2X4ff5tZSxku24B1QjZMwtnHotYN0dyKKk3cdinVGW
WY0dN58384YiIEsRmX7/+fHQcfWfSN4RfQX8RG8LCvFn6LhmD8Qx/OvhFc+AdZXnoq612WAavFIF
C0wE5pZkyb4MpDlP8tIuj6+Tr0ioe6O590wTJSEESDX+o5udXlWtF9Q8Q0lP2zQSptNylGMQizr6
XoUK6x/aBzrE1YZ2eh0yGRnGmIIPKy4IQVpG6e8+dMdsYGSY/oJYWDT2dee6CJ3k6y5e6Wt/+D7p
itZ8FoMlgq1+GaEgz2XgKiYz3K6SA9ZnMvaan/C87R92vfTlW12ATNc9bApnzWqWO39tD2tMQ/Bz
Di5h13DdDYnpFgYTGQQi/v/uvqDS8JcUdnv1udwSSkCNsFkSdbRiSfAVKXz36WoCNFFNdlC3XUXt
l+8qa4uKnk8uuJRciwXQfNOE4m4pOPj+jknBEDIpQqH8hD8HsXlb91dkAwy6dwuv8UGR3Oq937IT
jG9GwFEgKGQIIxHD9pNjFFieozBE4euR4XlTdQ2bY89KwlsbpJKUqzawfrZULBFyU4j6TmRvISwK
hw+5dubiXcvea+/qso5BaNblCftNLHNjL90a8jHs5gv/DZlX3QeU3ige1++m9gIPvhM3D3bz0nKY
26acWTKO6r8NR/9/SFpxhLMZqQzNkB93NbaVJUXnieHo9Qb+WwI0Cq++X44NDt03cowv5TDN/SFE
V8YBZw8MKEDwRXWC72m+B7SBz6m4fNlfMJHYyGDDjMrrzs59ZW+4e/xXlRft5AKKA4I7bSVfwm1T
T9wVWN7ZH5RirAkxbMivdoJvag5e7M7UPR74enhFB6lbsYXUFfGMqmb3PCfyHWPRqGaogY5frmQz
SuxadBU6VA0713RzJPO1ruEc9yg9LKVRrLEx21KiH1ZCJBurfD3kca/FnUoLqLmqhBLeQJ4vidR5
/gBc+eHGgOhB81Xre86AQQK2tiplXPhzzxmTuYlxMD7i38C5Aplh9zgc4A5VM2JaEOmbkQpyCqLk
KGH/g7QXM2cSEwsB4C95HT9CJGtLft3qXtx50Iflr+QU1NFwk5fFcjsWnmEyfZwyekEXnZcw3qJX
gVItiexx0yv8FNj8x2vMJRg7BY9vilHGYJzWyy5g5bWjcJksJBr+yrZ6wN0O34g2B/f7Fh/XGRtV
S8YLp8xZ7NFJ7buHvdZaikDQyg4MJ3D10Vzb2r0cPrU9fnQLIX9s/SPLvOSQI3PbR8cnAayld0PX
mQAEVL3vMnyAZNQdtWT54kiaAFeSiGxr6pdbGHmo6Pr7nkQgO9oqcbkSB6MdW3k0mk28Un0vWSs2
y2TjIaBebwKkUkpHMc/nlSIIHObQ9YgSatsvAiTy3Z8bD2Eop2cHnfaa2Rx1TTUAnybi/6594J8D
/hsGp3XyAsoxp+9W68rhaWqfJUqMCKUWNxcN9Jf6hT9YfNlxrC6to8OavzM155u9aXYj9cnOZ1Gk
gByzbwN/8bzdNmbHeLW9jqV/acdJsl8BF4Yq7+/X+W+JSZr3FMjV8Sbf5fLJupyVn3IuAOlHkdly
mwBsUYRSD5qNHLG4S0T6DX5/2I3k7i5D20xADYDnAIfykRv2ZL2sg6tKaiUh0kiCv6Ct418kCRYz
f7Rw4BIyvs6wJU34/RUea5Lm9dSJ6hUn29bDDX/5YmV2XoKiZI1OBFtpPB9cusTvRWXrVXKmCtnQ
HPIH8TKKBTMMYeyEzvV4p5ncPge2EyMenDthDcEIR1gyF42/BWaKcTRi3d1IeNdniglrd7hDZ6vg
VoCChx6K7ywHK3p7MnZftQ133KDuImkT2heMmhPdwmdCZW6Zc5OegTCi6QI3dS6XlopnzRe+8NFM
uQ+8XOJeBghAK/WITCwxkBTywQkN/722AJmJbLuEYkd5HEtDArPbR9MKf1uBkIgSVkQanXwx7oKO
DpDONW4+DHWR33Lgo16c6T1QX+u5Lg/kqoxlxZc32eSFXX4wZtmb3+F/NWWth/uBVKt3PXP/nYT1
ssBFAyKlD/ftAsKRGtubz3J9xstFC4GveW9D6tCgT4Q4JAyhqDE0OBRBcPkwRk+khnChXYoAz2Z4
p9FLDIFtMJqJjRAdyGiy3eFoMDE+ESHmGsHdeVHXXPS/GPogY9HUnwshTAlwRC9FuzBXnu70Zdw0
WWXRdfJRVCRtLB9xff494w0VYrbjs29EkPcRs7GYI0Fe43nus63pgiddbu3EXWzt795a4WH4q3Aa
xyMYA6TnwPpTsJx0jv9F7vxWJW91m5vWBgOG7YC44ltgLzco70gq5NCWXC5JBFpVretEIhOvtUF0
eXF6BsBoLTmCk/CwZcgPYADEko7+dmhUGvnguOjXEBKyclWzp5ER3bUuWYNljYMVpRIexe6tR3mw
o/jafn8NUzwQWdDeVKcZb4HLA32iGxbgWIKhbhsfQicuc2SkIwy+tsrsZeW9XfkpdO/aZij/NLOa
0dV6pgiq8Lh5x/NB8extmP3DC/tYe+gmwdQ5+/SITXfKG1AdpnpCdX2WNaBA5hRm9Zv0/CkQ7xos
UBIUUg5AhCQF99QRG/j7yZx1CgB1maNBjTNRlOrTSHEXR53ePOxyHU71fE09FsIw95/i3exojyu7
8KgrTfZQZUdFrnuoZTvgNNA+LhM9IrryS7tlZZYRojV0vGbfwe7gmP9Lhz7r7G1G0TRLEj/PPylG
mkSD7QOZ6FJVo5PAZmeDw/PoE/WRq8FEHNBjAEmCmR7XIqF08WqihBXPart29//UmCLQFFhwimde
N1IS+ubafZbrMNTCqu2JjDHlvGZW+inrot821P9c4vLKoGFaveCVoK94tBiupkyxyHKNccq4GPqP
5buWEzUdxAcQbtr6Aw+NDx+g1yevLZNwQgSL0GvY1VXWgpmUUKTXEHgwtiTYQSRB5Yvi0gw75gYh
IcacDzILTr44i66LBrLOUvY642dklqED6xmJIk4jOfs0o6oo6bPKORzb1tn68SQ/RVq4WV3oI4Gg
5xaXPFYxG+TnEX07+ny6gs86qTqxErd0b+WElTQx+ImO1Zb6f/XDm4O1bbJGLfCkv9v/lh/iC8w5
NpjeJsqMOYFJ/gNWg5A3xFzBmgCZaZ+FTD5kJn8rwjmhFQhQjKhY8xNikCnWFd42mVMzxpL9c4jn
NV/6NHHhCOdhCh/xnOVJ92HxYkZdKw8LqjPEPURQ799PYjiKWLM9YdBKFIDxqp6GCeX0evFKQov7
4dvC/JMya8QYeN9VesdeS4zvDMEv8eISB1rvN5cGDWipBY00xtm1Z3Rom+rxOIEcVe/OUiUvLwca
A/xb6V68bshfALoMXq0nFnKEZPm1Wdc0hYdv8ktH17ayVSzxCzoAw9CqkmW1TyblDCLd+XQLWrVE
/XNL06FrU678JO6ASOtmfBd2MwfkZnzNwoZFYok4nigBZVzib4r87xB6WEM98BAhrPZtOYyFaAMT
+FTe6Zo0UtMoolVZ/B7XBLPRdkXKwW5akozOlPDusBA40j9xmL7PsgONnEnpNzfDr1I4LX5bGc+g
qNoj1APz2pm5tPP5msA3PMzZQcGAVkZ6/JMXVs93IB+57o3nFjps6Jed2xFc+0Qw6TLI45nKi5L0
N9k1Py6Vz+QFnE/X/JR2SPnyaT09ygTasVU5q0z9BVCvCsILfhtnCEHIqYvIplzBUK8K8Y9/Phm0
fixSNP44OOHdFUzeeX9lXlR4QooWE0ApcYhkYtBm+vh/2OygB8YkQpc2y3LQNcJig34JQRE3ro0l
Fazm9JmuNd0+rKF9UXyDwQAl+nTEHNBdV73oCCeiU+s6hRQIxftgKhNOuhW+sDLZjrW7bUgR5wJn
b5+J2LV+cJSfe+gLiakhY1SO5raAYNm01DW9FlB1KM88tBoBU3/mROhsBWS6OAP+qBp1eUDxECL6
DHQGmYbh5EO8EG1jtesMa0A8/F0UEnWr5QtRd8dKyT0Hmsbrjci1iYpAXOEi6cs3D8CFSyKk22Ny
irw7NvjVDYaUMIZkkTKvGl9uNxdpHRcuztRpkehsFoKzwAMSN5+tTPThGdgjPtRsgueHWmCjVrot
ORk=
`protect end_protected
