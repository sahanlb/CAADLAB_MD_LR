-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
LBaSXNhi7LVwbZmALI5Am3mZw1h4ykaPYyQq7AXsQFGgXVApQXxLV/FXISsWkk0c
a+Q8Z6vJSEWrOIt+wU5Xsbb7VuAFRglghAuHce3g3FP1e0bkELeWcQKt9+VfU2E4
nLJHb7lD0fjr+jJL3tadTBze82WUj+c4GbYzCldY7qLj6xTNaNpbaw==
--pragma protect end_key_block
--pragma protect digest_block
V6Gu+lU2b5xtotuV4Gz7C7zD56A=
--pragma protect end_digest_block
--pragma protect data_block
FPOSAEgVrgoMA/SQLK7+7osKX+ZB7uu21ZBs7C+B8Nv7hzq1tKSGp20WFD23KdoE
SGEX2O6zy2IdQwSW9uLZzTdAGQzKE7j1Nk1U2lMJeRChApsRplrvnMmyLKyb+dic
quHsUS2fUXhNn5/y+PZL2TmLgXquQ/ZqdQvP95UTSKvQqUDUu+KEBRiwEbmdjV1C
kvuR9Q16CLVmfYW+XPIeHM96eR7ijopwXv+X37xx61PF/f/IRKuFc62e7an1q78J
ODNJMOe3R7/g9C8otkCdTN6VqbGJKsvO+asgDvT+s/jv11GbXzEOg/AsbU5BEOYI
dcIFMgjBW1pPvvHPSO/ARQ/ONQLxSQh55Cd8tfciMNRAO0NF1TUjbGe44XLcYhQK
SdugGx+Rp74jjdTlbyVk5f3XYUXZQtujs0JUJ+1kOy6sa48JOuIkys/7JrPzRmdL
Pvx3nCdW5AaILXNoHX/+x+niOQf+5v11foIr+GFBYmCN0OBoDXQf9OpTabdR09Zn
ubnh3aF0K7eM512NT5kiKU8PAuSVCRyhDxlgoNnor6B1CCfLJJ43AeTEXymzpvi1
U0D8u515BhpHit63zfFR5AJgXt11FHtOj2bartFUc/pCXwX8ilC7fjRqvYKXaWCI
cdqjycLl23CCl5iipi8eb8DMFQgtddD+16bdCmxpYzjUzC/KrkUD0GmM2w+NKbfG
QnT7nW8ksciGYXV04bOERUZHkrcM56iNcL/0RgZWhxAV7GBKLGKUp0ddw10UOx9P
AzosG6JLYa0utyXy7bU3CEkfSvVo8TeKdqXhoRBNFEkSJyF7g3aNFnEojibq8/KU
9ZN05kUJCkI4UHI7OZab8UCW+hap58PQIZWfHkQr1KkN1KnnCK2FCn5ciD2+EPdC
Nw7vsh7DaWhZbv8q+xteL7GjkRyWzVZpUHKHi9ml+8a2be0CZZCeCNuALaakFwIk
wBkDAu3uS/StDVqzucgjrbL9nWx4kJ3DrpsGNd8k26c3e+m/0MoK1jq+M/PhZXZ5
Q4TF3pYhRk3c18u2I70FsDqB+5qkqgTfisH5VjoU7oZgr1gtWmj11JX4QGyYNSCX
HFC8CRomvvY4Oeqszw5OcEj6WDRmZ0NiaiMqJ/6Xsuyf3rCawJImfaZFbdABT+LC
fmDynRENc5DN1Ckk3eKjYnLeK10aC91BpouWE5SppjGJN2T6xPS7fqAl+1vqP3pP
IvVm9jDUhnZjmC3afygMgpgt6fbG6nce0ktaMluMm31xIkJ+itaI0bUm9h7IIbQb
aqaW0qufhOkl8GXsa78/UZTUS9svHQuLmorquxBszjTdhdZYz9BPrneasOlJ1Lnh
wAyMmFoXyF+N2PzZMPKKSECwLt7G/9AfxF3YKxnnL+DCYH+JFqLW4n3OF3L0IHDI
0mTJrVBj51jzO0ezfCjZ2yBkurq5R/eTPqgI8cy3XRacFVnEXvd9nuEohWKdsw6b
AyGz+moh8nhiqlZQGGgJ1zqE32GWLmU/mKet3QfhBOssc5IwPMyd4JfLqlcfrtqj
/WTuKuYF8XsqNyrIsK4qpLH2TVn5Fq+7sE5Et6Med1XKOF6+0wUFK0uCQR55iQ0J
4UBxeckoBW2o0xrhZPJ+luwdyjPdNiIJvUhdUbYhz942S6csZJcb9iaPBOOmT9ka
0x2RR81OmyMaQeFw9t2GYRQIoTcMu/J81db6a7qJLP9hPfcP7uS6ENJwLMT1TjNY
hU4bpyBhI8CmmJ5yNbeoN3ZUrCJTgwoabytXQLk2b4OwB8JvTOTDJfhwF1qOV2+S
LCA0Oib72OAFVU2MXwpCixqp5usvdsm7E84IZPZijvmOyRcpKMtv7M7dR4gr6pTA
aubYPYyER3AivDWFiqHLLtAjpB6zTxuzZdjMHryCeFDmOfLQrQtjX1JVjgJgw7QR
IZGY/dr6WmhmevVDmpqAOEB1IwUV5vMNMpKIiKxyt9yu+ZMLmemhZKzZdgwDpI81
fo896Qzidc3B+w3/FclEO//a5PvETS/0YO3SCyiWvM2KHxuNga6SfBrztxOMdIcN
zSlKzxdg4AqRkOH9gDymOnL9yFveRYJ95rdkFkw9Ref+Rbj6++tqn2xG7DfKBQSr
O6wHTXXYMF8rzA/jveWdQg4JDyReavErBA5OjHj8on405edg8j3yzsSgiflHpJd0
D5qVo8LhcU0GrvKIsT9e2eLv+swsD6R2oiI3aJ8tW/PW3txSfMovxoWckgCaNpOK
2oc8oThEhebUOhcf0G02KyMjYpoMw5mQOyYs3xG+NRqmAwMyw6bS8ZD24pclK332
M3jaK6NRIcbu92bXayarsRQFQZ85XT2XEgjAGfQrZwsO0GcDy3vOPMnh4PgX8NWL
3fbNjpHacKEz4h+W8fNJE1V8czeXM+RRfu9EdFeIIR6UPB8e6FkygGMQmO3DpIkH
4jII8EdYwV9tXg+r/pbE3KlUKCLD7HuoZJtNIgLhBmhrAy+ikMMOPpsRjefUXIRq
X2qkrOSek3EesAVI0CkO/MrFgmtOmGc1Wenl8fCCruOxR0tOETo/pK8A1rdygJO9
+tFRn0UluI+OdXqyMSUlZfbt+k34XJ1WQxtyAdJbVLGuZCPZ9HpqWj3IMICpHCfn
chCWmO9kqdBWSjPHdD4HpTaUYd/VujFNczsPvog778BFJaIRsufIndTKlzFFtem0
9QQn74SQRdpiZmQfcyDJzmu9mvqzN8BaYg8Bhglx5cVPvAQVy5NlBn73KWiLeiFC
j9R1rqwCrlFaYriWySu+5JIsvv2p1InSk95TbLAtEiR3p2CsFpJjC73oADptizrg
1QQeBERnQV5VFiOmKPcG/e2NAucUIlXIAfPtwMEkmfMZf0jIYxmDtB9dhphsaWVf
2rZghTOkd2TO5JLdCXjfpYAaA2b4ARdmmjrmjgRQSsEgvLPXo9RfBtJ3D4NX5FZA
tPeLpaCBrSJKEHoaEpqJdf2TrWqCCJkN/qpxoZ1egOIMxMNjCuFht5DHBuNWRLYA
phmsmdw6ajDRir/4VNPotsGtMoGncsQtLK9/8EOBBOMhnBAsByN49YvYlrMmjtoz
qkwOi1RytM73pG8UjaZ1o0st3rng40YsZNFgxQq3kIORXYavxtPvT65BMrEZ9ZoD
XcfKzDfA0e2hktRBu7nV1LEUrzEsSNSFFC9nV1oN3p6vgM8YUeszxVQO3s6POMwL
y2zhlufa/RrjnyA01kWbqeH5socpyL+/yyQgFHJCU8DOK56zjilTxbhySGdJDXZ/
+oqdEcNi26OKjG/Zal5g+gu09QszTzKVwW7r0sOUEzkUx6UzzPY3xym6WaPbl+zL
m0MX4TMLLeDPfC/jE8QqrHxPiN9cnirfvJePK0kipQCo+3S92k162/z521E85rKg
ZUtPC7c/yGHr+oF8+AmJUvefFY0feMcQpbGvZaTiuEngn0ukgXP9JESzoEXpKXx6
7dbKzZhUwal9U3l5IGUJ/UEEKYTkDN9SYLVkrZVEFAUhep2jZ5vDaLuk0NcaK2ht
pjOcr03385u4/SkEV/uYwmmx0PMkWpzcpU0LJWBoTE69A2JwSkNbmnVJ9qa7NAl3
rr+iTqOyUHgPQx6ITNLoPocD6+V5dr7dpBwMJFxSLDuo/U3DafiQHTU7zBkH3lOu
D7Idj+2I1Nps4BOFn4sgrgJmI6eWiRsxoGyuQ1pQ/1AXGGz0Iw/C4rLEniayotY4
nYv8oy4+fspZJTtoekJe9bdNuvWKBYwRUnnvEW2dCKcL/R+OHg0CCDtMyFZ3iLTx
nm2qIwfVNaUk4+SJ76WtKJafTUDT9OwI4+UThiPoDULurcP9S6MtvxmwSnr6A0qH
UON1Mvc/QU8K9QfNKiaXLaHTUrTgDkPXWg3FlGgoGlsWTvLxYcXfaErasb53v53I
hNsdzv7DeriKlIe1oXFIpvErhy23Cov488krCvVFQQSLPvSUFikusMDZGuxNBh8r
CMyXu96X751/qRr1a0jOOmHYfbGFukJZJ8kbCgtA0KSYZP9h0UFWiCA+ClrQrYnp
s2vwTJKdvBZtdy17N/jvcr8gMsX99dCHqpSwGRilEut/zDAXyuwVnX54Wzftck75
nmL0T0Otil5PIa/otgyuucggqI730RUmunNp4tdPlm00oNbEocG1HcX0h4885/ka
vLJB6AYDCOzwrZBYkH5n3hL3c79qfaRSRDgt4LTBlboQs19GnVkkFRckQb8SUmDc
D+ukIOa0gjbQgzZsdvUAnCy3dMaEfxLScq/JRDugC0ww9RLpA+2rIQEjw60a0MO0
CCRu/8xJcvZKg6UNZwjulEo8fPhEAWtwF5mFwmPTUgkMtd5wXf4OTgb7GTG0RMbJ
hC/KVe4jByPIJ10TOtZWzkXFWYnlZlTVTP1jUVH48EGcIBjoOdnUOxIVjhTvrS2Q
hqUJUymvQtAa41OVGTheykM9yUDbKlGYUAlkowVUaT3zzNhtyxxmHIuUNg10zH3t
mRd7eudbV/a7MSJ21tUUQqSeiRLJywmneFfoGe5ovbKSpBUiakJYy8qPrSkVH1vD
yeGiIY0koj00Xg59GZ9xrHle6kALL7LONqqzY1Qs4WyvnSjCEe8iTtQBUyHH1N47
iLAIYruAiNvRf+97dkrVszA4Yvr9sRXeFXkGMD7p9oNATEgTejyotS8ZNgvzDlD0
FELYio1fUt98QuEnJp48i07JNIZ6O6OIOM3qzVZSoNmoMurdkyohZgs1yyC1stkC
pDA++47M3sqp3xOQczwuKSCFsj9qc4Ob9nAvpMDSev1XTlh36/3XD1/3KikZj48Y
DGv9S9r2CR8V6uuQXrKmNn7AjJ+XV1GEH1JrWO2K0wrpkh2Ez/FEcC5dhyBYsgxW
DMQbwwzayQ1a79545lPNDRntFwMlRkwNcYcPsBF8aeMnTw8vf5tojsv3MXvUh6bz
p1Oqv1cKb+av/SIwXZR7vw+xbc3RMX36Mpl61uqaqAKXeAz5hG/B6fiz80VXP4n+
1COyGi+hPwyLPSKpxb0VZMK+sC7Qkx5UMqaM2vpO7RIQyYrMJKA0bZqfH+IBBo+P
6hlNQ+/lmU7siKM+ywhjxf/JEqD9T6nA3AWUr9V+F3TU5XGgSYpAXiNV1i5dAXUt
HhxZJToETQkU3krWKtJ8GZMrlKwcEBbFa9LbpXUlhQpAtc9cqaZESvfYX06PiK3U
1kA48PHuDW9aqnncH1iyRYl0hZD9k277S7yfPnc9z7h6qKVZuQ+stbRdoEGQm4Wq
LZRPKladYGCCod7G0G5XGHhGodgp2eaE5Z/UC0NNpyz7DUMwujnaPqAtJZAe+4Lr
KwFUqDkT2ChofZ3KxIX3WKSA/fbUQwzaUX46QUgsefxhE87p+B1Af4CyA9Pa44nO
RqbOsPqMm4xPrmPDdxP5lZundb9O9YKjGSao4akPfBuZg93QwVwdlavngzvRriEr
HR5EF+fU/G9AAkNi6H32vCqgPK2El5XD/H3BayDRUVw8kxHGsiMWIo182EcMkRBT
g98sp+L6psiSYTi1CG4N0AytU9h25x1vVNn/4fWt/bQXw7j45Jtx66M/cI/LaV+N
YAPRGHckKxmm6GWK/bBXl80ZjroM9nLdl6OtFfBKyIA5oo+q98tATaOFYYEGg6ks
/Pc+iZ96rzoLGJ1nJSIarXSWhUUayoH3dSL/OLsThe3DMgQCltCVxjlGH8y4z3xQ
K52FOqzMnYQaOPGbWGTqYsxsyn448hA4fhJ0hvKdHktcXtwMNgo5IyXkMhkCFT/6
//TPi29M0UK6t7q1lBoLzEZlLDYWbUZTu4rLRK6HfSQRs8jaV83GjDuO2d+Qa+tn
gLt3kjmdYUZlv/aqWo2ptV15AWVrWW+y2ipRD1s+pg6OJhcHkzb+FCu0hsxTVtVU
h1GrHxY51c97cEWGsv2H9hpXTPkiNb72D4Ii6e7hJwYm1p01cf0lATr+fOkkGLod
K25O6gjpA40mLBwPP3/ouA7C4o/VuHJsO3tcJMQ9kykFSbRJha29QPE2BWdGLojp
MrdT7dUj0SZhX4YQxHcmYH90XSTn3sZnadSygQfo8zAF6vdPHtCLEGK0JGdoIzCj
nDmHJ4p61kCQZXHXjbyr1N6BKaxygcuLBffkrm2XeT/i0haCnLJQW+Vm4VRPLil9
BQA58UJkn0eIf5H1FT6hPXR7ZM8mu3e5fGyUuuBS2KGPvG0lqkNSaE9AunSHOnYj
8SmqKg2B22lxH2z4WJ6Ug2Gef05NM5l/nbn3xGuxozCw9ZaU19FLkQc3CjbJnKO1
U0p+iwkDQkoECMSPX5jeh4BzCXy438Jxsor94ifLg6sMscn2Umq08tFXr1ZiqJqL
KI6zgVYMgwuIY8g+nmvepqbQIqkVqxWY0njTrsunI+iOoDKoIhVZH0qyj/48tkQW
CK7BEfiK7I81lP0yOxJHVLE+5ZFIMpTg+2MsVM0WcfSnA1gI10gk1fgz1GuGxKyf
bnfUVEDvgAMBhOY2I4nClW8kzmgd20ut9l7SlQ/KcNrALGlDdIz6GvphPeq26h8m
yNnKbsceAaTwbxeQZXgI1rBhYV47tcs9sWXioVL4HqkccS8aTONwUkA1basF3bdJ
WrWWhGFXAQFmf5cZwedNAPIP13DabDT8xK6mk/j1kjDL+DAsh1oM0dXqKleD0N/X
kop3a1f1wI3KR2Sacf/DdN9vM48hyuOn7TQm+/Ge3GZfpjQd+lPy3DeVecxaSrIG
jw0/JPpQIGMih+cY1xFAcPXLC8g9cEpHHiS+OXihSpnSpa/xftWPupc3X2afeEr2
me7vPJs9ryBXNuo7jfKAJJXgI9DcdwBwxTbIaXV7NeX4ouKK2KL1aBoHeKWhPx4G
sdcCkPn5p7ZvjJmMXCcq57y0uphGju+pHPSTpUAAZOtKgpMxAjsto9sOBeKxqTVZ
soOwsS6tdRZVfUfzA2Xws0Ix2VvxwONFZeQtjYA3g0C//77S5OZJEzFcvUiVe1tf
KjMyAP+63oCWSrGdCK2rr0cc2EMfYHA1tJNImfSi3MjaGr51t0bBY4JBrG2Zgvwr
lZ7ChRD6Owff5sL1Xue9REb6Hci2i9yVnvBEz/+Dw9BI9bSbMXz2FR29zB2E6DHL
1bZzzKtqcfl0UtAWSfcHlgFumhxpIpBntmi1kG3nl9NIRaBYpVjTaa+VfXtY97HY
n6Lxu4N/vWFDAPoH9lNLj0kjeL+x4Dgv2zl89vW0Njped9Y4Or1Es0cv4aq7uhHm
BGifZ2nqGitrDY7Ugx5fSBhrj1ReBVI1iFOMALqP4EKfBz/1vR3FmDClaAMHqUxg
NwKZv5ah4Wm/LxzYIMruEfjyJpx52qg2SbGRk6XSr+byRN5ym52g3FCSuqn4bcQ9
JEe/st2SAghiHc73LWnnoifiyNyIlESJztWYU3padVPNt+TcW6zS6G+oEXKaQpZN
0oagd4kYK/nEgAzUVkmIx3x8Fj7X7jGW6/j1O50nQ/1ckv8q78lefx3p6CnHJDZb
eQnVhK9L0C9iLdfxLUsLFvn0eRNG5WQHlIy1A/VX5Z699XYg/kuQtyKcVEQ9ZTdN
2ohiozxkn67chn7fDy05V/hFg8pdjJy1agp2sAo4y6ieMDrxnBKnMf5PsbRFXmY+
AaG534sEgk+pmkmX0m5VdMErIN5Zn28871zp+sdh4FbDzHGo5mYrUo5ish5EhxgY
03mAJc7vcdCZs6djixpgu0n4u8pKou+23eux/jEjKElJW5qgwva2Pvhg0JaXgBDN
uIN4xnuPD1/FZHMO5qpcVm2rV/OazfetYPQTzdFgndmDrH9XqmJgBfSxbK/cAL4F
xVSPRv+f0Qheb1ILNuDsV/LKRa4MVTHbfaDbBE2jaJvQW0OG2Skk4MfCt93tJbVw
38Ln82rGr4B1p6AaHl8nWOqL7AnBiBfF1hNH715imaHzw6OFq6ZJRKC5qjVCcmPW
2ZlvUHMKIt1sMZ/X9BpqzD6VtLty8ryzNPDoCm1rGF2TLkPBxet1UELfok5vjAi9
+GPSDGJ52l0uybl3/chKY0xP6sT0PeAkL5tFQss7G6mTJpEd5HpDg3aU6x3nXh+B
yGMv5OlTjzx8ivlI0PrV7bzbLBmrZmrFzAExaMlX1Ce1T5unzjzb+BdtRTamOtd8
SrxGtad775k8fRSb2fI2Z+avvMMF4dY6U68qooWV/CQds37HcauVVGDjofslRTzm
qJgVZF9yYJ1F9D1vBRMpzPDKEarLKBVVtk2I7GjB0GKMy4eTnwSFrisW+u6Vz7ad
jgwXvG1UeQfFSdYESEW2Mpdpw1EDhV97CR8xe9QP95yZy25gJdo5xXZHcim3UFDA
VEKh7E/DbLzue08HLQKs1wF20o25IrzbeAudSpikvhGyYe3Ma0pwKLRGyaGkLWQR
tAWVW9GytI5R9+sMDH1RAXp8Tn2JqMJDg9/GxlMS+XMzSISkSjUuVKndg0SNYXmm
9SS4KFAVuddGobGCOveFr9ySFFgbk9VLVEfILmIzQab4D/wkcyCemEDYymtFbzb1
FJbEQA+HMM4HHNMunh8MI23yHuqVNRpQEtpKorTQx9BqcPELxnsyN9i1j3nHQQyT
Y0GYciACmesAPcMxDSTCDXa7cBqTjPuXwafP+J59kZKWoFchK5DoKsRXA8tXKO0B
44FqbnP4Gk9qYZPXfMB4swePxolK0CHxKtNleqIN2yWHecDypjQVr2GPIXXRyp8w
61pNCBOcguF6BiPOprsYrZm2eVHslGOmP07joujpnwO0H1mIUEpmyWX+1sc6Zn1R
JlQKOM/czmSIPgKHuYZ324j0Fb7UK75JLq/rhYiDhG2H4twdX6Tyc30LILDLIiam
/t1JK/l30v22fNULPIXuTmGVtcmSEblEwBH2gFtk7/wDwTDfjmBw8sEK3KnbXI5u
jRzm/RimjcOd2dQUtEDIIKwJHzTYXMkHk3hG3piDpi+Ck5VZMTRgkN/PIgWoY/hm
r75j7059NHHMp/bYKXzK6GqiNrH+8J1bAhsARnYV3SnfoRaJYmGXNmiQK7kPzdb4
4Hgz8xHCF0VBbJXy+A2cYhP0AhqKO+miZ6zs30/ttNxXxqpj0D+J7WAMdJszTee9
zXBHcYuU+l9S9mZG9imEMVMnowOt1sO7yeHHNG+UsTvj9SRbrcOLUATtSt34gd6R
Wbn03/EmNJAQ3dqe+WS10h+ZVY1Z6bTM/8O4FTxmCcR9FLUxH4nX8WciHdt6Odw7
OEJxwp5+swS/xftM5innzUriP/KyprH9nizeim2I45XjOGhaSTojNpQQmXv+M7XV
oAeAukZySttbB22rIU+Nml51+ngkbAvtVPOYrtJuMmAkQKkD8vWPLMovUlHpYkYq
mms1FLdCNUJ4XDw7KUnzhJfmjlfXw4uY5tSl8fE2lynakL/5uGYYenFNg+z7xyDL
KVah5TrdkJ+Nongqt985VNiDekpF+qiXgLKF6jYTMIrWM+NNE6i8GRy/0/dgrke4
jXTFeK4vX/btLSQlAhREqnjo+xyfbB6E3XuxFXtB8wwG+g/KX3HsvsOuoevLdwV1
uJzZs3oj6Cl6GKjmvkENa0hZ0Kk3d6IEvrlB1wBesie5Y6T7DWkO26VEOJf9E2Y9
gVXxHvcUkwCWZGy9ItQz7iWa3nWeGPPLQHisWAgDOm/GObFacOc10g22TPKksBHY
T5TojCFtb/+yfD0oM8083XPK71U4YIJplu/oeQVkKUojEBon+wymu91Xr0Kc8U4L
x1hY2qaM+079C0rHH/ixLTRq31hIbswmfMk6y9DXVW6ZNCy+NyHqs1RbzUvs8sMp
BU1SkWAu1Z5vGMlBku27nbvt6YtlGSHwSeYAOxzQBp8EIbyw+6guaXoQTBdyaHpL
GR+UzQ/dkrw5K6IhyRd48E6L+wSoxcV28oeA5RJzLUa3HfvAEqswtx9/Fp7kyCJv
4XaxxocuKJdknYJJFWY3z2U5QagMN5ub691JAK+ANsI+5hm8v4kVo/EwKWme5VkJ
OFiq3sFSbS9ohJxkEr4yinuJWLXIiwMjG20rYywRnBiX66csVqr6MO0cnCHEwdH+
7OByPxR8bFMJqPTGKHipoNQhJCgpyRiZT8Ewm1rYK4HsSlJiTChZWQz7YAJhHLgE
PBG2heeaVwBlHcqLqRYkgygNBuKueAVRbu1WQNFU0MXp6/s6rVho0E/y03PCj99J
EVQ3jH+YFpK+tYkZC/ixm2ifBAf3Rykpc0nymJYfwvUV3sHoSMs9Wl5s3+Zb7UQI
eLm8SuU2Io5au/3Q5bCn8OpGKRguIQzeycccxAR6WPl33BUIVU2nHQ58EqYhq4ci
lno2MvYYA3rZQZQJ5c+9C9bPJ1naS4quBEaO3f5M2udt6leIwweatu6S5ACp+DNX
5Ej/DtfRWkdtW+HMkV3i3OHbrdgb8Opx4draCqk+wsuPHEbW94/8i94aZEUaCZB0
dtMIZKY4d9VWzQO39D2O8z8fv8NiMzQ2xaI6IdiXuub70vELOBAMHQqo6xNh/tU0
AiBsrVgP1VFZovrY8ibEW3LhVPrRtr8LpQZi6wvKJzRN9DU7DZcKt+iQnVz9HcZH
TYLf61aAsBmqiTOc48WJKIMLib7orkLYrCTFzIYjbZNrBH8FcLMdlnkvyLtUTPzS
MYL3IdUMUEWRydGUKRa7gJlyi5ALA/HvV/erZAJnUzIp+e0CKjoA4xFZdyloVL7O
2lIgt0kJ8vRdpp1Tv86tH4HMTLRPRqKZ1qNbm/ELVuwNPAimqHkd0+2CUgKRgs5H
LnQ7WghMDOd6tg92PCgyYpFwho2xca4+UKCSpJCNBaAPkcLoUVKlt91olIfx/dID
QKr+aMOPPWZPH5LomaO+ZWSL8VrYTcYtfJVQ3Y2omiVCcpJO5cR1NJJDlnLm1VeG
bmuFWNT65ehPS6P5z4NxLUYUgC4VmWqqIf0j5xSAy0TM7S6HzL8G9yLLBvf8uCUS
cnJGJmsXBw3A1co1ZsRb7n+ZS56rlfrVrthtKjWLprJ6970WQSYE9Mn1/2WVpvmz
ZMHhrcYV7wxDVrPejJtbhwybdYzDwRr8+h1na7r9IHcMj8mKdpzc5ssvqfyP+f1Y
5x0XwZNFYIwcaDuHZ3Fs8hGdhpmq/5haPSrohGIx+pXgNhfQgUoFRMzGMhQRDd2u
3fO8s8DuW++M6zkYZq9eF6RZE/IZCosbE+kG/y9JY7+5k3/ZP7euj37QXpsNLYb/
676TwDqg+p20GtHEzshw886BvTFNa8r027x3W5cEAPFtGN2vxRoLmEPlLHp8J6s0
9R+cy0/hpXGs5KCoxZ3qquCLzDyeQyu/62Rfkx1TJ38JE/TS1MnMmKcwDUA5WLSW
kySCG3Dlogw98Yjd1qqrkVDVAnQsRoXRo2fPB+vPOk0fD8biOutm8+ED569q7qxx
Y4EyDdACMtES5M1e2d1XFMypMEnP6x+sIrvQlhh4xKRc25dAmOxB55ynAVVr6Szi
Jjzcgan8zmZvbXXprYl/bPRDokDBkM9aXP0BIUt7tnr19GwzJsUs9NfZCPOa1uAU
p0EWYzNwOy/ztle3JIEos5enR8h2rIDx2oiJZkMAow60VvMfbt76RN+3rH40ToDE
YhRoDkfeBS1V6PO7u1WGTRRMSbkk0t7paELatby6B+INQKdfBWKb7xr3YKokqjZ7
l7BwVMIvKmbhECET90+zUCd+glYH2htLDyjIekTAXkKOue4rCnw9deAzatxozNoq
jxGWWMYTYSQEY0o6NpYKegZiMHb93ELxU6yKivWS+7UKY6q2fSKny/Eapj3h1Ph1
PSp6Z+VtKKWNNR3TeehgBgOPXb9vUr/WKePe/K4N2/FUy+dbd5+tdPjS32o56/pU
jMoZpslm2kFwdgUE8HVxw61chwTQVXyKkqroSONHrJyDeV2mllqKIW67whSb1D0t
MU4FvpyzTSD9FfyY4d3nZrWH0KsoLBquWhWhjNB1qGICbNsrjI8zN73q1IG21zKG
9GyNN6feXcyHrrCZ2eAGb9gFa7u6UgEs7rKlMQNo56R8kL2Y4nazBZmXV89YY7dc
h5BcFl7AF9ybOuy4qoCw4mcpOsVm4K2BPPpEYuhIJN8P5HD7NX+GEGeQkXJbvqw7
uotT1Sq3Qhr+7ZqPAf44A0ZxHw7q8S+eTkWvNXWThbW/bGZKFW8Lfi/KLfMaEqRl
ZaWrAj0hzqDvo/Vbky54dqKgWMefyZp+oDNmAlG+0/03fum1a/KiNSsVgyHUpyJp
TFk5OqwvJni1G3FkfdWQz80neZ4YjGFYeyNiCZahUG+khaQUSoDBsiVTsI8ONZwc
dRmj9+qT8qTl9DCObAajCJhLGvBBiY7nq/H1OdRJfpvXQ4H17nK5XSwgqxwmGQVP
R2SWqPZ86gsw9WdL+pW9dlheFZKhvKw+zijrl/ISmSaeZDyOnzPUaPeEOG83bPej
cLuQhG8yNgTLsvfIopI3cSZUKxtDf9ftOQt+IPntmrIRbolLFNiXpeG0eHXYWc/n
AD4pBv5+I98YFqajQ2NsuLU6voqZZdU/SWgssmUNWH+V9AqmNqJHFStIc3KMvr63
Vo1aZg8hOo4ggXUpkqMTmGutxJCzTu1vAJVg3GtpcPeTbXJZjpRJ8I6tbyDUf3M4
48SfZaPxTv5x+myX8Fm5Dj20fBa/dnIHzPqRnJsgikf2mfnC1vVAn1SIhP1jBGly
BPJ9peSgjzzHllc+LdrgmcnUqiwD31Nwyj/kU+GPD8XYBl1A96NvYcj2Ur440Syc
vjwP2Gi01vldAWjj6AHrlzD/HYBzOqfCYc55Zrv6AKSeOtOyo8mz3iXR78AyNLaG
M4pUnX1/s0a8LQM07SvrbAK8Not9d/Guw551zj2Rd2tpk9vUevj2WcHfoXkWGVWm
zjoRXtsBePcyHYeew8DH9LUJMedWKTgEa2Cz4Ki8+sk1j5d+cUybzKDo1g4lrrcZ
Q/Pyr/Ufm8phJfkzpn141H5//olxFTYC6IlpilqXl2g=
--pragma protect end_data_block
--pragma protect digest_block
2qzmwTCTfRUYh2FnUoLr9AoIym4=
--pragma protect end_digest_block
--pragma protect end_protected
