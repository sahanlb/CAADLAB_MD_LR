-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
daMm2Newz54pCdg738+FgQnHGixG17GUxPDlTnXNNcxFEIqnci+wQ/1h2AyHO2bJNcEwYyiqFHlz
7tC26SubrlhGCztAGlFttCzMEdlRKz2pF/WCXhLbqjZhKL6DIsbn5utLHmq6pSoapF6ZfagoVp7x
IsZFyraszKOzTK4eVq/RYDVgfK6wR2BEH8OskrtZHjyp0IClalRhAH3Ot91qgZX/Qh7j2upbZbrf
ut5PZSB7ookQKxIMWW48RL0hOxNJmdyScRpuCbbUf+sj1/n9RfHaWF332zSkfUV0I4lQrMlI8FSr
9HtFPVa3DR+6PyIKzWQX/nb6A2XeRddTxKFV5A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 41984)
`protect data_block
+orCzknJF0sjellq+DXCIbDn6gMKmLFZCxtNibsh3WsnETiUSR0x6kLtMp+YjpKUKrve81/uv1H8
8rwluPeCIEkge8ykgD7EI2/JoHjIecAxID1d9jXl1atl6wivmY6BHC7Qm2WLROnhKpnoYV3daC6F
6Rnf0o4ZMeoRVmGmtLfSznlT5X+0e/Wy1Pi1CUy9DuEet68N8PsxWMoKxocuGXKLKKDHnKVx4KA/
ZwUzmCd3GSKmKSPHrNYQ1soekfa4Bux2+BcUInbvGf4N1kO4nFxt3CYnGgAF3YSb2QKtcePuCZ+s
ED/iibVZyNRkhf6htwX76AVNin0LIQEtlXsZOcYr4hjAid+NaWejDibi6qYu7vOjlC96xujAdPq1
wzSXGEZyL7T64lVE1PwijSnHhYsbGWBbq21sYz74d8Z6leYZkFT1WewP0xleTKob+2eGWOv2AMQL
eOL4pDRqn2sqMMar0vyV4ZvoSqDG4MuO/iLjF7DajeBxNJOm+LIc6xGo4R3r3MJ0pkBe9FrIYdUp
ZNBNJBZ0RiQTOoiWdT2f6luouA2uZs72UQCKqS9uJcqNE0uHoUGDwvf5kzGDj/OfSm2mKXjKy98X
U+eTQXe7zOpdhUjMaU06yaYwzEBwZa2mP2wQDQDOtICx4d8wQtjGDd6KjJzL6mhDE5yqXizE+k6Z
WBZeFzjR0/YZ34XZH8RCA2KXzXgNhRnSKomgXJVsDowszChXnubpgZqqitP/yMQtXNknyWDlkv9F
g4p4P6TfY9nFizwmskPpm5qx8aWErVUoguQbIiaCjncPApTPt+mNwf9RLgBtntJKQV+2I/WCHqBm
2xf+v9T6gctfFvdRpogUULrujI/JxIhUhN6AL1jIXdEMkfDKro34cxikh4qobjnZWGPkzmRV51qd
5O9Q3mVfQ0zQ6p6iN4rVzA3AbESiYIitxecerR23D399ll2RXtLEYssWMX4LC45p4NQFTcY11DFs
+vnfhtDwJ9GaQf26rAeq4/j6a93T6vuczGmyQEZ9iBevJfRGeW5GhVa9c+KglHMtFgUIZrK5nMEx
ASaqY60RO0XmaZ7aThdIUI+ITmUMXwnBZXHd/DOWTqTQ/7qTH99NxK+Kc1I1v4WxJHvSQP8+Ccs/
fGiUd7feTev3F0PoyWKR3do5znlYztKfBPpQVdsZqs+nL2DTCtrN+jEHwV8Q3MXA4lzuBd/0fhdz
u4LiFPNKRcuG1J4JzMjNnGEaYshTT+LOpqsktv0di1O5fO2xs6cZs3xJvrVdxx080L8KtWPwV9sh
Al9WfdnWAc4NMHZ3FlX+5Mele9GP2u8ZDIT30jWlHVIm3X+LFxAj1JZudzODOqzQp8y7ZZCpMRzg
0pPoqGI9ZBOuNHqddsU4zl/IRqLzy6Glh03sIXPnn+045o9Op9m+XJknPn9KcH5dMuabLbLdWuXm
HEtBSko4P0inDqppCeTdv0ritLbNZz4o/4MpqjrJKncNF6eo7rqAqTVTbLFSwGPT8Jw4lonKoWsk
hoq4gx1k8+fnHR09iKxotaVfAxPX2ArqUWUv3pg6FngbGv3aumt9vInPVsM1XN4wpGW9q0h0Gh3z
z3ADr34oov2inHHRu5tsT18Aq+/PDX+LwTxNDbrh3vvwBHGwU+QjT5LHTPCmX6xNAAScK701/Uu8
+AZDekXUet1RO9zVUTNwuzWH7Xu9iTuClXM7y6gVP1/WRk9JumJ3N7EKNLjLZKr2w1AyRzR1HMEi
ckHv+8c5IK6PlHPXtfoioE3YxzQ/p4foaXZPhUu0XgVteGOuaqsIE2SQewbwJW/1cSfY7bgIaIeb
Jou9ObJ4dlZ6eahONGYbW3azzln05i0ABaZo2d6xNhrGWdVbyuFLlnNgc1q+/mbfa02p2mY6zlxQ
xIOZYKAXYNHy8tgma4P001KxqK0GRkyaTusOjfRvK0EE9nlE8WNZOVA3b6PE13lM5mhqRYnt+WY3
gPsV+6c2Pet2QAIZ/2ip4PD7ipSWr25VYd2vFWjlGmMWiOy6mkn9kDdTHoB9zszR9AWBZh2cGkIB
IhWVlb785S/b0WOWqaK/XUbtvebd4VIaLK8jpWB+b8qAYVQCuYJTxkSVHqXo8moTzl/vAVq1f9XX
FW9RXF8oU6AaPz6TolAd76RD2Wo6Vq1jYHIGg6pGCzUqVUgKg7Ze21REzHtqC8QbiTSw4QXjajsH
xX4Ort/1NmJ5DSvyvhZSYzCenHEMujW6Nz2i/1I6zQAB0gzDvqXjV8kVE4I/B4ZflldmUwUuEkEj
mk1epfZqFO1h3PVSleHkT+3t4/8PdOT2dsZU8Hx4ow08tCK/tV92iDyrHRN4iFZwfK/0MTzf1nkP
kC/lPEl3v9M4j2ex/JnRy+fCofg1RRW/soAUP5aizeYaXRVwFUfVvpHTq90MsMAiIRIp+oOLNJyK
uqubkipYUOTUc4+C+MJdyycvWzpmjqs5zCpvpSx3RT96+KrAe9PG73wNhJmULFD7DOqVvZHQKFEv
UZEaEAwe1Inzpe4bLlW/D1fbd3XFBW9FAEbpKWV+FjEQ7z8SbhpACbSsVtWGyClE5U4is4AcixTh
j2lpbSST0hNOKBpF91WpoCcuuHkxty1XakG+geG7Fr/Bucro9LemYh3breYbrPcbBzayzoCBgeKI
sJQZO16/3e4dwnQuLcLbdU1wp+TutEQjLFReFox3uAa+nADIQh3sgGZ10DZ+JwV25qo2BAQGss2o
MTOHZCXLVAMecivdEV3BMH+ye+6WOkwu94J2+9HW2Fkg8J3jkuGc1L/Gus06VaR7pjRqbVfMzmtp
OKIti1Fj0f95U/PEH0N8XHWtW9g3KxTeYytXo1E7uQOWWbro4IGhuGPQ7NpZbPueoy9jZym7pPHd
DFyoq8n639o5a9+MofOYKAGXGArh2DqaeotO3dZ4ppbZ/VY9G74l5HTvAeGfZMaUkmo6VPdVsmfX
HzNUMNxfnLtjm248WuOrbz8CCYrfs/98GFwDRJbvFhwFwv06xKdNtgE38kNNq1kyZUoSohXOrzz9
feodG0cyY/t5AwEYlzdMPTbt0sFCM0OJbqDeogwhFRWu0s1wN73s9o9pgKOU+0G105p4mO+au76V
lM6/x9PPG9VXKsqX9ek/Yy4F5PN/H4+SwuNn7Q5m+pEQkG8KGl7RZPFOfK+JO0Ks0+VbJBFry+s2
f9Uatzgs2rdEDEUeMC9yA7r9k8Kk0/OubPqk94kqxgCcbeHMvMu0YJA486uXctTJpP2WwQwODRAM
EA9yfqZYi14B1GZBzhlObqsndch2ZrD1TAN0B3JCR+29QUQeSaom/m0hOWDyc+WcrnHY6bWcbZcb
SB8X2yXY+gYrAIOo+I4/wDzC4YwRQnQqJS96SP2cvrJOObBoRwQIk1PTpzw4Au9YQmxpX6VRQ09c
A3B+TgRtMYq6o40ye0f5XiNTAYxz3g8lBX8KMYFiLgppQ8GKhIrT0udj5JsRGQU+UcM3KkJ8PtUM
Spe0ST1AwQZRx3rVHVuaPcJB35pfKH+FNwqhjEkCHuzoQ40knZfTq4iJW4XahfMH1U2FW/p8j0ZU
Z0HQBLEbqd4zqavnuHYpXcbidmu9oiCoZsd1EI+YTbN6HfF7JRTeBDiMOG9M91DHbpDgt419tCcu
tTWdrgQDE6szM5ClC268pCeyPyislorHEK6SVLPUi11WlqjKjhbTiDDnL8nOB2Gs7rW6DkDtydqz
TGt1dF4P1KrJxUQmre0jdGyuegFFLNV4odlRM2Tp8uYZYypjFDOzUfR1+UvzWdSLBY7SRNJSVUtK
Xx13NUS8SFYv4pzAQZ7Q3E8Rf7z8mciJUUN/20Nx1Xbmtt6bEYh52Yy/wCK41DhqrYtX/Ht3TY71
MA8hd5r295n3qHLfAJTRCe6btyU860BzI+J+pxssJ1msfIz9OMvL8TqwvN6jsiMdevnfTe6G/GRH
GrJXd6/7c+4G7U09+n/NyDF7qN3BKlbKNkgIhqsHZwvIeL7AFhP8QA8xjm8aWyF+7jUohBaJJsts
UZaNKBqBo4KPxoH0skgMh00FLDOxEBxxRE6hI5bXtN8G7oPWZ5B5yRS86eIsUc1bayy5GKQWVEa5
trM9GiQqr8UMeq4iwl3efhh7jNxNnuef0Imhy3rdQpbBhNWYEGNjd6LLu+rkk/mfT9XEJ5rx9xQi
BeYeTDXHotxQ0P6GBh9v3w7MM0x+L6W04WgCgoZIHs36E67wnFWm3WSqiXFj1iTytaf3dGR/eg0s
OAPxrmHjBo3Kj0OH76f8JjSHVVSjO7X3RZRYXXOJw/SX+dyHJZHr41K6Qn2iRL6CbmoMoupSMHjR
fqcl2XaOA4Q4b4sx9gv/eU355Ys3+LZu/htmHBpV77RhyHUDHZiM9nPnTbN7U1f5XXm1Sacy/sve
vUCUYaXryYHepHmBtsGQ1jbjr6LZP+HORNCodcOFnY/dbJKJXonHfNcnyn+LUk6tJb8M24ns4sQk
hUZSt1XMyn1C6Vqpb0as/XqVAqlGWWtdWiGhBAKQqRSYhUnBWHTnGLXiwcj5Vg3OglP0Yj0dhkXR
tjDDCy4TLOP2g3Y1DL6CPCuIYgfY8Uchj71DhOErxBQM6On/Stp06TYvxbw9xNhEgjAxzmTF70TL
KxIDP2XCmaPZ+0Qt0OCPJ/UKCg71NaO7tx/X1YymEhIsH1EsXD3sJoGaA2LfWreTAhWZ5CjyZMGK
T0xfNSaWrscQWv4cOBgWrXfCPCVmuZwub9YaQz+jE1koHlM8ihKVsU3XGql+4eom+n7YjdgWMiT3
v0BLi3k1x4g0GC5MhLqjdwmqUnq8NJ9X1M4Uwb++U8Pb8BGU6u71WGpS5gjyEbGP6wTCyhj5AEqm
ygaUArxIGhig39OuLA+wPKkajhRxyviUkqqzDBEi5z5qqpiwhHGpqyaf1N3svnGb6PN8Ksro81/6
oYel9YZjzLwi71E/5aZu2wTlbVehNE8HSh+wP3AWR8i0nwO6awkZutH5sO0tXC1MArK2btl7FH5/
Er6QuOxaPw385gcO9ToERRL12OijMkkJHVP4ZZP/p5QicQ4mlxItp1sVvKDRM4T+a+Wv8nOVJNID
a2001s1KS6fpULl4g/wN6FQGHRa1BNTVisNo4DgmiqtuTfJAFvCfP4GlaGTchlCixtNk/qsr7KCP
A6raFs0o3L1+HLLgmUu0epT691/+kbs4EHruKB49oKevTMUeo7ifsy8C/Ba2s0tmxiOX4LTpjxsm
ddTwMtqnhLS5ITbmxxRt6PJj8EYT+PBdzVao0F4ui7b07utE4yc1cFjBPYzx59jNAQDPnFp3RZ07
MDNkYDG6p82K8YBxRGCppmggdK2W7ZT0LOHGFuTyznXATyQ/6Gey5TaVS9d6JrvCfRkRPAudkZyu
XviCv1CG55h72CdUiPft4m5qaUQbvO6wUiAvrU7R8yO05/3isIMPl4svwQv24Jtc2oWR85/RXhwk
oYXCJLHkDE7D3NgARl07wl1VuUu+W95msHaDoYzaV/eIjc7GHs84KoULLFP1ltKFig4Y2W2QXLfM
XvAjDCdmiKzBzaP3mbPI3xo+FGPpGMr+xdp8MkkJ7V5sVwsLJxuUPEdQbEzHQ9zcaEvKfgNsLwMF
tcyASlFJCGOKZVIekykg+uy3LsUC0YoQE9OQrsw7Uk95CCMo1ashPIbpfWASSEHO1lP31qeCMSRn
2uB+BHRfcWBJNkNWjHDOFdNBBkooF1NQn05QyLKdOXLmYTRrk56o1eQaI993qTexNj9qWC7nQYGG
mlJk5jQxaqCisylBsXQFNJ+eHboeDYfm3pmo368JBNYO0Mtb5/5JFEdxcxSIItTZ3kSvda5IkE5p
IVgvQNZEq0G7fSOpsAcIYWBT4azXIbjyGeWeceVQCL45VqqE9PCLj8ilKwjTv/eF6S02X8QhchNr
77opaojJPxFUIetIfuP8ZhKAsg5Rh2AYkmH/qQ96WylxWfJK9iEWudwabMTeYgONN+uyiczwJw0U
iDmA/30PDZYfpclC49EMa8ECbZiMZonYD2oLL6piog2i1eC/OV8jLRDHQFjGmrWFi298auRfdLdn
q6q4lnd+GyWgdD08awbS/SJm0k/ZuTlD8fF6D8lXSqYsMZySf0KyizSn+8x5xHAM0bYo9dGQ5ER4
WL1DDreuLqaVVXRtry7OU4vlzcpGWVynruGxOTXSPhrKeJ+a9Rr0ifn/kjhc+tAMhfIHMb54voKl
OBu4xpXSEF5eON/CNfK4+1NLRlujPY7eKvU8plP+aR61i/UOgQxmlGAHBcn2oEhz/zDgJi22fxvM
r3KpcyMLU5caFkdfn9eoevGf5R3+JmbG/DsP1NbDHPIPPI2ntdW7ONeNOMLACyeRQfxWc3/xX/Ej
KYQUmlJXDckir9oqlWryOUW2IOR3Qe01zr7CYHoa3TSLF1451yDavPnou4phmaHhyZY/y1gJQP2n
Me2Kxnu0NNu85tfX4mvfLJM8tD96MnGSSEEOMOrrNAzzqhKqrQvIsCts1J7UL31of+/UqdLAfY4f
f5WUh6NZSfdhwEWQe0eEW9Ht1+sIPJsmghsDFUvHoeJJhZXSxCJA53OETnnqbvHJdWakm6nk0iLR
4+BT5/SeevRUBQ59+ZOoVwkHC9zHVJARLJTV+w3Vmoq11mx0yMyfIO4jQ3xfzX4I+TMivAZuhFTo
3vlPt9UUaHFezjhf2ZDfVrkQ/q9szrphRNDf2DdiCFPZfkley46J84GB0eGN2E9ItKczx+pzcCNZ
z9OkaZk5vsndkuQfF05ZzFP7I2b3nC3EFhzCjYZ13HxWzRU15sQq1fiIK0yeT/n1csLAdy+eLiag
KGAeJD4kcF8Ny+qC3dvSfRpSJG6OJ1cIh7l0xeDv+9dOVGemSNLwVsXkt46N8i5vCvHGI152VvHb
ughSfiB8Yk2IKjiwPU+Fwu+wF/Ey90nHJlCCHr+rmDS8oz2UGGtVeJ+pv4YWkoEh8JMjo1BKsSYx
mspxdnnEuGK6GLNSpq8KUD6bn+Bjv6DB7GCxGXfpUKxTePlw5MkVNP+z52b4JNAg/3eeT338cviN
/csS42iSnd+BTgRVqWSne6K+t1Bw+ttSpsztXt1qPo+D1+AVzKMuNpUWrsaxyQlbyGr8shJzMZsq
onPmCEc2zZMl1ZE/Xfju2fzcdEedjS7vQrO6Oc8AsudGRhHowpe+73wRijCYGTYS28IGx3id+Yjp
l5UnYDuwcfdt/5Yj4WpNFS5oI8wY3FkH1eXhSSpbm/FGSyizdJaMVhFpkAZlBPUyVO3iKXVo1UmS
mvt+dEbJvN3lMbvYGbiH8iiPWV+iJBUGNxv1Q/X+skEYBZKlDP2FhoOldYHfbwwSbD0Qa0S5cNgf
lYDqy+c8t2HyX13Yjp4urGenN0xoRb6YtVwF3KejXrPgDBlbcbNsX+IsQUw7bA/pcgVQTiCJxoW0
oxTXXtTfPnhiAeXcCoc353LkZ2JHP65KUWkLCcEI/tZZo/AQDidrxxbngu57zKMT2irXqhrwbgkz
Q2KWfOi7NuQwCQdfS6B8okJ/Z6FBMKPUyoEXZVSUEzrVfqY2PwDGC5PFK8ZmAbe9q+jh8lS2hWGZ
m16JZ7ImrN4gmv1GQESBriA6nV8+Rej6JyUT8MmIaB/hH/zDpPwHXxmukAzWiISQV3AailRDQHKp
j2flyiy6jM30kh26PIPxqOjAfYdYSJ+64n6SyFmLMYV2LThXJT1WdoQ+OFtjMkHV8NQuonNAeRA/
46yTDeT5K1g+SL0mVEHJWZKwTocAOmt9xAb5Uz2wdwPFAzkEunXtZ5HeOi2F1Crod8RSHk2n//WN
OW/bh/fuZEPhRVg/o0Ka13NOS3H1lnQAZfzrUjCfJHNKfyTqDdQJLKrSpc1MryfJmAHw1sCNWHOU
gxMLvhb2PlsC8qCuq873rSmRRSVvFo9z1emUjRtILX+jvInvzMQ5/fTp0JNPigRsQGfCA/tHibAs
fx0CeQFW0RrPzZBXejK4f3aHBWZfjCVd+6rM3rBx/8HUtfzD5gxwnmOIHARjlPaSBIUkVN+L1AU1
XXGsuaZRUlEvzl+Xjigsp4OBe+MSMGxXY80WDk1loJgmpHjWPz0Rusv43EVbBvfajOG37wO9w+f+
47LoYJSI7hxilx3hRL6qduWeeOiRZoWrmhRVUsbgSVqgkt8ygKzWvdNRKeAf1CoW6pZukhItJuZ2
4gVxu28EdMJ6eVJQ6x69K7LzG23uk8alQ29Be1LMXF+SIjDqVM73Qbt19yCxxCvOIgPleWYtgvIP
YHg8GTH3nefTBSkxz27OMLMMxyv3et/ySp4eEEHpRxMJJE8R3WWLgVcb8gS6eJfTz7lYMRKNtkNt
L10bqwLhYwv3tPTbC7z3I9JvUe1zMkR89gZj2SLfax8qR3AVEm6kC3kVtTRXHZAMFs+t2uf61uwk
PjLHMGPJzNDvpv5vkPsEeIFFA9m8Y1UPb8wga43FR6esoZ4/JZtbs5HiVKcde49CuIhUuNgNRW8i
lvorp78l/AR3UBZ0xJCzPQjdTAWQGak0tMIUZ6cRSM03MrR4IEYL229Rsb/2defTcttUAnFrWHu2
6tGwAmZj877ArmfvaixRslQwZkjE26iSELCfVOfAqR+nSzQNgvN6I3TQM/VcWjPlJGRnq1GsP/N7
mPoOuYYMbuwGNNF41vOlNMfeAo0DquxLJJy2r6KxfCqWDYaYfEiZbNZuH3eb5gVrHMVLBrrzV1To
Kwh7CsQ0U32FQhZgJFRevPVyO+Esyl5kMaN8MvpdTYlQaxgALXVOKr6VUZ+BEyXS4rlzgu6onlE4
ynL1RpI+qOZ0n3jzjeaebM/Pw1d6z2LgTO/i7J1YK4d3c1V4kz1W392TPOZyJ1KnpmHuHFo3U5mg
WGYS2JIhAhc7Ua283ioOyFnyExK3/OTPGB5YJnElis3W7SA0gdpeWYXJ9yh6ehTlU21A78VAcN5o
hsDxLM//jfth8T7OK7ndy7cGwyFg47onxdsfvPE0uf4NWObEjvo1Oj6GS1Z6nozKZDlXmg657Zl+
NWGYcerlvqwMVdcmqqCf7KE7EVEeu2VxzzRifmxPO7qeEAhpFr5YJW5nEHtpexFl3/7AAqA6flow
4Xk/mW2ifX9m4iDQtVh4cK/vcK336hsisiURlilxIvFWun7+/7eJJ/XTI0RRicdvMbQ2PbPXPOCW
cP311BvD00hGP0GsjlowmcDKpbgDadN3c04XV5ehQmLM+IBnNmY5UO3OST1OOfng42vXkO7CEqm0
cNVnqgK7Av6hrkND3sZp835q+5VXTU7qoxk/2fimk5yJ7+bhXTnCe/6FUeZZGjWHCNOCLMS2/Goh
Tl2ctlYfhxv5MalPIpL3Iw7cGR4sQrT/XEdK9Oi88t/cF/ugOlzOVT/cbWA/TGqpHmXs8GFHvA4U
giQZRBqfDn0ky24ZhbdHDEjRAUW228arkt+Q+7ivapO30q2+IsbwKM6b5SH6mtcTqbTuc/RsQ+kj
i1paVDQadrfnvihiapkFhr9W0CZDh+AC3EO7OZsSjhkWi3Az0K5l+Z9UG+EOUIw5ZZ1t8efCX48x
c7pF8+hLwBrUZldsmn+TN1i2w7FElgpQzdGnndlMIIQEwPZ080LKBu/vuyOpLEN42P/6u974Pw+R
H/1vX/5OYJu8Mbh6ZJRT8aVw16auuIrHy63WT2H3dee5V7nHvWpu97UEBjGYncKMyVAPz8XRYemr
CQSZaMyvO+u+49yACGw63cji61U4C5sJTOz1yazmB4wdnb6D6QA1q+l8gK8ULEX2wt9SHM7oBZDe
Uvin/mqlPZ8QvemBLUfn5pBKIOk1EfWOvo+eOUn6qL21i3f/QSOJKFWlGJDPnrpWIvp30CwTdXVa
CmFxG+IE2JdnnAMHeW7l4s7J0Z1kt04Y0Qn3I/r2ObNEkmno28bNQxToPvLKiE80bYOooMzrN38p
hxRGygRCVZF8z1sCJHRWlxgwlcP3BD6cwTeg2SB2keQK4OvxDyt/Flr5DqX1s56pvmfALLQ3dOgk
g0L1qnJ2z/gYhe4rRnjPnVh+dmBCcLuMtQJGqzGmZRawthKM7kANgN/wZeatJ8CvyNeMLkwnMj1t
tTiBcnyp+bmK/DURRvQmhvxAs56zFhyCcZLgSLuLMBiuH9aR7wAdst4eh+XNjQsWo7RoJRYdrpnt
yy/At+Xs92F/valEF9GCL3XFIdWbRn5fSNx7SPD8xk+6i1BSJazEZClNzEZEOtto0E5kSzLLhKBO
I2jAwhLvAN+uXctBP0nKxRI3n1tT2xmeW6uQ8SV4gNk40Cq17qc/tOmEEqsEDbMS4FDV3c3RkjqG
P5ShOlzTPfzKFalDKmbIrhkNBYqr3BkWY5HFaCcmSwQ7UatMkSn8WWvop2+cmUktSEOnqfjDgH9D
W/+i653k81Km4+06gP1F2u/MbCzp1X68zZIzvmq76NVMBY70umeUW4ONJ7Lv0UFGW8UK5hibL04/
Bug5wZY4Auo3ao6EI1CQJ06hQIxEv6L9OMbR0vCPotoM0a3p213kzP7YVOGjEM5d82uyrSXltaCo
Cembfou++xWalBS/790x17xAE0Ppvj6G4fNFQpQSyBmnCWcn7tvAfA9XZlhWI/Y0wa7y9tvyvh8B
5O+Cp63nUM45+AHOJtOQgTTyD2Wv+MzWzqiix5bfl4Su+3dRKsmIfcQO6vTrP0MqUaKZJy95VJew
Cn+WdZ5axuxNW2pXGHidwuoLC15pP/FkYsjA2sIGs9JCaRj2p4EBqIMDnjo9JTSgnmFr/Ne4jEv+
qCAkl9RbHjj+mJei9PjRJ532MxRNfwabLsJK6YJbVvh7h/86KtvaxKYlztaIU9HlvaIFzl+ZMhS6
/nTfEBD5EtvvUhyo+GA7r0Jxfj8syn/Gbw0zrvsUsE1OimULiKZedVLviAs9yemjcZbt9q9J0g/i
u7iCNMjCMTvGeIkAMan6W/1CNExsa7/xcpqlf7+kWQEju7rVhranRnnciyrSAmRS6QziyCt2aLYj
92sZSwbTM3CnOlFuGqoYKtkW+/11wF8PlRzKclKyWBT/maRNZ1lS7bdij6NxLL9B921pTjPVr0fr
jH4wuB+wFF1buW1bHgx4ZEA6NSWOd4F/W2zkUr/svo3s3er3Lj2aRt0cq6tBCdwl4V1oE8pNRTFZ
76q1X/zsbBwslj3/W2HfYtCTmenjI/q531r0wsZVnhiSfGFfYTyviz+vjzuyuIxJTiy1cAZxHfS7
BlQQ93q26Yb17kASk6cYIOD5zEV94Mbie8wzbJWxQDdExWR3Qbh9smocy1tCB1lKZ4enwttF8c0p
4jR+oam/Xr4knci1HHL10Zs2vcdohoqm+shisBVRSg3jzyUbB+U2ntEvhDSD258PVvW/75CUxaTk
i4wiIp6plTFSSekwo2dv3QTK765SXn7z8bahffqGPTG8FOvBYe7klmCldMOkkN4UVbCRAII1tYRW
9eq8UFkqGZfx1Xh3SQffAhpkm59FKSXATfjwgfaHo+rGewCi6Ucpz279slg6cyOyAPJp8qCxWJKk
5BWfMPcYfp1E6dnV2PePOqdn/mcqkxpqouKhDMbsSgXwSTHzhhb5qnIVENdd3fV4tR9MVRS7M2k9
FglfPKovrHTGo2vGikdypuXktbHK2S0gDxcn1B3aVXJ2pyRUIqUjnRgMAfZzj69BM6DNYl1n3oS0
oWYgxVo4z9Nvxy6Be1CDC9gmXvWgjuPMp1w3WKBCVsy9d96fMg/eHantTWm3UGu0Io+aAu/DgKh9
XQEMkEljw5biWhWWN4GZlUsqvvUwj3euBRCjmNzGeOFWkyyBOq+za3Huhx7aTlqbNfiaxm0dAo/t
4YnqZgQh7tbSQSxLoFmS0AU9lYDY8kkMleMPrujmQal2SKFLOtI3v9Wq/LRI/Lyafvomzz+fb88w
TYF+0wD6HdqBsUrNWXTNF2JlzD2KuV9lL/0HY+Bp60Xat7hDzgdNuP/epSujeiiVoERT1lrcvzZW
ehPYZsGRH/cbzH1BAq7CGuuiy+s07Zy+xcLm2X5IH9XppjE2DeQxEbKxAbrxfclcLoqfqonaHTYJ
/VVoZb1ai8krmNmyhMw6FvTpjaYUKdHTmkGpJemuJvX9QYJWkEDcGwb3M1W3Mb+hA7ddTaxJ57S7
qhGgqL9d8FZ603yjm/y16+zzHTUeDYsrkC60XDemrzlNqUwe3zWXJzxQPK9KRp4U7jQFVSNdg64D
/jPLazfpnSPRs4FXV4Kgrrq2u/nCvGauKSIfQUsTzOrrjpSNTQ63ZXJgpFoNTJd+PKENpKcbrWwT
87c6MB/p5fBPnx96mnfXbyPPFCex1DphztYDL3CAp/xxUqZ9XdeJLsFh9XRsG7KxK2pXQGwL0zi7
LgOQBeGCP5nwHm+FFUpuHX7JaAzWC4VabDcqcgU3DXJY/CqMCPnw1JoLwQLSWEOMmYt8p68gK5iC
XH30jBuRlhvep+RMmwiAgSPlypadfHuWDGcgm9dEr53UkV1Mpp7lQ2bdshPPBUkcZZseNo/4XP9d
8CWvsDDPeKU8eb7tziC1/w2ArpGq1l+/OueiS6DpErvJI1m/dOnAltaP6o0fM/xkee/q+ETIG67y
mjjnsGmSOqq/kFtH2dr7y+J0CfHj27/MvK2IPualZm2yXS40bqu+OqZMJaL7FcYvHnYXXT8EKb2h
yovaTS9blnaK/oh3Zpx+B2AbhsloRW79s/f/0ISkAMYjuYNAY7YiqtWZksRCAkxW3lb1fIHKb9t/
2R2ckpdVDOm/OiSJFbvQ+KMXJqywas/IzEpK2EbLP7B9IqjVweZBW9XAGZtRKCiZ7paUt2SNSe9n
lHMUul3qamc7QobyCAS7ehaP/0hlUdAzf/uldMwaj9IyHxyXT5jD536mg9+ztcAcyHR8oChy2mlq
kzmK0j/6s5LJiC5msx6IP7i/P4YhKu9piz2q8pAB4XO4/gH66pFIckHzKvVbuVIi9zch8qeVh+QL
b5xd/hOEdpItjoSCzIwzkOSRjFFdVGIBL1noskzIEcznMRoNt9XHM7VsdsIQ5BW0I1D2nTHrQnVJ
5pXYtx/5zJp/bS98PvFAOtzJmSgRJXjLY3/UppfNEnZ2bLuArMamvVpVAt2j0UY3NLWZvmtnoCsg
OInF6g7vi5i9a3iQmKI8GdkIAujwQWIVMfckoRzY0GkAfE4ElSYM7qnU0IWNdcfU16m+mqCst9T/
SVDqr4htLenaf2uBlSPawT/SczAY9UqIEGrKoWyR7V6besz/+zFvvk7Fqp4TGqnGNaQJ3zVA6Kz/
htSLtTCDoFKJ6ToT8rACtJI4HWBxx44wN4aDi3MJ6zYFwt0aZyRnDsOtKEO9i0IuaB6pSDCvLXgM
fAgL5dwUsv/2YHPjIt3X21PGY7Z/f3Av3KmbEReIGcrgraem+kLqyAh5SJZ8rhxfj5J2zdZXC7y1
L2W/+QQLc7EYNjClGFnE4cQON+qhGAuwXbeJypss69Gdgpqn6IqzGib5ShyIlst06k+UnihvJEgi
Oasgfv3OtIxGaPIZTsNhqF4p/uFqOpa8rdTXC2RjPSlxu5PS+6txlhfQsXpHd8E4qCIP1soorbFt
uNzCIJ7ssrKrRjEXe33iqb5s2k4AkcDzkorGcXqEdjat/lmcU8qvR6nyUMDDSKn05v5B36ieXh8U
7yntT5Nd4LDsbjMtpGTZu9liXWXMNI3iEC1bCyL2Okt7I4tmpow24Y7TSfjReSef1YJXkoOicThz
XsLfTyBLEzUtQWtYWYbuohKGOX2JxdofWf8/6O3CGiOnI8pXs/j2NrRM0Ih4WtUYz/NEEMxyObph
n+HS01a82iyxiTRVbu+8cq5h+6XSkIzzW9vSejspu0rU0n0hEeTdo3htdWZzYtw3HwfwP+Dkb6yh
QxGGAQuMk+ByRjR7dvJ6ZUJ7gYQgVuPYZocWvXy13S8VZr2yr3Hg8ID+m9VWhPqhlYsReAEOsv0A
UPInSG8+1JfgGTxHOTro+9g8QIIffIBJW9dx9Q86L3jL5wDSrFM3yNaJdnFnXw8Cu8EmBeYu/1U9
Rllwqh7icz+gHpxYVp+lDEKO8UHpN7Qz3glrou795+9aWG8CjICK7cPTPk6TB0W9QfLDlgP9puuN
hgnXdZwU15SCpXvlmO85xTEEyVp0Ey+3LbM62djccFaJJFCseEDoC3zKA4pUd8tiaZxhADBM3G6o
Tn0VmwvCplSkJWJblHJGdzu01eVYQF+ln7JRelt2kvVBk3urPUk0JJ7gLFkuT3p7c7cDXcsrz581
D9xwL2RkEhS9AvvQxumLYcnTxzO/MPaV+Zg4FmmuS05YOl0BgM+1muohuDvN4cXYBKye32WSf4ct
atTpap9FDIja/rlLYM1J+yZX3RQS4VbImj9P351+TT4+iYVcie6F8K/K4MwT4C6JJkakjF7nDIRN
TAZQZNYd55Vu9XJAQrmjgYLP4HSp4pD2wveaG4/Tm8K7ZZtYSK2JiuKxwrR381SrpK1g32Brrl25
T+aroM/l6N2e280LKyupK2LFBTBCACRQDyNjAdsZK1Lh+tpSdWnfTLHewGek6gOOyi/yPnIiUZHj
JbHzdXOvWRZw+a7kg+QRwJZUUOOPPE6fKTQJOoFysLjQ+LSfXMFur5FQoupeBLQTvhvjQe0YCtGO
L5oaOeXPIOATblIwK52qeHBDVcfP42h9+HL44AqBlPM2NdiclzTdbdivQA5UnmDh7d3PkpQHZYDd
pQj05IZMPPMWElANPVCMhdwIKu7vmu3SYwyBdCG+f5p3b8h5k5atG35XjCGcq+KrkN6F03j+NOGM
maPPaQPe9Pe/zQnJ5fErBmAVB5MfbRj9krgqAW4pQthfMOHIle67fOx8Np7vyV8TCQkq1rsXewUz
GQSCpDVpfTTP7TtPxKy63LmWvkY/x7HKbtS9lB3ZcK/z6IYMhVIq/g2Tk6MWM+NkZnBKNa5PsX4P
2AfuLBhcbbQ89oXdkZm09U0MgmzyidUnq1fwZR5xcevBa+v0EAcQZcf5FdKsrtaGNyYIPyn7CKoQ
DEW3nWUQiFFQ/DlJ4WosY7ZTl/2SM5MiGqg+6mIfC5cicv5HYi4tlBILA94Xvlx20uIm8P1Kf3fA
sB9GsrsYazwQiSWJpeMV4rNssZOpXxqgTxUg0RaUs+1zm2UGYIjRy9qPeJlwd47Y4cnG9XRv03Ky
t4Qt9ep/klK6YCw0IcxsUQ+oklxwFiQ+Jh5P+Cy3c7yJSZq0lu8eluUo4osDPtK5IBTCSV7ss1Ts
rKEtOC7uPIuBAnM2XHrbzP7xVsS13EZLn6R2fIk/Wr0BsJnv5lVn1is5H9eML/cRt+nF8p5VzW64
OMAgsspI4WniZPbvc3Q5lTSBXE21jaRz6cAfr3L0cMl73qiIHO8Dn8IomJlrBSBmqNoT6UOa/WVK
eblqDOgdl6fZmJS3OwF6Vdp3yV7a0SjyeGcP6oYFj1gJ3nlcDn7k8wrm5pEPOr0/TIs9tOyUfAO9
2DFbc8viy8pwmRO4WZVhO0bJLlNWYO+57bI4DmOwziYU6CNequOPpYsXg6udFXrDBKlavRiMU9jV
oZI7Y35e1HArAClYnzTGlpe1N1PREe18BeZ9VgeQP6qq4Ts5PS/J4V3oG6c3CRd84qQmiRHSynVu
A3uGOZJhiQU7ZMXC+g/G8/GqmV7oLIV09FTvAddnz72T9welUTPjcNzc+Q+eaHeEZj4Zslj0otL1
L8tXz3yvWE1ZGegZtmyWogjZ/RVMg0Tsys4u2ToIreyMFEhFP+NptMddJUXTq3qJSuKN6/YIFFq0
Hn1doypPo0mdCxy5RetHNiBWEZ0N2mGuE1g5GbY8YWEcBlqd6UEr9Oo6eHeJifIddm1VOwPz1Qcw
VtUN7TVjL9ZOAnVEd25Zvrwck1hApX8ZQxUzSvPJM8C09NPQsj0K33Dx/nSULKI4mbtKOMoeN9b5
7amN2UDtqLyeOysED+rLSrnRDC4uY8fwmzdEKse/HtX+SjyU9i4Xq7xFVUzVydfZa7jV7HV5dokQ
o9mRTLEtxiE237zUHM87ZuupETH2FGJZmMhJ4VA6XJW09BtowT9D7zwK78n45au7LRNyh8HgFa/I
Xfu2w2pn72AWO3mqqnnaLcvSAsmQcuET8gYdZiHcCiPAkuZmOIZsIROuCllRXjB2flavEH4d5kHd
h8igDVvpghCW1nR/n9qgBBz1GjV+bMaGdKVMvHCpRVXRX+HckAkfy76T/ZyNAy82oOSMYwFDflBk
o5ftcEO2njNV+tswIuTpnnJBvhf4XQg2X6bMbyWl91O5GUsyP1B35xxChiA3sGJwYH0fdmGfF8hF
39QKwjD78RjjhmRubslO/8tElcfXrwV8KtLxYASHVBS4AkuJuB/z9xZwKmh9RIWJldmMurFPgbuH
H6EjB0hu/ORvSZU1PGgFg0kAR8h54LL05kjdonYfp+IT7Zc6Db8cvkbsI17Hc84hNddRDfnCvf9V
i0D6cQWYNG91+VnjFwQBKjk/8YfHK/H7fHKYpVQJh28KyYC97QkQbefW3NvCPXzbVOqXf2hhboK/
3nEnzbK6b7A6Xixi0dHoz0pvY7DS7dBJPY9PO7obYLziqOXC4EUKoPzseitbSSdv/4RscMHqlyo1
ImBb2uZPDAVbESYS1ytmbyuEP0NcF8PbX3NtrvPg0K+4KYKDGOByZYunhY0gRe2qmrbLkax6AFfz
M5/j76lJxwcDQCbgwlX+9ljf0dOYRDRVKcKkCAMPOC2cx4meW/xwYGjX2ptmS7tC960V/j92IPyg
Pcq+MlZoVBBDjFV87iX7JcJC3nJdhsppJffpo/3FupKE3gaDMTMp+ni2+aPBwMatty5NiPPTFtG8
Z54jepsekVAHW7i+NxR2npDlQo75+dBKX2dLxCDoTTP4PvbUBYiugOU1mtccHAt/MZjbtIN9qVFg
O05cCIy5ndonJFRVZpgIr46a4iZfMO3JZr8Um9kWy/O8NBxszJon+QaIBQv4xabK0eASNuE2+wVx
BoYbeyCDyRCgYtMxZhouc11OmmIqdsMGrQUc5yINpEcAfUd1qVy/9SRMbmjqO9WLVtaxwpA8HMn0
eZLFl72x5ydAJTG286qWSYLertVkWrPb1UFJWXe4PgjEF0D3SMvfcmHIf3sWgVJ4WXgVvsf8lvpY
CosteeuD13CUpGEAyLVMv7eOwOzmeGrKIkgtwwfAD79q5WRRgp2eSQELY90FD6+FIOhAwbwrh7LD
N5RBa1TDRTYMhzuLXFgeQH6LgEtgdUsYtBCR0UzcToP9OlIU8J9/gt6t2ysxRyF9nP8jVJgcctpJ
51YOJRS9hDkACXOZawUsciIxKxjKElalVU7gB9n/RxnnbTGQV50UZ4n5l5tP7AFUllrH5E7BGcqm
O78z9euVdRF6zoN2TnI+BADqtU+WEm+NpyrGMrMbZc7U097i3FyPKxV2UZd+j5O0Ev6i5GtWK/sQ
IZ2KOdE8rjQPtKAoOLz+VonfGaYZjWzNgmet3KHDIdguwLBD4jl5PbIupvWkxLO1B913LaP3IPWW
rpSe61FCA8pXwZNaRlG+dYbzAka62d3gihyuWn/kVDgVN0zTwbK82r3o2t9JjxrRxmY7oiqgeGv1
WmElcppbYsfPPbopbdbi7yJceGEQ2F3/aCJpSz3vaU4achovt6UMdpkd0QaMQ0YedVQI78hQEq/z
0ePE7dVbbAspDrDRGsClEewuUt50f2HcrQeU1Bv27Jvof/iZJLms+npZ6d4Il7Vx3GcagnBMgpoO
nyOtpTpD4ZGvxL+omUdVoYd5DAdWOuVd9VIPv6tOWN08a+56URxof6G7pUbW/uPnV1pYs5dV5W7N
sASecN8ZNylThKeBXef65FOm0q4jbscchVIYyte4L9hgutNRtOTguWw7xX4ufKXI3LnbYq/So5hj
RzAheRFvRjRlmT1Rck5/9mZ2vr5ceEwurKOKE7bjOw+1sTmWeEj0W8saq3m7Too4X/v49wImDbCU
gCBUuVxQfuzdh19r3RBEDRzeL8qw6uifoTcX37zLWQIM/HHj8QF4utQbD//eVTn9s2w9BCbfDpTw
JLu8+obKuiGXhRGBv1/GfkqzM7S88muGYg5dmrzIxfL7kRqfFZ23Prdobduesr7XaNxg3rLkEIA2
KotGoM//w+PtPkyzNt7naPfMrXP+Mxp425qW5Lno5yWHhCYRPQgBV+88kJnLk+W52bB8GLTsBRSn
wSdfCpkKoRhPC0ZbimFM/815beH4XWT00XM5YVC9cyz2KseTD/akjvqqJ2cKiJbl7cImRtcOWshY
JYeoMlo9DatWzITXPvI9b90xjFp+kEYwbVKLSjnsvBJyopeHei/o0xBc/RPBuxzV+fEvMRZJcVEU
f09nf3kTzMe+YX4rz5G248JcLZOHQEFMdfbrc5bSgbHeXWAAJZWWY6MJjppUYTWZxAQML0AyAQ1h
WY2MJQwsGganOZMBGl8dQgYMXQ8zmxnkeKm0x+uZHTJy/1K3MZfDMOpdOFKPCuAAT4ZWkSueXgA6
PC+93yNHWyub0KfG/fwjxcXPtK9DuZP1Fx83tHlH9CBIZj5S9IqhUcb2AZ/+5cW81bwj1wTR4ruM
IVYhdsAG/QWuYUw9utsIJpHwgRKM7ybpARHx8RRjgPdNrLKqMoYh2HXvOyHuVL0Bum2fmKMG28dL
EkPuvKgSJxfjmOo6CLyPblbLi08enZ9CIJoD9Ihle9EJq/AH7gvNxkBajHtBFMOpeYuc5TAXHfhz
zwq6OCl6PjpRjl0ViTHEivCwI/NA5i3+85jC502y0xbwB9k0AzPWVSx6ezyeyvy+5mAvImJB+l/G
cJ3UzBjLtRY1hMNAKe0KF7tE+ZH1g/Q4QwNDaTTvhzxzVrLDaWdaoTsgrctgtZvPSB0rtrSv+lRb
X9IyMdRVKQsmgRJz9KE8s02drPJNlryHAOP6t8FHE2Be2p9Vp7hX0lUxP5dSz0MHttioiW84SC4U
K9InqW1Bbt2XAzMSLZCEOX1vHkQSmTyQKUePwdgmMXOeI6wZwJlSUmv9G3Sx6VWsOusrBel3Yl8R
0E+YBaJVNgl74p+PKeoWHcnuiHacX1wIkHzK9Wdrx4TXcrdrfjGQnWhVd0rCR/iKONyEyw5PUrGY
KRpv8I0SXE3ky5a0PernXswtDPii0wYHzOuZsmzCa4lrDua4SP1S/bwAKnqzEMYODjlEFzSQYbNQ
W35OIm6P7FH49ukDQwlqGheeLGdbNzHulUTiTfFx8ozahq1zBFHqJ4ErSrV9ahMVlnzdn/4pOXiV
DbpKDocvmVQk4O6Wr+CfcrmOQ6Kxn1C5bgGTQ4Ul7+TUD/A+zQb42Q02EfNlPGoGUJlxwXXBjqmV
ybU7Kv+HZgV0smFJBTJELsP7cCZMR+M802TGdbn8LUXw8mHA2mvS6UIj12YSHzEx9atKUCsWnUJ9
vWS4lr5540n/j6qkleoTD8QcGi51TJFs21UHbn1IHk/e6YjeFtAdi2nvaOjQKWRkEzleX3rLyRRC
bomR8S/xamen3mzFfXjHC9qefsBNiBfYSrv+sFiGSXJ1UI+ryWAIJYMXWshtYW4Y/dmX+mVnlMtI
pvhGe3t7OcCyOzZ8pYqkZxj9yQyjU58+20AC/Od40HQhCQ9aYyzDekuuBbcssUDk0bTxA4W37hNq
A/OF5fw0sXpZDVh4StP+052M9wx6jdaR2uHo3k4AjfjVB3aNu1RojLEovEjUovj+aB61bKYG69lN
ZEPG3W1LCFgqZPtYCbD1m+kNiMV25tXuftiJf3/+MplUpO942lbCcfMhs1IGBq7Kp/VrmHqy6qYt
pC7+qnZfCYYtHACpRy4Awx24n35VMdDaobucI9rlt7nHj936zOwiskP3ojv9u8jaexWuWD1KkgmZ
BbjIQtVEEyPzHZppTlYD98wF+s88Q6a/XHo3YZ7iKQx5ESSvfFzbo8ZsX2rNDl6g0UPbA4gu+/Lk
5okyofQPw2nO7aAm45lywXjsaLHaeaeMTGESPfozMgvTLX3IAGdtf5GqYbHBuGdKNTBIg5xPXgti
qWNPWJF4bnOt0G56ehQkmSeCW7vFqrR0Vsfnhwcifm+pBrlnNPvPUVHOVAlnUAeEvmetYM6rJkBY
vgvPEsat6NCDovinb2mifvHzCQKnmy24dN9PYlVIIXZDC3foqm7vXt0WmQlQMoTmpKahGAWboQ+1
sV63wTj1fE96B3q202/ItgtT4cGjw6H49VIECMDLZANe4BTV9ifSkoZSjymwAijjCH9WU+ZxNagO
1qQy16M2/cMznQ9xi84GDc9suZUW1NmEDuo/SdXMLjAcZ0Pwh3xBI00PuppXjQRDndpIj1qxCy/s
h5oHqsoWFJL3Jw0PUbANUH2Z/LAtVT4Cu9n4STU7UO/iqH/05fjhPp2HuhGLHzABvygLawCJhq5D
rzN6p8paE4uG6ZJC1HV+auLpY27F1AaklFksEtYXbNS6qatdPC63infz06fXxkErdUaV8/f2j754
8mnrRI+mVVupltBTZ/g5YHCvrRrikLQlDqJJ3GEWdR60STNVkvgx/LqchmUGyDb32MKySFneYqw8
BPX5nsjaWCv3DE354cdGpxObtbsYY9adCoipix3m4OCBYULQ01zQv2xatfs7sVh68Sv6CqzoDS5u
yj7KnS3q17P9Cerbd4iR4CqpR1TL7FhYb09LpI3ThT0tBq6DhkXXyku3c9sYNScNDGYoIAgqQJ12
KFXh4VjUmMCNVd8s8uWww/E0X7OMJivuwpyeLgNfq7d8ndQP/JBortztHAyZNJyXrGRr2XgJ2G5/
UdHep4LJEfbA4NZxE2hWD4sWRmo4jh+gHYZe2EZUFqmFvrzt/H4HjBJGK32FnUnOWU3KyVoP2iBm
wviyEATdEUsoJ1H7zmci/YT6dTiqDzBsSmgo2ulVLE1HWbhAve/JFAWLaYHwGewiREI9czuTW9LZ
ByLghzI2/FE97f/Hz1HeIAND2cFIXbprVZKSmb1Cv0pYxaoa2D6gYwLlTjt+pcrRwmnnJ+YGrqeg
mzs8wm00zn8HPzc7C1SOgj4eBcTBZCOFa21/2YGbugQnd6H2fGWTbbZBlTk51OK0HyeS7di/Yhn6
x2ZrQjmLxwnTlzCy6rDJC06PJ73GjHpe3f2lWKD/nA05yF5PmbuzydU5q2CeNVaYpXOYMPd4/UeP
/859FOfYMa+LkKUeLX94yNdzirbuUqd/WbfbeHFO8UBM3TMureH8tpfQw+RnroVq4ONFUrN/qudk
YcJ5uvk4kC1/J/DN9B2S2D//t4DXA4RLZ40AKBuUB5i/70GC0zIKGLh1TZlOszs/tcrac+zQ7WO6
P3t8Tw9wBIfyEvFHEro3y48tqpy9fe1Nx8XAETbXWgu6u5LlwsZCPy/RMYtlzHX0RukPMF2Fz3tz
xAh+jY6g+QFDycsPefUdsPFCpj3asjc30yPbY2MY4ncZkgFSqxLUHw9IuqeaWo8EsVLVx6cJaiKV
idr9ZlV9Tfg+TJ8YUtOQEPvQ7nLtythpZInCQrbxCB04Q2TKdkLPA8/FZr7J3EmIyel3gC5QavQY
ExKyO0RsTFA/b2r2dTE1K8nbpJV5AGWvwhPk/Ob8Kr8SfNMD+QxBVih0Ea0lMZhEt7N4ky3pbZzd
X0B17dMu5Td8bnTdRuMw+iD77VEaPhnIAHP0Tz0+FVfz56enbC7rTQqGty23bGWrQ7ttuxLwHsOi
e/ixB7ca6oWKGUDB8vHA+Sh2n+9AbPUgaOyXruKPKa57/1R4RV+xPxC8H6XtZO5PyCe1SdzUFB2c
EmYYUOdjcRzVD3ZsW2fNDBKV5pbv5J9CrBOvyPRb6SDe3mseoKaOseDSOpZXGKRuuDYmMelCwxUt
ZyZqXnCVbZNS395QJoXgqi0QbMoRdv45b6pGVBvchXO+6httZXr9nrgV0aiDtL6aIaW5abn24sWf
N2on55HQgyKETPwL0I2IugssbTxv9YFD2tUH6sw92QervZl5gOHjgabO7Z5B2aMQ5PTMH5dYTdvM
gKTjFrhLbX5jgyHuogdXHgAGvCqZjsiuhPnpv3JmcenHYYznYFRZebxsgQB3UgYdV9X5cjmcHWFW
BnTT+6FksvMda5TjVD9m5vn2auV0i/1fAi6vDe4pStSPowxBwydmsk3e27nwG/gAf+s1Z6jZpItK
z7LrEuWmlZuRh6vEPxcFyubEh0zx+FYspiZ8QaUAGI3JLErQWFb0ubbcgaSsEAkazsYDQtY3Lftp
NximftTCUnBX2HF6PM0hrRpmGe6c2FeXetvz1wowG7FjwWfM2RlTxVRio5vRHRvccpMosyQW9DmY
/VnN8elOI5WiDXp39ETSxd5+ujy7kh1Fc2fhTdTSOw5kZG7sYGUVU+ZT/BobdQMSJvOKlDzo5Xc7
nOpaNNI9l+ubK+Z8xVkRxZ/fHXmIGjoK4ZNmMFsOiqiK4+B0yEOnQUFUMkJlg3RdenkHc9kxMOoK
pOo/gMcs+VCGTKOVZD+t4HQe1myOhi5juD4j55sFmlltXHsE7BGHNtDqXk3F8cuWa3qU0VRGf7MM
dNpkj86Vb5r++ZB0POAi7I53ECF3MMfY+KPL/++EhEmrmx2ZmtMr77sxyCvoKAyNTaHJWXtJ6tmC
F/eBHA7XRbSLqpVZaiRkx1S20btBBIBoFI1VgL/2C+iKRlFVQudxF90nlUlXLVtGWagYy6f6zji5
Pp0T91/M4gLnwijI1kY5dGK2OwVlbbokMWmtFaE7UaFaVRrTw3WguLQSRD3HyHOxbjbWYHa9Hxx/
3b0a9R8dgMh+wAsUudyoXCaHpXoMdp93YbEgfFcCv6tZrrOKcI5JwNxeOOjSrDuhkG/qXo7sidCP
q1wOfCwstgMe4QJAeqPOUod9f7WvyFW5JRLxMoPqTkjBemtLR7Q5iJTS9Iv9PIkHf+c5Y5l+LPQm
mwIwuccu17k57LD+t6267bHpLTWHDgkqVBpoWaheeqlcD7v3mAmeGSrvOPnqnuDqRdsvM8G8mvyn
iUwgFagzkptotpe7jSkqp+nbxNBPLuGadgLrtrqNyIGiR5JRoW+nVPbpaQJ8tUagzkuX5RCqfcNc
avIgPkb1enyA/oiAlLQqX7UkMn9yisljYHq1zyhKPbQmO57x89/GJW3Khr8VnRtnHth8Ked93GE/
m3aFhW27P1WzH0EgWnRPtcs83SMm+w8NCzF+BrxhPR7fsIwJJqc4cFyYfr4QsUP+moW6A4N2avzl
ge28+mZYulGoGQcNslBkm7LCeCsjBq+z9VR+8aYs70UJZZU0Ze6Ks8fVixUaV/vs34v96BpDCuT4
rjNZVZAx1bDKxu4U9StLyrT8NGLFdkwvrS3+POlvu7o/KQR+fx2Tp84qDnxVupN/3g/OybQ2Lkge
KvyyAvhHt+5B2DKxZxawXPGTGt3US5m1FR1dxzHBCPBM1CK0V96+0JI5G415/KvS7Vc2Fq3sODpP
pZ8ybfBMr+MygbgcMnVWDQT+yfC934kyWVTlDc0UaYqQU7I7X3XsofLuux87T0HkKwpqpG2cTP0V
rpHzSM82b8LetQ7jhZz3x5Prk6RpgTjUBjuhapBYoMvXMAVrW2oz2alJmNuBFZx4WAYm6cjdrCmZ
xFJpZSUnUe6uziG+Kk1xMHAglseodSPQBw36C6jXwXfgPSWEFPVOoKH7cAbv+iR+CTA6vXfNSOER
iGktMxcS4M0KyxDTDeaQBUtXHs/3FnKZmeXJCw3hcDJjmWfBk6Gvcy/hmqLAPfs/v5HigcDMXw9w
w9IyuliuU4YLpBCWIky9awaG3EeKTqiCHMF+T5O1+TQzKKGnHC0HlCIE/8ZuF2EpnDDG9jtOB0KZ
KtyLP3Rf+c/7JVdUxk+pNpBKqNuFeUzjVcF8BpvQPd5M26yNLZel8ceOfV+OSOa2FcNALxUeb+qA
A0mokNz5azccqwFO3mRoKLPRQNA13ZKuxMPcVsl0lCtdr64p88AppEjv/I5Pg5ureV1gHeG6/ghZ
yng7rPPqe1aRM0nQWkrIuBoumjawK6rSevYFhstsdXfw51yroVH6ETrw9Bzs1ke1rN+RAB2tlupC
jHne1dPvxZGAoaAy+jPgw0cjKnI0CxY1eNISNF2oxfSqTLPZ0cTUqLnJDN4f2CXwfijNu+Hbf2Tv
rd0uwe4D6EdaWFVWcewadN1aAxLm1RY7bWgyP+gQQ711DgkjUCgD43+uFUxotM0KDLUnayQRxTq2
vhAQW31KMcxuiTE5rgGyNYx2f2le3yN2l7VvNPOI28KDoJ9L2Twv6xVFP8QbqpeASwbLXjL9EVGE
siDtOmV512gyB6V01MPQ2/BLqkb/1KlbXfPWFhf2C3WHE12PBuIK+mSqYGr5Ffl4G0lUZy+Vk7oS
ck3kBF2z2faG51bHeQ0zcYr+2yoiR2PVKdjOdIdl0ZljIPzKC47in0DRYZRWR+bCWVnfg0QLmwYO
FKJ8ffPmdmacs9/qoJfuI57eZsgH1w6fwRRvI7ZYvXC0v9ixQmkdluMpTN4pnQg8oOC19wgpH7Q+
bR7z7ZwOqnY7A7UHO72SJmTSfUXSv8dl6uXNEO5wUI9xULjoSTbmQvDi4hcFLa5s5VkLBl2u4Gkl
a+uIxCeaZhzccKX7mWzlrm7j/bfZNvyYOGXAUfFIaoLT16ZnlKrQMJOXqL2j2YDOWY4pla/J+Iw1
j40EELpkQGWfNapwTUlx2sq1pqfbeFC31NgryNDG+dPMkkJ986j7Y+It8a/vLUxjbBmClLU35Ksg
0MMgKi8giTQhXkeBAmt9zLTC4JvsPaJZIaU77IVTWy9uJLafjC3VfpfYds2SqNmKBdomY8fVkKFL
tsqQfCYSkIFV9lIgvlYekhSf4Ou8jckkOPS81qJ34l80kLb/Fscnn7R3yiIJq8wPfe+qmXVsteqC
ERQM0480lTuTIceMmD8rnfgOFDeO6QnoPvmredJfZFzvOI3DubCwMerECOvHtv7WxTSjNoVKjRlU
Sd6zhRfnrr8YSpYJolj5B3261fpibF0GZPSYFjKAtXiq/OB7pgFeJM/oX39R96bPzR6tqJgkFIui
/kKO1Nq6uTb5J2Qr9C7SAH1aEmFQH3n/VTRO7lMcE6UxmSqz6J6QvipX4M+aBIgzgcfK6aP9v82E
A2IHhePcrIB0/LZ6ZDhuLu2/vcq2ttaZ6eMG8htVVYgoaahZPg7ytKpeylfAjCnxICdHIecqhCOc
/8ZxuQ7KS5/Z9huVbtRFx1gah4B9QEIKkxvjCoBTLIPtsYO1HKV1RF2vgyxgVEvmMpXfhN8wajET
tx/NcaH6HLTkekM4o+3G3fBwxKW3CyrshxcF0cWMHQ/8nKAtqw2rs6Nu7UB4gjFxXgsmi5cCHVgj
5rW2vS2oPv9CpMKD0HSoST20aI7uWjfNKPFfzXphcAVECAZRp3HthEZvXyICjeQxVl1HbSkznaSJ
q7WUIJxkWzOaq+GHSwqJfZtAwpFtliGbXOUcA/uWx8/tGS/4oiFVkRYylXLgmsLkKUPp9iJ50cA9
2JWyWlozwiirKAPqZK2xnxcTMpB9kkfQIpyP/sZvNp1ttEr68HUUxF4Cq9YAXMPdA9QtH6TBKK2W
kvbH9e63hGb8nnAeA0GNO3v7FD302NC5N8SWHyIZBLW7ZyyFk4lmnbsqOgfWEUvQzo7yDg5nZk0x
4xonxYWO5udvQUOZCRecEbq+Xn9w0Ai1ZfnqGbXKAal9S7RfweHE4CbMeVlpI0r5poGzSjij41PS
u9mbJL0J2D41kdJXpR7FY8nptlmHrqDdCq+3YR/dyugWSyfEyvCa5ZTaHL4iaQYesPXq8GqIuuAS
jOBcjJyxnKcTJxnJk6qEQLFYiGX6mKZqpIct0rzom6VEoL3hXF/RZEMyDGowAD97gxDmxqY94rkB
DowUm4aeec+Gs/OmFHHfr3mdeUPBg3G3Dw6EWGZQurwImUlB95AR1hfhmAXQR1geZjZ0HyFqqeaS
KwVKQaSPLzDJwWK8GB+1HNEMxgKv/HeVUpKFwAb0zbT6206SyzfmteGPgGPDuQbrSYzx6DV/+inv
pJTU3t0emgbInTQY8SLV8eOSnUCkKoiBWCgvmgkLmt2oPbCKkBEmHN82PACf8ts+xmWx8SjQqVwj
hBi1nWFlZ1PV8YhlltKIbWRXmHnHRWv3o4098FRkJTqLLv7mS7yL0vP4juMnwPYXz/R1s7OUASG2
IEt9JfQPmgGiSLlomZWeOHIW3mgZPsKugXxKvlz692ywrOMy0FFzE5HDhsrlxWYWFkJ8WjePbmsu
A9UbofHSpuUl2U4t4bZVKARPh+Rp92G0VOtmEzTAFY9GdPbdGLIlnG+U+ysozHVppZ137Z8h8yMX
CJ7jVLL8GAbdxYSuWNHVZ6EnD8FRd5giygOUtVMAlnGyTPJxC9DVEk4wHvkdA07QDEo3T7C3huFV
KB2aFtUvV7uEmKJEqnPqdCJ2I2DVyXhB8bj0ppuOPFOfawCVqqGSIp4XnVxZm6Ik10Hc8sjCmFIC
PNxnoeDoMI2uTj0ayafpxBpfrl/o9P3Kv4xu0FRBATFpA5Gx/dsOm9pAiUcNJnmM0vb03OW0Ekc6
m0i5uSO673BOisrHZHYtEnWy1GFRJQZmNchi8VDEIteMmzRQX/6lQAyXHAEYPsftUzusROj9kN1g
j5j324D/LN9zvNtE7c/o2Rf0OKRiiQVkFtieyuvIvyIAEvbIHnnizl9MoiyLMZVreygF6NJ300EB
ZlP9IxV3bL99V7N0PykvnD8VLARy1h4vFvV7EYB/b30379PlLL85bO9oYlnxLlwR1zXQbME+59kc
B4XRK//f6VPoEFFrZphm1kCAoLAhYtUfNVO9QqXMY6JHEOV0hqNRYovSJ2Byl7epXR1lG4pOfbyh
pt0TxADN9dmCq/91d7jvMY0DcrzRZ4duOCqBz2sVifAoxS9X8IFHoNizwtMqMxktD0tbRpVburXF
33Du4MuS97ikXtueWuPFPiHVALJNCAaIUt4s2ck2xUCL/Mmfjkv0PjNx/FT1JmqIA1xwPDDG9lR6
nk4XX8XBC1pUOr70NVrmkaqQSi3dMjrUWObK8DZul0RBo6h1jjdzJEg2Eg27YK0yERWIJBsEy9xx
CN1BYiXEaV2Kf1vJRvxjZ6Z9BWGmBJUQfUDanvEryKVZitZJD9TiuSqSlHf86GYl6OaPEk+F8VKO
8vSQS8PwVhLxZeu/fnnPjzw+3vuWMbObFyw+qRUqtzHH/QojfoBK0LY1+XwGLUn5Tszp83w7hILx
r3fn0xcvSsl+ROwuZQu8qIJwdjoxhp9lP2lOo9QUTXfsME/4VgGpWqhgKiXZYgudd5q+C/8hncuX
PSxS/2yLxgzMs7GyNYXz3d8QBvUOJ2J8WD4QI3Y1jfusSdUMcgEYIw+2DqrI+9lmQW93kHpdAyC3
QJmbwY+bxJ4hp4Rz+7UW9U3AUlZ4OSB7ssD1aihL9y2+Pc8S3P4wfFdH4hCJ+so/hhhcSxKw57ns
Idq/XfH01SH3ck8CDLnHYeF0FjRXINGO8Npq16KwseIYjqD0iSalwy8HoJld5ABoSZvfHif+Snqi
eyN4hxZu7WDbW/TUkGBJkz8ochDx5wZRb26Z7wA8PD7mzgvmxhoZpwB3amkZyQDm+7xtcTmzzhUZ
ypDdBbE4ksji0seORhSfQW6Vv9gSWgS7UR9oVW8N1OsgkQXuYJZIyoQW8DK/hhBlisKkVJ0o3eBl
RPrrFi3+fm/azNmKe86smKpezWszGKzOb9Qx68GlbIydo0KwJqQH2xZHC1rncKrnA8kvk7oE9ea8
DL4BiFD1WqorksYAJqo4uRBN8YXj0yrxlboVD4wVCnNamEKvd6tLr0dHOuzSajikxhZRqvK3HjSw
YeHM8WovtejRbB7gOwE7JLS9p0rVb+ZaLjg9RuagwPQEzlToirPnf3nm7QSYDDhlT6oCpM2lvmJ0
hA8bXpexkvMfNFOqcuMxFskXiSfqLCYwbX3PcTld83jBGdBgRLEpAsuSbYgFoftJaHmC1r5Htrjg
ivFP2KmqWiswBXBAwKtEPx1Nja0J0jzkb2BGgCg82Bq6Bal5KgI81LnMWwQXFiW2bUVVr9BW8p/P
g0b/rGiLO4jZyXchxqLIc5wRVyiTOLJ2hQYSdh/gzKpCcJCSFfdN475N+Z22ekVkhc7S9cWhZqiR
8a6OlqruPgUub82/y96onbShoTlz/aLOdM+e8eqXZvJ7Td9ulFhSTJqhAScdW11AUCfavUuVj/ff
WzfXOvJfI8TcQiRtvzoKlTuuUjWR+QzlU8162cUwWPdJx0UdVfVUqLY0Ghiz9+aMczx0bTLuVzbg
sx4nuOP1ZfzNUWmvg2ivNSV9Djlo2g3eJtwqe832Ys4qRQCVxmiVjd/WsGBGuvZb/Vngvivmlz0F
TQ512DU6OmtmmgvKbH6TmNNd+5o0D342bI0sor5uAtry1F9GXbS0qzMuDlZZbjw4T4gigtXOU9cl
yy3lGOyt/WdosycBoZyRDYBnCo8CccBKdoo9ODLvjQjZhterc1UHBnO6wFOIx1Ns3VvfWJ+LhZ0O
hDmVFEPRBXGpLwuLNipg5ieSCIu+amVeHzF9Cj2UtIeIgdr8sj6aG7oajHL+ElcjNPAFgAqfV6nF
jAb0jXxdEZLErZHPCRbMCahjzHxpf3WVDJ9Kvtcy2rC2H9mxRhQArAIopx2CBm0NpKZBhTzb+3+5
czh9pby7qCAAVTaTTUDASXyFX1/LskNqVlbqW8JpPU3Gqrpiw3TJ2gVjm2WRHB2WiqA9ZmkEklxk
RUnRkDLla9Yv96wqqwyo17fZKuwAvjMxTVE/D0UKdtOIU4oA7+k9hnf4pnsooi2rh63+nZQGATZY
7mdVx9chnFny/YqQI/53Zl/HwfznVRbWvRQjBNAl1apFYjfjMOvZIHVVQFWIHJSzYkbn30gUuQvp
R6QLGHqifbHrUA23Qv/quIdEXibrC5dHPaMJ4EbWhjHB5G7OLwXEUlbT5DE+ajrH+7c5q6bWDiBu
4pP8MD7QSzpTQGOHhMoZcAJ84xHLUAYt6ljCaLWs8PmkL1LZ505N+2sZNUODnWQ/7OGNhO1z8cnR
NJsNFMyZcp9eL7Tpet4AtxbzfJHFbYYtyA+HCENuJra3Z9OEExsN7utvtHXhrNWQneq/PosHvJ5T
MSQKY5PeNJ4dq/mZTwN3CCnatmxETcDvLUM6Qg/09HnpaaKPxPNxjQ1c8WUhwCYFja5lJDzIX0AA
OLpIGNIerLjjK9oi4Yhx1rD33g1sj5mjL1/VtmUVYcrV1cyUZgmm3L6bnvT3Wc/nEvl1qMq2UWrh
3ltZFryzSqfjtD/P3MwEZdFUXnTSai7PEp8Erw+V+1/cERCWeHU+p67BMegEC+4XiOBHq2lhgxTp
Bn7aZEX47V/yAd/2h9eVRLspz+U779G01Vl8vhGc0b9LnJiBZTcngmtilvbbAD0+f/QDDVyjCf4f
jDdrtMI/HnlCpLOhmeSXh5hlo69p79ITgkAQaK5JNw0TFatAilZQv3tgZ+Zwq/Oenb9jZQjXmIH4
5c5qk3LYm2aMGpMv0yfH12fXiASMD+aWT2WDrBg2jThlaVVYLa55W86mweqtsI0xrkHAynUXHH1q
TwGtUp7/27Wsp3DTz2kJDX5QsBEc1j6yME03KfmTAe99zcvyWszsq3l98tQSwPgqL4Ir3cshf3ir
ZCYVkHGrtS3utfwyhMnUiCyjEfhOQ4y/2LhfrOKIxC4rjLeEEXe+gtUmLCM7+NsiaskaMwZdIezp
ZHkPcy5iC8JpKpwWBGNfcFe5fS1r4h6hdTT7LtTMUDD+lAX9GxpWAhColfKZDH60KM8Y0+TXic1d
fgF8Vxs2KTNucIcMlJa6+60mQsVKnVlSQS+rJ1rAOLxWFPLTJwolGfV+O/15s71pyvEG7S9cSSaY
cnORoV9UaWXhBbe+7g09g4NslufJMrKg+6uTPsYkSHFgAJobO2BE7ElSfndramA+IGoq1gm3Hv1t
9dzV3kAlyiXISQO2NdgIpkPOTh3caakR+8deSBxqKmgyhyxLUTgZN+rmJN7XnsiYe92djKnEnFY7
8byFZZ1LGm+RqNWRY3l/zI2frNzkTbxJB2xmMRnxQlo5wl7D/eix2zdSigBQqUgtAXgJiq8UVGXk
6VGpXUmGG3ZN0Dx+gSxbASalJa03sz7Mu54/sFjwrh1f26XsNOrxCHOrk4K2z5ETTlOCxa60my2M
cQZkAipKNRA0yNA7heF+oBqWWQW4hG3thxouiffl6os4cRFtBgQjhkN+CI1awRoonWAdianfrxaP
woaYGRlwvue9Jb2ik9ZyeSRerXeSaS3wgrPe8ZZkwvhEorITNtzH0OvXS/waJrKHRqDfOkHYmc71
cDniX1avYfFWhA54P7w9fEVD6+VeRfPd1M/KWnZlzDfK5ZPsAYHPNx5ec0by8ZSDyXSVl1y46L2s
Pr1b3UyEXJV3PM1UbvnQZux2IeAJhnfg5phpum5zL05JO5H+B+jmULfPOwEUPc+dhjgkum5FyUZy
cSzBWTuhhPjTBiT2kg1fKFJPnkDOMuzgNJEiQMUO/ILmHvI3Wb9Tec6fKB8mUq3tqCIQVw9gQ6lE
P9t+l0JYh16ro1t1OkUV5h0zL3OmgW1Isrvuh1cg+nlrvROQ5AHCPQEwqMqrEDUFuwJMQfyOgVXw
rcXDvwiM1NHIWyi9pBZiwJLc3ENWvfbbk6hrwKad6lK9BAvAMUVIidshb8WeLC8n+jnEVYJA3d4N
rVgF4Iy2kmFohpCmoKDlhuCCL6XMsYIGayDn+5ssKFinYaFW6yX6jgD9AYY849XueXplM6UoYfO7
/gdVDbqiQ68Jv6ipOlGHEvdYLQr1ccgYkYdeoPn8udENZ0AUhz08cbCvKyIU982cu81EWwAeJr2v
OqwvoTsLniELf43BnW7Dgrih6QiTEgSaUvu6tj16/ye1VBD4g+P0vCxKXAmYqN7+P6wo4yIDc0Fn
d4uDiVfrkx64Ji3/fAXlOlE2Y6nNcM42kEIzN/5Rinz1m76NLArvMTOH9K7DRdjpoTZfcI5Hp8bC
/46cYGWe8qSLLpoLoxCydodTXVmQmosv0Uj0f1ATheYZTaA+Z6/1AX6oSDP08tZGTKP/dbfPC1Jj
YHlm13nXefB4K9i5yDy3aP42E8ZDxXcMyHvuWrMkPo17lhd+t3Tgt1XmjFUnKO4Ftfp975lmZ7Gy
I3886Um4ngSKtoAx80isSqLzvG4DA+oR7R2ePalv23C6xJHYohdfi2mEiho6oktbCQBEbHM1KV13
MRX5espwZfDJkFI6TAPEk+/M7B6kLB+50plQ/t88OufueOeKhPh5PWZA7X6ZL9UvaYxq1Ev8b9Lu
chynmFKAEtqqz4wJPqEHVl0NWot60dAn+BEJNZfAzBB4BeF+tJtsIfggReg4QnxYh5VTKk2uOuaA
7Uj27XYohBgc/wYPUO1t4BuW5C6YjKset8TZgL5LziFkGiA2JZpJ3aSK/WNemc8J2GNx+w97uwHV
E3XjzK4kLzapzpCpAp7Q8GLjUbh8A8js2Vn692c9+huGbIX8x5WxekOmnRg/hUBI5eyKLA/CWLSz
IARyqA76+EzydFicbPtdVdRoPFaFKaIHTkapkDybxNAb89jLJPotXjcOw5CTBYFlnz1blSS2O9MV
d+kNJc3KL90B9ufyxXv8gO2ICcVh7Nq1ga8cGff6ZyZz3qUOgJJdhRgs7uWJp4OsCs7I6uxFqmj1
PP6HIYzNHIpk6At26Hu959cRj3xzOWzQRF56XWzUJ56ImCblRuNw/u3efC5AnfhpJdhePnzgTA1t
nOcHzSdxQYDzldBzB4G0FtK38CJfS7AoNKb1VesNjC3TZbviJjEhYEh04QLzcYySK9opc4QExHeH
st82ZdwnE5N1zBBGFwDnCqC6WraevzFxTi4csWhI1/LjJr1B4dU27zenHdMNlZxq5x0cOtujz4Xa
27zBc2QGTpFwEw/4PCBHx/WmMqhVcjOL58a2cDg1e/r4wrh6iH5fRDwtNv95aOK+eOVFQH5mHXsV
iYeFA1iW2n0POvP3W5prHh+y3gyO/7d2hgVMZWT90cBVSf+cwPvRaHDfXzEh3hvWXdG0YiHopVoM
pioxQPmwZyymzc5ewHabVkw6GKpmvlN7jJsBNikitJB7XV0HLqiW44lCjO+qWY9pC8nvdbn0eWfc
/42d6UuXRQhxGIe5H51XQ7l4/omkoQvLiVB3MZtxcbpIhV9SXI7KW9mB/YC3+Cdp5szFfE+YQri1
E/WGiqvxk84S0Ldq9rQqsHAcMa1XMme/FI7R+ahL1dtX39FsPMYaCrX5fojpHxWRVWEZrsyvtPDu
5Hw1+B9xpVnH5FswTSFSbTlGFXrBcFPW/T+weiZwLVO2VKBQ5WPexZGEnV4PXE7yEDurW0SFRBB1
bLQkL9KTGks41uEIZOyz0ipjjTcHqqc7KezYp6zNW1UvGLabmreFBF4t8LLmWuSPIssscNYITcbr
mfrTkFzliGoZhHcZRaYPXNNJ4QprI8S+msmn8QG7qE1ULGL0ilmmE1Naf8gThZQlMb5Q6K94fYWg
8X6+y7COABvFnY5g27iqS7lR1oEdXrI6rlls1/fqP4Nj6XHZj8W9apiS1PO+ZgfzcF0NORbZdFpT
rN9n6I7icikdzGfrlEAq8yPWZ8wJkEVFB5+uY7xRFJdITNETo3E2KY5qjTWFogf3CUb3+hWVppqS
YwtgmVUfeH1mR+c037IyCxX3I+KW2WpYUFqvOyJemQIYUgZ+flEHEYTYQvZD1sw8QgmyXzX9pZW/
1CWgjb/RHrG1+0AjukBtoTU6vKl4bP6FwKok0oPk2+9RD0JXYXIgx5gHjYZaBaXxE8s8SFvH7tu+
z/kQr1y7Es+VavUC+Cezr5JpwT9bF4JIs0xtm5E6hbjKclMvJTwbKkN1sN+nsvRkh/oLLjEKFgz/
HAspOwFo8qQ8FabHm1oEQLRO6kQ0ZzpViijORdRXnzrIyzZbopFcu+Mr5DrRQVHdFK62cB+jy+Bf
F1Y9iaqhDfZpFAPZbtQju3TTXlDRydXW2/R1A8IcpUIGFCeFyYJjyS7PplLBc162N0VtGp3aTpKr
MMNE1WYP4mTLdoYqUKZWAbgAxrN2yf6+VnffN7pJTqa8OeJwKlnpuOWi9Ur+3mYppfw9w/8S1YVs
NYSQ7iy2hBobS34S6y0uKMGD1SaJtjxEEBMPX37SHrOU96D/FFjHe2EAhVtmqSMl9ANimlMVy/Px
ldWZ+GSHwjRcxxA8b4DLDyTBT0AdkyEhy7s2PWpdxhzWJ56tSSjPzoQJuWODie8VrBWOrqddiJIw
CVTnWlTHktYpyIevdRufwCPjyhQwL17aVQxpymeKuSP6J6FFhXXpQGDP9oD9D/XwDDwfIPW8LyeW
6K2RSWKarkm7h5d6cTx5VUzWqNZGGHwuoeFw84aR1Ii5ADhFWFqjVaAZhUfj49KF7i9GbuDI/E7T
p0pi9II9mh+fAED5g+TDC0HXo+jy7VHmWdAr1dK74ZyBc0YptrUPewBt8nBOTe45jwIMxbAQTER5
cMLTm7Z47hRowpj3v7DOznFtD6r02fV1IqvgerMC+rhqMq+XhQ3CnSHadfyzRIuaGeGVf9jkLBR6
DcQTLwhzzEh1CWF1VVeIYU8Z7wJ4JXuSSch7HzY4TqiPlGG6tzvl8faz3qjjGoBkRfSVa5YGh6oB
dfQ3nDXHSkyT0fSGYgaoltzJcuPIKzdRCPIx/w70izHcr46CMX4hVmhmuEeYdmCIciKP0S5+dMjo
sJSeI9ytaeLEhW21vLFSWDDfQRvgEa+GA9rw8eGIK0Ga0aC7QMF8EzNFgc1P8ASFkNQqA3+fHlDv
YMYxRc4AmZ40BgU4gOUeOvW1A8bs7CHjRtXcd+deAtRxRf7jc6BkwNLwFIXK8OQncou3c5UPolLC
3GwkkhskehnOGOMZq+H23myuO5FuJkMyU8vWof/XpXgF1MfUm8ibwd9Sqski27uh2ljJuB6fkF1u
bkHWtmztGbSdZRUgkCInAI6/f+4ZkWurQl0203yH1Z9/CpxI9EJSC+uz4p41AstuZMDwk+dizvXQ
nglW1oQZwRz7BFlv0dPlwtnuv5l/PsxviNxv9dym4V4shmAUjoArQy5yLGFFUq9h11BGlOPVUqpb
hCHfLrz43+Qi/OmFxfaOwwYTRSmNQxOWnZ4QdVyPNcJwh/hiTaqIIfE+2gxEtLLb16/oyCwvkjM0
x1JaG57brxnX/+eQcRD/yL4mIKO/gPVV1Pvp7AwmpXy6j+MjqPcn9NIzbon/X076WkKbY3FRsFlU
WSU9os6Ow8sA24yNjdErlG8/y5030/yYbVbmJETmhzNcWzHzLBLCEHtjK2rw1GtNQ2XKZNkslmOL
KXMiwpiEjnQX1suIgMgDWn/29H+3cnKAbnyIuJHlSSK1NAywkiEH13nL/RElSrti8at4obQF3gCM
89k86Zlhi5bCBguGndSZ5yOTupVXsjxEQ4DSd89+76usYNzASAE4G0PsZpUB80BkcMCQm+zKshj9
6gj483D8vFqeFCxhFGJ5rOzPIue+iK93d3h89N/X5aFOVSv6PDksutqbgbYbuxHrHnsIGccTIlPA
FHFI/CEgPtbbG/xIdmRa/yVrGkMNYWAPFupQ7vTkMWbXH5JzCSGoLKziQyVdpulfAACP0WqaIhY/
LbX3BzlXU8h0KbHekAltLzofC10lUHmyJ40UMQXp7Haqt1AAeoVm75BfZ/NnFjvjAEieXoPTGVe6
rRORaKz/twcvas1wFjZhmQHlgnkwRPckF47E0cOOiUTuixRqQVTfOamazp9PtX2TYKqwDacanZiq
99e1GRa3vRGQzSEZMkX6oO7QmeBHrqtxONEPGkgd0WgL6O9jrj6ufAHYkRh3j/vWtMjV63Eiic7E
5qH4tr44sb65saApimkKHF/xGplQwluYSL8JI4ffBFiVUXwaK7igtFZmhMvYjcx0c25h1POW9N7A
5pwNQXL3NNVzwRA9fnywR9a+in3uO9MWvOMEPwihNRhHDnx2E/4jszjzxMZl7Q6T6iUFl5CTiAtK
cTg0P33dX2zGRW9o+gNVhmThR6FGTuLzP5NY+Obm8RrRXX7CtkyV6oTOzubFAKzT+8G4fUBsN1Bq
KVbHedaYfywqjLRSHHg33Ms6tsMhBNfA92uhVbaXKC1BuNW9L+GYohsVyq6pUdjezUiIcuR9GrGm
UxlfbgFRHC8KAoODOXFGIQ+N8jwvNKMAffZiuDBOFgildyKYKD7t0wez9LEwuav5hFzhAF07lttl
pun3TFNZHTW1XuSOiqSON5Zb3HqWVwtTvbT8XAn9A1Vsv+ue6Nu3d3wO2o8/j6VZs6dDA/PnQHlr
oTtTIyXTswyDJhAqCfPX1NF8Zcx99TTK5Dl+AoA/9xULBMUH1PbUhm5QCLnaIS1zJj6hoiUnTGIK
gh5DvBC6+nwtbdY66SJpuqgeN5eQdLsK8l7JcKbBSvnFSNl6gHYhdKen2D/xRDy3IunnA92f4HQr
OlFe50LU0QReXUNL0ESGqCk3DqCxSRIomf0vo9CyiI93BptwwSf1kwdaNLP7uZNytRYqbYqzOlkq
BV07yMoO2+PngRzmDVBsNb4rEEto8wO63OOIR7NsG9/IbVd11NCUx4SmfMC+Gci3756xQeaagvJc
kmol23AOnz1UYAYmDD1Vt1SsvVUpdZ7EySpCcVAl3iND5T9HA7GTNpauBoLtUSHY1af+LMgTCdns
/P6gjc+7xuDbYjUp/uNK6bLCHN3VnbJgFExWpVtHq1Ci+SO+H5TN9iY1Gj2qjOu1vpFVgKhk5ktp
Kxy6jFIVetDTGPT/Fh9fT+ddFXMdVF1BCho+k2ezHstbjPJS6HiZPUY6zLtKMR/fiyfExIWCQO79
nmjMi7C1To6+vFSRcRjujFPCc8j9d4Oyij6PJKzogVVsABT5vkHLkkLJ75wmd5Jamx3oGgnrkrTn
R79POEQgA/ievghHMNvbt7N5lwzDQ4IXZFXDEdlRiG03SuPYiw7QfpDvAQtk6imyP6YwUDrahyGk
vKlt2uJr9Rkdq1ntUkbOY8ujZ3UCrcypd7gxnsT7aXvad6fNPARmVq7RzqoYUmsypjXjD+IZ878g
CZ7fMGn2EbElN2I82T2yS3rHRV+OlHb/Y8F8OAi9ZV17DpVoBK16noSbuiunokvz3FMxWjLeRknb
F2hfbDgLGocEvrHlHYPVn3CfiNEwDrGf1KaRDDe7u2JzQF3MEq56Xcx6/oHkadt11HmhZoP9+1oL
EQ32VwLFOjMBQlOyTJ4sBeKN3lyCfzL5n3mFpxXD0cqJJnaJnZbl4qQFHNWy91oAzZbYd8nI6GcS
xYVqr06otQBL5E/DrWsl1Whs6uhfY/KNFAGS8/73XaliR/iTaDsJxiN/cxSSuhvQtyi6NTqVnSjo
YuRz7Dz3MrDxEfR4HvsZ9mPf4gw+hN0PrrXf/4GvxAcutcrBzagDAFjoiYV1FgAJvpxm8eMLEkvS
oLam32NNqG0POdJ+8AcUaccemYl3vzQ+xtYVL0RcY/bE9KsJpJKp+e4QjJ7BfwZsEedkvD57e2k8
uU4U7ugkm848SzVTWQyVZexnJwcSS3FrBciR2WYNqXmPwYAc/x8V2k7cXeJVyyTr0smG2G7DLXry
8ejL13o73iXY5QIgOV7zeEi4HIj7WsLRx47Aly4mZpq45S2v6nG3pDW7VxIs9bgz59FYUq3UrULM
HbPtmPCvOwCzQyswTjGG1FNq5KOe738DYi2kF5TlTZh0djJmI7VZObweiYhHTzU+HYQYBrSw4rK4
0FejbR886mln2FOHinHPcfrANXg9o10RWnd6gZrh5NS0odMdMT9j6VoDnqMJXWMnt7qC8gk/rE9d
Vpmi1nygf74NClV0k2az/cEHEtvOdv6lZ1z7aCvGy6EK5ywIlqZIi8+qwujCfnvoKmTP8GqZybCF
bufLRCAxhEt/zby+WdiZf8dxkePBV+fHg8+POZR5rpHFYjkqXFDJkRLNPYm89De0mfyqi8FCpEEU
yHIon1/PD5HaIeml9YJuaahlONlyLUY7qeR11skQitl3fdiiVlLRLfkD3wRQnmoK6UPmZOlTmvk2
T1L1oIYPgdPfj8E8gbk395rEUUkp6b1iV4IBSUoW5ka8flFndg7MAqM70zBnnwMU5yWZQ4LGW+bG
sZWFk5ztbMEg5aJTrU5b7gWw5IDUjPJZ6yVk/fIauQhvst/RYY2iR15+CECxEz8PdHzy2JR1gCRm
iPurAvzjhx9lpO2PW8Y1zFcJjNDcnP6i17drcbTiNAh28S1/Zw/Gr9PR/6tBKBA3b623WqiBzJXM
lRolXoUVNzPA77mqlhq7OxMgLYWWHpzcFdM+9sJwhql8JGUpwr9SLMKPoqCGWWEszmXgVc3M0/d3
xkgA/maL801fwUHbXwN3gOLphH7WFj9QuR7iM4Mx7r80uhgaketJqHYjAptAwwekFsefW3DUvwMu
MfNNHauTq9KT1cdxzhaM8hZDbu1JLzdgErUqm7jReGiEG3sL2y2v/ac+uxdt8qQdTykXUWEqLJW2
BT6DpNC2xEjDXez5kQU4t8mPVzX1mRstdYXNHpu83hwRiGiI0HAP6Q3ujQqv63f9z9tkK4Jus/bn
09Tkwmraz0Mkv/pHJmmF7tYmzlN3GeBoZ0NzCyWf3Q6fLB4gWK3PrDqSNJXn4q1g4Tq3f1Mc/3kl
atN2ysLfpgVt8UwsSMLxTQcT7/TAq6verUM/3RL4KzZCUW1mhDW51DQ+R16Mqbx7SiMfm9CuZf/V
LVQ4xc+kABz4cvufm+O9sphXo2wFVtX6izPf5QYGpMoyM0Rr9dT/YwJ4TamEEYm0cMIvtNcBZ/Mj
9W9FN2kxzrKFmjgrEbQ0IJSIjzsNoPAtGIyR7HxUJSJQbbGRDzH7nRYX6/diBOgPvdDM3F2WM0/O
ZIJJMfBXqY85dJnuurpH2JpUcK1K2u5oCPdR3bxXhHo6I7baLDpOOnoXs4jKnu1g/5Cq0cli5GkF
Ovr47zbkHUCWsGiR/ld4htvtW+ALvgvokAg54EjhzIYz1AMtOLMQlqZ9FcijKJiiOPM1u2evgFX1
cz1i8/x0oFdtavpx9ES1IiyyIzge6218HNXaGxeUZ1zKBCNBaYcVLz1GWc+AqpNRzJQYdfhB4M6c
d+ZW6NiReUOePXqwRpTWOPv5Hm6ond2bdj6unDHgIngKhlwtGizedQgQje6yF0z2VgxscK9R14jC
dVJNxh4MhHY+yecy0H7B6yYz2p/74BE5nngP5BvbipnWyzju7V6olhJRiITov0zU7hiKWIhO3ETc
OQUcmlsGLyt3YDkTtBbbvrrcDDqVyg0CROR9oXDJ23pRy2Sv6vUconbk6s87n0ZxRUyRX8vI6tYW
TvvW16YG75SoM/PQeWjsvqvpMfKv2+/EI2YV2+273J69ixLQ8t5JoB5V75WVN+fVv2EdbcTjSWXX
FFbK94sVD/WY7PnhecZT/BobQUyJPsQjSbJA2w3hZwhWfoyyyBAYJ5zp3UxCkVx+qM5UpNc52Fcq
IOfKFxX1OGn9MQqjm39JzvPERCd3xX1kGKHuItUhuaXVh3vtR22ObNveQnb+s/mbk7j7WRc5+cbU
th7uOZ84gLNFm5B5AGqbrcxfzS8aJuXwfNATJCHLmUKGg8WZ4S2jC0zmwN5DrhP/WQykILg0C0ut
nQyeOJKiR4jUn5SyPiJ7BUqVrl4RKwn8z/8X2UpUIF3OmKU6b6geH6gbSubO7LqWuRNK+YEts+/e
ba9RB753A6wOerWTYVL9ZL3+kbLLOLLZalfr6WkAVH3i6IjKfRoo5TKf+0cJqbT9Of3mcjXWky8A
QwQ5hJtLqwbSWSEWtIQhbEPv292/BhNRkyFgChXcNnI6k33a1mZ324bTu3Ni/GGdhPQpprncZRpc
qZ2iyD+056tIsgL85MX/0uQQ1mfKyr+McpYErdnVRnQtfVkhhqbDsoa41NdrrzQGCQpF6BF+mMmL
5GTSS7cAQFZbtJ6/B65qzJm2YsfM682Bhj8r/07UvjoaZbgSvuSWklvYwDM+RAKSFVwG4Y0Of4eZ
tU1McZ0RcBxqgl+SZGWSOsBxVc7PxGIAGWb2UYw3I83uDRWHeulqYLZfPLVCRtJi7BV5ZuSexhrv
VHxmj5oKn2mpSqX6L+yLeQmXHOwASOTaOmFKnzASo4UaH+XKMlnyjyGgW+jMenwQ823ZVFTpfLM1
ofKB8JgmTP8rVxoJ026v7So8FEM2/dNqSmdJa4CPzIdfY8SBCSR0JH+YtXmATpk2t+i+YsfKoJvx
CPvJ93GPW34QTSrvHszPqibcufRyqSHrgRvYnzRw8m5QnHg3xB+OqOGgeBuY6djY0VlGu+YYk0wD
A2GF7w+0h28LHEuOKKJdI5yCeXA0xB115AduyMt/9gt+4NqCaUB2awDbBX9uBa1eFq3oS+wbqEXB
xpDbCu7BUH0A6rrlIGpQg2so71v0eipgjwTl7KrwzgBAABZugAiGdVIMSu3hLGd5MS28XIOagtW+
XG3HxNn0IK75XOh+ab9YygBVAsPjNdbmc9FSzYgGfGvT1tCCy1U10bdpBfNEckpVLXyHkHKPw5eM
PbIzQbmaoqwiCr3KTMy5DUtUEoUAQqMzS+em8LpI+5bZ2qNBxcQP8zQbaORAR4UUmI33SSVTojz2
vJgYbaRU9jFV1In4p4NGWt7XgjDPl2WLEmuDyhzEqg8pQBsS1fy2CwTpr/EIYiRxCD4OblcaFsev
ts5Volf0YBurXrt+Et/DZTT6wFqjs+NVlMEUs2LI9mHiG7PB0JCZqiGMIiPCR11icLbzAa0QmePJ
nzIrQnLZv2/RFNb8r+49yiROnNDfwHP/ssH3vLr2oU8lo0I2e9UTaR7YyACS99TXTtxmdXtQte3h
xPRWiJcjQLnhEjlj0J00gbhsKntSemcL0bQj//okn0kTyh77q6chQAj0ATuR4jaND8EtxBu5sYCT
oIFHpbCqWLLhzMVlRR/DbqrcVKB3GWFddnTJYT/FmuBOiUbbhykASW7QlmxXkfGp83Z5oNkldH9J
o/AJpyJvssxBScvtxvcebewxOUMO99i0ME695TXtZnR6rsbM0G2NHOArktQ+bcX/Kd9c7bcf8Zrz
beT2yExw3NaRaVZF39PfGBdr7hnvG2Cz8GH4jfcao10hIYiAP6SVH7x2CTczcxTWEbUOXWdV/bXb
AcNC2arzR0C5tBMf6HTRN5Mgroeadsek7Pze8NbAoBu6Z2LZgmipqgEQg+TWGVG76jLPaf8x829i
Mcd9E/vsELxPJTT0GBHzEgjvkC417U7XMEUkrMhLfYt48rSPFMXzMuxYmCIqYtmkAtfsTrVKQCaF
7E4yk5sw1Yq/ED/TaYcTKYHYXqgReMsavgCHg0WjXl5+05jJgnPlUz4n3E1Xvm7GlUUgns1FComo
druOCEdpB8QcWBQ2RcOQbhbhyjtbswq34c4RvKZTqEo9Pp+bW2jxBfv8uGbEKaFuq33Mbb8a0pxB
v/U+9lqSxVk4ocSERHiAZFcg0grArKE2VZy7T3Bccn/Lj4FIgCEpksp+1C74uriyLPYM6axx5ufy
L/75Qxi1et3GCHHqaiMUgdiwR/25eZaYTkl631+86X47b/606CNHVNtFwZc/c5l4Gf4ASSzSz1nl
vlVakJqVNUayHh3q7s/OWjl2WQjodhpk0/Di+SrdMn5TCYPeMUQtqjBUK8s2gX+avfBSKZAlMqmz
MRtprAw+KLL1Y/Hhc5LbtpLvePbmRzYFJUd5a0ra/MDXKpdACDhxNKjON10p94v56DCULyVJpYIN
S7vTMXqh1qb4YeAilVLsSgJJByBi8QmLRNK2jzKD73AoV9qi7+5k3ssJmmpwhKq5eOFT+4j+wzmL
ZNVF7mchln0xCZZfbmQNgJreR/WNBwF41ERT6G1wQcojxIC2HddscvtsMYWk3vioV/dIyRF2ZBOM
VbmsK5TzPCEojntD1GVTA8qJa2OxaUrkRGasO5hSj/9nhidxQUa4uXw6xPj7mkYIRwYcA8QGu7jw
wP3Az1tGTrdpgPd2u1PmxEI7fJHOGYl+9oWHYol35/wtEla/FPSBrkmoQnRELC6KnOn2rZ1u+p++
P919vnE7OuqJv7WuNEqtoon8fZeYATAGt0TLp3cmd7nhQlliTd2Pr2YZyFqDYSL8Ap8v2ZUdcXRz
cY31i4tNr5qeWJmpUm+egEGPLyJmSDFfM30llMUP9xm05cjZNViVPZIVnHuGYD2nXjP2HGIbwmEq
Cgg1CFalQILJd+SBA5os2/jA9OvDKV5gyBCWzlznkJoEJVqF8NnUXO2TmOm6q8oX5+prCcBFZjua
YUNUE8Zu2K0ubjq29Oiw/ZL6uCb8bXNzRlpsNOhv5I9fKYIwA4TbIlQed4WU7p2GFk764aySGvZK
iCPm911ISV4EJ8HnESKXo7bQdh9jdQ2xFmYs82PRQrDVcLBA/8PcELM/MCNeHVIqJHPJl7dl4okR
sw7h1yB4NiX/WjoRtMqwzrF8zGuVUVDzACafAeCbUGd2HClvmoOV+Dp8CWsXq3CBJ5Jon1ZPofI1
JwW99lzhs6jsnB1c9NXxWg7VyU60ZIWvmLXhzkNS8e3wfy5f1k6EeMf61IGbFHmDMdqIIK30ko21
hvD/fExr5CHkGFFxL0VHl9tRgSmVHJOJ011NEAx/QgwANWQmJXma6sxAlVYSzEhqzyaU/vDzhs83
IRhGoIVRRk8jofVp99K69cx8bTVOckXkAxtSRUUT4zgihTLRgDikrqUvqJC5PwxcNWr/8iirXWtT
tBdVs6IcEK1r37aIdZ0lPzRXE8Y/gBMkso1Zl9XWpwn3xzwOp/XpPVm3IYQe7McZHtig6+sOOlZ9
JLC3w30e6KetitxiilI83qE1YI1wIKTsV847YwI2wm/lsucR7gRVhSXjUAurNmCkb6D1SOPSoIfn
+AGxrQd/f9EGSs0YVidFRJ8lHxciZDE+mGja4PD+8bYT/FeGXeVxlRDKLWPP+eDVI8L+DZSf/XDq
bcwSroLX6qdB8bUmJVazVDpJOeEhcdGp8/OBg+wigmLVvGzH9Im5PZqoGJenIVD9KjJcujF/lvnM
S4ygoorSm1ExhL2lEqB5FN/+CLwPGyI8pWQt8pOZLO541j9iaPnQrRuPpP38d7rIo1fZ6/DHUPcX
qJfNtrk13JWM6Ml0yQanCtQHj4oQ8RQ1nggI+1IZjVvDJA7opxTX0UT63rVD5sVvW2597Rf4uuxw
D8A57WBQpChRs0RBS/gcEO+BPb78Sidq1+tT9Kr0BCjY8mAe27N9ZvwU4+UNG97vxkXfTMWtu5pt
LgG12sxcmBLVn9aYd/J2TQnD6AP2a8whdd+9xMCtAgwOV2fGN3IYgoYBODwCb+2pXPhDJUZWJYLA
h1V7R+AHW3f91eAnEXk/HcH2/b+9GSC77ObYwfharoucQWSfOHe5UWIvJkgG/oV1fjxhRiJKXoIs
cuJyKydNxdTFgEXDbK95hc1HePkr+btbAY5fGXl4Mq7edipl5CuLt+5O4erAKPDR9PwnL+G+Pz1Z
7bDqAFNfW+6a9sfYSrSbO8fWwb2oDAQC+jVRwodUbWVfu2atjh4cJstSV+wvOVqC8F0g+EdBOs2k
qG/hGZGTklBXo+hbDsLeNPEvX0f3ZIbzSSjSwclAi05Enx+cYxR+PeWT20d5xEQceaZcobT1oOxm
2uS2L7HXFGiq3+rQB7ThS/jOXUPsE8Oul/UXuGuYnX56SIiYsPYnDhtTqnSftlpXrS2opJFYoGh6
PdNtKENCbBwwU/MrEGLEunnZn3jbISJEnkc3CWK/goG+pevTmu1mOV9B/P6e9Jk6DQ2pfVzaHdzr
NA5WdrehamxRxQAW93Ee2XyBjWq3OhH6Ke/pisNEUhUrS54hBoveEmA9y5br4HpM+0vhIKLax694
zgfqAyQ2IiSJHK/xJv6VkDFaHOg2Ng5Am3H2f5L6glDcLhtNNb+j4R0bdqb4H72jU5yNSadbTqBZ
uumHCy9BNq3QbwzuE1dJf7qmN2oEkZFG4IiBxTxTQTzWkCgQ2M9/Ih3yafynMwpcC+a/pVBDLRjT
Ta9uFtjkbIu423etemQ+zEaOpD/1ioRGXdOZk/nK8nY5DzChLkg/ZLLyQ563IPD5H1A73b8s2ihV
NOCluYnT2Ex5PBRrFPFRr1a+hqo5ZyVLh0P/KbhpfHojeHH9fxCN3fdrXFpCtHmv0BUjuD+QXIQJ
OUMT1hDx/Udaseb4+kqzLn1bTuyNDqvuXx/KkXKKt9BWy+GbUhW5/mKtSZHufJSpGmpT+/G3vYMY
+P5tLNbLHsN6cFfcAbVeYurCySE1jDYtKsNgmy9QPIP0hn9f1JWBMKwxMs7tZo615Mou5caixazL
Ku37czjO6+G007tpiBAs/tXQgCRGYBaK04qPfPUmwo9qHBLOYhH59C5ezr5OfVGSGY5CN0TfFiU2
zapHvVU1mGorGddSkve98YFmO0LiSrXHr9JilgjFx/+/lQxJ4SfGJ3/imdoM1mpIZJ35DgsBz9h8
JcfEKoqfbUUADyEniev+fbSInPZKoQkV6HnDQq5fgF3Fd9hhiFOaJVS/bNTh6gRGr+U2OIa3GekD
lu+RiO6RPKR9LgT4Upt9XOd8qpgoEFktbQmCkZ4QD5HOZpBte9ykN3325R5C2DmpNta8o16q6nd3
tBkDjgiiqNMkIdA5sbKnOm88IhP7AVJ3Jm1JtC129SPxcnqp5PzyZIA/8rLRmugllC86XjrloABJ
UL0M17xV4QRdKm7blzeq4BIGi90QFHARYV+61onewhjCnNTi46MAOPu5zgZOA+gNder99Nl2quEH
9lLZP6TuzwiIE+SPffO5D1UyqSEBsGYc6f6IIzHgG2G3ERGSRwJtpapzZb4HAkvMWLt/gPeVtgPP
2haXwsxUr/Ojzg6QW3uk6Mw/ZndVpswAYi7CU8C9EkdZnBDyl+29inQ5z9ZMqt8xT8NCCW2BZMNk
0HwjjFT86Zv5oyKHJ4HwkjOsflB/hem5l16KJV4SKV/wIr6RYDz5c21v76RtHstIi6OloK+HvTEA
dy1/X3L8chW9zs/tXK5zqjZW1Jv9xn5tmcpNERbh74sPke/TExTfrGx6UKSOr44ujG+NoF7yxhnP
JkdSZQ4f+Ue3EoxG7m3r9YofaXWCuCHhdmgtvi5eSzSWKBJF0Ih/XbqzvXXhDVVaneu0nVpRPpnt
v4EC3p8j77Ac2823qRgGiM6pDScNK5g0rFCmSQFwcHh7rdpNuqG1bK0VkMoMx/S6BuaeItTqxi7w
aN4icgxKlEikSS4QAsFg2UqICsU0tDreujonGk0AB1UQFLeeeIi6ATlXFkss3L0Zk9Py1mO8F9jT
rrqV/n6wW26JOFz64W+FSXOObf1gbtuyzZKbwp0m+6u9WoK2naSvy1KUisH8Z4mSAOIYtZm9/5OS
17X9ACHkEM7cp3E0AelgSlU0EOXgVgqsuAES5GRpH/Jkpq//zZdtJgp1Sh2ErIdZ/FYI642L3PZr
ow9xPmJazvWlfMVB57WQlQci1eR9PrXOjflYTTdj6DoTVLTOBVjBkiHZCi6imO9P00nXV/c/wNX7
h7BjsQIp/R5fYmLcgaa0p2CSkpICTneAr6EbJPm+fkYAKxTAEhUZKQlecCVtR6a8EwVPAaXfI/hE
2jkv5aVTiMFRrhGSO1yPBuRXjrylTgFJyxsvsygoOh3kqDdiaHguQ3haaheqvUwhBylO3tCX22VZ
LST0TRq/OUjVGMScOh9v3NpL9pxTeLRsT1Xp1r1uPgQ7Yxri88WNEIqjKCT9wD6uGd6m0QRXu4VS
QLKd6kxCZQYN37S7NTWTht3DeiotGeni257kAilmiXJ90s6TJyVVd6bTh0dOzR1ZcUgnNeRQx/+P
H1/JM2ob8FgBkNmvX3cc5vargFi9/wolurH9NMK/RdzOXQgssZkrlJxCyIgByttylwL8jhuZsW7u
ZQx/v8o+huxKTTLKP+AIEWBfoSQhNuBfQZJFUIqwExPsUB6WMK2R6vxIXqjCQ/d0m3+JBBwQ+nTk
fnSKnhmxnfbAOHp7/K/7y54ecSWe7IkdhAilpxk4OfFKeubQN7qlruxYnyfUsQb4LfIGx+k21wjt
8Ga3YGpXwhDQPqgiVxstCmHDmEOLUTlqR2Zs2q+hmzk/ptGViysc+/UlwiTstK2QrkAXRS/Gb1PC
VYrOOf2wwNKyBuQnVQ+4UtbklYm/jn/jyBJYhOmoaeJrrBfJ8nOGPKSQT/ZkzCm+hgIFRnifkyxm
CJ4iqLnoAJhx0Ia+HZBuwtHb3dT5P7lBny0WO2boehR9QoAwGI5wii/Oaf+0tO8bCEJa+HW10AVa
x/ynnmtyddg4Xm2Y+FBM5JlRwi5xMQ4jdbuFrDuuonV32evv4BMPH0cGCslEP7+MDndkw6BnC/M2
kFTgNWaumL8TrH0aWMtsmyvx5IirUIBoqVXdMCEf/onI5Uf6bIvXyaGNAq2jbVGG8vS1q4Q7LgZf
kVM1AeMQLDBCgh8KAPz7t285qMXAIWPgi2Z7EE9uIAOE/0/IbpKZg+09A0ewjPno65HIveiO70y6
ZWkF+++XwN2ZSzr9LLbm7uul3vzfCJijcVJL73mUp+2YoxC2pqWXrqyEEDeoPY7TbJIlt0lG4K9x
enS1aOXgKHbIXEUiwyWVgaSdpYSU52+tET8lQ2Rk8dZHj2XLurjBG8t3ZLHGWlrxnnIFqnIhIWrh
/AOTCr6jJG3dFKH2a0o5idR4QEkh9oRIV1Xkkrh2jRKFeDQaQfuYY52PiXV+DQivvsgDDwhjjxJy
9mGCz41pDztlTdRoclarx574lIp4IwVKSpeENPNfv8JC458No79lL4paKdJisRfUPHMSgcvmo39T
L++JzIKXvCfTeQ0nO2dWSTWb2D/4NP5lHdDxtfCyfuSzlqAUnhXsu8GBaJVjWdObxtFTn0+HvEvj
9yti8Y2xdW4WTsjhv7Nz7AE8jVU5QFOVF5LSrsKAKV0ToiXHjiLaI1qWIpNkhTEq1FMoGvYrtr6r
NjvHttz0pdu9fNW7NV2LVDr5s6AuG1pWdrAKN7w+53FpBINfzDyOOfpDI1zh07Y4kkeA6LtctvmM
Y+sf3LfbYfycjFBO/3MkTPqYH/ZwjBxsY2I4mtfYvn+1P0Ap5N8tHOeTU9Xw3XvRGcfmEg5a5gLx
+zkcAZ78MY+Kd1eeaiHmRsU4aWXzDuGIol2N8g07fLounHVcVXbKq1FqPhMMGA+EBiP5iPDpF7DF
V0RE6AM7p1QWAmXDVN/4pbr68qxBdx8RsALI+jC410/HdWjRAy7yj9k2Qbp/9aPOQsg6+CGNFH6f
fOcT0G23T5Hm8aONJDzQzI/uxEreGdwtuBtHbGJ6mjRjBpkNR5HccbfG8kcu8C2jlgyOpvUcAucS
DmsVfoYMvRD8yFtI2Ei2JKdZ+O2F+glVtjd1em304trZc9/HJ4KhyPeVJXvu7/kxS+HT9PDixMzr
0m+XEYmULFmulNnTjDK0Y2Kg0ZCDTLaQK07p46Zd5Tzy1/fvIXNnNY/fs9jFqqDJiMQ7WwbdFKON
ekJZAXd5RiAeCJP5UMsN3HxxajOp0etgzQmvATQwRBAQNN0FQzshvqoHpSt5pZVNGXUipvsR+YUI
Wl51IKEyLITtwoU3gTTrhLUKuw8oi3ZrrHiX7VOx/TU6VhYakebUuQbGA9w2FIiVqKTIjgJ/S120
u6aTdX1KGrw8zmxV7gbNzq8sTc4ihoC2ui4xlWzSSoqfpX17RQ0MeyRqIckheM4tXqJA5PbLIHrf
cyEWmny5ziehAJhoKgdag5w/AZC8qLyEI0ENOgVgj1hyOGnAmkdd2lZ8ibHS6BqZ7wgykozXiSwz
p86+LD7Qwp00tpANhE+ELBE1B9uu5AxChXbj3nqFF0ErU6FjRj5xmICyAwBCXu83VWOYS24m16jr
Yrg7ag0zQcmI7myN7HmQl88laSfyIFJA/lDekHW5fr3f10Wex8RrtpvMkAIKHBE660zghZJzCOUl
pGpr/YHIN/iVxpQ52QyBa5kGx5RjYGU/2Z1b6Srq4q4wk9IfjdaT+qEb0fKWsCzCYM0eJNPofLXf
z1MORqlsAoBx5qDwRW17eU2FJYlNhLqNiim41W8kIWoAXHZZKF6Y8TfdpeDCZVMQ8PXSQYnasaZT
UGu/uxSxtZdnaLsluIGsEp2HEQigQJra1y71RPYzT6smh2FR4VOuNPaDOhZrt1o0irufV1PzgzfN
8/lyutioK417EInDkNjXxOKuba0d7Z0Rz8bciFKWSzBK32WTWeYdiFSLGMaxdD+GW+16/uyF13sI
zCooBs4ursVwWbGBD6c42/dZc4Thh4wNoaV7dTSo895qtxrZMfHgFX6jJKWId+uWwtgBnOR7XAkF
atGrZiI/HJmsrC0D4OODHYaiNka4KktfOb0A82JmkcsYSdV+pI8yX569rhWUbTZtCeFh3ThajBzB
KFb65MHmDZcwr4+dxHLtJbo+L6kpQRatUkTzgfy779pB340Mw7dDju2245Q+Cba0pTO+2KDIU5X2
tenmmecCWy2KV/hJMJND5R2CkkPiDz4XQActhxboFG2J1I7W2GsnysJpRm3jNRMFwKvkDzNtrUj6
nARCKCl9+AncKi6/aLrpLt545uNrskdLAFnLiicOLWixQT9/dBsZeB/zT5P0bL50H9qKNAU5lli8
TQpQUUpsGQ0SEurioadvTd3lH6aIShYWwoukDWTLRQqqkjB2thbFE001+72nQwF+rJ2y7+gUEPjw
Jr4n3fwrusIXEYJzBqQhuJVmQOpBRboNsYKqkIl15kQL+2Wm2n7TO87pVFC/L2wCT7Pf2E9EqK/E
oBHmByNhFtjzjxUNGO++5ou4H0Ix7cQcyN7mD0+lFh4s/OMVJ6gcSBJF6Gvqh5wX7fzmVjvfnPpJ
ifNemRGDZpbD3fCb6gLtjeDzHq5qSF+FLeGePO3v9mgbKNJCxtcDS9pdhJUNWTZHLRqChNmZ1SrU
s8i6FOekFkPUUFSnGy3OPE2LLjDaOorf9QXbiq1p2PlaHxOLAHz5EaOnVCr37s6vIkt/lIqy9MKz
4tp05HMCuD9E0QOxxXfg+T+KqCUb8bytqKc2NsZJIi+MVtsFwnV0CL0cUahaaqcXzWToZtmy1vcu
VegrnVGiLP9JB5oc3a6+CaB3X0ObShJJt8HhVcFl6MOAkJt/uHoxLsp2qPzYMGg+MmdBKQP9qG0E
2vmY6bcOvUTp/BY/wXS1rjDtnDZTFVhahBFZoYs6wNwFII6+RaeGkhE87bnH/opTxGQrVFZ/+GUw
pjmDUtmwEoLN7HLvxONiSAxShXGMiSFxJ48iEktW/VCtBj9G5EuNKlgl61qXDE0Dokn2g/oHSTQH
oEm6Ddc+o8Kxwi5FvxlrJ3isnHo/bWiWBlEpFR+icjZ9DQqmjA3t4sj1mVk4028qiICIQuT7c8ZZ
EWG2g0BTO8EQ6QAXcpiAnUgc5I2IdFJm+AXEq1nIiTYmFCQAgcv+moBXiB5gJRFfVXK9BDNsjsqH
QZnmoVmsdVaEuvMT/572b/FwSN6NbGORq1V718hTFVq+KETQIPK0F/HFrVVgALg7i+e437uw43Ho
HCRMT3VVS/gQKlFTdxHNYirDJZKxAww1rCfP7ATgtj3QIo1dlx+13oR7LVkD2juBFCa32FTBYWI2
zqW330w3JJaEmLKXls2wbUTSuXkScmNOtZHunt3nj2lO15SjSrN5yVyw+f2Rj4GAcpInoTzJpRWX
cCEwhG7wMvzdLkREe4pt9e2+RNwOJbkdROM2vWb0hLV/zaQHNKfBW+IGlu3VRzlxC0O2fSEAI+4J
6Di3IBh2ImZh+W7XaU1swdvutdq5lKGFUmzYy6YQoU+aQeBjvMqgrGNV1z9jj86+Al+JldhpfYvw
ARPsd9q2QC6pSrB3TgKPxbGcrrrR+jpySFwEdrHPYv7WrW6yStaAWliL0up71g+/pM4wzYnuZnES
Li/pZBzlwuQVL5EszCt0wa9MmSLnlscVDDJfV0REKzaF7lW3A/yQEOQlKf/vdPyUq8bAFO+IGkA5
sJGw+8VKDUhaccf44/OrAIKI1T/Sm0oeB7HMt7bAeVV1CNeRGrEsMeoocaQSt/7tMMCRi+FzX6RE
bhzViAbusagJty9IMPtKqn8RMAHCDKB0WQzrcWjXSXGY/qV6oOgvz86K3jdKBBAsuW2qOzbEI4iQ
1aoNyPfoWABWVg+lnGrmoYLgccAV2+NUgiZX8v1Qo+9/k7Htq6tfyTRHel4pPWPO5mBOHNuCXjLq
Slpvr84/ZS5LDGhmBC2FHIvE8D3DcbLWqUeXAcbeTiC84NXdw/Q/Y/iEMM3p2dlPxp0KfotUZDeb
GUaFBK889N9PZlzVyExxq6j15NhX0CgjLaJV8UtChl/VgGVE5/pAl6/V1WGeNMWA2uzKcimeDjp7
G+8+E9JBrM5k6ckUdNA4Kf1iU3mKJZWFqUczGMev0Lf2r+jsGQy3D3DKRAiR6PBsCWs0cZVBboV8
YLr69OGt5nAa9U1tegr5VAFYveEZoHDE1zuD5OxV61/QS0ia1q5UWc7OV2y07eQHKUWa8CfjI2QT
q7rKGNaDkdGNmeDbscpPsMaQTr1oqlC4sTwzXor9AVAlt7zf2WUdt8m2JFjtYFAAXrimI9p85juA
JQeP+uSr2/KjQzx7U9KoZkXYSeop5zbIwESu0aVvU+IOE3XW3PBd0WPV+vScTgCC0dpRgRhgnfaQ
AgBBCcLdApUhErJrzAMA1jPxXy4X67Iynarwdkh8vhZoFqJrHZ9c9hQi55D7UVVv0Oaay/UEZ66+
KHmB5SuXFx7DPuQAAMFAG5jt1FY+LCI4/jUhcxll56GCbZYCCqLv9WuP9nOogzG7sRs90dJHBZ+L
1ulrMsMxGQS3suyQnNeida+OJaDSU9uJ+ZBAqa2kzwngGTC0agNvEp0oTqcAxaXLaMGEvrJgHFA+
GtjWpjTsZvDZLQhwVPABw5E3Li8Jv3VczF3LsDFYFelu50RD26vKdQJBTCsole7shQEVFXfn4P17
E/OjIcjMv6s3cgcTV8zs87WLkGMf3PvlxULyloujrQQKux6BHqcGMCYO3bQtJ3EsEqVceltWwplh
SsnOqDfZFLR7120j3sEr18PhYXKSFRvDGV9KzUjYZssRGd1QVb/5Ong989fjkz9637NJdSm5BYQ8
j2ILi6akN6MWsPfouW+w1ELkSqcTIT5aqARhIkUkZwQ7yhnDaR8NAjF18buim99w4/45aRSLEUao
8OqCt3truPEv7ishDD9krD0gPDn9YENaMQ4zV7X/7YOwAlNyRa70Q4uJjUlvhAWE9wfcp5QZ820z
WE7QXr/3okF74Zp23KBOgTD2mOvqRcHagQjn6lLA3fGCE/wFSQzDNmaNRJMT5iVfbJBEqMsQ+wFq
08gMQKhjrV6feSVtz/sYeRoNPTCKCqVre25gsjEQNnR1Dnt7TqLPXKBnx/WpBElRJC70AsDwHq30
ZwCG+n+oIzDMMEK7k0J0WAmYqM+1DtEKN9RuT3dWFENxBt1SHoEEztcr7Sb21zCjxpHzSiRS4Fii
fInkXeA5WiL3pTkvgyLE/L44k5RtDyG4x5ygYGYXJzPgq00Zk3kk3HFTpgGCiJZMX67EtFvu9Rkq
Odz6lGlvsL505r3LZNBmgjma10JFc+IsBkcBRrLSJCkxi35hdsLuaOO7eolTLd1t/1DzZ2yXuJoo
UnnpPlezMphoOWRLP5YUXqu5JKgdjnyRdu/FwwVnbTHTae+KranhLdivKy7NtRAOub7Gi4xMLV61
iURwwAPowH+Y7kgUe2gi2Z9DGvXPs85Ld/HzS0ULcuqtXGPkf4G9vUymWtPs17NroqDlxuKnfHBB
QHfHdwzIKorFoWcPyZPA6vIgy1UEgOWQztyNH2FHrbPqJYAnbqkWelVDUcyZzsbtAI3DPosyv9PG
Q/LWyUmNe4CFgVYBZ1rItLfvqH9b6wfstrao9ZTKJRxuwj6CskpeJWrbVqfgfnorDfPiPJADZyHU
7GoWjei/K4wL9xTw2/jAjPWujNmyzeVwNVVnQTaWecUxNVtQDNIjE9JuKLCQJ4e5lKdVfnsyXm7E
TN7y3PX/9RgSKVmhmXgQrE9yOibOI0Ss2/fIo5Ez5OdRm5DpRo+Ww4KfqNQxUPPXM0vFKrj6uV6w
SGTtFG5tf3YzIXjB9KKBQDHOhAHEoKLwjc4LJ0Crfqn3k5QFAmeDIZklm6vOlg9qmEuhDYekaKNv
osauaYPcYcbVa51g/8NggRz0gy8pdLfvzPX926OXLjoLndF+4lSPHhiV2EkeQKXXnDH7BaXd0QiR
FnVKAoI1R0dW7DJLoW0p59Ah2t0lwjWXHC8a+zSzvqvvakC2vFX1cKZ/U5OMzVPuFRkOPaGNBrT1
V/1gNzHhw0JMUlSLL+gbS8/jk77aWlKkhIIcJmd9xEd7OT0PsF9knxrMQUimqe73JyWL+aeD6k9o
sgS6AVRFf1BgMTPrGQmHu/4mlIrBmXdCDcM4I8IYwwmikIzJx9M4c8kNB0TDIoqOdsrjydtiqDSl
IdOUNM8LZ90743pb6D5BhQNRpmoAby6wZ2pbZ++Ot9MeR7bqZBwwVsn7l73G5gjDKjrQMLZBa2tm
RFst7T1JXKyBu0/XJiVdavontcOls3Y3/a0Gi+pf4R0MN04qnqM48BXJkhDvGcRD7TSccp1f3rNg
ow0BVNS9OcXURm5YYJPtNb95Wa5clTG9TrrGTYEiV8ua5rAk0jZ/xHf7LtmRkzA9jw9umr6gZVGC
rWXXB9UxvnGVJxqbz1Itx1ayZcabJIieW55+fotLnyc4gjFhAL8WmHdceeL7kesKsnALRF+ZCq9I
G8sWcKJFoJiDGtpMs7OimWLrOPSLlJFqb/GOHIaR45KZto5WfYdxBORYzUV1Y3L29vHojTTpqtjU
HSkL7cLX/M8rxpvwXl9wFFOSR/KT438Mibgi+FwQFzpKm2Kx76IFTaotB5yNyl6DJ4KC2gitynmv
ucoSQO/MjSalEHypZg8OcckQGyCi7v/kuEYjAy+4fSGORkLJsi4vvsJR9ahN5U6A3REVJhKv19zQ
MWBtCzMKYRuRh8abFvh2MjX1RooyFo4zmFeWdmaSJFEuLjflAqQQ0vtmRQYYiq5t2ME6d4BZnneo
AvFpQt2sVkhurKoXmL0t/WUJLVeYamC5G/5h1OqWNehQwboTZWHoV8m2KeKVaotfJiihCHSgjWMB
51GbLCAuepHty8xzWBHMLza/7VRfrdcThW20iYbtwe77YQevjakfC5uidHEi5InOUriGky9LnDHW
R1OHfjIc3J8nWxxFpdbvRrmYWmf9QkorPdDa5cdq8iRlZ86PwWYzE1gqInAJwCGwt5X8M6970LLY
76xqGhEZhZoJnPaRLoB2OzOaUAom70Hp+u0eRSC/vZKzr74G0yeqCpM1kTBA2N3Ce/IM17uEnlYt
15hD1TS0ynmo7TyTQdW9hTjOICMQC7mrh4kkZFcbyWZEe6eE9fNGz+YVPMStc5qYdKGnm50y8q1X
C55Ykqw/PUjFgpfMCA4jzpuCxwGHjGS11bNr5AjRKDCVrZT6HEivNM5/uwRJiexYxTzqxEv5g+RK
H6r+Z7s+23JxjupsqzLLOyCtTLcB+o5PUtJJSNGmh6Htz+LPMg6taBPqxxdDmGq8j2LebHC0QlOG
mN41qEXEK22HeHFD1ulU3wZMlj7ldYfInDAETvMahvKzgHtws7K5qBY9E+WI6tJI9xv6diZY8VuR
TtxBRjSGyjmUR4eai10I50090JMfokimtdV93qHsdhGVDfLgfJPAP++YFAveRfWixy+iC3ykJ5tx
h0Vob7AS0melTASyiLohUv+Z75cICl6kuyLagOGffnx1Sc7YHDGq8wJAs4h7tI5Y7wm4cjMqMZsD
hBuMcJ58Cyw8ZFHBsx2EPn1emOjF8SyLi34L+L7LwX4qDL+1S8tShAa3IG7tA0B1N24Ybx6EXwL4
xf6ssQijBWtBsDnRp+OUQeX1IeN22gaJg4DN28gXKKiJ8O5VuZ3lPbRcL48OxlIEwCdX5OrX5ByS
XirPToz3Q6/2iKZ+yfRU3hrwp+6+3W+1IIboBwhOc/QrELNo/ru1xiyQ2KvLHEr06fHYprq3nHVl
vBZGRiqfSKMFt3MH0ifu2QnVzKvYgYFdBPB9ZqpQ0WeQj23FubD26G0qtKAlPcjU2duXPRlh8/zG
nY08mA/b3jgr0VI02z3F9UBZgCkUnuQRrGiq5dFXa39Jwc1jjCoUFm76692ZdmVseleKwjLRC4jz
2+PS/Wz5yPKYl3qK02t/SfNIa72p4ZWJvDkChsebJx8VO6w30EUY4MmiBEW6Rmp5Zmev5gqE3Fs3
Z43kBehQsu1fuKs3O5qhrRUjaykCyflNg0khrltZ1fhhPYv+LuqTMdejMP3w4d0XYISC3keq636R
LXFJFLtx1SsAa0kn2GOX3zlvBTRfwyR3fIGqDsHI3srXvzcNLRjbHjUh/+pgjMkPNxOb7bVeSkOy
Vb27TlbOcAZU8YXEgn4/r/txk3J+L1RY1gOS/FdGZGFl0LypYMRrqJIE8Rs/lanRZDwhJssSCyN6
BoTLhdi36YZNXReFZsdddUKssNzMyF38MVPl60j1NfBoXeIH2hrEjOvpHA9NCF0bYCGufI00jx2f
bqTLQ1qzP9mktgscEmkQR2tR2U1nx0HArplHt5hWIpoP3vlql6hdiMZYyiHaTHlm4aZPnxrKCITi
DkrTyz8oSbo1v1RpmEViUXWRbZFYgnGs/fIsEH14KPY2pLdXhG+CtRc5rSQAXKvWbvEuo+thy7c9
nNozjgbsvIqz96WANvGFHlEG4t+oyGen3fWt8T6x1Fao/wxxRPErYiEMtn6XurXUoPAgrlNVnTo8
aGpmesH0OMht0U6lVJ7hcAMhfMd//LOt7eMamv7BpCbQ1edjPxE+rMyI3nznYZs98LJ1F3Xp5XPs
vScXehFDusEXEPe32tYFGFlZl5A8xmLvx5FQtW5ti0zyaxbLNa7GAY+GfKXsDOeo1J4oDCZMr868
Q0oynOPuxUkrD+RXzQDJpC/8nz2ehE8zgg5JPggOoftdq9OGQfgjVr2YRWF15aHdrj3UO+UWKC/3
HFcxRVEAPkvIg3v8wwKLRzDZR301qJshOM4weryuK8EULALS+BrjDk+HsMsXJ51geFlk/xj+72SG
M0C6fwkDj7Sm1do3oNBRBfcBcJjC4xtLM1lRguJZhlBnnVRvi2hOLxGYcGzCWL2sBJql5EAjVYgq
z7llUH5ivnlvipQFVc6kyJw0h3pxWGxpvGeH35TUhXAtRcS1gjWXZN5wkU4W2hnPwPC0gtrvV2+s
R3YC5rE2f1k4hjmy2cuqbSpjrsD+E0N4cX3LZTp0+JknDiGy5UftFHhr3fU1+OYeGEnMTEjPgceB
3PYIjJgAgmHgbgMSUgL6hH+6AmCUUcEsUUtNWuku8ube3IEoac1v2CaVK5ojeGrpZSDg83VOnv89
si+Bjj0lxIQ+A50tpvzj1Leb2fX7567iU55VmYWgZSh9rjwkNoZ6oQFdGXpWxbLBs2GujCisMMlQ
WL1gNe2VX0IeWcFuL894pwwBS4P/tcUzDKLnrEjlUrhrz0JPcpTPlRrkXWeEFKHuVRw2YMM8I68e
+SB/4jlUAGhKvnLO4u/cS1sbsVarHNLL76awn6kgfQck+fIBLgGpYwQ1NjWBpDEnflWGFV9jKjC/
0FCA8HOwYS5TAJUDvkM8HOMsVG30lze7uti99EYk3B1q8zqdsiQ3/7pcYBS5oclvQOfbzO0lUkjD
K96PYfIp2qlSL806nEcy4k3KeyCBpSeVxEJmgZJFnGkAE9KvS1Idh5qIU1R2xVt8GB1fmwIrLBkT
qpHAPvXn1aP7sxGObhyYKVMeIKGA7QMkOyqwda1QcHYqhztIU0QBNLEDG/Bj0rPnS+Oi/HaszDkB
oEr91w6wJXCHSx9jhYq2CM+eJ9EgnanSsLMOgCP+3mIm2pKqV4Lo3E8hQYFHI3MKWO3fuYOUeYdE
oSh0NVAipIp7YYPpKrY5Fe6qOfeDCjD4rajWFV4JH+BL8JqUAK/zGnCUbHUVD9ksbmxTPThuCNOt
Er4A+3U+VP2N1SzTRm476Lok4tv1SwITPYfrPUSQ1ceIiViUmV6JCbdGNpCkKgWp6LsytgANudqu
biLyjaY3zRubeR7bRXX3q4NalACpVmwestfIPVr3ZYP1OC4yY8i3TDfGhzD0Cu+Xpnb+d07e+yRr
k7aEpzXemb/qksxKwFjUfWGF+Pyg7jJ898X+JczN7f6ouCSQwLkZInoKBbih3SGiyNG6zwTc20O9
of8VZqwyrvVxG7Kx5Z5HqHDgbG0omgCOBHITixnBI4a5OBUStvpjX9T4gqAdNNYT5xrHVFYJzKEU
jjt5+1Hu3ythowimYpvjoPWW1O+39eErcagL48GxZvY1RLOq+dcvLdVVwk91HyZTAuvUxkgBNQwx
MSx1u5T9iBmTqCX6Ma2Fho7Sl2eWB45MHBWqtWlZabLvwqR92sypdA4OU7+dipB2isZIVNQldjzv
P4W5It+A0KumTSXhXZ3kMYV/6GSirKcXyuv57jYCeFR6gG3H4MIyR6Xr1Ke7XHYdzXB3SVbluYiL
RCxIJ+HOmzk3kwYYTXBLgVTaMsDorQw0K0LexcnhSWhQSviy42vSN29yYHOYgjxxkYbp5e9c9UIT
gMq4iC+Zy+jEpYkKnHksLIHJxKFfRfr8+9l6oCKvW2ItF07SwZRn/dtRolZmqkpM99pAF00wE105
FlAvY+M0PCm2CqB912ucnPzFl+qYSd3K0BncmJ6i9oc=
`protect end_protected
