-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mj50H369BKNiO01JvS0o/lsA7vme0n4nzQL3jTRaSMPnlVqr0FuyepIG8oyEnytopvaLga5p8GW+
B/8GR8UmXiZC/fT0+AhxKQdCvZ4OPDkCZh8Z2VoQTFEGWuK5QawsLCf8Ddm4Hh2UbFzkcHsXdL5h
mweddJpWLTy1rmjpvYqxXlKrQJCG2iCxqaNkVEFKIksio+IVhoQvqx/r9K3aMeNK/RaT+aE2Jqvc
kfsqTKGUF3gfHOO7lxIhZocbEyj5+m9w9wUjz7eePTjJiZHHiqRJ/WIO+a6Hp9lMZrC6M9JRkxNi
9O2WNYu/Leps4GRcZ5fd2VDRgis3SfCxkxek7A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6880)
`protect data_block
inVuOH1PfMzFODVdP9xQJ4sGTqOV8bGZi5UQhDuJ62ruAo6gI7qbhWRoTp8C04zcDb4cYEJG+gwF
G1h1LHmJQhKIzGOHHFKlhFqLThXjwQKuMaEka2QFLnAkB2eKMNKxGjin6s1UOOjwXIJ755rx27Qb
Ri0cimzdF1CZ8s4EOMWiUxmRsqeIptDnSgW4w7sHdyfnZn51vH2/5SV2V+e1m9GoraJlNoY2go69
s7sBJ74bezEM36+O4MxMn9Z1qXiqc/oZymChG4fTx+f6YFaO1IEU/HEA0ubWIxqy77caeARlSVPh
EXN2uUKdcJwsp3FgDx4wPTEnpILXDChGGqyDMS27HiHOLRNEwu+nVZZW0Mx6gJFhJImOX72aVAPn
Vyk9V1O2KDyJg6dhtyK8hITVL2RCc0TeUZHEgyuYiquzdpZgbrfKgynz7bYco/ssKP5saioXheMq
IvIDSzrAR8G1FW/pwUenTmAUXMWOfBXrPuuDKo/RE3yXzMw6Txf82S+B4v0P4uC8OXiemnaTJ9Bk
CW25DZpAIDgIQC3wXY4+GrgNBCxh8BPRagr3CL80knP+k4Cq4WGG6MLlskWRsIFNqQTMFBl1/VjC
i3v7AEToxZOpSwfVuVBVgopmY9smv65Q7uyP+SjI4zvdd+zDzTkCGQotVGITJDoE+Lr2I2/IRr0L
V3Y5UGlr5P+EWXGAxhHfsbn2gNurKSU5dIpWRz7wd4rzA3tXc3xFeHazbEoVnw56/HGhQIiaZU9F
ZPBImhnsDH2r2pIpSI3CElzxwtaGV2HvbXVPAwVE9xy41QG3v60RHOCQZeRilZqP0iYdKCwI1ZUa
XryJH3daH226xQg9mLWtyeE6xPUQ5zZBIspIVdgCsIIJY/nfzmcyBreriA3hf9u5v1NnqMrJUoZ6
QfHi3YjQmke5WH66oBuMxxYHLE+o0WjI/8qkDNfK+ucCeViWLL2QgpZOoH2ReDxIboD52c9UFpaX
yFQ9L/N71g77Wdb9WQSVlwmD4+co1ixso6VgNhojbEakUYBFHan4C4XDPgEhY3FJb54/K8fmUofE
BSs6IEqSNkSoVk2+zZc+5kCx2rBBaN3oeJSFCocRxV3ZJuR0fakuSu1dg/TocxAotVLLdoIJ/6Jz
j76Ik5qTN7cT8I/Q64e0X7npCSj7YwYaTjU7h1eY/kK0g4OqWqPCBKiifOqr90uJ4r4m/d4TUeJp
KrtLly41WpAaFPZtpQXIQ2QK8hUk3NnmtQjYE+Rd8DSh4GupBaGoL1wOZNjdGbcfI/g5FYYEvE5T
jDYZ2oLL+X6pkBBDWeeBU4AIgrqaWP3AvTcMwiEapSaH3+mXl69X1oBQ1ozK66EfyeVwuKICfgCD
DIHpMT5+oyZ0iiggmqg1OSHgm/pZWWOfTlS3tRHIDS6q0Ihtyc29+3cjVZOOJj7a0VmiKbK11m66
rZhhyNLdK+bpAixLG5Ma9RfnY5jBeoKZRM/cE86CGtHi7edL8rGdtXFC2/CFvJ0STNe+zXZaQhAA
P6mdoLzooEoup+S0VMIG4NeofMnIc9NXUenGpXUFfrGPnWzdaAK2zdR2u2Ld3ESorn/rER4JjU6P
dpkOhzz3TKWS6QHl17WmyPmZGD0ZAQRrBUIeZzrMsq+PBCw4TA9kXs7PEfzGKGHA0CF9UMr8vAab
sYN4XzW4Kx2ykRqIqFGAXh/8sHXBZlOQ0M3lv2wgW+hC6Sa02bqwXH/z9Mgkef8GN+SER00ufKeg
3cSd7+TaVEqabMUbkamBuWlgE9qiQPgsR/RrYW6MXRR0vvDBZT257fPgP6FLgRs53SXHlvjSxvw4
I3O1yCPj/1TuvTLtaDl8zpHXu0OGqjYxq1WYkycuH3uEtbPyWsPJ6K/Qe3+qUg3GqBWfdzWtEvQK
FSoY3LQ1w6KAxAURm3geETITduEyJHDlVr4kLuMiBrDhb2ir0BVbgM2fn/uzdsS49nB/HwVtde7x
mueNnrVmC4QKghxcmkABgWPkTb5EYdA3/krzb8uACMTOvXX3mrFeXOPqHWnSQTrgZ/rAqk67PjzM
BQT9Nr3seoSHV1QZwGi+j2QxpYlPT5enyKkjj0BJa/p0E//Pjhj1Ioa1+VqS+ADSYjsqBHG2l7WW
yTEy/ftvqKTUxhH6j35f1GulI9hQXE6QrYfs25pDFK8Ow0Dkyyu8VzGeXmvk1GASe06L942hOxMK
5b86tHt5Q6fcdq2E0m2iUwfbUH0NE4RF9gbVlwY426jeqtQaA2L5+Jprx2OW8VYAj5N5SVzgEKeC
i2evtec25I60R6LjCvLY9mUoFtgV/EX2nmMiLnU8RuQvytlK0/fZac2qDfd55CMogJgFGQP6TUjs
hFHLBg2ahBqLedIa32+v/Y4JDJJbl0qI9Apt3+QbIkwI+uCd709ny3Or1PCOd15V2slJzYSjk4eN
u4lFKYJ+d18Tu/qSXk0sKxn/nYW3O28IDwsKTLGW15Rj/7HvEqv2JlpPRBg0yVmpN3iyAAkz1xI7
C2r5VPJRAEH8H0YmM4joRgzDQqMC6lUOsoTgONZH43ev2m9a/urG8qGQkAtgoEM3EIZ/+2hrU7AY
fIpa/lXklmdkoRLAGlOt6/b9/jyHUeD2jJkz0SQxSa3WJRMcJNxd3h4T7/Nt8Zwv0rr474qmFkZL
F4WHkpfm+ZZSCKwTYdFIqF3eWBGmmNVKUkPkfwtXWy2iBfQ8zbF+txInLdEwGudF94LWJni3TjMY
kHuJeyPqv7tlE3jOSEUXFKuH6SytQUNDFbNW6+BnJ1HPiPcX9pNHP71I2DCJ1aJV+Kfw9yxZ2AII
E9M8XV3ULGm+mPu3UO0EYidf9wPfQM1HlvypKJCa5D6LjmLdjcS+zcK5GRTgFNrnnFLLQogd1xNB
/AIXi4mctFZRLsf7YJvhHApvs/2ljxloAcka1JewOTg5Ua69d7afJjTMjQ0iGJDfRJXS21mCPDyt
esgmbg69X+bHhlU5M4TGP8YaUJ9P9SDpHTur124FPFCulSW/X/iNMNPOpV4UoWFu3NI7eeDjjy/M
PsDbcZOAZKCWmZDXUtIE6r0vXBFEbyYJfptBFbelnLWGOUzjFMM0s2N2LtiVBkj8S+1cNnHJwjNQ
HB+PScL+FLn4Gl2vM7rKx12ax/+crZYpnkwPCPM8+QQtCwpGu2OG2IXd5+2fIWVSS4kJIM+UQ2Em
vvIxxWrVTrKtt4e3zGjPCOg/8UCD+3MLCTVdWAUMJ1XcFcY804CQX4siIeIaiLs0OkPzwvTmLHqj
5fGbh7p4yijfAI5pP3CRlQsfq0kbm6hYe0++5kyUvU572mWpQBq/rYe8uvIZZXGRQ1AKTWC8xfLw
aJ38Jis7dBHJIJVx0uSOQRAPf+4dux2ZuGYvkgTkyYbuatyYwFlYNSs1y8C8GhFh34WoCCsRmy8m
KSf7PUHoHcNER0xD3EFlseI8nNn/eXmXBzhrCAyRyZTDoRJQV2XnQ1u9gDkNGi1DyMbXjAxe1WlM
8N7DxsTnyapRgIhE8sCAelSbnDk1bEMBs/fw5KoUGGJhDfC1hAaGvuIq79aloaJAhIf4T0Ci44+a
YCi2+/w4nobCGnczuCa/GUnh/L06qR2h7jQ9n5Sy6sRfALNJxgmx+zAT0Ol93vobyyMqYgLdQL8+
jpXI46NTi/BQ8FJQ31qEsawR2TloOoULliLkuRcYszO8Tp/JKCDzS/RsypM2ivvrY/rtALs+OmFl
5IPvKHMzTWS18tDJS4MZp9ZUN8UNLHfqWuFDyVj8cdSdp5lKUHCDxv5iMqtZw05NMMPjD+DeIv+g
OYvOG7KNlgbesoPmVWFM1s0hE80jma+05K2r+40w9O+clMkuabU1YDnJAcug7cKPv5Z10qX/0RkY
V1TfM9jB/QgXQM8nTDonJeQ9kChtTC9eaX/AtJ7uzDmUcw8SR/+gPrOYAB0zibU1tFvyO24+rjEp
QNAOyYT9gPGpcAavgUhYvXCJs3fui6b3BsQJDeTAXK3yvevgWjZ6CyhTlXNfsko8jrTx3zSTYdIk
bp7aH2Mn/ZH4W8x4bR7+md7y4k6qdFsKnJeAMAuy09MTJIWTTcN6Gf11rsPhjRkZDYxkDQdppi2L
L1VLOUM+zOQCw01qmEh2tMD3MoUazjOOFTSeXQN/zcRDJbe8AisxftZtwNTUEyeBZX6oBtkPmfqX
xcIt81YH1GmUVSPDbm7Q406F6uYfD/W5H1SAnVpY3LoJhBM8lR6APNG17IU7Po++PdWUmEE5nJP0
5OG7psnaqNj+3BfuVTcvFEBetHyEst+VLAH+300vVr/Dck1ybJBR+8YVrCRZRm5171Q4DaK2roXj
YpkPaPbRW0R/x89rJ16ib/dOgq9KIcSh+9q6AwK6acfbZ0vwpbb7y1MdLlmBnCBZzh8p1BZ6sZzB
7xSAVvO2m4vTXEP2ICLDlIugpHxHHPwGiXjviP4NFmHRe3Pt34QPv0nAkfc8udnmIS/V8Ai94y+x
0jxqkRABm+CmBLCBKPn0/VkAfXqqeeSHS2ypbd+g3cYDC3PVC8QMtlIF23DgPn2O2WIckmImiTK1
4a4wIl23nGsWS1wpF0e8tJuL4Mk4P8qGUqcTDXcTBea51JUNtWfW1vihwnDA+dgBmbMTvLl6oRaZ
yu9nq5FscI3tqx1wJEphs797boGTumYBkdYjwIMs5COhSDzJPBID56Fw3qtjDS1io0qureierPoS
rpKW9zmZfp4Bsmt1K+jFmXo7B2gp7Dfrx1teLg/vTu9aoytxO+6orGKx7vu4yxFLQTz1pJiR8klR
zz+lz4sCELMrSa7C2stGhmMj0OnY7PdqMlsY0VKzjFHXb5nSUCW9AixYWcyZFtBXRGLDHXe/BHBb
kcYILRZwpRvnLCXUhsiLRBuh6tTbJPzmrAZ8tE4djgCBAt0M5TIP4nzwrslOPxyY6ufBT1b1icuM
rihRA8fics9cmb7zGDjNJj6/n1nP676JQnp7s8OeaS6yzxJblLEf96edYtaDOEpZnu7QUGw6nevC
2TM0DFo0OnqrLu5K6r4fWtBh6kDDW3BUL7OA/HL+LZTzndpA4EYURyQoVJdPY+mDT5mQlYgzKhdL
kHXbP/+lJ3kT3z7IiKlNIVzEesxImFG+iqrN/gtSdyQvHYAZ2EBU0Uo8u+5S1oHtrYaEN74/ORdb
prd5bMtOJuVg5IyCd4bX2YX4VlzEasyE2Zi2wCceQVGKhQnCy0Gv884g859GG/41LDFiK7l+uBEt
Aiovi40pDBzCjipTMkes5spDK1GTowsJ+Hca/MI6zGpiTRh/A6+LUWr1lz417edIQNBCCDtXSEXx
LtVxGKMnLofxBIUSnxPqsnYZOZpSvoIu4YF8pSaUNLZQIzrOCRYrxcBpshhiz/hkCQN0eX9BlTfe
x0o9u7lSNtaUw0iPVUUVVeaN/tcdiEEEjCbOl7yUMWvmrbnWmcICrimpGGoA0MLIDcBT0HcMewLQ
nI3cx3XJ1FYVoohmm/6XdX9kVIJlXZo7WO29yGkIgLe06+3roRYm1jtL59jimBHrXTUUfHUqWkXp
ra0Ed4XllJqxoNJcnKI7nHiC8NoOEw+tIWCwqgYT/RR8NqlAmotFMfTBOlGkTCY1lHjLzeR1cf4j
r+O/fycspp8lKMojFM0bUSSwwds7FAQYDktFxKU6coDT1gzJVUg6bTHWQDQLnS5burwgoOAy+plm
Z1rZPmEKM4eHchvoi5EylPv82/jShT5LSrkHJc+kfeX3SH7xuCSo3z3iEx2HNsELDBAKXIdUy647
UQsoivCpUaJcZiTO5A5miorqtbkFhvSZ+XVZh4POJ7b9qiItUkCQp4wTTnl7XG3MkaYLMGyKhfFM
uknhvDwTRMJ/j1UgxbJg0HcgqgEquP7oDr7GUVLLtXeHf0lvmDKV0rfT5aOj+sZLMP9kqhfZuJnc
KcXKQ72MklLys1AwrB7yTWULroy/jFClenLhCfB+HC3KizUJVoulrsaSKYQDZyTp60via97D9CFQ
UfEZbmBHNSbbIZRhRpuXOW4C32x+TP9zm/qgy6hlV2ZUva2Y3Bjt6E8thWX+ZnPVtpjmsIs9CnIR
o0nrriZAOLNZsGlks43Q9n64lT+kYX/nF8DCZXM+VF3lADvM8h9z7i1pVb3ARE8G259j07aBW7xC
a188mhB5wT2XUvZVgaHGVwywF7EqDWqQomxBaV19wCghfxnAazcsG3PSbE80o7GqHV4NC/lngPzP
nEeDbJwS/A7S6uPBr7hJQgsbVdI8/zoTgGcwuo1qCvt2s5L67aKec3OMP+xoLYlx6+QY1XT42mHn
iwwntEejXyt3kFlFE2R0QdT3cqSgTpNKjNWWb1K4ZNQW0HPIxNsBq0tokVbPmEF9Fk9jpZXyrh50
X2HWKTOeS77m2VE7e7nFE54jDPNOI8x8+Aja3XlLfQm1T+1mHpnHwPH8b9l+9KV+UWppTWhFziZn
JbaxV3zxJE1Oi1JNQDVSRSHJjuHS7NRjV6NGccYZnV6vcT8zu4w1xDmZvTGdxOusIMpLBLNiia8i
0rCWoEW+IRiP1lPjzo3iSzyIeC1tH8oFF6Ok0eYDbPV9Kdi/XXGRxEJzJpotYMj14be2gUQN0vIp
1dychRHZlUJN+hZK/ncwAKetDij8LszaqLcnw61MdU0VPUrTwSw9PUn+1KQPNzHeVhfa6SiRXL/W
cJNu+izNy2sNxQ7S2odVa7U8eECGsaUkMJuKbHuhzJDk/cfVdDS15WCbIoBZNRQOn1w6waCQqieR
MMJj1nxEQ5dQlE7NvPRC7jjc73xrQk221Iqbr17kQYP8Z9q5Rr8j5J/dkn2Whvu/BZub4EtrIl2J
Dmnmv+hYJtS8rOQnDcYTEDT69YiUXjv6IRJirSNT1NRLs82PUzKGdri7DDklZHOFndr4XrCrmu/y
g3faQSdqIsH72TkWk0N7QQPN+za7eJEzDy5Qi2PBSDQs310m+DPTgwnf4iW3svyZSA2CSNXuOaV4
0zN3FGiDeYQtuEm30RfE2W1Z18Ln704NMRvHkeOd8cySzOn2f/qyogPeM23/3V9auB34oYE3bP8r
HanGJ7Me/NhQLfEm1dwQmBi3oQxoNzsVg5hn077/0wIFv7Yh3GsaRAIy2rTPhh0U76DYTkDCSV9y
Mhd82CJlv6arS+eMm8YjrOcE9ABaxyfOHLFt9sGzKBaVEwCcyKtID3pHEIbZkWKkZMwM4A4PD8GD
9L/3X4017k97ymiirO9m81LSqAXJ98imJTTd3WQqG9f89FfkVqzN0t40R4kaSzd+roX5qHxw+hdz
S94iRM6j+Q9Q2uJG3JwJoXw/wHDShc6qQCuwY9n10xQisg9Xyb/aj/y6B43RpRnOpjazFpxOQ4CA
dnKc4MJOQzEwAs/CvF9OYsQS/ThDgwQKNiUaLv9RdWTHpoG+WJBBS9GZVeM8FDiWcIkoaQ/Df4CN
uVJSaebdduWuMQYQftEkdh9UNAVqKZKWzB/DZ7Ekod5ARfLxeK4Qw0onL1aMz116mOnVGZqyI7pb
uU8ggGu7bL7TaL+gYefEaK27B+CLAWTWafEqCE3OCiNifxovNxlQpQwcwls0wKmstFwGcZGye8S7
3RtQL6Jdtfz2/CCG9/E07qAgVviDFh2PrfFFdkE/fAzWkGcnzdWNZNlTZmbHf+cvw+ttAuQM9AL+
UbnI3vFQZMAVXAs3PqtAXbGnMy083Dzn8EvPZqVtTFU4sprYhf6i4dfx/YEfoOHmr8JHTpCt+JQE
wlh9Qx5gxd9f/rbTDM09Mzu3mYZJMLSKGHC2/SHCYbm0l50s9luYJtzSaoCPzITPBz3MqMp90Dj6
SNb/AId1Jtm/aIwvRk62vbgCAvzBDpqTK8YFWobA/Y0uomVkwoZBoThcwUsZNtpiu2bHhW6uw8AI
U6KpsmlSF2mPKoe8ixeRuzMZylJkbfaDvWMpQfN5oIfeCnJAPOFZgrPb0ALpVfF6tYMUIgLXixPt
EjXbGQHy7ATn9E537y7NRfPNKWqnwqLn51hy5XD7cl60TE2CBIysOzQ4C5d8uhiH5D3InoHwCiAK
j1+QoB3UbmI+G8IUHLSdZ99FwESS5ifLNUh0pL66dxePl2lwhEGxoiV1GE0l7qFACAaf724CgOI7
mGlV/vuQo70Hr7jM5jA8dN4WpiL+MJATj8GD1o7lcOWHXYBY9sE4A+4eTEDaEyQ6cMDNRY/4uD37
mx426LL/nlTdgzGKZk+G0qAsVEdXJhhkOZlOtJJw+9hzrDPVKLoWY+C6StNJXBLUKfyCPDpyE14t
UtzhAQpQC/7PJYGzovpDX3A/N/W+NessBVYayMW3FXw2xqYQRrQXFBx4zviu8U0mBxTHhX2lyXbx
/pPpF9bBMPpQqze0Ehnk9SGbUWcOA7Tz3GhZSz0Z0DtBts6gpKH2dMqsuyk+tqfJHKq8wqbqIGqF
rTv8cLX560qWxaBHMKB1d8xUxZFUECZsQ1VUFSGH9XcMkzCbYpRgYl62AZqycK/+PB5zJGGt2YfC
qV4NStagyS7dvHdiMk/a/VVHVPlrn0PBEpYq1Ael3Eg9DJfunavhVB/o/vHbTpmUpGuDr+IpEK0B
tyC+S6ZNk6nFkgDadpWot3XHcx6VfF/50rN7uDsKgzfbF6598gVIC/AVe61GmfPJAUyTWkZeYJ5k
9aRjMIWIuPIoouB+gou90R29c/6q+M7frxUrFlkqk9he5yFV7jf656l3ryQHNRmKK2FvRCSq5rK2
FaWvr6l/mQsll8+TL2dLKKt7mTP7Rm/joID/xiOjdyHLWi3aPVdU0rub7y3DqqVe8kDa19QiZE/1
AbFappCzGRUXeQTE7m6ZfOHPdLXw4StvUnSFjQaPvS8iIWQ+U4NfRoW6Ah5jpOApx3rID7GdMs8Q
BT693eyyIPPlOFJdLxNxU59wK6o0eZwet8mrR/9aG5m+sfc/FlbgYuwg/rTKWlFltxkgbeiwJ9Vw
gPugjVvODEdtbkuOP5vAqgIVO+vPxCornqMDJDHxHRIimGOOKKtrALH2JYSjJ82zfJHavyrXFIoQ
jFmQKxeY1+SoUMmJ4kClFYAI1p8q/XH+9eseCa9nxA1Bi2Xd2Kh8EZnfRt31M8we6EUGahgGqG89
3q36xvUnosNjg5NOhxjUgvBq0cBzA2U+E1545nnkgVUxYAdfUkOmFA==
`protect end_protected
