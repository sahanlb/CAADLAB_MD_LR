-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QssYmAs4YGNlH8OWPNTiZ5EvKgp9/BUEy8PQVI+eEivdZfFDDYDAcPOCUubsk/Wv
n5KWIq4OaPgK3hmEPsmsYf+5gKJ66vJUdPvftWVaVYWZrTF4wIklnjsCVDyVyiTf
DZBQF38DeJW4tlx/oBUFIbNHFzk0BwquPZkvOvh0M8c=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6858)

`protect DATA_BLOCK
rAe4eoFHVL3T632oa+Do7PxZZO/Pqyjh/TNWs/1RPEF98O6COQHbfp+gc0t02AGt
D8Rqdu3qbMd0S3A+GEzSl0X5+ieLqWCGhkPG3J6flYhed65lFLNiasJKIp+vuXoQ
RuE6mD0f3Gujn+ovyU55H0yZgCuE6N5JwlC7MRBLuymEbcWVNVKSTnIesk1hWAXO
Kl5X/8JbRgurjlD/zVO3oCnSEZ8pg1hlB2kudt8spzmO17YWsYHFPEBRD98gwk1p
a+ybyEVVXlooUxustwrL+Du51BkGVYFaP2lNcYiSywODoHcjB8+mi4cmltkCQiTE
1LiRpTWI2Ekuc8ItrSViXBXjyS7ZZEns66HZJfR+k+dLSqw9AScWvnyrQaXEoMh6
HDu7aRBDBjJ+gNxfqpVTqkhPK8+1OBLAC1y/DUSncmtiovCErkS0Ru9C7J9OwYnX
Al2Mr/h9Vnstmu1hvQGwe3Zsbf3qN675RMSacePOgbio72jOesy+r7sM6d7/0EjF
RvzkJTjRZ39icytH2mFKvcmsE6DGLrOvRReyw2sHpcLGCirWng8DTvDcgGeMWdIz
Vc9UkEntANkuvVtenT828hfcHmNhZwprH5/HZqTjRzN4ZfDnV+YtavtAfkL+eqms
nED78ayJU/KwKOTeqVezlcoSm6Vwpbu9sK57e4fDP+Ekdq9p/+dn0KxqrssNBme8
bVRWOXOjITzjqqgHtnvZKMYqpvJj9XGTIUbaUI+58QcXQgG7puoGP/8rB1Avv76s
r9JWFeMlD0BPFxcSz/a8IyBsg3FBT5LfKc1niKHtwUx8pipHp9zcbRk778g1G7eQ
WVaosnEOraKBjTsyG9BKmly6reA0+4ZrMq5NjWA/oboTs/L9AiQLnv02U68rETUI
cwjv03jV59sNHJWQvoeCsESnyLe440cBlcE0qErq2zk9tHyJzic24O+bJxEA5hKf
AzihYEMVJ5TOw6Y80CdJkSu1fK+NEwo7Kl2LHcZ+vx5R7uDVYLoQ5B5qMbDMretw
KWCmt4s6oRG+Apj1kmNUJbXRpdQeU0EsuDv9lqN7KXOg1nucS95IgfTRrFr2Dbzi
RPvCSuN15foM3AudLK1WCDw6eF1bzz4i4rbYLQ8XVU/fJJJOritcjftsruE5+pS4
C+8sfxoMdRG+eTWiJF/6GI+dkGqX+btiZNAckBdLm6z5wgRsDKRNGSepeOMo/35I
dEUUYUKrcCEuKVM/L49jzz9D2xdILsp4Jw9QVJ8/OvJEO7v0TQoI9q8knmMil7Xr
4CYDQrBmznhmVbcPhfJ+pVb5htCmFFH1n4QRwvcik40Wo5njTgDbhX5FITX04wL1
erCC93c0Unyop2S9YGyaRzGj+ieNZvIQ2eGV2meYGjglOSEIQ16m58bfdzmIpbdK
h3XvV5i3LNP0/1/gnnI0dtuNgmdSXeIkslxLiB36WbveYKK2EsNl08KRRPTvn8JF
d9LAROzxXRRb+G5qXAv7D3wrF5+Q8iJqI/mbpHFVME6QoQgJLIwiLowZr2qxmZYA
y/0+jSY7yaURkv7YzCH59iZF44BpVb0gdfgpawW/GXP+lVNOqP9CgGQYUipisDhR
kP2nH5PdZ9sJFGnqIp9EZt2Z1iqacK5pqCk08l/5Bbs5NfJhoPl7DFyT1zmpma4f
Rr/aHIIAqA8KJnkEy3PMHKITErU1INX0HmjOOAK3I38j9Q/pIfG2giJMLEaCzmws
TkRZvXBVU5ph6fWdLtYm12KloDV5Ypjqd5aMF7atN/xUT6AnJN1OPu8a8I4wW/54
C/8cPWiZThbT6JRoEP8YmASncI9QLZV7gyFcHna4SVOavQcRXUFkTrdcK1JIv3Xm
bI2lXNJzrXBEOx5+mxKmf98AjTXOSn3KeaGV112DesnXEa0l/QBJ8uJciwoTCNfm
wb41cuvcF7RhevOLmpBWPttrwEkah9OJpSy5CHhSSofIbSSsXAdHA7gshTMhT+K3
BuiBgcezqq75T8wPA4vZM5gFZRWz4gsiiwOHqB5pQKtdMPW4nOm6wDr3ZHZcYslT
+rWOr0E4ED0LB/zAeXryfpLy798FYuSq08oi4rD/myRjxsMpeK72GrHuc/JmZwkS
WX5Rur+NyYS0eX0+eWNlOIf//TrXek41D+xewh96SVeHF6abUvslhQZeQ5wrZAdQ
Ec91l6O5oJAj3Aah3+lZKMrTIiQRlZcd7U36enURGftC00Hi5o2Pk4N151yGxenH
VR7CzWqOZyC76f4cZZvVjhY6MGDS8rnhXGOZlpEb0eSQzlbGBS1TBwFy8KAMCehY
Ca01StBsS9vKy9cv3sQQ3yjkR5n3PPdJJCf0jyE1Nuw6qVHPVU145TWLOifTazgR
Xu0vP/SbYZ/JRB0kG4K3RSoDkGLy3Rr3LnAxaS1xH47EbrCBxKD9vfAhXgvASqTW
1bLbFEMJxBmvDNEIy7xNbSVurU0jNjui6x4kPTLM4ox5m4DQo+hi/8QHtFSRnVIe
fIbgolzHdsRk3HGLwoRAEytxHUcvhvc28NiemQNPW0BPg5xdh++vFV393H9Qcri6
K4NNAXyCs/GTWlgM1w+ragUPVTyWUNYIdkO7/5zeHpq3hsF3Aedbbin57kYPm0mU
+o51OyCnRxmJ2dqxQsN1ztun1ToMemoAdJj5Lg366TQfvQiveTwWIT32Ksh0Ta71
NdmTeNvHrkNsXi2A0pXTVg9yeawTSldawQChIz3nbf7QY313Gk/tzejKf7eBO2Pf
M+W3Kbu2jJ/xqKxxVzOK27EZ7KDsSEJwaY28tkYWo0GvMjkA8jBz9/fbXvpKheHL
O4oZXqRXK/Z99PdogXYweteo61eSk9Tw3aHbFlAQ3YZ+j2EJpQCR1PzTjxcB4R5b
4iGaDfSpjmT/XZktLhm2riLrJwl03/D4XZ46YuwcWAQe2WOC8gNrHTw6CR1OHCcW
ACf9JG6uX7tv4jJPJ4esCobkfFNJB84nLgvxYu8ubukHukkR4syfsRk4c2DF9VWz
3IkZP2EXolMJXYlagmD0daIwJEfyYGIpYXVjbYB8v4LD9C712ZJzW25JfJKVAYAI
+Bvv05hEQYwt6wOpJpgi8qg96joJWE0qmICG6Ji2AyNX7G4fkiJybu819ISz+r0+
p/e/v/JwqO72jc5PcX3k+7xxyxa4866zlbmXBuEPUPvT32UpfJ7SgeYsmzHeV4U9
j7j2r5zvFkMxW5RqR8XRetBZydbO6Bo1S282J8feqKjCc9QDgH5ClRR3jPBbSL7O
Xn3KdkmwCu9/gBsEgixtMgbzJvO+XmgEqGka2yddGarKSlRD+WpPXaPigR5Ds+yU
Q+O4kwqkXsx6r+yKjQmdKjNB+fi/G2QHTY0NWMSLUPBZ2DskRmz/amy6fQDm7I1E
HOPceesNoJrwcZ6QpD2SomE7JiTenznOe0rkC5FVtI3B2hwHhApAI141Oj1yZB29
my6wY6mEZ9WNa+AfqL9xmlZsYabnBCF4o5kEXK6JPry3pvuVrfhPZGfqaouBkfIz
QLYW+uLzWMVuEag1XY3vxzQg9tH1mmnN4ukZrn44s7X2fuoO8j1qi9fZ8IXOGT2z
uAnk/qVjaEGmAcwHEmMDTFAFOwoEWoAs24ODbFa3a/V7mtax4AXvfYKXHfrkQL4C
5VUXSzkzD0GzX32XGPELNOSKpNiMwrFHBDNUDRn4Q+OFs1QT07fU0f6mXli3HErP
nDcbJ9sk3D5q6Vgkl6QcuaASONP0JkZfNbIrGfEUmP4UvwiWFv3ljodn9jq7K2xY
x+n4P8PcbkKQz1T0H4xZGaDNYSW9jY3bVrG7aPfCGbwQlrEu6C3oSH/tCcj+OwRQ
cuJ3ge0NEI5Hj4eqQCUGoERi2ngrqhKVm3R6p5SNISjMjW6ux+TtQsJQp7e0/ZmB
sTKV76tLgMkRcAaVQaRGTKxZBSk3ng4JbomnXkCvtYQng7xoyPUAC/UTwEppkuoA
ROYnk5pr8pXFSSwcY0b59yxmiH8Cb8D72aqEFdrv48E360J4WNfAbvlo2a+4Qkbr
272fytMOvTLEHtzD0+6hw7f+4a27SG1ryZjXCl3S8gfURl4aL04Vk6yR5ktNwEFd
IkOcU4aDyp4O5S3Eh+/z8WZYp+peM83lLsAt5LW0LKPeOpnHcqQJhsi+rnUnOzrS
jcqyeypc02CTeZP0h7TCpA30rlVt7642bpQNXUfP+xpluA++uOocbq7waesrQ8E8
qf30LRi6PDW4air/6wN6y4ZzWmQp+djL3Fe0oGX/8ouG6cVRSdFwTeG5XowPCJuG
kihB0VzlWhXQViY4R/EFAaHdJqmLEXVh15P952gmEAV9qCMAUw87Rq3v3Dg8IuxS
dzkGf/6lC2oqjNUEa+2PhB6rpBQgyrl1GvbsAZrqQ+K+6eEXNn5WMtEdT+1JfDVL
c/Fs+6FaruyAtsqmR2U0L59UwM0NvJN1LuhtMeN/LX7BR6yA0ucE0Pr3CCGmUjho
dAs0O+97qi084mgTKDaT8nyqg1b+LNsenAyEllIRqrgdM09ENscEDriOhB2RotaV
bM/gcD9FKXZBJH+oXrUwicJPHpd6hM08Ml/g4SQIcPvG7bN7JyPTdw+CH2W5Ik0k
OCMCdRn5HJNcoBgSjuiJdAtq4JkO6yNAtcZiVIadDum71NoK/al4zm5S+w7A7URW
TqBCTm5GWR8rC/W98a47jSUe9+WZ9Ez0EQcQKEwTKTaJKrNPHmPIYDdXVX3wVOtV
MUs9tdlJd1ojYv9nk+kWVuBmG26CWHtP0Z8XOGF4RgX0j+kQfDfXm0wj9J3eUFYX
0EBHS46gPZqF+KtkEb3FyFSjRpkho4HQekfYXhklmoDGBIedtRSihq0jCNbywuWx
35KZqC1EjWe9fwALmD9X1Y9hZQkuEH7kxLA6rKCOA/dTXIY1xh1T2FQqjBzxQ5P6
L2dt4pGEw0a3HUyetNyjZmRdl3rcRUfWH6py48xL5tJXFhkYc8JnmUhk2gNyPKJa
E+8wi7zPDaJ0fn/9Ok4S6VoSpAgcLfJnovSejUXtHFl8f90xqVU2lBW5mX/O52TP
xWUZzloGYHUzdWwlIix3x5nbvEchJ/6KqTKZgTuDewNZ+J7o7LJp92E3dbWH1x1B
ZKmwFb+8pH/xGVGB6QOFN53XiBZ900tMbO4Fy9x7BqvwNbWl5B0Tp+1LQm+YnllJ
RsjMeie3PKGnpeeHxEgd95bXEEi03fDlWJfyEnok+p2zQ5rXF02xX4c3O3ED8zFt
R96umiHcrjz3ZYkd7eLcofYBFcd1vhqvtP7pAVgrMrvHCSxn/qjXOR3CFBdDoWOo
cKJ6zsCyh6ULyEn//ogyY8QwxcB1rljVnmi57yw+9YqzK1ZneDo9NOAKiEpw4q3L
P++m88GT8vJ2aMhcxaQHiQO/lUxkXwjWvAJ9tqYuohNwnMJoCoVSz02+KewybL6E
PEz2GWqTglfHL7NRInDHh8qcGm9umfYoWTGsDp1IoCUviqFI1pCD18Tjp3ZWNao2
uMU6s7MGpDHkKcvYwwxXF2SKeD5OmEIoLaIpmOU9kU6x13xmynoa39VeMV8NxPGH
lzzXWFgFNtCplRERh7V/HfnNvSBav8lripTrURc1DwNdDVF6b8NkR+qbQpt7L7We
FIBbJNH92dAKn/muPEYEcqdlt0TKvWhW69eMQW98Un8rWJ0IxOk5vCSaUbVbTBU3
B3zJNFSTPhmHmDt9kNklmm3qJ33rqXQkaKpUR8vVJV8wS2BjibJSFlgH00j5A6+L
sRNq2lTJU33mm2OLdMA/nPHhdYt/46JSshaM6VwmSsE/NFBjWs+eGAUzfnzwCKoC
i54DeMf4MpbVWC/W/3sarJKxCKG3iVfS4+VLfycH65QbywLCy6x8DWlhJcpdNMif
lKC4HzpmeZG9QuQVVDSYKJVgjc7Qd43oFB4+IEl1y9Q7Hib2Wfk0DN3jfsn2yGeF
TaATuibLI5Qubeaq+8VfOWmanzkKYfRuPDsymZzvaMc5KbQ2EjXVXqm6l2LxKk6i
RoLlFoNI3EvkG5OHL8yQb4BFLVScH3jV5h/INErxpB3VAP0FLienfeZQ7eRoilGj
/qeMz1dm0XRgI1rnTpgOeXs1uvpV2mIkFbyn+keb0gQolbUBEjnYeKiaaOaZitJF
+SolKObT1JVvylhlS5jqErRCY8mKQeJWbq4aYYBhdijfot1zPMYk7NTQonSQAM2J
6WaMzGff1T5Weak8tBl+oV7ntBNqDPjTJLxXQj6Wuqg5vc6UouBp9seXgTOhS8AZ
IHY88j3jekryhaFW3ZB97jPu67leBPg8zR9BNwM4ZMbklwfN6pEhDMkwnkdUo9tI
Nhx8SVjj9QftKJxCQKpNQOnK3/5aG0gMV3h1gbq2jWjaV1YyGivTcWMZrOgTUpgP
FPGhiQ6y/yn27MobHVGWC8oWT9b2LAWlrgDrRMsDHL8fqLrhMnqjGHlp7KTbbl59
e5vncBGaA2yy0emrqG7DJXc2Xv1BX6PSsNsPtOupBUv3updqfwI2enRiUy3z3/7Y
wiuGGdOR3yYyYdsy2XF++VeTtVAJzOg7m9/k5lG8wGcrCWWAFqhku3VkB/o4gLYV
KmRUPXmFFGWQJ1E5zTFSSPSHUgAQ9n+/LWInN07L/85+G+qcSFO4M0RF+FU9m1gu
twBcfk51j1YfOOPCRe2Nh4SlVi9ukzr2oOpSzCK73eczw2gjly2d0xTJeT2zTHHl
AO++Fl/VE2iY0mitIAo9KnJf1DQ4MOnuer3rCK2B8MXCyx/btJJtJDywIZido1GP
YSGJunMxOSABDVa6aLheL31JFFKGmM6zptzNMaQVTIsUAeMFKUgvRYQRikEGeujb
1gZtrYfWDnHJEdQlvMKQFmD4xmFzQzzBeXY89ixLcmdCdHPFqp6zqKyXU9Jrm9uX
EAumtGl00QrN+7u9cDxmxgRUxRQH/h/rwHPecoL9a2q8EpwSJ0jxa8aobaSYCmck
liGB0kCf9r3X5DIgqENvyEekyonOTgSOU7/KrvX7FHSJ4XLOCHgumB85t2WZOG6X
BhfTyzL2YG+BPUBz1qNDMQ5WMdLBRANAPrOQHwC2/r/Bm4iMaZ/X46TOKPE7ELQu
cx7bpf4b1SgxT4z/uNAV1Qr5jTEh+98EF0GcIQK1844LJz4HkPLqjaOKlk+Qvatz
FI0e3sWJvo0V6E+wOXMVuoVrkJjrXZll4BKlfMmXs6WR9vp65QmC2hgUmPZhzO/Q
4xDAOynl4vnZqO1bY/AXZtCXZnDoz2jSx0j+sfl1b7kDPU6393qBrnfNKp07dI//
iARTgJBI04htybspg+rgAp5TaC7bs6juS7uZRUJkPBWZFgaU4TVj9q6TUqFr/yJk
PRAMbANBkrlb6KR1Dzf4nvSlLDR7MOU/3kOsj4fqWBsNftJvHMr1rnEJBTF++B1B
Qx9U11QO9oOwdJrOh8qoIb14msL1xGiPN4m6fdwZOVzBDDYdtlyDW2X/1WxqKOmG
MKelHPNRlxvi17sktzr/WmBvLHUt8T/08Y3yMzraNgk0zIQ5/Q5a4SimIGL5qxaP
PkwHsqN2GxwKgYaZObso3qAD6ke9/Gfw1qpeXM+kv/0QeQeQc1aRLLUobIfjI0n3
RtXiAgK7VX3Czhoh1s1TwNEe3ufiJ67/jqxPEn5aFRLON0CRWx9Y/Ouo/UiW/Pig
SliL6IKJL2uGDPD/RI4vVvSLwm5U94zJWhHfcQcRmaSDWolena422BwELOZMJInj
nqtYZB7ksLfgoo1AtIn5yPO/UrO+Wra5zJnxRiygLa1FdvCBCX4E9Ctr2d8OIPge
OEuLKEutoEKuV1Oj8Pi7y4Loso0OSETTQZfDpjnIitcNDFLkMeKQHD64WZJ5xDzp
qpGYtAVcQ4bUnqVBxs2mxoBAAtWJ/pnCCBJZo+YmEXPElF5WcApNr6/O7vPGBVhV
m+SVU69Fjqyg096HIiP6wsbA1zFFaR95x0NCQNK/TcfClGf6OxPgxZy3qGGQUMRZ
rSnaGfAsHnzPgSdhWV5vhf3iEuXEXGny12DqIKj0uhbeUvV7rWSOPaQ8bXNU0IO/
FXd1bEwt5DsyD0nRaNI3qnE3dXye8JLb5UFLSJSNE5CTzQeHKGKpUmU3nHMF9wX4
Ko51YtMe86Sx/j9eP+RQbvAmV1UuE9sLeNVF9ZywAxSp4SlJvPOmBsfqFpt4BX8I
9A7gY6NqGHlpnImjtPBJEjeGZCn6U62E7+qBi3zjXMmJT/TuBkKDVFoyw/TWXoVR
cbUBENxVcYV2ZmAxDSKA0f4HooeQc25Q1Lkx+M5FwGXwpXUc6o4rf0ipyy7Nh4gS
3ut5FeuUC36ZErYJE0B3Dumw8JENvwzqTYYRU6WJa77qL/osaC5LDYqSTc9JL0H3
TEYdQU6EHdQwjQZyhEUl0gc4zWVO5/T7APQfRKLtwWYtMyCRiepgjt/d534LNW3E
oOXpq5MXjEmPStsUAYZVjQVFr4JEBwvgTyoJVwG0cCmgpmh4qY/4fg3IzVlzj0y/
Ch+2uJ0dutuCpJHLv4lYrtgKKVZEYmGS/yhnyYa8BEF/m/Ps9jnrAqHywzqyFqLf
KIIt4qsJbxGEQeSwZrj81LPWMX6o2QYHsjKhDsmFcrNs4JSfhZVdRFuUgI9IPQ63
MGrC9Gj/g9aXjt5tDzZSXqQTjpQwwNerVYhQ6SdKqtKi45LlLrI/07Cw3NhsQYZs
TbGtUv3WgcIi5zGRAJWywx4aGfLB0y9DLwdTbc+C5VkGDJlyRGiqGWHjvL1Z2lY/
+1TkECns5SUcy1/McgRmKLG/LsA9PoDkEX4IlpM40ucwn2Cvg652ZWmN45Uogn/x
pEcJdXXA8E0MxDIk3xTHwzxebGnl7/pkCnNpWvbKiFcnwlzTsdSThkBn6i0JXsQk
wiyGuwNCcAHL1NpFSrVDWUG3dKPUFwKOvWU3BSjUEaQRAUOQ9pJ8GGFVcJAsV42U
H/ShpF/SrJvBK607XIGxp3Ivp8OemOFurluya0xXWgqiQszy80irMc1PzDZDB9d3
MWm1Pbd85OsqbbViiX6vboVc/D2rgevy2Ico4mGrRiNARCgMq88UQNmB4eSoYdLd
i5ruIJxkva3zmG9pypalF9Qk/ZVnvaYHPRXOK+nLnTJfPdduwyYr0WAQeD4AINsm
7kHJ4h3gLHlqRiqW/LpOlQ==
`protect END_PROTECTED