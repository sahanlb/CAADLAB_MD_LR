-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
U6xf+f4famSUEUO+OHRHv4r/ZNOS2WmkuuZNS8G3BOvKVWlIFYfq3iZVbDsM9oDU
ZSo+iNAO5v8K0oUl7zKjqnP6k8mLkXroLydjNxOAx8KtRKw5rz5hS81fhnkiTwG7
0G5LceQfUgDdNBADovWdYP5xUXXA/Y7X5hqPo48MmWI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7952)
`protect data_block
npWm6cVaZCnkNGSO9UaOVLTkP9i8GVzbyNEfBdvDaS+53c+Rek0AGW/YhVmZpi58
ru+m5QcBfp+oPCG98h/763+q9IxiZ2dmP0WGp4WYRQLtwyaTEFNVD3ccOCklp/0h
ca5NQFfvT5tvJKHnVwrIk4eazy31KygyW8ZRrJnt6Y0A9grs1NpZ5BdZ6OVN/OYq
tTzAf2Uax7h5dQPYGwRecEi4+O5U3quDTSHL0Zn8wuHUJFQgkr3sXE35Dqb01aRd
7/JUHGtJg5Yfl/VTadWJa7j2Tisd9ZC3XLe1BUjeSvvmRU6DUGsMoTGF6ycv7NyH
PXrsmwFX2hsUf1R+dK/CAPd/pdmXeRS4Rjo9UPDOozP8lkOnkhcoy6GENctvxlKj
S1Xxy0pXzZ47MBRKe9qOIji4322HF1ja3ZR+B9rTge1fwO7KI0Vd1iFQvxUW5YtK
Ja8XKCfSswDiPwtC5SbTctxHAImSCa4xYjadCc7KiX8WifzbAOS/zhbnVUGL6VDs
gY/hiJKjhRvHVn+WoYFMFghXLBQ6NrGBlucdLujZKPDNSAM2KRi+lLRYBJ8UO8mZ
lfPYAk42fjWYUmVfHhhfhmZL/PaI+1A/mXE+UmYqPYFIJqI/mGbUi6JhMANlZW9M
BSO+Y0ogF/kU3RRgmovMxKE58BO+KHIIQo7+E1q1acArsHQw6jq7nmphl+CW44wV
KsYOHvpZ6fjzbacQjGaaqxdowZLzeyyq6F1a0UB5yuiidfOaMGx16byKEgywBKhr
ktE2gJXLfl4VKxuuZKoi4RhjtvEoccJgKm5OC/6AUR9V/SE/IRHZn1T8ff0St4Nt
7YFmeFIwmLyEvWXJGirl+47Xmc8lEoBRW8a95aKBsJR/0Pul3mT0yMgsVPZ0h3Wh
i5kNxet79QPw8aDU9M4sWU+y0/MZbIb6Ejy6kr8ReHrG993b370mV0l0INOcrUzR
yLTJnYLV7SgPtjn+uvPatdoacvAuQ7OEDU+ZzF+uddYDlyu72gpCV+gyjQTnyfIe
3MzSvcBs66FL3YrKDkSTSTlkuVGNkaUCyyBJ/MzpIA27AsCmCQyPGaKZoYykLSxr
tKYyI3JqCROUuLI04q8+D8AnUcTMPzk/AqfDigqRpnKmsFaVTD+ElH7B/ZqGRCMe
gZRuU259jrT/xWaORiERP217vkFQPXYi6WdZu53xCE6XeybGX+mxFTsLOeaO+IU5
iE85AiEfRSJ/woQXBmHvUS96cIOMq+zZJFyhKHmUqy17ldkldZYOzg1w3BwqnNdP
OD1ROcYyk9ANprjfFczrKyk9BpDEvlNyZBEoBh2x0gNow4SmpyxIdbWkqtyogBaC
Mlfs0lnnizV3N7GFqkyit6MwULiTwwBMBB5c6Cqt1134yQWkbcOq3i1CJ30dRdgc
lFNjBIeN0fyPtQSDjG5/luJYt9iJIXkFQ5hdz6OGI/etKfu+V3eLcxQ+/XIGhx58
BlD8oeKrY6iSJcm4WBLe4J53P+/UAuHKmIpdYFCD12PAlbv+FNQcinltqpWpzOMT
j8BN5DnG3RjC2Z+beiD1owX/tClXpP4bZUoxt6vn3U0SWBaiAJ9+wuKa+rbJKmlg
F5+aolCEG0znYz3ETRbEy3KJ5ilhqbSAl2nOfuV+Zsa+tO9n+cGZqRKBSqW+8+Hp
Sr2eNUIkAh/szXQhToSthDALMrwF2n1LFoyP1xSSRgeWPGPODgB/IhctL9VNHoae
Wp7j4oA+avWlPodp3ZZABfiYythb6j7uVhqsyWMR0bHP+eoOsJy6IL6I3r/K4SsB
0CJeSmldF8YB+lOIMMnxiMzMtZuuBggzio4jzwLgmyx8AZS5OCxadzgdxD1XK2He
jPWOl9ZTNl0P2t7KuvnGcu/Vq0ApXkyR0DjYiB2tT8QkqZpL+MmJcJS2gIjyTbPi
Q+yKQW0s0MO7/WTcdZOkahVmKFwRulcf3xX7JazgROceSgahr/V5HBAv05pUU+oR
WYsndr02Bga9KvP6IiLnkldkz/L3saxUROBY6jS7CwtzpgmkkuYeUTDVS6dhOYGr
6LvE56NSDMUVgvJ0hwJ+AIq/sA1XchzSb51ihBdAZwxFBhGgZ4740fBEBLI5dhbt
E1x4RZtdvg2pdaSPn1DDcga5/IL/uzFLGmgFLs2zm7Ybz7x5tb51O0KmBiQjKhb4
MkMGHxLOJhcv3nljk8ni6X4Vbt7gZvyTrDv6RVysMtAQuiuvl/9jBYj+FEcfTwfM
WCnfobYJ7btw7f5bOz3s31X47fLFd+cn9xrDGedqIlyeSXf8+PNhjS9E4Y/PceiA
vpXCqNAfFTQi9bW/MPPwZSmUNOLMRH1LHiIupSuKw/xY42AvJkHJ53/6w1ihlQIl
jp3bMMpCfM3vqFwn/eUOk/whjIwY4H3GIGl/QqkZcLyGWp7/c5bmNbXVrdKelMNm
vCqySm2a2yAzso1GrylDyKuSC4UWfh+S5Z5W4gOBp5OntCXEkqgZM/0Hg/Ln+O3S
lruZftuNrOAh6sEqHYS+0nGL/iEIzmE5XaWzf5sxoVaTxLVFzWXaQn84cLRjb2gi
yawML0so0Kv7/P3K3GiCLwhNxc/vjKrZvVyWLypz4dhzyMDlBIwRAOx4rlRMcsWc
aIhnBEtU/e1i8BV44FfnF3E2aKm/f41CEK1rm2M7kNZqbQaYq9v8poQVBVe+eSfu
j16RnfqlqJ7VO+vHeHQloUv0uiuwgpWUHJNN9JR2iq8wkIq0XrSGh+k8OIBOVXZW
OOfbeG+yHZ6SOefOPv2ebikTCIyUVzyueijELaH0sBNT65slEHVdcpsrPY1vwD8w
roMwUVDdatE7gWZRdfIiEGsZbtL50/J0yq3MnUV6E7s2RIEEqr2hHGI7ABE6W3BT
o61TZEq6o7nky5aHoxXD4uqaDkHV8QbRBJLTTuerTzEsdCWC7TIF+TNdFon1MkYL
oTjzPV6zCBbt5Dn1tGX/8BjMJJcbX34slFf6p0GKjPOA0icW1qxPfo2ErxVn9ts8
hAoQS/OmR/TAJo3XvJWCaxG6XNKfA4lEccgRayAUrj5fMthPr9qt4TORW+jpxQqN
lu/hXF9gShvCMzwmn4Xr/+uHJsh3ZK5Ln43J589qB1RfNLDQrvkp4dIv4vc757CS
sSx/GLAL4YWTALzGKrkKdOS/1OWY0TBa1qaD1DrV4WvZuTThJuKqtnxQhLSml5fC
NuV5ONCzwB+7omzmhJoZb5GL81d1SlNQqAjHlbS945gI0syaSin7hg4dF3ZB/iyM
hNPXIY4DhqvA2fTimi8yhvm3G2veo6VfGZ8Jjk9CsIvtSTRu3RGhomQDgNV93CMG
zqz45uoNbMmi3n8rph+RHg9lVhPr0t5cHS1Hux93gL5P3EnlUub4rTaDYD/k5s3p
6SECIGG3X3bk7LRYGnEnMhPz2NFA/XiFSYIRqCGfCzpT6pfdFOpqxXdycyyyv2uX
GKbH99ITDz6siTwG5V5u+T3Y3/y1QF8flIO4bmxiKOZ50oazSl86jSr46tXX1ZPE
iByNJqWaijUG1unN7gABUv4y6TAVOjccAKoPgTDxxoAjHWI+NMU7js/EZyd9NZCY
Ssl4ETuWFqbWyis5HKMbeehzIpif0CKByx6EQ2LpyPDHZkqMoJQOtQHTYwuQ/+8S
iuLcDbme9p9I3eXxDM1+inmOLTHhnB6Cb8O7dz+NB7KxV+HOZSI2I74i0xmHMDVY
occGvJugLtU6TLGmOME7t/R9h4NwpIlGxJ1H92ULkFK2S+IrMRYbtoAPHQiTtdXK
jqy/jHtNexLWmJ8Wb/5k5AdiFy6B10olEOgcilfZop1Qm/0RONNgJ077AU20QBZv
awFIWAN3Qx2C1rvsAUwhaafr6hBWHcmrFNMgSSY1PN55R5FgtolyWfJbhlUuijWn
DLhsYtjJ5wwIUqFxpd57ZBmym/LJehpiflJLIEBvfn6GlZ6kOL7AfTRddEcLuukc
gkjicSwCl/fPP1SRkbEU85Fz3PfSxEQb4qFce3wh2cyskW6TQ5nqkmh/QjZEGz0r
k5LgCN2GiClsaqZv0tjm5sQ6WA2U5QpHuomKKxGO6FNp7HEL6HL3edYAhPPVs+Ub
/PNkJ1u3vioOPdaAY4EogC95ND8U1TT6KLkAsh4jQJ6YZodNAGmMKooW15yMLbtm
Lf1YNLvqInvzS5ETxZ60ckWlXvTZgqr6aEq3SdLQvaFO9/tgtp+gv5o8h/ebl9f/
Z4+IfQBK9IATD73tJagaxPhoyRmwJtfSMWavexdIs41UljXOsYgjpII9V9YEWTFV
HXmwhYgxNNLdB1Gbxa9ul1+ZrzycsnW/V9nTOgsS8N/qtRYGtzee1yGNOrjGYSBt
c1IFDUTgwON04nvpGc5FAFAeR+GKX65RPHpf8NdUr07+IMKpe4KegnrWiKUQnIyb
1QZmfNq7T8GJRRwNqiELlyogx+JcZV7+W8186sH0i8Z/e0hPf9GaYkD9k8ZHzniT
8lrqyZxX1KNhhm1mDa8CyzX6puQef6d/rFkyntCqAbdjdZIenm8VxL4LgOeIDoyO
vjFBrUzYn7QbitSgjxmfDc0BIOAQ2aCiCxQHa7zFJWDMvth5/KlPwctO+4UGlVXP
umrUlNR2MvO1ewbqGZeo5dFtWoN6YrBq+zcRJjNpuUBGBdHpr8WWs2tzRSlz7jwN
fZl4uURO4XmmLd/VIqsu0i7a6mFSiJD02mlxScp5CCYSRoUh3y2IXM4FDeAMXKJc
XIrPZWrOHepGX30QMoW1sEG45HVD7F0qMA8nVMtReSSTpCaBcGiYf152GWAmaLrI
gPX+h3JJNcNCFe6uGxjtqFjC7REUGMw/fzZzR5DqTpZLgFu+XxvvMXvPoQ1qfhBJ
1nbP9JDuPHyMxDK66pqtGQLh+NVgZ34T14xVmLalN1c1pKZpDEs5ZkvU52ixP7TP
FRMtg0xmPzrQClahngr0aOrNzFETF8SpyJxoEIDBrB/hChU12YzU7fTNNlyJOlQ9
CMtPxGRUMLm0Qm0tX/A8eLRmMvAmgrJSqQZ6e33rzQ9t0ssLyvJ8irpdV/h1ixZr
RgSGEV/Wx+ed8RS4CBvQYpAW6jlH0d77qz1BykY9svzctX2uzAHQukdYrA+sC+iq
uxJ7yqW/aismxa/VeJN1MLlcttxd2GaHzPHdvjDPogjuUob4SLrrJBsl0VlERYzm
U+bxgiBWmdxQ74vTi8WMJwl4zAH5umZccK7q/mI8t8DCo+S421JZ2yJFtl25lITl
gurgpcjE7SG2Bju8zRYobfTljgDkMZonBS8y2uOb54AEPUDYLgQvEkTdpqh7uZaS
rg9fFXWBo+FQTXIeTGvOUWD9UT/N1epYSCy0ipuj5nny4W+0CeDbhv7Plxd3OHVe
kssVxWaxyig7AIm0JyC7kIdTnq71JD7ZZFcw5VBnl356aAA/w1DqoLUcrnxIN0sO
BvPCD0jPUdjthwJnFAd8Zop4jybEHA8+bm6ZJMpbVpVyNtHukxTX6+3IO7PX9Ldo
h6KGlRZRI+E0cYkMyQ4CbCeMRX8Cd98fYe8o7BJijY629qp4as1SBa++iaofdoJl
it8t71cMNg/qM6TebM3rON0RiHVu8V8fHXHUfB9oBheEJaOw0WptQ+AaamzKjksB
2mCOQ9vgVPj8uVHnIGxVQTrazv0OWoYHWlUobv0ZW1ROeUhGrlv6PW8NdyW+/iB/
b1p/ez9dwd7pBRZdVjX/KtZxK3jZbxZiRUq0VUk9r1pPInxjqn99S9nP8OYw69+S
5y/EOhiEhPX0awKOrMulJZcWg2pI6JRC7h0ZIXxlcf7KmXGInKaYK6y/vXMkAFP8
Mx68xCuiqLeP1nFjcIcjD1kE8hvhdcc4pj4MxyPApYiUAZwhOyOiP+mNPfEXjCVf
nu4tGt7sKJjDlS6ujya5XOSTBoRRq/p0kVdHXHCX+mIZJwspPlhDaTgzHQl00ycf
b7ujUogs65hwz6c1QrLnmjZjRg3uIoDXuPqhSNQlfV3YBv1JTpFtyg7zNVFGXUqw
K8d5ftE6JEhVPpH+ZR4paLKe8TDHvbXNO1iiRAZMLf0QFaVFHv9Szi+RGqU114Fa
NfDkQMA0rtoEsI9pD0ID+YRUTqx+Us3Uk6ELW6vYxl/2mUE2U8qY6UYg4iUF7+Iz
DxvVLnN0Tq8E2yuAboqeSf8pARrpT5E0J77APNJ6Rx/AFD2Le1+pCLTqQHYgXVz4
SyADNEu8HZFcATjk+urJJivH9Lt6nzIIM7E+EyGHb8u5diEdago3fbnwvepKX318
aJU5qOy4MR/XQh2lCRdAF8VETN7MnogzgSUhP8bkIMTu4I/8ZLoLOdauXuMJ+YtE
rY9jPNRvQ2aVw+tFoWw8Ob3AIuxSjUQaYWvTvQbarS4X7RehReWdhnYye3fWr4jg
1yx3T/0Sg2mtnVcfmjyJi00wY/zY/yhRDskvOSUGzubCEcboygPBhGy83kFa+3ef
Pqi/rSKSJWx1oe+8g5s/UDMZcPfKItY/u0SeHq8VGtssNRMhYHxUxhvQXxY39KaO
HDh5QCLE0QTUOTCGeksDX65AdoHwPDT6xKpMsBWUsX95y2UXw+DB6nzCuDY//Nbw
3dZe7nxlzR5cDh7NAasvGuNdAKKi05OarQj6t+ZtYHLfyoxTV0O5J7kC3GAePUVL
uBkdxBvlTUIGCMBDBiqpEpZaAcSn9Duk+dXWoRdmc2uhkUoVawfqbctYXIGEACh+
Cs6hh2QF+ROX63NVYSaq0UIOU9jYvWUiaPddmKrAl8UuE98buNhT2gGuLEDSXuq5
FPfra3b88FzOYiLiWobE/OFaPhtPQK0gB1RRU44kDC5Mq2vjKddeAFrzBbVH7C3N
wkRFimW8jyTjskFkWC+gaajCwP5cIJApT/34EVmCTkI45fkdu+vnWEH4BenXr5mm
sm8dH53nQjzSK+Iyg9BDWlWdWW7n3BdogscweiJZhCv9NOGuKAjLFug3/cVS23Om
ENkvdsqomlj1XOsukcPydlXee2RQcdGABNdZ7F+wKaYVfAM5Gw2pfvxeZ9GROPBA
4QErJkreKEvHGqQ8ckJaGndtToWa/XniF++CChyty6QhG47ciEu0zKq6Ur9+KZRH
5zmK3mbdAHPooxu/L8InrKBu5ASzUbL4tAzH+iPs7jwPoVdeM6OqTDwpDi4xnE+O
V23N96TWBp6mJgS7cdni8BnsBuMStrNJGUUNhZyoqJeGMsnmeRM5Wsd1b3NkWACc
UyRdllMxR55Ao9PbLyFm4DH2vMYpw+UEsgrnMTfRazDT0BLSQBYGSNbDPbbtMDob
aMaEhb7hBahewPq0MoDmNySSdALZAMdBUcsczrrmiOaIhSDwe6BXTNfcGHxsMgrA
en6r6vyKsSC7r9uNX8PASGzGf6TQZV0ip6iYNjESNR7ncQjNTIt89GeiHEadksG1
U+0I+9cygnvg0uU+ymmXVVrKKIzWRgJlLtQ7OiN131R4TbqV3l5gxuRorcq5KJaG
7Di92XhkR6DfCTooaYJV5rYyjy0kJIA5+cVSsqcb5fSpAxPwaejMe1ATLlPMBGSd
XxlZI0Nwn1xiULhAshpanWAMOmRwKvFkXLfjf/nLPGsR+0X/by7ZF44Cu34BkqhG
oDJr9psdLl5jtf3UKVjLfSdOHiXtN2RyYFN1A/IG1FEFMlOI0meEAlfcsNf03oa3
HC59MH0IbWP8O3ptTszxjcYJK/mC+8o9qVKQZ46/9b3BauxPu7ue2q4lLY8BQNax
jVLhyx/QxENjqu5i31T9xAhCdnsNaBLFHa0LXYOX89i7BGMf9w4FQvob7H1Pj9T+
01Jdr6x1rYbXN05Jpsis+a0wgme5F2a/zqz54jmfhwq3kceHiO9YbNpJ56PKMzqq
aidqIYY5EMq3mxIw39FrR0DA6JBtXE5/5cekwJPCOb5gxJVReCY6okW2lRvR1PFf
A5qrQK+KHTHKbJmRP6Q0MVieHjLLCtvpRWGmR0PBFbv0mLaDtc7+cKlv/bB9YKwW
hm/6sbJcda91aRp9lC1CKhbEAJ3ARG0WiUVdXMoo4EYjSMpdvvKygyZ/RZkmkVcx
4LiR/m8nJBFtZTBln2pxc6f+tB2R/FshwlckOaBFpCIrlhyqtCHqCHvoXFp05v18
F1QxQ2llPOpXxRQ3UVS9eZDM4jEzOka9AQ6NsqouIJeiPimYCH2OCgDbkw7+5xJY
u7t15UeJSo/WIzQexuxHFjWyRZWvZB4bd9Tzix+Q+NHCMDmcqeYdx4XB68tfGbEw
5fUKfS4mxLNWX5vtWN150dsG+gkVRDu/pU2m2RR7fi2axkT6bpH8yAIU/BQoecmi
ovFKhaxSY/tiLwHPpvXnBYU2dfDaDu5btVkUe0V4CUd4aETW3mC5OLu4BROFjA/2
InNwG1o2VVw5pyWG+nbVZzYBhlXQaU9meCY4fRzaD8sTHUThgdMrpXMV0WipuwPL
2c0qettm7DOFLN4Qhh3lBPNL/FIUsA36ViozoQICtLL06YXfPNAWLkXFbUsHgUby
lTHRqHoVZQ5LXPorJvyA1BEJ6+cEZE4DOwmC76vZB9Aw/g4VQueMrblYCt3U8nQ0
hksAjCj0jsNQJlwrgxJuSX0HceUi43ebisrtGoyGs88/VDS2/QDH5Sw6OIGX9700
a5o1lHXu2j6GmSLYmNgC7xSPv6ZHDqkhZ3g57z/ZJasee385latyja4tC1er1F7T
VQAwjcnXsX2hG3qKqb2F7XtvHVvoL5mzU2w7aIgG2No/LTeqkpXUjHQtVeRQqe/W
PCNQTYm1Uo4Q29cXCzZ3e9zspt4uI/G0zbiWarUB0R0Rh4gZMujBQA2EdGKefIQO
c6/tUITtcCskUM2+Yb4ttIg9jxQcV6Y32mARFr54rI+UW7GcSsugmQc+aw9aMw5M
LSO66pCkLLHadpdbRTxik/LpW3C9fjQ2296GCMBwq8VwB19jjbLVK5vocC2Z2F0O
qQiBpGHe/PNNBN+niIcVOOJKpOCtK6PeY1SxSx2dugUam26xBc1Ytn95D+kW7uI0
8DQaelIdO92pAAzEhetsePfp1vEnaivcGZBknVvtc0NxQAYwzUrIP5RSKq+g6TOK
+qJdu35oWUxigZuupExQi22dUgskIhDCDUBL2olTPPS26PhLgkQAmJuh4e2wNY+l
sG3UfJ9O9Oak2zXj5lUB8KgOFkwOvPKcKJMWupo2pWbFN1mapF/6hXEcWoXQy65q
LrHfyNVfS3HhK82Bj02ZOCdvT+V6+3HVqbiGHtCJJGeQdvQ1hGb4hCxlO0gJpreu
djhMYRbHbuhTBmgNpvyyl4b3wO5BiA5teX4J4cbD+2vOe6VV/QVqusTiCw5FKsVO
w1+NCb3NLG9VP5UvtqKlhB4klIKSeUH9ZIfKC+7MgfONW5LqLXbVXhfP0Py1Gy3U
dIpE36lMFw5XYshR51o1v9/C86jXXFMyAisawwG04XxD6vScmCNMr8iJbIaFx3Gb
AmqZpsGF2Z/6rd5FP4HkC6Op+8cOG2MqJyj5xcaNE/HUDEp73UE5zwnFYcpoTBlV
ZTz7daNQdJ55UE0Ws1+VaHFkHSc/auGwavp3yjW3pWnTQLb2GuV7zYT/evthGfPH
d8tgYIfHTikBOrzAnfZlO1SV61MOVO9ABJ7YUG9+IsOtIA5TABAv0ncnPcTrevKt
qEg8k4P/1HzUTO6aqChluZ/pXvv0ckfK6rthW9xVNhv2+q18wAoomUJ8Qi0+5DcX
MQTVrzH5Ut8B0BBqBRkH80ofTJsqMFS9FqIkIdpB2R93okDA9xQarh9vGEA3bFWO
MYL0+yuKL9n96M+5p6ZbB1m4ZMu/7gxVaY5elAJXkGb8DIDTb3JyvV9LqT2FYZGy
erLiX1P0fM999mdEhe4z1UHyUN2OBHJZj/qI4ocgkmlAu8YeCaIYj4mk3xzU+L7A
C1eV7XU0/OhPQssa5eUeW9kZ7u6TCZLKdAiFmiAFBqc7rRBQFvggjrKE6dGjYutl
VwdQt78dYanbv3uNOaZ+1bRKmHagL+FqyMIm6HkAaFvdsKtrATV663hOyo2OJPZQ
cOkXW/KbwRR4TJDPxAgfxBXCVQYZK7Auqqzp2my0KdCqqmPqeekPqG28vOf10j0h
MZKgMKJWwBTfUSfAA21lWvgMvz5IE80jvC3UES9fpmIYRDb8Lj8KxaQQTknabogU
ATf6famAAtfLXO0jgSgd7j+9gccgi4CjaNUSiXuqnwpfs1A3ZcvQ/RCd2brbsgRQ
BllYrerQbirBW9/rOGeGsUux6HK10bYzz3eYA/jf/3xDZ4wgTWQ4ZQtS1iPMA4y9
B46bLd2Am+MrC8jMJkEX+5kuEF4C+jseLGbw80VLyHJFroW3jttm88OgGYD9ZUmY
kRFfpTfReWXuuXJ0faodMesTOVK0mViWGTD5I8/aiuw2BklsGVr0zXIKM+OjWXCm
ia1YWn5uSBl8BgwIj7TWIsSlzLwIyo+UvBgCtVUJmosjeXy/zdmZ+Jno+aWXfx31
GvjJEzYmrPmiUmyIkzu+/P0Nk7qINjU4faRLIbaaK68fHkfxxHV1N8853ajax92h
CU25mGyuKiXBbGrNaubtbfsBfN+DezrhyoJsxYZENCU=
`protect end_protected
