-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
H+ztwKonfJZ9rX0NFNsZOl5L+UPQtQAjQez6fNysXmmwyrxsuHtbr11LnMbryaxm
YMI1ngSYwTqAn732E1hc9hXaDeK8tCwE2oxWooV6C3K270L5kzzg/a6wEoh4Huum
6q0JJ4ac5XwWo/FJ9cz+ErNBxrdwBPHcZR24z2bYUdlFwqKIcaHVWw==
--pragma protect end_key_block
--pragma protect digest_block
PRV68AWOAl3JkI1KlMJsOUx12fI=
--pragma protect end_digest_block
--pragma protect data_block
vLFTw9dGuxkK+78EaSThbQuC97OXpnQlPFf3ViILHBwWrrEIA8Ad57JlANwXoibG
3WMiKt34h25lXeRM4NI/W3rZNz9u81zJYOZOGjMA5ep4dpdyEZ1zE/ov/omKf+HE
ZsY/KlhmWIOaUTFgokKF02AR1gVHUsNkmo0YNkTnNVxUIcYBop3JlexQH1vKZt9l
za2B5+sZaxa/dFv0XA310hPKswWMW5ef5bSd++hR/qKeRvjmfh+1UMiIX+ygl3Fz
5xuuMm6HZN+Ump0dh4diC4vmGCz+M/T4uoPvM0J1b7MY8MkdJAIntEFEIrKisDn8
IRAvwuhVaRC9C0sfngnOW50DntMtlRriUspViwSWPV+avH4UemWJgtOjYubx5wjB
bY1vUqBnEf4I05E9yVspluLREfT23U6w0fMG8ceI5n9KO32WGkztGfg8vG0zE0Z4
Fe6NU0oq0yXCjuH9jFE5EzjTPUVRbIqkc1lCKu1y6s34iGmZBOJGODkW7Y6xnAGw
sV8mbjknjhAyDlSEJOuKtPha2JdrXhroSltrTzFzZhhMg8CzY4aAaWPTA+S+VtZm
1zGopnzJ/G/UxgMCKKn/ka+ryIbWykbsQSLlGJLA3wHbP0W1/tUJcC4jWuj27tT1
/SktiUzlRO/iHU1i9vRDKw5vRQNE/XL7I+tVtktsTIN7R1342x6UsEz3CuNIHTAx
CDYGsDUJ0OX6uwi/MkDGQDHDiHPOxlr9ELzpEAQb2c2EUrix4mmHCl5kPx/Ld2Av
tOutCO1Xh2i1qkHjAds6AUYUmzxTZTfFZAvZC7LKMSuH8ReKhHFin1J3A0j7Y40y
ysVy8sQXbYjv07mdwRPN0fr+wnyKKF7CyaKGDj0a4Z58gRLHfRxTozud3F+3uqgV
xvrCMUz51pb8uvoYxlQ/bAeWOe6ia55uJV2cpCMfoHzm8tjdikDpn81CSpiXangw
rFkGyw0idINlUVnnoYuylXbQQ0AO6NgMSfzVqPXdtLGn2HGynw7h61cNC8aE7eeb
uAmzJuHCDoavKN4JZ5kFSH7Yt91v+ISOmiO0oOqRqHz7CCpPmvZy85N2A4Y2LhNO
Br0C/YQhHrRJ6PVm78XABzsEaFTg37DwOi3cXpWCy9sJZWQ/CoSoPErj5ulttBCU
eOSXvJ74Uo1VyP3lxxsCllUfXaDaBlJkTi4FpclEFU6ekiNQ4dS2Tjsek9ENgZmn
ZAmrQY1hUcqYW461g7piUx+F3i7z70wGF+4QtY+qEcK7RTFvjzGMnJG6pv7C8Gz9
Ceh5GdQ/wFsUDx0iIcl/VKTaYrMc84IPAXdBnF3tahao3aWYo9FnxFikD+4ooi67
4Je8yjNCCrt2daYwLQiz15R5BqYff3hp/6Wqjw9aVYMDu/wAWI98b6K5f+Wanuqo
8VpQx5WQozoBflWI+FVYAzz+JEspPCKVdOrsVQECdjyKJICf2UEBxLwxAiBt9umd
RkjKWGOFkEZYG0rxBMw44B+vYpEV1cfwmSY0oG49r86AqdxdNrPEqDHbsizbYD9x
b9TvJI3qQ1B+DvHmgiD6+fCrajPIk57A8/dSEW+/mgf+3t3p8SIJZEZqCXqgaVyo
m3owt1MitsKvg7+TzJjN0qhtKCmWJKjoMpfyv1GM45esQvHmYcsQbcN/8dk+fdxB
/3r9BxU4T3wtMiTtL8HVuzAtkKZRYXA8KIUECTPS71JVptJgcWow1IVxDTPSe2v8
xNt4nweSGoSr/n7BjVE/uM/X3G4w1uWtQUMT2xO/R+uNRA3EpSsLXemjdkakz5o3
/DMldr3ahjWrYv4cvh4ppZ94MwPm4jAEOvUn1XxtHKLoDmuEu0mQqxai2y8Wvi3N
aXQ6QzMzzYAAhLT9pR7PK6S3YOJgGv4keP0C8xmBPetdIn6t1IJqlfFBTxFMNhTf
0X2sbAYHUos5L/22UcPmtnfM+pGSQ2g34XY67zhSVYVl0b4zZs7kZhG65Lpb9ihF
j3EOjk5j6ZWr4EciiIrBtgjF74U6o1k0UPv7y2RCn+U61Z2/gd+AbOphx/nFtRi8
QKQHgSJqHoDQMJ11B7u7Af+waLZxgOXfWj3cgUwB+Ck2FHtfQG7hwVdF+3e3eoW9
wD1ajr4z3V8foxaS4iteQBl0+/chZnhbyL3usYEUvnvXMW2oE8kmeUb/RCG/rQ7r
0J3ypeanXsxBP13td3NPw2U2NlPOey/q+wTPxvHHxLRW/AObPWwiA1eCCb3KyMUB
QPpo22ycZETUq2JCngA3o5EXJP6obsxjFVHi+urE9y+CbKGHMbrb24V4Lt6Ushis
pgubDJEIavQXXYTp1eo2M4TLn28Yk5l/1X9FvRIsNCAx2ToLr3sf1t3PFNOtqaSH
oarHa9K5jvJvHdywVldCRREaA62BDM3l7Uj7UORNsWX4x5OaARTElph94qGoG5tI
2ysE7FHH3z2crdRBIz3MpWEr1f9gJxHhpiIOaOYILollWbqZnlqK4AMWUqaISDch
cKNfPbb28V8+s19CCizr+aVc7IWSlyQW9U7Cpkdpx2uMPgGHLgrbepUPzsrWUxr6
QcbtYo4TTF59mmDjLL3d740ncNOiN2EaOyIMUkvwTkDjG6YRKY08Xuu/Lrp3l+4N
J+uvWuNrzijXEbSOsGdT2/xKdk63K0xCd6pI9KvihgkGjG4ije+tBOST+eUWK6o0
zYY13XkBHSaf2kDrKPeq+TcecCyWgFc6yMO+Jcy/zHgBMuQW9K7xmeBf6L95oFPC
iDX5tkw2NI/LNd/LujLfb3gCm28ufZntJBlhV7Ib5VcVieOWgxI33+DHwj/1KTw8
ft6zxAdDeKhYu3R19Bors0KCrQWEqoNX2UYr1LxDZZZP8GfSLTLLA53axSD41hgD
c15fADZPkVppKav9KZrPxwNp0EApxZB05x91IS+b9uamU0Di1VVj2m54wqv4MLea
S6yhTQosVg4a4Ki7GgVElOINaeu/vOkzInYjFowdilBfcPE/NGEWlEZYnFwVj6K8
6mDQBZ3Asu/P/z+u9xhyqAr1ZJHBSqBCg+kSgRfNcRoYrMt+bsuCK3RiYKBXQoTD
QmVBWmvA7g5kcZu3QiBR0hyxKKHv6vHLvyJ0AIJWtX53DzwnUFhhpun47IXJm6/v
tzDzVcx+q1xYsfOwM+AuH3/9Spckba3Q7mfeFW8GIiwvNcWSBSWvcVC+atzxSzxL
H45U73v88qYBKjoXgA8dQuFSeWE30MUAQCR+9J24dNzurOg3FF27GG8Embm3KrQ/
oK/0htiL9gZsnqeb/H+9+IbkUOQ1LYuoaZjMaLDn7sqX3NT51PguBzXqu+sjz+B5
e6SU/+mHLCWxr11zI/JcouCgN7zzQHq5/IgX4CnydrtjuCryxYqySXSGjAoP+cRq
jlIc+2q8g57zvo5nJ/x4XFakMIZfwVZfYoWwmofos1Ula6chQ77+cdXHzNLk5MA8
FRlCmkPAgLI3QCk7QZuracvOu5mwYcNMOczxxBG2tYSnWrG+XyBfJxcb8V3ONHAG
FwaGIJUtRv3kOWuh8wfG94ekKUoRU29tou/Yb5C+u8vSFOh2PfPCxxsWaaIfk1pe
zRh3Xmv4ElZACFFBwkHG3GQOvF9+NUE79vTX50D9OV8vwlrSQAYrXa5p+VGQ9o4g
nv+SOyCdKq3m+DRkMM8xrCKe9EJ8hnf2AjUhmCWK8ht8xrYOsQbSGnWKGms1NDTv
0PF1NSdrgtww6eAgiCUrS66pj/myLjpTQPyCB804lFApSQPPixxe3yONjYAoigJY
tdj5/jiVIoksowrUEUzyAREKoTAt2McUFew5Wcc1JoboLyO5ODghBWqW4AuiuRMV
SqH17dvbm9o4chCN+lFp8svBwj87DXpl4bTSOBvgNgPC7Y2zOgdQJ8wrjoy3I66x
UCHfA9uA0BSFCnnppdVcPd147wv8qUrD6tnd0JSojseVmrsc40mIEDDhesrf8oYf
rje+OHIiAytn58w8e6LHGolnNPuhA3iCglW8d8ZWWAeiX6UmhQqqkFSKyYTF3v+p
i8kruwJdwL00tHoASCe1qk0gpQUTJVlJydvTUFfQyfbl6zBR54gOm3LV2O90Hz2Q
FTZlccpK1NHXOANmIzAqVeuD3nOYjDl3M3FQok8BhbXQwog0vWtU+qefEbgZ8E4q
HKCrDefWnKQ5e/odUgPSLG1hwYeiEK+9hp6zL9peoK8e3/RDpoc1ChBCTpKH+Dku
ctZ9WcyPYm1gAyL3pO75JT4OHsAjmBQER+7b2cB68USb6EIT3orN7XwTSox144Qw
mOpvcn5ILGWaRvYR/Ok5sQZ2UknioVfgfdFcAPxmsuCuWs3bK5Tt1Qfc84wHTYiX
ey0TZdKpf1w9/d/3TJpGPzIO+xNnIoppkBjkVfgSM8RjajHnCL7Gd5gFvBVoo1wa
HerE1LkXwe/NrlpvthGQHicOyPA34g1PW5eK568BInm/MYuxGAC8uB0nRid/PjSB
D7Z4HgdwE3d9G07X22wWx4cBaz1JlvX72htIZNQlkpyXaudnZE0rFsLceimodi7z
HpBP2xmWKcr1VMaKy1cGiFoySK4p4s4nvxGlJ09G+Xa4VGn78QGQLShfiEgcfkDi
x6EUXzFH8YI9QoNwTnh1u1RwUcVmnxq6B96TFU3ji0lQ0iZlB+ao6vemUdkoVlZb
QO9ptfggx97R5IsMPhh2EWikSkw0XceFsfJ6K6ohYFiua+dX7spGjtxhsTrIGAXT
208AqTl/fVDm2MB4+nUE6v6BRQ/0K7N8p9cXoRLfZsZjQLmTvinK7NTZQZGQocp0
lcsgMLfhSsUfK79KSy7TEtFxHN1gw5mZz5Xh37uRn+YXFrW3yrvAkz8D1ftaf/2Z
FQokAU8ZELyTlm8GQnRo9IWOErDIxBKBY8jZIgu3786iQOp8kZXKXupO7GRK2/kQ
JneX6sIGmvtPb+XIk1UF7ahohcHQH+HdfKEmIeQN5TiqZAsnycj264fvCsjc2/Q3
RsiPOfrPC7D3pwxhpknBG8hLWD+fX247xAPCLzmDVz8g9RZm2AUC3DiQAaSTe+8V
zxFBQUfVYzYJ1IL4hW3HUQuoMXrGZe4qmA9TqzXXIhtMX7OTnkdo3t0CwVni7+G0
Y6W7BtRlKIX+qdyD/DlRPy+P+h7G7+gM/VPz9TclM6qZsFTKNXdQxAvP7u9U/buo
Lt6nAZ0rwLfka13qBdPjo7NgIhJMBDtBPOeXgMn28/iap1B3zwqXcy7fIu5IHUov
DO1/20ZMyEpnYHBW/gCfNUX0B/I8xy1OC8eI6PQY/A23Vk6mViYlkhXCVmOFq8Mt
Or1TDeOnDWoAQoIDDwAr93WM1hv1CDDH8MfSxWLtyKXcsDf+MllbE1DyAWnuaEup
jwjor/th2gdo4P1S4CY2x/m3VLFBJvidTKBw7TleyWhahMcyx3m/idY3TGvRfZPb
wBoAm4lkcrrJHXCaFe0tCJQpChgE+7biEZQgDmkRfCG/JMsbTR5/mJHrhYyf3vxh
riZCY69TX3MpqvVm6yUq/9Kqpa4o7FXOTh+UniKN5N5lb2OvviWCu1siHZTivU63
6uXBtOIW8tBlL/6P1xOnZ9/ShBTI8qmRxFTrHqipzMxrdugTMfGQpokHwcPCK2tw
HU/B8q6JUTFEXcB5D8FTCV6V+h6dorZ4P+Y6tLSndsr9COSNm8P1IGMYkz70/Lo1
cOyKQO9ZPo2/dPuiD8s1iwv8EpTRKqxBvyOqbbMCIqjySSK5ACe7NIGe1NnOdycV
SdZcWfM9G4mS+McmUX2olaGTRdRFmBxVrwt+WJaFR/QF/z7LwyOLveEjaCb1GThQ
UhTFr/DjEnTGschipQLSu+LMtn63M4OKWUtZq5VYzRwKLdW+M4HcB0/GfRKBT+3N
0JygXuaz0KnN2T7ou1ZvjxcCVGjYph0jQvqsB1l1GrUI+Rb9GFcqfxsrNimAsWNc
NBjfQvbf1Zw+W/TNHuSJQXBseHpmU1DAYg7220vEiu3ikIuWeMSaHzP7S7Rk7Tyy
ugVbW978fmS3qubjHArH/BPfE5o7167LKPxi7E9vglVArpBizwL6cMHVCmH6FMqw
iLyFhS+ZO0j1L1LsndvuqIEQ8x5067sdGl035xL3BDKqZThQ6ThhounfRG51/0vi
/jYwphVMWcr8Sui1EX7I5Rk4PiyGv7NUvICBuvTwbpDfrSdfsStSf1LMKUxWcWBe
NN7+nwKtuMiahUGToIgy0+xMJiobn4TqmtOKSM/JFDN5uoOwgFaS5vH81PVl+7FW
l2H1rwOMUvy9/w4TdaZuPrzwy76qkiJ0+5qWnFc4xhjcgaSYYRiJRgKLoXCBOlT9
v5tx3ztkzYoBp4giPDA1WsDIt2II27eCLAviXfkthW1+WXKUKasBMRPzb+gHcVpo
O/pgnbYRGiIx/gkokYQYkNe3ZLkbzk2sRwhfsECZQ4lNkvWm/tq4QKS9R1zN5hZ/
kyhIsiw12RmDiNjAQ54vdU5rrypwHpwQddAXeq/94jOVP4k2kqCuXmWQyf/NKDnu
CylRjokLk8bhjWrznJH5wG0pgpoj7ScyU1YWT+mtQHT/2s6og1QZ0AGUt7IA0pxV
d2QrhH69U9ae7JkBCqk5ozCVrjzu6rGXD21uohfEXh+QVqRbg0jyxey37v8NJW3Z
aOkLP/cDp2mjjPo3m+Z9xw0BexbXapNWRjrbrgKRBOViP2tzrEZWxQZLcXoYo4TD
BP/qXvyN+fzfYVongs27GZRIJfdX35nFV6PjQPTYXsPXUZlcmNXxb/TD8apVByor
2Cm+K5uyAi3NNWahIY8v/tes6tTEPTkIjvcc8Ps2kVbpFe533VkYKkNDQqTZQFoh
wiyxeibsMMveGJqwhX6gzrIlqO8PHf3xR9LbN0m23rpnmC0zIbzV6weOD3F4UHOv
OsS2TuZu77SRvwjcRgxQJLNkHmxdYwkBtRZonsItdGpkfwwEB5FPh/dvZxlkgbuI
ynnUu8IeZAtLHN6a/5A2nmzgX41sDSe/gE1vWxcMlgJZ4dnIeJFfRSiJix2ZcDZm
adSerx7DsSFJmAZj4achrycREnLAeNtzydvzcAKQcMh63k1kcmXApHEftOXo4Q5E
EKwtXivJSIvgbV5gg/aK428yYUKPYRJPD54fg4Nvn5G7s7zCH/8xllS8W/q2gjS7
hMz++fXA42Fkf/eq/Eg0RJ/3KrVlXrTW5cSdclkptgPKAMalsRAj7Ot69WI5b4/j
lqXpf6jzjVKQFixvhJ84FVdpZTWUMZzl59tjVMt3cuWy4U60JagmSH/JAW8mFAyo
574jwYoRtcsBItuqUjpSqyMYImBYM5ZXlobCclRv4Rjlzx0nz7AgLid1uHQKmX9w
aho58DhTwotO5v6qvL/3dJgtiLQB52KACayXVplLnnRO2/rrTyHJAykAF0Ar2Luy
QKNStSeSRJzKqGbM0+fLnoqM9vFjtLKWLbKBgbu4f+2Wvy+MQotZvb/cMIAVcmQR
h1D5nq2Vm3DAYnuywQo6vNw0AdQbCyFP2EaxKyWjfDLyrtwDBSjedAM4wgrfHuQg
++XLd4hOO0N2ZWlCOF1XuS2ZiM+K9WE1+IgmZCIYXkv+dgjhd5ePz4wBPpMS2czx
OY8zjNVyf8+xfBO4w/FKWqqieSZZE1fSyYdWPRd4TOFuv6rU3tInKIm3uiUIb/Kq
tZ8r3NlUIsuQYwPVEhU8mO9EmnbS+PINdJbw+KELzWPkZ/iOC+MV9LF28aGzJxS1
+kjbZKmBwg0Wwy0HBICVYPw02N10dTC7J/n1laDMzr+aMhP7UmXnVjnpiG0KjaYV
ze16UG8b7agnEbtv25H2EttFhsS4Vxf9BPUxm786qtJmOTfVojedWZdQjKT+2Ubq
lXih1KxtX5+hYCxy1UTCG2bHodrFIu8qkfh+YE7XylmE31queZzOicijKWuL+YOd
Rn/EARPW3JW9LeKwAST87YrGJsrGROZ7G30wpk3zYTnBvuQUx/zjXBgHmcbGwh1z
CSBQIg7WpWKJLczyYQcD2KjOrJgYsnKLBauVFpp5p4Wex/fIVcx2HN6xZSGuLdH8
4avJxVcZqyLgaO6OWXos9VNjL2JxqYRljfklQdShn0p/m7yv9BMn+LVrrpFyA3XY
U6w347xUXq0DIlXeq4m5si+RsI4dm1OBfc602bHhA8bgmqPhZPj0mwUSRk3aw7sQ
WGUXZMrOyM3pMNH37j8mND6cfx2c4WymH1BghhmAicEst3y7g8OQik4vicpdCnp6
CWlgUAwRU3Zs/hho7gw27lVV5qPdjQAeQBFTJihuY5o=
--pragma protect end_data_block
--pragma protect digest_block
D5NJVBgLd2tHFR9GYE2miostHxw=
--pragma protect end_digest_block
--pragma protect end_protected
