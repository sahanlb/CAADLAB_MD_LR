-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PREFp6dG7dJTsehl3iJ96KOi+yfnCyPYPzSoaMzpkrHzfEhbG4pxaaCJtpDefewSLXP6QHaKwROC
OcDipa3VvDz9Il5cpS+bSrWrpVssVXQRqERx/UtBtDjeXMUKMAze5ms2TCAW/GshDnQrZxWDr5cQ
jK5sUsCGHn32bkt/WQdSDaxvU619j2hTnqOUpoiVEMxU5ns/84FOiOsjVHVTh+3M/n8g/EYBFwbi
dnSsg0jD0an7LFESpPK0tXWKxJOynwxvQvX5Xd4ZWeyT/mioV9BYAaCq/+B1jyiKI3p0l2fYp1lf
9tzHOr6onGH/CNK03LHAnkQwYh1bJYuy7tYQDg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5392)
`protect data_block
J5ifD/dNIERqPJa+L2EIBy1AvhTkwcI0xLx7wh2JngJT2vCxiIltQ6Ng+ntHSoG4o3MP4935zGG1
5Kae3YFRmXApXDdujC0M1HXgJ1YXhiVWR+gefxwB+hhSRLnDbfPn9ev8mwr3LPZqySq7ILZjRhkW
o4glur5sFSDUyJtUA98hYtGzAMsb1JAX1TFhxcPiCGsZmRKuO7/60+t9beHl4CSH6IzWTd4jaFKH
/cv6vfmFw7YwW/Gs0LXLuiMfKOZWJLH6hyBNC7Lksz1kC5vh93c2WoVfgzbbJlOAwIF5x230Je0I
bPu0wQw2HoUoRfMoxR7kpcyfd7uLlIkWl7rS0gSs1y1N4iAzmNz3XNRBMf1GRTLeefb6uMhyTgTF
im142QHgkXr+qFCgypofRgbMvDHiwER9k4kJA3VN3fZ27s+IC8PUIUvZ8q/M5YRjPy9Mfxd6azMR
Qb1yi4pR9GSTAJDv2Pgb5k0EEG/ozIV83TKQJQsUeoMSsTYysZkhItLsO0ES7ssDg1VTvwDKPPiX
TtDOs2eEVeIt7eoG63PZbOCUTB3+6529MeiwUhk3BeCofHYZ33HraZt0SaJ3tfQcDrGYTCMWQkaS
/Gk32oPE/TAabkcgoHVocNfM9Un5awZPclzLh3YU+2teXlBpKS/Z9POOZ6p1jeeBHlgMDwCcWRSE
GeutEPBTnz85mz8fwwLIkmCY4AIWfi2hl3eItu3Iec+DJVCCEuqjyeCHm+7568EEUnhrnuy1TRxg
gOusOUxfZZZ94Im0ZuModO0Qgea2wAPRLhxFSW0fZ5/oHWmTWZBJtNeoTju7up7fSH2xZC0p8xRl
eGVktb+59j1DC5joGgo2RpzTGAaKHRHXT84ayhS548bfSMOYS/jGjHZKPF09Q/e1NFsyIYXHyCve
3gxuKOqRtr43R6EPrq7/Z97fOnP6z37mtezqQrCmT5Jb7YyO2KzZ7BC+OzjunqpHJVuVrWi9b31t
wea5ktC6yrdk8GBRF+2DwgIBJ1IDFrq5bvkrVCd8HsQ/ewQR2vQFpudQSeuTbLmII7FhhQlf0ATP
chKhs9M8jo+gODJHZ3muKFFLiZ0Mgsvmn0Ibvux6nc55DBVX7JAG4N7AVKuG5pn7WJzLP1bsvWfF
2e0Ryojv0L9XULPtZnBXqntTdIUB28rrIEG/yB51HEsEB0ea3m54hzkgk6Wvee7bjTd3vtGDbxQw
8NJyixhUJV+PP5URMA9noGuVNaAUOJ/pW8R7j3H7st5L68ltEjG+l7mwLyZs8dLlrqiNw2RaTjrC
nGgS4sslboDC+VoWlCmCXCr7Hsu2A9Yh6zOzIeJi8rYDEg9Y+b9s/xZpcZcsVdG7DWiXZeJsMxu+
q6Dbt2LUjc7ChOzucElkFlW/SnmGbj4307gjVqzmgMIhJ1D50aiD/ssbwHiT9ThlNMdtjl8KIItA
7/0upKJQ3J9xlIZGOb2YQRVZA8DdLvPCANO9dlu4+MyTgm3enew5YVOg5prDxLLrdVrAAr5zyYOU
m8SO326LZ4hXeJkTTjkoa4Y3315wdjVgm7o0ZpeQWwxYOCvEhF37Q6jmqclk4lq87ZUhQTLB0Ws1
9GVl3yEu0Qz0KU8H1mCuaralRdTtILD3Y4vlpi9QHXuDCJ6Inud2hYRFaKkvMeqBHyn64qU5JOUg
ZDckWv5VJrVOTXCyVh5Rk9mFRmeJpcFvwFOOfdRQH6EpsMhfKRGqHFcXMJWXirXNs51pCDhVbSHQ
wX5twvnV315qYVZGnhVcXYm5okUz1afC7KGUxnkyScCYMUYddkQCFxzGlHBxqd8bC1s418hQAWqS
UTGAg3Rmcxtp8KUmGyNWjHYL6336hL4GzzVSO/x+h66DI46RA6rSlWUcNE89SqkO9i33CUq6ASH2
0fGMgt5+0L/dIjbPe34HoW1fRPe05A59S5LZtJJ4jLQvRxFlCtW7Bho11g+I0maQV7ti51hhvlLp
5man114JKEr8djzHROwQ0Tf4lk4VNpP1vgyozB1ek3kcGXo+wvQP0pUgRa0lYs53xcxmqzENAhv8
ZPINoMv3GUY3SKZVBgfaFxS9gkr8rZetHMYbKwcH0uhwJpwjXYbYXexmHsTfJrGdS24NnSgDe2y4
cN6wUmTA+degi1+Us2WIpb4LMKB+wUzYCcWoikktHQQjWm7dVdkivaUgFvr2VdswrgqX2Rc6UooO
UW9zP9cihMf3OwATbdnF2BnG5p9jGwSUrmC3+I0SU+FkGtX4TSjqILMblug3plDWkvT3o5qP8nwo
ln+LRdM2pIKUF+hYdC7ddMxgwdlU93u/npVCnrCOcQzs8sk08DaJ+9AVTELcjZUdwYfKgCCLgizF
jiHa7y1oiLCGafsipyREf4RPysuIqpBTY9ELpLoaWe0w9b8mvhUJHtJeyI1Lz+UD6I57Wi88NKvN
MawiAcjC6+yPLgdluHC4R8hxJ443KGFzywByegdARKxqC/DEilxUbBfTYr8m9XL6/S2jVBR3V7Ki
CfYAJ/Q074ue51T7Ijw6hEm+8VryPtMx9mMXRugEPo9d7SFKxQnVO6IJxy8uBGEI76+BLk4kiAhV
vjvP2vrLTifMl/farFNV0vXY0cqVwL0GLxnk6216X5esYeVffOpdUh/0lemfHrnncfhhDHFDKAxJ
FUV315adDygAmAtmt5/crjJf4+8mJEihfXLxYfLIOG+R8Odd9L76yy67aIxXQzMlZEsaE931huBH
SwINMwusQjf2pzOZVQnTURUXMK6vpVYdGtlkeKAUm6xt3V9SL0sCFD9ohVau1veEUFVkmRM4c1Bs
oj0xP1VRqAYV1OQcJhN/w7V04b0Lc6b8fyezQOc6t9QAaug4tnq1YFqxXJXgNv3g+d3VjrP1qDSy
cJCt+24g3Lwn/0dFrn4oTrM1oFu4WwfPxZacTRs5Cnh3BUr5LXSJhE2xOFhVfMlnzsNjlhH7F1TJ
r+0HoaHs63Y4e7TZlY4o0mPKf2uyeKyulSNqSzNFx0hUw8uEkPF0m6yyKOpG0ITpXfD9drezF2+M
iPSBvuenOqqabjzcDr4+LNtsBJ48oSbomAGg1aYEpLxSiUPMa5PEGKt5rhTOrdwT5l2M7bushJ0v
uvRbxMI0nI9RfuBIjjqwfLDqRP3IWjokY4xe3YS0fyqmI1xmWe2K1wt5joOa41dvekSgWhXqqfx0
X0iGRi3dN2q+1Gfki+yumQunbmjnjWQE3YKvni+AmK09LTe/CCSFvNmzMPiLA+JkbWj6gJbt3cnt
1BAyayjL54Zd3ryh84jbzLys4blUownfBREH5kep90+ydYXYFkitPj6ym7xryXVWEbXZza1iH8h0
9lzED1VxezOZ6to+eDLZzap2n1b39lDLKbGg0tDs8KEe3S5nCYW+S93jOPllIAdyDtnXp5Fq932z
leRxQk8yXIxqOBqbukOhqiYrcs8kJl7ipoDprCDhROiuMjVUOgkcIJwyajrdCqTPqtGml/Hostfu
RItFEFaP7o+qJ87elwYojIKGqhpb5S7maI1yaYJBzKqZHDAQ0PEAptAVpsSg2jC+uYxYlDPZvbgv
UDPnAJVcpj18XYpdzS3Fd/CBXFamFnut22ADlzt2w+MkAWzO+WTGC3Nfbgj1p7GfLEhUSVr4O3RH
2JA2aTd/ERF2X/J47FVjcjKZ9aKO8dYhHjr229rehYx8Asx+qQeIRnM3vbdsryuaVMxP5L80Qdud
AZ7rXFPD8ElnU9H+77Tp+z2OzPszxQ1UoM2+2pkGp3MfRgW4Kbqk0Ib0IdpuobS2aOQe2lLZXLAD
ZcmkTjn5bIRc+FFMNtSmp1hzq79j0EPlPFRnRmbXn/cfFg7/non/zLhxVW8UEN/4jWB3ngQMu4qc
x1W/af3tZjl3YAHGyMiDc5MzjtvTyEFO8+10+P2agSDMwiulCNs91sv52qofYhHa60chpuoPq0kj
Clg9PkDKXqBPefZjJycM3pjYUgbKeiVB4V9Qe1+CoU9uvV51h6hAy4ChZUDvSyhx6/lbNNwpexIe
BzgswV7QBvQniAhpQUbc4+NWfyMqnfYeP/Itq9b/3evhXjk71J5Ffxxz7yf21OieMbyWHaZWAqOW
3QUBJZ96bbvZuf/C64FvDemG5tbjM33keTyOZBdFaJkh30kEVl3iv/wM/X/r8/vVRqW6JZ3jDvWx
aKoHhDsXlQjrnEPF9Gs1T5hbwueABixUI/TlnbQwN9ZAZdG/uKUYe3KIWD8cXwLmP3p7bG/wyilg
nihBnbiREJIsqiIqM+PVpEwQHbAUSSbjWl5uMZyyPBNSGY6qR7SgwrdKW8mwXGywcrGIB+Xi3YDr
YJuZxwOotf52D5nxLCLknYl4LnDH4CcSE6Yu8pbPO2cw203YJECPZKnEngoxIlBfWFi95txGRdQR
t8QUvip287sK3YqKwFEdh+FAuEG8G9Y5wND10w4JvKYnwBHYV1Y9svFlPeoRcWYkLqE0OIfXTlae
EFZDtjVHAW/A7UdDY7Q9FQVmQHhmo3TyY4ESYnj8Sgb5RgJVuMGMwdwIe5t7vJFzJ1kEk8Ueu3nr
wMknlE7EGTOSrMSmSfMOeDk+WezjLvB5MR4MLg53jfjNigVLjXEI3C2exUaV46GbO9TSElOn1Hdz
m8gnBSH+kgbXOglxcVuSJYviLGyK7abUQUBcfkUKtVSQwLK+MeT1aQfro1uyzbVviRbBaJgpZKgD
N49BFOA4Gb2VW1LF4uL2yogboDPK/pmfK1fESXOfU9PXDGPcBVnaxMZQdeY/X0dkigpg5Qq7qNPM
DQvnQGw6qkjzSyUbya0CxIz7j581NffOtp6KqItpLoY5AFRtlEKQMJ1ncLLx337OpeLExPd/o0rf
REN7/SsREGy/ALjICMnp54VIBR7LguOdOh89oCrNcPX6BuQrxiXYsDv75yS78ElNpD0R5Bn3LqRJ
8njNTApyefENBy2G7ree4ATYsfySiP8t7zeG1NHi//v2VLV/jjQ8smaa5Mgoyxa8nopXL1mXahhZ
lOPNFotUPdAk+58V4M/A/hMY0/syw3nelfZMSfJgu9staMzyZMtDlvHKI4HrRDi1mcstnX3B/Evj
bI/xCd9QPfxJeaeL32qx9iGhMiHHeSZc4NrUSx23BBJamuZykdqve3+5h3c734YUkcIUwFu6FkTp
nY/I/uYIjXFNwMoQ2ElhH+3EwM4e/qnBdy9Qsbzdx6Na8K4xjJ2GmqrecDLiTzUgqpxWop9Hrt+/
8rO6KGEXHowFGFSpfzuNhUV5XCdzqoxqNWuOQH87qLDKccRe5ZHRzVB1LEwgGhbwGPg0u/pH5es/
B5/iPIhUAKyv5WxcUhtdt8iBgHlWYRaQQsJMRaE/6O/LYBsgFIxyaUJQ7L5R0zjqWBoANsBW4I2w
BLaMFyrdKV6shQY5mtPwRBGQ7sV5YDq9fG8Zd0f97rIC38tLnoG4j2NxmGyGyuxLr3+tTGkPAiA4
t1SM1BByd/KXWFHXCBlS2OZ2V0IgZ+nQP7eEI3znZw/6VAaGjMyQbeCX9JURr13PNhU5NSANinwg
xXWgDNhOQ4DSsszw74TL/xOCYeEmGF7NZ/s1JM/IQ/8oQ0dpEIbly1fpXbYi6ZeEzNvaNEwtz5qg
oXItYL9UW5ErdKNuvP0k4C3PvpRHvDQGOCkZ1VXCGcH4ITQJNvgyTXaqWlspDHJNew+htJqj/YvQ
iSJgo/21CEeFwJlgoBVrrNy3YWimPM8FwYL7KTSiYM5r1mSTSQpvVKyicvLWHyIqUwZmYJC5UKdJ
0qElI35cAyQTKCd/ccB/QCvTipwaUt6xGkkWOdUKWeqZUSCgOUXRqdZsdwlKZCah5swQkohjWuXg
qDBJ6L0HFbz1q/lymclhuIGQrceJWQB1U4whfFRamFw7DVpMtysi7dQoejyKEq4oblfeYe7u1oPv
5j6SDsmrptw0wi7his4k977ycwA7pzqKrx6E475xyGB/43f/6VDCdtazSYiCbtYUxwmmvsrcmw5X
fddmbxGCODdHJLYzYVo+yoe6FutnHc0WjENge2VMQVrtJ5Awtfx3Otu4sAGPJmjtq1cjuEGk+xyf
QQdcTAMe0rKoj+MDzMwB7qiMnTxXUKOMJVeoUmMmQ+jeDEJGbzTYwDqIr0nsR1o9v4bWkCU3qrjm
dgWSyV44ZAoJdpbt+AYuXR5HXxVhiJ2CuidxFpXxGt4BLFDvzuzu8LkfkZxVPRFWUadT68otksYr
JWeeV48gL4EjtiPTXt0nhxotcX4HJUJk8LqEpBenEOdft9sCoaGCh13VCmftULiBPrMrJTMYu1zd
vp+1Wh0WqyxHverVig/q4UTe6cDkMJoWtTXVB1yVbYSW+18Ey1BDg/Ispcw9Pk0GfDpPbBer93Nf
7xEFREnYdXWV0bQnxGW11vWaxb4NXcSvP2vvZcfEbjia4ouSx5FY/EOC31pBLNoUF1lXNuTlysZw
vTvY88XIiuyCcfR2NIxu6PV0NZoyYakwd8Z3OEyWo8w6NcTTjmtaXhLjVIqC0qkqQXFAuhHh0I+r
Jxf6AX3rRGVLg3jMxvnoKAYsEe1g7xvL3qzNiNIMG6zO3+dNZiwrP/kqL59Q8u0nI1QvHGC3a0Mj
Y3QbdPlI52XLpT9+YOMjPlXI+O5POZX8csxF+Nlsbdufy9c4PkmtvgxUtyGOibHPSIFewhSNzbF/
41blcSI9EpuHaitp9/nmBt8WNIRE446J1j7gx0te+4mOR0g1EJb84hrNc2DfrZJyx/nWq1eIWp5t
l4oH09tTKtn+x4FBmQguZsxPa85h0LYnf3INZ6irn/uMBpOKJW9B1M0Kul2bSQ1ddNUQrXrLXu6p
ROgNFmWd0a83tnD9cxFg6ASwlgohZdm2EE+raisJ1b4S9O8VgWDrj/YdkZSFca62QEZc2rWsU7dd
qgHvlFL31A712d8InF0vaoQILvY3YZtxd6n0pbdPAQITF5mUEcuf64cTaAUgONtNTW/HGdO/xB//
NHHY8VfdxhFCrf/M6IILO/SP/+0Fsbva0qZXUSetHeSzkqkKS7xTbEivHDPZsAu9y2g/nG08vTkm
wj8Qpqcwe9XRMy3fbr+d8A+CfsHdzAo74Y8j8/DP+FM5QlcQlzwkYFu8JXReQSChrUDfqc3hU5w8
t47xW/gir05MbQz1xxb75E81/Ki7T8hodCwcIcR6j5n9hQ==
`protect end_protected
