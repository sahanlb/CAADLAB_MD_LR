-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
zlwFqLcOjsn0kC/fZpiAmiX+SGtrzAsTJeCPmqaGaESujpCbhKvEEbklsGY5U0o6
Vr4biqzKcXGIklgdU4roZ3NtQt60KGg4LjHOxBH9twljryNNotbNUoKyNpRtQkje
kEH3SCDE7p/QpWLWcXY/hKjNv9+4ybIoc0Z+kQQozP/cJxStDDu8AQ==
--pragma protect end_key_block
--pragma protect digest_block
Ce/w1mEJ3s8HiYvzozlkeNkFneM=
--pragma protect end_digest_block
--pragma protect data_block
+wxakpPgd59ovjgxlS+F3k9TJdpYn2oikzUYST3J1M/28AssdAH5NvNR2pQLykqR
6o7UtRrMdsoL3HoMMWApUiey46JTZiAZJDH7DULAdW/wjPR9LLMNzDyTQGgF0bU8
l7HiZe11Zu8XveZNsWs6gLd8imgFq+7+yd53bI2xl/AKR60XDMLmZHl/8tTTKVeU
Y5oblhTjX6/7sXl9aMiaJDr5+BBpc5xvViQ24pg3F0S5F3ivn325O+h+khSCNbL5
gIseBCAxgSICyVrJYtsK59bWZbWU6uTCbMZuBq2zKq+3VhjtmJ9kYZ5huGxLr7zz
gLxwbsXJkUfynGbPkCF0TZPWUmZ2T+Icwtc1ejDm45i3vUtIUAh1YYlWxYMzmaaB
T7RwezWFVqiHNzdwuvGhiXBetuRUcHIz2qXG1JX/vQm+ewbgWVvXioH17u8txfok
HWEtahdTdqEc63js/avzoHj3mKIcXvLCKIQ1TKteqcZg2HhY7kTffscqUrVgci+E
pZYjU1HFrWQkWJS+l+kFQ3BqR3DSHeyPBiY8FlcChMJhxDZiUDSIVNVFinxbM9jv
qxgtR/2ujJ8a3KwMP1XgcQA/rpkwLeORTGnNEJuu12T11tF1VCCX5A8z8az2c+T2
B5qkDTTeFNipScRe/WomnuBO+irOnfDmTT3gbU56z6fFFPL7ceo63Nn6uimVzvgc
mHZWxKUevL/JsIBZ/cCD6NLgtj3s4FgARBn0uM/VpllAzIB4Ypy7qmFVFRfnyMJF
p2dy2G6sC2uX84QcjoIPDjx2iTU9iL02gprabWJJx1JVkcDI+N1cW/L/kc6xbzru
JVCJJbe/Tvd2O97y7HF17Qi57JAk6mEB3OekoqSjzJInWnWwxqK8gn+2hSaCbFZt
+k68rgnGk8cGStXFLKao04ox/iuT5C9P8ARPxQmdtvxxDL1V5cA9GL1VhB1pZjgJ
MDPbGBW8KosPeT8ugTQO5wdKAAdJtsbWsE9pSBhl3Adbbx2aYwuuw8DEiByMdSf2
bqb7u5tilyWVzVZ9xehJ2DEryexih/TUh/UEDWi8M/+U2EZEwmT0TjPAoml1HQ4c
xBW9CdHDFu0bzWH6WwgG6rV6n4YvdFT2OuEVOrBHISDWsn81oldStF+i2CKi1hRW
d/ifxsNqgB2++79mVY9Geb2uQui8+IauxtwbMocJFvoNGkFXXalewxvsFuawAaNy
ly2SPWG1mdaTqx2VnunR7TwZlajVbe4bK3TkOnsSfriSThQdK2DuuikzXwX3bhVO
oSMLCe+ygzB4HfK85m/MhGsAYuhSbeaPftsqsW4Ecy/bjpguHxHgJicSxV5P5dRb
9KckYQEspiNSqL/CBqPGN/nCF4uWEgm/OcTN192+5PL8W4C9oV96PHDp++A5NUdI
VyCnIhePKLhz1Nni8eDV9fe5nl7pr0cgEqFHrj0LxrvppBRAJ6+sfw8V/vH0k2V8
FI1E6s68U1J4FRChhse+8CywdNTczQRsToCqQwThGhxel6vqDwhI/L9i3zncWHji
72d5onF5fbayPRUopSPYuELNMHA8P//Jax10MT4UjeFLBCZ+31XuzvgnXLZnRymA
5TxN645XHmOywB7oZQztxs/7szuloipl2naguuOfZbduFcPBJqeU1TcTZ6AOVhW2
Kq2kkL/wzECfylWcPb9mgsuaZdTCIPh4DecQUpxXHEEXHfFRQ/YyzCzdd4QfQj6B
vQVV2Tf8quVsOUAOvQFh5q10L0X1tB9/gS8GIsYQC0PmKsCazy0aGATNCzLUk+Zk
X3bJyfKgaMFCOl9Kkdu45972shUie5Xdea/7r8SedqRJWf07zw8wQEsINk6m0MZB
WMPLOPT/dkSKiLJC4F8K8sCyS6WDtBuiooRKn5ZbaAP+kyTaydAoyhQMbvw+RadK
c3IGWpRKBCO3v884m1OeHZIuiiEfIttGlqQIoFIWJ9wnIAY1xG3aNwObNbpmVc+r
zyvontcIrcmDSDIpW+OyUdcxmYTZ8PgLGvjRIkzCt6aj2eeYkXcIxmmhIjBcPIV+
8YmvWhIG3d8o0/fSyAebhm0kpxZBQcvbZg55ospaO3eGpZfs1IY80B4KRVHkgpCM
zQCCiWYzIQbSYvNuLXlkPvvc2M3nnmSpBDFW3v8UXoQcBSBj+hoO76YKenDQQmVB
v0eseLGEuEd+NcQKpBOAXaQyV2SobleTMzwM638KVVhdLenY+zLXFNaqBYIoBVXh
40yhqlWxD4Ji6CqrJpZgQJuO9NelaE2VIQ8L/fpnEpj4M6XZR+6+bQihTEFzzKXF
rnAxGU6Sjk2moi5roQSP49WIqVojyVjwv/qOnIDwnUPFjL4IYw8d7H1jeM6RZY2X
EHrsLhVONUzqA2vQTHh6HcWwotin42+gtooMxvMwcWD7af8w2f3DUyRXLKyzMt9n
PN2fhn2bDPYZhPc1dyJzXipTafWa348fDnayNXzyhrlopjAPyD4gqUboO02zGTE4
4pPV5TFVyeMNTpeGlg58BLK4F3hUYc5PPyAnWKCEENHgy6HA0tmQLXCjlvY0rwF5
OcSmRVNvzH5dosiwoNkXpkdAGHyLGzDnOxrrQq8ycsWdenEMvJ82YXOibnL4Uj5w
mNiWAQa13tZaj/4EGCcltH6HU8vHPHvNqrr52oAAHWLqPPXnnAneZbY2KatzcnMw
uujLj18IGwKFuvO9RwsHqDnHvn1/f3KVWfpwkunOYCYcQYbAxP4DcWbDrOf8I7rl
FBp3CsNtWl2QIxGGP3K71wMefFt2nB4i7L52eEsCWWyr6ux276IMF6nfRWWVlbdy
CJrpmCZ2Y8lRDN9yqCcqn0/VBvKdcdaP3hsbM6wFv3Ml4lhvmVukVdlYIh6kO7v4
Mjp1SEQtRFj5MpQe/brH0QRcHXY7t0szKOrPuRDXYTCXPx2SrvlrLF471Xx7bMkm
KUVRHIGPiK4hs5AdHrBsUKCSorDNT4QtNVOLLKBdIeO4U00FZt6uSWB/PypvSI0Y
lKVilh+0dIGcTGcm+VoBU/u9m6zOeOhDLH8pD9Yzw6NbZWsjvhtw6oPhNAR5ceAW
0m0QjxPGTlY3dJKZP6SZmOwy3nEVWhRLjnZ9ZYwKFm6aAibTtlWRWPnpOaGjuh65
tHLWHb6xCbzfOu3HjmTP+NNh3QqA0TYOMMQ0M4AgfVu8KFUw3raqcayunwNww3+S
9fFV6FuR7VRmTmrPMT8AVTIx8jDN+0u4ReEpLg10R/+0ylbKzT+KqSk5ShzAIDGc
NCQVNsx9/QGg1bAzaHfrH270mOKRmR7ey2aOYHEB9JdRDxmNt/eR/wuuKIEZLydF
QlLWD625fBkjlY/3lquXP1ubnlo5anvghsC9cipppBQZwCTQYF1fLDWRFrcBH1MH
GSTjHFb24gOQ56h1u5SKikKNZZO/y6Vd1A4mQOaUZvidCnLQ0P3OUpDt2KLyWtSK
HYv+iVurDp8QR23qFgjA6pswOHJKbTVT97iNSkV8GpY/hd990mhwlPeSroxJAHYD
k9PzrALz6Bx6y+KgNJQK0ljwa6OVBy6pZDgiwhoQ+hdE7JiNZv6Vcl+6ix2P2hMW
q4Q7HXwwAeMGblDBSxicBbb5mXyvf/Di6jRCLHBd2Pxyuc9bg+wQVSbjse9wSNpZ
7HklUhfHOAiVWq/lIxmpGIsEUfJu8312LVLlwMP2BP1u69iAkmcELYB1w8w1x6zO
dhSWPtTpYTamoCl8AgPjAatX3WaiijE5EcMIYJa+uoSv7Mkhf7mzNBZxnDJtOtAE
J8hx0GIlBGM/Vc8+i/CePOLUdJH7I99m1ysNugAQTJ85ajUWXPkF8NAhj5HnfDWK
Yuk6wBcN5Q8lpGKCOp8o/TtNS3ZuDtpL7UTqO92JQY7s2RTIppEuK/QsEbM2F7ta
JmWGy9mgrH0hpWiVTE7Izcl201OIm8Xiw6StUbsZQUlDQnoQsqphaGIUZrlaAqjT
5KkOZWW0UdAxgK9SCpnAngmUiNokT/8/aY1RDI2wE/UZhUtogSUq6/+oP9tnZYJR
nNSxoGtZBVm+I0P4w5gU6FKcv1ISEQYvBlN4t+CL4468mPMb3fOw7N0aemwwCZ0R
WAZiSvbXioCw226wUQMqmDJ3OiO45yykFc7CitLa1YkQgjLKkUuAbHriRVJ333aH
/uRhwdhLSWKEDAYtIJvLoO3ylweyavRK347MY0ScNEe8n7qKJ7uCdAikaterPOZy
41h3ff1j56AHBppXrWBkoh5BavBf4uOfWEdUjjIgHMFiHtEkMcNk7s7Dp/cGhS71
SkAzzHo+Df0QOf3ZdUSCEf6WwAkS0puuvR+t6OLvc5WISZTn2RMVndbBujoeQZMh
N6sZd3btneoK3/S6J/nV4aMuGRciRqoNCiS/kPbnFxsVw28CwMj7lMVXqU+jDx7g
vqFPhrLxlPGAkCn1VqfCoR0ZY5H1bLOMBYyulNzJxl2jIstz3e5vdzmF6Nazm6mo
GN0s5iXmQZZt8fxYSmviGqbsro1L+aNp69o54gSrCnTEydnxSYX6Hew285kvOkml
3MEdjHeA2mcgUDMk/gy0+wGf08DaLaEzDY6WsepQk/u2zmOkmQo1YEFo+TUA7sDg
vBdswfDh5l4VfE81zoJ72wwVYRucOP1IBOow3E48rdwcU/el/3eKb5FQQ02/BTwk
qwspUVW4m78FIo2sT5ddhyrW90Qp7CTcCu7vvPn8/kjguygl8gsutC8MUjQJmzQf
KBqFUgYD/4BF58DGl3Kis0j1VlkR10n0sRqQnWCk8vHmWAmfi8xh2HQSYcISHFVq
wlXKzLzRGhK0hggHRp4YRer4OExlrhhnfduZ8jWykWi/MLtalUYYz+0LTqbjsg4l
KL+m0jKtLCNwGDm4UE4Hy9A/7UgPIVY04uiIwen7qBxzMtza9C1NCrsw+iq+LG/6
w7Tyb3743oEoVPARCV4WoH0NgiiUEjF7wuxBY2oOvvJKQ8q8aHG5mr3bmNTf2o0K
Zic9GhlrMoAcTvHXLhgpLBdso/6vnc0hFT1+Sa6HbGqFCJFeqNw6tfUIcxkbu5GM
lXliMmTv3s6qsOADBXSYIBCIOqT39mGrttOIw2V6VcuLBV/f4kTM+rvj7H/kDMjb
H2rr+Rl7Khc4V+sRM88JYlCMnZRaUTgiBrcEZhgFVxY/mo4hRYnr9TL8RKyhPvHm
fSSBUqWBP67sXJBc4NZC0IgCVGRZDZEHEj30yhKcTpzJBZ7kOj7cGUpYH7iYhWvo
0ZjCQSgzCtsD1yJMF18NR6fh7m+k1aoO+Sj0Bh2dAXYfeq6ZSGdRtUYoLNah75Nk
iaqPViinz5Wi/v78kb7ve5+0DLLeR2X6j5xWiylk3iXQQgMH/xMT7HoKxeDnAEvS
OZDfe7+aFIzpyoAhshvjBeAe3URG+gEZuPRqpFmZ6Yrrb2SNaGiUoea3h9lIxJx4
jYawo8+UQZ5dhThwwop3PDMoT9owfsT5ToPPOKddNqEXE+bgSw81J3Nbpll9q30W
Tr+eZGWcq1zuQtpiotP+GtiSnk6Cl7sh9+LQ0YoEBggkByJbz+vjohjj/gOMVv/1
N/RnIPtkwqFdMuxlIlkeKrLIBWxwuskq6vgMJ8V6LDEzMPJ0yx2pxmfpHwgU6goX
XoRbcQw+ybEoyl2OaI0VVKO2qFOC2VLVnIhdc3A/fZ5nN8QvwdXqSV8D5uIDWqwJ
nBBcjhsL6NCu9/vboDMGqNeSuW8byEr63ElLecSRiWV2ThLfCLTcQbXbFUypC4rg
qBvKTipkL+nTJni7t3TqJeJ3qmA4rQBbmcynyZYWOF7p0InHAFgSN/At8VHM+Xn2
BQSBtcxXMw5Nhd4BBzCQfAm3kafFBOCTXXNkR6EJtaFAeQKS1L+M91mYsKLODYti
xXAQ7NQW+/ju3GUDsoOc8k7dnRh1QVWPG5yPzyX9iStZNBA7Z6znez9f17rXM9nM
1nPcj+3bqRKtz6Y8wbjkqfsjoE7+dds5s97sF/af3V+hPlx3X+EVZ4ovHy8phlsx
yxA1JaIW05OBArE6mnjbYGyhLuZVbfH3kQV4OFFaXWBg77N+qZF8RPmSDcTU4uzR
5DP36b8hYAQl+oll/5NhGOES7diYSqDDJh8BFrsh20FTYx6dBiABYJ1hQZjyLLyE
7srJee+SgxbNDvVw1OttlP/FliOc/6T16b9FjFW6tvtiUmZvRXe/CQ2H03uytQUU
VqibyFmK1pa4yCNS35aw2L5/d2xW41qKxUl5Y5t9SZaqObXIhtY7kj9oZOL9lObf
1YOj8c2Igr0egZbIEsYOQjpYAOb9pg6vKs6Dwuy4Yu0Ljn+ocukSUysYSNvp78cD
RBg8vii8zg7BC+U3uQ0w7j6KmLVk0W8rR8zMcgHY9+rbCaR61C5nromxcJDuSSCv
BlP6j8Hrv1LmuMQEA8t8KsPoV1/newC1BO+U1USSKn/uXSEmEtIMKVaih1V+c363
IHPgZdipa1g87yrJh23AILX1XkUdK0s2PBo151Y9Y+apUNATFzpympaZnk6MOWid
XlETzogYokS7t1NpTJ8oGi2lxHqBHdD+xs+YQWAci+I5Z1L78gzX+E+Cm8FRope1
fUjIsPNP9Mhr+8FpDIjRgCTQej9zIAl2jrj9UMFLLjj4IjCrfIACX9SSZzVIxCwN
J+iTBYor/dJh03AwcGFTqiP5Fea5V7QmKD0K/6TyNoCSsI8i65a2Uf02BYt0ZQAL
CrcpFJx0IZnRU+j5ON0dfJpvrH5nS8gjhQ2ieKzCGMUu9cq71eHc39laZpuCBm9S
51bV9K0hB3zNEW+nuGiODUC+d2HKyrbvas2mzjwCLcTD7s1FLrgvkFs+jVjxiQgL
0Ujf5fnqFOObhNTNHffiM4D+cqoK66sSDTitLYEWd+iZtJIwmHn8vAMcQFzuJ1lz
+Ntmqn7TopAOUkDfhQcOoID3Qsxd8ZrlxM2CN1T7EcXIXYp0+KyifFqPDQDBQc1s
jzizN/SmcoBb9w3llsVLwNgGHPYFSvnsFRwqHkaQiBDusHDVYxL9oS0Tv+si4kve
sgNWgyCnzL6LCrzlPFbvzBDgGb1nbkKJ1e5RfcRAbJwTklYs1rU8rMy9qA0vPtW+
CLeymn2cVmz+VF/oTZ8Fr4gbfVVTmgNkk+GeNTDoS6/Cu4Yh8ZZxkfp3f4C6g2pn
lmjD6iml/pRRHbv2XFIR1QWlvX/hDOm0JI3KhrW8vL7x3IY9JhFRDO7W43VpZbLa
xQzQ8YQuSz7MkQgNKsju7E18ONiqiDG/9jT0LrQsnLhV5+ZT7KAfe8d7Kkx0sqwb
qwGGP/1ZvBa6ZhSJGhkPufu8cTCGTHFVT3ez9sPAukxSnCkZmrV8XH9NRkC8EFf5
Y3MUc2VTRGu51GnAyQHvM5KYM/bad8i6/mfk2hq/tKaYMSVaPBFTQRzGVmURiifP
buxyedNQEuJsjxtaVbcmrPZHp0SpT8KaUd4abjLxmUiuNOZZzqpXTy/Ys7Wv5EkJ
SmH8T9FWlcpATRWBNqB4D1OTlECc22TX8tvd17VUg3Y0BI/6OXYYQit/jSBUjPvS
7lQhQm2iJH0dWmTQDDsCfm+Co0agpZQR5/E0+p34wWacFm47JkxcF52nEUcUCqV0
vhNS4aqH7J3+mZRqhR/EGFBjWf0A2BYihyzn/YkPVLJKLVJU9KiJHegIKN+wsyFC
wUjOH6n2ULPwqEKL6JRpUxUYet9qgoaDH3vdsiwQzQuMJNE+ly9PpScxmEIzsu3t
4w1QLdSC7PAK4ZGO5VTTeZmtGldf8esLyZEVQBTZyWnEUU0TzezXbVTJ9GrsJxdj
oU+0WmpSBHvsFppEKL/yKhxzmobgHKOeC1Yieg0R1Y00nJoY+TMYjovrmE+DtBgS
Pi6mhs70DZAhs5MdnIrCh2h4xh3e6FbJR9UGqvOkvzbzLwwfgjjRCqj6gUyDf+9D
flUWVIO1TjiRpdhfkor+NAiRTj+NADZ/hJIim/wtQ58f2ltlrFvEYVA82vPkScag
yAHVAh7KR3WUAjSaZwBXMN7MFFiPrY1TSlHpVRMxG4nnkIam9gUokk579k3Gml3K
zA9zREfYLSQ3jA6Erv7dhlnv69v1+8ALEYBOgBqUBxAbDhytbYb01iNeu8mjepTd
gFUkN70TbxJb8letgxnBHXI+omyImpg9UclUteQU607uqHGNp9Wx0e/VczFGagGd
wGPzTZXhrHNLg3aKe8/dHRiLgIzSze3mYoOzkS59jigqS+qPiDb90VUr/4yM9I/b
vmK+TMT+SxlGgdz9Vlw/Y4qwgoJbP5mhOygR+eoF+dTdaHogB2TUBgobRY5gRXbl
MHgehNCOInNkStUoE8MgCC6aEfVABo3B8cl1WPcv1fSvMffzTKGqjtnxJ+h36wSS
J5yGs8zwEmZkoWBAKRIMvjXs906NrVjIuaVU5tQGtG/xVdNVUV65JAEMvUZcXCks
wY8N6qzKWYMrzF7Kf7E9YYrs3u8CBlnG+OhJs2fmwJae/Yv5aoNmGMftrj2FfI4R
9CmZO3yeBwaMFubjmgsjhmftPOy/cNSYiZMe/eX4EAeVhr2uYYvuz+IwJnVhnbYS
1zdzWsYkfovhkhiPCNzlOGg5KGCKipyUkhxgfoZxI4PfQjqchK8RNHwKsbwDBews
v2cpPk/XSFvuWAdUhZSuduQNOHVpXGDhkidykTUnZhxDmPJccl60znzp26azZ5KU
RJnT2qdn8J31qV0OlgiKRqJkxC6zg0QUsgJLqJkKy8eHO0sl31e3N5/s0NHlvbng
VmOrUOgjljsidGkq2j2wKuqhwiU8f+8QFz0WBIqXlzN1ef+Bzk6vxTbUn4H8YmXG
d53vJYOiVviEAIpqx2AEjy9TrNXdhEyDGQSKYxOkKsv44jwM20QlToZlfrv3WFub
epjC+v3R3v9MSYttQUPMQRyDUdIiOl5dG4UfDKES2+b1mHXjyH/x0cQJXNp2Rdg+
fIc4pT2naWYFZKE0icIC7e970+pyjmjMquQhBbBQ33EP+WpM9INgzmRNnFvTWR53
+5XO8gUoowVUnca0ZB5IzjGpbzh4+AIgxP9Axi7iBkaAmW2GaanNoM93ZRvr0KQb
d65dvGMQoVFUCO3huMUts+rIkgYpWMAki1iWxmGXx8dLzx0JYC8eqsL8hR/fLkOJ
P2p5AFx+IN6NeqI38E1z7U8oqt7AAJODBQ4F7E8ZjENj2tiXdPL1GRhgRGqlmDG5
etHc8EeIUz21XuLei0XafWtiNoVNTdphuOaMbSYk0FZXHhN8vWP/DwZbfYcoYCVX
llZLaUgEk5ddYtZ3/xJQGlWZcB40s5sd287i09nlvr7fJo/oALw2SobZWi0+lJoM
S9yeJNwY6E44qRN9N0ElZR9djMEcnS7sfmu9IfVqq06CR683Jc+8co+HZ/KpGj6R
MaXfi6A7Jz6LIiSE9JuKXewaqfNm2vCnJ1fEfX9VlEJQrkMmz8pk26mRG5HYfVYA
vRTKY1WLs0jfB9bJHfbj/vtGsnZBicbfNtjfQgLAI1IQV47pIExKv5zkv/ynXoG/
HF7AQaMeHBz1KRJdjj0Hc+1FxqP4comsTUJSUUNambfkJPV4OKxWwVRcbiGZTUM1
b+2u/RQPGPXgZLayb/W3dctsWI3PnJRUIXABDUjxfPA+pooulqDoKYnssXvZzknN
p2FbPHtwjhgF6WjJNt6Tabj9PDOU/DiHcQ615pNrDXUXmaZJpyYaMx/yoChNUxF/
CyzywnFKs92CdLbirbedTbJ0lFL7WoolmzD1Mvs4y3mDX+mK+i88jX+3kfJ2WGTN
hVPa+If1AUdzogNe4NaYM3WWsvlhPameV/G/t5wOiKogStSj4rjBTyk8M5iDUYig
C/OhxnPX4toyRH8PMs4JpkN66uJPjoN+jmb0CFcDBkVEpxAFCKlhObHOBfGl8BaE
Au3+iCRL1AojQad1VM0/Mq9XBut6XDNGlhDSSFK6kc/1zMv0a3tWFgK2zUXcW0xM
CI40d6CMhZV1xAjHjoFE7DXi4hkl1OQuN1GYdU0LRpBnqyaXU4wxygPTWujkFDOc
2oaFPz8TGcSslHPXC+XaBrh+dl4RsqIXRPwJRYK8ZBkcOPne6SLFEsa+j3S1h0+M
d+JT7s9wAtLOOLW71lv3UDximNANplwW8ZWA3Z9ZlgvYnL2f4VGuZAfTjUcpKxt4
8iwecncQY8t7Dp6fJc3NijEewhjMtbpda+tELlgofOsmMvmUF1P9TKPGGThF2s/r
ks39IbPeTG1ScEd9gssRLCtJllz8XBIhfc9cSi/SNNCxph2PTdsWgZBr4ejVorKB
uGUWFIJmIPOvszth1LJvcZ8nW3xlwms7v3PmedxA8XLMX0jqvwaEwlftj2l+HMYz
fz1rRI2IIVBDEBdrKELr8TC918xEZsfAK8gbiVHwMsJtFDFKysCgceZ+DX0tTKaN
Wwx8pGkLpZ/xUSVrzPiKSIf9tb1CxLjJZxAtT+0KL9tT0RsVKqS/W4g0r0dMUTO+
X047BY2mvNlf1ARpE+CRBo4dPkiJ4DOnQ+iiekp78qn4wevRhY+VHGkTa1byHRgq
iFaNNueDqIhIxgbno5YgnkBb2B+Py6nRIZ+R5w0ftjrS7ge9eu7U3aboSdybzvbD
LGUKFB7somFZy2cue51ZPfGqhGPc4Xg1IjQfflGsO8aXG9fCuRyydrJ2L/oqmmcb
4nkPrRvsaNMEUHth+4+PXGmV7k28+prVI9mCmKbJk37lbRvFZVl/9ZzqjnsBx15x
e8V8ogYxms4t+qe1Lcnkhu6tFiZLmJweE1zb9GglapJP5NBDFK+fw9ElH841EqxU
rBN6/NFQQontoeplfaM6DU/hRE3o5OeDtowZx9gio1lyuGZqR0os31zlXcmSFmJa
oksPAvcbWeZMWjRtYY9P2+WlBAb0AIV4hj4pT3O0bepPA01rE3mD/1gubEbqC5qV
nVC4VUrrhJNTv+CK/S9bvFsw4qhBIcRcAeubJDd0AD+oDSyn0i7WefrAvFWCZ49B
Dx5wdXXJE80fz+m49JiVsAYiT1ZGnlbDFPr+ggYwredN9P11LB8Zg8THLbMokQYb
UUZNBD+Eq4k70oOMl0R00Cgt85lrcndgKGVRJ617XJ8MXYy2/t3FOfRtWW9OsSN8
MHeYihiiz/CkP66sg1WuD+mhGCjM8XVYpRovtNn59v5c1r7pUMlcHyf6RnZH3hG/
6s+vVxHh8VSkZjqHfAu+vMlui61iYnBfU//AThdql0bXUm54hUYk1FM59fDK3jqt
bNcFbSWIY9drS5dzlr8DkXMgwEcJ8zdpuOFPdoS9jnR5CMTpTMQEYg4sy1fVNC08
QfoSmltrGqAh7zmmMN+BG3EzcmpJqACRfpuVtES3TjIF4quWVOrsG5INysZmD842
5KQ+7IOTrbp6qm36BlfG/f3UpBNT04aOwkQNTgaHa25NMvFz1rDAtFLZndPTg1pu
G27WxDTE8rBYO/uDbJy3XLk1xLrwpvZDIHKlJaPZ0eIwy43l41Ok0UtNY4iaru1m
sNVGRwicE9/molL+qR+qA9rxNWqxBLhx2VBz1RLN+gskk7z0jPnXMgdVe3YJchBV
8kMn7auxFP1ZCb85lSpeSG1YgVSvTUOWTzviH6TwVChPVckXyRP7+3HCCtLqtoEy
7Em1vJFb7Y4V/9NL78bu0V2osoSVzsVfNAHAK0njdaw692e19wWvSGiLnQDh5+AS
GiRCfPRmgG87vsb5kxFAOyDTCIkrQCQuD7dkWoJbr2fFXTYkUdBT7MzaVc1+tusd
+HMA5Tgb+JG1mDrMk1MMAQ4PUMIC9b95+uZQKPS8HT2YqahhGKpkubDZpyft8Hc5
avb3NinQzAhdURB0bx0O5ix5f05ygfOkcd78POvKf8acPtI4AYIdN6+BcEJ6CWrC
jo2XzhkidSEYh0Bc6jLCBe0WvpA0DAiG8skm9Vt3R6Gwi8vcpVvkYSV5kZzQa9mv
ld74p+NTilHwHEv0htuTs4LHm5DS9RSvfm1XEYopncSevl528OYcPgkHY6frnbvt
vDjC6erU3zFq1OnUatB3fXOZFEc467Tqxoga+7BdOGG2QiBqL9naFrCBSRMRKQ2l
lp+nhhP5pa4h9O4NnpLQgmutATjYMB7J6Thm3CauP+pfdcNLbH2y5LibCXGNzFt0
me6xUbZhMJb6VbVggtMPkKpmU1cExCwRdCvuousQ6x8Cy1VXQZQk9PzEeodSKtWz
HmFSfVZIsNByoFS9OlfdyMmhgrfajnGNfJA2RQWfFijwNt6X+obz6zoiDjCYms32
BJMUtTP6eUSc0THiImYhhl8P3EJFODd9nwMLat2T0oAY3OT1Z7OfYpxfjAxl8ovR
M8iMnX2WYrp02d/mp6Jy4Se66rJAWrJNIB7D8jWYjScAYqWCRO9vDW1vmuccjFz+
B7j7aaC/BEXAVu7ZYKAOqgaxc6U9WjCwraO5qcLZR3TPB64Qj5vC/iQoTNRdR+Cq
HZ+7K+xpwDhCZF9AXY9U5ViH+Y3XrVE3u47Jl1Y5Ji6lYsqDOjQGc5LmFDFzfwt+
1WUai5e0+1yDCGEN1uk8snxl8yzakiNL4Ez0xIge6OnRKof7/4MTMISBqfuz5myY
dTmxUt5zAALGU83jC27VVjbzzJfD+a99wuxe42t8PoqTAh+UCFTYRi18tz5wP7yH
gOrL5GhT4IQmZ/PxviLlVRSvFou4ajZtbPqlraHWdMuD3AsCZJu+SW4gUzfTBT9W
1h8ygKII/UrnmQhE6+slQ0f5/l4D6dNYfHlUKc+vgSFjA0ffu25dv+ZrpxeGK4BT
Fxk+DKHGC2NR7CwQlQrMAVStVPRADFVmJzPoOei5nJ3dRCtpnI3g8XYnNC4on5kL
eDbqX79v/OElaa18pxur4YVfTEr40FN/6yjCcrvQEU07q7Ma5fnBsyxMIiRg3JJx
nqOc2sQAMnGuGFf55F/667C9qi2Qb43adzJtNcaK6XyEzqog90OQ+BiN9Si8AYZi
EmbTQwpbdQQvH0r/vVAvi7mXVvqdJnfjXkGlSOxBhvk6q7FCzTuiN6fXqOM4eMB3
jYNTpcSSUoBlj/6OO5ZilICCOsoCbFJmMVqea0CNY260dIqm8/Vu+QZ0czt9Lg0X
Q71jpBY/XzhKBQ5cPihbtsMWUsJ6SB05VPES1+1NowH81B0OZpIlYrWB8ylSdPvG
c6VLWhfr2OoX/076puAJCMn4WbZ+jWQq9N2JIhwGO8FSs6IEcR/jFbwInSmxkzQK
BtrrmCXEL6DqVpOaQGg/L6FyWBbfAUy//7leMktz+AWpq4ylE0aYiRvvLzi3/3HO
B4b4aJDKvq2OBFUyMEyt3lfH/XNZconO0enOqmCfpOBaNItSmleRsqi1fcQwajh1
ECTS+lUYZLe9oYfDItEDpvP7NbyW10YhH1A9ByY1nuLjMeBx4cqgeCuh5JIqFPlm
ueoIqfmNd0eGnzmEV3hXe1BqCcCwbau7cQG+PPKdQi1BaYpFvHNtC7sP3kTa1I8Y
lKuOPfC5+aQgaKBs4yiBBtMbTxwNPt52ypa4aClMKZ9WKfNba3S5seJGVyCkta3k
araiy8npjiJtKxGrSc1y4j0mnDyQw9uE3iBovTmlJU0JMieH0oOf1GI2kxGPpkwB
ZjOm/FeNYRt2LUz4Q4Udw+HPrX2A6QYIZagLLmlJU3BPvTI5ek/TH7OrmfNtUvT1
SUkcQ1SNqhqx+6UvyK4RWFB7x9wiW6m2SQn5wrBWPNnGdC6paWduR8mSWlH2LRvW
uKDvTwOLnMTtaCV8rCUxd9K71KdxOUkxa0wdvg5sq8nxgieNhozovFlkIlLt3NYG
Iok243Tjd9qBPbiMGJjwVdSXFoMnUHLguCfxYGBTGpNy0AGpxTlZBcjmC2dHmG6A
StRgxv8cxOYBY/AheVPzgEFMnuNjCCcPpvDverLTTZRFmpRvpTMDnFDUHutz3RlF
dqsDyM+ohIsHJMp+hHwW8S3llgbuvj6PvrwGg1hhPhVKfJsOjwgGUrIDFNjsAfdZ
RUcZPMvV4auncZe+GhGRANoXfq2T+aqpbruSlgjFOiP2TEQNvdXrTuA1fYpAQ2Cj
Azv90Nfa/wjtu+PHpl0+vG1xtT8SOxEtCMvsqv6/2DiKdpaAaOuzt5ZaMBlFfDSw
uhtR8k8AaQZzhnL5RBJHKwgwX6CjgREHBJAzUd4DGoFAHGISMv6icqK0jx0/a99U
Odyvnqn8e9n8+JWDQ4eHZSjJm5j1jjMZmGY6k0mIJzbFuC5Ard7OUvsF9p5J5Vg4
HbbNk6Pk2VnNrMOwALV5x1/UlMgVXJas/xESEf4weOipI153+o76bQgDFfxEE6sP
ERiy1D1yiUA/QqWZ+842Vk9mw1sYNocdva9Ryl/nWnUVTEZ2p3p3PccvCpC5ltv6
lRAS8QhsDph3IXjUMj7bw+VQB6SqpLQiP0IMvMuplb9EXRRzrjslLTMW/cia24I4
D/4sF0o3kzlzYiG8n70Rfh02fRw7Q7KHkMKG8209TmlZfYs35GolSfLDyoHEK+8l
xx+MhcYu0FKRjs4Hlu3VTf057Irf5xa/HJEnLxV0B0ZLfgr9YmWtLXOLOJutVqpG
XW+WNIabBtOyUSvlFI/unyPGSXwQud/40YtkVskzoyBy4HxC8FaP+yoYHHNG6lby
TxJ9mT+/98I4gxtwRADbDGQLsJYOomKDMqgY2M+Tz2CwG3yQTrPPDkDdtpuAtVSt
ZCx5u6iPOy9xcrDedW2OgtDH7qGE9W9D1ktSliWAI8FyOXa/1u0Hs9L8PFSe4K1Z
omecOFEEsEh1pA0h/n8A2QPF4PKYUZJQ3WkreFFd6mCQj7m6gNeuCss/e8fNwsf4
LSfw4BPOUUM3GKwx8+J0WlH7xzxTR20Slj/NlHnA6HcvfvsyhJF8guAtdzrrwSIJ
ilAitWpOp1M1g4MBwK2bpiE/x44FEyVbOlIo5r1nsIMQ0LVpGaoz2Q/wCFKfeuQ4
pK0RzBa/5YqRS/UJ9EX5GKda8wf4Paut4eDclD4wirM9XRhz21wvqu7+ninm3oWu
aLRGqMud4e+ED7Vy03Ue6uqxCRKmz3TxVZzCjbn0rsaBdCsIjuUoho2CsP/PqHKI
D3pxNyaM9ROCqoHRcCAik/lMBX2hoMbFECepxQJLggJeIcil0k3x31yMcR2kbtDP
y3NvQTd5HiUNw1RrUr67Gr2GolpBzVq0+rcdhQnWDdfYaVX7f3Ah0D9pKMrXji6n
2cighgKBZmrIy0lQtgWKRJ3mpWC5xpu1/+RJULQuKW68aQR8kywBCA+ufkBNo8dw
cEfQ8dy6t1StCdIWUagLC6HZnXnv3+gnpDfzGT8PG4KSTdi6hfosWXQc/LXxC0i6
VSaK4XB5nimBi28jM4swQNCpUQ8n1AZiyHp3fICsFN6cq+QQI8vanFIo12ufPdAp
IjdFMgwFrLXJJ4N747ti+3VJM8BK7dKkj/aQ2r8cQc3057r1w+/u1z59/B848I0Y
WtAYpiqm9qAt2gIMXPViVFN26lkZH7Q97ZEMoQJjikO1WjxnLbwJ7aJE9UmQWrTa
oyAXAsPhZ7aZHIiE99AWfP1Kc+HJcmzvBOC8Zv7FtTUw21EnL8wPr3T3A2kai5Ow
TbAajl6m/X66ymTawSxDtl6tpp/OdAmjsz7lUSkNGyaN4MLlB+bS9i3FNlhBjrGo
7NlGTXmZZgwwBpq3gZYIzg==
--pragma protect end_data_block
--pragma protect digest_block
AcPW4Pw4k379DqCoko+ANg/mf/M=
--pragma protect end_digest_block
--pragma protect end_protected
