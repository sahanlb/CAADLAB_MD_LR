-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
KLYyU3m2c6Hhu4xb6kafnGDZvUlSRRXxxjFhgfmIQiMeaNv8Hj850wx6qLc1Ju+x
ir33rDDVafmpl8LMIgFMsg9UcLu6IE14QPfSvD0tCHsVQyusa4bCHXNYzV0E+RNs
KYZHw2hi5hj6RY0JX2vUwvT5MgYZZV9s07h9E45Cmv0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 47967)

`protect DATA_BLOCK
ppQUc7R1X/qjemjmGgYtyIB35bA+tQrURnTwuC4IwZP9b4ULO02MxsRPc8ambRV0
7Ohp5o1PCumGM2qeZjkeagE7kvZGQVzCZmJPocyqntTO4ktwxhkegWkdjy7Jh37J
xFM4JlfHj21/r0PMREMbGi/A/IQ+KdI9muDv91CVlY7wGD/ptY2u8YOirBhNUfYj
DyByOm1CSD57xDVWaWZXBGcm6ufXeoMgwdIIz82jZesiiqag8r3wDImp8VZFVkV7
+Dnrp2XNGRj/HrWBDpsOgPZZYjmGM9JRM96N4cOvMMJAaPI0L1hYInKnu8N4Cz8r
PYxVVYne+aiUGwHTILjE1uOvttn2JUDYfSJi/WyzTQ/HddTEKfUO4t+AAMHkEsEz
KXOmZdvaWtv+P8BlaspyuLyjpFuAO7QJgMvlnEjyKHGcXwoi85ubZLTH1n8+M/N/
CSh/TNm0uMx1eX5nooXD1YwlPT4qwh83fHbFF6R5UQqRIt/rIkxoXP6eTZclhYMX
pQok27oNiv1dfVf99+XSEFSdawupwTCXgbu6i74ZKYRQtiEhxiozmWyZtRQIdZsG
VXFvg4RrudhzGyIQe4zCc1qu6R8sCLNqYVhe2sga+Qz6/BsG/Ogel/AJn68QbwLL
4aBlRAbzBspjk0H5UTZYHaaD/IfFjfNjy7sLo2x8YFxkA6bEfv7PpGnZGA18Z+A+
7C3oaKDJaZYc42Yb1LKS658aVYn2Qgz/ofz8CrDWN0qCmU7HY78MsEDQEDMs05tD
5d6qr/toRZjxwh0Tk2bFjTEm67alEP7Sg6/u8hbnWr+L3QwsdPXzG+1cJ6a92Ytx
FLJxRENmb0Q9I9rXCk+VgmBWTEhScQBG39ywsjM810btXz1SP4ET23EjUfqWF4iP
xyIonRgT/9JUelF092WkIl1sUvS/O6aHamvMmFD9qyHr2YmVEECij9g7vb5pVr8M
mVvIAPTMnsB6jcj3dtJDXNeezGjICxs4Mv45sEqXOXk7fWAbRnoqTE3W74rC+q7R
dAK7Coq32U/RSKvQnrR6bVK6Hwo6pyar9FbGme5i7fdwCkZyAqnEIr4WpiMUSVbz
f0pXC4Z84NtpyQnnUAa2bzgGrM4awfNL8HVeSU/3tUxNL2J2NYjOgmrqe3rbDw7V
OowWlw2ATmjm99pARTnHto4OXcnPHFLBw6P1c/DNhmD7WawOXQLG7YBJgGqSZbaO
PJ9a2oHjoxdIXQwjNM8tYyQvv+lTfV2TL5XHMR01yOWyiJYJziPgN4YOP4ZiNMXW
o4zvFmS7FaYX/6PjX8qjWT0swTUQYQJ2mFQNezYCdRPH1ngHRyd5Ttb2iBk1gmqu
+KCmDCbP+75uShfVH0EW5qYETxmcWNoaQZKDVcjmioZopqBCEm/8vZchLDnpOzFD
+mEPoq/GFYGmYcMbCmdw6JJsTUYsI2zGpWG3YErTVy8dK051hvb6MyXGPhf3/4fx
/lS5Xpjbe5s18zAhNuvJfqrTwVmuWK4215m4nAAqBvhkrEfMp5m1kynRfOxA8LqS
0Vt+I054G3bvsVWcZzzNjouX70kAg7tNdCUunRvWSor9PpJAJamy41JHgCTOHKnX
FcrmyaBUAFG3XPy9QoU1C7gs9dXOdfqtzvMwlOCvFKdUowFgEFwuqDSHfv3rsyGZ
9o7vTFypJiBRyartfDXha6DItMYXRHH8FqRdrJ1D7RJB08wDMx5YfQA5iTdkMQ5t
LxQRHisntaBXZPpUzig3Vg3fnvzJs2kpptMy0W+ivPfbrgP4pkGFqCAzCBufgQew
LkZuOFNDP4cNc3DsX9J/pQMhwT569n6ZBP0JPvKvSPHruZMyk1jCRi87GZ8Q6wam
GYVmlcRTFnbzIzdY9LcSXoZ7TCR0oK9QLhp5AN7e1NZNT2bfnz59yfPAQ1sl4KbF
lmlHH/xB501jX0q5bvN6H4o1n4T+uHSSgi7KMWo7t5TSqKOOT8cQg2w8imLMWAq5
NjNucs31hiCQubHvTAwHgtY0xQp5eTACCex40H4pl1tQ7k2XpxfwV9d83UM6n1yh
CymbOzOKfzfIC/RdUtFd5UzPP1rOQh/QzEWZdPFzAp65hr/9WO3p7HVPuEqXaWqu
LjPV/ydNz3gVfoNf/RJxAcndoGy0Ku4N4HeNQR3AiNiJJecL4TLssqie2DWTW8B/
GCGO82J804P+nhwYseb36hBKXsuYQXzY6Vg35yIIJOuRLsLspOKivXjn8egcZJ01
R+25FUkoGoV8HltoGlQAK/TylDeW3tDPLWUmlpr4G5GB6mbRk+EPZ2Q2O63xx/Pj
bpWntskAsTwXygTGEBbxaNy9N1O2H9oC4Ueach+8RHwanmuGWQfnqHSG7mwLe6xy
QPtJ7iMeCCNeAvvPgogDui0iWSFk7BocAhrYEzI8218NmaTy8yKtGR05W6RhpBo5
2JX5x1LcXGheuYweqtqWxPRiMGlbq/RVGsDSwvfjXTkzdIFNAtiucm2tQoNLwuVM
pNTD4D0X1uVUNkQwW8Wa309Fo2vkrpqkPVwy28kP145aNPcRnZ9WHuOjpQaICsNy
9wGDzT+bkHSajIAa2CXqiN0gVEAOGYqZal7rkCcyebC4QMRFWUYeCfIM9lenxkVo
d2RgkBEcYkXvzQTV/t5PiaaGhrhZu0C0+vJDEDcaFTmG0oLv5wv9Ff2iSZpZYv/J
jPR1yYYQ4+ftvSGhj+Zq4X/HA8aG8k1Bd9p2nwy9ogfq4g87LwV5h+hAGWurZBGK
xqUuLBGkHOKwV5UzvWyGO3Z7mo4OuIjx1HReYW7ZcTNu1wwpUdaCUYCjf7WY6Hz0
+gpQVR2116V9Ta0H9pS7CH9rZwH1qf17U7jomj5hrnqcJXw5Y8xkjzhjY0DAV1VC
tksiKvjV4+9skTYEoXMoHpV0z/UvZwqaP5Qa7ljgi+rhgkr6Yz/V2FOgxuyPBXEz
TblVNJCc8LvcH8cm3gXiH7A3bpPx8B0srabXkNPhkW/XwRU+s6jgNJ6+nFzXu3Wu
O8ja36rJ0cddj/lXjT1WispOOvzNmNzMPYqMiD/ZdFA9ws03ADYR5EXg9bws7whF
N5egNZEMkpvov/t0PCbTdfG8nOVMhNnS7qTXwQS4SBUhwHWoCtAsNlmcrghcK5Rk
UyQhxfrN08+yT/LJGKfwctYIJAP/CqoLtmtbshtNxR4xEB1m2xY/KIjWA0wJkAAw
+ZnZIme3D8TdKQL6/EpbbxOsb2ZHEgNjowHomrzJqoZGhIS33KzbJPV3P9uW6NEc
xi7YDvcGoKhH+d96CBZSCq8vEdp0P9nxkOQweL46K5CF0zuLYRO0Eumi/EYZhuP9
GnTLCTOY2oAFW7zO5bzmYCdJn4D5lNsndNn654dM675C27esHXUYo8hOwvGCv9TJ
0cG5AefBSokWaVjOhpEN2TJNIlt/wXib5fMmh7RYJJGvfEHgcZXYCi6E8eqwXMkm
U3DRvYNfSkIq3tpe02bgs4Vi9MBjLERCz38M3BnPjjdGtwYa03LkXrv7xN0W06mE
Kx9uloM6AvEXGmlGl+nvuG6ahlLWE2c0fAwU+mlMvobbKXM1q8AmldpehWnEE2M5
7BXX4BT3qEJhrXauYlTWrj5DvlgerhkMqQ4qeJ5VuByuhZOAtm6pUPAzGLs8f3hd
dyQPYHnNs2wFQLF/6es7olwJj+Eqj1NmFZmTpwsfh3DqS+vAROZVXdS7/Iv5BM7x
FBPucp1reP50L9fFrcVtn5Icz17aVlFe8bXPFSvlh8KiQaHQagpGzH8po1BC1vdj
SiOSIuRJxgPz3vkJw4qpu8PuSZUTnmEtrTP1Qrlm4W5tEmszLaUZbSoFO1kGONwb
uwkZ5k1/aape+0f3xFXkn2GH8Bh8cW2PL44fw387GSDJFTf0/Le5u6FPQ33v/MVK
3c84ZyUVeDwuZPJljiwlcemHddSyeGp2rKGRWtDpWu1+k+ctXOWynyKhEqiQrklZ
p7v8Oy5kx2/ns8PNpT0Gf+lwP7BVUGsIFox4kNtYQAoDWOoiDdSXWVDNv4s1zUoy
xXFErWtpGNiBcWmx1k7wS5s3/dVgajzt0rcMDXcN8hrpwnuDtrbk0pE0id8fExmQ
jAAXAPs7WbJ1eMXh+v21KoEPeUEKKgfF83LCfpT0xGmpu4drf8r8pxqJxHp+bEYZ
6AT9Lb41q/zJKtDJYnpFEFBo/3RYRqidlydyAXEGuyLpQYM/EyQ/JgOtwH15zaKv
WsN92Jl+Pdqg1nvxJyFgSMp1ziNL6DvnE9Mf4AOuGjFK8EKuAjvzQvdpH+31Nndq
ZQjg6RGOZXEt+VMEPgpmNXZ4NrC8trW0fzuLE18bKsh/ZTwhxSOlS3oHUQN4p8+J
T9X7KOhDLghM/zGfJ+uDCglhZO1gMBRmoSrrNP9g5KUOmEhDvRlmZsFA31dXo+05
bbBULk4kmyVlfQvrcZIGTy+s+q96WHQSRSyH9eSB2pWira0wggs1LDosfV2/Pci2
UeOghOYZMoGMxqxb3sezg4FEqvHlZT+DlN3lDC56gl0Q89IPk8Zf14QLn/KP+0UZ
/3F+B+sSCc9M9fhFdy9hqK4OBlvQmiJN4d5zWvoODNhkiJ94bA+2+X9we+IYpowA
vw3a4NwopAPovNA4rLtUiftYmi0ENtTxqMS39W0mg55ELuKE2tMtXP7Vt9xAbNUz
bhoh4CB+mu4C5UOOaXY8M4JKrz0diUQQQPp/A3xg/sNNNggwsTu9oNCXxqQtxZP2
kY80B+eY0bxbCQN5cc0EMxRYnHc/BJJ6X18UbQxW3CUbYbNKWKJKzxFnXNmCarmp
ZlTvExy1l9Pd9F6Tn91wd+duQc5oaqtT9f/g6DxHdggtaUcWgbhoblPZvRH/4fdz
4BajBxwzDmJ7TOHV2m8SHfMGxSvNN9odrQJGtWAosakP4cUx8s8zhL3ZgTgQywrr
U5lC7MHyW1Rr/I87QFfvCS52hJzWXfnEn5LGPmuhdHiIk/cmXmwYtdKiU2hBMyaU
dAgKmk6aUb8yl0J7tQhdl6YeIhwzTIQEv0pzbcXaGXoKRcWRA2y2aTmuIYaRmIDo
7NPy4cRMe81CWToJMX7IDe4TcVTQxE75iswOwAHIh9HyMd52lNUFfhUuJjb0UEJz
y+ayC9TS1KlH1qdaOco0b9NLcnWafzzLUe32gnRkK2krSpU3hjg0lnn4lB5jIWuZ
BV4h2MQGSSMQabrzUmGJxd0bmnxpbXHfwH/Yaq/sEaBqG3EZFUjmlPWHByBVxiEW
QN8bIZzhJw1snLjWc2bevBvhIiUa2ollMF4nOojfIAJB6U4FmqTGlAOYIYU+qxv0
jl6FDarCm85zWLM6VX3qNsn/dUvRmFmy76MpxrHMQggzglRs6GYDQ+XsVvWHXdwg
CqmB01jWKWfMgjaGCfwQXACHxFhCTtinylMXu+DWKfq36fHJ9+JfMsvCZkUvVWvr
yyRRONF9BVCP+Sy+JoSVrZkKEwO0T0HmY6y7XBQ44FJgL5JYCEMokMjM3oaLToTI
JHDiHfYokgIKThAqn2s0+Gs80dS4AQ4pSVrfadHlP2jcKvQ4a9W95KyNJbx1lmI1
h5RtD+22azBIyTjuZWdoBB60ebjsvuc1vPZ+nhMJZBnS2XFTva5VjLONqVhsX06P
YGtfz+gs4/Ybbzi4w+hPErPE/lc0zeAeZpnd35uFYyN4a1yahyjcbTQllJOV/hGP
Kg6jQLTmS8wT4rcocg3dqMY9O3jgG+34/ZnnVIf7hzJbmKlgabgwcLukNJqgybB9
0IAqqf2Hxtomvz2w8oE3J4/umoQIzbyI2HYtvZM+kyvmhKIkNWK7dj1fAqI9Yl1V
5E4sLlgx5kzbFvFq9JXyfrOYx7suBrTL57wtP3tqKM0ClnNwr/WN/AtrvOVYGsBY
e/HP82sixl8ydz+/JfdMqdCOKyuuQbaA2HmKprR0NtLzkaSRnSJQZK80lKs0m3M/
WQqUhnsV4nEgqIfB0woykK4vXwvJC/7RsDIvRjHWqZpgjkt4FKmK6ckEakTJrU7z
MNK0+r28NN/QQeb5O/LYALgqBVYLBwM7uFpO8MEdzXD1ZPw7ZmE+v/GyY7IMMP89
KQZCU2CB8xJAeunN8Eq/yg6jUtDVv2Am84O9n6d3FLDq5NZPrZ2o/x20UyqGZFc5
8Cg/yHo1HtqyJK1mEBmvYiQ5O/hUjVCbMg9ruP/CPPmemARiHA77xhUIwpqoSuAE
3K1VvpFODaMEUzG/+CmirneXvHjCH1Ym1NTSah+oIAbSVxmKRoYQJqtDemT3vbvv
7fKkmw7WsyM4XAlzwPBu2dWCSDgN9TTnLgpYQvnGLiNcLO9BUwtVJiXm8mpRt9mS
mTRaKuO+g1LVj+epnmMh3DxaohPbVtikV8IG0Unp4DNGl8sPtPOmOsf5QvBR1Qpe
lucB5AfT+x1hFag/aVLwQWOS5MlIFfA3cPos9nCWd8X2uphiX2CVATTGsaKMoub+
mk/uptApAxreYzYfUbNNYzk5kP1LeHyMNv9LB+S2u9htN9Y43FKbybhr6pft/ymI
hEdhbQJu7wmwRgDeAMejJxa3Q8GtO8ZJKwSb5NUKqD+s7wCYXgWq0lQN+UEglwE2
1Mj2QYzs7VwcqPyeJYLQ8XSj6kWIk7FlMSxWyeEWMK0oztLVO6soVOuCuJ012zt6
DasYrTgODmssMQNGnhYWRPtBu2x7Xp74TqfjCPNjhHCLcdzZCDIO89essjN9Xfg0
1SKafgafp0Mk63odZTXKnuvSp1oCrSKpXNyp/1/Qxta9CweH/5VF/RcrMX3DFE7c
ZQLsvPJRBwL5qW6t7nvx6/a52NvF7eEM3/zcnXkM/6VIWektVCyIL+V2zgOH/F+K
RzMSwng3NML+yvGqhDUw39Iy4Z5g8u9fg00slWxdmdNn+VHlbEGam2VGd6YkHOmZ
MzVYZuUljhN+2uCVvmnN9ds/N4BgQb/lRogU+CZL9BMXtAGWbxQBnIWEsU2y5HZX
pmCpbQ2QxpPj3XzLWVfJCd+zpJNP1wbVnP520fSVrMZo6S8xMet1EbEhkzoHqraj
hpnkhxze6IPWzvmdFpspTaLn/q0vwqmkOazB2nmvBs3ibhXMb/R4Raqa7UwBk9cF
2RJy/lLM+Pchvk2CNVdwl4UzXkATnrD2LeRkScE/RXd08R+P+e08BWCQXXvNBn+h
zTwvq3dkfMCjBJGQvupKxQGc6mahOQJUWxzQjBpNS8Ux5L2hpU7AAk25trW5B6Cn
YOMqSxM3/osBtecRX8Zp+QZZIF92p2Y8uMmUE2ey6F2swaV2cWMKDmC80hBbPZOC
w9i5LePqKu9EVJQktmq0yjfoVKdGmN4R0vwamJd8bMr7zJio5WK6PEZoDFFAIpxT
Uwc8TPlYNdQCHrqUnMHeA+aUjDEeyUSGm8WQ4Ek1nMRKi06Ye3l14J126emukpyu
dleV+N4pbMtqtMpckFRxHNsn1xN7ZzvnlLZ7qIeUTJdu2YYdNDU4923974slk+0m
6HnEd9lonZxXOVM6XPb4sTlIqT64GgdfjIwvttzlUw5Mfg23g1igsStA7gjJ6wgR
CFvbCOlvLlisIJxYDbjHdeKDv/iuOlG1t492AXeO7+jOK9k7jk2cWsPqiO5qkwK/
RTWGV3T4zGSSUONr7OulZBm0eq2lZsNctJGXWMy7MOEXeutZnIMGvcBPEPUg1I6y
LSrjEAV0xdmgGv/+dzJwvoMIbKHyDrYZVUlZIqer8S61dHd/k6nTrw9lU/sNzw7b
EMdpA6CYPCDhHB/kqzvL/weuqeiY7cXkSBnadsWSUZxhnTebz7+zgIXHBqS0uIXg
fuXThdWLv+cuWIz4lGlZ9LC00OZ4nIx3xNQ3kGF2n/ACtn6oiuGsD15leCmZ4Azn
hbLTAoM+0T7G2fOgi0OpagFRwEZxhMyQO6S6QCmdlNGqWGMHAuupA7uFIKoK3rag
WNBiBRKStzSPHV/omsNERdkVlMh0MOmPF4IUZTK5bPIFCv239ePYpapEH3vtyLtE
CEPm3XDoAQB7mIQgP7MbSlbOOZeUy5tuFw+7L+ro6Wm72bugu87pnLI/xkmYXgF4
8eZrBnKifq8yvWQc0xOPPRboAA1/rI15CYtOsiWhPCajBo4tau86cufHa8kIKzaX
pXjbsM0sX7tyEiXh5+ziT1wW6Kp8QESsjvEC1sDxFgiWwcWxrOPl8zBNMrH9nTwF
tuHJ8C2rGVgMYeqKEFLu/5m80lvWznkgWcH4WlYakpgMV91yzbrme+/9lJNBl70O
x22RZdYCSOZwzlrMdDT2GuECSArF158FjR17Qjn9DW4huPpvodC5axczk4p+UBa9
5qaZExk5O/vjXPxDy7l0cPZoM9w3FdVqQNJqdyQ2NwbtI/B6S+BkyWHFxTEes9HP
awTNnMIZBQmCCFYhOCrnGTi1NNyuKtfkNLot86sWm9K0ybvlW4deu5vdmNEOZsWj
3u3rFUi0WpRiJpyd3r77bx7O/9HbSldk0gKL9kXQ1tyGjxOkaIaD8zAZaTwRb+0v
Lahw0a1MG0jwBEDFT6rFJdVNan0K9XVqgAg4ou673pNeCY8RPsMum2EXwLiBIwrG
PX4KXe4o60q7vu51f5o753YM0NpFNxvCnSTEW72kKYd/X1V+IGdKYWu5t7cK0UNE
BMJmYR7dNCWSN/cgQ6QKlfd5EJzXLvAzxTFuw3iAE26J2ii2Se8FmHQUWO5Z5y6k
9WvTLas4SmeRqm26oaMyWdTviaeJ235S6kxmYDadIHjOLXpNBzVbX1/n6OJVY6ky
KEEAaH6bOXogARBkCYgoSd+Vzv7Mx+4Glj3MXReHUkzZezGDaKNhqfaswHQMAZpT
zTjNgZJB1BAWK3uW3fS9iSHK4sI2PVyhDI9F7HwPXRJeWnj2BGZxc+RxWPX+rIG0
Ggtt/t7b/4Gvc9753cnyTumBDQMcdPFTfUTA0ZKZE94BE1QXUGLjdIjr4hiCQ/QL
wLApQVV6jnu7fWVkcr30kbJgSkvXuikiOo8PWe55FE3t53vkEWg36uol1/Q5llJo
086VUVof7956qs1eN8S5WDjV64kGR0eP2xirZJuhMN5h2HYdJ76fQ/3I8ILROHgu
dWAfpr83t3/YplSID9XBaLBT3pBj8cocHjSzpnRWxHkUx7XGtZkOxDJKZAjMe9wS
Dg2vGAyUej7ytCMYche3i+2OulTZMS1JV47WWQ4aZyToVTbjwToYqggoPUDV+B6i
J/2LifeP2GX2xHxURaImBKWPUD0hdSQbOYZLTBMTats54wDGh89W/K8nIZquUtih
NMl5alYi/9vfrqZeEFdDvdGCERaQBAkWIsMyByGqUbV1b+PCmcgeukUQWfFLJd2P
HNeLltJAnKAgh3NxBkb9rWwByfv2sv69iVZ8GUxHECxfLslxTofZArWiouAnwmC0
0uGA9ZnyCpjMGf69SowIn5JW46luVwIXPhYb7AtyYGLQQj/R7LOV5M7+1Lq+aEs6
lvDL6doeAyABqlzcuITUDkS7Xc2e26bSBC6OqgW7ZnPVgX1b4jvCzmFWgkzklLlg
hIcgqBq5egeRevumUnyfJSW2fG0Lh+Yg+OeLKgI5hmP9KXL8C8lx9S3ZkhAJ6BEV
isjqYo26PACgsZdujgQBy85RArLKUdmo/zoGtS9L48eW6u+60g0tKOPcu6Ac+Erc
zkEF9OQUzbuvzm/ZNjxI1kwg9akmhsdY8PtL2AC3+gapBXanQpfNIACGCtU6WT2N
RaMlc5quxcJGVmPtoZwdX+fJIO1avHqxGERnpydEbbGsnmDDCP1x3QkTXprw5Wx4
5lPF8dTSrGp+xzD8QfAT1xO8EiX5e6fEJWvcq1z1jAjphrUHSM6UeuhAXfs+wq4X
ze+MtKLKg2aVXwRjuiks8EkAgExu4n2+i+sH1WJFRUyI1UiPxySiJAKsbJYx+Vnh
uBIu4XfFKzoFdc4cANQUbn4F6PnRMoPp7bKTFyTb9JiWqLdZvCSe1fRPSzAEDI0E
nuamJQHUd3U0wPcqjWGxq+9Khpo7V5x9N3fs7uhcp3PeMBOjGHO7u0rmcbCK9rSv
3TxqI2/g+LMylM/rM2PHIgAZ8ppN3IoyP4qtvBGSPYfx6hXAla7UCTVnmNzasf+U
jnTmvXbhcBI2PofOT4giVzPTDsalAaq2I0sSbq9KrbswTJf8v9IJh3sjNg15tjnB
NKW/fRghaeCx6HGNzF1IdD+QLoSefDXuwxEIGnjWyya23KhIWjdQVlsenv3B+EVp
hYM7lAi7Fp4XfNqFJ5YioY7+xweX1a6OpmIzTeRSQ1NQpE3l9Ag0qtLciHCGB/Q9
c7e2NA8e3eWYM0rl1fTI6CgPUl3v3o8ei0tzCzFuEtFwZhzdnI35HOc0fFJv1uss
TFrYbddIzrI1ad4Yc8SYHinCB5EuYIYzYS+CuimtjvVKKIVJhhXhPJ8ZfQgNAT99
wXj9YYQ2kEoHFA9GK65ot12CSK+UQ4B48MM80sbcxammInkRSjVGW6OML4W1OrDN
Q8BRD0eFZoYCL0xZTAxA59Rq9RRR0pyGkg6SSmnI+a2cTEEg+FKNBN3JEKrDZSI0
tTHwulfZkTqSMSC+nFgm5geYgkyAaKcRC4PEyZLTcSSkp/lkNlZjZczzZJfPOrzI
EnXWaB6Uj7LjB45L0d2tv3l6UG4yAmZgXo/TnZILSsSIG6ITsuc8Xh6fbAOBDdO2
khEeA9Fmcp9GQZfbmeX8EC0MRs8tIIrLkq9IztauRrm+GtlLadvGMo56Gkq0IOiX
jWJ3/q3rys/W1kbfNfT8iLwpFUSg8HdcCkge4dEdrkOjJWVGclqjhUoBWyyoc2sr
T86CwkBrF1BNVDUZvC/J6yHK8beZbQpRfd9frmcZmr8UQHQH/5vErt3d5ZAMHOT1
gO3UIuwhX8QbUVHb27nU0tIcD3U4LJj2A8gbB1QBWoKy4lbf6mXMAvl7/koR6e6g
ge3kiv/inv5RpbHtZFaftEg3hhMUg/Ojdg+/cah3tQl1rE91kcYEl1qhWcjG8AMN
FYpdrr5HHaqg0nbYAYRPfTUzRNoM+jbcziFKAAdbbqxBZ+0L0rR4KzLBWxaVGDLH
LA2Vn06+YrCy2+FfcbjPIkV9x3auQC7JfOVnRoEwBTbp4JAfKny+cyoIhaZYJiYs
pSezrJD2YFXTNdSTI6RWCWxgW/GYeuxwJPt/jUUbLptNgM/1pBYa35haG681eOFb
VuWZadqElA6P6yjBmM5Ml2Gxx3Tff3pfUalJj4V/EenUxxtA8nshOt0fAHqAory3
JR/WFAaD9vfPS1Ue7Ie75SWAAqV1Z9sW/tYg37pqqZjTQuPkPMK+/i2LDd/KF1NQ
j+zRyHK+XIpJf9UudQWL5MFMKXs1IRWkZaQfg3BB3Hb8J1gh+SWrs9TDy8OMjNhv
9J+fpVb/tjAzbJO+5dFW9fCgmNYuT4cW+kIWUs8CijuyOW7xztJG9VRDlchJa/fI
tazQHlETmLxNh++pKtfnO7vmwfsHjeZtTqFG5ZkRXUdhu0Kkp9RLHbLqzX0WqUKe
534UCvjPH+X9Ca9FfzV8I9aIF/ntzNbHg7b7PItxWo0Bhi1rVWvkGz1m4BLCZfaw
yLk111mP4C3ov5B5m09cKOSsBKt89noHFzZ5pUcG2RQAqStOhOCfAwiuojGWfIY6
8NteEl13xqdAcPPJnTsYLPuvdkDc17SSVneK6nCrPeJAZB0+987S37JiEYzFQ3Dc
/2qpbkq+PWqjkHPyjKxWLb6OhulZmDqWEh9f9K42rflFOhXOqnrDnyCGjJazBRiR
Rlvf7SkBrq4RuLOVmSolYOqZCEg51PaBoZ3u9p3wh22hZKJdVyYVWlToqLEVJggz
c8XIftiI9oxcN5ICuAv/TMdE1iS74pKVT+TStWuNNYwiCSMR9GliAvz7hnjSaPih
Rui/avKlEhL3+6tfNn6fYqepnBcPR63ksERQXgV46khpco9O/Wyo+JdVZpaqVZA2
u4nCGOkH1ZEc1ouTD+vXdmmqG64TC4bapeA+u9kXWuVdzyuQv3+9oAHW4RIKLrKe
nocyqU5k2mTA15xjPC4zdCSmLFTnL4GU79C478Py+kYwAXQ0Y4l1o+A9IOKiUIsn
hEeyEvJujooqh8MiUBXgCozekDDMirnDt80SCpLOIQMH2hBoJH28M+JOwdXaN3Lf
mvbny9r7PeGuWYsVJioEXrT04NoYFZ5VmGCqVhuK+W+WkCFZffh5S2U+jvbKFPCg
lJ632xjTV8fbLchMJalS5EWZiRQRafhSv4RDfB+fG2lbXTokz5NXVZlMSsX/tr86
8OMUhS4J8KZzzqrr/0UbCW/bMdZtJVCok26LOgH7T9Ry6Bo3ksLORBM1iOn2uv3r
O97OAipR6ia0VbBVC6VIl2RVYw1fHDwz1h3OT+mrIdeiygE7bOoVmoyt4/FBop9S
Z26sArV8ZS6Le2SBNgPC93pnaQgKHPXWS2j/ZOn6z7niQ+beAhmYlzY8VNIoLWy+
/QXCRuyvu27FRN10qnxQkr06fMQagINyqyAjc1hrsa6BgJuXH5ksERv8VLGhYKIE
QQHwKhyypUcetl6SPhBGPi8y7grDRDTOCBSBk5iHG4h3dfdMMhUKQLHqOneXVAdB
Yyh19uVcUsLe0B6OFLKDonJbeEd/3ZYNjbrVraqtJUPxQMdcIhYaz6b8/+BLRGid
OS+9BfZMd6Uvwzn/XNPAFujiQ3/U2JORfKMvbo3N0EL2aUpWiIHyAViMgdDtmTJ8
HxZ2l4AAPHF+c+Kw3t78jv3LqiAlVLfP36JgRSnnsokojxVTG/uA+A8LTaSBEAed
LxQVSqX/6ZCKq+UuAlJxyc+m28dKB00M15rWqvaX58A41GCO0VHG2sz79E7Zfo/H
qghpj2pZO2vX4ickF4thzoYxR3GHPAq2nxGG6JF9SQhXIF6lGCHgnFb/rClLKmWU
Wn4r38zMG5kn3WGOxkbhDhRFuSNa0yll/2+bC6oevVsQC7a448dDyYzgFVjU+rz2
km1w8/VxYF62VkLVQYkuwt8sTPOUZg1hnnDriUiOmVstL7lVs6ATxdFHTjJq8Rna
olu2H2bvdi+HJbXx0McUed/x8drhY6nSOzDxbm+j3QlpKb0Uhhjhz83R+Xr/i3Mp
NjwC6ll8WvVNZW7Vv96PGRkcJ6QJqHP7g4iOc5nsZ9RARpqwEnRoljPoiSV98sqx
7ouhzKMbsAg4DWqrsl1eu0n8Y7sZ3124ZzkTAUUSr3D4TuP//puRKccQd7MNHry3
F7oV6ls2DYmr2nnuSMDaTU8KEQu2+9OFMYDxDzqa3J5azWrNz72QjGF55yf3lq/K
bDvBBlkqcVmZJzcsg8MgwMXVJsAyPpOrHnsGs9hX5v5Iie80krG0gw+vBW9qCJlD
KdG2ne4ZtWXFUDssj/ufTyO5+gjKrhBQg5AR3BA25+I7Pfz5ML6D+LZtoBKMNneG
qpkN7IeguNZM+DbdDc3B4BkJI4KwIBgnvkt4cXmBc9Siu+KIP2cZr866HmPiFTPY
ka4/RzrY5fbub1MUnWqJ/yeJUOyJBdsFP4Kool8XdqXoHJvjMP8rNatYxgLfC3rd
2qOfzmVl4tSlI6z3FUkbhho463lJGjzz/ESF++lNYISGaJpkSxAidP3XqduU8IOy
NWJXThL/o75/LFIbVqqIKRf7Bed7SDz0vN0FhF7RltgCNaN3terX+U4bKpQquckp
UeVuxoq1gfXpjnNurjNteBRNA83ruvUgv8Qtc+j+ug6XZf81smxqXl8ygStgfSOt
V87rXvseSTAC1AdGo+/XppXyp2M+6LI/PUk5HJrvHocUvYeyszWGbzupWgJOCWwQ
QQTY/W/noe7ESmdfc1fsmkqST4KCnGrEiGZoNSqiB8Da4q2i5InzDkN8QraF0vpm
jYcUh4Z7aoIGoO4Nrv1XEa+GIdWpp6+wUTkMUwQ0jbSbRVh+ffRm9+lxLRwWYnbH
5Vf+gAk/s3zSfvVYzYZd3s4lBwGq8nr02HrrlWpYh4vIytAns0Ir4Dg8N6dwppLf
yPZI9oZOWIvHumOft4A9OjJx8Wo76xSejMxce45lvSuoUuy3lj36yUA9eHHGYHB0
XIxstHAVz/OWFgwsgSNJYYo4b13YpIm/VN2grE2kKCjlWgROo1t9xm7vlDsQk27M
fR1CDqXQJaRsjALfi08Di6k1KrM6HKcLhexQKPDdrFp9EZ7uIADKZAetURnMRkVj
L1XzaBs6ZeJuiab67AcDz90v2mvfSeT5hLb4DR7qGdfR9uf9CGTNT3UCs02ur6SK
88uhbvll5cWTUUU1MzJw6DPPKvFjtqD9anXHZhdZXRCrIrPD4JstLwp21YuOLpPO
PNjYUp2a+Jzdec2IJPeuoB4Q9bibIyADT58oioY1oM4FiltCRmO8gdPVXtGTwOyv
3bHfq9yn90KTlkayQ4j+g3nQAsO5j0PGwEhFBc2gv8c0SgR9VVKUpCBfX9GfBgFv
vAVsmofebIs6BQJbW8ELPOWp7TfkPcP01uMdYqY84UZ/xAFsLIPoaTYNzHeAKSq1
aB/NiAXvimIj6Egl6ryqzuRRtg5duZjmi1DC0gbpf+ciC6N/HALuXk5qWpjZKLki
dsj+zlKziSkl4QU23udL0qtJxPWTB2wMavngh7XFAeQnk41A1CiQtqrKX4t2Tpko
WFuvI+S54UnowpHIqY7EjaluAmfE9RJfJCxD33SvCmYNuZr0VlWnxXgASBuhTAJQ
Rw+6AH5r5zNciOyxBefmgcFWYQZPCZ08E34nSQJjAzL2+KdXfIOsK80z9MIxlHZf
ZBIpwDMvAx/YwDzeSiT8OOzSvhalSD3y/QbL60ytPGRimZd4wOg18ipH0erV7UYR
V7co53p8QUpPe5qar+ovIvySVdi5ue2W9bMUyP7RHMema+r74TVa85ZSmpbKrmSi
ZQZ1wjyYdbOJyc15yUJw7TCFt04qCga8sy95FPl/jHoSOcJnMKEOBZYJsROuextX
A+xtq1GiEfncqJY7a0hOY6NzTLDm4taCrR5SU+5Wx8k4jB7soV1Mp8h0Oras6u8d
8N0Y9UXh8F9fwjm5ffH81YnqLbBuogPmlRxs1/R6M5tvKnf1Fr21OdkEmZyKOJAA
sx1sQjH3qPTSfi1i5wfJL5KThHfPNLF1K7znUrfhkQQHI7Il/d9lR9Y7Cpfy90xQ
y6UyVc10UBVPCOPzt9zciw+JRL7oO81O5xThVaKsJAi6/zzsn2/YpUdQRTfuWaEN
/wgcsG3E6Ly+K4hqZ2Rfa7pjqC/kdcM/wHk6wNEbJfPxskHAFCyQwQHDQ3jADsNF
Tsh18Mha+USzpMhuUNABcPrrMeoYnbj9vhPBbWE/hgkq1No1iGx6n7MzlQFrTg3U
oFt2YTaeDPnNUdov3d25lt6IHRKzpmDVxm50hDMDxBWCih04OtszsO0LfYxAyxFA
7bhzzrxz/f29rQFwoV2G0ZmA3P6m5nQ+6EfgT/f2RJjpJuezN7kbIu6rWIFpyE2z
EiWPOTJn7EQVPGltpdx1pxVS7IwQVtiVW+Ush9My3jZJxMh4O86mbc/HNrX7MoxS
iKbmHXzeLdQuNXiWtEw1navyvramPGWWETzmA8m2eqN/UWuFcqeoj4UhQIXW2JWc
WtVGsTZ0loBY6b1hMVAstlqAd4w5/Mv4LBtefwpiFbAr7L0L0EZKkLc+HwAXuFEO
Vo/8+6r7rmdMUiH6Tm2iNKQQfvKRJgN5+T5uabdDcXTDkaSKlaXVC43+4cOqNsyA
uY8Uyn0hZWljc8BwKPTyiLHj57gIE9KdCyNX2ypfTMm3Q8WVmcZZtTswB4JnECEw
RbxXHdF8d9TZLK52GIHiMQYnZXDvG27ZAsdyTV3atJORvbGgaCVsjgNwlyl8abRb
56+UTOENygZySm9es+IFr7vued5K+1l8MDksWnfMFI9HyR6qKNWGPtsHKlGChuoE
Pmgj+UoRHuCciCO0MwnNqi6nVmW5MKOI9OoT0TR7N5x0tNlo8xaZ/Pt1UVpawtcv
xDegHHZlK7B72baRHTUSCeBhAy8DRlZOvpQgTa2mbJiWx0KNVjU9+/qCXM8gKsn+
WY7Bbp1Gc/Y/TNFurArfaVLYVCHZbijs7DdpvwrZxIbFg2MpRdiqRhGhCicHO07X
kbLY7yL57wS6ZuaNkP1DAljMt1qzcf1Qz6a7nctzQvkCUmP19uBY5jmB+na9mFxl
POwrZvI8gEg0P3u8IypKMO8KQA8wA3lZIFFfOvTN3QahVS5n8h2ctSPLnK0q/SUg
N2H2HOH7wfuFjx72aKRV+AztPUeQ35Nar4oy/StEhxghNgwqzFtbh0qjsUlmOur5
7E7UUlB4ulC8bTF18sz8Er8wVnRGBhtoM66da/jGOOSIsiRs5g0O4bEjK1mxrUul
U4cefxGJj8ZtqTHOTT1bslO8mqNC9zkYAzZfLEo9Lf6YS9dHm4jQartpLcI59tIK
QmEcXU1A6N0gJ1zZ9A2bhsMHyoLsqbuomsVN1a/SoX2AXmQT0Rcn3omvnIhVSMu9
tOUlRqsENe7fgCZDxKjgOC2Qac2TSMl0grFLuEKeG2U9cMib/de6yPRIdnHuXc7n
RgWRFRnVeDmaQmZVL1dAt93j0t6MIKY2EjiPg2fyCDjj8DnBGZOq7EGorhg1Ryt1
LwvEZ69Y/ezr9M/pHeTJl310xMCmTP71DgIoolNPhw4FPONqLaT2BuQT8feTbDNg
J/Lv9hs3xbpV2Cg4fGe/bGYTfMqbBaZe6PZKOnmLbz4qD3kul3QOpNxF0GtWKydb
qiZIgIN/Wgsx/rqiz5XJ+qQuj6r9JbiBhcux8pdsqgHvpCNDtcUjJCrkKARBEe83
Q3PyIB8diLRXcu8UeyDrqnl+jbhFlSBaB/WXJcfhHn3GiuBW9VEAg2UcORhSg/Wk
6eCz0oGCAZbHB989G11OblZSasZyurht8XuUXn1ZclUEiHf3DhS+nLpqG23vWD14
5uPPhCj9zwR2roYL/Fv1sNSqBE+3jCP+ajtJEaXDJSSc6Q0TKCg7xzCwwJVnjKjR
lWvmoiOPXHrzKJloraZHvV0HolEFZFRr+7sA8Zbulqc7Gz+02w97vPltfsBbNpf4
GvdK/MO5aOdqGHAmQ2b9cgyMlicWveTcbJjuJOahrMv8a5bqXHmXeoOBe7wV6+rQ
WbVMBdYVfuiy/uALkQ5thV+G1Dxx1cCQu3zFuKxIO74FUlK39E2HesgxV6qEwcV4
xZtHJ8irV7ALBiTEyMpAVWFoGqHoIxVRHUuuP9Gg8+egPqMno4gCd8ea67TT3Zk5
+x/2rS6fdSS+x9WG2t1pPz3Z2l2R0WQXOfVnY7f9AnDOdJymQ5wsGk4ghzew/AUh
0g0WkO6l+0Gk9Tf5LqzoQSfx9xz1tpy4AVuMwGDUNpYh7DQ6LjVMycoyKbTfIJAo
R/2iv1XCqtS8GnfXudTpQcASCWR76utHwh/CnI5U0qfeBHTVKdtHOzlxVrUNm1GD
Cvs7x67WBPv935pedUyi4biH3EYUzKH+9yExmH6owuCQ+i1TbSFyNIzT90Xz2OPY
ilp/0l4G8GEMonoa+FdYKVI6N7hccghXXZs0L9wHnpdnHJ87ev/LLpr2ZbvnoRh1
ggKt9PwosODN1iuPqE9WiBDwUIWl1p0RJ5efBAFiLcBQN7QrqPh14nPrVeBq51pU
xxMLZQ5S+EmoVaWyHNOqf3jJCXQG2JNaq3TUwq3ietxQmvACRTJvnxMUAPiuQksB
YjLqTxnSfKYbOG7ZBXc4zjDCfMNF699ZZ06cDtlTechXM9LxjoZJu6vhM9GUhfOO
xnxU6d9U03nxR668w/ODM0kKE8rKpWTtQ7cmYZm/Pn18YRrhtETKrL0WCkP4eIE8
153JODZq4M1Lb1tHKxbttZHik5pOznJYPKHz4cXEaHCuXT0SKIn+6DS6Q996btpc
CzjSx0OZ3qSDyyKknj0as7MbIbq8kVPE628Z3qMSp+/lc9Lfos3q5vf9Y6gCyWrl
DBupQOTC/TwoKGLuMNJDupVbPp1Cvaluf8dWUpQHrRcg+b0Mk1A4/+pQp9gqGORi
w2hTZ9cxB8FbJ2+Psnk8qTyJ414/AlhdQrKcz2ArpF/lqioXN1VIKDGtK3REYncB
+evjkG0vpjih0crfXC7fB5T/MW/oJc39Lu8yCiBf2sEKTErzHyQKEjH1oifhuXVp
18gHgIFbxPR5k37UOdYkwNi74zkXoqT5y/vI4YftECqnagz1K5lZgzIOGTGnwVfX
DEqNVABtoFEr/haZ41Bk/BBPUaYzOsCcBEvupmWTJr+fhEDHVUVr+kdOAM6MIMFa
aaYllPdZUakmFKUW6XqJtdDRuKsxrUTiOOBPNccFbkb/5c+a6qs6TVpvGtiXtMnJ
ULr6Xd4y0ep5lDjR5gySLZ0Nv8HCN6zLOgLGpYzOTsu6SpiFOAYdSCy8Fv658O4G
lSG/w0iGHt+k7Y8RkRECxQ8KPW7OAc1uO1C0fT7rNEwrCSyYyRvlmcw+5Sq9gs1u
9p+9gmlct7U+nG1RaR+FIJqFr8AsSgboFaWW2Y52LILR8lKFhEbE/tKP0BC7dgPv
7MihLb5eWupgc2wMouE4qkcl9vnTBvPSck1/thKN7WSmFFqvmT+cuJZaq05kB20C
ZBxQ2ecUItgmwaNNv+b2/a1PZqtyX5h0ZCHOmTnzuEL7L7GQ1tjo4OQ1sItMlhnD
bIQUzC1SJF1wjeZIMsuTXE54zbJmLOv6Xltv5wMsrMSihXPcxdfC53U+sP5mM2Ae
vkY8uymACxUJ22Gf5GuboZ7MAf4dSHLvJPj89+RP2hLjw8lh+Xs3uXYobkty5kuP
BSXE2ge7zghnWUb4n7kMQMXvuj5HoBZCkXAA8tWHjJhBv/YsmYydwqeHCOaz4xiP
MihjzRVU4gkAWHm7hWWOcUkzlZJF4GDkD9YGPkcG+ckh/rRbKZrE1RuSWQP8iM9v
5se6IvAaodfplUmPyKm7OHhAyYV1WVU1WPgEqXHYgIpq9iPRKgMTMn9yKDV/wOic
dQKwgytAcshAdv6gDNENWLAP9SMvL6+eo2Exxl0Ssmzp7E1ZVhTuqhZ9Nw3SuWR/
xVQGG7MC9RluntXgm6VYXs1GhUpidoFw4a6XFmuY6L69M9fLlWoBb5bCg/LOEQlK
7tTKgB13qZJfsW/rY+0WsH+BLfLAnZ2SBqWO/MZxd4Rv7/bFhmNavM0t6gIeXnq5
OobhdHaCzbYevbXkckyz5C+v7MlmpPSD8qwrBekc+Iayuq2bNvnzD1GVQywCKcCl
IzGapD+0w+DBJv19P7Q4xxJgxJxv85HsNZdNQ/tehSTo/Z75K1BcUqFe8pIhwOf0
XMfVsVxAVNanqB75DKtbGk4ax+OmRBk1f2RhvgZZRO47fxJbA0hUcowKRMl0ZmxE
0JzQ3VwZbNeDzNr6ag45ba20FSqHYP7zh/hMN8RLKzZO7/eyq4ej1YnL9xah/tud
cDI+cQgpso5ZkceENhS69ilrxddTlOaA/22OyWbTi8a3n4g83eps3R8VXtkmr0Tq
LF8b3mOb2WcHLtTmdTgMRH30hsy3pUfHbxNk0mhKgH7D6E6B+XzBrnPzTLmY5xNA
kKtNMjUpBLG0PbSNOocDLXjsPfNUDNzv+arrXf4aFjE08dVt/vpXpGTwIe9ITkCY
anyvjdRapAUHJsmSatDlYPjDMwz6S8rOVyf3EyoSFv4i2oTD7u0xvv24lGz92byI
HwW0rQ7g9Il08zAppO1Gs/nImEOCKc4NvvgISCE4K52thSW8+7u+KdI3F05U22Hz
RgJM89+5i1gtYRV4vBBN18SH9KWaHltR0/rppkGMVRz8GOa1vtrSRkH4r/VVwsJ3
7RDfCC4RRMXOVZjZeA4Hh8iiMj4AgwSlKPrCGQ+rUL8BhszztApr1TRQ25wi4gIh
FkfBoqrwLi596ICPbnR59lbRVdpR04S1ZK5nInMK78ZtMPv87trjgzhJCCqempCu
OFfeBphiAzB9ahHsFZvAxUAXF6IavciAbTiOIMvOeoH0eB6Gt3cbUPFvflIOX5Ry
WIpkx/GIV6+qfxtN4lGyjTBMNIeqExPJWUhInEiOzIolBsfcSJ44dzz+HD7oLAKm
9CiQ/OhNP4ZotNQwLp78z8ldHazwq8e9wYc5j4Wy+sou0J2VE1FEo6uj1a/KPFCl
vsD/MvIwXEHGNvz6iuubd3/UdeIpOpc8k1mgj9sL4pBBsHMXl+A4flDks2gyrkU5
Dt4vY94XruVsVk+J8I8NFOpo+P8HaWsxhvcYDqShyteJI0R9oum/x53HjKlLqvrn
MVnn0lAmClYMz8fAclodcIbYccilqcIx4TtFaaqd0+Pn9WxDFIQyXN31vjDdeWGY
dCZOjupy63F/Plt8b7HR6iDS+LWj9EVBNkMt8nMDniBI8bpcDGLEHOCI/TFT8HFM
AHPU356CSiqC4whdHGYooIIZmG3DauYm3ao1OW8yaWZQ6JWSMzoMZTmtzvzFwRSZ
OCElqopved0lgBNCJ1lOQGM2VZzHHGCjUaWEC25sH2aEpF76CStEOIpHM5sv/3Af
P0V+oq/vtp3wZKwvL9ZGKlopTvMlbyrQneKNmfNrbJPZsF/u6lv6cgk8eCisikMw
ZnuDBeTrXts9+lJjTAwDZC3/ok9ef0JJ4aiiNmPCDR5hoc95Cd0ye3ZvXv5H9B1j
ypY5BFydEKV2qa+FZJU47QqIjabSTT5ZzxQlg922/vI/hUtv1h29fvtwI2mHll/S
7w+jI9NscmgEiOqOVjhQoIqfFH7mYrlyvSx4AVhY9z8x9O9dhK7YuEHHFRPFKDJi
2bjzEZAZqhZCgaRArAT+yM64wu1+dBACw71CtcINF1LQLuYgDNSVctlp8O+8j3RY
Vt5dfHAXfCdx7vsY2wP2ocWq3NuD5yF7SRlLNo31vS+Y2BllQ1drT6cR+NW9Jmoj
VHbvJ/cH3jI0yksawYt+qgj/topF6GMkLn9cLdAZObeUKg2uCTxfvlLpAoio8KQu
9LvDskbkzrjPlRePAFjFPEqZYLEu3Rms9LrkwMBRy0M3evNbr4xjJID8GU60GVs2
EyYahzKeLGOPClWpI+/u/s+7vQWDG7PY8QKNJqVokLgD+zt+RSrzbS8A+T3JHaEe
/mcgQga6e1offyC5yRRF4XA3OhEjuqyYNrpI7VvgvH4yIzvUrT1zoceOQWBlp4qG
vmBIK+BysxCTlLhxNnnfwVwDkd47N3/QeTSStpjWHb9HpLDWwa4/tCOt1GP//mJ9
TgfKLTpfXhHVEaSf2zVn2BiFTmKME3gXVM9Ayi2CKSRhwKa0/58RYYFKQ75cBgnX
Z9HTD4LIdaQ7zfrj9mWCKdAm0pXeDCUVlaBEG6x0mp/EfXc25dlWI8yP/3Dyx/9i
KdlrDdXZwM+G01yQtTDL+MmyEL1YKfJGP+OQCBIh9AuUlt1cO8koS9iNjdApx4KW
TYZDfNCUsd0SDxZDB3cru0Y7xQOWnYEfUIjImKtTitJ8GJnQiWvk9BAYsrcW075N
N5x5aj7ETHbLmsdSqF9lCyzKfJoMve/hd+fUePUX2ENEX4sYBU/7d/eJUCgMmWRe
8PWMJ08W9z1VxvxlJxfaIzHA//GYiCwirOL/lXZ3zeKljj7yYDHrIo0YcXA+cTfI
4U3Dnlb6uxQ9zKWf7Xs5GxbgEeEvpW4lgQRdqVoDtu6SJkMp0EevqNjei1FoYL5k
eIynrBxqTQ3BDRjCLSXjzvjhuKGeeikOFA/jBY8TCCrSk7pPowA0p70/ufoKnJHP
RIGUkNFH9AL8vTplxYkYamHdiGKoP/8sAexljAiEHzxUzQrByIu3KnzKjlpmJ1d1
lZyaHuXKfe/Z1uA1Hp34GuFfII7Y4bbRjkeZsfWF6edI5QeSGOasebVfoPoUeh+n
bOJl5EBGuXk349Uom+D7IoFY+p8qjN7nH15PAmuHgyEbUfqMIQzsJQs0+MWcRlxY
zo4mYmUuJCXSuCPeKzSLQSXCXnfRR4hXp9HYq6er1YE4EqATNJWf+8U4cHQDuJrK
s4tGjnBuTPka6WuJJsEWQ4RJrhYAHPkDfhUzu526sfGTzyu5vevrPAU6+tm2Zfss
tskzdLXuV0jMD+1SB+NCqodbSN2Gocbt5HUXBUJCc5YJF7VDL7NxnIAmi5x8moUD
BpLBbURdFTgjWfDOnGaT+v49crvDRpl+hdy70qqog4xA2ukUXTpUku1cdkUpxmw2
hKALXsKKbEho+5qNMtXkvlefvV9KE5H79TTYjbBmtknGhxp7odV4TZZTpSdBzy77
+NRBsnLbjC4Ls7R4ZWfo63n2uPILZzn06EPuoKkQtjZBh2RQNPNvBwYnRAe+XS51
+2snRzhX3AZ0pexoyAY/OeVboHx/30BteqlimKYQaNY6beuyLWipG/ztZoQPMybZ
cM+lGJnFRdzgD8Rba1eLZ63CmMjzSYz8WdcJsjUm7Ky40x9o7PESbm/bA3FqxovG
BSzmd38TvpHn6stRRDVPviNdmWWGjYRr1rt8Rcr7dfbU0M9/VaEIAU6XHj3yHT31
2OK73Rr5AE9bpdEOTcwSTo9sVEem1c4Dw4R7XrNsjKcUBZrUmHzRhVQfN9W29ehm
BmQ+zU+ewpjficNANZZ+ETUGq33uvUDHFQqpUf7X2fLs240kOYgTOsVDLIz8LMIz
xLd59FA1/zHJZm3efcr910A5jh28PDe7+V00aOBxJflVac4mFbg8Zn7d8pjHyF4d
3vVQ1zY8q1IeyTCp/IVGz11T+NORxBLkK8gZZrktcLkRz0Nj0R8/lbgJwREMhXE7
iECiTANzC106iXKlPHM429cJVc8n9TMTwqEbFzZlwjOm1Ozq3UEOXKwr+glvaKf2
OZUV3z2qvWG45EPcq1l5FsUCh3GxnvzqVOMsnL971XDLUbr9fcZBPeHsb1tkPVRN
0Zi59QB+9gFY8872JMvsXtP5DhmtIEUO7UuJsx5nJEF5BvepdT8YhACv4qwgKpuT
TvsqePiHJrUlXvrRQ0TCaFH1aZ/WUKcSAv3lJovpKJA2uvmkAUKKoOHaUL/BQUBT
0KQ0PWwSuaKrUvQ2SwJQKGzfFlPUl2Wo6xhqThLguGq/xlHJxKsLfXGdavb9Com/
bWbBin2Qls53ZA0Tz+4Cf911RN/UnhwETlAyW+mNBxbDsXOR6XpNaeZJKnuxjr7z
4RTvx2RyKhFlVX8dqHpKGfgtX3GLhDZTiLhMhRzupM5+rj003/jVPVqPfW5yhi5w
k6JoCXGV6Og8w7uGTHWPtD072+20eLOYqnyGsS1GICdBkS7YKDPN4JykCYFe7Qae
Vp07cBXvrMY4XUb8TvhN8ZcLIRtsjVwl3pL8Dn8iSfjcK/K/WryFH5BEWeEWVzb3
5S1S9McIVQRDKRqSg3SCSo4Go1n530audxtSnRNryo0w/sg1AvMVSi65sFXcmgZ3
pnVfpTjZMLCXwdFWoOCwZRgUdemFx+Vtxx/Fla5euPcE2j1lR2C+8xiJmudVvzRf
Oq9++cTN6LarR7ZcDtt2KhMGkq7jpZv6/gQmxDL7EhwOLTnlWUYUndYDuj5KULEb
7eSgHrSxxG26r/1FGlu9KGTZPQnIRrN1VM4LaQfwRY4bYyloe//bZi4LLZHYs1El
g1Q0wxLZiFaEVWdwDpJsRjPDhNkfkP0MtZLxQXABl5r6Oq64HpN/JroywQR2j/80
liZT+WFRurNFeMS1WPvst0mvygStXffoks2z4r90KCwoNTV6RUKL05IPa5HYZcU0
lLIX2DjmnR0WVj4awbMAIlVSO0poBV6PlVyWva5kJZwxpLUvXFHx7RsdQEyr+yWd
X9h3LPneo3hFPHxKmRM+AvoADDnCABYSciR/+KZ/IvznmHlj0OWo0awEQPNafOsC
AuR/prd4jqzMl+Ef/XP+4zH/SIQEiir5gw2nny5SK3whmvQJVYpzPV5WMleVktez
xfpLD31K1O8E9X2rP9QI0vI1oVTvQtvEagLC++WJ8IHUpLDXYGgLBlmGobGuam1Q
rzdzne7+7PNB1zOkwH8t/oVs6j2iNYGkAVzo7ehmrWebvEFHeLO2+N2I8cWqwzcJ
wZeBnVG3vq5qpyCQV5x156xzVWbuphb8JsDB04K4OxYwc5q4oqbDsqsVx2WTTC2t
ijVNRIbX5Pp76NsKi5Z0AeOeJ2/BX2vK8kVjIvCvc9lGprHqrOMpLQY9WlqbrIpJ
wOyxWBVzdUkpH369v+NAJBqu+DOinsnPoLmXUe96FNqk9oWBuVh9eRqMv573c7S9
OF/fFIJqvuR41ufvfcYsbxYUx+4yuK2QDwwuPDsbeUKpx9XiUqHJKwTMvMXcRZfr
D0iu929GeyQA2GUpar/jqzSoH7NxVio1WDtxlLUQc4mRi8HkaiHyXMoByrEWN/yp
eLdUJZdcj9KhuCibbRz3ddNrlYT31koHPgrgCbEfx46PV4QndgZV7YizE1ldHLaq
Hi2VoT/Ai8GGAMk2lmWtTZUhVuhCnSwEGSpSYZePMFtGs9JoOjpsdSYLGsrBNtx+
PFCsEiJDP19VMTfdHpu3mYQnMQ1K50DAhDcMSN0j5MwUtYNOHJiMvgr2+lKEgiPB
j+c0+uIEsh8npDRkZexixe8/+LXiw0qAdSe4VRzgCqWcmuR1WQZPTZva4O4WyTqg
h4UzaC3IGesGKjg/fEftl+w/s+Lo+tIdzmTy3907k5g9fuzrQq/ox2/qJz26ss53
yBX5/zzfoBuS/u0fzbabscVw2ujWEzpexhLwW9jgIEvtLj7m8q3hFjDa1QMwt6dZ
xejnCageTZ7LlwIFOMZ/R8Zubdo7flVqX8D+2sJsLvYfAVvDfwMMG4PSAgPJUevQ
SR7ScElOrbH3LE5IQjnSt+3lMKT14WAICfcwFVQJ8sEE7vc2d5zhRYM4dMuc2HHJ
PVue3mdEDqdGAoR8Zb68SBcqYzG6yZ0jZHlnt6GxzSl8R4plGzhbV+BG81Bgc4Mm
VqYFIHkk2UTNkcJy9wvP11dzbNh0YbRIUDwnj4vKrv9ZyhyhEz6Tz1179uZ8a8Dh
y4fSF6o4qIyPLX8QXVYfyIa6U2T3EBf9MKrwM6bIR+sU3dFG4q974TdyfIoMXHnb
4kV0+r45TJqFfaQ05fiFFp1TRWvc9TPTIjL0YR5270dkD9CfRyitK4ibByZkrBEE
TgQ5He1G9/S59Ln2PNPXSP95za40EVY8gvixFuZVvgzsmbs/nS92mW3HI1IqkOVc
UVpPoJNdhlNBtKdKSwM29/Hq29mtXzcDTRSdB7McpnzHYFD6ifTKpwPOXeiScV2n
QsNJWar9YnhlOqN1XLA7Z8wD8KnHF8F3UuuBIs1I10/icIuOOWU5L4BuYqBg/mMf
a1EERux2RGxhXjMN/BtK7NXhvCe3+ivkPOfnP3iF9v2crxTq2CJXBTMEYU7FA6fw
sZOVatNnJFaRqM6nZI1QdNGcrNNB2iM/BprCFzi9My4BIOYXCEAv42ojck0Rzt69
BOdCLx5mSgtjBqhuTht/9sbKwv2LVOxjLpSq88yy5pZOf+XkrXdKSq9pdME/biuT
xYRyASIta5DI6WiegjB8xLij1Bpk1L8ufrxLfmmSDh9VMZlMicxlNfgMH3eVWLt5
YrvoB3FRxYeABlgg7bRJpkXalMe7N4U9xcNyHn8KkUkD7kg4c4CldZl5+FvqyQqU
KPXm7+DH/ZPcadszaA+HbiWuc0GjdfZux53YTLl9jbq25IX7Wc9jsykrclBoSpvu
JlQ7j0ohzrZc7UpXsuBHMyYbsoz+4RmzYx3fwKtTovNz1JL+EBWcNw9aPs3sTxc7
2iyq8AgjzZ3d9Ch7saEOyG+PkVUIlYX/DLcKPj4u+VQW4Ez/sH2Up5ItvVwC1GCr
vd0eI2I/G3nhh5zPMb4bUaw2DvbrWcvUIJSriytKpG5CuXmRADTqP/+NiCRaWr8h
4jhsNwDNapceWrt0qvS9eV1APp0KXoCLF5XAXfYwsF8elBBYeaXLwJpidvEhtcPI
Joe6UgsAmPXy2d+l0AdE045K94zapYE1DEhzTqHRLX/8wX4EWfcUJJPdK3u7LQar
dRsF47yBzO6iEHiaHWx+OgJTlbz5MH8cIwP3gzOyrhMFTyrEbG+xIkpAHA6fHpDq
IPKbCD4tMkfWh+Hwd42RWcZZbIjBD3oOsYd20LPRp5FVYKH80s95tNh98u4ZN7HI
9tsv6Dd4QnyBo4fokCzt/lvTyg9/7fITPcEObd4YX2PB51vU6CEtzMzZg0as122O
UVrVSp+FoavpGItAFe2cy+BtT9m0VnpnkZ5p/tY/Tc67nr6MAIplyTYua02SaeSY
FDnB0eSFbyiENUMnwPR/+X9j3ldShM7O1e709ptlGb/G9mNaliT3/E/Hy71y8y0D
lBrSsGxRmrZ2W1WwO0gMvVsDTlcyOhTnZUULM/Kh0pvmkCxzBy865EXY0e0xQbwg
Z4sn31Bh3xYjz25O3u/wTzDnlwqk9PYnX8KSfAIJwNpz57bjep2LFXXfTpNmQjnI
tsIamSCuB6oC2ooZjpYdrYgv2CJb7PA547ROgCadwS7ZJYRP9QnGQevBDzPb6vDM
BWnbqMQc5R+42v11BNfdJ83usArsNZePuvjdRYaklAYogrAZn4DXpYNjPo0PKXvJ
B1UamshUllYiuP2CxRfwtXvIL32kAPajCsx2adE5bb/OMiiTg6WpTuKw/crIPkz7
2b7CP80Iq+QfgkC/eu6POti9u8ykWqDYpybwswrBZ7ATky+TZ+CAyy39HcQ+EGZU
r21gFbTcgI+wPkOO39Wccdg8kwqyUmLttgw2macX0mtZKr8hvPJuPZ1GzdHWyCm4
zqczFv+eLv+7sZt1LaZP/PZq2HX29qaBJvWMFAqQxpT6SBt6sLjkFKB2QCizs8zR
1aLlwj8PW8JTNQjCYJgaSdoH6nVlxQA7eU9jc84FyRRVEzrMfRWfhZJmG2o//FQg
4D0Vb10yGQcw6jqvF2/kmCdwp1xDakBlOGgjDOX7Oq2xpEhIzsy7552s/yRypZrn
BgIBRdkKCMQOjNaozVs4/hhDqXkAIv6/M/yUl135PWMcZAgt17khGbb+xM3+SXTb
Lrw34za31Ij9v26mvlpD/KKzIraQ1IkZlbxVQ2fao2iSjMi6JFCnN97XVi6rbbX4
/BlqpIXKXzyBKazlkKU+Pcgaoxiwqk+omP8oRS2ztAkINZwfkGlb/Hk+fYneoWGv
Ga4/ms5I+/jRy4hEAa7vbhgZEgnlkW+lE9i/m/VyzMz0w1/58LjLf5LEyOQE5hjl
beDM5m978N5H42NtXKNZWbJVrI7/O6yEfJA32vX3hCG/5ewjArOldvOYeVMZ0iFJ
Z+bRgZhaJB8d9Bd10T6RMG3w6U4lA1ZLQV39tSIXgvtDSrMxSKJzIR8lwaxARakT
KcpBy4XyN3mo1VU13KJ4Pj1THlwqAAxU5D9f8YC9QQ9+SoxUqmTCTjfLpF8NrojM
kmRXyoHdn6S+G5505LdQyni3kJ/sLyv01aHLG+ef2vGMPnI8wgl57VvcWwrqCGx5
R7ztNUmzaMHInYBW8icKGPP2KULTg+D9hr+NzuWrktIVM7tOV6BIpyZI++fwfkzC
Rbc/HHuB0P49Uv7Ul39w4RmVM+JQXpOra0QRAErPeX/Jm+gXaCPU394plLYzCSr7
lh4YnIvhPzFZ6TU7sHXro6eBbInrms4GpoRIX4/8dohl0BfePSTFXiHLv7NDmzza
jognTDrqowlnGP9Y2pEAp/xV2kek9CfbmR3Q9KSsY/snTZTsGDmHYZMEA9S361dM
9JvyMsldp7LSjDkmBsQm0UF4WXBYuJJJNri0zBmM+yliOEx9YXRJy4mG/D3S/15N
6mUFV9oK0JrpN3FS1FtWwXPea+VxtBgVzBv5NYQfVDJfIriT7KxGxSwKojHA8jwq
AEZe9MKcV5viGNbJjIChO/qzmfetKdjUotbFplhmJDu7KuY8UT6e4+ky10Q+G57h
z4uuPUcpMV7NtUsXoItX8OXT0/2yi2HJjnSqvJ1gqdfpR1wSTcSlxTUGYvXwCbX/
Wrnf9LlD7GUWo6VROD7wvyPg80wLLTh5I+RHN6XQK+d37MecvJciTyOsmxDXsrrq
+cDEye9OrI8vkJ691CwU61QQxNP/hXSxVhws46v0yDFrgpzmDTS6o/13XPiiQQ9/
etfjIxhAnoEvmxsxX94aQbnaQpseqGHGJDKLE5K/FBfvLCqtSPPHPppm7cuA6ytM
rFVJG6qLVm+9OJgelirAmVkmQiKQEIbGR9e1ZC5tkOVMWawx2wxNzCXWmtVU4M6s
vIL/+L9eT7K0ej03EEYL2wuOVl2/wdDg81qxMpOMoeemIaDfHvKIHwWvpU1WZAXC
jXkabo0optD8PxfjRmFmdB4QHnWPv/g7vxICgQS3AbHdRk3BFzh0JEiBAMznoOwh
9aU5T/F499cNc4d3Nf2US3MhGLlgFcLceE49nywbzUUW4tO0JghKhMJCnSoCxkrA
SWjA1uov6OvumpxaNG8sS4XPi2AchlpuW6m7cbw50vJMwn3AlAayPc+a6Lza4fZ/
D/TACFTvoRKoYnGHX5qqAAliBTHJB2oSNY+Mb7/pvlzK/osg7i6W/x8utm6yka7N
18k/xk/BjBmea7+BAq1Ro3AKArauol3VofcHgHDV5SjB4jSkSy5/KTVCY8p0Arlz
R69aevPGUvoItbrLbY+WzkzhtinjFWJCcHHKPktGJiVKAHhpwRJPEq/XJwDGEhEM
kD3Ji64TprLHNwH8Tpq/zkyfgZoWq6TcEAaVhrudiGrkBkb7bLmJBYnsl0bSPH8O
mRaskJ9hNtYmUA6JF1jr4HvSZypTC5UVo0IHkXmnqF3hUGmVL5482VZBNX487m+c
sTmZKN+p+KBPKGeQZ4twmSCgF+NHGfpykAwtz49iL5rFbwDsasKgQDty/0Tw+A1B
TNeclStqlPywa0TM+a/DpDLYhnbF3LKpRYOaxDwwMGL1ZtW4rTKr/n6PHPX3GM63
d4fn4VXmWNoTuw0ZM5OCvSOB3IothKhV1y/9cG5RqbqnsaSc/0EPpeL9iFJYVPBp
2fR/1OGpwQjDhOlpmnCGY4Nxa9NFO9dMSe90kj/6lGxhc6piyhk7GUiDY/Nde+nT
FXa/ilVq25d95N6GweOBtVYtiiD4NrfCmQYKGuJslQ1Y9RhCwU7Eqvak5aoCTx5z
K7amUghB10Iy6RC8zi4vkduXHfAidcvws5+x4s4q7e/ciGiri+WgdID96eNAf3ST
pOvCp9fcb9Dh9sFhtyg4Qz81hdc1enbpETza1xJq4rXNLJZhK2JGszC47dr0UkYm
omktHXv/NhukoW4EBV/UwdlTXjoe1E7J7lDRS2VyPef0ohW11K6qfrN5QAp1Bogi
URuLSheueikS32LdcAf/cS6I5FwZiKEktwhIDuzL+Z58T4P0pvdOiNf0n1iaz/OF
4sZEwupN5tFgef43Cswsjt5NKeNt5bI0PvHSMaB4LNFyk1gcfDXE+KwJ90OlLdgU
dQlfsixRVHmKdUnQZM0E4dI4FjklYWijaGgs14wzKI1lUbYm8h+4NPUgnbXW0Uol
wM6myfZwLACyyyBwVj0QU3k7we+7u0HEOVF8zgfIE+z92iNuGcS2U5N7IeONhfsV
TxU2bSO/Rs+lWZZ6KtcTtaYh6xwKTjMPrG1SFJsREnFkrOCZOWqINloXJdVTXeVj
eLWhB3utyq6ucqqxSYoqvdWdkWJHIsBOpVkr16743Q4YbywptnhgromvETrTEkDB
7D91qokuSzladQsjpjpL+VVL54/uypeecr3/jdJ0C/4YwjZ5+FfQyNy3LsQBq428
pg01nhUUD3/GiCtsL1uInOsjJbsQY38elc0d8cnRpaZXC7kZvMrGV9hBc++vbh2p
XbP5mo+BTTUkkWGImgdFhUZht7fiLJ4v8E90Tu/zH8YNjV4jOfQhFr2ldVI3y4M9
EXIjSaZXxK0kxUJ+utg5SH6JPVlG+JwA0Ui22ZiShd/yu4r0P+hg9Fq0H9BhOrHN
KP7uM//vbyi2v68Wj+fQhWpwTJ6qzaZTdwAiFkhxfvcEBBh3w8ALWPvf738HBlQK
ApwBZGDTSpc5RgtOKIGU2f0IQHXzPSPTpEy/F1IASQhGv5SDVONu+Du0sgYNnq/w
xc3fFidXGuwd/5BYSGe1sud2MN7kNQYOT8bltF8At8AuY3ARsrTQqxMExJ9PoVG4
YLq5tFmmLycapsLwS/556ahB/9bIrGoYeXcmvMp3mjqW0KSf0Lq1uyZGIPgjwlAc
R56z3G81kaiQRk40wFOyJmmspaoP4o3TatMYblf0AqbEV17AfWi1W8VdHWBM7Ilx
Bo4R+cDUtcbaJV+OmCrY5zWoZrLlMbUfjrpkGYl8z5xcCf1bijCWu77eTXzsVSaX
wMIiePT4ilF2aL9NnJ1vseaanbgBVuV8+8zwwdBUNakQXyOkDcQh1zOTOb+N5SBj
RLY+i3W2u/UmKNQQK8XVFvZNNEBDJB2kj0ALKaYSW/ASOXbw78E1fy7tcjhvPo/y
u6i2kYBZQTdtV9YHIDAgWbZhEXSehvb6NOErKZoov2F8lfLwBrQR7jYuNPwZ52ul
ZiQcPwsnES/RnJzJCJcjU/6z1JZqXGvrnCAP1h6GoQQChNbjBIF6Mbe0vS6ZDubU
xHVZORMXc5CGGY4BpaULA3Pdgp+mQsYzkMjKJqu4emiN/jr98IlBW+wFvA2ndHxh
DB+qCqnVMdPzN8faxLKyKUYVSPpyAlkmGZ7yP3hPsOSTt35xnSukPa7zyIba3Ipy
qCaGaqiFszS5XIAq6pJEvbyaon0jJ5bIHFjHxD8+s+6RNklpyOVloq+0Z8s9ygXL
tg5jxcmyr0Y08PoDmn11T7sZ3RutUIj252c+YVuYCR+5r1OWGx2xDzYjLQ1QkOla
lIL4qfZWAWqIhVDQ41kB9kEADEnx5LShGta3X7ZX4Jvxrf4ypVT89ScEl2Zqolyf
YSQCsPE7k6+WFBUcqEb1Y72lqlL69B3gOZYdTGR3jpQF6K3dpFRMKcTlcu86EY+y
i5mJbtkXGNMf3TowL9s8/FeGdvPxUvcpbkM/M2Gajlw2FTp0LMcrgA74PNxeiIcj
pTvl6L650ye9JhjEM8ckrzpVMSbgraQqq3SUsBsIobgKgvi0otVFOOfy/MEXqeve
XIqpdli6bnPoQQpo1/S1EgTZWlJCIeq5ZOv2mayTrwFZaiXYpFXerdN6Ca3KQAbL
n0rE79HD0K8bI5fmiqe+NAkTyqN+gYpFAhsaaKHBim7b3pNei6QFr6XVjSaiTUS4
9HD6rotMvU0BFpJg50xPd8Sqm96WoYHQRchxHnUgJekYDrudxsjOpZHoBAaYeMgG
Yu3D4cVECtZ1JEy80XocI+1jxkovYZaFhJoXchxBKAoaTP/vYhZBrHyzZ2x8maLz
PXKPa5yL+io6gOW4SxgaXjA3ghBSiQJQ+wGIoXQiLrSCyyX7ooDdUnRRRGbF+ydr
U3QdasD1fgr2n2+ACj58CarM/FEseKgF5Rf9Y3kxE2nhXrwQSks3NjJe6LySPNbs
TX2B4WjxWvGRZU60pktu0zWKbpNZfUCxnH5Xllq4+SkDb5m8MxeL/fpeSZ/+5cMu
4TAlIkCqSao3A9Kz7xyhKPLo3QsN9+7H53i1AnNXgzU0i1dXEeEWeHnJOiK4JDmd
5S0b0pWeOuxkDlaHT/mccp3LdDN6r/TLRC77zoGpkwuPUlnk/+OdFyKUsyGQLmFu
Bmdk2oU10nvf468m24ijli/NZLKTrOryNIXu6+D9+ulEwW0ZNJFjOmZ6ZlFAzWjR
lhQERIyYz+o7h1VqImDw6WqUi7tkbJZ5dkXxzNyoYG29L19uoiBuIkueha8tzliF
zK0k8KXKqfd6fMNlamgSxzH1DWT2m1rc9/pS8rPXPVH0pF9Q46TTPXCnPvU7DJ6Z
5/t9qgltvTDLsV6cZNbI6MYLd0tY54teE/6yfNY5OAfYRdk1ldvu2jbYS+3uJT3K
DQtHvSh9v7OYuMYAGsUybYsY6JvS7wKMHTpysMCRAakqCU81ADeL69TWCPQU2/Nh
ZYYyVrO15AxEd3Q6I9TNoQcud+s9MUXVXWtKpQlxUzV/yXDPkYJZvU0xgB8HPg6X
F6kNPC85ygnAuwbO1efDYan/MUtuMChHCKZdFqPsa7qTaN4hmnc4Y8KtKONMmYfx
7IYuASmdpZvWQf3U+NqR5oGkgFPVozVQysh3f/EsUjmA17JN50Y2RbTp2+HMNikC
MDkIlCOCsoIDlVwN2j6zh3pzq+aY2Jxf9BIw8b9rxv4wsTiMQPB7UDM+FdPPrmi3
WSr7YYk4lUAkJQQp6dXjMDh/q/jl0q6T7INxVSc+Ibvsx916tWHsVCmDt5+x68Bx
1BbXitaScDKFDudnwwMpVrDMxaF4AIPjTQPHx4USKyjC40pR7b/v2ykaxlJcsykV
EtAYVBur2umvZG90NyGCyKIq70vEzS6ae3UJVMY4BkeGRA4la6b+hLuaMDpPzfRT
J4d4UgTdKdH4yR0SI8Yj4VhJvaGNxuz8sg/IYNsVR79bb6kGXeghzQLRXa5KQlLB
ehQxGw0+6Yz/MHlLzP41GCmVn6iHzO13WzQcAlkyZUj1eR6sZb0XzRkqjL1xJK8C
v7kBERIV2bjmbdFvVJiUX9kK/6k4xbTYi0xEffwmOHzK585C/sTSZCRMZXB2h2Jo
1GoI2Xv/dJVe08lD1+uMgjY6g/vJ8oL0HDBMfPFv5nK/LnlWd5UJdVPCqVcb38au
KapRXLSoPo2zbCoSiTnQi1uyDlk9TDH7naO7O9ztDFY1aYAwYOZYI0LwunFqSV13
zPpYU7ljgPD1hbuaTo2RDb+FO77e7OnGnxjvqz7ibTY4ClPrZHiP4p8X2VJuW02o
bBRcAJns8jYalid1ZyD9q+2nGHYGA3gtff4obQCqCoSpgRk3IE6YKb1IR1DCMg4x
aPOOByC9cz8GrnqvN5LmD3ggHVBoy0zao6CY1PQFJkYmY6p6CwtuQ8rZ39bsi+s6
rM+mfc8++AUCrM2C/dVchNVYQmEnpRQPUaLWfsquUgODoXRRGrC7thkC5lCJ04g2
nvVlQzhsue3PVaelSB3L21WFD+ISLSTjybTMVRPXhYxBAsooDqFNH1LQFrlQuzyN
3Aq6JOoQ7e5/KHgqAMQ2ToCLXA+ixxCjC38hzNLoP/mRBR1sZgadz+I1eQt+3hED
qjlR74h7k2vN5AGw8nJCp/Li91s9Yahp9/AIjNm1Epg0ljffI30PbXUISa37xFRU
ZaFJHPewoGSnXz6JIO2lNIvK2x7XlrHraug7od+QWpdRg7kRCQ6KTmF2gfrvFMl2
ZmBC6wqHX6d+j/0EhZVI1s4GZ81ZCwQVGAH6kDvSEVO0hAGoyRpTabgpmp7LZRCY
0MS+BIonAwZ4jf/cZPIiorq4xb/Z/s3mZ8TbJj2jWSSB4wDf+1mxMI7cZQx187Aq
BKY3Chj4qCiz1meap5Ra7VdfPViK7au1bB5CfiluHVvcJ5cipMaMXobdrGzy9GI8
WA+O6QD9MCoQ6rrLUW72Cb+JU/lOsSfn8865D3efSMQI6pOlA21lAYa5KLKhz4xz
k0jzf0/bsOndMI/wktMKZNltv7Y0r2Wfii2sMpTNP1n4POBUCX9COeb0Lnklwfv3
N17+SQj7ZgrdfJgDbPWDEQ3wTdPLX3/ECLfuQtdIjTUHNETPUVnfxe7dMRad3eOy
puNGIQw+z6BvQTFMhMb8oL8QkAayZ1WhFDMoNj/BfFStzsdVSA74x7dlmoXw8WMv
B+O6gva7C4p9Mwfg202LY5Ox7FZ5DQNbRh9LvKtqvUnrO+zsZATfq+fNbflj1kqm
wtZg5iXbvYN/OavQk8PTV9We4jYh/dRKGxlxH/CD4VdfxkccAEc9Z8XhN5vj1AE1
XEZzfXNCVVtXMwVD65aPvdDOdJ0/BXTiVF+1UZ8zhKVkZFQwK470nukQyknvy7KB
HEAKRZUsZdzKieJdkV2rKuQ8TJYpuFGNvhvODi4EJQUmxo5JTxAviEGDln2Ry7WY
qqbJRoJFaoZTKh700wA17tHBqzR24YNXTQr0MO22y0YTRrwRXVsVIzcR7F69DoWe
otPU2V89Ew3ZLqGndInkGs7X5KDeje/NpLwum21odIEiZVbMRACJMD9zP5epZjBF
ZynholVa1P7pENXFVLngoXoymC6PuLJfdsnbUBJUqRYzlMP8dQSfuElj5FZaYqQG
beo47JvZQKSGP9cgfw/MSdAPCO+F63zxl2ItToDZHbUg6JwmCIbHQN8DuRjKZrBD
raDINsD0/gARwVpNlsKU3IYauRpMugir19oTY9SsmuBIj5Si53ZgSwPhON3HRTHt
GffxK7mW9jaZxv94dRSveESMj2wYEM1lr/fUxQVv8sY/05JujtaGMx9h+a3Oda16
uGR/FKCfzPTYb0uZRNITTGPK0kqUBD2z6YGHUVHJcFFPuk8BrWUWKHQdSX7innib
UPWhZGn/L7r65gVhlDQA0lRL3pp1QYE97zQyp9Qx0OVZ4mU0IdugSI0CLOlRDnCl
YycidPmPzuOzb+EEt89QqJGRjiVN2XjxS7cIxXRhegm0lmqn0AnM6qb/Nk5g1arT
KFB8Wt5oAc5sz2zxLJy02TbaIM18HPkHbAeuXaa0fjNiwIJIpYh487ndrFNfIjUF
R/HjVr2JGKmcVhkm9xTs/VPCaA4WEd/AhUpQSq07MMYFj/m19oVKhj4grI+ASxB4
T46u/oiK9TZ5Ad3C5BRuv7EOk21YJhIf1pi0484CHs6o9SUhBQ48DScoQjGcdJoy
n3FNHyG58GQoNU6kNt2cjbEDV+gU1TRzx9iPHMJodBlWcUoJNR3yW2UdUFIsegxD
wigruxXYbLyMvRlyf4WLPJnYA3WnVx0GNGBCQKcF0Dc0ghH39bwyxm4/8FObfdJ6
v7F5gqGgZ2ssIIx8pP1K1hx25mzIJDdC82TiVoB645JMl/LYGRgc4oLsq2CMLJLX
94fAMHgZYo9WfuoFWiLLhSjakqpgGY7MkvMgMnJPuV4D5IfM8kTbAc9BD6NW4QEh
Tk4zX7Etv/xogo8Jf3M3w/YnCHO5hQi+5TzgkYisNRMX98CKZCa9nOvppHYcdM1t
ypYz6JZL0TjtrXkkgN0T91XQXLt1M3wOQ7KmbswyCopGeG5PNsVeiM/hq4+UJWmU
g8gPRzgg/b4EkC55Z2tts1vRxTz1fCveLlfBDwONc+pO9znyrOJbPaLvM9URHSPG
MHCRdh7+8CkNjqicTJCW/HJm875So4X4I4n61yygDBRVPeiDerutvxo8Q2H/vUFS
brUQlkPoMSOLPZDQWCDAJ4qZCUMLHuWHcj9v+y7kfPnFtP5n4C+6GKomCfh2pT/h
ooIoSZHHEEFQONFKM1i98A/+AKAPJhzFG5iGVvITYEqYXg/Ub4wXntWUyqTOd793
rRs0HfVKUeqDqCxIh518qV8AcUKl0j/5j7Bz6gJg/j427i0kl1cU2kuUc8VJyp+h
QfhtToZOzJKdrlO+vCEEM/Fo3G1IDEKieF2GcMN/UPblOKPQmAa6jNLwME9zT2Pb
ZsNjXDcodjI0KERkQv45v1OZGda98+AxBf+JBy4DaAXwEjYj1d9Ru+uW5NOfzGad
uOfeOSSqixCJ8bfU7lLjJXPlCMRIoFHTNF5Ml/fqEp5WfVJTPzXRmqzPQmnz0U8s
Y0G/2n7oVuvi59pFJZ3yFIlOdMn4WpmJw83hTlynpxzQmVS8UivEVlbbzVNI4iSH
ka613OVZ1ICE9swIw6Ot3yukK0HwcGWifIOAqyg/28ntEdMWHrWFLG3WJf6mPht+
ojJmY1vDy52n3GAoXwmQ0olmp/tdFyuy8Asj4NL4lXb1PAmQKSo5l6VlrW3ZmYB8
egL4b6AHTcRrng5Sy9k9/tLH7HVZFsRU8uMqtFVzpziTL174ud8NHN3ViN5jYZ0F
gJFeQiUQESaHUyYpd0JNTnjIOEheBAOKMpKdA6ETmuFUSTfWd0k2xOsNhmhv07MC
OW4P4O6Lxv7mN4Qat83MdzMpiDPWVk6Jv1w7f2LNXy5lz2MioOz86ocrEs2GT9Es
y1ShmpV3fyPdLW3HE8QXPnHla+VkJ787jUR6/38D0Pw7CK52be8llRPyWotcpJM+
MuV/AertwVB9XnQCVxT7ahqXCn4vzLkdOPeJbO4KKN9wtQp95tdkyum5zXBkWScs
EFQR5IwgP5FFJC3hsauu5gTEOBd7i6fkU2gFxnNSZ3obwR3kDLUekdM96Yn4a/cp
U8srDOgTtSZmnFZYhgW1Rv/xxJMR/HWb5vGOJVDkihWffrf0oGasBr+5NIeXPRGh
3y49yd4iUMNrqmOIMdXuoDZUxpNqLacY7zggx1tyK6w11kvCz2Wav/y3cr4q85+3
4aTZZo5+5YshNSPW3J+12D7b0OACbh19sYnFVVdkIDbu3pc1MHFB+bcVsFP6N5Wb
ufGYfkTJlE2ECWpllukESmQKX5pneL7446j5EVANeRszti6H2VW8iYVq2JgmL05F
Ly4wQBI/MaOcO3cSxnPgG4z+9hm4lVu0zcl1DwwgHBYnHqMF7Pp0Cpgf+iPtP57s
tSMSyZMyZSnV2BJGYOHsGYDf6arzwp8IUzXPD7vzurVT9VumYCe9a+WacthQybhF
3Mb4IwpVv8cPJKKexI1yqrXx7839+EWEUiIL8ybzKnbkbpKUSMgetuQ7BAlZvASJ
bmTR0aYZG08+w+MrsXDUPINa/c9wMtO7xYDnFBh6/j1O3k7Ar9pWozTAgAY4si2q
YXxP5fUV+X2FcHtk+cvTWJCk3nMw5M4ILBwJNNRGKLCyKKm66/O6jQ/eeATxjejs
p6vANEwqOSCeYHnM1bwOkXt58OQ3lLcGiXHU5aQm3FC5ogXbjpE87yrv27ivyd9V
wG2EPydtWq/R/M4c3vU6jXld0JauJ6MuvpERf/pmeI+98g8NpS8wcKgUfEJ3cbCJ
eNUBuzm2R4sayzhjGVQ+yKRFq8iXv1VEcqFNlECZ6ZJ6SAS81FW/3oxpmZJ06vm5
MOxvcs7QzhWA5fwNIwREqAKyuX7kHUskgL8I0gil3DWuXame0ONnUknLvPTLJxU3
ilvixIjhsDzOIaZdq0/oX7XgGqniuV5Y+5e7U4sMqvxbYImZA6paAjdyVEjvyXlO
Y64L7dUuVUOEk7gJptBuHUZzR9+8NLAJeKkuRaPMWFptEmHCfhrookg5If6bbApS
FzRdZDiAHHJaiSu4ORL8KusBdFcjVtnGUplPN3LctGatXzTFLd3XHcmr8nf6lnfc
w5jQ2OPgYhJyLRf5R8WyvoNrFixkcBj0qepSvu9C1hhZ4pigqjMLP1iNZa6zTtqC
0DDpcUOkRcdBfrKJpiNSsDsAASf1YiYHsdhKS5H1FsWMMTfVaVYgtzJOHTMuLO50
R0OMC1yEAs7MTv4h28KwTBAsglPTQHqfQzcLKrjqjHP5Y7iUVQop5tZq+oirR6rd
EuPxyAxY/QtzQQxUtps2LZDj9zk06qIP2hrQjO++VSmNdKYyKrUWLcIoqkw5AMu3
w+is8neF2HouYR0cBHT9MnE+YKW2K8vR2nQzhpQ9t0fsHqWibeBgGHw+teZeNkaw
Xygu+0+SM33Tv7cLkdydD9yhueHOJxEEvHTfeX+AoxZ5g5YO5X9PsRigFv9rOb9k
nz++3QHRkqKIw2Vw+rbUbCM6tLDvpbm0yTOK8PBPYfjljBRmbJ7uXppYtGhGMHMz
MID8uYGPzCxTKHm0Decwp92gyTGn6T03lvUzRTJgfDtor64duLzdBbZfLZvFlpWX
6m8tNj0yZqGIl7EJFwsnFejLFaCDYfMmMjIq+S8ng8J0VPiieWapNHtlvVF7idZ5
khCcdPtO2lA2FPpAjnSICIYjDbpTGYgRraxq/ERMzewcuI9Bdpv22ekTLtQgTajk
rKjklJZwMtEEqW30jMCziiVNLnyjzFIS0paaWVVOeWMlsIjTHyu5fhN69zPesh6P
xiv2vtKEqq02wNsLx3yVJZA8+MhJJDSloNoc7fcufblyejRaoZ7ZRT0ssinDNMl6
m/WcMPe4sGKgbcmyCpr+DTeATAfIakWIRGVUNFFuHlxY3SSqYJy28usHenKTslJQ
ARQ1ows0TsAW5AeJYFsYZFcdszx54Yw+V3CFNSx1v8Oof0m3uElWR1q2enm5SyZB
TqBMIs8Kf8aUt+MpArLXa/4ZL0BeQgpn9uU9a73SdDr1YcPqZZmfZTl84zdP+MD/
J32XP05yxOLYiZA8KWATmqqc1JuzsKrQyYUdTw9d2/jGsVxFjY4Wj7S+CTgyxJ/G
OmpNIwsBKmAoAAzNmngjOzorTnTF2Q4+0XMOzxDEFLtWuH1AKA39Qw62lUsEuOep
eaGx/eSohmJS69Vm+GBIE6pHpMYuG+O9CNsejfn001TthsFp692LMlNEN6hB0nNo
QyIqg3+sMiwkc/JmXq6b+O3/iO0e09vkJVMeEptQJgn1tIgzMrAtU+jotDMGY4BW
wlwEhDynsnYmVuNjUzn2kn615kAVG/gxCbMhEmWMePGikmQL8A7v+WbvvxNDOHYV
Wvj+YerZrDSA/4LwKKkNZdQcaJpdWluNmy0zSkRmSkShKN+0EVljaSqaMkKmo9QP
0WdHHTjWD9mqzztAeGBHGaG5E9YpToSifskDSo9NoVTWd1a0eYBlBQM7NWkgOS8C
X4DNJ6jCUnAdwmVq5yAKm2TLsSkbxjvg84KdbsjgEYbVGmebocHVilfo8GhOr8Cb
n67sTp/FBX2R2958i2jGu7vJetQtkXriRqBWXJcuHCqZHYw6lHvPeibuW3BWwbsk
45pUNxOnj3DJEst+Wd1ghnB078qanCvbtQk2SuNlu5BN5qDNTXjbggWrl+p4RPHt
dfR70l32F9tMjzhZJ/IUxPXdPsm4AneMrT76fKfATigNiH1SJ7upx1wgBd8/eu3N
w0kvQ3u94FjsPJGmvqHVQ4jA53IVHlBwL0DV+9Q7g7XAyi9jtJKc1Pw+Y8BbCvmf
PFcXq+WpZEIrtpaa/Y6uBBkeN9P3DWNaZypBuKvxQrs0bSzwtMg4LfUOUgeFvOHz
kVifzv3Sa3XgqHsh287u+em8/iSeHrHfXIDBPFwLJ+XiEmOY5LuKCOZttXdEZ20g
vWIym6g3erQUGfaQIoBeiZmLZchM1MnNy9kiBKDQIn25bOFguDMhIeZiIjAwyDJC
yahXD8zmw1/ZsJTM0BlHm8O0KDG3ABan9qibFlTquFt9Mb12S8c6PYcaAVL42nul
XcIUI8Agj+c4Kh5OmlzgtIJUSt9yBm75pQ8hIy7JaJPNBo7VZBj58Ezqhk3cjGvr
9DafqM2San8NLxIRtHO0zjzwftuzglM46gDSgKd7hqbFWAGQCzw+WHxZkwkH3kYl
3JdrxtWK8udVZBXwshjytz+s7W5ntYC60eNnPDAx+SETnsNpR2yAQSSnTBkAsrHN
Aj3/HauJwU4F9KmiYuKhnlUzDnj8cP81m2tmJEquWEeRLJAh5APcphEtvIe/aOLL
1jXeuigkZ9Suf8euxEEtkUFRYNG+bDPzST6PjSXKLcUYgioMbYD1V1GJmeHyo9oW
riI09ZqzLWPS5nyB4qr6u7xrbsQYDDjjjBkuQCCRDscI/n2jFiTgkJ/ajoeCi7S5
0NuBD7vkYYkCgRemZh5BDwm8Mbm8z6AAeFdBtVxjFhG/kAdqo5SvihzqYF+Ir4HZ
CKF8dRwbiHnkogwmArTwmRyxzQRZfZokes5aWCejxQYXlKY/OH1InmMat00fbYCm
8BEqvuUz5wzAwk2mRSkWM/JvohpdJeDzgOnvik/77zWY1XrYykBjSJnUGgFhaWuu
GgI/6waMWhuyjmFXj2U6uafbQ53sUtOdzXrQSnvuK60rK2AdxEEOFaTQBw3BX/fp
W2Rr2a3HtqMbf0FIciz4mGH7mZL2xV7RFM7azrK67YJ/NymMPkOUy9cYRiOz1eLz
6yeak1QM/xsOBex09rTzB1UhSKOUJuGTln8LwO1xje7x8u723UNgfo1hsJioff6r
HRup6bHBeUhoKgK8jPY5eRxrKCKC6Ddj7tRtDjvA9F/JNYSjlwRH3NFjl/R+zf7S
waG0S+GPRMt1Jeo2wqKYf2P3NoxVH+gsh4RVByzKtrVgseTRRhcDOhg7UprJJGwn
3opNcTsvEW9AA9if0CrcEfrCzJUuZHTd5hZ7UwCMZMy494zEc+GKp+HOfpfByeBQ
TjZHlYehYaKNUmHqz5Rj7NqRTvvnTvNdFP/uf9+U8nLjRw3Tml1lKVxA0fXVH9kt
HKhvrmqdOgwyPUcm0lh46cPZjZ2SfEgCekffS594zO/dn6P+iyRNPK1wbTG7DV11
S+Xnu4e3rdM7mPgvaRjPh/WOrFrKGobGDXBMNrCbEZbgew+vdfZS+scJ9yCmYUkk
gJwGSLagUgSWPfaxDoICDMgX6ABdXXiamfKoOX30+MNGoNPBD8voXEssrjFhku0L
lFX0TZsiAnGg94SJRsmWmiotepe2s50QUj7jebmoUlLHqAoUL6raSLfg2IEl17IL
VOHWqztvav2xd1VWVr0Pw5lnnfkiY7wcAU+nXaCeHtZ1/MHLYaoxq9u+BxnXufuj
sHSntHwI/g4Zmin8OEymAT22LJbznu1Lw2D3ZH0Rm8aDfWmyT3DjbDVmOkx36ket
bW3R5DdV2Mz5tYMYuqaU1W1zaMXVTP6kaDP0s9Cl2PJnS/HkadjBqvceOLwzFhrj
9ZGd3HllIAm/RycwOgf9JQ3UY/oVSjKgHusnV1Q/3Xy3jTrTyo8A6GQzrm/6VCZH
/WV3rKwkY2nCph+K8ebYB6BqKWepj7lByFY4+MR6Lp6/b4Mt3IwEXS63xYtrVeLz
MoL8KZf4bfItRfM4FzupCe8ATAHqD9TgEo+g7rkJ92cNwx74mjLtuCVjSZtzKPTR
eb1a+dVdFhxVrELrPxt4XIcYh1WE/vCIugcQEp4ZuPVNLhZKEB+RdTN8S8+tg1cB
6GuURuApKTFPsbmiQ+uif3n24mrK4j1x136VGa5EEizD8CpV0zzj40O64aCDDp8l
SDKdq6fq8++8ZQafxlgCc0STdIMVmQ2qyRndPXVoohRqjEVsmvx3Swx71vNYcq6l
14OIqSvTulHbIoDC7M5Fo50eFoEeHWy3jH1pBMsneuTy3QoUzqQPnVhkdRXMz5TX
DMfVPbRs972c1xXFqnkAvaEfryUC9INigue3MQo+Z4M2+ao9Qi6Fxdh8d9FNV8jw
BGutaZ64awviwaHgthRNnuiV2gC/0jStSNEoKiIPd/FS4JJz8M5kW62cRx+T8Mai
YCtwlvndeJl5jAiZaGygVVkRUHFH8KfYEkcK4zBkZhhq3K7+688WrSsSplmdayGm
fmkgd8iR40hECueKdtIr2wUn4KKm5yBM+KweRK5ZTdHNu6l9NlZYwBBKW7cqTnpy
0U1wLBbc7PgyfvFIqg5n0OL9IuX/aoZDtthkURwxbA2ce5MIU9ZUCHMXF8jZwMWO
RU12EhsMeGtZMgrCfrMpYlWrkIQ59eupuUHBNCIvX1AUUk/vOZn1KInEp6f/WHuV
j0iZD68V/f9oxKKfu+MbXIaPOLrOkPOaa6+BOz5UZwj1yu5T3DMfTKrx51+eO/jV
+pNSUsfUh1Yk0wjQ2CMbl7d7q0Us6UOG/8ztxmI97oxnzLkmkoju/n/ry3gVtkNc
tGvaC32MGWBpqD+Q6HTyJsIzvlWYACY+4HIzUtaS6s38CQIW1yTkVzPFo4AgZlsu
39dbJhY1o7GIzbPtDNXg06I27bGF/O/XqD2Dh+5mlI/TKWCoCRXMcli42GpNQ6F8
fMz5ADiqf6VM15xTEIbSGJeWjFL2wVIbsJpwR04GQ1ZhGGZU6+6Ee1sMyji/zqJS
LSaoNYQ4fcimLzX+PfF6lkWrbpAdAvaM1vMU5Hoe1yVyJaRH/75wOsChki2sKCiW
W8fDA7hUt89kHiIbpy1/sExIKYvlVv2HueLwT8ySvh2HaHC3ZXA4FRla5ZyAPk56
4nDLBZs86wOOTK+Rkj7IKONlJzW2ZF6T5DPmN3bq/DTcESzJs0ll+XWfFHHXOL//
GZzf/0Ldnn35Epa91P7u4xZim47UiKuCT0uOIZQ+2WSgNY9wP+ns1jQUMe+tmEqX
BWCDwd2lXAgFSjZfqdsnuBJQA8cvTuXjSbnNiMvkZ2FNSOQMPCtMNA9Ha9utJE80
PkQN4fshTa2ZaAQuzwJqP1guweGrtFybIx8cK65YH9lewAzRknwBWwD1d1PDuhN5
Y1kYndTEZojR46N5wxH0ZbsbhnoVHvJAM5tIp8rBkK9LW40QJqou1Mh/Gor4/Pct
HMAeu22k4uyMSW0rdSrgmF47V7TABkOBJ9PMbGYgrIj0IW5z5cYhi2mCVZVX8hF9
SxYUeLmwEzj5dF59ZsgSHewGRR7B2idWm5Xp25pTjM3g0MSfI0WvXPk//JoD8v4c
+1mkQySUHUrwxoenl1kbn0iDM2zD5wUcSBfeBOS5+Fy82S87zgLS4RCpAbspO7YP
iQv1MBrgVIouAIurv390WB0bZi/+VxdxjPJCs3MAQwJRvtrgsIq939l4g1Crxleq
y9KEVC0iMl02tiHYZhJUZKUzwW8eWMRJsI+svLCcT+mtjay+AObq7K6uWqhZEFAL
4jb01IL5tIO5VqKoGn9TPRxglkTq7GeC+mDM71qhNMLJvHjU8vEKKZZUY/KFvvVf
0QHrM3LRr2Dn5qp4vZCMugj5GpV/EuklL/Yzj9NZhdl6Wjr8V4BF+SeDA3xwCRND
oqZ09GX4s2BoShlybZjMvuwk5xNXMSWLQEVfNQmZLOF1FCeOilloCpTOr437ZiaJ
nafJVGzK+Z9oFGYubowF/B/qvfCWIpbIvcLDEg+e4F+rUjPsHC9dBDYOTOM+BqhI
OQFE8KTIB1Q4X2y82UE4ss9VHFkQTBTEKUFWdOCS99naKOQPtQ9pdvxZQKNak9cu
5O43Nwg9QeCd1A/lNfIoXSZK0e1sy4YziQtlVKjoUGsLNAdqfzvSKhaIVTlqoXWs
p4M6m2XUXvnHjE9KjdJgOBfHyKogVK8mSy7YWaLgD7DVB9ApfzzOxK+FRGAB/gqy
KIL6JKDsuY3COitT6Sxs1eyy2GA6lXOhRV23cnUtuI04HPxlRFq4H7k0qJtW/bKO
IXNVmjDkIO4cK1FQRX/kK79BUCc15TiJ16E7e9mkgDcR24Hsck/XVsWI3PGbRedN
e4O4dOCrsYVjfLzExh6+kV05qpazsTT5ooStE3RiSV+/CCy0S9F/b/VPhImca3Er
RVds5de2dsdgWkr9/qGU8+zut9WkrGaDSrKL0mp7AfNYaUFlfNzA2gglgTwUDziE
nIOw0p1oVpmDKr7LnV+oxV2WSNgt+hRNeL9N+7DHADpPex+MCarVQ9k9hcv1akfD
aXxadWUpdk5QUOjIbCmrPkZeKk72hzXhxzM4QxZ1Jnp/Je0S0FF/v/r67fvf50yU
DR7O35cRH8G4nI9DgmBrNBIKh3qa3ymva+2CgsWVV+q/PMfYdiTVyy+Tpymr7hbh
zr2HuBzh1n0LBVjhVzbQ13eb3Oex0srt3gXtf+BAz0A6b4uIcGpTP4n5ovAMOOFO
zDlgkx1950K8RYvA+cGD9/HclBMo7RNC6QYqTkzHxn3SfdS1ftoewPpq0MxBhv6g
SM300u5vk9PSA4LjRaWYJwbevHbt+jNkOGSRddLznETZsg61Dpf6krdjfcV3ESf1
GR7zG/w2fLI/9jN5pRlbOeFyXXTncUyeGBjHQkuLK6615/1nT9l9EMNoSNtPoQSm
un0ulmQr+p01t5dVJyWXfuWvAFPDCFNEmTC5kmn0cKG53hsAdWEg8/vO4x+jSjIc
Kv72LAT+3NgfZxI0fFsx+WWwrnE8fFZ5eFHPkrOb+lw4UAUU8oX7uzF2nJX87IYd
Eg3wy68cSztFyz8APEmCRgWjva6ixl0lndYV2epdEYCdoecXd1hyMclyrEiUkgv+
35RCrb363mG+95tZbPYHou3FlXVt4CLTX/cBR/j60IqyIE+JJbC2VXbqRAvbd8Vv
uTEQZRvPWpytAm+tDiw37o9ryITfTF8waW12TZA4EC5HLPhPlIvd4qllchu5glnQ
O7B6HtoxsM9NSdKCMtvZWnjGKIFRpZRGvskmRCawvkQv3cfzWb9Rt41y9qvivumD
Ua1cClhh82mserqXqmemjhYu6GBM1eu8UorFtXlnE5DY1hLwphFwbT3U8uyiPzEn
rwhqqinrTiwg/GzTbuWhvlKZT7Lgn+nTEo5ltNTivt23ZuBfTZmmFrxw1t4FQCPP
1sdQagBklKFodhRB4h7KGDbUr39Dt+BEgJfb0Q/M+pWKECaKtyqEL2SCFf5lf/sU
M2OI/rEtOtlJ580ek6oOTm7WSJofmAvlfDfsA7WqWBG6iM9eVH9el0VFAmPc/Gku
THyhrAlwHmtWZAEyjujp1lV+rO4Wd/l27NDBimGNxrgCmxW5yzicfbGQTP30bcTr
k9GQloxjGTTOeGlK7WPAweLknHWiI62u4Mco0qQyjiHf/MSs+rBBXmApr7U5TRhQ
Y4Mmy7BbRND+gvlBRZhRsLnTnEalIL08wXffVbXlvZxwxW55gCUbP54LMUs78pzA
+nVwNQaRzD1wNu7ZpalSp0cxzw3Fr1BdaVNBSyAECDDhMNShLjD85Ta0mB9QILnT
DSVrvYglWZLs3L4F2Q3GCMny6adQnXy455RsMAZ/rl7f/gS0DZHkQDgR2iHw6djH
wQdroz6H0mN1xOIuerhTOROfp0gzudgzUBEUmNo+Tbb74yvYgkExyvOLro1LJXRH
Cx/R777IUlkO66YKVV/pxwbFsXc22gyOdqcIwUo9a+c2Ztzi17eKDpSOr5Voo/EI
xpDipUFRxXf0YR3m0Tqw2wiyEhOB+FzqKZVISC1Z9SJGcvhWAs9M1F5MRuYTzvRe
CByQbxaowuUzq7Ogkf77bgYiZkt1eSiYtAC2aAugFtBFlZOC91hmTwRuII800eaJ
9vSTkR6THI3BQbdVan3FVUA1vAMK+hXq0SXgiwKjwHsN2YYj8ir8Iny1RmITkN1R
rkEqfRh7v1Ul3XXnF+YFGw9/9fPvh1h/bkIIeV5XfDy9BACz/E4vKlZ9+f1GJd8k
BDTaNQTI2wVxUO4Wu2zDiP/L5a6euVqF0s/dKwD9LPIw/gnLJ28eanV6taO3KxY3
GW4z0dYgGy+K5kWp8w7iGKDUrLBatALEFUv0u6JwcOAVtK+qV6K0vmeGhuohsFN5
hlqKTupuxUU7G5u5m2Boes8CEX/++9Rye5GT1wzAwZSYXDthXwDoZrKf+n64m149
ZyxFVkhVdu7M1Bfy0dCppTi22a+61q7EDksu8V1t/BBYFhuk7VSqPPphfcQCRXJw
vuXOZMEPruRQfViE0f7yNId6lNL2b+/1iubWVMeSHnnqkJmJ4Hn2w+UnJGuxEnwX
RaqsSJ+SmMJqfgGezQMztUEWfp5sQ4GCPmtOo4kGWbr1UB+cvv2ovzyG0WgttvVK
Q7n/1IjXODoN5AmK0mTcFjiPCqpodZdoNsERhOnASiRWsmI1zJv70SilgVnZiQS1
+K+/jWgqyXEWaQTsAjPOcb5o5co+V5lySTq6P+0M21QaClNbJOmqzN/RYYcRaKpC
Iq19ok1k1yEGfGNNzm8NkKHR7z+rojhxAfWYw6KoRm0ir1l/mE77mfD8jESljkBL
CB3r6LOex7mZcqsEjzhXz9xgZ4xbSbrymgvaOZSalDJJiGpvZm0yk/jB2FNHIpZb
ZlCQwLsf/qZs3L7Q8fmlu6HITct26nwExOtxicMyXP5fiB0Jxhx56Evk8TLOJIgK
Pykq/aSOL0CZNh/skZpT40PIEmaC2GA3dIwg/fEb1ggOnSo4GyaarCgNpTEARXe2
NltW2PD6fhUlPRD9zqwBqm9xJ8vpjAZQ7/yimpivxEz5/07kS1QWPkdcbu4kiB2e
LmkU7KFF/KAhDh6oWS9eGMpPWsGr14vDgA0WsTHJPTU5+JqKRppWQcrrdTygGLPk
rW3+NCw51+qz+6kOz6JeyQKHGbpUcIb+0Dd0DjI/LnuQlZszm2rtdjkJYvpjIHCY
USJGkXYM4Uc1u3akJBBEMv7d0zOGeOdTNtJynE1ixehj/7BhlRw6pwSNH4FYrwwT
imQvY+fqLXwDYVPLbx0xh1VOs/em7u75jmjTPOnEq8VsKst+lItCokdIIVTEU/23
pix2wB8WHVHL5axX4R6686uzvOMUNuSgk0sw3hjpjubMRK2feSyQCxrXLdetQtMk
RFbXm1FJXlUcpvVjJ+mbCskd9eWh6TqDORwtjVyqUc4kmiHbK8CB/Nv56V6UjuQG
dVxQdKbH46RDX0a9Y0HnmPvVeLDuDvvHsmX0OCd3ttfx5FS1YdtGuM+ohV7yfYJj
6gk2rtrHADp/K5vBLEb/Fw1nQUjFZTYQwaLypBwdM/vS7yO3tGOlHY0gXxIIrswo
ZR0pt5ENyOOCQ3y4AY7KliFx1gfXX1nSE/zlsfrpgasNRuLhAAhpZ+duacSKZygC
eletoww2okfs+jikHZZP4jRitnLe98Mnap6smao+BrYHiVYB/dzE2+mso/D0YMLF
bbREJwaWWl67ViaIAQtwJP4NpTrkNrwoKSveguzWEQ2tQaf5fytbDv0RSdth392A
LgihLL4LzEfxdDpZKUz7ppXNZOdk2dTf0YgbtRA37obKszh8y9VHefiWFXRVXRCB
5dlyiIjUuzPBMMCB0TxsANxSA41JlZKxZ7ECCqtkI0GdiVSGZfkgBjmMWoDfff5X
Z8To9asls8bXhTnZJwPd+6X1qRILE+ag0i+VBAxPrhG4ZcG5RgM01y08X5gwmjcL
T5d3iLDVg9Y7jMSBWdj2Prg7oCQ/A1EnYK+iM/GB/6nItJ7apKU5aZa8FLwM4I8e
CJ3PdZ1qgAxb6esC09ius45zeoST/d2MUT4ci9N82pN3YuvLdQBZyzw+IzWnGVWF
2QL1djtwyGobbfwqTEReHkE8mxAflpkp3g8jl/F2CX5WJZOZaA13NWP3PIYqU14U
JCvyPy5G3iUKrMrIEnOdNQm/r/n55NKLwQM1bSs0jOBWqnz1SZaCoTX6sDV2C/jr
LKSImmxsdtubvCSY//eVVrxvrm9IPniwma2qwc9weU+rnGNTCU0RUmqOyjNpmI4P
CQHZmo0eF2oQt/rJC8Q0WmHE4yo9sRj/xSh/+qRNChZsFmB3FOsaPdY/YKHvRIYS
CK/kkf3OPHKlMXVT9KDJ5JkMJi0OOzgVjjf7T+8d2gKhDUyJkaT6gmjj80EHkpwj
OSyVzmeNHLl3dh5aSyK1wT6Rb0PRWxzudlBfUEZghleSfcbHnau0ZvuiKXxYDbOz
XMoqbZ4xucOFL3dQ5ZbDSGbIPqULXIKIN28hx3fUPX1D9OQPFqlnZqVvCssOeUgN
ymVpv1U1we9mijiyLlNtO8eSEuD0doD+2mJjq/gPyR1ZA0ReUlR1vMk9UGC5xgwO
6avWiI8l/pUGlxSz7gkYnBSY34i7cIreAnSEkteRc7JS8kIJlRtY3OfwGYRjVSaj
C1Fll57xEJLYu1byf6mFQqcYBh44ClthMZsY+Pj+r6v1kHIpqznZs9Au5YRn85FF
X9b3MOanibjmos/vJZ8y6s1Flwyn6a5Rj9EhXJen4aHbi1/yCHdWUWRtuXlh8COd
anmpL/bFnKP6kJ51eng9Awg/EDSOvZIrWnFmWjtkr70bhO91CQozx1s8MqZq/LFG
2UCP+0Cx4uKMSUBvYGoGL9EfM5ZYZl355oG1R4f/5zyLSFuUlE61UkWLEfVv3y0K
ciUJZ3X6wdYwISo4XM+RIbZ7SEW1smx74I+vcaHH4zA0ctHFxO6+xD6ORnuWL0gq
pPn1MfakIQMD4W6vM1ckq5tFrsekRqaVPNe3hu8rAeqrOu/xtHI9fYAJsA8bGMiO
7j904gRqsq2URjnEPmDl6orqAd4pZjfzhEgRfhMnlkZXQ3y7pahd5hbYkdayPSC/
F/sKnONFU3xVvnf0gR74B6VlMkp1WFqA/x1vBQpOZ4O83tfsafYa1WOTtR8NSMYa
SJt6Y6+P22dttyC+4tXvuPKKH2qyoO1l5/fJDsveB6WcyaQtOZmgqjJ2++TGezHT
wD4iK3ZvAKjou91ysebSfYRSA59+5wOsGpnrUM4hnYBmMzgfj5Wj4TaSKNenh2J4
wUQqGM2EKZNBJB8laaBwiu3np+xX8a3mOYYDLQUR7PF5OGsqpJYVH4Vd5L+vXjKs
WHGJcKND6/lYCM4CY76udKbs5NTL42ZNK4T4Ol7G9N9Qa7nQCOfhBwhg3YyPJtqI
hpTBfWTrl72z73vNTEg2l00g4Vr/b2xi+k5Faysp3+d3LsD8rUXZxodErn5OE3e5
gB/Ngaeqhm5KeqBYBqwgbNjnkInYwZ+MsX+T9/2FpVGP0DteJymNsV8tWA41YHu6
7NBCAr8kFjkZ2s16kp6+SJHCi1iJPsRZbP4qG91tCf3rgYOowXLeE7qhr5uVT2ys
XqmcgZBNpRS8wetACEO0D6bJ9zIIaQOGZW9DOjAZn5JW3fhlkp4RbjqgJ29fesWw
3E0HWP862cSwEsVWThFKQ3kdnkPg4lAKb2bbeC0Yy9EuZoZnHm7sKh0CsBU0Y59h
r84yxklT3UNY3aRkPmEy0s4j2m9mF31urmXJXDSv0CUl6SdrVrm6uYTm9OIvvEFk
QMo7yqQFyYgHNsmiha//gmF/DlcYHMFPksSjoXKr3Dmahq6yN2Z0Lsmmju5gxQFF
1S6/5dHEDGc4PzGVkvf3Y4sb1DGooce0r9xCGpdBD92h1UIDDlkgWPdOXVrHVNaM
ZWh7WTu7sK1PGdTCye2qZYksNt9+3pUY5kwf7WgHMU8iCf6SyVCr27Pt4ibhDApa
KWa8H1jatisyoWtKA41TnbIax1/pbcyNeTNB7VVPIvuz8oNsd3/Dm5h3hy727XI3
9A/qmZFdDMCUq6d1a7QlYRAtDTohM3JtASlxfgUcM566UvGRv2Bcp+KrH4UKcU53
7SBXEHZ6zJcvR3reoDFbyG1B1qlY19TSMAb9aYy43mDymnPVCAuPVzGkf4V4zH1Y
X6rqBbMGU++fzL0WGj+atrADktQuNPheD7sXQtUXnHd+PPUUDKcpJIYwV2llM+Hi
joE+FlLq8d9behvY7bz4zfwWnkpF28hVEiL7QrAY/fLVyx90nQ0AmdzaZfIyk3og
+AW/A90UIE2iSEC5d3Pk7qpQN4APSLzyTiqkEOoaaG3GcA61IvFDi9dgwp4JyOQ2
vbKxcNu5fY8v764+CZC8ktFyEUbHrLXFKEr/wZ9SmA7bTXACAztIsjHKImxd24E4
fgAZ9bsh7Mk/azdEVVnWnKOGVya0jFksFoCeJGLfBGq/dz1/9poeaZ7Su+pkV5yl
FBgwp/Cc9Nn3FyegRe6Xzs/J8DS8HgjQLppDHtH8uijtCzsgR9y1gcoev9C74y/u
n6U5DR+aA1m6wvoEuRVD9xbyTXpdDbXeKPQCUSDwbtDFRQkAfcaITWPRzWLcBvnO
eajoUlRomDfaLgvULUNgjnUh3zlkoUzpa7YWYs41VqwKHLbArXkc+IkvHw2AA/jA
RcgkAUOCVLJ1NrspKPyaovJ7HMuLKOnjUraSD2jhncujBAS8MSFMf1mwkVzID/iM
TnxtiMX0AnI8ESQAlyWhGrL73lpnBBuvrl9FosY99rTXntJX6SJZ9ObJHxoGPy9c
E0SudYiJ/0S3wcK9oVjDYHWyY1ZVtsZrJxBvugBevjMmk6U9E0RcAZMTINJ7zFMQ
pA2UEofg+B//8QPBXpFuTCVuihPzS3cXDTUbc3+0JN03Yyk7JzLYAuShsMgdei14
Qc4yJy+pIx/OwSRdaT7fU6arkWbEvgMb4uZBHmKi9V5hDw+O261ah2jWDuvsXw7Q
c3+DoHfuOXLWzlJfHaTis3KRdmIV4ALtLLsQ4Y6sX84ioy2ROeLO8eLyNOZloNwT
fR+0mkktJQ9UF/aXrRSBi8tb5MXzTGjJ9TuftLT6t2xfWHLPSsqfJASsiQo8PTYw
oHz65v6eJ3wnuqG9WotFpPy2kpZnzSZ3JnH+qZwjCcb6/180X6yqopFmdPEmFlXy
arJdz6wuG0biAU4tony1tmUXjMb9/Xz6ZnAMBPAQS8TPNmQrcdt9+3WMO13gRAeU
5YDfBQX/uE0Hw0BwrhHi3otxZoiXuFPHiMHeMld76JYmYbOrOWCK9EiaQFkrRjgf
oCihjdlNE8ZqCn5gtTFnxBmiXCm433zVKpJotqr43qYCQECEWpa5r6PBeYiFKm2i
aYj9szELv/u4MtZJRtcbwadGeMk6EKFuylopQarTV8ICB44OWjnNpRWBe0HmSZPf
I0cYV6hdpk2D7cZXXjFi1Tln3C7CLuNM4HX897B2OFBlA8RBWF5M0ka6HDcFD+j1
DKG0INrNhsLXbEv+CwYnNTk7Pof8+vrPKrKIp6fGNd64TaXQXaWqbogwPCuQ1CDZ
uT5qFuA6WRKjnJ5QyN8NkMV9VQmkuk3PzfjNY1MXj42qVnTJM00QLWVehadfPL6x
VCTVYAW6vA5xbpXM93EIY0zuRNMtmjbYkwLn22KbbSvoMDJVyzZ/BXggp2vv596E
kBTXUHfHj3DRD8bbhRk4K4Jib4VV09EW7agu/l7voiYsSeUCFCF+Y3d8OaAQnjRV
OugwbxUc2low0JpL14t3mmdPuE6e4sjprBYRHT4imsuaxmNZL/OO609azvWKXCCt
8g+ISMslum6UCEGvs/SO1E0ctUyGdx6nq5rfxHmyhu4bbWgVHVZgf3u6cHcIp1+W
bopvtL9kQK+YPxEUpO0ufxrYJANcp2dn+Np7qrXdzaVx0yQ2fQ8DJ9uCBb5BELg2
+mrzrX0g0t1ZHDJNDu7aTOCIuy/ltzPVfLuQqaMrEoaxgq0lE+tJ/UshBKPfZGyk
Okg3QGgrwGQdmWrg9QEWkTAlpXajWEMyrTTb1lltwTQkUXaB/Nxgf59bZBpJDtJ6
qqp2NnvY9v0wwq/GXCuvKiZVfLXPhPGME7sGHc3GC4AHU23zRfkY27wtK0Ht/WHd
kGUORDcCx4bb0q8j+ZPskdi+QFMKT+LTT6VWQ8oIbR5kaODByVPGczkl25QGvlxM
aBe0oV6j8Sp6badA4TYpfpwXdLeQ58RtW0Azy7ZFHKNy60TW6RM8m4geRX5hbvtF
+9mkJezSnptCQ5wpc26zXO8Ydy/1iVS2qWGMr2n4HXIAH4IScWBD8nUfD9BoDJg1
qAfE86bf1yaI1za/vhjsI6qWjAcavLiErk1kztVp64CuNxsaeaFuPjRnakWC0mO2
NzKxuFGmbNRXyEKZaHK5fFkXsxmB8zvH/O+7p/kagsW4xwFaa2ReUM9fTQlk5xyL
za0GC80KJeNYYA+uM2lSGi6B2+4Rg5xRwLQ9zMPKJHOE52KIo2ypcFKX1gQ1IwBK
lIXRj8+tbJ0E8xImBR+3vOrFBQUwPc7MOPMlvUGHMUPKZ2NnHJw25nI0+WA1hP9u
g7LrWTMbAQPaG2DeFY20TaLhSRnMuunuVvchnjjGT+KaLiGdfDxfLT8ucs6OWXTV
wIPIf3i5EvZBwz0pDfHWiJ2sZU6R5Gj9qtu8WjIMCzxwi/McCWsAq9jHwdMlTKC7
zquSq/ZLFgg0curRYqQ7VMia3e9CnACXkCzH9kkqM5zsekylmzNkDna7osTxrcpq
jOsdQeHWAkU+IJu2NYZe1J77q8+dmlTlaNPZV/mAY0jCnjErPMvVn+Pcab+688cL
j/t5IdLfHP2a7KazssvXI0702JT/GRnTRZNoJPVBdvluTNNPnFxaUeP7jX/2YURv
E8wheHAbxQ99358RZbEtyN0Zzm08lqFnN8sWZHmS8uo6dNjhGbGi7AlGb81jsMFh
qy7KwWUDwLctJNVr55LMSz7SzVr8M6TwVa0XbNh0ZxueNvOs846k868HCyvTfAP8
GS/G8JV3w/a7R+6ZPFix185CfKQLLRoy2g/h5dslKFGxL2dWdX9RwnAKLmdOx0uP
QuemSG9S0SzWwzV+k7NlhOSBH26DJi2C8HA5MMYbsAsTgnXFAKV5hsQkvuLaNsev
665xih/s46rMm+3EXMoWJZdY8/PaHNlvy5haCTx9tZhrHOk/uhPPeEBK8QE5TFq/
iDio3+7QqD84VjmPRlj0qeUQTbqoJa1N+OZ/GrxyFtzv8sDxZHSQCM5kk5/bop2v
L07O0zZuL24aK6S2qRt/Xlaby6cHfHOV/PllQWNr9xNMKd3N8FDrrtR6OGEmfUsu
T7zXUYuLMLvLgLN1SmezZ2s5PiqLqqWpdXFY33d6wIyYLp+Yxe4MePMxrQ5Ok8ZT
NmESGuC0X1Yk4gEQq8SXwg2yQXYP5G6URfD9jfYcsgFo4b175NwHLJCTgIn/SOTi
EZsUzKvJ6tREK3nMcr8Va1iu4Ecbzg42Jc+F9kFHilfi0A51DZauyd7nuOt3xsZz
R4Yp0IdBHmlfUyWICFtyba3HS1I+PTwJOO0ZNseb1sVaOvbMTDfMw92HA286OmfT
yne08SFpvHgwgeneObBrBAbek+1YRKjSwc+PR6RY5tpHCDQ6FysCZrqxwmzKIqGF
VDOptSfHiO2dNP4XwQdwxnEckZJpS3bUUVxVSxtGw8xl2eqOIDBfgUTE7qRXeZxe
3XrvJAAv49rQDi/HuHltF37z9jUCcN8HtSoj3o6frDFfmjwi3nYHT6MHI+BRU/zg
JNPDUTt+vTHDEiTVgZ7ATZWzWkfBivo/7iiF+1VOKSq3DtHkTpedR01wvmBDe6MM
qzjO8KNOTIZzJdt80JSUGQOJXPRn+IKGM62Sr+ySDI/QG0TX9srv0IY/ROaYi4lA
AVRQEI6jElaEePOK+3X1jLzIqPOxj9hqnvURbaddmOFDrQxRxaFC6yZhdTf5PBRN
sggMMTntm2fJDeGY6Ni737ljAxUe4R+SiGooeVo6IfgorTIL2k89SGIVDxDYiFmg
4il32LVP2UIZqob1h9vRwuHXKQCFnexoeLgXywar40vXb2pAPnJf8q1sTyvcHta8
xV5xAsgtJZGW8YRK7MWhucCMy/w/e0bnWEnou+/DNaDd8Lk9ZfWVUZuhSgCsVDVX
BMq0LBnb+eFVCZBc/ADwWceGZwpUhbYgymxY+veE+qzt3cTL7W7AcQIU1lQn6IwL
WIH5PVtw2ThXJcTQfN5y9ZkkNC5W66KWXZllY1AASb0qgs1IV2LaJDWY8ItrpGGL
4ORxCyodSaQpm/HAkzpHA6d9rtUz781sLLJdSKaf2foo1PaVrKFZTq/2YZqdhGUN
LCoB7Bn8p1ZK0ta1YwmnP2miz9quIO3AlwjMTXYIW+qalLFlMM2f/132ss3uImqV
RBsfok04Y/gg9UOf/QCS6z0GJTzBcd+kDyMBwrdPKpYg36A62I0+j34Opqv4VqCs
bpBxR4nQS4K6gf2zIzvd22fSFu4sACl8UXmkdCp6nv382bb0wpGjJdSFsFrBTUpS
IstwqyVXLy870TnZQnTqAPPlhjafmYunWszKzZnltKPSM2yMCqo47cDiHCNKXsjg
MN9Tah0dnx5HRW2f9w+/AOFj8kxAG7qzGhDdsR9rkHN/Nmgvg2kkAnKyo66w/gcK
P+jjz3J+1Sbamxh8Ig4hRrbIvy9EcxWcbdXvya5ZJpW9opxeE9L81XQQnvOclBKO
1B2QcmcNzgbGusMAE5xPYto2kSECvBLKX7jcl3k4O8zWJhOCpuK4MYLsPzn57zaR
mgYLVtLgoyLcVpNm+sghCSP7/RolMm08g06KV1d/Cu58VEqi5jVSoUwqPrRxpAow
V3HLmiV686TQzlgRU7Ap+KSTdI7hrCPBwUgLXXh6iengOIsyhM2GHAbJrAEy2NWa
L6tg8Pc0JnGw9twWIv8QOviRyfeep4Nu7C3JIKwgvIheYmtnSN4HL0C5D0a9ZVTf
h1AYnyolo63yUEu1HJ/xEad3wPU1lTgRAZ0WIYbEJ31rZMqUX/cu8DrLRzwLitvx
XhfrUp1dzTB/3+OydJKqXiXrTp8/gyqY3RjJivxzWhRqPZthgCnyhmWbGhWgDY0h
66Q8/NEF4O/4Yps2iH6LUN8Y40vpobSnErhYI4VQryFXNqKi8+H0RPoLjc5MaEdI
OwkYmYfQM8O0RJI+Q1boVlDTfq8TDt8ekNrwWaRSQpQwvCNiEEL/YH4MCsc0Q+dy
U4kqc7sZN1xpd4aTSG2oin5hXt1kmS28z6jM/4/ngvMwCAgTcd3r6drivy46NWlc
rtPjyXnypFdEq9vGHW5CT7G+RHtaV0vlxxxZr1OlXQNOR3QDFyHOOgWKTJoOxTyc
pup0f0WAxKBFt4L7tdiIbaQ4LS6OV+8HLwKpwbpVAiYqQwfqSTXaVoAkTFd+P6b1
/pZK6wVXh4Czd2/iI3tm9IpSJmLnTeSuEe0o7UjK/7E7hAF5QeSKsyVbV/y74XiA
AyO0Lhv0UaF0NULtCjqhgf6mSfQG4EWNk/qyFDu2+PNZOMkkeqUrYs6uYYzpSIo6
58yEExBJmd0Iqv0PlzsFDZ4K1HeetAUsP03Xa5g8kqpu5pjMw5t1o0TTxdmc7Zka
JOIXX5cUZ9d3toK6G/6fmj+ianoeupK9HxqzFzewsCg4h3t3fwPFhRkZfomFIbsb
9edVbFLOOEu9QnZEy014UqMrY9318TNUOCoQvfFDkRmRAtr+APgOdUqMEUsFxO/g
lF32VqZzoPggNGExPicFqPAOu5UAh56F2WmqUCwqIFDPB6rmEUb4CImJ279BXzb5
97kz7Iy6FmCKs+heUvbDEJRHcAm9bOP3MgVdsLIIu5qXK6Xam5WKpk2X9tlNZ4VP
GhbUzNuw4N4boI2vGdvT6cpv6iHlZZDGkH3IcjSFf6rGy8y6L6LEQlMrKaR9tn3n
8lPveYF1yRRdttq2XSQColCrX+uGUNo/tg5VGZPyJ1hjPW2Dqjxjm9UljTiEHP+w
sS36VR9RmMzl5cTM/IpZpjGlRUKqxb3Ki+HZZ4GdZEA3efg9pPAzgEWfuDH8M+rp
6m1FF/JtQTWkI3dUwkGAJBKrTqcp1egeUBReaSA9IwXZ6KOZml7niQ8IavWIdGSc
2pn/gxAZA3Cz9buLkXiK0XPonsrWp8ZgcYpFJIxKT21KMiFAzr5j9tmCBTeqs99k
G1i90gwVFZU898z02YHLmcuVLvdcfZNHTq7E1XeBqFTOCfDLB4CB+C7ig2ytZaMB
FIwmJxwqB+wFiGMCLmcnC3qKVWsFJ+IdcEmsO7Btw+SNlmgQupZPNwpH+3LGaB7p
2SSu91zQPZaLcb5iCbTUw1wfSB4+2q3ulQxTOSS1XEBbvCsodfBG3l0QUruDs7y5
kxb9rrZ7pKM/j0whqwNhcSEKQJ9ECmr/DpxR6yNCMVGaTqOmb7LyM+vbHEwvmPdh
GSRxHpwibPPBqzhWtUdzKHiLYJxJSFwdUTHzZro8IKHcXgHzDcuJ9Tq6EzuXUwIc
zh7r4+cu6UeOnGWsElRfrFfLe6ppyaHw1FaiJLTddsKORtLfhqMhuerd3hx4pkil
1sefbkAmA/5T5qrMPWiD/PceNwwMIzejS91mFodRG3S3XBJyOrcuZTgB79XplzTD
JqgxdJ46onOvrRXGsIbLRhWC/KzYYNG5F+tHd2hfTzYFRcdsxfgoOghSBT895h05
xAoaIg48sBcoCfTqXwQsIUw3nVTImSZqth210Vmjrdska8rbMACxdBWOLTUrr8Er
B0phMm0vhocb3Xf/lomp3OUaPZ4/vi+a1pP+IRcsKGEdetGG9MS5j3z4ZJAIB96m
YqNlS5cRmCDc5lzJKFgY0nXhiT1V73ED1/mcPiHunW7Tue+cjKpul28Mj8Md+Md9
i06WMQeCwdI3+16p9iVV2q4O06HRO2jx/nD9S1fdyjlLGtt+ffpjMt55PWLn9pn4
MfxqvSSC0xT/ZspTuyarVw3z/pGCPGugh/Zu4hVYgFYpMP3+csdVELw20gDDS9A2
OetzwvIL62aLEaYVIXSz0IBMvNuSDP46xNyrJv4KCdn3oc7LMXNul99BQHZyNjRf
B4uaHVt45Z+jPp+I1+cBZ1fj1nf0sQsEsv2JdUR0IZQtO8Y4cUV8wXc2+IDAQ+p4
z+bnQz6rx+ImjDJLVsI6HTuta/MMX07wfiwZBUx7zpw4ksgMb+HE1ANi3Ooceou7
0ejjhunJbXTzJHFRmVFqLFIqdyUxV+U7H2pOx92kLjgFScSG5WLWLwS8fDDFLr08
j/jl38SagwvjtJQfQRh3US7Ypz3QykOSQNEi3i0+w85hgVmBqVR7ki4W7k7cQ9Ke
79j4DJa6AlrBOTgfOZSJ/5ZNxCt1xIERq3mZrGb+NKZZ9yS8p+BHzKta77cPMrV4
UHdcwF6cVk8e7vPxTchA8iw2osxOwdXENtq53NAlFf8KfS4L3S6mzzwdwYHhU3wn
Ib1Ri2C10vArYgroHUh8tgd8PqXrZwxd6ojQT3tqk17qVBD5p0Ivxm8MpvYIUxcc
/ZH9s5tpjuAsEy8lXepndIoWeMjBN91izhARy6J+dGB+9NQZUVmRykL3/kQ/O3VS
xMgMpY29MDQI2RcXL2LoELN76AnWCpn1oWWFJNJM9Cp6vCeL6shAx957nSA4iWwn
4O0d3FCEquoq1PxI7c0er2D8Mv7OUtb4WYUzJtcA5N00AyERSyUvpLsf6ENDnG9Z
MswAxS0Xuo0vfqntv4hnt6ClhS85iGonDZCMA4Cq9ERpzVZoLfUSs1x+DU8aXMDC
dvK9axMkX1yODm+xf1P75I4piZcSqV1qFHuACwzgIHNxf+KO1fEu2Lwfoy7s3cJP
2jpItFtmPEJfL/CuT+m+BctqiyFoWc09atGZgvnMkQwlrJj/eZnaRWydkI0JmPXh
wpjlQabiNChXKCFYe848s6+talrP+g+5yNxOxDFvwAi/xZMX/acEqcvLryNgTVc2
O3URyTYyB3Z5J+v/BA9zsp/gQ/t8t5T90eEuJahDuyvrC3soas4AGYrpNnaC7B0d
VNbYYPidcsv+bw5Ax6jq1gXFWYYYknrwRReBULrEs1bv2GbrX1qq9CSVA5sayVyq
d/JFm0EY7cdR41whdwNLrfaiiayJ3zN7IKeQ7yuO2iFuesn1TLSqD3Rx1aOR2YV1
Ijm9ObIxYCp5zMoh0JBxGrjE7zMVGHo5q7FHl4/yLdsf3eZ75jR5zE/pYfUNWxvg
hT0LR7aTO6UUyTuRS5ddd/5Q9ILzANaIjzpOYxbWlXUgnDofFYQ0ucso28nsB76S
n8pn7dRxiEGcTrL1OyeMnHB13BS+fq07eAFMT8jMrhnMVtgb6o4D4JIaX7+p/Zqf
1FOogEgvTl8AslCTA2VgvFOr9wDiVOCCmzBQpTRjAAyHih+I8HVfQFq/XIT0Wm/G
dmyFMzbqSFM/YQc4n3yZHAm2ENzQjrsmrpa0XQrhoy22ba6GGPJa+ULjSIEintUr
xQRzXHy2/6V0UzuCbHaXtPNiHJotzxeIYHc5PYFu1WsUCJwfvGIhyMqCYMs7nYpc
40YQQewblmPq+zYkS35Dy/W3GwfrPY+XbldHPrOaBurEGZ6HS7BJHU/T+VIoh3HY
aP2hDgI9HUl/lBhjhaVAtzBDrFmR82tJuYDSh1kQJWNFIHigmtmUX1zSjXsmd1Lz
ooua0iB+jKa9SxPf/vta8hfO8LEZkc5uWLr/oTOwp67CwXqnF7/vvAHUv1n0BYVK
dEnTtfMIwOLtTLO+FfjjwXiQxZF8tZ21tiMkHbbd/lyyrQl4l1EuyM7ju2/54msR
pbEdEkUdJDv8ZgvtyQB+c9NHsSK/LXjmrrYgY6jIPBqbV2N/vVq5vOQcyef/MDnl
mjxRJ3o37RNc1rT9J8GJQGaF8JijDEHccTWWTpnedVj2cTyWvwHm0o5xgZX41tXm
odd4WZhkwJdBbZePIgKagVyh360WWmZapOGguEAS2PVWmzYcURkw/4TmMqWfU1RY
lmamIqaLIe4fvhSx6yGbGKfRykSK34ehtVlJZ/UKkeBFn98C3cAuYqdZrN0vh/pJ
kDJEa8mIPST+lqKZsezFZk6bcmXsd27E2t6MZTTPabPp+VNcMfd8ZVZyemZs7NCc
VyN5/wbNTcApzGAZiFm8KdReDGyjVcxzUS8zuImTlOUsGj5Xqy+WWGQkCdHUjWl5
C2IZHSH4XmJ+Qmz7zNL4comB5uDvhuWY3OZhAhpHtYlaW5a5Y54K2ngnEqDRoj+c
SmSLHCyM8nFJ69iJdn1gZxUoRyTg3X+cghSbaZ5pRTH0MX7bJNvCqoy6el5JYu0j
4xalvBCbc6az4/JFf8Y1D8fbwZ+B+AsbHbyjJJFOqLu6KfrFpPnm/yVGk3rLtiVK
yW/X2oMKYHDSimJxBbHy+ITPSB6Ml3ang/ekCMCtOifL1L0qfIrTgrr83LMwMkkU
fSSxTnunXx+5pcgnBMLEQ6Fb9wv9r/DhYx/z32uzvZI0xJkxO7vtI/kr24HpU+K3
itM38EoCLBTswocAbNoUWGN2WlHtEU6KT+u9tt/BAIL3HMKw16PD8Zs1R2CSIoje
oZXjcgSiOTrjSkcrsmXxOmFKyKA8Gb0hGUxSERL9RFFvfe+W1MUIPaOyzt2lsuSw
x1taLppzMOxzPYsv+ElQEHv9x6lgmUVlkBMorOZbkbruO94A3ir+9+SVo6xRcEAq
8Is1SKKMNJ0hBeyEWH6XoI9MneCzYu/ZuT43GBq7LinXW6ELASQxOt+F98Q0fHva
msu17UnP8N6upVtzmB1fkBVkQ2iVmmU0+oAW2QSSz+eHM+s6YyspSHZJSBssNtKz
s2qsnMl1B3UDSL3CSg64NTakPcEQdjz1nHwKKOWmTgpRGbHFPDEqnTiB8MuTbzr2
f+RGJrxtc4KdJnwqtEhk6n7LXFpOH5h9xvGCfn103ymge9flAnpctmx27kBCmAZE
mUemEQgATunUapNJbs0ZMjqeCeZH2LUhbgM2q7IZqfBKkVlEQsgZrOLnDZX58J/f
bnqiaYqQp3X6i3KtShHc1be/66TabxFZv4fCByvauzSB8xPyR0WZZNT8lE54V/zE
scnNmsGrmpoCwJ6B5V1n090OBsywdiYsvj1HmP+8+1Iz2YpMJNQqp4/AamPZCF7E
vrEVKBcqITSuIHCsHd7TSZR0LsRV/PaxGxBPlyVvL7OoUt+Um4sCIJ/bBKLJut2p
IYc3fM84DDtywRzEjDLbEeTRpFPUrLnAXxBFsWvtIu0Q7I741G8KYEOkpYo7hMP8
RjF0gdCkafd2B2P6/CmPxAAIrUcN3Zasi7ZIJKPU1istm/tnS8X9GjSMqmBHEu1k
3NyFwQatNP9fsv29g6B/Q5qEo/9eK3k0dr5fEVk+bvm1ktvcnVbITfU4gzF73E3m
4ct8RyDLEj9apDGwLcjsFlSh+4oYTfHFzvPl5Flb8pye3MywftSl/rQPbKHYJySL
qAHb3QsxcjHgzPsfeLzH2sio4PLvX3LiyBFIHPBxHEApgw30MgvEH/TIuHG4WiFv
FhhVZhoRGXr/mC+0FBgUbADqJ2nePO5kSrXp9ZxP29SiTtW4ZZsSBVH/qw5glxx9
HC//0Ny4hLcdh70EK68IEF57uRwPOFcmp9EqdxIE4HE+ipuLv0VNJR7DuAi/IWtL
i8zEaLILqnltjaBwxB3D4r7wF/P3LQxXoLoqpAMj+CcXARMIcAQvAcd9hc24rFyE
AK+AdLpFADd9HzNsiNehTh6lhm0t5ouKGbTE6qlJsyoAaoRKu2BQWblIr0D7TkoW
YtVnfMUmtum8WeJCklcmeEHaoqdimhjxgEiB/4sicDDY4M+iy3u0Y8FBwQJDDfa1
FTm9kxyKr6igtCerkLTgThrozH2DUnsJtLy+zWzlMXwZjtPMsequAzvDkoumOOPM
Y5k/H/vufEI8Y3vXEBDIqtgw5QRKGYnWLOf4K7CuXHrmrhqrPa7eflDEVsBr6Gxq
MRerD6MoJnoDMYY5AeZcaj5QTUxb3WKWwMewLqiW2N4qyItW1iyiw6PgqUIU/hnh
GcKctTKhsroCFEEz5XW6B/n5zofSBKRKG8AEQ6/zYOdxLO4xqWvd+gUgNFwoLgwK
CXbJKjEvfxsQWhReSaWvyYzfqGCOgcccStn7T8K5tp/pUBFhxRr7WD1CvFDlabdj
COcZRYRS7s9A+97AtrDBRz1C/fFB6zPvVSyFmrw+JMJZTUj/1EWZXcFkPVBfni5A
iA4Vb2Sj49J+cq1Fke1ytz+u0kqwCUBeGTpSO83VzSlzZ2nk4gl8MkBZgRpacct+
SYH6IxcNhirsBm/ULwMVhgYL0A+rdKAv4ithdvJtUPH3er7c/d6OrDvUSFlBMqYZ
EjhCVpIA6nG8ALufQSQoJKjQTCxHwx2BvWvhq/xiZNt+iS7slxnY5kJ7vw07GXAj
qJo6UhbIOZ4Rghap4bhIMtj8YQ7mLB1FBY9T407DRjDyy9qLtYyzg8nIHwS8I1fY
nRyiGI4NLnhn5uREPr/TJE/Axu4AhFu0NAqC5/dRwwpTQ9AykKuWel3D9LRSCHvN
lYCa/YbHaaWUUOCUHucYYgmWIJGoJIDs9d4z5tYfJZxxsPO20IUsMqEcoZEsALrm
T3rknA1HU/ZZWAt66K0yXpxgTNeTX6wGhZl/mdZCXEyqcZM7uWxFLGf3TIyTey8b
iuBzTD6bmU2jWk7+MSoejfE6BZao2WaLZnkoMqGVFz8oZBXGA7jjM5J0YIMT6jTz
DqMqItoGS4Ja1di11EiMer3a8UK0Cw55xoIjm7CCQSRSS1QVGBUxJ3Vd8Js3DGuw
+xX9wDGmPQEUmxuSyoQuiIjF90oSvkwiAKwuowKNA/4dnSJmdjCvoY8I/HUnMGgG
YpLFwp6b3YCbrX1OT3QoHqFaFqBHMCmAXBRZRZR/aOMZGn4GLvTrHLyzyIkatSQX
9acqYb0teIHcFyWc7U2L/xx72A/D0cnZR9OZIjjWZaQllcehzsxlIp8w5Zo9lPBD
ltugLiTEX5/rzE84f4en5As/tYR64V3hDT29h+oG3EursfhPiJblB1S0e0VwV5/v
juos5vk05Njn9h4/qwoIDBCM7bsMhbtsc/ycqrEtRCwI6bjEQQL4UZ59iM+gRdvO
bwBR80cSOFUYEbNLhvG1LjJO092TzP30vTQtYZ2Tng7gGLV4QIa1X23jOw8971nL
464mkIzVNcd/cs+R9rgllIJJotYqZH78ElUuVrsvpsNo6iRTKUzaFRMFeHafmPi5
ZSgfvz5uKgE4eIIXRyAkj/4zBSlZqp3U2+T1nRrbxUo8pq6wOK9ACVxFJAzz+PBC
wMiGLDLCBKNQ/6Q+c3pJkWpSUJ6nhZxAYAWXXCA7DPiuhkg04jd2uS3/CWItt/fH
K1Dr5fTKTHgSncox79tSWwLeqGsGc3aUWxz2R2ktTp1qdKhVIIo9XbslE86dWmce
TIxCJDI1JHWcJLHIG9aA08mASju8NDTlC1KMj/+DtAQ9fBv+HfyiUvKj79hQlMla
zu1hCNA26atOu+G1Cyromxz0yG6SQ7sRl/P2dcZ9a3xRPcLYFlyyeXZONMu/nqQ+
1AuvOjwWbD5GDItOJdLLY6rm49x/rK4eJiFOp8O0189MKHPA+dbaieqjoiwQv1aw
DSsXUM3M4BaBJ1d2lCswWD+ck7NWTJ+uScQnnCHw8BxzlyVJtEpxm9nUrobwHlvI
41MWDT9lf9jK9jUWHZMpVfhLKyzgOQdCtxHiWKCDrXmlVDU1o9Iiw1E7zsHv/Aoi
bmXa5f8yIqF7NAAzcEmIdmKZBnzL60rob5mWUZjfOf1DeE12luSwHrHlE6tslk4Z
E8+BvNdWk/mUEJ1ZapYjnqNJ1/bEP0v7r3oX9JPKPSfGXTu0dX0WQ1OouHTe7JD5
7YPujl7S9itMYcMbeScG4ImzNdCGiFdl+BwVj3be3agOF0FXy+yX0fgVkixk9Zyj
oGkO1j5F6TgBp0NLQpT195LV7e0vNYMHrsy+lZuh1+L9lcr0zv7zsoYn0l+xjIbc
Mr7HAeKytfGHp6U0jPS1NVQoJN/c9juk2fzszqaX9L3CXZS1Zc9MWeMsEz/v2iYD
0u/bxMfJiEOMPCutkzvHxxQ0i6UbotMFwAKqpy0lgZZHeHllRDXeKxVTh+CNTuwy
LP3PKOB9QLr4hazog8Y2kXwJVyvZdyj6dSodoeESaFxRvHty1tdbRgE/q4GEZv0n
nXMa2ckLkZfPLk7YBqhhD3fms6NU3vzDGmEmdxh42UQ5TWsIK/vHoGqUDmgs3Vk3
XY3ySQnCaAn3Kmg5EmizzoxpRKnxdBkOrshr3MP8STZMJHZqSolKozdzMvcDeYRo
kjnY69jY59in39mVjjBFrit7GttmHlM7Bw3GDDmB+DLCXJdzWNFa56i1Vilt/7nG
m66eJjJKoq22NI9goWpAkR2vEDNO6bzess0LEC8ZCDenjazHzzV/u2XzpKD+DTXn
KMI6pOi+8y2kLZzeJ5KzWD2DhKABJd69E5YicEidelOv//roOk35LG5mxLFNOpNr
Uxd04te3MxUp3eyAnfHJC54Y0roPiUCFxcS9DiMIiRSzP+/vXY8tqjU57pPkIpzq
elY4OuHSYMjohnM6NZi3srheKbGM/Lq//x7Qm6NhJhhXmEU1NyxtSDblVptYWWE1
UMrUr0C2vmB4Pd5AcNB8nHacb70Pw2/BTeD/UFXsuhTupDuJMLoY8OXD9TuNGzSd
uxGPr3VltPMIN2eftEecP6fgQ4kYSMMiPWO1ziz0lqIze9AI9c6emEpVgZ0L1Me5
N1RtrTbbXbCR19Gi1YjANQlceoeDBSfYZkzQdrBCkMW9X1wggfob0tumtBgbApov
Hz0H2MaEgYe7l6kNbEidYgRldvlZJ0hB58wVTWz7ZJCrG2wqR7/34tqijpuneGDX
yF6bLkpzMEjkkRr6e7bX91NzH9x0JigdxWiR5uJxYixJrV+klBoyNaZ4gXgczMe9
I2eGJanLrmkjBlYMJhlvBUbQX2oFLp8W+sMjNnwCnwBWpZrHdkqg2FRZrWJvJIdz
ftAOkxCwVNc/P/quC0rDc7ak+Er4f2uA48o2MKOb22XaSCbZj4XuitZI1yBLmAe8
KK8S1toGiGjNu2J/yr8wkX2iyCJ8UpgI+WPEyOuBQ41Bg4ISLcbjw/F2b76I/lyp
6F8vHh6PABgVBR5Ynu6NWi7NY+pId5J6ZpyzoLmtwY6Iuoy74F02OoGAj80yliGM
nFL6m/k6BwWCT6Vi2WzeVf/eVFpwmec7znYI77IRKxyST3s9Altli9ZLxXVkIJD9
OPaxmLuLlDVBcZFTUb9rLNQZTg9anU0d1MkRaEXvAnUCqTIsJ46nw+KOL+6T4Ver
0RJU3CvT5gaVrlMb91m9NqS+plfNOzOkOG3p/rxItCRG1qDl5+nrnZ9FCTkZ7PXl
DKR3U3+Z4rv/huv1le68A7UULlERg8D1/u/5t4zmSBu014v1Tss2mBeoG9Cqde1b
YWeM0bH4m+R0RrjB9GwmVyUc6RypUsfbVpj0bdqcdIC3VuIwj5BmYRapsHzM2ShM
6N6GftrjeYu6iUq/qaVaxOAxTa2fPZr7w9xzmyAG9+uFFedG7aKJXZaRglCSCmhN
bDYUMn4XMQRn8/madf1grRwkzkfUV27F2uCtsqq1oswVok6MrALi3F33vW+SV7jl
M1HXQD12hh6xsXySOOtVkxyPj3URlib8e94R2qlgX7hBHwETKLarTCFYyoRY3W05
hbXwogu7PIt4yHtoqTikrFE3KrhlKh+UrHgOBrVKyr8BRz+NK0Wj2KI8xuyPm8b6
7o/MpHcIDVxN72iA4dB9yWMy9+iUHzMY7259pCWK5z3Z1F9ndbo6magk+n0KNkvs
AalRfEuTp5BnBgISOcMI9lUXmulb+6GpTdQKvYDDWno=
`protect END_PROTECTED