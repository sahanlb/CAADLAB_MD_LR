-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
iZR9sIrMlA9wrEQp+tWOUZ4q/vv8Zt2jVi3lmhHcwA/vOtfyFfcAbYikROm6remr
s4TjEGR/mGIp6UcAzrotLTKFzClgnPEe+5bDT/1gC8C04NqKV3KMyBd2HrmIn1Bp
Q2r9F1G6gdV0A2/K7LlkGja8cDuCcusUr1vMUQbuWZ8nRI3tmrs8Kw==
--pragma protect end_key_block
--pragma protect digest_block
Z4fWgeeXe5Wc+gdJoHqelc+VRZs=
--pragma protect end_digest_block
--pragma protect data_block
3iN7ouY1onyzQLiXelUonf9zOLK76PhNVOEZ9eT5ahqUUtSIsyTeqKO4hn6aBmbP
whvYAIXap4c4ANExy1jSQvdEhodbeJeTSnSzH7aimbXyzSzhXqsVdji2kDMi55zI
Ipq+n/TP1fcvpfG4pqMqw1duBUQy/sHu+36V8uleXXeO3I12cYvOH5Tfw3f+43k7
VXcqSHtMwqxaTErHW3OWdeujF8x9YmPcib0nuTBh+NNQpZujYMU7ZUB4Q40VXKln
O4h7bjCaxyxBquphlZtdoabEpYiwghi7sqHozkUDf/+lpofPdrJKbax0kicom46x
ydfbtettEwlZK1VkJ+aF2r0RCc3zgrJAql2KJVfrJZ4WaV1rQgIegJJy2miLvXUC
N50isTnBc1hMPcPBKvqvH/mGDsByeLTKydhJ/42aB0glrJ4ep5k5KGiG0Q1YznUQ
Sxz4DKgvJTECngxCxEv+pKJ0jeDwenpvXB0O/yth3cDblybLadyamoWHDxRATcGd
qfIdQHCsmvD4qKP5zZ9FgJXEk7w1Z/ma3TE23ai31zGjjmV6+Prpc6FqTYYE8XsV
Tmd/BH1g8/JF+P5YQxp0bCd//WWZ7NRImVvq2oG56Tx0tpGb6VoFLZgrezF2TC1K
pfti81GJpmEmEr0Mw9J0koOZEfoa5LnMB44Q29tJgpjEseh2t4tB7Mt2CU1itNjd
/Nc2oUZGLuPOI8cAUBOr4uVobccSALwxJZ7c1qz/qfjb5ZGIV6Mjn0XcwJJ/Mmwi
CQQnbP76/RP8cNMinpRf4OQkFfyvR9tFygTmylTUQ67HvcXhijnPbO+aZ1dmFZCH
Eradd4VzHRvNI4p2UixuA1al3AM2A3giZevwzyff6UR6Wl+ZVw9NJ+8OVHJcgo+3
E0uQsjZi4nE4btmF7BGAGmLdhrlinsM2c1repNRSlf6+rEw6dmfXq92Us4bO3lAt
Wy3TxIf8iHeNCl0JQpfe2Kj66zweI75L+k1NHjvBvKkhaX65GxJ+6GYe1bdTSL15
98V/plVeVh2e1aGnDUeKtzAYKaAWld7X1VgJsggWCdPlHiFxPe/WF+8qXGIZOl50
RhezjCUHVUDrEoTH2MEnUsRozwVSs645xo7vseMCfqazTF++KykuyU6tLr/Rck/j
I4nVUYfDuDVTrO/vgGdJ8L58CtfXeRiPsyCLhjuqAxhYvHBPMfeFwt9TZRUKgpbm
DHv/cYiCBBF+0KXBgItKfxUAx4s9W9w7iFSaeHtKL2JSaf2xVIwEwg+rxa+Yq+4e
pFm4StQctEHZv+E1bedjiZiitfVxYWb4DF1I5AfqdjmyKRXPrhfQUQ8zpwNV/RVp
TLx7qcz/VDeuUte3MBggqDlmbCHxfS0lnEmK5eK0GXD96esWpZOekauwIdWv4QgG
pQmFJkBC2mutYsm93VWn2U84yA1fFTM7FOYBO8yRvfvbcC5D3vwQFwZzBUzP6wR5
0kgx3wd/5VwPh8POW+68AW9QMfoHYMwaZIqBLTLGfx60f8PoJhLvwt9NMeMOxBMU
XM0i6lrC2bDaxIxIK6vw9VwVO/1PXAaOnOLwb5aOGuSlyHY1TX9mDOHYxXh7U3ir
zK2dQrhQrCVmnsXXic+xcZH3wrRd8Rfyvxh12U1ykaqEydI73qv5wajY7t73LTHt
wE3dxb9aTQjpmhQ48mwM/HVA0s+jBfsWc4PJ5TMb0fOgM4mVADLTAPKr8wiKC2xQ
taXLHGmEPM69DHCBgtmIahGfsOVNCVd+fcnCS37zp0Nm9BuQYZKgVCXlp1842r+F
hd3qiaWBC02fSNGM0iUuoC8bOOvsZXnrU2+V0LVeIAWi5h31TMIhtiUeG18jdhEy
FUDP0iz8mpQue3LQHyqj+NpQcSjIHCP4V0A928i37QIa5ryyX7m83wHqkPytGAAO
BKmWDpFW2azFPUGK4bYxyOg3TlQ/jWUPKXS/nt3kdkNOLjwwrXJBz8fB2Lpm//3M
edy8L8jO1p6FRg/3OnsA8FMIXljzzC5CRs10RsxOoAjHR3VhEd0jyyE/IUnqFJTw
cJPIsQHCT7f6S2osH+TLYZ5VVuGv2Wg0gzDmLq0F6wwLUepk5+1xLX5EKpotWsRb
Mg9F/OdNea/OlcWrDsPz10Dao3UGUuwoxCclTw/BI4I+CAUD7Sf6APZVKdmuEUE5
Kqp/aTCHOto5vG6KunHD4TLmewO3Q8d0hHW3LLGk/DEao59CgDphO3geJ7Ku3U7m
Tb/fpEC7c2VQTbPtwrxonJ6jOxmqWjYkIRRJJybhA+EO5M+gYtdTRsrQRkCHTdhv
Ff4+8ToB/s2tL7SK6kB5vHMt6B1uZhCoP9xpklk0owVYQ16pGta+9/5EMXxz/5r3
BmnBHNaHVfuZshsOiPwqfB4YaKfEoKRs8pqq1jjDk4KrSQGZHkPVxHXX0KYOfkuz
4mvU3/zZeFr1jkKgn9rt+dl0onJjFPqyyHidxl8s2HAhjqwK9sncBQuROXs2VRny
Ve3agrOKKb+TC+RAg9+vuX9fhrcBVNMEH1tp/abELRxb+YJAXPHnosu6I31YvsT5
CfnNbeCoYCuysCSdIY8k4R0fXQ1ZQSylYB2yyJCHbYvchQoJIOkcsrmY/MRhZnU/
n9N9Cng13ZdhZmVPejWxk/l7lcEW0q0EOqowQw9M9I8tLKCvsUyRTbCtKldXuVwb
p0u11IOHMu9O7Y5W1EknFy4JdRgPqKOx+N/qs2evhGMr464xXJPqOJbhH6YLCMkC
//RCdo3mq46JIx/9sIZPn8q0Z+T4W0CSRcchPkKFOgK0Ip9ruR6oZOr9xWpBY7gN
ESmGvNCNu7vJHI1BTX6IUh7tJFUbbf6BGNewMWu9isW/n/niMPZF4rHxF185yQU+
4MYzTuTOs1KezZX6wCtuaMnL5ilai4+SmMfGVEINPQzMpWZ99gDF99bKHbafKn9s
44xx2WeazupkuvM8kO2cBU3uxUxwbDJ4V3eVFEGrToc7+8206NOUfuP+Qc9LpvvG
IeACwm/qH79h1XNgpF6fAup+zKie+nQ6nLq9xosj05laE+XBRPv7RZ5YQILHnnbn
lRcm1r16u+eQ0I2s3EgV2gJaGuyEjoJtFmecONxXZeDfztJiygY48ca6FyD1ZPM8
FlKPZmW9qU/9COmRJPwnuy8CbZTKRao0kXIEVe+JGR3D1rvFoPAT2Xoyh+R5wtmf
dZDlq3OzzRzBmsjBN12zF2Od3IrfrRUA5Wvb7/W9ly3S71WHnlxP6bfvY0YvXnLZ
sRaFJqbfJ7n8wNEAyYYWvqAJxmF00uNnoTpCsiVpB2nRmmZ4x0yfE74cq3QA5Lf2
gtOLoweVuZRYF6MYZnZ/Pc+l7PwPDlqShz7VOtzQOB+yJWQLI8F2/2xF2jDog8Eb
FYpGvU2qsrLXG7Wu3UKOIf8pjkYCD6jL3MaN2WO/2da4hLPaBfJDlKSEPNT3GtVj
015KKyXXzjUt51/15t7Psl3eIFQxYhbQzErxQzq7IZL2wswTiwYR4Mzsn/WMaAP0
+3y1vZCtLZszKM8i+iGWehvxMsHW9WzO4vTQWb577wud9Aq//+mM899fmSr+rLiR
5juDWRqhfxiFgoQylZnT5qKBUquh8M4jwGfaern7eilHEs7PBZLbIRWE1JBNutlB
tWncHoOSJO4zpaW4LEEoWGgFB0W8yIsS/KdUnqCEkXz4nZFcOMiHjgsxBDpaKnEm
NDf8vFX+A9X8Di67csMgH0iVaEr+6TEDYDopeMwR9vfJ/zJ0au8iwBwCtKVH6nyh
XnfmHQCnaEX+cRbvcU1f8IUbiqaJHn7DHXWfJk9N/0bMvW7O2WoItWQ4r8roXVl9
CSz0jXVUZx1/uUVC+pDbDERpVNodObiE/SpMPYTGuULDjgEm4ADkV3utjpwEf60f
+OM+4FMQRURUj08JspOc5cI+xpo6L/IFlzX9Rr0Xj8igzzD9+nQ7j5C27t8LOe7T
ufMk4oxDL9SnxesfPm74UtoDMzqP7/LgJLBdd3dl0Dp5s0eqz933OMfOhHnOuXVH
AEmYo3Xku3OEudIXP6cGJ27JhaLCxPrfBHuvGLS5QCgi8hHNLNT3VLSVawKvCEDc
O7QZ85+guC8wqmg3LMEA9HT2mJMY8rUPwJ2OhimPHsv/oMiTuvOkkEvHqdbFh82K
NmuFFmib9XtuVttplBUvCqXYnPCWM2KjlnW4IRmrP4lkqTHMuYKLvTz1sCvX5gXh
7NGnNRytjjtGaJfVFLSVYgDlDqdwpc4LQBx+dQxQ1AEqipyIiv8yMHtb2vmGspJH
C3MX1kVU5usFZHI/cjlXh5jwIY2ZRc+NB+ev6sP5UiOjGYCI/6Cu+/CIhzBbk8Gu
ZXphqGg1F8Cu8jeQpVsyGc/3HC/LV2IHDHWd1+4vPedCslgOJ2FnSe2lRQpAVSwn
+fk7WFBHYYvJRrFk4JQjYoeO9hKs8n2LriqZe+KXoNz3fZDEDtDj1+pcvmwhcG+/
oiDPkGIfG1OiT9S9z7hquJbUL8nYZRMMOtZBYK8qlfX7heTBBlhcnLLF8EBdcMou
3bTIKlbSbOZ5eDjWxaf4gABQ+ylVWeD1UJ8z964GC/UhQ6k1ta+6KE4C6SUMDr3L
+KpaUCtzt3X3Twncik36U7xGaUXQX1HXafG4IdiQIy5yDyfeALHv1ydn7FlS2CHA
RSSm8XA9IPKa6MyxTg6eIzQSlqX1oHeMa3zoP5Y6OAsOd4CToj5vBrW8Hi48O3Bh
Aq+eVxISLJF1J0f53Ld7ZqJjj3JXN0pK8VyTqImzOcZ0C/89f8Skst2ycvDnCshm
EibKP+ImQ7N8RxN4ENdcPr0Jh90a2HU5Pq4W4f7Pf5E6NXVKRzU7U994jivT77Ts
svhnf/u1nKH3dPKJZgrkVvLJOgTfam4qfM6jqkyhUsytSMPj8A9YXWwG/kRxOHd7
j2ueqIQZDpOy9b6rb7K3DCclIO6tZ1wTfH4vl6Qt+IkonJzYx/lYbFhbkbVUL6sY
Bu47TIkC74bM+8T9iM4jlxsC1r1mpRSV69fEWITJTH2gDIreRcYpWHG60JG6sd9N
rsVQw03Mv9jr6N9dr+uAjYVgDfPI+Vulxnlm8N9e2sbIuCbW9txeQQj/085xW5b3
Z+ab5di6OZNshE1HZynDCm4q/5x7qLDpZWDz1C2APVgcs0qYQCR1BFwiGLFRJIPM
F3Bn53RzGs6RRC87CsP404zPOVh8ZbQcI34ODBC20t30CZF3mcdyNEgzCeZJQQsB
qaLd8cvXuSrv/mckLtY+uOPEp1TxRM7U+bDxFrEHdGgd2RUY/o2CZDSgBXHrbfxi
RFmAGCY+z9z4NmHmkz4NCRzhfR+f44Ou+Z/SZOM/oXWHLSTcfwc0L0APj9zitfTT
KNuA2LcphNkd9yk0NeMJEqSscCpyjBl+th9iyFfhts/nVus4JcG333p9v3j6ctDA
zuKxRaK/Zur+s8h2sxYqcrxXwnst89IMtP7SJbiIe3WY1T5LAgcxrS0hARiKbh27
eBBRmcSNSZHB65T5wDUDpMmKDNGc30XAHxQ0AykWSFXRJ4NXI+i1OCtbtT+tuY7X
N2nO9E0Nh0rYeeoBHGolfOzr+FxqAxmAputWPEFS3l3rBpjq6qPdnQixniVXr318
o+SDmBj2ONRQV1KIz5f+NQ4lzMcZMeqYAi8toasWZGnXVZ560xirNEal3EwuafFI
5avnzjD/fygp6AOX7+oKjzvzyas4UyDAeQ3FsjWr1S3cG70fG70dyNxbD43q9/x2
Nt98XIFWbPafKpwe+pTGbe+NTa/a1YqamhDWUfdITKikP/smD+Rn4NxCPpwC/mqn
0DM0zGxQexc7q4+dtQowoCtkIkjU8OAuscb8rbgSOFw38E/oh8AcM8Ro0Lb79uBh
1C8YLqMdGE348YI9wfpwDT+Ng4WIj4MRMIaaAwukqyC8RG1IgrUzqR9pvNDgb/PJ
vn2jEU1geK50mBmel9nSmXy4swFYNL+Oo7Xv10PJw3pqwZIjo3gMSe5vsQBsfHgM
DTIbqgZRo2JWuQEy+9VbpQS08VHjwuq71AwLQacA9DxnTsaDcq2i/yssi4pT0MyH
+yHxLtnu057DWKczb/GNU/zoNGbJ3mGY+oln5zS/mmdeLsLLQ00zCafUTVwYPzVL
K4X7XB+dL2tZj2dXtXe7K/mmIbtQXuQASoNXY10VBNKpMy5uK51ThZ2+8sKeTF3q
Ld/8KtdJSjZxWh0YYzHZRidXNCt5waBj+Os03N97Bn4SYbfBlhK1PfVP3KT/Drhm
TkRcrXLDcqemZtIHNjvE69o5CEY6uYafgjI6qHspW4InvNTVEvZdcJ37JF09ayas
xRz6s9uGkw5KA95PQ7QQsgSU0sHiiLMU2RonL6ROAC2S0KJKc0AYy+u2mZBuRb5L
qwiMXJbkE/ZA+OFFj4h7TCH0fC4cTuijB7+IBAM0RXl66pDperr9kux3qBzYeqAz
jgCtDO0rSn0kHUw44uNI+t12Lf6rLep23l7SrbML2HPvW2soPJ4krlSkleSXtY2p
iBmgKi+is4pNKP0poVf7qzMM7yzhunVM/O61JC3tsmkPvSI7LBz2ReCBiWaOPHMi
M6nnl4M1dbgrO22yDZkZOuHMpOuda0UanP6/P9B2TyR20f/nUjVpYNMUm7QaMhhD
w1a92Vx75g76/InzsRfSZWzQoKQ5rIEGjvlE77L9gRn+wbHaFKy9oab5HWrY9ivj
kC3Bmv64lF73RoiVstl1l9GdlmFm2wgw7cZrTrZbuuD1b8w96f9nCyj9hRumwT1w
QTe2SiKAuWnPXvLUJDAs8Gx6krKnTAh71SGKaNoWgqVNJSfkqG6xkTL9prjf/C/P
0Ubqf3+CpPt+A2fAF9D/A5CVGpfIVOUveJdz47jt/ISDtmzwTy8uLxAQ9hq4S8QK
N6Yzjz9kZDwD15pVsXfcNS7DYucab/xXTNW2PEhhUn5w+kePBnYtsskbH3Tv9pK5
bvbrba9OhmMUaMYSjPhfyVLgxvxeKjnj+iFESZtYes1AKKLYiE/0Ap4kQ//B+LEp
VChdB4zJ9YA7Jy7+i2dBDU3cn9xskW8LMGxBpx9hWXX+8Mr3OCAxqkjFsztZ2VAd
FWX/8FSj2ZeuW9mNEc4R8A0clM1r9jDeWuDnUlrGOIE7s1RpM6OXZMmOPfpV5mOu
CpdRrjkxTnW3SFn7yqulKKSE5O7WTCllBq9Um+/CE4y/3lSBm00Aw8k1QhtP4dGT
C6HmfS6fsoYW4ed20IdXCnAHak8618gjwKpFoR71hJP1bWOKwJghPItfy8rdRD1C
7HJDpHCZdliLeZAaNqdifT6V6wqOTMSQzgI7vOrcVW7I/9AR6wvBeKU7mtSu2BNS
wllFo/RkgLYc0nMWsrV0nwz0UqqTpAcSFCsJ6vddMSnB6Lv/vK0GhL0izYii4FsE
qb9hNLNuKvhU7N0bg5KMcBI3pblEQWlTthxm/XoxLGBavJcKRMS+H88l8pGvCZfq
Hsmwci9XxiHisoLl53h6L2jJRV+niDKc8BbUBstqAaZCoH9sgaYxrxU2m4uZW4r0
abTJ/r9gDRtsQX31cKidZfdf8Tw79z/PB3vb7nhISmCZNOeaRxKlLUJrB6FUKDif
wMFbAafC/lvKh9nMcoxqatK4gErXhtelHx8FadLwKa9ThI4v6QE/5rq6ABeXRG4D
cMZg5HcQkW+okCw3s2SnZnqxrnf9Q6xziPNrIZOlQ1fVSg9O7vg6GZ0EjTG7GNdz
FzkkPjkfPHSauL55hyyn9fJkMj0fE7HCME5MKKKoF1zN3gJvj2851RPh78dRVh+r
1krGCjnbauy8odMcZX2lyyLhsFCyeDS/VIGtvXzZDehZbTcztjqsbsSQSs0X0hX3
xl+77zR8naJPrPktmfr0lJ8THv+HYbgdOAVnVouRUiQL+6xXOq3tqDWgIMdM5z1w
gCZlrA52mYPODP4dIOd4tTdFtKToEAyWbqVhZtEvbbE3mzZuQtl0thq8DpkonOLY
KTNnkSoZhAJQdd0XXH1vFwuYwQ78xRjp/mfKXiUi6bLHCSg2F/FTdQWihwsRWEUy
pK3a7lyzn2h5l+jl421Hw0FZZlfqDNgLMiOCX1i3yI9g1sdv7BqbO30WbAmpJHGj
mxtL8KDXnVRz7FjDLwsPnh1vBeMPbPVQLlky+n+IUl7DLzGz/dD8FTyXejv+Zj+1
2spYZKA/WZtMnYMyL8xY1urNIEYWfGeuGwNc1II+T4O1p+KiPwM7UEdiBQQBmupc
MDsfPrOInGnuuuF8Aof0qCTNSdvoLCr8IVuYUMtEqPgdruimJ3p5+LanT2oy6GdM
oQyS/X3YtPNo3VAHGOMo3IXoXtqPxJqIH7c5PqGEre6dXBBf2lDqPcc81AnsJecW
gjVZuObAE1t5aHYWAXNxxSKXyK2xm0MqenK6Cd7D8PGnXxWRC1sHyxtO4yhyah+L
WKrtCieOrwXaK98ah4mmGOjPNEs2FbVvN0e30kx+/xKltgNKIPwYek03r+bOkOmd
tSEtbafrpW22QMD+b57icrm4o3LY/k0UKyyIKDlW90qTEGCNomcRatopqhpxleqz
kgW2XuQV3wOyXs69+2Vr9RzE0R2qPiorn0N39jaV0sSMVus6OTXeBzrYI9O6Oasx
6HbhF4D8qhU5hdFc8M/SQekFbxkLPvPfV5wH/Mxy75kc+rxVWyeTOIU1fynucCVc
UjJuzdzqPeFwczchW29uU3fiDnWgvoRGXtmHVdMMwWIHN6F8ikLJLK0FtSgeMusC
i6kXKpeER1KHKr4lpuS2/grxvqcWGXMg9vmFivnvPdO/sF80t05SfGbo3o5ExNYg
jDrRwZnAAJidXeO/qwJfr1+Q1BacfSwmu3s8u/04JC03u7r4qKPeeuF7H6SEIEr4
XFEaSoLDNlxrMe3dwld0n9bB+eFellsGJ+Ubz13baodP796syl7N39VVO+Ic3qFb
C3S4l0Ixm5AoqPDZrRm0ZoEd2wKkJydApeFX8tfWBML9KFTUM+eHoQ4juTCaLYhZ
pO3m9upwjNxRCpqN0nbDQbNq3Q4L2rausdMZXpYRsF4UEt+sIzsNkEbM8H6hN3SF
RRvtvPrI977+4RZetVlSRGpX/G4hM9Gfxp5UrhkbaaI9YMMX+aCb5A+V73Xn5BPw
PYIGPZmIu/dVLUA9rsYYwh0lVwNfUIEfxcDxz0CPfiNT9GGOZyI51jQ3x3vrITi1
2dprz4J5/ReQ4/HtrpdU0SzoFWl3NRXq5nD7Aip9ZNOAPgVQhHVLCJGMV1M1sfSj
fLesbMrc5pNVIwt333qepjQvt5ISKbwlCIH5SjmL1vpR5yo23hKP6Gl8jIB2HeDG
fj7tdUSNaTFZeROssGAvBKxEpTxGr0y+dkbONaKP/4W0hYHCelmAr+KCEzG7X2gx
O4zVLTmXy2KTOZJ5cXML+9KMpwT/dQ+hVLcO7XMMn7n4rj0WxljEARviQ6hMMnLV
vy7rq4tjWCFOUVhHfzJTPoBO52qpwRogJm+33AVSJWJnnDwX3Hxl9A9TV4Q9mRn8
WcyBbZJvsDY9Rm1J1deKWEmF5ZlMcUdYWeD618wdRrS8SfWPC9F8lkPlX6Pj7qjY
1L5OoJ/96ADzTBu/tesLg0nxC6amhd3w5nwlWAVlW+TPJby+a/l1AwJor4/Q1zBq
0VrhicdZ30tAGmE1LG+Pwk45Jr4iGGoA5zIbCjCYWsirzafMDXIM7c4VhLlD17D0
pwHlKAb9I3jqRl8K7/M8P7ldhtZEKb+47jq4lDUm9bzMMceoRmNf7QCbU9IYJ1k/
mDWtGCvm8TuBLQUu6nxBXsCmQqfQ96mU3KEOtNCDN5MCCKgydSCGRJWs8f1Slbkj
S0Ee4WB6SvCBHnXatp1SpZmRjJ7IjU9U7D4UGThfwSNqPhQfulk8oTw9mjHeaa3o
WfDbQOF/IT6Gg4MMBkdCnvQREYVrrpW65mMIixJrtH77i+ov65noP1tj55+ZWJ+g
GG4x9Gz9kq7iH9Ln2AqgXIxg+46PgczQ9d+BzUkpVXTMvn4Oam6QFXYLTRaFlIp5
H4Au/eIuefUNRI3IxMeFSLrz/qAeuFD/P0F8eIDtyW5M1jxHuotFv8lfIhOeDrJf
AhbWPI6Nejv6kf8Oto2X2h0rx24w7nU5wAhQDc7ZFEa+6a4foOZhI0cNSgb17ErV
N8V7OJcY0NKNtpe/C/dH72ac4yGmtz5a87QkWRFdyzrpxAogvhnGJ4bfiGdLogKW
tdjIB8mUwPTTNPmXPjYYCpwTCK0gGMGkejVhNvA7xdYGOSs0HcccWOy6/OQL2u57
7SIbF/dAXrQNSxv7FZ+x6dyNCydyUYGROidlIO+N0xRsmkLq2Fm1qZQGSAKLedWV
UPKqYjr8hBSZfeLQY6SbRAKuoiNp6qptndhJ/4AzL2rk1JmmgXaH/o+sPhG18mF/
GpL6nriqIHQO5asYXkXJDoSwVY4V4x0XRLxQAwZGKWswsOWdUQf7FNGMdQeBdo8s
TYdhll2hEFuUDmDAuDcmVYQ2R6WRE+eKr/wPg+ouxbGjxfNS82WeMlv0ablFoZ7I
hPPUIwciSjRC5KM/k55xiGYuNwK0TNtBcg2iLWgC7bG/WU9n4jPzE39gYGaby5T4
GzaLVpr1vOMUOfI3ZJtFIH+6n0BEknTDMH0d0Phjfza2tsM43Jyz3xuWwYo3NMKM
jBBsPmPWDLwUcar7fzmetFCCEcQ1K+O6TVOwdvgFSriVJJyksqF4Du4wYGu1aU9G
4b3HTzOHeCHghmaFhBhUstpaqrmeS/BoUYq59PYBQQcyZXnk25dGtOmVx1vZxTEY
gdx0lcjcccLGcNtOgLXP3fA85bQISdU49Kx2+I0ynOBd7UbUKcas6ihfukdFR5Bm
IP9NyPRJaa/8u0lNZQrHix1L4qVY4Up+aSjEvjCBUr8df4lYhGJWFMsDq3g2taW0
28yc0JRvXHYL3cV5VBSiFVI67BJTEip6houB35CsgRTk+cCXLYM/nK72UOgxp0BZ
MTbFAhfbajtvJadHsPvbIvsv1r5Px9fYjJBuhAAi8y4x9ETNFyvJIgju8mYQgm1r
vNI5soPnmK0UvocI3C5FjAbBWejDNnwhHtHIV+kDxHBLaVp0j6TqQyjphgJ3HjQH
S0JHYoi7w74ygn7Qg4kwdO55e7gqkgD8yrQnPUbB6M8+Jap0c4lIJXcnZnK+bZwL
5g/mswf154BGeTI55n5XaSkYl68QgCjNGEPI1IgvhO4JeLMLtEvSPnUtDyTcpIwr
tvjXXxNmnXAHyEtCoCu/u77tKP8p9EjC0Y6JMunBoXGShpyTFvzp9Cl0HHGB2MLL
nfsIyfANQ5x3TSUavWAJ1Xfq/OblyI3rXFDv9zLtQGyeBFbYu+qaRBHe2FoeTkqY
ttbV9riNlKKcxh90U5HgymK5h9agnuG9ugP7CGe6p8kWbMYR6uWBE1fh/qfRaQTt
6+zdAB8LhFZPuu/jOdOaQP8Sy1Qe13LkHSqRhpi7wuTnh3TmqyX0udJwZchpcofE
tmZSsi9BBe5ubO5gStppbQHchciVEV1SRijtB9ctaJOO3+SC6tr/nW5WBmbOM19k
jO5+0M/E3bX+RYxNJoU01/xCO2JJqXYV14ucROjePChryEUKRSofEpOHWD8ASPrR
cz3KW3ty0KvLyLXBZsUUrrwXtvkUauy8oGbDh2SebgwY6f6Ss9U4VIXNuZCkHsEA
lyIakojt52vztunJ/a0obMKY/aPDLQXEQVMLUU2wpf9HE6sqOUfzMVKIpBFCOnjq
ttjfIDfdWhFN+l8ISsVUJ6TdJvcbi+IUoxaf02FbRH4+mMJ2RNLeePaswEKUoitG
xqoTAnZX3V6MmfZlTYuHr+tLuAilLR/At663aBd3h03lAWbH6iwmWDzNUA6nt8W6
jjTA/2qzeqTt7L+qdjBbjmLWPC0rn7ZUiWIJ9GxwUXAPSgc3qMVVm9k3Sb6A4VW3
jZI2572yV2FaA2xZ0LlmQRUTxAwm29pRrIloNR5bdbINb+6UaGUpLcAAAkIyb+0x
LyqPWskq8AxKgdmaJZ7VTWJ1+zzJuEQ5E/9zlpZiEWQOdfkEZ3zsfOUUcOm/plQC
CA7aekFkXxejZ3+A7Ch3B8/ueHJ7h3377gzK6C/1oUeNFLr+a31JpdrdHp8wBTie
ap1Eu5WfnBWkZNDhxJz6i30nB4OmVdJmawtZUL8EEeCOAxtBq4TEfy/M6YXfDXr9
ECV61ERTFwzSWc/LHQDt8UvEmFo2L6kTzpP+gXPjEG2c0qzQIrd1omPHXTab0Iz9
ZvSkkNj3r3hv5iXzOwnf13IPO5CeArbDHc3rRD3OHoRbhvo+H8Z+hzkarnO/Xj7w
JWeB8WuAcjE551ipztFixOXuEC0qNW7qdkLe1mcYwCZOqzVXOlBIzyuMFKdGKDk2
kB/ZG/+xuLLmlWj9hobOMqUPO4qW/KQ5pII5RQBTUMsrygfD+vFq9dvqplDSiTCO
TJz5Nr0bbE4VvwlesO/nMno0tgMeLyGJLTFK1FxfbnTAKyZPCtMEyA3ZWF7/YgwC
vCK+nuXvoVBtSecfd9WNmEQMazIvfZ+y2z/0gsNKquzKI5j4TyKnQRU2BeqTVwOf
ZZQIZDxElcbpRoz/R/4sGovOjwN1MW961Gz9jGim8zucLgk0HmLG4DfN3SYw/Myj
peltb4nbJaAnznF+lAy/tvbcLEsZpbMqG4NxvVt3TtZwcmwevRNLZaUtblxQm7l6
+ycWebCXygFOl5kDxxjMJ8rgoDf3nAyzN60l+nDoHJlO88Qi77ZDHX+a4hcSGeIN
tDaqZnYEOLqbH/NnfOTjTVBneZ2oL15sUx1kdxSjC4cIQ93ofH+hjDjj6Rv/1vU4
ibEkNgorkJZswRQqNdNAcperEDEwytSkbIP/JVM+YDa4Z3+ir9T9lWqLu1NblW2F
+3IyDVbA0Y5aMIed1xNk2Wi9e6IqwLtvgX8XyGB8ZyZ1qGwuy9KjUoJEI+UQb4bh
poXWXB93dGKeJsiNKMuRRvweWyn4KVscMTUAk01Umkvjg19RkzrmiQofbKZJ6Pi3
s7JFtua8gVgxVi4p9m9Eu0GbC1ncrEV3h5yxCH2ycjkid+F7FbALCg8kc4nczkGp
DtSOGVkQm2blgAdgq+Wy8r/T1j/+q+Za9+walBJ6FCLfTCkM79l5vhpV6SZV1DzT
VvQmTsLXul2yS9GwX+1T3lWLJVNpd5Bl0O2a2JsJkjxnXlcoqtrxz2l4Un4lAjt7
+J7msY65iUez2fGUsCvmsuTeMCk4PbHgspP5OD0gDsL9fl4DRR27RORdkabyVnr+
ZjVNCgXH9KWNmfJ8JlCdhlLEqILjVWRHeMBvB/qkdrxYXMrVBJgA/qFmzqGyVVaD
YlJ0ks8aXgSE2NKMz0Z3L3QnlhL8AcqBHHZuZ37nVCrRwOzPrLheAs1rA798iXtw
vuat3z2tPoxmMKVADtDPxw==
--pragma protect end_data_block
--pragma protect digest_block
zfFUoZ6Bigq0jgfNatx5KV68N48=
--pragma protect end_digest_block
--pragma protect end_protected
