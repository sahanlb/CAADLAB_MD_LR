-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
wWs8GNsPeDcOU4sSJ7qz8chi/MQRAvTm+zRs9mNgoFekaJ7KUAGdNYJP/WBpsVlk
L7TCCjNpuPNJjWOiA4lv+7/QCJ8Vo1RgbgkFsVvbFXywSSkqzENQdglepxYQoZpU
OyZPZoH5PMRDC2WUUC11XiJcBn7H25ABSlWAECJzCvI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 17136)
`protect data_block
7dArJ3v2FbCjvqfWmFcxvgclT/eCLCeeR6pq1v1fAmUntZ93puG9ddutrCBhXWTl
Edk/fgpTXgfwC157A6rOrRaFKU25pr9sSTqtQLVysL2yFMQgggqdVb/hbJMQWoZH
ACI1NZUUZZU15BgR5OmgDo+OtT6VmvQodTGJHqghVAXB/NaJaBRwkjb/qaP6nAMn
XpoTDRTHfh+00MRUuwhY+EGbiCmwxjX3MD5xwU3Sp7QOfOzQIZecmpleZHqKyJHH
ZL4HZPZaL2dBjxR1llfcZKGKXsUFn5BCYHFOpwYjKMNkxZuOHkStGTW2Hcecd7br
BWTPYpOlD9OSnckdTULbzh1eLoBvRZ9cjpB/kPiAv7TjOrcdk6LtzCcZ58d/LcSA
cX7yhmvgrY1gdfjYel2E/MwcbDXGTGaPVNbKAiA2Guj/xXz7czDtlNpQBkOvAtIy
LTUz7NuUoAIZNUJRyA/eMoVBtxYY+xfOJGCd1OqwkwoxgHP4xl4VsnP9/N03KhWI
LtxzDolaPAxxuyYfV2ujRpBn39HW3jOiksIvLJI1E/1M8YqN2P2YcxbCcAXKTxqC
T4q3e8d3WUkrnfdrgSs3IiZaHmvhfe95keNUtegVlBaKeL7QrxHB1rdF5FAkFGie
Ng8dYvYo1C4LPULkmRRfNd5gCPBBQGo2MiMkeuKcMllNsVO3qIeT4TE4Wcxbz4JZ
woWjiVXKLqEyKuaJJxwzfNroNhXQ7Im5kbo0MDrYMw3aWEmSYbgnDTdNeS7qCGKH
3wsoAfIPCstKlcAVAo8FYmH/e8tlRRYFqOM0wg/+v/fdxTZ7mdN71mLh67eHJn6s
QLcxO2N/ttb9kRSk+H7lA0g3vJE3PFz6uPXvy8red2XngvtnWm4r6fo2rcE7k7/M
YPz8MUYeCyYRpVSVkDm7GVigTcA9xiF0E8lh5+y+7tSc+j77iIGHWyLAFyCMV6Gz
EI15IL/wdqEzF6h5qDDo3f4HBvrZjw//hAdbgFQNMptwSkQnTot2xvAP/YNKgRu2
fE3+bYVJNCiAICc0m2mbpKOmbUXC/9X6ZfAxAS55HT4RfSrJN0a8DYTfP8zNNGvP
uDPCRw9bwx+RBbiPRaxT/j0Hg18PPYC/+wD97K/mkPlmewoLvl9JenSdqM6wvnzS
uA93BAD303768FoTZJiaemHCH9kb03w+au3IQBaJmg9oUL+8RkBblNyukyftb83F
BtCdWsRjfNDgqkQ56x0ZlOg43QF9dSjQY17hqlTFT/R3U+mntdEwGv1YjOiS8/OX
W1aDgVRfJG7FNLgJl0y+qdoEv/G9aD6SUNx+k28fKCOOfdBa5d/eNdFWyxtus5VE
Xr4fGNDrHYbJ0dKN0uhpsPZOZCbtdGWZiusTRI19v2JJseUidh1eFAj/0Jc76Urb
fX1PUGNxLDBVjYnlPMpseePIS3I1522PXfYKg6HHftrPyBpZH+5tNOJkC9JIapgI
4Anxeij1vQXbcgqNldjdCiH/yU+1/WVGpW+CxRZvuM6iNxGIt3TbN28IkIVRzAf/
3FOvQddHPdQJWyl5gMvOYATThjbmaEzzbXpDlVs4nuCJxQT4BxGX2EJ4qVIHMlEP
LTTDswj3JI3JsoOMVcA10o1Dg4db8w893nFw5qPGDIAMYcn3k5ABAlIYZNAaCPgk
U7hhgr4e53sFEKY7qyCkyOQRrpz3c5Uu+T94lDlTVnb4xmWpxJJ13B3/Svtcibna
MoSd60SvcOf4ZcL5WPgZ0b+sDD4T9wkbW2qJ3r7Y/vBCrAYvpNloYK0nNIsPxbbP
FMIoA1kJ31vkNO0HICZCZMzxMNyq3XpMZlf5aMgJA+wXmMEiMazUI2Unxd4aBC0n
MjO0+GqDT8qy6mchwXAvWG1lbZtQzUf1pfLIdR0gUvIH1hdOuEixs8enPNSldfgG
F1qCw31i1pFCpYK36r3g6Y9x17+bWcMC7eIEVIRZa6Zhn141o6jsRLKnWPf3L2ie
vOoLugPoCw+flq3xQQIHmysdA3HYuCUHsW0CKgc3c+ULvZTroa6gkeQrFbQR/STM
OlNN243ufej5Ih3153tO1yiL4M7Ghy7mT/tQ0EmZnyMpxk+eR1qun8cnrl9KQY9j
MgZbSG8yD+muYx8Qq7xFHlPnGb5HMzBcgpyaEHhUbd2F3+xIxCswZVsYHzyB5ndu
CuLqBAbYq6az4BK5gqhANlDJgyYF2ikpTNMi+bwswUE71q3Y4N8PfJoD8KAAWOuS
mXnsvc118BZaQX57Q4BSAc74ID2E9k8HO5CJHsNj1BCh/QKpOmg3H0Wnr/iKOmrN
h+Ge7TGAZjAvl+fMqNMafb3ZnyJVcU/gF2tUrgGFhoW2Yk7fMWaaNiWk3tRErugz
PGu8Du0fZJavVywFxCa9wBKHs1RBLRoCdpzHB3LR252jsChI/58XChH5lo2UhRgz
SqXcFesxveT+Bq4gAr+sbKaKJYlu0q8saoqo1rrbJ3MVWh0mc0O7qoFqE+yZmgg5
36okRjQ1FckU+j0av7rir5H6a1TIDRT01axtDR64PLeE1ikCMqU9GXnqL3WoyeHx
RM1FEcPfPjEg0fXUBBKS2idM1P9nAGPN6z6y9T3dRT7/tqsAh4zsakYvy/kcAQwF
tLI945pBbbjnK0O0flKv/3lQEn75M01XgTRqpLZ8/QUTV2X7e47PRZ+mo5vS5nsX
eMvb+k1cMcUbS/JRHhrdomxkBpNWa9y4KCAxkkiAuFuNyxShXUCuBBKNMjxquTtV
xdfaa5E7JudWC+zM5dplqEBUvryg17sWqwhT4kFG8kMR4s1rJUVeOmqdT6p6btl9
asZ6y93Ww169Lf/hwrcS+Zw/EMn3PdZJ3nJvTj0T5YUnmee56tiqGrr1CGGhu8dx
oCMXACUTVBJXA+D5rYf4D389GQSS1R3aMX3kirgg7D5LNK/xskZm+axv3pumI6ZL
LF0o4o2s4t16uMjG1OHa8Vfi+49aoMh79h+upVqPSNSoRZC7JwvFTrH1I5aF+Wjr
RrLsVO56ehlswgqr+DdUZHq20xwb0Ggxbk71CQ3XtOs4QvKKs2TXm+Q0vsCnma9K
HoEk/Nul/+Q0HIWMMGBt+wN7R8liesESIoQsOQV37wShWLrx3R4ACUxk1vH4SeSj
rSv6dM208pD7qXbYD0Mt5OQSrq7mlL/RHsUFQ+wfz9Pg5k4BW1JvbuifQKbyo6Is
bfYDDqeSGEhC+igIHCt4KCVbdDUHOSiS7mDwemC3VFftzJeRLMItpiOaT7ksiAOx
bKSRQU/CuT5prOh/gGT4h7se6FQGWRufVj0b5Mw654+3N05X6rZ4fcomCGPA9Zwx
/lEQrREt7CnkuEry41AXcM084eiIUtvaAwDoxrto97UkLC1FOJQWEtrFGCEAmKyJ
c5jpFYExDlCQUvmuft7wgkbM1cKQPukA3xNVp5DI2htHuaaWauVMEWCC+M/f8VDB
Gmo3bd0iYCSKGQJkSb1bnYshh0st/HmIjbCCg7f/GCg4LrzKYV7AqfQYKIPugkdZ
Clw9LcFuC4vIicfEPHiLR3k/hAzCMzZ/0/QFG0Nnl9y/FetmZK0M7Iamzv2R3otR
HhRabaEzPGM3kCvZ/4NX4LHj0dtKGnc8yGy8ccu8TlqdAEH2xbXcagp8+5UzsQAU
gs9DHgfsBQ0rmmAk5EkgB6sU4OKTnZINONhwP70kr0+LIvOLaUlCqnjemA6wZwec
TrwT34LAuEs6Jsah6ke3h28YrqAylf44xrpByor2RK8M+jdPL+UzZ3ZCqivyAwiX
wwBibxpNMujXpT94YOI9eXe7c1ZAeDLcsHaId2e+LVSTougjyCCyarlFTV5BKVhx
ILDHm85TuCj9lououDL/t94tt6uoCdNUWqGlMrOMTFiJA/nyKCeMdIzWu/zvJMeD
rm4GU1AOpkbdPW3XI11Plj3HZZvlvF+8CtlhbIbBXrlvJmlX/An5IqbdCLKfffxS
doU/4IEoVIriZGHgbQtkM38DUu1tQKXiQaJXLori1xrK0haDRU0lYx5CjFqVX+FY
JohivWihW4Y3MO9QZrxXN7LIbJzkzLmF3oZ2d3bdgeY7UoDP006MctXyZHKdYOoz
4DM6yQ01g7eWn2IcOX7rJzc5I9Kv1N4UA6Hl/ngjSxqab4Lx2QUHWatAuXEuWMy1
S1Qd1bbynzhg9p4I4/s6eI8rHZcnH1EKsS6ApDKN4GazdIjoPpX9umWQoLd7kLa5
uHeqp2lMryLOOIJervb8LwFp4L04cPbovjI6EBxila94GhoKRmN02po8DrH6+v/j
BwqqJOmDyrqEFV6TwGk4cg9TCvNDeJq0HOqR/u/I7Ol0ybERN7f4es+8XxprEOYT
h1hjtc06KmPBoyRC+0TKTp5MI+AmBo5ymjTb5NbbuiVUrMlYkxV/cw3YGCLAkAkO
6/bh7tcFGG77EMGPc5K8MY9wGdpwbZtuxKEUpV4uX8XtcXp4Wuh6Gj1L4hahfaxP
E92MzvSA9UOfcimWGwEMawZ6w5ahF5rgNTMKioZeSadgoIWSW4IvhFU7Y0A/k4ro
S7V50Xy67M/vqTdNIdCOd+sY2mBqiqOOE3tfbvBuDVmS9tsAR+JE98X2Vn/PAONR
jINDGdo62nHvwPYqYAXSzA6mLF2NPe07RW2TcIKNorueDlJjrhEv0Juh3utXycSX
xUGCoKbmkOsgEpvfc3AXEgaeFJffacnRQWvyeo4YMJrKDy3fLGxoF+Vf1Gq34W6j
7FoJJWySMF5h0+xLjGl76Z/eiIu13Kmf9uxOtI5mmqGYJn7DEeQXWhPF6VljEm1G
JymfjBQHLNFMZj6P8FqAt4b3Zi1UhAdq9TSw2AFrQC3yPrq8HYvRgkq8WnCoADqw
qzRO6Z4tt3uHq+CWet+qLjaIkDu6wcXi5taQ9MVfE41u9kTzhALDF6HBQeekDLIn
2EbMPDo5yzrm5GiEyJp0eWtYM6FItvelRcEd9KhJ22H93RDFRMd2jbq1XqbQjTM8
Gg97v3n5kYXkF7WqA8aJ4UrremaCKw5lzEdur2hKCGJ2H/bNm7Ln1X4kOw1s2m4V
MYfeRq2Q2QXfkXzlSvxmxjjMRZVyaG1Q7vld+gn6Hu9l7PDQU/DIKnF4XiK0mykD
AznbEBED2MgfCXvt2Pq+CxhRO1REaydhKEpQ8SLRxF2klrYqizK9qk9pnX4ZswlH
t8cop4UrSaAGzxuaamB4Xe6alYOVM4COEOU9ZSG1/mlpM7VTWcvTztKl1jwkDkRm
l8qXVfIa0DNggFq6bLCpHExl+H0dnnOUkVfcjXnFXlElxS/p6rKRSo1UysuyfI3w
ay7wzB5gOVo+4QfE5Xq4q/7G4RREs63klketH8J/p1On3MXMYx/jIt73OF3OgiKn
FKwuuyng2ZwA7yl8MkEYAa3TOO8m1AONJveh5Xl8G7/KU7+UKu7uF1Ckpr3dsaCc
wB4gCmg04IIfWF5eAKLpt4puBlvJQ+e3xiM0YC7hAg+Q0qDCIMA0dkAWmlHc7/9V
BlN6fUHHU2S+0Jz5AWD5uI8nWdv6lbQn1PbvL59neDvwbAo+0wN443B6Dey3R/fe
tGALDKvz+MItDlW0OkZrryu4FEzGBZ8V/DWIZBrzWfXweB6vWB65J+5TT8g9HrIn
Vi0LrqigAuyPyHZvs9NiYHgLMuKv8VkQ0ixgBmXg3TBmzwp2ufaORr0UhwioQsAa
N1WKzT+L5ewNSI6oJjNqB+kjwrTihruNVEFMnbJKUD67W1WF1LfEWhlo+BYXsiVi
b1SpdjKexGQqOVDUidEO/NkB1eX4jvUDwYrRDTtFQwq/MvSSXHP4zZBDakiBkajj
nObl5TyL7tDxR2SJMWKKIjpEjr0gEpKHNpmrwgoTc7jcdXQeT4HNYeAo3X1IpmD/
uzgC5mnxfabLDhmMJtorQoeQVmsRbmXSqMA7Uj+0kATbahLy5ko311+O7tXBxL4l
fMmr5g7uOnk0AKKyUfMzgT97w+H5oc86dLr7nLuOU/KoVSWThBTU51a0QYpf/fN+
wqYoivYAPxPdwmddr+L/geDZyGlX9Dnxinfrm00h6L+lndUpDxbGSMs66tlHcgMx
X5a/fJUqCt06wgVpaPpCZ+q0VwexoxSxpqCzQQSo/2n3lku8TjPgd1QBqrEDvf5n
1cQODvkLDCWyCO9bn9PX5uI6fw1U+IzYMN+LjFPZsHJil1S4SrXxM9tLHAq0CWP3
GlmJuYzAyn7S9prV4nK8IB5akM+Dt+LgZI4gXXsGkAkIY/G4pXZCfL9GGJuXbo1K
cdUlCmsLWFCooNERXWyoBoeJeBf8OnOyYpArGMUr7C179eSWemk5+ix5KRecsMpX
HL2xIEHCefm8SJc9H0+0nztJqo2SkK/0u1fygjx/SiEu/9vy5/WhKnPsqlWUzLaf
rToVBTDIDKx30vIBrWQEtcqXFjU3m8HRNrwcDU4whHU/EYw+ZMjl1U5UMRaOJdJ/
SAF2/4y0C+W233AshIe+man1UF/Ir4ZAoQPQiWLkeAoGB3MTHhqPcLvbMUacuQES
hgdFpEr3z0cMX4LHldc8OPKj9Vx4TeAPMEZIa42ahtQs7QiQC6xTevnG5d2qo1KK
xr1FOE4hokWe7XSVDFxjePZt/+3Q+UOztHHdkeuYA1MVfR2ETA6hudUMLrJWu+ao
ATCFP21VmtyQPCR0z1JURn9ZcehpnN+D2Zj7iPZjBLXxTPrbHNF8AGghhYBH8wce
HXsc4DJhtHnf6rCMgHgEsSlsLViMIYvy5j3fDoaFplmZ9nb9PbuB1YXCJmJIfbX+
W6J/RVmXrc9GR61eTOhbeJek8jvg354e3CTjo1jlWLwgzQMWi/RRkTg49/svtguW
2tSfbJov4zVCTyIHxf4iQGmM13yHYmiL/UhPWxqWacgy9P/dR0Y5D5fFNDnAxSKg
V0s0ERWX6SHqFsZHVQOoaPHaIZDhlByRyoAfEv7wQVEQG6VkZkkb0x7ln1447N1d
Dy0fLXnNKZosywSqDs1Es10rMUjzbcsQ63kplJ/xGh4aPauZ8pFUwU/nPH8ehwFG
YMsz77DL1KfcGuUIZfKnSKU/pJ1jSfgdeH0usicovJWsUuHg1ngj4AbUQkIYgNEN
hNmXNoSUv61X8et8M208WOz0+CJzpBf0X0HzljO0Zs9uSRF0x7qa0vT+yszQvXiZ
dr3Ug26qk5L2y519Mf5E8LwRIMhiRziW4/C3e5HatPk8vj8T63pB3OwTZEVBaiq4
9Yj1FmmQIQ6ZA1jzboB479QHQx9sxib0xcoldG2Y7wWG8QKpF6+CkQnSBzJpNN5J
MRh7D+0KMEc2aLlyaH/USGXlun9TWZlUBnL8VL62MvlxEISofa5xO7QgXJr4h5f/
ybd9TchQhXkcG/waQabOeqpLwhXgQszoTVVwj0jUEUfTJwcnuprAilOWq8dCKZ79
NgUXwAWz+/zFGSV718sHFx4t8YAgGmAH824ppJjfT/8c7VceOVEoG+Or3wETzwBJ
GI2G0XUGl2rUGlNhsLR2l0R55HeLGkoci3sK79InQ2pb++ljXdqpQun1u3oKdtRA
imPv/EXSwuaa6xNyPnUpyhSR16n64MpN/faV1X6ZmpcUtt0/VDhofRyrT807msVt
wnipfRQnVFOuYc3jBara2fAX04ftY6ovtVBLsm5CyTEPg/aWgkG/jNlXBdGOqu1g
lO5wA5oXTjdLysVHCphg1ZiiIW/IH0zWY+yBxi3t9GBagp3/44V4sZTWJAvJ1kKn
An4GSeQxkgfuWt87f/2TLaq5Mi/NMt1uqVD69THqYcZY+oOSzZ8uABwbkSfHdD0X
sVKGXYMP3zm0aos7ORWPYS+sZu0bS+vxydlsiKv8I5gEC0/uhRoVFSIbJuQUmfkd
VdbqKZDGx5Njyl6Db3lRBUi19GuX4/mm1r0boHDrpIalLhVJ55KzWF1lqxm4UNlS
4cjugy4R/jaQ+6DyJxKY+ip/EB4hekTbKlcyXt8/T2o0xJV5lq5Hds7cPGfTvUQ2
BWZzqJrk50LZi83sGeN/K85h1isdcd6Wt1eDJO+3Sd3G7tXcUN88FoSzSml/YE/6
6yl0Xw8wWw6xVfAJpDJFIwS1JpAbn1Y+t9AnsE+EcG/xm4zv1vgFygm597oDNcm1
yCBhzJ8MJeMTCiC4rn7Q5nhR3ptfwBc9HJlYhNlv8UnZRRoMaufla38IMS7wPaJz
sIM8qCf6aj0kG+QdJeBBPVAe3J+i4akb+NVDZaanr+a6no/REYnU5EN45ehPxJUE
N/scau0rtMjED1bJ0C+pU7jSUVFvaPeoe3jhjLwpTZE9lQTy1sKp1vFVC4NqNlIx
BmOcNq1w4G1ETihJeaE9KDp84f17ZHNGTkHxkiTsjZ0CBebZhpi3q7RfwVRWDnKO
2GWTOpuzWpJKDGzTqjn77G7BKTmIaMaPo04E6GIoekACElDgL7Bozx33B7+kQklB
X6Y8iER6KFexk0T58eeSgMq7tZY3PyCiO7xeBosnfy6SfJ9LxYouJ5C6qMukdBK9
d+ekK6fMHJIbDPsKwxkw0idqxQKqZQ+VPwlDzYm3WeeX5ChFxgi/P2xq/JlJkQYz
9jpwNUZyt4ae7m8Tu1AtqMPMYVfzkcDK6ghCD2LAa6NXN8/sfGyg0NqVLOqA7ae8
7Cce/VPPX5Dq8dyObo7x3DY+VseQEPRwm/W/MgEPiA/GRpKig23lnYzJSuJLxEap
x2OgSGEvcAGeMIfZErEjw17sndnGPnjhyfXG0Iyo3YjNyf4xrQdNb+3YBeIMJZkL
K2FE6IeuRK7MYmw0SsYCjZbzIl64/Koui/auan73h5IZRuZDhDuNr9twylDxNzGj
59zT+bGG8j2S/oO6LQE2p5k/DvxI4RB2isSLaGw+TMAcHZh1TlxM7uClIy4tVrHv
YxXIqzq2AefUX3MZaSjBfSqugP4DCdXozj51JzcNYL4t52lIc3J+UQgxN3Wq79bn
rA/Kg3j2hcNzy08o7C5MkDXwYcd6teEkFx7NqJlguu9mro8I2vPRcIE3K3wesjs7
G0KoEZWgG8LC0BBqiNIR8CF06QVYRdLA7G0VfUWKiMq5+cRKefwPOwTqbJ/CcVxZ
CpDZ84Cxt02QcyiTgc97LadlDp4cYBKEC4AvFrJHKplWuiAfu+us+y7piqgFbOcq
zz03DGZg1ZHSnB5K/1CVkAdwP0Ek3KrKKIta4yCRW6H6G47nHaWL1JDkOYHSeEng
3SCvA9379zmSdS8cT0u3b+riZEYtisyUx/rcs7jTujXtcmIyWSs0HRDZfG/UEUzP
y7aXD5P9IRjWU9WtoJQpNKTr1ptHikoidT32vgqUD3rzRRCInU6hxgWgZtelzPWU
e8z7M68d7aJw+zLm83m4xL5U+XDsbFbrYxrqJ3mB1CtNiolta0gLs6Q/UBqHQhrO
u+LJoqNRliSN6ZmUFZI+TRhkUCsne+XuFSavtuaUKhUORnN3nzEJx9cCtWMIA1ym
YCoyvk+wW76/SfPcifzZU4LMYkeRviO08T/PZCW8G7q+MeVxNWijyhVmTZW9D2eJ
sg+JNfYb7TeqnPo2wSVgm7rAcREPhSaL5fOb3y0UC87Yg/ztYUTLE3vVuFN6+wml
kPy/c+MNl7RmjG6hzOYTbQxYnHb7C6h5uADU9umR7R1dd3+2Af3ksU2O8V71fGYp
HTXwBb/CLeeTHJrRRbsTVbCbHe2AeVeNI+JGcJ4cWmxLho0mIGfTLqz8G0GKOL9Z
8p1HB1l4Q8dHIsWE1zFPzAKhab5pOBp+jN0DkhgdgRH8eyLZPbeqLGSMw4s4SQsu
VW4sCtz9KdexcrVBw0c9Nz723PpV0ZHKFzysu7/JNciS7IrdILejusbyHJnnBoyX
gMzS4L+TmkgT4DgogiVA5PelBc61q230QADBguLfzm19B9x5KFwzYqcuTDZISbGl
y9a4tJrYXN7sQN7ShvpAnCz+6UPT7A2aKIYk11IWESCwzP12toEqMAUUJxSvBbKu
nus6WW9xr173ZA2uiGHGixOuQGmjtgIe9vcsHoek8CjO2/fSGYFp8J/B5nOcVeQz
+LZ/fZ/tQE7ooZHJllHDoXSVZU5ppf3uQ8fHrMlrEsE7gHMEN92GMb3ahdOUD7RI
IPq5UHgr/cTChlQ3L3dPFDyKE0tJtkvtR7kb6JX7VNMV62+A5B3pfbobGKRs4i+L
EA73lconYEhcluHcyKftNMM2LoKWBZhYCiS1TGEwGjqTYKPKd43aBeWt1iku4d1C
/r7G7EEOhXEO7UJV+AY05Dw2q/QoPdNl93+oMVK55ftJwsUeA7tlPPZ6QG1HHl1J
inr/B+gc0zfoaz/b7E954gJXa72DewvwK45n9sN8VDet4s881e01KF7gkXkSqNR9
W5QgqlH1NXGRsY868wwvgFNIjvG3L+eUst3lKPMoreKog/jFczlCJKFH/QktIJJJ
/qfmih0cN557nOEX8nXPQULDzfV0gk+dK9O2S7GtK1sLRBBoWGpU0Z7V8/JP6tmg
QRDm+HcZhn6p1I8807Leb2Q5OaqsAyI4Kd+1eG6jGE9saeDLjX3L3gSnkir8qRt4
aV9FNnjoSknx0D8kfAUvHdn2fPuzwf99NBHW6BrWUZ1mPP4h40pCnZapQ3uIXA47
uxVeIoO5IAfEbXVUgS8ptcARU/6JUG8YZ7neMHtN1b8hIsLilo0CryEeJa/sI3s/
gB9x/CmV6HQyVl2Bw7a8nVSsjQTJFRVztrE9elFZays0OJh7mvu06sYXzo14YdgI
1vlBBJ6RPjVUlD/hFi8ETk+YUaAVm9YeVDb0Al7D1jrHfqgu5tEGDZH8ITsk3jQv
uKJ1Z8k9wSOxYSBvm2TA2mpfmgik2Z24nkvipBZal7uJC/rkyY+hUrWKFFaFCKax
eHB6JIp2M5Yvfwo4T9sudDiJjNW+Z1hds2z28Ve9sPcxWHT0QSF9qOF1xgC/siyE
6VznJ/19WUYoLirEqFnH9aZT249aMVD6//tM7yW/glPHi+HUyp0XuTHJNWIHf632
vl0T3T1qplK3+v5o23Reb15cN455OYwVzaASbkd8P034yAUFB9IftEKz7UdiP2Gi
lHqIIc4dMZ+Iy9iEmq8fojwwDMLE8xmZFxUbpao6ttqHRRYQjwdojMv20jR9H4wW
KOoDPhvAoEHHgou6C/MWF4vkujdpVem/R03vuytFh+6Oj9KbAXhThckx/VjirzpA
dMOWD2NhAMYDRin32bYOCBLvtZsjxgYhKuABlVyvqSFLyuNMlGCfQBFXLIEemnde
NIgmTetFH3BdYUCmMYcLqXfUf67ZSqNUe12HOU83Vc8UbuqrDjtPPbzzoYhrIij8
2G4iODqk3TX1PNiwoF6xmP+f5gX5VhL2pW/3/0JLTMZMV4GkI1QgulaOxjB0cpZC
js52AgksVvWeNuB9T/Le2xf67iLiIhMoTiw6xT8MbHO1zaruoBtJgUmsLi9EkI9J
jutIB3AVaUvz6Up+nonNqVoCta/2L2vXK85Dpu7jqzZGuLve7FVSzxy3N8kgDwpg
0gegceu3/rGh/lWKDEi4sU8j2AEii9w1yBLWmokqhLSCsBlQgsYligQbqvpB8PRv
zOOmhwk0EReK5sGCfAPEgMSFwakz/AKK56o9OsJsAkxluA+O3uk4JgutEi/roazo
7yYAD71xXpHTY0CNq9ZDomBVnBxZ/acZSx9Cj5aeIK+dATb20k+NVuOWZoGVz6Of
9ijxwtzG6ghdR/oT4zw+JOJY91IYY5LcDofa/Mz0NTs+gl6NgOkBupjUJypnHLNw
olF0jJeea/tXoe/OHpC/vCg22VWHiudd1oVfJ/V9bU+4TUVzMlz8/WizVp5+Y1Zo
fOMAozKv+77WIFeQiTlGy0B0p2RJ6MqGWRmdE+FfM2TGWwGhsOAg9oBb4uPtFChw
QGvAU1CAJPRO6BfUfSytuy6R6FDTbcA50+P7NjNtZAccmTOZ88K+BykKDDfzvIj8
AakD5RvPC/hGzrTe+/Htl0SnnsErQMfVTbBAPeMLvExC4tEDKEL3TvURLYL8oOHI
CKMtu+G3yDT93dKj5kfnhBTIfOCegRUgzA/Xrt7Y3dTj9oUE3oAPx1iksxPivPV/
oWS9Z4pmbnh+2P7OB+t5o/8tMCj6ItpmjQd0nHOD6tba4tMVLQK1rvRcpOtPTLQH
Pcsf9c9iNXoX8MjW/KHwGXg5WWLNoJa4kX0M3k33lHqpiRwecVQ4+S57SBqEAOo4
yOnNuXUTSGxsFcCDIC890nY2GrrEE8pC31yTCQ3A6qE+w3D6SncrYSTDv+k0hLtI
hkf9SrMUWXA4/xtaPzjGxxnvCPOHbfk226umKUyQJCH91Kpx5jw0W+o4y9AbVvs7
Y+GuACzlGNYs8MOjrrReNPIl0PA807ZpjcHVakr2N1iodrhQrz9sUXR2bSOiwL0k
Vl8SGB+7dcMjyx74cn3fUw/+63OLaQ5JnzdvKjKkkLeU64/cFwB8WGMh7INFRN8F
1SeJDVo+C556VY3vWZenXt6ypPh4MPoeLODr+lKCuH3NJ/5cZWqtIez+qXpvbJ64
9dNvHmNmR8+FCleaCkTEsHQWW7fWfe0nxPuO6N/0vSjrjIGBWRycs+caFWElWLr9
sATZ30nSMxqLF5gAJYReQcwmdpaZ+4vzDhAZ/zXmI92rn9J+BReHROVh48ynqJZB
wb9O2LHUzpiK0e+tgDwStiwvyAddJOEssDD1EjK1NqdRhBrwQh5kJ8A9SIndsClu
7FsxhBC+Mvj70FVexNZSCNJaTV+Lo2trqV6oIUlWvFbdCRBK1H4FdqCz2L6tUp88
4+4aehyxb8BTbpkKuzLQ4M0YBDnFNaj4p2xbeRbCd+h+Y6IJI5IarAkvVslZ5UN8
TXmCYHh+nrcJErjUIllPxFw0sUv1TZ/vyQzJrTYoiR2l1iLi2vqGWi01sG9hpKXk
+S9XxHieGDUkknLj0KECJHuh6tw09MqucT/rTD2nSXJbZvT6fo/0p/8v7+LRA6NO
phuprazto3yo17awk9OSplIkSCfB821TFemiB+JGGSAq2PQKRLYAeK0nVybCufvO
TTfLSNF0NDnm0DZkzF3k05vDtGUcIReiN26wV8t7Euq3ngTBx+tw7f9Y/KYcv3ox
J7NcnwKxpwEU5T8unxgI8vu+c/GBhokCr2ycJJXFCqFf94Fwy2wH7g0g1ACkzdC9
n+/7hs4tGQ1Cah02GYRqVr9gCNgw4CBMuSRP8x6oOVkNtT3vFGVIAyOeV8WnOJ5y
iEanCtiA+PrsbtCqZMwZGpmwWSv1k1ndvienh3Bzf8pGUXlU64YtwWM20zD+vkLA
ZerqwPCmDBC+qjpKwx3WAeOeVUi361N4ZPQRJ4no8RvctwLws5Yy7WpfzLtGmFoW
2OKoPdql9Z/0Np5yhXjrJZCTUh4TLusMeF+2V0XBLfX6sP5dMq+pg4LgbGRduvJj
NScXWRQ6duLKGOi6OSleiy4Ezxdb/dWCUgtgwtlhs2DG/zJJFE+HW6mYjZBEhvOS
cS9hWwm1YGtRvZYpBb33W+NeB2INj6xhltxnZNfEicNyVJHuehvHnTsO2TkZ7JwR
mj6D+m2QGiEMLpi7XIqtLs152cYkGCtNIHwYTraU1lBIa9iAhpHtShD0+yiV0DOl
e7kPrFnwIVAjFsbHc/oQ0oXauwmp279pX2JwGv0syAjgs7vLCUnp7UZj3X2Cei+7
MWFzg9J6Y/2YL1m1G7DHkye5pFGWSinsRJOQwii8iNrvo1h/Mim+7Z8c4y3YnX+4
JRR7EA9Zx7HaCemT6kyQINK3F+ve8BlRPyt8YNoWDfWQ4CFViHaQkFJm8KDkYaUi
4FTaY5QoUVWXvsww3KtighqRP9oOLWW65ZwWnNKMgsjiSDz3wzcetsbvwTP+dlvE
xqNBXlq024EB+dsHuNMazqqOjak+SWSWBKCKzMTPuXNqmpqchsEWpdG8YMwkM6Sy
FJAWTc3drSJZ64xGJwBNl184TaMRUaH364GnPzHxhhQ/HcU0DGcO31Vd4yOUBNVm
poQBLxakebwMdHdVglO6lvHzCgaA38g6dBdgGg+Ew6aF4HhYdRSMFOEJn/Yz+9/O
TtA7HuSbJ2g5UoNzUvtZ7oxJNPf3nCsJa65cISJJc43y6ANc5ACK/ET1iJILUcZu
4L2dE5GP8pJedE5ubu28liHjNW21pjasLIMBDEHOPv8iVBZ2HPGejAh33GU2AI5j
x4Vep7vXX7Dk8X4OsUEyPf3bD1vBSO6jPipkL38FFdmjlcznqp2UmyjygIaqekje
iFgM3OiSY/xm5dXHE9KOjP4KaqgomwYAfe0Do38g3V9Og5Zl3S7MZJEXoiOI7WJq
KApmiemynvakbSdfARwCDKNkC62LYRkiGlHGirwfsbtHa9wWtIShJcoEkzjUA5qw
GGbvYZlzBuJ+4dof7AmYKXQVFBhe+ZAAHaqJMxCuUXKt4om2qtyb/r8U4O0uB2dN
AIYIlRf2NOpbDPWZ6NyC3kQk+sgwmpBvWlOGquRt/XHxx/wzDV1NuC3EN+31P+6n
zYYQ1Sj5aBlaYT5brFe52q9SUG1A844rKQs6ulCGY/PkCPuD3Ds0sMqHcp6rLU9n
rW+hxDKlLvDb7yvo5T1rWWy5jDoXHwHmT/W69tD8/GImqcsZpnnyBD4kBLJapgoW
2k6fm/pBfkE3Ocbo6QkKLMwB1pYoOL+jdM7wDloBX9d4EBh9eeHEV0YGuiVKtaHC
IbE2TSqV6mBVDQj77PPeij5OWcvZr42i2CPoNYupH1kme2jUAeaU0Wb5gOZ1aCu+
NIVCzZYD/fCOfhRN0SEfZEUjNBXYp16fbeQfmxGHfbdOOrrlrZxXzanYbtMR76P0
WUPe0iKrdhJ6KUV8q45JuK9RO7ez5kQXcI53KvUXjdPaQTrhy41dAC0lT5JrqcWp
wHDlFjdvl+El++dXZT9oUGLIgrG6IY0lT5gN5BEWuJwyotqTNvbQa++n+ro2I6VK
I/xlNT5E1/f7u1C1OUuorH+2NWS9QY4Iem0Drdkbr97fXKv9w6t/HahzaWMtCqGQ
Xc3QhsKoRiaPPwyV4Ob/V829EfciQ36+DOMyQH+yIWEDzL3xCzOny0hsjVsbFnGv
88YMFOvQYdGH3RrI2vKm5jvz0zh2I33qXhD66Vpp0Rx1JGOwikJw57GIZFeJf71a
uQpVit0tG/BBloYLnB7PjfsS+nyfM1C3PmqP83Y39DPxgoxPS5LeqzWwlUtq6uQX
c6frT4LXImAddLeA3Gp6V0IwP8Ry16GTUkJPws11GYEmJy85OC+evXO2fvqpx2j7
Fb+nZO/jHVy5OigOxhHx+0YSiIKHATSIjALM7m/ydRZqAufG71HHpRNIqsLDDsqp
e8f30ID5pz3mqW0Dlz9rQBXRlgSmbOe0DfECgFh7nUpFw7H4s878MgOK13FoaFwd
4WofgNz/gYI3jSED23PMsNg9GUOPvymbJScnWfxc136KBNEKMoLkrvv6NUF6APi7
H7ultWtS4tbxEKDGWwcg5z00JCyxKTAph+3OiCq2HbIlhGx8R6jrWZQayicnbQFa
k6Vg2A9LSPM+ooS+9Fnq7uzbKH5USIFq/uOWQETBdrHIXiZgmLf7EyLhU5AytyCh
PYYcTEkvoTE25wj4VV8hX2Gm0LMW6/UHxqgZ9uFeYMAYYSLbOxpuPNhek69CRKpj
ph9vRYJ0Q/8SHP61FGX9ul7eHRIRK/VuyeYOsf70WC7PFIKUqxxrpD7WPzSsrad4
fZUeMvkHr3jqkzXn2/m/pRp0r9iJtU7mB+d9fccTAd/3SugHYSdb0Yua0YIqoFek
kwOQnFM53292D2Ce0f8+nb2a794fnR6xzOwhIZ34oAXFCSbwWIv8CEFsyX76Gy2w
Qc7Mu+TByh7o7ccFlJbXdEmjxqWe7CdhX7YJ7LnHHbPY+K58ys4UwjeZPLw0qXMs
7UIYCg2ZBEq4mjHv85kYtqFmcfH9eO7KKikpcwheVkABr8Q6aUIOgCThyzJU3O6H
MOm1CTay+cn5aTR0e5uIo1AnKVU22kopDwYpiwgUZZmgZX58mWdUi28txid8Vhxb
rBb6+Sy03J8HAS1KWLirJ+R4WVvJ6JQlduJa3CUTqHPH6nZ77WNkCpLRJ9gg5iA4
IG6v/YX+Jows8LJ2pxV/f9ht7DgnDfzkjmfwe4RcFwNb/YQDA/eGcRHdub/yskBd
sVAeWuBk9Fbkv0BDmSa73613UiUAOoGRNsdRzUaFeTPLF1aL1/isOu/Xa2FWKT7R
w4AM5rE8pNXCC//ZKRNdMgPxX0zdPxMo7B80bTPlTH2LXkJ/owa+YlrMrQx0e5Ok
/uGcg02N2VU9qkGnABZWcgB/wp9lgb8Uo7XP2nh2Si+7AbctUhFjX/g2o+FXjL6B
tELkIBEFAN5FCECEuMUcuJrAuWcCCNB1tf11LcRqQhUzhJOqzjYLt9ymuVQAi6ZD
8wOJEnGplNpB1O3eg8ckGT7S0GPln5OUbB9rUeXSSJlQOpBzqxmN1Nte/6o6rBh0
Bwy3CUVXOPCqFa0Z3sjwcm+GYa6qlB4/BQLZn80CB8+nEV2YVy1ww80bn7f3yv5Z
ZUiMGHE7NjWeTJW/h2UEnYLQDassn/9mjKbXCxrVuM3v1OMEd9yhx42c3AKUga3U
pqQ63mxKs4RCcvoa7scq6t4gaZzf7l+PdlGR3XD/6L6PDrW8Eo8IldvBUxukUBpI
IT1tOKpLZlBOQFQWVWMX+ERqbWjMb96w45SUNr8OxkNnhIe8h1FVDP2hOUDe424t
EeAywUp87VEMXVdyrgjS157IlpQXmYYrqCEizI26WZsBRYFnegQF2XHAQUn8K23T
boB7phozL5JAHeJNyN9MUT5x69Fn42Fl9gc4+/N1+RUdOFqP4P6yiQAjtZNVEksy
fxtVksanSxjTfumckrLlvO95NeZvsP1xZnn6xKGTzyKvlRtyBPGPG38n78GyThE5
9KcV+LuDNIPKfx0G6OJ4N5xYzZqYZrG5KGs+CPJ4B182mJ6GcuCpU9+Jopf+i83X
YjDWB43HrUXbsCZb6SOAMlj3JH5yI1xRkbD0f3RiW8KaslSkswYK7vOPQJMh/2EL
U8uOuGUq0Q/dkWYgqHJeRDn4WgY41m62xDb3YgwNY8WjbywbLlkY0371FSmnLnFj
A74HFZHunXUFYdgHzkAIUAVosd+PFbIzqvRoqYcrKP0dOMY1KujnNghHsvlO5Tzi
aXPp/PsApIOb10r3ZF5A4jyMRWG4aCbrx5kQgS+9k2nZuBKfbMRIuSpt5cDUhGUD
b2q1/otq/gEphvy6U7Fzy+amn9xAOikhk6mVNXnz/f2g0cbR0RHcMwJTrGbvF29u
nkQsC4vFm3coXifdPhFihbY7R+q4SBLM/d/iGMfnh2D4sujXZcp4lbia/YBa3Ykp
6KhJ3ONX8ZL8bCbv+bMwA7IQ53gzjWJ+bGHot4E3aX3UwV8hjd724OSR4gK/gP+k
5TRECARi0IdvZ0+df9lcqpHs8azmjDPQ+MKAwLagNMjZkJGl68qFWfxoUatwGXSb
v/B+gxbl4BbV+te6enPzEwIMRwGUUpW7r21gDBuvbgf2L2DPER05bDLIoHRxkq4G
UmzQj4vtfGqRYScQ4QKvQA8doItcC/pE57qkLvMan0/gr4bMOt+vZAQl6s9l2itE
teO8WrLTj+jKibZx2JCAHR40AJZYYvLM0bsC35YmlbD6fVCGTWy4zhyySuT1EAJW
rkY4GrSxHQVU7WuWCXhkir/N4a1groDf0S1osIsyRvB8zra7r5wqbc6foRflXz2f
uTGLjYstsmVCb80kWylukyI/dZuAa+HaORnftYK3hes3zT032tLS6GS2Eh4fXHsc
mpghvv0GMEiymx0e0i5+3uUKJvPkn34flijgMOpK775Cp0d2zTqTsC9o7QdKCQNG
bpHKETx052ixk9SoPudFj1VeZOMN9P1HNFi+5FYlSfNa7g//jEPwPIyGRtgiuEzq
IF2bYSOCZvNhics/adKfFNYsor2oXA2hxa7gz32ErQWMG8gW80o0KNe7EkDP04ZZ
+RgNCWSuuRMoYc0hLGp9Gy4hYhB4i2KV5EMaw4jh0CF7payfnIiLGDQUP6nTwgXB
D6SJ08Ajt7y3Xb6JXb61hPLoWYrKfBV5AoqF4tIl/v87uIGJgd03iQmsCBRIpy2e
7/1YA3YCKaMQXIZt1gUlGInV/v6CP6/wWUil2JZBEja0Cc8mmvA3jgROrSvB3L+R
ndEaGqVweIBiTGMfIZYYEaZqCmXvfK07XbOghJCWQPual8qdqy45OHNfCxoZHhuy
vZbEoG2RXRyx3mhwRUTudBtChafDlYlDC4QclMSnWiZEWUp4fyruJqAjiYs1kbSG
WLyvcxtBL1tKbg47gFWZ9Ah555bNBRfv8pOMY2ER1VmdvdEnUyAfQYCu2BHe9vdu
tBU5rZebv3VpuQh08uFXO48rKe/tH1ky5KJ5B0bNUUddRJW8n0xhCp87JPU+wg+p
qMKoeSb+xz8wTj03t3omnxkFT0j0//sQVJPluJsDLJW91W1VEYZjha7b3J0TP1AI
AMLVMwNksZab6vGKDtjzH8ECf80Q/JsPvZrsSqCLOHIN+vR3dLVPYWrOtWjYFVTq
d7ruZhkyzaWjvlsLKRcwPemCQ6uLghHp/Gcn2jQ5cuSCzLkoPWnZoGCV2U0j/k7f
b1HiiPPxwi7J+wNCMOlNBqK/bBRl0iL3EXtspIgv84wq5D62q4ucV9JpakwcEtxX
VUVaewXc1lkiHB7kBnxbaWR8hNhXdROylt55iglzQcJYwuLUhXJyWb+xkV9Be4yQ
hOdyu0LiiPDTEj8qRypCYlMJ0Dp1Z9w0pwl4LEu/gp1xAHRATYeerlKlemBfGUyP
dR7JLWN8fNEFLRCppKmuAaG4isrhF4FBMPiSo3yC+rJXG83OHmnzBD7m56fHLSn8
aTeq6Xi5gxwrOyiDeA0heKlXeV8vqBOY13GepzATC6HRAGB8rEsjxGleJ+XURV86
zzX5OIBkzNNaUI0mLc1gVEEF59hasFsMU6bJOAksdfnCMqhi1Y2/GNsWRwInvhzQ
MEEdmvKbMz9c+TbLKdWx/dDGVW7xtPjJ2wUw59UruuX6MJ8c85CuNZWKcF70RQbR
dO8m3kF1KA6Wh9pi28fBubcTnGz07u7i4S3vPhvEXLH3wcgacPnrPQbczSZ7/y8A
zhslxfEY4WWh3I+f1Z3GEDJLBkt6U8jtFvg66JM/PLGDHLVidBJjeAK7rkUZAKKU
FMcRfNSCMT4HjfyV+UJxI3ondOjye+WpBnq3VlEDEZLs19ZDCs0SBLqLr1mF6jtd
JID4m2y24hMeurRvsV0q+/MKmW4uXuhEMrB+5OaCaSjb70N9cgb7Y6TA9s/oq8L8
Jm1cVKA4bVRtLBenIL8NFC9KOuN7W2P9TUIkzlWj98dp4h22HfWNx42cIzyPzWCh
irMkIb8hVgzv0j8GT6E1OJrOGAO1j2jGk2qXJndqv8XRFnh7bjSgVyFsS3Kgg4Sr
uOIhS9Xr3WkyKEtWdBS1/A39UjFFS4KhjznDs/3WgJ57EXhSmOA9FvKMv7SvPVB6
5ublUtXyd89THNwOkSwE5mzOXnj3PEqOz1oY+7LoFqRYLdNzw2ECcUo4OzL0jijX
mCYIgLpmO/Fy4YQmKLsMmMCt1BmOo9IcDYSbPJajWc1wVU+cvD1DoJkGP085gpWl
zW6V4jv0vN7Npoo8EsZxWYCxgEKHBjcI0L3StrCO2z4Rktpefx+S7Nayq7vE1G95
OhybkPn70VmGegxtmir3Wik0epS35p5tW8wtGHHjsttgJwfcJNvEII/4Kt04TW0X
8Baqgn3sprmYNA3zRkb2HGmr+5p0aw0VS76Z765RIDNSijzd4YJYfte5zW7Zap53
Qk959GeBffEVUaSJ4iNkATQz71rEc2Evv4Omk7fGXBr15ya4nsK195UcTNlxxZt4
ksrQdTKm+jFaREcGArVtzB4jG6WgeT9Tc5k+LvehlRjroU/v0qVjTsS+bnwWkzUQ
tnJgoHuWkj6c6jqgrhZxOmFjwUoQ8RblLykD/OdbJmeJ0pYE4DzjpkZySGgspVo6
e67W/8TRZJHXeXO/DqgtuCob2GWenyz6PzLcPeyS/RPYVN0Ejd80QO1Y7f4SBTsP
GE59t8zlB8mv0IPbFOWBc8kI+a7e1HEUlrBdfOhWRfs2CiNvRI6gurXpPplRZp9J
PSXV+5HLLQVxh5xgcvecgWg13fclFBLX9YhPyQOnRw2GSlmAVTN7YzUHi38+PZf8
f/MvBF9kngrzPv7de3tMvGxSTMw9f474kEd/YVbrMRf5ZBZd3LWDdA4soEoBGcX/
ST06G1yBKjEicpluqTNFJ/YWRdpP48zc49itKEQZ03co0WgiLwYKc0EBZkav3fVR
4tdYcKZWA489PL7i+w5vTxZ9SHJRUEmYdeScguV9aUxnLNs3u/ex2q3/db08S1++
D62e0LfNwfibzZQ5EsJ6eCx6t3MuwmTRoAJ4DnW9306nd3mqKi15JWmogGS34VfM
KNpyIt8tjvsOR6bwzaAkhtx7jLSHl+Fdgb9nWH36LFSgMVm11jo2J/32oUU9iS9v
uuInf89ySg8dz4Eiw4FUneGahsuOSDYZ+sHFo7VjdpheVz3s8nZ1giBEPTexX0I7
aM/+ZPdETNDxeCwfteOHbAzMcidsAnlMR5J+VIAjcQ5ty+fOXgHWNDnsC7UKP0tF
Uha0e9r+OTM8oYQNqATq8SYEshMl11wVCmIO8qE1WRwmYNjhPzD9I/D61cm4zlET
5HzSBnQEZHpmsbx20ipXtCyHdU2+DEfC0ceeQ6OuYgwc9HnjCRZg2zHeTdsQpqo1
WwWh8tuR2WMaOAN+2CKRXcrdxb915bhh6JqL2xKmndOiUWLDk3LYpKyVrkCFwrxG
d0D6PyfM8JTsxIjRv00p99tfmtLw6h87sFeHX8ISyGfiC59k+d38SRqFaia6g1wX
cGBgUFucPVnzDrLGQ9DxEvOY4UqDYRJmsLxt1boQtOBo5vVIugeDfh0Fl+GQVVza
0yk4LV1kTH6BbKHMeB3Dm5RDtNcgf+bM0dTPyXs3hq7U/4960saRDxYD3t6GwXco
Rm4ChVdQu0SR2vGLLePh1iGlZYdAQ2zxWUS11s6vZmp2KDZ6nkAZBL0uTCoZgEvI
KZnMjWGa3dBeFzyMqS29U6FNi+YMxubSX81758HHWzqC2e0XD35YQHdBr0Kbe7sZ
duOmSXobQ0Ma7ChsePc6SWk5OGqwWA5hKpYEUD9MZPj6lLefcrzMZwRPMwzjo6JO
MnOFOEA9Y3A0v96NJI5i8sjeA8UwRsI+/rOSzPMZJd5G0bzlTJG33/I6hnNpXiXK
QN2UZGKEz3PxhguxjxFrT6cYdLz2yHXnYqMPRsN8XqZxZRUkuSIiAGrSM20UzWcr
t/HI3j1d8tXhogsfycRj6khmL/Van4sd9ZUi3cXBiv62sXwUS4YXhMYC/U+A2M7x
QAlFG28oo0AN1kHATxHUtqlxkLwb6sMXUXlb5aWylTaB/jGKECwyj8sdSpYcKhFg
FZ12uXph+xaTBzyFsQ6t35ao4nxgwwHRpnI117dUwHLroXuJjL3Ip1jhQhLbBCGD
6tMeJdQacb0/e/JuSBK4nAbvx6YY6OKI6Met9UGpBM53SKa4jWpYIhm9jT7Xeeez
s6Zj5N/VvoEIpY/KeDuDGZQhw3B6nfCXOA+stQasCkBxmzDoYWpji43z9eNIAhD+
7YRNqZwAVjSsb+Wbfhi4r/E2WTodqHFEr6Jwb9PXsp1YtSuTjPOEH0ppCiAPy1c+
jcvPOnmapgUw3zkLJIig0RAiHzwXTtJ9UwK49glMt2e41m5V0QvmfR+5AIdRk2ix
jO4jRLt2e+BDwz0/3YQaB9xkw4HdJLIURXV17mlfg7+HuuIV+EF71Z3NHluYQJ0i
BwVc2cqgtzEwbnxG0CDhU/Rx9A96Tvu2ETDXmqhf0aT1GNePk9q1sdVOscXZVC4K
qY58AAXUkfBh1F+8YbkarGMvZ2Cf7IqzS+pnE22JIj0RpHEM9t8fnZcmfJ0cyVE/
g/nfgDeKUtUvFwRRD47dRR1a7hLDR6J4t4ktm0mzzhNbVo4iCfZ/s8gwX2g/223y
dYVYAChSjkQWMWyDj83ue1+x7lUGBICLbROWnKyM5wYaQoJ9Yu3GvoEEZkae3Sz/
JPP/rQ4yebyv2N5Druymn2rgj9SmhT7B0my2o+kOXDcj31PXKQ141/0TcaV+Gkyv
vD6Lj/5kRSKJBR52DD5npA0jxcPjdBMbICLqLkytmP1FBMdCvkxQB6FhHMVr9QEo
A/sVsQ2imflnAnYv0HqOvV98aIT6aa0RbAhEJZFeZYATC81wpWI8TPAH1S5IpTA4
O3HQhSBl2WWvluiB4cRYiAy5MrjW1xtEUupFU3ZmbAq6NXDn7w3CiVu1QNJXkLqs
G9k0BLl6GYItgZ3RErsuJ250C/NwZCJbWG0m/DI4xF/bkBmGx8cSBXBJ42MoCP6V
WB+6nAZ6p6i+Pb3GJx+8e2Jen+rVycFRvLxrPcbsZYskuBtjseqAkTKmizvnAgBl
QbzZokIq6KcSgMObBZmzz/+Rd11+xOZ/frztvlW61rzNDGQuzKGsp4HvjmfyFMp1
JrMImDA/DeVBuVfwjeEOakUf+jbXtcH751AJSgiztqNMl5fE2ONB6P8r73idYcM5
03BlgL+5evEAN/t1Xt2M9wTmqoQIP9bzefU4iEourHkq3foTxPLiPwaJjjNM1c9k
s3v1ZMEKL0kx6yL0LYDghKgvCknpYS9rfVApICB/61E81rUJaXab1ixYHmPVQWmd
`protect end_protected
