-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JriggO9kJT8C4yxzvwr8w99AlhY4prPulzNJLkbZ61a185TOaw67lgLm8cm3tnIem/b/GoG86hkD
OurnxynVw400BKwa/oFvpkcM3vYRAWo81Q6XG/HgU/RW7ixyjqi1xVIQLjSVK1FGc0L672VXzaYO
08VlxZHIr+VgzLAXs30HuP6zSsRS9uU3dXkm6tYxjFCIIGJFyOhzk0h65fG+x0xJEaVxE5Zo7Lng
Bu411cjeKPzbhCyZLp9LnQkX+bU/TxEfox1d7v7vSOfIzWSIjsEQbBP6C9Uz9lBwSRIg9tO5uRH3
B5w5qHkoMBJ4XlaWItwneqcQsAB55OpwpzMWyQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47984)
`protect data_block
HBITiKShqqNZTK87HNloF6v4qi8Us957HWwKN3iKRvrNlcmZcjZdDKfBmxFgHzrqaD65JAHChL47
+LySH5JyMg+m+uJ2zLDFvyHPOqxUAEvDHJgfF1aHpHct88RCKkZI/2td4O2ijNZ7RQgq3LgaevlB
oM4DdYpE4uiI2RyWLNJLD9BHihxfGK7xiVbeun1+FfHUQeybIHEw4QX4uP12jpcZEO3JMtA6mBk1
xKKs6q1W7Me8KxFQlBsgX3bpE+tchMUlTZKxL53TGdaW1RYLfuFFZ4zsLZNPPozwDaIXzjbf0Dyq
KyTWYXMFht2KunXb5C/wM6gT6XbkA1pgpkxdGXHhTsDFq2MDxROFwcVUtTsWuQsFUuLZwt9aleEG
v+ZKTiX9Rs/V3khdIGN23DQtCM8XQZqpJm3mLB77+9kUXz+CNBTux6Cdzmws/Vif0WfL5h6u3iP2
5g3rd+jDzebZp2ydb5Jxwegz4BKt03ZH9MvKqMPCX0ws569LTTicRmQV/JsPwdO5cOhnvZOm8PwR
SAJ+z4sZG7qBbiAOmEbxf5bbNeNSxIp0eDukiBU9UqjSz3P1I8CM+MVrzLAtUB8HH0QQ3KVVv6u4
WwZl7ZImKhoKg8fhP+IFZVYQKhuN48lS/Df0kNaPX0f7DVy6hCt+lsJXkrVnyjyAi5Z5r52++XOH
/umjadj1JfLybp1dVD362/ucX/WfGQm3ugewIdJDpg5FBXffWswvWmJ7q2mADFO4qj0XG1O3KsPL
9xfjk5QexBsL0RoI2jeWZVPkSfUmGRB7E2kmhGeQjL4uMQEODYz1+tY05hsLqx1PSOmLn45vgowt
FGlPidC29O/AQ2N2JwHpgr9Okkwk62+aLBCp3Gzz2fR7tJUTrZ87ObK5DqFsgZYbR5+AiDOS0Gkn
0L/iTcDVnS0M70HwItMYtVRIGRnIYb9PnJIZOangVkQOAxgV9Uk5fkZBveL2nTZ/LdN2KHdgN3zn
jTEeUnmo0j3HRt6BFC4sYJLUjm3cClqeWhr8DLjHPobwf4A8BSLAixKJH/fcb3+Y5DUqHJI7SQB0
vCWo6My0yYrZmZByD4E+YDJHFx2Etu2Lb3dLC18tI9x+II1eYw/iLl5+3nwzK3r6qu1F6CV2Mbk9
XQfuqBF4Pv7hzD+lqJ+/fSWmaa1Ar6k+ER1kfH5wj9iw8Ltd1EybtA0YkEAZw0fngpKCJ9iQDO/Q
pIDz4+ONOm/A/BHh8LvVZubfdTQS9vhpedAmDDiDsCPbwZpV5PWybk3Iqth5U871/9thIovYE3HV
uDFXXVjqxfDtSw1KL8RCeiDKgmG2myZuqBEhmM0vQC+uwbU7wP6GYVFsyVTwpdv4zrYYtiVzHq4a
9OR0GTVATAgM9Mmazly8UplC5kap7SIPyCzy2+gB+Ycas9KcsceudBqGJU22QkcJTO02m6e+zSoU
k/xJBFGPiXCPd3QavhusmvReB+/1zIbJUxRRtOSOxRxDbD4puXGZpAVY3cpJPS5lPMktmjHSLOBd
RX5x0TWCSwcDQgdq+G7Q0l648YRA9voRRQmCmT2kOdQEK2LJ5NN8b82ctTWj8Us8LiZt/gm0cKML
ZIkGUh19yAA9SFMmWBPa0C4pRy0wW8LH2N9gFZadcplkuHgwQOEZg2rZcGRT1TegSkJTrX5CbhiN
2QAzXnnA9QIC4YAI0ujKlLz/p4zIgFdT+tCNYXc9saGtQDuKLtu6x82xEuBn6YGiHBf20M/U0nRf
Zj+yo90pN5fgXalKJU+7yU2DMBaEGP+B6zfax/566H856mpZEdqLPmkgkTgIamJ36XzgwpBnNhIc
fVI/giJr8b9hdJgMishLjv1jrAiiLDaKXkllP77d6NrolK4FOOXoNL2QRg9rEQNlPf8hFU7LCI5C
Nlb+O4AoYlVbNSBfIFuKMAAqnwl8K2hzm7lQhjYN3RCs6ddyNuGVuYMK7LKu9SSONJZJngXFAxpP
4xJ1smsUjENXwDHVVCY8cctWLsyNHXWADPhxPN+Bg6UdVVS/B36l7QhzFp8ChFeKxtvnXoH7Fggf
Ayxz70U85sCMVfy82cbqcKcbgG+V4aZvLQgg3JtS1kZ/oN9USdBKjEDFDUeoHKK8qYuV77rjlCqg
cSkKdYx3Tv88sTHP1nZo0zQ5qP0M+MwSZcpX3gPxStSLfUrsSAmx4tMb9PIiXaDgShQsehuFxkx0
ZrO9Vjkx3A5AIGT2RftRgps8iudThYri4CNCAsXMJx0oXpBaOkC51VqIHQjqWVu0FMUHCZGgw+Pu
WXpinDcwLSITbH+ugffu/GdHrtZXq7LL3tnmCYA1QnEewMlNFanzJQ43usyjAOQxPHYzwUyUeyrV
N6GZ66pLhWngx0mI/qA4/v4z3Fa8Kw+MiV4dy5gNmPsez0P+UNfSgTZ3yfcD58Npa6wojUQWNYJX
Up3njkrzTFrJuJw4Xtah7z70UD93RwE7+Zq+DqlZ2hjIdl+EvIIDvKbecShLZhpWqaus/DFznjhl
BwE/oL5dXrdlR8zy+OojcG9bjLqErHs+OXFTD9zli7eNLRWB5QkC+h/b8NG6b9Tpu/TuqwiQ6mY0
73voZqlDOeOSCnnD+zq4x3mGLUyiEvw1PfmkWWV9YxvBbhOsRGATvP60oeVqgwNI0++nfNFBA44U
GqEc09J7boL17n53fGxQKI268WVfRJDM7fyPPNMYoTc+M1szbzy6ORM1d6wryqcDxbVO6PC3TW7U
okj3Oi/lf9E5jMA8tEpawO64MljilzkEgFjOZCRMx0YN6EBfiadFtwWxRC0eoDZMfSAtf6ke+UJo
syFJ32wlQRVAi63WvEFw0OUAs/CsYnsTxSe+ZsWewPDXHUWFKklrsOb+FomBtJLH+KFIre6lsijw
jCnrOVWVNov+0RfvOAIygxb0PxvsUpa8yY8jcPiKEEbR/TUuaU0xtZJ2DN2jX8YTXXy+oddZhOUI
Q6acVsnnnB6CnoWNBAEWrJmhENgZk2nRZPKcOqTlDKrfYbHWjOYR8xCoaKA0egHPIN7xRA85wVAA
OOqyjC7LOTbCvVC5Qv7w8z+7Gs6IYhntOQad5dKjz5PX9VG3ZHEwK4ESZs5Af8I9nNYGId/017Eh
zRlx3G9/bIYfFN2MTXf/2QNoFP9G168wa7C/7DxjZ1EO1OhLGmf0LBI+1FKeLtblgp8gmNNdKeh1
jguHsSP92Bp+mDbhQZxI4FEpD+B7L0dgSXlvw03iIr9AMvJsQarFKH8y3i3DmPOJlCzpJBH/A6wr
P2h7TXx4sciR+BucsWNQggJ4wxkA5Ulkc1XcPaycRSi9NiURqusE9fHuGmnzpMzgjulATIgMXbb3
H9+P7YqJQxMV/gtg6k+nFOX0JJV8HPxefQrjiexFsCMZYsOPqplCegXDPbW5eS1tY38Xw0AbUn4Q
o4WHuvPErnZsXw4gFzuu1CmdpNzOX349PPaz3CCdEO0l6Guxdm8snjcF0V/fl7D4lTmJWOkdzPv/
JD32RAHcnh5CNInvhxSe17bMMbzlLbal+L4UnGlqztDHTifvTxGO2mED/w3RtZu1WAVgzvM1/7BF
YhonYCUea5XStWEOIyLRhJRoHNhcgP8/nsqgl/zgBGJR6VgPbcdOWHpCgb+ou2hGF37pZGYFBhba
iB8Q+sdC/P1L5doG1pyaHvEekTum8T3vXp9YOcjxoeWT3RDsK9A20jKEYf/NTjNuLxb7vOVjJzOa
5f4LWwMeUIo2A/J1GEj/d8pScPfTF4GQDW1iaX1mXbQbSgPErvjNRl3mLDFR1pdCheX3XwlR5Y14
jwaZJWNUtiQZPPnEhRlu9+iAkpt8FNdT3yRDv/TJfq7nZ4BCovPMaxbMGFdjYOjZIlb0bwZH4/2X
W8cB9KZRHf3WsMX4z7aJQh0bRWardktDnh5SosipU7ofyOaUVMy19IJqXA1nGgB+V9abQvl3Axef
kXZVvzoPyjdBpGq8p8xbK76l2aOHHIgR3kuXBKJhQy/ggE62JIPa3Bk5B+6WhBc4CbE7diCWb9hh
gmp4T8gJyHrhIbmmtQeOZ2H4fR0CJdCtl0KBob8L21gRqyzuLGIAUne5dFJJENSrIX9LnPRNPqMb
VXyUAC/ndkSTySfoNnGJg+sONAS+gJIcKyQ9pH/joqP7CjFZAhAImwbwPedstcNIOOcYAqTD/Kdo
42Dt8McDU6GJMKCzeRFduDsfzg6I09vwJwQP/ty7JwRrpSg/X1mEmBUJ/6LeWWdqAPCcQJMVEsDW
zV3jf19NCQSN/0MY/J2jTYm61/2wV0WKUsh7RUfLj2pf7B8kKS5UsBQLKt3FSFRH8zUuD8NjRuLg
21TLdRk+7MdSFBKRsGl9sM22JvVBMT48gvmcEZWxLz7iUhYG0uS/CRuVEBlwLGGRuDBxOgvz2APw
3sBOeaJCu1P6qiS9TlMgKPoeRavGVrZMABigb6P3rL28zzY3batBs9kg2oRO4r4Kf4krfW51x2RU
GaCrn6QOigT3Jl6Ag6AH6ghyJMRi3gcy/Ix/MDULw0+vR7inE/Q0fYa02n+Xj2hXiMcSSn1DfUyD
W5AZBa99HItuDiVIozQmCz2bm7yz0QIbKyKeGH3vBCNHe4YgHa2TddUueAPkkib9NVGN9OQwH9ya
KMGbeI/XsOodmHwrudeztuRoonuv5vZX/vPluM1aPmwD9HpHC0Sauzo2CsoJirm++cVS6s6dKwH+
zEUiXeUoIwwlvAUd4UugLjMbnrsgMvjhL1cBsZdeEP6qZH4S10uloyyGkuKdQEYnx1fpDg1ecNyJ
czzJQ9n8OUYrNOWNmpcEPvzx18pyherbBKnj4PAWNg6nEPYFMeTGTLRyj2m/I5bSkWEjXg351Wb0
pCdGh7EspiTxUeW7OLUn+38EYMuk8aGyGo9wfawF2tCYpcNecZjd1RlGUWccmfs1A5JULZkedrKO
iVsYFPGsoGhpGL9nhe2nUxUnoGRhJLAmRBYMiTY4P6pQKmvX56bKNg1yK6x5T5W3tpkJoHm6j1GQ
NLfbWiVp350C2RqJpRm0BsCN0vekcofLtPYlhMxJ/RPJwcVP5/Hw1F7IfBUc/lRNiDU4LV6VJBYs
paBv1glFa2T3H8xNkxFfeApg2Gz+ao/RI1sjNpGwE3Po5uZqJhWDhwPhz6SzlJKwP2Pfd5zMAdVn
7gPTwVJGhIQvzv0SaF2aeC/yRl6UtYaYZYDbhyzQwrcaflRPWOtVE7xGB+MCydiOZr+f0HI2GSxT
EUgtZhNODvDOVFMaLdOHezpvN9esbx00pK+wsI8SHTYa5uJLy5ZFUWco33rWzdoyp47XS2jUBZtV
TA/nNjeiA6KRk5b7wx8+3e2KgdwoxYyjvE3Siziun7nkdZ3A0H+EiXJaFKFPzoR4SocESv0hYt/n
srZHSfFMDIwDgnGKhJESHR4Um0Va2HboEtHy14LGJfjk/JJELas40Kfv3YWYlG8shcQDfl4cl2gG
hw1CIx4WRpVer26Sre61YvZfbNmTA2wkZKFn8coU/8HSnPE5KLkIQVg92vIv7NzR+IX21NXCd5rI
79iymF2EZ3RGUmUdB/ZQo/KD+oy2d86eE5OCf8anD2q/2h6IWzeQEnqg/5FG6OswojUdKaNniAWn
0lcSbJ5HX0zpsfXt3l90VqyO60wYJNfX4UfmMPj5LUTRuBgct6Rpwq1a7xby2cG/4zeZPTYR4oFm
1X9UTo52NwcOABGeEACFLLaQUle4NDHhC+m4BPBdmnrPOYp5FYOMcblMy0uDuygiicovuGFyM0pi
MVhNpc9R9h09aJEjrlHoiuR0+rkYqDbnobfq1pd4qT2I1hQof949JVsmzUQeQipaEYz2n/aZk5lT
2XkB7vscKLCq6Fa1wya02HJZAzbGPKTJ8FYPm2bcrKRjccwSq+2Mz4twp3Ll4qz6EmavrJU+bXKc
3sX+ZWg2TYW3vGtqpd478gxKQsheMS1JszxyDGQ0zzttHmYYpavPZnkMJS/KPbrZaDmC2vV3/3t5
5/C2BAuiGikiILCbuqfLw+bGQsu5UgGCVsycOtxFTVOZ+HfkwPQiu9woXPCLsbwpcOiP8xDERZZN
dQvunv+GUjWRAwUvnP2xtA2YtX0xUP92BiSh5cd8Hbq/7jTqu7gPrgjvrQdA62CpK5g17CPDAMQa
DKluxjKNhWJLCcpRI8ZQwgCL6N2ZlTMZGbNuMNHZI95VJsuW3oTkHRymEIlsrgOUixWFzxXtwcwT
1OzV/m369AqzwPIJirseYh8C0ipLGwMipOUy+ZOBWWV6SEITDkNgDbwTmBTizEbEbCUxT6woGBWW
PJcYVbEP0l06tNV34Do9XL0m2vV0/kziV15ICYnWlD5HG2ggu5sOU874NhDcw/q7U8PDdISHOuKK
20+I8elbT2nd/YGmsiBibANL4v3WriGPs3OIIooa5yNnnTpe53SHokifCxwLW1Dbw8oo4b25GACg
SZzGSzRgmeXQDFVo29Jpx4e+Rqe+5/QkkHjMag/kswCsKYMJtDhVdoE9P0lRhx7AtB8hdMIJwULO
ibUdpTCskcD5MzTGIOETonzAHduMXmpOmVyMiQgkntexHSQmRrs3jO/dAmIh1NGHsOMb8cPknokr
Oe1Xlt+/PCMsjDJqj93Y1BHdAI8pSoc3YjhOoWXQJkoO+Rx0M/kgbIxVzKhM2xTjS6EloRCaXaNX
prDiNiRvfPdfAoZMq29YjM0BzLpq2hJAayeCEaUTHa9zIaw+NTcT6xdq/Kz28J8T0yq6SYu84TRj
u5v9KaOfOCzo1LVXr8egJ4ptSMRKs7XkwURaQxO+vcKNHcXgOLpTAVRtwd/7dqiFjB9/KjVbX89E
8KQ0H5KrXts8ph6DEc+0OrpeEsinDu479cvQvyYbveOgWoVBRJMo/SsZixw1qAZsVM0ve60yyf6h
Rrk0T531nZr8Bm2x0uWoXmLh6nD9o+izdPdLCeCHcJL61+TDuoUdH0uji3pj9e67KWcl77kq0CmM
ZywxCV3fd3FH8qTLQO9N05k1Dtww1oyhzDopm27dqR+KvIFjdPZ0V+gK3IAUUNKYwas53RPradcs
tH+6P8y2pGIdHT5zYE+snW/x6JmPy86SWHTkzqdijzPo2msSW8S7XIu7rJMdMtTr7u1evBtlqKz/
qcljQ+JfFGDAafUZaLbAa9MS3edNtQ83+RhIgmDoHG0B6YAdqXwxr8Z3eV89zP5PY+TDaR6h5CAB
WyRId8s9B8cNo8R1cQOy686jEec7O3WKCT+UmnfNdiaUF3rZ+omjgwFE2g5SapL1sfHtIlq5hzeO
4KgXoHbaIiVg5nJ4uaYZDdF/3qN97Een29ESjOjBqCpIRhpd8zs6H0ubuAP1PW1YNfaZglH7Uic4
Iqx9tbRJIRwl8TGvvLrsIA2SaU89d4gDRpUVlwq4oIB5zguOKVuzDrW2xGqNrNkhRGKluXGAgsod
Esj16wWyFrbbulgUhU4oq1vGDnc2rc6lUsQk1lUc+AsfqzAo8yPrj3XMvnmmARFuqmLKl96Fk8Xt
O2LVUqjnTdOdzW4eybgHmshaJJEBnggUWTriKk6zh/6dGtDbs9oy9QEFGBB+5/FKCTSRg1IZP7HX
uSWRQ/nlosThNSjyxszCsnx63BEmgODaqNiZyh9Un0RGdoKpRekRSxflVdzCpxzxzRd9LmMwMYKc
iX25znsjp3ire3iLLB5Q6l+6GndngEqETB5qFtyzwvC+5ArOmkdn1QTYihY9bSuvFzkDqyVr/fFm
nCkPJXe+/L2ZBn0wbUsYPUTCtAjcFIqk8WaCQ4nf5R2Ptwehta2hG9ZHmSBGMXzq5faqQ72X4szd
isbMHPFwlSnMQu+ZygEHMj7ouKETTqdtviVk2xlqqvktcXq8VHg9jXY4wfw9OOB3GMNqGPPLdBzn
gfgPPClyo6QXn118Kz9h3PY+3tJZJ1ayRky54Oa+jAm8dXtp11QpM6Ht/DMW6S/Ix8Ak09nB0yZC
QdabzfrjxhdJ+Ju1VXhaUUVAPcz+H7uFkPbuONRrrA546o3gSsAlzxDUWpOMikVGppSTCsDfoCBw
BRkV79YSQmLZJL5gX8zh3s4R96xS+HWc1HsGQI3QJKDajz+IuDgLkxaDFLpg9sNE7l+VfJGkgOi+
TFAUoCdDEDDl5GX7RNN2LzvHpVexSWOQfaY+DP863+qWu/KUCiN6uVAh+W9Y/5CgNaf06zNicyKR
ygVgpG5rdGWAmbkEi/5q6ivwW8GrD14u23iuCEmxh2hYiS4GvW5PYbNI4GfVRzK5K6ReOqDmpa91
KCcv72w4jGnw+KrDPzfxpZ0X43PK3ckFKLKpjHtBWuN8PPGMDvCPc3KAOi7HxvzS3OpbKCKLjVQm
pZeYRuObAd1Apicgr+OM/vE8MK3/686iXda44hkmWT3tf19fvp3cBwMR2Zb9CrSyqHA5Q7kexyjs
8f2bfLJAbPyLvN7ucwXGlmRKgdYhKGHUuEmL+zWrlJ3sS5Nx3XudWzFB98K9YBizjj+IcAn6/sjA
xO5MxJxb1PNPXLnhVGPmys7MeAl0XodzULSv/9jMqCcvVvQ94kAm4nsGjRJjDQV8wHMtCDkm3UEv
Bf3gCjRAKM+DlRRcqJw9ViszeC3l5Vm3Qbto/vt+Lmxx4YFf9SgV+AWuMGUfqVCJnjeYf9eUc7pU
Ug3+HUq9ZcvMdmCACbrJZD1KdEcuPfaIuwMQbmLNAJzuGO2pWyUoW9BTuVWE92oUgU/lnb99wAKg
T5LUQiqyv7LpngxJZUI5DNuU0WWmNtq3/vZv1WbAozbXCPBoWBHqEzBjHtfTe589mBz0/flNNjRK
E0LY19kv6K0Nw4paLHZvsr7H+YToj8z3NhvfuMCH16ltEIX8SpmrL1XNoEs3tsFE/5ke0jl/STIE
sLE3qUFk3L04l5bhvIZRTXMvMYjYSD/CxmPK6nvX3K8hTF4eFX36K94t3a6kgGOGNkga35J34V4j
kXVSNzAr28kDkhKbEJhNv/iLuNZlwNo4VceI+Br81QJDbBWzEa6Ymjf2MEZeIPYezpBfll3484+O
L51utTlYLH/u4SZLrcxUW3bsSgxYzQqEE5v5d8AWxh6uEVqb4Dt5WaWHp1brGfz7e3yiX3MghMhW
W1nKw/kJtHLZgN0O904Lk2Z4XwPkhkdEoS4PwyDqi4pE0063vYd67SFL87Kngy8JlpqB8PamNqnT
OLxsaQaxd9o6+6/H78HmXDI6DtiaZEt0bLmiIPs5BEc/CQNGXkFnnS6A4Y+XREjB5J48cK3N32sp
7iC0t5ff3zLbsE0uuXfZ3fv+lXMzDsJTR32Om0NhlsbnDaFEfVP8zuL2vHLvWLlwCE9FEHYAL6mb
H/8w5cb3EYINEFc2Aee/HpnvX6UEaoc8erd87ISPmTByIeVJ2djiHc4oyTu22SHA2K07K2YbFQlX
V1wo0UlLKgNmHNLHAcbOzc9wE3eVOzibV9+1YbD8o6sLBBdw3g6YX0g0Za/WgXS+mvYE+1DQ1Wiz
hi7bKPdUljFwYPzjWyX+jhZdUJfGoIiGSXuRXPAW6MAuVF7TaTrDbTWVMNj9SSoabchTm6ANUNEZ
836tkIXKcwrdoBrWMZ4EbigVjh6cxfIBo8B9bKUISoJ1+DJU0aytKE3S5HUhzTabRImRuS4CMe+x
5lUJHmXNfEftDoX1OOj1vJFt3lNua5RrzTekChtCeeXx2T78wrdcY0HcUEGOp+uL81W6gh3GM8ch
vDiQnIJdA8X2mC5dPxV/QAm97+i0EGFWIFOnjmUfROdTf6CjqAC1F17OiqG9Dq1L6e4uhi8SMpG9
1dQHKYpD2FC7WR9wqUaIOuovyISE0offd53jqFniKU9kxjeQSZYxL/KdUOEoUX2h5khtvzWI//aD
O7Em83+PI9UBtifcGp4O0Id+/5B1TtL06oPxmJPNtGaiwfKf/euAYum/Yd7FtAcJhKQnfDwRuOzL
ybOty8Z3T7RucXebmw7kvC0RCDwJFugVJfCdA7B9WuKXx+AuGNJyWXgdCv5VNmIzTl9YMhJbgf4M
l0nHeSZmAKupuVW5/2S683dwuQZSyVaTuQz+NpWk95xCmEtF6oQCFr+Jzo3JggdludMtSP10BNo3
klpYSD+ZxeCHa5OQl704OGMqHUhi6WLnvWldsakKPn0ACoJx9sXstuez+5Qxb37ldm93RlWQUfHX
uh25zbJvAcz6NWjPXHOKaieYt+zHdDznZS7fmTMRsZSQBiW5UhwZ/QTYkTY0drMksM0y54k1pb5s
RqmTHG6x2NgfayeUr3cafIo7OPNMSKQPIxN0fqTRl+ogZPhXNXeSeVzHpvRWVoBLXe41dbPzqJ9m
5xIetYSCuU6OAUWo2z0lbmCLNRcUyucPyBY0xjWO6UTnRpHDZpZJSMzI6aBpyfkIufkeQnGmeNiT
179vV5YLujG9yyiQ6yGr2ytPDTFM7ALqKf5VKJzcBaO30KDvqTNLuyrI3kwofdtEyKh+d4MOKwx8
pjyTdog5xpDxBY2lFjqbrpaE0G/IP9hEuRCBD6ZIRoTLvE0MpIMkqZktyLYhpmEiZbm92zYT/qcP
D/8tSjLsQyLdf6dGu28dLDp5JKtgv8lNQs0EwFBkrlZOwJtAkVgfeBjoybtIr/p3GhsVL7dlcikU
RVPIuHoUxmMx6JLIMmFC51iEXZ3LOCQ+v9JYNAc5belOCSwnjZ+pf6Y0WigisAfzKJe6TljcUv5C
mNpsrIeYJGDNYtBjWuABb3nT4xfChMw6F7mXCbQGiLsoLQBPsTKfZ6vt+ZmO5+qJAw4cx6pE1eOh
Q8bg8vv2iuFLy8wHlWa0KI8NZoDyyyRCP58Mbzj6iCrqyXMDjy3yRbW9O84Frfr0VN2NNSZ2xr6i
0Q9CNT+EiMwH96SRP5sLIFShyCEVLQ5mIR5lH3Et81+PirEfBtKipvxVDy2lAaF6AgF2y4z8gOFw
My1mHFy+bRKRtjHtQoIf9tLWQGZVPFIPY64GV3kwjnyq5foO6FDfrmyLQHfqL+Wb6Gf4pmE3rUoe
Oa7ADdT7hTK+gSwDB4fbh0z6LbOtXqgTGRtj1axmVcAsrarzIHtcVUAAOgJ4R4S3ozowIkN0eyWk
Y8KnEC74XCPl6lcmg26q284B/phGuby5sUOwHdngI2H2bs0XJZmqtVWQ32a6wldLJklsEt8Uszyj
LruB1Q0MAo1FwSP4aa4KuOGj57Z7+uHYmNeyhjqQ8BGg8uT3dDHpRRme7O5hE7wHTUjQfCszvr5e
qIM3LDlAE/xTzEpgLj0wcb9F3fQY8MlwCF9WBpw88ToG6gBnNY2zAeSqaq8BoCmmFCXcx/4FV+Un
NAFZAIT4RudmYlF0j4ePRDEw40YJWnQ4osUZR1VUoxxHex2z1cRaQjX4C2bEGfJ99s6LRbNtcr0p
kDzg1y/2BgbhU/Bl0+Z472seq+HymJyv4ObE2oemlRcHRDZV9O9jRMa8C52UXKkPDFLu1hLxEHIW
Rov4wE1SE/h8NCfxzDaUvqL7kkSyiIdOW4E5FFTk6ppS4sZlclG4cEzZNDWKwb+ypVt4RxcliVml
ByJaK5OKzf1bjILlkCSP/rwU3F+5WRnIuCed/3gcwbKhqMEsGpPJ+AyTqTJ3eMkGOUB2E3CSyZIT
SHoSpEnz/3jOJm6Pq/ZOWF1MyMSDlARa1rPCMvr7UGyXaTNpv+R8XlzYe5inAub5G2oaIn8Cr0UX
NRaICd7FKJ8cD7Dsz0JSmZOq7PyoQfZvt9+j4TQQCnFxXedCE3K7JXn+X0AUQiwWUwTQRFY4OFuf
ZVLvzZ0WDHwD7i38w8DduXHWFAr+psGuW9Tsn/c2J3HiMtfSUveRbO/aBkxUV2cE+K6E7rsGjSlX
KhehqyNRaCYXC5rxvAnEAkjorODpi49Voj1aVDz/1pL83+O7q5ka5tgMqIAXpRmxWVXVHBIw5qEO
eIXJ1gBYa4Z/hlXmEUbosHd//7xOCKV4CK8xVxsULH5xxb+1qVp8E5wwITrOZLo2uofTnEY0+zjC
M8xTwAK0GOzCrK3eolzxp3Uk6Depu9XarIwsp2hAsuujkeXK2aev1UpEHfSdYuCXooDYjD/s0Fqr
s4++4a37eOBeWxYCD0B7nVyZFSOnVWS+VcSAFyfYTYjczG+3c9IuhxOni/k9P6vv/+CkIxfzCNpT
/oBgPkz1ukJkbRDmSDJ91bdngY7MFAmVcjN/tGZ0qnatFhJMZcPZ7kfnfXcBOcEm6MulteNFwTx+
TQd0Avwek62sThuIK2FzWG430owXQwKSIRJL8Za1rWiAmophozoLrOPBa9HGFeR0USvx6Rn/krMh
tw+5/T1nS7yvk+8ioWZlxaqmMeW0nu95+a2uTphei7MQ+kiKOG1RU4NaKzg8jIp/VWoKXBT8YwRk
u7aHD1DvXhdXYE3767IsRjeM/rIyFullrSeh7o4fXJMatimWDjD46BlUq3EKaBj6xEzTyGowaO+5
ugC8zJtTgkle8/QdEHGDSXgcgQ2IAasfKKEqAWzZdq3RyaN6qNyvl/+vdcyNBIV5hQqG+KJ48Vfg
44iE8X5EQX/tFEhxgVE4osSg2tJ2qmR3c6Hj8bH4ZW37hKy5p8b86UuRz9z/aFIxBamHwWro+NUd
jJ5Dy15WW/zXBETVfwuC3iF5X1csr4qSWxM7g4zCaMVAtvwIj/pjz5BjPesrBg6W11xmR1R8ftyv
wv8Yz8UgSguMXIgvMT6LDX/75H4cvjI85GRw+upqLddbVDsjf0oRAuA9iRBcUO9gQ+dRKrZdPZiM
GLTe9eSQq6NFrDVxBsd2I/f5ygQg+zT3VG4esLtqa7ZmahXABu5qIGbSr4BU27IJJSzzyef+jkMK
yXAGp1vEFc7lB0/8dax7tZpISNnDdT3QpjKmvYTGYRq8D/rWzXAuUQ61ed1FovC4DGRl5A9uTUf5
mYJujMTuKbPuT0jvImeU/eKQIjLVFOMr45fkLy1GQ6cMUP2mt17uR4vpVSaDTyzjmV83UWdRfZSU
uZKgB73aQ9wHOaDDk5OBDl6DHYolP9InFSNpsqR/fwZuy08HCQUj2UqkosRxWK/bTLRUbNzJUZLm
908md7soSdUMIgsHv1gqlCEP/Kh4ECZOa0ShQsGJR3AAs/OzdS7Riqi8ywKTqJzr370KqHp4whdP
8MX6bxb2w1bVHCuJRXYSOL1eeYkYcZSOCpjIrIB2XtIuud4M50gauGmXemrc/HqElo9JuMQRjviX
dfi2rFW1XziPjvNtreU4u4MYga9lV2P8ymWb3PlBnOxNAlvslWXCQTq/+i05+B/VOlO4I85gQ41o
tQDi+vfG8AeQmuncA8YW0Qs1l3PHu28acM8EgHtAGo+IL//Cku/KIKqQkazTCAhhyabysO650SMI
gODFGw+9CXND/TEDJSMwI/ZnsudZ6WypU3EO8Nl5ZvmSx28mlP3kS1pTyY8L9kRPX+ZIagCb1Xz+
WIJiha7sfrhwwFLMYVF2QJ4PxTAKAXp69aVJgoMH4i1y5VhafWXOOsLpKvPz4swRR+AA1AqMmbJM
5zgdlVWx8II3ejmOVwEbMi4aiHQJCuNNauBCSg7RelvGdPM70JJ+1sFpHr1NOWPpG/z1RONqkScC
rYh7qntOzVAgUV0DWSoVLqqN85GXJPV2qlzNhwm4GGt3lLReSTyMSOdcoasjsu5/SkqFfsgEFAvM
C0KiV1XcNQjS0aKurkoF0dVBRWLUIzNYkNtjBpgt2JT6WH7ULyO9+orHAaW4OsURSON4Dx6F94ai
whzT/ChvftJN6ttKiXc2Lu6smRkxRvcOfO4sbjo1bobRCWB+fq085vQvxput0jS4FVdi1owIJJTG
qrSaiEljsyXGZXS4jX5zofg4IQcqIn2kC29ac7E7ybWb1hGPeCljWem/BVTGOSzf6rwPQ5NsZF/4
evBjCc2FzMlUeUi/CoaHqGP9pM/4h9xnYx17x2b4BFFSJDFrp/FiePcPDgEWPhHXee0k/0tkoWTo
CiEMn5nc5uE/Wx36yRCSrdNJJhMJYMlvmVml1qIFwW7731rcxgpiTGp9IrfW2fBslb3Ka5F+thVB
kPtZnYO8t5puutVOywnBd3oM0dO6D4IFVLocq8bqecr7DbhXE9LtT8ZtQ7CLHp6Xi/dLfm15PQOL
RtHsAtgHZoIY8ijyx+kIZZABnVQ/YMN5HG8f9jazuzilOWQOabuEKOCqN4seUvVLyO/D113GOK9M
4hC2sf/mRrZWIybcYb+W00GVxwzh7b9iMc17rTuVx39x50//1jpmTm9bMfWZVL5uE7ulQKDKosTY
6ojWk8d2eKdPBQmbiCr0qPZZOg2sem9KfapSm0unWUEOPV9oCZmARXd62hnntTUYYv9EpChs7t4u
/1k0LpiA2uM9jL9WvcmTSs7qARsGu1n81KIN8PKPFMUf8sYi891eQoIP5LhPapz5vSP0JXmRGKgF
5WO/7uor+VaucnCZrFmes20NcsZ2MWpJHABN4Uo/G+aeFfyTaFUSWfd1Tyx2fyD7hfdGBdkKJAxa
9KE6ZhL2aYQlU24L0F8l/u3DwJsqIFt80SydhohMYgGJ9OV7TQMA1+qJeVYsKkwf97cubHWHelHX
CyVYf71BsX9SYNCOT1jQf8yoq/oUriJmHS8gaGuOI2FreDQwhzDIYIhrJAfKnY2oOntAZjsLbIxd
BNAZj6jm0YmWbZDuUfHuCFYwjF6v/NY5gzmzuR6kEHQ7UCNFeD+fsWBaEj/dSFI5ONowSRjnrVol
i/FPufOAhE/TgnEd7oUKu3ii3jfHicA0qfazeQIq8AhLB0KDXwtloTersnZtvviqiC7d1M56fsJI
EWcoNTkUjXnkGAhZd21fmxtyyrAjL8XLvg8ZrSSrw963a7IUzOAFR6hBi/uFinlNT/iD9UJEFrzq
TfyPNFjDMq/n414On1rkadlFbl0VCvWZtyUY8SvuSPIW3vwiOgPV07aL2Y7huPzKa+S2fFmkVQfn
KaQjZZgMXiVEeh2sqYb+2MYZTNXjiW6uxkHZbsHndTweNXgL2h+qVZ7iLH+jdaJTTJdFXi/qVAXL
RUX6nIS55m3qOB3p93dfv7iHn7apfFkz9UoVUnFjpmzZl3f1p2/d1LJD7QlZFEkgHKKngTlgsesr
Zmlz2h01ZwB/5uBMfXoJtC9kvb2AwCjbUOJEHkVTTAyHKvphRumWlkbiVtIAeQdDXYeqD7w8Ue/e
2rYeYgulnh2P6m49YkU6ioknojpXmp0DVl4ErjgWh1mW9e6g386lN36W9mYWG7eRvv+jOkmR8W4Y
U81kVuWVjIGtyW0CjYTEv/rUcG5CSEzM0YV/kgJ/NGfbcKCnhoo7SzPBpyaQQKM2dF/iB43dUp3b
pTNXLmYkiZ5n6HWYXyT/tfFT0Rvrd99pzY4ksAj/883JGw9Mc3zHXOO2kwFd81J11CcngQb1ycGs
g+SNQKtrTJveeTNUDUkzBxYFjrLfdJ3nwKHmhCdcCt6urth7iom/6bAql6K0VembIppFuzyue8Mb
DkfnCtKtOuIdhPU2q+mtptF2YOyz/RGrZd6hlvmG6OwXq2Ib91Ds3gCCEV6uCcSAKT9q92te4fs3
rygK+4nWNhZeGMR/Gs0vYs5MMDexl5RrZiuD5ia5m05LivaPduRiSHDCiCAIZj7a037K4PkYldDr
u0Nq+JQoSy0UEqXRIm7xgTqYoe2e7nmmrQgowZ5xtqbWfWFCDtRf4qpiQtXPv8dF0RUct24CNt7b
kwZjBNFmoy3falpa5Lz2clFzoUVcZHU/Vvi5LC5cHJ+3drYvte1aBQC8O/3r07kkce9EG5FiJ50i
lBbg97ML1zuO5ecblatWViN0S6XqAH0yrpnU9NhnbpB+aVEfyPcTbFuVRI6ujFvx52Mvi+2vzWyj
E4XQmGUg0161+F5ncuhIvOsSMGgHwQLh9aBbZdY65J2eKeHlWZBpi0DDhC1LrLdDd7y5dSp9o4kc
hTHnnLXI0T1r95RLrBhY3fw551piRM+vrjl+tLuDU1h1xRiVg29m6tQsLImUzHCFzEKC6XgSKskK
35BKHpeiyeWdvm60VTFy3CzFXs8z9bBHcVRjqHuCrG7tOM2T8AmPJu2BwDWLOoM574UO+ktYRPDM
iW1ykJ0MAVThUx7q6MWG4XcjEJ9BfKudoHHhpFmW3LR1o6Kr9Bcbv5i05V+QuE1y+xwfUsJmb6NK
YM78uo2nHBiy4JDmhwhW00s8jqwxg/q+mbiR4u98+0M0YPUnrApQtvj1mGzdTcojdu+9s2zp3R56
9QCwksdZ6xqE2DTHQ6iUwMNF0qofIQ9w6NetvXU4xBvuUTVaJhwnjW4pRPpV6birokV5EaOhJHpc
B0krcY9/5gvXRBQUzLVxFAJvdxGpx7WyxLBgmVwyWtuMG0AQsetCgPzBOHRQHFdKi70vfkt6Xaw4
PLrjDN/z01qpL8jkTDVj5jqLWGztsEgzAK9kIUhmYBcEhEQzVHswHxw4zpsq+jfv4FxeraqwUKSb
pYRKawPfR5FtPo8ijlzTPvrmVwdDOoVrTa8j5qQUwGmVxZg9tS9Ry8vKIreE7mEggF2uavB1v7D0
fbVLdChxni+XdjnMF+U6SdQs5BKEATgFQhmrTCpg88In1822d1pUpUhQj67lArPlCZ4x+FcWPKPT
9WgH4ritgeDI4jf65JdJaN4PWd7It6X5lyDkl5AYqWoFMGAbhO7tdZ/kgNXHsz2C+SXXN8NJJ5A7
n4oAX6XAQHBylaS7SStwKau6NrkozZ43wBNy384JBcYzccqsGKhyfQGf1N4jRRgWX2CEescyIhRv
cYEAgFZGk2uSxiVhtcGEO28bvs+lvLhdDMT68XMR0H4BcaoZZsFqKSF6AUkGERc5NQ4UlxMAvHV6
tWkz1K4MTiuP2r2dSDE4tYyJGfia7JBwGPWm1a8JWZI/TvBS6w+g22qGh441MxT9TVHp/ngEjeS1
Qq0ynXSGNO8eoemX3PJWzF0aFCIBTiPLmarCEzGAEg3nx7asYHZx4mYtRhQlUXCFvgXY/p6rsBAt
53Mg2TIB7HcihuvSPN8adF+HFWBPoBFg7pP2xIc5iq+O440+uKaABbf/mTX9116YC/rsnjSjlzOB
y+eYsEOEvypuf/vIajy5Ow11qopq+V4L/JvD0d0fgxusRhHNZt/JmtFtCEyV2UEvQhvoNve+VWB0
SXYWNFgr4IshT3DEg77yHm04Tj3pbWc+guzCgcwzqWvGONX3tL6GvqnQ5jDQ4JDpZtQxAlX/Xdgk
rhYBvfdc/kJbm4LOaVlVfgVqaw3x9Jhx5y54LcDhDNLruLnYMJYTXFF1l4p52CrzMWLyt7w/QpI0
vuVmaQQTTrE+LUT9t+wZr2KzgnR3/pg0GjYFxavEg2QibgrHvKAOSI4xlIXT1ffZVrw7s3WI8tMY
Yhkku6s+5Jvbmp/dxTKgkUAgIdAZqQ8Ym6Azw+i4dTMMhqcqJ3hQzpFydfrhiSferGoEFYecjfEj
s5U3ZHUL8ZkmC2vIBJyHtkkJL+RXSEFyEcod+ila1g7rdxGdVI+qVtG5h9OifnuA/AZ7czAofmt/
IzaxNmHoyBXm0FZq/HZ21aHDtU+A26TBnC7LKx4SNizHiZqCKCnYbMkTmvjVcaT4YVABAQLEtF9G
tCUUH3hmkRfDbWl8Nkr3b2JQ7EH8oUYAbufiKWj+WyCDKtvOKBtYJeNszrkoMH6wMUAg73xI8Q7M
6HiTiheWuu4Gis6SI1IywpxW6F9a4EuYf5Vf2vXOZLmtqMmvE+0VMx8n1MtNURwFV4NqkLjnD3rF
RrRGpu6OL7THc3pyZDLfi/Nxzqf20xkZweFQSM+5Q27IWnwfmMB74mOpQQvArYBkI4tMhK9iHiir
oXrs5Nu+f/S3CHOiL/W8Vmj7Tpq6JHkUHG0G2xfUGzBgDC2hP1r/+SEg8PTBkWyX6ri8SaS3O11f
tCS6FAjGqkpyLlv685b6SecQttxNicVo3UrQ6zfWdky6Bth8KVCMguYHIYAxWoIwlzB+7GUs0gwq
Wvyt4YI8R/b+SEeGF0I0SwShz3OQwMQu0iFdVHBUO6cnoE1FKARbOAqQ4XAtriOvef6mrpf108Cg
kxA9td2fSsms/dq4M5a2u/up0Al20L9NFNsctkqYpEcuH5nf3nqii1N2WJ5hPyyXembkvD5g8gVa
e/j4oBPbjIOhmMxp1xc9f/EBPNlWvGKQLdVSOCfwNFMLjpIwFEi1u2tx2vBeMRZ01WuVxHXQNeKy
2QsTRJh7W7oDUztMbfZcnDnkKQQcdQH6tcozzkjIqlkSqcm/xTX7kxrc2ABucfFlwX36JjCLN0yg
+DRU4lq3rMfrY5OZje//gYDoRyNLXlTm+oWIjSRMdQj/AfGtuWx5G/ANdMhJGXOZWpat1z++B7WH
UV9HlCnl3VKjN0s4B2DUT3iAJn3/9q9wKUP4Wp13VO6SAzv7fPcf4Hby5YppfuVyMo0WQVK3MAku
n1OgnjsgnHbEJte6EIMjwaKgKq7uOPIe5j+fi5C3HQBiECsCbuwybOW08i7Fyv04VS6FN1liv7KQ
nUY4YpZI1o9xn7FalfTGUFBq62T2ZgZM6zX1QG9qEgTYqZw3kwJLQNr/N4Ur6+Wp0nJDjfdCMY3S
uqJ3CWAt1H2Io+frxBNkRYWjPHT/mg/xiha6JYRZZcdHXnr1ZhLdXNXHKVvU4FdszzNI0hBApcs1
Kpumt7wYxSLYWvnsPIe6sZ7PNNVLLV+XyssmBG1HFvIdgHwCGdc/c6IKbtnHjaj5UVjDd1VUpmK4
8HmP0Jy/lhFeXsPrgijp+lvH/PSmmUCB+GN+1v8RQYDHv2URnTosJbLYEh36P5IADwmMe+3TsXxE
uDN/y8Sm4zz98bHoWNPRX4GlOQc3rX6MXD4OExePEYS9vGWo3TKP5D149v5T0OKxJ50z1vqY+ajq
yO0nxrb1qJlxUQWi7gxne7hoBuyzd2cNf/XDoAHvrGnOrioTdX5ECn2H3aTIBpvok5ja4ab25P8v
4HOi/dm1hbrAw2VOHYquf8YQLQS28U4XKC8MsdjqVjPv2qX9LPukFYP98tygJkmykha3f4Z+XslK
nzReb6sUOwWqlq/3v+JLFChRWxmwUCQ2moOBjLYYuKpgmn5vKRwLfXQBGRdyLOUODymLvS/Vap9S
mhYrQblZyiTO/8PoFs39xsbvO5OTC+H5hSiYKKnq6pbYH2daYtru7OcFJNo0lJlCwOsiWJ0erggu
u0nKyB5aWHHerdIF1gjXq/9HjNEdG0KXIkx6wTxav71F8N+tYijCjndFvci8u5oae+TsYGaiQejR
843UH3h6HaRIgeD7TtdeaHlgJgYPaEIlb0NO58qEalZFwiKuiZNCHOC6FaawZg8rvVa1ABYEwGfW
Vt7WC7dPqnLOsYg3NUJJywORaEbwZyJHM/TYhZPlSW57vy7cQCIZxz59ddjvFc9Is5cMN0ZxvSwq
ihAjaFcNCuJgizHxuEn7biY9qfyeE+X/ZuQu6g+jfg9bASudoDmiyDzHqcO3/6oUDIEfntatxEZ0
/aDQa+t94IqLAu/0Rrpy6e8acI0sxzK00pbnrB/3Kvu1wVFOl5eC/VG+5Yw/dhS4jdSxvNa8DQJP
gpNEE/O0cw2+UsE0WVgBL9dwpcrdVA1oyFBgqEEMkiPk9H5Lt1Z8dY+N8Ar3lMGDa9gAHVk37O7g
5+LdOBImdN+7SomqjnlbrBF7AVH+rcUniylNrtNrbj3yUQjumFMNPBiA07nWdQyL5eatFHqHsX5w
xvnhuwIzXYZGcBZnEI6W34bipHxwow2DvEEzIcB6459dYs2dONyuoNg8hBPah98NFantqlj1mcI5
eIJ0mXplb1hQVA3DHT0lM7vu7XLAV9O5uAIfa1hjr4eM4XmfYC5srOO9T1QyY72GBN4/X5nUlHtW
+/FZzmaUMoxhOzDekrL8nYQb1vKY04b7b2JB/y2SgmJOu1ub+qt6Da0Cpg48MSJ/iOdg4+3Dpuyf
cyh8+SYvgJCM51nwn+jXImPlefXOLR9C5bp3WOMc6+EHltj9/K8SXxLTeUu2nVIOyvNWldocMIu6
r2zjydrdWcEWnIgFymX+NYjtHoihhoz+qXGG8yj4M7f2LdrB0nGlVkYvAdXyVD1/nNC0JTXIx1XP
2bxcrKaTKSnCCrCTeDH69Iwd/ugfyljnRaMZdtoV1DmqRGYrVGk2JP6YkzKy5Nux2CubKvseW6s/
zizgl8pccIjCPn/uAu2sK4JeNuPK9ewjI4BUIe+QBS9JTBdRabAkPEfOsuOnYnR3BOstSd+GDTq6
JS4RwsgB1LePkd2Pq2atHc7XqfvtvX0TiTZ0IgtWDE783P3zKyRbXEyUtU19FW76RX5/3hmDVOUA
eoogTCjvhoJAK8uHlKyl+IVuKSMnb3OYwXv7rNmOq/JTxzYPkYmVyGRdLK9x6AgCE19PDJEp392v
W35mfCVmtvwaitgMXhqc2Pb/Hsv3FGYY8oSsgCEGms43jF2rALS4h6ZB5WO4iSaYwe/sX5ZeSjjE
JQRJuXq4xzaMNHKhIjnFeeIsjmaoQRUMhtUcx2sI7fR2Vb8nedUqXHlOPFEbRQ6APVff1iJKD5Ev
0IEPeBcl4jAc8bvvCKKmUU9RCCQYgOtqRLeeAW5HLR/dwMxZaj76bOZJ6QPFUlEPU1jiN+XDXDwy
gEnmmtJ3gcCvK8U7OVff03hyOs0lwqd4Do533UxFUvgjpQQmrN2VVbf5uZbF6smHFLNnq6t+T4lH
c2/1x8zbZ9GcbUmf3IfhtpQD0KT4zBypxG4biTWg3t8a/JEhdIaPGeOW4VUkoaIvO5vHbKzSByqs
2BF0LOUggWcJN3H6tJKyO0h0dU1SOfCisNX4oKElNkydFoNpgiETyV4ZJRrnyRFRydfOAko2rx/r
Tlcof28VmUfsWFa6Ea/Zhf+yd4LUgV8sPf0N3LIveXhmfJrafH9ICD3fL6t3jAIz3nzgzwdVKngV
rVE2ESbu8p5pIbreRjs2wSpsx1jxfT3TGDuTCwq1SvhzQfA2HfImLYdiSqHeMiMqv2LH8cV3SR3M
5CMStEi4FRLHsjRqlo92f2VKdkI4D9C7rqa1EM84RaeYCtG9Y7PlG4Z3K5vWapxP2ARHU8rOo6NS
K+nEK2+1XaMcKcxHBiLWBdowqiSjBTrJ+6eoCUGrmwcYRQ0D8oF1nGhgYkel64cunoOqUnNdYKIy
3NBH3/qAlkF2O7oBJpG27JGjZ8VczB3g+vcCgA6OSK17KW2S+BYDZghDXBVewtz5B4xhQbsr4wj2
goxOnaw3SwAA39L1kdVVnee9xodDGpk0/dif3Rz0JlXLcmjiXe515pJOFFnbEXcjUQQWAsPpJCyc
P2x46eeOsqjp71u1MYOor51mD7BTULuyO2j2J9qdxwVM8fv9K9U8oKXe94WYD3GdPjZYi/kHIkcq
OlFFgoJgtl0XNMA+tHs110LEorwTPEt+pz2um8xMeBiRSRPOMBAdMK8rz0gEY1IjlYtnXvNz4Pgv
QhFMX1CWDtRh5BGduu3cLBGvm6Hw4EZe0DLU0oHMYDCnDis2fPUFjUb6EwQs3m+wSsHx6r/W17Pu
Yrg3iGtJmf++8jp9uzivSiK/EF+eY5L/ig77XkmDV47OqXbVcvo/zvMegG//bUpozTAXTrmUD/HR
bCHy190+m/XBFTZlf50X5qSYITODe57yXKVlNPC/uBDpSgfRUMx3HzT/DF7UxHqr8fUX8oV7U0pu
2C3C36xeRIxNSw27TXLJuw/f+zxsfoWIcFlX5GV7TRH8qhDpRMv0eARY2qG5BZnRiDMsSJGaWib/
2Xqf/KRDLTyGqZd3klJEwYqWIwPPxBO/XXtRQfgRwIpsPNSmtOEZhWwsUSEcfUDiIdyJMY2h8PGU
v0rwW3c3llzl+uhMn/fAHD1Hsd50Mk9KMbgQpenrqBb5mODrqmINMjYnyNOO+Qdd4Q1f9CvoNnQ1
ABkR5bCAVyvvEH7/TukO3ARgz0ZiED7yw/kmSPQU3mracM1JjoopqeTa1rPNtueajOk7E+BAJoO9
Lke25urLIGJVrb1YOirInPr1ONiBi8PH6VZ1SqviQX02wN/hbD7nwayvl7KXklCSTnMghS5JhaF+
ZEtOcGPy87YD8SL12FYEI/qyWq6/0cXo1yeKuUMnPVM133Mp0AQXFpWH+9FvGTjEbKb0O8QI/RFf
VQw3F9orO0v4RCPA9dxyUDB2l6yanEkMT1U4budoRmmEd8GrYo25P1YP8ELuyO1hQLSiqaj4Eik4
iu9NBz3y5tJVQ15vzlQeQ6zQhKkMlIHlPIzYQfYgZr3/OrHt/TjlMREDB46UtBH2e6xxjfGARR5m
gxNhni/N1AXSeIoNspgOa9TduUzKFmDAqEtHUvP8RR4bPsn6zNkL37YcrNF0vBZ2wzLxaMYeJGl9
Bxp+Mvpdy7ymM+17rrD0iX+qnVuuq4yWPNuDm9mfN01bByWghxUrFMyWdheAQ9Sf45vQFc9X4ZDz
GdVP25wLNr2L0DwZEKRMISzAiLgo/1SRKu/oZHKstmZT6gGW1RKBkdyiktYrfgqKZCQwQvKo4bbv
K0DrDjaYCx/x6K4zydr91nOwqPJk4mPFUl/Pxa7ehCxUryrO/hPQXy0CfiW7uz+w3P1CiHQ7l5iS
Eo6oLxA1YLBuSzafqWrjOjk0WKsB0heznefP1i6PYXfS3PuSsfDgmtAQXfC7IG0JRBS1FEuFHapN
BA+8m2U3VzeS4/Mzu5L6hr80MD+j9nLkX8L6eJYPCIliNEJ9+LDDfenN9fIutMTyz5sbm6l7xtWo
f+kvq2BPXl4Nxi4BEEou0DRE6MZBSFvhKqfbK+lBN8SVrq7PfLyMtu+c5eNwRcBdFpDO/LY6EgqO
ZzDBoOKlDadsKSrE76zox5vdrpd6obs7efXp1phVYcc3nZ/yLkecG4TiINGV4lfNd4IYnKouPhFv
yvgZI84KZRt4d765nz5NRpsoHTVjOQa1264YOv7TuZu3PFPzVRQPXMXXpT8nf4Zr+U2qif1iLSK7
RhqTmo6USgC/Kgp6ElAEQ/anM8JDDGcyEh4AbXiIfj6ZuiBymdsLdK+s+bNyIwNpgbL1T01WKWUX
NP+q3Vffg5UlHFiDoHe0flMnpCS+J4sFDLgJFTQHYrKe2B69B9WM18XAYS/bMhEDPB1lRQ/LyBU/
56a98ltMrhj0but9xJ5l3TYkBEx9gAIwdmP2i89gP46/9U21ivMd/F4RPZiu5wexW1l74jxEheJC
lk+KTmVof2ZqZ9g95Dar0afxQFrYMDqg19XWhWPtZ2Sz7lH19baZhmmSF/KGZG+7Nz5DockQh64n
XUI8tO+CCG2GcBctF6rH2m+mE0GKiDNd1BroPaLsrxgw7Lmt1bu9jXgnXJmtTfIFP9jWpEPvDcwv
8gwZv6s3jZhkkwBCfz540qdrG9hmdFP5k1bmSlQ0nAVeMIuEgtEqDDSO6SXMrOqw52E4N+zGzSSU
sv63hPPZO3RK+NK9pywlgQKa69GUgxJ2d+9sVuI1fPY61OfoIW1CnetIOYYekeDIWtyWH2RKu9ie
3wLbMknrVZ87vHoxAcdDF8wAEEMfmloocaBqwvxY6TMnKuS3uW9S76fu7L8Bgf57LuJU4z408ke1
aVmMl2yUCgeN9vkwEFYE8RT4Ff0EAjxTd3QyFkWhsu/g5NZthQ1n7l9S/OjW12A4ud8mfn1Tc/gd
OISx0JYfeI2KyJ3pi96vaRHhd988uug8MfDuCAz+59bDyx1Kw8IwucqmcCjUoqHeIrgXNonEYsdb
TTz/LQGhPpBUA1o8dIP38cX7RpKVfc+zNyt+AfIrLLFPyK/AlyAKw7yp7LawuQJF7NzRE3v3J1RA
jIUwPnJqCkNqkuu18uxe/NNuIQGSVkp51zcKfmD7nh+w6oiq9FlXbM9qe1UjzeDSJkL/IiKf89Kk
js4Y9vIxD2LgJN6WNEdpryxhbRwVP0lIYz10PMtPX7RysqwCwNWJVXWwgGUUkpLh1zec4yQENmO1
DVXleLIU+j4T9BRbH9DvUzu0LTSiZNyylbtDZzHjCirHGQ0mWIf7hWKNKocODV/8bN5Hpd2AM3FI
Hd1heUyWwn0QpgYZpdz/DQCJmmwkFT2R+hpbHWD2GgaOq5e8SsM8IWJ5WmIEovdCr6qa9c8/m56w
MzUsChPbTS3YBemsBEsIIe82RE+1md6Z/ImkxI2vC/EBhRcdA6BmzJrajgTRcgn0l+BD7uqP1Ju9
zrs1i/VBjzU+3SK4O/yygVAFx/SQAt0tNzcnPBMTb5i2HHlobfDXi4hmYHkifTiYLrr2WA9niCUR
+7GnDYSf1GxWNL3fCWRZbL/Eja6Uza6Bx9pt1qhQ+dB7B1BFz9eqMdaFZmSgrYDedCsWV01mjrwy
K+tQtyMiU7lMrwaJKR1uGS+MSuk65IOnerUEu71GROgoJVxaGIVQ4MejglekFiAqAkln4GqJyPrM
I+3RKfxXduqYIhV2nisFuVkPU+BJTuj69n8HcHieE6/pJiKcY06cimuYEa2j4OwnSKZ/PV+Ghwk1
tPgDg4e/D90lBp4ZePvPl3TMSrEH+kSV+RIXoCROiQ7tmLujuyjSM6heyqOrOMicZHCzB1Sln79f
SKDBmdpxiQtVpsh2C1qsVjsmJco31pV4ePonDhOEQ8LXNQDzu/VFElLhu+nxkMiNMSBva1Frpr1U
WNl6a0b9SH+ry3jIT+Tkhr5il6LBAUxg10XUkNWVJ4guxKdHSdRW4E277v8W0ATAZKe2HLFmo+SG
uoOERhHEDWRwQ3aihJbR/U0ZMbOMSYWeMKVJ2Bs3e7p5QLfh8ANX4ynfuCyNPm1iryufDFkRxhnq
ktSRRN2itEKMqFi0xHja+nh2Vppnou6OdgZlq7SEQ1M3/TeEKX8jgNRc4CEii7sB/OjEY8jSzOq/
zjxFE9DCpuEl1tI1ByOd1wQHYgK1EL6Xw1ujvBW3SRkJUBtfU/UwtV4j6a5xpg6oRDLB8jxOuZ/P
2+aNSBSp7UzBSmM+jMn+HbgjRjRBmnhYIzkOYRAMOo57tcRpWhj79H0SEPWmJ7aY/ok+fsj8y2cz
fYU02wSzw1yHsXNeMtEsA9/TmgIfPzEwxqTfhCAXpQYZtsrM5EuoR9lknh7yW+2W98ElBPqodF1x
b/72mvrVT3sAdxwqlNhIHAY/lORJhRD7FvtV1KasG+2LHHsRVtQaf4wpTy/kSvYGCDeokjt6HS5K
sLXlz9CRtfDtWQR2WmgJ/s5yJNcsCGfwCPbMInFy+S6IlEvVh1bhgERA+kkqw0F7iGnZ4dOaj893
NP5Cd/DtICJPbPf0J4BEI9gjFHCt500wwPxyJlbhrhymyXVAacwACh5xJNbroznr9AUMDSMfSanG
p8hj+upSoFUJ3QG2mw5v0d64OP33r693uolpwPGEY+pEC3CUtKvEFtUc0EGK03r9Qw4N+1ynPEBJ
VGPcYWF3BHYE2dSjPWVy6PrzEjLB00Ik6O8mAiiLHWcXP5gPvewYOK2w6Vp40Lfwsqy5S2GAL5gh
f8zjFHbYHCR3fapP8snhz58mz/LI//4eUvwe3HT4aCAkK7eFsbPaRL8QwY8lLGRTQXvU6cl7GNkk
CWIyYU1po/wL56DCMIlKaKy4hkrzuZKLUg4dFR0F6BHztR08RSqaaSmDwcfBJiuvlEo6kbz9+uD9
+8RyT9n5ZEVjsOxhm5HN6Tn8D/WSyia22uaS4UrKwr/M+l07Votc7uQOxnh7Pxa/OP/iklAjawhE
nZzViBJw9z4/PXZXxwwyZEMLWxBlnE0pqinMSn4O7TxdK9UtstraMpbubcvO6jiRxMp41ZtVh9Kp
d7z3MlLsgoW41lJ6SdROqMnjoDrAREXHfP/qsWQ98afH58JuOyZ6zlxtCS2HcgyxPl/qJ35pX2ur
3UxkQpEfUf9txp0PEaR+1NTPw9LOtx+IhQdNqSj/L8684yhhPfw4hxDr9sbvfx+zD4UsxmdMBikV
MBjJNcbndC/PC43lfP48wwQIGMknkmHL2CyNpmFdKXkdx5bHvDNMOelakU8v9ZyD8a7i/f+I7ewG
scC2J1d9UXF63KvjqQ5X5WTJJFZP9yEw+FtMnb/9UfbVjnvN4sSF0v0JHp6AkUogKJzp38nEU7Xv
jt5t0Swf5t+IVkwZb7Z89wl7CEtJT/sdgPxOkYt3dZAXeR0oTGh6VPTa4WM7eAdBELYcyWFJmg09
xSFILmrHKELsWIqbLInW65L7sNwtpoyzJG1JpdDZFALDFRcAzIhJnnrnSzczBLKyfHF8XsEwjWYd
Xxf8Lt+MFkh5bzu0zUePN7+eItI+eY3O+yC3DpM8xr2mp+UAXU1jGDWGBVsqFkfaB1u39KMDFgTb
qZPplVOmvaXxvJdZFPfsoRpQB1gQkeITwgzgZfp2tDf/QILelUbU25+Zx1wkEAy5QRMBolZldl0J
Xm7sjdjBM+BuFoEJ3IdMDzgMUBz3gs4cbi/UnKoM38+0lqU/nw9o1GMZDReYjnT4auFWVwlQD0RH
ECrJI+WVg1iCzCmmF2IPYsJ0qDdkkeAahGNsyar3lFpqU/IoLNOdpnaD62Bwkarz8DZC8tbPQV7i
+h0AJcKCrFzQQJ9oBVOL80uwt6VIf8L/2tlcuWVl+HgQAFJrFiNYqq9rmsut/YMiR0PLOiQ6+02p
4nIq+CmgpHSdXxjvoNw0pXfKTriAKdwJaDyizIj/gXY56aOk2p1NMeMH1SKh9yxmKMP80Q1a8e1K
TVEnv0dEurnM3amulppfcbAYSEMXqJPk8QACL03UAIUQqEW/l3jMYtVGZ22NSXzMhNpz8MH1OqS9
kebbpgSaIqaRjg+G7leRrIjxPimhb0itrS6PEZOai5UImqGgDlz+UonbcGK+6FRZBPCBUEsE/pLL
iYQKdlQkTiV7ShnYbZYRrRvFd2zfwGz4VAqPwHFqroTaCBTtvkxKGDxoamO+Qt2TOvZ/qwGKuz3Y
Hp7VJ1qiD5AXfqDVvbqM9cSUVqeWwOiGDbxkHK5SLdpSG70TQdDtnR0iKIYmF07anjUvYltlsw7x
xpCCy6q8xntH9KEoO0z9+6ADcSlSW0OEFq4JZQc+kLNPWeapFt2xsKeTqW8cjy8GnGOImbJt9acC
2OsBdCdP/hmIyEGjvic91094/5FDC+2YAjA0aY4DEEFXf3FtIkmzDxuXwHwVhxcV+s4t7iMpJWUr
pvuIQ+jHYBGidxp9OX1uTOPqEUVWXiuFrh48tWcMHETDSOBe+cgVZoPV9lWB5hrkPO7emCI1bLz1
xdt9DDrMksIoQs1EOXjwc3qSMD6jwcrylQgxLJrBqcN8HO6rkRiry45d1u2hD6G+iFQrgd3OLboE
iPPTOz1vQ012NKBiQm+D97b6TGAtY3w1cWzRFB6eoXG79JY3Oq/GdwQokSFwwvoIfVHW7VsNiWCN
jqqxk86pQD9Ow8cHBff+oeH8uixJQzjBBzeMjDM5UJc3J/yVVCcg5XHAIgbR0fMsVK8mCh0st4Cy
dwnMmzaVv9xZ9AFoFL7eI9phniPix4xZKbRZcIWqDBY2ojDfL1vdx+ifuBpZU5+dwUvR5MgXoAjA
jUJlBebVaz6CZyeWb+Im/i5P3j/SXymuwzGd3nX/y1mJHakQdGfHdnfzdT+nXMNFYddImTdBcWOY
d+l8HyovTRXIhufdaMThnPey0Bss9LZ+KMLPzUtRif2OWDhvLsNHX6EmxVUNwj/P7CvjeryYnOqy
74mOf7/mKHU0eWW0d/jI0T7VZoJf2WwLijRDSvhru/mLb/V9LLqakopGHsClmIu65REuB/QZFDPc
otK0WXyKHh5E71Eci3dWBFJ7knCfbDMkP2cD2fvOX7PtRr7DuIBzrGcVhXhMSx7d7AiV8FQ6eN/f
c4t6BnN5VR9+q30M/2sRc13DpMEnoMLJTeo5Z7KfFseXR1xO0zx5Graz0pOEDLx7Jg2OzJBPcV4M
GuAXGmaWDFGDQy2MxbcVmgLKFck2tPf6V6C/mTwRiDxBa4Rc+bt3/cRm8L5t8uUk0YncHgXf0O8a
IlMvpMzsw2DAtuk/33suRsR+bQnBfaDI+NOrIvWLzIDWI1JZCFUeOvXjIMuHVHg6tY6XxL7gmj9S
Qt4rbeHWbGMrDiHOIYhlHHndGLGE5PSa7mBTRsqFTOWNEvdV0fBwxyTQxYMiiJp0h9ChAilZ1pdw
neghVs7EIkOWBWlyozSskw4GlYQ6YrLv42aXh8xDEZvf//6VmEBZJqyn6q7CzKWByEwxii50mRia
3wVXweCo5rkfEiXClVGhuc1tFZuHTDsB03tlXHYRKd9rOl927PDSxjuhflvRa/ypLRzpaWQIzWOG
QO8Um+1la56dqCqdWIRmwXFDvaxFOB5E0i1RQaOc/qW4JqbyPD6Suu2cp5UTvNQ7chOt5iFqcpnT
2Eqkn3c0t6B1PoUm1QjrQzUwRFtEjKrBR4Kc8DcXjdhTuFFBmQoywu3KQqRAoAVX9govXH3Xg/DD
+iBMnKGKlA//wwR7HpbwrNwbDJ2c91J4yeA7fr4GhthWGjzK3WNuu4St2B+T/7b2as6QBWHcdb2e
ReCWpNXp30vdsU54EZomnsSf4jINhrAy5sTWBla3avOpZPOlDrYmDSvt5FfeKrwqL9WL2drZ37CR
VAi/Zo6CZwUau5vqgS0P2s5/y0zI60pzfv4Litt2RsP9827TIyIdwqCY+N9tjgj4US9Zd3hG2qZE
55xAUlM6em08Z2KbMd9TYSbQsXnGlySBLQ90oPr7aZU+a/sJbL4ZqEaaobGk+nOv6gYWoi4kXDEl
GWjaO4G22zpElWrhEWEXZjOP0m3nkdgzxF0IHGTOzXo8FxHYI6QRZkmKtHhhepOu68sRkFEQz3KA
00iuarlr6NirJFj4k84EkwYp6stRMX29ajlAwLDTFOPqlKOQlqFzd0DdrggVPxrLbTHzSRBlZULp
bJyN92AJCXInYlvV8GMA8jmklIi5cbeET51wfncRL3wq3OqE/NhtfzjaYMs1bEPuT0NAwR3K4Eru
vP68cA2YyjdoswGwTzcyNqkYlrCrSYU+Pw0QdUK1o4ct7N4QsvpDkeDdSmZQPNJd/ysNdlN+hZQu
DoxkfXZ7ELjDfdMJU8dDeNSkTxZyX/QHWwytGYT8wDiN0F7ExOJVUvptRK0Vk1a/Jd1FgiuLe67o
s0ryzRkFOoubymIlLnaIzKUGy/B7AK8r1fO5pgJv8aZNjWWLppOOymR3JnHzLs7jYF7zqgC0VQG+
cLosO/zcWnKF+AOVn4ek6MIZNkuikBT9jNrI8yS9qv7hSVicUfeW44J947oY8wZrT5wpMDRvxt0G
NWDWRkg7bfEu39xooPU5cguVnO3u1PuJibOUKMTh7W8QNz7buUlrRfHxcig9JwgVjOoZ20ngRIGZ
VzuO8DXp+Cx2ofGZKAb55l8idH+ZTveMmawWpH8MpWWQ2wgsAyTfqmEW6eQsVSfogP6Dnag8CY47
+2QcV56GDrF8ptfGEt/xeneQNhommfFPE4/KMBkk7JjWhgdPaxpguEWaYZKOEg+OUb7LU6oKBoA7
bVLyLrCBsmyzE8VuKv21d+FT/URVfB8MpqatkCJPyVryNJQS0APYcrXZn+RaBLaNvurLw12+vZgg
Rh8tLwyrjrEbWvtEoLTe6OWCgXu7gq/Sd6cMTabog1DzIQHCHQy/r6uACS3rMr80zWDFylKgN8mg
gVboZIyIQeIEly6ulYC2+7UfsUOrsKvXFHLyb74qxD7MnzMvGelO8KnPckxaY9TRHP7xAT1ezmyd
AeJh/p+GoGVjYEtD7mj6EzO4cJ8tCtfNX3g0GBU1YuqgOVw2rkKtfAnXUO0p613OOqaAqxnq88gG
fz1hpfnASLs6uSdwUmmZgUYeHfz8vSyJgH+tqekHvVMgC6f3Jd3QQdrRpEv8KxbSmJdRIEQQkMyv
o3tf4y9C/N/yV+7gn0XHvdSzFVCs0wEY53w5WkJzQKXmdq5udeL00hdY4IBMMmcN25si59vGdJrj
Uf1ZCJTCw8wF4dvLeICJZ86Ucr826NTZmN1KUm1/26oZi7tmFzaYwDsrQeyCRouFGI0w9REOFcdb
aXGOrzC3ffqu+iAsPFUscx3eJPWjsabKLdaJGrfu1JhLiWzEzi++aFWBPvZQioYVLjypiBA1SiSF
zg2av8Xi+gAg/fBvEs7lLyLW6de9Pw+9olwRvKSU6oIbtb4w4N6fOvXnSMoxysriwwBwwJmEFr2i
xdzMdEVH1v6bNn4FCs6JyiT0SxcGWo3TXwfSFLsEA458g6dfSBD1lObEKK6korGPYhfhz734yXpi
wrdCs5UmMHdGPEJwrvNYVXbJKs6Hzm13x7j8JPjSUQJh3MyrfrqjrBH8KFFlGk1Cc9Iocp7Vttm5
gAcsKwBc4uXAYTtjJofuatK2Kzd/3+nJwpALgQVr/KOWvvn5kOjLDfI4mRPSW8H1+aPThfGpE/4m
bdspM728f/18msPYcAfcLBOlwffaFT//2IdpiozcX28eXj8kGkoOywb6LhD0pWHwvk2MTgMTueP3
wPzcyFD0fKF9J/uaFMU5p0WKxaXSoA0q2KSu5IzdPEnws4dOQ30G9j9LmxfOkjJONDVcqjCaQd5o
AND18gusnDp3HXRgvpisKSFOKIpLB3gtKn+bSdi85c8og18kXXPB6iPAw77qEM/yjfRRzkJS6b3+
Bp/FsRActLWDQXDsBJwiKlBO7vOUVt/+EQTpVMz/dNhto/KDD1NZk1Lqe8rRJCYN3THjbKtUYeb3
JaGGueP7TVHhqKqzVivzKsQFFc+kc0WrXZpPInCjhZGmMx0l87IMQvo23Ryak57u7hQxsNJUKar3
UltoRYnhZCPld9UCE3ywz6GCgYoJJxNJ6PHOjEqI0QKchVSZ26vY+905mdMSuWYZPbQaDpbhgbXf
c2bt8zkMwBZSoJmq6t30vLEShMmTDTk5nsEeoY+Ihr1KCoQ0ltba3Q07zOQ/UI5PvpdupayZFJyg
GBT7DrbVUoqdZ28MP1ujDdLJwEozcg+twlApHzQpSOYkz8Kn1sKPasEinj32KLBX8+iHl0gCmlVt
FrnIkwQVZyx1e9TEXUAxPZZkKoIjMxCJA5PIiKAmh8vlbKoMZKPZABb+Z47fI3/Yms+dM2aUtq7D
mF2pGQc9GSSUCBJfZ1vyKEZ8m2X8T+Usv6eIgYWYK+CSgsAQCcwZp7lFc7K/GiW+FG8fJKvNDSKQ
vsmyRD1sdGV9blHUyCTyTt6BXxwWkOzQ0WRsMlmakLxn5LGCIklAMEDm7gdTNFQHncaXhFq4ys4a
3WZr0Vh5hsNTjVvDxGLLu93NppwV6tICFiSnCQ5oV3oPRjZJSJHpcucs2YgF1cfD/ibL0R/7tuYc
6BMdmVJGyayNmHis2Sa3U7HKB5/jtNJODNCG6m/AUZgMDHohm5Bf9zJaLAyZdLqQTy3hVh3iGunx
hcUcG0Ea7ILt1HNyT/5NkXtu7bZurkWAIIAS/R+gm9NyRyuKvAC5ZcfOD8V0K5npTb005CYDPBiZ
fpYTmRbSJifLByLfXB1utFxhfgYzKYzRtxH9LSkXDv2gUZVLT7TDi8VMkgOz7WTWVSxICMDZ45Mg
4/uTlXQ6FBzuJrGf9t7Z4OHFOqxDYV93NaOmLgBUhG4lE5KNu9VtqS1CgSOFMEzCu3JWQiin5eay
KNlSYkfg1Nb7utSL3F/+K2vb7C8TK3aw7VyFNVYDDKVnTTEqnNcnoJ3U74bKkHf5h6X+PRngPx5b
CHfyEXGuTgo5rFXg3n5l8kC6a78LwhKC3QeibQdwN2bOUSATa7AlHD8sAaa2uC9Wvf+88kYqYZ8L
4vneVhArcFHRCfq9Bj8SOgew47FiP/dijt7atrIDwH3qWqCy5vGcbnnIncW8n3p5gbEe2LqtgAsn
J8JTce+WgrQwQao2deAYhyZpmpW1O3eWGgk5kqlI2yQ21CwjjpGI6KMlJ74xqoO5mvHxzF37GF5Z
6K81daT60bcFC2r28W/4rzjv01qs/CY2qpB77KXrCnkJ09vTsMZmql8XZHIaDnzsX2DfvtBde9iK
FxmOYiDB7Lt5LyQIXCyRbbLq7/5TPM3aLd1XjiIxfLv9Q1LFSaXCUlaHAIm54InTeSxnipO1flW8
8twXRNPIefU7NSxCXnxygOno8ng3BqNZD4TsgU8KTfPYHKCHjA9yUsyo0HqTeWRxwdrZcDJHei7Y
PtZSEhV9H477QjHmGTdRVZ4c3kNDfJijF1c7yzH0cH5xPlaM3xqHFzss92JmCY+Mq26vFKDhlR0k
9RQAZpoLxLAInoEa/QSvHUjMko3m7OZcuXZihblcfw2EJh6oi0/baMAZnwgHknoit5l42y00OhaC
/0WhB5c0goRr/Fju6jOrXxeo5gOIgylq4zaOnPkCfH5pGFZ2GeiRHbUpqXwIZSYdiF0B/vKPojfF
aC5P0m4vBGhag253nSU+fSCUNe2oVW38TCVorU80DuNvXH9Lt6+2Je+3bLs9pSk7uoGwZ2ekgktt
ZJhKKNDsKPJBdyDRNADJA49GRc3lt5WPPrHl+araKCzu2zLP03QFzFu+lvhOEpNGVFVxv75nOTzh
mqJX/4vKMUbPaMAB6FoNO91JssytN5bdGP9jmLk4yqS8KpnTUPFNJaI4d1/hb73WtZcUsAvBciOG
Jy27p097LWxtqwNmJdn0IdCTPV1mL+fToKoEv0pqYGBAT3hLefeWq7d5YEvhyM7Nt77SXwbAYv3w
yc79UVQypv2kwX1Fs0cJoeC+gyWdQtaoBJFhbTQfhrp3YFoA6YnD7hwcI5jYwBzDMPo029anZdXB
5Mx6NhRLbDc+em//JAbxkS1Fyiu4rRD5GjYRb1x/c0B3ga1kfotJu9zOWmsW8zJfZc9MZn5CCAAl
txVCvGqc+WUrGjW/XgDa4jq83r6AbgL89ZDICjpCGGsQbBIW+NGXREezOpx4Zl8yj5ChDI2mntKJ
DORWJf1BNGIflSp/rDS9xz8jnkucrChmlDyyuBDEsqumNBTrpXVvxoZ6aj6fBMwH6dj5435V/YS6
11JX6nTCc3lXe2cY+PvVOmBUpcldxIj4J8A3+srnVVGyhe9OZACjhYoLxDIV3J0eEh6A+O7u+v18
zIaVxpbRCQ9hBib8Q98D8IZgCcMxt+QYPdUMj127H+uSykhJ96VtqPkP+ZVefPfqI6Jv/jgADHYa
/ekB+q4kOem7f5G1vzbW5k7AnU2ZbNEgUCHym4WWCpiI/43M34TgG84AHsJ8KChlQHeTexIIJcMA
aL+BZoSUqP82171UzHwpbhUUqwgmmsafKgKDMrFRzDxg8EK9VzgODkqkZndEFx0mD+9OFamtfMCg
ggj5AH27WPY8P6qVwAjoowN07puKEbL7jk2roVGW/fL5uSmnUcQdYDZHgmIhxbOkLYE4YU6VQnhl
gSq5Sb+sUJ5IoGXif0dhbFFygh1r5Z9ZfukFxkGHPxYGyBYrttbHNEMiUrBU7HHcS+Jv3t6fvKm4
0ugfDJrEFP8Ww6TUR3BdRWTG6v5OD5cf2lOPDbi6zENSJO/VquNfG7YJrzhTRg2YMLhwM2ah58j+
KaxmhQTvBF9GcHaecmngwN9G7dab1UF4IV8q6co5eQDYNBHg468UOz58Nzwl5h8Dg/7EVVvO8JrT
9L3xr/yb4Cvy+jJOwJOkENPsZaqecBaFzbOJInCauhOtzXB7QZOdeZWommpMF0PmE432xwemaXtU
E8DMfPeE5D0s076V1l4IgQRjBub3sYjqFSHQVrsRj91ciDuYZ0uOwIMUYspx2mTyE967r4J/1Fhi
icbySJjDBNCtirSn7dOcctUtm47jLLN82SmEWmqR3HsAkERJSpSoXO0rWcFrupaKqXbcz4Lq9V1X
cZO1NNtKxhSpIsyFjB9NFW/hWG+DZcjGF72Nce1E02LNoNoNzgEXbXH3U5NBnUiwrDt+BP8+YTiY
ASxBxImYpI1p2exWng1qDPq4BcV8OFmZF+Hf5Xp3nkeIR8k/qrX+jO+61tGw5O+8pfvA3ynP3Thp
qW9ZrpljzFCJbXaXclhwy3BZ3UTbxCneNOqR4z4Ys8pF1UhBfUD8+9N/r84eENBLQstTgJFSOUnq
nnvZ6NQdBvk3kKMLqsjT1RYM6dxHRhbYS+4E8P2IwMYqDVV5czqhDJvl6SulMW3vCWR0A97wk3sX
CEadPMbnPWtqvj7FQSzDALa0cj4VBqTiJ7Zkzn0otUx5zrf/G0r+IffZ2DZpApzjPiri5XSaS+FR
vVl6MGTkhAwmPlL2nLkBuwHlsmKoxv4dRxvjPgEIeLBzLRy2KiKW+6yPu+qp5uKsHu/FxE0/VAtN
rv1uUjC5PoWH1wHUIhkdE/tS0lwk3LhLOf/dQaxTXRH4y/Jh8DJSElyWPbqw1AW4mtASGkLwpcpg
Az/pvaZ/TWVX4B8aycASvZMEIXx3Ko5lYQbpok/dJRtGlHyFGtHOgJGZ5bm/1i3riuz+wGemXlSm
QxhVBPSahb3r7AxIA07/x+eTOCqiRjK42Al7FLtPoHTm4WGk5mBxRdKnOSAMb8wo5MUu/bNJfWFt
RjsAl3i0faI29ifN1vZRFDY1FE5AIaf2/6nAkoGlONWYe3dISyxJ0MXH94zJvnkgVUxtrZPZQeqU
tfoqcaeBvsMSppLutuEf6D6vn7/lA6Ony5thv4faFBmUL49USsXeU+gvBr30jrPjE7oTaALMMNZ0
j8GBOME0KtCJFvwAUecWYa8A3XG291FvxfX+N9z70ULnVJEHlj3exaN9i/I/g1fh+wVvxl8ijeND
95vXgswNj/pgt5iJ8J+sQjxN+RTq3vPDdQcGzPDYKJxVG0PQh10OyQ06Kya5ww4YaCdxIUiQs1Di
ZN34GlpdObIystsp8w+WCxGZkJMMSvMM9E7HgFX67SDP5CUnxJ8HoBDBvINPpP1UWf1jQatwefUv
WledUka3iwuQOQLaCLi9oeIx2Hk19kdu4Rghhd9vrS32+QyZfE2gcCW5d3MWQV3TfdKaGsmJQ+3U
LgobY39vkhFt5HOorEBpDnFC5RY+Ve9kVBAfev/lx6DS0M8P22R3MBst9Im6mX1EB8BExciT8qMs
sEeT/5eo0H7ZIjjbSHjRa1sqyxZHsRG1w6xQ5NbaAC/PTMbfvEsK+TN9D0Da7dg3nyiNaH/xTZO1
s9odxni98uJvNvheoMmso6gJdg2Ln42eJKi5VjHQbwsK5c+9pzFUS29KjXzng4ZNN6SrmjQ+omC0
QgbXuJqVUFBZOmO55d/k2IY7WyDSlsFGlCAEQmvSK5sqB2oYBI/fXOiC8H2FpfwCN36pQx3IAFpA
iN8PmnrXC2mGI/OET4Uyb1ICwK7Xj3oAzBeZxf6wnoZjGr+Tipl0pCtyLAmiEdL60ZVIr3ZgwjzS
T5vhEqM8uiO0qh57PLA1KdydRg597i6u1eoPM02jP6uJmujiWW0cuiKZks4vBjM17UuHHm1Wf43i
s4/lxr962+i7dr9KGAGzrAQT+OC1XxrRLtKAxNAa5qkRPSNVFHDerUZENFTTiKOz8X9mEGRzGSZe
InIXATDNzfIDAIxGMVnDW17n3uBEA9Q+qwtn19k97rvVb/jBBy89oeQlq3eTFjJ9Nw6zOriCjoS5
tkPIgGIjXsL6rh9uJjfLamz2uhDleraVBlkgcN5afzGRr+5INI/ITwaIfeeNkl5Wmq23Fz81dgyI
Wh0JtBweFAFVE5GXZGp0/UltxpjR/T3YyAmLnE2kG81qv5jNX/s6YY4J6/hWIaBKtcK9Y/LlD0Aa
1dc/d2AHS4kMJRttynMrj+9gHkbMpWrkQg/yFLE4anc9DbNUYiOLnsozg0T+QnhZODI3VWLzNJVm
ekUdYLOOGLAJMONUw5VBSjRVjM220Qao/8pqrgLDDIOChd1ZDzRnzqTi5HCekyhdoV0UCfgufvte
rmJTShbHX6LEw7XQUHpB1/KfnG/tFP2z4+oLW5kIx/Zf2h4nZ/Tq76KvslDQb+wR85F0nqQ7W3oX
8NjnW69aL4xI/T2+JmwNptSdULMxNNckL/DbKzlJARPyrmcLRAh34VAS/MpZUfCkSqgNExdtgSHp
omLHRIouj9tX4aKzV6sCXb+EqD97AJZHQlK9R3gFL0+ruw95t+LAmtTauV/mkSTlzU3mfAbiw5CQ
1vEgUenaBF/c0vBXsCQ0EYTqcl3iiFVrbyyoLQQCZKUa18r0bJ4OTU5JgGBbgkWfiPSPdaBIUwY7
tkX3MajsSQG4hmCvvcg/jUZ/U/UyaeWCtoFhhXBCUFin+kahXGMveEZH/c2yczUkrHhqjEK0BvrO
68nECDjc1qrnzVQSGXBE16y1VGu5NTq1o3HoI/y+qU9UNhr3kSnTNnrxYoosUnf8Jp9fzrsywMlm
c2da0xFeE9ioVvavYBTdLIkomZUg3uV7gFlsNIDbIDJIMLmpdNg3d8BQ9mXY/ZS36lHnPhYGp+5x
tw5/dy7Xvi0TXzLhyTd/kIYSytSY6pt85DkvxjUQrk3gRcKIdO0yO1NMcLH1MXdz8t0aAU/xnULl
yyDciq+rIgMnZ1SKw1bglZIxjRCLaHwuyHyK7/G8VU109zpiVLQufgAm4tU+ZnLKEgDwMWTwioDn
Lghip+2186fO1FzhnAfgQ7cf7qQuuWmcUy9Q/sFTc8QzbJOYIQAp5JGxHuRL6bvfNak1UfelJN6p
o0GyfgW87j8xV2g6oQAxFAmukm4UIvh18QrLUdPsJ4M75ULctp4LcxVqcwE8M18jJwas4N4HvZqO
N0QuhLM6RYOl4JDQs0Uitjl4fNsJFgoHZuhUbohZ/FkdxXtq0k+CkdaPVei7ICJUahfpbGlE3aXF
XpEUwB9xy8Eyd5a7lSNQpUu/atEzzYNiQzRuSGlL3D4Lu/wJ2poXqHZyvi3F2Pk2rKiOKEDPLmIC
iA+pO+H+jAFZfz6+zJ+j2s/+X9tykuvs7awCknwSzZaI70HeVD/UDaE0Yp/qlLB97luXs6+evtMB
L6KKzvNDM/k/gfQxxr5YfuPS3U9qvWnJ6Bc5HhshYpKpz/ux2H/dcNJb+z7ddbBD180MyNR2OpJc
vBdFai4+MXsdXIUWy9GnVg5wglDX6NlqfBILcJLWak/Tm7pFvAEhxtXUmhymWtfXccyp+BPK/fYg
Iczy1MERUPhG4rqUdsYXkvQSRPxxEWTEnQXo3B6F0JRSzXKm8/qoNawxDgLiDViVBHXhGphGk9My
WOCOglCcKs/LHn7qU7euTlIuXDqT5RNac8M7k9dBywsRRHIO8prklXPtCW/HDDmp6ZeiaDIbZEnu
HIAqK/OpvfQVObkZv9mWrwWdX5mghIi6LjDUMHc2nw81OsdSzAI01lFGbrO31K5q8itsdIREYO1u
rZ/mQXH9HdBVnrYj2qKh3JowgmQgPp5ZybktUToZQALjI4JhmtD+PvQ+ymggXpdk1gj1A1rx26K4
3mADsBDQtCnedoRwdtvq3bnjMn6gJCOoUVktEXMUjeliBflOw1cgpbqGTE670C+G5pnMk7kQAP5l
c3TRSVSgGASPIqfTcNtJaJ7Ms1TIL5VylPEH1ookk1kQNX2/0Ud59rs5BhwRcd5dB03UEZd4NCxg
dIvyBQRJil12KW1P4e0udBnkb/yicsfZMPCs8VYnBGncLpCSH7/faysUWKfXqlsjcmA2wnQZjch7
wMebrVKvB1oVL9N2Dh4fIkouQcv4RvmlFDN0eSQJ9cYvKGIYmzvoCVIEK/MFP7ky3HmqU1Ec0skc
okBEz/zrbraq+kmHuPZrfQHzzDXXFcKt6FM7nx/9loVyR8xAkiJQLKITiLAJwlhuu7i9Fq4XSBGt
fIqCpEWV+wxH0zajAlTvVHy/+Fwk5BLfsWaU97tRKgShzKXRjwv1pmEmQDr4BVMcia0vjhHNT99L
0rIOOubFX6q7SpjQQ9sCKabbcAa9M9lpu2RnY1JOg4fgu/pKeGLEsuaGftWtzGvXzubGAcYwFgSr
15RKbO4NXr8TuLeYRpJ1EUPzgNdH6G65G8jpaz6/AoXstI68hjnglofyEPboqkIjTmjzOKUl5hUu
nLHO2E3d0WqfJSW/R51C8nt5TnZEE2qKXZWD3PKkAQzoWkkVjfAf1KXMvtghPlo3oDzoN4toVmcD
kaeOKOUJtvExhF32HueLspNEqshLnFXpfaoj4tfIZjLIejjvChCJMgaeUWOIlnoIGslNIa63bCWs
gIR0LDU46sUqIzV77gvaXshwt+rxLcq3KsC4jJleAAbSTqrWwQANMFE4pjKyUj8L6mwriJWU43fK
yXvloIK9Jo6uEyj7L88KZ8v8No3jOlfq6mj4yMTMT9wYoF5dE4fM+1JkdBVCyjYZXnuCueGSKoGU
cZGEDtWVfPgCXuMg0QywrJE8M7r0W/YQOsqW+4KKO1rqAzlybtjVnv37PGCVAJoImCV8BOdRw8GH
tB6RRVs9NW9Tk1Ewqlbq6v5ivprK/Q/TQyp++awBKMnDH7m2ef/O8T79zT4spl0QketRJv56Do8W
aR7dmSzEput6L8kWAkyn2mBqOezCD8qjWhGiS34tFtsHxPslocWa2varawmgfwcpZTuwwchowvLK
aHRC0U/PAPAbtlCE4H5zLT+c7eZ1We/96ha1k2B/04NwWIXpV1GA6+ncVNzyf2pd7lFceAO5wk8K
kIxQ3TfhzF6wSgvC7IFCq/zvhhowKdBydrOACIserkdb+ckriK8zWFfPTnbEmxVGOzCSV/lwOVvc
AjJ9qDuITcaGzKtbPDXtikqv4ctxufwyfsw0TUwKKP1NumTmV1450wZj8Co5X0s/qG5roKx2C+Bn
MYHZnuKHXopypDRtD6fY3iBJaJPWuEipOY15Az0LsFVaQoZO3X+r0Ebl1W3nHQ12vNPw5+AyMhu1
Oy9vaaSLu8GlGbc2N870PqsDQu2vztpIoFlaKFjf0zzKywNG/aXgd6BM8NPRDNkvrr7Cl3HHmi/q
ln/ST/NdL+4Cg0KFyaqhDF6emhQWTdmdFRXw/JSUATw5bvyU5Xav98U7kcorZXGL30tnKbmaygqT
3CxgVPlzf1YSkKkh4AJsTbcN61DXA4KFple4KsLnQSdZ8lk9hLejmzvAI9GqkUsclZMJBgwCwXmJ
oYZtlg5lsdnyKVgUj74thbEaHkffg6huJMd88tgFvyuzmAcre65apB8+qh1DAgGUY60qfcN6WycT
Us1S+gLqI5kCtTOwHYSB+fEWo/WZrUkCW/hwBlbPmZLg7y8LSu9gqoTM6M2I5PvbbLSQfuEwFZM1
FZQ5OBhwWNGrvyOEpXUcTO9PKJg75cMWcGD1x5uo7dEwDo64lxFysC3rO/2R7a6tmM7ZUHx3srPu
ediS3F5+Q+khV+FocZ43byCUR2IG4xxKvvrqIrj01nc+CbFyKItJC5eqeAcpNDQa9wh31LyGraM0
6UItp8EaPMRykxFndvBEu4MFzIZJ6xXC5gJAA8y1hr6N7fYjnA37ooJTNSG5m2IyLdWBjQX+PB2P
HblyJgF52QCbXU+MOr1p3M/XCYAYW99zh35ZuN3sgdIRyB2kW4z6GBxnK6AMirT2/8+chDH2oto2
mdS/IwiH54XBm/7cs6RU7C241oU9245RvRz7+OIrOv5xkelNowySoegxrhh8hUoNPJ0NxUgimUBn
3SAhDhjnJfljwCUKX+tW2g9is4u7QIuxS32FxB2rN4zHrhpM6EyDJtYbrcwjsQGIo91/F+eVprNK
0aghRwqJhD7K4C8MBKJxVTfBCAptzro21KhJwNFI72Xstywl4kQ9seF3yHj55BMuR2tCIzGdzrEU
ckAW0HWrPlpJOiUWhOHX/q5yircviJVCUACATZJY6cufs3k8fhv0vFAQXxavHEpZ1cRtDOali7rZ
MHQnWCAQv0/DcLrIBtnnEuxl/PFSru/nSbQFC1za27CbHuY2B1Yw0+nzmpsjbza6p9CpuButr96T
AoabpKeVSwZ3Q6hwf+E19kFkf0lB00n91JB/85WIyMan/yLeDs7mrhVc9eKLc7kOBWsaLlNfm2xh
52lBjh93+t4R9X78I89Pi8k3NIBQ9o8TB5lvkBDVIhgZGypgYcrnh8H0sYpEpOhRoJqU1li7SB18
kqhfdk8eYRVbdY4ZD3ysFQCSWOhB0l4Z/TUtpD5gsaVxZMGTscbdZqrsZ1Ymup3pSMAS1+v9hqul
5D+yYso5FOLDhTEzK3EMg8U25hbpv+CTslfXdmrM+FghkhRU3OA2dWM8yB1KfaMbQFjBKxJGjkWk
25KKwabroLd3fyspuNTP1gmQC3orYY2BpVABM+ybF9Qfu4tyKSDYo9Sda+4AOulvxB5DsV+L/XeU
UBXi9KW1gQSPy91FYLbXzj1EWdkJvnPjWp17LVCMW0Kj9ScVugRuhrtsTeWdJYWH7yR30V2A2vo3
Jm8s2DtHaB8Z3zcb5SsEL4r06D2LGd29zLNhyEFo4MhAxgODSZsbibWu/V1RPZv2qZxzWBB4wEGU
JMdRA9A57HeIGj76CL2YwqgCO8phUhsGhtz3SdNJTmZUmg67uqSCAA9MPyJT7JkTLs9JdncKgB5+
3EiVNGUxuZDNUGLLnHzVm4MfyjLhgy841otVtuK19Dy6Lava1IOwBuzUTqDG8tbBlDY///Ktq+58
Pek4LxXEWjy9yB2NrnWk8LqXHvLjElt+hDpo5FeSJQb7T/q1ccoeQelGdNE0wRIDdA3ru5HPvx5f
C2/axaLRd12CPwylsKx7ABbtTHLEQ0P4CtjJTfiplJ/08hpxkrJF7t/doQbpDLhh4JmDvMtuuOjN
hv4G0Uc+Dk+4zgNaYnX3vlvD3uFlsOC9bAXq9bRilsTJS1okQnFQ3yVBkYQsIhv9or7AIvqiH1em
6rfXYJrt7xaN/JroGMcoK6/qXpcS9jThlaozAntdeQQKTHpJy00MaTiSk4mH4qZPb9kmIu6NKeCb
1ABvxGNMniPX3UXyVa3oC+H9SZ61ouvsO7BmnaXW1ft273GWV0ZZInH+QoTBf0gZGbAFWcGDz9KY
zXVa+p9vSN/dDaxmR9bEYRGCLRxBYGBGlFF7dAy/29eo235RliywVTRZgCfOOZNpcRRsuU5fVyGN
YgHLLe5rJnlg53Pq5z2rpYn7o+94wEw41ewl8dFwgJLTJxq8KbgiE1znl8DEAo7uBNvOSKz7A31p
7nGKgn+j8b/mRXHz4/JtFT6vgtKqFvjoj9GUBVGRdUiJauSCCVpMCzinxH9ibfX9yBhjx2ICiswN
mM25DaPs+a6xfaFfkJ1YE0EV6/dgjnVUgR44mR4AlDY9xg68TOPuofdk4J5ReBtbUM+qgVtXxby5
WPOGAKxw+Q10JRhGtOQtQ/gpu4PKr/4vU+ope7hhB9NaiSS9fpXweGROsn/d3KwfgiKHEnz8l138
ii8qswuOuhEvYdZextRgmbte43RljjOLUPkdSpvR1zP5CHUCi9FkKJw/pp3suHy2hkEbVEELm73p
exjkdb0QE46Yl2RcpSNz/C59YtepZUs5r2tVVCxjw5jcAJ8qV3anrOkYFm5fvJyXsbpOC7hfFHZh
nDZBGWx8adHM73Li8ZhVkMUKrPmS9bOXmG4Sm3M8MGVRfWsKC/zcfld7oov5Ijr4Qppreaars3xa
rHiq+zrUh7/Ux71QihUyJJrzXhApszFLQMKy4j9Xe82yYQUbXojOHV0igJ57G8UEg3d+BdAkYeM0
7ACbDuv5b+G+/ODWpx5SQn3zmNoeq4ZYETy1aWGTjYK8a0y760L0FBrC/SvSpBhNhli1V5yalrsr
++eWmS1suRlnD2dRVvKh9TyfmtmjEAn8apk5TMu9jbiVCuTQX3Dx6JCXxVHMfGQN6hfVf7IYf4oP
OTMO0gLCcOoetRUEoWkBV8T57lQUwx9WinrD/+R0e813ayqlral9IfmnRXreOh6hHJv1VNmtr/yw
+z4+xSEBnLiF9MDUvK3th+Sv9cFVsV5wN6Z8cwMMT/Xm2M5nN0dnBT9gZaQyC+IG37gGG/XnJ538
xArTglemycsiWPAv16piKxF+E1rbSCI1/i7fzMbvqPCCihEBtfexcSl9NUPCSLz8Ib6uhBa4a9WP
FCnC3JH39MLLHatB4Ttez7xavblsCfSbs1wrdw7EnhwwIWVq/LmEBBWmgW/MDy5/fioLF4Xecze4
3UCuyMGbYnPUwF3iPgCPHjFxq2besyacBL0gzE45hohjBPTknkefjzYXzMxZ8FpLLOViWayxQfN6
LgS4Idvg3ltMDb41L7o1lk25ggkT8YxRkUSZahuvlvFKCwZcMaRyFXscv4Wvei+VlvYCgZQDhnUV
6a73jfYkwxsdXbE8HaqyJRETx/jsbGZFlwLBby4w1eiThV55/Lp5KzNWmYr1eEUQdrk9zaBrfeXI
+I1mrWJ1rkVgO3tt8KKHC4c5NROXUYzsIqlxh9982hYSc6lBeO0Io4yQ1IjZvlnUkL5lbDuGJTGk
PLo4BqWuVe0rR/ADMW3obBbYlqFx13Y482w6rhjN6RuGjAa6FHQiWEOrO06GjQGgDg18wL7jlxEI
9RHPkfj0UbLsKqBl1P2MLbeo4ii4JWlI+p/KQpjiGFAzTcaQHC8k/TM8p086d8VJGaUTBCv4ElMi
Z8LpeBQPN9JzmJMO1PeorWPbl3NSBLQAdi3kJkhlv9KiaHzsHMBeDwwDamOb97i/xqESieEUzRiw
A/J3O+X1d527n/cHXy7//BrRwNQs5HkuYTT5y2PCfAEnR3k6qYJEeoXVQtL0yp5ARwW2SMW7X1uT
9LxSAQxlo1gdAHdncZzROB1/ZhW5MI0nSCyjGrgYI69U7MUbUO/X6+ag9hvyR1bhtqOxhGi7ifYq
3/RIoJe1qjNZdsXA//4fnOn643Cnmu8vUpF6hkEAkVAaDgSYhBh0UqK0iFz8cZJstUAmE0OekazC
kcgfmJli6ayLiKittxwfSrvi5DiLD6hIQehIzSg0gHG6nhN6Fjnr3mxDb+5E/H4JbRksFN2D4gMZ
xkKIxvdx3+ZVynE4v+05kwk9XLGZ26Q30SehDpWeJGQzeH0ZBCTTD/arVyEseGKbkGIbRfENdmgt
TpQVzDl95MgD9kyAM6INfwAorbCzhJnGcvvMLeigJ19DPBaE4P7f8l8MOMa5Ehd3NdS4RQicJPy5
uEFqPHjrcufgYVL1fqJbVHcG9SEka0F1N/+lqyi1/y7EqCer0eSVYS+EltGBqKlZ33i8zFpP1vdK
YNqFVITb7tETlavR8okqAISLgAFeMuyiRXWzkYTVrckDmrkvkK/RFsNmL1qL8RRWFhZt/ET0Z2U2
JiD7pECdvTk6adBstQ7G2ddpl0KWLdLFRxoH5aQbnZ52OEcHKCHQafFDdRyYefStlssSbyka87jc
FWEvegGx1G8cwazNcUyufDMtRwsTe4RBk2V8LhCC1f69viu9G2+MgdWFLUJFGxBjbqMciXoEG6YV
/i6YBb3zByueq/qvSSX8EyaMWTCIHgryKBAeclNho4XezDJfF3CC7fr+NYN02USeUA6omLMJE0Cd
V54z3g3mb1OTCRD4SQ4dAk7j+W/hbHFH3FLI/rA8b1oQsP0UG6aPxGNubnAybAx3HWjrr/D8cCK9
osHjq5IslKsYUNQ+TNys/UHSErzP62oRPth+8smFZt8UE22AvpdjAUXeqnotJmxPMeq7+hnZJl9y
h21u8ReZohwXeC3TParfVUV9CwN8g4VATA9bjRfJ36Uv03kW6t+2m38DhXijTwi3HC25S6/cN8wn
DQHtGiGQ1E4ol93ti0zSpK6Q+2PQqOfTOb37zK9XZGqxjTFirBzUA1/mTcCdGQZxSPMsG2t4J+DE
kwrhZ1KBq+NKneIT/kQ/PrrgLTWPdt4r0DN2hJja15C/dKMH2Ism0s+DlpnvXkY8alHeF76BkHbX
AVeBO9LNnZcj+eB0m/itTlnLpjaneEwXvNdfkGwAUBnXs52P09LyF16mS+c8NBlUNNHgPbNEa/3Y
hnr03JXNyxx6UdbC+t7JMfQ5cfEbapbgeIKSHXZYdfwXc1f2rnJcX4dM9wAR6liBFMRVmGjEtSLq
kLroOpO94nXdWcbKI8e5eKj5j8snUqtEQTA+9xuSJWND6VfO7o1baQKRPiapJlFkvdVPogMqrLYp
svG7XvesgZ51M0LtJf54SXZYCrL8+gQrcldvAz5Y/he8Cu+4tWZCqrdM+JfWE9EUgvm4KrObWCVQ
uHZzZrY343td/13JHLCWKot/TIKkWKCiN3hXlZrIFOLUo8CCLk9/JMH3cIv/EvXLTfhqLzCtDg87
GvghNFtrkz2ebpNL1nxqusC+6QQj8jWJF42L1wJxG6xjf+Kh3T80yCI4PyRBCW3Dt0VvHAPL/OdC
p7V/+4cemjyVQvFJUkCh1D/hVPD4nwbu3m55g2uShWHJQ4H6a4JTRiA8b161+0M4RtjGGGtOmTDe
ywjB0fCx2Kr/6RZdSEiaBKiUODfBz3aDdGclguokVduD7pK6KBjLQB5eJ7McnpTRo5xoLdb1DWm9
9yhnuDRJLs0xbyaNeuAo+v8OMP2JsZ5Gey+iOOxWgMVGUBDOI8AKioUy8yTXVL1+R2WVtGHsb/qW
CphN1EOimZsKG2zApn7m0BH6V9fSkeUuf3qbH9/ZCezN3wmzmce/7fHbmdjo+WyWpNCMVHPDMW8d
PZoCZq6JNIcp0UzRHuDgtxBaARuTU+Imy1wzbgYJm234GCAORDUkgobmhqG0MANhnUK8HbX2uOU8
3moOCvhs/FoKOe47TI1Zqwi9HwuwvzBNE5ddjWN4XNUGXJ/NqewxZ36k60kTqXXqu2wB3qem7a/+
lfmC++R2FdFGUK/DhXO7ZjN/6v9E5QAcXujp3MHOQLa7/N47KeNIM7xKGKcANe1E0SVyv6rlXDPP
iiu3u1EYGdUj606I5PLsFwxF5OWnu68GNn9AWVmRRHLPS4UV5d6Go2vO9o4ecnioqnW3kk/EkGqJ
TAgWwyfkA03TD2+Aj/any4oLYh4u/nNk1Jo1P8PDbB6xCbezFkJObxxQIc88lD41anl+0n2rC9qX
wCWmcbiFD4wIh+cffJVkk0adlkNz5ypSCfxEGSZoCIWBFVm7n6UHeqQDFYKrXRQ3OXDhCLQxJj3+
qg1o1xAsNjqSPYf4LB0ghTuf7ZZmODvfhRfr3cuFAPA7KpYlgWxvoILncCe5+Sezrp7mGlVyJobN
xWHANpemiH6okc2FiydUCOxLL4dnJYcwQqJuR+xK34T+Z/yQHyTv+Co9oJ0lg0Bi7B2Bck3Ls68U
137zdc2uS7rV5sl9ye/6vgVZ1DQvvXHd2g/c/XSn2aGqFEMht0ZFJ49Jk3aAaPY+6nlWBhZFkPb8
5l/Hsj9Z2XsvDqI9tqwGbRTn0N6/ykCx/wx6gsqtiAz/jSDrP0c2EWFYVc4KlgVUl/gaU4DNdZR+
DEbwrGT9mCfSugEhK6rDZa+WdzmZPUouDTFn+lC0LpexIlLhU4t3XbztMIQBIgG2NdN+m+PAMt95
jFm69u5dXVl8om7dKtUhDTuAACD1U04seaf4Co0Iwahw8LoVOPLJMmboz5GHHvDh24nLArfomG/F
EEi0bKAJSoClPwO0Y+xIprJ51Ki9e85vG2UidRGPz/bt7pGoQ0W6yj+RF5RE44iDDcbOHFlglk+S
RRVSZOj12lkBfrNkUt0ruJYXzKVv99SE/7at0xHRBpt8mCNRRkCjOwRj2y8BGePzI5RKja9U0PUO
5AJ8zYOLqXTDnvek1j9FnRE2iiTR9NbB8SW85/+4Di9BqlVwnrJmovuqQhepdmZ65exvp2OaIk1a
G2eqDv48nXR+xnFBdZcNM8zM67+iG+9owAXL/1xg6NG/yGlc4flWNDXzpRx7cTVl38W8jYPzruti
1R/Uyd3CWRelqW8fslqZHiCEG/cYvS7hYAsAsO/8An98XrEP7RlBpTg9rg2JUw+PBWyNM22iuVa4
ILAG3wQ2TzX6xWDKh4IEnnxDo8ZP0BjAzSnqNHDa/jJfdZ/ckBSyvEeZOIcaIvQkmHMdwqnWN8K3
VEaSYWXXP3gm/l0ZPuvLQSX0piMEPJHRBK6I4zm71MCPah1wLdYhWfbQd2VXpLAFf+KWGpsuMWqw
7l1H2ngFn54E3XcvgO0CnwgxQ4Z3n+/SwMQ/Hnsl7Z5mqIbCiVsHZU25qdagCEajU9nuIc26IzZB
fb1FTX3HE17U95erA/ab0FoFbN13dsKTcIxWhQpC2tjiu8Ti2lio2aon9K+lruhyRRq7NptKdQdw
Rm/Ez0Tfhp2QkEXJQZUxUQlr7OhUFBEEdaNB4/zXwzauj+1Aa+M7LqxsO4QTuKF6MJViBjsl8kNz
Mdetly+zAFLkijCpHBBxicgtIGFPUZ/rcZ+UNXqg02+VOOZZU6DyfxXm4NCX3SuLpywtcI2DiyCX
UQKJip2r7F/kKGcG2EjNNsX7p/6AjNQvZfLMA0B/0xlg/qUlscJD4sTz0zwTzxAhjmIwVDiJOsHV
TtVQrPl9ysmZTznTnpjNujD5NEHQYfVR7CCbUUAtCuk4s8Yfp8QD9wrm+cGwvzxEVchtnLThDMwe
MXBS9Qxn0wGo8FmaaInEScNWur5XQj49t6tMSw+/jqhSyvw15Qi2ab3Xpq12h7CGSW1BdrHFeVB2
KdgEu+H1lSZE7/zlMtLYSXiAAl1M3vyyOJqkiH0Dme4nYuBvwunF8XiVQrUr2NbvzCO2IX31nSId
ryd678L7D5xTop2Rnor9oSkDop9EyRgt2xsKDPHjCLSn29M/s4Gbmu637w7FA8DopTE8lIQI+qZi
Y1V1XhRgkb5P0vNFpQS4F6VqA89d8HlqjTljVGgIXyX0zQ3JN0OCLySKJveNfo7CCZb/J37r2OPO
7VlSgCA6liP8CfmEqp/2vxQqX9hEmDLG8tOs1dkX2S4MclHc+HFmjMz+neX+ewMt4YrPhi0sHb+0
KoWfEOfDMxIftTW3wbmNuw3pzX3ovfiXmA4ajcwcJip2+t4UMLnJ2WkQ5K/RlwmPoI8cR02SkKq8
OfMGMObCMA3ClOrxtEwUHSEE3RnaCVsNXr1jekbjL8i0YxFLnwDMIucV5PW15F5HwV/BkVVRp1Um
Th/5l0lTvKVy3M+q0+cJcqli46JgvoWsY8zgbQ2PS+mZ9YupG2Bqxnx0ATohJ07CnIx0fQSuJhjf
J5gppWNoQmGoYJQAKTIfNR6JgGCr5+REsLCbaQCfmrM7jiD7/kvzS3wf+MfqegDoZqKSqVCm4G3e
wqvxCKCHNALcGv+2ftw2PFlw/6BrtV5cDk7hoOZsIS+68y6ImX4zg6I0748YDN1TQhE71NxT+Efm
DXht2HhcXEMhO8oOQqQIcJO1eL+NGl1r6K6MtoyOySWxjXWwLUe0iO8tcZusImwBYpDnh35WSlgz
MRHMGQszvfh2+FmjXk1C55Zbo0wOlaB1l3iLJODTqvnV83GSKx1XTfYCJVXgcLbgiN/Y81jLfyjm
S9LZd/OQPkIEOlKqBaXGtCxyM7o1/tSasn1T1hJ1ix/R2nQfUfXwOGKkRkPJpSESgHd8GHtXbmZI
rbSy8tOo6W7Z2FR2NjMFh8MOp5O8BiXjFeOY35qFKVnu72sBhsU7nEm5Fmcjp9EGndKj6bMoPQwr
Nzo/x+vUVZD5VeONRW5ha2GfDH6+TgXxLSFICTz3HzLcbKS0t5DDTrnJOuJLQeHcZs3IfO/+y12F
Moo5v53xJiaxjVCZB7W2TSZwTSzXIJLP/Ru+U6es1tE/x4xPuonxIvQaYercswoRCUrZEm9U4YQ0
tb2oAMrq8YVFS3Bb21Ft6f/W8/jL9+TWWzKdD1mJJAQ8AaCMXVhQz6JFmM6fLCRFwOXhiO5b+dty
WPGwYxYHV7oY+e0qu3Vuztk6ji/I+kBDX8R9NZGww9oWB1m52uLhB2RMwX5W8Mmxhsw2garVXqqN
bEcZpLfzdSZkdWWlHhV4XOhuUiZvGI81AtwNhTKcuazzY280TLYP5qq3hR7kusn5f6bzIFE1ZZmo
/mGvQeLUdvwbqq0TFETslSWXf40jo8fImB1IKOOUm4dYJAmrB11ABctw12tE1xGKbvvRgHOCC1V+
eRUp6OAcR3gXtdBl1O/Sv0lIVkjtCQsZi6oZ/kt7ll+3WZR3Mj7rpxOPxNx6o6JlwTeR98nKjLYj
BtxWgbDN6bWZYyVAvNlrkuJVoO8+47TRQUGJROCKuaY9IUB8eSpUzTLq4XiJ5W/iTF4J+Ib5FGFi
PLsf0j/2DNoE0N75ntpn1LWQAbB5fPTq8J3Nk3Lb1ok1n1gXgQKVheDSuL/vVGafurBtZpSTb2Il
O0KyGsyMbA2hq5zvdjR0jUzPLXtWB+S3YGlHtdDSbN6jnsSWMyyAO2ijoRdy3acUbkT346X8RM4v
iW11F76m+ZaS8qj4EUcUYis005jnMGWwtAC9rDhvLf/6YjXcti3xmCeA4Z2E2208hN7ca9biASZA
29dLNekCiKMrwDXONAa1nPJFFyGPTxqbAxffG1nGx2uCM4Jsqlf/gTsjrW+i8zAHPeKBiB002lFe
2III5jx8k/mnpYSUtQBswnMzp6nYss285/jZohUEdiLpO/BAAfX5ba6gBu3MLvo2nhRudPiGfn7W
y90GkaFH6/ew15bVbLjFtTR27PrNKOcK8W78n6CmOZpmub9rPIAQUiv3laoi+DMri9IKzuJQ5zM2
LBWNQcwJA/w0ZfrA5kWRWMBexFOjB6uJxuc+IIwgwH5aelEvMaUiDtEeCDyn/WiM7IIb1K9EygwA
vMoT/91xEVbwSATiMeiXZINCyEGRP/+k0BdJIGsVSbbgR++GPNFOhEbYAnzyJS2XZbC59zm0Yc8r
G+9ZQBDBVrq+FED+8LI9Ff7qDdqSQC+xS+ONsteJ931fmr0+T5P9sDWAy/4vuOcVDvZQkxw7z/yK
iotomKKshmkyMWVh7P7Cmfd48HX8WCsa0+QBbhpq4hiF/C9JwR5vDU9EjCj1VlXmKc+Cah3iWdhC
zSQih/7cI0dhD5ps1kQxzK+EKe/EYPjBqK7pVosMtzAGtE9TWb2WAoQaPUVTqTtjcSh3cV0TYqgC
DW5Z/9opOmHgYWksRA8qLgLmOKcIp8cwneu9cHBSoDGrhirQfyhKpIlg4KisyySTUWXZWKj5C3EG
yT2A9k8sMRd79EcasXdCKx3L0lvdLmhL9Mt7A2eT6LFmRJTVyD+rOfy+c+crDnUYEsqg/7MnGvfF
A4adbaxvJfU9AIAIIMGZaAYVdxtBjAkh+mVFIWOPUi3xBY8zqvDkt4dpVh4WNTiLp9Cak2keAF2i
1aUDnZ+OcMXGN37cBTjEfNTto6aTXj3lD60a/9Tkx0g0CcRaVtlh5ORZEw/peuNphM9Z/C0wASsG
PM8K927bEhTVfyIrEkX4IBtzX94ECrr9HggtwNYvPMor8W2mK9UBxY7KCnAKbvUqncQ+BqPuPvr6
tckGagkUrsesDQFTyFT2aLBSW0OXXrgeI1mlh4fT5zcc2e3a00vc2ln1qfJWR5dKLNiPIYQvKrMg
pNpiUFMaQZWna4/2U0v2n9Jo/SMLkotaGIh6rFFHMjTdc/jtA81BOOGThBLPgTxC18y2Zv7MnhrO
u828znB2mg23tickd50kaReB9CCoFgK4s6BNx87iwzH++HHNb/xv5hBL3cA11pO8EQHnSm7YgXU5
pxw4jIwMpbAukphCTN8omSKvcLvECM3MdLQ8DUA48EaYPG+itzdmYrQbZVJWp67dwgzwE2YxKuUp
oTw34dAW0QfFjP+TvayxIsafv3gKLx7dw1U52XHuYgNJOEmNzNrt/WZB+NgseKCXk3C0Ud2BodFA
vGsAu2Wnv4E6SsH/pGtngC7Qy/DC1Ovv3IpT0rFuQHYCZzxq0hTXRz3iQyQ8SoXcmzUwhABxv+39
5enZ32R0lUX3OkDGWcINQYH00wSGe4EqEJN9Qo09x0RwmEmWO+fwIXt2TzNgCSN8dE66HD7NsGpl
vo8PwtF3OlSnSLCPQxr8bQ/4BUEOj74J5zoLHcWrcqRU4xeNo+nr4clbhkQ0HvkL/qfpXn4fHZBw
pM1pDGjdIQaBpu6cpNCs1tWtAAGs8nZCQkAEG2Apk6zz7v5XpEL7HRQn5m7g36hKnRVTkGANa0vi
vWlft5T1cSypBhKh3EEPLREED61xdz8jovlTqwSyRo0MP2it4M7KqUiBKiRbCzgqQ2CptqAxzXS1
zHXvAxkqIVRpXZpU9arCSZYldonMvd2zjSpGagCDWYVEofHqrIEgclOBth2S/03QMHgusLYPVViP
F7tWNstR+b7WRyuWu5zUjS8JSMAigz4LhEgjfziYCrsBrPGbpBMCYjeniAjI39XoaBE6W7rs2ijm
3kHxC2o1WYo66WOlTJccCVA1n1pYYOUnu37pke423u1JQnMRTQNnkMDgLRbtal5NXimOvPT8uV/I
asp0T1WEW23sWmMZQ5TUiGZhnn1WMzSRsCEQvC9tGZTQaKZxq3+Du5h7Py9XsOCKO7VpokExgMoc
rSjG2QMczoPjesrsJL4sMKt7hNGA4mm/HK5jdcfd/psfcbNPuBHiOrTPK0rtzNnaKNo5pL2rC3RE
E2+lCiIb1Pal/WeXiwJakizvS3L/6cnqk1s8s4F2YbRAC0iABe6Nb74JRLV4ebkBPB1MnYgQrwdi
W9+eK3+UykR8sxq+pjb948ntRhd8Q/fOLHtykDdAz7yynuM7t9ql9vIwr62umwitiQMRZhNoDWVz
81HgjYRotYdtXNPpcZUql5ZZNlN/BRVYb8B6TTGRHJisdDsoEF78UJcLslosdGdkFaoRGlj4/Cpf
U9iBIQzkBOjHRGUTkzzdU6TBVst9b0oky3SucHyqHsrsbZmyCs5ClIUXd6b8G7navqy+eu7TCi69
RS4E4EQabB6LzgC08/+XwgRk3srXK1/CnJH8Dr5bAZBmA8zUQYw/xnpkMRQJw12f6yYrgR1Haiel
6kYdFK1ULzBAO3wjZ6R0IZH1c52VIzVl47ME0mGlqR0n+jBdx4pGkCjll6RzaZWTmGJPDqWkJpHi
CbfQpbL0+1oSs2oqgzx0/ck0bus0HpqQST9nwaAvIZDqrJ/clrBudUJmSqhbPUuu+HYUlR+AntxH
OANlv2UbiOTXc/BESbyDNUzbvqj5FUS+npdNglUz0vsOCKaDvImbeiKUrDUlxXW0mlDOTrtBjIkl
NtWjDUxKg0VdCZOR34cepc/vjjPsi6OcvmZTXpAFcX8iPmZJSymMKWm4eGKKQFOdrpvvYhQhNQRt
0lyWJRgxp7FT80Sp7mywG/wpwRuWX0c0lKKEP+DyAbkdMxG/KlY7rV3N+YCJbz1CqlpcB1PG047Z
GsMkKfJPYpdRW6CQo01Y9v9gUR5a2NgJ8c0cC66CNKjImxUM8JgmHMC3ebkc+lL4Hfz9PcULIQbG
btN7BW1Qu11azeZ/e2yN4VlZjMvrUEBBbefW6jHOb/WR8EjChlSKTyTITOVqrMtJND+RLL09MUZo
gg4fa7bhRLnORccpzt2ckSy8f+uErcIrGgR8miydwSCB+XXl6RyarbnRqfnK3/ni5MS7RaZp2vqp
eFM3ZPXVZMWMhWJcHj97CS8HDKHedDXc4j1FS0p1U9Q7jFJzuDLT9AFyKcm8KRFwg7hmgbcf/gL9
cYAHVBS5hhAn15CjCOyuUzzhjCMZmVAt4sWk/vFdMX03hn174xKuzI92BMp94yzoBw98OJjrlEtR
0+RsxvxzuZwSmrqdcJ/sn0f4guAcUWmlfsJzhhjH/WzPZjXepZGMMQ4siGoBzLSZmAJ7+sCujJAt
bXIoXzuF5K9cXZeze6KGTqkKAIpbNQijW58DXdkPfZcocFt4zd+KM+eA7flEgr62Av8kn35x/qoF
gS4zVI24VPx2nHraGySwl20VK68cIwKSzYztKHqA52Ixf2htvYPyiJL/Pq5I9EGcwOxo78LV/OPO
0ZJixsgDk6W+Y444PbEvwTOAatnZ7FaOcvWsnYkXkU/fsrNNK0dzUc4wwpfUQuGIZYKPKPVYnYNX
P5ipd4DMBl+kcStgzBy3UGaekCUEtAQbnZynQ6wNfFS5ORD5B8Mn6NkiQoXH7unhON5C8kdMDo68
X75ppy0fgYFaGk3CKceYCS72sVp7rDPhLJNPSfPtk9UDbFIh6WahF9hdGsAj8RyLWjrPl9HTmskd
EmxBqO2ErGeSsP9x/IW9k+NrSei+oeO32fpcZn5kuzUrWEma37ckSNyJtPiz/DT/cPGpyz+zcQ/c
DA9EcCFmkE2r5gnRj85o5LbtX0MJj60juPuqUZPdtoOxwVNoYwmKpqdrFXHoJy3mMCe+7fP1no7R
xaSCGjYaFJP80LLvAd+oZAXM9u5YlLAToW7YEf//SbPYExEdf+Z+ijHfIpAfpKdFxLs5lJKgB5x7
5Mj69a39W6ynCCC0LgfyN1rQ4UrBtrw+xe/+a2yxokLjKA2QTaxhp1rOYs8gyLOg5eWdWk+JV3Fs
rrOjw5IvRrs8ljfnXmIQvSYw/IiGIL+of8+E2pauWe8S/I+P+ue0rGdGVpTZ0134KpWmRJZf5Beg
AUoppQSPWyS27Szf/MP/II70Yuz5GQA/Jd08bDgf0GWzps9kVEHa5r94PkaT+ZQMKrFPVtAZjpmr
THio2T/fJE4iFhXAA+U1ETnXxS+itnhUizATQwlEeqZOiXKKhgk/6/FK/3QqkrNG7wJZpoyw0yy2
i9jNTdy9U56PEFU4eO47+am/DiteG41vRq9QE79mbEPSPkzhtK/P1dL/hpdGAjpLSouXWj3SqOT0
JiuD8RPbTfmZ/8dCObDTNZCXjIaGVJLO2wicWNCYmh+/UWON8BGQwIeFmsUpc1xCBkDaN0UBkDFf
8FumJTMITxGZtcFQfVcwUKATI9nMoQvkjtYaUoc9xINtdSzrypwEx6Q8NqCjovUhZQEsaFpJyCf5
1R14fYstuELD7aZG5n3tklxCPq43UbZmfISNUnNHVdm0yOXpyCEeh2CW8+TSEnIePhEI7I8y0qXh
HsPXgtBP5WmlwPNXR8xaSQBjCads+nIefqpm6Vl2UgbH1wP2pa2xTScakWt6QA41+B7ZoklVBwRX
sQjImpJsoXLbd1EZbXcjioKKknmjpk8zoc4UghdGbdVNPC7cf6eW1O2GeMmwuuHIE5i+Ib83ftTo
dBUFcb/FZN51DtHI//o7C3rCi8JuadpntYUCED0JQRQmJmS9hnEVUPAXk+Zl+1BDj/WmcAaE/5XZ
dZ0iihtfQNBu4Ty1thMuRhpDo/JF5rMdLB1KauyHv3yvYkkhfDUNdwQOo+PDR4QNTWYZmRJw6GAa
zFeEQ4A6tG0rb2d5GWCOVRINHcL5NdgKFoMVGcAUFn7VqtHaiZltZ+opQu7/8MdR66Mz8iE6N6c8
qEjKEfOsUCdIWX3JBza/6BWqGUr1xlD4PG3lZv84tofHLaUbMeO7Xm3ddxXPOdYQgnMb9i6OtE31
epyetyKLIebun9zuxCoWNUF7tdzyhRgdxf6LrQnT5feSUJUIllRC2asPKoEgQcBRUoFcwmR2U3tb
eQRhrJ2eQJRYzwRv18AaP1ofLdjz9gdO1mquvMSHX/Eq00MNCDIYvYlP6WstKBHYSYouMbBpJz7y
ZKLOn5cNi1/QamEiMOpVAxoxCVHm7c03NBBSt1HOcYW6Vj06Y5P2D5c1P4vmwuPqwGrjL5tkC/Ye
kPGxZ0U2nnYZlSEqrfPPLSPXeOTzyXFESnIQgsiXcFu7VBTaV1L6iKdSMTiLWK4fBqY+dIJ4t1+O
DD+g6WkPwTvYxkxAMYROhTLc5edekNpbNajZ4cAwblXaYLWaHAri4vOEWkdT9OrD094XdEtY4FoE
h1p7BEVmTOYNl3ipZnb8xgqfK20LCek67inq/3Jhmf5TYnp91NYAOuta1UDphsijUZm96Om+cnW/
kQRf4eKWqbIreXiaIUcJGCqrw9MRBJR9LyDzQOQJVW5R9qxUV/dA0Z2YC380unUeiMwVYmWEw0MZ
fMiRKGTesisOao54EiPBkmsTcJq4vo8YyuvmOhzuvukQYRvbwtlwdOdQHCfEIun624mp/Kxk+fS6
EyxAddJf8U4p5lHOZY4T26/0fv+nIi/AkIvpPiXlAPHr68SAU4n0LIJmDCxyQ2blF2Dmw/xEW66K
wk+lMoVw/nvPodzl25sTpW+TMdirvhVYW5lifrR0xKHa5aiIjuhMsQmRXwMo0kKj30q/dEEE7VLq
Cp1iaAHbjEVU828Xkd6GaxzWTiGwAyXKZZ+cjWKxb0zdqRDpzS7rzZ5PgJoQxwmdQ74qAR0hsRBM
93MynMyar1swEERkMGqMF+KBpcGVGyZ9609OPntLdoyY0JIJGBFS+I8dDn5alI1zxAqGXm6pe/Yc
S4NQR3v7fMXa/T+EFDvb0LaBYPeRTSBjaH1N2vpxoxJG8n7SlDO8dn5criip1I2goOmzDzn7pIhB
/1XViMxMRNjxT6MlZk2cuBEU2IMYwLh6A/YtVgmXIXiV2HZ1JbTlroGemkqasgOKUn4A/vU/nSr1
VT6AcD6R3lzRH7VXTQxCLelFw5JEesj66wZAzHbSgCschchw4E/4zymcItgaxYHZ98859FsKeu0y
g0JvPAK1PnaGgmVoshB4IVyWGLGkWclI7RypaMoieqWcPokI1xzyAy+DkGCZx2Z/FxyX9XRQpTTz
uyxTUh1b4yDTXv73jAW3y3PISkMo0f5tiYy5cVOAojHEinShA/h+Q9xht5zaknaFEGEwqWOC8jeG
AQYDDW+6OWuf792TxiFwn5AKNNANEzanwfXDXDo2tcFrXMeGGUWzuwDLycEs3v3lJoX1nJZ+Wby2
XCGmWRloU55JBu/l5lVeBHMOs/pc6GqCLJa2ft7aFjymOEgnHIxKTEl4edlV1VeS+6i+5vjZN3X/
VUYTBERuJu2+eIz/0cBS1VRiKizvEHpHRtivHqM/gfzPnul/KC0fGUKvJFATGorm5QdvCAUCPvkg
FlOt+n8dkAQ80R31Uch4+3dFSz0bRlD7PcWL6ExmEL3z9qIrqlA2QgGnpo3foWnTn7ilYVpIHogO
Qjbzu2dG7tReKjLRW52rl0BnvIQjkBf13pE3AMJy7rn8fYmRf19qWeYMnQFIQUiDv6WbY1LCAtC3
D0069Xd7FuZ3LHHpc9bPgdRPCyyoLdGtN41jmXFpNuXl3h+mZTI6ONLggmP+nefWGnMPsI1/amDm
zEswPUstzlmPNlA23/2yFmoPjNCiCyQMHzCzgJiSpljKI00Il3+yQ1IGnU+sNbRnJo52NKB2y7VX
paOTvwNdcZXeo3cAI/cGDvfq8nnaL2ISlCBf4nZPzPDCdYA4ZQdsxvChj7DepjPOt2KabpL2JhhY
fLeD9MN84tb0Qi5gvjKuKUNMygS244qLUGRILq+8sU1ShaZCTzBwVnmtcobWxPzRf6WJbqTl9Gto
cOL5tOziRXB+URE4AzNCoDHJ1NS9zDvRuOaChqmG4+6A4M6XmNs/cCF1H9R11cCHM1Xx1FIlox1V
JiRuQtRx9xwa+z9ChBqN6NcreIeHM+0ceepaAteVzALAgCor7odix5WS1X72SiD7fU/q2DbkOYtU
VHobrwPG+SHc6aahQQV0syAi2J8iaBvCI7DW4JZhIderGv7u1/qBbtSjVIg4MWm/+DktBvPckQlC
RaWejlNrPhc4Eyq1SJLwPqiEuln8tTF6Z6lPTw8fFcqYrmiYloFoxWSMT2PuD0UkTq67w45q5utZ
2/qiBAmbkWGt+TMHJ6GlQd6zrLLsngynq1YbnpV9rUqM3UcVtEKkyZT/TXT37d628IMwwYIw0ohZ
HIgpBMfcfIofYifv9ExJas+y715OWmzf1n0JoMUALHc/e66JoVtsRJHKjE+dxKLci5oEtY5YONmN
st4tJNT2yxaDO+C4MLoM7YAHaWX4nt97kMdLPfWjDnoHzISFsG0BtCYNaMwcL/tq2avydXPpvO57
wurJo95P60iYaJT/Ti/oqiLOWrN/acK7aMqKouBaDltZFBLhkmOer7lDNztliJm7bbehj28WZM+V
1VNgCudukCa+v9kUTCy+dpiAwqvtLTpTsSRjnaJ+sFv5D85mwhVNZMP6bhurXlGv10BlQxEN2d3X
X6qghEvpXZ1ZrYNgEWAUJsgEYYsyIoa1qUtsIZUWsr0zv8zqcduCIaC6RhAWzt6ZtQi+3cmU0TBG
MCy5MEhpDaAN3JiZ/lR8lrqUCpXq3lslmgKQeGU94hd1Kl5vNesEFpLJQEFVIbpjUWwhtIbs09nH
lds/LAhsRVwhCdJSKgFLXVTOuNQmX8IA11qUaenAlpZDzWzx79YVHtVKTqAdWkVk+gENM8580Oli
DGh12geVD7welGdPa87UgIm6VypZ2o+MEPaKbLme/DXAbov5YJm/Kc1DtptN5Tjb8UCIMXeokSL+
goy/2kZBXnyHXI16DZOdZOy7eVdnSfCJxilGfanZPxs397iDwWNKCFLpm+Zycy7wbMd5ZTkMW2E4
QhDiNsAx6gUxptw/vChLcZIgXnNbclePEM1Eg1GpCz24cvo+gd4HMWup/SEvKROudybfHCU5wNTB
xDMm1eZ7j/uDQyYNlFClnJWpb+mdMYAFiWQlfUnK9Quu64jntrlL2oXejXt0cfG4jY6hbPrSmt9v
40vPhX9abfVt4ypPumMkzXK9Ab8KUHwRAt58SjCwtIubMdBrVQbdYzbfmoxRMnMm/u+O09qz24QA
FTrmSXbojps2Y6XlutxljlXKNtHoP3pf06ZRGu1pGxqD7V3oO7tClzgKZzh2bbrSVpB6CHLBPur9
lw+8Zo6BL/UvreBytW7FsxgqjjlFGTJ15A3ABuyOfzBkhZI60MZTKjo//mLBse3mGAImUwYKW51X
1hBZdLtWBjBlrdUhyqLWtZQouhrfQ6TnV0Fg+WH+rolEuPJqI2USPbK/VjwlB+eGo3wJVjEGwwfI
PF+suVP9FgAFMFslYfpsAXKSf5IhH5nIeum0pU7NfsAQ4O/tt5Ak0tl2rDW1kxwK/PwrvBaEheEt
ldECHbIzrMHZbysFc821fwrQhjlEbPgUdClcprqw55M/5w/ue2o9BlgaBa6z6XnM03vaQX8A9o4n
pleLJPBqcf9OFc/fQJ/1Gjy2Q/lHPxyGx30UIJ8YXkI6CP+p9CCaegLygX0Bflvy8KTPn6PASMcy
A9t8/qrJFG2ciq8FtcwUyXhDNoAlDX0cKB+4XZPr5+sx9R1C3eWjjnf6HN+9UANd575UCDUHPTZt
/686EWYYnPBqpg1HWRvl1W42DKRpBiRppFGfNOrQRZWBpxQEimqf54kbdsWGIjEjZtEN4lEQGLmI
c4xmDIkxMtJPc0Q7NOsE66OYKLcUH+uXkhDJsX5kLm0G/a4LEObJ7FNyBFStZgJ0KAtvEoXq4ms0
/4z/vDjMErLJMXp5V4+hS17r3QRWyy67gddKcQdLVjgtaFqN1rj+4gsjjCmvMOtkZpidXk3khMwn
2IXqrXHYAY7aow+jkDhcMYGaLxz8fRox0pvhPVsTgQMvHCUC8Lx1w08XX3eOkm3cF5dDpchpIwYS
dXqUeRAx54Knrneq3DdrwJ0fXbmBb8FaJJ2QjAJaz/GGSZMhRjdX4Urg1m21JHuGt6l2nTDkzccB
1dNmdXogIwuYSuKMLis33kOK0zH4yoFUqFtY9Is3q/HP6bOU1BYqZoO74mPD2hwlybAHOEWQlyu4
rjaJJVMIFiCxCxP1/AxHjQWDK6yMaFOsz9/Roej8HJhaA1VL/F0bFS3GX3RnLsx+EVa9Dwu+f5YR
xknrz85d7isf07DlrymFQX8Alv+kyPHVHt2heV5mEdrdkjOUquB8CAXHyNisGGvmtOdK+EAUI+q9
K+fjf7efvHawIZZZKqqH8YpUZTV6P7XdWJzniZLqdNauyiopv3WzCa+Q81b9Z3/uwm0OG/OV42pe
VqPTpUMEOWTGrbE2BOUKxRnHqYMXmn8e21fxxDns1pSD5igTeFZ42akHb1N4Ms1JOsviiG3jwOHF
yU6Zaf4p/MeAZFwBSbbstdJeD+AccJrS0C3OlIGcOPvTq25dxMetXg9UquuZu9zgvRCtukBFPxjW
UGE6elvdYlWVddCVJO2te3lUoYIZnMCqWj9ArtN6OubXYVXCC3AQFTVh2zJuXkbhGjin0GaWxuB1
himlNDVbS1Cdq2kMT3lsLDj9EJa/mI51nNPWopaBnT0O13/vKh1lcoLi7URwy++LvgRZoZkmmFqR
QoYqAX6AqwxseLFb9Uq8s21g+xH40Vhkl8f2ddLByVLtsLL3Sd6yBc10Ft+ZAoQOgG35y4phP8Ic
uIfpxawtvzKo9yQO4waauEc+1RwUDEk4wM83I7udb8yQb9W1uj/bcF5M+AGotnRq4fvKgIx2irHm
tqlHXDvSectAK7lVnTTseZFxC1EWsp1J8s2B/hshfZEyAmbMNxn+eBLToJnv41u8ud/7uM99ptpj
1p/w5k7WnEt1xdefWh/sobH+TkctIdb/XMhM9EaImq+R5FX7hI7NP5pEyHcdyuZfmEfK0xqQ51ep
maN6+6U7MX1sg3iD0WWrtgpnrpskGOJrjvgoHglns4xyir3mAmjSOsaSQ3aQOPiKGuhmNYfpr31W
2iLnalg24WC2XUn7UHs8cSNdrvShGQGtjMZ+4ZcTFkD2NRNxz/ZfmS/9vcOslK+MXr8KwPMxZ+OU
/at1Rs9m+aAiS97LbC6rqG61LhpuwKnHcHUSQwsXSXG4pOxXV23MBG+9bY+RGVBRrFcsv5mSYDnX
SHUrSeRbcvYK0wTtg5slZEsr6373DUEcU9rsE9kvs87eBYMQhcZgcF0RGN6wQEoFU9e632LmhY2i
BpqBBFP5pyNyfixmDxO7ZWUpjOPnhnszZc7dWYA/pZYm5F1dhskTCQx84X0T8yCm5hBqJr0pYAgY
zVSNJFg3TPs2jrzzEWXOHpuSdU2YPmahhjI70bryPZdGw3HFEggGHtIow55xrgjhHnY9ijLT/bWb
xLTNeqxgPVMHJ4f9N5B4oeZDlBsWU1u5N2Vf4rRphODKCPub3zYMCFS2f8rMZWwO8Hm0ltwvC288
EAlj72BR5zhalmo+Jp3UnTtNmaykVhisv+XvXOm5/YejIIJBle9sCX4/K7JvS3umQu1AyRki90ht
D7A/EDJzHjF/qvkgtxgxPYfPylS0Q1Lh7H+HV5QS3AIKyvt/fvYIwPFXzCLnh0IFlhU7QVfVxk+Z
cKLYHXhEs0cJJT7EL2qLJx/iCtU0ONlab0eQCitaf+sjZPCyteX47KTBedgrURuzMJRRr/lY62Jv
A+5S/OvNWrQVBTIVewxJMuwh6M9EpXOymx+Myz6boeuMIilLDN46UFlS8xccaInu+M5JVAc82/o2
ULKl5oC7WzTrpHp/U6q3eH8T1BAPexqJk/hk1s79J+dUhSZ8Ofh3qa5H5k9V9iiMb7kzqgRaMc92
/Y1Lx9nF8nfQN4DF8yg+X8YPh30KJNj1ZjyRmqbK0NMb2aC1r+b0yse3Quw9TOrUuJwZ2+d+oeOf
tTkZ5mqPE3ypG9aWOuBH+Kltpa7wi6gpWP2XIVf1z9lrcEvmYxrJdrxfD/e4f8jXHEE3zSGdqRv1
njp5bsMnEUnB9lVlFHjT9Dj/+i7DUJ4uILSkX2XoR9NUkSjmdF60G5f7ojUxxAnsCYJx83azdigD
9bHXz/Bai7PzlPHJrOwBiunyK0BcAkSUyvGVmQk98QlY5xPKrYIAMLk5EtPgwW+IYNVX66ttFKfV
+9Mk02n8gEU38exxaA/gjzum/ty5Hnfdr3l9jLB26JI3qQPLMfy0/PK+QL4TP9BMqynxA85pqecp
WlsWCFs2F6Rtq9v3pngdyYOEGbg3J8E0d6YIpNwo1kBgoBb7IHLKqO8cAzBABpyeechdDO+fPDsY
IpswGrTK2P/QElKEYPdlDvw/UAY89nrAazVdDUMZ7uPGkUgj4vTs9abW4EDRebbZxuq+GhmmVfcY
QokmSpV6c8fm8c1RU/oAzmSYIgXGfl7nD6fkm0RIpI3xTzUO283tqhSw+KRf20Sfh6Mpza8erfOQ
ukcLFMDzwp4kbT8QKg4oIPSjMDjNFmDqAgEhTtTIOk29ojj9XVkQKMeUhnEIV4JTnaLHGPzJFFiz
KqNzslNdn7to2r0yOw7QHYSITTlNo2uSIYdu/psW8muXjtdYRu2mzfaByMhrJhgQxlyFg5c+4/f9
wRGZZzUB4S6JCSeoX8opwek7luqMojciRtCTh+qea8WnNP9KW5V+8usy9xh9m3Z5uzN6f5+SmP8i
CTkHIqp9p7MnJawGYS1V30LQlPZOCT7D1P44W0jM7Ptkqq9B1qYWGTBiBA3S4r5L41LZ6GU7Z/WW
Mpim3r+j0itQiEA0vVPSKNjx7eR6SqEw/Rxzb9dwrSp8FrfmDR0vYskyX9/7ZhYjBbR9b8EHJ7Pa
1kJ8wTugxfIkMBBpOKeSvGm3wqIWh6k+SowZimpL2n5q4ifIQGx0DKcHtUt3AWYj8C6BkDIp0qXY
Wmt6z/kxCTnwnzSugQpGTskER8dWpcG6TFgmc9J8+9WMQPWmUWn0Ruroc1Hs5PKGLftklvZKFDQX
/+JyDRcfmDZFjYevnLMjumeF4GbJ9MaigK3XT+kZZWdmRycc2/csZKxaCH6/UZeqmK2p9N/4xfQ/
yRMUGn9pyUK5SOXglo6mGU0gLttfr+luRIihEJKLPMpu8yJ7/nSUM8B/FH0+AkqyOc0A7ZN1mvwM
BfxqbhS9QvYgmG4yrJyth4oZnczkVPdd6qkGx16sX54t8cvzTJnewlkFDfWh5GStwPfAeUPG4IOu
NMq5jmaaxbnQqD71gDH1J3Kse0Ml9i4KhNnt0t+EEQQQwNNf/hFrTr2BDREcUvDAprTbeZAEPAyo
kUheFZrtRleQD73KOaFKyo1edDasMj9eymdFyvwJt0VYnRjSbrdQb0EvLLnaBam7A6CSKlrC6Wbb
wCapSMTfdhPT6M57EQ3vJEE6DSaizpIwWFYapQBmqb1rCgFBSPOKpzcgd9kaQxxTpPiOmRa91pg7
43IhvFSRC2a+UgxC26XHfXvlKgFuz8lTM1ZYsE7A207SfHZmp+8/EJ/7ttR2olQw1l83hHg8hSTD
wVq3KtRsk80hhNuqAdW2dM9m6PpcdSg1iBKbQK2tJrCKOrAWYqNDRUdAAq99UQaper47uCpynqcg
86rziRsIA0lRqn2GJYtjN0GPAo/5jFJZwQCeBOef44Io0as0SBFIwA3CWVOzS1M2RGK3fAP/NhWj
fso7Z0PquBIzInSs+lLAv0KDx2FYqe5wSrraQvNprvvWu8u99IDeuuEC6dn967jGTvtsSnGGlgX0
oX+JosPcGIry9C9K0lXk5IOGbIyIYZmUWe51BubVMQ8aFe/QsOI1D3cbh80hizC7Tr6I7XaYygTF
K2DJltP3+JXTBBEDJlhOyZQ1aQ2qT+L7tynvgu06lHVOkXgsxrkT9PeM23+DgYZQ9FdZ8pVb7QjS
VVGnH7rl8TkEKBHEqQfQVcAjiyY3MBDXisXDhlS2DZ0ebRjew6fRnJY+E37AGwVl4+iT//T1R246
8mO4VMJLFrYc4ZZpGCy5FIY+hGb490zgusS6BTwPNTrbp1uJRzGq3WTtnTg8gF+vo7ZBeQwg9JZ1
eMadJzVuHHZ3o/epucKlKAaMM6C+ANWPDz+i4ldlPEa9bP6ylT4JOMPoAa3C8GUyCiPoi/ebsDOb
ombKvuElQmYfLU3MfjhRcegqm3/kLPUyI5Vk1U5bqkKqJtm00NT9A/h+k6DhVTMBW6t3uWzxocBW
OAQS6AhpRfjwI/vGZHTi03IvcAhnvX8mrozIP6L3u7P1I4ZWinghFHXRR4emdfW68e8qM9ibGKQ4
KL/oLVqk19DQJ13rR8Fegy7xZ2RY7qcmzpSwAAN0HBMNqRC7nxBDgnmw13axCssRIq2QoWRmoYJ3
yQw1YzSDLRKyVF0WBlcfLTVpQQxYYUOvYr7NVgnhn2Y0NcgrFtZurm14hlVIMWhJvmGE7vOva7zL
2v1tT8zOZSZlMH4nadrbffl4O1jjlUW0eX9njJy1VcREwpFXT6z86U7a3+iGH9hgqgFzxhh1T2Wx
++FDCy/4A7j8zlnYWGCa7zS1xN6GwPjl+ws18fBJ123oQvNKWRAx7cm9gQfzcNGEFMWkaAVMHgC0
0UoIXO/kNvQPSpX0903n4hlj3E4pm6Mt1fnRKFRX/xTVLpMIzFAIs+/8SDzPXGwGVhZM79XHYsVI
it9RVSrqgNWg0KIqVevLbNwDzACivoyo6M0A16+EfJSXX8sdVssezeyjnKA+bdrOMXgNSlj/aNvM
zgu0ky6FrWbseAI5XqnElOSMuKmjFiuNlCT1uVxNkriI/vBeQ0FdyK2C7dc26BTT8lo9KQmgn2ZB
c5hXH1n9m61Au+Y1ky6uORQfbkQjpHp1RR3OReDo7WJ5iYvuzBlkvXNIRQpXzBxkTjdmrWUehM18
iche27AJcjgCo3NQ6uWbO6K2sjRIkENvfgKdpodxaAY74P5X+hVcttLQhnSU7wCJlZ7gKQfFFoUx
zNNEZd2gD01xkol16fod53sdzJv2gnFGLJM+8uosmcjwv4tisJK2qdv8jSWWsDnU46fU/u5mEm3L
aCiVTqjjdSOGW0b0ZXFxWa65ccyLBFlN82hwjGvvbYjkeYIKIC01apnX01KITUA+253nBATjuR3y
ZazN9zAndpixGx5zqQZBxW2soP2cwe1WuCwPjpnRU3CzR23Qtaat6vGx/sBRiGaRC54qx1spvH+F
CXSdjiT0pVJYbEVwkayz/Nww06P8IssM5sby0mwjbijhTQ0RQrZgrBoJ2yaaK1t4qg2phlVdtUjQ
iiMxeJ9MCzGMF7g0VpAStFKuaJnL2ik1hoYDLP+7+xwBKeYzLSpUrah/lp4Yib5IJB84UffJ6AeT
f1Pi11ULex4jI5RmHTqFAv/qAt3jWZhZbkkYq5NaGpTqouuEnoh0bVGmnJIm6f8jhsgO77rQ6M4o
unermA64ViLQKYkmSAS8fSLzzeit5wWlq4Ikocfk3HchSv9MGoIVH62idz7RdQOEiY7szqlaqilO
kujhWWAytp+n3IqtgoBS/FeL0ssggYvtXGEWYY8szEd4u/LAUQjoZ48a9iC7m9/31svdlGUAjnWO
GYWXZ9XFYBXILD6ew4pGfFIj2mKvSnA6sAZAwjOr9qWPPok3ZxQqrPsk5S+fW4mSbKdBZW0934CU
w4W2Tu1+W5qI6ybsGycCkcSfMEhzSKkZ8sWLvxQOu2+EY9JbGUG3X1OHYe7haEGRd6mKWe22rIZk
wiNLxBaMMPSaGH3PXkVmQZFy3CbzDDO806LiXwaoQE2SBcqQ31lSksehvYJUc8/e36fOJD7hIGGQ
r2oWM6VWwMxEHFCDP4Fyr6GFvB5g/FVprMuXyKFpxV8Aw/VRBnCxl5jnzazfts6BuJEuZVahGv41
BhG3DapSZb3rgkcUUjmr5N/9oCaaC+h0xi8qFDcCV9h5F+6si7okVJYf5yMzBD4IOuLgLm74u1qt
dhQ1uiQ7NjpJ0k2g4phocHU45vVI3M7ZQb38XEp6xMdIIUK9/GEIT1XFwzSlxJcxfVZpfWWlFKzg
/5sdOvTEZ6u2YwoMB1Ydbvz9qbPPzsPRZfpVZsaR+yQk7MkZAc4uyIvTbVH4R39+oQr2Mbq5iryX
MHE4Vqd1smVurK5yd5jdgZMtugz2bMpRcOGQkbQY2wLz3BZG48EqdH74hPU2nNuIIzM8F1RgI0d1
87CfDtbOmDbHP3s3pcW8riEGDag5ye5N8ZVDHntoGwkAEewYb9BW3nRXiTJbHIpRCt0BkPW22L+L
MOisL9V7EwNr18pa/ZtYVBll663KEzg5NrrX/k4waxq9pkLl/enYdjwn7+7TcrA=
`protect end_protected
