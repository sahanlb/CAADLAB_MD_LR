// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
MDAf+1BySKoOGYp4+MMaLqRUWobCgp4xvcGlCkrsRj1r5LsWu/RgMi8JDSGV8AnR
hgjbNP8QdlQWXsyUrd+Kq4aapP1ukkwQetLzqiSNzUqYS1ZNavBY5TzgQ4zzt4gO
qgYIMOmKyfANyE3HPyw0b8kincYqJKHD11DYSJI7oFs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7728 )
`pragma protect data_block
J3oV9XS7a+qoW0dpUMnRYf+iHzz86yTjJ5xf/rc70vun2UTpDjh8h9YBJVDPAiWs
uRMLaKM3wgj7Dpk9jCYtenGy8i86X6m6aIdIsbUXbwoaXcYK/y/8rVPyWqAU7Wb4
Cx+5PfLpdmGCr0foA6DqkXPxr+mCa16sz+joyA6GRnSDyzJgMh2mAPoecH7V0aPE
jcOu2hdvdMk12XHhesOlQ4H28btsQqUI4l8LqMPgMQC3FlRuKmn6uznNAkoyyaAl
24GfY6gs/x/ziveS7vOnm/ns+pMVyJ5lYHUt3wsNumqtkGscmjmX+lfSc9JIQG1t
T3SMtQykM3TX6Q3mIrWL6higR1XXS+bmYee9x/jkmx8u/IxPMljBxxDHYCJU0aTO
Rp3xeUxrFEutYLLW7tGPoqo0bDXRHpykhLq8canWgUU0QO6fzn19qJ2lVXVfU/AF
8anqDfV1BzL/9fLZTZkd4EeNcypXQ4QkCzBLl/9nHHeMHzDbTau29chM3tEXTBkv
qknweHnNuG3ObfTk83eEoU+7aIu9ir/Nr8Iudc3U98uTVQSrzvoVVPndzsDTYPiT
rxRE6/hMeDL4n8tDhyLiAefSZaK49SJIBVb9qzb+Nr8lO6R/l085yKQdsn1+SMPC
u4UJAxNqrOcIKU5f2gPuljFI+ZUj6PMS/Ghs4y/CpxPbsKs4QyWMLBqvpkTtL6CS
DrnrWZOu97GrmgLoXIuqMtpEZSI12LAivPJjVXJhuICqWLBHgpPkSt+tILTPdwbP
b1A/T5bH5rhrtsdt8jBiW4OB4kEO5fTzIhKS+RgFiJPFHBS61h7JdNSfOnab1KnP
r6D83XKTI7YzS5GowHAphlGbX1Cv0D9IP6rk3E+sSB8shIoQq2vz0BL+QBe3uEhs
rWKc0bYFp8bgz0Y9GN7DYkJgakb1amgRj+bNrZ+hGkrJV3O+ad3Vs21eYaVvsi2X
FDLJgnZOS19GI6yzb7vlVjq4enD1dUKn06F8HvRTYBmPOVJ8LK1VDAYFvnpSeRAT
NLyWyLzHsJp+3gkPvvGEpShaa0nulQLVmBJxQqGwyjkE1D17HJgMUu+cbWsJIZ+B
4FdG44BHZMMZEBRxekT4890Eou/274ZxO1vTkGpQPexQUvTJGYJCo2vy0sjzu/AM
nNamjLJE1i5A8LE7RkO4ELYObXJSaEL91FpYb5SML6RQHsnmFIzuV9oS+SK3d/Zf
xxp99N62qJbn0XPeZmLL0zdntJYmmLabgwXLQzz9xsBMjT7mIdd5kgHHETqWpH3b
3o41yn4pP925MQ3El5/kqVTYRJ4+X/AD2HNOUrPR6wUOQj7uGtmZZ52V596d+Dxv
nyLU2dnQp9+skYWhn8C5vCVMmnDgc0hngnhbIzHr8udSxRSqCtmaUSM7x8NDXM6s
S+DYLAL+vDDEG5FwgH5Jczk1MeCnWIM/uAtC0GYfJW/6DnjwpVifamdcA3cNqnpg
+qiIGTV1F4KYUWKkPjdNN6UBtwaA/dojh/fEHtLHMxqeb/gIJOcJZsr3jW8aqa0w
0jkmhTVJUuivjvBLFZOrAvBdZ3VBqAU3NOvY9ZHqV0+qPrMlWEiISk6VUWLoTFhi
7vm73YaMhqqb+DKiCLZIkVIR6pFdppXQh7y2dNxBGrJBKx2nfwmOeckGYHBycVHu
KpHFrh12OHosqfUN3m7qwLgr9nmVKj5cHXCKisuYa9+RRK+3PrliktjDmVN/vXlS
CMB4nbfmQEztrfLSQKEwQ64psnJT9dxxYN1mJ0Qprv6WU3jMrfsb1YxzwYg2xlNj
CSRoRGeeV8u7a/MqLy3cbAC2lThpgJx74kyeuD+MavRyGbhhYkkzZ4IeVaQ395gI
0kwQQERvUFX0QvVrrWW6y/S201KNe426Amumwli9H5ZWU0N6GxuIoeodCp35DBWF
tIzLR44h2fII7Fs4W7J8rPbtx3jkZpyxWmqXRCWcGSLHATldBFY0b/LxM1urFCmn
+k3gIc32SdgSmc8Phmj6SurG+ph1Llc7k7NAJkmjUHw9W6metK+HLKyTZRysGXKd
INLeeA2CatuzuFOJGBS99t1DlFCI1tcuBmrXD2y85Mdc1OQ9G/KSoyUWwFmCSHQV
YZ/ZM6RFN+ysmSaQ7lfYxZcvhXZD3KDkLiqgRHPvlfq5Wh4urI37mBggkCFav3N1
beRKx3AIc6vuEvDuXSg1XEkmUP+NmbwjWoik+pFiHYY68yXdNIEfcPIDEpNkzdyC
Q7ed+8ToAc90C9+101tQ7beW2XbyG47hprwqo8H2L8exkOSTyyYLgosrRsVWsFwq
hQSvifZCwoe/IVcPTN/zAtASMgOiX7D7//MqND8X9VJTkuCKRn4ENHGVCLMGO26o
Sg1R9wOOJvOhtSaXQ5gbb6bC1Oa9YfQ/YUgXg3ijZTGrNF8rjpnhKnM8ekR01/ds
05lzVs3sKOgcbZdlgndL3PPeTDXhfF6jwASUuLWwc8TZpm81DV9KyKQRUQxADgCp
2kB63Ppn9F6QtKoicxYPFmf67ZxwgX7h2SLSG58UjQG06tHIa9B8FdYkzJA7QRcE
J/Kou7fK+8aIuaBWSsIlGi2d4fG+VdlP3WTw1IGAMwJL5qleYCAHaP0KzwT/1Zu4
zW+sGTot983lbk9T9Zgbu+6kUcQjiEY2ZnriEj4BthLWdPcHeGRmp3PfiZNFJSKW
sOR3meQMiT6mBSz/djGyHLPSOZUDQoAy1/G/76prY/0ODoX86Sx66SAzdX/r8+22
gIq8mzzb2TEzU121DEES0hmNjBXYpqUA9mvH4GzhhJ4HCmdiRge6I/ybQawgtOLe
E6fw55PAGJUrsf2MTNWbosxU+RsHT/4zbNICSTrwCuEAGVQdfXv6QOVpYwLVUzw+
Yr4CtaKzfWFUU1AL3/MdglBfUG0GjHzDnWMCYo/GXWBBo3H9qxqTpXrQlr6bIJ7t
M0EiM6uKiVgftUmHYFPhmPlbHcw/9pMXlvuCWV6OtmSO6/ZFvOiWjjcskn0JSEW8
G7OFlYtFpPq0ADyl8mSf2+mWTQwaW543grUQVXzhkE1aFelRMBHpPl8U/lnWZ8FR
t1RQT2xZjVy46GEwI8/5gDmnNPSWAlR/aQCGOdM+UmRnDNkiHMOMBWf5/TsVOfTK
MqRQKpC/kbE6WNKtnMNePbilaBONK+x7BANI05SGBVCRKVewggjacfwUNbIXmiuV
z4JELJcymgUUNyDwVl55EtZTkJ/B7zidGNzk9d2EksFs8yQ8Qt646DZIrN560iOT
SOOJ17/L2kXFnL5fMbEKSc6L232K+aLETYsoEIEngMkmTKkxWKaWDHnuiAfyFK0Q
O3pHQdyzQgWsjNJGeii5vVROK5jOJqbGuKlqjQ4fNaR9Hno6VhAWViVhbdS32B+L
H51Chryvqfy32whNWYP9WN9z8w9wcni3oaQb7rkYQq5mw62+S7K0BRoguK2hrg1i
+g/mh/GyEvpwvJPHkMkH/q0sIDhQZ3Af3zWGvy31EhfcDAKZtQw2f2E8aLSEDetj
gdk0oBgKQCAQlrUrZTKBzysncNPRgcV3oqlHP1eVYJWzTF7jPkrUM01eTBZYUy9R
l/fsLrcQTUr5BUzavVRwLyovroV0yOyCWjqdeVD9bqQEWoAMJhIJelySLEQQrhir
L2mnllruSRSjWCr6PeJyYj6uRltQao0sHbJbWXxBe6CC+DtFf+IsmzID1a1GJP+z
cSZn/2Ua99022Ne01dcPbPlwtbK02/Mtw3jEaKXwctVTzCyBplxXniEdvNrY0ByE
LK2/nk6Ffm9eoGYOGIIA4ArphSaa4kuH9BfeA6TBNz9l9qwGonkMxlY4V9EPcmCR
36aJKmYayxgLgmYM30Go1NWIEnq8afboBISN/IarrhmewCxIP8PLAHfKNb5V4GW4
PzgkWjWEGi6xO7QokhQIj+ceLS+mydL7JhHddxfiDLRLLO/Iz34Sy/BpeJqoNkM3
EI8iTy/P8KaxwO+PMWT8mHlB2hz+8t38r+Qe0AeNGtgbkwcmuLDvTzjqiLvx5N9t
+yucjvq5hM4K8R3ma5deKC+/7U9m87WCiqE0ghuZUu3xzK80rH5oqq4nl159UzHA
40W6JJ1sPvXWwWJiaE6eKWEscRuT9v3rAZ8ofpYBVrI4cxxdXsM4VZJcavufB+1A
wHncT6xm49waX/H4ohAoAggt8t5vpsE35teK38S5zYi8V3+OSLjD+gX/NlGViVuD
bmGXJkZi9kYOBKp4pq88DJ0VvLcvBcWQPFi4LRryYmNj8Zf6jeS35hEdH6CLg4FT
IPnn743ZHMh4rTn0WyyP0xq40jY9R/FdBRrcY+fJaPZ6MtkIWwdCTBK0UbnoFTtx
FyQfineesKBJJneiX8fJm7WymTwTXPGl0LCUtE4mbhaDZVSotiKb5PudhtnNvEOF
H9SUJSMdUPFNL6rd1xWxScbdcLXWSQ/1Hy1c8WGvbxJx7+91mSZt6126cnvdaIvf
rQ1GUfUS+bD9XTY1WwQgSDSgnupg7tJyMWXorlnxwww3khfj/b1jDZWzZviHJtFK
nPpwnJOZ0YLP/XR1maxiKsbYb6NRcFL5hhpz1+mhb/uIFjYXSDHoEtN+zgzwsji1
LE3Oc/Xdl19rSMedDejCXMcEuK8yFrjCYBZsS5xKpkXLtLwIX5zkSMQxA4wrlc35
Btt/VfuvwtRE/8nYjuruPYbA8yQ9UvishadFia2FNwUBzHwA02j/N6ZCHygNbcYR
4/ZB6pmhHpAdDywJkXaBp13fPly0X5a4CC2Szmknf6KGP5w471JF8ZGCV2xf1UDW
a1a6Jdmpeg97IyBuBUtmU3lPydrSt4VivIbXbqYYrzGiWYvGAwR7LUbGu7cNoStK
xg1ltw4yR5X0rv+mK+rzFD2mNWUQHwFG9iAR1pIEVAYTKX90WA9k16isI+kAA+v0
DOP1fak0w0g5J8fekIXcwdwZnQtQPz0RC7f7I3gD/nej991VP2NDaJJ0KkSNmo/U
PsOeSkGM1WJahJLqvzZm/oQj+ZDTDpHYBfFdzTpJ8G7TaMJg0N8eR6fM/cjxjeqR
5fZWrukcLlCFyPUKrToC/XvCWfjakP2BOt7NnT52PTVEvgXBkhJ5ETDVAe80FEDt
uSNCF1cP92+/07hsdRUKwqBf/6xcXFLnH7fpE4DyUUokkDR+uMk4ryPQrgjPT3pw
I5plAW522x7TQJ0JRFZp6Q1UV7BGVog1jX9PSR6xY2GrektE8HtvyaxOBDHUqoeK
6nq0CnDvg3soxxpVzGyhCDp4lt2D7nAKlYINIur3yZMLyYPsCYsdSn7B8VuolczX
PB3rNfhqxnAMw5TnZgDNKGd36deLTwzWtpUnC13NRuSvW7r0xW8yzPuQ6ZWC8OBA
fV7Zq6B8SnXVXJkW9afH3gzx15rQA0Vl3wRpIZuX8GqnpaR8sQ44gUukjop9lmDw
vt48DTFAK+PL90FCnOYLNa6EnDxZ5PGl0KXjuSvZuImBaoEbEPdpUtBt3k3zMar4
hQhO+oABLZypWDaVsq7V6eJLqqp7TImUZ80/bx2OJpJUUIONf5TJdH4Uzw7U6xeq
bmCspkc2Q9eu+WIBLnxwydqoEeXQhE/7tY1HQOO/E0KiX6bcT1zhkk1rquMdYkrr
MPMY7JAk9S31fvv2A6Bhw0cq5TkJf57MRkk3Cnu1PaaPxOFWq7yJ1TgbyRoDrAi6
M9MoKbnVJuM+LzzrFA1t90YT4uk2U2NobL4t1yUW6OJ18QAdItkhaGiaaJ4cRGlJ
zn/DTD7OFl+5cjrU42m8x0PTduN5WGhvvfPmoscdGKQPifaOC/HvQgJ8rP4VoV1G
PyDWcD44+jfm/k/qUA081PpOsL5q61nQgyYpO1+vora4D+kiKDb0TaFNMou1ipQO
6ctY8yOGqT4dg/XFRiekuLhGHtzZ4Fwa28HvTvLYoClJa+/UTk+KK7Os5w/3nXye
6F9qC4vGoCuJbhHXSn4ESkDnrCbwKHHvEktI5WyL1Tqu/nS89SFnOrgsf8vLZXCd
RwFHSbENe2+Z09uKSjiIfO95dGaxEXLLhgs9hH+fc4AhQAGtosgGu8lVTRM3Eyz2
cCgzg4k5A438b6AgQAZpwTEv+8oNvo9cqkaYo0+RTWnbKOGtC9kNMf5qVFYlUUdm
FO9vSm1FuGX25iBcSnaIU/tR7BjeJt2dilDAlODNrdwRR2y2M/QHeyikpqB3DHI0
qnYHH4d5lQC02Pa9dSD/LMCiFJARYYiMhqt/PiLic0XqCpPHXlsztkAG602LGa1I
bQt8ue9ikfGZiXzD0RO+pqucZV8YD74E6uGvwSCzWyqUhi6HemCoIvDT6oM4t2ZJ
TTfRnlI8bNqxEIorarzc9JavBSky2ro47ecJ0mk8jTylhqfoR7/xGO8wIWGxVhYf
WGJO68WU8dSWbIGEEhckGoQmY/NxhpnLztriuQ4PbpltM3Jab8yg+tkhGoqF1MoK
NVQuLXZGm5yEhVGYfhf0AGNs/51D9eb4Zcu4vmP89Bv1Ol1VRjefUc/IQB+MLGiE
kLtEf3cMKgeFLwS1X2OqeZFvuaPGBI+opM/CmIBqXGzrf3BdCID/2lJ0VMpv+h+8
Y6mxYcto1pNypuX4ZJ/x0YvXKvnQk+2XDYvOqLNJ/sjsAUcQ3iw4wKdKluljsh0e
6FK6IcyYqbO74ogJ0LGNqWuLvgY8EtgSmGWa35bJAtf5+gl0nXTJb+aqsIMeEQ8I
wB9rgU4YAEIsOvtub2uIiUt9T3Ppx8EO9ESdZ/G/Hj/JFrEITBgI8RbKXCaG0lJR
ialo1efHfhPYKZtbiXkrhsTChmww6QKGflU0L0NnQl/Tubfp5olh670Or7mQ9jUr
fJ5grwAiAnvsPmJg//Lvj/8MlBxITj4O2Xg3wq9JYAkUwtIo6TmEjMcpIjTfN/xg
rfIXe5gCcUHOzT4BaNtEYeRB0bcxV7U+ZNguD4YlgWLC+Smk+kBqk3GdDOwrV6sh
0SgUowyDKMg/DqYbSkSSLOd9Cqmg69mZKEv3a70Wbu2IrE+R/pOfaCKG0VxkCr39
RCG8qpuB9It1ikPMHlsvqkK5cnSN6xA5Z5Uplr9U4kHikurh4/p7cur+guXCScRS
+7jE8IJ7Ymghe93a+kBPP+5gYAC9lEn1OdUNUoxbPaus0M5QuHz5/BFWbxMSp6kE
nuCsKaIr4sREkXj+Txhv5r9NwDLvHb0eLqI68OZNVg3A07xHZS8q//VNhOjgRtU2
CqSDo4+NW7yS3eab1A8HWck1zTCnJr9TuxqLSbhK/TA2edrflhMMKBwiWezrnhK9
bKFjfYR3PM5CAnhU9aosuxsICcTaMai53cAjwIShkP2AQChj77VZGDsx4uXTWgcY
sTalhdyED8EiZ0j2S3cpCGgbGVdUgUX3TPQM/TieAtZe5MfovYlBpmaXJMMXbR4j
GMX7q7bGwLyrep2AYoXcJmsQuziqgPC0HpanjNwYEVYg6O4vRXi3OEtLyLjRUoXx
P9NVfoRA9gXdGXaizWonAZ3YTCZfMDbUQXT921/bicZICMxOomZN1bOkMa6VlkaA
1MPN3v4lerHmbO60Ce4+bt9YL4RJOEb6L63uHZJ1JdV8H0x/kbP7UZY5n6uEw0L3
UG755BcZRoZb1Y6FQb9OEMctV8OmkEFLEWuqJXCe9qOhlIhKdaW+Mk/S+XzN5vun
c47Yb54gzBEc4n8DXZmNoRUSvOpUgH8uZFSLggBTzOxzYTfZIvXXflYa7RDaJjN7
dAGZeoHo4miWIcPjzyuIB+Lb59dbXqfck3S53E9N61zsj35pW55Xk210k1wdLqGq
GtDNQ6WJXHotOHSg5CqFdROFt/WxUhrbRmwnqxfFw+eLNowsTbCoOskLwleHewy7
BagHpJODGoXTgtOvPdydbGNvti8HYdMRRaRS2oDXPrU0/TJC+0v8GDy1caF/pg6M
N/4q4e2l1Dl5hAQU6GrxIBEGOOe9X4b1XmTvrMW9Synbl0QCs5mQCuLneGZ0uxmN
uaNaaHiJIAZWvNzFhQ2cwmwBTLyBT0d/QFLVDLWaApQydRaE100F8f8PHIdsymXF
r26Lc2AzCpL7dyvMt0JsbOAk6sozQVkmynZN4SvCKwuMPOySln2bkbRWZ7nfD45K
8u3FprjrNJRw6BEXXvnd26aXEGa0GCXpeBiR0uxjFxh0g2xn3KvarZrE/GK4DC+J
YLQbNkHU88Hb9BShxrp0r3zMgAPsswmqK/qriCfZ/ivAYUsayKN6xZxDdsq1FKG0
D0IE9v5Kv6Y+5Ax/NVkpv9lOvucn59pBt3UnEAPBmAadUYdmQOrwk6oXQbdJrh5o
4Pn4fIVqKQDdJw3zrxMYplY6L1eryWGSHGcrA5RZuDYVWgeGBHDgP57w3UwIOzsZ
yJdfTuBisExJkQOxWMFPpZxP85q3t+MvZvgYj9gqeZLbRBGqMLhpeqUuMnDy/zcC
Lblcmtx+KuIKncLh/DXOdNkZNQ+BSS8adofFpRa++Mi0wt1VBIRvmJKbUGGcwk6c
iGNuC3AFn2qCGiZaTgM637upqm0U8xIEwmyU26aM2VAVhHEMc59fnSD2CSrtTEQv
2qIJaterdYyXZ0Ba23RymgHUq+SlalDaJiPOlkLF8zLS8ZoIEdYZStVomidfUwt8
vxA3/jtrAd9j9vNP8OQ30pIaueYUYVs/Qy5wqAgXCTBqj1coPIoBStF4wZEiOPor
eBBmdcz2HZz9NOSaUHZhD6bhxg4CvlmPblVx+d8tQXtFUiChkLz/PZMKspv4mPZX
0ZcG14AyQi/FNFfPFCTk12BaIlhnMZhSsr001+I1/CF8TvC2zixg1CNGa/jeEoMx
lZDyr9uvFpcIByHYn1j7TTLlms0IWlny5w2Gd706yjtGTKEoS4/0xY62MQ1mVIxZ
zgIjoaYn9JNk2duDvLh+Cj3MbFIQWal6Q61Qm5aMXgvqKnSJmpT/PoFjwkZh+kGy
NF8r/pG9G+FT0vCnpO2ZtU8CGVDZmbCye2w5CXX5njwKdnREcIdiRYMnEAHFqyV5
GF6JH0VBDjDvmQuAbHDH69oeF49RNpS4743PDFh55LRoroUZwCeRoGjsbbuqaplG
GE2skYMYE4baSQ7JpFzyIIGiCUXCda0yY8gcwuDzwWLu8LY4UZgyUZV/sj8QMeB/
wRpw0QKzDE0L9oME/lgeeVcW+AxNTy0OjuSem3b+q3v+87O4tsWjvBqOQqLU9WZ7
ONWVnB7PnjAHu+GntyUrd8m/HXD9IQcdSb7LOZHbtQxd7tm3J1k4alsq2/rj+gwJ
8yeuivmjWeI+0u8qAzzB4yPG/DMCNHqfcW2cNAxJGBxeE+W6gVVEnKBMUvyjhnST
Keb/PpE1zYKvWHbcqoCOJiwknEuTxmIZdyJ/VrsjX17h8tQ1heRp4TW/06kD2kuk
7fSoXBLdd3pB4teayGsp+HaJaAHzNKAzqSsEiM9tztgDc4G5SRn89rYiIBDZeO9K
n3f+ftiCtbktjW9Lb0MJX902VvjVT9uzLJ0zQIRLwpZFC4qm9nAWiZ9vA9U5yn0o
EDx3cm+r5fpud5tP79TTCNJrbk08uwQ0BxCRkv4vqymfJTiBzIWXJQddOdVgf25L
Gy6lVbw8ulcxvxup10dun6J9rQrM3CEtI8gNUjvBDZQt0GlHBJ3W+hr0DZu6nHfC
6tcnPK01KpArfVtY7nv1CHHv2/UhfHVrpl4EPOadAuK/9FfFsbSkvbgxlD3uDrX9
LOqNUMYY5tCh7jNfpMdL8TL1JmyfjVQh8JvgxIi3Qg+PdRwZnNjXVgvh0p537DMp
MziXhv5jtnU/j/9FE+IHjgL4oEnAyzU6LNKNu5Mi2tQ/w/QPWQZrPIzXjxErqTvj
TyxTnE3j+jXeE3bDnrplWOGy93kd8h4gny0Emy02c4S+DrtTHxRqMNGSLaAvrw8Z
kufPw9kW5aviWrpYx2JYTNRhsaC2S4Ik7fbhe1/mg2P39fwePs47b2a9pbtkLD4j
XZsmg0uoWEHXQr9ovGl986QGAfkIRBhPBKsS+aktiyglkao3q8ReUIRCELmM2UOJ
upKnA/Iua9fdhXTSjw2Q+jypGaEpxuJct5PAOu53qQ/iUcd6bwYwtq///+UxWkHC
dhGwbh2b/9aJD4U+noBy1Hy2iTV/wpv+HHgxjj1eMhC14NTkscq2WG4J/m3QarNx
OwY4L8Oo+EEQkYxONFvb9W4fGaWLP3KDex0SOSWpqY0/pqzkDiiAkDQ4vl29tPKq
aebykpUImIod+aAsqRG3m0Hz/SPLD0o+gAMBEcp/qO7wltuWnGJsfawin8c8gf2/

`pragma protect end_protected
