-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
fhVqtt/ZPVgXJ7nu9+Ge1+XVMFMb6mR3ysv7KfNQKDS+PcL368LuJYz5wSeoWmOA
mew8wNCDVzBaXIsjAQZW68cnjkMFMkiLGkoF4F6ZhnlEofMJbRVB9bjn4p9CEJxO
s47a3sT6xACEG91dcGDJzYXBD6oHmgDjopql4aLngqw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 4160)
`protect data_block
ehSX6gpaBEAvW+Pxe9xARhJuQshPouBqQ5/BnF/9NNYlXeZkdrK24bs0Mmt0ouAZ
OLuKKgPR2o3gZmQP4zvMeKbKhFAxUPxgE8BwytmyyBbjMtTdhs513L8UoAIN9pjE
TsV+WevsRteOwuyYe4hga0Sb0hD7uLOPsvRygBdljQu3yEUjXNkqn066FN56fZF/
kAlK7sY4hOdTuDOkS8SDPjBZNRPji6dXMzACDeIUYotfbr4pROziZYTuRnqtCY5Z
hVEeqph5sdmGZx8jsPh7ksQv4CJNOlrEOPiuretrTpwC6yHgzuzHLmk6Qqy+mG7n
Op3MiMeRGATVYMfswkEOqxdpd1Ds6YgULzh3iQj5PPdfp15nM8p9WuWiJnFZNuBu
B3G4ouVxCoQ9muOMBLEjHZnY+dXXQ/SM5cphC48BOZu4yMlWT7PUh3tMiRCgmUlR
mekZJxWKhMdZ1Qy2IkBEmzDkQC/rkq9MXHMKvwB5w45c9kmIIAn//fOYcRnUPgfF
2WqQpe2jA2TjzSdGMQ5QG+wg99zLJrJEqVl5Gj7epXCop1CknqiU0vo+vTX4IIC2
4BP1UANwzX0POF77P5Lk8CC++KeXYEwZik/Jv7YPYyZ+3a1gNX7zgDm5aoGqe6UL
0DZETa0OxU6nc2skRvogBfiAdbrQl7HBWvlI7lNQ2oy/ar/FO6suVL5+1Mml5X3w
elORQU2UkIoH3TxPIlfzRX4t7RYXDg060n2NJ6YXbsbRk0wLPHy0JVaGuK6gpdYR
BhdF3CZD7d7IZOmEZ9WGGsc93/banRypZl5l2F7LzFT8dhfe8BPvaJpX5yUb2EoC
jnjq/1GzVeOq2UpG3/FFwyKE5dNxNGJcQfqxsKqbQIopx3G3qy3JTCv1WKJoTvw/
ac7cuNFR17leza31u1VkxK58wIEQT5aU0R5lM1cAkQ4Xlfns5r2UcSdl1FJRju2o
/huSQ1C4O2xaySdSGWQpaRQoFz38rFYuV30kz0fCzutw4C7gIxRn7E+DW0sZ5mJI
V5wTKrNyl8kItnXuZkrGOsX+645sMcqRdxslHJo7JWKxLtQR+o6cbqqptDQhf3nR
+027z7iu870nCFhl4UghU3q26C6VKHlypkXr/G4zDUfEYwCUcQtN2c5fVvHdQ+WG
n34dzc1FcAt03qRnoRTsI9Up3K+ToF3R21pINn1vaRoODnJUKZT46++SZXUn5HxU
j5B4EqMlN1qRUsxB7IM1pdhEopF7WLlt/4SDTxpMktz9MuM2+3uYrMwGCHXs1Guk
RNw/lH1LohfvH21qh9wLvwuoK9TOe8V6Nnev+zXpX227pM1Wcztje4au8+9yDgUS
bpLn6PiE/R97X/MDKhuYLK9jchnuLTtug0JyGAw4Jsm+hw27tAYq2J4DSmiKqdAC
G50HD2x/Nse2OBP+7V2EyBOwyyK8AXvNGQrdF0oy7rmYgkepd/GtbtzlUGi/hFXM
oYhk4U+VY6rEgyinKG1iC4sFb6Ass+K8E9uiGcphDGJWt2IAiLzc/+UPyHisonrO
TDRef1GIs2GUZ13QyJAj9hRS8JgBeuxTPCBBQE2PAxICznFLcNLIRKLwFRfSmNrt
9Cy1rioqFItwnMfhp6pjlmOMCcZkazYaFt8FJ61meWg12Z2SGiOC/SoVAUZDJFBl
g3qi8Dsjitd/txjoCvyXwnekV6jYCqZxhf6e82hV0z48n82d/1U/gD7WIbTnnlt/
lKiBQcX+Etayp5UcvvmM3En1GGhpgoX9xjN0FG8kiMhaMreDgCp5iYomQkAq7ut1
KbyfGCwnga4MLR9BTjDN64KQ+EprtQ2qNHGtV/l4pOOhTKoUgYCtFLedugNRSYqQ
HJZODlKeTBY95MEfiXnO9t6f00Aat6o+DOUCS92tQBOZAGIUtgqclyIbZ57p9NlG
aa54MHT1nULqXCJ3VrNP11Vppi0S+V+sncww2XmccdQcg1CuFFo2+edg9AsHd4ZK
Pqm/W5En4/sGoTh0QPcfzLszJkcUWOdxnZJbfQ7sTomNOXmX8KwCxrzdMmkGYnev
ZKF55ikQyp6RZTZadrE3iDOLsiJOLP+AX9U287t6MwRYw6KZPqUHL5fqLpdBkaVc
X2fzONY+WOAHlRHkvGSmLOTmFmGd59Jo4j2A5v3ZYMVS1MqHfqEtePgS0EiRcCfQ
yB0Vu0FqDOva2T5Yrwg3ak7fl9oDN1eJHS+PdaPu2jhMKSl4DCGBgG/+b2Tra0MU
qYUMTiVuZ1I0s6lmKmo53mVmMUudY2+0WYNIx9bYhjjjYjkokeeMMpXHOsKtncRm
+CkqGTdCNu4sp+sQK6ViBuDOyWJRMohZ+4oOZQc9kRsZSGVE+PqtCWVFSPPmI+LV
a1vNxfm4bkhgsFgaDicV4oTrTgM7RanQ657h26xEiteWaQdhD3WbgapepMapGEV+
Qc++GvtcC4G3keM5SN/B65oid6cs0zsOAsKyT4oHWuyxUI+3Kq3iHhyGosiBcbFx
oloq4mkcZQlOaXrfcdGuwPEJY5XRLUYLmQwnQjGHhmhn6Ygx/qcx9IxV4ImHaqUV
9cDQ1hdvAZ1/xJ6kVeix/iLUVOI32R/+URgtcZ+yMUxnP9hRlACOCnM8n/PXXHoR
+RxtpOtjr2bE3QIyqxawPVxVc8zQuXYwgJoO4qLwZbNsf8YitssmshaYRLvixjar
8OJfTMI9Y/2QYkpbkd24XFnTOOOwFWkwQYKPPt+sWFSN90uniFbaQym6OQYbY5F9
rPqGKYP+xAq8kvEC8hqGK/cgzoko4nd/lBpirDlblnfoq2sDS6jqD+N4ilan6fNh
nFR+hRvk/PLmt90wyocZllFTDTyWJSOROgF0pSJKQPG15SkJ6abqpvMAx59TWt/C
TzEaGPQi2VrOpUcyzA6u9IREtZDKTLcgCqK6AKLX1cKuqwQwB/WtRMUtUvSRBVsk
Tlqtuuu7FVLhogh3M1JG2H1MCK8bgPamLtumsnDObf/4e+00NizjZwH5o7Vho0Sr
vUKQ1rzLVWQV0U22Pzy7Cmf/dQXFomR4vNUoK0b0C9WbNECan4B4QhodYky2v64S
mcK88WN+4JoF+x2lW91j/So2BRNopB8wLCZUBDEGBoUTLeiuW2LfR6d5drNzLD+8
W7/FR8hDRmOJGqQH5dNaTwHjIxhsUklgvjGiRfrQWxZNTVOY83QjQgMuzWjsoSP9
eNeT/iK3Ur+jfWuiF9qL4V3bWOiKBg7B818JsIURz2iRuumlMeTNGk1RI2Lvaj4N
yXiK2inhWKu5/lC0lEQ4JmsjxKwoFKWwjrAAx+9j1Ayl3oyhpPKfVlW6uK0OcLt2
b+iTznNlFuHwElMNwBCKHzhDtbmDRU5DUZ2d2Tryi66xuzkkHp2ftQFsYvTb0NSx
/5oNsTsQ+Ya0mTvfbM6Ru4/6fQ81hMg7JYLfIGnae9VImEGUQV5K2tzV8IEjZc4U
EAS6nljr2TEmJ2AIFxz3/RIBngM40vxfYhNb9OxEP2XWjmo7ZiOGbJy5vr6qcCBY
NSRlukgmBI1lvJLcqWpqnnhCtAzZ/F4XeGd2jS9lXSjHi1An4/8CyBadiA/ewgpF
ZWSt6Q0YCQSXdu7xYoWlgbSR6Oyrm6nXMcIejZqrAYOtPcz9lHr0fbc4S6+dW5oO
Xoecslab5tTb0l8xQIQNKFXe5q4yciZOgEez/fiNIdFuXvVZOANwAEiMSg4yzrCN
2ftWKjrnm6lqmWVzsuj9YmGF9ftHAV8dIrexgjAn3RRb/NnQfhbabSJ3iXEQ/yyD
APepI32CCEKJnGkwynjH/Nyh91C9i6S6/BaW6EUO5WAPV90JJKU2j2+/jGbCpuoo
q/9ZL0Xit6wvySRH+HsC2z2982144eFZNJYA2+VDtgPK29ou7XHzzTN58QyZFDVF
gyin2NbHZwS34jEWlFfKVbYuO1ujmWC6IafGFNHq/+7qfM7qYmIBlaCTTvh00xS9
iqdhmG2RmkEqcVpgwqXK3jQccX2z2mwIaMVZLhUfdW9bI/DZSGWu+yAHO/CFgzrS
gSzS0mGhfg1Fu0jH0duQhgXVKhWUAuMiPdSJpBP3YuBVkm4Ff9pZO/1n5dOXcQN3
53KM1vxXnv4WrQjd1J2Mg36T0N+XA3DR7qYpAzfeIBgyfbPyNId80UWcRfRu1Zld
awyNtaQLiVKFZ6GEB2m2Ck2lEpAfYaqLx/+9bp2E874Y6P9amwo1Hjx4b3Cw0ARy
dwMVSYPx+sglfZ6bmj/pUJ9Zypco98PjpEJ1ZSmhg99/yaxyQy01ZIdwsIgOTbYF
0xNxiJhcM+LpunFMvsSrDJKIuyBEoJiL9m5V2eqCLeNHFBcCyvVkgSbCArkYgbpD
RqySkKpSnSkgSeOFAqEMXcAt7bdwtAxmtdCf081XyFAyt/hJzuWdijIizDu3ddpL
mlYJzLjRU/YgFxvouLc4nx9uft3LxYJZ32i3rkbsPsQwR5PzEISTTWk978IwBclJ
ZjsV2uicyU1hRq8MSR8R8mdJdWSUD/89AohcDA6OprTqlMnUK43rEcrts10Jk3fC
x7d2C0BYZsWjo7MVAnLNGL1/+BsPICbe0oAuL6ww+h6LSLXBo9F1sX6QWhydJStj
0k8jjepp+xvYRYMPQduDqjZ4vt39waumimqAifdbvWsoJZtHxzkhWlarebAI+gf+
gC5yAoujd9GpT8AqLhqVN32/dmXRag3tGFh9kmPK1zMwJenkp0eFy+x2PkTfLQy1
HgFJ2d2Xtg/4CrA4KLjyJzDk5uZ4W8LNa0BE8Bw/OuV8sVORYDxbgtIlphGxnQNo
on6mhNh9RfK2SWjTN3u1Fl0lb4VNuRlJQ+TV/krM2pCBb6qNap3+39POa8xYQScy
e6qiMa+w6/rSCk1hNCjyCM6BQJH6iR5M0Rm0G+g9AiKUD3ZsG6lzdkunF/fHksrC
hEGcSnHDIcd2It+lW37EU/w3uP89+mluj2RgauNM/6/DqqYRmaPMpQkHyf0lx0hu
n1nZ4nu2ZrXl/UTewr2mceuV8CEdxNiU1VJkzgViPx9Qi8Qo6pT6HlIp4Nv0fsoV
eBUBsZkMIS0c2gLQsaG3D093bQBVEmgKDQCysR+ljR/DujqutE2mLbiyzODCOH0O
ox4dNyIvrZ66BkdooMoEbhuy8CWhFgh8YnJusEOgG2s8jyz5uaXonQl0WKV45VPU
GoVGYlpae0JUw385o6FPNSiYQaKh/7mHCtZtFSmSAZ1d8zB8AXS+cCBSJO34oqab
32HHg3QHBG8AIj72plwK4AwiJSfkvyYVmdEYnlzxT2+bcF9eFLVhC2Ok3gTBbIz1
EFK/VQaPKNkL8Eg5/TjIShDqGhaOZP4PZTi5EdNcDx6hEamO12S3RMlXbceuHJLL
SsiH9ND6RYdNooD+efsQ06Wh8Lz56dqhEauQNcTHkpDg7KnJPkngH8wJ63owG0Ph
rSxnvxuZWWxbtsaxEYwwXGHq3M3U8trC1LoDoU22HHAatWB+Kelo2s4zXwY9+duz
SZciqJrNmdg4ljna6JxqSV/+peeodpu5vNhQD+Si/qU=
`protect end_protected
