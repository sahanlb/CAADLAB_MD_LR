-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
azeLv9IvUpD2oETL9egITEdaHEQYCakVZEpAI+RATVnENo5BCDapvEbuDWqy7rxcitPS15n8CWAo
HYTLRgWCetJg6A1ozZmC0Tc343a7zM+Yoj829tPPNNz7e6EnQCWQ2m34FN1ui56hxWP0fa5jXWzQ
x5LwcmjV5So2fMmZTtuzJEpUZDDYvBxN5FX8EIANuhnRSaaHDvE/F+NYc8+nxJt226VP6hefeUu/
wJNgcHCbrXrXa7mxqmF0oUiwaW5l33FR1CxC90YGWQrvq38pe0CdXM6VKn71KI4CcmDzI7tsKvAb
Be5qmi4FnuguOU2k8+LAFkatdJ6TlhXlbwG3fg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17136)
`protect data_block
QOb1B30nYhVk2CJOTeyeNmByfxHm0kbC0JbylBwT+SAgi6oYWwNo9WLmF5lwYprPuJ1j1Dh/W2yp
P0adqWMq3vAj8yv0nyHzh/P8al7jQ4Ho8k8htZj27I2uzqW6uBzWZHOPJhoOlkVIJlVdtckGAj8U
2Ui2D5pgue5q1fTkZ/X5NpZINTkukHKksSeLk4WRViJVbzmREkv/F6kXn0GxzP4FkakLcu0fl3XI
9F6gI7J/tqI4etdyIcSaYfjof0oEZU1k1TQjbHGAXYI+w6CYjmqIy5S9o66I4oRKbYE4CoCV7TEK
Puo8TglZNUf/rlXJzWl+93RlcLgKfrnoSoi2n5rn86y2OrWBVrXT/imtXIozIiUZGeqQBm0t5r0U
nSWimo/y7IAVyUbwacJhdA8m27DFBXrdj5UJl6uJhrLmRQr+tq3IKlFlcOTRuXkDUfo4gq33xaBd
l59sLziFFjk9TE1L2hlIxQvJgoAvWp5T9UsEzYaBgop3441RQeDDfdtjar5LnaykSNEUyex89pLS
FPF3hogSjRHqIwx3Fj22AQiyXq/GlKaEI3PUHV1Iejq/XY6F9q0D7ATMw0oDm4Ghmrk6Vq4KL7/k
yQnQrm0x3Kpj2vAgs3GbY+RjigKhUCIHAQkm0AW17cbuSXQUWb7JC8733dyT9q5nwd5GXEK6mVC3
1EiznNCr9q4depEkRNZBfe59At+ChZ5XmnzumRbgPbzyNGbJ8KohqeK9ImnA2TwFEVzJB06hoJKa
CP9xO4HwUFPjP1EqAr/IYXZ+h4F8NeDb01EAuL88d2kok12K/6J0iilK96IKo9Mv76//4vj9I0rV
8Vk7YJmkb+GyR6SUrjBlMB6qM+kKm9hW5Jibj83vpt68VUYVmrNVmIN3nLqFiUP6gLRKjYKtr/Kc
jc3lvZ8cv3JTccONylkTeB8dG3EFDUgy0CrErLSPtPRvzVqW7z4qdDnaJnoFJlEzIZX6GgQKi+F+
0NNjIjIh1N5zapJD+/PP6IwGis1XF+Gnup7UmG3OtGdH19LQkjrB+XEx2TNoE+117NOoD0SsiQE+
pXNjSFfkZ0eYdrXrQmssGmYPsadeDNxXx9/ITE/O5daq270BMBAjrMjW3V/EoQB6K/ALHHvPiQuR
MTb5B72aR/cJ3KG2y3Fk6emZ3/pbC4CwT2cW2YgXvev765hTOP62KYklYEnX2jrprgwIYTgJyT6t
/oZJGdvS4UPW5ZWLSkF0eF23rRQu+5X7qvtXcs95rKU30MXwx4WaVoTk6uGasg/PRap9BFL8r3yI
IvbfnMtPrkje7+MGVCCfiffKPjzNL1i09VU3oZy6UPSjwUEW9tN5talTqKtvq9IuIgchl4Zp8Ikb
8vHLHMNC2Tb6XHrXDa50FQD0KcDaKzyqw/pVEzeCrgqBVgpEtQFyXhkBLvPdo3lBCwAtQG5VRCgE
kOFogqw/5nTTMgPA7V2UhDKQd9C5Xa5baYq6HPr036XyLvCNtb56dMTudalEyPZajASdAo5a3A08
lP3lyEIJ+WgosU+8YS+dSjO+bFTwkuLEyWjkbwCp96UC61sofsDQNL2ZXK/obrQ4d+m4HVAntIZV
eHiNprTnPs+zO5fDHqNNfHCw1m38U6EYt5l6JE9Y9LlfBzCV+QGpYJyMTfLJYSDG0iecD4C6z3AU
6K37MXtG8jn28mIp+78rPu3Nm5x9wejkhTLLpKiZm04XqbDvGdIrCqzLRFw7R5/D8K04AVLQkW5C
sEZM3/7rVcmBL4t4znifCmLrV1g1j2NLB+1rnZ900A7BeDK/IgLTlQUMLtMTZgzG0Mx0UFoHoYpQ
vyUa2zpoV3Lvq59fdX+LTSkJlOTTVaBe9fSE1lMXpb95/9amwMF489xqtJQWPKBWF/HIVgbKScX1
A9mpdaVdTfo/PeGwEt5f+GMTUsqE5vmP6nXZTJUNdgvP9benvfaapdv9lJh3skCn5fpVSnZSW3nG
vdigIRu4L/gZRXC1AzJ+KOlP6Hcs7CvMekRe++HIBGbS8y0Y+RJEjXbSvMgsnUd+2os9DdkMmxFq
4JCU8K0J+A+1tQUi+818m0TuzhMPjugtnzVvfdMF999NyCRZI4IA6zWhYS8KwrkFpw3GjxtFdrQW
BPeHjD3z3EFyeq5z7VR5lxYbdTC3NFn7H6scnSbvExbt/yPIx3qAL00kHNDckyBdIe85rTXyyXvk
AC5ne5n+sxDP/x48m2nh1Y0X1A2ismvWMNeMsNI0FmqmFHsDPn1cb+8FYJEaVKwFibS3M0LUa4pB
/+Uzhl6VQJO0U1pMwhF7dKjLYrHujCGLL4TOiS44lue3+7lYow/ccF3n0meSSSWLwaUZfiCdFu3R
US2uAWPCTRwofB1s314dSO+LBwMDUrgaJyIYJgW8TtghmkKiwJfZgcraY8YIrCbv/8CV+MRClCWu
X4L/AQ23WnCAzStB6x/GLLfSPozTDgmm0YfLeaxT1AEDO9fB45CV5K6Whv+DIxQ5GJWcTKpoOtc6
L70xeVT86+AU6TnafOGHBe7fBhwZBOWpGUfIMyDBGWqFRX66Vk0UqN3O3tOXVirYbWdUDXxhGtWk
fx/EjrAo+Xy9LF4IHdvQTENlUVXJBYT36f0lAkWlQ+egWUJuz97+CB75yqVoLX5sL/XeuK1bjBJn
0Uv70dPbFAaZ+5/zPa21Ri1uxrZooKo1fTnvzQcKAFNZmIp3DPLr0Atf3seSsFGbHae+coh6Tqmy
Ucyn20ku2W1YG9Zz9OSjDggNc+XdTXmSyx1ost+DE0h8GAQUxQsNXyhWx2Qgm8WG03XltITY+aYy
t8WdWOZr0S9mg8si9IatowhZ2rn5pHCOHcDfWv3fOrj69LJd3w93UwFvM3QosmiN/CvBT8VLXi5C
9meLKLBQnJ9jW0xZnOlXrtdhofaUk6Sex9ysMU4e2bWmSotPWr8MUoVFzyPXXWTzyzXWCsmCFja0
LZlgjhmhIv1+wMaRksNArkpJ8U+lLMpnzveeGWLvoBAaqAruWUJX6+o8hTQlFSNEVKm6D4BdRbnD
IK/ca1GXuKstdaXm/S2T0qf4AFWjNQtfBmtYNM47FUcRP6PXpn/cUaf5ymGLuKnW7gEk5eLx2lEl
umMYEuawv88Ne0wOFFJoQ6kc0IJCj3jsHa2JGYzBOc2P6HhlQtBrxdM+G1adGl3YRdruY3KJmmVV
0yXXp4XEOnhEl9j0jTs5RlU3Py3wRdd6c9+lrfwrfR3GYqi35evQB5iPQpzPLntElf1hIeTChrZt
LchabAvbaiLHsNaexeGz8YQzobpxry5R0ScktIl5hhPuRnKsgZoXs/zu+A++WtQDzU/wtVpbdsaf
y7OXmLWrN8FUAAV43U/nnzxy3U1rSu2u7Usf9S8wm0DEOjw4tZqt1EPWEpN4AH8vuSxP0tQcLQbV
N86uML3AUf++vgNuUra48ZgKLS6Qa2HWyRhAl8uDDJcqK7i1F1Pwhs1/05MxcEaEE3SNh/OiNhnz
X5o+wSue5BprlunoTU+aBE/IMCHm0+DhJ8QmzMIKTuV9RznV76DbRWqPUPvpk55kIPwdB23l0cW6
fcDympK+LCX7zOL/VJsEA1yg7QYDBDsyAZi3P8OKd7cb4bmv0E2Wfn46S2VL8I0Y+Tw1QlVpzsCl
lJ3Hv5RXdUnNj0fZsJTJLoB0ZKbHEPjg18aLYygzYVh7Qboo/+jDEvCoq826wwQ+K896PyYkmZMk
Qb/3a9FBt4PPyxfWienrwOH2Yre0kvuC4P0G4HJUrfrTq74PgCiSoFd+nZKWyHhuIiXVwMitf3+3
YHnDaU10XiM3cXWsKXeaUljcWXeTzbbA9eSxhruq5bn2ntfeACBr+6dbgkjyY/Tmgp0k79ILrvSD
NdWpBBn7MFBH3BEklsWSJATSqF85PHjXm23n1nFY1wpFQ7xF18Fmz9z2U1pmkVPyLADXTG7l0Y+2
AJs1ZOp3muym2vTtT4WtgNXnl9cZvDEpBzzYUuTnYFDJH0XV0pzJ+oFuj2InsGKR5MWWkcQvzn07
NkbRzRjhCGOOSfp6VmTAIeGFnQe+28k9SXY3B+ufPHhPM/x6ul02Y01u6BztxZPv563XlCXksL8f
58k2NiIkxHbcL6KgNn8rZyckLKoeg6diml8MB3eggtKEd0XKLEFfoa/IRIPNgUlc2lTkoRgDmMvP
9nQROdixSm2evDd4Xq8Rf2ZECU17csKJPUr6IXA+jk3+NyqbnKnw/SpSDhWSMPRyPQ0MeXuRo44u
MSmPO35tlhuDSb3/Nx34mPR49xH5WJDhSe2hA7ks1p/x0CSLPnN8Dk480xV/sEgbwsjsqtEZDztO
AgTwozqllYMOdndylT4oivT/pvVKmRnQ9GGV1rIPBMNpqqvuSIqHjdpJn0F+E67mzw/9Lzx/LE8e
p0741CIRJrqRa9iQzOLrG0YJuuyNpY6TuTt5vBNttlY+nqc/wNoFDs2vFcJcfjmxgs92nvBTCaD7
Xvm3BBk/sr3IUni4zDjpaqLzxBa6D2JR/WRbKJr/VJ+KncOWGH3O7UBzYhxZUJJ8uHE4t7mWlcbb
w+Gcm03UNzTzXbucYJCTiJlfdJ2NWKoFxfQp+CWuVoYDZ8UMOCg5i4DbmuMGrPqi1HAW2GS3Zd4M
JPCvaq2uQAN25ptnh/Ub+7HjoTEDEFJ2GQrwuODXeNvyTHggN6R5MpjrQq/1jjcd682RJkvt5ZyI
BBDdozN0XIik5bgAtKW0Q5ABJbNEqF2yuovdLIFxKMCA4iQ0ANRiAE/hfSbSem8heXrcfC2kmxs5
PdypGMnrLujCgj8DelyC2Erx7aflQ4Z3j0ZgGo+ItFArDuQ+LStyxiprgA614GFVeA+lqtXfxzdc
pjZyw2xITye1wBAcq9lgnedHiPxlDFT154NTLHCeLU11dNQ7D/ydPJWHKkb+SQCAE+2vmQxzpwvJ
50NOK+QnC3a/ZEAp6c6kKxsQufAh/VCWytPpTeUk0Cfbv2u3E1ws2WIqzU0UVNrymGtzD8BmHsRE
soFuazewIlO/JtnM1dVxDcYs9O4wIGXgSAhtgUXRgvxFFkt/NhlMhAShVP6IF3zTH8k9hzsoFSqs
62oThzTJop6ZjkqnlBAH+8vpkOyxoiOBlEAbByv3p19tSW/+fz4lLSZ/VK0MLmGagBH3UwssWwyS
miDW7jO98eBM23L2tQi4pfNGynWC0Ve9dI5vs8v5orNk5N0ZgeJEZ6YuooBlq3DP0ZNpQI9odAXY
HNcfxtR/cVd4Bd5iM74jysmL5Fs90eIJcH9EoRQiL3rO+HD30/QkryU1w7lg0TVf7Gkb76R52KET
Rs/fY2YiW0C2HmZfQf1EGpneMEvATWZ5slfhyAko94FoymoTcE8tzex/tSC+eBAFyS533DkhVkKq
73LveC39UPIla+/oGnhyVQiuTPJcX8zL2e6pzXeo4OdsWBxWHAEda0yhxXBsoPqQOanJWPlUxtPB
9hNoEKoKkGqTLpymS9V6Gw7VFwSXCx1CE2XmtD/32m258uLoXcYZd9yZrViov3FJXj2g3Rc8tL0V
eDtQrCPIKGG6hcwBiYLSBd80Fvm/cvXM90gv6USoe3AM5xkkBEstKDN4yVH7QWY6ed34wYLRO94r
LxQ69M+Tcv51bxA8Zgsr0qLHUoTUlSfE0qM92jA4tE7vJ6klBROWh72VslfEoRUJXw/6fnvU273V
OZQzr39jG8lIS9ANSGF0dgUVPH6TFIsBewkZipSV8CAWn2GbzWeVnYxyYoPLTpJQZ931l/Dm58uA
dWCLK2R2Q2ZcBw/SF4AAbEiCV2KZ7mrL7bylejyOVnE93VyMYZ9l/GhQTdKeR6iZ9W+iATyNSZy9
tgyfpEF7rf1XUQT0J6TgLO5Es9glT/3YGe5IwM4TZJH1vTdNXZ2G8MydjzKQBflMcdvHS94kqDFC
H5d39xFOKUHI3ZAKJwu+obd4KGfCoRRm93LQM9OyQI7zJg6PDQOjyaZckkwaApOp2oQwuOduyCy2
kH7JUTj1XcAc71dzKv3TXx6Y67bn+Gqfjc3Bbo3oJmWzTnA9hdtG2JB6Yj5lhGxz6MfGxIg2J+yR
N8U30D9DgHql0Hd8GAjXRj8Zdk9udoID2kQmRSqgYRRLZ2YuHCm7IM5H2gAJ9E8SG1Dt96gv6/Y2
JHzBxzswgQ3Np/9QFdJrZBxX9iayI/Iwg/W5cQoLYYMxyZqLF7ISm4JjcIsUN0ZtDIxP8NXq+M8u
6Ge9qiftysxNZEekXQnAU6wo2qlI+XkeDEsKtZRhvw829BTUAfwdpRiWmbFzZlbdDRfZ++mhi/P3
Bi7BtFGEEMawsZcxobCZE7imwulsEE2fHJdvHaGn85a2ULCOQ3TUTt5P0mvmzW9uV2AKV3GdKHpX
T0s0yW82KtrNQiBCe4/3RnFNYjivPO/Midn021PeLB1Qhv1PuGLu23j9RqwaPxxzo/TFA3sqEfpK
OoYMqiWYf3uPkAvOw3KEFzg7GcLL/7WnmoTuhC3lJQwGOM3UDD8Ge7FOmDLedguCqVJFEr2cKBH4
1kkjdzdFxW6ljwa7I+cU6KonVWLvymzj3/VcXzc8avjRDQYWcY6oBkSkPrcKwHOqOw2IHo9RO0io
Ct1Tbe9Gy3nIw9MWnAkNHgY9SxHjDTadg2ZaiMRm+FPNStaZxFYMm7jFtHGbZL2lXC41LEWpKs+m
MnK3AIrije3AglwWriQ/meKGV+4FeAyxRvPUpZDvKPl4nf6Uow4hDmJdJQKT2v9YItidPA5jdqH+
L7eGG69WgwNfP88ClT+o1kzH+QIY/7uA3vMkav8TQ6OD5q0y8nEp2+EHQmGRZvAw4JDYnC/MhVz4
S+7rA4oqE0aarNuOMagpIUAu5GB8Yop+cSEUjl+peINfe5h5WLAxhjskAFk9WOq32vMGE1pueAqZ
MCQLySpE2BidT9HeVZ6z4LuyT+tqj+lXiRhQJvG5K1tKgZu6cyVIa5aKhDNVj9vXAvpx7E7D1KkC
kUgwF+4qgEytG+Ty41V4ZcvEho/XVrJDP9qOar34iQejF5e5KqaCw/8KcxNausjuQ/V9ZMABt4fK
m2Adgvkx37eu/cvZVOXCYP1Sahyd3Z5wVDtWGxe5rbr9ksblm6mMhjqcZ1teoAid68ztlrwRyzAc
+DRjXTxmCA8kRO3RfSyelBP5x7KgGRVES5nS7FNEcyVABVVMSLpvUteE897Q90bLit5W1/FoWGEo
WO/XEvTBV90wUfWigLnYSJOromNhyyRW0UpXmW46hJxm9FxixrA5DvauQnkyElP7RG+q+P/FcELg
ZzjHpFifQcjvz92UHS+XqrcJyxbM94Hs3mZpmvgsVzPzilaqfzpiAolsljWPnOugWRnYBF3kR5hs
Z8ICTw+c8npTZglBxFL3fEIKEcgfOlC4UYua+o1mjt2w2zsfiEBSVrhoSHE5AmL7nPOaBBbQT7Lt
ExLyzivWUKORU+F/lLE3F91dHiH6vJ28bLhpoP8rbHoIMi8uTH0Q8M2Gffmj3J3n/P1XvjyjuOR6
c7N690vOOvG1RV6+S2O7+P1GeVcu6VVl1/pga9KkhJtPHKsZDbHt07P+8z0et+zP/MsNfH3TJcZo
WGN/jCVapt86DOXWeAXyrDAqvDOa2FEfd0/4nFLKeUyFW5GYbPCSY04lLT+77W9Hn81hc8D1xBmQ
K0+ELrqA6S1JVvjmhhFhIllnEBPBTai+e/yMR9OZNQ1efXKksT1jAZGoj+IZg+mwzTLu1lIaZkpA
gYivA0K6bDXIrW2N99lzBPMYTcGEpNtOwoiLhRuGWOPB/d/CRChfD9F2PSgjvH+9Mqiag8y05X7m
eVeGs6/f6wiEDLjm2IBirfA5RkVJaqqDZ72EZekiw4UDxICqYnXb1j9e4nezxDt1p38II5JkFte5
30YZFktc4LtvSYOn3IN27+yPupmFAJetrIaJj2wBHNMpVI3iomDX+m6vjhg1MCTQLaOHLm6L0CXH
dzeVzeV0O82KLb9MluspN9yeR2i55yZ5lyUGJPZtR4rM47hcglP1y9Iyl+jY7A2Z7qCZj+5YAHNM
hT8/7QWXJSvHzTpwL3Lf8fbL2KArl+HMOK4/wXjxFZpHzPy+CTmuSh7xhSmmI5XtWpS2S3lxljtx
gEJXGu/ZUwkqSJfWxyZaVKx2wyjk7BYWIyei+fOmhCzagahK9qeU9se7N1wcyXbvOliTSZYhWg4i
PqhTFj8v/EVlZB3iju26QYWYr6h0I93dwdJ2EQZH1Jx8ZrlXCuhm6DQEEYaTmW7ICpnhqouFAukD
VBT2jBm16/7A/IjuSXKvrYH9IQEm1npZv33LTR6ZNI4kj0kkWngsJvWVNcnfnLnaOfGuE6juqPed
iF4z32thcfRpHGyqo6Fl4oeKHwD6XKyfuQ9tpsiQT8+3YABqed8r093wpkauJuKZW9NdK32FrIEv
Uv3WkZuHBtSXxh4dYO7SFSz0LqO6f9RMp/yhcl4T7ug/h6Hm8Q5xeHMK7n7sPYJLgE3NoJyZfmw3
l5oOGQrdvpC1lURpPpCcrpJwVEYu7PPWRK+f43W6nSiVRsYPeU1a/PAB6rFaLXsQb7HGXwNp8hT+
iW0FumBrIfSlKfTQ8fxSQsBC4k0tx3bZNe7G56B0To797WQVQZk1zKJRuHv6X89a6h/k6VCJwrZp
6llm2OYonQrb6y0nflbXeyISeTvtlyGzU/qvq5ubmJzmuMHkXP7r0FNCGR0/Y7mwGN2ub0BRzUIE
xd91PqEivs+HVzrzWyWLk+QyGExk+5ATrIoCeqBrw4oAr+2kbIKZKUptB936vLF+XToirfrLpfw6
xDL5ywvuCfxT5ExintL3/FBwLufqj1VB2axE6fMIe+HAgUUYIDjmI9vy4LVVYJjd8Mk0WqyUs2Vj
bBjwAJlJ+DVJXC+5Ovi/GdXxltlSgVlvsVsLGUtmbqDzLg8/DKZrrnTeJtp2D0iXNqB9nRXqsR16
zD9gmmoXq6Ik1upo9Vj5xBZvbOVdl0zIPhlL7AqxT1zsYovnWSZVkRmq1ye0DuQENSjr7kMf8YEB
iYcwwkwvNktsKg8yxQoD2sto7gp2ulPUlhDjv7lWwBDfyCAPC4NjOtCvwMRn3JxnJx1/MV6kBi0Q
hOqFpmhUnGo7vVHG7G+m8OWaiGH4oeQMFwpybNzcd7+fLMUel+GG2CrAH13OEZ948qKK62JwIYsE
gPRIJhEAF8VuK1NtIIlejBnq4XXCcVQ49dp8kxDCUdz1sLonpZuJBMYD18ZZmFk1ibrbhpUNQ5b+
mgie27wX6r6XsiaAEl8+0+1WJQPopHUvG88mKdsu2tQqY0USeAcLSGCOwEmNji1M6LHN62KR6jMP
hfsQsB854W0eorQg14lXsnKl35rUQxz5RewQUwyHfxcRKA+ErsdP2iGMn4ihhk9b0v2i1N6qPWs1
DTbKYPsSZeybJtOr39McozP66w6njRQnFg9twE5wiAmePrcd587/S0KxG073d5mGjRCGRkVtHyiL
+GuHDQFT+Ja3UzAMtZwqUERKeUkOjVRlHLmmxgIr4Ax4JLYNvDsnjyTumuuVFcyEZrDNTUkz/44p
oGxNZna2ENdn/7IBvRvKScv3T+3AnFgfaakZD7e3V+AfXUqo8lTX3+sy0dGDQJnBV+qfN4JF7N3w
dJVHALaxKo6Z+p+sNOSuC333LpectZMnokyUqKrCCBsQ/5kjejtHRSWsYDyr1MisXjbs6E5bFcUS
5JzuitFPXJTrc7oemkjdkBGXtItyB6qnu3Elv6Hhn5ifmE4MG3Knr7cqth+V9MD8mDYL614eZKlf
8B8TjyKMGLiJTX28d5jSRLeqxJs37BkwWgqP2N+jKk78xF/Jpc+BddwOsW+j/JG3MIoyGiptgbQa
NtT7Vg9Os3Kt0FdKlJ8+IUdxcN9Lv1sLSJAI5z7JKkmsu51l2stFUsp7V6A95jpwMzj0KA+OeWyT
YlN+yKG+Q8D7IUHxaiI2J3eszz8oq/SsWGpz67q/XqsXmIH4CnKolOMCHYkp9Og0Hk1iWtn+jALw
KMia2LKqxH5zzmEeTWf88921RruvrG2vVC/uOFWklCCpdif+ZocRrFyvokVlor1UqKDdNeNRGYoW
rxESRi3BfScDY54mRpkq0195KwEkdBRHzDBc/Sqk6cF5a2E9qCsO8PkTJawj9w7BIkbBnvkE+dFc
hTcZrEESBvEWq/VolsuXfy3TqMH4vzdo2tIOYplK9ujqHz51o4k6kqDM5CrlYW06Yjf4/FY87n9k
E3d57WTtDDnWdtevYEnIxiiNPs7JgjIFRHYVIZ5GQ++9OLnFcGPzALBbP9YeznzSsrDVZ3ih4/EG
409WdMWTedHTwJ/VIQv+DCsYdqfLPoIQtgKeeau+x/e//LOUdr25p3SRrCHsAuPtpk7WUuEV11bM
yxt9PNM1KWLTf4LcrEBYracHPaKooiDhQHu22pxK38a+MDvTxkfZJ5LI7Dih92xen3rwNcdFVpR3
wkjsB+Pt76ForbVgWnwrtcevBXH9gbug0qt87d8XRS+E5RtMY1CK2XHptz1LgdLF20vs39x+zowX
BXykVW8x0wsOQgcLpYP7H4dFkbdAx7s5ffRRKGCLnwxEfnGwmsULNz4B+NgBG68fm83Lz6yTJAl9
cGKafAHxElIiwKeQsU/myR97R6a1hwL+/ThVbZSrPgjHGSEqye+kJ2H93rz5mi9t04jYkOZXL9Wq
kTVrLgKYuJn/+AyT5HSh5Q9pVelrh2xGI/kiWSs/vmXvj8YhOh9XWWS3t1C7BPh6HKq6iozxEFhe
J8evMkZE/L23iw1rN+fiVg8FiUroMUgTRSc/LXqzUn40iyloH42JFDa6b/VqU/qgZU+JmYklBlZk
RCL8yKJpRI/4LPkctF530uk9fHblm+wqUyRx0uXaDLR+qGe4wi282aKLLYvcrFKN6Ty9cicVe4WG
iRBhOUrgQV44YTyeveZp1tKc/AbUsDFK4A6hc+ZV4h9bj1Q6kNjihTlY0zcWwRduqgf4L+kpDAZO
ZONyYXFoDCaVKBdxCNT2MWYLjbONmG6mtAJFWOJuAr/jxXhKBWjy4o9/mQZbtehVY6P5vXY3IAON
fInovy2MroNtR3sycaxhy1tQF2+BoihigXtfHT4+BdRhJr09lx/7Yz7/MuurNBneaUIJETcWjann
Yu+O0qf+yDECN2ab/Z7C0tU2/QMZ+Eai+Dgnnia32e3qBU9PFmpzPQL0V/tkEpFMv8/ILNoDL5E6
yIVyRJrqPY1I2WZsH+6Ob1RXLOalOVmOi889sfIlR2Qr6O7xBv0IRhXVWN5JTKJt49oXi1MReJcg
1F0UHgT9GLg8i5ZUip1Rg/cVO4AmXf7tMEMbPeURJJN3DpoipLvoKU9nyv+8zCZzLjKPjfgQMEGZ
Tjo5qIemLkPhy91ds/wUOu5zi6k+xJ4/zSP0/CDQjuJZnMGHFHg55tyY9Q7A/FshaAtF1aGMr2/M
iOJ/bX756v77qB98hlBnSNwkAwI/Lvs3Yw+Oxrgj57yhFhy7RcgOhzW1vaRWgY4oLYoYGh6OidaI
veZ3dD869sKRx8K0we2RjYYaZxnKfMGqh1hBYWxxQELli/ccUyms0xmG3MSJi11icOQQswv46LIR
sehya2S/DnbGhbWJLKR5adiZDvSDjulY5uNQNGoOe5yCKyR+x4RA/Q/quvhafU0EJQXI2lp6JSX8
9G4jsMmLAfrjQwPo8uyvF1qrcbr6uaKnKsXqULPncGKu7MgXsDtKDrn1MDLiHo4f9k3TMh0WVnsj
PJhkrouBcrVrbtBFkEOI8k/GzvmUd1Kx+3Gv9ia9IWD+eTm1bPgVsj47OVdg0gT+i91ZgURCdlZI
DDDLfaeaRfFSG2IyED+yP1HjbpSqafrqlGaEECeqLjRjn2OKRtURbBWnvbC+Sgy98U74/wIQoTWy
kBUsA8AIWmCFtbA+x+kZnRwFPb/t1hWnx+phK+Bw4Z20f3lUz3TelQ5pPZLvpdlOrVUKOrXlAHhL
tJGF8ZjjUUxKYcuhUQDJy91U7fQt8hlsM+MY2+04fxA2gGK6oOSIO5eMDt33D6OhPAxyWCVsUzWY
35PAIEn4SA5XsKTtjCWYeTqZTfkq2siCXzpY0qxzqWo1gpi6Q4qQ+Hzz3nM0zNfH2km3KjHQyKPA
lDU2A694xdH+Z2QkyCN6/vS6jzlkh59yIyB5bgD0T671b0RWpyJUbSrmqEcD2M6k5d+ERwwB4G9r
dQWM+gcCqY5hJFaiwAg+skAwafprpPog+yLWeUb0GOTLjWshbJWOz1EQ2yXVxQ978ZZb+AmPd0Z5
5+cTdp5Km87AHxm54boF9242/HQDdP7VwtWtNDqnT6/4nZJ+L/rs+DEbbtN58RyjHzAF7GylW6K9
80yuC8jSdK1tJD+9PzTy0dlBuuPFsf3kgQrz1fvtQrBvB+Sl3PkQHQVEz1bQq3LNAXjTJLU+mdh0
tXh7quSnRoUcINVrzyaLbhoRa34ggFgbIGBgoock2Kmo/IfTz+HWS/FN3zQln2VJEEMBcKka1NaI
dNAFa0mRihJswzv4MUMOqyBMhJVftPJflGp3sC/nGVmVMTocpectCgJrU+g0bgwPZ9Aa8hwOdhw9
FrDlHuo30xj0jqQ/ahMvh/YYoEsq47InjRFA3poEjWcGobMbr4NnI/sEtL3uY9DMt3JH4deFLXQM
UN+BeRfkDHpLZq6VviOf/mlKUHNuLFtq8EQ4Kt3SJaSXBFzmUio2cx27hyGUU4fA9qAwYc+GZSNx
kmL6r290MnSXHliRXloZLEI9wjkc6w/bvnJxDTxPmK6VrdYT0hmM6QVZT3HrqoT5KLZFiOYmQWm5
f7F5c9ECyx/oGs1c2rFcfU7uDG7J4fzE6+WnEyHCBIlLhIkoW4I6T+zK+N+cQFI5M9ea3MCoLJCN
8rEMRiFYgle98udCstUUXhkhR96rFO3n++31HU5EL78PUgq/M2nQebmh9Esmy+rFfSCJmDZO/3ma
cNZAPwFO5bbuWZ+ocvVIXtlalfM6jLXjScIbhtjy5Ku0L4g/86wm745OqEecGkJuK7xe8Z6hU20U
2lQgUY75JgFoHbiBu1/zDqaSLnsWI1drjqxsBR5eS1WkeTFcVOgA8cxvEktyFv+pf+XJBdC6LNdG
VmgFg/90EUgYQhWZbcPoa7K3ly8FHnCDkovbuLzw1LvL12KbA4/j/XlGWwv4RKpbjc+n1UEpEC5R
BBgTWNn20DfhOXw6J68nTQgXsxDs0q92rwEAHFtiM+Wb1Hz3uZmLxdfs1dUbvLOeTFD5zlnkEsKA
T18wXFoVsKYRGzKqplFTH1lsRrdzVG4WGMeTBW0YGwv3be0DB1Z74th+bRObTnyYAKzB09PghwMd
KkQFi3GP+xSGMaC2s5LXfItnt3+ei0W6iL5olMqejir6BTNKyqAFu+/kY+UYin/IGRDJSbuz4fCU
kDBND+vFR528CvZ9FuADv4/qNyu36fTkk/XoWuhTeedAq3+YzaTT9ERyNyjN6XsHAcmfUMgOL3t1
1G5it7ASC7s0ZQ8A3zAVrNjT/vtCadNHH3zf+437iIIeYm+lZhmvLlzoSuciGQF5tBn3d8BW4G2B
0J+VZcDuG2qXEeOMlxPDyibbOA1ZVNDhpRv2Qf4boXS7670CRaPGH5gDDJnJXknc18s8TaC4Byh/
OIu/8FpvEbUOxkEM5pImKRe0K8e3/sJlgvCePrTLg7ifj03dgdIW2diSx7Fjujro1fH/mUO0jnF2
zQKFzest2VDtB/wz/ZZ1uAGxxalauDvq2ak1NgmVDsLZBbjlSKH2MkKegOO+UeDiF2d4GFmjQx47
e8+DZV2AgttPnd7WMCeMA95RMC8NChCWNVUWDVkM8gJg3r59BGTMbFkv67N+ZZnflof7lwRBAHZj
lNyLlDIA6bBFpY+hs8x3Fxc4nMyBuYkXHXXfa2sCbkBMHtryxhD9pU6TxdwMZ/mKWdy1DUVotpNh
wdtAzdAx9s3GzH8rF8eiaERvw7cnyxXpgb2w3SMFI7INb5CBhZ2vthZ865wt2ysWbNqOGdwP82Zk
iSihZaFcqiWv0qxXjGzJDw2HB1zBHJaOz4+Rutfr9lqy1xmmRGH2iS4gyO2EFhOKXEGC4YTWkl7e
CQfYWhMujO/fet+epK/bCQBiX070F/JvL3cGpCbHRi3CJhXgts2zNVhTyzLRNg8kMYby4qe1cbhW
54uuoERuf7WouKy5RE9JL7d2jiIH2brqgV6CrTM3s47LPkt1P+t9dtDltUIaq+Iz1wtmTRzDQayX
giKQgIz4sG5cUVLT5y2VdEiI++TO5uwJOkwjWFMrdwjH4WF0Ew1yEV2YuDmBHlDIwtpTo3cRFIyC
+cxivh37e9GODtL3ATD3+x/c08M01iiZHc2DvcvHdWAs7JFTyJJIxCH6CkDu9uV5yRvNacEIxDyv
lieB3j74/+2lX7GTUe7glVIFaZ8FAt6Bn4IOoWtRYMz0MfwxQrd9umtN2JbBIpZVrGfe9g79CiKX
qNILb09/dBLBjAxpdPhoEHYETay2FQ3BZbqZqBQDohqMsqqY4zLi7qEi1RTcXdD8wQvhY1Ngxi7i
4aAkoK/PH8fJrchr/7q2IYr8W+kCuPzqt3VRpeMZPFWFixyQ+hB/rgdtrg7WVm77v7GkpJ3Ouc5F
FiNaIKUUDpqRckZgA+Go3k9s4YGHfas69cdKlQZhxfVhErXBb+F42EsiHI50qoqceTfX0XOqEbyI
Chvz90RkW9KVjbi5uSfeJi/ADMWf7T7sLGnxGnh0Z5jx/qaGNQBwB77xq20Bpub7Vc7jnX51PIrB
PLQ98/dOiLArAuYNMON7Yf9P/PPFaYUYYyzVzo0SzHPPio5kgdB0X5hD3n4RD7Xsz3iEAt9N3KQX
mbGBhOpf3mYsGrmnhKKxCL7E0WEJD2eWAsDHv+GdxaRwzZuTiqp1WRmYXL1n25QpOzNfN2ov74a/
eXlLYVzgfIvM1Mv1QG5tViEXlvfufF3k8vvLF3gSz4hEM1gZ+69wn+kQhgyziFCjZloI+97IUj76
W4cF3KVctQK08v+iAKgTU/GbblWUIz7g2l8MUWyf3rSsLYsBSliU2DbF8/uFm8zaBlyjeOL7hB6/
Hpp8FZ8M6Puh0sg/kyY6y1oJi13ekpxDdC4reEw9y6Sxkv3buyi86KeUVQvmoKTGvE9kbq8Ibe/U
wdnu2n7bvIq3pB9qyn6TxdR84fLJoLlo1tHzoLVBDnQQDqs5CaRmrM0S/enShQrHNoRCCnEFELjN
RckN7maN63iKdaGNU4depB5ZeZFNMPWcoN75ijuPQTMNRicXxxBs0YW6Y3nkiM7ZvMiO6/Hwy+ho
/n4x60H7VDjBwNPM6EqHXIUEJ09pPzfvQ55/7xhl+RRHZzVcPlnAgKrbvsQU34Lo4Vh0pTay4L/6
22jlrVBf1Z4qU5zvrqmYYEOvTGDUS1qdY4v2HvcLE5Ozw8Sm4mEEKItEoweH2fAlBAa2FyCwB6s/
clnztFgK6iOII3SBDdOM+sfa5wJrIds2Pi6g/tCydKTLWWnx6l+PHHo6blAJr6dvXpyt3yKD3x64
zHkEOFzRV9FjKRE5knsRTq7k+eHLUnxFMOEfnUiV/QMyYHsKBcxa4owc0sFMORT9k5cnATWm3K9P
w2Zz6HGwtbdVbbAJi0RDje9zKfNXhXmEJI11tMOSTod71WlIuDGzqBbaGuox8cR+qbeoPJyLtB0r
C3lnir71NK7SJ35h7S1+RK3RjGzzAWQ6Agr/AH021MRSe/gQRuNpbtyFl7PjH8pqACx2CzK2jIDr
9cZDoTN6WJRhBo2Zma+DwVLCSAvem3cUJE6bIU6NdSMg7PUmrBphGWNLrHRLaGxc6FtmliRiI59c
ehXUrF48tLOd/vkhtWym9eBcyci3VdVdKgCDU4oJttAJmEcjS5D7rnq2rLUC6ePfBDC4EMcH4YvG
lHkRzWvsRZhXBVVqoUXUbz8zcQfeFlhV9L/CV2Ed/WTzDipiXgU3flS82SKYtrGNn2PKEMPYo90m
fhd9QiJQL1xeLrteXDghLvH3ZmCvkJ4TD+XdpcW3S7eMV/FHL/JghRILaMKUo4H9kNBF6UIkBmCe
xaqY7nslB0OeDSdIotkyO13aCoPp2nruJ6pp7Vg/B8aqYkEq35Ri0+OI7I83LQGLE55c8+pZof8T
PPatw+91UVCan2F4Bu6cgrliUbgO7vhIsc5Z1dg5wKOXJcQ+NmaKcnO9VKDlzked6hO1r7RwfiHo
KMre0LXrirFqQfa2trvVmhK93tqkg+RJfqMiYmuv7iSC80pRxFaAvJwnlaD8cD5pi6CXHM1p/qRw
A1K5oX53vXq9vpdVa5fTXvryKCkBN88SJOd2r/TPxTmKnN7GU2BF33SK9EXCBe82qcNUNK4ZAp4V
f1uDDtwqsRCD40X/aw2DA+PItRtubiW0GbVA/uPZuK+a/jeq6yEmEiyL1aAK+TPuV7wnRqICmYY8
eZSiV6531zAUpaoWvhGqyMiV03T5H/84h42iGzIW/DsqXJcLjT7MHmsd6Ygj3IW3xKKnYMi4SfH5
Wa1EA83Jue3OYt1IwOJDTiq1lJp4ZbUQbrkRrHtbiNO/2O9ZnHSR2Bu695t914PJ9r1LDS7kplOh
JaaptbY/QyHx276anJrAP/OoTkNKTyx4cUS8nGrj1zHtzdJJ1IQ0rgksQDCajGIemrYNg/A5/hb7
ikBaO2iduQfQhsb8cyO+ZAVRKkdMxN7tC/S8sMqzTtJKPpu/JchOAuwdcEnfeBkPQA8ONL36Bmqz
fJxvJyi6UUQyLgHjbUdjN1w11A8gBaEgd4uOMNwBV5BQh9GOY9AQ4eeiKstzqbmN2A1KE3j3zmfd
N+gjXh9u9Qmr31vw2IauKLN+vqq3RjTzXgHB6mOMr+LDvA3gBnZFA5qANkc87gtuietL74BdMkKK
W4asYE6zn3QCPzUIyXeVE4UOCN0/Yzix9byt1Mkbci6qRAzkWsbqZmRs9ObPpg+9+QZVtyAUzMTa
KGfceskkPCedDrDg6r5NuZrjGrcDoFFmb1t5S9OqIJ8gMhPeg1VVcd68IoBhI/l+17AVvXxTMl4C
Fy02RCkuiprwvYL3Oo9BbF5d/mN43/n69QfBcfWdwLDRviim/rlFYfFoBqnuRIqYWyEAGP2k0KnL
nQzFTr8ncCiyjLZU8nZHPyY97WMSbtJGxuxvORynfkgAsyR7/4/Bh6/YMGU5XZk8gaZsD5kHInnv
VveGCpRnFZc59TwH2jllxa/SHrLeMsONnxjpVY3YMWWtuD4HOFybWk6ildf8SwzMIm6Lc/T5yUZG
Gfyy8uUDZnC3jUH3yV6+nJo9w3N5gpCrZ5gG4+sHZIXtxIdqGc+SGimpjHZszCD1sxeyHjKlFraW
dpIiuuaf5ssn6++FBddYfN5+PNkz2sHZ0NAqSNIiEFY/2C4c4YEBPAqkrkQzp3YZkuljgsWdhINz
Nm/h7te4Wm0EPSP8B5vn4V9ZsPthTyLtbqBAxSBtgpiJHgy598yY6+ijXcUHJV4GaBBfG31vAOov
7ENdPtL6p+lkvbktnavGKXRHCkYw/xCXXcrGitNuP+w7H5imwUudPIUTXRKEq3XOdQlsj0FVTrjr
AUcWYuYzrXd96B7pu2lFgdg1tCUPhLPJHdWqBpUOU1+0fwJYsMYhwcqs9txsMp+0YNEo4IXSb8Mc
3c2w0oaq80JxIwtEeCUqszRUd12otl8hV06c7/0WZklfV0nH6L9TpDk14sIYlRM/HKhhRy19FOr3
P2ijWb543SMgYtVpFl+mFaC+8xtN4FyXcBjXoe5FEvvc9VfneBVE6OHOaELWYQEVyCzflepq2pnf
M8+87p+HOoLS5IhejSrH0kuwKzSGTPa/PcDF2yjYQZzg2GsrmJJixYXPL+HRtssKWuziCg5cOJww
Kj4chAUaQVd6QrBn90bSv+HJo03cqxqo7+nomAol7JaTeurqMtGG+E5V0AAP6CglJHXP7sd32NZo
PUPg02V6NdSEWggwZ8vVHrDOeei5kBvS/c6RwLhlBe6OwhMLWbElY9476cxYxo7ZS40wG7InXXzH
f5MOQh4pcWp85hoDESB7g6EkXyWWhpf31GZPQDi4S8O9Rqtd0pfCFXdO4MTczZ2lJssPq/BJBYBo
RZOMOYxDiigFMiuXymnIgGbLQ1+swQZhRkMIbWq/ZfBPoqtPKsTUgDAfPRyspnfz8cGLD+OezVJO
bAFY5rhnw2TkoLOb3fqTgsEdL9aviMIuxEuK6HfxgnJZiEJqjGb7v9KEFo56zx+Mx1OZ4SvEWVWq
jebyngPBVOmDas3VJBysOPPhfzhS+ZLiT34m8wZ8RmkbjQCOpX9nr1Hfre5EcjiZuT3q3QaxLAGF
UeA6ANq8wctJArIPR6k6+/ETToRlBVqtVCM9pYANkhdbU7RfQmTWkJHyFuO7SLsUH4DSOycftFEB
WokkvU8byyXRC3CLeqa/PbOMG1LUIhd0J2HiqdcJHTprJagA2AfCS8ZxMlXgnFwKhaDUKxP9JtY/
0Y5LHEnC1ZanXv26dmhVTJdqnXqHsECvVFDhVz+I+u7ln+VGfrxAImb5xR8d6UwHHQPN1WUJMhKX
avO2w4uGKJsgYowJvdL3G8X+Fqr/RIyWGfGYv2Ak7OUx2hbD1HtTRuLInmKif8Smc4qOYRWEhZMK
JMo4aBdRtPW5R4iAJLbeEFvl3M5BC2LzaXmmzFYCqsPLhJS4C9v/wXXZdeyhgNAU/25roJyqAgNH
6F2yGj1BgfYrcr7XMWuBwW5jhX6sMQ+sbxQO5xO7R+yjPHBj13916oEBmZ+wjUK04BkNupWJgj++
DDj2RF2KYIiNgiERvzt+7A76YVuP29Wm09RJR0tZ+vdBFUTjiDydDub8Lnt3expUDvJVRRbRREke
x7mo6vNZoPtn0JcqDb9cprubmx4BvGkIka8+wT45wPiMWvJaXn+ZokRP8e4G1vVzbBDMzO16qePf
7kwfC/yCqWIl9E8T2LIbBimnVSTXic7fYPpTNpCVw36PTk95I0XtuKNsTEoY6i/nssRjViW4Kmkq
4RVImduf8f/WnfQ6jdfqPFtE1BosAF159Pbyqo0NUrywnffd1zFND2+PEDywc/aZs3Tr7Me2CkYX
RMmgacCgMCrMt6rPogNCVwcxjdQ57+yasZui1ZkFuZhn6FzB1SDJosSarxBw4yxHCMOaYXjOUFQX
KUUFuoTXc+07zKZe5bWhQV7hgI1HHpZY1l6+TjiLo4dID55O9I4NiWgmgUwQagWYJqYuIkSvkG6Q
8uoNRc94zvtbNoEYdQuhvG8eFhb/RDPKckoI43N0dXptq+frEHVnPWdoMuo9aySRVfTKnMkECYMU
dNDqlIx5zihM23dLQFd7biYfnE4wMtwI6EaAJNbMVbLvfsjMvFCYTcbnNSWDSozcqsWyD5e/rQMx
hrmCwrfuVgJub3vvAUQ63RtkK0q5O4VRJf8Z0/q6LjDKJE7VxoKha13VoQyUCkN0vMYJ0aA+24Ru
XtkgLl7VvSNVfQiDtCeVl01TFLmdmJNhTYxc96OOxOZJl8vxVrdwxhqJwYusqSsrdbqP4xdPwcDi
4nOH35FvC+Dnzu4HXGQhC3n3cGjGDQ4WDWtYQp4wuZcTgkD9Z/+WHwvVCR0WWRsRBE3Z6cQ1Ikdm
cjUTjkTwmpQ7R/ECViyF0Tcytu2kgQPTqipmGc57xj+Eeg7jtYdXiV0MvooCe9vc3QhfeJ4vxwU4
36X7h1QoQNjqz9VpUx/K4csXWxUfKJZ4USMdBDG15GM+ngFTKzHWs5eXEHcTFUqvAzJE7nxbuXZj
EnpPHPOXdVwUsd04ByjVO5qQdcsU96OAPHr8RUH1iiUwKq7kVkqmhvjPKMgbg5aOViA3Lz4cQPou
mSWdleICXcLVvr6s7/BE958bsgFh4Zn6XTosSE5KGojT5bZm0le7/VRlon4wkB4t0+AMVaNboK/Z
RJTcx+onz3Dne5patxLAXc9pGO+yO38BAK9KWqcBPzz1YryWszf6mZu6icBOpdxTlEEtz8Tx62Qo
LsMeViVtT8zE7o+FefROZmghV6RfvtJK5B8opO5SgCeYSwegHHMGrSyVsbPxVveA1BbETBG3690Z
32mris7fd/faiIySCq3q92SY0F/k382R6CTtS2v4lE5EYadiPEAzDR5NnfvSPPUREp8Ae0CaVYKo
fRGRWBj7uPId1JRwobAW2viOb9lqUVsoHm3WyvJlYfHpYLY7MHa4jtY3PZHpCX+VuX65Xeir5ucK
V2GqCG64aBOAcOCIHN92EPcrhquMc+6GVjiGJpH6sWUaiNZaxHDumNX5duYSyAm6GK3h4GDd2pI9
tyeboDsLSm1jT6OYHG828f/a8zuBYuIATh2RPqBoO8/mc1s2lALKe3NfXM+JkK9FZm2yhLTd6jL7
h0VOOjVElrDRgJgHu+gDCBm9JGVEKgYxSYd4ufBeig6fG/guc5LVkSDiuPfL06uKsNqf9bY6WeHL
lmTZbCesMKzEQWRUwManxSfewNl4GrefhEu3uskLsxqDPCRNCO+lQlw7DChj37w7FY4Ur9KErwnn
LRVw4L37PkBZYlXGQ/FD8c4aBXJApPyDr3vjZqZpGODJ0geDLdG2XfxmCdXc+VmXCixn0TzwCxrJ
+iEFavIImQV38Rx5SIvCzLPJp3dg1AImLxnme4EvbrWLNokunyzZSObXhRGaY9mIcZoU2yPsqi7t
1yUlnVNl3wEWcIMlHe3F1++m+ei2zbBCi7xvw1mxYO34LbCSJBe0QiB8UszYEoCFUe2XZ/ZyNX4t
pRVTf+s3PQEikiWAkMIx+WvHpBd/h1Srp36fOa3kd3U4Qk1jdJCe0Dswk4SUfmXIIMdtN59nKYRj
fE+E/5Fy9vBxfO90tmZ/jfFbutJ+St+7Eqg26Bu+qH223UyWIS9qs9AhgxD/SillA31ZYA3d+5FF
meiSyEGkxmbqSHbMUxTCBuv/UgqBOPZlw09i+e8zOAvVrbmtZ9b956dvrKggZeF3Pd19OEYQ/kUU
viD9w5mb9pzqiICCMl5pxLN8NpHZCgHbZhiTR01JqcLhbPditSHWb9yk0myrrNcPFvRMdK0fW6lH
BowEZMnS/fSvZ3sVqLC+kvTCo8LWtf0Tc/WqKgu4Wf1Bk/SafMNXr1OCnRnUnv/eYFOmuw+Gs5au
ytgkDqsoSJ9TiFlRZ+LbR41IRTI/pI4tGQESAGtLiibbZA/nUxyFU4UImbB/Rjb/IgHHx3J5DoFq
KjSqmpSE2I2LiEayCY8hvXMTX5MPh+7zc3+9KOfrWIVAOigcl/f44G9uutwYLDRc6WQqFDVXTwKr
CmcsX6oDeY4f2g2A/MgNDqriNRQwKWjRWyehq64xy3rAi29SblN2Ru6eAFwR8zgROksL1Rg/RhfL
egbStIIKlwG8H89pHq3u0sqkaugembySo/aU7nukH6gmICpB/bt3apieIQSK0zlzVm2wZMRrqWd3
6fOAQ3cD/opPqHGO9xGqG4Xkg4cZ/4kDWK5EyyymhBFpP1cYZLhfoLO+inukq53cTybHZWNTlV+G
x06Fj71xVY3cGaF0I2cS5LVGV4ksny2jKfLjTGQv/hwBNfW0pGPnpj3JTOwBiIMVuwmMcoAfZIvZ
j0QyvS6iQNMjUng5MjxQqgIbDisL0Nid7Chq1r+O/a+KK3QqZCkLuOQ92wvdfqq/FDhyLHgH/Dib
DDuFWe5mmSxFBQbNW0BugdFAxBq20KXw4SHBaNccl3o0wgub+ACo820vVuVcGl1LSkyZ30n8Ki86
beijS5HPQjpbULStJhfGg+aA1oEmGsFF7PaknN/SjRxVaFVgzD6mVs65DxVtpk1zRo9UxDivkEXJ
/PNuZn7ZqMerR26v7JOioVIdXzK203rv493tUMD6HJ8ABl9k3ft13w+eUL59+hBo/9AEBh6ulPo/
ed8UU1McCfdtxs2nmlICz7N29GZ8xBIy1ogoE7XONyANbzz63jSAOAtTmlkT00yHZr4IyjxR27t7
H8gSaawMyEtFlEROWq77u3s+CL4RAtS1SfETUi4S8wkhCs4b7T1B9wLF4/zHnW6q7jZwsx7ZTt76
HNThUwsO31ze1L9tkdchgBrEWzs8BzHC7/LzvNQADiM/av5An4wAGBaUplJjk4OKP1jZj3ssrzG7
DQoEicvdCZlW8q/QloM7lW6D3igkXDFWO3G0fJ+RPnBgicClG2gjPJJibW56jn82q/amTzu2wECy
e9NQYVQ+zUk0PDWuMNq7PwUNb+OJXs1IQWL9zn2NA48jQLICtU56lO1Cxfk8opndwcjIpa5GMP/O
/wLfCOLi6Z/rcafSQEOdsGf2J8mAgsfTHNwa/bI+kbdiJz7+1AEnTaBv1cRVHUHchLsjcVhDmDpN
e0E8Fr08iua8yXvywVYe2tuZhD3st/xfMf5ZeotkwZXHJSPQIrgm9yAy8aOne1Zr2Qf+J0nksCLc
FoZcHw4jxuW6Ucs4moxgSZpUZL1pNaV93tkLbBmoiavPNawaKeV0x5dzQv2JNMpPvQectN1DITzN
RdXPHLmlBsshJgwvDzkw+hENpI4Xy56gDsCfZDkpILFeqBjZ2zbdgU0vQsqk8lPPubm5/giM5L3u
+BEdpA77PpHQaBDeXG4LQPWnG+rwfcLkRypCaRjSM2qoJaDmskuw6H3cW/L3NFzuod3kfByxk1yt
5AuK+5GUFsdP+rMJEGjx/0kiYBu4unvc8mldlrhhgBFTS8mjcVmongmQlQwVgTOuNsflPsXaD44f
VsPrnk02pVz1+ExpdKLG6THKt6/qLhBfC43T90CvFs1wBK7a
`protect end_protected
