-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
//TBuLiT2Ixj8SiadVFj4giwxGYZnJ3oLDOgIWPVcdCvqwWU+bduGxI0XzC4SQ4k
RsOF1rs5IiLBfPX9u21v4hiwRxu6VOND3RJMAkNxdpgF6qWTfE5v+6lSNabOjO+S
puYHKj4pSZgLo3TjRHpm2QXZdlA6zPwf7F4QBzMc00i3S/0xwF/mMA==
--pragma protect end_key_block
--pragma protect digest_block
XbfXfN2L/Fw5DAbaa4irB8JkkTk=
--pragma protect end_digest_block
--pragma protect data_block
i/W0y0IUD6lzZo5mKP0sp4kZ8CbfIDW8maqzIWjAwArJekBVaRDuHh1WJabFCwL9
h8INDZkEPCZkxpNHNZvWCgdVgQAUo26c7R9bAs5OtpwKnuCE1rFxjSdwhP+71ii+
THiafozsf4A0qiMYfo0PFicUkUEtOB0JBhBU0kc3L6nNsWzgrE1QR7xhzWe3B1ui
xpOashLTVPaYoUiHBLlkyRcqNKCkQGl/5XEILIUecIi9wR/93bJ/EOXM6dRYFwM3
WNb9SFcbAG7CEiYHIGMDZl66xo3cBZfFpSlQkREYxZ1ScqpOOO1Orgj75BGqAz1D
MTr46MdTXF2uOJuP+c8nxOETcXXqwVDgIx9EKkyGwvu4XMX8gJuDpFAjjFhehvsj
90KufqdYTNAVblD0iw1DfyozM3KNsHtCdBKrD3RddL+r2r+uV05fxHm+EHQiTlwt
18P1SBWaeyYwWBeuIJeiLIElT7Kz8R3OiFCOukvwDgKz+VwxCoEoGrbdocD1T7TC
+ozrEH5KB4wjyXz9M/rucg3NyeziT5i7Rw352Fy+VKpSbo6eqVrt8wX8kIQ7L1RQ
uhCSIv06wqUxWHDilrLY1l8Zn/ezmBRtDsWosVYFos7selcsYVT0wjOwyOsTfzq3
L8pZ4fWeDRMmniuvgc8wctHI06c7RGZGUpo7THz6zawuNSq666V6UzxtAEPXXsD/
ueYdA7mF0Cl1x85OS2ZtBJJj8YIqeSbfIyWzRWx+Dfe4PIXR/mqw0fKJAW3PfN2A
uh7bBTPKD0Tssn1occiUoe36qdEaK8qPi2BdrGjR2LLhiALSnBr/FFbZ28F5I0R1
KWhqsEAAXMo/rBXF9M/pJ83GqvfShOXEI0gtI6KCCgbvIuzHw0Zj7Qzy9K7IglOl
d/fXbTFHDpXKZ/DW7ov4ipWjAKO+gm5+rVxfpsmxBuMl6oUS07i/0oBdOM1FfOI0
aDg7bQLb2/1dOGgQlra99LMJQDC4dRvG2a0ilJib0vG0VHEwEGRgKSGfu6YjwvTU
FY6zuqUIYCo7kkw54NHNi7VR4LQzRKSggCqQiW6VId+R8Op8egUN1fK6ZmE9h3/j
tGK70npheUGEk/5GH9CEE8rsDX3/N3g3dE1j7XLAJtO1McdRpQ5F/1TIm9yLM9Ch
2Sf6b2pcjFOw6cXS6CLUgaRy2vvg0EyB8zQHssQ29FClDUG8C0DGJes2ZyK48KuB
mxMmuc/xiDNhuzj82eX0j1NfA4xeBHcMvaiQ4YjQH7JWs/dsFrQJjHrR2zybPNDb
YjLEl2P2J9mRLdqm5hi791VDB13mIvQx6jrAt0MT1vLHsKw8Z+W7zvDB4vv4TlWd
hZYio2pjUgq2sJq2FW+/HENxaRfVE8dGEuZe+MDA5btJ3JPqRqlPrOvgz0osEwU4
E5xZOq7L7EtfLZ6JnmAerFoiIzPgmzS3P6sD/d4rHoXDnBRcVCXWip6NPwPNOgLS
v7LeXFEjorN6r8IGsTyZ1DNjaMaupVocFNdsNCeWHQcb+SLZcxlXot/7/ooRsPPR
DWF9paTdAqYOnzx5IWFaz3m4B+ChPRgZbuLohfXnIUIF1hl2Z0Dd3kGsQcqll4kz
eDJ5WN7QihQsXO5w1YaAKsiY9pL0hnaKLEeI4E1gI+JvA4fvmvbLJJlgMmBLR78d
UrE+6e0m6OaVh0Et0wVTLpTCuaOksWXmmA0oIxva/5SGLmdxXBwFP6tuM8tUqAMc
2v4FshA7tdRiZAIgrspEPpVpIeZEcrhuOF7QcPeANVZdOm1zOnCFqnWuaKd0psfi
r+BHb+3YvUxgurFeDmWWYexHOfi42e64ZwAKsevp8MwCbYnKXiIF7ye1Sls37Dwd
PH/bBa17Hk1q23gcpqtBsqL5UO5G8esOlWg3uuXnaOoyHkelLVakFvln/qfrpwK3
8YrFopJvIoIMZ0vq9ElhJAJatMfq0KbpR9qBlYbbiy7fdoTZnnPbFpKSL8rlxxoa
dOJ3UHsGhU5B05RDD75LDI9/pLYqhHHNAFSi7qrw0WXn55l+YJ7JW/FES6bynNKe
VMOESGnKWMnlN1UdFVYL2oBbgUGB/cPl2QgLkGX7g2yxFQm6g8ky5jpHzMAp/E43
Q6lE55AGt09pnxbjYIOG/4forxj4XGruZXgIzn3XTaRhsDBnxg/yFVNQuF4wdGUE
wUk1BytG6kC0r/O3phvReUXD96Gg681WFVo0AeMqEMx/zuwV1uEiuvAKut+bBnz2
CnGI+U/DpPHtZK55/RMCqXZ0UHVXqsXA9ZYAraYAI19TXJbYbRLk0C3IavvSolpX
dW4E1Mhl0eIkFS/PanN5zhfucEHtbERKzb9rPh0uyZlGwerscFs/pq9IXJw5Tq0E
TMqW/X5+I47iEmnWUidndkSAlpwm9sQBmF80zryDqb7MkUY7HtbLEQuBtpsoi5Li
rolzas3q+ZOx/AVOd5diF50eMy2mRBoEdo1JmcyY+doT9U4bwHLK1I71gsrF1XbK
TouJ6CqABCWzc53cI/zVhfR2UIyvbPDk4nq+7ScZ8/3H5x2ANXZLEmO3+2K/l/zp
/5hl4OP+07cnH5DDBnK3Wjoa79IipMlP0f+7BJ/7z5uVMem3dgEQ2h93FYoO2tqn
QGPWfuk7c+ijg1f+7COEDgaf5OhbxzMq5kkQ8QesGl8HA92UGmdzxzTrx3S5tCoq
mH+b+5CIJctOTYh4EpEM+EanjQtOtYdhIYj2DHfgEQhkK4xNyNVndiNObdLuCb4J
1MihB16gxtoqrQ2OCccRm3d4/JbRSjQyB/HmVYy8Zg4Z4LnmNF0ThQCQDH7ALbO7
hqc42DEQwT+9koOc914Dv44drG48y/BOYc/2aFOdCl1w+nJgsePnGcD4wOwir2jq
2mSRfTizvhIdw/D0pzs4feWdqo+UzUyvh7f/2SmXPVnHH/x4w7s51+JwYCi8+LZ+
kom7TMGzJ/WH3EWHwWLj5SAvc9zOfTVv1O9y1R01AhenXOZSUWqfGI0bm4MTqELE
K9btyoxXkdU+haX6C7TyIV7GwVmaqzMsklwaC8TJ0FdqyXDC2tgMeDj3c+MHlGMy
ZWiNZ0zKlgoM1R40rtDSW/EGvYkwsD37DOZpQpSjQXWiPXP3MbrVcJ1CsOHYQwwX
va3qEuP81K9di/RZHE2wYhKtRD+O59hawf7RHTXTM/0xH2lQ4NSrHtaUX6pkPeRA
hY7SIYwUJAZ71svkXcF3XMSLdNRiZtrguhdvv2p2E+HJVSeOZugg+AmsSGzoRh4g
+sZj0nostuijAQMSvX1+xzcYS9BjauMVkYIyFnlqfFvAF+Mh+0Rs//zybDhTVpmp
Kg7NlR+gS1lWOcskuR2Z2mry3r+ocdN6NGBJCr9/6mJScvN3mLvEZGJ5/E7I+xRX
t4Msxm4wAlRXQL32xlMFjEYkeRgfSp0V+LTvEWCeVIkseh6T1Qs0EK9q4MnRsmPN
nZFl17AsMEa+dKule7XB5S/YwS/vYBE4AcQr5+zYn2HwkfFBLJZwSL6w/kuUDKrP
FVNK4j85iY1WwM1726b2q5pMGbQC7l2HXKLrXVhfIyxB+DC5fL9FwSItd0w0oK2v
N6SReg73GK8ShDq/xUDqhoj14GY5+MuKocjWyu0RzhLU49Q7081jTz+Sdi9j2IrU
HOaPMOLO04B/mvacyn971qYXY5rregCd2jeddQm35niLyh3r0BHTdBjyLuXwSQ35
fZB+vbJvR5Bi1U53kq2VQWeOQbUNkPvP+WjGNo7x1WVfSj60QIwc5LWQZNxTltAn
AZvJ1A6xax7xD2RBVCjTf3+0W/Y/7OrCRAgYPckBGOg79msGxS/ijo/RWNRYkGqX
oqRTulyavsjgFvFG8Syc+2Omq8erfKVjVE8hiXM9EnfVeAYZdWBIEJna6O+praJg
9MEouoVYZgHWFq6Qr752v9LKgid0o8xfNfcwUPrVQhxMw9m1EZtx0Ba/QrgDam88
Pn0toG4l+cdZeVl7uN8OeQEl8Z5R4+lKzw6rRQwtRKLwyVWqmvLLu2yeJVBlXgQX
Qs0H3DMVGqgb/OeLCEb7csjMeLE9yaZmVIGvF1khjaeAep5aSiI07/cs5MlwV+H5
dKM76dYKjqGovbvcWrs92QSek0kRJTJWrxP3hlmxDIUr/hiuxnuKx1hMxV+h3okR
IQOO2m8qrB8RwUnvKNbWaNcAYMPjWawHO3vVhZ2krjUDHMhJ/Vp2bf2gzK1QV+tz
WAmHbMKAJGe3qCTlZIRVQoSWvAull7AfE2g60AZPWNvo5LMrt3O/UaRuYoaEuja8
qBkoYieq7bZlF592rtK7tzpFxMGzsQm59jN/K6AjKrc2ZczAL6wmLH7oa8eeLLnl
OyMrgsK23dYObVLKuPMi2fDh/z8tFC/4KUCDMtpFnhnXfQspE4acuGV2glIQurNH
y+INCpNugKbyqWtBOCULw/HudVrRQRMdWNVA2e11CsfBZ4ewhudFgTYz1DSdCHVA
qR3rkUSpZC8Yfe//LdrnoVcoZ0iXZAwH40bDDuUENpmRI+PZQnWgPmgaAVNeGvkv
JwiZjXCPt6N2lDak8bG9bERYMbIUhGn+NT1DMJW6fBxV9kXKUkfCmpZbBPHRoYGS
IAsS+QNf2/Uy3m00JWlU9/TQhYlhaDUozEF/y67aRMt+Z1vLoigoXZVhKRTxcu9o
zbdCN8FKy7ZV24d2Mo9N2tV6aZb+nitLmSYqsLGKIsQ0tDnY0K9xcDk7rFdSmZit
AhLBJAxE4kgg5mFUVx++gJebfPiDyQ4fMNwiRZYKrrisB32uknWlVMVDzhxiRg7g
pKr+dH+bI+84u8hvD2+Y87VUPNM4PMseRDjd9zC2Ko9ixaBusqcsoD2uHIC1p5xA
kAW/luY8zSlCT6Xy1PYF6mcP/fJ+peg/kFuhjutAR4McqreC6TdNlKnB8UCwNJ3T
ZsdzE/InqIvvPXlEVE22j0AbGCf5HXHi/XaiZ5n6RbhV3HUV5fpLWM1u5kMdIqDa
DqK9xIW7Uayr03PKbmhw/4G21eQdc/w2dVg4+SmniFHGgUe/93RPKTb2dP398mjR
MwDGSUqk+UJh+ENLZGqsVTG7USj3fLW/T3js5PjuLFcsi5jYGMBoX1QRGHFBni5K
VFsc/fIZsGBbGSnvWZKOEE9DxBrxQHO7TRGubJ8FVw5TsXCQP6xZ1j5V4R8UjIOH
IT5XOpAlnU8PZuUO4tJn+yD/PXK1gatJ6U35nCdmfOF3MvIS4MxltbA/fkLz3zmC
8U95J8C+dFaBD2PaHstyMbLX/ZK0wIsHjjp4EvlNAErCOaXRj+OXw2DNgxj8gcrT
vDkLwXYJFRPOgXnSO3Rnkv35GUeoLEbEQ2o098MkE/LZ3eqaFKR+6ksdc/MWrQLO
+JXgz7CWG2Pr6ttbPYa657BBTtirDsk7bAbu+vZOfsWN4izPrT6Pye+LZJwYehQM
WTpxryvLmLItGstg6xwtTx+ZDVZKOJyJiCu7WWKm+qxNtTQZc3UXEfQv3BzKTg5p
nUvOdxjR96+l1LQ6gMv9RCgKaleods5MjSTYZPuxf5yDj7RtKLR90J1TftWByZ2P
9Le0gc5LDNrBAmaeTVEo4TKIV0XrIU1yDJJIahszwDeSXb5+XZnOt8AIby0d+rp2
bCtfRNrv8PJaWXnpd/+T+BZIOK2E/99jAKWnqq5qQLjagF5Xy1TrDxW0lTlQh4eS
yUlBodnl9qYtFQ9gw95TEOd7pDi08HR5I3ZqDDEr/ldb7lhvb2/ro8V3qBpstzVi
Y//uNZp3nTJsanTGMPfj5duo6+SVPMR6OO/LKQ6vt0jXydsYxtc6F1aiWGKtJX4Z
idjC1WFGvBGvKuS9fEseOOBjQxQ6KYW/qU6687I/kAGYHZwn6XyDLewMtizDucdp
8Lqcp9brmjzcLbHECAPHxUkP/TBGUWCt7A6P8wYh2zXf6Fh329aCWR7j5ghzm7xd
7vZsBPdvnr5iEV1dWPhdnIEOratejIS40FVhkdngH16vk5YB8EH59Dk/XVomS7CZ
EQVl3bkPsidioMK/PsxJQ1rliNkM1kPZC1G86mJmi1cEyHNEzeV1SOhFO63J2TGk
McYXnqkazeHiN5Klkptd7XIgM58Tjo6xY08/kAMwN1PXE2Ym8LGnxKqnv/fgYI32
of3wst+apJQ+g7VksD/RJ2nnROBY0TsH5/og9/6iA5QVEDGx/VPMOv75QglCV1Oy
IFVzMTa1bVHNbgLAU4u7lL43YegvcmZ0vNn5ObINAdPJqDhFBqXi8Os5+iJqHLpW
WJyw7Jxd86M76KWktBXjOQQ7SgOn4YsWMYtXjpXodXv8Z24iOouYHepVjEL2GCzs
fouds76eaGANpje1zDTyX9zzRiikqnN41JJM+3EvWCeJz6ofr39fWmzhj1NUce6P
+u9ZP/ixCBfrxAvb4/fkwjLjRcyH1lwSpQMvQuUAbQO5WLEP8WK7U6WSoGNiXtwY
yl+o7WU3P41xvc7mdeweAtfDoxm6B24FocfCy6hPxrPwqBji72eV170vbXob/NYy
KBFf0QlwW3qKW9o3pH3pHyE6/TVgWADA21tkrCAV3ZjprBzh/hDodU1aJfV0VdjW
zPue8Zd+meECQ3JttSKkEvBrieSMqIg68nNojjWuSKkKctX2n9RAjMw/loXIIZKv
l3rYeZSvPM+MAEBnWR4Lt+oD+HmgSq25K4QDOHjBXZEig5WbX/SM2GUzbSY+mgoC
p8sOUjk8sMhJ7JQvcZIUp82YfEnmsDDUrVv0FU65O7ofbUtnMcHhW6wU+3noRmQQ
uXq4h4UdoLNgH6rG+H84QUio4jbTdurjrGUtrxEZSeczSpAIgWM5QjIf8vNhqYsf
wwgQIAV603nbadN34X9/2wIW1NlGEJD/KjGffWMxJIvaM8rkdP362rODDviKcHFN
Ojnb8cf+i3hxznd2stwb5cDy/4vPz4/2/Ahxyb+8YcyNWZe0GN00P76cmeNa+2pr
SzPDIKcIBJ4MkRDt/hYPQmG2SI1AUBnM1oao45vqmhG4vtedSa0kUz2uJRR0MI+/
fPEglUUt0uk/9H1faF3/v5B8WtZOa+8Tg6yGDPCQMbczP0/neb9Q9RSnnd9dN7pl
kygBe56KPCpZHJDQcJFXePYEizPdsjcP5euQIrxivGsVFJT41aLm67np4mkY+Yry
Y0YcJ0rrI1nJpGWTNDnm48amfOdLurQAYRAd/yLbwkvbFa8FFJauhiwSleYp8MvV
3THVdFt+lfmfE0aBTgB+G5hNT4InoTT81IbzRdEpF+vfBkV80aMEJnM/qAz9nNIS
H/+Seio+uwuzWY0X5JtoXALhbLHV8k/Fr2TqCxqbckxJfEQHpk9YFSU48y7IKE0Z
4lcZKd/qkjdmK2TG1QSTyeHEuRmCRBHVsUkmakWrSuFPeduPynKm7cclkGWTWZOy
pzcLz1z12fJ8WRH7OJsz2C+16EppeYIR29vsr6nnFrTX2OoSs2Bb3uxnvSy/3bIG
Ulbxj+69+npZZFc2BXGRwvkYpSqh4kHsAYsg26AKfW1EkxPN+HzSJ06GcfafzauJ
QLnbxqKTz7S3oGkZOfDomtrXR2BUJMESLGFleV9cBLpfBGrl1miTVO3RF7XQleLT
fuazW3qnSpHkIm86QGHCoZ22feU7XucxjYe216BaiIcZqAhAnET/V9yVahLc46Wk
rwC1/NxsBE05KRq7/h7ZyKycu6GFEqJWk53VJREFDa9+qSims4pdZDnOQacvJ32F
jDBzq1w7jGmSKaNfDXVxrVfl0zHcvqIEL6jZyI34cuUNY94ClLItsd1BAyp52j9y
jj8p18+SHxLelWSqjlxWq+rdgJZhgUaV+bU2ZopVj+kwE1JQCVIhe9TebPGeOAFu
OfdareMc8+7bdx0RpLQ0zZ/f8beVcNjRN+td/AAJW3rCh8o/8iMXDrlnDJTWDhKM
/a0Ma8Ra3LhznWtD8DAnRIZsByfSHqiaaOHjW0+oa/KNuEFmDxqVuZLBYqPJVSX4
DS27H0Ar7Uan8nAnqYDpOeihQmL0uLbpUru5p6a1KJxeVLdCXzR/J9Egsb2ZjaIZ
tllcCY7nJi6iunUDNRPex4OmS6mbGCNYgS5CCAfYHD45r7iZXGWVBt3KQFQ7BPC6
biDNeMPeEIfyfAex40BjbCYZX/+X7grrQd8A7Mlpa6oWiUILs8IHMzMHkSpbLWR1
Aw1C+w2L1tdZ25z3rja18N3uYc5lThtOkK5xOCapWC095Q1BLErbObMWniH6d+a8
TiXy6ypfCTOgTbeKkdpvdekqttZpytpAQDMSQP0fkukyNWxDlHYVPT+rJuNEsQAc
VHNOVi/aPLWkTUeo7uPHCzEx1kXLGlTYqz9+iVO3F93bPTV52u7EBC80xfwjMK9B
1RAKVtut8pPfmd28UjrhXcuvTxpCK0sAjX2hsQ+U0JZC0qA3TmnaAHTmBfuV5UBM
e319rmzDnxz3HAx7qFV1vY5/nsmPRHpu/cFgiSYVj969MCRQ7426m5AARNOg2a2O
mJ7kqEXHlEup/gk7bHZtvV8F9FmLG2EUuT4G0zmf+BamS4VGTdKtxaoaFMDOxKKv
8ewclQTosujlWRXhGb7j3IXAT2BoErFrb54XSOC3CmsPa4qcIr4pBdX7bd3HN9Pe
CzQ72htsI3IWN9PDwG3VDxpHwOLCvRDKUjPSJCPD+sJIxK9mLAqwxp2llDfQWAET
BTARQxzfg5if4n6ulkPQRlejpjn+SlzsL+FHd++hSm9ft/sl2pk/bJxVYlr1MJB2
ogdHHTAq1yfwNvfj+SM/cwk/BOLV/5FCH8hLRMtxGYl+yh18KlNoK73xzS1t5Itf
flXdl9spbMtWuHScYm/nbRdzAwM/NymR3R3fT2UgLMUVqngLMFhO38EMT3Jdglrr
bNyxWWoIbHqvwgUFU5AQOhUp5EjHe1z23qcScOa1bR0ytIz1TURMMdJuvRGTwdNd
DNehqbSuFJEjHA/gNBSJnxhuAE5CVzgTjVnwA4U8eGVT1kQtEvRHp5WAYFiB1bkr
4heiFwXJ0Nta65+M8l/tD6bDl2uDM/y72z4jYrPGUog0qMZ2vAjqkmWH+1Q8f8AN
7Lbq/P36rTQtVHdMVkToVgc3jCa8kzoLKP0TgTSyrszLlstjAaNlG87IbY3k7OSb
1oz1eucQQsHkCE1hDfGtOA+uVsGRXWe2q4t/XmdSj41lqiz5vufq8P5oniY/KwyE
KVjNyHFD+XXRH8rYray5PaIBQo77B4nulp93xKXOPGBjr5MhDVK97+EwjuQgYVPe
BueN6LTYAmRdKZv8Cf29wT0wktcL7Q6x0WQhQ58nm00UF2HSUCe7QDs6/zlZu2Ol
yGkmqn6UgKvrZFZJ6uF8SA6WMDDiGzZYvFYp4TIFMFFOBGEJGoj6S5sBbuNnbhzp
maxIQuZgc83H+AEP/qRDPdtpYrVN5UPToTV+xPM6F9a78mZllD6QEHsC4sY3VmB6
CLj034BT3WBFJv99+7P0Px4sk7yx8wy/djKMQzBrgAFJRn7toOuFXC7nWV4E/cKC
cZhKpFFKh+233E/0ZE/5iHwit5lZS23u1opP7gRlPoXtAxEghE5Jb3nEK769vcX6
ZHSl/NS4vIfbH+XY2rdTdTDKj/LrwuFg7ldWB5OXtnCenlTfzM7XA1g8foKjs9Zg
kfIjYAcevrA5cYOJY0kfiA1yDg+Rw7VCkq3ets97DmIYtSIkEUakkY8ZpFh77k1E
gLJe0D6Ai/pTUlTR2tmKPYiL/fc7xTyUMRfHQzpuzWUB7iRmGdfBsmfeUQb4C/N3
huwHLP2G8H4xQz5aQKTvxh+ramBy3rg3pYx9Qrp/XnGbumMIWkRUilzIx3KD75sf
g15CoWd4+Qa59riRlAbruN8N+HsLcFd91VJLiDAcuxHVVHzBqIcS+xsU6pxDs0hn
YtT/9B5b18Dk0f0J1sh1ZKHFuXp/DuOlkhaZteM2dPYI+Wu1qGnd62ts3Yf34NeG
5ic1Dx2CGfaZr9Xa5exnJtfLix+9y+VoW8TgUE6uWUy4nZXli+PLg2IbGjDXUFCz
J3njr+LA7jLWQ9O+wzi3rKwSZSjqbxjwEQoU+FESNALNWcm8NusxfvbRu46nOKW7
Oq97swnecwtpt4SWVWEV7Uwbc4L3egAoXZzqvVOPAei2rz34ekOT5dOQ66FTdOPf
ORTt5PfpbKWw1hl2qNIulH3WgyDCxkrayq5o95AZKTdAbyCFKSN7kUUJEFoj10HC
qa8+wZqAd5HnNKTJYFphkpMz8VkpAwHxrM7jTKiwHq9E3YSVB0mriNGgqgWUr8t3
dkQLaL9KQDp6n/YTPjpvKj4VlZP93OvStzX750E8t/jvQ4uvmenZNiqyDBBxfTh8
ivq+T+3lIaCyQHP2rHo/4ysqVR/ryc6UdqLZNzoVKclLEoSFNnMJfX6SlVRqK37l
bxe3RbOyM+87bAQVuDao//lOpPPu4TVR/27AivV1Uz8GQUchrSjlRXUgPdmyrneK
dK6EAaM79+Kh4uBWV1pQXzjAexe1vQApoyJ6Wh8CviQh1FrUB/LGoBmzhSoWUKSn
vPbfdjXncrmRlLmG4cmH6xIRR28tY/fPTqdyegFnycnZ5qkkOJFM/AbxAL/uF7WS
GsP5N0DdemqOBwjYGbyex4PAmLOViOh+agpwUAtdrn/9f5I3oJDVeWRFI4kKxuCG
hFVzWa93RTjhiHgKJVzV5Wy3ACN0mH2g1OZfLf+TJqz6KtHqkCwSMTVifQVz2yoy
be+pSbBTyqQEzgNLk6jrQu0L/bi5+xFUicS6IqSCy/qMIi6WHwNWsZMzBmkUteYY
me8jAVzReemFGUUCmVygfM1BJQBOZVTDnAu5ETLuHpFUaSGNxCktKrJCVDFIIil+
JljC1STYM4/qT73s4+tMvoqBQDXLmWiUEmo1WyMOv5ge0NG80203qX4NG1BRElej
Hygev5obD91LeuRgUFqX8onQHtDxb8tdssIa+X+u55n3r0OmKW2cZRfUML+qPEwE
Vp1L8Xw9uK32LTx070W92B8Pro72y4ToO/Pl8Ny+6Ef7GNj5O+5Z4/j5hZJfDZcM
lV1uxLvIwJxgD9IUBdsZC4HN+I3ru7u6GfjA1D6+VhWZJ+YgRBjKh0H3OTgCZKrg
HHoZz50oxCoegiGziRv3ysSVjDKxtolT9v6Uwj66upnInaUkyEz5/GalLwt1EXLq
97VGuyG8oFSRqc5eEY/W88osZFONAJvvC9v0YpSJJNgK9nX0JdPiDls5T2zjqIvQ
XTc8iIfIFhUpuWhJmJ1XfMmvUCNf+Er2TSuS0Q2Bu43ftsEv7c+IkQL29C7aeQNa
Eiw0K2SIx27R2XKXoxwLrRgr4+5iutTyEC/gY5n/fEq7HqABTAFxfUC4775Ca/QQ
nnUMoDLW8jMQP26WZfzGwMQIuGD7qzNYH7xOQF6mEdqnW2m0LXwJkPATpuVcylgv
59J8fiuYTgGe6FnCsqgnjn1S4Xk2PRWmS3fm1Jg6AfoLKYnnzMndo+5u3aPtaLsJ
pkJ+/TzqHsG9nZ7f/AGQtwkODm4/3IBoPb1apIegiIfxtl6wgyBkftKtFpbZjvEx
9HXjNof5atw+euy1WhCjSD/3EAk7LW6lwyujptv2SKhvZDMsLWvRViMFa5cjHlZu
KhshJvdBttvBcrhdD1izXv5OwTuD9peT+aVm1cl6rW/+/yslqGnTWPleUq6n/vrU
D4hIWBN1p2Nl1oQJLDwjT6R1y5qmZiRSEKFCEv6z+XUD9fEImC6jAjTfjD38lBOY
lL0ilS7xBrYHXFtBnIIhiRmHm3/BOW1nUyqwMw9Tp12lJiK1y/DjWFfrArgajskb
x+u6lWavSzb7M7jJHdqBYT/DnsrtDng3g2Qacy2XDV2ZZlSWvrRBc7hDlIw7NHsw
OzGfx0hXwPY90pNAPfXKcybpdvK1nTLo5l37P4OPYAMtpw6M21e25gXFV1eHuagU
rwtvrZhTn3QT7TqGL6j5909zQmxIfGGvaymtJJ62oObHQKXPD6QQiV+jki5mULU1
H5kytQzAknDssBjiF7E/sVcT1jRvl0zUH6QXlCuaCWUn0IXwxz2T0exrZXSNmi6U
b4IgTOQ8NVHgdyGPEselPGyx0BxxwEYwYSa6HzY4xlnCfFsgExSsCVBf9FaFFVMZ
/w2773jeSRzHL69gLEHrZ2lJ+g2ey4Cqn0Io5Lz4zR9RGSMQPCfdbWX5KqqR1F6K
j0bCl/CK6gsrk3M0HFg22629/4bZKOn2Ir2iaoQvMqtEP8AJM+mWxAoHnCPU5qUb
WDZ2JDOFFto/TQamiFDNYjqRPsW6GTKOxqcYdzLiTPy9Hrpeu3l7YB7mURyJw7pc
D+VZlHxbxROCOjSKk7TQbgol9P/CoQtZBg4/BkglnsfuzcYyTpbnMQRdt6t7na0N
9I0FGWi8q0jo3vqR5AAiwjZ9Xn+Q2Mc7rSkwn5Gn8hnjBjup2dkWdLhcfzSXd51u
ioG8nq6vrzXCnYI3YwzJqWf5aTqrDvs2tMy7ZOT9aGSN/HaocRCBuUAmpRiWhptJ
CcK9whlmyblx7ykI0C5ROdD0lQ69E5Yt8Im9dMEhdt+vT0gVWkbGKJI90W5h3b8M
wOM8LI4QLZxHiDS/DC41UOhmPwqgoxlvogTPwVLfhstwL9+0R97Zs5y75A6F0R4m
C4RDptLH+RmhApw6VoTZiReKS6Fur6V+7tmzlFrDZiAJB/cAwWgTfwpsK++tRTsV
ZBCa34V+K+DHva/8oTg6j+bxq5b6iHe+lAapHvRZ4AFANig1rhupqo059sywZGr7
naKzUIYrNhHbA4wJvRuJ0bfMy3ojuIKwh4VIJYTme4885Am9h7ZrIGOGCVvass5e
M1Kd8m7phIg96NYnsQyE0KhQeH9Ap/wGJmIEZ3424/IRzWWF9RqS+UyGKrQkz53t
Ootupp8lCk0YqreNKTzRDCupNmvFksJyq+KsjvvlefDUGpGs2MMPQazamkYmh2ED
W1d/Us1n3efpibgw7gjlpYjofZs1w0SujQtG2p/lfKYaXxJRB/RLMoFZlMo20Nxi
t5KJRG75w8RyxQyfyRvo3N9JuoCsnjhN7QItfATsNbTYQVBavTXh4jnJrB+QlCxT
kaNCm0PBeiuY1jsQG3QlIJrpn4UNoK0+uMnThlKMcEXehlmvcia3C6YE0rxkeRgJ
j9+JHZ7a4xdes7XZedvZ4o3aOblD05MzrCtSmceRoOSAkqRvv012oBFJI/WoO6SG
Jx5vA7WQ2kYd+prsaM1symbU8DTie4N2FIlOcndCNPt7lElT1qCbLFnuk5dTVx9k
rFO/5FU6phsg7Z5Dvzz4KBrLIA9TUmLOjFAms/4NjJqG+1GCTtfwtz+o9briOghV
w3f9rykxJ2zY4YPEhmlYYfG4OkMmnF5FL0SKPFKiuKN4b5f1PDSgwatF7xlrHF9t
kBNuLmtzIRqM5AOuMoZN9vyPWEYuRqBec+1Kj+1r6mbeTtgBuvfpnVpydiKt2wtn
PWJsYx+VnQvgq+ilUo2ePfBPMdeMK6gkRFuP4Th96QXLY5gDAjtVOJAhLc0rwXz7
UdrB8DSMsvJPXYU2xO3j+zJ5FjV72nUO/Ct8Ce38YZwuL6Ybss21ImprYd2fOwc2
ncAEVy6ggfyXI3EUXUqsEfQdEaT3vHBNXjsCWkWICNqX0Xt+igthhm9KjArcUuQf
wTwhWLBQe7sJuYGSKB8K6Z4d4fimlEorXyPCS4qnEVTI85GWzqlX9YcH/3KUfFk/
suFwl8bLkrjeNUwqUCODUtkEO4QterCZzpablyfezw95PLss6icsRz7C+GqZCkQf
tSi09qN/w+gwVtYv/LiIuBAPcET7y+x6Br+9+POOhTSueHks9S32hYFTXrHu7MUD
RuRo+THxf5Rdv5qXUUzc8fzib7jxb8FvlNzZIknrmQlRoUqkcoe+CCA4N421JwHA
eM+Shr7GfEjd9JpipsM1bEYDShVcRa6RhtlXYoUV65DUIbYHQC4BGD6CvaLH05AD
o+JKB92QHgBswoMMj48nWTapVbH629+4mc3SbGimVRxBljF0UsCLR9JPFPOY/zrY
EZrvMcZjdaLAW3ZLnu5YpGUXrUdEh8LU66iXmbHdg9sviuSOXIzcyVydEgXerBkm
nVZeai3kjdJxkRyNR81bFI6dgBigBLbiu92NYrMufv9Pk/duz2AuhYRvPjlBb6me
/G3w5rBH0SCLfEQWCZWfdJO1m1fxchsZpooWn9f54TSc2WcaVRRTSmLdEbbehxq9
HII+FwlN/ZoVj/RhJ0mYHxDx4J2paAeUihsXyMria2ysx/2QiYMNm2z5fAJtwXjm
s2rjE2+aHOlmNMmyLnhLHsBHZC01GU+6oRE27+321q0K3Zk65M0dyEpiqcS3Sky3
m+mpr5pbpLQG/p2JFF58HTaFgjPxu+JyqEZ1q1jM2+X4ebK+sFa+aJLgD1fMBA5d
EWlqjy5KzM2G6y4cRUUnxoxhifdYQH6oHrEi0U0aCLQcDQb0KfGZHetQs29ROsC0
vNAY4TEqjb3yCL88rwMZ8BcUvflimxfcY16UxivIu3oGBRvQfeU6GQBrUpkSi19G
6KTx8SUM9h6xTH/W/sb0KeEXmayEJfFvxmnAjCGuOr9va24Qk05cgH478/FyRl1k
Poeoi+cVxWkxhUwvdZ/0/wJIIPE6jzJBcvfZUPsOLlWYdy/mnJq9bNcaP6RJEoEO
eoaUFKe3ZmvJ4LMH95T+2vTgtE446jv+jmh3Kd1UzM6AU9b95SsQq1cE3cWv2h+l
xjmqOTm5rb8qz73g2ThGkXbQir7JzmULmmDtgR1WkILzetbv4F+DsMWFtvrU2qIt
dQgIT+bZvZtI1MaG5hEwt6ICSucF8QG7Qft5hQIQrCH9MEM4PvN3jo+5nEjFkJrc
ZrBRWfWUBwrxySM5tuJlo1zgXrMRQGlLgP8Hq/uBeWF5pN2iBtWq6UaR5NnL1D5C
J5rrgYbVNjEKed0p+WOMbmZMTHEEwiQTkp80U+zRNdSA0OVdUNQo1TjMhDnwX1PC
mcug3Yx8+2aenm+GBWz2C0jVYqh4y9V8vwi5vI5eMwsFnBTFw9duM2d93sjcrPVe
4w96yiREdFSfIDLN276PvPUbIzK1hHwGNp7wnQ6ifSGXPO2UJqEFxnf6TzliJWil
XT70cC0OgPbLfBaFAXtyftnJ55a9/jHurO/rI7hTKMNclktxV/m05gNEant9v8LM
E1eqdhqFTAvFKVj1ru/9AzRRkemo+EKI9fnr8bkliyxNsgR3j5TvoUkpvTRBj3a5
pli4JUZgjP809G8xfjP/IllxDOG3gXWLRr0+Zz6lONrozlk1qhHcnnuj8Gt0xp/V
6Kd1KNmY/9Xr5aSVoNCve2Y6jKR4ORCoRk4C2LrHoMODRCevlmNl1o8VW/rFGJjr
2oN1yIHSViXWsuMh6tZ/hNZD0KHr6R8Jocxu8UXDbCIoVL/28spedDK7klomivOX
EzgOJm8LzBJcnVmi43s8GT4o03zWTjvH1uc7UgFQmOyEz6/jjS9ZhyGircXD+JP5
XgZHP2diODP7/dIGJMU267+5+VClv/GuyTMv0TrzQSDbqTnP1am8HDZXW81lLHuY
zPCbB5MDKJlGZ4d2BfNc8oKGdUZ40j/QVmvGaPAAG6fi7hw9RmCR6LkICpNCIoZU
P8scB202hgK8zg4js70bzdgKdcfPOxB0yAQ+f/VeFjC5sfwV9EukFwFsLcu1QZgy
yNDE8BO5QlQScwIFBWkCSlmR/eRRz7413YW8vsmOWxXqN+eCagELnrMZ6yQEVHjf
3tSY8feie1webM2goF6nsr/7ohsv7NZn5r4jNT/PO07jYyweGV7WO5FZO76vtR1D
eX8+zqFRmgqMN41B3bErIE+hB9ivQtVfMZXTO3HYeFUSQ15ceHKkDuUnZEyseVsJ
hTTJnMc0a48ZoXZnRBiL5R7VxdEnObLs2xWIjlu8OtoCSW2G/ISQNWDqG9A5peds
1l4dmCdVvkvvu5sLe3HYH3JmnhMOKye1l8gRYh3e71eUZjunoZ8TXvhduMN8JKre
BuU3PrD22FgrribqoPZmR7TnCfwUinIM4+uL1+R3o+0JEiOijff6C1gcwB7kvC2k
TytFd8uX+DHbINJ+pxdHi0u1D1B29QR3dry1ODNGMwc61gRl5HeKx6wubwAH+2V7
QmJpqf/jmlMBRultiKkLXGYEOD1EMI4WmCJVCnV2q4zqP63khC1wq6hMHvZyyZdF
MtRgUnVR4282sz82B5sLAPKmCG0LnPDwyZsi2Zcd5j2MHmHj1zR5IufT3vnW5Aih
e/jNYvP+Z4+lF/odk3B7fy+Os7wQ2xcGwgORmwQjD63ZfcEUU7f2fG7n9VW/43se
Nb11XJ/Wl4PtUasvWoNO9PK9sRRY9Dt2KPaMdkjj+ZIv1IyKe+tXOIa7GIHYtb0O
vV6UbtNW5P5jvXMQ61nOWSy5NXIlvDd3OGpHzMI6uLRBshdoW90yBD+nZ3tOTsVp
Vv3ktOcugLsEIS/ykwxgiafR2HEXd1qovoMaS4lrCw3kQXdD+Ky6uVYxe3BGoCvP
pSX6bEZyAeQsz688bGsFN36y8K8XK6io0ViNd90ij7QLqjBumCOzOUWh8m7ldPrw
2qXmrjyXaMcLgTLsakgtL81dbOpVp3G9tAU15EYTBTJ5cR75vYwybDBJZyrs8Vd5
yqCoq8f24DbA7F1qqLM9vLHR2qG6Jmh8swm22Lk7BnOsJbT0p1Jrvm0Y65LPMMQH
xPax+sKrjS+ahu8UhAe8F9MjCJyDhwu1Pg9fklUsKH5ERXMENZ5NFjin8/xWWqQu
K9ZIHh2NDYLJ1FP+Psq1LL3J0oTpGOwJmQ3JgUM5FEmU4E920V1hL+pz92gdfjrL
Xav5ehjkCqN8eqi0d3zvXjRsFgUgd5L37ONKwDZecjOqCUEPv7ZSMFMJPoW/+l0D
Mut039S4PCYF2f5sMmiO0mYH20cCsrmUBc8/oSVhnled+CcrNbaFsRnMm/sPFvEt
2KJ+HDYoWhKERi2HWbmDzeJqzbVlFAiBBIqYB0K/M4OdGS5Vl5xd1FcT/D41cXCU
dC9Pzdbc3/lmqMQuyXItWlbOJuslYmekjmjNnayxSsRmfqWZW1Pu7QWXwy1Mj1+b
kP3ZTRoGmK0FHTUEYMQ6JdOVQKwrFleHHMtrwW2pM7bfHsNVYVSZzwuAeZvlRM/w
yb4cRF/DwPFqxL0uFjVwT7BDeMBhJo90QIvVwJ9sjEZgx3V3OU66rLEYjOHoZZFt
+c1+beAa/zq7/v3E7oibEGo+GBLCRKSA8+H6OTWK+J6wOBj128V4mKclsxkebrNZ
oNd5JgKZlGqXuPTBafe3NSwJOt6YddV/hxs7neE9C57lKa+qUPIvW0SUp+TSbwu7
nsEjzb77JRScd/em9WxvAKA2gNHXl7U42UN8srQw+NeHkeQub7qFozqrv9fRUx5R
eC3lQNJ0wiH9dhxvQu2ShPPXU7JduhuPSBHQ07U9UobMkv6TDt9J2YWoOUOFS6bT
VDK7hMiBJ234PoDN/KnGlB7j9d1u8lcqxG0h75xdhpTnjjtUsIYabokULyVC3NBd
2HN475ZIs1JVoS++lVluXdyWlqEUe7K5/ro2MXVOMN3g+CiV+zcojOZYcg7S45YQ
Jc7vZIC9QfgHGeUO8FnovISDoPsrlJfozFXmQkWLy8QK+bGmaL84Cq7vS87iIyRu
r2iAwEBDyS0XCrEmmldcrpk3OLv5GG/JAPlifvnteuB3a8zy3NEh0grqf6GBbXxh
QNgwnS3uR29o0Cp+vH4zYSmLA36Lg/xKDTD7AfnSTAcebTJu5X9f840Q1zzYlE7N
3TPrHZRGQiPvdzNEPmBJV10YRoWFRv5dc5RkvLbLchiiYHfIge9DG+YJ40Ux25SW
tqCvFlDmyqqTB1YY080tALdE4W2DSAu1sOgmITk1IXemu/e9+A2XFHWekW2gkXaB
CL2XPKmVJtIWn52+G1+wCWdXDfKjWUPEYRPx6NWdMOk35yLFukk2+YKxYPr+OvbV
6qXLZi8aZ2PDSkAhzttdLqQMBMhjDsKb9bfkfCio/7kvuR7uXQo0Oa+TnmBnW+Iv
zoZkdxKq7nGAQdx6yimE+w89gbvBt4ZZlUSe2GaEvu2+pqr54fJPm3EcZeDBHMWd
iuW7NZceOQcnsJvLN9YiPV9gUtxbR/dku45V5azhDFfWCVgurd1bKsmpZGc0etbC
izXg5ujgSh/hib7wtUooNeNjx5mxgPyF9FJxy9PaFFcsjLDirgDTPkaBzUlqA0fe
ka8ibxicgDBneGXIgvWa7FBPzcpedlWXNxuLEd0eaO6ZFKL/Z4S2u8MXxzecTyME
IJBTfvlIAphDWqznqDLXVot9NpJFVzFdwtx/cDIZ4bYuEqBPQtnMHNUoNIqh/p8F
XypyVTduvpbjLP0oEBTT7nxwh+Hz7m57X8oX7Vv9ty2mWTrspTq/4PEXCOrv8gkC
hB8mLS6RLBQUMgQxOkz8zA==
--pragma protect end_data_block
--pragma protect digest_block
hDEkV9177072CsqwotaoUkyeWNM=
--pragma protect end_digest_block
--pragma protect end_protected
