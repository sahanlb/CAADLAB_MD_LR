-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vwJ2PJxaA8faRmmqX3oWOSxaJydbbm4cE6IiyADimf1R0UdDOrMj9Fci8Gu4tmxVIOiVxd6O8ZQX
EAZOEwckqgW9oBphONuUX9BP1RP4J4uGlrkAnG35VmUjHcd0zimsKXs+YJvtQm5H6RAt/W32Z+22
GwmTQHo7x466jtags9/jcqb6Y+ZNrqtD8FFN6WRiRRJSntqGmRAD1EqZfu3eRgMc38eA+mfTRV4X
hPvct44SxCJJCv8MuTfVGQaLIqRibRRz2CRrb08RuXDq9i4qNvDLIdPM3y7vr4gSs1Nz3kCwqbKg
u0cYWDaTTBs7aRdWNIJWMc0hs9QJn6vNdd4/tg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5168)
`protect data_block
nyLONcJvO9DFNT+Ex+G0vfRBFLdBe5OqrHqhjsWgwLROPZX5zLj0+U8KkJG9ipRVi2D6iS1fY+4W
/7WuDGpCPK1HhUYWne8VSquiC/tHgeWtdKWSRA+OoEJJ6QF96eZv+0oIOQxzVQcfxZPGgbvF7O0V
oodFFCAF4tnv+0BhhMuMaJC3/TWkDD19/IrDfOi327OQWmBSFPmGJ9wUkZptf93VaYKDz2vIviJR
DI/bbxr3eIseLBky/Ap+cSpzrD/h3FjLqg3jN5bh+jnmRz5iRYFBmK24wY6GUKGMFXpWxjJg3aJJ
S5nLp9ghGaOicFms6zXBBAHp/TRTwVthzCgZiqATHO/saNXNuHHZ1ejm8wgXQWnrbSGAdru++hxi
sDthRSFv9xrAOgymipqIz1SfvUzRdrk0P0C8dxK30RGCi/obNobM7Kyezlule3iUQfeWNi4HNbfV
5/vcbyU0u7Tf6zTNyL1G+28MdMSWoKFLwKXemVAB9GBoSpBM3Xbq5ATXsrvLcd63pG3j472nrDe2
VVmkGALwAmwXCopYEbFsMbSS8lMjgfe484f1FpqJzIqugDRsriPdkv48DSONgapha5AL0HAG/41D
KG7QSy+MGrNZIpiJKbMg0T1tdV4yDml16Ozw8H8YraypjJDqQ6916AHAxZkYdI3erf4Ekg0z3bNV
2RekEXs0qD43jcdOiT4jKptMlyWBtMcLZKO4GOWx0GU8Bazgx0922kkQvLLvLTA3RroX/fyDU1Ln
Qw3qGyO2zo68iAhw9m+QBPQN5xn74370SgwnjQrwCI8R6GTImw7Xw8vzzLPPV2nvTTlJcC4xr1S/
bFy8iuG2eKCWRZWTZo+pyCvYQd70Mzu06dSJ9chJWq845yNQkzpNE7tpB2TLOKfrglwGR3EiaV3O
fRK8454M64ClXncdrg0QUtX7svoLqtGyuiHzKkPSYZCZfWbHEiY9U3W49fHiU3VQV48RbFFOzYeT
gApqLTfh9UBIxUb6wvcWeYjc0RXwjuIGOlKg/qprcUdHnheS7EPcBl2Xvaj+OMARkrdH9L0SXWjQ
ivBOUUnKwt3RhsbP+Q88w1DG5w5GoK0c5HX3855uAvEI5xzGFUvBEeE6iBEXQcA8Bd/BT6ieXxvh
AkMSG9BURgxLn+x5i1llv5pPEr2igCO2YAIte6GgnhaynvOL29DbWU3Z23X1BHKGkYm3eP2u8LYX
aDe1bYgQzkZPj45ii9zShAaVWI/BCXYy00SE46F0f4d5NSYGllfKdmEUMp8l9kIYRNxuT6i5yOf9
Q4yoCFl/B81IK1iCpXXc5CrAgr7vhb8g5sC3lJ+lOiXvmUozMZteOjXcQioHxZ13CzmbHiMOrh6i
2dztVSeWmq6Y0gpxzr69bN8aX/GpFGPmg+A6igXnB6V2+pl/3XpSbjx1eLP8/ZLPRfXmQWhLYwlu
RBXrKY0Rlr6iva6DZ49RIHDb3Ao2o/KF/np68J9X7gugJ9XfHvcAxyJdv3h2XoEaYjTGu74GeTcc
FX3D1jLMAsCq/6qlGC+8gVkCKI7q7j/VK2AUQRCC38ev3aaZUDi0XUDKFx/S8Sf78UxVhrxzgn8A
gPXUzNspZs3wX0vFamoc4H/7OH2F8B3cyJJ5EwcTxtUQ3KuB624dSGaEOVv5t+TTQ2dDfjLpKQsC
A9nb1tY33S1NIWNkkFiBRWn9iMRXM+VGVLBhE9UTMkQasCt/Rnv9N3k+v/QavUmYWN+0f0I1Ilw5
rSZylUP21X8oqH13mwfcG9eGrtEuxHtv0ZFi6bl/AryO64CQZvQ9sC/RzuSi7zowjmbVvpMX/oPb
Z9mJVGt+u1n4f9Gn4GYvHFHpudfyokNb6Q6VqkKNbAn0JZVClGTgsMJNWIwECevO5bmaTxxrZyef
Y/gCS1JD6xTjQsBSanwsfBB6w8sM30M29nWiV2a1JTT5ASoMa1G+15Hp+GqqEJKpv3ZO9sxw6940
mAxTIvaaagYZS76TIiF/+jcB13QSxcD8flowISUWmYgL4Z8if13H/NQNrMxxbMx4C7dKpKOCgpOn
KzPRhayipkGEQHbMPwlHu+0LXm28asMvNsEWoZOIgi7ej4lvlci1DP+okSPFhVfQ3cDJMZietsqw
1uYGLAT4QI1HYqIxCSFUOxJRoH2FLjlSGrcqOyiVbeWq9A1lojy2Tn/M49JWHfskb656JsBlQ78F
KkUejNyYus3dz0q4hQGdmXZlsPaJsbLVcwypMQQYEOPkoiv13QJ098ME2mLllxbYwvBBuVNitIFZ
4eNUEJTAJBC3OZc0S3HDs9OPRUyJ3xyywPHiZpaEC9TPW8l+Yg7/KBC5OzdWTZJHabKej7zO7bEv
SW3l27Nead9xBMpQ7wIY8r2Bbub5cOwp8+HJZHKUxlUo0ArT4yQOWgzcrXti45OeMObvksfbUubK
llF10MV2PQJy3UTmOlnyBePzEgEDZwlVDAaI6ps1sxrolYlNGhfwfHIRol97NY63k1pxbnJEx/Cq
SXOGl84YiVq+vEDW703vOrEUayJFMOtQ86TFlquC8hps43DZ1SDosgivkAmCqvrH1zG1lctbtENu
O/E7NaGRkzkgjKtnbbTx5lEOjJVqnj06cX6UqF/Vttw9fcQp9HaDPS1RTbaGu6nt7WakE2PsmqSk
/qss7cPUb7daG6bPjQ4i2nM/KIXi40P6v/lVOW+bj5cp8eJspZ4aVpc+uia+yN4hyg0iaA0npwnr
8ekpTzfU4+SEyjsNtwvjlS1PiQrFzBunZXIbK7r5ugeOGh0zvG73yh9k5bIA4WwkIJpO1nfc7XJD
7iBWpI6q+4JtnozrQlbeQg6vINou9DXO675M63yj6OvMndqTc45h1G4aEUtO2C0Mjg0FXlign7ex
YmbBI+JnmbX0d0/vqhStXeN/5wfAUEea7LV/niHj+HixrfUl50WA3jSEWXiiNMUa3qYfn7HbQh6D
ZTtbnwNP27/7VI+xi6LqgnXeRIXXXhQg24SQyLiXtheTPIveQ6YpM35Ez2VdDH2+9rDXRNyYI7GZ
MhQ/G4C/85ntWnJY9A7sCuADc1xP+pVjfmPN2BAdng39pgMgFjhyETjz2n8IgOupSZaqhAnVamTy
IB/8KwzpkP2zutW+hXos0WbBi9jVLEezne/6uHvmwEm1D8LQAsFs3icQYUliJJIH31u3zA0DGDxZ
wJKwr6Dp8GeoKTxZqttXRkjIsoH7KiCP1WJQ6/nwzMkWMFAmZ2opxjCimE2JbBbKWUtX+i1hmIwT
dDW0Y1Vv9I1EFSqouDSKoSNkaQFRuMtaIRdsrPEWEnxuqbLqlCecEURh8a63qQzM7ERQaohS6Kz8
j1l3+7HE0ONlFxqpOkniHF7upXfI646dP0LB4T/HaXHXu5dFGZfgptMi0xphoknI6x//4I6HzqM6
2UZyZ/E3Ri5wOvMSGMI7nZgonEaIgNqBu6AJ/CPJtSa3w+fHRc9eTDmwGumFlTol7h2JX330m+Ko
OXqIywUydlHplyYYKhZdEucg/E2vmf0rs9AjCec8JjPHjjuZ2uMFnqfHuUnQZDzrR8bQLyrmbID+
f90uLbA4A8K+g/2oRkUEfQTf91y4+Dx9lCfbRs16dR2Z0WMuRWf5m2f8fLXzTjPmvn0pcHaXsJ1j
ggo+j/h54xbHMPFC7zC14R1ugG8b5LbHpsmp3U8oNes5ZgAJnytK/Qj8gqQQdwKokdt9YZg+zpIa
kN8VV2TpOeiQKY/50XJnfEdDtjgWdES89t73hp/O2LIE9VGBz+Hn8HguxEVaXJkOx8DgIgzj7vTY
ixpxv+pL4ZkDbjZMXi3eGKhtzbvpnt86NrGFjhgP3S4eUwj21lPq6wAaYRQkKpgDgvKHexfjLR5H
e/aC6SuswJM+j7IBtfY2Ap/YzG8P2/VAIBSimYd4iORE6WSAYHXgH6GMDwxDwVm54bNn2lDZteux
a5J8dUrIHJ6DM4RQc8odDHnP1OCcJy62yfIx4zakkMIBRb/KRmhqcKkDZ3N9gwwMh8KQHaevLWIP
LQBJ7Co2cPGLTRqzhVBNbWaBuyNpVi4mRFMue9yFUHP/amNDSGKSPw9kB47FgyL/mh8SYe6obyG0
sFhyUhMXXzny6lZaaR0p6R5Kl8MFpnBMScM8C/LNPWUGdvL7UDyVqvsDasCEGErMIc7x3a5uR/SD
0Yq+RRi3NO5tmW4IMNUYk9nBu++n4QUh6XsNVN6XVgzOTT41TSj0S4IklHMia48bG8QtUZk71DoS
3gRn1+UJBaBVQ7XcpVeFNWARb14hCfEapSJUvP5orLA4RawUMZRJE1mClV/DbfRH83700BU/NFBl
+LBNVYY5c3wWqRhuh76LKgN0fBR/Ks2o/e9gpmdqiLtZPdYHg6jHJg20yJAzyz7Fw67o6clWt9+F
8jaTYwFRPL5P5xqSp42GfMMYTEhpcXIPzwLgQHs0CgsYdqZkWWwHyvuF+oPioXtMebKICGb3Ih99
5tCxk5VdSnEPv0Mb6e6yNDxIMhw/7EXvapjoQS8tIDNlBtPnm4hicfz3QcTtu6IEnKdP3Lx0VAjM
mtkZl9beAFzufzB2f7nlGWnBDO54t/iJ1lwcAJ7xolxO7sBbvELnbAaEU+3mexZfAMJ3uaVAZ0dd
Ccxv7kpi35PugZzikQ+vxX2DM6rSTI5m1Nsm739U8D5Hr6M4Ydnc89TiwY1GSaIkmPRD+5MunjAa
f5d4ZJCrAQKEervmydXw2c6lxzRfqSVEAfmL7nBxoeCLCSjTVW7hHD5lJ1IPqzhCi6zpxJo992fP
ADfbWBOqPFcOtRf+eSaWyCw4TUfoG1vuwU4mxWkizwrVKn1CfEkDZQRtkYnAo106ePue4x1T10RJ
CM1BdVedTJttyZKL1U9APcXelIrv/eH1Si/Xrultqima5pg3yJhQbcBEg606qq7QFGcnSdijHyFk
VQQhVdkgO5/eo1DIu25YrDS3Y824F+u75m2r+r569ygxK9DJNcaFzX2faJp7O65pMoVFnW6MS7wj
ylKvkHJYIfJCqgXBSBvW2n1Txz7FBVx7+dqQjPKCGMje9VadflhhD2ErZUJnn0slJXv1TpkmVeyA
RJ2QTtGXtLgUhsPhF8z9m2sRMIJa0a4vTEWjTCAOG5/LTtefidos19wVk1DsksHvuANpmIJNCVYC
poCpJ/Jls8EXO6DjSGZZACLfOKFjAy8UiK4Cbj1wtTogsFSQmHXeV+rfcJ+K/Ul0Fxh3agWkH8dM
9eE3KZCNv7QsEIprsO4nXBakw3oEZxTiCAOnHVVcf1wgMI/0EX9h9+ogiTVZZsdcQ6RITlKwBm1J
tlxtkKDKn6M6PkRHilLFj35cnPUtmCLoVNeANOQ2csUfoXrU1DeWBbW3TwSA60t0rnqjctqD+q6W
B/BQ4/Hxde3Wa2mhNJ+a0aV94L903SytlXaaQ5MX6Sg82ySA4fmhsY26psRvAFJbWiiLqXOoMtIy
RVt/A7r6L0aatyp/C070zH6y9gHv/dwjppWM7TMPvkqmsGkoWxeD8C4HB+Ij2H5A5+Vx49Dmc9Jb
RGEsbss/PdtaiVOMewlWzEvNjhNP2O7mI8rzwKtKmkSYPMvIKcm/iLrU0jmTPf2ZSsemGNrkrefg
0eVsiNNFmRfEsdo1r1nKbIu+bx1KxmDvLJocUDpfpoG1s8EkOVdF5DLNVQjuzRftXxh0pXfoxeSQ
/UqGErsZMQpuA9GNMKj12fpJdbxe2EnMV6QOxjyElun3djW1wbOOB2cbH43JMtYfAkfSZJKYUWTy
WQN5PEOVotjmVS6WkZSI/V0m9IKAKOHM4uVoVX2DgxpzPPhx2Cc8DuGUnFO0bfBgsAcLU5cURE1T
btYF6gVdum0lDyTmr0ITGJXIxuq39sIh/X8u6o0tmm1397vdZgF19I9vPYn/2ayD2JA3sVgwC4yZ
Qzla/9tJE4Ft42jtWueLAsFewR/w4GDX8u4HgdFQptk6PwZv5QcxmY3+fxN5Kp3qfhxuWPz+aPv8
21zepBwtWHFRfNEZDG/O7heOkXvGWM4NVckw4Y8TpcMZ17GPvi99uRBpesgUM+bkkhPyStwfrRD8
1BWpjFuL2+OJEUcv1GJiUvrfm8PNrGjlfU6+d3fhTL2Y0+ToiCsF2C3j7eBFwsx4uTE/C5Cf2pNT
x2lx31Qt932APXIRD30oXss0kOnrs/bqX2fYmm9ONh6OweTCPxRfMoCBmlAThCfH25PRq4aGzY/V
Ls9r8K8njE6aO860VgG/ICf6ek69RGJ0+PoomvQ1CornKZ7msyPGRptkXM/eyDbYTLKyFDV6qrlq
63uBOlzmpuEqWBGO2f2O7faS9pDqev0bS1Vn3eh8szWU1bSt+56RhnR48VYeaSP6zCfHMwuDOkCp
CD38B8DGlYaGgFF4/BEH5iDfl2UDQN5rp/Hn/w1J4AEByWpa5Do4zzojZhFvB/SPsOMD02TXflUj
oxA79skU6WfsArhutYPd+ydh8aUlhAV02qRSPItZPARDGs4AeiVr6Tk8Te92wNJ2Vqpf2i018ZI+
ZyI44hjRHcYIx2Tlc1JssXICTuC7czklgV9xCHsZb26qhRcgR9Vkj4G1okpMpDlv7hcKaWt4k1y3
ZA0AAriI0DaXHj3M3k1Sj4Jk/wLLjBO6AhVMsDvu9O0Xny8abQE8N/Sb5twoUJuXz4lUGRvbv/ZR
bqGl3znlWG3b+tb9Tolcf3J+Ptu8CAiSq99khVtgxzL2L5Fg2PLnpl2hxr9hpPz9r+E+FymMggJG
cs2Gbfvkq5DgOkH92EUP3AVFfEqfNYbCfV3DawoA65q9vUiY/i6YZcglhcr6fMSEAhwQFtzBTBMY
XQwFM1HFzWzAspk/9dshaaZAqGD5BPTTE7PQihYQmX80gio+RCw=
`protect end_protected
