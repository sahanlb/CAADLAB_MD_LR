-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
PSo81rx3pj288iEdtNr9JYXZY6AG255MYTuypgv0iKOHOuOAqaQZBE4Bc7K842ot
zRH7+xCKUQDgaS7U6aNXKvNnJRUt7GoxaTj90MaREDZbYemY/WKiJZwiCDehzsik
AUoh/sICPdXwktRim39JudEksmzJuNJTipCbtLFN0UB7O7GQPhIleA==
--pragma protect end_key_block
--pragma protect digest_block
nXBkZOELO6/9Vuh8Jj/vk1Ig3tQ=
--pragma protect end_digest_block
--pragma protect data_block
TaaJ0UCHYfp+vMSFfTz/fiybMK3gEWCehjz0cghvwKOCrfOxxHQL40Jg22I4TAp0
xYTlark9MX/YDwRwmt6geABn8X7Q6UsopKG0DSuMRQyURprkx6oUOh2Hgmfk2vke
NKL7zCRQFXVvB52ZVfrOxdShi8XDtLw8xVH0cpNMIbW8hJAYM5KY8dSyAOBIxpGL
HA/od5cAqWYXwrw2edCWiaAUsgPIeUJCV46iUBqqKEueGmQOYxV078nO8u89WPCF
ijJqsgwabDEygm48R7fDzXHRVGb2GpENx140HI9hpR0sLlv1gAOJEHD1eQbHwsT6
R8dxbVYw6VEPfTYOv+fU4EczuGmv81V+OyFXpTYjS+Jl5zIumF0QyKEcM2PhfQJl
6NpBChHl5p+lUsalwLlncNZtakxTBBKaivUg+qaXq1+qpC0XZFWxv+cCTjWKOLqR
S2fUfOpnLKob5cUwFjBYd8NkhmmzTE4xoqcgKRxwVYwwl0865ErsIy/O5UUyGxPa
xbENI2ve9a46lFpDVy0bgvlNu23aniyJW3LgHOnIFtyGqN6kVjWukg65vrhuRXkL
FCtrsKNIci5wh5LWMm0pTGUk+wVIq70hdTWz5tu7/TcDr0Xp8ayJ3IkwIoT5A0Lh
eDyhf70hADvNVj48cjPes4C+gZ6Rili58ptppZ/FM0RCL/2Wu1Up/zBH9i56Qtx4
7F+6MgsNEGVR2TastCqRVzEEG+Uf28/yzclNQV0sBSvMOV2Z4ZrXAgMJgWmohZ3n
86Q0sGP6KELhtzueXwNhYqnTdPAsw0JDp3YL32lTWwuk2WW+ewcMQplCRULRK01h
9KFhtpQqmUG+PoAtdzbeUkL1B8ZkZB6yyJRxAzuoF8HfXDwDprzKrjS8OHoTqGW0
I9KrZjFA+mZZDdOuePeN65NCmVQXJF1NwNUm2pbi7ltp8Yy1O+b0JUoagONykE/t
1V3yuOk+q7Kda9HNYsmdP4kk9ruuWaHb3gkk9rQoum5bK3mTKMmrJ1U2LkXy98cn
AVBqdGqq3qbjvZ4ip0YXMoDFmXTUQkZ+h+iTIKMSfF8rAywmrHwocHlOhBmZsdSO
RPwl/ioiEMqpqErfJwLEDeYbCeWsMmu2v1qmtIrhpxO4v9Mq1TU79SMFll7E1Hk+
YuZzDQyMGtzZQrVfV9cVsPnVqYvOkh5iAmD8NRQTvrxtqV95Hee2sJ5Pca7XYDoz
lCNRN40tz8O/VeKwmXFNNJUFPvcin1+Zzel+zA2yM3hRp5n6gde4b2eEf3SyDV3g
EoyflWv763p6DJQXRmbturluJLVRv6XqVY+3a9cuuKJy3pXXfAOgpWqexsMjJk1/
KVc/HUlIuNYbZ6zHiUw+P1+GfWe27mnMSLnUza9F/NL2f8ggl+1Xr8zseN1foRCn
sszOEK65BLl25qh16g4/43MrfHNHSEJuJsJz3OfEzrsU0qSPYN2mC6EJjc58rSy5
3535QKK1SmXU6+5tZuIuw8EODTwk/YQx8HUQ1THz/5J/eF7hU89y2XKPD48OIn68
zz1gZCxMJCpdsOt8miZm0HwyyvAKQcabaxgMZLXS2HkCuFWQwZkZRmQ7WRWYrHzT
RgBU6bbLgEf0HsDix0vvrN2hcz/79z9d44C06dRnmDS5vwWXp97Jh1Psbcu4BH8q
O53JJnhRw/6SoYmqKWmle+Vb1DMF6BhqEh2/atvA2Oi51MDBXzhmd0Our+SP0mLv
zZkm0153/fANQrh7JHKQXgy7FcxY5kLbndgVSKTPdj1JKtzLRPYwyF9fooqqXbh9
GJoe2Ec8DWfMaSHZvbyFiX2arolDWABVIb8SrydcUrGpfuwJ2dunnGHMMEeC7vC/
ZxDcBdnH5FKGn6875ZuADUFla5pYvCrGhaholePrC5WaseSNa0Hc/H+craT0SJmJ
zDd2U6vw/nnlmSWGkubpFUK1i+l1rab/4D1FWfwaJc7TuRvlhxca2oIlNq1nqWqx
0oZIlGdPPj1ni1YA4YpWx1DZ3t6PVzGNxiZdNl53jxsdVUxcl0cdPanbjkUl1LE5
xqizbp5liidOg1Y2FC6SocBVfK0l/GYijDmx33jBxVADsyQly5730NWMFfmhjroU
N6rmBMZ6vwu/Q8ngQ8y1dXS7IAaCyewiljv3Ot3OFPNCdc8NXn3gJeuhXnfxhJ8c
nKja7uPI5RiFJlwk0J5Uf0MeJRm3RFQvi6TcpAFiWdrrU8fjoMr5hlZwhhbGrQxA
6B9p5lKfNOMLo9ID9r+dnps+VoK8seY9Xrl0KoHTkpNyFB9imK4yryzd1XnDHbaB
qTTfoAoQU3ecltUU/ekqHXglSuf7d7hNQyF3/pug1dzxu3oyX/YP78lf6RJ/gCx6
xHHRKY284Qo6GJh39cOYkwiKihWwazFBFd6Zq4CjU6XvyagMm9mHfYTaRDCi09Mo
Wf6Glpx1BiF+HnroZjjnhA6n2akGhfR4E3No/fsmAIbmrREH9CrLfXHBtapNKeCy
FcE3iNGqjRIUSkaLv7qLvVR/9oSZCf4e6kHsvOCsIKXvyk8GuzxnsiEr73SASLQQ
+7M8QeKmf0I+E6dlvZCsdjpSPKbGIVtrtZo3BMIqBxp3vTCY6o+8kj1G4+db6N8m
dSaWM2lDNuQWVO+71Iz63OViX08r5kQoUGmR1lvBWrRQCvmH7n2h353ik69TAprr
fhxOB9dzBXnqwoNvUO1H7xAkmp5tKOf5TXdhwL4lAGOO0zTracuG7wWA1B8Fabr1
am3oMKl4afxV6RvK9xYkT2AZr0Nn2bh7zCDRLvTVUyVr6+glg7JHmuS6r2EqC44+
Cxk1rnQhznmm6sXZ/xuNqm2JAy0vbb7wVTniayQTIc0WZZWNiAEAvaVeJ9UtXpH5
0FKNBXsZfJO0ajwnBeaHLs6j4uPyEkwvBkUOCOry47Yon1VOZaAw+thMpSkzXdhA
XXnx0rYvKz3+wemuYGmkg26XZrrPyTPCUglUqVmfjwXJ6F3JCxddSlrQqdjVAV88
OVBkS1nuC2R+LoQDuQ/K0ftKDOYn4+Zu9J7OaCaeNaUeFEM+1xf71pZrPD2mxmfK
qI1s/54STcMQCuIFA4QVaWX4U5zbK6qdnqgDmKeUNrQfffQXz2hShE+PMeQivt9W
enm71AEUy44htHGxcj/i+F57OwJ35rquvcfD/C+ZniyrIWA2tj8AZ8ckVTQU+EpR
4jbL4ISw148NC16ekpm9kG2Sx/l9cVUpbrwbBfAj5Mrmwf0mWYuJow+sWwgXRv0r
u028am136krVttoXSjD/H3CDE2inY8iiS7KYiWux32N9tnvLCK/ACafsVI5bkLRD
B9t1TdTPpb6Qp9NTVHS8YYrJnO9EP0V/QAqZbQAk4FBsV378lQ2sfgbNCnqKHRrc
Mwng+hMQHFX/2eqFf0Eot2MjYT4MpLTRD9DHGhQvtWXk2jvQ/jOOj4Z0FZZi6rTo
Q6+gHcq332wNR2JTERkvl/PWcgy88oALiQOv+r2Is8XDlhdR7ymkAJJQpXip3z04
fSoI91V9IE6DaupqFAjcRYr0ND2kOevfsO8th8m0THPGGY30nOk9lLfqhmjqw3vj
M99/OT83stGEqiiJvVJys9P3xr7a6ZDyvytHS/d+iYnHsre7Jh1przwLBZ4Vu1cd
CoRk+IutknJpkPbZMLluvGwuAoRsrW0W9v03eRmKWcKMIogM8rlDAu59INluEMqX
I9vcnSs6P2JV38oOZ5zvP3ADm/s04el/o+0xAxMDm40MnoJtFm4FfScRKlzidhjV
2WqSdVDe4Xi3Av8MzJxpdUVsUuKoZQWvycpiCe8xbAkKZILfTSMaQ+ggpETdmsG9
FLtZpBCSXkc56EfxgHXNbJpc0qHCgxmy1+CI7KTGR/bOzFzREgVzCwHzVcM36U8c
hH8TWTwF3/+nI3m7kdPnJEHzYR7J6eV1yZogsEomHD5bf6Pie0XKUtWI+osnvkLx
QBEA7Kz8v5HqGB6pK0b5N8s9dZxgZEVog/8fhCnZEsx0REVVY11ULZL+/M9kn3gZ
UXjCaK9Ol6iiUaxh8Uu6zwEGAnXo7z6WrEGvPZcxQPmsapDG+Vv2fSYxcHpkzaTS
Y5hOnNkKPrL3mMfTGDWQB4thIVBTm/uIrzph8LCIsA2X2dRUJqPDhkoKaheH3Orn
8OEUrPhJ2npp+9WF4wDJubm4NFMJVpvGLcfKvxkBquDexUs+ujfcw9JjBNNk3ItQ
Kp/LQCtFnk4eV0aaYouhuCWfYv8eWy1SQpEnoI90ZPSND45rQE0KTeafl7ZbSCxU
SGS107clm1e0GdAdnxmf4+LK5WU6kr8Pn/+FZ1UE3juCyx1Ejh9P9hKLe10c4TRl
tFvRzYV+Y8gzxD2g48mT1/rCd18/2Mn+j32fQiAdXTYFSONSexkstDBOgaKLofZi
IaXHpobqg/YDovxLAwjJPZqfykprvdeDRre075BvGZBXXvWuRyn8BK0LakxCl+JH
C7DoHFubip/vb0xxP9E/v7jZIk9Iw/RPIh2USe/arKTYzKWIJZIGAvL9YBHtR4GF
lHqWtCSQsb7fhAiw+gsiD4i9xL2ZzRIiU/aPANiDdZsyjHCr6uTlHUYoxtQ+p97M
21lY6nj7yuFsbRIexmwinQfSwHwmQVKWvMMVKrtW805pf7VGwl2Al1euxg3iLFjR
FBzPzC8ZyOElyj+FJWNefzOZR9flI6KlYOQo62F947OlII5a+BwkPgOzR9NDMoWD
dej3LMsBGmDtD9JlADVoim1unuvAt/2owfdooWU+fwFk0bLINMTbEqMzqO+PG02P
ONaTTOkXIsHOmo/knC3tHZUvUMcHA4MlQxgnApJIxNPfzsprtYsaQ+bqH6Yi6ACl
coQxBIhSPaclFQpaquRcXKg4Y732wesbD7KMPqTXFSu2P28pDzGFFn/0DM8946TF
us7N7hTsn94bHAYxahgFd8pHBp8qOMLTCU8pqX628wYDiL2yLMXQC/9f2AruvADr
nwj1p3s6OREJM6ARldJ3NwBjAHgwuwYIW6Z8fe030UL5V4YRQCD2THFKRvIs6WPl
nWtWph0AURDlWYu0GrsAbHBcWepdNIIdlGtW18XNPHo4w40QHCWvj8SM1m4qu4Wx
dNUBrc+6SZoT7Ab0sfxk079BPNH8NwQDSvWlEqx3liOm30ltVYtpxyFbVkR3nHgG
0fsRYA+6yIvZVsmmklEZg6LGv+r8OknFB1+SQFmgFhz6nOGiROb081qiUwtJTCTm
RdKEx42dPUqSdxM+zlyaRYJG3dLkeQV1HHgkiccWnEeQROmB0toC3vnDofzQnglw
6Tr2LeIoFkjx6oKztpVUdHpQCIc3bcXUeS9vXfLecF7ngc4QmZoYeu5lRpe7a8AL
DT0XLl6nNOO323tg2prGWd3ebw6AC+us6pjYPd8Ha3ErPjkIccUzEuJpqq0+RIDB
AvjVVBpA4q9H/GQXOiYzSb9aflKEKbiLFlqlVNqf8nKhnhdKUaD1EdFAGMA3KqZ8
7YZUBpqfcFWgpqspO73xA8AMOmeqV7pUla8Ztl72WkARiIYEQ0KkOqu7uwznIXo1
LNk/9XMn3Meg6MySJRSF5KHHpkTxR0QUZObCm5BNdoZGyorOVb5zhfXkoPj3xX8i
9ghx9vyAVM+FbBJAJXfeoHiWMtIq7+dkCeF3nNaOXSKvH2WmGlUvmqEYUoeiTxmG
9bM4gzY57b3fJfiJe/fyDIe4WyHadOFpfGMs+6O/Xr1zqfVkosTM8nf1CTQl1jOk
Qq7bUgwq6TrpEHjHxBAa4HyjJWtHqLEsLaGcNa14RPA74fXWGbC4leifxKqraod6
FRG/qKiJiLa/8ltiYpgZuYn1IJFL6HMSyMu0aVzPJQN0xXkzO4dsQtHDWpunjVi5
azCBl9RD4isZcIhjqChD6L/bDFYhrzX2ayI1lDMpdIQ4zH+ZcKlEVM70oBcvJ6Mw
puB0/tWJVvNrMs6WlY8gPLaIm+/ojeXWSy8Bw1f4X9nIwLOAmBR3w++Sp4kCTqV+
pNlcmkoF8X//qy3qHVytDUy3h5HvSM/4lYN3bFRUcNQ=
--pragma protect end_data_block
--pragma protect digest_block
mMvMUt9aTpU09PmtffQsY/kyxTA=
--pragma protect end_digest_block
--pragma protect end_protected
