-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AB67bsAmeTEjgIpfOemG4JHr+yEogN0WMF/TrXWWDeJmTACrl5K0nqm9KRVqXnQbUFlgOoizCZJv
Z0INKp/3dIuvJxL1h51NDQPoFWcUIn0AcJ/3bZ1jmLr4NgGq/NI/XMdvqNwOW807QsTAobYru8AU
Y1iEobniIHXMEzqREcIEuTtlkqbWmffZAHQirLyVCXvNkcWfwip2cukj4yr1Fusxbsrjy8WFv/1N
6wZDVf0OqghbB7k6NgdJzPFMBarpiXKmyuR3/pl/xmo+HDlA6ac/LlqwiNqYINGRAT6fTlSfE0gx
h2ut4CG/k9z0JzHBYsIOK3bWlYxwxlMjRbEUJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13232)
`protect data_block
kdMAMCpSa4ZGWOe5+rX6+fkmuASNDZcP0Qf2bwlsxxTAhar4nG80tvQxNNRlE2+8bS+Boc8A1nHN
fAL0Vs0/VuBi/CEnKQ8n2vbj8gET0Nk1K1VCtxJRBNwa3aBUGJEbMsJH5KJoehsybslfvNELDd6q
lXJS176an2FiC7MDaWU5j14evNLAb4g+qGuzlRWmido68rqO5dogWOYafeGd4ExomVnAd0o0QavJ
z2PenN9DMmH5PfKARRUZ6pLAKVgAYWme+JK958Oi2BBLcXrLmOD3M2OoO0i2GjuMvv+dCs2dhbSq
9t/HPgZ7sWX/sBKgnVIdmGzKIcLEdFcc42Xx/cL5Yqh9Gh8+38Js+C9JJ+9kh5CK0SPEQ/ih1z0+
KoFSzmRRyORrU6re0ElgJjxfdvS00Ry34IxW/DvuikjfVrmI0MdpSFaiutP2iI7V/jK+XP55Ubx3
72y7dfWhwZN7e6NrSY846c/tgGKB538qlDkQYCOx2B/8aRAolRJ5DwfnwHIc0jBc+re+nfHGl6IZ
+MWHynq/RJKgGG3QerwdlXDI4IwY0O4pW7VNHkL1UxJcgKgA2SlLhb9UrrTGvW/8TrbNozIs7aLu
lbSrsvzoYCLMBmeh2ubzhPi6UQa4IWE5/Qxd3iAWuLGEUXZJoUEbrY0PxWBkMvUu7S/K4GVMYDks
cfqTx35v5xSqWba5d8EOWaZ0MQw9tgN7jw+IeZ7DAQyb5bVPSK4YxwK7bg/E7YML9rlAj7NpxBxl
fgoWosHRZaRTVGd1Uiy4CGBlQROfjidvlbwVHyXH/DD1YJTi+lUtlt1UbciTzP7IYV5pVKsKfIZk
nBn7G8mBdxXfv1s8wgb4Ls0o6KJ/Hy0x+I3OANYIy4nzpKA/ptMlstkZ9QZbEDSyIN/D2raJD7TD
Vq5w+WR/QcmdqiQ/y60xebEwZTp4f/3WLZDk3Q2LmxBqRPxgepUFnlT4jb7yKWU/d5RUeq1mqIEl
fA10GEjMUofIZSTjYza6VOEgWf9gUnoUtZSYzE3yGgWfd0GwYIcWac6aDZ91LvyPHmvhyxGiVMtm
v/ZRgaUWMV0cnQDSdRDCIxFNUzrKlvFGobPeFAswmC6Q+AJH2p4b8V+RAFe9piQNqJw8G2jgeMAG
7bqldFWkfrnrDd2HeTIlHChDafzL/hx1rVk1JwXYN/JtTDbzmql2Ek5WaPErXQo5RUwVqDxdkAno
QraTmvnVPSyZV5QVbZrcbKyLmDTm0410nPQ+0sDU/WUFmxzvLUgAjws97vER9FVwZec5+T4qdpla
nWZw3koWnhVqmKfWl7nypodSAV+4gtF6kRHZRC9rqtnP/noqfDAZASU71wqrHrfHhC0MnYMjOOBN
ouh54eeKVV1O9UyMAhncsqD6Hl4T2Mw1VQmVlZIIFMrh8JPy31XExLvAJkQJPy6X8867p+tvjdzh
ovbCO3BHqB3Sb0h9QNljAT3NzmOQuoeuMJK1213hEvfWipG9sqzbk8WXpd7jWYQsTc9ViRe73HbH
2imL5C+PM5ibkrtj4HnKPlf/paLEbhuLmw9USyq8qAL0Q97Rs0b0UzadlWXirbJ5cIwppi29oSLi
776Twj1FXR3wSB9UK7GDGVnVHlkeL145Odc788id1VtnrE6aTkMwxpiGf2MzR2TR0ib35Rby0pXC
U057Mj7fOC4sA/u0ta5kd2BzG1jN8+VB5QqXrLTOAk4PFoJNCKUU0NNrXba8ulZ7AiEyVH5j9KO2
URpqqoLlit7PrownL5737mHubb85LHwlTP+xH66k11PNRCoJu7jNuhZWAUsJS7PAxsFRAeaKQwAs
Q5O4b+BPjzH6eMEc3A+G65XBiaKSmAoNMr2Ki4ANA/rXqod2WyREwr8OIo/TtxVHEn1wjD9zS0ft
rGU0UZtHvZcCV6MjIoZHWXyaODq5jAKhNb8+bGUShAysAaOn+6p6xNEvXixRj24T0kDrZfaL9Gy7
6P8OQXJS6+MUxvvJL0exTQYphWxlEoAvteRK0GbWo0t+2sz5JMti9C7q0ClrIB7G3jA6Uuax+D7E
bTiwOAeUFL+KOQdl0u0UmHQjRTGPEqUCKNNau5mxeA014AfVcuf3ma/BPpmhqjvDSAD6HqeaVy4k
KXWI3TTCiGdzaUZWuKyweoDkxpyiYvgUqE36qQffodl09Zi/Y7MtdHW0EhH73mLM1M0Zjo/ZbVJX
OlGsnpYxaBLWwNzJu0X9RwyDFSgPxmCgZq7+KraTW0t0G5vyM8AqIMFWdrsg3zWCT7T5puI4mBFx
Wrvf1+u5VajGNFKpwk21hZJwBAarUmoxBLm+Votj3RO7S5qGiJ5C23vdG2pWItvXrny1xsnawvgx
AROOKnBs7eqfc3FkpzBHibAwc89Dljh1bicxCIcDLY2Cn9XtlUVLaGl2Aic8Fhuh66N4z1T8lCbJ
wIZwMjNskhKv/SKlHq3zTHsbWpdumIsGmESqFtOQykyJMixu6Ep+b6P/YMaEj3izByGDQxwkv+CV
WshYQWZYplHCVDjNAxl0PZFI9P0Zuu+5bFanK1oHKQ+6ypFWE4LTN7ItPctdsE6qaUvciQ1hI0JG
uUrBrfpXEtc2dpZ1gi8wkAiRZjLGBlGUbobAxH8N8rCQVjVv/CO5/Lgrr9ZQ0+GeWi6T0ojPXfKw
pIVq3GdPYOs4pcEdP/sEbwZ/Bb+npF5IOr4g3G9+JaqmCH8QXCqvtlXYSlhvLIl8a4JXcdeYrh/5
nkjZGDOc1GuVtuxUNDVMAjbHiLFtKbPuL72q6se8wB4bDahQRd2qXsNOZ71tdARc4RN82EPR6qN7
aZtdEyJL+3c5KNa2GEW22NAfSqUnai9R3DguzqMKlPO1fXFqheqdg5dvm9Kvj/llCDGhdZpR2IA1
vBCUxlNoX73xXeSIcx3OTV+fbTZTG0y+YFvBg6hBJVqStc8X/Dx1oL/aL+KPBjcXCuqW5YA6ZzJe
MpHIwTRINkG5ujX0ALwQX+rM6eCUKUxrPj8MMxXMupmlP445G5PJP+VQkPgnq4uydvuanJqnwL5T
j5abn6I9WsxbEkw28D5/0DaZGAKIWGVfART1dFQEmN1GJyTg5UbeJ0bgqEyIboKZWxpJJdYDIY7z
eAOVwaE16iSxFXhp9PVrTVJyF+78nD6gMftHngcZkN1HVzVzzNF5WRF4rFAzE+WKDzE3mzMR3Xi1
vF+HuHhtnTcpw4u3jAsNv8SnOzY1m+4J2T2EXq+F4AKLSfkEZxarOJYqjn9O2XiojcvruAc5ZFky
yv25G+JP6VQnr0dtywpO1G7SBef47vFvh6WfamjY++7UTQMg94/7nS99bmSTk9A3OtSbU0WnF9xC
mmSwWVwTFOa3RGOE536l/ry6RcTL6z6FUhfnhsRYdz6gRvFBXEFC0VCnwQ6PgN+NGHyWfSj0LzTz
FS8Ue6Iaq+L60luT9Guc4ZVWPwMPvhqdpXrWppK43NTBOf0SE6Akeb6JdgSpZpckuoIrTrUghV2Z
E+Vm+VANocxsPt1e1/EWBrO7dUtoJU8vNbzKEhgGgTq1pM+M7d2zwYHBJfwe/3CNYzigN7Q0FhLE
mlYWGi8DehhKqYAQmwmGd1FLTLKmdUS1X19lO0CC8lCYNtpzn1Es2q6sHrqdlnQniGa/S1nmELjW
4b5kySztST6n00HizGp3yZRlVmY9VD7o97rJCy9fEwpJar1q4RUgpIfDHgtQVifj0fS4fZz4pugS
tI/yXaXH9xQrrszroU6Cs5MgrxB4rCwLsOWBriEmOgFJfdgbHaWKCZcczxroPUeo6a9BiTYgS0PG
Op7awp1O8Ptf9mIX9g8RliRP2c6Lp0bXHsTLSBvMReRhN8vhkLmmdexqcxjLk41+nzoOrTpA528s
DW68KpvYezzXKH9q1FNGjwSsMUpABEddaVaYqsXNQ39BnzHA4AWeOcRBL5JD9OXC41VwhRIDafKh
vgN1FEAJbynjiCOPXwDPz3LbWto3rjveNdr/swxxr0+KkmrBQZjJUTR9Jd1AxLa2QO16Xt5LgYi1
K7K9D6xWEV8u/t92UmMBjH5zjflZ2i063Clpr27sHjtl2LdLJ5n44IQ7tuokp9+19MeXJJY0PHaE
o8qTEddTehdE8O19Vi4Canf5VqFGNFe9os0No99MTUkZMk1jEgcTKqzcsCkeGaMUEvo/Sr11ENwZ
CoSE9YGiaoRXNHxQ0Dw6F81oHiMLcCpMjvFo7EQ6aK+McFDfVQYf+ewWFhS1bu689WCGlek7F2aN
eZyt5fYwBzKQEvzQnRuJbLahYYRzEcZ3Z9CyIoaYInAcVQQCoD0po0/8Km8pmir573WRV7RvNIuB
LnLUG5h54PgMcdL3bwZj1SzXqx/znEu5lSket1Sv+Jcf/3N4w+QP7W7Tl/bLHx90pqAZuSza9M5r
64eqtjqBzEpAD3VYOWQssqJ6eM+cQ4wIC19blWInJCvVSrvR7DDHc1y2x5Y7fnDemo6yOrWy2+vv
iQTnXOexrt0GxqpCcFcsvdYUY5WPpAEcyaLPcNcgqrmuzDKXFNZvaSt8hWkMoFOOYGD9uVY3VGAw
obK47ZRCz4JXanhiFDrF010ciSlKBtO601EFfcPYRhFrIpMvsmwmnBug4bG3Cy5f3iB272z5gkIc
wO8dxwM2TgCv/pogdT2MkcmQ2WLn9fHJUvBuwGzCs2M2t+FIGYLsACo8yx8MGY6IV0SFewmfrZf3
HXR2fqIGDPyXfjVi6ArjSS+j2zyZuL4ee+PzeuMJpzSTV95grjJp++Rrf9epGbQE2eyxhuuVfX3w
9InvKTkuzAnxkz6FWDOwLg2G/h3i/PszcEBUkmwi+LWQUk+IxMUwS80nQu4BiHtBoXMASvw0QAOk
CukJbun8R0mloQvnWJ2xa1C/ClhrcCSsXsn1z8Fwdv4ja44U6zKc+1mErXOwr+3RsBYOnxyiB1eL
+OK3EeSwpz+//vKTX70x5raoblGwxv1/VtMzj4vp+tIhs4icIal/36kmN3W612e+qH56Ap48aBVz
CmVoz7Gqjdo5YxqHuEI8M1MyJcsv1T5Do+iuPTNvsTJNeLe8XiEKyzFx9i0zhT1CE6YPNoL5WZH0
K6xMOfezP27l/KDHKN5EfFzB2LXaKh07EqEsEKzrO76gu0wq+0V+qkIjbTqzfSNroW1YdEVm6Nyy
odp+4gpO6Jm9SRqouBhRplwZuNdC0cxM21fGrSBNEFeyy3gjag73VpOPBW9O0G17RHkEpu+TSvlj
IZoVW7TxUZwcW3mW0I+E6T/y0HHpKIwZ0ZWNhBbLOw6AJjpD81ukqaZKOVjrK+zihpaxYEWEePnt
omTAcyWc3axOLmOqZe7/vTtOCPVxQBXtoJZI14g5Pob9UWj4njf92/uPIA8CBG3PGE/uvY7Vgldc
4bGKQa8eO6CI4/ylKKopvsIvVx2SKkNS7OmyN+uwRxt9zL4s7WMP7u3Xm2fcDvMGwiCFhH5HQqtr
95+NrJ1Y68f5JLI9/iG9c+w6zY05xd7XCR8BFflSGo2NIUQakyvr7NuU3oBVieDzzl+tEZJXCQ9B
FPh/Ay95lD/ksQy3YTfsypARZkckcRYBBT7jTMOa+aga5UAYAqCEb9U80VmNdB+X0fnyU3hwCeb8
f+U3ZHF478gIOni8jC6czpd2cr2QodA+Aulst4gVzXAA4gHNtDfd+gSrSDaoGm73iR5TMAUzfc4H
APsLMaFYML+NUeQDOMjcqvy3+t/WBxMbKLvWgIp0n+asF0hnNRbgfiQ6dewhKPnzPmLsBBbP0bVP
LTZbsbovWQG+AXyrDVIh5KBcVTT3PcJ7QL2vGCdwV7VGn5D6fcL/htcBCOMfwp9qLpNhhd39OQG7
h3FJz3BwQT1WJZzVUHMBnDbHoNytlar+wIYaZXDome+xqdhvj0Xl0w1KKgn5EPD3Ie00aX3ECr4Z
Wcx69k0CSD98MpgvKHniS6kDY/SSS/V5yUFZ3mn/8OWoMo1ogG7zgX3Xm2dKly6GxAsd+YQqKuxq
A7B+NKfTHXMd/Uzk2YFrNd1kcdGICh1rt1RVb030qe3TCFjoflmQb97pNNgSywrAxe1KNqortLAZ
HufavnMKghXfkzbXUL9o2jGt/X6KCy51AD6xC1z4lZ9aIIkg1NVW9pIAvmEitLXyX+bHuflaIrH3
o7dg8svAjYrgBDdTYoLVhtFVFjNwgHl/jsxWy5je7HBXPvuDw0VJEsIpzneIHVlHbck1NeJIq5i2
6536JCZ3hRsxq0MLKBVhi3dHKaUashoF0xqB7twOirG7Vjj8e7c7LZO4haKQnEzEdIek0GrbA01n
hnSoP7Qduye4OugkjDfcHEShkJKskHPcG+ySDGsx5B20ISeLVebt1plDAZaqNre7QRX33b7d9s+V
26xDDeCdDOA7a1P0IVczjo0WpCLekXD7V1MGGR2aaCZTH5+hcgVgQjXYtuYqwiwKfDf94GQEAs7z
CznH4hO1Bb+K4PrX0D71p8OIOwXVZaABTm0o7xkBjpwF+wmfHyO/ZJs6RY8YvGDnAz8N7Mu2IDua
n10LGFkmSwKNK+FNoLMeYumpjNb1vAxxoFEhwCxHuqbSmeuLbkZYvEodFW/GysYTLuXK3N3UFCnb
BJ3tFTTICp1ZxGs67y3hAyVle6FP5JaDftidwWq8OOKVyXsLnij4oLg1wRPWRIJ+Bj1VSgwOR/WX
2HmRn4VODo7wI/2UiudUaXEk66ExfuUzuTrpggGj8mNhvsWeKoj2YH7ekjq8p8gmbgoXZBwApqJ5
4Gvpynu+bOGX+2+7ZTE/9lXbRfIr2ZNVS1FNx5kcEytJOLw65Ci5gTI8agSCmrNnIm7Sb4Ba424x
ak1i4EaHR4OGepAUAjxRF8+YBBZhd2BYX1YUucrYvE1adtst4w60JWMPtpL532liNLwJ+O6jX+93
ecvmwh61n/2WSmJX6P/Yq5PuHUKmu2MNewUN1Mrk4doQ2jqmKEVGTDbQ6YhfRzMj0pemhnrsaS4G
R6OgHu3GyDQQLVXMmX6FFoRXenEnJ/xxDtt2KfXu2eusTdkUJhFdiMGbC6loEyFd0OBXgW0k5E7C
lgPQyQZ1m0F4zJGhNcWMZ+0RD9YaU+NwEfkY5/KhelJl5rgARL5EkNgyWxO80DueCJAuxZBRw46n
6DQe/5b2U9YK45bIHnmiCbhmKv7m7f2Z7I7hYBVWAWS21Ti9Ry1s5eac4MKkSGkeA+seYTnHLpOH
PvdSTR7rGAsIZJJ5m+4IAZU2o3eg+0k7Z1Zahf1hn09z/t6DAsmsejxf3EZ2LR7C0MTlftkosP9h
uCDB9I5TV1VLBoO0spANMtoi8L8F03/lfRQ3XQ6nI7LdOBqJmtZsvp28btn9om0JeGAQDeQnLxsO
k4Uk7kqLLVWJTksKH/SGNne6egfP1isUPupQsuS5Xxl9dBvUegyevc5bWyat7mA1hf7UY10bkPkK
Hj73SyHoyytOJoah9BVf35I0PySbcF/8NFvfBtP6Fn+V0uN7J5uM/6pVPyoreBDbWu6hxvrNY/vm
GShEsiHR2T++/AmnxMF9LB1wtomiGYmxvZ7HuSuZtAGUQV+z7mVH+eAGZ1guixySzzEdI8BN4CNc
rFUu9dYUWQwTtV71tMkOBD0VEAE19FZq4XChj4SSTCIc9AGMxGldh3NtyFcYsFKzNwaKp8aWi55+
3fU3ahFrWgCM1YuAyBpSbYkDQuyB6wbikA/pZYsJX2ZKfJp39vCAkxRxqSyj3xse8kIfPiyw5Ch7
WRq36Lip6cNbqKglaEL3J1Ai979lRN6vk2R7kbMoQnEHOi27k+w43toww7MQCkVaKrEFFp6LJ4TY
YQNQIR6DfklT1aFqRacpx4+InPeBoAzKZuBgPyH5dKW/WALS5dAFxkq7CFDphmXduKgtKtn+zbSp
uPvMmy4pJbvdZjDi0DcSiu+KnE7xy63+9LqZqGyAA/c4uSh2kRzhRg2/xVIzQenicIcp2rq7CDKh
eykSBFn+dTy67Jhf8qHU6Ji0SqufAAjUIIM91I08KiGS9xpL8Uf2kMuOA4WJgpW0EifF1QkhrPks
dSGwRTC5NeC1OTUeNH8+pZ4ACbGqDhmzZRDDyuK0BD3oa7XgeQgKHGO00qhS34orHEBieZGIBBkD
ECsqD5i7JafaUR06bX9Nva9S4p7spPeN8k0qQxDXLiRmTMq6ZXIp10mO/Cuhb7FIKEhlE9VKUA87
vUenUkF6mOJbolxUxaif8yjJLIYvPT0qHM56MKAtq4znWGuCdv28q9gZoX/BWRX2VcfMYlojwkM+
ZAQK1RbJj/txXz25w9GeCKgusIn5xs/Ye/0yBwaqvKwLXRReUhrjveYR7CROyFqMVxK95Ge+DEbj
U+rMMnTuWwY3RPra0M74ihKqLgXeGrEWVoN/3FWknBRduMiZAg7dH6/3qyuVXaqIC5qGPIHtaqWW
Kil/LQ2eK7Z6sZE8gg/sadIfpI8/eyypad3gzBeDfaJ+kGVMjY9yoj0gpBYcjmQRjBZmjPXjX2gb
q69gIchrKMTUMkIK8CV6TF22d4C3a/DGv88Lfub6SjYw//GZXVTn37wx6uqiTzyLYnEyYBSyF8k2
mbK0g5PYvVe5VSVPilECbEnGYJKstbitLQki3OyHBO/yNfitfLd0taoBeQ/kRIspn8RiHmPfEI5w
WXEExn2QY8A1Wy5zhj7aGxDQy0ew11bHHr5ePDcNeMQWhIsSJ186iTJ64KsqAv9VlvJdA5hagVf/
4ozNn+Cn8KLyn5p9NZQX/mIU+wImnD3nCWX1LQ3C/ouXWEvqlzAMCz3fxdk3xNf59mYgY10xqlte
5lQiz7G1Qs8qxorWdJYok7/dZlHzP8q/kuG+9IaGjrPt4EGYv4KGrlc6FZB40ITRnDtYOeKp3i66
/XmcM3V71EGULZ9jQ+dKORHKK1KftR9QnLxyHhwk2LLgaEW7QGM5Mx1d6QuQdLoMvD5ztTwYZxFj
s93szinyeH5u/Be7+yQL8soARheWESYyWtql2J+6Tz9hHFpV9TJqDO94a5cwiEl01Aun50YAP6yN
/yss04WBMYFjO83zIk3CULYwiAUb1qGJqwGpHkfhE0o0qKaVi7E47+MKY2jUykHoBJcppCZlXfWv
2cEuTvB35xrBwoloccXBAmRVP+va2yOhtvzG/BA1iMh6n6HUxnwDX+hosPii+UYRsbRLREcJFyjF
UZjSSuEFgJrXlJjheH9duPw0kyHKTWJ8GBM3Kek7nyq03abeAsdvu4LO2mvIglzBmJ/BOSZpJhfw
ybcKgCcPq2wj71LZ6ES9mvGL8oMTx007yedTf0sF0j4gQYUryyJHJCyxi+ciA3AAES9yNCY5ffGl
cOO98RAq3bQCtUlK9xCfOR2Dl5HkwsoFTtGg9zeWQm4oduCRNFNsc5rtKngu8rRA5+v3e0Utlu6+
giCEU1ZfPivoNfsp3DfZM5t8KDv6qDwie6GlxCQiO8bDsTF7+jX2477VylHtf0V1vt9K7Gf+4vvf
h0+I8bgsC4uqhFmpg0k++pIOOs5hC5AQrFEgkTQTQZfbgqvuWPXrLUy+T85v4THkAMnG5WmLMiGb
qfnomw1KZfWXTZvy3+9Yk1QZarDb/xTv+cgn5/FGibh3cMp6292Crx6DtySEWqDwZirUzxrhP4fm
OPksGGxIBDvspx97qyES95a/MFyvP9x2i8B+dXjqUat7InT95g4F3ix9Jpoyex8pqCDJapcXixPe
6jk6rq+HYqEzdWEWH+iWyPoZVFR235GXc4WnT7jBxk/xEbAw/2RZdde8CHsRNeV++Uu9qwNeCrlY
pFQF3JkIEqdYXshcWPQN/y0TaozqBrrlKvTFjXL0v0wcjyQH14hcfyFBvPrBe1WIXlA0x2GgP9q2
4NyU6unicFcOR/juTyfxWSQvq8uZQGZ8KG+sE9fJFCHx0elwaj3MekyVuN4WsY1unMRCTgYG2WJp
j0lxWMG5Ix4N7WGGtSKGwC1PoVHXa6EBhcCkhal5VKZNHoNNeVyl2jxDAx3qr0moVnRkMqC7WSvh
v9fErU0fFPlxxAD93u8c6lloQxEz3fSIF6RFan3CEA2e1KnYrrhdKLwl84ORtrvSq+SF8yAfWnC7
W2CuAfw3b6S0W48YTd0sj/fC7zYesJvW8h3rxpUqEoqZIVtAEc3VM93MvmyfX21yzCaShAqYbR3h
mo9Dm271t4gbEP7I2GGo6Wx1mbFlhiV3/lwu68zzY5LFbGWXTujOjazM36HE2l3BNpRUaod7m1U2
lqvkEPDXa57m5Jn4fCc4Kubczx9C6psmyk3Omw7a6nCZaBR5cRV1duhgcjQJYR/5iq22z0ZlW4j8
RBfUrsTnKqjBJwXPqOEz3GO+SdqyCFBzCe/9+UHCaJ68ikS58EVNvz7QIVrpVTGfpy2Ll5Uzyaj8
Pcqbm0GR4UegvRWIt1YTvtpLwfz2AjzDlGXnrYbGfPC9Kw7XzAoyDsQ3S9dgZlJlpxJrMujK3HB8
QHhaFusYQQiNj4gYdTGz8MQEZgilgI5UJh0hfZX760fgmkn4wZsJdhvO9fI0YUJ0cZ4Ti0Gp0vOU
aD4Fx2SnQbMe3D9QTsIlx26AmB0fyk2KrKTpkkr61gRM0vmn9DGZ7Gt5fP5k0s1EiEx4ToSKf+Dt
KT3p02ZK30mWAvOaZNwk/9e/vQZxAkoKFhYaXajWxIh8yWW61IUQs/cH0UgJtIOB+YtrdWPyr3No
4PBz67q1nW1gaoNshDwT0wTwjMLm1hj2UGE56idNxtIM41EYBgk6+A07iSCq7MPKd5FmkgI3QMcJ
vhnmXQo3zm8dOFTJCUNvYAiDaUJvwln5YAFrJf/r8KM3et5Ly0LRpkbIDKpvMNlTe+zz12ssgOdW
TY2SMxv09nU/BdMW/WmLDxY+t8M99HKFGxizrI1mL3PV4T4mzlYTVzbZ3oPckE7EqoEuVGQrSFK7
mCxnBfg/nglXs0r5WAfWmhEyI2co1hA/h7G5IVcOsexfy3kUc41hZOznM5Y1vgIeA+bu6wodCEP0
Fg/bzzqi2ykrkmM9gMxtL1sNwLw+s89yWI6KfWGD95hxDjYd/ZuSxjmNmttajOuoBKFtVqL51CoM
iiI6VcBqlxC+GIzz1YhXDNOXE6lHvztLJvHVupHkVk+BwpzgXJxD29CA8t8czJlBPOmUv58zHBWG
txdHfOq4PGPcv1L0p8wFki/sNuMKcQCqfT1DP4dtzkrfJA3YZubiKAv9AoWNLZakAfTcjCGs98xC
8LQ6S8bC/5LPg2I79qRhtLVB8Vn4XUbF5GpNbuLFVdKoCsx2/d0Kt4AuurCOC+839taXm8+ooUAj
WtHwRtiTMV6uEVtw0sEzGf0N6+GMK6vJ0RAVJzkJ9K0uchMF4cO32EpWa7WtDvyzBKupFbUIOxSl
lpZoUR1VgNzbVUWbvVwMTh3EMZHVnGY+ooLiyxpzjb8mlCXxb4M3m038oG9lQUymwvq9QKUuYUsi
8FMQfpYA+OJEvPldNEqDMr2/hghhGLE8SNdEfVjMbzgUEYuO0e9lvkZ0Bpqi4hbqS0fpReUPZ3f7
wlrXR0aqLNQVzmY70sFrfVkeWoZ3hWFxT4qSJuHQDPF0Z1Hmj4tQg9qPwapqo3/kdC3crZp3EJ9p
3LUEJ4hOyV0msWgpZp1aQor632NrtWipDqvL4Np4++FWx2l1RJ4RqJjrJ3ur1PtXNaoOVB+VZ49u
n+vWiN6pAyir8TdZVlP7aZ6lt5dpb2QrnD7oLX9Ie5Dfnqup8nCrWOvtOtSv2jLSIuk3pD4Y5KVk
Gci7pea8wkKEW+c4IyqHd6y0UGc0RXxEAdCs8kYvdvDq/Sx4UfnvrUrScMU3ZJ4vRD47mNx2dUNV
IPi5Yx679Hqo46hcJxWt+uESh3LpQHRWh0Fxy10IWydUU0g7pUvl04iZPHSDuM+LwzpXqB9j87Y9
bMDmYPj1UH4SrCYdb7RUPo2s0Cpc75b9GuDGZwYuUSfGNyBn/9+Rc6CgIBG8259PlVmH69WPOGWJ
XLyM3D7sbHYsA+v0T40JUhJ6ftdnhQeHhS7PZYzxyKz1Ivtp/0nUiVqSj7CKBElOJ87AErZXyLct
CrZCS8d1HfqGm4G3khZ2lBIGMU2nCHGP2v/pY1k1yqEIwEQAaznBIFrTlOYP5nQ89QLN0ZcHt8zZ
fo+Y2IXwkCW+1175LqE+hF5oBr5Ig3P+sRCvkZU4QmU6TIWpdo32QaGvckNV0htHCQWhJQoOQ537
yVwAfSYGNTVsNjYTf+hoVPlj3A511WZwNPK77T2AVu6Uwx9yiCsADLVKpt6GXVUyI0xM9eYWGOH2
2aIbU/qMZAhJ97lmLaUdFrRazynTKOfVaPuof/vWXLoZNlZVYAvLqJkHpD/s9HhlEF7/tKV/3+Wf
SKvQd795RhwvQH+OBILZDAPEbbnPowSzzJdHkzSRPVbQMjVDI6I7hmu3w4qnmXzqPgrO0DBqHaqn
RFAo6Yr0ZS+68HPCVRQozOFN/wbJTuMm2NbGzQq3JmLWKVGPJCMbVlwk83p4PA1R+x75uZ8bM0A7
w9uw0e3fKX/9isGCYTWkQaI3kXIq8NXHryBgNFiEST3lRjPoMHfQIJXMaZpx0NqR0kqVcpyPLU/+
coawMhFtLKXHW3HFjHhL1dsktbIcnCbIku3WFkKIWGCBzkAxHkOpAaUOFvIs5BmqICThqL2D4zmg
vGtWzY8BTYMZRSSUDjL42TjyJJt49ayaR60JGF3+r2+kU37zCBAKJLhDBor/fRpyLp6fMGqpZ9+T
u/SgY4zm7opI6Bk4C+cHYOuXqHLOU+gaSw1Zi3meVn+8fv9G62o4IMpS5QxqqSttSZ/20KNGlmi/
7ii9/QMoV1loELMgtQu0WFTQq3LOvgKC9SI98ire2nwnehL9c4HyNq8CNRuzVNQOH2mTgWXTILm5
O5rbRcQzLFSkvQ7oKSTgavlu7VmT+pAUNH+9shQnrWaWvDduFvJvPsQFhhBMtXxj59WgaynEf7im
xt2QgZd/iN3Eb98LP79juMrFKoZ2Tg1DXh6Ibvj8elNkrv8jyS7BBfQGMgJi9vGDcaFjz84S1Mys
m7j3z40Sy/jYC/wPDeDIitluENNoUjUCRB4VOloDYTILc2WXfZV3qcdB1jfE6Ubhn37yT9OBftYs
DmPSmU+tiXNojpDxF5ujJo30FC9Pg90pmyC8ZZZCUrcgc13vxfT5/LwjbkU5aCP61dhWeePUhJl2
j0nDYdJb/25TAIbmbl88edyg7fx+7FUe5QL83SRprQf9GZVwyvhahdnzNa1Oylubnr2Nf1shwUmi
aj4uauvlJX+WvdESUmVRRtXOGFgju0QNbyfoM1oalsYGqDyt+NHBzDyhOsvUcPA3UnxecrOnUbrV
sh3NkRxecyp4jZU6m9vCSjjRPcljlV6hvXi970hXiCqPxF5I9esA+12lKOYWYP4sJ/lrH4WO84PT
07RXVAp94AWIGrywN8Q/6J9AWlLY7tKs5ekfKk6oPkYzk7QEqYkf22SkMgcoIgOmRFkKc8jmV6lM
i+NwAUGuICVx38VK1vI2I8un2htcObB5uh8B+Itz0GG0gimk3II3dzbQC/sMfrrXFQ6O7Yt1j1ta
E11qb6s9DXKn8FMy0jR6GIlDSNzpZSvRGMTAPSeQbbDtdPgAq0wDJoNjMjWMKDQMlaIvrPGdjbHn
qXduKxGpgESaDEymEzrIK0F2hkC5NwjvBC7gygv2gBR0/Vu+nWkWMyIFS7xpaWHDT+uYfOl+01qE
1MJlqp2SE90kNrlY2P6AoURVfKhZGLbDVP6VSKAdn0aRPjBNFmEITFi43SyON4kO+I/25ILDgYzj
8fG5NO+d5iDFXjHNlt6/5sAH+V6HawtWc0AZmOVbGN4aAKq6GvYJTxxLTC4fA+4PM/bv6vIcUpon
8zthbLWJ6OTKlRmPwfw4L6yEDZXNR3YmfqMXQxGjxua1Wp8PpbfJzkt5jLe86Yis0MyOjQwCphmg
WlfIEj408XCCDshCiv+AAhTVEbnh3qGfxnswX2tDUxAQXydWLsuHTDth4u+4IYpNJybGBly1cV2W
fhc1Rwym7jRasxgWh/cHw/Xkc0tBZhNQpXLIupy/i7WTcZ5TFbu8JN9N+XjPOHtadZzb/r37FDOk
/s6JpAYjzRIb2Q35usqYaVqTxebFM7IWi10xavEZt43TdPYJ3yuIdT493tp3fcwke2CYogEqPBmy
mKCrwEXulDnRAja03K6kDv6MB6i6QlbRGMdzF7wFdC4jeTddfxxwjxG/mt8rgEQEFWwv/Lt+OVVV
aNOmoyuxose404xb89KaXhVCI0DL+HKvpCKLGMv3uDRbXK8kVUboCKQ2hU1iLu4XRLfh29DkNR/E
sVfIos0+lD5ebzsnDSyVsMeuT9bNoo4cNDUdGaJ0Z8hcroZet/NXtrxh2j5staZF0EG03zK7wh4Z
cegt3Ur5q6RIiWdZAEbOXfSEat50+fmw7zLWmy60O+fA9pvB6k5x+73zyWwqNAmmijUU/VVKRa9c
uSJVS0jrobttMXid7J5TlU1ujP4QHHKeS6CZp9qasxw4YaS/hLdeXT3dYfW7gN0iJU+9c5Rx+Nct
Eh4YVgv14m5uh0oEkCIM4DUi2VxiXoNbRwcbvSult6JRxgbfmdIuwP+u8RhE46O+Of9fUXOPkkBV
XevXud3alWhSai4g+CvuH9JFZkFjjZNNdQBQVp1p4d9ZZN5FoL2VjsLIOe7MbD/jxeQ0bHY6DptB
58KqkhLHkkC5kUy01G9s2JE8iO35PJStBf6M+TKHQKDR2vYtVxvY1slBihyhRYRfVdyvy1i7LjC5
dp5v56lRXrQ5ypIgtuSP3UH/+kbY4/zAdXUgMqldHYkpPu/D4aVuygGZEPcmKQdP593y5D9yRRVF
5yZsXiT0BYMCvh0KdzKvlNuf6lUWRDrv0aYF1IHbuM4aExgwmHAsPSWKAza0n5EU5VdNdiyPi4bU
x764unEFQcw6oX9bQsvCtsULQvVAHsrYnSiLFcS+tM7OqW2ao3ZzKRxFKetfDzS8f5NCQfyt5ago
wJ3qGWVoKFweXjhEgfyT+G0xaBWp4NtNaI3SRF3oPQW048QHIbUlnTGNUUocT1t034DHQFJq93oW
4vCXZ/u5WNWG9yPmjjbn4OZgx+8K16YMOOKLq3Rw1N8I1wE3tq5pfqtD1+ebAW46F0VdZStP+v6Y
69Vpvd18HblopgqeM+7i0cBLgOCFHtxkRv6nhDVTv+Gy4y8SWmChhGr8Am/i1Mt9yeVkSdb+3aKm
H3LiOVXfOne6Lbk+uZ2wi9vSiE6OIMtaoOn7GRICFzrcGMHwlxzG4EQzUxVOs1ChFaMkBcW3jS//
hMsFJo3R0DrW2C2axpFaHQ86W6f68OHWAfoznZPoz4Ydus2aZvA5cGu4+F4qvCwh5I0UVpm44Wnw
JPh8z8GsSn2XXBCSAs7uOHOT/mCv4sI4dp0HZKAUjQXI0IvrDJmMY7YwN6e11v0l1ZAkldEtnWti
fcjiLmjqlsyHcY97wkBSKRhV1XVIIBSTLEdRuhiDrszaKfNOyWz1HVLqcXIz8gQ5FNMP0E+IQnxp
A3uBaY3BBVYSS/HvBWkUgfzlyFn0qpJbjphGjYWPYLjV51Cd1mwUeUDMEtmYIVZg9Qy3cEsbVsCT
aajmlh+8WI3DHbLAwdNThwuTsEdQHST6O6a1o4ZcHDV9AuydRNQqR6yZ2gmcoZuNQTS12cqn5GCL
0AQPkLCSrNJO1lXgnBeQYd103VgQgtFttTbMrtejxzwHCLbrNwsGHsikrD2RrGle8NwrbaC9BSn9
lIf+gQguNnuh0NreY59BRQgCvTXe2AJu+JfZ4Un1Kxwkg14uZwIlnkyda7FVJF7F5wICFSrkc2oO
ReCPFR8JfHZhD0qiElZ3EYVeqHkRfZw4slqUywr64Z5ZaEJ5pCu4/mTe72nuI+jls3KECFW+dbcm
6SXJHifj6pxeixrod83PIxWgxoBcrGhk9icJ4NWpAJnin8x5IIclfFGp+8YX+Q3ExmrTh9rTxVEe
usYLhA74T7NcPugKUPvLs89Qf0CbSV48urVUKRlg0K9H7vs4dwY5r/+mYhsqrWi4srQrDXet8M4g
7p7AEiAp8YjOjU5CJC/vq4+nlzVkvXUjDbWVlKJ3K4ChYjRcP1FRR+DtyDWBiTlDiSPSY3S5F+KR
w1z2M8f6eSjbt05I2t9fjzuIqlL7wgPfc3eaxwp+xdUpFdW0CF7/nlMc+UxaHr7zDq229B6tKhx0
LAekkCGAD4IujPrGj1rKVJvJYhQwMlxQR45FrgDsB7ZEPM5vb1AypvcDip0XUvRqb6NvtzHFOxhH
twE5MGVyCiZU9lIX4luoo1EKZ3HXtsNHut6Q3ScC6oB/D4OtCKCYQaFOC0Nq5zJBDybKAdaCRIb6
oRW5jh0XnaRaD2pg0yQrPBNF7BNT9rlbH2aZREAnSRtqexpbYZPLEh6Rke6Ih2PSdk60ZdU+tGMC
JnFhKVqEo8hxld0cU8xMt0SlhcbVpxaIN73TxAvST6/o3qcWSKudwgOl7+qt6QXllKwTbt6EoACl
X6H2p7tCoGRsottgoB7HnETNN0flrTW/GlPHooc8v68OVbh4BXhZZdRx/ArmDQlqXxgmL3iBPB40
WsKm6VxUmF/XujeM7muT/kmKlMyqi11OeRXr3WRgOtLzLlNvK3namyjY7mzmj9o8AAX8cZ3ZNJIY
nWWiEliLiJgcJaLU4q33jVSACsblpd0flmzofzzH9LBq+f4HnV13MuvTsZqBbBAYzXrXaka/QIp1
pUzVTVePeTRRDI49uZMEIhrKIZdUNPeEeQPic2dnM46FqNbrGFEppm5+5JFI10Cy6jGlD3sDRmq3
eKvukPd+carf1sO1V5uSTsBFykV8zNwelD0vCaqz3MsLkSpvo5zvZpt+EdqcKXXC/1uuL05PWTMh
e9/r9sZEcI4wIU9a5e1IUD6i0myUAsfK18MvVGTAnCTqpCa478EBp3ZB63X8PNHCItobcDBsSsK9
JGIHlJNAlDXgAE347balFGo1YyyZIFA3iyZ9RXcC6wtyoBPa5NNlKh7ZH/aEXTuwgeXNGpTXSxJq
HyFLWt3FN6e766/efBETmZ2TnVPtQiLdFoRq9Va7mpL4WZFPx1Rl7y8Fj8BW3lv9Vtz3SUKBQoRX
tAECvtp/S814eZOs7FvYS2i9/f2y/4eR5Mi3gvGilAjlrbVbg6s20VqLrvwUQEn6byeys/UxEBmR
gjbHbRSQWkdNgVF7XfpRQqLJlZx91uihDXu8pP9JlESuchmlknX4w2xndfrrbvufnb9UegmVKhPC
0riPq+q9+6dpN6Mx/JLQYui06+44ZQO9iXDskf168k1y87Jwh3MEfO7dT5f5KGOmKxezr/HmubLC
PJ1+ndRdUvCMSSE+kWvyl7NdJW9ruaOa4tRHN5R17YPtvIzh2xlN3ncisR3x59upxU6urRAcjhkK
zEgRxAgZzFQIG5jpkgxIclcFtGFaYcNdG6/2GPiVdTGYSUD3bHjktgBYHG2bGsovvLnpQknzABMf
DMWTNYVEu6uU4tilcbwIF0dRTHaehB2QBfheHWD3tcSGiCZmdm3boM0039z6H2JzVsIN6Ud+2I2b
vQid8moEE4g=
`protect end_protected
