-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tCnvgy57Tn0zPUpJ1w4mWHQXH1lKo/4Gw2qg57pfkUY3v5s5YPMuG5Dyj0Cga+sYTWTEKx34Q4X8
lk71rfU0ubEO7i3OiLYBvXHYUg1pCTsC+myUMk8/lR46iHWwpKNiTYcqx0o0+KY5uQWKb+spPJOi
NkvQiGGl+6SbMncI9Mhvak4j9uQk08BN2ciy89sL2uOFio+uhpd9sdHN2REGeUNU/TUndNbM0hYl
57MZ6q3ZknQO78Ddnt4GKAfVnlWAyDXc9IYZds1Sw7g/flSaAx+pl+4dAbBMBx9o9QofP89rl/v+
2Xn+1NKfjhqYpZZcvXOFfdHOoXnACgPqsY7pdQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 19728)
`protect data_block
qQt1WL6CpNb8MMqNqLiUpv0RaTIsuFepneEWMxx5lABUh2dS6/sF0ooCnXfx93mrUKXfmnHzzcjg
ewLHtwa/z6LJqkpYr5hujO4Ll4TYfJbzcGPDXg1lBaohXGivc073DHawMTImb15Lrip2Zua2Wzfo
r30TvAqCHdcPcZLzxGbt1R8xtdx+sHSFAyRfsA9I6BCCbeiH0pJmY91P71q9aZOgcJoMfxHmt0yC
yjtntaQVjp60mu3dOqSIkEguBhhqb1dNmizUDSw0A85TXSuUhkLucC+bta5TuhEo7TMb7fG5CBgX
Ikf/1DNC36w1vLowtpxTWWnM9htuTAl8+Zctrc5JRs047zJWDvIqMBZkr0lYJ8LU7C8reY5Yl42G
u7Y+lkkpkuRbDuuyfOtaqHoTEJu9AkKfpL9nJ03qvqneROSneyKZU5vj0BQ27CmYQXiMe7X7QkFj
dDdpRCyRHwadEk1SVNXTI8dLR3fABCBx68MTYOVJQaL/KnlJk/8Zhg3pEhJjmWJUDNV08HZCX554
WU1vNUNQBgvgIyUOeDBGbVqf8VklHRc5cifOqlkk60jb6NIwJKlGbAsRd0tAhxQzAPi+uALUMLxg
W/80dQdZLHTjEs4BGgD0iapzUh8t7+HfuawP3c7kOVZ/Nwgrj1RZS3d763SaWb0Dq59omBomf5rA
l2Esxm0en9LpVrv+GO3ZeyWuPJq2wjRZGUcDhrb5ak1Y3fvBckZlqmf9hIJQHH0r6MXcFI1jmsIB
nK52sE7mZkMt8kVVCWuqqUXwCC0KDSRrWsr8iCwrbsD/4WlcosvQWoeb6aLdp32idrUKl5cQcZ55
A8MrG4jQrkvuepSduYpk3c2+5U8rWQ15heqB7yp7GEiYsLl2DXRAcWZB6vFaG9PLLic6vUrJz5tT
6Y8ZY8tHaMUWzIs0CnMaz8XW51YcgEhbT375drz+ipvkZg1zB1wx7/zCO9K3qU/zLcYnmwDpRPq0
QySODigyRlJ2sMNkmguW5DTP3NOIs14KvinDvg1lZWcf+5mUIiUbur22BSTv9bFNnAiQnfuIfeKA
wqADA7362VTqQ74oRwRMxC3ZpGyQ46wHkefl1d8F0Fr203SsH9ECh1Mt0Bse+m0jSZ6xRGRLgth1
tRI9KZwSOl0U+eWUzzRr0N5atmr8RyDF2H2ui3F6FJDJy9ah8zdpbqdXv9K4E3DFySjfnJtTEZKK
khNr8t9w72jVKdzzAqMi6mTlq68Gtax7zvBlYbJV6cSVOSqdJQITb3dxPaXoPPxecK8gTiOEIiwu
Ss6pOJK/aEMF16gI6WvC8/Lff3Oi29a1NUrOz44eNcANYdwFb8BOpEV+f4YnjGcdqUTKcmk03AIb
expEHm+s9/zW/zZd09UciyWrzqLOK1As9SkWO5Lmfg8qhykedDSAQB9+Rk8o384HA3zoelAX9vaO
kChWkqtRUkC4tR5ToZ2BmJNDSVvAWaMfde2KQSgfvfdbHnAYhk6pBoS+iWmINqBy84z36nKYg+1L
nmBcjUHhBBj+6/jqIniRewit+LoV1oavEYgIo7nzimNUkx83bZsWBsWYzlvo7Bh2ioQFg3xWL0LJ
g6WIJusQ/Rm2CgF0TBaO/rItVTSVimYKY7gyx9sSFM126OdqCZhREO9eLwD2qngeXG0fnIg+247Z
QhQEK0uVMhyE8z1Pf12NOQ2hkxfVCViXBfOZzZ8dUvf1APpkcfrxQfppm5U8ytZ3AdRCXQoNQPYA
0SvMoNf0EgwGsBu97Cd3DjuxeJY7Ph9ax5GSHCXoD75UpKpCmLz9SJzmjvZ9jcoc2iIpHKG+IWla
69s6B8Y0TwUvfDCcIMjt/ZTpK6YMUfZdJ1QLiRO/oCtvIVtI97h5rwpIrjaPYU+pfQPb3HeyHE0o
ALfEVoKfSnH3kkIeKrw1PMD0dojooWnUkw5aKM9SdJj6Oevq9rCZxx3VWARaanWmdYr7jMSt5dPG
dxp+3PJPsjWD8XUMdAKQwNd+QHvV4BmBtnpGMZ/zLk1KvVcOMkd6ICjnkjo6czsIta7J9VG5kPgK
u4lBXBjOt2jENJCxZl3GPa8NxHQA1yVRFtit90/3JGeGClwVLweliXpFinfB4Ntl87a+CAhySnwA
Awa6+Z3PtQVDL3Hi2WNoTrqQQt9ru2kivmFkGs8RaBzR9CfhhJfFTvUNICQUlgkPverbkbCgBsUq
DTS9FhFWI5Cfda/ZPOTm8BbFZjNJAw7Q0t1fUdPGecFlWn8ZLdm5zkN/uDRhD65ZqBL6doq26lAq
7UZsT23BD4dVL7ECKRPZf2RgFBG11p7lcywk7NTcDU47q4m8AHLK9g32dm79gImbndSQp9r+RI9f
D3OTM2Ix3TTqlsgV6KL7tNVek0d+1xg+nrNttu9Tp+sNfGFhBvlCbqYpDxU9jr8UmcM60z5zv0l6
6j3EvFmwxeXePbeWahA6QsE3gMuRxpqS1grJkKfqPun/DmnyZ0LVE+vIX+IgoQR/8axBo8uJubQV
QelgW7c9lAOgXnpFbwvzBjR09CLtGFAKl9ANrKhdOxnuRahL7BHYPf1fU300pg+6on9tn6ZGiWoI
YewrUFNrPMqJdiqfHffUBOjwTpnj6lJF/ojy+gwgYS5uv8LBH/qfJi0NrYjmy7Wtq3r0ej1iPpRo
fEtQm8cdVOJmBLGnvgSosCoe/jP4G1ruIn1oP6zxmo/VcHLieXBNdlRK+ob4Z13h8mOnBNyniBif
epc6hko6g1elVQ6YmFqJhOj1F7V4OD6iXmdm2SdhDzymoFzMMehDhVWvb5KUHmOeesv+BExr9h1I
dUlJFu/Hv/re58G1AkqQN8N1NL/0rrLqjy6pkfvPUlGeoMAv9z7jWjak00J16y4oNJHHgU43ytJH
oQ/XquAvqFNT4uq/OfLuC7kkwZOFNIScHU4hpzlnCI3omCM8OP0jYJKQlxRnnQ+YQt/ovF/oqWAe
Kk8CRqdP/YJsfqIAatI+jPhucUHVV8xwb0y6b/P1Y06GqEqraIgHjhwSKHLj8+QOZzr+6zyB8MUB
vD1LNhjOzlhTs5YOhV7QQN8BX0K8WWf++KWygR3dZpcDgZVyGRkmZ5Mg9B+BO+2vNA4LTs2CM8XW
bWOTNnp7PP5GoMKJUCoQmdYssrqSGEjarjRirI5siJ+VKGdFzmttsx7SmS89hfh4xz0DAH2fTBvI
tFpSHllqWzigvUtinkGob/L1c6jTFUmdjX3JWd53BHlHY9oh+7mg+t33MZaQ82usCdCWjy7QBSXE
bylcT3ALzdY9JPv0G2dJFEIx1Ftm4UwOsrf/arAyJCfAwc7AcyF6qs03iNowRYia2CfqwHq491SM
RKkUdciNunCrbqxUxbLIA7iM8j12xAyPuDpNqpbIov0BOUm8zF84Ge1TlhIQAFSMl4xFDI15Vhat
k318fbYVU+euOgTGwMDfmKgM4JPs7aEEwAPpiuMq8baPOQ7V/r+omQ5aECuSX8WrCYhL1+qUf8DW
XJM22sqH6IeRUvbIK2hMSbVantufKyeHYRbL+ky43WU8b8EYLyqzO1Ah7fTmgiNpB5NToNEr39tN
7m+USagSiYPE8GSIYzAg8+WirucjODgX8k6wg4Cg4K4p7uvvmvyqiulC8t7gQ7aF3iTiHf5WKFbo
Y7fPa1NlRro6D2lSLBNpJZfU8bo/tLFqUclPE8RSEu67Zq5U6YelCisRyILXWXR/NY5kkF7qQBZf
qD/uLPL/s8a1lN5NYcvsfjq1j8WZjVPeQzGOPpzqdHsBwu/73So6LFuWHxyvFvBDBxqavr5NO3Pf
2O9+tybr4yEki0Rja2EW79FVe6AcARftAFd0sE9gKda4YS8m/JBNROOTC9ZXvgUEUbq7AohwW2AA
9TfHoXa/EE9D/n61ZYzGM+VaXvYKLATwu2UASigJqLl0yB4lmX1BcbQFEubc+LRZg+eQ57typ8xd
XzIziHCE+EntNMpuzdp2ypjGZQqeMV/Nz8A3v2If3MgpNMDDYMUY50+DgbqIhZq5IqX1m7UA//uX
vQRY7sHwZc9j5RuuPQAtoznxcSoCp2+PFf3RPJU4maVeBZ8MxE+AC0c11HrtXnkyrvGx4vDhsirf
YFSgSDRaYaJtD3PmXd9TqJs8TXyA/CXDEauduxDYcAP7RulITYmOmRQai8ILBQAeIv6VsRa2Dqas
F+H5wSyCCsjnmgCcS+2QP4/tG9VhHQg8vtJ8+O5VDV8RVlrtEWy6CPXFgKcsHJYv+FRiTR6VcHrt
JME7d7re8mh3pNaNpYoRHzE0u6UwAfjyKyivte8RiYkSqLka/08e+ITETvDg3pC1Q047VMD77S2M
EvbgTzvdMuEOsG6FKRPQVx29ZmO+mJFQp52woUgfNdPluGukzFdE9dyTKo0afP5XgF2Qf/Guptph
dJDlIWfkeYOHDQmQRqkYCTP1995BcXkhAfFIoJdJ8M/d7TVy/l/q5RroI84r/Ekj6dEA/PnMkdo7
IleKAhw8njXJZFEfoUQ6y2sJHOu1D2InWjTxE9BrbgK2QbMt6C4MDOLdSRT3HdQpGfpgyAlQPs+Q
Fin9mhM5kqj0Hfx6LOoO7kndy8WxrorWUfbCE0qZemielOgXzIvqV/QhhR+/IduV8bdnrNNmLkdy
XQf4wuMOVZCV5cJDEAwKSFysJqk2QD0n8LMnPMjjFE2NqJbmPvLm/sIbLxrtyPdsydDlw8KKevrp
wRzMSTgnjSU0Yz2yLvOlCvJqXqTgQJMkpqVJEZJubCnNEDJaAj5yS5l97ZRle/OmTacypXMTbsEq
9lhO4YlhTJ7pFhKmkYPLtm5KwX3KhkC8zNxhqKalmlMaW5NikhbTg2Jux5m9oEKz6eKOSUQ1v4do
wVaEr6bJLMYckUbyQ1fu97tZMITpB0BBMVo0Ndz+f++mNYZIMUgpgKW4dwUpVWdm7lVfkSss9zMp
/cHGvl7LUKFtUonynkE0ysNH9krftjp4E3sfZiFo76EZKc8VirAdmK+riBvGwZIT4hA7YXg7xH6L
+IkPG7BBkEAJVCGvhpIL4i/RkP7mEca4wTqNrCI3gFziNoclZacbAwbNk0kmjoPqNhIpRXZN5W2g
2vj7iom1EQvuFcfPKCHGL30NTgBdVGh20Gxb48BT1fyjVtkDRZsEDCnduRNX9OQ5NJBEN3y1HuLM
YKudRQDkDxt62PpBM4Woeb/9xck+p2kzXQ4aBv6LOUqbAXsyf43rKsUMazc05egLhx7F8Jv2xxV9
YHiFOJISstW80IYIaL5LEdyAzWq5islaTPMkjjyWF15/nU7OoHJWavmBbBexAlgcrkWqY2yeN9Ub
boeUCyv+CktQL/7o5Lkl7KAEqA6gTCDkxm4VFq1rjPpiJ/shOp1dcao4xVUcBKFnk4C8r2CDA1mm
27XgrsQzmLJXy7xhVomkU4kbiefGOTNk42zMfLv2xp7/fck1mjFLz+V/v0YBxKX6XuZMmNLy4rTC
vvZRaf9ZqOW1ID/HKQ2irDaaWgeWGFjgCrXRDq097rzsK9IbFrA6DOu1v+rDR8+jvfIP3D29BJvK
fAiYUEvoWB9oMAFP7vMZP9Su6sK+mgGRx3aWqzRy5BX2HNreCRvjpEGjKCuRCQOFWAgl5Bj+TP4P
aPmh5a+UdVypn3Z8KwBWn4WIQ0xSbt/GkerYwHd+fjy/CmvvV5iGObXd1JpfkfsCgx121IzFLMIN
zxmrQ6LouWV/MzZO9zYgEYP/R27n4A/hJDgMJYZxLE//E3CoZ0S5MaoOX8s6b8D+0QI4M9uXKPrF
NUv6U7GPYallXatjc6eAD9IAKsIPBQtxMoL4kv/lwgmgZ4vSA2MKImmNbu26wihK1s+v53+XVWGV
9t/d9txB2Sv63cwtl6lpyNB0AAQ1bhjGeTlN3eGJ0I9tNQSOpx7SRp6It84/1kl4HlYW+PV+17Q2
K/bXuMaw2gaN5NO1VbSBYOCz2AONOaX8UVV+/gs5Q7YxNiNgv0mVz9cA8qwOCDePln3ySQwG9ejf
8NzTaTpRBssCRSagTB1kAasIUw+5QMWwMuyXJv83h6bZBS4p6U5Ow97lp8oAs6M8VaTxPSc7X6K9
uXB1eFZx9/ToUP9qgTMaa2eu3AkEb03m3LLxbwh+HTpNP/cVtIPJ4IaG2b/hwsjg5nJy5JIUFNpa
pMDQvyWs3YBwY7zVvXDQUlNEy+m4hhtrrhVw2NhkLRnki55qXbuYvWMuo6B0nXNlFJPw5GUpyrbO
rWaSbkrLjbZc6MSUTDoLMeQ/t6aAAsQxEoS848ZSNvtcuKeohJySmkgI7eYmuwyJYHEqmN2gUSvI
DkyFvPHnRWCuDbGS6CSzTNmoQH85YNYeIzzWStKewIlZHEUL1CBkalZrFO44r47k1JaUEXfhmvHX
dWaKJV1E0VHMjY+jA067PmW4hqjX12iWI5J4rA/algQIm3687Sde+NVFE9Mp67hGowL86T4vAWI3
++K9HG2HFX2Xlxcx6I4jp/eTiEAz/3gtQJfecBcPT1Up6nQLaSYoa8oJOAoWrzfh1oOqqzcHUEM+
FXMsqTljKoICwMrlSEvi5zcP4PhAHsZ5DCX45crv+RUR81Gu5nGXRRPR5z9WN8iOxP8PpWMUOkYW
cIPDaEOdEu0xEn75iVu/fErh640st3Xn+16zYrG60+rk6UC4dNk/M9AkUplSSDy3JicuvVnk7Ghf
jm0O7RMxx0bl1Q5NJHSU1LYRB5CtmdFd2T9vxm6PibPzRlbPU/lLXBN707Lq2y2tmuW5XGobYnib
UQAcMpbEryfDAJi7oPGRJT0E/CysRn7OPdiX8OABXZl9BSChRW84enkGcIWurYOTV+WmTlnox0bV
Jh4OSGq8yYF4cCCZeJkhFKEqQocgjGGNHolZavNdoZUZmzyP31a9bZc3zarjipxSC2unHWybVFX+
7qw6cq5ZI2Qco8jzweBO77t11KKbJHUGG4JuDO67jydF5DD49edEjqsMJvZNDRU5tym+E9Zz+NNh
NeNKSIDKvYI5I+8OkQ+2Dy/KF5teQMyUrsRy6jAwGZT/YvpongB+ON2TeXmYTFKhcksFSWq0Lkzz
ioo46+Vgn5NwpZWbdqOmhGrt0qOzKQUdQdLHIrJsMxMZrz5YTVYagmIvwkF9aVpGq0XFZVxDVQcR
Clqd5NLKvacpcBA5z4Zvu+xsVecU5oH8nNn1LeSHm/whBPE8L4eLYN0szlr+t2Lt+/eE5LotLttu
1sUABT6kUUwBBJEzK5CA8F+kJSixBGlYIYiLYKlYQdir9+9075yNzl2N62QK5a8695MLEc8sCK8G
If1SWXCyFohentdgzJFoPHC0EfdOcvLorWa5KLgnoSkRArAfjHtUs+JIQEB7uExAJREtvTzW71bR
JWdcub6z9YH8QNWKP94c4Y3GZ+WLXaL6sbaXVgLm78iQLA5x4Rzg/+IBf4eUmHJhnKN7C7FRYhyy
5EiYOfhsMFb27vsordjQVH0EYPts83OKvHfSshPA85wYrdLTFJb9Fv/BMhZqYbCio2+JMtsDmD6R
tc7DB0AuBuO5LXvULlw/Kvt1E9+q+PesDto9CYPkHnPIPnZvOM895m9i+WndHah9dpTk7RQgfKrP
svh9UsMY2gShUkWZAGZ8w1MeF1lWMiihGuS9gDk5vLZTcIwP7arn0I9nSDHvMwACbN+jhMs+gzSZ
O7q3HrPYaJxjBZfo97K9NYyFdC1qu2mLmw4ncSygP3uNKVrBavkwB4hHF+8+6GoarQIQ5yeMpka0
5M1gm508CyBeCFxnw0OMpjWpl/4PykIIx5HouEspNu2l5D+0bKOqAIe7GzULWluOiiRZq1aYHzS6
duFY1kDzTSOGHYHm4Zz7ersTqPVLIcEmSWPva0pMACKZxMbauVcF/RIo8nw/2XZwM1pOM3Ww+pOZ
rmvvw3sqJY7ZKrOserJvqAs+1GSqaaZFbyA5pL/IPeP0QvG9Yqg4Bj1NOhy8yANEGXJFZtA6wrsT
mmH9gkIMxkNUxC320+R0lZRcjOLSzRYRtvwYP2WxLtVk9ZzSpc2yoWhHlLuC821Tu4wUH/ejHwpb
pXl3RcL71qfIFS80DEPqAX+C+CKfPSHEmqHmhN6rz9WfZQ5I6+mnnWsXWoY87VUpTtj5PaUsyw2B
FvhynKuc0hpuN3CKI4UrZ6d22WISa87lODJqvHOKUwRK5goexCdZ8Rx/gGXlJX/yOW25gqPW5H8E
aho5c6r/MY36bzNnTZ0W7HeQckrDkoPHPeXA9G4VNrN8b5v5ZzzuVdIO2ug3aHLRVzv+GlLSwZFT
8x0GW8zQW3ojkr9JJ1K2GnsbnbqrZGSYqxjwpyfNv03OLd5wsVpJGqqVkOoPpk8Jm43/wRSduBcF
lIoKJPkLKA8Lr4rdZtbyXteWt9vSjcYZmVmKVdl2L6qczxujHKKuLTeLF1dDZL4u8f7+8dvMymp+
nvY+PBbdGN3synJlxI51Qxm3NWpqtx579om87sfFuSKJBT4Wr1CIzyBZ6eRA2sSUh+LQC80Rxgyy
3RT8146VwoKy+pj10E0A5FvdmG06lsyQ6fEu7QbH9uByiSASPivQNHfHEXG4bf4oYh4uPrNQ8QuI
gyLlmH459OAO3aUg37/oMvzABXhPehjpq9904dvNPGzOjXKVsAw8+TtaBx7N3R3ViGa5mgpyXv8y
zVOEr8i3khfNUDoT+bWH2OUPrtXYt7OLsnrsKp86XrTYm+xu4SVTBLpTOW7iW7cv/jwrAM/Dt03w
bCDxz1jQIweWiMV4h5jhgfA+IvGidKxvNPCSBwMibMo0zQLG5lvXCjyhe4QwZ/aoBhF1+UVqoSsh
NX/852BjOSYXC9Lg8fIH6cXsEMLuwGiTJU4djTcdzdG1JbxK04Z8sN228zj6BhjWi0Q+z5eeIUyl
rSEzdtG53avEgj7KEmQO1ygn7DjAtSSi29ubpCzEIb8tPz3cJL+c5o24HCXmpjdtt2OEk02180pn
Nuq3jp4NXVpFGBmSv/w3fTABat9J8NMzmVx+ze55d0Tqz42pFuRipdNTdjpet5oTpwsbq1d7bEpy
1dPYCzMI5sS1J6CaitF8UIcm00CbziAw8wJmCDQzmdkFXLZequ5amekq4VOo6uIgFhvPrl6sEv2A
jhRsmxIND8c8/24AJ1wTK5zL3Fmp9JhlzlAh6oZyPtbN5hF6u6kyWkY9q/nWwJoqC/UcLftL3JDK
TzNsLxeBhrd39yvOa/7BNURsfUPLo1i1LB2zP0SFDEVrEpWG5VrzheW6IGYjjRlMDZ6lDQDC7Ocf
wbdW8hmKO4SuJAd7EOq502CXVqkRmmWXYGhs7osEKJiRB2PIHDYAPR+6l1clY9zF+zybPIjqte7/
D/JxieiSawWbzxauzwUDrxZ5Zv5F/fgfum7m8cPcp+JiQAoFqobr4lc88wqCq+lKTuS+2QtMJLkV
Xjka3aXbwXxleY+hT83eHibtl+Eu6YC8nyT6dpUiWMHPX1gHUWOwXe54/ktiD6MzA2YxSdmheJCj
7czuGlKskSDN9nXBa9uvyGjL4GCfzGUI2WD0QCk1ZFkl0zEaLREuYQ7g5iFISZrZS9dwvnvQnIxt
+iBZhDm26ZhYyH1m2/URfp7VzuclSPhaOSR5dnh/tNMlNXkf5Wk+96qoNzh0JmvvVLVed9R3e5F8
7CeaW81MbzPA+juQl70h7lpfglEGYI0H+3LcTt10JOPoVJwtCmlk833MMKLNMzW/L4weJTt6fyHA
e5XClOIkxuaDFRYDrtMoJ9Q9504pqLrChk773G4h5Zep1XSri93JSb5kwxAC8kr6QWVT2j8Ab4Ld
kSWZYebufB2H4jn8wr3NfbXPnDbTq3Vhu99Ofg8a4LF3vV6epM5fkaRw7qTr+BhVJ/sx+2w6wDlG
KKsFD0ZpZSwAncoDbpBW073i+cDfsrxwQDivA7cJBEyQQX3oWFlHDM+Xf8JJO2Svp6qkGU+wn2pU
ZGQV8TGVxH0fNlGBg0zoSjoDzQSQTumkL4T1UXk/deOKLSfTsJMgtAitjTzhYHFS6vl7drkJSGDn
fSNUmzEASS3DJPzQFDdZyv3BPC5kTGWGqRmCRNBYGd3rN4Ge4P+hn1zZLi+RPAFEfHdFKFP8DXJW
N4ESN/HUotfc+Man3S7nF50n/afqTITb7PBFU44cuVwvIi80Itteb8NSBrul/t+LBLCbuAhEweMs
JFwMcTvl3UnV+wcDXGemOId7eD8205tLGhaVKKfbjFHnXym5RAtAykdrnDrmy09cT0R/0pw9erMc
sa925Bc640EZwyJXp6xd238KRnLNb6TAnMlnKbUzfCs28Kg9Ba7ryhESq8vj2YYvevkmGHeRIJxy
+jMZutkvGjja9ldyRajfmoziP5TaTpnl/0UO8qg78W2TVUdt8sZ9H5uUT9sMiNnIOYEE3g5HVXgu
+lOSCy2RGEYDIXBZBCQ05Xg8xMylV2ETSEbxP+jfUFt09hmvCAAaSA31il8/WPwtGt5Vm6oyGz9T
IAwq5hu8YR1Twcc1Hi5OUI7+nN1fFa46K3wPYL7HNbNzqrPZrbArSm5sUWHyhO0P2sHxkWpSz51U
1xgVoBvdrAiiarX1RFcI29pGNSwfYtOpn6wjZqQhkDrCuci/Pxik4PVMQSMG4wiSwQis1tLeipLd
rCk2VzS1AWFAgDHkKODIsAemIJb+oand9b9h7iOweks4x/LR18g9+jXGXjWTtamNUtpg8vOsTsuC
3IrrHzWtWd0Eda6XQM7mr7r9CAT+OKfF/B53gFBEw62NJWp35sYtv0W1v8i+HzdWhevAvpVG267L
EsUUAmTdKr2N0OBLTC08LrHrhXs3QZOuWWYkBhEu016TphHgRWoVz4Ah2z4HkZhhs1fwPgFDkdRj
GUxAiuoU45auH6NnQhZljHahaZVcpnXJ8oMS2irhiaR/15k88xYtcc+jdG4FIAOwkLrorofpFUqD
Kb9LkfxccerdnfiBbO5sIHOGXzPvwi0o5NYrPocAGf3dQp9zOJlJzvX6oPBLIoiEQqt+03JdVVUA
pkKMacSmhgYg7WPltZovLk2QOgVssSK7aJSqW52Dp/ZNzptYm5OuNZc2nOgnROlbvb1+vXPoUtIP
/CJ4EbBEFObYV8gJ/kWmGBeE3lDR5/hs/g7p7nvXKvaNr3HLILCXjH2R1oSDUcUOd10zo9CpvSK7
zssETpY8Nsyk5guCEFp/G6iUCCN9hZ4p2N8sqQ6o7Ikydb1qQCk3T4hn1pwhLJqF5G1/gpOPmuPk
RnKEEOOg42SbUx7h31gC79rVqithOMc82eT67o9jsIozdIpZEo1/OdIajlCe6n3Z34XTBkjv+1ul
T7taase9nvSBCftuEWTpP+nteJ+t+B+Hgyii4aQLXP+eazMTJxbE35TkqNJyvs+nmdgjb2VtPV/F
Px/zppfV/tK40HinZ6RCVH5V3gkzVKfjTdtyGYRR+I/Qvpj4p20u38wEkiF1TC8kQ0ofmQm/+FJY
cnS/TzMqtBoVB0B/zC2yzfraxbEKL8M6ntdzyYxiPbyF3Qqo56H1BoHJ8G/n/Sh6O1oosbx+fMlR
cIJw5s3U621/QS82Z2DmaU7kXzwiG3xmdCeCnhA0fH/vNsZygpoInzHIrF0iJMrrLD0Ui9brWF7w
hQRs5oh3PjvtK0KRhZ4V4/Ey3OkcKLj/kvoot5K3CoKrdhQNWkc7y5PtHXN5NmAM8tQTohSQcv8k
PBo0/j4/CkD+R9gSu7y0oHpWGtYn7MVFN/KYYVjfK5WHlzZbZEEr2hucOTfgwLNA+xM9z4cNdPQk
dll3rqg3l/AkpLgGaw7wgySr6EIGgLgHn+9m4XJKZGMHFQN7ZERGK6yOE31XF4+oRZ9ftd43yOHL
hTqUyMF15oC/U2hNBo2H/T2nplg0tFi6rU8DwLRKX75cVXF7vdGVK84yN085f3kqtNmka21m/jtW
uX/l/rR5T86877XDISSQx2bAkSIYO21jo8ZQU2zjDvxqYtTtEOdhoGtWAJGu7pgqtCdJgYKJ9hbv
hs2vjCJ7mn/uBDLymPf7/4DjLhv8zpMaK/0CvW4WOWgQGiZhZ9ngxdS06rPvDhROtNPnoTHkMtgm
PnMeRPs3dwF2ksZm7fny9wOOUxiHOsvLk2IHKO6xZbdAb25DXeusnGSKwrtkIi7vW5v75k90lIjI
PyatKW7ZM26C13TYG9bg6ug1p8kaae7BmAm5HPF5KgTZJRLZlxEvZO4VtJCyZbrkKwUwGjyfGS14
sm2iKunjKoYrC8FsiCUNOReXXIvSDvCWTyhItdWxvLMVMmaBtnKMbsyQ7oMq/tHTtJTjTtqcErfq
PRvF6YMoo9/wwjTvvAchSZoKmL56XMBixc8yAmd6SAAQXWN7p3UO698HaYxO6/BWP7LKVCkkh9Gy
xxm+RwQF91EWMEDpun4+GuNTiSWSxX1IQIM8RtU6PYjwleNvLueI6NDho830EHcBkXjGaz1yStye
lR1dv3qTfFL2wkaFhj0dYPtESu52JcpH9Auc7jGCnWKkloZOASVPxZAAstzZ06PpuRkXg9fuXyYw
9uXgXfDklqFvv7pydvkAUBLvpSnyooCB4vwOOVzvfE7PrSQeHiFI9gF1QD0s6AIyqw8yxNKr5e7t
octTk+5cRcg71jLUhsHAjuLIBFVqSGPVdOqW5a1epCEsWQ7vhSC1qlI4USnpX6xxYNgM/WX7/5z/
Dy2877g+wYVfZyuPbmErW5S7EBvoCwG1dZzqi1ym1REH7gaeBEOYaWdaeDewyeFmJnk9yli4kuMy
cZn5QQEm5n0DYCLYZqeTb5DVgL/y7DAdVZZlBGIy6yICDupDKAiIRnkgRpk3yuTFe7ff72fFFq0x
eYxttuaJ/NfdM9Jn889TPA6kpq0CKHug5Re/AOdG6G1gTXkVaZg6UDxuLMENpeoOQNMzF8CCE8Hp
Pi0kEMTy/s4DzzY3JlhVNoSOsbpH+RqSubk+B3iPgGenZL0sYFeNAlCzy761VfR5gQxWOybjRVzk
rtddbhm4LtlzKzYKGDq7pbtoL1rMWoxXPznsezm3CRXfXV2tPfKacRVhZXpG6E8Kh7jGgJCGmOXw
xUBoGFfem8r6f2B1nGf5gIaCUXrpdsyNgdmQTvl4w6Ij1VFwHscqu5wNkSsbmhog4zUWGMQKjm5b
IJ2X3UgC1+I2CVyouW0ub1ET/LaV5up5W+P0WtM/p3KLqiCJTBFbCwbs3KQxA9OBBX/O5IzrOo2/
F9Ct80R6famW4KNq3v5K98rIX21Z6D9bVtL01CsmQk/DJYlaLIhg0AEX0mz9lZTjpWnP+jAfWYa/
GnRr/kLrZWE/wBS94PYBiuzeSyEtyIW2N1MYAHUtvW0i2/6JE6G6P7J+TJpCwunyQmmpDew9VI2+
K3KRdxwV4yrrdYNZpcQXvmIwsx/nwIleN+nC8u7FdbZnhRa4Mts8CY3ItVN10SdlOGq0dd+iOqDO
3ELQsft/2Zb8gDNS9ce0PFgrwcyYsJ0S1hGxK7CE+Z02nW34aBZXnxHKCHqp5Qp6Tbp8wG0a6Myf
z38IK62JGdEEnaPPVBk40YrG6MnYU225k43WrHoXBXwODVf8f7o7z3E0NoVLQkq+R7gucS2ZKL6q
PwBbmQE5h4chdqfIfeH+NfJx+8geDOR+aklQtuDUvZp0u0WfgvTAWJ5YsZY8d3s8cBEn8/Hm4Vsl
dzEXDwMrCMZK7BV1j6ingKQv9sSMQ7q8pMGR7CL4RxlpAt7ldF9TExEznTiBmx992ZKMuznOlbhP
Fu3NIWbfemzTpOuNuyAGYBaeNXnoB8L6hH4EbQOAyf2oMpITRi7FzzTbvhfv5lD7YLyHQI5yQEZf
UV9YbDnH77+EOmMpNiK5vaIGGioWbNQPhMANxK0FExlMWDl9js0qHkfwRsP68TqdCJ17vawYLW5o
c44rIw5fRDiutJnNBjK038qbXmCt1bLY4bwO0IZKKdD7BHihruz3vh2SF9h6GIUdthk28pOswF7+
kFXHtem6UDmAdBMM6x4bDCKhjwVUrsDcKmTAFP9zyo1ofbYxpcC9OWQTcakHSkykOWgTdmbeZ1in
dMHLz+Vw4E+Pmhz2IzbRndUR3qFCxE7GKgwxtv3qqXs0zItwiUjhsB5/yb6Fn+7eBOVSQm1RBdXA
1gJ9lUXy4EUmEErrV+0RQF/eLWliFtejLBeU5qE29BZ0j25Uv/v3Lp+rxF2J0qVm7fWxS0WSBaKB
nSq2xhCB1d2ERRm6zL015fGtf27yzxTa8J8vDTx1aTi98MTmnDo6X6cAN/YRxH8ZJtxiz7sEp6QR
lZkqP2VyJO7xtOozJj64qSQzPGsHzTIEFF6yE1P6CEVdsPyfjMwAgbMWAMHmxJFHbmHxJAiamUuE
7wYqeRJTGQNHFPqhmOlNH2Dib/SCUKpuubd46wNvlRHBifChUGn+SXLkUjdL/rTXUNThxfJM8n4v
sqP0cboloaV5JnBfQKg79Q8ZkXabpDpjN0KmRiZ6Ny/uIkFXn2Py5+x/nyMBrRkRtk3lPaZI3fU0
mywSXfv6yEcfA518KN3dgvQoa3lilkHMgnel6iqF09c1DIQXH2rq/W8PQRrIk1mCqYLn2WY+IH7U
lrTk8VjXvGKzeoSfOsvehcpRVpak3GbdsJYYpX0WWa4PVSY95eA/8oMkTk+BPHVE+2bn7GzmUDWy
UyjnM/ZxDUOKGzqN5TVYjpE6Dkr+zE4wAvfejqAGoXcyPZyfcB2ghdX3lW6/HTPHjWf6XlRHAOa1
Z4+Z9I6vo+NfttJflfOu+R1CDoXkCrMTTe+ZLxPylZzESc5XNsk5mDbJqIiksG9sokR0FOfYqCjd
soSr/Doivz23b1usOes6Yf18cJ2l48ACSCOIBwo2kW9Jqmt5cGjlnh8ZDYeiisYBuJd8WGeljU6l
WqzXmQpTqK+XdFNnZupl8FJ9AWJX1pP2kkgqZrccSfmxMxvFHGz5RUAlSz3fcpUyZizDsiq/gJQ+
+E1jUwYclIlkiyo4aZ3AerBPTzZajJwuTUH+EOw3yFjdusHTH5B8lpIWDH7ozf9TkbDj/bGQdA74
bCJFh3u31GHr9Ld6XAW4zUYFIWKd5bdQ3bxYfLNI9rdHbruCPemvNSXFq/h/YAug2gVKf1+GLcRB
xaeFz82uH4aPzdAY73UU2PJ9l4F9w+3JF27xMrtKL7RkHZZ0hkSlR/v4zswqxigPgN8P1VBNjUKV
gk6Lcp3ykcEx8/42aKa5sQCpwZzAARnCL18ZIFFBo/rRwrk69RJq8m+Hv3Ur1dyWA/bfxHH3rv0I
nEzZIb0OUQuOa1NoiLfVW5jH0lAoWulqw/5fz1r1hySp2mZiDdTtYfYiJenwffOcG04spciyZeNZ
sCCaf9ufibLBkDw6sIvT2bQ88i3NIb1MsWmNCzZcoATSR0m+RIliyWuN5Zd+PvDowmxKEmN5xGuv
2QuANaSCIcJkhAPFcdCTKUkI8lzpOG5/gXeOgI48ygkQsZYvKTaUbdJAsIZU5gIx1JYyWNQIqfKF
pou7XNTBcbRdxBFB0USG5rgCY2et7Oc1QxHNs6J41BW3IE4kquxJkX2QdTGjj9zfUnLL7nOdI/w1
Rn+aE3GyPb8YGjqMAEAz8AJ5BMw8qcIeeEcZvFwhw09Rcho8cV+Wy3fLycSrVqqXzzofmYYyZRND
WH75VSbzbj8fK2BBFMWxFoxyommrBNcRPtzQY/HMyMakg2aG8z1/3uLP5VVPm3odRLqUPEJxg5NW
IfAisb//hmQ+uWVlM1U5AfhR+Sbo2/1+LmYYrSmZaykJ4l4pC43nCtKXkK7fb/cHvOSGYfVmk342
4BvlsY5SxgalPqk5KIIVOcC1EdKUX3AvSTWy01iFnbIlzkBNx/xJg9v1AYGS3hB4LMXBr+c2oXQj
I5iWM7ivrdyU2Uu3KzY6KeVBcnboSUmp+rCAo0ZdTFi+wD4ViKSG5uO98NfvCF7a5M76DNFczT8E
iHCfYkSvEeghnvflrPq9sdbZ6hZ9ouxcI+i3jWcdPQROges4v+qKbCqsgWl3KAjtJlVFD0flo3mm
juapkwQ56EfopYia9O8+rPq4h3PvgHYzgnIIeG84vrsvL6tCGMGZIdVKcmUOjf8/aQhJWWSXLWoh
XFnsX7f2Sa+/FR5AYkx7JZz5F1SxlXlvbUB+gXE5BscqQ6j/KfgKwHIw3XzaUrAo4UbkuMq7xZOf
XRzOCGOgEPHTmj91CidCq+bUzNMY50GFDPflmEbvz2mFn/8eykzwZCx5dZ6Q1V6+llEtLR/BmFED
VvgKbhSb6ZEGPZxEBZ0OsYx62Fr0csE71vEEktHMzXH6WP2TaU860Lj/K5xfF/4A6eYxrQhmDzYX
9d5T6V0bWth5lVjdzyal8rjM5XLVq9Hwpn2JKjCsOOZ6VNnFMm4Ag3fG9DuU8A9W5hv4d6q3WiXt
Y7PhH13fq9zY5KKrVWMhDOjjiyYAXEGoHZD8XiPsULoYe4GNKYT9XsDGztFdfZ6O7zI67506OJ8B
QsduXejBBmlbkw7++qxbWWI8KR6wpx4uZNOcDzsVt4iBZR5znHs6iMu4rRZvzIuS8SryTMWI3ub1
sSsFxvZcMf2ojrU9M3Om49u60wXsQSdny71DeWpPBmqlQvJZFURTfRYd4cIDdsjHIfSXMf6gV+Ts
Y6ZPmQuB0gZjc03n1i9IFEnHe1R5xG5rTo11srTg1zBiP7HqE8DF80Ps87DD+BcDDyYgXfeHYzOl
Nt/TM4pBSWL3/9x7EM2DRJhBQL7CFCJnEDkz06QzDGVbRZiH196oqZjE4Z0r/2QwZSfVS+D/Ozc8
PLbPU6N6nLPyDrKfNRqACYWdcpLVe9U8wgYkmAJAZkES66C17a6Gq/ko0aUk73XltNNeD1BXeuEN
atb760uCLW5WOEFQ5c70MqCGL4OxhX3O9tUDfPZ5KdL6UtGxPqolf//RQ2+7D6jNRjBYq9MELZ3x
Znr0zmu7vrLaOAlMKU4xWmH6tcixUQbVfl0+wgDAHq9HMYVe26+MFtALGN89RRKOjG/U6OJDJ7xT
oWXayDCId8M9/XACO9qZ58k262u3WGpUVnX9ssgWqnki9BLya16KCdUzrHueNiYIZRn2hAxe1kaG
c7qJem3VLwxZTsfLdqm5ndzzFSTZf4769ewmW/CiulBrZBe364Vj9l4L/2N3WVfuvfA/efgjGWuU
xGxLEbZ4AY7jz+zakELb3VNzE7tIZE74EL2U6udaAvzg/rWx/lM6USmiSiqeuS2rgKOPlCUWHtEh
uoZVgLIOwAGV5RW0mKLJutN+h9KSe6GTmbylbqatmQr7vtEL7UP7JdnOdtMja2vvJAnTExmZS9Hs
VUMQdlwxrJ+kIAkN392rbipbptX4abl9bfYENdBzKKWSJK4e3EiBTSz048+vMJkhR4XIdsEstv6E
wgnBiavbh9OkOLojr11i2gWlGPE8GcRUdjw9jZWgb1BEwkV+TvLT3HN7F11ccXpNzoLv07B9PgjD
YOkLL3CthyP5PxsODPWnpDB5ZSGWygqT7neR/Hm7RHz2BEu8xT/2Xq62J7rx0kucqT1O4UURjWJb
OOxxoD9R5l8028m3KHtTDOPGLFRnfToDG9oZVqDSl810yqka+j/vcApRzi2Pe6RXC5EaFb72HTbp
cNwwV+433G5CFjmUB5r2TpzGZ15qoK6/in4877rHGqDxnNtnSVHNEQyp0CRliGZPNdjXfXJGlZN2
Ew3JZI9O8DEqLl4Ma41ikHfqBvoxwRulxQlOzz0mO0xdpum7QFzcyCOnddKkCKXjNPrfltmeSbOg
i/KM7ORBuqNUGqpVwo/gGPykehc+gDetYQLSJSqjWEGuwl/+Y39aO4iUc4nC7YvEnIrgwnuVB+2C
Yxlb92zRj0ZfvL/xoWsTO1uzsjCeETGANPsbyRrZmkV2bhBIUiTDeg6NCal1a0p/YlfxRFzB92GU
CuQ22IUgWrbiGyg+TASTUmG6YF+K2yOItqZYFxIkaVqSJBLbnVsOrzBm2luzCUiKS88GROaYvhKM
2M2wT7Fx3w4qI+GNaMhzgamFgRy2qzsIEdahbitv4ADEB+bIEGG1m8kSZj3GiINcfb/W+Pf1u3ku
4ZU9sXtkqJQbK4J2Dt9OQ50/cL3Lfktpa8aH6oUI/LvKD5C8eZFI5DHikDiS5m+BgI0Exz8d5G4/
nlf6ReI9levKRauLoSio9tQ0vSziCEMq9Kyc81JuapV/4BsEcT79A7W9BHHVJk+1dqAJgcbhrRQD
li1kjO6T4frOIjulS3s4ZIFxiBvS+dAkMPM+hSc/T2a2pPC8JSL1d01QsyemeO5tLLAhkh71v22V
BRaXvVzlt5NUsql5Ia5xg700J34qFhIQQVrvjrTqfm8l6X8NdeZrzQwCqSQ4h9iUtiOZtG0y5XIt
ULoMfxZ7QWCFmtU4NfHctwGBPippjAIhbT8WefdChN+MALS9W2nDyM6bpa+R3xKnaLGa9CDHjl52
8NnJ5jN48+PeQGUhxUcGPZrsf8hR9+L0eLIE3F4xA8aKWTj64y30ceNsfDw1kiTxHTmorqIiTg5j
VEjeMeLZGhbujKD1CH+oQNdNWizirXrEVzGpYuoCoHLZrXRn0DbzK5jslWBGK7xkJNaFWUvNsAj/
7Nbf0v8Mj2DDr4F5C1X4jDGd43xC0xvI/HV9TnmQPqfwBYoLXh9pG6eHqHWRBgUa+VX4tgNO9gFj
lBNg3oZkBBFeYOLTzKztUtmkXSSLvAkwfRGQTTzHB0JPPhKhut9wNDyaJtLVfLjUSK/dK+ZPLD3F
LbLImxaiKdJQJfzJy8VH3u9NSkETO4G6y/omGSUKmSegC3yDa3P8skMlnYTKabAOTOJu9UQxBvJH
DapuyXEynlxYeeCScx3/m/bdf4qKlRNC5Dnc3z1xIofnetFN/+gpPYtMI2PX4Nm5IXbYWMuvOB0/
aVDhIPSL487Oz+Oe0nljXFE0LnSeGwagO+Fb+xXstr4xJddpaprjEKNgEVNxDQaITlzFV17z0RaH
l/KYtIiph5+EtdaCHqbMhKBgV/dPiJZs2t/KuDYORbIL4OAj7dgOTMFkZNxWWUlwK2ro8N/EuOQu
AQrTA4wteJ31GdaShF7MxkMiUHcgUfadEvSDHxVBOX9npGx0B86zPE+TF+E0JaCvsgLt+du6S0Gq
rE0XF/ocfn0kj9vnJMuC6ozmeE0gY72BtGKl642MNgtuhXs5/08zf9l/HC+d6tJ+sfWsYXE49lAx
XPSwWaEMzisRqXXlQPqc+m2Bhuaf+BbN8ep65xa63nfagg852pDRN7joNlh1p1J01FqGjnFxN7gQ
tCQWLm3NHfp2N7TvSYTSflDw3PQ6CWQBhgBiPfKu37uFwLnvq55qVoZ94iDuPWQKSisHoW66Cuog
qh07968vfLegrk2QlQbRqp8zA9MJpzX6I1qi2TqSFH6ln5m3qbcWs0wJhwLENhsxXIGKWGCbdfNk
WN+gqBuJD9AjT8tcHTfKn3TeCHy7FekNuC/PhOuQm0lFEw5pzdYiXiCwIH4StGYkvM2DW1NN7pBv
qzJ49OpM5nS4ShdOj/LCBZFKKLJToniqgJhIZmHacS2Rdqmy6YEY9OgzA4t/6OODUmzA9Oy+3VsL
jliLDoksqSVWHSRwjlPo2JOqdkjRH6FAcMcBeflOGZLf3eyZ1CThIdSaMJ60qRQsZ0w3CtJ7STj/
HLFWDJ33eJ68Y65QIqlFJy/4JOe4HE56eNuHptJ37ICJgTyH0NK/LrKtyavl/CArs7cwpeX/047L
P2KSnEo3P5AuCnAAuhf/AR3yHn2Iu82ejFiNXHg6frfhqVuEERe35xOURrOJegsQUE84Y50ov7x9
x7VF6Z16eqyrBBukYU8BCTLHOAah+t+DBU4sCG4Y5ZCDRopS6ECtqGhMJf3j6dbnUaTf/c1GIQSS
JMQt8Q4gA/4i9SsCaUfxcrqWNzQCzkl3C3rmIBafl3lebDU5JHWQObYrywMuVVnin9pB8oDP3r3X
/3P8rL+BOoZAso1Oy5Rn8/ZuVqINiTPqsY9fprwgG5U9W7+9DY/I3fyeqHEmpuWBhQIp1LMfK/XE
Dso9hW58+7OBfNuKQyBvy0Ehq6NcelHYpAls4/99cnWD9ECTF0F785g45hI9gQsLN2koei+xwYdk
bdwhuTJ78QWj8yPikW/IYTRIME08ia/FgJhvrdzsXG4B8aJBdnNsSjv8Nm6EYK1g4oE8k7tSu7wg
TRkwR5SS1D9os2DwLBV5YuwyAMpJ0iVBIB3oyUKzCCwtl3Skk9r2v7QexKomGQ7Ikbi8YANaGAtf
s8B4tS2GS1yz9EKS64Na5kl2muycA0rQVHi7gTT2t3v/yUBJFP3qHlAi2rlZphoW45grKRqroaUh
2lR06AKjh/iDqOGioTWSYdaN2sXi1/UzzNTERI+yHNCBN9HC4/n+tzBbk2YqbL/PI4ZasOzGJcZc
3YA0a0FalVZqzgj+9wHldpDXQKks+q+m8g5Rfd2LXdp5dTzLipyEqCWjCE9sMYi53fyvEW9NQVoH
zJ89Sg8N6GBVlqAa03Z6mYTUrBkFLYI9x2Z6heE59YMXdkInhSwA5pYIYr4u9mJcFdJ4OYWRjx8u
VpxNKmOn0Avsvllrq9dmaeyr7ReJWXRxM/qvBHZ3CJFr8kGNrImy+ckd6o2QCZgdoqcbPb1z/m0r
v4tC7ZEsab3oR73ZQrkZ98OFpw+c/axlS+xcxcsk38C9/SSzipb5msjOvlC6wBeAOLaApC8j9VFJ
gmqlzAuMBTdt03WGVStG9uH27RYNyQgAOy/Z5xio4Ap0UygXsjeVzb/7rLDCMZJy6TtFkpo5AXyq
P1kM/YWo9YxV4LfdNEfRrjPl+bWVi2bjPKUyKsMoegpfDUwbCLw7h3keQKBM8C3mHaNAhUJVYV6l
SN09hsIxCiysYThtXtVA5tlT/ykRey+fsCTSEUyw2kGuNDsAqfX7pWG07BcYU0jTMhABsZZOwHVM
l6PkiZsre99X85bYjSaB6a+ha1F+gXX2BIBYeuVS5Df+uxQsG+x3M5Xbimh6+KcitakWGoh9ePZk
aAdMxBNv6w6Otny4f9FEMsho3rEr+Qn+2me5JDQrBym80oY5gkue/U7MBAPeSF2K9si0sNvSFarI
l21WR01z0LjiUL3mp1WyNMuJDnCJQNdvoibS8LySMpTv5I98yaH2LLKOKZUIEF3+K038SCttjn82
kTTyuorp0VKRT5aHodWQ0ePDhhv8q9nSGjDAmZPxn+rudzJKgQ8NXeHtNi49+6O/sp49MZ3SqSYj
ITGSeCrz+DJPjxwY6KLp2aLqUWNHeqLAn2AEKudV7sEnnq4VX7oGBnbXHc62O0TPly1yNxMt09VB
g5MWBp5UtMU9a5qKbUAA3SUjEshu/7eAmGEu1WLWAeBb6bZluqSGAGlDpP0HCqeoO71EbRIPA6zv
s3xHWHACFZ3wZ8DmEAJl9ogUeo8GMjcJYgXriuVR2AijeGYiZDqhXod8zSUVeHiZWYtpKun6mEyq
nhvWih0LVibUQBzvdMK5EaSDAk+9sf03BylZid3HfcuzEs8d+YP/wmS9ct2ttrSiDax5rFn3QJsH
MLHdRt5HpY8DHK0zJVr0ce9GBeenVQd3oEnoIjFIt/zHeUrTNatJSvgupe9f7Oc1EME/c0gxsX1l
JAoYqZqcoJYMNGCBcr/BXmryvn6JrCoPhn9hPspYlzX+S0WccSu0++zn3VUOuo+pcfHuovyUlxPT
ClswcpqueXsBAfCoG2vBvQzInzq1b2E82QHR+kqhrw1bCL9yPEZGB3bfhtmizv1guoLK8wtVmV3c
BLmjDb5jMdXoBOD6cZvtpO19rnplqNe6qh9B2Fc9NXVuEZB0f/OgDFKTdKmI2ac0oppadESbPzNo
kzu6zydsP/bvcwPPI04+KguM1Ak59kI37ztpgQiRWqBCFFxuETA13mNMOpEHqA2em5tn4cN/L6mH
1wxRP8+Q97AWQjtlK85WmVzM4UyAVOGP6fkJVp3S9i5KOr/QL5um9sn2OtYLV8fVfdrU+RuxedYE
DsMAPKknjkCkNjzexB1Ldb16fd+EAFsSwTtTcET8TALMwefcAVgYDweaUKuwADNWIWE9FCXJdJSE
JIfrmjZ7MPcozvNfVz1RkK4s/95tavlWRVipkJt65WywXeqAPCHNu6bbut1j0WXjtWTUynfQI373
pWlJb1mPmBTjgzNmKdHcSrYpC4d3tK3D+CNMc34OXD6C9bG4avwsJsHJoma4VFqyB7MBrIEUSIfe
XQD2GPfywehnz1YqzXO5ZNlizjh3wK70b+JgJx4jZ3uuhkDx7z/0+6hujSO7XZlnO5w+ZvRGhPSL
n+Zo0ixkSBhW2hZeNwGzQMdn6nSRnZalDOD1zcnxH0WNN8OaAdliwvWWnUyKgmRQ9oGtHhdoNos1
AE8wwY7p3Rxg9GRW83WLW2VkwPgDY1AsgvYN/5EBwddAt/nIG7fXMgfSn+IMQ3nGV0z8CNoag442
N1sGSdMdLpu0rtOfSl7aTndIsNWmqAVaw4NW7H0s/E9gEy7UAQAXCgILYOvhva3TPER4k803h6U6
ZJp4hPZq+CYhkGVVmNJbpl2ajXGPI5dNx06OjRlMahQtnQWTAHmMWG5+pxzd6EaySyrCMVfYZIs8
lNaDWoSjuOslxxC0U+kD/dysFLRmMqHLi20ZoAS8q8EX7PgqYQWpJIFf1cC4bxCsnvHOFZLKB3ku
c4u5KWtNMo4rKJu6jFGKjIr1Mm5pSgUUycKpVJLxOtz0Bm5jT4RNpuzn2dIHaGrMwfP6rV2qmHPf
x9eF1FgolA8pCU2v1kFDhLvzmLP4uQUJ0F/Iz9Px6vPYIlL/rWzY7Q9Ls55lJ7IO4W1R7cqEg5J9
u8qcBY9bV5hNeApRqRnV/Xbd5nrQZXmBmIyB+zZhgcOmtmd88DFCK/H5JCEgFftxWUhMXIlYiCe1
iMw+2U6EoN/h1USKZ93lc7rdbjJ+5hjF9XVUj89G41yUPrS8oXiW45xBHHnomIf+xOEilv1yhzLf
izQIJSJzraTGhnVaCLQSbz42fMCJPK4hwqh+Hn24rbwjYZ0/yD+iwoVAoRJysinEqT68iw5vi0w8
VX19f+FSTIdW1sqz5gQIYomw8Obxjah7sYFrdXqGNa4BwmpMhd9Z+IUQysZiFu/PWpA0SBY9wxgZ
BINicWFfVFkXGfOCj+IyuAikKKx29xav8MRdzFRWRf5vB9iuRjtA6h2GdEPu9KskSctX6DGPHiHw
rBVWTxeeTmE1JV6PqBL23F5udy1V66kDhu+nBztb9kRVuo//njcOEBE6Ci4+HZ9t1DTZ92MU5lXO
VIQXxv/ydKKKdgfYKsNdmtZlF54jjRonc+2C7K9igXCySwuZYTOk2uRgBS9j8s12kIQe2aMkb3Ij
yO59GME8onM4r9vsWG6ZLrbQb7f6QA+CruCsQBYRYGwkk+6lNWoFBF3nTFIAJYKxJ0b1C5KC6w3L
faX9iW3ey1arZt76Yqc1Q9Ci9x20RjM+ffklR3xSwpVQKHFuykia8Dwfv7wGDWRbiXr4tBYZcUTo
qBieUQ43tJ+e3Vq/MNmYn47OETatl1zYLhjx9omYKVPd7pd2Zbecosq5Wsk+/B+Lcr9hOyO2nrem
1lClg1yIBge4d03/Tw9hAmu7+NImXn9aCAkDbz6YfqwdhvTC6q2c3MdhND/rT8iQWuVHLkD0gdf3
K8WkN2mBBuv6XprhkPy2TNHFytGBlaaT6ZZgwh28mJHYowmUWH2OkTAoAP2Aqc3p8CBaKPm3H9PG
/T6Xu4xl+0Ue8z6cuXy6T0vEamtw1+1PPvtJY9xXJ+V+JV5dGVijxf0OxNJYDV3uNCZHr27Lz7jv
tDjThYhS4l3xhsAZunGkXjtPFpDWLFj9eNfr6EQ/vf7wfN1rXQ3E1b/r+O7mD4YbP0D94xRHAdZO
UmsJAEwMdvx4bdEgd+hpBlWXNGp64Ke1HhMUpZ1jK6EJ47/qfGOynIggKhtDKWGLU8ZjxF7eDXXF
kwgOClyjF+NbzWefK0bAyIkeQDM6eiaUzq+8DSwppbzSEs5d2ltG6pMhVce+1ov58tF8P0q/Gxb7
SRDzZ1LZ9QrupCfk+iDzIhMcrttuOFCdUR8+izF41sgXVxwCE5MIW5emlMpJyTZwychigc55zWyj
M57wpnEpmvnSvm+ogRv00NHJFSfvFFYeVWXu4FWHQSe9KgsdSm8hcZgMoxGwamxV+X3/3JGrF7vt
xN0tlEVcYLzImmbwp5EaNsFNEyNE21kQ7CwNJhcTovdIXC+hGZ2/MVCYuexW2jhw+enofJtO+Clg
90URU2RXCMNyC14exKlmhTvCETQJi2FJIE8NT64EQ1xjd0GNMdPNDWAm8JHiiyfKxwmwn4HokIG5
vRsM2izBOHxjoctE+HHvD3UJ3BALi/wsO22/Na5E3XH4PPOUayhN2NHE94hvE4Emrlu+pUHOH9ER
OXaQWyIaKRbQ2JmjRwieNWv7rW5xYJlmwRUVyu3ev/zJM1lFgG54Sjn1ex5+Xn+ab6kB+fiEGNrs
8yaeN/b+91pRGK1gC601gZZWYbFtCDwETYlavLQYBlfZ6BRvjDbmwJFLb7swNzc8T1RyCV6Z2Ymi
jFv0jlQyAPY4TYzRJlt7m4MXTqKQyvHU5D3u6vTP69EdCdvHL1yP/pGU1mJ1xZrY9tCOfOwOirBQ
X+RXdB5TgyeMjQPl5AXsOerP4zSzZU25QGqOTT5fS/4j2MqKpm/MsEJSK3IOSYlaN+eFMTfF9K9m
4dsrBs/RzFsWPja6shws4+rGDbweKATwcNliPmByfdvvFNCnWqpSeOHSLNd8M2OdN+skvhJC7Os8
DG3wIp2ILuN522IEptvAHnzIIXre4ghS9otofxQVGF6jWcIc2WYYBOPRS8JCyOUm8P7GsIo1lSWp
6R+GeVtqYPOcKDkOUGZMM2uxNndgaijAddJ4rcYfDKId3pM1Zmxgs6OuZEaWq780o0SPrwVk5yYN
5PmuFnxMNHecc9AhPvoC+9f0T9mJyc6VfmhMhInqq6S/XPpi1XwWeKNWchAh1ecvbUnZ1QWx/1pq
VdxO94vFt/8RiHoN7SAaShjPGEjTMhSD7VDeMPwtz1XNY1GrGgyxA1KJu7eQxBBCyOlbHoWV6UPf
iCoszY1nVKFo8mi0Y8lAMVBmpptXNT7UsbK0i8KxGNid1URUiT4D1li4hYZZsySTS7KX3jYP8Nli
1MU+pT/pfzpjHKYKHc6d76GvHhRnHBFlsIoIr+HWdwIxpbib8Vo4vKPSVEpnBVHBLz2SjaUNbl1A
kXTJFyOmo2hB6NYgySCJ6NByBId27xSR48dy91V+QGmPuvynGnf2Jeiw/8C/cdQHm2PS8DeyPYgU
g5IAlTRh08OhskV4ne5O3RkwUsOqE7y9ASXnwtvKlf2UgMElk6avy5DxpjA/fZPdVVmSHrFZJ0dD
VoPF1NYIQStVTrmXVgojVFupuWcWVKRUZZ6/3XPBb9XxrCxvSQ7Jo4mb+cAZfiRYfg+6vd6FHvGN
XRy3/qPc0nOmokeFTBWIFGUTewVN97F2mtKDYjWm6SHjGuhg0X7Ki7WDw3H0hfI0j0auLOhSj8md
oa+yDLe0xfvkkiUJQNRzGYXWm2cxtIAvQR4vDZFtglhCRaM6prPx+fwPN6HOCZVebmRGOx7w4oUG
t/FmRn4L+OQ/fDElp4aNatZHYtfYlS7RS1mZhMvT0QE8g2Uz8gFaG/GC0i4RJcrS0XRUIljcxJFK
//zi125JWO33Vk1b8yxUCC+YaKCQ+BKicLa7xhSKPlqj8Qy2JR34OMmJY4AjzmKu/XIGKd1MEyQt
skyHldAcSo3W6csi3QnONbu7nAiUWEpa4F01P4QiYLnaShK+fUj3JzWYqw0+EBx5RbPkonn7fT2a
Vvg3CPXAJ9H/M8sAt3odFkVdXb8I2zHjwRWPhzNX37iX7FanveEdf7c/u5RZJYVsnEWMDH17wxGX
knVfQCz6MyAEjOjFgnjvFy27HDBjqMACQWtGP6t4nUtfXXu6hKz3H6HkKNj8jfU+U1a4Hisybw04
lwXn+12O8F9l4dUrzM3tGG2zGr6rw7pcytudUY1gPwT++wnUHwHiONJX8dIMpXoldC6OduHA5lQ2
brU8Bc1ny+ohHdy14zWAInobWq4+GvX7C0J9vwbqqjvDcG8n7v2W18XlHIKmIiroMXkKSe11/Zf1
pnU84TOMtD49BDL+SYmTyT2wFtfOYa/MwulPp/BxLUH2s0fMlFSeeI/4Q100W5vXUrnplGqP6fl4
QBdyEz/Z
`protect end_protected
