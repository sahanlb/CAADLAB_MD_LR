-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
r7iE/sb4mnS+Fz28qSdWaCX++h1OwtSYFCcI88puxRji+BwIqebaBmd0y0BNyEzy
K4AUHE3mFuW871qwzGbRDUkxMoiHSrLg/vH5r/MfGHFjzeJFIjjne52md8zRAaoj
n83xOlkXYutNP+VRHEtxc2V1CR9l8Y/YRV/xrFLctVWN5FhO/hHRXg==
--pragma protect end_key_block
--pragma protect digest_block
R+ENhUz2eTxU7jlyr+BjkCq1d3k=
--pragma protect end_digest_block
--pragma protect data_block
ZGiqwTor/QZKf9/5mJTVA3fyRgYfhQ5pNRi6ZHitJoie5/c/ihFNe2wu5XLbdkyh
bh1oxkmAKEb14e4zJAT8P3xL16yoNPHtPbgm3q8DdkkBlaFc8dhGDyexEtELpV+O
08ayRDue6O+LONKdRTbAekfJmnGAQKzy32lX9VPVLoFyD2AYHjIMZaR3vDkudz12
1Ye5g0LYJqrbPzLzX1DVjFRXKA+L6l8oGRcsAkcEcPR3GwLK5dga84FER/R/9Cst
CXRG0NbkA0qO0bIsq0VxQAeI+yeFTX2saZyzES44W5kBwcDpkNWnQ5L2nPr5lXAL
zkfU7/y22wB5v8KDV9jJZyJFhU2k8pziuHin0GAQV3gfbykHUFpuaZksiOaM6dBI
cm9xxirvbmETW7cufgS5bsc0IoAEeESQ6Z8F1s01iO0haRgJHp3Mc0acbjoKgWck
6jpzAoXUeyR+vKVU4fX/2IMwHgrW/VvtNvXCcCcDh9pWf4D21CfrShCFvoEpndF6
68vnUFd2T2kyEDEpw1kl3OPl+7VhwIh1J4qXz0n/xo1uAsXqJrE/KbiIkWXFGIaF
flllMbBLtgVCwNYgqiS93Nm1SPg/9NlyLqIjJeCN+MWl/u9CBtoXF/FTzYSd5vP7
KKvResa5m2N3JZBQZEV/3zyTzyx9OsOnA0hwxbg66VDCpSWMIknh0PDV5U16pQbN
awBuCcGzIuqCX5PLJBZ/dxI2hdvZ7RIJF60tIcRHnb4+8UEIyDtxPUBUAb9qi6aY
xxC05lD8YkYJV1gHXCR6oa9ZT/MJQBNAJo2SM/rpHWtsF9diWyImA5CNacuMY89l
rDGVYj5vxXtgqVCqqKjJAq8aU8u5zVaweerNAQhpQHqo3WdYJNSyvP/qHNvgxq1R
egDDKROKKOGCjQXWb11x0/XZex/jrf11clkBCwk2MgR0Tb8kCepEHA4Z8cXGOFJG
Q6F7TKZh5gqSWdT3P6FgNA3oRnpsdhmzG+8xg9cMc7EmfTe+oESXSRzkNf5g9ySs
gLDrn8GVZ5xF18vBujqy3/PiRebAe0AZOFgOtdUCE10muMI8delx1/gh/2Z9HDpE
NHzR6YRdkEdDiCHEuMxj65S7tgR+TG+YU4cMJmXyP/QavDtxPRXUDjESp57GT5+i
D8tvN8SdeJu4Ly/Ic/BeAoPuhGLvG6ZW1RKs4etKt2UKzJEHQCraWDDIX42tMh76
8Q5y68+ZG0ICdAK0ty37vOrhxRaGO9pef9eCEpA4y1dNqqXcTe2fcN0W14fKJLLq
tbwsCXf5mv5BuX7xV8E/UvhHn82h775AsHz+IHCyH32SJ+1+m1RjTDRSvMiEmq2t
2LPrJ7iU0CjJS3occYI4snyQKcwvWXua0mZHXw7k+1cWDXgwX5mPVDPGs+hcDy/U
0B1ovr7BuAg1caflANtB3+2WUsyzYXIEjkEOAAritkPpzZZnwNldZ9oQ5yR/TCyY
cC+quwPy+FXxymLIugmFyycFJAtR3zaYeMZ5M+teCQL5OfwR9ozK0gqBbw6NBYIK
hipnG1qtyXF+eUbdWWqjTyoffVngY0NWKrYU3PnnF4Qp5OBQmUmHK6ZFK4VPhZ4O
YPBa4SLULgdAX7q9jgfAo10CHFOTgAHX/KXHVkQNDwxg3cKjai5cpaZku1zerJx+
w+twn/FxxpSZ9pddw2THa/YpRADCsZejDpesn+Kj/pqITFr/VTlIuNgWuvF2BMLM
TLrHbvUz9rMipFXL7FmxIULctdBt/KgPYmLepHOXIV61vf2g5HXptgYY7fNORh2F
rsKbFsDnEdzaA0/CMkUXKb/YJ11uIOW2RPI8+3AVcGS/bUZl+3ypgiRohibkIkoO
ZD/l4ma7nNyzVmvUHhYppmkQZLSQl/9Tq09ucfBR08qBFe0T3QblIB138QQxdvN3
lKTqIYp9cg0XjGhvF/sqbW6qUi5XX3qSM1Ch7PIdfayxdl0VIi70y87jtsGIdfX8
6wm4TjWotX1uSS/33E24tQ2S2dZWsb/qZeWEP1lEFQhEWvibLBujRxUSl+f4+Wdx
g5yRdZpSsVftcxu4V+2eqJrKS/HZXT5Zg5O7aiii/5n2jb+9GuVCDoQ9wIiVKZjH
RpcSCoe/+Qi1T3qiW6eOoMQ1NN5lSUXNF6wEB9dwXugBX+iYSh7nlwctt2x8NIz1
dagbke625Xqt6ETfTZm+uYt8k7+epI7XMZxLI+QPt0Sf0kLtdl6xEfirNQ6fFUw2
++g4XrYpDT5iiO+iyrpwT/wzXdNBurtBmSlfdIn4fjrR9Fa8kWLsiPoVKWDOUCUO
FlSgBQe0kzMrKq3e7Qc3NouRUcpSetqQZ8GeyWQVj8IVw1V3iKhRjAp7Hng8oHfh
BUxEO9AwDvSforCh9jesC9gOtNBQ0sTFtFffoCO5CU3TF2p85FxvD+wcNjRSohge
ICoWLNYf7yR0ar+8XCEhcfq3jM64Vuf2ORHYLpnLJP+cWQOXrVumjtQSC3e4PHBE
CFYjF0rdYoXS0chAYvLa6JUdrvkh43dO8XULxYfD/VTw9aZT2ED4GdqzrMpxmR2V
g0zxinmwz9tyKtxwo5WX7WVU5q3BPNc201lpagveyv5K+mDrdTdNlDSurrwKnyVA
j1WWWb78iCIIMucdY2eszxgL93EGZzONdY65MQ2VHZMOPOuBS2UkS5dojkfU8MVh
ChYZPPOirM3hMdspvRtbbTdkTJBwoZXNl5B9hcfT3VvZA8+hokz0kHwF2rOEnsY1
AIwKD6I38Yd1s3ZseMozDbaQY9ezJgUIs8vIOeZBOcCgdXY0NsZfuVsHDahM58Ts
WGhEArFgyhGFB8zbR9FJApR+jrK4HwbfywOb0VWwqxpXC+Boh/2OXZqgnHpaMhXW
qdbwW9AuqARrf7YQOBEgIEYSy/dDXXNkhW90uztwkabXve2MIRvLsyEDZ/MQVyZs
gOdQMI0DbVykwyuHgBZZAExh4pIoXXHJC/VRD7tH56cPh6rtaqJXrisOaD074v3c
4N7q63TLjmojt05XiwsWUUQquM5wD6TnOsgPkolhsmnITWZXl+tWa74j3V7OQLtH
up2McatrNJVk5B3KL9YRyzptKSR09FxUlT5lNSqEsEBGj0l3q1//RClMbxpUbok7
z/vi7ZxM9KosE+pIT2Hbcd41ari3qfoaTs4GGk+Otv+wwJhvu5FQkUGDT/dO/KBc
gKaSA+rK5GbL+TBI2B/+Up5birtEQqm6vYg2lCC5CsoyaBG/1yrPjiBvaiLcZ0ap
f8fUSrCz8ovALVQea7E0tO/pHSL3sSQ0oqijmMku4/5fsgDNH3eB5/dvIe8EXbif
jZiqqojidptkcvt5EHs0UrkCNij4J5593/RjHUqUud2hYnkL8CR7x7ECZa72xs5O
ZdRzexk+1ElcL/EDSyUEs/YSlZNIWruiJ3rus9LhSR9K57tg0b5K9mqGEyHjpQmE
40hjGtKDl9O2wFb4zvamu59euDHSclgSxFL8hoe2RUQ4RZAbCkrWkcWyzWOZ/dTD
5N0RVef76kKHSTxRSq6cc2fmQb1lWZKDw+NNu3RJ17DxsWSAWvEpnPj1fR1BFyAE
+fP43AIbcaFSwAtglu2pl2m+qUiHj4osfZ4KrzRpvqireRAuvg3LUtN6YAsj8LSJ
/alI5JfLrUNz7rQlnl6KjtOTd1ED9YZ+2W44y1sg+ECUCCaArKY31FZTkKtjQzMi
M7Ze2cYyZpBCL930/9CkdlQvpVp5SqrFSckynE2oChTw2POfr0cgxgxO6j8kWsZ0
paugL0bh1tI0pp78BQuctmbIegP7VKdyIFCsD9wVv6V9b5EUCGX3saPmiMISt8YA
5K1MFVCIxlcSQHMYRX/j502u5p3+7YCrpEIz+ot4NGfW5aJ6l2gtWu38jvpj6iyk
J9dMgDulxeLkSg9msQPMTSYbi6RsqzEt0WDSV2Z8wnHbkN037ckI+bI5Y5yIoGMy
JWmCRMPUbUqE68b8QrwBwSm1wtmB8XvpKie+HGhAI55qJVW/gdGU4U3pjfGBBHAy
DERe/A7d0RZhKKg2ybwj5oOgWLT5g8Wz3ZmYjLA7WHJZO8hVQR6PKsxdQzijb+49
pPaqMxxofCMPys52rHS+T543gVyaoFEQYBJPZkfw8tCg1Xmdv2YNBUTWdriWqyr1
9ljK2yDytJukyd5KBqapFP9wVpi5vbSBiJdhX2Z0BNIFBa4cgy/l/hMmiwLNZz9l
GAaYL/bgjvU07IBmhp7wop2AbM07/aYw9CH5n6fH28tyNMeZuCKK3YILcr671Jcn
SEkClk2XcsRzhqRTPd3qbSz2c8kqyhzQP2qNYpLtSh8kEz8fBioyVUIQjTu1ZiN1
QA+yvWmPO+W9/YCdeg16mVuxmDASmLovewxd+htYGUfjjReIK6ffTLPIJ/uMoNhH
NIBY7qhdF1WmL7YYuoC9xCYN6Z9ZOjopfdGzkqsKhw734NTzPG+VBkhtUr2PTsX/
+mlrF8wDZgh0Xk/iDzJX8QpbVmGyCtNZ8y0sD+4Flnj1Mbn+xSufWhkjk83y/wQw
Q17oFiuGQYGJL/g89xdjpeo4swoOZXOtFA8wMqtT0X3hDmBJlLg9Rhpr1Q+3nMWY
YjTrnY3AfacIEfN3DGeKBMfGAtS6CetmB1W3sqDQoRrwZvS/zPfgQy53jgdhUs+2
zF0bUT5c9ccnlrYOVUvoTC2qma7Bq9ldIQ77M97lG1P9IzOl7rnCwt45+gLTGODA
PqzhP6YtvN1gZv5SaYgd7RUIw6vbichjqpf8Hf0fkuJvbIZUbBHw4cM/CakrndvU
ODpF1p8H5noE+qZAXkKtqHor+pgu9BecT4dqMfeVVdSNpc+rr9r2dHPs50x2jmGq
pg46SXSlv/lCxzF4Pf/opGsCtwNEGGIf52YQNgG2rCa+FXi5Z4d6BwHYlrEx8KxH
xUojBlKcwcnCHztdFXixycYMr9sdNsDyRZwMiStV138uGR2vfQXpVo09nA8foin3
r5tJ+heZoubYRs/0wy9MKrKd4e0u7eKq8PDq1BavkyARCWAlG8L+Q/iymIxxXKqF
/D0a0iBsy9PcvFgtw29/uU2CuM4LazIpLL7ty0OFI3OR5846AkmVIrer89nmhluA
hAaChlb7H+m+s9YaX4L2T9W3kZ9XPMtIEGfT48o/NxuArvFq3N5LQKVxBSF0Mf25
+PT1OGHDyTia+AvTgZo0dDx978NnYVEdz8b5/L4/nndq2dPw+30uZCat6HRhViby
gA492Diw173s1I0u8IDHrkoGg4P0PLsiRUDnjYavCQY9D6IdHnG1QM8obIQ4vQEn
fjD1UKk6ze5qHJRyFiHD29OELkJOffxSkhr/C2/VU19vfMEwMcC2HmR0OedC5Urh
ffYNVSQEJN7GsfoKcmm/iWkfUgZBLz0Kf/xdOSKAZZ/NjW7sgrNrMmqXbh7/UDIl
JUUJsLJy7seIwDNhlDKzmtpjFdQu7/b95zbOkh9I299nynxCMNJxsJf+ZamHQkcQ
avEKITK3o4MyBS3DipyHGFo0QxeY4O3EjkORlQvwWlMyhYlfwVF82Jr6NY/Fsqo0
x4s1GsBimrUwDPFvV1kyd0mVFA0FahMbPMwI47iYFzQ/SVzQwa7Zhb+VJ8g25PMD
dDmYyxnOzU9XPIeyZndRsoW5pj0YLEtCr0UqS9O9chNdFuAdPu8qG6u6WxkvkbVb
XRcbuCYBueAj1hzpsTOyqzlG9cPset5XWScdNCS5M7oIPJ88/Gw9471l+tohrvrp
WerO/SncwGym1d2J4+af8vGiwWjwdNi+gyu5oI4VMAibbjjNN1u8h946RqVrEOXn
C6rjdI5SRt0c/4e41rfsIoCJlArB46yq5De0TIr3BRNSmDORWftRjGRF7tVpZzoa
QbXOUFvLr2DyRK2ArZ4gXDFKiirt7s0VGzHo93eSF3dFKeUSduwbHuTbDdqQtQbo
wQ457r07wieeOQ5MIWXGyI86G9oxP4EoU0ZZJ3V5twfhoZKi+aSitt6GQnttN2mM
zUmpcmw/AppRskvuuuGL+zUs5fux/3YG8xz0LYELzFaOY1+QE3NeXKjBq2Yscgre
jnDQq7A2DdPRxG4nW05vJnTuUTrDlafrOm7BMxdSOBzuPEq5DB4HussrR6FM3Tbv
Vsy2zgKu7dujJ7qr1ns0BKT04bS/ebpg8auWJl5iVj5Z4p6KH1aG+eCsgySPNHSQ
EmcD5FUOfdzWqprsouAm3lsxkyQn0a463FxRwSExpniCU1Asv+UdLJYYwtCXF7iQ
QfXBdtLVjoBVmWffr480wdqf+qHLuGlr21/bgm/Tsjb6BL8fq/+VQqjKrkN1N+GF
iPwZK/jme4E26TUTbYZcO/fRM6ypQEgU+3BJXygCkJCwbg5hIYxc0pCp5dzOIMTr
46m/ieg7wu9REfh7sBFeqRpmzBC2L+tkr3YySFs3q+OTxUgzihIQ+n63roAH776I
tQTDtzlv/LCjfU6kw5GbMU/eA5UkofzMnqZwrxeSwNiIqa4HwlPYv7G2xUquIDsO
+c/6OLGk+uNvgx45UPJ4uSb1fy7Ky0CAZi/5eni2tffqJIqFW0PQNA3nVLSdWn59
sI8yWUz2wIfz5RJsRDo6xlBH5X8cLJ7rhsPebTNa5sLF30G0puUKmIY9h/ph2XjY
8ABLfZkqRvZm2u2wzMLD0feCKYos9/vCj+dmB4HuykoO5JYXsC3ygEMNkEGim9hI
DhX0FK//ieA5i+8iRDjpA695Cjzl+WzWNGSp5qQ/kvZGyPBnQ+ZnYHk3ehyW4paG
HxGRDAkP+2NCHxSqSpzgbnmdIIsN+wpHRpbd0EclvS3FvPtUD+r6twE+xza5F8QS
zNDY2nfHDhsVlQA9w6c0H8qDXkZZfk0gdPcIhlCZXgY6jiElNrxsEadyPBGu1sVW
zYmhdR23WUsR1RZ5DH5TcPeIDxxLCtW013mdWFJJjQhDz5A34yJA4TqU457MnOVw
pgzkX4KGdzVFfl8WE2ciDw98M5yNGdhH5I0hdug/UUu9KOso/Y+KEmKStY8tdJnh
p2vWZWytBSsD20z0nJaCCOAzKsPKKlcl4VniH85Kb4Lfdu8H7NhrGEXL3LmWmhXp
sV9NYwpSH4IuUP66VnlB96b63RgkLIPxWEGQc9+/2glhpPDbnEzwNyDdxC/Smvuq
OrBkzQl2+fvFzVdxDSXfCS+sixg197m2MGyveYWYKYfb2dNE5tOdbgLty41aMYP5
MMJInNjP/eAOs365rVCBd19Cqy0h8X0HzFZERBov6l9jg6Rtqu6mDtfYGDzjoHm4
TdKvMp6IPb+G1n3d61KbK22vzac4NbjA0zE3rhDY6CBtRbH7TQP7/CEyFoMVbfX2
3SUq85TLesKyW41MVWOUzjhEVpMayMBPwONeyL+/WWAEHrfl1fhnJvWmuQnLoSlF
ZANzwyYV0AIn3RDX7FWgcGb/82fy28qjVj2YKUWzC2a1+6S8gOVQrm04Y6b8kuPg
aai6oByoQl1gEOf00LWQyhO41x4B3vXuKx4TVPExrx7zytO02IsD12JtiTnzT7E7
/CVF1LuxotDzl9LkBYud6NCSb6kVQFbZgRYtWMCk2XB+nmo3awgeD1WXvfzClxA3
57Yv7ruvUtXrl3nR1qJsnaT6yWrkYnoLW4gVblaRYHjsl7Pd0oy3Db9teIyrUkr9
N+qNxfOv+8rbzwYQ5cSOsgVpfRNFtH6qlPOm7/XiZHBHWNtGGqB2jevo/5T3Oc9o
QTs7A3/l6nEFKfScjKtlgF9nm68GbPby/jzMHSPwXvk1AEeD7gQ48hUXNpgs+ffI
YW461MLRBkVxlvIkjMR4i+queQB9bSgw3HHAqnp/Fdc=
--pragma protect end_data_block
--pragma protect digest_block
K0dQSr5m2J91kWIBiPfCeAf90Ks=
--pragma protect end_digest_block
--pragma protect end_protected
