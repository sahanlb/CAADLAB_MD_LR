-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
M1Pl/L0XVJJ1Xlf0jqfRruD1nbYGuNa0ppi4M7H0ibtEjyV3vRGtdCQkFTfO3CKR
5rLJICBVp+KHBwuBmu+SPcerJaYZxQnsq2Vx13eNfnJM/mdJZ4uBgcEzoBoApG0j
u+WWFfDeGkTIzTQU0mr/03gT1sBkBwlYwQyI319QEAY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 41962)

`protect DATA_BLOCK
k29Pg5/Mk/mS+Nh+HRe2cAhZ+i6yIGaGRecjM4QZo8mKqyK/d/dL5FD0hCESpUyI
MMkkoOBGERpD8QkujbCQHgkjlqD++Sw+vSjI7BLh8RxNep4Vb+prgyfItoKV5eH0
hOVMEg1pFR3NzHask6bOLrDAILcGYaCihJIXN+A7fnJFkOps0ZFGD7Iel861ZOTI
g3DF+jxhj6b+k1ZTFGR0xrJnh1DMabStQaMiG5pg7rSN6TnkN3QOLlAnvi+GEmyV
xFq7wGUaPqCUaoGlEC7m5bNlYiTpCK9GAc4tVeVpNoXXxT5WMT734xr5nvm6pM9q
Xaejkx5FLDEBDpbBGp8MajExDxNkQAU6B+oSr/yI2j6LkPyas5drBA9ozw/I0O3+
h13kzf9MHjbCVaTWkDSb/S0QecRHeC/Ort5FXoOdxKZTeXc2cOrKMV3kuqssa7a6
qUNhL546Cz5LFdW1CIsPc+hJ0+WdpsbWUHkZqo50E7ia7vNCO9WEo1V2ukuancXO
ZFwv+0vqnAFEfEquffObYc3fmXsyswfSvB04a95X70jmtIetD9hQGvgaTlrdQRN0
YO0gJK4ol6f7XyHHOqms6JnKttcG5bOH178C/yXV0iiMbM9uaqLrY0D8O+s2W3kQ
itktvxt9XnqhDN1HCnzPddNYOTQvqajM3AurBWbMyaBbHY8U9CCRr/ncTVLwuASW
ewGuUBs88ifWX8ZItiznf9XL2532O4whvxvTQIMU2KOzqvcGERE5VF9YrTYaWlYt
vK9mb3tC07dViduzx3t1YvyvTsIKAp37tq9BH/AD+6UgQji42oZ/dOCPtADw4Vh+
lCqxCYhlyKQcpK7IqPAY0VrTNEDcRZgopbwrJ+MtwrlpEXhpG/A3zF9I/XWTII4c
OJ40YhXsile4jqGAek3NKsUQs7JH4CKeg3GnuzsqWVfsieBBPNoxC+x/4hRFyQyQ
G1+xNsusxoaF/1F4pmGhB0G6gD0TWPk7hInxSSk+QlXHtIzmA45jDp7YlnmJosYS
3uD9eh/n+QSzGMlHEsgecliz78h0xm+LmhW9cF2FIpkLPRnZ8KUbU/4ERlYqBEHV
JCzYA4LLnDFpneoHSskEBjxbbqDb+dWSCJCSy72frC6cKNlwKcb/T4q11zmzFg/d
j6NeLr/P+i8AGrJZV5TBWmZEGCq1AzlG+xtjBMq5ewaViN2nYFyW95txr8/J/YCG
4sdHXvtLGy8sRt5/xWRLQZvt+Mx/3URkdN/aXgdVzpPXDBaMa0PE1JvkcbPVvjjO
fLL4JP1S2dq2hO2cgdRtyq26MQRvHwZqca4Cw5dbcJewth8k1ZkWzD/u35sEGgM7
Pr765YOxBsxC0iQEurOEPCp5pP1k8NjSX3W1sdp8c7VXe8MNlmNu3lu3TlJBkdqH
IcEWu3cwmRaHOWP3B+352FqDqKyOmFzNlPIDt1LSUurtyQYedvbetwYg1rvpLyVE
QWg89l4s6cF8aHhYeT82+Xc3Ecl9meKmMuf6nJaYu99KaJllu8/jCF1MvapNmtJZ
EGdMJWZPS622Ls9ndrfmQ3TmOX8UmkXR44yQXu4hy628n8rjwmT7LlCyEGZM16HV
bnSXQiX7M/NHAEUmwPgHxpxUKZn3i0FbLbjXlmXWaQs3ssa34Iqht/w7hbADDjeI
s1QbkASyvHkufP9NqBDV9ZrCQ7SMG+Xonr9ylKynFSNbQ4ZzP1pYOJx2AkMoWrn/
WXRHbLVg3PDSPqIgS2G7K4pyYRRcp7rxo21M+oAYwCAIfNYSqErkqSzlo8AOJVUE
QG+2tJAAmMJ3+mrp8EMjK5x7BL2niEqZ/C8l+yt5Iyk3EDf+Fh3r5qXr1gHGputl
v039/DkRYCFYCCuQnqBGtwe06aCyMZazHOiGLsLec/SXPCXbCO4MFLRIjSTEGEeP
9ep5ZM1vpndUlaKdaVCL6bTGDLbfdbert/fa94a4HCOK+XiwzHy2iGdcD2yPvmgA
QyiAjSyOJkFfibLE8jOwiH4Wp87iVa5P0T3ykxc0SRxGIPSRAH1OaC3d7N00Ka9m
jSZvAyaqFJ5xWF7oEbQVz8A7DDOhxyhTAWjoguPdMhq+nVptzed8W7KVliHEkRBH
gqwtxaK+J9ZMLq9GFUrKnX2SIf7V4jceEeZOBP1Pwesou+q2LQmJZTopQS0Tn9DG
o7tr4j+NqUiAVJp27PmBb0D3uSC1hL8qzfjpwd9DuLQ40F9pAVedVpHOp5dfAmO9
rqkDUwGjOPxbjlGnU2GH6mytUFdG0KITrGBt+UJccADv4W4sOwnoHS3ehD53TcRv
JdXB0CR+Gdp8pc9DKzidDL4xSzNc4bA4159j1UsihabIGHME9DlN6sWhg2FLaLsN
VxmXWeKVdzRohG68DdzKDgTesg+4nXwdWI2bcMfOu5AbKQsueF2K4SQf1eyXqxnI
fE/9VOhp8OP/HQdWEINKlBSVzG3P524C4WR2b+oBM576ftL8VafT4cDmHICL+Kgc
Z5SH5ze6fiPHcdWv9wStdOf6lytiBGKga5PjN+AolIbggyDYb/2Az2E9Aq3Ue4J/
Xvb8kIjatRBVNmRhd+jeNURwgIRLK8N3nyahHdhWkAysBdOKGub6X6hXog01kjc0
WzmVDNPxxJygDf6FKze4I/tBi6Gahl+4D6V8v2DwL6Zp466L6oGADlEpqT3ZvyJZ
jTwUFRbrLqyeHenXkaoA6nFN26Y3iM7zF9+RNLBfIh0FJI53kPlFN+Dwm42+fwYY
ZB/OzVDjCws111CWJFHhK7DmvEgpDGotNkdWOF5fuddZU8eXm2c682psLneb84iz
cO+ZTQWbrLlYuVTywec1Yb+52vI+RSfmSdEhWnNd2k0Cg2K0g291ZfZkgmpn/1hI
QyPBQkIM2xoozbFpQ/zPZd6n8hHJ3KHzP9GbWHy0/5r9OEPq4YyCP4T038Zq2yZn
w4NYGpai35AtVZVFiF37mImh4m3VwMH3+tPVChh/F4Nss5emQpP9ehShxpIq8Xpy
Wc8+SwImSWVueQCY5wMoSsrGXaTLhSp0/8wZx+HxO0M1L3PfEK2AXh8Jr5nA/9Zf
rP6vLySFbv61/9ovimaJgt7EOiAjdi0MVXjaKf3wJdo16KQBSgk6y+TdZIVdlhfz
OWtrPxRjmb6o8DBucZVHfhDSHOfJ5j3Jw5ZluhvcUAfdVjLT0kch9yX/NYJxismC
9hqBnSozgN/m1Fi6NoQ/Mm9tR1VRFJT9DHbVJI17e71h5BaiUZDfM+amCV+QkhVW
+MqIomWHbvhHTfmSkIWEpGBEd0K3/2cV+lY8qzFLsJT6hCis1jNUmYB9gdC8RWNC
RMM+b+x2lSlDePWEuZ3MVD2GyTnoKOJPTP1YUXj8YMZStBzKLxWJmWkTQ2MYGtll
yd3LJyWUGtUvPf/VrSR2FLSpQjvi4Lut5zPruh0rcqkOpufhXIvOpgCDIFZw/1VK
mdJXNe1uA01Dk8QDIEj6dfybS6C5fSZz6T2pZc7hZVNnmGFShUAb+SHvZTbVVUo2
nYlLI5h1pLc1G4PzLFHYf2a7yc/2F4OZdERs8Wv7YUzpNOiR75VvsVpChbvGHovS
3ZKhTmMWArfeTDOdk58LPjhjORDuT5OSxNfGa6w6a9TAKB3DxcxNr2pXw1WNh7Vj
ugBNmkr6vL6JT5A7FvWEQPdvKrmuI20Wuw8KVRdIc2ppjuDsYCpThmRFrTlWk6Wr
E5J+TwvoWMb/sYeohq4bOS4ux09MH3Bgymyoyf2yh6XNqPELp0nK6XsscnvZfdmF
BHM9GvhuCU9Puv6DnPv79hWb4Z85/0RyxWbGLNBK1apXfdQaalw0IeWNIvObKHlO
6A1jcPqba5ekqMkUQdyuDfFEjXHRR/+t8LFkbDqpNR1Hy+NZsuDGq1GsVPRz7NQJ
gzYQ6vq8aZoDWkoAa5cqlYMrTHEyss5C/RpWtcEdwBWsya16iEwNzitQRpnXEzsy
jQpCbZ3UZTQ9jg+82f+ESAqax6yeHj0TXKq75cQhjT0xvWZe+Y+K6D1f0TzQDLWK
bhs/4RxkDlZkv3LxZjlKl/Ff0AHV/o8ft/RQQdvBcZ+t4Oe5RheSZUIxzl6kemOf
+K9zI3b1zpHwg+F14xFDorwYLrHHefqGVRViD3L3ewwA5xrJpuID9Niv+7Rn5SUR
+QM3Zas/McbsGUDeynbLD8kutigoScM8C0sKVDO8w0NW6ttpdC4ABMhbjcOOQKbV
jeEqkh/J1kzrkomWe5VRdaCTsp3MIMvd8xFt/evbyWGc8zc6pxIU5UBX0De31Xyz
JD9zbiaKXPqJAnBGqWvPzreOEIHXTF+lNp9la2Pwbd3ykU/iP09/4O3tYPzVmoBn
hfJsLWGLwmbzNainmLNJwd9ALjPym0VUV+Pa7bn9BcOcZPGoLWU5FHFlHZgpElSy
aEgd2cC9B7hVwQ0sDc83JptBaz5rCy2MA7Er31jgM9itDG5yaPJ0NH7DozVQnVS+
glD9Md5H7ryNohCo4xgbvuRrmQ7OMx3ndtwq0aS0wRC2zG0xVWrxgOtCkZoUkLbk
dDbEombN1NJTic3j8PR60RmaaZ9iOZGR2uO0jRD0gJ/aBiv/8hfHAdTqlHLjfBkw
Srhfi3wMmdnG6KdpCceIPvnU42zemRcTftC5WTgDhxXKmfA5y0n+AnnJqCYxPLIw
LtKzJr9tpju0FdP2W81xhdSCGJFkFG510RWIztLDXjwZhkz06W6bFoUJuIVgKlA4
LrTmaZuv8++smD8kdHn/5sOcFIbQ4fCM8j8PYAlLgfpNl+A6B4pRtCtqjq6neA7n
AYDh/HY//3eSy1izbZ1zbA22aOmWgJAuZP5UKK221UfNCX0RQIKuBZ07lCwkUTUA
0MQyKxG2imN7CPjaE0OX1KKUXBw+OUYYIR3K2mAAnf70M8z8mN4eNq89RP5QKVqf
bZoOEiWPEYrOpN9smIOdpYJiJIuQjmM1lyh6LjwrBV17PLlYcXMZwsdNaxKMlS2P
MPrL2xYXWYOpBbgh7YCU1kWqFshIVa5DV4yfTV88YRxEYgPBy5xdR/Tu7NsUetA2
RhzlsswukEnyJkzeOyJvgaxPVedWx41JdYZ90YuZM2YP1uczANrJpxvHE6X3VgKT
FpY2lTHK3hiIF37Cj1nghn4JrhlrHLAGiJ1ypsrxWAGRppOQVlZAU/ilJkJqexon
guLjXfjwVbax2spCxT3zXHnATkX2JCdTKbDth+FsWJcmXJiS22f+BHVwKUB3pcXJ
8K5ELansHORtBD5EU+8jO8lXFOxS+75+r3TJ/Y/lZzi6N7xYYR10Mv3jdZqZL1Wr
lrFbMXThWP38fwPKFcAPKpAhpVMcmAIqHOpO5ZMqPiNyntSRzsn8gElx50fXB8m3
ZDYdq90JxZQlFF+lyKj1CpHPIWdd8wygsmCaxMn30yeMsm3oG+b6Ugj/AbmVMDwc
YdhrcMhODrjVil0m+dUsbIcihxyvzGJAYbG1sQ/tOjmH5Vm3VGl/y3t/Aq43ShJj
W40sp0o+z+U/huDdCjLfxfp3uhesNpDHDrh76B2FbrMFq0gav7/vZuW8F08VuV45
5EP9DwKOU6Ds0qc9+FZ7/cNaKgxqAmxEm42b8GI0GJc5hkvY0kAh8/p50pV7RlIJ
rwW3mU5os3DK/2VW4bszDMwUQro+vgUeUToEpuy1wW8/0SnKj+L+Gr3fPmivmpk5
ZOfC4kh0p3AI4WQ4FN/zzCkTk2oiEEOPLBpyYU9DqF+d2O7o1Nns10PQSXrDzduG
NKw0PTJL3jPAYG0c1e1Z+wBIR3Shpok48WYEDynLEvHT3xbBOe18W/u/DySkUVZW
Eabjd1lA3ut/1q/FTvqZisCURA4XsbDdMM+vgGxT4e1+qArQ+qbYEMkkcUH83gqU
S2XIECDyHYbvd8RJ7wspTT4kd2LkY7Zx41E5LD/ki8YIpoRqLUiPj7mV4uaboeq1
uIgmcPtJbQl3U57FBTdBrqzT9XzUFsN4WLBLYbX6CAxl0RexunQyy9/xttkBVVHn
5BpTujdRkoU1scRNFYsaztPPSPmHqo1leordLRkpouj+sjc5L5EfZlaxQY1hDXpf
SH2bERQLwlfkoMBcCFym/ioJKcmKtDh36/Nz4oH7HaH5drihL1zUb4xR53pIWlwp
dQld2crAw6r9VVesWc0jCuZgUDUxDb5OrmAMQr+DYLkQHXydOSO/lVc9hXEd7fJY
Ed1KhHT3cCSWtwNdA+ofiDGUu5qyEIDlLw6XljGTssUIVMC3Ok0AE/drrZvSSLwv
8GjRLCvqdRCubyhKs2ILt4Rz5+CiJ7uQfhgoDae2jV3ChDcDvaKPqr+aWWKr4FsK
Du+s/6KSrzw9mkuOCB9Vfdn1007iVS3ZLfoQcvUZ7Xl/TXSb1+5yZgUa9UhTjXDx
5/RCc0HrKqwmq/RClzAJwYp75q55lmmHfwaDPosBKohl4ZmS6FxPafInYcERArP6
mI9C6xhz2EnJ/Jc8x9rxfLN/XIA6eS4lrkpTAeAmLv6yP1GxJLxzuXU9TDgW+Icp
DM6ZAxZWgV+ZhJd1mtP9DpkvFuNcTIHoDHgbXAxe3VsiNIbg81eTkJXlkSwnokTu
7Jm7a8zkoRPQl+SQwj80T5ETxoIS1KAowF/OZItChKjQvyx+MGoeWo2PlvuL8g3u
tJZkHYJEo1/vKEwIJm1oExsLm6c6DkgfCUswlZoGalAz9Sdpp9Kw6UMgIpYPw5p8
VRN2XPPvaSQKeaXuxMKUT8bwrdzo9aeACHWCXpgr7z8810j7Ypq432O54UcCBO0K
2gI09gI7SV+qCvs0AwN2ueC21Znig9r3UXcU96lfoSUgYq9UWupHvAj+rWQ+yl5N
b4fkXBWsqR+lUisQfhleOfOl5SrYw/Du/KnC3SMdGkaRKF9CMpYdpZyuUN8PjBJK
Vhl6wPXWLWc3EC+pXWIYXfOtibVqq4wiJJeUtWVHnkkea7XZLJDmkSSP1bsEevN0
cPy0wJUfSM6DclkDEHtsk8HqZHQTe6TF5oCBpY7XN5aK9NQ5e6BP+Xp8/R2Tsnby
nhXLIzho1PxBkQne4vwrpOc4xVi3Wt7Epcg5SL/JaWzblFyEW0uqFrLLpqZ2sE7y
uY0grBEQj7Sdo5wPgQlTszL7zoi/4ZO/gQZ3ioN3kP60SFLPyvhSCr0Zup6gYy+G
g2TRoRW0oKtRCx18UgoGxZ0J6WK7KqKCKFM1eyjcB6wKZlVL+pqqjSa/Jkeu3FOm
GhyrwV3rzqbnDuSEAts5LQQ85yEScqvXHmkV2Zl4dkqR7zhPNKsnR3ZPwZtDPc8Q
qTLcYDRsZFqO5DavD3ZYHUS1eJD9hcVYx2IRtKRKzAwfgTTa7FMj61dwTl28VjjX
lV62hBRF+5TmEM8jp423R8SiyQvIZDfOdV8IPdy6OVfaEb7MBH8WDt0IQ0DsvB8z
Q/2gkLr+Ell1jWDHmgf5ZrT62nSWcg+IrLl8rWtu1Z/x/gZifWmA1hZksg34f3My
bw1YbcHYbtRovZss+478eRi+1hH9JG5CilaFzZChGdKMKY7/f1pXMAgv6HC+SO/r
sqsXNyY/lIkGBU6IlEbAM0NMqH/hJnv1C/NRpx5h+xov0c6THLYcLI5UyyaFi3JL
v1/FJmtglVY3xXAJoela6W7jmxDyHLcLi1b/N29ujWEGvMgGIldTmO9ZFgFD7fwL
A1+pbutU5HrdudcDy89pePxmDzka1+Jsln5eKwgits+oT1z32kBypdF2jE0vBZj0
8FJkfotE9A9hFRZaiOpmHcVq4cLpi5KfYlUqwaB3gDvnu/ld6ikLtb8qhCHwlFVR
rsMstKCNz0T7k9r9v7Myc24X0X2fyX1Pecy/XC/npl74ClPBNfzOnMJYhSEEKi5C
Eb8+z6b1brjOKCvkXEF0Blyw1wV17TESTRAuK80D9kOoHQrmVzrZMpTr/FLcR2ZG
pEwpu6nYeNOxphGfMiiJzlzX2UpV5u7CBAwjUkXkVBaSiBrwhHZ6izLhs+1csh69
IeNMU3MTOiQW5Pcge/E55cF8TogrssSZKti2iz/pyDF9FdDRqnAQrXUFdxxg1y41
mIzy2VHKU5C0BDbkf2Txuuymd8TpPFyplGpqHvwwviFex8souVORYkUQCOmxFPU1
O2dO1FxFP4Ve0VWckXvy3vaJ1RXvyTK7bLjxfZSnRWdY0j0mV2Vu1oGWNRmvrnAg
rKykGar5y0SDW2AWWKU0Y1MZSoTbMz/Ve70LEJpjIE1mOq80/A8zLvEGRAEUbUgu
fkC4z69oGcBKyWdAjeQsPTe7zD3ZWoUl4OJ+GWucpkM+YIzaRnBPJXcYxBB1yDrO
n9jf29/z1rvEI7hYRHDjyfH1PsjBOech+MK2BZO+qDDo5uc8EjxlODl3yYSRjnwE
km/P5TcODWnRUHu6PbB3sWttExJdO0UazDglE1rxrS1OBkMBNBwHPpxfsZhSdO9G
iNfdiPylHG5STr8Usado+1pL5NFddRuRNXBzAuSb1Q2RwsRCb2RfokgOYdmKnkQK
GQvneL3DE9QIR8OpYBQFXjoX8U8GlmiBNT4+MRv9boN5DmvUA9dToMt4YDkIX/7P
8r877m1JrRGheyZTNfKmCF/UoCjnnIViPGi+bUo/RoXwxLcQLaK7Tt/ZszUzZXCg
fa0szDZdD2kDDlBnn0oQOwVssutjjl3FZhxmBxEjo66hsBwIhXInHncSKNCz5b6C
kfm6lwtFIfKg6Otb80R5Fp+FfqRS/RxKXsY/e/Zw4g/sjO3UMWoAoGYgtTeHJhSz
+rgE7vmvjp1bgIg5vOcD7D+t8mYHIaNhZlcWq+8nhtW5tcHXfYoR5q4cRPS5NTjp
jSunTqY99rCapiwhE4L6UMgWTedyXUUN58osHBNiVaN8nqVArMDRbevSnrpplNmG
3js30+NAq4CTU4ElDxFUumzIj2Ak1u1ATUvdOzNSB28XqQEspaI346IEjEvOgpVp
nLvDMQZQ5WULMSgOi3axTqhAKizvC16omUZsw4ZWf8uSYtJuDNMvxA7X7F+FtGJT
QeBG+CsqUL3W3tglbIjHBBroOQ+OuPxjoTUOE3FNb4E60IhjYEi++iTifWhOpZlf
nuhsOI8PQMefP0k+YiWqHidYskLEfMS8YJ4+DNrXLkRYQFtBYvasnY9CnxZX3C79
GcO8QfGkaek56WnMhTAIK3ZGinVdiA/bhgnwzAEWv12HnCuW/jA513oKMZ7h8ykm
hFE+NOe/f2bmRODsZ7VGEdhAF7dopN/93RD7v7W+RFtsdV54BurQSrVf+d6KCIJl
C+tGnSOOHNzFXKFkMI+UTGo/oakX9nxM3eITcaMupYYBge8+nex8BEiGyck+jaXP
afknEh0QJXHBeYcuTvOCMtEYBbUPdnVe6To6Xs/AJf1jNhBPIly3r3rDzxJWiHK3
pFVIvcJpzlRGlM9wuz5pPK6UP+V8eVGsiXqift9TXIn+GKy2RHwWoN+UTRHLVXQf
0uqCxxuwTzaiZwht2OVte0kRCqUY8txdRNnj4cwm1NKFqDN3yl4nNHz81PpwhyDb
vTftPmatPBMK5PZ+eGcRF2RshziRLVXqj6+FTCDaW+9RTCSqRR5CSzle2SgPTJJ1
YbLwHRqm+WSWyn0YMDr4YX48PDw5p+l8ur3LBYyNUSnJFdjSL022hodPac8om4aF
G6SjH12yhwtYO633KwpfG8xsufZusTEblr8i0BH6tj1SJQTEriQyWVnSUAD3KdLc
cbuZVHzFxOPycDQkKm5j7K+sDASL3YBdBAKAiLpSOA9tpxTOc9vRE+7j7C2LruUt
yU3ZZ8OTHQowaneY9Wsh64oUS0Vkb8BqF5+ZUwRrlnS9kHdAkHMtX9B8cb4BOl0A
lhtkkCKU8adrBdB2Mx7exNBOvKRt7AjipijZWkjBWDtjHFQDlGl5RBOeQK6T3HC1
/A5OX/dCkIISWM45CpM/ThV0cTrtpnFZgs/jRbonpDsLFtry33BZa8TM4fKaRNxP
ZbLbmSFNffuKbvUa3hFHhHLILY5BWYyj+0ourDx3RVQ4+vXytRNuQjvZBlU8v8bu
f/wT4xRLXCan5KLIRFG5brzkFwOqAj0oDU+5R4zmwWVgrrrbFkbG38eXmjkmQdid
3l8oDDhY7vJDSjWg3xBcZH04gYIuRl4GLYFbNQ9HIWcEkZ9ReFyidmSbfSffN21Y
gpT2bBeDIJdbdWdfEoYV/4foVURa4WLutAmo8ZDIxpKUURvCF/PG/XM1YV14n3bS
bDmy1LFn1KWgtRKL3hscOrL1WTd42CTM+3FUqwyqbLnNEW1MoGm/eOpXxywPZtkq
3FTIGcHQCcx7LE8FkUyMVazHWxwRZL+sBsRI0FYFjLivk9lRHdz5f+RLRfyYPhnv
NTcQtfEftjva1be5wa75tsct2Rysi9uzJt2LiEmhb1qxMJhQLc7HlKK1zTHu58MJ
dj8wyFb9gEgf7xnp7TqJnB0wQwKZ+spJRC2+eeA5qFgGzXpyFtp9emxvsFRAn5up
HFKDEzxKge2WJgGx5IXHVob7dDwPMonjvFV8UFYalj0i0hrPpobt5DMudJNBgx8S
r6gziLA+h0HfA4TEE6LnqXpOpNdnfU12yjrzhRW5dZlr/wc18tT3kmcHbt//skfi
6oMwsaPmMm16OnmFdSm9stCcpKtKgQnPqbyjxbyO4DChRFjA9U937TkT5iO4J21A
AuP/DtaxWCgSBIio005OHiG1qrUAa12Z7cL7rxeHIPWwk6mg1f8sL2IHHStEX3DV
LKulLg1zcOCXkPfZ5Fh6ttjHQOAhGI3lGTc/5MHsXEgPdcC9suUTnEZdGEm7osJ8
R1wwK/O/8ukNOBkH34gQWqut4nlP0q/b1+Vqx7aDE/o6Jhz5/O93YZpMYKZLVJoP
UoiEOc93y2YqHEktgW9ZAuT+WHjaNbloZ8tU8+sIt8w/C8J8vie9xJwDOI4jfvfD
mf5BEhBMSFvhMfcwfknP6Wb85PaqUgWw7fNdTuplz4F/KK/rim+diYqypKIEr5XA
Z2fyy6jB3a8WjZhIoCgtOL8EEbZUtY70AC/euQ1zy9ndQf6rKVHslTIKvTnckFCK
fVPM1G3Ns/Y6sMFDfowLSoma8Kpi6dCEVhExsrM1yFZ4j1zXp+ZEZkS8IRIUOeqd
TPZBOVkrJXYxCWTId8bkdmPWXE86bOLwOrRGNFDy+Z1dSPDJwO9R4r8RBGEhKjzR
WfVhNX8OlByO09A3YRDq/lfw6xgbbgYSKmd+DH72IjKDdTBCj29KXGWw6VXOA0Z1
5ct02ycgp5adn9nKFUOTq+zlxZk4MbgcskrMsFujclEO6GIRClvVcRIwcSJDS+JV
Zt6PA+mIIzxLKHXvcGbbczU+/+3JIa2EYL2cFeSchsM5HW4s6pDgmOaw3zOxFdFf
wzOLgfqklIuwVZ9Ra6m5aErP0Pi0Z6CRLYhfqjY1hxT1gih0CaQAQHgAJ+9Krxbs
B3VXuUTkYHVVG5j8R7HWb7Nz1PlcZqxPes2pGnp0N3HCLt5gAGlZa/1ZnLCuPp2w
ueOqx3X7xb847nBq/ixKH9zXmhmGfQgj8XFLt7iH0KVlAVGnBdbkRoW5mcsavoQP
fOs2UWY7NzGhtAnDFOhCS1F67hbjIB2Jl1VrpIMlt+COuqX3hExYmoct/+tD+B2k
5GLZtAUWzjDl5n8rm3wDJuybu76DLnf6zLKljbHSpntgnx1x4LSpKgRDCtRwjUaz
k/etunrWjWSOrMZx1PeB/52bvoHSalyvpqAbTm40e3iXHaM99Ps2KI6Zbc1QRucc
ut4V5LDiaz+DELTpz5LxghqO59kkUMO3yVJ31wG+8TztcVmcYxOOqj3Lx2FmVS8X
/s0FqnI5PDncBqG8FiNVhPIDHabUW0Weiy0WwkKqgqbgNT7kZgKySlyfOWeo9LUj
PlbCixWPOmwsO3YyMAErFbv23ldZ7vcngjaHUsBLoPlRHTgKoZ9f1K5dU1m+xroT
q7r9G0q8/Kx/yj/u5/1zMW0nyFVDbIyw2ZU4sNTzpOtbtY5PppeUjufozwa/RnaW
V+nPQ7eaQGx+y5biuzRnPpP3CU0YbrVGFO+mOqtbRUWRDQKHERSKY/G2woQn0fCl
lU0PkZCI+uo04L9DY2RC6m6lBDoveWrGQ/1oqzrE9ZduWG/F3hcGfsID3HyaG4+t
PpvnznERUGEvnzzTvg0kf29iWZJnPDT1vy1GRjVcaUoov5tBzntpQrtjpswMbD3V
ErLpUOndYRlGbEyoLBhRzUaKJBZYncANOntapPhrh86rJAVMzNy6ZiwpEYTpduys
2qtEyLTeULRAvsRtV6Icx/CvwjjiAgLUMErerQ/waaXEsmmw00sW6reT2zH8xWbI
S1i/UjgVzpSaDbxNayIu0CabifWylpeHGqIKcAuiYoDIASPdEi57rM0tASghGxJt
xAOwaVk6aCy/bTW9inKOxAJk9aM0iYNlVxNj9D5TiTHAyWviqp/JxJiiYEfuyk5u
DbseWGLv0pQ+eHlvF/FbnlHDMM2vl66hKJYMdzmPJ1/rt+F9D0cabBxo1JZuGlWp
nzMMFDsRg9FQ4kE0IpQDhfVRHIo5Di/D4ylN4SNaUYHu/VncaVYnlHx3Ngq/35E8
0ff5Wmv49Sf6PY3EKL5hnp1KbbKl6g6wxbP/MKwb/9BtAMkp+E5qruzJ1WolhCt8
OLaX9HHaXJFN9zGcMoGbwlalYUBZX9G2dIoVEcx/N0gTbMAtNl7XgDtZmFjtuHCJ
HVR2oY6Pp/N5uyjrv+4MKlUYk3I5zWuLsDtqwzxWzk4kJESlFZMQNMxwuypk3dQk
AmlsZ0YHkc/9S+KQ/3SNNT5kPSwO5OvGS3BlHrF0CGKcmz3Ju0+hSCa6HG1smKbH
q5jYzf69YM3w3mtU/9x+lh5FIYKqLz9m753SEFkIjoQe5fMa0CIiFAh1UN7WJ3Id
RWe3cfZCqWLcFYOsYCBvy+XyTIOhT19lXNNXAn8qbDMarYX9MxzZelZUCJb51Kh1
ZukfWeoJtQceqmnvJGOWULJLBSRj37e8GwXvOjmEmzz67HfplY+41K05heGddUXC
gv1ww3VjrNktzHtlf3CuV5BX3wOg0ZuD3/O5fbZ7tc62R+QKBPqQLxi3Hc13ISyQ
bc5BTPvrAZLm3FEhSBAgcp0h42Ui8lNtWDZDEwCbG2rF85KqXO2hKryrA1jGR5YS
e3lDlauYhhoDGrgCBaPItvR6avuwqFBhsSUk7cHoD5eWdsPmcga+EZaK2lFdv7/j
Dlmm1EsgFaXlWLte9O5edknxnqATlL3GO7HBdGynPfnqCD6b+w94zinOLPDXYLK0
m4TAr5A/pbS8IFmT0gHgJ7jySxiECiN5YhWPgY8+DCEmpsp+UJYEIK92iHd1pSEs
5cS18yjrRvic9WkJ+LU5py6v7FMY9ue7vOzFKLx0i30ERh7jj44GAYNnoNbh6DQa
U23ij0CfytWTUwiT7wLzvwpg8XNYxGzPRRtAXye8oCOZ/VzltfwtdsjTLvxwgnqK
J1Md6br8O5J94pFKsozzXTX2Lyx9A2itSn1over4giwmkuEfrat7IlmBv9d196ZI
Hqx3lZ+LgqeFVYFMGuu1pmuWoJ/mvVGhPmbSuCCJoWyKyHH0AB6/IoWzQz5YpWt7
jMuqVLGhk8deL+Fd+6df+ZjNVnibQ34CRPcaezi+rrgUwEICGTO+BQUYbkWjRZ7U
z6IV6Fbpi+6IeRUQiaozdcZeD1LrG2LnGW89Q+DcuJquwqgN4c0l+MKeKI6S9kJl
Tk98WUM1TN3ah04HWQiAiFFRBB88V9BCWtHF2OYegJnJSRrP62eOnSey0U0+kBS/
R00Kk9T3Pj/Ds4m2Qg3AbAty5I0qEe/96w8+Pi0AemsqKgFwnuvCyqtkJCNi2b64
BxHHvHrH3Y/alvEyJtgEfFOfvv3e8XEcoLUZ4XMzLpwjh1v1NeYwwiMpGCRU5ke3
rOYBUqROignpxxB+L8kEAr6JwUkQoOJpgPiLLLcz3KL1PBZTdCP4PydK69HOFBO5
y3MLk7Qs6ErcfaRbymBWYxmXThiniWGXcoAH8UsWy208jBasGlWOk3jKEx/VoFvd
44qQfNCs9snpEuw3H4MtOEF03L6KgIXfPcvLC6l4dbKSC5PoQwssDhpHh0Xy471i
FEEz+bEhiCpGEk6QNkfP506oLcEeit/nSgn86n1cxF5+3/PihBo6bn9FxU2CQoTi
Orj0IWjapeqGsIEJX+X0CTmSlvroaKrQCLesFcx4PaE3AinZO68zERTgHleATWKr
n6aYyfVUio10zEJqMcempx69hAZ2Gz1JfFaSOMqHukJNzEFqLxRpFQx5pAbSqioV
0BCcFGYHYweKXa1QCDYV1e7ioXG+S5kksHwpfoTAIQW3dlqVZdmuNUk0fRU0MM0F
Zeyksj/epDdZGzlyp3q/kCjDclTKxtDXrjfmMt6RYtd+AuGFHL3p/8g598f6suC5
dpGn+2AnudyiqGCla2WVI0T2i+Rcs/YBipjEiCfqLM2nouB2AtN6ilHgduI56paN
Sadv8SrMTyRFGuNS6xYkB1D/RU4yr11NQpSkAhQhUzzXxPtmrKQ8wEZoXdGEWRn0
ThiGKk7DEXAkNe6uDesNoJ0mv8M4oEyWtvan4bP+vJmLPKpNuj5zNROPBf5uuvLX
P8kw4O1NfoJ9Gx1ECpdeUHHHV/CsgWDzBn8v3dM/5JnEEEKiAEp0GGs1ot811j8s
HNNKx0OBML+t6o6UpHF0KMBSYUKqhDFodI7ZEyvGDf16lvx7qGsVMi3Vb6PfVOiA
hTVGAoJTfGNfJhXhN00To+W4oPQRw1/hwvm8ad+EA7dVt1G68YH8j6LqfIjqj4Bq
eMLVKSegzOcoUl4dKK37T9ipeH/IgLIBMPaTkM0Tvrs6tA1MPms812L2Yj0ooABk
SgbGUXBe5r+3x/sWgitfCbs/FAwcu9mLmN4CUzjqc7QMx5+TZJMKLBUHkB0flrmP
C2b0jrvhKzOMbDnbWCd6wdWL6GcekKDogJTVGVXJRQ9oH7nR9Obi+i1mVYmjS9Ap
pnvtD+rX8OZZGMNY82UUmcEAY7zOWr4WGqgBURJTp/HWIlf1j9eKSnJfwEH4IPYQ
qmZCMGhMJAm9EhmJtdiPMCkW7BWlUE4EZ1FN6oXWNNm+OCEr7OdI+aimgIR64Cu4
hbslZ7gczQfgP6ma8s7Wubsn4m/j8znChlTXHyKUBqXEnY78vrw+liVdp7BYf4dn
OMvgVGntLndlF8xtAh4b+5fhlmRa3RsYn+dyQrJgowGxfNpL7/muADymX2vQc7Xs
ck1ZW0ubEervE2NQuMv74zQ2HSq/ecuEi6XcS3z2I+05ieZcbJkm8GBWaYw/EiLV
r2mtCIjlUkHeJYEFzio9e8eFqD2zTs0boOk3rr8y0B7OMpmZuMJ2eeFBETjqFgWn
y1xo4Ju0sO5ux7rJpYho5in97nNMUZMYk4VDsz9MxhA15tsi4XbV5l6PE6CkXPYT
DN2TAxkEuQxL4QT0FvBBb1soD/iDwiS+HfADEzXJuefEbpo+Y/ETdggDpcKLVD5o
V8y8hcgL+ifX5Cvv1tJEgGubKPxIwQD1rPxAUokJ7nEn4aPymM5bIfjIgmy0fRHd
0iHnAJJ1Puwjry4CaOtmu+T4bja9kliEadXK2bAOD//EUD1N7JnjbjiWpCDHOD1P
nq1Fjd+Mmb4p8T5epT1uLz62i1bhyTMrNw9hYSWqXYl5/obxVB3u1WwSNkWWYphs
LqtstzS+ZC3dWHqbuOyd4+bdsuW2f/zXCi7K6Nf/fldOU4zUshWN3RTuh8XmBvPy
HbTfv4nFOm0bE3E351BmoHk0dm2RlM0h3GdXEutEkt+8Nb3fwVImlSLYpRV9ghcz
Vr69ntn9ihOQFexVoq8MeNjAMUarv86r88WsAaCWfTMNRNxEIxnoe+pKearTiQPT
j/wtwvAeMeXzc8/M/tkXm7o3fxdyQ19/m8vygFR44EQL6vb8fzSJXzw/yDhnShXL
wXybTi30+GnRiszPQxiZEixkwh6sR5Ee+nn8RGNX9dTSCQ5tQ1gHJIGwBngov/5c
gfo9ohPVeu6WHRb4KbkQeihqBEqR2zo41h2Z97w2CAthk64Yn0vw5KhW+KlEHrnS
W+u9GKECJ5UPK+HOk1yEFsKfQYo87N6c8NNfUDMGfvpwRM9UqbcT639Kibjkalgb
RKZZDhrxIG8Jg3kBE+q421NayQ7IdrNx0BdbX4SLEeYw4S6wEeP4FBvjdcq7z6Fe
+X2QQ/GcPCnvTDzMWHpruG7Z39FfOIL2zImqOLkQKTrb1M43rngLYUx2AFM4RcIu
itGqrwzgsiifuWbEdQg7qDBFFJkX/dNkaxl3IXBXkcn4lnV/53joYga024Ddn8ga
p/S5V4g1yKWUlkbD0K2nPQ9xqyrx74W3fDJ1wI5pG2DlDOssVEQUq/J7S6ZytzjE
aYR8f8bEEyMQk7NQ5wGmgSEXFsWS4L+qF4S6XhITPcO0R+2UWdoo/gk1MOb1OT3P
Q9cdSQTS7wnhJHRxYYEp6WgmrW4RWu6dOIaQ7Fo26ZeJr4zFqQUD/GmXcVHZ+huI
vVmL4upgYzxvTTouff4FvOdCV6485kInq0YYgTo+yiBvnBZ4r8+YGenVKugVh2q4
wdzw8Jtewvspmi+dUWIjUvtjXvmc7EkUeVO0VM8Dd3tCI/sKkpFVQ5H4OsEi4GAb
OPNBjYR59FMB9Lw8FeVtZeYoMqgGlPETS/c8MMbtZ/QQCW/VH5Zduo3E9rdPGYy4
7ip+8imXQyqXV0hzk2a8hjcHB/x2spqEDs+uhflu9Dc/4SRvLRuCL86m1jPhstF/
ISkaIeYhrbivoCqTjpHjcOisU7WVJNjTzVi4CnITJhI7fX3P2UXoxVoRTFiUBtdQ
CSYrqEUQ3tGIWoTw0I34E5iZbQKVVThqOaN6gAqDHoURUd6gycEYV0wqW9kwPohm
F7voTtV0QO4sQf3JlLcbgohFFxJGvEN+6JlSimy0I++nEen0x/umHA84smUmbJWN
o5JbensLtol2DPoON1eG1n61ZE+FmjZZzw3YL0Hrs5DsTgLcK9AJvfJsNw/Ss9d7
PwZeo9k/ARlwnfSiIsPFLKaDS+tosSPdjzDddf5f0xO6DqIg8FS5AZz/pZTf6RCd
bY4LeCX9k6l4WqZHZNVAAztTL+riMLkpJXmIFUwMiHx6gZGOgwqcZf94z3OJD2K/
x5AikQsWUuV71Z3OG8B/aTCQJPQJovQFl7erftOzFKL4dh7W/TRR1sp+7AKYGPMQ
hYimW8iB1vSPhnLwkN3zhK6y+QMcUXW6bi7Y32aEw0VCcm9yXEG5jpwj1couRmCw
K1febEv+rud+dBlhIUYUR3ZJ/ybAJEFzGDLfuyWSUYaO9VjAGr9bSRaWkdGJghV8
dtSu/DE4R86gLXTDxa92/v5kWC2hy7wlD5J1a6x7UBV1NCG0RyafFY9PU9sRCwnA
HSM+Y87K+Fd87Dq/9qR7bJ/0922mogUpvlah9pRU/1UQOjx+2wf+GFqtWVqU0BQJ
4VT8vOlWdevWEjBOtXDVBYOmUv7sREyk0L9rN70EtoNQnTvBoqB0meFH+j8+u97n
rWBln0MEjg9Q8umdsZBmH5LuNhx6iHmYl5cPmgwu2tnwzK7ve5OceoaL0fTjskEf
XuaUiIv7wzmWyj49Dh/jPO4CJaRFSYot/7sbD21Ik8sNRpygi9Uaji5aIeUlX/8w
7+sIg7fTymJBZaTuOZIkc6sXaY5gICM7lui+e01wrJmQ87y0xeaFA+I55ppdrLYT
SCEQCCYT/lFcYbMU4OdhHxUO9DzPawRzU/092rHzhwOXLbodn4vM8pKVPArR2RoM
xRbZt/KIAE1T3BO+pTalf8cpgTD2wcTCEJ56yuIbbJzF/Gl7LwrNbBow8oteic1D
2TONf3O3eQZNv3KE0kU8MGKUGLyfw2pL8j0YBPoPW2FL3HSYAmd4mR+1WKRRdjAl
D4kRMzsW5QtU0wtJR4HmbKINsHdNDVHT6tiLAkFcHpKq2zJqBTIT50m1UPC/pmIh
XP/XCrmMyompFAM0rhzSys36ve0saR/xeTU5+vcwxNw64WuFc/DOlo9pSbphCgwo
spRuT9LbdkGCp5+7hpQQ0sHEsR8DfX/C1PMrb3J26SG3KjUfEIy0Bp0VNTaVDguD
3uNaPmPxl0ip78ugl4g0/JqgpHVa0atvXOLcN0HAX2i0La6C7tcHfYPSKoB1J2ou
NaC6tBJ3MYfvEIhBwc7s5vMhMh219KUtvWq10Q3xFPKFqD9J7on2FG9I34ivhsS6
aXfHTTwZZIlPxOsQodoh+/JhvD7kNF5ZU7zzROHEYRVDndrYMqfO35G+/E6ECS2S
fow1bbW1PAEfKVHAz8QcZR5eAy00enBAQOkGirUpVl6yfFTeABMqZuyVjLPvdtVq
EV22tKnRaTuaFveiiRR0FqOpCNrTS3MdZdjMQ3hOcAFAiECKSV/hIHyZHO4cBFBr
M9KUQ6uXf50Sw4Be256BOQVYJdVJs7v98wPB0dj+MfuOZb17xkOcSJqNT24EWzpi
S5POT5waq9+1Zt7pTrKthdDsOiKQ/J2QlhrqmG/b85kNGlircTAR5Iw1fD3CkagT
Oyo3BvxvaWZ5gzdn/c1AagQ5XZoWTe2/6XI78j1d8ZNYcJHzwr4bj/Wi8RvEm8r3
E2kiy9uUtJh8EiY+S3xxEUZraChM9MKx32LeWm+n4L1kSUSw/LP4n+4mNJA+O2ha
8oxdzat8fFLEFMP1HuJNa/YSinXDk9ij+2DMVTiX3V51MtL04Dxn7nF+o+n590nA
+jEH3DAbuV+7GoUEBWsPCG0Z4886R22hxstX/nqE/qsmVlpNGivaFU0ZBcTuwzVV
orisW+eWXnOOjXG7wWts4x+JRBl1DBTn+Tw93x1WJOdJNs4zVbW4Gu5yxqM+z47S
9Ni7+2DK/dqu/t+4/4Reiu67S4NXVNHt7xPqvLdhQlkYPc8oQXiOlhLlxt6O4R1a
V9GiwTDClhTFzqhMOLkrScew8wLi95/i/VCNFo07ucV3Le72fnZK5DNdLtMBrQVh
0HoWbBQwV2jVbAhsvXJHzVN8y/0mxwknm0FupKugUdbLhERChZhsDC6DxBgnve6R
urwqHmZRsiMEWruivrnogqpz6rE2aabu5NjmYhgUUk/KwgvRiJrqu2wOSXTZornC
7pDLwo3gzBu7OImtON6oFz03pztSLah6yDJZhoU87Cli76IbW4uhLLI5gQwPiak9
0FCbluFXQIY9+mkr7c5UXprYVF9kWX8vwvonLA8h4gKdRcwz6vYK5xxnV5rY0FU8
mCUwAgoJhhGXQdVbyQ8K1zPODdmsUsVQzNBoch0f8YGFEidrRyPYohOTmrGvMv4u
sGz+QNFJHVRp6kfCWoOFEJFBdrvu4LZbLwFHnMxK4zzYePwqHPmGh9LA+H7vDa+2
DwzMWyiB+oLcBdpiDmMOh2kKEvuYuhl2a3O2Rf4MnYEh64PdJu6ROXyMotWbJWVZ
6u3d3xvJeag609/FKcN76TwgkgvtGDA82waONugrkM0uCMK+ov7INwLR5YZkZcJ7
z/VZ+KqInC3u/VDwM+oZE2iYYpI6raJGAg4BLhXD8ZQ+97RcV1FacvlR0W21Vp7a
dYWIhXu9CnM6yUGcoNAfL8NilVsgkNPXOwM9ZAvFUysq6idtMKkYWxYkj2dCW/ae
HsTX27xvpYEKl5khs64HQ1J8awdF2qEX3s5mrFnTplWNjOTEpHIzSoox5TMkiytY
/MwA34L0JXbE5q+h+O/Kzjlaiir7lhsFf3aL5E/PtnccU3AS/1oav/RsvFgeaSBW
Xt8EGOdfBULdY7PIuPRCPVD6K5pDR0TWYQ2n9a32ArmckZ7cRkgrs36obxzYKOii
nQqvOmt51YLP7l22kbw/WXiNznLInhmOSBXcG0nA81L+Kf2k7k4hTHpcttxrniQ7
yFahsfd7G9nUGBx/4a63TqLsCGxL+IRr6Dg9Txf8M0SGgKUVzcFe7vpZ6vORcOUN
ZX5oK31eV8zgBrMWpHqv8mu4qsB2tDe0qvls4IHGfwR4nkr38EksnxZhwyGncJNP
8hXQfiZNLLpbVyLDIaBeR0LkH7BTuPw9HNnw4FEw09ybNNvEl3dsGuVkw7ZGExrt
TAmex7jqcb2PhL4QDTvndlRUyJ1XujILn3XscKSVAzQXcsc7hL6mY9a4ZIcaAmvf
JkFcJDkSHRtHlfQhndsUvJftBjaLYU24zi7bFEPvN2Dha0tpJJGv5poWx1WGNK2x
qR8fDk0goR9ibzlspVH4ogg0gxxjPr1M3ul/DSZOwrp9A23yYUYSns1HATQjQRJ/
UZhvhjSNqrOVcqtsomHtodbn+PwVXMi4JQxjuPVdxPXQ5atcsXnRODPFPJann6Cq
Wkuy6X1y6+3VcjW8FiRyiG9GxwRAJ7/iDf45+BX51xeqn1TnT6ft8xBDed3SoA4t
fdL2OXADysDJsDUpJrWLNJkyNYkkpO6qlXa05og4FBEszsvs6GiuenLY27eK/ey/
vtbE2j/teI8+9u+Y+VV1PO7q6JN4PCjqUHYI0z4LQjWfbkys113sER9zTkLFg6c1
kSo188QzHRCwB9Ru/ASjN9CT5p/SajTcQvFi8N+9E+PL2LvhiNiG3kcDEN5lmqa+
VWxspgg4IgJ7Wkw26CaTSvGNzof1G6CvberwtB4Ys2+I4wWR7RPwHMNMNVbW+P/k
R4zwhGSfAKafGoqrfHinPtudHmH0w0gewauMi8Ksx5hCqBftgXLLsqYWhuWx/u9g
LI2Q/y1kl0L30Z5HFe5XtxRmt2hn1r5DmodtSWbKJJgxcQaTqOW0qlD0NYj0CHgN
vWVlkm20n6osWM7D2csFnDYevkagrFHmGA9cQL2xGQmuRY1qzVRbDTRpMaQQBFSU
28N2HMFqSB4P1BTAugigPtynW1f13wrK/HzNQE65XFtR7lI8/SYJ6jVZPNRfaw48
EOT3mHIoQJBGq/usfZnX9v0Nm73GeWR8tjL/7BWatzVGl68Y3YgBPErnJ0XE+E3T
/M8RFV/FvVBi2PHa1FUeFAQ57SWUi+xZBYPLZeyd+mLxvF2vullL+mTgzvPgzFvS
5X1ZW9TJhokT2A1GmP6KFgkXHaZnSQgcFa46VhQwxmiUT4qDUpL9azf+XjAc0wX3
vqlbLDsnF5x1vtpT1v3cA83rxQhAZ11AH4xh7Mz1D87J2ort6O+BhpWV9Njo7x0f
L+lQLSPR02CQ8CrEtLOooXH/A8uMesZmQLWZHsMORot5vQxhd5DKsLlZZlSK6vgO
Nt8zNAJAgvIys7Pg+xyxaAAJleh1mi3uNc1UT4wgOJ3zafpDBOpHHAryWykBnWu6
8+MbuKTif67lzJiE9c6Wf1U3btSyE4jUU5uFaje8MnzSjT0QSb9sdzKSdaiECbex
xx78s9lfEe/+Qgg24bF3KAStJ1NpgXcI/3lM1emERUQTRGdgf6Vs4xYvNlJ3umhv
v9AbHexy4KqH63V4XYDYxlzPUA0DQ96H5yD83rhKmnfi+GYeF1PcathCNoK9x0AO
PjM5urYA1krrBRjg5mQkDwwT8fUvbTme9dUqFVDqdTf8OdbwcHXPwVu/hGVkLXkZ
1oFcD9pr6LE9tXr5/xKO0IyguuJ5EklRYqRdJEK8ZRepNeE4LxW3EaMqCuPk8RRx
dteOcJOhNklD96CQN7jpdgHtz7F3n4Rqra5WhnlvROluZytU61Dp2ymh/28t8Zjh
fPJtLkQmNgrhhQL8FzAobkPQHsMA3VsWzDvpN2tVGncASH5Uk7bOAYhK38/DFFJU
KdRLHmqhK63EE2vZDBj36LvC+0p08LGAk6y1GL8HD/k1lM6UNjNZetLCsbsY8eyP
3hQ/pUa0FP7PQutjFVIIY8MHkuMZzQ3mnLJbE3fWhskN51P72UpEqi8lIdpGN18P
6eXsskiRQXQ7kWyawi9Pres2drG6sU03rZbPJXYzMv+Hj2SBLIpFkxMnpoLpBi4g
oc1V9S7xaVlG0DYojyiyz+WJyHjGTxtOBV6Pl7yOUiIYgy1r9xa14fDeFHyD6o+T
yFNqlQsmM6YNxl5QqzVfngmSo60nOfWknR+/glU9xAJ7X1hMPPe2SAub+MQCwGil
3Y3Lp0WQ5LOh0UW6LdLNb6GXUziqPHKK5COZ2z+QHc3BQne/7BV4z5/1g39hDLSr
QCrqZp5QvqqFl3zF2lLpdCfWgjlhjndio70k7p1y0bU4EIuK8JlpvcfonT5wWSz9
NixofeSypRvEsl4Wpz47eqFIZ+YaVvS01t+RBn6YFJsEYKA3QhiFWTalPNO3nOt/
Hw48sfsEf3EE5mltj/ZI3gG6ZKaBpqmzp5Lr+78ILnpBMY5vF+3qfKOBtNvyHRVc
cQKGcbpeL6zUoVaKfK9ogbffTJ99zAFbtaZblmw+2mCGKcD9vMHdzfYeOVqEqukd
ENS7YO77/P2kPqYg7b6UZGuC61d+p+Wzam/QUXqC//muHp0Iq3iUJ01F1psW6FcV
e/9plLu7z2RGwK9FNiVc2jmAMUhS8pSsEHiHNc7n9P5qXTShyDeZFhrd/CwxkZ49
+eiLq1Xg7bJN237OihxMYZLdk37cL3w/jp4jCb/oyzvrNHRvzKnP74SbOb1QDpYj
+iZ8z16Y1UueXIofrB+aaxhv3H9tS+4ysRvUpXWtXbHG6m9rkN4orhm1R/Q9MXv1
lZTn1YGDS1kirDOLH6JaY2eoimWGrLH0G8aTOgD8e09E/myR7JuIadLiZQqC/rHw
RDNYecdgaFUFkLujPAnAYkf9weJZbjsBqa99oajfi+DPrGTx35luN2tQVx0z/wHi
DUgLq649Ee02EmGteW3KWnHmX2XH6UT8kqYQ4MNe31veAj5UWCAaHxrRbiWKXlbW
XpjGgIguxmKucOxXPmq591iyHe9XX3pmSyConHMO5xfIMybd++zYBsfbgo/+zlTu
DuAQp1DTGX6puSwL9Fi+VlJ/zTXcKV1gW7tws28de1zghatS7r3M5iQV9nOeQJA1
Axdg+A3Y+ugSxbOClHMd15T9s6QnXfL4oJqf1vWfpgPFEN0YmlyRD9fOagWVD+sf
uwNPVbsBW2KYgKEVy59be5RdcscLaIEj6pLjuNzeD37EMq+RUWGNxDqe+IdnQDW2
vtdby9z68XIYE6rlCM7vKwqwv+fduxtQ7yFvYfgJh9Mmv8wEBuPayH9sJpb2Wahe
WPtk+c/kCHFuIekIV3WRyeu/tC1QcmiM6nduLmGRls/93sL053J50tJk3UXU0uiF
BTaOIPNItwh5TQMO2R3JJNwMewt+lLT0NhQovrZZu/Mbb+gEtQgulSMz+oF4PZ9u
mjvo5wZMnQwSl8TEU+Xt9tqffCLKZ6W9GYF+V2hI78ATo+FZP/1Xj7HG5iRdJJ4T
aM5reBEd39TYr1ww5hulHlJSp0J51iQXwpG/9F2AGXi1QPDY4mXsXYOuKSmrlrGS
IzaA7VOMfHibV7FKls26U1g2eS859d3LCfGRrMPZfyiwhNX/3yOmO5B9rWD8wM5l
fLE8G2WpWegSWbhu4ZMyIcR6/MlDFJzu7FbG+3+EQfpinfY8FlpEEuwru3wz7aft
PHBGfiPp1fPK5PrBzS2j0FwkIaQZ8pS16Y8DrZN2AkUst09Z5NIShW9rjIkhOewl
U+RniOOFuQLM4aXviQuSX6irNNv8N0JWjd9ZWizVMklZDxsM4lsAuTrQ68exL4JP
RZSeFY5++7FgIM3xmRkEM//0i7pAm2VZT+NV5577uZJo//joJlm/hHwCSRzaD16A
NR3daGP2z9I6xgGA+Ipj8dIhc9wQLczFl/BCoHprWkRh5LQvEYufV0XQqE9BZ86D
Z25T80dGsYgRXZSe65ffZ+4GtmYu+vPPu3NPShmXboLZ9jCq7QhK/3fT3jNtGA1/
O1Od+WPeReDZL9DMNGb/9/c8uTSjTIok5sLvykkhGFmCpQfOkHPIi3qaKUu78pbE
uUqsbGWQ4Bz/ktUC7ByvNFy3e0GGkTlnnIoYrqDt8hEDtJbbKBjz/eZQ+uRBj9IO
03zesrI9rL3Mm8Gl3TLl5iikxrCqVFtjWuIJqi4RZfLi7e0pxIfkbCDQGbOF/2/K
bbh3/bGaZZ4JYf9nUUaRTGgslHl6AWA51Ce4P1oBPvYok+a/TRZBoAACsZjhQLI7
6zi54FZX5ZiZjarIDgn9LHC8EGyfJVHZrTdSfg6H9rwEehqnBqflFB9wUf4GdQ7K
gScBDsZjy+TQXjJcu0kO55J8M9axVBb/LdYrt3SjE3obJ1CuKwvE70x6M6mL2chu
8Ivmwrq0nSR4teHvZUICCTCs27yJJqIZTzplKnb2C8X12AV88EBFcsyNN7TLVlOB
8QLlXB0m15QfRGTJ7Wqu8TxS6n/c6Fb04TZQCAIIxygi2B8mlk4dqjfmZAnI6GQl
F21BNBgaVqkCk+hgBWvNfKwirpNVXXHMgwfGI4ef0R85F8l1m2hYQlan5C65yTJc
Q+igzCE8L8+zbBz9oW8AK6piB5z/K74zFC7Zs+yl6x8X9eHsHcZQBIJQD0drkyJK
625zmtRL6s3KG2ovaY8IA2u9ElAK6GHk3p2Pt3VIlpiRyYDwmdW4+nxEP8dhRo46
lnVd4Zgz74IQtBgy/7pX0sq9U6mSX9Ywpt7sFKP7t/FSE8Sud1XzyOMZ5/P3ZPz9
7QZM/oXuRFYM6RL6jYWlVcaA+FD9fm8bytMn2ehYKsneV8a77O8iMqwerc7pECPI
n1Vc57Hg9i8n2vFwbOtK0HgeILN7YD8v/q3cV8tMcWtT0NQnzGkZrgXwoPXkTIfG
M0o5DR9YgWrmB2ZrDArPwHFbpndUpt0LmCU/E2f2JhqsxGK4qlVCXuqubNoUmZV2
lgihGoaQTqkwjXIGEOdenUvGiUYzd39xGkhGJtyl1F/K9oo0DZvdyJ62mW4Qo1ly
ajUEDk+ERhe2Oj2eKYaa4t19JsBiFR9dpQoCVupBJqwk4ikN0nWeKXUKYGTgnV1H
sX2y1inoJakx6ZU8P06pb5hWS+Zu+Cf/R97NSRyPQ8Ep56MG21BbivcVzM1HU3gN
6n60cOdK6hUrylGTXuEq63AidxbyugbALPgAPgujkJOYGKocXH5TiOKdC21o3X7F
IYODTFUEA88/w6LaULQBUSy8BUmQI9pVgBIA1RA9jzhQAh8bYmS/K0mL49m2m78q
5V5dlaX1jqh4UzFI+L32fVHcbTi/z+k0w1A6NUL+wtJUYZl8v3ZtPQdL34nHkpkB
bzSTPCzRFFhAyw9aA23KY/Ve1LKx9VvI0bWw1XEcnEzNyCckFRAE4PpGa7L70zFe
QZ+AKsgLpCLK9enaaxkB7NjeCelO//WPs9lGJ1cyP9ViEdN3zebLbcp5lLxaf9oS
aArGWnlJhJ3+y3xbBV8/MutzLd17LOYCW0oKB4zDDHxauNWUBBvjgHyxXQPuLHfO
fitl4s6qaAEcsMhM3zToZVJmERASfvO8k7x4ujpCUxsJEJf61ienJnP0SRxV4xXt
OpnZ3QtFn3VsAjZBqH7Ns7sMzJ4XRAe6i8W5TUDBIAq1JdtBsI/eX+Yt3Ri5MsVj
32+mf3Dy05F9Jchfn6QoTVWP0bM40e5zTkA8Bkdg1YCYfAQO7Q0p4fvwFthrI/5K
gaaGBWfpB7rsFLcYDh19EUiTgzRu+wlpQBQ1pV5THcqhfB+E7KSB6yryxLk9/75u
aXk6sXPmoZQbIHMdGjxqcIVOCExeLPLT1QMw0YFtvPIiPmh6k6SWfbKwKeYKieug
uLnHAhAg793n7y5Y040kt901uJrxrAJ1UGsM0RWx90bAn0TQ4HHADHTsO9WeH5zS
LTuUlVElicET3kMbC4BCO6+CamQaUtCNlIWGR6T7Ng8ak/FyZnjYWhD4jeS2qDMB
vtz/OagIFEb3taAIipqldVVyUSiFUV9q8MsVKOvvKUnasW24DCbCyDNReoDIy/KJ
Th0zXXRTGdyg1loauobxJmIp+w2jdSP42Nsn6cV9BueY9tODG3h3K7QoF5wn/DFM
ZaKysUzPLqBQhYY0WG26FQnqvy0eZ03tR6j3w5D2lBjatp0LARotw9fPhHUTJQFQ
qmQp2wC+VzTiy+nQuNSDg9n7bQ30Q9uP3SFFUaKTvTRF7p4xC279Vpme90vd0z71
KCFVM73AI+mg06npBvSkRX8tXH6vAJFLJGbCQg7u0LFMyFxrLwr794iuEGMjSz2a
yyXusD46bt8SkV+uPdZeemQB2UxWFEwZaHwUJQ3AF/HAyVcboDH6BCmYX7qvT5Dq
Ibq1t6EEvN724UxDwTapBQ6z+vTl6vrnufzKAgyxKz71MTyUwzt96crX3KIi6z3t
mTbRYhdoEh87PYxQ4Qu6mRkBDS3/CP/Dfa2NiGtNeb7Z1gMpTOnZ01txLCx/QQA8
zjyQCPJROs0yEUfMyyHXxhK1UWtcboC2jffPmpHagLUNgWGyypTv+20iyojDayln
j5pbcd+uJB1GzagFksuFhLoW6jquq8DJoWnsmEcW+X991+fM97VIHjDavI0hJpZc
fP4+bMjrpD9dYgnKRvhlbV6c2iMIj8BZlss2U5QblXBDl4M0aU8QVUp90ZMqYTgZ
b24Ph+38YkPFNuGKBAhTxqo51uvgX3JkumpHt9WwDywZdZd2T7DnnTdTtwyqLPYq
dEwBiZiGwWE1t0oQp7W8SJKLSg0SZlAq3AqqoGgtRHDevIRHHB7otKuZXNU8jkHy
63V6WY0Ki/nM9IrUy1yjD5lWdYgl1xoD8Mx7lPFV5ICR+0evwcbf8Y7ftp+zaYR0
hcZkK6KDzxbnH6U3YNW5Z4TTEOZ1G1l+5UOcTLFjZtRSh2qTsy7zyIkzPCFVkJfb
ZKpigdRSzYJPU+GrQGBEMuCFTPJyVlnF6sXRsFtC1na9lJ0zRiyDg10Ywrydugav
gLR3Q1ZYmgmq0TQ8znKe/NVrmSmkooWuBNhX+EOZpp81etQKD5u5rfpUlxSi5HN8
dbvKiV8gKauOa6JLSbKIbpL5C9I9pu1WIv1v5B/Evw96GnDJLQH3E6ewsSw0eZ5R
9wfxekvzTHkrWwYUPo0RoJx/v8dPwSBMolSk90cgw8DRUjqjKPavjjcR7kMFsdeY
mCyC3Ud9Te8sB2Pw9Tv87jOYc9MaY/YOCQpbV2FCAb0dJPy0dBFMcA+nrZgC6MhB
zY6TW/72Yvay5xY879aELZPCdWcFvjJHu51wSGhhurRSCsLJrLK8X9KUPNN+bYqA
LI5zIiCzzX4APfT7z37FauKIPtMc9JJW7jIyiZdq/Lc9oaGhTF5yhbmSo6xm2J6B
Gnj4yLNmcR6yNjCDkzpj6fBEW2aX0DCA2+6G+o6SNqjpujBTRnKkFdFAfi5gBkvf
0etcQ7HRRrJrlJtFUZ5I3w+xnR0Adc+CfhLlaSE+Y6FHVvy8j0c5qPjZ4DpTZJ8K
QIwxQKFhjiy9EjKBljunV96u8UiEUCD6EEG8miexkIt43JyACghszIL7EhkWXoPX
LgTYLSz9z2OrlGcs2HVIYjCZ5uEc/xGDyBditqZ7uCNdaKGKv/JJ8Tr3bfOG0fF4
M47ySIVszN1vmsJlAgpKgWxk32x34tPcX/1W1/x1UtH9R0KNUOk0ad3jBlUO0noz
OX7GHaWeP5PjuzlnoPQa6UvdMQ2Cm/eprgrMMM/g+n87rW3CfcxIHI1xPgn+2n7h
lIIoBBQKgqO2wNQozpOdtiMsCYI6Bbkjehjj6GnpmYCH1ubCH4E5SceAfeHYKp/6
HsazdlAdU7r2Wt6MXQIcGuYp+tSGqESIRUzS/Vb0U3sPX3o4TfcRMGMAjAb94mAA
AbNassrzGMWtV1vUHrq8srD5evC4gSs0PAWtoEVBLNsWQmKEXgYvLwHlurxRwcbS
KCKiTSC+JPhpgBaXoLXQTjn5eW57QIcJJxFr4NUwTkVIRoiOPVRdLp1rcJYt3E+3
bPC1iEU7qKbaw/gILsHc2uQBeSWJ8Y6O3joYbdA9wBpgaRrHChgIqJjKIh94pj8i
tgNV5B1iIJcFC4SKyLQkZWuGGoJgmqVEaZcUbmg/HfRdyWHTTgBIWVCUfHvEIcDp
/f737TfQ+403D4JTtH/H9GJDdfmeTrNu0au30fjEHRWfyJPKlh8K0CQUq6LitBZu
sTIkYHGGuRgoU4LED7rVmrvt9XuViYj7Ma/qs6MSSrw4eImV1qvLSy8WUa24Bp2J
DyxiLncPjAWPXohYqqUc2bq3SDsFRN6QFFieIbB8QZi4we5GUa72b1sqseEBtUr6
UPzffAhQYDLTPXIBiZx7CAdcES1VRIcbJlKEyxfsZZVSzbLSgmL5yJm+1a8usMbz
zbt1NlolS6FaTA4ytuU1KEVcLd3m/8FKYojE3+7khBwjZ8bwatuq2TiEypoHnWiJ
Jehvg3ZNgYKDIV14nK6UJbfB/hDuqa2ZergCTXf2PWz4pXLo/sSp2jwfJFDxPJ5v
UDT2sSoTqCzS9nUHkTR3aBfPKOovHe7c1GBLXNiERJ/zJHl4hFUmUETKDXdcM8j+
KYiZM+2XHD4fZGcEqSU5krsQ1Yot0n6UCGJciGvrDX/IbCWJ70NvI5MltoDC8HFY
UhxYLHGUHpw3c9zm2QQK/g1pR1DJjMb7BtxnbKZwM3l5RAARIsS6rtsD99Mr0man
Ekc7lgTS6kdMmqqxznKOdIQEZiSulq3Tx0ESo704M5AxGkd0guQcbfL050bWuXVy
0sjyWZ2HN9Nqcb3uj90+tAFbo7iLhh9yDJB68oKyQ8Li3AzTEN2nOoLXJ9VB0H4+
yrjiFOX9Tj9y+eIreIsJ7KMlYXl1VgaTI2uYQKzWuGEQrPvqdZIPTh3nsyyhAQ0+
CYUWX1NcLggthuQFj2QOUXnq8hSlx8ffBczKTkvEfAWaCTvG9xfm5ZPoOoPz/ZuA
HKLlNKJCS1kWdwIWw5j00+dFGZWQqywVCJOsot9+4bz+3IR8g+3Ow6RGVht/FAIv
TmyclhQ/GWqm6BvJxXUEZMQ9w7rYBe6FT2+9gYrB4sv3UBkXQpdtn/uc8Ql8XO8d
OLlFN+QU7rllYrLgCfHZIt/2MDEne2kkUd9GxP62FdVxHoYxumoXHo5I0U8HNE8C
KRWzP0Dq3Ga9w7o+5oOe0t2gUeMpQ1XOaOOI8Qo8TGQNyoCXiBaW90Jx3nNiC3Mv
5rRJ9X1ruHvqi4aEWM2m4tqaSKNSQi+GIX9nKECHIlfLpKrzLlS37V54kW4/QlNh
fP8aNV+KczOgZHlVCWrRYZBAdUaVCFMF+KjdaX+JVkHtSveMcNL1AqO6Vehuhec7
rzeYsxXH/pFA5dzNM8GdFDuVHU1y0oj94Q+OJ8Th3PwQzwIp64p0XFz8wxhR2Yj0
kn9h1sk8eFC5RV/wSrF5tpKGfeRIONnEiH6DSfFzCLdcqoQYIxaFXk7RzGcEOhw6
8TJFklChpHzoJZRlI9Thq0s/pCGX+glFbSMFgzdBEDpj4tyBI60PC+MZE3Lrv9KB
FW67wSayvPvJMwNw5kEY9vEtLkJ2YIErOWUw+JqLWppCPI3wRayjx8ATbby3zG2h
4i3R+2dyzKTW2SVTXGx94Gzdd+SLyKYDxi+/3MBqepkNmrpDOL4904wR2vJrp8M9
Nu9Fomc8K/zvn64ptSxCI14WLUEBYIzBZbkkcz5OvHKjmMs8GA2QovTU6uy7aRfD
SOe/xFPpqB+gbOn51GiKbda2cWwQ3VigQ/WaJYeKQ/Jrpbes+CWCnpJescaCe+2m
Ek+RNd9OA0Edp0QwAJX6WkjWnjsmRbZCE97m1AOhMPYRt5tWXY1+/0kbIy+hHyoG
Kjkyyb25Hhnr69+5ziop+Kw17S6GtUklhY949Zr7gLn8x/uXH+kG8FKWXBJcoDlG
i0dX9uTD0pljUeBjmOKsHobTwduSlKsSFdxZiLHwNlj+noEPMT3OyP2HmaoBvJpb
fL/WrDnvwb4LwVceiIdQAubK5HqD8FcdreQNkgZx5goGWD+j9cWp1oS+aW6Hs4QU
L4uNFpOPV7TWjD89mJGBufS080l8orRiqmuMIB2ejz6Rpk+LydTefeTHV8NiYMwv
TfsoeeuuEcyZgIe26oKUNbzOO4p9/joDXs0wSeog9fYxGpz/WodYQDRbM8doqiWm
8qYkiEVB3eJ3g7oihqd0NylqyHLuS+ZFwfU8SC0yfBdfFmukGrRtmr71pT5/FPTj
hwwk/Q+4zfmVpFVpH0VgXKfXY++TlflJKNjTkbachfIyqCMZhw5XoK4NPuyW59U+
J9sVxy2RIAUXi2Bc7ezoWCBFLzR3aixhr31+oNJORI8KZdxNYlw/EyxPaN9ywPUU
ZNGeEUq3GlcFsf4IZOxeA+gwwZxCInP5AuXifxpiWka+qlie4To2AtMtBGPikrCx
HwL0sv08Qx9zG5Tevgli2qfGv60KNrmbTOKObAt8pgBJx/yBwrXvturyavFATSi7
K6vW38X5tCcWj12NDBNjTgnIZXAth5D6xk+fHZzj8oWLLXGsM5NUKSVr5UHyN/pe
ol7yeW6sYUp9aOnusRZamZqjbL7pmlr4pvKEvd+DOXuPAV0UwzCRonq+DW+nvjVM
vUz3zwbpFVZIDCACzl61Hf5tQINEh17IsQoD/kkosykqO+VwT3rtftKnrYvj7ROS
XQuQTTxqn/Mx4AXmYYHKCe/WXQho7Mkj01h1tQrTwXiRPXiyjZQKJ3b7B/G+0fjY
57VpGo/snyI+8AzC89CdfDrPb4ML8uPfiBxEcy8spRUucAB0raR3+9+3GLRzDm3B
Ois3Jvtknhp6XM0K05UM7xi3RBxtVO4NURZz8whl7Tfp8JmU84mbOZwyog8lVq3Y
W8tlRvYW+bheZIespuRIMQmHffbyrHVBWegt7Foul4uPlRnJV++QWdXuUK2rlQBB
yz3cLF4MWYU9ltu+qGI71XlF85FfA/uHDNS/b4GLxjy08uey3iEO2L0wjhrvoUsc
frOchojuhSByCLapo3sfiWL/0TXpDKIyUpI19jbAYTMnWk/AYch+aBrQoUIDkTkN
IyJVe1Sy/oOQ4P8WGVqVFdhFvzwzXIegUPcFcaYNMVKF/I7AwarkXjqGI+l9JR+i
Eum1I93igtRBG+qTgijX7CDUBFKqAvDpekN1rFoLskP3SdaNnEFY7A0XDpyNgMET
FQexUiiYA+CnRh2QhVJZrPBbJc0tF+GwuJls5jXezxI0oKBF32wq8+NEKCFkj6Ur
rnBtxIPRE+w0nolr7+lsfi9SppqOgrUoOuU9X3R+drzNe9+TreXav9BbGnNye8nd
s4Y2oYEDl5zjT4H9x6jvZetLVjeWIggrJB0aDc3zO+Lx6lNMAeUqNrZXRBKdVU1b
6uO5WNe/ru9QdwmtWSdKXP5t9ofd7fylMLtnfpqC6v4xuBZBBH/9617VWaJSjKXO
+KJvD9uFJHtgHjtGOavXGDVt9Cmq94hu96/OT8LSDJBi9kTBSYBfeMr7IcVFi7tt
0+/01osGxOtiS5EsRAIWz2V15qRF1o/X2Bg3pY+3JhdBPfgp3V5enhVrQxnf4Goy
KoqQx6xBQDjw5cPp6zckzNVAHpbgxox3RN4DA0SHizfwkQhBzniu2m3tE4Shy+Vv
avgBOuaxflIhVmRRFieLpS/IA4qH9V5Vbq2OiTUvG6bc5AFCv2r+29XIDs6ib4L+
YVxZTXAMcBnniAZ7iVhrD5A3i26pvcmci/1BURf/8p6Hn33kInAtz2a+UbGnCCYp
J23mrT3/krgpsXdKVhaS0e+Q5Y/xifY/foGcEZDQRrNiMqDJRPPzsWuIj7ExorZ4
+QouzO2xPV6G2mOXndep5Pkq+KyEG8+pwWcQkw13rQReFmW7BVXEvjxq8tTBhBIJ
/61j4xRhXAgXHijUCf+TXUCanDKh7vUoV1egJRhiGKKpb22hgtyE10JerHl7J1of
fDjnkyUyF0BDjQtMza31QHqhYxIdDtMC3r6RxN/fEPzuBs0Z8TC8fnn4CYkJ2GlT
sXfWXkxQQ5Zj6W6COn+fvihyYHCaWuNb37pRvs6tivkFEqcfSSaXBHMqVv4iYsVr
kd6Tm5280akS1RWMCpN6ndSgkx0UPZsulQiCMFM18qzQoBX3cjQTjGCaeNYxoj2t
nAYZ2lxc27blZ3I3Rf14sySTKbv34gr0loxbKzK4LYc7/9AUMuBYg9duVhcIV+oO
HZs4P1qXoUu9NbdsVFC9ieT3pZ7XNY43+1XXP4HbpqjB4E/1tq3OH8U2IAXKWNlI
DiZtek5FSeNyNhAsTRDoPopPSbeCEXuIypitOqi4aDKqMfMPvIuAbXmu/XcY4X9R
pHOhvk3+YeQdPwUJPdk251yXzgg/0XPbx0jDm+MYYgSwl41CI/APvy0GC3dTruWg
l5Fzanaq+KKwEPhpDLYZcF7p8HctDNEqJc8YIvUbl0wp25a+C20uQDUEd/QMJqMi
KfUkJRvnCZWBs1e573R9k5r+YnZfB+LPlrk6MgnhkY+vh/FcmdC0s1P1kFfufLFB
hJGpfvVXHWFgpzUuMpO4ly45crSlV+q+4kvzUOw8nhC/ANwpCOhQQWvAHKUvRMHn
h4jMZLA9Tcx1x9SRMdDiAcjR8NwebKv33Tb17iiSwNvYf03xIDbmYZ3YwiA2HXuW
mP8vw61r40PbTPcvUJQNX5UvHBg/lC740I/JQ00Yj6I1lgF/YjJRFkDsWx+iwq9y
eEZ+7btbK9EOC9oqA7y777KaopOhDiNWknKyq1KLcewV4DhioI8ynx3bwo5JnzUn
AW+KX8NisnmCZ8sW3RBFNUnNlj1PJ0Cb0PrDlo1e2M+SoEb/2Mn/2V4Okswqi4mb
Vk3hYO9IIn1xih1gJkSdCZ0liocYwHqdWeImkV98xtwZpBr5Cvnd9t4mK1dch/zh
+u72xvriFNIAr10hOQZk4jULUhvQuCgFQVGeHBV19wtPbA4WjV5VadKZVNZjwP0u
kaBGbmdHqJY21o+ynR/Vui6WkLZiN5GTEfJM733HrIvk4wPpHbJVVjoKu42pKCXB
/y898XgrOiC8Bjy9RMTso3DnhVN4aCu65Jy1E7bhbuaz/202qXYRReCh1ClphbYn
qZ9nmuWssM9UVIk+QMrxUvUm6ic3FrVPQQ3wBwIYaPH4jD6AVvMJceie+VCUS93w
zkQWG5OOwgJDg859Yfd//0E6mqzT9mhN9Pkf0oK90Nhai4Vw9fZGYtiO/pB1Qpb1
HjKhBhDeD0iXHkvtNQILdJJ7Ys6KclQe8LP4Rgeylqw/apJERhZthhDvWrLTfm76
cvOUlFD7C+flyMs1TEgBKRUZMgN6us4RQXj5Vpc862Sj6mzEhrF24m00YyAFsWjH
1nDcI20H2oVQNfn6yDhcD7z/z0NkqJWzXCir0BHAByfnDLGVQ91wIcxI0AAyyDAy
IgUbqPObteM+TVaPu2xAtFEYWECVrrywofqFnze/SZcSLPxi3QU0t3dQIGBeizfq
VWm0ZcfhwiU+rrt+pw+/DPH5Dw2ODexAel14BS+bfH/cmSDjI8vHCupxJcs0me4y
4lgMhlEHzEdA65ku+pd8FPPq0AtuQYuu5XfvhmvoRD4pdgbm2LdjudQgWCNHPASe
/4O2Vo55vs8W2+oiAzFscXQ3FUirpWn9CF3XJ++XHosZ5gzN8f+0IQpJwbNirBkV
UqJle1D7BSksqGFlPOJX7feGrpHppOaSAoGzae8up+THDqPbaxr3QPy41ag3WmGW
lIeVHwuRRlBwMxrBZ/KNQuTXOhTsY4pmbU8HGjgF0m8TOnYklrIkhxMb59qC7q48
CmeHtPbS0atoP8TlAx5Phsy+X40x0D5QU1pkxrT4t0B9ZZ9PTgsnOdwNl2/LpcgW
kIhbdvaZf4FzI35/nysJRpgp12bM/7O7dNZdKtZHZchB//RR+C9b24hFza57rRm8
QyRYcJbGN2q43y3bqU4VcmdP962GxXw85B7ORS1ieIvlLwDxkFmV5U7UBDlcpyA6
dT5Oad5QmSfK2SAMUok1jA5uGcjxnsQ4uraHEHEiuvMitHqzV+R3m6MWLFyp4UQI
0ziwMK5YN1sch3jsBupiEaZbdjKxSHUg87QHf5GrKJVBmDiLjh1ekLuJrS1DwAHp
8oRDeADiv4h3vPHD39Kn8ja88dOLn052/1/YS6PWSAkJ9J0+SWDcoPHPLbabX8Xn
7k6mST/PP8/dX2Z1ODgWCzsATf/KjAAWKO8OHWRD0oT5FgQ7qSkIdpZVuKry87Rv
tTciYBaebZJqXK53S8Z/7y84N0/7LtC+3SPTR82qsgEbebJ5ci0IUlnCIM+timUN
Chcnyms93kigYK7AZqEow7yCRNiDrAlsMqkUkpPEMqoOWS44gxf9v5lNkWkwY8FO
0i8U32PePy++Yt78IAhjk4tutNYbEsz2lTIktjJM/SZNKER39AzzGL7qrIIvuffd
nu2d495RIg0N8psskDzEvvhbR+jMy3EEwXoP4/h26lxbF11/69RdjxYXqhsUKIGx
OJ0GZMK2sBT8DxEzPyktWOLEf9UCy7WnbVtYjxIYFdzMdvoqCg7jGhg/wiHEGHTg
CU2+os8jE/XCMM8WdRSnQ+kc5uN+cuwrluO4895yMcCKe2LCNOBlQPSgOm/J7Ox2
NSBEqEiELH67WL8TCjw/ckotUQgKjoo6bZV+fE0QJ8UlLDl3el2yCERMI3jA4PDr
N9bcPuMlhXCxGzrw1eCdcl3SzbgtpV6xx7l6/EYSyGMqKgKeP2SHkKhP/OUVukmZ
30+215yfLD8qZy4C13olhKcAniO79Sdb/OKA98VZasGoArK9TWb7uOHqPyvLQ0BS
dpIjBypYux6bvcMBH9IywDOLVNUQG1C01OtD4n0Qp4Tu4m00hK4f4syVEz3mVBE0
boXCOTrYJllD4KZ/QhgLFdXEQoZjMT/7pcxdt5xA2qGkQFf3kfkLa65O6WnGxrGn
Uytaho7jxNgDfUYcwsiWrYr5qAusjvnhLrHGHh5wPEe0JYetxwE7wwsSzWGxrrmu
7grYi4v4nOO2TurXetqta2Toxarpd1I0VyN/h2ETsim/FJHiSN+FtHebq4oeMQNt
TBUWogXCxfyATntQXpBashyB0CsrAcp7b06i5xftZUlmwCgCC7avuQ4nFNNFgetv
k7m3y5kESCspV1nS9narbT2mVcgg3440y3tpktHwaMGnZGNAO25kC0rdtT2JWz9D
y99fxU1Gq8NzvQzkGbDu/0Ke5di5o/6oNPyJjyHJ/cbRaS8rF1fnsUaEALm9qOgI
IhjhWT7KSfgo7iB+CPkNIalKe3/YRFmteo3J8Mfo7m0u3NRqOjrwxwBSyZsx7yU+
Vn2Bwk9xpMsm/wk1A546NQ8axn/q0OBy6IXaxBjvZ9Hi3OhYgmeBPBnQOXXnVHnW
Tr2GkG+TXAYHrEA+W5+hXAYMJyt2GiAzI8foRozuBq4bjk9or0k6+wR9wU673mlE
8mzmASdvnolE828CxM1ikLSDOSSWXaEpBDsWQEpMulntqOtbZfZrImCPInkaAKtd
K2MQM9U9K+Yotq++dtpjvg3DjC5LjpLAVUgkxBMNv872WiV+ieJZuXcxCatEVIMN
YL4o7H7954mcG4tDExTdbg4S07nNhuohZ3qyc1sIvMrlK8H5FhM04i0zhCOq5wIx
b433AVa/7o20DfA9L+g/54IqE5MioACBSRJoSGAw6ecihcdCuhI46r6QEiwz+w5S
n+bNkUMFKKMBfxgfNrTPzL3xrs3CYIWEHk10oFZIFwVgZa9W0nTlLuRR5EjdZdiX
jGKOuRYOgsKvU9rTyvTTt1XkFzHbT+6UteDRYJY25DKfEUisWUKBFjXAJiCEq+Vm
7BRmWoNV8BkKDZz8v1QdBLoOky2M/kk/CGpcYRcTb/bt1h8xoMV6krFJjkXdwM9b
EHEWes6TpDDHyhQDGGRlDfsEjoiz/YZ3taJvnWumAsqYP0oQAEuPTh5EXlSjN/00
GAeOM1t8Tbz+5ssYKpyaQ6pLi7dD1PQApfXcPt2IVvnNagLrNQ4mBBmbTbjxKEkE
WwQYustqOmNrtr68FxumHx53xU/htMT6aYzJTbZdF2gNlCYUFhcHW8Yyj2lV8kOJ
OKMDi5nfDr7oxlbKykYepMY7DGlktvh2dAC7HA7Dzd70TZHnqtx7Bm2FhbDzbNlf
ox8TTY9vJixgeRYvwnLPT1tVkO1AVA59Ay05pALJOWyjIJAf8/Mm/Z0fzM0JfCSN
ZxEF8bDE6xf5TCQS224RB/d4WrN9/Kxu/kV6scqWrLMZ4TFKX8F7QNg2WYC8nWgc
3n6RQWMuznSWRjeNm0EKXV7V2yvfeFF0FBtAFlWeA75t/genkmnCnygq7kvr/YLX
v805C2a/D7IQOUTtC9vl7NHxmAdCziZowN+RK/5S9nLKfCSurTeEEvR2ZU4iIuWk
AZd6xPI0G1FdUPra/1L+pbfDExFbAOmsO8w9pI/F8a2sBKn5lOQyhJSgqVUgmixm
QnBJ2hXiK9l6GDUE8piYvBM+a4AB3pVkaj1pRR26I/8O/3r5BhQkGLZD2domePGc
+oMawKnKbdT84cCQknFU+wysxydrjm7vuL3VV01UbBhwgdT3LF8nBHH3qeG+lVbZ
V/z4liy2faFSjaB7g8B5fZy6v9xHmbYys1/vx3aH+tTqIFdm0Fst6tKf7Lu5oIW3
B2Fz5FFMc5STRXdV36UA0loGyQYYYKoUg9KB4Q60+NQ1r5PlACld5hQAqcSBAY1w
JTlvLk10oQT6ZPoL8dqu0Z/krSIKrHWtdaf9FQW6btIlrdHy2Rxof7AR+JkcOazc
59d37Mm0flL4u79y+0ryt5YZ1xThY6JhMw2FsQlQ6o5S5NNMYt7F9kI7CKhKVfQt
nHPx8CSpxTPgs3196PJg82Hsr+8An/slzgCNv1gkRPxrQ+RisKTKRfq0mEJwM67W
gmKdVYUtxSPyT/5NlXBBtXaq19P69VoKPY7ZTZykmznEXWL40sK5y027WwgllDlK
LW4tZ30sdni1FaiCDtOYChHzS0tjZn2+AKNhlx0SvJWSTujaJ9VCUT+s8HbdHq/V
5hC+E0rQ3Vcyjrq+TsEXG7i6HCDcelYQfWfLPA15yUBNz12Lrva3vVFDLdkTfRIT
MK2z2ejbWqd+UyFClrUcl/6/zgK0qHmyB5RulXUO/s79cSPXBNaVAfm3Ld/8WMzE
4q5X9VVNJYOqz1kd3wh+Y4ZA2IA5QAQu27IVWCttgfNCf/oc9rG6A1sy7eY9jUOB
gibNbEVlfA60AlvyTl/44NwcPmctoECQW95BATFNKVmx9IbpdunfNG+rVf9IYgzn
Gbb5IIqjRnqD0Owfrz6IEK0HCmYAk+sXuYG1qZyLeRNv/rHbJot5uF79Vl6zjF6s
SB7mLPmV+wEe0wk4fmDCNUYnaz7cH631qmXkrDAUO2FVdh6Fq7fTkKLvs5x1Jgdg
IwS4+7+6WIobBjnvnieK+UJf4A/5leTqxJu0kKLhWPk5hAQvLbCNAx3DmfGtAnrv
9mQDcxP8ilUKQHPLyXXCbtSUwgwEdYOjEIrejAKgBcWTwKSZwMWJPYzUPzEGJGd6
OXDuw5xU5El59hHztfLKLROgDv9ircqUxp8KBbYw7OETrKH4ph2bxgjJvigPfMlA
0gN1IRmNChAcfIeaNsWc+wbdZlub9VLQBM3BYfkRIW1q6QJwf3xQeL4zA1ZuPlF0
0zhOYAshbcX5YQjIhQLGuUw9JFWtVuKKRJkt6H45ClKHTYCQYVcaaTEclQvI19vS
Plp1CMS3ZCfO3I+vKGPCUSMXOWXLOuKhaNUWXjHR/MNAgx6mtgXuuU96PbV1Pq5D
/mqmWTf1+xpgsXeZGtZFGqz3os397UmWuCCKPR/7RKV/wCtdYWQbmyL9q23oqdMV
+1GVdy2SlsUo5ydToOUM6BZK+OYrcqO456JYDw0wgqOxE4trj908xwL++KrfC5H8
8O71SxItS2II2Q4OUgNey2P1Mf4OMlKKZCgkrgGnzeMKWt2fQ19q8zFhzi4KzHap
GuiwQWzU4rlscF1bbWmxsBzFzepuASiR9+n3gzZKDoCeiaD54rmmIEdEglyXa+W8
L6NIxyHjF7MiZGy7P6+xzYgxOCdSnD3VjxhrL4Ddjz/pwuwF/ACfv4C4AFZdSsmF
bDVtiPpPCcTcwBuyYPvrAEsqvzfpyGdkIWsFQBFiH6tfK8R5wMsvOEw8/AiUv7D/
caWwOhUcKVDArY9fWEqGs1APw0B1cs4hj19J/N8rLwusXXWvfIcH/Q5AH4YvkdSD
SallqlVgDtNnQioXqsPgxzrZ87oqUE+EWj+TGJuqGS95j8i02bB05eBURfC815L7
JmYsjLGXI+IWNbeO/Zs3I8fIss3ZH3ooALJLJYqfJUqwiwQwNohd7WzmtxNo54nO
cNlFlLGbSsk+EAJI2Vdr0zExVLYf2GWlSOoSt92+EYlsVIleDuPqEsZzE1TQBxOs
fyADLQVVFpbt5OzNHuSTlWjI9ffsZUiIf3yuLfh5l7zC5FE6Pu6wRI7Uo7J1xRQv
/S7jI73mHIFLjXVkRnIUum7VyiYbQkuHpBTbqh0ImLpfQASdE/EVt0tfblfF5Baj
uxGue48vOQPrtlB9idzPAnfP5GvrpJLOqA9G8H900zBIYlGKm+t93PZadkR2Rlma
i2gVx0UKjnJJwhMn5GxQhVULzrzzEAny2SfK+FbrSsm/1mad/N5098KMnbsOXC3C
PE/h0k/mSJtNVMWW7Fdw98Ko9LsSTP4pvwVgLh0Eqo9qWZI3ORHEg6HUATtfihPo
p+OXZqDmG1pHszS2Hm4jFhytfdiQhpWRrd52aSesFLpSNZ8rbqSlX0vMGunqfbTI
sdcHROQiz4hs62sPFkja8GzO2p/dBUAmJoGVB8rx8IXRK+3uCzAlAc/GzW1oUTeQ
TzwI6olNek6XadclGNsc/pQ8q0TsuIjgdS8K8LOiGt5ZOf8vSA51Df+6lkQAr848
oNa7DWU6wFl4zvtyNsGgcKH+/7K1O/eBPY+lhDsWcAmPqmMHYLVxBKVtcOkM6iau
oZSFG9tcamCAE/pEy0AQ367FJA4O0GZVOwO1J6EHZuNwpthCi9ATxL9vyn8eNHmT
+Hue1OxT5VEYnUMM9JD4FlzwfDO+W8nh/8kt/9nWehptaMtsBnn2PXPgW4jxHOH3
/ksTefTa7KxPIae6AIAAyLG2a7rQCYmUCMUPlLIKYb7wGLOdDWKj38YCvs+mkfHo
1a4v+Q2RDzHRInAR2utpfUTMfXhH0LPQEQttPAzh8Rjk47VwFn9fuiyqe4v6iXIX
o38tmHawXfI4QkVPG1PKSuPI2tv80xRNeWjVgH+P3rPxlrSSJlTFCcR37UxsgZHg
SprmmYrkuDodsMX0Jaygw/G9C3cTm8ggbmKT0pT3NvKWqPXeVR+9cbEaf1NRZLlI
526ixlSqrdHJjzPBTfHiyyg9UqYrtslo50yrHKc0zzkxgitm04/DCAq7o5xJcL1o
U0oyPyl6ysvdxXINL00Zr/RQPJSNnpvyGZFr+5sAqc0vvzEdPJKNZ/aY/QoHFAJA
BI4dD01pOKxCb52iWfDbbLFoiDTtBJ/72gqfMEYqTcRvV5yDVTHogSVRpuP+MC+T
VwD7TNgtNVLs6XTK6dwBt07TmyG0e2UlMaWjgAEA8Zl1VdCc9R880JfQ1MQtbDMX
QbYPQgtmnRO1syZCbI92dU4boJOxp7chYZahBHldzY6qpqw0SyNnGkpTSITzzwHA
o/NmtVYbkA/aVhwcJC++RvvUrNuJ+JFb8250zisfL9OwjQeNMR3VTjTKUs6Ymq//
izZsfTKrpoQydE+BXYPFxDWcAg9/9GkIUVqt6yhGJENa0qvG3boc186kP1pjcGu0
X0DMZOx0GFv4qN05c4xrsxLtbMaW+vJFfHPQM4VJ4oLRjLS5HtPaFAUn08g/u1Va
4dfOHmEeuGC0AMMV56+1fB8IkbRhyXIaACp17XG1aIyR1BQAyLJHL3vs/qEiK/Wf
DDxkziUJ+u9IUQwXNQXF+fUQ+F8aZzqC+k26h81w4dzD02Ua/nQ17fTOMwhxs6cu
ZSuZ8asqR3lmlEItDwjjvUr84TwEboSfOgl9KuKm6sVIul2M39+hUkgjAn+tlJkN
thpNnPBL1a2tQqCoPZt60leefpcyNGtHqLTYdYabdx9VLBk98tSMjXODRCdQCoK1
MRSn4JeOjUlNzJN+z/aIIYQVJys7UI/Pwcc6mi2qrzBgRdc5z+uqy94NGWAzTwe3
zEq82wuPK/h36J7yXsAZn1jL2PWRPiq1dEfT2YebnrsdlCrbUwsPnUJ5D30ERxA+
BE8I7KO9KnsCnJgw9a6CGCCI6eUKFrdVRL4KRnYHYRUFqHuDAKITtyIxi08XgiNu
LgQ3Az/VcGxERnAUzJn019j8gVJXF6bHqPZjcOPSVy/47DPlwtWl0VN8NCRo5IY2
OsXE42bZ0GrUYX95D6oFg+ikpinBOTF27Q+0tSbp3cnG77q8vuslTWGhve0fuxBd
84453fQAJfhN4t6cBjbdFxp0MgqlJdhCPGzqq7raWXwBf6NzlEnDb6l2k5gH5eWC
g96j2iFwcvOCQ5nfHywXtf5L4qk08zwpluNOjGvecb4rg4C5yMFyqUiL5nsWD0Do
bt4Nl72Hihyqv0F5MaC4vNAiYWni14ScFLXmYtA1GvohIZ+XyaxZ2iV8fw3RIP1s
ZUpxKL5AT5Vn+8+ghV/Elxtksx6h5ryBiFV/FAuzfzPRESoK+CS+/Jy45LzuICfL
8zbnAD+aW7g1hx7ejuFc/1axHMDLiSveC8yeySOcY1kdQBFv6P9eTub8hWcEFUif
Pt0n/Qb2UPVRy86nUW4rInSZ7d5Sja/56LIVXq0lLv5xXYtxSRdyvLTkBGa8MQ3V
0H3LtepoDBXUzBXgnq5xRcw9NoC5usVERiTwV58UqlV56TqLI5R8HdBMMSbnNvDl
lJYQYFhd/wjQ6HQPTdh8dK3iUKbM/D2iPoMZfARAyTLQ7cpVdp2/pNdt7huZB1ev
aVVQMjNBPNzIfqRV9NCSekAnp2HrspylbBW9hQJaZqIr+wg8W7FYqtdQ4xbHGscn
Y4N6LklU6X/x8Lg6r8Nn+O5k7iiDctcSJMIjNSgx7ijDGuN6GlhuUNrWIzd0EHCQ
bad5wBN/YQRQrfAnyProim67NOAJLPdkFKpCY+7Hz/nxOhzDZQ8xGasD8ok/k2mk
5oGCkXcLDjRu26oStCWGd8quGG5MnvKiNHnJ0/WgzOCZbtNQ16xRk9mFfINaaCFY
AZSSvIr1kLO9cdL74max2Z1pglMbiK+hVkdhdvdi93lesu8+Q6djsNJNrrekffag
Jt3O76rYXd85aiBEn16txPhPqjnrk+wlf3jRCneNkuwpRkYFWeTrg8OtauK46waG
6HJt1+6VaMIJIwnZd2KWlYt1m5wjKiyVnpRtVehOedX+1DB1lYv809Nx+9Q6iuv9
R6E+zLXhSB7Y0mUOj6JVFB6AQ2UuLW7IbX4N0RY9s/xBKpIMSw3E6dc16MgkkswI
WpSemKd00Ol5DoU1K4uoP4DH5rpNT+TWOri+TzAbvYpl59Mr4kjXjhF83ToT/YHA
TAi+++W6X5PrjSV3nw9hqa204mLcPleV+A2T0lyxpg5ch4RKq4IPCg4SPAYLjLMb
VxI3VmPtRlSOOIhop8Ljg1RmVWeBBROiql4w3sPZmJUv8hLP0aEgkrFasRlgoPe4
P7ziuDesUY8HLRv10cgy4j29WfwofYUN9W72wnriVdyPy5fihXDjvuaxpks2Q4VM
rEN5sKJQc0KhjdnFHYDkiADUeFYOjyaddWkHO8Xvx7cyVLd6Yef4FuxODkANR3gl
CVMlqMr++QXsy/cy58ozwq5mDobALoW2vDUATx5oIJ4sOld7hYwEQ/BdSUgSKuQ9
vEz5gClogkc17MUBA2zxjzr6Csy3+25OFLr62QIDSJT8MxiA+a0xRssHtG/qvt4W
n59qr2xJ3LDMZMMKIJpWwYMjwFHARhxgiqDvkO1g5kDY7nfGdCTArmIJw3wO1afk
IaXDyiDKFBnyty0oV7970LqnKWkJ0PCQ+BTJbut1fQoY7agYBMk9ZQPalnuvOK6+
b/xCFUMr7KqHu1QMvSKH7OdPD93EtqSRauw974GV0/U9/V76kjXq7RkERoOSOPXk
dbUfY3/aUdxCOnLo+APHIYotak8JdUt19zDp2aYYNczZcYgCw6NndT1V2eEgCIEg
96ZwAxfEMJf0ZHxMSBe6x8HgvoJis3OfnOubtOzPoA5kQoVipUCT4moQIirjvXi3
YZSrYwqEDrwjGfQBgCjgpgMWI+8PoWg2NgBB9ivriteU+xF0eXRTgU0EYgKhIGgF
E2F+45qREAH33HfQB0HkF1ZyNZM9V1C8HHjyOBASGEBCf0ifa1uKrlfs06GK/JYI
Y5R4SmTG0SlmUIJmppCsuZQhudwBwx3YM8fg24P56OGqkCPVseT8zAfvZ22+dYrT
OmUk3TQ6BtO9Y6mt9ZxRcd+mjyI0OvWkRXtqLxZil7IwbsJQ5HvBb8/Zx+hz/A2u
QqzkKXrySZ8HuTX6HM8FeH7G8NPrhuluy39xO1mz/iHeMpaAnNMq8y2GcHw7/pRm
GeSVO8PKaIi7yapi40oxw6JLMlVEM4ssFCyM8DbRB4rTOFQapLgEj3kpg4tV9Gp5
UCj1aiRR1FtI/KsPBaciidB6OWmKF21D9xEUvTRKAuJ/P0Xb6mty75y8ceuUT7Vy
6PwZe0kiDSqDvWe3isHBANaIbxWKoZkhnfI7lddjvWOcN7cz0vuzIcV7GR1bN29m
niz9zp+CO3YIInflhS8FQCKKSrX/AmWKFc5CiXQeVA9UU/rfJvZ2bRdcRoDoW98s
IsZu2ohygaq5IbozuGVwnbnu89WkfYNhHnmrjKm8T1BHjbu+PlblsYj9ntejfAOw
UJ9aCfulpEYAkdH4Ifj0D7X8p0SXYCM2XBH47QkWroGOpaZo0z8M99TfT/5yZyQW
Xgebsn+V0DWN4cPU9qHah5ahQFdLbEYJmY0ZDU8n8SMC7h7fgNAY30eYMCScGY+g
yONu7584Pswb6xWA5HNksI39r/v8/DEJOE19jk33qF9ITVoYWsspsDPpCnainMq/
JsilSucToGTahaKbJFweWn1MmKrKvmCvOrcUz+4S5ARWwYYaK6TJZbH2xsaoROfN
W9JNgL8E+mUOfA+y+dqXDurxfFwFzOw8XwfUukeKx8clKyh7lMTieFmHsnfjWZG3
ha4w2cYh2be64mY9awroRSLyJaXul/l2fmZZiS6hIEztefu7FNFDXc6eOgU8pjOR
YpcZipMYyom10cBN0cG4sKd5yPGUBt5p89kAup6RkTiUYPr9soLQ525VVFNVuPGi
dEPMf5qWfPFO8arhostrCQUeymuvvq8ft88PTXBZjvB2ZpnCj1nU5hfDosuiqG5q
cDWIPTcRPn2Fm/BRzfiAM3hjVYAaWY43DV8G6OV6jBQ6/gzjbGG69XUnpc/dO4xj
hQ/0qFqRo81HXu9PJiI/Mz3W7LCqmynYlgxwot6ibSt7i2S5438sbsHoZa/WPFc8
Xwc0Pb4Yi7M1FiuW5FtfnaJovHj5izw2TZadUseY9xPYvhTw3PDdhwHwNvRxL62B
dV/bPizHQaJPooUQoFRJeDl2GqKt+l5fQvjs6MYULdbztUlcy1l8+qGq5ZC79Q+K
X8wogxcWQ3EADbSnt6tfitJpc9lPLfRgO7DfNhiSUDVIjxUN81VSpYZQIzRrtzav
4cm9pF3SoE0884Rd0fwX64vWpzlLzFFlQYPBsXXX6szkvFQw7gZ5W/bOQK3Jo0b5
dOqKqjbJVmaJtwfQcQa/wNlr3OySm2zIav3DZW6DWIFbZmHlroQjt+1uxKnFtKX0
DIwgd4FLxuZj3j09Ckr4U9/st+ozVzSByAQ5mSXIPYlfUtlsJ8ZHs0TiYiR8giQF
c3nksIgcYSXcaLb5wPade0LRN7V+lgREViZxObaowDTTXe+ivv1HYKqzFMSwVFP4
maoSWhyNkUVdjWOAaXShXNIfxzWvl6zo6sC9Kgym2LEEVtgmC3Ix2zoPudEF9aPf
W0fJTqHjVyJvAmyd5PERTUjhmIf4k4izt6e6hpiTT0uSjEwYvywyRcZZuGuTW9B1
OcWJ/iYThQeG7c3OnT78CTGcyvc6/xE0ct+d5dbUifOen7WXTtCWLQYfDWKjz+mw
iaqjpPFV8fQ9CC2urFg5HpGf+vMb0MFFW9dNjVrkXNznc6uw2Q5LUZe6ORFhcf0W
qnelnJ+h9FZ1XRnNJmUyusu4OGasalW7V8WVOgN0WQAVgpIyP3INFSpLcNGGEqO0
vSMdVHY6IH8nOroXhv1S3mQLtZnCihVLUpLAbytQbk5OU76cYEZRXscPTOOArktM
j+JAxSoKBMhWa85DrRTjla9I71sS/oA4C7kMP3kVOdCr0wPtbNl7mKkVaU+j3W+z
jHBwZ6a+yUP7LX2Z2+GTv3FKn0h0cE0oClGw6/wYnDGyDszvwgY2hLm/YRgdrBjB
Se1qMJhixpNe3igiDzpyS7849S9IQ+c1Hb7uQZv7nOe37t5FFQuxQ2oOu3zbP09y
HgYPDHlMVoVqvDv3aKBQLzLFzvBdw0xpNkDUCzEMZkOPNtRiWzAI/htsPGpUBatG
s0Zotty/RVH/tY6R3uMhS/Cvomo2ggm17OWP2rHDX0PI/DoEN0rub6Yx0uQ8opJ5
93XylCtVgjuJx5oBo05cuSZ7BpRsMiDttoysmNNym4Jyx3Fh2cMX0KQcJh86rVSQ
51RReA3YF7tHL8e6yAUG3+w2yLRl8/XvTHPCWlRBJJtyKmqAiKxKqymXDf6VEoAI
9JM2anoetHJGH3fu4zOx+ibPTxEVBJMmlrD+kX8tXJYTtOqqSIFkp4gD+znQt/C6
cHODAxyyB49Jz6IOT5xdmq/od3pexMAcVMlOO0kNG0M9H85SHY2qmmZDNTlJqptI
hQi1YFfprDVxj0K1SZocnkEhzBxIf6opW5Jmv9HMCNLHmJtuncdoWPeCOr3obExf
a39nr1Z4QhLKvMoqt8qoSdkCWkqtlSpDWFJjbVUQNeJKq3qYNeXbTvpzu2YfQaNw
YkYrT/6Uo5BywofoLNxvLEV+ArRd9ll4On+Dz5TXCvpHbRXwqwPEevKnRzKS5tS/
ML6kcQOG1hQzgIzsEG59kHlPW5ktBOJ+5j97QwT8cLRAawHN/XfUpB5CNTzFAXx5
jo1/h/aEi8UmsIwGE93YS7TlprxCkI5ihwN1ejTve9mBHyMj2NMqZ9OlO1M4rmhk
DxNsBKtA6497Z1VUKsqRlSlPR33DbG3/BIMkV8ijdzdrCLiSNID1GXaCUqsfTcb9
rr5QJ3kBjTdBWwIEKpVZhwQrmdm3cvmTeOQqbvh5rTyyYe02/DPgxf7Q8yKDaaft
HYyYjujMtYMDdQMeSvtKdLcJlU0LSl5KkSLY5n5l4fxnK4rYe//1UPa/gJFu3dzt
w+FkcBn01AhOthrPkIN+nWG4jpTH1HYUhUokJfy+NVa5coL9U2uA5QmACGwgde8Q
iaReYStmiwpXndV048UoCBLwmQ02NA2MhydqRTrKLOz4suV8kdG0EAnYRXMt5YS0
Vw0AajzC7oHTxq9b7XCclkno78QDjYWFmNCdYvITcaBlzbG2S28gv3AimP69FXvg
pmc3zysj5GJPE+ZAKVUUVFJlTc9AmG+hOQ4F8Et5T8fjiKF/6cvW81RwKzLyJtvr
pvzUYHmrANh9OjEHk4/5Asjl1xuRA/eS/RCv9l98p/RE6P+GqSDalJMBOH2uq5q6
tFK8nngK3NPLqCfjkQI/CY3HGC+yghuVMnQZFYXKLLogrnaiPmzKB+GazNgYV4Pv
VSazf5YYPuKaL1Src7S1E0vWj2EMskRqhyNHudtQV8gAxnYjDXpElVYv2kjLi9fV
FBDES10VqvWcBhGjtSYy8y7Jcpr08TIUyFkrLGIKibTI78d5sTcIIUNCgOuH7z3+
NstKWV9CFuajybvgtDXNNu/SfKiGB0MPUsGTD/RluH8px4tRRosVDU5moutKJEjT
PZ1X1tesd93EJFVu4fhSNVDndJon5/s6VwSNt1RzFnyce3irpjrPEAscuHpkFKBH
XVcqcv4s8SpYPcG2zScJ4DZgY8OgJD58qrARiDzh1NugIaNMo19Q+zsjfGPBtWrf
iOEs8zyBxJrlWhIeU1j86/l892cDIrekHX/6jWcUNX153n1cm0liAvbtdI2RSxgR
A8s46WqHRBEjSoaqPezFMCTvsBDF1Y8mZnYShAXAQPuG0XS6lky8iJ3hqFplMJDs
zHMnRK7dkMpoVonwSqwITjeXCDKkIQ5ZJUiEjl7QjgnKUzRScZmidxBd1hGfPWlr
KN3jRAF3Lnp61lXVfT4kGYgt2Uue5RmU9TbXyoLUJEjzMubQ3hhEK9bhgg2r012M
xgrkXlm5V6W+Iyts/A3G0yQmYIVR1hlRt3v4bqBdPHYF4LWLNstnI6GHmdghaxgZ
ctt/FjovxX4uedSkdXM04NbhcTI9RK8vbjgnfqMS2rQgbT0ZlUztCODeht46j+e8
KUgqe4MZKHTN85/2cT5LuoDfKFg8VXHE9CqL91KB/QovPrwYFB8pMS7wKLUcNscn
Laj+jGqx5qwiuU6Wfj4RrlYuQbPVY8n1k3b9WIuUKdY9IjPeumjTSeu+xjxai4w/
8pE4OUtIEi9rYFW6+BDEZ1dUmyqi6V3pEOyptHbCKZXSzLmips3M1Zqzh1qfp/rm
qgouhA+gOYcbrfDhjAMbmSrxkKiLKpU41EHG8nvkd76vpHcfknRrTq4fOHyTvnd1
MousW8h4n+R8VjFd2fAQ0fZ9r6Kh6pJo3EMx63VrTnVgAm3aJD3nJ6lbWFhCGaU6
F3WjQB7DC7Fgu0AwZHDZ0v3nDkq0LiSfnYmnkcAII9IwrsewbUHULy9C4/tUscls
1rmSJxmNMlnBiba/Ms3zTrnFhIhemSWLZ7Zd8CAq3L/fyQuwRYJWTpPJ/1eAEayE
VlfClxq4nyryMfPhvgSKH3W6EASKghvInCNfYw+uneYcgaKx2kng8nrb1kYm6r73
o29++IFYlEYB0cr9u0sRbyBaTuqvtZk3xEnSOczRVfzg3AfVKXyOURh1Ev1C1iuW
d/45Nl3bmAK2GKcivLp5oBeEhCQ8A+0nYYtje2PG66GzLQD4tlKMej1rT9GHCVvU
SfU5AZUN3dPlKUDL+F/3NXV4AXMInLbON8DzpWqV7xQtKSFRGrd4iY9fkrnduyYT
mUvj9k+GFVQ0TtFfr4/seJmXoyt7xD95LzsIO6JhiLNO6wSA5f9Eua2z2ShWRU92
dJFDzpzqr7jpbg2mgCF0Qc/LXhAyBYtzbpW7WbzrDwv7ym4eK29uVSLpGzpH5pce
KXYw+AbtWXyTBlMzRKahFf8SvpIwpn8SomLzAE0HAItqdqrb5hRoxKLC8/Byiu1e
xmFASWoT9BMf0+C2Qat3yZg+4rflFkUYnOTFd7SQGZe+fwv4C/vDnHZlTZXoeE7+
7TLEKn0ojQd5NOWmG2V8y8DD4nKv6Xdo9/i8V44c+hjxDFrzv7VDZUTVm1H7wVh8
9MveoYVFvZNfBUhT23dPgVqR3P2xn7XNmp5EC7xn+cdgZOoXrzlQu55FdlNh55mX
OLbQagY0iAf2MfsWxE0ErgQoKV20Oz8f6V/A6eqEFihjd3wGJUsjPN0Zw0IGPI3D
P/Ll0aRpsCsSoH2dmiOCh3CVqkqsNQNpFla09REwQeyNdcLaU1U7mnfVfiT4k1pn
5n/YnFECuzh6+DnkIGkIbzVS2LURL+/+XfqHmacYDZ2kth1LnO784I2+F1Oq/guk
U5IESPQ8W2x2GlZs7pH3fo9esrBmIQgCiler7GqE6WCUiLYOqWfn+Mxv7mlgjC0Q
dXN6wMLyvKN3eYKQyB2WZZi2E5vcOJwc7f2EP2c9NRHBDyWvA0NLOCiwU5wvg0nV
XXMRKMb+ll92QtdMrzx77c5gWJAvRocQ986YjBh1PBCANZu08sm7nqibilVcBTQt
HX5yBfXqHQx5XXrLY9kU+ijDD8OR3gzNnYmyaqBZ5kGHDQXo1AfJVZAIcA73nvWM
wWtHVC17C2R1EFFLYhADOXC/YjGQOggq3tTB7aPP4kPsyvB2w8JCuUd38ekhL79p
FefwnCYiRizE87TA4r7pk5gb7IVxyGFqSDAkxDqsBvvp2qwsmyP0ZpyQg2e/rts0
SFDEB8wztsgluhypOBBFHU1rzmLKwv5ZJVpFb/f0nrQxqoMNdeW71+dfdVitZCvg
ndI5CPFPeM8W8CN2OxBhSn5og5IE7imF3tAyzeopxuefvUTtncWoOdoZ3muMjvTa
fvBgcGHQL6tU6snKudu8JiZkU0xIkCSTpm4PliPwIoprzv8/ERGHjJDWFjzE0VpA
nBdANUo6Uye/9WffvpNGG5eK1zjlNiEIoGWaEBdrucKGFfV1i2D2Vr3IsrFhY0xa
BDZD37cPLPFyPE5NSpKHbKoIPNXxX09cD9Qt0twHZGkBWVHjB1Gmp3z4VOdoD68C
JY/BWDjPV5krgOfeV43sTRaaQVQ+6yiARhbfK6jdYVoaSSlfwMafWuJjxX0d1EU4
McvDgvD49hpAiRtxMLWAcV6Zu4o8kGqelgsOul/XtxTgAAw9GZK1wp/fvXVrVZnw
s63uOkjz/tKnSanZGr5nmtX+AjYrkXcdIpGo5DHn85XTZ1lEtrwgy6+TyhrP9gMk
GIyuuDkLQiAKFu3prjuK37Yw41OBUBgeXGEdUBrZ5SxBb+JqeAkJAtcFVh7ILesb
icdjrx5vFhu6e6G9TKai+hlqLEU9rOgNQxcypIyH4YI563DcrPAvQrl8F0AEWzsu
cObwqOEqkBIJ9LkMp8ELs2kvbLQ40vSDoOiNChHvkXo07Rkx7vaYsu3tIR60qWq4
k91EiNwHLqCNqGForC27F9W00qghsVqcJ9a94e/acxeU5bzw/507iLMmGWwVcfEs
UXf+ja8wlqVeS4O4jk4ABnSwj/zEHFwzHb60RmAyN31UNzb9OYjt+UH65/fj60rS
/VupDh3jCwpBIyyxcFyB0+eR9xnpkdhMNfRJDxrdRzS3kH6BI55n3sz6jVdONswB
8U2LXBhnTLT8cDO1AqEXqhY77rhiKZps3l1c6ddnA2ISx6VW86aZoEDBLKVQpzAO
9MKFcusuWQD4R0UWL9h6ER2C+uPzhL+MfeqmLlcaulOTrYeLkfvfBHa/bOmdR8y4
kvNLIGa4piYgHTrwE7Ss6QvqzvZtjMo3pMqjVC1hUQER/ImKKeLPtbCbhmiRVkds
uJLRM32CyXhHUzcob8hMoxC06oFAP2UTvqeUrVG/LXj/kjDP0DBRn1nRYL+IEg4q
tZpU3vbkAV1qUfZxVteBYThNqMBzE7HwU5rddylRw4DmXYuEs3hHueV9t+45+3k+
JNgKEs0jMASg/Rhpy+Armdn3dKSvRxSj3L2IcQ/xskFuHgxTDjHlnhPy1vBA55o7
BA2VRltLbWFOa9TiHEmUCVt1RYd6k+ruKuUid7GeFfBHpOFXfZ9qDZf8e8frCz05
dZh7yBPiVpAglCB/bBsn5FsENQb0zYCiGuuy1znM3zKCPMPMsRLbzAB6a7RPPrAd
aJxUnV+ZA2dzhtoA96lF/jt2/aeWP6RuEBDDoKM8A/9EgPGlLn5zxFoyyO6YAMDr
yMys1eI0R9RsZo9f6QsuSOA5wsW72B/JrMMfHmSJwjQp3SOIDN9Rbuf+vqRaA5hD
yDykIfr/VVcW+VR9PHNcyBeZOguDov5iOHTTK7nDmqfdi1YDqNnpGUo+Pgo6Rk8G
QO+A0qSjp2rcPx3nBqjrC9KJBlSOLOA6h9rG20PKHO2Kl02EwRFLpnsJ4SimHiaV
fbNLDDrjjoFFULAsjSZALzcwx8P1u7sQxbua6NnKdkG/rAtZGrO391ClyyNjDKcZ
/FfamB5YK7EUMp+cTsIsBKwgXZptQuDNoxJKK2JxxACtMRDzxFkcT8lGsWZoS+yi
wlkkspYql+mjexOTsnbaIo2fEvlEWHPfqL8tPqXqNA9ptL145dXQxVCYPmJYAsFK
rBXAI6fFGQ0DrkJTGGiQBsFj7ohOko56YJcv2Uk/QlfosB0G7C35/oNLUlemv9VB
QMQ7tVSdAcsoyjCp9cfIRIaXS/livlrfC+f1RHblAH4xnde0s3uZmpJHKz0yjPo1
aYmdhFOiHCnclpARTSid4iVXQ1lSHuohfOrFelW3BjoyF0zLUWmoYMp0wxRIoylV
gYQLtqrAwUkeP+U8kQKseIUy5FicZRsn9bxti7ziQIOlIgAorzi4r12wBnag36oF
RrOBEkxdyCa8mkUtPBAMCE5BvmSVIYGbovTrxfp8NjC15KFvvXgUpoujL6Gvp1sL
p6VbLKb7QiTSr/V2jD05p+yVDqGtWpOzmw9d2OUx5bWDz0hAZfGEF52cbYwwcp0r
C+FkMoeLCziOgp3QbKFX3cBypd+mbnSMPqQb9RZQPa7G5nHXTZohsmTWuLc3SYt6
uwK6PQqrFaK5maLkMGyntK+lj0Gn3cgoZnQwBfKjeW4wmKaH7BtJvqwvH5PClRkG
bJxhSvvQOJMVNf9NDgOH2BA/HLE1yHRK2FdgRNeP56st7KUIRCI3yIWrp4zcD/CP
ob/6vB4Ut9AjEOZcWO3VR1SbR+6Ja39vzUX43TeJ2att1jMEneYeqpJ6hcZ9qF0Y
AJn3eoLJvPwnsix1smrYFOVXTXl6LpS1/Q870EdCXfjDpdmj7uIypPyP4xg94YDN
G+YF8sVOBO6InfE417WMjc0IYf3vFGKa6udksrGkWcKecsAkObkivnYegzG93vPH
pbZUlvBaqTV8Te8vOUGkWfypCyyUgPxcLwgfzCisOHdBLI5Yxby0eNQQ1tQF9WD3
iDr2K6ju4ul3IdBQBuljEE++oS2l6v/TNf6Rscs1mfV6jA+7IQbpcOCGw3xirPl2
iwEUt3Tp9ME9k1YCujMXcEEzFFczueAOd+tUtY9Koq5Z0kzoGhwypEgXStccKKIE
Ot5ZAwhaCAhMUwQ126O9vN/zmvM53KEG4fEMqd0PI9bFGNP9HH1LEVq0ncCGxZ4z
fJlYyKJqGu3/1VDItMyQ/qkvGodtMkviCQKfH96Ti2qu7v+9krq6AWb1gzZYwuEv
MCNZZ7+Ljcsi3BJA2BYJLYKryWOhYok/Xywd7ENA7Wo4JC9dXH1FB2hY9gVAbQOY
9234Jj1R7e2Q+FYSakBrI5QIAcWOdn3IV9M7nsMNW+EqcqkhHnZB5M8VNGpM8H3j
8eDPInPxXSSy0fmbnWLz4QBTP6scQt2VYlmBrxx7MV3KTPdyXYgyJjB+St4oJ57w
P9STc8Gms3KhVnE6N9mEILSxwQl/CFv8PQQkj7Oz+/52KkE+i2iaPuzDDuLO59VW
gAB1HQXQti5+fqXqIUtPJh19v+PDW7OqpIc5YQsiojjE7isyyFx1DL8LH3yc225K
zDqQGeJLmuZnQ6yyxSSw5rS1eWpJ2JZMI7SdFY1dN3mmALZsl75RU4bTnYSW4Rp9
gPlxQhOMdj9bZgy+VRiEf3MsI5ijlCt3M47Lmi13aIQ/rz98SsafotQHd7FnHe9l
iMURgm1Ri8zgxRp8t+VzPz4PIIjLqYISOlEjnFVz/ysUmmogZVg82Axf5EUNEwAa
VUlxHzWG+Ty1a97wlM4xr22EyZyMEXijoVgryHhuprXD7DMwMk/Aoq8x8qgdflL7
Z5LkwVkTAFtA3qimsn5HjOa+rl+fLc0ISInEn8huUYZOkAeq9VmcoMoTPiSkjxae
TLPoKqNC5x+ar9JPUDxUiw9Quz4Lxnqw+XOrc9h++6P8Iy8wIplc2+Hxiei9A0R2
92qY6CadjDnsQyllGfv8Bqzg95aqisv4zoSb94hDzMkJGjWw6aii1NkONO2McQrS
WX0Jy3Agz/eHWsyXybL+DH552kcew4jmpOifOg2c8VRy210znuPF1gFhDyn8oeTG
xT+WOyTx+dnuYyu1FBSKPNpu+W+OwjNpUJf6EHxGFdF5TtbKJztHjeeLn5B2NXcs
sJ+3RLI3iWYkDTorRphEZgjCefCyuzWC6v0PHkT0Wdu0ndz9I2jMezdCd31gZ0wQ
/nmYTOHUtSnZWn0/79RYPrhCkrAXu9pdG9HgCpgW9CCrw58vI838rKODK1J9qvH1
PorgxmMIwTQUDbmYuGcFRSWIhQMmWRHXqwcz8VmX9EDuysCA7MY6gqto7V8zyzA2
lsYOo7X51MNTd9WgkdJimFDk3CdWOPUP2RsFyXmHFjWkzCiORK7g+qQk+qPnyETB
IbRBprDFv+shMpcmSZqtpPktD+IWqVKSzYf2lOZlh2kunH48jntU4nAQa+EMaIZm
FHMNXewmGbvf/QMaa7P+mShza7vo1D6ZefL34AoDxZBA6s89pmxCCRnMeth/uqLX
6CXR5ZZCP7MowJKt3lqMtRQRj6NkBBVkcbtxBXYkvtWzBFfIIoUAMFAOpoEoocML
Qp+fAVmvYcdlBlNi+BxlHxF4fbZLhqy+3wOQxbdDJN26o76pFc7KOVNfUlrEj2ri
DoT8MfmJGuBvVstq4TgzMIBiQL9nryHt9JTs+Wdc2x6AmBLAOjp9n1rG/zfmjI2Y
CTKkswPdbW1/aTMeXA4kiwnU6rZYNtWfbCnaDgs7QMWnJir6UwNJz6Xlv/dMJ8Y+
P3WpErxJsCIBKYD2BONedrf9Ub6RVJL04ZLSUYs1TWfZX96lGoI/ZLvfgt/3LPMZ
jw/WfRS61XKQuB5vJPeiYnvZTb2T+f6PM3XKwTxr1Na9bkfbRrtVGq8qRtJ+G4va
oJiCkRRr5YiT0hir/T7246It0XQW7WVlrn0QwmMBKbHsAF1KRam5aBD3Q9028Mc3
aSLheMPwv75SFPUgZWzXbYLbPsUYLRR5s+nMXcGPIcwB3RpbiRNo3SycL8gSyYar
KjCI1ii+ZM4dS02s7R4yPP8uKdZz4tuiq8miLmQ+ateG1/7xZnnIxdG3RYrTviPD
3etgNY770pGTND49ij0+8c86X0QJ7aD6lkCxu2q52az6We10j/fhb3qwnI1z1nwg
MlL5e08UTqx8tlvduNKONjer/HcPs3hEapexigHD2n8jypFxr7Y1LSItvsFHMQrC
UBHORrAmKNZQF3O7ujGnZEiNSxG2cPq91H+iJVpskHfXWA+SRwvhPVTH9pV1+uvs
FQV8EqmUcTClcX1CodNe8XNEL4cJRthMX3P758g5eNZBxrM7Dy2zDO5lzxsTX8hW
7VkVczSf7ohKsbVSsRr++Ftcmh0KML4q4Po+xgOY44Y3w+we977dNo1FzTysfiRZ
3eDV3P78m+dCFzhYXOjGilGkqpwmz++mnYfQ6hSQ3B4vjpCKllQGew3lPYfA3BXi
NyfwseuTQkcq69Ro131aEynCUL4SeqLLYusNTbpgDJfSd+E/WmUPRcr9MA13/q1E
L4RLhFjn+2A0v65+7o9cjLxQvAV0zrK0CduNVrzfAaF7Xzcy6t//zFK6dp5ypYKo
WvDZ3QwkPUTF/FHfgu7jlrX0DsZJF6OaKdcblFaxb5HDY3Y0E03O67wpg+5LfTql
6TqBwgHcWRk2iaeIm4Y6rN7FLKLXhTR8Z8KyZVy3NTKGfA5ck1RruR/hkviBwvHf
V5iPJ4EdZ2S98Y5aL93TtUz53HuJHC/PjoANHhyQfaN8gpSwblO1ERl366ZTjFt5
MBJFap3PwX+mt2ACtG3WlGgZ1cUZ4rGWBzF3dxdxp3Tdmn9XtlnIv3Qanxa1YKGu
FdeWqeXCMyCAh1CKxlNKcrswjArkwrrujCQ0Vhe3OQD64jHFnxP8hAHFLsiWn5JY
5cHuPGkkzUf/2TgL/pwVlr8rp88ydLhATI/HTQHTEuqHECoX9pR0GhOlaz0VAZXN
7Ad7v+s+F2m1t2c+n7ExnWZs06A3sq15oXafdsSX0qOhVtzge0ZlyRPSCaWOsWWQ
06fisc0Q+hqQr3pnqsSboY/mi1xXk+mgCM35Ecw7eHdZkM5AkjdtnMM5VvVv7Xog
YLhxc+ma2gDA6H/TRGpFnd7b40kByrkFdxjPCTqXB52Tyd/6tZcfXA4D5x7MovIR
q9OZGyDToDDw5GnomTzgEfTSQD1H+Voy3O6pZp1+I2E4A5NQQu3lS2DzLMtSedi9
8BV/5jGUSDKEspIQOJ25s3txNZ8Em7CQPq4cORgXQh8ubdcNzToJFem9SrhbVEX6
qwju3priwnJA099rjpuOiLIqhj76nZE15JVDqy/oOCjg8AvuV9Awdoh0F87nRWs7
UROtgElQbiFL9TQf2Q5J8wC6AdGuyWtd/SQPop8xNj2GFZ3ndJdbvGzn8ioxApS6
+X6hhZs8Wd9ZNX54prSh1B79fkH9zzsVpzpSDuzUHkr3wDDypA44zIF6MD4CojcD
QM47lOOTaBwAmEblT9A1K4M6pdMenpoZhFUlUptFhBLjUVFFATfQKnq1HSv4c6uT
oHYKW74epSjdW1HrYYm1aZlv3Wi0Ar4Ny4Fld8IXltK961yzhoJzqbOtzcbTI+R/
VsKFXiJ5Rub1dG7u//eO2dBfO4UQwHyXKGL+apCorYEUxJ1cTRyVI+xbttAJHctP
CGyKDWLdNlM8dcS9b3iIgwS10YWA+V/0q7OIw3YTPEcL4Byolz+qpUGWno4r23RC
S9avnjlkRsLzrCPdhUe0WVAwHnpaoeNlXRJCB12kfhKWYqC/vM25sXG6XHcCMQN7
tD1vcDVkZ90VeSDafab5+RvVJ5EJdD9Lc30LTVMiTwkUa5ef8qiNZowEmJIR/jt9
fwocpfUW0D2jIIzQTL8pmF3a4lEIxPwqwCsEV69RyGNpaXJrVTKdmax9Bj1mbEoE
3Nka/oykgZlo5BEZxXKkqNOdeoddH8FIiYLQw0VMBr1RpNaHy0VhCdtl7dZjOWpW
NPRdsIF2c/FGE/DyQ3I8/OmP7VKF5T0M/16tDcqXCIyExk6EJf3GpD0prCWhyN77
q5zHBSWl9dqSBDNMZUB6DjRLsl3aO1cjnA/sDuPRZ7cIgnoDKjfsLFjziQHRkxKz
pffV1ioOkWd6v2/0QjCK5SrXTtRzTEQN1cbCZ814ZOelyNv8pQS56u6RzTgKtnHK
sBgSPWnCcaJ1hT0fpnJgTzow0qhEorayKayUUotuQFDOFA0IaHOOWyHfxIoeZy2j
av4Rgu4yznht2J2pJ1JR1LZ/XRY0N2JpEm7uTLXxmfjW/h0InRF9KwivyOizNC1C
LDJJMSb05Wl2lQqKg7+M9FKvl86//xHBzKSaUGqlj6h/lALVPzqug6FPHLCZu9WL
CkzKA7AW52mYAaOD6U2aBeey/BpM2IiYyXeDxCDXiiIrm701+xd9hq12j+skf+9O
/Ea18R49v9I8uYwxK8o+Mk3QVh4xijIovoaCH82U+zvk9mmismeiHN89oD0+rhFn
q7E6h3tKCxxTUeOp3Ma/uV/UuQV+bu10rTemnL3MKGsJGdueYdmaR0YHBj24X8/y
8aHCpE44yRMffekfE7WIGdXYaGdbB0LrQzd1qPwqN8XZa/8sPHXtwy9HwCgBPsT4
vOTD7XMvWzpVXL5DabEVXxaoIEDaUWZdaMQTIX0kDrEFKCka+0Q2fMRcKlG+WC4Z
VjQzX42uNjZ6CKkmRcKuDWKMaoKZ6qugO2ShIi5bVG/IO7x9M9DnO0vOwGZr8CcR
Ot8EPUfduS4uvSULjYoagmc4AVM0VzADNk2g64h0vL3IDII3TkGFClh0wpnYFhVW
hsaiDrMUs56AorT3+WiARSdShAHPoASYMXDpshH066E4TII+R9Bk7dsqfJgL4xiU
F/nIdZ3Pfv6p7t211buowOWyFfv6WwncW6jj3465SKYlHcYFnNSW/b/rFU1TVS2N
IMvCb/QDcWIUeIS4CIX4JZc+c9FiJrDtFiKd5u3g8L8=
`protect END_PROTECTED