localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTZ_CHK = {
  {32'h41deba66, 32'hc050ed40} /* (15, 15, 15) {real, imag} */,
  {32'hc2623ac4, 32'h414ed1ff} /* (15, 15, 14) {real, imag} */,
  {32'hc2a0fdfa, 32'hc11207fc} /* (15, 15, 13) {real, imag} */,
  {32'h4033b950, 32'hc195e4c9} /* (15, 15, 12) {real, imag} */,
  {32'hc1272329, 32'hc1caa356} /* (15, 15, 11) {real, imag} */,
  {32'h413149bf, 32'hc07b359a} /* (15, 15, 10) {real, imag} */,
  {32'hc158895a, 32'h417512b4} /* (15, 15, 9) {real, imag} */,
  {32'hc01669e8, 32'h40365bde} /* (15, 15, 8) {real, imag} */,
  {32'hc0545fe8, 32'h4128cbe4} /* (15, 15, 7) {real, imag} */,
  {32'h40e55c66, 32'h415a1830} /* (15, 15, 6) {real, imag} */,
  {32'h3fa05c08, 32'h41ac8992} /* (15, 15, 5) {real, imag} */,
  {32'h41208330, 32'h412cd9e6} /* (15, 15, 4) {real, imag} */,
  {32'hc0d7fd28, 32'hc24bb0bf} /* (15, 15, 3) {real, imag} */,
  {32'h42621a70, 32'h418e5ee4} /* (15, 15, 2) {real, imag} */,
  {32'hc0f2d4e0, 32'hc21cad88} /* (15, 15, 1) {real, imag} */,
  {32'h41455dba, 32'h4100577c} /* (15, 15, 0) {real, imag} */,
  {32'h413c106f, 32'hc0197463} /* (15, 14, 15) {real, imag} */,
  {32'h428ba3f8, 32'hbea99460} /* (15, 14, 14) {real, imag} */,
  {32'h4191188f, 32'hc011eb19} /* (15, 14, 13) {real, imag} */,
  {32'hc107ddfc, 32'hc123bafb} /* (15, 14, 12) {real, imag} */,
  {32'h41ae484f, 32'h41630963} /* (15, 14, 11) {real, imag} */,
  {32'hc0943f22, 32'h4063c807} /* (15, 14, 10) {real, imag} */,
  {32'hc167985a, 32'h40e89d49} /* (15, 14, 9) {real, imag} */,
  {32'h4147a852, 32'h3ff9b1f0} /* (15, 14, 8) {real, imag} */,
  {32'h40917224, 32'h4109b3ee} /* (15, 14, 7) {real, imag} */,
  {32'h4125851b, 32'hc1250502} /* (15, 14, 6) {real, imag} */,
  {32'hc139382a, 32'h41240075} /* (15, 14, 5) {real, imag} */,
  {32'h41e3f3e0, 32'hc113ea17} /* (15, 14, 4) {real, imag} */,
  {32'hc136e0aa, 32'hc0161803} /* (15, 14, 3) {real, imag} */,
  {32'hc17944ac, 32'hc15a8b99} /* (15, 14, 2) {real, imag} */,
  {32'hc201914d, 32'hc07be6bb} /* (15, 14, 1) {real, imag} */,
  {32'hc156161a, 32'h421e0c1c} /* (15, 14, 0) {real, imag} */,
  {32'hc1f1ea57, 32'hc1a6bc7a} /* (15, 13, 15) {real, imag} */,
  {32'h4205dd82, 32'h4106c969} /* (15, 13, 14) {real, imag} */,
  {32'h418b5563, 32'h4171b387} /* (15, 13, 13) {real, imag} */,
  {32'hc20f2ee4, 32'h41b1ab07} /* (15, 13, 12) {real, imag} */,
  {32'hc18ce007, 32'h3fc39740} /* (15, 13, 11) {real, imag} */,
  {32'hbfc7df64, 32'h41519cc1} /* (15, 13, 10) {real, imag} */,
  {32'hc0ab2b5c, 32'hc0b38d58} /* (15, 13, 9) {real, imag} */,
  {32'hc090ceda, 32'hc10f48fe} /* (15, 13, 8) {real, imag} */,
  {32'hc0f04c30, 32'hc0e90f48} /* (15, 13, 7) {real, imag} */,
  {32'h40972b0d, 32'h401d1bc4} /* (15, 13, 6) {real, imag} */,
  {32'hc195264b, 32'hc1440528} /* (15, 13, 5) {real, imag} */,
  {32'h4205918e, 32'hc17412c2} /* (15, 13, 4) {real, imag} */,
  {32'h41bd3d83, 32'hc1708125} /* (15, 13, 3) {real, imag} */,
  {32'h41100c8e, 32'hc200dc5d} /* (15, 13, 2) {real, imag} */,
  {32'hc2203f2e, 32'h42882ec6} /* (15, 13, 1) {real, imag} */,
  {32'hc10b146f, 32'hc1933f07} /* (15, 13, 0) {real, imag} */,
  {32'h41ffeef7, 32'h41a9d639} /* (15, 12, 15) {real, imag} */,
  {32'h411f5105, 32'hc0acc2a1} /* (15, 12, 14) {real, imag} */,
  {32'hc1995427, 32'hc016b050} /* (15, 12, 13) {real, imag} */,
  {32'hc19b0fa6, 32'hc0fb8500} /* (15, 12, 12) {real, imag} */,
  {32'hc06c6196, 32'h40bff698} /* (15, 12, 11) {real, imag} */,
  {32'h41183c35, 32'hc01e6817} /* (15, 12, 10) {real, imag} */,
  {32'hc0fcf496, 32'h405cef28} /* (15, 12, 9) {real, imag} */,
  {32'hbfe6dc98, 32'hc105dbe4} /* (15, 12, 8) {real, imag} */,
  {32'h4134ff3b, 32'h40aeb8f8} /* (15, 12, 7) {real, imag} */,
  {32'hc10e312f, 32'h40f77b66} /* (15, 12, 6) {real, imag} */,
  {32'hc198c5f5, 32'h40cbaa64} /* (15, 12, 5) {real, imag} */,
  {32'hc1cf483e, 32'hc24e5946} /* (15, 12, 4) {real, imag} */,
  {32'h410e03f6, 32'h41ae5bf1} /* (15, 12, 3) {real, imag} */,
  {32'hc18c3743, 32'hc1427d5a} /* (15, 12, 2) {real, imag} */,
  {32'h421da145, 32'hc0e6fec0} /* (15, 12, 1) {real, imag} */,
  {32'hc0a2f81a, 32'h41e8fbfe} /* (15, 12, 0) {real, imag} */,
  {32'h40c6cab3, 32'h41045cd9} /* (15, 11, 15) {real, imag} */,
  {32'hc1bd9cac, 32'hc0e6bd38} /* (15, 11, 14) {real, imag} */,
  {32'hc0ca770c, 32'h4153e173} /* (15, 11, 13) {real, imag} */,
  {32'hc028c110, 32'hc1043e3e} /* (15, 11, 12) {real, imag} */,
  {32'hbfd3d910, 32'hc161ad49} /* (15, 11, 11) {real, imag} */,
  {32'h409dea04, 32'h40d70a52} /* (15, 11, 10) {real, imag} */,
  {32'h40fe0b97, 32'hc10670c4} /* (15, 11, 9) {real, imag} */,
  {32'hc09b6035, 32'hc0c1c838} /* (15, 11, 8) {real, imag} */,
  {32'hc10fa538, 32'hc0964b38} /* (15, 11, 7) {real, imag} */,
  {32'hc0aa0dd0, 32'hbf16d790} /* (15, 11, 6) {real, imag} */,
  {32'h411725cc, 32'hc19b5a1b} /* (15, 11, 5) {real, imag} */,
  {32'h3f1632e0, 32'h40a825dd} /* (15, 11, 4) {real, imag} */,
  {32'hc0a873e8, 32'hbf648c10} /* (15, 11, 3) {real, imag} */,
  {32'h420b5762, 32'h42325717} /* (15, 11, 2) {real, imag} */,
  {32'hc19a74c3, 32'hbff91268} /* (15, 11, 1) {real, imag} */,
  {32'hc1201ffe, 32'hc24aed77} /* (15, 11, 0) {real, imag} */,
  {32'hc1a4e2f4, 32'hc0ddb6fc} /* (15, 10, 15) {real, imag} */,
  {32'hc160480e, 32'h3ffe1518} /* (15, 10, 14) {real, imag} */,
  {32'hc1cb6236, 32'h40e6f712} /* (15, 10, 13) {real, imag} */,
  {32'h41fd7889, 32'hc05e7ffc} /* (15, 10, 12) {real, imag} */,
  {32'h4179686c, 32'h3e307840} /* (15, 10, 11) {real, imag} */,
  {32'hbf98df76, 32'hbfd3dc08} /* (15, 10, 10) {real, imag} */,
  {32'hbf7cbfb8, 32'hc0a4a02c} /* (15, 10, 9) {real, imag} */,
  {32'h404b0720, 32'h40e2dfbf} /* (15, 10, 8) {real, imag} */,
  {32'h40a33b93, 32'h408b50a8} /* (15, 10, 7) {real, imag} */,
  {32'h3fba8306, 32'hc1432762} /* (15, 10, 6) {real, imag} */,
  {32'hbfbe3844, 32'h4108802f} /* (15, 10, 5) {real, imag} */,
  {32'hc0303038, 32'h414020ce} /* (15, 10, 4) {real, imag} */,
  {32'hbfb2c140, 32'h413dfc95} /* (15, 10, 3) {real, imag} */,
  {32'hc133c734, 32'hc11edcac} /* (15, 10, 2) {real, imag} */,
  {32'h40321310, 32'h40dd8b94} /* (15, 10, 1) {real, imag} */,
  {32'h419a7d0e, 32'hbfc9fb94} /* (15, 10, 0) {real, imag} */,
  {32'hbfec3326, 32'h417bd892} /* (15, 9, 15) {real, imag} */,
  {32'hc0c15234, 32'h3f78b914} /* (15, 9, 14) {real, imag} */,
  {32'h4004300a, 32'hc0c493b2} /* (15, 9, 13) {real, imag} */,
  {32'hc0efe391, 32'h402737ed} /* (15, 9, 12) {real, imag} */,
  {32'hc02926cd, 32'h40073867} /* (15, 9, 11) {real, imag} */,
  {32'hc1105a34, 32'h4037fc9d} /* (15, 9, 10) {real, imag} */,
  {32'h40167188, 32'h3fbbc778} /* (15, 9, 9) {real, imag} */,
  {32'hbe2a4400, 32'hbffbc8ae} /* (15, 9, 8) {real, imag} */,
  {32'hc10214ca, 32'hbf777740} /* (15, 9, 7) {real, imag} */,
  {32'h40040a4e, 32'hbfc61606} /* (15, 9, 6) {real, imag} */,
  {32'h3fe5331e, 32'hbee7b178} /* (15, 9, 5) {real, imag} */,
  {32'h419d0e88, 32'hc08397d4} /* (15, 9, 4) {real, imag} */,
  {32'h40434cf6, 32'hc0677f7c} /* (15, 9, 3) {real, imag} */,
  {32'hc017d7cd, 32'h40b80b46} /* (15, 9, 2) {real, imag} */,
  {32'h40710e45, 32'hbfb2e834} /* (15, 9, 1) {real, imag} */,
  {32'h412746ab, 32'hc06d51eb} /* (15, 9, 0) {real, imag} */,
  {32'hc12b8980, 32'h3f788f60} /* (15, 8, 15) {real, imag} */,
  {32'hc109b2ff, 32'hc104a25c} /* (15, 8, 14) {real, imag} */,
  {32'h40d21f16, 32'h40cae288} /* (15, 8, 13) {real, imag} */,
  {32'hc1170d1b, 32'hc0e3db31} /* (15, 8, 12) {real, imag} */,
  {32'h3fdd5e20, 32'hc07e0ecb} /* (15, 8, 11) {real, imag} */,
  {32'hc1000f21, 32'h403be0bc} /* (15, 8, 10) {real, imag} */,
  {32'h40899c52, 32'h40554f2f} /* (15, 8, 9) {real, imag} */,
  {32'h40152fe4, 32'h4055db4a} /* (15, 8, 8) {real, imag} */,
  {32'hbea196ec, 32'hc05a63b7} /* (15, 8, 7) {real, imag} */,
  {32'hc02d646f, 32'h3e98e984} /* (15, 8, 6) {real, imag} */,
  {32'h3fb8b778, 32'hc10ee2c5} /* (15, 8, 5) {real, imag} */,
  {32'hc0d67a0b, 32'h4070da36} /* (15, 8, 4) {real, imag} */,
  {32'hc02772b3, 32'h4183c2e8} /* (15, 8, 3) {real, imag} */,
  {32'hc0986560, 32'hc0eb4342} /* (15, 8, 2) {real, imag} */,
  {32'h40b7e93f, 32'h4113f22b} /* (15, 8, 1) {real, imag} */,
  {32'hc0ec8caa, 32'h40135892} /* (15, 8, 0) {real, imag} */,
  {32'h412a184a, 32'hc1516b06} /* (15, 7, 15) {real, imag} */,
  {32'h413907c9, 32'h414fe88d} /* (15, 7, 14) {real, imag} */,
  {32'hc037938e, 32'hc0b217f8} /* (15, 7, 13) {real, imag} */,
  {32'hc088ff92, 32'h41a09f62} /* (15, 7, 12) {real, imag} */,
  {32'hc0951dc1, 32'h40f33ec7} /* (15, 7, 11) {real, imag} */,
  {32'h40b0ef99, 32'h4084df52} /* (15, 7, 10) {real, imag} */,
  {32'hbf2ce6d3, 32'hbedf3240} /* (15, 7, 9) {real, imag} */,
  {32'h401a46b0, 32'hbff4a38c} /* (15, 7, 8) {real, imag} */,
  {32'h3e74f58c, 32'h40ccdacc} /* (15, 7, 7) {real, imag} */,
  {32'hbff789b5, 32'h404c19ac} /* (15, 7, 6) {real, imag} */,
  {32'h409be5a9, 32'hc0f7c011} /* (15, 7, 5) {real, imag} */,
  {32'h405754bf, 32'h40149158} /* (15, 7, 4) {real, imag} */,
  {32'hc02ff60e, 32'hc183d6c6} /* (15, 7, 3) {real, imag} */,
  {32'hc104d88b, 32'h40cc379a} /* (15, 7, 2) {real, imag} */,
  {32'h40fec014, 32'hc0ebe77b} /* (15, 7, 1) {real, imag} */,
  {32'h415b7c56, 32'h4109093e} /* (15, 7, 0) {real, imag} */,
  {32'h417eda64, 32'h41d22131} /* (15, 6, 15) {real, imag} */,
  {32'hbfd9be24, 32'h410fcf98} /* (15, 6, 14) {real, imag} */,
  {32'hbf544838, 32'h3fed7520} /* (15, 6, 13) {real, imag} */,
  {32'h4186e88c, 32'hc02da328} /* (15, 6, 12) {real, imag} */,
  {32'hc0c225e7, 32'hbf8e408c} /* (15, 6, 11) {real, imag} */,
  {32'hc13f6ccf, 32'h413100b2} /* (15, 6, 10) {real, imag} */,
  {32'hc0aced1a, 32'hc0c804ef} /* (15, 6, 9) {real, imag} */,
  {32'h40b29870, 32'h40024ac0} /* (15, 6, 8) {real, imag} */,
  {32'h400a873c, 32'h408ce803} /* (15, 6, 7) {real, imag} */,
  {32'h40985e22, 32'hc0f83755} /* (15, 6, 6) {real, imag} */,
  {32'hbfbbc674, 32'hc17b718e} /* (15, 6, 5) {real, imag} */,
  {32'hc1802ff4, 32'h4100fd66} /* (15, 6, 4) {real, imag} */,
  {32'hc0d29ba5, 32'h41c311a8} /* (15, 6, 3) {real, imag} */,
  {32'hc134e73a, 32'h4022e24b} /* (15, 6, 2) {real, imag} */,
  {32'h41af3d6a, 32'h41625c1e} /* (15, 6, 1) {real, imag} */,
  {32'h413a0220, 32'hbc49f800} /* (15, 6, 0) {real, imag} */,
  {32'h41cd3991, 32'h416aeb62} /* (15, 5, 15) {real, imag} */,
  {32'hc037e33e, 32'hc1a7ce35} /* (15, 5, 14) {real, imag} */,
  {32'h42211f65, 32'hc19f1e5a} /* (15, 5, 13) {real, imag} */,
  {32'hbf1843a4, 32'hc18b1fa6} /* (15, 5, 12) {real, imag} */,
  {32'h414b36d8, 32'hc03998e8} /* (15, 5, 11) {real, imag} */,
  {32'h40640f58, 32'hc0ff6309} /* (15, 5, 10) {real, imag} */,
  {32'h3fa3bf08, 32'h41115ebd} /* (15, 5, 9) {real, imag} */,
  {32'h402e64e8, 32'hc05eb708} /* (15, 5, 8) {real, imag} */,
  {32'h40ded75c, 32'hc0fea416} /* (15, 5, 7) {real, imag} */,
  {32'hc10b94f1, 32'hc12762d8} /* (15, 5, 6) {real, imag} */,
  {32'h40e763f1, 32'h41610fc0} /* (15, 5, 5) {real, imag} */,
  {32'h40c2d41e, 32'h3f310510} /* (15, 5, 4) {real, imag} */,
  {32'h416d716c, 32'h41031dcb} /* (15, 5, 3) {real, imag} */,
  {32'hc1547268, 32'hc110a312} /* (15, 5, 2) {real, imag} */,
  {32'h410a863e, 32'h41b0cc1b} /* (15, 5, 1) {real, imag} */,
  {32'hc191af2d, 32'hbf931c60} /* (15, 5, 0) {real, imag} */,
  {32'h412501f4, 32'h418a4176} /* (15, 4, 15) {real, imag} */,
  {32'h40bfade4, 32'hbf6986c0} /* (15, 4, 14) {real, imag} */,
  {32'h4096f502, 32'h40d35928} /* (15, 4, 13) {real, imag} */,
  {32'hc1226445, 32'h40038c26} /* (15, 4, 12) {real, imag} */,
  {32'hc13611d5, 32'hc1277387} /* (15, 4, 11) {real, imag} */,
  {32'h40e6ce56, 32'hc09fabf3} /* (15, 4, 10) {real, imag} */,
  {32'hc07c05b8, 32'h418a95e8} /* (15, 4, 9) {real, imag} */,
  {32'h401e2402, 32'hc0ad8c90} /* (15, 4, 8) {real, imag} */,
  {32'hc190be6e, 32'h40a368b6} /* (15, 4, 7) {real, imag} */,
  {32'hc00e4504, 32'h3f98de54} /* (15, 4, 6) {real, imag} */,
  {32'hbf893e58, 32'h41ba3e68} /* (15, 4, 5) {real, imag} */,
  {32'h41833910, 32'hc0e40467} /* (15, 4, 4) {real, imag} */,
  {32'hc13095b5, 32'hc220d047} /* (15, 4, 3) {real, imag} */,
  {32'hc25df15c, 32'hc1f797b0} /* (15, 4, 2) {real, imag} */,
  {32'h3f2377a0, 32'hc2a1c804} /* (15, 4, 1) {real, imag} */,
  {32'hc0994c85, 32'h42287cd6} /* (15, 4, 0) {real, imag} */,
  {32'h42216891, 32'hc0e01888} /* (15, 3, 15) {real, imag} */,
  {32'hc1a6fb5d, 32'hc23b09ce} /* (15, 3, 14) {real, imag} */,
  {32'hc165c1b2, 32'h426b8634} /* (15, 3, 13) {real, imag} */,
  {32'h416ced70, 32'hc12a200b} /* (15, 3, 12) {real, imag} */,
  {32'hc15b9b3c, 32'hc0e0b06b} /* (15, 3, 11) {real, imag} */,
  {32'h40cd8f0e, 32'h3f985520} /* (15, 3, 10) {real, imag} */,
  {32'h3f5c9598, 32'hc170746f} /* (15, 3, 9) {real, imag} */,
  {32'hc0d26726, 32'h418b343e} /* (15, 3, 8) {real, imag} */,
  {32'hc111bd5e, 32'hc1e84cdc} /* (15, 3, 7) {real, imag} */,
  {32'hbfac3850, 32'hc0ff2438} /* (15, 3, 6) {real, imag} */,
  {32'h40d1e588, 32'h41a5300f} /* (15, 3, 5) {real, imag} */,
  {32'hc205602e, 32'hc109bd05} /* (15, 3, 4) {real, imag} */,
  {32'hc13f527e, 32'hc2524ec8} /* (15, 3, 3) {real, imag} */,
  {32'hbf3b9260, 32'h41e76a14} /* (15, 3, 2) {real, imag} */,
  {32'h4204f4e7, 32'hc104f22e} /* (15, 3, 1) {real, imag} */,
  {32'hc1dfc068, 32'hc2357727} /* (15, 3, 0) {real, imag} */,
  {32'hc2bc284e, 32'h417e6fae} /* (15, 2, 15) {real, imag} */,
  {32'hc273f7b2, 32'h3e173200} /* (15, 2, 14) {real, imag} */,
  {32'h4219384e, 32'hc2384dbf} /* (15, 2, 13) {real, imag} */,
  {32'hc170eea1, 32'h41b5d092} /* (15, 2, 12) {real, imag} */,
  {32'hc16bc5ec, 32'hc116b4b0} /* (15, 2, 11) {real, imag} */,
  {32'hc1560f3e, 32'hc0e96586} /* (15, 2, 10) {real, imag} */,
  {32'h41d64b23, 32'hc1a83600} /* (15, 2, 9) {real, imag} */,
  {32'hc10c60d4, 32'hc04f3490} /* (15, 2, 8) {real, imag} */,
  {32'h41ec9c57, 32'h40a77af8} /* (15, 2, 7) {real, imag} */,
  {32'h40e2500c, 32'hc1acd13e} /* (15, 2, 6) {real, imag} */,
  {32'h40d11c83, 32'h41d90acc} /* (15, 2, 5) {real, imag} */,
  {32'hc1f70410, 32'hc138c824} /* (15, 2, 4) {real, imag} */,
  {32'hc15e5f76, 32'h41aa77da} /* (15, 2, 3) {real, imag} */,
  {32'hc22dff6c, 32'h4289d3a4} /* (15, 2, 2) {real, imag} */,
  {32'h42633134, 32'hc216e38c} /* (15, 2, 1) {real, imag} */,
  {32'h416d9004, 32'h422679af} /* (15, 2, 0) {real, imag} */,
  {32'hc18fa64e, 32'hc231dcf0} /* (15, 1, 15) {real, imag} */,
  {32'h424405ae, 32'hc2254000} /* (15, 1, 14) {real, imag} */,
  {32'hc1a113f6, 32'h41a43662} /* (15, 1, 13) {real, imag} */,
  {32'hc15c45d8, 32'h419f5caa} /* (15, 1, 12) {real, imag} */,
  {32'hc144f844, 32'hc19f8692} /* (15, 1, 11) {real, imag} */,
  {32'hc1528a7d, 32'h419c7cc5} /* (15, 1, 10) {real, imag} */,
  {32'h412cce0d, 32'hc07e2ce0} /* (15, 1, 9) {real, imag} */,
  {32'hc15d76f1, 32'h40b203e1} /* (15, 1, 8) {real, imag} */,
  {32'hbf003b50, 32'h41bfc5cb} /* (15, 1, 7) {real, imag} */,
  {32'h40fb1a32, 32'h41148c84} /* (15, 1, 6) {real, imag} */,
  {32'hc2177989, 32'hc1f4606a} /* (15, 1, 5) {real, imag} */,
  {32'hbf06f360, 32'hc19579aa} /* (15, 1, 4) {real, imag} */,
  {32'h41c66d2a, 32'h4116ddf1} /* (15, 1, 3) {real, imag} */,
  {32'hc0c02a5c, 32'hc218d838} /* (15, 1, 2) {real, imag} */,
  {32'hc10e3a29, 32'h411c7dc0} /* (15, 1, 1) {real, imag} */,
  {32'hc1a41ce8, 32'hc18c2583} /* (15, 1, 0) {real, imag} */,
  {32'h40f48020, 32'hc2a95903} /* (15, 0, 15) {real, imag} */,
  {32'h41f6d154, 32'h423fd0fb} /* (15, 0, 14) {real, imag} */,
  {32'hbf0b3660, 32'h42819c9d} /* (15, 0, 13) {real, imag} */,
  {32'hc141ec98, 32'hc1db4057} /* (15, 0, 12) {real, imag} */,
  {32'h41f888d5, 32'h416889a8} /* (15, 0, 11) {real, imag} */,
  {32'h41c7b1c2, 32'h40eba6a0} /* (15, 0, 10) {real, imag} */,
  {32'hc1c3c578, 32'h3fc17ad0} /* (15, 0, 9) {real, imag} */,
  {32'h4187f286, 32'h40843134} /* (15, 0, 8) {real, imag} */,
  {32'hc0d03b18, 32'hc1d84d47} /* (15, 0, 7) {real, imag} */,
  {32'hc1386e0c, 32'h425b90c4} /* (15, 0, 6) {real, imag} */,
  {32'h4135d946, 32'hc1632ee4} /* (15, 0, 5) {real, imag} */,
  {32'h42970c3f, 32'h41e51565} /* (15, 0, 4) {real, imag} */,
  {32'hc113e068, 32'h40d7266c} /* (15, 0, 3) {real, imag} */,
  {32'hc16fde50, 32'hc2758245} /* (15, 0, 2) {real, imag} */,
  {32'h41e38c9a, 32'h422a9b68} /* (15, 0, 1) {real, imag} */,
  {32'hc19fb956, 32'hc23e8d84} /* (15, 0, 0) {real, imag} */,
  {32'hc2b5b5de, 32'hc21d1354} /* (14, 15, 15) {real, imag} */,
  {32'h3dd6f800, 32'hc2500813} /* (14, 15, 14) {real, imag} */,
  {32'hc0895230, 32'h42248660} /* (14, 15, 13) {real, imag} */,
  {32'h4116018e, 32'h41a717a4} /* (14, 15, 12) {real, imag} */,
  {32'hc21ba7b0, 32'hc11469a2} /* (14, 15, 11) {real, imag} */,
  {32'hc0e7f490, 32'h3f1c8460} /* (14, 15, 10) {real, imag} */,
  {32'h4182e992, 32'hc085d39a} /* (14, 15, 9) {real, imag} */,
  {32'h3f0cd660, 32'h3f3552d8} /* (14, 15, 8) {real, imag} */,
  {32'h41029c28, 32'hc162440d} /* (14, 15, 7) {real, imag} */,
  {32'hc1c1012c, 32'hc093df00} /* (14, 15, 6) {real, imag} */,
  {32'h41289d04, 32'h407600c8} /* (14, 15, 5) {real, imag} */,
  {32'hc23bf07e, 32'hc1336e24} /* (14, 15, 4) {real, imag} */,
  {32'h4216ee1f, 32'h42845f5c} /* (14, 15, 3) {real, imag} */,
  {32'h41c40f08, 32'hc11c3a9c} /* (14, 15, 2) {real, imag} */,
  {32'hc0b93320, 32'h410114b7} /* (14, 15, 1) {real, imag} */,
  {32'h42179f5a, 32'hc0e214cd} /* (14, 15, 0) {real, imag} */,
  {32'hc0a21bcc, 32'hc209a987} /* (14, 14, 15) {real, imag} */,
  {32'hc1c08a3f, 32'hc1cb093c} /* (14, 14, 14) {real, imag} */,
  {32'h420c15b8, 32'hc1704b1e} /* (14, 14, 13) {real, imag} */,
  {32'h4262c19f, 32'hc22d035c} /* (14, 14, 12) {real, imag} */,
  {32'hc15eb149, 32'hc10a1eb2} /* (14, 14, 11) {real, imag} */,
  {32'hc1c91756, 32'hc18642bd} /* (14, 14, 10) {real, imag} */,
  {32'h3fa3edb8, 32'h41f575f6} /* (14, 14, 9) {real, imag} */,
  {32'hc10e4758, 32'hc0049bfc} /* (14, 14, 8) {real, imag} */,
  {32'hc0df6db2, 32'hc10dfe0c} /* (14, 14, 7) {real, imag} */,
  {32'h41390208, 32'h3e9843c0} /* (14, 14, 6) {real, imag} */,
  {32'h41297313, 32'h42066b28} /* (14, 14, 5) {real, imag} */,
  {32'h3ff4c6a0, 32'hc113600a} /* (14, 14, 4) {real, imag} */,
  {32'hc22d01b0, 32'hc23b58e6} /* (14, 14, 3) {real, imag} */,
  {32'hc28e554e, 32'h4237a0de} /* (14, 14, 2) {real, imag} */,
  {32'h41f54117, 32'h414956e4} /* (14, 14, 1) {real, imag} */,
  {32'h41508b10, 32'h412fab0b} /* (14, 14, 0) {real, imag} */,
  {32'h418a9696, 32'h4080c2a4} /* (14, 13, 15) {real, imag} */,
  {32'hbfe222b0, 32'h405bb78e} /* (14, 13, 14) {real, imag} */,
  {32'hc21b8a4d, 32'h40fb9d10} /* (14, 13, 13) {real, imag} */,
  {32'hc1e4ded3, 32'h41aab835} /* (14, 13, 12) {real, imag} */,
  {32'h40ac83ee, 32'h4187a796} /* (14, 13, 11) {real, imag} */,
  {32'hc08b52d8, 32'hc163df4e} /* (14, 13, 10) {real, imag} */,
  {32'hc0f915b5, 32'hc08629ff} /* (14, 13, 9) {real, imag} */,
  {32'hc0cc1618, 32'h40b74daf} /* (14, 13, 8) {real, imag} */,
  {32'hc13fcf34, 32'h4005ce92} /* (14, 13, 7) {real, imag} */,
  {32'hc1acde8c, 32'hc16daa8e} /* (14, 13, 6) {real, imag} */,
  {32'hc12ff221, 32'h413340bc} /* (14, 13, 5) {real, imag} */,
  {32'hc1be1bcb, 32'h41467be6} /* (14, 13, 4) {real, imag} */,
  {32'hc0cf6568, 32'h423352fa} /* (14, 13, 3) {real, imag} */,
  {32'h422665dc, 32'hc16bbf58} /* (14, 13, 2) {real, imag} */,
  {32'h41912412, 32'h41d645c7} /* (14, 13, 1) {real, imag} */,
  {32'hc22e979a, 32'h3f016a68} /* (14, 13, 0) {real, imag} */,
  {32'hc20645f7, 32'h40f102a7} /* (14, 12, 15) {real, imag} */,
  {32'hc21e8733, 32'h40a95f0e} /* (14, 12, 14) {real, imag} */,
  {32'hc2148acc, 32'h41e11630} /* (14, 12, 13) {real, imag} */,
  {32'h40ba0d58, 32'h4080e4aa} /* (14, 12, 12) {real, imag} */,
  {32'h4195237d, 32'hc10b8856} /* (14, 12, 11) {real, imag} */,
  {32'hc15c5c98, 32'hbf175330} /* (14, 12, 10) {real, imag} */,
  {32'h4142ba4e, 32'hc0a9b8f1} /* (14, 12, 9) {real, imag} */,
  {32'h3e8347c0, 32'hc099793f} /* (14, 12, 8) {real, imag} */,
  {32'h4113508e, 32'h40eb31ff} /* (14, 12, 7) {real, imag} */,
  {32'h40f779c0, 32'h417714b1} /* (14, 12, 6) {real, imag} */,
  {32'h40c7e6e4, 32'h4112a2ba} /* (14, 12, 5) {real, imag} */,
  {32'hc0902360, 32'h41a035f8} /* (14, 12, 4) {real, imag} */,
  {32'hc022fc50, 32'h4135df54} /* (14, 12, 3) {real, imag} */,
  {32'h40d5fe38, 32'hc1f5d21e} /* (14, 12, 2) {real, imag} */,
  {32'h4204d4ed, 32'hc081b4a9} /* (14, 12, 1) {real, imag} */,
  {32'hc20f8e40, 32'h411eb2dc} /* (14, 12, 0) {real, imag} */,
  {32'hc11d349b, 32'h41d14c36} /* (14, 11, 15) {real, imag} */,
  {32'h41d9534b, 32'hbf711f70} /* (14, 11, 14) {real, imag} */,
  {32'hbf77e068, 32'hc1bf78a0} /* (14, 11, 13) {real, imag} */,
  {32'h416500fa, 32'h41a66fb6} /* (14, 11, 12) {real, imag} */,
  {32'h40c1b4c2, 32'h4025c44c} /* (14, 11, 11) {real, imag} */,
  {32'hc18ac8c8, 32'h3fde7b68} /* (14, 11, 10) {real, imag} */,
  {32'hc05d3a92, 32'hbffb2478} /* (14, 11, 9) {real, imag} */,
  {32'h3fd92374, 32'hbf31b5a0} /* (14, 11, 8) {real, imag} */,
  {32'h40296416, 32'h411316b5} /* (14, 11, 7) {real, imag} */,
  {32'hc158c333, 32'hc1cd2b78} /* (14, 11, 6) {real, imag} */,
  {32'hc0208f87, 32'h4190f0f2} /* (14, 11, 5) {real, imag} */,
  {32'hc089d339, 32'h40526254} /* (14, 11, 4) {real, imag} */,
  {32'h412974b6, 32'hc1eaca14} /* (14, 11, 3) {real, imag} */,
  {32'h41172dfa, 32'hc0f389fa} /* (14, 11, 2) {real, imag} */,
  {32'hc1783311, 32'h405b0f3c} /* (14, 11, 1) {real, imag} */,
  {32'hc15623f2, 32'hc1cdc296} /* (14, 11, 0) {real, imag} */,
  {32'h3f1406a4, 32'hc1ba8e60} /* (14, 10, 15) {real, imag} */,
  {32'h40f24f91, 32'h3fd043c0} /* (14, 10, 14) {real, imag} */,
  {32'h416242aa, 32'h404b5140} /* (14, 10, 13) {real, imag} */,
  {32'hc1421f0e, 32'h4078e0ce} /* (14, 10, 12) {real, imag} */,
  {32'hc175298d, 32'h3fd40c14} /* (14, 10, 11) {real, imag} */,
  {32'hc09ee415, 32'hc17d3258} /* (14, 10, 10) {real, imag} */,
  {32'h3fd58bda, 32'h405d3fb7} /* (14, 10, 9) {real, imag} */,
  {32'h4081f344, 32'h3f8afadc} /* (14, 10, 8) {real, imag} */,
  {32'h3fec1886, 32'hc1294570} /* (14, 10, 7) {real, imag} */,
  {32'h40f823ef, 32'hc0df1864} /* (14, 10, 6) {real, imag} */,
  {32'hc1958dd2, 32'h3f3d5ec8} /* (14, 10, 5) {real, imag} */,
  {32'h4150ea0a, 32'hbe523b20} /* (14, 10, 4) {real, imag} */,
  {32'hc028a172, 32'hc03c8670} /* (14, 10, 3) {real, imag} */,
  {32'hbf13d898, 32'hc04c0a68} /* (14, 10, 2) {real, imag} */,
  {32'hc0b8cb28, 32'h41c3c440} /* (14, 10, 1) {real, imag} */,
  {32'hc0ca4958, 32'hc0f86df9} /* (14, 10, 0) {real, imag} */,
  {32'h40d46322, 32'hbf67a880} /* (14, 9, 15) {real, imag} */,
  {32'hc1a6cfa8, 32'hbef0f740} /* (14, 9, 14) {real, imag} */,
  {32'h3fdde53a, 32'hc14c68d6} /* (14, 9, 13) {real, imag} */,
  {32'h3fa3b94c, 32'hc0231eb8} /* (14, 9, 12) {real, imag} */,
  {32'h40e95275, 32'h3fbb07f8} /* (14, 9, 11) {real, imag} */,
  {32'h41585288, 32'hc01a78fc} /* (14, 9, 10) {real, imag} */,
  {32'hbf26e9c2, 32'h408f1b92} /* (14, 9, 9) {real, imag} */,
  {32'hbf1da458, 32'hbe127f50} /* (14, 9, 8) {real, imag} */,
  {32'h400e9404, 32'h4058e4ac} /* (14, 9, 7) {real, imag} */,
  {32'h40b13e3c, 32'h40df89b6} /* (14, 9, 6) {real, imag} */,
  {32'h40d3b02d, 32'hc011e9c0} /* (14, 9, 5) {real, imag} */,
  {32'hc100ec3a, 32'hc00f0418} /* (14, 9, 4) {real, imag} */,
  {32'h40b68ff4, 32'hc0db02fd} /* (14, 9, 3) {real, imag} */,
  {32'hc0875264, 32'h40e686b8} /* (14, 9, 2) {real, imag} */,
  {32'hc0d45fa8, 32'h40d38c9c} /* (14, 9, 1) {real, imag} */,
  {32'h4102d5ba, 32'h402fab11} /* (14, 9, 0) {real, imag} */,
  {32'h4180c725, 32'hbfd70f10} /* (14, 8, 15) {real, imag} */,
  {32'h409c996f, 32'h408ddc50} /* (14, 8, 14) {real, imag} */,
  {32'hc130f8f0, 32'h41037a49} /* (14, 8, 13) {real, imag} */,
  {32'hc0d41594, 32'hc166de5c} /* (14, 8, 12) {real, imag} */,
  {32'h4104e9ea, 32'hc084fea1} /* (14, 8, 11) {real, imag} */,
  {32'h405356bc, 32'hbfb69fd4} /* (14, 8, 10) {real, imag} */,
  {32'h3e05f430, 32'hbfb9c378} /* (14, 8, 9) {real, imag} */,
  {32'hbf3030ba, 32'h4000201e} /* (14, 8, 8) {real, imag} */,
  {32'h400fb2ef, 32'hc00f0fea} /* (14, 8, 7) {real, imag} */,
  {32'h3f72d420, 32'h3f3aae88} /* (14, 8, 6) {real, imag} */,
  {32'hc0c31c29, 32'hbfd78398} /* (14, 8, 5) {real, imag} */,
  {32'hc0ed7ed0, 32'hc0f4a250} /* (14, 8, 4) {real, imag} */,
  {32'hc1375e44, 32'h40742313} /* (14, 8, 3) {real, imag} */,
  {32'hc18b3c2c, 32'hc1846da2} /* (14, 8, 2) {real, imag} */,
  {32'hc11cf7d6, 32'h4026767a} /* (14, 8, 1) {real, imag} */,
  {32'h3f0f5002, 32'hc15c57cc} /* (14, 8, 0) {real, imag} */,
  {32'hc10520e2, 32'h3f39f2ba} /* (14, 7, 15) {real, imag} */,
  {32'hc01d46ec, 32'hc1196fa7} /* (14, 7, 14) {real, imag} */,
  {32'h4181ef6a, 32'hc07cf224} /* (14, 7, 13) {real, imag} */,
  {32'hc13cf89a, 32'hc0073dc6} /* (14, 7, 12) {real, imag} */,
  {32'hc129a284, 32'h3e2e90c0} /* (14, 7, 11) {real, imag} */,
  {32'hc0b28cdd, 32'hbf626d32} /* (14, 7, 10) {real, imag} */,
  {32'hbfa4b65b, 32'h3f25b396} /* (14, 7, 9) {real, imag} */,
  {32'h4083c091, 32'h402068ec} /* (14, 7, 8) {real, imag} */,
  {32'h3e466eb8, 32'h3e8a159d} /* (14, 7, 7) {real, imag} */,
  {32'hc0c772bd, 32'h4044d5ec} /* (14, 7, 6) {real, imag} */,
  {32'h3f5da9e8, 32'h4110cae3} /* (14, 7, 5) {real, imag} */,
  {32'h40bb633b, 32'h41007b94} /* (14, 7, 4) {real, imag} */,
  {32'h3fc3af9c, 32'h41243443} /* (14, 7, 3) {real, imag} */,
  {32'hbdd4f3f0, 32'h40c276fa} /* (14, 7, 2) {real, imag} */,
  {32'hc0d99dd5, 32'h3f6b6da2} /* (14, 7, 1) {real, imag} */,
  {32'h40d8a925, 32'h40b61f80} /* (14, 7, 0) {real, imag} */,
  {32'h41654eb5, 32'hbf9239e0} /* (14, 6, 15) {real, imag} */,
  {32'hc0d4571c, 32'h3f7f2df4} /* (14, 6, 14) {real, imag} */,
  {32'h4177af2e, 32'hc0a97d4a} /* (14, 6, 13) {real, imag} */,
  {32'hc12df440, 32'h412cb880} /* (14, 6, 12) {real, imag} */,
  {32'h40d9b746, 32'hc09424cc} /* (14, 6, 11) {real, imag} */,
  {32'h40a1d87d, 32'hbf82b83e} /* (14, 6, 10) {real, imag} */,
  {32'hbfb13d14, 32'h407e6d22} /* (14, 6, 9) {real, imag} */,
  {32'hc02a4e86, 32'h40228e52} /* (14, 6, 8) {real, imag} */,
  {32'hc03e041e, 32'h3fc330b1} /* (14, 6, 7) {real, imag} */,
  {32'hc0a6b21f, 32'hbebe276e} /* (14, 6, 6) {real, imag} */,
  {32'hc0030ec8, 32'h403f37c9} /* (14, 6, 5) {real, imag} */,
  {32'h404200d9, 32'hc17f8d38} /* (14, 6, 4) {real, imag} */,
  {32'hc10e48fe, 32'h3fb8954a} /* (14, 6, 3) {real, imag} */,
  {32'hc1ac8b91, 32'h406ee2a3} /* (14, 6, 2) {real, imag} */,
  {32'hc0e8ee06, 32'hc12e18ba} /* (14, 6, 1) {real, imag} */,
  {32'h414bc9d8, 32'hc0c185db} /* (14, 6, 0) {real, imag} */,
  {32'hbfd1bd78, 32'h41175bd7} /* (14, 5, 15) {real, imag} */,
  {32'hc1c4f90a, 32'hc11e2e06} /* (14, 5, 14) {real, imag} */,
  {32'hc0340200, 32'h41292e51} /* (14, 5, 13) {real, imag} */,
  {32'h4154740a, 32'h40ed4b0a} /* (14, 5, 12) {real, imag} */,
  {32'hc0b5530e, 32'hc007e77c} /* (14, 5, 11) {real, imag} */,
  {32'h4134c268, 32'hc00cb856} /* (14, 5, 10) {real, imag} */,
  {32'h40fddca6, 32'hc120cb93} /* (14, 5, 9) {real, imag} */,
  {32'h3ebcb670, 32'h4056ea0c} /* (14, 5, 8) {real, imag} */,
  {32'h409cd29a, 32'h40d62976} /* (14, 5, 7) {real, imag} */,
  {32'h4120dad8, 32'hc1414f38} /* (14, 5, 6) {real, imag} */,
  {32'hc0d5cb70, 32'hc1132347} /* (14, 5, 5) {real, imag} */,
  {32'hc11e5022, 32'h410741fc} /* (14, 5, 4) {real, imag} */,
  {32'hc04cf404, 32'hc14eecb3} /* (14, 5, 3) {real, imag} */,
  {32'h40ab9aa8, 32'h41a44720} /* (14, 5, 2) {real, imag} */,
  {32'h41e4b06a, 32'h421cf754} /* (14, 5, 1) {real, imag} */,
  {32'h4140625e, 32'hc1cddfc4} /* (14, 5, 0) {real, imag} */,
  {32'h4183ab64, 32'h42406d4a} /* (14, 4, 15) {real, imag} */,
  {32'hc0285aee, 32'h412ea678} /* (14, 4, 14) {real, imag} */,
  {32'h416e0e12, 32'h41ab5713} /* (14, 4, 13) {real, imag} */,
  {32'h41cca24d, 32'hc2316056} /* (14, 4, 12) {real, imag} */,
  {32'hbfb73a60, 32'h41c44544} /* (14, 4, 11) {real, imag} */,
  {32'h40e5df4c, 32'h40c75ed3} /* (14, 4, 10) {real, imag} */,
  {32'h40e72a73, 32'h41106a78} /* (14, 4, 9) {real, imag} */,
  {32'hc128eb9c, 32'hc04ab5ca} /* (14, 4, 8) {real, imag} */,
  {32'h3f9e286c, 32'hc04e3060} /* (14, 4, 7) {real, imag} */,
  {32'hc0d23bd2, 32'hc05c446e} /* (14, 4, 6) {real, imag} */,
  {32'h422570a8, 32'h4138bf74} /* (14, 4, 5) {real, imag} */,
  {32'hbfc63f90, 32'h4082c864} /* (14, 4, 4) {real, imag} */,
  {32'h40a82a24, 32'hc28ed2ab} /* (14, 4, 3) {real, imag} */,
  {32'hc10c658a, 32'h41567c88} /* (14, 4, 2) {real, imag} */,
  {32'hc065b022, 32'hc0a73d94} /* (14, 4, 1) {real, imag} */,
  {32'h40d46ab0, 32'hc13ca828} /* (14, 4, 0) {real, imag} */,
  {32'h41843379, 32'hc23130fd} /* (14, 3, 15) {real, imag} */,
  {32'h407df718, 32'hc17d1573} /* (14, 3, 14) {real, imag} */,
  {32'h3fc72570, 32'h41845f42} /* (14, 3, 13) {real, imag} */,
  {32'h40581f10, 32'hc21511ac} /* (14, 3, 12) {real, imag} */,
  {32'h417ab70e, 32'h41754c1d} /* (14, 3, 11) {real, imag} */,
  {32'h40e996d3, 32'h41694e56} /* (14, 3, 10) {real, imag} */,
  {32'h40ce278f, 32'hc136240d} /* (14, 3, 9) {real, imag} */,
  {32'hc0adea24, 32'hbff5ab00} /* (14, 3, 8) {real, imag} */,
  {32'hc155dcf0, 32'hc086f27e} /* (14, 3, 7) {real, imag} */,
  {32'hc0d11f1f, 32'hc09c8578} /* (14, 3, 6) {real, imag} */,
  {32'hc163d1fc, 32'h3f889c78} /* (14, 3, 5) {real, imag} */,
  {32'h42309db0, 32'hc12c76ae} /* (14, 3, 4) {real, imag} */,
  {32'h4225da82, 32'hc0e4da06} /* (14, 3, 3) {real, imag} */,
  {32'h40ae4b52, 32'hc09ea176} /* (14, 3, 2) {real, imag} */,
  {32'hc17d74b6, 32'h3e7daf00} /* (14, 3, 1) {real, imag} */,
  {32'hc0d4e114, 32'h40cd5258} /* (14, 3, 0) {real, imag} */,
  {32'h42380652, 32'h4289f407} /* (14, 2, 15) {real, imag} */,
  {32'h4235ef21, 32'h41d77a00} /* (14, 2, 14) {real, imag} */,
  {32'h40c48ad0, 32'h420bbe34} /* (14, 2, 13) {real, imag} */,
  {32'hc07dffbb, 32'hc202ab60} /* (14, 2, 12) {real, imag} */,
  {32'hc0be98d8, 32'hc0d33af0} /* (14, 2, 11) {real, imag} */,
  {32'h3e8c8640, 32'hc02ee1b8} /* (14, 2, 10) {real, imag} */,
  {32'hc047a8e0, 32'h4072e128} /* (14, 2, 9) {real, imag} */,
  {32'h3e0fde40, 32'h3f90a658} /* (14, 2, 8) {real, imag} */,
  {32'hbfc1d400, 32'hc0cdf774} /* (14, 2, 7) {real, imag} */,
  {32'h40376b30, 32'hc0cf3270} /* (14, 2, 6) {real, imag} */,
  {32'h4165dcd4, 32'hc11fab24} /* (14, 2, 5) {real, imag} */,
  {32'hc0c4b37e, 32'h418676ba} /* (14, 2, 4) {real, imag} */,
  {32'h428156bf, 32'hc131335c} /* (14, 2, 3) {real, imag} */,
  {32'h40a3e5a8, 32'hc20a919a} /* (14, 2, 2) {real, imag} */,
  {32'hc2ee3c8f, 32'hc13b1768} /* (14, 2, 1) {real, imag} */,
  {32'hc18178da, 32'h4120cbef} /* (14, 2, 0) {real, imag} */,
  {32'hc1d1700b, 32'hc19e1e8f} /* (14, 1, 15) {real, imag} */,
  {32'hc13a757e, 32'h41ad7761} /* (14, 1, 14) {real, imag} */,
  {32'hbd563200, 32'h41928b44} /* (14, 1, 13) {real, imag} */,
  {32'h4084d230, 32'hc288d994} /* (14, 1, 12) {real, imag} */,
  {32'hc04b8cc8, 32'hc0ba4967} /* (14, 1, 11) {real, imag} */,
  {32'h3fb669e0, 32'h4122051a} /* (14, 1, 10) {real, imag} */,
  {32'hc0d4a449, 32'hc17fac14} /* (14, 1, 9) {real, imag} */,
  {32'hc0909f30, 32'hbfb8a120} /* (14, 1, 8) {real, imag} */,
  {32'hbb77f800, 32'hc13082d6} /* (14, 1, 7) {real, imag} */,
  {32'hc08d6720, 32'hbed1c3d0} /* (14, 1, 6) {real, imag} */,
  {32'hc01ce18c, 32'hc00f5402} /* (14, 1, 5) {real, imag} */,
  {32'hc18e73f4, 32'hc0626170} /* (14, 1, 4) {real, imag} */,
  {32'h417b116b, 32'h41d7e04a} /* (14, 1, 3) {real, imag} */,
  {32'h428c82b2, 32'h40722588} /* (14, 1, 2) {real, imag} */,
  {32'h3e5b6980, 32'hc2223bfa} /* (14, 1, 1) {real, imag} */,
  {32'hc28fbf47, 32'h40f7aa88} /* (14, 1, 0) {real, imag} */,
  {32'h41c53440, 32'hc11637e8} /* (14, 0, 15) {real, imag} */,
  {32'hbf4462b0, 32'hbddd9f60} /* (14, 0, 14) {real, imag} */,
  {32'hc200a110, 32'h416e33cc} /* (14, 0, 13) {real, imag} */,
  {32'hc014a9e4, 32'h423f50d0} /* (14, 0, 12) {real, imag} */,
  {32'hc229e1ac, 32'h404c54e0} /* (14, 0, 11) {real, imag} */,
  {32'hc0a8bd46, 32'h3fe72888} /* (14, 0, 10) {real, imag} */,
  {32'h3e0f4090, 32'h400291b8} /* (14, 0, 9) {real, imag} */,
  {32'h41a96fdf, 32'hc10e932c} /* (14, 0, 8) {real, imag} */,
  {32'hc02e0ff9, 32'h413d6330} /* (14, 0, 7) {real, imag} */,
  {32'hc09cd18a, 32'hc1c714d2} /* (14, 0, 6) {real, imag} */,
  {32'h41afbebf, 32'h41041c09} /* (14, 0, 5) {real, imag} */,
  {32'hc197dbd8, 32'h40a1b388} /* (14, 0, 4) {real, imag} */,
  {32'h4232c714, 32'h413e5d94} /* (14, 0, 3) {real, imag} */,
  {32'hc1b89084, 32'hc0e77aee} /* (14, 0, 2) {real, imag} */,
  {32'h41059be1, 32'h41528ca6} /* (14, 0, 1) {real, imag} */,
  {32'h422db0f6, 32'h42c19ee2} /* (14, 0, 0) {real, imag} */,
  {32'hc22a0c99, 32'hc2044c5c} /* (13, 15, 15) {real, imag} */,
  {32'h41a5ac94, 32'h41673f47} /* (13, 15, 14) {real, imag} */,
  {32'h4237f9b7, 32'hc204cd18} /* (13, 15, 13) {real, imag} */,
  {32'hc0c750e4, 32'hc0b046ce} /* (13, 15, 12) {real, imag} */,
  {32'h40177234, 32'hc0d8a68a} /* (13, 15, 11) {real, imag} */,
  {32'h414fbc4e, 32'h41d3540c} /* (13, 15, 10) {real, imag} */,
  {32'h3f892850, 32'h406b92ac} /* (13, 15, 9) {real, imag} */,
  {32'hc005aa7c, 32'hc0ff2808} /* (13, 15, 8) {real, imag} */,
  {32'hc1ae5955, 32'h406d959c} /* (13, 15, 7) {real, imag} */,
  {32'hc0921318, 32'hc10a5b2d} /* (13, 15, 6) {real, imag} */,
  {32'hc10b8d8b, 32'hc06de004} /* (13, 15, 5) {real, imag} */,
  {32'h411cdefa, 32'h3dc32180} /* (13, 15, 4) {real, imag} */,
  {32'hc1a2230e, 32'h41c48822} /* (13, 15, 3) {real, imag} */,
  {32'hc2466422, 32'h414bee7b} /* (13, 15, 2) {real, imag} */,
  {32'h419510cc, 32'h419b8792} /* (13, 15, 1) {real, imag} */,
  {32'hc1c2af30, 32'hc21ac383} /* (13, 15, 0) {real, imag} */,
  {32'hc1994746, 32'hbe835800} /* (13, 14, 15) {real, imag} */,
  {32'h420ca311, 32'h4216ea6c} /* (13, 14, 14) {real, imag} */,
  {32'hc127ea23, 32'h4127964d} /* (13, 14, 13) {real, imag} */,
  {32'h41cc8714, 32'hc0cb016f} /* (13, 14, 12) {real, imag} */,
  {32'h418ef824, 32'h407b4c9c} /* (13, 14, 11) {real, imag} */,
  {32'hc0c77bc4, 32'hc04bb6d6} /* (13, 14, 10) {real, imag} */,
  {32'h3fb5fd66, 32'hbf403800} /* (13, 14, 9) {real, imag} */,
  {32'h406f3394, 32'hc07454fe} /* (13, 14, 8) {real, imag} */,
  {32'h3f979666, 32'h3f89fe10} /* (13, 14, 7) {real, imag} */,
  {32'h407f4db8, 32'hc0a966ab} /* (13, 14, 6) {real, imag} */,
  {32'hc103f459, 32'hc1f5620c} /* (13, 14, 5) {real, imag} */,
  {32'h41a21650, 32'h3ef4f7d0} /* (13, 14, 4) {real, imag} */,
  {32'h415e5d39, 32'h421f3039} /* (13, 14, 3) {real, imag} */,
  {32'h42415fcb, 32'hc2271aca} /* (13, 14, 2) {real, imag} */,
  {32'h41f6b1d4, 32'hc271093e} /* (13, 14, 1) {real, imag} */,
  {32'hc20b9ce1, 32'h4135dec6} /* (13, 14, 0) {real, imag} */,
  {32'hc1c5d7ce, 32'h41a11af8} /* (13, 13, 15) {real, imag} */,
  {32'h3ec20aa0, 32'hc1fbddfb} /* (13, 13, 14) {real, imag} */,
  {32'hc180c370, 32'h41009fcb} /* (13, 13, 13) {real, imag} */,
  {32'h40903314, 32'h41c71f22} /* (13, 13, 12) {real, imag} */,
  {32'hc201bf2a, 32'hc102a310} /* (13, 13, 11) {real, imag} */,
  {32'hbf3c5b40, 32'h41b42318} /* (13, 13, 10) {real, imag} */,
  {32'hc1338301, 32'h412a8609} /* (13, 13, 9) {real, imag} */,
  {32'h41159f56, 32'hbeff5470} /* (13, 13, 8) {real, imag} */,
  {32'hbf91afc8, 32'hc022e07c} /* (13, 13, 7) {real, imag} */,
  {32'hc13be8c4, 32'h40d7402a} /* (13, 13, 6) {real, imag} */,
  {32'h411a5c9a, 32'h41abbc04} /* (13, 13, 5) {real, imag} */,
  {32'hbfe0831e, 32'h419ca946} /* (13, 13, 4) {real, imag} */,
  {32'h4189716c, 32'hbf522bcc} /* (13, 13, 3) {real, imag} */,
  {32'h4174851b, 32'h4209a0f7} /* (13, 13, 2) {real, imag} */,
  {32'h4028b214, 32'h401d1ed4} /* (13, 13, 1) {real, imag} */,
  {32'h41c10305, 32'hc1594e96} /* (13, 13, 0) {real, imag} */,
  {32'h42634d01, 32'hc2015035} /* (13, 12, 15) {real, imag} */,
  {32'h3e5c2180, 32'h41746f8c} /* (13, 12, 14) {real, imag} */,
  {32'hc0cc4c12, 32'hc0d731bc} /* (13, 12, 13) {real, imag} */,
  {32'hc1952448, 32'hc0b7a1ac} /* (13, 12, 12) {real, imag} */,
  {32'hc15a9d88, 32'h3ff2f260} /* (13, 12, 11) {real, imag} */,
  {32'h417de4c2, 32'hc0498654} /* (13, 12, 10) {real, imag} */,
  {32'hbff761a8, 32'h40ef0582} /* (13, 12, 9) {real, imag} */,
  {32'h408c58e8, 32'hc0186ef8} /* (13, 12, 8) {real, imag} */,
  {32'hbfb27a78, 32'h40000aa4} /* (13, 12, 7) {real, imag} */,
  {32'h401dfec0, 32'h3ff59801} /* (13, 12, 6) {real, imag} */,
  {32'hbf167140, 32'hc106e53c} /* (13, 12, 5) {real, imag} */,
  {32'hbefea980, 32'h422332b0} /* (13, 12, 4) {real, imag} */,
  {32'hc0ac40be, 32'hc1dfc92f} /* (13, 12, 3) {real, imag} */,
  {32'h41f60936, 32'hc16b1660} /* (13, 12, 2) {real, imag} */,
  {32'h4139dc2c, 32'h3f5e9770} /* (13, 12, 1) {real, imag} */,
  {32'hc1f4f132, 32'h41c8a349} /* (13, 12, 0) {real, imag} */,
  {32'h40b7c010, 32'hc14de370} /* (13, 11, 15) {real, imag} */,
  {32'hc0989c85, 32'hc1074efa} /* (13, 11, 14) {real, imag} */,
  {32'hc0a48bf8, 32'h40ba4c30} /* (13, 11, 13) {real, imag} */,
  {32'hc206c270, 32'hc1bcf7e7} /* (13, 11, 12) {real, imag} */,
  {32'hc07f0f03, 32'h4067b304} /* (13, 11, 11) {real, imag} */,
  {32'h404c3761, 32'hc0c10dfb} /* (13, 11, 10) {real, imag} */,
  {32'hc06e2616, 32'hbec91950} /* (13, 11, 9) {real, imag} */,
  {32'h3f4ffb08, 32'h4023c060} /* (13, 11, 8) {real, imag} */,
  {32'h40e043d7, 32'hc033d08a} /* (13, 11, 7) {real, imag} */,
  {32'hc0b2e9ee, 32'hc0fde09f} /* (13, 11, 6) {real, imag} */,
  {32'hbe5430d0, 32'hc188798e} /* (13, 11, 5) {real, imag} */,
  {32'hbf802140, 32'hc085edb4} /* (13, 11, 4) {real, imag} */,
  {32'hc183ceb6, 32'h4217bb5c} /* (13, 11, 3) {real, imag} */,
  {32'h40564ebb, 32'hc09099a2} /* (13, 11, 2) {real, imag} */,
  {32'h41b4c7c9, 32'h41a32764} /* (13, 11, 1) {real, imag} */,
  {32'hc04c1e2a, 32'h421a2e60} /* (13, 11, 0) {real, imag} */,
  {32'h4098279c, 32'hc1761068} /* (13, 10, 15) {real, imag} */,
  {32'h40bba311, 32'h40ce70da} /* (13, 10, 14) {real, imag} */,
  {32'h3fe53647, 32'h3e8170c8} /* (13, 10, 13) {real, imag} */,
  {32'hc1268486, 32'hc182913a} /* (13, 10, 12) {real, imag} */,
  {32'h40dbfd55, 32'h3edbd1f0} /* (13, 10, 11) {real, imag} */,
  {32'h3f38f02c, 32'h3f9aed2f} /* (13, 10, 10) {real, imag} */,
  {32'h40acb052, 32'hc000aa1e} /* (13, 10, 9) {real, imag} */,
  {32'hc0009e8c, 32'h40899ed8} /* (13, 10, 8) {real, imag} */,
  {32'hbfe81970, 32'hc045eb02} /* (13, 10, 7) {real, imag} */,
  {32'h3f3ae0e0, 32'hc06fa8cc} /* (13, 10, 6) {real, imag} */,
  {32'h41008dbb, 32'h410b472a} /* (13, 10, 5) {real, imag} */,
  {32'hbf858b14, 32'h40a37dc2} /* (13, 10, 4) {real, imag} */,
  {32'hbf65474e, 32'h400fe015} /* (13, 10, 3) {real, imag} */,
  {32'h3f7de5c8, 32'h404cc454} /* (13, 10, 2) {real, imag} */,
  {32'hc1b25cb9, 32'h417714e0} /* (13, 10, 1) {real, imag} */,
  {32'hc1b169ee, 32'h3fa2563f} /* (13, 10, 0) {real, imag} */,
  {32'hc144b3f4, 32'h40dbea0a} /* (13, 9, 15) {real, imag} */,
  {32'h3f1167a0, 32'hc04f9a6f} /* (13, 9, 14) {real, imag} */,
  {32'h40ae8891, 32'h4157238e} /* (13, 9, 13) {real, imag} */,
  {32'h40a31d54, 32'h4072a9da} /* (13, 9, 12) {real, imag} */,
  {32'hc008e8d2, 32'hc00ee5b2} /* (13, 9, 11) {real, imag} */,
  {32'hc07c2e02, 32'h40132e18} /* (13, 9, 10) {real, imag} */,
  {32'h409460c2, 32'hbfe9059a} /* (13, 9, 9) {real, imag} */,
  {32'hc08543a3, 32'hbe21c470} /* (13, 9, 8) {real, imag} */,
  {32'hbece70d0, 32'hbfcbe05e} /* (13, 9, 7) {real, imag} */,
  {32'h407674c2, 32'hbedb956c} /* (13, 9, 6) {real, imag} */,
  {32'hbf36ada6, 32'h3f3f24e6} /* (13, 9, 5) {real, imag} */,
  {32'hc03b3bc0, 32'h3e147778} /* (13, 9, 4) {real, imag} */,
  {32'h40e8b9b7, 32'hc0dec6e3} /* (13, 9, 3) {real, imag} */,
  {32'h41906e87, 32'hc07eaa59} /* (13, 9, 2) {real, imag} */,
  {32'hc03269a8, 32'h4139026b} /* (13, 9, 1) {real, imag} */,
  {32'h3ddce840, 32'hbf7205c4} /* (13, 9, 0) {real, imag} */,
  {32'hc0980582, 32'h408b5f1d} /* (13, 8, 15) {real, imag} */,
  {32'hc041e014, 32'h4100df34} /* (13, 8, 14) {real, imag} */,
  {32'h40a76f64, 32'hc13b5e3a} /* (13, 8, 13) {real, imag} */,
  {32'h40e48276, 32'hc076e618} /* (13, 8, 12) {real, imag} */,
  {32'h4015e0c0, 32'h3f6159cc} /* (13, 8, 11) {real, imag} */,
  {32'hc022f94e, 32'hbf1f2040} /* (13, 8, 10) {real, imag} */,
  {32'h3fdf92b6, 32'hbecaf6e0} /* (13, 8, 9) {real, imag} */,
  {32'hc024b812, 32'h3e625f50} /* (13, 8, 8) {real, imag} */,
  {32'h4093f186, 32'h40cfeab6} /* (13, 8, 7) {real, imag} */,
  {32'h40488a2e, 32'h4058a754} /* (13, 8, 6) {real, imag} */,
  {32'hc1003160, 32'h4097ee6a} /* (13, 8, 5) {real, imag} */,
  {32'h40070231, 32'hbf0f6cee} /* (13, 8, 4) {real, imag} */,
  {32'hbf99c8b0, 32'hc08cd0b8} /* (13, 8, 3) {real, imag} */,
  {32'hc011cc2c, 32'hbf4b7310} /* (13, 8, 2) {real, imag} */,
  {32'h40dd2d56, 32'hc0f18d8b} /* (13, 8, 1) {real, imag} */,
  {32'h3fed900c, 32'h4096ef3a} /* (13, 8, 0) {real, imag} */,
  {32'h409da5f0, 32'h40ecd5c5} /* (13, 7, 15) {real, imag} */,
  {32'hc10d88d1, 32'h410278eb} /* (13, 7, 14) {real, imag} */,
  {32'hc0cf860a, 32'h41499380} /* (13, 7, 13) {real, imag} */,
  {32'hbffd435e, 32'hc0d913c5} /* (13, 7, 12) {real, imag} */,
  {32'h410c9b20, 32'hc061653c} /* (13, 7, 11) {real, imag} */,
  {32'h3f60da5c, 32'hc0e0bc5e} /* (13, 7, 10) {real, imag} */,
  {32'hbee49470, 32'hc04e1d66} /* (13, 7, 9) {real, imag} */,
  {32'hbf858790, 32'hc0074570} /* (13, 7, 8) {real, imag} */,
  {32'hbeb461e0, 32'h4098e476} /* (13, 7, 7) {real, imag} */,
  {32'h400cbd4b, 32'hc02c3a45} /* (13, 7, 6) {real, imag} */,
  {32'hc006db86, 32'h4043b780} /* (13, 7, 5) {real, imag} */,
  {32'hbfd947ca, 32'h40bd8057} /* (13, 7, 4) {real, imag} */,
  {32'h411513a3, 32'hbe718140} /* (13, 7, 3) {real, imag} */,
  {32'h40fbff46, 32'hc0d3cd36} /* (13, 7, 2) {real, imag} */,
  {32'h404eef29, 32'hc1427f4a} /* (13, 7, 1) {real, imag} */,
  {32'hc1317a88, 32'h3ff257d5} /* (13, 7, 0) {real, imag} */,
  {32'hc09ff3b4, 32'hc14b73a0} /* (13, 6, 15) {real, imag} */,
  {32'h41073174, 32'hc18dacff} /* (13, 6, 14) {real, imag} */,
  {32'h3f3c1140, 32'hc19c9c92} /* (13, 6, 13) {real, imag} */,
  {32'hc055e4b6, 32'h406a5cc0} /* (13, 6, 12) {real, imag} */,
  {32'hc0bf1d9c, 32'hc105efd7} /* (13, 6, 11) {real, imag} */,
  {32'h40b5dfd3, 32'h3fb439b8} /* (13, 6, 10) {real, imag} */,
  {32'h3f01c7c8, 32'h40ff80ea} /* (13, 6, 9) {real, imag} */,
  {32'hbfd61154, 32'h3f351124} /* (13, 6, 8) {real, imag} */,
  {32'h400ea384, 32'h3eb190e8} /* (13, 6, 7) {real, imag} */,
  {32'hc07878ca, 32'h410529b1} /* (13, 6, 6) {real, imag} */,
  {32'hc0448214, 32'hc0b8d3a8} /* (13, 6, 5) {real, imag} */,
  {32'hc1274dea, 32'h40d6c104} /* (13, 6, 4) {real, imag} */,
  {32'hc06be550, 32'hc1a72fb8} /* (13, 6, 3) {real, imag} */,
  {32'h3f1578d8, 32'h41271254} /* (13, 6, 2) {real, imag} */,
  {32'hc10c1cd8, 32'h411d31f6} /* (13, 6, 1) {real, imag} */,
  {32'h3efe14d0, 32'hc0cae7ea} /* (13, 6, 0) {real, imag} */,
  {32'h41efd3ca, 32'hc1cd2ef6} /* (13, 5, 15) {real, imag} */,
  {32'h3e7aef00, 32'hc150a40a} /* (13, 5, 14) {real, imag} */,
  {32'hc18b47b4, 32'h40a48342} /* (13, 5, 13) {real, imag} */,
  {32'hc11331cb, 32'h3f093978} /* (13, 5, 12) {real, imag} */,
  {32'h40732492, 32'h4166fa74} /* (13, 5, 11) {real, imag} */,
  {32'h412355ee, 32'h40afc334} /* (13, 5, 10) {real, imag} */,
  {32'h40ddce8e, 32'h40b1e9e4} /* (13, 5, 9) {real, imag} */,
  {32'h3e0837a0, 32'h3fb3b6a4} /* (13, 5, 8) {real, imag} */,
  {32'hc10cff71, 32'hc0ca0090} /* (13, 5, 7) {real, imag} */,
  {32'h3f2c3170, 32'h4121e0d0} /* (13, 5, 6) {real, imag} */,
  {32'hc04a2b7a, 32'hc0cf09d1} /* (13, 5, 5) {real, imag} */,
  {32'hc15ce405, 32'h412a1d66} /* (13, 5, 4) {real, imag} */,
  {32'hbf7fa840, 32'hbf962dc0} /* (13, 5, 3) {real, imag} */,
  {32'h420706c8, 32'hc116bea8} /* (13, 5, 2) {real, imag} */,
  {32'hc184391a, 32'hc19fa936} /* (13, 5, 1) {real, imag} */,
  {32'hc17c084e, 32'hc01a36a8} /* (13, 5, 0) {real, imag} */,
  {32'h41059c66, 32'h424b1372} /* (13, 4, 15) {real, imag} */,
  {32'h410c05c9, 32'hc07ead0b} /* (13, 4, 14) {real, imag} */,
  {32'h41f5bbfe, 32'hc087eca8} /* (13, 4, 13) {real, imag} */,
  {32'hc1d97a1e, 32'h3f06ee22} /* (13, 4, 12) {real, imag} */,
  {32'h3e5821c0, 32'hc14d4dd1} /* (13, 4, 11) {real, imag} */,
  {32'hc18e0f82, 32'hc138ce88} /* (13, 4, 10) {real, imag} */,
  {32'hbfddf0c4, 32'hbf992b50} /* (13, 4, 9) {real, imag} */,
  {32'hbf36fb74, 32'h40e1920c} /* (13, 4, 8) {real, imag} */,
  {32'h414b44b4, 32'h4022e958} /* (13, 4, 7) {real, imag} */,
  {32'hc145143c, 32'hc0a9e184} /* (13, 4, 6) {real, imag} */,
  {32'hc171db8d, 32'h41a9ad12} /* (13, 4, 5) {real, imag} */,
  {32'hbf7e85e0, 32'hc040590a} /* (13, 4, 4) {real, imag} */,
  {32'h41948262, 32'h4173b858} /* (13, 4, 3) {real, imag} */,
  {32'hbffcd8b0, 32'hc12aff49} /* (13, 4, 2) {real, imag} */,
  {32'h41be7e51, 32'hc0579128} /* (13, 4, 1) {real, imag} */,
  {32'hc0e3d25e, 32'hc08ea9e8} /* (13, 4, 0) {real, imag} */,
  {32'h41adeb40, 32'h409ef271} /* (13, 3, 15) {real, imag} */,
  {32'hc1f4c3fa, 32'h4107d570} /* (13, 3, 14) {real, imag} */,
  {32'h40db6f58, 32'h41d89311} /* (13, 3, 13) {real, imag} */,
  {32'hbf0e65c0, 32'hc0e9e79c} /* (13, 3, 12) {real, imag} */,
  {32'h41602739, 32'hc0c3c8fd} /* (13, 3, 11) {real, imag} */,
  {32'h419ae224, 32'hc13ebee6} /* (13, 3, 10) {real, imag} */,
  {32'h40635bea, 32'h40213b78} /* (13, 3, 9) {real, imag} */,
  {32'h41882aaa, 32'h3fadc4f0} /* (13, 3, 8) {real, imag} */,
  {32'h40a5e9a5, 32'hc094dc16} /* (13, 3, 7) {real, imag} */,
  {32'h40676840, 32'hc093a12f} /* (13, 3, 6) {real, imag} */,
  {32'hc13d209f, 32'h413c4152} /* (13, 3, 5) {real, imag} */,
  {32'h4245901d, 32'h4189a1cd} /* (13, 3, 4) {real, imag} */,
  {32'h41fa49ee, 32'hc1922899} /* (13, 3, 3) {real, imag} */,
  {32'hc166ca74, 32'h41cec1bc} /* (13, 3, 2) {real, imag} */,
  {32'hc18edeb4, 32'hc17d9994} /* (13, 3, 1) {real, imag} */,
  {32'hc1d595ba, 32'hbf1c4fa0} /* (13, 3, 0) {real, imag} */,
  {32'hc137aff6, 32'h4012888c} /* (13, 2, 15) {real, imag} */,
  {32'hc171fc4a, 32'h3ff66d70} /* (13, 2, 14) {real, imag} */,
  {32'h3f31ded4, 32'hc1820feb} /* (13, 2, 13) {real, imag} */,
  {32'h4177d1db, 32'hbf9175b0} /* (13, 2, 12) {real, imag} */,
  {32'h415ead48, 32'hc0a1687d} /* (13, 2, 11) {real, imag} */,
  {32'hc1d2a11b, 32'hc0a78c50} /* (13, 2, 10) {real, imag} */,
  {32'hc1649062, 32'h414ed2fc} /* (13, 2, 9) {real, imag} */,
  {32'hc0bffb26, 32'h4121c2c6} /* (13, 2, 8) {real, imag} */,
  {32'h3dc74d40, 32'hc0843d5d} /* (13, 2, 7) {real, imag} */,
  {32'hc0e725e4, 32'h3f1b4a5c} /* (13, 2, 6) {real, imag} */,
  {32'h4007522a, 32'h40de3613} /* (13, 2, 5) {real, imag} */,
  {32'hbda93080, 32'hc1ab1f01} /* (13, 2, 4) {real, imag} */,
  {32'h4078a271, 32'h4208744a} /* (13, 2, 3) {real, imag} */,
  {32'hc1e6d8d7, 32'h4146c688} /* (13, 2, 2) {real, imag} */,
  {32'h413a0966, 32'h41f00d38} /* (13, 2, 1) {real, imag} */,
  {32'h41d121bc, 32'hc0eefca3} /* (13, 2, 0) {real, imag} */,
  {32'hc2516937, 32'h41c49824} /* (13, 1, 15) {real, imag} */,
  {32'hc0f80fa0, 32'hc1993429} /* (13, 1, 14) {real, imag} */,
  {32'hc18b243a, 32'h41cbc81c} /* (13, 1, 13) {real, imag} */,
  {32'h41ab36b4, 32'hbe1be080} /* (13, 1, 12) {real, imag} */,
  {32'h418e661e, 32'h42271c3c} /* (13, 1, 11) {real, imag} */,
  {32'hc0bbc39e, 32'hc19347da} /* (13, 1, 10) {real, imag} */,
  {32'hc0f4cc7c, 32'hc0c87662} /* (13, 1, 9) {real, imag} */,
  {32'hc0dc9fde, 32'hc08c449a} /* (13, 1, 8) {real, imag} */,
  {32'h40019c78, 32'h40b75862} /* (13, 1, 7) {real, imag} */,
  {32'h41bf301c, 32'hc1733f78} /* (13, 1, 6) {real, imag} */,
  {32'h418d3566, 32'hc2112acc} /* (13, 1, 5) {real, imag} */,
  {32'h4049a2e8, 32'hc21ab26c} /* (13, 1, 4) {real, imag} */,
  {32'h418d1aca, 32'hc1a8beba} /* (13, 1, 3) {real, imag} */,
  {32'hc256087a, 32'h41b1094f} /* (13, 1, 2) {real, imag} */,
  {32'h40971120, 32'hc0205c84} /* (13, 1, 1) {real, imag} */,
  {32'h4174f80d, 32'h41159489} /* (13, 1, 0) {real, imag} */,
  {32'h41a704d9, 32'h420ba1cc} /* (13, 0, 15) {real, imag} */,
  {32'h40331420, 32'hc0b49636} /* (13, 0, 14) {real, imag} */,
  {32'hc10a0884, 32'hc1eb360d} /* (13, 0, 13) {real, imag} */,
  {32'hc0db4f48, 32'hc15c696d} /* (13, 0, 12) {real, imag} */,
  {32'hc0524c96, 32'h42586c30} /* (13, 0, 11) {real, imag} */,
  {32'hc1049e7a, 32'hc1065c71} /* (13, 0, 10) {real, imag} */,
  {32'h419aa66d, 32'hbd1cb300} /* (13, 0, 9) {real, imag} */,
  {32'hc093988a, 32'hc16a368e} /* (13, 0, 8) {real, imag} */,
  {32'h406319e6, 32'h40928dda} /* (13, 0, 7) {real, imag} */,
  {32'hbf965060, 32'hbf3ade50} /* (13, 0, 6) {real, imag} */,
  {32'h408867cb, 32'hc21c2e24} /* (13, 0, 5) {real, imag} */,
  {32'hc242f0eb, 32'h421875da} /* (13, 0, 4) {real, imag} */,
  {32'h41a27adc, 32'h4110fb86} /* (13, 0, 3) {real, imag} */,
  {32'h425544d8, 32'hc1ad18b8} /* (13, 0, 2) {real, imag} */,
  {32'hc05e9dc8, 32'hc25b8878} /* (13, 0, 1) {real, imag} */,
  {32'h41d7bf2c, 32'h4256a928} /* (13, 0, 0) {real, imag} */,
  {32'hc1c87d5b, 32'hc19262fe} /* (12, 15, 15) {real, imag} */,
  {32'h41f966ae, 32'hbf5ed1d4} /* (12, 15, 14) {real, imag} */,
  {32'hc11097f6, 32'hc1ef5f24} /* (12, 15, 13) {real, imag} */,
  {32'h41135992, 32'hbfe8efc8} /* (12, 15, 12) {real, imag} */,
  {32'hc1533dd2, 32'hc136e54c} /* (12, 15, 11) {real, imag} */,
  {32'hc0c966b2, 32'h3ecc8ec0} /* (12, 15, 10) {real, imag} */,
  {32'hbff46470, 32'hbff594a8} /* (12, 15, 9) {real, imag} */,
  {32'hc1016918, 32'hc04b7d36} /* (12, 15, 8) {real, imag} */,
  {32'h4042f6a8, 32'h3f96f948} /* (12, 15, 7) {real, imag} */,
  {32'h41062ca7, 32'hc191f4e9} /* (12, 15, 6) {real, imag} */,
  {32'hc120ca24, 32'h3f1508f8} /* (12, 15, 5) {real, imag} */,
  {32'h40b348c2, 32'h41b09574} /* (12, 15, 4) {real, imag} */,
  {32'hc18155ca, 32'h42168976} /* (12, 15, 3) {real, imag} */,
  {32'hc1cff37a, 32'hc088bfe0} /* (12, 15, 2) {real, imag} */,
  {32'h3ef49900, 32'hc25ab231} /* (12, 15, 1) {real, imag} */,
  {32'hc14a15dc, 32'h40ed6e25} /* (12, 15, 0) {real, imag} */,
  {32'h4119512f, 32'hc13699f6} /* (12, 14, 15) {real, imag} */,
  {32'h413eec6d, 32'h413d5404} /* (12, 14, 14) {real, imag} */,
  {32'h418facfb, 32'h417b8a63} /* (12, 14, 13) {real, imag} */,
  {32'hc02f1524, 32'h41bdf84c} /* (12, 14, 12) {real, imag} */,
  {32'hc03671c0, 32'h4108d5e8} /* (12, 14, 11) {real, imag} */,
  {32'h41795ce9, 32'hc14bb7da} /* (12, 14, 10) {real, imag} */,
  {32'hc1031bf9, 32'h4030a9bf} /* (12, 14, 9) {real, imag} */,
  {32'h415e0960, 32'hc032c804} /* (12, 14, 8) {real, imag} */,
  {32'hbfcace2a, 32'hc013b87f} /* (12, 14, 7) {real, imag} */,
  {32'hbf5e03f0, 32'h406e7778} /* (12, 14, 6) {real, imag} */,
  {32'h4156fbd8, 32'hc0dbe7d4} /* (12, 14, 5) {real, imag} */,
  {32'h408ee514, 32'hc13bd327} /* (12, 14, 4) {real, imag} */,
  {32'h4212f34c, 32'hc1826fd6} /* (12, 14, 3) {real, imag} */,
  {32'hc0f50116, 32'h42018560} /* (12, 14, 2) {real, imag} */,
  {32'h418e56e6, 32'hc1d9f9db} /* (12, 14, 1) {real, imag} */,
  {32'hc214d998, 32'h41bccf78} /* (12, 14, 0) {real, imag} */,
  {32'hc0e9873a, 32'hc1b5b49e} /* (12, 13, 15) {real, imag} */,
  {32'h412dda02, 32'hc124d9da} /* (12, 13, 14) {real, imag} */,
  {32'hbf151bb8, 32'h4148bead} /* (12, 13, 13) {real, imag} */,
  {32'hc1d9bd4a, 32'hc1069c84} /* (12, 13, 12) {real, imag} */,
  {32'h41a2cca4, 32'hc181baa4} /* (12, 13, 11) {real, imag} */,
  {32'h4146ef64, 32'hbfeb9318} /* (12, 13, 10) {real, imag} */,
  {32'hc05b4e06, 32'hc107fd96} /* (12, 13, 9) {real, imag} */,
  {32'h409ed4da, 32'h3f656e5e} /* (12, 13, 8) {real, imag} */,
  {32'h40de76d9, 32'hbfd6966e} /* (12, 13, 7) {real, imag} */,
  {32'h4150e01c, 32'h414c6744} /* (12, 13, 6) {real, imag} */,
  {32'h4126afa1, 32'hc0f1061e} /* (12, 13, 5) {real, imag} */,
  {32'hc0fcd7de, 32'h4126358a} /* (12, 13, 4) {real, imag} */,
  {32'hc16bce66, 32'h4178552f} /* (12, 13, 3) {real, imag} */,
  {32'h408955cd, 32'h40c06aec} /* (12, 13, 2) {real, imag} */,
  {32'hc1ba88b6, 32'hc0fcddde} /* (12, 13, 1) {real, imag} */,
  {32'h4154f2e7, 32'hc09c0e30} /* (12, 13, 0) {real, imag} */,
  {32'h414c27e4, 32'hc0e57e80} /* (12, 12, 15) {real, imag} */,
  {32'hc0cf3b80, 32'hc13a2e81} /* (12, 12, 14) {real, imag} */,
  {32'hc15ba2e7, 32'h411e7bc4} /* (12, 12, 13) {real, imag} */,
  {32'h41058a12, 32'hbfab3634} /* (12, 12, 12) {real, imag} */,
  {32'h41466f7a, 32'hbf4b3198} /* (12, 12, 11) {real, imag} */,
  {32'h404e5870, 32'h41068e82} /* (12, 12, 10) {real, imag} */,
  {32'h40793a5d, 32'h4033ba14} /* (12, 12, 9) {real, imag} */,
  {32'h4082e7fa, 32'h3ca01780} /* (12, 12, 8) {real, imag} */,
  {32'hbe2f31d0, 32'hc13a1a29} /* (12, 12, 7) {real, imag} */,
  {32'hc1a73206, 32'h40d18cff} /* (12, 12, 6) {real, imag} */,
  {32'h3fe41490, 32'hc109448a} /* (12, 12, 5) {real, imag} */,
  {32'h410f4a92, 32'hc10be3c6} /* (12, 12, 4) {real, imag} */,
  {32'hc0db8d6a, 32'hc1bea416} /* (12, 12, 3) {real, imag} */,
  {32'h4119b924, 32'hc15565cd} /* (12, 12, 2) {real, imag} */,
  {32'h41fd8e96, 32'h41346126} /* (12, 12, 1) {real, imag} */,
  {32'h417031f7, 32'hc0c9df82} /* (12, 12, 0) {real, imag} */,
  {32'h3f53e0a0, 32'hc1695ef2} /* (12, 11, 15) {real, imag} */,
  {32'hbe899a10, 32'h4150ddd8} /* (12, 11, 14) {real, imag} */,
  {32'hc1e79d0f, 32'hc1f618d7} /* (12, 11, 13) {real, imag} */,
  {32'h409fb588, 32'hc1243476} /* (12, 11, 12) {real, imag} */,
  {32'h4111bfaa, 32'h41215d8c} /* (12, 11, 11) {real, imag} */,
  {32'h402785e2, 32'hc0240b18} /* (12, 11, 10) {real, imag} */,
  {32'h409fb444, 32'hbfc7ac1c} /* (12, 11, 9) {real, imag} */,
  {32'h403ded21, 32'hc04fb243} /* (12, 11, 8) {real, imag} */,
  {32'h4097d764, 32'h3faa595c} /* (12, 11, 7) {real, imag} */,
  {32'hc04a961e, 32'h4112a584} /* (12, 11, 6) {real, imag} */,
  {32'hc16e1816, 32'hbff3847c} /* (12, 11, 5) {real, imag} */,
  {32'h40a7a624, 32'h412c5426} /* (12, 11, 4) {real, imag} */,
  {32'hc0ac9f7c, 32'h415f4efe} /* (12, 11, 3) {real, imag} */,
  {32'hc0af2901, 32'h4176c5a2} /* (12, 11, 2) {real, imag} */,
  {32'hc21df71e, 32'hc12677f6} /* (12, 11, 1) {real, imag} */,
  {32'hbe2cd4b0, 32'hc09ab82a} /* (12, 11, 0) {real, imag} */,
  {32'hbfdbf282, 32'h419d92ae} /* (12, 10, 15) {real, imag} */,
  {32'h419376df, 32'h40dc7408} /* (12, 10, 14) {real, imag} */,
  {32'hc0f6660a, 32'h4174bd40} /* (12, 10, 13) {real, imag} */,
  {32'h41383e3a, 32'hc1986434} /* (12, 10, 12) {real, imag} */,
  {32'hc069075d, 32'hc0a08110} /* (12, 10, 11) {real, imag} */,
  {32'h408c6557, 32'hbffd5712} /* (12, 10, 10) {real, imag} */,
  {32'hbf7dc595, 32'h3cd94e00} /* (12, 10, 9) {real, imag} */,
  {32'h40805e0d, 32'hc01f213c} /* (12, 10, 8) {real, imag} */,
  {32'hc0258bda, 32'h40ac5fd6} /* (12, 10, 7) {real, imag} */,
  {32'h4003e7c2, 32'hbeda9418} /* (12, 10, 6) {real, imag} */,
  {32'hc006c46f, 32'h3feae598} /* (12, 10, 5) {real, imag} */,
  {32'hc161b15c, 32'h4088421e} /* (12, 10, 4) {real, imag} */,
  {32'hbf622e24, 32'hbf9cf2e4} /* (12, 10, 3) {real, imag} */,
  {32'hbf9d0f50, 32'h41167734} /* (12, 10, 2) {real, imag} */,
  {32'hc0203b4b, 32'hc1f7a788} /* (12, 10, 1) {real, imag} */,
  {32'hc14a99aa, 32'hc1ed5bc4} /* (12, 10, 0) {real, imag} */,
  {32'h405a7f5d, 32'h413dcec0} /* (12, 9, 15) {real, imag} */,
  {32'h4118b0f2, 32'hc02b2af0} /* (12, 9, 14) {real, imag} */,
  {32'hc03a15df, 32'hc0b0ee18} /* (12, 9, 13) {real, imag} */,
  {32'hbf82423c, 32'hc09b0844} /* (12, 9, 12) {real, imag} */,
  {32'h40a05c26, 32'h4031b0d8} /* (12, 9, 11) {real, imag} */,
  {32'hc0da16db, 32'hc0240535} /* (12, 9, 10) {real, imag} */,
  {32'hbf3f1eec, 32'hc006ea6b} /* (12, 9, 9) {real, imag} */,
  {32'h3f808cd9, 32'hbebb8bc0} /* (12, 9, 8) {real, imag} */,
  {32'h4070cfb5, 32'hbfcefcf6} /* (12, 9, 7) {real, imag} */,
  {32'h3eba7050, 32'h406f0ceb} /* (12, 9, 6) {real, imag} */,
  {32'hbf6561cc, 32'hbf693092} /* (12, 9, 5) {real, imag} */,
  {32'hc176e5ac, 32'h3e3c3bc0} /* (12, 9, 4) {real, imag} */,
  {32'h4093edea, 32'h3fa79ca8} /* (12, 9, 3) {real, imag} */,
  {32'hc100d872, 32'hc0c46320} /* (12, 9, 2) {real, imag} */,
  {32'hbf49617c, 32'hc14fbfa8} /* (12, 9, 1) {real, imag} */,
  {32'h406142e8, 32'h4187b073} /* (12, 9, 0) {real, imag} */,
  {32'h40f349ab, 32'h3fa95f0d} /* (12, 8, 15) {real, imag} */,
  {32'h40c5a042, 32'h40d1c4a8} /* (12, 8, 14) {real, imag} */,
  {32'hbfc3da1d, 32'hc0980a1f} /* (12, 8, 13) {real, imag} */,
  {32'h4060d6f8, 32'h3fa0cc58} /* (12, 8, 12) {real, imag} */,
  {32'hc0ade486, 32'h409ba7f0} /* (12, 8, 11) {real, imag} */,
  {32'h409ed5ee, 32'hc03e18b2} /* (12, 8, 10) {real, imag} */,
  {32'hbed097ac, 32'hbe29c3b4} /* (12, 8, 9) {real, imag} */,
  {32'hbfdb6720, 32'hbf9fb3fa} /* (12, 8, 8) {real, imag} */,
  {32'h3ea4f3ec, 32'h3fc0f9e4} /* (12, 8, 7) {real, imag} */,
  {32'h40dfced6, 32'hc05f857e} /* (12, 8, 6) {real, imag} */,
  {32'hbfcb4e93, 32'hc04e3c88} /* (12, 8, 5) {real, imag} */,
  {32'hc09642bc, 32'hc10e15b5} /* (12, 8, 4) {real, imag} */,
  {32'hbfacc64f, 32'h400a8810} /* (12, 8, 3) {real, imag} */,
  {32'hc0a2a1b2, 32'hbedddb20} /* (12, 8, 2) {real, imag} */,
  {32'h41687344, 32'hbeb1e451} /* (12, 8, 1) {real, imag} */,
  {32'hc152d034, 32'hc012db7b} /* (12, 8, 0) {real, imag} */,
  {32'hc1acb8c7, 32'hc0cdaad2} /* (12, 7, 15) {real, imag} */,
  {32'h40c291ce, 32'h40a25fd4} /* (12, 7, 14) {real, imag} */,
  {32'hbefb29a8, 32'h407501eb} /* (12, 7, 13) {real, imag} */,
  {32'hc028de13, 32'h3d7616a0} /* (12, 7, 12) {real, imag} */,
  {32'hbfc87eab, 32'hc031c64c} /* (12, 7, 11) {real, imag} */,
  {32'h4025609d, 32'h40c7b2a8} /* (12, 7, 10) {real, imag} */,
  {32'hbf5b0778, 32'hbf134e53} /* (12, 7, 9) {real, imag} */,
  {32'h3f2f7b9a, 32'hc00718c4} /* (12, 7, 8) {real, imag} */,
  {32'hbe6f3b60, 32'h3cdf71a0} /* (12, 7, 7) {real, imag} */,
  {32'hbfa0a110, 32'hc09b1fac} /* (12, 7, 6) {real, imag} */,
  {32'h4084cfe6, 32'h3fda7c6c} /* (12, 7, 5) {real, imag} */,
  {32'h4067b209, 32'hc017f620} /* (12, 7, 4) {real, imag} */,
  {32'hc0d406a6, 32'h3f631f1c} /* (12, 7, 3) {real, imag} */,
  {32'hc0665015, 32'hc0cc807c} /* (12, 7, 2) {real, imag} */,
  {32'h40d1347b, 32'h401be7eb} /* (12, 7, 1) {real, imag} */,
  {32'h3d301e60, 32'h4048661c} /* (12, 7, 0) {real, imag} */,
  {32'h411f5a2a, 32'hc105ff69} /* (12, 6, 15) {real, imag} */,
  {32'h40a3e09e, 32'hc1afe2b8} /* (12, 6, 14) {real, imag} */,
  {32'h4144beb6, 32'hbfcf2068} /* (12, 6, 13) {real, imag} */,
  {32'h4056e09c, 32'h41006690} /* (12, 6, 12) {real, imag} */,
  {32'h4122071a, 32'h40dae88d} /* (12, 6, 11) {real, imag} */,
  {32'hc077008c, 32'hbfab8924} /* (12, 6, 10) {real, imag} */,
  {32'hbf99be10, 32'hbf54d212} /* (12, 6, 9) {real, imag} */,
  {32'hbf5c4020, 32'h401aa6f5} /* (12, 6, 8) {real, imag} */,
  {32'h3f375960, 32'hbfa2fbcb} /* (12, 6, 7) {real, imag} */,
  {32'hc1049fd5, 32'h3fdecca4} /* (12, 6, 6) {real, imag} */,
  {32'hc0766818, 32'hc055ba6a} /* (12, 6, 5) {real, imag} */,
  {32'hc0bef522, 32'hc0b413de} /* (12, 6, 4) {real, imag} */,
  {32'h40c3ee54, 32'h3e9d6680} /* (12, 6, 3) {real, imag} */,
  {32'h41db0ea8, 32'h40a55250} /* (12, 6, 2) {real, imag} */,
  {32'hc1dcee71, 32'hbfed5828} /* (12, 6, 1) {real, imag} */,
  {32'hc095c902, 32'h40c2239a} /* (12, 6, 0) {real, imag} */,
  {32'hc19aa46c, 32'h3beff000} /* (12, 5, 15) {real, imag} */,
  {32'h4101c12a, 32'hc145ba64} /* (12, 5, 14) {real, imag} */,
  {32'h401211ec, 32'h3fd6c916} /* (12, 5, 13) {real, imag} */,
  {32'h41031999, 32'h40b8dba6} /* (12, 5, 12) {real, imag} */,
  {32'h401fa6da, 32'hc06c01b1} /* (12, 5, 11) {real, imag} */,
  {32'hc0f56b64, 32'h401dd72a} /* (12, 5, 10) {real, imag} */,
  {32'hbfaac7c8, 32'hbf2fc8a0} /* (12, 5, 9) {real, imag} */,
  {32'h3f4b7d20, 32'hc0877a1c} /* (12, 5, 8) {real, imag} */,
  {32'hc0bd6b36, 32'h3ed1c760} /* (12, 5, 7) {real, imag} */,
  {32'h3f708100, 32'hc0631f32} /* (12, 5, 6) {real, imag} */,
  {32'h3f8984bc, 32'h40d82fe0} /* (12, 5, 5) {real, imag} */,
  {32'h41135861, 32'hc152c53f} /* (12, 5, 4) {real, imag} */,
  {32'hc187c666, 32'hc0f1c08e} /* (12, 5, 3) {real, imag} */,
  {32'hbfa6ad60, 32'h4195a684} /* (12, 5, 2) {real, imag} */,
  {32'hc21adf51, 32'h41b8d409} /* (12, 5, 1) {real, imag} */,
  {32'hc1849d7e, 32'hc1aef3c7} /* (12, 5, 0) {real, imag} */,
  {32'h418f4d03, 32'hc199d605} /* (12, 4, 15) {real, imag} */,
  {32'hc1cbb65c, 32'hc163b66c} /* (12, 4, 14) {real, imag} */,
  {32'h410db9b5, 32'hc159a24c} /* (12, 4, 13) {real, imag} */,
  {32'h3f8230e0, 32'hc0a13e1e} /* (12, 4, 12) {real, imag} */,
  {32'h40df55c3, 32'hc0d59dad} /* (12, 4, 11) {real, imag} */,
  {32'h415a65c3, 32'hc0f262e0} /* (12, 4, 10) {real, imag} */,
  {32'hbf5dca50, 32'h40bc709a} /* (12, 4, 9) {real, imag} */,
  {32'h40d645d0, 32'hbffbcee0} /* (12, 4, 8) {real, imag} */,
  {32'h40bbb21a, 32'hc0e480d2} /* (12, 4, 7) {real, imag} */,
  {32'hbeb15f60, 32'h3fc646a2} /* (12, 4, 6) {real, imag} */,
  {32'h40b3539b, 32'h3ff337f4} /* (12, 4, 5) {real, imag} */,
  {32'hc207d26d, 32'hbea2df60} /* (12, 4, 4) {real, imag} */,
  {32'h40af7e5c, 32'h4023655e} /* (12, 4, 3) {real, imag} */,
  {32'hc0ebe2fa, 32'h41bd6ce6} /* (12, 4, 2) {real, imag} */,
  {32'hbfbe40c0, 32'h4066cea0} /* (12, 4, 1) {real, imag} */,
  {32'hc0b12778, 32'hc15d507a} /* (12, 4, 0) {real, imag} */,
  {32'hc181ad80, 32'h415cd614} /* (12, 3, 15) {real, imag} */,
  {32'h4139aefd, 32'hc102fabc} /* (12, 3, 14) {real, imag} */,
  {32'hbfa3c100, 32'hc0ce10bc} /* (12, 3, 13) {real, imag} */,
  {32'h410a888b, 32'h3f8c14c4} /* (12, 3, 12) {real, imag} */,
  {32'h40faa19e, 32'h41b576e2} /* (12, 3, 11) {real, imag} */,
  {32'hc090aa31, 32'hc0e26337} /* (12, 3, 10) {real, imag} */,
  {32'hbfdd2d3c, 32'hc120e050} /* (12, 3, 9) {real, imag} */,
  {32'hc1019c76, 32'h3f6b1e38} /* (12, 3, 8) {real, imag} */,
  {32'hc10cfc66, 32'hc169794c} /* (12, 3, 7) {real, imag} */,
  {32'h4188bbb3, 32'h4115d508} /* (12, 3, 6) {real, imag} */,
  {32'hc10990fb, 32'hc0cbe56e} /* (12, 3, 5) {real, imag} */,
  {32'hc165af11, 32'hc0cc8e33} /* (12, 3, 4) {real, imag} */,
  {32'hc1260a4e, 32'h415bdbf6} /* (12, 3, 3) {real, imag} */,
  {32'hc13d4489, 32'hc1c52ba6} /* (12, 3, 2) {real, imag} */,
  {32'hc1868880, 32'hbe97dc50} /* (12, 3, 1) {real, imag} */,
  {32'h41296134, 32'hc08689a1} /* (12, 3, 0) {real, imag} */,
  {32'hc250856f, 32'h41a538eb} /* (12, 2, 15) {real, imag} */,
  {32'h42108e05, 32'hc0ac813e} /* (12, 2, 14) {real, imag} */,
  {32'hc117629f, 32'hc0857f76} /* (12, 2, 13) {real, imag} */,
  {32'hbf1b39b0, 32'h41bd5e46} /* (12, 2, 12) {real, imag} */,
  {32'hc0e5385e, 32'hc162efe9} /* (12, 2, 11) {real, imag} */,
  {32'h40272f42, 32'h41773f09} /* (12, 2, 10) {real, imag} */,
  {32'hc154c38b, 32'hc0232086} /* (12, 2, 9) {real, imag} */,
  {32'hc09423a4, 32'h41009b9c} /* (12, 2, 8) {real, imag} */,
  {32'hc089e82e, 32'h412e19ae} /* (12, 2, 7) {real, imag} */,
  {32'h41457fdc, 32'hc14882bb} /* (12, 2, 6) {real, imag} */,
  {32'hc155fb6d, 32'hc16b38ff} /* (12, 2, 5) {real, imag} */,
  {32'h4031bc7c, 32'h3e2998c0} /* (12, 2, 4) {real, imag} */,
  {32'hc10c686d, 32'hc1adb1f6} /* (12, 2, 3) {real, imag} */,
  {32'h41ddca80, 32'hc19f5f7a} /* (12, 2, 2) {real, imag} */,
  {32'h420dfc9d, 32'h4117957e} /* (12, 2, 1) {real, imag} */,
  {32'hc1a28221, 32'h425d2115} /* (12, 2, 0) {real, imag} */,
  {32'h42086af1, 32'h420ca0f6} /* (12, 1, 15) {real, imag} */,
  {32'hc22bf616, 32'h403e64ed} /* (12, 1, 14) {real, imag} */,
  {32'hc191d61a, 32'h40841248} /* (12, 1, 13) {real, imag} */,
  {32'h3f8d3d50, 32'hc0d006f4} /* (12, 1, 12) {real, imag} */,
  {32'hc19a0091, 32'h413040b4} /* (12, 1, 11) {real, imag} */,
  {32'hc0afe29b, 32'h40a19bca} /* (12, 1, 10) {real, imag} */,
  {32'h413a6e82, 32'h3f1bead8} /* (12, 1, 9) {real, imag} */,
  {32'hc0dff8e8, 32'hc100d31e} /* (12, 1, 8) {real, imag} */,
  {32'hc05a5d8e, 32'hc0d2adad} /* (12, 1, 7) {real, imag} */,
  {32'h3fd2b5c4, 32'h415af9bb} /* (12, 1, 6) {real, imag} */,
  {32'hc130331a, 32'h40328468} /* (12, 1, 5) {real, imag} */,
  {32'h41b88401, 32'h419ac937} /* (12, 1, 4) {real, imag} */,
  {32'hbf89ffe8, 32'hbf9e476e} /* (12, 1, 3) {real, imag} */,
  {32'h4191510c, 32'h40d857b4} /* (12, 1, 2) {real, imag} */,
  {32'h402435b0, 32'hc1366f82} /* (12, 1, 1) {real, imag} */,
  {32'h4299f14a, 32'hc237507c} /* (12, 1, 0) {real, imag} */,
  {32'h3f1ef1e0, 32'h420e657a} /* (12, 0, 15) {real, imag} */,
  {32'hc103774a, 32'h3fb57334} /* (12, 0, 14) {real, imag} */,
  {32'h406fd114, 32'h419c9117} /* (12, 0, 13) {real, imag} */,
  {32'hc1a8eb9e, 32'h41d4805c} /* (12, 0, 12) {real, imag} */,
  {32'hc03b14ec, 32'hc1ddfb76} /* (12, 0, 11) {real, imag} */,
  {32'hc1087b82, 32'h3f813251} /* (12, 0, 10) {real, imag} */,
  {32'hc02de12e, 32'h40f1aba8} /* (12, 0, 9) {real, imag} */,
  {32'hbf8e5470, 32'h3f9913ec} /* (12, 0, 8) {real, imag} */,
  {32'h412c7012, 32'h40808c5c} /* (12, 0, 7) {real, imag} */,
  {32'hc0ab4d57, 32'h3fc739af} /* (12, 0, 6) {real, imag} */,
  {32'h415df689, 32'h41a1b00a} /* (12, 0, 5) {real, imag} */,
  {32'h4144b7cc, 32'hc113c7a4} /* (12, 0, 4) {real, imag} */,
  {32'h41d0a76a, 32'hc21a2840} /* (12, 0, 3) {real, imag} */,
  {32'hc207aa2c, 32'h4106e6ea} /* (12, 0, 2) {real, imag} */,
  {32'hc23344c8, 32'h413b10c7} /* (12, 0, 1) {real, imag} */,
  {32'hc199457d, 32'hc028cad2} /* (12, 0, 0) {real, imag} */,
  {32'h414ae5b4, 32'h4113435e} /* (11, 15, 15) {real, imag} */,
  {32'h4136bffc, 32'hc1fd01b6} /* (11, 15, 14) {real, imag} */,
  {32'hc0bc54b2, 32'h4204a280} /* (11, 15, 13) {real, imag} */,
  {32'h40a0ef96, 32'h40928e32} /* (11, 15, 12) {real, imag} */,
  {32'hc041b11d, 32'h41be1ccf} /* (11, 15, 11) {real, imag} */,
  {32'h411f0e22, 32'hc0cc2306} /* (11, 15, 10) {real, imag} */,
  {32'h3fdbe650, 32'hbcc6e300} /* (11, 15, 9) {real, imag} */,
  {32'hc02320c2, 32'hbfd95e00} /* (11, 15, 8) {real, imag} */,
  {32'hc10e6b52, 32'hc0f1ef93} /* (11, 15, 7) {real, imag} */,
  {32'hbfd31a50, 32'h40fd1202} /* (11, 15, 6) {real, imag} */,
  {32'hc09b05b8, 32'hc0c34d1c} /* (11, 15, 5) {real, imag} */,
  {32'h4101feac, 32'hc1ad2abc} /* (11, 15, 4) {real, imag} */,
  {32'h413abc9f, 32'hc11bb53c} /* (11, 15, 3) {real, imag} */,
  {32'hc23c1972, 32'h41d157d8} /* (11, 15, 2) {real, imag} */,
  {32'h41dddb7e, 32'hc119d044} /* (11, 15, 1) {real, imag} */,
  {32'h4189bcc7, 32'hc1e41ccc} /* (11, 15, 0) {real, imag} */,
  {32'h423177de, 32'h4183895f} /* (11, 14, 15) {real, imag} */,
  {32'h4211a8a6, 32'h4184c17d} /* (11, 14, 14) {real, imag} */,
  {32'h41c5fb54, 32'h3fad3e0c} /* (11, 14, 13) {real, imag} */,
  {32'hc179ba15, 32'hc0b99348} /* (11, 14, 12) {real, imag} */,
  {32'hc12b22b9, 32'hbf97005c} /* (11, 14, 11) {real, imag} */,
  {32'h4091ea5d, 32'h40e0ff7e} /* (11, 14, 10) {real, imag} */,
  {32'hc0d169a2, 32'hbfe9c266} /* (11, 14, 9) {real, imag} */,
  {32'hbf8dca34, 32'h3e2f93e0} /* (11, 14, 8) {real, imag} */,
  {32'h3f128350, 32'h40ca663e} /* (11, 14, 7) {real, imag} */,
  {32'hc16aae9e, 32'hc152e8c5} /* (11, 14, 6) {real, imag} */,
  {32'h40693995, 32'hc1490b28} /* (11, 14, 5) {real, imag} */,
  {32'hc1169973, 32'h41da9614} /* (11, 14, 4) {real, imag} */,
  {32'hc1a9951c, 32'hc0ecad2f} /* (11, 14, 3) {real, imag} */,
  {32'hc0ad3d0c, 32'hc19fd043} /* (11, 14, 2) {real, imag} */,
  {32'h41c3cd6c, 32'hc196d6e5} /* (11, 14, 1) {real, imag} */,
  {32'h40ab4d79, 32'h402bf8c6} /* (11, 14, 0) {real, imag} */,
  {32'hc18188a1, 32'h3fca05ec} /* (11, 13, 15) {real, imag} */,
  {32'hc00fb39a, 32'hc0dfcc32} /* (11, 13, 14) {real, imag} */,
  {32'h41ac0f44, 32'hc19156be} /* (11, 13, 13) {real, imag} */,
  {32'hc1427622, 32'hc0335813} /* (11, 13, 12) {real, imag} */,
  {32'hc03da7e0, 32'h41af3f2e} /* (11, 13, 11) {real, imag} */,
  {32'h40ce635f, 32'h3e6a81d8} /* (11, 13, 10) {real, imag} */,
  {32'hbfff931e, 32'hc01c4052} /* (11, 13, 9) {real, imag} */,
  {32'hbf0a9c54, 32'hc0970d2b} /* (11, 13, 8) {real, imag} */,
  {32'hc061f723, 32'hc07bfe8e} /* (11, 13, 7) {real, imag} */,
  {32'h41483ae2, 32'h3f8ff313} /* (11, 13, 6) {real, imag} */,
  {32'h4188d17a, 32'hc096f100} /* (11, 13, 5) {real, imag} */,
  {32'h416ec6d8, 32'hc06aad09} /* (11, 13, 4) {real, imag} */,
  {32'h41581a44, 32'h40c06411} /* (11, 13, 3) {real, imag} */,
  {32'h40248272, 32'h3e9d17e0} /* (11, 13, 2) {real, imag} */,
  {32'h414787e5, 32'hc14f63a0} /* (11, 13, 1) {real, imag} */,
  {32'h40bb6f0e, 32'h411283c4} /* (11, 13, 0) {real, imag} */,
  {32'hc1a800e6, 32'h4129de94} /* (11, 12, 15) {real, imag} */,
  {32'hc19f2fad, 32'hc10184f0} /* (11, 12, 14) {real, imag} */,
  {32'hbfcd11c0, 32'h412a2774} /* (11, 12, 13) {real, imag} */,
  {32'hc1364822, 32'h3e384e10} /* (11, 12, 12) {real, imag} */,
  {32'h40dbd590, 32'h3ef752d0} /* (11, 12, 11) {real, imag} */,
  {32'hbf9b5abc, 32'h3d8d7630} /* (11, 12, 10) {real, imag} */,
  {32'h407f36ce, 32'hc0c12c32} /* (11, 12, 9) {real, imag} */,
  {32'hbf63799c, 32'hbc3bb600} /* (11, 12, 8) {real, imag} */,
  {32'h3f93cb5c, 32'h400487b4} /* (11, 12, 7) {real, imag} */,
  {32'h413ec9ae, 32'hc02d8ba6} /* (11, 12, 6) {real, imag} */,
  {32'hc0d8f172, 32'h40c71d03} /* (11, 12, 5) {real, imag} */,
  {32'h3fbd4860, 32'hc0f66f82} /* (11, 12, 4) {real, imag} */,
  {32'h40c006ca, 32'h4153d98e} /* (11, 12, 3) {real, imag} */,
  {32'h3fb52060, 32'h40cfdc08} /* (11, 12, 2) {real, imag} */,
  {32'hbf8152b8, 32'h42041884} /* (11, 12, 1) {real, imag} */,
  {32'hc0d9bcd4, 32'hc03ecd0a} /* (11, 12, 0) {real, imag} */,
  {32'h41b70204, 32'hc0eeb99a} /* (11, 11, 15) {real, imag} */,
  {32'hc13edc92, 32'h40bbea82} /* (11, 11, 14) {real, imag} */,
  {32'hc0416a54, 32'hc139b74b} /* (11, 11, 13) {real, imag} */,
  {32'h410b6d64, 32'h4118b278} /* (11, 11, 12) {real, imag} */,
  {32'h40dfe2ba, 32'h3f7da3e4} /* (11, 11, 11) {real, imag} */,
  {32'hc0c72c8c, 32'h3ff7a75c} /* (11, 11, 10) {real, imag} */,
  {32'hc0682b7a, 32'hbf6c9220} /* (11, 11, 9) {real, imag} */,
  {32'hbae74000, 32'h4056a8c3} /* (11, 11, 8) {real, imag} */,
  {32'h3f5b0348, 32'h40404028} /* (11, 11, 7) {real, imag} */,
  {32'h3fe335b6, 32'h4089d8e9} /* (11, 11, 6) {real, imag} */,
  {32'h3f6c630c, 32'h40da91de} /* (11, 11, 5) {real, imag} */,
  {32'hc06e7502, 32'h408947b3} /* (11, 11, 4) {real, imag} */,
  {32'hc0af7aa2, 32'hc1828dc5} /* (11, 11, 3) {real, imag} */,
  {32'hc014b50a, 32'hc1a94ffa} /* (11, 11, 2) {real, imag} */,
  {32'hbf98e3f8, 32'h417b1ac7} /* (11, 11, 1) {real, imag} */,
  {32'hc130ebf5, 32'h3f5359f4} /* (11, 11, 0) {real, imag} */,
  {32'hc1a50139, 32'hc0bdaf90} /* (11, 10, 15) {real, imag} */,
  {32'hbf8bea38, 32'hbe849a30} /* (11, 10, 14) {real, imag} */,
  {32'h40b9820c, 32'hc09239dc} /* (11, 10, 13) {real, imag} */,
  {32'h40118a72, 32'h411f9058} /* (11, 10, 12) {real, imag} */,
  {32'hc0df2864, 32'hbfd83806} /* (11, 10, 11) {real, imag} */,
  {32'hc099fb27, 32'hbf39236c} /* (11, 10, 10) {real, imag} */,
  {32'h3f909226, 32'hbebd7c9c} /* (11, 10, 9) {real, imag} */,
  {32'hbe9a40c0, 32'h4036ee7e} /* (11, 10, 8) {real, imag} */,
  {32'hc010293f, 32'hbfed18fd} /* (11, 10, 7) {real, imag} */,
  {32'hbf83095c, 32'h401a539d} /* (11, 10, 6) {real, imag} */,
  {32'h3f55a444, 32'hc0cb76b2} /* (11, 10, 5) {real, imag} */,
  {32'h4017442e, 32'h40815ba8} /* (11, 10, 4) {real, imag} */,
  {32'hc0dccd60, 32'h409ded3c} /* (11, 10, 3) {real, imag} */,
  {32'hc190d96e, 32'hbdaff100} /* (11, 10, 2) {real, imag} */,
  {32'hc0e5c6d4, 32'hc08092ec} /* (11, 10, 1) {real, imag} */,
  {32'h414f8b02, 32'h409a6211} /* (11, 10, 0) {real, imag} */,
  {32'hc0dcce66, 32'hc1087e7c} /* (11, 9, 15) {real, imag} */,
  {32'h404f8c46, 32'hc0a610a2} /* (11, 9, 14) {real, imag} */,
  {32'h40e27b27, 32'hc0194272} /* (11, 9, 13) {real, imag} */,
  {32'h4096b9b8, 32'h40f70a42} /* (11, 9, 12) {real, imag} */,
  {32'hbf6ee286, 32'h3f256abe} /* (11, 9, 11) {real, imag} */,
  {32'hc036cd10, 32'h4039630e} /* (11, 9, 10) {real, imag} */,
  {32'h4018f16a, 32'hbf811bb1} /* (11, 9, 9) {real, imag} */,
  {32'h3fe5e810, 32'hbfa9bd28} /* (11, 9, 8) {real, imag} */,
  {32'hbf872e1c, 32'h3fc5aa2f} /* (11, 9, 7) {real, imag} */,
  {32'hbff38279, 32'hbfde0a83} /* (11, 9, 6) {real, imag} */,
  {32'h40171630, 32'hc03901c6} /* (11, 9, 5) {real, imag} */,
  {32'hbff7bcf2, 32'h3f3f291c} /* (11, 9, 4) {real, imag} */,
  {32'h408ba5bd, 32'h40dbb1c3} /* (11, 9, 3) {real, imag} */,
  {32'hc04843a2, 32'hc04376c0} /* (11, 9, 2) {real, imag} */,
  {32'hc06d3ae0, 32'h3eff1d50} /* (11, 9, 1) {real, imag} */,
  {32'h3f832d34, 32'hc0c11ae2} /* (11, 9, 0) {real, imag} */,
  {32'h40619adc, 32'hc0e42176} /* (11, 8, 15) {real, imag} */,
  {32'hc0bb46aa, 32'h40516767} /* (11, 8, 14) {real, imag} */,
  {32'h4081f364, 32'hbfa440c9} /* (11, 8, 13) {real, imag} */,
  {32'hbfc6b82e, 32'h401a3e8d} /* (11, 8, 12) {real, imag} */,
  {32'h3a383000, 32'h3fdb0aaf} /* (11, 8, 11) {real, imag} */,
  {32'hbf5ea368, 32'hbd1f8f90} /* (11, 8, 10) {real, imag} */,
  {32'h3fe6befa, 32'h3f473b83} /* (11, 8, 9) {real, imag} */,
  {32'h3c4e7000, 32'hbf615734} /* (11, 8, 8) {real, imag} */,
  {32'hbfd97ee4, 32'hc0033b2d} /* (11, 8, 7) {real, imag} */,
  {32'hbfd554a8, 32'h3fb3d2e0} /* (11, 8, 6) {real, imag} */,
  {32'h4097d226, 32'h401eae8c} /* (11, 8, 5) {real, imag} */,
  {32'h40dce478, 32'hbe59b250} /* (11, 8, 4) {real, imag} */,
  {32'h40db2676, 32'hc0922cac} /* (11, 8, 3) {real, imag} */,
  {32'h404122fd, 32'h3f8514de} /* (11, 8, 2) {real, imag} */,
  {32'hbfc590c7, 32'h4135929b} /* (11, 8, 1) {real, imag} */,
  {32'hc0b22f8f, 32'hc0cd3830} /* (11, 8, 0) {real, imag} */,
  {32'h411dd7fc, 32'h40f259de} /* (11, 7, 15) {real, imag} */,
  {32'hc113786e, 32'hc03f04d4} /* (11, 7, 14) {real, imag} */,
  {32'hbf01cd1f, 32'h3fc8e938} /* (11, 7, 13) {real, imag} */,
  {32'h3ed359e4, 32'hc01ee6b0} /* (11, 7, 12) {real, imag} */,
  {32'hc043bbfa, 32'h3f9a0c02} /* (11, 7, 11) {real, imag} */,
  {32'h3fa3fe6e, 32'hbfc54cfb} /* (11, 7, 10) {real, imag} */,
  {32'hc017bdab, 32'h3f0ebfe4} /* (11, 7, 9) {real, imag} */,
  {32'hbf9d276b, 32'h403a126e} /* (11, 7, 8) {real, imag} */,
  {32'h3f5d7894, 32'h3f70d1a4} /* (11, 7, 7) {real, imag} */,
  {32'h3f24153c, 32'h40541c94} /* (11, 7, 6) {real, imag} */,
  {32'hbf5a2250, 32'hc021e932} /* (11, 7, 5) {real, imag} */,
  {32'hc0358b22, 32'hc0f48222} /* (11, 7, 4) {real, imag} */,
  {32'h400319d2, 32'h40bd1ee4} /* (11, 7, 3) {real, imag} */,
  {32'h402b2b61, 32'h3ff8f6dd} /* (11, 7, 2) {real, imag} */,
  {32'h3fd1589c, 32'h40483d2c} /* (11, 7, 1) {real, imag} */,
  {32'h3eef98ec, 32'hc1015bfc} /* (11, 7, 0) {real, imag} */,
  {32'hbf6db4b8, 32'hc187c5a4} /* (11, 6, 15) {real, imag} */,
  {32'h40609eb9, 32'hc0ae53b4} /* (11, 6, 14) {real, imag} */,
  {32'h3fd6717f, 32'hc11e66e6} /* (11, 6, 13) {real, imag} */,
  {32'h40b0d5d2, 32'h4094a086} /* (11, 6, 12) {real, imag} */,
  {32'h40802761, 32'h41034da2} /* (11, 6, 11) {real, imag} */,
  {32'hc0331107, 32'hbfb61b4a} /* (11, 6, 10) {real, imag} */,
  {32'h3ec66ec4, 32'h3fc0e2c6} /* (11, 6, 9) {real, imag} */,
  {32'h3dfadd00, 32'hbfcc49f6} /* (11, 6, 8) {real, imag} */,
  {32'hbfd6e431, 32'h3f67ccf4} /* (11, 6, 7) {real, imag} */,
  {32'h3f869436, 32'h3e6d8f8c} /* (11, 6, 6) {real, imag} */,
  {32'h409f88a7, 32'hc028a3d6} /* (11, 6, 5) {real, imag} */,
  {32'hc04e1a8d, 32'hc076c845} /* (11, 6, 4) {real, imag} */,
  {32'h4083d7c8, 32'hc0d2f894} /* (11, 6, 3) {real, imag} */,
  {32'h408d9132, 32'hc1169927} /* (11, 6, 2) {real, imag} */,
  {32'hc0ef5369, 32'hc0be0670} /* (11, 6, 1) {real, imag} */,
  {32'hc131abd6, 32'h40e58eb6} /* (11, 6, 0) {real, imag} */,
  {32'h403ce8ab, 32'hc10d3299} /* (11, 5, 15) {real, imag} */,
  {32'hc05697dd, 32'h41e77b99} /* (11, 5, 14) {real, imag} */,
  {32'h3f88ebc3, 32'hc1310452} /* (11, 5, 13) {real, imag} */,
  {32'h3fa36e9c, 32'hc0af0a34} /* (11, 5, 12) {real, imag} */,
  {32'h40eeb1c6, 32'h40683932} /* (11, 5, 11) {real, imag} */,
  {32'hc0d7cd2c, 32'hbf1fb718} /* (11, 5, 10) {real, imag} */,
  {32'hbecf2478, 32'h407aa596} /* (11, 5, 9) {real, imag} */,
  {32'hc031d19b, 32'h3ff04d3e} /* (11, 5, 8) {real, imag} */,
  {32'h3f97d591, 32'h40607956} /* (11, 5, 7) {real, imag} */,
  {32'h3ead8150, 32'hbee09b90} /* (11, 5, 6) {real, imag} */,
  {32'hbfcda008, 32'hc09d8ce1} /* (11, 5, 5) {real, imag} */,
  {32'hc0a15dca, 32'hc10fd5ef} /* (11, 5, 4) {real, imag} */,
  {32'hbf686e7a, 32'hc0268a6a} /* (11, 5, 3) {real, imag} */,
  {32'hc12faf87, 32'h416b5dee} /* (11, 5, 2) {real, imag} */,
  {32'h3fd5e242, 32'hc0d94058} /* (11, 5, 1) {real, imag} */,
  {32'h4127b3ee, 32'h40efb456} /* (11, 5, 0) {real, imag} */,
  {32'hc10b8888, 32'h40130dc6} /* (11, 4, 15) {real, imag} */,
  {32'hc1a97e67, 32'h3fcd6224} /* (11, 4, 14) {real, imag} */,
  {32'h408d16ef, 32'hc0f22bf1} /* (11, 4, 13) {real, imag} */,
  {32'hc08422e6, 32'h40cb14bc} /* (11, 4, 12) {real, imag} */,
  {32'hc10ed4ec, 32'hc134b198} /* (11, 4, 11) {real, imag} */,
  {32'h40c6700e, 32'h4102db9c} /* (11, 4, 10) {real, imag} */,
  {32'hc08afbec, 32'h409d5916} /* (11, 4, 9) {real, imag} */,
  {32'h401bc6bc, 32'hc0a26b7c} /* (11, 4, 8) {real, imag} */,
  {32'hc0d4e9d2, 32'hc0327698} /* (11, 4, 7) {real, imag} */,
  {32'h3fffadd8, 32'hc106bb20} /* (11, 4, 6) {real, imag} */,
  {32'hc00158be, 32'h410635e0} /* (11, 4, 5) {real, imag} */,
  {32'h41272e8b, 32'hbe800e10} /* (11, 4, 4) {real, imag} */,
  {32'h4093d191, 32'hc10a8c8c} /* (11, 4, 3) {real, imag} */,
  {32'h41a62a77, 32'h413a92c8} /* (11, 4, 2) {real, imag} */,
  {32'h4061df5a, 32'h3ff2cbeb} /* (11, 4, 1) {real, imag} */,
  {32'h414b867d, 32'hc106781c} /* (11, 4, 0) {real, imag} */,
  {32'hc0d5c1aa, 32'hbfe8f314} /* (11, 3, 15) {real, imag} */,
  {32'h419d5b8f, 32'h41e214b3} /* (11, 3, 14) {real, imag} */,
  {32'h40de663a, 32'hc153d80e} /* (11, 3, 13) {real, imag} */,
  {32'hc03d32bf, 32'h4157690e} /* (11, 3, 12) {real, imag} */,
  {32'h40e18266, 32'hc106126e} /* (11, 3, 11) {real, imag} */,
  {32'hc11f2b3c, 32'hbfeb4fa4} /* (11, 3, 10) {real, imag} */,
  {32'hbebe6bd0, 32'h3f2b1f12} /* (11, 3, 9) {real, imag} */,
  {32'h3f4a7c04, 32'hbf1eec2c} /* (11, 3, 8) {real, imag} */,
  {32'h3fbd4e28, 32'hc037217e} /* (11, 3, 7) {real, imag} */,
  {32'hc0244db6, 32'h4094d651} /* (11, 3, 6) {real, imag} */,
  {32'h415a5e27, 32'hc09f8094} /* (11, 3, 5) {real, imag} */,
  {32'h40bf5648, 32'h412d6c92} /* (11, 3, 4) {real, imag} */,
  {32'h40ee78bc, 32'h414fe35a} /* (11, 3, 3) {real, imag} */,
  {32'hc15f1702, 32'h40e63d9c} /* (11, 3, 2) {real, imag} */,
  {32'h412d3f6b, 32'hc1438168} /* (11, 3, 1) {real, imag} */,
  {32'hc0c5156e, 32'hc03f245d} /* (11, 3, 0) {real, imag} */,
  {32'h417539d2, 32'h40ae25c0} /* (11, 2, 15) {real, imag} */,
  {32'h4018aa02, 32'hc19cc161} /* (11, 2, 14) {real, imag} */,
  {32'hc1922c3b, 32'h41df0975} /* (11, 2, 13) {real, imag} */,
  {32'hc00043ac, 32'hc15c302f} /* (11, 2, 12) {real, imag} */,
  {32'h41286d96, 32'hc18b1232} /* (11, 2, 11) {real, imag} */,
  {32'h4183341f, 32'hc1132570} /* (11, 2, 10) {real, imag} */,
  {32'hbfa0e9c0, 32'h4080d47c} /* (11, 2, 9) {real, imag} */,
  {32'h40c02e46, 32'h4010f702} /* (11, 2, 8) {real, imag} */,
  {32'h413cfa52, 32'hc188fa2c} /* (11, 2, 7) {real, imag} */,
  {32'hc151cf36, 32'h40d90da8} /* (11, 2, 6) {real, imag} */,
  {32'hbffc74dc, 32'hc0a98b6e} /* (11, 2, 5) {real, imag} */,
  {32'h409a6d38, 32'hc19c6b26} /* (11, 2, 4) {real, imag} */,
  {32'hc1410518, 32'h41b821c7} /* (11, 2, 3) {real, imag} */,
  {32'hc1830cec, 32'h41623a4a} /* (11, 2, 2) {real, imag} */,
  {32'h3ff52c20, 32'h4191431f} /* (11, 2, 1) {real, imag} */,
  {32'hbfd31e78, 32'hc16587b0} /* (11, 2, 0) {real, imag} */,
  {32'h41a57cbf, 32'hc0b17f2e} /* (11, 1, 15) {real, imag} */,
  {32'h41c1c459, 32'h4049767a} /* (11, 1, 14) {real, imag} */,
  {32'hc09bbdf8, 32'h416dbf20} /* (11, 1, 13) {real, imag} */,
  {32'h41a121a3, 32'hc18b8dfa} /* (11, 1, 12) {real, imag} */,
  {32'hbf01ad60, 32'h4130be14} /* (11, 1, 11) {real, imag} */,
  {32'hc02bafa0, 32'hc00c922e} /* (11, 1, 10) {real, imag} */,
  {32'h4006303c, 32'hc066e28e} /* (11, 1, 9) {real, imag} */,
  {32'hbeffd970, 32'h3fe3493c} /* (11, 1, 8) {real, imag} */,
  {32'h40966f60, 32'h3fd5aadc} /* (11, 1, 7) {real, imag} */,
  {32'h41b23b8f, 32'h40650d1a} /* (11, 1, 6) {real, imag} */,
  {32'hc1c27f75, 32'hc1562e2c} /* (11, 1, 5) {real, imag} */,
  {32'h3ff1f930, 32'h407a0f5e} /* (11, 1, 4) {real, imag} */,
  {32'h41207495, 32'h40bdd28f} /* (11, 1, 3) {real, imag} */,
  {32'hc0816428, 32'h3fcc92d7} /* (11, 1, 2) {real, imag} */,
  {32'h41335302, 32'h418f2f24} /* (11, 1, 1) {real, imag} */,
  {32'h4147a58c, 32'h41028a20} /* (11, 1, 0) {real, imag} */,
  {32'h40f9db14, 32'h40551a44} /* (11, 0, 15) {real, imag} */,
  {32'hc1928d1e, 32'hbdcd46c0} /* (11, 0, 14) {real, imag} */,
  {32'hc127fd62, 32'h4133bdd9} /* (11, 0, 13) {real, imag} */,
  {32'h410a1875, 32'h41dc13c9} /* (11, 0, 12) {real, imag} */,
  {32'hc0d37655, 32'hc12707a8} /* (11, 0, 11) {real, imag} */,
  {32'h40c90ec8, 32'h40f4778a} /* (11, 0, 10) {real, imag} */,
  {32'hc0dc02e0, 32'h40147b0c} /* (11, 0, 9) {real, imag} */,
  {32'hc02470b4, 32'h3d8bc300} /* (11, 0, 8) {real, imag} */,
  {32'h407a0841, 32'h41063a8f} /* (11, 0, 7) {real, imag} */,
  {32'hbf9590e0, 32'h40f235e6} /* (11, 0, 6) {real, imag} */,
  {32'hc03bc31a, 32'h41eed974} /* (11, 0, 5) {real, imag} */,
  {32'h41592801, 32'h40ac52ec} /* (11, 0, 4) {real, imag} */,
  {32'hc11800b6, 32'hc10a337d} /* (11, 0, 3) {real, imag} */,
  {32'hc18347f2, 32'hc0f4c7b5} /* (11, 0, 2) {real, imag} */,
  {32'hc1551ea2, 32'hc190ae64} /* (11, 0, 1) {real, imag} */,
  {32'h41eb0f90, 32'h421d4f90} /* (11, 0, 0) {real, imag} */,
  {32'h41012070, 32'h410a3ac0} /* (10, 15, 15) {real, imag} */,
  {32'hc0d79028, 32'hc029f6ea} /* (10, 15, 14) {real, imag} */,
  {32'h40622464, 32'hc20572c7} /* (10, 15, 13) {real, imag} */,
  {32'h3fc2e7d8, 32'h4056b0d8} /* (10, 15, 12) {real, imag} */,
  {32'h40ab53c8, 32'hc139cfe4} /* (10, 15, 11) {real, imag} */,
  {32'h4151b8e3, 32'hc0939b26} /* (10, 15, 10) {real, imag} */,
  {32'hbf9c4938, 32'hbff21d4a} /* (10, 15, 9) {real, imag} */,
  {32'hc0253858, 32'h40521d28} /* (10, 15, 8) {real, imag} */,
  {32'h405cb852, 32'hc063fad5} /* (10, 15, 7) {real, imag} */,
  {32'hc0ae8f12, 32'h40de64d2} /* (10, 15, 6) {real, imag} */,
  {32'hc05e8e0d, 32'hc08fb771} /* (10, 15, 5) {real, imag} */,
  {32'h41a6063c, 32'hc1bde7db} /* (10, 15, 4) {real, imag} */,
  {32'hc1671223, 32'hc1a8e071} /* (10, 15, 3) {real, imag} */,
  {32'hc1ef4cf2, 32'hc07a52ec} /* (10, 15, 2) {real, imag} */,
  {32'hc13c7ea6, 32'hc1232252} /* (10, 15, 1) {real, imag} */,
  {32'h42015d2e, 32'h410420ce} /* (10, 15, 0) {real, imag} */,
  {32'hc23f251e, 32'hc11f54fb} /* (10, 14, 15) {real, imag} */,
  {32'hc0bc8a24, 32'hc0c99808} /* (10, 14, 14) {real, imag} */,
  {32'h4175949b, 32'h40885af4} /* (10, 14, 13) {real, imag} */,
  {32'hc108e3c6, 32'h41b51e84} /* (10, 14, 12) {real, imag} */,
  {32'h413c3ff0, 32'hc133f540} /* (10, 14, 11) {real, imag} */,
  {32'hbf9653c0, 32'h400ae8fb} /* (10, 14, 10) {real, imag} */,
  {32'h4094e1b5, 32'hc01009e2} /* (10, 14, 9) {real, imag} */,
  {32'h3fdc5610, 32'hc00fd300} /* (10, 14, 8) {real, imag} */,
  {32'hc00a028e, 32'hbe7f8058} /* (10, 14, 7) {real, imag} */,
  {32'h4013b0ec, 32'h4074010f} /* (10, 14, 6) {real, imag} */,
  {32'hc0f92f40, 32'h3f94e0f0} /* (10, 14, 5) {real, imag} */,
  {32'h3fe9475c, 32'hc14c665f} /* (10, 14, 4) {real, imag} */,
  {32'h4112a18b, 32'hbf515188} /* (10, 14, 3) {real, imag} */,
  {32'hc1ba6f15, 32'h40496143} /* (10, 14, 2) {real, imag} */,
  {32'h41ab9919, 32'hc185589c} /* (10, 14, 1) {real, imag} */,
  {32'h41de3027, 32'hc1a82527} /* (10, 14, 0) {real, imag} */,
  {32'hbfd78bfa, 32'h414c31a0} /* (10, 13, 15) {real, imag} */,
  {32'h3fb045a4, 32'hc1494e8e} /* (10, 13, 14) {real, imag} */,
  {32'hc1443bd8, 32'hc0f7fab7} /* (10, 13, 13) {real, imag} */,
  {32'h4104ef34, 32'hc0b40414} /* (10, 13, 12) {real, imag} */,
  {32'h3ffda861, 32'hc01bd498} /* (10, 13, 11) {real, imag} */,
  {32'hc094e50a, 32'h3e590380} /* (10, 13, 10) {real, imag} */,
  {32'h404b2912, 32'hc02f2578} /* (10, 13, 9) {real, imag} */,
  {32'hbf2a9be7, 32'hc00558d0} /* (10, 13, 8) {real, imag} */,
  {32'hbf895419, 32'hc0481b98} /* (10, 13, 7) {real, imag} */,
  {32'hbfe79c5a, 32'hc0220f96} /* (10, 13, 6) {real, imag} */,
  {32'h3f88b9e1, 32'h405ba004} /* (10, 13, 5) {real, imag} */,
  {32'h41092080, 32'hc05b7fb5} /* (10, 13, 4) {real, imag} */,
  {32'h40cbff00, 32'hc19210b2} /* (10, 13, 3) {real, imag} */,
  {32'hbecd5f80, 32'hc00327e0} /* (10, 13, 2) {real, imag} */,
  {32'hc1044736, 32'h40bad9e8} /* (10, 13, 1) {real, imag} */,
  {32'hbdde5f48, 32'h419e6910} /* (10, 13, 0) {real, imag} */,
  {32'h4150f488, 32'hc0678b54} /* (10, 12, 15) {real, imag} */,
  {32'h4174dca6, 32'hc1675579} /* (10, 12, 14) {real, imag} */,
  {32'hc06abf9f, 32'h40c2b944} /* (10, 12, 13) {real, imag} */,
  {32'hc189c87e, 32'h3f5b8f48} /* (10, 12, 12) {real, imag} */,
  {32'h3febed7f, 32'h3fdeb84e} /* (10, 12, 11) {real, imag} */,
  {32'h4062ea50, 32'hbff74b08} /* (10, 12, 10) {real, imag} */,
  {32'hc027bca0, 32'h3ffe8ccc} /* (10, 12, 9) {real, imag} */,
  {32'h3f219ee8, 32'h40e04612} /* (10, 12, 8) {real, imag} */,
  {32'h3e212980, 32'h4039255e} /* (10, 12, 7) {real, imag} */,
  {32'hc0bbf46a, 32'hbfb32d68} /* (10, 12, 6) {real, imag} */,
  {32'hc06c2516, 32'hbeb96218} /* (10, 12, 5) {real, imag} */,
  {32'h40963faf, 32'hbf6e8138} /* (10, 12, 4) {real, imag} */,
  {32'hc044d245, 32'hbfcfaabe} /* (10, 12, 3) {real, imag} */,
  {32'hc169c612, 32'hc0b637fa} /* (10, 12, 2) {real, imag} */,
  {32'h41694776, 32'h41643f6d} /* (10, 12, 1) {real, imag} */,
  {32'hc122826a, 32'hc0ff0d34} /* (10, 12, 0) {real, imag} */,
  {32'h41541f8a, 32'hbee87610} /* (10, 11, 15) {real, imag} */,
  {32'hbf4fea7e, 32'h41866600} /* (10, 11, 14) {real, imag} */,
  {32'h41262032, 32'h40e575c8} /* (10, 11, 13) {real, imag} */,
  {32'hc10a51e3, 32'hc02018d6} /* (10, 11, 12) {real, imag} */,
  {32'h3e3e33e8, 32'hc11451c0} /* (10, 11, 11) {real, imag} */,
  {32'hc08892ba, 32'hc02f6838} /* (10, 11, 10) {real, imag} */,
  {32'hc063f96f, 32'h40ab168a} /* (10, 11, 9) {real, imag} */,
  {32'hbff54976, 32'hc000cee4} /* (10, 11, 8) {real, imag} */,
  {32'hbfab091e, 32'h3ff75101} /* (10, 11, 7) {real, imag} */,
  {32'h3fe26090, 32'hbfae5ee1} /* (10, 11, 6) {real, imag} */,
  {32'h3fc36e9d, 32'hbf3df0f8} /* (10, 11, 5) {real, imag} */,
  {32'hc03f76a5, 32'h4110e6f2} /* (10, 11, 4) {real, imag} */,
  {32'hbf947890, 32'hc18b05ea} /* (10, 11, 3) {real, imag} */,
  {32'h3f6a0e3e, 32'h41168ef7} /* (10, 11, 2) {real, imag} */,
  {32'h3f688a80, 32'h3f7eebec} /* (10, 11, 1) {real, imag} */,
  {32'h4096a548, 32'hc150c93f} /* (10, 11, 0) {real, imag} */,
  {32'h408af368, 32'h40894f6f} /* (10, 10, 15) {real, imag} */,
  {32'h41053587, 32'h40f27f70} /* (10, 10, 14) {real, imag} */,
  {32'hbe85ccc4, 32'hbf45a926} /* (10, 10, 13) {real, imag} */,
  {32'hbfe6aed6, 32'hc0b872c1} /* (10, 10, 12) {real, imag} */,
  {32'h400528fe, 32'hbeafc518} /* (10, 10, 11) {real, imag} */,
  {32'h405b48d4, 32'hbfd71954} /* (10, 10, 10) {real, imag} */,
  {32'hbe733d98, 32'h3f83adfa} /* (10, 10, 9) {real, imag} */,
  {32'h3f208be8, 32'hbf7ddaa8} /* (10, 10, 8) {real, imag} */,
  {32'h4010f8b2, 32'hbf1e7fbc} /* (10, 10, 7) {real, imag} */,
  {32'h3fe39c34, 32'h4007db5c} /* (10, 10, 6) {real, imag} */,
  {32'hbf18ee32, 32'hc081ea6a} /* (10, 10, 5) {real, imag} */,
  {32'h409715fc, 32'hc0d2b00b} /* (10, 10, 4) {real, imag} */,
  {32'hc046bff6, 32'h3fdae669} /* (10, 10, 3) {real, imag} */,
  {32'hc0932572, 32'hc0075508} /* (10, 10, 2) {real, imag} */,
  {32'hc0b80b98, 32'h40e34cf9} /* (10, 10, 1) {real, imag} */,
  {32'hc1480b10, 32'h408e093d} /* (10, 10, 0) {real, imag} */,
  {32'hc0b34412, 32'hbe26b95c} /* (10, 9, 15) {real, imag} */,
  {32'hc097525a, 32'hc08930dc} /* (10, 9, 14) {real, imag} */,
  {32'hc0b0b691, 32'h3faf6eb0} /* (10, 9, 13) {real, imag} */,
  {32'hc028e89a, 32'hbfb6faa7} /* (10, 9, 12) {real, imag} */,
  {32'h3f9ec7fa, 32'h40c30988} /* (10, 9, 11) {real, imag} */,
  {32'h3fab3535, 32'hbf2116e5} /* (10, 9, 10) {real, imag} */,
  {32'hbe8a985c, 32'hbfa5129e} /* (10, 9, 9) {real, imag} */,
  {32'h400625ea, 32'h3fe0f512} /* (10, 9, 8) {real, imag} */,
  {32'hbfbf3f23, 32'h3f7260fc} /* (10, 9, 7) {real, imag} */,
  {32'hbfbc7c17, 32'hbf855e80} /* (10, 9, 6) {real, imag} */,
  {32'h3fbabb1a, 32'hc01e6314} /* (10, 9, 5) {real, imag} */,
  {32'h3e142158, 32'h400ec860} /* (10, 9, 4) {real, imag} */,
  {32'h40f09107, 32'h41155e55} /* (10, 9, 3) {real, imag} */,
  {32'hbf4312c0, 32'h3f741c94} /* (10, 9, 2) {real, imag} */,
  {32'hbf021920, 32'h3f98f58c} /* (10, 9, 1) {real, imag} */,
  {32'h40d7c4d7, 32'h3fffa2e4} /* (10, 9, 0) {real, imag} */,
  {32'h40d98366, 32'hbfdcdcaa} /* (10, 8, 15) {real, imag} */,
  {32'hc05fa027, 32'hc0d2683d} /* (10, 8, 14) {real, imag} */,
  {32'hbfe6658c, 32'h409fc4ea} /* (10, 8, 13) {real, imag} */,
  {32'h3f5c6b11, 32'hc02a9884} /* (10, 8, 12) {real, imag} */,
  {32'hc0158cc2, 32'h405ab94e} /* (10, 8, 11) {real, imag} */,
  {32'h40415a24, 32'hbf9bd30c} /* (10, 8, 10) {real, imag} */,
  {32'h3fa4de91, 32'hbf1b3e7c} /* (10, 8, 9) {real, imag} */,
  {32'hbe5e2440, 32'h3f0ff5fe} /* (10, 8, 8) {real, imag} */,
  {32'h3c958d40, 32'hbf8b7eb5} /* (10, 8, 7) {real, imag} */,
  {32'h3f322fb2, 32'h3fc85634} /* (10, 8, 6) {real, imag} */,
  {32'h40414102, 32'h3f5d089e} /* (10, 8, 5) {real, imag} */,
  {32'hbf7c780b, 32'h3fb1677b} /* (10, 8, 4) {real, imag} */,
  {32'h3cfef780, 32'hbfd0e2a6} /* (10, 8, 3) {real, imag} */,
  {32'h3fd705ea, 32'hc007a732} /* (10, 8, 2) {real, imag} */,
  {32'hc0825a96, 32'h3f2ef71b} /* (10, 8, 1) {real, imag} */,
  {32'h40333762, 32'hc083b770} /* (10, 8, 0) {real, imag} */,
  {32'h3fe23486, 32'hc07622fe} /* (10, 7, 15) {real, imag} */,
  {32'hc061770c, 32'h4107ca5a} /* (10, 7, 14) {real, imag} */,
  {32'h3e4e5c60, 32'hbf497b48} /* (10, 7, 13) {real, imag} */,
  {32'h3e55b6ec, 32'hc0da5915} /* (10, 7, 12) {real, imag} */,
  {32'hbfcc2e96, 32'hbf7378aa} /* (10, 7, 11) {real, imag} */,
  {32'hbdf65d08, 32'hbe070730} /* (10, 7, 10) {real, imag} */,
  {32'h3bf5bc80, 32'hbf064768} /* (10, 7, 9) {real, imag} */,
  {32'h3e832cd0, 32'h3f8aa0e8} /* (10, 7, 8) {real, imag} */,
  {32'hbf6b827f, 32'hbeb64d98} /* (10, 7, 7) {real, imag} */,
  {32'h3fb06352, 32'hc05950bb} /* (10, 7, 6) {real, imag} */,
  {32'h3fdd2842, 32'h3eb2086c} /* (10, 7, 5) {real, imag} */,
  {32'h3fdb75d8, 32'h3ff2acac} /* (10, 7, 4) {real, imag} */,
  {32'hc0b9450b, 32'h410eb300} /* (10, 7, 3) {real, imag} */,
  {32'h3f041cf2, 32'h3fc2b22c} /* (10, 7, 2) {real, imag} */,
  {32'hc0b87ea2, 32'hbff1b665} /* (10, 7, 1) {real, imag} */,
  {32'h40aa46af, 32'hc05ea30c} /* (10, 7, 0) {real, imag} */,
  {32'hc103ebea, 32'hbc9b76c0} /* (10, 6, 15) {real, imag} */,
  {32'hc0cf69c9, 32'h40514d7f} /* (10, 6, 14) {real, imag} */,
  {32'h4082e03a, 32'h40c486dc} /* (10, 6, 13) {real, imag} */,
  {32'hbf3a5780, 32'hc077eb39} /* (10, 6, 12) {real, imag} */,
  {32'hc0ea1a00, 32'hbf56296c} /* (10, 6, 11) {real, imag} */,
  {32'h3fc8f1cc, 32'hc06d8878} /* (10, 6, 10) {real, imag} */,
  {32'h4058766b, 32'hbf9308ff} /* (10, 6, 9) {real, imag} */,
  {32'hc00d6fe7, 32'hbfd1fb06} /* (10, 6, 8) {real, imag} */,
  {32'hbfe9e63a, 32'h4082171a} /* (10, 6, 7) {real, imag} */,
  {32'h409d6d1b, 32'hbee47e50} /* (10, 6, 6) {real, imag} */,
  {32'hc041f0c8, 32'h3eede658} /* (10, 6, 5) {real, imag} */,
  {32'h41623416, 32'h3ec569e8} /* (10, 6, 4) {real, imag} */,
  {32'hc0802df6, 32'hc07ebe59} /* (10, 6, 3) {real, imag} */,
  {32'hc13f308c, 32'h3fde054e} /* (10, 6, 2) {real, imag} */,
  {32'h40e0603c, 32'hbe8eea6c} /* (10, 6, 1) {real, imag} */,
  {32'hbfcd3152, 32'h401cb907} /* (10, 6, 0) {real, imag} */,
  {32'hbfe30d4f, 32'h411964be} /* (10, 5, 15) {real, imag} */,
  {32'hc000844f, 32'hc0a58ba9} /* (10, 5, 14) {real, imag} */,
  {32'hc14fb29e, 32'hbfb369d0} /* (10, 5, 13) {real, imag} */,
  {32'h403664da, 32'h4145e819} /* (10, 5, 12) {real, imag} */,
  {32'hc014f1ef, 32'hc073eb16} /* (10, 5, 11) {real, imag} */,
  {32'hbfc8c18e, 32'hc0be596d} /* (10, 5, 10) {real, imag} */,
  {32'h40118272, 32'h40caf874} /* (10, 5, 9) {real, imag} */,
  {32'hbfd97fba, 32'hc02342d1} /* (10, 5, 8) {real, imag} */,
  {32'hbfc3e00d, 32'h3f8dbfc2} /* (10, 5, 7) {real, imag} */,
  {32'hc07c30eb, 32'h40127a0a} /* (10, 5, 6) {real, imag} */,
  {32'h408f4326, 32'hc0379946} /* (10, 5, 5) {real, imag} */,
  {32'hbfa848c8, 32'hc0903e1e} /* (10, 5, 4) {real, imag} */,
  {32'hc094ea1d, 32'hc1027d81} /* (10, 5, 3) {real, imag} */,
  {32'hc09625fe, 32'hbf82e04c} /* (10, 5, 2) {real, imag} */,
  {32'h3fe41ac1, 32'hc09cb758} /* (10, 5, 1) {real, imag} */,
  {32'h410f7f01, 32'hc0eca824} /* (10, 5, 0) {real, imag} */,
  {32'hc1bc1522, 32'h40fbab94} /* (10, 4, 15) {real, imag} */,
  {32'h4019392a, 32'hc12b76c7} /* (10, 4, 14) {real, imag} */,
  {32'hc1b3a10e, 32'h41289ddd} /* (10, 4, 13) {real, imag} */,
  {32'h4112059c, 32'h41398500} /* (10, 4, 12) {real, imag} */,
  {32'hbede6e08, 32'h4066404c} /* (10, 4, 11) {real, imag} */,
  {32'h4019cfc1, 32'hbe1cb5b0} /* (10, 4, 10) {real, imag} */,
  {32'hc06cfea4, 32'hc06778fc} /* (10, 4, 9) {real, imag} */,
  {32'h40828cb3, 32'h3fdbd5f8} /* (10, 4, 8) {real, imag} */,
  {32'h3fe501b8, 32'hc019403c} /* (10, 4, 7) {real, imag} */,
  {32'hc044e00b, 32'h40dcd992} /* (10, 4, 6) {real, imag} */,
  {32'h40d86718, 32'hc15d3c77} /* (10, 4, 5) {real, imag} */,
  {32'hbf303d20, 32'h411c9fd0} /* (10, 4, 4) {real, imag} */,
  {32'hc1236317, 32'h4099f366} /* (10, 4, 3) {real, imag} */,
  {32'h3fac666f, 32'hbecf99a0} /* (10, 4, 2) {real, imag} */,
  {32'hbfebc1d8, 32'h4141fc76} /* (10, 4, 1) {real, imag} */,
  {32'h410f895e, 32'hc186b870} /* (10, 4, 0) {real, imag} */,
  {32'h415ffe46, 32'h4027d9ac} /* (10, 3, 15) {real, imag} */,
  {32'h41846a80, 32'h41674e15} /* (10, 3, 14) {real, imag} */,
  {32'h40e3ee26, 32'hc0d17a48} /* (10, 3, 13) {real, imag} */,
  {32'hbfebcf52, 32'h41897145} /* (10, 3, 12) {real, imag} */,
  {32'h3fe30ccc, 32'h403dab8c} /* (10, 3, 11) {real, imag} */,
  {32'h403acec6, 32'h40acbcdf} /* (10, 3, 10) {real, imag} */,
  {32'hc05f7a56, 32'hbfa6c068} /* (10, 3, 9) {real, imag} */,
  {32'h3e08e3c0, 32'hbf47f2a0} /* (10, 3, 8) {real, imag} */,
  {32'h3f6e2898, 32'hc060774c} /* (10, 3, 7) {real, imag} */,
  {32'h40221422, 32'h403a9c5a} /* (10, 3, 6) {real, imag} */,
  {32'h418a2b6b, 32'hc00a43ac} /* (10, 3, 5) {real, imag} */,
  {32'hc0ca9d94, 32'hc08d3221} /* (10, 3, 4) {real, imag} */,
  {32'hc0c35aec, 32'hc19cdb18} /* (10, 3, 3) {real, imag} */,
  {32'hc0bbf0fa, 32'hc104468b} /* (10, 3, 2) {real, imag} */,
  {32'h41a90053, 32'h4117ad65} /* (10, 3, 1) {real, imag} */,
  {32'hc188372c, 32'h419b2bab} /* (10, 3, 0) {real, imag} */,
  {32'h41818f70, 32'hc09714b2} /* (10, 2, 15) {real, imag} */,
  {32'hc0090f26, 32'hc0b612ae} /* (10, 2, 14) {real, imag} */,
  {32'h40fc57e6, 32'h3f167a00} /* (10, 2, 13) {real, imag} */,
  {32'h413bd2b0, 32'h412eb786} /* (10, 2, 12) {real, imag} */,
  {32'hc0650ba8, 32'hc0a33fd8} /* (10, 2, 11) {real, imag} */,
  {32'hbff3a8d4, 32'h410f8e29} /* (10, 2, 10) {real, imag} */,
  {32'hc0f13811, 32'h3ddebf80} /* (10, 2, 9) {real, imag} */,
  {32'h40fe3890, 32'h40164204} /* (10, 2, 8) {real, imag} */,
  {32'h40129d2a, 32'hc07c4f68} /* (10, 2, 7) {real, imag} */,
  {32'hc0d1e7af, 32'hbedc98e0} /* (10, 2, 6) {real, imag} */,
  {32'hc1345d14, 32'hc07225e8} /* (10, 2, 5) {real, imag} */,
  {32'h408cb911, 32'hc10f02c2} /* (10, 2, 4) {real, imag} */,
  {32'hbf773770, 32'h410c1db0} /* (10, 2, 3) {real, imag} */,
  {32'hc0efe241, 32'h41add86a} /* (10, 2, 2) {real, imag} */,
  {32'hc100b01c, 32'hc10428ee} /* (10, 2, 1) {real, imag} */,
  {32'h40b53228, 32'hc0f52cbc} /* (10, 2, 0) {real, imag} */,
  {32'h41cd9f92, 32'h403ae78a} /* (10, 1, 15) {real, imag} */,
  {32'h400a2a78, 32'hc1da7942} /* (10, 1, 14) {real, imag} */,
  {32'h3f1206a0, 32'h41041f2a} /* (10, 1, 13) {real, imag} */,
  {32'hc0bfa5b7, 32'h4061ab24} /* (10, 1, 12) {real, imag} */,
  {32'h3ffb551c, 32'hc05e5bc8} /* (10, 1, 11) {real, imag} */,
  {32'h408c355b, 32'h3f132fbe} /* (10, 1, 10) {real, imag} */,
  {32'h416edd7f, 32'hbfc4747e} /* (10, 1, 9) {real, imag} */,
  {32'hbfc4b558, 32'h4067f470} /* (10, 1, 8) {real, imag} */,
  {32'h405373d4, 32'h40d66806} /* (10, 1, 7) {real, imag} */,
  {32'hbf7bcf58, 32'hbf52e09e} /* (10, 1, 6) {real, imag} */,
  {32'h403c1d90, 32'h40a0f5ba} /* (10, 1, 5) {real, imag} */,
  {32'hc0af07ed, 32'h3ecb3d60} /* (10, 1, 4) {real, imag} */,
  {32'hc17c6462, 32'hc186d76f} /* (10, 1, 3) {real, imag} */,
  {32'h41a86fb9, 32'hc1a12d4e} /* (10, 1, 2) {real, imag} */,
  {32'hc0bddb56, 32'h40aadc87} /* (10, 1, 1) {real, imag} */,
  {32'hc1ff0e1e, 32'hc1867730} /* (10, 1, 0) {real, imag} */,
  {32'h40377f9b, 32'h4108968e} /* (10, 0, 15) {real, imag} */,
  {32'hc1d779ef, 32'h418f715e} /* (10, 0, 14) {real, imag} */,
  {32'hc0e3a5ce, 32'hc010d590} /* (10, 0, 13) {real, imag} */,
  {32'h4099b06f, 32'hc05856da} /* (10, 0, 12) {real, imag} */,
  {32'hc113954b, 32'h3f9fa0ea} /* (10, 0, 11) {real, imag} */,
  {32'hc0a0bc9a, 32'hc01a59bc} /* (10, 0, 10) {real, imag} */,
  {32'hc01110cd, 32'hbfb4a0ef} /* (10, 0, 9) {real, imag} */,
  {32'hc063a188, 32'h40354954} /* (10, 0, 8) {real, imag} */,
  {32'hbf0cac6c, 32'hbfe03491} /* (10, 0, 7) {real, imag} */,
  {32'h40dfc94e, 32'hbf7eb872} /* (10, 0, 6) {real, imag} */,
  {32'hc0d74ade, 32'hc0096aad} /* (10, 0, 5) {real, imag} */,
  {32'hc14b4386, 32'h41420c38} /* (10, 0, 4) {real, imag} */,
  {32'hc0ed6d86, 32'h4167cb4a} /* (10, 0, 3) {real, imag} */,
  {32'h41f272fb, 32'hc0d97dde} /* (10, 0, 2) {real, imag} */,
  {32'h412472e6, 32'h417241d2} /* (10, 0, 1) {real, imag} */,
  {32'h401f39a4, 32'hc0de6032} /* (10, 0, 0) {real, imag} */,
  {32'h41c84b0e, 32'hc1066ae1} /* (9, 15, 15) {real, imag} */,
  {32'h3f9d8f2a, 32'hbf1a564d} /* (9, 15, 14) {real, imag} */,
  {32'hc166f3c7, 32'h40b5324a} /* (9, 15, 13) {real, imag} */,
  {32'h3fd4aaa2, 32'hc16374ae} /* (9, 15, 12) {real, imag} */,
  {32'h41478243, 32'hc145fd3f} /* (9, 15, 11) {real, imag} */,
  {32'hc10d11ab, 32'hbfe21e1c} /* (9, 15, 10) {real, imag} */,
  {32'h3ee83dc0, 32'hc07ffa3b} /* (9, 15, 9) {real, imag} */,
  {32'h4009f253, 32'hc0514186} /* (9, 15, 8) {real, imag} */,
  {32'hbf2c8a40, 32'hc03c5fc1} /* (9, 15, 7) {real, imag} */,
  {32'h3fa5ec2e, 32'hbfc3b974} /* (9, 15, 6) {real, imag} */,
  {32'hc1156487, 32'h3fd625c8} /* (9, 15, 5) {real, imag} */,
  {32'hc0a26ebc, 32'h40b2fe9d} /* (9, 15, 4) {real, imag} */,
  {32'hc140f871, 32'hc06ab66d} /* (9, 15, 3) {real, imag} */,
  {32'h3fd1ce12, 32'hbfe60016} /* (9, 15, 2) {real, imag} */,
  {32'hc0534c38, 32'h4073eeb4} /* (9, 15, 1) {real, imag} */,
  {32'hbfc1255a, 32'h41419d94} /* (9, 15, 0) {real, imag} */,
  {32'h40f76c50, 32'h41495d85} /* (9, 14, 15) {real, imag} */,
  {32'hc18daf9b, 32'hc111b10a} /* (9, 14, 14) {real, imag} */,
  {32'hc0590458, 32'hbdced5c0} /* (9, 14, 13) {real, imag} */,
  {32'h3faff662, 32'h406ed3b2} /* (9, 14, 12) {real, imag} */,
  {32'hc11e22e6, 32'h40601c74} /* (9, 14, 11) {real, imag} */,
  {32'h4104517e, 32'h408bdda9} /* (9, 14, 10) {real, imag} */,
  {32'h3fda8b61, 32'hbf2fddec} /* (9, 14, 9) {real, imag} */,
  {32'h3fb35e34, 32'h4026a2c8} /* (9, 14, 8) {real, imag} */,
  {32'hc013fb8c, 32'hc0337f4b} /* (9, 14, 7) {real, imag} */,
  {32'h401c6553, 32'h3e799820} /* (9, 14, 6) {real, imag} */,
  {32'h410ff534, 32'h3f613ec0} /* (9, 14, 5) {real, imag} */,
  {32'hbf83da8a, 32'h410da558} /* (9, 14, 4) {real, imag} */,
  {32'h40ca2abc, 32'h40dd51a3} /* (9, 14, 3) {real, imag} */,
  {32'h406bbfba, 32'hbf055598} /* (9, 14, 2) {real, imag} */,
  {32'hc0209ccc, 32'hc0f13b9a} /* (9, 14, 1) {real, imag} */,
  {32'hc0b68235, 32'hc064f6d2} /* (9, 14, 0) {real, imag} */,
  {32'h40fcd9db, 32'h406505e6} /* (9, 13, 15) {real, imag} */,
  {32'hc093e20e, 32'h3f9e8250} /* (9, 13, 14) {real, imag} */,
  {32'h3fe1616e, 32'h40984574} /* (9, 13, 13) {real, imag} */,
  {32'h4108132c, 32'h3ff1a738} /* (9, 13, 12) {real, imag} */,
  {32'hbf247552, 32'h3f8aa4fc} /* (9, 13, 11) {real, imag} */,
  {32'hc08e6610, 32'hbf60b1b6} /* (9, 13, 10) {real, imag} */,
  {32'h3f5592b6, 32'hbfaaac62} /* (9, 13, 9) {real, imag} */,
  {32'h3f22ed78, 32'h3f5dcd98} /* (9, 13, 8) {real, imag} */,
  {32'h3f74c8b6, 32'h408a7cba} /* (9, 13, 7) {real, imag} */,
  {32'hc0d7951c, 32'hc001ceba} /* (9, 13, 6) {real, imag} */,
  {32'h3f42e3d6, 32'h3f3eb2a1} /* (9, 13, 5) {real, imag} */,
  {32'hc050420c, 32'h412a04a3} /* (9, 13, 4) {real, imag} */,
  {32'h40c8ea3c, 32'hc1081f7c} /* (9, 13, 3) {real, imag} */,
  {32'h4105b41d, 32'hc1060513} /* (9, 13, 2) {real, imag} */,
  {32'hc18ca5bb, 32'h400ff8c4} /* (9, 13, 1) {real, imag} */,
  {32'hc10db11c, 32'hc1468722} /* (9, 13, 0) {real, imag} */,
  {32'hc0e087fe, 32'h418695d8} /* (9, 12, 15) {real, imag} */,
  {32'h403471d4, 32'h40bc0abd} /* (9, 12, 14) {real, imag} */,
  {32'hc0886917, 32'hc1082dd8} /* (9, 12, 13) {real, imag} */,
  {32'h40028734, 32'hc0cc035e} /* (9, 12, 12) {real, imag} */,
  {32'hc095550a, 32'h406459ee} /* (9, 12, 11) {real, imag} */,
  {32'hc049d441, 32'h3d9ef598} /* (9, 12, 10) {real, imag} */,
  {32'hbf82ca90, 32'h3f0392b8} /* (9, 12, 9) {real, imag} */,
  {32'h3f985471, 32'h3fcfacfc} /* (9, 12, 8) {real, imag} */,
  {32'hbcd25800, 32'h3f5bfbd8} /* (9, 12, 7) {real, imag} */,
  {32'h40012497, 32'h3f12d065} /* (9, 12, 6) {real, imag} */,
  {32'h3fc0a3e4, 32'h40875fd5} /* (9, 12, 5) {real, imag} */,
  {32'hbfc937ac, 32'h401ea11b} /* (9, 12, 4) {real, imag} */,
  {32'h40190ae4, 32'hc0512b1e} /* (9, 12, 3) {real, imag} */,
  {32'h40333936, 32'h40bee42b} /* (9, 12, 2) {real, imag} */,
  {32'hc19e42d6, 32'hc0aada71} /* (9, 12, 1) {real, imag} */,
  {32'h408f046d, 32'h3fc0c364} /* (9, 12, 0) {real, imag} */,
  {32'h410c532f, 32'hc00e453e} /* (9, 11, 15) {real, imag} */,
  {32'hbf9a8455, 32'hc0cc6d47} /* (9, 11, 14) {real, imag} */,
  {32'h3fc6779c, 32'h40acbd2a} /* (9, 11, 13) {real, imag} */,
  {32'hbf4a4636, 32'h3ee0d1d0} /* (9, 11, 12) {real, imag} */,
  {32'h403130b7, 32'hc014f33e} /* (9, 11, 11) {real, imag} */,
  {32'hbf40717b, 32'h40019a53} /* (9, 11, 10) {real, imag} */,
  {32'h40498a4b, 32'hbfd3abed} /* (9, 11, 9) {real, imag} */,
  {32'hbf42e878, 32'hbf5557bc} /* (9, 11, 8) {real, imag} */,
  {32'h3f7fe664, 32'hbf492e02} /* (9, 11, 7) {real, imag} */,
  {32'h3f309e01, 32'hbfd94939} /* (9, 11, 6) {real, imag} */,
  {32'h408343c6, 32'h3fe142cc} /* (9, 11, 5) {real, imag} */,
  {32'h40227dc2, 32'hc0f4e71b} /* (9, 11, 4) {real, imag} */,
  {32'hc0eda3f5, 32'h40bc9fbe} /* (9, 11, 3) {real, imag} */,
  {32'hbfd03a8f, 32'h40a14bdb} /* (9, 11, 2) {real, imag} */,
  {32'h3fccf74e, 32'h40a53fba} /* (9, 11, 1) {real, imag} */,
  {32'hc159d26c, 32'h40429d78} /* (9, 11, 0) {real, imag} */,
  {32'h4031ceb0, 32'h40b857a2} /* (9, 10, 15) {real, imag} */,
  {32'h4069a0bb, 32'h404dd04f} /* (9, 10, 14) {real, imag} */,
  {32'hc0b03963, 32'h3ee55d30} /* (9, 10, 13) {real, imag} */,
  {32'hc03a517c, 32'h407e2d64} /* (9, 10, 12) {real, imag} */,
  {32'h3fa4381c, 32'hbdd91a30} /* (9, 10, 11) {real, imag} */,
  {32'hc0543e61, 32'hbf06f668} /* (9, 10, 10) {real, imag} */,
  {32'hbf21f4ec, 32'hbefb77a6} /* (9, 10, 9) {real, imag} */,
  {32'h3e709340, 32'hbfbc86ac} /* (9, 10, 8) {real, imag} */,
  {32'h3eac28d3, 32'h3ddb60e8} /* (9, 10, 7) {real, imag} */,
  {32'h40a613bc, 32'h408892d3} /* (9, 10, 6) {real, imag} */,
  {32'h3fc149bc, 32'h3f7ef2d4} /* (9, 10, 5) {real, imag} */,
  {32'hc0ac848c, 32'h3e1535c8} /* (9, 10, 4) {real, imag} */,
  {32'hc0b9167f, 32'h4085b9b6} /* (9, 10, 3) {real, imag} */,
  {32'h40de516a, 32'hc0a7230e} /* (9, 10, 2) {real, imag} */,
  {32'hbf8df31b, 32'hbfe5bd6e} /* (9, 10, 1) {real, imag} */,
  {32'h3fbd2a5a, 32'h410edd8c} /* (9, 10, 0) {real, imag} */,
  {32'hbfc50982, 32'h4024189a} /* (9, 9, 15) {real, imag} */,
  {32'hc0018a1c, 32'h40d9eb62} /* (9, 9, 14) {real, imag} */,
  {32'h40ad01dc, 32'hbd82a540} /* (9, 9, 13) {real, imag} */,
  {32'h400793d2, 32'hc00a2683} /* (9, 9, 12) {real, imag} */,
  {32'hc05fddd7, 32'hbf83a83c} /* (9, 9, 11) {real, imag} */,
  {32'h402c4f7c, 32'hbfa82c3c} /* (9, 9, 10) {real, imag} */,
  {32'hbf6d3b2c, 32'h3fdf5e58} /* (9, 9, 9) {real, imag} */,
  {32'hbe7295b0, 32'hbee1ed84} /* (9, 9, 8) {real, imag} */,
  {32'hbf81ed52, 32'h3ffe8f72} /* (9, 9, 7) {real, imag} */,
  {32'h3f838d58, 32'h3f5e561f} /* (9, 9, 6) {real, imag} */,
  {32'hbf1d429c, 32'h40607978} /* (9, 9, 5) {real, imag} */,
  {32'h406560a4, 32'hc043c1af} /* (9, 9, 4) {real, imag} */,
  {32'h3f6d862c, 32'h3f8a0869} /* (9, 9, 3) {real, imag} */,
  {32'hc0c9e48c, 32'hc0ae413e} /* (9, 9, 2) {real, imag} */,
  {32'hc0b5a8c2, 32'hbe1c7a78} /* (9, 9, 1) {real, imag} */,
  {32'h40870cec, 32'hc03608a6} /* (9, 9, 0) {real, imag} */,
  {32'hbf372308, 32'hbf307ae1} /* (9, 8, 15) {real, imag} */,
  {32'h404ead68, 32'h3fa2a16b} /* (9, 8, 14) {real, imag} */,
  {32'h40058a9a, 32'hc0511ebc} /* (9, 8, 13) {real, imag} */,
  {32'h3f6f6c86, 32'h40522369} /* (9, 8, 12) {real, imag} */,
  {32'hbfe979d2, 32'hbfdbdbf6} /* (9, 8, 11) {real, imag} */,
  {32'h3d4c30c0, 32'hbe5d5563} /* (9, 8, 10) {real, imag} */,
  {32'h3e0ecaa0, 32'h3f87f4e8} /* (9, 8, 9) {real, imag} */,
  {32'hbd350030, 32'h3f24de0e} /* (9, 8, 8) {real, imag} */,
  {32'hbe98d8c8, 32'hbf365b73} /* (9, 8, 7) {real, imag} */,
  {32'hbfc9fe7b, 32'h3e65101d} /* (9, 8, 6) {real, imag} */,
  {32'h4003ea8d, 32'hbfb33b52} /* (9, 8, 5) {real, imag} */,
  {32'h3fdfe339, 32'h403f3677} /* (9, 8, 4) {real, imag} */,
  {32'hbeed412c, 32'hc024a708} /* (9, 8, 3) {real, imag} */,
  {32'h3fdd7e88, 32'hbfe086a3} /* (9, 8, 2) {real, imag} */,
  {32'h40b0b6e5, 32'h3fa95746} /* (9, 8, 1) {real, imag} */,
  {32'h3fcb7f94, 32'h3fdda871} /* (9, 8, 0) {real, imag} */,
  {32'h40b81fa0, 32'h400be85a} /* (9, 7, 15) {real, imag} */,
  {32'h40d50cf8, 32'hbe66d1c2} /* (9, 7, 14) {real, imag} */,
  {32'h3f103764, 32'h3fad6106} /* (9, 7, 13) {real, imag} */,
  {32'hc09f61f3, 32'h3ea06a37} /* (9, 7, 12) {real, imag} */,
  {32'hbf71c18e, 32'hbf7b997b} /* (9, 7, 11) {real, imag} */,
  {32'hbd75d3c0, 32'hbf35a988} /* (9, 7, 10) {real, imag} */,
  {32'hbe95355a, 32'h3e30a190} /* (9, 7, 9) {real, imag} */,
  {32'h3df23ce0, 32'hbeb5d800} /* (9, 7, 8) {real, imag} */,
  {32'hbf9e4ef0, 32'hbf5c20c0} /* (9, 7, 7) {real, imag} */,
  {32'h3efa12d8, 32'hbe196c32} /* (9, 7, 6) {real, imag} */,
  {32'hbfc3c887, 32'hbe79f1b4} /* (9, 7, 5) {real, imag} */,
  {32'hbfc264b3, 32'hbe9bffb9} /* (9, 7, 4) {real, imag} */,
  {32'h3f7855c8, 32'hc0208871} /* (9, 7, 3) {real, imag} */,
  {32'h4004c9a5, 32'hbf998a1c} /* (9, 7, 2) {real, imag} */,
  {32'h4000670c, 32'h4076e44a} /* (9, 7, 1) {real, imag} */,
  {32'hc057800f, 32'hbfb2fe3e} /* (9, 7, 0) {real, imag} */,
  {32'h40d2df1c, 32'hc010a620} /* (9, 6, 15) {real, imag} */,
  {32'hbfc8ffe1, 32'h408ee5fd} /* (9, 6, 14) {real, imag} */,
  {32'h403e6c41, 32'h3f11ad40} /* (9, 6, 13) {real, imag} */,
  {32'h3f38776b, 32'h3f21a0ee} /* (9, 6, 12) {real, imag} */,
  {32'hc024bcfb, 32'h3fa8c444} /* (9, 6, 11) {real, imag} */,
  {32'hc016c547, 32'hbe6bd940} /* (9, 6, 10) {real, imag} */,
  {32'h3f50b1ac, 32'hbfb4a3db} /* (9, 6, 9) {real, imag} */,
  {32'h3f9d5f35, 32'h3f8f2dac} /* (9, 6, 8) {real, imag} */,
  {32'h3dc3bfe0, 32'hc007efb0} /* (9, 6, 7) {real, imag} */,
  {32'h3fefd9a2, 32'hc00a4020} /* (9, 6, 6) {real, imag} */,
  {32'h3f0a913c, 32'hc0675afa} /* (9, 6, 5) {real, imag} */,
  {32'h3f895720, 32'h408e91b5} /* (9, 6, 4) {real, imag} */,
  {32'hc0065b65, 32'hc0acd0e8} /* (9, 6, 3) {real, imag} */,
  {32'h4026c068, 32'hc08e3187} /* (9, 6, 2) {real, imag} */,
  {32'h3fa8cdfe, 32'hc06c6afa} /* (9, 6, 1) {real, imag} */,
  {32'h402ff814, 32'h40f38797} /* (9, 6, 0) {real, imag} */,
  {32'hc0c8e2b3, 32'h40f457d5} /* (9, 5, 15) {real, imag} */,
  {32'h3fa79967, 32'h3f80c294} /* (9, 5, 14) {real, imag} */,
  {32'hc08d5548, 32'h409c97c3} /* (9, 5, 13) {real, imag} */,
  {32'h3c64f700, 32'h3f2d2ae1} /* (9, 5, 12) {real, imag} */,
  {32'hc04dad9f, 32'hc021f2ca} /* (9, 5, 11) {real, imag} */,
  {32'h3e9d515a, 32'hbcc32680} /* (9, 5, 10) {real, imag} */,
  {32'hc0230f22, 32'hc07a7f9e} /* (9, 5, 9) {real, imag} */,
  {32'hbf544afc, 32'hbf385e5c} /* (9, 5, 8) {real, imag} */,
  {32'h3f9a85d5, 32'hbe58f358} /* (9, 5, 7) {real, imag} */,
  {32'h3fc3b816, 32'h3cb75e80} /* (9, 5, 6) {real, imag} */,
  {32'h3f1c099c, 32'hbd5a9840} /* (9, 5, 5) {real, imag} */,
  {32'h40fd7270, 32'hbfec5564} /* (9, 5, 4) {real, imag} */,
  {32'hbfaf3efa, 32'hbe17cd60} /* (9, 5, 3) {real, imag} */,
  {32'hbf3539fa, 32'hc10838aa} /* (9, 5, 2) {real, imag} */,
  {32'hc14f3200, 32'h417b832e} /* (9, 5, 1) {real, imag} */,
  {32'hbd29e4c0, 32'h406bc1b1} /* (9, 5, 0) {real, imag} */,
  {32'h40ddd4d1, 32'h4118d81d} /* (9, 4, 15) {real, imag} */,
  {32'h4029d198, 32'h40ba1874} /* (9, 4, 14) {real, imag} */,
  {32'hc0a4008a, 32'h3feef8fc} /* (9, 4, 13) {real, imag} */,
  {32'h404d6b21, 32'hc10b058d} /* (9, 4, 12) {real, imag} */,
  {32'h4040fa8c, 32'hc0b27ab4} /* (9, 4, 11) {real, imag} */,
  {32'h405a9d5a, 32'h40a9f498} /* (9, 4, 10) {real, imag} */,
  {32'h3fc89bbc, 32'h3df53f20} /* (9, 4, 9) {real, imag} */,
  {32'h3f8ee156, 32'hbf71dbc3} /* (9, 4, 8) {real, imag} */,
  {32'h3fb93d04, 32'h3f0f1a6c} /* (9, 4, 7) {real, imag} */,
  {32'h3f042f98, 32'hbfbd0d81} /* (9, 4, 6) {real, imag} */,
  {32'hbf797fc0, 32'h3ff92570} /* (9, 4, 5) {real, imag} */,
  {32'hbf1824fc, 32'h403a295d} /* (9, 4, 4) {real, imag} */,
  {32'h4136b8af, 32'hc0d1b0f9} /* (9, 4, 3) {real, imag} */,
  {32'hc0c4e150, 32'hc128a3c2} /* (9, 4, 2) {real, imag} */,
  {32'h417592a0, 32'h417f83f3} /* (9, 4, 1) {real, imag} */,
  {32'hbfb69fda, 32'hc0382831} /* (9, 4, 0) {real, imag} */,
  {32'hc120f401, 32'h3f21d4dc} /* (9, 3, 15) {real, imag} */,
  {32'h3f0faed0, 32'hc04898c0} /* (9, 3, 14) {real, imag} */,
  {32'hc09c7c06, 32'h4000a486} /* (9, 3, 13) {real, imag} */,
  {32'h40be338a, 32'hbe2a7660} /* (9, 3, 12) {real, imag} */,
  {32'h40f0017b, 32'hc0a4dd2a} /* (9, 3, 11) {real, imag} */,
  {32'hbfe00b1e, 32'h3fad14d6} /* (9, 3, 10) {real, imag} */,
  {32'hbf843238, 32'h3febe5ea} /* (9, 3, 9) {real, imag} */,
  {32'h4016569f, 32'hbf2489d0} /* (9, 3, 8) {real, imag} */,
  {32'hbf162b28, 32'h409075de} /* (9, 3, 7) {real, imag} */,
  {32'h3f896c1e, 32'h40221ce9} /* (9, 3, 6) {real, imag} */,
  {32'hc009fa2a, 32'hc039c364} /* (9, 3, 5) {real, imag} */,
  {32'hc033fb57, 32'h410da89e} /* (9, 3, 4) {real, imag} */,
  {32'h40004c6c, 32'h401ebc54} /* (9, 3, 3) {real, imag} */,
  {32'h4018ca06, 32'hc18aec82} /* (9, 3, 2) {real, imag} */,
  {32'h40084a6b, 32'hc02a467d} /* (9, 3, 1) {real, imag} */,
  {32'hc0ed0404, 32'hc10ac8c2} /* (9, 3, 0) {real, imag} */,
  {32'hc110e7cc, 32'hc1359d40} /* (9, 2, 15) {real, imag} */,
  {32'hc0e33294, 32'h41b07a42} /* (9, 2, 14) {real, imag} */,
  {32'hc0c1f2b4, 32'h408b327a} /* (9, 2, 13) {real, imag} */,
  {32'hc13f8da4, 32'hbeeb03d0} /* (9, 2, 12) {real, imag} */,
  {32'h41343960, 32'hc094b04d} /* (9, 2, 11) {real, imag} */,
  {32'h3e3973a8, 32'h3fc07ba4} /* (9, 2, 10) {real, imag} */,
  {32'h40147ca4, 32'hc0a1f7cc} /* (9, 2, 9) {real, imag} */,
  {32'h4073a32e, 32'h3f2b76e0} /* (9, 2, 8) {real, imag} */,
  {32'hbfc19110, 32'hc025b2bc} /* (9, 2, 7) {real, imag} */,
  {32'hbf96ebfb, 32'h3eb9d870} /* (9, 2, 6) {real, imag} */,
  {32'hbff31884, 32'h409fe5a3} /* (9, 2, 5) {real, imag} */,
  {32'h406dca28, 32'h4158cff2} /* (9, 2, 4) {real, imag} */,
  {32'hbd3480c0, 32'hc13a5ffb} /* (9, 2, 3) {real, imag} */,
  {32'h413cfa58, 32'hc07d3c50} /* (9, 2, 2) {real, imag} */,
  {32'hc0d1937e, 32'hc1754d8c} /* (9, 2, 1) {real, imag} */,
  {32'h410d1bba, 32'h40c641e3} /* (9, 2, 0) {real, imag} */,
  {32'hc171de82, 32'h418b1588} /* (9, 1, 15) {real, imag} */,
  {32'hc01514c4, 32'hc1aae62a} /* (9, 1, 14) {real, imag} */,
  {32'hc104c2c8, 32'hbf876bf4} /* (9, 1, 13) {real, imag} */,
  {32'h40ec9b50, 32'hc0be4cec} /* (9, 1, 12) {real, imag} */,
  {32'hbf8061d0, 32'h405d51fc} /* (9, 1, 11) {real, imag} */,
  {32'hbd83c360, 32'hc02e00f4} /* (9, 1, 10) {real, imag} */,
  {32'hbf1e8b48, 32'h4115af96} /* (9, 1, 9) {real, imag} */,
  {32'h3e825ac8, 32'h400e1232} /* (9, 1, 8) {real, imag} */,
  {32'hbf0fc5c8, 32'hbf018588} /* (9, 1, 7) {real, imag} */,
  {32'hc09d3792, 32'h41045857} /* (9, 1, 6) {real, imag} */,
  {32'h402e6588, 32'hc14abe35} /* (9, 1, 5) {real, imag} */,
  {32'hbf8d9a36, 32'hc09680a0} /* (9, 1, 4) {real, imag} */,
  {32'h41abd5d4, 32'h3f2b4088} /* (9, 1, 3) {real, imag} */,
  {32'hc1587a73, 32'h40cf0542} /* (9, 1, 2) {real, imag} */,
  {32'h419d35ff, 32'h41337aba} /* (9, 1, 1) {real, imag} */,
  {32'h400e1f51, 32'h40da91f3} /* (9, 1, 0) {real, imag} */,
  {32'h41867d91, 32'hc124878c} /* (9, 0, 15) {real, imag} */,
  {32'hc12b0db2, 32'hc13bffb4} /* (9, 0, 14) {real, imag} */,
  {32'h418ffd1b, 32'hbd930980} /* (9, 0, 13) {real, imag} */,
  {32'hc08a5298, 32'h3f45f76c} /* (9, 0, 12) {real, imag} */,
  {32'hc11a3128, 32'h3fd3b280} /* (9, 0, 11) {real, imag} */,
  {32'h40068261, 32'h4136496e} /* (9, 0, 10) {real, imag} */,
  {32'h40ac2455, 32'hbf907742} /* (9, 0, 9) {real, imag} */,
  {32'hc0d3aaaa, 32'h4090d97e} /* (9, 0, 8) {real, imag} */,
  {32'h401265d2, 32'hbf4bcbec} /* (9, 0, 7) {real, imag} */,
  {32'hbe3085b0, 32'h3feb3a3c} /* (9, 0, 6) {real, imag} */,
  {32'h3ee47f70, 32'hc11b3a54} /* (9, 0, 5) {real, imag} */,
  {32'hbef8f128, 32'hc091abf8} /* (9, 0, 4) {real, imag} */,
  {32'hc087eb9c, 32'h4185f596} /* (9, 0, 3) {real, imag} */,
  {32'h40d970f4, 32'h3f4a83c8} /* (9, 0, 2) {real, imag} */,
  {32'hc1330a6a, 32'hc16b42d4} /* (9, 0, 1) {real, imag} */,
  {32'h40901c58, 32'hc19b0e22} /* (9, 0, 0) {real, imag} */,
  {32'h400b9751, 32'hbed3d900} /* (8, 15, 15) {real, imag} */,
  {32'hc1660e40, 32'hc010cb68} /* (8, 15, 14) {real, imag} */,
  {32'h40870469, 32'h3ddd60c0} /* (8, 15, 13) {real, imag} */,
  {32'hc119ac72, 32'h3e115558} /* (8, 15, 12) {real, imag} */,
  {32'h400099a8, 32'hc08a9642} /* (8, 15, 11) {real, imag} */,
  {32'hc0c7a232, 32'hc00df7ac} /* (8, 15, 10) {real, imag} */,
  {32'h402abb2c, 32'h404fa06b} /* (8, 15, 9) {real, imag} */,
  {32'hbf3b979a, 32'h4002b61a} /* (8, 15, 8) {real, imag} */,
  {32'hc027e440, 32'hbefedc38} /* (8, 15, 7) {real, imag} */,
  {32'hc04ad530, 32'hbe95aea0} /* (8, 15, 6) {real, imag} */,
  {32'h409a09f4, 32'h401ed731} /* (8, 15, 5) {real, imag} */,
  {32'h40248dc2, 32'hbfb2025d} /* (8, 15, 4) {real, imag} */,
  {32'hc05719f6, 32'h41207d8a} /* (8, 15, 3) {real, imag} */,
  {32'h3f8d8968, 32'hc14c51c6} /* (8, 15, 2) {real, imag} */,
  {32'hc0f6cd26, 32'hc189945c} /* (8, 15, 1) {real, imag} */,
  {32'hc03beeec, 32'h404af126} /* (8, 15, 0) {real, imag} */,
  {32'hc09087c0, 32'hc1cdbc95} /* (8, 14, 15) {real, imag} */,
  {32'hc000ede8, 32'h4177c09b} /* (8, 14, 14) {real, imag} */,
  {32'hc0c88949, 32'hc07ad9ae} /* (8, 14, 13) {real, imag} */,
  {32'hc0069596, 32'hc10e92b0} /* (8, 14, 12) {real, imag} */,
  {32'h3fb2e559, 32'h41015046} /* (8, 14, 11) {real, imag} */,
  {32'h3f79cc10, 32'hc0210c46} /* (8, 14, 10) {real, imag} */,
  {32'h3e145cd0, 32'hbf30c760} /* (8, 14, 9) {real, imag} */,
  {32'hbf3bff22, 32'h4080148f} /* (8, 14, 8) {real, imag} */,
  {32'h40998bd2, 32'h4089a554} /* (8, 14, 7) {real, imag} */,
  {32'h4070ed98, 32'hbea48410} /* (8, 14, 6) {real, imag} */,
  {32'hbf5e587a, 32'h4119f85a} /* (8, 14, 5) {real, imag} */,
  {32'h410db0ba, 32'h40dd331c} /* (8, 14, 4) {real, imag} */,
  {32'hc0aae66f, 32'hc06392f4} /* (8, 14, 3) {real, imag} */,
  {32'hbf0bc428, 32'h4084c08e} /* (8, 14, 2) {real, imag} */,
  {32'h3cc0bd80, 32'hbf29fea0} /* (8, 14, 1) {real, imag} */,
  {32'hc02c0112, 32'h412e5bc0} /* (8, 14, 0) {real, imag} */,
  {32'hc1415404, 32'h404a0e14} /* (8, 13, 15) {real, imag} */,
  {32'hc0085aa4, 32'hbf9cc402} /* (8, 13, 14) {real, imag} */,
  {32'h404c9d50, 32'hc0b76f14} /* (8, 13, 13) {real, imag} */,
  {32'h403d395a, 32'h408f2493} /* (8, 13, 12) {real, imag} */,
  {32'hc0d24546, 32'h3f733e28} /* (8, 13, 11) {real, imag} */,
  {32'h3f5df5f8, 32'h4088fa6c} /* (8, 13, 10) {real, imag} */,
  {32'h405b2f74, 32'h4078cdaa} /* (8, 13, 9) {real, imag} */,
  {32'hbfdf51a8, 32'hbffa6ce7} /* (8, 13, 8) {real, imag} */,
  {32'h3f320830, 32'h4030d6a2} /* (8, 13, 7) {real, imag} */,
  {32'h4047f2c8, 32'hc08bd7ae} /* (8, 13, 6) {real, imag} */,
  {32'hc0042915, 32'h40a2f35f} /* (8, 13, 5) {real, imag} */,
  {32'h40473f14, 32'hc0a35ee3} /* (8, 13, 4) {real, imag} */,
  {32'hc1402a52, 32'h40578000} /* (8, 13, 3) {real, imag} */,
  {32'hbec8811e, 32'h4086728c} /* (8, 13, 2) {real, imag} */,
  {32'h404ca08a, 32'hc12b6b4f} /* (8, 13, 1) {real, imag} */,
  {32'hc0d1c342, 32'h3fe4e9ab} /* (8, 13, 0) {real, imag} */,
  {32'hc106e32c, 32'hc0c37b8c} /* (8, 12, 15) {real, imag} */,
  {32'h3f7ca410, 32'hc0974170} /* (8, 12, 14) {real, imag} */,
  {32'hbfaf12d1, 32'h40fd5288} /* (8, 12, 13) {real, imag} */,
  {32'h3f95b2dc, 32'h409ce8bc} /* (8, 12, 12) {real, imag} */,
  {32'h3fc5f9e3, 32'h3e522630} /* (8, 12, 11) {real, imag} */,
  {32'hbf0eac84, 32'hbfcf6374} /* (8, 12, 10) {real, imag} */,
  {32'h3d937ea0, 32'h3fc449f8} /* (8, 12, 9) {real, imag} */,
  {32'hc03893de, 32'hbfaf6e80} /* (8, 12, 8) {real, imag} */,
  {32'h404a8b35, 32'hc04866b2} /* (8, 12, 7) {real, imag} */,
  {32'h3f47d6c4, 32'hbf4c317c} /* (8, 12, 6) {real, imag} */,
  {32'h3fe1c5a5, 32'h3f7c6834} /* (8, 12, 5) {real, imag} */,
  {32'hbe8b1e82, 32'hc0c32610} /* (8, 12, 4) {real, imag} */,
  {32'h3ef61c84, 32'h40810b02} /* (8, 12, 3) {real, imag} */,
  {32'h413a618d, 32'hbff982e2} /* (8, 12, 2) {real, imag} */,
  {32'hc1147d98, 32'h415029c6} /* (8, 12, 1) {real, imag} */,
  {32'h40859d59, 32'hc13973c0} /* (8, 12, 0) {real, imag} */,
  {32'h40ac489a, 32'h40e84504} /* (8, 11, 15) {real, imag} */,
  {32'hc0e0dd97, 32'h40bdafe6} /* (8, 11, 14) {real, imag} */,
  {32'h410c17d3, 32'hc0a42c60} /* (8, 11, 13) {real, imag} */,
  {32'h404eea73, 32'h40162231} /* (8, 11, 12) {real, imag} */,
  {32'hbf85382a, 32'hbf882c4a} /* (8, 11, 11) {real, imag} */,
  {32'h3e6ddeb8, 32'h3e718930} /* (8, 11, 10) {real, imag} */,
  {32'hbe138e34, 32'h3ecae708} /* (8, 11, 9) {real, imag} */,
  {32'h3fc9b686, 32'hbf9af45e} /* (8, 11, 8) {real, imag} */,
  {32'hbf393b15, 32'h3ff92d3a} /* (8, 11, 7) {real, imag} */,
  {32'h3fb0f819, 32'h3fa4856e} /* (8, 11, 6) {real, imag} */,
  {32'h403b6133, 32'h400638c9} /* (8, 11, 5) {real, imag} */,
  {32'h40374ec1, 32'h3fd47c76} /* (8, 11, 4) {real, imag} */,
  {32'h40a341a6, 32'hbfed3b72} /* (8, 11, 3) {real, imag} */,
  {32'hc08a8131, 32'h40e04212} /* (8, 11, 2) {real, imag} */,
  {32'hc0a1b412, 32'h3fceb9f0} /* (8, 11, 1) {real, imag} */,
  {32'h40bef338, 32'hc08e3e50} /* (8, 11, 0) {real, imag} */,
  {32'hc0528d88, 32'hbfb7cb04} /* (8, 10, 15) {real, imag} */,
  {32'hc0af3cb5, 32'hc09dcd9e} /* (8, 10, 14) {real, imag} */,
  {32'hc02bb6a3, 32'hc0029d5e} /* (8, 10, 13) {real, imag} */,
  {32'h3f7d3f4c, 32'hbff4c676} /* (8, 10, 12) {real, imag} */,
  {32'h401c41ac, 32'h3f0c9892} /* (8, 10, 11) {real, imag} */,
  {32'hbff343fc, 32'hbf8f88dc} /* (8, 10, 10) {real, imag} */,
  {32'h3e8e8ac6, 32'h3fab27b0} /* (8, 10, 9) {real, imag} */,
  {32'h3f0cfca2, 32'h3efc0f4c} /* (8, 10, 8) {real, imag} */,
  {32'hbfa529d2, 32'h3dacd9a0} /* (8, 10, 7) {real, imag} */,
  {32'hbf002c8b, 32'h3fa663c4} /* (8, 10, 6) {real, imag} */,
  {32'hc01b3c36, 32'hbf641256} /* (8, 10, 5) {real, imag} */,
  {32'h3fbf35a4, 32'h4032fd03} /* (8, 10, 4) {real, imag} */,
  {32'h3e9f62b8, 32'hc04c8c5e} /* (8, 10, 3) {real, imag} */,
  {32'hbfcda74c, 32'h3e987b10} /* (8, 10, 2) {real, imag} */,
  {32'h40c9c034, 32'hbf8903a4} /* (8, 10, 1) {real, imag} */,
  {32'hbfff84bb, 32'h402787c0} /* (8, 10, 0) {real, imag} */,
  {32'hc075311d, 32'hbeebdc9e} /* (8, 9, 15) {real, imag} */,
  {32'h408ab798, 32'h4060153f} /* (8, 9, 14) {real, imag} */,
  {32'hbfdb0b03, 32'h407ee852} /* (8, 9, 13) {real, imag} */,
  {32'hbf96a707, 32'hc027055a} /* (8, 9, 12) {real, imag} */,
  {32'h3f9afb41, 32'h4000a796} /* (8, 9, 11) {real, imag} */,
  {32'hbf0fae32, 32'h3f89298f} /* (8, 9, 10) {real, imag} */,
  {32'h3f6abf4e, 32'hbe500834} /* (8, 9, 9) {real, imag} */,
  {32'hbf1cd788, 32'h3e81aa08} /* (8, 9, 8) {real, imag} */,
  {32'h3d774198, 32'hbfcda394} /* (8, 9, 7) {real, imag} */,
  {32'h3f9808d7, 32'h3f757072} /* (8, 9, 6) {real, imag} */,
  {32'h3fca3e8f, 32'hbeaf8b44} /* (8, 9, 5) {real, imag} */,
  {32'h3e340f28, 32'h3e54a100} /* (8, 9, 4) {real, imag} */,
  {32'hbe53c8a8, 32'hbebcd63c} /* (8, 9, 3) {real, imag} */,
  {32'hbfb2f261, 32'hc042caf1} /* (8, 9, 2) {real, imag} */,
  {32'h3fc91936, 32'h3fdb8ea0} /* (8, 9, 1) {real, imag} */,
  {32'h400bc6d8, 32'hc0860b02} /* (8, 9, 0) {real, imag} */,
  {32'h40cbd5c2, 32'h3f5e644c} /* (8, 8, 15) {real, imag} */,
  {32'hbe3769e6, 32'hbda38816} /* (8, 8, 14) {real, imag} */,
  {32'hbec784d2, 32'h3fe7a3a7} /* (8, 8, 13) {real, imag} */,
  {32'hbf82ef99, 32'hbfb25980} /* (8, 8, 12) {real, imag} */,
  {32'hbfcc1ae0, 32'hbe082b18} /* (8, 8, 11) {real, imag} */,
  {32'h3f8774d3, 32'h3e91da2a} /* (8, 8, 10) {real, imag} */,
  {32'hbfded7e6, 32'h3f154396} /* (8, 8, 9) {real, imag} */,
  {32'h3f31048c, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'hbfded7e6, 32'hbf154396} /* (8, 8, 7) {real, imag} */,
  {32'h3f8774d3, 32'hbe91da2a} /* (8, 8, 6) {real, imag} */,
  {32'hbfcc1ae0, 32'h3e082b18} /* (8, 8, 5) {real, imag} */,
  {32'hbf82ef99, 32'h3fb25980} /* (8, 8, 4) {real, imag} */,
  {32'hbec784d2, 32'hbfe7a3a7} /* (8, 8, 3) {real, imag} */,
  {32'hbe3769e6, 32'h3da38816} /* (8, 8, 2) {real, imag} */,
  {32'h40cbd5c2, 32'hbf5e644c} /* (8, 8, 1) {real, imag} */,
  {32'hbeedcc21, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h3fc91936, 32'hbfdb8ea0} /* (8, 7, 15) {real, imag} */,
  {32'hbfb2f261, 32'h4042caf1} /* (8, 7, 14) {real, imag} */,
  {32'hbe53c8a8, 32'h3ebcd63c} /* (8, 7, 13) {real, imag} */,
  {32'h3e340f28, 32'hbe54a100} /* (8, 7, 12) {real, imag} */,
  {32'h3fca3e8f, 32'h3eaf8b44} /* (8, 7, 11) {real, imag} */,
  {32'h3f9808d7, 32'hbf757072} /* (8, 7, 10) {real, imag} */,
  {32'h3d774198, 32'h3fcda394} /* (8, 7, 9) {real, imag} */,
  {32'hbf1cd788, 32'hbe81aa08} /* (8, 7, 8) {real, imag} */,
  {32'h3f6abf4e, 32'h3e500834} /* (8, 7, 7) {real, imag} */,
  {32'hbf0fae32, 32'hbf89298f} /* (8, 7, 6) {real, imag} */,
  {32'h3f9afb41, 32'hc000a796} /* (8, 7, 5) {real, imag} */,
  {32'hbf96a707, 32'h4027055a} /* (8, 7, 4) {real, imag} */,
  {32'hbfdb0b03, 32'hc07ee852} /* (8, 7, 3) {real, imag} */,
  {32'h408ab798, 32'hc060153f} /* (8, 7, 2) {real, imag} */,
  {32'hc075311d, 32'h3eebdc9e} /* (8, 7, 1) {real, imag} */,
  {32'h400bc6d8, 32'h40860b02} /* (8, 7, 0) {real, imag} */,
  {32'h40c9c034, 32'h3f8903a4} /* (8, 6, 15) {real, imag} */,
  {32'hbfcda74c, 32'hbe987b10} /* (8, 6, 14) {real, imag} */,
  {32'h3e9f62b8, 32'h404c8c5e} /* (8, 6, 13) {real, imag} */,
  {32'h3fbf35a4, 32'hc032fd03} /* (8, 6, 12) {real, imag} */,
  {32'hc01b3c36, 32'h3f641256} /* (8, 6, 11) {real, imag} */,
  {32'hbf002c8b, 32'hbfa663c4} /* (8, 6, 10) {real, imag} */,
  {32'hbfa529d2, 32'hbdacd9a0} /* (8, 6, 9) {real, imag} */,
  {32'h3f0cfca2, 32'hbefc0f4c} /* (8, 6, 8) {real, imag} */,
  {32'h3e8e8ac6, 32'hbfab27b0} /* (8, 6, 7) {real, imag} */,
  {32'hbff343fc, 32'h3f8f88dc} /* (8, 6, 6) {real, imag} */,
  {32'h401c41ac, 32'hbf0c9892} /* (8, 6, 5) {real, imag} */,
  {32'h3f7d3f4c, 32'h3ff4c676} /* (8, 6, 4) {real, imag} */,
  {32'hc02bb6a3, 32'h40029d5e} /* (8, 6, 3) {real, imag} */,
  {32'hc0af3cb5, 32'h409dcd9e} /* (8, 6, 2) {real, imag} */,
  {32'hc0528d88, 32'h3fb7cb04} /* (8, 6, 1) {real, imag} */,
  {32'hbfff84bb, 32'hc02787c0} /* (8, 6, 0) {real, imag} */,
  {32'hc0a1b412, 32'hbfceb9f0} /* (8, 5, 15) {real, imag} */,
  {32'hc08a8131, 32'hc0e04212} /* (8, 5, 14) {real, imag} */,
  {32'h40a341a6, 32'h3fed3b72} /* (8, 5, 13) {real, imag} */,
  {32'h40374ec1, 32'hbfd47c76} /* (8, 5, 12) {real, imag} */,
  {32'h403b6133, 32'hc00638c9} /* (8, 5, 11) {real, imag} */,
  {32'h3fb0f819, 32'hbfa4856e} /* (8, 5, 10) {real, imag} */,
  {32'hbf393b15, 32'hbff92d3a} /* (8, 5, 9) {real, imag} */,
  {32'h3fc9b686, 32'h3f9af45e} /* (8, 5, 8) {real, imag} */,
  {32'hbe138e34, 32'hbecae708} /* (8, 5, 7) {real, imag} */,
  {32'h3e6ddeb8, 32'hbe718930} /* (8, 5, 6) {real, imag} */,
  {32'hbf85382a, 32'h3f882c4a} /* (8, 5, 5) {real, imag} */,
  {32'h404eea73, 32'hc0162231} /* (8, 5, 4) {real, imag} */,
  {32'h410c17d3, 32'h40a42c60} /* (8, 5, 3) {real, imag} */,
  {32'hc0e0dd97, 32'hc0bdafe6} /* (8, 5, 2) {real, imag} */,
  {32'h40ac489a, 32'hc0e84504} /* (8, 5, 1) {real, imag} */,
  {32'h40bef338, 32'h408e3e50} /* (8, 5, 0) {real, imag} */,
  {32'hc1147d98, 32'hc15029c6} /* (8, 4, 15) {real, imag} */,
  {32'h413a618d, 32'h3ff982e2} /* (8, 4, 14) {real, imag} */,
  {32'h3ef61c84, 32'hc0810b02} /* (8, 4, 13) {real, imag} */,
  {32'hbe8b1e82, 32'h40c32610} /* (8, 4, 12) {real, imag} */,
  {32'h3fe1c5a5, 32'hbf7c6834} /* (8, 4, 11) {real, imag} */,
  {32'h3f47d6c4, 32'h3f4c317c} /* (8, 4, 10) {real, imag} */,
  {32'h404a8b35, 32'h404866b2} /* (8, 4, 9) {real, imag} */,
  {32'hc03893de, 32'h3faf6e80} /* (8, 4, 8) {real, imag} */,
  {32'h3d937ea0, 32'hbfc449f8} /* (8, 4, 7) {real, imag} */,
  {32'hbf0eac84, 32'h3fcf6374} /* (8, 4, 6) {real, imag} */,
  {32'h3fc5f9e3, 32'hbe522630} /* (8, 4, 5) {real, imag} */,
  {32'h3f95b2dc, 32'hc09ce8bc} /* (8, 4, 4) {real, imag} */,
  {32'hbfaf12d1, 32'hc0fd5288} /* (8, 4, 3) {real, imag} */,
  {32'h3f7ca410, 32'h40974170} /* (8, 4, 2) {real, imag} */,
  {32'hc106e32c, 32'h40c37b8c} /* (8, 4, 1) {real, imag} */,
  {32'h40859d59, 32'h413973c0} /* (8, 4, 0) {real, imag} */,
  {32'h404ca08a, 32'h412b6b4f} /* (8, 3, 15) {real, imag} */,
  {32'hbec8811e, 32'hc086728c} /* (8, 3, 14) {real, imag} */,
  {32'hc1402a52, 32'hc0578000} /* (8, 3, 13) {real, imag} */,
  {32'h40473f14, 32'h40a35ee3} /* (8, 3, 12) {real, imag} */,
  {32'hc0042915, 32'hc0a2f35f} /* (8, 3, 11) {real, imag} */,
  {32'h4047f2c8, 32'h408bd7ae} /* (8, 3, 10) {real, imag} */,
  {32'h3f320830, 32'hc030d6a2} /* (8, 3, 9) {real, imag} */,
  {32'hbfdf51a8, 32'h3ffa6ce7} /* (8, 3, 8) {real, imag} */,
  {32'h405b2f74, 32'hc078cdaa} /* (8, 3, 7) {real, imag} */,
  {32'h3f5df5f8, 32'hc088fa6c} /* (8, 3, 6) {real, imag} */,
  {32'hc0d24546, 32'hbf733e28} /* (8, 3, 5) {real, imag} */,
  {32'h403d395a, 32'hc08f2493} /* (8, 3, 4) {real, imag} */,
  {32'h404c9d50, 32'h40b76f14} /* (8, 3, 3) {real, imag} */,
  {32'hc0085aa4, 32'h3f9cc402} /* (8, 3, 2) {real, imag} */,
  {32'hc1415404, 32'hc04a0e14} /* (8, 3, 1) {real, imag} */,
  {32'hc0d1c342, 32'hbfe4e9ab} /* (8, 3, 0) {real, imag} */,
  {32'h3cc0bd80, 32'h3f29fea0} /* (8, 2, 15) {real, imag} */,
  {32'hbf0bc428, 32'hc084c08e} /* (8, 2, 14) {real, imag} */,
  {32'hc0aae66f, 32'h406392f4} /* (8, 2, 13) {real, imag} */,
  {32'h410db0ba, 32'hc0dd331c} /* (8, 2, 12) {real, imag} */,
  {32'hbf5e587a, 32'hc119f85a} /* (8, 2, 11) {real, imag} */,
  {32'h4070ed98, 32'h3ea48410} /* (8, 2, 10) {real, imag} */,
  {32'h40998bd2, 32'hc089a554} /* (8, 2, 9) {real, imag} */,
  {32'hbf3bff22, 32'hc080148f} /* (8, 2, 8) {real, imag} */,
  {32'h3e145cd0, 32'h3f30c760} /* (8, 2, 7) {real, imag} */,
  {32'h3f79cc10, 32'h40210c46} /* (8, 2, 6) {real, imag} */,
  {32'h3fb2e559, 32'hc1015046} /* (8, 2, 5) {real, imag} */,
  {32'hc0069596, 32'h410e92b0} /* (8, 2, 4) {real, imag} */,
  {32'hc0c88949, 32'h407ad9ae} /* (8, 2, 3) {real, imag} */,
  {32'hc000ede8, 32'hc177c09b} /* (8, 2, 2) {real, imag} */,
  {32'hc09087c0, 32'h41cdbc95} /* (8, 2, 1) {real, imag} */,
  {32'hc02c0112, 32'hc12e5bc0} /* (8, 2, 0) {real, imag} */,
  {32'hc0f6cd26, 32'h4189945c} /* (8, 1, 15) {real, imag} */,
  {32'h3f8d8968, 32'h414c51c6} /* (8, 1, 14) {real, imag} */,
  {32'hc05719f6, 32'hc1207d8a} /* (8, 1, 13) {real, imag} */,
  {32'h40248dc2, 32'h3fb2025d} /* (8, 1, 12) {real, imag} */,
  {32'h409a09f4, 32'hc01ed731} /* (8, 1, 11) {real, imag} */,
  {32'hc04ad530, 32'h3e95aea0} /* (8, 1, 10) {real, imag} */,
  {32'hc027e440, 32'h3efedc38} /* (8, 1, 9) {real, imag} */,
  {32'hbf3b979a, 32'hc002b61a} /* (8, 1, 8) {real, imag} */,
  {32'h402abb2c, 32'hc04fa06b} /* (8, 1, 7) {real, imag} */,
  {32'hc0c7a232, 32'h400df7ac} /* (8, 1, 6) {real, imag} */,
  {32'h400099a8, 32'h408a9642} /* (8, 1, 5) {real, imag} */,
  {32'hc119ac72, 32'hbe115558} /* (8, 1, 4) {real, imag} */,
  {32'h40870469, 32'hbddd60c0} /* (8, 1, 3) {real, imag} */,
  {32'hc1660e40, 32'h4010cb68} /* (8, 1, 2) {real, imag} */,
  {32'h400b9751, 32'h3ed3d900} /* (8, 1, 1) {real, imag} */,
  {32'hc03beeec, 32'hc04af126} /* (8, 1, 0) {real, imag} */,
  {32'h40a7f624, 32'hc084ab10} /* (8, 0, 15) {real, imag} */,
  {32'h40368b04, 32'hbfafedc8} /* (8, 0, 14) {real, imag} */,
  {32'h4071f099, 32'hc01030df} /* (8, 0, 13) {real, imag} */,
  {32'hc0812a3c, 32'hc0343c93} /* (8, 0, 12) {real, imag} */,
  {32'hbf2b8eec, 32'hbfcee4fe} /* (8, 0, 11) {real, imag} */,
  {32'h3fbe73a1, 32'h3fcc081a} /* (8, 0, 10) {real, imag} */,
  {32'hc04aa809, 32'hc013b5bc} /* (8, 0, 9) {real, imag} */,
  {32'h406a41d5, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'hc04aa809, 32'h4013b5bc} /* (8, 0, 7) {real, imag} */,
  {32'h3fbe73a1, 32'hbfcc081a} /* (8, 0, 6) {real, imag} */,
  {32'hbf2b8eec, 32'h3fcee4fe} /* (8, 0, 5) {real, imag} */,
  {32'hc0812a3c, 32'h40343c93} /* (8, 0, 4) {real, imag} */,
  {32'h4071f099, 32'h401030df} /* (8, 0, 3) {real, imag} */,
  {32'h40368b04, 32'h3fafedc8} /* (8, 0, 2) {real, imag} */,
  {32'h40a7f624, 32'h4084ab10} /* (8, 0, 1) {real, imag} */,
  {32'h408475a6, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h419d35ff, 32'hc1337aba} /* (7, 15, 15) {real, imag} */,
  {32'hc1587a73, 32'hc0cf0542} /* (7, 15, 14) {real, imag} */,
  {32'h41abd5d4, 32'hbf2b4088} /* (7, 15, 13) {real, imag} */,
  {32'hbf8d9a36, 32'h409680a0} /* (7, 15, 12) {real, imag} */,
  {32'h402e6588, 32'h414abe35} /* (7, 15, 11) {real, imag} */,
  {32'hc09d3792, 32'hc1045857} /* (7, 15, 10) {real, imag} */,
  {32'hbf0fc5c8, 32'h3f018588} /* (7, 15, 9) {real, imag} */,
  {32'h3e825ac8, 32'hc00e1232} /* (7, 15, 8) {real, imag} */,
  {32'hbf1e8b48, 32'hc115af96} /* (7, 15, 7) {real, imag} */,
  {32'hbd83c360, 32'h402e00f4} /* (7, 15, 6) {real, imag} */,
  {32'hbf8061d0, 32'hc05d51fc} /* (7, 15, 5) {real, imag} */,
  {32'h40ec9b50, 32'h40be4cec} /* (7, 15, 4) {real, imag} */,
  {32'hc104c2c8, 32'h3f876bf4} /* (7, 15, 3) {real, imag} */,
  {32'hc01514c4, 32'h41aae62a} /* (7, 15, 2) {real, imag} */,
  {32'hc171de82, 32'hc18b1588} /* (7, 15, 1) {real, imag} */,
  {32'h400e1f51, 32'hc0da91f3} /* (7, 15, 0) {real, imag} */,
  {32'hc0d1937e, 32'h41754d8c} /* (7, 14, 15) {real, imag} */,
  {32'h413cfa58, 32'h407d3c50} /* (7, 14, 14) {real, imag} */,
  {32'hbd3480c0, 32'h413a5ffb} /* (7, 14, 13) {real, imag} */,
  {32'h406dca28, 32'hc158cff2} /* (7, 14, 12) {real, imag} */,
  {32'hbff31884, 32'hc09fe5a3} /* (7, 14, 11) {real, imag} */,
  {32'hbf96ebfb, 32'hbeb9d870} /* (7, 14, 10) {real, imag} */,
  {32'hbfc19110, 32'h4025b2bc} /* (7, 14, 9) {real, imag} */,
  {32'h4073a32e, 32'hbf2b76e0} /* (7, 14, 8) {real, imag} */,
  {32'h40147ca4, 32'h40a1f7cc} /* (7, 14, 7) {real, imag} */,
  {32'h3e3973a8, 32'hbfc07ba4} /* (7, 14, 6) {real, imag} */,
  {32'h41343960, 32'h4094b04d} /* (7, 14, 5) {real, imag} */,
  {32'hc13f8da4, 32'h3eeb03d0} /* (7, 14, 4) {real, imag} */,
  {32'hc0c1f2b4, 32'hc08b327a} /* (7, 14, 3) {real, imag} */,
  {32'hc0e33294, 32'hc1b07a42} /* (7, 14, 2) {real, imag} */,
  {32'hc110e7cc, 32'h41359d40} /* (7, 14, 1) {real, imag} */,
  {32'h410d1bba, 32'hc0c641e3} /* (7, 14, 0) {real, imag} */,
  {32'h40084a6b, 32'h402a467d} /* (7, 13, 15) {real, imag} */,
  {32'h4018ca06, 32'h418aec82} /* (7, 13, 14) {real, imag} */,
  {32'h40004c6c, 32'hc01ebc54} /* (7, 13, 13) {real, imag} */,
  {32'hc033fb57, 32'hc10da89e} /* (7, 13, 12) {real, imag} */,
  {32'hc009fa2a, 32'h4039c364} /* (7, 13, 11) {real, imag} */,
  {32'h3f896c1e, 32'hc0221ce9} /* (7, 13, 10) {real, imag} */,
  {32'hbf162b28, 32'hc09075de} /* (7, 13, 9) {real, imag} */,
  {32'h4016569f, 32'h3f2489d0} /* (7, 13, 8) {real, imag} */,
  {32'hbf843238, 32'hbfebe5ea} /* (7, 13, 7) {real, imag} */,
  {32'hbfe00b1e, 32'hbfad14d6} /* (7, 13, 6) {real, imag} */,
  {32'h40f0017b, 32'h40a4dd2a} /* (7, 13, 5) {real, imag} */,
  {32'h40be338a, 32'h3e2a7660} /* (7, 13, 4) {real, imag} */,
  {32'hc09c7c06, 32'hc000a486} /* (7, 13, 3) {real, imag} */,
  {32'h3f0faed0, 32'h404898c0} /* (7, 13, 2) {real, imag} */,
  {32'hc120f401, 32'hbf21d4dc} /* (7, 13, 1) {real, imag} */,
  {32'hc0ed0404, 32'h410ac8c2} /* (7, 13, 0) {real, imag} */,
  {32'h417592a0, 32'hc17f83f3} /* (7, 12, 15) {real, imag} */,
  {32'hc0c4e150, 32'h4128a3c2} /* (7, 12, 14) {real, imag} */,
  {32'h4136b8af, 32'h40d1b0f9} /* (7, 12, 13) {real, imag} */,
  {32'hbf1824fc, 32'hc03a295d} /* (7, 12, 12) {real, imag} */,
  {32'hbf797fc0, 32'hbff92570} /* (7, 12, 11) {real, imag} */,
  {32'h3f042f98, 32'h3fbd0d81} /* (7, 12, 10) {real, imag} */,
  {32'h3fb93d04, 32'hbf0f1a6c} /* (7, 12, 9) {real, imag} */,
  {32'h3f8ee156, 32'h3f71dbc3} /* (7, 12, 8) {real, imag} */,
  {32'h3fc89bbc, 32'hbdf53f20} /* (7, 12, 7) {real, imag} */,
  {32'h405a9d5a, 32'hc0a9f498} /* (7, 12, 6) {real, imag} */,
  {32'h4040fa8c, 32'h40b27ab4} /* (7, 12, 5) {real, imag} */,
  {32'h404d6b21, 32'h410b058d} /* (7, 12, 4) {real, imag} */,
  {32'hc0a4008a, 32'hbfeef8fc} /* (7, 12, 3) {real, imag} */,
  {32'h4029d198, 32'hc0ba1874} /* (7, 12, 2) {real, imag} */,
  {32'h40ddd4d1, 32'hc118d81d} /* (7, 12, 1) {real, imag} */,
  {32'hbfb69fda, 32'h40382831} /* (7, 12, 0) {real, imag} */,
  {32'hc14f3200, 32'hc17b832e} /* (7, 11, 15) {real, imag} */,
  {32'hbf3539fa, 32'h410838aa} /* (7, 11, 14) {real, imag} */,
  {32'hbfaf3efa, 32'h3e17cd60} /* (7, 11, 13) {real, imag} */,
  {32'h40fd7270, 32'h3fec5564} /* (7, 11, 12) {real, imag} */,
  {32'h3f1c099c, 32'h3d5a9840} /* (7, 11, 11) {real, imag} */,
  {32'h3fc3b816, 32'hbcb75e80} /* (7, 11, 10) {real, imag} */,
  {32'h3f9a85d5, 32'h3e58f358} /* (7, 11, 9) {real, imag} */,
  {32'hbf544afc, 32'h3f385e5c} /* (7, 11, 8) {real, imag} */,
  {32'hc0230f22, 32'h407a7f9e} /* (7, 11, 7) {real, imag} */,
  {32'h3e9d515a, 32'h3cc32680} /* (7, 11, 6) {real, imag} */,
  {32'hc04dad9f, 32'h4021f2ca} /* (7, 11, 5) {real, imag} */,
  {32'h3c64f700, 32'hbf2d2ae1} /* (7, 11, 4) {real, imag} */,
  {32'hc08d5548, 32'hc09c97c3} /* (7, 11, 3) {real, imag} */,
  {32'h3fa79967, 32'hbf80c294} /* (7, 11, 2) {real, imag} */,
  {32'hc0c8e2b3, 32'hc0f457d5} /* (7, 11, 1) {real, imag} */,
  {32'hbd29e4c0, 32'hc06bc1b1} /* (7, 11, 0) {real, imag} */,
  {32'h3fa8cdfe, 32'h406c6afa} /* (7, 10, 15) {real, imag} */,
  {32'h4026c068, 32'h408e3187} /* (7, 10, 14) {real, imag} */,
  {32'hc0065b65, 32'h40acd0e8} /* (7, 10, 13) {real, imag} */,
  {32'h3f895720, 32'hc08e91b5} /* (7, 10, 12) {real, imag} */,
  {32'h3f0a913c, 32'h40675afa} /* (7, 10, 11) {real, imag} */,
  {32'h3fefd9a2, 32'h400a4020} /* (7, 10, 10) {real, imag} */,
  {32'h3dc3bfe0, 32'h4007efb0} /* (7, 10, 9) {real, imag} */,
  {32'h3f9d5f35, 32'hbf8f2dac} /* (7, 10, 8) {real, imag} */,
  {32'h3f50b1ac, 32'h3fb4a3db} /* (7, 10, 7) {real, imag} */,
  {32'hc016c547, 32'h3e6bd940} /* (7, 10, 6) {real, imag} */,
  {32'hc024bcfb, 32'hbfa8c444} /* (7, 10, 5) {real, imag} */,
  {32'h3f38776b, 32'hbf21a0ee} /* (7, 10, 4) {real, imag} */,
  {32'h403e6c41, 32'hbf11ad40} /* (7, 10, 3) {real, imag} */,
  {32'hbfc8ffe1, 32'hc08ee5fd} /* (7, 10, 2) {real, imag} */,
  {32'h40d2df1c, 32'h4010a620} /* (7, 10, 1) {real, imag} */,
  {32'h402ff814, 32'hc0f38797} /* (7, 10, 0) {real, imag} */,
  {32'h4000670c, 32'hc076e44a} /* (7, 9, 15) {real, imag} */,
  {32'h4004c9a5, 32'h3f998a1c} /* (7, 9, 14) {real, imag} */,
  {32'h3f7855c8, 32'h40208871} /* (7, 9, 13) {real, imag} */,
  {32'hbfc264b3, 32'h3e9bffb9} /* (7, 9, 12) {real, imag} */,
  {32'hbfc3c887, 32'h3e79f1b4} /* (7, 9, 11) {real, imag} */,
  {32'h3efa12d8, 32'h3e196c32} /* (7, 9, 10) {real, imag} */,
  {32'hbf9e4ef0, 32'h3f5c20c0} /* (7, 9, 9) {real, imag} */,
  {32'h3df23ce0, 32'h3eb5d800} /* (7, 9, 8) {real, imag} */,
  {32'hbe95355a, 32'hbe30a190} /* (7, 9, 7) {real, imag} */,
  {32'hbd75d3c0, 32'h3f35a988} /* (7, 9, 6) {real, imag} */,
  {32'hbf71c18e, 32'h3f7b997b} /* (7, 9, 5) {real, imag} */,
  {32'hc09f61f3, 32'hbea06a37} /* (7, 9, 4) {real, imag} */,
  {32'h3f103764, 32'hbfad6106} /* (7, 9, 3) {real, imag} */,
  {32'h40d50cf8, 32'h3e66d1c2} /* (7, 9, 2) {real, imag} */,
  {32'h40b81fa0, 32'hc00be85a} /* (7, 9, 1) {real, imag} */,
  {32'hc057800f, 32'h3fb2fe3e} /* (7, 9, 0) {real, imag} */,
  {32'h40b0b6e5, 32'hbfa95746} /* (7, 8, 15) {real, imag} */,
  {32'h3fdd7e88, 32'h3fe086a3} /* (7, 8, 14) {real, imag} */,
  {32'hbeed412c, 32'h4024a708} /* (7, 8, 13) {real, imag} */,
  {32'h3fdfe339, 32'hc03f3677} /* (7, 8, 12) {real, imag} */,
  {32'h4003ea8d, 32'h3fb33b52} /* (7, 8, 11) {real, imag} */,
  {32'hbfc9fe7b, 32'hbe65101d} /* (7, 8, 10) {real, imag} */,
  {32'hbe98d8c8, 32'h3f365b73} /* (7, 8, 9) {real, imag} */,
  {32'hbd350030, 32'hbf24de0e} /* (7, 8, 8) {real, imag} */,
  {32'h3e0ecaa0, 32'hbf87f4e8} /* (7, 8, 7) {real, imag} */,
  {32'h3d4c30c0, 32'h3e5d5563} /* (7, 8, 6) {real, imag} */,
  {32'hbfe979d2, 32'h3fdbdbf6} /* (7, 8, 5) {real, imag} */,
  {32'h3f6f6c86, 32'hc0522369} /* (7, 8, 4) {real, imag} */,
  {32'h40058a9a, 32'h40511ebc} /* (7, 8, 3) {real, imag} */,
  {32'h404ead68, 32'hbfa2a16b} /* (7, 8, 2) {real, imag} */,
  {32'hbf372308, 32'h3f307ae1} /* (7, 8, 1) {real, imag} */,
  {32'h3fcb7f94, 32'hbfdda871} /* (7, 8, 0) {real, imag} */,
  {32'hc0b5a8c2, 32'h3e1c7a78} /* (7, 7, 15) {real, imag} */,
  {32'hc0c9e48c, 32'h40ae413e} /* (7, 7, 14) {real, imag} */,
  {32'h3f6d862c, 32'hbf8a0869} /* (7, 7, 13) {real, imag} */,
  {32'h406560a4, 32'h4043c1af} /* (7, 7, 12) {real, imag} */,
  {32'hbf1d429c, 32'hc0607978} /* (7, 7, 11) {real, imag} */,
  {32'h3f838d58, 32'hbf5e561f} /* (7, 7, 10) {real, imag} */,
  {32'hbf81ed52, 32'hbffe8f72} /* (7, 7, 9) {real, imag} */,
  {32'hbe7295b0, 32'h3ee1ed84} /* (7, 7, 8) {real, imag} */,
  {32'hbf6d3b2c, 32'hbfdf5e58} /* (7, 7, 7) {real, imag} */,
  {32'h402c4f7c, 32'h3fa82c3c} /* (7, 7, 6) {real, imag} */,
  {32'hc05fddd7, 32'h3f83a83c} /* (7, 7, 5) {real, imag} */,
  {32'h400793d2, 32'h400a2683} /* (7, 7, 4) {real, imag} */,
  {32'h40ad01dc, 32'h3d82a540} /* (7, 7, 3) {real, imag} */,
  {32'hc0018a1c, 32'hc0d9eb62} /* (7, 7, 2) {real, imag} */,
  {32'hbfc50982, 32'hc024189a} /* (7, 7, 1) {real, imag} */,
  {32'h40870cec, 32'h403608a6} /* (7, 7, 0) {real, imag} */,
  {32'hbf8df31b, 32'h3fe5bd6e} /* (7, 6, 15) {real, imag} */,
  {32'h40de516a, 32'h40a7230e} /* (7, 6, 14) {real, imag} */,
  {32'hc0b9167f, 32'hc085b9b6} /* (7, 6, 13) {real, imag} */,
  {32'hc0ac848c, 32'hbe1535c8} /* (7, 6, 12) {real, imag} */,
  {32'h3fc149bc, 32'hbf7ef2d4} /* (7, 6, 11) {real, imag} */,
  {32'h40a613bc, 32'hc08892d3} /* (7, 6, 10) {real, imag} */,
  {32'h3eac28d3, 32'hbddb60e8} /* (7, 6, 9) {real, imag} */,
  {32'h3e709340, 32'h3fbc86ac} /* (7, 6, 8) {real, imag} */,
  {32'hbf21f4ec, 32'h3efb77a6} /* (7, 6, 7) {real, imag} */,
  {32'hc0543e61, 32'h3f06f668} /* (7, 6, 6) {real, imag} */,
  {32'h3fa4381c, 32'h3dd91a30} /* (7, 6, 5) {real, imag} */,
  {32'hc03a517c, 32'hc07e2d64} /* (7, 6, 4) {real, imag} */,
  {32'hc0b03963, 32'hbee55d30} /* (7, 6, 3) {real, imag} */,
  {32'h4069a0bb, 32'hc04dd04f} /* (7, 6, 2) {real, imag} */,
  {32'h4031ceb0, 32'hc0b857a2} /* (7, 6, 1) {real, imag} */,
  {32'h3fbd2a5a, 32'hc10edd8c} /* (7, 6, 0) {real, imag} */,
  {32'h3fccf74e, 32'hc0a53fba} /* (7, 5, 15) {real, imag} */,
  {32'hbfd03a8f, 32'hc0a14bdb} /* (7, 5, 14) {real, imag} */,
  {32'hc0eda3f5, 32'hc0bc9fbe} /* (7, 5, 13) {real, imag} */,
  {32'h40227dc2, 32'h40f4e71b} /* (7, 5, 12) {real, imag} */,
  {32'h408343c6, 32'hbfe142cc} /* (7, 5, 11) {real, imag} */,
  {32'h3f309e01, 32'h3fd94939} /* (7, 5, 10) {real, imag} */,
  {32'h3f7fe664, 32'h3f492e02} /* (7, 5, 9) {real, imag} */,
  {32'hbf42e878, 32'h3f5557bc} /* (7, 5, 8) {real, imag} */,
  {32'h40498a4b, 32'h3fd3abed} /* (7, 5, 7) {real, imag} */,
  {32'hbf40717b, 32'hc0019a53} /* (7, 5, 6) {real, imag} */,
  {32'h403130b7, 32'h4014f33e} /* (7, 5, 5) {real, imag} */,
  {32'hbf4a4636, 32'hbee0d1d0} /* (7, 5, 4) {real, imag} */,
  {32'h3fc6779c, 32'hc0acbd2a} /* (7, 5, 3) {real, imag} */,
  {32'hbf9a8455, 32'h40cc6d47} /* (7, 5, 2) {real, imag} */,
  {32'h410c532f, 32'h400e453e} /* (7, 5, 1) {real, imag} */,
  {32'hc159d26c, 32'hc0429d78} /* (7, 5, 0) {real, imag} */,
  {32'hc19e42d6, 32'h40aada71} /* (7, 4, 15) {real, imag} */,
  {32'h40333936, 32'hc0bee42b} /* (7, 4, 14) {real, imag} */,
  {32'h40190ae4, 32'h40512b1e} /* (7, 4, 13) {real, imag} */,
  {32'hbfc937ac, 32'hc01ea11b} /* (7, 4, 12) {real, imag} */,
  {32'h3fc0a3e4, 32'hc0875fd5} /* (7, 4, 11) {real, imag} */,
  {32'h40012497, 32'hbf12d065} /* (7, 4, 10) {real, imag} */,
  {32'hbcd25800, 32'hbf5bfbd8} /* (7, 4, 9) {real, imag} */,
  {32'h3f985471, 32'hbfcfacfc} /* (7, 4, 8) {real, imag} */,
  {32'hbf82ca90, 32'hbf0392b8} /* (7, 4, 7) {real, imag} */,
  {32'hc049d441, 32'hbd9ef598} /* (7, 4, 6) {real, imag} */,
  {32'hc095550a, 32'hc06459ee} /* (7, 4, 5) {real, imag} */,
  {32'h40028734, 32'h40cc035e} /* (7, 4, 4) {real, imag} */,
  {32'hc0886917, 32'h41082dd8} /* (7, 4, 3) {real, imag} */,
  {32'h403471d4, 32'hc0bc0abd} /* (7, 4, 2) {real, imag} */,
  {32'hc0e087fe, 32'hc18695d8} /* (7, 4, 1) {real, imag} */,
  {32'h408f046d, 32'hbfc0c364} /* (7, 4, 0) {real, imag} */,
  {32'hc18ca5bb, 32'hc00ff8c4} /* (7, 3, 15) {real, imag} */,
  {32'h4105b41d, 32'h41060513} /* (7, 3, 14) {real, imag} */,
  {32'h40c8ea3c, 32'h41081f7c} /* (7, 3, 13) {real, imag} */,
  {32'hc050420c, 32'hc12a04a3} /* (7, 3, 12) {real, imag} */,
  {32'h3f42e3d6, 32'hbf3eb2a1} /* (7, 3, 11) {real, imag} */,
  {32'hc0d7951c, 32'h4001ceba} /* (7, 3, 10) {real, imag} */,
  {32'h3f74c8b6, 32'hc08a7cba} /* (7, 3, 9) {real, imag} */,
  {32'h3f22ed78, 32'hbf5dcd98} /* (7, 3, 8) {real, imag} */,
  {32'h3f5592b6, 32'h3faaac62} /* (7, 3, 7) {real, imag} */,
  {32'hc08e6610, 32'h3f60b1b6} /* (7, 3, 6) {real, imag} */,
  {32'hbf247552, 32'hbf8aa4fc} /* (7, 3, 5) {real, imag} */,
  {32'h4108132c, 32'hbff1a738} /* (7, 3, 4) {real, imag} */,
  {32'h3fe1616e, 32'hc0984574} /* (7, 3, 3) {real, imag} */,
  {32'hc093e20e, 32'hbf9e8250} /* (7, 3, 2) {real, imag} */,
  {32'h40fcd9db, 32'hc06505e6} /* (7, 3, 1) {real, imag} */,
  {32'hc10db11c, 32'h41468722} /* (7, 3, 0) {real, imag} */,
  {32'hc0209ccc, 32'h40f13b9a} /* (7, 2, 15) {real, imag} */,
  {32'h406bbfba, 32'h3f055598} /* (7, 2, 14) {real, imag} */,
  {32'h40ca2abc, 32'hc0dd51a3} /* (7, 2, 13) {real, imag} */,
  {32'hbf83da8a, 32'hc10da558} /* (7, 2, 12) {real, imag} */,
  {32'h410ff534, 32'hbf613ec0} /* (7, 2, 11) {real, imag} */,
  {32'h401c6553, 32'hbe799820} /* (7, 2, 10) {real, imag} */,
  {32'hc013fb8c, 32'h40337f4b} /* (7, 2, 9) {real, imag} */,
  {32'h3fb35e34, 32'hc026a2c8} /* (7, 2, 8) {real, imag} */,
  {32'h3fda8b61, 32'h3f2fddec} /* (7, 2, 7) {real, imag} */,
  {32'h4104517e, 32'hc08bdda9} /* (7, 2, 6) {real, imag} */,
  {32'hc11e22e6, 32'hc0601c74} /* (7, 2, 5) {real, imag} */,
  {32'h3faff662, 32'hc06ed3b2} /* (7, 2, 4) {real, imag} */,
  {32'hc0590458, 32'h3dced5c0} /* (7, 2, 3) {real, imag} */,
  {32'hc18daf9b, 32'h4111b10a} /* (7, 2, 2) {real, imag} */,
  {32'h40f76c50, 32'hc1495d85} /* (7, 2, 1) {real, imag} */,
  {32'hc0b68235, 32'h4064f6d2} /* (7, 2, 0) {real, imag} */,
  {32'hc0534c38, 32'hc073eeb4} /* (7, 1, 15) {real, imag} */,
  {32'h3fd1ce12, 32'h3fe60016} /* (7, 1, 14) {real, imag} */,
  {32'hc140f871, 32'h406ab66d} /* (7, 1, 13) {real, imag} */,
  {32'hc0a26ebc, 32'hc0b2fe9d} /* (7, 1, 12) {real, imag} */,
  {32'hc1156487, 32'hbfd625c8} /* (7, 1, 11) {real, imag} */,
  {32'h3fa5ec2e, 32'h3fc3b974} /* (7, 1, 10) {real, imag} */,
  {32'hbf2c8a40, 32'h403c5fc1} /* (7, 1, 9) {real, imag} */,
  {32'h4009f253, 32'h40514186} /* (7, 1, 8) {real, imag} */,
  {32'h3ee83dc0, 32'h407ffa3b} /* (7, 1, 7) {real, imag} */,
  {32'hc10d11ab, 32'h3fe21e1c} /* (7, 1, 6) {real, imag} */,
  {32'h41478243, 32'h4145fd3f} /* (7, 1, 5) {real, imag} */,
  {32'h3fd4aaa2, 32'h416374ae} /* (7, 1, 4) {real, imag} */,
  {32'hc166f3c7, 32'hc0b5324a} /* (7, 1, 3) {real, imag} */,
  {32'h3f9d8f2a, 32'h3f1a564d} /* (7, 1, 2) {real, imag} */,
  {32'h41c84b0e, 32'h41066ae1} /* (7, 1, 1) {real, imag} */,
  {32'hbfc1255a, 32'hc1419d94} /* (7, 1, 0) {real, imag} */,
  {32'hc1330a6a, 32'h416b42d4} /* (7, 0, 15) {real, imag} */,
  {32'h40d970f4, 32'hbf4a83c8} /* (7, 0, 14) {real, imag} */,
  {32'hc087eb9c, 32'hc185f596} /* (7, 0, 13) {real, imag} */,
  {32'hbef8f128, 32'h4091abf8} /* (7, 0, 12) {real, imag} */,
  {32'h3ee47f70, 32'h411b3a54} /* (7, 0, 11) {real, imag} */,
  {32'hbe3085b0, 32'hbfeb3a3c} /* (7, 0, 10) {real, imag} */,
  {32'h401265d2, 32'h3f4bcbec} /* (7, 0, 9) {real, imag} */,
  {32'hc0d3aaaa, 32'hc090d97e} /* (7, 0, 8) {real, imag} */,
  {32'h40ac2455, 32'h3f907742} /* (7, 0, 7) {real, imag} */,
  {32'h40068261, 32'hc136496e} /* (7, 0, 6) {real, imag} */,
  {32'hc11a3128, 32'hbfd3b280} /* (7, 0, 5) {real, imag} */,
  {32'hc08a5298, 32'hbf45f76c} /* (7, 0, 4) {real, imag} */,
  {32'h418ffd1b, 32'h3d930980} /* (7, 0, 3) {real, imag} */,
  {32'hc12b0db2, 32'h413bffb4} /* (7, 0, 2) {real, imag} */,
  {32'h41867d91, 32'h4124878c} /* (7, 0, 1) {real, imag} */,
  {32'h40901c58, 32'h419b0e22} /* (7, 0, 0) {real, imag} */,
  {32'hc0bddb56, 32'hc0aadc87} /* (6, 15, 15) {real, imag} */,
  {32'h41a86fb9, 32'h41a12d4e} /* (6, 15, 14) {real, imag} */,
  {32'hc17c6462, 32'h4186d76f} /* (6, 15, 13) {real, imag} */,
  {32'hc0af07ed, 32'hbecb3d60} /* (6, 15, 12) {real, imag} */,
  {32'h403c1d90, 32'hc0a0f5ba} /* (6, 15, 11) {real, imag} */,
  {32'hbf7bcf58, 32'h3f52e09e} /* (6, 15, 10) {real, imag} */,
  {32'h405373d4, 32'hc0d66806} /* (6, 15, 9) {real, imag} */,
  {32'hbfc4b558, 32'hc067f470} /* (6, 15, 8) {real, imag} */,
  {32'h416edd7f, 32'h3fc4747e} /* (6, 15, 7) {real, imag} */,
  {32'h408c355b, 32'hbf132fbe} /* (6, 15, 6) {real, imag} */,
  {32'h3ffb551c, 32'h405e5bc8} /* (6, 15, 5) {real, imag} */,
  {32'hc0bfa5b7, 32'hc061ab24} /* (6, 15, 4) {real, imag} */,
  {32'h3f1206a0, 32'hc1041f2a} /* (6, 15, 3) {real, imag} */,
  {32'h400a2a78, 32'h41da7942} /* (6, 15, 2) {real, imag} */,
  {32'h41cd9f92, 32'hc03ae78a} /* (6, 15, 1) {real, imag} */,
  {32'hc1ff0e1e, 32'h41867730} /* (6, 15, 0) {real, imag} */,
  {32'hc100b01c, 32'h410428ee} /* (6, 14, 15) {real, imag} */,
  {32'hc0efe241, 32'hc1add86a} /* (6, 14, 14) {real, imag} */,
  {32'hbf773770, 32'hc10c1db0} /* (6, 14, 13) {real, imag} */,
  {32'h408cb911, 32'h410f02c2} /* (6, 14, 12) {real, imag} */,
  {32'hc1345d14, 32'h407225e8} /* (6, 14, 11) {real, imag} */,
  {32'hc0d1e7af, 32'h3edc98e0} /* (6, 14, 10) {real, imag} */,
  {32'h40129d2a, 32'h407c4f68} /* (6, 14, 9) {real, imag} */,
  {32'h40fe3890, 32'hc0164204} /* (6, 14, 8) {real, imag} */,
  {32'hc0f13811, 32'hbddebf80} /* (6, 14, 7) {real, imag} */,
  {32'hbff3a8d4, 32'hc10f8e29} /* (6, 14, 6) {real, imag} */,
  {32'hc0650ba8, 32'h40a33fd8} /* (6, 14, 5) {real, imag} */,
  {32'h413bd2b0, 32'hc12eb786} /* (6, 14, 4) {real, imag} */,
  {32'h40fc57e6, 32'hbf167a00} /* (6, 14, 3) {real, imag} */,
  {32'hc0090f26, 32'h40b612ae} /* (6, 14, 2) {real, imag} */,
  {32'h41818f70, 32'h409714b2} /* (6, 14, 1) {real, imag} */,
  {32'h40b53228, 32'h40f52cbc} /* (6, 14, 0) {real, imag} */,
  {32'h41a90053, 32'hc117ad65} /* (6, 13, 15) {real, imag} */,
  {32'hc0bbf0fa, 32'h4104468b} /* (6, 13, 14) {real, imag} */,
  {32'hc0c35aec, 32'h419cdb18} /* (6, 13, 13) {real, imag} */,
  {32'hc0ca9d94, 32'h408d3221} /* (6, 13, 12) {real, imag} */,
  {32'h418a2b6b, 32'h400a43ac} /* (6, 13, 11) {real, imag} */,
  {32'h40221422, 32'hc03a9c5a} /* (6, 13, 10) {real, imag} */,
  {32'h3f6e2898, 32'h4060774c} /* (6, 13, 9) {real, imag} */,
  {32'h3e08e3c0, 32'h3f47f2a0} /* (6, 13, 8) {real, imag} */,
  {32'hc05f7a56, 32'h3fa6c068} /* (6, 13, 7) {real, imag} */,
  {32'h403acec6, 32'hc0acbcdf} /* (6, 13, 6) {real, imag} */,
  {32'h3fe30ccc, 32'hc03dab8c} /* (6, 13, 5) {real, imag} */,
  {32'hbfebcf52, 32'hc1897145} /* (6, 13, 4) {real, imag} */,
  {32'h40e3ee26, 32'h40d17a48} /* (6, 13, 3) {real, imag} */,
  {32'h41846a80, 32'hc1674e15} /* (6, 13, 2) {real, imag} */,
  {32'h415ffe46, 32'hc027d9ac} /* (6, 13, 1) {real, imag} */,
  {32'hc188372c, 32'hc19b2bab} /* (6, 13, 0) {real, imag} */,
  {32'hbfebc1d8, 32'hc141fc76} /* (6, 12, 15) {real, imag} */,
  {32'h3fac666f, 32'h3ecf99a0} /* (6, 12, 14) {real, imag} */,
  {32'hc1236317, 32'hc099f366} /* (6, 12, 13) {real, imag} */,
  {32'hbf303d20, 32'hc11c9fd0} /* (6, 12, 12) {real, imag} */,
  {32'h40d86718, 32'h415d3c77} /* (6, 12, 11) {real, imag} */,
  {32'hc044e00b, 32'hc0dcd992} /* (6, 12, 10) {real, imag} */,
  {32'h3fe501b8, 32'h4019403c} /* (6, 12, 9) {real, imag} */,
  {32'h40828cb3, 32'hbfdbd5f8} /* (6, 12, 8) {real, imag} */,
  {32'hc06cfea4, 32'h406778fc} /* (6, 12, 7) {real, imag} */,
  {32'h4019cfc1, 32'h3e1cb5b0} /* (6, 12, 6) {real, imag} */,
  {32'hbede6e08, 32'hc066404c} /* (6, 12, 5) {real, imag} */,
  {32'h4112059c, 32'hc1398500} /* (6, 12, 4) {real, imag} */,
  {32'hc1b3a10e, 32'hc1289ddd} /* (6, 12, 3) {real, imag} */,
  {32'h4019392a, 32'h412b76c7} /* (6, 12, 2) {real, imag} */,
  {32'hc1bc1522, 32'hc0fbab94} /* (6, 12, 1) {real, imag} */,
  {32'h410f895e, 32'h4186b870} /* (6, 12, 0) {real, imag} */,
  {32'h3fe41ac1, 32'h409cb758} /* (6, 11, 15) {real, imag} */,
  {32'hc09625fe, 32'h3f82e04c} /* (6, 11, 14) {real, imag} */,
  {32'hc094ea1d, 32'h41027d81} /* (6, 11, 13) {real, imag} */,
  {32'hbfa848c8, 32'h40903e1e} /* (6, 11, 12) {real, imag} */,
  {32'h408f4326, 32'h40379946} /* (6, 11, 11) {real, imag} */,
  {32'hc07c30eb, 32'hc0127a0a} /* (6, 11, 10) {real, imag} */,
  {32'hbfc3e00d, 32'hbf8dbfc2} /* (6, 11, 9) {real, imag} */,
  {32'hbfd97fba, 32'h402342d1} /* (6, 11, 8) {real, imag} */,
  {32'h40118272, 32'hc0caf874} /* (6, 11, 7) {real, imag} */,
  {32'hbfc8c18e, 32'h40be596d} /* (6, 11, 6) {real, imag} */,
  {32'hc014f1ef, 32'h4073eb16} /* (6, 11, 5) {real, imag} */,
  {32'h403664da, 32'hc145e819} /* (6, 11, 4) {real, imag} */,
  {32'hc14fb29e, 32'h3fb369d0} /* (6, 11, 3) {real, imag} */,
  {32'hc000844f, 32'h40a58ba9} /* (6, 11, 2) {real, imag} */,
  {32'hbfe30d4f, 32'hc11964be} /* (6, 11, 1) {real, imag} */,
  {32'h410f7f01, 32'h40eca824} /* (6, 11, 0) {real, imag} */,
  {32'h40e0603c, 32'h3e8eea6c} /* (6, 10, 15) {real, imag} */,
  {32'hc13f308c, 32'hbfde054e} /* (6, 10, 14) {real, imag} */,
  {32'hc0802df6, 32'h407ebe59} /* (6, 10, 13) {real, imag} */,
  {32'h41623416, 32'hbec569e8} /* (6, 10, 12) {real, imag} */,
  {32'hc041f0c8, 32'hbeede658} /* (6, 10, 11) {real, imag} */,
  {32'h409d6d1b, 32'h3ee47e50} /* (6, 10, 10) {real, imag} */,
  {32'hbfe9e63a, 32'hc082171a} /* (6, 10, 9) {real, imag} */,
  {32'hc00d6fe7, 32'h3fd1fb06} /* (6, 10, 8) {real, imag} */,
  {32'h4058766b, 32'h3f9308ff} /* (6, 10, 7) {real, imag} */,
  {32'h3fc8f1cc, 32'h406d8878} /* (6, 10, 6) {real, imag} */,
  {32'hc0ea1a00, 32'h3f56296c} /* (6, 10, 5) {real, imag} */,
  {32'hbf3a5780, 32'h4077eb39} /* (6, 10, 4) {real, imag} */,
  {32'h4082e03a, 32'hc0c486dc} /* (6, 10, 3) {real, imag} */,
  {32'hc0cf69c9, 32'hc0514d7f} /* (6, 10, 2) {real, imag} */,
  {32'hc103ebea, 32'h3c9b76c0} /* (6, 10, 1) {real, imag} */,
  {32'hbfcd3152, 32'hc01cb907} /* (6, 10, 0) {real, imag} */,
  {32'hc0b87ea2, 32'h3ff1b665} /* (6, 9, 15) {real, imag} */,
  {32'h3f041cf2, 32'hbfc2b22c} /* (6, 9, 14) {real, imag} */,
  {32'hc0b9450b, 32'hc10eb300} /* (6, 9, 13) {real, imag} */,
  {32'h3fdb75d8, 32'hbff2acac} /* (6, 9, 12) {real, imag} */,
  {32'h3fdd2842, 32'hbeb2086c} /* (6, 9, 11) {real, imag} */,
  {32'h3fb06352, 32'h405950bb} /* (6, 9, 10) {real, imag} */,
  {32'hbf6b827f, 32'h3eb64d98} /* (6, 9, 9) {real, imag} */,
  {32'h3e832cd0, 32'hbf8aa0e8} /* (6, 9, 8) {real, imag} */,
  {32'h3bf5bc80, 32'h3f064768} /* (6, 9, 7) {real, imag} */,
  {32'hbdf65d08, 32'h3e070730} /* (6, 9, 6) {real, imag} */,
  {32'hbfcc2e96, 32'h3f7378aa} /* (6, 9, 5) {real, imag} */,
  {32'h3e55b6ec, 32'h40da5915} /* (6, 9, 4) {real, imag} */,
  {32'h3e4e5c60, 32'h3f497b48} /* (6, 9, 3) {real, imag} */,
  {32'hc061770c, 32'hc107ca5a} /* (6, 9, 2) {real, imag} */,
  {32'h3fe23486, 32'h407622fe} /* (6, 9, 1) {real, imag} */,
  {32'h40aa46af, 32'h405ea30c} /* (6, 9, 0) {real, imag} */,
  {32'hc0825a96, 32'hbf2ef71b} /* (6, 8, 15) {real, imag} */,
  {32'h3fd705ea, 32'h4007a732} /* (6, 8, 14) {real, imag} */,
  {32'h3cfef780, 32'h3fd0e2a6} /* (6, 8, 13) {real, imag} */,
  {32'hbf7c780b, 32'hbfb1677b} /* (6, 8, 12) {real, imag} */,
  {32'h40414102, 32'hbf5d089e} /* (6, 8, 11) {real, imag} */,
  {32'h3f322fb2, 32'hbfc85634} /* (6, 8, 10) {real, imag} */,
  {32'h3c958d40, 32'h3f8b7eb5} /* (6, 8, 9) {real, imag} */,
  {32'hbe5e2440, 32'hbf0ff5fe} /* (6, 8, 8) {real, imag} */,
  {32'h3fa4de91, 32'h3f1b3e7c} /* (6, 8, 7) {real, imag} */,
  {32'h40415a24, 32'h3f9bd30c} /* (6, 8, 6) {real, imag} */,
  {32'hc0158cc2, 32'hc05ab94e} /* (6, 8, 5) {real, imag} */,
  {32'h3f5c6b11, 32'h402a9884} /* (6, 8, 4) {real, imag} */,
  {32'hbfe6658c, 32'hc09fc4ea} /* (6, 8, 3) {real, imag} */,
  {32'hc05fa027, 32'h40d2683d} /* (6, 8, 2) {real, imag} */,
  {32'h40d98366, 32'h3fdcdcaa} /* (6, 8, 1) {real, imag} */,
  {32'h40333762, 32'h4083b770} /* (6, 8, 0) {real, imag} */,
  {32'hbf021920, 32'hbf98f58c} /* (6, 7, 15) {real, imag} */,
  {32'hbf4312c0, 32'hbf741c94} /* (6, 7, 14) {real, imag} */,
  {32'h40f09107, 32'hc1155e55} /* (6, 7, 13) {real, imag} */,
  {32'h3e142158, 32'hc00ec860} /* (6, 7, 12) {real, imag} */,
  {32'h3fbabb1a, 32'h401e6314} /* (6, 7, 11) {real, imag} */,
  {32'hbfbc7c17, 32'h3f855e80} /* (6, 7, 10) {real, imag} */,
  {32'hbfbf3f23, 32'hbf7260fc} /* (6, 7, 9) {real, imag} */,
  {32'h400625ea, 32'hbfe0f512} /* (6, 7, 8) {real, imag} */,
  {32'hbe8a985c, 32'h3fa5129e} /* (6, 7, 7) {real, imag} */,
  {32'h3fab3535, 32'h3f2116e5} /* (6, 7, 6) {real, imag} */,
  {32'h3f9ec7fa, 32'hc0c30988} /* (6, 7, 5) {real, imag} */,
  {32'hc028e89a, 32'h3fb6faa7} /* (6, 7, 4) {real, imag} */,
  {32'hc0b0b691, 32'hbfaf6eb0} /* (6, 7, 3) {real, imag} */,
  {32'hc097525a, 32'h408930dc} /* (6, 7, 2) {real, imag} */,
  {32'hc0b34412, 32'h3e26b95c} /* (6, 7, 1) {real, imag} */,
  {32'h40d7c4d7, 32'hbfffa2e4} /* (6, 7, 0) {real, imag} */,
  {32'hc0b80b98, 32'hc0e34cf9} /* (6, 6, 15) {real, imag} */,
  {32'hc0932572, 32'h40075508} /* (6, 6, 14) {real, imag} */,
  {32'hc046bff6, 32'hbfdae669} /* (6, 6, 13) {real, imag} */,
  {32'h409715fc, 32'h40d2b00b} /* (6, 6, 12) {real, imag} */,
  {32'hbf18ee32, 32'h4081ea6a} /* (6, 6, 11) {real, imag} */,
  {32'h3fe39c34, 32'hc007db5c} /* (6, 6, 10) {real, imag} */,
  {32'h4010f8b2, 32'h3f1e7fbc} /* (6, 6, 9) {real, imag} */,
  {32'h3f208be8, 32'h3f7ddaa8} /* (6, 6, 8) {real, imag} */,
  {32'hbe733d98, 32'hbf83adfa} /* (6, 6, 7) {real, imag} */,
  {32'h405b48d4, 32'h3fd71954} /* (6, 6, 6) {real, imag} */,
  {32'h400528fe, 32'h3eafc518} /* (6, 6, 5) {real, imag} */,
  {32'hbfe6aed6, 32'h40b872c1} /* (6, 6, 4) {real, imag} */,
  {32'hbe85ccc4, 32'h3f45a926} /* (6, 6, 3) {real, imag} */,
  {32'h41053587, 32'hc0f27f70} /* (6, 6, 2) {real, imag} */,
  {32'h408af368, 32'hc0894f6f} /* (6, 6, 1) {real, imag} */,
  {32'hc1480b10, 32'hc08e093d} /* (6, 6, 0) {real, imag} */,
  {32'h3f688a80, 32'hbf7eebec} /* (6, 5, 15) {real, imag} */,
  {32'h3f6a0e3e, 32'hc1168ef7} /* (6, 5, 14) {real, imag} */,
  {32'hbf947890, 32'h418b05ea} /* (6, 5, 13) {real, imag} */,
  {32'hc03f76a5, 32'hc110e6f2} /* (6, 5, 12) {real, imag} */,
  {32'h3fc36e9d, 32'h3f3df0f8} /* (6, 5, 11) {real, imag} */,
  {32'h3fe26090, 32'h3fae5ee1} /* (6, 5, 10) {real, imag} */,
  {32'hbfab091e, 32'hbff75101} /* (6, 5, 9) {real, imag} */,
  {32'hbff54976, 32'h4000cee4} /* (6, 5, 8) {real, imag} */,
  {32'hc063f96f, 32'hc0ab168a} /* (6, 5, 7) {real, imag} */,
  {32'hc08892ba, 32'h402f6838} /* (6, 5, 6) {real, imag} */,
  {32'h3e3e33e8, 32'h411451c0} /* (6, 5, 5) {real, imag} */,
  {32'hc10a51e3, 32'h402018d6} /* (6, 5, 4) {real, imag} */,
  {32'h41262032, 32'hc0e575c8} /* (6, 5, 3) {real, imag} */,
  {32'hbf4fea7e, 32'hc1866600} /* (6, 5, 2) {real, imag} */,
  {32'h41541f8a, 32'h3ee87610} /* (6, 5, 1) {real, imag} */,
  {32'h4096a548, 32'h4150c93f} /* (6, 5, 0) {real, imag} */,
  {32'h41694776, 32'hc1643f6d} /* (6, 4, 15) {real, imag} */,
  {32'hc169c612, 32'h40b637fa} /* (6, 4, 14) {real, imag} */,
  {32'hc044d245, 32'h3fcfaabe} /* (6, 4, 13) {real, imag} */,
  {32'h40963faf, 32'h3f6e8138} /* (6, 4, 12) {real, imag} */,
  {32'hc06c2516, 32'h3eb96218} /* (6, 4, 11) {real, imag} */,
  {32'hc0bbf46a, 32'h3fb32d68} /* (6, 4, 10) {real, imag} */,
  {32'h3e212980, 32'hc039255e} /* (6, 4, 9) {real, imag} */,
  {32'h3f219ee8, 32'hc0e04612} /* (6, 4, 8) {real, imag} */,
  {32'hc027bca0, 32'hbffe8ccc} /* (6, 4, 7) {real, imag} */,
  {32'h4062ea50, 32'h3ff74b08} /* (6, 4, 6) {real, imag} */,
  {32'h3febed7f, 32'hbfdeb84e} /* (6, 4, 5) {real, imag} */,
  {32'hc189c87e, 32'hbf5b8f48} /* (6, 4, 4) {real, imag} */,
  {32'hc06abf9f, 32'hc0c2b944} /* (6, 4, 3) {real, imag} */,
  {32'h4174dca6, 32'h41675579} /* (6, 4, 2) {real, imag} */,
  {32'h4150f488, 32'h40678b54} /* (6, 4, 1) {real, imag} */,
  {32'hc122826a, 32'h40ff0d34} /* (6, 4, 0) {real, imag} */,
  {32'hc1044736, 32'hc0bad9e8} /* (6, 3, 15) {real, imag} */,
  {32'hbecd5f80, 32'h400327e0} /* (6, 3, 14) {real, imag} */,
  {32'h40cbff00, 32'h419210b2} /* (6, 3, 13) {real, imag} */,
  {32'h41092080, 32'h405b7fb5} /* (6, 3, 12) {real, imag} */,
  {32'h3f88b9e1, 32'hc05ba004} /* (6, 3, 11) {real, imag} */,
  {32'hbfe79c5a, 32'h40220f96} /* (6, 3, 10) {real, imag} */,
  {32'hbf895419, 32'h40481b98} /* (6, 3, 9) {real, imag} */,
  {32'hbf2a9be7, 32'h400558d0} /* (6, 3, 8) {real, imag} */,
  {32'h404b2912, 32'h402f2578} /* (6, 3, 7) {real, imag} */,
  {32'hc094e50a, 32'hbe590380} /* (6, 3, 6) {real, imag} */,
  {32'h3ffda861, 32'h401bd498} /* (6, 3, 5) {real, imag} */,
  {32'h4104ef34, 32'h40b40414} /* (6, 3, 4) {real, imag} */,
  {32'hc1443bd8, 32'h40f7fab7} /* (6, 3, 3) {real, imag} */,
  {32'h3fb045a4, 32'h41494e8e} /* (6, 3, 2) {real, imag} */,
  {32'hbfd78bfa, 32'hc14c31a0} /* (6, 3, 1) {real, imag} */,
  {32'hbdde5f48, 32'hc19e6910} /* (6, 3, 0) {real, imag} */,
  {32'h41ab9919, 32'h4185589c} /* (6, 2, 15) {real, imag} */,
  {32'hc1ba6f15, 32'hc0496143} /* (6, 2, 14) {real, imag} */,
  {32'h4112a18b, 32'h3f515188} /* (6, 2, 13) {real, imag} */,
  {32'h3fe9475c, 32'h414c665f} /* (6, 2, 12) {real, imag} */,
  {32'hc0f92f40, 32'hbf94e0f0} /* (6, 2, 11) {real, imag} */,
  {32'h4013b0ec, 32'hc074010f} /* (6, 2, 10) {real, imag} */,
  {32'hc00a028e, 32'h3e7f8058} /* (6, 2, 9) {real, imag} */,
  {32'h3fdc5610, 32'h400fd300} /* (6, 2, 8) {real, imag} */,
  {32'h4094e1b5, 32'h401009e2} /* (6, 2, 7) {real, imag} */,
  {32'hbf9653c0, 32'hc00ae8fb} /* (6, 2, 6) {real, imag} */,
  {32'h413c3ff0, 32'h4133f540} /* (6, 2, 5) {real, imag} */,
  {32'hc108e3c6, 32'hc1b51e84} /* (6, 2, 4) {real, imag} */,
  {32'h4175949b, 32'hc0885af4} /* (6, 2, 3) {real, imag} */,
  {32'hc0bc8a24, 32'h40c99808} /* (6, 2, 2) {real, imag} */,
  {32'hc23f251e, 32'h411f54fb} /* (6, 2, 1) {real, imag} */,
  {32'h41de3027, 32'h41a82527} /* (6, 2, 0) {real, imag} */,
  {32'hc13c7ea6, 32'h41232252} /* (6, 1, 15) {real, imag} */,
  {32'hc1ef4cf2, 32'h407a52ec} /* (6, 1, 14) {real, imag} */,
  {32'hc1671223, 32'h41a8e071} /* (6, 1, 13) {real, imag} */,
  {32'h41a6063c, 32'h41bde7db} /* (6, 1, 12) {real, imag} */,
  {32'hc05e8e0d, 32'h408fb771} /* (6, 1, 11) {real, imag} */,
  {32'hc0ae8f12, 32'hc0de64d2} /* (6, 1, 10) {real, imag} */,
  {32'h405cb852, 32'h4063fad5} /* (6, 1, 9) {real, imag} */,
  {32'hc0253858, 32'hc0521d28} /* (6, 1, 8) {real, imag} */,
  {32'hbf9c4938, 32'h3ff21d4a} /* (6, 1, 7) {real, imag} */,
  {32'h4151b8e3, 32'h40939b26} /* (6, 1, 6) {real, imag} */,
  {32'h40ab53c8, 32'h4139cfe4} /* (6, 1, 5) {real, imag} */,
  {32'h3fc2e7d8, 32'hc056b0d8} /* (6, 1, 4) {real, imag} */,
  {32'h40622464, 32'h420572c7} /* (6, 1, 3) {real, imag} */,
  {32'hc0d79028, 32'h4029f6ea} /* (6, 1, 2) {real, imag} */,
  {32'h41012070, 32'hc10a3ac0} /* (6, 1, 1) {real, imag} */,
  {32'h42015d2e, 32'hc10420ce} /* (6, 1, 0) {real, imag} */,
  {32'h412472e6, 32'hc17241d2} /* (6, 0, 15) {real, imag} */,
  {32'h41f272fb, 32'h40d97dde} /* (6, 0, 14) {real, imag} */,
  {32'hc0ed6d86, 32'hc167cb4a} /* (6, 0, 13) {real, imag} */,
  {32'hc14b4386, 32'hc1420c38} /* (6, 0, 12) {real, imag} */,
  {32'hc0d74ade, 32'h40096aad} /* (6, 0, 11) {real, imag} */,
  {32'h40dfc94e, 32'h3f7eb872} /* (6, 0, 10) {real, imag} */,
  {32'hbf0cac6c, 32'h3fe03491} /* (6, 0, 9) {real, imag} */,
  {32'hc063a188, 32'hc0354954} /* (6, 0, 8) {real, imag} */,
  {32'hc01110cd, 32'h3fb4a0ef} /* (6, 0, 7) {real, imag} */,
  {32'hc0a0bc9a, 32'h401a59bc} /* (6, 0, 6) {real, imag} */,
  {32'hc113954b, 32'hbf9fa0ea} /* (6, 0, 5) {real, imag} */,
  {32'h4099b06f, 32'h405856da} /* (6, 0, 4) {real, imag} */,
  {32'hc0e3a5ce, 32'h4010d590} /* (6, 0, 3) {real, imag} */,
  {32'hc1d779ef, 32'hc18f715e} /* (6, 0, 2) {real, imag} */,
  {32'h40377f9b, 32'hc108968e} /* (6, 0, 1) {real, imag} */,
  {32'h401f39a4, 32'h40de6032} /* (6, 0, 0) {real, imag} */,
  {32'h41335302, 32'hc18f2f24} /* (5, 15, 15) {real, imag} */,
  {32'hc0816428, 32'hbfcc92d7} /* (5, 15, 14) {real, imag} */,
  {32'h41207495, 32'hc0bdd28f} /* (5, 15, 13) {real, imag} */,
  {32'h3ff1f930, 32'hc07a0f5e} /* (5, 15, 12) {real, imag} */,
  {32'hc1c27f75, 32'h41562e2c} /* (5, 15, 11) {real, imag} */,
  {32'h41b23b8f, 32'hc0650d1a} /* (5, 15, 10) {real, imag} */,
  {32'h40966f60, 32'hbfd5aadc} /* (5, 15, 9) {real, imag} */,
  {32'hbeffd970, 32'hbfe3493c} /* (5, 15, 8) {real, imag} */,
  {32'h4006303c, 32'h4066e28e} /* (5, 15, 7) {real, imag} */,
  {32'hc02bafa0, 32'h400c922e} /* (5, 15, 6) {real, imag} */,
  {32'hbf01ad60, 32'hc130be14} /* (5, 15, 5) {real, imag} */,
  {32'h41a121a3, 32'h418b8dfa} /* (5, 15, 4) {real, imag} */,
  {32'hc09bbdf8, 32'hc16dbf20} /* (5, 15, 3) {real, imag} */,
  {32'h41c1c459, 32'hc049767a} /* (5, 15, 2) {real, imag} */,
  {32'h41a57cbf, 32'h40b17f2e} /* (5, 15, 1) {real, imag} */,
  {32'h4147a58c, 32'hc1028a20} /* (5, 15, 0) {real, imag} */,
  {32'h3ff52c20, 32'hc191431f} /* (5, 14, 15) {real, imag} */,
  {32'hc1830cec, 32'hc1623a4a} /* (5, 14, 14) {real, imag} */,
  {32'hc1410518, 32'hc1b821c7} /* (5, 14, 13) {real, imag} */,
  {32'h409a6d38, 32'h419c6b26} /* (5, 14, 12) {real, imag} */,
  {32'hbffc74dc, 32'h40a98b6e} /* (5, 14, 11) {real, imag} */,
  {32'hc151cf36, 32'hc0d90da8} /* (5, 14, 10) {real, imag} */,
  {32'h413cfa52, 32'h4188fa2c} /* (5, 14, 9) {real, imag} */,
  {32'h40c02e46, 32'hc010f702} /* (5, 14, 8) {real, imag} */,
  {32'hbfa0e9c0, 32'hc080d47c} /* (5, 14, 7) {real, imag} */,
  {32'h4183341f, 32'h41132570} /* (5, 14, 6) {real, imag} */,
  {32'h41286d96, 32'h418b1232} /* (5, 14, 5) {real, imag} */,
  {32'hc00043ac, 32'h415c302f} /* (5, 14, 4) {real, imag} */,
  {32'hc1922c3b, 32'hc1df0975} /* (5, 14, 3) {real, imag} */,
  {32'h4018aa02, 32'h419cc161} /* (5, 14, 2) {real, imag} */,
  {32'h417539d2, 32'hc0ae25c0} /* (5, 14, 1) {real, imag} */,
  {32'hbfd31e78, 32'h416587b0} /* (5, 14, 0) {real, imag} */,
  {32'h412d3f6b, 32'h41438168} /* (5, 13, 15) {real, imag} */,
  {32'hc15f1702, 32'hc0e63d9c} /* (5, 13, 14) {real, imag} */,
  {32'h40ee78bc, 32'hc14fe35a} /* (5, 13, 13) {real, imag} */,
  {32'h40bf5648, 32'hc12d6c92} /* (5, 13, 12) {real, imag} */,
  {32'h415a5e27, 32'h409f8094} /* (5, 13, 11) {real, imag} */,
  {32'hc0244db6, 32'hc094d651} /* (5, 13, 10) {real, imag} */,
  {32'h3fbd4e28, 32'h4037217e} /* (5, 13, 9) {real, imag} */,
  {32'h3f4a7c04, 32'h3f1eec2c} /* (5, 13, 8) {real, imag} */,
  {32'hbebe6bd0, 32'hbf2b1f12} /* (5, 13, 7) {real, imag} */,
  {32'hc11f2b3c, 32'h3feb4fa4} /* (5, 13, 6) {real, imag} */,
  {32'h40e18266, 32'h4106126e} /* (5, 13, 5) {real, imag} */,
  {32'hc03d32bf, 32'hc157690e} /* (5, 13, 4) {real, imag} */,
  {32'h40de663a, 32'h4153d80e} /* (5, 13, 3) {real, imag} */,
  {32'h419d5b8f, 32'hc1e214b3} /* (5, 13, 2) {real, imag} */,
  {32'hc0d5c1aa, 32'h3fe8f314} /* (5, 13, 1) {real, imag} */,
  {32'hc0c5156e, 32'h403f245d} /* (5, 13, 0) {real, imag} */,
  {32'h4061df5a, 32'hbff2cbeb} /* (5, 12, 15) {real, imag} */,
  {32'h41a62a77, 32'hc13a92c8} /* (5, 12, 14) {real, imag} */,
  {32'h4093d191, 32'h410a8c8c} /* (5, 12, 13) {real, imag} */,
  {32'h41272e8b, 32'h3e800e10} /* (5, 12, 12) {real, imag} */,
  {32'hc00158be, 32'hc10635e0} /* (5, 12, 11) {real, imag} */,
  {32'h3fffadd8, 32'h4106bb20} /* (5, 12, 10) {real, imag} */,
  {32'hc0d4e9d2, 32'h40327698} /* (5, 12, 9) {real, imag} */,
  {32'h401bc6bc, 32'h40a26b7c} /* (5, 12, 8) {real, imag} */,
  {32'hc08afbec, 32'hc09d5916} /* (5, 12, 7) {real, imag} */,
  {32'h40c6700e, 32'hc102db9c} /* (5, 12, 6) {real, imag} */,
  {32'hc10ed4ec, 32'h4134b198} /* (5, 12, 5) {real, imag} */,
  {32'hc08422e6, 32'hc0cb14bc} /* (5, 12, 4) {real, imag} */,
  {32'h408d16ef, 32'h40f22bf1} /* (5, 12, 3) {real, imag} */,
  {32'hc1a97e67, 32'hbfcd6224} /* (5, 12, 2) {real, imag} */,
  {32'hc10b8888, 32'hc0130dc6} /* (5, 12, 1) {real, imag} */,
  {32'h414b867d, 32'h4106781c} /* (5, 12, 0) {real, imag} */,
  {32'h3fd5e242, 32'h40d94058} /* (5, 11, 15) {real, imag} */,
  {32'hc12faf87, 32'hc16b5dee} /* (5, 11, 14) {real, imag} */,
  {32'hbf686e7a, 32'h40268a6a} /* (5, 11, 13) {real, imag} */,
  {32'hc0a15dca, 32'h410fd5ef} /* (5, 11, 12) {real, imag} */,
  {32'hbfcda008, 32'h409d8ce1} /* (5, 11, 11) {real, imag} */,
  {32'h3ead8150, 32'h3ee09b90} /* (5, 11, 10) {real, imag} */,
  {32'h3f97d591, 32'hc0607956} /* (5, 11, 9) {real, imag} */,
  {32'hc031d19b, 32'hbff04d3e} /* (5, 11, 8) {real, imag} */,
  {32'hbecf2478, 32'hc07aa596} /* (5, 11, 7) {real, imag} */,
  {32'hc0d7cd2c, 32'h3f1fb718} /* (5, 11, 6) {real, imag} */,
  {32'h40eeb1c6, 32'hc0683932} /* (5, 11, 5) {real, imag} */,
  {32'h3fa36e9c, 32'h40af0a34} /* (5, 11, 4) {real, imag} */,
  {32'h3f88ebc3, 32'h41310452} /* (5, 11, 3) {real, imag} */,
  {32'hc05697dd, 32'hc1e77b99} /* (5, 11, 2) {real, imag} */,
  {32'h403ce8ab, 32'h410d3299} /* (5, 11, 1) {real, imag} */,
  {32'h4127b3ee, 32'hc0efb456} /* (5, 11, 0) {real, imag} */,
  {32'hc0ef5369, 32'h40be0670} /* (5, 10, 15) {real, imag} */,
  {32'h408d9132, 32'h41169927} /* (5, 10, 14) {real, imag} */,
  {32'h4083d7c8, 32'h40d2f894} /* (5, 10, 13) {real, imag} */,
  {32'hc04e1a8d, 32'h4076c845} /* (5, 10, 12) {real, imag} */,
  {32'h409f88a7, 32'h4028a3d6} /* (5, 10, 11) {real, imag} */,
  {32'h3f869436, 32'hbe6d8f8c} /* (5, 10, 10) {real, imag} */,
  {32'hbfd6e431, 32'hbf67ccf4} /* (5, 10, 9) {real, imag} */,
  {32'h3dfadd00, 32'h3fcc49f6} /* (5, 10, 8) {real, imag} */,
  {32'h3ec66ec4, 32'hbfc0e2c6} /* (5, 10, 7) {real, imag} */,
  {32'hc0331107, 32'h3fb61b4a} /* (5, 10, 6) {real, imag} */,
  {32'h40802761, 32'hc1034da2} /* (5, 10, 5) {real, imag} */,
  {32'h40b0d5d2, 32'hc094a086} /* (5, 10, 4) {real, imag} */,
  {32'h3fd6717f, 32'h411e66e6} /* (5, 10, 3) {real, imag} */,
  {32'h40609eb9, 32'h40ae53b4} /* (5, 10, 2) {real, imag} */,
  {32'hbf6db4b8, 32'h4187c5a4} /* (5, 10, 1) {real, imag} */,
  {32'hc131abd6, 32'hc0e58eb6} /* (5, 10, 0) {real, imag} */,
  {32'h3fd1589c, 32'hc0483d2c} /* (5, 9, 15) {real, imag} */,
  {32'h402b2b61, 32'hbff8f6dd} /* (5, 9, 14) {real, imag} */,
  {32'h400319d2, 32'hc0bd1ee4} /* (5, 9, 13) {real, imag} */,
  {32'hc0358b22, 32'h40f48222} /* (5, 9, 12) {real, imag} */,
  {32'hbf5a2250, 32'h4021e932} /* (5, 9, 11) {real, imag} */,
  {32'h3f24153c, 32'hc0541c94} /* (5, 9, 10) {real, imag} */,
  {32'h3f5d7894, 32'hbf70d1a4} /* (5, 9, 9) {real, imag} */,
  {32'hbf9d276b, 32'hc03a126e} /* (5, 9, 8) {real, imag} */,
  {32'hc017bdab, 32'hbf0ebfe4} /* (5, 9, 7) {real, imag} */,
  {32'h3fa3fe6e, 32'h3fc54cfb} /* (5, 9, 6) {real, imag} */,
  {32'hc043bbfa, 32'hbf9a0c02} /* (5, 9, 5) {real, imag} */,
  {32'h3ed359e4, 32'h401ee6b0} /* (5, 9, 4) {real, imag} */,
  {32'hbf01cd1f, 32'hbfc8e938} /* (5, 9, 3) {real, imag} */,
  {32'hc113786e, 32'h403f04d4} /* (5, 9, 2) {real, imag} */,
  {32'h411dd7fc, 32'hc0f259de} /* (5, 9, 1) {real, imag} */,
  {32'h3eef98ec, 32'h41015bfc} /* (5, 9, 0) {real, imag} */,
  {32'hbfc590c7, 32'hc135929b} /* (5, 8, 15) {real, imag} */,
  {32'h404122fd, 32'hbf8514de} /* (5, 8, 14) {real, imag} */,
  {32'h40db2676, 32'h40922cac} /* (5, 8, 13) {real, imag} */,
  {32'h40dce478, 32'h3e59b250} /* (5, 8, 12) {real, imag} */,
  {32'h4097d226, 32'hc01eae8c} /* (5, 8, 11) {real, imag} */,
  {32'hbfd554a8, 32'hbfb3d2e0} /* (5, 8, 10) {real, imag} */,
  {32'hbfd97ee4, 32'h40033b2d} /* (5, 8, 9) {real, imag} */,
  {32'h3c4e7000, 32'h3f615734} /* (5, 8, 8) {real, imag} */,
  {32'h3fe6befa, 32'hbf473b83} /* (5, 8, 7) {real, imag} */,
  {32'hbf5ea368, 32'h3d1f8f90} /* (5, 8, 6) {real, imag} */,
  {32'h3a383000, 32'hbfdb0aaf} /* (5, 8, 5) {real, imag} */,
  {32'hbfc6b82e, 32'hc01a3e8d} /* (5, 8, 4) {real, imag} */,
  {32'h4081f364, 32'h3fa440c9} /* (5, 8, 3) {real, imag} */,
  {32'hc0bb46aa, 32'hc0516767} /* (5, 8, 2) {real, imag} */,
  {32'h40619adc, 32'h40e42176} /* (5, 8, 1) {real, imag} */,
  {32'hc0b22f8f, 32'h40cd3830} /* (5, 8, 0) {real, imag} */,
  {32'hc06d3ae0, 32'hbeff1d50} /* (5, 7, 15) {real, imag} */,
  {32'hc04843a2, 32'h404376c0} /* (5, 7, 14) {real, imag} */,
  {32'h408ba5bd, 32'hc0dbb1c3} /* (5, 7, 13) {real, imag} */,
  {32'hbff7bcf2, 32'hbf3f291c} /* (5, 7, 12) {real, imag} */,
  {32'h40171630, 32'h403901c6} /* (5, 7, 11) {real, imag} */,
  {32'hbff38279, 32'h3fde0a83} /* (5, 7, 10) {real, imag} */,
  {32'hbf872e1c, 32'hbfc5aa2f} /* (5, 7, 9) {real, imag} */,
  {32'h3fe5e810, 32'h3fa9bd28} /* (5, 7, 8) {real, imag} */,
  {32'h4018f16a, 32'h3f811bb1} /* (5, 7, 7) {real, imag} */,
  {32'hc036cd10, 32'hc039630e} /* (5, 7, 6) {real, imag} */,
  {32'hbf6ee286, 32'hbf256abe} /* (5, 7, 5) {real, imag} */,
  {32'h4096b9b8, 32'hc0f70a42} /* (5, 7, 4) {real, imag} */,
  {32'h40e27b27, 32'h40194272} /* (5, 7, 3) {real, imag} */,
  {32'h404f8c46, 32'h40a610a2} /* (5, 7, 2) {real, imag} */,
  {32'hc0dcce66, 32'h41087e7c} /* (5, 7, 1) {real, imag} */,
  {32'h3f832d34, 32'h40c11ae2} /* (5, 7, 0) {real, imag} */,
  {32'hc0e5c6d4, 32'h408092ec} /* (5, 6, 15) {real, imag} */,
  {32'hc190d96e, 32'h3daff100} /* (5, 6, 14) {real, imag} */,
  {32'hc0dccd60, 32'hc09ded3c} /* (5, 6, 13) {real, imag} */,
  {32'h4017442e, 32'hc0815ba8} /* (5, 6, 12) {real, imag} */,
  {32'h3f55a444, 32'h40cb76b2} /* (5, 6, 11) {real, imag} */,
  {32'hbf83095c, 32'hc01a539d} /* (5, 6, 10) {real, imag} */,
  {32'hc010293f, 32'h3fed18fd} /* (5, 6, 9) {real, imag} */,
  {32'hbe9a40c0, 32'hc036ee7e} /* (5, 6, 8) {real, imag} */,
  {32'h3f909226, 32'h3ebd7c9c} /* (5, 6, 7) {real, imag} */,
  {32'hc099fb27, 32'h3f39236c} /* (5, 6, 6) {real, imag} */,
  {32'hc0df2864, 32'h3fd83806} /* (5, 6, 5) {real, imag} */,
  {32'h40118a72, 32'hc11f9058} /* (5, 6, 4) {real, imag} */,
  {32'h40b9820c, 32'h409239dc} /* (5, 6, 3) {real, imag} */,
  {32'hbf8bea38, 32'h3e849a30} /* (5, 6, 2) {real, imag} */,
  {32'hc1a50139, 32'h40bdaf90} /* (5, 6, 1) {real, imag} */,
  {32'h414f8b02, 32'hc09a6211} /* (5, 6, 0) {real, imag} */,
  {32'hbf98e3f8, 32'hc17b1ac7} /* (5, 5, 15) {real, imag} */,
  {32'hc014b50a, 32'h41a94ffa} /* (5, 5, 14) {real, imag} */,
  {32'hc0af7aa2, 32'h41828dc5} /* (5, 5, 13) {real, imag} */,
  {32'hc06e7502, 32'hc08947b3} /* (5, 5, 12) {real, imag} */,
  {32'h3f6c630c, 32'hc0da91de} /* (5, 5, 11) {real, imag} */,
  {32'h3fe335b6, 32'hc089d8e9} /* (5, 5, 10) {real, imag} */,
  {32'h3f5b0348, 32'hc0404028} /* (5, 5, 9) {real, imag} */,
  {32'hbae74000, 32'hc056a8c3} /* (5, 5, 8) {real, imag} */,
  {32'hc0682b7a, 32'h3f6c9220} /* (5, 5, 7) {real, imag} */,
  {32'hc0c72c8c, 32'hbff7a75c} /* (5, 5, 6) {real, imag} */,
  {32'h40dfe2ba, 32'hbf7da3e4} /* (5, 5, 5) {real, imag} */,
  {32'h410b6d64, 32'hc118b278} /* (5, 5, 4) {real, imag} */,
  {32'hc0416a54, 32'h4139b74b} /* (5, 5, 3) {real, imag} */,
  {32'hc13edc92, 32'hc0bbea82} /* (5, 5, 2) {real, imag} */,
  {32'h41b70204, 32'h40eeb99a} /* (5, 5, 1) {real, imag} */,
  {32'hc130ebf5, 32'hbf5359f4} /* (5, 5, 0) {real, imag} */,
  {32'hbf8152b8, 32'hc2041884} /* (5, 4, 15) {real, imag} */,
  {32'h3fb52060, 32'hc0cfdc08} /* (5, 4, 14) {real, imag} */,
  {32'h40c006ca, 32'hc153d98e} /* (5, 4, 13) {real, imag} */,
  {32'h3fbd4860, 32'h40f66f82} /* (5, 4, 12) {real, imag} */,
  {32'hc0d8f172, 32'hc0c71d03} /* (5, 4, 11) {real, imag} */,
  {32'h413ec9ae, 32'h402d8ba6} /* (5, 4, 10) {real, imag} */,
  {32'h3f93cb5c, 32'hc00487b4} /* (5, 4, 9) {real, imag} */,
  {32'hbf63799c, 32'h3c3bb600} /* (5, 4, 8) {real, imag} */,
  {32'h407f36ce, 32'h40c12c32} /* (5, 4, 7) {real, imag} */,
  {32'hbf9b5abc, 32'hbd8d7630} /* (5, 4, 6) {real, imag} */,
  {32'h40dbd590, 32'hbef752d0} /* (5, 4, 5) {real, imag} */,
  {32'hc1364822, 32'hbe384e10} /* (5, 4, 4) {real, imag} */,
  {32'hbfcd11c0, 32'hc12a2774} /* (5, 4, 3) {real, imag} */,
  {32'hc19f2fad, 32'h410184f0} /* (5, 4, 2) {real, imag} */,
  {32'hc1a800e6, 32'hc129de94} /* (5, 4, 1) {real, imag} */,
  {32'hc0d9bcd4, 32'h403ecd0a} /* (5, 4, 0) {real, imag} */,
  {32'h414787e5, 32'h414f63a0} /* (5, 3, 15) {real, imag} */,
  {32'h40248272, 32'hbe9d17e0} /* (5, 3, 14) {real, imag} */,
  {32'h41581a44, 32'hc0c06411} /* (5, 3, 13) {real, imag} */,
  {32'h416ec6d8, 32'h406aad09} /* (5, 3, 12) {real, imag} */,
  {32'h4188d17a, 32'h4096f100} /* (5, 3, 11) {real, imag} */,
  {32'h41483ae2, 32'hbf8ff313} /* (5, 3, 10) {real, imag} */,
  {32'hc061f723, 32'h407bfe8e} /* (5, 3, 9) {real, imag} */,
  {32'hbf0a9c54, 32'h40970d2b} /* (5, 3, 8) {real, imag} */,
  {32'hbfff931e, 32'h401c4052} /* (5, 3, 7) {real, imag} */,
  {32'h40ce635f, 32'hbe6a81d8} /* (5, 3, 6) {real, imag} */,
  {32'hc03da7e0, 32'hc1af3f2e} /* (5, 3, 5) {real, imag} */,
  {32'hc1427622, 32'h40335813} /* (5, 3, 4) {real, imag} */,
  {32'h41ac0f44, 32'h419156be} /* (5, 3, 3) {real, imag} */,
  {32'hc00fb39a, 32'h40dfcc32} /* (5, 3, 2) {real, imag} */,
  {32'hc18188a1, 32'hbfca05ec} /* (5, 3, 1) {real, imag} */,
  {32'h40bb6f0e, 32'hc11283c4} /* (5, 3, 0) {real, imag} */,
  {32'h41c3cd6c, 32'h4196d6e5} /* (5, 2, 15) {real, imag} */,
  {32'hc0ad3d0c, 32'h419fd043} /* (5, 2, 14) {real, imag} */,
  {32'hc1a9951c, 32'h40ecad2f} /* (5, 2, 13) {real, imag} */,
  {32'hc1169973, 32'hc1da9614} /* (5, 2, 12) {real, imag} */,
  {32'h40693995, 32'h41490b28} /* (5, 2, 11) {real, imag} */,
  {32'hc16aae9e, 32'h4152e8c5} /* (5, 2, 10) {real, imag} */,
  {32'h3f128350, 32'hc0ca663e} /* (5, 2, 9) {real, imag} */,
  {32'hbf8dca34, 32'hbe2f93e0} /* (5, 2, 8) {real, imag} */,
  {32'hc0d169a2, 32'h3fe9c266} /* (5, 2, 7) {real, imag} */,
  {32'h4091ea5d, 32'hc0e0ff7e} /* (5, 2, 6) {real, imag} */,
  {32'hc12b22b9, 32'h3f97005c} /* (5, 2, 5) {real, imag} */,
  {32'hc179ba15, 32'h40b99348} /* (5, 2, 4) {real, imag} */,
  {32'h41c5fb54, 32'hbfad3e0c} /* (5, 2, 3) {real, imag} */,
  {32'h4211a8a6, 32'hc184c17d} /* (5, 2, 2) {real, imag} */,
  {32'h423177de, 32'hc183895f} /* (5, 2, 1) {real, imag} */,
  {32'h40ab4d79, 32'hc02bf8c6} /* (5, 2, 0) {real, imag} */,
  {32'h41dddb7e, 32'h4119d044} /* (5, 1, 15) {real, imag} */,
  {32'hc23c1972, 32'hc1d157d8} /* (5, 1, 14) {real, imag} */,
  {32'h413abc9f, 32'h411bb53c} /* (5, 1, 13) {real, imag} */,
  {32'h4101feac, 32'h41ad2abc} /* (5, 1, 12) {real, imag} */,
  {32'hc09b05b8, 32'h40c34d1c} /* (5, 1, 11) {real, imag} */,
  {32'hbfd31a50, 32'hc0fd1202} /* (5, 1, 10) {real, imag} */,
  {32'hc10e6b52, 32'h40f1ef93} /* (5, 1, 9) {real, imag} */,
  {32'hc02320c2, 32'h3fd95e00} /* (5, 1, 8) {real, imag} */,
  {32'h3fdbe650, 32'h3cc6e300} /* (5, 1, 7) {real, imag} */,
  {32'h411f0e22, 32'h40cc2306} /* (5, 1, 6) {real, imag} */,
  {32'hc041b11d, 32'hc1be1ccf} /* (5, 1, 5) {real, imag} */,
  {32'h40a0ef96, 32'hc0928e32} /* (5, 1, 4) {real, imag} */,
  {32'hc0bc54b2, 32'hc204a280} /* (5, 1, 3) {real, imag} */,
  {32'h4136bffc, 32'h41fd01b6} /* (5, 1, 2) {real, imag} */,
  {32'h414ae5b4, 32'hc113435e} /* (5, 1, 1) {real, imag} */,
  {32'h4189bcc7, 32'h41e41ccc} /* (5, 1, 0) {real, imag} */,
  {32'hc1551ea2, 32'h4190ae64} /* (5, 0, 15) {real, imag} */,
  {32'hc18347f2, 32'h40f4c7b5} /* (5, 0, 14) {real, imag} */,
  {32'hc11800b6, 32'h410a337d} /* (5, 0, 13) {real, imag} */,
  {32'h41592801, 32'hc0ac52ec} /* (5, 0, 12) {real, imag} */,
  {32'hc03bc31a, 32'hc1eed974} /* (5, 0, 11) {real, imag} */,
  {32'hbf9590e0, 32'hc0f235e6} /* (5, 0, 10) {real, imag} */,
  {32'h407a0841, 32'hc1063a8f} /* (5, 0, 9) {real, imag} */,
  {32'hc02470b4, 32'hbd8bc300} /* (5, 0, 8) {real, imag} */,
  {32'hc0dc02e0, 32'hc0147b0c} /* (5, 0, 7) {real, imag} */,
  {32'h40c90ec8, 32'hc0f4778a} /* (5, 0, 6) {real, imag} */,
  {32'hc0d37655, 32'h412707a8} /* (5, 0, 5) {real, imag} */,
  {32'h410a1875, 32'hc1dc13c9} /* (5, 0, 4) {real, imag} */,
  {32'hc127fd62, 32'hc133bdd9} /* (5, 0, 3) {real, imag} */,
  {32'hc1928d1e, 32'h3dcd46c0} /* (5, 0, 2) {real, imag} */,
  {32'h40f9db14, 32'hc0551a44} /* (5, 0, 1) {real, imag} */,
  {32'h41eb0f90, 32'hc21d4f90} /* (5, 0, 0) {real, imag} */,
  {32'h402435b0, 32'h41366f82} /* (4, 15, 15) {real, imag} */,
  {32'h4191510c, 32'hc0d857b4} /* (4, 15, 14) {real, imag} */,
  {32'hbf89ffe8, 32'h3f9e476e} /* (4, 15, 13) {real, imag} */,
  {32'h41b88401, 32'hc19ac937} /* (4, 15, 12) {real, imag} */,
  {32'hc130331a, 32'hc0328468} /* (4, 15, 11) {real, imag} */,
  {32'h3fd2b5c4, 32'hc15af9bb} /* (4, 15, 10) {real, imag} */,
  {32'hc05a5d8e, 32'h40d2adad} /* (4, 15, 9) {real, imag} */,
  {32'hc0dff8e8, 32'h4100d31e} /* (4, 15, 8) {real, imag} */,
  {32'h413a6e82, 32'hbf1bead8} /* (4, 15, 7) {real, imag} */,
  {32'hc0afe29b, 32'hc0a19bca} /* (4, 15, 6) {real, imag} */,
  {32'hc19a0091, 32'hc13040b4} /* (4, 15, 5) {real, imag} */,
  {32'h3f8d3d50, 32'h40d006f4} /* (4, 15, 4) {real, imag} */,
  {32'hc191d61a, 32'hc0841248} /* (4, 15, 3) {real, imag} */,
  {32'hc22bf616, 32'hc03e64ed} /* (4, 15, 2) {real, imag} */,
  {32'h42086af1, 32'hc20ca0f6} /* (4, 15, 1) {real, imag} */,
  {32'h4299f14a, 32'h4237507c} /* (4, 15, 0) {real, imag} */,
  {32'h420dfc9d, 32'hc117957e} /* (4, 14, 15) {real, imag} */,
  {32'h41ddca80, 32'h419f5f7a} /* (4, 14, 14) {real, imag} */,
  {32'hc10c686d, 32'h41adb1f6} /* (4, 14, 13) {real, imag} */,
  {32'h4031bc7c, 32'hbe2998c0} /* (4, 14, 12) {real, imag} */,
  {32'hc155fb6d, 32'h416b38ff} /* (4, 14, 11) {real, imag} */,
  {32'h41457fdc, 32'h414882bb} /* (4, 14, 10) {real, imag} */,
  {32'hc089e82e, 32'hc12e19ae} /* (4, 14, 9) {real, imag} */,
  {32'hc09423a4, 32'hc1009b9c} /* (4, 14, 8) {real, imag} */,
  {32'hc154c38b, 32'h40232086} /* (4, 14, 7) {real, imag} */,
  {32'h40272f42, 32'hc1773f09} /* (4, 14, 6) {real, imag} */,
  {32'hc0e5385e, 32'h4162efe9} /* (4, 14, 5) {real, imag} */,
  {32'hbf1b39b0, 32'hc1bd5e46} /* (4, 14, 4) {real, imag} */,
  {32'hc117629f, 32'h40857f76} /* (4, 14, 3) {real, imag} */,
  {32'h42108e05, 32'h40ac813e} /* (4, 14, 2) {real, imag} */,
  {32'hc250856f, 32'hc1a538eb} /* (4, 14, 1) {real, imag} */,
  {32'hc1a28221, 32'hc25d2115} /* (4, 14, 0) {real, imag} */,
  {32'hc1868880, 32'h3e97dc50} /* (4, 13, 15) {real, imag} */,
  {32'hc13d4489, 32'h41c52ba6} /* (4, 13, 14) {real, imag} */,
  {32'hc1260a4e, 32'hc15bdbf6} /* (4, 13, 13) {real, imag} */,
  {32'hc165af11, 32'h40cc8e33} /* (4, 13, 12) {real, imag} */,
  {32'hc10990fb, 32'h40cbe56e} /* (4, 13, 11) {real, imag} */,
  {32'h4188bbb3, 32'hc115d508} /* (4, 13, 10) {real, imag} */,
  {32'hc10cfc66, 32'h4169794c} /* (4, 13, 9) {real, imag} */,
  {32'hc1019c76, 32'hbf6b1e38} /* (4, 13, 8) {real, imag} */,
  {32'hbfdd2d3c, 32'h4120e050} /* (4, 13, 7) {real, imag} */,
  {32'hc090aa31, 32'h40e26337} /* (4, 13, 6) {real, imag} */,
  {32'h40faa19e, 32'hc1b576e2} /* (4, 13, 5) {real, imag} */,
  {32'h410a888b, 32'hbf8c14c4} /* (4, 13, 4) {real, imag} */,
  {32'hbfa3c100, 32'h40ce10bc} /* (4, 13, 3) {real, imag} */,
  {32'h4139aefd, 32'h4102fabc} /* (4, 13, 2) {real, imag} */,
  {32'hc181ad80, 32'hc15cd614} /* (4, 13, 1) {real, imag} */,
  {32'h41296134, 32'h408689a1} /* (4, 13, 0) {real, imag} */,
  {32'hbfbe40c0, 32'hc066cea0} /* (4, 12, 15) {real, imag} */,
  {32'hc0ebe2fa, 32'hc1bd6ce6} /* (4, 12, 14) {real, imag} */,
  {32'h40af7e5c, 32'hc023655e} /* (4, 12, 13) {real, imag} */,
  {32'hc207d26d, 32'h3ea2df60} /* (4, 12, 12) {real, imag} */,
  {32'h40b3539b, 32'hbff337f4} /* (4, 12, 11) {real, imag} */,
  {32'hbeb15f60, 32'hbfc646a2} /* (4, 12, 10) {real, imag} */,
  {32'h40bbb21a, 32'h40e480d2} /* (4, 12, 9) {real, imag} */,
  {32'h40d645d0, 32'h3ffbcee0} /* (4, 12, 8) {real, imag} */,
  {32'hbf5dca50, 32'hc0bc709a} /* (4, 12, 7) {real, imag} */,
  {32'h415a65c3, 32'h40f262e0} /* (4, 12, 6) {real, imag} */,
  {32'h40df55c3, 32'h40d59dad} /* (4, 12, 5) {real, imag} */,
  {32'h3f8230e0, 32'h40a13e1e} /* (4, 12, 4) {real, imag} */,
  {32'h410db9b5, 32'h4159a24c} /* (4, 12, 3) {real, imag} */,
  {32'hc1cbb65c, 32'h4163b66c} /* (4, 12, 2) {real, imag} */,
  {32'h418f4d03, 32'h4199d605} /* (4, 12, 1) {real, imag} */,
  {32'hc0b12778, 32'h415d507a} /* (4, 12, 0) {real, imag} */,
  {32'hc21adf51, 32'hc1b8d409} /* (4, 11, 15) {real, imag} */,
  {32'hbfa6ad60, 32'hc195a684} /* (4, 11, 14) {real, imag} */,
  {32'hc187c666, 32'h40f1c08e} /* (4, 11, 13) {real, imag} */,
  {32'h41135861, 32'h4152c53f} /* (4, 11, 12) {real, imag} */,
  {32'h3f8984bc, 32'hc0d82fe0} /* (4, 11, 11) {real, imag} */,
  {32'h3f708100, 32'h40631f32} /* (4, 11, 10) {real, imag} */,
  {32'hc0bd6b36, 32'hbed1c760} /* (4, 11, 9) {real, imag} */,
  {32'h3f4b7d20, 32'h40877a1c} /* (4, 11, 8) {real, imag} */,
  {32'hbfaac7c8, 32'h3f2fc8a0} /* (4, 11, 7) {real, imag} */,
  {32'hc0f56b64, 32'hc01dd72a} /* (4, 11, 6) {real, imag} */,
  {32'h401fa6da, 32'h406c01b1} /* (4, 11, 5) {real, imag} */,
  {32'h41031999, 32'hc0b8dba6} /* (4, 11, 4) {real, imag} */,
  {32'h401211ec, 32'hbfd6c916} /* (4, 11, 3) {real, imag} */,
  {32'h4101c12a, 32'h4145ba64} /* (4, 11, 2) {real, imag} */,
  {32'hc19aa46c, 32'hbbeff000} /* (4, 11, 1) {real, imag} */,
  {32'hc1849d7e, 32'h41aef3c7} /* (4, 11, 0) {real, imag} */,
  {32'hc1dcee71, 32'h3fed5828} /* (4, 10, 15) {real, imag} */,
  {32'h41db0ea8, 32'hc0a55250} /* (4, 10, 14) {real, imag} */,
  {32'h40c3ee54, 32'hbe9d6680} /* (4, 10, 13) {real, imag} */,
  {32'hc0bef522, 32'h40b413de} /* (4, 10, 12) {real, imag} */,
  {32'hc0766818, 32'h4055ba6a} /* (4, 10, 11) {real, imag} */,
  {32'hc1049fd5, 32'hbfdecca4} /* (4, 10, 10) {real, imag} */,
  {32'h3f375960, 32'h3fa2fbcb} /* (4, 10, 9) {real, imag} */,
  {32'hbf5c4020, 32'hc01aa6f5} /* (4, 10, 8) {real, imag} */,
  {32'hbf99be10, 32'h3f54d212} /* (4, 10, 7) {real, imag} */,
  {32'hc077008c, 32'h3fab8924} /* (4, 10, 6) {real, imag} */,
  {32'h4122071a, 32'hc0dae88d} /* (4, 10, 5) {real, imag} */,
  {32'h4056e09c, 32'hc1006690} /* (4, 10, 4) {real, imag} */,
  {32'h4144beb6, 32'h3fcf2068} /* (4, 10, 3) {real, imag} */,
  {32'h40a3e09e, 32'h41afe2b8} /* (4, 10, 2) {real, imag} */,
  {32'h411f5a2a, 32'h4105ff69} /* (4, 10, 1) {real, imag} */,
  {32'hc095c902, 32'hc0c2239a} /* (4, 10, 0) {real, imag} */,
  {32'h40d1347b, 32'hc01be7eb} /* (4, 9, 15) {real, imag} */,
  {32'hc0665015, 32'h40cc807c} /* (4, 9, 14) {real, imag} */,
  {32'hc0d406a6, 32'hbf631f1c} /* (4, 9, 13) {real, imag} */,
  {32'h4067b209, 32'h4017f620} /* (4, 9, 12) {real, imag} */,
  {32'h4084cfe6, 32'hbfda7c6c} /* (4, 9, 11) {real, imag} */,
  {32'hbfa0a110, 32'h409b1fac} /* (4, 9, 10) {real, imag} */,
  {32'hbe6f3b60, 32'hbcdf71a0} /* (4, 9, 9) {real, imag} */,
  {32'h3f2f7b9a, 32'h400718c4} /* (4, 9, 8) {real, imag} */,
  {32'hbf5b0778, 32'h3f134e53} /* (4, 9, 7) {real, imag} */,
  {32'h4025609d, 32'hc0c7b2a8} /* (4, 9, 6) {real, imag} */,
  {32'hbfc87eab, 32'h4031c64c} /* (4, 9, 5) {real, imag} */,
  {32'hc028de13, 32'hbd7616a0} /* (4, 9, 4) {real, imag} */,
  {32'hbefb29a8, 32'hc07501eb} /* (4, 9, 3) {real, imag} */,
  {32'h40c291ce, 32'hc0a25fd4} /* (4, 9, 2) {real, imag} */,
  {32'hc1acb8c7, 32'h40cdaad2} /* (4, 9, 1) {real, imag} */,
  {32'h3d301e60, 32'hc048661c} /* (4, 9, 0) {real, imag} */,
  {32'h41687344, 32'h3eb1e451} /* (4, 8, 15) {real, imag} */,
  {32'hc0a2a1b2, 32'h3edddb20} /* (4, 8, 14) {real, imag} */,
  {32'hbfacc64f, 32'hc00a8810} /* (4, 8, 13) {real, imag} */,
  {32'hc09642bc, 32'h410e15b5} /* (4, 8, 12) {real, imag} */,
  {32'hbfcb4e93, 32'h404e3c88} /* (4, 8, 11) {real, imag} */,
  {32'h40dfced6, 32'h405f857e} /* (4, 8, 10) {real, imag} */,
  {32'h3ea4f3ec, 32'hbfc0f9e4} /* (4, 8, 9) {real, imag} */,
  {32'hbfdb6720, 32'h3f9fb3fa} /* (4, 8, 8) {real, imag} */,
  {32'hbed097ac, 32'h3e29c3b4} /* (4, 8, 7) {real, imag} */,
  {32'h409ed5ee, 32'h403e18b2} /* (4, 8, 6) {real, imag} */,
  {32'hc0ade486, 32'hc09ba7f0} /* (4, 8, 5) {real, imag} */,
  {32'h4060d6f8, 32'hbfa0cc58} /* (4, 8, 4) {real, imag} */,
  {32'hbfc3da1d, 32'h40980a1f} /* (4, 8, 3) {real, imag} */,
  {32'h40c5a042, 32'hc0d1c4a8} /* (4, 8, 2) {real, imag} */,
  {32'h40f349ab, 32'hbfa95f0d} /* (4, 8, 1) {real, imag} */,
  {32'hc152d034, 32'h4012db7b} /* (4, 8, 0) {real, imag} */,
  {32'hbf49617c, 32'h414fbfa8} /* (4, 7, 15) {real, imag} */,
  {32'hc100d872, 32'h40c46320} /* (4, 7, 14) {real, imag} */,
  {32'h4093edea, 32'hbfa79ca8} /* (4, 7, 13) {real, imag} */,
  {32'hc176e5ac, 32'hbe3c3bc0} /* (4, 7, 12) {real, imag} */,
  {32'hbf6561cc, 32'h3f693092} /* (4, 7, 11) {real, imag} */,
  {32'h3eba7050, 32'hc06f0ceb} /* (4, 7, 10) {real, imag} */,
  {32'h4070cfb5, 32'h3fcefcf6} /* (4, 7, 9) {real, imag} */,
  {32'h3f808cd9, 32'h3ebb8bc0} /* (4, 7, 8) {real, imag} */,
  {32'hbf3f1eec, 32'h4006ea6b} /* (4, 7, 7) {real, imag} */,
  {32'hc0da16db, 32'h40240535} /* (4, 7, 6) {real, imag} */,
  {32'h40a05c26, 32'hc031b0d8} /* (4, 7, 5) {real, imag} */,
  {32'hbf82423c, 32'h409b0844} /* (4, 7, 4) {real, imag} */,
  {32'hc03a15df, 32'h40b0ee18} /* (4, 7, 3) {real, imag} */,
  {32'h4118b0f2, 32'h402b2af0} /* (4, 7, 2) {real, imag} */,
  {32'h405a7f5d, 32'hc13dcec0} /* (4, 7, 1) {real, imag} */,
  {32'h406142e8, 32'hc187b073} /* (4, 7, 0) {real, imag} */,
  {32'hc0203b4b, 32'h41f7a788} /* (4, 6, 15) {real, imag} */,
  {32'hbf9d0f50, 32'hc1167734} /* (4, 6, 14) {real, imag} */,
  {32'hbf622e24, 32'h3f9cf2e4} /* (4, 6, 13) {real, imag} */,
  {32'hc161b15c, 32'hc088421e} /* (4, 6, 12) {real, imag} */,
  {32'hc006c46f, 32'hbfeae598} /* (4, 6, 11) {real, imag} */,
  {32'h4003e7c2, 32'h3eda9418} /* (4, 6, 10) {real, imag} */,
  {32'hc0258bda, 32'hc0ac5fd6} /* (4, 6, 9) {real, imag} */,
  {32'h40805e0d, 32'h401f213c} /* (4, 6, 8) {real, imag} */,
  {32'hbf7dc595, 32'hbcd94e00} /* (4, 6, 7) {real, imag} */,
  {32'h408c6557, 32'h3ffd5712} /* (4, 6, 6) {real, imag} */,
  {32'hc069075d, 32'h40a08110} /* (4, 6, 5) {real, imag} */,
  {32'h41383e3a, 32'h41986434} /* (4, 6, 4) {real, imag} */,
  {32'hc0f6660a, 32'hc174bd40} /* (4, 6, 3) {real, imag} */,
  {32'h419376df, 32'hc0dc7408} /* (4, 6, 2) {real, imag} */,
  {32'hbfdbf282, 32'hc19d92ae} /* (4, 6, 1) {real, imag} */,
  {32'hc14a99aa, 32'h41ed5bc4} /* (4, 6, 0) {real, imag} */,
  {32'hc21df71e, 32'h412677f6} /* (4, 5, 15) {real, imag} */,
  {32'hc0af2901, 32'hc176c5a2} /* (4, 5, 14) {real, imag} */,
  {32'hc0ac9f7c, 32'hc15f4efe} /* (4, 5, 13) {real, imag} */,
  {32'h40a7a624, 32'hc12c5426} /* (4, 5, 12) {real, imag} */,
  {32'hc16e1816, 32'h3ff3847c} /* (4, 5, 11) {real, imag} */,
  {32'hc04a961e, 32'hc112a584} /* (4, 5, 10) {real, imag} */,
  {32'h4097d764, 32'hbfaa595c} /* (4, 5, 9) {real, imag} */,
  {32'h403ded21, 32'h404fb243} /* (4, 5, 8) {real, imag} */,
  {32'h409fb444, 32'h3fc7ac1c} /* (4, 5, 7) {real, imag} */,
  {32'h402785e2, 32'h40240b18} /* (4, 5, 6) {real, imag} */,
  {32'h4111bfaa, 32'hc1215d8c} /* (4, 5, 5) {real, imag} */,
  {32'h409fb588, 32'h41243476} /* (4, 5, 4) {real, imag} */,
  {32'hc1e79d0f, 32'h41f618d7} /* (4, 5, 3) {real, imag} */,
  {32'hbe899a10, 32'hc150ddd8} /* (4, 5, 2) {real, imag} */,
  {32'h3f53e0a0, 32'h41695ef2} /* (4, 5, 1) {real, imag} */,
  {32'hbe2cd4b0, 32'h409ab82a} /* (4, 5, 0) {real, imag} */,
  {32'h41fd8e96, 32'hc1346126} /* (4, 4, 15) {real, imag} */,
  {32'h4119b924, 32'h415565cd} /* (4, 4, 14) {real, imag} */,
  {32'hc0db8d6a, 32'h41bea416} /* (4, 4, 13) {real, imag} */,
  {32'h410f4a92, 32'h410be3c6} /* (4, 4, 12) {real, imag} */,
  {32'h3fe41490, 32'h4109448a} /* (4, 4, 11) {real, imag} */,
  {32'hc1a73206, 32'hc0d18cff} /* (4, 4, 10) {real, imag} */,
  {32'hbe2f31d0, 32'h413a1a29} /* (4, 4, 9) {real, imag} */,
  {32'h4082e7fa, 32'hbca01780} /* (4, 4, 8) {real, imag} */,
  {32'h40793a5d, 32'hc033ba14} /* (4, 4, 7) {real, imag} */,
  {32'h404e5870, 32'hc1068e82} /* (4, 4, 6) {real, imag} */,
  {32'h41466f7a, 32'h3f4b3198} /* (4, 4, 5) {real, imag} */,
  {32'h41058a12, 32'h3fab3634} /* (4, 4, 4) {real, imag} */,
  {32'hc15ba2e7, 32'hc11e7bc4} /* (4, 4, 3) {real, imag} */,
  {32'hc0cf3b80, 32'h413a2e81} /* (4, 4, 2) {real, imag} */,
  {32'h414c27e4, 32'h40e57e80} /* (4, 4, 1) {real, imag} */,
  {32'h417031f7, 32'h40c9df82} /* (4, 4, 0) {real, imag} */,
  {32'hc1ba88b6, 32'h40fcddde} /* (4, 3, 15) {real, imag} */,
  {32'h408955cd, 32'hc0c06aec} /* (4, 3, 14) {real, imag} */,
  {32'hc16bce66, 32'hc178552f} /* (4, 3, 13) {real, imag} */,
  {32'hc0fcd7de, 32'hc126358a} /* (4, 3, 12) {real, imag} */,
  {32'h4126afa1, 32'h40f1061e} /* (4, 3, 11) {real, imag} */,
  {32'h4150e01c, 32'hc14c6744} /* (4, 3, 10) {real, imag} */,
  {32'h40de76d9, 32'h3fd6966e} /* (4, 3, 9) {real, imag} */,
  {32'h409ed4da, 32'hbf656e5e} /* (4, 3, 8) {real, imag} */,
  {32'hc05b4e06, 32'h4107fd96} /* (4, 3, 7) {real, imag} */,
  {32'h4146ef64, 32'h3feb9318} /* (4, 3, 6) {real, imag} */,
  {32'h41a2cca4, 32'h4181baa4} /* (4, 3, 5) {real, imag} */,
  {32'hc1d9bd4a, 32'h41069c84} /* (4, 3, 4) {real, imag} */,
  {32'hbf151bb8, 32'hc148bead} /* (4, 3, 3) {real, imag} */,
  {32'h412dda02, 32'h4124d9da} /* (4, 3, 2) {real, imag} */,
  {32'hc0e9873a, 32'h41b5b49e} /* (4, 3, 1) {real, imag} */,
  {32'h4154f2e7, 32'h409c0e30} /* (4, 3, 0) {real, imag} */,
  {32'h418e56e6, 32'h41d9f9db} /* (4, 2, 15) {real, imag} */,
  {32'hc0f50116, 32'hc2018560} /* (4, 2, 14) {real, imag} */,
  {32'h4212f34c, 32'h41826fd6} /* (4, 2, 13) {real, imag} */,
  {32'h408ee514, 32'h413bd327} /* (4, 2, 12) {real, imag} */,
  {32'h4156fbd8, 32'h40dbe7d4} /* (4, 2, 11) {real, imag} */,
  {32'hbf5e03f0, 32'hc06e7778} /* (4, 2, 10) {real, imag} */,
  {32'hbfcace2a, 32'h4013b87f} /* (4, 2, 9) {real, imag} */,
  {32'h415e0960, 32'h4032c804} /* (4, 2, 8) {real, imag} */,
  {32'hc1031bf9, 32'hc030a9bf} /* (4, 2, 7) {real, imag} */,
  {32'h41795ce9, 32'h414bb7da} /* (4, 2, 6) {real, imag} */,
  {32'hc03671c0, 32'hc108d5e8} /* (4, 2, 5) {real, imag} */,
  {32'hc02f1524, 32'hc1bdf84c} /* (4, 2, 4) {real, imag} */,
  {32'h418facfb, 32'hc17b8a63} /* (4, 2, 3) {real, imag} */,
  {32'h413eec6d, 32'hc13d5404} /* (4, 2, 2) {real, imag} */,
  {32'h4119512f, 32'h413699f6} /* (4, 2, 1) {real, imag} */,
  {32'hc214d998, 32'hc1bccf78} /* (4, 2, 0) {real, imag} */,
  {32'h3ef49900, 32'h425ab231} /* (4, 1, 15) {real, imag} */,
  {32'hc1cff37a, 32'h4088bfe0} /* (4, 1, 14) {real, imag} */,
  {32'hc18155ca, 32'hc2168976} /* (4, 1, 13) {real, imag} */,
  {32'h40b348c2, 32'hc1b09574} /* (4, 1, 12) {real, imag} */,
  {32'hc120ca24, 32'hbf1508f8} /* (4, 1, 11) {real, imag} */,
  {32'h41062ca7, 32'h4191f4e9} /* (4, 1, 10) {real, imag} */,
  {32'h4042f6a8, 32'hbf96f948} /* (4, 1, 9) {real, imag} */,
  {32'hc1016918, 32'h404b7d36} /* (4, 1, 8) {real, imag} */,
  {32'hbff46470, 32'h3ff594a8} /* (4, 1, 7) {real, imag} */,
  {32'hc0c966b2, 32'hbecc8ec0} /* (4, 1, 6) {real, imag} */,
  {32'hc1533dd2, 32'h4136e54c} /* (4, 1, 5) {real, imag} */,
  {32'h41135992, 32'h3fe8efc8} /* (4, 1, 4) {real, imag} */,
  {32'hc11097f6, 32'h41ef5f24} /* (4, 1, 3) {real, imag} */,
  {32'h41f966ae, 32'h3f5ed1d4} /* (4, 1, 2) {real, imag} */,
  {32'hc1c87d5b, 32'h419262fe} /* (4, 1, 1) {real, imag} */,
  {32'hc14a15dc, 32'hc0ed6e25} /* (4, 1, 0) {real, imag} */,
  {32'hc23344c8, 32'hc13b10c7} /* (4, 0, 15) {real, imag} */,
  {32'hc207aa2c, 32'hc106e6ea} /* (4, 0, 14) {real, imag} */,
  {32'h41d0a76a, 32'h421a2840} /* (4, 0, 13) {real, imag} */,
  {32'h4144b7cc, 32'h4113c7a4} /* (4, 0, 12) {real, imag} */,
  {32'h415df689, 32'hc1a1b00a} /* (4, 0, 11) {real, imag} */,
  {32'hc0ab4d57, 32'hbfc739af} /* (4, 0, 10) {real, imag} */,
  {32'h412c7012, 32'hc0808c5c} /* (4, 0, 9) {real, imag} */,
  {32'hbf8e5470, 32'hbf9913ec} /* (4, 0, 8) {real, imag} */,
  {32'hc02de12e, 32'hc0f1aba8} /* (4, 0, 7) {real, imag} */,
  {32'hc1087b82, 32'hbf813251} /* (4, 0, 6) {real, imag} */,
  {32'hc03b14ec, 32'h41ddfb76} /* (4, 0, 5) {real, imag} */,
  {32'hc1a8eb9e, 32'hc1d4805c} /* (4, 0, 4) {real, imag} */,
  {32'h406fd114, 32'hc19c9117} /* (4, 0, 3) {real, imag} */,
  {32'hc103774a, 32'hbfb57334} /* (4, 0, 2) {real, imag} */,
  {32'h3f1ef1e0, 32'hc20e657a} /* (4, 0, 1) {real, imag} */,
  {32'hc199457d, 32'h4028cad2} /* (4, 0, 0) {real, imag} */,
  {32'h40971120, 32'h40205c84} /* (3, 15, 15) {real, imag} */,
  {32'hc256087a, 32'hc1b1094f} /* (3, 15, 14) {real, imag} */,
  {32'h418d1aca, 32'h41a8beba} /* (3, 15, 13) {real, imag} */,
  {32'h4049a2e8, 32'h421ab26c} /* (3, 15, 12) {real, imag} */,
  {32'h418d3566, 32'h42112acc} /* (3, 15, 11) {real, imag} */,
  {32'h41bf301c, 32'h41733f78} /* (3, 15, 10) {real, imag} */,
  {32'h40019c78, 32'hc0b75862} /* (3, 15, 9) {real, imag} */,
  {32'hc0dc9fde, 32'h408c449a} /* (3, 15, 8) {real, imag} */,
  {32'hc0f4cc7c, 32'h40c87662} /* (3, 15, 7) {real, imag} */,
  {32'hc0bbc39e, 32'h419347da} /* (3, 15, 6) {real, imag} */,
  {32'h418e661e, 32'hc2271c3c} /* (3, 15, 5) {real, imag} */,
  {32'h41ab36b4, 32'h3e1be080} /* (3, 15, 4) {real, imag} */,
  {32'hc18b243a, 32'hc1cbc81c} /* (3, 15, 3) {real, imag} */,
  {32'hc0f80fa0, 32'h41993429} /* (3, 15, 2) {real, imag} */,
  {32'hc2516937, 32'hc1c49824} /* (3, 15, 1) {real, imag} */,
  {32'h4174f80d, 32'hc1159489} /* (3, 15, 0) {real, imag} */,
  {32'h413a0966, 32'hc1f00d38} /* (3, 14, 15) {real, imag} */,
  {32'hc1e6d8d7, 32'hc146c688} /* (3, 14, 14) {real, imag} */,
  {32'h4078a271, 32'hc208744a} /* (3, 14, 13) {real, imag} */,
  {32'hbda93080, 32'h41ab1f01} /* (3, 14, 12) {real, imag} */,
  {32'h4007522a, 32'hc0de3613} /* (3, 14, 11) {real, imag} */,
  {32'hc0e725e4, 32'hbf1b4a5c} /* (3, 14, 10) {real, imag} */,
  {32'h3dc74d40, 32'h40843d5d} /* (3, 14, 9) {real, imag} */,
  {32'hc0bffb26, 32'hc121c2c6} /* (3, 14, 8) {real, imag} */,
  {32'hc1649062, 32'hc14ed2fc} /* (3, 14, 7) {real, imag} */,
  {32'hc1d2a11b, 32'h40a78c50} /* (3, 14, 6) {real, imag} */,
  {32'h415ead48, 32'h40a1687d} /* (3, 14, 5) {real, imag} */,
  {32'h4177d1db, 32'h3f9175b0} /* (3, 14, 4) {real, imag} */,
  {32'h3f31ded4, 32'h41820feb} /* (3, 14, 3) {real, imag} */,
  {32'hc171fc4a, 32'hbff66d70} /* (3, 14, 2) {real, imag} */,
  {32'hc137aff6, 32'hc012888c} /* (3, 14, 1) {real, imag} */,
  {32'h41d121bc, 32'h40eefca3} /* (3, 14, 0) {real, imag} */,
  {32'hc18edeb4, 32'h417d9994} /* (3, 13, 15) {real, imag} */,
  {32'hc166ca74, 32'hc1cec1bc} /* (3, 13, 14) {real, imag} */,
  {32'h41fa49ee, 32'h41922899} /* (3, 13, 13) {real, imag} */,
  {32'h4245901d, 32'hc189a1cd} /* (3, 13, 12) {real, imag} */,
  {32'hc13d209f, 32'hc13c4152} /* (3, 13, 11) {real, imag} */,
  {32'h40676840, 32'h4093a12f} /* (3, 13, 10) {real, imag} */,
  {32'h40a5e9a5, 32'h4094dc16} /* (3, 13, 9) {real, imag} */,
  {32'h41882aaa, 32'hbfadc4f0} /* (3, 13, 8) {real, imag} */,
  {32'h40635bea, 32'hc0213b78} /* (3, 13, 7) {real, imag} */,
  {32'h419ae224, 32'h413ebee6} /* (3, 13, 6) {real, imag} */,
  {32'h41602739, 32'h40c3c8fd} /* (3, 13, 5) {real, imag} */,
  {32'hbf0e65c0, 32'h40e9e79c} /* (3, 13, 4) {real, imag} */,
  {32'h40db6f58, 32'hc1d89311} /* (3, 13, 3) {real, imag} */,
  {32'hc1f4c3fa, 32'hc107d570} /* (3, 13, 2) {real, imag} */,
  {32'h41adeb40, 32'hc09ef271} /* (3, 13, 1) {real, imag} */,
  {32'hc1d595ba, 32'h3f1c4fa0} /* (3, 13, 0) {real, imag} */,
  {32'h41be7e51, 32'h40579128} /* (3, 12, 15) {real, imag} */,
  {32'hbffcd8b0, 32'h412aff49} /* (3, 12, 14) {real, imag} */,
  {32'h41948262, 32'hc173b858} /* (3, 12, 13) {real, imag} */,
  {32'hbf7e85e0, 32'h4040590a} /* (3, 12, 12) {real, imag} */,
  {32'hc171db8d, 32'hc1a9ad12} /* (3, 12, 11) {real, imag} */,
  {32'hc145143c, 32'h40a9e184} /* (3, 12, 10) {real, imag} */,
  {32'h414b44b4, 32'hc022e958} /* (3, 12, 9) {real, imag} */,
  {32'hbf36fb74, 32'hc0e1920c} /* (3, 12, 8) {real, imag} */,
  {32'hbfddf0c4, 32'h3f992b50} /* (3, 12, 7) {real, imag} */,
  {32'hc18e0f82, 32'h4138ce88} /* (3, 12, 6) {real, imag} */,
  {32'h3e5821c0, 32'h414d4dd1} /* (3, 12, 5) {real, imag} */,
  {32'hc1d97a1e, 32'hbf06ee22} /* (3, 12, 4) {real, imag} */,
  {32'h41f5bbfe, 32'h4087eca8} /* (3, 12, 3) {real, imag} */,
  {32'h410c05c9, 32'h407ead0b} /* (3, 12, 2) {real, imag} */,
  {32'h41059c66, 32'hc24b1372} /* (3, 12, 1) {real, imag} */,
  {32'hc0e3d25e, 32'h408ea9e8} /* (3, 12, 0) {real, imag} */,
  {32'hc184391a, 32'h419fa936} /* (3, 11, 15) {real, imag} */,
  {32'h420706c8, 32'h4116bea8} /* (3, 11, 14) {real, imag} */,
  {32'hbf7fa840, 32'h3f962dc0} /* (3, 11, 13) {real, imag} */,
  {32'hc15ce405, 32'hc12a1d66} /* (3, 11, 12) {real, imag} */,
  {32'hc04a2b7a, 32'h40cf09d1} /* (3, 11, 11) {real, imag} */,
  {32'h3f2c3170, 32'hc121e0d0} /* (3, 11, 10) {real, imag} */,
  {32'hc10cff71, 32'h40ca0090} /* (3, 11, 9) {real, imag} */,
  {32'h3e0837a0, 32'hbfb3b6a4} /* (3, 11, 8) {real, imag} */,
  {32'h40ddce8e, 32'hc0b1e9e4} /* (3, 11, 7) {real, imag} */,
  {32'h412355ee, 32'hc0afc334} /* (3, 11, 6) {real, imag} */,
  {32'h40732492, 32'hc166fa74} /* (3, 11, 5) {real, imag} */,
  {32'hc11331cb, 32'hbf093978} /* (3, 11, 4) {real, imag} */,
  {32'hc18b47b4, 32'hc0a48342} /* (3, 11, 3) {real, imag} */,
  {32'h3e7aef00, 32'h4150a40a} /* (3, 11, 2) {real, imag} */,
  {32'h41efd3ca, 32'h41cd2ef6} /* (3, 11, 1) {real, imag} */,
  {32'hc17c084e, 32'h401a36a8} /* (3, 11, 0) {real, imag} */,
  {32'hc10c1cd8, 32'hc11d31f6} /* (3, 10, 15) {real, imag} */,
  {32'h3f1578d8, 32'hc1271254} /* (3, 10, 14) {real, imag} */,
  {32'hc06be550, 32'h41a72fb8} /* (3, 10, 13) {real, imag} */,
  {32'hc1274dea, 32'hc0d6c104} /* (3, 10, 12) {real, imag} */,
  {32'hc0448214, 32'h40b8d3a8} /* (3, 10, 11) {real, imag} */,
  {32'hc07878ca, 32'hc10529b1} /* (3, 10, 10) {real, imag} */,
  {32'h400ea384, 32'hbeb190e8} /* (3, 10, 9) {real, imag} */,
  {32'hbfd61154, 32'hbf351124} /* (3, 10, 8) {real, imag} */,
  {32'h3f01c7c8, 32'hc0ff80ea} /* (3, 10, 7) {real, imag} */,
  {32'h40b5dfd3, 32'hbfb439b8} /* (3, 10, 6) {real, imag} */,
  {32'hc0bf1d9c, 32'h4105efd7} /* (3, 10, 5) {real, imag} */,
  {32'hc055e4b6, 32'hc06a5cc0} /* (3, 10, 4) {real, imag} */,
  {32'h3f3c1140, 32'h419c9c92} /* (3, 10, 3) {real, imag} */,
  {32'h41073174, 32'h418dacff} /* (3, 10, 2) {real, imag} */,
  {32'hc09ff3b4, 32'h414b73a0} /* (3, 10, 1) {real, imag} */,
  {32'h3efe14d0, 32'h40cae7ea} /* (3, 10, 0) {real, imag} */,
  {32'h404eef29, 32'h41427f4a} /* (3, 9, 15) {real, imag} */,
  {32'h40fbff46, 32'h40d3cd36} /* (3, 9, 14) {real, imag} */,
  {32'h411513a3, 32'h3e718140} /* (3, 9, 13) {real, imag} */,
  {32'hbfd947ca, 32'hc0bd8057} /* (3, 9, 12) {real, imag} */,
  {32'hc006db86, 32'hc043b780} /* (3, 9, 11) {real, imag} */,
  {32'h400cbd4b, 32'h402c3a45} /* (3, 9, 10) {real, imag} */,
  {32'hbeb461e0, 32'hc098e476} /* (3, 9, 9) {real, imag} */,
  {32'hbf858790, 32'h40074570} /* (3, 9, 8) {real, imag} */,
  {32'hbee49470, 32'h404e1d66} /* (3, 9, 7) {real, imag} */,
  {32'h3f60da5c, 32'h40e0bc5e} /* (3, 9, 6) {real, imag} */,
  {32'h410c9b20, 32'h4061653c} /* (3, 9, 5) {real, imag} */,
  {32'hbffd435e, 32'h40d913c5} /* (3, 9, 4) {real, imag} */,
  {32'hc0cf860a, 32'hc1499380} /* (3, 9, 3) {real, imag} */,
  {32'hc10d88d1, 32'hc10278eb} /* (3, 9, 2) {real, imag} */,
  {32'h409da5f0, 32'hc0ecd5c5} /* (3, 9, 1) {real, imag} */,
  {32'hc1317a88, 32'hbff257d5} /* (3, 9, 0) {real, imag} */,
  {32'h40dd2d56, 32'h40f18d8b} /* (3, 8, 15) {real, imag} */,
  {32'hc011cc2c, 32'h3f4b7310} /* (3, 8, 14) {real, imag} */,
  {32'hbf99c8b0, 32'h408cd0b8} /* (3, 8, 13) {real, imag} */,
  {32'h40070231, 32'h3f0f6cee} /* (3, 8, 12) {real, imag} */,
  {32'hc1003160, 32'hc097ee6a} /* (3, 8, 11) {real, imag} */,
  {32'h40488a2e, 32'hc058a754} /* (3, 8, 10) {real, imag} */,
  {32'h4093f186, 32'hc0cfeab6} /* (3, 8, 9) {real, imag} */,
  {32'hc024b812, 32'hbe625f50} /* (3, 8, 8) {real, imag} */,
  {32'h3fdf92b6, 32'h3ecaf6e0} /* (3, 8, 7) {real, imag} */,
  {32'hc022f94e, 32'h3f1f2040} /* (3, 8, 6) {real, imag} */,
  {32'h4015e0c0, 32'hbf6159cc} /* (3, 8, 5) {real, imag} */,
  {32'h40e48276, 32'h4076e618} /* (3, 8, 4) {real, imag} */,
  {32'h40a76f64, 32'h413b5e3a} /* (3, 8, 3) {real, imag} */,
  {32'hc041e014, 32'hc100df34} /* (3, 8, 2) {real, imag} */,
  {32'hc0980582, 32'hc08b5f1d} /* (3, 8, 1) {real, imag} */,
  {32'h3fed900c, 32'hc096ef3a} /* (3, 8, 0) {real, imag} */,
  {32'hc03269a8, 32'hc139026b} /* (3, 7, 15) {real, imag} */,
  {32'h41906e87, 32'h407eaa59} /* (3, 7, 14) {real, imag} */,
  {32'h40e8b9b7, 32'h40dec6e3} /* (3, 7, 13) {real, imag} */,
  {32'hc03b3bc0, 32'hbe147778} /* (3, 7, 12) {real, imag} */,
  {32'hbf36ada6, 32'hbf3f24e6} /* (3, 7, 11) {real, imag} */,
  {32'h407674c2, 32'h3edb956c} /* (3, 7, 10) {real, imag} */,
  {32'hbece70d0, 32'h3fcbe05e} /* (3, 7, 9) {real, imag} */,
  {32'hc08543a3, 32'h3e21c470} /* (3, 7, 8) {real, imag} */,
  {32'h409460c2, 32'h3fe9059a} /* (3, 7, 7) {real, imag} */,
  {32'hc07c2e02, 32'hc0132e18} /* (3, 7, 6) {real, imag} */,
  {32'hc008e8d2, 32'h400ee5b2} /* (3, 7, 5) {real, imag} */,
  {32'h40a31d54, 32'hc072a9da} /* (3, 7, 4) {real, imag} */,
  {32'h40ae8891, 32'hc157238e} /* (3, 7, 3) {real, imag} */,
  {32'h3f1167a0, 32'h404f9a6f} /* (3, 7, 2) {real, imag} */,
  {32'hc144b3f4, 32'hc0dbea0a} /* (3, 7, 1) {real, imag} */,
  {32'h3ddce840, 32'h3f7205c4} /* (3, 7, 0) {real, imag} */,
  {32'hc1b25cb9, 32'hc17714e0} /* (3, 6, 15) {real, imag} */,
  {32'h3f7de5c8, 32'hc04cc454} /* (3, 6, 14) {real, imag} */,
  {32'hbf65474e, 32'hc00fe015} /* (3, 6, 13) {real, imag} */,
  {32'hbf858b14, 32'hc0a37dc2} /* (3, 6, 12) {real, imag} */,
  {32'h41008dbb, 32'hc10b472a} /* (3, 6, 11) {real, imag} */,
  {32'h3f3ae0e0, 32'h406fa8cc} /* (3, 6, 10) {real, imag} */,
  {32'hbfe81970, 32'h4045eb02} /* (3, 6, 9) {real, imag} */,
  {32'hc0009e8c, 32'hc0899ed8} /* (3, 6, 8) {real, imag} */,
  {32'h40acb052, 32'h4000aa1e} /* (3, 6, 7) {real, imag} */,
  {32'h3f38f02c, 32'hbf9aed2f} /* (3, 6, 6) {real, imag} */,
  {32'h40dbfd55, 32'hbedbd1f0} /* (3, 6, 5) {real, imag} */,
  {32'hc1268486, 32'h4182913a} /* (3, 6, 4) {real, imag} */,
  {32'h3fe53647, 32'hbe8170c8} /* (3, 6, 3) {real, imag} */,
  {32'h40bba311, 32'hc0ce70da} /* (3, 6, 2) {real, imag} */,
  {32'h4098279c, 32'h41761068} /* (3, 6, 1) {real, imag} */,
  {32'hc1b169ee, 32'hbfa2563f} /* (3, 6, 0) {real, imag} */,
  {32'h41b4c7c9, 32'hc1a32764} /* (3, 5, 15) {real, imag} */,
  {32'h40564ebb, 32'h409099a2} /* (3, 5, 14) {real, imag} */,
  {32'hc183ceb6, 32'hc217bb5c} /* (3, 5, 13) {real, imag} */,
  {32'hbf802140, 32'h4085edb4} /* (3, 5, 12) {real, imag} */,
  {32'hbe5430d0, 32'h4188798e} /* (3, 5, 11) {real, imag} */,
  {32'hc0b2e9ee, 32'h40fde09f} /* (3, 5, 10) {real, imag} */,
  {32'h40e043d7, 32'h4033d08a} /* (3, 5, 9) {real, imag} */,
  {32'h3f4ffb08, 32'hc023c060} /* (3, 5, 8) {real, imag} */,
  {32'hc06e2616, 32'h3ec91950} /* (3, 5, 7) {real, imag} */,
  {32'h404c3761, 32'h40c10dfb} /* (3, 5, 6) {real, imag} */,
  {32'hc07f0f03, 32'hc067b304} /* (3, 5, 5) {real, imag} */,
  {32'hc206c270, 32'h41bcf7e7} /* (3, 5, 4) {real, imag} */,
  {32'hc0a48bf8, 32'hc0ba4c30} /* (3, 5, 3) {real, imag} */,
  {32'hc0989c85, 32'h41074efa} /* (3, 5, 2) {real, imag} */,
  {32'h40b7c010, 32'h414de370} /* (3, 5, 1) {real, imag} */,
  {32'hc04c1e2a, 32'hc21a2e60} /* (3, 5, 0) {real, imag} */,
  {32'h4139dc2c, 32'hbf5e9770} /* (3, 4, 15) {real, imag} */,
  {32'h41f60936, 32'h416b1660} /* (3, 4, 14) {real, imag} */,
  {32'hc0ac40be, 32'h41dfc92f} /* (3, 4, 13) {real, imag} */,
  {32'hbefea980, 32'hc22332b0} /* (3, 4, 12) {real, imag} */,
  {32'hbf167140, 32'h4106e53c} /* (3, 4, 11) {real, imag} */,
  {32'h401dfec0, 32'hbff59801} /* (3, 4, 10) {real, imag} */,
  {32'hbfb27a78, 32'hc0000aa4} /* (3, 4, 9) {real, imag} */,
  {32'h408c58e8, 32'h40186ef8} /* (3, 4, 8) {real, imag} */,
  {32'hbff761a8, 32'hc0ef0582} /* (3, 4, 7) {real, imag} */,
  {32'h417de4c2, 32'h40498654} /* (3, 4, 6) {real, imag} */,
  {32'hc15a9d88, 32'hbff2f260} /* (3, 4, 5) {real, imag} */,
  {32'hc1952448, 32'h40b7a1ac} /* (3, 4, 4) {real, imag} */,
  {32'hc0cc4c12, 32'h40d731bc} /* (3, 4, 3) {real, imag} */,
  {32'h3e5c2180, 32'hc1746f8c} /* (3, 4, 2) {real, imag} */,
  {32'h42634d01, 32'h42015035} /* (3, 4, 1) {real, imag} */,
  {32'hc1f4f132, 32'hc1c8a349} /* (3, 4, 0) {real, imag} */,
  {32'h4028b214, 32'hc01d1ed4} /* (3, 3, 15) {real, imag} */,
  {32'h4174851b, 32'hc209a0f7} /* (3, 3, 14) {real, imag} */,
  {32'h4189716c, 32'h3f522bcc} /* (3, 3, 13) {real, imag} */,
  {32'hbfe0831e, 32'hc19ca946} /* (3, 3, 12) {real, imag} */,
  {32'h411a5c9a, 32'hc1abbc04} /* (3, 3, 11) {real, imag} */,
  {32'hc13be8c4, 32'hc0d7402a} /* (3, 3, 10) {real, imag} */,
  {32'hbf91afc8, 32'h4022e07c} /* (3, 3, 9) {real, imag} */,
  {32'h41159f56, 32'h3eff5470} /* (3, 3, 8) {real, imag} */,
  {32'hc1338301, 32'hc12a8609} /* (3, 3, 7) {real, imag} */,
  {32'hbf3c5b40, 32'hc1b42318} /* (3, 3, 6) {real, imag} */,
  {32'hc201bf2a, 32'h4102a310} /* (3, 3, 5) {real, imag} */,
  {32'h40903314, 32'hc1c71f22} /* (3, 3, 4) {real, imag} */,
  {32'hc180c370, 32'hc1009fcb} /* (3, 3, 3) {real, imag} */,
  {32'h3ec20aa0, 32'h41fbddfb} /* (3, 3, 2) {real, imag} */,
  {32'hc1c5d7ce, 32'hc1a11af8} /* (3, 3, 1) {real, imag} */,
  {32'h41c10305, 32'h41594e96} /* (3, 3, 0) {real, imag} */,
  {32'h41f6b1d4, 32'h4271093e} /* (3, 2, 15) {real, imag} */,
  {32'h42415fcb, 32'h42271aca} /* (3, 2, 14) {real, imag} */,
  {32'h415e5d39, 32'hc21f3039} /* (3, 2, 13) {real, imag} */,
  {32'h41a21650, 32'hbef4f7d0} /* (3, 2, 12) {real, imag} */,
  {32'hc103f459, 32'h41f5620c} /* (3, 2, 11) {real, imag} */,
  {32'h407f4db8, 32'h40a966ab} /* (3, 2, 10) {real, imag} */,
  {32'h3f979666, 32'hbf89fe10} /* (3, 2, 9) {real, imag} */,
  {32'h406f3394, 32'h407454fe} /* (3, 2, 8) {real, imag} */,
  {32'h3fb5fd66, 32'h3f403800} /* (3, 2, 7) {real, imag} */,
  {32'hc0c77bc4, 32'h404bb6d6} /* (3, 2, 6) {real, imag} */,
  {32'h418ef824, 32'hc07b4c9c} /* (3, 2, 5) {real, imag} */,
  {32'h41cc8714, 32'h40cb016f} /* (3, 2, 4) {real, imag} */,
  {32'hc127ea23, 32'hc127964d} /* (3, 2, 3) {real, imag} */,
  {32'h420ca311, 32'hc216ea6c} /* (3, 2, 2) {real, imag} */,
  {32'hc1994746, 32'h3e835800} /* (3, 2, 1) {real, imag} */,
  {32'hc20b9ce1, 32'hc135dec6} /* (3, 2, 0) {real, imag} */,
  {32'h419510cc, 32'hc19b8792} /* (3, 1, 15) {real, imag} */,
  {32'hc2466422, 32'hc14bee7b} /* (3, 1, 14) {real, imag} */,
  {32'hc1a2230e, 32'hc1c48822} /* (3, 1, 13) {real, imag} */,
  {32'h411cdefa, 32'hbdc32180} /* (3, 1, 12) {real, imag} */,
  {32'hc10b8d8b, 32'h406de004} /* (3, 1, 11) {real, imag} */,
  {32'hc0921318, 32'h410a5b2d} /* (3, 1, 10) {real, imag} */,
  {32'hc1ae5955, 32'hc06d959c} /* (3, 1, 9) {real, imag} */,
  {32'hc005aa7c, 32'h40ff2808} /* (3, 1, 8) {real, imag} */,
  {32'h3f892850, 32'hc06b92ac} /* (3, 1, 7) {real, imag} */,
  {32'h414fbc4e, 32'hc1d3540c} /* (3, 1, 6) {real, imag} */,
  {32'h40177234, 32'h40d8a68a} /* (3, 1, 5) {real, imag} */,
  {32'hc0c750e4, 32'h40b046ce} /* (3, 1, 4) {real, imag} */,
  {32'h4237f9b7, 32'h4204cd18} /* (3, 1, 3) {real, imag} */,
  {32'h41a5ac94, 32'hc1673f47} /* (3, 1, 2) {real, imag} */,
  {32'hc22a0c99, 32'h42044c5c} /* (3, 1, 1) {real, imag} */,
  {32'hc1c2af30, 32'h421ac383} /* (3, 1, 0) {real, imag} */,
  {32'hc05e9dc8, 32'h425b8878} /* (3, 0, 15) {real, imag} */,
  {32'h425544d8, 32'h41ad18b8} /* (3, 0, 14) {real, imag} */,
  {32'h41a27adc, 32'hc110fb86} /* (3, 0, 13) {real, imag} */,
  {32'hc242f0eb, 32'hc21875da} /* (3, 0, 12) {real, imag} */,
  {32'h408867cb, 32'h421c2e24} /* (3, 0, 11) {real, imag} */,
  {32'hbf965060, 32'h3f3ade50} /* (3, 0, 10) {real, imag} */,
  {32'h406319e6, 32'hc0928dda} /* (3, 0, 9) {real, imag} */,
  {32'hc093988a, 32'h416a368e} /* (3, 0, 8) {real, imag} */,
  {32'h419aa66d, 32'h3d1cb300} /* (3, 0, 7) {real, imag} */,
  {32'hc1049e7a, 32'h41065c71} /* (3, 0, 6) {real, imag} */,
  {32'hc0524c96, 32'hc2586c30} /* (3, 0, 5) {real, imag} */,
  {32'hc0db4f48, 32'h415c696d} /* (3, 0, 4) {real, imag} */,
  {32'hc10a0884, 32'h41eb360d} /* (3, 0, 3) {real, imag} */,
  {32'h40331420, 32'h40b49636} /* (3, 0, 2) {real, imag} */,
  {32'h41a704d9, 32'hc20ba1cc} /* (3, 0, 1) {real, imag} */,
  {32'h41d7bf2c, 32'hc256a928} /* (3, 0, 0) {real, imag} */,
  {32'h3e5b6980, 32'h42223bfa} /* (2, 15, 15) {real, imag} */,
  {32'h428c82b2, 32'hc0722588} /* (2, 15, 14) {real, imag} */,
  {32'h417b116b, 32'hc1d7e04a} /* (2, 15, 13) {real, imag} */,
  {32'hc18e73f4, 32'h40626170} /* (2, 15, 12) {real, imag} */,
  {32'hc01ce18c, 32'h400f5402} /* (2, 15, 11) {real, imag} */,
  {32'hc08d6720, 32'h3ed1c3d0} /* (2, 15, 10) {real, imag} */,
  {32'hbb77f800, 32'h413082d6} /* (2, 15, 9) {real, imag} */,
  {32'hc0909f30, 32'h3fb8a120} /* (2, 15, 8) {real, imag} */,
  {32'hc0d4a449, 32'h417fac14} /* (2, 15, 7) {real, imag} */,
  {32'h3fb669e0, 32'hc122051a} /* (2, 15, 6) {real, imag} */,
  {32'hc04b8cc8, 32'h40ba4967} /* (2, 15, 5) {real, imag} */,
  {32'h4084d230, 32'h4288d994} /* (2, 15, 4) {real, imag} */,
  {32'hbd563200, 32'hc1928b44} /* (2, 15, 3) {real, imag} */,
  {32'hc13a757e, 32'hc1ad7761} /* (2, 15, 2) {real, imag} */,
  {32'hc1d1700b, 32'h419e1e8f} /* (2, 15, 1) {real, imag} */,
  {32'hc28fbf47, 32'hc0f7aa88} /* (2, 15, 0) {real, imag} */,
  {32'hc2ee3c8f, 32'h413b1768} /* (2, 14, 15) {real, imag} */,
  {32'h40a3e5a8, 32'h420a919a} /* (2, 14, 14) {real, imag} */,
  {32'h428156bf, 32'h4131335c} /* (2, 14, 13) {real, imag} */,
  {32'hc0c4b37e, 32'hc18676ba} /* (2, 14, 12) {real, imag} */,
  {32'h4165dcd4, 32'h411fab24} /* (2, 14, 11) {real, imag} */,
  {32'h40376b30, 32'h40cf3270} /* (2, 14, 10) {real, imag} */,
  {32'hbfc1d400, 32'h40cdf774} /* (2, 14, 9) {real, imag} */,
  {32'h3e0fde40, 32'hbf90a658} /* (2, 14, 8) {real, imag} */,
  {32'hc047a8e0, 32'hc072e128} /* (2, 14, 7) {real, imag} */,
  {32'h3e8c8640, 32'h402ee1b8} /* (2, 14, 6) {real, imag} */,
  {32'hc0be98d8, 32'h40d33af0} /* (2, 14, 5) {real, imag} */,
  {32'hc07dffbb, 32'h4202ab60} /* (2, 14, 4) {real, imag} */,
  {32'h40c48ad0, 32'hc20bbe34} /* (2, 14, 3) {real, imag} */,
  {32'h4235ef21, 32'hc1d77a00} /* (2, 14, 2) {real, imag} */,
  {32'h42380652, 32'hc289f407} /* (2, 14, 1) {real, imag} */,
  {32'hc18178da, 32'hc120cbef} /* (2, 14, 0) {real, imag} */,
  {32'hc17d74b6, 32'hbe7daf00} /* (2, 13, 15) {real, imag} */,
  {32'h40ae4b52, 32'h409ea176} /* (2, 13, 14) {real, imag} */,
  {32'h4225da82, 32'h40e4da06} /* (2, 13, 13) {real, imag} */,
  {32'h42309db0, 32'h412c76ae} /* (2, 13, 12) {real, imag} */,
  {32'hc163d1fc, 32'hbf889c78} /* (2, 13, 11) {real, imag} */,
  {32'hc0d11f1f, 32'h409c8578} /* (2, 13, 10) {real, imag} */,
  {32'hc155dcf0, 32'h4086f27e} /* (2, 13, 9) {real, imag} */,
  {32'hc0adea24, 32'h3ff5ab00} /* (2, 13, 8) {real, imag} */,
  {32'h40ce278f, 32'h4136240d} /* (2, 13, 7) {real, imag} */,
  {32'h40e996d3, 32'hc1694e56} /* (2, 13, 6) {real, imag} */,
  {32'h417ab70e, 32'hc1754c1d} /* (2, 13, 5) {real, imag} */,
  {32'h40581f10, 32'h421511ac} /* (2, 13, 4) {real, imag} */,
  {32'h3fc72570, 32'hc1845f42} /* (2, 13, 3) {real, imag} */,
  {32'h407df718, 32'h417d1573} /* (2, 13, 2) {real, imag} */,
  {32'h41843379, 32'h423130fd} /* (2, 13, 1) {real, imag} */,
  {32'hc0d4e114, 32'hc0cd5258} /* (2, 13, 0) {real, imag} */,
  {32'hc065b022, 32'h40a73d94} /* (2, 12, 15) {real, imag} */,
  {32'hc10c658a, 32'hc1567c88} /* (2, 12, 14) {real, imag} */,
  {32'h40a82a24, 32'h428ed2ab} /* (2, 12, 13) {real, imag} */,
  {32'hbfc63f90, 32'hc082c864} /* (2, 12, 12) {real, imag} */,
  {32'h422570a8, 32'hc138bf74} /* (2, 12, 11) {real, imag} */,
  {32'hc0d23bd2, 32'h405c446e} /* (2, 12, 10) {real, imag} */,
  {32'h3f9e286c, 32'h404e3060} /* (2, 12, 9) {real, imag} */,
  {32'hc128eb9c, 32'h404ab5ca} /* (2, 12, 8) {real, imag} */,
  {32'h40e72a73, 32'hc1106a78} /* (2, 12, 7) {real, imag} */,
  {32'h40e5df4c, 32'hc0c75ed3} /* (2, 12, 6) {real, imag} */,
  {32'hbfb73a60, 32'hc1c44544} /* (2, 12, 5) {real, imag} */,
  {32'h41cca24d, 32'h42316056} /* (2, 12, 4) {real, imag} */,
  {32'h416e0e12, 32'hc1ab5713} /* (2, 12, 3) {real, imag} */,
  {32'hc0285aee, 32'hc12ea678} /* (2, 12, 2) {real, imag} */,
  {32'h4183ab64, 32'hc2406d4a} /* (2, 12, 1) {real, imag} */,
  {32'h40d46ab0, 32'h413ca828} /* (2, 12, 0) {real, imag} */,
  {32'h41e4b06a, 32'hc21cf754} /* (2, 11, 15) {real, imag} */,
  {32'h40ab9aa8, 32'hc1a44720} /* (2, 11, 14) {real, imag} */,
  {32'hc04cf404, 32'h414eecb3} /* (2, 11, 13) {real, imag} */,
  {32'hc11e5022, 32'hc10741fc} /* (2, 11, 12) {real, imag} */,
  {32'hc0d5cb70, 32'h41132347} /* (2, 11, 11) {real, imag} */,
  {32'h4120dad8, 32'h41414f38} /* (2, 11, 10) {real, imag} */,
  {32'h409cd29a, 32'hc0d62976} /* (2, 11, 9) {real, imag} */,
  {32'h3ebcb670, 32'hc056ea0c} /* (2, 11, 8) {real, imag} */,
  {32'h40fddca6, 32'h4120cb93} /* (2, 11, 7) {real, imag} */,
  {32'h4134c268, 32'h400cb856} /* (2, 11, 6) {real, imag} */,
  {32'hc0b5530e, 32'h4007e77c} /* (2, 11, 5) {real, imag} */,
  {32'h4154740a, 32'hc0ed4b0a} /* (2, 11, 4) {real, imag} */,
  {32'hc0340200, 32'hc1292e51} /* (2, 11, 3) {real, imag} */,
  {32'hc1c4f90a, 32'h411e2e06} /* (2, 11, 2) {real, imag} */,
  {32'hbfd1bd78, 32'hc1175bd7} /* (2, 11, 1) {real, imag} */,
  {32'h4140625e, 32'h41cddfc4} /* (2, 11, 0) {real, imag} */,
  {32'hc0e8ee06, 32'h412e18ba} /* (2, 10, 15) {real, imag} */,
  {32'hc1ac8b91, 32'hc06ee2a3} /* (2, 10, 14) {real, imag} */,
  {32'hc10e48fe, 32'hbfb8954a} /* (2, 10, 13) {real, imag} */,
  {32'h404200d9, 32'h417f8d38} /* (2, 10, 12) {real, imag} */,
  {32'hc0030ec8, 32'hc03f37c9} /* (2, 10, 11) {real, imag} */,
  {32'hc0a6b21f, 32'h3ebe276e} /* (2, 10, 10) {real, imag} */,
  {32'hc03e041e, 32'hbfc330b1} /* (2, 10, 9) {real, imag} */,
  {32'hc02a4e86, 32'hc0228e52} /* (2, 10, 8) {real, imag} */,
  {32'hbfb13d14, 32'hc07e6d22} /* (2, 10, 7) {real, imag} */,
  {32'h40a1d87d, 32'h3f82b83e} /* (2, 10, 6) {real, imag} */,
  {32'h40d9b746, 32'h409424cc} /* (2, 10, 5) {real, imag} */,
  {32'hc12df440, 32'hc12cb880} /* (2, 10, 4) {real, imag} */,
  {32'h4177af2e, 32'h40a97d4a} /* (2, 10, 3) {real, imag} */,
  {32'hc0d4571c, 32'hbf7f2df4} /* (2, 10, 2) {real, imag} */,
  {32'h41654eb5, 32'h3f9239e0} /* (2, 10, 1) {real, imag} */,
  {32'h414bc9d8, 32'h40c185db} /* (2, 10, 0) {real, imag} */,
  {32'hc0d99dd5, 32'hbf6b6da2} /* (2, 9, 15) {real, imag} */,
  {32'hbdd4f3f0, 32'hc0c276fa} /* (2, 9, 14) {real, imag} */,
  {32'h3fc3af9c, 32'hc1243443} /* (2, 9, 13) {real, imag} */,
  {32'h40bb633b, 32'hc1007b94} /* (2, 9, 12) {real, imag} */,
  {32'h3f5da9e8, 32'hc110cae3} /* (2, 9, 11) {real, imag} */,
  {32'hc0c772bd, 32'hc044d5ec} /* (2, 9, 10) {real, imag} */,
  {32'h3e466eb8, 32'hbe8a159d} /* (2, 9, 9) {real, imag} */,
  {32'h4083c091, 32'hc02068ec} /* (2, 9, 8) {real, imag} */,
  {32'hbfa4b65b, 32'hbf25b396} /* (2, 9, 7) {real, imag} */,
  {32'hc0b28cdd, 32'h3f626d32} /* (2, 9, 6) {real, imag} */,
  {32'hc129a284, 32'hbe2e90c0} /* (2, 9, 5) {real, imag} */,
  {32'hc13cf89a, 32'h40073dc6} /* (2, 9, 4) {real, imag} */,
  {32'h4181ef6a, 32'h407cf224} /* (2, 9, 3) {real, imag} */,
  {32'hc01d46ec, 32'h41196fa7} /* (2, 9, 2) {real, imag} */,
  {32'hc10520e2, 32'hbf39f2ba} /* (2, 9, 1) {real, imag} */,
  {32'h40d8a925, 32'hc0b61f80} /* (2, 9, 0) {real, imag} */,
  {32'hc11cf7d6, 32'hc026767a} /* (2, 8, 15) {real, imag} */,
  {32'hc18b3c2c, 32'h41846da2} /* (2, 8, 14) {real, imag} */,
  {32'hc1375e44, 32'hc0742313} /* (2, 8, 13) {real, imag} */,
  {32'hc0ed7ed0, 32'h40f4a250} /* (2, 8, 12) {real, imag} */,
  {32'hc0c31c29, 32'h3fd78398} /* (2, 8, 11) {real, imag} */,
  {32'h3f72d420, 32'hbf3aae88} /* (2, 8, 10) {real, imag} */,
  {32'h400fb2ef, 32'h400f0fea} /* (2, 8, 9) {real, imag} */,
  {32'hbf3030ba, 32'hc000201e} /* (2, 8, 8) {real, imag} */,
  {32'h3e05f430, 32'h3fb9c378} /* (2, 8, 7) {real, imag} */,
  {32'h405356bc, 32'h3fb69fd4} /* (2, 8, 6) {real, imag} */,
  {32'h4104e9ea, 32'h4084fea1} /* (2, 8, 5) {real, imag} */,
  {32'hc0d41594, 32'h4166de5c} /* (2, 8, 4) {real, imag} */,
  {32'hc130f8f0, 32'hc1037a49} /* (2, 8, 3) {real, imag} */,
  {32'h409c996f, 32'hc08ddc50} /* (2, 8, 2) {real, imag} */,
  {32'h4180c725, 32'h3fd70f10} /* (2, 8, 1) {real, imag} */,
  {32'h3f0f5002, 32'h415c57cc} /* (2, 8, 0) {real, imag} */,
  {32'hc0d45fa8, 32'hc0d38c9c} /* (2, 7, 15) {real, imag} */,
  {32'hc0875264, 32'hc0e686b8} /* (2, 7, 14) {real, imag} */,
  {32'h40b68ff4, 32'h40db02fd} /* (2, 7, 13) {real, imag} */,
  {32'hc100ec3a, 32'h400f0418} /* (2, 7, 12) {real, imag} */,
  {32'h40d3b02d, 32'h4011e9c0} /* (2, 7, 11) {real, imag} */,
  {32'h40b13e3c, 32'hc0df89b6} /* (2, 7, 10) {real, imag} */,
  {32'h400e9404, 32'hc058e4ac} /* (2, 7, 9) {real, imag} */,
  {32'hbf1da458, 32'h3e127f50} /* (2, 7, 8) {real, imag} */,
  {32'hbf26e9c2, 32'hc08f1b92} /* (2, 7, 7) {real, imag} */,
  {32'h41585288, 32'h401a78fc} /* (2, 7, 6) {real, imag} */,
  {32'h40e95275, 32'hbfbb07f8} /* (2, 7, 5) {real, imag} */,
  {32'h3fa3b94c, 32'h40231eb8} /* (2, 7, 4) {real, imag} */,
  {32'h3fdde53a, 32'h414c68d6} /* (2, 7, 3) {real, imag} */,
  {32'hc1a6cfa8, 32'h3ef0f740} /* (2, 7, 2) {real, imag} */,
  {32'h40d46322, 32'h3f67a880} /* (2, 7, 1) {real, imag} */,
  {32'h4102d5ba, 32'hc02fab11} /* (2, 7, 0) {real, imag} */,
  {32'hc0b8cb28, 32'hc1c3c440} /* (2, 6, 15) {real, imag} */,
  {32'hbf13d898, 32'h404c0a68} /* (2, 6, 14) {real, imag} */,
  {32'hc028a172, 32'h403c8670} /* (2, 6, 13) {real, imag} */,
  {32'h4150ea0a, 32'h3e523b20} /* (2, 6, 12) {real, imag} */,
  {32'hc1958dd2, 32'hbf3d5ec8} /* (2, 6, 11) {real, imag} */,
  {32'h40f823ef, 32'h40df1864} /* (2, 6, 10) {real, imag} */,
  {32'h3fec1886, 32'h41294570} /* (2, 6, 9) {real, imag} */,
  {32'h4081f344, 32'hbf8afadc} /* (2, 6, 8) {real, imag} */,
  {32'h3fd58bda, 32'hc05d3fb7} /* (2, 6, 7) {real, imag} */,
  {32'hc09ee415, 32'h417d3258} /* (2, 6, 6) {real, imag} */,
  {32'hc175298d, 32'hbfd40c14} /* (2, 6, 5) {real, imag} */,
  {32'hc1421f0e, 32'hc078e0ce} /* (2, 6, 4) {real, imag} */,
  {32'h416242aa, 32'hc04b5140} /* (2, 6, 3) {real, imag} */,
  {32'h40f24f91, 32'hbfd043c0} /* (2, 6, 2) {real, imag} */,
  {32'h3f1406a4, 32'h41ba8e60} /* (2, 6, 1) {real, imag} */,
  {32'hc0ca4958, 32'h40f86df9} /* (2, 6, 0) {real, imag} */,
  {32'hc1783311, 32'hc05b0f3c} /* (2, 5, 15) {real, imag} */,
  {32'h41172dfa, 32'h40f389fa} /* (2, 5, 14) {real, imag} */,
  {32'h412974b6, 32'h41eaca14} /* (2, 5, 13) {real, imag} */,
  {32'hc089d339, 32'hc0526254} /* (2, 5, 12) {real, imag} */,
  {32'hc0208f87, 32'hc190f0f2} /* (2, 5, 11) {real, imag} */,
  {32'hc158c333, 32'h41cd2b78} /* (2, 5, 10) {real, imag} */,
  {32'h40296416, 32'hc11316b5} /* (2, 5, 9) {real, imag} */,
  {32'h3fd92374, 32'h3f31b5a0} /* (2, 5, 8) {real, imag} */,
  {32'hc05d3a92, 32'h3ffb2478} /* (2, 5, 7) {real, imag} */,
  {32'hc18ac8c8, 32'hbfde7b68} /* (2, 5, 6) {real, imag} */,
  {32'h40c1b4c2, 32'hc025c44c} /* (2, 5, 5) {real, imag} */,
  {32'h416500fa, 32'hc1a66fb6} /* (2, 5, 4) {real, imag} */,
  {32'hbf77e068, 32'h41bf78a0} /* (2, 5, 3) {real, imag} */,
  {32'h41d9534b, 32'h3f711f70} /* (2, 5, 2) {real, imag} */,
  {32'hc11d349b, 32'hc1d14c36} /* (2, 5, 1) {real, imag} */,
  {32'hc15623f2, 32'h41cdc296} /* (2, 5, 0) {real, imag} */,
  {32'h4204d4ed, 32'h4081b4a9} /* (2, 4, 15) {real, imag} */,
  {32'h40d5fe38, 32'h41f5d21e} /* (2, 4, 14) {real, imag} */,
  {32'hc022fc50, 32'hc135df54} /* (2, 4, 13) {real, imag} */,
  {32'hc0902360, 32'hc1a035f8} /* (2, 4, 12) {real, imag} */,
  {32'h40c7e6e4, 32'hc112a2ba} /* (2, 4, 11) {real, imag} */,
  {32'h40f779c0, 32'hc17714b1} /* (2, 4, 10) {real, imag} */,
  {32'h4113508e, 32'hc0eb31ff} /* (2, 4, 9) {real, imag} */,
  {32'h3e8347c0, 32'h4099793f} /* (2, 4, 8) {real, imag} */,
  {32'h4142ba4e, 32'h40a9b8f1} /* (2, 4, 7) {real, imag} */,
  {32'hc15c5c98, 32'h3f175330} /* (2, 4, 6) {real, imag} */,
  {32'h4195237d, 32'h410b8856} /* (2, 4, 5) {real, imag} */,
  {32'h40ba0d58, 32'hc080e4aa} /* (2, 4, 4) {real, imag} */,
  {32'hc2148acc, 32'hc1e11630} /* (2, 4, 3) {real, imag} */,
  {32'hc21e8733, 32'hc0a95f0e} /* (2, 4, 2) {real, imag} */,
  {32'hc20645f7, 32'hc0f102a7} /* (2, 4, 1) {real, imag} */,
  {32'hc20f8e40, 32'hc11eb2dc} /* (2, 4, 0) {real, imag} */,
  {32'h41912412, 32'hc1d645c7} /* (2, 3, 15) {real, imag} */,
  {32'h422665dc, 32'h416bbf58} /* (2, 3, 14) {real, imag} */,
  {32'hc0cf6568, 32'hc23352fa} /* (2, 3, 13) {real, imag} */,
  {32'hc1be1bcb, 32'hc1467be6} /* (2, 3, 12) {real, imag} */,
  {32'hc12ff221, 32'hc13340bc} /* (2, 3, 11) {real, imag} */,
  {32'hc1acde8c, 32'h416daa8e} /* (2, 3, 10) {real, imag} */,
  {32'hc13fcf34, 32'hc005ce92} /* (2, 3, 9) {real, imag} */,
  {32'hc0cc1618, 32'hc0b74daf} /* (2, 3, 8) {real, imag} */,
  {32'hc0f915b5, 32'h408629ff} /* (2, 3, 7) {real, imag} */,
  {32'hc08b52d8, 32'h4163df4e} /* (2, 3, 6) {real, imag} */,
  {32'h40ac83ee, 32'hc187a796} /* (2, 3, 5) {real, imag} */,
  {32'hc1e4ded3, 32'hc1aab835} /* (2, 3, 4) {real, imag} */,
  {32'hc21b8a4d, 32'hc0fb9d10} /* (2, 3, 3) {real, imag} */,
  {32'hbfe222b0, 32'hc05bb78e} /* (2, 3, 2) {real, imag} */,
  {32'h418a9696, 32'hc080c2a4} /* (2, 3, 1) {real, imag} */,
  {32'hc22e979a, 32'hbf016a68} /* (2, 3, 0) {real, imag} */,
  {32'h41f54117, 32'hc14956e4} /* (2, 2, 15) {real, imag} */,
  {32'hc28e554e, 32'hc237a0de} /* (2, 2, 14) {real, imag} */,
  {32'hc22d01b0, 32'h423b58e6} /* (2, 2, 13) {real, imag} */,
  {32'h3ff4c6a0, 32'h4113600a} /* (2, 2, 12) {real, imag} */,
  {32'h41297313, 32'hc2066b28} /* (2, 2, 11) {real, imag} */,
  {32'h41390208, 32'hbe9843c0} /* (2, 2, 10) {real, imag} */,
  {32'hc0df6db2, 32'h410dfe0c} /* (2, 2, 9) {real, imag} */,
  {32'hc10e4758, 32'h40049bfc} /* (2, 2, 8) {real, imag} */,
  {32'h3fa3edb8, 32'hc1f575f6} /* (2, 2, 7) {real, imag} */,
  {32'hc1c91756, 32'h418642bd} /* (2, 2, 6) {real, imag} */,
  {32'hc15eb149, 32'h410a1eb2} /* (2, 2, 5) {real, imag} */,
  {32'h4262c19f, 32'h422d035c} /* (2, 2, 4) {real, imag} */,
  {32'h420c15b8, 32'h41704b1e} /* (2, 2, 3) {real, imag} */,
  {32'hc1c08a3f, 32'h41cb093c} /* (2, 2, 2) {real, imag} */,
  {32'hc0a21bcc, 32'h4209a987} /* (2, 2, 1) {real, imag} */,
  {32'h41508b10, 32'hc12fab0b} /* (2, 2, 0) {real, imag} */,
  {32'hc0b93320, 32'hc10114b7} /* (2, 1, 15) {real, imag} */,
  {32'h41c40f08, 32'h411c3a9c} /* (2, 1, 14) {real, imag} */,
  {32'h4216ee1f, 32'hc2845f5c} /* (2, 1, 13) {real, imag} */,
  {32'hc23bf07e, 32'h41336e24} /* (2, 1, 12) {real, imag} */,
  {32'h41289d04, 32'hc07600c8} /* (2, 1, 11) {real, imag} */,
  {32'hc1c1012c, 32'h4093df00} /* (2, 1, 10) {real, imag} */,
  {32'h41029c28, 32'h4162440d} /* (2, 1, 9) {real, imag} */,
  {32'h3f0cd660, 32'hbf3552d8} /* (2, 1, 8) {real, imag} */,
  {32'h4182e992, 32'h4085d39a} /* (2, 1, 7) {real, imag} */,
  {32'hc0e7f490, 32'hbf1c8460} /* (2, 1, 6) {real, imag} */,
  {32'hc21ba7b0, 32'h411469a2} /* (2, 1, 5) {real, imag} */,
  {32'h4116018e, 32'hc1a717a4} /* (2, 1, 4) {real, imag} */,
  {32'hc0895230, 32'hc2248660} /* (2, 1, 3) {real, imag} */,
  {32'h3dd6f800, 32'h42500813} /* (2, 1, 2) {real, imag} */,
  {32'hc2b5b5de, 32'h421d1354} /* (2, 1, 1) {real, imag} */,
  {32'h42179f5a, 32'h40e214cd} /* (2, 1, 0) {real, imag} */,
  {32'h41059be1, 32'hc1528ca6} /* (2, 0, 15) {real, imag} */,
  {32'hc1b89084, 32'h40e77aee} /* (2, 0, 14) {real, imag} */,
  {32'h4232c714, 32'hc13e5d94} /* (2, 0, 13) {real, imag} */,
  {32'hc197dbd8, 32'hc0a1b388} /* (2, 0, 12) {real, imag} */,
  {32'h41afbebf, 32'hc1041c09} /* (2, 0, 11) {real, imag} */,
  {32'hc09cd18a, 32'h41c714d2} /* (2, 0, 10) {real, imag} */,
  {32'hc02e0ff9, 32'hc13d6330} /* (2, 0, 9) {real, imag} */,
  {32'h41a96fdf, 32'h410e932c} /* (2, 0, 8) {real, imag} */,
  {32'h3e0f4090, 32'hc00291b8} /* (2, 0, 7) {real, imag} */,
  {32'hc0a8bd46, 32'hbfe72888} /* (2, 0, 6) {real, imag} */,
  {32'hc229e1ac, 32'hc04c54e0} /* (2, 0, 5) {real, imag} */,
  {32'hc014a9e4, 32'hc23f50d0} /* (2, 0, 4) {real, imag} */,
  {32'hc200a110, 32'hc16e33cc} /* (2, 0, 3) {real, imag} */,
  {32'hbf4462b0, 32'h3ddd9f60} /* (2, 0, 2) {real, imag} */,
  {32'h41c53440, 32'h411637e8} /* (2, 0, 1) {real, imag} */,
  {32'h422db0f6, 32'hc2c19ee2} /* (2, 0, 0) {real, imag} */,
  {32'hc10e3a29, 32'hc11c7dc0} /* (1, 15, 15) {real, imag} */,
  {32'hc0c02a5c, 32'h4218d838} /* (1, 15, 14) {real, imag} */,
  {32'h41c66d2a, 32'hc116ddf1} /* (1, 15, 13) {real, imag} */,
  {32'hbf06f360, 32'h419579aa} /* (1, 15, 12) {real, imag} */,
  {32'hc2177989, 32'h41f4606a} /* (1, 15, 11) {real, imag} */,
  {32'h40fb1a32, 32'hc1148c84} /* (1, 15, 10) {real, imag} */,
  {32'hbf003b50, 32'hc1bfc5cb} /* (1, 15, 9) {real, imag} */,
  {32'hc15d76f1, 32'hc0b203e1} /* (1, 15, 8) {real, imag} */,
  {32'h412cce0d, 32'h407e2ce0} /* (1, 15, 7) {real, imag} */,
  {32'hc1528a7d, 32'hc19c7cc5} /* (1, 15, 6) {real, imag} */,
  {32'hc144f844, 32'h419f8692} /* (1, 15, 5) {real, imag} */,
  {32'hc15c45d8, 32'hc19f5caa} /* (1, 15, 4) {real, imag} */,
  {32'hc1a113f6, 32'hc1a43662} /* (1, 15, 3) {real, imag} */,
  {32'h424405ae, 32'h42254000} /* (1, 15, 2) {real, imag} */,
  {32'hc18fa64e, 32'h4231dcf0} /* (1, 15, 1) {real, imag} */,
  {32'hc1a41ce8, 32'h418c2583} /* (1, 15, 0) {real, imag} */,
  {32'h42633134, 32'h4216e38c} /* (1, 14, 15) {real, imag} */,
  {32'hc22dff6c, 32'hc289d3a4} /* (1, 14, 14) {real, imag} */,
  {32'hc15e5f76, 32'hc1aa77da} /* (1, 14, 13) {real, imag} */,
  {32'hc1f70410, 32'h4138c824} /* (1, 14, 12) {real, imag} */,
  {32'h40d11c83, 32'hc1d90acc} /* (1, 14, 11) {real, imag} */,
  {32'h40e2500c, 32'h41acd13e} /* (1, 14, 10) {real, imag} */,
  {32'h41ec9c57, 32'hc0a77af8} /* (1, 14, 9) {real, imag} */,
  {32'hc10c60d4, 32'h404f3490} /* (1, 14, 8) {real, imag} */,
  {32'h41d64b23, 32'h41a83600} /* (1, 14, 7) {real, imag} */,
  {32'hc1560f3e, 32'h40e96586} /* (1, 14, 6) {real, imag} */,
  {32'hc16bc5ec, 32'h4116b4b0} /* (1, 14, 5) {real, imag} */,
  {32'hc170eea1, 32'hc1b5d092} /* (1, 14, 4) {real, imag} */,
  {32'h4219384e, 32'h42384dbf} /* (1, 14, 3) {real, imag} */,
  {32'hc273f7b2, 32'hbe173200} /* (1, 14, 2) {real, imag} */,
  {32'hc2bc284e, 32'hc17e6fae} /* (1, 14, 1) {real, imag} */,
  {32'h416d9004, 32'hc22679af} /* (1, 14, 0) {real, imag} */,
  {32'h4204f4e7, 32'h4104f22e} /* (1, 13, 15) {real, imag} */,
  {32'hbf3b9260, 32'hc1e76a14} /* (1, 13, 14) {real, imag} */,
  {32'hc13f527e, 32'h42524ec8} /* (1, 13, 13) {real, imag} */,
  {32'hc205602e, 32'h4109bd05} /* (1, 13, 12) {real, imag} */,
  {32'h40d1e588, 32'hc1a5300f} /* (1, 13, 11) {real, imag} */,
  {32'hbfac3850, 32'h40ff2438} /* (1, 13, 10) {real, imag} */,
  {32'hc111bd5e, 32'h41e84cdc} /* (1, 13, 9) {real, imag} */,
  {32'hc0d26726, 32'hc18b343e} /* (1, 13, 8) {real, imag} */,
  {32'h3f5c9598, 32'h4170746f} /* (1, 13, 7) {real, imag} */,
  {32'h40cd8f0e, 32'hbf985520} /* (1, 13, 6) {real, imag} */,
  {32'hc15b9b3c, 32'h40e0b06b} /* (1, 13, 5) {real, imag} */,
  {32'h416ced70, 32'h412a200b} /* (1, 13, 4) {real, imag} */,
  {32'hc165c1b2, 32'hc26b8634} /* (1, 13, 3) {real, imag} */,
  {32'hc1a6fb5d, 32'h423b09ce} /* (1, 13, 2) {real, imag} */,
  {32'h42216891, 32'h40e01888} /* (1, 13, 1) {real, imag} */,
  {32'hc1dfc068, 32'h42357727} /* (1, 13, 0) {real, imag} */,
  {32'h3f2377a0, 32'h42a1c804} /* (1, 12, 15) {real, imag} */,
  {32'hc25df15c, 32'h41f797b0} /* (1, 12, 14) {real, imag} */,
  {32'hc13095b5, 32'h4220d047} /* (1, 12, 13) {real, imag} */,
  {32'h41833910, 32'h40e40467} /* (1, 12, 12) {real, imag} */,
  {32'hbf893e58, 32'hc1ba3e68} /* (1, 12, 11) {real, imag} */,
  {32'hc00e4504, 32'hbf98de54} /* (1, 12, 10) {real, imag} */,
  {32'hc190be6e, 32'hc0a368b6} /* (1, 12, 9) {real, imag} */,
  {32'h401e2402, 32'h40ad8c90} /* (1, 12, 8) {real, imag} */,
  {32'hc07c05b8, 32'hc18a95e8} /* (1, 12, 7) {real, imag} */,
  {32'h40e6ce56, 32'h409fabf3} /* (1, 12, 6) {real, imag} */,
  {32'hc13611d5, 32'h41277387} /* (1, 12, 5) {real, imag} */,
  {32'hc1226445, 32'hc0038c26} /* (1, 12, 4) {real, imag} */,
  {32'h4096f502, 32'hc0d35928} /* (1, 12, 3) {real, imag} */,
  {32'h40bfade4, 32'h3f6986c0} /* (1, 12, 2) {real, imag} */,
  {32'h412501f4, 32'hc18a4176} /* (1, 12, 1) {real, imag} */,
  {32'hc0994c85, 32'hc2287cd6} /* (1, 12, 0) {real, imag} */,
  {32'h410a863e, 32'hc1b0cc1b} /* (1, 11, 15) {real, imag} */,
  {32'hc1547268, 32'h4110a312} /* (1, 11, 14) {real, imag} */,
  {32'h416d716c, 32'hc1031dcb} /* (1, 11, 13) {real, imag} */,
  {32'h40c2d41e, 32'hbf310510} /* (1, 11, 12) {real, imag} */,
  {32'h40e763f1, 32'hc1610fc0} /* (1, 11, 11) {real, imag} */,
  {32'hc10b94f1, 32'h412762d8} /* (1, 11, 10) {real, imag} */,
  {32'h40ded75c, 32'h40fea416} /* (1, 11, 9) {real, imag} */,
  {32'h402e64e8, 32'h405eb708} /* (1, 11, 8) {real, imag} */,
  {32'h3fa3bf08, 32'hc1115ebd} /* (1, 11, 7) {real, imag} */,
  {32'h40640f58, 32'h40ff6309} /* (1, 11, 6) {real, imag} */,
  {32'h414b36d8, 32'h403998e8} /* (1, 11, 5) {real, imag} */,
  {32'hbf1843a4, 32'h418b1fa6} /* (1, 11, 4) {real, imag} */,
  {32'h42211f65, 32'h419f1e5a} /* (1, 11, 3) {real, imag} */,
  {32'hc037e33e, 32'h41a7ce35} /* (1, 11, 2) {real, imag} */,
  {32'h41cd3991, 32'hc16aeb62} /* (1, 11, 1) {real, imag} */,
  {32'hc191af2d, 32'h3f931c60} /* (1, 11, 0) {real, imag} */,
  {32'h41af3d6a, 32'hc1625c1e} /* (1, 10, 15) {real, imag} */,
  {32'hc134e73a, 32'hc022e24b} /* (1, 10, 14) {real, imag} */,
  {32'hc0d29ba5, 32'hc1c311a8} /* (1, 10, 13) {real, imag} */,
  {32'hc1802ff4, 32'hc100fd66} /* (1, 10, 12) {real, imag} */,
  {32'hbfbbc674, 32'h417b718e} /* (1, 10, 11) {real, imag} */,
  {32'h40985e22, 32'h40f83755} /* (1, 10, 10) {real, imag} */,
  {32'h400a873c, 32'hc08ce803} /* (1, 10, 9) {real, imag} */,
  {32'h40b29870, 32'hc0024ac0} /* (1, 10, 8) {real, imag} */,
  {32'hc0aced1a, 32'h40c804ef} /* (1, 10, 7) {real, imag} */,
  {32'hc13f6ccf, 32'hc13100b2} /* (1, 10, 6) {real, imag} */,
  {32'hc0c225e7, 32'h3f8e408c} /* (1, 10, 5) {real, imag} */,
  {32'h4186e88c, 32'h402da328} /* (1, 10, 4) {real, imag} */,
  {32'hbf544838, 32'hbfed7520} /* (1, 10, 3) {real, imag} */,
  {32'hbfd9be24, 32'hc10fcf98} /* (1, 10, 2) {real, imag} */,
  {32'h417eda64, 32'hc1d22131} /* (1, 10, 1) {real, imag} */,
  {32'h413a0220, 32'h3c49f800} /* (1, 10, 0) {real, imag} */,
  {32'h40fec014, 32'h40ebe77b} /* (1, 9, 15) {real, imag} */,
  {32'hc104d88b, 32'hc0cc379a} /* (1, 9, 14) {real, imag} */,
  {32'hc02ff60e, 32'h4183d6c6} /* (1, 9, 13) {real, imag} */,
  {32'h405754bf, 32'hc0149158} /* (1, 9, 12) {real, imag} */,
  {32'h409be5a9, 32'h40f7c011} /* (1, 9, 11) {real, imag} */,
  {32'hbff789b5, 32'hc04c19ac} /* (1, 9, 10) {real, imag} */,
  {32'h3e74f58c, 32'hc0ccdacc} /* (1, 9, 9) {real, imag} */,
  {32'h401a46b0, 32'h3ff4a38c} /* (1, 9, 8) {real, imag} */,
  {32'hbf2ce6d3, 32'h3edf3240} /* (1, 9, 7) {real, imag} */,
  {32'h40b0ef99, 32'hc084df52} /* (1, 9, 6) {real, imag} */,
  {32'hc0951dc1, 32'hc0f33ec7} /* (1, 9, 5) {real, imag} */,
  {32'hc088ff92, 32'hc1a09f62} /* (1, 9, 4) {real, imag} */,
  {32'hc037938e, 32'h40b217f8} /* (1, 9, 3) {real, imag} */,
  {32'h413907c9, 32'hc14fe88d} /* (1, 9, 2) {real, imag} */,
  {32'h412a184a, 32'h41516b06} /* (1, 9, 1) {real, imag} */,
  {32'h415b7c56, 32'hc109093e} /* (1, 9, 0) {real, imag} */,
  {32'h40b7e93f, 32'hc113f22b} /* (1, 8, 15) {real, imag} */,
  {32'hc0986560, 32'h40eb4342} /* (1, 8, 14) {real, imag} */,
  {32'hc02772b3, 32'hc183c2e8} /* (1, 8, 13) {real, imag} */,
  {32'hc0d67a0b, 32'hc070da36} /* (1, 8, 12) {real, imag} */,
  {32'h3fb8b778, 32'h410ee2c5} /* (1, 8, 11) {real, imag} */,
  {32'hc02d646f, 32'hbe98e984} /* (1, 8, 10) {real, imag} */,
  {32'hbea196ec, 32'h405a63b7} /* (1, 8, 9) {real, imag} */,
  {32'h40152fe4, 32'hc055db4a} /* (1, 8, 8) {real, imag} */,
  {32'h40899c52, 32'hc0554f2f} /* (1, 8, 7) {real, imag} */,
  {32'hc1000f21, 32'hc03be0bc} /* (1, 8, 6) {real, imag} */,
  {32'h3fdd5e20, 32'h407e0ecb} /* (1, 8, 5) {real, imag} */,
  {32'hc1170d1b, 32'h40e3db31} /* (1, 8, 4) {real, imag} */,
  {32'h40d21f16, 32'hc0cae288} /* (1, 8, 3) {real, imag} */,
  {32'hc109b2ff, 32'h4104a25c} /* (1, 8, 2) {real, imag} */,
  {32'hc12b8980, 32'hbf788f60} /* (1, 8, 1) {real, imag} */,
  {32'hc0ec8caa, 32'hc0135892} /* (1, 8, 0) {real, imag} */,
  {32'h40710e45, 32'h3fb2e834} /* (1, 7, 15) {real, imag} */,
  {32'hc017d7cd, 32'hc0b80b46} /* (1, 7, 14) {real, imag} */,
  {32'h40434cf6, 32'h40677f7c} /* (1, 7, 13) {real, imag} */,
  {32'h419d0e88, 32'h408397d4} /* (1, 7, 12) {real, imag} */,
  {32'h3fe5331e, 32'h3ee7b178} /* (1, 7, 11) {real, imag} */,
  {32'h40040a4e, 32'h3fc61606} /* (1, 7, 10) {real, imag} */,
  {32'hc10214ca, 32'h3f777740} /* (1, 7, 9) {real, imag} */,
  {32'hbe2a4400, 32'h3ffbc8ae} /* (1, 7, 8) {real, imag} */,
  {32'h40167188, 32'hbfbbc778} /* (1, 7, 7) {real, imag} */,
  {32'hc1105a34, 32'hc037fc9d} /* (1, 7, 6) {real, imag} */,
  {32'hc02926cd, 32'hc0073867} /* (1, 7, 5) {real, imag} */,
  {32'hc0efe391, 32'hc02737ed} /* (1, 7, 4) {real, imag} */,
  {32'h4004300a, 32'h40c493b2} /* (1, 7, 3) {real, imag} */,
  {32'hc0c15234, 32'hbf78b914} /* (1, 7, 2) {real, imag} */,
  {32'hbfec3326, 32'hc17bd892} /* (1, 7, 1) {real, imag} */,
  {32'h412746ab, 32'h406d51eb} /* (1, 7, 0) {real, imag} */,
  {32'h40321310, 32'hc0dd8b94} /* (1, 6, 15) {real, imag} */,
  {32'hc133c734, 32'h411edcac} /* (1, 6, 14) {real, imag} */,
  {32'hbfb2c140, 32'hc13dfc95} /* (1, 6, 13) {real, imag} */,
  {32'hc0303038, 32'hc14020ce} /* (1, 6, 12) {real, imag} */,
  {32'hbfbe3844, 32'hc108802f} /* (1, 6, 11) {real, imag} */,
  {32'h3fba8306, 32'h41432762} /* (1, 6, 10) {real, imag} */,
  {32'h40a33b93, 32'hc08b50a8} /* (1, 6, 9) {real, imag} */,
  {32'h404b0720, 32'hc0e2dfbf} /* (1, 6, 8) {real, imag} */,
  {32'hbf7cbfb8, 32'h40a4a02c} /* (1, 6, 7) {real, imag} */,
  {32'hbf98df76, 32'h3fd3dc08} /* (1, 6, 6) {real, imag} */,
  {32'h4179686c, 32'hbe307840} /* (1, 6, 5) {real, imag} */,
  {32'h41fd7889, 32'h405e7ffc} /* (1, 6, 4) {real, imag} */,
  {32'hc1cb6236, 32'hc0e6f712} /* (1, 6, 3) {real, imag} */,
  {32'hc160480e, 32'hbffe1518} /* (1, 6, 2) {real, imag} */,
  {32'hc1a4e2f4, 32'h40ddb6fc} /* (1, 6, 1) {real, imag} */,
  {32'h419a7d0e, 32'h3fc9fb94} /* (1, 6, 0) {real, imag} */,
  {32'hc19a74c3, 32'h3ff91268} /* (1, 5, 15) {real, imag} */,
  {32'h420b5762, 32'hc2325717} /* (1, 5, 14) {real, imag} */,
  {32'hc0a873e8, 32'h3f648c10} /* (1, 5, 13) {real, imag} */,
  {32'h3f1632e0, 32'hc0a825dd} /* (1, 5, 12) {real, imag} */,
  {32'h411725cc, 32'h419b5a1b} /* (1, 5, 11) {real, imag} */,
  {32'hc0aa0dd0, 32'h3f16d790} /* (1, 5, 10) {real, imag} */,
  {32'hc10fa538, 32'h40964b38} /* (1, 5, 9) {real, imag} */,
  {32'hc09b6035, 32'h40c1c838} /* (1, 5, 8) {real, imag} */,
  {32'h40fe0b97, 32'h410670c4} /* (1, 5, 7) {real, imag} */,
  {32'h409dea04, 32'hc0d70a52} /* (1, 5, 6) {real, imag} */,
  {32'hbfd3d910, 32'h4161ad49} /* (1, 5, 5) {real, imag} */,
  {32'hc028c110, 32'h41043e3e} /* (1, 5, 4) {real, imag} */,
  {32'hc0ca770c, 32'hc153e173} /* (1, 5, 3) {real, imag} */,
  {32'hc1bd9cac, 32'h40e6bd38} /* (1, 5, 2) {real, imag} */,
  {32'h40c6cab3, 32'hc1045cd9} /* (1, 5, 1) {real, imag} */,
  {32'hc1201ffe, 32'h424aed77} /* (1, 5, 0) {real, imag} */,
  {32'h421da145, 32'h40e6fec0} /* (1, 4, 15) {real, imag} */,
  {32'hc18c3743, 32'h41427d5a} /* (1, 4, 14) {real, imag} */,
  {32'h410e03f6, 32'hc1ae5bf1} /* (1, 4, 13) {real, imag} */,
  {32'hc1cf483e, 32'h424e5946} /* (1, 4, 12) {real, imag} */,
  {32'hc198c5f5, 32'hc0cbaa64} /* (1, 4, 11) {real, imag} */,
  {32'hc10e312f, 32'hc0f77b66} /* (1, 4, 10) {real, imag} */,
  {32'h4134ff3b, 32'hc0aeb8f8} /* (1, 4, 9) {real, imag} */,
  {32'hbfe6dc98, 32'h4105dbe4} /* (1, 4, 8) {real, imag} */,
  {32'hc0fcf496, 32'hc05cef28} /* (1, 4, 7) {real, imag} */,
  {32'h41183c35, 32'h401e6817} /* (1, 4, 6) {real, imag} */,
  {32'hc06c6196, 32'hc0bff698} /* (1, 4, 5) {real, imag} */,
  {32'hc19b0fa6, 32'h40fb8500} /* (1, 4, 4) {real, imag} */,
  {32'hc1995427, 32'h4016b050} /* (1, 4, 3) {real, imag} */,
  {32'h411f5105, 32'h40acc2a1} /* (1, 4, 2) {real, imag} */,
  {32'h41ffeef7, 32'hc1a9d639} /* (1, 4, 1) {real, imag} */,
  {32'hc0a2f81a, 32'hc1e8fbfe} /* (1, 4, 0) {real, imag} */,
  {32'hc2203f2e, 32'hc2882ec6} /* (1, 3, 15) {real, imag} */,
  {32'h41100c8e, 32'h4200dc5d} /* (1, 3, 14) {real, imag} */,
  {32'h41bd3d83, 32'h41708125} /* (1, 3, 13) {real, imag} */,
  {32'h4205918e, 32'h417412c2} /* (1, 3, 12) {real, imag} */,
  {32'hc195264b, 32'h41440528} /* (1, 3, 11) {real, imag} */,
  {32'h40972b0d, 32'hc01d1bc4} /* (1, 3, 10) {real, imag} */,
  {32'hc0f04c30, 32'h40e90f48} /* (1, 3, 9) {real, imag} */,
  {32'hc090ceda, 32'h410f48fe} /* (1, 3, 8) {real, imag} */,
  {32'hc0ab2b5c, 32'h40b38d58} /* (1, 3, 7) {real, imag} */,
  {32'hbfc7df64, 32'hc1519cc1} /* (1, 3, 6) {real, imag} */,
  {32'hc18ce007, 32'hbfc39740} /* (1, 3, 5) {real, imag} */,
  {32'hc20f2ee4, 32'hc1b1ab07} /* (1, 3, 4) {real, imag} */,
  {32'h418b5563, 32'hc171b387} /* (1, 3, 3) {real, imag} */,
  {32'h4205dd82, 32'hc106c969} /* (1, 3, 2) {real, imag} */,
  {32'hc1f1ea57, 32'h41a6bc7a} /* (1, 3, 1) {real, imag} */,
  {32'hc10b146f, 32'h41933f07} /* (1, 3, 0) {real, imag} */,
  {32'hc201914d, 32'h407be6bb} /* (1, 2, 15) {real, imag} */,
  {32'hc17944ac, 32'h415a8b99} /* (1, 2, 14) {real, imag} */,
  {32'hc136e0aa, 32'h40161803} /* (1, 2, 13) {real, imag} */,
  {32'h41e3f3e0, 32'h4113ea17} /* (1, 2, 12) {real, imag} */,
  {32'hc139382a, 32'hc1240075} /* (1, 2, 11) {real, imag} */,
  {32'h4125851b, 32'h41250502} /* (1, 2, 10) {real, imag} */,
  {32'h40917224, 32'hc109b3ee} /* (1, 2, 9) {real, imag} */,
  {32'h4147a852, 32'hbff9b1f0} /* (1, 2, 8) {real, imag} */,
  {32'hc167985a, 32'hc0e89d49} /* (1, 2, 7) {real, imag} */,
  {32'hc0943f22, 32'hc063c807} /* (1, 2, 6) {real, imag} */,
  {32'h41ae484f, 32'hc1630963} /* (1, 2, 5) {real, imag} */,
  {32'hc107ddfc, 32'h4123bafb} /* (1, 2, 4) {real, imag} */,
  {32'h4191188f, 32'h4011eb19} /* (1, 2, 3) {real, imag} */,
  {32'h428ba3f8, 32'h3ea99460} /* (1, 2, 2) {real, imag} */,
  {32'h413c106f, 32'h40197463} /* (1, 2, 1) {real, imag} */,
  {32'hc156161a, 32'hc21e0c1c} /* (1, 2, 0) {real, imag} */,
  {32'hc0f2d4e0, 32'h421cad88} /* (1, 1, 15) {real, imag} */,
  {32'h42621a70, 32'hc18e5ee4} /* (1, 1, 14) {real, imag} */,
  {32'hc0d7fd28, 32'h424bb0bf} /* (1, 1, 13) {real, imag} */,
  {32'h41208330, 32'hc12cd9e6} /* (1, 1, 12) {real, imag} */,
  {32'h3fa05c08, 32'hc1ac8992} /* (1, 1, 11) {real, imag} */,
  {32'h40e55c66, 32'hc15a1830} /* (1, 1, 10) {real, imag} */,
  {32'hc0545fe8, 32'hc128cbe4} /* (1, 1, 9) {real, imag} */,
  {32'hc01669e8, 32'hc0365bde} /* (1, 1, 8) {real, imag} */,
  {32'hc158895a, 32'hc17512b4} /* (1, 1, 7) {real, imag} */,
  {32'h413149bf, 32'h407b359a} /* (1, 1, 6) {real, imag} */,
  {32'hc1272329, 32'h41caa356} /* (1, 1, 5) {real, imag} */,
  {32'h4033b950, 32'h4195e4c9} /* (1, 1, 4) {real, imag} */,
  {32'hc2a0fdfa, 32'h411207fc} /* (1, 1, 3) {real, imag} */,
  {32'hc2623ac4, 32'hc14ed1ff} /* (1, 1, 2) {real, imag} */,
  {32'h41deba66, 32'h4050ed40} /* (1, 1, 1) {real, imag} */,
  {32'h41455dba, 32'hc100577c} /* (1, 1, 0) {real, imag} */,
  {32'h41e38c9a, 32'hc22a9b68} /* (1, 0, 15) {real, imag} */,
  {32'hc16fde50, 32'h42758245} /* (1, 0, 14) {real, imag} */,
  {32'hc113e068, 32'hc0d7266c} /* (1, 0, 13) {real, imag} */,
  {32'h42970c3f, 32'hc1e51565} /* (1, 0, 12) {real, imag} */,
  {32'h4135d946, 32'h41632ee4} /* (1, 0, 11) {real, imag} */,
  {32'hc1386e0c, 32'hc25b90c4} /* (1, 0, 10) {real, imag} */,
  {32'hc0d03b18, 32'h41d84d47} /* (1, 0, 9) {real, imag} */,
  {32'h4187f286, 32'hc0843134} /* (1, 0, 8) {real, imag} */,
  {32'hc1c3c578, 32'hbfc17ad0} /* (1, 0, 7) {real, imag} */,
  {32'h41c7b1c2, 32'hc0eba6a0} /* (1, 0, 6) {real, imag} */,
  {32'h41f888d5, 32'hc16889a8} /* (1, 0, 5) {real, imag} */,
  {32'hc141ec98, 32'h41db4057} /* (1, 0, 4) {real, imag} */,
  {32'hbf0b3660, 32'hc2819c9d} /* (1, 0, 3) {real, imag} */,
  {32'h41f6d154, 32'hc23fd0fb} /* (1, 0, 2) {real, imag} */,
  {32'h40f48020, 32'h42a95903} /* (1, 0, 1) {real, imag} */,
  {32'hc19fb956, 32'h423e8d84} /* (1, 0, 0) {real, imag} */,
  {32'h41297f60, 32'hc22235ec} /* (0, 15, 15) {real, imag} */,
  {32'hc232c64e, 32'hc1ad9693} /* (0, 15, 14) {real, imag} */,
  {32'hc13b5b8b, 32'h41882c4d} /* (0, 15, 13) {real, imag} */,
  {32'h420934fc, 32'h40e82911} /* (0, 15, 12) {real, imag} */,
  {32'h40eb4f88, 32'h413ae3f4} /* (0, 15, 11) {real, imag} */,
  {32'h41862f04, 32'h3fc23c64} /* (0, 15, 10) {real, imag} */,
  {32'hbee50e50, 32'h40c677e2} /* (0, 15, 9) {real, imag} */,
  {32'h41525cad, 32'h41727c74} /* (0, 15, 8) {real, imag} */,
  {32'hc11d7afc, 32'h41aad5b6} /* (0, 15, 7) {real, imag} */,
  {32'h41c3fe3c, 32'h41388828} /* (0, 15, 6) {real, imag} */,
  {32'h404e8498, 32'h421db8ac} /* (0, 15, 5) {real, imag} */,
  {32'h4144da57, 32'hc0bbdfd7} /* (0, 15, 4) {real, imag} */,
  {32'h412f6d21, 32'hc26b1e5a} /* (0, 15, 3) {real, imag} */,
  {32'hc1f5e15f, 32'h4155320e} /* (0, 15, 2) {real, imag} */,
  {32'hc20d3090, 32'hc13b6735} /* (0, 15, 1) {real, imag} */,
  {32'hc1eba6d6, 32'hc1c23ae6} /* (0, 15, 0) {real, imag} */,
  {32'h41c70bc6, 32'hc111012a} /* (0, 14, 15) {real, imag} */,
  {32'hc2200368, 32'hc13dda87} /* (0, 14, 14) {real, imag} */,
  {32'h3e820288, 32'hc258d124} /* (0, 14, 13) {real, imag} */,
  {32'hc19135ea, 32'hc10f617b} /* (0, 14, 12) {real, imag} */,
  {32'hc187fb6e, 32'h40bb61ff} /* (0, 14, 11) {real, imag} */,
  {32'h40e55ff8, 32'hc19dd002} /* (0, 14, 10) {real, imag} */,
  {32'h400de32a, 32'hbfab1608} /* (0, 14, 9) {real, imag} */,
  {32'hc0a15b98, 32'hbfddc460} /* (0, 14, 8) {real, imag} */,
  {32'h3f977ab4, 32'hc00dc41c} /* (0, 14, 7) {real, imag} */,
  {32'hc1b9cc2e, 32'h41bf7ca2} /* (0, 14, 6) {real, imag} */,
  {32'h40e80c8a, 32'hc1028254} /* (0, 14, 5) {real, imag} */,
  {32'hc002837c, 32'h42064476} /* (0, 14, 4) {real, imag} */,
  {32'h40455075, 32'hc1fef8e7} /* (0, 14, 3) {real, imag} */,
  {32'h421b248e, 32'hc2273eb2} /* (0, 14, 2) {real, imag} */,
  {32'hc13249d8, 32'h4207c734} /* (0, 14, 1) {real, imag} */,
  {32'hc094fd30, 32'h422ddf11} /* (0, 14, 0) {real, imag} */,
  {32'h3f485c60, 32'h40c87994} /* (0, 13, 15) {real, imag} */,
  {32'hc1580cc8, 32'h4071981c} /* (0, 13, 14) {real, imag} */,
  {32'h3fe50850, 32'hc2332228} /* (0, 13, 13) {real, imag} */,
  {32'hc06213c0, 32'h425a035e} /* (0, 13, 12) {real, imag} */,
  {32'h41dd90ea, 32'h415919e4} /* (0, 13, 11) {real, imag} */,
  {32'hc1713cd0, 32'h40be35b1} /* (0, 13, 10) {real, imag} */,
  {32'hbfc0c1d8, 32'hc09f30da} /* (0, 13, 9) {real, imag} */,
  {32'h412413b0, 32'h3fc0c8b0} /* (0, 13, 8) {real, imag} */,
  {32'h3f811170, 32'h40c65d92} /* (0, 13, 7) {real, imag} */,
  {32'hc1cd39d0, 32'hc099895b} /* (0, 13, 6) {real, imag} */,
  {32'hc137e514, 32'h42127940} /* (0, 13, 5) {real, imag} */,
  {32'h4228f6d2, 32'hc15b1dc2} /* (0, 13, 4) {real, imag} */,
  {32'hc21e85ca, 32'h40d7ce88} /* (0, 13, 3) {real, imag} */,
  {32'hc1f0d41c, 32'hbfa07cb5} /* (0, 13, 2) {real, imag} */,
  {32'hc1e0eb63, 32'hc2879253} /* (0, 13, 1) {real, imag} */,
  {32'h4231ee4a, 32'hc24f9338} /* (0, 13, 0) {real, imag} */,
  {32'h40ec4db4, 32'hc161217f} /* (0, 12, 15) {real, imag} */,
  {32'h4090edd6, 32'h41c47958} /* (0, 12, 14) {real, imag} */,
  {32'hc1dbcff3, 32'h40e95f88} /* (0, 12, 13) {real, imag} */,
  {32'hc1a49ae6, 32'h4230411c} /* (0, 12, 12) {real, imag} */,
  {32'hc181eab3, 32'h41677a1e} /* (0, 12, 11) {real, imag} */,
  {32'hc00980fc, 32'hc1e8941e} /* (0, 12, 10) {real, imag} */,
  {32'hc03d40b4, 32'h3fcdb624} /* (0, 12, 9) {real, imag} */,
  {32'h407b2194, 32'h41203c1f} /* (0, 12, 8) {real, imag} */,
  {32'hc0be59c2, 32'hc1421060} /* (0, 12, 7) {real, imag} */,
  {32'h404d2878, 32'hc08b71fa} /* (0, 12, 6) {real, imag} */,
  {32'hc07e0f86, 32'h408c3a75} /* (0, 12, 5) {real, imag} */,
  {32'hbe708140, 32'hc1f9487c} /* (0, 12, 4) {real, imag} */,
  {32'hc2071dad, 32'h4216541c} /* (0, 12, 3) {real, imag} */,
  {32'hc0f21f20, 32'hc10671a9} /* (0, 12, 2) {real, imag} */,
  {32'h42782e6c, 32'hc1a9bed8} /* (0, 12, 1) {real, imag} */,
  {32'h41b94be8, 32'h42005658} /* (0, 12, 0) {real, imag} */,
  {32'hc1976988, 32'hc12fdb30} /* (0, 11, 15) {real, imag} */,
  {32'h41790d4a, 32'h41f83ca2} /* (0, 11, 14) {real, imag} */,
  {32'h411813f4, 32'hc0ad06f6} /* (0, 11, 13) {real, imag} */,
  {32'hbfedac6c, 32'h402a6e38} /* (0, 11, 12) {real, imag} */,
  {32'h415ff988, 32'hc143a24f} /* (0, 11, 11) {real, imag} */,
  {32'h407ed78e, 32'h3fe63ecb} /* (0, 11, 10) {real, imag} */,
  {32'h4015be1e, 32'h4025e544} /* (0, 11, 9) {real, imag} */,
  {32'h412e22f6, 32'h413b5d22} /* (0, 11, 8) {real, imag} */,
  {32'hc07a823a, 32'hc0d4ab7a} /* (0, 11, 7) {real, imag} */,
  {32'h416bbad2, 32'hc060d54a} /* (0, 11, 6) {real, imag} */,
  {32'hc0acf1d9, 32'hbeb320a0} /* (0, 11, 5) {real, imag} */,
  {32'h40e3b0e7, 32'hbf731780} /* (0, 11, 4) {real, imag} */,
  {32'hc1c89970, 32'hc1f17a58} /* (0, 11, 3) {real, imag} */,
  {32'h3f16e6c8, 32'hc21adecf} /* (0, 11, 2) {real, imag} */,
  {32'h41819bf0, 32'h3d1a4a00} /* (0, 11, 1) {real, imag} */,
  {32'h41cd1ccd, 32'h41b52b4f} /* (0, 11, 0) {real, imag} */,
  {32'h4191cecc, 32'h40b6264c} /* (0, 10, 15) {real, imag} */,
  {32'h417b78dd, 32'hc1830987} /* (0, 10, 14) {real, imag} */,
  {32'h40deb443, 32'h4152b367} /* (0, 10, 13) {real, imag} */,
  {32'hc144c8fd, 32'h415482dc} /* (0, 10, 12) {real, imag} */,
  {32'hc111f362, 32'h3e892b44} /* (0, 10, 11) {real, imag} */,
  {32'h401fa007, 32'h41103e90} /* (0, 10, 10) {real, imag} */,
  {32'h3fbc551c, 32'hc049f4b9} /* (0, 10, 9) {real, imag} */,
  {32'h3da87a80, 32'hc1363aca} /* (0, 10, 8) {real, imag} */,
  {32'h4096d7bb, 32'h40cd72b4} /* (0, 10, 7) {real, imag} */,
  {32'h40a2052a, 32'h408e44eb} /* (0, 10, 6) {real, imag} */,
  {32'hc10b08e8, 32'hc05cdbf8} /* (0, 10, 5) {real, imag} */,
  {32'h41137883, 32'h41485928} /* (0, 10, 4) {real, imag} */,
  {32'hc0d1211f, 32'h415514b5} /* (0, 10, 3) {real, imag} */,
  {32'h40695dac, 32'h4131ace1} /* (0, 10, 2) {real, imag} */,
  {32'hc1eabc14, 32'hc0e4f0c4} /* (0, 10, 1) {real, imag} */,
  {32'h41b0b9f2, 32'h3f981cec} /* (0, 10, 0) {real, imag} */,
  {32'h4190c361, 32'h41ab9be4} /* (0, 9, 15) {real, imag} */,
  {32'hc0ff1ca5, 32'h408e2baf} /* (0, 9, 14) {real, imag} */,
  {32'hc158400a, 32'h3fbe1880} /* (0, 9, 13) {real, imag} */,
  {32'h3f2c54f2, 32'hc129a16a} /* (0, 9, 12) {real, imag} */,
  {32'h3de92a40, 32'h3ff70e14} /* (0, 9, 11) {real, imag} */,
  {32'h4081a4c1, 32'hbfca3a02} /* (0, 9, 10) {real, imag} */,
  {32'h4009807f, 32'h402581eb} /* (0, 9, 9) {real, imag} */,
  {32'h3e8fcf64, 32'hbf93f004} /* (0, 9, 8) {real, imag} */,
  {32'hc008ba97, 32'h3fe2e466} /* (0, 9, 7) {real, imag} */,
  {32'h40b627b9, 32'h402952af} /* (0, 9, 6) {real, imag} */,
  {32'hc103c812, 32'hc09a5af9} /* (0, 9, 5) {real, imag} */,
  {32'h403856da, 32'h40d15961} /* (0, 9, 4) {real, imag} */,
  {32'hbf593a88, 32'hc17e3998} /* (0, 9, 3) {real, imag} */,
  {32'h40f44107, 32'hc03b592a} /* (0, 9, 2) {real, imag} */,
  {32'h4170cdf6, 32'hc0bca886} /* (0, 9, 1) {real, imag} */,
  {32'h4067ede4, 32'h3ff75bd0} /* (0, 9, 0) {real, imag} */,
  {32'h3ffcc758, 32'hbf940754} /* (0, 8, 15) {real, imag} */,
  {32'hbfc3c87d, 32'hc1a67bee} /* (0, 8, 14) {real, imag} */,
  {32'h40f97048, 32'hc1263abc} /* (0, 8, 13) {real, imag} */,
  {32'h41288aa2, 32'hbf9fb51c} /* (0, 8, 12) {real, imag} */,
  {32'h3f3509a4, 32'h3fb40dc0} /* (0, 8, 11) {real, imag} */,
  {32'hc003bd30, 32'h3eb606a0} /* (0, 8, 10) {real, imag} */,
  {32'hc017e476, 32'h3fa0edfc} /* (0, 8, 9) {real, imag} */,
  {32'hbe952e40, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hc017e476, 32'hbfa0edfc} /* (0, 8, 7) {real, imag} */,
  {32'hc003bd30, 32'hbeb606a0} /* (0, 8, 6) {real, imag} */,
  {32'h3f3509a4, 32'hbfb40dc0} /* (0, 8, 5) {real, imag} */,
  {32'h41288aa2, 32'h3f9fb51c} /* (0, 8, 4) {real, imag} */,
  {32'h40f97048, 32'h41263abc} /* (0, 8, 3) {real, imag} */,
  {32'hbfc3c87d, 32'h41a67bee} /* (0, 8, 2) {real, imag} */,
  {32'h3ffcc758, 32'h3f940754} /* (0, 8, 1) {real, imag} */,
  {32'hc1d36629, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h4170cdf6, 32'h40bca886} /* (0, 7, 15) {real, imag} */,
  {32'h40f44107, 32'h403b592a} /* (0, 7, 14) {real, imag} */,
  {32'hbf593a88, 32'h417e3998} /* (0, 7, 13) {real, imag} */,
  {32'h403856da, 32'hc0d15961} /* (0, 7, 12) {real, imag} */,
  {32'hc103c812, 32'h409a5af9} /* (0, 7, 11) {real, imag} */,
  {32'h40b627b9, 32'hc02952af} /* (0, 7, 10) {real, imag} */,
  {32'hc008ba97, 32'hbfe2e466} /* (0, 7, 9) {real, imag} */,
  {32'h3e8fcf64, 32'h3f93f004} /* (0, 7, 8) {real, imag} */,
  {32'h4009807f, 32'hc02581eb} /* (0, 7, 7) {real, imag} */,
  {32'h4081a4c1, 32'h3fca3a02} /* (0, 7, 6) {real, imag} */,
  {32'h3de92a40, 32'hbff70e14} /* (0, 7, 5) {real, imag} */,
  {32'h3f2c54f2, 32'h4129a16a} /* (0, 7, 4) {real, imag} */,
  {32'hc158400a, 32'hbfbe1880} /* (0, 7, 3) {real, imag} */,
  {32'hc0ff1ca5, 32'hc08e2baf} /* (0, 7, 2) {real, imag} */,
  {32'h4190c361, 32'hc1ab9be4} /* (0, 7, 1) {real, imag} */,
  {32'h4067ede4, 32'hbff75bd0} /* (0, 7, 0) {real, imag} */,
  {32'hc1eabc14, 32'h40e4f0c4} /* (0, 6, 15) {real, imag} */,
  {32'h40695dac, 32'hc131ace1} /* (0, 6, 14) {real, imag} */,
  {32'hc0d1211f, 32'hc15514b5} /* (0, 6, 13) {real, imag} */,
  {32'h41137883, 32'hc1485928} /* (0, 6, 12) {real, imag} */,
  {32'hc10b08e8, 32'h405cdbf8} /* (0, 6, 11) {real, imag} */,
  {32'h40a2052a, 32'hc08e44eb} /* (0, 6, 10) {real, imag} */,
  {32'h4096d7bb, 32'hc0cd72b4} /* (0, 6, 9) {real, imag} */,
  {32'h3da87a80, 32'h41363aca} /* (0, 6, 8) {real, imag} */,
  {32'h3fbc551c, 32'h4049f4b9} /* (0, 6, 7) {real, imag} */,
  {32'h401fa007, 32'hc1103e90} /* (0, 6, 6) {real, imag} */,
  {32'hc111f362, 32'hbe892b44} /* (0, 6, 5) {real, imag} */,
  {32'hc144c8fd, 32'hc15482dc} /* (0, 6, 4) {real, imag} */,
  {32'h40deb443, 32'hc152b367} /* (0, 6, 3) {real, imag} */,
  {32'h417b78dd, 32'h41830987} /* (0, 6, 2) {real, imag} */,
  {32'h4191cecc, 32'hc0b6264c} /* (0, 6, 1) {real, imag} */,
  {32'h41b0b9f2, 32'hbf981cec} /* (0, 6, 0) {real, imag} */,
  {32'h41819bf0, 32'hbd1a4a00} /* (0, 5, 15) {real, imag} */,
  {32'h3f16e6c8, 32'h421adecf} /* (0, 5, 14) {real, imag} */,
  {32'hc1c89970, 32'h41f17a58} /* (0, 5, 13) {real, imag} */,
  {32'h40e3b0e7, 32'h3f731780} /* (0, 5, 12) {real, imag} */,
  {32'hc0acf1d9, 32'h3eb320a0} /* (0, 5, 11) {real, imag} */,
  {32'h416bbad2, 32'h4060d54a} /* (0, 5, 10) {real, imag} */,
  {32'hc07a823a, 32'h40d4ab7a} /* (0, 5, 9) {real, imag} */,
  {32'h412e22f6, 32'hc13b5d22} /* (0, 5, 8) {real, imag} */,
  {32'h4015be1e, 32'hc025e544} /* (0, 5, 7) {real, imag} */,
  {32'h407ed78e, 32'hbfe63ecb} /* (0, 5, 6) {real, imag} */,
  {32'h415ff988, 32'h4143a24f} /* (0, 5, 5) {real, imag} */,
  {32'hbfedac6c, 32'hc02a6e38} /* (0, 5, 4) {real, imag} */,
  {32'h411813f4, 32'h40ad06f6} /* (0, 5, 3) {real, imag} */,
  {32'h41790d4a, 32'hc1f83ca2} /* (0, 5, 2) {real, imag} */,
  {32'hc1976988, 32'h412fdb30} /* (0, 5, 1) {real, imag} */,
  {32'h41cd1ccd, 32'hc1b52b4f} /* (0, 5, 0) {real, imag} */,
  {32'h42782e6c, 32'h41a9bed8} /* (0, 4, 15) {real, imag} */,
  {32'hc0f21f20, 32'h410671a9} /* (0, 4, 14) {real, imag} */,
  {32'hc2071dad, 32'hc216541c} /* (0, 4, 13) {real, imag} */,
  {32'hbe708140, 32'h41f9487c} /* (0, 4, 12) {real, imag} */,
  {32'hc07e0f86, 32'hc08c3a75} /* (0, 4, 11) {real, imag} */,
  {32'h404d2878, 32'h408b71fa} /* (0, 4, 10) {real, imag} */,
  {32'hc0be59c2, 32'h41421060} /* (0, 4, 9) {real, imag} */,
  {32'h407b2194, 32'hc1203c1f} /* (0, 4, 8) {real, imag} */,
  {32'hc03d40b4, 32'hbfcdb624} /* (0, 4, 7) {real, imag} */,
  {32'hc00980fc, 32'h41e8941e} /* (0, 4, 6) {real, imag} */,
  {32'hc181eab3, 32'hc1677a1e} /* (0, 4, 5) {real, imag} */,
  {32'hc1a49ae6, 32'hc230411c} /* (0, 4, 4) {real, imag} */,
  {32'hc1dbcff3, 32'hc0e95f88} /* (0, 4, 3) {real, imag} */,
  {32'h4090edd6, 32'hc1c47958} /* (0, 4, 2) {real, imag} */,
  {32'h40ec4db4, 32'h4161217f} /* (0, 4, 1) {real, imag} */,
  {32'h41b94be8, 32'hc2005658} /* (0, 4, 0) {real, imag} */,
  {32'hc1e0eb63, 32'h42879253} /* (0, 3, 15) {real, imag} */,
  {32'hc1f0d41c, 32'h3fa07cb5} /* (0, 3, 14) {real, imag} */,
  {32'hc21e85ca, 32'hc0d7ce88} /* (0, 3, 13) {real, imag} */,
  {32'h4228f6d2, 32'h415b1dc2} /* (0, 3, 12) {real, imag} */,
  {32'hc137e514, 32'hc2127940} /* (0, 3, 11) {real, imag} */,
  {32'hc1cd39d0, 32'h4099895b} /* (0, 3, 10) {real, imag} */,
  {32'h3f811170, 32'hc0c65d92} /* (0, 3, 9) {real, imag} */,
  {32'h412413b0, 32'hbfc0c8b0} /* (0, 3, 8) {real, imag} */,
  {32'hbfc0c1d8, 32'h409f30da} /* (0, 3, 7) {real, imag} */,
  {32'hc1713cd0, 32'hc0be35b1} /* (0, 3, 6) {real, imag} */,
  {32'h41dd90ea, 32'hc15919e4} /* (0, 3, 5) {real, imag} */,
  {32'hc06213c0, 32'hc25a035e} /* (0, 3, 4) {real, imag} */,
  {32'h3fe50850, 32'h42332228} /* (0, 3, 3) {real, imag} */,
  {32'hc1580cc8, 32'hc071981c} /* (0, 3, 2) {real, imag} */,
  {32'h3f485c60, 32'hc0c87994} /* (0, 3, 1) {real, imag} */,
  {32'h4231ee4a, 32'h424f9338} /* (0, 3, 0) {real, imag} */,
  {32'hc13249d8, 32'hc207c734} /* (0, 2, 15) {real, imag} */,
  {32'h421b248e, 32'h42273eb2} /* (0, 2, 14) {real, imag} */,
  {32'h40455075, 32'h41fef8e7} /* (0, 2, 13) {real, imag} */,
  {32'hc002837c, 32'hc2064476} /* (0, 2, 12) {real, imag} */,
  {32'h40e80c8a, 32'h41028254} /* (0, 2, 11) {real, imag} */,
  {32'hc1b9cc2e, 32'hc1bf7ca2} /* (0, 2, 10) {real, imag} */,
  {32'h3f977ab4, 32'h400dc41c} /* (0, 2, 9) {real, imag} */,
  {32'hc0a15b98, 32'h3fddc460} /* (0, 2, 8) {real, imag} */,
  {32'h400de32a, 32'h3fab1608} /* (0, 2, 7) {real, imag} */,
  {32'h40e55ff8, 32'h419dd002} /* (0, 2, 6) {real, imag} */,
  {32'hc187fb6e, 32'hc0bb61ff} /* (0, 2, 5) {real, imag} */,
  {32'hc19135ea, 32'h410f617b} /* (0, 2, 4) {real, imag} */,
  {32'h3e820288, 32'h4258d124} /* (0, 2, 3) {real, imag} */,
  {32'hc2200368, 32'h413dda87} /* (0, 2, 2) {real, imag} */,
  {32'h41c70bc6, 32'h4111012a} /* (0, 2, 1) {real, imag} */,
  {32'hc094fd30, 32'hc22ddf11} /* (0, 2, 0) {real, imag} */,
  {32'hc20d3090, 32'h413b6735} /* (0, 1, 15) {real, imag} */,
  {32'hc1f5e15f, 32'hc155320e} /* (0, 1, 14) {real, imag} */,
  {32'h412f6d21, 32'h426b1e5a} /* (0, 1, 13) {real, imag} */,
  {32'h4144da57, 32'h40bbdfd7} /* (0, 1, 12) {real, imag} */,
  {32'h404e8498, 32'hc21db8ac} /* (0, 1, 11) {real, imag} */,
  {32'h41c3fe3c, 32'hc1388828} /* (0, 1, 10) {real, imag} */,
  {32'hc11d7afc, 32'hc1aad5b6} /* (0, 1, 9) {real, imag} */,
  {32'h41525cad, 32'hc1727c74} /* (0, 1, 8) {real, imag} */,
  {32'hbee50e50, 32'hc0c677e2} /* (0, 1, 7) {real, imag} */,
  {32'h41862f04, 32'hbfc23c64} /* (0, 1, 6) {real, imag} */,
  {32'h40eb4f88, 32'hc13ae3f4} /* (0, 1, 5) {real, imag} */,
  {32'h420934fc, 32'hc0e82911} /* (0, 1, 4) {real, imag} */,
  {32'hc13b5b8b, 32'hc1882c4d} /* (0, 1, 3) {real, imag} */,
  {32'hc232c64e, 32'h41ad9693} /* (0, 1, 2) {real, imag} */,
  {32'h41297f60, 32'h422235ec} /* (0, 1, 1) {real, imag} */,
  {32'hc1eba6d6, 32'h41c23ae6} /* (0, 1, 0) {real, imag} */,
  {32'hc144dcba, 32'hc0b10114} /* (0, 0, 15) {real, imag} */,
  {32'h414bf09c, 32'hc253b2e0} /* (0, 0, 14) {real, imag} */,
  {32'h42721bcd, 32'h412763e8} /* (0, 0, 13) {real, imag} */,
  {32'h4275e5d2, 32'hc15e4e4a} /* (0, 0, 12) {real, imag} */,
  {32'h4209ea07, 32'h41662474} /* (0, 0, 11) {real, imag} */,
  {32'hc120481e, 32'h423cb140} /* (0, 0, 10) {real, imag} */,
  {32'h41ac2355, 32'hc0f43234} /* (0, 0, 9) {real, imag} */,
  {32'hc1ff3c15, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h41ac2355, 32'h40f43234} /* (0, 0, 7) {real, imag} */,
  {32'hc120481e, 32'hc23cb140} /* (0, 0, 6) {real, imag} */,
  {32'h4209ea07, 32'hc1662474} /* (0, 0, 5) {real, imag} */,
  {32'h4275e5d2, 32'h415e4e4a} /* (0, 0, 4) {real, imag} */,
  {32'h42721bcd, 32'hc12763e8} /* (0, 0, 3) {real, imag} */,
  {32'h414bf09c, 32'h4253b2e0} /* (0, 0, 2) {real, imag} */,
  {32'hc144dcba, 32'h40b10114} /* (0, 0, 1) {real, imag} */,
  {32'hb6c00000, 32'h00000000} /* (0, 0, 0) {real, imag} */};
