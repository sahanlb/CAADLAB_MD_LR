-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
B4huNYGThBgeBGYXx0Y+6F1KFUP6RCyVxCyCUOzQnevM0K5IUvY9v+8bzBe60zI5
Nfs4+JWDG4vYykSg/VajaKSSoBUgSgQ7X76qUf0IVQGJdtg97Oz4WGdv6Btcu2X/
o0LKVxwLNjwz6VyH64CtkEZG8ncHajlTlv+FzYLq/CM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7685)

`protect DATA_BLOCK
0l4eXpPkEC1SNKVcqyaT6VroV4G4pNRGdBT3MRmYQfekTV6eX7QJW+PqwQ+fK5MS
JodLvoayyB5huCqHNdQghfECiVCovtZM/4Zb/rH1J8B9r8RcXv52m1ABr6gG4iLU
S87iPVItt6zGELzRzWud8Yps1QF+EhmHnt91V+XP/o0voQFYVnLZ60yRf8mZBvmN
8fxwDXj7h4WxbBK/hTJLSf2FMhmHPxx9xgLFJkw9cIroUt7CfrCY9Rj7Ypeyn+BE
5ygO8/4rHa1sFyqt/3O+a7fMZaOTEShbeHmzvQH/D71Oj9aG50Npw7qCVkTSUdru
V45llg1VL02obGwu2QN4/Y8FHDoi/2hg4PsYaqkT37WGahwgHbjEZRwsZgFjKcTv
EyibJxa6tmM7UuBGZnCe+8Pvu2+D33PNSfnntkn71cl1aXkAfFU0Fj3kCDRdwzAH
pIaqOdKKrTsKssFgfG0fr3HnptGL1QGetZ4JaT6rpaRJ6308eAbfsrp256EbDYkB
OHWzNqSdO5C/1tfivb4nZoEl5z10IKmPE8LH2zVGubQQ1dwVFf7ozflHj4FQ6OqB
CUs2rfb63+R5paETzW9kAeBh+UCrNaQWLpybdjVLYzti7dwZgMdfWAvj8VxJK/9F
P6Ig2R18Dc2Ymiu+M/ZuFdaNsB5DczbEOEUBztqXGpt3EzDsgBOCwcmSm8/8u1Im
Hyj6cm2SKq1dNFQMCzsCwLLJOLf7/1e5RFiqSJRUmjWnQVJskqsG+T3lsvydHtDF
mNOFlTgDu0/un74uENg14GwzH0VAXn1yAx/1Vg8zR/oYe7fZpquEON+Ejj32vvpj
DKhLZJkQd8eB/9sGySLsdp3HVfyYEkN6i7IKYi485IEr2gnel+oXvHVGEa2NOL4q
fK0k5FzOtwD4O+O7i4u0UxNZGL+eAQARkuQKiKD6N2HUzyS0gESLvAm5tS2L5rOG
heBLphc5SJTu/w/2Y660LfHHro+CmTuVaGoowzWuW4CFt/BXLeQL4DGo86UQ8bqT
fFadoT7zFgxzCBUL/sSX7mdVJf3genuOwo+CJDn5UFPKJkmWpmMZvytMoVFMj9Gu
Dmv5jnmDxCrUAuEFYk5rEhgVHWkAN0zX6Mr2sE+7go0Y9YKvD/xgNwCaCFzcs0Fq
F76ymF8JQ0QQeie6b2UQPxyXcSU48EMQdhV+ggRnslYM9x1VTJyvpk47lNcz8at8
v7cgkXAkdW4h6mP5UwgJjA2rFpoKN/leJb13vm6lpMdkU8t2FZVbTY5531hbXgTE
AVIQGoHE6aL5C/jRQtk5FywGjFCHHtO3eV0gdhyBOTUZEyumRlIftGB1YoLMnLbT
E1KevKQGVXvYHP9cSqc3mqaTiVT9r+kVoXTHdy9xfEYCYzjwiyNr7DocGzXwxPxf
osChqp4QCDFdYIeTtkdDy/NB2tzGJWOGaxz28Ni7lhP/SMseWotAv1ftPWFJRtnb
M0iMBFi5euOx0W09Ves5n1qCCmgoyKmr7Vfganyd/h7kaRSCCnFBPE7nV1BnFHV4
pRJdTVTowP6aJDCgq+FtyLQ1jU3o7oXBqLGHtzzBLePyY2scs/QvECsdTDOxrFyB
ELOecEPPrU7EqJQPedAEAJAOxLcuA656OgnHaMkaUc9sT+tG9yYW77erBlPx8edM
jF4Fu2KTzqLCxkWTQHR6hHHDNI46luD3tWjZaPhqFq3E1MF3Zg00rGnnbO82cRo3
l2Smi0C1QMAwOF4J3d1glfUS4Iq5UVzcRn7hiGTutDZd35Ms7dNHIxTiV8R/+0lv
em4zehIdU3MwvXJ+SDPNGjJZ5jL6WldwDEXi+J9eUNr0VrpOiE5JqExwi1naRGH7
ekbj+zPN8Nbs0Qq9MopniZzDHxD0NGCOmRyvVM8X3SYO5YHW9Z6+7Sv570zb1Vc4
DCyB5QQjzcSMG3Uv5RXL1Wyz2ncsD2dhF3kKVruLAYCe3JEeH11MFgvhPLW1uEvU
oLPy1/ya2Fr7G92sajUH9riJSMxGRIpqqKIhHuaYerBc4dy9zb8fPyhWg7JCvua2
OMxOqPL9MgTGbqFdqdNAveb6gY2eaEtTS2XBev5eACicnVO6hryg8/daxdiNeS/p
K4A8i+Y0Oer8BDcdY33BcFwDe6ioKyoN5Ywirt3OD4+ZXleNqRVeviXMy9BIlHim
NUsCatcUF1wOdVYja74t2BO+IBxtjGsB2/Aj8vCeBMh4Z6StxPmKg4SJsBTk3jbl
bIiJOde4m8omOSoDGyYSOQkKwG4g81msbTsunOd7Ma0i1AxuzuitIN8pyofuav7L
uWKGLiqJEkEWVTwV79YbHRyrDNMneLqbcvXfDi+Ht1feu4Y4tehIdOhHdSA9IJRX
Xl8DwfyoN7ba82i+3ErVe6G5wosed8SFzdtRSVSFKzo0hCBJY20dyS+nXWLISGBV
RIhl3bXgmIcNINZHjitCutFtqphgAulsAg3xsYB8DXQRUbBwvNIg2K5Hq6WYJFkT
xXHGUGV5GCq7/W16YccShKbK/kCDWPkEySOnNIuedaugN2vLGNltbT5wEN95AkQS
ce6EG1RWWDEDLHP6X/H6fgpqx7PV9QMMgXjZWcTwqI8HqURNA6kE93w+iW8vNUFS
Ed/EgKUTh45WzipHN/RrA1hU2io+LqgqWpNebLr5dh97ZP7YfDT2VDMKftlDYsCB
jE6P0O0KwCszMScYXINFS5HA9jtKK7mylBqwzJ5JXibxYaV6rJXGIevkDZX+U8Vg
zg8jDkD/68uYzpaJ8r0XKzDBcT9mluRxGqy/VJgIIwwYAKKNflDpNhG0xEVumKMv
eaZaSKeshvYRWcZtddi3gkC2UOgMO86H9hoi+wKlkNyBEkDNYUBlS6njXBj7q45S
A6K8iyfNfAmOITiaLGOGNgMujd/WRbK+ylZHghefD7nhKBkqAwR/2OH3u5t5KpKd
WCGfi3u1cknMPBTKUXxr2RYaCidfEc+W6k7RNVvggIx+IlB9o1WvdfO5xQeg9Ekr
1SM839OX+no0G+eq4UfqeErk98iOcqNejElZPkoeXaaaOZgiLR5Rm6sB/w1xGw+1
0icv7U/MB+qLEB7RpX+3LG6jpi0/GCxBWD7HAME45LBt5h/e0Kr36HGq3kDFXIWA
3HszCYHeeaTpj0J5zmh7/Zgi6izEXC0hWaY/6xjJQLeoOA4tDFDp2ygamGfNs+lV
uKs30hmCXlEYoCplbN664G9knq77Myztf1bbNude0e7rKDWU6FHmp64e7pqbRW6B
mQk44AgcbBugQSy+t1YaadrBDQ5CK9x+RshDzJukqTdPxMt527R0qtz7mtK8LWEB
lcRiBDMJ1CrEhlDeag1mke59g2SFF9Iwdxb49GRP3HW2JyuL0/RPgAdPnCVxR8Zw
iZOU5mDa3thBsQRqB1MRjYgYXcbAWDvg6Rh0CRYddRRKVe9ABlHRY3+KP1LgFLDo
KyoqYHU0AQaXzCyg6AMQ7IPf2MEHyp7+f0F9iDT6sTNeRaCnrQq6kCNXCy/gNy8r
bN4B8BO7ng+xYxBFLnwcILvn7I85Pe2Mp/fuuarjeU2Y2h1ODRRDKfkVTEv3Z3nc
3JLBN2giqCw6SQnql7YOJeZVdgYft9WmeqyYG60lg/mwQT/Y6wXuXiMmPW+FNpCN
FjgkNdFQSI0ZsbLJLwVU8b+UPI38bPdAINq3mB+nW1W8IFZ03/UJWqdXCd8YrD+O
AV8hrOJoTphuHb30jPITwdTnMhwPnYG+2jl3Z/YsCT8TnLyOupuFhHFnUsRTrfe0
9jUZQImzTBERj/zb6qfyXOQ22o8noKIRxjreG5s55L4I8yWfRwVrXVnci9qihKTD
5OvlFhEsE4L7PzMhVXgJIwUd2R3AnOauETS4gCKIj2LULHehj58Ze0X1//Zj1WIZ
NmjXNkQ2k00NgVtlJFgGqGZfp5JOpOB22obdfCGxV41uGMmkV9/k9aj3dTcxEQXn
mIGhXF9jrOrBcA26wBQ9Bg2iUISAMTccFUcWGpBpenGPE3S9dCAcYEogVtWxvO/s
0mJO1DVmOmBQ/UDWT1aRdId1JazbN/iUeuGPNGCYjncjDd8Z63+Bq/klYdni8EJm
rv8pvOw9dL6SINg8X1WHVtOXyFNzBVw8SDCmSeMs6T0FyV4eJThT+043eAE4iQ0m
6OH1j/atvXtnFYqaCw9XreQv20bKyf9pQWjKRQZsgrckj/51AdiIQEMVPESSitnh
0lX0mdzPCuMPfS0rkFh2b7elK26YlLLGfF+5iOh4aZaX1HnRP7OOVp8rMnViXxrN
nKYtc23f+PSjVPan66KhvRLt+Ax1S5nJH3X9fdQ+Njc2aufLy/TLR7pQ/AapMT5h
zP8N8rVejhM5i2jEgddDR9F8onoNZI+jkUi/YlhWpftNF4DOJyaxZJoj/DiOy1mW
vRoZNJAEpfFAdTfl9QoXVeGQZNHSIDH5E8bEz2V3EU/jjAaX5jjXOEH/pE2xoQGq
fJqHhkNKtRqfB0tEPDXwN17jYYBsaxwOwBK/e/2RF+2duST/EoEE4uRp/Cp0L7mV
QanwMP4pRkMrB5UPPERY2dWR7PTCn4gD9Ip48n9/0CpkTui3cnTZIsRwVUIjt4Ft
zi1wIz/8kWPtvxrbX7w8W5r+FWQ6gC+d004ed8xAepY6GjvZIN1S4suAbI941ctx
yqkwCQeWHmI+lp+XvQTYfL182r+DLqZ5ZksVpyRwWXZ4AsgWefPb9nXOGiLyvcaO
aCq4Mnmo5DXcQFAKvIg4eJMBjEzo0VzXHA/CaKCj3rXAv/UXRLUwv7C3+hea3UEP
d/15lDXT+1CiZaOnVgb6ZVEBmHPhrgrwF8vk6iwzAgTNtVnyFy97nrKZOhjW3ncf
wF3MXQNFuI7xI/7A4+uYcyoz1coQv6KX/Kw7jzpdzyTqa13IMQI/BnmAavh0IQm4
lj2DL0a19QWCT8sYh63Z3oRC2+0J/KDpqhuzIxELUyuMPRwymG4ZhZaqAQAqACq8
2C9jGYdDL+KZQ+7My0bCGv6Xfp/fhvvWAaadaCU6AsovG1Ceb0UY5RJhN0sCZDKr
wMHJSQTgwEDg093SjvNxvcsbhLmxUfoEY+p9LG59ajBPirO5bPRnRG7Vk6OjRrFe
xv631/PTvrJEAOsKxsPEKtkqnW790zaLbd7vaCuoKYuuop3OqznZNKk2v3AEGCQF
9XmwYsF2+G32jmub9F6K/mI129eOAmSqhQOsGDO33ZcebfZqRGAQJ9GDutk3oZpZ
biR8YarulN8EL/IPQLsB6tmF05v5WujxPyv/BsJcrKp++ZGE8pPL/F9PFUjbF63p
uRg/qrvr16J3L2ypAnTc+yCHmBRCchBh+Ji/SjhVoQ7xY/kE1TtZQF3jYaNY1qKf
+G01qs7hfgkAau2p+mio8OjhxXL1mcBV4X2fv/z4bWzxEj509MSn7BZArmFTiaCs
sw7n2r/zKUDXzZqNywWcxhcTER13eR+Uh4JpRSfD7OrvmYLyXzjwq8jh1Pz+Li/I
8OVKqt+P1d9+z+DWEljU1ercstUCw8+p6YdOGpnu9x57bQtb0AEKb7sMOqO61pfc
L3BRpMc+Dcko+I6YQmwney3e0LfhLVOWPvZ74NA4Fo9SbB8cFP+LpGXwzfltZ2pV
1pOiVJpcEuxKvIWIPlEo19rhLOKd2ownjJ66clQ1F+IpjpRGd3j70x6semFBfSR1
tNEeDD+MrdUBvTEsm95jm6mmFRm0ucf44BFbjLImOaDRTHXP0PqEpKz30SF5X5fz
AkTbjrCNKDqYnczI093ibs+JKZuJtsApAPdopymGU6V7jRn45CogixoenFPFBAvh
grzMR1TCINu0LgzoInOkqyEgX5ZAnI5pTtCKAknC+genk9f9E82KyP0P1NKiBw7I
j1k3r++XZdoY9LojWYQlZGttSXmBrxYjTdBkx8d46ztrzvycrenmRvogMvvnQboi
QlDcDL6Z/1YCByAJhhgWsWA2VCAhbWcDMRXnNoNOxYHGJ5iHEnKDFJT3uUjBcBLO
u/SQraORTxmsNo3DLkBmsiyQyUIF3GsiZSUWVzMKuCpX6MZaDWhOErnDtlW29RnU
kgnayV+4c+Zt9l98bhC95+rac+MgkjXcLSuiKSGHxp96feIZa58y7i5C6MhA49Kq
/JsKD5OUTMbZGg0a3rC9w9Ho9LLD0he1SJAXbhCJqthjA88VjqYYe09knHLMGeDa
cPEoMHUW3/v0bOX7F2btI8mo43CL8/3MzxB7imHkLd2A0A0XIBkqaT4rlkXwKS95
5w75ntIQtcNi8AtL/HVlI+GWek2k2CkAx3ok7w9ZOmJH2Fk6doFFeMmm4C6owmaj
SG6cgVOlpSdwF+H1av5axhbBVgQ4n57kBPqua5/1IOyojot3tSicFBT4F4Ky/ThH
wP6FgdHjvqahIo0Tk+c4NX+Mt7KGu5vOtk33F72BAbPltLO09GDDElyhqb7KFeeY
PPedBqNsfP6GNFC9tWV+7ubfv1/Hi5SHUTV/+/0DX03DIswZ9Qk8Z1cxLEmNBgB0
1jTzXg4mSa/K38oOzs1akPnkImYHkxH8OKDgZmvU/Am/G1qhNam3htsC3cADivW7
0aLB5xt4g71pg40lZrV8zMVWwCqgDigKWCHkveyewcUHZ02sUU2lO9H02/9DbtI4
GaXvmrT1SRN/vm22PlLaPT17jDlOscCHikH8l0PMboyBi+VcJcNxz0TXhIazhEiR
fVAN0ICvtFnQLPekhRb6K0tcHWub50vH+kIpch49zNP1+88vkr5pAKi/BaGUx8ke
NWk3FIKU53zWf/3wMDvEKZU51IuHthcfPdRMsh80oeYmcL0HtK+ZJ5Whzjplbu7b
Qc/B7Aoqr5o+PONX6WCABUkzoX3Vb0b+lmpXNeoCKDqpDyrDlfyrYOkp+BUhW25p
Pih1Wgi3rK6rBssRu54yk2SmJg5j74OgKLL1GwuKD0BM8bessemUFGmjlgS2hn5t
zf6sqBu6ag2S37OBCkS0jGB/lHKJ56O3wvlh8hGdaETIV+eurRRMnCfmDFYAI/Mx
0hgn64McLuTS2WK6VxwlAMWET7KxGBl1SVP78n3mrKGFemuE24r28owdN/opRx6t
/4YCVGi4b1vDOcPRAnUfMj7E2oXQYOea0S/6MDoUdAPiZwdXoFDRjyyOqAv+h3OW
TDggA1oQeJwZs2+kmeorBcnzJ0e/oOi+wR7iMOsnUFK1Wu3t2FqSY04AaXCAdB81
CntZ770htRnptU94VqTANn2uoFvvONWl/6y8zoMqK+LjeSZoxGGk7Snh9knxoYsd
0lp9DvljZpNuQ0XLDGWjQxDv+bMc6wcB2Fe1l3ltwHw5Ig74PEBbf/4VgwwF2RUE
bYAplXsgBS2wOG0nIIHeOYk+8+smQx00W4eWeTvvp+cm3ItZYXqX+Hj+dCcvNCjX
5V2Vlr5i/RQa0R/Z6WsymfVHXNcLudwn+wDnE40RC7pdp/7/o8YrQ5eO0uKPgte1
fZmYqcGhybqrl1wNhqnADDEtT+soozFw/XXn6OU7NLsf9qju27QF9YIi32kQBLBh
kSeg9EuxXCki1+kefr2gQLqoG0N5+iv/1cGFEQB+tTxKkkJ9ZRYbN0HTQzTA33jC
Vvb6WIGBVDichHtlHKNw9hGRyVvZrQiHFgTwetadmYqqtuSRJeflzR4ul4BXqm0k
PqetUdxImaoRYsOXI4MksNfz3T9rpEQ4pdXHN6eFP15+ZvLWlSPHc5qA6hE98/49
npop2A2Shn7GhSUxE7GLwiZN8bPkd8CpwkYgppEpEtXllJ1EKu/TxMSNSKq3S6CZ
K8VboGKUHAQk2dmlUo4FFqOSPZtzpw5vCSguzcyLE7Azwxo4HrYPMqkcDSlL+SZF
/JikPaPYYFjkjuO4xqhoUEDUtBjRWIv9WzVnBPWfEMl/NnPRqNVeQQR6AQmuegUm
Qx43H0XwsPbUU3A7X0npmSkIWpnNCQ5MuvkPapFEtJzpqaDyn48eCTALoIF2iIjn
ypmRNDF9k8kVcrJRCz8cdYDfz2xNeYJRIZaVwrwf8TSltJWH5JyhSzRLLNwKqW+F
RWnvEqJJDyJx0Ay5is5jehze05wbiIg/YZTI+0MicAO/28ctVnX3MdRSLyDQXW/A
RHnvohyaiPQlLIBSTgtEQa725SOOph176WFQbQn8iOzvOiY6d+si8Iqe5zOgKRwj
AmfvXqoSiSMGASb1SQRI916Uh7Y4V6wfMeyBzao1ObQ+PuSM6hMLE3c2abUulQHq
suHeJxvOFkTOothWhMoJsIxMzamw1TonhFT9eLmztXWJdZPhpMT0xeyRcCFcLSJ4
MxjuZXLXzllu2rgAatCo/Ms/hLK0oxBrpN+0XxK9qn1mA/vU2gz5TjRzm1EUj7nw
FBc1zqdP8Frb8OQvEGkVg/IBhabUqK6Se/IvRuNTF8Sn1DvFSvB0o5faiUkLJvzv
Oui4RRm6GWu1J5vJjTPX4cVBYuJ4jmQxAgu2L/dr8hPfEZlJTf71VDYkyoTBCVbB
9H1Huc5DhLCoartk3mHvuGJKSXuc2oIN5Y7wd45Rn6ztMk/IPPFOqQfRO5R/9RuN
wcifQG0lEFrQM0qcgYToQkV3TMLMxzdlYJnG7r7fdeK5nJhZEVN627XtVfLCZCJd
HOcs6sktoeXADLTAFohMr+jfQCBGMa2MpSNnoR5Ok2Mkfdfe+Swyl/XJZ24/ZC+7
HXdF+XzM0dGWvBQDFLlclvPk5+Rnm2UIHXJ9ozpEe1GTtwK7Nx5qUcgE4NjhWfwc
yJCA1Dv2w0rS306IAOMWj0mUalshBWQsz2X0gVaBanYWsPIptJ6TERvpF21wknLC
qWIgYZWlNcP6aJmnaLMH9djrKaVwl8vWXncf/FJaSqdSUbUAvRPNaxtCRtS71YEY
1vIeR8mc3zwZUsfIcZCW8Pr+X5x9pIe8chc3VXqUaUY/zHE7+WNdWKzIiN4aYEOM
Gra+Iben2eZ2NZWTs160PveiEheGK1qejMWQwuZ6BfQoU+dM80NYFeq+8MzYvNoR
+6ms3LnN+nu6rz+1FvT7hwq2gAHnOTyPnQBVhmBQaODa4TJgj5TSwhvuexZMm2ef
l4W/kq/9xXbRyMoGROX//HdD24RanDiJsnhA4M6Oams1yEx7zEKzywVNh8i2Pfzo
zZeHATXOwqOdlnkTM19mj3pLxX+B9c651v1ocFCHCjqNOObEdH3vnOo3j9pEmSIr
aG0OgldHgoZrcIoaTaXdjpU7WHnkKDvUBjl37OLxkVaELGEAmh+5tk/Ga0DCX4dV
zlHrXrTBmkVku/rbqSFiUePDb2Ng8sd0u0uojWR58jQXHaxIOb0RmbY1pTmEIEXh
NDYY+0qVp1/FiQoSVKZpJ8tiRAa26Iqb/n+Y1tcT3Yjg2ZQE4kBGxQG1MjmpVGH6
kjbu3JJ6gQ0JQUtv5KGnwBIY+QNV7zGpFZUs5hUvrX1xWk6lZ3EWdkpx7uiykd/B
LygyP0iychpqbPqFxwKXUDYMZkYQlJ9sRl97spQjKOP2VGbMxXAaKh4oJnR75Hz7
PLCennbTIHmTf9bxJZmzPO5pUn5yLR0savc7/hH+ZIyExRXhwB7e52FjIlSfeNJF
VWlN30kxSwpT7ZCDsYRLowUk5a1/3jBPeHCvFWO88WD0D3NLxYHlhYm2wNCOV373
2DPKtGD1O2ee9PQZPOmfWUKxUk/1o1byH7a5TTvgENQizuHjGBGvCd3l4oGCVqps
HNeCRiuxDlYpxhJJtpFqhditb8otGbJw/Qg/y3UEyllSHO8hLn3QRZqL9J8Z2L52
pTEHkFfwU8zOR9tMxvN5Um4+GP9xKwvf2IS3D8pJ1dCPd/6ePi1i4K9fDmBqVy9H
PM9Kt3fcMwL06MB1CY+uo+HiNmxwTmlVttl7z+qVSRaQoZIOtQMq+0nodatkFYjK
4LGYPFs9dcFZkeNKjeOXtd9g6jItotAqFgOWZt2Bfkn5CR+cixW5Y94cfCEu4Huy
Xfd+zyTzvCeimXLvZtxVp99Gi+Wm6YSfSObvg5zESdXPRTiOIoTzP64rgf9GQ+0v
g1NecXeTRY+aiNgjPvVxZfnmdkIroy+eJNvOiF9ADoreHfe9PL++h+CiR4mdl59t
52alvfI0M9h3snlqfZZ1d4q6MShhLLdX0RUchPAGm3cc/G4ofz53dNGfA2JT+7z7
bQH6cTK4kabrF4NMV1K/G3zlf8o6g7qMMoPA4Jax1Q0fdE2NqQ+SBpVG3d/6m6ka
5i/63t4cFjXTWtTuG89kM4LDC99d/QqTRsXsDoSPLx4=
`protect END_PROTECTED