-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Cl/5KlTYEykhcH7k93eVF4rcXvEhhDdj3Vckh4iZXyftABV74ORiyBTaXG//3p6R
AKFdMWoVrNIu35HOa29Y1Ni7SWcbcAZcJVnLES1lVYZSbXkg1bTscPDsCosmaVkM
1w4rNYwsIktDy2OtAQZ48b5NwaPL9aCzZQ5wAyMmMm0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5374)

`protect DATA_BLOCK
OA/eNa9Ti7RGojTe8D04SUAHc7Dv34bpsioKbt706TYR5UOEmsRVJJRekYK3Fm5F
9j1+syv94+6cYmUuZm6eopN/0qMMbMogSIS0vtsJIRvebDP4ZRFF6GNaGeb/KXdq
osHbQzD/o2SVrmwrt1uBXPCmkZNYvCE02FkMGOqjwwVcOhiSntoJ23w3l0ja8TUA
f8bMG8wWq4eBNIOxAGfkd9s11aNlsxrRCtob0NzQOAM1dqXGPT+asH5K4gYAHsBv
Ht/Vc5f/gnaQaxbMCPSJtnrGKSVBD0lD/Q71ZEMcOVqy0sD88yEMl//wtxL/BtS7
W5BEhdMZCp+FPSt82Qv5kKLSuFIEu2gJQVMDreM3Yhug05snQMc2wbocOX/AIlE9
BzSt4jb2k3O00vyJb0CFE5jWADxDtoaflUt3rXIZc/vuPjS1yM9Q9ci60uSi01lN
yzZy2SIXftkqhXZrcd+lHmbXNBI6aK1fBt5VblyOzMwO1rMCmOH53E22VAiE4nFf
jhNvSiVlTg4eyIbdJYV7IC+cfWm0crtztWPdT/LYWbZMvBtKk9Pyw7W7HneMfZcy
Ta+9F+6utLMbD4GJHzrhGj+fdHwpfpeUBRa1Ta6OmcMdy2yS/uqDfPrRAN8qaHHc
0z3SxqeXGGlpz13FudkYS3F3lbt1dF7T89S6nrSw2wEjLPLkZXjzagbo4EerjzR+
Let4YDTFh1uKHs0oU3m/nwlipGYxK/xSZyGR6JHQOOop5kdJe2K9tNZeL30VuRrg
GAkF4A/Dj3KaCXEVQVvVhnYol+D9CT9bBI1WMQH43Dz0j2J4/trnW16ysbAKsdkV
wcfVxEiCC2uwVp2GxLMA1jg4o5Ip8cC54WCj/Xza6HqqLIjaYgu5riTHSarCZFZS
8Mrt+Frqoxm4Fv4XuH7i8PBe7EetWA4+brC1TLBVIVZxDqBaWGtIdChgQULLtnut
GZOsfiaD52waoBTZf1wLfZ3GrfJUcQ2HonmSjLAK0Iz7dztpbAvbAq9FW7jEf3ip
pytPghjwQG4QrGHQXtbIDVPFQJpd/AYWH7L+83v0k1tU7kSiG1VIp9/7CXZuHJDn
dd1LDEkA1+uqn8YH3DZ58FTLf6XtuuXBpNy7EVQZ5EbAOhZ+1Q7+xSZ3h8aQal+i
s0QVMwj4rVhMI+PHo4JCyjHFPOhewydyJIJCiY2EpFNu+XxDKGZMzLxIEF+G6BkH
/gzI1POVvgOe8Yi9NDbNEuv6MrtUrQOPFjnhmv0J8So6AqBVt71NpkYu1aPNiiVY
nVtNToa/528ekke9h3//LD7N0x9MMjSI/qx+iKfHhYtFLvNnRGiIhZaw0S/0kNgk
segzsqe1II0yMmvey+AiDtd/N0PQHnyKi1s5GMKM45QUHg85HCTIKqo7qt1wJsd3
ttIhTtKQ5OXK4XO7FIgG44iXRaWR54Bonnd51OHXWTpv5U4mZC4qMm8JkfG4pGLm
3z7gLzlvUt7WMEDTKaOwYdQqbFAHuIDm1tCkni8mUx01yRrJWw10r+DPOIa7tVFQ
JvUG/UXhhW075Bi2/3iFpLBCyLTalidssA+NceGbrtptI8e8b8moPsO1xZn9BYRz
+P93zgcBCFbnkcbBQ+ShUWTaPS0t8/t0CHB5YOQH4K/jXhwUcZ4/AdUvzRlPknNL
UinjjnFWERzPqRtRog98j0kJbcvOWfgS2Gfn1oignPp8VEzVjWxCZP61YNyFrxSn
ODI6YI4j94uxhSX/ol1E8iFAUb4z3winGiXDw4/uaJQ2WApbM6bEcPCZ5j5JyecP
m3carn0ryryKVs65xCJ/qhrXtG0qvN/MhOrSs93QtDDmPLsPTz39rnWnC/tCIetx
NcFCxZDedBRZqylBgWW/5kWIdesaST5+c7055Ftytz6cjOOl5/nGp2onQ+ydZCmT
oq17blydehsPl7kuiWGVH2DLPk/sMCeo6SF3kDfkXIg/Rn0YMygEn5Ey3V80nsj+
d2NArRiDyPcld4N22A42IaqcScu+u1OEZDnZQqKe7DP6k2AVxZG6IhjfDPYMAfkn
wKvkcskR89fUPaxbUqydjTwXYZwem6ev8DoZLoGpkg6yyRowdWNXU4DNzPYb1PGY
gmnG3JwpK4CMCz13Ke5bU3z1srvEXsAJfs0uImMgq1JMcEhx0+g5aaVtKyKmBdGc
COohFZar0wUYdoIorfjgoWvtHx6aFZt/JBIg1+zkM5xMYmVHw1JIuwds2z3wM22G
E618FeQcU4salSDPxYe6axczWbe4ddsJ1MDfaHUnXtCoO1+/XqyoLvv7ujUaHJCi
kpTAIsnIX/hVKuYwQ7/oxDNerTDWkywH45aagM4pgPGL7F613/wwGcwnyGGRKuvV
InYoCt+eau04mAakNkvfQ28wSJbVa8gbi8YBNelTSdgJZ1Yo6KBqVodS7awxVDmj
DoLnXDeEpGIlPIdzflmNo3Qw4fbsMkO9Xj8+bRN/1nM8d/PQ2lfFc3xt4HYlZ+rs
gUkcX2yAz7hkGIkgUf4iRHFu0aSiMiKWXtwjbFB4evzlAb0w94HCHHbudLCWgirD
1XnYWkjC4BF1XaEWILq7b6+AQCQs7t7wgV4lhlgjgvE+QCCbp+epg87kglSA8RKX
v6etWQTEbjrzF8BQ4dHcpfXamkzt/tVgPZlXWG9KJuNbK0aZw0UIMBgodN+9dBrd
xsymzvE/vyhTyCbL8h7rYcBkkD1EwEUxzS3mndCbAt5aCeD9+wNTPRV5hnETMnlw
IPKjv8iLSqf1JEWTSeOrJOz3G33giGjpqvp0Wd0/c859H4yyCPGfFQI/Slon9+JI
2IDr0A2BfJNgg8YEEbMGy9PzplR8inlo0+8UfaxbXacYhg+iblHy5PYB8XwZ5hsL
T11ATgnGOcdqWgJ3OJ3/8KJixfiyKGkAKg7zHgy5BWn0zlw8IobFkEs08txJInuN
Bhm2GxfRHFOPWaodm2/ogpjKObnqNeA6pbzd0O3mQgRLzgIER2w5tUK3LtSsC0XU
g3NOqABOoMon2CxanGk3Ascgq8IVyjpqJXhTswGwy3Hiq69Jraqun9YJxkR3sTfI
+iFqPUcOegArhQnfrxZTqIWDB5/YOjrKe9TMZUUz8Z1Bic/3g5zqi69ISYTvnJr2
O2VoXKQHoEzeoU0se39SsEFo6Cx/GshFQrJ5mYSjM7g7jsFP0xNUdR/mwghjA+6F
1PL7THPZ6TFhFp12kffxOIenwzmcXTQDZpbMI8LwMrGJNMiiYeQAvkfi3nucmBmP
8+zMEj3roqlUA+fQ8m6O72bWwhoJozDMxJvGRQlFE5k6UTAQCCt8jus/VyJgcuQi
iy1ztOK18zREHDGqTUYFhCFUBP8+RWaqwxwOCKj2pGMdZ9RLeDvialnFrzyzOd2M
UXhOkn/u5n3oHWCE0OaFi7l5XokRUXOFJMfMfufmsl6q0S6KQmQl234qtENN81XU
PWpqxF+0Ro+s2sIwWZNyxPMQVxx8vsi1MMNBDlcFPr23RVeP2qn+8OxAj564pdgv
SJTrQTnLk243qSSXg2OB330yUSNqR4SOlD/tlopOwmPclkimMjvgClys0Otu8jrz
nboQzvb2GvdatY0zawC4rTp5vaPFZC/ipfYR/cUO3uXaogaDU3wSOXull/5x0Jhi
ICGpGAtLrCSkU8sONgqpt0F0F0uwRvzxXhGN43CIOfZgmwP/RmsaHefT2Ujuccgg
ZN37I0770ku7B3m/pUk+vRYclUaNJ5iTDeJu+RH1m3tgazOqeB+kS0tvDh9jmoGv
nWRGL+p3YTkYvWhrpKudnSdstw8vuPagzViCZDWd2/92nsztkcQiMt6KKcL7z51Q
cz8DjepYHIh80N3vMo3IPbv4MpXd5wfvTR9RIl/Otb7VQL/eDNjoTZcXS5bILAP2
6PU0bYFuz43jNLqEEy/XnJ70T07PRvD0uJBs49RFWoDpN0Tfc4M7Ga8Pd5FsyD2n
luMxk4KDHblkK8beDOP0ECNpRYmRFGGsMcThBXm7i03UApSuwQs6xMSZXB5ZeHbU
fZ5td+GO7sbEDq0eYs059fB69yK5sLdlFUSq2pIOHzkpoyHNoauEtC16GWH34orK
1lyyukqgQvq/CRKGrPL2DdByXARNJ/htOU6hfv+8xYtp9XFchFgXB56AvwiG0OBj
QIZeaSjlRqFYknNNmzSHuekfbiLmmxhSCdYEnwlAOyBqoX0RjgpuUocHYl8Lu2Mq
WmICMh59v7jGplM2QovHsIxUSAog5LSTA52eZXbR1reSdkNoPynuZRYFYVyi7QEf
Lbsb4MyQlcCdBSs1V8wBiPniBtRBoEPOekdjoMwBL3/8LZa9IcXcnXjVKWzepX2Y
3K7APf7fTP+Zfatkq4qRxftSFcM7bgpRIkibJXnvbpPxGuRklnwqCXq7T4/C9YP+
k8EuTEHDaAlSen8BPj6h8O05CV9raXzBgYarWEBvZzkVDzXFls1kVLUdeYnMA3ao
wV9wrjiMMIPWXUkYeuuN76nI/GmJDHfwywxmBCal4tjtVp2w5XIQ4MVX3p7aEWHD
ztIZiTrbxXbIKad3KJm2NGasISe0xPHaNop6VFr3x+YkDzpQMy7U12Js4GTGFUwM
wvQAG5fHKDEuqGMRWOortY8uniSaDi7wBChFI7CoMKhw34iklgQU7HKyMrWKM1+Q
Sz3oNKaYuwAWW9R3VPYPS2AOqtfMxdujG3ir9ruxejtzEPeaHivjf3Z/motpbTNe
8N1XD2w+3n1C0AlAUb6ZTnJhCQOsislMM4ccbDm7BSTPD/RpUwzmviGmcEO9fiYR
HER5ilR1Cc1XxYUhJd1lD/IKxtrRKxMAUGdBO8QRXsohsyzwAaiCiDVRoN5aYOvF
gcqNX4v6Uwf0XD5f9VIZbrjdqR4pTusrBM/uE+/VlIIqsEKVoJqeR3IwDbX1Xc05
5V7DRzKQOAEaD/jYMOm9WrilVH3LmvWF10IDM1LBDd+nfLQlwW8Wy2DEkAaDQdnW
1dzz9kag/DrSfyhJVIhrMWSk7r0rL5S7YlU1mDiEj2UqRDE00LJrn76jsEg+hijm
GHiUNOIlLbOHpghhDa5Hz+OMtXRtRKRhgo+e4GDEippTWTIXKsdSTaJt7Hhz2AuP
r/bz68dk3rk0LHjAzXEYrhk+Pb9Lf6rePgTMrCfJ6r1Hz9BAhlNEmP7O+1JaFGe2
bB+/0mUjDadte5uNLXCwS7fbKmde9v62Wektoh3evqRZhSESQ3Ve/O5yX6l58jzP
qKUWY51Hftlu+ZEwu0HySJMaA63JGpmEtRm9e8Mm92OUXInIV2SRSYveffXDgs45
Q2hqM0doI1rP192IFg+QFgPJrFOautMiSWDP0GNV8iMemsOHnPdgvycEY2c+TiEo
Zap2+iiQydHPXehAfQ8npdeA8X2JZZbDloFibUDmD0IQilqff337r4Oz0F9NMrOY
BP2g9z9GVHXqh86Y3yUnA4cjYhDR6zauUJqLhdHLZBeex5vOG9vpuzPu4l25nYQU
l+e3tprVUOdLZXyo/hI/NdL61z7ZxsxQ1oKybZeJhuELb7pbtUJMHqVtX1JSEaZL
l4KWZijc5A1IDqlXsNTbApGSKqQD2sHIhMpisHXahqso+kqr334miI+OQSDY6DL6
mcYJ9rvrs2DTdStJINbOsgbephhyLjKzRC/aTByasENyEYbxccdy7OrOTP1jRWFS
ktD1WHmGdGoONwZPThNcbGHU767+B22CPc56qbVLTQ3MA+j7W3+SFFgh+Eq5BoAO
aMo/joGzc0rEkapbL8SEj6mnpnou8ZBEiKi3GywlL/e5EL122BzS2nB15O2B12l7
1BlzN0tsiHba0faTOyY3MBbJld5ruw3+Xi5Yh0MgVG1YhG63ocrtyGFGO3EVofQI
XrnTxyrOopN6cAZ/lY6mdQGT1f9c0A9Ie0MM5wCYXgE3Ma4XxqEOE+Y347FRD7n4
V54l+D+SPfxI4vYG5YbwDXDG1IDWaXTNsroiuE90Rra/BAUwWOKxvEckw9zfE9ob
t6eEeqeP/9PAOEH9NYckJ9532a8nyn3PQjAytN46nZYkde3kCTaMduz+UCN/IWVO
vqDea8VHk6uM+X8BGzdSu6nT8v2uRKfm2Uf5M2AFBDxg4mEjvfir/s/AO5tTztgW
YxvJ7YBf2smOxjbE2t3uADktzszUXhYJksvGnCokSOScZyKQZAoi8zAreUTtz8xc
D0QFP96leKW36HyYvu0kA5KcfHR0RvTJnqgdD1EEnIWgEDw9vQ7igJ+Czj5zwniA
6sGH3AWxy2VGLrukHAH3gLcRycWiudtpOK75KCAs8AyqPU5I+Or0eqNTF579+1oR
k0eXYIMbBAACbG58u7e93nhD2kGsn6Z0bIdqohK5FxXoRa5EAyooRPjZ9hnTKbe4
AOdIzo/YLP7V/aY3UY5qImEZWEsvuwD/0GPrM4Dvw14ZT4Qj2y9tMZEDb5jgoDiC
EM50AcV5FF8zzO4RbL4jFkFo9yH1kmpUjqH9EeZ193BS3EuZnCR+5NToyDDerou0
Jr6tOSytBwABiD8OO+VjQ71FpmjGFEKPeQ6KRkNforwPnbp9b+5pa/qCOFCamsqD
BTQxAE2s7SPrOXERwYb5LhIP5QzMYhvXDZMB0cLEyBwBJ8AQPuTIRWKlvkcZDh4o
TMk6puuSDJx2GMESTsGDkV2nrpx9IaUWvsgqnwiizRNIPpz/xen9a3hF/E6dOins
TBBK1tFRl8h4GDDLoiJ+2QZsQRlCxF2kpHOBiB6gTyPQiTGrWvbwO06LsXh9QMbh
na3+x45ptdyiQgV+qbPSV5Wr8cYLS/LRJbvYDoV2XvsSQhIYnIznHYyQxXmcjNOE
R9Jt2svN3NIjNIFrjAKjUFyk8Qv5PanDj44vDLpEe66AI5hgMoYDWHeTep2NPML6
f4Fd/IRh7m/i3xKk6y8Dtx8qgHGSxHu5bo0ZbfesCvmqMpQAAbuPmFnNWsEiDi+Y
Y8BJWjlEsSyuIFn5fKJ6t43mVm/g8WK9lzDmB5HWY99AA+YGTG6z0/U0pdqCIMBG
hi1vAqtdL3KE3LaCi2BpYjtJ6RdKk3S3LFKQFBDn5Oof4oDkBifYuObWoT/bFhsG
ferW5weZ0gXyrQ6ORFknI/b6cLVZr0Ouk4fJ4tHFt7H3aYMzRsnHHQJHY8QbGJdD
ypfX2/TV4kLr9bMvEAPerw==
`protect END_PROTECTED