-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
cDS/UuzOZNvMzfqD9zDq9BjbGcFaEXpjgwfQnMlnsS/pS/yigWIdLIIkJWljMh1D
XjBhQDf2s3GobcOSOVjRPTqGm1zbXEPzdDnuufJWKjBCNrleFtHlZ2K2X5zW6WWy
ga83IORNIV41osim2hndW69LjXojWpxKkR0GiAGrKsg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1650)

`protect DATA_BLOCK
cyHv5OqIAPXFuZ/4+YY/jQMSoRdIxt4s3kNU9flipM1l66x5XFaDSxFS5+o1waSv
eda65OdGqhX5uZDEo3bxLqRHbo1KZx0lEEQbHrmpholFYFmAAlXu0CPmj8uwUEUR
A6nBgR7rTGrpQZ5AIqjk7++JXF5XcGOPSQ9qvAye+f2w9IU57U5qQ7bvUilFQfhz
jnKzsfxec1INo5igzueoFbJrcJFONxAr/A2OGMeFUJQ8GvuCwJeecxqJmM2kFSbb
aPTTS1FelO09izDHPpwYbSSKCZuzZc49uhEQSAnkPQ06VUHCdDfBjMpaw7MZPCkD
ec+UqUIFMa0iffiGblZ3F1tF7N3SAVfdkgcDBcVsOYA7V2d+Dl+o4ZIyyrgapuWr
l3nAwIirpv8SCAfCceEFwvCrIkxSf4uxsEo7qS2Xs4WxcQg9V2jPRiMaZN1DbZJH
8Qonx/PjdbxpgoDAjnOcm1672ciJ1+vPH7ZtmPynApKJvCJpy+N1V6ej5DwNTZgL
mAFOLOfGq1f1Lk44/R+kFvFZ+lAgX7A4aGSNxF9bawMFk4+NkG+AKZ3DN333Cl3l
BgyNGdG9DGCfp7WzGA0cK30jBeKt5FfIPWT+ovXvVC2BAyzjyGhSEP8OjA01pvTW
vnzjjCtyHkUn2mekTjv59uDadB8H1eIKJaJw/o8Hu+YzRQHLK08JqhzzgGXroY63
XbzLcyb8SaxwbXMjQKgbTTcZvDY/cDrSSvZ1TTP3a8t05hWTRCEgttYRs+wmiPD+
ixYFI4nZb55FIHy/RPHOODJMlSw2MMhH6aW8L7V8/uOO1Z8Js+ayTUz2ZmrTz56N
fI9XQzNoIAwqPvG/EAxl39ytBpCPPT5t6QpXZoLRNSBR1G3y7ojRcoWWZvtMROck
gGh8QNKt0MvmDRBOQqadeUpJacQBJ+zYC6tP1cyHJl2gFzfrpf+ZkHnFlRjZGQAF
3KNc3RtLEjpdJRiGKv2+AAMNFKDq09ZaK7GOBd2qpExbZF2gXZFutnTzFErapnfo
J2qw8/XCGuz52qrGBByIBSHNyGp2WPkrOgKikOhyUqzLgeXHiBDsaw0jQTaBdKkF
Cj5VQI7wIoWEeQHV+Rr1kvJ/Ic1gDEJxKlOh6RReg61dN+SgKnvNMTPRUjBUoPY4
tdfksjMeUiyTAGqtQlvkfxsANvwK0vKiQRZzUwIMoI6NcTwmJpLstIcPDTH7erBC
zRoCUHXtKdWLZ+o1ydrwYNc4JP7vo7ad7jArsMWjoMBDFN0BeiB6mRUHhNRmWCGg
9KFq28s97LLfUDckI80Wk20Y3TbLHrhdK2s0WLOKhMzWCyUtYzqcS0PqFKpfOJAj
0Uzimd0fyPphU+bIwVBix7Z0HDs/+8howq27ssmC4DIZWik/UYgfA4WZGf+XGtAK
Teeen6L42shOipkVMH6AkEJqtFt7kSWsyJyLrBa9nTxR4bYtzWoGwuSL/RT+hHrf
jAjYZ9A243L6nt3RXKxddaUVrdp9Qiyjo1uhePbQPJeW4IuEfb/uUoXaDRT5kTbs
jQM2Gs1KrhXfMSIy15bncPfjQxW4cl2B4SWMa13PLst9l0qGYH4mIqzaewwXSKu8
cJDZCuIQXKXgvqmo0Gcg77BXorIc7MT7QjNxQ9dT4PBqUM29/p51QLqCfy3nmh/t
rd4WFOZYXy/K59fchp4UADbSoHvo/2nyV5z1Ynt6Ufk4kwpeykp6N3qeb82xPrBA
VeFaXuhmUgHTHOUE37qt9P1Y3NHQ8QT7R6NtTiNnfKHZIvLUzXIr5Zs4/dXDuS/P
lhwSVFHEt9nOE0ZDg+xnbZ1cHqh+urVDCF3ZFREwVTmWAfCxHxXqdWbvCiY/VeDg
sS1GnQgQUgqVv0mf+9Ua4qjTupscY1FM8mobFHimIsqggoVjWYKJU5LskHI4U7Q2
wu2bDyM7Spej3ZDdTI5GbDXdkR8wVdofB1iI5albpUqpnQN3ApDI+N7VdzTj4xwY
WlE+nMErq7+pCJ3C8tO12/88GHGYW+ND9P19NVsAsWTw1MGt6W6PnpEVO61StEoy
K+LflPI7rsy/8soJjjAMGusLZDNUeOqGGr4IB+BNhMaBlsuPq54+MDWRZ9xQAcxL
17/5QeTyeriTQi6a/rRG+ZrLdeJkp8zEAamJCB/3qR94gpmpR0Za73jyL5FxGxak
WR9pfESMZ8wzji7XsBOANpb24lUABkFAIZmOD49uxmgFrouLwiIwgtkjHPtmuImY
`protect END_PROTECTED