-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
JPKiZAIyDLebyWm2JSTKVPUYozUg9ZDhkErrOosG63JtaVHv3uoj1V+x12aM2rSc
DTEQuNm89XiEfuVDEPqlZaD5iKLnXQbqvEq094A3Ptk/L2kDMCcCgbDEPHIiHDnF
HDRRmjWqjYLepy+QHI8lHE0MTbUDb8ZWKqX2NGPQMs8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 42951)

`protect DATA_BLOCK
UBELohvKsvynJHOZDRb8xnyIo2PFSMf94L/sa2SLigban0VPmB0crolsxtEqHymI
EfERcaUe98x5btDB8OWMO003DFRGPdJ1G6JNaiTm2JnGrSQtqNNASOiHhx6nOg7m
aeEDC70xkybwWjMMZIVisYHaqG+dg5U/qErW5ZLgALeyLsJpULthVPbNnOQnuLSH
BcuW2J9bDEAYsy51TiHthGC3oA0/l9AgAadIdtl81HlCWhWUxeYRdpJK3hU5tFRT
H/37INScxTbST6gnj2i1WZifm+HomS+xK1z2sPvJEYLHDrTJ8MQlvY8YiHfj8Rt/
kNZdTMgqK7KyVh4KQaIswVpAbUMlqk/RyffVlxkXxvHSBxt15zQkAsF2J7iptcUE
xk2C7NVpZ8Wkm0UnGeAUc2Wr85zfu5fGCxF1vDhxvFBxJq80+xP+m/5jDXZwd6Bk
CeXu7d5qX7sWcctTE8dwP+m7q0gi30ZkKMGvUsybOFObAu71uTYqQDKtdcvzjN+6
IsECBN0KfGCJS6Sdk4yAzOsXCKYT4ZAzch80rjCNb3FV6T4euHHSn5XUfAQ8CoV/
dHjt3O29sqKzX3nWexKyeKCePO7Uu9BnOfYuUV/BcsRDi5eH/HqF2OIGq9NN+T94
sRgG2hWU1cvujRSC50xdmT9QVHOxR/bHEf9kuw+n9kroxRoSDN98QQbdxY1ItBwR
6UYabObVaEaH/x8enHy7oDMnME40IuCVBIOOqU4hB0i/azLrbJYt1ISIbIKHmpa9
VXjGDkZ278DDTiL+EmVpuZSx4M8oYuvPcl8HNY+n2NVZB0/xbTpK+4VTkNtz691Y
gvF63Lzit6Ci4PtKQLtQ8vfUwyieotHkmUu4L36D8X43rvGP6c8/ZdaCy/mUxiRo
vl/NI6UvZ6uYMWQD5xFaDwmabk1RV+urE75lNH0OEb4rsMlE1fs3XpHN7qkgKOal
XKT/PTEznLm36fk3n5yHrB+uCTgmODFgEW8CRVdY6FQeHiNib00QN6I5bWwTR1lU
YQJkvg+GjoEmvTPl0uHXaW84Kc+KEv6I/Y995jET4f4PVnaTLBtqHjHL04NrRbtW
uEyQauiVv0XdAR6biYeFDBTuzWSCA8aA9Tbj66MA6Fj3NjzCahmH4LzTG3wxT6Ef
ZXxyaEY6WAa0VseNAeotWw9TpKL+0i9be3OAeRVtsIRfAlQKvDaScve3xbAhcUrq
tTokqQ/KgMoGI1OBITEqnJ3umvjoVD34AkwcEHHhXYbVslCDg0nZPvFof14YXzNF
xXlOTrXPdWI73gIZcexEcsmOWbTI3AZPzSAMxjPhsdeCLsBcUdOXvXBO09m2UQLO
Rsl85shjy47zB82tYntpHviNpBCgMgq1AauPcHLgvUpedh8j9RvRq0mYNWFzfaz0
AnKhuc/q+LuLXCIIEsjV88c+X0NTtHUple1rJBNnIC4AlvIvXuG4lhsZFiztsn+U
TpXJ2sAunUyuO4w+kGCFVbrjKf+sQ+dHRkjZOJ2y9aH5S8GXzbmJmG3TzlkmSsAP
+3Rfk7uXTy9GjfLOQIUDwdesgvRQu9tbsiex0bqSs9Ymf3nTHPlI/VHpE8xXwJok
gnr8lnEA+21WIIy43hddY0sLkxSM6TCnfGWf6pansF+JKzSlNpdygglBQKVyp/L7
gfVLUfOBmMQ0go/ci0MnfgpNM/3M9mJVgHy5hQVZAl0Ebdcaqxj7okhFOmfKSpxZ
vcUmRDKat9KbCEZV9YvCijWYstJ7JeGWVHncJJRuqkiRVUFzsY1k0hBDwuOJ2b7b
N8vwKi8M46Om13pPockBsFfKUhvgtY8FtyLsN5+0nL+9hfV3Yjt69CkJNHkBPGQ3
1lYg6pe9L0c1wWlITd22Wladym5pcSLdu3IuNTXak3YDioDDjPXBXxLmzt3zQ7aE
ywFhUUgRx/leqHjUqDH0wOlIY+DiCwSmHkdIsbDAcPrge/h2LTIkWcf8vxABJbmM
Bu7TX11CG+W93WAINbzrQjoRaxTrlWhq31C6jwWePkAnTGlfe88nrD425kGasOKs
LsRs6RLpYqZjM2Dmnwpq5QMHNfR8c43/JNFgjR0NGU1MAIc+Sw5BXEae7tpdrrh0
suqeSnbxlIEff1ZBtyU16I95ygPwHrmKRpvMdlscAub/iEE0IhVBLU2VX8kSDpqF
vSXD2XVwdvSowpBiwfcWHnuND92jCAjY3YTD9DXJPy/RUsY6cZ4tHsQs0duUdO0W
T4Jz7zxPAFRirVFJmI1oNBNXOhGBVgjSh9wqW20E84voTshYaU1v1aSBYcKnY/62
cY9oYAJYc6L6kLKL+cgQTRKqeX/dItwJoW7KEGaZkQ4aApbskHo4J0BcU7XcrWvg
if9UCsoPTITQH/RKbjT1+VtWt6Ir+QxnOHIY2rqmtHuT+KQpuWpxNOW5kJD2rBYA
1ga+UMniS8ObIrwSEDWRNKtYbUJGs/vSjZriDpGFWsDFHWgeA+H1Tsu6wfMYJh5j
aJgGhFKh3v3ZD1Z9ExMqzu3ndYJCpsw2AoKalvTodWkKXOXJWAiYy8u7ofHl1n9p
/M/DuRqB5I8gdjber47Rndh3VC5NRR5Z5V3tNeXUX5T0lbCT5UQIlE1HEJWlIUX1
3qZM2ub358zTReG72tlFLKJAvn/gqpcRUh+aaspwWkh4dFkARSfZRh9wetmQ7O32
xBhp82TgpMAWuuLPlSfdKAz/0Ik5Stbm5wmy97BV9OhXNqv4Vu7cQstVMZ0nsfwY
ViaAJnlD/YTekIkKXufvV/9P7WmKdOCpAkCUcAwRXOSNGNw0r52/bP4V5UOn/gJp
rTrePXFIaFrHhxhwNsx/iNK44oZzwYfrqwGWOYf0QPTq9+p99TfY+vYSXJJdLXeN
X+gnw/i9auaq+Y5GND3RNURqOTkuPrf+hNYruEoNMyJ1QW7iOpa6Xl9B+E6Vn4YI
quoDD6KxmBC51KG7lHjFczYAmjAoN8jFj4w17lhZsfzrzAH30l8k/E72I4iGiynD
4XlFaIBBsnh/2EG20w5jzhUn30w/V03duRP1XZQv0+ZI9WxlhPODBi77Si9Bxdwu
AZzOTFdWkoAyy/MPxhFYCGixfeamEgmeUk6ylMr+zuhHhtzUvij8C5PUzXUYPT/V
kn4DJd6u0qFPH74YI5+MQSWssO01ALm6qNzmebR/iQJpVsFmWUCI98Cs2BL1j8GP
cdiqqM2VW+rdPQDVoch3ef3yCfyvnYKFwgde0NKEGnteB0sCDLNIe2RtcX7Jigpj
4ipCWTuUZI3da2Zndf2eX8BU3OunnFVlu66bpk62zLli5rx3Fh+bJmUYleIySjbz
gannmDYhdHmT1XrV//EqmOni6Cu9DWWNYfK3KDypHgNgnfMt7MIA8Avyt2kMiMIY
XXojCk9eU+gcBjxf7So762INRr3Lp8knTQdULWwiiROrbjh9iZoOKWPD/I6Dji8Q
v4AKxut7Xq70zME6mvZqajuw0HecYgB2Vpl0jl6r1ZrvBEkPkfCeJhZPbyl9KfSD
wZPhfLyp4hBp9lQOLpou+dELKjOaAvNkcpfwVA4wtzBvZLWy9hswHRdFn68ChVNY
0yQM/d7zxPMgHHLc7FE6MPlKsqfTT+1sCDEJkpHreZzW0TZ68Z9OPNuJbSNS6BzT
PtjBG53yVv+NYhgXsf+9kg+K96P5R4rdE418ASlv3kbUBO1kKDLpHG4s1trnlvKK
ioEChs3Y8npWhTlDo3OJvXAfsNTzuS0zgLBJaDFGKdaMSqQjg75O/16AfAP+/7Ab
Try0ps4K3oYXggDsZOuXFcbwKSRLhy1dFNBZzDE1t+HXJAWVryUNstalabBTG/3N
cOHHeTbgRqwmLLGQ1M8jqLdV1yuk7LnTJuq5jjnjtRrrenFGEmoz24Ph59JdU3Ne
mdvLjkjBs4vehhtyp1R8IdIpjvKtOfKleIQGE6dlI7vhqOd1juJFbb5CfiK025Qo
e4hIwkxvHM5AcR+cdSw4a3WoP9/6kwPFyg3gTyDbP3I82s8AbzeWv+B1GnnqQ9Ob
EoVewY3R7ab4VBUVWoX+OdsxRaRO9RRLXURVmDuKN3DhwzDq0EWWPx4I8JTFWSvx
VuAA62xmwDlj1ocT6W4QlhAqWmUk0K9nhftBkkNrjNqznoi4n+aK6zw9RwY4q0Ee
rnDb9VyS12JkSNn1osKrRqaXjDyPUkI9B7hfhcT/letdVLhzztKdmKPp/S9jmTXe
ArQBb43CbXZE1eISdCP0UEcWIPBHivbu2ndOT1371rQduaEF0uqxlt0pywl2V64O
eboZsbIL1EJPT2+tCMR71gldLDrY2JF8guF6Ik21NX3QLH/WvsJQmmxvcv0zvDgt
0MGmu5hCI7g9/OV+u+llHxLAPJd/fb4PPKthGKZG9tu9cYCnyYhVRU7X6Bb4sRtw
aP1l5KH9lxdgpXjUtmb3jUs/d+ZPeq+jxGbMKa48macAHaovvS9mDa3N6BCxdBgz
xpsyYIN9N9oq0M4F9w9cW8ClKpL1+KwijX2UACpV2kG7YtjFSMcl6myQXd8ubZmQ
Y93YCMshL3u6UVca6lW/sPsvnIbpmgC4WRRydKgpbk6hzYOrvLP0JuKyPNfxpw3n
rGiPwmFedKELc5KEtxZwc5LyghiQH4SWw4RDUTDbkHQSgQtrVAauTInJR938B2wz
gsPzAKNvEjgwhVc6Zu6vgWJqay6+YSwZ1gVVlpWIsxEY4KdPLsmhxHZ579G8DedE
f/8Yb+FQ7GDYTGJNcj0/uVkepFo+y25GYUj5lDsqq8uhoFw9qXRQno146ZxB+0Da
zqzvFil8RwXinzYm/kkaJit8ar0vR9HNUk1lEZyVx8fbe3AgN1GwIkxEMibAfTgO
V7DFC3ucbAFNeGfJBuP0wJzKX1wSoziHv0s6bMAkDICvTslt4OJMOoKjoGtmHmXy
j8vZNmgS4HXBjXWZHynI+R3Pehi/qMdbpbBKbNQK8jGCSH9r+d2K338CdB4kbbOB
BSW/m0dY6UJ9ItzpUq483+48rFXy3pnrmX32TflFtEc/4uOpMmL3OeDgOmBT7/xO
z2+d/MGIHP4+T0o+p/LsYn62vy6cC/P0mMhWmT0PwNkj5cJmh5E5/eBPSpZg+5nP
t/ZSoFMLfMPwGhMjnL6UY8H/NNezIN5QVurRif/lf/UQoeZC8+vea8A0OhZ7zZ9k
NRKhpYMC/qPdqiP5TJAOyE6JoXwAGaLlmpemU4XdXfiZIdsWnj/a05dbkUDlp5rb
Ej1Rim5j4g6RY220OCs3Q7ualt8NTgJ+fFx5EfL3TofbyMwE0bK0E0dCK9djuTDM
v8c9YOlYvPttpQuU5dpze1r2OpA45UUsyFaVIEO/xkGPwZuYHFViYNhYXrTTt9Ng
LY65GFM85kmNswg+mPWmpEv/U2VMcVIvBFbCf8lTEjO3n/qnhZ4m2hbMTUxEbnCa
LIfddnc8mBM2l7b19xe4keBaZzr5793I1fda2bVE1X+xw+46LpWz4WSLeK+I8/nD
OUOKSfpbm/ut8NDOIDHqlipyeR5mDn0ZDYOXLP+mEbJ/yddRwa3287HGcem3StWH
S0JkRM+10kPAciBz6PLPH3gQWCwZ+HCg2fC3SA8FUw9qgMBWqAm0SKf82tnQG74x
QJyfAPm7T82z8vqVTYPV8gHszrwhrjpZQOo7Jq0PK41VVlsvbnO2kQPD+V4Jwa01
ZlgUmfGEQUPHN04S/6kowz4xoA+dNi/61/OTPr+DU4GMLcN4sJfN8hEMofsLNc6n
ES6Qpg0N+uJ8F79z35yGto6BaWL7P+mYw43Mk8NP3LpQMrD1u7EaJtNEz2cJd13C
7lo+X59aJUdfYqVevdCKzgR2oU6dEfBJHsKdRcrhX3zfzcU7UEjt1DD83bpjbVDY
m0lczOd7hZCyDDTAQX1vGdCghSK++A/Vgay0dOODK3KjrBczX4qURwfp++uq80Wa
6brSIX6n6nRiLdWEeKtLpVxyUo9PLZ+ROno2EcSJbg+vV2m44QJBa6STAg/v34Lq
HgI8e38fJCajGDFi/Weyd2xwFysCn2ilU1hVseAn6anV3Gm1KN1MUm93yuGgn+31
CIYVoSm4GhsQrVRJOKgBESW0Ep8JDN6aqD1Bao41n2+NMA9UbMWYW1yGfUmaVKTx
y0qd/ppF+TNfkmDevTtRqFQUtW9wdPuamFiBDUX9e73NEZ3SdDKhLekHaEv2owzB
GvxPdWArFDXn9L5/IfX4Okx7NhCVuFT77T0EScOG3Z1jfpH6gFf4ckQN/xbTT24Z
Cm5HdAG47i+kyEUJ6lZtY/UzSIwM/1IJYnWNKwmjSyjgKsx9Fc0n7AYZU5funXqy
3ajTdwiG2kVKzTDuzwxwxx5y5YkaybC6Fwvn43dqU1Eo72wt8e1Clp2WlbEqA/Dh
BqKD0VGI+ypfKxAdN1Tyv0o2o2j1HT1/enkY186/iyOn8CZMmSHpcN1aOJr66QM3
bxdnnY+w0/+vmgsekaBmnsdZf3qel7XJPFy1T0dBb8Gc1CM4We566taUCK4KNZ94
f6QnoRf3Qi9BokMDa/FfQQ8Zd9mMazZA2J4jmGLUNw3CQ7sElCw4gsd1gHug0GKK
ad7WdJ5+lYs+napCzx73RaJB8bj1Q9kWVaug0JkNVbjueGuiopFloK2+WT24cNdj
liesSKF9RHsWRIt9lU7edMPDHTXaIBUM3VYav8bFS2PyB0qhiRglqWfCefh7YNAc
W8TA0MW45v49KfvLqWjPM2yQ5J3fPtPzFXlOajIxX1c8s3bhNkZ6po6OpzgQR689
cXjhIfQTWXE7NFk4YuJ6bpaWafC2dGU968bup7MKk0UbppZIhhyLjcnSH0P0K9I1
ztodQDiwfpBqf417SeWVHbm4/7Jb6yTKt+/HbIIOx13tDATiQsHOs30XY7EQdTaB
yvISGJWsKeoWB6GkQ8hGLShPUnYNoGAe5HT6Ay+uvKnoWRg+KDR2RuYW97c5rRhi
xsAibN2N2ildHURssunzRYQWqHWr0wOwcat/trjI6Rn8D/EJzkUYphsRAiFzPWd4
gvuKElzGXxsU9MMev2bI9FKjQu3IOdXof4sLwAGiKZYUE1uiP61mORW5g7K31DpR
lVsBRH+KwJqOFL+GkNHgkAujOIiKO51i/Rml4ms3mFGx6Q5ZmYcKhxdeLREGZ4WD
9m8RKw5WoPGriHIW91zFOhpQ1sEbg6Joomfy9TVntyndkBkVq4f98ry72xoHvS5K
YYXghkH71odsAJSChUTJ3c/Moa/2vMzI573zYRn0BR7VZlTSakU83zITQA5srQMF
WD5Ki5EXJB6Ug7bUqLUqsE6uLpBc4bz35caW7dicjOg3+nIs94j3OrLAoNH5mg21
yVT9Xjvt80wSG3ocrAJPpEmstl4/ycCeDUEKIH9yWdy7yE0WOh1B2oZPzKuKOANs
2OlquJM57A+MwC6y51o7d6rU0Cej2YieSLeptxuxyP4XWLidSUP5vL8mFczJwGhh
yQZmNK39sdkz+4EaYdyOzfShH1uvKCEQy8AI2Y5Bvh5a01Oet1Zv1Vdpcg2GNQTb
YEsSHcuAIcU7BA8RDWMCfU7VZ0BbBL2Qnw4hsUqKQ0cflFwgqw8AnXgVAXvBW6jB
ff44gM59Mfxr4I0pZuNyrMniG2PsKwCt4KhQrxhanzKdbOMSOZesVKY6uk4ok9Jz
4cMsvt7aAuJVemss1MFLo/pQpufTrwHzZ6yD5IPklNPmXFZAWy9oGeQjypUF93ql
ZE+UfY6cMZG4XkUF92v8aMw74LOhW4f93BnzyFXB6Q3ZT9Pt1dj+uE1LOexJL6OI
r320PO9oucPyTgGNRZbYyurjVNGn/6DFCrjLxH5O5xvr/gPxnOrARUrUBaXidPVL
jD5/+otCh+AzomwecHa+s7TlQZzElcOd1b8Kp56+uzmh/zyy/Mw9JhjbhSx1BHRX
ntKq0MoBMAEd17So6OXOGgsHgb2BpEpUvrJIbrPXPjvZ9h2u8mc61EPQgSCqUZ+H
Hp3MAjO999R01uuXyyxFlrHtKEc5jACJOuKiVcJR8qrakzjr/i/gnK9KeUVEZx8N
04kxUfWpVZ/W3ZkRQ7w3vXZ8dZYhLyENHWPZvBKFMZe3naoee6VOu8dR60FO8kcB
vNLOrcDYJ9oNofwF6TGzXg29otsM700JdkmyZH/PmWnk3ndXfUJMDyUSC8ABiAOn
9/f5HbHdBxv+fi+VlK6plFjKhAUWv4gyt+CEVRIVgTvmDfGTrYpB+I5NkUP45zJ6
ZPBQCCpbk27NuGyIcOHSU0Yymkh6mpbp59LRcfx+o45NrUumaJ2bU/1h6cv8EDYW
FvOiqiBh3moV+NFkJ67rF0ePGLWZq/rf0PVE3yxjVPFTe/WYIEOTSBXqVgUU4ipW
ziJSlzLRxYUnAtfPswrOjGZzXsLb3MLubMlrrjWb84SYWsHaFNbc4hIlff9u/nRu
+zheoeTDhzTvSNrvFInojHwkbLz/lnTn1HM0n6RL3qdXWhZ5Pc8S68Ma6yxmKplm
GD8dJtwRBGp6h5zAXyMNDHg0ZjZc3ggSScyApM8ejZ4Mv/lPlE8RCBao0fS4vqlw
vgS/tqXs3+eF34djXB6ywsZ9IKMUFT3zyMnVGSMHeQnE8HMBbry8e484U+/j+aU2
wOqaSTIDzt66ALXWuevorYhATXwAfxQqBp3p9CLfwfMhPJ7L4lRJBBw1dzKADlvZ
jQWpl4mD72KkYYy6shbnvWpA5pcSvVXsJXfvPpxggeag7w8rBbXZL/0tt0qLETj3
6Bn71e/C5vIIAM2Z5qsKcL76XQyFC3h7wS7CKSG+UWqdYVEwCI+bVMk1qeqe+AbM
BdWPQNHhJyYgLTYdIg1l+Wy/i0WbcnPqTuNLliI+a+3Z3lB5491791AZLqmoJdSY
tdd8TBvju9aaBnCH2VXsOaf/ck912wwswGtEXh7TFKe0CEnw1lPFts9RxT9EJyvA
YkDtMwAH0ACYm7YFGojqt7YHuzPm9UqiuZJYdClM6O+hVG1Apx7Y80C4qKOVBcsE
ZlqjQQ8NNJ4r3Dmkuh11fAoqpLfSkwtCjGQIZUinYFSL+TKFQ8RCS4HtExQ7XX4k
lmWenKpNjD3sEFxTmG+bwuiKADQ2jxGuMsbJve9AdkyHYQpHYDMHvxaaVGv2X13u
GvAdw8cMRRAiXbpmIBvVkmYPaFO0tQMAETJLOCEPm/SjugTVIZqitx99IdIUNR/J
IeDFsT4U1umOE7RvfWR1zMUndYcx5w3Ou6oFFuZf2zg6K1bcZa0m3TWyhk8Jp9Fo
rJyDqaHJo2IL92geXMpYCB4elW7FyhbwO9RWLaXUxtTtJ3EMDBOhHcfSW2LiEXng
wjxo9MJPQds+XgBJVS7p3qv7bNMMJW1ZewPPrDFm3sbq2ufWWcmDsMhssN1WYF4v
xzOYzxeIRDfFN1BuSBDigf+zHO3G8dzlGFj1aJyA4VPrJ2CRK/Epxx0O9VcWt0hO
TIELszE9ZfHMoW+DH1zNH27ETipY6ymhs5i4DnbGg39O0ihzlgQdg9yguWa/Hs8G
bYYVReSv0ayWa4i7n9JT+bxPNcOOuZQKv7l80LPdNzkIj1ESag8cuC4HWbPB9iHg
/xHZvYy09EpimpZTbaC/JyUyISKFdvQdai3YiHJnbY1UGQXADFEEvKYRjzeyqUpG
BJpxJ4IQJzuPLp0TdmGNF1w0tL+oYrKa6gvJD3W5UuSNMs5xxeIM1vUCHPbSwQKH
aE10goPuf5VsDWF17v9OOw/TBPX+sGKiFUFHvh0aRTZP+RHtWCM5WBebLUOVW0O8
sfnvMnR7g6BVSiqPKwtJg0zsBFIRTF5VLsZFdvjlJhaT5ku6bEYU8vxWAG4itJjU
dIFCRpYh2uYgCuUF78ojLWNhd6A3KpCQAg5FPcWXfnrgqNsAuBsz01KDfaim/QM/
/dT76P3zWZU2Os5cIrEvBfoWskkI+E8acFVtJc6hbBlDCxcaD1674gGrGjjSoWHi
XLAk7j2Dho2PkD9Uvm3gOF8GyrCCL1opFPooDieokAMh/Ma53UDqtz17atxhW9F1
VJyMFc5Oa3VoXbnt2jthuRYw/kfkb6Nvf7b5X/yDttSdoOka7u6cBJW9YWjb+B26
pJIn/h4TiiX+TWcs158BCWiFE3P1/w4gniysk0Ys9fEdsG4zz0FVdaXg2icVHzSE
mXPvS67EG6yLtQfzE7+0UoCfLOB7zyPdONRS1KIsy23kA7LYuR3zUxApfEdQbF/4
9KbaeUfbh2h/FbDPVarMtIu6cbbjovE+QMkKGX/ViNuQuZOhB1fcG+vxBM/pzn9a
lcbXLODWet2m7UZKt5WVxNEHhFT04/GqD2n0JMQ49F0eukB4uP5SXGxBdjm04P/L
3Rm+aJJtaUeuFFyCELdxk5p202yIpp6jN+RdoxC9q1mX5kAOvMGe8A9JZhCPtf+z
JtKLul3+WMMEpl2PmDIj4v4bc+PmR7SZ2Gdyj3Tkw6uM9BqC0n+TAyP2xLeCxmjm
b1wOaeS9alse1KaJXWwoCey6Zek6rD8Fvrqh0dfYJVQUrAG0iKzNDUNPosfcbAnI
LOAsUSHq4LAat7r8qtXAnvgFPa9CtyPdz2nXwFZoUfIOKpdcDZ4r6TlOj3ZKK3zY
HbPrqAWIWTzhdzN8rKP8le2CurGHvFUGq02GsMr6AndEL0bbQkxcXl3NNW6LUrgX
GxfKtQowTzNW0yKyfKGoSZEC+ygfYr4ZH1U+Er5CG0iZvmxh1HMJJcGQ/xltQCoG
eTMzZUayL0ZgDAyW7D+37wp1m6noyq+rCjpizmDFaNI+t5DMrBTpEDZP28rqPqtu
kFFabqjU4y3wp0wyqK+zLoqfN6kU/MX0xNdXwjBrxy/Wpi9fACc6MyGYNkTo/v9h
jeH1QAer67sk2CpuJ2uLnpHhDAcBTmwDzahs72u2ImAXNu0A05vZMFTRl31yeY+F
7GVOHjmci8buszYx8tWxUhEa41rza2QKDHvn4/ticdeaUegAV8avizbIyoUknVA2
DNwDFF3NjLTgwwfu7K1KCfrr4G3E42LhNwqsOfFYSSiVp7GKQNiw0LUambzRq6D1
/8+S86i8Uk3uQBercuqmb1ZDhzyL3imVBQFstpu+y43+YQd2mT3/1+u+mEz8Astz
q8RtfRz4DLw1coL/abOOHgmolsPb0xYO45Tn8dlY1qdXwH76rJeDJXZ2+/wZNXPF
sHW4ir2G70gKP3oC0GZWnLNuYAWrRZocbKvA6BAh+4cAyU32VFinm95R/N1+fX+p
YEs/hzNdTLtqq5ZmidwkWWD3XhxqW5ww9Yr7oa6AAkgI0Fl2JgxRzgtJmoswVZMj
N94iXLrw9w7r7HgXI/Npwm3oLLLmCHKR8AKFHhh2uHIWCvymjjPRzws70vHUtbX1
Ub/hBVACtLn1gbUAT+yRZlo9gI8TLuK+7VziTzjpZNXoucFt1/VmzrGDbvFROKcy
qf3GNPuEK/ErR9vyGUThU+oknybvdrDgYUOkoklv91xTgc6BnloJf4/iBRr362oC
QyNSZ671JKoXMw4HAYoFnInvJv0wLGdzQWw+ivlsdCz8A5ppqY6+aZrKKPePC3/6
7iRGF5+KVwgm2158x2hAVwNfw36YCqPNHJ3+Qjz5DrDvLkmeB82v9dttEPS2SXM3
2QeryU9LLrz6m6qzipKuy17+0yjjTnaQBmUuQFqYyVIYFNtWtdsGeyTv/WZyXJkV
CV66iMmTghMtA4a1twwdni1o0xo+Dwscpk9r0aaAx26CCeuy6lvXvYh7ieuxsEiZ
K5oozpnKjPhd0VpAZ473gH0YeH5slvfuFKlRQkzlceD1YulfUqUV0KoW3eeh/3gM
SrEv0y6hf2Cd+YilM/3ReTXsTv+CwN7M7l42xIwylcrGHiSl0IV3RKUG8AHKOdVK
Z/Os8Qg88+P6b4LRO+ct+yUzlEtWsriN2ycgCCoNYAh6jTokIwBt38QBDOPAaj3N
tCB90lO5sspL7vjQBx7aiebp8uVxLJhDvnBtJoavPD8x9Iy+yhqp6JcmleIqZjBU
a6i+YQ942nzZ/8wToZEgsLUNpr1FCZxC8OYXxf/UgZzPdo5aFlmhpDZaCtwwQ3NR
UrRwgNp+9/w1ciywQ3TWJIuoW7jVHqahir55ts+0eaDj8N2UB6hbNhukxxXJAKDc
zH3sV4mmrS/d+uFQu9Re2uSKutuJYEN9eNnIDAU1i+LGyge8NaIxiwdF01MAm1zd
7iHjpY+c/iiNmVYjFtzz7d3XTqmsRiBTOuxNU08hmgGnI/aAoHQEOsZvStFWy1do
hdtufawLVXsK9wKxllU1cTVtKZaOi5nqNUM+Ay3vp8TTb5vtCCWwZgZoU7OXT0Z/
VvVrqHDjLx0dTkX+3SkGG/j4PJTPzkLD+JPQnP8bZ1oLzj4hLnt6HeTiaC9Zorco
fzsfjcblJQ9gMpGWnmX1fa3VGSR9tfgnXrZmSFvkmWOh/TMdJzmRhsmH5dw3Qrqj
a2FMTDsvb6PmZC2c7ZqeqM5hYZJ4VJu7nN+TwS5wHh4PIq9Bqq1F0oEtDYIKM98t
wUPiZ/NG4YNqcq13XAy7jQkP0qlCG3rvF7SbO39f6Ajsvf/YQGAr43cVYbkXZWMd
IexXSBurdjpVZgymDGOjf5HAO+7DHLrVCcSruvjTP/qk00leGotdoDZRe6wxtR//
4xBTeY79lN8/IqZnqErAllSSkoiMHpJLvbfEZ+ZX0gVHnLnK3yxy6Gv/+vRutGJH
Q7jABPqpUfrrp50M94wsa6MXwC/UIEhzV0nw6DOC45GZ/EdVkoBQ+DclsAVDHTiG
wCzv6HUtvJYrsXPbXtIyhR4o5Z/19aySnhsxlo164f6xl3C3KMnd9EEe6Bodc6Dp
IbfUPTZ3N4Hxcw1yl2F7qn0HCMSQgYPqCxt5uwYrObm/dpdSwYc5+gb2IPILzJAu
+Ykr4LCm7Z58xfIuEd0osmdvX9keFYmy4ffGpxawXeHPf4H6LUJ0CHakQtvr0R+c
Ug3xWn88pmk0uh3CVYCuRrrJac3Tcimm+m+cXvi3nPXUx2iZcJGD0olV+NKbQ4BG
RGjHcsM2+uti1mKJ/Pn9BGHOuVNbw/yHMpRD6rihdWL4seUtSngljr0WakEbsUVR
HQ/bLl6sp4TtGbgX75XIGTforyY0VpxcL9NrTA6JelB+Jodcu8FRUVoZM6+t3Isr
pDyCnb0O2nMWzIB7QLAXa8EKrb1CC8khKmKaxSmz1qB3JdhleSHbtQfZfJhTqtL9
49bLuNSUXW/jlswab1UnXrlSGzJt1IhFD3egv2cK3LEVsa1GfGWW9vxPqn2/R8cb
Z7AarNmZjBn7YnI0OmrtP5Y6104ma5z2gjCY0Kn4LfOcE1YHBPGzE6o3sUP0oqgs
ZmVTa+BcTT3H3+z885i/a2kHlffLrEykaEWfLPdyUWlC1EBbXRWi1YEOyB6GyuVG
XZhDj507CFLv0BHpOMSoswMLi4ydneewHql5eT0JVikcltv41v9oDp4xPOP9Z820
UiIiWklyNO6OO/ElzSRBG3ptZ/lYD0z+7phRPX0paaqgcKCh0s9FqPlZXgi88pWB
pq2x+niO8q797gtbrysLh9JGF3nuE9mFPnk+L0HvZWpNchjdAsNrF0nUqs+hli09
9Nf7yCbzb4BiX71kxS5F7exq143S9e6i2lIzwCQrgMw7TaU7ZhW1+BGzSYOjPgxE
bmqzN0ydlljXt10XwztkFh4k/OQnbitf8cOpWITzXbUpfDiBCR3KYTZI+klslSLJ
wlHPb7YE/T63Ye5Irj0FYtyUfe+e+UwNt1N+tRF4NDK6uIlAndfirYWnEv1sTbns
NQHDPch8kXYjT8lewBFJvT525sS0Xvi4gVMjvMu3h7TKLHBmwx2wWuh0QVFezDTy
i7Ao1sNTILehaMEBQZQwLaweBypZ5BXL3F97V/C64EVHfDbVFEp1bYM6ZizCsMQJ
+M2uvdD1HMgHlTg/wt+Fahm+WMuj7rCwX237Shcu37iCjAji22589kg2xSam8LSF
9XAUGn9QoKcmFahJgmZ2jcHsHrbQ2XKGaJZEu0ts9Pxpa6R9DCmd8Gefiz00hchH
WuNVUOLXssiRzJHWCPUVWydfmi/NJuCWdns8bRBz7ANVmjzzQBpgPkIztB0g5N9G
q/bHqurq4Pn3KxaiH7b1Lx0UzYK/1lIF7Ogsm5sQqFGCI2VOV4stBkk582sB54KQ
BOXQB4SLAHnB/BQeUUWO+SPJxGLAwXyJgw6DeReU1+1ZU1rKpQZglC/I1WAJ1rA7
+hZHB01/psMtX2Y7D96PLLDgRJ2ZYKMUPRrog2fIvK8Gj7ZSoop4FzsQrOCVhXls
QRG4UzrAfEq4DHvsSYcarGiHzJGYFKqiD0mAxXsBsfg2N/DlbjwqbVdCuhtDDtif
pMBIeaolmWhpWzZhmxjdYIOVWxUw44s4TAGIBk02WZz6oTBULkApTGSDKZ9uor4E
ANLQQlORPTC6hgDFQEKnL/5fx7+cw+Awzheu4hkCEejbWhrDPgxWHzQg0jDEDfAx
msIVeMGUu5LPlujLKDvV0OCE5XeFR6L6qF2P0Nuj3lzfY9qVeq38LPy+1IxYTaBd
32uoiTvrD8dMDz3Vkd2MYwrdSXX/w8nFzTuoRuQoC8Qb3e1hfFNrBgihaBeBieK8
E+M+qbgBi3lv3oCZH0G9+6WKxUeiaJi+M/Y5MZAbMP/Bzv/ECxifl2KPkQ2+ZRS2
DZihzp6c/SCZ5aa0qCADqITnpY5s3NcWxMDmKnSkRrwQ0s6XtGR/HDm8IQD5iA6z
mvCmPrVKE4fb2HIhohkfaZF9XJVXKh6ulc1EjkuuHcAYCdn00kvMt5vXtUkyK2tn
eavtrJzX6L3ogGM0opBhHq8EwevU9Ps5D40KvHAULyMslRhue+4fYFZ3KJkMiAeJ
THKziBbwzF3wYtICOpZGfg2EzWXeHl30UeRvFYLsNQ7qjytV59hLi5NnGOtcf5mP
f5bw/2yHLR1FVCtD31fe4hLG6oX1Ik4S7xAVHqfNyDGLUGdlw2p+pgZcoLpfFW9A
2N0Q2+UAsCmWbstRPYAdR96/SUQv2vhWmsFNenx2mK6ZMMH/lMj6Lw0Exkub6NmN
lXWIt5nBCxPvGOGjgArYnjejqLdEIgeQjgeHyFgXck29e8LHndzWfZ/4C3p/4aYm
nOk9SkFfhLVNClN6EMiIm7fWcrK7B7JAQKvCWhGJaDsJyCCMwtvX2GdNBmo0YJYA
TKb8ei/240zxrmpOzqVh+0wYz0AEnR2D18kVqgnwYJU/jcjQwzje9IDaVBm0Xj6K
MsEs29VEiCXVj+hLdiTIXw53t0H7lBS5US9miAK2EAxRg6ivdVTZflLXONgAeOw8
FZtlOYldE36OwdJWFrspJG0KTc5aIkJlOY0Mgt8Rcr9qrikewnnJU74LfF9An7vv
YopiGMvMePIu1Y3hnQ78k0kgYkBJfLBYHsNpiLGiAspFK5MrpXf8FaL6WfoVWS0M
M2VQxO9RhnArcxUHSLstYyGpJUnGTw/umVsU60QSalwSqFaVGRa7VNVdau+rlg8T
TQ69n4lO4HcuIZTwdwXWEaVdpXLBK9fasP19o1v1SNFA5s32fjADfYyDsCEHeNgv
URAOKsQ3gkaMTSlwJWqpGazNM1TBiihcAHy1bZE3ZQdPxRv0wk/ymyHOzE2gEtTx
1WE7crudzMnwPbMbm0sXaa2hi/S+pX3a+Ht2JLitbDETFUdU8uIZWwbbcIQeJgiV
sqHu9utAkaOh6jTDNLUzfpJH5DleskJuaoRTz8JofJRr7fBlpUfMJYy7acs0Ryyi
Dem4pguzFmGPLoaGsdH1sZDTRESqB5h7nF71aenYqbthmgw5jNUlRTXk1iKO2l+y
N3jjzeR0Pkq0I9V7WharBYWRmaNGkd8+UzP/r79wbxXRwOp0r3QyihaKt7aJbQno
QR7aCaeF2+y7+U51/DcaLeGLwycxPc521kQx9aHjnWWU0aghF72KbM4qhMGz22RV
RQO6cxA/vQ8MMWWXD4kAqoX3R6TIkPTpD147MlqW6u0yJrBYANdq0uQMs+TalhJS
dqJQuq2tgrecmN9zq6yMNqlDrDGiFOd/9UYJQns64J6Ly/dA54EYNyvctcSMP4q5
LXP8TQpLL51NDIYHaUt0wMncx/w/K2ipX4Jj46ppBU9KS1a8A24IG1psFLrhF8nj
Pk3jzdHE9pyl7Qv/KYVV/PSYhsaiDX6t/Vbyc32/d+AvButNy1ERvJ2H6baQU0FR
gsbJiFdg5UssWuXmaTTpKD5kyYgbYpt1RPmybxdQgP1Ac59eTM1WCRGP31y316iE
71OF/6hu0D0+Pq0ah9yc+TTLXnUpcn3lBp1W1R2D+exxbcJV1O5Ls0H7YDZgIgBa
JUx5B589U9LllaZTa6wVf37McAADXLKxRuX6ewbYG6yJCP8tRVLdywmMlGRfWa3/
/q6I9QLNo1xt7IZJorVB/DhNNxcwpd+oO6/HOJf0kklVrKuHEHCDx8kcbQCkywF1
2Rk29ODN6fRgUXflzkcA0kfHqIV75s5NwILNywM1iafiy3H8nkZFdCBo+Xg7WEyX
xDFyuso0Fox1qegSvCrGAqAnbCPodMCbOX/63YUpHPOzOCTP6rQJIMuzoFEH5LKK
EQv20yQLegyL2qa7HTzA6meAEmggFbqTf+vPZmF5ic1X5AcsjyW6nmVLCvVpeKFV
MZehmBX7jevdbMaF75X3VRXBDEBqzfiocfXEK4qan3FcjRbQi/dn6QcqmhLMNSIv
8XuURjHB4p+l0HEn4SigK4t6ugkbspc2PCZmxSCR8nGRSjcYkD9cOyl4tqgRwMnr
uX9A0tk0VedOGyJIXqZfk2aoyrOat6TSCkebkT1p0Og9GDYXO+x62nSHcn2zavIv
c6UWeWEHTpH06VwMqakIxF+B9xFAHqET8Tw9aFefGDIV2e90FUsuWfRhGf3ICfnV
AAgSd7FCwFVl1XcrXfVhGZEP9If/AcfL+ZLvjcM6ECEc2pZRh7IkoQTKs3J+qFDY
aqEZyIp8zUFloDvGEqNhOPWE1A0zCxAm17bZ52rsAx7ZbMcXuP6jlnk8B6PEnkwV
5CiPZpk0ZjYNTkiE0KfaXLS7G2MZPSV1agFliYuB5RSXtNRYNsL/iT7ULGpF/rik
ROMzfPQ2SFF0cN8SPqd5Eh7nmgEBy4bwefpLlL3g8CL/v/+BltRWCGtWVJdW7vB2
f8xU858EMi3WbsUbhJlUm83MOSJd1qLIL0Rap8GBDPkYKidtCtciHjzlZfaDQ8UW
h7uyJxrpzK/ANFtUOBOag23oZr9Xi4ojizbTihben4AP+BOh4JOM37UyNTvLGjOp
FfRse05tAajZj0SZi8FHEwLtuQi59sMwbgCEtYA/sR8npLr5WHRlYoxOEWCPGxHR
mwehEoVW0dPO46fTNwkzPqKx0RzlVU2cqP0/2vAUuh1O+Wn6Yn4rXUYDzhU/1jHq
J9S9a/x00ceCzFqg4gubWSKG9hBZac3STM7CcyJF4UvfcNwKkGOlxCunzKXPOG2r
aPN+nYGY+BbKmfUxhD3GHvZL0FGIzx4iJxye0KTI019vCvr+J7VbdA0K1Ki7wP+1
ns/emv0qVeRn6OW8FlBRDXLAHl9Caosudw66cnkcKGXt1RCznHj8KTcuEix+jq9D
rtEa/4i9/QWJ8JXsCDTWP0E5gb6tU3WptakvmrXv5efisHV5UC5Lbz9ci/otZ0rj
UhWJUacpekv0G2t5i7THknbpmGAEpvwjmuUF3+cZLyGFn481ygZyNABY4jzvfcq7
UHmGWX8x7lmIGmM2umUo3J7Hb2+jBcxxTfUVwAoKti1Ek6i+zOdsTyrHNZ2jkvAt
fp9E23UevcQjM06mEqa4oJv8ImiU/B/KFYgubfpPre7ucTimLOwUnbQ4NtKxbIPC
sEptMElk6gVKnHOFis0U/qkhzjMTUfTTGI4kO9/xEQBoR97+g2nPIteaW727vnIa
szkjZfcJcVOGnwfSOvkbE+t3EmZiBtrfflvRQYUxDCHbnZG2fkhOKVEXsCDiMysA
ey61y4I+ZtEoJlvNJa/fr/RAWvyd4UDT2d0mfS5XY8OENktiNh39Lhf3pOCuqNiZ
KRRAHxIRrbo7ZpIPnLD3oHRnG/e1ZDle1ZOBbGWJGM/jYr7qD8Hsrb9J8TT9A84O
LvLN5aIjBJ5t0yPUJFcZ1SSSv6S5EMX/w8uWs8AHxg944qXpg2f9OjKjHc0+pOl4
ON7L2+wEoGZxgD/8Itgxyp30tkt0qBDh7DsW4ELNvOId83JU6LD2TCMjZ4xeWH7F
v88pEn9hVKwECmBhts7ey24MCY0ZXQ7EQ2qWdbSNN/Jik2InER/E/he5XSPF8Y4V
rXdF7Vn/JZu6OS1x7lH6hYL/4egp1wbltvhvsjCJZjXdifSpdaVk6iBFNDvy34KF
8ObhIZV2qxUDZ/r4LEBVFNyrDuMWcV7NCIR4u0+j7EQcUsdoOdv2rgw2ODYFBu99
FnMr+rpW72T4h347aBCbZnucV1lmLQu7g7Ckne9ZPx5PxnxcCtrEhdAdRtqocDGc
szt+IhgT0gTP+ySMOy08e0PT57f9om8G3yVvvpFku6nbPuCdwZb7EUBj8olefeMF
2iW+sLYpEduXvYQjt3dJ0+InnzB8Q9HY0AJTuPeMl88QWr9EKZK4zyhEqTPvh2J0
IAHAMvY3Sod5FXlz/FeHMVjC5HoHv+OzYTlZ2+N+057FMiYBFmyNZ7LA9RmY8cwv
QxNVaf/kgmSvyuWP0bPohNfv0MHsLtcs2v92AcTqMOzyPq7ZDpD4pkDLbVj85rJ4
+l3xAumqkV6c9dytNAVkQhhPNz4WT/l1JLlZXddZ6nC53NA7X5E9j32pFoIpKYUG
utUn2lQxoFihB5qwHqzRbL2cNB4BLkFvIhtizL+XiioD+9cvGN47lR8hMluGCBsH
2kBzN/qNVuZCPMSgNiGg0yeWoyDc28tyFq4t05jwEuBCgZhQhuV66cHWCDouEk0V
XtFM8FjnkvoZImwi9x/aRrHZGgW41E6JHmkAgtMFWncenriVxI4gjzug+GrX/V6r
R3+qxUJLpIGqpAVsG8CMGKuN6W3b8N6vlMZnQBpOuWC8ifW7+ED0ugf/ne+tiGzJ
ltQxLlhnvX1xU0KJqbgL23U4qDho+LnrEyuVoOA+5L6Fr/QBPDYeP+YJ89bqzOlk
4yVGaUKwzOzn7tn2QCDz429lkfq2gQMN83OgsNqsUlrxdkDcV5aSD+vwbGnE5kp0
B2+dkxYNuq+w0PZlgaCwTurLdiuzuufm9XiwC2EzRbSfghYnNMz7PsXNyMMGn2UD
e+nt3gnIQIg52y/8PniRtMd72+XlRdjT3LLnXMdM4hxjC809cHI0ikZurxZusJxc
bhEgFLa/9eLcz2pd+Bz35Sq+boffD1nxFrLogIa1oX7JGxV0MHaJ3ndK4EJANyxL
374YXigLw4uqnDDYszR8QNJRgWxwcghvm0QB3zfoOfNlM4bI2axuZq6lsVEnOaYg
7N4enAp3nC/AhxDKfxVOesoN3QyB4yTFUOuGCuZfttSnSzfPPVOxug2wfZCS7MJP
AAvsJ/8t8vaafPEUQVHwMSmsqagEqzrHpkXyoBG0Xr5VUGCyb7s/bMmNrH9LicfB
EVObolEhBJCe3agZxaHyk4r8kDY9iesXm0sCZ3uXBu4aGpSAWiccqFXX8GHRm6rG
Aet8LHSqzHcM5tJ8frfAUapCYgaUAIo/iUQcslk7GUUzP49HxpOlXYYeM13rS2fR
eGmQdmaSt9hECSZhBc38szNcXiQWifxGHIdCchsZ0g1elZMBbCxusvhW98kJ0cp/
75YKeLMYhdOCKBTbeVACQI648nVg+jdqcckJb+CS3xYBUbLsLBH2u5e7jqUp6oOk
FnRGpv/5Y7eLymPgDeRtT/Nubm5/IKrfzsWP8gNEN616aakvibh26AnAZ2OB+Lbl
M5g7e3FnOB6W4LkFjp8ZzOgCYG05dCDyIcKGk/K6LFydyqfXFRzlY1nzP5PgpUS9
bIsO43Euaj6v9Ochry9hAIdL3B8TPJM5JhRpX7K9ztwWJsPkx2gnjqDVxFke5lZy
eKGFbZFXS1c6OsImGv26ivAOLkzrHZ63iwSmB4NnM2Y+IGZ8wO1REhAxDtvqmHJm
Ui7nO38jx6vEAyG0kyqiku1WQKdfsUnS3UlaacGaKjBymfV7nLcVwXG++wtfmRSv
Ef0AlPyiefsp3ThUC9BqESS8osnDbJIVTDiRhdVWZfAvlPUS4bX/fCNAOG5dmtf6
q3E7gtBUHS6F18aBX3YqU/3AvCPIcU3cNBBAmDAnUKTZF70KzNApSXN2D2qAigM7
cSH4BMCA8QhdES7rSPpuv414fQxh3IOQlH2/y+OtUujDjUhWyBdn8/q2hITWj7Pu
tR6l5LPc4nsaRDGAlsgka6N6U7p19GWhjU6hg6n8dE/OzV7tvjzldMGYnks0okmb
RVlTMh9S+vuLz10N/XJJyrHW4Fjgd6UPuThC1I7FgP4FGhPEtTeRDsArRoOXo+GA
xZXVcHWfP38G2KiosLKtm+YZwswW5vDw9NRQ298bm8MMjrqJHoss6MkTWNKbEDgo
fwoVVkyyALeGzSh8x8PBnBsBLyle2d0tOifRNzuxDqvVmOy64zqfhstUlKstYyIC
bJRkEFoGDXYs5jjm5pkRkkRgsQ+TcSrQJ+mb5VAkhCxvtbFZvMMjAs1ManAb/bLW
djaahr014UaHYAL5odXbfdfaRyVr0HylxJ4fRhyx/ZF8UR2dqsLchX+/qRqBLdug
GJthmhWMbFbM2bj+IDdgb9OQSh6Wrq8KAy9bgjbHJAXrQffmJd9f88qjExjHht5j
XmQ71C61Y4n9HjOby1gEtU3Wn26S/eEKoE1665OMpVEdkBfBwd970r5ut7gsXmX/
r8IgOR7oK2Ppb92+UVi5Ulb3zVS5SFAZS2/sosYJRfK0cFnOawpqFemgKFKVfEiT
fUU8pLYE6GIdO+5K0W4szaifMuAH8+9GSnpzw+d0UDE+xslSVrPsLRPn8tRBn644
xr9aIH/qdKIumXPjGRM1Ep3g57k7OxLARXq+QbEbRqIvkwCOr/mN0V/2K7393CMo
PONK+EVMRzuoM78yb+oTBvMwo4KZFblNtPTdRRLwZB5HW87kPJSJPwCXfXTKkRaA
H+8FqvoNKJkinvsKYaKJyDSHTSOoXiQaaOhmtktgwxskrHx4dPB/DEfRBYMs2QZe
Wm/bCz55lvdefCRQSgwUCFKuCq+bTJQdYrn8Ews7EHFU3qq33dpdAMjT4WRU65MW
pQFSzssWsPblHTslvcuouOmczXCbVIrK4vc0hPYvpwLMPuUJ8oN3wEoWob9VrOF0
KYidJCi3Tyh5PuFMmnsKJpSu31r6lfjt55SYS2nLekalojTCM3HdQ8Q7gd456KBZ
LTqGrplSDxkOHPNJpMW9oAF92jIqBKOfhMgnBnxsXu2Ho/c8KLmA9eBvSaQHXQcc
bqCtjtC/upg5d3UpuWTCOmDU+F6B+2BrdlZpL9Zva3hq4/BOTC/ovTPFTISGVYb5
mYTK28tj8ZWzwevAml3b2N4sQV4Zc0qaq3rTBTnA509lQ7jHXRp7LCT36azhjOMG
/ogzUcxJL2Z/PQz0BMgMEpTUTC2e+0ItlL2TdcrZiFGkdHmqsZxq8SHg+SqU+fBw
arW20IrRG8Taxyo+wsWURQxHgZWLS0acCBWySEq61FxaoZ8VbGwmrTbAHvTZyO6n
FHzszX31CpkDnysNegcqbylosObUhM+e6w94pP6wJUxs+/FlLx/ZHOafFqnsDc7o
3UTfolp3D1f1lTs0K/rexr5w29Wffoqrlu+KOtHDf0h62aRcBxEvunGrUVvfbJ2X
86g9nZiUoBCQ/qyZjDYEQ3RjmzUSmYPFRrKWzYJ4nhBTNmoLPKMywgq743whJv6/
ipoa0KQwAI9hYbE/FVrzO66ScfBM8Su9Uaen76uLON9DIQU4YEqyUqA8otteouL9
JYR10rRu3kDYB+rMw4C4QtNSm38+buO/sA4ECd0Lh8RtW/RTZEOf6DjW9t33L4aK
1MSgLqroI6IyxvAHK54iYvISl4L7q+wixgSW0ICHuJ7e+T25KvOHpjiQQ9vB8VBA
MoWRG+0G1VHvc+hlbndjYgp/flr1bHqYaShwEZa0/R9PjhjL38oRQVBqU5ahjJB/
0mM4J0U45oNHZgO1eOxSf3XRkZd6qg/68TbcomXbdp8WC8t6urPP+Kxyb77DcBZS
g5C0KXIDAHayfHhJX1Vv8BI9OMGUyJUKfLG2uTcXsA4s2wQU5yagow21cFQ0fBUy
sDJvK00usECXL9ATmmNermeXLcmaKymzz5QBzpgA0P41XaBIP9UlvpFtJQ0LBHA6
WMqF5JJpGD4wS5uzI9NmQmf+8qOFacsXjVWBgS1mT/5M2BZDyoqQtHG+N522DM3j
NsIKtDNWQs7dMkGUepy9VZBJJlbn0mUN5rmr/tjLTVO1rXfGKx5JojXIEyhtNezg
ha538tv8lQLKwh4AJCC0AuFir28S3FOjzUPkMGTlTj68v11VGsieLKD+JwNpGUju
O63Go2BVHFVsH2stRz8yf2nxO1H8VZg2fCcadVdCldknNxjdr/2sNUl+W/NQC9bQ
V1dN5KNsFl/597DwAA04y16lawspan7IRA875P5y76EKrXeUe3oGx+fqoVlrkA8I
T5ynauUX2Gtfe87pzOJZ1gsC9XstRsxjm8b9akNFVkbHfwRMBwSaVO22RIy31g+m
dFqWFY+7Z9yVedVyX+048DPEJUp95giN/VO3epOH6nmMMdFuUGL9L+Vql4qiqNDV
HcTni56Alw9Pah6VxT10W7ln5lyUFg0OnOI3pJqBIR2OYR/ulf/twLWch1nM/hIS
Lxf9hWEVZMfr+YnHbkD9pK9lIzcWY4OqFeF8+BO5JUBiIepUa+uax2AvyP1eAUwY
uN4OSoEywiMMQWk2/GJrte19ccGcTwBQ6cmYBXibo/6F/c07N1buDK862qjX0d82
4YP5pSI+C5B+e6UHJwiL6Ghhg1MxxjRb+MPj7zLvkQ9EHQzhz8Zm1aNHiKGLvAMP
J06Ow+3Eg0YafzhqbCWeucltgZfB9REvSRN09gWgOJ1aNjcy3f3Jl2lDqxPXSO3k
He60gTjF4uifl3GgNLiNoEIWqHVTL9Q7rRAV2tpx6x6zFFPUq8sHROIvFLwrxi84
e8T1cRGU/4WTBch0hEh/pGZzZ5JQotyRDehT5UuMnDf50/XDDxOY1xIIo+Mfjk+6
BHSf10YSTRsJul2fmz+VOJV8RQOLCAsh/RYp+5+Dt/tDaJlWg0BGncHVpZzvh1hR
FsGile0z4t7pzElXLRhNfj6bzHBXO2CiAbGITxFu8aQtrRfaP8k0rTy1H5D68g4r
79ktQqGuFaHeYozwjwcVt38riShJRFczf4z0BmJG6mqRmAVs8xlSJ8QK/TBGUZ8C
ZVhMCHj115ng0q/IHMIEKP3ej9MWvZT8Ve4BOEPqOthkv7A8D0zcihplqdySA/KZ
dEsasKbcebIb2HilxnoB84iNAxxebKrrb8X9v9wktUU4prW8sM1dN7N0KffBcZdg
ml3ZqrWNaByHllfTeOV9KFKwJds+lFM7WHEPMJmUDc5f9WXMPnDEORI0hGL0uE3Q
ePzWiZoGXdkx4TkDnt3tWQAUAz7yRn9KtHop94M22Dv4ya8Isb6sGBJTvr5Awi2P
lA9W43QPj5yhr6sGjVwsM6ARDiUqVCFizXbjTbzrlVLbC3mlOhkPlGOFd3UuApah
/iB2p33XoYBv12wdnZ/1j65C6UaaV4iY3Q63ry2vjcAT8BxFMSbUBz1H895/F5x+
OL8mcXVOE+WTAdFrdPOFkiK2ysn2Yl5uD95k94IwTLjcqQFOYeQsRAqbmrEaqQHz
/uwbFiVYan3sDHkYtOj6oWQVR2iQhaBznNhhMPuT4Ypq0LRlUCjE6PaOaV+ZUY4J
ubK4MPmNNz8+49JZgDaSiuSrv6eDvGR/4bHx+YX2tWE5cMR8PvEUIcgOfHehXI/o
rS+EW/uaQmLVPUJT1z7WBaEggzbqF+MsEyvncO/U2KF0hUpmKU6en4PU0FgxD0My
DTqyWXgtnXx/n0/ac/MTM0ml3ku+CRPLpNvONes6CaSuULSMTRxGqHTfcyFtnfD9
GDHbpldLhAojf+kXykIoE4K8mkEZ4z3mUEdE74IpK5V8gELOvWg6i+YNqnz2NOX8
b6ze2QPvx+kHRu7XxNffVwkd7JVM1K3pRc4SKPrlmcHHc0njENGBttGdBMY13VpK
AuI9gj+BkXsOBb7S1yvGH+27BBbwsomF1sjH8UKAAEwf0TK2ypg8hZok9TwcB8gw
nTINxFIODoxShWfRFust4SD+I3jId6VeklPSKKvDvVbusAovGaiQ/4dxzJ+UXifh
cpnAmO107V5UNlmf/4Sh4VvqyG+oaHrtrlsmI/LsxtrJ8SRM1d7RkVKe9hzmo4OL
FE9Vk8PyIFlQ0qK9vHw3+T/ICKU06EATRk27ewu6aa0/9z3UsJka2urMcDoISmn7
cwGvK0PxGqQc/bID5anC4/S7b5aiD1RL5LNv3HwCTCqQzCigq0wH4umcROCfma0+
iNJJthcUpzabm0BfApVFNNTzL6UB/T7Th76SaJWRfKqFIWOnMk09SQgraieAo9YN
ZooqmDLV5HdkRF7+hOkAZMML+2jeUCJBmBYKfsGfNXwkByRtRQnzA8mbL0Fr5Bwz
iOGM2BZCnHvG5g/X+Me+uwGiBhxk4aF2cAAF8i83ZTbYgdNDM51wkY33xHIOqH2z
OcerCnfyIpE40YChz/SyhlyN77vDWE/hGIt2B/Dq4GOqcRoNFCAthtSsTh967UZZ
HE6Ytw1JXKTniCYNMm2IasN+LqLRRs3fqPWcHk/kFh3gJNxtTU3g+R27OyFcLQiN
7zjHO/Rc34XFdm7jvq+soFFssfSBuX9mupm4T6D+/WKBEPmdSXpkbPWIm9fZNzHH
R0h+ZqJJ1VBZqswjxTrjmvDmsCQcUgufQSNMGqc4MVbIVCHKRrlAix8blV2S1Ngy
w4V6B/XmVUH/4UN7X/eGxPSBEP8cuyYIwPI7Je7H2nTslzW3ZBD7LEzgHNy4ZRV/
jLP4vCK7/+xckXQ+yveGjSjVY4c/hr7BIHI38/KV6Ww6RAY2/tg6no9bk0izYHSJ
hHyoIk68J5jZ94y8K7YaJ+Quvh17weo8DUuHPBFEzdINS/NX52WXhXojtm0ddvNe
fY2ZUi46BR/2RDbxuPktO9/vqRVwm6a7euBndqVro6jxdcsk/fL1n46l0/cmxGvw
9xCTxOFwHMduawBovbafE+oNtUIIC8/T+S3wLN1jHY/zX/EBZOOXbJHf9zJNAwfT
7NsGSEEt/tfwG8rDCSGx8w3ly0GwGdHAYWBNtb11tlEEgwQBti9bnk1QClImOpKZ
pEEmKQkET0phcBn3p/cQAq7WjUHmZpICi+CspG9uAE11JctZgXE/VFSPyFjRwXKH
dNHvBAhot/7JDjzgsLYGG6PSFgJM5odmbPj5T9xH3rc66yJOti6qK3fmqgCAaMNJ
rOKhRHcd5+dkHCLr9ycyahDtvxd99PYp1Z9Jj8XgYUAnQ9va/ZtoCgJtZ/r5OOKV
I66mYQnipG+pC/3VGTgd5oByqPHGTOF1Ik1EZoQ64dIqZYlkBmU4+HirahjnmEHj
s/wpLCH3UiVzNiMYP2l1oC2jFD9/vVBd5jfdOuq3ERSFOq3XXkXWY/LmfK7yj1xS
eTBgiR69gXTek0iS+wDUZIOAT/0MwwZTotE6rO+7KvhU/RARMnR2VhNMQdCB1etQ
lE3mEx2jjDtFQoNIRXlR5PBTbZOFvF2UQhzK6KkhSTSW68mQgdjkoUGHNGvIM14v
Qstyelk3MSyaNtNRQU/95AYCq1J8Br9+dJWx6UDOSUpiZV26HWu9INSeb4m3O0Yq
VvI4QWVm3I7z24djPq2pv5fKSGZqcLl4fIUowa4eXS2/1pTVr79cuKCDB9J4TGJx
+c0TNWNaGjZlDcm3PRDC/P+KHssm34Y5PhJ5J08ppcWuEZfRNd9SogVbtQYw2Xw/
iMCl+tUgVGZK+KlSwhin9xAB8cKUjcm1gP3oTLp4HtqRJql8m2EhuFiLCBlZsuCW
290QFbF4Vlzej/AFna8/7rIEgBT1R1b4Ney3QTu8gDK0/6LK9WjFWFvyRKetp3pM
lQo3wdXofGjFd5GFHBt2NtjoBYYAln2i+hTPK/hnS8lc22CJPynA8tUb3yOpvAc8
awLRtRDjdyZ43/STnnkAXZPZ6VSGb5Pd4JqXGNRqK4oFvlAU1GI3rkJssuuVPBXi
sIo6yZ3moHYD73r3D/7dQ2d2ThWPO/4SAkdipnMZdVs+Lx4g09URTnYJIvmUL9wF
ME9AmrSnE/xemQl5ei5pe405mMtVO4RIMj6DUFuMa4Z6zNs9TVkHm7l8iXD121me
BTE5jXUneI812uq9mLSq2R151fxAX/QG7n+EuQxXlSsBcf75SsSHd86DvBloyLmb
Z7INHEIBnJxyPf1rvO9bzU+sbr6f4rRgdGiJAcbYOz3EwZlkBrM83k0Mp62GUnt0
FoalGcYAnAU3kec6NUBLRsfs1gyuqPHDLYgXRPSRUjz3Ej+9SZ9bhSE6TYub+MDz
h12r3+nmHuqfPZVnHL6zBzvwny1+mt1sVjmgVPGTUfuFKXh97SCtRdJmExxCJemR
EfU9k4CxzVATZJn6msWw3Z06dfN+lAlQcljFivWQHDW/DfdhbKLARL/0Op5vETgd
zgnjUSxqoWDxcwYoon/yBVTIix6JcH3CHrdJstvj2U49K6fNjgo61tng77FdVXnf
OYAxDBay03x71iQDgQpcerSIKrp7cofxhqz1vaDdTHZUiBEUvIiUBTBBkv399qkM
i18NMUr9RSgNq5hkwo+8gkCb0zBVU+V0lHZ7n8Gjpq5GeEku7otnTYEDesOmePXb
2nEYEtYV0wak8K1A1NP20B5Q4RPPwpC0sBvqN8k/lvJRG+2AqH6zN958vQX35zif
gHVQGrYYAbL+58Oql4rggqaypYp9bTfZhdtophnEroBsoSdKNdZOHUqXDnt7XD2k
IkDrRLQZuo7vCeulam4gSdJKquHdNvVwEzIlRj+aldFGs7RFaxVfFSikvvsIewAd
ab6TLYdiSjfEJSlOMzCDT+Ukfz84V+cFY2VbKLZ9nTP6p5f55Mge67S0HVJrXey2
VepR50XIm7kuSSOBtN0nhNWhpoWPihxj064JLjmWS8GyzKjipir3X1hAjpKlnmfZ
GkRhOaUzyuQEI5hr/+Jv07PMcpfEXGfyLMB+f1V4yHUAV7R4Yeuti0KZF6XBjIt3
ge1pYpo5x3xR6ZPJuzNWGKkZl+9n5mwRp5JYabRHdv0b5CjDORPzmc75AqMKQm9D
w2pkF3pNn0hMIeNoFHGsmc87jz5oFKyECQ0AHUl2vj/Hno//QH9609QhVNiuf4qK
feUEVnLXu4GDa6sayFTsIDGCwWGFqdSUQq8u/1zxRz1Bno+w3vl7IAmNrQTm4/0k
fOJyWu8wP1Q2mJDrNQe1zvfxKCh+IiUECiGGHaPiQ7oBzU6Q5eSFbk325bd4moEV
0NY8+z2lDTO5klv2vPlOsT+SZWcampb/UPB82t+zCcKYsy1d5kE77Ut52Xz47+4B
OSb0vJGRUAu/VO8GMVRg+Bh1eLy7TMQUNFOeSmslVXr94nnPCrzOqKnQsJptqdE3
jw3Pv5qzUgmTc1hZwdVWXCXE0Ft5F44DflPzJa6Ynt740uBuFiMq8NND/2gMHAKr
DKkwl6dVHUK31lywRf5Xk8iNtgzXvy6YeVBQu+4W8E/G/lGDcYuZNPJayIVF6xRK
D44h5jJ4cBoU1jd7rqG0TeERIurKV+QUKUSmJwfmHRpZfM4/koytTWIK+QSaX7Rn
4srV17fyON2nzk5HB7LvqZwceTnulYLg28EXAGGG+leOmxGZoHuADnK8L+6BvTce
4/5SU3I0RkDnZhHw/w5NnZvlUkPtOYmF6E5r91VNAG9mC03HqhpzkYVeC3UWDvGw
/ksNYklTziMqOyMHZ1eO2pg395d/yUtaAwyUZjo3Tl0WctqL/50XGPl0CAgiM+w8
xW9dR/7SOVNpD6U1kP5IaA5F5rdPF2+5eQde7xYgxHC3+wqhAHDUzylTTvmkwOVC
KY4BgcTEBqJu1ItweIg9x5PW5ve8R4D1zvssTc5vjvSq7vKbnRtIulouro3EA26P
++7Hse0F/hgzvR7ahiJ8G572j4xpdo4LNUtk2tH/IQ6cqK/7YFXLedqd4nPjxKh7
Ex7Sy+hZNNvoGW4IVSj2zHudUZ0ligXi7vJlg4SBqjgOnD8+/7Js/V/kmBRo6QCX
ttRC8kZP8xhZFrhYtITybltZnFRkOC3e9NWDtM5qEsMhuaz7JIXxkz7J5P5meM8E
err3ucA9OOMPYUEgjsOVL0wCB/Wzi+xY21EMMENh+lKbuXSOEUwwYFxfy63nIUQC
97gvktkKuQaLTmeeljBfl2t4yEotoPX0ZHOpvCdIoCCbXwdNLKMYPv4c87G7e1Qw
SUB+X4H5/Fv2F8PCM3Q0drFVRgLfX9RdvBpEaNxFYo0jMvmcTZzrRBZNZa2Fc0Fo
pE/l1zcic/sHj9XE0eRLvLQSo4EozOzy8qu0aBkmEfAf5ZU9ZxP/S3aCmM5Odup6
F05H3XDVmoU580DjXNldBJ9tAnCaDTUkz8G7vBjsgXSUAR93bu1EpXsIYmeIP9GT
lYNwu4rOEm4mZCOii+pEEKGMkYggsYY6TqCoE9aVktvtNQq6kN7EbQWIJEfZEx0M
0g1t6mObE4d3F7kroJO5/4L1qoalOhlwok2v0yxCB2Q6cetszbl0LCv8dxwvYahv
52ey78LRe9A7ZBg+MgTuYUepSKftuD/1Rqr8egOJ5W6JrJeOQI667K4Uh51b2AuL
EcbxQbJuU21RHxhLYYgsKV924ztu9WJn9bq/9ZXiJNsOeKVQ9b73NzQznt68wK7b
NoQuBEG3ujgQQkU0hAlc0CATfrykwnsA9R4P6dmzdR3q4SJGIELYy/y1DBgjWdlx
Y1vJXt9i/VH4qFaGE2787UMg+GxyttXc5d/mf7F/i00DBL9p/jNHCF0guBUpaIto
n5j+suQDyfU8M9V1Kv6MlXAVP1R6s1i+y4RVNBLecoNRI543Qjf7kqnnNX2kHn/1
HrqoPJo41GS42HLOx1hlllFeIanD7Q9wOR1iuyOKyu22FTWFBilbOewDt75zNws8
nOyInrVz20P9Mfz+NXOG+QwSECVDafHYjtoTwuQnEer1RTmPygEcURTM7iTp9wjk
zBZPTPVE5IqGoxYAGgDmbVxOmmXNt1L32gyyXkmhwsqzRPZphHyDL2cPr9xalVtv
7HCbXi/6NwxgPhYyLomu1gyItiLdxKLmgu/s4m2rVRIfunTr0+jJW0Nc9DsnaId8
OKq5lcBPCikK9LpaU5ZYJpnZr8QSEWVbpiG4m9m6Pr+0R52j+B7Ibk8jXWoE1jrt
tV68iQ7KBhAOyKXUmp57dyslbqfW3EX78kBK/Upl7yiOdyEvKpkAV9AZ9kz+Scnf
5fk80o50iSW5TpcIs6xtzjSNGN75ywfnOZS20xYtKzk8kNrvbgzOR0jNASmkv+fR
bs0AKnepSq/ONofcvLwqm2TotcQ8NnKk94V8HR75RyysVAsteu8Z7PjAANFdt1Qi
12IKM7EjxLFzzSeSLuv63nqFISabOoPxHfnozbdYq35UWNpFg2hQQyONpp7q4KqZ
6xeDhoUTHhaG46bMeV+c9H/Qs5sy7k0IptaJdQZocZiFXUOJhisu9Zwdp3ReNts5
jPl7e05W2Rw3rMG1uzxYUQ2RfFwWfM0pH9oqdjuht1+wHp22LrqUZ7iXtKrBrEce
7okLL1mpZN2yxcg4ijyg8kwW8pe475LmahRXOd8b0wI0joSLpBbxAulnn4lDArft
NwHR7TaodW0b3uK3kSqxIj/JKuFdm4JGd52j3+CUhOuH2Cz99QKI9XSUo87G9OQl
7VP8nAEJ75CimSusYrgGHYbJQgAmWz4Xpot9Wm5IMOAxnybGl5pq9YwGhST38Zze
JnbnJ6MlU4zpSGbMgOrSk6jGa7OfGHpeu0il7F/L3ADmZY4fnR2AX0Itj/CTGOu1
pFLDyAxizILhLU0pmIi1FKa/k0gj5hq7v5X/B42rcBztbDllBXyEb5A/l64WhLD9
xYQKVICjev1SIcnuwL6y99wm9CbefEYyeT8LzvgzVny4NJuOmUuWVt9arm5wWY+N
KTetf/nYTJ2BaZHrDZVuIUdA1i209ab70zEAWV49XO8+5u2IMOWFYkmouXwc2w6j
lQMPws+VxLCUmfaAl7miTVkmB1EmSKtbk9UY/6q0gCl554+x6wcj4GZqjMfcZF1Y
PaW3osccX/al47jmLdJLqjQ9bQ03bUqmRFjENqE9BaXdqg8tdYkdoYCcR3ehXKNN
GUJV8T1AorpRHCF1sTEsJcyE5cW6pQhrTEGua/YsQZ98EtgFtDQyXz0P7G79fV9Y
voOdYLjMnD3j+q73yr9JRIs9AQNfmOn8/U+xQlleDl6AjhniPJHqY3Tv8nih2LhE
yi06yuoVCqginjt4DUhIh1eTgYpcG7pLoz2tvdeKXzZg2d/jp2A84HDFKA+vdO8l
L0h56COIQsN31H729ZWpcfHe48reABwY7YAaOCDnIN321+UpAWRRN2uuUrInJ+/8
0YoRvc3cmrQLM3i7ydRhfp3LLs0ha3TlNc/LLPXrH0t6HZUs8wUzbU0ABBv1ghk7
bxjtiWHUQEaqhQ8WmfMmxGbwWYiFLAPolW6RthocuzOUemim42ehiWbvEvC2MuVI
u58c3WWApLlGF+sb7KcHfB851dFJWlcgjRN8W0RuK7N09OKH+Z6cfaO4GAak6Cog
ErwHWSG2gT9yaHhyby42JQ5IB4W3UAthJ1HwsUEICE2IntK0UrB3hZLLJSMy2ZOO
tOl2AVZuF5jx6YgYmahoXEnCsYjgzcSM3S+h4uxvMs0bDE7OGBjrD7OEwRCYxN3J
6F4RtRMmJqD2ABpnc+dM74r/trF0g2eOEay4FIJeWNsezbJin2e18OeukzBot+IF
Z9eSh53xZibTujT2qUmmu0Avuy4ta68awKQKjzlc/dpZX2hSGjN1iVhSL+3JSdbj
TADTXstMEjkJV4/XKLLtFb9D1qCYZRcTn7cimP6MS6lIR1DPlVXePEIQrb+02jW+
UgVOAlZsCDwTpRb7lkex7JuOyd7fjVtkrkzKFS4TJsVhxmZtMjE3t4xXrN5KA6oB
82yzliz/psRWNiSWOdhi6TIqAHBXO8VYNEfw2lkgrHCUaOUf4QRbD72MAnXhVdae
Ovhz31YFjSDjdfHyrhyyTUjugdkR9WJwldcr5gkKmr/8MAnBYoKcANCu2YEDZq5a
TS0s4kfNa2qfGCPQa81k5xdwjl27qa6dmOJJ23e045sSn2gklMqKx7BtStMckGK6
W3n+HvqGitek5iuaSc81C8VM9SodRLjTLC1EG6fIcaLxeJSi+2FtyPL5nZAsMRto
p7O8vIXbTBZ9Z4Y16tGVEdoDdQjTBb5gHS2H2dZLgRZTSgacJo5rq42TPjPQp2pK
iLLxckNcv81g2MsU/WzDXg/Q82HsaGb96ZQtu+9pb4FjUltU8UKQK/5Pfuqq9D9w
SAktitCu7nfFXz1Ty1347y9MtsDrROmQ11gBUiAO/dBmWxO8dgJzIVCPY3rRewEc
qtlOgIqUmjkx+z7NxYTyQH/Hu/XgCT0mXYYsWZjEYBAaJ7K7Pq7W+JlD2dTv5GqN
VQ9a4MXP6XIb8O/wWHZQxvq0yxY36vc3VTgMZdl8aPCa1e7VCK3NC+w0H4Wn8ERe
UJZZ1t81Cww5Vw8KHsP98JfZvTukzDeDm8wfErHG60kcBb44ZWJXtLy1B30WgMDS
MkSDuv60iApTV3SlwF1vQmR9C7OvhP63qDU/9FLTs7k8yV8bQDwoE3uDDOVP7d+Z
3irsJ9WyA66/JND73LLSjUncrVslmbpj6GbN9rtQmzjyAXauEYS6mpjj5mf+ihW6
v38CaCdwuXbYaXozq4B57YN6r4r0qmUG8ks3DKIWrctSa1nB33tcfTMylvuBWoIW
N8e3NOR+4Gi93P1L/EY7A7MeWIxpJVr2lRd8+M3G7EBNdbUNdeeZNWYJ/Q5hZ4V9
BwgF/8m8Y+ZDw7pRkV9B4EvZzgqid8Te9MpVry3R6fDFxG8yZBDkyi5duUwSjPXZ
bJk6SZbcja2NVHRXzZvNltHh5NJp/3Q/h8HJ7/3ExEseSIvz0lqwTZxhIIPcX1d9
v+HWKeyQZwSYMq4svPO4IPMeB95AuB1eHx3Y2vFwNZ8oMp42BPL5xLxUlw1ZWyKc
Lh9qIf/UEHffeNPQruRUlSM4b27Gor9wSu/srvJb+8l6INSKF1hI6ULQxFUybT+p
PCkdIeiDgQ/633XokWhFom82KcbAROPSZhD7sM1iz6TG9Bc2FFHA/BnGA93WJ68z
lzsXcD7zzUtc0uOo52PVOyqW7kUogIsVNt9x8S8yTJEtqSppNGQgPl7HJhd1q0AP
k3I8LWdDz3TVscHmsXS259p/mktLVVcfhK5VoiQcx4rBzQIbvaAHe7yCuzvxhd8W
/40IK0IcYKhM+WpKG8UpCKeQHjZE4gyMwJ3TvKiDSkm/YI3NaRwQT7ioWNghE3Hl
cRj9EFhVoBgibzezVrA3gVzL0HM/TTaQiNnO7NPhUsJKwC8T0p5I+Gt6c33Op1+a
GXHFI4ebdRn++H2zgPUbVOhwucT2U4v5zEt8mEGVj7fvRar78bJmomR1bKcynVpS
kVIj+dBAunaWGFf+NrNgvxHdJhH88gM/eQGNzVC0WgiHdlrIDg/JmQipxwQDNc7C
2FiJA63PwPWQKHquf/RpYjQYPUJHUCprNbyDGcxFJavTaR8zPiuQ5aDXfh0PNRvi
wxs8TQIN9IAOtKy6PI/Q5p1KrkSVGSIpY7irWrvLnXLEBgCSmXysLwbF7piESAdd
bAodMM8qBXxe4QoSun/gFRp4f818jb9G9dN4kbcGghcL0hxX6K3HwRTsqJxOE0Dp
yI2WIjPSlTx5uQwxMBhowWYymqdaAUAc5zh1fGwUY147smuiv/DcEYR01lXTMSky
DRqWHrHt2mmiZRZVnmaKePb5zmnmJzKzVrjml1hsOacWRSEO8BbWeE7mCnGfkAQI
lo+atYcZ8U476TfJkD8RqL+KxJR5wb/sFG2EITo6KF0Fw1SSyIvEnRG2hZgfPiiF
ZRnt0JDdUaUsKdKNdTU5lLXW7nWBOYT0weQu5hSmPU27wekL/yr4pmpiTK2gWnvX
PAS7Z3rfL11xlv3AiWOx9RcyydaLnLfTBys4mW4infgFoKazHUz7707DrIcYm2dQ
y3tHBvJ8Qbg3xYgEYQyd8sIBuhlioTqc11jFfLBPiO37rMfxaOYKqsufGS755hYG
5N2eXt7IqwDoYh1x9D7cPSlP6voGzzCSeZiZDiJXMH9r76Sk1uzut7ulnjVHjLfr
/zQd2RJr+p4/TkYXQBmkcFRYxF9NQEQhhswqo7VJ9KON/UATp8j8Wpk6DQBInu2c
+dggxgVDPyXFSYTxpvK9bVfCG7i5IH9AHSVKHewcDfqfm8Uz4R8SEamU6bkWe1hq
OYi2Qj4MyehItm3/EHzgIYSpiXLGu0Wj6oVOeOHSgs3z8cQDFkj/LMGopWzcKK6Z
iHasvzb1uxHOKHznzgjaz44L+chqfuFfpQyk3bQkQP1UcmYjnaCcJlZafh9yPqhS
scYcUmzZrjcNun7KfizpJ2sGDDzQBGCHNgHYraS2G+zSQaJ26x+Ar+Vql3OYsfQd
ixzbt3mF3yjZq2/GzefeC+qHsBP+rYskn+KocSh3Dp9650KLh7IB0rHhYcko1Sxb
SemN6y4KYNFXRS1wcGBWW7CNndNyf3shLtpS5jV86ZFUolNQ3xdIEYWUlroxndn9
D7Ps27CuI/1/5byLQBkEnzTDoYgyimoXviH3pw1eigV3R21NC2ZcjqG9X9it/4dq
yeXAaknPIjuUwOaodi7OvLP82PV8hY4VlfHXOaYS4fOKnuJv7mua0tmhm3mN0sZV
wzQqPJZC72ycljxv60YhAR370bKr+vmKw6g7m9Vzdu7VjnexWSu888cZOBvn3f6o
dZq/3SR8dkprwXrxdTlaAiF6ufiiJhIBBZ2PSBfrAlCFkQVrFpQOJKUXUppOb94V
g9ina2E+pcuXOOrDpZKalD/4CkN4lVThqQHy/DNsCqAVa7jLajADMiuoqvZuIMa2
nmtKlkXaAT9I8eqGxK2gZf+cAOnfXJIVzSSTzQSlpNSfd2T2X7mG9SQRg8CUQF3U
zTMZWVjKzhOhKQWcu3WBLFFuOd9C4SPfkR8hQyPRMsSsfKhn0pcsVhOv/jBgEJbT
Ud21O5d6lYSSYc+AogAoyners5+qoHmEEJaEhNXUxvZcSHYxQF9Q67EfY2GlLr2/
bYulJgx7VQxNJHEjO9yA42WMLQfvT3O1mjOBzj2ieH7QMeKZ2X44ZN0s6/Cwr1nQ
kLjFN0WUZNB1wXl2cqTwaMyVxz7+VAsU9w1izr9O4Fv8LsboC9SlqVIXvgSZLOiI
H356b+MpbN0L4BbDQ2xzQ3G3YnxDIJSisrRjBkNzHwlrBRlOG140zvSGtfczZecV
RTCkET9qa28DTs4fqz53hPEXZ8iz0OLHXvzIqqL3ajaEQG18uFCNSEueKp24GVbp
g8TE+XBsDt09XUezOcJn+SulwLwa/GD9YFIIz3hkvMaGc9c7FIxWCZZpVTv0R+gc
V8adz4cIHYfOlNYdotN0TwMS2YPrnLyaON314ZFTo62FviChjZPROhVUUZPwBAUD
jdA0x42rLAnJuqS9rVHASC5vkJZximRc3iaS87Ob43beL4tMdhCkK0u9mOdLf61Z
k5Oaq8gFy6RK3xi2QhF10SQKMkVg14p24YRGAd4QQ6nQlXu5ZhJL3wI2Ht0Ct98i
iH0+KgDZcl5TDOdiS4JrBgky8FBqexV0iohXtQjQUlReM6wtS0a16etgERBM1UD2
I6k7MjSnzJ5gKtAQc6XmIF+72ftKQ/S+D4VI4KGzKSFoazxlQzd9TniH5625HQFc
aOgSDj/cw3eeXQ6q40J45oZsJk7Eb93KIqHsCGdcmYQmXOoj+k2Pat49pgdeBfKP
2c3o2h3oxRnFqJBsNxdcggtmI7XYNjj/QgN8WdiY29zPo7cEbgQXq9U6tqWaZ7wE
5pv5gL6S9jGqPaTO3ZRQ1wJXomeZJvzce64y0KIKlPcCIYvCLAJ8DEvsSABNt2O3
fYzeo1zY4f7h+YFAnLGjMuLjZOWX/fgGUbLWuprI/6bAUueKesXoRALAs6PCAcs3
vF8KtKJMjU6Z8FZ/ThLrEhlvZpM58ebOmVX4W/7flAmSwqaHsk4gvEaykFz9sQlg
y4Jh9OW9rKRHwcGK77qQuKPMSVrQBtnKXP27z3K3CvXTE/TCfma5FTHbV7OWbloh
qyBS2J8xbH3n+ssBSyT/Q+t1ALETtjEY6m+e1B9BE4DMRfGFDWuQYOD98AhHk/Wc
bpX45oWDPvp0By7vOLtU4yCxZ9lFu36P4NGvEjI4+D1zE4OSjeYWX6MefC+bTFge
i34/veL7y+C+eujSH44iyenFg+rwEHLYaqKglVnTOyDkEyDMdO0pJE4xwGRLKtav
VvrUG7ceHeNR0bLyTGeTlYtUEcj82LNY7q2s3Y1W9tQqcICeKxYVkA/WrcpYevSi
gWEXLih8rG0Fn80OKxCZMGYs+T3HE+WHQGLRx/KnF6sho73g8qaFGbPbUNE+MX83
Q7BlAE7GJ1iVEwfEilIvJ5Ogh0wxIXWfamDTGtbynlpCg4V4lo5dR2C1NOVyzphG
k9wT92aAWlc5AVkYCzT8iyp9BLdWAC+F0RujJo+VizAlxlBeyXjpHlftzpIKRR2Y
cXeNdNBC8b7yisl6xuplON6UZokygp7PCsTSOcQ8G0VX1pjLq7MyllJHJTbbIwcT
QkkSDVvui/swlOEesQVPrrzED6XcFh81K0mhK+26h3gDWgUoI/NSz8AiDgmdRW6T
VIPyDtCmjshFRjav5FihpAm302GdLUBBlWp591lX0XXiL9wjuPg1gc8cyPc9TcNb
CMHa1CCqiNKgC8Y0Inagutn6Nr7fkva1UjmnCLFE6K0bJZeZmJur9GxwcjWWyC1p
UZ7X6WKmya44XPZ3biXLqUU1a+pvhhGiQIK3UmYuRyv+ez0JEozp/3sqM3+ee5F+
UPR1M8/cHAELKOWhJzq7NVGnK7DIT6DGRfhlfkULFFzeowSLiQ7uKJeS2kmD+8Dn
jJ8du9dSaPjdObqQDp769dkSc1abyXcz/RlwQA6twLOtTUJAEyv/zmpO+UUy6FbY
Gl1H/AyyNhMvEv9w9hdu/JAiFLbIPbcABCXcmcmCNiS4Yy7ZSkyUR2vjUjybFjxM
VZ/rgiFXMOppQAGNRTx2hdipbyrSRPfUYL1x4AUq8+5DpE8tR+45jwS0u7n8gXN2
FURLVGCCeMYqNtKAM+pkfpvR4eniv9qzzzFt/fyUQ3haTMgHiBzz5AkLU3da8X0J
2gNrmnwo9QtQjXE1ZYHmIXYyW4oCso6XlyK6RBJSCm+whF/9WR4cS5m89e561S5Q
4irUp6jEEDNdBwNAgxsI/ZTfdFWzQ/HlUFxtvGKf4GYG9rvaibBbwvKusyS0LbtD
LmEEGjL67JMUvuN8JpEM/QxhM8XmQD6uMLnz9JjzubXg/yMIaDmBhSGcYYAfVkdD
xTZnexkaKqdbRMs3ZWXbN796eEM/1Hr/+TefhDnFRRiMVzd+/QtIK6oExYKJCV/w
W/+HxBhMbBAb9+kFxJLoFEFnMhsLtkjc3oOxm13swEeY56J7C7t5oNeMIhS+oSDP
tQyGhj+2PrH3r7oCC25FtxFd6VYtHRHoM05kM+uN0fO6b722vVLwGDMp0ARwbPE+
naVX+8GaoHYNPtkea7BG9DBAzujQwISRK0SATV0BBW0BYGfWA4waz5K1+OCLREul
1pNsXIS0DMRohORny33rFYLzUMYt0Q+mdQ8+zDt+AYRaPuHlFnRCDbzC5IVoO5Kw
0yXwRXndx93l8piGuAsWpbrtdgEISubJHp7mxuPQwrc20froXvt9nzziORJsUCfX
pnTdVNdKVhb9tTPUkospPTlQbCMY1JtWjxew2ulxGKsbVZ8yI9MddpoKQ8wFTjdP
xpCsZs+DfW2Uvxn+v/q6I7YIXU3lUX0gcinHyi1u2dXVan49Y330cSa60YYGQmqS
CZkQkjX4bOKPQDspCgwj3l8ZNCExusUZEorsk7OT6b0lqg7iXyNtWyZoWweA22av
D3O/pKPtUfxsJUHxKVlKOCApTwOs9dDrqm9C8/2aQs7l82ht8ParqLtFbjnXpzIN
J/szfJ9y9P8XqI5mx6OE2RO23X3pWi+GdMfmMp0XCv+k9NQLVMfooW5DW6lBx5Zq
6/pymC6mGvdcTuymeDyA6qBR5VarwWRap9UnDDoY5kG61ae5CERuYVvYUAwDP7qM
yciJDYrw/AmuOIdqAK9cHRqy9TyOaztaPZqgZX3/1VktOZ6Mnhx2xI1UeyRA8TtT
K0vOgpw9zJTItWA5IU63VqCQazvaCN1I716LkmwV17kml9gWHJhQoMCVAkUJWRo/
A+VcmNdK07hTt+aoJrN+oITa3vLDVqa8jcGTqc/NcDmMPMU61FFuwoi31O/PUd2V
wiGBDXq+CmbEhRf/Pu/XNAB11HO/sCEhKoPXBCx//1HJDpEha5eGGUAUmEDgKZFd
j4HdR0Dug/rDeH4IpBaECsspOjyLMFdCvgEQP5N4N1bso5A+XbNhLhmlKmMvj4he
mUIxYVW3IuNRVH4HZgJPBMh4v0N3y8jsfelO0xvSwLDTq6o/rnnF33tTQnORE9tN
TnA5rMhJ2N8NXPK/upU9JQg9kzjfbFgbJzhtRukf6ZEWnxAgkNxDHV+U2NlitguQ
FW8tlF9fSOElizmjBceCfdKznGlxX6yuffNI9c+EJEfXn+bnDspISiuBk4ZxVxHn
AYdATO6qSepDWY5quP1rJ1IzkocHLJy346TPBzkJIdxzQNi5Lr2azIpsbrfkK3Gr
BVOyLBLGRvL3/kI1zZeXCy7E8SBBkhP66EHHy07YXGh1JeXK8AKJGJyNCx0fmBWT
+LyeRMmqFVvVLdZevaTVCNRyp4+1VEl9rvN3aEn88gzObYeMD0xpJf1Ecvcq2HV5
2et8ZnDI3G5U3Mbk4Lw1UIBe8ouDj92XgV6u0QF/KKl+xthgAUDnoGsEaEkjijYt
Iy6V/uoy/LKizXc3xqKgtF6oK/1q9KVwX4DOI+lrDXzC7dBVipq0mRfdJSlBDvmc
8qe356Tz+Mx8+1eiIKvIvEM0upSEBAG4f8YamJmXInua8f4FtXDSfvh9yzQ8U8A/
kUKUkeyE47dtzFK0D+eogBByvD/MBS9TrkJQWDuqxnD4+TNo750QhxCaxD3jN7vP
ydWrk9mRezo1kZ+lcePn0E8VfHYn1kCdfReJomsFDsB+yp18H0WlBp/AAONUOq13
NlYUJUv9u3wWyP/dv3BhT38urqx6B8tlkUZyvMzo1U+Z/znZM8uKjMqRQoL+JBvQ
ufJcEOcGf9dRTCtYB3B0osIEUCpTyQOljyIsYxlOMjCBpTwbxODM/uAvO22Yy5jU
MTElpcmy1xbYOUHG/a4Zi8Yi3Xjb9wxa3VoyjmFk0lMyFRK9kFzLIsdTWH0IC1dS
g3G4yJrIa8nKV/AzX0XacQQrxRTH+Yg82KiVwuYc9q+TBoGp+M9Yqnd1R+nSs/uh
7nOhRfVFE/pXi/YB2KolNU1rUgA+9pd01BJg+VrQ362ILj6EPvXGQhK0VfV6mvIY
APxLQbAircZl5Ej8KUMP6q9hWszAyiP3Fb3ZmlHvZkwJmwurBenkbHqghaAKXpmE
zZ9g29RqjmC4PGFbg5KmQqMZjEreNPr9BIfa8nx1EzgeHECr3Q+o0sdJl0VIBSXb
u505S17iFNL3Fhfzo4LAqBN6AoIXGp2eg+s0jLkf2W+MvZMCeFF7TK5+HYCgP30q
53y2djXvxbx0Fl6W2/CljSin8gvjC+yxm+zbN5G2uSBOlsslCO9/caYJchj3AelE
0HabpKuN40kXCRXS9QEXi7BnnURYHonNZxLBFqgMoBxfqmyV60YWBrCkeA3F/9JV
ktBQG0fk+cUQWy419k1KtdCnwwGLjbjvnlLjCVQjRUFeijQESdoor8qKVxteokxR
A005jZJIw+HlQIiHEp9GGWyvX86ACyyiQeOyFY3W/4FiqFswYf+xzOOHb3ADNduY
iLtlVJV+Bn4Fp1oStFHC2l1cBOlJDlZphggKffvGn3xpvsx7MUxbSVM2J5CM2Mak
sbApPMeQB8Jw9GNCvOc+NHM0q3gcsvf8lH8lRK+j6WSN0px+GqhPP6tZnIWM8/Bp
CbWMaIJZKRWWj2AjT+z2XgmqOYLAF59njOBJZ0ETPrCTMZXKArn+boQSCW4jUjEV
AyeG/PHVjv4VEYgx/0zA4qcZJntY/fmX8w9NSfC/m/9hT0jz0OpjNbcKcQhW6yN1
C3Mb77Q/ljGUxK+QbWAaTBbElCFMvouVSokGsYpZ2zDHcDA61oQaGwOIo9OCq6s3
zDwYoIff2qyuu9oKOuSsy73Q7ehzLk7i4kR1C5LAR1QNnzspkrR0fuPGsZfV75/2
T3OKVp+DvxGgPFHPZrZUHzeuXfVSrppMuQYRlTFHlyGbAPDLRAL4ZQJWHyDp93mB
pIFbznKYO6hEhX4XBoKLSvxOtC+lwMLtoxa3g5LKzOOekoraMYaClvzxdpL+6Orf
qHk6P3WR/9Q/OKiYOL01Qi/vl1g7hgjXCCiL6EPTrnxMGTCD0BLAE/byiqc+e4Az
MOZVtaXIlWeS5Ee2PuPsx8BQDAj+9+POmkOwdwDivj2Q9r0BxP9L3nzVfR4C3Omt
SydymtPKED/eiBMIJq2OJjXN3FRUyADLXCelXVg9es4tZ8hSaVKcKJZfxydS/mnV
VX/qCync1E7TQy6k1NRgiJteC39Sn/Jzfyuh7OjKkC7WtjdAlbijgoVb3EpbnkKU
5nvIDgA6O+003CYoqOUHsoeoGEwPMxOohtm5vtT+lGebwAsDZcIQ8nB7gqbtfnXY
kHCDU5m+nFIGTqnRCJdhUttz/Tp0aZEabz0frODlQ5p/xWfI7u26Z4hc7LPKA9Zi
njoNJLsmnPT2jXpkK7Dkihb1wD2krDfsaCr2H7MhQx4puBhe67i87l/TtT08t/5k
d6+AHe4Dd+wcnKNBnLWUt1Lbbx0Pe5sI0SLf5F26fTja/tj2a/pJ8bdcQwKZODQn
3zUUYQChvwZBb6v9LZ1iSXnDpZAzu70J7B2qsGXoaMxTkiw7mpFXkNq4mQDGQSw2
WLZsiOSE6Lv4LyT9Su0A++40UCt3btXqGKOWCvf+x2FqKB7veTIw+NS0izXBWzLv
d+A9vIJ1dqU2iFV0t0HZuagvdwqZgT5jTaQrLdygjyIJdtEo3NdPXaf0evfH4yRJ
wnyo3C4BzCfM2oQmuPYkFT6FJ/wHKODnAw7OqUNz6Z4u9biN7HloILttk0RGfFwt
Ru+IHjdrPGPFkuzmSwFp833WSwaHs6pDtG7/mF86wmNmPPDVivKwsnkCEB9g+6R+
7x+6XRUQpTGv+grbs9HIMSwhAtYhsuRrD5J1MoBjtzprQBXAP+WAFpfxoQotW/j+
c7NWYdVLaEYuPWk7sQSaT+vd291+g4QnwbL1OkQtvLHI9WezzsDBh00zRGpPDe65
St8S4xPyBkD7Ll6zNxbrvsOGQWmqWKl4oHrYUJJdb+pEeO/Yq2Dp0QW5/Bkf+6/A
rqaSHWcy6mLKr2oByuSLpomA0y/Bg7VgGmMh7Xkz+IkKI7n3b/5uF8k9T7gDS+29
rrhWVTAp3QdKrRFwBBxWpBvSlkc50gxbG9IJVRi3tucabVi9uJPW2uCBLefu6/s9
c4fuzmpUuLKua6lvMiHTC4VABC/sFTb7dJXRhwEl68YwplPJyf/iyqK3/ZWHlZVf
NpB0mWM6tLwblD2m0EE8HMqVVjaZEyER7WoSm8BIz6CZAUYdZWhCa0IIXYFdH/C6
P5konY+OjnZZSp0pi9vApyoLG/KIhqtkXp6YhupahCSj6LUT6AVofNdX1tKBp/8p
qZSJZO0XLptfxcNYdEmxPGgBrmIJx8hE1+DNv3vlBMSHb0dp+w6paKv2L+ilwxjq
k3cF08cqfcOto7gZkETyQB/5rPRuRiRMJBoZl2IDcLVVIYOCUDacjXeEZLPOgHKT
iaclFT3Lp1ET1Sslk7pctBOARoawy+nNdD9uwR5OXgrgKuifPVk1Xnsx2cQPwl7i
bIfa9LewwI2VQTyuFqO/icY3XMviwVM9QOBCgrRHZ/87fW++vxLVLntam2/W6xmV
w3VJoW0Ie6RTrE3yaXbPBuRJ9MLqAky44SyQ0f7Wb9z0eMm69nzTQ9shotEnXYDZ
lgoocIdv7hH4qfGv/8cg9HRUTymU3ILfYUFX1GaZOKJErPAhvQy6zdGkYzCCZX/L
7GFgPIcVcJWRhpw9ouWUQqeKIgypZNKc5Y+lpO2smXaGsvN4Z7qlSXCIBh9TD6Sq
f63eyDa58c/riPKLILOtpHXGWF338g2O8T+M7YRVkk5J68s3JEIaFHq0oS7EDqK8
MqnfKdBfTlLUkymZ7s/yMfS/yDZ1RksCf43PqDzijS22y2G/z7I89ddrh+9b2wHD
7trwYI5GTha1qq4+tOFoumLeB52UzmnU5ib9PgCi9hAPY07pCQMwEYHQ3T+3931z
KMO2MsrnDKpBg9ewFtuP9NCoI0wSJ6fH+WA/jb8a3Sjpu0UMmb8qApYq3RZaT+fZ
F7P0pexFgCiorOgZ7V8BWijOh7Nmlu1bkMd4t/j1n0cBg5lrcmTK2gq6QEt5kn6z
48LnOaYX6vHK6rI5T/UDrDYpEyGgvgfk65q++W5jwUquWjFwLJ0zAiQCYZZOUOVU
7EZVqwzWVxQJ17li8TneWby8sbvvy0gMOCSy79Tt9fpzOm/sTT8rR3XPlvU3EGok
0rw1BTYCb3K2bnjg0ZKKlc6il9jkZZJmnpwqA8W1EA8jtd+bgT2UTU/gofVJy38x
U0mTOLx8OMM4sxmX3UVNStmHoaUQt/NPPvr5Y8YxccaHab+IiNhWHD6KbW0FvK4J
BYmmIenXN/kjQXAobBTZmonZsP5sdGPRK/sNj3vUrnS0J5cJhTCx7Ru3RtQyXH+s
V7Eg8ZBZjJgm2tLlB9LghhEODOjTUztMtTP6L+23nJQCa4n28jegqFRSpRo4ZKrq
3SnhnUi24xyrlwLUocCiMCrWkJmOVXge03JTGmq2P9bqDz0wT0GOJKwS3dd8JZuB
SaB2/DQOAkJ5p+0ZPWpnFJjaOvcPQCU//6AObNzUyMUFwzmxuGe3lNxN7/dGBggD
AYVw3xmEk5LLO8xex+mSIo6gejzv/GhdbOyNt3srtLD8BI1OPy+raRF0vXsnssuw
SXpOSECK1oc+mDJw5hDRdMdNYGwofY6Aad+YnKCEJKP10cYSaCVzbvwJ8vXAwLsQ
04aye8r4sGxLHDy5dBN+RwPbcvSR2syMCpPcc5Ob7kfZWmBAANql7GJxJNURCFzJ
OTMKAmElvUEt0k1vTRiLQ7dFDY+3v0uJGyf3YydbQFAkpF6P386MFrKurgIYdoN3
JwZtZeJoYLHSyJV4I8YJ4LQF6DbPkh2tW9mXZmPQQZqanMX9iVhSZqNCcRZjZ2RC
zQpG+1teEE7IFtXNmktyXi7i3zfCxz8UmInDUbeZ302i9av7COWMkgZILAf/f4mS
SJLMQJIiO0uDo5VSbt6MApEK9f32eovqXZGp/a31mdU0bI9yNXZEm99KksXyxDGE
FkqDfD0wbv7WxfVk+9bRTqXyQY2kBzEkeREsE1FszVn3zxTt1EpcBmjC0T86Ax0i
yBGplByzTs0pqpX1ZPsh5TEk9knNEUevk4vMPwCMG46qK+FnICXI/KmkZqRvCa89
kfs53w7JjSBtBJG3eKrqaoYRpQXCn0qPXPDquwSDb7PWeddajuoOV7lWM+Cxz7d3
hROU01h1pvvXO3t2op5Xi8070PUQRWk0lDxctqNVWidtM6Brj65RtEDd25+Qqqw7
1HGamDbK2piH9PjK4q3/1fXbXj0azTsVLirwP40nyhRZJJj7Afa7B8cjWMLMC66/
tpaAeBt+du9LRp/NWzyfYKAgY+FzpVIAh6tJICjSwDQQol51nhJPCg5pEwtSxhqp
R0fYscw+WzuU2xHA/5Kk8W7ZZIHNCk5qRrpc7d2bUq2w+OiUMCOpTOCH5MjUJqm/
1r/M15PD/Xs5RnOWMcN6xDBsfRwcPlgxo+vdWrGJA9uSCmI8IHtChwqJwQF8wTiV
o5v0saYPOuLkdh+/KsLDJ7gRqlrBRwE7Nt9UqWVB+Yo8fFosBm/Vf5ocoiMTN/tE
liMRXFzibIP4iPimk2Clj4vWHIWetP5iysfaTM0fl2DH1Dhk3eF3aiTRetLUcdTu
ev3+/LFz6d26VmJDWnxP6XZnJ0UaFeyZq45qPbix9/dTDdvH5VA0wkUYi/zPVuL7
EdMWDYeJ12rKlzQvLBJNLB1q6/TW0Qt0ieID3Ev9+ZBvcrGPmABwaFBE+hf8sFYp
wNikUEes4Vo6gr1OJodWSYLIZJfOCUVWDJmDPeSpg46KsHd2inrJTDoao38NChoH
1QgtxBfnY7P3pKlsPq5v7TwMq34d+hidMdV6g+C2vxyRkP2bv7v5QJI16VimIQiP
VqS4vn+O1wc9+GdqH5EOgU+dhLUMIqKufBuKRk59ON9G+Wy2VRmR4qzSwYvjhujt
76pB5EnSGM/tx/Qq9QPuwfHYA9Az+ewDl0E7IQ30ol18hM++8iI21FK0vZ4ZbDia
JIGaiaLALkQGw55/OgN1Q1J+m8z5rgthbTbZbPLOzMJh45lHaxtcu3u6+fsPTYKD
J5wNnt0jIhqqKWNrLEebY91ugfbfNfF60BfU9BcL16qNwBrLXek/wrzl4hk5Aev/
Fnyv5cNSi/owRlVRqsevINBSjM2FLZpcQaFC6Yed5zCt6GfbE2tPoH2SaMznk0DU
2lwgskECYRE0gb8MtGhTl0oSW0pEQXvCVof6RmVEFPmGJ3Z7h1L+71QX5FAqhCp6
YLhebEsRkBm0c3k0yGCXBGwsOg/Oa46c8mrKsCZ0Fra9OEWPHZQQ/KjmXUHjDD55
f655n/SxHyvZbk9kwVovgjjguqHJuAsJYUrQZ72wOHh3qq/YJ1PpDbgd4r8vNTxP
mzPnd7sHhA/jJZAtmUfQKYfDc7RrNoGdJ0Yv9IStuhbKuOVe6IjWcm/fXB5TYniN
WgOGlLko7mlKIZSlozJIPFMpcNp3NfFzRfMnGlJrlH/eIouA4P0y8ie39RpDc0aK
d1WeWDWEBb6HpCKVEb1jXS3JCpAjcI3iKriSXYyKvukc9aM0nSfZhDUaYxL/l9wK
BroLAGqqtGZwoqP+19uCIiEQbhnypUytUnkzN+VLek8uqE1T4qyen9bMfayesZ9N
VPWzqRKMu17Ont28UTYJpkXCrmatVEJEcaY6xo3Jmqiv4Xazjt5+kG9K2ZMMfEzh
JVnOqJWZf5XtjctG3o0S5tg84xD9FTmhBMYkW0y62IZKoHnXQIAC179dxeDzNXgB
ZNKqN28/KMCveixNs+bhsZyPqksFqQu6X0EMxodmj3hhqK/8NV3jDFSwNc2ONJXd
ZTKIPOdnwcI9psMy2aKR4Ndyp8eXhT+I/v+jvAwrttx04UyCqc5D5UJ9bwao/G+6
11xT5FGDvjv6k7+Ov03IGatZjJXFq90Z0VM4S1UmeIdq2bI6LDaVATh8g7gNqVC6
c4mRUqAUt0MEtfNNyGTeP+RaSmo5SqbZiltl+WWT72PUH4xFFv6rf1ZPUK6OcYES
1GJv8FQnAS128+FWNl9UuUs+s2V14Zi3kB6xpathIgLFoBYEe9OMoFTvHYheiaTG
4PTfFtX1c5tjTMB2H/4Phfg9Al1iOuI1s2hNEpM0U9iPsbrLUCQC7Iiu2ywv++5e
6nZkNt52mXXgXnxvl0TqozT37QSjY+oaZ4NzHkz06H8YDJJb4DbIi3L7RMZHsKQ/
ByKsSngO6kQh45IRHBne+AXr2xEejnyeuTf6D6NYUYg+llJAzEsVO1LtkWozcUeS
yoPRNBzX7wAxAy5KZXhP0Q/wN96ehnMzH5scC3G0r54C3Ivgfglu9cUrXEacy1vP
Rckix7sb5+EQmkFENiiumZe3CvdYuDrejivHxrELlkPAHqrITuERK5ELD5P1aUwL
675ZFjnK6rtd+DVrU9SBhlerng3MnjxTn4bq1M4liEgiGM8a/xTTu0Y2Z69cMEe5
++to46yeGztm+lRYq18kcLTGHHLn+AP7evC6C8QLJsNTQugUQUqns2c6Q8rYxis7
TWKyMil2LuNxNFKBqVjq3sPYOBt+3LC+FzFhN5/gqEBTcOF8VVgECSoACSOisvXl
4ukJVmjmbJYyZgtR+ZhD2VOuNMz/9mYxoLstSUEWWU+Co9Zx2KHt3rSiHi+d/jSb
oVARpF4DiqiX6mdRYl03fOPIWwEVhiVYVV0DRineMfM0yiLohLiWKQsmQcQjf4ag
xyHVXa6XnY5146Qw1JaBcHUcVwBGwlp634V/kr3FkIE9ZkTDvQh6Rx+skS3VbRmq
dIyhZhEZ8Vdm3IPPbbcx/0EM+M9lB61MsHnp4NgstRMpBsHCdhPjwrB50lnNbuaG
rRjyO+15nMLyvaD5dnjP6MYiy6rnT2xnjGPQJTXQRYTD1bQ3OYCyAJc0q7Wg26oP
foHOSoR8DDnj+ypFCsyPgRe9IdBNt6BNZS/Ltx0rEHuhK5E+ztoXXlnUPCmPHvij
I3pSfKEA1pmhKl5gF9mDfw5y5hKTeld9mWtX8Dx1TUxqDsmR4GvhJ2ay+qZj9fkx
zrRlS9a2E8JAgBrgRoec5lpFDYCLFKIAyn7kdcpdazRhiTiWuIdKiiIk5nXxaQck
nRy/4+wv6VvacJlbSaM9TKLO+gru+tHrYldhOen6rVuh90p2duaipvjtnsHPIDYI
vK8h+JUePb/UHIjt9OCysVcUliUwjfG8NmDgFkgypuxmka8YfNCJ07vnjgm0+/y2
GaB/h9czrqvkYmXMmv155ueCOCgtRJDCHwSANKX/kmMb4h4tpwwX1ZGdICh8ScLq
0c6buVkWnoS5CeR/bSu2qFnCWuAfYID5cHV+N1t2FcWzeaZdYlNQkvjzMRqqIsCn
smr4giPGX8TOSbZd0PGSWl+i+gkK4OUzgVqgNYyFDo/9Vlvl6ixz6yBgFftyCo3+
yH/ixRLdwlaQzyKwhTqdUhfo2sKD+Qr4CD/rqRKbdrFDOb9s3chV534Ev56iKU5p
Mcy4MT3zyNa+262rje2lLzQU03CEDoOUuEUT29weaFO2H0wjFiwOcBEca3lYxs2J
opgXpamVKt9VXU8cJyAo/fBZwAGSvCtPb8JDmzsGih0v+1AzPXc9qLazj4YAmGDy
jDyBP4IbYWpgzrgBbvsD8oH1PUrq2OTq6y3wshhfIM7KBCnTAy6HAMLFVxn6vt4j
LdjSnaNOTvA1lVjw/qiEHx1fD4oV/XR44C+8Sr7YeBhgaLLIUQEX22iCSOezc+yf
jXBX5WsjbRtV2miFS+CKSiC5EFLbKUN4BY41P5ZTroyUrFM1/0jOPq368gGjufYp
RVCSqw642h0OrP00KfGJ92s7NN6Qs+6tZYgZTFjdWzJOo9RS40gbXxj1qYOl36h5
P76HaUeZ51i/7Qiw2LEcMdGznWer72Dsqyf1ixe7NKg9soP93lRhH+seL0CfOR2u
aIdBr/j4n7JeHgSnqsZCQ5BRwa1XuwvE0d18euWtyfx73pxQ/hDKcNvNTMd7NyWs
N/nqWA8d9T1ZlJMgqPX3YEghdheLlXhqwuZo8uQt9qi06+JCv39OJWMqf2FNxvvE
UwPda7OCwwDYiosydND9b9fNrp7EwETdRpVrw5/xDFduc5QmDHcepDGWUEPxuRlr
fWnqRtVHAhAAoi0zaDkSB/UfGIp+DZaETM9sPTUUn+3aUH4Mnp/QDshXt/IrowT2
zYkSIU9PmPnQMaPdcCqzwfniBt4efbpkFmfW2uZ6wl2jYn+bmd9Sry5tlR4sXyqF
J82LjkgLpFgv9wjQrDlWok5FEhd0nqXFfsJ5ijJGCZXqP3cJjVNUD4l7vbpoCwX5
QKuJ/FQNEnL3/nYqDVpciBc49W4E47L5S1WU9sOGF4EIqYh8Aw/HU2urJUpc3pfv
jgsot//Fgr9D9qsjfEgeN2e1HBXsWiYmWT7r9ihuTBRpgilTlOMyluPZ4w68fItI
40rmWrx42ZFWTYHrn7J6Do5VklU0YlF/3e+TcHMyHcfssGUMpJHfJ9k30xcsS0nL
qcjGJgr5ifpe5FPKa8Tad7p3vOMX6/BGvm2soyiWOt4GmjItqCrSc2Ra0W1eudqL
wEEyhHvNw1/c+9JZEMB8BaeeVHV+zCnuLE6ya2fkknglQAIHkmKKwPK6X+ttbB64
/sKZS4SVEvgKBcPzkYQxQRPwMKyQy1xBlw/GhKVCIjgdBlhe8ItkEQnC1JcYvZhu
Ow9DboolL2tVEJZPtRLWHltlzTmpwIAZripY7ge4if3DK2I7bMhwVNrjxC0983mq
mPGlPorvgrCzqdauUMgLAlADBkJxvQLvdfbtym7d8hmZJ1127xCSwEler105YOaj
vWC1PVkNbvPWVOqXht+w7Cx+z9m6ZPv1VE0RUyBnaOHoK5hbP3xPRjJ663KXFrjz
st1P781nD9rGO9dZeaF5BTxbw+yEj5X5GgLQBPH7bVGkM3E8qF4tcSRGAlJ/BLm2
K+TEMU9cyN/VRS1rnCakq8HjZwTdV7OhqgOgo44phqs2prVNCkZWpeCJbBzNQFmC
W9jId384Ho8WSeUOEeMZyvDk6aujlY+JmV+7Gvlc4yorr47kqnqXo5jiLqBB6tjX
KjHZ/dPfCaWR7kxHl1W5AIu6yhyw7Bb8zDukPQe6GcOd/JUbPQSBAmjdIW9WJBo3
2kS442SMWIpFpJ1HApn6dqWU6GnqaSrPoXrQ660WCVJoYW6GkNaiIEAv/s6ZeKe9
rYSgAILoRfN9R6M4BBen3aQuXwsu5Le3cNotiOKpCYjd/LHhlCjw5sUTXzfksoI8
juOC1b7BRlZB6mYbBMdEVcL9Xc3oh1F7L8SOjq8HRkv/JRTPK504Taq92QQ42uKC
aYADEH9Y2VRjSiDb/f3CFEvOhi1mLeWZdNUCc7upH1f0Pb0naT8A6HVYjhQdYXYu
4rv9+CeAHtfpUX1vG/EnUYDmrPvaqUub1GTqZK7XAy8+gGtbwh4ZbffUpS6Arcas
UfApF+hoG//+3TC3NvtUQzehkFyDHSN4xtbqXY0s8UnXpUm18og+IuF/JI7C75L2
Vb6yxPHX9UzlUurUXpM98cLF0pt512SRzM5GrrbTWvbKQKHKi4ZOvIbro5UvQqGz
IadoW0uEH0Nd4rvAkeRJKtNh2OX8kl27DYVC9LPLAw+pCfotlD3moVgufQNuVZue
6y4UgnnV7IbGMfv8QwrnSWE0PnkY0E92jeLCmHsCuz2IZvC4V1kDTMZB/nfahvno
gkwn34nWJzel4JsEg8gNUCnyIQnLB1NEq+USpexlUFOH/ctObyUoio2si9A9TBx4
onJK+srhOA8RUMpQhxUVlIXY+SmU9kxmmBoYZArrAUB6KMsU2Ly1T2w1ki+BPyoo
hisxzTRd5DI7EN/cmkP7zuG7KyYm7sKEEYTYSVhrKb+2Murlm8EIg5fM1CdENWZ6
rqeMjFMKBZ50oh/mp12ecAY9UEElcukSWBUpCSqPBoJnZ3KcRRMZzGFjTBYWh3yR
8bkvBvfM3+h+QmRwZJaAhH0PTrfj19mrAObpgexBN/UOnkGYbU0INrASp2cWIO6x
UMQn5gucHzJOfOjWTJ1xQD0hhROEazzX4/aYverfAWD3XRfIDWeG6X87hEie2Ogq
vpc3Q0lzPzZifjHW3TbYuaInl+YChU2Dwh8dX4TUro2d1iBCC+FM4kAi0jsb+MMS
hea6WRGz5ps/gmZz7CqgxpmkCAUS7g4w/PLqBfGlK/fA190OOtAIwMwJiA2SKXiN
z0jYOsr8FQqIf4EXeopUn+G+PRjG9HOs7wy+esCrVcWMmbcVi2tGdrYlHzps7M2K
3k366wIdqmQBASL75QSSqByyUS2lc3xivt7oNDyILQyfoIO7Z2rELYiZWbmxM1p+
oBONjjpgq3wQTwE0Jp1DaEqjKvfm716ZZkaen26sNzKwrHdv5i8Jb8LOxg2HI3Ph
sRsLentm3e8k5FxaDXXSZxNLW/IEwc6XTUG7TWxf+OYkvKaDE2QsObjH9Gpbh1mY
NHgwKLyrSonultZxmcf+q4gNjm8hpQAQP5eqjN3NwegAUHwwJyQykNqcsrUez5Zf
3ne9kCD3sGhqEtzvifb70V9vxVsQifnD9H77o/EhhXIBDA/5OFqGvR723qPJJdxx
l8/318kzmVpENqFN0GyjB3A8T0AUSbSEynMO2HjnIeiOYfyjzgaGihky2QU3bwkI
TNwqZFKvPkjd+mNq+GDqfUu4H5kkCO1PTkMEh9f/Kl34BTMj6/uIeKgNchb2DEcp
h6heWudTpVenq0V8Al27Y4zIXjtgpbfWiiTPrIsMaRw/3wbWTdSjANb7XalTUJ8i
AztFwazFjqGyfxQSY0ETKPoabjod2tSJXfRdNoHHKonRLKrEEO+DjR/pDuOjdX0O
i+VbA8lcg1JBVum+CxCQyCyXwSX0ugYaRrJcqmSggL1YJ/gbwj10mPGqbR6mcMWe
Fj5yud6NSZFd3NyUsjs02Db3OyLq6tfrnX1j1Pa0wM4/jErNvyikYsIqN/Va/wVf
tccm4e+tfLj7JHz1+NrRxIFx+/Wufj8o7pNYQ0DDYueZURzPuL5/eeRykiX/lfAT
+jF0Wrs+CYaQA8sdLK17j7965RKUKI2aVwBLWfrX6ohHvLhV4pgKpgI+AkblU1Ip
HEto+f9ZYtPK1QFsQxzwrGipwKdvSYmqU2cSq3xalobeX+fk16X/RTFO2jSfYs9r
5gRITVFCrnankgTgbH3B6pUFjHZG8uo+JCUO3YVaEt7r/m5g6gB9tVsVgdN0qTDG
laHtIxfZr+vX3VqU6Kgf35QgdSKC64tkGfBQGNw7C1Co+GgNeiiyiI9+telK5qI/
UtOq6wy/u6PFIV7K+igjUaSJFq9QKVVoTUgIxVIUHkzDom3/XIVvNuMuIgwbOlqD
BRFEYp7hzpswD6XkfNHB90h0sj3zovX7/4kOQDuTFjPfud3L9iAP51OiFVer/4gW
TCHYJ44X2quREfs4rOHuK2Mmp09YL6yp9Rd8+Z+xSSXwyud/KA5FD8VqSnbExYHM
p+0BxOcKz+RqLEN+IJKDahUf6bNMSzPlRu4G68d52mNIAFz0bwhZsi3Eixe2eKXR
IxcR7om3v+Ai6r5qfLHg8ZMbuP2vP+XGOoaFWDj96Lf7GzNdDIMJkC+zUD8D8VYz
UEvAGMilT+XaB2Xc90+T6xzmDETd38xUIuWfZgPXr6jFuREMbu4dUI+p/B+nLUBl
gaFR3SekfuX9nYy2+/IirgXk5bgdbacojj7sEkabXB2ok9cdvp8qUT2VmbE8biTF
hRC4nD3zHPImerOL5HOOhSIaKGoN22PW7S0Y+IreC4lzmEzcHsb84W0ssUnSv4SY
8lhrC/WIHBCVmYc3fFmRexJ00uu13Ggp6JUd59C0fUJKatPG5CL+kvPA8LHDBrwt
fLpZdOA8kVUdJjN15Rx/KdxVVG6h3Cm4prr1OaEL1oiNRdj9huzJt5JCvBpm9Fb7
1cIrmf/cMBeJPfn4ugerlLwXLxJGC+lHTDXI4Cbroo7cfZ8CL/c/9oYErbha4xh6
OnWJRZgoY718sklnwe8hU8ciDnOGGajPpuTwJhcTt33fwFKblj85yCGJN/Prqc/9
u41EFzit9o1TWAJxo5NGU4qZVOyYJopo0QRc08BgOiyi+BFDE3xN4Ewio9xAkC7N
WGh7bVarWae3D+WQZwKxdTinM26bRZNOFmRRIuUYmmH2RvIB1Zs7zWuXUHztxM0C
lcJeDfgag1o7OT7zkFCwkfYxM2SkBUGpP/a/7WKbtNS5G/g5apCsDYCx1GB7LkZO
HrRboA+ZpooPRKSwduQOarbiyrkVEwlAZNb+9msCa0D3MpS9XMYXpuCNnDA9YGG/
MzMZsqWQ/LBX6eu5ESz9K/PC1NV8Cm/ZEXqnI4zIXLXb1lbbRxNgi1X/+e5FySzA
b7bDrJJchqjgE1Kz4gC9iVmjLxy0gJLtuDuO0jn19lazGny/4YADUwhfqPX4P5Cd
N2C6cH9yS1dySaePICVBiF+KLsoZZvDjijxSBifQFvzGS6vqE7Qn7oWeyv0rHr3v
QkGAtGGuillrDhz9nU39qHblzn7Ii1r2IdnV+1erWxhY6XLOtA0Hc4hIblZckGlb
ndDl1R4TbxPcGTsbt6AocxaE8+/iFk87vGvSXnvc6YbHMiE/q7ohVyxCw4QCigta
gmYmb5QYIwZGjKv96V/BG/KKDi5W7GmRcLaEWJ3QRuV1x44oKEDpIsU+qSrvy0kK
/8+2qOdKlSIXgC+1CTY3nC7Mwp9fm4pgDQTqxQX67BDdiH1YsuYvMa+XPuuyULim
dVgqrCnadvUBKVSyx7yWKiKhmgZeXCI3hX4m5aEmrJAQY+TqY/KxBa5X3qdaqgsm
JktmuQpj/OemnDlmsFYSGUDDzmoxCuKozujj0fzPMN+mrJlODauG9cDLSqxNTnMJ
nEerhZ3CRDgFD7sn7kfNYprg4cQj7SiksrBgkW3Zsj7Ebnn3lwOKR5TmC/eAa/Be
KRaaUyS0VVwtQmYteroC/UrnmXz9hG8oqO0bo+3Sj9kYsHYt1JCDEJrwcRe+hMNu
2GcaTpAn5xpzuYREr6UAgTMEd6c0ylOF13nZi2r+W0qlHZJIbfj5Fv9kOjJOXYFB
OGbCkAwwjpU2hUcnAlehki6Lg+K+kReH1OIVF/oPKzHPnbz8iUhsnVJTi/FTT9CH
Nnl0/tOx3joSqi9gs2KUneY0MqWbriXzFwBsDXydFoQQSdCaeYnsis6tU0Q9xQrS
cCqCdeykFkMut0Q543u5pZW3ulS+W3NrmYdGnJ07IDDmH8UlUYiFCSPy+uyISNDd
EM3XYoK0T0M6BJGATthdAd+v4dgLZloeV1bDR1OFvhxu1saGH6z1b2KfpQb1Liw8
m+ljrWm89dEhVwtfi2AZ9DtcPx1HR5kmPgcUyZ6LNNz3uJhPG7bp8a3BvQ1kxhC5
2xNksD+0ND7LDolKmOGtFb0UKHEhHwYZpsaf9H/CNwraSxVDEpblq3zpe8tqmVxN
s5d42GhRobkxATvlmg4zMJMT94+m4cv15wqJ7BXGRcujL4vVFnYXom+v2oQxbUWP
i1U/LXuGwW6Bzment254oh3BDlzf4bg8Zk5sasZp1OZ+TtAFdOPgmwpJup8olMQL
zXmPdbZiHvJzEWF54uiY23co7qTJjSoifLHcO9n77o7OTIW5UnpoS0t3YNX4A0Nv
X1DH1PXVEFzDRajKok1uJcSsYpSVIOnH2fkQkpqi50Cd/cPEs5Yqm/cyeP9+WHFZ
2leWnmH2DAmEcQ6zrhJ4QdqD9DDzEcarauIsuTEt6ScH33dE9sPOa5uLLmtIOP5s
XTf/VZGFxpciNK97jOS6YChnEuzymdvOPtWN01vO2mqWBZpmxu2ZU4dr6XR0dbJ3
vd3UkwAmXRxhMCaenLvPk6bvrCbJc81wbXvaRUvsfgodA8quiRlsba/JO93hPx9O
zZFWNxIw7csYRCuc3k2oYEFb2VRQ7nLkUVfOAgAf7HAXXE6iH0D9QHq75ED7jOB5
8HW0aQT1wnpSw6+2jmnofkSPk4ykHQOBaA5XVRflHEm1fm8AiKo4vtGIJsYXYAdI
kOwFUxOuOGu8v1PqOemFWVOdVYbALOgZupEA2KCRheoI+Cvz5yCc0NZKlPrH3X6y
0Rra6ar8QLl042YtdNGTvzTw1eOZsEnzIkseiKm16LblMJH4K5P6aR9TQiWZKlSs
f0xjlXM0+3ls8pQfhOJkTsK2a56KcIIaZ4ziqT6roY+k6QtroybP5VbgrqwxRBIk
JH7eRvDXwscl0K+/DLIdilmUNW+OPlUO7jV8ak6NICXsAomJHsp90T8k+5Fgg4Fb
ZG3ZSGweffc+t+Sx6HW5/c4C54FEg7uBa7Fatvbb8kMyBCHCq9c65IIs/gCj8Hrp
GA8N5nBJ4l5to5gmxXK32h55BR5/cNmgVW6lfNdaAgyBPU9CHTTa1YJU9H528Haj
4X/bBtUwh5exR8X4uiw01MIGiTwiG+uyoJfl/1eWVJV9BQQYF94VEpw8xOwiNsjb
GSapG60F8QmTh/vqenh86dNh8ccUkwCn0IqMe4SNRpm3UYCQcXraJqYXAH2L40re
5jezVUlMD33x74qTSj/oQLkooKawuVsSIBKeRzOB4MxsY797GFNY33lnRqQr3lmE
Ysmi/X+w5gqMG8W+9/61Hilhbfncb9o90nf5SU9xksBe3RUE0xGZV8cOhfCjWlTh
ZOGNNFGtdtQzXh4wZB1f9kh9C2edR8i2GJ7l6Az7QM/eloP9s6aTaFlxk2veDkyq
TpZWW7SLrcO9kso+34R46EWCAggQrNczGtFn8O8N78RO5gF9RfqYZ39Vl6TgDGFK
+6km6IwDvNXXfL8xEqq0Pbi/7CUnqtepdDUTI3wYrQUQQhhEgvZt/avExxeB/z19
8tIl85etA2jnI+ek+bhI1D1N3tQQXZLr4LZkx74xY1GzGXlWemT6gN1Rs7SM8Oh+
I1A1SEhEYfTUpYsh2FXACwCJ0AsW9P2vzOjjgMke2V3Se4u/jnOt9rkHcEwFmIBz
kyx83NV1iNRL2bl+5Q4CM7ZLqMrUzbDCxCkodbc781HdWrZlIFsdSuKVsWRzJ9k9
Y0jLQ3fJIs89F06gDIDWLJLEgeapIiQBCZ7oN3WGzgP1KHRtI+IAQxYYyn0n3hwl
/TGok7JZCklP0TFp16aROFAf782WQHDKkW9PkTvQEy4oXK881NSR6Le4b5PIPlwk
xACHMU/Gtey386B5ah4AuQ4TD6W3qbuXm0Lg65u1vsiWNBzziz06WwBSf4rvkFAX
Ozr/Xn3bM4PbKlYc4facDo2vJKsJgNVC34hYocUdODvOf9UdA5OOiMRqWZdJLE3v
pqM9AXZUoJu5yaGEYxEcqW5CaSwFsSXfDqkhJ/MDeZqHsjyM/kkpR+FuZmMBgH/7
itBCLj1Z0ASTtAzCpOjfCZdOVSh1tc5l5fIqT7OSE2ASqqYP4/SxEK8cVqzgqaCR
mPXwJwpucZJ4ndcTvSMTuG0ROxDddeVQoHnrz+lvt3gPKyeu06GneLARt3r6Ag7p
zNdR3Z02Mlm8I+l/02E46yg6aVqJEQqKasaSE87sGNXmvmTONmw1asOACVvLTIYS
V5gp283mVCxgU2UPNRF50YVsTy+bY1h5Xx8jdaFA4iIPoopVPAH5+zGDR9OSiUuh
LTDPdOz2eSBMtnJKJZPosYHGFzkj/DQ6IEN7Ca4M4v06pVO4zhKMDN+Ue5z9G76k
BZlkOcqs98clbfd1boyN8Jqr8X88baJSWi50bxBIDc2Dw910qF1AUuuLO8NqSqdc
vbb6eg8VppyHHVos140RYJXT3IJvM1CKWtg6UYvm6BiOypypZCfIErDHYCr1ZXm/
M9h6hBTpE5I+xffjLcJphivG9S5TRxuLdGDjsq2yYmwN1cwi5VbCDy2UTGOx/NEs
3bm3vkuHZ1+ovf2fLqlN2fluGzV3/syZQ8DS+DyGKqZx6lf8WwRNA/qUoYeOShvT
UFIEicd/FPx59ALXOKcftjq0LfDby5E1Ok6DefbMzvio/NUYpqOhFsE3qfkQr5YE
8fIvy30JaaN0d9cTuQNj6aYBLR15bbo/zuDEn1okE3p02UpGqGthxOvj6RtwOaSw
9Z8CSLwzxTe75CTvvCsNHO4bs9A0LiXr3yHpEzA5MXnYZmhe0e2uGHoHgpmwbq8D
UKtCrMv4jv7ggnrh7OWNeUCkOr+CWp+GZk5JGonlPEyViiXyMpSxA6Ujl8YEJa2r
dKjddKWoZt38V0m85zpJYkV7VhEAA6DcFbbQfxAyFRYEBmxgkioMbPH6xPQap7FX
ehYFJYV4Bhmr30htZlgeaP5GOkKd9ENAaJHOGlZ0W0M14W5+ZgB/8O6oDiPOTB7L
gkEMdugzMmHinZK9AwmUagoCEdKXKXFCjuqowDzliCpCKAdncp2tZKQQXszxaTMA
mmYWFtleum9AyWlsCcyHJsMV4ejlr88sz5y1L+xF0ZbalSsnfE/FbWIToGAlx2o5
BIaWpPvRtNO7nqfpnLzXWbGXVOjUTcM42TaNZwEyHjuKfyf5/Sf+vXpCkIL2YJnx
JKz/XF6Rh6cmuT0Mt2Dbtu5N7y+vwPTNoj8hS5ID359QzAqfESpLka1FxbfpDHJ2
XOuM+YBBbW7bYRHHlWR7QInHYNtcXpjsG57vDJVfhfhyxTTLqgRaPXFe/GPvvNNh
tZE2XmWfFd9wms15BZR7e+ERI3eKlon/rP6vX07iSGYbsNJeHsDA0hSUc9v+uMOh
n0JX+K/Vg6Bd39SBgIuXew5o1drZnwGfOQU0C03XGOh4NRIKOdNjK45TuCZ//E0J
cfv0pznG8pRriw13KElmKB4XNTZ/hPgldhRYMvs5udxdkDWAysQxWM7o3D14E3FV
nH3A47KSACMQcZS7EQtZ+7egGy5eyzXKC5k5dmWmr3GogDrpmCf8y+hUviBRY2O8
SYv8Q/BxjuQTb1Gl32nCaVtcqjMiO1UwTRQyLzXxMzM5Tf5V1ZfzVPrrbEkYA+o+
Py9IInSEa6mqMC4PbOTARP8c1fb0D7TiVBXzRhKEA5CNdLHl6na6IdSRxDfNawg+
CVwJPMo69aLlvEtiumFxmxOiGbUHBNwAQVKnZePPpKKMNh31WiAqxFgafRznSQ8r
tmvoSd2hBTXOW1e5FoDk2strEdXP8rTV3PB4LM56yJ+LsK8wgdtQPE/a7WmDlzu7
zpVvLwCWl8O6pbO01sQ2yjm96KXSa6fW7I/aYBT+8UuX/zdDJx2vXApymK29GqRs
dO9DEmxjGFwL8gz9uJFT5e+rD90jyx57NoFPW16A2ZQayBwE+hSxOJ239cI5CYJ/
DC+mGHX969Ru9X4VA3D8ZR7sKuIfBFyv+oJUTI51mT/snF+UCas/vgP9GEjy05DC
j9f9UczcT1otl0opdJZX6SWhUEMkvStgwkMiQ1DvEj0Kx0jsl8cfuOFtQ5sI/d8/
NHEtUpyndq45olgz5XCXZlHUvd/V+wwVM4OogHWpYMZu3pW1Ut8lH1vyTyaP0JyR
6tDx5su2PMFJdtPqBN0KkE2hjUurOYVpil54CFxJjJ2pFqUy6CNU91unZ4w49cta
CeVGyVbL99mdjgtjXNXzWa0yVd9AzgiVqFnGhFecK7JvmckHU4c8OlQd8hig4V0E
rrFioxmsgGVn/XdhR+3geAUtxFqJaFVTmQ5pQNORF60iDaWksQHtiYccTYzAB9O+
wUML3j6ss7OyOL6s9nx+CjBt+eAEKlvDWHVdpGUFKkKlqZq4dDAqZ6cqlAXHd81p
276xCZii94puypuNU9MLdn14GAorZ11Jfyr5hkOv7rJC1VvCyjqnffqeERzPWSZ7
VD0KLOb2Gb9rvuvEEQG1zA5NMDL3AWpyLmDepmZpzzgFtbVbk4i5lySRF34e2C5c
Kk9bq5WW33t30o0ODKT4eaSs5eLfMnahNugI6F+/8WsTnXn2iva8DTZ0fdIri17y
0JFrlfUKq/TSeOp6xKTWNMil1TbL+Udq/JAvXTvE1gTfPwEcQnnsGYrYWmdOWw4y
pcjXYVYhzHCidpiimG+Jk1lCyLc0SFHa5osCSgzmDYuqc4hVwYxkXxQIOc1Q2zuu
9h43ozHQZs8qwjRypG8qLGXfRNWX4XanLuE2ND+l/AzAX3uubGg0uLBZXTZnUARd
4cdgIRbgL24eCCr03/qiqw0XjU+WfizVwZXfNjiI4X50saOf9kagVh9qdMF0gsD0
0O+DCfOp7PGm6iScTsM5GQ==
`protect END_PROTECTED