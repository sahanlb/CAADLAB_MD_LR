localparam [NNN1D-1:0][NNN1D-1:0][NNN1D-1:0][BMEMD-1:0][31:0] ROMVAL = {
  32'h3ec3aed4 /* (31, 31, 31) */,
  32'h3d6890ff /* (27, 31, 31) */,
  32'h3d11a602 /* (23, 31, 31) */,
  32'h3d1e42f1 /* (19, 31, 31) */,
  32'h3d167d01 /* (15, 31, 31) */,
  32'h3d151591 /* (11, 31, 31) */,
  32'h3d2402bf /* (7, 31, 31) */,
  32'h3deb372d /* (3, 31, 31) */,
  32'h3d6890ff /* (31, 27, 31) */,
  32'h3d249f29 /* (27, 27, 31) */,
  32'h3d170f20 /* (23, 27, 31) */,
  32'h3d398f3f /* (19, 27, 31) */,
  32'h3d35f880 /* (15, 27, 31) */,
  32'h3d26c9db /* (11, 27, 31) */,
  32'h3d151e01 /* (7, 27, 31) */,
  32'h3d45ae9a /* (3, 27, 31) */,
  32'h3d11a602 /* (31, 23, 31) */,
  32'h3d170f20 /* (27, 23, 31) */,
  32'h3d3ee791 /* (23, 23, 31) */,
  32'h3d8ac476 /* (19, 23, 31) */,
  32'h3d8f3655 /* (15, 23, 31) */,
  32'h3d68852c /* (11, 23, 31) */,
  32'h3d245baa /* (7, 23, 31) */,
  32'h3d126006 /* (3, 23, 31) */,
  32'h3d1e42f1 /* (31, 19, 31) */,
  32'h3d398f3f /* (27, 19, 31) */,
  32'h3d8ac476 /* (23, 19, 31) */,
  32'h3de602d9 /* (19, 19, 31) */,
  32'h3df92d6c /* (15, 19, 31) */,
  32'h3db58f74 /* (11, 19, 31) */,
  32'h3d5c17b6 /* (7, 19, 31) */,
  32'h3d269671 /* (3, 19, 31) */,
  32'h3d167d01 /* (31, 15, 31) */,
  32'h3d35f880 /* (27, 15, 31) */,
  32'h3d8f3655 /* (23, 15, 31) */,
  32'h3df92d6c /* (19, 15, 31) */,
  32'h3e09bd27 /* (15, 15, 31) */,
  32'h3dc031e4 /* (11, 15, 31) */,
  32'h3d5d3ed0 /* (7, 15, 31) */,
  32'h3d202be8 /* (3, 15, 31) */,
  32'h3d151591 /* (31, 11, 31) */,
  32'h3d26c9db /* (27, 11, 31) */,
  32'h3d68852c /* (23, 11, 31) */,
  32'h3db58f74 /* (19, 11, 31) */,
  32'h3dc031e4 /* (15, 11, 31) */,
  32'h3d9352ec /* (11, 11, 31) */,
  32'h3d3efe62 /* (7, 11, 31) */,
  32'h3d1a3ccf /* (3, 11, 31) */,
  32'h3d2402bf /* (31, 7, 31) */,
  32'h3d151e01 /* (27, 7, 31) */,
  32'h3d245baa /* (23, 7, 31) */,
  32'h3d5c17b6 /* (19, 7, 31) */,
  32'h3d5d3ed0 /* (15, 7, 31) */,
  32'h3d3efe62 /* (11, 7, 31) */,
  32'h3d167b79 /* (7, 7, 31) */,
  32'h3d1c3652 /* (3, 7, 31) */,
  32'h3deb372d /* (31, 3, 31) */,
  32'h3d45ae9a /* (27, 3, 31) */,
  32'h3d126006 /* (23, 3, 31) */,
  32'h3d269671 /* (19, 3, 31) */,
  32'h3d202be8 /* (15, 3, 31) */,
  32'h3d1a3ccf /* (11, 3, 31) */,
  32'h3d1c3652 /* (7, 3, 31) */,
  32'h3d960c3c /* (3, 3, 31) */,
  32'h3d6890ff /* (31, 31, 27) */,
  32'h3d249f29 /* (27, 31, 27) */,
  32'h3d170f20 /* (23, 31, 27) */,
  32'h3d398f3f /* (19, 31, 27) */,
  32'h3d35f880 /* (15, 31, 27) */,
  32'h3d26c9db /* (11, 31, 27) */,
  32'h3d151e01 /* (7, 31, 27) */,
  32'h3d45ae9a /* (3, 31, 27) */,
  32'h3d249f29 /* (31, 27, 27) */,
  32'h3d15ac37 /* (27, 27, 27) */,
  32'h3d24f869 /* (23, 27, 27) */,
  32'h3d5ce99d /* (19, 27, 27) */,
  32'h3d5e11d0 /* (15, 27, 27) */,
  32'h3d3fb488 /* (11, 27, 27) */,
  32'h3d170afd /* (7, 27, 27) */,
  32'h3d1ccb4c /* (3, 27, 27) */,
  32'h3d170f20 /* (31, 23, 27) */,
  32'h3d24f869 /* (27, 23, 27) */,
  32'h3d5e7d3b /* (23, 23, 27) */,
  32'h3da95898 /* (19, 23, 27) */,
  32'h3db198fc /* (15, 23, 27) */,
  32'h3d8b02ad /* (11, 23, 27) */,
  32'h3d39ba58 /* (7, 23, 27) */,
  32'h3d1addce /* (3, 23, 27) */,
  32'h3d398f3f /* (31, 19, 27) */,
  32'h3d5ce99d /* (27, 19, 27) */,
  32'h3da95898 /* (23, 19, 27) */,
  32'h3e0f99f2 /* (19, 19, 27) */,
  32'h3e1d0a10 /* (15, 19, 27) */,
  32'h3de04254 /* (11, 19, 27) */,
  32'h3d849ae2 /* (7, 19, 27) */,
  32'h3d4466f8 /* (3, 19, 27) */,
  32'h3d35f880 /* (31, 15, 27) */,
  32'h3d5e11d0 /* (27, 15, 27) */,
  32'h3db198fc /* (23, 15, 27) */,
  32'h3e1d0a10 /* (19, 15, 27) */,
  32'h3e2edbb4 /* (15, 15, 27) */,
  32'h3df05994 /* (11, 15, 27) */,
  32'h3d880917 /* (7, 15, 27) */,
  32'h3d424fe8 /* (3, 15, 27) */,
  32'h3d26c9db /* (31, 11, 27) */,
  32'h3d3fb488 /* (27, 11, 27) */,
  32'h3d8b02ad /* (23, 11, 27) */,
  32'h3de04254 /* (19, 11, 27) */,
  32'h3df05994 /* (15, 11, 27) */,
  32'h3db345e2 /* (11, 11, 27) */,
  32'h3d5ff008 /* (7, 11, 27) */,
  32'h3d2e4aa1 /* (3, 11, 27) */,
  32'h3d151e01 /* (31, 7, 27) */,
  32'h3d170afd /* (27, 7, 27) */,
  32'h3d39ba58 /* (23, 7, 27) */,
  32'h3d849ae2 /* (19, 7, 27) */,
  32'h3d880917 /* (15, 7, 27) */,
  32'h3d5ff008 /* (11, 7, 27) */,
  32'h3d21f168 /* (7, 7, 27) */,
  32'h3d147808 /* (3, 7, 27) */,
  32'h3d45ae9a /* (31, 3, 27) */,
  32'h3d1ccb4c /* (27, 3, 27) */,
  32'h3d1addce /* (23, 3, 27) */,
  32'h3d4466f8 /* (19, 3, 27) */,
  32'h3d424fe8 /* (15, 3, 27) */,
  32'h3d2e4aa1 /* (11, 3, 27) */,
  32'h3d147808 /* (7, 3, 27) */,
  32'h3d314afb /* (3, 3, 27) */,
  32'h3d11a602 /* (31, 31, 23) */,
  32'h3d170f20 /* (27, 31, 23) */,
  32'h3d3ee791 /* (23, 31, 23) */,
  32'h3d8ac476 /* (19, 31, 23) */,
  32'h3d8f3655 /* (15, 31, 23) */,
  32'h3d68852c /* (11, 31, 23) */,
  32'h3d245baa /* (7, 31, 23) */,
  32'h3d126006 /* (3, 31, 23) */,
  32'h3d170f20 /* (31, 27, 23) */,
  32'h3d24f869 /* (27, 27, 23) */,
  32'h3d5e7d3b /* (23, 27, 23) */,
  32'h3da95898 /* (19, 27, 23) */,
  32'h3db198fc /* (15, 27, 23) */,
  32'h3d8b02ad /* (11, 27, 23) */,
  32'h3d39ba58 /* (7, 27, 23) */,
  32'h3d1addce /* (3, 27, 23) */,
  32'h3d3ee791 /* (31, 23, 23) */,
  32'h3d5e7d3b /* (27, 23, 23) */,
  32'h3da4cfbf /* (23, 23, 23) */,
  32'h3e076ebd /* (19, 23, 23) */,
  32'h3e123783 /* (15, 23, 23) */,
  32'h3dd6aa1b /* (11, 23, 23) */,
  32'h3d8354ed /* (7, 23, 23) */,
  32'h3d48821f /* (3, 23, 23) */,
  32'h3d8ac476 /* (31, 19, 23) */,
  32'h3da95898 /* (27, 19, 23) */,
  32'h3e076ebd /* (23, 19, 23) */,
  32'h3e6f82ab /* (19, 19, 23) */,
  32'h3e8557f4 /* (15, 19, 23) */,
  32'h3e37494b /* (11, 19, 23) */,
  32'h3dcf79e9 /* (7, 19, 23) */,
  32'h3d942dc4 /* (3, 19, 23) */,
  32'h3d8f3655 /* (31, 15, 23) */,
  32'h3db198fc /* (27, 15, 23) */,
  32'h3e123783 /* (23, 15, 23) */,
  32'h3e8557f4 /* (19, 15, 23) */,
  32'h3e969108 /* (15, 15, 23) */,
  32'h3e49046a /* (11, 15, 23) */,
  32'h3ddc94c6 /* (7, 15, 23) */,
  32'h3d99caa3 /* (3, 15, 23) */,
  32'h3d68852c /* (31, 11, 23) */,
  32'h3d8b02ad /* (27, 11, 23) */,
  32'h3dd6aa1b /* (23, 11, 23) */,
  32'h3e37494b /* (19, 11, 23) */,
  32'h3e49046a /* (15, 11, 23) */,
  32'h3e0ea5fd /* (11, 11, 23) */,
  32'h3da777c1 /* (7, 11, 23) */,
  32'h3d767d5d /* (3, 11, 23) */,
  32'h3d245baa /* (31, 7, 23) */,
  32'h3d39ba58 /* (27, 7, 23) */,
  32'h3d8354ed /* (23, 7, 23) */,
  32'h3dcf79e9 /* (19, 7, 23) */,
  32'h3ddc94c6 /* (15, 7, 23) */,
  32'h3da777c1 /* (11, 7, 23) */,
  32'h3d563bcb /* (7, 7, 23) */,
  32'h3d2aad03 /* (3, 7, 23) */,
  32'h3d126006 /* (31, 3, 23) */,
  32'h3d1addce /* (27, 3, 23) */,
  32'h3d48821f /* (23, 3, 23) */,
  32'h3d942dc4 /* (19, 3, 23) */,
  32'h3d99caa3 /* (15, 3, 23) */,
  32'h3d767d5d /* (11, 3, 23) */,
  32'h3d2aad03 /* (7, 3, 23) */,
  32'h3d144047 /* (3, 3, 23) */,
  32'h3d1e42f1 /* (31, 31, 19) */,
  32'h3d398f3f /* (27, 31, 19) */,
  32'h3d8ac476 /* (23, 31, 19) */,
  32'h3de602d9 /* (19, 31, 19) */,
  32'h3df92d6c /* (15, 31, 19) */,
  32'h3db58f74 /* (11, 31, 19) */,
  32'h3d5c17b6 /* (7, 31, 19) */,
  32'h3d269671 /* (3, 31, 19) */,
  32'h3d398f3f /* (31, 27, 19) */,
  32'h3d5ce99d /* (27, 27, 19) */,
  32'h3da95898 /* (23, 27, 19) */,
  32'h3e0f99f2 /* (19, 27, 19) */,
  32'h3e1d0a10 /* (15, 27, 19) */,
  32'h3de04254 /* (11, 27, 19) */,
  32'h3d849ae2 /* (7, 27, 19) */,
  32'h3d4466f8 /* (3, 27, 19) */,
  32'h3d8ac476 /* (31, 23, 19) */,
  32'h3da95898 /* (27, 23, 19) */,
  32'h3e076ebd /* (23, 23, 19) */,
  32'h3e6f82ab /* (19, 23, 19) */,
  32'h3e8557f4 /* (15, 23, 19) */,
  32'h3e37494b /* (11, 23, 19) */,
  32'h3dcf79e9 /* (7, 23, 19) */,
  32'h3d942dc4 /* (3, 23, 19) */,
  32'h3de602d9 /* (31, 19, 19) */,
  32'h3e0f99f2 /* (27, 19, 19) */,
  32'h3e6f82ab /* (23, 19, 19) */,
  32'h3edd8ee5 /* (19, 19, 19) */,
  32'h3efbd9fe /* (15, 19, 19) */,
  32'h3ea5d30f /* (11, 19, 19) */,
  32'h3e336d1b /* (7, 19, 19) */,
  32'h3df79892 /* (3, 19, 19) */,
  32'h3df92d6c /* (31, 15, 19) */,
  32'h3e1d0a10 /* (27, 15, 19) */,
  32'h3e8557f4 /* (23, 15, 19) */,
  32'h3efbd9fe /* (19, 15, 19) */,
  32'h3f1092e5 /* (15, 15, 19) */,
  32'h3eba8e90 /* (11, 15, 19) */,
  32'h3e45db44 /* (7, 15, 19) */,
  32'h3e068db8 /* (3, 15, 19) */,
  32'h3db58f74 /* (31, 11, 19) */,
  32'h3de04254 /* (27, 11, 19) */,
  32'h3e37494b /* (23, 11, 19) */,
  32'h3ea5d30f /* (19, 11, 19) */,
  32'h3eba8e90 /* (15, 11, 19) */,
  32'h3e7af74d /* (11, 11, 19) */,
  32'h3e0aca9a /* (7, 11, 19) */,
  32'h3dc2b35d /* (3, 11, 19) */,
  32'h3d5c17b6 /* (31, 7, 19) */,
  32'h3d849ae2 /* (27, 7, 19) */,
  32'h3dcf79e9 /* (23, 7, 19) */,
  32'h3e336d1b /* (19, 7, 19) */,
  32'h3e45db44 /* (15, 7, 19) */,
  32'h3e0aca9a /* (11, 7, 19) */,
  32'h3da0c360 /* (7, 7, 19) */,
  32'h3d69f6ae /* (3, 7, 19) */,
  32'h3d269671 /* (31, 3, 19) */,
  32'h3d4466f8 /* (27, 3, 19) */,
  32'h3d942dc4 /* (23, 3, 19) */,
  32'h3df79892 /* (19, 3, 19) */,
  32'h3e068db8 /* (15, 3, 19) */,
  32'h3dc2b35d /* (11, 3, 19) */,
  32'h3d69f6ae /* (7, 3, 19) */,
  32'h3d2fb3ed /* (3, 3, 19) */,
  32'h3d167d01 /* (31, 31, 15) */,
  32'h3d35f880 /* (27, 31, 15) */,
  32'h3d8f3655 /* (23, 31, 15) */,
  32'h3df92d6c /* (19, 31, 15) */,
  32'h3e09bd27 /* (15, 31, 15) */,
  32'h3dc031e4 /* (11, 31, 15) */,
  32'h3d5d3ed0 /* (7, 31, 15) */,
  32'h3d202be8 /* (3, 31, 15) */,
  32'h3d35f880 /* (31, 27, 15) */,
  32'h3d5e11d0 /* (27, 27, 15) */,
  32'h3db198fc /* (23, 27, 15) */,
  32'h3e1d0a10 /* (19, 27, 15) */,
  32'h3e2edbb4 /* (15, 27, 15) */,
  32'h3df05994 /* (11, 27, 15) */,
  32'h3d880917 /* (7, 27, 15) */,
  32'h3d424fe8 /* (3, 27, 15) */,
  32'h3d8f3655 /* (31, 23, 15) */,
  32'h3db198fc /* (27, 23, 15) */,
  32'h3e123783 /* (23, 23, 15) */,
  32'h3e8557f4 /* (19, 23, 15) */,
  32'h3e969108 /* (15, 23, 15) */,
  32'h3e49046a /* (11, 23, 15) */,
  32'h3ddc94c6 /* (7, 23, 15) */,
  32'h3d99caa3 /* (3, 23, 15) */,
  32'h3df92d6c /* (31, 19, 15) */,
  32'h3e1d0a10 /* (27, 19, 15) */,
  32'h3e8557f4 /* (23, 19, 15) */,
  32'h3efbd9fe /* (19, 19, 15) */,
  32'h3f1092e5 /* (15, 19, 15) */,
  32'h3eba8e90 /* (11, 19, 15) */,
  32'h3e45db44 /* (7, 19, 15) */,
  32'h3e068db8 /* (3, 19, 15) */,
  32'h3e09bd27 /* (31, 15, 15) */,
  32'h3e2edbb4 /* (27, 15, 15) */,
  32'h3e969108 /* (23, 15, 15) */,
  32'h3f1092e5 /* (19, 15, 15) */,
  32'h3f275a64 /* (15, 15, 15) */,
  32'h3ed4648a /* (11, 15, 15) */,
  32'h3e5db918 /* (7, 15, 15) */,
  32'h3e151f83 /* (3, 15, 15) */,
  32'h3dc031e4 /* (31, 11, 15) */,
  32'h3df05994 /* (27, 11, 15) */,
  32'h3e49046a /* (23, 11, 15) */,
  32'h3eba8e90 /* (19, 11, 15) */,
  32'h3ed4648a /* (15, 11, 15) */,
  32'h3e8b66c2 /* (11, 11, 15) */,
  32'h3e165b49 /* (7, 11, 15) */,
  32'h3dceffa6 /* (3, 11, 15) */,
  32'h3d5d3ed0 /* (31, 7, 15) */,
  32'h3d880917 /* (27, 7, 15) */,
  32'h3ddc94c6 /* (23, 7, 15) */,
  32'h3e45db44 /* (19, 7, 15) */,
  32'h3e5db918 /* (15, 7, 15) */,
  32'h3e165b49 /* (11, 7, 15) */,
  32'h3da7bf05 /* (7, 7, 15) */,
  32'h3d6ce397 /* (3, 7, 15) */,
  32'h3d202be8 /* (31, 3, 15) */,
  32'h3d424fe8 /* (27, 3, 15) */,
  32'h3d99caa3 /* (23, 3, 15) */,
  32'h3e068db8 /* (19, 3, 15) */,
  32'h3e151f83 /* (15, 3, 15) */,
  32'h3dceffa6 /* (11, 3, 15) */,
  32'h3d6ce397 /* (7, 3, 15) */,
  32'h3d2aacf2 /* (3, 3, 15) */,
  32'h3d151591 /* (31, 31, 11) */,
  32'h3d26c9db /* (27, 31, 11) */,
  32'h3d68852c /* (23, 31, 11) */,
  32'h3db58f74 /* (19, 31, 11) */,
  32'h3dc031e4 /* (15, 31, 11) */,
  32'h3d9352ec /* (11, 31, 11) */,
  32'h3d3efe62 /* (7, 31, 11) */,
  32'h3d1a3ccf /* (3, 31, 11) */,
  32'h3d26c9db /* (31, 27, 11) */,
  32'h3d3fb488 /* (27, 27, 11) */,
  32'h3d8b02ad /* (23, 27, 11) */,
  32'h3de04254 /* (19, 27, 11) */,
  32'h3df05994 /* (15, 27, 11) */,
  32'h3db345e2 /* (11, 27, 11) */,
  32'h3d5ff008 /* (7, 27, 11) */,
  32'h3d2e4aa1 /* (3, 27, 11) */,
  32'h3d68852c /* (31, 23, 11) */,
  32'h3d8b02ad /* (27, 23, 11) */,
  32'h3dd6aa1b /* (23, 23, 11) */,
  32'h3e37494b /* (19, 23, 11) */,
  32'h3e49046a /* (15, 23, 11) */,
  32'h3e0ea5fd /* (11, 23, 11) */,
  32'h3da777c1 /* (7, 23, 11) */,
  32'h3d767d5d /* (3, 23, 11) */,
  32'h3db58f74 /* (31, 19, 11) */,
  32'h3de04254 /* (27, 19, 11) */,
  32'h3e37494b /* (23, 19, 11) */,
  32'h3ea5d30f /* (19, 19, 11) */,
  32'h3eba8e90 /* (15, 19, 11) */,
  32'h3e7af74d /* (11, 19, 11) */,
  32'h3e0aca9a /* (7, 19, 11) */,
  32'h3dc2b35d /* (3, 19, 11) */,
  32'h3dc031e4 /* (31, 15, 11) */,
  32'h3df05994 /* (27, 15, 11) */,
  32'h3e49046a /* (23, 15, 11) */,
  32'h3eba8e90 /* (19, 15, 11) */,
  32'h3ed4648a /* (15, 15, 11) */,
  32'h3e8b66c2 /* (11, 15, 11) */,
  32'h3e165b49 /* (7, 15, 11) */,
  32'h3dceffa6 /* (3, 15, 11) */,
  32'h3d9352ec /* (31, 11, 11) */,
  32'h3db345e2 /* (27, 11, 11) */,
  32'h3e0ea5fd /* (23, 11, 11) */,
  32'h3e7af74d /* (19, 11, 11) */,
  32'h3e8b66c2 /* (15, 11, 11) */,
  32'h3e4089a2 /* (11, 11, 11) */,
  32'h3ddb1c7f /* (7, 11, 11) */,
  32'h3d9d27e1 /* (3, 11, 11) */,
  32'h3d3efe62 /* (31, 7, 11) */,
  32'h3d5ff008 /* (27, 7, 11) */,
  32'h3da777c1 /* (23, 7, 11) */,
  32'h3e0aca9a /* (19, 7, 11) */,
  32'h3e165b49 /* (15, 7, 11) */,
  32'h3ddb1c7f /* (11, 7, 11) */,
  32'h3d84ce75 /* (7, 7, 11) */,
  32'h3d490aba /* (3, 7, 11) */,
  32'h3d1a3ccf /* (31, 3, 11) */,
  32'h3d2e4aa1 /* (27, 3, 11) */,
  32'h3d767d5d /* (23, 3, 11) */,
  32'h3dc2b35d /* (19, 3, 11) */,
  32'h3dceffa6 /* (15, 3, 11) */,
  32'h3d9d27e1 /* (11, 3, 11) */,
  32'h3d490aba /* (7, 3, 11) */,
  32'h3d202a91 /* (3, 3, 11) */,
  32'h3d2402bf /* (31, 31, 7) */,
  32'h3d151e01 /* (27, 31, 7) */,
  32'h3d245baa /* (23, 31, 7) */,
  32'h3d5c17b6 /* (19, 31, 7) */,
  32'h3d5d3ed0 /* (15, 31, 7) */,
  32'h3d3efe62 /* (11, 31, 7) */,
  32'h3d167b79 /* (7, 31, 7) */,
  32'h3d1c3652 /* (3, 31, 7) */,
  32'h3d151e01 /* (31, 27, 7) */,
  32'h3d170afd /* (27, 27, 7) */,
  32'h3d39ba58 /* (23, 27, 7) */,
  32'h3d849ae2 /* (19, 27, 7) */,
  32'h3d880917 /* (15, 27, 7) */,
  32'h3d5ff008 /* (11, 27, 7) */,
  32'h3d21f168 /* (7, 27, 7) */,
  32'h3d147808 /* (3, 27, 7) */,
  32'h3d245baa /* (31, 23, 7) */,
  32'h3d39ba58 /* (27, 23, 7) */,
  32'h3d8354ed /* (23, 23, 7) */,
  32'h3dcf79e9 /* (19, 23, 7) */,
  32'h3ddc94c6 /* (15, 23, 7) */,
  32'h3da777c1 /* (11, 23, 7) */,
  32'h3d563bcb /* (7, 23, 7) */,
  32'h3d2aad03 /* (3, 23, 7) */,
  32'h3d5c17b6 /* (31, 19, 7) */,
  32'h3d849ae2 /* (27, 19, 7) */,
  32'h3dcf79e9 /* (23, 19, 7) */,
  32'h3e336d1b /* (19, 19, 7) */,
  32'h3e45db44 /* (15, 19, 7) */,
  32'h3e0aca9a /* (11, 19, 7) */,
  32'h3da0c360 /* (7, 19, 7) */,
  32'h3d69f6ae /* (3, 19, 7) */,
  32'h3d5d3ed0 /* (31, 15, 7) */,
  32'h3d880917 /* (27, 15, 7) */,
  32'h3ddc94c6 /* (23, 15, 7) */,
  32'h3e45db44 /* (19, 15, 7) */,
  32'h3e5db918 /* (15, 15, 7) */,
  32'h3e165b49 /* (11, 15, 7) */,
  32'h3da7bf05 /* (7, 15, 7) */,
  32'h3d6ce397 /* (3, 15, 7) */,
  32'h3d3efe62 /* (31, 11, 7) */,
  32'h3d5ff008 /* (27, 11, 7) */,
  32'h3da777c1 /* (23, 11, 7) */,
  32'h3e0aca9a /* (19, 11, 7) */,
  32'h3e165b49 /* (15, 11, 7) */,
  32'h3ddb1c7f /* (11, 11, 7) */,
  32'h3d84ce75 /* (7, 11, 7) */,
  32'h3d490aba /* (3, 11, 7) */,
  32'h3d167b79 /* (31, 7, 7) */,
  32'h3d21f168 /* (27, 7, 7) */,
  32'h3d563bcb /* (23, 7, 7) */,
  32'h3da0c360 /* (19, 7, 7) */,
  32'h3da7bf05 /* (15, 7, 7) */,
  32'h3d84ce75 /* (11, 7, 7) */,
  32'h3d348078 /* (7, 7, 7) */,
  32'h3d1969a9 /* (3, 7, 7) */,
  32'h3d1c3652 /* (31, 3, 7) */,
  32'h3d147808 /* (27, 3, 7) */,
  32'h3d2aad03 /* (23, 3, 7) */,
  32'h3d69f6ae /* (19, 3, 7) */,
  32'h3d6ce397 /* (15, 3, 7) */,
  32'h3d490aba /* (11, 3, 7) */,
  32'h3d1969a9 /* (7, 3, 7) */,
  32'h3d179239 /* (3, 3, 7) */,
  32'h3deb372d /* (31, 31, 3) */,
  32'h3d45ae9a /* (27, 31, 3) */,
  32'h3d126006 /* (23, 31, 3) */,
  32'h3d269671 /* (19, 31, 3) */,
  32'h3d202be8 /* (15, 31, 3) */,
  32'h3d1a3ccf /* (11, 31, 3) */,
  32'h3d1c3652 /* (7, 31, 3) */,
  32'h3d960c3c /* (3, 31, 3) */,
  32'h3d45ae9a /* (31, 27, 3) */,
  32'h3d1ccb4c /* (27, 27, 3) */,
  32'h3d1addce /* (23, 27, 3) */,
  32'h3d4466f8 /* (19, 27, 3) */,
  32'h3d424fe8 /* (15, 27, 3) */,
  32'h3d2e4aa1 /* (11, 27, 3) */,
  32'h3d147808 /* (7, 27, 3) */,
  32'h3d314afb /* (3, 27, 3) */,
  32'h3d126006 /* (31, 23, 3) */,
  32'h3d1addce /* (27, 23, 3) */,
  32'h3d48821f /* (23, 23, 3) */,
  32'h3d942dc4 /* (19, 23, 3) */,
  32'h3d99caa3 /* (15, 23, 3) */,
  32'h3d767d5d /* (11, 23, 3) */,
  32'h3d2aad03 /* (7, 23, 3) */,
  32'h3d144047 /* (3, 23, 3) */,
  32'h3d269671 /* (31, 19, 3) */,
  32'h3d4466f8 /* (27, 19, 3) */,
  32'h3d942dc4 /* (23, 19, 3) */,
  32'h3df79892 /* (19, 19, 3) */,
  32'h3e068db8 /* (15, 19, 3) */,
  32'h3dc2b35d /* (11, 19, 3) */,
  32'h3d69f6ae /* (7, 19, 3) */,
  32'h3d2fb3ed /* (3, 19, 3) */,
  32'h3d202be8 /* (31, 15, 3) */,
  32'h3d424fe8 /* (27, 15, 3) */,
  32'h3d99caa3 /* (23, 15, 3) */,
  32'h3e068db8 /* (19, 15, 3) */,
  32'h3e151f83 /* (15, 15, 3) */,
  32'h3dceffa6 /* (11, 15, 3) */,
  32'h3d6ce397 /* (7, 15, 3) */,
  32'h3d2aacf2 /* (3, 15, 3) */,
  32'h3d1a3ccf /* (31, 11, 3) */,
  32'h3d2e4aa1 /* (27, 11, 3) */,
  32'h3d767d5d /* (23, 11, 3) */,
  32'h3dc2b35d /* (19, 11, 3) */,
  32'h3dceffa6 /* (15, 11, 3) */,
  32'h3d9d27e1 /* (11, 11, 3) */,
  32'h3d490aba /* (7, 11, 3) */,
  32'h3d202a91 /* (3, 11, 3) */,
  32'h3d1c3652 /* (31, 7, 3) */,
  32'h3d147808 /* (27, 7, 3) */,
  32'h3d2aad03 /* (23, 7, 3) */,
  32'h3d69f6ae /* (19, 7, 3) */,
  32'h3d6ce397 /* (15, 7, 3) */,
  32'h3d490aba /* (11, 7, 3) */,
  32'h3d1969a9 /* (7, 7, 3) */,
  32'h3d179239 /* (3, 7, 3) */,
  32'h3d960c3c /* (31, 3, 3) */,
  32'h3d314afb /* (27, 3, 3) */,
  32'h3d144047 /* (23, 3, 3) */,
  32'h3d2fb3ed /* (19, 3, 3) */,
  32'h3d2aacf2 /* (15, 3, 3) */,
  32'h3d202a91 /* (11, 3, 3) */,
  32'h3d179239 /* (7, 3, 3) */,
  32'h3d68b01f /* (3, 3, 3) */,
  32'h3e4aeee2 /* (30, 31, 31) */,
  32'h3d3c9698 /* (26, 31, 31) */,
  32'h3d119771 /* (22, 31, 31) */,
  32'h3d1e0bb6 /* (18, 31, 31) */,
  32'h3d1e0bb6 /* (14, 31, 31) */,
  32'h3d119771 /* (10, 31, 31) */,
  32'h3d3c9698 /* (6, 31, 31) */,
  32'h3e4aeee2 /* (2, 31, 31) */,
  32'h3d59109a /* (30, 27, 31) */,
  32'h3d1a8b5a /* (26, 27, 31) */,
  32'h3d1d9589 /* (22, 27, 31) */,
  32'h3d3c7841 /* (18, 27, 31) */,
  32'h3d3c7841 /* (14, 27, 31) */,
  32'h3d1d9589 /* (10, 27, 31) */,
  32'h3d1a8b5a /* (6, 27, 31) */,
  32'h3d59109a /* (2, 27, 31) */,
  32'h3d11c69f /* (30, 23, 31) */,
  32'h3d1c53e8 /* (26, 23, 31) */,
  32'h3d52081f /* (22, 23, 31) */,
  32'h3d90dff9 /* (18, 23, 31) */,
  32'h3d90dff9 /* (14, 23, 31) */,
  32'h3d52081f /* (10, 23, 31) */,
  32'h3d1c53e8 /* (6, 23, 31) */,
  32'h3d11c69f /* (2, 23, 31) */,
  32'h3d214ba3 /* (30, 19, 31) */,
  32'h3d4876ff /* (26, 19, 31) */,
  32'h3d9e7894 /* (22, 19, 31) */,
  32'h3df65860 /* (18, 19, 31) */,
  32'h3df65860 /* (14, 19, 31) */,
  32'h3d9e7894 /* (10, 19, 31) */,
  32'h3d4876ff /* (6, 19, 31) */,
  32'h3d214ba3 /* (2, 19, 31) */,
  32'h3d1a0745 /* (30, 15, 31) */,
  32'h3d46f53f /* (26, 15, 31) */,
  32'h3da5ac70 /* (22, 15, 31) */,
  32'h3e06d8bb /* (18, 15, 31) */,
  32'h3e06d8bb /* (14, 15, 31) */,
  32'h3da5ac70 /* (10, 15, 31) */,
  32'h3d46f53f /* (6, 15, 31) */,
  32'h3d1a0745 /* (2, 15, 31) */,
  32'h3d16ed42 /* (30, 11, 31) */,
  32'h3d31191b /* (26, 11, 31) */,
  32'h3d829849 /* (22, 11, 31) */,
  32'h3dc01db4 /* (18, 11, 31) */,
  32'h3dc01db4 /* (14, 11, 31) */,
  32'h3d829849 /* (10, 11, 31) */,
  32'h3d31191b /* (6, 11, 31) */,
  32'h3d16ed42 /* (2, 11, 31) */,
  32'h3d20a35e /* (30, 7, 31) */,
  32'h3d146a43 /* (26, 7, 31) */,
  32'h3d305430 /* (22, 7, 31) */,
  32'h3d62906c /* (18, 7, 31) */,
  32'h3d62906c /* (14, 7, 31) */,
  32'h3d305430 /* (10, 7, 31) */,
  32'h3d146a43 /* (6, 7, 31) */,
  32'h3d20a35e /* (2, 7, 31) */,
  32'h3dbfa8df /* (30, 3, 31) */,
  32'h3d2ba889 /* (26, 3, 31) */,
  32'h3d14c0fd /* (22, 3, 31) */,
  32'h3d276174 /* (18, 3, 31) */,
  32'h3d276174 /* (14, 3, 31) */,
  32'h3d14c0fd /* (10, 3, 31) */,
  32'h3d2ba889 /* (6, 3, 31) */,
  32'h3dbfa8df /* (2, 3, 31) */,
  32'h3d59109a /* (30, 31, 27) */,
  32'h3d1a8b5a /* (26, 31, 27) */,
  32'h3d1d9589 /* (22, 31, 27) */,
  32'h3d3c7841 /* (18, 31, 27) */,
  32'h3d3c7841 /* (14, 31, 27) */,
  32'h3d1d9589 /* (10, 31, 27) */,
  32'h3d1a8b5a /* (6, 31, 27) */,
  32'h3d59109a /* (2, 31, 27) */,
  32'h3d213c91 /* (30, 27, 27) */,
  32'h3d14f7ce /* (26, 27, 27) */,
  32'h3d30fc5a /* (22, 27, 27) */,
  32'h3d63687e /* (18, 27, 27) */,
  32'h3d63687e /* (14, 27, 27) */,
  32'h3d30fc5a /* (10, 27, 27) */,
  32'h3d14f7ce /* (6, 27, 27) */,
  32'h3d213c91 /* (2, 27, 27) */,
  32'h3d18622e /* (30, 23, 27) */,
  32'h3d2db0cc /* (26, 23, 27) */,
  32'h3d781ae6 /* (22, 23, 27) */,
  32'h3db24f8e /* (18, 23, 27) */,
  32'h3db24f8e /* (14, 23, 27) */,
  32'h3d781ae6 /* (10, 23, 27) */,
  32'h3d2db0cc /* (6, 23, 27) */,
  32'h3d18622e /* (2, 23, 27) */,
  32'h3d3d84de /* (30, 19, 27) */,
  32'h3d700ffa /* (26, 19, 27) */,
  32'h3dc29629 /* (22, 19, 27) */,
  32'h3e1a8d8c /* (18, 19, 27) */,
  32'h3e1a8d8c /* (14, 19, 27) */,
  32'h3dc29629 /* (10, 19, 27) */,
  32'h3d700ffa /* (6, 19, 27) */,
  32'h3d3d84de /* (2, 19, 27) */,
  32'h3d3a7be5 /* (30, 15, 27) */,
  32'h3d73b16f /* (26, 15, 27) */,
  32'h3dce52e6 /* (22, 15, 27) */,
  32'h3e2a981c /* (18, 15, 27) */,
  32'h3e2a981c /* (14, 15, 27) */,
  32'h3dce52e6 /* (10, 15, 27) */,
  32'h3d73b16f /* (6, 15, 27) */,
  32'h3d3a7be5 /* (2, 15, 27) */,
  32'h3d29823f /* (30, 11, 27) */,
  32'h3d4d9045 /* (26, 11, 27) */,
  32'h3d9d9380 /* (22, 11, 27) */,
  32'h3deed79f /* (18, 11, 27) */,
  32'h3deed79f /* (14, 11, 27) */,
  32'h3d9d9380 /* (10, 11, 27) */,
  32'h3d4d9045 /* (6, 11, 27) */,
  32'h3d29823f /* (2, 11, 27) */,
  32'h3d14b1c0 /* (30, 7, 27) */,
  32'h3d1b2471 /* (26, 7, 27) */,
  32'h3d4b3dc7 /* (22, 7, 27) */,
  32'h3d8a0000 /* (18, 7, 27) */,
  32'h3d8a0000 /* (14, 7, 27) */,
  32'h3d4b3dc7 /* (10, 7, 27) */,
  32'h3d1b2471 /* (6, 7, 27) */,
  32'h3d14b1c0 /* (2, 7, 27) */,
  32'h3d3cd255 /* (30, 3, 27) */,
  32'h3d16d305 /* (26, 3, 27) */,
  32'h3d2344c4 /* (22, 3, 27) */,
  32'h3d487174 /* (18, 3, 27) */,
  32'h3d487174 /* (14, 3, 27) */,
  32'h3d2344c4 /* (10, 3, 27) */,
  32'h3d16d305 /* (6, 3, 27) */,
  32'h3d3cd255 /* (2, 3, 27) */,
  32'h3d11c69f /* (30, 31, 23) */,
  32'h3d1c53e8 /* (26, 31, 23) */,
  32'h3d52081f /* (22, 31, 23) */,
  32'h3d90dff9 /* (18, 31, 23) */,
  32'h3d90dff9 /* (14, 31, 23) */,
  32'h3d52081f /* (10, 31, 23) */,
  32'h3d1c53e8 /* (6, 31, 23) */,
  32'h3d11c69f /* (2, 31, 23) */,
  32'h3d18622e /* (30, 27, 23) */,
  32'h3d2db0cc /* (26, 27, 23) */,
  32'h3d781ae6 /* (22, 27, 23) */,
  32'h3db24f8e /* (18, 27, 23) */,
  32'h3db24f8e /* (14, 27, 23) */,
  32'h3d781ae6 /* (10, 27, 23) */,
  32'h3d2db0cc /* (6, 27, 23) */,
  32'h3d18622e /* (2, 27, 23) */,
  32'h3d42665b /* (30, 23, 23) */,
  32'h3d6fd024 /* (26, 23, 23) */,
  32'h3dbbc730 /* (22, 23, 23) */,
  32'h3e10cac5 /* (18, 23, 23) */,
  32'h3e10cac5 /* (14, 23, 23) */,
  32'h3dbbc730 /* (10, 23, 23) */,
  32'h3d6fd024 /* (6, 23, 23) */,
  32'h3d42665b /* (2, 23, 23) */,
  32'h3d8e358b /* (30, 19, 23) */,
  32'h3db9d5f4 /* (26, 19, 23) */,
  32'h3e1d56b2 /* (22, 19, 23) */,
  32'h3e821787 /* (18, 19, 23) */,
  32'h3e821787 /* (14, 19, 23) */,
  32'h3e1d56b2 /* (10, 19, 23) */,
  32'h3db9d5f4 /* (6, 19, 23) */,
  32'h3d8e358b /* (2, 19, 23) */,
  32'h3d9314c2 /* (30, 15, 23) */,
  32'h3dc42ad0 /* (26, 15, 23) */,
  32'h3e2b3653 /* (22, 15, 23) */,
  32'h3e91e4f8 /* (18, 15, 23) */,
  32'h3e91e4f8 /* (14, 15, 23) */,
  32'h3e2b3653 /* (10, 15, 23) */,
  32'h3dc42ad0 /* (6, 15, 23) */,
  32'h3d9314c2 /* (2, 15, 23) */,
  32'h3d6d9fa3 /* (30, 11, 23) */,
  32'h3d9750ce /* (26, 11, 23) */,
  32'h3df71c69 /* (22, 11, 23) */,
  32'h3e458f30 /* (18, 11, 23) */,
  32'h3e458f30 /* (14, 11, 23) */,
  32'h3df71c69 /* (10, 11, 23) */,
  32'h3d9750ce /* (6, 11, 23) */,
  32'h3d6d9fa3 /* (2, 11, 23) */,
  32'h3d26a1b5 /* (30, 7, 23) */,
  32'h3d45eb5b /* (26, 7, 23) */,
  32'h3d94014f /* (22, 7, 23) */,
  32'h3ddc09d8 /* (18, 7, 23) */,
  32'h3ddc09d8 /* (14, 7, 23) */,
  32'h3d94014f /* (10, 7, 23) */,
  32'h3d45eb5b /* (6, 7, 23) */,
  32'h3d26a1b5 /* (2, 7, 23) */,
  32'h3d12f42a /* (30, 3, 23) */,
  32'h3d215063 /* (26, 3, 23) */,
  32'h3d5dae2c /* (22, 3, 23) */,
  32'h3d9b2a7b /* (18, 3, 23) */,
  32'h3d9b2a7b /* (14, 3, 23) */,
  32'h3d5dae2c /* (10, 3, 23) */,
  32'h3d215063 /* (6, 3, 23) */,
  32'h3d12f42a /* (2, 3, 23) */,
  32'h3d214ba3 /* (30, 31, 19) */,
  32'h3d4876ff /* (26, 31, 19) */,
  32'h3d9e7894 /* (22, 31, 19) */,
  32'h3df65860 /* (18, 31, 19) */,
  32'h3df65860 /* (14, 31, 19) */,
  32'h3d9e7894 /* (10, 31, 19) */,
  32'h3d4876ff /* (6, 31, 19) */,
  32'h3d214ba3 /* (2, 31, 19) */,
  32'h3d3d84de /* (30, 27, 19) */,
  32'h3d700ffa /* (26, 27, 19) */,
  32'h3dc29629 /* (22, 27, 19) */,
  32'h3e1a8d8c /* (18, 27, 19) */,
  32'h3e1a8d8c /* (14, 27, 19) */,
  32'h3dc29629 /* (10, 27, 19) */,
  32'h3d700ffa /* (6, 27, 19) */,
  32'h3d3d84de /* (2, 27, 19) */,
  32'h3d8e358b /* (30, 23, 19) */,
  32'h3db9d5f4 /* (26, 23, 19) */,
  32'h3e1d56b2 /* (22, 23, 19) */,
  32'h3e821787 /* (18, 23, 19) */,
  32'h3e821787 /* (14, 23, 19) */,
  32'h3e1d56b2 /* (10, 23, 19) */,
  32'h3db9d5f4 /* (6, 23, 19) */,
  32'h3d8e358b /* (2, 23, 19) */,
  32'h3dec70da /* (30, 19, 19) */,
  32'h3e1f113d /* (26, 19, 19) */,
  32'h3e8cbae1 /* (22, 19, 19) */,
  32'h3ef33ce4 /* (18, 19, 19) */,
  32'h3ef33ce4 /* (14, 19, 19) */,
  32'h3e8cbae1 /* (10, 19, 19) */,
  32'h3e1f113d /* (6, 19, 19) */,
  32'h3dec70da /* (2, 19, 19) */,
  32'h3e003b1e /* (30, 15, 19) */,
  32'h3e2ea39a /* (26, 15, 19) */,
  32'h3e9d80fb /* (22, 15, 19) */,
  32'h3f0af24f /* (18, 15, 19) */,
  32'h3f0af24f /* (14, 15, 19) */,
  32'h3e9d80fb /* (10, 15, 19) */,
  32'h3e2ea39a /* (6, 15, 19) */,
  32'h3e003b1e /* (2, 15, 19) */,
  32'h3dba5db4 /* (30, 11, 19) */,
  32'h3df74dbc /* (26, 11, 19) */,
  32'h3e562fb1 /* (22, 11, 19) */,
  32'h3eb517ce /* (18, 11, 19) */,
  32'h3eb517ce /* (14, 11, 19) */,
  32'h3e562fb1 /* (10, 11, 19) */,
  32'h3df74dbc /* (6, 11, 19) */,
  32'h3dba5db4 /* (2, 11, 19) */,
  32'h3d6129ae /* (30, 7, 19) */,
  32'h3d90c8a7 /* (26, 7, 19) */,
  32'h3defa49b /* (22, 7, 19) */,
  32'h3e41f14c /* (18, 7, 19) */,
  32'h3e41f14c /* (14, 7, 19) */,
  32'h3defa49b /* (10, 7, 19) */,
  32'h3d90c8a7 /* (6, 7, 19) */,
  32'h3d6129ae /* (2, 7, 19) */,
  32'h3d29e985 /* (30, 3, 19) */,
  32'h3d54a03b /* (26, 3, 19) */,
  32'h3da99659 /* (22, 3, 19) */,
  32'h3e04d0b8 /* (18, 3, 19) */,
  32'h3e04d0b8 /* (14, 3, 19) */,
  32'h3da99659 /* (10, 3, 19) */,
  32'h3d54a03b /* (6, 3, 19) */,
  32'h3d29e985 /* (2, 3, 19) */,
  32'h3d1a0745 /* (30, 31, 15) */,
  32'h3d46f53f /* (26, 31, 15) */,
  32'h3da5ac70 /* (22, 31, 15) */,
  32'h3e06d8bb /* (18, 31, 15) */,
  32'h3e06d8bb /* (14, 31, 15) */,
  32'h3da5ac70 /* (10, 31, 15) */,
  32'h3d46f53f /* (6, 31, 15) */,
  32'h3d1a0745 /* (2, 31, 15) */,
  32'h3d3a7be5 /* (30, 27, 15) */,
  32'h3d73b16f /* (26, 27, 15) */,
  32'h3dce52e6 /* (22, 27, 15) */,
  32'h3e2a981c /* (18, 27, 15) */,
  32'h3e2a981c /* (14, 27, 15) */,
  32'h3dce52e6 /* (10, 27, 15) */,
  32'h3d73b16f /* (6, 27, 15) */,
  32'h3d3a7be5 /* (2, 27, 15) */,
  32'h3d9314c2 /* (30, 23, 15) */,
  32'h3dc42ad0 /* (26, 23, 15) */,
  32'h3e2b3653 /* (22, 23, 15) */,
  32'h3e91e4f8 /* (18, 23, 15) */,
  32'h3e91e4f8 /* (14, 23, 15) */,
  32'h3e2b3653 /* (10, 23, 15) */,
  32'h3dc42ad0 /* (6, 23, 15) */,
  32'h3d9314c2 /* (2, 23, 15) */,
  32'h3e003b1e /* (30, 19, 15) */,
  32'h3e2ea39a /* (26, 19, 15) */,
  32'h3e9d80fb /* (22, 19, 15) */,
  32'h3f0af24f /* (18, 19, 15) */,
  32'h3f0af24f /* (14, 19, 15) */,
  32'h3e9d80fb /* (10, 19, 15) */,
  32'h3e2ea39a /* (6, 19, 15) */,
  32'h3e003b1e /* (2, 19, 15) */,
  32'h3e0de5f8 /* (30, 15, 15) */,
  32'h3e430b11 /* (26, 15, 15) */,
  32'h3eb2925b /* (22, 15, 15) */,
  32'h3f202f9a /* (18, 15, 15) */,
  32'h3f202f9a /* (14, 15, 15) */,
  32'h3eb2925b /* (10, 15, 15) */,
  32'h3e430b11 /* (6, 15, 15) */,
  32'h3e0de5f8 /* (2, 15, 15) */,
  32'h3dc59b81 /* (30, 11, 15) */,
  32'h3e0533d0 /* (26, 11, 15) */,
  32'h3e6c6ac0 /* (22, 11, 15) */,
  32'h3eccf8ff /* (18, 11, 15) */,
  32'h3eccf8ff /* (14, 11, 15) */,
  32'h3e6c6ac0 /* (10, 11, 15) */,
  32'h3e0533d0 /* (6, 11, 15) */,
  32'h3dc59b81 /* (2, 11, 15) */,
  32'h3d62f778 /* (30, 7, 15) */,
  32'h3d95be73 /* (26, 7, 15) */,
  32'h3e009a19 /* (22, 7, 15) */,
  32'h3e57a44b /* (18, 7, 15) */,
  32'h3e57a44b /* (14, 7, 15) */,
  32'h3e009a19 /* (10, 7, 15) */,
  32'h3d95be73 /* (6, 7, 15) */,
  32'h3d62f778 /* (2, 7, 15) */,
  32'h3d240321 /* (30, 3, 15) */,
  32'h3d54ba37 /* (26, 3, 15) */,
  32'h3db22d06 /* (22, 3, 15) */,
  32'h3e11d12f /* (18, 3, 15) */,
  32'h3e11d12f /* (14, 3, 15) */,
  32'h3db22d06 /* (10, 3, 15) */,
  32'h3d54ba37 /* (6, 3, 15) */,
  32'h3d240321 /* (2, 3, 15) */,
  32'h3d16ed42 /* (30, 31, 11) */,
  32'h3d31191b /* (26, 31, 11) */,
  32'h3d829849 /* (22, 31, 11) */,
  32'h3dc01db4 /* (18, 31, 11) */,
  32'h3dc01db4 /* (14, 31, 11) */,
  32'h3d829849 /* (10, 31, 11) */,
  32'h3d31191b /* (6, 31, 11) */,
  32'h3d16ed42 /* (2, 31, 11) */,
  32'h3d29823f /* (30, 27, 11) */,
  32'h3d4d9045 /* (26, 27, 11) */,
  32'h3d9d9380 /* (22, 27, 11) */,
  32'h3deed79f /* (18, 27, 11) */,
  32'h3deed79f /* (14, 27, 11) */,
  32'h3d9d9380 /* (10, 27, 11) */,
  32'h3d4d9045 /* (6, 27, 11) */,
  32'h3d29823f /* (2, 27, 11) */,
  32'h3d6d9fa3 /* (30, 23, 11) */,
  32'h3d9750ce /* (26, 23, 11) */,
  32'h3df71c69 /* (22, 23, 11) */,
  32'h3e458f30 /* (18, 23, 11) */,
  32'h3e458f30 /* (14, 23, 11) */,
  32'h3df71c69 /* (10, 23, 11) */,
  32'h3d9750ce /* (6, 23, 11) */,
  32'h3d6d9fa3 /* (2, 23, 11) */,
  32'h3dba5db4 /* (30, 19, 11) */,
  32'h3df74dbc /* (26, 19, 11) */,
  32'h3e562fb1 /* (22, 19, 11) */,
  32'h3eb517ce /* (18, 19, 11) */,
  32'h3eb517ce /* (14, 19, 11) */,
  32'h3e562fb1 /* (10, 19, 11) */,
  32'h3df74dbc /* (6, 19, 11) */,
  32'h3dba5db4 /* (2, 19, 11) */,
  32'h3dc59b81 /* (30, 15, 11) */,
  32'h3e0533d0 /* (26, 15, 11) */,
  32'h3e6c6ac0 /* (22, 15, 11) */,
  32'h3eccf8ff /* (18, 15, 11) */,
  32'h3eccf8ff /* (14, 15, 11) */,
  32'h3e6c6ac0 /* (10, 15, 11) */,
  32'h3e0533d0 /* (6, 15, 11) */,
  32'h3dc59b81 /* (2, 15, 11) */,
  32'h3d96eb50 /* (30, 11, 11) */,
  32'h3dc480ba /* (26, 11, 11) */,
  32'h3e257fc6 /* (22, 11, 11) */,
  32'h3e882756 /* (18, 11, 11) */,
  32'h3e882756 /* (14, 11, 11) */,
  32'h3e257fc6 /* (10, 11, 11) */,
  32'h3dc480ba /* (6, 11, 11) */,
  32'h3d96eb50 /* (2, 11, 11) */,
  32'h3d42a7b8 /* (30, 7, 11) */,
  32'h3d71ecf9 /* (26, 7, 11) */,
  32'h3dbf3f1d /* (22, 7, 11) */,
  32'h3e14a5c9 /* (18, 7, 11) */,
  32'h3e14a5c9 /* (14, 7, 11) */,
  32'h3dbf3f1d /* (10, 7, 11) */,
  32'h3d71ecf9 /* (6, 7, 11) */,
  32'h3d42a7b8 /* (2, 7, 11) */,
  32'h3d1c5f03 /* (30, 3, 11) */,
  32'h3d39bb76 /* (26, 3, 11) */,
  32'h3d8ae43c /* (22, 3, 11) */,
  32'h3dce7d45 /* (18, 3, 11) */,
  32'h3dce7d45 /* (14, 3, 11) */,
  32'h3d8ae43c /* (10, 3, 11) */,
  32'h3d39bb76 /* (6, 3, 11) */,
  32'h3d1c5f03 /* (2, 3, 11) */,
  32'h3d20a35e /* (30, 31, 7) */,
  32'h3d146a43 /* (26, 31, 7) */,
  32'h3d305430 /* (22, 31, 7) */,
  32'h3d62906c /* (18, 31, 7) */,
  32'h3d62906c /* (14, 31, 7) */,
  32'h3d305430 /* (10, 31, 7) */,
  32'h3d146a43 /* (6, 31, 7) */,
  32'h3d20a35e /* (2, 31, 7) */,
  32'h3d14b1c0 /* (30, 27, 7) */,
  32'h3d1b2471 /* (26, 27, 7) */,
  32'h3d4b3dc7 /* (22, 27, 7) */,
  32'h3d8a0000 /* (18, 27, 7) */,
  32'h3d8a0000 /* (14, 27, 7) */,
  32'h3d4b3dc7 /* (10, 27, 7) */,
  32'h3d1b2471 /* (6, 27, 7) */,
  32'h3d14b1c0 /* (2, 27, 7) */,
  32'h3d26a1b5 /* (30, 23, 7) */,
  32'h3d45eb5b /* (26, 23, 7) */,
  32'h3d94014f /* (22, 23, 7) */,
  32'h3ddc09d8 /* (18, 23, 7) */,
  32'h3ddc09d8 /* (14, 23, 7) */,
  32'h3d94014f /* (10, 23, 7) */,
  32'h3d45eb5b /* (6, 23, 7) */,
  32'h3d26a1b5 /* (2, 23, 7) */,
  32'h3d6129ae /* (30, 19, 7) */,
  32'h3d90c8a7 /* (26, 19, 7) */,
  32'h3defa49b /* (22, 19, 7) */,
  32'h3e41f14c /* (18, 19, 7) */,
  32'h3e41f14c /* (14, 19, 7) */,
  32'h3defa49b /* (10, 19, 7) */,
  32'h3d90c8a7 /* (6, 19, 7) */,
  32'h3d6129ae /* (2, 19, 7) */,
  32'h3d62f778 /* (30, 15, 7) */,
  32'h3d95be73 /* (26, 15, 7) */,
  32'h3e009a19 /* (22, 15, 7) */,
  32'h3e57a44b /* (18, 15, 7) */,
  32'h3e57a44b /* (14, 15, 7) */,
  32'h3e009a19 /* (10, 15, 7) */,
  32'h3d95be73 /* (6, 15, 7) */,
  32'h3d62f778 /* (2, 15, 7) */,
  32'h3d42a7b8 /* (30, 11, 7) */,
  32'h3d71ecf9 /* (26, 11, 7) */,
  32'h3dbf3f1d /* (22, 11, 7) */,
  32'h3e14a5c9 /* (18, 11, 7) */,
  32'h3e14a5c9 /* (14, 11, 7) */,
  32'h3dbf3f1d /* (10, 11, 7) */,
  32'h3d71ecf9 /* (6, 11, 7) */,
  32'h3d42a7b8 /* (2, 11, 7) */,
  32'h3d1777c7 /* (30, 7, 7) */,
  32'h3d29a602 /* (26, 7, 7) */,
  32'h3d6deb12 /* (22, 7, 7) */,
  32'h3da8d240 /* (18, 7, 7) */,
  32'h3da8d240 /* (14, 7, 7) */,
  32'h3d6deb12 /* (10, 7, 7) */,
  32'h3d29a602 /* (6, 7, 7) */,
  32'h3d1777c7 /* (2, 7, 7) */,
  32'h3d1a2949 /* (30, 3, 7) */,
  32'h3d159d44 /* (26, 3, 7) */,
  32'h3d387393 /* (22, 3, 7) */,
  32'h3d71c736 /* (18, 3, 7) */,
  32'h3d71c736 /* (14, 3, 7) */,
  32'h3d387393 /* (10, 3, 7) */,
  32'h3d159d44 /* (6, 3, 7) */,
  32'h3d1a2949 /* (2, 3, 7) */,
  32'h3dbfa8df /* (30, 31, 3) */,
  32'h3d2ba889 /* (26, 31, 3) */,
  32'h3d14c0fd /* (22, 31, 3) */,
  32'h3d276174 /* (18, 31, 3) */,
  32'h3d276174 /* (14, 31, 3) */,
  32'h3d14c0fd /* (10, 31, 3) */,
  32'h3d2ba889 /* (6, 31, 3) */,
  32'h3dbfa8df /* (2, 31, 3) */,
  32'h3d3cd255 /* (30, 27, 3) */,
  32'h3d16d305 /* (26, 27, 3) */,
  32'h3d2344c4 /* (22, 27, 3) */,
  32'h3d487174 /* (18, 27, 3) */,
  32'h3d487174 /* (14, 27, 3) */,
  32'h3d2344c4 /* (10, 27, 3) */,
  32'h3d16d305 /* (6, 27, 3) */,
  32'h3d3cd255 /* (2, 27, 3) */,
  32'h3d12f42a /* (30, 23, 3) */,
  32'h3d215063 /* (26, 23, 3) */,
  32'h3d5dae2c /* (22, 23, 3) */,
  32'h3d9b2a7b /* (18, 23, 3) */,
  32'h3d9b2a7b /* (14, 23, 3) */,
  32'h3d5dae2c /* (10, 23, 3) */,
  32'h3d215063 /* (6, 23, 3) */,
  32'h3d12f42a /* (2, 23, 3) */,
  32'h3d29e985 /* (30, 19, 3) */,
  32'h3d54a03b /* (26, 19, 3) */,
  32'h3da99659 /* (22, 19, 3) */,
  32'h3e04d0b8 /* (18, 19, 3) */,
  32'h3e04d0b8 /* (14, 19, 3) */,
  32'h3da99659 /* (10, 19, 3) */,
  32'h3d54a03b /* (6, 19, 3) */,
  32'h3d29e985 /* (2, 19, 3) */,
  32'h3d240321 /* (30, 15, 3) */,
  32'h3d54ba37 /* (26, 15, 3) */,
  32'h3db22d06 /* (22, 15, 3) */,
  32'h3e11d12f /* (18, 15, 3) */,
  32'h3e11d12f /* (14, 15, 3) */,
  32'h3db22d06 /* (10, 15, 3) */,
  32'h3d54ba37 /* (6, 15, 3) */,
  32'h3d240321 /* (2, 15, 3) */,
  32'h3d1c5f03 /* (30, 11, 3) */,
  32'h3d39bb76 /* (26, 11, 3) */,
  32'h3d8ae43c /* (22, 11, 3) */,
  32'h3dce7d45 /* (18, 11, 3) */,
  32'h3dce7d45 /* (14, 11, 3) */,
  32'h3d8ae43c /* (10, 11, 3) */,
  32'h3d39bb76 /* (6, 11, 3) */,
  32'h3d1c5f03 /* (2, 11, 3) */,
  32'h3d1a2949 /* (30, 7, 3) */,
  32'h3d159d44 /* (26, 7, 3) */,
  32'h3d387393 /* (22, 7, 3) */,
  32'h3d71c736 /* (18, 7, 3) */,
  32'h3d71c736 /* (14, 7, 3) */,
  32'h3d387393 /* (10, 7, 3) */,
  32'h3d159d44 /* (6, 7, 3) */,
  32'h3d1a2949 /* (2, 7, 3) */,
  32'h3d866355 /* (30, 3, 3) */,
  32'h3d211f1b /* (26, 3, 3) */,
  32'h3d18cb02 /* (22, 3, 3) */,
  32'h3d3188e3 /* (18, 3, 3) */,
  32'h3d3188e3 /* (14, 3, 3) */,
  32'h3d18cb02 /* (10, 3, 3) */,
  32'h3d211f1b /* (6, 3, 3) */,
  32'h3d866355 /* (2, 3, 3) */,
  32'h3deb372d /* (29, 31, 31) */,
  32'h3d2402bf /* (25, 31, 31) */,
  32'h3d151591 /* (21, 31, 31) */,
  32'h3d167d01 /* (17, 31, 31) */,
  32'h3d1e42f1 /* (13, 31, 31) */,
  32'h3d11a602 /* (9, 31, 31) */,
  32'h3d6890ff /* (5, 31, 31) */,
  32'h3ec3aed4 /* (1, 31, 31) */,
  32'h3d45ae9a /* (29, 27, 31) */,
  32'h3d151e01 /* (25, 27, 31) */,
  32'h3d26c9db /* (21, 27, 31) */,
  32'h3d35f880 /* (17, 27, 31) */,
  32'h3d398f3f /* (13, 27, 31) */,
  32'h3d170f20 /* (9, 27, 31) */,
  32'h3d249f29 /* (5, 27, 31) */,
  32'h3d6890ff /* (1, 27, 31) */,
  32'h3d126006 /* (29, 23, 31) */,
  32'h3d245baa /* (25, 23, 31) */,
  32'h3d68852c /* (21, 23, 31) */,
  32'h3d8f3655 /* (17, 23, 31) */,
  32'h3d8ac476 /* (13, 23, 31) */,
  32'h3d3ee791 /* (9, 23, 31) */,
  32'h3d170f20 /* (5, 23, 31) */,
  32'h3d11a602 /* (1, 23, 31) */,
  32'h3d269671 /* (29, 19, 31) */,
  32'h3d5c17b6 /* (25, 19, 31) */,
  32'h3db58f74 /* (21, 19, 31) */,
  32'h3df92d6c /* (17, 19, 31) */,
  32'h3de602d9 /* (13, 19, 31) */,
  32'h3d8ac476 /* (9, 19, 31) */,
  32'h3d398f3f /* (5, 19, 31) */,
  32'h3d1e42f1 /* (1, 19, 31) */,
  32'h3d202be8 /* (29, 15, 31) */,
  32'h3d5d3ed0 /* (25, 15, 31) */,
  32'h3dc031e4 /* (21, 15, 31) */,
  32'h3e09bd27 /* (17, 15, 31) */,
  32'h3df92d6c /* (13, 15, 31) */,
  32'h3d8f3655 /* (9, 15, 31) */,
  32'h3d35f880 /* (5, 15, 31) */,
  32'h3d167d01 /* (1, 15, 31) */,
  32'h3d1a3ccf /* (29, 11, 31) */,
  32'h3d3efe62 /* (25, 11, 31) */,
  32'h3d9352ec /* (21, 11, 31) */,
  32'h3dc031e4 /* (17, 11, 31) */,
  32'h3db58f74 /* (13, 11, 31) */,
  32'h3d68852c /* (9, 11, 31) */,
  32'h3d26c9db /* (5, 11, 31) */,
  32'h3d151591 /* (1, 11, 31) */,
  32'h3d1c3652 /* (29, 7, 31) */,
  32'h3d167b79 /* (25, 7, 31) */,
  32'h3d3efe62 /* (21, 7, 31) */,
  32'h3d5d3ed0 /* (17, 7, 31) */,
  32'h3d5c17b6 /* (13, 7, 31) */,
  32'h3d245baa /* (9, 7, 31) */,
  32'h3d151e01 /* (5, 7, 31) */,
  32'h3d2402bf /* (1, 7, 31) */,
  32'h3d960c3c /* (29, 3, 31) */,
  32'h3d1c3652 /* (25, 3, 31) */,
  32'h3d1a3ccf /* (21, 3, 31) */,
  32'h3d202be8 /* (17, 3, 31) */,
  32'h3d269671 /* (13, 3, 31) */,
  32'h3d126006 /* (9, 3, 31) */,
  32'h3d45ae9a /* (5, 3, 31) */,
  32'h3deb372d /* (1, 3, 31) */,
  32'h3d45ae9a /* (29, 31, 27) */,
  32'h3d151e01 /* (25, 31, 27) */,
  32'h3d26c9db /* (21, 31, 27) */,
  32'h3d35f880 /* (17, 31, 27) */,
  32'h3d398f3f /* (13, 31, 27) */,
  32'h3d170f20 /* (9, 31, 27) */,
  32'h3d249f29 /* (5, 31, 27) */,
  32'h3d6890ff /* (1, 31, 27) */,
  32'h3d1ccb4c /* (29, 27, 27) */,
  32'h3d170afd /* (25, 27, 27) */,
  32'h3d3fb488 /* (21, 27, 27) */,
  32'h3d5e11d0 /* (17, 27, 27) */,
  32'h3d5ce99d /* (13, 27, 27) */,
  32'h3d24f869 /* (9, 27, 27) */,
  32'h3d15ac37 /* (5, 27, 27) */,
  32'h3d249f29 /* (1, 27, 27) */,
  32'h3d1addce /* (29, 23, 27) */,
  32'h3d39ba58 /* (25, 23, 27) */,
  32'h3d8b02ad /* (21, 23, 27) */,
  32'h3db198fc /* (17, 23, 27) */,
  32'h3da95898 /* (13, 23, 27) */,
  32'h3d5e7d3b /* (9, 23, 27) */,
  32'h3d24f869 /* (5, 23, 27) */,
  32'h3d170f20 /* (1, 23, 27) */,
  32'h3d4466f8 /* (29, 19, 27) */,
  32'h3d849ae2 /* (25, 19, 27) */,
  32'h3de04254 /* (21, 19, 27) */,
  32'h3e1d0a10 /* (17, 19, 27) */,
  32'h3e0f99f2 /* (13, 19, 27) */,
  32'h3da95898 /* (9, 19, 27) */,
  32'h3d5ce99d /* (5, 19, 27) */,
  32'h3d398f3f /* (1, 19, 27) */,
  32'h3d424fe8 /* (29, 15, 27) */,
  32'h3d880917 /* (25, 15, 27) */,
  32'h3df05994 /* (21, 15, 27) */,
  32'h3e2edbb4 /* (17, 15, 27) */,
  32'h3e1d0a10 /* (13, 15, 27) */,
  32'h3db198fc /* (9, 15, 27) */,
  32'h3d5e11d0 /* (5, 15, 27) */,
  32'h3d35f880 /* (1, 15, 27) */,
  32'h3d2e4aa1 /* (29, 11, 27) */,
  32'h3d5ff008 /* (25, 11, 27) */,
  32'h3db345e2 /* (21, 11, 27) */,
  32'h3df05994 /* (17, 11, 27) */,
  32'h3de04254 /* (13, 11, 27) */,
  32'h3d8b02ad /* (9, 11, 27) */,
  32'h3d3fb488 /* (5, 11, 27) */,
  32'h3d26c9db /* (1, 11, 27) */,
  32'h3d147808 /* (29, 7, 27) */,
  32'h3d21f168 /* (25, 7, 27) */,
  32'h3d5ff008 /* (21, 7, 27) */,
  32'h3d880917 /* (17, 7, 27) */,
  32'h3d849ae2 /* (13, 7, 27) */,
  32'h3d39ba58 /* (9, 7, 27) */,
  32'h3d170afd /* (5, 7, 27) */,
  32'h3d151e01 /* (1, 7, 27) */,
  32'h3d314afb /* (29, 3, 27) */,
  32'h3d147808 /* (25, 3, 27) */,
  32'h3d2e4aa1 /* (21, 3, 27) */,
  32'h3d424fe8 /* (17, 3, 27) */,
  32'h3d4466f8 /* (13, 3, 27) */,
  32'h3d1addce /* (9, 3, 27) */,
  32'h3d1ccb4c /* (5, 3, 27) */,
  32'h3d45ae9a /* (1, 3, 27) */,
  32'h3d126006 /* (29, 31, 23) */,
  32'h3d245baa /* (25, 31, 23) */,
  32'h3d68852c /* (21, 31, 23) */,
  32'h3d8f3655 /* (17, 31, 23) */,
  32'h3d8ac476 /* (13, 31, 23) */,
  32'h3d3ee791 /* (9, 31, 23) */,
  32'h3d170f20 /* (5, 31, 23) */,
  32'h3d11a602 /* (1, 31, 23) */,
  32'h3d1addce /* (29, 27, 23) */,
  32'h3d39ba58 /* (25, 27, 23) */,
  32'h3d8b02ad /* (21, 27, 23) */,
  32'h3db198fc /* (17, 27, 23) */,
  32'h3da95898 /* (13, 27, 23) */,
  32'h3d5e7d3b /* (9, 27, 23) */,
  32'h3d24f869 /* (5, 27, 23) */,
  32'h3d170f20 /* (1, 27, 23) */,
  32'h3d48821f /* (29, 23, 23) */,
  32'h3d8354ed /* (25, 23, 23) */,
  32'h3dd6aa1b /* (21, 23, 23) */,
  32'h3e123783 /* (17, 23, 23) */,
  32'h3e076ebd /* (13, 23, 23) */,
  32'h3da4cfbf /* (9, 23, 23) */,
  32'h3d5e7d3b /* (5, 23, 23) */,
  32'h3d3ee791 /* (1, 23, 23) */,
  32'h3d942dc4 /* (29, 19, 23) */,
  32'h3dcf79e9 /* (25, 19, 23) */,
  32'h3e37494b /* (21, 19, 23) */,
  32'h3e8557f4 /* (17, 19, 23) */,
  32'h3e6f82ab /* (13, 19, 23) */,
  32'h3e076ebd /* (9, 19, 23) */,
  32'h3da95898 /* (5, 19, 23) */,
  32'h3d8ac476 /* (1, 19, 23) */,
  32'h3d99caa3 /* (29, 15, 23) */,
  32'h3ddc94c6 /* (25, 15, 23) */,
  32'h3e49046a /* (21, 15, 23) */,
  32'h3e969108 /* (17, 15, 23) */,
  32'h3e8557f4 /* (13, 15, 23) */,
  32'h3e123783 /* (9, 15, 23) */,
  32'h3db198fc /* (5, 15, 23) */,
  32'h3d8f3655 /* (1, 15, 23) */,
  32'h3d767d5d /* (29, 11, 23) */,
  32'h3da777c1 /* (25, 11, 23) */,
  32'h3e0ea5fd /* (21, 11, 23) */,
  32'h3e49046a /* (17, 11, 23) */,
  32'h3e37494b /* (13, 11, 23) */,
  32'h3dd6aa1b /* (9, 11, 23) */,
  32'h3d8b02ad /* (5, 11, 23) */,
  32'h3d68852c /* (1, 11, 23) */,
  32'h3d2aad03 /* (29, 7, 23) */,
  32'h3d563bcb /* (25, 7, 23) */,
  32'h3da777c1 /* (21, 7, 23) */,
  32'h3ddc94c6 /* (17, 7, 23) */,
  32'h3dcf79e9 /* (13, 7, 23) */,
  32'h3d8354ed /* (9, 7, 23) */,
  32'h3d39ba58 /* (5, 7, 23) */,
  32'h3d245baa /* (1, 7, 23) */,
  32'h3d144047 /* (29, 3, 23) */,
  32'h3d2aad03 /* (25, 3, 23) */,
  32'h3d767d5d /* (21, 3, 23) */,
  32'h3d99caa3 /* (17, 3, 23) */,
  32'h3d942dc4 /* (13, 3, 23) */,
  32'h3d48821f /* (9, 3, 23) */,
  32'h3d1addce /* (5, 3, 23) */,
  32'h3d126006 /* (1, 3, 23) */,
  32'h3d269671 /* (29, 31, 19) */,
  32'h3d5c17b6 /* (25, 31, 19) */,
  32'h3db58f74 /* (21, 31, 19) */,
  32'h3df92d6c /* (17, 31, 19) */,
  32'h3de602d9 /* (13, 31, 19) */,
  32'h3d8ac476 /* (9, 31, 19) */,
  32'h3d398f3f /* (5, 31, 19) */,
  32'h3d1e42f1 /* (1, 31, 19) */,
  32'h3d4466f8 /* (29, 27, 19) */,
  32'h3d849ae2 /* (25, 27, 19) */,
  32'h3de04254 /* (21, 27, 19) */,
  32'h3e1d0a10 /* (17, 27, 19) */,
  32'h3e0f99f2 /* (13, 27, 19) */,
  32'h3da95898 /* (9, 27, 19) */,
  32'h3d5ce99d /* (5, 27, 19) */,
  32'h3d398f3f /* (1, 27, 19) */,
  32'h3d942dc4 /* (29, 23, 19) */,
  32'h3dcf79e9 /* (25, 23, 19) */,
  32'h3e37494b /* (21, 23, 19) */,
  32'h3e8557f4 /* (17, 23, 19) */,
  32'h3e6f82ab /* (13, 23, 19) */,
  32'h3e076ebd /* (9, 23, 19) */,
  32'h3da95898 /* (5, 23, 19) */,
  32'h3d8ac476 /* (1, 23, 19) */,
  32'h3df79892 /* (29, 19, 19) */,
  32'h3e336d1b /* (25, 19, 19) */,
  32'h3ea5d30f /* (21, 19, 19) */,
  32'h3efbd9fe /* (17, 19, 19) */,
  32'h3edd8ee5 /* (13, 19, 19) */,
  32'h3e6f82ab /* (9, 19, 19) */,
  32'h3e0f99f2 /* (5, 19, 19) */,
  32'h3de602d9 /* (1, 19, 19) */,
  32'h3e068db8 /* (29, 15, 19) */,
  32'h3e45db44 /* (25, 15, 19) */,
  32'h3eba8e90 /* (21, 15, 19) */,
  32'h3f1092e5 /* (17, 15, 19) */,
  32'h3efbd9fe /* (13, 15, 19) */,
  32'h3e8557f4 /* (9, 15, 19) */,
  32'h3e1d0a10 /* (5, 15, 19) */,
  32'h3df92d6c /* (1, 15, 19) */,
  32'h3dc2b35d /* (29, 11, 19) */,
  32'h3e0aca9a /* (25, 11, 19) */,
  32'h3e7af74d /* (21, 11, 19) */,
  32'h3eba8e90 /* (17, 11, 19) */,
  32'h3ea5d30f /* (13, 11, 19) */,
  32'h3e37494b /* (9, 11, 19) */,
  32'h3de04254 /* (5, 11, 19) */,
  32'h3db58f74 /* (1, 11, 19) */,
  32'h3d69f6ae /* (29, 7, 19) */,
  32'h3da0c360 /* (25, 7, 19) */,
  32'h3e0aca9a /* (21, 7, 19) */,
  32'h3e45db44 /* (17, 7, 19) */,
  32'h3e336d1b /* (13, 7, 19) */,
  32'h3dcf79e9 /* (9, 7, 19) */,
  32'h3d849ae2 /* (5, 7, 19) */,
  32'h3d5c17b6 /* (1, 7, 19) */,
  32'h3d2fb3ed /* (29, 3, 19) */,
  32'h3d69f6ae /* (25, 3, 19) */,
  32'h3dc2b35d /* (21, 3, 19) */,
  32'h3e068db8 /* (17, 3, 19) */,
  32'h3df79892 /* (13, 3, 19) */,
  32'h3d942dc4 /* (9, 3, 19) */,
  32'h3d4466f8 /* (5, 3, 19) */,
  32'h3d269671 /* (1, 3, 19) */,
  32'h3d202be8 /* (29, 31, 15) */,
  32'h3d5d3ed0 /* (25, 31, 15) */,
  32'h3dc031e4 /* (21, 31, 15) */,
  32'h3e09bd27 /* (17, 31, 15) */,
  32'h3df92d6c /* (13, 31, 15) */,
  32'h3d8f3655 /* (9, 31, 15) */,
  32'h3d35f880 /* (5, 31, 15) */,
  32'h3d167d01 /* (1, 31, 15) */,
  32'h3d424fe8 /* (29, 27, 15) */,
  32'h3d880917 /* (25, 27, 15) */,
  32'h3df05994 /* (21, 27, 15) */,
  32'h3e2edbb4 /* (17, 27, 15) */,
  32'h3e1d0a10 /* (13, 27, 15) */,
  32'h3db198fc /* (9, 27, 15) */,
  32'h3d5e11d0 /* (5, 27, 15) */,
  32'h3d35f880 /* (1, 27, 15) */,
  32'h3d99caa3 /* (29, 23, 15) */,
  32'h3ddc94c6 /* (25, 23, 15) */,
  32'h3e49046a /* (21, 23, 15) */,
  32'h3e969108 /* (17, 23, 15) */,
  32'h3e8557f4 /* (13, 23, 15) */,
  32'h3e123783 /* (9, 23, 15) */,
  32'h3db198fc /* (5, 23, 15) */,
  32'h3d8f3655 /* (1, 23, 15) */,
  32'h3e068db8 /* (29, 19, 15) */,
  32'h3e45db44 /* (25, 19, 15) */,
  32'h3eba8e90 /* (21, 19, 15) */,
  32'h3f1092e5 /* (17, 19, 15) */,
  32'h3efbd9fe /* (13, 19, 15) */,
  32'h3e8557f4 /* (9, 19, 15) */,
  32'h3e1d0a10 /* (5, 19, 15) */,
  32'h3df92d6c /* (1, 19, 15) */,
  32'h3e151f83 /* (29, 15, 15) */,
  32'h3e5db918 /* (25, 15, 15) */,
  32'h3ed4648a /* (21, 15, 15) */,
  32'h3f275a64 /* (17, 15, 15) */,
  32'h3f1092e5 /* (13, 15, 15) */,
  32'h3e969108 /* (9, 15, 15) */,
  32'h3e2edbb4 /* (5, 15, 15) */,
  32'h3e09bd27 /* (1, 15, 15) */,
  32'h3dceffa6 /* (29, 11, 15) */,
  32'h3e165b49 /* (25, 11, 15) */,
  32'h3e8b66c2 /* (21, 11, 15) */,
  32'h3ed4648a /* (17, 11, 15) */,
  32'h3eba8e90 /* (13, 11, 15) */,
  32'h3e49046a /* (9, 11, 15) */,
  32'h3df05994 /* (5, 11, 15) */,
  32'h3dc031e4 /* (1, 11, 15) */,
  32'h3d6ce397 /* (29, 7, 15) */,
  32'h3da7bf05 /* (25, 7, 15) */,
  32'h3e165b49 /* (21, 7, 15) */,
  32'h3e5db918 /* (17, 7, 15) */,
  32'h3e45db44 /* (13, 7, 15) */,
  32'h3ddc94c6 /* (9, 7, 15) */,
  32'h3d880917 /* (5, 7, 15) */,
  32'h3d5d3ed0 /* (1, 7, 15) */,
  32'h3d2aacf2 /* (29, 3, 15) */,
  32'h3d6ce397 /* (25, 3, 15) */,
  32'h3dceffa6 /* (21, 3, 15) */,
  32'h3e151f83 /* (17, 3, 15) */,
  32'h3e068db8 /* (13, 3, 15) */,
  32'h3d99caa3 /* (9, 3, 15) */,
  32'h3d424fe8 /* (5, 3, 15) */,
  32'h3d202be8 /* (1, 3, 15) */,
  32'h3d1a3ccf /* (29, 31, 11) */,
  32'h3d3efe62 /* (25, 31, 11) */,
  32'h3d9352ec /* (21, 31, 11) */,
  32'h3dc031e4 /* (17, 31, 11) */,
  32'h3db58f74 /* (13, 31, 11) */,
  32'h3d68852c /* (9, 31, 11) */,
  32'h3d26c9db /* (5, 31, 11) */,
  32'h3d151591 /* (1, 31, 11) */,
  32'h3d2e4aa1 /* (29, 27, 11) */,
  32'h3d5ff008 /* (25, 27, 11) */,
  32'h3db345e2 /* (21, 27, 11) */,
  32'h3df05994 /* (17, 27, 11) */,
  32'h3de04254 /* (13, 27, 11) */,
  32'h3d8b02ad /* (9, 27, 11) */,
  32'h3d3fb488 /* (5, 27, 11) */,
  32'h3d26c9db /* (1, 27, 11) */,
  32'h3d767d5d /* (29, 23, 11) */,
  32'h3da777c1 /* (25, 23, 11) */,
  32'h3e0ea5fd /* (21, 23, 11) */,
  32'h3e49046a /* (17, 23, 11) */,
  32'h3e37494b /* (13, 23, 11) */,
  32'h3dd6aa1b /* (9, 23, 11) */,
  32'h3d8b02ad /* (5, 23, 11) */,
  32'h3d68852c /* (1, 23, 11) */,
  32'h3dc2b35d /* (29, 19, 11) */,
  32'h3e0aca9a /* (25, 19, 11) */,
  32'h3e7af74d /* (21, 19, 11) */,
  32'h3eba8e90 /* (17, 19, 11) */,
  32'h3ea5d30f /* (13, 19, 11) */,
  32'h3e37494b /* (9, 19, 11) */,
  32'h3de04254 /* (5, 19, 11) */,
  32'h3db58f74 /* (1, 19, 11) */,
  32'h3dceffa6 /* (29, 15, 11) */,
  32'h3e165b49 /* (25, 15, 11) */,
  32'h3e8b66c2 /* (21, 15, 11) */,
  32'h3ed4648a /* (17, 15, 11) */,
  32'h3eba8e90 /* (13, 15, 11) */,
  32'h3e49046a /* (9, 15, 11) */,
  32'h3df05994 /* (5, 15, 11) */,
  32'h3dc031e4 /* (1, 15, 11) */,
  32'h3d9d27e1 /* (29, 11, 11) */,
  32'h3ddb1c7f /* (25, 11, 11) */,
  32'h3e4089a2 /* (21, 11, 11) */,
  32'h3e8b66c2 /* (17, 11, 11) */,
  32'h3e7af74d /* (13, 11, 11) */,
  32'h3e0ea5fd /* (9, 11, 11) */,
  32'h3db345e2 /* (5, 11, 11) */,
  32'h3d9352ec /* (1, 11, 11) */,
  32'h3d490aba /* (29, 7, 11) */,
  32'h3d84ce75 /* (25, 7, 11) */,
  32'h3ddb1c7f /* (21, 7, 11) */,
  32'h3e165b49 /* (17, 7, 11) */,
  32'h3e0aca9a /* (13, 7, 11) */,
  32'h3da777c1 /* (9, 7, 11) */,
  32'h3d5ff008 /* (5, 7, 11) */,
  32'h3d3efe62 /* (1, 7, 11) */,
  32'h3d202a91 /* (29, 3, 11) */,
  32'h3d490aba /* (25, 3, 11) */,
  32'h3d9d27e1 /* (21, 3, 11) */,
  32'h3dceffa6 /* (17, 3, 11) */,
  32'h3dc2b35d /* (13, 3, 11) */,
  32'h3d767d5d /* (9, 3, 11) */,
  32'h3d2e4aa1 /* (5, 3, 11) */,
  32'h3d1a3ccf /* (1, 3, 11) */,
  32'h3d1c3652 /* (29, 31, 7) */,
  32'h3d167b79 /* (25, 31, 7) */,
  32'h3d3efe62 /* (21, 31, 7) */,
  32'h3d5d3ed0 /* (17, 31, 7) */,
  32'h3d5c17b6 /* (13, 31, 7) */,
  32'h3d245baa /* (9, 31, 7) */,
  32'h3d151e01 /* (5, 31, 7) */,
  32'h3d2402bf /* (1, 31, 7) */,
  32'h3d147808 /* (29, 27, 7) */,
  32'h3d21f168 /* (25, 27, 7) */,
  32'h3d5ff008 /* (21, 27, 7) */,
  32'h3d880917 /* (17, 27, 7) */,
  32'h3d849ae2 /* (13, 27, 7) */,
  32'h3d39ba58 /* (9, 27, 7) */,
  32'h3d170afd /* (5, 27, 7) */,
  32'h3d151e01 /* (1, 27, 7) */,
  32'h3d2aad03 /* (29, 23, 7) */,
  32'h3d563bcb /* (25, 23, 7) */,
  32'h3da777c1 /* (21, 23, 7) */,
  32'h3ddc94c6 /* (17, 23, 7) */,
  32'h3dcf79e9 /* (13, 23, 7) */,
  32'h3d8354ed /* (9, 23, 7) */,
  32'h3d39ba58 /* (5, 23, 7) */,
  32'h3d245baa /* (1, 23, 7) */,
  32'h3d69f6ae /* (29, 19, 7) */,
  32'h3da0c360 /* (25, 19, 7) */,
  32'h3e0aca9a /* (21, 19, 7) */,
  32'h3e45db44 /* (17, 19, 7) */,
  32'h3e336d1b /* (13, 19, 7) */,
  32'h3dcf79e9 /* (9, 19, 7) */,
  32'h3d849ae2 /* (5, 19, 7) */,
  32'h3d5c17b6 /* (1, 19, 7) */,
  32'h3d6ce397 /* (29, 15, 7) */,
  32'h3da7bf05 /* (25, 15, 7) */,
  32'h3e165b49 /* (21, 15, 7) */,
  32'h3e5db918 /* (17, 15, 7) */,
  32'h3e45db44 /* (13, 15, 7) */,
  32'h3ddc94c6 /* (9, 15, 7) */,
  32'h3d880917 /* (5, 15, 7) */,
  32'h3d5d3ed0 /* (1, 15, 7) */,
  32'h3d490aba /* (29, 11, 7) */,
  32'h3d84ce75 /* (25, 11, 7) */,
  32'h3ddb1c7f /* (21, 11, 7) */,
  32'h3e165b49 /* (17, 11, 7) */,
  32'h3e0aca9a /* (13, 11, 7) */,
  32'h3da777c1 /* (9, 11, 7) */,
  32'h3d5ff008 /* (5, 11, 7) */,
  32'h3d3efe62 /* (1, 11, 7) */,
  32'h3d1969a9 /* (29, 7, 7) */,
  32'h3d348078 /* (25, 7, 7) */,
  32'h3d84ce75 /* (21, 7, 7) */,
  32'h3da7bf05 /* (17, 7, 7) */,
  32'h3da0c360 /* (13, 7, 7) */,
  32'h3d563bcb /* (9, 7, 7) */,
  32'h3d21f168 /* (5, 7, 7) */,
  32'h3d167b79 /* (1, 7, 7) */,
  32'h3d179239 /* (29, 3, 7) */,
  32'h3d1969a9 /* (25, 3, 7) */,
  32'h3d490aba /* (21, 3, 7) */,
  32'h3d6ce397 /* (17, 3, 7) */,
  32'h3d69f6ae /* (13, 3, 7) */,
  32'h3d2aad03 /* (9, 3, 7) */,
  32'h3d147808 /* (5, 3, 7) */,
  32'h3d1c3652 /* (1, 3, 7) */,
  32'h3d960c3c /* (29, 31, 3) */,
  32'h3d1c3652 /* (25, 31, 3) */,
  32'h3d1a3ccf /* (21, 31, 3) */,
  32'h3d202be8 /* (17, 31, 3) */,
  32'h3d269671 /* (13, 31, 3) */,
  32'h3d126006 /* (9, 31, 3) */,
  32'h3d45ae9a /* (5, 31, 3) */,
  32'h3deb372d /* (1, 31, 3) */,
  32'h3d314afb /* (29, 27, 3) */,
  32'h3d147808 /* (25, 27, 3) */,
  32'h3d2e4aa1 /* (21, 27, 3) */,
  32'h3d424fe8 /* (17, 27, 3) */,
  32'h3d4466f8 /* (13, 27, 3) */,
  32'h3d1addce /* (9, 27, 3) */,
  32'h3d1ccb4c /* (5, 27, 3) */,
  32'h3d45ae9a /* (1, 27, 3) */,
  32'h3d144047 /* (29, 23, 3) */,
  32'h3d2aad03 /* (25, 23, 3) */,
  32'h3d767d5d /* (21, 23, 3) */,
  32'h3d99caa3 /* (17, 23, 3) */,
  32'h3d942dc4 /* (13, 23, 3) */,
  32'h3d48821f /* (9, 23, 3) */,
  32'h3d1addce /* (5, 23, 3) */,
  32'h3d126006 /* (1, 23, 3) */,
  32'h3d2fb3ed /* (29, 19, 3) */,
  32'h3d69f6ae /* (25, 19, 3) */,
  32'h3dc2b35d /* (21, 19, 3) */,
  32'h3e068db8 /* (17, 19, 3) */,
  32'h3df79892 /* (13, 19, 3) */,
  32'h3d942dc4 /* (9, 19, 3) */,
  32'h3d4466f8 /* (5, 19, 3) */,
  32'h3d269671 /* (1, 19, 3) */,
  32'h3d2aacf2 /* (29, 15, 3) */,
  32'h3d6ce397 /* (25, 15, 3) */,
  32'h3dceffa6 /* (21, 15, 3) */,
  32'h3e151f83 /* (17, 15, 3) */,
  32'h3e068db8 /* (13, 15, 3) */,
  32'h3d99caa3 /* (9, 15, 3) */,
  32'h3d424fe8 /* (5, 15, 3) */,
  32'h3d202be8 /* (1, 15, 3) */,
  32'h3d202a91 /* (29, 11, 3) */,
  32'h3d490aba /* (25, 11, 3) */,
  32'h3d9d27e1 /* (21, 11, 3) */,
  32'h3dceffa6 /* (17, 11, 3) */,
  32'h3dc2b35d /* (13, 11, 3) */,
  32'h3d767d5d /* (9, 11, 3) */,
  32'h3d2e4aa1 /* (5, 11, 3) */,
  32'h3d1a3ccf /* (1, 11, 3) */,
  32'h3d179239 /* (29, 7, 3) */,
  32'h3d1969a9 /* (25, 7, 3) */,
  32'h3d490aba /* (21, 7, 3) */,
  32'h3d6ce397 /* (17, 7, 3) */,
  32'h3d69f6ae /* (13, 7, 3) */,
  32'h3d2aad03 /* (9, 7, 3) */,
  32'h3d147808 /* (5, 7, 3) */,
  32'h3d1c3652 /* (1, 7, 3) */,
  32'h3d68b01f /* (29, 3, 3) */,
  32'h3d179239 /* (25, 3, 3) */,
  32'h3d202a91 /* (21, 3, 3) */,
  32'h3d2aacf2 /* (17, 3, 3) */,
  32'h3d2fb3ed /* (13, 3, 3) */,
  32'h3d144047 /* (9, 3, 3) */,
  32'h3d314afb /* (5, 3, 3) */,
  32'h3d960c3c /* (1, 3, 3) */,
  32'h3d9c757b /* (28, 31, 31) */,
  32'h3d1704d7 /* (24, 31, 31) */,
  32'h3d1a2df1 /* (20, 31, 31) */,
  32'h3d067e68 /* (16, 31, 31) */,
  32'h3d1a2df1 /* (12, 31, 31) */,
  32'h3d1704d7 /* (8, 31, 31) */,
  32'h3d9c757b /* (4, 31, 31) */,
  32'h3f10fe39 /* (0, 31, 31) */,
  32'h3d334ee4 /* (28, 27, 31) */,
  32'h3d1412fd /* (24, 27, 31) */,
  32'h3d310ad3 /* (20, 27, 31) */,
  32'h3d24852f /* (16, 27, 31) */,
  32'h3d310ad3 /* (12, 27, 31) */,
  32'h3d1412fd /* (8, 27, 31) */,
  32'h3d334ee4 /* (4, 27, 31) */,
  32'h3d6e9998 /* (0, 27, 31) */,
  32'h3d13f199 /* (28, 23, 31) */,
  32'h3d2fba80 /* (24, 23, 31) */,
  32'h3d803124 /* (20, 23, 31) */,
  32'h3d8420c9 /* (16, 23, 31) */,
  32'h3d803124 /* (12, 23, 31) */,
  32'h3d2fba80 /* (8, 23, 31) */,
  32'h3d13f199 /* (4, 23, 31) */,
  32'h3d11a5c6 /* (0, 23, 31) */,
  32'h3d2e802a /* (28, 19, 31) */,
  32'h3d7573b6 /* (24, 19, 31) */,
  32'h3dce8d02 /* (20, 19, 31) */,
  32'h3deaafef /* (16, 19, 31) */,
  32'h3dce8d02 /* (12, 19, 31) */,
  32'h3d7573b6 /* (8, 19, 31) */,
  32'h3d2e802a /* (4, 19, 31) */,
  32'h3d1d4601 /* (0, 19, 31) */,
  32'h3d294c4b /* (28, 15, 31) */,
  32'h3d7a003f /* (24, 15, 31) */,
  32'h3ddd43c2 /* (20, 15, 31) */,
  32'h3e02e976 /* (16, 15, 31) */,
  32'h3ddd43c2 /* (12, 15, 31) */,
  32'h3d7a003f /* (8, 15, 31) */,
  32'h3d294c4b /* (4, 15, 31) */,
  32'h3d155505 /* (0, 15, 31) */,
  32'h3d1f5dc3 /* (28, 11, 31) */,
  32'h3d513c3d /* (24, 11, 31) */,
  32'h3da53628 /* (20, 11, 31) */,
  32'h3db336e0 /* (16, 11, 31) */,
  32'h3da53628 /* (12, 11, 31) */,
  32'h3d513c3d /* (8, 11, 31) */,
  32'h3d1f5dc3 /* (4, 11, 31) */,
  32'h3d147e90 /* (0, 11, 31) */,
  32'h3d17ff6b /* (28, 7, 31) */,
  32'h3d1bb8b6 /* (24, 7, 31) */,
  32'h3d4ea8e5 /* (20, 7, 31) */,
  32'h3d49f75a /* (16, 7, 31) */,
  32'h3d4ea8e5 /* (12, 7, 31) */,
  32'h3d1bb8b6 /* (8, 7, 31) */,
  32'h3d17ff6b /* (4, 7, 31) */,
  32'h3d25463b /* (0, 7, 31) */,
  32'h3d6eb36b /* (28, 3, 31) */,
  32'h3d146963 /* (24, 3, 31) */,
  32'h3d210eee /* (20, 3, 31) */,
  32'h3d0fbc59 /* (16, 3, 31) */,
  32'h3d210eee /* (12, 3, 31) */,
  32'h3d146963 /* (8, 3, 31) */,
  32'h3d6eb36b /* (4, 3, 31) */,
  32'h3dff9e3f /* (0, 3, 31) */,
  32'h3d334ee4 /* (28, 31, 27) */,
  32'h3d1412fd /* (24, 31, 27) */,
  32'h3d310ad3 /* (20, 31, 27) */,
  32'h3d24852f /* (16, 31, 27) */,
  32'h3d310ad3 /* (12, 31, 27) */,
  32'h3d1412fd /* (8, 31, 27) */,
  32'h3d334ee4 /* (4, 31, 27) */,
  32'h3d6e9998 /* (0, 31, 27) */,
  32'h3d189061 /* (28, 27, 27) */,
  32'h3d1c4d38 /* (24, 27, 27) */,
  32'h3d4f6dfc /* (20, 27, 27) */,
  32'h3d4ab7f7 /* (16, 27, 27) */,
  32'h3d4f6dfc /* (12, 27, 27) */,
  32'h3d1c4d38 /* (8, 27, 27) */,
  32'h3d189061 /* (4, 27, 27) */,
  32'h3d25e3da /* (0, 27, 27) */,
  32'h3d1ee50b /* (28, 23, 27) */,
  32'h3d49c96c /* (24, 23, 27) */,
  32'h3d9af1c2 /* (20, 23, 27) */,
  32'h3da4f2f4 /* (16, 23, 27) */,
  32'h3d9af1c2 /* (12, 23, 27) */,
  32'h3d49c96c /* (8, 23, 27) */,
  32'h3d1ee50b /* (4, 23, 27) */,
  32'h3d16a564 /* (0, 23, 27) */,
  32'h3d4ea6a0 /* (28, 19, 27) */,
  32'h3d94d380 /* (24, 19, 27) */,
  32'h3e00477d /* (20, 19, 27) */,
  32'h3e1486b7 /* (16, 19, 27) */,
  32'h3e00477d /* (12, 19, 27) */,
  32'h3d94d380 /* (8, 19, 27) */,
  32'h3d4ea6a0 /* (4, 19, 27) */,
  32'h3d384488 /* (0, 19, 27) */,
  32'h3d4def9b /* (28, 15, 27) */,
  32'h3d9a5b6b /* (24, 15, 27) */,
  32'h3e0ae903 /* (20, 15, 27) */,
  32'h3e26bbbb /* (16, 15, 27) */,
  32'h3e0ae903 /* (12, 15, 27) */,
  32'h3d9a5b6b /* (8, 15, 27) */,
  32'h3d4def9b /* (4, 15, 27) */,
  32'h3d347f0a /* (0, 15, 27) */,
  32'h3d358341 /* (28, 11, 27) */,
  32'h3d77c8fd /* (24, 11, 27) */,
  32'h3dca9d53 /* (20, 11, 27) */,
  32'h3de14ffa /* (16, 11, 27) */,
  32'h3dca9d53 /* (12, 11, 27) */,
  32'h3d77c8fd /* (8, 11, 27) */,
  32'h3d358341 /* (4, 11, 27) */,
  32'h3d25e815 /* (0, 11, 27) */,
  32'h3d1508af /* (28, 7, 27) */,
  32'h3d2bff3e /* (24, 7, 27) */,
  32'h3d75e4d4 /* (20, 7, 27) */,
  32'h3d7a662c /* (16, 7, 27) */,
  32'h3d75e4d4 /* (12, 7, 27) */,
  32'h3d2bff3e /* (8, 7, 27) */,
  32'h3d1508af /* (4, 7, 27) */,
  32'h3d154f7b /* (0, 7, 27) */,
  32'h3d25f5ce /* (28, 3, 27) */,
  32'h3d15d660 /* (24, 3, 27) */,
  32'h3d3a4ebb /* (20, 3, 27) */,
  32'h3d3046d8 /* (16, 3, 27) */,
  32'h3d3a4ebb /* (12, 3, 27) */,
  32'h3d15d660 /* (8, 3, 27) */,
  32'h3d25f5ce /* (4, 3, 27) */,
  32'h3d490b0e /* (0, 3, 27) */,
  32'h3d13f199 /* (28, 31, 23) */,
  32'h3d2fba80 /* (24, 31, 23) */,
  32'h3d803124 /* (20, 31, 23) */,
  32'h3d8420c9 /* (16, 31, 23) */,
  32'h3d803124 /* (12, 31, 23) */,
  32'h3d2fba80 /* (8, 31, 23) */,
  32'h3d13f199 /* (4, 31, 23) */,
  32'h3d11a5c6 /* (0, 31, 23) */,
  32'h3d1ee50b /* (28, 27, 23) */,
  32'h3d49c96c /* (24, 27, 23) */,
  32'h3d9af1c2 /* (20, 27, 23) */,
  32'h3da4f2f4 /* (16, 27, 23) */,
  32'h3d9af1c2 /* (12, 27, 23) */,
  32'h3d49c96c /* (8, 27, 23) */,
  32'h3d1ee50b /* (4, 27, 23) */,
  32'h3d16a564 /* (0, 27, 23) */,
  32'h3d51a9d2 /* (28, 23, 23) */,
  32'h3d921bde /* (24, 23, 23) */,
  32'h3df3b4f2 /* (20, 23, 23) */,
  32'h3e0981d7 /* (16, 23, 23) */,
  32'h3df3b4f2 /* (12, 23, 23) */,
  32'h3d921bde /* (8, 23, 23) */,
  32'h3d51a9d2 /* (4, 23, 23) */,
  32'h3d3dc47d /* (0, 23, 23) */,
  32'h3d9d0afa /* (28, 19, 23) */,
  32'h3deb6b6d /* (24, 19, 23) */,
  32'h3e53dc51 /* (20, 19, 23) */,
  32'h3e7e4b9d /* (16, 19, 23) */,
  32'h3e53dc51 /* (12, 19, 23) */,
  32'h3deb6b6d /* (8, 19, 23) */,
  32'h3d9d0afa /* (4, 19, 23) */,
  32'h3d89a49e /* (0, 19, 23) */,
  32'h3da3c1ed /* (28, 15, 23) */,
  32'h3dfc30a3 /* (24, 15, 23) */,
  32'h3e6a25fd /* (20, 15, 23) */,
  32'h3e908107 /* (16, 15, 23) */,
  32'h3e6a25fd /* (12, 15, 23) */,
  32'h3dfc30a3 /* (8, 15, 23) */,
  32'h3da3c1ed /* (4, 15, 23) */,
  32'h3d8df2c1 /* (0, 15, 23) */,
  32'h3d81d711 /* (28, 11, 23) */,
  32'h3dbc4d73 /* (24, 11, 23) */,
  32'h3e23781b /* (20, 11, 23) */,
  32'h3e3e5da7 /* (16, 11, 23) */,
  32'h3e23781b /* (12, 11, 23) */,
  32'h3dbc4d73 /* (8, 11, 23) */,
  32'h3d81d711 /* (4, 11, 23) */,
  32'h3d66dac1 /* (0, 11, 23) */,
  32'h3d30de15 /* (28, 7, 23) */,
  32'h3d6b8b35 /* (24, 7, 23) */,
  32'h3dbc51f9 /* (20, 7, 23) */,
  32'h3dce1075 /* (16, 7, 23) */,
  32'h3dbc51f9 /* (12, 7, 23) */,
  32'h3d6b8b35 /* (8, 7, 23) */,
  32'h3d30de15 /* (4, 7, 23) */,
  32'h3d23a039 /* (0, 7, 23) */,
  32'h3d16b5b2 /* (28, 3, 23) */,
  32'h3d37919e /* (24, 3, 23) */,
  32'h3d886b82 /* (20, 3, 23) */,
  32'h3d8e3848 /* (16, 3, 23) */,
  32'h3d886b82 /* (12, 3, 23) */,
  32'h3d37919e /* (8, 3, 23) */,
  32'h3d16b5b2 /* (4, 3, 23) */,
  32'h3d1237a7 /* (0, 3, 23) */,
  32'h3d2e802a /* (28, 31, 19) */,
  32'h3d7573b6 /* (24, 31, 19) */,
  32'h3dce8d02 /* (20, 31, 19) */,
  32'h3deaafef /* (16, 31, 19) */,
  32'h3dce8d02 /* (12, 31, 19) */,
  32'h3d7573b6 /* (8, 31, 19) */,
  32'h3d2e802a /* (4, 31, 19) */,
  32'h3d1d4601 /* (0, 31, 19) */,
  32'h3d4ea6a0 /* (28, 27, 19) */,
  32'h3d94d380 /* (24, 27, 19) */,
  32'h3e00477d /* (20, 27, 19) */,
  32'h3e1486b7 /* (16, 27, 19) */,
  32'h3e00477d /* (12, 27, 19) */,
  32'h3d94d380 /* (8, 27, 19) */,
  32'h3d4ea6a0 /* (4, 27, 19) */,
  32'h3d384488 /* (0, 27, 19) */,
  32'h3d9d0afa /* (28, 23, 19) */,
  32'h3deb6b6d /* (24, 23, 19) */,
  32'h3e53dc51 /* (20, 23, 19) */,
  32'h3e7e4b9d /* (16, 23, 19) */,
  32'h3e53dc51 /* (12, 23, 19) */,
  32'h3deb6b6d /* (8, 23, 19) */,
  32'h3d9d0afa /* (4, 23, 19) */,
  32'h3d89a49e /* (0, 23, 19) */,
  32'h3e0415cb /* (28, 19, 19) */,
  32'h3e4dd3dc /* (24, 19, 19) */,
  32'h3ec1d890 /* (20, 19, 19) */,
  32'h3ef27895 /* (16, 19, 19) */,
  32'h3ec1d890 /* (12, 19, 19) */,
  32'h3e4dd3dc /* (8, 19, 19) */,
  32'h3e0415cb /* (4, 19, 19) */,
  32'h3de3e928 /* (0, 19, 19) */,
  32'h3e0ff4ce /* (28, 15, 19) */,
  32'h3e640ba2 /* (24, 15, 19) */,
  32'h3edb3822 /* (20, 15, 19) */,
  32'h3f0bd969 /* (16, 15, 19) */,
  32'h3edb3822 /* (12, 15, 19) */,
  32'h3e640ba2 /* (8, 15, 19) */,
  32'h3e0ff4ce /* (4, 15, 19) */,
  32'h3df6cc6d /* (0, 15, 19) */,
  32'h3dcf13a3 /* (28, 11, 19) */,
  32'h3e1e607d /* (24, 11, 19) */,
  32'h3e91dfe2 /* (20, 11, 19) */,
  32'h3eb2bd2a /* (16, 11, 19) */,
  32'h3e91dfe2 /* (12, 11, 19) */,
  32'h3e1e607d /* (8, 11, 19) */,
  32'h3dcf13a3 /* (4, 11, 19) */,
  32'h3db3fd83 /* (0, 11, 19) */,
  32'h3d770afc /* (28, 7, 19) */,
  32'h3db56072 /* (24, 7, 19) */,
  32'h3e1f8cbf /* (20, 7, 19) */,
  32'h3e3bd4ee /* (16, 7, 19) */,
  32'h3e1f8cbf /* (12, 7, 19) */,
  32'h3db56072 /* (8, 7, 19) */,
  32'h3d770afc /* (4, 7, 19) */,
  32'h3d5a6fdd /* (0, 7, 19) */,
  32'h3d385879 /* (28, 3, 19) */,
  32'h3d82c188 /* (24, 3, 19) */,
  32'h3dddef48 /* (20, 3, 19) */,
  32'h3dfdd31f /* (16, 3, 19) */,
  32'h3dddef48 /* (12, 3, 19) */,
  32'h3d82c188 /* (8, 3, 19) */,
  32'h3d385879 /* (4, 3, 19) */,
  32'h3d258110 /* (0, 3, 19) */,
  32'h3d294c4b /* (28, 31, 15) */,
  32'h3d7a003f /* (24, 31, 15) */,
  32'h3ddd43c2 /* (20, 31, 15) */,
  32'h3e02e976 /* (16, 31, 15) */,
  32'h3ddd43c2 /* (12, 31, 15) */,
  32'h3d7a003f /* (8, 31, 15) */,
  32'h3d294c4b /* (4, 31, 15) */,
  32'h3d155505 /* (0, 31, 15) */,
  32'h3d4def9b /* (28, 27, 15) */,
  32'h3d9a5b6b /* (24, 27, 15) */,
  32'h3e0ae903 /* (20, 27, 15) */,
  32'h3e26bbbb /* (16, 27, 15) */,
  32'h3e0ae903 /* (12, 27, 15) */,
  32'h3d9a5b6b /* (8, 27, 15) */,
  32'h3d4def9b /* (4, 27, 15) */,
  32'h3d347f0a /* (0, 27, 15) */,
  32'h3da3c1ed /* (28, 23, 15) */,
  32'h3dfc30a3 /* (24, 23, 15) */,
  32'h3e6a25fd /* (20, 23, 15) */,
  32'h3e908107 /* (16, 23, 15) */,
  32'h3e6a25fd /* (12, 23, 15) */,
  32'h3dfc30a3 /* (8, 23, 15) */,
  32'h3da3c1ed /* (4, 23, 15) */,
  32'h3d8df2c1 /* (0, 23, 15) */,
  32'h3e0ff4ce /* (28, 19, 15) */,
  32'h3e640ba2 /* (24, 19, 15) */,
  32'h3edb3822 /* (20, 19, 15) */,
  32'h3f0bd969 /* (16, 19, 15) */,
  32'h3edb3822 /* (12, 19, 15) */,
  32'h3e640ba2 /* (8, 19, 15) */,
  32'h3e0ff4ce /* (4, 19, 15) */,
  32'h3df6cc6d /* (0, 19, 15) */,
  32'h3e1fe07e /* (28, 15, 15) */,
  32'h3e803f85 /* (24, 15, 15) */,
  32'h3efaa119 /* (20, 15, 15) */,
  32'h3f2286f8 /* (16, 15, 15) */,
  32'h3efaa119 /* (12, 15, 15) */,
  32'h3e803f85 /* (8, 15, 15) */,
  32'h3e1fe07e /* (4, 15, 15) */,
  32'h3e086183 /* (0, 15, 15) */,
  32'h3ddcf428 /* (28, 11, 15) */,
  32'h3e2c9c6c /* (24, 11, 15) */,
  32'h3ea31756 /* (20, 11, 15) */,
  32'h3ecca1ac /* (16, 11, 15) */,
  32'h3ea31756 /* (12, 11, 15) */,
  32'h3e2c9c6c /* (8, 11, 15) */,
  32'h3ddcf428 /* (4, 11, 15) */,
  32'h3dbe6d47 /* (0, 11, 15) */,
  32'h3d7b9f11 /* (28, 7, 15) */,
  32'h3dbf0444 /* (24, 7, 15) */,
  32'h3e2e6a71 /* (20, 7, 15) */,
  32'h3e540b9b /* (16, 7, 15) */,
  32'h3e2e6a71 /* (12, 7, 15) */,
  32'h3dbf0444 /* (8, 7, 15) */,
  32'h3d7b9f11 /* (4, 7, 15) */,
  32'h3d5b6048 /* (0, 7, 15) */,
  32'h3d349293 /* (28, 3, 15) */,
  32'h3d8608f0 /* (24, 3, 15) */,
  32'h3deea44d /* (20, 3, 15) */,
  32'h3e0de417 /* (16, 3, 15) */,
  32'h3deea44d /* (12, 3, 15) */,
  32'h3d8608f0 /* (8, 3, 15) */,
  32'h3d349293 /* (4, 3, 15) */,
  32'h3d1eeabe /* (0, 3, 15) */,
  32'h3d1f5dc3 /* (28, 31, 11) */,
  32'h3d513c3d /* (24, 31, 11) */,
  32'h3da53628 /* (20, 31, 11) */,
  32'h3db336e0 /* (16, 31, 11) */,
  32'h3da53628 /* (12, 31, 11) */,
  32'h3d513c3d /* (8, 31, 11) */,
  32'h3d1f5dc3 /* (4, 31, 11) */,
  32'h3d147e90 /* (0, 31, 11) */,
  32'h3d358341 /* (28, 27, 11) */,
  32'h3d77c8fd /* (24, 27, 11) */,
  32'h3dca9d53 /* (20, 27, 11) */,
  32'h3de14ffa /* (16, 27, 11) */,
  32'h3dca9d53 /* (12, 27, 11) */,
  32'h3d77c8fd /* (8, 27, 11) */,
  32'h3d358341 /* (4, 27, 11) */,
  32'h3d25e815 /* (0, 27, 11) */,
  32'h3d81d711 /* (28, 23, 11) */,
  32'h3dbc4d73 /* (24, 23, 11) */,
  32'h3e23781b /* (20, 23, 11) */,
  32'h3e3e5da7 /* (16, 23, 11) */,
  32'h3e23781b /* (12, 23, 11) */,
  32'h3dbc4d73 /* (8, 23, 11) */,
  32'h3d81d711 /* (4, 23, 11) */,
  32'h3d66dac1 /* (0, 23, 11) */,
  32'h3dcf13a3 /* (28, 19, 11) */,
  32'h3e1e607d /* (24, 19, 11) */,
  32'h3e91dfe2 /* (20, 19, 11) */,
  32'h3eb2bd2a /* (16, 19, 11) */,
  32'h3e91dfe2 /* (12, 19, 11) */,
  32'h3e1e607d /* (8, 19, 11) */,
  32'h3dcf13a3 /* (4, 19, 11) */,
  32'h3db3fd83 /* (0, 19, 11) */,
  32'h3ddcf428 /* (28, 15, 11) */,
  32'h3e2c9c6c /* (24, 15, 11) */,
  32'h3ea31756 /* (20, 15, 11) */,
  32'h3ecca1ac /* (16, 15, 11) */,
  32'h3ea31756 /* (12, 15, 11) */,
  32'h3e2c9c6c /* (8, 15, 11) */,
  32'h3ddcf428 /* (4, 15, 11) */,
  32'h3dbe6d47 /* (0, 15, 11) */,
  32'h3da66ad4 /* (28, 11, 11) */,
  32'h3df84bb3 /* (24, 11, 11) */,
  32'h3e5e44ac /* (20, 11, 11) */,
  32'h3e84c8e0 /* (16, 11, 11) */,
  32'h3e5e44ac /* (12, 11, 11) */,
  32'h3df84bb3 /* (8, 11, 11) */,
  32'h3da66ad4 /* (4, 11, 11) */,
  32'h3d922642 /* (0, 11, 11) */,
  32'h3d52976b /* (28, 7, 11) */,
  32'h3d941bce /* (24, 7, 11) */,
  32'h3df94537 /* (20, 7, 11) */,
  32'h3e0d9cf0 /* (16, 7, 11) */,
  32'h3df94537 /* (12, 7, 11) */,
  32'h3d941bce /* (8, 7, 11) */,
  32'h3d52976b /* (4, 7, 11) */,
  32'h3d3dcd22 /* (0, 7, 11) */,
  32'h3d25fa09 /* (28, 3, 11) */,
  32'h3d5d0a38 /* (24, 3, 11) */,
  32'h3db0b965 /* (20, 3, 11) */,
  32'h3dc1602b /* (16, 3, 11) */,
  32'h3db0b965 /* (12, 3, 11) */,
  32'h3d5d0a38 /* (8, 3, 11) */,
  32'h3d25fa09 /* (4, 3, 11) */,
  32'h3d198ce9 /* (0, 3, 11) */,
  32'h3d17ff6b /* (28, 31, 7) */,
  32'h3d1bb8b6 /* (24, 31, 7) */,
  32'h3d4ea8e5 /* (20, 31, 7) */,
  32'h3d49f75a /* (16, 31, 7) */,
  32'h3d4ea8e5 /* (12, 31, 7) */,
  32'h3d1bb8b6 /* (8, 31, 7) */,
  32'h3d17ff6b /* (4, 31, 7) */,
  32'h3d25463b /* (0, 31, 7) */,
  32'h3d1508af /* (28, 27, 7) */,
  32'h3d2bff3e /* (24, 27, 7) */,
  32'h3d75e4d4 /* (20, 27, 7) */,
  32'h3d7a662c /* (16, 27, 7) */,
  32'h3d75e4d4 /* (12, 27, 7) */,
  32'h3d2bff3e /* (8, 27, 7) */,
  32'h3d1508af /* (4, 27, 7) */,
  32'h3d154f7b /* (0, 27, 7) */,
  32'h3d30de15 /* (28, 23, 7) */,
  32'h3d6b8b35 /* (24, 23, 7) */,
  32'h3dbc51f9 /* (20, 23, 7) */,
  32'h3dce1075 /* (16, 23, 7) */,
  32'h3dbc51f9 /* (12, 23, 7) */,
  32'h3d6b8b35 /* (8, 23, 7) */,
  32'h3d30de15 /* (4, 23, 7) */,
  32'h3d23a039 /* (0, 23, 7) */,
  32'h3d770afc /* (28, 19, 7) */,
  32'h3db56072 /* (24, 19, 7) */,
  32'h3e1f8cbf /* (20, 19, 7) */,
  32'h3e3bd4ee /* (16, 19, 7) */,
  32'h3e1f8cbf /* (12, 19, 7) */,
  32'h3db56072 /* (8, 19, 7) */,
  32'h3d770afc /* (4, 19, 7) */,
  32'h3d5a6fdd /* (0, 19, 7) */,
  32'h3d7b9f11 /* (28, 15, 7) */,
  32'h3dbf0444 /* (24, 15, 7) */,
  32'h3e2e6a71 /* (20, 15, 7) */,
  32'h3e540b9b /* (16, 15, 7) */,
  32'h3e2e6a71 /* (12, 15, 7) */,
  32'h3dbf0444 /* (8, 15, 7) */,
  32'h3d7b9f11 /* (4, 15, 7) */,
  32'h3d5b6048 /* (0, 15, 7) */,
  32'h3d52976b /* (28, 11, 7) */,
  32'h3d941bce /* (24, 11, 7) */,
  32'h3df94537 /* (20, 11, 7) */,
  32'h3e0d9cf0 /* (16, 11, 7) */,
  32'h3df94537 /* (12, 11, 7) */,
  32'h3d941bce /* (8, 11, 7) */,
  32'h3d52976b /* (4, 11, 7) */,
  32'h3d3dcd22 /* (0, 11, 7) */,
  32'h3d1cbb18 /* (28, 7, 7) */,
  32'h3d432bf1 /* (24, 7, 7) */,
  32'h3d938890 /* (20, 7, 7) */,
  32'h3d9b7830 /* (16, 7, 7) */,
  32'h3d938890 /* (12, 7, 7) */,
  32'h3d432bf1 /* (8, 7, 7) */,
  32'h3d1cbb18 /* (4, 7, 7) */,
  32'h3d162f74 /* (0, 7, 7) */,
  32'h3d155fa4 /* (28, 3, 7) */,
  32'h3d2054cd /* (24, 3, 7) */,
  32'h3d5ab0e1 /* (20, 3, 7) */,
  32'h3d58de26 /* (16, 3, 7) */,
  32'h3d5ab0e1 /* (12, 3, 7) */,
  32'h3d2054cd /* (8, 3, 7) */,
  32'h3d155fa4 /* (4, 3, 7) */,
  32'h3d1cfd70 /* (0, 3, 7) */,
  32'h3d6eb36b /* (28, 31, 3) */,
  32'h3d146963 /* (24, 31, 3) */,
  32'h3d210eee /* (20, 31, 3) */,
  32'h3d0fbc59 /* (16, 31, 3) */,
  32'h3d210eee /* (12, 31, 3) */,
  32'h3d146963 /* (8, 31, 3) */,
  32'h3d6eb36b /* (4, 31, 3) */,
  32'h3dff9e3f /* (0, 31, 3) */,
  32'h3d25f5ce /* (28, 27, 3) */,
  32'h3d15d660 /* (24, 27, 3) */,
  32'h3d3a4ebb /* (20, 27, 3) */,
  32'h3d3046d8 /* (16, 27, 3) */,
  32'h3d3a4ebb /* (12, 27, 3) */,
  32'h3d15d660 /* (8, 27, 3) */,
  32'h3d25f5ce /* (4, 27, 3) */,
  32'h3d490b0e /* (0, 27, 3) */,
  32'h3d16b5b2 /* (28, 23, 3) */,
  32'h3d37919e /* (24, 23, 3) */,
  32'h3d886b82 /* (20, 23, 3) */,
  32'h3d8e3848 /* (16, 23, 3) */,
  32'h3d886b82 /* (12, 23, 3) */,
  32'h3d37919e /* (8, 23, 3) */,
  32'h3d16b5b2 /* (4, 23, 3) */,
  32'h3d1237a7 /* (0, 23, 3) */,
  32'h3d385879 /* (28, 19, 3) */,
  32'h3d82c188 /* (24, 19, 3) */,
  32'h3dddef48 /* (20, 19, 3) */,
  32'h3dfdd31f /* (16, 19, 3) */,
  32'h3dddef48 /* (12, 19, 3) */,
  32'h3d82c188 /* (8, 19, 3) */,
  32'h3d385879 /* (4, 19, 3) */,
  32'h3d258110 /* (0, 19, 3) */,
  32'h3d349293 /* (28, 15, 3) */,
  32'h3d8608f0 /* (24, 15, 3) */,
  32'h3deea44d /* (20, 15, 3) */,
  32'h3e0de417 /* (16, 15, 3) */,
  32'h3deea44d /* (12, 15, 3) */,
  32'h3d8608f0 /* (8, 15, 3) */,
  32'h3d349293 /* (4, 15, 3) */,
  32'h3d1eeabe /* (0, 15, 3) */,
  32'h3d25fa09 /* (28, 11, 3) */,
  32'h3d5d0a38 /* (24, 11, 3) */,
  32'h3db0b965 /* (20, 11, 3) */,
  32'h3dc1602b /* (16, 11, 3) */,
  32'h3db0b965 /* (12, 11, 3) */,
  32'h3d5d0a38 /* (8, 11, 3) */,
  32'h3d25fa09 /* (4, 11, 3) */,
  32'h3d198ce9 /* (0, 11, 3) */,
  32'h3d155fa4 /* (28, 7, 3) */,
  32'h3d2054cd /* (24, 7, 3) */,
  32'h3d5ab0e1 /* (20, 7, 3) */,
  32'h3d58de26 /* (16, 7, 3) */,
  32'h3d5ab0e1 /* (12, 7, 3) */,
  32'h3d2054cd /* (8, 7, 3) */,
  32'h3d155fa4 /* (4, 7, 3) */,
  32'h3d1cfd70 /* (0, 7, 3) */,
  32'h3d4920d0 /* (28, 3, 3) */,
  32'h3d1392fe /* (24, 3, 3) */,
  32'h3d28b308 /* (20, 3, 3) */,
  32'h3d19c07a /* (16, 3, 3) */,
  32'h3d28b308 /* (12, 3, 3) */,
  32'h3d1392fe /* (8, 3, 3) */,
  32'h3d4920d0 /* (4, 3, 3) */,
  32'h3d9c797c /* (0, 3, 3) */,
  32'h3e4aeee2 /* (31, 30, 31) */,
  32'h3d59109a /* (27, 30, 31) */,
  32'h3d11c69f /* (23, 30, 31) */,
  32'h3d214ba3 /* (19, 30, 31) */,
  32'h3d1a0745 /* (15, 30, 31) */,
  32'h3d16ed42 /* (11, 30, 31) */,
  32'h3d20a35e /* (7, 30, 31) */,
  32'h3dbfa8df /* (3, 30, 31) */,
  32'h3d3c9698 /* (31, 26, 31) */,
  32'h3d1a8b5a /* (27, 26, 31) */,
  32'h3d1c53e8 /* (23, 26, 31) */,
  32'h3d4876ff /* (19, 26, 31) */,
  32'h3d46f53f /* (15, 26, 31) */,
  32'h3d31191b /* (11, 26, 31) */,
  32'h3d146a43 /* (7, 26, 31) */,
  32'h3d2ba889 /* (3, 26, 31) */,
  32'h3d119771 /* (31, 22, 31) */,
  32'h3d1d9589 /* (27, 22, 31) */,
  32'h3d52081f /* (23, 22, 31) */,
  32'h3d9e7894 /* (19, 22, 31) */,
  32'h3da5ac70 /* (15, 22, 31) */,
  32'h3d829849 /* (11, 22, 31) */,
  32'h3d305430 /* (7, 22, 31) */,
  32'h3d14c0fd /* (3, 22, 31) */,
  32'h3d1e0bb6 /* (31, 18, 31) */,
  32'h3d3c7841 /* (27, 18, 31) */,
  32'h3d90dff9 /* (23, 18, 31) */,
  32'h3df65860 /* (19, 18, 31) */,
  32'h3e06d8bb /* (15, 18, 31) */,
  32'h3dc01db4 /* (11, 18, 31) */,
  32'h3d62906c /* (7, 18, 31) */,
  32'h3d276174 /* (3, 18, 31) */,
  32'h3d1e0bb6 /* (31, 14, 31) */,
  32'h3d3c7841 /* (27, 14, 31) */,
  32'h3d90dff9 /* (23, 14, 31) */,
  32'h3df65860 /* (19, 14, 31) */,
  32'h3e06d8bb /* (15, 14, 31) */,
  32'h3dc01db4 /* (11, 14, 31) */,
  32'h3d62906c /* (7, 14, 31) */,
  32'h3d276174 /* (3, 14, 31) */,
  32'h3d119771 /* (31, 10, 31) */,
  32'h3d1d9589 /* (27, 10, 31) */,
  32'h3d52081f /* (23, 10, 31) */,
  32'h3d9e7894 /* (19, 10, 31) */,
  32'h3da5ac70 /* (15, 10, 31) */,
  32'h3d829849 /* (11, 10, 31) */,
  32'h3d305430 /* (7, 10, 31) */,
  32'h3d14c0fd /* (3, 10, 31) */,
  32'h3d3c9698 /* (31, 6, 31) */,
  32'h3d1a8b5a /* (27, 6, 31) */,
  32'h3d1c53e8 /* (23, 6, 31) */,
  32'h3d4876ff /* (19, 6, 31) */,
  32'h3d46f53f /* (15, 6, 31) */,
  32'h3d31191b /* (11, 6, 31) */,
  32'h3d146a43 /* (7, 6, 31) */,
  32'h3d2ba889 /* (3, 6, 31) */,
  32'h3e4aeee2 /* (31, 2, 31) */,
  32'h3d59109a /* (27, 2, 31) */,
  32'h3d11c69f /* (23, 2, 31) */,
  32'h3d214ba3 /* (19, 2, 31) */,
  32'h3d1a0745 /* (15, 2, 31) */,
  32'h3d16ed42 /* (11, 2, 31) */,
  32'h3d20a35e /* (7, 2, 31) */,
  32'h3dbfa8df /* (3, 2, 31) */,
  32'h3d59109a /* (31, 30, 27) */,
  32'h3d213c91 /* (27, 30, 27) */,
  32'h3d18622e /* (23, 30, 27) */,
  32'h3d3d84de /* (19, 30, 27) */,
  32'h3d3a7be5 /* (15, 30, 27) */,
  32'h3d29823f /* (11, 30, 27) */,
  32'h3d14b1c0 /* (7, 30, 27) */,
  32'h3d3cd255 /* (3, 30, 27) */,
  32'h3d1a8b5a /* (31, 26, 27) */,
  32'h3d14f7ce /* (27, 26, 27) */,
  32'h3d2db0cc /* (23, 26, 27) */,
  32'h3d700ffa /* (19, 26, 27) */,
  32'h3d73b16f /* (15, 26, 27) */,
  32'h3d4d9045 /* (11, 26, 27) */,
  32'h3d1b2471 /* (7, 26, 27) */,
  32'h3d16d305 /* (3, 26, 27) */,
  32'h3d1d9589 /* (31, 22, 27) */,
  32'h3d30fc5a /* (27, 22, 27) */,
  32'h3d781ae6 /* (23, 22, 27) */,
  32'h3dc29629 /* (19, 22, 27) */,
  32'h3dce52e6 /* (15, 22, 27) */,
  32'h3d9d9380 /* (11, 22, 27) */,
  32'h3d4b3dc7 /* (7, 22, 27) */,
  32'h3d2344c4 /* (3, 22, 27) */,
  32'h3d3c7841 /* (31, 18, 27) */,
  32'h3d63687e /* (27, 18, 27) */,
  32'h3db24f8e /* (23, 18, 27) */,
  32'h3e1a8d8c /* (19, 18, 27) */,
  32'h3e2a981c /* (15, 18, 27) */,
  32'h3deed79f /* (11, 18, 27) */,
  32'h3d8a0000 /* (7, 18, 27) */,
  32'h3d487174 /* (3, 18, 27) */,
  32'h3d3c7841 /* (31, 14, 27) */,
  32'h3d63687e /* (27, 14, 27) */,
  32'h3db24f8e /* (23, 14, 27) */,
  32'h3e1a8d8c /* (19, 14, 27) */,
  32'h3e2a981c /* (15, 14, 27) */,
  32'h3deed79f /* (11, 14, 27) */,
  32'h3d8a0000 /* (7, 14, 27) */,
  32'h3d487174 /* (3, 14, 27) */,
  32'h3d1d9589 /* (31, 10, 27) */,
  32'h3d30fc5a /* (27, 10, 27) */,
  32'h3d781ae6 /* (23, 10, 27) */,
  32'h3dc29629 /* (19, 10, 27) */,
  32'h3dce52e6 /* (15, 10, 27) */,
  32'h3d9d9380 /* (11, 10, 27) */,
  32'h3d4b3dc7 /* (7, 10, 27) */,
  32'h3d2344c4 /* (3, 10, 27) */,
  32'h3d1a8b5a /* (31, 6, 27) */,
  32'h3d14f7ce /* (27, 6, 27) */,
  32'h3d2db0cc /* (23, 6, 27) */,
  32'h3d700ffa /* (19, 6, 27) */,
  32'h3d73b16f /* (15, 6, 27) */,
  32'h3d4d9045 /* (11, 6, 27) */,
  32'h3d1b2471 /* (7, 6, 27) */,
  32'h3d16d305 /* (3, 6, 27) */,
  32'h3d59109a /* (31, 2, 27) */,
  32'h3d213c91 /* (27, 2, 27) */,
  32'h3d18622e /* (23, 2, 27) */,
  32'h3d3d84de /* (19, 2, 27) */,
  32'h3d3a7be5 /* (15, 2, 27) */,
  32'h3d29823f /* (11, 2, 27) */,
  32'h3d14b1c0 /* (7, 2, 27) */,
  32'h3d3cd255 /* (3, 2, 27) */,
  32'h3d11c69f /* (31, 30, 23) */,
  32'h3d18622e /* (27, 30, 23) */,
  32'h3d42665b /* (23, 30, 23) */,
  32'h3d8e358b /* (19, 30, 23) */,
  32'h3d9314c2 /* (15, 30, 23) */,
  32'h3d6d9fa3 /* (11, 30, 23) */,
  32'h3d26a1b5 /* (7, 30, 23) */,
  32'h3d12f42a /* (3, 30, 23) */,
  32'h3d1c53e8 /* (31, 26, 23) */,
  32'h3d2db0cc /* (27, 26, 23) */,
  32'h3d6fd024 /* (23, 26, 23) */,
  32'h3db9d5f4 /* (19, 26, 23) */,
  32'h3dc42ad0 /* (15, 26, 23) */,
  32'h3d9750ce /* (11, 26, 23) */,
  32'h3d45eb5b /* (7, 26, 23) */,
  32'h3d215063 /* (3, 26, 23) */,
  32'h3d52081f /* (31, 22, 23) */,
  32'h3d781ae6 /* (27, 22, 23) */,
  32'h3dbbc730 /* (23, 22, 23) */,
  32'h3e1d56b2 /* (19, 22, 23) */,
  32'h3e2b3653 /* (15, 22, 23) */,
  32'h3df71c69 /* (11, 22, 23) */,
  32'h3d94014f /* (7, 22, 23) */,
  32'h3d5dae2c /* (3, 22, 23) */,
  32'h3d90dff9 /* (31, 18, 23) */,
  32'h3db24f8e /* (27, 18, 23) */,
  32'h3e10cac5 /* (23, 18, 23) */,
  32'h3e821787 /* (19, 18, 23) */,
  32'h3e91e4f8 /* (15, 18, 23) */,
  32'h3e458f30 /* (11, 18, 23) */,
  32'h3ddc09d8 /* (7, 18, 23) */,
  32'h3d9b2a7b /* (3, 18, 23) */,
  32'h3d90dff9 /* (31, 14, 23) */,
  32'h3db24f8e /* (27, 14, 23) */,
  32'h3e10cac5 /* (23, 14, 23) */,
  32'h3e821787 /* (19, 14, 23) */,
  32'h3e91e4f8 /* (15, 14, 23) */,
  32'h3e458f30 /* (11, 14, 23) */,
  32'h3ddc09d8 /* (7, 14, 23) */,
  32'h3d9b2a7b /* (3, 14, 23) */,
  32'h3d52081f /* (31, 10, 23) */,
  32'h3d781ae6 /* (27, 10, 23) */,
  32'h3dbbc730 /* (23, 10, 23) */,
  32'h3e1d56b2 /* (19, 10, 23) */,
  32'h3e2b3653 /* (15, 10, 23) */,
  32'h3df71c69 /* (11, 10, 23) */,
  32'h3d94014f /* (7, 10, 23) */,
  32'h3d5dae2c /* (3, 10, 23) */,
  32'h3d1c53e8 /* (31, 6, 23) */,
  32'h3d2db0cc /* (27, 6, 23) */,
  32'h3d6fd024 /* (23, 6, 23) */,
  32'h3db9d5f4 /* (19, 6, 23) */,
  32'h3dc42ad0 /* (15, 6, 23) */,
  32'h3d9750ce /* (11, 6, 23) */,
  32'h3d45eb5b /* (7, 6, 23) */,
  32'h3d215063 /* (3, 6, 23) */,
  32'h3d11c69f /* (31, 2, 23) */,
  32'h3d18622e /* (27, 2, 23) */,
  32'h3d42665b /* (23, 2, 23) */,
  32'h3d8e358b /* (19, 2, 23) */,
  32'h3d9314c2 /* (15, 2, 23) */,
  32'h3d6d9fa3 /* (11, 2, 23) */,
  32'h3d26a1b5 /* (7, 2, 23) */,
  32'h3d12f42a /* (3, 2, 23) */,
  32'h3d214ba3 /* (31, 30, 19) */,
  32'h3d3d84de /* (27, 30, 19) */,
  32'h3d8e358b /* (23, 30, 19) */,
  32'h3dec70da /* (19, 30, 19) */,
  32'h3e003b1e /* (15, 30, 19) */,
  32'h3dba5db4 /* (11, 30, 19) */,
  32'h3d6129ae /* (7, 30, 19) */,
  32'h3d29e985 /* (3, 30, 19) */,
  32'h3d4876ff /* (31, 26, 19) */,
  32'h3d700ffa /* (27, 26, 19) */,
  32'h3db9d5f4 /* (23, 26, 19) */,
  32'h3e1f113d /* (19, 26, 19) */,
  32'h3e2ea39a /* (15, 26, 19) */,
  32'h3df74dbc /* (11, 26, 19) */,
  32'h3d90c8a7 /* (7, 26, 19) */,
  32'h3d54a03b /* (3, 26, 19) */,
  32'h3d9e7894 /* (31, 22, 19) */,
  32'h3dc29629 /* (27, 22, 19) */,
  32'h3e1d56b2 /* (23, 22, 19) */,
  32'h3e8cbae1 /* (19, 22, 19) */,
  32'h3e9d80fb /* (15, 22, 19) */,
  32'h3e562fb1 /* (11, 22, 19) */,
  32'h3defa49b /* (7, 22, 19) */,
  32'h3da99659 /* (3, 22, 19) */,
  32'h3df65860 /* (31, 18, 19) */,
  32'h3e1a8d8c /* (27, 18, 19) */,
  32'h3e821787 /* (23, 18, 19) */,
  32'h3ef33ce4 /* (19, 18, 19) */,
  32'h3f0af24f /* (15, 18, 19) */,
  32'h3eb517ce /* (11, 18, 19) */,
  32'h3e41f14c /* (7, 18, 19) */,
  32'h3e04d0b8 /* (3, 18, 19) */,
  32'h3df65860 /* (31, 14, 19) */,
  32'h3e1a8d8c /* (27, 14, 19) */,
  32'h3e821787 /* (23, 14, 19) */,
  32'h3ef33ce4 /* (19, 14, 19) */,
  32'h3f0af24f /* (15, 14, 19) */,
  32'h3eb517ce /* (11, 14, 19) */,
  32'h3e41f14c /* (7, 14, 19) */,
  32'h3e04d0b8 /* (3, 14, 19) */,
  32'h3d9e7894 /* (31, 10, 19) */,
  32'h3dc29629 /* (27, 10, 19) */,
  32'h3e1d56b2 /* (23, 10, 19) */,
  32'h3e8cbae1 /* (19, 10, 19) */,
  32'h3e9d80fb /* (15, 10, 19) */,
  32'h3e562fb1 /* (11, 10, 19) */,
  32'h3defa49b /* (7, 10, 19) */,
  32'h3da99659 /* (3, 10, 19) */,
  32'h3d4876ff /* (31, 6, 19) */,
  32'h3d700ffa /* (27, 6, 19) */,
  32'h3db9d5f4 /* (23, 6, 19) */,
  32'h3e1f113d /* (19, 6, 19) */,
  32'h3e2ea39a /* (15, 6, 19) */,
  32'h3df74dbc /* (11, 6, 19) */,
  32'h3d90c8a7 /* (7, 6, 19) */,
  32'h3d54a03b /* (3, 6, 19) */,
  32'h3d214ba3 /* (31, 2, 19) */,
  32'h3d3d84de /* (27, 2, 19) */,
  32'h3d8e358b /* (23, 2, 19) */,
  32'h3dec70da /* (19, 2, 19) */,
  32'h3e003b1e /* (15, 2, 19) */,
  32'h3dba5db4 /* (11, 2, 19) */,
  32'h3d6129ae /* (7, 2, 19) */,
  32'h3d29e985 /* (3, 2, 19) */,
  32'h3d1a0745 /* (31, 30, 15) */,
  32'h3d3a7be5 /* (27, 30, 15) */,
  32'h3d9314c2 /* (23, 30, 15) */,
  32'h3e003b1e /* (19, 30, 15) */,
  32'h3e0de5f8 /* (15, 30, 15) */,
  32'h3dc59b81 /* (11, 30, 15) */,
  32'h3d62f778 /* (7, 30, 15) */,
  32'h3d240321 /* (3, 30, 15) */,
  32'h3d46f53f /* (31, 26, 15) */,
  32'h3d73b16f /* (27, 26, 15) */,
  32'h3dc42ad0 /* (23, 26, 15) */,
  32'h3e2ea39a /* (19, 26, 15) */,
  32'h3e430b11 /* (15, 26, 15) */,
  32'h3e0533d0 /* (11, 26, 15) */,
  32'h3d95be73 /* (7, 26, 15) */,
  32'h3d54ba37 /* (3, 26, 15) */,
  32'h3da5ac70 /* (31, 22, 15) */,
  32'h3dce52e6 /* (27, 22, 15) */,
  32'h3e2b3653 /* (23, 22, 15) */,
  32'h3e9d80fb /* (19, 22, 15) */,
  32'h3eb2925b /* (15, 22, 15) */,
  32'h3e6c6ac0 /* (11, 22, 15) */,
  32'h3e009a19 /* (7, 22, 15) */,
  32'h3db22d06 /* (3, 22, 15) */,
  32'h3e06d8bb /* (31, 18, 15) */,
  32'h3e2a981c /* (27, 18, 15) */,
  32'h3e91e4f8 /* (23, 18, 15) */,
  32'h3f0af24f /* (19, 18, 15) */,
  32'h3f202f9a /* (15, 18, 15) */,
  32'h3eccf8ff /* (11, 18, 15) */,
  32'h3e57a44b /* (7, 18, 15) */,
  32'h3e11d12f /* (3, 18, 15) */,
  32'h3e06d8bb /* (31, 14, 15) */,
  32'h3e2a981c /* (27, 14, 15) */,
  32'h3e91e4f8 /* (23, 14, 15) */,
  32'h3f0af24f /* (19, 14, 15) */,
  32'h3f202f9a /* (15, 14, 15) */,
  32'h3eccf8ff /* (11, 14, 15) */,
  32'h3e57a44b /* (7, 14, 15) */,
  32'h3e11d12f /* (3, 14, 15) */,
  32'h3da5ac70 /* (31, 10, 15) */,
  32'h3dce52e6 /* (27, 10, 15) */,
  32'h3e2b3653 /* (23, 10, 15) */,
  32'h3e9d80fb /* (19, 10, 15) */,
  32'h3eb2925b /* (15, 10, 15) */,
  32'h3e6c6ac0 /* (11, 10, 15) */,
  32'h3e009a19 /* (7, 10, 15) */,
  32'h3db22d06 /* (3, 10, 15) */,
  32'h3d46f53f /* (31, 6, 15) */,
  32'h3d73b16f /* (27, 6, 15) */,
  32'h3dc42ad0 /* (23, 6, 15) */,
  32'h3e2ea39a /* (19, 6, 15) */,
  32'h3e430b11 /* (15, 6, 15) */,
  32'h3e0533d0 /* (11, 6, 15) */,
  32'h3d95be73 /* (7, 6, 15) */,
  32'h3d54ba37 /* (3, 6, 15) */,
  32'h3d1a0745 /* (31, 2, 15) */,
  32'h3d3a7be5 /* (27, 2, 15) */,
  32'h3d9314c2 /* (23, 2, 15) */,
  32'h3e003b1e /* (19, 2, 15) */,
  32'h3e0de5f8 /* (15, 2, 15) */,
  32'h3dc59b81 /* (11, 2, 15) */,
  32'h3d62f778 /* (7, 2, 15) */,
  32'h3d240321 /* (3, 2, 15) */,
  32'h3d16ed42 /* (31, 30, 11) */,
  32'h3d29823f /* (27, 30, 11) */,
  32'h3d6d9fa3 /* (23, 30, 11) */,
  32'h3dba5db4 /* (19, 30, 11) */,
  32'h3dc59b81 /* (15, 30, 11) */,
  32'h3d96eb50 /* (11, 30, 11) */,
  32'h3d42a7b8 /* (7, 30, 11) */,
  32'h3d1c5f03 /* (3, 30, 11) */,
  32'h3d31191b /* (31, 26, 11) */,
  32'h3d4d9045 /* (27, 26, 11) */,
  32'h3d9750ce /* (23, 26, 11) */,
  32'h3df74dbc /* (19, 26, 11) */,
  32'h3e0533d0 /* (15, 26, 11) */,
  32'h3dc480ba /* (11, 26, 11) */,
  32'h3d71ecf9 /* (7, 26, 11) */,
  32'h3d39bb76 /* (3, 26, 11) */,
  32'h3d829849 /* (31, 22, 11) */,
  32'h3d9d9380 /* (27, 22, 11) */,
  32'h3df71c69 /* (23, 22, 11) */,
  32'h3e562fb1 /* (19, 22, 11) */,
  32'h3e6c6ac0 /* (15, 22, 11) */,
  32'h3e257fc6 /* (11, 22, 11) */,
  32'h3dbf3f1d /* (7, 22, 11) */,
  32'h3d8ae43c /* (3, 22, 11) */,
  32'h3dc01db4 /* (31, 18, 11) */,
  32'h3deed79f /* (27, 18, 11) */,
  32'h3e458f30 /* (23, 18, 11) */,
  32'h3eb517ce /* (19, 18, 11) */,
  32'h3eccf8ff /* (15, 18, 11) */,
  32'h3e882756 /* (11, 18, 11) */,
  32'h3e14a5c9 /* (7, 18, 11) */,
  32'h3dce7d45 /* (3, 18, 11) */,
  32'h3dc01db4 /* (31, 14, 11) */,
  32'h3deed79f /* (27, 14, 11) */,
  32'h3e458f30 /* (23, 14, 11) */,
  32'h3eb517ce /* (19, 14, 11) */,
  32'h3eccf8ff /* (15, 14, 11) */,
  32'h3e882756 /* (11, 14, 11) */,
  32'h3e14a5c9 /* (7, 14, 11) */,
  32'h3dce7d45 /* (3, 14, 11) */,
  32'h3d829849 /* (31, 10, 11) */,
  32'h3d9d9380 /* (27, 10, 11) */,
  32'h3df71c69 /* (23, 10, 11) */,
  32'h3e562fb1 /* (19, 10, 11) */,
  32'h3e6c6ac0 /* (15, 10, 11) */,
  32'h3e257fc6 /* (11, 10, 11) */,
  32'h3dbf3f1d /* (7, 10, 11) */,
  32'h3d8ae43c /* (3, 10, 11) */,
  32'h3d31191b /* (31, 6, 11) */,
  32'h3d4d9045 /* (27, 6, 11) */,
  32'h3d9750ce /* (23, 6, 11) */,
  32'h3df74dbc /* (19, 6, 11) */,
  32'h3e0533d0 /* (15, 6, 11) */,
  32'h3dc480ba /* (11, 6, 11) */,
  32'h3d71ecf9 /* (7, 6, 11) */,
  32'h3d39bb76 /* (3, 6, 11) */,
  32'h3d16ed42 /* (31, 2, 11) */,
  32'h3d29823f /* (27, 2, 11) */,
  32'h3d6d9fa3 /* (23, 2, 11) */,
  32'h3dba5db4 /* (19, 2, 11) */,
  32'h3dc59b81 /* (15, 2, 11) */,
  32'h3d96eb50 /* (11, 2, 11) */,
  32'h3d42a7b8 /* (7, 2, 11) */,
  32'h3d1c5f03 /* (3, 2, 11) */,
  32'h3d20a35e /* (31, 30, 7) */,
  32'h3d14b1c0 /* (27, 30, 7) */,
  32'h3d26a1b5 /* (23, 30, 7) */,
  32'h3d6129ae /* (19, 30, 7) */,
  32'h3d62f778 /* (15, 30, 7) */,
  32'h3d42a7b8 /* (11, 30, 7) */,
  32'h3d1777c7 /* (7, 30, 7) */,
  32'h3d1a2949 /* (3, 30, 7) */,
  32'h3d146a43 /* (31, 26, 7) */,
  32'h3d1b2471 /* (27, 26, 7) */,
  32'h3d45eb5b /* (23, 26, 7) */,
  32'h3d90c8a7 /* (19, 26, 7) */,
  32'h3d95be73 /* (15, 26, 7) */,
  32'h3d71ecf9 /* (11, 26, 7) */,
  32'h3d29a602 /* (7, 26, 7) */,
  32'h3d159d44 /* (3, 26, 7) */,
  32'h3d305430 /* (31, 22, 7) */,
  32'h3d4b3dc7 /* (27, 22, 7) */,
  32'h3d94014f /* (23, 22, 7) */,
  32'h3defa49b /* (19, 22, 7) */,
  32'h3e009a19 /* (15, 22, 7) */,
  32'h3dbf3f1d /* (11, 22, 7) */,
  32'h3d6deb12 /* (7, 22, 7) */,
  32'h3d387393 /* (3, 22, 7) */,
  32'h3d62906c /* (31, 18, 7) */,
  32'h3d8a0000 /* (27, 18, 7) */,
  32'h3ddc09d8 /* (23, 18, 7) */,
  32'h3e41f14c /* (19, 18, 7) */,
  32'h3e57a44b /* (15, 18, 7) */,
  32'h3e14a5c9 /* (11, 18, 7) */,
  32'h3da8d240 /* (7, 18, 7) */,
  32'h3d71c736 /* (3, 18, 7) */,
  32'h3d62906c /* (31, 14, 7) */,
  32'h3d8a0000 /* (27, 14, 7) */,
  32'h3ddc09d8 /* (23, 14, 7) */,
  32'h3e41f14c /* (19, 14, 7) */,
  32'h3e57a44b /* (15, 14, 7) */,
  32'h3e14a5c9 /* (11, 14, 7) */,
  32'h3da8d240 /* (7, 14, 7) */,
  32'h3d71c736 /* (3, 14, 7) */,
  32'h3d305430 /* (31, 10, 7) */,
  32'h3d4b3dc7 /* (27, 10, 7) */,
  32'h3d94014f /* (23, 10, 7) */,
  32'h3defa49b /* (19, 10, 7) */,
  32'h3e009a19 /* (15, 10, 7) */,
  32'h3dbf3f1d /* (11, 10, 7) */,
  32'h3d6deb12 /* (7, 10, 7) */,
  32'h3d387393 /* (3, 10, 7) */,
  32'h3d146a43 /* (31, 6, 7) */,
  32'h3d1b2471 /* (27, 6, 7) */,
  32'h3d45eb5b /* (23, 6, 7) */,
  32'h3d90c8a7 /* (19, 6, 7) */,
  32'h3d95be73 /* (15, 6, 7) */,
  32'h3d71ecf9 /* (11, 6, 7) */,
  32'h3d29a602 /* (7, 6, 7) */,
  32'h3d159d44 /* (3, 6, 7) */,
  32'h3d20a35e /* (31, 2, 7) */,
  32'h3d14b1c0 /* (27, 2, 7) */,
  32'h3d26a1b5 /* (23, 2, 7) */,
  32'h3d6129ae /* (19, 2, 7) */,
  32'h3d62f778 /* (15, 2, 7) */,
  32'h3d42a7b8 /* (11, 2, 7) */,
  32'h3d1777c7 /* (7, 2, 7) */,
  32'h3d1a2949 /* (3, 2, 7) */,
  32'h3dbfa8df /* (31, 30, 3) */,
  32'h3d3cd255 /* (27, 30, 3) */,
  32'h3d12f42a /* (23, 30, 3) */,
  32'h3d29e985 /* (19, 30, 3) */,
  32'h3d240321 /* (15, 30, 3) */,
  32'h3d1c5f03 /* (11, 30, 3) */,
  32'h3d1a2949 /* (7, 30, 3) */,
  32'h3d866355 /* (3, 30, 3) */,
  32'h3d2ba889 /* (31, 26, 3) */,
  32'h3d16d305 /* (27, 26, 3) */,
  32'h3d215063 /* (23, 26, 3) */,
  32'h3d54a03b /* (19, 26, 3) */,
  32'h3d54ba37 /* (15, 26, 3) */,
  32'h3d39bb76 /* (11, 26, 3) */,
  32'h3d159d44 /* (7, 26, 3) */,
  32'h3d211f1b /* (3, 26, 3) */,
  32'h3d14c0fd /* (31, 22, 3) */,
  32'h3d2344c4 /* (27, 22, 3) */,
  32'h3d5dae2c /* (23, 22, 3) */,
  32'h3da99659 /* (19, 22, 3) */,
  32'h3db22d06 /* (15, 22, 3) */,
  32'h3d8ae43c /* (11, 22, 3) */,
  32'h3d387393 /* (7, 22, 3) */,
  32'h3d18cb02 /* (3, 22, 3) */,
  32'h3d276174 /* (31, 18, 3) */,
  32'h3d487174 /* (27, 18, 3) */,
  32'h3d9b2a7b /* (23, 18, 3) */,
  32'h3e04d0b8 /* (19, 18, 3) */,
  32'h3e11d12f /* (15, 18, 3) */,
  32'h3dce7d45 /* (11, 18, 3) */,
  32'h3d71c736 /* (7, 18, 3) */,
  32'h3d3188e3 /* (3, 18, 3) */,
  32'h3d276174 /* (31, 14, 3) */,
  32'h3d487174 /* (27, 14, 3) */,
  32'h3d9b2a7b /* (23, 14, 3) */,
  32'h3e04d0b8 /* (19, 14, 3) */,
  32'h3e11d12f /* (15, 14, 3) */,
  32'h3dce7d45 /* (11, 14, 3) */,
  32'h3d71c736 /* (7, 14, 3) */,
  32'h3d3188e3 /* (3, 14, 3) */,
  32'h3d14c0fd /* (31, 10, 3) */,
  32'h3d2344c4 /* (27, 10, 3) */,
  32'h3d5dae2c /* (23, 10, 3) */,
  32'h3da99659 /* (19, 10, 3) */,
  32'h3db22d06 /* (15, 10, 3) */,
  32'h3d8ae43c /* (11, 10, 3) */,
  32'h3d387393 /* (7, 10, 3) */,
  32'h3d18cb02 /* (3, 10, 3) */,
  32'h3d2ba889 /* (31, 6, 3) */,
  32'h3d16d305 /* (27, 6, 3) */,
  32'h3d215063 /* (23, 6, 3) */,
  32'h3d54a03b /* (19, 6, 3) */,
  32'h3d54ba37 /* (15, 6, 3) */,
  32'h3d39bb76 /* (11, 6, 3) */,
  32'h3d159d44 /* (7, 6, 3) */,
  32'h3d211f1b /* (3, 6, 3) */,
  32'h3dbfa8df /* (31, 2, 3) */,
  32'h3d3cd255 /* (27, 2, 3) */,
  32'h3d12f42a /* (23, 2, 3) */,
  32'h3d29e985 /* (19, 2, 3) */,
  32'h3d240321 /* (15, 2, 3) */,
  32'h3d1c5f03 /* (11, 2, 3) */,
  32'h3d1a2949 /* (7, 2, 3) */,
  32'h3d866355 /* (3, 2, 3) */,
  32'h3e0c4d23 /* (30, 30, 31) */,
  32'h3d3543e4 /* (26, 30, 31) */,
  32'h3d12ac07 /* (22, 30, 31) */,
  32'h3d217487 /* (18, 30, 31) */,
  32'h3d217487 /* (14, 30, 31) */,
  32'h3d12ac07 /* (10, 30, 31) */,
  32'h3d3543e4 /* (6, 30, 31) */,
  32'h3e0c4d23 /* (2, 30, 31) */,
  32'h3d3543e4 /* (30, 26, 31) */,
  32'h3d15cc97 /* (26, 26, 31) */,
  32'h3d2567ce /* (22, 26, 31) */,
  32'h3d4cf093 /* (18, 26, 31) */,
  32'h3d4cf093 /* (14, 26, 31) */,
  32'h3d2567ce /* (10, 26, 31) */,
  32'h3d15cc97 /* (6, 26, 31) */,
  32'h3d3543e4 /* (2, 26, 31) */,
  32'h3d12ac07 /* (30, 22, 31) */,
  32'h3d2567ce /* (26, 22, 31) */,
  32'h3d699f13 /* (22, 22, 31) */,
  32'h3da6958f /* (18, 22, 31) */,
  32'h3da6958f /* (14, 22, 31) */,
  32'h3d699f13 /* (10, 22, 31) */,
  32'h3d2567ce /* (6, 22, 31) */,
  32'h3d12ac07 /* (2, 22, 31) */,
  32'h3d217487 /* (30, 18, 31) */,
  32'h3d4cf093 /* (26, 18, 31) */,
  32'h3da6958f /* (22, 18, 31) */,
  32'h3e04a438 /* (18, 18, 31) */,
  32'h3e04a438 /* (14, 18, 31) */,
  32'h3da6958f /* (10, 18, 31) */,
  32'h3d4cf093 /* (6, 18, 31) */,
  32'h3d217487 /* (2, 18, 31) */,
  32'h3d217487 /* (30, 14, 31) */,
  32'h3d4cf093 /* (26, 14, 31) */,
  32'h3da6958f /* (22, 14, 31) */,
  32'h3e04a438 /* (18, 14, 31) */,
  32'h3e04a438 /* (14, 14, 31) */,
  32'h3da6958f /* (10, 14, 31) */,
  32'h3d4cf093 /* (6, 14, 31) */,
  32'h3d217487 /* (2, 14, 31) */,
  32'h3d12ac07 /* (30, 10, 31) */,
  32'h3d2567ce /* (26, 10, 31) */,
  32'h3d699f13 /* (22, 10, 31) */,
  32'h3da6958f /* (18, 10, 31) */,
  32'h3da6958f /* (14, 10, 31) */,
  32'h3d699f13 /* (10, 10, 31) */,
  32'h3d2567ce /* (6, 10, 31) */,
  32'h3d12ac07 /* (2, 10, 31) */,
  32'h3d3543e4 /* (30, 6, 31) */,
  32'h3d15cc97 /* (26, 6, 31) */,
  32'h3d2567ce /* (22, 6, 31) */,
  32'h3d4cf093 /* (18, 6, 31) */,
  32'h3d4cf093 /* (14, 6, 31) */,
  32'h3d2567ce /* (10, 6, 31) */,
  32'h3d15cc97 /* (6, 6, 31) */,
  32'h3d3543e4 /* (2, 6, 31) */,
  32'h3e0c4d23 /* (30, 2, 31) */,
  32'h3d3543e4 /* (26, 2, 31) */,
  32'h3d12ac07 /* (22, 2, 31) */,
  32'h3d217487 /* (18, 2, 31) */,
  32'h3d217487 /* (14, 2, 31) */,
  32'h3d12ac07 /* (10, 2, 31) */,
  32'h3d3543e4 /* (6, 2, 31) */,
  32'h3e0c4d23 /* (2, 2, 31) */,
  32'h3d4ca49b /* (30, 30, 27) */,
  32'h3d18df8d /* (26, 30, 27) */,
  32'h3d1f9f49 /* (22, 30, 27) */,
  32'h3d40d8bf /* (18, 30, 27) */,
  32'h3d40d8bf /* (14, 30, 27) */,
  32'h3d1f9f49 /* (10, 30, 27) */,
  32'h3d18df8d /* (6, 30, 27) */,
  32'h3d4ca49b /* (2, 30, 27) */,
  32'h3d18df8d /* (30, 26, 27) */,
  32'h3d16bb8b /* (26, 26, 27) */,
  32'h3d3c300c /* (22, 26, 27) */,
  32'h3d786cd6 /* (18, 26, 27) */,
  32'h3d786cd6 /* (14, 26, 27) */,
  32'h3d3c300c /* (10, 26, 27) */,
  32'h3d16bb8b /* (6, 26, 27) */,
  32'h3d18df8d /* (2, 26, 27) */,
  32'h3d1f9f49 /* (30, 22, 27) */,
  32'h3d3c300c /* (26, 22, 27) */,
  32'h3d8b85a2 /* (22, 22, 27) */,
  32'h3dce13fe /* (18, 22, 27) */,
  32'h3dce13fe /* (14, 22, 27) */,
  32'h3d8b85a2 /* (10, 22, 27) */,
  32'h3d3c300c /* (6, 22, 27) */,
  32'h3d1f9f49 /* (2, 22, 27) */,
  32'h3d40d8bf /* (30, 18, 27) */,
  32'h3d786cd6 /* (26, 18, 27) */,
  32'h3dce13fe /* (22, 18, 27) */,
  32'h3e27240a /* (18, 18, 27) */,
  32'h3e27240a /* (14, 18, 27) */,
  32'h3dce13fe /* (10, 18, 27) */,
  32'h3d786cd6 /* (6, 18, 27) */,
  32'h3d40d8bf /* (2, 18, 27) */,
  32'h3d40d8bf /* (30, 14, 27) */,
  32'h3d786cd6 /* (26, 14, 27) */,
  32'h3dce13fe /* (22, 14, 27) */,
  32'h3e27240a /* (18, 14, 27) */,
  32'h3e27240a /* (14, 14, 27) */,
  32'h3dce13fe /* (10, 14, 27) */,
  32'h3d786cd6 /* (6, 14, 27) */,
  32'h3d40d8bf /* (2, 14, 27) */,
  32'h3d1f9f49 /* (30, 10, 27) */,
  32'h3d3c300c /* (26, 10, 27) */,
  32'h3d8b85a2 /* (22, 10, 27) */,
  32'h3dce13fe /* (18, 10, 27) */,
  32'h3dce13fe /* (14, 10, 27) */,
  32'h3d8b85a2 /* (10, 10, 27) */,
  32'h3d3c300c /* (6, 10, 27) */,
  32'h3d1f9f49 /* (2, 10, 27) */,
  32'h3d18df8d /* (30, 6, 27) */,
  32'h3d16bb8b /* (26, 6, 27) */,
  32'h3d3c300c /* (22, 6, 27) */,
  32'h3d786cd6 /* (18, 6, 27) */,
  32'h3d786cd6 /* (14, 6, 27) */,
  32'h3d3c300c /* (10, 6, 27) */,
  32'h3d16bb8b /* (6, 6, 27) */,
  32'h3d18df8d /* (2, 6, 27) */,
  32'h3d4ca49b /* (30, 2, 27) */,
  32'h3d18df8d /* (26, 2, 27) */,
  32'h3d1f9f49 /* (22, 2, 27) */,
  32'h3d40d8bf /* (18, 2, 27) */,
  32'h3d40d8bf /* (14, 2, 27) */,
  32'h3d1f9f49 /* (10, 2, 27) */,
  32'h3d18df8d /* (6, 2, 27) */,
  32'h3d4ca49b /* (2, 2, 27) */,
  32'h3d1214c5 /* (30, 30, 23) */,
  32'h3d1e19af /* (26, 30, 23) */,
  32'h3d56480e /* (22, 30, 23) */,
  32'h3d94a37c /* (18, 30, 23) */,
  32'h3d94a37c /* (14, 30, 23) */,
  32'h3d56480e /* (10, 30, 23) */,
  32'h3d1e19af /* (6, 30, 23) */,
  32'h3d1214c5 /* (2, 30, 23) */,
  32'h3d1e19af /* (30, 26, 23) */,
  32'h3d37f9d0 /* (26, 26, 23) */,
  32'h3d866682 /* (22, 26, 23) */,
  32'h3dc45939 /* (18, 26, 23) */,
  32'h3dc45939 /* (14, 26, 23) */,
  32'h3d866682 /* (10, 26, 23) */,
  32'h3d37f9d0 /* (6, 26, 23) */,
  32'h3d1e19af /* (2, 26, 23) */,
  32'h3d56480e /* (30, 22, 23) */,
  32'h3d866682 /* (26, 22, 23) */,
  32'h3dd7137d /* (22, 22, 23) */,
  32'h3e28e750 /* (18, 22, 23) */,
  32'h3e28e750 /* (14, 22, 23) */,
  32'h3dd7137d /* (10, 22, 23) */,
  32'h3d866682 /* (6, 22, 23) */,
  32'h3d56480e /* (2, 22, 23) */,
  32'h3d94a37c /* (30, 18, 23) */,
  32'h3dc45939 /* (26, 18, 23) */,
  32'h3e28e750 /* (22, 18, 23) */,
  32'h3e8dd733 /* (18, 18, 23) */,
  32'h3e8dd733 /* (14, 18, 23) */,
  32'h3e28e750 /* (10, 18, 23) */,
  32'h3dc45939 /* (6, 18, 23) */,
  32'h3d94a37c /* (2, 18, 23) */,
  32'h3d94a37c /* (30, 14, 23) */,
  32'h3dc45939 /* (26, 14, 23) */,
  32'h3e28e750 /* (22, 14, 23) */,
  32'h3e8dd733 /* (18, 14, 23) */,
  32'h3e8dd733 /* (14, 14, 23) */,
  32'h3e28e750 /* (10, 14, 23) */,
  32'h3dc45939 /* (6, 14, 23) */,
  32'h3d94a37c /* (2, 14, 23) */,
  32'h3d56480e /* (30, 10, 23) */,
  32'h3d866682 /* (26, 10, 23) */,
  32'h3dd7137d /* (22, 10, 23) */,
  32'h3e28e750 /* (18, 10, 23) */,
  32'h3e28e750 /* (14, 10, 23) */,
  32'h3dd7137d /* (10, 10, 23) */,
  32'h3d866682 /* (6, 10, 23) */,
  32'h3d56480e /* (2, 10, 23) */,
  32'h3d1e19af /* (30, 6, 23) */,
  32'h3d37f9d0 /* (26, 6, 23) */,
  32'h3d866682 /* (22, 6, 23) */,
  32'h3dc45939 /* (18, 6, 23) */,
  32'h3dc45939 /* (14, 6, 23) */,
  32'h3d866682 /* (10, 6, 23) */,
  32'h3d37f9d0 /* (6, 6, 23) */,
  32'h3d1e19af /* (2, 6, 23) */,
  32'h3d1214c5 /* (30, 2, 23) */,
  32'h3d1e19af /* (26, 2, 23) */,
  32'h3d56480e /* (22, 2, 23) */,
  32'h3d94a37c /* (18, 2, 23) */,
  32'h3d94a37c /* (14, 2, 23) */,
  32'h3d56480e /* (10, 2, 23) */,
  32'h3d1e19af /* (6, 2, 23) */,
  32'h3d1214c5 /* (2, 2, 23) */,
  32'h3d246fbd /* (30, 30, 19) */,
  32'h3d4ce87b /* (26, 30, 19) */,
  32'h3da2895a /* (22, 30, 19) */,
  32'h3dfd653f /* (18, 30, 19) */,
  32'h3dfd653f /* (14, 30, 19) */,
  32'h3da2895a /* (10, 30, 19) */,
  32'h3d4ce87b /* (6, 30, 19) */,
  32'h3d246fbd /* (2, 30, 19) */,
  32'h3d4ce87b /* (30, 26, 19) */,
  32'h3d82bc35 /* (26, 26, 19) */,
  32'h3dd610ea /* (22, 26, 19) */,
  32'h3e2b8c37 /* (18, 26, 19) */,
  32'h3e2b8c37 /* (14, 26, 19) */,
  32'h3dd610ea /* (10, 26, 19) */,
  32'h3d82bc35 /* (6, 26, 19) */,
  32'h3d4ce87b /* (2, 26, 19) */,
  32'h3da2895a /* (30, 22, 19) */,
  32'h3dd610ea /* (26, 22, 19) */,
  32'h3e37540b /* (22, 22, 19) */,
  32'h3e994798 /* (18, 22, 19) */,
  32'h3e994798 /* (14, 22, 19) */,
  32'h3e37540b /* (10, 22, 19) */,
  32'h3dd610ea /* (6, 22, 19) */,
  32'h3da2895a /* (2, 22, 19) */,
  32'h3dfd653f /* (30, 18, 19) */,
  32'h3e2b8c37 /* (26, 18, 19) */,
  32'h3e994798 /* (22, 18, 19) */,
  32'h3f05dc96 /* (18, 18, 19) */,
  32'h3f05dc96 /* (14, 18, 19) */,
  32'h3e994798 /* (10, 18, 19) */,
  32'h3e2b8c37 /* (6, 18, 19) */,
  32'h3dfd653f /* (2, 18, 19) */,
  32'h3dfd653f /* (30, 14, 19) */,
  32'h3e2b8c37 /* (26, 14, 19) */,
  32'h3e994798 /* (22, 14, 19) */,
  32'h3f05dc96 /* (18, 14, 19) */,
  32'h3f05dc96 /* (14, 14, 19) */,
  32'h3e994798 /* (10, 14, 19) */,
  32'h3e2b8c37 /* (6, 14, 19) */,
  32'h3dfd653f /* (2, 14, 19) */,
  32'h3da2895a /* (30, 10, 19) */,
  32'h3dd610ea /* (26, 10, 19) */,
  32'h3e37540b /* (22, 10, 19) */,
  32'h3e994798 /* (18, 10, 19) */,
  32'h3e994798 /* (14, 10, 19) */,
  32'h3e37540b /* (10, 10, 19) */,
  32'h3dd610ea /* (6, 10, 19) */,
  32'h3da2895a /* (2, 10, 19) */,
  32'h3d4ce87b /* (30, 6, 19) */,
  32'h3d82bc35 /* (26, 6, 19) */,
  32'h3dd610ea /* (22, 6, 19) */,
  32'h3e2b8c37 /* (18, 6, 19) */,
  32'h3e2b8c37 /* (14, 6, 19) */,
  32'h3dd610ea /* (10, 6, 19) */,
  32'h3d82bc35 /* (6, 6, 19) */,
  32'h3d4ce87b /* (2, 6, 19) */,
  32'h3d246fbd /* (30, 2, 19) */,
  32'h3d4ce87b /* (26, 2, 19) */,
  32'h3da2895a /* (22, 2, 19) */,
  32'h3dfd653f /* (18, 2, 19) */,
  32'h3dfd653f /* (14, 2, 19) */,
  32'h3da2895a /* (10, 2, 19) */,
  32'h3d4ce87b /* (6, 2, 19) */,
  32'h3d246fbd /* (2, 2, 19) */,
  32'h3d1dadb9 /* (30, 30, 15) */,
  32'h3d4bfe66 /* (26, 30, 15) */,
  32'h3daa3ec9 /* (22, 30, 15) */,
  32'h3e0adb0d /* (18, 30, 15) */,
  32'h3e0adb0d /* (14, 30, 15) */,
  32'h3daa3ec9 /* (10, 30, 15) */,
  32'h3d4bfe66 /* (6, 30, 15) */,
  32'h3d1dadb9 /* (2, 30, 15) */,
  32'h3d4bfe66 /* (30, 26, 15) */,
  32'h3d85e8bf /* (26, 26, 15) */,
  32'h3de44bb3 /* (22, 26, 15) */,
  32'h3e3e01e0 /* (18, 26, 15) */,
  32'h3e3e01e0 /* (14, 26, 15) */,
  32'h3de44bb3 /* (10, 26, 15) */,
  32'h3d85e8bf /* (6, 26, 15) */,
  32'h3d4bfe66 /* (2, 26, 15) */,
  32'h3daa3ec9 /* (30, 22, 15) */,
  32'h3de44bb3 /* (26, 22, 15) */,
  32'h3e48eba4 /* (22, 22, 15) */,
  32'h3eacaf9b /* (18, 22, 15) */,
  32'h3eacaf9b /* (14, 22, 15) */,
  32'h3e48eba4 /* (10, 22, 15) */,
  32'h3de44bb3 /* (6, 22, 15) */,
  32'h3daa3ec9 /* (2, 22, 15) */,
  32'h3e0adb0d /* (30, 18, 15) */,
  32'h3e3e01e0 /* (26, 18, 15) */,
  32'h3eacaf9b /* (22, 18, 15) */,
  32'h3f19a2a7 /* (18, 18, 15) */,
  32'h3f19a2a7 /* (14, 18, 15) */,
  32'h3eacaf9b /* (10, 18, 15) */,
  32'h3e3e01e0 /* (6, 18, 15) */,
  32'h3e0adb0d /* (2, 18, 15) */,
  32'h3e0adb0d /* (30, 14, 15) */,
  32'h3e3e01e0 /* (26, 14, 15) */,
  32'h3eacaf9b /* (22, 14, 15) */,
  32'h3f19a2a7 /* (18, 14, 15) */,
  32'h3f19a2a7 /* (14, 14, 15) */,
  32'h3eacaf9b /* (10, 14, 15) */,
  32'h3e3e01e0 /* (6, 14, 15) */,
  32'h3e0adb0d /* (2, 14, 15) */,
  32'h3daa3ec9 /* (30, 10, 15) */,
  32'h3de44bb3 /* (26, 10, 15) */,
  32'h3e48eba4 /* (22, 10, 15) */,
  32'h3eacaf9b /* (18, 10, 15) */,
  32'h3eacaf9b /* (14, 10, 15) */,
  32'h3e48eba4 /* (10, 10, 15) */,
  32'h3de44bb3 /* (6, 10, 15) */,
  32'h3daa3ec9 /* (2, 10, 15) */,
  32'h3d4bfe66 /* (30, 6, 15) */,
  32'h3d85e8bf /* (26, 6, 15) */,
  32'h3de44bb3 /* (22, 6, 15) */,
  32'h3e3e01e0 /* (18, 6, 15) */,
  32'h3e3e01e0 /* (14, 6, 15) */,
  32'h3de44bb3 /* (10, 6, 15) */,
  32'h3d85e8bf /* (6, 6, 15) */,
  32'h3d4bfe66 /* (2, 6, 15) */,
  32'h3d1dadb9 /* (30, 2, 15) */,
  32'h3d4bfe66 /* (26, 2, 15) */,
  32'h3daa3ec9 /* (22, 2, 15) */,
  32'h3e0adb0d /* (18, 2, 15) */,
  32'h3e0adb0d /* (14, 2, 15) */,
  32'h3daa3ec9 /* (10, 2, 15) */,
  32'h3d4bfe66 /* (6, 2, 15) */,
  32'h3d1dadb9 /* (2, 2, 15) */,
  32'h3d18e0f8 /* (30, 30, 11) */,
  32'h3d343ccb /* (26, 30, 11) */,
  32'h3d85a0b3 /* (22, 30, 11) */,
  32'h3dc55f41 /* (18, 30, 11) */,
  32'h3dc55f41 /* (14, 30, 11) */,
  32'h3d85a0b3 /* (10, 30, 11) */,
  32'h3d343ccb /* (6, 30, 11) */,
  32'h3d18e0f8 /* (2, 30, 11) */,
  32'h3d343ccb /* (30, 26, 11) */,
  32'h3d5d3b5c /* (26, 26, 11) */,
  32'h3dac23aa /* (22, 26, 11) */,
  32'h3e040b60 /* (18, 26, 11) */,
  32'h3e040b60 /* (14, 26, 11) */,
  32'h3dac23aa /* (10, 26, 11) */,
  32'h3d5d3b5c /* (6, 26, 11) */,
  32'h3d343ccb /* (2, 26, 11) */,
  32'h3d85a0b3 /* (30, 22, 11) */,
  32'h3dac23aa /* (26, 22, 11) */,
  32'h3e0ecbcd /* (22, 22, 11) */,
  32'h3e67a191 /* (18, 22, 11) */,
  32'h3e67a191 /* (14, 22, 11) */,
  32'h3e0ecbcd /* (10, 22, 11) */,
  32'h3dac23aa /* (6, 22, 11) */,
  32'h3d85a0b3 /* (2, 22, 11) */,
  32'h3dc55f41 /* (30, 18, 11) */,
  32'h3e040b60 /* (26, 18, 11) */,
  32'h3e67a191 /* (22, 18, 11) */,
  32'h3ec66134 /* (18, 18, 11) */,
  32'h3ec66134 /* (14, 18, 11) */,
  32'h3e67a191 /* (10, 18, 11) */,
  32'h3e040b60 /* (6, 18, 11) */,
  32'h3dc55f41 /* (2, 18, 11) */,
  32'h3dc55f41 /* (30, 14, 11) */,
  32'h3e040b60 /* (26, 14, 11) */,
  32'h3e67a191 /* (22, 14, 11) */,
  32'h3ec66134 /* (18, 14, 11) */,
  32'h3ec66134 /* (14, 14, 11) */,
  32'h3e67a191 /* (10, 14, 11) */,
  32'h3e040b60 /* (6, 14, 11) */,
  32'h3dc55f41 /* (2, 14, 11) */,
  32'h3d85a0b3 /* (30, 10, 11) */,
  32'h3dac23aa /* (26, 10, 11) */,
  32'h3e0ecbcd /* (22, 10, 11) */,
  32'h3e67a191 /* (18, 10, 11) */,
  32'h3e67a191 /* (14, 10, 11) */,
  32'h3e0ecbcd /* (10, 10, 11) */,
  32'h3dac23aa /* (6, 10, 11) */,
  32'h3d85a0b3 /* (2, 10, 11) */,
  32'h3d343ccb /* (30, 6, 11) */,
  32'h3d5d3b5c /* (26, 6, 11) */,
  32'h3dac23aa /* (22, 6, 11) */,
  32'h3e040b60 /* (18, 6, 11) */,
  32'h3e040b60 /* (14, 6, 11) */,
  32'h3dac23aa /* (10, 6, 11) */,
  32'h3d5d3b5c /* (6, 6, 11) */,
  32'h3d343ccb /* (2, 6, 11) */,
  32'h3d18e0f8 /* (30, 2, 11) */,
  32'h3d343ccb /* (26, 2, 11) */,
  32'h3d85a0b3 /* (22, 2, 11) */,
  32'h3dc55f41 /* (18, 2, 11) */,
  32'h3dc55f41 /* (14, 2, 11) */,
  32'h3d85a0b3 /* (10, 2, 11) */,
  32'h3d343ccb /* (6, 2, 11) */,
  32'h3d18e0f8 /* (2, 2, 11) */,
  32'h3d1dd271 /* (30, 30, 7) */,
  32'h3d14b9d3 /* (26, 30, 7) */,
  32'h3d3346c6 /* (22, 30, 7) */,
  32'h3d6820b1 /* (18, 30, 7) */,
  32'h3d6820b1 /* (14, 30, 7) */,
  32'h3d3346c6 /* (10, 30, 7) */,
  32'h3d14b9d3 /* (6, 30, 7) */,
  32'h3d1dd271 /* (2, 30, 7) */,
  32'h3d14b9d3 /* (30, 26, 7) */,
  32'h3d20f672 /* (26, 26, 7) */,
  32'h3d5a2934 /* (22, 26, 7) */,
  32'h3d975464 /* (18, 26, 7) */,
  32'h3d975464 /* (14, 26, 7) */,
  32'h3d5a2934 /* (10, 26, 7) */,
  32'h3d20f672 /* (6, 26, 7) */,
  32'h3d14b9d3 /* (2, 26, 7) */,
  32'h3d3346c6 /* (30, 22, 7) */,
  32'h3d5a2934 /* (26, 22, 7) */,
  32'h3da7f0fb /* (22, 22, 7) */,
  32'h3dff6ab3 /* (18, 22, 7) */,
  32'h3dff6ab3 /* (14, 22, 7) */,
  32'h3da7f0fb /* (10, 22, 7) */,
  32'h3d5a2934 /* (6, 22, 7) */,
  32'h3d3346c6 /* (2, 22, 7) */,
  32'h3d6820b1 /* (30, 18, 7) */,
  32'h3d975464 /* (26, 18, 7) */,
  32'h3dff6ab3 /* (22, 18, 7) */,
  32'h3e528761 /* (18, 18, 7) */,
  32'h3e528761 /* (14, 18, 7) */,
  32'h3dff6ab3 /* (10, 18, 7) */,
  32'h3d975464 /* (6, 18, 7) */,
  32'h3d6820b1 /* (2, 18, 7) */,
  32'h3d6820b1 /* (30, 14, 7) */,
  32'h3d975464 /* (26, 14, 7) */,
  32'h3dff6ab3 /* (22, 14, 7) */,
  32'h3e528761 /* (18, 14, 7) */,
  32'h3e528761 /* (14, 14, 7) */,
  32'h3dff6ab3 /* (10, 14, 7) */,
  32'h3d975464 /* (6, 14, 7) */,
  32'h3d6820b1 /* (2, 14, 7) */,
  32'h3d3346c6 /* (30, 10, 7) */,
  32'h3d5a2934 /* (26, 10, 7) */,
  32'h3da7f0fb /* (22, 10, 7) */,
  32'h3dff6ab3 /* (18, 10, 7) */,
  32'h3dff6ab3 /* (14, 10, 7) */,
  32'h3da7f0fb /* (10, 10, 7) */,
  32'h3d5a2934 /* (6, 10, 7) */,
  32'h3d3346c6 /* (2, 10, 7) */,
  32'h3d14b9d3 /* (30, 6, 7) */,
  32'h3d20f672 /* (26, 6, 7) */,
  32'h3d5a2934 /* (22, 6, 7) */,
  32'h3d975464 /* (18, 6, 7) */,
  32'h3d975464 /* (14, 6, 7) */,
  32'h3d5a2934 /* (10, 6, 7) */,
  32'h3d20f672 /* (6, 6, 7) */,
  32'h3d14b9d3 /* (2, 6, 7) */,
  32'h3d1dd271 /* (30, 2, 7) */,
  32'h3d14b9d3 /* (26, 2, 7) */,
  32'h3d3346c6 /* (22, 2, 7) */,
  32'h3d6820b1 /* (18, 2, 7) */,
  32'h3d6820b1 /* (14, 2, 7) */,
  32'h3d3346c6 /* (10, 2, 7) */,
  32'h3d14b9d3 /* (6, 2, 7) */,
  32'h3d1dd271 /* (2, 2, 7) */,
  32'h3da3af74 /* (30, 30, 3) */,
  32'h3d271e8d /* (26, 30, 3) */,
  32'h3d162b76 /* (22, 30, 3) */,
  32'h3d2b1735 /* (18, 30, 3) */,
  32'h3d2b1735 /* (14, 30, 3) */,
  32'h3d162b76 /* (10, 30, 3) */,
  32'h3d271e8d /* (6, 30, 3) */,
  32'h3da3af74 /* (2, 30, 3) */,
  32'h3d271e8d /* (30, 26, 3) */,
  32'h3d14c14d /* (26, 26, 3) */,
  32'h3d2c3293 /* (22, 26, 3) */,
  32'h3d5a5169 /* (18, 26, 3) */,
  32'h3d5a5169 /* (14, 26, 3) */,
  32'h3d2c3293 /* (10, 26, 3) */,
  32'h3d14c14d /* (6, 26, 3) */,
  32'h3d271e8d /* (2, 26, 3) */,
  32'h3d162b76 /* (30, 22, 3) */,
  32'h3d2c3293 /* (26, 22, 3) */,
  32'h3d77904c /* (22, 22, 3) */,
  32'h3db2bcb9 /* (18, 22, 3) */,
  32'h3db2bcb9 /* (14, 22, 3) */,
  32'h3d77904c /* (10, 22, 3) */,
  32'h3d2c3293 /* (6, 22, 3) */,
  32'h3d162b76 /* (2, 22, 3) */,
  32'h3d2b1735 /* (30, 18, 3) */,
  32'h3d5a5169 /* (26, 18, 3) */,
  32'h3db2bcb9 /* (22, 18, 3) */,
  32'h3e0f3c67 /* (18, 18, 3) */,
  32'h3e0f3c67 /* (14, 18, 3) */,
  32'h3db2bcb9 /* (10, 18, 3) */,
  32'h3d5a5169 /* (6, 18, 3) */,
  32'h3d2b1735 /* (2, 18, 3) */,
  32'h3d2b1735 /* (30, 14, 3) */,
  32'h3d5a5169 /* (26, 14, 3) */,
  32'h3db2bcb9 /* (22, 14, 3) */,
  32'h3e0f3c67 /* (18, 14, 3) */,
  32'h3e0f3c67 /* (14, 14, 3) */,
  32'h3db2bcb9 /* (10, 14, 3) */,
  32'h3d5a5169 /* (6, 14, 3) */,
  32'h3d2b1735 /* (2, 14, 3) */,
  32'h3d162b76 /* (30, 10, 3) */,
  32'h3d2c3293 /* (26, 10, 3) */,
  32'h3d77904c /* (22, 10, 3) */,
  32'h3db2bcb9 /* (18, 10, 3) */,
  32'h3db2bcb9 /* (14, 10, 3) */,
  32'h3d77904c /* (10, 10, 3) */,
  32'h3d2c3293 /* (6, 10, 3) */,
  32'h3d162b76 /* (2, 10, 3) */,
  32'h3d271e8d /* (30, 6, 3) */,
  32'h3d14c14d /* (26, 6, 3) */,
  32'h3d2c3293 /* (22, 6, 3) */,
  32'h3d5a5169 /* (18, 6, 3) */,
  32'h3d5a5169 /* (14, 6, 3) */,
  32'h3d2c3293 /* (10, 6, 3) */,
  32'h3d14c14d /* (6, 6, 3) */,
  32'h3d271e8d /* (2, 6, 3) */,
  32'h3da3af74 /* (30, 2, 3) */,
  32'h3d271e8d /* (26, 2, 3) */,
  32'h3d162b76 /* (22, 2, 3) */,
  32'h3d2b1735 /* (18, 2, 3) */,
  32'h3d2b1735 /* (14, 2, 3) */,
  32'h3d162b76 /* (10, 2, 3) */,
  32'h3d271e8d /* (6, 2, 3) */,
  32'h3da3af74 /* (2, 2, 3) */,
  32'h3dbfa8df /* (29, 30, 31) */,
  32'h3d20a35e /* (25, 30, 31) */,
  32'h3d16ed42 /* (21, 30, 31) */,
  32'h3d1a0745 /* (17, 30, 31) */,
  32'h3d214ba3 /* (13, 30, 31) */,
  32'h3d11c69f /* (9, 30, 31) */,
  32'h3d59109a /* (5, 30, 31) */,
  32'h3e4aeee2 /* (1, 30, 31) */,
  32'h3d2ba889 /* (29, 26, 31) */,
  32'h3d146a43 /* (25, 26, 31) */,
  32'h3d31191b /* (21, 26, 31) */,
  32'h3d46f53f /* (17, 26, 31) */,
  32'h3d4876ff /* (13, 26, 31) */,
  32'h3d1c53e8 /* (9, 26, 31) */,
  32'h3d1a8b5a /* (5, 26, 31) */,
  32'h3d3c9698 /* (1, 26, 31) */,
  32'h3d14c0fd /* (29, 22, 31) */,
  32'h3d305430 /* (25, 22, 31) */,
  32'h3d829849 /* (21, 22, 31) */,
  32'h3da5ac70 /* (17, 22, 31) */,
  32'h3d9e7894 /* (13, 22, 31) */,
  32'h3d52081f /* (9, 22, 31) */,
  32'h3d1d9589 /* (5, 22, 31) */,
  32'h3d119771 /* (1, 22, 31) */,
  32'h3d276174 /* (29, 18, 31) */,
  32'h3d62906c /* (25, 18, 31) */,
  32'h3dc01db4 /* (21, 18, 31) */,
  32'h3e06d8bb /* (17, 18, 31) */,
  32'h3df65860 /* (13, 18, 31) */,
  32'h3d90dff9 /* (9, 18, 31) */,
  32'h3d3c7841 /* (5, 18, 31) */,
  32'h3d1e0bb6 /* (1, 18, 31) */,
  32'h3d276174 /* (29, 14, 31) */,
  32'h3d62906c /* (25, 14, 31) */,
  32'h3dc01db4 /* (21, 14, 31) */,
  32'h3e06d8bb /* (17, 14, 31) */,
  32'h3df65860 /* (13, 14, 31) */,
  32'h3d90dff9 /* (9, 14, 31) */,
  32'h3d3c7841 /* (5, 14, 31) */,
  32'h3d1e0bb6 /* (1, 14, 31) */,
  32'h3d14c0fd /* (29, 10, 31) */,
  32'h3d305430 /* (25, 10, 31) */,
  32'h3d829849 /* (21, 10, 31) */,
  32'h3da5ac70 /* (17, 10, 31) */,
  32'h3d9e7894 /* (13, 10, 31) */,
  32'h3d52081f /* (9, 10, 31) */,
  32'h3d1d9589 /* (5, 10, 31) */,
  32'h3d119771 /* (1, 10, 31) */,
  32'h3d2ba889 /* (29, 6, 31) */,
  32'h3d146a43 /* (25, 6, 31) */,
  32'h3d31191b /* (21, 6, 31) */,
  32'h3d46f53f /* (17, 6, 31) */,
  32'h3d4876ff /* (13, 6, 31) */,
  32'h3d1c53e8 /* (9, 6, 31) */,
  32'h3d1a8b5a /* (5, 6, 31) */,
  32'h3d3c9698 /* (1, 6, 31) */,
  32'h3dbfa8df /* (29, 2, 31) */,
  32'h3d20a35e /* (25, 2, 31) */,
  32'h3d16ed42 /* (21, 2, 31) */,
  32'h3d1a0745 /* (17, 2, 31) */,
  32'h3d214ba3 /* (13, 2, 31) */,
  32'h3d11c69f /* (9, 2, 31) */,
  32'h3d59109a /* (5, 2, 31) */,
  32'h3e4aeee2 /* (1, 2, 31) */,
  32'h3d3cd255 /* (29, 30, 27) */,
  32'h3d14b1c0 /* (25, 30, 27) */,
  32'h3d29823f /* (21, 30, 27) */,
  32'h3d3a7be5 /* (17, 30, 27) */,
  32'h3d3d84de /* (13, 30, 27) */,
  32'h3d18622e /* (9, 30, 27) */,
  32'h3d213c91 /* (5, 30, 27) */,
  32'h3d59109a /* (1, 30, 27) */,
  32'h3d16d305 /* (29, 26, 27) */,
  32'h3d1b2471 /* (25, 26, 27) */,
  32'h3d4d9045 /* (21, 26, 27) */,
  32'h3d73b16f /* (17, 26, 27) */,
  32'h3d700ffa /* (13, 26, 27) */,
  32'h3d2db0cc /* (9, 26, 27) */,
  32'h3d14f7ce /* (5, 26, 27) */,
  32'h3d1a8b5a /* (1, 26, 27) */,
  32'h3d2344c4 /* (29, 22, 27) */,
  32'h3d4b3dc7 /* (25, 22, 27) */,
  32'h3d9d9380 /* (21, 22, 27) */,
  32'h3dce52e6 /* (17, 22, 27) */,
  32'h3dc29629 /* (13, 22, 27) */,
  32'h3d781ae6 /* (9, 22, 27) */,
  32'h3d30fc5a /* (5, 22, 27) */,
  32'h3d1d9589 /* (1, 22, 27) */,
  32'h3d487174 /* (29, 18, 27) */,
  32'h3d8a0000 /* (25, 18, 27) */,
  32'h3deed79f /* (21, 18, 27) */,
  32'h3e2a981c /* (17, 18, 27) */,
  32'h3e1a8d8c /* (13, 18, 27) */,
  32'h3db24f8e /* (9, 18, 27) */,
  32'h3d63687e /* (5, 18, 27) */,
  32'h3d3c7841 /* (1, 18, 27) */,
  32'h3d487174 /* (29, 14, 27) */,
  32'h3d8a0000 /* (25, 14, 27) */,
  32'h3deed79f /* (21, 14, 27) */,
  32'h3e2a981c /* (17, 14, 27) */,
  32'h3e1a8d8c /* (13, 14, 27) */,
  32'h3db24f8e /* (9, 14, 27) */,
  32'h3d63687e /* (5, 14, 27) */,
  32'h3d3c7841 /* (1, 14, 27) */,
  32'h3d2344c4 /* (29, 10, 27) */,
  32'h3d4b3dc7 /* (25, 10, 27) */,
  32'h3d9d9380 /* (21, 10, 27) */,
  32'h3dce52e6 /* (17, 10, 27) */,
  32'h3dc29629 /* (13, 10, 27) */,
  32'h3d781ae6 /* (9, 10, 27) */,
  32'h3d30fc5a /* (5, 10, 27) */,
  32'h3d1d9589 /* (1, 10, 27) */,
  32'h3d16d305 /* (29, 6, 27) */,
  32'h3d1b2471 /* (25, 6, 27) */,
  32'h3d4d9045 /* (21, 6, 27) */,
  32'h3d73b16f /* (17, 6, 27) */,
  32'h3d700ffa /* (13, 6, 27) */,
  32'h3d2db0cc /* (9, 6, 27) */,
  32'h3d14f7ce /* (5, 6, 27) */,
  32'h3d1a8b5a /* (1, 6, 27) */,
  32'h3d3cd255 /* (29, 2, 27) */,
  32'h3d14b1c0 /* (25, 2, 27) */,
  32'h3d29823f /* (21, 2, 27) */,
  32'h3d3a7be5 /* (17, 2, 27) */,
  32'h3d3d84de /* (13, 2, 27) */,
  32'h3d18622e /* (9, 2, 27) */,
  32'h3d213c91 /* (5, 2, 27) */,
  32'h3d59109a /* (1, 2, 27) */,
  32'h3d12f42a /* (29, 30, 23) */,
  32'h3d26a1b5 /* (25, 30, 23) */,
  32'h3d6d9fa3 /* (21, 30, 23) */,
  32'h3d9314c2 /* (17, 30, 23) */,
  32'h3d8e358b /* (13, 30, 23) */,
  32'h3d42665b /* (9, 30, 23) */,
  32'h3d18622e /* (5, 30, 23) */,
  32'h3d11c69f /* (1, 30, 23) */,
  32'h3d215063 /* (29, 26, 23) */,
  32'h3d45eb5b /* (25, 26, 23) */,
  32'h3d9750ce /* (21, 26, 23) */,
  32'h3dc42ad0 /* (17, 26, 23) */,
  32'h3db9d5f4 /* (13, 26, 23) */,
  32'h3d6fd024 /* (9, 26, 23) */,
  32'h3d2db0cc /* (5, 26, 23) */,
  32'h3d1c53e8 /* (1, 26, 23) */,
  32'h3d5dae2c /* (29, 22, 23) */,
  32'h3d94014f /* (25, 22, 23) */,
  32'h3df71c69 /* (21, 22, 23) */,
  32'h3e2b3653 /* (17, 22, 23) */,
  32'h3e1d56b2 /* (13, 22, 23) */,
  32'h3dbbc730 /* (9, 22, 23) */,
  32'h3d781ae6 /* (5, 22, 23) */,
  32'h3d52081f /* (1, 22, 23) */,
  32'h3d9b2a7b /* (29, 18, 23) */,
  32'h3ddc09d8 /* (25, 18, 23) */,
  32'h3e458f30 /* (21, 18, 23) */,
  32'h3e91e4f8 /* (17, 18, 23) */,
  32'h3e821787 /* (13, 18, 23) */,
  32'h3e10cac5 /* (9, 18, 23) */,
  32'h3db24f8e /* (5, 18, 23) */,
  32'h3d90dff9 /* (1, 18, 23) */,
  32'h3d9b2a7b /* (29, 14, 23) */,
  32'h3ddc09d8 /* (25, 14, 23) */,
  32'h3e458f30 /* (21, 14, 23) */,
  32'h3e91e4f8 /* (17, 14, 23) */,
  32'h3e821787 /* (13, 14, 23) */,
  32'h3e10cac5 /* (9, 14, 23) */,
  32'h3db24f8e /* (5, 14, 23) */,
  32'h3d90dff9 /* (1, 14, 23) */,
  32'h3d5dae2c /* (29, 10, 23) */,
  32'h3d94014f /* (25, 10, 23) */,
  32'h3df71c69 /* (21, 10, 23) */,
  32'h3e2b3653 /* (17, 10, 23) */,
  32'h3e1d56b2 /* (13, 10, 23) */,
  32'h3dbbc730 /* (9, 10, 23) */,
  32'h3d781ae6 /* (5, 10, 23) */,
  32'h3d52081f /* (1, 10, 23) */,
  32'h3d215063 /* (29, 6, 23) */,
  32'h3d45eb5b /* (25, 6, 23) */,
  32'h3d9750ce /* (21, 6, 23) */,
  32'h3dc42ad0 /* (17, 6, 23) */,
  32'h3db9d5f4 /* (13, 6, 23) */,
  32'h3d6fd024 /* (9, 6, 23) */,
  32'h3d2db0cc /* (5, 6, 23) */,
  32'h3d1c53e8 /* (1, 6, 23) */,
  32'h3d12f42a /* (29, 2, 23) */,
  32'h3d26a1b5 /* (25, 2, 23) */,
  32'h3d6d9fa3 /* (21, 2, 23) */,
  32'h3d9314c2 /* (17, 2, 23) */,
  32'h3d8e358b /* (13, 2, 23) */,
  32'h3d42665b /* (9, 2, 23) */,
  32'h3d18622e /* (5, 2, 23) */,
  32'h3d11c69f /* (1, 2, 23) */,
  32'h3d29e985 /* (29, 30, 19) */,
  32'h3d6129ae /* (25, 30, 19) */,
  32'h3dba5db4 /* (21, 30, 19) */,
  32'h3e003b1e /* (17, 30, 19) */,
  32'h3dec70da /* (13, 30, 19) */,
  32'h3d8e358b /* (9, 30, 19) */,
  32'h3d3d84de /* (5, 30, 19) */,
  32'h3d214ba3 /* (1, 30, 19) */,
  32'h3d54a03b /* (29, 26, 19) */,
  32'h3d90c8a7 /* (25, 26, 19) */,
  32'h3df74dbc /* (21, 26, 19) */,
  32'h3e2ea39a /* (17, 26, 19) */,
  32'h3e1f113d /* (13, 26, 19) */,
  32'h3db9d5f4 /* (9, 26, 19) */,
  32'h3d700ffa /* (5, 26, 19) */,
  32'h3d4876ff /* (1, 26, 19) */,
  32'h3da99659 /* (29, 22, 19) */,
  32'h3defa49b /* (25, 22, 19) */,
  32'h3e562fb1 /* (21, 22, 19) */,
  32'h3e9d80fb /* (17, 22, 19) */,
  32'h3e8cbae1 /* (13, 22, 19) */,
  32'h3e1d56b2 /* (9, 22, 19) */,
  32'h3dc29629 /* (5, 22, 19) */,
  32'h3d9e7894 /* (1, 22, 19) */,
  32'h3e04d0b8 /* (29, 18, 19) */,
  32'h3e41f14c /* (25, 18, 19) */,
  32'h3eb517ce /* (21, 18, 19) */,
  32'h3f0af24f /* (17, 18, 19) */,
  32'h3ef33ce4 /* (13, 18, 19) */,
  32'h3e821787 /* (9, 18, 19) */,
  32'h3e1a8d8c /* (5, 18, 19) */,
  32'h3df65860 /* (1, 18, 19) */,
  32'h3e04d0b8 /* (29, 14, 19) */,
  32'h3e41f14c /* (25, 14, 19) */,
  32'h3eb517ce /* (21, 14, 19) */,
  32'h3f0af24f /* (17, 14, 19) */,
  32'h3ef33ce4 /* (13, 14, 19) */,
  32'h3e821787 /* (9, 14, 19) */,
  32'h3e1a8d8c /* (5, 14, 19) */,
  32'h3df65860 /* (1, 14, 19) */,
  32'h3da99659 /* (29, 10, 19) */,
  32'h3defa49b /* (25, 10, 19) */,
  32'h3e562fb1 /* (21, 10, 19) */,
  32'h3e9d80fb /* (17, 10, 19) */,
  32'h3e8cbae1 /* (13, 10, 19) */,
  32'h3e1d56b2 /* (9, 10, 19) */,
  32'h3dc29629 /* (5, 10, 19) */,
  32'h3d9e7894 /* (1, 10, 19) */,
  32'h3d54a03b /* (29, 6, 19) */,
  32'h3d90c8a7 /* (25, 6, 19) */,
  32'h3df74dbc /* (21, 6, 19) */,
  32'h3e2ea39a /* (17, 6, 19) */,
  32'h3e1f113d /* (13, 6, 19) */,
  32'h3db9d5f4 /* (9, 6, 19) */,
  32'h3d700ffa /* (5, 6, 19) */,
  32'h3d4876ff /* (1, 6, 19) */,
  32'h3d29e985 /* (29, 2, 19) */,
  32'h3d6129ae /* (25, 2, 19) */,
  32'h3dba5db4 /* (21, 2, 19) */,
  32'h3e003b1e /* (17, 2, 19) */,
  32'h3dec70da /* (13, 2, 19) */,
  32'h3d8e358b /* (9, 2, 19) */,
  32'h3d3d84de /* (5, 2, 19) */,
  32'h3d214ba3 /* (1, 2, 19) */,
  32'h3d240321 /* (29, 30, 15) */,
  32'h3d62f778 /* (25, 30, 15) */,
  32'h3dc59b81 /* (21, 30, 15) */,
  32'h3e0de5f8 /* (17, 30, 15) */,
  32'h3e003b1e /* (13, 30, 15) */,
  32'h3d9314c2 /* (9, 30, 15) */,
  32'h3d3a7be5 /* (5, 30, 15) */,
  32'h3d1a0745 /* (1, 30, 15) */,
  32'h3d54ba37 /* (29, 26, 15) */,
  32'h3d95be73 /* (25, 26, 15) */,
  32'h3e0533d0 /* (21, 26, 15) */,
  32'h3e430b11 /* (17, 26, 15) */,
  32'h3e2ea39a /* (13, 26, 15) */,
  32'h3dc42ad0 /* (9, 26, 15) */,
  32'h3d73b16f /* (5, 26, 15) */,
  32'h3d46f53f /* (1, 26, 15) */,
  32'h3db22d06 /* (29, 22, 15) */,
  32'h3e009a19 /* (25, 22, 15) */,
  32'h3e6c6ac0 /* (21, 22, 15) */,
  32'h3eb2925b /* (17, 22, 15) */,
  32'h3e9d80fb /* (13, 22, 15) */,
  32'h3e2b3653 /* (9, 22, 15) */,
  32'h3dce52e6 /* (5, 22, 15) */,
  32'h3da5ac70 /* (1, 22, 15) */,
  32'h3e11d12f /* (29, 18, 15) */,
  32'h3e57a44b /* (25, 18, 15) */,
  32'h3eccf8ff /* (21, 18, 15) */,
  32'h3f202f9a /* (17, 18, 15) */,
  32'h3f0af24f /* (13, 18, 15) */,
  32'h3e91e4f8 /* (9, 18, 15) */,
  32'h3e2a981c /* (5, 18, 15) */,
  32'h3e06d8bb /* (1, 18, 15) */,
  32'h3e11d12f /* (29, 14, 15) */,
  32'h3e57a44b /* (25, 14, 15) */,
  32'h3eccf8ff /* (21, 14, 15) */,
  32'h3f202f9a /* (17, 14, 15) */,
  32'h3f0af24f /* (13, 14, 15) */,
  32'h3e91e4f8 /* (9, 14, 15) */,
  32'h3e2a981c /* (5, 14, 15) */,
  32'h3e06d8bb /* (1, 14, 15) */,
  32'h3db22d06 /* (29, 10, 15) */,
  32'h3e009a19 /* (25, 10, 15) */,
  32'h3e6c6ac0 /* (21, 10, 15) */,
  32'h3eb2925b /* (17, 10, 15) */,
  32'h3e9d80fb /* (13, 10, 15) */,
  32'h3e2b3653 /* (9, 10, 15) */,
  32'h3dce52e6 /* (5, 10, 15) */,
  32'h3da5ac70 /* (1, 10, 15) */,
  32'h3d54ba37 /* (29, 6, 15) */,
  32'h3d95be73 /* (25, 6, 15) */,
  32'h3e0533d0 /* (21, 6, 15) */,
  32'h3e430b11 /* (17, 6, 15) */,
  32'h3e2ea39a /* (13, 6, 15) */,
  32'h3dc42ad0 /* (9, 6, 15) */,
  32'h3d73b16f /* (5, 6, 15) */,
  32'h3d46f53f /* (1, 6, 15) */,
  32'h3d240321 /* (29, 2, 15) */,
  32'h3d62f778 /* (25, 2, 15) */,
  32'h3dc59b81 /* (21, 2, 15) */,
  32'h3e0de5f8 /* (17, 2, 15) */,
  32'h3e003b1e /* (13, 2, 15) */,
  32'h3d9314c2 /* (9, 2, 15) */,
  32'h3d3a7be5 /* (5, 2, 15) */,
  32'h3d1a0745 /* (1, 2, 15) */,
  32'h3d1c5f03 /* (29, 30, 11) */,
  32'h3d42a7b8 /* (25, 30, 11) */,
  32'h3d96eb50 /* (21, 30, 11) */,
  32'h3dc59b81 /* (17, 30, 11) */,
  32'h3dba5db4 /* (13, 30, 11) */,
  32'h3d6d9fa3 /* (9, 30, 11) */,
  32'h3d29823f /* (5, 30, 11) */,
  32'h3d16ed42 /* (1, 30, 11) */,
  32'h3d39bb76 /* (29, 26, 11) */,
  32'h3d71ecf9 /* (25, 26, 11) */,
  32'h3dc480ba /* (21, 26, 11) */,
  32'h3e0533d0 /* (17, 26, 11) */,
  32'h3df74dbc /* (13, 26, 11) */,
  32'h3d9750ce /* (9, 26, 11) */,
  32'h3d4d9045 /* (5, 26, 11) */,
  32'h3d31191b /* (1, 26, 11) */,
  32'h3d8ae43c /* (29, 22, 11) */,
  32'h3dbf3f1d /* (25, 22, 11) */,
  32'h3e257fc6 /* (21, 22, 11) */,
  32'h3e6c6ac0 /* (17, 22, 11) */,
  32'h3e562fb1 /* (13, 22, 11) */,
  32'h3df71c69 /* (9, 22, 11) */,
  32'h3d9d9380 /* (5, 22, 11) */,
  32'h3d829849 /* (1, 22, 11) */,
  32'h3dce7d45 /* (29, 18, 11) */,
  32'h3e14a5c9 /* (25, 18, 11) */,
  32'h3e882756 /* (21, 18, 11) */,
  32'h3eccf8ff /* (17, 18, 11) */,
  32'h3eb517ce /* (13, 18, 11) */,
  32'h3e458f30 /* (9, 18, 11) */,
  32'h3deed79f /* (5, 18, 11) */,
  32'h3dc01db4 /* (1, 18, 11) */,
  32'h3dce7d45 /* (29, 14, 11) */,
  32'h3e14a5c9 /* (25, 14, 11) */,
  32'h3e882756 /* (21, 14, 11) */,
  32'h3eccf8ff /* (17, 14, 11) */,
  32'h3eb517ce /* (13, 14, 11) */,
  32'h3e458f30 /* (9, 14, 11) */,
  32'h3deed79f /* (5, 14, 11) */,
  32'h3dc01db4 /* (1, 14, 11) */,
  32'h3d8ae43c /* (29, 10, 11) */,
  32'h3dbf3f1d /* (25, 10, 11) */,
  32'h3e257fc6 /* (21, 10, 11) */,
  32'h3e6c6ac0 /* (17, 10, 11) */,
  32'h3e562fb1 /* (13, 10, 11) */,
  32'h3df71c69 /* (9, 10, 11) */,
  32'h3d9d9380 /* (5, 10, 11) */,
  32'h3d829849 /* (1, 10, 11) */,
  32'h3d39bb76 /* (29, 6, 11) */,
  32'h3d71ecf9 /* (25, 6, 11) */,
  32'h3dc480ba /* (21, 6, 11) */,
  32'h3e0533d0 /* (17, 6, 11) */,
  32'h3df74dbc /* (13, 6, 11) */,
  32'h3d9750ce /* (9, 6, 11) */,
  32'h3d4d9045 /* (5, 6, 11) */,
  32'h3d31191b /* (1, 6, 11) */,
  32'h3d1c5f03 /* (29, 2, 11) */,
  32'h3d42a7b8 /* (25, 2, 11) */,
  32'h3d96eb50 /* (21, 2, 11) */,
  32'h3dc59b81 /* (17, 2, 11) */,
  32'h3dba5db4 /* (13, 2, 11) */,
  32'h3d6d9fa3 /* (9, 2, 11) */,
  32'h3d29823f /* (5, 2, 11) */,
  32'h3d16ed42 /* (1, 2, 11) */,
  32'h3d1a2949 /* (29, 30, 7) */,
  32'h3d1777c7 /* (25, 30, 7) */,
  32'h3d42a7b8 /* (21, 30, 7) */,
  32'h3d62f778 /* (17, 30, 7) */,
  32'h3d6129ae /* (13, 30, 7) */,
  32'h3d26a1b5 /* (9, 30, 7) */,
  32'h3d14b1c0 /* (5, 30, 7) */,
  32'h3d20a35e /* (1, 30, 7) */,
  32'h3d159d44 /* (29, 26, 7) */,
  32'h3d29a602 /* (25, 26, 7) */,
  32'h3d71ecf9 /* (21, 26, 7) */,
  32'h3d95be73 /* (17, 26, 7) */,
  32'h3d90c8a7 /* (13, 26, 7) */,
  32'h3d45eb5b /* (9, 26, 7) */,
  32'h3d1b2471 /* (5, 26, 7) */,
  32'h3d146a43 /* (1, 26, 7) */,
  32'h3d387393 /* (29, 22, 7) */,
  32'h3d6deb12 /* (25, 22, 7) */,
  32'h3dbf3f1d /* (21, 22, 7) */,
  32'h3e009a19 /* (17, 22, 7) */,
  32'h3defa49b /* (13, 22, 7) */,
  32'h3d94014f /* (9, 22, 7) */,
  32'h3d4b3dc7 /* (5, 22, 7) */,
  32'h3d305430 /* (1, 22, 7) */,
  32'h3d71c736 /* (29, 18, 7) */,
  32'h3da8d240 /* (25, 18, 7) */,
  32'h3e14a5c9 /* (21, 18, 7) */,
  32'h3e57a44b /* (17, 18, 7) */,
  32'h3e41f14c /* (13, 18, 7) */,
  32'h3ddc09d8 /* (9, 18, 7) */,
  32'h3d8a0000 /* (5, 18, 7) */,
  32'h3d62906c /* (1, 18, 7) */,
  32'h3d71c736 /* (29, 14, 7) */,
  32'h3da8d240 /* (25, 14, 7) */,
  32'h3e14a5c9 /* (21, 14, 7) */,
  32'h3e57a44b /* (17, 14, 7) */,
  32'h3e41f14c /* (13, 14, 7) */,
  32'h3ddc09d8 /* (9, 14, 7) */,
  32'h3d8a0000 /* (5, 14, 7) */,
  32'h3d62906c /* (1, 14, 7) */,
  32'h3d387393 /* (29, 10, 7) */,
  32'h3d6deb12 /* (25, 10, 7) */,
  32'h3dbf3f1d /* (21, 10, 7) */,
  32'h3e009a19 /* (17, 10, 7) */,
  32'h3defa49b /* (13, 10, 7) */,
  32'h3d94014f /* (9, 10, 7) */,
  32'h3d4b3dc7 /* (5, 10, 7) */,
  32'h3d305430 /* (1, 10, 7) */,
  32'h3d159d44 /* (29, 6, 7) */,
  32'h3d29a602 /* (25, 6, 7) */,
  32'h3d71ecf9 /* (21, 6, 7) */,
  32'h3d95be73 /* (17, 6, 7) */,
  32'h3d90c8a7 /* (13, 6, 7) */,
  32'h3d45eb5b /* (9, 6, 7) */,
  32'h3d1b2471 /* (5, 6, 7) */,
  32'h3d146a43 /* (1, 6, 7) */,
  32'h3d1a2949 /* (29, 2, 7) */,
  32'h3d1777c7 /* (25, 2, 7) */,
  32'h3d42a7b8 /* (21, 2, 7) */,
  32'h3d62f778 /* (17, 2, 7) */,
  32'h3d6129ae /* (13, 2, 7) */,
  32'h3d26a1b5 /* (9, 2, 7) */,
  32'h3d14b1c0 /* (5, 2, 7) */,
  32'h3d20a35e /* (1, 2, 7) */,
  32'h3d866355 /* (29, 30, 3) */,
  32'h3d1a2949 /* (25, 30, 3) */,
  32'h3d1c5f03 /* (21, 30, 3) */,
  32'h3d240321 /* (17, 30, 3) */,
  32'h3d29e985 /* (13, 30, 3) */,
  32'h3d12f42a /* (9, 30, 3) */,
  32'h3d3cd255 /* (5, 30, 3) */,
  32'h3dbfa8df /* (1, 30, 3) */,
  32'h3d211f1b /* (29, 26, 3) */,
  32'h3d159d44 /* (25, 26, 3) */,
  32'h3d39bb76 /* (21, 26, 3) */,
  32'h3d54ba37 /* (17, 26, 3) */,
  32'h3d54a03b /* (13, 26, 3) */,
  32'h3d215063 /* (9, 26, 3) */,
  32'h3d16d305 /* (5, 26, 3) */,
  32'h3d2ba889 /* (1, 26, 3) */,
  32'h3d18cb02 /* (29, 22, 3) */,
  32'h3d387393 /* (25, 22, 3) */,
  32'h3d8ae43c /* (21, 22, 3) */,
  32'h3db22d06 /* (17, 22, 3) */,
  32'h3da99659 /* (13, 22, 3) */,
  32'h3d5dae2c /* (9, 22, 3) */,
  32'h3d2344c4 /* (5, 22, 3) */,
  32'h3d14c0fd /* (1, 22, 3) */,
  32'h3d3188e3 /* (29, 18, 3) */,
  32'h3d71c736 /* (25, 18, 3) */,
  32'h3dce7d45 /* (21, 18, 3) */,
  32'h3e11d12f /* (17, 18, 3) */,
  32'h3e04d0b8 /* (13, 18, 3) */,
  32'h3d9b2a7b /* (9, 18, 3) */,
  32'h3d487174 /* (5, 18, 3) */,
  32'h3d276174 /* (1, 18, 3) */,
  32'h3d3188e3 /* (29, 14, 3) */,
  32'h3d71c736 /* (25, 14, 3) */,
  32'h3dce7d45 /* (21, 14, 3) */,
  32'h3e11d12f /* (17, 14, 3) */,
  32'h3e04d0b8 /* (13, 14, 3) */,
  32'h3d9b2a7b /* (9, 14, 3) */,
  32'h3d487174 /* (5, 14, 3) */,
  32'h3d276174 /* (1, 14, 3) */,
  32'h3d18cb02 /* (29, 10, 3) */,
  32'h3d387393 /* (25, 10, 3) */,
  32'h3d8ae43c /* (21, 10, 3) */,
  32'h3db22d06 /* (17, 10, 3) */,
  32'h3da99659 /* (13, 10, 3) */,
  32'h3d5dae2c /* (9, 10, 3) */,
  32'h3d2344c4 /* (5, 10, 3) */,
  32'h3d14c0fd /* (1, 10, 3) */,
  32'h3d211f1b /* (29, 6, 3) */,
  32'h3d159d44 /* (25, 6, 3) */,
  32'h3d39bb76 /* (21, 6, 3) */,
  32'h3d54ba37 /* (17, 6, 3) */,
  32'h3d54a03b /* (13, 6, 3) */,
  32'h3d215063 /* (9, 6, 3) */,
  32'h3d16d305 /* (5, 6, 3) */,
  32'h3d2ba889 /* (1, 6, 3) */,
  32'h3d866355 /* (29, 2, 3) */,
  32'h3d1a2949 /* (25, 2, 3) */,
  32'h3d1c5f03 /* (21, 2, 3) */,
  32'h3d240321 /* (17, 2, 3) */,
  32'h3d29e985 /* (13, 2, 3) */,
  32'h3d12f42a /* (9, 2, 3) */,
  32'h3d3cd255 /* (5, 2, 3) */,
  32'h3dbfa8df /* (1, 2, 3) */,
  32'h3d8b1391 /* (28, 30, 31) */,
  32'h3d15ce12 /* (24, 30, 31) */,
  32'h3d1cac31 /* (20, 30, 31) */,
  32'h3d09dfab /* (16, 30, 31) */,
  32'h3d1cac31 /* (12, 30, 31) */,
  32'h3d15ce12 /* (8, 30, 31) */,
  32'h3d8b1391 /* (4, 30, 31) */,
  32'h3e709592 /* (0, 30, 31) */,
  32'h3d222a9c /* (28, 26, 31) */,
  32'h3d169650 /* (24, 26, 31) */,
  32'h3d3dc5f0 /* (20, 26, 31) */,
  32'h3d34b66a /* (16, 26, 31) */,
  32'h3d3dc5f0 /* (12, 26, 31) */,
  32'h3d169650 /* (8, 26, 31) */,
  32'h3d222a9c /* (4, 26, 31) */,
  32'h3d3f59b8 /* (0, 26, 31) */,
  32'h3d1839e3 /* (28, 22, 31) */,
  32'h3d3f0366 /* (24, 22, 31) */,
  32'h3d91435f /* (20, 22, 31) */,
  32'h3d99ac24 /* (16, 22, 31) */,
  32'h3d91435f /* (12, 22, 31) */,
  32'h3d3f0366 /* (8, 22, 31) */,
  32'h3d1839e3 /* (4, 22, 31) */,
  32'h3d1142bb /* (0, 22, 31) */,
  32'h3d303352 /* (28, 18, 31) */,
  32'h3d7e759f /* (24, 18, 31) */,
  32'h3ddbed5a /* (20, 18, 31) */,
  32'h3dff32bb /* (16, 18, 31) */,
  32'h3ddbed5a /* (12, 18, 31) */,
  32'h3d7e759f /* (8, 18, 31) */,
  32'h3d303352 /* (4, 18, 31) */,
  32'h3d1ceee6 /* (0, 18, 31) */,
  32'h3d303352 /* (28, 14, 31) */,
  32'h3d7e759f /* (24, 14, 31) */,
  32'h3ddbed5a /* (20, 14, 31) */,
  32'h3dff32bb /* (16, 14, 31) */,
  32'h3ddbed5a /* (12, 14, 31) */,
  32'h3d7e759f /* (8, 14, 31) */,
  32'h3d303352 /* (4, 14, 31) */,
  32'h3d1ceee6 /* (0, 14, 31) */,
  32'h3d1839e3 /* (28, 10, 31) */,
  32'h3d3f0366 /* (24, 10, 31) */,
  32'h3d91435f /* (20, 10, 31) */,
  32'h3d99ac24 /* (16, 10, 31) */,
  32'h3d91435f /* (12, 10, 31) */,
  32'h3d3f0366 /* (8, 10, 31) */,
  32'h3d1839e3 /* (4, 10, 31) */,
  32'h3d1142bb /* (0, 10, 31) */,
  32'h3d222a9c /* (28, 6, 31) */,
  32'h3d169650 /* (24, 6, 31) */,
  32'h3d3dc5f0 /* (20, 6, 31) */,
  32'h3d34b66a /* (16, 6, 31) */,
  32'h3d3dc5f0 /* (12, 6, 31) */,
  32'h3d169650 /* (8, 6, 31) */,
  32'h3d222a9c /* (4, 6, 31) */,
  32'h3d3f59b8 /* (0, 6, 31) */,
  32'h3d8b1391 /* (28, 2, 31) */,
  32'h3d15ce12 /* (24, 2, 31) */,
  32'h3d1cac31 /* (20, 2, 31) */,
  32'h3d09dfab /* (16, 2, 31) */,
  32'h3d1cac31 /* (12, 2, 31) */,
  32'h3d15ce12 /* (8, 2, 31) */,
  32'h3d8b1391 /* (4, 2, 31) */,
  32'h3e709592 /* (0, 2, 31) */,
  32'h3d2d8e0e /* (28, 30, 27) */,
  32'h3d149b5c /* (24, 30, 27) */,
  32'h3d346b02 /* (20, 30, 27) */,
  32'h3d28d1e5 /* (16, 30, 27) */,
  32'h3d346b02 /* (12, 30, 27) */,
  32'h3d149b5c /* (8, 30, 27) */,
  32'h3d2d8e0e /* (4, 30, 27) */,
  32'h3d5dd7d1 /* (0, 30, 27) */,
  32'h3d153e19 /* (28, 26, 27) */,
  32'h3d22af34 /* (24, 26, 27) */,
  32'h3d6007ad /* (20, 26, 27) */,
  32'h3d5f53fb /* (16, 26, 27) */,
  32'h3d6007ad /* (12, 26, 27) */,
  32'h3d22af34 /* (8, 26, 27) */,
  32'h3d153e19 /* (4, 26, 27) */,
  32'h3d1b2f33 /* (0, 26, 27) */,
  32'h3d28e3b2 /* (28, 22, 27) */,
  32'h3d5ef675 /* (24, 22, 27) */,
  32'h3db0e528 /* (20, 22, 27) */,
  32'h3dc0863e /* (16, 22, 27) */,
  32'h3db0e528 /* (12, 22, 27) */,
  32'h3d5ef675 /* (8, 22, 27) */,
  32'h3d28e3b2 /* (4, 22, 27) */,
  32'h3d1cee15 /* (0, 22, 27) */,
  32'h3d53bb31 /* (28, 18, 27) */,
  32'h3d9bc970 /* (24, 18, 27) */,
  32'h3e095be4 /* (20, 18, 27) */,
  32'h3e2205a1 /* (16, 18, 27) */,
  32'h3e095be4 /* (12, 18, 27) */,
  32'h3d9bc970 /* (8, 18, 27) */,
  32'h3d53bb31 /* (4, 18, 27) */,
  32'h3d3b0a55 /* (0, 18, 27) */,
  32'h3d53bb31 /* (28, 14, 27) */,
  32'h3d9bc970 /* (24, 14, 27) */,
  32'h3e095be4 /* (20, 14, 27) */,
  32'h3e2205a1 /* (16, 14, 27) */,
  32'h3e095be4 /* (12, 14, 27) */,
  32'h3d9bc970 /* (8, 14, 27) */,
  32'h3d53bb31 /* (4, 14, 27) */,
  32'h3d3b0a55 /* (0, 14, 27) */,
  32'h3d28e3b2 /* (28, 10, 27) */,
  32'h3d5ef675 /* (24, 10, 27) */,
  32'h3db0e528 /* (20, 10, 27) */,
  32'h3dc0863e /* (16, 10, 27) */,
  32'h3db0e528 /* (12, 10, 27) */,
  32'h3d5ef675 /* (8, 10, 27) */,
  32'h3d28e3b2 /* (4, 10, 27) */,
  32'h3d1cee15 /* (0, 10, 27) */,
  32'h3d153e19 /* (28, 6, 27) */,
  32'h3d22af34 /* (24, 6, 27) */,
  32'h3d6007ad /* (20, 6, 27) */,
  32'h3d5f53fb /* (16, 6, 27) */,
  32'h3d6007ad /* (12, 6, 27) */,
  32'h3d22af34 /* (8, 6, 27) */,
  32'h3d153e19 /* (4, 6, 27) */,
  32'h3d1b2f33 /* (0, 6, 27) */,
  32'h3d2d8e0e /* (28, 2, 27) */,
  32'h3d149b5c /* (24, 2, 27) */,
  32'h3d346b02 /* (20, 2, 27) */,
  32'h3d28d1e5 /* (16, 2, 27) */,
  32'h3d346b02 /* (12, 2, 27) */,
  32'h3d149b5c /* (8, 2, 27) */,
  32'h3d2d8e0e /* (4, 2, 27) */,
  32'h3d5dd7d1 /* (0, 2, 27) */,
  32'h3d14de35 /* (28, 30, 23) */,
  32'h3d3291f6 /* (24, 30, 23) */,
  32'h3d833332 /* (20, 30, 23) */,
  32'h3d87d16b /* (16, 30, 23) */,
  32'h3d833332 /* (12, 30, 23) */,
  32'h3d3291f6 /* (8, 30, 23) */,
  32'h3d14de35 /* (4, 30, 23) */,
  32'h3d11b684 /* (0, 30, 23) */,
  32'h3d2657dd /* (28, 26, 23) */,
  32'h3d584c0c /* (24, 26, 23) */,
  32'h3da96159 /* (20, 26, 23) */,
  32'h3db6b309 /* (16, 26, 23) */,
  32'h3da96159 /* (12, 26, 23) */,
  32'h3d584c0c /* (8, 26, 23) */,
  32'h3d2657dd /* (4, 26, 23) */,
  32'h3d1bc36a /* (0, 26, 23) */,
  32'h3d68b7a2 /* (28, 22, 23) */,
  32'h3da590e9 /* (24, 22, 23) */,
  32'h3e0cf021 /* (20, 22, 23) */,
  32'h3e21930d /* (16, 22, 23) */,
  32'h3e0cf021 /* (12, 22, 23) */,
  32'h3da590e9 /* (8, 22, 23) */,
  32'h3d68b7a2 /* (4, 22, 23) */,
  32'h3d50a575 /* (0, 22, 23) */,
  32'h3da4db8a /* (28, 18, 23) */,
  32'h3dfaaa60 /* (24, 18, 23) */,
  32'h3e654448 /* (20, 18, 23) */,
  32'h3e8b9344 /* (16, 18, 23) */,
  32'h3e654448 /* (12, 18, 23) */,
  32'h3dfaaa60 /* (8, 18, 23) */,
  32'h3da4db8a /* (4, 18, 23) */,
  32'h3d8fa52c /* (0, 18, 23) */,
  32'h3da4db8a /* (28, 14, 23) */,
  32'h3dfaaa60 /* (24, 14, 23) */,
  32'h3e654448 /* (20, 14, 23) */,
  32'h3e8b9344 /* (16, 14, 23) */,
  32'h3e654448 /* (12, 14, 23) */,
  32'h3dfaaa60 /* (8, 14, 23) */,
  32'h3da4db8a /* (4, 14, 23) */,
  32'h3d8fa52c /* (0, 14, 23) */,
  32'h3d68b7a2 /* (28, 10, 23) */,
  32'h3da590e9 /* (24, 10, 23) */,
  32'h3e0cf021 /* (20, 10, 23) */,
  32'h3e21930d /* (16, 10, 23) */,
  32'h3e0cf021 /* (12, 10, 23) */,
  32'h3da590e9 /* (8, 10, 23) */,
  32'h3d68b7a2 /* (4, 10, 23) */,
  32'h3d50a575 /* (0, 10, 23) */,
  32'h3d2657dd /* (28, 6, 23) */,
  32'h3d584c0c /* (24, 6, 23) */,
  32'h3da96159 /* (20, 6, 23) */,
  32'h3db6b309 /* (16, 6, 23) */,
  32'h3da96159 /* (12, 6, 23) */,
  32'h3d584c0c /* (8, 6, 23) */,
  32'h3d2657dd /* (4, 6, 23) */,
  32'h3d1bc36a /* (0, 6, 23) */,
  32'h3d14de35 /* (28, 2, 23) */,
  32'h3d3291f6 /* (24, 2, 23) */,
  32'h3d833332 /* (20, 2, 23) */,
  32'h3d87d16b /* (16, 2, 23) */,
  32'h3d833332 /* (12, 2, 23) */,
  32'h3d3291f6 /* (8, 2, 23) */,
  32'h3d14de35 /* (4, 2, 23) */,
  32'h3d11b684 /* (0, 2, 23) */,
  32'h3d3217f4 /* (28, 30, 19) */,
  32'h3d7b52f8 /* (24, 30, 19) */,
  32'h3dd42d31 /* (20, 30, 19) */,
  32'h3df1ae3d /* (16, 30, 19) */,
  32'h3dd42d31 /* (12, 30, 19) */,
  32'h3d7b52f8 /* (8, 30, 19) */,
  32'h3d3217f4 /* (4, 30, 19) */,
  32'h3d2045b1 /* (0, 30, 19) */,
  32'h3d601ae9 /* (28, 26, 19) */,
  32'h3da2e7a9 /* (24, 26, 19) */,
  32'h3e0dc95f /* (20, 26, 19) */,
  32'h3e2576a9 /* (16, 26, 19) */,
  32'h3e0dc95f /* (12, 26, 19) */,
  32'h3da2e7a9 /* (8, 26, 19) */,
  32'h3d601ae9 /* (4, 26, 19) */,
  32'h3d4703b2 /* (0, 26, 19) */,
  32'h3db40e50 /* (28, 22, 19) */,
  32'h3e085939 /* (24, 22, 19) */,
  32'h3e7848b5 /* (20, 22, 19) */,
  32'h3e968a40 /* (16, 22, 19) */,
  32'h3e7848b5 /* (12, 22, 19) */,
  32'h3e085939 /* (8, 22, 19) */,
  32'h3db40e50 /* (4, 22, 19) */,
  32'h3d9d248b /* (0, 22, 19) */,
  32'h3e0de89e /* (28, 18, 19) */,
  32'h3e5f05ce /* (24, 18, 19) */,
  32'h3ed441df /* (20, 18, 19) */,
  32'h3f06176f /* (16, 18, 19) */,
  32'h3ed441df /* (12, 18, 19) */,
  32'h3e5f05ce /* (8, 18, 19) */,
  32'h3e0de89e /* (4, 18, 19) */,
  32'h3df40add /* (0, 18, 19) */,
  32'h3e0de89e /* (28, 14, 19) */,
  32'h3e5f05ce /* (24, 14, 19) */,
  32'h3ed441df /* (20, 14, 19) */,
  32'h3f06176f /* (16, 14, 19) */,
  32'h3ed441df /* (12, 14, 19) */,
  32'h3e5f05ce /* (8, 14, 19) */,
  32'h3e0de89e /* (4, 14, 19) */,
  32'h3df40add /* (0, 14, 19) */,
  32'h3db40e50 /* (28, 10, 19) */,
  32'h3e085939 /* (24, 10, 19) */,
  32'h3e7848b5 /* (20, 10, 19) */,
  32'h3e968a40 /* (16, 10, 19) */,
  32'h3e7848b5 /* (12, 10, 19) */,
  32'h3e085939 /* (8, 10, 19) */,
  32'h3db40e50 /* (4, 10, 19) */,
  32'h3d9d248b /* (0, 10, 19) */,
  32'h3d601ae9 /* (28, 6, 19) */,
  32'h3da2e7a9 /* (24, 6, 19) */,
  32'h3e0dc95f /* (20, 6, 19) */,
  32'h3e2576a9 /* (16, 6, 19) */,
  32'h3e0dc95f /* (12, 6, 19) */,
  32'h3da2e7a9 /* (8, 6, 19) */,
  32'h3d601ae9 /* (4, 6, 19) */,
  32'h3d4703b2 /* (0, 6, 19) */,
  32'h3d3217f4 /* (28, 2, 19) */,
  32'h3d7b52f8 /* (24, 2, 19) */,
  32'h3dd42d31 /* (20, 2, 19) */,
  32'h3df1ae3d /* (16, 2, 19) */,
  32'h3dd42d31 /* (12, 2, 19) */,
  32'h3d7b52f8 /* (8, 2, 19) */,
  32'h3d3217f4 /* (4, 2, 19) */,
  32'h3d2045b1 /* (0, 2, 19) */,
  32'h3d2d6bba /* (28, 30, 15) */,
  32'h3d804df8 /* (24, 30, 15) */,
  32'h3de39dff /* (20, 30, 15) */,
  32'h3e06ec2e /* (16, 30, 15) */,
  32'h3de39dff /* (12, 30, 15) */,
  32'h3d804df8 /* (8, 30, 15) */,
  32'h3d2d6bba /* (4, 30, 15) */,
  32'h3d18d610 /* (0, 30, 15) */,
  32'h3d61b1de /* (28, 26, 15) */,
  32'h3daa3349 /* (24, 26, 15) */,
  32'h3e1a3a56 /* (20, 26, 15) */,
  32'h3e3a3d1a /* (16, 26, 15) */,
  32'h3e1a3a56 /* (12, 26, 15) */,
  32'h3daa3349 /* (8, 26, 15) */,
  32'h3d61b1de /* (4, 26, 15) */,
  32'h3d455011 /* (0, 26, 15) */,
  32'h3dbdf4f8 /* (28, 22, 15) */,
  32'h3e135573 /* (24, 22, 15) */,
  32'h3e89fde5 /* (20, 22, 15) */,
  32'h3eabb572 /* (16, 22, 15) */,
  32'h3e89fde5 /* (12, 22, 15) */,
  32'h3e135573 /* (8, 22, 15) */,
  32'h3dbdf4f8 /* (4, 22, 15) */,
  32'h3da42e1b /* (0, 22, 15) */,
  32'h3e1c2ca1 /* (28, 18, 15) */,
  32'h3e79034c /* (24, 18, 15) */,
  32'h3ef15f91 /* (20, 18, 15) */,
  32'h3f1b42bd /* (16, 18, 15) */,
  32'h3ef15f91 /* (12, 18, 15) */,
  32'h3e79034c /* (8, 18, 15) */,
  32'h3e1c2ca1 /* (4, 18, 15) */,
  32'h3e05899d /* (0, 18, 15) */,
  32'h3e1c2ca1 /* (28, 14, 15) */,
  32'h3e79034c /* (24, 14, 15) */,
  32'h3ef15f91 /* (20, 14, 15) */,
  32'h3f1b42bd /* (16, 14, 15) */,
  32'h3ef15f91 /* (12, 14, 15) */,
  32'h3e79034c /* (8, 14, 15) */,
  32'h3e1c2ca1 /* (4, 14, 15) */,
  32'h3e05899d /* (0, 14, 15) */,
  32'h3dbdf4f8 /* (28, 10, 15) */,
  32'h3e135573 /* (24, 10, 15) */,
  32'h3e89fde5 /* (20, 10, 15) */,
  32'h3eabb572 /* (16, 10, 15) */,
  32'h3e89fde5 /* (12, 10, 15) */,
  32'h3e135573 /* (8, 10, 15) */,
  32'h3dbdf4f8 /* (4, 10, 15) */,
  32'h3da42e1b /* (0, 10, 15) */,
  32'h3d61b1de /* (28, 6, 15) */,
  32'h3daa3349 /* (24, 6, 15) */,
  32'h3e1a3a56 /* (20, 6, 15) */,
  32'h3e3a3d1a /* (16, 6, 15) */,
  32'h3e1a3a56 /* (12, 6, 15) */,
  32'h3daa3349 /* (8, 6, 15) */,
  32'h3d61b1de /* (4, 6, 15) */,
  32'h3d455011 /* (0, 6, 15) */,
  32'h3d2d6bba /* (28, 2, 15) */,
  32'h3d804df8 /* (24, 2, 15) */,
  32'h3de39dff /* (20, 2, 15) */,
  32'h3e06ec2e /* (16, 2, 15) */,
  32'h3de39dff /* (12, 2, 15) */,
  32'h3d804df8 /* (8, 2, 15) */,
  32'h3d2d6bba /* (4, 2, 15) */,
  32'h3d18d610 /* (0, 2, 15) */,
  32'h3d21c128 /* (28, 30, 11) */,
  32'h3d558b1c /* (24, 30, 11) */,
  32'h3da96c08 /* (20, 30, 11) */,
  32'h3db86416 /* (16, 30, 11) */,
  32'h3da96c08 /* (12, 30, 11) */,
  32'h3d558b1c /* (8, 30, 11) */,
  32'h3d21c128 /* (4, 30, 11) */,
  32'h3d164ce1 /* (0, 30, 11) */,
  32'h3d41fb9f /* (28, 26, 11) */,
  32'h3d865b59 /* (24, 26, 11) */,
  32'h3ddec971 /* (20, 26, 11) */,
  32'h3dfa4afe /* (16, 26, 11) */,
  32'h3ddec971 /* (12, 26, 11) */,
  32'h3d865b59 /* (8, 26, 11) */,
  32'h3d41fb9f /* (4, 26, 11) */,
  32'h3d3013e2 /* (0, 26, 11) */,
  32'h3d92b699 /* (28, 22, 11) */,
  32'h3dd7e578 /* (24, 22, 11) */,
  32'h3e3e5baf /* (20, 22, 11) */,
  32'h3e60898b /* (16, 22, 11) */,
  32'h3e3e5baf /* (12, 22, 11) */,
  32'h3dd7e578 /* (8, 22, 11) */,
  32'h3d92b699 /* (4, 22, 11) */,
  32'h3d819abc /* (0, 22, 11) */,
  32'h3ddc0819 /* (28, 18, 11) */,
  32'h3e2a27e4 /* (24, 18, 11) */,
  32'h3e9ecc49 /* (20, 18, 11) */,
  32'h3ec4f0a1 /* (16, 18, 11) */,
  32'h3e9ecc49 /* (12, 18, 11) */,
  32'h3e2a27e4 /* (8, 18, 11) */,
  32'h3ddc0819 /* (4, 18, 11) */,
  32'h3dbe661f /* (0, 18, 11) */,
  32'h3ddc0819 /* (28, 14, 11) */,
  32'h3e2a27e4 /* (24, 14, 11) */,
  32'h3e9ecc49 /* (20, 14, 11) */,
  32'h3ec4f0a1 /* (16, 14, 11) */,
  32'h3e9ecc49 /* (12, 14, 11) */,
  32'h3e2a27e4 /* (8, 14, 11) */,
  32'h3ddc0819 /* (4, 14, 11) */,
  32'h3dbe661f /* (0, 14, 11) */,
  32'h3d92b699 /* (28, 10, 11) */,
  32'h3dd7e578 /* (24, 10, 11) */,
  32'h3e3e5baf /* (20, 10, 11) */,
  32'h3e60898b /* (16, 10, 11) */,
  32'h3e3e5baf /* (12, 10, 11) */,
  32'h3dd7e578 /* (8, 10, 11) */,
  32'h3d92b699 /* (4, 10, 11) */,
  32'h3d819abc /* (0, 10, 11) */,
  32'h3d41fb9f /* (28, 6, 11) */,
  32'h3d865b59 /* (24, 6, 11) */,
  32'h3ddec971 /* (20, 6, 11) */,
  32'h3dfa4afe /* (16, 6, 11) */,
  32'h3ddec971 /* (12, 6, 11) */,
  32'h3d865b59 /* (8, 6, 11) */,
  32'h3d41fb9f /* (4, 6, 11) */,
  32'h3d3013e2 /* (0, 6, 11) */,
  32'h3d21c128 /* (28, 2, 11) */,
  32'h3d558b1c /* (24, 2, 11) */,
  32'h3da96c08 /* (20, 2, 11) */,
  32'h3db86416 /* (16, 2, 11) */,
  32'h3da96c08 /* (12, 2, 11) */,
  32'h3d558b1c /* (8, 2, 11) */,
  32'h3d21c128 /* (4, 2, 11) */,
  32'h3d164ce1 /* (0, 2, 11) */,
  32'h3d16c6a3 /* (28, 30, 7) */,
  32'h3d1d59b0 /* (24, 30, 7) */,
  32'h3d530d8e /* (20, 30, 7) */,
  32'h3d4f6a6e /* (16, 30, 7) */,
  32'h3d530d8e /* (12, 30, 7) */,
  32'h3d1d59b0 /* (8, 30, 7) */,
  32'h3d16c6a3 /* (4, 30, 7) */,
  32'h3d21b235 /* (0, 30, 7) */,
  32'h3d17902e /* (28, 26, 7) */,
  32'h3d35cd98 /* (24, 26, 7) */,
  32'h3d859348 /* (20, 26, 7) */,
  32'h3d8a46e7 /* (16, 26, 7) */,
  32'h3d859348 /* (12, 26, 7) */,
  32'h3d35cd98 /* (8, 26, 7) */,
  32'h3d17902e /* (4, 26, 7) */,
  32'h3d1459dd /* (0, 26, 7) */,
  32'h3d404057 /* (28, 22, 7) */,
  32'h3d83c517 /* (24, 22, 7) */,
  32'h3dd85675 /* (20, 22, 7) */,
  32'h3df142da /* (16, 22, 7) */,
  32'h3dd85675 /* (12, 22, 7) */,
  32'h3d83c517 /* (8, 22, 7) */,
  32'h3d404057 /* (4, 22, 7) */,
  32'h3d2f5f5a /* (0, 22, 7) */,
  32'h3d800deb /* (28, 18, 7) */,
  32'h3dbf672f /* (24, 18, 7) */,
  32'h3e2baf50 /* (20, 18, 7) */,
  32'h3e4d7ce8 /* (16, 18, 7) */,
  32'h3e2baf50 /* (12, 18, 7) */,
  32'h3dbf672f /* (8, 18, 7) */,
  32'h3d800deb /* (4, 18, 7) */,
  32'h3d60bf24 /* (0, 18, 7) */,
  32'h3d800deb /* (28, 14, 7) */,
  32'h3dbf672f /* (24, 14, 7) */,
  32'h3e2baf50 /* (20, 14, 7) */,
  32'h3e4d7ce8 /* (16, 14, 7) */,
  32'h3e2baf50 /* (12, 14, 7) */,
  32'h3dbf672f /* (8, 14, 7) */,
  32'h3d800deb /* (4, 14, 7) */,
  32'h3d60bf24 /* (0, 14, 7) */,
  32'h3d404057 /* (28, 10, 7) */,
  32'h3d83c517 /* (24, 10, 7) */,
  32'h3dd85675 /* (20, 10, 7) */,
  32'h3df142da /* (16, 10, 7) */,
  32'h3dd85675 /* (12, 10, 7) */,
  32'h3d83c517 /* (8, 10, 7) */,
  32'h3d404057 /* (4, 10, 7) */,
  32'h3d2f5f5a /* (0, 10, 7) */,
  32'h3d17902e /* (28, 6, 7) */,
  32'h3d35cd98 /* (24, 6, 7) */,
  32'h3d859348 /* (20, 6, 7) */,
  32'h3d8a46e7 /* (16, 6, 7) */,
  32'h3d859348 /* (12, 6, 7) */,
  32'h3d35cd98 /* (8, 6, 7) */,
  32'h3d17902e /* (4, 6, 7) */,
  32'h3d1459dd /* (0, 6, 7) */,
  32'h3d16c6a3 /* (28, 2, 7) */,
  32'h3d1d59b0 /* (24, 2, 7) */,
  32'h3d530d8e /* (20, 2, 7) */,
  32'h3d4f6a6e /* (16, 2, 7) */,
  32'h3d530d8e /* (12, 2, 7) */,
  32'h3d1d59b0 /* (8, 2, 7) */,
  32'h3d16c6a3 /* (4, 2, 7) */,
  32'h3d21b235 /* (0, 2, 7) */,
  32'h3d5defd3 /* (28, 30, 3) */,
  32'h3d13e9f7 /* (24, 30, 3) */,
  32'h3d23d587 /* (20, 30, 3) */,
  32'h3d13661d /* (16, 30, 3) */,
  32'h3d23d587 /* (12, 30, 3) */,
  32'h3d13e9f7 /* (8, 30, 3) */,
  32'h3d5defd3 /* (4, 30, 3) */,
  32'h3dcbea25 /* (0, 30, 3) */,
  32'h3d1b3fff /* (28, 26, 3) */,
  32'h3d19bf4b /* (24, 26, 3) */,
  32'h3d48406d /* (20, 26, 3) */,
  32'h3d41d3ae /* (16, 26, 3) */,
  32'h3d48406d /* (12, 26, 3) */,
  32'h3d19bf4b /* (8, 26, 3) */,
  32'h3d1b3fff /* (4, 26, 3) */,
  32'h3d2d5b95 /* (0, 26, 3) */,
  32'h3d1cff11 /* (28, 22, 3) */,
  32'h3d48bc7e /* (24, 22, 3) */,
  32'h3d9aff71 /* (20, 22, 3) */,
  32'h3da59d10 /* (16, 22, 3) */,
  32'h3d9aff71 /* (12, 22, 3) */,
  32'h3d48bc7e /* (8, 22, 3) */,
  32'h3d1cff11 /* (4, 22, 3) */,
  32'h3d144f19 /* (0, 22, 3) */,
  32'h3d3b1e93 /* (28, 18, 3) */,
  32'h3d880501 /* (24, 18, 3) */,
  32'h3decc5e8 /* (20, 18, 3) */,
  32'h3e0a27e7 /* (16, 18, 3) */,
  32'h3decc5e8 /* (12, 18, 3) */,
  32'h3d880501 /* (8, 18, 3) */,
  32'h3d3b1e93 /* (4, 18, 3) */,
  32'h3d262b6e /* (0, 18, 3) */,
  32'h3d3b1e93 /* (28, 14, 3) */,
  32'h3d880501 /* (24, 14, 3) */,
  32'h3decc5e8 /* (20, 14, 3) */,
  32'h3e0a27e7 /* (16, 14, 3) */,
  32'h3decc5e8 /* (12, 14, 3) */,
  32'h3d880501 /* (8, 14, 3) */,
  32'h3d3b1e93 /* (4, 14, 3) */,
  32'h3d262b6e /* (0, 14, 3) */,
  32'h3d1cff11 /* (28, 10, 3) */,
  32'h3d48bc7e /* (24, 10, 3) */,
  32'h3d9aff71 /* (20, 10, 3) */,
  32'h3da59d10 /* (16, 10, 3) */,
  32'h3d9aff71 /* (12, 10, 3) */,
  32'h3d48bc7e /* (8, 10, 3) */,
  32'h3d1cff11 /* (4, 10, 3) */,
  32'h3d144f19 /* (0, 10, 3) */,
  32'h3d1b3fff /* (28, 6, 3) */,
  32'h3d19bf4b /* (24, 6, 3) */,
  32'h3d48406d /* (20, 6, 3) */,
  32'h3d41d3ae /* (16, 6, 3) */,
  32'h3d48406d /* (12, 6, 3) */,
  32'h3d19bf4b /* (8, 6, 3) */,
  32'h3d1b3fff /* (4, 6, 3) */,
  32'h3d2d5b95 /* (0, 6, 3) */,
  32'h3d5defd3 /* (28, 2, 3) */,
  32'h3d13e9f7 /* (24, 2, 3) */,
  32'h3d23d587 /* (20, 2, 3) */,
  32'h3d13661d /* (16, 2, 3) */,
  32'h3d23d587 /* (12, 2, 3) */,
  32'h3d13e9f7 /* (8, 2, 3) */,
  32'h3d5defd3 /* (4, 2, 3) */,
  32'h3dcbea25 /* (0, 2, 3) */,
  32'h3deb372d /* (31, 29, 31) */,
  32'h3d45ae9a /* (27, 29, 31) */,
  32'h3d126006 /* (23, 29, 31) */,
  32'h3d269671 /* (19, 29, 31) */,
  32'h3d202be8 /* (15, 29, 31) */,
  32'h3d1a3ccf /* (11, 29, 31) */,
  32'h3d1c3652 /* (7, 29, 31) */,
  32'h3d960c3c /* (3, 29, 31) */,
  32'h3d2402bf /* (31, 25, 31) */,
  32'h3d151e01 /* (27, 25, 31) */,
  32'h3d245baa /* (23, 25, 31) */,
  32'h3d5c17b6 /* (19, 25, 31) */,
  32'h3d5d3ed0 /* (15, 25, 31) */,
  32'h3d3efe62 /* (11, 25, 31) */,
  32'h3d167b79 /* (7, 25, 31) */,
  32'h3d1c3652 /* (3, 25, 31) */,
  32'h3d151591 /* (31, 21, 31) */,
  32'h3d26c9db /* (27, 21, 31) */,
  32'h3d68852c /* (23, 21, 31) */,
  32'h3db58f74 /* (19, 21, 31) */,
  32'h3dc031e4 /* (15, 21, 31) */,
  32'h3d9352ec /* (11, 21, 31) */,
  32'h3d3efe62 /* (7, 21, 31) */,
  32'h3d1a3ccf /* (3, 21, 31) */,
  32'h3d167d01 /* (31, 17, 31) */,
  32'h3d35f880 /* (27, 17, 31) */,
  32'h3d8f3655 /* (23, 17, 31) */,
  32'h3df92d6c /* (19, 17, 31) */,
  32'h3e09bd27 /* (15, 17, 31) */,
  32'h3dc031e4 /* (11, 17, 31) */,
  32'h3d5d3ed0 /* (7, 17, 31) */,
  32'h3d202be8 /* (3, 17, 31) */,
  32'h3d1e42f1 /* (31, 13, 31) */,
  32'h3d398f3f /* (27, 13, 31) */,
  32'h3d8ac476 /* (23, 13, 31) */,
  32'h3de602d9 /* (19, 13, 31) */,
  32'h3df92d6c /* (15, 13, 31) */,
  32'h3db58f74 /* (11, 13, 31) */,
  32'h3d5c17b6 /* (7, 13, 31) */,
  32'h3d269671 /* (3, 13, 31) */,
  32'h3d11a602 /* (31, 9, 31) */,
  32'h3d170f20 /* (27, 9, 31) */,
  32'h3d3ee791 /* (23, 9, 31) */,
  32'h3d8ac476 /* (19, 9, 31) */,
  32'h3d8f3655 /* (15, 9, 31) */,
  32'h3d68852c /* (11, 9, 31) */,
  32'h3d245baa /* (7, 9, 31) */,
  32'h3d126006 /* (3, 9, 31) */,
  32'h3d6890ff /* (31, 5, 31) */,
  32'h3d249f29 /* (27, 5, 31) */,
  32'h3d170f20 /* (23, 5, 31) */,
  32'h3d398f3f /* (19, 5, 31) */,
  32'h3d35f880 /* (15, 5, 31) */,
  32'h3d26c9db /* (11, 5, 31) */,
  32'h3d151e01 /* (7, 5, 31) */,
  32'h3d45ae9a /* (3, 5, 31) */,
  32'h3ec3aed4 /* (31, 1, 31) */,
  32'h3d6890ff /* (27, 1, 31) */,
  32'h3d11a602 /* (23, 1, 31) */,
  32'h3d1e42f1 /* (19, 1, 31) */,
  32'h3d167d01 /* (15, 1, 31) */,
  32'h3d151591 /* (11, 1, 31) */,
  32'h3d2402bf /* (7, 1, 31) */,
  32'h3deb372d /* (3, 1, 31) */,
  32'h3d45ae9a /* (31, 29, 27) */,
  32'h3d1ccb4c /* (27, 29, 27) */,
  32'h3d1addce /* (23, 29, 27) */,
  32'h3d4466f8 /* (19, 29, 27) */,
  32'h3d424fe8 /* (15, 29, 27) */,
  32'h3d2e4aa1 /* (11, 29, 27) */,
  32'h3d147808 /* (7, 29, 27) */,
  32'h3d314afb /* (3, 29, 27) */,
  32'h3d151e01 /* (31, 25, 27) */,
  32'h3d170afd /* (27, 25, 27) */,
  32'h3d39ba58 /* (23, 25, 27) */,
  32'h3d849ae2 /* (19, 25, 27) */,
  32'h3d880917 /* (15, 25, 27) */,
  32'h3d5ff008 /* (11, 25, 27) */,
  32'h3d21f168 /* (7, 25, 27) */,
  32'h3d147808 /* (3, 25, 27) */,
  32'h3d26c9db /* (31, 21, 27) */,
  32'h3d3fb488 /* (27, 21, 27) */,
  32'h3d8b02ad /* (23, 21, 27) */,
  32'h3de04254 /* (19, 21, 27) */,
  32'h3df05994 /* (15, 21, 27) */,
  32'h3db345e2 /* (11, 21, 27) */,
  32'h3d5ff008 /* (7, 21, 27) */,
  32'h3d2e4aa1 /* (3, 21, 27) */,
  32'h3d35f880 /* (31, 17, 27) */,
  32'h3d5e11d0 /* (27, 17, 27) */,
  32'h3db198fc /* (23, 17, 27) */,
  32'h3e1d0a10 /* (19, 17, 27) */,
  32'h3e2edbb4 /* (15, 17, 27) */,
  32'h3df05994 /* (11, 17, 27) */,
  32'h3d880917 /* (7, 17, 27) */,
  32'h3d424fe8 /* (3, 17, 27) */,
  32'h3d398f3f /* (31, 13, 27) */,
  32'h3d5ce99d /* (27, 13, 27) */,
  32'h3da95898 /* (23, 13, 27) */,
  32'h3e0f99f2 /* (19, 13, 27) */,
  32'h3e1d0a10 /* (15, 13, 27) */,
  32'h3de04254 /* (11, 13, 27) */,
  32'h3d849ae2 /* (7, 13, 27) */,
  32'h3d4466f8 /* (3, 13, 27) */,
  32'h3d170f20 /* (31, 9, 27) */,
  32'h3d24f869 /* (27, 9, 27) */,
  32'h3d5e7d3b /* (23, 9, 27) */,
  32'h3da95898 /* (19, 9, 27) */,
  32'h3db198fc /* (15, 9, 27) */,
  32'h3d8b02ad /* (11, 9, 27) */,
  32'h3d39ba58 /* (7, 9, 27) */,
  32'h3d1addce /* (3, 9, 27) */,
  32'h3d249f29 /* (31, 5, 27) */,
  32'h3d15ac37 /* (27, 5, 27) */,
  32'h3d24f869 /* (23, 5, 27) */,
  32'h3d5ce99d /* (19, 5, 27) */,
  32'h3d5e11d0 /* (15, 5, 27) */,
  32'h3d3fb488 /* (11, 5, 27) */,
  32'h3d170afd /* (7, 5, 27) */,
  32'h3d1ccb4c /* (3, 5, 27) */,
  32'h3d6890ff /* (31, 1, 27) */,
  32'h3d249f29 /* (27, 1, 27) */,
  32'h3d170f20 /* (23, 1, 27) */,
  32'h3d398f3f /* (19, 1, 27) */,
  32'h3d35f880 /* (15, 1, 27) */,
  32'h3d26c9db /* (11, 1, 27) */,
  32'h3d151e01 /* (7, 1, 27) */,
  32'h3d45ae9a /* (3, 1, 27) */,
  32'h3d126006 /* (31, 29, 23) */,
  32'h3d1addce /* (27, 29, 23) */,
  32'h3d48821f /* (23, 29, 23) */,
  32'h3d942dc4 /* (19, 29, 23) */,
  32'h3d99caa3 /* (15, 29, 23) */,
  32'h3d767d5d /* (11, 29, 23) */,
  32'h3d2aad03 /* (7, 29, 23) */,
  32'h3d144047 /* (3, 29, 23) */,
  32'h3d245baa /* (31, 25, 23) */,
  32'h3d39ba58 /* (27, 25, 23) */,
  32'h3d8354ed /* (23, 25, 23) */,
  32'h3dcf79e9 /* (19, 25, 23) */,
  32'h3ddc94c6 /* (15, 25, 23) */,
  32'h3da777c1 /* (11, 25, 23) */,
  32'h3d563bcb /* (7, 25, 23) */,
  32'h3d2aad03 /* (3, 25, 23) */,
  32'h3d68852c /* (31, 21, 23) */,
  32'h3d8b02ad /* (27, 21, 23) */,
  32'h3dd6aa1b /* (23, 21, 23) */,
  32'h3e37494b /* (19, 21, 23) */,
  32'h3e49046a /* (15, 21, 23) */,
  32'h3e0ea5fd /* (11, 21, 23) */,
  32'h3da777c1 /* (7, 21, 23) */,
  32'h3d767d5d /* (3, 21, 23) */,
  32'h3d8f3655 /* (31, 17, 23) */,
  32'h3db198fc /* (27, 17, 23) */,
  32'h3e123783 /* (23, 17, 23) */,
  32'h3e8557f4 /* (19, 17, 23) */,
  32'h3e969108 /* (15, 17, 23) */,
  32'h3e49046a /* (11, 17, 23) */,
  32'h3ddc94c6 /* (7, 17, 23) */,
  32'h3d99caa3 /* (3, 17, 23) */,
  32'h3d8ac476 /* (31, 13, 23) */,
  32'h3da95898 /* (27, 13, 23) */,
  32'h3e076ebd /* (23, 13, 23) */,
  32'h3e6f82ab /* (19, 13, 23) */,
  32'h3e8557f4 /* (15, 13, 23) */,
  32'h3e37494b /* (11, 13, 23) */,
  32'h3dcf79e9 /* (7, 13, 23) */,
  32'h3d942dc4 /* (3, 13, 23) */,
  32'h3d3ee791 /* (31, 9, 23) */,
  32'h3d5e7d3b /* (27, 9, 23) */,
  32'h3da4cfbf /* (23, 9, 23) */,
  32'h3e076ebd /* (19, 9, 23) */,
  32'h3e123783 /* (15, 9, 23) */,
  32'h3dd6aa1b /* (11, 9, 23) */,
  32'h3d8354ed /* (7, 9, 23) */,
  32'h3d48821f /* (3, 9, 23) */,
  32'h3d170f20 /* (31, 5, 23) */,
  32'h3d24f869 /* (27, 5, 23) */,
  32'h3d5e7d3b /* (23, 5, 23) */,
  32'h3da95898 /* (19, 5, 23) */,
  32'h3db198fc /* (15, 5, 23) */,
  32'h3d8b02ad /* (11, 5, 23) */,
  32'h3d39ba58 /* (7, 5, 23) */,
  32'h3d1addce /* (3, 5, 23) */,
  32'h3d11a602 /* (31, 1, 23) */,
  32'h3d170f20 /* (27, 1, 23) */,
  32'h3d3ee791 /* (23, 1, 23) */,
  32'h3d8ac476 /* (19, 1, 23) */,
  32'h3d8f3655 /* (15, 1, 23) */,
  32'h3d68852c /* (11, 1, 23) */,
  32'h3d245baa /* (7, 1, 23) */,
  32'h3d126006 /* (3, 1, 23) */,
  32'h3d269671 /* (31, 29, 19) */,
  32'h3d4466f8 /* (27, 29, 19) */,
  32'h3d942dc4 /* (23, 29, 19) */,
  32'h3df79892 /* (19, 29, 19) */,
  32'h3e068db8 /* (15, 29, 19) */,
  32'h3dc2b35d /* (11, 29, 19) */,
  32'h3d69f6ae /* (7, 29, 19) */,
  32'h3d2fb3ed /* (3, 29, 19) */,
  32'h3d5c17b6 /* (31, 25, 19) */,
  32'h3d849ae2 /* (27, 25, 19) */,
  32'h3dcf79e9 /* (23, 25, 19) */,
  32'h3e336d1b /* (19, 25, 19) */,
  32'h3e45db44 /* (15, 25, 19) */,
  32'h3e0aca9a /* (11, 25, 19) */,
  32'h3da0c360 /* (7, 25, 19) */,
  32'h3d69f6ae /* (3, 25, 19) */,
  32'h3db58f74 /* (31, 21, 19) */,
  32'h3de04254 /* (27, 21, 19) */,
  32'h3e37494b /* (23, 21, 19) */,
  32'h3ea5d30f /* (19, 21, 19) */,
  32'h3eba8e90 /* (15, 21, 19) */,
  32'h3e7af74d /* (11, 21, 19) */,
  32'h3e0aca9a /* (7, 21, 19) */,
  32'h3dc2b35d /* (3, 21, 19) */,
  32'h3df92d6c /* (31, 17, 19) */,
  32'h3e1d0a10 /* (27, 17, 19) */,
  32'h3e8557f4 /* (23, 17, 19) */,
  32'h3efbd9fe /* (19, 17, 19) */,
  32'h3f1092e5 /* (15, 17, 19) */,
  32'h3eba8e90 /* (11, 17, 19) */,
  32'h3e45db44 /* (7, 17, 19) */,
  32'h3e068db8 /* (3, 17, 19) */,
  32'h3de602d9 /* (31, 13, 19) */,
  32'h3e0f99f2 /* (27, 13, 19) */,
  32'h3e6f82ab /* (23, 13, 19) */,
  32'h3edd8ee5 /* (19, 13, 19) */,
  32'h3efbd9fe /* (15, 13, 19) */,
  32'h3ea5d30f /* (11, 13, 19) */,
  32'h3e336d1b /* (7, 13, 19) */,
  32'h3df79892 /* (3, 13, 19) */,
  32'h3d8ac476 /* (31, 9, 19) */,
  32'h3da95898 /* (27, 9, 19) */,
  32'h3e076ebd /* (23, 9, 19) */,
  32'h3e6f82ab /* (19, 9, 19) */,
  32'h3e8557f4 /* (15, 9, 19) */,
  32'h3e37494b /* (11, 9, 19) */,
  32'h3dcf79e9 /* (7, 9, 19) */,
  32'h3d942dc4 /* (3, 9, 19) */,
  32'h3d398f3f /* (31, 5, 19) */,
  32'h3d5ce99d /* (27, 5, 19) */,
  32'h3da95898 /* (23, 5, 19) */,
  32'h3e0f99f2 /* (19, 5, 19) */,
  32'h3e1d0a10 /* (15, 5, 19) */,
  32'h3de04254 /* (11, 5, 19) */,
  32'h3d849ae2 /* (7, 5, 19) */,
  32'h3d4466f8 /* (3, 5, 19) */,
  32'h3d1e42f1 /* (31, 1, 19) */,
  32'h3d398f3f /* (27, 1, 19) */,
  32'h3d8ac476 /* (23, 1, 19) */,
  32'h3de602d9 /* (19, 1, 19) */,
  32'h3df92d6c /* (15, 1, 19) */,
  32'h3db58f74 /* (11, 1, 19) */,
  32'h3d5c17b6 /* (7, 1, 19) */,
  32'h3d269671 /* (3, 1, 19) */,
  32'h3d202be8 /* (31, 29, 15) */,
  32'h3d424fe8 /* (27, 29, 15) */,
  32'h3d99caa3 /* (23, 29, 15) */,
  32'h3e068db8 /* (19, 29, 15) */,
  32'h3e151f83 /* (15, 29, 15) */,
  32'h3dceffa6 /* (11, 29, 15) */,
  32'h3d6ce397 /* (7, 29, 15) */,
  32'h3d2aacf2 /* (3, 29, 15) */,
  32'h3d5d3ed0 /* (31, 25, 15) */,
  32'h3d880917 /* (27, 25, 15) */,
  32'h3ddc94c6 /* (23, 25, 15) */,
  32'h3e45db44 /* (19, 25, 15) */,
  32'h3e5db918 /* (15, 25, 15) */,
  32'h3e165b49 /* (11, 25, 15) */,
  32'h3da7bf05 /* (7, 25, 15) */,
  32'h3d6ce397 /* (3, 25, 15) */,
  32'h3dc031e4 /* (31, 21, 15) */,
  32'h3df05994 /* (27, 21, 15) */,
  32'h3e49046a /* (23, 21, 15) */,
  32'h3eba8e90 /* (19, 21, 15) */,
  32'h3ed4648a /* (15, 21, 15) */,
  32'h3e8b66c2 /* (11, 21, 15) */,
  32'h3e165b49 /* (7, 21, 15) */,
  32'h3dceffa6 /* (3, 21, 15) */,
  32'h3e09bd27 /* (31, 17, 15) */,
  32'h3e2edbb4 /* (27, 17, 15) */,
  32'h3e969108 /* (23, 17, 15) */,
  32'h3f1092e5 /* (19, 17, 15) */,
  32'h3f275a64 /* (15, 17, 15) */,
  32'h3ed4648a /* (11, 17, 15) */,
  32'h3e5db918 /* (7, 17, 15) */,
  32'h3e151f83 /* (3, 17, 15) */,
  32'h3df92d6c /* (31, 13, 15) */,
  32'h3e1d0a10 /* (27, 13, 15) */,
  32'h3e8557f4 /* (23, 13, 15) */,
  32'h3efbd9fe /* (19, 13, 15) */,
  32'h3f1092e5 /* (15, 13, 15) */,
  32'h3eba8e90 /* (11, 13, 15) */,
  32'h3e45db44 /* (7, 13, 15) */,
  32'h3e068db8 /* (3, 13, 15) */,
  32'h3d8f3655 /* (31, 9, 15) */,
  32'h3db198fc /* (27, 9, 15) */,
  32'h3e123783 /* (23, 9, 15) */,
  32'h3e8557f4 /* (19, 9, 15) */,
  32'h3e969108 /* (15, 9, 15) */,
  32'h3e49046a /* (11, 9, 15) */,
  32'h3ddc94c6 /* (7, 9, 15) */,
  32'h3d99caa3 /* (3, 9, 15) */,
  32'h3d35f880 /* (31, 5, 15) */,
  32'h3d5e11d0 /* (27, 5, 15) */,
  32'h3db198fc /* (23, 5, 15) */,
  32'h3e1d0a10 /* (19, 5, 15) */,
  32'h3e2edbb4 /* (15, 5, 15) */,
  32'h3df05994 /* (11, 5, 15) */,
  32'h3d880917 /* (7, 5, 15) */,
  32'h3d424fe8 /* (3, 5, 15) */,
  32'h3d167d01 /* (31, 1, 15) */,
  32'h3d35f880 /* (27, 1, 15) */,
  32'h3d8f3655 /* (23, 1, 15) */,
  32'h3df92d6c /* (19, 1, 15) */,
  32'h3e09bd27 /* (15, 1, 15) */,
  32'h3dc031e4 /* (11, 1, 15) */,
  32'h3d5d3ed0 /* (7, 1, 15) */,
  32'h3d202be8 /* (3, 1, 15) */,
  32'h3d1a3ccf /* (31, 29, 11) */,
  32'h3d2e4aa1 /* (27, 29, 11) */,
  32'h3d767d5d /* (23, 29, 11) */,
  32'h3dc2b35d /* (19, 29, 11) */,
  32'h3dceffa6 /* (15, 29, 11) */,
  32'h3d9d27e1 /* (11, 29, 11) */,
  32'h3d490aba /* (7, 29, 11) */,
  32'h3d202a91 /* (3, 29, 11) */,
  32'h3d3efe62 /* (31, 25, 11) */,
  32'h3d5ff008 /* (27, 25, 11) */,
  32'h3da777c1 /* (23, 25, 11) */,
  32'h3e0aca9a /* (19, 25, 11) */,
  32'h3e165b49 /* (15, 25, 11) */,
  32'h3ddb1c7f /* (11, 25, 11) */,
  32'h3d84ce75 /* (7, 25, 11) */,
  32'h3d490aba /* (3, 25, 11) */,
  32'h3d9352ec /* (31, 21, 11) */,
  32'h3db345e2 /* (27, 21, 11) */,
  32'h3e0ea5fd /* (23, 21, 11) */,
  32'h3e7af74d /* (19, 21, 11) */,
  32'h3e8b66c2 /* (15, 21, 11) */,
  32'h3e4089a2 /* (11, 21, 11) */,
  32'h3ddb1c7f /* (7, 21, 11) */,
  32'h3d9d27e1 /* (3, 21, 11) */,
  32'h3dc031e4 /* (31, 17, 11) */,
  32'h3df05994 /* (27, 17, 11) */,
  32'h3e49046a /* (23, 17, 11) */,
  32'h3eba8e90 /* (19, 17, 11) */,
  32'h3ed4648a /* (15, 17, 11) */,
  32'h3e8b66c2 /* (11, 17, 11) */,
  32'h3e165b49 /* (7, 17, 11) */,
  32'h3dceffa6 /* (3, 17, 11) */,
  32'h3db58f74 /* (31, 13, 11) */,
  32'h3de04254 /* (27, 13, 11) */,
  32'h3e37494b /* (23, 13, 11) */,
  32'h3ea5d30f /* (19, 13, 11) */,
  32'h3eba8e90 /* (15, 13, 11) */,
  32'h3e7af74d /* (11, 13, 11) */,
  32'h3e0aca9a /* (7, 13, 11) */,
  32'h3dc2b35d /* (3, 13, 11) */,
  32'h3d68852c /* (31, 9, 11) */,
  32'h3d8b02ad /* (27, 9, 11) */,
  32'h3dd6aa1b /* (23, 9, 11) */,
  32'h3e37494b /* (19, 9, 11) */,
  32'h3e49046a /* (15, 9, 11) */,
  32'h3e0ea5fd /* (11, 9, 11) */,
  32'h3da777c1 /* (7, 9, 11) */,
  32'h3d767d5d /* (3, 9, 11) */,
  32'h3d26c9db /* (31, 5, 11) */,
  32'h3d3fb488 /* (27, 5, 11) */,
  32'h3d8b02ad /* (23, 5, 11) */,
  32'h3de04254 /* (19, 5, 11) */,
  32'h3df05994 /* (15, 5, 11) */,
  32'h3db345e2 /* (11, 5, 11) */,
  32'h3d5ff008 /* (7, 5, 11) */,
  32'h3d2e4aa1 /* (3, 5, 11) */,
  32'h3d151591 /* (31, 1, 11) */,
  32'h3d26c9db /* (27, 1, 11) */,
  32'h3d68852c /* (23, 1, 11) */,
  32'h3db58f74 /* (19, 1, 11) */,
  32'h3dc031e4 /* (15, 1, 11) */,
  32'h3d9352ec /* (11, 1, 11) */,
  32'h3d3efe62 /* (7, 1, 11) */,
  32'h3d1a3ccf /* (3, 1, 11) */,
  32'h3d1c3652 /* (31, 29, 7) */,
  32'h3d147808 /* (27, 29, 7) */,
  32'h3d2aad03 /* (23, 29, 7) */,
  32'h3d69f6ae /* (19, 29, 7) */,
  32'h3d6ce397 /* (15, 29, 7) */,
  32'h3d490aba /* (11, 29, 7) */,
  32'h3d1969a9 /* (7, 29, 7) */,
  32'h3d179239 /* (3, 29, 7) */,
  32'h3d167b79 /* (31, 25, 7) */,
  32'h3d21f168 /* (27, 25, 7) */,
  32'h3d563bcb /* (23, 25, 7) */,
  32'h3da0c360 /* (19, 25, 7) */,
  32'h3da7bf05 /* (15, 25, 7) */,
  32'h3d84ce75 /* (11, 25, 7) */,
  32'h3d348078 /* (7, 25, 7) */,
  32'h3d1969a9 /* (3, 25, 7) */,
  32'h3d3efe62 /* (31, 21, 7) */,
  32'h3d5ff008 /* (27, 21, 7) */,
  32'h3da777c1 /* (23, 21, 7) */,
  32'h3e0aca9a /* (19, 21, 7) */,
  32'h3e165b49 /* (15, 21, 7) */,
  32'h3ddb1c7f /* (11, 21, 7) */,
  32'h3d84ce75 /* (7, 21, 7) */,
  32'h3d490aba /* (3, 21, 7) */,
  32'h3d5d3ed0 /* (31, 17, 7) */,
  32'h3d880917 /* (27, 17, 7) */,
  32'h3ddc94c6 /* (23, 17, 7) */,
  32'h3e45db44 /* (19, 17, 7) */,
  32'h3e5db918 /* (15, 17, 7) */,
  32'h3e165b49 /* (11, 17, 7) */,
  32'h3da7bf05 /* (7, 17, 7) */,
  32'h3d6ce397 /* (3, 17, 7) */,
  32'h3d5c17b6 /* (31, 13, 7) */,
  32'h3d849ae2 /* (27, 13, 7) */,
  32'h3dcf79e9 /* (23, 13, 7) */,
  32'h3e336d1b /* (19, 13, 7) */,
  32'h3e45db44 /* (15, 13, 7) */,
  32'h3e0aca9a /* (11, 13, 7) */,
  32'h3da0c360 /* (7, 13, 7) */,
  32'h3d69f6ae /* (3, 13, 7) */,
  32'h3d245baa /* (31, 9, 7) */,
  32'h3d39ba58 /* (27, 9, 7) */,
  32'h3d8354ed /* (23, 9, 7) */,
  32'h3dcf79e9 /* (19, 9, 7) */,
  32'h3ddc94c6 /* (15, 9, 7) */,
  32'h3da777c1 /* (11, 9, 7) */,
  32'h3d563bcb /* (7, 9, 7) */,
  32'h3d2aad03 /* (3, 9, 7) */,
  32'h3d151e01 /* (31, 5, 7) */,
  32'h3d170afd /* (27, 5, 7) */,
  32'h3d39ba58 /* (23, 5, 7) */,
  32'h3d849ae2 /* (19, 5, 7) */,
  32'h3d880917 /* (15, 5, 7) */,
  32'h3d5ff008 /* (11, 5, 7) */,
  32'h3d21f168 /* (7, 5, 7) */,
  32'h3d147808 /* (3, 5, 7) */,
  32'h3d2402bf /* (31, 1, 7) */,
  32'h3d151e01 /* (27, 1, 7) */,
  32'h3d245baa /* (23, 1, 7) */,
  32'h3d5c17b6 /* (19, 1, 7) */,
  32'h3d5d3ed0 /* (15, 1, 7) */,
  32'h3d3efe62 /* (11, 1, 7) */,
  32'h3d167b79 /* (7, 1, 7) */,
  32'h3d1c3652 /* (3, 1, 7) */,
  32'h3d960c3c /* (31, 29, 3) */,
  32'h3d314afb /* (27, 29, 3) */,
  32'h3d144047 /* (23, 29, 3) */,
  32'h3d2fb3ed /* (19, 29, 3) */,
  32'h3d2aacf2 /* (15, 29, 3) */,
  32'h3d202a91 /* (11, 29, 3) */,
  32'h3d179239 /* (7, 29, 3) */,
  32'h3d68b01f /* (3, 29, 3) */,
  32'h3d1c3652 /* (31, 25, 3) */,
  32'h3d147808 /* (27, 25, 3) */,
  32'h3d2aad03 /* (23, 25, 3) */,
  32'h3d69f6ae /* (19, 25, 3) */,
  32'h3d6ce397 /* (15, 25, 3) */,
  32'h3d490aba /* (11, 25, 3) */,
  32'h3d1969a9 /* (7, 25, 3) */,
  32'h3d179239 /* (3, 25, 3) */,
  32'h3d1a3ccf /* (31, 21, 3) */,
  32'h3d2e4aa1 /* (27, 21, 3) */,
  32'h3d767d5d /* (23, 21, 3) */,
  32'h3dc2b35d /* (19, 21, 3) */,
  32'h3dceffa6 /* (15, 21, 3) */,
  32'h3d9d27e1 /* (11, 21, 3) */,
  32'h3d490aba /* (7, 21, 3) */,
  32'h3d202a91 /* (3, 21, 3) */,
  32'h3d202be8 /* (31, 17, 3) */,
  32'h3d424fe8 /* (27, 17, 3) */,
  32'h3d99caa3 /* (23, 17, 3) */,
  32'h3e068db8 /* (19, 17, 3) */,
  32'h3e151f83 /* (15, 17, 3) */,
  32'h3dceffa6 /* (11, 17, 3) */,
  32'h3d6ce397 /* (7, 17, 3) */,
  32'h3d2aacf2 /* (3, 17, 3) */,
  32'h3d269671 /* (31, 13, 3) */,
  32'h3d4466f8 /* (27, 13, 3) */,
  32'h3d942dc4 /* (23, 13, 3) */,
  32'h3df79892 /* (19, 13, 3) */,
  32'h3e068db8 /* (15, 13, 3) */,
  32'h3dc2b35d /* (11, 13, 3) */,
  32'h3d69f6ae /* (7, 13, 3) */,
  32'h3d2fb3ed /* (3, 13, 3) */,
  32'h3d126006 /* (31, 9, 3) */,
  32'h3d1addce /* (27, 9, 3) */,
  32'h3d48821f /* (23, 9, 3) */,
  32'h3d942dc4 /* (19, 9, 3) */,
  32'h3d99caa3 /* (15, 9, 3) */,
  32'h3d767d5d /* (11, 9, 3) */,
  32'h3d2aad03 /* (7, 9, 3) */,
  32'h3d144047 /* (3, 9, 3) */,
  32'h3d45ae9a /* (31, 5, 3) */,
  32'h3d1ccb4c /* (27, 5, 3) */,
  32'h3d1addce /* (23, 5, 3) */,
  32'h3d4466f8 /* (19, 5, 3) */,
  32'h3d424fe8 /* (15, 5, 3) */,
  32'h3d2e4aa1 /* (11, 5, 3) */,
  32'h3d147808 /* (7, 5, 3) */,
  32'h3d314afb /* (3, 5, 3) */,
  32'h3deb372d /* (31, 1, 3) */,
  32'h3d45ae9a /* (27, 1, 3) */,
  32'h3d126006 /* (23, 1, 3) */,
  32'h3d269671 /* (19, 1, 3) */,
  32'h3d202be8 /* (15, 1, 3) */,
  32'h3d1a3ccf /* (11, 1, 3) */,
  32'h3d1c3652 /* (7, 1, 3) */,
  32'h3d960c3c /* (3, 1, 3) */,
  32'h3dbfa8df /* (30, 29, 31) */,
  32'h3d2ba889 /* (26, 29, 31) */,
  32'h3d14c0fd /* (22, 29, 31) */,
  32'h3d276174 /* (18, 29, 31) */,
  32'h3d276174 /* (14, 29, 31) */,
  32'h3d14c0fd /* (10, 29, 31) */,
  32'h3d2ba889 /* (6, 29, 31) */,
  32'h3dbfa8df /* (2, 29, 31) */,
  32'h3d20a35e /* (30, 25, 31) */,
  32'h3d146a43 /* (26, 25, 31) */,
  32'h3d305430 /* (22, 25, 31) */,
  32'h3d62906c /* (18, 25, 31) */,
  32'h3d62906c /* (14, 25, 31) */,
  32'h3d305430 /* (10, 25, 31) */,
  32'h3d146a43 /* (6, 25, 31) */,
  32'h3d20a35e /* (2, 25, 31) */,
  32'h3d16ed42 /* (30, 21, 31) */,
  32'h3d31191b /* (26, 21, 31) */,
  32'h3d829849 /* (22, 21, 31) */,
  32'h3dc01db4 /* (18, 21, 31) */,
  32'h3dc01db4 /* (14, 21, 31) */,
  32'h3d829849 /* (10, 21, 31) */,
  32'h3d31191b /* (6, 21, 31) */,
  32'h3d16ed42 /* (2, 21, 31) */,
  32'h3d1a0745 /* (30, 17, 31) */,
  32'h3d46f53f /* (26, 17, 31) */,
  32'h3da5ac70 /* (22, 17, 31) */,
  32'h3e06d8bb /* (18, 17, 31) */,
  32'h3e06d8bb /* (14, 17, 31) */,
  32'h3da5ac70 /* (10, 17, 31) */,
  32'h3d46f53f /* (6, 17, 31) */,
  32'h3d1a0745 /* (2, 17, 31) */,
  32'h3d214ba3 /* (30, 13, 31) */,
  32'h3d4876ff /* (26, 13, 31) */,
  32'h3d9e7894 /* (22, 13, 31) */,
  32'h3df65860 /* (18, 13, 31) */,
  32'h3df65860 /* (14, 13, 31) */,
  32'h3d9e7894 /* (10, 13, 31) */,
  32'h3d4876ff /* (6, 13, 31) */,
  32'h3d214ba3 /* (2, 13, 31) */,
  32'h3d11c69f /* (30, 9, 31) */,
  32'h3d1c53e8 /* (26, 9, 31) */,
  32'h3d52081f /* (22, 9, 31) */,
  32'h3d90dff9 /* (18, 9, 31) */,
  32'h3d90dff9 /* (14, 9, 31) */,
  32'h3d52081f /* (10, 9, 31) */,
  32'h3d1c53e8 /* (6, 9, 31) */,
  32'h3d11c69f /* (2, 9, 31) */,
  32'h3d59109a /* (30, 5, 31) */,
  32'h3d1a8b5a /* (26, 5, 31) */,
  32'h3d1d9589 /* (22, 5, 31) */,
  32'h3d3c7841 /* (18, 5, 31) */,
  32'h3d3c7841 /* (14, 5, 31) */,
  32'h3d1d9589 /* (10, 5, 31) */,
  32'h3d1a8b5a /* (6, 5, 31) */,
  32'h3d59109a /* (2, 5, 31) */,
  32'h3e4aeee2 /* (30, 1, 31) */,
  32'h3d3c9698 /* (26, 1, 31) */,
  32'h3d119771 /* (22, 1, 31) */,
  32'h3d1e0bb6 /* (18, 1, 31) */,
  32'h3d1e0bb6 /* (14, 1, 31) */,
  32'h3d119771 /* (10, 1, 31) */,
  32'h3d3c9698 /* (6, 1, 31) */,
  32'h3e4aeee2 /* (2, 1, 31) */,
  32'h3d3cd255 /* (30, 29, 27) */,
  32'h3d16d305 /* (26, 29, 27) */,
  32'h3d2344c4 /* (22, 29, 27) */,
  32'h3d487174 /* (18, 29, 27) */,
  32'h3d487174 /* (14, 29, 27) */,
  32'h3d2344c4 /* (10, 29, 27) */,
  32'h3d16d305 /* (6, 29, 27) */,
  32'h3d3cd255 /* (2, 29, 27) */,
  32'h3d14b1c0 /* (30, 25, 27) */,
  32'h3d1b2471 /* (26, 25, 27) */,
  32'h3d4b3dc7 /* (22, 25, 27) */,
  32'h3d8a0000 /* (18, 25, 27) */,
  32'h3d8a0000 /* (14, 25, 27) */,
  32'h3d4b3dc7 /* (10, 25, 27) */,
  32'h3d1b2471 /* (6, 25, 27) */,
  32'h3d14b1c0 /* (2, 25, 27) */,
  32'h3d29823f /* (30, 21, 27) */,
  32'h3d4d9045 /* (26, 21, 27) */,
  32'h3d9d9380 /* (22, 21, 27) */,
  32'h3deed79f /* (18, 21, 27) */,
  32'h3deed79f /* (14, 21, 27) */,
  32'h3d9d9380 /* (10, 21, 27) */,
  32'h3d4d9045 /* (6, 21, 27) */,
  32'h3d29823f /* (2, 21, 27) */,
  32'h3d3a7be5 /* (30, 17, 27) */,
  32'h3d73b16f /* (26, 17, 27) */,
  32'h3dce52e6 /* (22, 17, 27) */,
  32'h3e2a981c /* (18, 17, 27) */,
  32'h3e2a981c /* (14, 17, 27) */,
  32'h3dce52e6 /* (10, 17, 27) */,
  32'h3d73b16f /* (6, 17, 27) */,
  32'h3d3a7be5 /* (2, 17, 27) */,
  32'h3d3d84de /* (30, 13, 27) */,
  32'h3d700ffa /* (26, 13, 27) */,
  32'h3dc29629 /* (22, 13, 27) */,
  32'h3e1a8d8c /* (18, 13, 27) */,
  32'h3e1a8d8c /* (14, 13, 27) */,
  32'h3dc29629 /* (10, 13, 27) */,
  32'h3d700ffa /* (6, 13, 27) */,
  32'h3d3d84de /* (2, 13, 27) */,
  32'h3d18622e /* (30, 9, 27) */,
  32'h3d2db0cc /* (26, 9, 27) */,
  32'h3d781ae6 /* (22, 9, 27) */,
  32'h3db24f8e /* (18, 9, 27) */,
  32'h3db24f8e /* (14, 9, 27) */,
  32'h3d781ae6 /* (10, 9, 27) */,
  32'h3d2db0cc /* (6, 9, 27) */,
  32'h3d18622e /* (2, 9, 27) */,
  32'h3d213c91 /* (30, 5, 27) */,
  32'h3d14f7ce /* (26, 5, 27) */,
  32'h3d30fc5a /* (22, 5, 27) */,
  32'h3d63687e /* (18, 5, 27) */,
  32'h3d63687e /* (14, 5, 27) */,
  32'h3d30fc5a /* (10, 5, 27) */,
  32'h3d14f7ce /* (6, 5, 27) */,
  32'h3d213c91 /* (2, 5, 27) */,
  32'h3d59109a /* (30, 1, 27) */,
  32'h3d1a8b5a /* (26, 1, 27) */,
  32'h3d1d9589 /* (22, 1, 27) */,
  32'h3d3c7841 /* (18, 1, 27) */,
  32'h3d3c7841 /* (14, 1, 27) */,
  32'h3d1d9589 /* (10, 1, 27) */,
  32'h3d1a8b5a /* (6, 1, 27) */,
  32'h3d59109a /* (2, 1, 27) */,
  32'h3d12f42a /* (30, 29, 23) */,
  32'h3d215063 /* (26, 29, 23) */,
  32'h3d5dae2c /* (22, 29, 23) */,
  32'h3d9b2a7b /* (18, 29, 23) */,
  32'h3d9b2a7b /* (14, 29, 23) */,
  32'h3d5dae2c /* (10, 29, 23) */,
  32'h3d215063 /* (6, 29, 23) */,
  32'h3d12f42a /* (2, 29, 23) */,
  32'h3d26a1b5 /* (30, 25, 23) */,
  32'h3d45eb5b /* (26, 25, 23) */,
  32'h3d94014f /* (22, 25, 23) */,
  32'h3ddc09d8 /* (18, 25, 23) */,
  32'h3ddc09d8 /* (14, 25, 23) */,
  32'h3d94014f /* (10, 25, 23) */,
  32'h3d45eb5b /* (6, 25, 23) */,
  32'h3d26a1b5 /* (2, 25, 23) */,
  32'h3d6d9fa3 /* (30, 21, 23) */,
  32'h3d9750ce /* (26, 21, 23) */,
  32'h3df71c69 /* (22, 21, 23) */,
  32'h3e458f30 /* (18, 21, 23) */,
  32'h3e458f30 /* (14, 21, 23) */,
  32'h3df71c69 /* (10, 21, 23) */,
  32'h3d9750ce /* (6, 21, 23) */,
  32'h3d6d9fa3 /* (2, 21, 23) */,
  32'h3d9314c2 /* (30, 17, 23) */,
  32'h3dc42ad0 /* (26, 17, 23) */,
  32'h3e2b3653 /* (22, 17, 23) */,
  32'h3e91e4f8 /* (18, 17, 23) */,
  32'h3e91e4f8 /* (14, 17, 23) */,
  32'h3e2b3653 /* (10, 17, 23) */,
  32'h3dc42ad0 /* (6, 17, 23) */,
  32'h3d9314c2 /* (2, 17, 23) */,
  32'h3d8e358b /* (30, 13, 23) */,
  32'h3db9d5f4 /* (26, 13, 23) */,
  32'h3e1d56b2 /* (22, 13, 23) */,
  32'h3e821787 /* (18, 13, 23) */,
  32'h3e821787 /* (14, 13, 23) */,
  32'h3e1d56b2 /* (10, 13, 23) */,
  32'h3db9d5f4 /* (6, 13, 23) */,
  32'h3d8e358b /* (2, 13, 23) */,
  32'h3d42665b /* (30, 9, 23) */,
  32'h3d6fd024 /* (26, 9, 23) */,
  32'h3dbbc730 /* (22, 9, 23) */,
  32'h3e10cac5 /* (18, 9, 23) */,
  32'h3e10cac5 /* (14, 9, 23) */,
  32'h3dbbc730 /* (10, 9, 23) */,
  32'h3d6fd024 /* (6, 9, 23) */,
  32'h3d42665b /* (2, 9, 23) */,
  32'h3d18622e /* (30, 5, 23) */,
  32'h3d2db0cc /* (26, 5, 23) */,
  32'h3d781ae6 /* (22, 5, 23) */,
  32'h3db24f8e /* (18, 5, 23) */,
  32'h3db24f8e /* (14, 5, 23) */,
  32'h3d781ae6 /* (10, 5, 23) */,
  32'h3d2db0cc /* (6, 5, 23) */,
  32'h3d18622e /* (2, 5, 23) */,
  32'h3d11c69f /* (30, 1, 23) */,
  32'h3d1c53e8 /* (26, 1, 23) */,
  32'h3d52081f /* (22, 1, 23) */,
  32'h3d90dff9 /* (18, 1, 23) */,
  32'h3d90dff9 /* (14, 1, 23) */,
  32'h3d52081f /* (10, 1, 23) */,
  32'h3d1c53e8 /* (6, 1, 23) */,
  32'h3d11c69f /* (2, 1, 23) */,
  32'h3d29e985 /* (30, 29, 19) */,
  32'h3d54a03b /* (26, 29, 19) */,
  32'h3da99659 /* (22, 29, 19) */,
  32'h3e04d0b8 /* (18, 29, 19) */,
  32'h3e04d0b8 /* (14, 29, 19) */,
  32'h3da99659 /* (10, 29, 19) */,
  32'h3d54a03b /* (6, 29, 19) */,
  32'h3d29e985 /* (2, 29, 19) */,
  32'h3d6129ae /* (30, 25, 19) */,
  32'h3d90c8a7 /* (26, 25, 19) */,
  32'h3defa49b /* (22, 25, 19) */,
  32'h3e41f14c /* (18, 25, 19) */,
  32'h3e41f14c /* (14, 25, 19) */,
  32'h3defa49b /* (10, 25, 19) */,
  32'h3d90c8a7 /* (6, 25, 19) */,
  32'h3d6129ae /* (2, 25, 19) */,
  32'h3dba5db4 /* (30, 21, 19) */,
  32'h3df74dbc /* (26, 21, 19) */,
  32'h3e562fb1 /* (22, 21, 19) */,
  32'h3eb517ce /* (18, 21, 19) */,
  32'h3eb517ce /* (14, 21, 19) */,
  32'h3e562fb1 /* (10, 21, 19) */,
  32'h3df74dbc /* (6, 21, 19) */,
  32'h3dba5db4 /* (2, 21, 19) */,
  32'h3e003b1e /* (30, 17, 19) */,
  32'h3e2ea39a /* (26, 17, 19) */,
  32'h3e9d80fb /* (22, 17, 19) */,
  32'h3f0af24f /* (18, 17, 19) */,
  32'h3f0af24f /* (14, 17, 19) */,
  32'h3e9d80fb /* (10, 17, 19) */,
  32'h3e2ea39a /* (6, 17, 19) */,
  32'h3e003b1e /* (2, 17, 19) */,
  32'h3dec70da /* (30, 13, 19) */,
  32'h3e1f113d /* (26, 13, 19) */,
  32'h3e8cbae1 /* (22, 13, 19) */,
  32'h3ef33ce4 /* (18, 13, 19) */,
  32'h3ef33ce4 /* (14, 13, 19) */,
  32'h3e8cbae1 /* (10, 13, 19) */,
  32'h3e1f113d /* (6, 13, 19) */,
  32'h3dec70da /* (2, 13, 19) */,
  32'h3d8e358b /* (30, 9, 19) */,
  32'h3db9d5f4 /* (26, 9, 19) */,
  32'h3e1d56b2 /* (22, 9, 19) */,
  32'h3e821787 /* (18, 9, 19) */,
  32'h3e821787 /* (14, 9, 19) */,
  32'h3e1d56b2 /* (10, 9, 19) */,
  32'h3db9d5f4 /* (6, 9, 19) */,
  32'h3d8e358b /* (2, 9, 19) */,
  32'h3d3d84de /* (30, 5, 19) */,
  32'h3d700ffa /* (26, 5, 19) */,
  32'h3dc29629 /* (22, 5, 19) */,
  32'h3e1a8d8c /* (18, 5, 19) */,
  32'h3e1a8d8c /* (14, 5, 19) */,
  32'h3dc29629 /* (10, 5, 19) */,
  32'h3d700ffa /* (6, 5, 19) */,
  32'h3d3d84de /* (2, 5, 19) */,
  32'h3d214ba3 /* (30, 1, 19) */,
  32'h3d4876ff /* (26, 1, 19) */,
  32'h3d9e7894 /* (22, 1, 19) */,
  32'h3df65860 /* (18, 1, 19) */,
  32'h3df65860 /* (14, 1, 19) */,
  32'h3d9e7894 /* (10, 1, 19) */,
  32'h3d4876ff /* (6, 1, 19) */,
  32'h3d214ba3 /* (2, 1, 19) */,
  32'h3d240321 /* (30, 29, 15) */,
  32'h3d54ba37 /* (26, 29, 15) */,
  32'h3db22d06 /* (22, 29, 15) */,
  32'h3e11d12f /* (18, 29, 15) */,
  32'h3e11d12f /* (14, 29, 15) */,
  32'h3db22d06 /* (10, 29, 15) */,
  32'h3d54ba37 /* (6, 29, 15) */,
  32'h3d240321 /* (2, 29, 15) */,
  32'h3d62f778 /* (30, 25, 15) */,
  32'h3d95be73 /* (26, 25, 15) */,
  32'h3e009a19 /* (22, 25, 15) */,
  32'h3e57a44b /* (18, 25, 15) */,
  32'h3e57a44b /* (14, 25, 15) */,
  32'h3e009a19 /* (10, 25, 15) */,
  32'h3d95be73 /* (6, 25, 15) */,
  32'h3d62f778 /* (2, 25, 15) */,
  32'h3dc59b81 /* (30, 21, 15) */,
  32'h3e0533d0 /* (26, 21, 15) */,
  32'h3e6c6ac0 /* (22, 21, 15) */,
  32'h3eccf8ff /* (18, 21, 15) */,
  32'h3eccf8ff /* (14, 21, 15) */,
  32'h3e6c6ac0 /* (10, 21, 15) */,
  32'h3e0533d0 /* (6, 21, 15) */,
  32'h3dc59b81 /* (2, 21, 15) */,
  32'h3e0de5f8 /* (30, 17, 15) */,
  32'h3e430b11 /* (26, 17, 15) */,
  32'h3eb2925b /* (22, 17, 15) */,
  32'h3f202f9a /* (18, 17, 15) */,
  32'h3f202f9a /* (14, 17, 15) */,
  32'h3eb2925b /* (10, 17, 15) */,
  32'h3e430b11 /* (6, 17, 15) */,
  32'h3e0de5f8 /* (2, 17, 15) */,
  32'h3e003b1e /* (30, 13, 15) */,
  32'h3e2ea39a /* (26, 13, 15) */,
  32'h3e9d80fb /* (22, 13, 15) */,
  32'h3f0af24f /* (18, 13, 15) */,
  32'h3f0af24f /* (14, 13, 15) */,
  32'h3e9d80fb /* (10, 13, 15) */,
  32'h3e2ea39a /* (6, 13, 15) */,
  32'h3e003b1e /* (2, 13, 15) */,
  32'h3d9314c2 /* (30, 9, 15) */,
  32'h3dc42ad0 /* (26, 9, 15) */,
  32'h3e2b3653 /* (22, 9, 15) */,
  32'h3e91e4f8 /* (18, 9, 15) */,
  32'h3e91e4f8 /* (14, 9, 15) */,
  32'h3e2b3653 /* (10, 9, 15) */,
  32'h3dc42ad0 /* (6, 9, 15) */,
  32'h3d9314c2 /* (2, 9, 15) */,
  32'h3d3a7be5 /* (30, 5, 15) */,
  32'h3d73b16f /* (26, 5, 15) */,
  32'h3dce52e6 /* (22, 5, 15) */,
  32'h3e2a981c /* (18, 5, 15) */,
  32'h3e2a981c /* (14, 5, 15) */,
  32'h3dce52e6 /* (10, 5, 15) */,
  32'h3d73b16f /* (6, 5, 15) */,
  32'h3d3a7be5 /* (2, 5, 15) */,
  32'h3d1a0745 /* (30, 1, 15) */,
  32'h3d46f53f /* (26, 1, 15) */,
  32'h3da5ac70 /* (22, 1, 15) */,
  32'h3e06d8bb /* (18, 1, 15) */,
  32'h3e06d8bb /* (14, 1, 15) */,
  32'h3da5ac70 /* (10, 1, 15) */,
  32'h3d46f53f /* (6, 1, 15) */,
  32'h3d1a0745 /* (2, 1, 15) */,
  32'h3d1c5f03 /* (30, 29, 11) */,
  32'h3d39bb76 /* (26, 29, 11) */,
  32'h3d8ae43c /* (22, 29, 11) */,
  32'h3dce7d45 /* (18, 29, 11) */,
  32'h3dce7d45 /* (14, 29, 11) */,
  32'h3d8ae43c /* (10, 29, 11) */,
  32'h3d39bb76 /* (6, 29, 11) */,
  32'h3d1c5f03 /* (2, 29, 11) */,
  32'h3d42a7b8 /* (30, 25, 11) */,
  32'h3d71ecf9 /* (26, 25, 11) */,
  32'h3dbf3f1d /* (22, 25, 11) */,
  32'h3e14a5c9 /* (18, 25, 11) */,
  32'h3e14a5c9 /* (14, 25, 11) */,
  32'h3dbf3f1d /* (10, 25, 11) */,
  32'h3d71ecf9 /* (6, 25, 11) */,
  32'h3d42a7b8 /* (2, 25, 11) */,
  32'h3d96eb50 /* (30, 21, 11) */,
  32'h3dc480ba /* (26, 21, 11) */,
  32'h3e257fc6 /* (22, 21, 11) */,
  32'h3e882756 /* (18, 21, 11) */,
  32'h3e882756 /* (14, 21, 11) */,
  32'h3e257fc6 /* (10, 21, 11) */,
  32'h3dc480ba /* (6, 21, 11) */,
  32'h3d96eb50 /* (2, 21, 11) */,
  32'h3dc59b81 /* (30, 17, 11) */,
  32'h3e0533d0 /* (26, 17, 11) */,
  32'h3e6c6ac0 /* (22, 17, 11) */,
  32'h3eccf8ff /* (18, 17, 11) */,
  32'h3eccf8ff /* (14, 17, 11) */,
  32'h3e6c6ac0 /* (10, 17, 11) */,
  32'h3e0533d0 /* (6, 17, 11) */,
  32'h3dc59b81 /* (2, 17, 11) */,
  32'h3dba5db4 /* (30, 13, 11) */,
  32'h3df74dbc /* (26, 13, 11) */,
  32'h3e562fb1 /* (22, 13, 11) */,
  32'h3eb517ce /* (18, 13, 11) */,
  32'h3eb517ce /* (14, 13, 11) */,
  32'h3e562fb1 /* (10, 13, 11) */,
  32'h3df74dbc /* (6, 13, 11) */,
  32'h3dba5db4 /* (2, 13, 11) */,
  32'h3d6d9fa3 /* (30, 9, 11) */,
  32'h3d9750ce /* (26, 9, 11) */,
  32'h3df71c69 /* (22, 9, 11) */,
  32'h3e458f30 /* (18, 9, 11) */,
  32'h3e458f30 /* (14, 9, 11) */,
  32'h3df71c69 /* (10, 9, 11) */,
  32'h3d9750ce /* (6, 9, 11) */,
  32'h3d6d9fa3 /* (2, 9, 11) */,
  32'h3d29823f /* (30, 5, 11) */,
  32'h3d4d9045 /* (26, 5, 11) */,
  32'h3d9d9380 /* (22, 5, 11) */,
  32'h3deed79f /* (18, 5, 11) */,
  32'h3deed79f /* (14, 5, 11) */,
  32'h3d9d9380 /* (10, 5, 11) */,
  32'h3d4d9045 /* (6, 5, 11) */,
  32'h3d29823f /* (2, 5, 11) */,
  32'h3d16ed42 /* (30, 1, 11) */,
  32'h3d31191b /* (26, 1, 11) */,
  32'h3d829849 /* (22, 1, 11) */,
  32'h3dc01db4 /* (18, 1, 11) */,
  32'h3dc01db4 /* (14, 1, 11) */,
  32'h3d829849 /* (10, 1, 11) */,
  32'h3d31191b /* (6, 1, 11) */,
  32'h3d16ed42 /* (2, 1, 11) */,
  32'h3d1a2949 /* (30, 29, 7) */,
  32'h3d159d44 /* (26, 29, 7) */,
  32'h3d387393 /* (22, 29, 7) */,
  32'h3d71c736 /* (18, 29, 7) */,
  32'h3d71c736 /* (14, 29, 7) */,
  32'h3d387393 /* (10, 29, 7) */,
  32'h3d159d44 /* (6, 29, 7) */,
  32'h3d1a2949 /* (2, 29, 7) */,
  32'h3d1777c7 /* (30, 25, 7) */,
  32'h3d29a602 /* (26, 25, 7) */,
  32'h3d6deb12 /* (22, 25, 7) */,
  32'h3da8d240 /* (18, 25, 7) */,
  32'h3da8d240 /* (14, 25, 7) */,
  32'h3d6deb12 /* (10, 25, 7) */,
  32'h3d29a602 /* (6, 25, 7) */,
  32'h3d1777c7 /* (2, 25, 7) */,
  32'h3d42a7b8 /* (30, 21, 7) */,
  32'h3d71ecf9 /* (26, 21, 7) */,
  32'h3dbf3f1d /* (22, 21, 7) */,
  32'h3e14a5c9 /* (18, 21, 7) */,
  32'h3e14a5c9 /* (14, 21, 7) */,
  32'h3dbf3f1d /* (10, 21, 7) */,
  32'h3d71ecf9 /* (6, 21, 7) */,
  32'h3d42a7b8 /* (2, 21, 7) */,
  32'h3d62f778 /* (30, 17, 7) */,
  32'h3d95be73 /* (26, 17, 7) */,
  32'h3e009a19 /* (22, 17, 7) */,
  32'h3e57a44b /* (18, 17, 7) */,
  32'h3e57a44b /* (14, 17, 7) */,
  32'h3e009a19 /* (10, 17, 7) */,
  32'h3d95be73 /* (6, 17, 7) */,
  32'h3d62f778 /* (2, 17, 7) */,
  32'h3d6129ae /* (30, 13, 7) */,
  32'h3d90c8a7 /* (26, 13, 7) */,
  32'h3defa49b /* (22, 13, 7) */,
  32'h3e41f14c /* (18, 13, 7) */,
  32'h3e41f14c /* (14, 13, 7) */,
  32'h3defa49b /* (10, 13, 7) */,
  32'h3d90c8a7 /* (6, 13, 7) */,
  32'h3d6129ae /* (2, 13, 7) */,
  32'h3d26a1b5 /* (30, 9, 7) */,
  32'h3d45eb5b /* (26, 9, 7) */,
  32'h3d94014f /* (22, 9, 7) */,
  32'h3ddc09d8 /* (18, 9, 7) */,
  32'h3ddc09d8 /* (14, 9, 7) */,
  32'h3d94014f /* (10, 9, 7) */,
  32'h3d45eb5b /* (6, 9, 7) */,
  32'h3d26a1b5 /* (2, 9, 7) */,
  32'h3d14b1c0 /* (30, 5, 7) */,
  32'h3d1b2471 /* (26, 5, 7) */,
  32'h3d4b3dc7 /* (22, 5, 7) */,
  32'h3d8a0000 /* (18, 5, 7) */,
  32'h3d8a0000 /* (14, 5, 7) */,
  32'h3d4b3dc7 /* (10, 5, 7) */,
  32'h3d1b2471 /* (6, 5, 7) */,
  32'h3d14b1c0 /* (2, 5, 7) */,
  32'h3d20a35e /* (30, 1, 7) */,
  32'h3d146a43 /* (26, 1, 7) */,
  32'h3d305430 /* (22, 1, 7) */,
  32'h3d62906c /* (18, 1, 7) */,
  32'h3d62906c /* (14, 1, 7) */,
  32'h3d305430 /* (10, 1, 7) */,
  32'h3d146a43 /* (6, 1, 7) */,
  32'h3d20a35e /* (2, 1, 7) */,
  32'h3d866355 /* (30, 29, 3) */,
  32'h3d211f1b /* (26, 29, 3) */,
  32'h3d18cb02 /* (22, 29, 3) */,
  32'h3d3188e3 /* (18, 29, 3) */,
  32'h3d3188e3 /* (14, 29, 3) */,
  32'h3d18cb02 /* (10, 29, 3) */,
  32'h3d211f1b /* (6, 29, 3) */,
  32'h3d866355 /* (2, 29, 3) */,
  32'h3d1a2949 /* (30, 25, 3) */,
  32'h3d159d44 /* (26, 25, 3) */,
  32'h3d387393 /* (22, 25, 3) */,
  32'h3d71c736 /* (18, 25, 3) */,
  32'h3d71c736 /* (14, 25, 3) */,
  32'h3d387393 /* (10, 25, 3) */,
  32'h3d159d44 /* (6, 25, 3) */,
  32'h3d1a2949 /* (2, 25, 3) */,
  32'h3d1c5f03 /* (30, 21, 3) */,
  32'h3d39bb76 /* (26, 21, 3) */,
  32'h3d8ae43c /* (22, 21, 3) */,
  32'h3dce7d45 /* (18, 21, 3) */,
  32'h3dce7d45 /* (14, 21, 3) */,
  32'h3d8ae43c /* (10, 21, 3) */,
  32'h3d39bb76 /* (6, 21, 3) */,
  32'h3d1c5f03 /* (2, 21, 3) */,
  32'h3d240321 /* (30, 17, 3) */,
  32'h3d54ba37 /* (26, 17, 3) */,
  32'h3db22d06 /* (22, 17, 3) */,
  32'h3e11d12f /* (18, 17, 3) */,
  32'h3e11d12f /* (14, 17, 3) */,
  32'h3db22d06 /* (10, 17, 3) */,
  32'h3d54ba37 /* (6, 17, 3) */,
  32'h3d240321 /* (2, 17, 3) */,
  32'h3d29e985 /* (30, 13, 3) */,
  32'h3d54a03b /* (26, 13, 3) */,
  32'h3da99659 /* (22, 13, 3) */,
  32'h3e04d0b8 /* (18, 13, 3) */,
  32'h3e04d0b8 /* (14, 13, 3) */,
  32'h3da99659 /* (10, 13, 3) */,
  32'h3d54a03b /* (6, 13, 3) */,
  32'h3d29e985 /* (2, 13, 3) */,
  32'h3d12f42a /* (30, 9, 3) */,
  32'h3d215063 /* (26, 9, 3) */,
  32'h3d5dae2c /* (22, 9, 3) */,
  32'h3d9b2a7b /* (18, 9, 3) */,
  32'h3d9b2a7b /* (14, 9, 3) */,
  32'h3d5dae2c /* (10, 9, 3) */,
  32'h3d215063 /* (6, 9, 3) */,
  32'h3d12f42a /* (2, 9, 3) */,
  32'h3d3cd255 /* (30, 5, 3) */,
  32'h3d16d305 /* (26, 5, 3) */,
  32'h3d2344c4 /* (22, 5, 3) */,
  32'h3d487174 /* (18, 5, 3) */,
  32'h3d487174 /* (14, 5, 3) */,
  32'h3d2344c4 /* (10, 5, 3) */,
  32'h3d16d305 /* (6, 5, 3) */,
  32'h3d3cd255 /* (2, 5, 3) */,
  32'h3dbfa8df /* (30, 1, 3) */,
  32'h3d2ba889 /* (26, 1, 3) */,
  32'h3d14c0fd /* (22, 1, 3) */,
  32'h3d276174 /* (18, 1, 3) */,
  32'h3d276174 /* (14, 1, 3) */,
  32'h3d14c0fd /* (10, 1, 3) */,
  32'h3d2ba889 /* (6, 1, 3) */,
  32'h3dbfa8df /* (2, 1, 3) */,
  32'h3d960c3c /* (29, 29, 31) */,
  32'h3d1c3652 /* (25, 29, 31) */,
  32'h3d1a3ccf /* (21, 29, 31) */,
  32'h3d202be8 /* (17, 29, 31) */,
  32'h3d269671 /* (13, 29, 31) */,
  32'h3d126006 /* (9, 29, 31) */,
  32'h3d45ae9a /* (5, 29, 31) */,
  32'h3deb372d /* (1, 29, 31) */,
  32'h3d1c3652 /* (29, 25, 31) */,
  32'h3d167b79 /* (25, 25, 31) */,
  32'h3d3efe62 /* (21, 25, 31) */,
  32'h3d5d3ed0 /* (17, 25, 31) */,
  32'h3d5c17b6 /* (13, 25, 31) */,
  32'h3d245baa /* (9, 25, 31) */,
  32'h3d151e01 /* (5, 25, 31) */,
  32'h3d2402bf /* (1, 25, 31) */,
  32'h3d1a3ccf /* (29, 21, 31) */,
  32'h3d3efe62 /* (25, 21, 31) */,
  32'h3d9352ec /* (21, 21, 31) */,
  32'h3dc031e4 /* (17, 21, 31) */,
  32'h3db58f74 /* (13, 21, 31) */,
  32'h3d68852c /* (9, 21, 31) */,
  32'h3d26c9db /* (5, 21, 31) */,
  32'h3d151591 /* (1, 21, 31) */,
  32'h3d202be8 /* (29, 17, 31) */,
  32'h3d5d3ed0 /* (25, 17, 31) */,
  32'h3dc031e4 /* (21, 17, 31) */,
  32'h3e09bd27 /* (17, 17, 31) */,
  32'h3df92d6c /* (13, 17, 31) */,
  32'h3d8f3655 /* (9, 17, 31) */,
  32'h3d35f880 /* (5, 17, 31) */,
  32'h3d167d01 /* (1, 17, 31) */,
  32'h3d269671 /* (29, 13, 31) */,
  32'h3d5c17b6 /* (25, 13, 31) */,
  32'h3db58f74 /* (21, 13, 31) */,
  32'h3df92d6c /* (17, 13, 31) */,
  32'h3de602d9 /* (13, 13, 31) */,
  32'h3d8ac476 /* (9, 13, 31) */,
  32'h3d398f3f /* (5, 13, 31) */,
  32'h3d1e42f1 /* (1, 13, 31) */,
  32'h3d126006 /* (29, 9, 31) */,
  32'h3d245baa /* (25, 9, 31) */,
  32'h3d68852c /* (21, 9, 31) */,
  32'h3d8f3655 /* (17, 9, 31) */,
  32'h3d8ac476 /* (13, 9, 31) */,
  32'h3d3ee791 /* (9, 9, 31) */,
  32'h3d170f20 /* (5, 9, 31) */,
  32'h3d11a602 /* (1, 9, 31) */,
  32'h3d45ae9a /* (29, 5, 31) */,
  32'h3d151e01 /* (25, 5, 31) */,
  32'h3d26c9db /* (21, 5, 31) */,
  32'h3d35f880 /* (17, 5, 31) */,
  32'h3d398f3f /* (13, 5, 31) */,
  32'h3d170f20 /* (9, 5, 31) */,
  32'h3d249f29 /* (5, 5, 31) */,
  32'h3d6890ff /* (1, 5, 31) */,
  32'h3deb372d /* (29, 1, 31) */,
  32'h3d2402bf /* (25, 1, 31) */,
  32'h3d151591 /* (21, 1, 31) */,
  32'h3d167d01 /* (17, 1, 31) */,
  32'h3d1e42f1 /* (13, 1, 31) */,
  32'h3d11a602 /* (9, 1, 31) */,
  32'h3d6890ff /* (5, 1, 31) */,
  32'h3ec3aed4 /* (1, 1, 31) */,
  32'h3d314afb /* (29, 29, 27) */,
  32'h3d147808 /* (25, 29, 27) */,
  32'h3d2e4aa1 /* (21, 29, 27) */,
  32'h3d424fe8 /* (17, 29, 27) */,
  32'h3d4466f8 /* (13, 29, 27) */,
  32'h3d1addce /* (9, 29, 27) */,
  32'h3d1ccb4c /* (5, 29, 27) */,
  32'h3d45ae9a /* (1, 29, 27) */,
  32'h3d147808 /* (29, 25, 27) */,
  32'h3d21f168 /* (25, 25, 27) */,
  32'h3d5ff008 /* (21, 25, 27) */,
  32'h3d880917 /* (17, 25, 27) */,
  32'h3d849ae2 /* (13, 25, 27) */,
  32'h3d39ba58 /* (9, 25, 27) */,
  32'h3d170afd /* (5, 25, 27) */,
  32'h3d151e01 /* (1, 25, 27) */,
  32'h3d2e4aa1 /* (29, 21, 27) */,
  32'h3d5ff008 /* (25, 21, 27) */,
  32'h3db345e2 /* (21, 21, 27) */,
  32'h3df05994 /* (17, 21, 27) */,
  32'h3de04254 /* (13, 21, 27) */,
  32'h3d8b02ad /* (9, 21, 27) */,
  32'h3d3fb488 /* (5, 21, 27) */,
  32'h3d26c9db /* (1, 21, 27) */,
  32'h3d424fe8 /* (29, 17, 27) */,
  32'h3d880917 /* (25, 17, 27) */,
  32'h3df05994 /* (21, 17, 27) */,
  32'h3e2edbb4 /* (17, 17, 27) */,
  32'h3e1d0a10 /* (13, 17, 27) */,
  32'h3db198fc /* (9, 17, 27) */,
  32'h3d5e11d0 /* (5, 17, 27) */,
  32'h3d35f880 /* (1, 17, 27) */,
  32'h3d4466f8 /* (29, 13, 27) */,
  32'h3d849ae2 /* (25, 13, 27) */,
  32'h3de04254 /* (21, 13, 27) */,
  32'h3e1d0a10 /* (17, 13, 27) */,
  32'h3e0f99f2 /* (13, 13, 27) */,
  32'h3da95898 /* (9, 13, 27) */,
  32'h3d5ce99d /* (5, 13, 27) */,
  32'h3d398f3f /* (1, 13, 27) */,
  32'h3d1addce /* (29, 9, 27) */,
  32'h3d39ba58 /* (25, 9, 27) */,
  32'h3d8b02ad /* (21, 9, 27) */,
  32'h3db198fc /* (17, 9, 27) */,
  32'h3da95898 /* (13, 9, 27) */,
  32'h3d5e7d3b /* (9, 9, 27) */,
  32'h3d24f869 /* (5, 9, 27) */,
  32'h3d170f20 /* (1, 9, 27) */,
  32'h3d1ccb4c /* (29, 5, 27) */,
  32'h3d170afd /* (25, 5, 27) */,
  32'h3d3fb488 /* (21, 5, 27) */,
  32'h3d5e11d0 /* (17, 5, 27) */,
  32'h3d5ce99d /* (13, 5, 27) */,
  32'h3d24f869 /* (9, 5, 27) */,
  32'h3d15ac37 /* (5, 5, 27) */,
  32'h3d249f29 /* (1, 5, 27) */,
  32'h3d45ae9a /* (29, 1, 27) */,
  32'h3d151e01 /* (25, 1, 27) */,
  32'h3d26c9db /* (21, 1, 27) */,
  32'h3d35f880 /* (17, 1, 27) */,
  32'h3d398f3f /* (13, 1, 27) */,
  32'h3d170f20 /* (9, 1, 27) */,
  32'h3d249f29 /* (5, 1, 27) */,
  32'h3d6890ff /* (1, 1, 27) */,
  32'h3d144047 /* (29, 29, 23) */,
  32'h3d2aad03 /* (25, 29, 23) */,
  32'h3d767d5d /* (21, 29, 23) */,
  32'h3d99caa3 /* (17, 29, 23) */,
  32'h3d942dc4 /* (13, 29, 23) */,
  32'h3d48821f /* (9, 29, 23) */,
  32'h3d1addce /* (5, 29, 23) */,
  32'h3d126006 /* (1, 29, 23) */,
  32'h3d2aad03 /* (29, 25, 23) */,
  32'h3d563bcb /* (25, 25, 23) */,
  32'h3da777c1 /* (21, 25, 23) */,
  32'h3ddc94c6 /* (17, 25, 23) */,
  32'h3dcf79e9 /* (13, 25, 23) */,
  32'h3d8354ed /* (9, 25, 23) */,
  32'h3d39ba58 /* (5, 25, 23) */,
  32'h3d245baa /* (1, 25, 23) */,
  32'h3d767d5d /* (29, 21, 23) */,
  32'h3da777c1 /* (25, 21, 23) */,
  32'h3e0ea5fd /* (21, 21, 23) */,
  32'h3e49046a /* (17, 21, 23) */,
  32'h3e37494b /* (13, 21, 23) */,
  32'h3dd6aa1b /* (9, 21, 23) */,
  32'h3d8b02ad /* (5, 21, 23) */,
  32'h3d68852c /* (1, 21, 23) */,
  32'h3d99caa3 /* (29, 17, 23) */,
  32'h3ddc94c6 /* (25, 17, 23) */,
  32'h3e49046a /* (21, 17, 23) */,
  32'h3e969108 /* (17, 17, 23) */,
  32'h3e8557f4 /* (13, 17, 23) */,
  32'h3e123783 /* (9, 17, 23) */,
  32'h3db198fc /* (5, 17, 23) */,
  32'h3d8f3655 /* (1, 17, 23) */,
  32'h3d942dc4 /* (29, 13, 23) */,
  32'h3dcf79e9 /* (25, 13, 23) */,
  32'h3e37494b /* (21, 13, 23) */,
  32'h3e8557f4 /* (17, 13, 23) */,
  32'h3e6f82ab /* (13, 13, 23) */,
  32'h3e076ebd /* (9, 13, 23) */,
  32'h3da95898 /* (5, 13, 23) */,
  32'h3d8ac476 /* (1, 13, 23) */,
  32'h3d48821f /* (29, 9, 23) */,
  32'h3d8354ed /* (25, 9, 23) */,
  32'h3dd6aa1b /* (21, 9, 23) */,
  32'h3e123783 /* (17, 9, 23) */,
  32'h3e076ebd /* (13, 9, 23) */,
  32'h3da4cfbf /* (9, 9, 23) */,
  32'h3d5e7d3b /* (5, 9, 23) */,
  32'h3d3ee791 /* (1, 9, 23) */,
  32'h3d1addce /* (29, 5, 23) */,
  32'h3d39ba58 /* (25, 5, 23) */,
  32'h3d8b02ad /* (21, 5, 23) */,
  32'h3db198fc /* (17, 5, 23) */,
  32'h3da95898 /* (13, 5, 23) */,
  32'h3d5e7d3b /* (9, 5, 23) */,
  32'h3d24f869 /* (5, 5, 23) */,
  32'h3d170f20 /* (1, 5, 23) */,
  32'h3d126006 /* (29, 1, 23) */,
  32'h3d245baa /* (25, 1, 23) */,
  32'h3d68852c /* (21, 1, 23) */,
  32'h3d8f3655 /* (17, 1, 23) */,
  32'h3d8ac476 /* (13, 1, 23) */,
  32'h3d3ee791 /* (9, 1, 23) */,
  32'h3d170f20 /* (5, 1, 23) */,
  32'h3d11a602 /* (1, 1, 23) */,
  32'h3d2fb3ed /* (29, 29, 19) */,
  32'h3d69f6ae /* (25, 29, 19) */,
  32'h3dc2b35d /* (21, 29, 19) */,
  32'h3e068db8 /* (17, 29, 19) */,
  32'h3df79892 /* (13, 29, 19) */,
  32'h3d942dc4 /* (9, 29, 19) */,
  32'h3d4466f8 /* (5, 29, 19) */,
  32'h3d269671 /* (1, 29, 19) */,
  32'h3d69f6ae /* (29, 25, 19) */,
  32'h3da0c360 /* (25, 25, 19) */,
  32'h3e0aca9a /* (21, 25, 19) */,
  32'h3e45db44 /* (17, 25, 19) */,
  32'h3e336d1b /* (13, 25, 19) */,
  32'h3dcf79e9 /* (9, 25, 19) */,
  32'h3d849ae2 /* (5, 25, 19) */,
  32'h3d5c17b6 /* (1, 25, 19) */,
  32'h3dc2b35d /* (29, 21, 19) */,
  32'h3e0aca9a /* (25, 21, 19) */,
  32'h3e7af74d /* (21, 21, 19) */,
  32'h3eba8e90 /* (17, 21, 19) */,
  32'h3ea5d30f /* (13, 21, 19) */,
  32'h3e37494b /* (9, 21, 19) */,
  32'h3de04254 /* (5, 21, 19) */,
  32'h3db58f74 /* (1, 21, 19) */,
  32'h3e068db8 /* (29, 17, 19) */,
  32'h3e45db44 /* (25, 17, 19) */,
  32'h3eba8e90 /* (21, 17, 19) */,
  32'h3f1092e5 /* (17, 17, 19) */,
  32'h3efbd9fe /* (13, 17, 19) */,
  32'h3e8557f4 /* (9, 17, 19) */,
  32'h3e1d0a10 /* (5, 17, 19) */,
  32'h3df92d6c /* (1, 17, 19) */,
  32'h3df79892 /* (29, 13, 19) */,
  32'h3e336d1b /* (25, 13, 19) */,
  32'h3ea5d30f /* (21, 13, 19) */,
  32'h3efbd9fe /* (17, 13, 19) */,
  32'h3edd8ee5 /* (13, 13, 19) */,
  32'h3e6f82ab /* (9, 13, 19) */,
  32'h3e0f99f2 /* (5, 13, 19) */,
  32'h3de602d9 /* (1, 13, 19) */,
  32'h3d942dc4 /* (29, 9, 19) */,
  32'h3dcf79e9 /* (25, 9, 19) */,
  32'h3e37494b /* (21, 9, 19) */,
  32'h3e8557f4 /* (17, 9, 19) */,
  32'h3e6f82ab /* (13, 9, 19) */,
  32'h3e076ebd /* (9, 9, 19) */,
  32'h3da95898 /* (5, 9, 19) */,
  32'h3d8ac476 /* (1, 9, 19) */,
  32'h3d4466f8 /* (29, 5, 19) */,
  32'h3d849ae2 /* (25, 5, 19) */,
  32'h3de04254 /* (21, 5, 19) */,
  32'h3e1d0a10 /* (17, 5, 19) */,
  32'h3e0f99f2 /* (13, 5, 19) */,
  32'h3da95898 /* (9, 5, 19) */,
  32'h3d5ce99d /* (5, 5, 19) */,
  32'h3d398f3f /* (1, 5, 19) */,
  32'h3d269671 /* (29, 1, 19) */,
  32'h3d5c17b6 /* (25, 1, 19) */,
  32'h3db58f74 /* (21, 1, 19) */,
  32'h3df92d6c /* (17, 1, 19) */,
  32'h3de602d9 /* (13, 1, 19) */,
  32'h3d8ac476 /* (9, 1, 19) */,
  32'h3d398f3f /* (5, 1, 19) */,
  32'h3d1e42f1 /* (1, 1, 19) */,
  32'h3d2aacf2 /* (29, 29, 15) */,
  32'h3d6ce397 /* (25, 29, 15) */,
  32'h3dceffa6 /* (21, 29, 15) */,
  32'h3e151f83 /* (17, 29, 15) */,
  32'h3e068db8 /* (13, 29, 15) */,
  32'h3d99caa3 /* (9, 29, 15) */,
  32'h3d424fe8 /* (5, 29, 15) */,
  32'h3d202be8 /* (1, 29, 15) */,
  32'h3d6ce397 /* (29, 25, 15) */,
  32'h3da7bf05 /* (25, 25, 15) */,
  32'h3e165b49 /* (21, 25, 15) */,
  32'h3e5db918 /* (17, 25, 15) */,
  32'h3e45db44 /* (13, 25, 15) */,
  32'h3ddc94c6 /* (9, 25, 15) */,
  32'h3d880917 /* (5, 25, 15) */,
  32'h3d5d3ed0 /* (1, 25, 15) */,
  32'h3dceffa6 /* (29, 21, 15) */,
  32'h3e165b49 /* (25, 21, 15) */,
  32'h3e8b66c2 /* (21, 21, 15) */,
  32'h3ed4648a /* (17, 21, 15) */,
  32'h3eba8e90 /* (13, 21, 15) */,
  32'h3e49046a /* (9, 21, 15) */,
  32'h3df05994 /* (5, 21, 15) */,
  32'h3dc031e4 /* (1, 21, 15) */,
  32'h3e151f83 /* (29, 17, 15) */,
  32'h3e5db918 /* (25, 17, 15) */,
  32'h3ed4648a /* (21, 17, 15) */,
  32'h3f275a64 /* (17, 17, 15) */,
  32'h3f1092e5 /* (13, 17, 15) */,
  32'h3e969108 /* (9, 17, 15) */,
  32'h3e2edbb4 /* (5, 17, 15) */,
  32'h3e09bd27 /* (1, 17, 15) */,
  32'h3e068db8 /* (29, 13, 15) */,
  32'h3e45db44 /* (25, 13, 15) */,
  32'h3eba8e90 /* (21, 13, 15) */,
  32'h3f1092e5 /* (17, 13, 15) */,
  32'h3efbd9fe /* (13, 13, 15) */,
  32'h3e8557f4 /* (9, 13, 15) */,
  32'h3e1d0a10 /* (5, 13, 15) */,
  32'h3df92d6c /* (1, 13, 15) */,
  32'h3d99caa3 /* (29, 9, 15) */,
  32'h3ddc94c6 /* (25, 9, 15) */,
  32'h3e49046a /* (21, 9, 15) */,
  32'h3e969108 /* (17, 9, 15) */,
  32'h3e8557f4 /* (13, 9, 15) */,
  32'h3e123783 /* (9, 9, 15) */,
  32'h3db198fc /* (5, 9, 15) */,
  32'h3d8f3655 /* (1, 9, 15) */,
  32'h3d424fe8 /* (29, 5, 15) */,
  32'h3d880917 /* (25, 5, 15) */,
  32'h3df05994 /* (21, 5, 15) */,
  32'h3e2edbb4 /* (17, 5, 15) */,
  32'h3e1d0a10 /* (13, 5, 15) */,
  32'h3db198fc /* (9, 5, 15) */,
  32'h3d5e11d0 /* (5, 5, 15) */,
  32'h3d35f880 /* (1, 5, 15) */,
  32'h3d202be8 /* (29, 1, 15) */,
  32'h3d5d3ed0 /* (25, 1, 15) */,
  32'h3dc031e4 /* (21, 1, 15) */,
  32'h3e09bd27 /* (17, 1, 15) */,
  32'h3df92d6c /* (13, 1, 15) */,
  32'h3d8f3655 /* (9, 1, 15) */,
  32'h3d35f880 /* (5, 1, 15) */,
  32'h3d167d01 /* (1, 1, 15) */,
  32'h3d202a91 /* (29, 29, 11) */,
  32'h3d490aba /* (25, 29, 11) */,
  32'h3d9d27e1 /* (21, 29, 11) */,
  32'h3dceffa6 /* (17, 29, 11) */,
  32'h3dc2b35d /* (13, 29, 11) */,
  32'h3d767d5d /* (9, 29, 11) */,
  32'h3d2e4aa1 /* (5, 29, 11) */,
  32'h3d1a3ccf /* (1, 29, 11) */,
  32'h3d490aba /* (29, 25, 11) */,
  32'h3d84ce75 /* (25, 25, 11) */,
  32'h3ddb1c7f /* (21, 25, 11) */,
  32'h3e165b49 /* (17, 25, 11) */,
  32'h3e0aca9a /* (13, 25, 11) */,
  32'h3da777c1 /* (9, 25, 11) */,
  32'h3d5ff008 /* (5, 25, 11) */,
  32'h3d3efe62 /* (1, 25, 11) */,
  32'h3d9d27e1 /* (29, 21, 11) */,
  32'h3ddb1c7f /* (25, 21, 11) */,
  32'h3e4089a2 /* (21, 21, 11) */,
  32'h3e8b66c2 /* (17, 21, 11) */,
  32'h3e7af74d /* (13, 21, 11) */,
  32'h3e0ea5fd /* (9, 21, 11) */,
  32'h3db345e2 /* (5, 21, 11) */,
  32'h3d9352ec /* (1, 21, 11) */,
  32'h3dceffa6 /* (29, 17, 11) */,
  32'h3e165b49 /* (25, 17, 11) */,
  32'h3e8b66c2 /* (21, 17, 11) */,
  32'h3ed4648a /* (17, 17, 11) */,
  32'h3eba8e90 /* (13, 17, 11) */,
  32'h3e49046a /* (9, 17, 11) */,
  32'h3df05994 /* (5, 17, 11) */,
  32'h3dc031e4 /* (1, 17, 11) */,
  32'h3dc2b35d /* (29, 13, 11) */,
  32'h3e0aca9a /* (25, 13, 11) */,
  32'h3e7af74d /* (21, 13, 11) */,
  32'h3eba8e90 /* (17, 13, 11) */,
  32'h3ea5d30f /* (13, 13, 11) */,
  32'h3e37494b /* (9, 13, 11) */,
  32'h3de04254 /* (5, 13, 11) */,
  32'h3db58f74 /* (1, 13, 11) */,
  32'h3d767d5d /* (29, 9, 11) */,
  32'h3da777c1 /* (25, 9, 11) */,
  32'h3e0ea5fd /* (21, 9, 11) */,
  32'h3e49046a /* (17, 9, 11) */,
  32'h3e37494b /* (13, 9, 11) */,
  32'h3dd6aa1b /* (9, 9, 11) */,
  32'h3d8b02ad /* (5, 9, 11) */,
  32'h3d68852c /* (1, 9, 11) */,
  32'h3d2e4aa1 /* (29, 5, 11) */,
  32'h3d5ff008 /* (25, 5, 11) */,
  32'h3db345e2 /* (21, 5, 11) */,
  32'h3df05994 /* (17, 5, 11) */,
  32'h3de04254 /* (13, 5, 11) */,
  32'h3d8b02ad /* (9, 5, 11) */,
  32'h3d3fb488 /* (5, 5, 11) */,
  32'h3d26c9db /* (1, 5, 11) */,
  32'h3d1a3ccf /* (29, 1, 11) */,
  32'h3d3efe62 /* (25, 1, 11) */,
  32'h3d9352ec /* (21, 1, 11) */,
  32'h3dc031e4 /* (17, 1, 11) */,
  32'h3db58f74 /* (13, 1, 11) */,
  32'h3d68852c /* (9, 1, 11) */,
  32'h3d26c9db /* (5, 1, 11) */,
  32'h3d151591 /* (1, 1, 11) */,
  32'h3d179239 /* (29, 29, 7) */,
  32'h3d1969a9 /* (25, 29, 7) */,
  32'h3d490aba /* (21, 29, 7) */,
  32'h3d6ce397 /* (17, 29, 7) */,
  32'h3d69f6ae /* (13, 29, 7) */,
  32'h3d2aad03 /* (9, 29, 7) */,
  32'h3d147808 /* (5, 29, 7) */,
  32'h3d1c3652 /* (1, 29, 7) */,
  32'h3d1969a9 /* (29, 25, 7) */,
  32'h3d348078 /* (25, 25, 7) */,
  32'h3d84ce75 /* (21, 25, 7) */,
  32'h3da7bf05 /* (17, 25, 7) */,
  32'h3da0c360 /* (13, 25, 7) */,
  32'h3d563bcb /* (9, 25, 7) */,
  32'h3d21f168 /* (5, 25, 7) */,
  32'h3d167b79 /* (1, 25, 7) */,
  32'h3d490aba /* (29, 21, 7) */,
  32'h3d84ce75 /* (25, 21, 7) */,
  32'h3ddb1c7f /* (21, 21, 7) */,
  32'h3e165b49 /* (17, 21, 7) */,
  32'h3e0aca9a /* (13, 21, 7) */,
  32'h3da777c1 /* (9, 21, 7) */,
  32'h3d5ff008 /* (5, 21, 7) */,
  32'h3d3efe62 /* (1, 21, 7) */,
  32'h3d6ce397 /* (29, 17, 7) */,
  32'h3da7bf05 /* (25, 17, 7) */,
  32'h3e165b49 /* (21, 17, 7) */,
  32'h3e5db918 /* (17, 17, 7) */,
  32'h3e45db44 /* (13, 17, 7) */,
  32'h3ddc94c6 /* (9, 17, 7) */,
  32'h3d880917 /* (5, 17, 7) */,
  32'h3d5d3ed0 /* (1, 17, 7) */,
  32'h3d69f6ae /* (29, 13, 7) */,
  32'h3da0c360 /* (25, 13, 7) */,
  32'h3e0aca9a /* (21, 13, 7) */,
  32'h3e45db44 /* (17, 13, 7) */,
  32'h3e336d1b /* (13, 13, 7) */,
  32'h3dcf79e9 /* (9, 13, 7) */,
  32'h3d849ae2 /* (5, 13, 7) */,
  32'h3d5c17b6 /* (1, 13, 7) */,
  32'h3d2aad03 /* (29, 9, 7) */,
  32'h3d563bcb /* (25, 9, 7) */,
  32'h3da777c1 /* (21, 9, 7) */,
  32'h3ddc94c6 /* (17, 9, 7) */,
  32'h3dcf79e9 /* (13, 9, 7) */,
  32'h3d8354ed /* (9, 9, 7) */,
  32'h3d39ba58 /* (5, 9, 7) */,
  32'h3d245baa /* (1, 9, 7) */,
  32'h3d147808 /* (29, 5, 7) */,
  32'h3d21f168 /* (25, 5, 7) */,
  32'h3d5ff008 /* (21, 5, 7) */,
  32'h3d880917 /* (17, 5, 7) */,
  32'h3d849ae2 /* (13, 5, 7) */,
  32'h3d39ba58 /* (9, 5, 7) */,
  32'h3d170afd /* (5, 5, 7) */,
  32'h3d151e01 /* (1, 5, 7) */,
  32'h3d1c3652 /* (29, 1, 7) */,
  32'h3d167b79 /* (25, 1, 7) */,
  32'h3d3efe62 /* (21, 1, 7) */,
  32'h3d5d3ed0 /* (17, 1, 7) */,
  32'h3d5c17b6 /* (13, 1, 7) */,
  32'h3d245baa /* (9, 1, 7) */,
  32'h3d151e01 /* (5, 1, 7) */,
  32'h3d2402bf /* (1, 1, 7) */,
  32'h3d68b01f /* (29, 29, 3) */,
  32'h3d179239 /* (25, 29, 3) */,
  32'h3d202a91 /* (21, 29, 3) */,
  32'h3d2aacf2 /* (17, 29, 3) */,
  32'h3d2fb3ed /* (13, 29, 3) */,
  32'h3d144047 /* (9, 29, 3) */,
  32'h3d314afb /* (5, 29, 3) */,
  32'h3d960c3c /* (1, 29, 3) */,
  32'h3d179239 /* (29, 25, 3) */,
  32'h3d1969a9 /* (25, 25, 3) */,
  32'h3d490aba /* (21, 25, 3) */,
  32'h3d6ce397 /* (17, 25, 3) */,
  32'h3d69f6ae /* (13, 25, 3) */,
  32'h3d2aad03 /* (9, 25, 3) */,
  32'h3d147808 /* (5, 25, 3) */,
  32'h3d1c3652 /* (1, 25, 3) */,
  32'h3d202a91 /* (29, 21, 3) */,
  32'h3d490aba /* (25, 21, 3) */,
  32'h3d9d27e1 /* (21, 21, 3) */,
  32'h3dceffa6 /* (17, 21, 3) */,
  32'h3dc2b35d /* (13, 21, 3) */,
  32'h3d767d5d /* (9, 21, 3) */,
  32'h3d2e4aa1 /* (5, 21, 3) */,
  32'h3d1a3ccf /* (1, 21, 3) */,
  32'h3d2aacf2 /* (29, 17, 3) */,
  32'h3d6ce397 /* (25, 17, 3) */,
  32'h3dceffa6 /* (21, 17, 3) */,
  32'h3e151f83 /* (17, 17, 3) */,
  32'h3e068db8 /* (13, 17, 3) */,
  32'h3d99caa3 /* (9, 17, 3) */,
  32'h3d424fe8 /* (5, 17, 3) */,
  32'h3d202be8 /* (1, 17, 3) */,
  32'h3d2fb3ed /* (29, 13, 3) */,
  32'h3d69f6ae /* (25, 13, 3) */,
  32'h3dc2b35d /* (21, 13, 3) */,
  32'h3e068db8 /* (17, 13, 3) */,
  32'h3df79892 /* (13, 13, 3) */,
  32'h3d942dc4 /* (9, 13, 3) */,
  32'h3d4466f8 /* (5, 13, 3) */,
  32'h3d269671 /* (1, 13, 3) */,
  32'h3d144047 /* (29, 9, 3) */,
  32'h3d2aad03 /* (25, 9, 3) */,
  32'h3d767d5d /* (21, 9, 3) */,
  32'h3d99caa3 /* (17, 9, 3) */,
  32'h3d942dc4 /* (13, 9, 3) */,
  32'h3d48821f /* (9, 9, 3) */,
  32'h3d1addce /* (5, 9, 3) */,
  32'h3d126006 /* (1, 9, 3) */,
  32'h3d314afb /* (29, 5, 3) */,
  32'h3d147808 /* (25, 5, 3) */,
  32'h3d2e4aa1 /* (21, 5, 3) */,
  32'h3d424fe8 /* (17, 5, 3) */,
  32'h3d4466f8 /* (13, 5, 3) */,
  32'h3d1addce /* (9, 5, 3) */,
  32'h3d1ccb4c /* (5, 5, 3) */,
  32'h3d45ae9a /* (1, 5, 3) */,
  32'h3d960c3c /* (29, 1, 3) */,
  32'h3d1c3652 /* (25, 1, 3) */,
  32'h3d1a3ccf /* (21, 1, 3) */,
  32'h3d202be8 /* (17, 1, 3) */,
  32'h3d269671 /* (13, 1, 3) */,
  32'h3d126006 /* (9, 1, 3) */,
  32'h3d45ae9a /* (5, 1, 3) */,
  32'h3deb372d /* (1, 1, 3) */,
  32'h3d6eb36b /* (28, 29, 31) */,
  32'h3d146963 /* (24, 29, 31) */,
  32'h3d210eee /* (20, 29, 31) */,
  32'h3d0fbc59 /* (16, 29, 31) */,
  32'h3d210eee /* (12, 29, 31) */,
  32'h3d146963 /* (8, 29, 31) */,
  32'h3d6eb36b /* (4, 29, 31) */,
  32'h3dff9e3f /* (0, 29, 31) */,
  32'h3d17ff6b /* (28, 25, 31) */,
  32'h3d1bb8b6 /* (24, 25, 31) */,
  32'h3d4ea8e5 /* (20, 25, 31) */,
  32'h3d49f75a /* (16, 25, 31) */,
  32'h3d4ea8e5 /* (12, 25, 31) */,
  32'h3d1bb8b6 /* (8, 25, 31) */,
  32'h3d17ff6b /* (4, 25, 31) */,
  32'h3d25463b /* (0, 25, 31) */,
  32'h3d1f5dc3 /* (28, 21, 31) */,
  32'h3d513c3d /* (24, 21, 31) */,
  32'h3da53628 /* (20, 21, 31) */,
  32'h3db336e0 /* (16, 21, 31) */,
  32'h3da53628 /* (12, 21, 31) */,
  32'h3d513c3d /* (8, 21, 31) */,
  32'h3d1f5dc3 /* (4, 21, 31) */,
  32'h3d147e90 /* (0, 21, 31) */,
  32'h3d294c4b /* (28, 17, 31) */,
  32'h3d7a003f /* (24, 17, 31) */,
  32'h3ddd43c2 /* (20, 17, 31) */,
  32'h3e02e976 /* (16, 17, 31) */,
  32'h3ddd43c2 /* (12, 17, 31) */,
  32'h3d7a003f /* (8, 17, 31) */,
  32'h3d294c4b /* (4, 17, 31) */,
  32'h3d155505 /* (0, 17, 31) */,
  32'h3d2e802a /* (28, 13, 31) */,
  32'h3d7573b6 /* (24, 13, 31) */,
  32'h3dce8d02 /* (20, 13, 31) */,
  32'h3deaafef /* (16, 13, 31) */,
  32'h3dce8d02 /* (12, 13, 31) */,
  32'h3d7573b6 /* (8, 13, 31) */,
  32'h3d2e802a /* (4, 13, 31) */,
  32'h3d1d4601 /* (0, 13, 31) */,
  32'h3d13f199 /* (28, 9, 31) */,
  32'h3d2fba80 /* (24, 9, 31) */,
  32'h3d803124 /* (20, 9, 31) */,
  32'h3d8420c9 /* (16, 9, 31) */,
  32'h3d803124 /* (12, 9, 31) */,
  32'h3d2fba80 /* (8, 9, 31) */,
  32'h3d13f199 /* (4, 9, 31) */,
  32'h3d11a5c6 /* (0, 9, 31) */,
  32'h3d334ee4 /* (28, 5, 31) */,
  32'h3d1412fd /* (24, 5, 31) */,
  32'h3d310ad3 /* (20, 5, 31) */,
  32'h3d24852f /* (16, 5, 31) */,
  32'h3d310ad3 /* (12, 5, 31) */,
  32'h3d1412fd /* (8, 5, 31) */,
  32'h3d334ee4 /* (4, 5, 31) */,
  32'h3d6e9998 /* (0, 5, 31) */,
  32'h3d9c757b /* (28, 1, 31) */,
  32'h3d1704d7 /* (24, 1, 31) */,
  32'h3d1a2df1 /* (20, 1, 31) */,
  32'h3d067e68 /* (16, 1, 31) */,
  32'h3d1a2df1 /* (12, 1, 31) */,
  32'h3d1704d7 /* (8, 1, 31) */,
  32'h3d9c757b /* (4, 1, 31) */,
  32'h3f10fe39 /* (0, 1, 31) */,
  32'h3d25f5ce /* (28, 29, 27) */,
  32'h3d15d660 /* (24, 29, 27) */,
  32'h3d3a4ebb /* (20, 29, 27) */,
  32'h3d3046d8 /* (16, 29, 27) */,
  32'h3d3a4ebb /* (12, 29, 27) */,
  32'h3d15d660 /* (8, 29, 27) */,
  32'h3d25f5ce /* (4, 29, 27) */,
  32'h3d490b0e /* (0, 29, 27) */,
  32'h3d1508af /* (28, 25, 27) */,
  32'h3d2bff3e /* (24, 25, 27) */,
  32'h3d75e4d4 /* (20, 25, 27) */,
  32'h3d7a662c /* (16, 25, 27) */,
  32'h3d75e4d4 /* (12, 25, 27) */,
  32'h3d2bff3e /* (8, 25, 27) */,
  32'h3d1508af /* (4, 25, 27) */,
  32'h3d154f7b /* (0, 25, 27) */,
  32'h3d358341 /* (28, 21, 27) */,
  32'h3d77c8fd /* (24, 21, 27) */,
  32'h3dca9d53 /* (20, 21, 27) */,
  32'h3de14ffa /* (16, 21, 27) */,
  32'h3dca9d53 /* (12, 21, 27) */,
  32'h3d77c8fd /* (8, 21, 27) */,
  32'h3d358341 /* (4, 21, 27) */,
  32'h3d25e815 /* (0, 21, 27) */,
  32'h3d4def9b /* (28, 17, 27) */,
  32'h3d9a5b6b /* (24, 17, 27) */,
  32'h3e0ae903 /* (20, 17, 27) */,
  32'h3e26bbbb /* (16, 17, 27) */,
  32'h3e0ae903 /* (12, 17, 27) */,
  32'h3d9a5b6b /* (8, 17, 27) */,
  32'h3d4def9b /* (4, 17, 27) */,
  32'h3d347f0a /* (0, 17, 27) */,
  32'h3d4ea6a0 /* (28, 13, 27) */,
  32'h3d94d380 /* (24, 13, 27) */,
  32'h3e00477d /* (20, 13, 27) */,
  32'h3e1486b7 /* (16, 13, 27) */,
  32'h3e00477d /* (12, 13, 27) */,
  32'h3d94d380 /* (8, 13, 27) */,
  32'h3d4ea6a0 /* (4, 13, 27) */,
  32'h3d384488 /* (0, 13, 27) */,
  32'h3d1ee50b /* (28, 9, 27) */,
  32'h3d49c96c /* (24, 9, 27) */,
  32'h3d9af1c2 /* (20, 9, 27) */,
  32'h3da4f2f4 /* (16, 9, 27) */,
  32'h3d9af1c2 /* (12, 9, 27) */,
  32'h3d49c96c /* (8, 9, 27) */,
  32'h3d1ee50b /* (4, 9, 27) */,
  32'h3d16a564 /* (0, 9, 27) */,
  32'h3d189061 /* (28, 5, 27) */,
  32'h3d1c4d38 /* (24, 5, 27) */,
  32'h3d4f6dfc /* (20, 5, 27) */,
  32'h3d4ab7f7 /* (16, 5, 27) */,
  32'h3d4f6dfc /* (12, 5, 27) */,
  32'h3d1c4d38 /* (8, 5, 27) */,
  32'h3d189061 /* (4, 5, 27) */,
  32'h3d25e3da /* (0, 5, 27) */,
  32'h3d334ee4 /* (28, 1, 27) */,
  32'h3d1412fd /* (24, 1, 27) */,
  32'h3d310ad3 /* (20, 1, 27) */,
  32'h3d24852f /* (16, 1, 27) */,
  32'h3d310ad3 /* (12, 1, 27) */,
  32'h3d1412fd /* (8, 1, 27) */,
  32'h3d334ee4 /* (4, 1, 27) */,
  32'h3d6e9998 /* (0, 1, 27) */,
  32'h3d16b5b2 /* (28, 29, 23) */,
  32'h3d37919e /* (24, 29, 23) */,
  32'h3d886b82 /* (20, 29, 23) */,
  32'h3d8e3848 /* (16, 29, 23) */,
  32'h3d886b82 /* (12, 29, 23) */,
  32'h3d37919e /* (8, 29, 23) */,
  32'h3d16b5b2 /* (4, 29, 23) */,
  32'h3d1237a7 /* (0, 29, 23) */,
  32'h3d30de15 /* (28, 25, 23) */,
  32'h3d6b8b35 /* (24, 25, 23) */,
  32'h3dbc51f9 /* (20, 25, 23) */,
  32'h3dce1075 /* (16, 25, 23) */,
  32'h3dbc51f9 /* (12, 25, 23) */,
  32'h3d6b8b35 /* (8, 25, 23) */,
  32'h3d30de15 /* (4, 25, 23) */,
  32'h3d23a039 /* (0, 25, 23) */,
  32'h3d81d711 /* (28, 21, 23) */,
  32'h3dbc4d73 /* (24, 21, 23) */,
  32'h3e23781b /* (20, 21, 23) */,
  32'h3e3e5da7 /* (16, 21, 23) */,
  32'h3e23781b /* (12, 21, 23) */,
  32'h3dbc4d73 /* (8, 21, 23) */,
  32'h3d81d711 /* (4, 21, 23) */,
  32'h3d66dac1 /* (0, 21, 23) */,
  32'h3da3c1ed /* (28, 17, 23) */,
  32'h3dfc30a3 /* (24, 17, 23) */,
  32'h3e6a25fd /* (20, 17, 23) */,
  32'h3e908107 /* (16, 17, 23) */,
  32'h3e6a25fd /* (12, 17, 23) */,
  32'h3dfc30a3 /* (8, 17, 23) */,
  32'h3da3c1ed /* (4, 17, 23) */,
  32'h3d8df2c1 /* (0, 17, 23) */,
  32'h3d9d0afa /* (28, 13, 23) */,
  32'h3deb6b6d /* (24, 13, 23) */,
  32'h3e53dc51 /* (20, 13, 23) */,
  32'h3e7e4b9d /* (16, 13, 23) */,
  32'h3e53dc51 /* (12, 13, 23) */,
  32'h3deb6b6d /* (8, 13, 23) */,
  32'h3d9d0afa /* (4, 13, 23) */,
  32'h3d89a49e /* (0, 13, 23) */,
  32'h3d51a9d2 /* (28, 9, 23) */,
  32'h3d921bde /* (24, 9, 23) */,
  32'h3df3b4f2 /* (20, 9, 23) */,
  32'h3e0981d7 /* (16, 9, 23) */,
  32'h3df3b4f2 /* (12, 9, 23) */,
  32'h3d921bde /* (8, 9, 23) */,
  32'h3d51a9d2 /* (4, 9, 23) */,
  32'h3d3dc47d /* (0, 9, 23) */,
  32'h3d1ee50b /* (28, 5, 23) */,
  32'h3d49c96c /* (24, 5, 23) */,
  32'h3d9af1c2 /* (20, 5, 23) */,
  32'h3da4f2f4 /* (16, 5, 23) */,
  32'h3d9af1c2 /* (12, 5, 23) */,
  32'h3d49c96c /* (8, 5, 23) */,
  32'h3d1ee50b /* (4, 5, 23) */,
  32'h3d16a564 /* (0, 5, 23) */,
  32'h3d13f199 /* (28, 1, 23) */,
  32'h3d2fba80 /* (24, 1, 23) */,
  32'h3d803124 /* (20, 1, 23) */,
  32'h3d8420c9 /* (16, 1, 23) */,
  32'h3d803124 /* (12, 1, 23) */,
  32'h3d2fba80 /* (8, 1, 23) */,
  32'h3d13f199 /* (4, 1, 23) */,
  32'h3d11a5c6 /* (0, 1, 23) */,
  32'h3d385879 /* (28, 29, 19) */,
  32'h3d82c188 /* (24, 29, 19) */,
  32'h3dddef48 /* (20, 29, 19) */,
  32'h3dfdd31f /* (16, 29, 19) */,
  32'h3dddef48 /* (12, 29, 19) */,
  32'h3d82c188 /* (8, 29, 19) */,
  32'h3d385879 /* (4, 29, 19) */,
  32'h3d258110 /* (0, 29, 19) */,
  32'h3d770afc /* (28, 25, 19) */,
  32'h3db56072 /* (24, 25, 19) */,
  32'h3e1f8cbf /* (20, 25, 19) */,
  32'h3e3bd4ee /* (16, 25, 19) */,
  32'h3e1f8cbf /* (12, 25, 19) */,
  32'h3db56072 /* (8, 25, 19) */,
  32'h3d770afc /* (4, 25, 19) */,
  32'h3d5a6fdd /* (0, 25, 19) */,
  32'h3dcf13a3 /* (28, 21, 19) */,
  32'h3e1e607d /* (24, 21, 19) */,
  32'h3e91dfe2 /* (20, 21, 19) */,
  32'h3eb2bd2a /* (16, 21, 19) */,
  32'h3e91dfe2 /* (12, 21, 19) */,
  32'h3e1e607d /* (8, 21, 19) */,
  32'h3dcf13a3 /* (4, 21, 19) */,
  32'h3db3fd83 /* (0, 21, 19) */,
  32'h3e0ff4ce /* (28, 17, 19) */,
  32'h3e640ba2 /* (24, 17, 19) */,
  32'h3edb3822 /* (20, 17, 19) */,
  32'h3f0bd969 /* (16, 17, 19) */,
  32'h3edb3822 /* (12, 17, 19) */,
  32'h3e640ba2 /* (8, 17, 19) */,
  32'h3e0ff4ce /* (4, 17, 19) */,
  32'h3df6cc6d /* (0, 17, 19) */,
  32'h3e0415cb /* (28, 13, 19) */,
  32'h3e4dd3dc /* (24, 13, 19) */,
  32'h3ec1d890 /* (20, 13, 19) */,
  32'h3ef27895 /* (16, 13, 19) */,
  32'h3ec1d890 /* (12, 13, 19) */,
  32'h3e4dd3dc /* (8, 13, 19) */,
  32'h3e0415cb /* (4, 13, 19) */,
  32'h3de3e928 /* (0, 13, 19) */,
  32'h3d9d0afa /* (28, 9, 19) */,
  32'h3deb6b6d /* (24, 9, 19) */,
  32'h3e53dc51 /* (20, 9, 19) */,
  32'h3e7e4b9d /* (16, 9, 19) */,
  32'h3e53dc51 /* (12, 9, 19) */,
  32'h3deb6b6d /* (8, 9, 19) */,
  32'h3d9d0afa /* (4, 9, 19) */,
  32'h3d89a49e /* (0, 9, 19) */,
  32'h3d4ea6a0 /* (28, 5, 19) */,
  32'h3d94d380 /* (24, 5, 19) */,
  32'h3e00477d /* (20, 5, 19) */,
  32'h3e1486b7 /* (16, 5, 19) */,
  32'h3e00477d /* (12, 5, 19) */,
  32'h3d94d380 /* (8, 5, 19) */,
  32'h3d4ea6a0 /* (4, 5, 19) */,
  32'h3d384488 /* (0, 5, 19) */,
  32'h3d2e802a /* (28, 1, 19) */,
  32'h3d7573b6 /* (24, 1, 19) */,
  32'h3dce8d02 /* (20, 1, 19) */,
  32'h3deaafef /* (16, 1, 19) */,
  32'h3dce8d02 /* (12, 1, 19) */,
  32'h3d7573b6 /* (8, 1, 19) */,
  32'h3d2e802a /* (4, 1, 19) */,
  32'h3d1d4601 /* (0, 1, 19) */,
  32'h3d349293 /* (28, 29, 15) */,
  32'h3d8608f0 /* (24, 29, 15) */,
  32'h3deea44d /* (20, 29, 15) */,
  32'h3e0de417 /* (16, 29, 15) */,
  32'h3deea44d /* (12, 29, 15) */,
  32'h3d8608f0 /* (8, 29, 15) */,
  32'h3d349293 /* (4, 29, 15) */,
  32'h3d1eeabe /* (0, 29, 15) */,
  32'h3d7b9f11 /* (28, 25, 15) */,
  32'h3dbf0444 /* (24, 25, 15) */,
  32'h3e2e6a71 /* (20, 25, 15) */,
  32'h3e540b9b /* (16, 25, 15) */,
  32'h3e2e6a71 /* (12, 25, 15) */,
  32'h3dbf0444 /* (8, 25, 15) */,
  32'h3d7b9f11 /* (4, 25, 15) */,
  32'h3d5b6048 /* (0, 25, 15) */,
  32'h3ddcf428 /* (28, 21, 15) */,
  32'h3e2c9c6c /* (24, 21, 15) */,
  32'h3ea31756 /* (20, 21, 15) */,
  32'h3ecca1ac /* (16, 21, 15) */,
  32'h3ea31756 /* (12, 21, 15) */,
  32'h3e2c9c6c /* (8, 21, 15) */,
  32'h3ddcf428 /* (4, 21, 15) */,
  32'h3dbe6d47 /* (0, 21, 15) */,
  32'h3e1fe07e /* (28, 17, 15) */,
  32'h3e803f85 /* (24, 17, 15) */,
  32'h3efaa119 /* (20, 17, 15) */,
  32'h3f2286f8 /* (16, 17, 15) */,
  32'h3efaa119 /* (12, 17, 15) */,
  32'h3e803f85 /* (8, 17, 15) */,
  32'h3e1fe07e /* (4, 17, 15) */,
  32'h3e086183 /* (0, 17, 15) */,
  32'h3e0ff4ce /* (28, 13, 15) */,
  32'h3e640ba2 /* (24, 13, 15) */,
  32'h3edb3822 /* (20, 13, 15) */,
  32'h3f0bd969 /* (16, 13, 15) */,
  32'h3edb3822 /* (12, 13, 15) */,
  32'h3e640ba2 /* (8, 13, 15) */,
  32'h3e0ff4ce /* (4, 13, 15) */,
  32'h3df6cc6d /* (0, 13, 15) */,
  32'h3da3c1ed /* (28, 9, 15) */,
  32'h3dfc30a3 /* (24, 9, 15) */,
  32'h3e6a25fd /* (20, 9, 15) */,
  32'h3e908107 /* (16, 9, 15) */,
  32'h3e6a25fd /* (12, 9, 15) */,
  32'h3dfc30a3 /* (8, 9, 15) */,
  32'h3da3c1ed /* (4, 9, 15) */,
  32'h3d8df2c1 /* (0, 9, 15) */,
  32'h3d4def9b /* (28, 5, 15) */,
  32'h3d9a5b6b /* (24, 5, 15) */,
  32'h3e0ae903 /* (20, 5, 15) */,
  32'h3e26bbbb /* (16, 5, 15) */,
  32'h3e0ae903 /* (12, 5, 15) */,
  32'h3d9a5b6b /* (8, 5, 15) */,
  32'h3d4def9b /* (4, 5, 15) */,
  32'h3d347f0a /* (0, 5, 15) */,
  32'h3d294c4b /* (28, 1, 15) */,
  32'h3d7a003f /* (24, 1, 15) */,
  32'h3ddd43c2 /* (20, 1, 15) */,
  32'h3e02e976 /* (16, 1, 15) */,
  32'h3ddd43c2 /* (12, 1, 15) */,
  32'h3d7a003f /* (8, 1, 15) */,
  32'h3d294c4b /* (4, 1, 15) */,
  32'h3d155505 /* (0, 1, 15) */,
  32'h3d25fa09 /* (28, 29, 11) */,
  32'h3d5d0a38 /* (24, 29, 11) */,
  32'h3db0b965 /* (20, 29, 11) */,
  32'h3dc1602b /* (16, 29, 11) */,
  32'h3db0b965 /* (12, 29, 11) */,
  32'h3d5d0a38 /* (8, 29, 11) */,
  32'h3d25fa09 /* (4, 29, 11) */,
  32'h3d198ce9 /* (0, 29, 11) */,
  32'h3d52976b /* (28, 25, 11) */,
  32'h3d941bce /* (24, 25, 11) */,
  32'h3df94537 /* (20, 25, 11) */,
  32'h3e0d9cf0 /* (16, 25, 11) */,
  32'h3df94537 /* (12, 25, 11) */,
  32'h3d941bce /* (8, 25, 11) */,
  32'h3d52976b /* (4, 25, 11) */,
  32'h3d3dcd22 /* (0, 25, 11) */,
  32'h3da66ad4 /* (28, 21, 11) */,
  32'h3df84bb3 /* (24, 21, 11) */,
  32'h3e5e44ac /* (20, 21, 11) */,
  32'h3e84c8e0 /* (16, 21, 11) */,
  32'h3e5e44ac /* (12, 21, 11) */,
  32'h3df84bb3 /* (8, 21, 11) */,
  32'h3da66ad4 /* (4, 21, 11) */,
  32'h3d922642 /* (0, 21, 11) */,
  32'h3ddcf428 /* (28, 17, 11) */,
  32'h3e2c9c6c /* (24, 17, 11) */,
  32'h3ea31756 /* (20, 17, 11) */,
  32'h3ecca1ac /* (16, 17, 11) */,
  32'h3ea31756 /* (12, 17, 11) */,
  32'h3e2c9c6c /* (8, 17, 11) */,
  32'h3ddcf428 /* (4, 17, 11) */,
  32'h3dbe6d47 /* (0, 17, 11) */,
  32'h3dcf13a3 /* (28, 13, 11) */,
  32'h3e1e607d /* (24, 13, 11) */,
  32'h3e91dfe2 /* (20, 13, 11) */,
  32'h3eb2bd2a /* (16, 13, 11) */,
  32'h3e91dfe2 /* (12, 13, 11) */,
  32'h3e1e607d /* (8, 13, 11) */,
  32'h3dcf13a3 /* (4, 13, 11) */,
  32'h3db3fd83 /* (0, 13, 11) */,
  32'h3d81d711 /* (28, 9, 11) */,
  32'h3dbc4d73 /* (24, 9, 11) */,
  32'h3e23781b /* (20, 9, 11) */,
  32'h3e3e5da7 /* (16, 9, 11) */,
  32'h3e23781b /* (12, 9, 11) */,
  32'h3dbc4d73 /* (8, 9, 11) */,
  32'h3d81d711 /* (4, 9, 11) */,
  32'h3d66dac1 /* (0, 9, 11) */,
  32'h3d358341 /* (28, 5, 11) */,
  32'h3d77c8fd /* (24, 5, 11) */,
  32'h3dca9d53 /* (20, 5, 11) */,
  32'h3de14ffa /* (16, 5, 11) */,
  32'h3dca9d53 /* (12, 5, 11) */,
  32'h3d77c8fd /* (8, 5, 11) */,
  32'h3d358341 /* (4, 5, 11) */,
  32'h3d25e815 /* (0, 5, 11) */,
  32'h3d1f5dc3 /* (28, 1, 11) */,
  32'h3d513c3d /* (24, 1, 11) */,
  32'h3da53628 /* (20, 1, 11) */,
  32'h3db336e0 /* (16, 1, 11) */,
  32'h3da53628 /* (12, 1, 11) */,
  32'h3d513c3d /* (8, 1, 11) */,
  32'h3d1f5dc3 /* (4, 1, 11) */,
  32'h3d147e90 /* (0, 1, 11) */,
  32'h3d155fa4 /* (28, 29, 7) */,
  32'h3d2054cd /* (24, 29, 7) */,
  32'h3d5ab0e1 /* (20, 29, 7) */,
  32'h3d58de26 /* (16, 29, 7) */,
  32'h3d5ab0e1 /* (12, 29, 7) */,
  32'h3d2054cd /* (8, 29, 7) */,
  32'h3d155fa4 /* (4, 29, 7) */,
  32'h3d1cfd70 /* (0, 29, 7) */,
  32'h3d1cbb18 /* (28, 25, 7) */,
  32'h3d432bf1 /* (24, 25, 7) */,
  32'h3d938890 /* (20, 25, 7) */,
  32'h3d9b7830 /* (16, 25, 7) */,
  32'h3d938890 /* (12, 25, 7) */,
  32'h3d432bf1 /* (8, 25, 7) */,
  32'h3d1cbb18 /* (4, 25, 7) */,
  32'h3d162f74 /* (0, 25, 7) */,
  32'h3d52976b /* (28, 21, 7) */,
  32'h3d941bce /* (24, 21, 7) */,
  32'h3df94537 /* (20, 21, 7) */,
  32'h3e0d9cf0 /* (16, 21, 7) */,
  32'h3df94537 /* (12, 21, 7) */,
  32'h3d941bce /* (8, 21, 7) */,
  32'h3d52976b /* (4, 21, 7) */,
  32'h3d3dcd22 /* (0, 21, 7) */,
  32'h3d7b9f11 /* (28, 17, 7) */,
  32'h3dbf0444 /* (24, 17, 7) */,
  32'h3e2e6a71 /* (20, 17, 7) */,
  32'h3e540b9b /* (16, 17, 7) */,
  32'h3e2e6a71 /* (12, 17, 7) */,
  32'h3dbf0444 /* (8, 17, 7) */,
  32'h3d7b9f11 /* (4, 17, 7) */,
  32'h3d5b6048 /* (0, 17, 7) */,
  32'h3d770afc /* (28, 13, 7) */,
  32'h3db56072 /* (24, 13, 7) */,
  32'h3e1f8cbf /* (20, 13, 7) */,
  32'h3e3bd4ee /* (16, 13, 7) */,
  32'h3e1f8cbf /* (12, 13, 7) */,
  32'h3db56072 /* (8, 13, 7) */,
  32'h3d770afc /* (4, 13, 7) */,
  32'h3d5a6fdd /* (0, 13, 7) */,
  32'h3d30de15 /* (28, 9, 7) */,
  32'h3d6b8b35 /* (24, 9, 7) */,
  32'h3dbc51f9 /* (20, 9, 7) */,
  32'h3dce1075 /* (16, 9, 7) */,
  32'h3dbc51f9 /* (12, 9, 7) */,
  32'h3d6b8b35 /* (8, 9, 7) */,
  32'h3d30de15 /* (4, 9, 7) */,
  32'h3d23a039 /* (0, 9, 7) */,
  32'h3d1508af /* (28, 5, 7) */,
  32'h3d2bff3e /* (24, 5, 7) */,
  32'h3d75e4d4 /* (20, 5, 7) */,
  32'h3d7a662c /* (16, 5, 7) */,
  32'h3d75e4d4 /* (12, 5, 7) */,
  32'h3d2bff3e /* (8, 5, 7) */,
  32'h3d1508af /* (4, 5, 7) */,
  32'h3d154f7b /* (0, 5, 7) */,
  32'h3d17ff6b /* (28, 1, 7) */,
  32'h3d1bb8b6 /* (24, 1, 7) */,
  32'h3d4ea8e5 /* (20, 1, 7) */,
  32'h3d49f75a /* (16, 1, 7) */,
  32'h3d4ea8e5 /* (12, 1, 7) */,
  32'h3d1bb8b6 /* (8, 1, 7) */,
  32'h3d17ff6b /* (4, 1, 7) */,
  32'h3d25463b /* (0, 1, 7) */,
  32'h3d4920d0 /* (28, 29, 3) */,
  32'h3d1392fe /* (24, 29, 3) */,
  32'h3d28b308 /* (20, 29, 3) */,
  32'h3d19c07a /* (16, 29, 3) */,
  32'h3d28b308 /* (12, 29, 3) */,
  32'h3d1392fe /* (8, 29, 3) */,
  32'h3d4920d0 /* (4, 29, 3) */,
  32'h3d9c797c /* (0, 29, 3) */,
  32'h3d155fa4 /* (28, 25, 3) */,
  32'h3d2054cd /* (24, 25, 3) */,
  32'h3d5ab0e1 /* (20, 25, 3) */,
  32'h3d58de26 /* (16, 25, 3) */,
  32'h3d5ab0e1 /* (12, 25, 3) */,
  32'h3d2054cd /* (8, 25, 3) */,
  32'h3d155fa4 /* (4, 25, 3) */,
  32'h3d1cfd70 /* (0, 25, 3) */,
  32'h3d25fa09 /* (28, 21, 3) */,
  32'h3d5d0a38 /* (24, 21, 3) */,
  32'h3db0b965 /* (20, 21, 3) */,
  32'h3dc1602b /* (16, 21, 3) */,
  32'h3db0b965 /* (12, 21, 3) */,
  32'h3d5d0a38 /* (8, 21, 3) */,
  32'h3d25fa09 /* (4, 21, 3) */,
  32'h3d198ce9 /* (0, 21, 3) */,
  32'h3d349293 /* (28, 17, 3) */,
  32'h3d8608f0 /* (24, 17, 3) */,
  32'h3deea44d /* (20, 17, 3) */,
  32'h3e0de417 /* (16, 17, 3) */,
  32'h3deea44d /* (12, 17, 3) */,
  32'h3d8608f0 /* (8, 17, 3) */,
  32'h3d349293 /* (4, 17, 3) */,
  32'h3d1eeabe /* (0, 17, 3) */,
  32'h3d385879 /* (28, 13, 3) */,
  32'h3d82c188 /* (24, 13, 3) */,
  32'h3dddef48 /* (20, 13, 3) */,
  32'h3dfdd31f /* (16, 13, 3) */,
  32'h3dddef48 /* (12, 13, 3) */,
  32'h3d82c188 /* (8, 13, 3) */,
  32'h3d385879 /* (4, 13, 3) */,
  32'h3d258110 /* (0, 13, 3) */,
  32'h3d16b5b2 /* (28, 9, 3) */,
  32'h3d37919e /* (24, 9, 3) */,
  32'h3d886b82 /* (20, 9, 3) */,
  32'h3d8e3848 /* (16, 9, 3) */,
  32'h3d886b82 /* (12, 9, 3) */,
  32'h3d37919e /* (8, 9, 3) */,
  32'h3d16b5b2 /* (4, 9, 3) */,
  32'h3d1237a7 /* (0, 9, 3) */,
  32'h3d25f5ce /* (28, 5, 3) */,
  32'h3d15d660 /* (24, 5, 3) */,
  32'h3d3a4ebb /* (20, 5, 3) */,
  32'h3d3046d8 /* (16, 5, 3) */,
  32'h3d3a4ebb /* (12, 5, 3) */,
  32'h3d15d660 /* (8, 5, 3) */,
  32'h3d25f5ce /* (4, 5, 3) */,
  32'h3d490b0e /* (0, 5, 3) */,
  32'h3d6eb36b /* (28, 1, 3) */,
  32'h3d146963 /* (24, 1, 3) */,
  32'h3d210eee /* (20, 1, 3) */,
  32'h3d0fbc59 /* (16, 1, 3) */,
  32'h3d210eee /* (12, 1, 3) */,
  32'h3d146963 /* (8, 1, 3) */,
  32'h3d6eb36b /* (4, 1, 3) */,
  32'h3dff9e3f /* (0, 1, 3) */,
  32'h3d9c757b /* (31, 28, 31) */,
  32'h3d334ee4 /* (27, 28, 31) */,
  32'h3d13f199 /* (23, 28, 31) */,
  32'h3d2e802a /* (19, 28, 31) */,
  32'h3d294c4b /* (15, 28, 31) */,
  32'h3d1f5dc3 /* (11, 28, 31) */,
  32'h3d17ff6b /* (7, 28, 31) */,
  32'h3d6eb36b /* (3, 28, 31) */,
  32'h3d1704d7 /* (31, 24, 31) */,
  32'h3d1412fd /* (27, 24, 31) */,
  32'h3d2fba80 /* (23, 24, 31) */,
  32'h3d7573b6 /* (19, 24, 31) */,
  32'h3d7a003f /* (15, 24, 31) */,
  32'h3d513c3d /* (11, 24, 31) */,
  32'h3d1bb8b6 /* (7, 24, 31) */,
  32'h3d146963 /* (3, 24, 31) */,
  32'h3d1a2df1 /* (31, 20, 31) */,
  32'h3d310ad3 /* (27, 20, 31) */,
  32'h3d803124 /* (23, 20, 31) */,
  32'h3dce8d02 /* (19, 20, 31) */,
  32'h3ddd43c2 /* (15, 20, 31) */,
  32'h3da53628 /* (11, 20, 31) */,
  32'h3d4ea8e5 /* (7, 20, 31) */,
  32'h3d210eee /* (3, 20, 31) */,
  32'h3d067e68 /* (31, 16, 31) */,
  32'h3d24852f /* (27, 16, 31) */,
  32'h3d8420c9 /* (23, 16, 31) */,
  32'h3deaafef /* (19, 16, 31) */,
  32'h3e02e976 /* (15, 16, 31) */,
  32'h3db336e0 /* (11, 16, 31) */,
  32'h3d49f75a /* (7, 16, 31) */,
  32'h3d0fbc59 /* (3, 16, 31) */,
  32'h3d1a2df1 /* (31, 12, 31) */,
  32'h3d310ad3 /* (27, 12, 31) */,
  32'h3d803124 /* (23, 12, 31) */,
  32'h3dce8d02 /* (19, 12, 31) */,
  32'h3ddd43c2 /* (15, 12, 31) */,
  32'h3da53628 /* (11, 12, 31) */,
  32'h3d4ea8e5 /* (7, 12, 31) */,
  32'h3d210eee /* (3, 12, 31) */,
  32'h3d1704d7 /* (31, 8, 31) */,
  32'h3d1412fd /* (27, 8, 31) */,
  32'h3d2fba80 /* (23, 8, 31) */,
  32'h3d7573b6 /* (19, 8, 31) */,
  32'h3d7a003f /* (15, 8, 31) */,
  32'h3d513c3d /* (11, 8, 31) */,
  32'h3d1bb8b6 /* (7, 8, 31) */,
  32'h3d146963 /* (3, 8, 31) */,
  32'h3d9c757b /* (31, 4, 31) */,
  32'h3d334ee4 /* (27, 4, 31) */,
  32'h3d13f199 /* (23, 4, 31) */,
  32'h3d2e802a /* (19, 4, 31) */,
  32'h3d294c4b /* (15, 4, 31) */,
  32'h3d1f5dc3 /* (11, 4, 31) */,
  32'h3d17ff6b /* (7, 4, 31) */,
  32'h3d6eb36b /* (3, 4, 31) */,
  32'h3f10fe39 /* (31, 0, 31) */,
  32'h3d6e9998 /* (27, 0, 31) */,
  32'h3d11a5c6 /* (23, 0, 31) */,
  32'h3d1d4601 /* (19, 0, 31) */,
  32'h3d155505 /* (15, 0, 31) */,
  32'h3d147e90 /* (11, 0, 31) */,
  32'h3d25463b /* (7, 0, 31) */,
  32'h3dff9e3f /* (3, 0, 31) */,
  32'h3d334ee4 /* (31, 28, 27) */,
  32'h3d189061 /* (27, 28, 27) */,
  32'h3d1ee50b /* (23, 28, 27) */,
  32'h3d4ea6a0 /* (19, 28, 27) */,
  32'h3d4def9b /* (15, 28, 27) */,
  32'h3d358341 /* (11, 28, 27) */,
  32'h3d1508af /* (7, 28, 27) */,
  32'h3d25f5ce /* (3, 28, 27) */,
  32'h3d1412fd /* (31, 24, 27) */,
  32'h3d1c4d38 /* (27, 24, 27) */,
  32'h3d49c96c /* (23, 24, 27) */,
  32'h3d94d380 /* (19, 24, 27) */,
  32'h3d9a5b6b /* (15, 24, 27) */,
  32'h3d77c8fd /* (11, 24, 27) */,
  32'h3d2bff3e /* (7, 24, 27) */,
  32'h3d15d660 /* (3, 24, 27) */,
  32'h3d310ad3 /* (31, 20, 27) */,
  32'h3d4f6dfc /* (27, 20, 27) */,
  32'h3d9af1c2 /* (23, 20, 27) */,
  32'h3e00477d /* (19, 20, 27) */,
  32'h3e0ae903 /* (15, 20, 27) */,
  32'h3dca9d53 /* (11, 20, 27) */,
  32'h3d75e4d4 /* (7, 20, 27) */,
  32'h3d3a4ebb /* (3, 20, 27) */,
  32'h3d24852f /* (31, 16, 27) */,
  32'h3d4ab7f7 /* (27, 16, 27) */,
  32'h3da4f2f4 /* (23, 16, 27) */,
  32'h3e1486b7 /* (19, 16, 27) */,
  32'h3e26bbbb /* (15, 16, 27) */,
  32'h3de14ffa /* (11, 16, 27) */,
  32'h3d7a662c /* (7, 16, 27) */,
  32'h3d3046d8 /* (3, 16, 27) */,
  32'h3d310ad3 /* (31, 12, 27) */,
  32'h3d4f6dfc /* (27, 12, 27) */,
  32'h3d9af1c2 /* (23, 12, 27) */,
  32'h3e00477d /* (19, 12, 27) */,
  32'h3e0ae903 /* (15, 12, 27) */,
  32'h3dca9d53 /* (11, 12, 27) */,
  32'h3d75e4d4 /* (7, 12, 27) */,
  32'h3d3a4ebb /* (3, 12, 27) */,
  32'h3d1412fd /* (31, 8, 27) */,
  32'h3d1c4d38 /* (27, 8, 27) */,
  32'h3d49c96c /* (23, 8, 27) */,
  32'h3d94d380 /* (19, 8, 27) */,
  32'h3d9a5b6b /* (15, 8, 27) */,
  32'h3d77c8fd /* (11, 8, 27) */,
  32'h3d2bff3e /* (7, 8, 27) */,
  32'h3d15d660 /* (3, 8, 27) */,
  32'h3d334ee4 /* (31, 4, 27) */,
  32'h3d189061 /* (27, 4, 27) */,
  32'h3d1ee50b /* (23, 4, 27) */,
  32'h3d4ea6a0 /* (19, 4, 27) */,
  32'h3d4def9b /* (15, 4, 27) */,
  32'h3d358341 /* (11, 4, 27) */,
  32'h3d1508af /* (7, 4, 27) */,
  32'h3d25f5ce /* (3, 4, 27) */,
  32'h3d6e9998 /* (31, 0, 27) */,
  32'h3d25e3da /* (27, 0, 27) */,
  32'h3d16a564 /* (23, 0, 27) */,
  32'h3d384488 /* (19, 0, 27) */,
  32'h3d347f0a /* (15, 0, 27) */,
  32'h3d25e815 /* (11, 0, 27) */,
  32'h3d154f7b /* (7, 0, 27) */,
  32'h3d490b0e /* (3, 0, 27) */,
  32'h3d13f199 /* (31, 28, 23) */,
  32'h3d1ee50b /* (27, 28, 23) */,
  32'h3d51a9d2 /* (23, 28, 23) */,
  32'h3d9d0afa /* (19, 28, 23) */,
  32'h3da3c1ed /* (15, 28, 23) */,
  32'h3d81d711 /* (11, 28, 23) */,
  32'h3d30de15 /* (7, 28, 23) */,
  32'h3d16b5b2 /* (3, 28, 23) */,
  32'h3d2fba80 /* (31, 24, 23) */,
  32'h3d49c96c /* (27, 24, 23) */,
  32'h3d921bde /* (23, 24, 23) */,
  32'h3deb6b6d /* (19, 24, 23) */,
  32'h3dfc30a3 /* (15, 24, 23) */,
  32'h3dbc4d73 /* (11, 24, 23) */,
  32'h3d6b8b35 /* (7, 24, 23) */,
  32'h3d37919e /* (3, 24, 23) */,
  32'h3d803124 /* (31, 20, 23) */,
  32'h3d9af1c2 /* (27, 20, 23) */,
  32'h3df3b4f2 /* (23, 20, 23) */,
  32'h3e53dc51 /* (19, 20, 23) */,
  32'h3e6a25fd /* (15, 20, 23) */,
  32'h3e23781b /* (11, 20, 23) */,
  32'h3dbc51f9 /* (7, 20, 23) */,
  32'h3d886b82 /* (3, 20, 23) */,
  32'h3d8420c9 /* (31, 16, 23) */,
  32'h3da4f2f4 /* (27, 16, 23) */,
  32'h3e0981d7 /* (23, 16, 23) */,
  32'h3e7e4b9d /* (19, 16, 23) */,
  32'h3e908107 /* (15, 16, 23) */,
  32'h3e3e5da7 /* (11, 16, 23) */,
  32'h3dce1075 /* (7, 16, 23) */,
  32'h3d8e3848 /* (3, 16, 23) */,
  32'h3d803124 /* (31, 12, 23) */,
  32'h3d9af1c2 /* (27, 12, 23) */,
  32'h3df3b4f2 /* (23, 12, 23) */,
  32'h3e53dc51 /* (19, 12, 23) */,
  32'h3e6a25fd /* (15, 12, 23) */,
  32'h3e23781b /* (11, 12, 23) */,
  32'h3dbc51f9 /* (7, 12, 23) */,
  32'h3d886b82 /* (3, 12, 23) */,
  32'h3d2fba80 /* (31, 8, 23) */,
  32'h3d49c96c /* (27, 8, 23) */,
  32'h3d921bde /* (23, 8, 23) */,
  32'h3deb6b6d /* (19, 8, 23) */,
  32'h3dfc30a3 /* (15, 8, 23) */,
  32'h3dbc4d73 /* (11, 8, 23) */,
  32'h3d6b8b35 /* (7, 8, 23) */,
  32'h3d37919e /* (3, 8, 23) */,
  32'h3d13f199 /* (31, 4, 23) */,
  32'h3d1ee50b /* (27, 4, 23) */,
  32'h3d51a9d2 /* (23, 4, 23) */,
  32'h3d9d0afa /* (19, 4, 23) */,
  32'h3da3c1ed /* (15, 4, 23) */,
  32'h3d81d711 /* (11, 4, 23) */,
  32'h3d30de15 /* (7, 4, 23) */,
  32'h3d16b5b2 /* (3, 4, 23) */,
  32'h3d11a5c6 /* (31, 0, 23) */,
  32'h3d16a564 /* (27, 0, 23) */,
  32'h3d3dc47d /* (23, 0, 23) */,
  32'h3d89a49e /* (19, 0, 23) */,
  32'h3d8df2c1 /* (15, 0, 23) */,
  32'h3d66dac1 /* (11, 0, 23) */,
  32'h3d23a039 /* (7, 0, 23) */,
  32'h3d1237a7 /* (3, 0, 23) */,
  32'h3d2e802a /* (31, 28, 19) */,
  32'h3d4ea6a0 /* (27, 28, 19) */,
  32'h3d9d0afa /* (23, 28, 19) */,
  32'h3e0415cb /* (19, 28, 19) */,
  32'h3e0ff4ce /* (15, 28, 19) */,
  32'h3dcf13a3 /* (11, 28, 19) */,
  32'h3d770afc /* (7, 28, 19) */,
  32'h3d385879 /* (3, 28, 19) */,
  32'h3d7573b6 /* (31, 24, 19) */,
  32'h3d94d380 /* (27, 24, 19) */,
  32'h3deb6b6d /* (23, 24, 19) */,
  32'h3e4dd3dc /* (19, 24, 19) */,
  32'h3e640ba2 /* (15, 24, 19) */,
  32'h3e1e607d /* (11, 24, 19) */,
  32'h3db56072 /* (7, 24, 19) */,
  32'h3d82c188 /* (3, 24, 19) */,
  32'h3dce8d02 /* (31, 20, 19) */,
  32'h3e00477d /* (27, 20, 19) */,
  32'h3e53dc51 /* (23, 20, 19) */,
  32'h3ec1d890 /* (19, 20, 19) */,
  32'h3edb3822 /* (15, 20, 19) */,
  32'h3e91dfe2 /* (11, 20, 19) */,
  32'h3e1f8cbf /* (7, 20, 19) */,
  32'h3dddef48 /* (3, 20, 19) */,
  32'h3deaafef /* (31, 16, 19) */,
  32'h3e1486b7 /* (27, 16, 19) */,
  32'h3e7e4b9d /* (23, 16, 19) */,
  32'h3ef27895 /* (19, 16, 19) */,
  32'h3f0bd969 /* (15, 16, 19) */,
  32'h3eb2bd2a /* (11, 16, 19) */,
  32'h3e3bd4ee /* (7, 16, 19) */,
  32'h3dfdd31f /* (3, 16, 19) */,
  32'h3dce8d02 /* (31, 12, 19) */,
  32'h3e00477d /* (27, 12, 19) */,
  32'h3e53dc51 /* (23, 12, 19) */,
  32'h3ec1d890 /* (19, 12, 19) */,
  32'h3edb3822 /* (15, 12, 19) */,
  32'h3e91dfe2 /* (11, 12, 19) */,
  32'h3e1f8cbf /* (7, 12, 19) */,
  32'h3dddef48 /* (3, 12, 19) */,
  32'h3d7573b6 /* (31, 8, 19) */,
  32'h3d94d380 /* (27, 8, 19) */,
  32'h3deb6b6d /* (23, 8, 19) */,
  32'h3e4dd3dc /* (19, 8, 19) */,
  32'h3e640ba2 /* (15, 8, 19) */,
  32'h3e1e607d /* (11, 8, 19) */,
  32'h3db56072 /* (7, 8, 19) */,
  32'h3d82c188 /* (3, 8, 19) */,
  32'h3d2e802a /* (31, 4, 19) */,
  32'h3d4ea6a0 /* (27, 4, 19) */,
  32'h3d9d0afa /* (23, 4, 19) */,
  32'h3e0415cb /* (19, 4, 19) */,
  32'h3e0ff4ce /* (15, 4, 19) */,
  32'h3dcf13a3 /* (11, 4, 19) */,
  32'h3d770afc /* (7, 4, 19) */,
  32'h3d385879 /* (3, 4, 19) */,
  32'h3d1d4601 /* (31, 0, 19) */,
  32'h3d384488 /* (27, 0, 19) */,
  32'h3d89a49e /* (23, 0, 19) */,
  32'h3de3e928 /* (19, 0, 19) */,
  32'h3df6cc6d /* (15, 0, 19) */,
  32'h3db3fd83 /* (11, 0, 19) */,
  32'h3d5a6fdd /* (7, 0, 19) */,
  32'h3d258110 /* (3, 0, 19) */,
  32'h3d294c4b /* (31, 28, 15) */,
  32'h3d4def9b /* (27, 28, 15) */,
  32'h3da3c1ed /* (23, 28, 15) */,
  32'h3e0ff4ce /* (19, 28, 15) */,
  32'h3e1fe07e /* (15, 28, 15) */,
  32'h3ddcf428 /* (11, 28, 15) */,
  32'h3d7b9f11 /* (7, 28, 15) */,
  32'h3d349293 /* (3, 28, 15) */,
  32'h3d7a003f /* (31, 24, 15) */,
  32'h3d9a5b6b /* (27, 24, 15) */,
  32'h3dfc30a3 /* (23, 24, 15) */,
  32'h3e640ba2 /* (19, 24, 15) */,
  32'h3e803f85 /* (15, 24, 15) */,
  32'h3e2c9c6c /* (11, 24, 15) */,
  32'h3dbf0444 /* (7, 24, 15) */,
  32'h3d8608f0 /* (3, 24, 15) */,
  32'h3ddd43c2 /* (31, 20, 15) */,
  32'h3e0ae903 /* (27, 20, 15) */,
  32'h3e6a25fd /* (23, 20, 15) */,
  32'h3edb3822 /* (19, 20, 15) */,
  32'h3efaa119 /* (15, 20, 15) */,
  32'h3ea31756 /* (11, 20, 15) */,
  32'h3e2e6a71 /* (7, 20, 15) */,
  32'h3deea44d /* (3, 20, 15) */,
  32'h3e02e976 /* (31, 16, 15) */,
  32'h3e26bbbb /* (27, 16, 15) */,
  32'h3e908107 /* (23, 16, 15) */,
  32'h3f0bd969 /* (19, 16, 15) */,
  32'h3f2286f8 /* (15, 16, 15) */,
  32'h3ecca1ac /* (11, 16, 15) */,
  32'h3e540b9b /* (7, 16, 15) */,
  32'h3e0de417 /* (3, 16, 15) */,
  32'h3ddd43c2 /* (31, 12, 15) */,
  32'h3e0ae903 /* (27, 12, 15) */,
  32'h3e6a25fd /* (23, 12, 15) */,
  32'h3edb3822 /* (19, 12, 15) */,
  32'h3efaa119 /* (15, 12, 15) */,
  32'h3ea31756 /* (11, 12, 15) */,
  32'h3e2e6a71 /* (7, 12, 15) */,
  32'h3deea44d /* (3, 12, 15) */,
  32'h3d7a003f /* (31, 8, 15) */,
  32'h3d9a5b6b /* (27, 8, 15) */,
  32'h3dfc30a3 /* (23, 8, 15) */,
  32'h3e640ba2 /* (19, 8, 15) */,
  32'h3e803f85 /* (15, 8, 15) */,
  32'h3e2c9c6c /* (11, 8, 15) */,
  32'h3dbf0444 /* (7, 8, 15) */,
  32'h3d8608f0 /* (3, 8, 15) */,
  32'h3d294c4b /* (31, 4, 15) */,
  32'h3d4def9b /* (27, 4, 15) */,
  32'h3da3c1ed /* (23, 4, 15) */,
  32'h3e0ff4ce /* (19, 4, 15) */,
  32'h3e1fe07e /* (15, 4, 15) */,
  32'h3ddcf428 /* (11, 4, 15) */,
  32'h3d7b9f11 /* (7, 4, 15) */,
  32'h3d349293 /* (3, 4, 15) */,
  32'h3d155505 /* (31, 0, 15) */,
  32'h3d347f0a /* (27, 0, 15) */,
  32'h3d8df2c1 /* (23, 0, 15) */,
  32'h3df6cc6d /* (19, 0, 15) */,
  32'h3e086183 /* (15, 0, 15) */,
  32'h3dbe6d47 /* (11, 0, 15) */,
  32'h3d5b6048 /* (7, 0, 15) */,
  32'h3d1eeabe /* (3, 0, 15) */,
  32'h3d1f5dc3 /* (31, 28, 11) */,
  32'h3d358341 /* (27, 28, 11) */,
  32'h3d81d711 /* (23, 28, 11) */,
  32'h3dcf13a3 /* (19, 28, 11) */,
  32'h3ddcf428 /* (15, 28, 11) */,
  32'h3da66ad4 /* (11, 28, 11) */,
  32'h3d52976b /* (7, 28, 11) */,
  32'h3d25fa09 /* (3, 28, 11) */,
  32'h3d513c3d /* (31, 24, 11) */,
  32'h3d77c8fd /* (27, 24, 11) */,
  32'h3dbc4d73 /* (23, 24, 11) */,
  32'h3e1e607d /* (19, 24, 11) */,
  32'h3e2c9c6c /* (15, 24, 11) */,
  32'h3df84bb3 /* (11, 24, 11) */,
  32'h3d941bce /* (7, 24, 11) */,
  32'h3d5d0a38 /* (3, 24, 11) */,
  32'h3da53628 /* (31, 20, 11) */,
  32'h3dca9d53 /* (27, 20, 11) */,
  32'h3e23781b /* (23, 20, 11) */,
  32'h3e91dfe2 /* (19, 20, 11) */,
  32'h3ea31756 /* (15, 20, 11) */,
  32'h3e5e44ac /* (11, 20, 11) */,
  32'h3df94537 /* (7, 20, 11) */,
  32'h3db0b965 /* (3, 20, 11) */,
  32'h3db336e0 /* (31, 16, 11) */,
  32'h3de14ffa /* (27, 16, 11) */,
  32'h3e3e5da7 /* (23, 16, 11) */,
  32'h3eb2bd2a /* (19, 16, 11) */,
  32'h3ecca1ac /* (15, 16, 11) */,
  32'h3e84c8e0 /* (11, 16, 11) */,
  32'h3e0d9cf0 /* (7, 16, 11) */,
  32'h3dc1602b /* (3, 16, 11) */,
  32'h3da53628 /* (31, 12, 11) */,
  32'h3dca9d53 /* (27, 12, 11) */,
  32'h3e23781b /* (23, 12, 11) */,
  32'h3e91dfe2 /* (19, 12, 11) */,
  32'h3ea31756 /* (15, 12, 11) */,
  32'h3e5e44ac /* (11, 12, 11) */,
  32'h3df94537 /* (7, 12, 11) */,
  32'h3db0b965 /* (3, 12, 11) */,
  32'h3d513c3d /* (31, 8, 11) */,
  32'h3d77c8fd /* (27, 8, 11) */,
  32'h3dbc4d73 /* (23, 8, 11) */,
  32'h3e1e607d /* (19, 8, 11) */,
  32'h3e2c9c6c /* (15, 8, 11) */,
  32'h3df84bb3 /* (11, 8, 11) */,
  32'h3d941bce /* (7, 8, 11) */,
  32'h3d5d0a38 /* (3, 8, 11) */,
  32'h3d1f5dc3 /* (31, 4, 11) */,
  32'h3d358341 /* (27, 4, 11) */,
  32'h3d81d711 /* (23, 4, 11) */,
  32'h3dcf13a3 /* (19, 4, 11) */,
  32'h3ddcf428 /* (15, 4, 11) */,
  32'h3da66ad4 /* (11, 4, 11) */,
  32'h3d52976b /* (7, 4, 11) */,
  32'h3d25fa09 /* (3, 4, 11) */,
  32'h3d147e90 /* (31, 0, 11) */,
  32'h3d25e815 /* (27, 0, 11) */,
  32'h3d66dac1 /* (23, 0, 11) */,
  32'h3db3fd83 /* (19, 0, 11) */,
  32'h3dbe6d47 /* (15, 0, 11) */,
  32'h3d922642 /* (11, 0, 11) */,
  32'h3d3dcd22 /* (7, 0, 11) */,
  32'h3d198ce9 /* (3, 0, 11) */,
  32'h3d17ff6b /* (31, 28, 7) */,
  32'h3d1508af /* (27, 28, 7) */,
  32'h3d30de15 /* (23, 28, 7) */,
  32'h3d770afc /* (19, 28, 7) */,
  32'h3d7b9f11 /* (15, 28, 7) */,
  32'h3d52976b /* (11, 28, 7) */,
  32'h3d1cbb18 /* (7, 28, 7) */,
  32'h3d155fa4 /* (3, 28, 7) */,
  32'h3d1bb8b6 /* (31, 24, 7) */,
  32'h3d2bff3e /* (27, 24, 7) */,
  32'h3d6b8b35 /* (23, 24, 7) */,
  32'h3db56072 /* (19, 24, 7) */,
  32'h3dbf0444 /* (15, 24, 7) */,
  32'h3d941bce /* (11, 24, 7) */,
  32'h3d432bf1 /* (7, 24, 7) */,
  32'h3d2054cd /* (3, 24, 7) */,
  32'h3d4ea8e5 /* (31, 20, 7) */,
  32'h3d75e4d4 /* (27, 20, 7) */,
  32'h3dbc51f9 /* (23, 20, 7) */,
  32'h3e1f8cbf /* (19, 20, 7) */,
  32'h3e2e6a71 /* (15, 20, 7) */,
  32'h3df94537 /* (11, 20, 7) */,
  32'h3d938890 /* (7, 20, 7) */,
  32'h3d5ab0e1 /* (3, 20, 7) */,
  32'h3d49f75a /* (31, 16, 7) */,
  32'h3d7a662c /* (27, 16, 7) */,
  32'h3dce1075 /* (23, 16, 7) */,
  32'h3e3bd4ee /* (19, 16, 7) */,
  32'h3e540b9b /* (15, 16, 7) */,
  32'h3e0d9cf0 /* (11, 16, 7) */,
  32'h3d9b7830 /* (7, 16, 7) */,
  32'h3d58de26 /* (3, 16, 7) */,
  32'h3d4ea8e5 /* (31, 12, 7) */,
  32'h3d75e4d4 /* (27, 12, 7) */,
  32'h3dbc51f9 /* (23, 12, 7) */,
  32'h3e1f8cbf /* (19, 12, 7) */,
  32'h3e2e6a71 /* (15, 12, 7) */,
  32'h3df94537 /* (11, 12, 7) */,
  32'h3d938890 /* (7, 12, 7) */,
  32'h3d5ab0e1 /* (3, 12, 7) */,
  32'h3d1bb8b6 /* (31, 8, 7) */,
  32'h3d2bff3e /* (27, 8, 7) */,
  32'h3d6b8b35 /* (23, 8, 7) */,
  32'h3db56072 /* (19, 8, 7) */,
  32'h3dbf0444 /* (15, 8, 7) */,
  32'h3d941bce /* (11, 8, 7) */,
  32'h3d432bf1 /* (7, 8, 7) */,
  32'h3d2054cd /* (3, 8, 7) */,
  32'h3d17ff6b /* (31, 4, 7) */,
  32'h3d1508af /* (27, 4, 7) */,
  32'h3d30de15 /* (23, 4, 7) */,
  32'h3d770afc /* (19, 4, 7) */,
  32'h3d7b9f11 /* (15, 4, 7) */,
  32'h3d52976b /* (11, 4, 7) */,
  32'h3d1cbb18 /* (7, 4, 7) */,
  32'h3d155fa4 /* (3, 4, 7) */,
  32'h3d25463b /* (31, 0, 7) */,
  32'h3d154f7b /* (27, 0, 7) */,
  32'h3d23a039 /* (23, 0, 7) */,
  32'h3d5a6fdd /* (19, 0, 7) */,
  32'h3d5b6048 /* (15, 0, 7) */,
  32'h3d3dcd22 /* (11, 0, 7) */,
  32'h3d162f74 /* (7, 0, 7) */,
  32'h3d1cfd70 /* (3, 0, 7) */,
  32'h3d6eb36b /* (31, 28, 3) */,
  32'h3d25f5ce /* (27, 28, 3) */,
  32'h3d16b5b2 /* (23, 28, 3) */,
  32'h3d385879 /* (19, 28, 3) */,
  32'h3d349293 /* (15, 28, 3) */,
  32'h3d25fa09 /* (11, 28, 3) */,
  32'h3d155fa4 /* (7, 28, 3) */,
  32'h3d4920d0 /* (3, 28, 3) */,
  32'h3d146963 /* (31, 24, 3) */,
  32'h3d15d660 /* (27, 24, 3) */,
  32'h3d37919e /* (23, 24, 3) */,
  32'h3d82c188 /* (19, 24, 3) */,
  32'h3d8608f0 /* (15, 24, 3) */,
  32'h3d5d0a38 /* (11, 24, 3) */,
  32'h3d2054cd /* (7, 24, 3) */,
  32'h3d1392fe /* (3, 24, 3) */,
  32'h3d210eee /* (31, 20, 3) */,
  32'h3d3a4ebb /* (27, 20, 3) */,
  32'h3d886b82 /* (23, 20, 3) */,
  32'h3dddef48 /* (19, 20, 3) */,
  32'h3deea44d /* (15, 20, 3) */,
  32'h3db0b965 /* (11, 20, 3) */,
  32'h3d5ab0e1 /* (7, 20, 3) */,
  32'h3d28b308 /* (3, 20, 3) */,
  32'h3d0fbc59 /* (31, 16, 3) */,
  32'h3d3046d8 /* (27, 16, 3) */,
  32'h3d8e3848 /* (23, 16, 3) */,
  32'h3dfdd31f /* (19, 16, 3) */,
  32'h3e0de417 /* (15, 16, 3) */,
  32'h3dc1602b /* (11, 16, 3) */,
  32'h3d58de26 /* (7, 16, 3) */,
  32'h3d19c07a /* (3, 16, 3) */,
  32'h3d210eee /* (31, 12, 3) */,
  32'h3d3a4ebb /* (27, 12, 3) */,
  32'h3d886b82 /* (23, 12, 3) */,
  32'h3dddef48 /* (19, 12, 3) */,
  32'h3deea44d /* (15, 12, 3) */,
  32'h3db0b965 /* (11, 12, 3) */,
  32'h3d5ab0e1 /* (7, 12, 3) */,
  32'h3d28b308 /* (3, 12, 3) */,
  32'h3d146963 /* (31, 8, 3) */,
  32'h3d15d660 /* (27, 8, 3) */,
  32'h3d37919e /* (23, 8, 3) */,
  32'h3d82c188 /* (19, 8, 3) */,
  32'h3d8608f0 /* (15, 8, 3) */,
  32'h3d5d0a38 /* (11, 8, 3) */,
  32'h3d2054cd /* (7, 8, 3) */,
  32'h3d1392fe /* (3, 8, 3) */,
  32'h3d6eb36b /* (31, 4, 3) */,
  32'h3d25f5ce /* (27, 4, 3) */,
  32'h3d16b5b2 /* (23, 4, 3) */,
  32'h3d385879 /* (19, 4, 3) */,
  32'h3d349293 /* (15, 4, 3) */,
  32'h3d25fa09 /* (11, 4, 3) */,
  32'h3d155fa4 /* (7, 4, 3) */,
  32'h3d4920d0 /* (3, 4, 3) */,
  32'h3dff9e3f /* (31, 0, 3) */,
  32'h3d490b0e /* (27, 0, 3) */,
  32'h3d1237a7 /* (23, 0, 3) */,
  32'h3d258110 /* (19, 0, 3) */,
  32'h3d1eeabe /* (15, 0, 3) */,
  32'h3d198ce9 /* (11, 0, 3) */,
  32'h3d1cfd70 /* (7, 0, 3) */,
  32'h3d9c797c /* (3, 0, 3) */,
  32'h3d8b1391 /* (30, 28, 31) */,
  32'h3d222a9c /* (26, 28, 31) */,
  32'h3d1839e3 /* (22, 28, 31) */,
  32'h3d303352 /* (18, 28, 31) */,
  32'h3d303352 /* (14, 28, 31) */,
  32'h3d1839e3 /* (10, 28, 31) */,
  32'h3d222a9c /* (6, 28, 31) */,
  32'h3d8b1391 /* (2, 28, 31) */,
  32'h3d15ce12 /* (30, 24, 31) */,
  32'h3d169650 /* (26, 24, 31) */,
  32'h3d3f0366 /* (22, 24, 31) */,
  32'h3d7e759f /* (18, 24, 31) */,
  32'h3d7e759f /* (14, 24, 31) */,
  32'h3d3f0366 /* (10, 24, 31) */,
  32'h3d169650 /* (6, 24, 31) */,
  32'h3d15ce12 /* (2, 24, 31) */,
  32'h3d1cac31 /* (30, 20, 31) */,
  32'h3d3dc5f0 /* (26, 20, 31) */,
  32'h3d91435f /* (22, 20, 31) */,
  32'h3ddbed5a /* (18, 20, 31) */,
  32'h3ddbed5a /* (14, 20, 31) */,
  32'h3d91435f /* (10, 20, 31) */,
  32'h3d3dc5f0 /* (6, 20, 31) */,
  32'h3d1cac31 /* (2, 20, 31) */,
  32'h3d09dfab /* (30, 16, 31) */,
  32'h3d34b66a /* (26, 16, 31) */,
  32'h3d99ac24 /* (22, 16, 31) */,
  32'h3dff32bb /* (18, 16, 31) */,
  32'h3dff32bb /* (14, 16, 31) */,
  32'h3d99ac24 /* (10, 16, 31) */,
  32'h3d34b66a /* (6, 16, 31) */,
  32'h3d09dfab /* (2, 16, 31) */,
  32'h3d1cac31 /* (30, 12, 31) */,
  32'h3d3dc5f0 /* (26, 12, 31) */,
  32'h3d91435f /* (22, 12, 31) */,
  32'h3ddbed5a /* (18, 12, 31) */,
  32'h3ddbed5a /* (14, 12, 31) */,
  32'h3d91435f /* (10, 12, 31) */,
  32'h3d3dc5f0 /* (6, 12, 31) */,
  32'h3d1cac31 /* (2, 12, 31) */,
  32'h3d15ce12 /* (30, 8, 31) */,
  32'h3d169650 /* (26, 8, 31) */,
  32'h3d3f0366 /* (22, 8, 31) */,
  32'h3d7e759f /* (18, 8, 31) */,
  32'h3d7e759f /* (14, 8, 31) */,
  32'h3d3f0366 /* (10, 8, 31) */,
  32'h3d169650 /* (6, 8, 31) */,
  32'h3d15ce12 /* (2, 8, 31) */,
  32'h3d8b1391 /* (30, 4, 31) */,
  32'h3d222a9c /* (26, 4, 31) */,
  32'h3d1839e3 /* (22, 4, 31) */,
  32'h3d303352 /* (18, 4, 31) */,
  32'h3d303352 /* (14, 4, 31) */,
  32'h3d1839e3 /* (10, 4, 31) */,
  32'h3d222a9c /* (6, 4, 31) */,
  32'h3d8b1391 /* (2, 4, 31) */,
  32'h3e709592 /* (30, 0, 31) */,
  32'h3d3f59b8 /* (26, 0, 31) */,
  32'h3d1142bb /* (22, 0, 31) */,
  32'h3d1ceee6 /* (18, 0, 31) */,
  32'h3d1ceee6 /* (14, 0, 31) */,
  32'h3d1142bb /* (10, 0, 31) */,
  32'h3d3f59b8 /* (6, 0, 31) */,
  32'h3e709592 /* (2, 0, 31) */,
  32'h3d2d8e0e /* (30, 28, 27) */,
  32'h3d153e19 /* (26, 28, 27) */,
  32'h3d28e3b2 /* (22, 28, 27) */,
  32'h3d53bb31 /* (18, 28, 27) */,
  32'h3d53bb31 /* (14, 28, 27) */,
  32'h3d28e3b2 /* (10, 28, 27) */,
  32'h3d153e19 /* (6, 28, 27) */,
  32'h3d2d8e0e /* (2, 28, 27) */,
  32'h3d149b5c /* (30, 24, 27) */,
  32'h3d22af34 /* (26, 24, 27) */,
  32'h3d5ef675 /* (22, 24, 27) */,
  32'h3d9bc970 /* (18, 24, 27) */,
  32'h3d9bc970 /* (14, 24, 27) */,
  32'h3d5ef675 /* (10, 24, 27) */,
  32'h3d22af34 /* (6, 24, 27) */,
  32'h3d149b5c /* (2, 24, 27) */,
  32'h3d346b02 /* (30, 20, 27) */,
  32'h3d6007ad /* (26, 20, 27) */,
  32'h3db0e528 /* (22, 20, 27) */,
  32'h3e095be4 /* (18, 20, 27) */,
  32'h3e095be4 /* (14, 20, 27) */,
  32'h3db0e528 /* (10, 20, 27) */,
  32'h3d6007ad /* (6, 20, 27) */,
  32'h3d346b02 /* (2, 20, 27) */,
  32'h3d28d1e5 /* (30, 16, 27) */,
  32'h3d5f53fb /* (26, 16, 27) */,
  32'h3dc0863e /* (22, 16, 27) */,
  32'h3e2205a1 /* (18, 16, 27) */,
  32'h3e2205a1 /* (14, 16, 27) */,
  32'h3dc0863e /* (10, 16, 27) */,
  32'h3d5f53fb /* (6, 16, 27) */,
  32'h3d28d1e5 /* (2, 16, 27) */,
  32'h3d346b02 /* (30, 12, 27) */,
  32'h3d6007ad /* (26, 12, 27) */,
  32'h3db0e528 /* (22, 12, 27) */,
  32'h3e095be4 /* (18, 12, 27) */,
  32'h3e095be4 /* (14, 12, 27) */,
  32'h3db0e528 /* (10, 12, 27) */,
  32'h3d6007ad /* (6, 12, 27) */,
  32'h3d346b02 /* (2, 12, 27) */,
  32'h3d149b5c /* (30, 8, 27) */,
  32'h3d22af34 /* (26, 8, 27) */,
  32'h3d5ef675 /* (22, 8, 27) */,
  32'h3d9bc970 /* (18, 8, 27) */,
  32'h3d9bc970 /* (14, 8, 27) */,
  32'h3d5ef675 /* (10, 8, 27) */,
  32'h3d22af34 /* (6, 8, 27) */,
  32'h3d149b5c /* (2, 8, 27) */,
  32'h3d2d8e0e /* (30, 4, 27) */,
  32'h3d153e19 /* (26, 4, 27) */,
  32'h3d28e3b2 /* (22, 4, 27) */,
  32'h3d53bb31 /* (18, 4, 27) */,
  32'h3d53bb31 /* (14, 4, 27) */,
  32'h3d28e3b2 /* (10, 4, 27) */,
  32'h3d153e19 /* (6, 4, 27) */,
  32'h3d2d8e0e /* (2, 4, 27) */,
  32'h3d5dd7d1 /* (30, 0, 27) */,
  32'h3d1b2f33 /* (26, 0, 27) */,
  32'h3d1cee15 /* (22, 0, 27) */,
  32'h3d3b0a55 /* (18, 0, 27) */,
  32'h3d3b0a55 /* (14, 0, 27) */,
  32'h3d1cee15 /* (10, 0, 27) */,
  32'h3d1b2f33 /* (6, 0, 27) */,
  32'h3d5dd7d1 /* (2, 0, 27) */,
  32'h3d14de35 /* (30, 28, 23) */,
  32'h3d2657dd /* (26, 28, 23) */,
  32'h3d68b7a2 /* (22, 28, 23) */,
  32'h3da4db8a /* (18, 28, 23) */,
  32'h3da4db8a /* (14, 28, 23) */,
  32'h3d68b7a2 /* (10, 28, 23) */,
  32'h3d2657dd /* (6, 28, 23) */,
  32'h3d14de35 /* (2, 28, 23) */,
  32'h3d3291f6 /* (30, 24, 23) */,
  32'h3d584c0c /* (26, 24, 23) */,
  32'h3da590e9 /* (22, 24, 23) */,
  32'h3dfaaa60 /* (18, 24, 23) */,
  32'h3dfaaa60 /* (14, 24, 23) */,
  32'h3da590e9 /* (10, 24, 23) */,
  32'h3d584c0c /* (6, 24, 23) */,
  32'h3d3291f6 /* (2, 24, 23) */,
  32'h3d833332 /* (30, 20, 23) */,
  32'h3da96159 /* (26, 20, 23) */,
  32'h3e0cf021 /* (22, 20, 23) */,
  32'h3e654448 /* (18, 20, 23) */,
  32'h3e654448 /* (14, 20, 23) */,
  32'h3e0cf021 /* (10, 20, 23) */,
  32'h3da96159 /* (6, 20, 23) */,
  32'h3d833332 /* (2, 20, 23) */,
  32'h3d87d16b /* (30, 16, 23) */,
  32'h3db6b309 /* (26, 16, 23) */,
  32'h3e21930d /* (22, 16, 23) */,
  32'h3e8b9344 /* (18, 16, 23) */,
  32'h3e8b9344 /* (14, 16, 23) */,
  32'h3e21930d /* (10, 16, 23) */,
  32'h3db6b309 /* (6, 16, 23) */,
  32'h3d87d16b /* (2, 16, 23) */,
  32'h3d833332 /* (30, 12, 23) */,
  32'h3da96159 /* (26, 12, 23) */,
  32'h3e0cf021 /* (22, 12, 23) */,
  32'h3e654448 /* (18, 12, 23) */,
  32'h3e654448 /* (14, 12, 23) */,
  32'h3e0cf021 /* (10, 12, 23) */,
  32'h3da96159 /* (6, 12, 23) */,
  32'h3d833332 /* (2, 12, 23) */,
  32'h3d3291f6 /* (30, 8, 23) */,
  32'h3d584c0c /* (26, 8, 23) */,
  32'h3da590e9 /* (22, 8, 23) */,
  32'h3dfaaa60 /* (18, 8, 23) */,
  32'h3dfaaa60 /* (14, 8, 23) */,
  32'h3da590e9 /* (10, 8, 23) */,
  32'h3d584c0c /* (6, 8, 23) */,
  32'h3d3291f6 /* (2, 8, 23) */,
  32'h3d14de35 /* (30, 4, 23) */,
  32'h3d2657dd /* (26, 4, 23) */,
  32'h3d68b7a2 /* (22, 4, 23) */,
  32'h3da4db8a /* (18, 4, 23) */,
  32'h3da4db8a /* (14, 4, 23) */,
  32'h3d68b7a2 /* (10, 4, 23) */,
  32'h3d2657dd /* (6, 4, 23) */,
  32'h3d14de35 /* (2, 4, 23) */,
  32'h3d11b684 /* (30, 0, 23) */,
  32'h3d1bc36a /* (26, 0, 23) */,
  32'h3d50a575 /* (22, 0, 23) */,
  32'h3d8fa52c /* (18, 0, 23) */,
  32'h3d8fa52c /* (14, 0, 23) */,
  32'h3d50a575 /* (10, 0, 23) */,
  32'h3d1bc36a /* (6, 0, 23) */,
  32'h3d11b684 /* (2, 0, 23) */,
  32'h3d3217f4 /* (30, 28, 19) */,
  32'h3d601ae9 /* (26, 28, 19) */,
  32'h3db40e50 /* (22, 28, 19) */,
  32'h3e0de89e /* (18, 28, 19) */,
  32'h3e0de89e /* (14, 28, 19) */,
  32'h3db40e50 /* (10, 28, 19) */,
  32'h3d601ae9 /* (6, 28, 19) */,
  32'h3d3217f4 /* (2, 28, 19) */,
  32'h3d7b52f8 /* (30, 24, 19) */,
  32'h3da2e7a9 /* (26, 24, 19) */,
  32'h3e085939 /* (22, 24, 19) */,
  32'h3e5f05ce /* (18, 24, 19) */,
  32'h3e5f05ce /* (14, 24, 19) */,
  32'h3e085939 /* (10, 24, 19) */,
  32'h3da2e7a9 /* (6, 24, 19) */,
  32'h3d7b52f8 /* (2, 24, 19) */,
  32'h3dd42d31 /* (30, 20, 19) */,
  32'h3e0dc95f /* (26, 20, 19) */,
  32'h3e7848b5 /* (22, 20, 19) */,
  32'h3ed441df /* (18, 20, 19) */,
  32'h3ed441df /* (14, 20, 19) */,
  32'h3e7848b5 /* (10, 20, 19) */,
  32'h3e0dc95f /* (6, 20, 19) */,
  32'h3dd42d31 /* (2, 20, 19) */,
  32'h3df1ae3d /* (30, 16, 19) */,
  32'h3e2576a9 /* (26, 16, 19) */,
  32'h3e968a40 /* (22, 16, 19) */,
  32'h3f06176f /* (18, 16, 19) */,
  32'h3f06176f /* (14, 16, 19) */,
  32'h3e968a40 /* (10, 16, 19) */,
  32'h3e2576a9 /* (6, 16, 19) */,
  32'h3df1ae3d /* (2, 16, 19) */,
  32'h3dd42d31 /* (30, 12, 19) */,
  32'h3e0dc95f /* (26, 12, 19) */,
  32'h3e7848b5 /* (22, 12, 19) */,
  32'h3ed441df /* (18, 12, 19) */,
  32'h3ed441df /* (14, 12, 19) */,
  32'h3e7848b5 /* (10, 12, 19) */,
  32'h3e0dc95f /* (6, 12, 19) */,
  32'h3dd42d31 /* (2, 12, 19) */,
  32'h3d7b52f8 /* (30, 8, 19) */,
  32'h3da2e7a9 /* (26, 8, 19) */,
  32'h3e085939 /* (22, 8, 19) */,
  32'h3e5f05ce /* (18, 8, 19) */,
  32'h3e5f05ce /* (14, 8, 19) */,
  32'h3e085939 /* (10, 8, 19) */,
  32'h3da2e7a9 /* (6, 8, 19) */,
  32'h3d7b52f8 /* (2, 8, 19) */,
  32'h3d3217f4 /* (30, 4, 19) */,
  32'h3d601ae9 /* (26, 4, 19) */,
  32'h3db40e50 /* (22, 4, 19) */,
  32'h3e0de89e /* (18, 4, 19) */,
  32'h3e0de89e /* (14, 4, 19) */,
  32'h3db40e50 /* (10, 4, 19) */,
  32'h3d601ae9 /* (6, 4, 19) */,
  32'h3d3217f4 /* (2, 4, 19) */,
  32'h3d2045b1 /* (30, 0, 19) */,
  32'h3d4703b2 /* (26, 0, 19) */,
  32'h3d9d248b /* (22, 0, 19) */,
  32'h3df40add /* (18, 0, 19) */,
  32'h3df40add /* (14, 0, 19) */,
  32'h3d9d248b /* (10, 0, 19) */,
  32'h3d4703b2 /* (6, 0, 19) */,
  32'h3d2045b1 /* (2, 0, 19) */,
  32'h3d2d6bba /* (30, 28, 15) */,
  32'h3d61b1de /* (26, 28, 15) */,
  32'h3dbdf4f8 /* (22, 28, 15) */,
  32'h3e1c2ca1 /* (18, 28, 15) */,
  32'h3e1c2ca1 /* (14, 28, 15) */,
  32'h3dbdf4f8 /* (10, 28, 15) */,
  32'h3d61b1de /* (6, 28, 15) */,
  32'h3d2d6bba /* (2, 28, 15) */,
  32'h3d804df8 /* (30, 24, 15) */,
  32'h3daa3349 /* (26, 24, 15) */,
  32'h3e135573 /* (22, 24, 15) */,
  32'h3e79034c /* (18, 24, 15) */,
  32'h3e79034c /* (14, 24, 15) */,
  32'h3e135573 /* (10, 24, 15) */,
  32'h3daa3349 /* (6, 24, 15) */,
  32'h3d804df8 /* (2, 24, 15) */,
  32'h3de39dff /* (30, 20, 15) */,
  32'h3e1a3a56 /* (26, 20, 15) */,
  32'h3e89fde5 /* (22, 20, 15) */,
  32'h3ef15f91 /* (18, 20, 15) */,
  32'h3ef15f91 /* (14, 20, 15) */,
  32'h3e89fde5 /* (10, 20, 15) */,
  32'h3e1a3a56 /* (6, 20, 15) */,
  32'h3de39dff /* (2, 20, 15) */,
  32'h3e06ec2e /* (30, 16, 15) */,
  32'h3e3a3d1a /* (26, 16, 15) */,
  32'h3eabb572 /* (22, 16, 15) */,
  32'h3f1b42bd /* (18, 16, 15) */,
  32'h3f1b42bd /* (14, 16, 15) */,
  32'h3eabb572 /* (10, 16, 15) */,
  32'h3e3a3d1a /* (6, 16, 15) */,
  32'h3e06ec2e /* (2, 16, 15) */,
  32'h3de39dff /* (30, 12, 15) */,
  32'h3e1a3a56 /* (26, 12, 15) */,
  32'h3e89fde5 /* (22, 12, 15) */,
  32'h3ef15f91 /* (18, 12, 15) */,
  32'h3ef15f91 /* (14, 12, 15) */,
  32'h3e89fde5 /* (10, 12, 15) */,
  32'h3e1a3a56 /* (6, 12, 15) */,
  32'h3de39dff /* (2, 12, 15) */,
  32'h3d804df8 /* (30, 8, 15) */,
  32'h3daa3349 /* (26, 8, 15) */,
  32'h3e135573 /* (22, 8, 15) */,
  32'h3e79034c /* (18, 8, 15) */,
  32'h3e79034c /* (14, 8, 15) */,
  32'h3e135573 /* (10, 8, 15) */,
  32'h3daa3349 /* (6, 8, 15) */,
  32'h3d804df8 /* (2, 8, 15) */,
  32'h3d2d6bba /* (30, 4, 15) */,
  32'h3d61b1de /* (26, 4, 15) */,
  32'h3dbdf4f8 /* (22, 4, 15) */,
  32'h3e1c2ca1 /* (18, 4, 15) */,
  32'h3e1c2ca1 /* (14, 4, 15) */,
  32'h3dbdf4f8 /* (10, 4, 15) */,
  32'h3d61b1de /* (6, 4, 15) */,
  32'h3d2d6bba /* (2, 4, 15) */,
  32'h3d18d610 /* (30, 0, 15) */,
  32'h3d455011 /* (26, 0, 15) */,
  32'h3da42e1b /* (22, 0, 15) */,
  32'h3e05899d /* (18, 0, 15) */,
  32'h3e05899d /* (14, 0, 15) */,
  32'h3da42e1b /* (10, 0, 15) */,
  32'h3d455011 /* (6, 0, 15) */,
  32'h3d18d610 /* (2, 0, 15) */,
  32'h3d21c128 /* (30, 28, 11) */,
  32'h3d41fb9f /* (26, 28, 11) */,
  32'h3d92b699 /* (22, 28, 11) */,
  32'h3ddc0819 /* (18, 28, 11) */,
  32'h3ddc0819 /* (14, 28, 11) */,
  32'h3d92b699 /* (10, 28, 11) */,
  32'h3d41fb9f /* (6, 28, 11) */,
  32'h3d21c128 /* (2, 28, 11) */,
  32'h3d558b1c /* (30, 24, 11) */,
  32'h3d865b59 /* (26, 24, 11) */,
  32'h3dd7e578 /* (22, 24, 11) */,
  32'h3e2a27e4 /* (18, 24, 11) */,
  32'h3e2a27e4 /* (14, 24, 11) */,
  32'h3dd7e578 /* (10, 24, 11) */,
  32'h3d865b59 /* (6, 24, 11) */,
  32'h3d558b1c /* (2, 24, 11) */,
  32'h3da96c08 /* (30, 20, 11) */,
  32'h3ddec971 /* (26, 20, 11) */,
  32'h3e3e5baf /* (22, 20, 11) */,
  32'h3e9ecc49 /* (18, 20, 11) */,
  32'h3e9ecc49 /* (14, 20, 11) */,
  32'h3e3e5baf /* (10, 20, 11) */,
  32'h3ddec971 /* (6, 20, 11) */,
  32'h3da96c08 /* (2, 20, 11) */,
  32'h3db86416 /* (30, 16, 11) */,
  32'h3dfa4afe /* (26, 16, 11) */,
  32'h3e60898b /* (22, 16, 11) */,
  32'h3ec4f0a1 /* (18, 16, 11) */,
  32'h3ec4f0a1 /* (14, 16, 11) */,
  32'h3e60898b /* (10, 16, 11) */,
  32'h3dfa4afe /* (6, 16, 11) */,
  32'h3db86416 /* (2, 16, 11) */,
  32'h3da96c08 /* (30, 12, 11) */,
  32'h3ddec971 /* (26, 12, 11) */,
  32'h3e3e5baf /* (22, 12, 11) */,
  32'h3e9ecc49 /* (18, 12, 11) */,
  32'h3e9ecc49 /* (14, 12, 11) */,
  32'h3e3e5baf /* (10, 12, 11) */,
  32'h3ddec971 /* (6, 12, 11) */,
  32'h3da96c08 /* (2, 12, 11) */,
  32'h3d558b1c /* (30, 8, 11) */,
  32'h3d865b59 /* (26, 8, 11) */,
  32'h3dd7e578 /* (22, 8, 11) */,
  32'h3e2a27e4 /* (18, 8, 11) */,
  32'h3e2a27e4 /* (14, 8, 11) */,
  32'h3dd7e578 /* (10, 8, 11) */,
  32'h3d865b59 /* (6, 8, 11) */,
  32'h3d558b1c /* (2, 8, 11) */,
  32'h3d21c128 /* (30, 4, 11) */,
  32'h3d41fb9f /* (26, 4, 11) */,
  32'h3d92b699 /* (22, 4, 11) */,
  32'h3ddc0819 /* (18, 4, 11) */,
  32'h3ddc0819 /* (14, 4, 11) */,
  32'h3d92b699 /* (10, 4, 11) */,
  32'h3d41fb9f /* (6, 4, 11) */,
  32'h3d21c128 /* (2, 4, 11) */,
  32'h3d164ce1 /* (30, 0, 11) */,
  32'h3d3013e2 /* (26, 0, 11) */,
  32'h3d819abc /* (22, 0, 11) */,
  32'h3dbe661f /* (18, 0, 11) */,
  32'h3dbe661f /* (14, 0, 11) */,
  32'h3d819abc /* (10, 0, 11) */,
  32'h3d3013e2 /* (6, 0, 11) */,
  32'h3d164ce1 /* (2, 0, 11) */,
  32'h3d16c6a3 /* (30, 28, 7) */,
  32'h3d17902e /* (26, 28, 7) */,
  32'h3d404057 /* (22, 28, 7) */,
  32'h3d800deb /* (18, 28, 7) */,
  32'h3d800deb /* (14, 28, 7) */,
  32'h3d404057 /* (10, 28, 7) */,
  32'h3d17902e /* (6, 28, 7) */,
  32'h3d16c6a3 /* (2, 28, 7) */,
  32'h3d1d59b0 /* (30, 24, 7) */,
  32'h3d35cd98 /* (26, 24, 7) */,
  32'h3d83c517 /* (22, 24, 7) */,
  32'h3dbf672f /* (18, 24, 7) */,
  32'h3dbf672f /* (14, 24, 7) */,
  32'h3d83c517 /* (10, 24, 7) */,
  32'h3d35cd98 /* (6, 24, 7) */,
  32'h3d1d59b0 /* (2, 24, 7) */,
  32'h3d530d8e /* (30, 20, 7) */,
  32'h3d859348 /* (26, 20, 7) */,
  32'h3dd85675 /* (22, 20, 7) */,
  32'h3e2baf50 /* (18, 20, 7) */,
  32'h3e2baf50 /* (14, 20, 7) */,
  32'h3dd85675 /* (10, 20, 7) */,
  32'h3d859348 /* (6, 20, 7) */,
  32'h3d530d8e /* (2, 20, 7) */,
  32'h3d4f6a6e /* (30, 16, 7) */,
  32'h3d8a46e7 /* (26, 16, 7) */,
  32'h3df142da /* (22, 16, 7) */,
  32'h3e4d7ce8 /* (18, 16, 7) */,
  32'h3e4d7ce8 /* (14, 16, 7) */,
  32'h3df142da /* (10, 16, 7) */,
  32'h3d8a46e7 /* (6, 16, 7) */,
  32'h3d4f6a6e /* (2, 16, 7) */,
  32'h3d530d8e /* (30, 12, 7) */,
  32'h3d859348 /* (26, 12, 7) */,
  32'h3dd85675 /* (22, 12, 7) */,
  32'h3e2baf50 /* (18, 12, 7) */,
  32'h3e2baf50 /* (14, 12, 7) */,
  32'h3dd85675 /* (10, 12, 7) */,
  32'h3d859348 /* (6, 12, 7) */,
  32'h3d530d8e /* (2, 12, 7) */,
  32'h3d1d59b0 /* (30, 8, 7) */,
  32'h3d35cd98 /* (26, 8, 7) */,
  32'h3d83c517 /* (22, 8, 7) */,
  32'h3dbf672f /* (18, 8, 7) */,
  32'h3dbf672f /* (14, 8, 7) */,
  32'h3d83c517 /* (10, 8, 7) */,
  32'h3d35cd98 /* (6, 8, 7) */,
  32'h3d1d59b0 /* (2, 8, 7) */,
  32'h3d16c6a3 /* (30, 4, 7) */,
  32'h3d17902e /* (26, 4, 7) */,
  32'h3d404057 /* (22, 4, 7) */,
  32'h3d800deb /* (18, 4, 7) */,
  32'h3d800deb /* (14, 4, 7) */,
  32'h3d404057 /* (10, 4, 7) */,
  32'h3d17902e /* (6, 4, 7) */,
  32'h3d16c6a3 /* (2, 4, 7) */,
  32'h3d21b235 /* (30, 0, 7) */,
  32'h3d1459dd /* (26, 0, 7) */,
  32'h3d2f5f5a /* (22, 0, 7) */,
  32'h3d60bf24 /* (18, 0, 7) */,
  32'h3d60bf24 /* (14, 0, 7) */,
  32'h3d2f5f5a /* (10, 0, 7) */,
  32'h3d1459dd /* (6, 0, 7) */,
  32'h3d21b235 /* (2, 0, 7) */,
  32'h3d5defd3 /* (30, 28, 3) */,
  32'h3d1b3fff /* (26, 28, 3) */,
  32'h3d1cff11 /* (22, 28, 3) */,
  32'h3d3b1e93 /* (18, 28, 3) */,
  32'h3d3b1e93 /* (14, 28, 3) */,
  32'h3d1cff11 /* (10, 28, 3) */,
  32'h3d1b3fff /* (6, 28, 3) */,
  32'h3d5defd3 /* (2, 28, 3) */,
  32'h3d13e9f7 /* (30, 24, 3) */,
  32'h3d19bf4b /* (26, 24, 3) */,
  32'h3d48bc7e /* (22, 24, 3) */,
  32'h3d880501 /* (18, 24, 3) */,
  32'h3d880501 /* (14, 24, 3) */,
  32'h3d48bc7e /* (10, 24, 3) */,
  32'h3d19bf4b /* (6, 24, 3) */,
  32'h3d13e9f7 /* (2, 24, 3) */,
  32'h3d23d587 /* (30, 20, 3) */,
  32'h3d48406d /* (26, 20, 3) */,
  32'h3d9aff71 /* (22, 20, 3) */,
  32'h3decc5e8 /* (18, 20, 3) */,
  32'h3decc5e8 /* (14, 20, 3) */,
  32'h3d9aff71 /* (10, 20, 3) */,
  32'h3d48406d /* (6, 20, 3) */,
  32'h3d23d587 /* (2, 20, 3) */,
  32'h3d13661d /* (30, 16, 3) */,
  32'h3d41d3ae /* (26, 16, 3) */,
  32'h3da59d10 /* (22, 16, 3) */,
  32'h3e0a27e7 /* (18, 16, 3) */,
  32'h3e0a27e7 /* (14, 16, 3) */,
  32'h3da59d10 /* (10, 16, 3) */,
  32'h3d41d3ae /* (6, 16, 3) */,
  32'h3d13661d /* (2, 16, 3) */,
  32'h3d23d587 /* (30, 12, 3) */,
  32'h3d48406d /* (26, 12, 3) */,
  32'h3d9aff71 /* (22, 12, 3) */,
  32'h3decc5e8 /* (18, 12, 3) */,
  32'h3decc5e8 /* (14, 12, 3) */,
  32'h3d9aff71 /* (10, 12, 3) */,
  32'h3d48406d /* (6, 12, 3) */,
  32'h3d23d587 /* (2, 12, 3) */,
  32'h3d13e9f7 /* (30, 8, 3) */,
  32'h3d19bf4b /* (26, 8, 3) */,
  32'h3d48bc7e /* (22, 8, 3) */,
  32'h3d880501 /* (18, 8, 3) */,
  32'h3d880501 /* (14, 8, 3) */,
  32'h3d48bc7e /* (10, 8, 3) */,
  32'h3d19bf4b /* (6, 8, 3) */,
  32'h3d13e9f7 /* (2, 8, 3) */,
  32'h3d5defd3 /* (30, 4, 3) */,
  32'h3d1b3fff /* (26, 4, 3) */,
  32'h3d1cff11 /* (22, 4, 3) */,
  32'h3d3b1e93 /* (18, 4, 3) */,
  32'h3d3b1e93 /* (14, 4, 3) */,
  32'h3d1cff11 /* (10, 4, 3) */,
  32'h3d1b3fff /* (6, 4, 3) */,
  32'h3d5defd3 /* (2, 4, 3) */,
  32'h3dcbea25 /* (30, 0, 3) */,
  32'h3d2d5b95 /* (26, 0, 3) */,
  32'h3d144f19 /* (22, 0, 3) */,
  32'h3d262b6e /* (18, 0, 3) */,
  32'h3d262b6e /* (14, 0, 3) */,
  32'h3d144f19 /* (10, 0, 3) */,
  32'h3d2d5b95 /* (6, 0, 3) */,
  32'h3dcbea25 /* (2, 0, 3) */,
  32'h3d6eb36b /* (29, 28, 31) */,
  32'h3d17ff6b /* (25, 28, 31) */,
  32'h3d1f5dc3 /* (21, 28, 31) */,
  32'h3d294c4b /* (17, 28, 31) */,
  32'h3d2e802a /* (13, 28, 31) */,
  32'h3d13f199 /* (9, 28, 31) */,
  32'h3d334ee4 /* (5, 28, 31) */,
  32'h3d9c757b /* (1, 28, 31) */,
  32'h3d146963 /* (29, 24, 31) */,
  32'h3d1bb8b6 /* (25, 24, 31) */,
  32'h3d513c3d /* (21, 24, 31) */,
  32'h3d7a003f /* (17, 24, 31) */,
  32'h3d7573b6 /* (13, 24, 31) */,
  32'h3d2fba80 /* (9, 24, 31) */,
  32'h3d1412fd /* (5, 24, 31) */,
  32'h3d1704d7 /* (1, 24, 31) */,
  32'h3d210eee /* (29, 20, 31) */,
  32'h3d4ea8e5 /* (25, 20, 31) */,
  32'h3da53628 /* (21, 20, 31) */,
  32'h3ddd43c2 /* (17, 20, 31) */,
  32'h3dce8d02 /* (13, 20, 31) */,
  32'h3d803124 /* (9, 20, 31) */,
  32'h3d310ad3 /* (5, 20, 31) */,
  32'h3d1a2df1 /* (1, 20, 31) */,
  32'h3d0fbc59 /* (29, 16, 31) */,
  32'h3d49f75a /* (25, 16, 31) */,
  32'h3db336e0 /* (21, 16, 31) */,
  32'h3e02e976 /* (17, 16, 31) */,
  32'h3deaafef /* (13, 16, 31) */,
  32'h3d8420c9 /* (9, 16, 31) */,
  32'h3d24852f /* (5, 16, 31) */,
  32'h3d067e68 /* (1, 16, 31) */,
  32'h3d210eee /* (29, 12, 31) */,
  32'h3d4ea8e5 /* (25, 12, 31) */,
  32'h3da53628 /* (21, 12, 31) */,
  32'h3ddd43c2 /* (17, 12, 31) */,
  32'h3dce8d02 /* (13, 12, 31) */,
  32'h3d803124 /* (9, 12, 31) */,
  32'h3d310ad3 /* (5, 12, 31) */,
  32'h3d1a2df1 /* (1, 12, 31) */,
  32'h3d146963 /* (29, 8, 31) */,
  32'h3d1bb8b6 /* (25, 8, 31) */,
  32'h3d513c3d /* (21, 8, 31) */,
  32'h3d7a003f /* (17, 8, 31) */,
  32'h3d7573b6 /* (13, 8, 31) */,
  32'h3d2fba80 /* (9, 8, 31) */,
  32'h3d1412fd /* (5, 8, 31) */,
  32'h3d1704d7 /* (1, 8, 31) */,
  32'h3d6eb36b /* (29, 4, 31) */,
  32'h3d17ff6b /* (25, 4, 31) */,
  32'h3d1f5dc3 /* (21, 4, 31) */,
  32'h3d294c4b /* (17, 4, 31) */,
  32'h3d2e802a /* (13, 4, 31) */,
  32'h3d13f199 /* (9, 4, 31) */,
  32'h3d334ee4 /* (5, 4, 31) */,
  32'h3d9c757b /* (1, 4, 31) */,
  32'h3dff9e3f /* (29, 0, 31) */,
  32'h3d25463b /* (25, 0, 31) */,
  32'h3d147e90 /* (21, 0, 31) */,
  32'h3d155505 /* (17, 0, 31) */,
  32'h3d1d4601 /* (13, 0, 31) */,
  32'h3d11a5c6 /* (9, 0, 31) */,
  32'h3d6e9998 /* (5, 0, 31) */,
  32'h3f10fe39 /* (1, 0, 31) */,
  32'h3d25f5ce /* (29, 28, 27) */,
  32'h3d1508af /* (25, 28, 27) */,
  32'h3d358341 /* (21, 28, 27) */,
  32'h3d4def9b /* (17, 28, 27) */,
  32'h3d4ea6a0 /* (13, 28, 27) */,
  32'h3d1ee50b /* (9, 28, 27) */,
  32'h3d189061 /* (5, 28, 27) */,
  32'h3d334ee4 /* (1, 28, 27) */,
  32'h3d15d660 /* (29, 24, 27) */,
  32'h3d2bff3e /* (25, 24, 27) */,
  32'h3d77c8fd /* (21, 24, 27) */,
  32'h3d9a5b6b /* (17, 24, 27) */,
  32'h3d94d380 /* (13, 24, 27) */,
  32'h3d49c96c /* (9, 24, 27) */,
  32'h3d1c4d38 /* (5, 24, 27) */,
  32'h3d1412fd /* (1, 24, 27) */,
  32'h3d3a4ebb /* (29, 20, 27) */,
  32'h3d75e4d4 /* (25, 20, 27) */,
  32'h3dca9d53 /* (21, 20, 27) */,
  32'h3e0ae903 /* (17, 20, 27) */,
  32'h3e00477d /* (13, 20, 27) */,
  32'h3d9af1c2 /* (9, 20, 27) */,
  32'h3d4f6dfc /* (5, 20, 27) */,
  32'h3d310ad3 /* (1, 20, 27) */,
  32'h3d3046d8 /* (29, 16, 27) */,
  32'h3d7a662c /* (25, 16, 27) */,
  32'h3de14ffa /* (21, 16, 27) */,
  32'h3e26bbbb /* (17, 16, 27) */,
  32'h3e1486b7 /* (13, 16, 27) */,
  32'h3da4f2f4 /* (9, 16, 27) */,
  32'h3d4ab7f7 /* (5, 16, 27) */,
  32'h3d24852f /* (1, 16, 27) */,
  32'h3d3a4ebb /* (29, 12, 27) */,
  32'h3d75e4d4 /* (25, 12, 27) */,
  32'h3dca9d53 /* (21, 12, 27) */,
  32'h3e0ae903 /* (17, 12, 27) */,
  32'h3e00477d /* (13, 12, 27) */,
  32'h3d9af1c2 /* (9, 12, 27) */,
  32'h3d4f6dfc /* (5, 12, 27) */,
  32'h3d310ad3 /* (1, 12, 27) */,
  32'h3d15d660 /* (29, 8, 27) */,
  32'h3d2bff3e /* (25, 8, 27) */,
  32'h3d77c8fd /* (21, 8, 27) */,
  32'h3d9a5b6b /* (17, 8, 27) */,
  32'h3d94d380 /* (13, 8, 27) */,
  32'h3d49c96c /* (9, 8, 27) */,
  32'h3d1c4d38 /* (5, 8, 27) */,
  32'h3d1412fd /* (1, 8, 27) */,
  32'h3d25f5ce /* (29, 4, 27) */,
  32'h3d1508af /* (25, 4, 27) */,
  32'h3d358341 /* (21, 4, 27) */,
  32'h3d4def9b /* (17, 4, 27) */,
  32'h3d4ea6a0 /* (13, 4, 27) */,
  32'h3d1ee50b /* (9, 4, 27) */,
  32'h3d189061 /* (5, 4, 27) */,
  32'h3d334ee4 /* (1, 4, 27) */,
  32'h3d490b0e /* (29, 0, 27) */,
  32'h3d154f7b /* (25, 0, 27) */,
  32'h3d25e815 /* (21, 0, 27) */,
  32'h3d347f0a /* (17, 0, 27) */,
  32'h3d384488 /* (13, 0, 27) */,
  32'h3d16a564 /* (9, 0, 27) */,
  32'h3d25e3da /* (5, 0, 27) */,
  32'h3d6e9998 /* (1, 0, 27) */,
  32'h3d16b5b2 /* (29, 28, 23) */,
  32'h3d30de15 /* (25, 28, 23) */,
  32'h3d81d711 /* (21, 28, 23) */,
  32'h3da3c1ed /* (17, 28, 23) */,
  32'h3d9d0afa /* (13, 28, 23) */,
  32'h3d51a9d2 /* (9, 28, 23) */,
  32'h3d1ee50b /* (5, 28, 23) */,
  32'h3d13f199 /* (1, 28, 23) */,
  32'h3d37919e /* (29, 24, 23) */,
  32'h3d6b8b35 /* (25, 24, 23) */,
  32'h3dbc4d73 /* (21, 24, 23) */,
  32'h3dfc30a3 /* (17, 24, 23) */,
  32'h3deb6b6d /* (13, 24, 23) */,
  32'h3d921bde /* (9, 24, 23) */,
  32'h3d49c96c /* (5, 24, 23) */,
  32'h3d2fba80 /* (1, 24, 23) */,
  32'h3d886b82 /* (29, 20, 23) */,
  32'h3dbc51f9 /* (25, 20, 23) */,
  32'h3e23781b /* (21, 20, 23) */,
  32'h3e6a25fd /* (17, 20, 23) */,
  32'h3e53dc51 /* (13, 20, 23) */,
  32'h3df3b4f2 /* (9, 20, 23) */,
  32'h3d9af1c2 /* (5, 20, 23) */,
  32'h3d803124 /* (1, 20, 23) */,
  32'h3d8e3848 /* (29, 16, 23) */,
  32'h3dce1075 /* (25, 16, 23) */,
  32'h3e3e5da7 /* (21, 16, 23) */,
  32'h3e908107 /* (17, 16, 23) */,
  32'h3e7e4b9d /* (13, 16, 23) */,
  32'h3e0981d7 /* (9, 16, 23) */,
  32'h3da4f2f4 /* (5, 16, 23) */,
  32'h3d8420c9 /* (1, 16, 23) */,
  32'h3d886b82 /* (29, 12, 23) */,
  32'h3dbc51f9 /* (25, 12, 23) */,
  32'h3e23781b /* (21, 12, 23) */,
  32'h3e6a25fd /* (17, 12, 23) */,
  32'h3e53dc51 /* (13, 12, 23) */,
  32'h3df3b4f2 /* (9, 12, 23) */,
  32'h3d9af1c2 /* (5, 12, 23) */,
  32'h3d803124 /* (1, 12, 23) */,
  32'h3d37919e /* (29, 8, 23) */,
  32'h3d6b8b35 /* (25, 8, 23) */,
  32'h3dbc4d73 /* (21, 8, 23) */,
  32'h3dfc30a3 /* (17, 8, 23) */,
  32'h3deb6b6d /* (13, 8, 23) */,
  32'h3d921bde /* (9, 8, 23) */,
  32'h3d49c96c /* (5, 8, 23) */,
  32'h3d2fba80 /* (1, 8, 23) */,
  32'h3d16b5b2 /* (29, 4, 23) */,
  32'h3d30de15 /* (25, 4, 23) */,
  32'h3d81d711 /* (21, 4, 23) */,
  32'h3da3c1ed /* (17, 4, 23) */,
  32'h3d9d0afa /* (13, 4, 23) */,
  32'h3d51a9d2 /* (9, 4, 23) */,
  32'h3d1ee50b /* (5, 4, 23) */,
  32'h3d13f199 /* (1, 4, 23) */,
  32'h3d1237a7 /* (29, 0, 23) */,
  32'h3d23a039 /* (25, 0, 23) */,
  32'h3d66dac1 /* (21, 0, 23) */,
  32'h3d8df2c1 /* (17, 0, 23) */,
  32'h3d89a49e /* (13, 0, 23) */,
  32'h3d3dc47d /* (9, 0, 23) */,
  32'h3d16a564 /* (5, 0, 23) */,
  32'h3d11a5c6 /* (1, 0, 23) */,
  32'h3d385879 /* (29, 28, 19) */,
  32'h3d770afc /* (25, 28, 19) */,
  32'h3dcf13a3 /* (21, 28, 19) */,
  32'h3e0ff4ce /* (17, 28, 19) */,
  32'h3e0415cb /* (13, 28, 19) */,
  32'h3d9d0afa /* (9, 28, 19) */,
  32'h3d4ea6a0 /* (5, 28, 19) */,
  32'h3d2e802a /* (1, 28, 19) */,
  32'h3d82c188 /* (29, 24, 19) */,
  32'h3db56072 /* (25, 24, 19) */,
  32'h3e1e607d /* (21, 24, 19) */,
  32'h3e640ba2 /* (17, 24, 19) */,
  32'h3e4dd3dc /* (13, 24, 19) */,
  32'h3deb6b6d /* (9, 24, 19) */,
  32'h3d94d380 /* (5, 24, 19) */,
  32'h3d7573b6 /* (1, 24, 19) */,
  32'h3dddef48 /* (29, 20, 19) */,
  32'h3e1f8cbf /* (25, 20, 19) */,
  32'h3e91dfe2 /* (21, 20, 19) */,
  32'h3edb3822 /* (17, 20, 19) */,
  32'h3ec1d890 /* (13, 20, 19) */,
  32'h3e53dc51 /* (9, 20, 19) */,
  32'h3e00477d /* (5, 20, 19) */,
  32'h3dce8d02 /* (1, 20, 19) */,
  32'h3dfdd31f /* (29, 16, 19) */,
  32'h3e3bd4ee /* (25, 16, 19) */,
  32'h3eb2bd2a /* (21, 16, 19) */,
  32'h3f0bd969 /* (17, 16, 19) */,
  32'h3ef27895 /* (13, 16, 19) */,
  32'h3e7e4b9d /* (9, 16, 19) */,
  32'h3e1486b7 /* (5, 16, 19) */,
  32'h3deaafef /* (1, 16, 19) */,
  32'h3dddef48 /* (29, 12, 19) */,
  32'h3e1f8cbf /* (25, 12, 19) */,
  32'h3e91dfe2 /* (21, 12, 19) */,
  32'h3edb3822 /* (17, 12, 19) */,
  32'h3ec1d890 /* (13, 12, 19) */,
  32'h3e53dc51 /* (9, 12, 19) */,
  32'h3e00477d /* (5, 12, 19) */,
  32'h3dce8d02 /* (1, 12, 19) */,
  32'h3d82c188 /* (29, 8, 19) */,
  32'h3db56072 /* (25, 8, 19) */,
  32'h3e1e607d /* (21, 8, 19) */,
  32'h3e640ba2 /* (17, 8, 19) */,
  32'h3e4dd3dc /* (13, 8, 19) */,
  32'h3deb6b6d /* (9, 8, 19) */,
  32'h3d94d380 /* (5, 8, 19) */,
  32'h3d7573b6 /* (1, 8, 19) */,
  32'h3d385879 /* (29, 4, 19) */,
  32'h3d770afc /* (25, 4, 19) */,
  32'h3dcf13a3 /* (21, 4, 19) */,
  32'h3e0ff4ce /* (17, 4, 19) */,
  32'h3e0415cb /* (13, 4, 19) */,
  32'h3d9d0afa /* (9, 4, 19) */,
  32'h3d4ea6a0 /* (5, 4, 19) */,
  32'h3d2e802a /* (1, 4, 19) */,
  32'h3d258110 /* (29, 0, 19) */,
  32'h3d5a6fdd /* (25, 0, 19) */,
  32'h3db3fd83 /* (21, 0, 19) */,
  32'h3df6cc6d /* (17, 0, 19) */,
  32'h3de3e928 /* (13, 0, 19) */,
  32'h3d89a49e /* (9, 0, 19) */,
  32'h3d384488 /* (5, 0, 19) */,
  32'h3d1d4601 /* (1, 0, 19) */,
  32'h3d349293 /* (29, 28, 15) */,
  32'h3d7b9f11 /* (25, 28, 15) */,
  32'h3ddcf428 /* (21, 28, 15) */,
  32'h3e1fe07e /* (17, 28, 15) */,
  32'h3e0ff4ce /* (13, 28, 15) */,
  32'h3da3c1ed /* (9, 28, 15) */,
  32'h3d4def9b /* (5, 28, 15) */,
  32'h3d294c4b /* (1, 28, 15) */,
  32'h3d8608f0 /* (29, 24, 15) */,
  32'h3dbf0444 /* (25, 24, 15) */,
  32'h3e2c9c6c /* (21, 24, 15) */,
  32'h3e803f85 /* (17, 24, 15) */,
  32'h3e640ba2 /* (13, 24, 15) */,
  32'h3dfc30a3 /* (9, 24, 15) */,
  32'h3d9a5b6b /* (5, 24, 15) */,
  32'h3d7a003f /* (1, 24, 15) */,
  32'h3deea44d /* (29, 20, 15) */,
  32'h3e2e6a71 /* (25, 20, 15) */,
  32'h3ea31756 /* (21, 20, 15) */,
  32'h3efaa119 /* (17, 20, 15) */,
  32'h3edb3822 /* (13, 20, 15) */,
  32'h3e6a25fd /* (9, 20, 15) */,
  32'h3e0ae903 /* (5, 20, 15) */,
  32'h3ddd43c2 /* (1, 20, 15) */,
  32'h3e0de417 /* (29, 16, 15) */,
  32'h3e540b9b /* (25, 16, 15) */,
  32'h3ecca1ac /* (21, 16, 15) */,
  32'h3f2286f8 /* (17, 16, 15) */,
  32'h3f0bd969 /* (13, 16, 15) */,
  32'h3e908107 /* (9, 16, 15) */,
  32'h3e26bbbb /* (5, 16, 15) */,
  32'h3e02e976 /* (1, 16, 15) */,
  32'h3deea44d /* (29, 12, 15) */,
  32'h3e2e6a71 /* (25, 12, 15) */,
  32'h3ea31756 /* (21, 12, 15) */,
  32'h3efaa119 /* (17, 12, 15) */,
  32'h3edb3822 /* (13, 12, 15) */,
  32'h3e6a25fd /* (9, 12, 15) */,
  32'h3e0ae903 /* (5, 12, 15) */,
  32'h3ddd43c2 /* (1, 12, 15) */,
  32'h3d8608f0 /* (29, 8, 15) */,
  32'h3dbf0444 /* (25, 8, 15) */,
  32'h3e2c9c6c /* (21, 8, 15) */,
  32'h3e803f85 /* (17, 8, 15) */,
  32'h3e640ba2 /* (13, 8, 15) */,
  32'h3dfc30a3 /* (9, 8, 15) */,
  32'h3d9a5b6b /* (5, 8, 15) */,
  32'h3d7a003f /* (1, 8, 15) */,
  32'h3d349293 /* (29, 4, 15) */,
  32'h3d7b9f11 /* (25, 4, 15) */,
  32'h3ddcf428 /* (21, 4, 15) */,
  32'h3e1fe07e /* (17, 4, 15) */,
  32'h3e0ff4ce /* (13, 4, 15) */,
  32'h3da3c1ed /* (9, 4, 15) */,
  32'h3d4def9b /* (5, 4, 15) */,
  32'h3d294c4b /* (1, 4, 15) */,
  32'h3d1eeabe /* (29, 0, 15) */,
  32'h3d5b6048 /* (25, 0, 15) */,
  32'h3dbe6d47 /* (21, 0, 15) */,
  32'h3e086183 /* (17, 0, 15) */,
  32'h3df6cc6d /* (13, 0, 15) */,
  32'h3d8df2c1 /* (9, 0, 15) */,
  32'h3d347f0a /* (5, 0, 15) */,
  32'h3d155505 /* (1, 0, 15) */,
  32'h3d25fa09 /* (29, 28, 11) */,
  32'h3d52976b /* (25, 28, 11) */,
  32'h3da66ad4 /* (21, 28, 11) */,
  32'h3ddcf428 /* (17, 28, 11) */,
  32'h3dcf13a3 /* (13, 28, 11) */,
  32'h3d81d711 /* (9, 28, 11) */,
  32'h3d358341 /* (5, 28, 11) */,
  32'h3d1f5dc3 /* (1, 28, 11) */,
  32'h3d5d0a38 /* (29, 24, 11) */,
  32'h3d941bce /* (25, 24, 11) */,
  32'h3df84bb3 /* (21, 24, 11) */,
  32'h3e2c9c6c /* (17, 24, 11) */,
  32'h3e1e607d /* (13, 24, 11) */,
  32'h3dbc4d73 /* (9, 24, 11) */,
  32'h3d77c8fd /* (5, 24, 11) */,
  32'h3d513c3d /* (1, 24, 11) */,
  32'h3db0b965 /* (29, 20, 11) */,
  32'h3df94537 /* (25, 20, 11) */,
  32'h3e5e44ac /* (21, 20, 11) */,
  32'h3ea31756 /* (17, 20, 11) */,
  32'h3e91dfe2 /* (13, 20, 11) */,
  32'h3e23781b /* (9, 20, 11) */,
  32'h3dca9d53 /* (5, 20, 11) */,
  32'h3da53628 /* (1, 20, 11) */,
  32'h3dc1602b /* (29, 16, 11) */,
  32'h3e0d9cf0 /* (25, 16, 11) */,
  32'h3e84c8e0 /* (21, 16, 11) */,
  32'h3ecca1ac /* (17, 16, 11) */,
  32'h3eb2bd2a /* (13, 16, 11) */,
  32'h3e3e5da7 /* (9, 16, 11) */,
  32'h3de14ffa /* (5, 16, 11) */,
  32'h3db336e0 /* (1, 16, 11) */,
  32'h3db0b965 /* (29, 12, 11) */,
  32'h3df94537 /* (25, 12, 11) */,
  32'h3e5e44ac /* (21, 12, 11) */,
  32'h3ea31756 /* (17, 12, 11) */,
  32'h3e91dfe2 /* (13, 12, 11) */,
  32'h3e23781b /* (9, 12, 11) */,
  32'h3dca9d53 /* (5, 12, 11) */,
  32'h3da53628 /* (1, 12, 11) */,
  32'h3d5d0a38 /* (29, 8, 11) */,
  32'h3d941bce /* (25, 8, 11) */,
  32'h3df84bb3 /* (21, 8, 11) */,
  32'h3e2c9c6c /* (17, 8, 11) */,
  32'h3e1e607d /* (13, 8, 11) */,
  32'h3dbc4d73 /* (9, 8, 11) */,
  32'h3d77c8fd /* (5, 8, 11) */,
  32'h3d513c3d /* (1, 8, 11) */,
  32'h3d25fa09 /* (29, 4, 11) */,
  32'h3d52976b /* (25, 4, 11) */,
  32'h3da66ad4 /* (21, 4, 11) */,
  32'h3ddcf428 /* (17, 4, 11) */,
  32'h3dcf13a3 /* (13, 4, 11) */,
  32'h3d81d711 /* (9, 4, 11) */,
  32'h3d358341 /* (5, 4, 11) */,
  32'h3d1f5dc3 /* (1, 4, 11) */,
  32'h3d198ce9 /* (29, 0, 11) */,
  32'h3d3dcd22 /* (25, 0, 11) */,
  32'h3d922642 /* (21, 0, 11) */,
  32'h3dbe6d47 /* (17, 0, 11) */,
  32'h3db3fd83 /* (13, 0, 11) */,
  32'h3d66dac1 /* (9, 0, 11) */,
  32'h3d25e815 /* (5, 0, 11) */,
  32'h3d147e90 /* (1, 0, 11) */,
  32'h3d155fa4 /* (29, 28, 7) */,
  32'h3d1cbb18 /* (25, 28, 7) */,
  32'h3d52976b /* (21, 28, 7) */,
  32'h3d7b9f11 /* (17, 28, 7) */,
  32'h3d770afc /* (13, 28, 7) */,
  32'h3d30de15 /* (9, 28, 7) */,
  32'h3d1508af /* (5, 28, 7) */,
  32'h3d17ff6b /* (1, 28, 7) */,
  32'h3d2054cd /* (29, 24, 7) */,
  32'h3d432bf1 /* (25, 24, 7) */,
  32'h3d941bce /* (21, 24, 7) */,
  32'h3dbf0444 /* (17, 24, 7) */,
  32'h3db56072 /* (13, 24, 7) */,
  32'h3d6b8b35 /* (9, 24, 7) */,
  32'h3d2bff3e /* (5, 24, 7) */,
  32'h3d1bb8b6 /* (1, 24, 7) */,
  32'h3d5ab0e1 /* (29, 20, 7) */,
  32'h3d938890 /* (25, 20, 7) */,
  32'h3df94537 /* (21, 20, 7) */,
  32'h3e2e6a71 /* (17, 20, 7) */,
  32'h3e1f8cbf /* (13, 20, 7) */,
  32'h3dbc51f9 /* (9, 20, 7) */,
  32'h3d75e4d4 /* (5, 20, 7) */,
  32'h3d4ea8e5 /* (1, 20, 7) */,
  32'h3d58de26 /* (29, 16, 7) */,
  32'h3d9b7830 /* (25, 16, 7) */,
  32'h3e0d9cf0 /* (21, 16, 7) */,
  32'h3e540b9b /* (17, 16, 7) */,
  32'h3e3bd4ee /* (13, 16, 7) */,
  32'h3dce1075 /* (9, 16, 7) */,
  32'h3d7a662c /* (5, 16, 7) */,
  32'h3d49f75a /* (1, 16, 7) */,
  32'h3d5ab0e1 /* (29, 12, 7) */,
  32'h3d938890 /* (25, 12, 7) */,
  32'h3df94537 /* (21, 12, 7) */,
  32'h3e2e6a71 /* (17, 12, 7) */,
  32'h3e1f8cbf /* (13, 12, 7) */,
  32'h3dbc51f9 /* (9, 12, 7) */,
  32'h3d75e4d4 /* (5, 12, 7) */,
  32'h3d4ea8e5 /* (1, 12, 7) */,
  32'h3d2054cd /* (29, 8, 7) */,
  32'h3d432bf1 /* (25, 8, 7) */,
  32'h3d941bce /* (21, 8, 7) */,
  32'h3dbf0444 /* (17, 8, 7) */,
  32'h3db56072 /* (13, 8, 7) */,
  32'h3d6b8b35 /* (9, 8, 7) */,
  32'h3d2bff3e /* (5, 8, 7) */,
  32'h3d1bb8b6 /* (1, 8, 7) */,
  32'h3d155fa4 /* (29, 4, 7) */,
  32'h3d1cbb18 /* (25, 4, 7) */,
  32'h3d52976b /* (21, 4, 7) */,
  32'h3d7b9f11 /* (17, 4, 7) */,
  32'h3d770afc /* (13, 4, 7) */,
  32'h3d30de15 /* (9, 4, 7) */,
  32'h3d1508af /* (5, 4, 7) */,
  32'h3d17ff6b /* (1, 4, 7) */,
  32'h3d1cfd70 /* (29, 0, 7) */,
  32'h3d162f74 /* (25, 0, 7) */,
  32'h3d3dcd22 /* (21, 0, 7) */,
  32'h3d5b6048 /* (17, 0, 7) */,
  32'h3d5a6fdd /* (13, 0, 7) */,
  32'h3d23a039 /* (9, 0, 7) */,
  32'h3d154f7b /* (5, 0, 7) */,
  32'h3d25463b /* (1, 0, 7) */,
  32'h3d4920d0 /* (29, 28, 3) */,
  32'h3d155fa4 /* (25, 28, 3) */,
  32'h3d25fa09 /* (21, 28, 3) */,
  32'h3d349293 /* (17, 28, 3) */,
  32'h3d385879 /* (13, 28, 3) */,
  32'h3d16b5b2 /* (9, 28, 3) */,
  32'h3d25f5ce /* (5, 28, 3) */,
  32'h3d6eb36b /* (1, 28, 3) */,
  32'h3d1392fe /* (29, 24, 3) */,
  32'h3d2054cd /* (25, 24, 3) */,
  32'h3d5d0a38 /* (21, 24, 3) */,
  32'h3d8608f0 /* (17, 24, 3) */,
  32'h3d82c188 /* (13, 24, 3) */,
  32'h3d37919e /* (9, 24, 3) */,
  32'h3d15d660 /* (5, 24, 3) */,
  32'h3d146963 /* (1, 24, 3) */,
  32'h3d28b308 /* (29, 20, 3) */,
  32'h3d5ab0e1 /* (25, 20, 3) */,
  32'h3db0b965 /* (21, 20, 3) */,
  32'h3deea44d /* (17, 20, 3) */,
  32'h3dddef48 /* (13, 20, 3) */,
  32'h3d886b82 /* (9, 20, 3) */,
  32'h3d3a4ebb /* (5, 20, 3) */,
  32'h3d210eee /* (1, 20, 3) */,
  32'h3d19c07a /* (29, 16, 3) */,
  32'h3d58de26 /* (25, 16, 3) */,
  32'h3dc1602b /* (21, 16, 3) */,
  32'h3e0de417 /* (17, 16, 3) */,
  32'h3dfdd31f /* (13, 16, 3) */,
  32'h3d8e3848 /* (9, 16, 3) */,
  32'h3d3046d8 /* (5, 16, 3) */,
  32'h3d0fbc59 /* (1, 16, 3) */,
  32'h3d28b308 /* (29, 12, 3) */,
  32'h3d5ab0e1 /* (25, 12, 3) */,
  32'h3db0b965 /* (21, 12, 3) */,
  32'h3deea44d /* (17, 12, 3) */,
  32'h3dddef48 /* (13, 12, 3) */,
  32'h3d886b82 /* (9, 12, 3) */,
  32'h3d3a4ebb /* (5, 12, 3) */,
  32'h3d210eee /* (1, 12, 3) */,
  32'h3d1392fe /* (29, 8, 3) */,
  32'h3d2054cd /* (25, 8, 3) */,
  32'h3d5d0a38 /* (21, 8, 3) */,
  32'h3d8608f0 /* (17, 8, 3) */,
  32'h3d82c188 /* (13, 8, 3) */,
  32'h3d37919e /* (9, 8, 3) */,
  32'h3d15d660 /* (5, 8, 3) */,
  32'h3d146963 /* (1, 8, 3) */,
  32'h3d4920d0 /* (29, 4, 3) */,
  32'h3d155fa4 /* (25, 4, 3) */,
  32'h3d25fa09 /* (21, 4, 3) */,
  32'h3d349293 /* (17, 4, 3) */,
  32'h3d385879 /* (13, 4, 3) */,
  32'h3d16b5b2 /* (9, 4, 3) */,
  32'h3d25f5ce /* (5, 4, 3) */,
  32'h3d6eb36b /* (1, 4, 3) */,
  32'h3d9c797c /* (29, 0, 3) */,
  32'h3d1cfd70 /* (25, 0, 3) */,
  32'h3d198ce9 /* (21, 0, 3) */,
  32'h3d1eeabe /* (17, 0, 3) */,
  32'h3d258110 /* (13, 0, 3) */,
  32'h3d1237a7 /* (9, 0, 3) */,
  32'h3d490b0e /* (5, 0, 3) */,
  32'h3dff9e3f /* (1, 0, 3) */,
  32'h3d4cb45d /* (28, 28, 31) */,
  32'h3d139499 /* (24, 28, 31) */,
  32'h3d27af27 /* (20, 28, 31) */,
  32'h3d18708b /* (16, 28, 31) */,
  32'h3d27af27 /* (12, 28, 31) */,
  32'h3d139499 /* (8, 28, 31) */,
  32'h3d4cb45d /* (4, 28, 31) */,
  32'h3da3aa58 /* (0, 28, 31) */,
  32'h3d139499 /* (28, 24, 31) */,
  32'h3d23fb6f /* (24, 24, 31) */,
  32'h3d649547 /* (20, 24, 31) */,
  32'h3d656b11 /* (16, 24, 31) */,
  32'h3d649547 /* (12, 24, 31) */,
  32'h3d23fb6f /* (8, 24, 31) */,
  32'h3d139499 /* (4, 24, 31) */,
  32'h3d177e6a /* (0, 24, 31) */,
  32'h3d27af27 /* (28, 20, 31) */,
  32'h3d649547 /* (24, 20, 31) */,
  32'h3dbaaaa9 /* (20, 20, 31) */,
  32'h3dcf60c6 /* (16, 20, 31) */,
  32'h3dbaaaa9 /* (12, 20, 31) */,
  32'h3d649547 /* (8, 20, 31) */,
  32'h3d27af27 /* (4, 20, 31) */,
  32'h3d195f14 /* (0, 20, 31) */,
  32'h3d18708b /* (28, 16, 31) */,
  32'h3d656b11 /* (24, 16, 31) */,
  32'h3dcf60c6 /* (20, 16, 31) */,
  32'h3df9e164 /* (16, 16, 31) */,
  32'h3dcf60c6 /* (12, 16, 31) */,
  32'h3d656b11 /* (8, 16, 31) */,
  32'h3d18708b /* (4, 16, 31) */,
  32'h3d0563b9 /* (0, 16, 31) */,
  32'h3d27af27 /* (28, 12, 31) */,
  32'h3d649547 /* (24, 12, 31) */,
  32'h3dbaaaa9 /* (20, 12, 31) */,
  32'h3dcf60c6 /* (16, 12, 31) */,
  32'h3dbaaaa9 /* (12, 12, 31) */,
  32'h3d649547 /* (8, 12, 31) */,
  32'h3d27af27 /* (4, 12, 31) */,
  32'h3d195f14 /* (0, 12, 31) */,
  32'h3d139499 /* (28, 8, 31) */,
  32'h3d23fb6f /* (24, 8, 31) */,
  32'h3d649547 /* (20, 8, 31) */,
  32'h3d656b11 /* (16, 8, 31) */,
  32'h3d649547 /* (12, 8, 31) */,
  32'h3d23fb6f /* (8, 8, 31) */,
  32'h3d139499 /* (4, 8, 31) */,
  32'h3d177e6a /* (0, 8, 31) */,
  32'h3d4cb45d /* (28, 4, 31) */,
  32'h3d139499 /* (24, 4, 31) */,
  32'h3d27af27 /* (20, 4, 31) */,
  32'h3d18708b /* (16, 4, 31) */,
  32'h3d27af27 /* (12, 4, 31) */,
  32'h3d139499 /* (8, 4, 31) */,
  32'h3d4cb45d /* (4, 4, 31) */,
  32'h3da3aa58 /* (0, 4, 31) */,
  32'h3da3aa58 /* (28, 0, 31) */,
  32'h3d177e6a /* (24, 0, 31) */,
  32'h3d195f14 /* (20, 0, 31) */,
  32'h3d0563b9 /* (16, 0, 31) */,
  32'h3d195f14 /* (12, 0, 31) */,
  32'h3d177e6a /* (8, 0, 31) */,
  32'h3da3aa58 /* (4, 0, 31) */,
  32'h3f8f3ec8 /* (0, 0, 31) */,
  32'h3d1e7527 /* (28, 28, 27) */,
  32'h3d183845 /* (24, 28, 27) */,
  32'h3d431db1 /* (20, 28, 27) */,
  32'h3d3b5943 /* (16, 28, 27) */,
  32'h3d431db1 /* (12, 28, 27) */,
  32'h3d183845 /* (8, 28, 27) */,
  32'h3d1e7527 /* (4, 28, 27) */,
  32'h3d3577a5 /* (0, 28, 27) */,
  32'h3d183845 /* (28, 24, 27) */,
  32'h3d38dbff /* (24, 24, 27) */,
  32'h3d89129f /* (20, 24, 27) */,
  32'h3d8eb3bf /* (16, 24, 27) */,
  32'h3d89129f /* (12, 24, 27) */,
  32'h3d38dbff /* (8, 24, 27) */,
  32'h3d183845 /* (4, 24, 27) */,
  32'h3d13eed3 /* (0, 24, 27) */,
  32'h3d431db1 /* (28, 20, 27) */,
  32'h3d89129f /* (24, 20, 27) */,
  32'h3de671da /* (20, 20, 27) */,
  32'h3e02cee2 /* (16, 20, 27) */,
  32'h3de671da /* (12, 20, 27) */,
  32'h3d89129f /* (8, 20, 27) */,
  32'h3d431db1 /* (4, 20, 27) */,
  32'h3d2ff16f /* (0, 20, 27) */,
  32'h3d3b5943 /* (28, 16, 27) */,
  32'h3d8eb3bf /* (24, 16, 27) */,
  32'h3e02cee2 /* (20, 16, 27) */,
  32'h3e1f95bf /* (16, 16, 27) */,
  32'h3e02cee2 /* (12, 16, 27) */,
  32'h3d8eb3bf /* (8, 16, 27) */,
  32'h3d3b5943 /* (4, 16, 27) */,
  32'h3d231d8f /* (0, 16, 27) */,
  32'h3d431db1 /* (28, 12, 27) */,
  32'h3d89129f /* (24, 12, 27) */,
  32'h3de671da /* (20, 12, 27) */,
  32'h3e02cee2 /* (16, 12, 27) */,
  32'h3de671da /* (12, 12, 27) */,
  32'h3d89129f /* (8, 12, 27) */,
  32'h3d431db1 /* (4, 12, 27) */,
  32'h3d2ff16f /* (0, 12, 27) */,
  32'h3d183845 /* (28, 8, 27) */,
  32'h3d38dbff /* (24, 8, 27) */,
  32'h3d89129f /* (20, 8, 27) */,
  32'h3d8eb3bf /* (16, 8, 27) */,
  32'h3d89129f /* (12, 8, 27) */,
  32'h3d38dbff /* (8, 8, 27) */,
  32'h3d183845 /* (4, 8, 27) */,
  32'h3d13eed3 /* (0, 8, 27) */,
  32'h3d1e7527 /* (28, 4, 27) */,
  32'h3d183845 /* (24, 4, 27) */,
  32'h3d431db1 /* (20, 4, 27) */,
  32'h3d3b5943 /* (16, 4, 27) */,
  32'h3d431db1 /* (12, 4, 27) */,
  32'h3d183845 /* (8, 4, 27) */,
  32'h3d1e7527 /* (4, 4, 27) */,
  32'h3d3577a5 /* (0, 4, 27) */,
  32'h3d3577a5 /* (28, 0, 27) */,
  32'h3d13eed3 /* (24, 0, 27) */,
  32'h3d2ff16f /* (20, 0, 27) */,
  32'h3d231d8f /* (16, 0, 27) */,
  32'h3d2ff16f /* (12, 0, 27) */,
  32'h3d13eed3 /* (8, 0, 27) */,
  32'h3d3577a5 /* (4, 0, 27) */,
  32'h3d75271a /* (0, 0, 27) */,
  32'h3d19e157 /* (28, 28, 23) */,
  32'h3d3f1eea /* (24, 28, 23) */,
  32'h3d902ce0 /* (20, 28, 23) */,
  32'h3d97bb42 /* (16, 28, 23) */,
  32'h3d902ce0 /* (12, 28, 23) */,
  32'h3d3f1eea /* (8, 28, 23) */,
  32'h3d19e157 /* (4, 28, 23) */,
  32'h3d13aacb /* (0, 28, 23) */,
  32'h3d3f1eea /* (28, 24, 23) */,
  32'h3d824402 /* (24, 24, 23) */,
  32'h3dd4c19e /* (20, 24, 23) */,
  32'h3dec5cc9 /* (16, 24, 23) */,
  32'h3dd4c19e /* (12, 24, 23) */,
  32'h3d824402 /* (8, 24, 23) */,
  32'h3d3f1eea /* (4, 24, 23) */,
  32'h3d2eceba /* (0, 24, 23) */,
  32'h3d902ce0 /* (28, 20, 23) */,
  32'h3dd4c19e /* (24, 20, 23) */,
  32'h3e3c290c /* (20, 20, 23) */,
  32'h3e5e82df /* (16, 20, 23) */,
  32'h3e3c290c /* (12, 20, 23) */,
  32'h3dd4c19e /* (8, 20, 23) */,
  32'h3d902ce0 /* (4, 20, 23) */,
  32'h3d7e6b4b /* (0, 20, 23) */,
  32'h3d97bb42 /* (28, 16, 23) */,
  32'h3dec5cc9 /* (24, 16, 23) */,
  32'h3e5e82df /* (20, 16, 23) */,
  32'h3e8b1bdf /* (16, 16, 23) */,
  32'h3e5e82df /* (12, 16, 23) */,
  32'h3dec5cc9 /* (8, 16, 23) */,
  32'h3d97bb42 /* (4, 16, 23) */,
  32'h3d82ec35 /* (0, 16, 23) */,
  32'h3d902ce0 /* (28, 12, 23) */,
  32'h3dd4c19e /* (24, 12, 23) */,
  32'h3e3c290c /* (20, 12, 23) */,
  32'h3e5e82df /* (16, 12, 23) */,
  32'h3e3c290c /* (12, 12, 23) */,
  32'h3dd4c19e /* (8, 12, 23) */,
  32'h3d902ce0 /* (4, 12, 23) */,
  32'h3d7e6b4b /* (0, 12, 23) */,
  32'h3d3f1eea /* (28, 8, 23) */,
  32'h3d824402 /* (24, 8, 23) */,
  32'h3dd4c19e /* (20, 8, 23) */,
  32'h3dec5cc9 /* (16, 8, 23) */,
  32'h3dd4c19e /* (12, 8, 23) */,
  32'h3d824402 /* (8, 8, 23) */,
  32'h3d3f1eea /* (4, 8, 23) */,
  32'h3d2eceba /* (0, 8, 23) */,
  32'h3d19e157 /* (28, 4, 23) */,
  32'h3d3f1eea /* (24, 4, 23) */,
  32'h3d902ce0 /* (20, 4, 23) */,
  32'h3d97bb42 /* (16, 4, 23) */,
  32'h3d902ce0 /* (12, 4, 23) */,
  32'h3d3f1eea /* (8, 4, 23) */,
  32'h3d19e157 /* (4, 4, 23) */,
  32'h3d13aacb /* (0, 4, 23) */,
  32'h3d13aacb /* (28, 0, 23) */,
  32'h3d2eceba /* (24, 0, 23) */,
  32'h3d7e6b4b /* (20, 0, 23) */,
  32'h3d82ec35 /* (16, 0, 23) */,
  32'h3d7e6b4b /* (12, 0, 23) */,
  32'h3d2eceba /* (8, 0, 23) */,
  32'h3d13aacb /* (4, 0, 23) */,
  32'h3d11ab15 /* (0, 0, 23) */,
  32'h3d41aa67 /* (28, 28, 19) */,
  32'h3d8a5278 /* (24, 28, 19) */,
  32'h3dec6d9f /* (20, 28, 19) */,
  32'h3e07f264 /* (16, 28, 19) */,
  32'h3dec6d9f /* (12, 28, 19) */,
  32'h3d8a5278 /* (8, 28, 19) */,
  32'h3d41aa67 /* (4, 28, 19) */,
  32'h3d2d543a /* (0, 28, 19) */,
  32'h3d8a5278 /* (28, 24, 19) */,
  32'h3dcd36cb /* (24, 24, 19) */,
  32'h3e368e5b /* (20, 24, 19) */,
  32'h3e58f4b1 /* (16, 24, 19) */,
  32'h3e368e5b /* (12, 24, 19) */,
  32'h3dcd36cb /* (8, 24, 19) */,
  32'h3d8a5278 /* (4, 24, 19) */,
  32'h3d7388b1 /* (0, 24, 19) */,
  32'h3dec6d9f /* (28, 20, 19) */,
  32'h3e368e5b /* (24, 20, 19) */,
  32'h3eaa0eb2 /* (20, 20, 19) */,
  32'h3ed28b29 /* (16, 20, 19) */,
  32'h3eaa0eb2 /* (12, 20, 19) */,
  32'h3e368e5b /* (8, 20, 19) */,
  32'h3dec6d9f /* (4, 20, 19) */,
  32'h3dccb681 /* (0, 20, 19) */,
  32'h3e07f264 /* (28, 16, 19) */,
  32'h3e58f4b1 /* (24, 16, 19) */,
  32'h3ed28b29 /* (20, 16, 19) */,
  32'h3f079668 /* (16, 16, 19) */,
  32'h3ed28b29 /* (12, 16, 19) */,
  32'h3e58f4b1 /* (8, 16, 19) */,
  32'h3e07f264 /* (4, 16, 19) */,
  32'h3de8675d /* (0, 16, 19) */,
  32'h3dec6d9f /* (28, 12, 19) */,
  32'h3e368e5b /* (24, 12, 19) */,
  32'h3eaa0eb2 /* (20, 12, 19) */,
  32'h3ed28b29 /* (16, 12, 19) */,
  32'h3eaa0eb2 /* (12, 12, 19) */,
  32'h3e368e5b /* (8, 12, 19) */,
  32'h3dec6d9f /* (4, 12, 19) */,
  32'h3dccb681 /* (0, 12, 19) */,
  32'h3d8a5278 /* (28, 8, 19) */,
  32'h3dcd36cb /* (24, 8, 19) */,
  32'h3e368e5b /* (20, 8, 19) */,
  32'h3e58f4b1 /* (16, 8, 19) */,
  32'h3e368e5b /* (12, 8, 19) */,
  32'h3dcd36cb /* (8, 8, 19) */,
  32'h3d8a5278 /* (4, 8, 19) */,
  32'h3d7388b1 /* (0, 8, 19) */,
  32'h3d41aa67 /* (28, 4, 19) */,
  32'h3d8a5278 /* (24, 4, 19) */,
  32'h3dec6d9f /* (20, 4, 19) */,
  32'h3e07f264 /* (16, 4, 19) */,
  32'h3dec6d9f /* (12, 4, 19) */,
  32'h3d8a5278 /* (8, 4, 19) */,
  32'h3d41aa67 /* (4, 4, 19) */,
  32'h3d2d543a /* (0, 4, 19) */,
  32'h3d2d543a /* (28, 0, 19) */,
  32'h3d7388b1 /* (24, 0, 19) */,
  32'h3dccb681 /* (20, 0, 19) */,
  32'h3de8675d /* (16, 0, 19) */,
  32'h3dccb681 /* (12, 0, 19) */,
  32'h3d7388b1 /* (8, 0, 19) */,
  32'h3d2d543a /* (4, 0, 19) */,
  32'h3d1c4c09 /* (0, 0, 19) */,
  32'h3d3f317e /* (28, 28, 15) */,
  32'h3d8e8b3a /* (24, 28, 15) */,
  32'h3dff07bf /* (20, 28, 15) */,
  32'h3e18449a /* (16, 28, 15) */,
  32'h3dff07bf /* (12, 28, 15) */,
  32'h3d8e8b3a /* (8, 28, 15) */,
  32'h3d3f317e /* (4, 28, 15) */,
  32'h3d27f384 /* (0, 28, 15) */,
  32'h3d8e8b3a /* (28, 24, 15) */,
  32'h3dd9f1d0 /* (24, 24, 15) */,
  32'h3e48a298 /* (20, 24, 15) */,
  32'h3e75b861 /* (16, 24, 15) */,
  32'h3e48a298 /* (12, 24, 15) */,
  32'h3dd9f1d0 /* (8, 24, 15) */,
  32'h3d8e8b3a /* (4, 24, 15) */,
  32'h3d77d78b /* (0, 24, 15) */,
  32'h3dff07bf /* (28, 20, 15) */,
  32'h3e48a298 /* (24, 20, 15) */,
  32'h3ebf3a63 /* (20, 20, 15) */,
  32'h3ef1f40b /* (16, 20, 15) */,
  32'h3ebf3a63 /* (12, 20, 15) */,
  32'h3e48a298 /* (8, 20, 15) */,
  32'h3dff07bf /* (4, 20, 15) */,
  32'h3ddb309a /* (0, 20, 15) */,
  32'h3e18449a /* (28, 16, 15) */,
  32'h3e75b861 /* (24, 16, 15) */,
  32'h3ef1f40b /* (20, 16, 15) */,
  32'h3f1e253a /* (16, 16, 15) */,
  32'h3ef1f40b /* (12, 16, 15) */,
  32'h3e75b861 /* (8, 16, 15) */,
  32'h3e18449a /* (4, 16, 15) */,
  32'h3e019a4f /* (0, 16, 15) */,
  32'h3dff07bf /* (28, 12, 15) */,
  32'h3e48a298 /* (24, 12, 15) */,
  32'h3ebf3a63 /* (20, 12, 15) */,
  32'h3ef1f40b /* (16, 12, 15) */,
  32'h3ebf3a63 /* (12, 12, 15) */,
  32'h3e48a298 /* (8, 12, 15) */,
  32'h3dff07bf /* (4, 12, 15) */,
  32'h3ddb309a /* (0, 12, 15) */,
  32'h3d8e8b3a /* (28, 8, 15) */,
  32'h3dd9f1d0 /* (24, 8, 15) */,
  32'h3e48a298 /* (20, 8, 15) */,
  32'h3e75b861 /* (16, 8, 15) */,
  32'h3e48a298 /* (12, 8, 15) */,
  32'h3dd9f1d0 /* (8, 8, 15) */,
  32'h3d8e8b3a /* (4, 8, 15) */,
  32'h3d77d78b /* (0, 8, 15) */,
  32'h3d3f317e /* (28, 4, 15) */,
  32'h3d8e8b3a /* (24, 4, 15) */,
  32'h3dff07bf /* (20, 4, 15) */,
  32'h3e18449a /* (16, 4, 15) */,
  32'h3dff07bf /* (12, 4, 15) */,
  32'h3d8e8b3a /* (8, 4, 15) */,
  32'h3d3f317e /* (4, 4, 15) */,
  32'h3d27f384 /* (0, 4, 15) */,
  32'h3d27f384 /* (28, 0, 15) */,
  32'h3d77d78b /* (24, 0, 15) */,
  32'h3ddb309a /* (20, 0, 15) */,
  32'h3e019a4f /* (16, 0, 15) */,
  32'h3ddb309a /* (12, 0, 15) */,
  32'h3d77d78b /* (8, 0, 15) */,
  32'h3d27f384 /* (4, 0, 15) */,
  32'h3d14300c /* (0, 0, 15) */,
  32'h3d2c64eb /* (28, 28, 11) */,
  32'h3d683712 /* (24, 28, 11) */,
  32'h3dbb90ec /* (20, 28, 11) */,
  32'h3dcebbc1 /* (16, 28, 11) */,
  32'h3dbb90ec /* (12, 28, 11) */,
  32'h3d683712 /* (8, 28, 11) */,
  32'h3d2c64eb /* (4, 28, 11) */,
  32'h3d1e982c /* (0, 28, 11) */,
  32'h3d683712 /* (28, 24, 11) */,
  32'h3da5dafd /* (24, 24, 11) */,
  32'h3e0dbead /* (20, 24, 11) */,
  32'h3e2301df /* (16, 24, 11) */,
  32'h3e0dbead /* (12, 24, 11) */,
  32'h3da5dafd /* (8, 24, 11) */,
  32'h3d683712 /* (4, 24, 11) */,
  32'h3d4fd499 /* (0, 24, 11) */,
  32'h3dbb90ec /* (28, 20, 11) */,
  32'h3e0dbead /* (24, 20, 11) */,
  32'h3e80c082 /* (20, 20, 11) */,
  32'h3e9bce24 /* (16, 20, 11) */,
  32'h3e80c082 /* (12, 20, 11) */,
  32'h3e0dbead /* (8, 20, 11) */,
  32'h3dbb90ec /* (4, 20, 11) */,
  32'h3da3d600 /* (0, 20, 11) */,
  32'h3dcebbc1 /* (28, 16, 11) */,
  32'h3e2301df /* (24, 16, 11) */,
  32'h3e9bce24 /* (20, 16, 11) */,
  32'h3ec5ad99 /* (16, 16, 11) */,
  32'h3e9bce24 /* (12, 16, 11) */,
  32'h3e2301df /* (8, 16, 11) */,
  32'h3dcebbc1 /* (4, 16, 11) */,
  32'h3db1860e /* (0, 16, 11) */,
  32'h3dbb90ec /* (28, 12, 11) */,
  32'h3e0dbead /* (24, 12, 11) */,
  32'h3e80c082 /* (20, 12, 11) */,
  32'h3e9bce24 /* (16, 12, 11) */,
  32'h3e80c082 /* (12, 12, 11) */,
  32'h3e0dbead /* (8, 12, 11) */,
  32'h3dbb90ec /* (4, 12, 11) */,
  32'h3da3d600 /* (0, 12, 11) */,
  32'h3d683712 /* (28, 8, 11) */,
  32'h3da5dafd /* (24, 8, 11) */,
  32'h3e0dbead /* (20, 8, 11) */,
  32'h3e2301df /* (16, 8, 11) */,
  32'h3e0dbead /* (12, 8, 11) */,
  32'h3da5dafd /* (8, 8, 11) */,
  32'h3d683712 /* (4, 8, 11) */,
  32'h3d4fd499 /* (0, 8, 11) */,
  32'h3d2c64eb /* (28, 4, 11) */,
  32'h3d683712 /* (24, 4, 11) */,
  32'h3dbb90ec /* (20, 4, 11) */,
  32'h3dcebbc1 /* (16, 4, 11) */,
  32'h3dbb90ec /* (12, 4, 11) */,
  32'h3d683712 /* (8, 4, 11) */,
  32'h3d2c64eb /* (4, 4, 11) */,
  32'h3d1e982c /* (0, 4, 11) */,
  32'h3d1e982c /* (28, 0, 11) */,
  32'h3d4fd499 /* (24, 0, 11) */,
  32'h3da3d600 /* (20, 0, 11) */,
  32'h3db1860e /* (16, 0, 11) */,
  32'h3da3d600 /* (12, 0, 11) */,
  32'h3d4fd499 /* (8, 0, 11) */,
  32'h3d1e982c /* (4, 0, 11) */,
  32'h3d13eab3 /* (0, 0, 11) */,
  32'h3d148979 /* (28, 28, 7) */,
  32'h3d250b86 /* (24, 28, 7) */,
  32'h3d66108f /* (20, 28, 7) */,
  32'h3d66e7bc /* (16, 28, 7) */,
  32'h3d66108f /* (12, 28, 7) */,
  32'h3d250b86 /* (8, 28, 7) */,
  32'h3d148979 /* (4, 28, 7) */,
  32'h3d1879c9 /* (0, 28, 7) */,
  32'h3d250b86 /* (28, 24, 7) */,
  32'h3d54dbd1 /* (24, 24, 7) */,
  32'h3da58a7f /* (20, 24, 7) */,
  32'h3db1ba44 /* (16, 24, 7) */,
  32'h3da58a7f /* (12, 24, 7) */,
  32'h3d54dbd1 /* (8, 24, 7) */,
  32'h3d250b86 /* (4, 24, 7) */,
  32'h3d1b34b2 /* (0, 24, 7) */,
  32'h3d66108f /* (28, 20, 7) */,
  32'h3da58a7f /* (24, 20, 7) */,
  32'h3e0e8e1e /* (20, 20, 7) */,
  32'h3e24eefd /* (16, 20, 7) */,
  32'h3e0e8e1e /* (12, 20, 7) */,
  32'h3da58a7f /* (8, 20, 7) */,
  32'h3d66108f /* (4, 20, 7) */,
  32'h3d4d39f8 /* (0, 20, 7) */,
  32'h3d66e7bc /* (28, 16, 7) */,
  32'h3db1ba44 /* (24, 16, 7) */,
  32'h3e24eefd /* (20, 16, 7) */,
  32'h3e4b7c7a /* (16, 16, 7) */,
  32'h3e24eefd /* (12, 16, 7) */,
  32'h3db1ba44 /* (8, 16, 7) */,
  32'h3d66e7bc /* (4, 16, 7) */,
  32'h3d482f92 /* (0, 16, 7) */,
  32'h3d66108f /* (28, 12, 7) */,
  32'h3da58a7f /* (24, 12, 7) */,
  32'h3e0e8e1e /* (20, 12, 7) */,
  32'h3e24eefd /* (16, 12, 7) */,
  32'h3e0e8e1e /* (12, 12, 7) */,
  32'h3da58a7f /* (8, 12, 7) */,
  32'h3d66108f /* (4, 12, 7) */,
  32'h3d4d39f8 /* (0, 12, 7) */,
  32'h3d250b86 /* (28, 8, 7) */,
  32'h3d54dbd1 /* (24, 8, 7) */,
  32'h3da58a7f /* (20, 8, 7) */,
  32'h3db1ba44 /* (16, 8, 7) */,
  32'h3da58a7f /* (12, 8, 7) */,
  32'h3d54dbd1 /* (8, 8, 7) */,
  32'h3d250b86 /* (4, 8, 7) */,
  32'h3d1b34b2 /* (0, 8, 7) */,
  32'h3d148979 /* (28, 4, 7) */,
  32'h3d250b86 /* (24, 4, 7) */,
  32'h3d66108f /* (20, 4, 7) */,
  32'h3d66e7bc /* (16, 4, 7) */,
  32'h3d66108f /* (12, 4, 7) */,
  32'h3d250b86 /* (8, 4, 7) */,
  32'h3d148979 /* (4, 4, 7) */,
  32'h3d1879c9 /* (0, 4, 7) */,
  32'h3d1879c9 /* (28, 0, 7) */,
  32'h3d1b34b2 /* (24, 0, 7) */,
  32'h3d4d39f8 /* (20, 0, 7) */,
  32'h3d482f92 /* (16, 0, 7) */,
  32'h3d4d39f8 /* (12, 0, 7) */,
  32'h3d1b34b2 /* (8, 0, 7) */,
  32'h3d1879c9 /* (4, 0, 7) */,
  32'h3d269d45 /* (0, 0, 7) */,
  32'h3d358b49 /* (28, 28, 3) */,
  32'h3d13fed6 /* (24, 28, 3) */,
  32'h3d30047a /* (20, 28, 3) */,
  32'h3d232f37 /* (16, 28, 3) */,
  32'h3d30047a /* (12, 28, 3) */,
  32'h3d13fed6 /* (8, 28, 3) */,
  32'h3d358b49 /* (4, 28, 3) */,
  32'h3d7541a2 /* (0, 28, 3) */,
  32'h3d13fed6 /* (28, 24, 3) */,
  32'h3d2a2238 /* (24, 24, 3) */,
  32'h3d729483 /* (20, 24, 3) */,
  32'h3d76a38f /* (16, 24, 3) */,
  32'h3d729483 /* (12, 24, 3) */,
  32'h3d2a2238 /* (8, 24, 3) */,
  32'h3d13fed6 /* (4, 24, 3) */,
  32'h3d14a194 /* (0, 24, 3) */,
  32'h3d30047a /* (28, 20, 3) */,
  32'h3d729483 /* (24, 20, 3) */,
  32'h3dc823b1 /* (20, 20, 3) */,
  32'h3de007f6 /* (16, 20, 3) */,
  32'h3dc823b1 /* (12, 20, 3) */,
  32'h3d729483 /* (8, 20, 3) */,
  32'h3d30047a /* (4, 20, 3) */,
  32'h3d202826 /* (0, 20, 3) */,
  32'h3d232f37 /* (28, 16, 3) */,
  32'h3d76a38f /* (24, 16, 3) */,
  32'h3de007f6 /* (20, 16, 3) */,
  32'h3e078d5a /* (16, 16, 3) */,
  32'h3de007f6 /* (12, 16, 3) */,
  32'h3d76a38f /* (8, 16, 3) */,
  32'h3d232f37 /* (4, 16, 3) */,
  32'h3d0e89f8 /* (0, 16, 3) */,
  32'h3d30047a /* (28, 12, 3) */,
  32'h3d729483 /* (24, 12, 3) */,
  32'h3dc823b1 /* (20, 12, 3) */,
  32'h3de007f6 /* (16, 12, 3) */,
  32'h3dc823b1 /* (12, 12, 3) */,
  32'h3d729483 /* (8, 12, 3) */,
  32'h3d30047a /* (4, 12, 3) */,
  32'h3d202826 /* (0, 12, 3) */,
  32'h3d13fed6 /* (28, 8, 3) */,
  32'h3d2a2238 /* (24, 8, 3) */,
  32'h3d729483 /* (20, 8, 3) */,
  32'h3d76a38f /* (16, 8, 3) */,
  32'h3d729483 /* (12, 8, 3) */,
  32'h3d2a2238 /* (8, 8, 3) */,
  32'h3d13fed6 /* (4, 8, 3) */,
  32'h3d14a194 /* (0, 8, 3) */,
  32'h3d358b49 /* (28, 4, 3) */,
  32'h3d13fed6 /* (24, 4, 3) */,
  32'h3d30047a /* (20, 4, 3) */,
  32'h3d232f37 /* (16, 4, 3) */,
  32'h3d30047a /* (12, 4, 3) */,
  32'h3d13fed6 /* (8, 4, 3) */,
  32'h3d358b49 /* (4, 4, 3) */,
  32'h3d7541a2 /* (0, 4, 3) */,
  32'h3d7541a2 /* (28, 0, 3) */,
  32'h3d14a194 /* (24, 0, 3) */,
  32'h3d202826 /* (20, 0, 3) */,
  32'h3d0e89f8 /* (16, 0, 3) */,
  32'h3d202826 /* (12, 0, 3) */,
  32'h3d14a194 /* (8, 0, 3) */,
  32'h3d7541a2 /* (4, 0, 3) */,
  32'h3e0c4c59 /* (0, 0, 3) */,
  32'h3e4aeee2 /* (31, 31, 30) */,
  32'h3d59109a /* (27, 31, 30) */,
  32'h3d11c69f /* (23, 31, 30) */,
  32'h3d214ba3 /* (19, 31, 30) */,
  32'h3d1a0745 /* (15, 31, 30) */,
  32'h3d16ed42 /* (11, 31, 30) */,
  32'h3d20a35e /* (7, 31, 30) */,
  32'h3dbfa8df /* (3, 31, 30) */,
  32'h3d59109a /* (31, 27, 30) */,
  32'h3d213c91 /* (27, 27, 30) */,
  32'h3d18622e /* (23, 27, 30) */,
  32'h3d3d84de /* (19, 27, 30) */,
  32'h3d3a7be5 /* (15, 27, 30) */,
  32'h3d29823f /* (11, 27, 30) */,
  32'h3d14b1c0 /* (7, 27, 30) */,
  32'h3d3cd255 /* (3, 27, 30) */,
  32'h3d11c69f /* (31, 23, 30) */,
  32'h3d18622e /* (27, 23, 30) */,
  32'h3d42665b /* (23, 23, 30) */,
  32'h3d8e358b /* (19, 23, 30) */,
  32'h3d9314c2 /* (15, 23, 30) */,
  32'h3d6d9fa3 /* (11, 23, 30) */,
  32'h3d26a1b5 /* (7, 23, 30) */,
  32'h3d12f42a /* (3, 23, 30) */,
  32'h3d214ba3 /* (31, 19, 30) */,
  32'h3d3d84de /* (27, 19, 30) */,
  32'h3d8e358b /* (23, 19, 30) */,
  32'h3dec70da /* (19, 19, 30) */,
  32'h3e003b1e /* (15, 19, 30) */,
  32'h3dba5db4 /* (11, 19, 30) */,
  32'h3d6129ae /* (7, 19, 30) */,
  32'h3d29e985 /* (3, 19, 30) */,
  32'h3d1a0745 /* (31, 15, 30) */,
  32'h3d3a7be5 /* (27, 15, 30) */,
  32'h3d9314c2 /* (23, 15, 30) */,
  32'h3e003b1e /* (19, 15, 30) */,
  32'h3e0de5f8 /* (15, 15, 30) */,
  32'h3dc59b81 /* (11, 15, 30) */,
  32'h3d62f778 /* (7, 15, 30) */,
  32'h3d240321 /* (3, 15, 30) */,
  32'h3d16ed42 /* (31, 11, 30) */,
  32'h3d29823f /* (27, 11, 30) */,
  32'h3d6d9fa3 /* (23, 11, 30) */,
  32'h3dba5db4 /* (19, 11, 30) */,
  32'h3dc59b81 /* (15, 11, 30) */,
  32'h3d96eb50 /* (11, 11, 30) */,
  32'h3d42a7b8 /* (7, 11, 30) */,
  32'h3d1c5f03 /* (3, 11, 30) */,
  32'h3d20a35e /* (31, 7, 30) */,
  32'h3d14b1c0 /* (27, 7, 30) */,
  32'h3d26a1b5 /* (23, 7, 30) */,
  32'h3d6129ae /* (19, 7, 30) */,
  32'h3d62f778 /* (15, 7, 30) */,
  32'h3d42a7b8 /* (11, 7, 30) */,
  32'h3d1777c7 /* (7, 7, 30) */,
  32'h3d1a2949 /* (3, 7, 30) */,
  32'h3dbfa8df /* (31, 3, 30) */,
  32'h3d3cd255 /* (27, 3, 30) */,
  32'h3d12f42a /* (23, 3, 30) */,
  32'h3d29e985 /* (19, 3, 30) */,
  32'h3d240321 /* (15, 3, 30) */,
  32'h3d1c5f03 /* (11, 3, 30) */,
  32'h3d1a2949 /* (7, 3, 30) */,
  32'h3d866355 /* (3, 3, 30) */,
  32'h3d3c9698 /* (31, 31, 26) */,
  32'h3d1a8b5a /* (27, 31, 26) */,
  32'h3d1c53e8 /* (23, 31, 26) */,
  32'h3d4876ff /* (19, 31, 26) */,
  32'h3d46f53f /* (15, 31, 26) */,
  32'h3d31191b /* (11, 31, 26) */,
  32'h3d146a43 /* (7, 31, 26) */,
  32'h3d2ba889 /* (3, 31, 26) */,
  32'h3d1a8b5a /* (31, 27, 26) */,
  32'h3d14f7ce /* (27, 27, 26) */,
  32'h3d2db0cc /* (23, 27, 26) */,
  32'h3d700ffa /* (19, 27, 26) */,
  32'h3d73b16f /* (15, 27, 26) */,
  32'h3d4d9045 /* (11, 27, 26) */,
  32'h3d1b2471 /* (7, 27, 26) */,
  32'h3d16d305 /* (3, 27, 26) */,
  32'h3d1c53e8 /* (31, 23, 26) */,
  32'h3d2db0cc /* (27, 23, 26) */,
  32'h3d6fd024 /* (23, 23, 26) */,
  32'h3db9d5f4 /* (19, 23, 26) */,
  32'h3dc42ad0 /* (15, 23, 26) */,
  32'h3d9750ce /* (11, 23, 26) */,
  32'h3d45eb5b /* (7, 23, 26) */,
  32'h3d215063 /* (3, 23, 26) */,
  32'h3d4876ff /* (31, 19, 26) */,
  32'h3d700ffa /* (27, 19, 26) */,
  32'h3db9d5f4 /* (23, 19, 26) */,
  32'h3e1f113d /* (19, 19, 26) */,
  32'h3e2ea39a /* (15, 19, 26) */,
  32'h3df74dbc /* (11, 19, 26) */,
  32'h3d90c8a7 /* (7, 19, 26) */,
  32'h3d54a03b /* (3, 19, 26) */,
  32'h3d46f53f /* (31, 15, 26) */,
  32'h3d73b16f /* (27, 15, 26) */,
  32'h3dc42ad0 /* (23, 15, 26) */,
  32'h3e2ea39a /* (19, 15, 26) */,
  32'h3e430b11 /* (15, 15, 26) */,
  32'h3e0533d0 /* (11, 15, 26) */,
  32'h3d95be73 /* (7, 15, 26) */,
  32'h3d54ba37 /* (3, 15, 26) */,
  32'h3d31191b /* (31, 11, 26) */,
  32'h3d4d9045 /* (27, 11, 26) */,
  32'h3d9750ce /* (23, 11, 26) */,
  32'h3df74dbc /* (19, 11, 26) */,
  32'h3e0533d0 /* (15, 11, 26) */,
  32'h3dc480ba /* (11, 11, 26) */,
  32'h3d71ecf9 /* (7, 11, 26) */,
  32'h3d39bb76 /* (3, 11, 26) */,
  32'h3d146a43 /* (31, 7, 26) */,
  32'h3d1b2471 /* (27, 7, 26) */,
  32'h3d45eb5b /* (23, 7, 26) */,
  32'h3d90c8a7 /* (19, 7, 26) */,
  32'h3d95be73 /* (15, 7, 26) */,
  32'h3d71ecf9 /* (11, 7, 26) */,
  32'h3d29a602 /* (7, 7, 26) */,
  32'h3d159d44 /* (3, 7, 26) */,
  32'h3d2ba889 /* (31, 3, 26) */,
  32'h3d16d305 /* (27, 3, 26) */,
  32'h3d215063 /* (23, 3, 26) */,
  32'h3d54a03b /* (19, 3, 26) */,
  32'h3d54ba37 /* (15, 3, 26) */,
  32'h3d39bb76 /* (11, 3, 26) */,
  32'h3d159d44 /* (7, 3, 26) */,
  32'h3d211f1b /* (3, 3, 26) */,
  32'h3d119771 /* (31, 31, 22) */,
  32'h3d1d9589 /* (27, 31, 22) */,
  32'h3d52081f /* (23, 31, 22) */,
  32'h3d9e7894 /* (19, 31, 22) */,
  32'h3da5ac70 /* (15, 31, 22) */,
  32'h3d829849 /* (11, 31, 22) */,
  32'h3d305430 /* (7, 31, 22) */,
  32'h3d14c0fd /* (3, 31, 22) */,
  32'h3d1d9589 /* (31, 27, 22) */,
  32'h3d30fc5a /* (27, 27, 22) */,
  32'h3d781ae6 /* (23, 27, 22) */,
  32'h3dc29629 /* (19, 27, 22) */,
  32'h3dce52e6 /* (15, 27, 22) */,
  32'h3d9d9380 /* (11, 27, 22) */,
  32'h3d4b3dc7 /* (7, 27, 22) */,
  32'h3d2344c4 /* (3, 27, 22) */,
  32'h3d52081f /* (31, 23, 22) */,
  32'h3d781ae6 /* (27, 23, 22) */,
  32'h3dbbc730 /* (23, 23, 22) */,
  32'h3e1d56b2 /* (19, 23, 22) */,
  32'h3e2b3653 /* (15, 23, 22) */,
  32'h3df71c69 /* (11, 23, 22) */,
  32'h3d94014f /* (7, 23, 22) */,
  32'h3d5dae2c /* (3, 23, 22) */,
  32'h3d9e7894 /* (31, 19, 22) */,
  32'h3dc29629 /* (27, 19, 22) */,
  32'h3e1d56b2 /* (23, 19, 22) */,
  32'h3e8cbae1 /* (19, 19, 22) */,
  32'h3e9d80fb /* (15, 19, 22) */,
  32'h3e562fb1 /* (11, 19, 22) */,
  32'h3defa49b /* (7, 19, 22) */,
  32'h3da99659 /* (3, 19, 22) */,
  32'h3da5ac70 /* (31, 15, 22) */,
  32'h3dce52e6 /* (27, 15, 22) */,
  32'h3e2b3653 /* (23, 15, 22) */,
  32'h3e9d80fb /* (19, 15, 22) */,
  32'h3eb2925b /* (15, 15, 22) */,
  32'h3e6c6ac0 /* (11, 15, 22) */,
  32'h3e009a19 /* (7, 15, 22) */,
  32'h3db22d06 /* (3, 15, 22) */,
  32'h3d829849 /* (31, 11, 22) */,
  32'h3d9d9380 /* (27, 11, 22) */,
  32'h3df71c69 /* (23, 11, 22) */,
  32'h3e562fb1 /* (19, 11, 22) */,
  32'h3e6c6ac0 /* (15, 11, 22) */,
  32'h3e257fc6 /* (11, 11, 22) */,
  32'h3dbf3f1d /* (7, 11, 22) */,
  32'h3d8ae43c /* (3, 11, 22) */,
  32'h3d305430 /* (31, 7, 22) */,
  32'h3d4b3dc7 /* (27, 7, 22) */,
  32'h3d94014f /* (23, 7, 22) */,
  32'h3defa49b /* (19, 7, 22) */,
  32'h3e009a19 /* (15, 7, 22) */,
  32'h3dbf3f1d /* (11, 7, 22) */,
  32'h3d6deb12 /* (7, 7, 22) */,
  32'h3d387393 /* (3, 7, 22) */,
  32'h3d14c0fd /* (31, 3, 22) */,
  32'h3d2344c4 /* (27, 3, 22) */,
  32'h3d5dae2c /* (23, 3, 22) */,
  32'h3da99659 /* (19, 3, 22) */,
  32'h3db22d06 /* (15, 3, 22) */,
  32'h3d8ae43c /* (11, 3, 22) */,
  32'h3d387393 /* (7, 3, 22) */,
  32'h3d18cb02 /* (3, 3, 22) */,
  32'h3d1e0bb6 /* (31, 31, 18) */,
  32'h3d3c7841 /* (27, 31, 18) */,
  32'h3d90dff9 /* (23, 31, 18) */,
  32'h3df65860 /* (19, 31, 18) */,
  32'h3e06d8bb /* (15, 31, 18) */,
  32'h3dc01db4 /* (11, 31, 18) */,
  32'h3d62906c /* (7, 31, 18) */,
  32'h3d276174 /* (3, 31, 18) */,
  32'h3d3c7841 /* (31, 27, 18) */,
  32'h3d63687e /* (27, 27, 18) */,
  32'h3db24f8e /* (23, 27, 18) */,
  32'h3e1a8d8c /* (19, 27, 18) */,
  32'h3e2a981c /* (15, 27, 18) */,
  32'h3deed79f /* (11, 27, 18) */,
  32'h3d8a0000 /* (7, 27, 18) */,
  32'h3d487174 /* (3, 27, 18) */,
  32'h3d90dff9 /* (31, 23, 18) */,
  32'h3db24f8e /* (27, 23, 18) */,
  32'h3e10cac5 /* (23, 23, 18) */,
  32'h3e821787 /* (19, 23, 18) */,
  32'h3e91e4f8 /* (15, 23, 18) */,
  32'h3e458f30 /* (11, 23, 18) */,
  32'h3ddc09d8 /* (7, 23, 18) */,
  32'h3d9b2a7b /* (3, 23, 18) */,
  32'h3df65860 /* (31, 19, 18) */,
  32'h3e1a8d8c /* (27, 19, 18) */,
  32'h3e821787 /* (23, 19, 18) */,
  32'h3ef33ce4 /* (19, 19, 18) */,
  32'h3f0af24f /* (15, 19, 18) */,
  32'h3eb517ce /* (11, 19, 18) */,
  32'h3e41f14c /* (7, 19, 18) */,
  32'h3e04d0b8 /* (3, 19, 18) */,
  32'h3e06d8bb /* (31, 15, 18) */,
  32'h3e2a981c /* (27, 15, 18) */,
  32'h3e91e4f8 /* (23, 15, 18) */,
  32'h3f0af24f /* (19, 15, 18) */,
  32'h3f202f9a /* (15, 15, 18) */,
  32'h3eccf8ff /* (11, 15, 18) */,
  32'h3e57a44b /* (7, 15, 18) */,
  32'h3e11d12f /* (3, 15, 18) */,
  32'h3dc01db4 /* (31, 11, 18) */,
  32'h3deed79f /* (27, 11, 18) */,
  32'h3e458f30 /* (23, 11, 18) */,
  32'h3eb517ce /* (19, 11, 18) */,
  32'h3eccf8ff /* (15, 11, 18) */,
  32'h3e882756 /* (11, 11, 18) */,
  32'h3e14a5c9 /* (7, 11, 18) */,
  32'h3dce7d45 /* (3, 11, 18) */,
  32'h3d62906c /* (31, 7, 18) */,
  32'h3d8a0000 /* (27, 7, 18) */,
  32'h3ddc09d8 /* (23, 7, 18) */,
  32'h3e41f14c /* (19, 7, 18) */,
  32'h3e57a44b /* (15, 7, 18) */,
  32'h3e14a5c9 /* (11, 7, 18) */,
  32'h3da8d240 /* (7, 7, 18) */,
  32'h3d71c736 /* (3, 7, 18) */,
  32'h3d276174 /* (31, 3, 18) */,
  32'h3d487174 /* (27, 3, 18) */,
  32'h3d9b2a7b /* (23, 3, 18) */,
  32'h3e04d0b8 /* (19, 3, 18) */,
  32'h3e11d12f /* (15, 3, 18) */,
  32'h3dce7d45 /* (11, 3, 18) */,
  32'h3d71c736 /* (7, 3, 18) */,
  32'h3d3188e3 /* (3, 3, 18) */,
  32'h3d1e0bb6 /* (31, 31, 14) */,
  32'h3d3c7841 /* (27, 31, 14) */,
  32'h3d90dff9 /* (23, 31, 14) */,
  32'h3df65860 /* (19, 31, 14) */,
  32'h3e06d8bb /* (15, 31, 14) */,
  32'h3dc01db4 /* (11, 31, 14) */,
  32'h3d62906c /* (7, 31, 14) */,
  32'h3d276174 /* (3, 31, 14) */,
  32'h3d3c7841 /* (31, 27, 14) */,
  32'h3d63687e /* (27, 27, 14) */,
  32'h3db24f8e /* (23, 27, 14) */,
  32'h3e1a8d8c /* (19, 27, 14) */,
  32'h3e2a981c /* (15, 27, 14) */,
  32'h3deed79f /* (11, 27, 14) */,
  32'h3d8a0000 /* (7, 27, 14) */,
  32'h3d487174 /* (3, 27, 14) */,
  32'h3d90dff9 /* (31, 23, 14) */,
  32'h3db24f8e /* (27, 23, 14) */,
  32'h3e10cac5 /* (23, 23, 14) */,
  32'h3e821787 /* (19, 23, 14) */,
  32'h3e91e4f8 /* (15, 23, 14) */,
  32'h3e458f30 /* (11, 23, 14) */,
  32'h3ddc09d8 /* (7, 23, 14) */,
  32'h3d9b2a7b /* (3, 23, 14) */,
  32'h3df65860 /* (31, 19, 14) */,
  32'h3e1a8d8c /* (27, 19, 14) */,
  32'h3e821787 /* (23, 19, 14) */,
  32'h3ef33ce4 /* (19, 19, 14) */,
  32'h3f0af24f /* (15, 19, 14) */,
  32'h3eb517ce /* (11, 19, 14) */,
  32'h3e41f14c /* (7, 19, 14) */,
  32'h3e04d0b8 /* (3, 19, 14) */,
  32'h3e06d8bb /* (31, 15, 14) */,
  32'h3e2a981c /* (27, 15, 14) */,
  32'h3e91e4f8 /* (23, 15, 14) */,
  32'h3f0af24f /* (19, 15, 14) */,
  32'h3f202f9a /* (15, 15, 14) */,
  32'h3eccf8ff /* (11, 15, 14) */,
  32'h3e57a44b /* (7, 15, 14) */,
  32'h3e11d12f /* (3, 15, 14) */,
  32'h3dc01db4 /* (31, 11, 14) */,
  32'h3deed79f /* (27, 11, 14) */,
  32'h3e458f30 /* (23, 11, 14) */,
  32'h3eb517ce /* (19, 11, 14) */,
  32'h3eccf8ff /* (15, 11, 14) */,
  32'h3e882756 /* (11, 11, 14) */,
  32'h3e14a5c9 /* (7, 11, 14) */,
  32'h3dce7d45 /* (3, 11, 14) */,
  32'h3d62906c /* (31, 7, 14) */,
  32'h3d8a0000 /* (27, 7, 14) */,
  32'h3ddc09d8 /* (23, 7, 14) */,
  32'h3e41f14c /* (19, 7, 14) */,
  32'h3e57a44b /* (15, 7, 14) */,
  32'h3e14a5c9 /* (11, 7, 14) */,
  32'h3da8d240 /* (7, 7, 14) */,
  32'h3d71c736 /* (3, 7, 14) */,
  32'h3d276174 /* (31, 3, 14) */,
  32'h3d487174 /* (27, 3, 14) */,
  32'h3d9b2a7b /* (23, 3, 14) */,
  32'h3e04d0b8 /* (19, 3, 14) */,
  32'h3e11d12f /* (15, 3, 14) */,
  32'h3dce7d45 /* (11, 3, 14) */,
  32'h3d71c736 /* (7, 3, 14) */,
  32'h3d3188e3 /* (3, 3, 14) */,
  32'h3d119771 /* (31, 31, 10) */,
  32'h3d1d9589 /* (27, 31, 10) */,
  32'h3d52081f /* (23, 31, 10) */,
  32'h3d9e7894 /* (19, 31, 10) */,
  32'h3da5ac70 /* (15, 31, 10) */,
  32'h3d829849 /* (11, 31, 10) */,
  32'h3d305430 /* (7, 31, 10) */,
  32'h3d14c0fd /* (3, 31, 10) */,
  32'h3d1d9589 /* (31, 27, 10) */,
  32'h3d30fc5a /* (27, 27, 10) */,
  32'h3d781ae6 /* (23, 27, 10) */,
  32'h3dc29629 /* (19, 27, 10) */,
  32'h3dce52e6 /* (15, 27, 10) */,
  32'h3d9d9380 /* (11, 27, 10) */,
  32'h3d4b3dc7 /* (7, 27, 10) */,
  32'h3d2344c4 /* (3, 27, 10) */,
  32'h3d52081f /* (31, 23, 10) */,
  32'h3d781ae6 /* (27, 23, 10) */,
  32'h3dbbc730 /* (23, 23, 10) */,
  32'h3e1d56b2 /* (19, 23, 10) */,
  32'h3e2b3653 /* (15, 23, 10) */,
  32'h3df71c69 /* (11, 23, 10) */,
  32'h3d94014f /* (7, 23, 10) */,
  32'h3d5dae2c /* (3, 23, 10) */,
  32'h3d9e7894 /* (31, 19, 10) */,
  32'h3dc29629 /* (27, 19, 10) */,
  32'h3e1d56b2 /* (23, 19, 10) */,
  32'h3e8cbae1 /* (19, 19, 10) */,
  32'h3e9d80fb /* (15, 19, 10) */,
  32'h3e562fb1 /* (11, 19, 10) */,
  32'h3defa49b /* (7, 19, 10) */,
  32'h3da99659 /* (3, 19, 10) */,
  32'h3da5ac70 /* (31, 15, 10) */,
  32'h3dce52e6 /* (27, 15, 10) */,
  32'h3e2b3653 /* (23, 15, 10) */,
  32'h3e9d80fb /* (19, 15, 10) */,
  32'h3eb2925b /* (15, 15, 10) */,
  32'h3e6c6ac0 /* (11, 15, 10) */,
  32'h3e009a19 /* (7, 15, 10) */,
  32'h3db22d06 /* (3, 15, 10) */,
  32'h3d829849 /* (31, 11, 10) */,
  32'h3d9d9380 /* (27, 11, 10) */,
  32'h3df71c69 /* (23, 11, 10) */,
  32'h3e562fb1 /* (19, 11, 10) */,
  32'h3e6c6ac0 /* (15, 11, 10) */,
  32'h3e257fc6 /* (11, 11, 10) */,
  32'h3dbf3f1d /* (7, 11, 10) */,
  32'h3d8ae43c /* (3, 11, 10) */,
  32'h3d305430 /* (31, 7, 10) */,
  32'h3d4b3dc7 /* (27, 7, 10) */,
  32'h3d94014f /* (23, 7, 10) */,
  32'h3defa49b /* (19, 7, 10) */,
  32'h3e009a19 /* (15, 7, 10) */,
  32'h3dbf3f1d /* (11, 7, 10) */,
  32'h3d6deb12 /* (7, 7, 10) */,
  32'h3d387393 /* (3, 7, 10) */,
  32'h3d14c0fd /* (31, 3, 10) */,
  32'h3d2344c4 /* (27, 3, 10) */,
  32'h3d5dae2c /* (23, 3, 10) */,
  32'h3da99659 /* (19, 3, 10) */,
  32'h3db22d06 /* (15, 3, 10) */,
  32'h3d8ae43c /* (11, 3, 10) */,
  32'h3d387393 /* (7, 3, 10) */,
  32'h3d18cb02 /* (3, 3, 10) */,
  32'h3d3c9698 /* (31, 31, 6) */,
  32'h3d1a8b5a /* (27, 31, 6) */,
  32'h3d1c53e8 /* (23, 31, 6) */,
  32'h3d4876ff /* (19, 31, 6) */,
  32'h3d46f53f /* (15, 31, 6) */,
  32'h3d31191b /* (11, 31, 6) */,
  32'h3d146a43 /* (7, 31, 6) */,
  32'h3d2ba889 /* (3, 31, 6) */,
  32'h3d1a8b5a /* (31, 27, 6) */,
  32'h3d14f7ce /* (27, 27, 6) */,
  32'h3d2db0cc /* (23, 27, 6) */,
  32'h3d700ffa /* (19, 27, 6) */,
  32'h3d73b16f /* (15, 27, 6) */,
  32'h3d4d9045 /* (11, 27, 6) */,
  32'h3d1b2471 /* (7, 27, 6) */,
  32'h3d16d305 /* (3, 27, 6) */,
  32'h3d1c53e8 /* (31, 23, 6) */,
  32'h3d2db0cc /* (27, 23, 6) */,
  32'h3d6fd024 /* (23, 23, 6) */,
  32'h3db9d5f4 /* (19, 23, 6) */,
  32'h3dc42ad0 /* (15, 23, 6) */,
  32'h3d9750ce /* (11, 23, 6) */,
  32'h3d45eb5b /* (7, 23, 6) */,
  32'h3d215063 /* (3, 23, 6) */,
  32'h3d4876ff /* (31, 19, 6) */,
  32'h3d700ffa /* (27, 19, 6) */,
  32'h3db9d5f4 /* (23, 19, 6) */,
  32'h3e1f113d /* (19, 19, 6) */,
  32'h3e2ea39a /* (15, 19, 6) */,
  32'h3df74dbc /* (11, 19, 6) */,
  32'h3d90c8a7 /* (7, 19, 6) */,
  32'h3d54a03b /* (3, 19, 6) */,
  32'h3d46f53f /* (31, 15, 6) */,
  32'h3d73b16f /* (27, 15, 6) */,
  32'h3dc42ad0 /* (23, 15, 6) */,
  32'h3e2ea39a /* (19, 15, 6) */,
  32'h3e430b11 /* (15, 15, 6) */,
  32'h3e0533d0 /* (11, 15, 6) */,
  32'h3d95be73 /* (7, 15, 6) */,
  32'h3d54ba37 /* (3, 15, 6) */,
  32'h3d31191b /* (31, 11, 6) */,
  32'h3d4d9045 /* (27, 11, 6) */,
  32'h3d9750ce /* (23, 11, 6) */,
  32'h3df74dbc /* (19, 11, 6) */,
  32'h3e0533d0 /* (15, 11, 6) */,
  32'h3dc480ba /* (11, 11, 6) */,
  32'h3d71ecf9 /* (7, 11, 6) */,
  32'h3d39bb76 /* (3, 11, 6) */,
  32'h3d146a43 /* (31, 7, 6) */,
  32'h3d1b2471 /* (27, 7, 6) */,
  32'h3d45eb5b /* (23, 7, 6) */,
  32'h3d90c8a7 /* (19, 7, 6) */,
  32'h3d95be73 /* (15, 7, 6) */,
  32'h3d71ecf9 /* (11, 7, 6) */,
  32'h3d29a602 /* (7, 7, 6) */,
  32'h3d159d44 /* (3, 7, 6) */,
  32'h3d2ba889 /* (31, 3, 6) */,
  32'h3d16d305 /* (27, 3, 6) */,
  32'h3d215063 /* (23, 3, 6) */,
  32'h3d54a03b /* (19, 3, 6) */,
  32'h3d54ba37 /* (15, 3, 6) */,
  32'h3d39bb76 /* (11, 3, 6) */,
  32'h3d159d44 /* (7, 3, 6) */,
  32'h3d211f1b /* (3, 3, 6) */,
  32'h3e4aeee2 /* (31, 31, 2) */,
  32'h3d59109a /* (27, 31, 2) */,
  32'h3d11c69f /* (23, 31, 2) */,
  32'h3d214ba3 /* (19, 31, 2) */,
  32'h3d1a0745 /* (15, 31, 2) */,
  32'h3d16ed42 /* (11, 31, 2) */,
  32'h3d20a35e /* (7, 31, 2) */,
  32'h3dbfa8df /* (3, 31, 2) */,
  32'h3d59109a /* (31, 27, 2) */,
  32'h3d213c91 /* (27, 27, 2) */,
  32'h3d18622e /* (23, 27, 2) */,
  32'h3d3d84de /* (19, 27, 2) */,
  32'h3d3a7be5 /* (15, 27, 2) */,
  32'h3d29823f /* (11, 27, 2) */,
  32'h3d14b1c0 /* (7, 27, 2) */,
  32'h3d3cd255 /* (3, 27, 2) */,
  32'h3d11c69f /* (31, 23, 2) */,
  32'h3d18622e /* (27, 23, 2) */,
  32'h3d42665b /* (23, 23, 2) */,
  32'h3d8e358b /* (19, 23, 2) */,
  32'h3d9314c2 /* (15, 23, 2) */,
  32'h3d6d9fa3 /* (11, 23, 2) */,
  32'h3d26a1b5 /* (7, 23, 2) */,
  32'h3d12f42a /* (3, 23, 2) */,
  32'h3d214ba3 /* (31, 19, 2) */,
  32'h3d3d84de /* (27, 19, 2) */,
  32'h3d8e358b /* (23, 19, 2) */,
  32'h3dec70da /* (19, 19, 2) */,
  32'h3e003b1e /* (15, 19, 2) */,
  32'h3dba5db4 /* (11, 19, 2) */,
  32'h3d6129ae /* (7, 19, 2) */,
  32'h3d29e985 /* (3, 19, 2) */,
  32'h3d1a0745 /* (31, 15, 2) */,
  32'h3d3a7be5 /* (27, 15, 2) */,
  32'h3d9314c2 /* (23, 15, 2) */,
  32'h3e003b1e /* (19, 15, 2) */,
  32'h3e0de5f8 /* (15, 15, 2) */,
  32'h3dc59b81 /* (11, 15, 2) */,
  32'h3d62f778 /* (7, 15, 2) */,
  32'h3d240321 /* (3, 15, 2) */,
  32'h3d16ed42 /* (31, 11, 2) */,
  32'h3d29823f /* (27, 11, 2) */,
  32'h3d6d9fa3 /* (23, 11, 2) */,
  32'h3dba5db4 /* (19, 11, 2) */,
  32'h3dc59b81 /* (15, 11, 2) */,
  32'h3d96eb50 /* (11, 11, 2) */,
  32'h3d42a7b8 /* (7, 11, 2) */,
  32'h3d1c5f03 /* (3, 11, 2) */,
  32'h3d20a35e /* (31, 7, 2) */,
  32'h3d14b1c0 /* (27, 7, 2) */,
  32'h3d26a1b5 /* (23, 7, 2) */,
  32'h3d6129ae /* (19, 7, 2) */,
  32'h3d62f778 /* (15, 7, 2) */,
  32'h3d42a7b8 /* (11, 7, 2) */,
  32'h3d1777c7 /* (7, 7, 2) */,
  32'h3d1a2949 /* (3, 7, 2) */,
  32'h3dbfa8df /* (31, 3, 2) */,
  32'h3d3cd255 /* (27, 3, 2) */,
  32'h3d12f42a /* (23, 3, 2) */,
  32'h3d29e985 /* (19, 3, 2) */,
  32'h3d240321 /* (15, 3, 2) */,
  32'h3d1c5f03 /* (11, 3, 2) */,
  32'h3d1a2949 /* (7, 3, 2) */,
  32'h3d866355 /* (3, 3, 2) */,
  32'h3e0c4d23 /* (30, 31, 30) */,
  32'h3d3543e4 /* (26, 31, 30) */,
  32'h3d12ac07 /* (22, 31, 30) */,
  32'h3d217487 /* (18, 31, 30) */,
  32'h3d217487 /* (14, 31, 30) */,
  32'h3d12ac07 /* (10, 31, 30) */,
  32'h3d3543e4 /* (6, 31, 30) */,
  32'h3e0c4d23 /* (2, 31, 30) */,
  32'h3d4ca49b /* (30, 27, 30) */,
  32'h3d18df8d /* (26, 27, 30) */,
  32'h3d1f9f49 /* (22, 27, 30) */,
  32'h3d40d8bf /* (18, 27, 30) */,
  32'h3d40d8bf /* (14, 27, 30) */,
  32'h3d1f9f49 /* (10, 27, 30) */,
  32'h3d18df8d /* (6, 27, 30) */,
  32'h3d4ca49b /* (2, 27, 30) */,
  32'h3d1214c5 /* (30, 23, 30) */,
  32'h3d1e19af /* (26, 23, 30) */,
  32'h3d56480e /* (22, 23, 30) */,
  32'h3d94a37c /* (18, 23, 30) */,
  32'h3d94a37c /* (14, 23, 30) */,
  32'h3d56480e /* (10, 23, 30) */,
  32'h3d1e19af /* (6, 23, 30) */,
  32'h3d1214c5 /* (2, 23, 30) */,
  32'h3d246fbd /* (30, 19, 30) */,
  32'h3d4ce87b /* (26, 19, 30) */,
  32'h3da2895a /* (22, 19, 30) */,
  32'h3dfd653f /* (18, 19, 30) */,
  32'h3dfd653f /* (14, 19, 30) */,
  32'h3da2895a /* (10, 19, 30) */,
  32'h3d4ce87b /* (6, 19, 30) */,
  32'h3d246fbd /* (2, 19, 30) */,
  32'h3d1dadb9 /* (30, 15, 30) */,
  32'h3d4bfe66 /* (26, 15, 30) */,
  32'h3daa3ec9 /* (22, 15, 30) */,
  32'h3e0adb0d /* (18, 15, 30) */,
  32'h3e0adb0d /* (14, 15, 30) */,
  32'h3daa3ec9 /* (10, 15, 30) */,
  32'h3d4bfe66 /* (6, 15, 30) */,
  32'h3d1dadb9 /* (2, 15, 30) */,
  32'h3d18e0f8 /* (30, 11, 30) */,
  32'h3d343ccb /* (26, 11, 30) */,
  32'h3d85a0b3 /* (22, 11, 30) */,
  32'h3dc55f41 /* (18, 11, 30) */,
  32'h3dc55f41 /* (14, 11, 30) */,
  32'h3d85a0b3 /* (10, 11, 30) */,
  32'h3d343ccb /* (6, 11, 30) */,
  32'h3d18e0f8 /* (2, 11, 30) */,
  32'h3d1dd271 /* (30, 7, 30) */,
  32'h3d14b9d3 /* (26, 7, 30) */,
  32'h3d3346c6 /* (22, 7, 30) */,
  32'h3d6820b1 /* (18, 7, 30) */,
  32'h3d6820b1 /* (14, 7, 30) */,
  32'h3d3346c6 /* (10, 7, 30) */,
  32'h3d14b9d3 /* (6, 7, 30) */,
  32'h3d1dd271 /* (2, 7, 30) */,
  32'h3da3af74 /* (30, 3, 30) */,
  32'h3d271e8d /* (26, 3, 30) */,
  32'h3d162b76 /* (22, 3, 30) */,
  32'h3d2b1735 /* (18, 3, 30) */,
  32'h3d2b1735 /* (14, 3, 30) */,
  32'h3d162b76 /* (10, 3, 30) */,
  32'h3d271e8d /* (6, 3, 30) */,
  32'h3da3af74 /* (2, 3, 30) */,
  32'h3d3543e4 /* (30, 31, 26) */,
  32'h3d15cc97 /* (26, 31, 26) */,
  32'h3d2567ce /* (22, 31, 26) */,
  32'h3d4cf093 /* (18, 31, 26) */,
  32'h3d4cf093 /* (14, 31, 26) */,
  32'h3d2567ce /* (10, 31, 26) */,
  32'h3d15cc97 /* (6, 31, 26) */,
  32'h3d3543e4 /* (2, 31, 26) */,
  32'h3d18df8d /* (30, 27, 26) */,
  32'h3d16bb8b /* (26, 27, 26) */,
  32'h3d3c300c /* (22, 27, 26) */,
  32'h3d786cd6 /* (18, 27, 26) */,
  32'h3d786cd6 /* (14, 27, 26) */,
  32'h3d3c300c /* (10, 27, 26) */,
  32'h3d16bb8b /* (6, 27, 26) */,
  32'h3d18df8d /* (2, 27, 26) */,
  32'h3d1e19af /* (30, 23, 26) */,
  32'h3d37f9d0 /* (26, 23, 26) */,
  32'h3d866682 /* (22, 23, 26) */,
  32'h3dc45939 /* (18, 23, 26) */,
  32'h3dc45939 /* (14, 23, 26) */,
  32'h3d866682 /* (10, 23, 26) */,
  32'h3d37f9d0 /* (6, 23, 26) */,
  32'h3d1e19af /* (2, 23, 26) */,
  32'h3d4ce87b /* (30, 19, 26) */,
  32'h3d82bc35 /* (26, 19, 26) */,
  32'h3dd610ea /* (22, 19, 26) */,
  32'h3e2b8c37 /* (18, 19, 26) */,
  32'h3e2b8c37 /* (14, 19, 26) */,
  32'h3dd610ea /* (10, 19, 26) */,
  32'h3d82bc35 /* (6, 19, 26) */,
  32'h3d4ce87b /* (2, 19, 26) */,
  32'h3d4bfe66 /* (30, 15, 26) */,
  32'h3d85e8bf /* (26, 15, 26) */,
  32'h3de44bb3 /* (22, 15, 26) */,
  32'h3e3e01e0 /* (18, 15, 26) */,
  32'h3e3e01e0 /* (14, 15, 26) */,
  32'h3de44bb3 /* (10, 15, 26) */,
  32'h3d85e8bf /* (6, 15, 26) */,
  32'h3d4bfe66 /* (2, 15, 26) */,
  32'h3d343ccb /* (30, 11, 26) */,
  32'h3d5d3b5c /* (26, 11, 26) */,
  32'h3dac23aa /* (22, 11, 26) */,
  32'h3e040b60 /* (18, 11, 26) */,
  32'h3e040b60 /* (14, 11, 26) */,
  32'h3dac23aa /* (10, 11, 26) */,
  32'h3d5d3b5c /* (6, 11, 26) */,
  32'h3d343ccb /* (2, 11, 26) */,
  32'h3d14b9d3 /* (30, 7, 26) */,
  32'h3d20f672 /* (26, 7, 26) */,
  32'h3d5a2934 /* (22, 7, 26) */,
  32'h3d975464 /* (18, 7, 26) */,
  32'h3d975464 /* (14, 7, 26) */,
  32'h3d5a2934 /* (10, 7, 26) */,
  32'h3d20f672 /* (6, 7, 26) */,
  32'h3d14b9d3 /* (2, 7, 26) */,
  32'h3d271e8d /* (30, 3, 26) */,
  32'h3d14c14d /* (26, 3, 26) */,
  32'h3d2c3293 /* (22, 3, 26) */,
  32'h3d5a5169 /* (18, 3, 26) */,
  32'h3d5a5169 /* (14, 3, 26) */,
  32'h3d2c3293 /* (10, 3, 26) */,
  32'h3d14c14d /* (6, 3, 26) */,
  32'h3d271e8d /* (2, 3, 26) */,
  32'h3d12ac07 /* (30, 31, 22) */,
  32'h3d2567ce /* (26, 31, 22) */,
  32'h3d699f13 /* (22, 31, 22) */,
  32'h3da6958f /* (18, 31, 22) */,
  32'h3da6958f /* (14, 31, 22) */,
  32'h3d699f13 /* (10, 31, 22) */,
  32'h3d2567ce /* (6, 31, 22) */,
  32'h3d12ac07 /* (2, 31, 22) */,
  32'h3d1f9f49 /* (30, 27, 22) */,
  32'h3d3c300c /* (26, 27, 22) */,
  32'h3d8b85a2 /* (22, 27, 22) */,
  32'h3dce13fe /* (18, 27, 22) */,
  32'h3dce13fe /* (14, 27, 22) */,
  32'h3d8b85a2 /* (10, 27, 22) */,
  32'h3d3c300c /* (6, 27, 22) */,
  32'h3d1f9f49 /* (2, 27, 22) */,
  32'h3d56480e /* (30, 23, 22) */,
  32'h3d866682 /* (26, 23, 22) */,
  32'h3dd7137d /* (22, 23, 22) */,
  32'h3e28e750 /* (18, 23, 22) */,
  32'h3e28e750 /* (14, 23, 22) */,
  32'h3dd7137d /* (10, 23, 22) */,
  32'h3d866682 /* (6, 23, 22) */,
  32'h3d56480e /* (2, 23, 22) */,
  32'h3da2895a /* (30, 19, 22) */,
  32'h3dd610ea /* (26, 19, 22) */,
  32'h3e37540b /* (22, 19, 22) */,
  32'h3e994798 /* (18, 19, 22) */,
  32'h3e994798 /* (14, 19, 22) */,
  32'h3e37540b /* (10, 19, 22) */,
  32'h3dd610ea /* (6, 19, 22) */,
  32'h3da2895a /* (2, 19, 22) */,
  32'h3daa3ec9 /* (30, 15, 22) */,
  32'h3de44bb3 /* (26, 15, 22) */,
  32'h3e48eba4 /* (22, 15, 22) */,
  32'h3eacaf9b /* (18, 15, 22) */,
  32'h3eacaf9b /* (14, 15, 22) */,
  32'h3e48eba4 /* (10, 15, 22) */,
  32'h3de44bb3 /* (6, 15, 22) */,
  32'h3daa3ec9 /* (2, 15, 22) */,
  32'h3d85a0b3 /* (30, 11, 22) */,
  32'h3dac23aa /* (26, 11, 22) */,
  32'h3e0ecbcd /* (22, 11, 22) */,
  32'h3e67a191 /* (18, 11, 22) */,
  32'h3e67a191 /* (14, 11, 22) */,
  32'h3e0ecbcd /* (10, 11, 22) */,
  32'h3dac23aa /* (6, 11, 22) */,
  32'h3d85a0b3 /* (2, 11, 22) */,
  32'h3d3346c6 /* (30, 7, 22) */,
  32'h3d5a2934 /* (26, 7, 22) */,
  32'h3da7f0fb /* (22, 7, 22) */,
  32'h3dff6ab3 /* (18, 7, 22) */,
  32'h3dff6ab3 /* (14, 7, 22) */,
  32'h3da7f0fb /* (10, 7, 22) */,
  32'h3d5a2934 /* (6, 7, 22) */,
  32'h3d3346c6 /* (2, 7, 22) */,
  32'h3d162b76 /* (30, 3, 22) */,
  32'h3d2c3293 /* (26, 3, 22) */,
  32'h3d77904c /* (22, 3, 22) */,
  32'h3db2bcb9 /* (18, 3, 22) */,
  32'h3db2bcb9 /* (14, 3, 22) */,
  32'h3d77904c /* (10, 3, 22) */,
  32'h3d2c3293 /* (6, 3, 22) */,
  32'h3d162b76 /* (2, 3, 22) */,
  32'h3d217487 /* (30, 31, 18) */,
  32'h3d4cf093 /* (26, 31, 18) */,
  32'h3da6958f /* (22, 31, 18) */,
  32'h3e04a438 /* (18, 31, 18) */,
  32'h3e04a438 /* (14, 31, 18) */,
  32'h3da6958f /* (10, 31, 18) */,
  32'h3d4cf093 /* (6, 31, 18) */,
  32'h3d217487 /* (2, 31, 18) */,
  32'h3d40d8bf /* (30, 27, 18) */,
  32'h3d786cd6 /* (26, 27, 18) */,
  32'h3dce13fe /* (22, 27, 18) */,
  32'h3e27240a /* (18, 27, 18) */,
  32'h3e27240a /* (14, 27, 18) */,
  32'h3dce13fe /* (10, 27, 18) */,
  32'h3d786cd6 /* (6, 27, 18) */,
  32'h3d40d8bf /* (2, 27, 18) */,
  32'h3d94a37c /* (30, 23, 18) */,
  32'h3dc45939 /* (26, 23, 18) */,
  32'h3e28e750 /* (22, 23, 18) */,
  32'h3e8dd733 /* (18, 23, 18) */,
  32'h3e8dd733 /* (14, 23, 18) */,
  32'h3e28e750 /* (10, 23, 18) */,
  32'h3dc45939 /* (6, 23, 18) */,
  32'h3d94a37c /* (2, 23, 18) */,
  32'h3dfd653f /* (30, 19, 18) */,
  32'h3e2b8c37 /* (26, 19, 18) */,
  32'h3e994798 /* (22, 19, 18) */,
  32'h3f05dc96 /* (18, 19, 18) */,
  32'h3f05dc96 /* (14, 19, 18) */,
  32'h3e994798 /* (10, 19, 18) */,
  32'h3e2b8c37 /* (6, 19, 18) */,
  32'h3dfd653f /* (2, 19, 18) */,
  32'h3e0adb0d /* (30, 15, 18) */,
  32'h3e3e01e0 /* (26, 15, 18) */,
  32'h3eacaf9b /* (22, 15, 18) */,
  32'h3f19a2a7 /* (18, 15, 18) */,
  32'h3f19a2a7 /* (14, 15, 18) */,
  32'h3eacaf9b /* (10, 15, 18) */,
  32'h3e3e01e0 /* (6, 15, 18) */,
  32'h3e0adb0d /* (2, 15, 18) */,
  32'h3dc55f41 /* (30, 11, 18) */,
  32'h3e040b60 /* (26, 11, 18) */,
  32'h3e67a191 /* (22, 11, 18) */,
  32'h3ec66134 /* (18, 11, 18) */,
  32'h3ec66134 /* (14, 11, 18) */,
  32'h3e67a191 /* (10, 11, 18) */,
  32'h3e040b60 /* (6, 11, 18) */,
  32'h3dc55f41 /* (2, 11, 18) */,
  32'h3d6820b1 /* (30, 7, 18) */,
  32'h3d975464 /* (26, 7, 18) */,
  32'h3dff6ab3 /* (22, 7, 18) */,
  32'h3e528761 /* (18, 7, 18) */,
  32'h3e528761 /* (14, 7, 18) */,
  32'h3dff6ab3 /* (10, 7, 18) */,
  32'h3d975464 /* (6, 7, 18) */,
  32'h3d6820b1 /* (2, 7, 18) */,
  32'h3d2b1735 /* (30, 3, 18) */,
  32'h3d5a5169 /* (26, 3, 18) */,
  32'h3db2bcb9 /* (22, 3, 18) */,
  32'h3e0f3c67 /* (18, 3, 18) */,
  32'h3e0f3c67 /* (14, 3, 18) */,
  32'h3db2bcb9 /* (10, 3, 18) */,
  32'h3d5a5169 /* (6, 3, 18) */,
  32'h3d2b1735 /* (2, 3, 18) */,
  32'h3d217487 /* (30, 31, 14) */,
  32'h3d4cf093 /* (26, 31, 14) */,
  32'h3da6958f /* (22, 31, 14) */,
  32'h3e04a438 /* (18, 31, 14) */,
  32'h3e04a438 /* (14, 31, 14) */,
  32'h3da6958f /* (10, 31, 14) */,
  32'h3d4cf093 /* (6, 31, 14) */,
  32'h3d217487 /* (2, 31, 14) */,
  32'h3d40d8bf /* (30, 27, 14) */,
  32'h3d786cd6 /* (26, 27, 14) */,
  32'h3dce13fe /* (22, 27, 14) */,
  32'h3e27240a /* (18, 27, 14) */,
  32'h3e27240a /* (14, 27, 14) */,
  32'h3dce13fe /* (10, 27, 14) */,
  32'h3d786cd6 /* (6, 27, 14) */,
  32'h3d40d8bf /* (2, 27, 14) */,
  32'h3d94a37c /* (30, 23, 14) */,
  32'h3dc45939 /* (26, 23, 14) */,
  32'h3e28e750 /* (22, 23, 14) */,
  32'h3e8dd733 /* (18, 23, 14) */,
  32'h3e8dd733 /* (14, 23, 14) */,
  32'h3e28e750 /* (10, 23, 14) */,
  32'h3dc45939 /* (6, 23, 14) */,
  32'h3d94a37c /* (2, 23, 14) */,
  32'h3dfd653f /* (30, 19, 14) */,
  32'h3e2b8c37 /* (26, 19, 14) */,
  32'h3e994798 /* (22, 19, 14) */,
  32'h3f05dc96 /* (18, 19, 14) */,
  32'h3f05dc96 /* (14, 19, 14) */,
  32'h3e994798 /* (10, 19, 14) */,
  32'h3e2b8c37 /* (6, 19, 14) */,
  32'h3dfd653f /* (2, 19, 14) */,
  32'h3e0adb0d /* (30, 15, 14) */,
  32'h3e3e01e0 /* (26, 15, 14) */,
  32'h3eacaf9b /* (22, 15, 14) */,
  32'h3f19a2a7 /* (18, 15, 14) */,
  32'h3f19a2a7 /* (14, 15, 14) */,
  32'h3eacaf9b /* (10, 15, 14) */,
  32'h3e3e01e0 /* (6, 15, 14) */,
  32'h3e0adb0d /* (2, 15, 14) */,
  32'h3dc55f41 /* (30, 11, 14) */,
  32'h3e040b60 /* (26, 11, 14) */,
  32'h3e67a191 /* (22, 11, 14) */,
  32'h3ec66134 /* (18, 11, 14) */,
  32'h3ec66134 /* (14, 11, 14) */,
  32'h3e67a191 /* (10, 11, 14) */,
  32'h3e040b60 /* (6, 11, 14) */,
  32'h3dc55f41 /* (2, 11, 14) */,
  32'h3d6820b1 /* (30, 7, 14) */,
  32'h3d975464 /* (26, 7, 14) */,
  32'h3dff6ab3 /* (22, 7, 14) */,
  32'h3e528761 /* (18, 7, 14) */,
  32'h3e528761 /* (14, 7, 14) */,
  32'h3dff6ab3 /* (10, 7, 14) */,
  32'h3d975464 /* (6, 7, 14) */,
  32'h3d6820b1 /* (2, 7, 14) */,
  32'h3d2b1735 /* (30, 3, 14) */,
  32'h3d5a5169 /* (26, 3, 14) */,
  32'h3db2bcb9 /* (22, 3, 14) */,
  32'h3e0f3c67 /* (18, 3, 14) */,
  32'h3e0f3c67 /* (14, 3, 14) */,
  32'h3db2bcb9 /* (10, 3, 14) */,
  32'h3d5a5169 /* (6, 3, 14) */,
  32'h3d2b1735 /* (2, 3, 14) */,
  32'h3d12ac07 /* (30, 31, 10) */,
  32'h3d2567ce /* (26, 31, 10) */,
  32'h3d699f13 /* (22, 31, 10) */,
  32'h3da6958f /* (18, 31, 10) */,
  32'h3da6958f /* (14, 31, 10) */,
  32'h3d699f13 /* (10, 31, 10) */,
  32'h3d2567ce /* (6, 31, 10) */,
  32'h3d12ac07 /* (2, 31, 10) */,
  32'h3d1f9f49 /* (30, 27, 10) */,
  32'h3d3c300c /* (26, 27, 10) */,
  32'h3d8b85a2 /* (22, 27, 10) */,
  32'h3dce13fe /* (18, 27, 10) */,
  32'h3dce13fe /* (14, 27, 10) */,
  32'h3d8b85a2 /* (10, 27, 10) */,
  32'h3d3c300c /* (6, 27, 10) */,
  32'h3d1f9f49 /* (2, 27, 10) */,
  32'h3d56480e /* (30, 23, 10) */,
  32'h3d866682 /* (26, 23, 10) */,
  32'h3dd7137d /* (22, 23, 10) */,
  32'h3e28e750 /* (18, 23, 10) */,
  32'h3e28e750 /* (14, 23, 10) */,
  32'h3dd7137d /* (10, 23, 10) */,
  32'h3d866682 /* (6, 23, 10) */,
  32'h3d56480e /* (2, 23, 10) */,
  32'h3da2895a /* (30, 19, 10) */,
  32'h3dd610ea /* (26, 19, 10) */,
  32'h3e37540b /* (22, 19, 10) */,
  32'h3e994798 /* (18, 19, 10) */,
  32'h3e994798 /* (14, 19, 10) */,
  32'h3e37540b /* (10, 19, 10) */,
  32'h3dd610ea /* (6, 19, 10) */,
  32'h3da2895a /* (2, 19, 10) */,
  32'h3daa3ec9 /* (30, 15, 10) */,
  32'h3de44bb3 /* (26, 15, 10) */,
  32'h3e48eba4 /* (22, 15, 10) */,
  32'h3eacaf9b /* (18, 15, 10) */,
  32'h3eacaf9b /* (14, 15, 10) */,
  32'h3e48eba4 /* (10, 15, 10) */,
  32'h3de44bb3 /* (6, 15, 10) */,
  32'h3daa3ec9 /* (2, 15, 10) */,
  32'h3d85a0b3 /* (30, 11, 10) */,
  32'h3dac23aa /* (26, 11, 10) */,
  32'h3e0ecbcd /* (22, 11, 10) */,
  32'h3e67a191 /* (18, 11, 10) */,
  32'h3e67a191 /* (14, 11, 10) */,
  32'h3e0ecbcd /* (10, 11, 10) */,
  32'h3dac23aa /* (6, 11, 10) */,
  32'h3d85a0b3 /* (2, 11, 10) */,
  32'h3d3346c6 /* (30, 7, 10) */,
  32'h3d5a2934 /* (26, 7, 10) */,
  32'h3da7f0fb /* (22, 7, 10) */,
  32'h3dff6ab3 /* (18, 7, 10) */,
  32'h3dff6ab3 /* (14, 7, 10) */,
  32'h3da7f0fb /* (10, 7, 10) */,
  32'h3d5a2934 /* (6, 7, 10) */,
  32'h3d3346c6 /* (2, 7, 10) */,
  32'h3d162b76 /* (30, 3, 10) */,
  32'h3d2c3293 /* (26, 3, 10) */,
  32'h3d77904c /* (22, 3, 10) */,
  32'h3db2bcb9 /* (18, 3, 10) */,
  32'h3db2bcb9 /* (14, 3, 10) */,
  32'h3d77904c /* (10, 3, 10) */,
  32'h3d2c3293 /* (6, 3, 10) */,
  32'h3d162b76 /* (2, 3, 10) */,
  32'h3d3543e4 /* (30, 31, 6) */,
  32'h3d15cc97 /* (26, 31, 6) */,
  32'h3d2567ce /* (22, 31, 6) */,
  32'h3d4cf093 /* (18, 31, 6) */,
  32'h3d4cf093 /* (14, 31, 6) */,
  32'h3d2567ce /* (10, 31, 6) */,
  32'h3d15cc97 /* (6, 31, 6) */,
  32'h3d3543e4 /* (2, 31, 6) */,
  32'h3d18df8d /* (30, 27, 6) */,
  32'h3d16bb8b /* (26, 27, 6) */,
  32'h3d3c300c /* (22, 27, 6) */,
  32'h3d786cd6 /* (18, 27, 6) */,
  32'h3d786cd6 /* (14, 27, 6) */,
  32'h3d3c300c /* (10, 27, 6) */,
  32'h3d16bb8b /* (6, 27, 6) */,
  32'h3d18df8d /* (2, 27, 6) */,
  32'h3d1e19af /* (30, 23, 6) */,
  32'h3d37f9d0 /* (26, 23, 6) */,
  32'h3d866682 /* (22, 23, 6) */,
  32'h3dc45939 /* (18, 23, 6) */,
  32'h3dc45939 /* (14, 23, 6) */,
  32'h3d866682 /* (10, 23, 6) */,
  32'h3d37f9d0 /* (6, 23, 6) */,
  32'h3d1e19af /* (2, 23, 6) */,
  32'h3d4ce87b /* (30, 19, 6) */,
  32'h3d82bc35 /* (26, 19, 6) */,
  32'h3dd610ea /* (22, 19, 6) */,
  32'h3e2b8c37 /* (18, 19, 6) */,
  32'h3e2b8c37 /* (14, 19, 6) */,
  32'h3dd610ea /* (10, 19, 6) */,
  32'h3d82bc35 /* (6, 19, 6) */,
  32'h3d4ce87b /* (2, 19, 6) */,
  32'h3d4bfe66 /* (30, 15, 6) */,
  32'h3d85e8bf /* (26, 15, 6) */,
  32'h3de44bb3 /* (22, 15, 6) */,
  32'h3e3e01e0 /* (18, 15, 6) */,
  32'h3e3e01e0 /* (14, 15, 6) */,
  32'h3de44bb3 /* (10, 15, 6) */,
  32'h3d85e8bf /* (6, 15, 6) */,
  32'h3d4bfe66 /* (2, 15, 6) */,
  32'h3d343ccb /* (30, 11, 6) */,
  32'h3d5d3b5c /* (26, 11, 6) */,
  32'h3dac23aa /* (22, 11, 6) */,
  32'h3e040b60 /* (18, 11, 6) */,
  32'h3e040b60 /* (14, 11, 6) */,
  32'h3dac23aa /* (10, 11, 6) */,
  32'h3d5d3b5c /* (6, 11, 6) */,
  32'h3d343ccb /* (2, 11, 6) */,
  32'h3d14b9d3 /* (30, 7, 6) */,
  32'h3d20f672 /* (26, 7, 6) */,
  32'h3d5a2934 /* (22, 7, 6) */,
  32'h3d975464 /* (18, 7, 6) */,
  32'h3d975464 /* (14, 7, 6) */,
  32'h3d5a2934 /* (10, 7, 6) */,
  32'h3d20f672 /* (6, 7, 6) */,
  32'h3d14b9d3 /* (2, 7, 6) */,
  32'h3d271e8d /* (30, 3, 6) */,
  32'h3d14c14d /* (26, 3, 6) */,
  32'h3d2c3293 /* (22, 3, 6) */,
  32'h3d5a5169 /* (18, 3, 6) */,
  32'h3d5a5169 /* (14, 3, 6) */,
  32'h3d2c3293 /* (10, 3, 6) */,
  32'h3d14c14d /* (6, 3, 6) */,
  32'h3d271e8d /* (2, 3, 6) */,
  32'h3e0c4d23 /* (30, 31, 2) */,
  32'h3d3543e4 /* (26, 31, 2) */,
  32'h3d12ac07 /* (22, 31, 2) */,
  32'h3d217487 /* (18, 31, 2) */,
  32'h3d217487 /* (14, 31, 2) */,
  32'h3d12ac07 /* (10, 31, 2) */,
  32'h3d3543e4 /* (6, 31, 2) */,
  32'h3e0c4d23 /* (2, 31, 2) */,
  32'h3d4ca49b /* (30, 27, 2) */,
  32'h3d18df8d /* (26, 27, 2) */,
  32'h3d1f9f49 /* (22, 27, 2) */,
  32'h3d40d8bf /* (18, 27, 2) */,
  32'h3d40d8bf /* (14, 27, 2) */,
  32'h3d1f9f49 /* (10, 27, 2) */,
  32'h3d18df8d /* (6, 27, 2) */,
  32'h3d4ca49b /* (2, 27, 2) */,
  32'h3d1214c5 /* (30, 23, 2) */,
  32'h3d1e19af /* (26, 23, 2) */,
  32'h3d56480e /* (22, 23, 2) */,
  32'h3d94a37c /* (18, 23, 2) */,
  32'h3d94a37c /* (14, 23, 2) */,
  32'h3d56480e /* (10, 23, 2) */,
  32'h3d1e19af /* (6, 23, 2) */,
  32'h3d1214c5 /* (2, 23, 2) */,
  32'h3d246fbd /* (30, 19, 2) */,
  32'h3d4ce87b /* (26, 19, 2) */,
  32'h3da2895a /* (22, 19, 2) */,
  32'h3dfd653f /* (18, 19, 2) */,
  32'h3dfd653f /* (14, 19, 2) */,
  32'h3da2895a /* (10, 19, 2) */,
  32'h3d4ce87b /* (6, 19, 2) */,
  32'h3d246fbd /* (2, 19, 2) */,
  32'h3d1dadb9 /* (30, 15, 2) */,
  32'h3d4bfe66 /* (26, 15, 2) */,
  32'h3daa3ec9 /* (22, 15, 2) */,
  32'h3e0adb0d /* (18, 15, 2) */,
  32'h3e0adb0d /* (14, 15, 2) */,
  32'h3daa3ec9 /* (10, 15, 2) */,
  32'h3d4bfe66 /* (6, 15, 2) */,
  32'h3d1dadb9 /* (2, 15, 2) */,
  32'h3d18e0f8 /* (30, 11, 2) */,
  32'h3d343ccb /* (26, 11, 2) */,
  32'h3d85a0b3 /* (22, 11, 2) */,
  32'h3dc55f41 /* (18, 11, 2) */,
  32'h3dc55f41 /* (14, 11, 2) */,
  32'h3d85a0b3 /* (10, 11, 2) */,
  32'h3d343ccb /* (6, 11, 2) */,
  32'h3d18e0f8 /* (2, 11, 2) */,
  32'h3d1dd271 /* (30, 7, 2) */,
  32'h3d14b9d3 /* (26, 7, 2) */,
  32'h3d3346c6 /* (22, 7, 2) */,
  32'h3d6820b1 /* (18, 7, 2) */,
  32'h3d6820b1 /* (14, 7, 2) */,
  32'h3d3346c6 /* (10, 7, 2) */,
  32'h3d14b9d3 /* (6, 7, 2) */,
  32'h3d1dd271 /* (2, 7, 2) */,
  32'h3da3af74 /* (30, 3, 2) */,
  32'h3d271e8d /* (26, 3, 2) */,
  32'h3d162b76 /* (22, 3, 2) */,
  32'h3d2b1735 /* (18, 3, 2) */,
  32'h3d2b1735 /* (14, 3, 2) */,
  32'h3d162b76 /* (10, 3, 2) */,
  32'h3d271e8d /* (6, 3, 2) */,
  32'h3da3af74 /* (2, 3, 2) */,
  32'h3dbfa8df /* (29, 31, 30) */,
  32'h3d20a35e /* (25, 31, 30) */,
  32'h3d16ed42 /* (21, 31, 30) */,
  32'h3d1a0745 /* (17, 31, 30) */,
  32'h3d214ba3 /* (13, 31, 30) */,
  32'h3d11c69f /* (9, 31, 30) */,
  32'h3d59109a /* (5, 31, 30) */,
  32'h3e4aeee2 /* (1, 31, 30) */,
  32'h3d3cd255 /* (29, 27, 30) */,
  32'h3d14b1c0 /* (25, 27, 30) */,
  32'h3d29823f /* (21, 27, 30) */,
  32'h3d3a7be5 /* (17, 27, 30) */,
  32'h3d3d84de /* (13, 27, 30) */,
  32'h3d18622e /* (9, 27, 30) */,
  32'h3d213c91 /* (5, 27, 30) */,
  32'h3d59109a /* (1, 27, 30) */,
  32'h3d12f42a /* (29, 23, 30) */,
  32'h3d26a1b5 /* (25, 23, 30) */,
  32'h3d6d9fa3 /* (21, 23, 30) */,
  32'h3d9314c2 /* (17, 23, 30) */,
  32'h3d8e358b /* (13, 23, 30) */,
  32'h3d42665b /* (9, 23, 30) */,
  32'h3d18622e /* (5, 23, 30) */,
  32'h3d11c69f /* (1, 23, 30) */,
  32'h3d29e985 /* (29, 19, 30) */,
  32'h3d6129ae /* (25, 19, 30) */,
  32'h3dba5db4 /* (21, 19, 30) */,
  32'h3e003b1e /* (17, 19, 30) */,
  32'h3dec70da /* (13, 19, 30) */,
  32'h3d8e358b /* (9, 19, 30) */,
  32'h3d3d84de /* (5, 19, 30) */,
  32'h3d214ba3 /* (1, 19, 30) */,
  32'h3d240321 /* (29, 15, 30) */,
  32'h3d62f778 /* (25, 15, 30) */,
  32'h3dc59b81 /* (21, 15, 30) */,
  32'h3e0de5f8 /* (17, 15, 30) */,
  32'h3e003b1e /* (13, 15, 30) */,
  32'h3d9314c2 /* (9, 15, 30) */,
  32'h3d3a7be5 /* (5, 15, 30) */,
  32'h3d1a0745 /* (1, 15, 30) */,
  32'h3d1c5f03 /* (29, 11, 30) */,
  32'h3d42a7b8 /* (25, 11, 30) */,
  32'h3d96eb50 /* (21, 11, 30) */,
  32'h3dc59b81 /* (17, 11, 30) */,
  32'h3dba5db4 /* (13, 11, 30) */,
  32'h3d6d9fa3 /* (9, 11, 30) */,
  32'h3d29823f /* (5, 11, 30) */,
  32'h3d16ed42 /* (1, 11, 30) */,
  32'h3d1a2949 /* (29, 7, 30) */,
  32'h3d1777c7 /* (25, 7, 30) */,
  32'h3d42a7b8 /* (21, 7, 30) */,
  32'h3d62f778 /* (17, 7, 30) */,
  32'h3d6129ae /* (13, 7, 30) */,
  32'h3d26a1b5 /* (9, 7, 30) */,
  32'h3d14b1c0 /* (5, 7, 30) */,
  32'h3d20a35e /* (1, 7, 30) */,
  32'h3d866355 /* (29, 3, 30) */,
  32'h3d1a2949 /* (25, 3, 30) */,
  32'h3d1c5f03 /* (21, 3, 30) */,
  32'h3d240321 /* (17, 3, 30) */,
  32'h3d29e985 /* (13, 3, 30) */,
  32'h3d12f42a /* (9, 3, 30) */,
  32'h3d3cd255 /* (5, 3, 30) */,
  32'h3dbfa8df /* (1, 3, 30) */,
  32'h3d2ba889 /* (29, 31, 26) */,
  32'h3d146a43 /* (25, 31, 26) */,
  32'h3d31191b /* (21, 31, 26) */,
  32'h3d46f53f /* (17, 31, 26) */,
  32'h3d4876ff /* (13, 31, 26) */,
  32'h3d1c53e8 /* (9, 31, 26) */,
  32'h3d1a8b5a /* (5, 31, 26) */,
  32'h3d3c9698 /* (1, 31, 26) */,
  32'h3d16d305 /* (29, 27, 26) */,
  32'h3d1b2471 /* (25, 27, 26) */,
  32'h3d4d9045 /* (21, 27, 26) */,
  32'h3d73b16f /* (17, 27, 26) */,
  32'h3d700ffa /* (13, 27, 26) */,
  32'h3d2db0cc /* (9, 27, 26) */,
  32'h3d14f7ce /* (5, 27, 26) */,
  32'h3d1a8b5a /* (1, 27, 26) */,
  32'h3d215063 /* (29, 23, 26) */,
  32'h3d45eb5b /* (25, 23, 26) */,
  32'h3d9750ce /* (21, 23, 26) */,
  32'h3dc42ad0 /* (17, 23, 26) */,
  32'h3db9d5f4 /* (13, 23, 26) */,
  32'h3d6fd024 /* (9, 23, 26) */,
  32'h3d2db0cc /* (5, 23, 26) */,
  32'h3d1c53e8 /* (1, 23, 26) */,
  32'h3d54a03b /* (29, 19, 26) */,
  32'h3d90c8a7 /* (25, 19, 26) */,
  32'h3df74dbc /* (21, 19, 26) */,
  32'h3e2ea39a /* (17, 19, 26) */,
  32'h3e1f113d /* (13, 19, 26) */,
  32'h3db9d5f4 /* (9, 19, 26) */,
  32'h3d700ffa /* (5, 19, 26) */,
  32'h3d4876ff /* (1, 19, 26) */,
  32'h3d54ba37 /* (29, 15, 26) */,
  32'h3d95be73 /* (25, 15, 26) */,
  32'h3e0533d0 /* (21, 15, 26) */,
  32'h3e430b11 /* (17, 15, 26) */,
  32'h3e2ea39a /* (13, 15, 26) */,
  32'h3dc42ad0 /* (9, 15, 26) */,
  32'h3d73b16f /* (5, 15, 26) */,
  32'h3d46f53f /* (1, 15, 26) */,
  32'h3d39bb76 /* (29, 11, 26) */,
  32'h3d71ecf9 /* (25, 11, 26) */,
  32'h3dc480ba /* (21, 11, 26) */,
  32'h3e0533d0 /* (17, 11, 26) */,
  32'h3df74dbc /* (13, 11, 26) */,
  32'h3d9750ce /* (9, 11, 26) */,
  32'h3d4d9045 /* (5, 11, 26) */,
  32'h3d31191b /* (1, 11, 26) */,
  32'h3d159d44 /* (29, 7, 26) */,
  32'h3d29a602 /* (25, 7, 26) */,
  32'h3d71ecf9 /* (21, 7, 26) */,
  32'h3d95be73 /* (17, 7, 26) */,
  32'h3d90c8a7 /* (13, 7, 26) */,
  32'h3d45eb5b /* (9, 7, 26) */,
  32'h3d1b2471 /* (5, 7, 26) */,
  32'h3d146a43 /* (1, 7, 26) */,
  32'h3d211f1b /* (29, 3, 26) */,
  32'h3d159d44 /* (25, 3, 26) */,
  32'h3d39bb76 /* (21, 3, 26) */,
  32'h3d54ba37 /* (17, 3, 26) */,
  32'h3d54a03b /* (13, 3, 26) */,
  32'h3d215063 /* (9, 3, 26) */,
  32'h3d16d305 /* (5, 3, 26) */,
  32'h3d2ba889 /* (1, 3, 26) */,
  32'h3d14c0fd /* (29, 31, 22) */,
  32'h3d305430 /* (25, 31, 22) */,
  32'h3d829849 /* (21, 31, 22) */,
  32'h3da5ac70 /* (17, 31, 22) */,
  32'h3d9e7894 /* (13, 31, 22) */,
  32'h3d52081f /* (9, 31, 22) */,
  32'h3d1d9589 /* (5, 31, 22) */,
  32'h3d119771 /* (1, 31, 22) */,
  32'h3d2344c4 /* (29, 27, 22) */,
  32'h3d4b3dc7 /* (25, 27, 22) */,
  32'h3d9d9380 /* (21, 27, 22) */,
  32'h3dce52e6 /* (17, 27, 22) */,
  32'h3dc29629 /* (13, 27, 22) */,
  32'h3d781ae6 /* (9, 27, 22) */,
  32'h3d30fc5a /* (5, 27, 22) */,
  32'h3d1d9589 /* (1, 27, 22) */,
  32'h3d5dae2c /* (29, 23, 22) */,
  32'h3d94014f /* (25, 23, 22) */,
  32'h3df71c69 /* (21, 23, 22) */,
  32'h3e2b3653 /* (17, 23, 22) */,
  32'h3e1d56b2 /* (13, 23, 22) */,
  32'h3dbbc730 /* (9, 23, 22) */,
  32'h3d781ae6 /* (5, 23, 22) */,
  32'h3d52081f /* (1, 23, 22) */,
  32'h3da99659 /* (29, 19, 22) */,
  32'h3defa49b /* (25, 19, 22) */,
  32'h3e562fb1 /* (21, 19, 22) */,
  32'h3e9d80fb /* (17, 19, 22) */,
  32'h3e8cbae1 /* (13, 19, 22) */,
  32'h3e1d56b2 /* (9, 19, 22) */,
  32'h3dc29629 /* (5, 19, 22) */,
  32'h3d9e7894 /* (1, 19, 22) */,
  32'h3db22d06 /* (29, 15, 22) */,
  32'h3e009a19 /* (25, 15, 22) */,
  32'h3e6c6ac0 /* (21, 15, 22) */,
  32'h3eb2925b /* (17, 15, 22) */,
  32'h3e9d80fb /* (13, 15, 22) */,
  32'h3e2b3653 /* (9, 15, 22) */,
  32'h3dce52e6 /* (5, 15, 22) */,
  32'h3da5ac70 /* (1, 15, 22) */,
  32'h3d8ae43c /* (29, 11, 22) */,
  32'h3dbf3f1d /* (25, 11, 22) */,
  32'h3e257fc6 /* (21, 11, 22) */,
  32'h3e6c6ac0 /* (17, 11, 22) */,
  32'h3e562fb1 /* (13, 11, 22) */,
  32'h3df71c69 /* (9, 11, 22) */,
  32'h3d9d9380 /* (5, 11, 22) */,
  32'h3d829849 /* (1, 11, 22) */,
  32'h3d387393 /* (29, 7, 22) */,
  32'h3d6deb12 /* (25, 7, 22) */,
  32'h3dbf3f1d /* (21, 7, 22) */,
  32'h3e009a19 /* (17, 7, 22) */,
  32'h3defa49b /* (13, 7, 22) */,
  32'h3d94014f /* (9, 7, 22) */,
  32'h3d4b3dc7 /* (5, 7, 22) */,
  32'h3d305430 /* (1, 7, 22) */,
  32'h3d18cb02 /* (29, 3, 22) */,
  32'h3d387393 /* (25, 3, 22) */,
  32'h3d8ae43c /* (21, 3, 22) */,
  32'h3db22d06 /* (17, 3, 22) */,
  32'h3da99659 /* (13, 3, 22) */,
  32'h3d5dae2c /* (9, 3, 22) */,
  32'h3d2344c4 /* (5, 3, 22) */,
  32'h3d14c0fd /* (1, 3, 22) */,
  32'h3d276174 /* (29, 31, 18) */,
  32'h3d62906c /* (25, 31, 18) */,
  32'h3dc01db4 /* (21, 31, 18) */,
  32'h3e06d8bb /* (17, 31, 18) */,
  32'h3df65860 /* (13, 31, 18) */,
  32'h3d90dff9 /* (9, 31, 18) */,
  32'h3d3c7841 /* (5, 31, 18) */,
  32'h3d1e0bb6 /* (1, 31, 18) */,
  32'h3d487174 /* (29, 27, 18) */,
  32'h3d8a0000 /* (25, 27, 18) */,
  32'h3deed79f /* (21, 27, 18) */,
  32'h3e2a981c /* (17, 27, 18) */,
  32'h3e1a8d8c /* (13, 27, 18) */,
  32'h3db24f8e /* (9, 27, 18) */,
  32'h3d63687e /* (5, 27, 18) */,
  32'h3d3c7841 /* (1, 27, 18) */,
  32'h3d9b2a7b /* (29, 23, 18) */,
  32'h3ddc09d8 /* (25, 23, 18) */,
  32'h3e458f30 /* (21, 23, 18) */,
  32'h3e91e4f8 /* (17, 23, 18) */,
  32'h3e821787 /* (13, 23, 18) */,
  32'h3e10cac5 /* (9, 23, 18) */,
  32'h3db24f8e /* (5, 23, 18) */,
  32'h3d90dff9 /* (1, 23, 18) */,
  32'h3e04d0b8 /* (29, 19, 18) */,
  32'h3e41f14c /* (25, 19, 18) */,
  32'h3eb517ce /* (21, 19, 18) */,
  32'h3f0af24f /* (17, 19, 18) */,
  32'h3ef33ce4 /* (13, 19, 18) */,
  32'h3e821787 /* (9, 19, 18) */,
  32'h3e1a8d8c /* (5, 19, 18) */,
  32'h3df65860 /* (1, 19, 18) */,
  32'h3e11d12f /* (29, 15, 18) */,
  32'h3e57a44b /* (25, 15, 18) */,
  32'h3eccf8ff /* (21, 15, 18) */,
  32'h3f202f9a /* (17, 15, 18) */,
  32'h3f0af24f /* (13, 15, 18) */,
  32'h3e91e4f8 /* (9, 15, 18) */,
  32'h3e2a981c /* (5, 15, 18) */,
  32'h3e06d8bb /* (1, 15, 18) */,
  32'h3dce7d45 /* (29, 11, 18) */,
  32'h3e14a5c9 /* (25, 11, 18) */,
  32'h3e882756 /* (21, 11, 18) */,
  32'h3eccf8ff /* (17, 11, 18) */,
  32'h3eb517ce /* (13, 11, 18) */,
  32'h3e458f30 /* (9, 11, 18) */,
  32'h3deed79f /* (5, 11, 18) */,
  32'h3dc01db4 /* (1, 11, 18) */,
  32'h3d71c736 /* (29, 7, 18) */,
  32'h3da8d240 /* (25, 7, 18) */,
  32'h3e14a5c9 /* (21, 7, 18) */,
  32'h3e57a44b /* (17, 7, 18) */,
  32'h3e41f14c /* (13, 7, 18) */,
  32'h3ddc09d8 /* (9, 7, 18) */,
  32'h3d8a0000 /* (5, 7, 18) */,
  32'h3d62906c /* (1, 7, 18) */,
  32'h3d3188e3 /* (29, 3, 18) */,
  32'h3d71c736 /* (25, 3, 18) */,
  32'h3dce7d45 /* (21, 3, 18) */,
  32'h3e11d12f /* (17, 3, 18) */,
  32'h3e04d0b8 /* (13, 3, 18) */,
  32'h3d9b2a7b /* (9, 3, 18) */,
  32'h3d487174 /* (5, 3, 18) */,
  32'h3d276174 /* (1, 3, 18) */,
  32'h3d276174 /* (29, 31, 14) */,
  32'h3d62906c /* (25, 31, 14) */,
  32'h3dc01db4 /* (21, 31, 14) */,
  32'h3e06d8bb /* (17, 31, 14) */,
  32'h3df65860 /* (13, 31, 14) */,
  32'h3d90dff9 /* (9, 31, 14) */,
  32'h3d3c7841 /* (5, 31, 14) */,
  32'h3d1e0bb6 /* (1, 31, 14) */,
  32'h3d487174 /* (29, 27, 14) */,
  32'h3d8a0000 /* (25, 27, 14) */,
  32'h3deed79f /* (21, 27, 14) */,
  32'h3e2a981c /* (17, 27, 14) */,
  32'h3e1a8d8c /* (13, 27, 14) */,
  32'h3db24f8e /* (9, 27, 14) */,
  32'h3d63687e /* (5, 27, 14) */,
  32'h3d3c7841 /* (1, 27, 14) */,
  32'h3d9b2a7b /* (29, 23, 14) */,
  32'h3ddc09d8 /* (25, 23, 14) */,
  32'h3e458f30 /* (21, 23, 14) */,
  32'h3e91e4f8 /* (17, 23, 14) */,
  32'h3e821787 /* (13, 23, 14) */,
  32'h3e10cac5 /* (9, 23, 14) */,
  32'h3db24f8e /* (5, 23, 14) */,
  32'h3d90dff9 /* (1, 23, 14) */,
  32'h3e04d0b8 /* (29, 19, 14) */,
  32'h3e41f14c /* (25, 19, 14) */,
  32'h3eb517ce /* (21, 19, 14) */,
  32'h3f0af24f /* (17, 19, 14) */,
  32'h3ef33ce4 /* (13, 19, 14) */,
  32'h3e821787 /* (9, 19, 14) */,
  32'h3e1a8d8c /* (5, 19, 14) */,
  32'h3df65860 /* (1, 19, 14) */,
  32'h3e11d12f /* (29, 15, 14) */,
  32'h3e57a44b /* (25, 15, 14) */,
  32'h3eccf8ff /* (21, 15, 14) */,
  32'h3f202f9a /* (17, 15, 14) */,
  32'h3f0af24f /* (13, 15, 14) */,
  32'h3e91e4f8 /* (9, 15, 14) */,
  32'h3e2a981c /* (5, 15, 14) */,
  32'h3e06d8bb /* (1, 15, 14) */,
  32'h3dce7d45 /* (29, 11, 14) */,
  32'h3e14a5c9 /* (25, 11, 14) */,
  32'h3e882756 /* (21, 11, 14) */,
  32'h3eccf8ff /* (17, 11, 14) */,
  32'h3eb517ce /* (13, 11, 14) */,
  32'h3e458f30 /* (9, 11, 14) */,
  32'h3deed79f /* (5, 11, 14) */,
  32'h3dc01db4 /* (1, 11, 14) */,
  32'h3d71c736 /* (29, 7, 14) */,
  32'h3da8d240 /* (25, 7, 14) */,
  32'h3e14a5c9 /* (21, 7, 14) */,
  32'h3e57a44b /* (17, 7, 14) */,
  32'h3e41f14c /* (13, 7, 14) */,
  32'h3ddc09d8 /* (9, 7, 14) */,
  32'h3d8a0000 /* (5, 7, 14) */,
  32'h3d62906c /* (1, 7, 14) */,
  32'h3d3188e3 /* (29, 3, 14) */,
  32'h3d71c736 /* (25, 3, 14) */,
  32'h3dce7d45 /* (21, 3, 14) */,
  32'h3e11d12f /* (17, 3, 14) */,
  32'h3e04d0b8 /* (13, 3, 14) */,
  32'h3d9b2a7b /* (9, 3, 14) */,
  32'h3d487174 /* (5, 3, 14) */,
  32'h3d276174 /* (1, 3, 14) */,
  32'h3d14c0fd /* (29, 31, 10) */,
  32'h3d305430 /* (25, 31, 10) */,
  32'h3d829849 /* (21, 31, 10) */,
  32'h3da5ac70 /* (17, 31, 10) */,
  32'h3d9e7894 /* (13, 31, 10) */,
  32'h3d52081f /* (9, 31, 10) */,
  32'h3d1d9589 /* (5, 31, 10) */,
  32'h3d119771 /* (1, 31, 10) */,
  32'h3d2344c4 /* (29, 27, 10) */,
  32'h3d4b3dc7 /* (25, 27, 10) */,
  32'h3d9d9380 /* (21, 27, 10) */,
  32'h3dce52e6 /* (17, 27, 10) */,
  32'h3dc29629 /* (13, 27, 10) */,
  32'h3d781ae6 /* (9, 27, 10) */,
  32'h3d30fc5a /* (5, 27, 10) */,
  32'h3d1d9589 /* (1, 27, 10) */,
  32'h3d5dae2c /* (29, 23, 10) */,
  32'h3d94014f /* (25, 23, 10) */,
  32'h3df71c69 /* (21, 23, 10) */,
  32'h3e2b3653 /* (17, 23, 10) */,
  32'h3e1d56b2 /* (13, 23, 10) */,
  32'h3dbbc730 /* (9, 23, 10) */,
  32'h3d781ae6 /* (5, 23, 10) */,
  32'h3d52081f /* (1, 23, 10) */,
  32'h3da99659 /* (29, 19, 10) */,
  32'h3defa49b /* (25, 19, 10) */,
  32'h3e562fb1 /* (21, 19, 10) */,
  32'h3e9d80fb /* (17, 19, 10) */,
  32'h3e8cbae1 /* (13, 19, 10) */,
  32'h3e1d56b2 /* (9, 19, 10) */,
  32'h3dc29629 /* (5, 19, 10) */,
  32'h3d9e7894 /* (1, 19, 10) */,
  32'h3db22d06 /* (29, 15, 10) */,
  32'h3e009a19 /* (25, 15, 10) */,
  32'h3e6c6ac0 /* (21, 15, 10) */,
  32'h3eb2925b /* (17, 15, 10) */,
  32'h3e9d80fb /* (13, 15, 10) */,
  32'h3e2b3653 /* (9, 15, 10) */,
  32'h3dce52e6 /* (5, 15, 10) */,
  32'h3da5ac70 /* (1, 15, 10) */,
  32'h3d8ae43c /* (29, 11, 10) */,
  32'h3dbf3f1d /* (25, 11, 10) */,
  32'h3e257fc6 /* (21, 11, 10) */,
  32'h3e6c6ac0 /* (17, 11, 10) */,
  32'h3e562fb1 /* (13, 11, 10) */,
  32'h3df71c69 /* (9, 11, 10) */,
  32'h3d9d9380 /* (5, 11, 10) */,
  32'h3d829849 /* (1, 11, 10) */,
  32'h3d387393 /* (29, 7, 10) */,
  32'h3d6deb12 /* (25, 7, 10) */,
  32'h3dbf3f1d /* (21, 7, 10) */,
  32'h3e009a19 /* (17, 7, 10) */,
  32'h3defa49b /* (13, 7, 10) */,
  32'h3d94014f /* (9, 7, 10) */,
  32'h3d4b3dc7 /* (5, 7, 10) */,
  32'h3d305430 /* (1, 7, 10) */,
  32'h3d18cb02 /* (29, 3, 10) */,
  32'h3d387393 /* (25, 3, 10) */,
  32'h3d8ae43c /* (21, 3, 10) */,
  32'h3db22d06 /* (17, 3, 10) */,
  32'h3da99659 /* (13, 3, 10) */,
  32'h3d5dae2c /* (9, 3, 10) */,
  32'h3d2344c4 /* (5, 3, 10) */,
  32'h3d14c0fd /* (1, 3, 10) */,
  32'h3d2ba889 /* (29, 31, 6) */,
  32'h3d146a43 /* (25, 31, 6) */,
  32'h3d31191b /* (21, 31, 6) */,
  32'h3d46f53f /* (17, 31, 6) */,
  32'h3d4876ff /* (13, 31, 6) */,
  32'h3d1c53e8 /* (9, 31, 6) */,
  32'h3d1a8b5a /* (5, 31, 6) */,
  32'h3d3c9698 /* (1, 31, 6) */,
  32'h3d16d305 /* (29, 27, 6) */,
  32'h3d1b2471 /* (25, 27, 6) */,
  32'h3d4d9045 /* (21, 27, 6) */,
  32'h3d73b16f /* (17, 27, 6) */,
  32'h3d700ffa /* (13, 27, 6) */,
  32'h3d2db0cc /* (9, 27, 6) */,
  32'h3d14f7ce /* (5, 27, 6) */,
  32'h3d1a8b5a /* (1, 27, 6) */,
  32'h3d215063 /* (29, 23, 6) */,
  32'h3d45eb5b /* (25, 23, 6) */,
  32'h3d9750ce /* (21, 23, 6) */,
  32'h3dc42ad0 /* (17, 23, 6) */,
  32'h3db9d5f4 /* (13, 23, 6) */,
  32'h3d6fd024 /* (9, 23, 6) */,
  32'h3d2db0cc /* (5, 23, 6) */,
  32'h3d1c53e8 /* (1, 23, 6) */,
  32'h3d54a03b /* (29, 19, 6) */,
  32'h3d90c8a7 /* (25, 19, 6) */,
  32'h3df74dbc /* (21, 19, 6) */,
  32'h3e2ea39a /* (17, 19, 6) */,
  32'h3e1f113d /* (13, 19, 6) */,
  32'h3db9d5f4 /* (9, 19, 6) */,
  32'h3d700ffa /* (5, 19, 6) */,
  32'h3d4876ff /* (1, 19, 6) */,
  32'h3d54ba37 /* (29, 15, 6) */,
  32'h3d95be73 /* (25, 15, 6) */,
  32'h3e0533d0 /* (21, 15, 6) */,
  32'h3e430b11 /* (17, 15, 6) */,
  32'h3e2ea39a /* (13, 15, 6) */,
  32'h3dc42ad0 /* (9, 15, 6) */,
  32'h3d73b16f /* (5, 15, 6) */,
  32'h3d46f53f /* (1, 15, 6) */,
  32'h3d39bb76 /* (29, 11, 6) */,
  32'h3d71ecf9 /* (25, 11, 6) */,
  32'h3dc480ba /* (21, 11, 6) */,
  32'h3e0533d0 /* (17, 11, 6) */,
  32'h3df74dbc /* (13, 11, 6) */,
  32'h3d9750ce /* (9, 11, 6) */,
  32'h3d4d9045 /* (5, 11, 6) */,
  32'h3d31191b /* (1, 11, 6) */,
  32'h3d159d44 /* (29, 7, 6) */,
  32'h3d29a602 /* (25, 7, 6) */,
  32'h3d71ecf9 /* (21, 7, 6) */,
  32'h3d95be73 /* (17, 7, 6) */,
  32'h3d90c8a7 /* (13, 7, 6) */,
  32'h3d45eb5b /* (9, 7, 6) */,
  32'h3d1b2471 /* (5, 7, 6) */,
  32'h3d146a43 /* (1, 7, 6) */,
  32'h3d211f1b /* (29, 3, 6) */,
  32'h3d159d44 /* (25, 3, 6) */,
  32'h3d39bb76 /* (21, 3, 6) */,
  32'h3d54ba37 /* (17, 3, 6) */,
  32'h3d54a03b /* (13, 3, 6) */,
  32'h3d215063 /* (9, 3, 6) */,
  32'h3d16d305 /* (5, 3, 6) */,
  32'h3d2ba889 /* (1, 3, 6) */,
  32'h3dbfa8df /* (29, 31, 2) */,
  32'h3d20a35e /* (25, 31, 2) */,
  32'h3d16ed42 /* (21, 31, 2) */,
  32'h3d1a0745 /* (17, 31, 2) */,
  32'h3d214ba3 /* (13, 31, 2) */,
  32'h3d11c69f /* (9, 31, 2) */,
  32'h3d59109a /* (5, 31, 2) */,
  32'h3e4aeee2 /* (1, 31, 2) */,
  32'h3d3cd255 /* (29, 27, 2) */,
  32'h3d14b1c0 /* (25, 27, 2) */,
  32'h3d29823f /* (21, 27, 2) */,
  32'h3d3a7be5 /* (17, 27, 2) */,
  32'h3d3d84de /* (13, 27, 2) */,
  32'h3d18622e /* (9, 27, 2) */,
  32'h3d213c91 /* (5, 27, 2) */,
  32'h3d59109a /* (1, 27, 2) */,
  32'h3d12f42a /* (29, 23, 2) */,
  32'h3d26a1b5 /* (25, 23, 2) */,
  32'h3d6d9fa3 /* (21, 23, 2) */,
  32'h3d9314c2 /* (17, 23, 2) */,
  32'h3d8e358b /* (13, 23, 2) */,
  32'h3d42665b /* (9, 23, 2) */,
  32'h3d18622e /* (5, 23, 2) */,
  32'h3d11c69f /* (1, 23, 2) */,
  32'h3d29e985 /* (29, 19, 2) */,
  32'h3d6129ae /* (25, 19, 2) */,
  32'h3dba5db4 /* (21, 19, 2) */,
  32'h3e003b1e /* (17, 19, 2) */,
  32'h3dec70da /* (13, 19, 2) */,
  32'h3d8e358b /* (9, 19, 2) */,
  32'h3d3d84de /* (5, 19, 2) */,
  32'h3d214ba3 /* (1, 19, 2) */,
  32'h3d240321 /* (29, 15, 2) */,
  32'h3d62f778 /* (25, 15, 2) */,
  32'h3dc59b81 /* (21, 15, 2) */,
  32'h3e0de5f8 /* (17, 15, 2) */,
  32'h3e003b1e /* (13, 15, 2) */,
  32'h3d9314c2 /* (9, 15, 2) */,
  32'h3d3a7be5 /* (5, 15, 2) */,
  32'h3d1a0745 /* (1, 15, 2) */,
  32'h3d1c5f03 /* (29, 11, 2) */,
  32'h3d42a7b8 /* (25, 11, 2) */,
  32'h3d96eb50 /* (21, 11, 2) */,
  32'h3dc59b81 /* (17, 11, 2) */,
  32'h3dba5db4 /* (13, 11, 2) */,
  32'h3d6d9fa3 /* (9, 11, 2) */,
  32'h3d29823f /* (5, 11, 2) */,
  32'h3d16ed42 /* (1, 11, 2) */,
  32'h3d1a2949 /* (29, 7, 2) */,
  32'h3d1777c7 /* (25, 7, 2) */,
  32'h3d42a7b8 /* (21, 7, 2) */,
  32'h3d62f778 /* (17, 7, 2) */,
  32'h3d6129ae /* (13, 7, 2) */,
  32'h3d26a1b5 /* (9, 7, 2) */,
  32'h3d14b1c0 /* (5, 7, 2) */,
  32'h3d20a35e /* (1, 7, 2) */,
  32'h3d866355 /* (29, 3, 2) */,
  32'h3d1a2949 /* (25, 3, 2) */,
  32'h3d1c5f03 /* (21, 3, 2) */,
  32'h3d240321 /* (17, 3, 2) */,
  32'h3d29e985 /* (13, 3, 2) */,
  32'h3d12f42a /* (9, 3, 2) */,
  32'h3d3cd255 /* (5, 3, 2) */,
  32'h3dbfa8df /* (1, 3, 2) */,
  32'h3d8b1391 /* (28, 31, 30) */,
  32'h3d15ce12 /* (24, 31, 30) */,
  32'h3d1cac31 /* (20, 31, 30) */,
  32'h3d09dfab /* (16, 31, 30) */,
  32'h3d1cac31 /* (12, 31, 30) */,
  32'h3d15ce12 /* (8, 31, 30) */,
  32'h3d8b1391 /* (4, 31, 30) */,
  32'h3e709592 /* (0, 31, 30) */,
  32'h3d2d8e0e /* (28, 27, 30) */,
  32'h3d149b5c /* (24, 27, 30) */,
  32'h3d346b02 /* (20, 27, 30) */,
  32'h3d28d1e5 /* (16, 27, 30) */,
  32'h3d346b02 /* (12, 27, 30) */,
  32'h3d149b5c /* (8, 27, 30) */,
  32'h3d2d8e0e /* (4, 27, 30) */,
  32'h3d5dd7d1 /* (0, 27, 30) */,
  32'h3d14de35 /* (28, 23, 30) */,
  32'h3d3291f6 /* (24, 23, 30) */,
  32'h3d833332 /* (20, 23, 30) */,
  32'h3d87d16b /* (16, 23, 30) */,
  32'h3d833332 /* (12, 23, 30) */,
  32'h3d3291f6 /* (8, 23, 30) */,
  32'h3d14de35 /* (4, 23, 30) */,
  32'h3d11b684 /* (0, 23, 30) */,
  32'h3d3217f4 /* (28, 19, 30) */,
  32'h3d7b52f8 /* (24, 19, 30) */,
  32'h3dd42d31 /* (20, 19, 30) */,
  32'h3df1ae3d /* (16, 19, 30) */,
  32'h3dd42d31 /* (12, 19, 30) */,
  32'h3d7b52f8 /* (8, 19, 30) */,
  32'h3d3217f4 /* (4, 19, 30) */,
  32'h3d2045b1 /* (0, 19, 30) */,
  32'h3d2d6bba /* (28, 15, 30) */,
  32'h3d804df8 /* (24, 15, 30) */,
  32'h3de39dff /* (20, 15, 30) */,
  32'h3e06ec2e /* (16, 15, 30) */,
  32'h3de39dff /* (12, 15, 30) */,
  32'h3d804df8 /* (8, 15, 30) */,
  32'h3d2d6bba /* (4, 15, 30) */,
  32'h3d18d610 /* (0, 15, 30) */,
  32'h3d21c128 /* (28, 11, 30) */,
  32'h3d558b1c /* (24, 11, 30) */,
  32'h3da96c08 /* (20, 11, 30) */,
  32'h3db86416 /* (16, 11, 30) */,
  32'h3da96c08 /* (12, 11, 30) */,
  32'h3d558b1c /* (8, 11, 30) */,
  32'h3d21c128 /* (4, 11, 30) */,
  32'h3d164ce1 /* (0, 11, 30) */,
  32'h3d16c6a3 /* (28, 7, 30) */,
  32'h3d1d59b0 /* (24, 7, 30) */,
  32'h3d530d8e /* (20, 7, 30) */,
  32'h3d4f6a6e /* (16, 7, 30) */,
  32'h3d530d8e /* (12, 7, 30) */,
  32'h3d1d59b0 /* (8, 7, 30) */,
  32'h3d16c6a3 /* (4, 7, 30) */,
  32'h3d21b235 /* (0, 7, 30) */,
  32'h3d5defd3 /* (28, 3, 30) */,
  32'h3d13e9f7 /* (24, 3, 30) */,
  32'h3d23d587 /* (20, 3, 30) */,
  32'h3d13661d /* (16, 3, 30) */,
  32'h3d23d587 /* (12, 3, 30) */,
  32'h3d13e9f7 /* (8, 3, 30) */,
  32'h3d5defd3 /* (4, 3, 30) */,
  32'h3dcbea25 /* (0, 3, 30) */,
  32'h3d222a9c /* (28, 31, 26) */,
  32'h3d169650 /* (24, 31, 26) */,
  32'h3d3dc5f0 /* (20, 31, 26) */,
  32'h3d34b66a /* (16, 31, 26) */,
  32'h3d3dc5f0 /* (12, 31, 26) */,
  32'h3d169650 /* (8, 31, 26) */,
  32'h3d222a9c /* (4, 31, 26) */,
  32'h3d3f59b8 /* (0, 31, 26) */,
  32'h3d153e19 /* (28, 27, 26) */,
  32'h3d22af34 /* (24, 27, 26) */,
  32'h3d6007ad /* (20, 27, 26) */,
  32'h3d5f53fb /* (16, 27, 26) */,
  32'h3d6007ad /* (12, 27, 26) */,
  32'h3d22af34 /* (8, 27, 26) */,
  32'h3d153e19 /* (4, 27, 26) */,
  32'h3d1b2f33 /* (0, 27, 26) */,
  32'h3d2657dd /* (28, 23, 26) */,
  32'h3d584c0c /* (24, 23, 26) */,
  32'h3da96159 /* (20, 23, 26) */,
  32'h3db6b309 /* (16, 23, 26) */,
  32'h3da96159 /* (12, 23, 26) */,
  32'h3d584c0c /* (8, 23, 26) */,
  32'h3d2657dd /* (4, 23, 26) */,
  32'h3d1bc36a /* (0, 23, 26) */,
  32'h3d601ae9 /* (28, 19, 26) */,
  32'h3da2e7a9 /* (24, 19, 26) */,
  32'h3e0dc95f /* (20, 19, 26) */,
  32'h3e2576a9 /* (16, 19, 26) */,
  32'h3e0dc95f /* (12, 19, 26) */,
  32'h3da2e7a9 /* (8, 19, 26) */,
  32'h3d601ae9 /* (4, 19, 26) */,
  32'h3d4703b2 /* (0, 19, 26) */,
  32'h3d61b1de /* (28, 15, 26) */,
  32'h3daa3349 /* (24, 15, 26) */,
  32'h3e1a3a56 /* (20, 15, 26) */,
  32'h3e3a3d1a /* (16, 15, 26) */,
  32'h3e1a3a56 /* (12, 15, 26) */,
  32'h3daa3349 /* (8, 15, 26) */,
  32'h3d61b1de /* (4, 15, 26) */,
  32'h3d455011 /* (0, 15, 26) */,
  32'h3d41fb9f /* (28, 11, 26) */,
  32'h3d865b59 /* (24, 11, 26) */,
  32'h3ddec971 /* (20, 11, 26) */,
  32'h3dfa4afe /* (16, 11, 26) */,
  32'h3ddec971 /* (12, 11, 26) */,
  32'h3d865b59 /* (8, 11, 26) */,
  32'h3d41fb9f /* (4, 11, 26) */,
  32'h3d3013e2 /* (0, 11, 26) */,
  32'h3d17902e /* (28, 7, 26) */,
  32'h3d35cd98 /* (24, 7, 26) */,
  32'h3d859348 /* (20, 7, 26) */,
  32'h3d8a46e7 /* (16, 7, 26) */,
  32'h3d859348 /* (12, 7, 26) */,
  32'h3d35cd98 /* (8, 7, 26) */,
  32'h3d17902e /* (4, 7, 26) */,
  32'h3d1459dd /* (0, 7, 26) */,
  32'h3d1b3fff /* (28, 3, 26) */,
  32'h3d19bf4b /* (24, 3, 26) */,
  32'h3d48406d /* (20, 3, 26) */,
  32'h3d41d3ae /* (16, 3, 26) */,
  32'h3d48406d /* (12, 3, 26) */,
  32'h3d19bf4b /* (8, 3, 26) */,
  32'h3d1b3fff /* (4, 3, 26) */,
  32'h3d2d5b95 /* (0, 3, 26) */,
  32'h3d1839e3 /* (28, 31, 22) */,
  32'h3d3f0366 /* (24, 31, 22) */,
  32'h3d91435f /* (20, 31, 22) */,
  32'h3d99ac24 /* (16, 31, 22) */,
  32'h3d91435f /* (12, 31, 22) */,
  32'h3d3f0366 /* (8, 31, 22) */,
  32'h3d1839e3 /* (4, 31, 22) */,
  32'h3d1142bb /* (0, 31, 22) */,
  32'h3d28e3b2 /* (28, 27, 22) */,
  32'h3d5ef675 /* (24, 27, 22) */,
  32'h3db0e528 /* (20, 27, 22) */,
  32'h3dc0863e /* (16, 27, 22) */,
  32'h3db0e528 /* (12, 27, 22) */,
  32'h3d5ef675 /* (8, 27, 22) */,
  32'h3d28e3b2 /* (4, 27, 22) */,
  32'h3d1cee15 /* (0, 27, 22) */,
  32'h3d68b7a2 /* (28, 23, 22) */,
  32'h3da590e9 /* (24, 23, 22) */,
  32'h3e0cf021 /* (20, 23, 22) */,
  32'h3e21930d /* (16, 23, 22) */,
  32'h3e0cf021 /* (12, 23, 22) */,
  32'h3da590e9 /* (8, 23, 22) */,
  32'h3d68b7a2 /* (4, 23, 22) */,
  32'h3d50a575 /* (0, 23, 22) */,
  32'h3db40e50 /* (28, 19, 22) */,
  32'h3e085939 /* (24, 19, 22) */,
  32'h3e7848b5 /* (20, 19, 22) */,
  32'h3e968a40 /* (16, 19, 22) */,
  32'h3e7848b5 /* (12, 19, 22) */,
  32'h3e085939 /* (8, 19, 22) */,
  32'h3db40e50 /* (4, 19, 22) */,
  32'h3d9d248b /* (0, 19, 22) */,
  32'h3dbdf4f8 /* (28, 15, 22) */,
  32'h3e135573 /* (24, 15, 22) */,
  32'h3e89fde5 /* (20, 15, 22) */,
  32'h3eabb572 /* (16, 15, 22) */,
  32'h3e89fde5 /* (12, 15, 22) */,
  32'h3e135573 /* (8, 15, 22) */,
  32'h3dbdf4f8 /* (4, 15, 22) */,
  32'h3da42e1b /* (0, 15, 22) */,
  32'h3d92b699 /* (28, 11, 22) */,
  32'h3dd7e578 /* (24, 11, 22) */,
  32'h3e3e5baf /* (20, 11, 22) */,
  32'h3e60898b /* (16, 11, 22) */,
  32'h3e3e5baf /* (12, 11, 22) */,
  32'h3dd7e578 /* (8, 11, 22) */,
  32'h3d92b699 /* (4, 11, 22) */,
  32'h3d819abc /* (0, 11, 22) */,
  32'h3d404057 /* (28, 7, 22) */,
  32'h3d83c517 /* (24, 7, 22) */,
  32'h3dd85675 /* (20, 7, 22) */,
  32'h3df142da /* (16, 7, 22) */,
  32'h3dd85675 /* (12, 7, 22) */,
  32'h3d83c517 /* (8, 7, 22) */,
  32'h3d404057 /* (4, 7, 22) */,
  32'h3d2f5f5a /* (0, 7, 22) */,
  32'h3d1cff11 /* (28, 3, 22) */,
  32'h3d48bc7e /* (24, 3, 22) */,
  32'h3d9aff71 /* (20, 3, 22) */,
  32'h3da59d10 /* (16, 3, 22) */,
  32'h3d9aff71 /* (12, 3, 22) */,
  32'h3d48bc7e /* (8, 3, 22) */,
  32'h3d1cff11 /* (4, 3, 22) */,
  32'h3d144f19 /* (0, 3, 22) */,
  32'h3d303352 /* (28, 31, 18) */,
  32'h3d7e759f /* (24, 31, 18) */,
  32'h3ddbed5a /* (20, 31, 18) */,
  32'h3dff32bb /* (16, 31, 18) */,
  32'h3ddbed5a /* (12, 31, 18) */,
  32'h3d7e759f /* (8, 31, 18) */,
  32'h3d303352 /* (4, 31, 18) */,
  32'h3d1ceee6 /* (0, 31, 18) */,
  32'h3d53bb31 /* (28, 27, 18) */,
  32'h3d9bc970 /* (24, 27, 18) */,
  32'h3e095be4 /* (20, 27, 18) */,
  32'h3e2205a1 /* (16, 27, 18) */,
  32'h3e095be4 /* (12, 27, 18) */,
  32'h3d9bc970 /* (8, 27, 18) */,
  32'h3d53bb31 /* (4, 27, 18) */,
  32'h3d3b0a55 /* (0, 27, 18) */,
  32'h3da4db8a /* (28, 23, 18) */,
  32'h3dfaaa60 /* (24, 23, 18) */,
  32'h3e654448 /* (20, 23, 18) */,
  32'h3e8b9344 /* (16, 23, 18) */,
  32'h3e654448 /* (12, 23, 18) */,
  32'h3dfaaa60 /* (8, 23, 18) */,
  32'h3da4db8a /* (4, 23, 18) */,
  32'h3d8fa52c /* (0, 23, 18) */,
  32'h3e0de89e /* (28, 19, 18) */,
  32'h3e5f05ce /* (24, 19, 18) */,
  32'h3ed441df /* (20, 19, 18) */,
  32'h3f06176f /* (16, 19, 18) */,
  32'h3ed441df /* (12, 19, 18) */,
  32'h3e5f05ce /* (8, 19, 18) */,
  32'h3e0de89e /* (4, 19, 18) */,
  32'h3df40add /* (0, 19, 18) */,
  32'h3e1c2ca1 /* (28, 15, 18) */,
  32'h3e79034c /* (24, 15, 18) */,
  32'h3ef15f91 /* (20, 15, 18) */,
  32'h3f1b42bd /* (16, 15, 18) */,
  32'h3ef15f91 /* (12, 15, 18) */,
  32'h3e79034c /* (8, 15, 18) */,
  32'h3e1c2ca1 /* (4, 15, 18) */,
  32'h3e05899d /* (0, 15, 18) */,
  32'h3ddc0819 /* (28, 11, 18) */,
  32'h3e2a27e4 /* (24, 11, 18) */,
  32'h3e9ecc49 /* (20, 11, 18) */,
  32'h3ec4f0a1 /* (16, 11, 18) */,
  32'h3e9ecc49 /* (12, 11, 18) */,
  32'h3e2a27e4 /* (8, 11, 18) */,
  32'h3ddc0819 /* (4, 11, 18) */,
  32'h3dbe661f /* (0, 11, 18) */,
  32'h3d800deb /* (28, 7, 18) */,
  32'h3dbf672f /* (24, 7, 18) */,
  32'h3e2baf50 /* (20, 7, 18) */,
  32'h3e4d7ce8 /* (16, 7, 18) */,
  32'h3e2baf50 /* (12, 7, 18) */,
  32'h3dbf672f /* (8, 7, 18) */,
  32'h3d800deb /* (4, 7, 18) */,
  32'h3d60bf24 /* (0, 7, 18) */,
  32'h3d3b1e93 /* (28, 3, 18) */,
  32'h3d880501 /* (24, 3, 18) */,
  32'h3decc5e8 /* (20, 3, 18) */,
  32'h3e0a27e7 /* (16, 3, 18) */,
  32'h3decc5e8 /* (12, 3, 18) */,
  32'h3d880501 /* (8, 3, 18) */,
  32'h3d3b1e93 /* (4, 3, 18) */,
  32'h3d262b6e /* (0, 3, 18) */,
  32'h3d303352 /* (28, 31, 14) */,
  32'h3d7e759f /* (24, 31, 14) */,
  32'h3ddbed5a /* (20, 31, 14) */,
  32'h3dff32bb /* (16, 31, 14) */,
  32'h3ddbed5a /* (12, 31, 14) */,
  32'h3d7e759f /* (8, 31, 14) */,
  32'h3d303352 /* (4, 31, 14) */,
  32'h3d1ceee6 /* (0, 31, 14) */,
  32'h3d53bb31 /* (28, 27, 14) */,
  32'h3d9bc970 /* (24, 27, 14) */,
  32'h3e095be4 /* (20, 27, 14) */,
  32'h3e2205a1 /* (16, 27, 14) */,
  32'h3e095be4 /* (12, 27, 14) */,
  32'h3d9bc970 /* (8, 27, 14) */,
  32'h3d53bb31 /* (4, 27, 14) */,
  32'h3d3b0a55 /* (0, 27, 14) */,
  32'h3da4db8a /* (28, 23, 14) */,
  32'h3dfaaa60 /* (24, 23, 14) */,
  32'h3e654448 /* (20, 23, 14) */,
  32'h3e8b9344 /* (16, 23, 14) */,
  32'h3e654448 /* (12, 23, 14) */,
  32'h3dfaaa60 /* (8, 23, 14) */,
  32'h3da4db8a /* (4, 23, 14) */,
  32'h3d8fa52c /* (0, 23, 14) */,
  32'h3e0de89e /* (28, 19, 14) */,
  32'h3e5f05ce /* (24, 19, 14) */,
  32'h3ed441df /* (20, 19, 14) */,
  32'h3f06176f /* (16, 19, 14) */,
  32'h3ed441df /* (12, 19, 14) */,
  32'h3e5f05ce /* (8, 19, 14) */,
  32'h3e0de89e /* (4, 19, 14) */,
  32'h3df40add /* (0, 19, 14) */,
  32'h3e1c2ca1 /* (28, 15, 14) */,
  32'h3e79034c /* (24, 15, 14) */,
  32'h3ef15f91 /* (20, 15, 14) */,
  32'h3f1b42bd /* (16, 15, 14) */,
  32'h3ef15f91 /* (12, 15, 14) */,
  32'h3e79034c /* (8, 15, 14) */,
  32'h3e1c2ca1 /* (4, 15, 14) */,
  32'h3e05899d /* (0, 15, 14) */,
  32'h3ddc0819 /* (28, 11, 14) */,
  32'h3e2a27e4 /* (24, 11, 14) */,
  32'h3e9ecc49 /* (20, 11, 14) */,
  32'h3ec4f0a1 /* (16, 11, 14) */,
  32'h3e9ecc49 /* (12, 11, 14) */,
  32'h3e2a27e4 /* (8, 11, 14) */,
  32'h3ddc0819 /* (4, 11, 14) */,
  32'h3dbe661f /* (0, 11, 14) */,
  32'h3d800deb /* (28, 7, 14) */,
  32'h3dbf672f /* (24, 7, 14) */,
  32'h3e2baf50 /* (20, 7, 14) */,
  32'h3e4d7ce8 /* (16, 7, 14) */,
  32'h3e2baf50 /* (12, 7, 14) */,
  32'h3dbf672f /* (8, 7, 14) */,
  32'h3d800deb /* (4, 7, 14) */,
  32'h3d60bf24 /* (0, 7, 14) */,
  32'h3d3b1e93 /* (28, 3, 14) */,
  32'h3d880501 /* (24, 3, 14) */,
  32'h3decc5e8 /* (20, 3, 14) */,
  32'h3e0a27e7 /* (16, 3, 14) */,
  32'h3decc5e8 /* (12, 3, 14) */,
  32'h3d880501 /* (8, 3, 14) */,
  32'h3d3b1e93 /* (4, 3, 14) */,
  32'h3d262b6e /* (0, 3, 14) */,
  32'h3d1839e3 /* (28, 31, 10) */,
  32'h3d3f0366 /* (24, 31, 10) */,
  32'h3d91435f /* (20, 31, 10) */,
  32'h3d99ac24 /* (16, 31, 10) */,
  32'h3d91435f /* (12, 31, 10) */,
  32'h3d3f0366 /* (8, 31, 10) */,
  32'h3d1839e3 /* (4, 31, 10) */,
  32'h3d1142bb /* (0, 31, 10) */,
  32'h3d28e3b2 /* (28, 27, 10) */,
  32'h3d5ef675 /* (24, 27, 10) */,
  32'h3db0e528 /* (20, 27, 10) */,
  32'h3dc0863e /* (16, 27, 10) */,
  32'h3db0e528 /* (12, 27, 10) */,
  32'h3d5ef675 /* (8, 27, 10) */,
  32'h3d28e3b2 /* (4, 27, 10) */,
  32'h3d1cee15 /* (0, 27, 10) */,
  32'h3d68b7a2 /* (28, 23, 10) */,
  32'h3da590e9 /* (24, 23, 10) */,
  32'h3e0cf021 /* (20, 23, 10) */,
  32'h3e21930d /* (16, 23, 10) */,
  32'h3e0cf021 /* (12, 23, 10) */,
  32'h3da590e9 /* (8, 23, 10) */,
  32'h3d68b7a2 /* (4, 23, 10) */,
  32'h3d50a575 /* (0, 23, 10) */,
  32'h3db40e50 /* (28, 19, 10) */,
  32'h3e085939 /* (24, 19, 10) */,
  32'h3e7848b5 /* (20, 19, 10) */,
  32'h3e968a40 /* (16, 19, 10) */,
  32'h3e7848b5 /* (12, 19, 10) */,
  32'h3e085939 /* (8, 19, 10) */,
  32'h3db40e50 /* (4, 19, 10) */,
  32'h3d9d248b /* (0, 19, 10) */,
  32'h3dbdf4f8 /* (28, 15, 10) */,
  32'h3e135573 /* (24, 15, 10) */,
  32'h3e89fde5 /* (20, 15, 10) */,
  32'h3eabb572 /* (16, 15, 10) */,
  32'h3e89fde5 /* (12, 15, 10) */,
  32'h3e135573 /* (8, 15, 10) */,
  32'h3dbdf4f8 /* (4, 15, 10) */,
  32'h3da42e1b /* (0, 15, 10) */,
  32'h3d92b699 /* (28, 11, 10) */,
  32'h3dd7e578 /* (24, 11, 10) */,
  32'h3e3e5baf /* (20, 11, 10) */,
  32'h3e60898b /* (16, 11, 10) */,
  32'h3e3e5baf /* (12, 11, 10) */,
  32'h3dd7e578 /* (8, 11, 10) */,
  32'h3d92b699 /* (4, 11, 10) */,
  32'h3d819abc /* (0, 11, 10) */,
  32'h3d404057 /* (28, 7, 10) */,
  32'h3d83c517 /* (24, 7, 10) */,
  32'h3dd85675 /* (20, 7, 10) */,
  32'h3df142da /* (16, 7, 10) */,
  32'h3dd85675 /* (12, 7, 10) */,
  32'h3d83c517 /* (8, 7, 10) */,
  32'h3d404057 /* (4, 7, 10) */,
  32'h3d2f5f5a /* (0, 7, 10) */,
  32'h3d1cff11 /* (28, 3, 10) */,
  32'h3d48bc7e /* (24, 3, 10) */,
  32'h3d9aff71 /* (20, 3, 10) */,
  32'h3da59d10 /* (16, 3, 10) */,
  32'h3d9aff71 /* (12, 3, 10) */,
  32'h3d48bc7e /* (8, 3, 10) */,
  32'h3d1cff11 /* (4, 3, 10) */,
  32'h3d144f19 /* (0, 3, 10) */,
  32'h3d222a9c /* (28, 31, 6) */,
  32'h3d169650 /* (24, 31, 6) */,
  32'h3d3dc5f0 /* (20, 31, 6) */,
  32'h3d34b66a /* (16, 31, 6) */,
  32'h3d3dc5f0 /* (12, 31, 6) */,
  32'h3d169650 /* (8, 31, 6) */,
  32'h3d222a9c /* (4, 31, 6) */,
  32'h3d3f59b8 /* (0, 31, 6) */,
  32'h3d153e19 /* (28, 27, 6) */,
  32'h3d22af34 /* (24, 27, 6) */,
  32'h3d6007ad /* (20, 27, 6) */,
  32'h3d5f53fb /* (16, 27, 6) */,
  32'h3d6007ad /* (12, 27, 6) */,
  32'h3d22af34 /* (8, 27, 6) */,
  32'h3d153e19 /* (4, 27, 6) */,
  32'h3d1b2f33 /* (0, 27, 6) */,
  32'h3d2657dd /* (28, 23, 6) */,
  32'h3d584c0c /* (24, 23, 6) */,
  32'h3da96159 /* (20, 23, 6) */,
  32'h3db6b309 /* (16, 23, 6) */,
  32'h3da96159 /* (12, 23, 6) */,
  32'h3d584c0c /* (8, 23, 6) */,
  32'h3d2657dd /* (4, 23, 6) */,
  32'h3d1bc36a /* (0, 23, 6) */,
  32'h3d601ae9 /* (28, 19, 6) */,
  32'h3da2e7a9 /* (24, 19, 6) */,
  32'h3e0dc95f /* (20, 19, 6) */,
  32'h3e2576a9 /* (16, 19, 6) */,
  32'h3e0dc95f /* (12, 19, 6) */,
  32'h3da2e7a9 /* (8, 19, 6) */,
  32'h3d601ae9 /* (4, 19, 6) */,
  32'h3d4703b2 /* (0, 19, 6) */,
  32'h3d61b1de /* (28, 15, 6) */,
  32'h3daa3349 /* (24, 15, 6) */,
  32'h3e1a3a56 /* (20, 15, 6) */,
  32'h3e3a3d1a /* (16, 15, 6) */,
  32'h3e1a3a56 /* (12, 15, 6) */,
  32'h3daa3349 /* (8, 15, 6) */,
  32'h3d61b1de /* (4, 15, 6) */,
  32'h3d455011 /* (0, 15, 6) */,
  32'h3d41fb9f /* (28, 11, 6) */,
  32'h3d865b59 /* (24, 11, 6) */,
  32'h3ddec971 /* (20, 11, 6) */,
  32'h3dfa4afe /* (16, 11, 6) */,
  32'h3ddec971 /* (12, 11, 6) */,
  32'h3d865b59 /* (8, 11, 6) */,
  32'h3d41fb9f /* (4, 11, 6) */,
  32'h3d3013e2 /* (0, 11, 6) */,
  32'h3d17902e /* (28, 7, 6) */,
  32'h3d35cd98 /* (24, 7, 6) */,
  32'h3d859348 /* (20, 7, 6) */,
  32'h3d8a46e7 /* (16, 7, 6) */,
  32'h3d859348 /* (12, 7, 6) */,
  32'h3d35cd98 /* (8, 7, 6) */,
  32'h3d17902e /* (4, 7, 6) */,
  32'h3d1459dd /* (0, 7, 6) */,
  32'h3d1b3fff /* (28, 3, 6) */,
  32'h3d19bf4b /* (24, 3, 6) */,
  32'h3d48406d /* (20, 3, 6) */,
  32'h3d41d3ae /* (16, 3, 6) */,
  32'h3d48406d /* (12, 3, 6) */,
  32'h3d19bf4b /* (8, 3, 6) */,
  32'h3d1b3fff /* (4, 3, 6) */,
  32'h3d2d5b95 /* (0, 3, 6) */,
  32'h3d8b1391 /* (28, 31, 2) */,
  32'h3d15ce12 /* (24, 31, 2) */,
  32'h3d1cac31 /* (20, 31, 2) */,
  32'h3d09dfab /* (16, 31, 2) */,
  32'h3d1cac31 /* (12, 31, 2) */,
  32'h3d15ce12 /* (8, 31, 2) */,
  32'h3d8b1391 /* (4, 31, 2) */,
  32'h3e709592 /* (0, 31, 2) */,
  32'h3d2d8e0e /* (28, 27, 2) */,
  32'h3d149b5c /* (24, 27, 2) */,
  32'h3d346b02 /* (20, 27, 2) */,
  32'h3d28d1e5 /* (16, 27, 2) */,
  32'h3d346b02 /* (12, 27, 2) */,
  32'h3d149b5c /* (8, 27, 2) */,
  32'h3d2d8e0e /* (4, 27, 2) */,
  32'h3d5dd7d1 /* (0, 27, 2) */,
  32'h3d14de35 /* (28, 23, 2) */,
  32'h3d3291f6 /* (24, 23, 2) */,
  32'h3d833332 /* (20, 23, 2) */,
  32'h3d87d16b /* (16, 23, 2) */,
  32'h3d833332 /* (12, 23, 2) */,
  32'h3d3291f6 /* (8, 23, 2) */,
  32'h3d14de35 /* (4, 23, 2) */,
  32'h3d11b684 /* (0, 23, 2) */,
  32'h3d3217f4 /* (28, 19, 2) */,
  32'h3d7b52f8 /* (24, 19, 2) */,
  32'h3dd42d31 /* (20, 19, 2) */,
  32'h3df1ae3d /* (16, 19, 2) */,
  32'h3dd42d31 /* (12, 19, 2) */,
  32'h3d7b52f8 /* (8, 19, 2) */,
  32'h3d3217f4 /* (4, 19, 2) */,
  32'h3d2045b1 /* (0, 19, 2) */,
  32'h3d2d6bba /* (28, 15, 2) */,
  32'h3d804df8 /* (24, 15, 2) */,
  32'h3de39dff /* (20, 15, 2) */,
  32'h3e06ec2e /* (16, 15, 2) */,
  32'h3de39dff /* (12, 15, 2) */,
  32'h3d804df8 /* (8, 15, 2) */,
  32'h3d2d6bba /* (4, 15, 2) */,
  32'h3d18d610 /* (0, 15, 2) */,
  32'h3d21c128 /* (28, 11, 2) */,
  32'h3d558b1c /* (24, 11, 2) */,
  32'h3da96c08 /* (20, 11, 2) */,
  32'h3db86416 /* (16, 11, 2) */,
  32'h3da96c08 /* (12, 11, 2) */,
  32'h3d558b1c /* (8, 11, 2) */,
  32'h3d21c128 /* (4, 11, 2) */,
  32'h3d164ce1 /* (0, 11, 2) */,
  32'h3d16c6a3 /* (28, 7, 2) */,
  32'h3d1d59b0 /* (24, 7, 2) */,
  32'h3d530d8e /* (20, 7, 2) */,
  32'h3d4f6a6e /* (16, 7, 2) */,
  32'h3d530d8e /* (12, 7, 2) */,
  32'h3d1d59b0 /* (8, 7, 2) */,
  32'h3d16c6a3 /* (4, 7, 2) */,
  32'h3d21b235 /* (0, 7, 2) */,
  32'h3d5defd3 /* (28, 3, 2) */,
  32'h3d13e9f7 /* (24, 3, 2) */,
  32'h3d23d587 /* (20, 3, 2) */,
  32'h3d13661d /* (16, 3, 2) */,
  32'h3d23d587 /* (12, 3, 2) */,
  32'h3d13e9f7 /* (8, 3, 2) */,
  32'h3d5defd3 /* (4, 3, 2) */,
  32'h3dcbea25 /* (0, 3, 2) */,
  32'h3e0c4d23 /* (31, 30, 30) */,
  32'h3d4ca49b /* (27, 30, 30) */,
  32'h3d1214c5 /* (23, 30, 30) */,
  32'h3d246fbd /* (19, 30, 30) */,
  32'h3d1dadb9 /* (15, 30, 30) */,
  32'h3d18e0f8 /* (11, 30, 30) */,
  32'h3d1dd271 /* (7, 30, 30) */,
  32'h3da3af74 /* (3, 30, 30) */,
  32'h3d3543e4 /* (31, 26, 30) */,
  32'h3d18df8d /* (27, 26, 30) */,
  32'h3d1e19af /* (23, 26, 30) */,
  32'h3d4ce87b /* (19, 26, 30) */,
  32'h3d4bfe66 /* (15, 26, 30) */,
  32'h3d343ccb /* (11, 26, 30) */,
  32'h3d14b9d3 /* (7, 26, 30) */,
  32'h3d271e8d /* (3, 26, 30) */,
  32'h3d12ac07 /* (31, 22, 30) */,
  32'h3d1f9f49 /* (27, 22, 30) */,
  32'h3d56480e /* (23, 22, 30) */,
  32'h3da2895a /* (19, 22, 30) */,
  32'h3daa3ec9 /* (15, 22, 30) */,
  32'h3d85a0b3 /* (11, 22, 30) */,
  32'h3d3346c6 /* (7, 22, 30) */,
  32'h3d162b76 /* (3, 22, 30) */,
  32'h3d217487 /* (31, 18, 30) */,
  32'h3d40d8bf /* (27, 18, 30) */,
  32'h3d94a37c /* (23, 18, 30) */,
  32'h3dfd653f /* (19, 18, 30) */,
  32'h3e0adb0d /* (15, 18, 30) */,
  32'h3dc55f41 /* (11, 18, 30) */,
  32'h3d6820b1 /* (7, 18, 30) */,
  32'h3d2b1735 /* (3, 18, 30) */,
  32'h3d217487 /* (31, 14, 30) */,
  32'h3d40d8bf /* (27, 14, 30) */,
  32'h3d94a37c /* (23, 14, 30) */,
  32'h3dfd653f /* (19, 14, 30) */,
  32'h3e0adb0d /* (15, 14, 30) */,
  32'h3dc55f41 /* (11, 14, 30) */,
  32'h3d6820b1 /* (7, 14, 30) */,
  32'h3d2b1735 /* (3, 14, 30) */,
  32'h3d12ac07 /* (31, 10, 30) */,
  32'h3d1f9f49 /* (27, 10, 30) */,
  32'h3d56480e /* (23, 10, 30) */,
  32'h3da2895a /* (19, 10, 30) */,
  32'h3daa3ec9 /* (15, 10, 30) */,
  32'h3d85a0b3 /* (11, 10, 30) */,
  32'h3d3346c6 /* (7, 10, 30) */,
  32'h3d162b76 /* (3, 10, 30) */,
  32'h3d3543e4 /* (31, 6, 30) */,
  32'h3d18df8d /* (27, 6, 30) */,
  32'h3d1e19af /* (23, 6, 30) */,
  32'h3d4ce87b /* (19, 6, 30) */,
  32'h3d4bfe66 /* (15, 6, 30) */,
  32'h3d343ccb /* (11, 6, 30) */,
  32'h3d14b9d3 /* (7, 6, 30) */,
  32'h3d271e8d /* (3, 6, 30) */,
  32'h3e0c4d23 /* (31, 2, 30) */,
  32'h3d4ca49b /* (27, 2, 30) */,
  32'h3d1214c5 /* (23, 2, 30) */,
  32'h3d246fbd /* (19, 2, 30) */,
  32'h3d1dadb9 /* (15, 2, 30) */,
  32'h3d18e0f8 /* (11, 2, 30) */,
  32'h3d1dd271 /* (7, 2, 30) */,
  32'h3da3af74 /* (3, 2, 30) */,
  32'h3d3543e4 /* (31, 30, 26) */,
  32'h3d18df8d /* (27, 30, 26) */,
  32'h3d1e19af /* (23, 30, 26) */,
  32'h3d4ce87b /* (19, 30, 26) */,
  32'h3d4bfe66 /* (15, 30, 26) */,
  32'h3d343ccb /* (11, 30, 26) */,
  32'h3d14b9d3 /* (7, 30, 26) */,
  32'h3d271e8d /* (3, 30, 26) */,
  32'h3d15cc97 /* (31, 26, 26) */,
  32'h3d16bb8b /* (27, 26, 26) */,
  32'h3d37f9d0 /* (23, 26, 26) */,
  32'h3d82bc35 /* (19, 26, 26) */,
  32'h3d85e8bf /* (15, 26, 26) */,
  32'h3d5d3b5c /* (11, 26, 26) */,
  32'h3d20f672 /* (7, 26, 26) */,
  32'h3d14c14d /* (3, 26, 26) */,
  32'h3d2567ce /* (31, 22, 26) */,
  32'h3d3c300c /* (27, 22, 26) */,
  32'h3d866682 /* (23, 22, 26) */,
  32'h3dd610ea /* (19, 22, 26) */,
  32'h3de44bb3 /* (15, 22, 26) */,
  32'h3dac23aa /* (11, 22, 26) */,
  32'h3d5a2934 /* (7, 22, 26) */,
  32'h3d2c3293 /* (3, 22, 26) */,
  32'h3d4cf093 /* (31, 18, 26) */,
  32'h3d786cd6 /* (27, 18, 26) */,
  32'h3dc45939 /* (23, 18, 26) */,
  32'h3e2b8c37 /* (19, 18, 26) */,
  32'h3e3e01e0 /* (15, 18, 26) */,
  32'h3e040b60 /* (11, 18, 26) */,
  32'h3d975464 /* (7, 18, 26) */,
  32'h3d5a5169 /* (3, 18, 26) */,
  32'h3d4cf093 /* (31, 14, 26) */,
  32'h3d786cd6 /* (27, 14, 26) */,
  32'h3dc45939 /* (23, 14, 26) */,
  32'h3e2b8c37 /* (19, 14, 26) */,
  32'h3e3e01e0 /* (15, 14, 26) */,
  32'h3e040b60 /* (11, 14, 26) */,
  32'h3d975464 /* (7, 14, 26) */,
  32'h3d5a5169 /* (3, 14, 26) */,
  32'h3d2567ce /* (31, 10, 26) */,
  32'h3d3c300c /* (27, 10, 26) */,
  32'h3d866682 /* (23, 10, 26) */,
  32'h3dd610ea /* (19, 10, 26) */,
  32'h3de44bb3 /* (15, 10, 26) */,
  32'h3dac23aa /* (11, 10, 26) */,
  32'h3d5a2934 /* (7, 10, 26) */,
  32'h3d2c3293 /* (3, 10, 26) */,
  32'h3d15cc97 /* (31, 6, 26) */,
  32'h3d16bb8b /* (27, 6, 26) */,
  32'h3d37f9d0 /* (23, 6, 26) */,
  32'h3d82bc35 /* (19, 6, 26) */,
  32'h3d85e8bf /* (15, 6, 26) */,
  32'h3d5d3b5c /* (11, 6, 26) */,
  32'h3d20f672 /* (7, 6, 26) */,
  32'h3d14c14d /* (3, 6, 26) */,
  32'h3d3543e4 /* (31, 2, 26) */,
  32'h3d18df8d /* (27, 2, 26) */,
  32'h3d1e19af /* (23, 2, 26) */,
  32'h3d4ce87b /* (19, 2, 26) */,
  32'h3d4bfe66 /* (15, 2, 26) */,
  32'h3d343ccb /* (11, 2, 26) */,
  32'h3d14b9d3 /* (7, 2, 26) */,
  32'h3d271e8d /* (3, 2, 26) */,
  32'h3d12ac07 /* (31, 30, 22) */,
  32'h3d1f9f49 /* (27, 30, 22) */,
  32'h3d56480e /* (23, 30, 22) */,
  32'h3da2895a /* (19, 30, 22) */,
  32'h3daa3ec9 /* (15, 30, 22) */,
  32'h3d85a0b3 /* (11, 30, 22) */,
  32'h3d3346c6 /* (7, 30, 22) */,
  32'h3d162b76 /* (3, 30, 22) */,
  32'h3d2567ce /* (31, 26, 22) */,
  32'h3d3c300c /* (27, 26, 22) */,
  32'h3d866682 /* (23, 26, 22) */,
  32'h3dd610ea /* (19, 26, 22) */,
  32'h3de44bb3 /* (15, 26, 22) */,
  32'h3dac23aa /* (11, 26, 22) */,
  32'h3d5a2934 /* (7, 26, 22) */,
  32'h3d2c3293 /* (3, 26, 22) */,
  32'h3d699f13 /* (31, 22, 22) */,
  32'h3d8b85a2 /* (27, 22, 22) */,
  32'h3dd7137d /* (23, 22, 22) */,
  32'h3e37540b /* (19, 22, 22) */,
  32'h3e48eba4 /* (15, 22, 22) */,
  32'h3e0ecbcd /* (11, 22, 22) */,
  32'h3da7f0fb /* (7, 22, 22) */,
  32'h3d77904c /* (3, 22, 22) */,
  32'h3da6958f /* (31, 18, 22) */,
  32'h3dce13fe /* (27, 18, 22) */,
  32'h3e28e750 /* (23, 18, 22) */,
  32'h3e994798 /* (19, 18, 22) */,
  32'h3eacaf9b /* (15, 18, 22) */,
  32'h3e67a191 /* (11, 18, 22) */,
  32'h3dff6ab3 /* (7, 18, 22) */,
  32'h3db2bcb9 /* (3, 18, 22) */,
  32'h3da6958f /* (31, 14, 22) */,
  32'h3dce13fe /* (27, 14, 22) */,
  32'h3e28e750 /* (23, 14, 22) */,
  32'h3e994798 /* (19, 14, 22) */,
  32'h3eacaf9b /* (15, 14, 22) */,
  32'h3e67a191 /* (11, 14, 22) */,
  32'h3dff6ab3 /* (7, 14, 22) */,
  32'h3db2bcb9 /* (3, 14, 22) */,
  32'h3d699f13 /* (31, 10, 22) */,
  32'h3d8b85a2 /* (27, 10, 22) */,
  32'h3dd7137d /* (23, 10, 22) */,
  32'h3e37540b /* (19, 10, 22) */,
  32'h3e48eba4 /* (15, 10, 22) */,
  32'h3e0ecbcd /* (11, 10, 22) */,
  32'h3da7f0fb /* (7, 10, 22) */,
  32'h3d77904c /* (3, 10, 22) */,
  32'h3d2567ce /* (31, 6, 22) */,
  32'h3d3c300c /* (27, 6, 22) */,
  32'h3d866682 /* (23, 6, 22) */,
  32'h3dd610ea /* (19, 6, 22) */,
  32'h3de44bb3 /* (15, 6, 22) */,
  32'h3dac23aa /* (11, 6, 22) */,
  32'h3d5a2934 /* (7, 6, 22) */,
  32'h3d2c3293 /* (3, 6, 22) */,
  32'h3d12ac07 /* (31, 2, 22) */,
  32'h3d1f9f49 /* (27, 2, 22) */,
  32'h3d56480e /* (23, 2, 22) */,
  32'h3da2895a /* (19, 2, 22) */,
  32'h3daa3ec9 /* (15, 2, 22) */,
  32'h3d85a0b3 /* (11, 2, 22) */,
  32'h3d3346c6 /* (7, 2, 22) */,
  32'h3d162b76 /* (3, 2, 22) */,
  32'h3d217487 /* (31, 30, 18) */,
  32'h3d40d8bf /* (27, 30, 18) */,
  32'h3d94a37c /* (23, 30, 18) */,
  32'h3dfd653f /* (19, 30, 18) */,
  32'h3e0adb0d /* (15, 30, 18) */,
  32'h3dc55f41 /* (11, 30, 18) */,
  32'h3d6820b1 /* (7, 30, 18) */,
  32'h3d2b1735 /* (3, 30, 18) */,
  32'h3d4cf093 /* (31, 26, 18) */,
  32'h3d786cd6 /* (27, 26, 18) */,
  32'h3dc45939 /* (23, 26, 18) */,
  32'h3e2b8c37 /* (19, 26, 18) */,
  32'h3e3e01e0 /* (15, 26, 18) */,
  32'h3e040b60 /* (11, 26, 18) */,
  32'h3d975464 /* (7, 26, 18) */,
  32'h3d5a5169 /* (3, 26, 18) */,
  32'h3da6958f /* (31, 22, 18) */,
  32'h3dce13fe /* (27, 22, 18) */,
  32'h3e28e750 /* (23, 22, 18) */,
  32'h3e994798 /* (19, 22, 18) */,
  32'h3eacaf9b /* (15, 22, 18) */,
  32'h3e67a191 /* (11, 22, 18) */,
  32'h3dff6ab3 /* (7, 22, 18) */,
  32'h3db2bcb9 /* (3, 22, 18) */,
  32'h3e04a438 /* (31, 18, 18) */,
  32'h3e27240a /* (27, 18, 18) */,
  32'h3e8dd733 /* (23, 18, 18) */,
  32'h3f05dc96 /* (19, 18, 18) */,
  32'h3f19a2a7 /* (15, 18, 18) */,
  32'h3ec66134 /* (11, 18, 18) */,
  32'h3e528761 /* (7, 18, 18) */,
  32'h3e0f3c67 /* (3, 18, 18) */,
  32'h3e04a438 /* (31, 14, 18) */,
  32'h3e27240a /* (27, 14, 18) */,
  32'h3e8dd733 /* (23, 14, 18) */,
  32'h3f05dc96 /* (19, 14, 18) */,
  32'h3f19a2a7 /* (15, 14, 18) */,
  32'h3ec66134 /* (11, 14, 18) */,
  32'h3e528761 /* (7, 14, 18) */,
  32'h3e0f3c67 /* (3, 14, 18) */,
  32'h3da6958f /* (31, 10, 18) */,
  32'h3dce13fe /* (27, 10, 18) */,
  32'h3e28e750 /* (23, 10, 18) */,
  32'h3e994798 /* (19, 10, 18) */,
  32'h3eacaf9b /* (15, 10, 18) */,
  32'h3e67a191 /* (11, 10, 18) */,
  32'h3dff6ab3 /* (7, 10, 18) */,
  32'h3db2bcb9 /* (3, 10, 18) */,
  32'h3d4cf093 /* (31, 6, 18) */,
  32'h3d786cd6 /* (27, 6, 18) */,
  32'h3dc45939 /* (23, 6, 18) */,
  32'h3e2b8c37 /* (19, 6, 18) */,
  32'h3e3e01e0 /* (15, 6, 18) */,
  32'h3e040b60 /* (11, 6, 18) */,
  32'h3d975464 /* (7, 6, 18) */,
  32'h3d5a5169 /* (3, 6, 18) */,
  32'h3d217487 /* (31, 2, 18) */,
  32'h3d40d8bf /* (27, 2, 18) */,
  32'h3d94a37c /* (23, 2, 18) */,
  32'h3dfd653f /* (19, 2, 18) */,
  32'h3e0adb0d /* (15, 2, 18) */,
  32'h3dc55f41 /* (11, 2, 18) */,
  32'h3d6820b1 /* (7, 2, 18) */,
  32'h3d2b1735 /* (3, 2, 18) */,
  32'h3d217487 /* (31, 30, 14) */,
  32'h3d40d8bf /* (27, 30, 14) */,
  32'h3d94a37c /* (23, 30, 14) */,
  32'h3dfd653f /* (19, 30, 14) */,
  32'h3e0adb0d /* (15, 30, 14) */,
  32'h3dc55f41 /* (11, 30, 14) */,
  32'h3d6820b1 /* (7, 30, 14) */,
  32'h3d2b1735 /* (3, 30, 14) */,
  32'h3d4cf093 /* (31, 26, 14) */,
  32'h3d786cd6 /* (27, 26, 14) */,
  32'h3dc45939 /* (23, 26, 14) */,
  32'h3e2b8c37 /* (19, 26, 14) */,
  32'h3e3e01e0 /* (15, 26, 14) */,
  32'h3e040b60 /* (11, 26, 14) */,
  32'h3d975464 /* (7, 26, 14) */,
  32'h3d5a5169 /* (3, 26, 14) */,
  32'h3da6958f /* (31, 22, 14) */,
  32'h3dce13fe /* (27, 22, 14) */,
  32'h3e28e750 /* (23, 22, 14) */,
  32'h3e994798 /* (19, 22, 14) */,
  32'h3eacaf9b /* (15, 22, 14) */,
  32'h3e67a191 /* (11, 22, 14) */,
  32'h3dff6ab3 /* (7, 22, 14) */,
  32'h3db2bcb9 /* (3, 22, 14) */,
  32'h3e04a438 /* (31, 18, 14) */,
  32'h3e27240a /* (27, 18, 14) */,
  32'h3e8dd733 /* (23, 18, 14) */,
  32'h3f05dc96 /* (19, 18, 14) */,
  32'h3f19a2a7 /* (15, 18, 14) */,
  32'h3ec66134 /* (11, 18, 14) */,
  32'h3e528761 /* (7, 18, 14) */,
  32'h3e0f3c67 /* (3, 18, 14) */,
  32'h3e04a438 /* (31, 14, 14) */,
  32'h3e27240a /* (27, 14, 14) */,
  32'h3e8dd733 /* (23, 14, 14) */,
  32'h3f05dc96 /* (19, 14, 14) */,
  32'h3f19a2a7 /* (15, 14, 14) */,
  32'h3ec66134 /* (11, 14, 14) */,
  32'h3e528761 /* (7, 14, 14) */,
  32'h3e0f3c67 /* (3, 14, 14) */,
  32'h3da6958f /* (31, 10, 14) */,
  32'h3dce13fe /* (27, 10, 14) */,
  32'h3e28e750 /* (23, 10, 14) */,
  32'h3e994798 /* (19, 10, 14) */,
  32'h3eacaf9b /* (15, 10, 14) */,
  32'h3e67a191 /* (11, 10, 14) */,
  32'h3dff6ab3 /* (7, 10, 14) */,
  32'h3db2bcb9 /* (3, 10, 14) */,
  32'h3d4cf093 /* (31, 6, 14) */,
  32'h3d786cd6 /* (27, 6, 14) */,
  32'h3dc45939 /* (23, 6, 14) */,
  32'h3e2b8c37 /* (19, 6, 14) */,
  32'h3e3e01e0 /* (15, 6, 14) */,
  32'h3e040b60 /* (11, 6, 14) */,
  32'h3d975464 /* (7, 6, 14) */,
  32'h3d5a5169 /* (3, 6, 14) */,
  32'h3d217487 /* (31, 2, 14) */,
  32'h3d40d8bf /* (27, 2, 14) */,
  32'h3d94a37c /* (23, 2, 14) */,
  32'h3dfd653f /* (19, 2, 14) */,
  32'h3e0adb0d /* (15, 2, 14) */,
  32'h3dc55f41 /* (11, 2, 14) */,
  32'h3d6820b1 /* (7, 2, 14) */,
  32'h3d2b1735 /* (3, 2, 14) */,
  32'h3d12ac07 /* (31, 30, 10) */,
  32'h3d1f9f49 /* (27, 30, 10) */,
  32'h3d56480e /* (23, 30, 10) */,
  32'h3da2895a /* (19, 30, 10) */,
  32'h3daa3ec9 /* (15, 30, 10) */,
  32'h3d85a0b3 /* (11, 30, 10) */,
  32'h3d3346c6 /* (7, 30, 10) */,
  32'h3d162b76 /* (3, 30, 10) */,
  32'h3d2567ce /* (31, 26, 10) */,
  32'h3d3c300c /* (27, 26, 10) */,
  32'h3d866682 /* (23, 26, 10) */,
  32'h3dd610ea /* (19, 26, 10) */,
  32'h3de44bb3 /* (15, 26, 10) */,
  32'h3dac23aa /* (11, 26, 10) */,
  32'h3d5a2934 /* (7, 26, 10) */,
  32'h3d2c3293 /* (3, 26, 10) */,
  32'h3d699f13 /* (31, 22, 10) */,
  32'h3d8b85a2 /* (27, 22, 10) */,
  32'h3dd7137d /* (23, 22, 10) */,
  32'h3e37540b /* (19, 22, 10) */,
  32'h3e48eba4 /* (15, 22, 10) */,
  32'h3e0ecbcd /* (11, 22, 10) */,
  32'h3da7f0fb /* (7, 22, 10) */,
  32'h3d77904c /* (3, 22, 10) */,
  32'h3da6958f /* (31, 18, 10) */,
  32'h3dce13fe /* (27, 18, 10) */,
  32'h3e28e750 /* (23, 18, 10) */,
  32'h3e994798 /* (19, 18, 10) */,
  32'h3eacaf9b /* (15, 18, 10) */,
  32'h3e67a191 /* (11, 18, 10) */,
  32'h3dff6ab3 /* (7, 18, 10) */,
  32'h3db2bcb9 /* (3, 18, 10) */,
  32'h3da6958f /* (31, 14, 10) */,
  32'h3dce13fe /* (27, 14, 10) */,
  32'h3e28e750 /* (23, 14, 10) */,
  32'h3e994798 /* (19, 14, 10) */,
  32'h3eacaf9b /* (15, 14, 10) */,
  32'h3e67a191 /* (11, 14, 10) */,
  32'h3dff6ab3 /* (7, 14, 10) */,
  32'h3db2bcb9 /* (3, 14, 10) */,
  32'h3d699f13 /* (31, 10, 10) */,
  32'h3d8b85a2 /* (27, 10, 10) */,
  32'h3dd7137d /* (23, 10, 10) */,
  32'h3e37540b /* (19, 10, 10) */,
  32'h3e48eba4 /* (15, 10, 10) */,
  32'h3e0ecbcd /* (11, 10, 10) */,
  32'h3da7f0fb /* (7, 10, 10) */,
  32'h3d77904c /* (3, 10, 10) */,
  32'h3d2567ce /* (31, 6, 10) */,
  32'h3d3c300c /* (27, 6, 10) */,
  32'h3d866682 /* (23, 6, 10) */,
  32'h3dd610ea /* (19, 6, 10) */,
  32'h3de44bb3 /* (15, 6, 10) */,
  32'h3dac23aa /* (11, 6, 10) */,
  32'h3d5a2934 /* (7, 6, 10) */,
  32'h3d2c3293 /* (3, 6, 10) */,
  32'h3d12ac07 /* (31, 2, 10) */,
  32'h3d1f9f49 /* (27, 2, 10) */,
  32'h3d56480e /* (23, 2, 10) */,
  32'h3da2895a /* (19, 2, 10) */,
  32'h3daa3ec9 /* (15, 2, 10) */,
  32'h3d85a0b3 /* (11, 2, 10) */,
  32'h3d3346c6 /* (7, 2, 10) */,
  32'h3d162b76 /* (3, 2, 10) */,
  32'h3d3543e4 /* (31, 30, 6) */,
  32'h3d18df8d /* (27, 30, 6) */,
  32'h3d1e19af /* (23, 30, 6) */,
  32'h3d4ce87b /* (19, 30, 6) */,
  32'h3d4bfe66 /* (15, 30, 6) */,
  32'h3d343ccb /* (11, 30, 6) */,
  32'h3d14b9d3 /* (7, 30, 6) */,
  32'h3d271e8d /* (3, 30, 6) */,
  32'h3d15cc97 /* (31, 26, 6) */,
  32'h3d16bb8b /* (27, 26, 6) */,
  32'h3d37f9d0 /* (23, 26, 6) */,
  32'h3d82bc35 /* (19, 26, 6) */,
  32'h3d85e8bf /* (15, 26, 6) */,
  32'h3d5d3b5c /* (11, 26, 6) */,
  32'h3d20f672 /* (7, 26, 6) */,
  32'h3d14c14d /* (3, 26, 6) */,
  32'h3d2567ce /* (31, 22, 6) */,
  32'h3d3c300c /* (27, 22, 6) */,
  32'h3d866682 /* (23, 22, 6) */,
  32'h3dd610ea /* (19, 22, 6) */,
  32'h3de44bb3 /* (15, 22, 6) */,
  32'h3dac23aa /* (11, 22, 6) */,
  32'h3d5a2934 /* (7, 22, 6) */,
  32'h3d2c3293 /* (3, 22, 6) */,
  32'h3d4cf093 /* (31, 18, 6) */,
  32'h3d786cd6 /* (27, 18, 6) */,
  32'h3dc45939 /* (23, 18, 6) */,
  32'h3e2b8c37 /* (19, 18, 6) */,
  32'h3e3e01e0 /* (15, 18, 6) */,
  32'h3e040b60 /* (11, 18, 6) */,
  32'h3d975464 /* (7, 18, 6) */,
  32'h3d5a5169 /* (3, 18, 6) */,
  32'h3d4cf093 /* (31, 14, 6) */,
  32'h3d786cd6 /* (27, 14, 6) */,
  32'h3dc45939 /* (23, 14, 6) */,
  32'h3e2b8c37 /* (19, 14, 6) */,
  32'h3e3e01e0 /* (15, 14, 6) */,
  32'h3e040b60 /* (11, 14, 6) */,
  32'h3d975464 /* (7, 14, 6) */,
  32'h3d5a5169 /* (3, 14, 6) */,
  32'h3d2567ce /* (31, 10, 6) */,
  32'h3d3c300c /* (27, 10, 6) */,
  32'h3d866682 /* (23, 10, 6) */,
  32'h3dd610ea /* (19, 10, 6) */,
  32'h3de44bb3 /* (15, 10, 6) */,
  32'h3dac23aa /* (11, 10, 6) */,
  32'h3d5a2934 /* (7, 10, 6) */,
  32'h3d2c3293 /* (3, 10, 6) */,
  32'h3d15cc97 /* (31, 6, 6) */,
  32'h3d16bb8b /* (27, 6, 6) */,
  32'h3d37f9d0 /* (23, 6, 6) */,
  32'h3d82bc35 /* (19, 6, 6) */,
  32'h3d85e8bf /* (15, 6, 6) */,
  32'h3d5d3b5c /* (11, 6, 6) */,
  32'h3d20f672 /* (7, 6, 6) */,
  32'h3d14c14d /* (3, 6, 6) */,
  32'h3d3543e4 /* (31, 2, 6) */,
  32'h3d18df8d /* (27, 2, 6) */,
  32'h3d1e19af /* (23, 2, 6) */,
  32'h3d4ce87b /* (19, 2, 6) */,
  32'h3d4bfe66 /* (15, 2, 6) */,
  32'h3d343ccb /* (11, 2, 6) */,
  32'h3d14b9d3 /* (7, 2, 6) */,
  32'h3d271e8d /* (3, 2, 6) */,
  32'h3e0c4d23 /* (31, 30, 2) */,
  32'h3d4ca49b /* (27, 30, 2) */,
  32'h3d1214c5 /* (23, 30, 2) */,
  32'h3d246fbd /* (19, 30, 2) */,
  32'h3d1dadb9 /* (15, 30, 2) */,
  32'h3d18e0f8 /* (11, 30, 2) */,
  32'h3d1dd271 /* (7, 30, 2) */,
  32'h3da3af74 /* (3, 30, 2) */,
  32'h3d3543e4 /* (31, 26, 2) */,
  32'h3d18df8d /* (27, 26, 2) */,
  32'h3d1e19af /* (23, 26, 2) */,
  32'h3d4ce87b /* (19, 26, 2) */,
  32'h3d4bfe66 /* (15, 26, 2) */,
  32'h3d343ccb /* (11, 26, 2) */,
  32'h3d14b9d3 /* (7, 26, 2) */,
  32'h3d271e8d /* (3, 26, 2) */,
  32'h3d12ac07 /* (31, 22, 2) */,
  32'h3d1f9f49 /* (27, 22, 2) */,
  32'h3d56480e /* (23, 22, 2) */,
  32'h3da2895a /* (19, 22, 2) */,
  32'h3daa3ec9 /* (15, 22, 2) */,
  32'h3d85a0b3 /* (11, 22, 2) */,
  32'h3d3346c6 /* (7, 22, 2) */,
  32'h3d162b76 /* (3, 22, 2) */,
  32'h3d217487 /* (31, 18, 2) */,
  32'h3d40d8bf /* (27, 18, 2) */,
  32'h3d94a37c /* (23, 18, 2) */,
  32'h3dfd653f /* (19, 18, 2) */,
  32'h3e0adb0d /* (15, 18, 2) */,
  32'h3dc55f41 /* (11, 18, 2) */,
  32'h3d6820b1 /* (7, 18, 2) */,
  32'h3d2b1735 /* (3, 18, 2) */,
  32'h3d217487 /* (31, 14, 2) */,
  32'h3d40d8bf /* (27, 14, 2) */,
  32'h3d94a37c /* (23, 14, 2) */,
  32'h3dfd653f /* (19, 14, 2) */,
  32'h3e0adb0d /* (15, 14, 2) */,
  32'h3dc55f41 /* (11, 14, 2) */,
  32'h3d6820b1 /* (7, 14, 2) */,
  32'h3d2b1735 /* (3, 14, 2) */,
  32'h3d12ac07 /* (31, 10, 2) */,
  32'h3d1f9f49 /* (27, 10, 2) */,
  32'h3d56480e /* (23, 10, 2) */,
  32'h3da2895a /* (19, 10, 2) */,
  32'h3daa3ec9 /* (15, 10, 2) */,
  32'h3d85a0b3 /* (11, 10, 2) */,
  32'h3d3346c6 /* (7, 10, 2) */,
  32'h3d162b76 /* (3, 10, 2) */,
  32'h3d3543e4 /* (31, 6, 2) */,
  32'h3d18df8d /* (27, 6, 2) */,
  32'h3d1e19af /* (23, 6, 2) */,
  32'h3d4ce87b /* (19, 6, 2) */,
  32'h3d4bfe66 /* (15, 6, 2) */,
  32'h3d343ccb /* (11, 6, 2) */,
  32'h3d14b9d3 /* (7, 6, 2) */,
  32'h3d271e8d /* (3, 6, 2) */,
  32'h3e0c4d23 /* (31, 2, 2) */,
  32'h3d4ca49b /* (27, 2, 2) */,
  32'h3d1214c5 /* (23, 2, 2) */,
  32'h3d246fbd /* (19, 2, 2) */,
  32'h3d1dadb9 /* (15, 2, 2) */,
  32'h3d18e0f8 /* (11, 2, 2) */,
  32'h3d1dd271 /* (7, 2, 2) */,
  32'h3da3af74 /* (3, 2, 2) */,
  32'h3dda3fd8 /* (30, 30, 30) */,
  32'h3d2f2a11 /* (26, 30, 30) */,
  32'h3d13e191 /* (22, 30, 30) */,
  32'h3d24f995 /* (18, 30, 30) */,
  32'h3d24f995 /* (14, 30, 30) */,
  32'h3d13e191 /* (10, 30, 30) */,
  32'h3d2f2a11 /* (6, 30, 30) */,
  32'h3dda3fd8 /* (2, 30, 30) */,
  32'h3d2f2a11 /* (30, 26, 30) */,
  32'h3d153797 /* (26, 26, 30) */,
  32'h3d27dbb1 /* (22, 26, 30) */,
  32'h3d51d4cc /* (18, 26, 30) */,
  32'h3d51d4cc /* (14, 26, 30) */,
  32'h3d27dbb1 /* (10, 26, 30) */,
  32'h3d153797 /* (6, 26, 30) */,
  32'h3d2f2a11 /* (2, 26, 30) */,
  32'h3d13e191 /* (30, 22, 30) */,
  32'h3d27dbb1 /* (26, 22, 30) */,
  32'h3d6eb6e0 /* (22, 22, 30) */,
  32'h3dab075b /* (18, 22, 30) */,
  32'h3dab075b /* (14, 22, 30) */,
  32'h3d6eb6e0 /* (10, 22, 30) */,
  32'h3d27dbb1 /* (6, 22, 30) */,
  32'h3d13e191 /* (2, 22, 30) */,
  32'h3d24f995 /* (30, 18, 30) */,
  32'h3d51d4cc /* (26, 18, 30) */,
  32'h3dab075b /* (22, 18, 30) */,
  32'h3e08838c /* (18, 18, 30) */,
  32'h3e08838c /* (14, 18, 30) */,
  32'h3dab075b /* (10, 18, 30) */,
  32'h3d51d4cc /* (6, 18, 30) */,
  32'h3d24f995 /* (2, 18, 30) */,
  32'h3d24f995 /* (30, 14, 30) */,
  32'h3d51d4cc /* (26, 14, 30) */,
  32'h3dab075b /* (22, 14, 30) */,
  32'h3e08838c /* (18, 14, 30) */,
  32'h3e08838c /* (14, 14, 30) */,
  32'h3dab075b /* (10, 14, 30) */,
  32'h3d51d4cc /* (6, 14, 30) */,
  32'h3d24f995 /* (2, 14, 30) */,
  32'h3d13e191 /* (30, 10, 30) */,
  32'h3d27dbb1 /* (26, 10, 30) */,
  32'h3d6eb6e0 /* (22, 10, 30) */,
  32'h3dab075b /* (18, 10, 30) */,
  32'h3dab075b /* (14, 10, 30) */,
  32'h3d6eb6e0 /* (10, 10, 30) */,
  32'h3d27dbb1 /* (6, 10, 30) */,
  32'h3d13e191 /* (2, 10, 30) */,
  32'h3d2f2a11 /* (30, 6, 30) */,
  32'h3d153797 /* (26, 6, 30) */,
  32'h3d27dbb1 /* (22, 6, 30) */,
  32'h3d51d4cc /* (18, 6, 30) */,
  32'h3d51d4cc /* (14, 6, 30) */,
  32'h3d27dbb1 /* (10, 6, 30) */,
  32'h3d153797 /* (6, 6, 30) */,
  32'h3d2f2a11 /* (2, 6, 30) */,
  32'h3dda3fd8 /* (30, 2, 30) */,
  32'h3d2f2a11 /* (26, 2, 30) */,
  32'h3d13e191 /* (22, 2, 30) */,
  32'h3d24f995 /* (18, 2, 30) */,
  32'h3d24f995 /* (14, 2, 30) */,
  32'h3d13e191 /* (10, 2, 30) */,
  32'h3d2f2a11 /* (6, 2, 30) */,
  32'h3dda3fd8 /* (2, 2, 30) */,
  32'h3d2f2a11 /* (30, 30, 26) */,
  32'h3d153797 /* (26, 30, 26) */,
  32'h3d27dbb1 /* (22, 30, 26) */,
  32'h3d51d4cc /* (18, 30, 26) */,
  32'h3d51d4cc /* (14, 30, 26) */,
  32'h3d27dbb1 /* (10, 30, 26) */,
  32'h3d153797 /* (6, 30, 26) */,
  32'h3d2f2a11 /* (2, 30, 26) */,
  32'h3d153797 /* (30, 26, 26) */,
  32'h3d1a814a /* (26, 26, 26) */,
  32'h3d49097c /* (22, 26, 26) */,
  32'h3d87f0f8 /* (18, 26, 26) */,
  32'h3d87f0f8 /* (14, 26, 26) */,
  32'h3d49097c /* (10, 26, 26) */,
  32'h3d1a814a /* (6, 26, 26) */,
  32'h3d153797 /* (2, 26, 26) */,
  32'h3d27dbb1 /* (30, 22, 26) */,
  32'h3d49097c /* (26, 22, 26) */,
  32'h3d97cf64 /* (22, 22, 26) */,
  32'h3de365d7 /* (18, 22, 26) */,
  32'h3de365d7 /* (14, 22, 26) */,
  32'h3d97cf64 /* (10, 22, 26) */,
  32'h3d49097c /* (6, 22, 26) */,
  32'h3d27dbb1 /* (2, 22, 26) */,
  32'h3d51d4cc /* (30, 18, 26) */,
  32'h3d87f0f8 /* (26, 18, 26) */,
  32'h3de365d7 /* (22, 18, 26) */,
  32'h3e39d98f /* (18, 18, 26) */,
  32'h3e39d98f /* (14, 18, 26) */,
  32'h3de365d7 /* (10, 18, 26) */,
  32'h3d87f0f8 /* (6, 18, 26) */,
  32'h3d51d4cc /* (2, 18, 26) */,
  32'h3d51d4cc /* (30, 14, 26) */,
  32'h3d87f0f8 /* (26, 14, 26) */,
  32'h3de365d7 /* (22, 14, 26) */,
  32'h3e39d98f /* (18, 14, 26) */,
  32'h3e39d98f /* (14, 14, 26) */,
  32'h3de365d7 /* (10, 14, 26) */,
  32'h3d87f0f8 /* (6, 14, 26) */,
  32'h3d51d4cc /* (2, 14, 26) */,
  32'h3d27dbb1 /* (30, 10, 26) */,
  32'h3d49097c /* (26, 10, 26) */,
  32'h3d97cf64 /* (22, 10, 26) */,
  32'h3de365d7 /* (18, 10, 26) */,
  32'h3de365d7 /* (14, 10, 26) */,
  32'h3d97cf64 /* (10, 10, 26) */,
  32'h3d49097c /* (6, 10, 26) */,
  32'h3d27dbb1 /* (2, 10, 26) */,
  32'h3d153797 /* (30, 6, 26) */,
  32'h3d1a814a /* (26, 6, 26) */,
  32'h3d49097c /* (22, 6, 26) */,
  32'h3d87f0f8 /* (18, 6, 26) */,
  32'h3d87f0f8 /* (14, 6, 26) */,
  32'h3d49097c /* (10, 6, 26) */,
  32'h3d1a814a /* (6, 6, 26) */,
  32'h3d153797 /* (2, 6, 26) */,
  32'h3d2f2a11 /* (30, 2, 26) */,
  32'h3d153797 /* (26, 2, 26) */,
  32'h3d27dbb1 /* (22, 2, 26) */,
  32'h3d51d4cc /* (18, 2, 26) */,
  32'h3d51d4cc /* (14, 2, 26) */,
  32'h3d27dbb1 /* (10, 2, 26) */,
  32'h3d153797 /* (6, 2, 26) */,
  32'h3d2f2a11 /* (2, 2, 26) */,
  32'h3d13e191 /* (30, 30, 22) */,
  32'h3d27dbb1 /* (26, 30, 22) */,
  32'h3d6eb6e0 /* (22, 30, 22) */,
  32'h3dab075b /* (18, 30, 22) */,
  32'h3dab075b /* (14, 30, 22) */,
  32'h3d6eb6e0 /* (10, 30, 22) */,
  32'h3d27dbb1 /* (6, 30, 22) */,
  32'h3d13e191 /* (2, 30, 22) */,
  32'h3d27dbb1 /* (30, 26, 22) */,
  32'h3d49097c /* (26, 26, 22) */,
  32'h3d97cf64 /* (22, 26, 22) */,
  32'h3de365d7 /* (18, 26, 22) */,
  32'h3de365d7 /* (14, 26, 22) */,
  32'h3d97cf64 /* (10, 26, 22) */,
  32'h3d49097c /* (6, 26, 22) */,
  32'h3d27dbb1 /* (2, 26, 22) */,
  32'h3d6eb6e0 /* (30, 22, 22) */,
  32'h3d97cf64 /* (26, 22, 22) */,
  32'h3df7795b /* (22, 22, 22) */,
  32'h3e45882e /* (18, 22, 22) */,
  32'h3e45882e /* (14, 22, 22) */,
  32'h3df7795b /* (10, 22, 22) */,
  32'h3d97cf64 /* (6, 22, 22) */,
  32'h3d6eb6e0 /* (2, 22, 22) */,
  32'h3dab075b /* (30, 18, 22) */,
  32'h3de365d7 /* (26, 18, 22) */,
  32'h3e45882e /* (22, 18, 22) */,
  32'h3ea78361 /* (18, 18, 22) */,
  32'h3ea78361 /* (14, 18, 22) */,
  32'h3e45882e /* (10, 18, 22) */,
  32'h3de365d7 /* (6, 18, 22) */,
  32'h3dab075b /* (2, 18, 22) */,
  32'h3dab075b /* (30, 14, 22) */,
  32'h3de365d7 /* (26, 14, 22) */,
  32'h3e45882e /* (22, 14, 22) */,
  32'h3ea78361 /* (18, 14, 22) */,
  32'h3ea78361 /* (14, 14, 22) */,
  32'h3e45882e /* (10, 14, 22) */,
  32'h3de365d7 /* (6, 14, 22) */,
  32'h3dab075b /* (2, 14, 22) */,
  32'h3d6eb6e0 /* (30, 10, 22) */,
  32'h3d97cf64 /* (26, 10, 22) */,
  32'h3df7795b /* (22, 10, 22) */,
  32'h3e45882e /* (18, 10, 22) */,
  32'h3e45882e /* (14, 10, 22) */,
  32'h3df7795b /* (10, 10, 22) */,
  32'h3d97cf64 /* (6, 10, 22) */,
  32'h3d6eb6e0 /* (2, 10, 22) */,
  32'h3d27dbb1 /* (30, 6, 22) */,
  32'h3d49097c /* (26, 6, 22) */,
  32'h3d97cf64 /* (22, 6, 22) */,
  32'h3de365d7 /* (18, 6, 22) */,
  32'h3de365d7 /* (14, 6, 22) */,
  32'h3d97cf64 /* (10, 6, 22) */,
  32'h3d49097c /* (6, 6, 22) */,
  32'h3d27dbb1 /* (2, 6, 22) */,
  32'h3d13e191 /* (30, 2, 22) */,
  32'h3d27dbb1 /* (26, 2, 22) */,
  32'h3d6eb6e0 /* (22, 2, 22) */,
  32'h3dab075b /* (18, 2, 22) */,
  32'h3dab075b /* (14, 2, 22) */,
  32'h3d6eb6e0 /* (10, 2, 22) */,
  32'h3d27dbb1 /* (6, 2, 22) */,
  32'h3d13e191 /* (2, 2, 22) */,
  32'h3d24f995 /* (30, 30, 18) */,
  32'h3d51d4cc /* (26, 30, 18) */,
  32'h3dab075b /* (22, 30, 18) */,
  32'h3e08838c /* (18, 30, 18) */,
  32'h3e08838c /* (14, 30, 18) */,
  32'h3dab075b /* (10, 30, 18) */,
  32'h3d51d4cc /* (6, 30, 18) */,
  32'h3d24f995 /* (2, 30, 18) */,
  32'h3d51d4cc /* (30, 26, 18) */,
  32'h3d87f0f8 /* (26, 26, 18) */,
  32'h3de365d7 /* (22, 26, 18) */,
  32'h3e39d98f /* (18, 26, 18) */,
  32'h3e39d98f /* (14, 26, 18) */,
  32'h3de365d7 /* (10, 26, 18) */,
  32'h3d87f0f8 /* (6, 26, 18) */,
  32'h3d51d4cc /* (2, 26, 18) */,
  32'h3dab075b /* (30, 22, 18) */,
  32'h3de365d7 /* (26, 22, 18) */,
  32'h3e45882e /* (22, 22, 18) */,
  32'h3ea78361 /* (18, 22, 18) */,
  32'h3ea78361 /* (14, 22, 18) */,
  32'h3e45882e /* (10, 22, 18) */,
  32'h3de365d7 /* (6, 22, 18) */,
  32'h3dab075b /* (2, 22, 18) */,
  32'h3e08838c /* (30, 18, 18) */,
  32'h3e39d98f /* (26, 18, 18) */,
  32'h3ea78361 /* (22, 18, 18) */,
  32'h3f13adcc /* (18, 18, 18) */,
  32'h3f13adcc /* (14, 18, 18) */,
  32'h3ea78361 /* (10, 18, 18) */,
  32'h3e39d98f /* (6, 18, 18) */,
  32'h3e08838c /* (2, 18, 18) */,
  32'h3e08838c /* (30, 14, 18) */,
  32'h3e39d98f /* (26, 14, 18) */,
  32'h3ea78361 /* (22, 14, 18) */,
  32'h3f13adcc /* (18, 14, 18) */,
  32'h3f13adcc /* (14, 14, 18) */,
  32'h3ea78361 /* (10, 14, 18) */,
  32'h3e39d98f /* (6, 14, 18) */,
  32'h3e08838c /* (2, 14, 18) */,
  32'h3dab075b /* (30, 10, 18) */,
  32'h3de365d7 /* (26, 10, 18) */,
  32'h3e45882e /* (22, 10, 18) */,
  32'h3ea78361 /* (18, 10, 18) */,
  32'h3ea78361 /* (14, 10, 18) */,
  32'h3e45882e /* (10, 10, 18) */,
  32'h3de365d7 /* (6, 10, 18) */,
  32'h3dab075b /* (2, 10, 18) */,
  32'h3d51d4cc /* (30, 6, 18) */,
  32'h3d87f0f8 /* (26, 6, 18) */,
  32'h3de365d7 /* (22, 6, 18) */,
  32'h3e39d98f /* (18, 6, 18) */,
  32'h3e39d98f /* (14, 6, 18) */,
  32'h3de365d7 /* (10, 6, 18) */,
  32'h3d87f0f8 /* (6, 6, 18) */,
  32'h3d51d4cc /* (2, 6, 18) */,
  32'h3d24f995 /* (30, 2, 18) */,
  32'h3d51d4cc /* (26, 2, 18) */,
  32'h3dab075b /* (22, 2, 18) */,
  32'h3e08838c /* (18, 2, 18) */,
  32'h3e08838c /* (14, 2, 18) */,
  32'h3dab075b /* (10, 2, 18) */,
  32'h3d51d4cc /* (6, 2, 18) */,
  32'h3d24f995 /* (2, 2, 18) */,
  32'h3d24f995 /* (30, 30, 14) */,
  32'h3d51d4cc /* (26, 30, 14) */,
  32'h3dab075b /* (22, 30, 14) */,
  32'h3e08838c /* (18, 30, 14) */,
  32'h3e08838c /* (14, 30, 14) */,
  32'h3dab075b /* (10, 30, 14) */,
  32'h3d51d4cc /* (6, 30, 14) */,
  32'h3d24f995 /* (2, 30, 14) */,
  32'h3d51d4cc /* (30, 26, 14) */,
  32'h3d87f0f8 /* (26, 26, 14) */,
  32'h3de365d7 /* (22, 26, 14) */,
  32'h3e39d98f /* (18, 26, 14) */,
  32'h3e39d98f /* (14, 26, 14) */,
  32'h3de365d7 /* (10, 26, 14) */,
  32'h3d87f0f8 /* (6, 26, 14) */,
  32'h3d51d4cc /* (2, 26, 14) */,
  32'h3dab075b /* (30, 22, 14) */,
  32'h3de365d7 /* (26, 22, 14) */,
  32'h3e45882e /* (22, 22, 14) */,
  32'h3ea78361 /* (18, 22, 14) */,
  32'h3ea78361 /* (14, 22, 14) */,
  32'h3e45882e /* (10, 22, 14) */,
  32'h3de365d7 /* (6, 22, 14) */,
  32'h3dab075b /* (2, 22, 14) */,
  32'h3e08838c /* (30, 18, 14) */,
  32'h3e39d98f /* (26, 18, 14) */,
  32'h3ea78361 /* (22, 18, 14) */,
  32'h3f13adcc /* (18, 18, 14) */,
  32'h3f13adcc /* (14, 18, 14) */,
  32'h3ea78361 /* (10, 18, 14) */,
  32'h3e39d98f /* (6, 18, 14) */,
  32'h3e08838c /* (2, 18, 14) */,
  32'h3e08838c /* (30, 14, 14) */,
  32'h3e39d98f /* (26, 14, 14) */,
  32'h3ea78361 /* (22, 14, 14) */,
  32'h3f13adcc /* (18, 14, 14) */,
  32'h3f13adcc /* (14, 14, 14) */,
  32'h3ea78361 /* (10, 14, 14) */,
  32'h3e39d98f /* (6, 14, 14) */,
  32'h3e08838c /* (2, 14, 14) */,
  32'h3dab075b /* (30, 10, 14) */,
  32'h3de365d7 /* (26, 10, 14) */,
  32'h3e45882e /* (22, 10, 14) */,
  32'h3ea78361 /* (18, 10, 14) */,
  32'h3ea78361 /* (14, 10, 14) */,
  32'h3e45882e /* (10, 10, 14) */,
  32'h3de365d7 /* (6, 10, 14) */,
  32'h3dab075b /* (2, 10, 14) */,
  32'h3d51d4cc /* (30, 6, 14) */,
  32'h3d87f0f8 /* (26, 6, 14) */,
  32'h3de365d7 /* (22, 6, 14) */,
  32'h3e39d98f /* (18, 6, 14) */,
  32'h3e39d98f /* (14, 6, 14) */,
  32'h3de365d7 /* (10, 6, 14) */,
  32'h3d87f0f8 /* (6, 6, 14) */,
  32'h3d51d4cc /* (2, 6, 14) */,
  32'h3d24f995 /* (30, 2, 14) */,
  32'h3d51d4cc /* (26, 2, 14) */,
  32'h3dab075b /* (22, 2, 14) */,
  32'h3e08838c /* (18, 2, 14) */,
  32'h3e08838c /* (14, 2, 14) */,
  32'h3dab075b /* (10, 2, 14) */,
  32'h3d51d4cc /* (6, 2, 14) */,
  32'h3d24f995 /* (2, 2, 14) */,
  32'h3d13e191 /* (30, 30, 10) */,
  32'h3d27dbb1 /* (26, 30, 10) */,
  32'h3d6eb6e0 /* (22, 30, 10) */,
  32'h3dab075b /* (18, 30, 10) */,
  32'h3dab075b /* (14, 30, 10) */,
  32'h3d6eb6e0 /* (10, 30, 10) */,
  32'h3d27dbb1 /* (6, 30, 10) */,
  32'h3d13e191 /* (2, 30, 10) */,
  32'h3d27dbb1 /* (30, 26, 10) */,
  32'h3d49097c /* (26, 26, 10) */,
  32'h3d97cf64 /* (22, 26, 10) */,
  32'h3de365d7 /* (18, 26, 10) */,
  32'h3de365d7 /* (14, 26, 10) */,
  32'h3d97cf64 /* (10, 26, 10) */,
  32'h3d49097c /* (6, 26, 10) */,
  32'h3d27dbb1 /* (2, 26, 10) */,
  32'h3d6eb6e0 /* (30, 22, 10) */,
  32'h3d97cf64 /* (26, 22, 10) */,
  32'h3df7795b /* (22, 22, 10) */,
  32'h3e45882e /* (18, 22, 10) */,
  32'h3e45882e /* (14, 22, 10) */,
  32'h3df7795b /* (10, 22, 10) */,
  32'h3d97cf64 /* (6, 22, 10) */,
  32'h3d6eb6e0 /* (2, 22, 10) */,
  32'h3dab075b /* (30, 18, 10) */,
  32'h3de365d7 /* (26, 18, 10) */,
  32'h3e45882e /* (22, 18, 10) */,
  32'h3ea78361 /* (18, 18, 10) */,
  32'h3ea78361 /* (14, 18, 10) */,
  32'h3e45882e /* (10, 18, 10) */,
  32'h3de365d7 /* (6, 18, 10) */,
  32'h3dab075b /* (2, 18, 10) */,
  32'h3dab075b /* (30, 14, 10) */,
  32'h3de365d7 /* (26, 14, 10) */,
  32'h3e45882e /* (22, 14, 10) */,
  32'h3ea78361 /* (18, 14, 10) */,
  32'h3ea78361 /* (14, 14, 10) */,
  32'h3e45882e /* (10, 14, 10) */,
  32'h3de365d7 /* (6, 14, 10) */,
  32'h3dab075b /* (2, 14, 10) */,
  32'h3d6eb6e0 /* (30, 10, 10) */,
  32'h3d97cf64 /* (26, 10, 10) */,
  32'h3df7795b /* (22, 10, 10) */,
  32'h3e45882e /* (18, 10, 10) */,
  32'h3e45882e /* (14, 10, 10) */,
  32'h3df7795b /* (10, 10, 10) */,
  32'h3d97cf64 /* (6, 10, 10) */,
  32'h3d6eb6e0 /* (2, 10, 10) */,
  32'h3d27dbb1 /* (30, 6, 10) */,
  32'h3d49097c /* (26, 6, 10) */,
  32'h3d97cf64 /* (22, 6, 10) */,
  32'h3de365d7 /* (18, 6, 10) */,
  32'h3de365d7 /* (14, 6, 10) */,
  32'h3d97cf64 /* (10, 6, 10) */,
  32'h3d49097c /* (6, 6, 10) */,
  32'h3d27dbb1 /* (2, 6, 10) */,
  32'h3d13e191 /* (30, 2, 10) */,
  32'h3d27dbb1 /* (26, 2, 10) */,
  32'h3d6eb6e0 /* (22, 2, 10) */,
  32'h3dab075b /* (18, 2, 10) */,
  32'h3dab075b /* (14, 2, 10) */,
  32'h3d6eb6e0 /* (10, 2, 10) */,
  32'h3d27dbb1 /* (6, 2, 10) */,
  32'h3d13e191 /* (2, 2, 10) */,
  32'h3d2f2a11 /* (30, 30, 6) */,
  32'h3d153797 /* (26, 30, 6) */,
  32'h3d27dbb1 /* (22, 30, 6) */,
  32'h3d51d4cc /* (18, 30, 6) */,
  32'h3d51d4cc /* (14, 30, 6) */,
  32'h3d27dbb1 /* (10, 30, 6) */,
  32'h3d153797 /* (6, 30, 6) */,
  32'h3d2f2a11 /* (2, 30, 6) */,
  32'h3d153797 /* (30, 26, 6) */,
  32'h3d1a814a /* (26, 26, 6) */,
  32'h3d49097c /* (22, 26, 6) */,
  32'h3d87f0f8 /* (18, 26, 6) */,
  32'h3d87f0f8 /* (14, 26, 6) */,
  32'h3d49097c /* (10, 26, 6) */,
  32'h3d1a814a /* (6, 26, 6) */,
  32'h3d153797 /* (2, 26, 6) */,
  32'h3d27dbb1 /* (30, 22, 6) */,
  32'h3d49097c /* (26, 22, 6) */,
  32'h3d97cf64 /* (22, 22, 6) */,
  32'h3de365d7 /* (18, 22, 6) */,
  32'h3de365d7 /* (14, 22, 6) */,
  32'h3d97cf64 /* (10, 22, 6) */,
  32'h3d49097c /* (6, 22, 6) */,
  32'h3d27dbb1 /* (2, 22, 6) */,
  32'h3d51d4cc /* (30, 18, 6) */,
  32'h3d87f0f8 /* (26, 18, 6) */,
  32'h3de365d7 /* (22, 18, 6) */,
  32'h3e39d98f /* (18, 18, 6) */,
  32'h3e39d98f /* (14, 18, 6) */,
  32'h3de365d7 /* (10, 18, 6) */,
  32'h3d87f0f8 /* (6, 18, 6) */,
  32'h3d51d4cc /* (2, 18, 6) */,
  32'h3d51d4cc /* (30, 14, 6) */,
  32'h3d87f0f8 /* (26, 14, 6) */,
  32'h3de365d7 /* (22, 14, 6) */,
  32'h3e39d98f /* (18, 14, 6) */,
  32'h3e39d98f /* (14, 14, 6) */,
  32'h3de365d7 /* (10, 14, 6) */,
  32'h3d87f0f8 /* (6, 14, 6) */,
  32'h3d51d4cc /* (2, 14, 6) */,
  32'h3d27dbb1 /* (30, 10, 6) */,
  32'h3d49097c /* (26, 10, 6) */,
  32'h3d97cf64 /* (22, 10, 6) */,
  32'h3de365d7 /* (18, 10, 6) */,
  32'h3de365d7 /* (14, 10, 6) */,
  32'h3d97cf64 /* (10, 10, 6) */,
  32'h3d49097c /* (6, 10, 6) */,
  32'h3d27dbb1 /* (2, 10, 6) */,
  32'h3d153797 /* (30, 6, 6) */,
  32'h3d1a814a /* (26, 6, 6) */,
  32'h3d49097c /* (22, 6, 6) */,
  32'h3d87f0f8 /* (18, 6, 6) */,
  32'h3d87f0f8 /* (14, 6, 6) */,
  32'h3d49097c /* (10, 6, 6) */,
  32'h3d1a814a /* (6, 6, 6) */,
  32'h3d153797 /* (2, 6, 6) */,
  32'h3d2f2a11 /* (30, 2, 6) */,
  32'h3d153797 /* (26, 2, 6) */,
  32'h3d27dbb1 /* (22, 2, 6) */,
  32'h3d51d4cc /* (18, 2, 6) */,
  32'h3d51d4cc /* (14, 2, 6) */,
  32'h3d27dbb1 /* (10, 2, 6) */,
  32'h3d153797 /* (6, 2, 6) */,
  32'h3d2f2a11 /* (2, 2, 6) */,
  32'h3dda3fd8 /* (30, 30, 2) */,
  32'h3d2f2a11 /* (26, 30, 2) */,
  32'h3d13e191 /* (22, 30, 2) */,
  32'h3d24f995 /* (18, 30, 2) */,
  32'h3d24f995 /* (14, 30, 2) */,
  32'h3d13e191 /* (10, 30, 2) */,
  32'h3d2f2a11 /* (6, 30, 2) */,
  32'h3dda3fd8 /* (2, 30, 2) */,
  32'h3d2f2a11 /* (30, 26, 2) */,
  32'h3d153797 /* (26, 26, 2) */,
  32'h3d27dbb1 /* (22, 26, 2) */,
  32'h3d51d4cc /* (18, 26, 2) */,
  32'h3d51d4cc /* (14, 26, 2) */,
  32'h3d27dbb1 /* (10, 26, 2) */,
  32'h3d153797 /* (6, 26, 2) */,
  32'h3d2f2a11 /* (2, 26, 2) */,
  32'h3d13e191 /* (30, 22, 2) */,
  32'h3d27dbb1 /* (26, 22, 2) */,
  32'h3d6eb6e0 /* (22, 22, 2) */,
  32'h3dab075b /* (18, 22, 2) */,
  32'h3dab075b /* (14, 22, 2) */,
  32'h3d6eb6e0 /* (10, 22, 2) */,
  32'h3d27dbb1 /* (6, 22, 2) */,
  32'h3d13e191 /* (2, 22, 2) */,
  32'h3d24f995 /* (30, 18, 2) */,
  32'h3d51d4cc /* (26, 18, 2) */,
  32'h3dab075b /* (22, 18, 2) */,
  32'h3e08838c /* (18, 18, 2) */,
  32'h3e08838c /* (14, 18, 2) */,
  32'h3dab075b /* (10, 18, 2) */,
  32'h3d51d4cc /* (6, 18, 2) */,
  32'h3d24f995 /* (2, 18, 2) */,
  32'h3d24f995 /* (30, 14, 2) */,
  32'h3d51d4cc /* (26, 14, 2) */,
  32'h3dab075b /* (22, 14, 2) */,
  32'h3e08838c /* (18, 14, 2) */,
  32'h3e08838c /* (14, 14, 2) */,
  32'h3dab075b /* (10, 14, 2) */,
  32'h3d51d4cc /* (6, 14, 2) */,
  32'h3d24f995 /* (2, 14, 2) */,
  32'h3d13e191 /* (30, 10, 2) */,
  32'h3d27dbb1 /* (26, 10, 2) */,
  32'h3d6eb6e0 /* (22, 10, 2) */,
  32'h3dab075b /* (18, 10, 2) */,
  32'h3dab075b /* (14, 10, 2) */,
  32'h3d6eb6e0 /* (10, 10, 2) */,
  32'h3d27dbb1 /* (6, 10, 2) */,
  32'h3d13e191 /* (2, 10, 2) */,
  32'h3d2f2a11 /* (30, 6, 2) */,
  32'h3d153797 /* (26, 6, 2) */,
  32'h3d27dbb1 /* (22, 6, 2) */,
  32'h3d51d4cc /* (18, 6, 2) */,
  32'h3d51d4cc /* (14, 6, 2) */,
  32'h3d27dbb1 /* (10, 6, 2) */,
  32'h3d153797 /* (6, 6, 2) */,
  32'h3d2f2a11 /* (2, 6, 2) */,
  32'h3dda3fd8 /* (30, 2, 2) */,
  32'h3d2f2a11 /* (26, 2, 2) */,
  32'h3d13e191 /* (22, 2, 2) */,
  32'h3d24f995 /* (18, 2, 2) */,
  32'h3d24f995 /* (14, 2, 2) */,
  32'h3d13e191 /* (10, 2, 2) */,
  32'h3d2f2a11 /* (6, 2, 2) */,
  32'h3dda3fd8 /* (2, 2, 2) */,
  32'h3da3af74 /* (29, 30, 30) */,
  32'h3d1dd271 /* (25, 30, 30) */,
  32'h3d18e0f8 /* (21, 30, 30) */,
  32'h3d1dadb9 /* (17, 30, 30) */,
  32'h3d246fbd /* (13, 30, 30) */,
  32'h3d1214c5 /* (9, 30, 30) */,
  32'h3d4ca49b /* (5, 30, 30) */,
  32'h3e0c4d23 /* (1, 30, 30) */,
  32'h3d271e8d /* (29, 26, 30) */,
  32'h3d14b9d3 /* (25, 26, 30) */,
  32'h3d343ccb /* (21, 26, 30) */,
  32'h3d4bfe66 /* (17, 26, 30) */,
  32'h3d4ce87b /* (13, 26, 30) */,
  32'h3d1e19af /* (9, 26, 30) */,
  32'h3d18df8d /* (5, 26, 30) */,
  32'h3d3543e4 /* (1, 26, 30) */,
  32'h3d162b76 /* (29, 22, 30) */,
  32'h3d3346c6 /* (25, 22, 30) */,
  32'h3d85a0b3 /* (21, 22, 30) */,
  32'h3daa3ec9 /* (17, 22, 30) */,
  32'h3da2895a /* (13, 22, 30) */,
  32'h3d56480e /* (9, 22, 30) */,
  32'h3d1f9f49 /* (5, 22, 30) */,
  32'h3d12ac07 /* (1, 22, 30) */,
  32'h3d2b1735 /* (29, 18, 30) */,
  32'h3d6820b1 /* (25, 18, 30) */,
  32'h3dc55f41 /* (21, 18, 30) */,
  32'h3e0adb0d /* (17, 18, 30) */,
  32'h3dfd653f /* (13, 18, 30) */,
  32'h3d94a37c /* (9, 18, 30) */,
  32'h3d40d8bf /* (5, 18, 30) */,
  32'h3d217487 /* (1, 18, 30) */,
  32'h3d2b1735 /* (29, 14, 30) */,
  32'h3d6820b1 /* (25, 14, 30) */,
  32'h3dc55f41 /* (21, 14, 30) */,
  32'h3e0adb0d /* (17, 14, 30) */,
  32'h3dfd653f /* (13, 14, 30) */,
  32'h3d94a37c /* (9, 14, 30) */,
  32'h3d40d8bf /* (5, 14, 30) */,
  32'h3d217487 /* (1, 14, 30) */,
  32'h3d162b76 /* (29, 10, 30) */,
  32'h3d3346c6 /* (25, 10, 30) */,
  32'h3d85a0b3 /* (21, 10, 30) */,
  32'h3daa3ec9 /* (17, 10, 30) */,
  32'h3da2895a /* (13, 10, 30) */,
  32'h3d56480e /* (9, 10, 30) */,
  32'h3d1f9f49 /* (5, 10, 30) */,
  32'h3d12ac07 /* (1, 10, 30) */,
  32'h3d271e8d /* (29, 6, 30) */,
  32'h3d14b9d3 /* (25, 6, 30) */,
  32'h3d343ccb /* (21, 6, 30) */,
  32'h3d4bfe66 /* (17, 6, 30) */,
  32'h3d4ce87b /* (13, 6, 30) */,
  32'h3d1e19af /* (9, 6, 30) */,
  32'h3d18df8d /* (5, 6, 30) */,
  32'h3d3543e4 /* (1, 6, 30) */,
  32'h3da3af74 /* (29, 2, 30) */,
  32'h3d1dd271 /* (25, 2, 30) */,
  32'h3d18e0f8 /* (21, 2, 30) */,
  32'h3d1dadb9 /* (17, 2, 30) */,
  32'h3d246fbd /* (13, 2, 30) */,
  32'h3d1214c5 /* (9, 2, 30) */,
  32'h3d4ca49b /* (5, 2, 30) */,
  32'h3e0c4d23 /* (1, 2, 30) */,
  32'h3d271e8d /* (29, 30, 26) */,
  32'h3d14b9d3 /* (25, 30, 26) */,
  32'h3d343ccb /* (21, 30, 26) */,
  32'h3d4bfe66 /* (17, 30, 26) */,
  32'h3d4ce87b /* (13, 30, 26) */,
  32'h3d1e19af /* (9, 30, 26) */,
  32'h3d18df8d /* (5, 30, 26) */,
  32'h3d3543e4 /* (1, 30, 26) */,
  32'h3d14c14d /* (29, 26, 26) */,
  32'h3d20f672 /* (25, 26, 26) */,
  32'h3d5d3b5c /* (21, 26, 26) */,
  32'h3d85e8bf /* (17, 26, 26) */,
  32'h3d82bc35 /* (13, 26, 26) */,
  32'h3d37f9d0 /* (9, 26, 26) */,
  32'h3d16bb8b /* (5, 26, 26) */,
  32'h3d15cc97 /* (1, 26, 26) */,
  32'h3d2c3293 /* (29, 22, 26) */,
  32'h3d5a2934 /* (25, 22, 26) */,
  32'h3dac23aa /* (21, 22, 26) */,
  32'h3de44bb3 /* (17, 22, 26) */,
  32'h3dd610ea /* (13, 22, 26) */,
  32'h3d866682 /* (9, 22, 26) */,
  32'h3d3c300c /* (5, 22, 26) */,
  32'h3d2567ce /* (1, 22, 26) */,
  32'h3d5a5169 /* (29, 18, 26) */,
  32'h3d975464 /* (25, 18, 26) */,
  32'h3e040b60 /* (21, 18, 26) */,
  32'h3e3e01e0 /* (17, 18, 26) */,
  32'h3e2b8c37 /* (13, 18, 26) */,
  32'h3dc45939 /* (9, 18, 26) */,
  32'h3d786cd6 /* (5, 18, 26) */,
  32'h3d4cf093 /* (1, 18, 26) */,
  32'h3d5a5169 /* (29, 14, 26) */,
  32'h3d975464 /* (25, 14, 26) */,
  32'h3e040b60 /* (21, 14, 26) */,
  32'h3e3e01e0 /* (17, 14, 26) */,
  32'h3e2b8c37 /* (13, 14, 26) */,
  32'h3dc45939 /* (9, 14, 26) */,
  32'h3d786cd6 /* (5, 14, 26) */,
  32'h3d4cf093 /* (1, 14, 26) */,
  32'h3d2c3293 /* (29, 10, 26) */,
  32'h3d5a2934 /* (25, 10, 26) */,
  32'h3dac23aa /* (21, 10, 26) */,
  32'h3de44bb3 /* (17, 10, 26) */,
  32'h3dd610ea /* (13, 10, 26) */,
  32'h3d866682 /* (9, 10, 26) */,
  32'h3d3c300c /* (5, 10, 26) */,
  32'h3d2567ce /* (1, 10, 26) */,
  32'h3d14c14d /* (29, 6, 26) */,
  32'h3d20f672 /* (25, 6, 26) */,
  32'h3d5d3b5c /* (21, 6, 26) */,
  32'h3d85e8bf /* (17, 6, 26) */,
  32'h3d82bc35 /* (13, 6, 26) */,
  32'h3d37f9d0 /* (9, 6, 26) */,
  32'h3d16bb8b /* (5, 6, 26) */,
  32'h3d15cc97 /* (1, 6, 26) */,
  32'h3d271e8d /* (29, 2, 26) */,
  32'h3d14b9d3 /* (25, 2, 26) */,
  32'h3d343ccb /* (21, 2, 26) */,
  32'h3d4bfe66 /* (17, 2, 26) */,
  32'h3d4ce87b /* (13, 2, 26) */,
  32'h3d1e19af /* (9, 2, 26) */,
  32'h3d18df8d /* (5, 2, 26) */,
  32'h3d3543e4 /* (1, 2, 26) */,
  32'h3d162b76 /* (29, 30, 22) */,
  32'h3d3346c6 /* (25, 30, 22) */,
  32'h3d85a0b3 /* (21, 30, 22) */,
  32'h3daa3ec9 /* (17, 30, 22) */,
  32'h3da2895a /* (13, 30, 22) */,
  32'h3d56480e /* (9, 30, 22) */,
  32'h3d1f9f49 /* (5, 30, 22) */,
  32'h3d12ac07 /* (1, 30, 22) */,
  32'h3d2c3293 /* (29, 26, 22) */,
  32'h3d5a2934 /* (25, 26, 22) */,
  32'h3dac23aa /* (21, 26, 22) */,
  32'h3de44bb3 /* (17, 26, 22) */,
  32'h3dd610ea /* (13, 26, 22) */,
  32'h3d866682 /* (9, 26, 22) */,
  32'h3d3c300c /* (5, 26, 22) */,
  32'h3d2567ce /* (1, 26, 22) */,
  32'h3d77904c /* (29, 22, 22) */,
  32'h3da7f0fb /* (25, 22, 22) */,
  32'h3e0ecbcd /* (21, 22, 22) */,
  32'h3e48eba4 /* (17, 22, 22) */,
  32'h3e37540b /* (13, 22, 22) */,
  32'h3dd7137d /* (9, 22, 22) */,
  32'h3d8b85a2 /* (5, 22, 22) */,
  32'h3d699f13 /* (1, 22, 22) */,
  32'h3db2bcb9 /* (29, 18, 22) */,
  32'h3dff6ab3 /* (25, 18, 22) */,
  32'h3e67a191 /* (21, 18, 22) */,
  32'h3eacaf9b /* (17, 18, 22) */,
  32'h3e994798 /* (13, 18, 22) */,
  32'h3e28e750 /* (9, 18, 22) */,
  32'h3dce13fe /* (5, 18, 22) */,
  32'h3da6958f /* (1, 18, 22) */,
  32'h3db2bcb9 /* (29, 14, 22) */,
  32'h3dff6ab3 /* (25, 14, 22) */,
  32'h3e67a191 /* (21, 14, 22) */,
  32'h3eacaf9b /* (17, 14, 22) */,
  32'h3e994798 /* (13, 14, 22) */,
  32'h3e28e750 /* (9, 14, 22) */,
  32'h3dce13fe /* (5, 14, 22) */,
  32'h3da6958f /* (1, 14, 22) */,
  32'h3d77904c /* (29, 10, 22) */,
  32'h3da7f0fb /* (25, 10, 22) */,
  32'h3e0ecbcd /* (21, 10, 22) */,
  32'h3e48eba4 /* (17, 10, 22) */,
  32'h3e37540b /* (13, 10, 22) */,
  32'h3dd7137d /* (9, 10, 22) */,
  32'h3d8b85a2 /* (5, 10, 22) */,
  32'h3d699f13 /* (1, 10, 22) */,
  32'h3d2c3293 /* (29, 6, 22) */,
  32'h3d5a2934 /* (25, 6, 22) */,
  32'h3dac23aa /* (21, 6, 22) */,
  32'h3de44bb3 /* (17, 6, 22) */,
  32'h3dd610ea /* (13, 6, 22) */,
  32'h3d866682 /* (9, 6, 22) */,
  32'h3d3c300c /* (5, 6, 22) */,
  32'h3d2567ce /* (1, 6, 22) */,
  32'h3d162b76 /* (29, 2, 22) */,
  32'h3d3346c6 /* (25, 2, 22) */,
  32'h3d85a0b3 /* (21, 2, 22) */,
  32'h3daa3ec9 /* (17, 2, 22) */,
  32'h3da2895a /* (13, 2, 22) */,
  32'h3d56480e /* (9, 2, 22) */,
  32'h3d1f9f49 /* (5, 2, 22) */,
  32'h3d12ac07 /* (1, 2, 22) */,
  32'h3d2b1735 /* (29, 30, 18) */,
  32'h3d6820b1 /* (25, 30, 18) */,
  32'h3dc55f41 /* (21, 30, 18) */,
  32'h3e0adb0d /* (17, 30, 18) */,
  32'h3dfd653f /* (13, 30, 18) */,
  32'h3d94a37c /* (9, 30, 18) */,
  32'h3d40d8bf /* (5, 30, 18) */,
  32'h3d217487 /* (1, 30, 18) */,
  32'h3d5a5169 /* (29, 26, 18) */,
  32'h3d975464 /* (25, 26, 18) */,
  32'h3e040b60 /* (21, 26, 18) */,
  32'h3e3e01e0 /* (17, 26, 18) */,
  32'h3e2b8c37 /* (13, 26, 18) */,
  32'h3dc45939 /* (9, 26, 18) */,
  32'h3d786cd6 /* (5, 26, 18) */,
  32'h3d4cf093 /* (1, 26, 18) */,
  32'h3db2bcb9 /* (29, 22, 18) */,
  32'h3dff6ab3 /* (25, 22, 18) */,
  32'h3e67a191 /* (21, 22, 18) */,
  32'h3eacaf9b /* (17, 22, 18) */,
  32'h3e994798 /* (13, 22, 18) */,
  32'h3e28e750 /* (9, 22, 18) */,
  32'h3dce13fe /* (5, 22, 18) */,
  32'h3da6958f /* (1, 22, 18) */,
  32'h3e0f3c67 /* (29, 18, 18) */,
  32'h3e528761 /* (25, 18, 18) */,
  32'h3ec66134 /* (21, 18, 18) */,
  32'h3f19a2a7 /* (17, 18, 18) */,
  32'h3f05dc96 /* (13, 18, 18) */,
  32'h3e8dd733 /* (9, 18, 18) */,
  32'h3e27240a /* (5, 18, 18) */,
  32'h3e04a438 /* (1, 18, 18) */,
  32'h3e0f3c67 /* (29, 14, 18) */,
  32'h3e528761 /* (25, 14, 18) */,
  32'h3ec66134 /* (21, 14, 18) */,
  32'h3f19a2a7 /* (17, 14, 18) */,
  32'h3f05dc96 /* (13, 14, 18) */,
  32'h3e8dd733 /* (9, 14, 18) */,
  32'h3e27240a /* (5, 14, 18) */,
  32'h3e04a438 /* (1, 14, 18) */,
  32'h3db2bcb9 /* (29, 10, 18) */,
  32'h3dff6ab3 /* (25, 10, 18) */,
  32'h3e67a191 /* (21, 10, 18) */,
  32'h3eacaf9b /* (17, 10, 18) */,
  32'h3e994798 /* (13, 10, 18) */,
  32'h3e28e750 /* (9, 10, 18) */,
  32'h3dce13fe /* (5, 10, 18) */,
  32'h3da6958f /* (1, 10, 18) */,
  32'h3d5a5169 /* (29, 6, 18) */,
  32'h3d975464 /* (25, 6, 18) */,
  32'h3e040b60 /* (21, 6, 18) */,
  32'h3e3e01e0 /* (17, 6, 18) */,
  32'h3e2b8c37 /* (13, 6, 18) */,
  32'h3dc45939 /* (9, 6, 18) */,
  32'h3d786cd6 /* (5, 6, 18) */,
  32'h3d4cf093 /* (1, 6, 18) */,
  32'h3d2b1735 /* (29, 2, 18) */,
  32'h3d6820b1 /* (25, 2, 18) */,
  32'h3dc55f41 /* (21, 2, 18) */,
  32'h3e0adb0d /* (17, 2, 18) */,
  32'h3dfd653f /* (13, 2, 18) */,
  32'h3d94a37c /* (9, 2, 18) */,
  32'h3d40d8bf /* (5, 2, 18) */,
  32'h3d217487 /* (1, 2, 18) */,
  32'h3d2b1735 /* (29, 30, 14) */,
  32'h3d6820b1 /* (25, 30, 14) */,
  32'h3dc55f41 /* (21, 30, 14) */,
  32'h3e0adb0d /* (17, 30, 14) */,
  32'h3dfd653f /* (13, 30, 14) */,
  32'h3d94a37c /* (9, 30, 14) */,
  32'h3d40d8bf /* (5, 30, 14) */,
  32'h3d217487 /* (1, 30, 14) */,
  32'h3d5a5169 /* (29, 26, 14) */,
  32'h3d975464 /* (25, 26, 14) */,
  32'h3e040b60 /* (21, 26, 14) */,
  32'h3e3e01e0 /* (17, 26, 14) */,
  32'h3e2b8c37 /* (13, 26, 14) */,
  32'h3dc45939 /* (9, 26, 14) */,
  32'h3d786cd6 /* (5, 26, 14) */,
  32'h3d4cf093 /* (1, 26, 14) */,
  32'h3db2bcb9 /* (29, 22, 14) */,
  32'h3dff6ab3 /* (25, 22, 14) */,
  32'h3e67a191 /* (21, 22, 14) */,
  32'h3eacaf9b /* (17, 22, 14) */,
  32'h3e994798 /* (13, 22, 14) */,
  32'h3e28e750 /* (9, 22, 14) */,
  32'h3dce13fe /* (5, 22, 14) */,
  32'h3da6958f /* (1, 22, 14) */,
  32'h3e0f3c67 /* (29, 18, 14) */,
  32'h3e528761 /* (25, 18, 14) */,
  32'h3ec66134 /* (21, 18, 14) */,
  32'h3f19a2a7 /* (17, 18, 14) */,
  32'h3f05dc96 /* (13, 18, 14) */,
  32'h3e8dd733 /* (9, 18, 14) */,
  32'h3e27240a /* (5, 18, 14) */,
  32'h3e04a438 /* (1, 18, 14) */,
  32'h3e0f3c67 /* (29, 14, 14) */,
  32'h3e528761 /* (25, 14, 14) */,
  32'h3ec66134 /* (21, 14, 14) */,
  32'h3f19a2a7 /* (17, 14, 14) */,
  32'h3f05dc96 /* (13, 14, 14) */,
  32'h3e8dd733 /* (9, 14, 14) */,
  32'h3e27240a /* (5, 14, 14) */,
  32'h3e04a438 /* (1, 14, 14) */,
  32'h3db2bcb9 /* (29, 10, 14) */,
  32'h3dff6ab3 /* (25, 10, 14) */,
  32'h3e67a191 /* (21, 10, 14) */,
  32'h3eacaf9b /* (17, 10, 14) */,
  32'h3e994798 /* (13, 10, 14) */,
  32'h3e28e750 /* (9, 10, 14) */,
  32'h3dce13fe /* (5, 10, 14) */,
  32'h3da6958f /* (1, 10, 14) */,
  32'h3d5a5169 /* (29, 6, 14) */,
  32'h3d975464 /* (25, 6, 14) */,
  32'h3e040b60 /* (21, 6, 14) */,
  32'h3e3e01e0 /* (17, 6, 14) */,
  32'h3e2b8c37 /* (13, 6, 14) */,
  32'h3dc45939 /* (9, 6, 14) */,
  32'h3d786cd6 /* (5, 6, 14) */,
  32'h3d4cf093 /* (1, 6, 14) */,
  32'h3d2b1735 /* (29, 2, 14) */,
  32'h3d6820b1 /* (25, 2, 14) */,
  32'h3dc55f41 /* (21, 2, 14) */,
  32'h3e0adb0d /* (17, 2, 14) */,
  32'h3dfd653f /* (13, 2, 14) */,
  32'h3d94a37c /* (9, 2, 14) */,
  32'h3d40d8bf /* (5, 2, 14) */,
  32'h3d217487 /* (1, 2, 14) */,
  32'h3d162b76 /* (29, 30, 10) */,
  32'h3d3346c6 /* (25, 30, 10) */,
  32'h3d85a0b3 /* (21, 30, 10) */,
  32'h3daa3ec9 /* (17, 30, 10) */,
  32'h3da2895a /* (13, 30, 10) */,
  32'h3d56480e /* (9, 30, 10) */,
  32'h3d1f9f49 /* (5, 30, 10) */,
  32'h3d12ac07 /* (1, 30, 10) */,
  32'h3d2c3293 /* (29, 26, 10) */,
  32'h3d5a2934 /* (25, 26, 10) */,
  32'h3dac23aa /* (21, 26, 10) */,
  32'h3de44bb3 /* (17, 26, 10) */,
  32'h3dd610ea /* (13, 26, 10) */,
  32'h3d866682 /* (9, 26, 10) */,
  32'h3d3c300c /* (5, 26, 10) */,
  32'h3d2567ce /* (1, 26, 10) */,
  32'h3d77904c /* (29, 22, 10) */,
  32'h3da7f0fb /* (25, 22, 10) */,
  32'h3e0ecbcd /* (21, 22, 10) */,
  32'h3e48eba4 /* (17, 22, 10) */,
  32'h3e37540b /* (13, 22, 10) */,
  32'h3dd7137d /* (9, 22, 10) */,
  32'h3d8b85a2 /* (5, 22, 10) */,
  32'h3d699f13 /* (1, 22, 10) */,
  32'h3db2bcb9 /* (29, 18, 10) */,
  32'h3dff6ab3 /* (25, 18, 10) */,
  32'h3e67a191 /* (21, 18, 10) */,
  32'h3eacaf9b /* (17, 18, 10) */,
  32'h3e994798 /* (13, 18, 10) */,
  32'h3e28e750 /* (9, 18, 10) */,
  32'h3dce13fe /* (5, 18, 10) */,
  32'h3da6958f /* (1, 18, 10) */,
  32'h3db2bcb9 /* (29, 14, 10) */,
  32'h3dff6ab3 /* (25, 14, 10) */,
  32'h3e67a191 /* (21, 14, 10) */,
  32'h3eacaf9b /* (17, 14, 10) */,
  32'h3e994798 /* (13, 14, 10) */,
  32'h3e28e750 /* (9, 14, 10) */,
  32'h3dce13fe /* (5, 14, 10) */,
  32'h3da6958f /* (1, 14, 10) */,
  32'h3d77904c /* (29, 10, 10) */,
  32'h3da7f0fb /* (25, 10, 10) */,
  32'h3e0ecbcd /* (21, 10, 10) */,
  32'h3e48eba4 /* (17, 10, 10) */,
  32'h3e37540b /* (13, 10, 10) */,
  32'h3dd7137d /* (9, 10, 10) */,
  32'h3d8b85a2 /* (5, 10, 10) */,
  32'h3d699f13 /* (1, 10, 10) */,
  32'h3d2c3293 /* (29, 6, 10) */,
  32'h3d5a2934 /* (25, 6, 10) */,
  32'h3dac23aa /* (21, 6, 10) */,
  32'h3de44bb3 /* (17, 6, 10) */,
  32'h3dd610ea /* (13, 6, 10) */,
  32'h3d866682 /* (9, 6, 10) */,
  32'h3d3c300c /* (5, 6, 10) */,
  32'h3d2567ce /* (1, 6, 10) */,
  32'h3d162b76 /* (29, 2, 10) */,
  32'h3d3346c6 /* (25, 2, 10) */,
  32'h3d85a0b3 /* (21, 2, 10) */,
  32'h3daa3ec9 /* (17, 2, 10) */,
  32'h3da2895a /* (13, 2, 10) */,
  32'h3d56480e /* (9, 2, 10) */,
  32'h3d1f9f49 /* (5, 2, 10) */,
  32'h3d12ac07 /* (1, 2, 10) */,
  32'h3d271e8d /* (29, 30, 6) */,
  32'h3d14b9d3 /* (25, 30, 6) */,
  32'h3d343ccb /* (21, 30, 6) */,
  32'h3d4bfe66 /* (17, 30, 6) */,
  32'h3d4ce87b /* (13, 30, 6) */,
  32'h3d1e19af /* (9, 30, 6) */,
  32'h3d18df8d /* (5, 30, 6) */,
  32'h3d3543e4 /* (1, 30, 6) */,
  32'h3d14c14d /* (29, 26, 6) */,
  32'h3d20f672 /* (25, 26, 6) */,
  32'h3d5d3b5c /* (21, 26, 6) */,
  32'h3d85e8bf /* (17, 26, 6) */,
  32'h3d82bc35 /* (13, 26, 6) */,
  32'h3d37f9d0 /* (9, 26, 6) */,
  32'h3d16bb8b /* (5, 26, 6) */,
  32'h3d15cc97 /* (1, 26, 6) */,
  32'h3d2c3293 /* (29, 22, 6) */,
  32'h3d5a2934 /* (25, 22, 6) */,
  32'h3dac23aa /* (21, 22, 6) */,
  32'h3de44bb3 /* (17, 22, 6) */,
  32'h3dd610ea /* (13, 22, 6) */,
  32'h3d866682 /* (9, 22, 6) */,
  32'h3d3c300c /* (5, 22, 6) */,
  32'h3d2567ce /* (1, 22, 6) */,
  32'h3d5a5169 /* (29, 18, 6) */,
  32'h3d975464 /* (25, 18, 6) */,
  32'h3e040b60 /* (21, 18, 6) */,
  32'h3e3e01e0 /* (17, 18, 6) */,
  32'h3e2b8c37 /* (13, 18, 6) */,
  32'h3dc45939 /* (9, 18, 6) */,
  32'h3d786cd6 /* (5, 18, 6) */,
  32'h3d4cf093 /* (1, 18, 6) */,
  32'h3d5a5169 /* (29, 14, 6) */,
  32'h3d975464 /* (25, 14, 6) */,
  32'h3e040b60 /* (21, 14, 6) */,
  32'h3e3e01e0 /* (17, 14, 6) */,
  32'h3e2b8c37 /* (13, 14, 6) */,
  32'h3dc45939 /* (9, 14, 6) */,
  32'h3d786cd6 /* (5, 14, 6) */,
  32'h3d4cf093 /* (1, 14, 6) */,
  32'h3d2c3293 /* (29, 10, 6) */,
  32'h3d5a2934 /* (25, 10, 6) */,
  32'h3dac23aa /* (21, 10, 6) */,
  32'h3de44bb3 /* (17, 10, 6) */,
  32'h3dd610ea /* (13, 10, 6) */,
  32'h3d866682 /* (9, 10, 6) */,
  32'h3d3c300c /* (5, 10, 6) */,
  32'h3d2567ce /* (1, 10, 6) */,
  32'h3d14c14d /* (29, 6, 6) */,
  32'h3d20f672 /* (25, 6, 6) */,
  32'h3d5d3b5c /* (21, 6, 6) */,
  32'h3d85e8bf /* (17, 6, 6) */,
  32'h3d82bc35 /* (13, 6, 6) */,
  32'h3d37f9d0 /* (9, 6, 6) */,
  32'h3d16bb8b /* (5, 6, 6) */,
  32'h3d15cc97 /* (1, 6, 6) */,
  32'h3d271e8d /* (29, 2, 6) */,
  32'h3d14b9d3 /* (25, 2, 6) */,
  32'h3d343ccb /* (21, 2, 6) */,
  32'h3d4bfe66 /* (17, 2, 6) */,
  32'h3d4ce87b /* (13, 2, 6) */,
  32'h3d1e19af /* (9, 2, 6) */,
  32'h3d18df8d /* (5, 2, 6) */,
  32'h3d3543e4 /* (1, 2, 6) */,
  32'h3da3af74 /* (29, 30, 2) */,
  32'h3d1dd271 /* (25, 30, 2) */,
  32'h3d18e0f8 /* (21, 30, 2) */,
  32'h3d1dadb9 /* (17, 30, 2) */,
  32'h3d246fbd /* (13, 30, 2) */,
  32'h3d1214c5 /* (9, 30, 2) */,
  32'h3d4ca49b /* (5, 30, 2) */,
  32'h3e0c4d23 /* (1, 30, 2) */,
  32'h3d271e8d /* (29, 26, 2) */,
  32'h3d14b9d3 /* (25, 26, 2) */,
  32'h3d343ccb /* (21, 26, 2) */,
  32'h3d4bfe66 /* (17, 26, 2) */,
  32'h3d4ce87b /* (13, 26, 2) */,
  32'h3d1e19af /* (9, 26, 2) */,
  32'h3d18df8d /* (5, 26, 2) */,
  32'h3d3543e4 /* (1, 26, 2) */,
  32'h3d162b76 /* (29, 22, 2) */,
  32'h3d3346c6 /* (25, 22, 2) */,
  32'h3d85a0b3 /* (21, 22, 2) */,
  32'h3daa3ec9 /* (17, 22, 2) */,
  32'h3da2895a /* (13, 22, 2) */,
  32'h3d56480e /* (9, 22, 2) */,
  32'h3d1f9f49 /* (5, 22, 2) */,
  32'h3d12ac07 /* (1, 22, 2) */,
  32'h3d2b1735 /* (29, 18, 2) */,
  32'h3d6820b1 /* (25, 18, 2) */,
  32'h3dc55f41 /* (21, 18, 2) */,
  32'h3e0adb0d /* (17, 18, 2) */,
  32'h3dfd653f /* (13, 18, 2) */,
  32'h3d94a37c /* (9, 18, 2) */,
  32'h3d40d8bf /* (5, 18, 2) */,
  32'h3d217487 /* (1, 18, 2) */,
  32'h3d2b1735 /* (29, 14, 2) */,
  32'h3d6820b1 /* (25, 14, 2) */,
  32'h3dc55f41 /* (21, 14, 2) */,
  32'h3e0adb0d /* (17, 14, 2) */,
  32'h3dfd653f /* (13, 14, 2) */,
  32'h3d94a37c /* (9, 14, 2) */,
  32'h3d40d8bf /* (5, 14, 2) */,
  32'h3d217487 /* (1, 14, 2) */,
  32'h3d162b76 /* (29, 10, 2) */,
  32'h3d3346c6 /* (25, 10, 2) */,
  32'h3d85a0b3 /* (21, 10, 2) */,
  32'h3daa3ec9 /* (17, 10, 2) */,
  32'h3da2895a /* (13, 10, 2) */,
  32'h3d56480e /* (9, 10, 2) */,
  32'h3d1f9f49 /* (5, 10, 2) */,
  32'h3d12ac07 /* (1, 10, 2) */,
  32'h3d271e8d /* (29, 6, 2) */,
  32'h3d14b9d3 /* (25, 6, 2) */,
  32'h3d343ccb /* (21, 6, 2) */,
  32'h3d4bfe66 /* (17, 6, 2) */,
  32'h3d4ce87b /* (13, 6, 2) */,
  32'h3d1e19af /* (9, 6, 2) */,
  32'h3d18df8d /* (5, 6, 2) */,
  32'h3d3543e4 /* (1, 6, 2) */,
  32'h3da3af74 /* (29, 2, 2) */,
  32'h3d1dd271 /* (25, 2, 2) */,
  32'h3d18e0f8 /* (21, 2, 2) */,
  32'h3d1dadb9 /* (17, 2, 2) */,
  32'h3d246fbd /* (13, 2, 2) */,
  32'h3d1214c5 /* (9, 2, 2) */,
  32'h3d4ca49b /* (5, 2, 2) */,
  32'h3e0c4d23 /* (1, 2, 2) */,
  32'h3d7c66bd /* (28, 30, 30) */,
  32'h3d14e1d9 /* (24, 30, 30) */,
  32'h3d1f454c /* (20, 30, 30) */,
  32'h3d0d5b74 /* (16, 30, 30) */,
  32'h3d1f454c /* (12, 30, 30) */,
  32'h3d14e1d9 /* (8, 30, 30) */,
  32'h3d7c66bd /* (4, 30, 30) */,
  32'h3e1befb2 /* (0, 30, 30) */,
  32'h3d1f2a5d /* (28, 26, 30) */,
  32'h3d17a967 /* (24, 26, 30) */,
  32'h3d41987e /* (20, 26, 30) */,
  32'h3d39823a /* (16, 26, 30) */,
  32'h3d41987e /* (12, 26, 30) */,
  32'h3d17a967 /* (8, 26, 30) */,
  32'h3d1f2a5d /* (4, 26, 30) */,
  32'h3d378ea1 /* (0, 26, 30) */,
  32'h3d19eb69 /* (28, 22, 30) */,
  32'h3d428d9a /* (24, 22, 30) */,
  32'h3d94d2ae /* (20, 22, 30) */,
  32'h3d9e09be /* (16, 22, 30) */,
  32'h3d94d2ae /* (12, 22, 30) */,
  32'h3d428d9a /* (8, 22, 30) */,
  32'h3d19eb69 /* (4, 22, 30) */,
  32'h3d124c17 /* (0, 22, 30) */,
  32'h3d3430e1 /* (28, 18, 30) */,
  32'h3d8271c0 /* (24, 18, 30) */,
  32'h3de2162b /* (20, 18, 30) */,
  32'h3e0374c7 /* (16, 18, 30) */,
  32'h3de2162b /* (12, 18, 30) */,
  32'h3d8271c0 /* (8, 18, 30) */,
  32'h3d3430e1 /* (4, 18, 30) */,
  32'h3d204e75 /* (0, 18, 30) */,
  32'h3d3430e1 /* (28, 14, 30) */,
  32'h3d8271c0 /* (24, 14, 30) */,
  32'h3de2162b /* (20, 14, 30) */,
  32'h3e0374c7 /* (16, 14, 30) */,
  32'h3de2162b /* (12, 14, 30) */,
  32'h3d8271c0 /* (8, 14, 30) */,
  32'h3d3430e1 /* (4, 14, 30) */,
  32'h3d204e75 /* (0, 14, 30) */,
  32'h3d19eb69 /* (28, 10, 30) */,
  32'h3d428d9a /* (24, 10, 30) */,
  32'h3d94d2ae /* (20, 10, 30) */,
  32'h3d9e09be /* (16, 10, 30) */,
  32'h3d94d2ae /* (12, 10, 30) */,
  32'h3d428d9a /* (8, 10, 30) */,
  32'h3d19eb69 /* (4, 10, 30) */,
  32'h3d124c17 /* (0, 10, 30) */,
  32'h3d1f2a5d /* (28, 6, 30) */,
  32'h3d17a967 /* (24, 6, 30) */,
  32'h3d41987e /* (20, 6, 30) */,
  32'h3d39823a /* (16, 6, 30) */,
  32'h3d41987e /* (12, 6, 30) */,
  32'h3d17a967 /* (8, 6, 30) */,
  32'h3d1f2a5d /* (4, 6, 30) */,
  32'h3d378ea1 /* (0, 6, 30) */,
  32'h3d7c66bd /* (28, 2, 30) */,
  32'h3d14e1d9 /* (24, 2, 30) */,
  32'h3d1f454c /* (20, 2, 30) */,
  32'h3d0d5b74 /* (16, 2, 30) */,
  32'h3d1f454c /* (12, 2, 30) */,
  32'h3d14e1d9 /* (8, 2, 30) */,
  32'h3d7c66bd /* (4, 2, 30) */,
  32'h3e1befb2 /* (0, 2, 30) */,
  32'h3d1f2a5d /* (28, 30, 26) */,
  32'h3d17a967 /* (24, 30, 26) */,
  32'h3d41987e /* (20, 30, 26) */,
  32'h3d39823a /* (16, 30, 26) */,
  32'h3d41987e /* (12, 30, 26) */,
  32'h3d17a967 /* (8, 30, 26) */,
  32'h3d1f2a5d /* (4, 30, 26) */,
  32'h3d378ea1 /* (0, 30, 26) */,
  32'h3d1508f6 /* (28, 26, 26) */,
  32'h3d2aa638 /* (24, 26, 26) */,
  32'h3d72a853 /* (20, 26, 26) */,
  32'h3d765452 /* (16, 26, 26) */,
  32'h3d72a853 /* (12, 26, 26) */,
  32'h3d2aa638 /* (8, 26, 26) */,
  32'h3d1508f6 /* (4, 26, 26) */,
  32'h3d160c85 /* (0, 26, 26) */,
  32'h3d32cc97 /* (28, 22, 26) */,
  32'h3d7076ff /* (24, 22, 26) */,
  32'h3dc1f419 /* (20, 22, 26) */,
  32'h3dd58e62 /* (16, 22, 26) */,
  32'h3dc1f419 /* (12, 22, 26) */,
  32'h3d7076ff /* (8, 22, 26) */,
  32'h3d32cc97 /* (4, 22, 26) */,
  32'h3d249cf9 /* (0, 22, 26) */,
  32'h3d66ec8b /* (28, 18, 26) */,
  32'h3dab2ff1 /* (24, 18, 26) */,
  32'h3e182d5a /* (20, 18, 26) */,
  32'h3e34be0d /* (16, 18, 26) */,
  32'h3e182d5a /* (12, 18, 26) */,
  32'h3dab2ff1 /* (8, 18, 26) */,
  32'h3d66ec8b /* (4, 18, 26) */,
  32'h3d4b578e /* (0, 18, 26) */,
  32'h3d66ec8b /* (28, 14, 26) */,
  32'h3dab2ff1 /* (24, 14, 26) */,
  32'h3e182d5a /* (20, 14, 26) */,
  32'h3e34be0d /* (16, 14, 26) */,
  32'h3e182d5a /* (12, 14, 26) */,
  32'h3dab2ff1 /* (8, 14, 26) */,
  32'h3d66ec8b /* (4, 14, 26) */,
  32'h3d4b578e /* (0, 14, 26) */,
  32'h3d32cc97 /* (28, 10, 26) */,
  32'h3d7076ff /* (24, 10, 26) */,
  32'h3dc1f419 /* (20, 10, 26) */,
  32'h3dd58e62 /* (16, 10, 26) */,
  32'h3dc1f419 /* (12, 10, 26) */,
  32'h3d7076ff /* (8, 10, 26) */,
  32'h3d32cc97 /* (4, 10, 26) */,
  32'h3d249cf9 /* (0, 10, 26) */,
  32'h3d1508f6 /* (28, 6, 26) */,
  32'h3d2aa638 /* (24, 6, 26) */,
  32'h3d72a853 /* (20, 6, 26) */,
  32'h3d765452 /* (16, 6, 26) */,
  32'h3d72a853 /* (12, 6, 26) */,
  32'h3d2aa638 /* (8, 6, 26) */,
  32'h3d1508f6 /* (4, 6, 26) */,
  32'h3d160c85 /* (0, 6, 26) */,
  32'h3d1f2a5d /* (28, 2, 26) */,
  32'h3d17a967 /* (24, 2, 26) */,
  32'h3d41987e /* (20, 2, 26) */,
  32'h3d39823a /* (16, 2, 26) */,
  32'h3d41987e /* (12, 2, 26) */,
  32'h3d17a967 /* (8, 2, 26) */,
  32'h3d1f2a5d /* (4, 2, 26) */,
  32'h3d378ea1 /* (0, 2, 26) */,
  32'h3d19eb69 /* (28, 30, 22) */,
  32'h3d428d9a /* (24, 30, 22) */,
  32'h3d94d2ae /* (20, 30, 22) */,
  32'h3d9e09be /* (16, 30, 22) */,
  32'h3d94d2ae /* (12, 30, 22) */,
  32'h3d428d9a /* (8, 30, 22) */,
  32'h3d19eb69 /* (4, 30, 22) */,
  32'h3d124c17 /* (0, 30, 22) */,
  32'h3d32cc97 /* (28, 26, 22) */,
  32'h3d7076ff /* (24, 26, 22) */,
  32'h3dc1f419 /* (20, 26, 22) */,
  32'h3dd58e62 /* (16, 26, 22) */,
  32'h3dc1f419 /* (12, 26, 22) */,
  32'h3d7076ff /* (8, 26, 22) */,
  32'h3d32cc97 /* (4, 26, 22) */,
  32'h3d249cf9 /* (0, 26, 22) */,
  32'h3d825da2 /* (28, 22, 22) */,
  32'h3dbcbfdf /* (24, 22, 22) */,
  32'h3e239217 /* (20, 22, 22) */,
  32'h3e3e36ae /* (16, 22, 22) */,
  32'h3e239217 /* (12, 22, 22) */,
  32'h3dbcbfdf /* (8, 22, 22) */,
  32'h3d825da2 /* (4, 22, 22) */,
  32'h3d67f590 /* (0, 22, 22) */,
  32'h3dbe2f24 /* (28, 18, 22) */,
  32'h3e11d65f /* (24, 18, 22) */,
  32'h3e86bd25 /* (20, 18, 22) */,
  32'h3ea58eba /* (16, 18, 22) */,
  32'h3e86bd25 /* (12, 18, 22) */,
  32'h3e11d65f /* (8, 18, 22) */,
  32'h3dbe2f24 /* (4, 18, 22) */,
  32'h3da521d3 /* (0, 18, 22) */,
  32'h3dbe2f24 /* (28, 14, 22) */,
  32'h3e11d65f /* (24, 14, 22) */,
  32'h3e86bd25 /* (20, 14, 22) */,
  32'h3ea58eba /* (16, 14, 22) */,
  32'h3e86bd25 /* (12, 14, 22) */,
  32'h3e11d65f /* (8, 14, 22) */,
  32'h3dbe2f24 /* (4, 14, 22) */,
  32'h3da521d3 /* (0, 14, 22) */,
  32'h3d825da2 /* (28, 10, 22) */,
  32'h3dbcbfdf /* (24, 10, 22) */,
  32'h3e239217 /* (20, 10, 22) */,
  32'h3e3e36ae /* (16, 10, 22) */,
  32'h3e239217 /* (12, 10, 22) */,
  32'h3dbcbfdf /* (8, 10, 22) */,
  32'h3d825da2 /* (4, 10, 22) */,
  32'h3d67f590 /* (0, 10, 22) */,
  32'h3d32cc97 /* (28, 6, 22) */,
  32'h3d7076ff /* (24, 6, 22) */,
  32'h3dc1f419 /* (20, 6, 22) */,
  32'h3dd58e62 /* (16, 6, 22) */,
  32'h3dc1f419 /* (12, 6, 22) */,
  32'h3d7076ff /* (8, 6, 22) */,
  32'h3d32cc97 /* (4, 6, 22) */,
  32'h3d249cf9 /* (0, 6, 22) */,
  32'h3d19eb69 /* (28, 2, 22) */,
  32'h3d428d9a /* (24, 2, 22) */,
  32'h3d94d2ae /* (20, 2, 22) */,
  32'h3d9e09be /* (16, 2, 22) */,
  32'h3d94d2ae /* (12, 2, 22) */,
  32'h3d428d9a /* (8, 2, 22) */,
  32'h3d19eb69 /* (4, 2, 22) */,
  32'h3d124c17 /* (0, 2, 22) */,
  32'h3d3430e1 /* (28, 30, 18) */,
  32'h3d8271c0 /* (24, 30, 18) */,
  32'h3de2162b /* (20, 30, 18) */,
  32'h3e0374c7 /* (16, 30, 18) */,
  32'h3de2162b /* (12, 30, 18) */,
  32'h3d8271c0 /* (8, 30, 18) */,
  32'h3d3430e1 /* (4, 30, 18) */,
  32'h3d204e75 /* (0, 30, 18) */,
  32'h3d66ec8b /* (28, 26, 18) */,
  32'h3dab2ff1 /* (24, 26, 18) */,
  32'h3e182d5a /* (20, 26, 18) */,
  32'h3e34be0d /* (16, 26, 18) */,
  32'h3e182d5a /* (12, 26, 18) */,
  32'h3dab2ff1 /* (8, 26, 18) */,
  32'h3d66ec8b /* (4, 26, 18) */,
  32'h3d4b578e /* (0, 26, 18) */,
  32'h3dbe2f24 /* (28, 22, 18) */,
  32'h3e11d65f /* (24, 22, 18) */,
  32'h3e86bd25 /* (20, 22, 18) */,
  32'h3ea58eba /* (16, 22, 18) */,
  32'h3e86bd25 /* (12, 22, 18) */,
  32'h3e11d65f /* (8, 22, 18) */,
  32'h3dbe2f24 /* (4, 22, 18) */,
  32'h3da521d3 /* (0, 22, 18) */,
  32'h3e193b79 /* (28, 18, 18) */,
  32'h3e729d82 /* (24, 18, 18) */,
  32'h3ee912bc /* (20, 18, 18) */,
  32'h3f14977b /* (16, 18, 18) */,
  32'h3ee912bc /* (12, 18, 18) */,
  32'h3e729d82 /* (8, 18, 18) */,
  32'h3e193b79 /* (4, 18, 18) */,
  32'h3e036079 /* (0, 18, 18) */,
  32'h3e193b79 /* (28, 14, 18) */,
  32'h3e729d82 /* (24, 14, 18) */,
  32'h3ee912bc /* (20, 14, 18) */,
  32'h3f14977b /* (16, 14, 18) */,
  32'h3ee912bc /* (12, 14, 18) */,
  32'h3e729d82 /* (8, 14, 18) */,
  32'h3e193b79 /* (4, 14, 18) */,
  32'h3e036079 /* (0, 14, 18) */,
  32'h3dbe2f24 /* (28, 10, 18) */,
  32'h3e11d65f /* (24, 10, 18) */,
  32'h3e86bd25 /* (20, 10, 18) */,
  32'h3ea58eba /* (16, 10, 18) */,
  32'h3e86bd25 /* (12, 10, 18) */,
  32'h3e11d65f /* (8, 10, 18) */,
  32'h3dbe2f24 /* (4, 10, 18) */,
  32'h3da521d3 /* (0, 10, 18) */,
  32'h3d66ec8b /* (28, 6, 18) */,
  32'h3dab2ff1 /* (24, 6, 18) */,
  32'h3e182d5a /* (20, 6, 18) */,
  32'h3e34be0d /* (16, 6, 18) */,
  32'h3e182d5a /* (12, 6, 18) */,
  32'h3dab2ff1 /* (8, 6, 18) */,
  32'h3d66ec8b /* (4, 6, 18) */,
  32'h3d4b578e /* (0, 6, 18) */,
  32'h3d3430e1 /* (28, 2, 18) */,
  32'h3d8271c0 /* (24, 2, 18) */,
  32'h3de2162b /* (20, 2, 18) */,
  32'h3e0374c7 /* (16, 2, 18) */,
  32'h3de2162b /* (12, 2, 18) */,
  32'h3d8271c0 /* (8, 2, 18) */,
  32'h3d3430e1 /* (4, 2, 18) */,
  32'h3d204e75 /* (0, 2, 18) */,
  32'h3d3430e1 /* (28, 30, 14) */,
  32'h3d8271c0 /* (24, 30, 14) */,
  32'h3de2162b /* (20, 30, 14) */,
  32'h3e0374c7 /* (16, 30, 14) */,
  32'h3de2162b /* (12, 30, 14) */,
  32'h3d8271c0 /* (8, 30, 14) */,
  32'h3d3430e1 /* (4, 30, 14) */,
  32'h3d204e75 /* (0, 30, 14) */,
  32'h3d66ec8b /* (28, 26, 14) */,
  32'h3dab2ff1 /* (24, 26, 14) */,
  32'h3e182d5a /* (20, 26, 14) */,
  32'h3e34be0d /* (16, 26, 14) */,
  32'h3e182d5a /* (12, 26, 14) */,
  32'h3dab2ff1 /* (8, 26, 14) */,
  32'h3d66ec8b /* (4, 26, 14) */,
  32'h3d4b578e /* (0, 26, 14) */,
  32'h3dbe2f24 /* (28, 22, 14) */,
  32'h3e11d65f /* (24, 22, 14) */,
  32'h3e86bd25 /* (20, 22, 14) */,
  32'h3ea58eba /* (16, 22, 14) */,
  32'h3e86bd25 /* (12, 22, 14) */,
  32'h3e11d65f /* (8, 22, 14) */,
  32'h3dbe2f24 /* (4, 22, 14) */,
  32'h3da521d3 /* (0, 22, 14) */,
  32'h3e193b79 /* (28, 18, 14) */,
  32'h3e729d82 /* (24, 18, 14) */,
  32'h3ee912bc /* (20, 18, 14) */,
  32'h3f14977b /* (16, 18, 14) */,
  32'h3ee912bc /* (12, 18, 14) */,
  32'h3e729d82 /* (8, 18, 14) */,
  32'h3e193b79 /* (4, 18, 14) */,
  32'h3e036079 /* (0, 18, 14) */,
  32'h3e193b79 /* (28, 14, 14) */,
  32'h3e729d82 /* (24, 14, 14) */,
  32'h3ee912bc /* (20, 14, 14) */,
  32'h3f14977b /* (16, 14, 14) */,
  32'h3ee912bc /* (12, 14, 14) */,
  32'h3e729d82 /* (8, 14, 14) */,
  32'h3e193b79 /* (4, 14, 14) */,
  32'h3e036079 /* (0, 14, 14) */,
  32'h3dbe2f24 /* (28, 10, 14) */,
  32'h3e11d65f /* (24, 10, 14) */,
  32'h3e86bd25 /* (20, 10, 14) */,
  32'h3ea58eba /* (16, 10, 14) */,
  32'h3e86bd25 /* (12, 10, 14) */,
  32'h3e11d65f /* (8, 10, 14) */,
  32'h3dbe2f24 /* (4, 10, 14) */,
  32'h3da521d3 /* (0, 10, 14) */,
  32'h3d66ec8b /* (28, 6, 14) */,
  32'h3dab2ff1 /* (24, 6, 14) */,
  32'h3e182d5a /* (20, 6, 14) */,
  32'h3e34be0d /* (16, 6, 14) */,
  32'h3e182d5a /* (12, 6, 14) */,
  32'h3dab2ff1 /* (8, 6, 14) */,
  32'h3d66ec8b /* (4, 6, 14) */,
  32'h3d4b578e /* (0, 6, 14) */,
  32'h3d3430e1 /* (28, 2, 14) */,
  32'h3d8271c0 /* (24, 2, 14) */,
  32'h3de2162b /* (20, 2, 14) */,
  32'h3e0374c7 /* (16, 2, 14) */,
  32'h3de2162b /* (12, 2, 14) */,
  32'h3d8271c0 /* (8, 2, 14) */,
  32'h3d3430e1 /* (4, 2, 14) */,
  32'h3d204e75 /* (0, 2, 14) */,
  32'h3d19eb69 /* (28, 30, 10) */,
  32'h3d428d9a /* (24, 30, 10) */,
  32'h3d94d2ae /* (20, 30, 10) */,
  32'h3d9e09be /* (16, 30, 10) */,
  32'h3d94d2ae /* (12, 30, 10) */,
  32'h3d428d9a /* (8, 30, 10) */,
  32'h3d19eb69 /* (4, 30, 10) */,
  32'h3d124c17 /* (0, 30, 10) */,
  32'h3d32cc97 /* (28, 26, 10) */,
  32'h3d7076ff /* (24, 26, 10) */,
  32'h3dc1f419 /* (20, 26, 10) */,
  32'h3dd58e62 /* (16, 26, 10) */,
  32'h3dc1f419 /* (12, 26, 10) */,
  32'h3d7076ff /* (8, 26, 10) */,
  32'h3d32cc97 /* (4, 26, 10) */,
  32'h3d249cf9 /* (0, 26, 10) */,
  32'h3d825da2 /* (28, 22, 10) */,
  32'h3dbcbfdf /* (24, 22, 10) */,
  32'h3e239217 /* (20, 22, 10) */,
  32'h3e3e36ae /* (16, 22, 10) */,
  32'h3e239217 /* (12, 22, 10) */,
  32'h3dbcbfdf /* (8, 22, 10) */,
  32'h3d825da2 /* (4, 22, 10) */,
  32'h3d67f590 /* (0, 22, 10) */,
  32'h3dbe2f24 /* (28, 18, 10) */,
  32'h3e11d65f /* (24, 18, 10) */,
  32'h3e86bd25 /* (20, 18, 10) */,
  32'h3ea58eba /* (16, 18, 10) */,
  32'h3e86bd25 /* (12, 18, 10) */,
  32'h3e11d65f /* (8, 18, 10) */,
  32'h3dbe2f24 /* (4, 18, 10) */,
  32'h3da521d3 /* (0, 18, 10) */,
  32'h3dbe2f24 /* (28, 14, 10) */,
  32'h3e11d65f /* (24, 14, 10) */,
  32'h3e86bd25 /* (20, 14, 10) */,
  32'h3ea58eba /* (16, 14, 10) */,
  32'h3e86bd25 /* (12, 14, 10) */,
  32'h3e11d65f /* (8, 14, 10) */,
  32'h3dbe2f24 /* (4, 14, 10) */,
  32'h3da521d3 /* (0, 14, 10) */,
  32'h3d825da2 /* (28, 10, 10) */,
  32'h3dbcbfdf /* (24, 10, 10) */,
  32'h3e239217 /* (20, 10, 10) */,
  32'h3e3e36ae /* (16, 10, 10) */,
  32'h3e239217 /* (12, 10, 10) */,
  32'h3dbcbfdf /* (8, 10, 10) */,
  32'h3d825da2 /* (4, 10, 10) */,
  32'h3d67f590 /* (0, 10, 10) */,
  32'h3d32cc97 /* (28, 6, 10) */,
  32'h3d7076ff /* (24, 6, 10) */,
  32'h3dc1f419 /* (20, 6, 10) */,
  32'h3dd58e62 /* (16, 6, 10) */,
  32'h3dc1f419 /* (12, 6, 10) */,
  32'h3d7076ff /* (8, 6, 10) */,
  32'h3d32cc97 /* (4, 6, 10) */,
  32'h3d249cf9 /* (0, 6, 10) */,
  32'h3d19eb69 /* (28, 2, 10) */,
  32'h3d428d9a /* (24, 2, 10) */,
  32'h3d94d2ae /* (20, 2, 10) */,
  32'h3d9e09be /* (16, 2, 10) */,
  32'h3d94d2ae /* (12, 2, 10) */,
  32'h3d428d9a /* (8, 2, 10) */,
  32'h3d19eb69 /* (4, 2, 10) */,
  32'h3d124c17 /* (0, 2, 10) */,
  32'h3d1f2a5d /* (28, 30, 6) */,
  32'h3d17a967 /* (24, 30, 6) */,
  32'h3d41987e /* (20, 30, 6) */,
  32'h3d39823a /* (16, 30, 6) */,
  32'h3d41987e /* (12, 30, 6) */,
  32'h3d17a967 /* (8, 30, 6) */,
  32'h3d1f2a5d /* (4, 30, 6) */,
  32'h3d378ea1 /* (0, 30, 6) */,
  32'h3d1508f6 /* (28, 26, 6) */,
  32'h3d2aa638 /* (24, 26, 6) */,
  32'h3d72a853 /* (20, 26, 6) */,
  32'h3d765452 /* (16, 26, 6) */,
  32'h3d72a853 /* (12, 26, 6) */,
  32'h3d2aa638 /* (8, 26, 6) */,
  32'h3d1508f6 /* (4, 26, 6) */,
  32'h3d160c85 /* (0, 26, 6) */,
  32'h3d32cc97 /* (28, 22, 6) */,
  32'h3d7076ff /* (24, 22, 6) */,
  32'h3dc1f419 /* (20, 22, 6) */,
  32'h3dd58e62 /* (16, 22, 6) */,
  32'h3dc1f419 /* (12, 22, 6) */,
  32'h3d7076ff /* (8, 22, 6) */,
  32'h3d32cc97 /* (4, 22, 6) */,
  32'h3d249cf9 /* (0, 22, 6) */,
  32'h3d66ec8b /* (28, 18, 6) */,
  32'h3dab2ff1 /* (24, 18, 6) */,
  32'h3e182d5a /* (20, 18, 6) */,
  32'h3e34be0d /* (16, 18, 6) */,
  32'h3e182d5a /* (12, 18, 6) */,
  32'h3dab2ff1 /* (8, 18, 6) */,
  32'h3d66ec8b /* (4, 18, 6) */,
  32'h3d4b578e /* (0, 18, 6) */,
  32'h3d66ec8b /* (28, 14, 6) */,
  32'h3dab2ff1 /* (24, 14, 6) */,
  32'h3e182d5a /* (20, 14, 6) */,
  32'h3e34be0d /* (16, 14, 6) */,
  32'h3e182d5a /* (12, 14, 6) */,
  32'h3dab2ff1 /* (8, 14, 6) */,
  32'h3d66ec8b /* (4, 14, 6) */,
  32'h3d4b578e /* (0, 14, 6) */,
  32'h3d32cc97 /* (28, 10, 6) */,
  32'h3d7076ff /* (24, 10, 6) */,
  32'h3dc1f419 /* (20, 10, 6) */,
  32'h3dd58e62 /* (16, 10, 6) */,
  32'h3dc1f419 /* (12, 10, 6) */,
  32'h3d7076ff /* (8, 10, 6) */,
  32'h3d32cc97 /* (4, 10, 6) */,
  32'h3d249cf9 /* (0, 10, 6) */,
  32'h3d1508f6 /* (28, 6, 6) */,
  32'h3d2aa638 /* (24, 6, 6) */,
  32'h3d72a853 /* (20, 6, 6) */,
  32'h3d765452 /* (16, 6, 6) */,
  32'h3d72a853 /* (12, 6, 6) */,
  32'h3d2aa638 /* (8, 6, 6) */,
  32'h3d1508f6 /* (4, 6, 6) */,
  32'h3d160c85 /* (0, 6, 6) */,
  32'h3d1f2a5d /* (28, 2, 6) */,
  32'h3d17a967 /* (24, 2, 6) */,
  32'h3d41987e /* (20, 2, 6) */,
  32'h3d39823a /* (16, 2, 6) */,
  32'h3d41987e /* (12, 2, 6) */,
  32'h3d17a967 /* (8, 2, 6) */,
  32'h3d1f2a5d /* (4, 2, 6) */,
  32'h3d378ea1 /* (0, 2, 6) */,
  32'h3d7c66bd /* (28, 30, 2) */,
  32'h3d14e1d9 /* (24, 30, 2) */,
  32'h3d1f454c /* (20, 30, 2) */,
  32'h3d0d5b74 /* (16, 30, 2) */,
  32'h3d1f454c /* (12, 30, 2) */,
  32'h3d14e1d9 /* (8, 30, 2) */,
  32'h3d7c66bd /* (4, 30, 2) */,
  32'h3e1befb2 /* (0, 30, 2) */,
  32'h3d1f2a5d /* (28, 26, 2) */,
  32'h3d17a967 /* (24, 26, 2) */,
  32'h3d41987e /* (20, 26, 2) */,
  32'h3d39823a /* (16, 26, 2) */,
  32'h3d41987e /* (12, 26, 2) */,
  32'h3d17a967 /* (8, 26, 2) */,
  32'h3d1f2a5d /* (4, 26, 2) */,
  32'h3d378ea1 /* (0, 26, 2) */,
  32'h3d19eb69 /* (28, 22, 2) */,
  32'h3d428d9a /* (24, 22, 2) */,
  32'h3d94d2ae /* (20, 22, 2) */,
  32'h3d9e09be /* (16, 22, 2) */,
  32'h3d94d2ae /* (12, 22, 2) */,
  32'h3d428d9a /* (8, 22, 2) */,
  32'h3d19eb69 /* (4, 22, 2) */,
  32'h3d124c17 /* (0, 22, 2) */,
  32'h3d3430e1 /* (28, 18, 2) */,
  32'h3d8271c0 /* (24, 18, 2) */,
  32'h3de2162b /* (20, 18, 2) */,
  32'h3e0374c7 /* (16, 18, 2) */,
  32'h3de2162b /* (12, 18, 2) */,
  32'h3d8271c0 /* (8, 18, 2) */,
  32'h3d3430e1 /* (4, 18, 2) */,
  32'h3d204e75 /* (0, 18, 2) */,
  32'h3d3430e1 /* (28, 14, 2) */,
  32'h3d8271c0 /* (24, 14, 2) */,
  32'h3de2162b /* (20, 14, 2) */,
  32'h3e0374c7 /* (16, 14, 2) */,
  32'h3de2162b /* (12, 14, 2) */,
  32'h3d8271c0 /* (8, 14, 2) */,
  32'h3d3430e1 /* (4, 14, 2) */,
  32'h3d204e75 /* (0, 14, 2) */,
  32'h3d19eb69 /* (28, 10, 2) */,
  32'h3d428d9a /* (24, 10, 2) */,
  32'h3d94d2ae /* (20, 10, 2) */,
  32'h3d9e09be /* (16, 10, 2) */,
  32'h3d94d2ae /* (12, 10, 2) */,
  32'h3d428d9a /* (8, 10, 2) */,
  32'h3d19eb69 /* (4, 10, 2) */,
  32'h3d124c17 /* (0, 10, 2) */,
  32'h3d1f2a5d /* (28, 6, 2) */,
  32'h3d17a967 /* (24, 6, 2) */,
  32'h3d41987e /* (20, 6, 2) */,
  32'h3d39823a /* (16, 6, 2) */,
  32'h3d41987e /* (12, 6, 2) */,
  32'h3d17a967 /* (8, 6, 2) */,
  32'h3d1f2a5d /* (4, 6, 2) */,
  32'h3d378ea1 /* (0, 6, 2) */,
  32'h3d7c66bd /* (28, 2, 2) */,
  32'h3d14e1d9 /* (24, 2, 2) */,
  32'h3d1f454c /* (20, 2, 2) */,
  32'h3d0d5b74 /* (16, 2, 2) */,
  32'h3d1f454c /* (12, 2, 2) */,
  32'h3d14e1d9 /* (8, 2, 2) */,
  32'h3d7c66bd /* (4, 2, 2) */,
  32'h3e1befb2 /* (0, 2, 2) */,
  32'h3dbfa8df /* (31, 29, 30) */,
  32'h3d3cd255 /* (27, 29, 30) */,
  32'h3d12f42a /* (23, 29, 30) */,
  32'h3d29e985 /* (19, 29, 30) */,
  32'h3d240321 /* (15, 29, 30) */,
  32'h3d1c5f03 /* (11, 29, 30) */,
  32'h3d1a2949 /* (7, 29, 30) */,
  32'h3d866355 /* (3, 29, 30) */,
  32'h3d20a35e /* (31, 25, 30) */,
  32'h3d14b1c0 /* (27, 25, 30) */,
  32'h3d26a1b5 /* (23, 25, 30) */,
  32'h3d6129ae /* (19, 25, 30) */,
  32'h3d62f778 /* (15, 25, 30) */,
  32'h3d42a7b8 /* (11, 25, 30) */,
  32'h3d1777c7 /* (7, 25, 30) */,
  32'h3d1a2949 /* (3, 25, 30) */,
  32'h3d16ed42 /* (31, 21, 30) */,
  32'h3d29823f /* (27, 21, 30) */,
  32'h3d6d9fa3 /* (23, 21, 30) */,
  32'h3dba5db4 /* (19, 21, 30) */,
  32'h3dc59b81 /* (15, 21, 30) */,
  32'h3d96eb50 /* (11, 21, 30) */,
  32'h3d42a7b8 /* (7, 21, 30) */,
  32'h3d1c5f03 /* (3, 21, 30) */,
  32'h3d1a0745 /* (31, 17, 30) */,
  32'h3d3a7be5 /* (27, 17, 30) */,
  32'h3d9314c2 /* (23, 17, 30) */,
  32'h3e003b1e /* (19, 17, 30) */,
  32'h3e0de5f8 /* (15, 17, 30) */,
  32'h3dc59b81 /* (11, 17, 30) */,
  32'h3d62f778 /* (7, 17, 30) */,
  32'h3d240321 /* (3, 17, 30) */,
  32'h3d214ba3 /* (31, 13, 30) */,
  32'h3d3d84de /* (27, 13, 30) */,
  32'h3d8e358b /* (23, 13, 30) */,
  32'h3dec70da /* (19, 13, 30) */,
  32'h3e003b1e /* (15, 13, 30) */,
  32'h3dba5db4 /* (11, 13, 30) */,
  32'h3d6129ae /* (7, 13, 30) */,
  32'h3d29e985 /* (3, 13, 30) */,
  32'h3d11c69f /* (31, 9, 30) */,
  32'h3d18622e /* (27, 9, 30) */,
  32'h3d42665b /* (23, 9, 30) */,
  32'h3d8e358b /* (19, 9, 30) */,
  32'h3d9314c2 /* (15, 9, 30) */,
  32'h3d6d9fa3 /* (11, 9, 30) */,
  32'h3d26a1b5 /* (7, 9, 30) */,
  32'h3d12f42a /* (3, 9, 30) */,
  32'h3d59109a /* (31, 5, 30) */,
  32'h3d213c91 /* (27, 5, 30) */,
  32'h3d18622e /* (23, 5, 30) */,
  32'h3d3d84de /* (19, 5, 30) */,
  32'h3d3a7be5 /* (15, 5, 30) */,
  32'h3d29823f /* (11, 5, 30) */,
  32'h3d14b1c0 /* (7, 5, 30) */,
  32'h3d3cd255 /* (3, 5, 30) */,
  32'h3e4aeee2 /* (31, 1, 30) */,
  32'h3d59109a /* (27, 1, 30) */,
  32'h3d11c69f /* (23, 1, 30) */,
  32'h3d214ba3 /* (19, 1, 30) */,
  32'h3d1a0745 /* (15, 1, 30) */,
  32'h3d16ed42 /* (11, 1, 30) */,
  32'h3d20a35e /* (7, 1, 30) */,
  32'h3dbfa8df /* (3, 1, 30) */,
  32'h3d2ba889 /* (31, 29, 26) */,
  32'h3d16d305 /* (27, 29, 26) */,
  32'h3d215063 /* (23, 29, 26) */,
  32'h3d54a03b /* (19, 29, 26) */,
  32'h3d54ba37 /* (15, 29, 26) */,
  32'h3d39bb76 /* (11, 29, 26) */,
  32'h3d159d44 /* (7, 29, 26) */,
  32'h3d211f1b /* (3, 29, 26) */,
  32'h3d146a43 /* (31, 25, 26) */,
  32'h3d1b2471 /* (27, 25, 26) */,
  32'h3d45eb5b /* (23, 25, 26) */,
  32'h3d90c8a7 /* (19, 25, 26) */,
  32'h3d95be73 /* (15, 25, 26) */,
  32'h3d71ecf9 /* (11, 25, 26) */,
  32'h3d29a602 /* (7, 25, 26) */,
  32'h3d159d44 /* (3, 25, 26) */,
  32'h3d31191b /* (31, 21, 26) */,
  32'h3d4d9045 /* (27, 21, 26) */,
  32'h3d9750ce /* (23, 21, 26) */,
  32'h3df74dbc /* (19, 21, 26) */,
  32'h3e0533d0 /* (15, 21, 26) */,
  32'h3dc480ba /* (11, 21, 26) */,
  32'h3d71ecf9 /* (7, 21, 26) */,
  32'h3d39bb76 /* (3, 21, 26) */,
  32'h3d46f53f /* (31, 17, 26) */,
  32'h3d73b16f /* (27, 17, 26) */,
  32'h3dc42ad0 /* (23, 17, 26) */,
  32'h3e2ea39a /* (19, 17, 26) */,
  32'h3e430b11 /* (15, 17, 26) */,
  32'h3e0533d0 /* (11, 17, 26) */,
  32'h3d95be73 /* (7, 17, 26) */,
  32'h3d54ba37 /* (3, 17, 26) */,
  32'h3d4876ff /* (31, 13, 26) */,
  32'h3d700ffa /* (27, 13, 26) */,
  32'h3db9d5f4 /* (23, 13, 26) */,
  32'h3e1f113d /* (19, 13, 26) */,
  32'h3e2ea39a /* (15, 13, 26) */,
  32'h3df74dbc /* (11, 13, 26) */,
  32'h3d90c8a7 /* (7, 13, 26) */,
  32'h3d54a03b /* (3, 13, 26) */,
  32'h3d1c53e8 /* (31, 9, 26) */,
  32'h3d2db0cc /* (27, 9, 26) */,
  32'h3d6fd024 /* (23, 9, 26) */,
  32'h3db9d5f4 /* (19, 9, 26) */,
  32'h3dc42ad0 /* (15, 9, 26) */,
  32'h3d9750ce /* (11, 9, 26) */,
  32'h3d45eb5b /* (7, 9, 26) */,
  32'h3d215063 /* (3, 9, 26) */,
  32'h3d1a8b5a /* (31, 5, 26) */,
  32'h3d14f7ce /* (27, 5, 26) */,
  32'h3d2db0cc /* (23, 5, 26) */,
  32'h3d700ffa /* (19, 5, 26) */,
  32'h3d73b16f /* (15, 5, 26) */,
  32'h3d4d9045 /* (11, 5, 26) */,
  32'h3d1b2471 /* (7, 5, 26) */,
  32'h3d16d305 /* (3, 5, 26) */,
  32'h3d3c9698 /* (31, 1, 26) */,
  32'h3d1a8b5a /* (27, 1, 26) */,
  32'h3d1c53e8 /* (23, 1, 26) */,
  32'h3d4876ff /* (19, 1, 26) */,
  32'h3d46f53f /* (15, 1, 26) */,
  32'h3d31191b /* (11, 1, 26) */,
  32'h3d146a43 /* (7, 1, 26) */,
  32'h3d2ba889 /* (3, 1, 26) */,
  32'h3d14c0fd /* (31, 29, 22) */,
  32'h3d2344c4 /* (27, 29, 22) */,
  32'h3d5dae2c /* (23, 29, 22) */,
  32'h3da99659 /* (19, 29, 22) */,
  32'h3db22d06 /* (15, 29, 22) */,
  32'h3d8ae43c /* (11, 29, 22) */,
  32'h3d387393 /* (7, 29, 22) */,
  32'h3d18cb02 /* (3, 29, 22) */,
  32'h3d305430 /* (31, 25, 22) */,
  32'h3d4b3dc7 /* (27, 25, 22) */,
  32'h3d94014f /* (23, 25, 22) */,
  32'h3defa49b /* (19, 25, 22) */,
  32'h3e009a19 /* (15, 25, 22) */,
  32'h3dbf3f1d /* (11, 25, 22) */,
  32'h3d6deb12 /* (7, 25, 22) */,
  32'h3d387393 /* (3, 25, 22) */,
  32'h3d829849 /* (31, 21, 22) */,
  32'h3d9d9380 /* (27, 21, 22) */,
  32'h3df71c69 /* (23, 21, 22) */,
  32'h3e562fb1 /* (19, 21, 22) */,
  32'h3e6c6ac0 /* (15, 21, 22) */,
  32'h3e257fc6 /* (11, 21, 22) */,
  32'h3dbf3f1d /* (7, 21, 22) */,
  32'h3d8ae43c /* (3, 21, 22) */,
  32'h3da5ac70 /* (31, 17, 22) */,
  32'h3dce52e6 /* (27, 17, 22) */,
  32'h3e2b3653 /* (23, 17, 22) */,
  32'h3e9d80fb /* (19, 17, 22) */,
  32'h3eb2925b /* (15, 17, 22) */,
  32'h3e6c6ac0 /* (11, 17, 22) */,
  32'h3e009a19 /* (7, 17, 22) */,
  32'h3db22d06 /* (3, 17, 22) */,
  32'h3d9e7894 /* (31, 13, 22) */,
  32'h3dc29629 /* (27, 13, 22) */,
  32'h3e1d56b2 /* (23, 13, 22) */,
  32'h3e8cbae1 /* (19, 13, 22) */,
  32'h3e9d80fb /* (15, 13, 22) */,
  32'h3e562fb1 /* (11, 13, 22) */,
  32'h3defa49b /* (7, 13, 22) */,
  32'h3da99659 /* (3, 13, 22) */,
  32'h3d52081f /* (31, 9, 22) */,
  32'h3d781ae6 /* (27, 9, 22) */,
  32'h3dbbc730 /* (23, 9, 22) */,
  32'h3e1d56b2 /* (19, 9, 22) */,
  32'h3e2b3653 /* (15, 9, 22) */,
  32'h3df71c69 /* (11, 9, 22) */,
  32'h3d94014f /* (7, 9, 22) */,
  32'h3d5dae2c /* (3, 9, 22) */,
  32'h3d1d9589 /* (31, 5, 22) */,
  32'h3d30fc5a /* (27, 5, 22) */,
  32'h3d781ae6 /* (23, 5, 22) */,
  32'h3dc29629 /* (19, 5, 22) */,
  32'h3dce52e6 /* (15, 5, 22) */,
  32'h3d9d9380 /* (11, 5, 22) */,
  32'h3d4b3dc7 /* (7, 5, 22) */,
  32'h3d2344c4 /* (3, 5, 22) */,
  32'h3d119771 /* (31, 1, 22) */,
  32'h3d1d9589 /* (27, 1, 22) */,
  32'h3d52081f /* (23, 1, 22) */,
  32'h3d9e7894 /* (19, 1, 22) */,
  32'h3da5ac70 /* (15, 1, 22) */,
  32'h3d829849 /* (11, 1, 22) */,
  32'h3d305430 /* (7, 1, 22) */,
  32'h3d14c0fd /* (3, 1, 22) */,
  32'h3d276174 /* (31, 29, 18) */,
  32'h3d487174 /* (27, 29, 18) */,
  32'h3d9b2a7b /* (23, 29, 18) */,
  32'h3e04d0b8 /* (19, 29, 18) */,
  32'h3e11d12f /* (15, 29, 18) */,
  32'h3dce7d45 /* (11, 29, 18) */,
  32'h3d71c736 /* (7, 29, 18) */,
  32'h3d3188e3 /* (3, 29, 18) */,
  32'h3d62906c /* (31, 25, 18) */,
  32'h3d8a0000 /* (27, 25, 18) */,
  32'h3ddc09d8 /* (23, 25, 18) */,
  32'h3e41f14c /* (19, 25, 18) */,
  32'h3e57a44b /* (15, 25, 18) */,
  32'h3e14a5c9 /* (11, 25, 18) */,
  32'h3da8d240 /* (7, 25, 18) */,
  32'h3d71c736 /* (3, 25, 18) */,
  32'h3dc01db4 /* (31, 21, 18) */,
  32'h3deed79f /* (27, 21, 18) */,
  32'h3e458f30 /* (23, 21, 18) */,
  32'h3eb517ce /* (19, 21, 18) */,
  32'h3eccf8ff /* (15, 21, 18) */,
  32'h3e882756 /* (11, 21, 18) */,
  32'h3e14a5c9 /* (7, 21, 18) */,
  32'h3dce7d45 /* (3, 21, 18) */,
  32'h3e06d8bb /* (31, 17, 18) */,
  32'h3e2a981c /* (27, 17, 18) */,
  32'h3e91e4f8 /* (23, 17, 18) */,
  32'h3f0af24f /* (19, 17, 18) */,
  32'h3f202f9a /* (15, 17, 18) */,
  32'h3eccf8ff /* (11, 17, 18) */,
  32'h3e57a44b /* (7, 17, 18) */,
  32'h3e11d12f /* (3, 17, 18) */,
  32'h3df65860 /* (31, 13, 18) */,
  32'h3e1a8d8c /* (27, 13, 18) */,
  32'h3e821787 /* (23, 13, 18) */,
  32'h3ef33ce4 /* (19, 13, 18) */,
  32'h3f0af24f /* (15, 13, 18) */,
  32'h3eb517ce /* (11, 13, 18) */,
  32'h3e41f14c /* (7, 13, 18) */,
  32'h3e04d0b8 /* (3, 13, 18) */,
  32'h3d90dff9 /* (31, 9, 18) */,
  32'h3db24f8e /* (27, 9, 18) */,
  32'h3e10cac5 /* (23, 9, 18) */,
  32'h3e821787 /* (19, 9, 18) */,
  32'h3e91e4f8 /* (15, 9, 18) */,
  32'h3e458f30 /* (11, 9, 18) */,
  32'h3ddc09d8 /* (7, 9, 18) */,
  32'h3d9b2a7b /* (3, 9, 18) */,
  32'h3d3c7841 /* (31, 5, 18) */,
  32'h3d63687e /* (27, 5, 18) */,
  32'h3db24f8e /* (23, 5, 18) */,
  32'h3e1a8d8c /* (19, 5, 18) */,
  32'h3e2a981c /* (15, 5, 18) */,
  32'h3deed79f /* (11, 5, 18) */,
  32'h3d8a0000 /* (7, 5, 18) */,
  32'h3d487174 /* (3, 5, 18) */,
  32'h3d1e0bb6 /* (31, 1, 18) */,
  32'h3d3c7841 /* (27, 1, 18) */,
  32'h3d90dff9 /* (23, 1, 18) */,
  32'h3df65860 /* (19, 1, 18) */,
  32'h3e06d8bb /* (15, 1, 18) */,
  32'h3dc01db4 /* (11, 1, 18) */,
  32'h3d62906c /* (7, 1, 18) */,
  32'h3d276174 /* (3, 1, 18) */,
  32'h3d276174 /* (31, 29, 14) */,
  32'h3d487174 /* (27, 29, 14) */,
  32'h3d9b2a7b /* (23, 29, 14) */,
  32'h3e04d0b8 /* (19, 29, 14) */,
  32'h3e11d12f /* (15, 29, 14) */,
  32'h3dce7d45 /* (11, 29, 14) */,
  32'h3d71c736 /* (7, 29, 14) */,
  32'h3d3188e3 /* (3, 29, 14) */,
  32'h3d62906c /* (31, 25, 14) */,
  32'h3d8a0000 /* (27, 25, 14) */,
  32'h3ddc09d8 /* (23, 25, 14) */,
  32'h3e41f14c /* (19, 25, 14) */,
  32'h3e57a44b /* (15, 25, 14) */,
  32'h3e14a5c9 /* (11, 25, 14) */,
  32'h3da8d240 /* (7, 25, 14) */,
  32'h3d71c736 /* (3, 25, 14) */,
  32'h3dc01db4 /* (31, 21, 14) */,
  32'h3deed79f /* (27, 21, 14) */,
  32'h3e458f30 /* (23, 21, 14) */,
  32'h3eb517ce /* (19, 21, 14) */,
  32'h3eccf8ff /* (15, 21, 14) */,
  32'h3e882756 /* (11, 21, 14) */,
  32'h3e14a5c9 /* (7, 21, 14) */,
  32'h3dce7d45 /* (3, 21, 14) */,
  32'h3e06d8bb /* (31, 17, 14) */,
  32'h3e2a981c /* (27, 17, 14) */,
  32'h3e91e4f8 /* (23, 17, 14) */,
  32'h3f0af24f /* (19, 17, 14) */,
  32'h3f202f9a /* (15, 17, 14) */,
  32'h3eccf8ff /* (11, 17, 14) */,
  32'h3e57a44b /* (7, 17, 14) */,
  32'h3e11d12f /* (3, 17, 14) */,
  32'h3df65860 /* (31, 13, 14) */,
  32'h3e1a8d8c /* (27, 13, 14) */,
  32'h3e821787 /* (23, 13, 14) */,
  32'h3ef33ce4 /* (19, 13, 14) */,
  32'h3f0af24f /* (15, 13, 14) */,
  32'h3eb517ce /* (11, 13, 14) */,
  32'h3e41f14c /* (7, 13, 14) */,
  32'h3e04d0b8 /* (3, 13, 14) */,
  32'h3d90dff9 /* (31, 9, 14) */,
  32'h3db24f8e /* (27, 9, 14) */,
  32'h3e10cac5 /* (23, 9, 14) */,
  32'h3e821787 /* (19, 9, 14) */,
  32'h3e91e4f8 /* (15, 9, 14) */,
  32'h3e458f30 /* (11, 9, 14) */,
  32'h3ddc09d8 /* (7, 9, 14) */,
  32'h3d9b2a7b /* (3, 9, 14) */,
  32'h3d3c7841 /* (31, 5, 14) */,
  32'h3d63687e /* (27, 5, 14) */,
  32'h3db24f8e /* (23, 5, 14) */,
  32'h3e1a8d8c /* (19, 5, 14) */,
  32'h3e2a981c /* (15, 5, 14) */,
  32'h3deed79f /* (11, 5, 14) */,
  32'h3d8a0000 /* (7, 5, 14) */,
  32'h3d487174 /* (3, 5, 14) */,
  32'h3d1e0bb6 /* (31, 1, 14) */,
  32'h3d3c7841 /* (27, 1, 14) */,
  32'h3d90dff9 /* (23, 1, 14) */,
  32'h3df65860 /* (19, 1, 14) */,
  32'h3e06d8bb /* (15, 1, 14) */,
  32'h3dc01db4 /* (11, 1, 14) */,
  32'h3d62906c /* (7, 1, 14) */,
  32'h3d276174 /* (3, 1, 14) */,
  32'h3d14c0fd /* (31, 29, 10) */,
  32'h3d2344c4 /* (27, 29, 10) */,
  32'h3d5dae2c /* (23, 29, 10) */,
  32'h3da99659 /* (19, 29, 10) */,
  32'h3db22d06 /* (15, 29, 10) */,
  32'h3d8ae43c /* (11, 29, 10) */,
  32'h3d387393 /* (7, 29, 10) */,
  32'h3d18cb02 /* (3, 29, 10) */,
  32'h3d305430 /* (31, 25, 10) */,
  32'h3d4b3dc7 /* (27, 25, 10) */,
  32'h3d94014f /* (23, 25, 10) */,
  32'h3defa49b /* (19, 25, 10) */,
  32'h3e009a19 /* (15, 25, 10) */,
  32'h3dbf3f1d /* (11, 25, 10) */,
  32'h3d6deb12 /* (7, 25, 10) */,
  32'h3d387393 /* (3, 25, 10) */,
  32'h3d829849 /* (31, 21, 10) */,
  32'h3d9d9380 /* (27, 21, 10) */,
  32'h3df71c69 /* (23, 21, 10) */,
  32'h3e562fb1 /* (19, 21, 10) */,
  32'h3e6c6ac0 /* (15, 21, 10) */,
  32'h3e257fc6 /* (11, 21, 10) */,
  32'h3dbf3f1d /* (7, 21, 10) */,
  32'h3d8ae43c /* (3, 21, 10) */,
  32'h3da5ac70 /* (31, 17, 10) */,
  32'h3dce52e6 /* (27, 17, 10) */,
  32'h3e2b3653 /* (23, 17, 10) */,
  32'h3e9d80fb /* (19, 17, 10) */,
  32'h3eb2925b /* (15, 17, 10) */,
  32'h3e6c6ac0 /* (11, 17, 10) */,
  32'h3e009a19 /* (7, 17, 10) */,
  32'h3db22d06 /* (3, 17, 10) */,
  32'h3d9e7894 /* (31, 13, 10) */,
  32'h3dc29629 /* (27, 13, 10) */,
  32'h3e1d56b2 /* (23, 13, 10) */,
  32'h3e8cbae1 /* (19, 13, 10) */,
  32'h3e9d80fb /* (15, 13, 10) */,
  32'h3e562fb1 /* (11, 13, 10) */,
  32'h3defa49b /* (7, 13, 10) */,
  32'h3da99659 /* (3, 13, 10) */,
  32'h3d52081f /* (31, 9, 10) */,
  32'h3d781ae6 /* (27, 9, 10) */,
  32'h3dbbc730 /* (23, 9, 10) */,
  32'h3e1d56b2 /* (19, 9, 10) */,
  32'h3e2b3653 /* (15, 9, 10) */,
  32'h3df71c69 /* (11, 9, 10) */,
  32'h3d94014f /* (7, 9, 10) */,
  32'h3d5dae2c /* (3, 9, 10) */,
  32'h3d1d9589 /* (31, 5, 10) */,
  32'h3d30fc5a /* (27, 5, 10) */,
  32'h3d781ae6 /* (23, 5, 10) */,
  32'h3dc29629 /* (19, 5, 10) */,
  32'h3dce52e6 /* (15, 5, 10) */,
  32'h3d9d9380 /* (11, 5, 10) */,
  32'h3d4b3dc7 /* (7, 5, 10) */,
  32'h3d2344c4 /* (3, 5, 10) */,
  32'h3d119771 /* (31, 1, 10) */,
  32'h3d1d9589 /* (27, 1, 10) */,
  32'h3d52081f /* (23, 1, 10) */,
  32'h3d9e7894 /* (19, 1, 10) */,
  32'h3da5ac70 /* (15, 1, 10) */,
  32'h3d829849 /* (11, 1, 10) */,
  32'h3d305430 /* (7, 1, 10) */,
  32'h3d14c0fd /* (3, 1, 10) */,
  32'h3d2ba889 /* (31, 29, 6) */,
  32'h3d16d305 /* (27, 29, 6) */,
  32'h3d215063 /* (23, 29, 6) */,
  32'h3d54a03b /* (19, 29, 6) */,
  32'h3d54ba37 /* (15, 29, 6) */,
  32'h3d39bb76 /* (11, 29, 6) */,
  32'h3d159d44 /* (7, 29, 6) */,
  32'h3d211f1b /* (3, 29, 6) */,
  32'h3d146a43 /* (31, 25, 6) */,
  32'h3d1b2471 /* (27, 25, 6) */,
  32'h3d45eb5b /* (23, 25, 6) */,
  32'h3d90c8a7 /* (19, 25, 6) */,
  32'h3d95be73 /* (15, 25, 6) */,
  32'h3d71ecf9 /* (11, 25, 6) */,
  32'h3d29a602 /* (7, 25, 6) */,
  32'h3d159d44 /* (3, 25, 6) */,
  32'h3d31191b /* (31, 21, 6) */,
  32'h3d4d9045 /* (27, 21, 6) */,
  32'h3d9750ce /* (23, 21, 6) */,
  32'h3df74dbc /* (19, 21, 6) */,
  32'h3e0533d0 /* (15, 21, 6) */,
  32'h3dc480ba /* (11, 21, 6) */,
  32'h3d71ecf9 /* (7, 21, 6) */,
  32'h3d39bb76 /* (3, 21, 6) */,
  32'h3d46f53f /* (31, 17, 6) */,
  32'h3d73b16f /* (27, 17, 6) */,
  32'h3dc42ad0 /* (23, 17, 6) */,
  32'h3e2ea39a /* (19, 17, 6) */,
  32'h3e430b11 /* (15, 17, 6) */,
  32'h3e0533d0 /* (11, 17, 6) */,
  32'h3d95be73 /* (7, 17, 6) */,
  32'h3d54ba37 /* (3, 17, 6) */,
  32'h3d4876ff /* (31, 13, 6) */,
  32'h3d700ffa /* (27, 13, 6) */,
  32'h3db9d5f4 /* (23, 13, 6) */,
  32'h3e1f113d /* (19, 13, 6) */,
  32'h3e2ea39a /* (15, 13, 6) */,
  32'h3df74dbc /* (11, 13, 6) */,
  32'h3d90c8a7 /* (7, 13, 6) */,
  32'h3d54a03b /* (3, 13, 6) */,
  32'h3d1c53e8 /* (31, 9, 6) */,
  32'h3d2db0cc /* (27, 9, 6) */,
  32'h3d6fd024 /* (23, 9, 6) */,
  32'h3db9d5f4 /* (19, 9, 6) */,
  32'h3dc42ad0 /* (15, 9, 6) */,
  32'h3d9750ce /* (11, 9, 6) */,
  32'h3d45eb5b /* (7, 9, 6) */,
  32'h3d215063 /* (3, 9, 6) */,
  32'h3d1a8b5a /* (31, 5, 6) */,
  32'h3d14f7ce /* (27, 5, 6) */,
  32'h3d2db0cc /* (23, 5, 6) */,
  32'h3d700ffa /* (19, 5, 6) */,
  32'h3d73b16f /* (15, 5, 6) */,
  32'h3d4d9045 /* (11, 5, 6) */,
  32'h3d1b2471 /* (7, 5, 6) */,
  32'h3d16d305 /* (3, 5, 6) */,
  32'h3d3c9698 /* (31, 1, 6) */,
  32'h3d1a8b5a /* (27, 1, 6) */,
  32'h3d1c53e8 /* (23, 1, 6) */,
  32'h3d4876ff /* (19, 1, 6) */,
  32'h3d46f53f /* (15, 1, 6) */,
  32'h3d31191b /* (11, 1, 6) */,
  32'h3d146a43 /* (7, 1, 6) */,
  32'h3d2ba889 /* (3, 1, 6) */,
  32'h3dbfa8df /* (31, 29, 2) */,
  32'h3d3cd255 /* (27, 29, 2) */,
  32'h3d12f42a /* (23, 29, 2) */,
  32'h3d29e985 /* (19, 29, 2) */,
  32'h3d240321 /* (15, 29, 2) */,
  32'h3d1c5f03 /* (11, 29, 2) */,
  32'h3d1a2949 /* (7, 29, 2) */,
  32'h3d866355 /* (3, 29, 2) */,
  32'h3d20a35e /* (31, 25, 2) */,
  32'h3d14b1c0 /* (27, 25, 2) */,
  32'h3d26a1b5 /* (23, 25, 2) */,
  32'h3d6129ae /* (19, 25, 2) */,
  32'h3d62f778 /* (15, 25, 2) */,
  32'h3d42a7b8 /* (11, 25, 2) */,
  32'h3d1777c7 /* (7, 25, 2) */,
  32'h3d1a2949 /* (3, 25, 2) */,
  32'h3d16ed42 /* (31, 21, 2) */,
  32'h3d29823f /* (27, 21, 2) */,
  32'h3d6d9fa3 /* (23, 21, 2) */,
  32'h3dba5db4 /* (19, 21, 2) */,
  32'h3dc59b81 /* (15, 21, 2) */,
  32'h3d96eb50 /* (11, 21, 2) */,
  32'h3d42a7b8 /* (7, 21, 2) */,
  32'h3d1c5f03 /* (3, 21, 2) */,
  32'h3d1a0745 /* (31, 17, 2) */,
  32'h3d3a7be5 /* (27, 17, 2) */,
  32'h3d9314c2 /* (23, 17, 2) */,
  32'h3e003b1e /* (19, 17, 2) */,
  32'h3e0de5f8 /* (15, 17, 2) */,
  32'h3dc59b81 /* (11, 17, 2) */,
  32'h3d62f778 /* (7, 17, 2) */,
  32'h3d240321 /* (3, 17, 2) */,
  32'h3d214ba3 /* (31, 13, 2) */,
  32'h3d3d84de /* (27, 13, 2) */,
  32'h3d8e358b /* (23, 13, 2) */,
  32'h3dec70da /* (19, 13, 2) */,
  32'h3e003b1e /* (15, 13, 2) */,
  32'h3dba5db4 /* (11, 13, 2) */,
  32'h3d6129ae /* (7, 13, 2) */,
  32'h3d29e985 /* (3, 13, 2) */,
  32'h3d11c69f /* (31, 9, 2) */,
  32'h3d18622e /* (27, 9, 2) */,
  32'h3d42665b /* (23, 9, 2) */,
  32'h3d8e358b /* (19, 9, 2) */,
  32'h3d9314c2 /* (15, 9, 2) */,
  32'h3d6d9fa3 /* (11, 9, 2) */,
  32'h3d26a1b5 /* (7, 9, 2) */,
  32'h3d12f42a /* (3, 9, 2) */,
  32'h3d59109a /* (31, 5, 2) */,
  32'h3d213c91 /* (27, 5, 2) */,
  32'h3d18622e /* (23, 5, 2) */,
  32'h3d3d84de /* (19, 5, 2) */,
  32'h3d3a7be5 /* (15, 5, 2) */,
  32'h3d29823f /* (11, 5, 2) */,
  32'h3d14b1c0 /* (7, 5, 2) */,
  32'h3d3cd255 /* (3, 5, 2) */,
  32'h3e4aeee2 /* (31, 1, 2) */,
  32'h3d59109a /* (27, 1, 2) */,
  32'h3d11c69f /* (23, 1, 2) */,
  32'h3d214ba3 /* (19, 1, 2) */,
  32'h3d1a0745 /* (15, 1, 2) */,
  32'h3d16ed42 /* (11, 1, 2) */,
  32'h3d20a35e /* (7, 1, 2) */,
  32'h3dbfa8df /* (3, 1, 2) */,
  32'h3da3af74 /* (30, 29, 30) */,
  32'h3d271e8d /* (26, 29, 30) */,
  32'h3d162b76 /* (22, 29, 30) */,
  32'h3d2b1735 /* (18, 29, 30) */,
  32'h3d2b1735 /* (14, 29, 30) */,
  32'h3d162b76 /* (10, 29, 30) */,
  32'h3d271e8d /* (6, 29, 30) */,
  32'h3da3af74 /* (2, 29, 30) */,
  32'h3d1dd271 /* (30, 25, 30) */,
  32'h3d14b9d3 /* (26, 25, 30) */,
  32'h3d3346c6 /* (22, 25, 30) */,
  32'h3d6820b1 /* (18, 25, 30) */,
  32'h3d6820b1 /* (14, 25, 30) */,
  32'h3d3346c6 /* (10, 25, 30) */,
  32'h3d14b9d3 /* (6, 25, 30) */,
  32'h3d1dd271 /* (2, 25, 30) */,
  32'h3d18e0f8 /* (30, 21, 30) */,
  32'h3d343ccb /* (26, 21, 30) */,
  32'h3d85a0b3 /* (22, 21, 30) */,
  32'h3dc55f41 /* (18, 21, 30) */,
  32'h3dc55f41 /* (14, 21, 30) */,
  32'h3d85a0b3 /* (10, 21, 30) */,
  32'h3d343ccb /* (6, 21, 30) */,
  32'h3d18e0f8 /* (2, 21, 30) */,
  32'h3d1dadb9 /* (30, 17, 30) */,
  32'h3d4bfe66 /* (26, 17, 30) */,
  32'h3daa3ec9 /* (22, 17, 30) */,
  32'h3e0adb0d /* (18, 17, 30) */,
  32'h3e0adb0d /* (14, 17, 30) */,
  32'h3daa3ec9 /* (10, 17, 30) */,
  32'h3d4bfe66 /* (6, 17, 30) */,
  32'h3d1dadb9 /* (2, 17, 30) */,
  32'h3d246fbd /* (30, 13, 30) */,
  32'h3d4ce87b /* (26, 13, 30) */,
  32'h3da2895a /* (22, 13, 30) */,
  32'h3dfd653f /* (18, 13, 30) */,
  32'h3dfd653f /* (14, 13, 30) */,
  32'h3da2895a /* (10, 13, 30) */,
  32'h3d4ce87b /* (6, 13, 30) */,
  32'h3d246fbd /* (2, 13, 30) */,
  32'h3d1214c5 /* (30, 9, 30) */,
  32'h3d1e19af /* (26, 9, 30) */,
  32'h3d56480e /* (22, 9, 30) */,
  32'h3d94a37c /* (18, 9, 30) */,
  32'h3d94a37c /* (14, 9, 30) */,
  32'h3d56480e /* (10, 9, 30) */,
  32'h3d1e19af /* (6, 9, 30) */,
  32'h3d1214c5 /* (2, 9, 30) */,
  32'h3d4ca49b /* (30, 5, 30) */,
  32'h3d18df8d /* (26, 5, 30) */,
  32'h3d1f9f49 /* (22, 5, 30) */,
  32'h3d40d8bf /* (18, 5, 30) */,
  32'h3d40d8bf /* (14, 5, 30) */,
  32'h3d1f9f49 /* (10, 5, 30) */,
  32'h3d18df8d /* (6, 5, 30) */,
  32'h3d4ca49b /* (2, 5, 30) */,
  32'h3e0c4d23 /* (30, 1, 30) */,
  32'h3d3543e4 /* (26, 1, 30) */,
  32'h3d12ac07 /* (22, 1, 30) */,
  32'h3d217487 /* (18, 1, 30) */,
  32'h3d217487 /* (14, 1, 30) */,
  32'h3d12ac07 /* (10, 1, 30) */,
  32'h3d3543e4 /* (6, 1, 30) */,
  32'h3e0c4d23 /* (2, 1, 30) */,
  32'h3d271e8d /* (30, 29, 26) */,
  32'h3d14c14d /* (26, 29, 26) */,
  32'h3d2c3293 /* (22, 29, 26) */,
  32'h3d5a5169 /* (18, 29, 26) */,
  32'h3d5a5169 /* (14, 29, 26) */,
  32'h3d2c3293 /* (10, 29, 26) */,
  32'h3d14c14d /* (6, 29, 26) */,
  32'h3d271e8d /* (2, 29, 26) */,
  32'h3d14b9d3 /* (30, 25, 26) */,
  32'h3d20f672 /* (26, 25, 26) */,
  32'h3d5a2934 /* (22, 25, 26) */,
  32'h3d975464 /* (18, 25, 26) */,
  32'h3d975464 /* (14, 25, 26) */,
  32'h3d5a2934 /* (10, 25, 26) */,
  32'h3d20f672 /* (6, 25, 26) */,
  32'h3d14b9d3 /* (2, 25, 26) */,
  32'h3d343ccb /* (30, 21, 26) */,
  32'h3d5d3b5c /* (26, 21, 26) */,
  32'h3dac23aa /* (22, 21, 26) */,
  32'h3e040b60 /* (18, 21, 26) */,
  32'h3e040b60 /* (14, 21, 26) */,
  32'h3dac23aa /* (10, 21, 26) */,
  32'h3d5d3b5c /* (6, 21, 26) */,
  32'h3d343ccb /* (2, 21, 26) */,
  32'h3d4bfe66 /* (30, 17, 26) */,
  32'h3d85e8bf /* (26, 17, 26) */,
  32'h3de44bb3 /* (22, 17, 26) */,
  32'h3e3e01e0 /* (18, 17, 26) */,
  32'h3e3e01e0 /* (14, 17, 26) */,
  32'h3de44bb3 /* (10, 17, 26) */,
  32'h3d85e8bf /* (6, 17, 26) */,
  32'h3d4bfe66 /* (2, 17, 26) */,
  32'h3d4ce87b /* (30, 13, 26) */,
  32'h3d82bc35 /* (26, 13, 26) */,
  32'h3dd610ea /* (22, 13, 26) */,
  32'h3e2b8c37 /* (18, 13, 26) */,
  32'h3e2b8c37 /* (14, 13, 26) */,
  32'h3dd610ea /* (10, 13, 26) */,
  32'h3d82bc35 /* (6, 13, 26) */,
  32'h3d4ce87b /* (2, 13, 26) */,
  32'h3d1e19af /* (30, 9, 26) */,
  32'h3d37f9d0 /* (26, 9, 26) */,
  32'h3d866682 /* (22, 9, 26) */,
  32'h3dc45939 /* (18, 9, 26) */,
  32'h3dc45939 /* (14, 9, 26) */,
  32'h3d866682 /* (10, 9, 26) */,
  32'h3d37f9d0 /* (6, 9, 26) */,
  32'h3d1e19af /* (2, 9, 26) */,
  32'h3d18df8d /* (30, 5, 26) */,
  32'h3d16bb8b /* (26, 5, 26) */,
  32'h3d3c300c /* (22, 5, 26) */,
  32'h3d786cd6 /* (18, 5, 26) */,
  32'h3d786cd6 /* (14, 5, 26) */,
  32'h3d3c300c /* (10, 5, 26) */,
  32'h3d16bb8b /* (6, 5, 26) */,
  32'h3d18df8d /* (2, 5, 26) */,
  32'h3d3543e4 /* (30, 1, 26) */,
  32'h3d15cc97 /* (26, 1, 26) */,
  32'h3d2567ce /* (22, 1, 26) */,
  32'h3d4cf093 /* (18, 1, 26) */,
  32'h3d4cf093 /* (14, 1, 26) */,
  32'h3d2567ce /* (10, 1, 26) */,
  32'h3d15cc97 /* (6, 1, 26) */,
  32'h3d3543e4 /* (2, 1, 26) */,
  32'h3d162b76 /* (30, 29, 22) */,
  32'h3d2c3293 /* (26, 29, 22) */,
  32'h3d77904c /* (22, 29, 22) */,
  32'h3db2bcb9 /* (18, 29, 22) */,
  32'h3db2bcb9 /* (14, 29, 22) */,
  32'h3d77904c /* (10, 29, 22) */,
  32'h3d2c3293 /* (6, 29, 22) */,
  32'h3d162b76 /* (2, 29, 22) */,
  32'h3d3346c6 /* (30, 25, 22) */,
  32'h3d5a2934 /* (26, 25, 22) */,
  32'h3da7f0fb /* (22, 25, 22) */,
  32'h3dff6ab3 /* (18, 25, 22) */,
  32'h3dff6ab3 /* (14, 25, 22) */,
  32'h3da7f0fb /* (10, 25, 22) */,
  32'h3d5a2934 /* (6, 25, 22) */,
  32'h3d3346c6 /* (2, 25, 22) */,
  32'h3d85a0b3 /* (30, 21, 22) */,
  32'h3dac23aa /* (26, 21, 22) */,
  32'h3e0ecbcd /* (22, 21, 22) */,
  32'h3e67a191 /* (18, 21, 22) */,
  32'h3e67a191 /* (14, 21, 22) */,
  32'h3e0ecbcd /* (10, 21, 22) */,
  32'h3dac23aa /* (6, 21, 22) */,
  32'h3d85a0b3 /* (2, 21, 22) */,
  32'h3daa3ec9 /* (30, 17, 22) */,
  32'h3de44bb3 /* (26, 17, 22) */,
  32'h3e48eba4 /* (22, 17, 22) */,
  32'h3eacaf9b /* (18, 17, 22) */,
  32'h3eacaf9b /* (14, 17, 22) */,
  32'h3e48eba4 /* (10, 17, 22) */,
  32'h3de44bb3 /* (6, 17, 22) */,
  32'h3daa3ec9 /* (2, 17, 22) */,
  32'h3da2895a /* (30, 13, 22) */,
  32'h3dd610ea /* (26, 13, 22) */,
  32'h3e37540b /* (22, 13, 22) */,
  32'h3e994798 /* (18, 13, 22) */,
  32'h3e994798 /* (14, 13, 22) */,
  32'h3e37540b /* (10, 13, 22) */,
  32'h3dd610ea /* (6, 13, 22) */,
  32'h3da2895a /* (2, 13, 22) */,
  32'h3d56480e /* (30, 9, 22) */,
  32'h3d866682 /* (26, 9, 22) */,
  32'h3dd7137d /* (22, 9, 22) */,
  32'h3e28e750 /* (18, 9, 22) */,
  32'h3e28e750 /* (14, 9, 22) */,
  32'h3dd7137d /* (10, 9, 22) */,
  32'h3d866682 /* (6, 9, 22) */,
  32'h3d56480e /* (2, 9, 22) */,
  32'h3d1f9f49 /* (30, 5, 22) */,
  32'h3d3c300c /* (26, 5, 22) */,
  32'h3d8b85a2 /* (22, 5, 22) */,
  32'h3dce13fe /* (18, 5, 22) */,
  32'h3dce13fe /* (14, 5, 22) */,
  32'h3d8b85a2 /* (10, 5, 22) */,
  32'h3d3c300c /* (6, 5, 22) */,
  32'h3d1f9f49 /* (2, 5, 22) */,
  32'h3d12ac07 /* (30, 1, 22) */,
  32'h3d2567ce /* (26, 1, 22) */,
  32'h3d699f13 /* (22, 1, 22) */,
  32'h3da6958f /* (18, 1, 22) */,
  32'h3da6958f /* (14, 1, 22) */,
  32'h3d699f13 /* (10, 1, 22) */,
  32'h3d2567ce /* (6, 1, 22) */,
  32'h3d12ac07 /* (2, 1, 22) */,
  32'h3d2b1735 /* (30, 29, 18) */,
  32'h3d5a5169 /* (26, 29, 18) */,
  32'h3db2bcb9 /* (22, 29, 18) */,
  32'h3e0f3c67 /* (18, 29, 18) */,
  32'h3e0f3c67 /* (14, 29, 18) */,
  32'h3db2bcb9 /* (10, 29, 18) */,
  32'h3d5a5169 /* (6, 29, 18) */,
  32'h3d2b1735 /* (2, 29, 18) */,
  32'h3d6820b1 /* (30, 25, 18) */,
  32'h3d975464 /* (26, 25, 18) */,
  32'h3dff6ab3 /* (22, 25, 18) */,
  32'h3e528761 /* (18, 25, 18) */,
  32'h3e528761 /* (14, 25, 18) */,
  32'h3dff6ab3 /* (10, 25, 18) */,
  32'h3d975464 /* (6, 25, 18) */,
  32'h3d6820b1 /* (2, 25, 18) */,
  32'h3dc55f41 /* (30, 21, 18) */,
  32'h3e040b60 /* (26, 21, 18) */,
  32'h3e67a191 /* (22, 21, 18) */,
  32'h3ec66134 /* (18, 21, 18) */,
  32'h3ec66134 /* (14, 21, 18) */,
  32'h3e67a191 /* (10, 21, 18) */,
  32'h3e040b60 /* (6, 21, 18) */,
  32'h3dc55f41 /* (2, 21, 18) */,
  32'h3e0adb0d /* (30, 17, 18) */,
  32'h3e3e01e0 /* (26, 17, 18) */,
  32'h3eacaf9b /* (22, 17, 18) */,
  32'h3f19a2a7 /* (18, 17, 18) */,
  32'h3f19a2a7 /* (14, 17, 18) */,
  32'h3eacaf9b /* (10, 17, 18) */,
  32'h3e3e01e0 /* (6, 17, 18) */,
  32'h3e0adb0d /* (2, 17, 18) */,
  32'h3dfd653f /* (30, 13, 18) */,
  32'h3e2b8c37 /* (26, 13, 18) */,
  32'h3e994798 /* (22, 13, 18) */,
  32'h3f05dc96 /* (18, 13, 18) */,
  32'h3f05dc96 /* (14, 13, 18) */,
  32'h3e994798 /* (10, 13, 18) */,
  32'h3e2b8c37 /* (6, 13, 18) */,
  32'h3dfd653f /* (2, 13, 18) */,
  32'h3d94a37c /* (30, 9, 18) */,
  32'h3dc45939 /* (26, 9, 18) */,
  32'h3e28e750 /* (22, 9, 18) */,
  32'h3e8dd733 /* (18, 9, 18) */,
  32'h3e8dd733 /* (14, 9, 18) */,
  32'h3e28e750 /* (10, 9, 18) */,
  32'h3dc45939 /* (6, 9, 18) */,
  32'h3d94a37c /* (2, 9, 18) */,
  32'h3d40d8bf /* (30, 5, 18) */,
  32'h3d786cd6 /* (26, 5, 18) */,
  32'h3dce13fe /* (22, 5, 18) */,
  32'h3e27240a /* (18, 5, 18) */,
  32'h3e27240a /* (14, 5, 18) */,
  32'h3dce13fe /* (10, 5, 18) */,
  32'h3d786cd6 /* (6, 5, 18) */,
  32'h3d40d8bf /* (2, 5, 18) */,
  32'h3d217487 /* (30, 1, 18) */,
  32'h3d4cf093 /* (26, 1, 18) */,
  32'h3da6958f /* (22, 1, 18) */,
  32'h3e04a438 /* (18, 1, 18) */,
  32'h3e04a438 /* (14, 1, 18) */,
  32'h3da6958f /* (10, 1, 18) */,
  32'h3d4cf093 /* (6, 1, 18) */,
  32'h3d217487 /* (2, 1, 18) */,
  32'h3d2b1735 /* (30, 29, 14) */,
  32'h3d5a5169 /* (26, 29, 14) */,
  32'h3db2bcb9 /* (22, 29, 14) */,
  32'h3e0f3c67 /* (18, 29, 14) */,
  32'h3e0f3c67 /* (14, 29, 14) */,
  32'h3db2bcb9 /* (10, 29, 14) */,
  32'h3d5a5169 /* (6, 29, 14) */,
  32'h3d2b1735 /* (2, 29, 14) */,
  32'h3d6820b1 /* (30, 25, 14) */,
  32'h3d975464 /* (26, 25, 14) */,
  32'h3dff6ab3 /* (22, 25, 14) */,
  32'h3e528761 /* (18, 25, 14) */,
  32'h3e528761 /* (14, 25, 14) */,
  32'h3dff6ab3 /* (10, 25, 14) */,
  32'h3d975464 /* (6, 25, 14) */,
  32'h3d6820b1 /* (2, 25, 14) */,
  32'h3dc55f41 /* (30, 21, 14) */,
  32'h3e040b60 /* (26, 21, 14) */,
  32'h3e67a191 /* (22, 21, 14) */,
  32'h3ec66134 /* (18, 21, 14) */,
  32'h3ec66134 /* (14, 21, 14) */,
  32'h3e67a191 /* (10, 21, 14) */,
  32'h3e040b60 /* (6, 21, 14) */,
  32'h3dc55f41 /* (2, 21, 14) */,
  32'h3e0adb0d /* (30, 17, 14) */,
  32'h3e3e01e0 /* (26, 17, 14) */,
  32'h3eacaf9b /* (22, 17, 14) */,
  32'h3f19a2a7 /* (18, 17, 14) */,
  32'h3f19a2a7 /* (14, 17, 14) */,
  32'h3eacaf9b /* (10, 17, 14) */,
  32'h3e3e01e0 /* (6, 17, 14) */,
  32'h3e0adb0d /* (2, 17, 14) */,
  32'h3dfd653f /* (30, 13, 14) */,
  32'h3e2b8c37 /* (26, 13, 14) */,
  32'h3e994798 /* (22, 13, 14) */,
  32'h3f05dc96 /* (18, 13, 14) */,
  32'h3f05dc96 /* (14, 13, 14) */,
  32'h3e994798 /* (10, 13, 14) */,
  32'h3e2b8c37 /* (6, 13, 14) */,
  32'h3dfd653f /* (2, 13, 14) */,
  32'h3d94a37c /* (30, 9, 14) */,
  32'h3dc45939 /* (26, 9, 14) */,
  32'h3e28e750 /* (22, 9, 14) */,
  32'h3e8dd733 /* (18, 9, 14) */,
  32'h3e8dd733 /* (14, 9, 14) */,
  32'h3e28e750 /* (10, 9, 14) */,
  32'h3dc45939 /* (6, 9, 14) */,
  32'h3d94a37c /* (2, 9, 14) */,
  32'h3d40d8bf /* (30, 5, 14) */,
  32'h3d786cd6 /* (26, 5, 14) */,
  32'h3dce13fe /* (22, 5, 14) */,
  32'h3e27240a /* (18, 5, 14) */,
  32'h3e27240a /* (14, 5, 14) */,
  32'h3dce13fe /* (10, 5, 14) */,
  32'h3d786cd6 /* (6, 5, 14) */,
  32'h3d40d8bf /* (2, 5, 14) */,
  32'h3d217487 /* (30, 1, 14) */,
  32'h3d4cf093 /* (26, 1, 14) */,
  32'h3da6958f /* (22, 1, 14) */,
  32'h3e04a438 /* (18, 1, 14) */,
  32'h3e04a438 /* (14, 1, 14) */,
  32'h3da6958f /* (10, 1, 14) */,
  32'h3d4cf093 /* (6, 1, 14) */,
  32'h3d217487 /* (2, 1, 14) */,
  32'h3d162b76 /* (30, 29, 10) */,
  32'h3d2c3293 /* (26, 29, 10) */,
  32'h3d77904c /* (22, 29, 10) */,
  32'h3db2bcb9 /* (18, 29, 10) */,
  32'h3db2bcb9 /* (14, 29, 10) */,
  32'h3d77904c /* (10, 29, 10) */,
  32'h3d2c3293 /* (6, 29, 10) */,
  32'h3d162b76 /* (2, 29, 10) */,
  32'h3d3346c6 /* (30, 25, 10) */,
  32'h3d5a2934 /* (26, 25, 10) */,
  32'h3da7f0fb /* (22, 25, 10) */,
  32'h3dff6ab3 /* (18, 25, 10) */,
  32'h3dff6ab3 /* (14, 25, 10) */,
  32'h3da7f0fb /* (10, 25, 10) */,
  32'h3d5a2934 /* (6, 25, 10) */,
  32'h3d3346c6 /* (2, 25, 10) */,
  32'h3d85a0b3 /* (30, 21, 10) */,
  32'h3dac23aa /* (26, 21, 10) */,
  32'h3e0ecbcd /* (22, 21, 10) */,
  32'h3e67a191 /* (18, 21, 10) */,
  32'h3e67a191 /* (14, 21, 10) */,
  32'h3e0ecbcd /* (10, 21, 10) */,
  32'h3dac23aa /* (6, 21, 10) */,
  32'h3d85a0b3 /* (2, 21, 10) */,
  32'h3daa3ec9 /* (30, 17, 10) */,
  32'h3de44bb3 /* (26, 17, 10) */,
  32'h3e48eba4 /* (22, 17, 10) */,
  32'h3eacaf9b /* (18, 17, 10) */,
  32'h3eacaf9b /* (14, 17, 10) */,
  32'h3e48eba4 /* (10, 17, 10) */,
  32'h3de44bb3 /* (6, 17, 10) */,
  32'h3daa3ec9 /* (2, 17, 10) */,
  32'h3da2895a /* (30, 13, 10) */,
  32'h3dd610ea /* (26, 13, 10) */,
  32'h3e37540b /* (22, 13, 10) */,
  32'h3e994798 /* (18, 13, 10) */,
  32'h3e994798 /* (14, 13, 10) */,
  32'h3e37540b /* (10, 13, 10) */,
  32'h3dd610ea /* (6, 13, 10) */,
  32'h3da2895a /* (2, 13, 10) */,
  32'h3d56480e /* (30, 9, 10) */,
  32'h3d866682 /* (26, 9, 10) */,
  32'h3dd7137d /* (22, 9, 10) */,
  32'h3e28e750 /* (18, 9, 10) */,
  32'h3e28e750 /* (14, 9, 10) */,
  32'h3dd7137d /* (10, 9, 10) */,
  32'h3d866682 /* (6, 9, 10) */,
  32'h3d56480e /* (2, 9, 10) */,
  32'h3d1f9f49 /* (30, 5, 10) */,
  32'h3d3c300c /* (26, 5, 10) */,
  32'h3d8b85a2 /* (22, 5, 10) */,
  32'h3dce13fe /* (18, 5, 10) */,
  32'h3dce13fe /* (14, 5, 10) */,
  32'h3d8b85a2 /* (10, 5, 10) */,
  32'h3d3c300c /* (6, 5, 10) */,
  32'h3d1f9f49 /* (2, 5, 10) */,
  32'h3d12ac07 /* (30, 1, 10) */,
  32'h3d2567ce /* (26, 1, 10) */,
  32'h3d699f13 /* (22, 1, 10) */,
  32'h3da6958f /* (18, 1, 10) */,
  32'h3da6958f /* (14, 1, 10) */,
  32'h3d699f13 /* (10, 1, 10) */,
  32'h3d2567ce /* (6, 1, 10) */,
  32'h3d12ac07 /* (2, 1, 10) */,
  32'h3d271e8d /* (30, 29, 6) */,
  32'h3d14c14d /* (26, 29, 6) */,
  32'h3d2c3293 /* (22, 29, 6) */,
  32'h3d5a5169 /* (18, 29, 6) */,
  32'h3d5a5169 /* (14, 29, 6) */,
  32'h3d2c3293 /* (10, 29, 6) */,
  32'h3d14c14d /* (6, 29, 6) */,
  32'h3d271e8d /* (2, 29, 6) */,
  32'h3d14b9d3 /* (30, 25, 6) */,
  32'h3d20f672 /* (26, 25, 6) */,
  32'h3d5a2934 /* (22, 25, 6) */,
  32'h3d975464 /* (18, 25, 6) */,
  32'h3d975464 /* (14, 25, 6) */,
  32'h3d5a2934 /* (10, 25, 6) */,
  32'h3d20f672 /* (6, 25, 6) */,
  32'h3d14b9d3 /* (2, 25, 6) */,
  32'h3d343ccb /* (30, 21, 6) */,
  32'h3d5d3b5c /* (26, 21, 6) */,
  32'h3dac23aa /* (22, 21, 6) */,
  32'h3e040b60 /* (18, 21, 6) */,
  32'h3e040b60 /* (14, 21, 6) */,
  32'h3dac23aa /* (10, 21, 6) */,
  32'h3d5d3b5c /* (6, 21, 6) */,
  32'h3d343ccb /* (2, 21, 6) */,
  32'h3d4bfe66 /* (30, 17, 6) */,
  32'h3d85e8bf /* (26, 17, 6) */,
  32'h3de44bb3 /* (22, 17, 6) */,
  32'h3e3e01e0 /* (18, 17, 6) */,
  32'h3e3e01e0 /* (14, 17, 6) */,
  32'h3de44bb3 /* (10, 17, 6) */,
  32'h3d85e8bf /* (6, 17, 6) */,
  32'h3d4bfe66 /* (2, 17, 6) */,
  32'h3d4ce87b /* (30, 13, 6) */,
  32'h3d82bc35 /* (26, 13, 6) */,
  32'h3dd610ea /* (22, 13, 6) */,
  32'h3e2b8c37 /* (18, 13, 6) */,
  32'h3e2b8c37 /* (14, 13, 6) */,
  32'h3dd610ea /* (10, 13, 6) */,
  32'h3d82bc35 /* (6, 13, 6) */,
  32'h3d4ce87b /* (2, 13, 6) */,
  32'h3d1e19af /* (30, 9, 6) */,
  32'h3d37f9d0 /* (26, 9, 6) */,
  32'h3d866682 /* (22, 9, 6) */,
  32'h3dc45939 /* (18, 9, 6) */,
  32'h3dc45939 /* (14, 9, 6) */,
  32'h3d866682 /* (10, 9, 6) */,
  32'h3d37f9d0 /* (6, 9, 6) */,
  32'h3d1e19af /* (2, 9, 6) */,
  32'h3d18df8d /* (30, 5, 6) */,
  32'h3d16bb8b /* (26, 5, 6) */,
  32'h3d3c300c /* (22, 5, 6) */,
  32'h3d786cd6 /* (18, 5, 6) */,
  32'h3d786cd6 /* (14, 5, 6) */,
  32'h3d3c300c /* (10, 5, 6) */,
  32'h3d16bb8b /* (6, 5, 6) */,
  32'h3d18df8d /* (2, 5, 6) */,
  32'h3d3543e4 /* (30, 1, 6) */,
  32'h3d15cc97 /* (26, 1, 6) */,
  32'h3d2567ce /* (22, 1, 6) */,
  32'h3d4cf093 /* (18, 1, 6) */,
  32'h3d4cf093 /* (14, 1, 6) */,
  32'h3d2567ce /* (10, 1, 6) */,
  32'h3d15cc97 /* (6, 1, 6) */,
  32'h3d3543e4 /* (2, 1, 6) */,
  32'h3da3af74 /* (30, 29, 2) */,
  32'h3d271e8d /* (26, 29, 2) */,
  32'h3d162b76 /* (22, 29, 2) */,
  32'h3d2b1735 /* (18, 29, 2) */,
  32'h3d2b1735 /* (14, 29, 2) */,
  32'h3d162b76 /* (10, 29, 2) */,
  32'h3d271e8d /* (6, 29, 2) */,
  32'h3da3af74 /* (2, 29, 2) */,
  32'h3d1dd271 /* (30, 25, 2) */,
  32'h3d14b9d3 /* (26, 25, 2) */,
  32'h3d3346c6 /* (22, 25, 2) */,
  32'h3d6820b1 /* (18, 25, 2) */,
  32'h3d6820b1 /* (14, 25, 2) */,
  32'h3d3346c6 /* (10, 25, 2) */,
  32'h3d14b9d3 /* (6, 25, 2) */,
  32'h3d1dd271 /* (2, 25, 2) */,
  32'h3d18e0f8 /* (30, 21, 2) */,
  32'h3d343ccb /* (26, 21, 2) */,
  32'h3d85a0b3 /* (22, 21, 2) */,
  32'h3dc55f41 /* (18, 21, 2) */,
  32'h3dc55f41 /* (14, 21, 2) */,
  32'h3d85a0b3 /* (10, 21, 2) */,
  32'h3d343ccb /* (6, 21, 2) */,
  32'h3d18e0f8 /* (2, 21, 2) */,
  32'h3d1dadb9 /* (30, 17, 2) */,
  32'h3d4bfe66 /* (26, 17, 2) */,
  32'h3daa3ec9 /* (22, 17, 2) */,
  32'h3e0adb0d /* (18, 17, 2) */,
  32'h3e0adb0d /* (14, 17, 2) */,
  32'h3daa3ec9 /* (10, 17, 2) */,
  32'h3d4bfe66 /* (6, 17, 2) */,
  32'h3d1dadb9 /* (2, 17, 2) */,
  32'h3d246fbd /* (30, 13, 2) */,
  32'h3d4ce87b /* (26, 13, 2) */,
  32'h3da2895a /* (22, 13, 2) */,
  32'h3dfd653f /* (18, 13, 2) */,
  32'h3dfd653f /* (14, 13, 2) */,
  32'h3da2895a /* (10, 13, 2) */,
  32'h3d4ce87b /* (6, 13, 2) */,
  32'h3d246fbd /* (2, 13, 2) */,
  32'h3d1214c5 /* (30, 9, 2) */,
  32'h3d1e19af /* (26, 9, 2) */,
  32'h3d56480e /* (22, 9, 2) */,
  32'h3d94a37c /* (18, 9, 2) */,
  32'h3d94a37c /* (14, 9, 2) */,
  32'h3d56480e /* (10, 9, 2) */,
  32'h3d1e19af /* (6, 9, 2) */,
  32'h3d1214c5 /* (2, 9, 2) */,
  32'h3d4ca49b /* (30, 5, 2) */,
  32'h3d18df8d /* (26, 5, 2) */,
  32'h3d1f9f49 /* (22, 5, 2) */,
  32'h3d40d8bf /* (18, 5, 2) */,
  32'h3d40d8bf /* (14, 5, 2) */,
  32'h3d1f9f49 /* (10, 5, 2) */,
  32'h3d18df8d /* (6, 5, 2) */,
  32'h3d4ca49b /* (2, 5, 2) */,
  32'h3e0c4d23 /* (30, 1, 2) */,
  32'h3d3543e4 /* (26, 1, 2) */,
  32'h3d12ac07 /* (22, 1, 2) */,
  32'h3d217487 /* (18, 1, 2) */,
  32'h3d217487 /* (14, 1, 2) */,
  32'h3d12ac07 /* (10, 1, 2) */,
  32'h3d3543e4 /* (6, 1, 2) */,
  32'h3e0c4d23 /* (2, 1, 2) */,
  32'h3d866355 /* (29, 29, 30) */,
  32'h3d1a2949 /* (25, 29, 30) */,
  32'h3d1c5f03 /* (21, 29, 30) */,
  32'h3d240321 /* (17, 29, 30) */,
  32'h3d29e985 /* (13, 29, 30) */,
  32'h3d12f42a /* (9, 29, 30) */,
  32'h3d3cd255 /* (5, 29, 30) */,
  32'h3dbfa8df /* (1, 29, 30) */,
  32'h3d1a2949 /* (29, 25, 30) */,
  32'h3d1777c7 /* (25, 25, 30) */,
  32'h3d42a7b8 /* (21, 25, 30) */,
  32'h3d62f778 /* (17, 25, 30) */,
  32'h3d6129ae /* (13, 25, 30) */,
  32'h3d26a1b5 /* (9, 25, 30) */,
  32'h3d14b1c0 /* (5, 25, 30) */,
  32'h3d20a35e /* (1, 25, 30) */,
  32'h3d1c5f03 /* (29, 21, 30) */,
  32'h3d42a7b8 /* (25, 21, 30) */,
  32'h3d96eb50 /* (21, 21, 30) */,
  32'h3dc59b81 /* (17, 21, 30) */,
  32'h3dba5db4 /* (13, 21, 30) */,
  32'h3d6d9fa3 /* (9, 21, 30) */,
  32'h3d29823f /* (5, 21, 30) */,
  32'h3d16ed42 /* (1, 21, 30) */,
  32'h3d240321 /* (29, 17, 30) */,
  32'h3d62f778 /* (25, 17, 30) */,
  32'h3dc59b81 /* (21, 17, 30) */,
  32'h3e0de5f8 /* (17, 17, 30) */,
  32'h3e003b1e /* (13, 17, 30) */,
  32'h3d9314c2 /* (9, 17, 30) */,
  32'h3d3a7be5 /* (5, 17, 30) */,
  32'h3d1a0745 /* (1, 17, 30) */,
  32'h3d29e985 /* (29, 13, 30) */,
  32'h3d6129ae /* (25, 13, 30) */,
  32'h3dba5db4 /* (21, 13, 30) */,
  32'h3e003b1e /* (17, 13, 30) */,
  32'h3dec70da /* (13, 13, 30) */,
  32'h3d8e358b /* (9, 13, 30) */,
  32'h3d3d84de /* (5, 13, 30) */,
  32'h3d214ba3 /* (1, 13, 30) */,
  32'h3d12f42a /* (29, 9, 30) */,
  32'h3d26a1b5 /* (25, 9, 30) */,
  32'h3d6d9fa3 /* (21, 9, 30) */,
  32'h3d9314c2 /* (17, 9, 30) */,
  32'h3d8e358b /* (13, 9, 30) */,
  32'h3d42665b /* (9, 9, 30) */,
  32'h3d18622e /* (5, 9, 30) */,
  32'h3d11c69f /* (1, 9, 30) */,
  32'h3d3cd255 /* (29, 5, 30) */,
  32'h3d14b1c0 /* (25, 5, 30) */,
  32'h3d29823f /* (21, 5, 30) */,
  32'h3d3a7be5 /* (17, 5, 30) */,
  32'h3d3d84de /* (13, 5, 30) */,
  32'h3d18622e /* (9, 5, 30) */,
  32'h3d213c91 /* (5, 5, 30) */,
  32'h3d59109a /* (1, 5, 30) */,
  32'h3dbfa8df /* (29, 1, 30) */,
  32'h3d20a35e /* (25, 1, 30) */,
  32'h3d16ed42 /* (21, 1, 30) */,
  32'h3d1a0745 /* (17, 1, 30) */,
  32'h3d214ba3 /* (13, 1, 30) */,
  32'h3d11c69f /* (9, 1, 30) */,
  32'h3d59109a /* (5, 1, 30) */,
  32'h3e4aeee2 /* (1, 1, 30) */,
  32'h3d211f1b /* (29, 29, 26) */,
  32'h3d159d44 /* (25, 29, 26) */,
  32'h3d39bb76 /* (21, 29, 26) */,
  32'h3d54ba37 /* (17, 29, 26) */,
  32'h3d54a03b /* (13, 29, 26) */,
  32'h3d215063 /* (9, 29, 26) */,
  32'h3d16d305 /* (5, 29, 26) */,
  32'h3d2ba889 /* (1, 29, 26) */,
  32'h3d159d44 /* (29, 25, 26) */,
  32'h3d29a602 /* (25, 25, 26) */,
  32'h3d71ecf9 /* (21, 25, 26) */,
  32'h3d95be73 /* (17, 25, 26) */,
  32'h3d90c8a7 /* (13, 25, 26) */,
  32'h3d45eb5b /* (9, 25, 26) */,
  32'h3d1b2471 /* (5, 25, 26) */,
  32'h3d146a43 /* (1, 25, 26) */,
  32'h3d39bb76 /* (29, 21, 26) */,
  32'h3d71ecf9 /* (25, 21, 26) */,
  32'h3dc480ba /* (21, 21, 26) */,
  32'h3e0533d0 /* (17, 21, 26) */,
  32'h3df74dbc /* (13, 21, 26) */,
  32'h3d9750ce /* (9, 21, 26) */,
  32'h3d4d9045 /* (5, 21, 26) */,
  32'h3d31191b /* (1, 21, 26) */,
  32'h3d54ba37 /* (29, 17, 26) */,
  32'h3d95be73 /* (25, 17, 26) */,
  32'h3e0533d0 /* (21, 17, 26) */,
  32'h3e430b11 /* (17, 17, 26) */,
  32'h3e2ea39a /* (13, 17, 26) */,
  32'h3dc42ad0 /* (9, 17, 26) */,
  32'h3d73b16f /* (5, 17, 26) */,
  32'h3d46f53f /* (1, 17, 26) */,
  32'h3d54a03b /* (29, 13, 26) */,
  32'h3d90c8a7 /* (25, 13, 26) */,
  32'h3df74dbc /* (21, 13, 26) */,
  32'h3e2ea39a /* (17, 13, 26) */,
  32'h3e1f113d /* (13, 13, 26) */,
  32'h3db9d5f4 /* (9, 13, 26) */,
  32'h3d700ffa /* (5, 13, 26) */,
  32'h3d4876ff /* (1, 13, 26) */,
  32'h3d215063 /* (29, 9, 26) */,
  32'h3d45eb5b /* (25, 9, 26) */,
  32'h3d9750ce /* (21, 9, 26) */,
  32'h3dc42ad0 /* (17, 9, 26) */,
  32'h3db9d5f4 /* (13, 9, 26) */,
  32'h3d6fd024 /* (9, 9, 26) */,
  32'h3d2db0cc /* (5, 9, 26) */,
  32'h3d1c53e8 /* (1, 9, 26) */,
  32'h3d16d305 /* (29, 5, 26) */,
  32'h3d1b2471 /* (25, 5, 26) */,
  32'h3d4d9045 /* (21, 5, 26) */,
  32'h3d73b16f /* (17, 5, 26) */,
  32'h3d700ffa /* (13, 5, 26) */,
  32'h3d2db0cc /* (9, 5, 26) */,
  32'h3d14f7ce /* (5, 5, 26) */,
  32'h3d1a8b5a /* (1, 5, 26) */,
  32'h3d2ba889 /* (29, 1, 26) */,
  32'h3d146a43 /* (25, 1, 26) */,
  32'h3d31191b /* (21, 1, 26) */,
  32'h3d46f53f /* (17, 1, 26) */,
  32'h3d4876ff /* (13, 1, 26) */,
  32'h3d1c53e8 /* (9, 1, 26) */,
  32'h3d1a8b5a /* (5, 1, 26) */,
  32'h3d3c9698 /* (1, 1, 26) */,
  32'h3d18cb02 /* (29, 29, 22) */,
  32'h3d387393 /* (25, 29, 22) */,
  32'h3d8ae43c /* (21, 29, 22) */,
  32'h3db22d06 /* (17, 29, 22) */,
  32'h3da99659 /* (13, 29, 22) */,
  32'h3d5dae2c /* (9, 29, 22) */,
  32'h3d2344c4 /* (5, 29, 22) */,
  32'h3d14c0fd /* (1, 29, 22) */,
  32'h3d387393 /* (29, 25, 22) */,
  32'h3d6deb12 /* (25, 25, 22) */,
  32'h3dbf3f1d /* (21, 25, 22) */,
  32'h3e009a19 /* (17, 25, 22) */,
  32'h3defa49b /* (13, 25, 22) */,
  32'h3d94014f /* (9, 25, 22) */,
  32'h3d4b3dc7 /* (5, 25, 22) */,
  32'h3d305430 /* (1, 25, 22) */,
  32'h3d8ae43c /* (29, 21, 22) */,
  32'h3dbf3f1d /* (25, 21, 22) */,
  32'h3e257fc6 /* (21, 21, 22) */,
  32'h3e6c6ac0 /* (17, 21, 22) */,
  32'h3e562fb1 /* (13, 21, 22) */,
  32'h3df71c69 /* (9, 21, 22) */,
  32'h3d9d9380 /* (5, 21, 22) */,
  32'h3d829849 /* (1, 21, 22) */,
  32'h3db22d06 /* (29, 17, 22) */,
  32'h3e009a19 /* (25, 17, 22) */,
  32'h3e6c6ac0 /* (21, 17, 22) */,
  32'h3eb2925b /* (17, 17, 22) */,
  32'h3e9d80fb /* (13, 17, 22) */,
  32'h3e2b3653 /* (9, 17, 22) */,
  32'h3dce52e6 /* (5, 17, 22) */,
  32'h3da5ac70 /* (1, 17, 22) */,
  32'h3da99659 /* (29, 13, 22) */,
  32'h3defa49b /* (25, 13, 22) */,
  32'h3e562fb1 /* (21, 13, 22) */,
  32'h3e9d80fb /* (17, 13, 22) */,
  32'h3e8cbae1 /* (13, 13, 22) */,
  32'h3e1d56b2 /* (9, 13, 22) */,
  32'h3dc29629 /* (5, 13, 22) */,
  32'h3d9e7894 /* (1, 13, 22) */,
  32'h3d5dae2c /* (29, 9, 22) */,
  32'h3d94014f /* (25, 9, 22) */,
  32'h3df71c69 /* (21, 9, 22) */,
  32'h3e2b3653 /* (17, 9, 22) */,
  32'h3e1d56b2 /* (13, 9, 22) */,
  32'h3dbbc730 /* (9, 9, 22) */,
  32'h3d781ae6 /* (5, 9, 22) */,
  32'h3d52081f /* (1, 9, 22) */,
  32'h3d2344c4 /* (29, 5, 22) */,
  32'h3d4b3dc7 /* (25, 5, 22) */,
  32'h3d9d9380 /* (21, 5, 22) */,
  32'h3dce52e6 /* (17, 5, 22) */,
  32'h3dc29629 /* (13, 5, 22) */,
  32'h3d781ae6 /* (9, 5, 22) */,
  32'h3d30fc5a /* (5, 5, 22) */,
  32'h3d1d9589 /* (1, 5, 22) */,
  32'h3d14c0fd /* (29, 1, 22) */,
  32'h3d305430 /* (25, 1, 22) */,
  32'h3d829849 /* (21, 1, 22) */,
  32'h3da5ac70 /* (17, 1, 22) */,
  32'h3d9e7894 /* (13, 1, 22) */,
  32'h3d52081f /* (9, 1, 22) */,
  32'h3d1d9589 /* (5, 1, 22) */,
  32'h3d119771 /* (1, 1, 22) */,
  32'h3d3188e3 /* (29, 29, 18) */,
  32'h3d71c736 /* (25, 29, 18) */,
  32'h3dce7d45 /* (21, 29, 18) */,
  32'h3e11d12f /* (17, 29, 18) */,
  32'h3e04d0b8 /* (13, 29, 18) */,
  32'h3d9b2a7b /* (9, 29, 18) */,
  32'h3d487174 /* (5, 29, 18) */,
  32'h3d276174 /* (1, 29, 18) */,
  32'h3d71c736 /* (29, 25, 18) */,
  32'h3da8d240 /* (25, 25, 18) */,
  32'h3e14a5c9 /* (21, 25, 18) */,
  32'h3e57a44b /* (17, 25, 18) */,
  32'h3e41f14c /* (13, 25, 18) */,
  32'h3ddc09d8 /* (9, 25, 18) */,
  32'h3d8a0000 /* (5, 25, 18) */,
  32'h3d62906c /* (1, 25, 18) */,
  32'h3dce7d45 /* (29, 21, 18) */,
  32'h3e14a5c9 /* (25, 21, 18) */,
  32'h3e882756 /* (21, 21, 18) */,
  32'h3eccf8ff /* (17, 21, 18) */,
  32'h3eb517ce /* (13, 21, 18) */,
  32'h3e458f30 /* (9, 21, 18) */,
  32'h3deed79f /* (5, 21, 18) */,
  32'h3dc01db4 /* (1, 21, 18) */,
  32'h3e11d12f /* (29, 17, 18) */,
  32'h3e57a44b /* (25, 17, 18) */,
  32'h3eccf8ff /* (21, 17, 18) */,
  32'h3f202f9a /* (17, 17, 18) */,
  32'h3f0af24f /* (13, 17, 18) */,
  32'h3e91e4f8 /* (9, 17, 18) */,
  32'h3e2a981c /* (5, 17, 18) */,
  32'h3e06d8bb /* (1, 17, 18) */,
  32'h3e04d0b8 /* (29, 13, 18) */,
  32'h3e41f14c /* (25, 13, 18) */,
  32'h3eb517ce /* (21, 13, 18) */,
  32'h3f0af24f /* (17, 13, 18) */,
  32'h3ef33ce4 /* (13, 13, 18) */,
  32'h3e821787 /* (9, 13, 18) */,
  32'h3e1a8d8c /* (5, 13, 18) */,
  32'h3df65860 /* (1, 13, 18) */,
  32'h3d9b2a7b /* (29, 9, 18) */,
  32'h3ddc09d8 /* (25, 9, 18) */,
  32'h3e458f30 /* (21, 9, 18) */,
  32'h3e91e4f8 /* (17, 9, 18) */,
  32'h3e821787 /* (13, 9, 18) */,
  32'h3e10cac5 /* (9, 9, 18) */,
  32'h3db24f8e /* (5, 9, 18) */,
  32'h3d90dff9 /* (1, 9, 18) */,
  32'h3d487174 /* (29, 5, 18) */,
  32'h3d8a0000 /* (25, 5, 18) */,
  32'h3deed79f /* (21, 5, 18) */,
  32'h3e2a981c /* (17, 5, 18) */,
  32'h3e1a8d8c /* (13, 5, 18) */,
  32'h3db24f8e /* (9, 5, 18) */,
  32'h3d63687e /* (5, 5, 18) */,
  32'h3d3c7841 /* (1, 5, 18) */,
  32'h3d276174 /* (29, 1, 18) */,
  32'h3d62906c /* (25, 1, 18) */,
  32'h3dc01db4 /* (21, 1, 18) */,
  32'h3e06d8bb /* (17, 1, 18) */,
  32'h3df65860 /* (13, 1, 18) */,
  32'h3d90dff9 /* (9, 1, 18) */,
  32'h3d3c7841 /* (5, 1, 18) */,
  32'h3d1e0bb6 /* (1, 1, 18) */,
  32'h3d3188e3 /* (29, 29, 14) */,
  32'h3d71c736 /* (25, 29, 14) */,
  32'h3dce7d45 /* (21, 29, 14) */,
  32'h3e11d12f /* (17, 29, 14) */,
  32'h3e04d0b8 /* (13, 29, 14) */,
  32'h3d9b2a7b /* (9, 29, 14) */,
  32'h3d487174 /* (5, 29, 14) */,
  32'h3d276174 /* (1, 29, 14) */,
  32'h3d71c736 /* (29, 25, 14) */,
  32'h3da8d240 /* (25, 25, 14) */,
  32'h3e14a5c9 /* (21, 25, 14) */,
  32'h3e57a44b /* (17, 25, 14) */,
  32'h3e41f14c /* (13, 25, 14) */,
  32'h3ddc09d8 /* (9, 25, 14) */,
  32'h3d8a0000 /* (5, 25, 14) */,
  32'h3d62906c /* (1, 25, 14) */,
  32'h3dce7d45 /* (29, 21, 14) */,
  32'h3e14a5c9 /* (25, 21, 14) */,
  32'h3e882756 /* (21, 21, 14) */,
  32'h3eccf8ff /* (17, 21, 14) */,
  32'h3eb517ce /* (13, 21, 14) */,
  32'h3e458f30 /* (9, 21, 14) */,
  32'h3deed79f /* (5, 21, 14) */,
  32'h3dc01db4 /* (1, 21, 14) */,
  32'h3e11d12f /* (29, 17, 14) */,
  32'h3e57a44b /* (25, 17, 14) */,
  32'h3eccf8ff /* (21, 17, 14) */,
  32'h3f202f9a /* (17, 17, 14) */,
  32'h3f0af24f /* (13, 17, 14) */,
  32'h3e91e4f8 /* (9, 17, 14) */,
  32'h3e2a981c /* (5, 17, 14) */,
  32'h3e06d8bb /* (1, 17, 14) */,
  32'h3e04d0b8 /* (29, 13, 14) */,
  32'h3e41f14c /* (25, 13, 14) */,
  32'h3eb517ce /* (21, 13, 14) */,
  32'h3f0af24f /* (17, 13, 14) */,
  32'h3ef33ce4 /* (13, 13, 14) */,
  32'h3e821787 /* (9, 13, 14) */,
  32'h3e1a8d8c /* (5, 13, 14) */,
  32'h3df65860 /* (1, 13, 14) */,
  32'h3d9b2a7b /* (29, 9, 14) */,
  32'h3ddc09d8 /* (25, 9, 14) */,
  32'h3e458f30 /* (21, 9, 14) */,
  32'h3e91e4f8 /* (17, 9, 14) */,
  32'h3e821787 /* (13, 9, 14) */,
  32'h3e10cac5 /* (9, 9, 14) */,
  32'h3db24f8e /* (5, 9, 14) */,
  32'h3d90dff9 /* (1, 9, 14) */,
  32'h3d487174 /* (29, 5, 14) */,
  32'h3d8a0000 /* (25, 5, 14) */,
  32'h3deed79f /* (21, 5, 14) */,
  32'h3e2a981c /* (17, 5, 14) */,
  32'h3e1a8d8c /* (13, 5, 14) */,
  32'h3db24f8e /* (9, 5, 14) */,
  32'h3d63687e /* (5, 5, 14) */,
  32'h3d3c7841 /* (1, 5, 14) */,
  32'h3d276174 /* (29, 1, 14) */,
  32'h3d62906c /* (25, 1, 14) */,
  32'h3dc01db4 /* (21, 1, 14) */,
  32'h3e06d8bb /* (17, 1, 14) */,
  32'h3df65860 /* (13, 1, 14) */,
  32'h3d90dff9 /* (9, 1, 14) */,
  32'h3d3c7841 /* (5, 1, 14) */,
  32'h3d1e0bb6 /* (1, 1, 14) */,
  32'h3d18cb02 /* (29, 29, 10) */,
  32'h3d387393 /* (25, 29, 10) */,
  32'h3d8ae43c /* (21, 29, 10) */,
  32'h3db22d06 /* (17, 29, 10) */,
  32'h3da99659 /* (13, 29, 10) */,
  32'h3d5dae2c /* (9, 29, 10) */,
  32'h3d2344c4 /* (5, 29, 10) */,
  32'h3d14c0fd /* (1, 29, 10) */,
  32'h3d387393 /* (29, 25, 10) */,
  32'h3d6deb12 /* (25, 25, 10) */,
  32'h3dbf3f1d /* (21, 25, 10) */,
  32'h3e009a19 /* (17, 25, 10) */,
  32'h3defa49b /* (13, 25, 10) */,
  32'h3d94014f /* (9, 25, 10) */,
  32'h3d4b3dc7 /* (5, 25, 10) */,
  32'h3d305430 /* (1, 25, 10) */,
  32'h3d8ae43c /* (29, 21, 10) */,
  32'h3dbf3f1d /* (25, 21, 10) */,
  32'h3e257fc6 /* (21, 21, 10) */,
  32'h3e6c6ac0 /* (17, 21, 10) */,
  32'h3e562fb1 /* (13, 21, 10) */,
  32'h3df71c69 /* (9, 21, 10) */,
  32'h3d9d9380 /* (5, 21, 10) */,
  32'h3d829849 /* (1, 21, 10) */,
  32'h3db22d06 /* (29, 17, 10) */,
  32'h3e009a19 /* (25, 17, 10) */,
  32'h3e6c6ac0 /* (21, 17, 10) */,
  32'h3eb2925b /* (17, 17, 10) */,
  32'h3e9d80fb /* (13, 17, 10) */,
  32'h3e2b3653 /* (9, 17, 10) */,
  32'h3dce52e6 /* (5, 17, 10) */,
  32'h3da5ac70 /* (1, 17, 10) */,
  32'h3da99659 /* (29, 13, 10) */,
  32'h3defa49b /* (25, 13, 10) */,
  32'h3e562fb1 /* (21, 13, 10) */,
  32'h3e9d80fb /* (17, 13, 10) */,
  32'h3e8cbae1 /* (13, 13, 10) */,
  32'h3e1d56b2 /* (9, 13, 10) */,
  32'h3dc29629 /* (5, 13, 10) */,
  32'h3d9e7894 /* (1, 13, 10) */,
  32'h3d5dae2c /* (29, 9, 10) */,
  32'h3d94014f /* (25, 9, 10) */,
  32'h3df71c69 /* (21, 9, 10) */,
  32'h3e2b3653 /* (17, 9, 10) */,
  32'h3e1d56b2 /* (13, 9, 10) */,
  32'h3dbbc730 /* (9, 9, 10) */,
  32'h3d781ae6 /* (5, 9, 10) */,
  32'h3d52081f /* (1, 9, 10) */,
  32'h3d2344c4 /* (29, 5, 10) */,
  32'h3d4b3dc7 /* (25, 5, 10) */,
  32'h3d9d9380 /* (21, 5, 10) */,
  32'h3dce52e6 /* (17, 5, 10) */,
  32'h3dc29629 /* (13, 5, 10) */,
  32'h3d781ae6 /* (9, 5, 10) */,
  32'h3d30fc5a /* (5, 5, 10) */,
  32'h3d1d9589 /* (1, 5, 10) */,
  32'h3d14c0fd /* (29, 1, 10) */,
  32'h3d305430 /* (25, 1, 10) */,
  32'h3d829849 /* (21, 1, 10) */,
  32'h3da5ac70 /* (17, 1, 10) */,
  32'h3d9e7894 /* (13, 1, 10) */,
  32'h3d52081f /* (9, 1, 10) */,
  32'h3d1d9589 /* (5, 1, 10) */,
  32'h3d119771 /* (1, 1, 10) */,
  32'h3d211f1b /* (29, 29, 6) */,
  32'h3d159d44 /* (25, 29, 6) */,
  32'h3d39bb76 /* (21, 29, 6) */,
  32'h3d54ba37 /* (17, 29, 6) */,
  32'h3d54a03b /* (13, 29, 6) */,
  32'h3d215063 /* (9, 29, 6) */,
  32'h3d16d305 /* (5, 29, 6) */,
  32'h3d2ba889 /* (1, 29, 6) */,
  32'h3d159d44 /* (29, 25, 6) */,
  32'h3d29a602 /* (25, 25, 6) */,
  32'h3d71ecf9 /* (21, 25, 6) */,
  32'h3d95be73 /* (17, 25, 6) */,
  32'h3d90c8a7 /* (13, 25, 6) */,
  32'h3d45eb5b /* (9, 25, 6) */,
  32'h3d1b2471 /* (5, 25, 6) */,
  32'h3d146a43 /* (1, 25, 6) */,
  32'h3d39bb76 /* (29, 21, 6) */,
  32'h3d71ecf9 /* (25, 21, 6) */,
  32'h3dc480ba /* (21, 21, 6) */,
  32'h3e0533d0 /* (17, 21, 6) */,
  32'h3df74dbc /* (13, 21, 6) */,
  32'h3d9750ce /* (9, 21, 6) */,
  32'h3d4d9045 /* (5, 21, 6) */,
  32'h3d31191b /* (1, 21, 6) */,
  32'h3d54ba37 /* (29, 17, 6) */,
  32'h3d95be73 /* (25, 17, 6) */,
  32'h3e0533d0 /* (21, 17, 6) */,
  32'h3e430b11 /* (17, 17, 6) */,
  32'h3e2ea39a /* (13, 17, 6) */,
  32'h3dc42ad0 /* (9, 17, 6) */,
  32'h3d73b16f /* (5, 17, 6) */,
  32'h3d46f53f /* (1, 17, 6) */,
  32'h3d54a03b /* (29, 13, 6) */,
  32'h3d90c8a7 /* (25, 13, 6) */,
  32'h3df74dbc /* (21, 13, 6) */,
  32'h3e2ea39a /* (17, 13, 6) */,
  32'h3e1f113d /* (13, 13, 6) */,
  32'h3db9d5f4 /* (9, 13, 6) */,
  32'h3d700ffa /* (5, 13, 6) */,
  32'h3d4876ff /* (1, 13, 6) */,
  32'h3d215063 /* (29, 9, 6) */,
  32'h3d45eb5b /* (25, 9, 6) */,
  32'h3d9750ce /* (21, 9, 6) */,
  32'h3dc42ad0 /* (17, 9, 6) */,
  32'h3db9d5f4 /* (13, 9, 6) */,
  32'h3d6fd024 /* (9, 9, 6) */,
  32'h3d2db0cc /* (5, 9, 6) */,
  32'h3d1c53e8 /* (1, 9, 6) */,
  32'h3d16d305 /* (29, 5, 6) */,
  32'h3d1b2471 /* (25, 5, 6) */,
  32'h3d4d9045 /* (21, 5, 6) */,
  32'h3d73b16f /* (17, 5, 6) */,
  32'h3d700ffa /* (13, 5, 6) */,
  32'h3d2db0cc /* (9, 5, 6) */,
  32'h3d14f7ce /* (5, 5, 6) */,
  32'h3d1a8b5a /* (1, 5, 6) */,
  32'h3d2ba889 /* (29, 1, 6) */,
  32'h3d146a43 /* (25, 1, 6) */,
  32'h3d31191b /* (21, 1, 6) */,
  32'h3d46f53f /* (17, 1, 6) */,
  32'h3d4876ff /* (13, 1, 6) */,
  32'h3d1c53e8 /* (9, 1, 6) */,
  32'h3d1a8b5a /* (5, 1, 6) */,
  32'h3d3c9698 /* (1, 1, 6) */,
  32'h3d866355 /* (29, 29, 2) */,
  32'h3d1a2949 /* (25, 29, 2) */,
  32'h3d1c5f03 /* (21, 29, 2) */,
  32'h3d240321 /* (17, 29, 2) */,
  32'h3d29e985 /* (13, 29, 2) */,
  32'h3d12f42a /* (9, 29, 2) */,
  32'h3d3cd255 /* (5, 29, 2) */,
  32'h3dbfa8df /* (1, 29, 2) */,
  32'h3d1a2949 /* (29, 25, 2) */,
  32'h3d1777c7 /* (25, 25, 2) */,
  32'h3d42a7b8 /* (21, 25, 2) */,
  32'h3d62f778 /* (17, 25, 2) */,
  32'h3d6129ae /* (13, 25, 2) */,
  32'h3d26a1b5 /* (9, 25, 2) */,
  32'h3d14b1c0 /* (5, 25, 2) */,
  32'h3d20a35e /* (1, 25, 2) */,
  32'h3d1c5f03 /* (29, 21, 2) */,
  32'h3d42a7b8 /* (25, 21, 2) */,
  32'h3d96eb50 /* (21, 21, 2) */,
  32'h3dc59b81 /* (17, 21, 2) */,
  32'h3dba5db4 /* (13, 21, 2) */,
  32'h3d6d9fa3 /* (9, 21, 2) */,
  32'h3d29823f /* (5, 21, 2) */,
  32'h3d16ed42 /* (1, 21, 2) */,
  32'h3d240321 /* (29, 17, 2) */,
  32'h3d62f778 /* (25, 17, 2) */,
  32'h3dc59b81 /* (21, 17, 2) */,
  32'h3e0de5f8 /* (17, 17, 2) */,
  32'h3e003b1e /* (13, 17, 2) */,
  32'h3d9314c2 /* (9, 17, 2) */,
  32'h3d3a7be5 /* (5, 17, 2) */,
  32'h3d1a0745 /* (1, 17, 2) */,
  32'h3d29e985 /* (29, 13, 2) */,
  32'h3d6129ae /* (25, 13, 2) */,
  32'h3dba5db4 /* (21, 13, 2) */,
  32'h3e003b1e /* (17, 13, 2) */,
  32'h3dec70da /* (13, 13, 2) */,
  32'h3d8e358b /* (9, 13, 2) */,
  32'h3d3d84de /* (5, 13, 2) */,
  32'h3d214ba3 /* (1, 13, 2) */,
  32'h3d12f42a /* (29, 9, 2) */,
  32'h3d26a1b5 /* (25, 9, 2) */,
  32'h3d6d9fa3 /* (21, 9, 2) */,
  32'h3d9314c2 /* (17, 9, 2) */,
  32'h3d8e358b /* (13, 9, 2) */,
  32'h3d42665b /* (9, 9, 2) */,
  32'h3d18622e /* (5, 9, 2) */,
  32'h3d11c69f /* (1, 9, 2) */,
  32'h3d3cd255 /* (29, 5, 2) */,
  32'h3d14b1c0 /* (25, 5, 2) */,
  32'h3d29823f /* (21, 5, 2) */,
  32'h3d3a7be5 /* (17, 5, 2) */,
  32'h3d3d84de /* (13, 5, 2) */,
  32'h3d18622e /* (9, 5, 2) */,
  32'h3d213c91 /* (5, 5, 2) */,
  32'h3d59109a /* (1, 5, 2) */,
  32'h3dbfa8df /* (29, 1, 2) */,
  32'h3d20a35e /* (25, 1, 2) */,
  32'h3d16ed42 /* (21, 1, 2) */,
  32'h3d1a0745 /* (17, 1, 2) */,
  32'h3d214ba3 /* (13, 1, 2) */,
  32'h3d11c69f /* (9, 1, 2) */,
  32'h3d59109a /* (5, 1, 2) */,
  32'h3e4aeee2 /* (1, 1, 2) */,
  32'h3d5defd3 /* (28, 29, 30) */,
  32'h3d13e9f7 /* (24, 29, 30) */,
  32'h3d23d587 /* (20, 29, 30) */,
  32'h3d13661d /* (16, 29, 30) */,
  32'h3d23d587 /* (12, 29, 30) */,
  32'h3d13e9f7 /* (8, 29, 30) */,
  32'h3d5defd3 /* (4, 29, 30) */,
  32'h3dcbea25 /* (0, 29, 30) */,
  32'h3d16c6a3 /* (28, 25, 30) */,
  32'h3d1d59b0 /* (24, 25, 30) */,
  32'h3d530d8e /* (20, 25, 30) */,
  32'h3d4f6a6e /* (16, 25, 30) */,
  32'h3d530d8e /* (12, 25, 30) */,
  32'h3d1d59b0 /* (8, 25, 30) */,
  32'h3d16c6a3 /* (4, 25, 30) */,
  32'h3d21b235 /* (0, 25, 30) */,
  32'h3d21c128 /* (28, 21, 30) */,
  32'h3d558b1c /* (24, 21, 30) */,
  32'h3da96c08 /* (20, 21, 30) */,
  32'h3db86416 /* (16, 21, 30) */,
  32'h3da96c08 /* (12, 21, 30) */,
  32'h3d558b1c /* (8, 21, 30) */,
  32'h3d21c128 /* (4, 21, 30) */,
  32'h3d164ce1 /* (0, 21, 30) */,
  32'h3d2d6bba /* (28, 17, 30) */,
  32'h3d804df8 /* (24, 17, 30) */,
  32'h3de39dff /* (20, 17, 30) */,
  32'h3e06ec2e /* (16, 17, 30) */,
  32'h3de39dff /* (12, 17, 30) */,
  32'h3d804df8 /* (8, 17, 30) */,
  32'h3d2d6bba /* (4, 17, 30) */,
  32'h3d18d610 /* (0, 17, 30) */,
  32'h3d3217f4 /* (28, 13, 30) */,
  32'h3d7b52f8 /* (24, 13, 30) */,
  32'h3dd42d31 /* (20, 13, 30) */,
  32'h3df1ae3d /* (16, 13, 30) */,
  32'h3dd42d31 /* (12, 13, 30) */,
  32'h3d7b52f8 /* (8, 13, 30) */,
  32'h3d3217f4 /* (4, 13, 30) */,
  32'h3d2045b1 /* (0, 13, 30) */,
  32'h3d14de35 /* (28, 9, 30) */,
  32'h3d3291f6 /* (24, 9, 30) */,
  32'h3d833332 /* (20, 9, 30) */,
  32'h3d87d16b /* (16, 9, 30) */,
  32'h3d833332 /* (12, 9, 30) */,
  32'h3d3291f6 /* (8, 9, 30) */,
  32'h3d14de35 /* (4, 9, 30) */,
  32'h3d11b684 /* (0, 9, 30) */,
  32'h3d2d8e0e /* (28, 5, 30) */,
  32'h3d149b5c /* (24, 5, 30) */,
  32'h3d346b02 /* (20, 5, 30) */,
  32'h3d28d1e5 /* (16, 5, 30) */,
  32'h3d346b02 /* (12, 5, 30) */,
  32'h3d149b5c /* (8, 5, 30) */,
  32'h3d2d8e0e /* (4, 5, 30) */,
  32'h3d5dd7d1 /* (0, 5, 30) */,
  32'h3d8b1391 /* (28, 1, 30) */,
  32'h3d15ce12 /* (24, 1, 30) */,
  32'h3d1cac31 /* (20, 1, 30) */,
  32'h3d09dfab /* (16, 1, 30) */,
  32'h3d1cac31 /* (12, 1, 30) */,
  32'h3d15ce12 /* (8, 1, 30) */,
  32'h3d8b1391 /* (4, 1, 30) */,
  32'h3e709592 /* (0, 1, 30) */,
  32'h3d1b3fff /* (28, 29, 26) */,
  32'h3d19bf4b /* (24, 29, 26) */,
  32'h3d48406d /* (20, 29, 26) */,
  32'h3d41d3ae /* (16, 29, 26) */,
  32'h3d48406d /* (12, 29, 26) */,
  32'h3d19bf4b /* (8, 29, 26) */,
  32'h3d1b3fff /* (4, 29, 26) */,
  32'h3d2d5b95 /* (0, 29, 26) */,
  32'h3d17902e /* (28, 25, 26) */,
  32'h3d35cd98 /* (24, 25, 26) */,
  32'h3d859348 /* (20, 25, 26) */,
  32'h3d8a46e7 /* (16, 25, 26) */,
  32'h3d859348 /* (12, 25, 26) */,
  32'h3d35cd98 /* (8, 25, 26) */,
  32'h3d17902e /* (4, 25, 26) */,
  32'h3d1459dd /* (0, 25, 26) */,
  32'h3d41fb9f /* (28, 21, 26) */,
  32'h3d865b59 /* (24, 21, 26) */,
  32'h3ddec971 /* (20, 21, 26) */,
  32'h3dfa4afe /* (16, 21, 26) */,
  32'h3ddec971 /* (12, 21, 26) */,
  32'h3d865b59 /* (8, 21, 26) */,
  32'h3d41fb9f /* (4, 21, 26) */,
  32'h3d3013e2 /* (0, 21, 26) */,
  32'h3d61b1de /* (28, 17, 26) */,
  32'h3daa3349 /* (24, 17, 26) */,
  32'h3e1a3a56 /* (20, 17, 26) */,
  32'h3e3a3d1a /* (16, 17, 26) */,
  32'h3e1a3a56 /* (12, 17, 26) */,
  32'h3daa3349 /* (8, 17, 26) */,
  32'h3d61b1de /* (4, 17, 26) */,
  32'h3d455011 /* (0, 17, 26) */,
  32'h3d601ae9 /* (28, 13, 26) */,
  32'h3da2e7a9 /* (24, 13, 26) */,
  32'h3e0dc95f /* (20, 13, 26) */,
  32'h3e2576a9 /* (16, 13, 26) */,
  32'h3e0dc95f /* (12, 13, 26) */,
  32'h3da2e7a9 /* (8, 13, 26) */,
  32'h3d601ae9 /* (4, 13, 26) */,
  32'h3d4703b2 /* (0, 13, 26) */,
  32'h3d2657dd /* (28, 9, 26) */,
  32'h3d584c0c /* (24, 9, 26) */,
  32'h3da96159 /* (20, 9, 26) */,
  32'h3db6b309 /* (16, 9, 26) */,
  32'h3da96159 /* (12, 9, 26) */,
  32'h3d584c0c /* (8, 9, 26) */,
  32'h3d2657dd /* (4, 9, 26) */,
  32'h3d1bc36a /* (0, 9, 26) */,
  32'h3d153e19 /* (28, 5, 26) */,
  32'h3d22af34 /* (24, 5, 26) */,
  32'h3d6007ad /* (20, 5, 26) */,
  32'h3d5f53fb /* (16, 5, 26) */,
  32'h3d6007ad /* (12, 5, 26) */,
  32'h3d22af34 /* (8, 5, 26) */,
  32'h3d153e19 /* (4, 5, 26) */,
  32'h3d1b2f33 /* (0, 5, 26) */,
  32'h3d222a9c /* (28, 1, 26) */,
  32'h3d169650 /* (24, 1, 26) */,
  32'h3d3dc5f0 /* (20, 1, 26) */,
  32'h3d34b66a /* (16, 1, 26) */,
  32'h3d3dc5f0 /* (12, 1, 26) */,
  32'h3d169650 /* (8, 1, 26) */,
  32'h3d222a9c /* (4, 1, 26) */,
  32'h3d3f59b8 /* (0, 1, 26) */,
  32'h3d1cff11 /* (28, 29, 22) */,
  32'h3d48bc7e /* (24, 29, 22) */,
  32'h3d9aff71 /* (20, 29, 22) */,
  32'h3da59d10 /* (16, 29, 22) */,
  32'h3d9aff71 /* (12, 29, 22) */,
  32'h3d48bc7e /* (8, 29, 22) */,
  32'h3d1cff11 /* (4, 29, 22) */,
  32'h3d144f19 /* (0, 29, 22) */,
  32'h3d404057 /* (28, 25, 22) */,
  32'h3d83c517 /* (24, 25, 22) */,
  32'h3dd85675 /* (20, 25, 22) */,
  32'h3df142da /* (16, 25, 22) */,
  32'h3dd85675 /* (12, 25, 22) */,
  32'h3d83c517 /* (8, 25, 22) */,
  32'h3d404057 /* (4, 25, 22) */,
  32'h3d2f5f5a /* (0, 25, 22) */,
  32'h3d92b699 /* (28, 21, 22) */,
  32'h3dd7e578 /* (24, 21, 22) */,
  32'h3e3e5baf /* (20, 21, 22) */,
  32'h3e60898b /* (16, 21, 22) */,
  32'h3e3e5baf /* (12, 21, 22) */,
  32'h3dd7e578 /* (8, 21, 22) */,
  32'h3d92b699 /* (4, 21, 22) */,
  32'h3d819abc /* (0, 21, 22) */,
  32'h3dbdf4f8 /* (28, 17, 22) */,
  32'h3e135573 /* (24, 17, 22) */,
  32'h3e89fde5 /* (20, 17, 22) */,
  32'h3eabb572 /* (16, 17, 22) */,
  32'h3e89fde5 /* (12, 17, 22) */,
  32'h3e135573 /* (8, 17, 22) */,
  32'h3dbdf4f8 /* (4, 17, 22) */,
  32'h3da42e1b /* (0, 17, 22) */,
  32'h3db40e50 /* (28, 13, 22) */,
  32'h3e085939 /* (24, 13, 22) */,
  32'h3e7848b5 /* (20, 13, 22) */,
  32'h3e968a40 /* (16, 13, 22) */,
  32'h3e7848b5 /* (12, 13, 22) */,
  32'h3e085939 /* (8, 13, 22) */,
  32'h3db40e50 /* (4, 13, 22) */,
  32'h3d9d248b /* (0, 13, 22) */,
  32'h3d68b7a2 /* (28, 9, 22) */,
  32'h3da590e9 /* (24, 9, 22) */,
  32'h3e0cf021 /* (20, 9, 22) */,
  32'h3e21930d /* (16, 9, 22) */,
  32'h3e0cf021 /* (12, 9, 22) */,
  32'h3da590e9 /* (8, 9, 22) */,
  32'h3d68b7a2 /* (4, 9, 22) */,
  32'h3d50a575 /* (0, 9, 22) */,
  32'h3d28e3b2 /* (28, 5, 22) */,
  32'h3d5ef675 /* (24, 5, 22) */,
  32'h3db0e528 /* (20, 5, 22) */,
  32'h3dc0863e /* (16, 5, 22) */,
  32'h3db0e528 /* (12, 5, 22) */,
  32'h3d5ef675 /* (8, 5, 22) */,
  32'h3d28e3b2 /* (4, 5, 22) */,
  32'h3d1cee15 /* (0, 5, 22) */,
  32'h3d1839e3 /* (28, 1, 22) */,
  32'h3d3f0366 /* (24, 1, 22) */,
  32'h3d91435f /* (20, 1, 22) */,
  32'h3d99ac24 /* (16, 1, 22) */,
  32'h3d91435f /* (12, 1, 22) */,
  32'h3d3f0366 /* (8, 1, 22) */,
  32'h3d1839e3 /* (4, 1, 22) */,
  32'h3d1142bb /* (0, 1, 22) */,
  32'h3d3b1e93 /* (28, 29, 18) */,
  32'h3d880501 /* (24, 29, 18) */,
  32'h3decc5e8 /* (20, 29, 18) */,
  32'h3e0a27e7 /* (16, 29, 18) */,
  32'h3decc5e8 /* (12, 29, 18) */,
  32'h3d880501 /* (8, 29, 18) */,
  32'h3d3b1e93 /* (4, 29, 18) */,
  32'h3d262b6e /* (0, 29, 18) */,
  32'h3d800deb /* (28, 25, 18) */,
  32'h3dbf672f /* (24, 25, 18) */,
  32'h3e2baf50 /* (20, 25, 18) */,
  32'h3e4d7ce8 /* (16, 25, 18) */,
  32'h3e2baf50 /* (12, 25, 18) */,
  32'h3dbf672f /* (8, 25, 18) */,
  32'h3d800deb /* (4, 25, 18) */,
  32'h3d60bf24 /* (0, 25, 18) */,
  32'h3ddc0819 /* (28, 21, 18) */,
  32'h3e2a27e4 /* (24, 21, 18) */,
  32'h3e9ecc49 /* (20, 21, 18) */,
  32'h3ec4f0a1 /* (16, 21, 18) */,
  32'h3e9ecc49 /* (12, 21, 18) */,
  32'h3e2a27e4 /* (8, 21, 18) */,
  32'h3ddc0819 /* (4, 21, 18) */,
  32'h3dbe661f /* (0, 21, 18) */,
  32'h3e1c2ca1 /* (28, 17, 18) */,
  32'h3e79034c /* (24, 17, 18) */,
  32'h3ef15f91 /* (20, 17, 18) */,
  32'h3f1b42bd /* (16, 17, 18) */,
  32'h3ef15f91 /* (12, 17, 18) */,
  32'h3e79034c /* (8, 17, 18) */,
  32'h3e1c2ca1 /* (4, 17, 18) */,
  32'h3e05899d /* (0, 17, 18) */,
  32'h3e0de89e /* (28, 13, 18) */,
  32'h3e5f05ce /* (24, 13, 18) */,
  32'h3ed441df /* (20, 13, 18) */,
  32'h3f06176f /* (16, 13, 18) */,
  32'h3ed441df /* (12, 13, 18) */,
  32'h3e5f05ce /* (8, 13, 18) */,
  32'h3e0de89e /* (4, 13, 18) */,
  32'h3df40add /* (0, 13, 18) */,
  32'h3da4db8a /* (28, 9, 18) */,
  32'h3dfaaa60 /* (24, 9, 18) */,
  32'h3e654448 /* (20, 9, 18) */,
  32'h3e8b9344 /* (16, 9, 18) */,
  32'h3e654448 /* (12, 9, 18) */,
  32'h3dfaaa60 /* (8, 9, 18) */,
  32'h3da4db8a /* (4, 9, 18) */,
  32'h3d8fa52c /* (0, 9, 18) */,
  32'h3d53bb31 /* (28, 5, 18) */,
  32'h3d9bc970 /* (24, 5, 18) */,
  32'h3e095be4 /* (20, 5, 18) */,
  32'h3e2205a1 /* (16, 5, 18) */,
  32'h3e095be4 /* (12, 5, 18) */,
  32'h3d9bc970 /* (8, 5, 18) */,
  32'h3d53bb31 /* (4, 5, 18) */,
  32'h3d3b0a55 /* (0, 5, 18) */,
  32'h3d303352 /* (28, 1, 18) */,
  32'h3d7e759f /* (24, 1, 18) */,
  32'h3ddbed5a /* (20, 1, 18) */,
  32'h3dff32bb /* (16, 1, 18) */,
  32'h3ddbed5a /* (12, 1, 18) */,
  32'h3d7e759f /* (8, 1, 18) */,
  32'h3d303352 /* (4, 1, 18) */,
  32'h3d1ceee6 /* (0, 1, 18) */,
  32'h3d3b1e93 /* (28, 29, 14) */,
  32'h3d880501 /* (24, 29, 14) */,
  32'h3decc5e8 /* (20, 29, 14) */,
  32'h3e0a27e7 /* (16, 29, 14) */,
  32'h3decc5e8 /* (12, 29, 14) */,
  32'h3d880501 /* (8, 29, 14) */,
  32'h3d3b1e93 /* (4, 29, 14) */,
  32'h3d262b6e /* (0, 29, 14) */,
  32'h3d800deb /* (28, 25, 14) */,
  32'h3dbf672f /* (24, 25, 14) */,
  32'h3e2baf50 /* (20, 25, 14) */,
  32'h3e4d7ce8 /* (16, 25, 14) */,
  32'h3e2baf50 /* (12, 25, 14) */,
  32'h3dbf672f /* (8, 25, 14) */,
  32'h3d800deb /* (4, 25, 14) */,
  32'h3d60bf24 /* (0, 25, 14) */,
  32'h3ddc0819 /* (28, 21, 14) */,
  32'h3e2a27e4 /* (24, 21, 14) */,
  32'h3e9ecc49 /* (20, 21, 14) */,
  32'h3ec4f0a1 /* (16, 21, 14) */,
  32'h3e9ecc49 /* (12, 21, 14) */,
  32'h3e2a27e4 /* (8, 21, 14) */,
  32'h3ddc0819 /* (4, 21, 14) */,
  32'h3dbe661f /* (0, 21, 14) */,
  32'h3e1c2ca1 /* (28, 17, 14) */,
  32'h3e79034c /* (24, 17, 14) */,
  32'h3ef15f91 /* (20, 17, 14) */,
  32'h3f1b42bd /* (16, 17, 14) */,
  32'h3ef15f91 /* (12, 17, 14) */,
  32'h3e79034c /* (8, 17, 14) */,
  32'h3e1c2ca1 /* (4, 17, 14) */,
  32'h3e05899d /* (0, 17, 14) */,
  32'h3e0de89e /* (28, 13, 14) */,
  32'h3e5f05ce /* (24, 13, 14) */,
  32'h3ed441df /* (20, 13, 14) */,
  32'h3f06176f /* (16, 13, 14) */,
  32'h3ed441df /* (12, 13, 14) */,
  32'h3e5f05ce /* (8, 13, 14) */,
  32'h3e0de89e /* (4, 13, 14) */,
  32'h3df40add /* (0, 13, 14) */,
  32'h3da4db8a /* (28, 9, 14) */,
  32'h3dfaaa60 /* (24, 9, 14) */,
  32'h3e654448 /* (20, 9, 14) */,
  32'h3e8b9344 /* (16, 9, 14) */,
  32'h3e654448 /* (12, 9, 14) */,
  32'h3dfaaa60 /* (8, 9, 14) */,
  32'h3da4db8a /* (4, 9, 14) */,
  32'h3d8fa52c /* (0, 9, 14) */,
  32'h3d53bb31 /* (28, 5, 14) */,
  32'h3d9bc970 /* (24, 5, 14) */,
  32'h3e095be4 /* (20, 5, 14) */,
  32'h3e2205a1 /* (16, 5, 14) */,
  32'h3e095be4 /* (12, 5, 14) */,
  32'h3d9bc970 /* (8, 5, 14) */,
  32'h3d53bb31 /* (4, 5, 14) */,
  32'h3d3b0a55 /* (0, 5, 14) */,
  32'h3d303352 /* (28, 1, 14) */,
  32'h3d7e759f /* (24, 1, 14) */,
  32'h3ddbed5a /* (20, 1, 14) */,
  32'h3dff32bb /* (16, 1, 14) */,
  32'h3ddbed5a /* (12, 1, 14) */,
  32'h3d7e759f /* (8, 1, 14) */,
  32'h3d303352 /* (4, 1, 14) */,
  32'h3d1ceee6 /* (0, 1, 14) */,
  32'h3d1cff11 /* (28, 29, 10) */,
  32'h3d48bc7e /* (24, 29, 10) */,
  32'h3d9aff71 /* (20, 29, 10) */,
  32'h3da59d10 /* (16, 29, 10) */,
  32'h3d9aff71 /* (12, 29, 10) */,
  32'h3d48bc7e /* (8, 29, 10) */,
  32'h3d1cff11 /* (4, 29, 10) */,
  32'h3d144f19 /* (0, 29, 10) */,
  32'h3d404057 /* (28, 25, 10) */,
  32'h3d83c517 /* (24, 25, 10) */,
  32'h3dd85675 /* (20, 25, 10) */,
  32'h3df142da /* (16, 25, 10) */,
  32'h3dd85675 /* (12, 25, 10) */,
  32'h3d83c517 /* (8, 25, 10) */,
  32'h3d404057 /* (4, 25, 10) */,
  32'h3d2f5f5a /* (0, 25, 10) */,
  32'h3d92b699 /* (28, 21, 10) */,
  32'h3dd7e578 /* (24, 21, 10) */,
  32'h3e3e5baf /* (20, 21, 10) */,
  32'h3e60898b /* (16, 21, 10) */,
  32'h3e3e5baf /* (12, 21, 10) */,
  32'h3dd7e578 /* (8, 21, 10) */,
  32'h3d92b699 /* (4, 21, 10) */,
  32'h3d819abc /* (0, 21, 10) */,
  32'h3dbdf4f8 /* (28, 17, 10) */,
  32'h3e135573 /* (24, 17, 10) */,
  32'h3e89fde5 /* (20, 17, 10) */,
  32'h3eabb572 /* (16, 17, 10) */,
  32'h3e89fde5 /* (12, 17, 10) */,
  32'h3e135573 /* (8, 17, 10) */,
  32'h3dbdf4f8 /* (4, 17, 10) */,
  32'h3da42e1b /* (0, 17, 10) */,
  32'h3db40e50 /* (28, 13, 10) */,
  32'h3e085939 /* (24, 13, 10) */,
  32'h3e7848b5 /* (20, 13, 10) */,
  32'h3e968a40 /* (16, 13, 10) */,
  32'h3e7848b5 /* (12, 13, 10) */,
  32'h3e085939 /* (8, 13, 10) */,
  32'h3db40e50 /* (4, 13, 10) */,
  32'h3d9d248b /* (0, 13, 10) */,
  32'h3d68b7a2 /* (28, 9, 10) */,
  32'h3da590e9 /* (24, 9, 10) */,
  32'h3e0cf021 /* (20, 9, 10) */,
  32'h3e21930d /* (16, 9, 10) */,
  32'h3e0cf021 /* (12, 9, 10) */,
  32'h3da590e9 /* (8, 9, 10) */,
  32'h3d68b7a2 /* (4, 9, 10) */,
  32'h3d50a575 /* (0, 9, 10) */,
  32'h3d28e3b2 /* (28, 5, 10) */,
  32'h3d5ef675 /* (24, 5, 10) */,
  32'h3db0e528 /* (20, 5, 10) */,
  32'h3dc0863e /* (16, 5, 10) */,
  32'h3db0e528 /* (12, 5, 10) */,
  32'h3d5ef675 /* (8, 5, 10) */,
  32'h3d28e3b2 /* (4, 5, 10) */,
  32'h3d1cee15 /* (0, 5, 10) */,
  32'h3d1839e3 /* (28, 1, 10) */,
  32'h3d3f0366 /* (24, 1, 10) */,
  32'h3d91435f /* (20, 1, 10) */,
  32'h3d99ac24 /* (16, 1, 10) */,
  32'h3d91435f /* (12, 1, 10) */,
  32'h3d3f0366 /* (8, 1, 10) */,
  32'h3d1839e3 /* (4, 1, 10) */,
  32'h3d1142bb /* (0, 1, 10) */,
  32'h3d1b3fff /* (28, 29, 6) */,
  32'h3d19bf4b /* (24, 29, 6) */,
  32'h3d48406d /* (20, 29, 6) */,
  32'h3d41d3ae /* (16, 29, 6) */,
  32'h3d48406d /* (12, 29, 6) */,
  32'h3d19bf4b /* (8, 29, 6) */,
  32'h3d1b3fff /* (4, 29, 6) */,
  32'h3d2d5b95 /* (0, 29, 6) */,
  32'h3d17902e /* (28, 25, 6) */,
  32'h3d35cd98 /* (24, 25, 6) */,
  32'h3d859348 /* (20, 25, 6) */,
  32'h3d8a46e7 /* (16, 25, 6) */,
  32'h3d859348 /* (12, 25, 6) */,
  32'h3d35cd98 /* (8, 25, 6) */,
  32'h3d17902e /* (4, 25, 6) */,
  32'h3d1459dd /* (0, 25, 6) */,
  32'h3d41fb9f /* (28, 21, 6) */,
  32'h3d865b59 /* (24, 21, 6) */,
  32'h3ddec971 /* (20, 21, 6) */,
  32'h3dfa4afe /* (16, 21, 6) */,
  32'h3ddec971 /* (12, 21, 6) */,
  32'h3d865b59 /* (8, 21, 6) */,
  32'h3d41fb9f /* (4, 21, 6) */,
  32'h3d3013e2 /* (0, 21, 6) */,
  32'h3d61b1de /* (28, 17, 6) */,
  32'h3daa3349 /* (24, 17, 6) */,
  32'h3e1a3a56 /* (20, 17, 6) */,
  32'h3e3a3d1a /* (16, 17, 6) */,
  32'h3e1a3a56 /* (12, 17, 6) */,
  32'h3daa3349 /* (8, 17, 6) */,
  32'h3d61b1de /* (4, 17, 6) */,
  32'h3d455011 /* (0, 17, 6) */,
  32'h3d601ae9 /* (28, 13, 6) */,
  32'h3da2e7a9 /* (24, 13, 6) */,
  32'h3e0dc95f /* (20, 13, 6) */,
  32'h3e2576a9 /* (16, 13, 6) */,
  32'h3e0dc95f /* (12, 13, 6) */,
  32'h3da2e7a9 /* (8, 13, 6) */,
  32'h3d601ae9 /* (4, 13, 6) */,
  32'h3d4703b2 /* (0, 13, 6) */,
  32'h3d2657dd /* (28, 9, 6) */,
  32'h3d584c0c /* (24, 9, 6) */,
  32'h3da96159 /* (20, 9, 6) */,
  32'h3db6b309 /* (16, 9, 6) */,
  32'h3da96159 /* (12, 9, 6) */,
  32'h3d584c0c /* (8, 9, 6) */,
  32'h3d2657dd /* (4, 9, 6) */,
  32'h3d1bc36a /* (0, 9, 6) */,
  32'h3d153e19 /* (28, 5, 6) */,
  32'h3d22af34 /* (24, 5, 6) */,
  32'h3d6007ad /* (20, 5, 6) */,
  32'h3d5f53fb /* (16, 5, 6) */,
  32'h3d6007ad /* (12, 5, 6) */,
  32'h3d22af34 /* (8, 5, 6) */,
  32'h3d153e19 /* (4, 5, 6) */,
  32'h3d1b2f33 /* (0, 5, 6) */,
  32'h3d222a9c /* (28, 1, 6) */,
  32'h3d169650 /* (24, 1, 6) */,
  32'h3d3dc5f0 /* (20, 1, 6) */,
  32'h3d34b66a /* (16, 1, 6) */,
  32'h3d3dc5f0 /* (12, 1, 6) */,
  32'h3d169650 /* (8, 1, 6) */,
  32'h3d222a9c /* (4, 1, 6) */,
  32'h3d3f59b8 /* (0, 1, 6) */,
  32'h3d5defd3 /* (28, 29, 2) */,
  32'h3d13e9f7 /* (24, 29, 2) */,
  32'h3d23d587 /* (20, 29, 2) */,
  32'h3d13661d /* (16, 29, 2) */,
  32'h3d23d587 /* (12, 29, 2) */,
  32'h3d13e9f7 /* (8, 29, 2) */,
  32'h3d5defd3 /* (4, 29, 2) */,
  32'h3dcbea25 /* (0, 29, 2) */,
  32'h3d16c6a3 /* (28, 25, 2) */,
  32'h3d1d59b0 /* (24, 25, 2) */,
  32'h3d530d8e /* (20, 25, 2) */,
  32'h3d4f6a6e /* (16, 25, 2) */,
  32'h3d530d8e /* (12, 25, 2) */,
  32'h3d1d59b0 /* (8, 25, 2) */,
  32'h3d16c6a3 /* (4, 25, 2) */,
  32'h3d21b235 /* (0, 25, 2) */,
  32'h3d21c128 /* (28, 21, 2) */,
  32'h3d558b1c /* (24, 21, 2) */,
  32'h3da96c08 /* (20, 21, 2) */,
  32'h3db86416 /* (16, 21, 2) */,
  32'h3da96c08 /* (12, 21, 2) */,
  32'h3d558b1c /* (8, 21, 2) */,
  32'h3d21c128 /* (4, 21, 2) */,
  32'h3d164ce1 /* (0, 21, 2) */,
  32'h3d2d6bba /* (28, 17, 2) */,
  32'h3d804df8 /* (24, 17, 2) */,
  32'h3de39dff /* (20, 17, 2) */,
  32'h3e06ec2e /* (16, 17, 2) */,
  32'h3de39dff /* (12, 17, 2) */,
  32'h3d804df8 /* (8, 17, 2) */,
  32'h3d2d6bba /* (4, 17, 2) */,
  32'h3d18d610 /* (0, 17, 2) */,
  32'h3d3217f4 /* (28, 13, 2) */,
  32'h3d7b52f8 /* (24, 13, 2) */,
  32'h3dd42d31 /* (20, 13, 2) */,
  32'h3df1ae3d /* (16, 13, 2) */,
  32'h3dd42d31 /* (12, 13, 2) */,
  32'h3d7b52f8 /* (8, 13, 2) */,
  32'h3d3217f4 /* (4, 13, 2) */,
  32'h3d2045b1 /* (0, 13, 2) */,
  32'h3d14de35 /* (28, 9, 2) */,
  32'h3d3291f6 /* (24, 9, 2) */,
  32'h3d833332 /* (20, 9, 2) */,
  32'h3d87d16b /* (16, 9, 2) */,
  32'h3d833332 /* (12, 9, 2) */,
  32'h3d3291f6 /* (8, 9, 2) */,
  32'h3d14de35 /* (4, 9, 2) */,
  32'h3d11b684 /* (0, 9, 2) */,
  32'h3d2d8e0e /* (28, 5, 2) */,
  32'h3d149b5c /* (24, 5, 2) */,
  32'h3d346b02 /* (20, 5, 2) */,
  32'h3d28d1e5 /* (16, 5, 2) */,
  32'h3d346b02 /* (12, 5, 2) */,
  32'h3d149b5c /* (8, 5, 2) */,
  32'h3d2d8e0e /* (4, 5, 2) */,
  32'h3d5dd7d1 /* (0, 5, 2) */,
  32'h3d8b1391 /* (28, 1, 2) */,
  32'h3d15ce12 /* (24, 1, 2) */,
  32'h3d1cac31 /* (20, 1, 2) */,
  32'h3d09dfab /* (16, 1, 2) */,
  32'h3d1cac31 /* (12, 1, 2) */,
  32'h3d15ce12 /* (8, 1, 2) */,
  32'h3d8b1391 /* (4, 1, 2) */,
  32'h3e709592 /* (0, 1, 2) */,
  32'h3d8b1391 /* (31, 28, 30) */,
  32'h3d2d8e0e /* (27, 28, 30) */,
  32'h3d14de35 /* (23, 28, 30) */,
  32'h3d3217f4 /* (19, 28, 30) */,
  32'h3d2d6bba /* (15, 28, 30) */,
  32'h3d21c128 /* (11, 28, 30) */,
  32'h3d16c6a3 /* (7, 28, 30) */,
  32'h3d5defd3 /* (3, 28, 30) */,
  32'h3d15ce12 /* (31, 24, 30) */,
  32'h3d149b5c /* (27, 24, 30) */,
  32'h3d3291f6 /* (23, 24, 30) */,
  32'h3d7b52f8 /* (19, 24, 30) */,
  32'h3d804df8 /* (15, 24, 30) */,
  32'h3d558b1c /* (11, 24, 30) */,
  32'h3d1d59b0 /* (7, 24, 30) */,
  32'h3d13e9f7 /* (3, 24, 30) */,
  32'h3d1cac31 /* (31, 20, 30) */,
  32'h3d346b02 /* (27, 20, 30) */,
  32'h3d833332 /* (23, 20, 30) */,
  32'h3dd42d31 /* (19, 20, 30) */,
  32'h3de39dff /* (15, 20, 30) */,
  32'h3da96c08 /* (11, 20, 30) */,
  32'h3d530d8e /* (7, 20, 30) */,
  32'h3d23d587 /* (3, 20, 30) */,
  32'h3d09dfab /* (31, 16, 30) */,
  32'h3d28d1e5 /* (27, 16, 30) */,
  32'h3d87d16b /* (23, 16, 30) */,
  32'h3df1ae3d /* (19, 16, 30) */,
  32'h3e06ec2e /* (15, 16, 30) */,
  32'h3db86416 /* (11, 16, 30) */,
  32'h3d4f6a6e /* (7, 16, 30) */,
  32'h3d13661d /* (3, 16, 30) */,
  32'h3d1cac31 /* (31, 12, 30) */,
  32'h3d346b02 /* (27, 12, 30) */,
  32'h3d833332 /* (23, 12, 30) */,
  32'h3dd42d31 /* (19, 12, 30) */,
  32'h3de39dff /* (15, 12, 30) */,
  32'h3da96c08 /* (11, 12, 30) */,
  32'h3d530d8e /* (7, 12, 30) */,
  32'h3d23d587 /* (3, 12, 30) */,
  32'h3d15ce12 /* (31, 8, 30) */,
  32'h3d149b5c /* (27, 8, 30) */,
  32'h3d3291f6 /* (23, 8, 30) */,
  32'h3d7b52f8 /* (19, 8, 30) */,
  32'h3d804df8 /* (15, 8, 30) */,
  32'h3d558b1c /* (11, 8, 30) */,
  32'h3d1d59b0 /* (7, 8, 30) */,
  32'h3d13e9f7 /* (3, 8, 30) */,
  32'h3d8b1391 /* (31, 4, 30) */,
  32'h3d2d8e0e /* (27, 4, 30) */,
  32'h3d14de35 /* (23, 4, 30) */,
  32'h3d3217f4 /* (19, 4, 30) */,
  32'h3d2d6bba /* (15, 4, 30) */,
  32'h3d21c128 /* (11, 4, 30) */,
  32'h3d16c6a3 /* (7, 4, 30) */,
  32'h3d5defd3 /* (3, 4, 30) */,
  32'h3e709592 /* (31, 0, 30) */,
  32'h3d5dd7d1 /* (27, 0, 30) */,
  32'h3d11b684 /* (23, 0, 30) */,
  32'h3d2045b1 /* (19, 0, 30) */,
  32'h3d18d610 /* (15, 0, 30) */,
  32'h3d164ce1 /* (11, 0, 30) */,
  32'h3d21b235 /* (7, 0, 30) */,
  32'h3dcbea25 /* (3, 0, 30) */,
  32'h3d222a9c /* (31, 28, 26) */,
  32'h3d153e19 /* (27, 28, 26) */,
  32'h3d2657dd /* (23, 28, 26) */,
  32'h3d601ae9 /* (19, 28, 26) */,
  32'h3d61b1de /* (15, 28, 26) */,
  32'h3d41fb9f /* (11, 28, 26) */,
  32'h3d17902e /* (7, 28, 26) */,
  32'h3d1b3fff /* (3, 28, 26) */,
  32'h3d169650 /* (31, 24, 26) */,
  32'h3d22af34 /* (27, 24, 26) */,
  32'h3d584c0c /* (23, 24, 26) */,
  32'h3da2e7a9 /* (19, 24, 26) */,
  32'h3daa3349 /* (15, 24, 26) */,
  32'h3d865b59 /* (11, 24, 26) */,
  32'h3d35cd98 /* (7, 24, 26) */,
  32'h3d19bf4b /* (3, 24, 26) */,
  32'h3d3dc5f0 /* (31, 20, 26) */,
  32'h3d6007ad /* (27, 20, 26) */,
  32'h3da96159 /* (23, 20, 26) */,
  32'h3e0dc95f /* (19, 20, 26) */,
  32'h3e1a3a56 /* (15, 20, 26) */,
  32'h3ddec971 /* (11, 20, 26) */,
  32'h3d859348 /* (7, 20, 26) */,
  32'h3d48406d /* (3, 20, 26) */,
  32'h3d34b66a /* (31, 16, 26) */,
  32'h3d5f53fb /* (27, 16, 26) */,
  32'h3db6b309 /* (23, 16, 26) */,
  32'h3e2576a9 /* (19, 16, 26) */,
  32'h3e3a3d1a /* (15, 16, 26) */,
  32'h3dfa4afe /* (11, 16, 26) */,
  32'h3d8a46e7 /* (7, 16, 26) */,
  32'h3d41d3ae /* (3, 16, 26) */,
  32'h3d3dc5f0 /* (31, 12, 26) */,
  32'h3d6007ad /* (27, 12, 26) */,
  32'h3da96159 /* (23, 12, 26) */,
  32'h3e0dc95f /* (19, 12, 26) */,
  32'h3e1a3a56 /* (15, 12, 26) */,
  32'h3ddec971 /* (11, 12, 26) */,
  32'h3d859348 /* (7, 12, 26) */,
  32'h3d48406d /* (3, 12, 26) */,
  32'h3d169650 /* (31, 8, 26) */,
  32'h3d22af34 /* (27, 8, 26) */,
  32'h3d584c0c /* (23, 8, 26) */,
  32'h3da2e7a9 /* (19, 8, 26) */,
  32'h3daa3349 /* (15, 8, 26) */,
  32'h3d865b59 /* (11, 8, 26) */,
  32'h3d35cd98 /* (7, 8, 26) */,
  32'h3d19bf4b /* (3, 8, 26) */,
  32'h3d222a9c /* (31, 4, 26) */,
  32'h3d153e19 /* (27, 4, 26) */,
  32'h3d2657dd /* (23, 4, 26) */,
  32'h3d601ae9 /* (19, 4, 26) */,
  32'h3d61b1de /* (15, 4, 26) */,
  32'h3d41fb9f /* (11, 4, 26) */,
  32'h3d17902e /* (7, 4, 26) */,
  32'h3d1b3fff /* (3, 4, 26) */,
  32'h3d3f59b8 /* (31, 0, 26) */,
  32'h3d1b2f33 /* (27, 0, 26) */,
  32'h3d1bc36a /* (23, 0, 26) */,
  32'h3d4703b2 /* (19, 0, 26) */,
  32'h3d455011 /* (15, 0, 26) */,
  32'h3d3013e2 /* (11, 0, 26) */,
  32'h3d1459dd /* (7, 0, 26) */,
  32'h3d2d5b95 /* (3, 0, 26) */,
  32'h3d1839e3 /* (31, 28, 22) */,
  32'h3d28e3b2 /* (27, 28, 22) */,
  32'h3d68b7a2 /* (23, 28, 22) */,
  32'h3db40e50 /* (19, 28, 22) */,
  32'h3dbdf4f8 /* (15, 28, 22) */,
  32'h3d92b699 /* (11, 28, 22) */,
  32'h3d404057 /* (7, 28, 22) */,
  32'h3d1cff11 /* (3, 28, 22) */,
  32'h3d3f0366 /* (31, 24, 22) */,
  32'h3d5ef675 /* (27, 24, 22) */,
  32'h3da590e9 /* (23, 24, 22) */,
  32'h3e085939 /* (19, 24, 22) */,
  32'h3e135573 /* (15, 24, 22) */,
  32'h3dd7e578 /* (11, 24, 22) */,
  32'h3d83c517 /* (7, 24, 22) */,
  32'h3d48bc7e /* (3, 24, 22) */,
  32'h3d91435f /* (31, 20, 22) */,
  32'h3db0e528 /* (27, 20, 22) */,
  32'h3e0cf021 /* (23, 20, 22) */,
  32'h3e7848b5 /* (19, 20, 22) */,
  32'h3e89fde5 /* (15, 20, 22) */,
  32'h3e3e5baf /* (11, 20, 22) */,
  32'h3dd85675 /* (7, 20, 22) */,
  32'h3d9aff71 /* (3, 20, 22) */,
  32'h3d99ac24 /* (31, 16, 22) */,
  32'h3dc0863e /* (27, 16, 22) */,
  32'h3e21930d /* (23, 16, 22) */,
  32'h3e968a40 /* (19, 16, 22) */,
  32'h3eabb572 /* (15, 16, 22) */,
  32'h3e60898b /* (11, 16, 22) */,
  32'h3df142da /* (7, 16, 22) */,
  32'h3da59d10 /* (3, 16, 22) */,
  32'h3d91435f /* (31, 12, 22) */,
  32'h3db0e528 /* (27, 12, 22) */,
  32'h3e0cf021 /* (23, 12, 22) */,
  32'h3e7848b5 /* (19, 12, 22) */,
  32'h3e89fde5 /* (15, 12, 22) */,
  32'h3e3e5baf /* (11, 12, 22) */,
  32'h3dd85675 /* (7, 12, 22) */,
  32'h3d9aff71 /* (3, 12, 22) */,
  32'h3d3f0366 /* (31, 8, 22) */,
  32'h3d5ef675 /* (27, 8, 22) */,
  32'h3da590e9 /* (23, 8, 22) */,
  32'h3e085939 /* (19, 8, 22) */,
  32'h3e135573 /* (15, 8, 22) */,
  32'h3dd7e578 /* (11, 8, 22) */,
  32'h3d83c517 /* (7, 8, 22) */,
  32'h3d48bc7e /* (3, 8, 22) */,
  32'h3d1839e3 /* (31, 4, 22) */,
  32'h3d28e3b2 /* (27, 4, 22) */,
  32'h3d68b7a2 /* (23, 4, 22) */,
  32'h3db40e50 /* (19, 4, 22) */,
  32'h3dbdf4f8 /* (15, 4, 22) */,
  32'h3d92b699 /* (11, 4, 22) */,
  32'h3d404057 /* (7, 4, 22) */,
  32'h3d1cff11 /* (3, 4, 22) */,
  32'h3d1142bb /* (31, 0, 22) */,
  32'h3d1cee15 /* (27, 0, 22) */,
  32'h3d50a575 /* (23, 0, 22) */,
  32'h3d9d248b /* (19, 0, 22) */,
  32'h3da42e1b /* (15, 0, 22) */,
  32'h3d819abc /* (11, 0, 22) */,
  32'h3d2f5f5a /* (7, 0, 22) */,
  32'h3d144f19 /* (3, 0, 22) */,
  32'h3d303352 /* (31, 28, 18) */,
  32'h3d53bb31 /* (27, 28, 18) */,
  32'h3da4db8a /* (23, 28, 18) */,
  32'h3e0de89e /* (19, 28, 18) */,
  32'h3e1c2ca1 /* (15, 28, 18) */,
  32'h3ddc0819 /* (11, 28, 18) */,
  32'h3d800deb /* (7, 28, 18) */,
  32'h3d3b1e93 /* (3, 28, 18) */,
  32'h3d7e759f /* (31, 24, 18) */,
  32'h3d9bc970 /* (27, 24, 18) */,
  32'h3dfaaa60 /* (23, 24, 18) */,
  32'h3e5f05ce /* (19, 24, 18) */,
  32'h3e79034c /* (15, 24, 18) */,
  32'h3e2a27e4 /* (11, 24, 18) */,
  32'h3dbf672f /* (7, 24, 18) */,
  32'h3d880501 /* (3, 24, 18) */,
  32'h3ddbed5a /* (31, 20, 18) */,
  32'h3e095be4 /* (27, 20, 18) */,
  32'h3e654448 /* (23, 20, 18) */,
  32'h3ed441df /* (19, 20, 18) */,
  32'h3ef15f91 /* (15, 20, 18) */,
  32'h3e9ecc49 /* (11, 20, 18) */,
  32'h3e2baf50 /* (7, 20, 18) */,
  32'h3decc5e8 /* (3, 20, 18) */,
  32'h3dff32bb /* (31, 16, 18) */,
  32'h3e2205a1 /* (27, 16, 18) */,
  32'h3e8b9344 /* (23, 16, 18) */,
  32'h3f06176f /* (19, 16, 18) */,
  32'h3f1b42bd /* (15, 16, 18) */,
  32'h3ec4f0a1 /* (11, 16, 18) */,
  32'h3e4d7ce8 /* (7, 16, 18) */,
  32'h3e0a27e7 /* (3, 16, 18) */,
  32'h3ddbed5a /* (31, 12, 18) */,
  32'h3e095be4 /* (27, 12, 18) */,
  32'h3e654448 /* (23, 12, 18) */,
  32'h3ed441df /* (19, 12, 18) */,
  32'h3ef15f91 /* (15, 12, 18) */,
  32'h3e9ecc49 /* (11, 12, 18) */,
  32'h3e2baf50 /* (7, 12, 18) */,
  32'h3decc5e8 /* (3, 12, 18) */,
  32'h3d7e759f /* (31, 8, 18) */,
  32'h3d9bc970 /* (27, 8, 18) */,
  32'h3dfaaa60 /* (23, 8, 18) */,
  32'h3e5f05ce /* (19, 8, 18) */,
  32'h3e79034c /* (15, 8, 18) */,
  32'h3e2a27e4 /* (11, 8, 18) */,
  32'h3dbf672f /* (7, 8, 18) */,
  32'h3d880501 /* (3, 8, 18) */,
  32'h3d303352 /* (31, 4, 18) */,
  32'h3d53bb31 /* (27, 4, 18) */,
  32'h3da4db8a /* (23, 4, 18) */,
  32'h3e0de89e /* (19, 4, 18) */,
  32'h3e1c2ca1 /* (15, 4, 18) */,
  32'h3ddc0819 /* (11, 4, 18) */,
  32'h3d800deb /* (7, 4, 18) */,
  32'h3d3b1e93 /* (3, 4, 18) */,
  32'h3d1ceee6 /* (31, 0, 18) */,
  32'h3d3b0a55 /* (27, 0, 18) */,
  32'h3d8fa52c /* (23, 0, 18) */,
  32'h3df40add /* (19, 0, 18) */,
  32'h3e05899d /* (15, 0, 18) */,
  32'h3dbe661f /* (11, 0, 18) */,
  32'h3d60bf24 /* (7, 0, 18) */,
  32'h3d262b6e /* (3, 0, 18) */,
  32'h3d303352 /* (31, 28, 14) */,
  32'h3d53bb31 /* (27, 28, 14) */,
  32'h3da4db8a /* (23, 28, 14) */,
  32'h3e0de89e /* (19, 28, 14) */,
  32'h3e1c2ca1 /* (15, 28, 14) */,
  32'h3ddc0819 /* (11, 28, 14) */,
  32'h3d800deb /* (7, 28, 14) */,
  32'h3d3b1e93 /* (3, 28, 14) */,
  32'h3d7e759f /* (31, 24, 14) */,
  32'h3d9bc970 /* (27, 24, 14) */,
  32'h3dfaaa60 /* (23, 24, 14) */,
  32'h3e5f05ce /* (19, 24, 14) */,
  32'h3e79034c /* (15, 24, 14) */,
  32'h3e2a27e4 /* (11, 24, 14) */,
  32'h3dbf672f /* (7, 24, 14) */,
  32'h3d880501 /* (3, 24, 14) */,
  32'h3ddbed5a /* (31, 20, 14) */,
  32'h3e095be4 /* (27, 20, 14) */,
  32'h3e654448 /* (23, 20, 14) */,
  32'h3ed441df /* (19, 20, 14) */,
  32'h3ef15f91 /* (15, 20, 14) */,
  32'h3e9ecc49 /* (11, 20, 14) */,
  32'h3e2baf50 /* (7, 20, 14) */,
  32'h3decc5e8 /* (3, 20, 14) */,
  32'h3dff32bb /* (31, 16, 14) */,
  32'h3e2205a1 /* (27, 16, 14) */,
  32'h3e8b9344 /* (23, 16, 14) */,
  32'h3f06176f /* (19, 16, 14) */,
  32'h3f1b42bd /* (15, 16, 14) */,
  32'h3ec4f0a1 /* (11, 16, 14) */,
  32'h3e4d7ce8 /* (7, 16, 14) */,
  32'h3e0a27e7 /* (3, 16, 14) */,
  32'h3ddbed5a /* (31, 12, 14) */,
  32'h3e095be4 /* (27, 12, 14) */,
  32'h3e654448 /* (23, 12, 14) */,
  32'h3ed441df /* (19, 12, 14) */,
  32'h3ef15f91 /* (15, 12, 14) */,
  32'h3e9ecc49 /* (11, 12, 14) */,
  32'h3e2baf50 /* (7, 12, 14) */,
  32'h3decc5e8 /* (3, 12, 14) */,
  32'h3d7e759f /* (31, 8, 14) */,
  32'h3d9bc970 /* (27, 8, 14) */,
  32'h3dfaaa60 /* (23, 8, 14) */,
  32'h3e5f05ce /* (19, 8, 14) */,
  32'h3e79034c /* (15, 8, 14) */,
  32'h3e2a27e4 /* (11, 8, 14) */,
  32'h3dbf672f /* (7, 8, 14) */,
  32'h3d880501 /* (3, 8, 14) */,
  32'h3d303352 /* (31, 4, 14) */,
  32'h3d53bb31 /* (27, 4, 14) */,
  32'h3da4db8a /* (23, 4, 14) */,
  32'h3e0de89e /* (19, 4, 14) */,
  32'h3e1c2ca1 /* (15, 4, 14) */,
  32'h3ddc0819 /* (11, 4, 14) */,
  32'h3d800deb /* (7, 4, 14) */,
  32'h3d3b1e93 /* (3, 4, 14) */,
  32'h3d1ceee6 /* (31, 0, 14) */,
  32'h3d3b0a55 /* (27, 0, 14) */,
  32'h3d8fa52c /* (23, 0, 14) */,
  32'h3df40add /* (19, 0, 14) */,
  32'h3e05899d /* (15, 0, 14) */,
  32'h3dbe661f /* (11, 0, 14) */,
  32'h3d60bf24 /* (7, 0, 14) */,
  32'h3d262b6e /* (3, 0, 14) */,
  32'h3d1839e3 /* (31, 28, 10) */,
  32'h3d28e3b2 /* (27, 28, 10) */,
  32'h3d68b7a2 /* (23, 28, 10) */,
  32'h3db40e50 /* (19, 28, 10) */,
  32'h3dbdf4f8 /* (15, 28, 10) */,
  32'h3d92b699 /* (11, 28, 10) */,
  32'h3d404057 /* (7, 28, 10) */,
  32'h3d1cff11 /* (3, 28, 10) */,
  32'h3d3f0366 /* (31, 24, 10) */,
  32'h3d5ef675 /* (27, 24, 10) */,
  32'h3da590e9 /* (23, 24, 10) */,
  32'h3e085939 /* (19, 24, 10) */,
  32'h3e135573 /* (15, 24, 10) */,
  32'h3dd7e578 /* (11, 24, 10) */,
  32'h3d83c517 /* (7, 24, 10) */,
  32'h3d48bc7e /* (3, 24, 10) */,
  32'h3d91435f /* (31, 20, 10) */,
  32'h3db0e528 /* (27, 20, 10) */,
  32'h3e0cf021 /* (23, 20, 10) */,
  32'h3e7848b5 /* (19, 20, 10) */,
  32'h3e89fde5 /* (15, 20, 10) */,
  32'h3e3e5baf /* (11, 20, 10) */,
  32'h3dd85675 /* (7, 20, 10) */,
  32'h3d9aff71 /* (3, 20, 10) */,
  32'h3d99ac24 /* (31, 16, 10) */,
  32'h3dc0863e /* (27, 16, 10) */,
  32'h3e21930d /* (23, 16, 10) */,
  32'h3e968a40 /* (19, 16, 10) */,
  32'h3eabb572 /* (15, 16, 10) */,
  32'h3e60898b /* (11, 16, 10) */,
  32'h3df142da /* (7, 16, 10) */,
  32'h3da59d10 /* (3, 16, 10) */,
  32'h3d91435f /* (31, 12, 10) */,
  32'h3db0e528 /* (27, 12, 10) */,
  32'h3e0cf021 /* (23, 12, 10) */,
  32'h3e7848b5 /* (19, 12, 10) */,
  32'h3e89fde5 /* (15, 12, 10) */,
  32'h3e3e5baf /* (11, 12, 10) */,
  32'h3dd85675 /* (7, 12, 10) */,
  32'h3d9aff71 /* (3, 12, 10) */,
  32'h3d3f0366 /* (31, 8, 10) */,
  32'h3d5ef675 /* (27, 8, 10) */,
  32'h3da590e9 /* (23, 8, 10) */,
  32'h3e085939 /* (19, 8, 10) */,
  32'h3e135573 /* (15, 8, 10) */,
  32'h3dd7e578 /* (11, 8, 10) */,
  32'h3d83c517 /* (7, 8, 10) */,
  32'h3d48bc7e /* (3, 8, 10) */,
  32'h3d1839e3 /* (31, 4, 10) */,
  32'h3d28e3b2 /* (27, 4, 10) */,
  32'h3d68b7a2 /* (23, 4, 10) */,
  32'h3db40e50 /* (19, 4, 10) */,
  32'h3dbdf4f8 /* (15, 4, 10) */,
  32'h3d92b699 /* (11, 4, 10) */,
  32'h3d404057 /* (7, 4, 10) */,
  32'h3d1cff11 /* (3, 4, 10) */,
  32'h3d1142bb /* (31, 0, 10) */,
  32'h3d1cee15 /* (27, 0, 10) */,
  32'h3d50a575 /* (23, 0, 10) */,
  32'h3d9d248b /* (19, 0, 10) */,
  32'h3da42e1b /* (15, 0, 10) */,
  32'h3d819abc /* (11, 0, 10) */,
  32'h3d2f5f5a /* (7, 0, 10) */,
  32'h3d144f19 /* (3, 0, 10) */,
  32'h3d222a9c /* (31, 28, 6) */,
  32'h3d153e19 /* (27, 28, 6) */,
  32'h3d2657dd /* (23, 28, 6) */,
  32'h3d601ae9 /* (19, 28, 6) */,
  32'h3d61b1de /* (15, 28, 6) */,
  32'h3d41fb9f /* (11, 28, 6) */,
  32'h3d17902e /* (7, 28, 6) */,
  32'h3d1b3fff /* (3, 28, 6) */,
  32'h3d169650 /* (31, 24, 6) */,
  32'h3d22af34 /* (27, 24, 6) */,
  32'h3d584c0c /* (23, 24, 6) */,
  32'h3da2e7a9 /* (19, 24, 6) */,
  32'h3daa3349 /* (15, 24, 6) */,
  32'h3d865b59 /* (11, 24, 6) */,
  32'h3d35cd98 /* (7, 24, 6) */,
  32'h3d19bf4b /* (3, 24, 6) */,
  32'h3d3dc5f0 /* (31, 20, 6) */,
  32'h3d6007ad /* (27, 20, 6) */,
  32'h3da96159 /* (23, 20, 6) */,
  32'h3e0dc95f /* (19, 20, 6) */,
  32'h3e1a3a56 /* (15, 20, 6) */,
  32'h3ddec971 /* (11, 20, 6) */,
  32'h3d859348 /* (7, 20, 6) */,
  32'h3d48406d /* (3, 20, 6) */,
  32'h3d34b66a /* (31, 16, 6) */,
  32'h3d5f53fb /* (27, 16, 6) */,
  32'h3db6b309 /* (23, 16, 6) */,
  32'h3e2576a9 /* (19, 16, 6) */,
  32'h3e3a3d1a /* (15, 16, 6) */,
  32'h3dfa4afe /* (11, 16, 6) */,
  32'h3d8a46e7 /* (7, 16, 6) */,
  32'h3d41d3ae /* (3, 16, 6) */,
  32'h3d3dc5f0 /* (31, 12, 6) */,
  32'h3d6007ad /* (27, 12, 6) */,
  32'h3da96159 /* (23, 12, 6) */,
  32'h3e0dc95f /* (19, 12, 6) */,
  32'h3e1a3a56 /* (15, 12, 6) */,
  32'h3ddec971 /* (11, 12, 6) */,
  32'h3d859348 /* (7, 12, 6) */,
  32'h3d48406d /* (3, 12, 6) */,
  32'h3d169650 /* (31, 8, 6) */,
  32'h3d22af34 /* (27, 8, 6) */,
  32'h3d584c0c /* (23, 8, 6) */,
  32'h3da2e7a9 /* (19, 8, 6) */,
  32'h3daa3349 /* (15, 8, 6) */,
  32'h3d865b59 /* (11, 8, 6) */,
  32'h3d35cd98 /* (7, 8, 6) */,
  32'h3d19bf4b /* (3, 8, 6) */,
  32'h3d222a9c /* (31, 4, 6) */,
  32'h3d153e19 /* (27, 4, 6) */,
  32'h3d2657dd /* (23, 4, 6) */,
  32'h3d601ae9 /* (19, 4, 6) */,
  32'h3d61b1de /* (15, 4, 6) */,
  32'h3d41fb9f /* (11, 4, 6) */,
  32'h3d17902e /* (7, 4, 6) */,
  32'h3d1b3fff /* (3, 4, 6) */,
  32'h3d3f59b8 /* (31, 0, 6) */,
  32'h3d1b2f33 /* (27, 0, 6) */,
  32'h3d1bc36a /* (23, 0, 6) */,
  32'h3d4703b2 /* (19, 0, 6) */,
  32'h3d455011 /* (15, 0, 6) */,
  32'h3d3013e2 /* (11, 0, 6) */,
  32'h3d1459dd /* (7, 0, 6) */,
  32'h3d2d5b95 /* (3, 0, 6) */,
  32'h3d8b1391 /* (31, 28, 2) */,
  32'h3d2d8e0e /* (27, 28, 2) */,
  32'h3d14de35 /* (23, 28, 2) */,
  32'h3d3217f4 /* (19, 28, 2) */,
  32'h3d2d6bba /* (15, 28, 2) */,
  32'h3d21c128 /* (11, 28, 2) */,
  32'h3d16c6a3 /* (7, 28, 2) */,
  32'h3d5defd3 /* (3, 28, 2) */,
  32'h3d15ce12 /* (31, 24, 2) */,
  32'h3d149b5c /* (27, 24, 2) */,
  32'h3d3291f6 /* (23, 24, 2) */,
  32'h3d7b52f8 /* (19, 24, 2) */,
  32'h3d804df8 /* (15, 24, 2) */,
  32'h3d558b1c /* (11, 24, 2) */,
  32'h3d1d59b0 /* (7, 24, 2) */,
  32'h3d13e9f7 /* (3, 24, 2) */,
  32'h3d1cac31 /* (31, 20, 2) */,
  32'h3d346b02 /* (27, 20, 2) */,
  32'h3d833332 /* (23, 20, 2) */,
  32'h3dd42d31 /* (19, 20, 2) */,
  32'h3de39dff /* (15, 20, 2) */,
  32'h3da96c08 /* (11, 20, 2) */,
  32'h3d530d8e /* (7, 20, 2) */,
  32'h3d23d587 /* (3, 20, 2) */,
  32'h3d09dfab /* (31, 16, 2) */,
  32'h3d28d1e5 /* (27, 16, 2) */,
  32'h3d87d16b /* (23, 16, 2) */,
  32'h3df1ae3d /* (19, 16, 2) */,
  32'h3e06ec2e /* (15, 16, 2) */,
  32'h3db86416 /* (11, 16, 2) */,
  32'h3d4f6a6e /* (7, 16, 2) */,
  32'h3d13661d /* (3, 16, 2) */,
  32'h3d1cac31 /* (31, 12, 2) */,
  32'h3d346b02 /* (27, 12, 2) */,
  32'h3d833332 /* (23, 12, 2) */,
  32'h3dd42d31 /* (19, 12, 2) */,
  32'h3de39dff /* (15, 12, 2) */,
  32'h3da96c08 /* (11, 12, 2) */,
  32'h3d530d8e /* (7, 12, 2) */,
  32'h3d23d587 /* (3, 12, 2) */,
  32'h3d15ce12 /* (31, 8, 2) */,
  32'h3d149b5c /* (27, 8, 2) */,
  32'h3d3291f6 /* (23, 8, 2) */,
  32'h3d7b52f8 /* (19, 8, 2) */,
  32'h3d804df8 /* (15, 8, 2) */,
  32'h3d558b1c /* (11, 8, 2) */,
  32'h3d1d59b0 /* (7, 8, 2) */,
  32'h3d13e9f7 /* (3, 8, 2) */,
  32'h3d8b1391 /* (31, 4, 2) */,
  32'h3d2d8e0e /* (27, 4, 2) */,
  32'h3d14de35 /* (23, 4, 2) */,
  32'h3d3217f4 /* (19, 4, 2) */,
  32'h3d2d6bba /* (15, 4, 2) */,
  32'h3d21c128 /* (11, 4, 2) */,
  32'h3d16c6a3 /* (7, 4, 2) */,
  32'h3d5defd3 /* (3, 4, 2) */,
  32'h3e709592 /* (31, 0, 2) */,
  32'h3d5dd7d1 /* (27, 0, 2) */,
  32'h3d11b684 /* (23, 0, 2) */,
  32'h3d2045b1 /* (19, 0, 2) */,
  32'h3d18d610 /* (15, 0, 2) */,
  32'h3d164ce1 /* (11, 0, 2) */,
  32'h3d21b235 /* (7, 0, 2) */,
  32'h3dcbea25 /* (3, 0, 2) */,
  32'h3d7c66bd /* (30, 28, 30) */,
  32'h3d1f2a5d /* (26, 28, 30) */,
  32'h3d19eb69 /* (22, 28, 30) */,
  32'h3d3430e1 /* (18, 28, 30) */,
  32'h3d3430e1 /* (14, 28, 30) */,
  32'h3d19eb69 /* (10, 28, 30) */,
  32'h3d1f2a5d /* (6, 28, 30) */,
  32'h3d7c66bd /* (2, 28, 30) */,
  32'h3d14e1d9 /* (30, 24, 30) */,
  32'h3d17a967 /* (26, 24, 30) */,
  32'h3d428d9a /* (22, 24, 30) */,
  32'h3d8271c0 /* (18, 24, 30) */,
  32'h3d8271c0 /* (14, 24, 30) */,
  32'h3d428d9a /* (10, 24, 30) */,
  32'h3d17a967 /* (6, 24, 30) */,
  32'h3d14e1d9 /* (2, 24, 30) */,
  32'h3d1f454c /* (30, 20, 30) */,
  32'h3d41987e /* (26, 20, 30) */,
  32'h3d94d2ae /* (22, 20, 30) */,
  32'h3de2162b /* (18, 20, 30) */,
  32'h3de2162b /* (14, 20, 30) */,
  32'h3d94d2ae /* (10, 20, 30) */,
  32'h3d41987e /* (6, 20, 30) */,
  32'h3d1f454c /* (2, 20, 30) */,
  32'h3d0d5b74 /* (30, 16, 30) */,
  32'h3d39823a /* (26, 16, 30) */,
  32'h3d9e09be /* (22, 16, 30) */,
  32'h3e0374c7 /* (18, 16, 30) */,
  32'h3e0374c7 /* (14, 16, 30) */,
  32'h3d9e09be /* (10, 16, 30) */,
  32'h3d39823a /* (6, 16, 30) */,
  32'h3d0d5b74 /* (2, 16, 30) */,
  32'h3d1f454c /* (30, 12, 30) */,
  32'h3d41987e /* (26, 12, 30) */,
  32'h3d94d2ae /* (22, 12, 30) */,
  32'h3de2162b /* (18, 12, 30) */,
  32'h3de2162b /* (14, 12, 30) */,
  32'h3d94d2ae /* (10, 12, 30) */,
  32'h3d41987e /* (6, 12, 30) */,
  32'h3d1f454c /* (2, 12, 30) */,
  32'h3d14e1d9 /* (30, 8, 30) */,
  32'h3d17a967 /* (26, 8, 30) */,
  32'h3d428d9a /* (22, 8, 30) */,
  32'h3d8271c0 /* (18, 8, 30) */,
  32'h3d8271c0 /* (14, 8, 30) */,
  32'h3d428d9a /* (10, 8, 30) */,
  32'h3d17a967 /* (6, 8, 30) */,
  32'h3d14e1d9 /* (2, 8, 30) */,
  32'h3d7c66bd /* (30, 4, 30) */,
  32'h3d1f2a5d /* (26, 4, 30) */,
  32'h3d19eb69 /* (22, 4, 30) */,
  32'h3d3430e1 /* (18, 4, 30) */,
  32'h3d3430e1 /* (14, 4, 30) */,
  32'h3d19eb69 /* (10, 4, 30) */,
  32'h3d1f2a5d /* (6, 4, 30) */,
  32'h3d7c66bd /* (2, 4, 30) */,
  32'h3e1befb2 /* (30, 0, 30) */,
  32'h3d378ea1 /* (26, 0, 30) */,
  32'h3d124c17 /* (22, 0, 30) */,
  32'h3d204e75 /* (18, 0, 30) */,
  32'h3d204e75 /* (14, 0, 30) */,
  32'h3d124c17 /* (10, 0, 30) */,
  32'h3d378ea1 /* (6, 0, 30) */,
  32'h3e1befb2 /* (2, 0, 30) */,
  32'h3d1f2a5d /* (30, 28, 26) */,
  32'h3d1508f6 /* (26, 28, 26) */,
  32'h3d32cc97 /* (22, 28, 26) */,
  32'h3d66ec8b /* (18, 28, 26) */,
  32'h3d66ec8b /* (14, 28, 26) */,
  32'h3d32cc97 /* (10, 28, 26) */,
  32'h3d1508f6 /* (6, 28, 26) */,
  32'h3d1f2a5d /* (2, 28, 26) */,
  32'h3d17a967 /* (30, 24, 26) */,
  32'h3d2aa638 /* (26, 24, 26) */,
  32'h3d7076ff /* (22, 24, 26) */,
  32'h3dab2ff1 /* (18, 24, 26) */,
  32'h3dab2ff1 /* (14, 24, 26) */,
  32'h3d7076ff /* (10, 24, 26) */,
  32'h3d2aa638 /* (6, 24, 26) */,
  32'h3d17a967 /* (2, 24, 26) */,
  32'h3d41987e /* (30, 20, 26) */,
  32'h3d72a853 /* (26, 20, 26) */,
  32'h3dc1f419 /* (22, 20, 26) */,
  32'h3e182d5a /* (18, 20, 26) */,
  32'h3e182d5a /* (14, 20, 26) */,
  32'h3dc1f419 /* (10, 20, 26) */,
  32'h3d72a853 /* (6, 20, 26) */,
  32'h3d41987e /* (2, 20, 26) */,
  32'h3d39823a /* (30, 16, 26) */,
  32'h3d765452 /* (26, 16, 26) */,
  32'h3dd58e62 /* (22, 16, 26) */,
  32'h3e34be0d /* (18, 16, 26) */,
  32'h3e34be0d /* (14, 16, 26) */,
  32'h3dd58e62 /* (10, 16, 26) */,
  32'h3d765452 /* (6, 16, 26) */,
  32'h3d39823a /* (2, 16, 26) */,
  32'h3d41987e /* (30, 12, 26) */,
  32'h3d72a853 /* (26, 12, 26) */,
  32'h3dc1f419 /* (22, 12, 26) */,
  32'h3e182d5a /* (18, 12, 26) */,
  32'h3e182d5a /* (14, 12, 26) */,
  32'h3dc1f419 /* (10, 12, 26) */,
  32'h3d72a853 /* (6, 12, 26) */,
  32'h3d41987e /* (2, 12, 26) */,
  32'h3d17a967 /* (30, 8, 26) */,
  32'h3d2aa638 /* (26, 8, 26) */,
  32'h3d7076ff /* (22, 8, 26) */,
  32'h3dab2ff1 /* (18, 8, 26) */,
  32'h3dab2ff1 /* (14, 8, 26) */,
  32'h3d7076ff /* (10, 8, 26) */,
  32'h3d2aa638 /* (6, 8, 26) */,
  32'h3d17a967 /* (2, 8, 26) */,
  32'h3d1f2a5d /* (30, 4, 26) */,
  32'h3d1508f6 /* (26, 4, 26) */,
  32'h3d32cc97 /* (22, 4, 26) */,
  32'h3d66ec8b /* (18, 4, 26) */,
  32'h3d66ec8b /* (14, 4, 26) */,
  32'h3d32cc97 /* (10, 4, 26) */,
  32'h3d1508f6 /* (6, 4, 26) */,
  32'h3d1f2a5d /* (2, 4, 26) */,
  32'h3d378ea1 /* (30, 0, 26) */,
  32'h3d160c85 /* (26, 0, 26) */,
  32'h3d249cf9 /* (22, 0, 26) */,
  32'h3d4b578e /* (18, 0, 26) */,
  32'h3d4b578e /* (14, 0, 26) */,
  32'h3d249cf9 /* (10, 0, 26) */,
  32'h3d160c85 /* (6, 0, 26) */,
  32'h3d378ea1 /* (2, 0, 26) */,
  32'h3d19eb69 /* (30, 28, 22) */,
  32'h3d32cc97 /* (26, 28, 22) */,
  32'h3d825da2 /* (22, 28, 22) */,
  32'h3dbe2f24 /* (18, 28, 22) */,
  32'h3dbe2f24 /* (14, 28, 22) */,
  32'h3d825da2 /* (10, 28, 22) */,
  32'h3d32cc97 /* (6, 28, 22) */,
  32'h3d19eb69 /* (2, 28, 22) */,
  32'h3d428d9a /* (30, 24, 22) */,
  32'h3d7076ff /* (26, 24, 22) */,
  32'h3dbcbfdf /* (22, 24, 22) */,
  32'h3e11d65f /* (18, 24, 22) */,
  32'h3e11d65f /* (14, 24, 22) */,
  32'h3dbcbfdf /* (10, 24, 22) */,
  32'h3d7076ff /* (6, 24, 22) */,
  32'h3d428d9a /* (2, 24, 22) */,
  32'h3d94d2ae /* (30, 20, 22) */,
  32'h3dc1f419 /* (26, 20, 22) */,
  32'h3e239217 /* (22, 20, 22) */,
  32'h3e86bd25 /* (18, 20, 22) */,
  32'h3e86bd25 /* (14, 20, 22) */,
  32'h3e239217 /* (10, 20, 22) */,
  32'h3dc1f419 /* (6, 20, 22) */,
  32'h3d94d2ae /* (2, 20, 22) */,
  32'h3d9e09be /* (30, 16, 22) */,
  32'h3dd58e62 /* (26, 16, 22) */,
  32'h3e3e36ae /* (22, 16, 22) */,
  32'h3ea58eba /* (18, 16, 22) */,
  32'h3ea58eba /* (14, 16, 22) */,
  32'h3e3e36ae /* (10, 16, 22) */,
  32'h3dd58e62 /* (6, 16, 22) */,
  32'h3d9e09be /* (2, 16, 22) */,
  32'h3d94d2ae /* (30, 12, 22) */,
  32'h3dc1f419 /* (26, 12, 22) */,
  32'h3e239217 /* (22, 12, 22) */,
  32'h3e86bd25 /* (18, 12, 22) */,
  32'h3e86bd25 /* (14, 12, 22) */,
  32'h3e239217 /* (10, 12, 22) */,
  32'h3dc1f419 /* (6, 12, 22) */,
  32'h3d94d2ae /* (2, 12, 22) */,
  32'h3d428d9a /* (30, 8, 22) */,
  32'h3d7076ff /* (26, 8, 22) */,
  32'h3dbcbfdf /* (22, 8, 22) */,
  32'h3e11d65f /* (18, 8, 22) */,
  32'h3e11d65f /* (14, 8, 22) */,
  32'h3dbcbfdf /* (10, 8, 22) */,
  32'h3d7076ff /* (6, 8, 22) */,
  32'h3d428d9a /* (2, 8, 22) */,
  32'h3d19eb69 /* (30, 4, 22) */,
  32'h3d32cc97 /* (26, 4, 22) */,
  32'h3d825da2 /* (22, 4, 22) */,
  32'h3dbe2f24 /* (18, 4, 22) */,
  32'h3dbe2f24 /* (14, 4, 22) */,
  32'h3d825da2 /* (10, 4, 22) */,
  32'h3d32cc97 /* (6, 4, 22) */,
  32'h3d19eb69 /* (2, 4, 22) */,
  32'h3d124c17 /* (30, 0, 22) */,
  32'h3d249cf9 /* (26, 0, 22) */,
  32'h3d67f590 /* (22, 0, 22) */,
  32'h3da521d3 /* (18, 0, 22) */,
  32'h3da521d3 /* (14, 0, 22) */,
  32'h3d67f590 /* (10, 0, 22) */,
  32'h3d249cf9 /* (6, 0, 22) */,
  32'h3d124c17 /* (2, 0, 22) */,
  32'h3d3430e1 /* (30, 28, 18) */,
  32'h3d66ec8b /* (26, 28, 18) */,
  32'h3dbe2f24 /* (22, 28, 18) */,
  32'h3e193b79 /* (18, 28, 18) */,
  32'h3e193b79 /* (14, 28, 18) */,
  32'h3dbe2f24 /* (10, 28, 18) */,
  32'h3d66ec8b /* (6, 28, 18) */,
  32'h3d3430e1 /* (2, 28, 18) */,
  32'h3d8271c0 /* (30, 24, 18) */,
  32'h3dab2ff1 /* (26, 24, 18) */,
  32'h3e11d65f /* (22, 24, 18) */,
  32'h3e729d82 /* (18, 24, 18) */,
  32'h3e729d82 /* (14, 24, 18) */,
  32'h3e11d65f /* (10, 24, 18) */,
  32'h3dab2ff1 /* (6, 24, 18) */,
  32'h3d8271c0 /* (2, 24, 18) */,
  32'h3de2162b /* (30, 20, 18) */,
  32'h3e182d5a /* (26, 20, 18) */,
  32'h3e86bd25 /* (22, 20, 18) */,
  32'h3ee912bc /* (18, 20, 18) */,
  32'h3ee912bc /* (14, 20, 18) */,
  32'h3e86bd25 /* (10, 20, 18) */,
  32'h3e182d5a /* (6, 20, 18) */,
  32'h3de2162b /* (2, 20, 18) */,
  32'h3e0374c7 /* (30, 16, 18) */,
  32'h3e34be0d /* (26, 16, 18) */,
  32'h3ea58eba /* (22, 16, 18) */,
  32'h3f14977b /* (18, 16, 18) */,
  32'h3f14977b /* (14, 16, 18) */,
  32'h3ea58eba /* (10, 16, 18) */,
  32'h3e34be0d /* (6, 16, 18) */,
  32'h3e0374c7 /* (2, 16, 18) */,
  32'h3de2162b /* (30, 12, 18) */,
  32'h3e182d5a /* (26, 12, 18) */,
  32'h3e86bd25 /* (22, 12, 18) */,
  32'h3ee912bc /* (18, 12, 18) */,
  32'h3ee912bc /* (14, 12, 18) */,
  32'h3e86bd25 /* (10, 12, 18) */,
  32'h3e182d5a /* (6, 12, 18) */,
  32'h3de2162b /* (2, 12, 18) */,
  32'h3d8271c0 /* (30, 8, 18) */,
  32'h3dab2ff1 /* (26, 8, 18) */,
  32'h3e11d65f /* (22, 8, 18) */,
  32'h3e729d82 /* (18, 8, 18) */,
  32'h3e729d82 /* (14, 8, 18) */,
  32'h3e11d65f /* (10, 8, 18) */,
  32'h3dab2ff1 /* (6, 8, 18) */,
  32'h3d8271c0 /* (2, 8, 18) */,
  32'h3d3430e1 /* (30, 4, 18) */,
  32'h3d66ec8b /* (26, 4, 18) */,
  32'h3dbe2f24 /* (22, 4, 18) */,
  32'h3e193b79 /* (18, 4, 18) */,
  32'h3e193b79 /* (14, 4, 18) */,
  32'h3dbe2f24 /* (10, 4, 18) */,
  32'h3d66ec8b /* (6, 4, 18) */,
  32'h3d3430e1 /* (2, 4, 18) */,
  32'h3d204e75 /* (30, 0, 18) */,
  32'h3d4b578e /* (26, 0, 18) */,
  32'h3da521d3 /* (22, 0, 18) */,
  32'h3e036079 /* (18, 0, 18) */,
  32'h3e036079 /* (14, 0, 18) */,
  32'h3da521d3 /* (10, 0, 18) */,
  32'h3d4b578e /* (6, 0, 18) */,
  32'h3d204e75 /* (2, 0, 18) */,
  32'h3d3430e1 /* (30, 28, 14) */,
  32'h3d66ec8b /* (26, 28, 14) */,
  32'h3dbe2f24 /* (22, 28, 14) */,
  32'h3e193b79 /* (18, 28, 14) */,
  32'h3e193b79 /* (14, 28, 14) */,
  32'h3dbe2f24 /* (10, 28, 14) */,
  32'h3d66ec8b /* (6, 28, 14) */,
  32'h3d3430e1 /* (2, 28, 14) */,
  32'h3d8271c0 /* (30, 24, 14) */,
  32'h3dab2ff1 /* (26, 24, 14) */,
  32'h3e11d65f /* (22, 24, 14) */,
  32'h3e729d82 /* (18, 24, 14) */,
  32'h3e729d82 /* (14, 24, 14) */,
  32'h3e11d65f /* (10, 24, 14) */,
  32'h3dab2ff1 /* (6, 24, 14) */,
  32'h3d8271c0 /* (2, 24, 14) */,
  32'h3de2162b /* (30, 20, 14) */,
  32'h3e182d5a /* (26, 20, 14) */,
  32'h3e86bd25 /* (22, 20, 14) */,
  32'h3ee912bc /* (18, 20, 14) */,
  32'h3ee912bc /* (14, 20, 14) */,
  32'h3e86bd25 /* (10, 20, 14) */,
  32'h3e182d5a /* (6, 20, 14) */,
  32'h3de2162b /* (2, 20, 14) */,
  32'h3e0374c7 /* (30, 16, 14) */,
  32'h3e34be0d /* (26, 16, 14) */,
  32'h3ea58eba /* (22, 16, 14) */,
  32'h3f14977b /* (18, 16, 14) */,
  32'h3f14977b /* (14, 16, 14) */,
  32'h3ea58eba /* (10, 16, 14) */,
  32'h3e34be0d /* (6, 16, 14) */,
  32'h3e0374c7 /* (2, 16, 14) */,
  32'h3de2162b /* (30, 12, 14) */,
  32'h3e182d5a /* (26, 12, 14) */,
  32'h3e86bd25 /* (22, 12, 14) */,
  32'h3ee912bc /* (18, 12, 14) */,
  32'h3ee912bc /* (14, 12, 14) */,
  32'h3e86bd25 /* (10, 12, 14) */,
  32'h3e182d5a /* (6, 12, 14) */,
  32'h3de2162b /* (2, 12, 14) */,
  32'h3d8271c0 /* (30, 8, 14) */,
  32'h3dab2ff1 /* (26, 8, 14) */,
  32'h3e11d65f /* (22, 8, 14) */,
  32'h3e729d82 /* (18, 8, 14) */,
  32'h3e729d82 /* (14, 8, 14) */,
  32'h3e11d65f /* (10, 8, 14) */,
  32'h3dab2ff1 /* (6, 8, 14) */,
  32'h3d8271c0 /* (2, 8, 14) */,
  32'h3d3430e1 /* (30, 4, 14) */,
  32'h3d66ec8b /* (26, 4, 14) */,
  32'h3dbe2f24 /* (22, 4, 14) */,
  32'h3e193b79 /* (18, 4, 14) */,
  32'h3e193b79 /* (14, 4, 14) */,
  32'h3dbe2f24 /* (10, 4, 14) */,
  32'h3d66ec8b /* (6, 4, 14) */,
  32'h3d3430e1 /* (2, 4, 14) */,
  32'h3d204e75 /* (30, 0, 14) */,
  32'h3d4b578e /* (26, 0, 14) */,
  32'h3da521d3 /* (22, 0, 14) */,
  32'h3e036079 /* (18, 0, 14) */,
  32'h3e036079 /* (14, 0, 14) */,
  32'h3da521d3 /* (10, 0, 14) */,
  32'h3d4b578e /* (6, 0, 14) */,
  32'h3d204e75 /* (2, 0, 14) */,
  32'h3d19eb69 /* (30, 28, 10) */,
  32'h3d32cc97 /* (26, 28, 10) */,
  32'h3d825da2 /* (22, 28, 10) */,
  32'h3dbe2f24 /* (18, 28, 10) */,
  32'h3dbe2f24 /* (14, 28, 10) */,
  32'h3d825da2 /* (10, 28, 10) */,
  32'h3d32cc97 /* (6, 28, 10) */,
  32'h3d19eb69 /* (2, 28, 10) */,
  32'h3d428d9a /* (30, 24, 10) */,
  32'h3d7076ff /* (26, 24, 10) */,
  32'h3dbcbfdf /* (22, 24, 10) */,
  32'h3e11d65f /* (18, 24, 10) */,
  32'h3e11d65f /* (14, 24, 10) */,
  32'h3dbcbfdf /* (10, 24, 10) */,
  32'h3d7076ff /* (6, 24, 10) */,
  32'h3d428d9a /* (2, 24, 10) */,
  32'h3d94d2ae /* (30, 20, 10) */,
  32'h3dc1f419 /* (26, 20, 10) */,
  32'h3e239217 /* (22, 20, 10) */,
  32'h3e86bd25 /* (18, 20, 10) */,
  32'h3e86bd25 /* (14, 20, 10) */,
  32'h3e239217 /* (10, 20, 10) */,
  32'h3dc1f419 /* (6, 20, 10) */,
  32'h3d94d2ae /* (2, 20, 10) */,
  32'h3d9e09be /* (30, 16, 10) */,
  32'h3dd58e62 /* (26, 16, 10) */,
  32'h3e3e36ae /* (22, 16, 10) */,
  32'h3ea58eba /* (18, 16, 10) */,
  32'h3ea58eba /* (14, 16, 10) */,
  32'h3e3e36ae /* (10, 16, 10) */,
  32'h3dd58e62 /* (6, 16, 10) */,
  32'h3d9e09be /* (2, 16, 10) */,
  32'h3d94d2ae /* (30, 12, 10) */,
  32'h3dc1f419 /* (26, 12, 10) */,
  32'h3e239217 /* (22, 12, 10) */,
  32'h3e86bd25 /* (18, 12, 10) */,
  32'h3e86bd25 /* (14, 12, 10) */,
  32'h3e239217 /* (10, 12, 10) */,
  32'h3dc1f419 /* (6, 12, 10) */,
  32'h3d94d2ae /* (2, 12, 10) */,
  32'h3d428d9a /* (30, 8, 10) */,
  32'h3d7076ff /* (26, 8, 10) */,
  32'h3dbcbfdf /* (22, 8, 10) */,
  32'h3e11d65f /* (18, 8, 10) */,
  32'h3e11d65f /* (14, 8, 10) */,
  32'h3dbcbfdf /* (10, 8, 10) */,
  32'h3d7076ff /* (6, 8, 10) */,
  32'h3d428d9a /* (2, 8, 10) */,
  32'h3d19eb69 /* (30, 4, 10) */,
  32'h3d32cc97 /* (26, 4, 10) */,
  32'h3d825da2 /* (22, 4, 10) */,
  32'h3dbe2f24 /* (18, 4, 10) */,
  32'h3dbe2f24 /* (14, 4, 10) */,
  32'h3d825da2 /* (10, 4, 10) */,
  32'h3d32cc97 /* (6, 4, 10) */,
  32'h3d19eb69 /* (2, 4, 10) */,
  32'h3d124c17 /* (30, 0, 10) */,
  32'h3d249cf9 /* (26, 0, 10) */,
  32'h3d67f590 /* (22, 0, 10) */,
  32'h3da521d3 /* (18, 0, 10) */,
  32'h3da521d3 /* (14, 0, 10) */,
  32'h3d67f590 /* (10, 0, 10) */,
  32'h3d249cf9 /* (6, 0, 10) */,
  32'h3d124c17 /* (2, 0, 10) */,
  32'h3d1f2a5d /* (30, 28, 6) */,
  32'h3d1508f6 /* (26, 28, 6) */,
  32'h3d32cc97 /* (22, 28, 6) */,
  32'h3d66ec8b /* (18, 28, 6) */,
  32'h3d66ec8b /* (14, 28, 6) */,
  32'h3d32cc97 /* (10, 28, 6) */,
  32'h3d1508f6 /* (6, 28, 6) */,
  32'h3d1f2a5d /* (2, 28, 6) */,
  32'h3d17a967 /* (30, 24, 6) */,
  32'h3d2aa638 /* (26, 24, 6) */,
  32'h3d7076ff /* (22, 24, 6) */,
  32'h3dab2ff1 /* (18, 24, 6) */,
  32'h3dab2ff1 /* (14, 24, 6) */,
  32'h3d7076ff /* (10, 24, 6) */,
  32'h3d2aa638 /* (6, 24, 6) */,
  32'h3d17a967 /* (2, 24, 6) */,
  32'h3d41987e /* (30, 20, 6) */,
  32'h3d72a853 /* (26, 20, 6) */,
  32'h3dc1f419 /* (22, 20, 6) */,
  32'h3e182d5a /* (18, 20, 6) */,
  32'h3e182d5a /* (14, 20, 6) */,
  32'h3dc1f419 /* (10, 20, 6) */,
  32'h3d72a853 /* (6, 20, 6) */,
  32'h3d41987e /* (2, 20, 6) */,
  32'h3d39823a /* (30, 16, 6) */,
  32'h3d765452 /* (26, 16, 6) */,
  32'h3dd58e62 /* (22, 16, 6) */,
  32'h3e34be0d /* (18, 16, 6) */,
  32'h3e34be0d /* (14, 16, 6) */,
  32'h3dd58e62 /* (10, 16, 6) */,
  32'h3d765452 /* (6, 16, 6) */,
  32'h3d39823a /* (2, 16, 6) */,
  32'h3d41987e /* (30, 12, 6) */,
  32'h3d72a853 /* (26, 12, 6) */,
  32'h3dc1f419 /* (22, 12, 6) */,
  32'h3e182d5a /* (18, 12, 6) */,
  32'h3e182d5a /* (14, 12, 6) */,
  32'h3dc1f419 /* (10, 12, 6) */,
  32'h3d72a853 /* (6, 12, 6) */,
  32'h3d41987e /* (2, 12, 6) */,
  32'h3d17a967 /* (30, 8, 6) */,
  32'h3d2aa638 /* (26, 8, 6) */,
  32'h3d7076ff /* (22, 8, 6) */,
  32'h3dab2ff1 /* (18, 8, 6) */,
  32'h3dab2ff1 /* (14, 8, 6) */,
  32'h3d7076ff /* (10, 8, 6) */,
  32'h3d2aa638 /* (6, 8, 6) */,
  32'h3d17a967 /* (2, 8, 6) */,
  32'h3d1f2a5d /* (30, 4, 6) */,
  32'h3d1508f6 /* (26, 4, 6) */,
  32'h3d32cc97 /* (22, 4, 6) */,
  32'h3d66ec8b /* (18, 4, 6) */,
  32'h3d66ec8b /* (14, 4, 6) */,
  32'h3d32cc97 /* (10, 4, 6) */,
  32'h3d1508f6 /* (6, 4, 6) */,
  32'h3d1f2a5d /* (2, 4, 6) */,
  32'h3d378ea1 /* (30, 0, 6) */,
  32'h3d160c85 /* (26, 0, 6) */,
  32'h3d249cf9 /* (22, 0, 6) */,
  32'h3d4b578e /* (18, 0, 6) */,
  32'h3d4b578e /* (14, 0, 6) */,
  32'h3d249cf9 /* (10, 0, 6) */,
  32'h3d160c85 /* (6, 0, 6) */,
  32'h3d378ea1 /* (2, 0, 6) */,
  32'h3d7c66bd /* (30, 28, 2) */,
  32'h3d1f2a5d /* (26, 28, 2) */,
  32'h3d19eb69 /* (22, 28, 2) */,
  32'h3d3430e1 /* (18, 28, 2) */,
  32'h3d3430e1 /* (14, 28, 2) */,
  32'h3d19eb69 /* (10, 28, 2) */,
  32'h3d1f2a5d /* (6, 28, 2) */,
  32'h3d7c66bd /* (2, 28, 2) */,
  32'h3d14e1d9 /* (30, 24, 2) */,
  32'h3d17a967 /* (26, 24, 2) */,
  32'h3d428d9a /* (22, 24, 2) */,
  32'h3d8271c0 /* (18, 24, 2) */,
  32'h3d8271c0 /* (14, 24, 2) */,
  32'h3d428d9a /* (10, 24, 2) */,
  32'h3d17a967 /* (6, 24, 2) */,
  32'h3d14e1d9 /* (2, 24, 2) */,
  32'h3d1f454c /* (30, 20, 2) */,
  32'h3d41987e /* (26, 20, 2) */,
  32'h3d94d2ae /* (22, 20, 2) */,
  32'h3de2162b /* (18, 20, 2) */,
  32'h3de2162b /* (14, 20, 2) */,
  32'h3d94d2ae /* (10, 20, 2) */,
  32'h3d41987e /* (6, 20, 2) */,
  32'h3d1f454c /* (2, 20, 2) */,
  32'h3d0d5b74 /* (30, 16, 2) */,
  32'h3d39823a /* (26, 16, 2) */,
  32'h3d9e09be /* (22, 16, 2) */,
  32'h3e0374c7 /* (18, 16, 2) */,
  32'h3e0374c7 /* (14, 16, 2) */,
  32'h3d9e09be /* (10, 16, 2) */,
  32'h3d39823a /* (6, 16, 2) */,
  32'h3d0d5b74 /* (2, 16, 2) */,
  32'h3d1f454c /* (30, 12, 2) */,
  32'h3d41987e /* (26, 12, 2) */,
  32'h3d94d2ae /* (22, 12, 2) */,
  32'h3de2162b /* (18, 12, 2) */,
  32'h3de2162b /* (14, 12, 2) */,
  32'h3d94d2ae /* (10, 12, 2) */,
  32'h3d41987e /* (6, 12, 2) */,
  32'h3d1f454c /* (2, 12, 2) */,
  32'h3d14e1d9 /* (30, 8, 2) */,
  32'h3d17a967 /* (26, 8, 2) */,
  32'h3d428d9a /* (22, 8, 2) */,
  32'h3d8271c0 /* (18, 8, 2) */,
  32'h3d8271c0 /* (14, 8, 2) */,
  32'h3d428d9a /* (10, 8, 2) */,
  32'h3d17a967 /* (6, 8, 2) */,
  32'h3d14e1d9 /* (2, 8, 2) */,
  32'h3d7c66bd /* (30, 4, 2) */,
  32'h3d1f2a5d /* (26, 4, 2) */,
  32'h3d19eb69 /* (22, 4, 2) */,
  32'h3d3430e1 /* (18, 4, 2) */,
  32'h3d3430e1 /* (14, 4, 2) */,
  32'h3d19eb69 /* (10, 4, 2) */,
  32'h3d1f2a5d /* (6, 4, 2) */,
  32'h3d7c66bd /* (2, 4, 2) */,
  32'h3e1befb2 /* (30, 0, 2) */,
  32'h3d378ea1 /* (26, 0, 2) */,
  32'h3d124c17 /* (22, 0, 2) */,
  32'h3d204e75 /* (18, 0, 2) */,
  32'h3d204e75 /* (14, 0, 2) */,
  32'h3d124c17 /* (10, 0, 2) */,
  32'h3d378ea1 /* (6, 0, 2) */,
  32'h3e1befb2 /* (2, 0, 2) */,
  32'h3d5defd3 /* (29, 28, 30) */,
  32'h3d16c6a3 /* (25, 28, 30) */,
  32'h3d21c128 /* (21, 28, 30) */,
  32'h3d2d6bba /* (17, 28, 30) */,
  32'h3d3217f4 /* (13, 28, 30) */,
  32'h3d14de35 /* (9, 28, 30) */,
  32'h3d2d8e0e /* (5, 28, 30) */,
  32'h3d8b1391 /* (1, 28, 30) */,
  32'h3d13e9f7 /* (29, 24, 30) */,
  32'h3d1d59b0 /* (25, 24, 30) */,
  32'h3d558b1c /* (21, 24, 30) */,
  32'h3d804df8 /* (17, 24, 30) */,
  32'h3d7b52f8 /* (13, 24, 30) */,
  32'h3d3291f6 /* (9, 24, 30) */,
  32'h3d149b5c /* (5, 24, 30) */,
  32'h3d15ce12 /* (1, 24, 30) */,
  32'h3d23d587 /* (29, 20, 30) */,
  32'h3d530d8e /* (25, 20, 30) */,
  32'h3da96c08 /* (21, 20, 30) */,
  32'h3de39dff /* (17, 20, 30) */,
  32'h3dd42d31 /* (13, 20, 30) */,
  32'h3d833332 /* (9, 20, 30) */,
  32'h3d346b02 /* (5, 20, 30) */,
  32'h3d1cac31 /* (1, 20, 30) */,
  32'h3d13661d /* (29, 16, 30) */,
  32'h3d4f6a6e /* (25, 16, 30) */,
  32'h3db86416 /* (21, 16, 30) */,
  32'h3e06ec2e /* (17, 16, 30) */,
  32'h3df1ae3d /* (13, 16, 30) */,
  32'h3d87d16b /* (9, 16, 30) */,
  32'h3d28d1e5 /* (5, 16, 30) */,
  32'h3d09dfab /* (1, 16, 30) */,
  32'h3d23d587 /* (29, 12, 30) */,
  32'h3d530d8e /* (25, 12, 30) */,
  32'h3da96c08 /* (21, 12, 30) */,
  32'h3de39dff /* (17, 12, 30) */,
  32'h3dd42d31 /* (13, 12, 30) */,
  32'h3d833332 /* (9, 12, 30) */,
  32'h3d346b02 /* (5, 12, 30) */,
  32'h3d1cac31 /* (1, 12, 30) */,
  32'h3d13e9f7 /* (29, 8, 30) */,
  32'h3d1d59b0 /* (25, 8, 30) */,
  32'h3d558b1c /* (21, 8, 30) */,
  32'h3d804df8 /* (17, 8, 30) */,
  32'h3d7b52f8 /* (13, 8, 30) */,
  32'h3d3291f6 /* (9, 8, 30) */,
  32'h3d149b5c /* (5, 8, 30) */,
  32'h3d15ce12 /* (1, 8, 30) */,
  32'h3d5defd3 /* (29, 4, 30) */,
  32'h3d16c6a3 /* (25, 4, 30) */,
  32'h3d21c128 /* (21, 4, 30) */,
  32'h3d2d6bba /* (17, 4, 30) */,
  32'h3d3217f4 /* (13, 4, 30) */,
  32'h3d14de35 /* (9, 4, 30) */,
  32'h3d2d8e0e /* (5, 4, 30) */,
  32'h3d8b1391 /* (1, 4, 30) */,
  32'h3dcbea25 /* (29, 0, 30) */,
  32'h3d21b235 /* (25, 0, 30) */,
  32'h3d164ce1 /* (21, 0, 30) */,
  32'h3d18d610 /* (17, 0, 30) */,
  32'h3d2045b1 /* (13, 0, 30) */,
  32'h3d11b684 /* (9, 0, 30) */,
  32'h3d5dd7d1 /* (5, 0, 30) */,
  32'h3e709592 /* (1, 0, 30) */,
  32'h3d1b3fff /* (29, 28, 26) */,
  32'h3d17902e /* (25, 28, 26) */,
  32'h3d41fb9f /* (21, 28, 26) */,
  32'h3d61b1de /* (17, 28, 26) */,
  32'h3d601ae9 /* (13, 28, 26) */,
  32'h3d2657dd /* (9, 28, 26) */,
  32'h3d153e19 /* (5, 28, 26) */,
  32'h3d222a9c /* (1, 28, 26) */,
  32'h3d19bf4b /* (29, 24, 26) */,
  32'h3d35cd98 /* (25, 24, 26) */,
  32'h3d865b59 /* (21, 24, 26) */,
  32'h3daa3349 /* (17, 24, 26) */,
  32'h3da2e7a9 /* (13, 24, 26) */,
  32'h3d584c0c /* (9, 24, 26) */,
  32'h3d22af34 /* (5, 24, 26) */,
  32'h3d169650 /* (1, 24, 26) */,
  32'h3d48406d /* (29, 20, 26) */,
  32'h3d859348 /* (25, 20, 26) */,
  32'h3ddec971 /* (21, 20, 26) */,
  32'h3e1a3a56 /* (17, 20, 26) */,
  32'h3e0dc95f /* (13, 20, 26) */,
  32'h3da96159 /* (9, 20, 26) */,
  32'h3d6007ad /* (5, 20, 26) */,
  32'h3d3dc5f0 /* (1, 20, 26) */,
  32'h3d41d3ae /* (29, 16, 26) */,
  32'h3d8a46e7 /* (25, 16, 26) */,
  32'h3dfa4afe /* (21, 16, 26) */,
  32'h3e3a3d1a /* (17, 16, 26) */,
  32'h3e2576a9 /* (13, 16, 26) */,
  32'h3db6b309 /* (9, 16, 26) */,
  32'h3d5f53fb /* (5, 16, 26) */,
  32'h3d34b66a /* (1, 16, 26) */,
  32'h3d48406d /* (29, 12, 26) */,
  32'h3d859348 /* (25, 12, 26) */,
  32'h3ddec971 /* (21, 12, 26) */,
  32'h3e1a3a56 /* (17, 12, 26) */,
  32'h3e0dc95f /* (13, 12, 26) */,
  32'h3da96159 /* (9, 12, 26) */,
  32'h3d6007ad /* (5, 12, 26) */,
  32'h3d3dc5f0 /* (1, 12, 26) */,
  32'h3d19bf4b /* (29, 8, 26) */,
  32'h3d35cd98 /* (25, 8, 26) */,
  32'h3d865b59 /* (21, 8, 26) */,
  32'h3daa3349 /* (17, 8, 26) */,
  32'h3da2e7a9 /* (13, 8, 26) */,
  32'h3d584c0c /* (9, 8, 26) */,
  32'h3d22af34 /* (5, 8, 26) */,
  32'h3d169650 /* (1, 8, 26) */,
  32'h3d1b3fff /* (29, 4, 26) */,
  32'h3d17902e /* (25, 4, 26) */,
  32'h3d41fb9f /* (21, 4, 26) */,
  32'h3d61b1de /* (17, 4, 26) */,
  32'h3d601ae9 /* (13, 4, 26) */,
  32'h3d2657dd /* (9, 4, 26) */,
  32'h3d153e19 /* (5, 4, 26) */,
  32'h3d222a9c /* (1, 4, 26) */,
  32'h3d2d5b95 /* (29, 0, 26) */,
  32'h3d1459dd /* (25, 0, 26) */,
  32'h3d3013e2 /* (21, 0, 26) */,
  32'h3d455011 /* (17, 0, 26) */,
  32'h3d4703b2 /* (13, 0, 26) */,
  32'h3d1bc36a /* (9, 0, 26) */,
  32'h3d1b2f33 /* (5, 0, 26) */,
  32'h3d3f59b8 /* (1, 0, 26) */,
  32'h3d1cff11 /* (29, 28, 22) */,
  32'h3d404057 /* (25, 28, 22) */,
  32'h3d92b699 /* (21, 28, 22) */,
  32'h3dbdf4f8 /* (17, 28, 22) */,
  32'h3db40e50 /* (13, 28, 22) */,
  32'h3d68b7a2 /* (9, 28, 22) */,
  32'h3d28e3b2 /* (5, 28, 22) */,
  32'h3d1839e3 /* (1, 28, 22) */,
  32'h3d48bc7e /* (29, 24, 22) */,
  32'h3d83c517 /* (25, 24, 22) */,
  32'h3dd7e578 /* (21, 24, 22) */,
  32'h3e135573 /* (17, 24, 22) */,
  32'h3e085939 /* (13, 24, 22) */,
  32'h3da590e9 /* (9, 24, 22) */,
  32'h3d5ef675 /* (5, 24, 22) */,
  32'h3d3f0366 /* (1, 24, 22) */,
  32'h3d9aff71 /* (29, 20, 22) */,
  32'h3dd85675 /* (25, 20, 22) */,
  32'h3e3e5baf /* (21, 20, 22) */,
  32'h3e89fde5 /* (17, 20, 22) */,
  32'h3e7848b5 /* (13, 20, 22) */,
  32'h3e0cf021 /* (9, 20, 22) */,
  32'h3db0e528 /* (5, 20, 22) */,
  32'h3d91435f /* (1, 20, 22) */,
  32'h3da59d10 /* (29, 16, 22) */,
  32'h3df142da /* (25, 16, 22) */,
  32'h3e60898b /* (21, 16, 22) */,
  32'h3eabb572 /* (17, 16, 22) */,
  32'h3e968a40 /* (13, 16, 22) */,
  32'h3e21930d /* (9, 16, 22) */,
  32'h3dc0863e /* (5, 16, 22) */,
  32'h3d99ac24 /* (1, 16, 22) */,
  32'h3d9aff71 /* (29, 12, 22) */,
  32'h3dd85675 /* (25, 12, 22) */,
  32'h3e3e5baf /* (21, 12, 22) */,
  32'h3e89fde5 /* (17, 12, 22) */,
  32'h3e7848b5 /* (13, 12, 22) */,
  32'h3e0cf021 /* (9, 12, 22) */,
  32'h3db0e528 /* (5, 12, 22) */,
  32'h3d91435f /* (1, 12, 22) */,
  32'h3d48bc7e /* (29, 8, 22) */,
  32'h3d83c517 /* (25, 8, 22) */,
  32'h3dd7e578 /* (21, 8, 22) */,
  32'h3e135573 /* (17, 8, 22) */,
  32'h3e085939 /* (13, 8, 22) */,
  32'h3da590e9 /* (9, 8, 22) */,
  32'h3d5ef675 /* (5, 8, 22) */,
  32'h3d3f0366 /* (1, 8, 22) */,
  32'h3d1cff11 /* (29, 4, 22) */,
  32'h3d404057 /* (25, 4, 22) */,
  32'h3d92b699 /* (21, 4, 22) */,
  32'h3dbdf4f8 /* (17, 4, 22) */,
  32'h3db40e50 /* (13, 4, 22) */,
  32'h3d68b7a2 /* (9, 4, 22) */,
  32'h3d28e3b2 /* (5, 4, 22) */,
  32'h3d1839e3 /* (1, 4, 22) */,
  32'h3d144f19 /* (29, 0, 22) */,
  32'h3d2f5f5a /* (25, 0, 22) */,
  32'h3d819abc /* (21, 0, 22) */,
  32'h3da42e1b /* (17, 0, 22) */,
  32'h3d9d248b /* (13, 0, 22) */,
  32'h3d50a575 /* (9, 0, 22) */,
  32'h3d1cee15 /* (5, 0, 22) */,
  32'h3d1142bb /* (1, 0, 22) */,
  32'h3d3b1e93 /* (29, 28, 18) */,
  32'h3d800deb /* (25, 28, 18) */,
  32'h3ddc0819 /* (21, 28, 18) */,
  32'h3e1c2ca1 /* (17, 28, 18) */,
  32'h3e0de89e /* (13, 28, 18) */,
  32'h3da4db8a /* (9, 28, 18) */,
  32'h3d53bb31 /* (5, 28, 18) */,
  32'h3d303352 /* (1, 28, 18) */,
  32'h3d880501 /* (29, 24, 18) */,
  32'h3dbf672f /* (25, 24, 18) */,
  32'h3e2a27e4 /* (21, 24, 18) */,
  32'h3e79034c /* (17, 24, 18) */,
  32'h3e5f05ce /* (13, 24, 18) */,
  32'h3dfaaa60 /* (9, 24, 18) */,
  32'h3d9bc970 /* (5, 24, 18) */,
  32'h3d7e759f /* (1, 24, 18) */,
  32'h3decc5e8 /* (29, 20, 18) */,
  32'h3e2baf50 /* (25, 20, 18) */,
  32'h3e9ecc49 /* (21, 20, 18) */,
  32'h3ef15f91 /* (17, 20, 18) */,
  32'h3ed441df /* (13, 20, 18) */,
  32'h3e654448 /* (9, 20, 18) */,
  32'h3e095be4 /* (5, 20, 18) */,
  32'h3ddbed5a /* (1, 20, 18) */,
  32'h3e0a27e7 /* (29, 16, 18) */,
  32'h3e4d7ce8 /* (25, 16, 18) */,
  32'h3ec4f0a1 /* (21, 16, 18) */,
  32'h3f1b42bd /* (17, 16, 18) */,
  32'h3f06176f /* (13, 16, 18) */,
  32'h3e8b9344 /* (9, 16, 18) */,
  32'h3e2205a1 /* (5, 16, 18) */,
  32'h3dff32bb /* (1, 16, 18) */,
  32'h3decc5e8 /* (29, 12, 18) */,
  32'h3e2baf50 /* (25, 12, 18) */,
  32'h3e9ecc49 /* (21, 12, 18) */,
  32'h3ef15f91 /* (17, 12, 18) */,
  32'h3ed441df /* (13, 12, 18) */,
  32'h3e654448 /* (9, 12, 18) */,
  32'h3e095be4 /* (5, 12, 18) */,
  32'h3ddbed5a /* (1, 12, 18) */,
  32'h3d880501 /* (29, 8, 18) */,
  32'h3dbf672f /* (25, 8, 18) */,
  32'h3e2a27e4 /* (21, 8, 18) */,
  32'h3e79034c /* (17, 8, 18) */,
  32'h3e5f05ce /* (13, 8, 18) */,
  32'h3dfaaa60 /* (9, 8, 18) */,
  32'h3d9bc970 /* (5, 8, 18) */,
  32'h3d7e759f /* (1, 8, 18) */,
  32'h3d3b1e93 /* (29, 4, 18) */,
  32'h3d800deb /* (25, 4, 18) */,
  32'h3ddc0819 /* (21, 4, 18) */,
  32'h3e1c2ca1 /* (17, 4, 18) */,
  32'h3e0de89e /* (13, 4, 18) */,
  32'h3da4db8a /* (9, 4, 18) */,
  32'h3d53bb31 /* (5, 4, 18) */,
  32'h3d303352 /* (1, 4, 18) */,
  32'h3d262b6e /* (29, 0, 18) */,
  32'h3d60bf24 /* (25, 0, 18) */,
  32'h3dbe661f /* (21, 0, 18) */,
  32'h3e05899d /* (17, 0, 18) */,
  32'h3df40add /* (13, 0, 18) */,
  32'h3d8fa52c /* (9, 0, 18) */,
  32'h3d3b0a55 /* (5, 0, 18) */,
  32'h3d1ceee6 /* (1, 0, 18) */,
  32'h3d3b1e93 /* (29, 28, 14) */,
  32'h3d800deb /* (25, 28, 14) */,
  32'h3ddc0819 /* (21, 28, 14) */,
  32'h3e1c2ca1 /* (17, 28, 14) */,
  32'h3e0de89e /* (13, 28, 14) */,
  32'h3da4db8a /* (9, 28, 14) */,
  32'h3d53bb31 /* (5, 28, 14) */,
  32'h3d303352 /* (1, 28, 14) */,
  32'h3d880501 /* (29, 24, 14) */,
  32'h3dbf672f /* (25, 24, 14) */,
  32'h3e2a27e4 /* (21, 24, 14) */,
  32'h3e79034c /* (17, 24, 14) */,
  32'h3e5f05ce /* (13, 24, 14) */,
  32'h3dfaaa60 /* (9, 24, 14) */,
  32'h3d9bc970 /* (5, 24, 14) */,
  32'h3d7e759f /* (1, 24, 14) */,
  32'h3decc5e8 /* (29, 20, 14) */,
  32'h3e2baf50 /* (25, 20, 14) */,
  32'h3e9ecc49 /* (21, 20, 14) */,
  32'h3ef15f91 /* (17, 20, 14) */,
  32'h3ed441df /* (13, 20, 14) */,
  32'h3e654448 /* (9, 20, 14) */,
  32'h3e095be4 /* (5, 20, 14) */,
  32'h3ddbed5a /* (1, 20, 14) */,
  32'h3e0a27e7 /* (29, 16, 14) */,
  32'h3e4d7ce8 /* (25, 16, 14) */,
  32'h3ec4f0a1 /* (21, 16, 14) */,
  32'h3f1b42bd /* (17, 16, 14) */,
  32'h3f06176f /* (13, 16, 14) */,
  32'h3e8b9344 /* (9, 16, 14) */,
  32'h3e2205a1 /* (5, 16, 14) */,
  32'h3dff32bb /* (1, 16, 14) */,
  32'h3decc5e8 /* (29, 12, 14) */,
  32'h3e2baf50 /* (25, 12, 14) */,
  32'h3e9ecc49 /* (21, 12, 14) */,
  32'h3ef15f91 /* (17, 12, 14) */,
  32'h3ed441df /* (13, 12, 14) */,
  32'h3e654448 /* (9, 12, 14) */,
  32'h3e095be4 /* (5, 12, 14) */,
  32'h3ddbed5a /* (1, 12, 14) */,
  32'h3d880501 /* (29, 8, 14) */,
  32'h3dbf672f /* (25, 8, 14) */,
  32'h3e2a27e4 /* (21, 8, 14) */,
  32'h3e79034c /* (17, 8, 14) */,
  32'h3e5f05ce /* (13, 8, 14) */,
  32'h3dfaaa60 /* (9, 8, 14) */,
  32'h3d9bc970 /* (5, 8, 14) */,
  32'h3d7e759f /* (1, 8, 14) */,
  32'h3d3b1e93 /* (29, 4, 14) */,
  32'h3d800deb /* (25, 4, 14) */,
  32'h3ddc0819 /* (21, 4, 14) */,
  32'h3e1c2ca1 /* (17, 4, 14) */,
  32'h3e0de89e /* (13, 4, 14) */,
  32'h3da4db8a /* (9, 4, 14) */,
  32'h3d53bb31 /* (5, 4, 14) */,
  32'h3d303352 /* (1, 4, 14) */,
  32'h3d262b6e /* (29, 0, 14) */,
  32'h3d60bf24 /* (25, 0, 14) */,
  32'h3dbe661f /* (21, 0, 14) */,
  32'h3e05899d /* (17, 0, 14) */,
  32'h3df40add /* (13, 0, 14) */,
  32'h3d8fa52c /* (9, 0, 14) */,
  32'h3d3b0a55 /* (5, 0, 14) */,
  32'h3d1ceee6 /* (1, 0, 14) */,
  32'h3d1cff11 /* (29, 28, 10) */,
  32'h3d404057 /* (25, 28, 10) */,
  32'h3d92b699 /* (21, 28, 10) */,
  32'h3dbdf4f8 /* (17, 28, 10) */,
  32'h3db40e50 /* (13, 28, 10) */,
  32'h3d68b7a2 /* (9, 28, 10) */,
  32'h3d28e3b2 /* (5, 28, 10) */,
  32'h3d1839e3 /* (1, 28, 10) */,
  32'h3d48bc7e /* (29, 24, 10) */,
  32'h3d83c517 /* (25, 24, 10) */,
  32'h3dd7e578 /* (21, 24, 10) */,
  32'h3e135573 /* (17, 24, 10) */,
  32'h3e085939 /* (13, 24, 10) */,
  32'h3da590e9 /* (9, 24, 10) */,
  32'h3d5ef675 /* (5, 24, 10) */,
  32'h3d3f0366 /* (1, 24, 10) */,
  32'h3d9aff71 /* (29, 20, 10) */,
  32'h3dd85675 /* (25, 20, 10) */,
  32'h3e3e5baf /* (21, 20, 10) */,
  32'h3e89fde5 /* (17, 20, 10) */,
  32'h3e7848b5 /* (13, 20, 10) */,
  32'h3e0cf021 /* (9, 20, 10) */,
  32'h3db0e528 /* (5, 20, 10) */,
  32'h3d91435f /* (1, 20, 10) */,
  32'h3da59d10 /* (29, 16, 10) */,
  32'h3df142da /* (25, 16, 10) */,
  32'h3e60898b /* (21, 16, 10) */,
  32'h3eabb572 /* (17, 16, 10) */,
  32'h3e968a40 /* (13, 16, 10) */,
  32'h3e21930d /* (9, 16, 10) */,
  32'h3dc0863e /* (5, 16, 10) */,
  32'h3d99ac24 /* (1, 16, 10) */,
  32'h3d9aff71 /* (29, 12, 10) */,
  32'h3dd85675 /* (25, 12, 10) */,
  32'h3e3e5baf /* (21, 12, 10) */,
  32'h3e89fde5 /* (17, 12, 10) */,
  32'h3e7848b5 /* (13, 12, 10) */,
  32'h3e0cf021 /* (9, 12, 10) */,
  32'h3db0e528 /* (5, 12, 10) */,
  32'h3d91435f /* (1, 12, 10) */,
  32'h3d48bc7e /* (29, 8, 10) */,
  32'h3d83c517 /* (25, 8, 10) */,
  32'h3dd7e578 /* (21, 8, 10) */,
  32'h3e135573 /* (17, 8, 10) */,
  32'h3e085939 /* (13, 8, 10) */,
  32'h3da590e9 /* (9, 8, 10) */,
  32'h3d5ef675 /* (5, 8, 10) */,
  32'h3d3f0366 /* (1, 8, 10) */,
  32'h3d1cff11 /* (29, 4, 10) */,
  32'h3d404057 /* (25, 4, 10) */,
  32'h3d92b699 /* (21, 4, 10) */,
  32'h3dbdf4f8 /* (17, 4, 10) */,
  32'h3db40e50 /* (13, 4, 10) */,
  32'h3d68b7a2 /* (9, 4, 10) */,
  32'h3d28e3b2 /* (5, 4, 10) */,
  32'h3d1839e3 /* (1, 4, 10) */,
  32'h3d144f19 /* (29, 0, 10) */,
  32'h3d2f5f5a /* (25, 0, 10) */,
  32'h3d819abc /* (21, 0, 10) */,
  32'h3da42e1b /* (17, 0, 10) */,
  32'h3d9d248b /* (13, 0, 10) */,
  32'h3d50a575 /* (9, 0, 10) */,
  32'h3d1cee15 /* (5, 0, 10) */,
  32'h3d1142bb /* (1, 0, 10) */,
  32'h3d1b3fff /* (29, 28, 6) */,
  32'h3d17902e /* (25, 28, 6) */,
  32'h3d41fb9f /* (21, 28, 6) */,
  32'h3d61b1de /* (17, 28, 6) */,
  32'h3d601ae9 /* (13, 28, 6) */,
  32'h3d2657dd /* (9, 28, 6) */,
  32'h3d153e19 /* (5, 28, 6) */,
  32'h3d222a9c /* (1, 28, 6) */,
  32'h3d19bf4b /* (29, 24, 6) */,
  32'h3d35cd98 /* (25, 24, 6) */,
  32'h3d865b59 /* (21, 24, 6) */,
  32'h3daa3349 /* (17, 24, 6) */,
  32'h3da2e7a9 /* (13, 24, 6) */,
  32'h3d584c0c /* (9, 24, 6) */,
  32'h3d22af34 /* (5, 24, 6) */,
  32'h3d169650 /* (1, 24, 6) */,
  32'h3d48406d /* (29, 20, 6) */,
  32'h3d859348 /* (25, 20, 6) */,
  32'h3ddec971 /* (21, 20, 6) */,
  32'h3e1a3a56 /* (17, 20, 6) */,
  32'h3e0dc95f /* (13, 20, 6) */,
  32'h3da96159 /* (9, 20, 6) */,
  32'h3d6007ad /* (5, 20, 6) */,
  32'h3d3dc5f0 /* (1, 20, 6) */,
  32'h3d41d3ae /* (29, 16, 6) */,
  32'h3d8a46e7 /* (25, 16, 6) */,
  32'h3dfa4afe /* (21, 16, 6) */,
  32'h3e3a3d1a /* (17, 16, 6) */,
  32'h3e2576a9 /* (13, 16, 6) */,
  32'h3db6b309 /* (9, 16, 6) */,
  32'h3d5f53fb /* (5, 16, 6) */,
  32'h3d34b66a /* (1, 16, 6) */,
  32'h3d48406d /* (29, 12, 6) */,
  32'h3d859348 /* (25, 12, 6) */,
  32'h3ddec971 /* (21, 12, 6) */,
  32'h3e1a3a56 /* (17, 12, 6) */,
  32'h3e0dc95f /* (13, 12, 6) */,
  32'h3da96159 /* (9, 12, 6) */,
  32'h3d6007ad /* (5, 12, 6) */,
  32'h3d3dc5f0 /* (1, 12, 6) */,
  32'h3d19bf4b /* (29, 8, 6) */,
  32'h3d35cd98 /* (25, 8, 6) */,
  32'h3d865b59 /* (21, 8, 6) */,
  32'h3daa3349 /* (17, 8, 6) */,
  32'h3da2e7a9 /* (13, 8, 6) */,
  32'h3d584c0c /* (9, 8, 6) */,
  32'h3d22af34 /* (5, 8, 6) */,
  32'h3d169650 /* (1, 8, 6) */,
  32'h3d1b3fff /* (29, 4, 6) */,
  32'h3d17902e /* (25, 4, 6) */,
  32'h3d41fb9f /* (21, 4, 6) */,
  32'h3d61b1de /* (17, 4, 6) */,
  32'h3d601ae9 /* (13, 4, 6) */,
  32'h3d2657dd /* (9, 4, 6) */,
  32'h3d153e19 /* (5, 4, 6) */,
  32'h3d222a9c /* (1, 4, 6) */,
  32'h3d2d5b95 /* (29, 0, 6) */,
  32'h3d1459dd /* (25, 0, 6) */,
  32'h3d3013e2 /* (21, 0, 6) */,
  32'h3d455011 /* (17, 0, 6) */,
  32'h3d4703b2 /* (13, 0, 6) */,
  32'h3d1bc36a /* (9, 0, 6) */,
  32'h3d1b2f33 /* (5, 0, 6) */,
  32'h3d3f59b8 /* (1, 0, 6) */,
  32'h3d5defd3 /* (29, 28, 2) */,
  32'h3d16c6a3 /* (25, 28, 2) */,
  32'h3d21c128 /* (21, 28, 2) */,
  32'h3d2d6bba /* (17, 28, 2) */,
  32'h3d3217f4 /* (13, 28, 2) */,
  32'h3d14de35 /* (9, 28, 2) */,
  32'h3d2d8e0e /* (5, 28, 2) */,
  32'h3d8b1391 /* (1, 28, 2) */,
  32'h3d13e9f7 /* (29, 24, 2) */,
  32'h3d1d59b0 /* (25, 24, 2) */,
  32'h3d558b1c /* (21, 24, 2) */,
  32'h3d804df8 /* (17, 24, 2) */,
  32'h3d7b52f8 /* (13, 24, 2) */,
  32'h3d3291f6 /* (9, 24, 2) */,
  32'h3d149b5c /* (5, 24, 2) */,
  32'h3d15ce12 /* (1, 24, 2) */,
  32'h3d23d587 /* (29, 20, 2) */,
  32'h3d530d8e /* (25, 20, 2) */,
  32'h3da96c08 /* (21, 20, 2) */,
  32'h3de39dff /* (17, 20, 2) */,
  32'h3dd42d31 /* (13, 20, 2) */,
  32'h3d833332 /* (9, 20, 2) */,
  32'h3d346b02 /* (5, 20, 2) */,
  32'h3d1cac31 /* (1, 20, 2) */,
  32'h3d13661d /* (29, 16, 2) */,
  32'h3d4f6a6e /* (25, 16, 2) */,
  32'h3db86416 /* (21, 16, 2) */,
  32'h3e06ec2e /* (17, 16, 2) */,
  32'h3df1ae3d /* (13, 16, 2) */,
  32'h3d87d16b /* (9, 16, 2) */,
  32'h3d28d1e5 /* (5, 16, 2) */,
  32'h3d09dfab /* (1, 16, 2) */,
  32'h3d23d587 /* (29, 12, 2) */,
  32'h3d530d8e /* (25, 12, 2) */,
  32'h3da96c08 /* (21, 12, 2) */,
  32'h3de39dff /* (17, 12, 2) */,
  32'h3dd42d31 /* (13, 12, 2) */,
  32'h3d833332 /* (9, 12, 2) */,
  32'h3d346b02 /* (5, 12, 2) */,
  32'h3d1cac31 /* (1, 12, 2) */,
  32'h3d13e9f7 /* (29, 8, 2) */,
  32'h3d1d59b0 /* (25, 8, 2) */,
  32'h3d558b1c /* (21, 8, 2) */,
  32'h3d804df8 /* (17, 8, 2) */,
  32'h3d7b52f8 /* (13, 8, 2) */,
  32'h3d3291f6 /* (9, 8, 2) */,
  32'h3d149b5c /* (5, 8, 2) */,
  32'h3d15ce12 /* (1, 8, 2) */,
  32'h3d5defd3 /* (29, 4, 2) */,
  32'h3d16c6a3 /* (25, 4, 2) */,
  32'h3d21c128 /* (21, 4, 2) */,
  32'h3d2d6bba /* (17, 4, 2) */,
  32'h3d3217f4 /* (13, 4, 2) */,
  32'h3d14de35 /* (9, 4, 2) */,
  32'h3d2d8e0e /* (5, 4, 2) */,
  32'h3d8b1391 /* (1, 4, 2) */,
  32'h3dcbea25 /* (29, 0, 2) */,
  32'h3d21b235 /* (25, 0, 2) */,
  32'h3d164ce1 /* (21, 0, 2) */,
  32'h3d18d610 /* (17, 0, 2) */,
  32'h3d2045b1 /* (13, 0, 2) */,
  32'h3d11b684 /* (9, 0, 2) */,
  32'h3d5dd7d1 /* (5, 0, 2) */,
  32'h3e709592 /* (1, 0, 2) */,
  32'h3d429928 /* (28, 28, 30) */,
  32'h3d139519 /* (24, 28, 30) */,
  32'h3d2ab74a /* (20, 28, 30) */,
  32'h3d1c5e8a /* (16, 28, 30) */,
  32'h3d2ab74a /* (12, 28, 30) */,
  32'h3d139519 /* (8, 28, 30) */,
  32'h3d429928 /* (4, 28, 30) */,
  32'h3d90451b /* (0, 28, 30) */,
  32'h3d139519 /* (28, 24, 30) */,
  32'h3d263161 /* (24, 24, 30) */,
  32'h3d69b2a3 /* (20, 24, 30) */,
  32'h3d6bb726 /* (16, 24, 30) */,
  32'h3d69b2a3 /* (12, 24, 30) */,
  32'h3d263161 /* (8, 24, 30) */,
  32'h3d139519 /* (4, 24, 30) */,
  32'h3d162cf4 /* (0, 24, 30) */,
  32'h3d2ab74a /* (28, 20, 30) */,
  32'h3d69b2a3 /* (24, 20, 30) */,
  32'h3dbf980c /* (20, 20, 30) */,
  32'h3dd576ed /* (16, 20, 30) */,
  32'h3dbf980c /* (12, 20, 30) */,
  32'h3d69b2a3 /* (8, 20, 30) */,
  32'h3d2ab74a /* (4, 20, 30) */,
  32'h3d1bd472 /* (0, 20, 30) */,
  32'h3d1c5e8a /* (28, 16, 30) */,
  32'h3d6bb726 /* (24, 16, 30) */,
  32'h3dd576ed /* (20, 16, 30) */,
  32'h3e00d0e8 /* (16, 16, 30) */,
  32'h3dd576ed /* (12, 16, 30) */,
  32'h3d6bb726 /* (8, 16, 30) */,
  32'h3d1c5e8a /* (4, 16, 30) */,
  32'h3d08bc50 /* (0, 16, 30) */,
  32'h3d2ab74a /* (28, 12, 30) */,
  32'h3d69b2a3 /* (24, 12, 30) */,
  32'h3dbf980c /* (20, 12, 30) */,
  32'h3dd576ed /* (16, 12, 30) */,
  32'h3dbf980c /* (12, 12, 30) */,
  32'h3d69b2a3 /* (8, 12, 30) */,
  32'h3d2ab74a /* (4, 12, 30) */,
  32'h3d1bd472 /* (0, 12, 30) */,
  32'h3d139519 /* (28, 8, 30) */,
  32'h3d263161 /* (24, 8, 30) */,
  32'h3d69b2a3 /* (20, 8, 30) */,
  32'h3d6bb726 /* (16, 8, 30) */,
  32'h3d69b2a3 /* (12, 8, 30) */,
  32'h3d263161 /* (8, 8, 30) */,
  32'h3d139519 /* (4, 8, 30) */,
  32'h3d162cf4 /* (0, 8, 30) */,
  32'h3d429928 /* (28, 4, 30) */,
  32'h3d139519 /* (24, 4, 30) */,
  32'h3d2ab74a /* (20, 4, 30) */,
  32'h3d1c5e8a /* (16, 4, 30) */,
  32'h3d2ab74a /* (12, 4, 30) */,
  32'h3d139519 /* (8, 4, 30) */,
  32'h3d429928 /* (4, 4, 30) */,
  32'h3d90451b /* (0, 4, 30) */,
  32'h3d90451b /* (28, 0, 30) */,
  32'h3d162cf4 /* (24, 0, 30) */,
  32'h3d1bd472 /* (20, 0, 30) */,
  32'h3d08bc50 /* (16, 0, 30) */,
  32'h3d1bd472 /* (12, 0, 30) */,
  32'h3d162cf4 /* (8, 0, 30) */,
  32'h3d90451b /* (4, 0, 30) */,
  32'h3e948d77 /* (0, 0, 30) */,
  32'h3d1796af /* (28, 28, 26) */,
  32'h3d1d3fef /* (24, 28, 26) */,
  32'h3d522ea6 /* (20, 28, 26) */,
  32'h3d4e2dc2 /* (16, 28, 26) */,
  32'h3d522ea6 /* (12, 28, 26) */,
  32'h3d1d3fef /* (8, 28, 26) */,
  32'h3d1796af /* (4, 28, 26) */,
  32'h3d234ae8 /* (0, 28, 26) */,
  32'h3d1d3fef /* (28, 24, 26) */,
  32'h3d44d2c5 /* (24, 24, 26) */,
  32'h3d95625b /* (20, 24, 26) */,
  32'h3d9dd43f /* (16, 24, 26) */,
  32'h3d95625b /* (12, 24, 26) */,
  32'h3d44d2c5 /* (8, 24, 26) */,
  32'h3d1d3fef /* (4, 24, 26) */,
  32'h3d164277 /* (0, 24, 26) */,
  32'h3d522ea6 /* (28, 20, 26) */,
  32'h3d95625b /* (24, 20, 26) */,
  32'h3dfe11f4 /* (20, 20, 26) */,
  32'h3e11854b /* (16, 20, 26) */,
  32'h3dfe11f4 /* (12, 20, 26) */,
  32'h3d95625b /* (8, 20, 26) */,
  32'h3d522ea6 /* (4, 20, 26) */,
  32'h3d3c86f4 /* (0, 20, 26) */,
  32'h3d4e2dc2 /* (28, 16, 26) */,
  32'h3d9dd43f /* (24, 16, 26) */,
  32'h3e11854b /* (20, 16, 26) */,
  32'h3e327927 /* (16, 16, 26) */,
  32'h3e11854b /* (12, 16, 26) */,
  32'h3d9dd43f /* (8, 16, 26) */,
  32'h3d4e2dc2 /* (4, 16, 26) */,
  32'h3d332545 /* (0, 16, 26) */,
  32'h3d522ea6 /* (28, 12, 26) */,
  32'h3d95625b /* (24, 12, 26) */,
  32'h3dfe11f4 /* (20, 12, 26) */,
  32'h3e11854b /* (16, 12, 26) */,
  32'h3dfe11f4 /* (12, 12, 26) */,
  32'h3d95625b /* (8, 12, 26) */,
  32'h3d522ea6 /* (4, 12, 26) */,
  32'h3d3c86f4 /* (0, 12, 26) */,
  32'h3d1d3fef /* (28, 8, 26) */,
  32'h3d44d2c5 /* (24, 8, 26) */,
  32'h3d95625b /* (20, 8, 26) */,
  32'h3d9dd43f /* (16, 8, 26) */,
  32'h3d95625b /* (12, 8, 26) */,
  32'h3d44d2c5 /* (8, 8, 26) */,
  32'h3d1d3fef /* (4, 8, 26) */,
  32'h3d164277 /* (0, 8, 26) */,
  32'h3d1796af /* (28, 4, 26) */,
  32'h3d1d3fef /* (24, 4, 26) */,
  32'h3d522ea6 /* (20, 4, 26) */,
  32'h3d4e2dc2 /* (16, 4, 26) */,
  32'h3d522ea6 /* (12, 4, 26) */,
  32'h3d1d3fef /* (8, 4, 26) */,
  32'h3d1796af /* (4, 4, 26) */,
  32'h3d234ae8 /* (0, 4, 26) */,
  32'h3d234ae8 /* (28, 0, 26) */,
  32'h3d164277 /* (24, 0, 26) */,
  32'h3d3c86f4 /* (20, 0, 26) */,
  32'h3d332545 /* (16, 0, 26) */,
  32'h3d3c86f4 /* (12, 0, 26) */,
  32'h3d164277 /* (8, 0, 26) */,
  32'h3d234ae8 /* (4, 0, 26) */,
  32'h3d424b89 /* (0, 0, 26) */,
  32'h3d21d2a4 /* (28, 28, 22) */,
  32'h3d51ff4c /* (24, 28, 22) */,
  32'h3da42ada /* (20, 28, 22) */,
  32'h3db0df4f /* (16, 28, 22) */,
  32'h3da42ada /* (12, 28, 22) */,
  32'h3d51ff4c /* (8, 28, 22) */,
  32'h3d21d2a4 /* (4, 28, 22) */,
  32'h3d17b006 /* (0, 28, 22) */,
  32'h3d51ff4c /* (28, 24, 22) */,
  32'h3d92b00e /* (24, 24, 22) */,
  32'h3df53c17 /* (20, 24, 22) */,
  32'h3e0a9c46 /* (16, 24, 22) */,
  32'h3df53c17 /* (12, 24, 22) */,
  32'h3d92b00e /* (8, 24, 22) */,
  32'h3d51ff4c /* (4, 24, 22) */,
  32'h3d3ddc84 /* (0, 24, 22) */,
  32'h3da42ada /* (28, 20, 22) */,
  32'h3df53c17 /* (24, 20, 22) */,
  32'h3e5bd2f1 /* (20, 20, 22) */,
  32'h3e837a14 /* (16, 20, 22) */,
  32'h3e5bd2f1 /* (12, 20, 22) */,
  32'h3df53c17 /* (8, 20, 22) */,
  32'h3da42ada /* (4, 20, 22) */,
  32'h3d9019ab /* (0, 20, 22) */,
  32'h3db0df4f /* (28, 16, 22) */,
  32'h3e0a9c46 /* (24, 16, 22) */,
  32'h3e837a14 /* (20, 16, 22) */,
  32'h3ea594bb /* (16, 16, 22) */,
  32'h3e837a14 /* (12, 16, 22) */,
  32'h3e0a9c46 /* (8, 16, 22) */,
  32'h3db0df4f /* (4, 16, 22) */,
  32'h3d983f17 /* (0, 16, 22) */,
  32'h3da42ada /* (28, 12, 22) */,
  32'h3df53c17 /* (24, 12, 22) */,
  32'h3e5bd2f1 /* (20, 12, 22) */,
  32'h3e837a14 /* (16, 12, 22) */,
  32'h3e5bd2f1 /* (12, 12, 22) */,
  32'h3df53c17 /* (8, 12, 22) */,
  32'h3da42ada /* (4, 12, 22) */,
  32'h3d9019ab /* (0, 12, 22) */,
  32'h3d51ff4c /* (28, 8, 22) */,
  32'h3d92b00e /* (24, 8, 22) */,
  32'h3df53c17 /* (20, 8, 22) */,
  32'h3e0a9c46 /* (16, 8, 22) */,
  32'h3df53c17 /* (12, 8, 22) */,
  32'h3d92b00e /* (8, 8, 22) */,
  32'h3d51ff4c /* (4, 8, 22) */,
  32'h3d3ddc84 /* (0, 8, 22) */,
  32'h3d21d2a4 /* (28, 4, 22) */,
  32'h3d51ff4c /* (24, 4, 22) */,
  32'h3da42ada /* (20, 4, 22) */,
  32'h3db0df4f /* (16, 4, 22) */,
  32'h3da42ada /* (12, 4, 22) */,
  32'h3d51ff4c /* (8, 4, 22) */,
  32'h3d21d2a4 /* (4, 4, 22) */,
  32'h3d17b006 /* (0, 4, 22) */,
  32'h3d17b006 /* (28, 0, 22) */,
  32'h3d3ddc84 /* (24, 0, 22) */,
  32'h3d9019ab /* (20, 0, 22) */,
  32'h3d983f17 /* (16, 0, 22) */,
  32'h3d9019ab /* (12, 0, 22) */,
  32'h3d3ddc84 /* (8, 0, 22) */,
  32'h3d17b006 /* (4, 0, 22) */,
  32'h3d10f1da /* (0, 0, 22) */,
  32'h3d456b70 /* (28, 28, 18) */,
  32'h3d904c26 /* (24, 28, 18) */,
  32'h3dfca6c8 /* (20, 28, 18) */,
  32'h3e1420e4 /* (16, 28, 18) */,
  32'h3dfca6c8 /* (12, 28, 18) */,
  32'h3d904c26 /* (8, 28, 18) */,
  32'h3d456b70 /* (4, 28, 18) */,
  32'h3d2ee5c8 /* (0, 28, 18) */,
  32'h3d904c26 /* (28, 24, 18) */,
  32'h3dd9849b /* (24, 24, 18) */,
  32'h3e44fc23 /* (20, 24, 18) */,
  32'h3e6dbe20 /* (16, 24, 18) */,
  32'h3e44fc23 /* (12, 24, 18) */,
  32'h3dd9849b /* (8, 24, 18) */,
  32'h3d904c26 /* (4, 24, 18) */,
  32'h3d7c5be6 /* (0, 24, 18) */,
  32'h3dfca6c8 /* (28, 20, 18) */,
  32'h3e44fc23 /* (24, 20, 18) */,
  32'h3eb9abaa /* (20, 20, 18) */,
  32'h3ee86d0e /* (16, 20, 18) */,
  32'h3eb9abaa /* (12, 20, 18) */,
  32'h3e44fc23 /* (8, 20, 18) */,
  32'h3dfca6c8 /* (4, 20, 18) */,
  32'h3dd9ea44 /* (0, 20, 18) */,
  32'h3e1420e4 /* (28, 16, 18) */,
  32'h3e6dbe20 /* (24, 16, 18) */,
  32'h3ee86d0e /* (20, 16, 18) */,
  32'h3f16cd97 /* (16, 16, 18) */,
  32'h3ee86d0e /* (12, 16, 18) */,
  32'h3e6dbe20 /* (8, 16, 18) */,
  32'h3e1420e4 /* (4, 16, 18) */,
  32'h3dfcae00 /* (0, 16, 18) */,
  32'h3dfca6c8 /* (28, 12, 18) */,
  32'h3e44fc23 /* (24, 12, 18) */,
  32'h3eb9abaa /* (20, 12, 18) */,
  32'h3ee86d0e /* (16, 12, 18) */,
  32'h3eb9abaa /* (12, 12, 18) */,
  32'h3e44fc23 /* (8, 12, 18) */,
  32'h3dfca6c8 /* (4, 12, 18) */,
  32'h3dd9ea44 /* (0, 12, 18) */,
  32'h3d904c26 /* (28, 8, 18) */,
  32'h3dd9849b /* (24, 8, 18) */,
  32'h3e44fc23 /* (20, 8, 18) */,
  32'h3e6dbe20 /* (16, 8, 18) */,
  32'h3e44fc23 /* (12, 8, 18) */,
  32'h3dd9849b /* (8, 8, 18) */,
  32'h3d904c26 /* (4, 8, 18) */,
  32'h3d7c5be6 /* (0, 8, 18) */,
  32'h3d456b70 /* (28, 4, 18) */,
  32'h3d904c26 /* (24, 4, 18) */,
  32'h3dfca6c8 /* (20, 4, 18) */,
  32'h3e1420e4 /* (16, 4, 18) */,
  32'h3dfca6c8 /* (12, 4, 18) */,
  32'h3d904c26 /* (8, 4, 18) */,
  32'h3d456b70 /* (4, 4, 18) */,
  32'h3d2ee5c8 /* (0, 4, 18) */,
  32'h3d2ee5c8 /* (28, 0, 18) */,
  32'h3d7c5be6 /* (24, 0, 18) */,
  32'h3dd9ea44 /* (20, 0, 18) */,
  32'h3dfcae00 /* (16, 0, 18) */,
  32'h3dd9ea44 /* (12, 0, 18) */,
  32'h3d7c5be6 /* (8, 0, 18) */,
  32'h3d2ee5c8 /* (4, 0, 18) */,
  32'h3d1bd51d /* (0, 0, 18) */,
  32'h3d456b70 /* (28, 28, 14) */,
  32'h3d904c26 /* (24, 28, 14) */,
  32'h3dfca6c8 /* (20, 28, 14) */,
  32'h3e1420e4 /* (16, 28, 14) */,
  32'h3dfca6c8 /* (12, 28, 14) */,
  32'h3d904c26 /* (8, 28, 14) */,
  32'h3d456b70 /* (4, 28, 14) */,
  32'h3d2ee5c8 /* (0, 28, 14) */,
  32'h3d904c26 /* (28, 24, 14) */,
  32'h3dd9849b /* (24, 24, 14) */,
  32'h3e44fc23 /* (20, 24, 14) */,
  32'h3e6dbe20 /* (16, 24, 14) */,
  32'h3e44fc23 /* (12, 24, 14) */,
  32'h3dd9849b /* (8, 24, 14) */,
  32'h3d904c26 /* (4, 24, 14) */,
  32'h3d7c5be6 /* (0, 24, 14) */,
  32'h3dfca6c8 /* (28, 20, 14) */,
  32'h3e44fc23 /* (24, 20, 14) */,
  32'h3eb9abaa /* (20, 20, 14) */,
  32'h3ee86d0e /* (16, 20, 14) */,
  32'h3eb9abaa /* (12, 20, 14) */,
  32'h3e44fc23 /* (8, 20, 14) */,
  32'h3dfca6c8 /* (4, 20, 14) */,
  32'h3dd9ea44 /* (0, 20, 14) */,
  32'h3e1420e4 /* (28, 16, 14) */,
  32'h3e6dbe20 /* (24, 16, 14) */,
  32'h3ee86d0e /* (20, 16, 14) */,
  32'h3f16cd97 /* (16, 16, 14) */,
  32'h3ee86d0e /* (12, 16, 14) */,
  32'h3e6dbe20 /* (8, 16, 14) */,
  32'h3e1420e4 /* (4, 16, 14) */,
  32'h3dfcae00 /* (0, 16, 14) */,
  32'h3dfca6c8 /* (28, 12, 14) */,
  32'h3e44fc23 /* (24, 12, 14) */,
  32'h3eb9abaa /* (20, 12, 14) */,
  32'h3ee86d0e /* (16, 12, 14) */,
  32'h3eb9abaa /* (12, 12, 14) */,
  32'h3e44fc23 /* (8, 12, 14) */,
  32'h3dfca6c8 /* (4, 12, 14) */,
  32'h3dd9ea44 /* (0, 12, 14) */,
  32'h3d904c26 /* (28, 8, 14) */,
  32'h3dd9849b /* (24, 8, 14) */,
  32'h3e44fc23 /* (20, 8, 14) */,
  32'h3e6dbe20 /* (16, 8, 14) */,
  32'h3e44fc23 /* (12, 8, 14) */,
  32'h3dd9849b /* (8, 8, 14) */,
  32'h3d904c26 /* (4, 8, 14) */,
  32'h3d7c5be6 /* (0, 8, 14) */,
  32'h3d456b70 /* (28, 4, 14) */,
  32'h3d904c26 /* (24, 4, 14) */,
  32'h3dfca6c8 /* (20, 4, 14) */,
  32'h3e1420e4 /* (16, 4, 14) */,
  32'h3dfca6c8 /* (12, 4, 14) */,
  32'h3d904c26 /* (8, 4, 14) */,
  32'h3d456b70 /* (4, 4, 14) */,
  32'h3d2ee5c8 /* (0, 4, 14) */,
  32'h3d2ee5c8 /* (28, 0, 14) */,
  32'h3d7c5be6 /* (24, 0, 14) */,
  32'h3dd9ea44 /* (20, 0, 14) */,
  32'h3dfcae00 /* (16, 0, 14) */,
  32'h3dd9ea44 /* (12, 0, 14) */,
  32'h3d7c5be6 /* (8, 0, 14) */,
  32'h3d2ee5c8 /* (4, 0, 14) */,
  32'h3d1bd51d /* (0, 0, 14) */,
  32'h3d21d2a4 /* (28, 28, 10) */,
  32'h3d51ff4c /* (24, 28, 10) */,
  32'h3da42ada /* (20, 28, 10) */,
  32'h3db0df4f /* (16, 28, 10) */,
  32'h3da42ada /* (12, 28, 10) */,
  32'h3d51ff4c /* (8, 28, 10) */,
  32'h3d21d2a4 /* (4, 28, 10) */,
  32'h3d17b006 /* (0, 28, 10) */,
  32'h3d51ff4c /* (28, 24, 10) */,
  32'h3d92b00e /* (24, 24, 10) */,
  32'h3df53c17 /* (20, 24, 10) */,
  32'h3e0a9c46 /* (16, 24, 10) */,
  32'h3df53c17 /* (12, 24, 10) */,
  32'h3d92b00e /* (8, 24, 10) */,
  32'h3d51ff4c /* (4, 24, 10) */,
  32'h3d3ddc84 /* (0, 24, 10) */,
  32'h3da42ada /* (28, 20, 10) */,
  32'h3df53c17 /* (24, 20, 10) */,
  32'h3e5bd2f1 /* (20, 20, 10) */,
  32'h3e837a14 /* (16, 20, 10) */,
  32'h3e5bd2f1 /* (12, 20, 10) */,
  32'h3df53c17 /* (8, 20, 10) */,
  32'h3da42ada /* (4, 20, 10) */,
  32'h3d9019ab /* (0, 20, 10) */,
  32'h3db0df4f /* (28, 16, 10) */,
  32'h3e0a9c46 /* (24, 16, 10) */,
  32'h3e837a14 /* (20, 16, 10) */,
  32'h3ea594bb /* (16, 16, 10) */,
  32'h3e837a14 /* (12, 16, 10) */,
  32'h3e0a9c46 /* (8, 16, 10) */,
  32'h3db0df4f /* (4, 16, 10) */,
  32'h3d983f17 /* (0, 16, 10) */,
  32'h3da42ada /* (28, 12, 10) */,
  32'h3df53c17 /* (24, 12, 10) */,
  32'h3e5bd2f1 /* (20, 12, 10) */,
  32'h3e837a14 /* (16, 12, 10) */,
  32'h3e5bd2f1 /* (12, 12, 10) */,
  32'h3df53c17 /* (8, 12, 10) */,
  32'h3da42ada /* (4, 12, 10) */,
  32'h3d9019ab /* (0, 12, 10) */,
  32'h3d51ff4c /* (28, 8, 10) */,
  32'h3d92b00e /* (24, 8, 10) */,
  32'h3df53c17 /* (20, 8, 10) */,
  32'h3e0a9c46 /* (16, 8, 10) */,
  32'h3df53c17 /* (12, 8, 10) */,
  32'h3d92b00e /* (8, 8, 10) */,
  32'h3d51ff4c /* (4, 8, 10) */,
  32'h3d3ddc84 /* (0, 8, 10) */,
  32'h3d21d2a4 /* (28, 4, 10) */,
  32'h3d51ff4c /* (24, 4, 10) */,
  32'h3da42ada /* (20, 4, 10) */,
  32'h3db0df4f /* (16, 4, 10) */,
  32'h3da42ada /* (12, 4, 10) */,
  32'h3d51ff4c /* (8, 4, 10) */,
  32'h3d21d2a4 /* (4, 4, 10) */,
  32'h3d17b006 /* (0, 4, 10) */,
  32'h3d17b006 /* (28, 0, 10) */,
  32'h3d3ddc84 /* (24, 0, 10) */,
  32'h3d9019ab /* (20, 0, 10) */,
  32'h3d983f17 /* (16, 0, 10) */,
  32'h3d9019ab /* (12, 0, 10) */,
  32'h3d3ddc84 /* (8, 0, 10) */,
  32'h3d17b006 /* (4, 0, 10) */,
  32'h3d10f1da /* (0, 0, 10) */,
  32'h3d1796af /* (28, 28, 6) */,
  32'h3d1d3fef /* (24, 28, 6) */,
  32'h3d522ea6 /* (20, 28, 6) */,
  32'h3d4e2dc2 /* (16, 28, 6) */,
  32'h3d522ea6 /* (12, 28, 6) */,
  32'h3d1d3fef /* (8, 28, 6) */,
  32'h3d1796af /* (4, 28, 6) */,
  32'h3d234ae8 /* (0, 28, 6) */,
  32'h3d1d3fef /* (28, 24, 6) */,
  32'h3d44d2c5 /* (24, 24, 6) */,
  32'h3d95625b /* (20, 24, 6) */,
  32'h3d9dd43f /* (16, 24, 6) */,
  32'h3d95625b /* (12, 24, 6) */,
  32'h3d44d2c5 /* (8, 24, 6) */,
  32'h3d1d3fef /* (4, 24, 6) */,
  32'h3d164277 /* (0, 24, 6) */,
  32'h3d522ea6 /* (28, 20, 6) */,
  32'h3d95625b /* (24, 20, 6) */,
  32'h3dfe11f4 /* (20, 20, 6) */,
  32'h3e11854b /* (16, 20, 6) */,
  32'h3dfe11f4 /* (12, 20, 6) */,
  32'h3d95625b /* (8, 20, 6) */,
  32'h3d522ea6 /* (4, 20, 6) */,
  32'h3d3c86f4 /* (0, 20, 6) */,
  32'h3d4e2dc2 /* (28, 16, 6) */,
  32'h3d9dd43f /* (24, 16, 6) */,
  32'h3e11854b /* (20, 16, 6) */,
  32'h3e327927 /* (16, 16, 6) */,
  32'h3e11854b /* (12, 16, 6) */,
  32'h3d9dd43f /* (8, 16, 6) */,
  32'h3d4e2dc2 /* (4, 16, 6) */,
  32'h3d332545 /* (0, 16, 6) */,
  32'h3d522ea6 /* (28, 12, 6) */,
  32'h3d95625b /* (24, 12, 6) */,
  32'h3dfe11f4 /* (20, 12, 6) */,
  32'h3e11854b /* (16, 12, 6) */,
  32'h3dfe11f4 /* (12, 12, 6) */,
  32'h3d95625b /* (8, 12, 6) */,
  32'h3d522ea6 /* (4, 12, 6) */,
  32'h3d3c86f4 /* (0, 12, 6) */,
  32'h3d1d3fef /* (28, 8, 6) */,
  32'h3d44d2c5 /* (24, 8, 6) */,
  32'h3d95625b /* (20, 8, 6) */,
  32'h3d9dd43f /* (16, 8, 6) */,
  32'h3d95625b /* (12, 8, 6) */,
  32'h3d44d2c5 /* (8, 8, 6) */,
  32'h3d1d3fef /* (4, 8, 6) */,
  32'h3d164277 /* (0, 8, 6) */,
  32'h3d1796af /* (28, 4, 6) */,
  32'h3d1d3fef /* (24, 4, 6) */,
  32'h3d522ea6 /* (20, 4, 6) */,
  32'h3d4e2dc2 /* (16, 4, 6) */,
  32'h3d522ea6 /* (12, 4, 6) */,
  32'h3d1d3fef /* (8, 4, 6) */,
  32'h3d1796af /* (4, 4, 6) */,
  32'h3d234ae8 /* (0, 4, 6) */,
  32'h3d234ae8 /* (28, 0, 6) */,
  32'h3d164277 /* (24, 0, 6) */,
  32'h3d3c86f4 /* (20, 0, 6) */,
  32'h3d332545 /* (16, 0, 6) */,
  32'h3d3c86f4 /* (12, 0, 6) */,
  32'h3d164277 /* (8, 0, 6) */,
  32'h3d234ae8 /* (4, 0, 6) */,
  32'h3d424b89 /* (0, 0, 6) */,
  32'h3d429928 /* (28, 28, 2) */,
  32'h3d139519 /* (24, 28, 2) */,
  32'h3d2ab74a /* (20, 28, 2) */,
  32'h3d1c5e8a /* (16, 28, 2) */,
  32'h3d2ab74a /* (12, 28, 2) */,
  32'h3d139519 /* (8, 28, 2) */,
  32'h3d429928 /* (4, 28, 2) */,
  32'h3d90451b /* (0, 28, 2) */,
  32'h3d139519 /* (28, 24, 2) */,
  32'h3d263161 /* (24, 24, 2) */,
  32'h3d69b2a3 /* (20, 24, 2) */,
  32'h3d6bb726 /* (16, 24, 2) */,
  32'h3d69b2a3 /* (12, 24, 2) */,
  32'h3d263161 /* (8, 24, 2) */,
  32'h3d139519 /* (4, 24, 2) */,
  32'h3d162cf4 /* (0, 24, 2) */,
  32'h3d2ab74a /* (28, 20, 2) */,
  32'h3d69b2a3 /* (24, 20, 2) */,
  32'h3dbf980c /* (20, 20, 2) */,
  32'h3dd576ed /* (16, 20, 2) */,
  32'h3dbf980c /* (12, 20, 2) */,
  32'h3d69b2a3 /* (8, 20, 2) */,
  32'h3d2ab74a /* (4, 20, 2) */,
  32'h3d1bd472 /* (0, 20, 2) */,
  32'h3d1c5e8a /* (28, 16, 2) */,
  32'h3d6bb726 /* (24, 16, 2) */,
  32'h3dd576ed /* (20, 16, 2) */,
  32'h3e00d0e8 /* (16, 16, 2) */,
  32'h3dd576ed /* (12, 16, 2) */,
  32'h3d6bb726 /* (8, 16, 2) */,
  32'h3d1c5e8a /* (4, 16, 2) */,
  32'h3d08bc50 /* (0, 16, 2) */,
  32'h3d2ab74a /* (28, 12, 2) */,
  32'h3d69b2a3 /* (24, 12, 2) */,
  32'h3dbf980c /* (20, 12, 2) */,
  32'h3dd576ed /* (16, 12, 2) */,
  32'h3dbf980c /* (12, 12, 2) */,
  32'h3d69b2a3 /* (8, 12, 2) */,
  32'h3d2ab74a /* (4, 12, 2) */,
  32'h3d1bd472 /* (0, 12, 2) */,
  32'h3d139519 /* (28, 8, 2) */,
  32'h3d263161 /* (24, 8, 2) */,
  32'h3d69b2a3 /* (20, 8, 2) */,
  32'h3d6bb726 /* (16, 8, 2) */,
  32'h3d69b2a3 /* (12, 8, 2) */,
  32'h3d263161 /* (8, 8, 2) */,
  32'h3d139519 /* (4, 8, 2) */,
  32'h3d162cf4 /* (0, 8, 2) */,
  32'h3d429928 /* (28, 4, 2) */,
  32'h3d139519 /* (24, 4, 2) */,
  32'h3d2ab74a /* (20, 4, 2) */,
  32'h3d1c5e8a /* (16, 4, 2) */,
  32'h3d2ab74a /* (12, 4, 2) */,
  32'h3d139519 /* (8, 4, 2) */,
  32'h3d429928 /* (4, 4, 2) */,
  32'h3d90451b /* (0, 4, 2) */,
  32'h3d90451b /* (28, 0, 2) */,
  32'h3d162cf4 /* (24, 0, 2) */,
  32'h3d1bd472 /* (20, 0, 2) */,
  32'h3d08bc50 /* (16, 0, 2) */,
  32'h3d1bd472 /* (12, 0, 2) */,
  32'h3d162cf4 /* (8, 0, 2) */,
  32'h3d90451b /* (4, 0, 2) */,
  32'h3e948d77 /* (0, 0, 2) */,
  32'h3deb372d /* (31, 31, 29) */,
  32'h3d45ae9a /* (27, 31, 29) */,
  32'h3d126006 /* (23, 31, 29) */,
  32'h3d269671 /* (19, 31, 29) */,
  32'h3d202be8 /* (15, 31, 29) */,
  32'h3d1a3ccf /* (11, 31, 29) */,
  32'h3d1c3652 /* (7, 31, 29) */,
  32'h3d960c3c /* (3, 31, 29) */,
  32'h3d45ae9a /* (31, 27, 29) */,
  32'h3d1ccb4c /* (27, 27, 29) */,
  32'h3d1addce /* (23, 27, 29) */,
  32'h3d4466f8 /* (19, 27, 29) */,
  32'h3d424fe8 /* (15, 27, 29) */,
  32'h3d2e4aa1 /* (11, 27, 29) */,
  32'h3d147808 /* (7, 27, 29) */,
  32'h3d314afb /* (3, 27, 29) */,
  32'h3d126006 /* (31, 23, 29) */,
  32'h3d1addce /* (27, 23, 29) */,
  32'h3d48821f /* (23, 23, 29) */,
  32'h3d942dc4 /* (19, 23, 29) */,
  32'h3d99caa3 /* (15, 23, 29) */,
  32'h3d767d5d /* (11, 23, 29) */,
  32'h3d2aad03 /* (7, 23, 29) */,
  32'h3d144047 /* (3, 23, 29) */,
  32'h3d269671 /* (31, 19, 29) */,
  32'h3d4466f8 /* (27, 19, 29) */,
  32'h3d942dc4 /* (23, 19, 29) */,
  32'h3df79892 /* (19, 19, 29) */,
  32'h3e068db8 /* (15, 19, 29) */,
  32'h3dc2b35d /* (11, 19, 29) */,
  32'h3d69f6ae /* (7, 19, 29) */,
  32'h3d2fb3ed /* (3, 19, 29) */,
  32'h3d202be8 /* (31, 15, 29) */,
  32'h3d424fe8 /* (27, 15, 29) */,
  32'h3d99caa3 /* (23, 15, 29) */,
  32'h3e068db8 /* (19, 15, 29) */,
  32'h3e151f83 /* (15, 15, 29) */,
  32'h3dceffa6 /* (11, 15, 29) */,
  32'h3d6ce397 /* (7, 15, 29) */,
  32'h3d2aacf2 /* (3, 15, 29) */,
  32'h3d1a3ccf /* (31, 11, 29) */,
  32'h3d2e4aa1 /* (27, 11, 29) */,
  32'h3d767d5d /* (23, 11, 29) */,
  32'h3dc2b35d /* (19, 11, 29) */,
  32'h3dceffa6 /* (15, 11, 29) */,
  32'h3d9d27e1 /* (11, 11, 29) */,
  32'h3d490aba /* (7, 11, 29) */,
  32'h3d202a91 /* (3, 11, 29) */,
  32'h3d1c3652 /* (31, 7, 29) */,
  32'h3d147808 /* (27, 7, 29) */,
  32'h3d2aad03 /* (23, 7, 29) */,
  32'h3d69f6ae /* (19, 7, 29) */,
  32'h3d6ce397 /* (15, 7, 29) */,
  32'h3d490aba /* (11, 7, 29) */,
  32'h3d1969a9 /* (7, 7, 29) */,
  32'h3d179239 /* (3, 7, 29) */,
  32'h3d960c3c /* (31, 3, 29) */,
  32'h3d314afb /* (27, 3, 29) */,
  32'h3d144047 /* (23, 3, 29) */,
  32'h3d2fb3ed /* (19, 3, 29) */,
  32'h3d2aacf2 /* (15, 3, 29) */,
  32'h3d202a91 /* (11, 3, 29) */,
  32'h3d179239 /* (7, 3, 29) */,
  32'h3d68b01f /* (3, 3, 29) */,
  32'h3d2402bf /* (31, 31, 25) */,
  32'h3d151e01 /* (27, 31, 25) */,
  32'h3d245baa /* (23, 31, 25) */,
  32'h3d5c17b6 /* (19, 31, 25) */,
  32'h3d5d3ed0 /* (15, 31, 25) */,
  32'h3d3efe62 /* (11, 31, 25) */,
  32'h3d167b79 /* (7, 31, 25) */,
  32'h3d1c3652 /* (3, 31, 25) */,
  32'h3d151e01 /* (31, 27, 25) */,
  32'h3d170afd /* (27, 27, 25) */,
  32'h3d39ba58 /* (23, 27, 25) */,
  32'h3d849ae2 /* (19, 27, 25) */,
  32'h3d880917 /* (15, 27, 25) */,
  32'h3d5ff008 /* (11, 27, 25) */,
  32'h3d21f168 /* (7, 27, 25) */,
  32'h3d147808 /* (3, 27, 25) */,
  32'h3d245baa /* (31, 23, 25) */,
  32'h3d39ba58 /* (27, 23, 25) */,
  32'h3d8354ed /* (23, 23, 25) */,
  32'h3dcf79e9 /* (19, 23, 25) */,
  32'h3ddc94c6 /* (15, 23, 25) */,
  32'h3da777c1 /* (11, 23, 25) */,
  32'h3d563bcb /* (7, 23, 25) */,
  32'h3d2aad03 /* (3, 23, 25) */,
  32'h3d5c17b6 /* (31, 19, 25) */,
  32'h3d849ae2 /* (27, 19, 25) */,
  32'h3dcf79e9 /* (23, 19, 25) */,
  32'h3e336d1b /* (19, 19, 25) */,
  32'h3e45db44 /* (15, 19, 25) */,
  32'h3e0aca9a /* (11, 19, 25) */,
  32'h3da0c360 /* (7, 19, 25) */,
  32'h3d69f6ae /* (3, 19, 25) */,
  32'h3d5d3ed0 /* (31, 15, 25) */,
  32'h3d880917 /* (27, 15, 25) */,
  32'h3ddc94c6 /* (23, 15, 25) */,
  32'h3e45db44 /* (19, 15, 25) */,
  32'h3e5db918 /* (15, 15, 25) */,
  32'h3e165b49 /* (11, 15, 25) */,
  32'h3da7bf05 /* (7, 15, 25) */,
  32'h3d6ce397 /* (3, 15, 25) */,
  32'h3d3efe62 /* (31, 11, 25) */,
  32'h3d5ff008 /* (27, 11, 25) */,
  32'h3da777c1 /* (23, 11, 25) */,
  32'h3e0aca9a /* (19, 11, 25) */,
  32'h3e165b49 /* (15, 11, 25) */,
  32'h3ddb1c7f /* (11, 11, 25) */,
  32'h3d84ce75 /* (7, 11, 25) */,
  32'h3d490aba /* (3, 11, 25) */,
  32'h3d167b79 /* (31, 7, 25) */,
  32'h3d21f168 /* (27, 7, 25) */,
  32'h3d563bcb /* (23, 7, 25) */,
  32'h3da0c360 /* (19, 7, 25) */,
  32'h3da7bf05 /* (15, 7, 25) */,
  32'h3d84ce75 /* (11, 7, 25) */,
  32'h3d348078 /* (7, 7, 25) */,
  32'h3d1969a9 /* (3, 7, 25) */,
  32'h3d1c3652 /* (31, 3, 25) */,
  32'h3d147808 /* (27, 3, 25) */,
  32'h3d2aad03 /* (23, 3, 25) */,
  32'h3d69f6ae /* (19, 3, 25) */,
  32'h3d6ce397 /* (15, 3, 25) */,
  32'h3d490aba /* (11, 3, 25) */,
  32'h3d1969a9 /* (7, 3, 25) */,
  32'h3d179239 /* (3, 3, 25) */,
  32'h3d151591 /* (31, 31, 21) */,
  32'h3d26c9db /* (27, 31, 21) */,
  32'h3d68852c /* (23, 31, 21) */,
  32'h3db58f74 /* (19, 31, 21) */,
  32'h3dc031e4 /* (15, 31, 21) */,
  32'h3d9352ec /* (11, 31, 21) */,
  32'h3d3efe62 /* (7, 31, 21) */,
  32'h3d1a3ccf /* (3, 31, 21) */,
  32'h3d26c9db /* (31, 27, 21) */,
  32'h3d3fb488 /* (27, 27, 21) */,
  32'h3d8b02ad /* (23, 27, 21) */,
  32'h3de04254 /* (19, 27, 21) */,
  32'h3df05994 /* (15, 27, 21) */,
  32'h3db345e2 /* (11, 27, 21) */,
  32'h3d5ff008 /* (7, 27, 21) */,
  32'h3d2e4aa1 /* (3, 27, 21) */,
  32'h3d68852c /* (31, 23, 21) */,
  32'h3d8b02ad /* (27, 23, 21) */,
  32'h3dd6aa1b /* (23, 23, 21) */,
  32'h3e37494b /* (19, 23, 21) */,
  32'h3e49046a /* (15, 23, 21) */,
  32'h3e0ea5fd /* (11, 23, 21) */,
  32'h3da777c1 /* (7, 23, 21) */,
  32'h3d767d5d /* (3, 23, 21) */,
  32'h3db58f74 /* (31, 19, 21) */,
  32'h3de04254 /* (27, 19, 21) */,
  32'h3e37494b /* (23, 19, 21) */,
  32'h3ea5d30f /* (19, 19, 21) */,
  32'h3eba8e90 /* (15, 19, 21) */,
  32'h3e7af74d /* (11, 19, 21) */,
  32'h3e0aca9a /* (7, 19, 21) */,
  32'h3dc2b35d /* (3, 19, 21) */,
  32'h3dc031e4 /* (31, 15, 21) */,
  32'h3df05994 /* (27, 15, 21) */,
  32'h3e49046a /* (23, 15, 21) */,
  32'h3eba8e90 /* (19, 15, 21) */,
  32'h3ed4648a /* (15, 15, 21) */,
  32'h3e8b66c2 /* (11, 15, 21) */,
  32'h3e165b49 /* (7, 15, 21) */,
  32'h3dceffa6 /* (3, 15, 21) */,
  32'h3d9352ec /* (31, 11, 21) */,
  32'h3db345e2 /* (27, 11, 21) */,
  32'h3e0ea5fd /* (23, 11, 21) */,
  32'h3e7af74d /* (19, 11, 21) */,
  32'h3e8b66c2 /* (15, 11, 21) */,
  32'h3e4089a2 /* (11, 11, 21) */,
  32'h3ddb1c7f /* (7, 11, 21) */,
  32'h3d9d27e1 /* (3, 11, 21) */,
  32'h3d3efe62 /* (31, 7, 21) */,
  32'h3d5ff008 /* (27, 7, 21) */,
  32'h3da777c1 /* (23, 7, 21) */,
  32'h3e0aca9a /* (19, 7, 21) */,
  32'h3e165b49 /* (15, 7, 21) */,
  32'h3ddb1c7f /* (11, 7, 21) */,
  32'h3d84ce75 /* (7, 7, 21) */,
  32'h3d490aba /* (3, 7, 21) */,
  32'h3d1a3ccf /* (31, 3, 21) */,
  32'h3d2e4aa1 /* (27, 3, 21) */,
  32'h3d767d5d /* (23, 3, 21) */,
  32'h3dc2b35d /* (19, 3, 21) */,
  32'h3dceffa6 /* (15, 3, 21) */,
  32'h3d9d27e1 /* (11, 3, 21) */,
  32'h3d490aba /* (7, 3, 21) */,
  32'h3d202a91 /* (3, 3, 21) */,
  32'h3d167d01 /* (31, 31, 17) */,
  32'h3d35f880 /* (27, 31, 17) */,
  32'h3d8f3655 /* (23, 31, 17) */,
  32'h3df92d6c /* (19, 31, 17) */,
  32'h3e09bd27 /* (15, 31, 17) */,
  32'h3dc031e4 /* (11, 31, 17) */,
  32'h3d5d3ed0 /* (7, 31, 17) */,
  32'h3d202be8 /* (3, 31, 17) */,
  32'h3d35f880 /* (31, 27, 17) */,
  32'h3d5e11d0 /* (27, 27, 17) */,
  32'h3db198fc /* (23, 27, 17) */,
  32'h3e1d0a10 /* (19, 27, 17) */,
  32'h3e2edbb4 /* (15, 27, 17) */,
  32'h3df05994 /* (11, 27, 17) */,
  32'h3d880917 /* (7, 27, 17) */,
  32'h3d424fe8 /* (3, 27, 17) */,
  32'h3d8f3655 /* (31, 23, 17) */,
  32'h3db198fc /* (27, 23, 17) */,
  32'h3e123783 /* (23, 23, 17) */,
  32'h3e8557f4 /* (19, 23, 17) */,
  32'h3e969108 /* (15, 23, 17) */,
  32'h3e49046a /* (11, 23, 17) */,
  32'h3ddc94c6 /* (7, 23, 17) */,
  32'h3d99caa3 /* (3, 23, 17) */,
  32'h3df92d6c /* (31, 19, 17) */,
  32'h3e1d0a10 /* (27, 19, 17) */,
  32'h3e8557f4 /* (23, 19, 17) */,
  32'h3efbd9fe /* (19, 19, 17) */,
  32'h3f1092e5 /* (15, 19, 17) */,
  32'h3eba8e90 /* (11, 19, 17) */,
  32'h3e45db44 /* (7, 19, 17) */,
  32'h3e068db8 /* (3, 19, 17) */,
  32'h3e09bd27 /* (31, 15, 17) */,
  32'h3e2edbb4 /* (27, 15, 17) */,
  32'h3e969108 /* (23, 15, 17) */,
  32'h3f1092e5 /* (19, 15, 17) */,
  32'h3f275a64 /* (15, 15, 17) */,
  32'h3ed4648a /* (11, 15, 17) */,
  32'h3e5db918 /* (7, 15, 17) */,
  32'h3e151f83 /* (3, 15, 17) */,
  32'h3dc031e4 /* (31, 11, 17) */,
  32'h3df05994 /* (27, 11, 17) */,
  32'h3e49046a /* (23, 11, 17) */,
  32'h3eba8e90 /* (19, 11, 17) */,
  32'h3ed4648a /* (15, 11, 17) */,
  32'h3e8b66c2 /* (11, 11, 17) */,
  32'h3e165b49 /* (7, 11, 17) */,
  32'h3dceffa6 /* (3, 11, 17) */,
  32'h3d5d3ed0 /* (31, 7, 17) */,
  32'h3d880917 /* (27, 7, 17) */,
  32'h3ddc94c6 /* (23, 7, 17) */,
  32'h3e45db44 /* (19, 7, 17) */,
  32'h3e5db918 /* (15, 7, 17) */,
  32'h3e165b49 /* (11, 7, 17) */,
  32'h3da7bf05 /* (7, 7, 17) */,
  32'h3d6ce397 /* (3, 7, 17) */,
  32'h3d202be8 /* (31, 3, 17) */,
  32'h3d424fe8 /* (27, 3, 17) */,
  32'h3d99caa3 /* (23, 3, 17) */,
  32'h3e068db8 /* (19, 3, 17) */,
  32'h3e151f83 /* (15, 3, 17) */,
  32'h3dceffa6 /* (11, 3, 17) */,
  32'h3d6ce397 /* (7, 3, 17) */,
  32'h3d2aacf2 /* (3, 3, 17) */,
  32'h3d1e42f1 /* (31, 31, 13) */,
  32'h3d398f3f /* (27, 31, 13) */,
  32'h3d8ac476 /* (23, 31, 13) */,
  32'h3de602d9 /* (19, 31, 13) */,
  32'h3df92d6c /* (15, 31, 13) */,
  32'h3db58f74 /* (11, 31, 13) */,
  32'h3d5c17b6 /* (7, 31, 13) */,
  32'h3d269671 /* (3, 31, 13) */,
  32'h3d398f3f /* (31, 27, 13) */,
  32'h3d5ce99d /* (27, 27, 13) */,
  32'h3da95898 /* (23, 27, 13) */,
  32'h3e0f99f2 /* (19, 27, 13) */,
  32'h3e1d0a10 /* (15, 27, 13) */,
  32'h3de04254 /* (11, 27, 13) */,
  32'h3d849ae2 /* (7, 27, 13) */,
  32'h3d4466f8 /* (3, 27, 13) */,
  32'h3d8ac476 /* (31, 23, 13) */,
  32'h3da95898 /* (27, 23, 13) */,
  32'h3e076ebd /* (23, 23, 13) */,
  32'h3e6f82ab /* (19, 23, 13) */,
  32'h3e8557f4 /* (15, 23, 13) */,
  32'h3e37494b /* (11, 23, 13) */,
  32'h3dcf79e9 /* (7, 23, 13) */,
  32'h3d942dc4 /* (3, 23, 13) */,
  32'h3de602d9 /* (31, 19, 13) */,
  32'h3e0f99f2 /* (27, 19, 13) */,
  32'h3e6f82ab /* (23, 19, 13) */,
  32'h3edd8ee5 /* (19, 19, 13) */,
  32'h3efbd9fe /* (15, 19, 13) */,
  32'h3ea5d30f /* (11, 19, 13) */,
  32'h3e336d1b /* (7, 19, 13) */,
  32'h3df79892 /* (3, 19, 13) */,
  32'h3df92d6c /* (31, 15, 13) */,
  32'h3e1d0a10 /* (27, 15, 13) */,
  32'h3e8557f4 /* (23, 15, 13) */,
  32'h3efbd9fe /* (19, 15, 13) */,
  32'h3f1092e5 /* (15, 15, 13) */,
  32'h3eba8e90 /* (11, 15, 13) */,
  32'h3e45db44 /* (7, 15, 13) */,
  32'h3e068db8 /* (3, 15, 13) */,
  32'h3db58f74 /* (31, 11, 13) */,
  32'h3de04254 /* (27, 11, 13) */,
  32'h3e37494b /* (23, 11, 13) */,
  32'h3ea5d30f /* (19, 11, 13) */,
  32'h3eba8e90 /* (15, 11, 13) */,
  32'h3e7af74d /* (11, 11, 13) */,
  32'h3e0aca9a /* (7, 11, 13) */,
  32'h3dc2b35d /* (3, 11, 13) */,
  32'h3d5c17b6 /* (31, 7, 13) */,
  32'h3d849ae2 /* (27, 7, 13) */,
  32'h3dcf79e9 /* (23, 7, 13) */,
  32'h3e336d1b /* (19, 7, 13) */,
  32'h3e45db44 /* (15, 7, 13) */,
  32'h3e0aca9a /* (11, 7, 13) */,
  32'h3da0c360 /* (7, 7, 13) */,
  32'h3d69f6ae /* (3, 7, 13) */,
  32'h3d269671 /* (31, 3, 13) */,
  32'h3d4466f8 /* (27, 3, 13) */,
  32'h3d942dc4 /* (23, 3, 13) */,
  32'h3df79892 /* (19, 3, 13) */,
  32'h3e068db8 /* (15, 3, 13) */,
  32'h3dc2b35d /* (11, 3, 13) */,
  32'h3d69f6ae /* (7, 3, 13) */,
  32'h3d2fb3ed /* (3, 3, 13) */,
  32'h3d11a602 /* (31, 31, 9) */,
  32'h3d170f20 /* (27, 31, 9) */,
  32'h3d3ee791 /* (23, 31, 9) */,
  32'h3d8ac476 /* (19, 31, 9) */,
  32'h3d8f3655 /* (15, 31, 9) */,
  32'h3d68852c /* (11, 31, 9) */,
  32'h3d245baa /* (7, 31, 9) */,
  32'h3d126006 /* (3, 31, 9) */,
  32'h3d170f20 /* (31, 27, 9) */,
  32'h3d24f869 /* (27, 27, 9) */,
  32'h3d5e7d3b /* (23, 27, 9) */,
  32'h3da95898 /* (19, 27, 9) */,
  32'h3db198fc /* (15, 27, 9) */,
  32'h3d8b02ad /* (11, 27, 9) */,
  32'h3d39ba58 /* (7, 27, 9) */,
  32'h3d1addce /* (3, 27, 9) */,
  32'h3d3ee791 /* (31, 23, 9) */,
  32'h3d5e7d3b /* (27, 23, 9) */,
  32'h3da4cfbf /* (23, 23, 9) */,
  32'h3e076ebd /* (19, 23, 9) */,
  32'h3e123783 /* (15, 23, 9) */,
  32'h3dd6aa1b /* (11, 23, 9) */,
  32'h3d8354ed /* (7, 23, 9) */,
  32'h3d48821f /* (3, 23, 9) */,
  32'h3d8ac476 /* (31, 19, 9) */,
  32'h3da95898 /* (27, 19, 9) */,
  32'h3e076ebd /* (23, 19, 9) */,
  32'h3e6f82ab /* (19, 19, 9) */,
  32'h3e8557f4 /* (15, 19, 9) */,
  32'h3e37494b /* (11, 19, 9) */,
  32'h3dcf79e9 /* (7, 19, 9) */,
  32'h3d942dc4 /* (3, 19, 9) */,
  32'h3d8f3655 /* (31, 15, 9) */,
  32'h3db198fc /* (27, 15, 9) */,
  32'h3e123783 /* (23, 15, 9) */,
  32'h3e8557f4 /* (19, 15, 9) */,
  32'h3e969108 /* (15, 15, 9) */,
  32'h3e49046a /* (11, 15, 9) */,
  32'h3ddc94c6 /* (7, 15, 9) */,
  32'h3d99caa3 /* (3, 15, 9) */,
  32'h3d68852c /* (31, 11, 9) */,
  32'h3d8b02ad /* (27, 11, 9) */,
  32'h3dd6aa1b /* (23, 11, 9) */,
  32'h3e37494b /* (19, 11, 9) */,
  32'h3e49046a /* (15, 11, 9) */,
  32'h3e0ea5fd /* (11, 11, 9) */,
  32'h3da777c1 /* (7, 11, 9) */,
  32'h3d767d5d /* (3, 11, 9) */,
  32'h3d245baa /* (31, 7, 9) */,
  32'h3d39ba58 /* (27, 7, 9) */,
  32'h3d8354ed /* (23, 7, 9) */,
  32'h3dcf79e9 /* (19, 7, 9) */,
  32'h3ddc94c6 /* (15, 7, 9) */,
  32'h3da777c1 /* (11, 7, 9) */,
  32'h3d563bcb /* (7, 7, 9) */,
  32'h3d2aad03 /* (3, 7, 9) */,
  32'h3d126006 /* (31, 3, 9) */,
  32'h3d1addce /* (27, 3, 9) */,
  32'h3d48821f /* (23, 3, 9) */,
  32'h3d942dc4 /* (19, 3, 9) */,
  32'h3d99caa3 /* (15, 3, 9) */,
  32'h3d767d5d /* (11, 3, 9) */,
  32'h3d2aad03 /* (7, 3, 9) */,
  32'h3d144047 /* (3, 3, 9) */,
  32'h3d6890ff /* (31, 31, 5) */,
  32'h3d249f29 /* (27, 31, 5) */,
  32'h3d170f20 /* (23, 31, 5) */,
  32'h3d398f3f /* (19, 31, 5) */,
  32'h3d35f880 /* (15, 31, 5) */,
  32'h3d26c9db /* (11, 31, 5) */,
  32'h3d151e01 /* (7, 31, 5) */,
  32'h3d45ae9a /* (3, 31, 5) */,
  32'h3d249f29 /* (31, 27, 5) */,
  32'h3d15ac37 /* (27, 27, 5) */,
  32'h3d24f869 /* (23, 27, 5) */,
  32'h3d5ce99d /* (19, 27, 5) */,
  32'h3d5e11d0 /* (15, 27, 5) */,
  32'h3d3fb488 /* (11, 27, 5) */,
  32'h3d170afd /* (7, 27, 5) */,
  32'h3d1ccb4c /* (3, 27, 5) */,
  32'h3d170f20 /* (31, 23, 5) */,
  32'h3d24f869 /* (27, 23, 5) */,
  32'h3d5e7d3b /* (23, 23, 5) */,
  32'h3da95898 /* (19, 23, 5) */,
  32'h3db198fc /* (15, 23, 5) */,
  32'h3d8b02ad /* (11, 23, 5) */,
  32'h3d39ba58 /* (7, 23, 5) */,
  32'h3d1addce /* (3, 23, 5) */,
  32'h3d398f3f /* (31, 19, 5) */,
  32'h3d5ce99d /* (27, 19, 5) */,
  32'h3da95898 /* (23, 19, 5) */,
  32'h3e0f99f2 /* (19, 19, 5) */,
  32'h3e1d0a10 /* (15, 19, 5) */,
  32'h3de04254 /* (11, 19, 5) */,
  32'h3d849ae2 /* (7, 19, 5) */,
  32'h3d4466f8 /* (3, 19, 5) */,
  32'h3d35f880 /* (31, 15, 5) */,
  32'h3d5e11d0 /* (27, 15, 5) */,
  32'h3db198fc /* (23, 15, 5) */,
  32'h3e1d0a10 /* (19, 15, 5) */,
  32'h3e2edbb4 /* (15, 15, 5) */,
  32'h3df05994 /* (11, 15, 5) */,
  32'h3d880917 /* (7, 15, 5) */,
  32'h3d424fe8 /* (3, 15, 5) */,
  32'h3d26c9db /* (31, 11, 5) */,
  32'h3d3fb488 /* (27, 11, 5) */,
  32'h3d8b02ad /* (23, 11, 5) */,
  32'h3de04254 /* (19, 11, 5) */,
  32'h3df05994 /* (15, 11, 5) */,
  32'h3db345e2 /* (11, 11, 5) */,
  32'h3d5ff008 /* (7, 11, 5) */,
  32'h3d2e4aa1 /* (3, 11, 5) */,
  32'h3d151e01 /* (31, 7, 5) */,
  32'h3d170afd /* (27, 7, 5) */,
  32'h3d39ba58 /* (23, 7, 5) */,
  32'h3d849ae2 /* (19, 7, 5) */,
  32'h3d880917 /* (15, 7, 5) */,
  32'h3d5ff008 /* (11, 7, 5) */,
  32'h3d21f168 /* (7, 7, 5) */,
  32'h3d147808 /* (3, 7, 5) */,
  32'h3d45ae9a /* (31, 3, 5) */,
  32'h3d1ccb4c /* (27, 3, 5) */,
  32'h3d1addce /* (23, 3, 5) */,
  32'h3d4466f8 /* (19, 3, 5) */,
  32'h3d424fe8 /* (15, 3, 5) */,
  32'h3d2e4aa1 /* (11, 3, 5) */,
  32'h3d147808 /* (7, 3, 5) */,
  32'h3d314afb /* (3, 3, 5) */,
  32'h3ec3aed4 /* (31, 31, 1) */,
  32'h3d6890ff /* (27, 31, 1) */,
  32'h3d11a602 /* (23, 31, 1) */,
  32'h3d1e42f1 /* (19, 31, 1) */,
  32'h3d167d01 /* (15, 31, 1) */,
  32'h3d151591 /* (11, 31, 1) */,
  32'h3d2402bf /* (7, 31, 1) */,
  32'h3deb372d /* (3, 31, 1) */,
  32'h3d6890ff /* (31, 27, 1) */,
  32'h3d249f29 /* (27, 27, 1) */,
  32'h3d170f20 /* (23, 27, 1) */,
  32'h3d398f3f /* (19, 27, 1) */,
  32'h3d35f880 /* (15, 27, 1) */,
  32'h3d26c9db /* (11, 27, 1) */,
  32'h3d151e01 /* (7, 27, 1) */,
  32'h3d45ae9a /* (3, 27, 1) */,
  32'h3d11a602 /* (31, 23, 1) */,
  32'h3d170f20 /* (27, 23, 1) */,
  32'h3d3ee791 /* (23, 23, 1) */,
  32'h3d8ac476 /* (19, 23, 1) */,
  32'h3d8f3655 /* (15, 23, 1) */,
  32'h3d68852c /* (11, 23, 1) */,
  32'h3d245baa /* (7, 23, 1) */,
  32'h3d126006 /* (3, 23, 1) */,
  32'h3d1e42f1 /* (31, 19, 1) */,
  32'h3d398f3f /* (27, 19, 1) */,
  32'h3d8ac476 /* (23, 19, 1) */,
  32'h3de602d9 /* (19, 19, 1) */,
  32'h3df92d6c /* (15, 19, 1) */,
  32'h3db58f74 /* (11, 19, 1) */,
  32'h3d5c17b6 /* (7, 19, 1) */,
  32'h3d269671 /* (3, 19, 1) */,
  32'h3d167d01 /* (31, 15, 1) */,
  32'h3d35f880 /* (27, 15, 1) */,
  32'h3d8f3655 /* (23, 15, 1) */,
  32'h3df92d6c /* (19, 15, 1) */,
  32'h3e09bd27 /* (15, 15, 1) */,
  32'h3dc031e4 /* (11, 15, 1) */,
  32'h3d5d3ed0 /* (7, 15, 1) */,
  32'h3d202be8 /* (3, 15, 1) */,
  32'h3d151591 /* (31, 11, 1) */,
  32'h3d26c9db /* (27, 11, 1) */,
  32'h3d68852c /* (23, 11, 1) */,
  32'h3db58f74 /* (19, 11, 1) */,
  32'h3dc031e4 /* (15, 11, 1) */,
  32'h3d9352ec /* (11, 11, 1) */,
  32'h3d3efe62 /* (7, 11, 1) */,
  32'h3d1a3ccf /* (3, 11, 1) */,
  32'h3d2402bf /* (31, 7, 1) */,
  32'h3d151e01 /* (27, 7, 1) */,
  32'h3d245baa /* (23, 7, 1) */,
  32'h3d5c17b6 /* (19, 7, 1) */,
  32'h3d5d3ed0 /* (15, 7, 1) */,
  32'h3d3efe62 /* (11, 7, 1) */,
  32'h3d167b79 /* (7, 7, 1) */,
  32'h3d1c3652 /* (3, 7, 1) */,
  32'h3deb372d /* (31, 3, 1) */,
  32'h3d45ae9a /* (27, 3, 1) */,
  32'h3d126006 /* (23, 3, 1) */,
  32'h3d269671 /* (19, 3, 1) */,
  32'h3d202be8 /* (15, 3, 1) */,
  32'h3d1a3ccf /* (11, 3, 1) */,
  32'h3d1c3652 /* (7, 3, 1) */,
  32'h3d960c3c /* (3, 3, 1) */,
  32'h3dbfa8df /* (30, 31, 29) */,
  32'h3d2ba889 /* (26, 31, 29) */,
  32'h3d14c0fd /* (22, 31, 29) */,
  32'h3d276174 /* (18, 31, 29) */,
  32'h3d276174 /* (14, 31, 29) */,
  32'h3d14c0fd /* (10, 31, 29) */,
  32'h3d2ba889 /* (6, 31, 29) */,
  32'h3dbfa8df /* (2, 31, 29) */,
  32'h3d3cd255 /* (30, 27, 29) */,
  32'h3d16d305 /* (26, 27, 29) */,
  32'h3d2344c4 /* (22, 27, 29) */,
  32'h3d487174 /* (18, 27, 29) */,
  32'h3d487174 /* (14, 27, 29) */,
  32'h3d2344c4 /* (10, 27, 29) */,
  32'h3d16d305 /* (6, 27, 29) */,
  32'h3d3cd255 /* (2, 27, 29) */,
  32'h3d12f42a /* (30, 23, 29) */,
  32'h3d215063 /* (26, 23, 29) */,
  32'h3d5dae2c /* (22, 23, 29) */,
  32'h3d9b2a7b /* (18, 23, 29) */,
  32'h3d9b2a7b /* (14, 23, 29) */,
  32'h3d5dae2c /* (10, 23, 29) */,
  32'h3d215063 /* (6, 23, 29) */,
  32'h3d12f42a /* (2, 23, 29) */,
  32'h3d29e985 /* (30, 19, 29) */,
  32'h3d54a03b /* (26, 19, 29) */,
  32'h3da99659 /* (22, 19, 29) */,
  32'h3e04d0b8 /* (18, 19, 29) */,
  32'h3e04d0b8 /* (14, 19, 29) */,
  32'h3da99659 /* (10, 19, 29) */,
  32'h3d54a03b /* (6, 19, 29) */,
  32'h3d29e985 /* (2, 19, 29) */,
  32'h3d240321 /* (30, 15, 29) */,
  32'h3d54ba37 /* (26, 15, 29) */,
  32'h3db22d06 /* (22, 15, 29) */,
  32'h3e11d12f /* (18, 15, 29) */,
  32'h3e11d12f /* (14, 15, 29) */,
  32'h3db22d06 /* (10, 15, 29) */,
  32'h3d54ba37 /* (6, 15, 29) */,
  32'h3d240321 /* (2, 15, 29) */,
  32'h3d1c5f03 /* (30, 11, 29) */,
  32'h3d39bb76 /* (26, 11, 29) */,
  32'h3d8ae43c /* (22, 11, 29) */,
  32'h3dce7d45 /* (18, 11, 29) */,
  32'h3dce7d45 /* (14, 11, 29) */,
  32'h3d8ae43c /* (10, 11, 29) */,
  32'h3d39bb76 /* (6, 11, 29) */,
  32'h3d1c5f03 /* (2, 11, 29) */,
  32'h3d1a2949 /* (30, 7, 29) */,
  32'h3d159d44 /* (26, 7, 29) */,
  32'h3d387393 /* (22, 7, 29) */,
  32'h3d71c736 /* (18, 7, 29) */,
  32'h3d71c736 /* (14, 7, 29) */,
  32'h3d387393 /* (10, 7, 29) */,
  32'h3d159d44 /* (6, 7, 29) */,
  32'h3d1a2949 /* (2, 7, 29) */,
  32'h3d866355 /* (30, 3, 29) */,
  32'h3d211f1b /* (26, 3, 29) */,
  32'h3d18cb02 /* (22, 3, 29) */,
  32'h3d3188e3 /* (18, 3, 29) */,
  32'h3d3188e3 /* (14, 3, 29) */,
  32'h3d18cb02 /* (10, 3, 29) */,
  32'h3d211f1b /* (6, 3, 29) */,
  32'h3d866355 /* (2, 3, 29) */,
  32'h3d20a35e /* (30, 31, 25) */,
  32'h3d146a43 /* (26, 31, 25) */,
  32'h3d305430 /* (22, 31, 25) */,
  32'h3d62906c /* (18, 31, 25) */,
  32'h3d62906c /* (14, 31, 25) */,
  32'h3d305430 /* (10, 31, 25) */,
  32'h3d146a43 /* (6, 31, 25) */,
  32'h3d20a35e /* (2, 31, 25) */,
  32'h3d14b1c0 /* (30, 27, 25) */,
  32'h3d1b2471 /* (26, 27, 25) */,
  32'h3d4b3dc7 /* (22, 27, 25) */,
  32'h3d8a0000 /* (18, 27, 25) */,
  32'h3d8a0000 /* (14, 27, 25) */,
  32'h3d4b3dc7 /* (10, 27, 25) */,
  32'h3d1b2471 /* (6, 27, 25) */,
  32'h3d14b1c0 /* (2, 27, 25) */,
  32'h3d26a1b5 /* (30, 23, 25) */,
  32'h3d45eb5b /* (26, 23, 25) */,
  32'h3d94014f /* (22, 23, 25) */,
  32'h3ddc09d8 /* (18, 23, 25) */,
  32'h3ddc09d8 /* (14, 23, 25) */,
  32'h3d94014f /* (10, 23, 25) */,
  32'h3d45eb5b /* (6, 23, 25) */,
  32'h3d26a1b5 /* (2, 23, 25) */,
  32'h3d6129ae /* (30, 19, 25) */,
  32'h3d90c8a7 /* (26, 19, 25) */,
  32'h3defa49b /* (22, 19, 25) */,
  32'h3e41f14c /* (18, 19, 25) */,
  32'h3e41f14c /* (14, 19, 25) */,
  32'h3defa49b /* (10, 19, 25) */,
  32'h3d90c8a7 /* (6, 19, 25) */,
  32'h3d6129ae /* (2, 19, 25) */,
  32'h3d62f778 /* (30, 15, 25) */,
  32'h3d95be73 /* (26, 15, 25) */,
  32'h3e009a19 /* (22, 15, 25) */,
  32'h3e57a44b /* (18, 15, 25) */,
  32'h3e57a44b /* (14, 15, 25) */,
  32'h3e009a19 /* (10, 15, 25) */,
  32'h3d95be73 /* (6, 15, 25) */,
  32'h3d62f778 /* (2, 15, 25) */,
  32'h3d42a7b8 /* (30, 11, 25) */,
  32'h3d71ecf9 /* (26, 11, 25) */,
  32'h3dbf3f1d /* (22, 11, 25) */,
  32'h3e14a5c9 /* (18, 11, 25) */,
  32'h3e14a5c9 /* (14, 11, 25) */,
  32'h3dbf3f1d /* (10, 11, 25) */,
  32'h3d71ecf9 /* (6, 11, 25) */,
  32'h3d42a7b8 /* (2, 11, 25) */,
  32'h3d1777c7 /* (30, 7, 25) */,
  32'h3d29a602 /* (26, 7, 25) */,
  32'h3d6deb12 /* (22, 7, 25) */,
  32'h3da8d240 /* (18, 7, 25) */,
  32'h3da8d240 /* (14, 7, 25) */,
  32'h3d6deb12 /* (10, 7, 25) */,
  32'h3d29a602 /* (6, 7, 25) */,
  32'h3d1777c7 /* (2, 7, 25) */,
  32'h3d1a2949 /* (30, 3, 25) */,
  32'h3d159d44 /* (26, 3, 25) */,
  32'h3d387393 /* (22, 3, 25) */,
  32'h3d71c736 /* (18, 3, 25) */,
  32'h3d71c736 /* (14, 3, 25) */,
  32'h3d387393 /* (10, 3, 25) */,
  32'h3d159d44 /* (6, 3, 25) */,
  32'h3d1a2949 /* (2, 3, 25) */,
  32'h3d16ed42 /* (30, 31, 21) */,
  32'h3d31191b /* (26, 31, 21) */,
  32'h3d829849 /* (22, 31, 21) */,
  32'h3dc01db4 /* (18, 31, 21) */,
  32'h3dc01db4 /* (14, 31, 21) */,
  32'h3d829849 /* (10, 31, 21) */,
  32'h3d31191b /* (6, 31, 21) */,
  32'h3d16ed42 /* (2, 31, 21) */,
  32'h3d29823f /* (30, 27, 21) */,
  32'h3d4d9045 /* (26, 27, 21) */,
  32'h3d9d9380 /* (22, 27, 21) */,
  32'h3deed79f /* (18, 27, 21) */,
  32'h3deed79f /* (14, 27, 21) */,
  32'h3d9d9380 /* (10, 27, 21) */,
  32'h3d4d9045 /* (6, 27, 21) */,
  32'h3d29823f /* (2, 27, 21) */,
  32'h3d6d9fa3 /* (30, 23, 21) */,
  32'h3d9750ce /* (26, 23, 21) */,
  32'h3df71c69 /* (22, 23, 21) */,
  32'h3e458f30 /* (18, 23, 21) */,
  32'h3e458f30 /* (14, 23, 21) */,
  32'h3df71c69 /* (10, 23, 21) */,
  32'h3d9750ce /* (6, 23, 21) */,
  32'h3d6d9fa3 /* (2, 23, 21) */,
  32'h3dba5db4 /* (30, 19, 21) */,
  32'h3df74dbc /* (26, 19, 21) */,
  32'h3e562fb1 /* (22, 19, 21) */,
  32'h3eb517ce /* (18, 19, 21) */,
  32'h3eb517ce /* (14, 19, 21) */,
  32'h3e562fb1 /* (10, 19, 21) */,
  32'h3df74dbc /* (6, 19, 21) */,
  32'h3dba5db4 /* (2, 19, 21) */,
  32'h3dc59b81 /* (30, 15, 21) */,
  32'h3e0533d0 /* (26, 15, 21) */,
  32'h3e6c6ac0 /* (22, 15, 21) */,
  32'h3eccf8ff /* (18, 15, 21) */,
  32'h3eccf8ff /* (14, 15, 21) */,
  32'h3e6c6ac0 /* (10, 15, 21) */,
  32'h3e0533d0 /* (6, 15, 21) */,
  32'h3dc59b81 /* (2, 15, 21) */,
  32'h3d96eb50 /* (30, 11, 21) */,
  32'h3dc480ba /* (26, 11, 21) */,
  32'h3e257fc6 /* (22, 11, 21) */,
  32'h3e882756 /* (18, 11, 21) */,
  32'h3e882756 /* (14, 11, 21) */,
  32'h3e257fc6 /* (10, 11, 21) */,
  32'h3dc480ba /* (6, 11, 21) */,
  32'h3d96eb50 /* (2, 11, 21) */,
  32'h3d42a7b8 /* (30, 7, 21) */,
  32'h3d71ecf9 /* (26, 7, 21) */,
  32'h3dbf3f1d /* (22, 7, 21) */,
  32'h3e14a5c9 /* (18, 7, 21) */,
  32'h3e14a5c9 /* (14, 7, 21) */,
  32'h3dbf3f1d /* (10, 7, 21) */,
  32'h3d71ecf9 /* (6, 7, 21) */,
  32'h3d42a7b8 /* (2, 7, 21) */,
  32'h3d1c5f03 /* (30, 3, 21) */,
  32'h3d39bb76 /* (26, 3, 21) */,
  32'h3d8ae43c /* (22, 3, 21) */,
  32'h3dce7d45 /* (18, 3, 21) */,
  32'h3dce7d45 /* (14, 3, 21) */,
  32'h3d8ae43c /* (10, 3, 21) */,
  32'h3d39bb76 /* (6, 3, 21) */,
  32'h3d1c5f03 /* (2, 3, 21) */,
  32'h3d1a0745 /* (30, 31, 17) */,
  32'h3d46f53f /* (26, 31, 17) */,
  32'h3da5ac70 /* (22, 31, 17) */,
  32'h3e06d8bb /* (18, 31, 17) */,
  32'h3e06d8bb /* (14, 31, 17) */,
  32'h3da5ac70 /* (10, 31, 17) */,
  32'h3d46f53f /* (6, 31, 17) */,
  32'h3d1a0745 /* (2, 31, 17) */,
  32'h3d3a7be5 /* (30, 27, 17) */,
  32'h3d73b16f /* (26, 27, 17) */,
  32'h3dce52e6 /* (22, 27, 17) */,
  32'h3e2a981c /* (18, 27, 17) */,
  32'h3e2a981c /* (14, 27, 17) */,
  32'h3dce52e6 /* (10, 27, 17) */,
  32'h3d73b16f /* (6, 27, 17) */,
  32'h3d3a7be5 /* (2, 27, 17) */,
  32'h3d9314c2 /* (30, 23, 17) */,
  32'h3dc42ad0 /* (26, 23, 17) */,
  32'h3e2b3653 /* (22, 23, 17) */,
  32'h3e91e4f8 /* (18, 23, 17) */,
  32'h3e91e4f8 /* (14, 23, 17) */,
  32'h3e2b3653 /* (10, 23, 17) */,
  32'h3dc42ad0 /* (6, 23, 17) */,
  32'h3d9314c2 /* (2, 23, 17) */,
  32'h3e003b1e /* (30, 19, 17) */,
  32'h3e2ea39a /* (26, 19, 17) */,
  32'h3e9d80fb /* (22, 19, 17) */,
  32'h3f0af24f /* (18, 19, 17) */,
  32'h3f0af24f /* (14, 19, 17) */,
  32'h3e9d80fb /* (10, 19, 17) */,
  32'h3e2ea39a /* (6, 19, 17) */,
  32'h3e003b1e /* (2, 19, 17) */,
  32'h3e0de5f8 /* (30, 15, 17) */,
  32'h3e430b11 /* (26, 15, 17) */,
  32'h3eb2925b /* (22, 15, 17) */,
  32'h3f202f9a /* (18, 15, 17) */,
  32'h3f202f9a /* (14, 15, 17) */,
  32'h3eb2925b /* (10, 15, 17) */,
  32'h3e430b11 /* (6, 15, 17) */,
  32'h3e0de5f8 /* (2, 15, 17) */,
  32'h3dc59b81 /* (30, 11, 17) */,
  32'h3e0533d0 /* (26, 11, 17) */,
  32'h3e6c6ac0 /* (22, 11, 17) */,
  32'h3eccf8ff /* (18, 11, 17) */,
  32'h3eccf8ff /* (14, 11, 17) */,
  32'h3e6c6ac0 /* (10, 11, 17) */,
  32'h3e0533d0 /* (6, 11, 17) */,
  32'h3dc59b81 /* (2, 11, 17) */,
  32'h3d62f778 /* (30, 7, 17) */,
  32'h3d95be73 /* (26, 7, 17) */,
  32'h3e009a19 /* (22, 7, 17) */,
  32'h3e57a44b /* (18, 7, 17) */,
  32'h3e57a44b /* (14, 7, 17) */,
  32'h3e009a19 /* (10, 7, 17) */,
  32'h3d95be73 /* (6, 7, 17) */,
  32'h3d62f778 /* (2, 7, 17) */,
  32'h3d240321 /* (30, 3, 17) */,
  32'h3d54ba37 /* (26, 3, 17) */,
  32'h3db22d06 /* (22, 3, 17) */,
  32'h3e11d12f /* (18, 3, 17) */,
  32'h3e11d12f /* (14, 3, 17) */,
  32'h3db22d06 /* (10, 3, 17) */,
  32'h3d54ba37 /* (6, 3, 17) */,
  32'h3d240321 /* (2, 3, 17) */,
  32'h3d214ba3 /* (30, 31, 13) */,
  32'h3d4876ff /* (26, 31, 13) */,
  32'h3d9e7894 /* (22, 31, 13) */,
  32'h3df65860 /* (18, 31, 13) */,
  32'h3df65860 /* (14, 31, 13) */,
  32'h3d9e7894 /* (10, 31, 13) */,
  32'h3d4876ff /* (6, 31, 13) */,
  32'h3d214ba3 /* (2, 31, 13) */,
  32'h3d3d84de /* (30, 27, 13) */,
  32'h3d700ffa /* (26, 27, 13) */,
  32'h3dc29629 /* (22, 27, 13) */,
  32'h3e1a8d8c /* (18, 27, 13) */,
  32'h3e1a8d8c /* (14, 27, 13) */,
  32'h3dc29629 /* (10, 27, 13) */,
  32'h3d700ffa /* (6, 27, 13) */,
  32'h3d3d84de /* (2, 27, 13) */,
  32'h3d8e358b /* (30, 23, 13) */,
  32'h3db9d5f4 /* (26, 23, 13) */,
  32'h3e1d56b2 /* (22, 23, 13) */,
  32'h3e821787 /* (18, 23, 13) */,
  32'h3e821787 /* (14, 23, 13) */,
  32'h3e1d56b2 /* (10, 23, 13) */,
  32'h3db9d5f4 /* (6, 23, 13) */,
  32'h3d8e358b /* (2, 23, 13) */,
  32'h3dec70da /* (30, 19, 13) */,
  32'h3e1f113d /* (26, 19, 13) */,
  32'h3e8cbae1 /* (22, 19, 13) */,
  32'h3ef33ce4 /* (18, 19, 13) */,
  32'h3ef33ce4 /* (14, 19, 13) */,
  32'h3e8cbae1 /* (10, 19, 13) */,
  32'h3e1f113d /* (6, 19, 13) */,
  32'h3dec70da /* (2, 19, 13) */,
  32'h3e003b1e /* (30, 15, 13) */,
  32'h3e2ea39a /* (26, 15, 13) */,
  32'h3e9d80fb /* (22, 15, 13) */,
  32'h3f0af24f /* (18, 15, 13) */,
  32'h3f0af24f /* (14, 15, 13) */,
  32'h3e9d80fb /* (10, 15, 13) */,
  32'h3e2ea39a /* (6, 15, 13) */,
  32'h3e003b1e /* (2, 15, 13) */,
  32'h3dba5db4 /* (30, 11, 13) */,
  32'h3df74dbc /* (26, 11, 13) */,
  32'h3e562fb1 /* (22, 11, 13) */,
  32'h3eb517ce /* (18, 11, 13) */,
  32'h3eb517ce /* (14, 11, 13) */,
  32'h3e562fb1 /* (10, 11, 13) */,
  32'h3df74dbc /* (6, 11, 13) */,
  32'h3dba5db4 /* (2, 11, 13) */,
  32'h3d6129ae /* (30, 7, 13) */,
  32'h3d90c8a7 /* (26, 7, 13) */,
  32'h3defa49b /* (22, 7, 13) */,
  32'h3e41f14c /* (18, 7, 13) */,
  32'h3e41f14c /* (14, 7, 13) */,
  32'h3defa49b /* (10, 7, 13) */,
  32'h3d90c8a7 /* (6, 7, 13) */,
  32'h3d6129ae /* (2, 7, 13) */,
  32'h3d29e985 /* (30, 3, 13) */,
  32'h3d54a03b /* (26, 3, 13) */,
  32'h3da99659 /* (22, 3, 13) */,
  32'h3e04d0b8 /* (18, 3, 13) */,
  32'h3e04d0b8 /* (14, 3, 13) */,
  32'h3da99659 /* (10, 3, 13) */,
  32'h3d54a03b /* (6, 3, 13) */,
  32'h3d29e985 /* (2, 3, 13) */,
  32'h3d11c69f /* (30, 31, 9) */,
  32'h3d1c53e8 /* (26, 31, 9) */,
  32'h3d52081f /* (22, 31, 9) */,
  32'h3d90dff9 /* (18, 31, 9) */,
  32'h3d90dff9 /* (14, 31, 9) */,
  32'h3d52081f /* (10, 31, 9) */,
  32'h3d1c53e8 /* (6, 31, 9) */,
  32'h3d11c69f /* (2, 31, 9) */,
  32'h3d18622e /* (30, 27, 9) */,
  32'h3d2db0cc /* (26, 27, 9) */,
  32'h3d781ae6 /* (22, 27, 9) */,
  32'h3db24f8e /* (18, 27, 9) */,
  32'h3db24f8e /* (14, 27, 9) */,
  32'h3d781ae6 /* (10, 27, 9) */,
  32'h3d2db0cc /* (6, 27, 9) */,
  32'h3d18622e /* (2, 27, 9) */,
  32'h3d42665b /* (30, 23, 9) */,
  32'h3d6fd024 /* (26, 23, 9) */,
  32'h3dbbc730 /* (22, 23, 9) */,
  32'h3e10cac5 /* (18, 23, 9) */,
  32'h3e10cac5 /* (14, 23, 9) */,
  32'h3dbbc730 /* (10, 23, 9) */,
  32'h3d6fd024 /* (6, 23, 9) */,
  32'h3d42665b /* (2, 23, 9) */,
  32'h3d8e358b /* (30, 19, 9) */,
  32'h3db9d5f4 /* (26, 19, 9) */,
  32'h3e1d56b2 /* (22, 19, 9) */,
  32'h3e821787 /* (18, 19, 9) */,
  32'h3e821787 /* (14, 19, 9) */,
  32'h3e1d56b2 /* (10, 19, 9) */,
  32'h3db9d5f4 /* (6, 19, 9) */,
  32'h3d8e358b /* (2, 19, 9) */,
  32'h3d9314c2 /* (30, 15, 9) */,
  32'h3dc42ad0 /* (26, 15, 9) */,
  32'h3e2b3653 /* (22, 15, 9) */,
  32'h3e91e4f8 /* (18, 15, 9) */,
  32'h3e91e4f8 /* (14, 15, 9) */,
  32'h3e2b3653 /* (10, 15, 9) */,
  32'h3dc42ad0 /* (6, 15, 9) */,
  32'h3d9314c2 /* (2, 15, 9) */,
  32'h3d6d9fa3 /* (30, 11, 9) */,
  32'h3d9750ce /* (26, 11, 9) */,
  32'h3df71c69 /* (22, 11, 9) */,
  32'h3e458f30 /* (18, 11, 9) */,
  32'h3e458f30 /* (14, 11, 9) */,
  32'h3df71c69 /* (10, 11, 9) */,
  32'h3d9750ce /* (6, 11, 9) */,
  32'h3d6d9fa3 /* (2, 11, 9) */,
  32'h3d26a1b5 /* (30, 7, 9) */,
  32'h3d45eb5b /* (26, 7, 9) */,
  32'h3d94014f /* (22, 7, 9) */,
  32'h3ddc09d8 /* (18, 7, 9) */,
  32'h3ddc09d8 /* (14, 7, 9) */,
  32'h3d94014f /* (10, 7, 9) */,
  32'h3d45eb5b /* (6, 7, 9) */,
  32'h3d26a1b5 /* (2, 7, 9) */,
  32'h3d12f42a /* (30, 3, 9) */,
  32'h3d215063 /* (26, 3, 9) */,
  32'h3d5dae2c /* (22, 3, 9) */,
  32'h3d9b2a7b /* (18, 3, 9) */,
  32'h3d9b2a7b /* (14, 3, 9) */,
  32'h3d5dae2c /* (10, 3, 9) */,
  32'h3d215063 /* (6, 3, 9) */,
  32'h3d12f42a /* (2, 3, 9) */,
  32'h3d59109a /* (30, 31, 5) */,
  32'h3d1a8b5a /* (26, 31, 5) */,
  32'h3d1d9589 /* (22, 31, 5) */,
  32'h3d3c7841 /* (18, 31, 5) */,
  32'h3d3c7841 /* (14, 31, 5) */,
  32'h3d1d9589 /* (10, 31, 5) */,
  32'h3d1a8b5a /* (6, 31, 5) */,
  32'h3d59109a /* (2, 31, 5) */,
  32'h3d213c91 /* (30, 27, 5) */,
  32'h3d14f7ce /* (26, 27, 5) */,
  32'h3d30fc5a /* (22, 27, 5) */,
  32'h3d63687e /* (18, 27, 5) */,
  32'h3d63687e /* (14, 27, 5) */,
  32'h3d30fc5a /* (10, 27, 5) */,
  32'h3d14f7ce /* (6, 27, 5) */,
  32'h3d213c91 /* (2, 27, 5) */,
  32'h3d18622e /* (30, 23, 5) */,
  32'h3d2db0cc /* (26, 23, 5) */,
  32'h3d781ae6 /* (22, 23, 5) */,
  32'h3db24f8e /* (18, 23, 5) */,
  32'h3db24f8e /* (14, 23, 5) */,
  32'h3d781ae6 /* (10, 23, 5) */,
  32'h3d2db0cc /* (6, 23, 5) */,
  32'h3d18622e /* (2, 23, 5) */,
  32'h3d3d84de /* (30, 19, 5) */,
  32'h3d700ffa /* (26, 19, 5) */,
  32'h3dc29629 /* (22, 19, 5) */,
  32'h3e1a8d8c /* (18, 19, 5) */,
  32'h3e1a8d8c /* (14, 19, 5) */,
  32'h3dc29629 /* (10, 19, 5) */,
  32'h3d700ffa /* (6, 19, 5) */,
  32'h3d3d84de /* (2, 19, 5) */,
  32'h3d3a7be5 /* (30, 15, 5) */,
  32'h3d73b16f /* (26, 15, 5) */,
  32'h3dce52e6 /* (22, 15, 5) */,
  32'h3e2a981c /* (18, 15, 5) */,
  32'h3e2a981c /* (14, 15, 5) */,
  32'h3dce52e6 /* (10, 15, 5) */,
  32'h3d73b16f /* (6, 15, 5) */,
  32'h3d3a7be5 /* (2, 15, 5) */,
  32'h3d29823f /* (30, 11, 5) */,
  32'h3d4d9045 /* (26, 11, 5) */,
  32'h3d9d9380 /* (22, 11, 5) */,
  32'h3deed79f /* (18, 11, 5) */,
  32'h3deed79f /* (14, 11, 5) */,
  32'h3d9d9380 /* (10, 11, 5) */,
  32'h3d4d9045 /* (6, 11, 5) */,
  32'h3d29823f /* (2, 11, 5) */,
  32'h3d14b1c0 /* (30, 7, 5) */,
  32'h3d1b2471 /* (26, 7, 5) */,
  32'h3d4b3dc7 /* (22, 7, 5) */,
  32'h3d8a0000 /* (18, 7, 5) */,
  32'h3d8a0000 /* (14, 7, 5) */,
  32'h3d4b3dc7 /* (10, 7, 5) */,
  32'h3d1b2471 /* (6, 7, 5) */,
  32'h3d14b1c0 /* (2, 7, 5) */,
  32'h3d3cd255 /* (30, 3, 5) */,
  32'h3d16d305 /* (26, 3, 5) */,
  32'h3d2344c4 /* (22, 3, 5) */,
  32'h3d487174 /* (18, 3, 5) */,
  32'h3d487174 /* (14, 3, 5) */,
  32'h3d2344c4 /* (10, 3, 5) */,
  32'h3d16d305 /* (6, 3, 5) */,
  32'h3d3cd255 /* (2, 3, 5) */,
  32'h3e4aeee2 /* (30, 31, 1) */,
  32'h3d3c9698 /* (26, 31, 1) */,
  32'h3d119771 /* (22, 31, 1) */,
  32'h3d1e0bb6 /* (18, 31, 1) */,
  32'h3d1e0bb6 /* (14, 31, 1) */,
  32'h3d119771 /* (10, 31, 1) */,
  32'h3d3c9698 /* (6, 31, 1) */,
  32'h3e4aeee2 /* (2, 31, 1) */,
  32'h3d59109a /* (30, 27, 1) */,
  32'h3d1a8b5a /* (26, 27, 1) */,
  32'h3d1d9589 /* (22, 27, 1) */,
  32'h3d3c7841 /* (18, 27, 1) */,
  32'h3d3c7841 /* (14, 27, 1) */,
  32'h3d1d9589 /* (10, 27, 1) */,
  32'h3d1a8b5a /* (6, 27, 1) */,
  32'h3d59109a /* (2, 27, 1) */,
  32'h3d11c69f /* (30, 23, 1) */,
  32'h3d1c53e8 /* (26, 23, 1) */,
  32'h3d52081f /* (22, 23, 1) */,
  32'h3d90dff9 /* (18, 23, 1) */,
  32'h3d90dff9 /* (14, 23, 1) */,
  32'h3d52081f /* (10, 23, 1) */,
  32'h3d1c53e8 /* (6, 23, 1) */,
  32'h3d11c69f /* (2, 23, 1) */,
  32'h3d214ba3 /* (30, 19, 1) */,
  32'h3d4876ff /* (26, 19, 1) */,
  32'h3d9e7894 /* (22, 19, 1) */,
  32'h3df65860 /* (18, 19, 1) */,
  32'h3df65860 /* (14, 19, 1) */,
  32'h3d9e7894 /* (10, 19, 1) */,
  32'h3d4876ff /* (6, 19, 1) */,
  32'h3d214ba3 /* (2, 19, 1) */,
  32'h3d1a0745 /* (30, 15, 1) */,
  32'h3d46f53f /* (26, 15, 1) */,
  32'h3da5ac70 /* (22, 15, 1) */,
  32'h3e06d8bb /* (18, 15, 1) */,
  32'h3e06d8bb /* (14, 15, 1) */,
  32'h3da5ac70 /* (10, 15, 1) */,
  32'h3d46f53f /* (6, 15, 1) */,
  32'h3d1a0745 /* (2, 15, 1) */,
  32'h3d16ed42 /* (30, 11, 1) */,
  32'h3d31191b /* (26, 11, 1) */,
  32'h3d829849 /* (22, 11, 1) */,
  32'h3dc01db4 /* (18, 11, 1) */,
  32'h3dc01db4 /* (14, 11, 1) */,
  32'h3d829849 /* (10, 11, 1) */,
  32'h3d31191b /* (6, 11, 1) */,
  32'h3d16ed42 /* (2, 11, 1) */,
  32'h3d20a35e /* (30, 7, 1) */,
  32'h3d146a43 /* (26, 7, 1) */,
  32'h3d305430 /* (22, 7, 1) */,
  32'h3d62906c /* (18, 7, 1) */,
  32'h3d62906c /* (14, 7, 1) */,
  32'h3d305430 /* (10, 7, 1) */,
  32'h3d146a43 /* (6, 7, 1) */,
  32'h3d20a35e /* (2, 7, 1) */,
  32'h3dbfa8df /* (30, 3, 1) */,
  32'h3d2ba889 /* (26, 3, 1) */,
  32'h3d14c0fd /* (22, 3, 1) */,
  32'h3d276174 /* (18, 3, 1) */,
  32'h3d276174 /* (14, 3, 1) */,
  32'h3d14c0fd /* (10, 3, 1) */,
  32'h3d2ba889 /* (6, 3, 1) */,
  32'h3dbfa8df /* (2, 3, 1) */,
  32'h3d960c3c /* (29, 31, 29) */,
  32'h3d1c3652 /* (25, 31, 29) */,
  32'h3d1a3ccf /* (21, 31, 29) */,
  32'h3d202be8 /* (17, 31, 29) */,
  32'h3d269671 /* (13, 31, 29) */,
  32'h3d126006 /* (9, 31, 29) */,
  32'h3d45ae9a /* (5, 31, 29) */,
  32'h3deb372d /* (1, 31, 29) */,
  32'h3d314afb /* (29, 27, 29) */,
  32'h3d147808 /* (25, 27, 29) */,
  32'h3d2e4aa1 /* (21, 27, 29) */,
  32'h3d424fe8 /* (17, 27, 29) */,
  32'h3d4466f8 /* (13, 27, 29) */,
  32'h3d1addce /* (9, 27, 29) */,
  32'h3d1ccb4c /* (5, 27, 29) */,
  32'h3d45ae9a /* (1, 27, 29) */,
  32'h3d144047 /* (29, 23, 29) */,
  32'h3d2aad03 /* (25, 23, 29) */,
  32'h3d767d5d /* (21, 23, 29) */,
  32'h3d99caa3 /* (17, 23, 29) */,
  32'h3d942dc4 /* (13, 23, 29) */,
  32'h3d48821f /* (9, 23, 29) */,
  32'h3d1addce /* (5, 23, 29) */,
  32'h3d126006 /* (1, 23, 29) */,
  32'h3d2fb3ed /* (29, 19, 29) */,
  32'h3d69f6ae /* (25, 19, 29) */,
  32'h3dc2b35d /* (21, 19, 29) */,
  32'h3e068db8 /* (17, 19, 29) */,
  32'h3df79892 /* (13, 19, 29) */,
  32'h3d942dc4 /* (9, 19, 29) */,
  32'h3d4466f8 /* (5, 19, 29) */,
  32'h3d269671 /* (1, 19, 29) */,
  32'h3d2aacf2 /* (29, 15, 29) */,
  32'h3d6ce397 /* (25, 15, 29) */,
  32'h3dceffa6 /* (21, 15, 29) */,
  32'h3e151f83 /* (17, 15, 29) */,
  32'h3e068db8 /* (13, 15, 29) */,
  32'h3d99caa3 /* (9, 15, 29) */,
  32'h3d424fe8 /* (5, 15, 29) */,
  32'h3d202be8 /* (1, 15, 29) */,
  32'h3d202a91 /* (29, 11, 29) */,
  32'h3d490aba /* (25, 11, 29) */,
  32'h3d9d27e1 /* (21, 11, 29) */,
  32'h3dceffa6 /* (17, 11, 29) */,
  32'h3dc2b35d /* (13, 11, 29) */,
  32'h3d767d5d /* (9, 11, 29) */,
  32'h3d2e4aa1 /* (5, 11, 29) */,
  32'h3d1a3ccf /* (1, 11, 29) */,
  32'h3d179239 /* (29, 7, 29) */,
  32'h3d1969a9 /* (25, 7, 29) */,
  32'h3d490aba /* (21, 7, 29) */,
  32'h3d6ce397 /* (17, 7, 29) */,
  32'h3d69f6ae /* (13, 7, 29) */,
  32'h3d2aad03 /* (9, 7, 29) */,
  32'h3d147808 /* (5, 7, 29) */,
  32'h3d1c3652 /* (1, 7, 29) */,
  32'h3d68b01f /* (29, 3, 29) */,
  32'h3d179239 /* (25, 3, 29) */,
  32'h3d202a91 /* (21, 3, 29) */,
  32'h3d2aacf2 /* (17, 3, 29) */,
  32'h3d2fb3ed /* (13, 3, 29) */,
  32'h3d144047 /* (9, 3, 29) */,
  32'h3d314afb /* (5, 3, 29) */,
  32'h3d960c3c /* (1, 3, 29) */,
  32'h3d1c3652 /* (29, 31, 25) */,
  32'h3d167b79 /* (25, 31, 25) */,
  32'h3d3efe62 /* (21, 31, 25) */,
  32'h3d5d3ed0 /* (17, 31, 25) */,
  32'h3d5c17b6 /* (13, 31, 25) */,
  32'h3d245baa /* (9, 31, 25) */,
  32'h3d151e01 /* (5, 31, 25) */,
  32'h3d2402bf /* (1, 31, 25) */,
  32'h3d147808 /* (29, 27, 25) */,
  32'h3d21f168 /* (25, 27, 25) */,
  32'h3d5ff008 /* (21, 27, 25) */,
  32'h3d880917 /* (17, 27, 25) */,
  32'h3d849ae2 /* (13, 27, 25) */,
  32'h3d39ba58 /* (9, 27, 25) */,
  32'h3d170afd /* (5, 27, 25) */,
  32'h3d151e01 /* (1, 27, 25) */,
  32'h3d2aad03 /* (29, 23, 25) */,
  32'h3d563bcb /* (25, 23, 25) */,
  32'h3da777c1 /* (21, 23, 25) */,
  32'h3ddc94c6 /* (17, 23, 25) */,
  32'h3dcf79e9 /* (13, 23, 25) */,
  32'h3d8354ed /* (9, 23, 25) */,
  32'h3d39ba58 /* (5, 23, 25) */,
  32'h3d245baa /* (1, 23, 25) */,
  32'h3d69f6ae /* (29, 19, 25) */,
  32'h3da0c360 /* (25, 19, 25) */,
  32'h3e0aca9a /* (21, 19, 25) */,
  32'h3e45db44 /* (17, 19, 25) */,
  32'h3e336d1b /* (13, 19, 25) */,
  32'h3dcf79e9 /* (9, 19, 25) */,
  32'h3d849ae2 /* (5, 19, 25) */,
  32'h3d5c17b6 /* (1, 19, 25) */,
  32'h3d6ce397 /* (29, 15, 25) */,
  32'h3da7bf05 /* (25, 15, 25) */,
  32'h3e165b49 /* (21, 15, 25) */,
  32'h3e5db918 /* (17, 15, 25) */,
  32'h3e45db44 /* (13, 15, 25) */,
  32'h3ddc94c6 /* (9, 15, 25) */,
  32'h3d880917 /* (5, 15, 25) */,
  32'h3d5d3ed0 /* (1, 15, 25) */,
  32'h3d490aba /* (29, 11, 25) */,
  32'h3d84ce75 /* (25, 11, 25) */,
  32'h3ddb1c7f /* (21, 11, 25) */,
  32'h3e165b49 /* (17, 11, 25) */,
  32'h3e0aca9a /* (13, 11, 25) */,
  32'h3da777c1 /* (9, 11, 25) */,
  32'h3d5ff008 /* (5, 11, 25) */,
  32'h3d3efe62 /* (1, 11, 25) */,
  32'h3d1969a9 /* (29, 7, 25) */,
  32'h3d348078 /* (25, 7, 25) */,
  32'h3d84ce75 /* (21, 7, 25) */,
  32'h3da7bf05 /* (17, 7, 25) */,
  32'h3da0c360 /* (13, 7, 25) */,
  32'h3d563bcb /* (9, 7, 25) */,
  32'h3d21f168 /* (5, 7, 25) */,
  32'h3d167b79 /* (1, 7, 25) */,
  32'h3d179239 /* (29, 3, 25) */,
  32'h3d1969a9 /* (25, 3, 25) */,
  32'h3d490aba /* (21, 3, 25) */,
  32'h3d6ce397 /* (17, 3, 25) */,
  32'h3d69f6ae /* (13, 3, 25) */,
  32'h3d2aad03 /* (9, 3, 25) */,
  32'h3d147808 /* (5, 3, 25) */,
  32'h3d1c3652 /* (1, 3, 25) */,
  32'h3d1a3ccf /* (29, 31, 21) */,
  32'h3d3efe62 /* (25, 31, 21) */,
  32'h3d9352ec /* (21, 31, 21) */,
  32'h3dc031e4 /* (17, 31, 21) */,
  32'h3db58f74 /* (13, 31, 21) */,
  32'h3d68852c /* (9, 31, 21) */,
  32'h3d26c9db /* (5, 31, 21) */,
  32'h3d151591 /* (1, 31, 21) */,
  32'h3d2e4aa1 /* (29, 27, 21) */,
  32'h3d5ff008 /* (25, 27, 21) */,
  32'h3db345e2 /* (21, 27, 21) */,
  32'h3df05994 /* (17, 27, 21) */,
  32'h3de04254 /* (13, 27, 21) */,
  32'h3d8b02ad /* (9, 27, 21) */,
  32'h3d3fb488 /* (5, 27, 21) */,
  32'h3d26c9db /* (1, 27, 21) */,
  32'h3d767d5d /* (29, 23, 21) */,
  32'h3da777c1 /* (25, 23, 21) */,
  32'h3e0ea5fd /* (21, 23, 21) */,
  32'h3e49046a /* (17, 23, 21) */,
  32'h3e37494b /* (13, 23, 21) */,
  32'h3dd6aa1b /* (9, 23, 21) */,
  32'h3d8b02ad /* (5, 23, 21) */,
  32'h3d68852c /* (1, 23, 21) */,
  32'h3dc2b35d /* (29, 19, 21) */,
  32'h3e0aca9a /* (25, 19, 21) */,
  32'h3e7af74d /* (21, 19, 21) */,
  32'h3eba8e90 /* (17, 19, 21) */,
  32'h3ea5d30f /* (13, 19, 21) */,
  32'h3e37494b /* (9, 19, 21) */,
  32'h3de04254 /* (5, 19, 21) */,
  32'h3db58f74 /* (1, 19, 21) */,
  32'h3dceffa6 /* (29, 15, 21) */,
  32'h3e165b49 /* (25, 15, 21) */,
  32'h3e8b66c2 /* (21, 15, 21) */,
  32'h3ed4648a /* (17, 15, 21) */,
  32'h3eba8e90 /* (13, 15, 21) */,
  32'h3e49046a /* (9, 15, 21) */,
  32'h3df05994 /* (5, 15, 21) */,
  32'h3dc031e4 /* (1, 15, 21) */,
  32'h3d9d27e1 /* (29, 11, 21) */,
  32'h3ddb1c7f /* (25, 11, 21) */,
  32'h3e4089a2 /* (21, 11, 21) */,
  32'h3e8b66c2 /* (17, 11, 21) */,
  32'h3e7af74d /* (13, 11, 21) */,
  32'h3e0ea5fd /* (9, 11, 21) */,
  32'h3db345e2 /* (5, 11, 21) */,
  32'h3d9352ec /* (1, 11, 21) */,
  32'h3d490aba /* (29, 7, 21) */,
  32'h3d84ce75 /* (25, 7, 21) */,
  32'h3ddb1c7f /* (21, 7, 21) */,
  32'h3e165b49 /* (17, 7, 21) */,
  32'h3e0aca9a /* (13, 7, 21) */,
  32'h3da777c1 /* (9, 7, 21) */,
  32'h3d5ff008 /* (5, 7, 21) */,
  32'h3d3efe62 /* (1, 7, 21) */,
  32'h3d202a91 /* (29, 3, 21) */,
  32'h3d490aba /* (25, 3, 21) */,
  32'h3d9d27e1 /* (21, 3, 21) */,
  32'h3dceffa6 /* (17, 3, 21) */,
  32'h3dc2b35d /* (13, 3, 21) */,
  32'h3d767d5d /* (9, 3, 21) */,
  32'h3d2e4aa1 /* (5, 3, 21) */,
  32'h3d1a3ccf /* (1, 3, 21) */,
  32'h3d202be8 /* (29, 31, 17) */,
  32'h3d5d3ed0 /* (25, 31, 17) */,
  32'h3dc031e4 /* (21, 31, 17) */,
  32'h3e09bd27 /* (17, 31, 17) */,
  32'h3df92d6c /* (13, 31, 17) */,
  32'h3d8f3655 /* (9, 31, 17) */,
  32'h3d35f880 /* (5, 31, 17) */,
  32'h3d167d01 /* (1, 31, 17) */,
  32'h3d424fe8 /* (29, 27, 17) */,
  32'h3d880917 /* (25, 27, 17) */,
  32'h3df05994 /* (21, 27, 17) */,
  32'h3e2edbb4 /* (17, 27, 17) */,
  32'h3e1d0a10 /* (13, 27, 17) */,
  32'h3db198fc /* (9, 27, 17) */,
  32'h3d5e11d0 /* (5, 27, 17) */,
  32'h3d35f880 /* (1, 27, 17) */,
  32'h3d99caa3 /* (29, 23, 17) */,
  32'h3ddc94c6 /* (25, 23, 17) */,
  32'h3e49046a /* (21, 23, 17) */,
  32'h3e969108 /* (17, 23, 17) */,
  32'h3e8557f4 /* (13, 23, 17) */,
  32'h3e123783 /* (9, 23, 17) */,
  32'h3db198fc /* (5, 23, 17) */,
  32'h3d8f3655 /* (1, 23, 17) */,
  32'h3e068db8 /* (29, 19, 17) */,
  32'h3e45db44 /* (25, 19, 17) */,
  32'h3eba8e90 /* (21, 19, 17) */,
  32'h3f1092e5 /* (17, 19, 17) */,
  32'h3efbd9fe /* (13, 19, 17) */,
  32'h3e8557f4 /* (9, 19, 17) */,
  32'h3e1d0a10 /* (5, 19, 17) */,
  32'h3df92d6c /* (1, 19, 17) */,
  32'h3e151f83 /* (29, 15, 17) */,
  32'h3e5db918 /* (25, 15, 17) */,
  32'h3ed4648a /* (21, 15, 17) */,
  32'h3f275a64 /* (17, 15, 17) */,
  32'h3f1092e5 /* (13, 15, 17) */,
  32'h3e969108 /* (9, 15, 17) */,
  32'h3e2edbb4 /* (5, 15, 17) */,
  32'h3e09bd27 /* (1, 15, 17) */,
  32'h3dceffa6 /* (29, 11, 17) */,
  32'h3e165b49 /* (25, 11, 17) */,
  32'h3e8b66c2 /* (21, 11, 17) */,
  32'h3ed4648a /* (17, 11, 17) */,
  32'h3eba8e90 /* (13, 11, 17) */,
  32'h3e49046a /* (9, 11, 17) */,
  32'h3df05994 /* (5, 11, 17) */,
  32'h3dc031e4 /* (1, 11, 17) */,
  32'h3d6ce397 /* (29, 7, 17) */,
  32'h3da7bf05 /* (25, 7, 17) */,
  32'h3e165b49 /* (21, 7, 17) */,
  32'h3e5db918 /* (17, 7, 17) */,
  32'h3e45db44 /* (13, 7, 17) */,
  32'h3ddc94c6 /* (9, 7, 17) */,
  32'h3d880917 /* (5, 7, 17) */,
  32'h3d5d3ed0 /* (1, 7, 17) */,
  32'h3d2aacf2 /* (29, 3, 17) */,
  32'h3d6ce397 /* (25, 3, 17) */,
  32'h3dceffa6 /* (21, 3, 17) */,
  32'h3e151f83 /* (17, 3, 17) */,
  32'h3e068db8 /* (13, 3, 17) */,
  32'h3d99caa3 /* (9, 3, 17) */,
  32'h3d424fe8 /* (5, 3, 17) */,
  32'h3d202be8 /* (1, 3, 17) */,
  32'h3d269671 /* (29, 31, 13) */,
  32'h3d5c17b6 /* (25, 31, 13) */,
  32'h3db58f74 /* (21, 31, 13) */,
  32'h3df92d6c /* (17, 31, 13) */,
  32'h3de602d9 /* (13, 31, 13) */,
  32'h3d8ac476 /* (9, 31, 13) */,
  32'h3d398f3f /* (5, 31, 13) */,
  32'h3d1e42f1 /* (1, 31, 13) */,
  32'h3d4466f8 /* (29, 27, 13) */,
  32'h3d849ae2 /* (25, 27, 13) */,
  32'h3de04254 /* (21, 27, 13) */,
  32'h3e1d0a10 /* (17, 27, 13) */,
  32'h3e0f99f2 /* (13, 27, 13) */,
  32'h3da95898 /* (9, 27, 13) */,
  32'h3d5ce99d /* (5, 27, 13) */,
  32'h3d398f3f /* (1, 27, 13) */,
  32'h3d942dc4 /* (29, 23, 13) */,
  32'h3dcf79e9 /* (25, 23, 13) */,
  32'h3e37494b /* (21, 23, 13) */,
  32'h3e8557f4 /* (17, 23, 13) */,
  32'h3e6f82ab /* (13, 23, 13) */,
  32'h3e076ebd /* (9, 23, 13) */,
  32'h3da95898 /* (5, 23, 13) */,
  32'h3d8ac476 /* (1, 23, 13) */,
  32'h3df79892 /* (29, 19, 13) */,
  32'h3e336d1b /* (25, 19, 13) */,
  32'h3ea5d30f /* (21, 19, 13) */,
  32'h3efbd9fe /* (17, 19, 13) */,
  32'h3edd8ee5 /* (13, 19, 13) */,
  32'h3e6f82ab /* (9, 19, 13) */,
  32'h3e0f99f2 /* (5, 19, 13) */,
  32'h3de602d9 /* (1, 19, 13) */,
  32'h3e068db8 /* (29, 15, 13) */,
  32'h3e45db44 /* (25, 15, 13) */,
  32'h3eba8e90 /* (21, 15, 13) */,
  32'h3f1092e5 /* (17, 15, 13) */,
  32'h3efbd9fe /* (13, 15, 13) */,
  32'h3e8557f4 /* (9, 15, 13) */,
  32'h3e1d0a10 /* (5, 15, 13) */,
  32'h3df92d6c /* (1, 15, 13) */,
  32'h3dc2b35d /* (29, 11, 13) */,
  32'h3e0aca9a /* (25, 11, 13) */,
  32'h3e7af74d /* (21, 11, 13) */,
  32'h3eba8e90 /* (17, 11, 13) */,
  32'h3ea5d30f /* (13, 11, 13) */,
  32'h3e37494b /* (9, 11, 13) */,
  32'h3de04254 /* (5, 11, 13) */,
  32'h3db58f74 /* (1, 11, 13) */,
  32'h3d69f6ae /* (29, 7, 13) */,
  32'h3da0c360 /* (25, 7, 13) */,
  32'h3e0aca9a /* (21, 7, 13) */,
  32'h3e45db44 /* (17, 7, 13) */,
  32'h3e336d1b /* (13, 7, 13) */,
  32'h3dcf79e9 /* (9, 7, 13) */,
  32'h3d849ae2 /* (5, 7, 13) */,
  32'h3d5c17b6 /* (1, 7, 13) */,
  32'h3d2fb3ed /* (29, 3, 13) */,
  32'h3d69f6ae /* (25, 3, 13) */,
  32'h3dc2b35d /* (21, 3, 13) */,
  32'h3e068db8 /* (17, 3, 13) */,
  32'h3df79892 /* (13, 3, 13) */,
  32'h3d942dc4 /* (9, 3, 13) */,
  32'h3d4466f8 /* (5, 3, 13) */,
  32'h3d269671 /* (1, 3, 13) */,
  32'h3d126006 /* (29, 31, 9) */,
  32'h3d245baa /* (25, 31, 9) */,
  32'h3d68852c /* (21, 31, 9) */,
  32'h3d8f3655 /* (17, 31, 9) */,
  32'h3d8ac476 /* (13, 31, 9) */,
  32'h3d3ee791 /* (9, 31, 9) */,
  32'h3d170f20 /* (5, 31, 9) */,
  32'h3d11a602 /* (1, 31, 9) */,
  32'h3d1addce /* (29, 27, 9) */,
  32'h3d39ba58 /* (25, 27, 9) */,
  32'h3d8b02ad /* (21, 27, 9) */,
  32'h3db198fc /* (17, 27, 9) */,
  32'h3da95898 /* (13, 27, 9) */,
  32'h3d5e7d3b /* (9, 27, 9) */,
  32'h3d24f869 /* (5, 27, 9) */,
  32'h3d170f20 /* (1, 27, 9) */,
  32'h3d48821f /* (29, 23, 9) */,
  32'h3d8354ed /* (25, 23, 9) */,
  32'h3dd6aa1b /* (21, 23, 9) */,
  32'h3e123783 /* (17, 23, 9) */,
  32'h3e076ebd /* (13, 23, 9) */,
  32'h3da4cfbf /* (9, 23, 9) */,
  32'h3d5e7d3b /* (5, 23, 9) */,
  32'h3d3ee791 /* (1, 23, 9) */,
  32'h3d942dc4 /* (29, 19, 9) */,
  32'h3dcf79e9 /* (25, 19, 9) */,
  32'h3e37494b /* (21, 19, 9) */,
  32'h3e8557f4 /* (17, 19, 9) */,
  32'h3e6f82ab /* (13, 19, 9) */,
  32'h3e076ebd /* (9, 19, 9) */,
  32'h3da95898 /* (5, 19, 9) */,
  32'h3d8ac476 /* (1, 19, 9) */,
  32'h3d99caa3 /* (29, 15, 9) */,
  32'h3ddc94c6 /* (25, 15, 9) */,
  32'h3e49046a /* (21, 15, 9) */,
  32'h3e969108 /* (17, 15, 9) */,
  32'h3e8557f4 /* (13, 15, 9) */,
  32'h3e123783 /* (9, 15, 9) */,
  32'h3db198fc /* (5, 15, 9) */,
  32'h3d8f3655 /* (1, 15, 9) */,
  32'h3d767d5d /* (29, 11, 9) */,
  32'h3da777c1 /* (25, 11, 9) */,
  32'h3e0ea5fd /* (21, 11, 9) */,
  32'h3e49046a /* (17, 11, 9) */,
  32'h3e37494b /* (13, 11, 9) */,
  32'h3dd6aa1b /* (9, 11, 9) */,
  32'h3d8b02ad /* (5, 11, 9) */,
  32'h3d68852c /* (1, 11, 9) */,
  32'h3d2aad03 /* (29, 7, 9) */,
  32'h3d563bcb /* (25, 7, 9) */,
  32'h3da777c1 /* (21, 7, 9) */,
  32'h3ddc94c6 /* (17, 7, 9) */,
  32'h3dcf79e9 /* (13, 7, 9) */,
  32'h3d8354ed /* (9, 7, 9) */,
  32'h3d39ba58 /* (5, 7, 9) */,
  32'h3d245baa /* (1, 7, 9) */,
  32'h3d144047 /* (29, 3, 9) */,
  32'h3d2aad03 /* (25, 3, 9) */,
  32'h3d767d5d /* (21, 3, 9) */,
  32'h3d99caa3 /* (17, 3, 9) */,
  32'h3d942dc4 /* (13, 3, 9) */,
  32'h3d48821f /* (9, 3, 9) */,
  32'h3d1addce /* (5, 3, 9) */,
  32'h3d126006 /* (1, 3, 9) */,
  32'h3d45ae9a /* (29, 31, 5) */,
  32'h3d151e01 /* (25, 31, 5) */,
  32'h3d26c9db /* (21, 31, 5) */,
  32'h3d35f880 /* (17, 31, 5) */,
  32'h3d398f3f /* (13, 31, 5) */,
  32'h3d170f20 /* (9, 31, 5) */,
  32'h3d249f29 /* (5, 31, 5) */,
  32'h3d6890ff /* (1, 31, 5) */,
  32'h3d1ccb4c /* (29, 27, 5) */,
  32'h3d170afd /* (25, 27, 5) */,
  32'h3d3fb488 /* (21, 27, 5) */,
  32'h3d5e11d0 /* (17, 27, 5) */,
  32'h3d5ce99d /* (13, 27, 5) */,
  32'h3d24f869 /* (9, 27, 5) */,
  32'h3d15ac37 /* (5, 27, 5) */,
  32'h3d249f29 /* (1, 27, 5) */,
  32'h3d1addce /* (29, 23, 5) */,
  32'h3d39ba58 /* (25, 23, 5) */,
  32'h3d8b02ad /* (21, 23, 5) */,
  32'h3db198fc /* (17, 23, 5) */,
  32'h3da95898 /* (13, 23, 5) */,
  32'h3d5e7d3b /* (9, 23, 5) */,
  32'h3d24f869 /* (5, 23, 5) */,
  32'h3d170f20 /* (1, 23, 5) */,
  32'h3d4466f8 /* (29, 19, 5) */,
  32'h3d849ae2 /* (25, 19, 5) */,
  32'h3de04254 /* (21, 19, 5) */,
  32'h3e1d0a10 /* (17, 19, 5) */,
  32'h3e0f99f2 /* (13, 19, 5) */,
  32'h3da95898 /* (9, 19, 5) */,
  32'h3d5ce99d /* (5, 19, 5) */,
  32'h3d398f3f /* (1, 19, 5) */,
  32'h3d424fe8 /* (29, 15, 5) */,
  32'h3d880917 /* (25, 15, 5) */,
  32'h3df05994 /* (21, 15, 5) */,
  32'h3e2edbb4 /* (17, 15, 5) */,
  32'h3e1d0a10 /* (13, 15, 5) */,
  32'h3db198fc /* (9, 15, 5) */,
  32'h3d5e11d0 /* (5, 15, 5) */,
  32'h3d35f880 /* (1, 15, 5) */,
  32'h3d2e4aa1 /* (29, 11, 5) */,
  32'h3d5ff008 /* (25, 11, 5) */,
  32'h3db345e2 /* (21, 11, 5) */,
  32'h3df05994 /* (17, 11, 5) */,
  32'h3de04254 /* (13, 11, 5) */,
  32'h3d8b02ad /* (9, 11, 5) */,
  32'h3d3fb488 /* (5, 11, 5) */,
  32'h3d26c9db /* (1, 11, 5) */,
  32'h3d147808 /* (29, 7, 5) */,
  32'h3d21f168 /* (25, 7, 5) */,
  32'h3d5ff008 /* (21, 7, 5) */,
  32'h3d880917 /* (17, 7, 5) */,
  32'h3d849ae2 /* (13, 7, 5) */,
  32'h3d39ba58 /* (9, 7, 5) */,
  32'h3d170afd /* (5, 7, 5) */,
  32'h3d151e01 /* (1, 7, 5) */,
  32'h3d314afb /* (29, 3, 5) */,
  32'h3d147808 /* (25, 3, 5) */,
  32'h3d2e4aa1 /* (21, 3, 5) */,
  32'h3d424fe8 /* (17, 3, 5) */,
  32'h3d4466f8 /* (13, 3, 5) */,
  32'h3d1addce /* (9, 3, 5) */,
  32'h3d1ccb4c /* (5, 3, 5) */,
  32'h3d45ae9a /* (1, 3, 5) */,
  32'h3deb372d /* (29, 31, 1) */,
  32'h3d2402bf /* (25, 31, 1) */,
  32'h3d151591 /* (21, 31, 1) */,
  32'h3d167d01 /* (17, 31, 1) */,
  32'h3d1e42f1 /* (13, 31, 1) */,
  32'h3d11a602 /* (9, 31, 1) */,
  32'h3d6890ff /* (5, 31, 1) */,
  32'h3ec3aed4 /* (1, 31, 1) */,
  32'h3d45ae9a /* (29, 27, 1) */,
  32'h3d151e01 /* (25, 27, 1) */,
  32'h3d26c9db /* (21, 27, 1) */,
  32'h3d35f880 /* (17, 27, 1) */,
  32'h3d398f3f /* (13, 27, 1) */,
  32'h3d170f20 /* (9, 27, 1) */,
  32'h3d249f29 /* (5, 27, 1) */,
  32'h3d6890ff /* (1, 27, 1) */,
  32'h3d126006 /* (29, 23, 1) */,
  32'h3d245baa /* (25, 23, 1) */,
  32'h3d68852c /* (21, 23, 1) */,
  32'h3d8f3655 /* (17, 23, 1) */,
  32'h3d8ac476 /* (13, 23, 1) */,
  32'h3d3ee791 /* (9, 23, 1) */,
  32'h3d170f20 /* (5, 23, 1) */,
  32'h3d11a602 /* (1, 23, 1) */,
  32'h3d269671 /* (29, 19, 1) */,
  32'h3d5c17b6 /* (25, 19, 1) */,
  32'h3db58f74 /* (21, 19, 1) */,
  32'h3df92d6c /* (17, 19, 1) */,
  32'h3de602d9 /* (13, 19, 1) */,
  32'h3d8ac476 /* (9, 19, 1) */,
  32'h3d398f3f /* (5, 19, 1) */,
  32'h3d1e42f1 /* (1, 19, 1) */,
  32'h3d202be8 /* (29, 15, 1) */,
  32'h3d5d3ed0 /* (25, 15, 1) */,
  32'h3dc031e4 /* (21, 15, 1) */,
  32'h3e09bd27 /* (17, 15, 1) */,
  32'h3df92d6c /* (13, 15, 1) */,
  32'h3d8f3655 /* (9, 15, 1) */,
  32'h3d35f880 /* (5, 15, 1) */,
  32'h3d167d01 /* (1, 15, 1) */,
  32'h3d1a3ccf /* (29, 11, 1) */,
  32'h3d3efe62 /* (25, 11, 1) */,
  32'h3d9352ec /* (21, 11, 1) */,
  32'h3dc031e4 /* (17, 11, 1) */,
  32'h3db58f74 /* (13, 11, 1) */,
  32'h3d68852c /* (9, 11, 1) */,
  32'h3d26c9db /* (5, 11, 1) */,
  32'h3d151591 /* (1, 11, 1) */,
  32'h3d1c3652 /* (29, 7, 1) */,
  32'h3d167b79 /* (25, 7, 1) */,
  32'h3d3efe62 /* (21, 7, 1) */,
  32'h3d5d3ed0 /* (17, 7, 1) */,
  32'h3d5c17b6 /* (13, 7, 1) */,
  32'h3d245baa /* (9, 7, 1) */,
  32'h3d151e01 /* (5, 7, 1) */,
  32'h3d2402bf /* (1, 7, 1) */,
  32'h3d960c3c /* (29, 3, 1) */,
  32'h3d1c3652 /* (25, 3, 1) */,
  32'h3d1a3ccf /* (21, 3, 1) */,
  32'h3d202be8 /* (17, 3, 1) */,
  32'h3d269671 /* (13, 3, 1) */,
  32'h3d126006 /* (9, 3, 1) */,
  32'h3d45ae9a /* (5, 3, 1) */,
  32'h3deb372d /* (1, 3, 1) */,
  32'h3d6eb36b /* (28, 31, 29) */,
  32'h3d146963 /* (24, 31, 29) */,
  32'h3d210eee /* (20, 31, 29) */,
  32'h3d0fbc59 /* (16, 31, 29) */,
  32'h3d210eee /* (12, 31, 29) */,
  32'h3d146963 /* (8, 31, 29) */,
  32'h3d6eb36b /* (4, 31, 29) */,
  32'h3dff9e3f /* (0, 31, 29) */,
  32'h3d25f5ce /* (28, 27, 29) */,
  32'h3d15d660 /* (24, 27, 29) */,
  32'h3d3a4ebb /* (20, 27, 29) */,
  32'h3d3046d8 /* (16, 27, 29) */,
  32'h3d3a4ebb /* (12, 27, 29) */,
  32'h3d15d660 /* (8, 27, 29) */,
  32'h3d25f5ce /* (4, 27, 29) */,
  32'h3d490b0e /* (0, 27, 29) */,
  32'h3d16b5b2 /* (28, 23, 29) */,
  32'h3d37919e /* (24, 23, 29) */,
  32'h3d886b82 /* (20, 23, 29) */,
  32'h3d8e3848 /* (16, 23, 29) */,
  32'h3d886b82 /* (12, 23, 29) */,
  32'h3d37919e /* (8, 23, 29) */,
  32'h3d16b5b2 /* (4, 23, 29) */,
  32'h3d1237a7 /* (0, 23, 29) */,
  32'h3d385879 /* (28, 19, 29) */,
  32'h3d82c188 /* (24, 19, 29) */,
  32'h3dddef48 /* (20, 19, 29) */,
  32'h3dfdd31f /* (16, 19, 29) */,
  32'h3dddef48 /* (12, 19, 29) */,
  32'h3d82c188 /* (8, 19, 29) */,
  32'h3d385879 /* (4, 19, 29) */,
  32'h3d258110 /* (0, 19, 29) */,
  32'h3d349293 /* (28, 15, 29) */,
  32'h3d8608f0 /* (24, 15, 29) */,
  32'h3deea44d /* (20, 15, 29) */,
  32'h3e0de417 /* (16, 15, 29) */,
  32'h3deea44d /* (12, 15, 29) */,
  32'h3d8608f0 /* (8, 15, 29) */,
  32'h3d349293 /* (4, 15, 29) */,
  32'h3d1eeabe /* (0, 15, 29) */,
  32'h3d25fa09 /* (28, 11, 29) */,
  32'h3d5d0a38 /* (24, 11, 29) */,
  32'h3db0b965 /* (20, 11, 29) */,
  32'h3dc1602b /* (16, 11, 29) */,
  32'h3db0b965 /* (12, 11, 29) */,
  32'h3d5d0a38 /* (8, 11, 29) */,
  32'h3d25fa09 /* (4, 11, 29) */,
  32'h3d198ce9 /* (0, 11, 29) */,
  32'h3d155fa4 /* (28, 7, 29) */,
  32'h3d2054cd /* (24, 7, 29) */,
  32'h3d5ab0e1 /* (20, 7, 29) */,
  32'h3d58de26 /* (16, 7, 29) */,
  32'h3d5ab0e1 /* (12, 7, 29) */,
  32'h3d2054cd /* (8, 7, 29) */,
  32'h3d155fa4 /* (4, 7, 29) */,
  32'h3d1cfd70 /* (0, 7, 29) */,
  32'h3d4920d0 /* (28, 3, 29) */,
  32'h3d1392fe /* (24, 3, 29) */,
  32'h3d28b308 /* (20, 3, 29) */,
  32'h3d19c07a /* (16, 3, 29) */,
  32'h3d28b308 /* (12, 3, 29) */,
  32'h3d1392fe /* (8, 3, 29) */,
  32'h3d4920d0 /* (4, 3, 29) */,
  32'h3d9c797c /* (0, 3, 29) */,
  32'h3d17ff6b /* (28, 31, 25) */,
  32'h3d1bb8b6 /* (24, 31, 25) */,
  32'h3d4ea8e5 /* (20, 31, 25) */,
  32'h3d49f75a /* (16, 31, 25) */,
  32'h3d4ea8e5 /* (12, 31, 25) */,
  32'h3d1bb8b6 /* (8, 31, 25) */,
  32'h3d17ff6b /* (4, 31, 25) */,
  32'h3d25463b /* (0, 31, 25) */,
  32'h3d1508af /* (28, 27, 25) */,
  32'h3d2bff3e /* (24, 27, 25) */,
  32'h3d75e4d4 /* (20, 27, 25) */,
  32'h3d7a662c /* (16, 27, 25) */,
  32'h3d75e4d4 /* (12, 27, 25) */,
  32'h3d2bff3e /* (8, 27, 25) */,
  32'h3d1508af /* (4, 27, 25) */,
  32'h3d154f7b /* (0, 27, 25) */,
  32'h3d30de15 /* (28, 23, 25) */,
  32'h3d6b8b35 /* (24, 23, 25) */,
  32'h3dbc51f9 /* (20, 23, 25) */,
  32'h3dce1075 /* (16, 23, 25) */,
  32'h3dbc51f9 /* (12, 23, 25) */,
  32'h3d6b8b35 /* (8, 23, 25) */,
  32'h3d30de15 /* (4, 23, 25) */,
  32'h3d23a039 /* (0, 23, 25) */,
  32'h3d770afc /* (28, 19, 25) */,
  32'h3db56072 /* (24, 19, 25) */,
  32'h3e1f8cbf /* (20, 19, 25) */,
  32'h3e3bd4ee /* (16, 19, 25) */,
  32'h3e1f8cbf /* (12, 19, 25) */,
  32'h3db56072 /* (8, 19, 25) */,
  32'h3d770afc /* (4, 19, 25) */,
  32'h3d5a6fdd /* (0, 19, 25) */,
  32'h3d7b9f11 /* (28, 15, 25) */,
  32'h3dbf0444 /* (24, 15, 25) */,
  32'h3e2e6a71 /* (20, 15, 25) */,
  32'h3e540b9b /* (16, 15, 25) */,
  32'h3e2e6a71 /* (12, 15, 25) */,
  32'h3dbf0444 /* (8, 15, 25) */,
  32'h3d7b9f11 /* (4, 15, 25) */,
  32'h3d5b6048 /* (0, 15, 25) */,
  32'h3d52976b /* (28, 11, 25) */,
  32'h3d941bce /* (24, 11, 25) */,
  32'h3df94537 /* (20, 11, 25) */,
  32'h3e0d9cf0 /* (16, 11, 25) */,
  32'h3df94537 /* (12, 11, 25) */,
  32'h3d941bce /* (8, 11, 25) */,
  32'h3d52976b /* (4, 11, 25) */,
  32'h3d3dcd22 /* (0, 11, 25) */,
  32'h3d1cbb18 /* (28, 7, 25) */,
  32'h3d432bf1 /* (24, 7, 25) */,
  32'h3d938890 /* (20, 7, 25) */,
  32'h3d9b7830 /* (16, 7, 25) */,
  32'h3d938890 /* (12, 7, 25) */,
  32'h3d432bf1 /* (8, 7, 25) */,
  32'h3d1cbb18 /* (4, 7, 25) */,
  32'h3d162f74 /* (0, 7, 25) */,
  32'h3d155fa4 /* (28, 3, 25) */,
  32'h3d2054cd /* (24, 3, 25) */,
  32'h3d5ab0e1 /* (20, 3, 25) */,
  32'h3d58de26 /* (16, 3, 25) */,
  32'h3d5ab0e1 /* (12, 3, 25) */,
  32'h3d2054cd /* (8, 3, 25) */,
  32'h3d155fa4 /* (4, 3, 25) */,
  32'h3d1cfd70 /* (0, 3, 25) */,
  32'h3d1f5dc3 /* (28, 31, 21) */,
  32'h3d513c3d /* (24, 31, 21) */,
  32'h3da53628 /* (20, 31, 21) */,
  32'h3db336e0 /* (16, 31, 21) */,
  32'h3da53628 /* (12, 31, 21) */,
  32'h3d513c3d /* (8, 31, 21) */,
  32'h3d1f5dc3 /* (4, 31, 21) */,
  32'h3d147e90 /* (0, 31, 21) */,
  32'h3d358341 /* (28, 27, 21) */,
  32'h3d77c8fd /* (24, 27, 21) */,
  32'h3dca9d53 /* (20, 27, 21) */,
  32'h3de14ffa /* (16, 27, 21) */,
  32'h3dca9d53 /* (12, 27, 21) */,
  32'h3d77c8fd /* (8, 27, 21) */,
  32'h3d358341 /* (4, 27, 21) */,
  32'h3d25e815 /* (0, 27, 21) */,
  32'h3d81d711 /* (28, 23, 21) */,
  32'h3dbc4d73 /* (24, 23, 21) */,
  32'h3e23781b /* (20, 23, 21) */,
  32'h3e3e5da7 /* (16, 23, 21) */,
  32'h3e23781b /* (12, 23, 21) */,
  32'h3dbc4d73 /* (8, 23, 21) */,
  32'h3d81d711 /* (4, 23, 21) */,
  32'h3d66dac1 /* (0, 23, 21) */,
  32'h3dcf13a3 /* (28, 19, 21) */,
  32'h3e1e607d /* (24, 19, 21) */,
  32'h3e91dfe2 /* (20, 19, 21) */,
  32'h3eb2bd2a /* (16, 19, 21) */,
  32'h3e91dfe2 /* (12, 19, 21) */,
  32'h3e1e607d /* (8, 19, 21) */,
  32'h3dcf13a3 /* (4, 19, 21) */,
  32'h3db3fd83 /* (0, 19, 21) */,
  32'h3ddcf428 /* (28, 15, 21) */,
  32'h3e2c9c6c /* (24, 15, 21) */,
  32'h3ea31756 /* (20, 15, 21) */,
  32'h3ecca1ac /* (16, 15, 21) */,
  32'h3ea31756 /* (12, 15, 21) */,
  32'h3e2c9c6c /* (8, 15, 21) */,
  32'h3ddcf428 /* (4, 15, 21) */,
  32'h3dbe6d47 /* (0, 15, 21) */,
  32'h3da66ad4 /* (28, 11, 21) */,
  32'h3df84bb3 /* (24, 11, 21) */,
  32'h3e5e44ac /* (20, 11, 21) */,
  32'h3e84c8e0 /* (16, 11, 21) */,
  32'h3e5e44ac /* (12, 11, 21) */,
  32'h3df84bb3 /* (8, 11, 21) */,
  32'h3da66ad4 /* (4, 11, 21) */,
  32'h3d922642 /* (0, 11, 21) */,
  32'h3d52976b /* (28, 7, 21) */,
  32'h3d941bce /* (24, 7, 21) */,
  32'h3df94537 /* (20, 7, 21) */,
  32'h3e0d9cf0 /* (16, 7, 21) */,
  32'h3df94537 /* (12, 7, 21) */,
  32'h3d941bce /* (8, 7, 21) */,
  32'h3d52976b /* (4, 7, 21) */,
  32'h3d3dcd22 /* (0, 7, 21) */,
  32'h3d25fa09 /* (28, 3, 21) */,
  32'h3d5d0a38 /* (24, 3, 21) */,
  32'h3db0b965 /* (20, 3, 21) */,
  32'h3dc1602b /* (16, 3, 21) */,
  32'h3db0b965 /* (12, 3, 21) */,
  32'h3d5d0a38 /* (8, 3, 21) */,
  32'h3d25fa09 /* (4, 3, 21) */,
  32'h3d198ce9 /* (0, 3, 21) */,
  32'h3d294c4b /* (28, 31, 17) */,
  32'h3d7a003f /* (24, 31, 17) */,
  32'h3ddd43c2 /* (20, 31, 17) */,
  32'h3e02e976 /* (16, 31, 17) */,
  32'h3ddd43c2 /* (12, 31, 17) */,
  32'h3d7a003f /* (8, 31, 17) */,
  32'h3d294c4b /* (4, 31, 17) */,
  32'h3d155505 /* (0, 31, 17) */,
  32'h3d4def9b /* (28, 27, 17) */,
  32'h3d9a5b6b /* (24, 27, 17) */,
  32'h3e0ae903 /* (20, 27, 17) */,
  32'h3e26bbbb /* (16, 27, 17) */,
  32'h3e0ae903 /* (12, 27, 17) */,
  32'h3d9a5b6b /* (8, 27, 17) */,
  32'h3d4def9b /* (4, 27, 17) */,
  32'h3d347f0a /* (0, 27, 17) */,
  32'h3da3c1ed /* (28, 23, 17) */,
  32'h3dfc30a3 /* (24, 23, 17) */,
  32'h3e6a25fd /* (20, 23, 17) */,
  32'h3e908107 /* (16, 23, 17) */,
  32'h3e6a25fd /* (12, 23, 17) */,
  32'h3dfc30a3 /* (8, 23, 17) */,
  32'h3da3c1ed /* (4, 23, 17) */,
  32'h3d8df2c1 /* (0, 23, 17) */,
  32'h3e0ff4ce /* (28, 19, 17) */,
  32'h3e640ba2 /* (24, 19, 17) */,
  32'h3edb3822 /* (20, 19, 17) */,
  32'h3f0bd969 /* (16, 19, 17) */,
  32'h3edb3822 /* (12, 19, 17) */,
  32'h3e640ba2 /* (8, 19, 17) */,
  32'h3e0ff4ce /* (4, 19, 17) */,
  32'h3df6cc6d /* (0, 19, 17) */,
  32'h3e1fe07e /* (28, 15, 17) */,
  32'h3e803f85 /* (24, 15, 17) */,
  32'h3efaa119 /* (20, 15, 17) */,
  32'h3f2286f8 /* (16, 15, 17) */,
  32'h3efaa119 /* (12, 15, 17) */,
  32'h3e803f85 /* (8, 15, 17) */,
  32'h3e1fe07e /* (4, 15, 17) */,
  32'h3e086183 /* (0, 15, 17) */,
  32'h3ddcf428 /* (28, 11, 17) */,
  32'h3e2c9c6c /* (24, 11, 17) */,
  32'h3ea31756 /* (20, 11, 17) */,
  32'h3ecca1ac /* (16, 11, 17) */,
  32'h3ea31756 /* (12, 11, 17) */,
  32'h3e2c9c6c /* (8, 11, 17) */,
  32'h3ddcf428 /* (4, 11, 17) */,
  32'h3dbe6d47 /* (0, 11, 17) */,
  32'h3d7b9f11 /* (28, 7, 17) */,
  32'h3dbf0444 /* (24, 7, 17) */,
  32'h3e2e6a71 /* (20, 7, 17) */,
  32'h3e540b9b /* (16, 7, 17) */,
  32'h3e2e6a71 /* (12, 7, 17) */,
  32'h3dbf0444 /* (8, 7, 17) */,
  32'h3d7b9f11 /* (4, 7, 17) */,
  32'h3d5b6048 /* (0, 7, 17) */,
  32'h3d349293 /* (28, 3, 17) */,
  32'h3d8608f0 /* (24, 3, 17) */,
  32'h3deea44d /* (20, 3, 17) */,
  32'h3e0de417 /* (16, 3, 17) */,
  32'h3deea44d /* (12, 3, 17) */,
  32'h3d8608f0 /* (8, 3, 17) */,
  32'h3d349293 /* (4, 3, 17) */,
  32'h3d1eeabe /* (0, 3, 17) */,
  32'h3d2e802a /* (28, 31, 13) */,
  32'h3d7573b6 /* (24, 31, 13) */,
  32'h3dce8d02 /* (20, 31, 13) */,
  32'h3deaafef /* (16, 31, 13) */,
  32'h3dce8d02 /* (12, 31, 13) */,
  32'h3d7573b6 /* (8, 31, 13) */,
  32'h3d2e802a /* (4, 31, 13) */,
  32'h3d1d4601 /* (0, 31, 13) */,
  32'h3d4ea6a0 /* (28, 27, 13) */,
  32'h3d94d380 /* (24, 27, 13) */,
  32'h3e00477d /* (20, 27, 13) */,
  32'h3e1486b7 /* (16, 27, 13) */,
  32'h3e00477d /* (12, 27, 13) */,
  32'h3d94d380 /* (8, 27, 13) */,
  32'h3d4ea6a0 /* (4, 27, 13) */,
  32'h3d384488 /* (0, 27, 13) */,
  32'h3d9d0afa /* (28, 23, 13) */,
  32'h3deb6b6d /* (24, 23, 13) */,
  32'h3e53dc51 /* (20, 23, 13) */,
  32'h3e7e4b9d /* (16, 23, 13) */,
  32'h3e53dc51 /* (12, 23, 13) */,
  32'h3deb6b6d /* (8, 23, 13) */,
  32'h3d9d0afa /* (4, 23, 13) */,
  32'h3d89a49e /* (0, 23, 13) */,
  32'h3e0415cb /* (28, 19, 13) */,
  32'h3e4dd3dc /* (24, 19, 13) */,
  32'h3ec1d890 /* (20, 19, 13) */,
  32'h3ef27895 /* (16, 19, 13) */,
  32'h3ec1d890 /* (12, 19, 13) */,
  32'h3e4dd3dc /* (8, 19, 13) */,
  32'h3e0415cb /* (4, 19, 13) */,
  32'h3de3e928 /* (0, 19, 13) */,
  32'h3e0ff4ce /* (28, 15, 13) */,
  32'h3e640ba2 /* (24, 15, 13) */,
  32'h3edb3822 /* (20, 15, 13) */,
  32'h3f0bd969 /* (16, 15, 13) */,
  32'h3edb3822 /* (12, 15, 13) */,
  32'h3e640ba2 /* (8, 15, 13) */,
  32'h3e0ff4ce /* (4, 15, 13) */,
  32'h3df6cc6d /* (0, 15, 13) */,
  32'h3dcf13a3 /* (28, 11, 13) */,
  32'h3e1e607d /* (24, 11, 13) */,
  32'h3e91dfe2 /* (20, 11, 13) */,
  32'h3eb2bd2a /* (16, 11, 13) */,
  32'h3e91dfe2 /* (12, 11, 13) */,
  32'h3e1e607d /* (8, 11, 13) */,
  32'h3dcf13a3 /* (4, 11, 13) */,
  32'h3db3fd83 /* (0, 11, 13) */,
  32'h3d770afc /* (28, 7, 13) */,
  32'h3db56072 /* (24, 7, 13) */,
  32'h3e1f8cbf /* (20, 7, 13) */,
  32'h3e3bd4ee /* (16, 7, 13) */,
  32'h3e1f8cbf /* (12, 7, 13) */,
  32'h3db56072 /* (8, 7, 13) */,
  32'h3d770afc /* (4, 7, 13) */,
  32'h3d5a6fdd /* (0, 7, 13) */,
  32'h3d385879 /* (28, 3, 13) */,
  32'h3d82c188 /* (24, 3, 13) */,
  32'h3dddef48 /* (20, 3, 13) */,
  32'h3dfdd31f /* (16, 3, 13) */,
  32'h3dddef48 /* (12, 3, 13) */,
  32'h3d82c188 /* (8, 3, 13) */,
  32'h3d385879 /* (4, 3, 13) */,
  32'h3d258110 /* (0, 3, 13) */,
  32'h3d13f199 /* (28, 31, 9) */,
  32'h3d2fba80 /* (24, 31, 9) */,
  32'h3d803124 /* (20, 31, 9) */,
  32'h3d8420c9 /* (16, 31, 9) */,
  32'h3d803124 /* (12, 31, 9) */,
  32'h3d2fba80 /* (8, 31, 9) */,
  32'h3d13f199 /* (4, 31, 9) */,
  32'h3d11a5c6 /* (0, 31, 9) */,
  32'h3d1ee50b /* (28, 27, 9) */,
  32'h3d49c96c /* (24, 27, 9) */,
  32'h3d9af1c2 /* (20, 27, 9) */,
  32'h3da4f2f4 /* (16, 27, 9) */,
  32'h3d9af1c2 /* (12, 27, 9) */,
  32'h3d49c96c /* (8, 27, 9) */,
  32'h3d1ee50b /* (4, 27, 9) */,
  32'h3d16a564 /* (0, 27, 9) */,
  32'h3d51a9d2 /* (28, 23, 9) */,
  32'h3d921bde /* (24, 23, 9) */,
  32'h3df3b4f2 /* (20, 23, 9) */,
  32'h3e0981d7 /* (16, 23, 9) */,
  32'h3df3b4f2 /* (12, 23, 9) */,
  32'h3d921bde /* (8, 23, 9) */,
  32'h3d51a9d2 /* (4, 23, 9) */,
  32'h3d3dc47d /* (0, 23, 9) */,
  32'h3d9d0afa /* (28, 19, 9) */,
  32'h3deb6b6d /* (24, 19, 9) */,
  32'h3e53dc51 /* (20, 19, 9) */,
  32'h3e7e4b9d /* (16, 19, 9) */,
  32'h3e53dc51 /* (12, 19, 9) */,
  32'h3deb6b6d /* (8, 19, 9) */,
  32'h3d9d0afa /* (4, 19, 9) */,
  32'h3d89a49e /* (0, 19, 9) */,
  32'h3da3c1ed /* (28, 15, 9) */,
  32'h3dfc30a3 /* (24, 15, 9) */,
  32'h3e6a25fd /* (20, 15, 9) */,
  32'h3e908107 /* (16, 15, 9) */,
  32'h3e6a25fd /* (12, 15, 9) */,
  32'h3dfc30a3 /* (8, 15, 9) */,
  32'h3da3c1ed /* (4, 15, 9) */,
  32'h3d8df2c1 /* (0, 15, 9) */,
  32'h3d81d711 /* (28, 11, 9) */,
  32'h3dbc4d73 /* (24, 11, 9) */,
  32'h3e23781b /* (20, 11, 9) */,
  32'h3e3e5da7 /* (16, 11, 9) */,
  32'h3e23781b /* (12, 11, 9) */,
  32'h3dbc4d73 /* (8, 11, 9) */,
  32'h3d81d711 /* (4, 11, 9) */,
  32'h3d66dac1 /* (0, 11, 9) */,
  32'h3d30de15 /* (28, 7, 9) */,
  32'h3d6b8b35 /* (24, 7, 9) */,
  32'h3dbc51f9 /* (20, 7, 9) */,
  32'h3dce1075 /* (16, 7, 9) */,
  32'h3dbc51f9 /* (12, 7, 9) */,
  32'h3d6b8b35 /* (8, 7, 9) */,
  32'h3d30de15 /* (4, 7, 9) */,
  32'h3d23a039 /* (0, 7, 9) */,
  32'h3d16b5b2 /* (28, 3, 9) */,
  32'h3d37919e /* (24, 3, 9) */,
  32'h3d886b82 /* (20, 3, 9) */,
  32'h3d8e3848 /* (16, 3, 9) */,
  32'h3d886b82 /* (12, 3, 9) */,
  32'h3d37919e /* (8, 3, 9) */,
  32'h3d16b5b2 /* (4, 3, 9) */,
  32'h3d1237a7 /* (0, 3, 9) */,
  32'h3d334ee4 /* (28, 31, 5) */,
  32'h3d1412fd /* (24, 31, 5) */,
  32'h3d310ad3 /* (20, 31, 5) */,
  32'h3d24852f /* (16, 31, 5) */,
  32'h3d310ad3 /* (12, 31, 5) */,
  32'h3d1412fd /* (8, 31, 5) */,
  32'h3d334ee4 /* (4, 31, 5) */,
  32'h3d6e9998 /* (0, 31, 5) */,
  32'h3d189061 /* (28, 27, 5) */,
  32'h3d1c4d38 /* (24, 27, 5) */,
  32'h3d4f6dfc /* (20, 27, 5) */,
  32'h3d4ab7f7 /* (16, 27, 5) */,
  32'h3d4f6dfc /* (12, 27, 5) */,
  32'h3d1c4d38 /* (8, 27, 5) */,
  32'h3d189061 /* (4, 27, 5) */,
  32'h3d25e3da /* (0, 27, 5) */,
  32'h3d1ee50b /* (28, 23, 5) */,
  32'h3d49c96c /* (24, 23, 5) */,
  32'h3d9af1c2 /* (20, 23, 5) */,
  32'h3da4f2f4 /* (16, 23, 5) */,
  32'h3d9af1c2 /* (12, 23, 5) */,
  32'h3d49c96c /* (8, 23, 5) */,
  32'h3d1ee50b /* (4, 23, 5) */,
  32'h3d16a564 /* (0, 23, 5) */,
  32'h3d4ea6a0 /* (28, 19, 5) */,
  32'h3d94d380 /* (24, 19, 5) */,
  32'h3e00477d /* (20, 19, 5) */,
  32'h3e1486b7 /* (16, 19, 5) */,
  32'h3e00477d /* (12, 19, 5) */,
  32'h3d94d380 /* (8, 19, 5) */,
  32'h3d4ea6a0 /* (4, 19, 5) */,
  32'h3d384488 /* (0, 19, 5) */,
  32'h3d4def9b /* (28, 15, 5) */,
  32'h3d9a5b6b /* (24, 15, 5) */,
  32'h3e0ae903 /* (20, 15, 5) */,
  32'h3e26bbbb /* (16, 15, 5) */,
  32'h3e0ae903 /* (12, 15, 5) */,
  32'h3d9a5b6b /* (8, 15, 5) */,
  32'h3d4def9b /* (4, 15, 5) */,
  32'h3d347f0a /* (0, 15, 5) */,
  32'h3d358341 /* (28, 11, 5) */,
  32'h3d77c8fd /* (24, 11, 5) */,
  32'h3dca9d53 /* (20, 11, 5) */,
  32'h3de14ffa /* (16, 11, 5) */,
  32'h3dca9d53 /* (12, 11, 5) */,
  32'h3d77c8fd /* (8, 11, 5) */,
  32'h3d358341 /* (4, 11, 5) */,
  32'h3d25e815 /* (0, 11, 5) */,
  32'h3d1508af /* (28, 7, 5) */,
  32'h3d2bff3e /* (24, 7, 5) */,
  32'h3d75e4d4 /* (20, 7, 5) */,
  32'h3d7a662c /* (16, 7, 5) */,
  32'h3d75e4d4 /* (12, 7, 5) */,
  32'h3d2bff3e /* (8, 7, 5) */,
  32'h3d1508af /* (4, 7, 5) */,
  32'h3d154f7b /* (0, 7, 5) */,
  32'h3d25f5ce /* (28, 3, 5) */,
  32'h3d15d660 /* (24, 3, 5) */,
  32'h3d3a4ebb /* (20, 3, 5) */,
  32'h3d3046d8 /* (16, 3, 5) */,
  32'h3d3a4ebb /* (12, 3, 5) */,
  32'h3d15d660 /* (8, 3, 5) */,
  32'h3d25f5ce /* (4, 3, 5) */,
  32'h3d490b0e /* (0, 3, 5) */,
  32'h3d9c757b /* (28, 31, 1) */,
  32'h3d1704d7 /* (24, 31, 1) */,
  32'h3d1a2df1 /* (20, 31, 1) */,
  32'h3d067e68 /* (16, 31, 1) */,
  32'h3d1a2df1 /* (12, 31, 1) */,
  32'h3d1704d7 /* (8, 31, 1) */,
  32'h3d9c757b /* (4, 31, 1) */,
  32'h3f10fe39 /* (0, 31, 1) */,
  32'h3d334ee4 /* (28, 27, 1) */,
  32'h3d1412fd /* (24, 27, 1) */,
  32'h3d310ad3 /* (20, 27, 1) */,
  32'h3d24852f /* (16, 27, 1) */,
  32'h3d310ad3 /* (12, 27, 1) */,
  32'h3d1412fd /* (8, 27, 1) */,
  32'h3d334ee4 /* (4, 27, 1) */,
  32'h3d6e9998 /* (0, 27, 1) */,
  32'h3d13f199 /* (28, 23, 1) */,
  32'h3d2fba80 /* (24, 23, 1) */,
  32'h3d803124 /* (20, 23, 1) */,
  32'h3d8420c9 /* (16, 23, 1) */,
  32'h3d803124 /* (12, 23, 1) */,
  32'h3d2fba80 /* (8, 23, 1) */,
  32'h3d13f199 /* (4, 23, 1) */,
  32'h3d11a5c6 /* (0, 23, 1) */,
  32'h3d2e802a /* (28, 19, 1) */,
  32'h3d7573b6 /* (24, 19, 1) */,
  32'h3dce8d02 /* (20, 19, 1) */,
  32'h3deaafef /* (16, 19, 1) */,
  32'h3dce8d02 /* (12, 19, 1) */,
  32'h3d7573b6 /* (8, 19, 1) */,
  32'h3d2e802a /* (4, 19, 1) */,
  32'h3d1d4601 /* (0, 19, 1) */,
  32'h3d294c4b /* (28, 15, 1) */,
  32'h3d7a003f /* (24, 15, 1) */,
  32'h3ddd43c2 /* (20, 15, 1) */,
  32'h3e02e976 /* (16, 15, 1) */,
  32'h3ddd43c2 /* (12, 15, 1) */,
  32'h3d7a003f /* (8, 15, 1) */,
  32'h3d294c4b /* (4, 15, 1) */,
  32'h3d155505 /* (0, 15, 1) */,
  32'h3d1f5dc3 /* (28, 11, 1) */,
  32'h3d513c3d /* (24, 11, 1) */,
  32'h3da53628 /* (20, 11, 1) */,
  32'h3db336e0 /* (16, 11, 1) */,
  32'h3da53628 /* (12, 11, 1) */,
  32'h3d513c3d /* (8, 11, 1) */,
  32'h3d1f5dc3 /* (4, 11, 1) */,
  32'h3d147e90 /* (0, 11, 1) */,
  32'h3d17ff6b /* (28, 7, 1) */,
  32'h3d1bb8b6 /* (24, 7, 1) */,
  32'h3d4ea8e5 /* (20, 7, 1) */,
  32'h3d49f75a /* (16, 7, 1) */,
  32'h3d4ea8e5 /* (12, 7, 1) */,
  32'h3d1bb8b6 /* (8, 7, 1) */,
  32'h3d17ff6b /* (4, 7, 1) */,
  32'h3d25463b /* (0, 7, 1) */,
  32'h3d6eb36b /* (28, 3, 1) */,
  32'h3d146963 /* (24, 3, 1) */,
  32'h3d210eee /* (20, 3, 1) */,
  32'h3d0fbc59 /* (16, 3, 1) */,
  32'h3d210eee /* (12, 3, 1) */,
  32'h3d146963 /* (8, 3, 1) */,
  32'h3d6eb36b /* (4, 3, 1) */,
  32'h3dff9e3f /* (0, 3, 1) */,
  32'h3dbfa8df /* (31, 30, 29) */,
  32'h3d3cd255 /* (27, 30, 29) */,
  32'h3d12f42a /* (23, 30, 29) */,
  32'h3d29e985 /* (19, 30, 29) */,
  32'h3d240321 /* (15, 30, 29) */,
  32'h3d1c5f03 /* (11, 30, 29) */,
  32'h3d1a2949 /* (7, 30, 29) */,
  32'h3d866355 /* (3, 30, 29) */,
  32'h3d2ba889 /* (31, 26, 29) */,
  32'h3d16d305 /* (27, 26, 29) */,
  32'h3d215063 /* (23, 26, 29) */,
  32'h3d54a03b /* (19, 26, 29) */,
  32'h3d54ba37 /* (15, 26, 29) */,
  32'h3d39bb76 /* (11, 26, 29) */,
  32'h3d159d44 /* (7, 26, 29) */,
  32'h3d211f1b /* (3, 26, 29) */,
  32'h3d14c0fd /* (31, 22, 29) */,
  32'h3d2344c4 /* (27, 22, 29) */,
  32'h3d5dae2c /* (23, 22, 29) */,
  32'h3da99659 /* (19, 22, 29) */,
  32'h3db22d06 /* (15, 22, 29) */,
  32'h3d8ae43c /* (11, 22, 29) */,
  32'h3d387393 /* (7, 22, 29) */,
  32'h3d18cb02 /* (3, 22, 29) */,
  32'h3d276174 /* (31, 18, 29) */,
  32'h3d487174 /* (27, 18, 29) */,
  32'h3d9b2a7b /* (23, 18, 29) */,
  32'h3e04d0b8 /* (19, 18, 29) */,
  32'h3e11d12f /* (15, 18, 29) */,
  32'h3dce7d45 /* (11, 18, 29) */,
  32'h3d71c736 /* (7, 18, 29) */,
  32'h3d3188e3 /* (3, 18, 29) */,
  32'h3d276174 /* (31, 14, 29) */,
  32'h3d487174 /* (27, 14, 29) */,
  32'h3d9b2a7b /* (23, 14, 29) */,
  32'h3e04d0b8 /* (19, 14, 29) */,
  32'h3e11d12f /* (15, 14, 29) */,
  32'h3dce7d45 /* (11, 14, 29) */,
  32'h3d71c736 /* (7, 14, 29) */,
  32'h3d3188e3 /* (3, 14, 29) */,
  32'h3d14c0fd /* (31, 10, 29) */,
  32'h3d2344c4 /* (27, 10, 29) */,
  32'h3d5dae2c /* (23, 10, 29) */,
  32'h3da99659 /* (19, 10, 29) */,
  32'h3db22d06 /* (15, 10, 29) */,
  32'h3d8ae43c /* (11, 10, 29) */,
  32'h3d387393 /* (7, 10, 29) */,
  32'h3d18cb02 /* (3, 10, 29) */,
  32'h3d2ba889 /* (31, 6, 29) */,
  32'h3d16d305 /* (27, 6, 29) */,
  32'h3d215063 /* (23, 6, 29) */,
  32'h3d54a03b /* (19, 6, 29) */,
  32'h3d54ba37 /* (15, 6, 29) */,
  32'h3d39bb76 /* (11, 6, 29) */,
  32'h3d159d44 /* (7, 6, 29) */,
  32'h3d211f1b /* (3, 6, 29) */,
  32'h3dbfa8df /* (31, 2, 29) */,
  32'h3d3cd255 /* (27, 2, 29) */,
  32'h3d12f42a /* (23, 2, 29) */,
  32'h3d29e985 /* (19, 2, 29) */,
  32'h3d240321 /* (15, 2, 29) */,
  32'h3d1c5f03 /* (11, 2, 29) */,
  32'h3d1a2949 /* (7, 2, 29) */,
  32'h3d866355 /* (3, 2, 29) */,
  32'h3d20a35e /* (31, 30, 25) */,
  32'h3d14b1c0 /* (27, 30, 25) */,
  32'h3d26a1b5 /* (23, 30, 25) */,
  32'h3d6129ae /* (19, 30, 25) */,
  32'h3d62f778 /* (15, 30, 25) */,
  32'h3d42a7b8 /* (11, 30, 25) */,
  32'h3d1777c7 /* (7, 30, 25) */,
  32'h3d1a2949 /* (3, 30, 25) */,
  32'h3d146a43 /* (31, 26, 25) */,
  32'h3d1b2471 /* (27, 26, 25) */,
  32'h3d45eb5b /* (23, 26, 25) */,
  32'h3d90c8a7 /* (19, 26, 25) */,
  32'h3d95be73 /* (15, 26, 25) */,
  32'h3d71ecf9 /* (11, 26, 25) */,
  32'h3d29a602 /* (7, 26, 25) */,
  32'h3d159d44 /* (3, 26, 25) */,
  32'h3d305430 /* (31, 22, 25) */,
  32'h3d4b3dc7 /* (27, 22, 25) */,
  32'h3d94014f /* (23, 22, 25) */,
  32'h3defa49b /* (19, 22, 25) */,
  32'h3e009a19 /* (15, 22, 25) */,
  32'h3dbf3f1d /* (11, 22, 25) */,
  32'h3d6deb12 /* (7, 22, 25) */,
  32'h3d387393 /* (3, 22, 25) */,
  32'h3d62906c /* (31, 18, 25) */,
  32'h3d8a0000 /* (27, 18, 25) */,
  32'h3ddc09d8 /* (23, 18, 25) */,
  32'h3e41f14c /* (19, 18, 25) */,
  32'h3e57a44b /* (15, 18, 25) */,
  32'h3e14a5c9 /* (11, 18, 25) */,
  32'h3da8d240 /* (7, 18, 25) */,
  32'h3d71c736 /* (3, 18, 25) */,
  32'h3d62906c /* (31, 14, 25) */,
  32'h3d8a0000 /* (27, 14, 25) */,
  32'h3ddc09d8 /* (23, 14, 25) */,
  32'h3e41f14c /* (19, 14, 25) */,
  32'h3e57a44b /* (15, 14, 25) */,
  32'h3e14a5c9 /* (11, 14, 25) */,
  32'h3da8d240 /* (7, 14, 25) */,
  32'h3d71c736 /* (3, 14, 25) */,
  32'h3d305430 /* (31, 10, 25) */,
  32'h3d4b3dc7 /* (27, 10, 25) */,
  32'h3d94014f /* (23, 10, 25) */,
  32'h3defa49b /* (19, 10, 25) */,
  32'h3e009a19 /* (15, 10, 25) */,
  32'h3dbf3f1d /* (11, 10, 25) */,
  32'h3d6deb12 /* (7, 10, 25) */,
  32'h3d387393 /* (3, 10, 25) */,
  32'h3d146a43 /* (31, 6, 25) */,
  32'h3d1b2471 /* (27, 6, 25) */,
  32'h3d45eb5b /* (23, 6, 25) */,
  32'h3d90c8a7 /* (19, 6, 25) */,
  32'h3d95be73 /* (15, 6, 25) */,
  32'h3d71ecf9 /* (11, 6, 25) */,
  32'h3d29a602 /* (7, 6, 25) */,
  32'h3d159d44 /* (3, 6, 25) */,
  32'h3d20a35e /* (31, 2, 25) */,
  32'h3d14b1c0 /* (27, 2, 25) */,
  32'h3d26a1b5 /* (23, 2, 25) */,
  32'h3d6129ae /* (19, 2, 25) */,
  32'h3d62f778 /* (15, 2, 25) */,
  32'h3d42a7b8 /* (11, 2, 25) */,
  32'h3d1777c7 /* (7, 2, 25) */,
  32'h3d1a2949 /* (3, 2, 25) */,
  32'h3d16ed42 /* (31, 30, 21) */,
  32'h3d29823f /* (27, 30, 21) */,
  32'h3d6d9fa3 /* (23, 30, 21) */,
  32'h3dba5db4 /* (19, 30, 21) */,
  32'h3dc59b81 /* (15, 30, 21) */,
  32'h3d96eb50 /* (11, 30, 21) */,
  32'h3d42a7b8 /* (7, 30, 21) */,
  32'h3d1c5f03 /* (3, 30, 21) */,
  32'h3d31191b /* (31, 26, 21) */,
  32'h3d4d9045 /* (27, 26, 21) */,
  32'h3d9750ce /* (23, 26, 21) */,
  32'h3df74dbc /* (19, 26, 21) */,
  32'h3e0533d0 /* (15, 26, 21) */,
  32'h3dc480ba /* (11, 26, 21) */,
  32'h3d71ecf9 /* (7, 26, 21) */,
  32'h3d39bb76 /* (3, 26, 21) */,
  32'h3d829849 /* (31, 22, 21) */,
  32'h3d9d9380 /* (27, 22, 21) */,
  32'h3df71c69 /* (23, 22, 21) */,
  32'h3e562fb1 /* (19, 22, 21) */,
  32'h3e6c6ac0 /* (15, 22, 21) */,
  32'h3e257fc6 /* (11, 22, 21) */,
  32'h3dbf3f1d /* (7, 22, 21) */,
  32'h3d8ae43c /* (3, 22, 21) */,
  32'h3dc01db4 /* (31, 18, 21) */,
  32'h3deed79f /* (27, 18, 21) */,
  32'h3e458f30 /* (23, 18, 21) */,
  32'h3eb517ce /* (19, 18, 21) */,
  32'h3eccf8ff /* (15, 18, 21) */,
  32'h3e882756 /* (11, 18, 21) */,
  32'h3e14a5c9 /* (7, 18, 21) */,
  32'h3dce7d45 /* (3, 18, 21) */,
  32'h3dc01db4 /* (31, 14, 21) */,
  32'h3deed79f /* (27, 14, 21) */,
  32'h3e458f30 /* (23, 14, 21) */,
  32'h3eb517ce /* (19, 14, 21) */,
  32'h3eccf8ff /* (15, 14, 21) */,
  32'h3e882756 /* (11, 14, 21) */,
  32'h3e14a5c9 /* (7, 14, 21) */,
  32'h3dce7d45 /* (3, 14, 21) */,
  32'h3d829849 /* (31, 10, 21) */,
  32'h3d9d9380 /* (27, 10, 21) */,
  32'h3df71c69 /* (23, 10, 21) */,
  32'h3e562fb1 /* (19, 10, 21) */,
  32'h3e6c6ac0 /* (15, 10, 21) */,
  32'h3e257fc6 /* (11, 10, 21) */,
  32'h3dbf3f1d /* (7, 10, 21) */,
  32'h3d8ae43c /* (3, 10, 21) */,
  32'h3d31191b /* (31, 6, 21) */,
  32'h3d4d9045 /* (27, 6, 21) */,
  32'h3d9750ce /* (23, 6, 21) */,
  32'h3df74dbc /* (19, 6, 21) */,
  32'h3e0533d0 /* (15, 6, 21) */,
  32'h3dc480ba /* (11, 6, 21) */,
  32'h3d71ecf9 /* (7, 6, 21) */,
  32'h3d39bb76 /* (3, 6, 21) */,
  32'h3d16ed42 /* (31, 2, 21) */,
  32'h3d29823f /* (27, 2, 21) */,
  32'h3d6d9fa3 /* (23, 2, 21) */,
  32'h3dba5db4 /* (19, 2, 21) */,
  32'h3dc59b81 /* (15, 2, 21) */,
  32'h3d96eb50 /* (11, 2, 21) */,
  32'h3d42a7b8 /* (7, 2, 21) */,
  32'h3d1c5f03 /* (3, 2, 21) */,
  32'h3d1a0745 /* (31, 30, 17) */,
  32'h3d3a7be5 /* (27, 30, 17) */,
  32'h3d9314c2 /* (23, 30, 17) */,
  32'h3e003b1e /* (19, 30, 17) */,
  32'h3e0de5f8 /* (15, 30, 17) */,
  32'h3dc59b81 /* (11, 30, 17) */,
  32'h3d62f778 /* (7, 30, 17) */,
  32'h3d240321 /* (3, 30, 17) */,
  32'h3d46f53f /* (31, 26, 17) */,
  32'h3d73b16f /* (27, 26, 17) */,
  32'h3dc42ad0 /* (23, 26, 17) */,
  32'h3e2ea39a /* (19, 26, 17) */,
  32'h3e430b11 /* (15, 26, 17) */,
  32'h3e0533d0 /* (11, 26, 17) */,
  32'h3d95be73 /* (7, 26, 17) */,
  32'h3d54ba37 /* (3, 26, 17) */,
  32'h3da5ac70 /* (31, 22, 17) */,
  32'h3dce52e6 /* (27, 22, 17) */,
  32'h3e2b3653 /* (23, 22, 17) */,
  32'h3e9d80fb /* (19, 22, 17) */,
  32'h3eb2925b /* (15, 22, 17) */,
  32'h3e6c6ac0 /* (11, 22, 17) */,
  32'h3e009a19 /* (7, 22, 17) */,
  32'h3db22d06 /* (3, 22, 17) */,
  32'h3e06d8bb /* (31, 18, 17) */,
  32'h3e2a981c /* (27, 18, 17) */,
  32'h3e91e4f8 /* (23, 18, 17) */,
  32'h3f0af24f /* (19, 18, 17) */,
  32'h3f202f9a /* (15, 18, 17) */,
  32'h3eccf8ff /* (11, 18, 17) */,
  32'h3e57a44b /* (7, 18, 17) */,
  32'h3e11d12f /* (3, 18, 17) */,
  32'h3e06d8bb /* (31, 14, 17) */,
  32'h3e2a981c /* (27, 14, 17) */,
  32'h3e91e4f8 /* (23, 14, 17) */,
  32'h3f0af24f /* (19, 14, 17) */,
  32'h3f202f9a /* (15, 14, 17) */,
  32'h3eccf8ff /* (11, 14, 17) */,
  32'h3e57a44b /* (7, 14, 17) */,
  32'h3e11d12f /* (3, 14, 17) */,
  32'h3da5ac70 /* (31, 10, 17) */,
  32'h3dce52e6 /* (27, 10, 17) */,
  32'h3e2b3653 /* (23, 10, 17) */,
  32'h3e9d80fb /* (19, 10, 17) */,
  32'h3eb2925b /* (15, 10, 17) */,
  32'h3e6c6ac0 /* (11, 10, 17) */,
  32'h3e009a19 /* (7, 10, 17) */,
  32'h3db22d06 /* (3, 10, 17) */,
  32'h3d46f53f /* (31, 6, 17) */,
  32'h3d73b16f /* (27, 6, 17) */,
  32'h3dc42ad0 /* (23, 6, 17) */,
  32'h3e2ea39a /* (19, 6, 17) */,
  32'h3e430b11 /* (15, 6, 17) */,
  32'h3e0533d0 /* (11, 6, 17) */,
  32'h3d95be73 /* (7, 6, 17) */,
  32'h3d54ba37 /* (3, 6, 17) */,
  32'h3d1a0745 /* (31, 2, 17) */,
  32'h3d3a7be5 /* (27, 2, 17) */,
  32'h3d9314c2 /* (23, 2, 17) */,
  32'h3e003b1e /* (19, 2, 17) */,
  32'h3e0de5f8 /* (15, 2, 17) */,
  32'h3dc59b81 /* (11, 2, 17) */,
  32'h3d62f778 /* (7, 2, 17) */,
  32'h3d240321 /* (3, 2, 17) */,
  32'h3d214ba3 /* (31, 30, 13) */,
  32'h3d3d84de /* (27, 30, 13) */,
  32'h3d8e358b /* (23, 30, 13) */,
  32'h3dec70da /* (19, 30, 13) */,
  32'h3e003b1e /* (15, 30, 13) */,
  32'h3dba5db4 /* (11, 30, 13) */,
  32'h3d6129ae /* (7, 30, 13) */,
  32'h3d29e985 /* (3, 30, 13) */,
  32'h3d4876ff /* (31, 26, 13) */,
  32'h3d700ffa /* (27, 26, 13) */,
  32'h3db9d5f4 /* (23, 26, 13) */,
  32'h3e1f113d /* (19, 26, 13) */,
  32'h3e2ea39a /* (15, 26, 13) */,
  32'h3df74dbc /* (11, 26, 13) */,
  32'h3d90c8a7 /* (7, 26, 13) */,
  32'h3d54a03b /* (3, 26, 13) */,
  32'h3d9e7894 /* (31, 22, 13) */,
  32'h3dc29629 /* (27, 22, 13) */,
  32'h3e1d56b2 /* (23, 22, 13) */,
  32'h3e8cbae1 /* (19, 22, 13) */,
  32'h3e9d80fb /* (15, 22, 13) */,
  32'h3e562fb1 /* (11, 22, 13) */,
  32'h3defa49b /* (7, 22, 13) */,
  32'h3da99659 /* (3, 22, 13) */,
  32'h3df65860 /* (31, 18, 13) */,
  32'h3e1a8d8c /* (27, 18, 13) */,
  32'h3e821787 /* (23, 18, 13) */,
  32'h3ef33ce4 /* (19, 18, 13) */,
  32'h3f0af24f /* (15, 18, 13) */,
  32'h3eb517ce /* (11, 18, 13) */,
  32'h3e41f14c /* (7, 18, 13) */,
  32'h3e04d0b8 /* (3, 18, 13) */,
  32'h3df65860 /* (31, 14, 13) */,
  32'h3e1a8d8c /* (27, 14, 13) */,
  32'h3e821787 /* (23, 14, 13) */,
  32'h3ef33ce4 /* (19, 14, 13) */,
  32'h3f0af24f /* (15, 14, 13) */,
  32'h3eb517ce /* (11, 14, 13) */,
  32'h3e41f14c /* (7, 14, 13) */,
  32'h3e04d0b8 /* (3, 14, 13) */,
  32'h3d9e7894 /* (31, 10, 13) */,
  32'h3dc29629 /* (27, 10, 13) */,
  32'h3e1d56b2 /* (23, 10, 13) */,
  32'h3e8cbae1 /* (19, 10, 13) */,
  32'h3e9d80fb /* (15, 10, 13) */,
  32'h3e562fb1 /* (11, 10, 13) */,
  32'h3defa49b /* (7, 10, 13) */,
  32'h3da99659 /* (3, 10, 13) */,
  32'h3d4876ff /* (31, 6, 13) */,
  32'h3d700ffa /* (27, 6, 13) */,
  32'h3db9d5f4 /* (23, 6, 13) */,
  32'h3e1f113d /* (19, 6, 13) */,
  32'h3e2ea39a /* (15, 6, 13) */,
  32'h3df74dbc /* (11, 6, 13) */,
  32'h3d90c8a7 /* (7, 6, 13) */,
  32'h3d54a03b /* (3, 6, 13) */,
  32'h3d214ba3 /* (31, 2, 13) */,
  32'h3d3d84de /* (27, 2, 13) */,
  32'h3d8e358b /* (23, 2, 13) */,
  32'h3dec70da /* (19, 2, 13) */,
  32'h3e003b1e /* (15, 2, 13) */,
  32'h3dba5db4 /* (11, 2, 13) */,
  32'h3d6129ae /* (7, 2, 13) */,
  32'h3d29e985 /* (3, 2, 13) */,
  32'h3d11c69f /* (31, 30, 9) */,
  32'h3d18622e /* (27, 30, 9) */,
  32'h3d42665b /* (23, 30, 9) */,
  32'h3d8e358b /* (19, 30, 9) */,
  32'h3d9314c2 /* (15, 30, 9) */,
  32'h3d6d9fa3 /* (11, 30, 9) */,
  32'h3d26a1b5 /* (7, 30, 9) */,
  32'h3d12f42a /* (3, 30, 9) */,
  32'h3d1c53e8 /* (31, 26, 9) */,
  32'h3d2db0cc /* (27, 26, 9) */,
  32'h3d6fd024 /* (23, 26, 9) */,
  32'h3db9d5f4 /* (19, 26, 9) */,
  32'h3dc42ad0 /* (15, 26, 9) */,
  32'h3d9750ce /* (11, 26, 9) */,
  32'h3d45eb5b /* (7, 26, 9) */,
  32'h3d215063 /* (3, 26, 9) */,
  32'h3d52081f /* (31, 22, 9) */,
  32'h3d781ae6 /* (27, 22, 9) */,
  32'h3dbbc730 /* (23, 22, 9) */,
  32'h3e1d56b2 /* (19, 22, 9) */,
  32'h3e2b3653 /* (15, 22, 9) */,
  32'h3df71c69 /* (11, 22, 9) */,
  32'h3d94014f /* (7, 22, 9) */,
  32'h3d5dae2c /* (3, 22, 9) */,
  32'h3d90dff9 /* (31, 18, 9) */,
  32'h3db24f8e /* (27, 18, 9) */,
  32'h3e10cac5 /* (23, 18, 9) */,
  32'h3e821787 /* (19, 18, 9) */,
  32'h3e91e4f8 /* (15, 18, 9) */,
  32'h3e458f30 /* (11, 18, 9) */,
  32'h3ddc09d8 /* (7, 18, 9) */,
  32'h3d9b2a7b /* (3, 18, 9) */,
  32'h3d90dff9 /* (31, 14, 9) */,
  32'h3db24f8e /* (27, 14, 9) */,
  32'h3e10cac5 /* (23, 14, 9) */,
  32'h3e821787 /* (19, 14, 9) */,
  32'h3e91e4f8 /* (15, 14, 9) */,
  32'h3e458f30 /* (11, 14, 9) */,
  32'h3ddc09d8 /* (7, 14, 9) */,
  32'h3d9b2a7b /* (3, 14, 9) */,
  32'h3d52081f /* (31, 10, 9) */,
  32'h3d781ae6 /* (27, 10, 9) */,
  32'h3dbbc730 /* (23, 10, 9) */,
  32'h3e1d56b2 /* (19, 10, 9) */,
  32'h3e2b3653 /* (15, 10, 9) */,
  32'h3df71c69 /* (11, 10, 9) */,
  32'h3d94014f /* (7, 10, 9) */,
  32'h3d5dae2c /* (3, 10, 9) */,
  32'h3d1c53e8 /* (31, 6, 9) */,
  32'h3d2db0cc /* (27, 6, 9) */,
  32'h3d6fd024 /* (23, 6, 9) */,
  32'h3db9d5f4 /* (19, 6, 9) */,
  32'h3dc42ad0 /* (15, 6, 9) */,
  32'h3d9750ce /* (11, 6, 9) */,
  32'h3d45eb5b /* (7, 6, 9) */,
  32'h3d215063 /* (3, 6, 9) */,
  32'h3d11c69f /* (31, 2, 9) */,
  32'h3d18622e /* (27, 2, 9) */,
  32'h3d42665b /* (23, 2, 9) */,
  32'h3d8e358b /* (19, 2, 9) */,
  32'h3d9314c2 /* (15, 2, 9) */,
  32'h3d6d9fa3 /* (11, 2, 9) */,
  32'h3d26a1b5 /* (7, 2, 9) */,
  32'h3d12f42a /* (3, 2, 9) */,
  32'h3d59109a /* (31, 30, 5) */,
  32'h3d213c91 /* (27, 30, 5) */,
  32'h3d18622e /* (23, 30, 5) */,
  32'h3d3d84de /* (19, 30, 5) */,
  32'h3d3a7be5 /* (15, 30, 5) */,
  32'h3d29823f /* (11, 30, 5) */,
  32'h3d14b1c0 /* (7, 30, 5) */,
  32'h3d3cd255 /* (3, 30, 5) */,
  32'h3d1a8b5a /* (31, 26, 5) */,
  32'h3d14f7ce /* (27, 26, 5) */,
  32'h3d2db0cc /* (23, 26, 5) */,
  32'h3d700ffa /* (19, 26, 5) */,
  32'h3d73b16f /* (15, 26, 5) */,
  32'h3d4d9045 /* (11, 26, 5) */,
  32'h3d1b2471 /* (7, 26, 5) */,
  32'h3d16d305 /* (3, 26, 5) */,
  32'h3d1d9589 /* (31, 22, 5) */,
  32'h3d30fc5a /* (27, 22, 5) */,
  32'h3d781ae6 /* (23, 22, 5) */,
  32'h3dc29629 /* (19, 22, 5) */,
  32'h3dce52e6 /* (15, 22, 5) */,
  32'h3d9d9380 /* (11, 22, 5) */,
  32'h3d4b3dc7 /* (7, 22, 5) */,
  32'h3d2344c4 /* (3, 22, 5) */,
  32'h3d3c7841 /* (31, 18, 5) */,
  32'h3d63687e /* (27, 18, 5) */,
  32'h3db24f8e /* (23, 18, 5) */,
  32'h3e1a8d8c /* (19, 18, 5) */,
  32'h3e2a981c /* (15, 18, 5) */,
  32'h3deed79f /* (11, 18, 5) */,
  32'h3d8a0000 /* (7, 18, 5) */,
  32'h3d487174 /* (3, 18, 5) */,
  32'h3d3c7841 /* (31, 14, 5) */,
  32'h3d63687e /* (27, 14, 5) */,
  32'h3db24f8e /* (23, 14, 5) */,
  32'h3e1a8d8c /* (19, 14, 5) */,
  32'h3e2a981c /* (15, 14, 5) */,
  32'h3deed79f /* (11, 14, 5) */,
  32'h3d8a0000 /* (7, 14, 5) */,
  32'h3d487174 /* (3, 14, 5) */,
  32'h3d1d9589 /* (31, 10, 5) */,
  32'h3d30fc5a /* (27, 10, 5) */,
  32'h3d781ae6 /* (23, 10, 5) */,
  32'h3dc29629 /* (19, 10, 5) */,
  32'h3dce52e6 /* (15, 10, 5) */,
  32'h3d9d9380 /* (11, 10, 5) */,
  32'h3d4b3dc7 /* (7, 10, 5) */,
  32'h3d2344c4 /* (3, 10, 5) */,
  32'h3d1a8b5a /* (31, 6, 5) */,
  32'h3d14f7ce /* (27, 6, 5) */,
  32'h3d2db0cc /* (23, 6, 5) */,
  32'h3d700ffa /* (19, 6, 5) */,
  32'h3d73b16f /* (15, 6, 5) */,
  32'h3d4d9045 /* (11, 6, 5) */,
  32'h3d1b2471 /* (7, 6, 5) */,
  32'h3d16d305 /* (3, 6, 5) */,
  32'h3d59109a /* (31, 2, 5) */,
  32'h3d213c91 /* (27, 2, 5) */,
  32'h3d18622e /* (23, 2, 5) */,
  32'h3d3d84de /* (19, 2, 5) */,
  32'h3d3a7be5 /* (15, 2, 5) */,
  32'h3d29823f /* (11, 2, 5) */,
  32'h3d14b1c0 /* (7, 2, 5) */,
  32'h3d3cd255 /* (3, 2, 5) */,
  32'h3e4aeee2 /* (31, 30, 1) */,
  32'h3d59109a /* (27, 30, 1) */,
  32'h3d11c69f /* (23, 30, 1) */,
  32'h3d214ba3 /* (19, 30, 1) */,
  32'h3d1a0745 /* (15, 30, 1) */,
  32'h3d16ed42 /* (11, 30, 1) */,
  32'h3d20a35e /* (7, 30, 1) */,
  32'h3dbfa8df /* (3, 30, 1) */,
  32'h3d3c9698 /* (31, 26, 1) */,
  32'h3d1a8b5a /* (27, 26, 1) */,
  32'h3d1c53e8 /* (23, 26, 1) */,
  32'h3d4876ff /* (19, 26, 1) */,
  32'h3d46f53f /* (15, 26, 1) */,
  32'h3d31191b /* (11, 26, 1) */,
  32'h3d146a43 /* (7, 26, 1) */,
  32'h3d2ba889 /* (3, 26, 1) */,
  32'h3d119771 /* (31, 22, 1) */,
  32'h3d1d9589 /* (27, 22, 1) */,
  32'h3d52081f /* (23, 22, 1) */,
  32'h3d9e7894 /* (19, 22, 1) */,
  32'h3da5ac70 /* (15, 22, 1) */,
  32'h3d829849 /* (11, 22, 1) */,
  32'h3d305430 /* (7, 22, 1) */,
  32'h3d14c0fd /* (3, 22, 1) */,
  32'h3d1e0bb6 /* (31, 18, 1) */,
  32'h3d3c7841 /* (27, 18, 1) */,
  32'h3d90dff9 /* (23, 18, 1) */,
  32'h3df65860 /* (19, 18, 1) */,
  32'h3e06d8bb /* (15, 18, 1) */,
  32'h3dc01db4 /* (11, 18, 1) */,
  32'h3d62906c /* (7, 18, 1) */,
  32'h3d276174 /* (3, 18, 1) */,
  32'h3d1e0bb6 /* (31, 14, 1) */,
  32'h3d3c7841 /* (27, 14, 1) */,
  32'h3d90dff9 /* (23, 14, 1) */,
  32'h3df65860 /* (19, 14, 1) */,
  32'h3e06d8bb /* (15, 14, 1) */,
  32'h3dc01db4 /* (11, 14, 1) */,
  32'h3d62906c /* (7, 14, 1) */,
  32'h3d276174 /* (3, 14, 1) */,
  32'h3d119771 /* (31, 10, 1) */,
  32'h3d1d9589 /* (27, 10, 1) */,
  32'h3d52081f /* (23, 10, 1) */,
  32'h3d9e7894 /* (19, 10, 1) */,
  32'h3da5ac70 /* (15, 10, 1) */,
  32'h3d829849 /* (11, 10, 1) */,
  32'h3d305430 /* (7, 10, 1) */,
  32'h3d14c0fd /* (3, 10, 1) */,
  32'h3d3c9698 /* (31, 6, 1) */,
  32'h3d1a8b5a /* (27, 6, 1) */,
  32'h3d1c53e8 /* (23, 6, 1) */,
  32'h3d4876ff /* (19, 6, 1) */,
  32'h3d46f53f /* (15, 6, 1) */,
  32'h3d31191b /* (11, 6, 1) */,
  32'h3d146a43 /* (7, 6, 1) */,
  32'h3d2ba889 /* (3, 6, 1) */,
  32'h3e4aeee2 /* (31, 2, 1) */,
  32'h3d59109a /* (27, 2, 1) */,
  32'h3d11c69f /* (23, 2, 1) */,
  32'h3d214ba3 /* (19, 2, 1) */,
  32'h3d1a0745 /* (15, 2, 1) */,
  32'h3d16ed42 /* (11, 2, 1) */,
  32'h3d20a35e /* (7, 2, 1) */,
  32'h3dbfa8df /* (3, 2, 1) */,
  32'h3da3af74 /* (30, 30, 29) */,
  32'h3d271e8d /* (26, 30, 29) */,
  32'h3d162b76 /* (22, 30, 29) */,
  32'h3d2b1735 /* (18, 30, 29) */,
  32'h3d2b1735 /* (14, 30, 29) */,
  32'h3d162b76 /* (10, 30, 29) */,
  32'h3d271e8d /* (6, 30, 29) */,
  32'h3da3af74 /* (2, 30, 29) */,
  32'h3d271e8d /* (30, 26, 29) */,
  32'h3d14c14d /* (26, 26, 29) */,
  32'h3d2c3293 /* (22, 26, 29) */,
  32'h3d5a5169 /* (18, 26, 29) */,
  32'h3d5a5169 /* (14, 26, 29) */,
  32'h3d2c3293 /* (10, 26, 29) */,
  32'h3d14c14d /* (6, 26, 29) */,
  32'h3d271e8d /* (2, 26, 29) */,
  32'h3d162b76 /* (30, 22, 29) */,
  32'h3d2c3293 /* (26, 22, 29) */,
  32'h3d77904c /* (22, 22, 29) */,
  32'h3db2bcb9 /* (18, 22, 29) */,
  32'h3db2bcb9 /* (14, 22, 29) */,
  32'h3d77904c /* (10, 22, 29) */,
  32'h3d2c3293 /* (6, 22, 29) */,
  32'h3d162b76 /* (2, 22, 29) */,
  32'h3d2b1735 /* (30, 18, 29) */,
  32'h3d5a5169 /* (26, 18, 29) */,
  32'h3db2bcb9 /* (22, 18, 29) */,
  32'h3e0f3c67 /* (18, 18, 29) */,
  32'h3e0f3c67 /* (14, 18, 29) */,
  32'h3db2bcb9 /* (10, 18, 29) */,
  32'h3d5a5169 /* (6, 18, 29) */,
  32'h3d2b1735 /* (2, 18, 29) */,
  32'h3d2b1735 /* (30, 14, 29) */,
  32'h3d5a5169 /* (26, 14, 29) */,
  32'h3db2bcb9 /* (22, 14, 29) */,
  32'h3e0f3c67 /* (18, 14, 29) */,
  32'h3e0f3c67 /* (14, 14, 29) */,
  32'h3db2bcb9 /* (10, 14, 29) */,
  32'h3d5a5169 /* (6, 14, 29) */,
  32'h3d2b1735 /* (2, 14, 29) */,
  32'h3d162b76 /* (30, 10, 29) */,
  32'h3d2c3293 /* (26, 10, 29) */,
  32'h3d77904c /* (22, 10, 29) */,
  32'h3db2bcb9 /* (18, 10, 29) */,
  32'h3db2bcb9 /* (14, 10, 29) */,
  32'h3d77904c /* (10, 10, 29) */,
  32'h3d2c3293 /* (6, 10, 29) */,
  32'h3d162b76 /* (2, 10, 29) */,
  32'h3d271e8d /* (30, 6, 29) */,
  32'h3d14c14d /* (26, 6, 29) */,
  32'h3d2c3293 /* (22, 6, 29) */,
  32'h3d5a5169 /* (18, 6, 29) */,
  32'h3d5a5169 /* (14, 6, 29) */,
  32'h3d2c3293 /* (10, 6, 29) */,
  32'h3d14c14d /* (6, 6, 29) */,
  32'h3d271e8d /* (2, 6, 29) */,
  32'h3da3af74 /* (30, 2, 29) */,
  32'h3d271e8d /* (26, 2, 29) */,
  32'h3d162b76 /* (22, 2, 29) */,
  32'h3d2b1735 /* (18, 2, 29) */,
  32'h3d2b1735 /* (14, 2, 29) */,
  32'h3d162b76 /* (10, 2, 29) */,
  32'h3d271e8d /* (6, 2, 29) */,
  32'h3da3af74 /* (2, 2, 29) */,
  32'h3d1dd271 /* (30, 30, 25) */,
  32'h3d14b9d3 /* (26, 30, 25) */,
  32'h3d3346c6 /* (22, 30, 25) */,
  32'h3d6820b1 /* (18, 30, 25) */,
  32'h3d6820b1 /* (14, 30, 25) */,
  32'h3d3346c6 /* (10, 30, 25) */,
  32'h3d14b9d3 /* (6, 30, 25) */,
  32'h3d1dd271 /* (2, 30, 25) */,
  32'h3d14b9d3 /* (30, 26, 25) */,
  32'h3d20f672 /* (26, 26, 25) */,
  32'h3d5a2934 /* (22, 26, 25) */,
  32'h3d975464 /* (18, 26, 25) */,
  32'h3d975464 /* (14, 26, 25) */,
  32'h3d5a2934 /* (10, 26, 25) */,
  32'h3d20f672 /* (6, 26, 25) */,
  32'h3d14b9d3 /* (2, 26, 25) */,
  32'h3d3346c6 /* (30, 22, 25) */,
  32'h3d5a2934 /* (26, 22, 25) */,
  32'h3da7f0fb /* (22, 22, 25) */,
  32'h3dff6ab3 /* (18, 22, 25) */,
  32'h3dff6ab3 /* (14, 22, 25) */,
  32'h3da7f0fb /* (10, 22, 25) */,
  32'h3d5a2934 /* (6, 22, 25) */,
  32'h3d3346c6 /* (2, 22, 25) */,
  32'h3d6820b1 /* (30, 18, 25) */,
  32'h3d975464 /* (26, 18, 25) */,
  32'h3dff6ab3 /* (22, 18, 25) */,
  32'h3e528761 /* (18, 18, 25) */,
  32'h3e528761 /* (14, 18, 25) */,
  32'h3dff6ab3 /* (10, 18, 25) */,
  32'h3d975464 /* (6, 18, 25) */,
  32'h3d6820b1 /* (2, 18, 25) */,
  32'h3d6820b1 /* (30, 14, 25) */,
  32'h3d975464 /* (26, 14, 25) */,
  32'h3dff6ab3 /* (22, 14, 25) */,
  32'h3e528761 /* (18, 14, 25) */,
  32'h3e528761 /* (14, 14, 25) */,
  32'h3dff6ab3 /* (10, 14, 25) */,
  32'h3d975464 /* (6, 14, 25) */,
  32'h3d6820b1 /* (2, 14, 25) */,
  32'h3d3346c6 /* (30, 10, 25) */,
  32'h3d5a2934 /* (26, 10, 25) */,
  32'h3da7f0fb /* (22, 10, 25) */,
  32'h3dff6ab3 /* (18, 10, 25) */,
  32'h3dff6ab3 /* (14, 10, 25) */,
  32'h3da7f0fb /* (10, 10, 25) */,
  32'h3d5a2934 /* (6, 10, 25) */,
  32'h3d3346c6 /* (2, 10, 25) */,
  32'h3d14b9d3 /* (30, 6, 25) */,
  32'h3d20f672 /* (26, 6, 25) */,
  32'h3d5a2934 /* (22, 6, 25) */,
  32'h3d975464 /* (18, 6, 25) */,
  32'h3d975464 /* (14, 6, 25) */,
  32'h3d5a2934 /* (10, 6, 25) */,
  32'h3d20f672 /* (6, 6, 25) */,
  32'h3d14b9d3 /* (2, 6, 25) */,
  32'h3d1dd271 /* (30, 2, 25) */,
  32'h3d14b9d3 /* (26, 2, 25) */,
  32'h3d3346c6 /* (22, 2, 25) */,
  32'h3d6820b1 /* (18, 2, 25) */,
  32'h3d6820b1 /* (14, 2, 25) */,
  32'h3d3346c6 /* (10, 2, 25) */,
  32'h3d14b9d3 /* (6, 2, 25) */,
  32'h3d1dd271 /* (2, 2, 25) */,
  32'h3d18e0f8 /* (30, 30, 21) */,
  32'h3d343ccb /* (26, 30, 21) */,
  32'h3d85a0b3 /* (22, 30, 21) */,
  32'h3dc55f41 /* (18, 30, 21) */,
  32'h3dc55f41 /* (14, 30, 21) */,
  32'h3d85a0b3 /* (10, 30, 21) */,
  32'h3d343ccb /* (6, 30, 21) */,
  32'h3d18e0f8 /* (2, 30, 21) */,
  32'h3d343ccb /* (30, 26, 21) */,
  32'h3d5d3b5c /* (26, 26, 21) */,
  32'h3dac23aa /* (22, 26, 21) */,
  32'h3e040b60 /* (18, 26, 21) */,
  32'h3e040b60 /* (14, 26, 21) */,
  32'h3dac23aa /* (10, 26, 21) */,
  32'h3d5d3b5c /* (6, 26, 21) */,
  32'h3d343ccb /* (2, 26, 21) */,
  32'h3d85a0b3 /* (30, 22, 21) */,
  32'h3dac23aa /* (26, 22, 21) */,
  32'h3e0ecbcd /* (22, 22, 21) */,
  32'h3e67a191 /* (18, 22, 21) */,
  32'h3e67a191 /* (14, 22, 21) */,
  32'h3e0ecbcd /* (10, 22, 21) */,
  32'h3dac23aa /* (6, 22, 21) */,
  32'h3d85a0b3 /* (2, 22, 21) */,
  32'h3dc55f41 /* (30, 18, 21) */,
  32'h3e040b60 /* (26, 18, 21) */,
  32'h3e67a191 /* (22, 18, 21) */,
  32'h3ec66134 /* (18, 18, 21) */,
  32'h3ec66134 /* (14, 18, 21) */,
  32'h3e67a191 /* (10, 18, 21) */,
  32'h3e040b60 /* (6, 18, 21) */,
  32'h3dc55f41 /* (2, 18, 21) */,
  32'h3dc55f41 /* (30, 14, 21) */,
  32'h3e040b60 /* (26, 14, 21) */,
  32'h3e67a191 /* (22, 14, 21) */,
  32'h3ec66134 /* (18, 14, 21) */,
  32'h3ec66134 /* (14, 14, 21) */,
  32'h3e67a191 /* (10, 14, 21) */,
  32'h3e040b60 /* (6, 14, 21) */,
  32'h3dc55f41 /* (2, 14, 21) */,
  32'h3d85a0b3 /* (30, 10, 21) */,
  32'h3dac23aa /* (26, 10, 21) */,
  32'h3e0ecbcd /* (22, 10, 21) */,
  32'h3e67a191 /* (18, 10, 21) */,
  32'h3e67a191 /* (14, 10, 21) */,
  32'h3e0ecbcd /* (10, 10, 21) */,
  32'h3dac23aa /* (6, 10, 21) */,
  32'h3d85a0b3 /* (2, 10, 21) */,
  32'h3d343ccb /* (30, 6, 21) */,
  32'h3d5d3b5c /* (26, 6, 21) */,
  32'h3dac23aa /* (22, 6, 21) */,
  32'h3e040b60 /* (18, 6, 21) */,
  32'h3e040b60 /* (14, 6, 21) */,
  32'h3dac23aa /* (10, 6, 21) */,
  32'h3d5d3b5c /* (6, 6, 21) */,
  32'h3d343ccb /* (2, 6, 21) */,
  32'h3d18e0f8 /* (30, 2, 21) */,
  32'h3d343ccb /* (26, 2, 21) */,
  32'h3d85a0b3 /* (22, 2, 21) */,
  32'h3dc55f41 /* (18, 2, 21) */,
  32'h3dc55f41 /* (14, 2, 21) */,
  32'h3d85a0b3 /* (10, 2, 21) */,
  32'h3d343ccb /* (6, 2, 21) */,
  32'h3d18e0f8 /* (2, 2, 21) */,
  32'h3d1dadb9 /* (30, 30, 17) */,
  32'h3d4bfe66 /* (26, 30, 17) */,
  32'h3daa3ec9 /* (22, 30, 17) */,
  32'h3e0adb0d /* (18, 30, 17) */,
  32'h3e0adb0d /* (14, 30, 17) */,
  32'h3daa3ec9 /* (10, 30, 17) */,
  32'h3d4bfe66 /* (6, 30, 17) */,
  32'h3d1dadb9 /* (2, 30, 17) */,
  32'h3d4bfe66 /* (30, 26, 17) */,
  32'h3d85e8bf /* (26, 26, 17) */,
  32'h3de44bb3 /* (22, 26, 17) */,
  32'h3e3e01e0 /* (18, 26, 17) */,
  32'h3e3e01e0 /* (14, 26, 17) */,
  32'h3de44bb3 /* (10, 26, 17) */,
  32'h3d85e8bf /* (6, 26, 17) */,
  32'h3d4bfe66 /* (2, 26, 17) */,
  32'h3daa3ec9 /* (30, 22, 17) */,
  32'h3de44bb3 /* (26, 22, 17) */,
  32'h3e48eba4 /* (22, 22, 17) */,
  32'h3eacaf9b /* (18, 22, 17) */,
  32'h3eacaf9b /* (14, 22, 17) */,
  32'h3e48eba4 /* (10, 22, 17) */,
  32'h3de44bb3 /* (6, 22, 17) */,
  32'h3daa3ec9 /* (2, 22, 17) */,
  32'h3e0adb0d /* (30, 18, 17) */,
  32'h3e3e01e0 /* (26, 18, 17) */,
  32'h3eacaf9b /* (22, 18, 17) */,
  32'h3f19a2a7 /* (18, 18, 17) */,
  32'h3f19a2a7 /* (14, 18, 17) */,
  32'h3eacaf9b /* (10, 18, 17) */,
  32'h3e3e01e0 /* (6, 18, 17) */,
  32'h3e0adb0d /* (2, 18, 17) */,
  32'h3e0adb0d /* (30, 14, 17) */,
  32'h3e3e01e0 /* (26, 14, 17) */,
  32'h3eacaf9b /* (22, 14, 17) */,
  32'h3f19a2a7 /* (18, 14, 17) */,
  32'h3f19a2a7 /* (14, 14, 17) */,
  32'h3eacaf9b /* (10, 14, 17) */,
  32'h3e3e01e0 /* (6, 14, 17) */,
  32'h3e0adb0d /* (2, 14, 17) */,
  32'h3daa3ec9 /* (30, 10, 17) */,
  32'h3de44bb3 /* (26, 10, 17) */,
  32'h3e48eba4 /* (22, 10, 17) */,
  32'h3eacaf9b /* (18, 10, 17) */,
  32'h3eacaf9b /* (14, 10, 17) */,
  32'h3e48eba4 /* (10, 10, 17) */,
  32'h3de44bb3 /* (6, 10, 17) */,
  32'h3daa3ec9 /* (2, 10, 17) */,
  32'h3d4bfe66 /* (30, 6, 17) */,
  32'h3d85e8bf /* (26, 6, 17) */,
  32'h3de44bb3 /* (22, 6, 17) */,
  32'h3e3e01e0 /* (18, 6, 17) */,
  32'h3e3e01e0 /* (14, 6, 17) */,
  32'h3de44bb3 /* (10, 6, 17) */,
  32'h3d85e8bf /* (6, 6, 17) */,
  32'h3d4bfe66 /* (2, 6, 17) */,
  32'h3d1dadb9 /* (30, 2, 17) */,
  32'h3d4bfe66 /* (26, 2, 17) */,
  32'h3daa3ec9 /* (22, 2, 17) */,
  32'h3e0adb0d /* (18, 2, 17) */,
  32'h3e0adb0d /* (14, 2, 17) */,
  32'h3daa3ec9 /* (10, 2, 17) */,
  32'h3d4bfe66 /* (6, 2, 17) */,
  32'h3d1dadb9 /* (2, 2, 17) */,
  32'h3d246fbd /* (30, 30, 13) */,
  32'h3d4ce87b /* (26, 30, 13) */,
  32'h3da2895a /* (22, 30, 13) */,
  32'h3dfd653f /* (18, 30, 13) */,
  32'h3dfd653f /* (14, 30, 13) */,
  32'h3da2895a /* (10, 30, 13) */,
  32'h3d4ce87b /* (6, 30, 13) */,
  32'h3d246fbd /* (2, 30, 13) */,
  32'h3d4ce87b /* (30, 26, 13) */,
  32'h3d82bc35 /* (26, 26, 13) */,
  32'h3dd610ea /* (22, 26, 13) */,
  32'h3e2b8c37 /* (18, 26, 13) */,
  32'h3e2b8c37 /* (14, 26, 13) */,
  32'h3dd610ea /* (10, 26, 13) */,
  32'h3d82bc35 /* (6, 26, 13) */,
  32'h3d4ce87b /* (2, 26, 13) */,
  32'h3da2895a /* (30, 22, 13) */,
  32'h3dd610ea /* (26, 22, 13) */,
  32'h3e37540b /* (22, 22, 13) */,
  32'h3e994798 /* (18, 22, 13) */,
  32'h3e994798 /* (14, 22, 13) */,
  32'h3e37540b /* (10, 22, 13) */,
  32'h3dd610ea /* (6, 22, 13) */,
  32'h3da2895a /* (2, 22, 13) */,
  32'h3dfd653f /* (30, 18, 13) */,
  32'h3e2b8c37 /* (26, 18, 13) */,
  32'h3e994798 /* (22, 18, 13) */,
  32'h3f05dc96 /* (18, 18, 13) */,
  32'h3f05dc96 /* (14, 18, 13) */,
  32'h3e994798 /* (10, 18, 13) */,
  32'h3e2b8c37 /* (6, 18, 13) */,
  32'h3dfd653f /* (2, 18, 13) */,
  32'h3dfd653f /* (30, 14, 13) */,
  32'h3e2b8c37 /* (26, 14, 13) */,
  32'h3e994798 /* (22, 14, 13) */,
  32'h3f05dc96 /* (18, 14, 13) */,
  32'h3f05dc96 /* (14, 14, 13) */,
  32'h3e994798 /* (10, 14, 13) */,
  32'h3e2b8c37 /* (6, 14, 13) */,
  32'h3dfd653f /* (2, 14, 13) */,
  32'h3da2895a /* (30, 10, 13) */,
  32'h3dd610ea /* (26, 10, 13) */,
  32'h3e37540b /* (22, 10, 13) */,
  32'h3e994798 /* (18, 10, 13) */,
  32'h3e994798 /* (14, 10, 13) */,
  32'h3e37540b /* (10, 10, 13) */,
  32'h3dd610ea /* (6, 10, 13) */,
  32'h3da2895a /* (2, 10, 13) */,
  32'h3d4ce87b /* (30, 6, 13) */,
  32'h3d82bc35 /* (26, 6, 13) */,
  32'h3dd610ea /* (22, 6, 13) */,
  32'h3e2b8c37 /* (18, 6, 13) */,
  32'h3e2b8c37 /* (14, 6, 13) */,
  32'h3dd610ea /* (10, 6, 13) */,
  32'h3d82bc35 /* (6, 6, 13) */,
  32'h3d4ce87b /* (2, 6, 13) */,
  32'h3d246fbd /* (30, 2, 13) */,
  32'h3d4ce87b /* (26, 2, 13) */,
  32'h3da2895a /* (22, 2, 13) */,
  32'h3dfd653f /* (18, 2, 13) */,
  32'h3dfd653f /* (14, 2, 13) */,
  32'h3da2895a /* (10, 2, 13) */,
  32'h3d4ce87b /* (6, 2, 13) */,
  32'h3d246fbd /* (2, 2, 13) */,
  32'h3d1214c5 /* (30, 30, 9) */,
  32'h3d1e19af /* (26, 30, 9) */,
  32'h3d56480e /* (22, 30, 9) */,
  32'h3d94a37c /* (18, 30, 9) */,
  32'h3d94a37c /* (14, 30, 9) */,
  32'h3d56480e /* (10, 30, 9) */,
  32'h3d1e19af /* (6, 30, 9) */,
  32'h3d1214c5 /* (2, 30, 9) */,
  32'h3d1e19af /* (30, 26, 9) */,
  32'h3d37f9d0 /* (26, 26, 9) */,
  32'h3d866682 /* (22, 26, 9) */,
  32'h3dc45939 /* (18, 26, 9) */,
  32'h3dc45939 /* (14, 26, 9) */,
  32'h3d866682 /* (10, 26, 9) */,
  32'h3d37f9d0 /* (6, 26, 9) */,
  32'h3d1e19af /* (2, 26, 9) */,
  32'h3d56480e /* (30, 22, 9) */,
  32'h3d866682 /* (26, 22, 9) */,
  32'h3dd7137d /* (22, 22, 9) */,
  32'h3e28e750 /* (18, 22, 9) */,
  32'h3e28e750 /* (14, 22, 9) */,
  32'h3dd7137d /* (10, 22, 9) */,
  32'h3d866682 /* (6, 22, 9) */,
  32'h3d56480e /* (2, 22, 9) */,
  32'h3d94a37c /* (30, 18, 9) */,
  32'h3dc45939 /* (26, 18, 9) */,
  32'h3e28e750 /* (22, 18, 9) */,
  32'h3e8dd733 /* (18, 18, 9) */,
  32'h3e8dd733 /* (14, 18, 9) */,
  32'h3e28e750 /* (10, 18, 9) */,
  32'h3dc45939 /* (6, 18, 9) */,
  32'h3d94a37c /* (2, 18, 9) */,
  32'h3d94a37c /* (30, 14, 9) */,
  32'h3dc45939 /* (26, 14, 9) */,
  32'h3e28e750 /* (22, 14, 9) */,
  32'h3e8dd733 /* (18, 14, 9) */,
  32'h3e8dd733 /* (14, 14, 9) */,
  32'h3e28e750 /* (10, 14, 9) */,
  32'h3dc45939 /* (6, 14, 9) */,
  32'h3d94a37c /* (2, 14, 9) */,
  32'h3d56480e /* (30, 10, 9) */,
  32'h3d866682 /* (26, 10, 9) */,
  32'h3dd7137d /* (22, 10, 9) */,
  32'h3e28e750 /* (18, 10, 9) */,
  32'h3e28e750 /* (14, 10, 9) */,
  32'h3dd7137d /* (10, 10, 9) */,
  32'h3d866682 /* (6, 10, 9) */,
  32'h3d56480e /* (2, 10, 9) */,
  32'h3d1e19af /* (30, 6, 9) */,
  32'h3d37f9d0 /* (26, 6, 9) */,
  32'h3d866682 /* (22, 6, 9) */,
  32'h3dc45939 /* (18, 6, 9) */,
  32'h3dc45939 /* (14, 6, 9) */,
  32'h3d866682 /* (10, 6, 9) */,
  32'h3d37f9d0 /* (6, 6, 9) */,
  32'h3d1e19af /* (2, 6, 9) */,
  32'h3d1214c5 /* (30, 2, 9) */,
  32'h3d1e19af /* (26, 2, 9) */,
  32'h3d56480e /* (22, 2, 9) */,
  32'h3d94a37c /* (18, 2, 9) */,
  32'h3d94a37c /* (14, 2, 9) */,
  32'h3d56480e /* (10, 2, 9) */,
  32'h3d1e19af /* (6, 2, 9) */,
  32'h3d1214c5 /* (2, 2, 9) */,
  32'h3d4ca49b /* (30, 30, 5) */,
  32'h3d18df8d /* (26, 30, 5) */,
  32'h3d1f9f49 /* (22, 30, 5) */,
  32'h3d40d8bf /* (18, 30, 5) */,
  32'h3d40d8bf /* (14, 30, 5) */,
  32'h3d1f9f49 /* (10, 30, 5) */,
  32'h3d18df8d /* (6, 30, 5) */,
  32'h3d4ca49b /* (2, 30, 5) */,
  32'h3d18df8d /* (30, 26, 5) */,
  32'h3d16bb8b /* (26, 26, 5) */,
  32'h3d3c300c /* (22, 26, 5) */,
  32'h3d786cd6 /* (18, 26, 5) */,
  32'h3d786cd6 /* (14, 26, 5) */,
  32'h3d3c300c /* (10, 26, 5) */,
  32'h3d16bb8b /* (6, 26, 5) */,
  32'h3d18df8d /* (2, 26, 5) */,
  32'h3d1f9f49 /* (30, 22, 5) */,
  32'h3d3c300c /* (26, 22, 5) */,
  32'h3d8b85a2 /* (22, 22, 5) */,
  32'h3dce13fe /* (18, 22, 5) */,
  32'h3dce13fe /* (14, 22, 5) */,
  32'h3d8b85a2 /* (10, 22, 5) */,
  32'h3d3c300c /* (6, 22, 5) */,
  32'h3d1f9f49 /* (2, 22, 5) */,
  32'h3d40d8bf /* (30, 18, 5) */,
  32'h3d786cd6 /* (26, 18, 5) */,
  32'h3dce13fe /* (22, 18, 5) */,
  32'h3e27240a /* (18, 18, 5) */,
  32'h3e27240a /* (14, 18, 5) */,
  32'h3dce13fe /* (10, 18, 5) */,
  32'h3d786cd6 /* (6, 18, 5) */,
  32'h3d40d8bf /* (2, 18, 5) */,
  32'h3d40d8bf /* (30, 14, 5) */,
  32'h3d786cd6 /* (26, 14, 5) */,
  32'h3dce13fe /* (22, 14, 5) */,
  32'h3e27240a /* (18, 14, 5) */,
  32'h3e27240a /* (14, 14, 5) */,
  32'h3dce13fe /* (10, 14, 5) */,
  32'h3d786cd6 /* (6, 14, 5) */,
  32'h3d40d8bf /* (2, 14, 5) */,
  32'h3d1f9f49 /* (30, 10, 5) */,
  32'h3d3c300c /* (26, 10, 5) */,
  32'h3d8b85a2 /* (22, 10, 5) */,
  32'h3dce13fe /* (18, 10, 5) */,
  32'h3dce13fe /* (14, 10, 5) */,
  32'h3d8b85a2 /* (10, 10, 5) */,
  32'h3d3c300c /* (6, 10, 5) */,
  32'h3d1f9f49 /* (2, 10, 5) */,
  32'h3d18df8d /* (30, 6, 5) */,
  32'h3d16bb8b /* (26, 6, 5) */,
  32'h3d3c300c /* (22, 6, 5) */,
  32'h3d786cd6 /* (18, 6, 5) */,
  32'h3d786cd6 /* (14, 6, 5) */,
  32'h3d3c300c /* (10, 6, 5) */,
  32'h3d16bb8b /* (6, 6, 5) */,
  32'h3d18df8d /* (2, 6, 5) */,
  32'h3d4ca49b /* (30, 2, 5) */,
  32'h3d18df8d /* (26, 2, 5) */,
  32'h3d1f9f49 /* (22, 2, 5) */,
  32'h3d40d8bf /* (18, 2, 5) */,
  32'h3d40d8bf /* (14, 2, 5) */,
  32'h3d1f9f49 /* (10, 2, 5) */,
  32'h3d18df8d /* (6, 2, 5) */,
  32'h3d4ca49b /* (2, 2, 5) */,
  32'h3e0c4d23 /* (30, 30, 1) */,
  32'h3d3543e4 /* (26, 30, 1) */,
  32'h3d12ac07 /* (22, 30, 1) */,
  32'h3d217487 /* (18, 30, 1) */,
  32'h3d217487 /* (14, 30, 1) */,
  32'h3d12ac07 /* (10, 30, 1) */,
  32'h3d3543e4 /* (6, 30, 1) */,
  32'h3e0c4d23 /* (2, 30, 1) */,
  32'h3d3543e4 /* (30, 26, 1) */,
  32'h3d15cc97 /* (26, 26, 1) */,
  32'h3d2567ce /* (22, 26, 1) */,
  32'h3d4cf093 /* (18, 26, 1) */,
  32'h3d4cf093 /* (14, 26, 1) */,
  32'h3d2567ce /* (10, 26, 1) */,
  32'h3d15cc97 /* (6, 26, 1) */,
  32'h3d3543e4 /* (2, 26, 1) */,
  32'h3d12ac07 /* (30, 22, 1) */,
  32'h3d2567ce /* (26, 22, 1) */,
  32'h3d699f13 /* (22, 22, 1) */,
  32'h3da6958f /* (18, 22, 1) */,
  32'h3da6958f /* (14, 22, 1) */,
  32'h3d699f13 /* (10, 22, 1) */,
  32'h3d2567ce /* (6, 22, 1) */,
  32'h3d12ac07 /* (2, 22, 1) */,
  32'h3d217487 /* (30, 18, 1) */,
  32'h3d4cf093 /* (26, 18, 1) */,
  32'h3da6958f /* (22, 18, 1) */,
  32'h3e04a438 /* (18, 18, 1) */,
  32'h3e04a438 /* (14, 18, 1) */,
  32'h3da6958f /* (10, 18, 1) */,
  32'h3d4cf093 /* (6, 18, 1) */,
  32'h3d217487 /* (2, 18, 1) */,
  32'h3d217487 /* (30, 14, 1) */,
  32'h3d4cf093 /* (26, 14, 1) */,
  32'h3da6958f /* (22, 14, 1) */,
  32'h3e04a438 /* (18, 14, 1) */,
  32'h3e04a438 /* (14, 14, 1) */,
  32'h3da6958f /* (10, 14, 1) */,
  32'h3d4cf093 /* (6, 14, 1) */,
  32'h3d217487 /* (2, 14, 1) */,
  32'h3d12ac07 /* (30, 10, 1) */,
  32'h3d2567ce /* (26, 10, 1) */,
  32'h3d699f13 /* (22, 10, 1) */,
  32'h3da6958f /* (18, 10, 1) */,
  32'h3da6958f /* (14, 10, 1) */,
  32'h3d699f13 /* (10, 10, 1) */,
  32'h3d2567ce /* (6, 10, 1) */,
  32'h3d12ac07 /* (2, 10, 1) */,
  32'h3d3543e4 /* (30, 6, 1) */,
  32'h3d15cc97 /* (26, 6, 1) */,
  32'h3d2567ce /* (22, 6, 1) */,
  32'h3d4cf093 /* (18, 6, 1) */,
  32'h3d4cf093 /* (14, 6, 1) */,
  32'h3d2567ce /* (10, 6, 1) */,
  32'h3d15cc97 /* (6, 6, 1) */,
  32'h3d3543e4 /* (2, 6, 1) */,
  32'h3e0c4d23 /* (30, 2, 1) */,
  32'h3d3543e4 /* (26, 2, 1) */,
  32'h3d12ac07 /* (22, 2, 1) */,
  32'h3d217487 /* (18, 2, 1) */,
  32'h3d217487 /* (14, 2, 1) */,
  32'h3d12ac07 /* (10, 2, 1) */,
  32'h3d3543e4 /* (6, 2, 1) */,
  32'h3e0c4d23 /* (2, 2, 1) */,
  32'h3d866355 /* (29, 30, 29) */,
  32'h3d1a2949 /* (25, 30, 29) */,
  32'h3d1c5f03 /* (21, 30, 29) */,
  32'h3d240321 /* (17, 30, 29) */,
  32'h3d29e985 /* (13, 30, 29) */,
  32'h3d12f42a /* (9, 30, 29) */,
  32'h3d3cd255 /* (5, 30, 29) */,
  32'h3dbfa8df /* (1, 30, 29) */,
  32'h3d211f1b /* (29, 26, 29) */,
  32'h3d159d44 /* (25, 26, 29) */,
  32'h3d39bb76 /* (21, 26, 29) */,
  32'h3d54ba37 /* (17, 26, 29) */,
  32'h3d54a03b /* (13, 26, 29) */,
  32'h3d215063 /* (9, 26, 29) */,
  32'h3d16d305 /* (5, 26, 29) */,
  32'h3d2ba889 /* (1, 26, 29) */,
  32'h3d18cb02 /* (29, 22, 29) */,
  32'h3d387393 /* (25, 22, 29) */,
  32'h3d8ae43c /* (21, 22, 29) */,
  32'h3db22d06 /* (17, 22, 29) */,
  32'h3da99659 /* (13, 22, 29) */,
  32'h3d5dae2c /* (9, 22, 29) */,
  32'h3d2344c4 /* (5, 22, 29) */,
  32'h3d14c0fd /* (1, 22, 29) */,
  32'h3d3188e3 /* (29, 18, 29) */,
  32'h3d71c736 /* (25, 18, 29) */,
  32'h3dce7d45 /* (21, 18, 29) */,
  32'h3e11d12f /* (17, 18, 29) */,
  32'h3e04d0b8 /* (13, 18, 29) */,
  32'h3d9b2a7b /* (9, 18, 29) */,
  32'h3d487174 /* (5, 18, 29) */,
  32'h3d276174 /* (1, 18, 29) */,
  32'h3d3188e3 /* (29, 14, 29) */,
  32'h3d71c736 /* (25, 14, 29) */,
  32'h3dce7d45 /* (21, 14, 29) */,
  32'h3e11d12f /* (17, 14, 29) */,
  32'h3e04d0b8 /* (13, 14, 29) */,
  32'h3d9b2a7b /* (9, 14, 29) */,
  32'h3d487174 /* (5, 14, 29) */,
  32'h3d276174 /* (1, 14, 29) */,
  32'h3d18cb02 /* (29, 10, 29) */,
  32'h3d387393 /* (25, 10, 29) */,
  32'h3d8ae43c /* (21, 10, 29) */,
  32'h3db22d06 /* (17, 10, 29) */,
  32'h3da99659 /* (13, 10, 29) */,
  32'h3d5dae2c /* (9, 10, 29) */,
  32'h3d2344c4 /* (5, 10, 29) */,
  32'h3d14c0fd /* (1, 10, 29) */,
  32'h3d211f1b /* (29, 6, 29) */,
  32'h3d159d44 /* (25, 6, 29) */,
  32'h3d39bb76 /* (21, 6, 29) */,
  32'h3d54ba37 /* (17, 6, 29) */,
  32'h3d54a03b /* (13, 6, 29) */,
  32'h3d215063 /* (9, 6, 29) */,
  32'h3d16d305 /* (5, 6, 29) */,
  32'h3d2ba889 /* (1, 6, 29) */,
  32'h3d866355 /* (29, 2, 29) */,
  32'h3d1a2949 /* (25, 2, 29) */,
  32'h3d1c5f03 /* (21, 2, 29) */,
  32'h3d240321 /* (17, 2, 29) */,
  32'h3d29e985 /* (13, 2, 29) */,
  32'h3d12f42a /* (9, 2, 29) */,
  32'h3d3cd255 /* (5, 2, 29) */,
  32'h3dbfa8df /* (1, 2, 29) */,
  32'h3d1a2949 /* (29, 30, 25) */,
  32'h3d1777c7 /* (25, 30, 25) */,
  32'h3d42a7b8 /* (21, 30, 25) */,
  32'h3d62f778 /* (17, 30, 25) */,
  32'h3d6129ae /* (13, 30, 25) */,
  32'h3d26a1b5 /* (9, 30, 25) */,
  32'h3d14b1c0 /* (5, 30, 25) */,
  32'h3d20a35e /* (1, 30, 25) */,
  32'h3d159d44 /* (29, 26, 25) */,
  32'h3d29a602 /* (25, 26, 25) */,
  32'h3d71ecf9 /* (21, 26, 25) */,
  32'h3d95be73 /* (17, 26, 25) */,
  32'h3d90c8a7 /* (13, 26, 25) */,
  32'h3d45eb5b /* (9, 26, 25) */,
  32'h3d1b2471 /* (5, 26, 25) */,
  32'h3d146a43 /* (1, 26, 25) */,
  32'h3d387393 /* (29, 22, 25) */,
  32'h3d6deb12 /* (25, 22, 25) */,
  32'h3dbf3f1d /* (21, 22, 25) */,
  32'h3e009a19 /* (17, 22, 25) */,
  32'h3defa49b /* (13, 22, 25) */,
  32'h3d94014f /* (9, 22, 25) */,
  32'h3d4b3dc7 /* (5, 22, 25) */,
  32'h3d305430 /* (1, 22, 25) */,
  32'h3d71c736 /* (29, 18, 25) */,
  32'h3da8d240 /* (25, 18, 25) */,
  32'h3e14a5c9 /* (21, 18, 25) */,
  32'h3e57a44b /* (17, 18, 25) */,
  32'h3e41f14c /* (13, 18, 25) */,
  32'h3ddc09d8 /* (9, 18, 25) */,
  32'h3d8a0000 /* (5, 18, 25) */,
  32'h3d62906c /* (1, 18, 25) */,
  32'h3d71c736 /* (29, 14, 25) */,
  32'h3da8d240 /* (25, 14, 25) */,
  32'h3e14a5c9 /* (21, 14, 25) */,
  32'h3e57a44b /* (17, 14, 25) */,
  32'h3e41f14c /* (13, 14, 25) */,
  32'h3ddc09d8 /* (9, 14, 25) */,
  32'h3d8a0000 /* (5, 14, 25) */,
  32'h3d62906c /* (1, 14, 25) */,
  32'h3d387393 /* (29, 10, 25) */,
  32'h3d6deb12 /* (25, 10, 25) */,
  32'h3dbf3f1d /* (21, 10, 25) */,
  32'h3e009a19 /* (17, 10, 25) */,
  32'h3defa49b /* (13, 10, 25) */,
  32'h3d94014f /* (9, 10, 25) */,
  32'h3d4b3dc7 /* (5, 10, 25) */,
  32'h3d305430 /* (1, 10, 25) */,
  32'h3d159d44 /* (29, 6, 25) */,
  32'h3d29a602 /* (25, 6, 25) */,
  32'h3d71ecf9 /* (21, 6, 25) */,
  32'h3d95be73 /* (17, 6, 25) */,
  32'h3d90c8a7 /* (13, 6, 25) */,
  32'h3d45eb5b /* (9, 6, 25) */,
  32'h3d1b2471 /* (5, 6, 25) */,
  32'h3d146a43 /* (1, 6, 25) */,
  32'h3d1a2949 /* (29, 2, 25) */,
  32'h3d1777c7 /* (25, 2, 25) */,
  32'h3d42a7b8 /* (21, 2, 25) */,
  32'h3d62f778 /* (17, 2, 25) */,
  32'h3d6129ae /* (13, 2, 25) */,
  32'h3d26a1b5 /* (9, 2, 25) */,
  32'h3d14b1c0 /* (5, 2, 25) */,
  32'h3d20a35e /* (1, 2, 25) */,
  32'h3d1c5f03 /* (29, 30, 21) */,
  32'h3d42a7b8 /* (25, 30, 21) */,
  32'h3d96eb50 /* (21, 30, 21) */,
  32'h3dc59b81 /* (17, 30, 21) */,
  32'h3dba5db4 /* (13, 30, 21) */,
  32'h3d6d9fa3 /* (9, 30, 21) */,
  32'h3d29823f /* (5, 30, 21) */,
  32'h3d16ed42 /* (1, 30, 21) */,
  32'h3d39bb76 /* (29, 26, 21) */,
  32'h3d71ecf9 /* (25, 26, 21) */,
  32'h3dc480ba /* (21, 26, 21) */,
  32'h3e0533d0 /* (17, 26, 21) */,
  32'h3df74dbc /* (13, 26, 21) */,
  32'h3d9750ce /* (9, 26, 21) */,
  32'h3d4d9045 /* (5, 26, 21) */,
  32'h3d31191b /* (1, 26, 21) */,
  32'h3d8ae43c /* (29, 22, 21) */,
  32'h3dbf3f1d /* (25, 22, 21) */,
  32'h3e257fc6 /* (21, 22, 21) */,
  32'h3e6c6ac0 /* (17, 22, 21) */,
  32'h3e562fb1 /* (13, 22, 21) */,
  32'h3df71c69 /* (9, 22, 21) */,
  32'h3d9d9380 /* (5, 22, 21) */,
  32'h3d829849 /* (1, 22, 21) */,
  32'h3dce7d45 /* (29, 18, 21) */,
  32'h3e14a5c9 /* (25, 18, 21) */,
  32'h3e882756 /* (21, 18, 21) */,
  32'h3eccf8ff /* (17, 18, 21) */,
  32'h3eb517ce /* (13, 18, 21) */,
  32'h3e458f30 /* (9, 18, 21) */,
  32'h3deed79f /* (5, 18, 21) */,
  32'h3dc01db4 /* (1, 18, 21) */,
  32'h3dce7d45 /* (29, 14, 21) */,
  32'h3e14a5c9 /* (25, 14, 21) */,
  32'h3e882756 /* (21, 14, 21) */,
  32'h3eccf8ff /* (17, 14, 21) */,
  32'h3eb517ce /* (13, 14, 21) */,
  32'h3e458f30 /* (9, 14, 21) */,
  32'h3deed79f /* (5, 14, 21) */,
  32'h3dc01db4 /* (1, 14, 21) */,
  32'h3d8ae43c /* (29, 10, 21) */,
  32'h3dbf3f1d /* (25, 10, 21) */,
  32'h3e257fc6 /* (21, 10, 21) */,
  32'h3e6c6ac0 /* (17, 10, 21) */,
  32'h3e562fb1 /* (13, 10, 21) */,
  32'h3df71c69 /* (9, 10, 21) */,
  32'h3d9d9380 /* (5, 10, 21) */,
  32'h3d829849 /* (1, 10, 21) */,
  32'h3d39bb76 /* (29, 6, 21) */,
  32'h3d71ecf9 /* (25, 6, 21) */,
  32'h3dc480ba /* (21, 6, 21) */,
  32'h3e0533d0 /* (17, 6, 21) */,
  32'h3df74dbc /* (13, 6, 21) */,
  32'h3d9750ce /* (9, 6, 21) */,
  32'h3d4d9045 /* (5, 6, 21) */,
  32'h3d31191b /* (1, 6, 21) */,
  32'h3d1c5f03 /* (29, 2, 21) */,
  32'h3d42a7b8 /* (25, 2, 21) */,
  32'h3d96eb50 /* (21, 2, 21) */,
  32'h3dc59b81 /* (17, 2, 21) */,
  32'h3dba5db4 /* (13, 2, 21) */,
  32'h3d6d9fa3 /* (9, 2, 21) */,
  32'h3d29823f /* (5, 2, 21) */,
  32'h3d16ed42 /* (1, 2, 21) */,
  32'h3d240321 /* (29, 30, 17) */,
  32'h3d62f778 /* (25, 30, 17) */,
  32'h3dc59b81 /* (21, 30, 17) */,
  32'h3e0de5f8 /* (17, 30, 17) */,
  32'h3e003b1e /* (13, 30, 17) */,
  32'h3d9314c2 /* (9, 30, 17) */,
  32'h3d3a7be5 /* (5, 30, 17) */,
  32'h3d1a0745 /* (1, 30, 17) */,
  32'h3d54ba37 /* (29, 26, 17) */,
  32'h3d95be73 /* (25, 26, 17) */,
  32'h3e0533d0 /* (21, 26, 17) */,
  32'h3e430b11 /* (17, 26, 17) */,
  32'h3e2ea39a /* (13, 26, 17) */,
  32'h3dc42ad0 /* (9, 26, 17) */,
  32'h3d73b16f /* (5, 26, 17) */,
  32'h3d46f53f /* (1, 26, 17) */,
  32'h3db22d06 /* (29, 22, 17) */,
  32'h3e009a19 /* (25, 22, 17) */,
  32'h3e6c6ac0 /* (21, 22, 17) */,
  32'h3eb2925b /* (17, 22, 17) */,
  32'h3e9d80fb /* (13, 22, 17) */,
  32'h3e2b3653 /* (9, 22, 17) */,
  32'h3dce52e6 /* (5, 22, 17) */,
  32'h3da5ac70 /* (1, 22, 17) */,
  32'h3e11d12f /* (29, 18, 17) */,
  32'h3e57a44b /* (25, 18, 17) */,
  32'h3eccf8ff /* (21, 18, 17) */,
  32'h3f202f9a /* (17, 18, 17) */,
  32'h3f0af24f /* (13, 18, 17) */,
  32'h3e91e4f8 /* (9, 18, 17) */,
  32'h3e2a981c /* (5, 18, 17) */,
  32'h3e06d8bb /* (1, 18, 17) */,
  32'h3e11d12f /* (29, 14, 17) */,
  32'h3e57a44b /* (25, 14, 17) */,
  32'h3eccf8ff /* (21, 14, 17) */,
  32'h3f202f9a /* (17, 14, 17) */,
  32'h3f0af24f /* (13, 14, 17) */,
  32'h3e91e4f8 /* (9, 14, 17) */,
  32'h3e2a981c /* (5, 14, 17) */,
  32'h3e06d8bb /* (1, 14, 17) */,
  32'h3db22d06 /* (29, 10, 17) */,
  32'h3e009a19 /* (25, 10, 17) */,
  32'h3e6c6ac0 /* (21, 10, 17) */,
  32'h3eb2925b /* (17, 10, 17) */,
  32'h3e9d80fb /* (13, 10, 17) */,
  32'h3e2b3653 /* (9, 10, 17) */,
  32'h3dce52e6 /* (5, 10, 17) */,
  32'h3da5ac70 /* (1, 10, 17) */,
  32'h3d54ba37 /* (29, 6, 17) */,
  32'h3d95be73 /* (25, 6, 17) */,
  32'h3e0533d0 /* (21, 6, 17) */,
  32'h3e430b11 /* (17, 6, 17) */,
  32'h3e2ea39a /* (13, 6, 17) */,
  32'h3dc42ad0 /* (9, 6, 17) */,
  32'h3d73b16f /* (5, 6, 17) */,
  32'h3d46f53f /* (1, 6, 17) */,
  32'h3d240321 /* (29, 2, 17) */,
  32'h3d62f778 /* (25, 2, 17) */,
  32'h3dc59b81 /* (21, 2, 17) */,
  32'h3e0de5f8 /* (17, 2, 17) */,
  32'h3e003b1e /* (13, 2, 17) */,
  32'h3d9314c2 /* (9, 2, 17) */,
  32'h3d3a7be5 /* (5, 2, 17) */,
  32'h3d1a0745 /* (1, 2, 17) */,
  32'h3d29e985 /* (29, 30, 13) */,
  32'h3d6129ae /* (25, 30, 13) */,
  32'h3dba5db4 /* (21, 30, 13) */,
  32'h3e003b1e /* (17, 30, 13) */,
  32'h3dec70da /* (13, 30, 13) */,
  32'h3d8e358b /* (9, 30, 13) */,
  32'h3d3d84de /* (5, 30, 13) */,
  32'h3d214ba3 /* (1, 30, 13) */,
  32'h3d54a03b /* (29, 26, 13) */,
  32'h3d90c8a7 /* (25, 26, 13) */,
  32'h3df74dbc /* (21, 26, 13) */,
  32'h3e2ea39a /* (17, 26, 13) */,
  32'h3e1f113d /* (13, 26, 13) */,
  32'h3db9d5f4 /* (9, 26, 13) */,
  32'h3d700ffa /* (5, 26, 13) */,
  32'h3d4876ff /* (1, 26, 13) */,
  32'h3da99659 /* (29, 22, 13) */,
  32'h3defa49b /* (25, 22, 13) */,
  32'h3e562fb1 /* (21, 22, 13) */,
  32'h3e9d80fb /* (17, 22, 13) */,
  32'h3e8cbae1 /* (13, 22, 13) */,
  32'h3e1d56b2 /* (9, 22, 13) */,
  32'h3dc29629 /* (5, 22, 13) */,
  32'h3d9e7894 /* (1, 22, 13) */,
  32'h3e04d0b8 /* (29, 18, 13) */,
  32'h3e41f14c /* (25, 18, 13) */,
  32'h3eb517ce /* (21, 18, 13) */,
  32'h3f0af24f /* (17, 18, 13) */,
  32'h3ef33ce4 /* (13, 18, 13) */,
  32'h3e821787 /* (9, 18, 13) */,
  32'h3e1a8d8c /* (5, 18, 13) */,
  32'h3df65860 /* (1, 18, 13) */,
  32'h3e04d0b8 /* (29, 14, 13) */,
  32'h3e41f14c /* (25, 14, 13) */,
  32'h3eb517ce /* (21, 14, 13) */,
  32'h3f0af24f /* (17, 14, 13) */,
  32'h3ef33ce4 /* (13, 14, 13) */,
  32'h3e821787 /* (9, 14, 13) */,
  32'h3e1a8d8c /* (5, 14, 13) */,
  32'h3df65860 /* (1, 14, 13) */,
  32'h3da99659 /* (29, 10, 13) */,
  32'h3defa49b /* (25, 10, 13) */,
  32'h3e562fb1 /* (21, 10, 13) */,
  32'h3e9d80fb /* (17, 10, 13) */,
  32'h3e8cbae1 /* (13, 10, 13) */,
  32'h3e1d56b2 /* (9, 10, 13) */,
  32'h3dc29629 /* (5, 10, 13) */,
  32'h3d9e7894 /* (1, 10, 13) */,
  32'h3d54a03b /* (29, 6, 13) */,
  32'h3d90c8a7 /* (25, 6, 13) */,
  32'h3df74dbc /* (21, 6, 13) */,
  32'h3e2ea39a /* (17, 6, 13) */,
  32'h3e1f113d /* (13, 6, 13) */,
  32'h3db9d5f4 /* (9, 6, 13) */,
  32'h3d700ffa /* (5, 6, 13) */,
  32'h3d4876ff /* (1, 6, 13) */,
  32'h3d29e985 /* (29, 2, 13) */,
  32'h3d6129ae /* (25, 2, 13) */,
  32'h3dba5db4 /* (21, 2, 13) */,
  32'h3e003b1e /* (17, 2, 13) */,
  32'h3dec70da /* (13, 2, 13) */,
  32'h3d8e358b /* (9, 2, 13) */,
  32'h3d3d84de /* (5, 2, 13) */,
  32'h3d214ba3 /* (1, 2, 13) */,
  32'h3d12f42a /* (29, 30, 9) */,
  32'h3d26a1b5 /* (25, 30, 9) */,
  32'h3d6d9fa3 /* (21, 30, 9) */,
  32'h3d9314c2 /* (17, 30, 9) */,
  32'h3d8e358b /* (13, 30, 9) */,
  32'h3d42665b /* (9, 30, 9) */,
  32'h3d18622e /* (5, 30, 9) */,
  32'h3d11c69f /* (1, 30, 9) */,
  32'h3d215063 /* (29, 26, 9) */,
  32'h3d45eb5b /* (25, 26, 9) */,
  32'h3d9750ce /* (21, 26, 9) */,
  32'h3dc42ad0 /* (17, 26, 9) */,
  32'h3db9d5f4 /* (13, 26, 9) */,
  32'h3d6fd024 /* (9, 26, 9) */,
  32'h3d2db0cc /* (5, 26, 9) */,
  32'h3d1c53e8 /* (1, 26, 9) */,
  32'h3d5dae2c /* (29, 22, 9) */,
  32'h3d94014f /* (25, 22, 9) */,
  32'h3df71c69 /* (21, 22, 9) */,
  32'h3e2b3653 /* (17, 22, 9) */,
  32'h3e1d56b2 /* (13, 22, 9) */,
  32'h3dbbc730 /* (9, 22, 9) */,
  32'h3d781ae6 /* (5, 22, 9) */,
  32'h3d52081f /* (1, 22, 9) */,
  32'h3d9b2a7b /* (29, 18, 9) */,
  32'h3ddc09d8 /* (25, 18, 9) */,
  32'h3e458f30 /* (21, 18, 9) */,
  32'h3e91e4f8 /* (17, 18, 9) */,
  32'h3e821787 /* (13, 18, 9) */,
  32'h3e10cac5 /* (9, 18, 9) */,
  32'h3db24f8e /* (5, 18, 9) */,
  32'h3d90dff9 /* (1, 18, 9) */,
  32'h3d9b2a7b /* (29, 14, 9) */,
  32'h3ddc09d8 /* (25, 14, 9) */,
  32'h3e458f30 /* (21, 14, 9) */,
  32'h3e91e4f8 /* (17, 14, 9) */,
  32'h3e821787 /* (13, 14, 9) */,
  32'h3e10cac5 /* (9, 14, 9) */,
  32'h3db24f8e /* (5, 14, 9) */,
  32'h3d90dff9 /* (1, 14, 9) */,
  32'h3d5dae2c /* (29, 10, 9) */,
  32'h3d94014f /* (25, 10, 9) */,
  32'h3df71c69 /* (21, 10, 9) */,
  32'h3e2b3653 /* (17, 10, 9) */,
  32'h3e1d56b2 /* (13, 10, 9) */,
  32'h3dbbc730 /* (9, 10, 9) */,
  32'h3d781ae6 /* (5, 10, 9) */,
  32'h3d52081f /* (1, 10, 9) */,
  32'h3d215063 /* (29, 6, 9) */,
  32'h3d45eb5b /* (25, 6, 9) */,
  32'h3d9750ce /* (21, 6, 9) */,
  32'h3dc42ad0 /* (17, 6, 9) */,
  32'h3db9d5f4 /* (13, 6, 9) */,
  32'h3d6fd024 /* (9, 6, 9) */,
  32'h3d2db0cc /* (5, 6, 9) */,
  32'h3d1c53e8 /* (1, 6, 9) */,
  32'h3d12f42a /* (29, 2, 9) */,
  32'h3d26a1b5 /* (25, 2, 9) */,
  32'h3d6d9fa3 /* (21, 2, 9) */,
  32'h3d9314c2 /* (17, 2, 9) */,
  32'h3d8e358b /* (13, 2, 9) */,
  32'h3d42665b /* (9, 2, 9) */,
  32'h3d18622e /* (5, 2, 9) */,
  32'h3d11c69f /* (1, 2, 9) */,
  32'h3d3cd255 /* (29, 30, 5) */,
  32'h3d14b1c0 /* (25, 30, 5) */,
  32'h3d29823f /* (21, 30, 5) */,
  32'h3d3a7be5 /* (17, 30, 5) */,
  32'h3d3d84de /* (13, 30, 5) */,
  32'h3d18622e /* (9, 30, 5) */,
  32'h3d213c91 /* (5, 30, 5) */,
  32'h3d59109a /* (1, 30, 5) */,
  32'h3d16d305 /* (29, 26, 5) */,
  32'h3d1b2471 /* (25, 26, 5) */,
  32'h3d4d9045 /* (21, 26, 5) */,
  32'h3d73b16f /* (17, 26, 5) */,
  32'h3d700ffa /* (13, 26, 5) */,
  32'h3d2db0cc /* (9, 26, 5) */,
  32'h3d14f7ce /* (5, 26, 5) */,
  32'h3d1a8b5a /* (1, 26, 5) */,
  32'h3d2344c4 /* (29, 22, 5) */,
  32'h3d4b3dc7 /* (25, 22, 5) */,
  32'h3d9d9380 /* (21, 22, 5) */,
  32'h3dce52e6 /* (17, 22, 5) */,
  32'h3dc29629 /* (13, 22, 5) */,
  32'h3d781ae6 /* (9, 22, 5) */,
  32'h3d30fc5a /* (5, 22, 5) */,
  32'h3d1d9589 /* (1, 22, 5) */,
  32'h3d487174 /* (29, 18, 5) */,
  32'h3d8a0000 /* (25, 18, 5) */,
  32'h3deed79f /* (21, 18, 5) */,
  32'h3e2a981c /* (17, 18, 5) */,
  32'h3e1a8d8c /* (13, 18, 5) */,
  32'h3db24f8e /* (9, 18, 5) */,
  32'h3d63687e /* (5, 18, 5) */,
  32'h3d3c7841 /* (1, 18, 5) */,
  32'h3d487174 /* (29, 14, 5) */,
  32'h3d8a0000 /* (25, 14, 5) */,
  32'h3deed79f /* (21, 14, 5) */,
  32'h3e2a981c /* (17, 14, 5) */,
  32'h3e1a8d8c /* (13, 14, 5) */,
  32'h3db24f8e /* (9, 14, 5) */,
  32'h3d63687e /* (5, 14, 5) */,
  32'h3d3c7841 /* (1, 14, 5) */,
  32'h3d2344c4 /* (29, 10, 5) */,
  32'h3d4b3dc7 /* (25, 10, 5) */,
  32'h3d9d9380 /* (21, 10, 5) */,
  32'h3dce52e6 /* (17, 10, 5) */,
  32'h3dc29629 /* (13, 10, 5) */,
  32'h3d781ae6 /* (9, 10, 5) */,
  32'h3d30fc5a /* (5, 10, 5) */,
  32'h3d1d9589 /* (1, 10, 5) */,
  32'h3d16d305 /* (29, 6, 5) */,
  32'h3d1b2471 /* (25, 6, 5) */,
  32'h3d4d9045 /* (21, 6, 5) */,
  32'h3d73b16f /* (17, 6, 5) */,
  32'h3d700ffa /* (13, 6, 5) */,
  32'h3d2db0cc /* (9, 6, 5) */,
  32'h3d14f7ce /* (5, 6, 5) */,
  32'h3d1a8b5a /* (1, 6, 5) */,
  32'h3d3cd255 /* (29, 2, 5) */,
  32'h3d14b1c0 /* (25, 2, 5) */,
  32'h3d29823f /* (21, 2, 5) */,
  32'h3d3a7be5 /* (17, 2, 5) */,
  32'h3d3d84de /* (13, 2, 5) */,
  32'h3d18622e /* (9, 2, 5) */,
  32'h3d213c91 /* (5, 2, 5) */,
  32'h3d59109a /* (1, 2, 5) */,
  32'h3dbfa8df /* (29, 30, 1) */,
  32'h3d20a35e /* (25, 30, 1) */,
  32'h3d16ed42 /* (21, 30, 1) */,
  32'h3d1a0745 /* (17, 30, 1) */,
  32'h3d214ba3 /* (13, 30, 1) */,
  32'h3d11c69f /* (9, 30, 1) */,
  32'h3d59109a /* (5, 30, 1) */,
  32'h3e4aeee2 /* (1, 30, 1) */,
  32'h3d2ba889 /* (29, 26, 1) */,
  32'h3d146a43 /* (25, 26, 1) */,
  32'h3d31191b /* (21, 26, 1) */,
  32'h3d46f53f /* (17, 26, 1) */,
  32'h3d4876ff /* (13, 26, 1) */,
  32'h3d1c53e8 /* (9, 26, 1) */,
  32'h3d1a8b5a /* (5, 26, 1) */,
  32'h3d3c9698 /* (1, 26, 1) */,
  32'h3d14c0fd /* (29, 22, 1) */,
  32'h3d305430 /* (25, 22, 1) */,
  32'h3d829849 /* (21, 22, 1) */,
  32'h3da5ac70 /* (17, 22, 1) */,
  32'h3d9e7894 /* (13, 22, 1) */,
  32'h3d52081f /* (9, 22, 1) */,
  32'h3d1d9589 /* (5, 22, 1) */,
  32'h3d119771 /* (1, 22, 1) */,
  32'h3d276174 /* (29, 18, 1) */,
  32'h3d62906c /* (25, 18, 1) */,
  32'h3dc01db4 /* (21, 18, 1) */,
  32'h3e06d8bb /* (17, 18, 1) */,
  32'h3df65860 /* (13, 18, 1) */,
  32'h3d90dff9 /* (9, 18, 1) */,
  32'h3d3c7841 /* (5, 18, 1) */,
  32'h3d1e0bb6 /* (1, 18, 1) */,
  32'h3d276174 /* (29, 14, 1) */,
  32'h3d62906c /* (25, 14, 1) */,
  32'h3dc01db4 /* (21, 14, 1) */,
  32'h3e06d8bb /* (17, 14, 1) */,
  32'h3df65860 /* (13, 14, 1) */,
  32'h3d90dff9 /* (9, 14, 1) */,
  32'h3d3c7841 /* (5, 14, 1) */,
  32'h3d1e0bb6 /* (1, 14, 1) */,
  32'h3d14c0fd /* (29, 10, 1) */,
  32'h3d305430 /* (25, 10, 1) */,
  32'h3d829849 /* (21, 10, 1) */,
  32'h3da5ac70 /* (17, 10, 1) */,
  32'h3d9e7894 /* (13, 10, 1) */,
  32'h3d52081f /* (9, 10, 1) */,
  32'h3d1d9589 /* (5, 10, 1) */,
  32'h3d119771 /* (1, 10, 1) */,
  32'h3d2ba889 /* (29, 6, 1) */,
  32'h3d146a43 /* (25, 6, 1) */,
  32'h3d31191b /* (21, 6, 1) */,
  32'h3d46f53f /* (17, 6, 1) */,
  32'h3d4876ff /* (13, 6, 1) */,
  32'h3d1c53e8 /* (9, 6, 1) */,
  32'h3d1a8b5a /* (5, 6, 1) */,
  32'h3d3c9698 /* (1, 6, 1) */,
  32'h3dbfa8df /* (29, 2, 1) */,
  32'h3d20a35e /* (25, 2, 1) */,
  32'h3d16ed42 /* (21, 2, 1) */,
  32'h3d1a0745 /* (17, 2, 1) */,
  32'h3d214ba3 /* (13, 2, 1) */,
  32'h3d11c69f /* (9, 2, 1) */,
  32'h3d59109a /* (5, 2, 1) */,
  32'h3e4aeee2 /* (1, 2, 1) */,
  32'h3d5defd3 /* (28, 30, 29) */,
  32'h3d13e9f7 /* (24, 30, 29) */,
  32'h3d23d587 /* (20, 30, 29) */,
  32'h3d13661d /* (16, 30, 29) */,
  32'h3d23d587 /* (12, 30, 29) */,
  32'h3d13e9f7 /* (8, 30, 29) */,
  32'h3d5defd3 /* (4, 30, 29) */,
  32'h3dcbea25 /* (0, 30, 29) */,
  32'h3d1b3fff /* (28, 26, 29) */,
  32'h3d19bf4b /* (24, 26, 29) */,
  32'h3d48406d /* (20, 26, 29) */,
  32'h3d41d3ae /* (16, 26, 29) */,
  32'h3d48406d /* (12, 26, 29) */,
  32'h3d19bf4b /* (8, 26, 29) */,
  32'h3d1b3fff /* (4, 26, 29) */,
  32'h3d2d5b95 /* (0, 26, 29) */,
  32'h3d1cff11 /* (28, 22, 29) */,
  32'h3d48bc7e /* (24, 22, 29) */,
  32'h3d9aff71 /* (20, 22, 29) */,
  32'h3da59d10 /* (16, 22, 29) */,
  32'h3d9aff71 /* (12, 22, 29) */,
  32'h3d48bc7e /* (8, 22, 29) */,
  32'h3d1cff11 /* (4, 22, 29) */,
  32'h3d144f19 /* (0, 22, 29) */,
  32'h3d3b1e93 /* (28, 18, 29) */,
  32'h3d880501 /* (24, 18, 29) */,
  32'h3decc5e8 /* (20, 18, 29) */,
  32'h3e0a27e7 /* (16, 18, 29) */,
  32'h3decc5e8 /* (12, 18, 29) */,
  32'h3d880501 /* (8, 18, 29) */,
  32'h3d3b1e93 /* (4, 18, 29) */,
  32'h3d262b6e /* (0, 18, 29) */,
  32'h3d3b1e93 /* (28, 14, 29) */,
  32'h3d880501 /* (24, 14, 29) */,
  32'h3decc5e8 /* (20, 14, 29) */,
  32'h3e0a27e7 /* (16, 14, 29) */,
  32'h3decc5e8 /* (12, 14, 29) */,
  32'h3d880501 /* (8, 14, 29) */,
  32'h3d3b1e93 /* (4, 14, 29) */,
  32'h3d262b6e /* (0, 14, 29) */,
  32'h3d1cff11 /* (28, 10, 29) */,
  32'h3d48bc7e /* (24, 10, 29) */,
  32'h3d9aff71 /* (20, 10, 29) */,
  32'h3da59d10 /* (16, 10, 29) */,
  32'h3d9aff71 /* (12, 10, 29) */,
  32'h3d48bc7e /* (8, 10, 29) */,
  32'h3d1cff11 /* (4, 10, 29) */,
  32'h3d144f19 /* (0, 10, 29) */,
  32'h3d1b3fff /* (28, 6, 29) */,
  32'h3d19bf4b /* (24, 6, 29) */,
  32'h3d48406d /* (20, 6, 29) */,
  32'h3d41d3ae /* (16, 6, 29) */,
  32'h3d48406d /* (12, 6, 29) */,
  32'h3d19bf4b /* (8, 6, 29) */,
  32'h3d1b3fff /* (4, 6, 29) */,
  32'h3d2d5b95 /* (0, 6, 29) */,
  32'h3d5defd3 /* (28, 2, 29) */,
  32'h3d13e9f7 /* (24, 2, 29) */,
  32'h3d23d587 /* (20, 2, 29) */,
  32'h3d13661d /* (16, 2, 29) */,
  32'h3d23d587 /* (12, 2, 29) */,
  32'h3d13e9f7 /* (8, 2, 29) */,
  32'h3d5defd3 /* (4, 2, 29) */,
  32'h3dcbea25 /* (0, 2, 29) */,
  32'h3d16c6a3 /* (28, 30, 25) */,
  32'h3d1d59b0 /* (24, 30, 25) */,
  32'h3d530d8e /* (20, 30, 25) */,
  32'h3d4f6a6e /* (16, 30, 25) */,
  32'h3d530d8e /* (12, 30, 25) */,
  32'h3d1d59b0 /* (8, 30, 25) */,
  32'h3d16c6a3 /* (4, 30, 25) */,
  32'h3d21b235 /* (0, 30, 25) */,
  32'h3d17902e /* (28, 26, 25) */,
  32'h3d35cd98 /* (24, 26, 25) */,
  32'h3d859348 /* (20, 26, 25) */,
  32'h3d8a46e7 /* (16, 26, 25) */,
  32'h3d859348 /* (12, 26, 25) */,
  32'h3d35cd98 /* (8, 26, 25) */,
  32'h3d17902e /* (4, 26, 25) */,
  32'h3d1459dd /* (0, 26, 25) */,
  32'h3d404057 /* (28, 22, 25) */,
  32'h3d83c517 /* (24, 22, 25) */,
  32'h3dd85675 /* (20, 22, 25) */,
  32'h3df142da /* (16, 22, 25) */,
  32'h3dd85675 /* (12, 22, 25) */,
  32'h3d83c517 /* (8, 22, 25) */,
  32'h3d404057 /* (4, 22, 25) */,
  32'h3d2f5f5a /* (0, 22, 25) */,
  32'h3d800deb /* (28, 18, 25) */,
  32'h3dbf672f /* (24, 18, 25) */,
  32'h3e2baf50 /* (20, 18, 25) */,
  32'h3e4d7ce8 /* (16, 18, 25) */,
  32'h3e2baf50 /* (12, 18, 25) */,
  32'h3dbf672f /* (8, 18, 25) */,
  32'h3d800deb /* (4, 18, 25) */,
  32'h3d60bf24 /* (0, 18, 25) */,
  32'h3d800deb /* (28, 14, 25) */,
  32'h3dbf672f /* (24, 14, 25) */,
  32'h3e2baf50 /* (20, 14, 25) */,
  32'h3e4d7ce8 /* (16, 14, 25) */,
  32'h3e2baf50 /* (12, 14, 25) */,
  32'h3dbf672f /* (8, 14, 25) */,
  32'h3d800deb /* (4, 14, 25) */,
  32'h3d60bf24 /* (0, 14, 25) */,
  32'h3d404057 /* (28, 10, 25) */,
  32'h3d83c517 /* (24, 10, 25) */,
  32'h3dd85675 /* (20, 10, 25) */,
  32'h3df142da /* (16, 10, 25) */,
  32'h3dd85675 /* (12, 10, 25) */,
  32'h3d83c517 /* (8, 10, 25) */,
  32'h3d404057 /* (4, 10, 25) */,
  32'h3d2f5f5a /* (0, 10, 25) */,
  32'h3d17902e /* (28, 6, 25) */,
  32'h3d35cd98 /* (24, 6, 25) */,
  32'h3d859348 /* (20, 6, 25) */,
  32'h3d8a46e7 /* (16, 6, 25) */,
  32'h3d859348 /* (12, 6, 25) */,
  32'h3d35cd98 /* (8, 6, 25) */,
  32'h3d17902e /* (4, 6, 25) */,
  32'h3d1459dd /* (0, 6, 25) */,
  32'h3d16c6a3 /* (28, 2, 25) */,
  32'h3d1d59b0 /* (24, 2, 25) */,
  32'h3d530d8e /* (20, 2, 25) */,
  32'h3d4f6a6e /* (16, 2, 25) */,
  32'h3d530d8e /* (12, 2, 25) */,
  32'h3d1d59b0 /* (8, 2, 25) */,
  32'h3d16c6a3 /* (4, 2, 25) */,
  32'h3d21b235 /* (0, 2, 25) */,
  32'h3d21c128 /* (28, 30, 21) */,
  32'h3d558b1c /* (24, 30, 21) */,
  32'h3da96c08 /* (20, 30, 21) */,
  32'h3db86416 /* (16, 30, 21) */,
  32'h3da96c08 /* (12, 30, 21) */,
  32'h3d558b1c /* (8, 30, 21) */,
  32'h3d21c128 /* (4, 30, 21) */,
  32'h3d164ce1 /* (0, 30, 21) */,
  32'h3d41fb9f /* (28, 26, 21) */,
  32'h3d865b59 /* (24, 26, 21) */,
  32'h3ddec971 /* (20, 26, 21) */,
  32'h3dfa4afe /* (16, 26, 21) */,
  32'h3ddec971 /* (12, 26, 21) */,
  32'h3d865b59 /* (8, 26, 21) */,
  32'h3d41fb9f /* (4, 26, 21) */,
  32'h3d3013e2 /* (0, 26, 21) */,
  32'h3d92b699 /* (28, 22, 21) */,
  32'h3dd7e578 /* (24, 22, 21) */,
  32'h3e3e5baf /* (20, 22, 21) */,
  32'h3e60898b /* (16, 22, 21) */,
  32'h3e3e5baf /* (12, 22, 21) */,
  32'h3dd7e578 /* (8, 22, 21) */,
  32'h3d92b699 /* (4, 22, 21) */,
  32'h3d819abc /* (0, 22, 21) */,
  32'h3ddc0819 /* (28, 18, 21) */,
  32'h3e2a27e4 /* (24, 18, 21) */,
  32'h3e9ecc49 /* (20, 18, 21) */,
  32'h3ec4f0a1 /* (16, 18, 21) */,
  32'h3e9ecc49 /* (12, 18, 21) */,
  32'h3e2a27e4 /* (8, 18, 21) */,
  32'h3ddc0819 /* (4, 18, 21) */,
  32'h3dbe661f /* (0, 18, 21) */,
  32'h3ddc0819 /* (28, 14, 21) */,
  32'h3e2a27e4 /* (24, 14, 21) */,
  32'h3e9ecc49 /* (20, 14, 21) */,
  32'h3ec4f0a1 /* (16, 14, 21) */,
  32'h3e9ecc49 /* (12, 14, 21) */,
  32'h3e2a27e4 /* (8, 14, 21) */,
  32'h3ddc0819 /* (4, 14, 21) */,
  32'h3dbe661f /* (0, 14, 21) */,
  32'h3d92b699 /* (28, 10, 21) */,
  32'h3dd7e578 /* (24, 10, 21) */,
  32'h3e3e5baf /* (20, 10, 21) */,
  32'h3e60898b /* (16, 10, 21) */,
  32'h3e3e5baf /* (12, 10, 21) */,
  32'h3dd7e578 /* (8, 10, 21) */,
  32'h3d92b699 /* (4, 10, 21) */,
  32'h3d819abc /* (0, 10, 21) */,
  32'h3d41fb9f /* (28, 6, 21) */,
  32'h3d865b59 /* (24, 6, 21) */,
  32'h3ddec971 /* (20, 6, 21) */,
  32'h3dfa4afe /* (16, 6, 21) */,
  32'h3ddec971 /* (12, 6, 21) */,
  32'h3d865b59 /* (8, 6, 21) */,
  32'h3d41fb9f /* (4, 6, 21) */,
  32'h3d3013e2 /* (0, 6, 21) */,
  32'h3d21c128 /* (28, 2, 21) */,
  32'h3d558b1c /* (24, 2, 21) */,
  32'h3da96c08 /* (20, 2, 21) */,
  32'h3db86416 /* (16, 2, 21) */,
  32'h3da96c08 /* (12, 2, 21) */,
  32'h3d558b1c /* (8, 2, 21) */,
  32'h3d21c128 /* (4, 2, 21) */,
  32'h3d164ce1 /* (0, 2, 21) */,
  32'h3d2d6bba /* (28, 30, 17) */,
  32'h3d804df8 /* (24, 30, 17) */,
  32'h3de39dff /* (20, 30, 17) */,
  32'h3e06ec2e /* (16, 30, 17) */,
  32'h3de39dff /* (12, 30, 17) */,
  32'h3d804df8 /* (8, 30, 17) */,
  32'h3d2d6bba /* (4, 30, 17) */,
  32'h3d18d610 /* (0, 30, 17) */,
  32'h3d61b1de /* (28, 26, 17) */,
  32'h3daa3349 /* (24, 26, 17) */,
  32'h3e1a3a56 /* (20, 26, 17) */,
  32'h3e3a3d1a /* (16, 26, 17) */,
  32'h3e1a3a56 /* (12, 26, 17) */,
  32'h3daa3349 /* (8, 26, 17) */,
  32'h3d61b1de /* (4, 26, 17) */,
  32'h3d455011 /* (0, 26, 17) */,
  32'h3dbdf4f8 /* (28, 22, 17) */,
  32'h3e135573 /* (24, 22, 17) */,
  32'h3e89fde5 /* (20, 22, 17) */,
  32'h3eabb572 /* (16, 22, 17) */,
  32'h3e89fde5 /* (12, 22, 17) */,
  32'h3e135573 /* (8, 22, 17) */,
  32'h3dbdf4f8 /* (4, 22, 17) */,
  32'h3da42e1b /* (0, 22, 17) */,
  32'h3e1c2ca1 /* (28, 18, 17) */,
  32'h3e79034c /* (24, 18, 17) */,
  32'h3ef15f91 /* (20, 18, 17) */,
  32'h3f1b42bd /* (16, 18, 17) */,
  32'h3ef15f91 /* (12, 18, 17) */,
  32'h3e79034c /* (8, 18, 17) */,
  32'h3e1c2ca1 /* (4, 18, 17) */,
  32'h3e05899d /* (0, 18, 17) */,
  32'h3e1c2ca1 /* (28, 14, 17) */,
  32'h3e79034c /* (24, 14, 17) */,
  32'h3ef15f91 /* (20, 14, 17) */,
  32'h3f1b42bd /* (16, 14, 17) */,
  32'h3ef15f91 /* (12, 14, 17) */,
  32'h3e79034c /* (8, 14, 17) */,
  32'h3e1c2ca1 /* (4, 14, 17) */,
  32'h3e05899d /* (0, 14, 17) */,
  32'h3dbdf4f8 /* (28, 10, 17) */,
  32'h3e135573 /* (24, 10, 17) */,
  32'h3e89fde5 /* (20, 10, 17) */,
  32'h3eabb572 /* (16, 10, 17) */,
  32'h3e89fde5 /* (12, 10, 17) */,
  32'h3e135573 /* (8, 10, 17) */,
  32'h3dbdf4f8 /* (4, 10, 17) */,
  32'h3da42e1b /* (0, 10, 17) */,
  32'h3d61b1de /* (28, 6, 17) */,
  32'h3daa3349 /* (24, 6, 17) */,
  32'h3e1a3a56 /* (20, 6, 17) */,
  32'h3e3a3d1a /* (16, 6, 17) */,
  32'h3e1a3a56 /* (12, 6, 17) */,
  32'h3daa3349 /* (8, 6, 17) */,
  32'h3d61b1de /* (4, 6, 17) */,
  32'h3d455011 /* (0, 6, 17) */,
  32'h3d2d6bba /* (28, 2, 17) */,
  32'h3d804df8 /* (24, 2, 17) */,
  32'h3de39dff /* (20, 2, 17) */,
  32'h3e06ec2e /* (16, 2, 17) */,
  32'h3de39dff /* (12, 2, 17) */,
  32'h3d804df8 /* (8, 2, 17) */,
  32'h3d2d6bba /* (4, 2, 17) */,
  32'h3d18d610 /* (0, 2, 17) */,
  32'h3d3217f4 /* (28, 30, 13) */,
  32'h3d7b52f8 /* (24, 30, 13) */,
  32'h3dd42d31 /* (20, 30, 13) */,
  32'h3df1ae3d /* (16, 30, 13) */,
  32'h3dd42d31 /* (12, 30, 13) */,
  32'h3d7b52f8 /* (8, 30, 13) */,
  32'h3d3217f4 /* (4, 30, 13) */,
  32'h3d2045b1 /* (0, 30, 13) */,
  32'h3d601ae9 /* (28, 26, 13) */,
  32'h3da2e7a9 /* (24, 26, 13) */,
  32'h3e0dc95f /* (20, 26, 13) */,
  32'h3e2576a9 /* (16, 26, 13) */,
  32'h3e0dc95f /* (12, 26, 13) */,
  32'h3da2e7a9 /* (8, 26, 13) */,
  32'h3d601ae9 /* (4, 26, 13) */,
  32'h3d4703b2 /* (0, 26, 13) */,
  32'h3db40e50 /* (28, 22, 13) */,
  32'h3e085939 /* (24, 22, 13) */,
  32'h3e7848b5 /* (20, 22, 13) */,
  32'h3e968a40 /* (16, 22, 13) */,
  32'h3e7848b5 /* (12, 22, 13) */,
  32'h3e085939 /* (8, 22, 13) */,
  32'h3db40e50 /* (4, 22, 13) */,
  32'h3d9d248b /* (0, 22, 13) */,
  32'h3e0de89e /* (28, 18, 13) */,
  32'h3e5f05ce /* (24, 18, 13) */,
  32'h3ed441df /* (20, 18, 13) */,
  32'h3f06176f /* (16, 18, 13) */,
  32'h3ed441df /* (12, 18, 13) */,
  32'h3e5f05ce /* (8, 18, 13) */,
  32'h3e0de89e /* (4, 18, 13) */,
  32'h3df40add /* (0, 18, 13) */,
  32'h3e0de89e /* (28, 14, 13) */,
  32'h3e5f05ce /* (24, 14, 13) */,
  32'h3ed441df /* (20, 14, 13) */,
  32'h3f06176f /* (16, 14, 13) */,
  32'h3ed441df /* (12, 14, 13) */,
  32'h3e5f05ce /* (8, 14, 13) */,
  32'h3e0de89e /* (4, 14, 13) */,
  32'h3df40add /* (0, 14, 13) */,
  32'h3db40e50 /* (28, 10, 13) */,
  32'h3e085939 /* (24, 10, 13) */,
  32'h3e7848b5 /* (20, 10, 13) */,
  32'h3e968a40 /* (16, 10, 13) */,
  32'h3e7848b5 /* (12, 10, 13) */,
  32'h3e085939 /* (8, 10, 13) */,
  32'h3db40e50 /* (4, 10, 13) */,
  32'h3d9d248b /* (0, 10, 13) */,
  32'h3d601ae9 /* (28, 6, 13) */,
  32'h3da2e7a9 /* (24, 6, 13) */,
  32'h3e0dc95f /* (20, 6, 13) */,
  32'h3e2576a9 /* (16, 6, 13) */,
  32'h3e0dc95f /* (12, 6, 13) */,
  32'h3da2e7a9 /* (8, 6, 13) */,
  32'h3d601ae9 /* (4, 6, 13) */,
  32'h3d4703b2 /* (0, 6, 13) */,
  32'h3d3217f4 /* (28, 2, 13) */,
  32'h3d7b52f8 /* (24, 2, 13) */,
  32'h3dd42d31 /* (20, 2, 13) */,
  32'h3df1ae3d /* (16, 2, 13) */,
  32'h3dd42d31 /* (12, 2, 13) */,
  32'h3d7b52f8 /* (8, 2, 13) */,
  32'h3d3217f4 /* (4, 2, 13) */,
  32'h3d2045b1 /* (0, 2, 13) */,
  32'h3d14de35 /* (28, 30, 9) */,
  32'h3d3291f6 /* (24, 30, 9) */,
  32'h3d833332 /* (20, 30, 9) */,
  32'h3d87d16b /* (16, 30, 9) */,
  32'h3d833332 /* (12, 30, 9) */,
  32'h3d3291f6 /* (8, 30, 9) */,
  32'h3d14de35 /* (4, 30, 9) */,
  32'h3d11b684 /* (0, 30, 9) */,
  32'h3d2657dd /* (28, 26, 9) */,
  32'h3d584c0c /* (24, 26, 9) */,
  32'h3da96159 /* (20, 26, 9) */,
  32'h3db6b309 /* (16, 26, 9) */,
  32'h3da96159 /* (12, 26, 9) */,
  32'h3d584c0c /* (8, 26, 9) */,
  32'h3d2657dd /* (4, 26, 9) */,
  32'h3d1bc36a /* (0, 26, 9) */,
  32'h3d68b7a2 /* (28, 22, 9) */,
  32'h3da590e9 /* (24, 22, 9) */,
  32'h3e0cf021 /* (20, 22, 9) */,
  32'h3e21930d /* (16, 22, 9) */,
  32'h3e0cf021 /* (12, 22, 9) */,
  32'h3da590e9 /* (8, 22, 9) */,
  32'h3d68b7a2 /* (4, 22, 9) */,
  32'h3d50a575 /* (0, 22, 9) */,
  32'h3da4db8a /* (28, 18, 9) */,
  32'h3dfaaa60 /* (24, 18, 9) */,
  32'h3e654448 /* (20, 18, 9) */,
  32'h3e8b9344 /* (16, 18, 9) */,
  32'h3e654448 /* (12, 18, 9) */,
  32'h3dfaaa60 /* (8, 18, 9) */,
  32'h3da4db8a /* (4, 18, 9) */,
  32'h3d8fa52c /* (0, 18, 9) */,
  32'h3da4db8a /* (28, 14, 9) */,
  32'h3dfaaa60 /* (24, 14, 9) */,
  32'h3e654448 /* (20, 14, 9) */,
  32'h3e8b9344 /* (16, 14, 9) */,
  32'h3e654448 /* (12, 14, 9) */,
  32'h3dfaaa60 /* (8, 14, 9) */,
  32'h3da4db8a /* (4, 14, 9) */,
  32'h3d8fa52c /* (0, 14, 9) */,
  32'h3d68b7a2 /* (28, 10, 9) */,
  32'h3da590e9 /* (24, 10, 9) */,
  32'h3e0cf021 /* (20, 10, 9) */,
  32'h3e21930d /* (16, 10, 9) */,
  32'h3e0cf021 /* (12, 10, 9) */,
  32'h3da590e9 /* (8, 10, 9) */,
  32'h3d68b7a2 /* (4, 10, 9) */,
  32'h3d50a575 /* (0, 10, 9) */,
  32'h3d2657dd /* (28, 6, 9) */,
  32'h3d584c0c /* (24, 6, 9) */,
  32'h3da96159 /* (20, 6, 9) */,
  32'h3db6b309 /* (16, 6, 9) */,
  32'h3da96159 /* (12, 6, 9) */,
  32'h3d584c0c /* (8, 6, 9) */,
  32'h3d2657dd /* (4, 6, 9) */,
  32'h3d1bc36a /* (0, 6, 9) */,
  32'h3d14de35 /* (28, 2, 9) */,
  32'h3d3291f6 /* (24, 2, 9) */,
  32'h3d833332 /* (20, 2, 9) */,
  32'h3d87d16b /* (16, 2, 9) */,
  32'h3d833332 /* (12, 2, 9) */,
  32'h3d3291f6 /* (8, 2, 9) */,
  32'h3d14de35 /* (4, 2, 9) */,
  32'h3d11b684 /* (0, 2, 9) */,
  32'h3d2d8e0e /* (28, 30, 5) */,
  32'h3d149b5c /* (24, 30, 5) */,
  32'h3d346b02 /* (20, 30, 5) */,
  32'h3d28d1e5 /* (16, 30, 5) */,
  32'h3d346b02 /* (12, 30, 5) */,
  32'h3d149b5c /* (8, 30, 5) */,
  32'h3d2d8e0e /* (4, 30, 5) */,
  32'h3d5dd7d1 /* (0, 30, 5) */,
  32'h3d153e19 /* (28, 26, 5) */,
  32'h3d22af34 /* (24, 26, 5) */,
  32'h3d6007ad /* (20, 26, 5) */,
  32'h3d5f53fb /* (16, 26, 5) */,
  32'h3d6007ad /* (12, 26, 5) */,
  32'h3d22af34 /* (8, 26, 5) */,
  32'h3d153e19 /* (4, 26, 5) */,
  32'h3d1b2f33 /* (0, 26, 5) */,
  32'h3d28e3b2 /* (28, 22, 5) */,
  32'h3d5ef675 /* (24, 22, 5) */,
  32'h3db0e528 /* (20, 22, 5) */,
  32'h3dc0863e /* (16, 22, 5) */,
  32'h3db0e528 /* (12, 22, 5) */,
  32'h3d5ef675 /* (8, 22, 5) */,
  32'h3d28e3b2 /* (4, 22, 5) */,
  32'h3d1cee15 /* (0, 22, 5) */,
  32'h3d53bb31 /* (28, 18, 5) */,
  32'h3d9bc970 /* (24, 18, 5) */,
  32'h3e095be4 /* (20, 18, 5) */,
  32'h3e2205a1 /* (16, 18, 5) */,
  32'h3e095be4 /* (12, 18, 5) */,
  32'h3d9bc970 /* (8, 18, 5) */,
  32'h3d53bb31 /* (4, 18, 5) */,
  32'h3d3b0a55 /* (0, 18, 5) */,
  32'h3d53bb31 /* (28, 14, 5) */,
  32'h3d9bc970 /* (24, 14, 5) */,
  32'h3e095be4 /* (20, 14, 5) */,
  32'h3e2205a1 /* (16, 14, 5) */,
  32'h3e095be4 /* (12, 14, 5) */,
  32'h3d9bc970 /* (8, 14, 5) */,
  32'h3d53bb31 /* (4, 14, 5) */,
  32'h3d3b0a55 /* (0, 14, 5) */,
  32'h3d28e3b2 /* (28, 10, 5) */,
  32'h3d5ef675 /* (24, 10, 5) */,
  32'h3db0e528 /* (20, 10, 5) */,
  32'h3dc0863e /* (16, 10, 5) */,
  32'h3db0e528 /* (12, 10, 5) */,
  32'h3d5ef675 /* (8, 10, 5) */,
  32'h3d28e3b2 /* (4, 10, 5) */,
  32'h3d1cee15 /* (0, 10, 5) */,
  32'h3d153e19 /* (28, 6, 5) */,
  32'h3d22af34 /* (24, 6, 5) */,
  32'h3d6007ad /* (20, 6, 5) */,
  32'h3d5f53fb /* (16, 6, 5) */,
  32'h3d6007ad /* (12, 6, 5) */,
  32'h3d22af34 /* (8, 6, 5) */,
  32'h3d153e19 /* (4, 6, 5) */,
  32'h3d1b2f33 /* (0, 6, 5) */,
  32'h3d2d8e0e /* (28, 2, 5) */,
  32'h3d149b5c /* (24, 2, 5) */,
  32'h3d346b02 /* (20, 2, 5) */,
  32'h3d28d1e5 /* (16, 2, 5) */,
  32'h3d346b02 /* (12, 2, 5) */,
  32'h3d149b5c /* (8, 2, 5) */,
  32'h3d2d8e0e /* (4, 2, 5) */,
  32'h3d5dd7d1 /* (0, 2, 5) */,
  32'h3d8b1391 /* (28, 30, 1) */,
  32'h3d15ce12 /* (24, 30, 1) */,
  32'h3d1cac31 /* (20, 30, 1) */,
  32'h3d09dfab /* (16, 30, 1) */,
  32'h3d1cac31 /* (12, 30, 1) */,
  32'h3d15ce12 /* (8, 30, 1) */,
  32'h3d8b1391 /* (4, 30, 1) */,
  32'h3e709592 /* (0, 30, 1) */,
  32'h3d222a9c /* (28, 26, 1) */,
  32'h3d169650 /* (24, 26, 1) */,
  32'h3d3dc5f0 /* (20, 26, 1) */,
  32'h3d34b66a /* (16, 26, 1) */,
  32'h3d3dc5f0 /* (12, 26, 1) */,
  32'h3d169650 /* (8, 26, 1) */,
  32'h3d222a9c /* (4, 26, 1) */,
  32'h3d3f59b8 /* (0, 26, 1) */,
  32'h3d1839e3 /* (28, 22, 1) */,
  32'h3d3f0366 /* (24, 22, 1) */,
  32'h3d91435f /* (20, 22, 1) */,
  32'h3d99ac24 /* (16, 22, 1) */,
  32'h3d91435f /* (12, 22, 1) */,
  32'h3d3f0366 /* (8, 22, 1) */,
  32'h3d1839e3 /* (4, 22, 1) */,
  32'h3d1142bb /* (0, 22, 1) */,
  32'h3d303352 /* (28, 18, 1) */,
  32'h3d7e759f /* (24, 18, 1) */,
  32'h3ddbed5a /* (20, 18, 1) */,
  32'h3dff32bb /* (16, 18, 1) */,
  32'h3ddbed5a /* (12, 18, 1) */,
  32'h3d7e759f /* (8, 18, 1) */,
  32'h3d303352 /* (4, 18, 1) */,
  32'h3d1ceee6 /* (0, 18, 1) */,
  32'h3d303352 /* (28, 14, 1) */,
  32'h3d7e759f /* (24, 14, 1) */,
  32'h3ddbed5a /* (20, 14, 1) */,
  32'h3dff32bb /* (16, 14, 1) */,
  32'h3ddbed5a /* (12, 14, 1) */,
  32'h3d7e759f /* (8, 14, 1) */,
  32'h3d303352 /* (4, 14, 1) */,
  32'h3d1ceee6 /* (0, 14, 1) */,
  32'h3d1839e3 /* (28, 10, 1) */,
  32'h3d3f0366 /* (24, 10, 1) */,
  32'h3d91435f /* (20, 10, 1) */,
  32'h3d99ac24 /* (16, 10, 1) */,
  32'h3d91435f /* (12, 10, 1) */,
  32'h3d3f0366 /* (8, 10, 1) */,
  32'h3d1839e3 /* (4, 10, 1) */,
  32'h3d1142bb /* (0, 10, 1) */,
  32'h3d222a9c /* (28, 6, 1) */,
  32'h3d169650 /* (24, 6, 1) */,
  32'h3d3dc5f0 /* (20, 6, 1) */,
  32'h3d34b66a /* (16, 6, 1) */,
  32'h3d3dc5f0 /* (12, 6, 1) */,
  32'h3d169650 /* (8, 6, 1) */,
  32'h3d222a9c /* (4, 6, 1) */,
  32'h3d3f59b8 /* (0, 6, 1) */,
  32'h3d8b1391 /* (28, 2, 1) */,
  32'h3d15ce12 /* (24, 2, 1) */,
  32'h3d1cac31 /* (20, 2, 1) */,
  32'h3d09dfab /* (16, 2, 1) */,
  32'h3d1cac31 /* (12, 2, 1) */,
  32'h3d15ce12 /* (8, 2, 1) */,
  32'h3d8b1391 /* (4, 2, 1) */,
  32'h3e709592 /* (0, 2, 1) */,
  32'h3d960c3c /* (31, 29, 29) */,
  32'h3d314afb /* (27, 29, 29) */,
  32'h3d144047 /* (23, 29, 29) */,
  32'h3d2fb3ed /* (19, 29, 29) */,
  32'h3d2aacf2 /* (15, 29, 29) */,
  32'h3d202a91 /* (11, 29, 29) */,
  32'h3d179239 /* (7, 29, 29) */,
  32'h3d68b01f /* (3, 29, 29) */,
  32'h3d1c3652 /* (31, 25, 29) */,
  32'h3d147808 /* (27, 25, 29) */,
  32'h3d2aad03 /* (23, 25, 29) */,
  32'h3d69f6ae /* (19, 25, 29) */,
  32'h3d6ce397 /* (15, 25, 29) */,
  32'h3d490aba /* (11, 25, 29) */,
  32'h3d1969a9 /* (7, 25, 29) */,
  32'h3d179239 /* (3, 25, 29) */,
  32'h3d1a3ccf /* (31, 21, 29) */,
  32'h3d2e4aa1 /* (27, 21, 29) */,
  32'h3d767d5d /* (23, 21, 29) */,
  32'h3dc2b35d /* (19, 21, 29) */,
  32'h3dceffa6 /* (15, 21, 29) */,
  32'h3d9d27e1 /* (11, 21, 29) */,
  32'h3d490aba /* (7, 21, 29) */,
  32'h3d202a91 /* (3, 21, 29) */,
  32'h3d202be8 /* (31, 17, 29) */,
  32'h3d424fe8 /* (27, 17, 29) */,
  32'h3d99caa3 /* (23, 17, 29) */,
  32'h3e068db8 /* (19, 17, 29) */,
  32'h3e151f83 /* (15, 17, 29) */,
  32'h3dceffa6 /* (11, 17, 29) */,
  32'h3d6ce397 /* (7, 17, 29) */,
  32'h3d2aacf2 /* (3, 17, 29) */,
  32'h3d269671 /* (31, 13, 29) */,
  32'h3d4466f8 /* (27, 13, 29) */,
  32'h3d942dc4 /* (23, 13, 29) */,
  32'h3df79892 /* (19, 13, 29) */,
  32'h3e068db8 /* (15, 13, 29) */,
  32'h3dc2b35d /* (11, 13, 29) */,
  32'h3d69f6ae /* (7, 13, 29) */,
  32'h3d2fb3ed /* (3, 13, 29) */,
  32'h3d126006 /* (31, 9, 29) */,
  32'h3d1addce /* (27, 9, 29) */,
  32'h3d48821f /* (23, 9, 29) */,
  32'h3d942dc4 /* (19, 9, 29) */,
  32'h3d99caa3 /* (15, 9, 29) */,
  32'h3d767d5d /* (11, 9, 29) */,
  32'h3d2aad03 /* (7, 9, 29) */,
  32'h3d144047 /* (3, 9, 29) */,
  32'h3d45ae9a /* (31, 5, 29) */,
  32'h3d1ccb4c /* (27, 5, 29) */,
  32'h3d1addce /* (23, 5, 29) */,
  32'h3d4466f8 /* (19, 5, 29) */,
  32'h3d424fe8 /* (15, 5, 29) */,
  32'h3d2e4aa1 /* (11, 5, 29) */,
  32'h3d147808 /* (7, 5, 29) */,
  32'h3d314afb /* (3, 5, 29) */,
  32'h3deb372d /* (31, 1, 29) */,
  32'h3d45ae9a /* (27, 1, 29) */,
  32'h3d126006 /* (23, 1, 29) */,
  32'h3d269671 /* (19, 1, 29) */,
  32'h3d202be8 /* (15, 1, 29) */,
  32'h3d1a3ccf /* (11, 1, 29) */,
  32'h3d1c3652 /* (7, 1, 29) */,
  32'h3d960c3c /* (3, 1, 29) */,
  32'h3d1c3652 /* (31, 29, 25) */,
  32'h3d147808 /* (27, 29, 25) */,
  32'h3d2aad03 /* (23, 29, 25) */,
  32'h3d69f6ae /* (19, 29, 25) */,
  32'h3d6ce397 /* (15, 29, 25) */,
  32'h3d490aba /* (11, 29, 25) */,
  32'h3d1969a9 /* (7, 29, 25) */,
  32'h3d179239 /* (3, 29, 25) */,
  32'h3d167b79 /* (31, 25, 25) */,
  32'h3d21f168 /* (27, 25, 25) */,
  32'h3d563bcb /* (23, 25, 25) */,
  32'h3da0c360 /* (19, 25, 25) */,
  32'h3da7bf05 /* (15, 25, 25) */,
  32'h3d84ce75 /* (11, 25, 25) */,
  32'h3d348078 /* (7, 25, 25) */,
  32'h3d1969a9 /* (3, 25, 25) */,
  32'h3d3efe62 /* (31, 21, 25) */,
  32'h3d5ff008 /* (27, 21, 25) */,
  32'h3da777c1 /* (23, 21, 25) */,
  32'h3e0aca9a /* (19, 21, 25) */,
  32'h3e165b49 /* (15, 21, 25) */,
  32'h3ddb1c7f /* (11, 21, 25) */,
  32'h3d84ce75 /* (7, 21, 25) */,
  32'h3d490aba /* (3, 21, 25) */,
  32'h3d5d3ed0 /* (31, 17, 25) */,
  32'h3d880917 /* (27, 17, 25) */,
  32'h3ddc94c6 /* (23, 17, 25) */,
  32'h3e45db44 /* (19, 17, 25) */,
  32'h3e5db918 /* (15, 17, 25) */,
  32'h3e165b49 /* (11, 17, 25) */,
  32'h3da7bf05 /* (7, 17, 25) */,
  32'h3d6ce397 /* (3, 17, 25) */,
  32'h3d5c17b6 /* (31, 13, 25) */,
  32'h3d849ae2 /* (27, 13, 25) */,
  32'h3dcf79e9 /* (23, 13, 25) */,
  32'h3e336d1b /* (19, 13, 25) */,
  32'h3e45db44 /* (15, 13, 25) */,
  32'h3e0aca9a /* (11, 13, 25) */,
  32'h3da0c360 /* (7, 13, 25) */,
  32'h3d69f6ae /* (3, 13, 25) */,
  32'h3d245baa /* (31, 9, 25) */,
  32'h3d39ba58 /* (27, 9, 25) */,
  32'h3d8354ed /* (23, 9, 25) */,
  32'h3dcf79e9 /* (19, 9, 25) */,
  32'h3ddc94c6 /* (15, 9, 25) */,
  32'h3da777c1 /* (11, 9, 25) */,
  32'h3d563bcb /* (7, 9, 25) */,
  32'h3d2aad03 /* (3, 9, 25) */,
  32'h3d151e01 /* (31, 5, 25) */,
  32'h3d170afd /* (27, 5, 25) */,
  32'h3d39ba58 /* (23, 5, 25) */,
  32'h3d849ae2 /* (19, 5, 25) */,
  32'h3d880917 /* (15, 5, 25) */,
  32'h3d5ff008 /* (11, 5, 25) */,
  32'h3d21f168 /* (7, 5, 25) */,
  32'h3d147808 /* (3, 5, 25) */,
  32'h3d2402bf /* (31, 1, 25) */,
  32'h3d151e01 /* (27, 1, 25) */,
  32'h3d245baa /* (23, 1, 25) */,
  32'h3d5c17b6 /* (19, 1, 25) */,
  32'h3d5d3ed0 /* (15, 1, 25) */,
  32'h3d3efe62 /* (11, 1, 25) */,
  32'h3d167b79 /* (7, 1, 25) */,
  32'h3d1c3652 /* (3, 1, 25) */,
  32'h3d1a3ccf /* (31, 29, 21) */,
  32'h3d2e4aa1 /* (27, 29, 21) */,
  32'h3d767d5d /* (23, 29, 21) */,
  32'h3dc2b35d /* (19, 29, 21) */,
  32'h3dceffa6 /* (15, 29, 21) */,
  32'h3d9d27e1 /* (11, 29, 21) */,
  32'h3d490aba /* (7, 29, 21) */,
  32'h3d202a91 /* (3, 29, 21) */,
  32'h3d3efe62 /* (31, 25, 21) */,
  32'h3d5ff008 /* (27, 25, 21) */,
  32'h3da777c1 /* (23, 25, 21) */,
  32'h3e0aca9a /* (19, 25, 21) */,
  32'h3e165b49 /* (15, 25, 21) */,
  32'h3ddb1c7f /* (11, 25, 21) */,
  32'h3d84ce75 /* (7, 25, 21) */,
  32'h3d490aba /* (3, 25, 21) */,
  32'h3d9352ec /* (31, 21, 21) */,
  32'h3db345e2 /* (27, 21, 21) */,
  32'h3e0ea5fd /* (23, 21, 21) */,
  32'h3e7af74d /* (19, 21, 21) */,
  32'h3e8b66c2 /* (15, 21, 21) */,
  32'h3e4089a2 /* (11, 21, 21) */,
  32'h3ddb1c7f /* (7, 21, 21) */,
  32'h3d9d27e1 /* (3, 21, 21) */,
  32'h3dc031e4 /* (31, 17, 21) */,
  32'h3df05994 /* (27, 17, 21) */,
  32'h3e49046a /* (23, 17, 21) */,
  32'h3eba8e90 /* (19, 17, 21) */,
  32'h3ed4648a /* (15, 17, 21) */,
  32'h3e8b66c2 /* (11, 17, 21) */,
  32'h3e165b49 /* (7, 17, 21) */,
  32'h3dceffa6 /* (3, 17, 21) */,
  32'h3db58f74 /* (31, 13, 21) */,
  32'h3de04254 /* (27, 13, 21) */,
  32'h3e37494b /* (23, 13, 21) */,
  32'h3ea5d30f /* (19, 13, 21) */,
  32'h3eba8e90 /* (15, 13, 21) */,
  32'h3e7af74d /* (11, 13, 21) */,
  32'h3e0aca9a /* (7, 13, 21) */,
  32'h3dc2b35d /* (3, 13, 21) */,
  32'h3d68852c /* (31, 9, 21) */,
  32'h3d8b02ad /* (27, 9, 21) */,
  32'h3dd6aa1b /* (23, 9, 21) */,
  32'h3e37494b /* (19, 9, 21) */,
  32'h3e49046a /* (15, 9, 21) */,
  32'h3e0ea5fd /* (11, 9, 21) */,
  32'h3da777c1 /* (7, 9, 21) */,
  32'h3d767d5d /* (3, 9, 21) */,
  32'h3d26c9db /* (31, 5, 21) */,
  32'h3d3fb488 /* (27, 5, 21) */,
  32'h3d8b02ad /* (23, 5, 21) */,
  32'h3de04254 /* (19, 5, 21) */,
  32'h3df05994 /* (15, 5, 21) */,
  32'h3db345e2 /* (11, 5, 21) */,
  32'h3d5ff008 /* (7, 5, 21) */,
  32'h3d2e4aa1 /* (3, 5, 21) */,
  32'h3d151591 /* (31, 1, 21) */,
  32'h3d26c9db /* (27, 1, 21) */,
  32'h3d68852c /* (23, 1, 21) */,
  32'h3db58f74 /* (19, 1, 21) */,
  32'h3dc031e4 /* (15, 1, 21) */,
  32'h3d9352ec /* (11, 1, 21) */,
  32'h3d3efe62 /* (7, 1, 21) */,
  32'h3d1a3ccf /* (3, 1, 21) */,
  32'h3d202be8 /* (31, 29, 17) */,
  32'h3d424fe8 /* (27, 29, 17) */,
  32'h3d99caa3 /* (23, 29, 17) */,
  32'h3e068db8 /* (19, 29, 17) */,
  32'h3e151f83 /* (15, 29, 17) */,
  32'h3dceffa6 /* (11, 29, 17) */,
  32'h3d6ce397 /* (7, 29, 17) */,
  32'h3d2aacf2 /* (3, 29, 17) */,
  32'h3d5d3ed0 /* (31, 25, 17) */,
  32'h3d880917 /* (27, 25, 17) */,
  32'h3ddc94c6 /* (23, 25, 17) */,
  32'h3e45db44 /* (19, 25, 17) */,
  32'h3e5db918 /* (15, 25, 17) */,
  32'h3e165b49 /* (11, 25, 17) */,
  32'h3da7bf05 /* (7, 25, 17) */,
  32'h3d6ce397 /* (3, 25, 17) */,
  32'h3dc031e4 /* (31, 21, 17) */,
  32'h3df05994 /* (27, 21, 17) */,
  32'h3e49046a /* (23, 21, 17) */,
  32'h3eba8e90 /* (19, 21, 17) */,
  32'h3ed4648a /* (15, 21, 17) */,
  32'h3e8b66c2 /* (11, 21, 17) */,
  32'h3e165b49 /* (7, 21, 17) */,
  32'h3dceffa6 /* (3, 21, 17) */,
  32'h3e09bd27 /* (31, 17, 17) */,
  32'h3e2edbb4 /* (27, 17, 17) */,
  32'h3e969108 /* (23, 17, 17) */,
  32'h3f1092e5 /* (19, 17, 17) */,
  32'h3f275a64 /* (15, 17, 17) */,
  32'h3ed4648a /* (11, 17, 17) */,
  32'h3e5db918 /* (7, 17, 17) */,
  32'h3e151f83 /* (3, 17, 17) */,
  32'h3df92d6c /* (31, 13, 17) */,
  32'h3e1d0a10 /* (27, 13, 17) */,
  32'h3e8557f4 /* (23, 13, 17) */,
  32'h3efbd9fe /* (19, 13, 17) */,
  32'h3f1092e5 /* (15, 13, 17) */,
  32'h3eba8e90 /* (11, 13, 17) */,
  32'h3e45db44 /* (7, 13, 17) */,
  32'h3e068db8 /* (3, 13, 17) */,
  32'h3d8f3655 /* (31, 9, 17) */,
  32'h3db198fc /* (27, 9, 17) */,
  32'h3e123783 /* (23, 9, 17) */,
  32'h3e8557f4 /* (19, 9, 17) */,
  32'h3e969108 /* (15, 9, 17) */,
  32'h3e49046a /* (11, 9, 17) */,
  32'h3ddc94c6 /* (7, 9, 17) */,
  32'h3d99caa3 /* (3, 9, 17) */,
  32'h3d35f880 /* (31, 5, 17) */,
  32'h3d5e11d0 /* (27, 5, 17) */,
  32'h3db198fc /* (23, 5, 17) */,
  32'h3e1d0a10 /* (19, 5, 17) */,
  32'h3e2edbb4 /* (15, 5, 17) */,
  32'h3df05994 /* (11, 5, 17) */,
  32'h3d880917 /* (7, 5, 17) */,
  32'h3d424fe8 /* (3, 5, 17) */,
  32'h3d167d01 /* (31, 1, 17) */,
  32'h3d35f880 /* (27, 1, 17) */,
  32'h3d8f3655 /* (23, 1, 17) */,
  32'h3df92d6c /* (19, 1, 17) */,
  32'h3e09bd27 /* (15, 1, 17) */,
  32'h3dc031e4 /* (11, 1, 17) */,
  32'h3d5d3ed0 /* (7, 1, 17) */,
  32'h3d202be8 /* (3, 1, 17) */,
  32'h3d269671 /* (31, 29, 13) */,
  32'h3d4466f8 /* (27, 29, 13) */,
  32'h3d942dc4 /* (23, 29, 13) */,
  32'h3df79892 /* (19, 29, 13) */,
  32'h3e068db8 /* (15, 29, 13) */,
  32'h3dc2b35d /* (11, 29, 13) */,
  32'h3d69f6ae /* (7, 29, 13) */,
  32'h3d2fb3ed /* (3, 29, 13) */,
  32'h3d5c17b6 /* (31, 25, 13) */,
  32'h3d849ae2 /* (27, 25, 13) */,
  32'h3dcf79e9 /* (23, 25, 13) */,
  32'h3e336d1b /* (19, 25, 13) */,
  32'h3e45db44 /* (15, 25, 13) */,
  32'h3e0aca9a /* (11, 25, 13) */,
  32'h3da0c360 /* (7, 25, 13) */,
  32'h3d69f6ae /* (3, 25, 13) */,
  32'h3db58f74 /* (31, 21, 13) */,
  32'h3de04254 /* (27, 21, 13) */,
  32'h3e37494b /* (23, 21, 13) */,
  32'h3ea5d30f /* (19, 21, 13) */,
  32'h3eba8e90 /* (15, 21, 13) */,
  32'h3e7af74d /* (11, 21, 13) */,
  32'h3e0aca9a /* (7, 21, 13) */,
  32'h3dc2b35d /* (3, 21, 13) */,
  32'h3df92d6c /* (31, 17, 13) */,
  32'h3e1d0a10 /* (27, 17, 13) */,
  32'h3e8557f4 /* (23, 17, 13) */,
  32'h3efbd9fe /* (19, 17, 13) */,
  32'h3f1092e5 /* (15, 17, 13) */,
  32'h3eba8e90 /* (11, 17, 13) */,
  32'h3e45db44 /* (7, 17, 13) */,
  32'h3e068db8 /* (3, 17, 13) */,
  32'h3de602d9 /* (31, 13, 13) */,
  32'h3e0f99f2 /* (27, 13, 13) */,
  32'h3e6f82ab /* (23, 13, 13) */,
  32'h3edd8ee5 /* (19, 13, 13) */,
  32'h3efbd9fe /* (15, 13, 13) */,
  32'h3ea5d30f /* (11, 13, 13) */,
  32'h3e336d1b /* (7, 13, 13) */,
  32'h3df79892 /* (3, 13, 13) */,
  32'h3d8ac476 /* (31, 9, 13) */,
  32'h3da95898 /* (27, 9, 13) */,
  32'h3e076ebd /* (23, 9, 13) */,
  32'h3e6f82ab /* (19, 9, 13) */,
  32'h3e8557f4 /* (15, 9, 13) */,
  32'h3e37494b /* (11, 9, 13) */,
  32'h3dcf79e9 /* (7, 9, 13) */,
  32'h3d942dc4 /* (3, 9, 13) */,
  32'h3d398f3f /* (31, 5, 13) */,
  32'h3d5ce99d /* (27, 5, 13) */,
  32'h3da95898 /* (23, 5, 13) */,
  32'h3e0f99f2 /* (19, 5, 13) */,
  32'h3e1d0a10 /* (15, 5, 13) */,
  32'h3de04254 /* (11, 5, 13) */,
  32'h3d849ae2 /* (7, 5, 13) */,
  32'h3d4466f8 /* (3, 5, 13) */,
  32'h3d1e42f1 /* (31, 1, 13) */,
  32'h3d398f3f /* (27, 1, 13) */,
  32'h3d8ac476 /* (23, 1, 13) */,
  32'h3de602d9 /* (19, 1, 13) */,
  32'h3df92d6c /* (15, 1, 13) */,
  32'h3db58f74 /* (11, 1, 13) */,
  32'h3d5c17b6 /* (7, 1, 13) */,
  32'h3d269671 /* (3, 1, 13) */,
  32'h3d126006 /* (31, 29, 9) */,
  32'h3d1addce /* (27, 29, 9) */,
  32'h3d48821f /* (23, 29, 9) */,
  32'h3d942dc4 /* (19, 29, 9) */,
  32'h3d99caa3 /* (15, 29, 9) */,
  32'h3d767d5d /* (11, 29, 9) */,
  32'h3d2aad03 /* (7, 29, 9) */,
  32'h3d144047 /* (3, 29, 9) */,
  32'h3d245baa /* (31, 25, 9) */,
  32'h3d39ba58 /* (27, 25, 9) */,
  32'h3d8354ed /* (23, 25, 9) */,
  32'h3dcf79e9 /* (19, 25, 9) */,
  32'h3ddc94c6 /* (15, 25, 9) */,
  32'h3da777c1 /* (11, 25, 9) */,
  32'h3d563bcb /* (7, 25, 9) */,
  32'h3d2aad03 /* (3, 25, 9) */,
  32'h3d68852c /* (31, 21, 9) */,
  32'h3d8b02ad /* (27, 21, 9) */,
  32'h3dd6aa1b /* (23, 21, 9) */,
  32'h3e37494b /* (19, 21, 9) */,
  32'h3e49046a /* (15, 21, 9) */,
  32'h3e0ea5fd /* (11, 21, 9) */,
  32'h3da777c1 /* (7, 21, 9) */,
  32'h3d767d5d /* (3, 21, 9) */,
  32'h3d8f3655 /* (31, 17, 9) */,
  32'h3db198fc /* (27, 17, 9) */,
  32'h3e123783 /* (23, 17, 9) */,
  32'h3e8557f4 /* (19, 17, 9) */,
  32'h3e969108 /* (15, 17, 9) */,
  32'h3e49046a /* (11, 17, 9) */,
  32'h3ddc94c6 /* (7, 17, 9) */,
  32'h3d99caa3 /* (3, 17, 9) */,
  32'h3d8ac476 /* (31, 13, 9) */,
  32'h3da95898 /* (27, 13, 9) */,
  32'h3e076ebd /* (23, 13, 9) */,
  32'h3e6f82ab /* (19, 13, 9) */,
  32'h3e8557f4 /* (15, 13, 9) */,
  32'h3e37494b /* (11, 13, 9) */,
  32'h3dcf79e9 /* (7, 13, 9) */,
  32'h3d942dc4 /* (3, 13, 9) */,
  32'h3d3ee791 /* (31, 9, 9) */,
  32'h3d5e7d3b /* (27, 9, 9) */,
  32'h3da4cfbf /* (23, 9, 9) */,
  32'h3e076ebd /* (19, 9, 9) */,
  32'h3e123783 /* (15, 9, 9) */,
  32'h3dd6aa1b /* (11, 9, 9) */,
  32'h3d8354ed /* (7, 9, 9) */,
  32'h3d48821f /* (3, 9, 9) */,
  32'h3d170f20 /* (31, 5, 9) */,
  32'h3d24f869 /* (27, 5, 9) */,
  32'h3d5e7d3b /* (23, 5, 9) */,
  32'h3da95898 /* (19, 5, 9) */,
  32'h3db198fc /* (15, 5, 9) */,
  32'h3d8b02ad /* (11, 5, 9) */,
  32'h3d39ba58 /* (7, 5, 9) */,
  32'h3d1addce /* (3, 5, 9) */,
  32'h3d11a602 /* (31, 1, 9) */,
  32'h3d170f20 /* (27, 1, 9) */,
  32'h3d3ee791 /* (23, 1, 9) */,
  32'h3d8ac476 /* (19, 1, 9) */,
  32'h3d8f3655 /* (15, 1, 9) */,
  32'h3d68852c /* (11, 1, 9) */,
  32'h3d245baa /* (7, 1, 9) */,
  32'h3d126006 /* (3, 1, 9) */,
  32'h3d45ae9a /* (31, 29, 5) */,
  32'h3d1ccb4c /* (27, 29, 5) */,
  32'h3d1addce /* (23, 29, 5) */,
  32'h3d4466f8 /* (19, 29, 5) */,
  32'h3d424fe8 /* (15, 29, 5) */,
  32'h3d2e4aa1 /* (11, 29, 5) */,
  32'h3d147808 /* (7, 29, 5) */,
  32'h3d314afb /* (3, 29, 5) */,
  32'h3d151e01 /* (31, 25, 5) */,
  32'h3d170afd /* (27, 25, 5) */,
  32'h3d39ba58 /* (23, 25, 5) */,
  32'h3d849ae2 /* (19, 25, 5) */,
  32'h3d880917 /* (15, 25, 5) */,
  32'h3d5ff008 /* (11, 25, 5) */,
  32'h3d21f168 /* (7, 25, 5) */,
  32'h3d147808 /* (3, 25, 5) */,
  32'h3d26c9db /* (31, 21, 5) */,
  32'h3d3fb488 /* (27, 21, 5) */,
  32'h3d8b02ad /* (23, 21, 5) */,
  32'h3de04254 /* (19, 21, 5) */,
  32'h3df05994 /* (15, 21, 5) */,
  32'h3db345e2 /* (11, 21, 5) */,
  32'h3d5ff008 /* (7, 21, 5) */,
  32'h3d2e4aa1 /* (3, 21, 5) */,
  32'h3d35f880 /* (31, 17, 5) */,
  32'h3d5e11d0 /* (27, 17, 5) */,
  32'h3db198fc /* (23, 17, 5) */,
  32'h3e1d0a10 /* (19, 17, 5) */,
  32'h3e2edbb4 /* (15, 17, 5) */,
  32'h3df05994 /* (11, 17, 5) */,
  32'h3d880917 /* (7, 17, 5) */,
  32'h3d424fe8 /* (3, 17, 5) */,
  32'h3d398f3f /* (31, 13, 5) */,
  32'h3d5ce99d /* (27, 13, 5) */,
  32'h3da95898 /* (23, 13, 5) */,
  32'h3e0f99f2 /* (19, 13, 5) */,
  32'h3e1d0a10 /* (15, 13, 5) */,
  32'h3de04254 /* (11, 13, 5) */,
  32'h3d849ae2 /* (7, 13, 5) */,
  32'h3d4466f8 /* (3, 13, 5) */,
  32'h3d170f20 /* (31, 9, 5) */,
  32'h3d24f869 /* (27, 9, 5) */,
  32'h3d5e7d3b /* (23, 9, 5) */,
  32'h3da95898 /* (19, 9, 5) */,
  32'h3db198fc /* (15, 9, 5) */,
  32'h3d8b02ad /* (11, 9, 5) */,
  32'h3d39ba58 /* (7, 9, 5) */,
  32'h3d1addce /* (3, 9, 5) */,
  32'h3d249f29 /* (31, 5, 5) */,
  32'h3d15ac37 /* (27, 5, 5) */,
  32'h3d24f869 /* (23, 5, 5) */,
  32'h3d5ce99d /* (19, 5, 5) */,
  32'h3d5e11d0 /* (15, 5, 5) */,
  32'h3d3fb488 /* (11, 5, 5) */,
  32'h3d170afd /* (7, 5, 5) */,
  32'h3d1ccb4c /* (3, 5, 5) */,
  32'h3d6890ff /* (31, 1, 5) */,
  32'h3d249f29 /* (27, 1, 5) */,
  32'h3d170f20 /* (23, 1, 5) */,
  32'h3d398f3f /* (19, 1, 5) */,
  32'h3d35f880 /* (15, 1, 5) */,
  32'h3d26c9db /* (11, 1, 5) */,
  32'h3d151e01 /* (7, 1, 5) */,
  32'h3d45ae9a /* (3, 1, 5) */,
  32'h3deb372d /* (31, 29, 1) */,
  32'h3d45ae9a /* (27, 29, 1) */,
  32'h3d126006 /* (23, 29, 1) */,
  32'h3d269671 /* (19, 29, 1) */,
  32'h3d202be8 /* (15, 29, 1) */,
  32'h3d1a3ccf /* (11, 29, 1) */,
  32'h3d1c3652 /* (7, 29, 1) */,
  32'h3d960c3c /* (3, 29, 1) */,
  32'h3d2402bf /* (31, 25, 1) */,
  32'h3d151e01 /* (27, 25, 1) */,
  32'h3d245baa /* (23, 25, 1) */,
  32'h3d5c17b6 /* (19, 25, 1) */,
  32'h3d5d3ed0 /* (15, 25, 1) */,
  32'h3d3efe62 /* (11, 25, 1) */,
  32'h3d167b79 /* (7, 25, 1) */,
  32'h3d1c3652 /* (3, 25, 1) */,
  32'h3d151591 /* (31, 21, 1) */,
  32'h3d26c9db /* (27, 21, 1) */,
  32'h3d68852c /* (23, 21, 1) */,
  32'h3db58f74 /* (19, 21, 1) */,
  32'h3dc031e4 /* (15, 21, 1) */,
  32'h3d9352ec /* (11, 21, 1) */,
  32'h3d3efe62 /* (7, 21, 1) */,
  32'h3d1a3ccf /* (3, 21, 1) */,
  32'h3d167d01 /* (31, 17, 1) */,
  32'h3d35f880 /* (27, 17, 1) */,
  32'h3d8f3655 /* (23, 17, 1) */,
  32'h3df92d6c /* (19, 17, 1) */,
  32'h3e09bd27 /* (15, 17, 1) */,
  32'h3dc031e4 /* (11, 17, 1) */,
  32'h3d5d3ed0 /* (7, 17, 1) */,
  32'h3d202be8 /* (3, 17, 1) */,
  32'h3d1e42f1 /* (31, 13, 1) */,
  32'h3d398f3f /* (27, 13, 1) */,
  32'h3d8ac476 /* (23, 13, 1) */,
  32'h3de602d9 /* (19, 13, 1) */,
  32'h3df92d6c /* (15, 13, 1) */,
  32'h3db58f74 /* (11, 13, 1) */,
  32'h3d5c17b6 /* (7, 13, 1) */,
  32'h3d269671 /* (3, 13, 1) */,
  32'h3d11a602 /* (31, 9, 1) */,
  32'h3d170f20 /* (27, 9, 1) */,
  32'h3d3ee791 /* (23, 9, 1) */,
  32'h3d8ac476 /* (19, 9, 1) */,
  32'h3d8f3655 /* (15, 9, 1) */,
  32'h3d68852c /* (11, 9, 1) */,
  32'h3d245baa /* (7, 9, 1) */,
  32'h3d126006 /* (3, 9, 1) */,
  32'h3d6890ff /* (31, 5, 1) */,
  32'h3d249f29 /* (27, 5, 1) */,
  32'h3d170f20 /* (23, 5, 1) */,
  32'h3d398f3f /* (19, 5, 1) */,
  32'h3d35f880 /* (15, 5, 1) */,
  32'h3d26c9db /* (11, 5, 1) */,
  32'h3d151e01 /* (7, 5, 1) */,
  32'h3d45ae9a /* (3, 5, 1) */,
  32'h3ec3aed4 /* (31, 1, 1) */,
  32'h3d6890ff /* (27, 1, 1) */,
  32'h3d11a602 /* (23, 1, 1) */,
  32'h3d1e42f1 /* (19, 1, 1) */,
  32'h3d167d01 /* (15, 1, 1) */,
  32'h3d151591 /* (11, 1, 1) */,
  32'h3d2402bf /* (7, 1, 1) */,
  32'h3deb372d /* (3, 1, 1) */,
  32'h3d866355 /* (30, 29, 29) */,
  32'h3d211f1b /* (26, 29, 29) */,
  32'h3d18cb02 /* (22, 29, 29) */,
  32'h3d3188e3 /* (18, 29, 29) */,
  32'h3d3188e3 /* (14, 29, 29) */,
  32'h3d18cb02 /* (10, 29, 29) */,
  32'h3d211f1b /* (6, 29, 29) */,
  32'h3d866355 /* (2, 29, 29) */,
  32'h3d1a2949 /* (30, 25, 29) */,
  32'h3d159d44 /* (26, 25, 29) */,
  32'h3d387393 /* (22, 25, 29) */,
  32'h3d71c736 /* (18, 25, 29) */,
  32'h3d71c736 /* (14, 25, 29) */,
  32'h3d387393 /* (10, 25, 29) */,
  32'h3d159d44 /* (6, 25, 29) */,
  32'h3d1a2949 /* (2, 25, 29) */,
  32'h3d1c5f03 /* (30, 21, 29) */,
  32'h3d39bb76 /* (26, 21, 29) */,
  32'h3d8ae43c /* (22, 21, 29) */,
  32'h3dce7d45 /* (18, 21, 29) */,
  32'h3dce7d45 /* (14, 21, 29) */,
  32'h3d8ae43c /* (10, 21, 29) */,
  32'h3d39bb76 /* (6, 21, 29) */,
  32'h3d1c5f03 /* (2, 21, 29) */,
  32'h3d240321 /* (30, 17, 29) */,
  32'h3d54ba37 /* (26, 17, 29) */,
  32'h3db22d06 /* (22, 17, 29) */,
  32'h3e11d12f /* (18, 17, 29) */,
  32'h3e11d12f /* (14, 17, 29) */,
  32'h3db22d06 /* (10, 17, 29) */,
  32'h3d54ba37 /* (6, 17, 29) */,
  32'h3d240321 /* (2, 17, 29) */,
  32'h3d29e985 /* (30, 13, 29) */,
  32'h3d54a03b /* (26, 13, 29) */,
  32'h3da99659 /* (22, 13, 29) */,
  32'h3e04d0b8 /* (18, 13, 29) */,
  32'h3e04d0b8 /* (14, 13, 29) */,
  32'h3da99659 /* (10, 13, 29) */,
  32'h3d54a03b /* (6, 13, 29) */,
  32'h3d29e985 /* (2, 13, 29) */,
  32'h3d12f42a /* (30, 9, 29) */,
  32'h3d215063 /* (26, 9, 29) */,
  32'h3d5dae2c /* (22, 9, 29) */,
  32'h3d9b2a7b /* (18, 9, 29) */,
  32'h3d9b2a7b /* (14, 9, 29) */,
  32'h3d5dae2c /* (10, 9, 29) */,
  32'h3d215063 /* (6, 9, 29) */,
  32'h3d12f42a /* (2, 9, 29) */,
  32'h3d3cd255 /* (30, 5, 29) */,
  32'h3d16d305 /* (26, 5, 29) */,
  32'h3d2344c4 /* (22, 5, 29) */,
  32'h3d487174 /* (18, 5, 29) */,
  32'h3d487174 /* (14, 5, 29) */,
  32'h3d2344c4 /* (10, 5, 29) */,
  32'h3d16d305 /* (6, 5, 29) */,
  32'h3d3cd255 /* (2, 5, 29) */,
  32'h3dbfa8df /* (30, 1, 29) */,
  32'h3d2ba889 /* (26, 1, 29) */,
  32'h3d14c0fd /* (22, 1, 29) */,
  32'h3d276174 /* (18, 1, 29) */,
  32'h3d276174 /* (14, 1, 29) */,
  32'h3d14c0fd /* (10, 1, 29) */,
  32'h3d2ba889 /* (6, 1, 29) */,
  32'h3dbfa8df /* (2, 1, 29) */,
  32'h3d1a2949 /* (30, 29, 25) */,
  32'h3d159d44 /* (26, 29, 25) */,
  32'h3d387393 /* (22, 29, 25) */,
  32'h3d71c736 /* (18, 29, 25) */,
  32'h3d71c736 /* (14, 29, 25) */,
  32'h3d387393 /* (10, 29, 25) */,
  32'h3d159d44 /* (6, 29, 25) */,
  32'h3d1a2949 /* (2, 29, 25) */,
  32'h3d1777c7 /* (30, 25, 25) */,
  32'h3d29a602 /* (26, 25, 25) */,
  32'h3d6deb12 /* (22, 25, 25) */,
  32'h3da8d240 /* (18, 25, 25) */,
  32'h3da8d240 /* (14, 25, 25) */,
  32'h3d6deb12 /* (10, 25, 25) */,
  32'h3d29a602 /* (6, 25, 25) */,
  32'h3d1777c7 /* (2, 25, 25) */,
  32'h3d42a7b8 /* (30, 21, 25) */,
  32'h3d71ecf9 /* (26, 21, 25) */,
  32'h3dbf3f1d /* (22, 21, 25) */,
  32'h3e14a5c9 /* (18, 21, 25) */,
  32'h3e14a5c9 /* (14, 21, 25) */,
  32'h3dbf3f1d /* (10, 21, 25) */,
  32'h3d71ecf9 /* (6, 21, 25) */,
  32'h3d42a7b8 /* (2, 21, 25) */,
  32'h3d62f778 /* (30, 17, 25) */,
  32'h3d95be73 /* (26, 17, 25) */,
  32'h3e009a19 /* (22, 17, 25) */,
  32'h3e57a44b /* (18, 17, 25) */,
  32'h3e57a44b /* (14, 17, 25) */,
  32'h3e009a19 /* (10, 17, 25) */,
  32'h3d95be73 /* (6, 17, 25) */,
  32'h3d62f778 /* (2, 17, 25) */,
  32'h3d6129ae /* (30, 13, 25) */,
  32'h3d90c8a7 /* (26, 13, 25) */,
  32'h3defa49b /* (22, 13, 25) */,
  32'h3e41f14c /* (18, 13, 25) */,
  32'h3e41f14c /* (14, 13, 25) */,
  32'h3defa49b /* (10, 13, 25) */,
  32'h3d90c8a7 /* (6, 13, 25) */,
  32'h3d6129ae /* (2, 13, 25) */,
  32'h3d26a1b5 /* (30, 9, 25) */,
  32'h3d45eb5b /* (26, 9, 25) */,
  32'h3d94014f /* (22, 9, 25) */,
  32'h3ddc09d8 /* (18, 9, 25) */,
  32'h3ddc09d8 /* (14, 9, 25) */,
  32'h3d94014f /* (10, 9, 25) */,
  32'h3d45eb5b /* (6, 9, 25) */,
  32'h3d26a1b5 /* (2, 9, 25) */,
  32'h3d14b1c0 /* (30, 5, 25) */,
  32'h3d1b2471 /* (26, 5, 25) */,
  32'h3d4b3dc7 /* (22, 5, 25) */,
  32'h3d8a0000 /* (18, 5, 25) */,
  32'h3d8a0000 /* (14, 5, 25) */,
  32'h3d4b3dc7 /* (10, 5, 25) */,
  32'h3d1b2471 /* (6, 5, 25) */,
  32'h3d14b1c0 /* (2, 5, 25) */,
  32'h3d20a35e /* (30, 1, 25) */,
  32'h3d146a43 /* (26, 1, 25) */,
  32'h3d305430 /* (22, 1, 25) */,
  32'h3d62906c /* (18, 1, 25) */,
  32'h3d62906c /* (14, 1, 25) */,
  32'h3d305430 /* (10, 1, 25) */,
  32'h3d146a43 /* (6, 1, 25) */,
  32'h3d20a35e /* (2, 1, 25) */,
  32'h3d1c5f03 /* (30, 29, 21) */,
  32'h3d39bb76 /* (26, 29, 21) */,
  32'h3d8ae43c /* (22, 29, 21) */,
  32'h3dce7d45 /* (18, 29, 21) */,
  32'h3dce7d45 /* (14, 29, 21) */,
  32'h3d8ae43c /* (10, 29, 21) */,
  32'h3d39bb76 /* (6, 29, 21) */,
  32'h3d1c5f03 /* (2, 29, 21) */,
  32'h3d42a7b8 /* (30, 25, 21) */,
  32'h3d71ecf9 /* (26, 25, 21) */,
  32'h3dbf3f1d /* (22, 25, 21) */,
  32'h3e14a5c9 /* (18, 25, 21) */,
  32'h3e14a5c9 /* (14, 25, 21) */,
  32'h3dbf3f1d /* (10, 25, 21) */,
  32'h3d71ecf9 /* (6, 25, 21) */,
  32'h3d42a7b8 /* (2, 25, 21) */,
  32'h3d96eb50 /* (30, 21, 21) */,
  32'h3dc480ba /* (26, 21, 21) */,
  32'h3e257fc6 /* (22, 21, 21) */,
  32'h3e882756 /* (18, 21, 21) */,
  32'h3e882756 /* (14, 21, 21) */,
  32'h3e257fc6 /* (10, 21, 21) */,
  32'h3dc480ba /* (6, 21, 21) */,
  32'h3d96eb50 /* (2, 21, 21) */,
  32'h3dc59b81 /* (30, 17, 21) */,
  32'h3e0533d0 /* (26, 17, 21) */,
  32'h3e6c6ac0 /* (22, 17, 21) */,
  32'h3eccf8ff /* (18, 17, 21) */,
  32'h3eccf8ff /* (14, 17, 21) */,
  32'h3e6c6ac0 /* (10, 17, 21) */,
  32'h3e0533d0 /* (6, 17, 21) */,
  32'h3dc59b81 /* (2, 17, 21) */,
  32'h3dba5db4 /* (30, 13, 21) */,
  32'h3df74dbc /* (26, 13, 21) */,
  32'h3e562fb1 /* (22, 13, 21) */,
  32'h3eb517ce /* (18, 13, 21) */,
  32'h3eb517ce /* (14, 13, 21) */,
  32'h3e562fb1 /* (10, 13, 21) */,
  32'h3df74dbc /* (6, 13, 21) */,
  32'h3dba5db4 /* (2, 13, 21) */,
  32'h3d6d9fa3 /* (30, 9, 21) */,
  32'h3d9750ce /* (26, 9, 21) */,
  32'h3df71c69 /* (22, 9, 21) */,
  32'h3e458f30 /* (18, 9, 21) */,
  32'h3e458f30 /* (14, 9, 21) */,
  32'h3df71c69 /* (10, 9, 21) */,
  32'h3d9750ce /* (6, 9, 21) */,
  32'h3d6d9fa3 /* (2, 9, 21) */,
  32'h3d29823f /* (30, 5, 21) */,
  32'h3d4d9045 /* (26, 5, 21) */,
  32'h3d9d9380 /* (22, 5, 21) */,
  32'h3deed79f /* (18, 5, 21) */,
  32'h3deed79f /* (14, 5, 21) */,
  32'h3d9d9380 /* (10, 5, 21) */,
  32'h3d4d9045 /* (6, 5, 21) */,
  32'h3d29823f /* (2, 5, 21) */,
  32'h3d16ed42 /* (30, 1, 21) */,
  32'h3d31191b /* (26, 1, 21) */,
  32'h3d829849 /* (22, 1, 21) */,
  32'h3dc01db4 /* (18, 1, 21) */,
  32'h3dc01db4 /* (14, 1, 21) */,
  32'h3d829849 /* (10, 1, 21) */,
  32'h3d31191b /* (6, 1, 21) */,
  32'h3d16ed42 /* (2, 1, 21) */,
  32'h3d240321 /* (30, 29, 17) */,
  32'h3d54ba37 /* (26, 29, 17) */,
  32'h3db22d06 /* (22, 29, 17) */,
  32'h3e11d12f /* (18, 29, 17) */,
  32'h3e11d12f /* (14, 29, 17) */,
  32'h3db22d06 /* (10, 29, 17) */,
  32'h3d54ba37 /* (6, 29, 17) */,
  32'h3d240321 /* (2, 29, 17) */,
  32'h3d62f778 /* (30, 25, 17) */,
  32'h3d95be73 /* (26, 25, 17) */,
  32'h3e009a19 /* (22, 25, 17) */,
  32'h3e57a44b /* (18, 25, 17) */,
  32'h3e57a44b /* (14, 25, 17) */,
  32'h3e009a19 /* (10, 25, 17) */,
  32'h3d95be73 /* (6, 25, 17) */,
  32'h3d62f778 /* (2, 25, 17) */,
  32'h3dc59b81 /* (30, 21, 17) */,
  32'h3e0533d0 /* (26, 21, 17) */,
  32'h3e6c6ac0 /* (22, 21, 17) */,
  32'h3eccf8ff /* (18, 21, 17) */,
  32'h3eccf8ff /* (14, 21, 17) */,
  32'h3e6c6ac0 /* (10, 21, 17) */,
  32'h3e0533d0 /* (6, 21, 17) */,
  32'h3dc59b81 /* (2, 21, 17) */,
  32'h3e0de5f8 /* (30, 17, 17) */,
  32'h3e430b11 /* (26, 17, 17) */,
  32'h3eb2925b /* (22, 17, 17) */,
  32'h3f202f9a /* (18, 17, 17) */,
  32'h3f202f9a /* (14, 17, 17) */,
  32'h3eb2925b /* (10, 17, 17) */,
  32'h3e430b11 /* (6, 17, 17) */,
  32'h3e0de5f8 /* (2, 17, 17) */,
  32'h3e003b1e /* (30, 13, 17) */,
  32'h3e2ea39a /* (26, 13, 17) */,
  32'h3e9d80fb /* (22, 13, 17) */,
  32'h3f0af24f /* (18, 13, 17) */,
  32'h3f0af24f /* (14, 13, 17) */,
  32'h3e9d80fb /* (10, 13, 17) */,
  32'h3e2ea39a /* (6, 13, 17) */,
  32'h3e003b1e /* (2, 13, 17) */,
  32'h3d9314c2 /* (30, 9, 17) */,
  32'h3dc42ad0 /* (26, 9, 17) */,
  32'h3e2b3653 /* (22, 9, 17) */,
  32'h3e91e4f8 /* (18, 9, 17) */,
  32'h3e91e4f8 /* (14, 9, 17) */,
  32'h3e2b3653 /* (10, 9, 17) */,
  32'h3dc42ad0 /* (6, 9, 17) */,
  32'h3d9314c2 /* (2, 9, 17) */,
  32'h3d3a7be5 /* (30, 5, 17) */,
  32'h3d73b16f /* (26, 5, 17) */,
  32'h3dce52e6 /* (22, 5, 17) */,
  32'h3e2a981c /* (18, 5, 17) */,
  32'h3e2a981c /* (14, 5, 17) */,
  32'h3dce52e6 /* (10, 5, 17) */,
  32'h3d73b16f /* (6, 5, 17) */,
  32'h3d3a7be5 /* (2, 5, 17) */,
  32'h3d1a0745 /* (30, 1, 17) */,
  32'h3d46f53f /* (26, 1, 17) */,
  32'h3da5ac70 /* (22, 1, 17) */,
  32'h3e06d8bb /* (18, 1, 17) */,
  32'h3e06d8bb /* (14, 1, 17) */,
  32'h3da5ac70 /* (10, 1, 17) */,
  32'h3d46f53f /* (6, 1, 17) */,
  32'h3d1a0745 /* (2, 1, 17) */,
  32'h3d29e985 /* (30, 29, 13) */,
  32'h3d54a03b /* (26, 29, 13) */,
  32'h3da99659 /* (22, 29, 13) */,
  32'h3e04d0b8 /* (18, 29, 13) */,
  32'h3e04d0b8 /* (14, 29, 13) */,
  32'h3da99659 /* (10, 29, 13) */,
  32'h3d54a03b /* (6, 29, 13) */,
  32'h3d29e985 /* (2, 29, 13) */,
  32'h3d6129ae /* (30, 25, 13) */,
  32'h3d90c8a7 /* (26, 25, 13) */,
  32'h3defa49b /* (22, 25, 13) */,
  32'h3e41f14c /* (18, 25, 13) */,
  32'h3e41f14c /* (14, 25, 13) */,
  32'h3defa49b /* (10, 25, 13) */,
  32'h3d90c8a7 /* (6, 25, 13) */,
  32'h3d6129ae /* (2, 25, 13) */,
  32'h3dba5db4 /* (30, 21, 13) */,
  32'h3df74dbc /* (26, 21, 13) */,
  32'h3e562fb1 /* (22, 21, 13) */,
  32'h3eb517ce /* (18, 21, 13) */,
  32'h3eb517ce /* (14, 21, 13) */,
  32'h3e562fb1 /* (10, 21, 13) */,
  32'h3df74dbc /* (6, 21, 13) */,
  32'h3dba5db4 /* (2, 21, 13) */,
  32'h3e003b1e /* (30, 17, 13) */,
  32'h3e2ea39a /* (26, 17, 13) */,
  32'h3e9d80fb /* (22, 17, 13) */,
  32'h3f0af24f /* (18, 17, 13) */,
  32'h3f0af24f /* (14, 17, 13) */,
  32'h3e9d80fb /* (10, 17, 13) */,
  32'h3e2ea39a /* (6, 17, 13) */,
  32'h3e003b1e /* (2, 17, 13) */,
  32'h3dec70da /* (30, 13, 13) */,
  32'h3e1f113d /* (26, 13, 13) */,
  32'h3e8cbae1 /* (22, 13, 13) */,
  32'h3ef33ce4 /* (18, 13, 13) */,
  32'h3ef33ce4 /* (14, 13, 13) */,
  32'h3e8cbae1 /* (10, 13, 13) */,
  32'h3e1f113d /* (6, 13, 13) */,
  32'h3dec70da /* (2, 13, 13) */,
  32'h3d8e358b /* (30, 9, 13) */,
  32'h3db9d5f4 /* (26, 9, 13) */,
  32'h3e1d56b2 /* (22, 9, 13) */,
  32'h3e821787 /* (18, 9, 13) */,
  32'h3e821787 /* (14, 9, 13) */,
  32'h3e1d56b2 /* (10, 9, 13) */,
  32'h3db9d5f4 /* (6, 9, 13) */,
  32'h3d8e358b /* (2, 9, 13) */,
  32'h3d3d84de /* (30, 5, 13) */,
  32'h3d700ffa /* (26, 5, 13) */,
  32'h3dc29629 /* (22, 5, 13) */,
  32'h3e1a8d8c /* (18, 5, 13) */,
  32'h3e1a8d8c /* (14, 5, 13) */,
  32'h3dc29629 /* (10, 5, 13) */,
  32'h3d700ffa /* (6, 5, 13) */,
  32'h3d3d84de /* (2, 5, 13) */,
  32'h3d214ba3 /* (30, 1, 13) */,
  32'h3d4876ff /* (26, 1, 13) */,
  32'h3d9e7894 /* (22, 1, 13) */,
  32'h3df65860 /* (18, 1, 13) */,
  32'h3df65860 /* (14, 1, 13) */,
  32'h3d9e7894 /* (10, 1, 13) */,
  32'h3d4876ff /* (6, 1, 13) */,
  32'h3d214ba3 /* (2, 1, 13) */,
  32'h3d12f42a /* (30, 29, 9) */,
  32'h3d215063 /* (26, 29, 9) */,
  32'h3d5dae2c /* (22, 29, 9) */,
  32'h3d9b2a7b /* (18, 29, 9) */,
  32'h3d9b2a7b /* (14, 29, 9) */,
  32'h3d5dae2c /* (10, 29, 9) */,
  32'h3d215063 /* (6, 29, 9) */,
  32'h3d12f42a /* (2, 29, 9) */,
  32'h3d26a1b5 /* (30, 25, 9) */,
  32'h3d45eb5b /* (26, 25, 9) */,
  32'h3d94014f /* (22, 25, 9) */,
  32'h3ddc09d8 /* (18, 25, 9) */,
  32'h3ddc09d8 /* (14, 25, 9) */,
  32'h3d94014f /* (10, 25, 9) */,
  32'h3d45eb5b /* (6, 25, 9) */,
  32'h3d26a1b5 /* (2, 25, 9) */,
  32'h3d6d9fa3 /* (30, 21, 9) */,
  32'h3d9750ce /* (26, 21, 9) */,
  32'h3df71c69 /* (22, 21, 9) */,
  32'h3e458f30 /* (18, 21, 9) */,
  32'h3e458f30 /* (14, 21, 9) */,
  32'h3df71c69 /* (10, 21, 9) */,
  32'h3d9750ce /* (6, 21, 9) */,
  32'h3d6d9fa3 /* (2, 21, 9) */,
  32'h3d9314c2 /* (30, 17, 9) */,
  32'h3dc42ad0 /* (26, 17, 9) */,
  32'h3e2b3653 /* (22, 17, 9) */,
  32'h3e91e4f8 /* (18, 17, 9) */,
  32'h3e91e4f8 /* (14, 17, 9) */,
  32'h3e2b3653 /* (10, 17, 9) */,
  32'h3dc42ad0 /* (6, 17, 9) */,
  32'h3d9314c2 /* (2, 17, 9) */,
  32'h3d8e358b /* (30, 13, 9) */,
  32'h3db9d5f4 /* (26, 13, 9) */,
  32'h3e1d56b2 /* (22, 13, 9) */,
  32'h3e821787 /* (18, 13, 9) */,
  32'h3e821787 /* (14, 13, 9) */,
  32'h3e1d56b2 /* (10, 13, 9) */,
  32'h3db9d5f4 /* (6, 13, 9) */,
  32'h3d8e358b /* (2, 13, 9) */,
  32'h3d42665b /* (30, 9, 9) */,
  32'h3d6fd024 /* (26, 9, 9) */,
  32'h3dbbc730 /* (22, 9, 9) */,
  32'h3e10cac5 /* (18, 9, 9) */,
  32'h3e10cac5 /* (14, 9, 9) */,
  32'h3dbbc730 /* (10, 9, 9) */,
  32'h3d6fd024 /* (6, 9, 9) */,
  32'h3d42665b /* (2, 9, 9) */,
  32'h3d18622e /* (30, 5, 9) */,
  32'h3d2db0cc /* (26, 5, 9) */,
  32'h3d781ae6 /* (22, 5, 9) */,
  32'h3db24f8e /* (18, 5, 9) */,
  32'h3db24f8e /* (14, 5, 9) */,
  32'h3d781ae6 /* (10, 5, 9) */,
  32'h3d2db0cc /* (6, 5, 9) */,
  32'h3d18622e /* (2, 5, 9) */,
  32'h3d11c69f /* (30, 1, 9) */,
  32'h3d1c53e8 /* (26, 1, 9) */,
  32'h3d52081f /* (22, 1, 9) */,
  32'h3d90dff9 /* (18, 1, 9) */,
  32'h3d90dff9 /* (14, 1, 9) */,
  32'h3d52081f /* (10, 1, 9) */,
  32'h3d1c53e8 /* (6, 1, 9) */,
  32'h3d11c69f /* (2, 1, 9) */,
  32'h3d3cd255 /* (30, 29, 5) */,
  32'h3d16d305 /* (26, 29, 5) */,
  32'h3d2344c4 /* (22, 29, 5) */,
  32'h3d487174 /* (18, 29, 5) */,
  32'h3d487174 /* (14, 29, 5) */,
  32'h3d2344c4 /* (10, 29, 5) */,
  32'h3d16d305 /* (6, 29, 5) */,
  32'h3d3cd255 /* (2, 29, 5) */,
  32'h3d14b1c0 /* (30, 25, 5) */,
  32'h3d1b2471 /* (26, 25, 5) */,
  32'h3d4b3dc7 /* (22, 25, 5) */,
  32'h3d8a0000 /* (18, 25, 5) */,
  32'h3d8a0000 /* (14, 25, 5) */,
  32'h3d4b3dc7 /* (10, 25, 5) */,
  32'h3d1b2471 /* (6, 25, 5) */,
  32'h3d14b1c0 /* (2, 25, 5) */,
  32'h3d29823f /* (30, 21, 5) */,
  32'h3d4d9045 /* (26, 21, 5) */,
  32'h3d9d9380 /* (22, 21, 5) */,
  32'h3deed79f /* (18, 21, 5) */,
  32'h3deed79f /* (14, 21, 5) */,
  32'h3d9d9380 /* (10, 21, 5) */,
  32'h3d4d9045 /* (6, 21, 5) */,
  32'h3d29823f /* (2, 21, 5) */,
  32'h3d3a7be5 /* (30, 17, 5) */,
  32'h3d73b16f /* (26, 17, 5) */,
  32'h3dce52e6 /* (22, 17, 5) */,
  32'h3e2a981c /* (18, 17, 5) */,
  32'h3e2a981c /* (14, 17, 5) */,
  32'h3dce52e6 /* (10, 17, 5) */,
  32'h3d73b16f /* (6, 17, 5) */,
  32'h3d3a7be5 /* (2, 17, 5) */,
  32'h3d3d84de /* (30, 13, 5) */,
  32'h3d700ffa /* (26, 13, 5) */,
  32'h3dc29629 /* (22, 13, 5) */,
  32'h3e1a8d8c /* (18, 13, 5) */,
  32'h3e1a8d8c /* (14, 13, 5) */,
  32'h3dc29629 /* (10, 13, 5) */,
  32'h3d700ffa /* (6, 13, 5) */,
  32'h3d3d84de /* (2, 13, 5) */,
  32'h3d18622e /* (30, 9, 5) */,
  32'h3d2db0cc /* (26, 9, 5) */,
  32'h3d781ae6 /* (22, 9, 5) */,
  32'h3db24f8e /* (18, 9, 5) */,
  32'h3db24f8e /* (14, 9, 5) */,
  32'h3d781ae6 /* (10, 9, 5) */,
  32'h3d2db0cc /* (6, 9, 5) */,
  32'h3d18622e /* (2, 9, 5) */,
  32'h3d213c91 /* (30, 5, 5) */,
  32'h3d14f7ce /* (26, 5, 5) */,
  32'h3d30fc5a /* (22, 5, 5) */,
  32'h3d63687e /* (18, 5, 5) */,
  32'h3d63687e /* (14, 5, 5) */,
  32'h3d30fc5a /* (10, 5, 5) */,
  32'h3d14f7ce /* (6, 5, 5) */,
  32'h3d213c91 /* (2, 5, 5) */,
  32'h3d59109a /* (30, 1, 5) */,
  32'h3d1a8b5a /* (26, 1, 5) */,
  32'h3d1d9589 /* (22, 1, 5) */,
  32'h3d3c7841 /* (18, 1, 5) */,
  32'h3d3c7841 /* (14, 1, 5) */,
  32'h3d1d9589 /* (10, 1, 5) */,
  32'h3d1a8b5a /* (6, 1, 5) */,
  32'h3d59109a /* (2, 1, 5) */,
  32'h3dbfa8df /* (30, 29, 1) */,
  32'h3d2ba889 /* (26, 29, 1) */,
  32'h3d14c0fd /* (22, 29, 1) */,
  32'h3d276174 /* (18, 29, 1) */,
  32'h3d276174 /* (14, 29, 1) */,
  32'h3d14c0fd /* (10, 29, 1) */,
  32'h3d2ba889 /* (6, 29, 1) */,
  32'h3dbfa8df /* (2, 29, 1) */,
  32'h3d20a35e /* (30, 25, 1) */,
  32'h3d146a43 /* (26, 25, 1) */,
  32'h3d305430 /* (22, 25, 1) */,
  32'h3d62906c /* (18, 25, 1) */,
  32'h3d62906c /* (14, 25, 1) */,
  32'h3d305430 /* (10, 25, 1) */,
  32'h3d146a43 /* (6, 25, 1) */,
  32'h3d20a35e /* (2, 25, 1) */,
  32'h3d16ed42 /* (30, 21, 1) */,
  32'h3d31191b /* (26, 21, 1) */,
  32'h3d829849 /* (22, 21, 1) */,
  32'h3dc01db4 /* (18, 21, 1) */,
  32'h3dc01db4 /* (14, 21, 1) */,
  32'h3d829849 /* (10, 21, 1) */,
  32'h3d31191b /* (6, 21, 1) */,
  32'h3d16ed42 /* (2, 21, 1) */,
  32'h3d1a0745 /* (30, 17, 1) */,
  32'h3d46f53f /* (26, 17, 1) */,
  32'h3da5ac70 /* (22, 17, 1) */,
  32'h3e06d8bb /* (18, 17, 1) */,
  32'h3e06d8bb /* (14, 17, 1) */,
  32'h3da5ac70 /* (10, 17, 1) */,
  32'h3d46f53f /* (6, 17, 1) */,
  32'h3d1a0745 /* (2, 17, 1) */,
  32'h3d214ba3 /* (30, 13, 1) */,
  32'h3d4876ff /* (26, 13, 1) */,
  32'h3d9e7894 /* (22, 13, 1) */,
  32'h3df65860 /* (18, 13, 1) */,
  32'h3df65860 /* (14, 13, 1) */,
  32'h3d9e7894 /* (10, 13, 1) */,
  32'h3d4876ff /* (6, 13, 1) */,
  32'h3d214ba3 /* (2, 13, 1) */,
  32'h3d11c69f /* (30, 9, 1) */,
  32'h3d1c53e8 /* (26, 9, 1) */,
  32'h3d52081f /* (22, 9, 1) */,
  32'h3d90dff9 /* (18, 9, 1) */,
  32'h3d90dff9 /* (14, 9, 1) */,
  32'h3d52081f /* (10, 9, 1) */,
  32'h3d1c53e8 /* (6, 9, 1) */,
  32'h3d11c69f /* (2, 9, 1) */,
  32'h3d59109a /* (30, 5, 1) */,
  32'h3d1a8b5a /* (26, 5, 1) */,
  32'h3d1d9589 /* (22, 5, 1) */,
  32'h3d3c7841 /* (18, 5, 1) */,
  32'h3d3c7841 /* (14, 5, 1) */,
  32'h3d1d9589 /* (10, 5, 1) */,
  32'h3d1a8b5a /* (6, 5, 1) */,
  32'h3d59109a /* (2, 5, 1) */,
  32'h3e4aeee2 /* (30, 1, 1) */,
  32'h3d3c9698 /* (26, 1, 1) */,
  32'h3d119771 /* (22, 1, 1) */,
  32'h3d1e0bb6 /* (18, 1, 1) */,
  32'h3d1e0bb6 /* (14, 1, 1) */,
  32'h3d119771 /* (10, 1, 1) */,
  32'h3d3c9698 /* (6, 1, 1) */,
  32'h3e4aeee2 /* (2, 1, 1) */,
  32'h3d68b01f /* (29, 29, 29) */,
  32'h3d179239 /* (25, 29, 29) */,
  32'h3d202a91 /* (21, 29, 29) */,
  32'h3d2aacf2 /* (17, 29, 29) */,
  32'h3d2fb3ed /* (13, 29, 29) */,
  32'h3d144047 /* (9, 29, 29) */,
  32'h3d314afb /* (5, 29, 29) */,
  32'h3d960c3c /* (1, 29, 29) */,
  32'h3d179239 /* (29, 25, 29) */,
  32'h3d1969a9 /* (25, 25, 29) */,
  32'h3d490aba /* (21, 25, 29) */,
  32'h3d6ce397 /* (17, 25, 29) */,
  32'h3d69f6ae /* (13, 25, 29) */,
  32'h3d2aad03 /* (9, 25, 29) */,
  32'h3d147808 /* (5, 25, 29) */,
  32'h3d1c3652 /* (1, 25, 29) */,
  32'h3d202a91 /* (29, 21, 29) */,
  32'h3d490aba /* (25, 21, 29) */,
  32'h3d9d27e1 /* (21, 21, 29) */,
  32'h3dceffa6 /* (17, 21, 29) */,
  32'h3dc2b35d /* (13, 21, 29) */,
  32'h3d767d5d /* (9, 21, 29) */,
  32'h3d2e4aa1 /* (5, 21, 29) */,
  32'h3d1a3ccf /* (1, 21, 29) */,
  32'h3d2aacf2 /* (29, 17, 29) */,
  32'h3d6ce397 /* (25, 17, 29) */,
  32'h3dceffa6 /* (21, 17, 29) */,
  32'h3e151f83 /* (17, 17, 29) */,
  32'h3e068db8 /* (13, 17, 29) */,
  32'h3d99caa3 /* (9, 17, 29) */,
  32'h3d424fe8 /* (5, 17, 29) */,
  32'h3d202be8 /* (1, 17, 29) */,
  32'h3d2fb3ed /* (29, 13, 29) */,
  32'h3d69f6ae /* (25, 13, 29) */,
  32'h3dc2b35d /* (21, 13, 29) */,
  32'h3e068db8 /* (17, 13, 29) */,
  32'h3df79892 /* (13, 13, 29) */,
  32'h3d942dc4 /* (9, 13, 29) */,
  32'h3d4466f8 /* (5, 13, 29) */,
  32'h3d269671 /* (1, 13, 29) */,
  32'h3d144047 /* (29, 9, 29) */,
  32'h3d2aad03 /* (25, 9, 29) */,
  32'h3d767d5d /* (21, 9, 29) */,
  32'h3d99caa3 /* (17, 9, 29) */,
  32'h3d942dc4 /* (13, 9, 29) */,
  32'h3d48821f /* (9, 9, 29) */,
  32'h3d1addce /* (5, 9, 29) */,
  32'h3d126006 /* (1, 9, 29) */,
  32'h3d314afb /* (29, 5, 29) */,
  32'h3d147808 /* (25, 5, 29) */,
  32'h3d2e4aa1 /* (21, 5, 29) */,
  32'h3d424fe8 /* (17, 5, 29) */,
  32'h3d4466f8 /* (13, 5, 29) */,
  32'h3d1addce /* (9, 5, 29) */,
  32'h3d1ccb4c /* (5, 5, 29) */,
  32'h3d45ae9a /* (1, 5, 29) */,
  32'h3d960c3c /* (29, 1, 29) */,
  32'h3d1c3652 /* (25, 1, 29) */,
  32'h3d1a3ccf /* (21, 1, 29) */,
  32'h3d202be8 /* (17, 1, 29) */,
  32'h3d269671 /* (13, 1, 29) */,
  32'h3d126006 /* (9, 1, 29) */,
  32'h3d45ae9a /* (5, 1, 29) */,
  32'h3deb372d /* (1, 1, 29) */,
  32'h3d179239 /* (29, 29, 25) */,
  32'h3d1969a9 /* (25, 29, 25) */,
  32'h3d490aba /* (21, 29, 25) */,
  32'h3d6ce397 /* (17, 29, 25) */,
  32'h3d69f6ae /* (13, 29, 25) */,
  32'h3d2aad03 /* (9, 29, 25) */,
  32'h3d147808 /* (5, 29, 25) */,
  32'h3d1c3652 /* (1, 29, 25) */,
  32'h3d1969a9 /* (29, 25, 25) */,
  32'h3d348078 /* (25, 25, 25) */,
  32'h3d84ce75 /* (21, 25, 25) */,
  32'h3da7bf05 /* (17, 25, 25) */,
  32'h3da0c360 /* (13, 25, 25) */,
  32'h3d563bcb /* (9, 25, 25) */,
  32'h3d21f168 /* (5, 25, 25) */,
  32'h3d167b79 /* (1, 25, 25) */,
  32'h3d490aba /* (29, 21, 25) */,
  32'h3d84ce75 /* (25, 21, 25) */,
  32'h3ddb1c7f /* (21, 21, 25) */,
  32'h3e165b49 /* (17, 21, 25) */,
  32'h3e0aca9a /* (13, 21, 25) */,
  32'h3da777c1 /* (9, 21, 25) */,
  32'h3d5ff008 /* (5, 21, 25) */,
  32'h3d3efe62 /* (1, 21, 25) */,
  32'h3d6ce397 /* (29, 17, 25) */,
  32'h3da7bf05 /* (25, 17, 25) */,
  32'h3e165b49 /* (21, 17, 25) */,
  32'h3e5db918 /* (17, 17, 25) */,
  32'h3e45db44 /* (13, 17, 25) */,
  32'h3ddc94c6 /* (9, 17, 25) */,
  32'h3d880917 /* (5, 17, 25) */,
  32'h3d5d3ed0 /* (1, 17, 25) */,
  32'h3d69f6ae /* (29, 13, 25) */,
  32'h3da0c360 /* (25, 13, 25) */,
  32'h3e0aca9a /* (21, 13, 25) */,
  32'h3e45db44 /* (17, 13, 25) */,
  32'h3e336d1b /* (13, 13, 25) */,
  32'h3dcf79e9 /* (9, 13, 25) */,
  32'h3d849ae2 /* (5, 13, 25) */,
  32'h3d5c17b6 /* (1, 13, 25) */,
  32'h3d2aad03 /* (29, 9, 25) */,
  32'h3d563bcb /* (25, 9, 25) */,
  32'h3da777c1 /* (21, 9, 25) */,
  32'h3ddc94c6 /* (17, 9, 25) */,
  32'h3dcf79e9 /* (13, 9, 25) */,
  32'h3d8354ed /* (9, 9, 25) */,
  32'h3d39ba58 /* (5, 9, 25) */,
  32'h3d245baa /* (1, 9, 25) */,
  32'h3d147808 /* (29, 5, 25) */,
  32'h3d21f168 /* (25, 5, 25) */,
  32'h3d5ff008 /* (21, 5, 25) */,
  32'h3d880917 /* (17, 5, 25) */,
  32'h3d849ae2 /* (13, 5, 25) */,
  32'h3d39ba58 /* (9, 5, 25) */,
  32'h3d170afd /* (5, 5, 25) */,
  32'h3d151e01 /* (1, 5, 25) */,
  32'h3d1c3652 /* (29, 1, 25) */,
  32'h3d167b79 /* (25, 1, 25) */,
  32'h3d3efe62 /* (21, 1, 25) */,
  32'h3d5d3ed0 /* (17, 1, 25) */,
  32'h3d5c17b6 /* (13, 1, 25) */,
  32'h3d245baa /* (9, 1, 25) */,
  32'h3d151e01 /* (5, 1, 25) */,
  32'h3d2402bf /* (1, 1, 25) */,
  32'h3d202a91 /* (29, 29, 21) */,
  32'h3d490aba /* (25, 29, 21) */,
  32'h3d9d27e1 /* (21, 29, 21) */,
  32'h3dceffa6 /* (17, 29, 21) */,
  32'h3dc2b35d /* (13, 29, 21) */,
  32'h3d767d5d /* (9, 29, 21) */,
  32'h3d2e4aa1 /* (5, 29, 21) */,
  32'h3d1a3ccf /* (1, 29, 21) */,
  32'h3d490aba /* (29, 25, 21) */,
  32'h3d84ce75 /* (25, 25, 21) */,
  32'h3ddb1c7f /* (21, 25, 21) */,
  32'h3e165b49 /* (17, 25, 21) */,
  32'h3e0aca9a /* (13, 25, 21) */,
  32'h3da777c1 /* (9, 25, 21) */,
  32'h3d5ff008 /* (5, 25, 21) */,
  32'h3d3efe62 /* (1, 25, 21) */,
  32'h3d9d27e1 /* (29, 21, 21) */,
  32'h3ddb1c7f /* (25, 21, 21) */,
  32'h3e4089a2 /* (21, 21, 21) */,
  32'h3e8b66c2 /* (17, 21, 21) */,
  32'h3e7af74d /* (13, 21, 21) */,
  32'h3e0ea5fd /* (9, 21, 21) */,
  32'h3db345e2 /* (5, 21, 21) */,
  32'h3d9352ec /* (1, 21, 21) */,
  32'h3dceffa6 /* (29, 17, 21) */,
  32'h3e165b49 /* (25, 17, 21) */,
  32'h3e8b66c2 /* (21, 17, 21) */,
  32'h3ed4648a /* (17, 17, 21) */,
  32'h3eba8e90 /* (13, 17, 21) */,
  32'h3e49046a /* (9, 17, 21) */,
  32'h3df05994 /* (5, 17, 21) */,
  32'h3dc031e4 /* (1, 17, 21) */,
  32'h3dc2b35d /* (29, 13, 21) */,
  32'h3e0aca9a /* (25, 13, 21) */,
  32'h3e7af74d /* (21, 13, 21) */,
  32'h3eba8e90 /* (17, 13, 21) */,
  32'h3ea5d30f /* (13, 13, 21) */,
  32'h3e37494b /* (9, 13, 21) */,
  32'h3de04254 /* (5, 13, 21) */,
  32'h3db58f74 /* (1, 13, 21) */,
  32'h3d767d5d /* (29, 9, 21) */,
  32'h3da777c1 /* (25, 9, 21) */,
  32'h3e0ea5fd /* (21, 9, 21) */,
  32'h3e49046a /* (17, 9, 21) */,
  32'h3e37494b /* (13, 9, 21) */,
  32'h3dd6aa1b /* (9, 9, 21) */,
  32'h3d8b02ad /* (5, 9, 21) */,
  32'h3d68852c /* (1, 9, 21) */,
  32'h3d2e4aa1 /* (29, 5, 21) */,
  32'h3d5ff008 /* (25, 5, 21) */,
  32'h3db345e2 /* (21, 5, 21) */,
  32'h3df05994 /* (17, 5, 21) */,
  32'h3de04254 /* (13, 5, 21) */,
  32'h3d8b02ad /* (9, 5, 21) */,
  32'h3d3fb488 /* (5, 5, 21) */,
  32'h3d26c9db /* (1, 5, 21) */,
  32'h3d1a3ccf /* (29, 1, 21) */,
  32'h3d3efe62 /* (25, 1, 21) */,
  32'h3d9352ec /* (21, 1, 21) */,
  32'h3dc031e4 /* (17, 1, 21) */,
  32'h3db58f74 /* (13, 1, 21) */,
  32'h3d68852c /* (9, 1, 21) */,
  32'h3d26c9db /* (5, 1, 21) */,
  32'h3d151591 /* (1, 1, 21) */,
  32'h3d2aacf2 /* (29, 29, 17) */,
  32'h3d6ce397 /* (25, 29, 17) */,
  32'h3dceffa6 /* (21, 29, 17) */,
  32'h3e151f83 /* (17, 29, 17) */,
  32'h3e068db8 /* (13, 29, 17) */,
  32'h3d99caa3 /* (9, 29, 17) */,
  32'h3d424fe8 /* (5, 29, 17) */,
  32'h3d202be8 /* (1, 29, 17) */,
  32'h3d6ce397 /* (29, 25, 17) */,
  32'h3da7bf05 /* (25, 25, 17) */,
  32'h3e165b49 /* (21, 25, 17) */,
  32'h3e5db918 /* (17, 25, 17) */,
  32'h3e45db44 /* (13, 25, 17) */,
  32'h3ddc94c6 /* (9, 25, 17) */,
  32'h3d880917 /* (5, 25, 17) */,
  32'h3d5d3ed0 /* (1, 25, 17) */,
  32'h3dceffa6 /* (29, 21, 17) */,
  32'h3e165b49 /* (25, 21, 17) */,
  32'h3e8b66c2 /* (21, 21, 17) */,
  32'h3ed4648a /* (17, 21, 17) */,
  32'h3eba8e90 /* (13, 21, 17) */,
  32'h3e49046a /* (9, 21, 17) */,
  32'h3df05994 /* (5, 21, 17) */,
  32'h3dc031e4 /* (1, 21, 17) */,
  32'h3e151f83 /* (29, 17, 17) */,
  32'h3e5db918 /* (25, 17, 17) */,
  32'h3ed4648a /* (21, 17, 17) */,
  32'h3f275a64 /* (17, 17, 17) */,
  32'h3f1092e5 /* (13, 17, 17) */,
  32'h3e969108 /* (9, 17, 17) */,
  32'h3e2edbb4 /* (5, 17, 17) */,
  32'h3e09bd27 /* (1, 17, 17) */,
  32'h3e068db8 /* (29, 13, 17) */,
  32'h3e45db44 /* (25, 13, 17) */,
  32'h3eba8e90 /* (21, 13, 17) */,
  32'h3f1092e5 /* (17, 13, 17) */,
  32'h3efbd9fe /* (13, 13, 17) */,
  32'h3e8557f4 /* (9, 13, 17) */,
  32'h3e1d0a10 /* (5, 13, 17) */,
  32'h3df92d6c /* (1, 13, 17) */,
  32'h3d99caa3 /* (29, 9, 17) */,
  32'h3ddc94c6 /* (25, 9, 17) */,
  32'h3e49046a /* (21, 9, 17) */,
  32'h3e969108 /* (17, 9, 17) */,
  32'h3e8557f4 /* (13, 9, 17) */,
  32'h3e123783 /* (9, 9, 17) */,
  32'h3db198fc /* (5, 9, 17) */,
  32'h3d8f3655 /* (1, 9, 17) */,
  32'h3d424fe8 /* (29, 5, 17) */,
  32'h3d880917 /* (25, 5, 17) */,
  32'h3df05994 /* (21, 5, 17) */,
  32'h3e2edbb4 /* (17, 5, 17) */,
  32'h3e1d0a10 /* (13, 5, 17) */,
  32'h3db198fc /* (9, 5, 17) */,
  32'h3d5e11d0 /* (5, 5, 17) */,
  32'h3d35f880 /* (1, 5, 17) */,
  32'h3d202be8 /* (29, 1, 17) */,
  32'h3d5d3ed0 /* (25, 1, 17) */,
  32'h3dc031e4 /* (21, 1, 17) */,
  32'h3e09bd27 /* (17, 1, 17) */,
  32'h3df92d6c /* (13, 1, 17) */,
  32'h3d8f3655 /* (9, 1, 17) */,
  32'h3d35f880 /* (5, 1, 17) */,
  32'h3d167d01 /* (1, 1, 17) */,
  32'h3d2fb3ed /* (29, 29, 13) */,
  32'h3d69f6ae /* (25, 29, 13) */,
  32'h3dc2b35d /* (21, 29, 13) */,
  32'h3e068db8 /* (17, 29, 13) */,
  32'h3df79892 /* (13, 29, 13) */,
  32'h3d942dc4 /* (9, 29, 13) */,
  32'h3d4466f8 /* (5, 29, 13) */,
  32'h3d269671 /* (1, 29, 13) */,
  32'h3d69f6ae /* (29, 25, 13) */,
  32'h3da0c360 /* (25, 25, 13) */,
  32'h3e0aca9a /* (21, 25, 13) */,
  32'h3e45db44 /* (17, 25, 13) */,
  32'h3e336d1b /* (13, 25, 13) */,
  32'h3dcf79e9 /* (9, 25, 13) */,
  32'h3d849ae2 /* (5, 25, 13) */,
  32'h3d5c17b6 /* (1, 25, 13) */,
  32'h3dc2b35d /* (29, 21, 13) */,
  32'h3e0aca9a /* (25, 21, 13) */,
  32'h3e7af74d /* (21, 21, 13) */,
  32'h3eba8e90 /* (17, 21, 13) */,
  32'h3ea5d30f /* (13, 21, 13) */,
  32'h3e37494b /* (9, 21, 13) */,
  32'h3de04254 /* (5, 21, 13) */,
  32'h3db58f74 /* (1, 21, 13) */,
  32'h3e068db8 /* (29, 17, 13) */,
  32'h3e45db44 /* (25, 17, 13) */,
  32'h3eba8e90 /* (21, 17, 13) */,
  32'h3f1092e5 /* (17, 17, 13) */,
  32'h3efbd9fe /* (13, 17, 13) */,
  32'h3e8557f4 /* (9, 17, 13) */,
  32'h3e1d0a10 /* (5, 17, 13) */,
  32'h3df92d6c /* (1, 17, 13) */,
  32'h3df79892 /* (29, 13, 13) */,
  32'h3e336d1b /* (25, 13, 13) */,
  32'h3ea5d30f /* (21, 13, 13) */,
  32'h3efbd9fe /* (17, 13, 13) */,
  32'h3edd8ee5 /* (13, 13, 13) */,
  32'h3e6f82ab /* (9, 13, 13) */,
  32'h3e0f99f2 /* (5, 13, 13) */,
  32'h3de602d9 /* (1, 13, 13) */,
  32'h3d942dc4 /* (29, 9, 13) */,
  32'h3dcf79e9 /* (25, 9, 13) */,
  32'h3e37494b /* (21, 9, 13) */,
  32'h3e8557f4 /* (17, 9, 13) */,
  32'h3e6f82ab /* (13, 9, 13) */,
  32'h3e076ebd /* (9, 9, 13) */,
  32'h3da95898 /* (5, 9, 13) */,
  32'h3d8ac476 /* (1, 9, 13) */,
  32'h3d4466f8 /* (29, 5, 13) */,
  32'h3d849ae2 /* (25, 5, 13) */,
  32'h3de04254 /* (21, 5, 13) */,
  32'h3e1d0a10 /* (17, 5, 13) */,
  32'h3e0f99f2 /* (13, 5, 13) */,
  32'h3da95898 /* (9, 5, 13) */,
  32'h3d5ce99d /* (5, 5, 13) */,
  32'h3d398f3f /* (1, 5, 13) */,
  32'h3d269671 /* (29, 1, 13) */,
  32'h3d5c17b6 /* (25, 1, 13) */,
  32'h3db58f74 /* (21, 1, 13) */,
  32'h3df92d6c /* (17, 1, 13) */,
  32'h3de602d9 /* (13, 1, 13) */,
  32'h3d8ac476 /* (9, 1, 13) */,
  32'h3d398f3f /* (5, 1, 13) */,
  32'h3d1e42f1 /* (1, 1, 13) */,
  32'h3d144047 /* (29, 29, 9) */,
  32'h3d2aad03 /* (25, 29, 9) */,
  32'h3d767d5d /* (21, 29, 9) */,
  32'h3d99caa3 /* (17, 29, 9) */,
  32'h3d942dc4 /* (13, 29, 9) */,
  32'h3d48821f /* (9, 29, 9) */,
  32'h3d1addce /* (5, 29, 9) */,
  32'h3d126006 /* (1, 29, 9) */,
  32'h3d2aad03 /* (29, 25, 9) */,
  32'h3d563bcb /* (25, 25, 9) */,
  32'h3da777c1 /* (21, 25, 9) */,
  32'h3ddc94c6 /* (17, 25, 9) */,
  32'h3dcf79e9 /* (13, 25, 9) */,
  32'h3d8354ed /* (9, 25, 9) */,
  32'h3d39ba58 /* (5, 25, 9) */,
  32'h3d245baa /* (1, 25, 9) */,
  32'h3d767d5d /* (29, 21, 9) */,
  32'h3da777c1 /* (25, 21, 9) */,
  32'h3e0ea5fd /* (21, 21, 9) */,
  32'h3e49046a /* (17, 21, 9) */,
  32'h3e37494b /* (13, 21, 9) */,
  32'h3dd6aa1b /* (9, 21, 9) */,
  32'h3d8b02ad /* (5, 21, 9) */,
  32'h3d68852c /* (1, 21, 9) */,
  32'h3d99caa3 /* (29, 17, 9) */,
  32'h3ddc94c6 /* (25, 17, 9) */,
  32'h3e49046a /* (21, 17, 9) */,
  32'h3e969108 /* (17, 17, 9) */,
  32'h3e8557f4 /* (13, 17, 9) */,
  32'h3e123783 /* (9, 17, 9) */,
  32'h3db198fc /* (5, 17, 9) */,
  32'h3d8f3655 /* (1, 17, 9) */,
  32'h3d942dc4 /* (29, 13, 9) */,
  32'h3dcf79e9 /* (25, 13, 9) */,
  32'h3e37494b /* (21, 13, 9) */,
  32'h3e8557f4 /* (17, 13, 9) */,
  32'h3e6f82ab /* (13, 13, 9) */,
  32'h3e076ebd /* (9, 13, 9) */,
  32'h3da95898 /* (5, 13, 9) */,
  32'h3d8ac476 /* (1, 13, 9) */,
  32'h3d48821f /* (29, 9, 9) */,
  32'h3d8354ed /* (25, 9, 9) */,
  32'h3dd6aa1b /* (21, 9, 9) */,
  32'h3e123783 /* (17, 9, 9) */,
  32'h3e076ebd /* (13, 9, 9) */,
  32'h3da4cfbf /* (9, 9, 9) */,
  32'h3d5e7d3b /* (5, 9, 9) */,
  32'h3d3ee791 /* (1, 9, 9) */,
  32'h3d1addce /* (29, 5, 9) */,
  32'h3d39ba58 /* (25, 5, 9) */,
  32'h3d8b02ad /* (21, 5, 9) */,
  32'h3db198fc /* (17, 5, 9) */,
  32'h3da95898 /* (13, 5, 9) */,
  32'h3d5e7d3b /* (9, 5, 9) */,
  32'h3d24f869 /* (5, 5, 9) */,
  32'h3d170f20 /* (1, 5, 9) */,
  32'h3d126006 /* (29, 1, 9) */,
  32'h3d245baa /* (25, 1, 9) */,
  32'h3d68852c /* (21, 1, 9) */,
  32'h3d8f3655 /* (17, 1, 9) */,
  32'h3d8ac476 /* (13, 1, 9) */,
  32'h3d3ee791 /* (9, 1, 9) */,
  32'h3d170f20 /* (5, 1, 9) */,
  32'h3d11a602 /* (1, 1, 9) */,
  32'h3d314afb /* (29, 29, 5) */,
  32'h3d147808 /* (25, 29, 5) */,
  32'h3d2e4aa1 /* (21, 29, 5) */,
  32'h3d424fe8 /* (17, 29, 5) */,
  32'h3d4466f8 /* (13, 29, 5) */,
  32'h3d1addce /* (9, 29, 5) */,
  32'h3d1ccb4c /* (5, 29, 5) */,
  32'h3d45ae9a /* (1, 29, 5) */,
  32'h3d147808 /* (29, 25, 5) */,
  32'h3d21f168 /* (25, 25, 5) */,
  32'h3d5ff008 /* (21, 25, 5) */,
  32'h3d880917 /* (17, 25, 5) */,
  32'h3d849ae2 /* (13, 25, 5) */,
  32'h3d39ba58 /* (9, 25, 5) */,
  32'h3d170afd /* (5, 25, 5) */,
  32'h3d151e01 /* (1, 25, 5) */,
  32'h3d2e4aa1 /* (29, 21, 5) */,
  32'h3d5ff008 /* (25, 21, 5) */,
  32'h3db345e2 /* (21, 21, 5) */,
  32'h3df05994 /* (17, 21, 5) */,
  32'h3de04254 /* (13, 21, 5) */,
  32'h3d8b02ad /* (9, 21, 5) */,
  32'h3d3fb488 /* (5, 21, 5) */,
  32'h3d26c9db /* (1, 21, 5) */,
  32'h3d424fe8 /* (29, 17, 5) */,
  32'h3d880917 /* (25, 17, 5) */,
  32'h3df05994 /* (21, 17, 5) */,
  32'h3e2edbb4 /* (17, 17, 5) */,
  32'h3e1d0a10 /* (13, 17, 5) */,
  32'h3db198fc /* (9, 17, 5) */,
  32'h3d5e11d0 /* (5, 17, 5) */,
  32'h3d35f880 /* (1, 17, 5) */,
  32'h3d4466f8 /* (29, 13, 5) */,
  32'h3d849ae2 /* (25, 13, 5) */,
  32'h3de04254 /* (21, 13, 5) */,
  32'h3e1d0a10 /* (17, 13, 5) */,
  32'h3e0f99f2 /* (13, 13, 5) */,
  32'h3da95898 /* (9, 13, 5) */,
  32'h3d5ce99d /* (5, 13, 5) */,
  32'h3d398f3f /* (1, 13, 5) */,
  32'h3d1addce /* (29, 9, 5) */,
  32'h3d39ba58 /* (25, 9, 5) */,
  32'h3d8b02ad /* (21, 9, 5) */,
  32'h3db198fc /* (17, 9, 5) */,
  32'h3da95898 /* (13, 9, 5) */,
  32'h3d5e7d3b /* (9, 9, 5) */,
  32'h3d24f869 /* (5, 9, 5) */,
  32'h3d170f20 /* (1, 9, 5) */,
  32'h3d1ccb4c /* (29, 5, 5) */,
  32'h3d170afd /* (25, 5, 5) */,
  32'h3d3fb488 /* (21, 5, 5) */,
  32'h3d5e11d0 /* (17, 5, 5) */,
  32'h3d5ce99d /* (13, 5, 5) */,
  32'h3d24f869 /* (9, 5, 5) */,
  32'h3d15ac37 /* (5, 5, 5) */,
  32'h3d249f29 /* (1, 5, 5) */,
  32'h3d45ae9a /* (29, 1, 5) */,
  32'h3d151e01 /* (25, 1, 5) */,
  32'h3d26c9db /* (21, 1, 5) */,
  32'h3d35f880 /* (17, 1, 5) */,
  32'h3d398f3f /* (13, 1, 5) */,
  32'h3d170f20 /* (9, 1, 5) */,
  32'h3d249f29 /* (5, 1, 5) */,
  32'h3d6890ff /* (1, 1, 5) */,
  32'h3d960c3c /* (29, 29, 1) */,
  32'h3d1c3652 /* (25, 29, 1) */,
  32'h3d1a3ccf /* (21, 29, 1) */,
  32'h3d202be8 /* (17, 29, 1) */,
  32'h3d269671 /* (13, 29, 1) */,
  32'h3d126006 /* (9, 29, 1) */,
  32'h3d45ae9a /* (5, 29, 1) */,
  32'h3deb372d /* (1, 29, 1) */,
  32'h3d1c3652 /* (29, 25, 1) */,
  32'h3d167b79 /* (25, 25, 1) */,
  32'h3d3efe62 /* (21, 25, 1) */,
  32'h3d5d3ed0 /* (17, 25, 1) */,
  32'h3d5c17b6 /* (13, 25, 1) */,
  32'h3d245baa /* (9, 25, 1) */,
  32'h3d151e01 /* (5, 25, 1) */,
  32'h3d2402bf /* (1, 25, 1) */,
  32'h3d1a3ccf /* (29, 21, 1) */,
  32'h3d3efe62 /* (25, 21, 1) */,
  32'h3d9352ec /* (21, 21, 1) */,
  32'h3dc031e4 /* (17, 21, 1) */,
  32'h3db58f74 /* (13, 21, 1) */,
  32'h3d68852c /* (9, 21, 1) */,
  32'h3d26c9db /* (5, 21, 1) */,
  32'h3d151591 /* (1, 21, 1) */,
  32'h3d202be8 /* (29, 17, 1) */,
  32'h3d5d3ed0 /* (25, 17, 1) */,
  32'h3dc031e4 /* (21, 17, 1) */,
  32'h3e09bd27 /* (17, 17, 1) */,
  32'h3df92d6c /* (13, 17, 1) */,
  32'h3d8f3655 /* (9, 17, 1) */,
  32'h3d35f880 /* (5, 17, 1) */,
  32'h3d167d01 /* (1, 17, 1) */,
  32'h3d269671 /* (29, 13, 1) */,
  32'h3d5c17b6 /* (25, 13, 1) */,
  32'h3db58f74 /* (21, 13, 1) */,
  32'h3df92d6c /* (17, 13, 1) */,
  32'h3de602d9 /* (13, 13, 1) */,
  32'h3d8ac476 /* (9, 13, 1) */,
  32'h3d398f3f /* (5, 13, 1) */,
  32'h3d1e42f1 /* (1, 13, 1) */,
  32'h3d126006 /* (29, 9, 1) */,
  32'h3d245baa /* (25, 9, 1) */,
  32'h3d68852c /* (21, 9, 1) */,
  32'h3d8f3655 /* (17, 9, 1) */,
  32'h3d8ac476 /* (13, 9, 1) */,
  32'h3d3ee791 /* (9, 9, 1) */,
  32'h3d170f20 /* (5, 9, 1) */,
  32'h3d11a602 /* (1, 9, 1) */,
  32'h3d45ae9a /* (29, 5, 1) */,
  32'h3d151e01 /* (25, 5, 1) */,
  32'h3d26c9db /* (21, 5, 1) */,
  32'h3d35f880 /* (17, 5, 1) */,
  32'h3d398f3f /* (13, 5, 1) */,
  32'h3d170f20 /* (9, 5, 1) */,
  32'h3d249f29 /* (5, 5, 1) */,
  32'h3d6890ff /* (1, 5, 1) */,
  32'h3deb372d /* (29, 1, 1) */,
  32'h3d2402bf /* (25, 1, 1) */,
  32'h3d151591 /* (21, 1, 1) */,
  32'h3d167d01 /* (17, 1, 1) */,
  32'h3d1e42f1 /* (13, 1, 1) */,
  32'h3d11a602 /* (9, 1, 1) */,
  32'h3d6890ff /* (5, 1, 1) */,
  32'h3ec3aed4 /* (1, 1, 1) */,
  32'h3d4920d0 /* (28, 29, 29) */,
  32'h3d1392fe /* (24, 29, 29) */,
  32'h3d28b308 /* (20, 29, 29) */,
  32'h3d19c07a /* (16, 29, 29) */,
  32'h3d28b308 /* (12, 29, 29) */,
  32'h3d1392fe /* (8, 29, 29) */,
  32'h3d4920d0 /* (4, 29, 29) */,
  32'h3d9c797c /* (0, 29, 29) */,
  32'h3d155fa4 /* (28, 25, 29) */,
  32'h3d2054cd /* (24, 25, 29) */,
  32'h3d5ab0e1 /* (20, 25, 29) */,
  32'h3d58de26 /* (16, 25, 29) */,
  32'h3d5ab0e1 /* (12, 25, 29) */,
  32'h3d2054cd /* (8, 25, 29) */,
  32'h3d155fa4 /* (4, 25, 29) */,
  32'h3d1cfd70 /* (0, 25, 29) */,
  32'h3d25fa09 /* (28, 21, 29) */,
  32'h3d5d0a38 /* (24, 21, 29) */,
  32'h3db0b965 /* (20, 21, 29) */,
  32'h3dc1602b /* (16, 21, 29) */,
  32'h3db0b965 /* (12, 21, 29) */,
  32'h3d5d0a38 /* (8, 21, 29) */,
  32'h3d25fa09 /* (4, 21, 29) */,
  32'h3d198ce9 /* (0, 21, 29) */,
  32'h3d349293 /* (28, 17, 29) */,
  32'h3d8608f0 /* (24, 17, 29) */,
  32'h3deea44d /* (20, 17, 29) */,
  32'h3e0de417 /* (16, 17, 29) */,
  32'h3deea44d /* (12, 17, 29) */,
  32'h3d8608f0 /* (8, 17, 29) */,
  32'h3d349293 /* (4, 17, 29) */,
  32'h3d1eeabe /* (0, 17, 29) */,
  32'h3d385879 /* (28, 13, 29) */,
  32'h3d82c188 /* (24, 13, 29) */,
  32'h3dddef48 /* (20, 13, 29) */,
  32'h3dfdd31f /* (16, 13, 29) */,
  32'h3dddef48 /* (12, 13, 29) */,
  32'h3d82c188 /* (8, 13, 29) */,
  32'h3d385879 /* (4, 13, 29) */,
  32'h3d258110 /* (0, 13, 29) */,
  32'h3d16b5b2 /* (28, 9, 29) */,
  32'h3d37919e /* (24, 9, 29) */,
  32'h3d886b82 /* (20, 9, 29) */,
  32'h3d8e3848 /* (16, 9, 29) */,
  32'h3d886b82 /* (12, 9, 29) */,
  32'h3d37919e /* (8, 9, 29) */,
  32'h3d16b5b2 /* (4, 9, 29) */,
  32'h3d1237a7 /* (0, 9, 29) */,
  32'h3d25f5ce /* (28, 5, 29) */,
  32'h3d15d660 /* (24, 5, 29) */,
  32'h3d3a4ebb /* (20, 5, 29) */,
  32'h3d3046d8 /* (16, 5, 29) */,
  32'h3d3a4ebb /* (12, 5, 29) */,
  32'h3d15d660 /* (8, 5, 29) */,
  32'h3d25f5ce /* (4, 5, 29) */,
  32'h3d490b0e /* (0, 5, 29) */,
  32'h3d6eb36b /* (28, 1, 29) */,
  32'h3d146963 /* (24, 1, 29) */,
  32'h3d210eee /* (20, 1, 29) */,
  32'h3d0fbc59 /* (16, 1, 29) */,
  32'h3d210eee /* (12, 1, 29) */,
  32'h3d146963 /* (8, 1, 29) */,
  32'h3d6eb36b /* (4, 1, 29) */,
  32'h3dff9e3f /* (0, 1, 29) */,
  32'h3d155fa4 /* (28, 29, 25) */,
  32'h3d2054cd /* (24, 29, 25) */,
  32'h3d5ab0e1 /* (20, 29, 25) */,
  32'h3d58de26 /* (16, 29, 25) */,
  32'h3d5ab0e1 /* (12, 29, 25) */,
  32'h3d2054cd /* (8, 29, 25) */,
  32'h3d155fa4 /* (4, 29, 25) */,
  32'h3d1cfd70 /* (0, 29, 25) */,
  32'h3d1cbb18 /* (28, 25, 25) */,
  32'h3d432bf1 /* (24, 25, 25) */,
  32'h3d938890 /* (20, 25, 25) */,
  32'h3d9b7830 /* (16, 25, 25) */,
  32'h3d938890 /* (12, 25, 25) */,
  32'h3d432bf1 /* (8, 25, 25) */,
  32'h3d1cbb18 /* (4, 25, 25) */,
  32'h3d162f74 /* (0, 25, 25) */,
  32'h3d52976b /* (28, 21, 25) */,
  32'h3d941bce /* (24, 21, 25) */,
  32'h3df94537 /* (20, 21, 25) */,
  32'h3e0d9cf0 /* (16, 21, 25) */,
  32'h3df94537 /* (12, 21, 25) */,
  32'h3d941bce /* (8, 21, 25) */,
  32'h3d52976b /* (4, 21, 25) */,
  32'h3d3dcd22 /* (0, 21, 25) */,
  32'h3d7b9f11 /* (28, 17, 25) */,
  32'h3dbf0444 /* (24, 17, 25) */,
  32'h3e2e6a71 /* (20, 17, 25) */,
  32'h3e540b9b /* (16, 17, 25) */,
  32'h3e2e6a71 /* (12, 17, 25) */,
  32'h3dbf0444 /* (8, 17, 25) */,
  32'h3d7b9f11 /* (4, 17, 25) */,
  32'h3d5b6048 /* (0, 17, 25) */,
  32'h3d770afc /* (28, 13, 25) */,
  32'h3db56072 /* (24, 13, 25) */,
  32'h3e1f8cbf /* (20, 13, 25) */,
  32'h3e3bd4ee /* (16, 13, 25) */,
  32'h3e1f8cbf /* (12, 13, 25) */,
  32'h3db56072 /* (8, 13, 25) */,
  32'h3d770afc /* (4, 13, 25) */,
  32'h3d5a6fdd /* (0, 13, 25) */,
  32'h3d30de15 /* (28, 9, 25) */,
  32'h3d6b8b35 /* (24, 9, 25) */,
  32'h3dbc51f9 /* (20, 9, 25) */,
  32'h3dce1075 /* (16, 9, 25) */,
  32'h3dbc51f9 /* (12, 9, 25) */,
  32'h3d6b8b35 /* (8, 9, 25) */,
  32'h3d30de15 /* (4, 9, 25) */,
  32'h3d23a039 /* (0, 9, 25) */,
  32'h3d1508af /* (28, 5, 25) */,
  32'h3d2bff3e /* (24, 5, 25) */,
  32'h3d75e4d4 /* (20, 5, 25) */,
  32'h3d7a662c /* (16, 5, 25) */,
  32'h3d75e4d4 /* (12, 5, 25) */,
  32'h3d2bff3e /* (8, 5, 25) */,
  32'h3d1508af /* (4, 5, 25) */,
  32'h3d154f7b /* (0, 5, 25) */,
  32'h3d17ff6b /* (28, 1, 25) */,
  32'h3d1bb8b6 /* (24, 1, 25) */,
  32'h3d4ea8e5 /* (20, 1, 25) */,
  32'h3d49f75a /* (16, 1, 25) */,
  32'h3d4ea8e5 /* (12, 1, 25) */,
  32'h3d1bb8b6 /* (8, 1, 25) */,
  32'h3d17ff6b /* (4, 1, 25) */,
  32'h3d25463b /* (0, 1, 25) */,
  32'h3d25fa09 /* (28, 29, 21) */,
  32'h3d5d0a38 /* (24, 29, 21) */,
  32'h3db0b965 /* (20, 29, 21) */,
  32'h3dc1602b /* (16, 29, 21) */,
  32'h3db0b965 /* (12, 29, 21) */,
  32'h3d5d0a38 /* (8, 29, 21) */,
  32'h3d25fa09 /* (4, 29, 21) */,
  32'h3d198ce9 /* (0, 29, 21) */,
  32'h3d52976b /* (28, 25, 21) */,
  32'h3d941bce /* (24, 25, 21) */,
  32'h3df94537 /* (20, 25, 21) */,
  32'h3e0d9cf0 /* (16, 25, 21) */,
  32'h3df94537 /* (12, 25, 21) */,
  32'h3d941bce /* (8, 25, 21) */,
  32'h3d52976b /* (4, 25, 21) */,
  32'h3d3dcd22 /* (0, 25, 21) */,
  32'h3da66ad4 /* (28, 21, 21) */,
  32'h3df84bb3 /* (24, 21, 21) */,
  32'h3e5e44ac /* (20, 21, 21) */,
  32'h3e84c8e0 /* (16, 21, 21) */,
  32'h3e5e44ac /* (12, 21, 21) */,
  32'h3df84bb3 /* (8, 21, 21) */,
  32'h3da66ad4 /* (4, 21, 21) */,
  32'h3d922642 /* (0, 21, 21) */,
  32'h3ddcf428 /* (28, 17, 21) */,
  32'h3e2c9c6c /* (24, 17, 21) */,
  32'h3ea31756 /* (20, 17, 21) */,
  32'h3ecca1ac /* (16, 17, 21) */,
  32'h3ea31756 /* (12, 17, 21) */,
  32'h3e2c9c6c /* (8, 17, 21) */,
  32'h3ddcf428 /* (4, 17, 21) */,
  32'h3dbe6d47 /* (0, 17, 21) */,
  32'h3dcf13a3 /* (28, 13, 21) */,
  32'h3e1e607d /* (24, 13, 21) */,
  32'h3e91dfe2 /* (20, 13, 21) */,
  32'h3eb2bd2a /* (16, 13, 21) */,
  32'h3e91dfe2 /* (12, 13, 21) */,
  32'h3e1e607d /* (8, 13, 21) */,
  32'h3dcf13a3 /* (4, 13, 21) */,
  32'h3db3fd83 /* (0, 13, 21) */,
  32'h3d81d711 /* (28, 9, 21) */,
  32'h3dbc4d73 /* (24, 9, 21) */,
  32'h3e23781b /* (20, 9, 21) */,
  32'h3e3e5da7 /* (16, 9, 21) */,
  32'h3e23781b /* (12, 9, 21) */,
  32'h3dbc4d73 /* (8, 9, 21) */,
  32'h3d81d711 /* (4, 9, 21) */,
  32'h3d66dac1 /* (0, 9, 21) */,
  32'h3d358341 /* (28, 5, 21) */,
  32'h3d77c8fd /* (24, 5, 21) */,
  32'h3dca9d53 /* (20, 5, 21) */,
  32'h3de14ffa /* (16, 5, 21) */,
  32'h3dca9d53 /* (12, 5, 21) */,
  32'h3d77c8fd /* (8, 5, 21) */,
  32'h3d358341 /* (4, 5, 21) */,
  32'h3d25e815 /* (0, 5, 21) */,
  32'h3d1f5dc3 /* (28, 1, 21) */,
  32'h3d513c3d /* (24, 1, 21) */,
  32'h3da53628 /* (20, 1, 21) */,
  32'h3db336e0 /* (16, 1, 21) */,
  32'h3da53628 /* (12, 1, 21) */,
  32'h3d513c3d /* (8, 1, 21) */,
  32'h3d1f5dc3 /* (4, 1, 21) */,
  32'h3d147e90 /* (0, 1, 21) */,
  32'h3d349293 /* (28, 29, 17) */,
  32'h3d8608f0 /* (24, 29, 17) */,
  32'h3deea44d /* (20, 29, 17) */,
  32'h3e0de417 /* (16, 29, 17) */,
  32'h3deea44d /* (12, 29, 17) */,
  32'h3d8608f0 /* (8, 29, 17) */,
  32'h3d349293 /* (4, 29, 17) */,
  32'h3d1eeabe /* (0, 29, 17) */,
  32'h3d7b9f11 /* (28, 25, 17) */,
  32'h3dbf0444 /* (24, 25, 17) */,
  32'h3e2e6a71 /* (20, 25, 17) */,
  32'h3e540b9b /* (16, 25, 17) */,
  32'h3e2e6a71 /* (12, 25, 17) */,
  32'h3dbf0444 /* (8, 25, 17) */,
  32'h3d7b9f11 /* (4, 25, 17) */,
  32'h3d5b6048 /* (0, 25, 17) */,
  32'h3ddcf428 /* (28, 21, 17) */,
  32'h3e2c9c6c /* (24, 21, 17) */,
  32'h3ea31756 /* (20, 21, 17) */,
  32'h3ecca1ac /* (16, 21, 17) */,
  32'h3ea31756 /* (12, 21, 17) */,
  32'h3e2c9c6c /* (8, 21, 17) */,
  32'h3ddcf428 /* (4, 21, 17) */,
  32'h3dbe6d47 /* (0, 21, 17) */,
  32'h3e1fe07e /* (28, 17, 17) */,
  32'h3e803f85 /* (24, 17, 17) */,
  32'h3efaa119 /* (20, 17, 17) */,
  32'h3f2286f8 /* (16, 17, 17) */,
  32'h3efaa119 /* (12, 17, 17) */,
  32'h3e803f85 /* (8, 17, 17) */,
  32'h3e1fe07e /* (4, 17, 17) */,
  32'h3e086183 /* (0, 17, 17) */,
  32'h3e0ff4ce /* (28, 13, 17) */,
  32'h3e640ba2 /* (24, 13, 17) */,
  32'h3edb3822 /* (20, 13, 17) */,
  32'h3f0bd969 /* (16, 13, 17) */,
  32'h3edb3822 /* (12, 13, 17) */,
  32'h3e640ba2 /* (8, 13, 17) */,
  32'h3e0ff4ce /* (4, 13, 17) */,
  32'h3df6cc6d /* (0, 13, 17) */,
  32'h3da3c1ed /* (28, 9, 17) */,
  32'h3dfc30a3 /* (24, 9, 17) */,
  32'h3e6a25fd /* (20, 9, 17) */,
  32'h3e908107 /* (16, 9, 17) */,
  32'h3e6a25fd /* (12, 9, 17) */,
  32'h3dfc30a3 /* (8, 9, 17) */,
  32'h3da3c1ed /* (4, 9, 17) */,
  32'h3d8df2c1 /* (0, 9, 17) */,
  32'h3d4def9b /* (28, 5, 17) */,
  32'h3d9a5b6b /* (24, 5, 17) */,
  32'h3e0ae903 /* (20, 5, 17) */,
  32'h3e26bbbb /* (16, 5, 17) */,
  32'h3e0ae903 /* (12, 5, 17) */,
  32'h3d9a5b6b /* (8, 5, 17) */,
  32'h3d4def9b /* (4, 5, 17) */,
  32'h3d347f0a /* (0, 5, 17) */,
  32'h3d294c4b /* (28, 1, 17) */,
  32'h3d7a003f /* (24, 1, 17) */,
  32'h3ddd43c2 /* (20, 1, 17) */,
  32'h3e02e976 /* (16, 1, 17) */,
  32'h3ddd43c2 /* (12, 1, 17) */,
  32'h3d7a003f /* (8, 1, 17) */,
  32'h3d294c4b /* (4, 1, 17) */,
  32'h3d155505 /* (0, 1, 17) */,
  32'h3d385879 /* (28, 29, 13) */,
  32'h3d82c188 /* (24, 29, 13) */,
  32'h3dddef48 /* (20, 29, 13) */,
  32'h3dfdd31f /* (16, 29, 13) */,
  32'h3dddef48 /* (12, 29, 13) */,
  32'h3d82c188 /* (8, 29, 13) */,
  32'h3d385879 /* (4, 29, 13) */,
  32'h3d258110 /* (0, 29, 13) */,
  32'h3d770afc /* (28, 25, 13) */,
  32'h3db56072 /* (24, 25, 13) */,
  32'h3e1f8cbf /* (20, 25, 13) */,
  32'h3e3bd4ee /* (16, 25, 13) */,
  32'h3e1f8cbf /* (12, 25, 13) */,
  32'h3db56072 /* (8, 25, 13) */,
  32'h3d770afc /* (4, 25, 13) */,
  32'h3d5a6fdd /* (0, 25, 13) */,
  32'h3dcf13a3 /* (28, 21, 13) */,
  32'h3e1e607d /* (24, 21, 13) */,
  32'h3e91dfe2 /* (20, 21, 13) */,
  32'h3eb2bd2a /* (16, 21, 13) */,
  32'h3e91dfe2 /* (12, 21, 13) */,
  32'h3e1e607d /* (8, 21, 13) */,
  32'h3dcf13a3 /* (4, 21, 13) */,
  32'h3db3fd83 /* (0, 21, 13) */,
  32'h3e0ff4ce /* (28, 17, 13) */,
  32'h3e640ba2 /* (24, 17, 13) */,
  32'h3edb3822 /* (20, 17, 13) */,
  32'h3f0bd969 /* (16, 17, 13) */,
  32'h3edb3822 /* (12, 17, 13) */,
  32'h3e640ba2 /* (8, 17, 13) */,
  32'h3e0ff4ce /* (4, 17, 13) */,
  32'h3df6cc6d /* (0, 17, 13) */,
  32'h3e0415cb /* (28, 13, 13) */,
  32'h3e4dd3dc /* (24, 13, 13) */,
  32'h3ec1d890 /* (20, 13, 13) */,
  32'h3ef27895 /* (16, 13, 13) */,
  32'h3ec1d890 /* (12, 13, 13) */,
  32'h3e4dd3dc /* (8, 13, 13) */,
  32'h3e0415cb /* (4, 13, 13) */,
  32'h3de3e928 /* (0, 13, 13) */,
  32'h3d9d0afa /* (28, 9, 13) */,
  32'h3deb6b6d /* (24, 9, 13) */,
  32'h3e53dc51 /* (20, 9, 13) */,
  32'h3e7e4b9d /* (16, 9, 13) */,
  32'h3e53dc51 /* (12, 9, 13) */,
  32'h3deb6b6d /* (8, 9, 13) */,
  32'h3d9d0afa /* (4, 9, 13) */,
  32'h3d89a49e /* (0, 9, 13) */,
  32'h3d4ea6a0 /* (28, 5, 13) */,
  32'h3d94d380 /* (24, 5, 13) */,
  32'h3e00477d /* (20, 5, 13) */,
  32'h3e1486b7 /* (16, 5, 13) */,
  32'h3e00477d /* (12, 5, 13) */,
  32'h3d94d380 /* (8, 5, 13) */,
  32'h3d4ea6a0 /* (4, 5, 13) */,
  32'h3d384488 /* (0, 5, 13) */,
  32'h3d2e802a /* (28, 1, 13) */,
  32'h3d7573b6 /* (24, 1, 13) */,
  32'h3dce8d02 /* (20, 1, 13) */,
  32'h3deaafef /* (16, 1, 13) */,
  32'h3dce8d02 /* (12, 1, 13) */,
  32'h3d7573b6 /* (8, 1, 13) */,
  32'h3d2e802a /* (4, 1, 13) */,
  32'h3d1d4601 /* (0, 1, 13) */,
  32'h3d16b5b2 /* (28, 29, 9) */,
  32'h3d37919e /* (24, 29, 9) */,
  32'h3d886b82 /* (20, 29, 9) */,
  32'h3d8e3848 /* (16, 29, 9) */,
  32'h3d886b82 /* (12, 29, 9) */,
  32'h3d37919e /* (8, 29, 9) */,
  32'h3d16b5b2 /* (4, 29, 9) */,
  32'h3d1237a7 /* (0, 29, 9) */,
  32'h3d30de15 /* (28, 25, 9) */,
  32'h3d6b8b35 /* (24, 25, 9) */,
  32'h3dbc51f9 /* (20, 25, 9) */,
  32'h3dce1075 /* (16, 25, 9) */,
  32'h3dbc51f9 /* (12, 25, 9) */,
  32'h3d6b8b35 /* (8, 25, 9) */,
  32'h3d30de15 /* (4, 25, 9) */,
  32'h3d23a039 /* (0, 25, 9) */,
  32'h3d81d711 /* (28, 21, 9) */,
  32'h3dbc4d73 /* (24, 21, 9) */,
  32'h3e23781b /* (20, 21, 9) */,
  32'h3e3e5da7 /* (16, 21, 9) */,
  32'h3e23781b /* (12, 21, 9) */,
  32'h3dbc4d73 /* (8, 21, 9) */,
  32'h3d81d711 /* (4, 21, 9) */,
  32'h3d66dac1 /* (0, 21, 9) */,
  32'h3da3c1ed /* (28, 17, 9) */,
  32'h3dfc30a3 /* (24, 17, 9) */,
  32'h3e6a25fd /* (20, 17, 9) */,
  32'h3e908107 /* (16, 17, 9) */,
  32'h3e6a25fd /* (12, 17, 9) */,
  32'h3dfc30a3 /* (8, 17, 9) */,
  32'h3da3c1ed /* (4, 17, 9) */,
  32'h3d8df2c1 /* (0, 17, 9) */,
  32'h3d9d0afa /* (28, 13, 9) */,
  32'h3deb6b6d /* (24, 13, 9) */,
  32'h3e53dc51 /* (20, 13, 9) */,
  32'h3e7e4b9d /* (16, 13, 9) */,
  32'h3e53dc51 /* (12, 13, 9) */,
  32'h3deb6b6d /* (8, 13, 9) */,
  32'h3d9d0afa /* (4, 13, 9) */,
  32'h3d89a49e /* (0, 13, 9) */,
  32'h3d51a9d2 /* (28, 9, 9) */,
  32'h3d921bde /* (24, 9, 9) */,
  32'h3df3b4f2 /* (20, 9, 9) */,
  32'h3e0981d7 /* (16, 9, 9) */,
  32'h3df3b4f2 /* (12, 9, 9) */,
  32'h3d921bde /* (8, 9, 9) */,
  32'h3d51a9d2 /* (4, 9, 9) */,
  32'h3d3dc47d /* (0, 9, 9) */,
  32'h3d1ee50b /* (28, 5, 9) */,
  32'h3d49c96c /* (24, 5, 9) */,
  32'h3d9af1c2 /* (20, 5, 9) */,
  32'h3da4f2f4 /* (16, 5, 9) */,
  32'h3d9af1c2 /* (12, 5, 9) */,
  32'h3d49c96c /* (8, 5, 9) */,
  32'h3d1ee50b /* (4, 5, 9) */,
  32'h3d16a564 /* (0, 5, 9) */,
  32'h3d13f199 /* (28, 1, 9) */,
  32'h3d2fba80 /* (24, 1, 9) */,
  32'h3d803124 /* (20, 1, 9) */,
  32'h3d8420c9 /* (16, 1, 9) */,
  32'h3d803124 /* (12, 1, 9) */,
  32'h3d2fba80 /* (8, 1, 9) */,
  32'h3d13f199 /* (4, 1, 9) */,
  32'h3d11a5c6 /* (0, 1, 9) */,
  32'h3d25f5ce /* (28, 29, 5) */,
  32'h3d15d660 /* (24, 29, 5) */,
  32'h3d3a4ebb /* (20, 29, 5) */,
  32'h3d3046d8 /* (16, 29, 5) */,
  32'h3d3a4ebb /* (12, 29, 5) */,
  32'h3d15d660 /* (8, 29, 5) */,
  32'h3d25f5ce /* (4, 29, 5) */,
  32'h3d490b0e /* (0, 29, 5) */,
  32'h3d1508af /* (28, 25, 5) */,
  32'h3d2bff3e /* (24, 25, 5) */,
  32'h3d75e4d4 /* (20, 25, 5) */,
  32'h3d7a662c /* (16, 25, 5) */,
  32'h3d75e4d4 /* (12, 25, 5) */,
  32'h3d2bff3e /* (8, 25, 5) */,
  32'h3d1508af /* (4, 25, 5) */,
  32'h3d154f7b /* (0, 25, 5) */,
  32'h3d358341 /* (28, 21, 5) */,
  32'h3d77c8fd /* (24, 21, 5) */,
  32'h3dca9d53 /* (20, 21, 5) */,
  32'h3de14ffa /* (16, 21, 5) */,
  32'h3dca9d53 /* (12, 21, 5) */,
  32'h3d77c8fd /* (8, 21, 5) */,
  32'h3d358341 /* (4, 21, 5) */,
  32'h3d25e815 /* (0, 21, 5) */,
  32'h3d4def9b /* (28, 17, 5) */,
  32'h3d9a5b6b /* (24, 17, 5) */,
  32'h3e0ae903 /* (20, 17, 5) */,
  32'h3e26bbbb /* (16, 17, 5) */,
  32'h3e0ae903 /* (12, 17, 5) */,
  32'h3d9a5b6b /* (8, 17, 5) */,
  32'h3d4def9b /* (4, 17, 5) */,
  32'h3d347f0a /* (0, 17, 5) */,
  32'h3d4ea6a0 /* (28, 13, 5) */,
  32'h3d94d380 /* (24, 13, 5) */,
  32'h3e00477d /* (20, 13, 5) */,
  32'h3e1486b7 /* (16, 13, 5) */,
  32'h3e00477d /* (12, 13, 5) */,
  32'h3d94d380 /* (8, 13, 5) */,
  32'h3d4ea6a0 /* (4, 13, 5) */,
  32'h3d384488 /* (0, 13, 5) */,
  32'h3d1ee50b /* (28, 9, 5) */,
  32'h3d49c96c /* (24, 9, 5) */,
  32'h3d9af1c2 /* (20, 9, 5) */,
  32'h3da4f2f4 /* (16, 9, 5) */,
  32'h3d9af1c2 /* (12, 9, 5) */,
  32'h3d49c96c /* (8, 9, 5) */,
  32'h3d1ee50b /* (4, 9, 5) */,
  32'h3d16a564 /* (0, 9, 5) */,
  32'h3d189061 /* (28, 5, 5) */,
  32'h3d1c4d38 /* (24, 5, 5) */,
  32'h3d4f6dfc /* (20, 5, 5) */,
  32'h3d4ab7f7 /* (16, 5, 5) */,
  32'h3d4f6dfc /* (12, 5, 5) */,
  32'h3d1c4d38 /* (8, 5, 5) */,
  32'h3d189061 /* (4, 5, 5) */,
  32'h3d25e3da /* (0, 5, 5) */,
  32'h3d334ee4 /* (28, 1, 5) */,
  32'h3d1412fd /* (24, 1, 5) */,
  32'h3d310ad3 /* (20, 1, 5) */,
  32'h3d24852f /* (16, 1, 5) */,
  32'h3d310ad3 /* (12, 1, 5) */,
  32'h3d1412fd /* (8, 1, 5) */,
  32'h3d334ee4 /* (4, 1, 5) */,
  32'h3d6e9998 /* (0, 1, 5) */,
  32'h3d6eb36b /* (28, 29, 1) */,
  32'h3d146963 /* (24, 29, 1) */,
  32'h3d210eee /* (20, 29, 1) */,
  32'h3d0fbc59 /* (16, 29, 1) */,
  32'h3d210eee /* (12, 29, 1) */,
  32'h3d146963 /* (8, 29, 1) */,
  32'h3d6eb36b /* (4, 29, 1) */,
  32'h3dff9e3f /* (0, 29, 1) */,
  32'h3d17ff6b /* (28, 25, 1) */,
  32'h3d1bb8b6 /* (24, 25, 1) */,
  32'h3d4ea8e5 /* (20, 25, 1) */,
  32'h3d49f75a /* (16, 25, 1) */,
  32'h3d4ea8e5 /* (12, 25, 1) */,
  32'h3d1bb8b6 /* (8, 25, 1) */,
  32'h3d17ff6b /* (4, 25, 1) */,
  32'h3d25463b /* (0, 25, 1) */,
  32'h3d1f5dc3 /* (28, 21, 1) */,
  32'h3d513c3d /* (24, 21, 1) */,
  32'h3da53628 /* (20, 21, 1) */,
  32'h3db336e0 /* (16, 21, 1) */,
  32'h3da53628 /* (12, 21, 1) */,
  32'h3d513c3d /* (8, 21, 1) */,
  32'h3d1f5dc3 /* (4, 21, 1) */,
  32'h3d147e90 /* (0, 21, 1) */,
  32'h3d294c4b /* (28, 17, 1) */,
  32'h3d7a003f /* (24, 17, 1) */,
  32'h3ddd43c2 /* (20, 17, 1) */,
  32'h3e02e976 /* (16, 17, 1) */,
  32'h3ddd43c2 /* (12, 17, 1) */,
  32'h3d7a003f /* (8, 17, 1) */,
  32'h3d294c4b /* (4, 17, 1) */,
  32'h3d155505 /* (0, 17, 1) */,
  32'h3d2e802a /* (28, 13, 1) */,
  32'h3d7573b6 /* (24, 13, 1) */,
  32'h3dce8d02 /* (20, 13, 1) */,
  32'h3deaafef /* (16, 13, 1) */,
  32'h3dce8d02 /* (12, 13, 1) */,
  32'h3d7573b6 /* (8, 13, 1) */,
  32'h3d2e802a /* (4, 13, 1) */,
  32'h3d1d4601 /* (0, 13, 1) */,
  32'h3d13f199 /* (28, 9, 1) */,
  32'h3d2fba80 /* (24, 9, 1) */,
  32'h3d803124 /* (20, 9, 1) */,
  32'h3d8420c9 /* (16, 9, 1) */,
  32'h3d803124 /* (12, 9, 1) */,
  32'h3d2fba80 /* (8, 9, 1) */,
  32'h3d13f199 /* (4, 9, 1) */,
  32'h3d11a5c6 /* (0, 9, 1) */,
  32'h3d334ee4 /* (28, 5, 1) */,
  32'h3d1412fd /* (24, 5, 1) */,
  32'h3d310ad3 /* (20, 5, 1) */,
  32'h3d24852f /* (16, 5, 1) */,
  32'h3d310ad3 /* (12, 5, 1) */,
  32'h3d1412fd /* (8, 5, 1) */,
  32'h3d334ee4 /* (4, 5, 1) */,
  32'h3d6e9998 /* (0, 5, 1) */,
  32'h3d9c757b /* (28, 1, 1) */,
  32'h3d1704d7 /* (24, 1, 1) */,
  32'h3d1a2df1 /* (20, 1, 1) */,
  32'h3d067e68 /* (16, 1, 1) */,
  32'h3d1a2df1 /* (12, 1, 1) */,
  32'h3d1704d7 /* (8, 1, 1) */,
  32'h3d9c757b /* (4, 1, 1) */,
  32'h3f10fe39 /* (0, 1, 1) */,
  32'h3d6eb36b /* (31, 28, 29) */,
  32'h3d25f5ce /* (27, 28, 29) */,
  32'h3d16b5b2 /* (23, 28, 29) */,
  32'h3d385879 /* (19, 28, 29) */,
  32'h3d349293 /* (15, 28, 29) */,
  32'h3d25fa09 /* (11, 28, 29) */,
  32'h3d155fa4 /* (7, 28, 29) */,
  32'h3d4920d0 /* (3, 28, 29) */,
  32'h3d146963 /* (31, 24, 29) */,
  32'h3d15d660 /* (27, 24, 29) */,
  32'h3d37919e /* (23, 24, 29) */,
  32'h3d82c188 /* (19, 24, 29) */,
  32'h3d8608f0 /* (15, 24, 29) */,
  32'h3d5d0a38 /* (11, 24, 29) */,
  32'h3d2054cd /* (7, 24, 29) */,
  32'h3d1392fe /* (3, 24, 29) */,
  32'h3d210eee /* (31, 20, 29) */,
  32'h3d3a4ebb /* (27, 20, 29) */,
  32'h3d886b82 /* (23, 20, 29) */,
  32'h3dddef48 /* (19, 20, 29) */,
  32'h3deea44d /* (15, 20, 29) */,
  32'h3db0b965 /* (11, 20, 29) */,
  32'h3d5ab0e1 /* (7, 20, 29) */,
  32'h3d28b308 /* (3, 20, 29) */,
  32'h3d0fbc59 /* (31, 16, 29) */,
  32'h3d3046d8 /* (27, 16, 29) */,
  32'h3d8e3848 /* (23, 16, 29) */,
  32'h3dfdd31f /* (19, 16, 29) */,
  32'h3e0de417 /* (15, 16, 29) */,
  32'h3dc1602b /* (11, 16, 29) */,
  32'h3d58de26 /* (7, 16, 29) */,
  32'h3d19c07a /* (3, 16, 29) */,
  32'h3d210eee /* (31, 12, 29) */,
  32'h3d3a4ebb /* (27, 12, 29) */,
  32'h3d886b82 /* (23, 12, 29) */,
  32'h3dddef48 /* (19, 12, 29) */,
  32'h3deea44d /* (15, 12, 29) */,
  32'h3db0b965 /* (11, 12, 29) */,
  32'h3d5ab0e1 /* (7, 12, 29) */,
  32'h3d28b308 /* (3, 12, 29) */,
  32'h3d146963 /* (31, 8, 29) */,
  32'h3d15d660 /* (27, 8, 29) */,
  32'h3d37919e /* (23, 8, 29) */,
  32'h3d82c188 /* (19, 8, 29) */,
  32'h3d8608f0 /* (15, 8, 29) */,
  32'h3d5d0a38 /* (11, 8, 29) */,
  32'h3d2054cd /* (7, 8, 29) */,
  32'h3d1392fe /* (3, 8, 29) */,
  32'h3d6eb36b /* (31, 4, 29) */,
  32'h3d25f5ce /* (27, 4, 29) */,
  32'h3d16b5b2 /* (23, 4, 29) */,
  32'h3d385879 /* (19, 4, 29) */,
  32'h3d349293 /* (15, 4, 29) */,
  32'h3d25fa09 /* (11, 4, 29) */,
  32'h3d155fa4 /* (7, 4, 29) */,
  32'h3d4920d0 /* (3, 4, 29) */,
  32'h3dff9e3f /* (31, 0, 29) */,
  32'h3d490b0e /* (27, 0, 29) */,
  32'h3d1237a7 /* (23, 0, 29) */,
  32'h3d258110 /* (19, 0, 29) */,
  32'h3d1eeabe /* (15, 0, 29) */,
  32'h3d198ce9 /* (11, 0, 29) */,
  32'h3d1cfd70 /* (7, 0, 29) */,
  32'h3d9c797c /* (3, 0, 29) */,
  32'h3d17ff6b /* (31, 28, 25) */,
  32'h3d1508af /* (27, 28, 25) */,
  32'h3d30de15 /* (23, 28, 25) */,
  32'h3d770afc /* (19, 28, 25) */,
  32'h3d7b9f11 /* (15, 28, 25) */,
  32'h3d52976b /* (11, 28, 25) */,
  32'h3d1cbb18 /* (7, 28, 25) */,
  32'h3d155fa4 /* (3, 28, 25) */,
  32'h3d1bb8b6 /* (31, 24, 25) */,
  32'h3d2bff3e /* (27, 24, 25) */,
  32'h3d6b8b35 /* (23, 24, 25) */,
  32'h3db56072 /* (19, 24, 25) */,
  32'h3dbf0444 /* (15, 24, 25) */,
  32'h3d941bce /* (11, 24, 25) */,
  32'h3d432bf1 /* (7, 24, 25) */,
  32'h3d2054cd /* (3, 24, 25) */,
  32'h3d4ea8e5 /* (31, 20, 25) */,
  32'h3d75e4d4 /* (27, 20, 25) */,
  32'h3dbc51f9 /* (23, 20, 25) */,
  32'h3e1f8cbf /* (19, 20, 25) */,
  32'h3e2e6a71 /* (15, 20, 25) */,
  32'h3df94537 /* (11, 20, 25) */,
  32'h3d938890 /* (7, 20, 25) */,
  32'h3d5ab0e1 /* (3, 20, 25) */,
  32'h3d49f75a /* (31, 16, 25) */,
  32'h3d7a662c /* (27, 16, 25) */,
  32'h3dce1075 /* (23, 16, 25) */,
  32'h3e3bd4ee /* (19, 16, 25) */,
  32'h3e540b9b /* (15, 16, 25) */,
  32'h3e0d9cf0 /* (11, 16, 25) */,
  32'h3d9b7830 /* (7, 16, 25) */,
  32'h3d58de26 /* (3, 16, 25) */,
  32'h3d4ea8e5 /* (31, 12, 25) */,
  32'h3d75e4d4 /* (27, 12, 25) */,
  32'h3dbc51f9 /* (23, 12, 25) */,
  32'h3e1f8cbf /* (19, 12, 25) */,
  32'h3e2e6a71 /* (15, 12, 25) */,
  32'h3df94537 /* (11, 12, 25) */,
  32'h3d938890 /* (7, 12, 25) */,
  32'h3d5ab0e1 /* (3, 12, 25) */,
  32'h3d1bb8b6 /* (31, 8, 25) */,
  32'h3d2bff3e /* (27, 8, 25) */,
  32'h3d6b8b35 /* (23, 8, 25) */,
  32'h3db56072 /* (19, 8, 25) */,
  32'h3dbf0444 /* (15, 8, 25) */,
  32'h3d941bce /* (11, 8, 25) */,
  32'h3d432bf1 /* (7, 8, 25) */,
  32'h3d2054cd /* (3, 8, 25) */,
  32'h3d17ff6b /* (31, 4, 25) */,
  32'h3d1508af /* (27, 4, 25) */,
  32'h3d30de15 /* (23, 4, 25) */,
  32'h3d770afc /* (19, 4, 25) */,
  32'h3d7b9f11 /* (15, 4, 25) */,
  32'h3d52976b /* (11, 4, 25) */,
  32'h3d1cbb18 /* (7, 4, 25) */,
  32'h3d155fa4 /* (3, 4, 25) */,
  32'h3d25463b /* (31, 0, 25) */,
  32'h3d154f7b /* (27, 0, 25) */,
  32'h3d23a039 /* (23, 0, 25) */,
  32'h3d5a6fdd /* (19, 0, 25) */,
  32'h3d5b6048 /* (15, 0, 25) */,
  32'h3d3dcd22 /* (11, 0, 25) */,
  32'h3d162f74 /* (7, 0, 25) */,
  32'h3d1cfd70 /* (3, 0, 25) */,
  32'h3d1f5dc3 /* (31, 28, 21) */,
  32'h3d358341 /* (27, 28, 21) */,
  32'h3d81d711 /* (23, 28, 21) */,
  32'h3dcf13a3 /* (19, 28, 21) */,
  32'h3ddcf428 /* (15, 28, 21) */,
  32'h3da66ad4 /* (11, 28, 21) */,
  32'h3d52976b /* (7, 28, 21) */,
  32'h3d25fa09 /* (3, 28, 21) */,
  32'h3d513c3d /* (31, 24, 21) */,
  32'h3d77c8fd /* (27, 24, 21) */,
  32'h3dbc4d73 /* (23, 24, 21) */,
  32'h3e1e607d /* (19, 24, 21) */,
  32'h3e2c9c6c /* (15, 24, 21) */,
  32'h3df84bb3 /* (11, 24, 21) */,
  32'h3d941bce /* (7, 24, 21) */,
  32'h3d5d0a38 /* (3, 24, 21) */,
  32'h3da53628 /* (31, 20, 21) */,
  32'h3dca9d53 /* (27, 20, 21) */,
  32'h3e23781b /* (23, 20, 21) */,
  32'h3e91dfe2 /* (19, 20, 21) */,
  32'h3ea31756 /* (15, 20, 21) */,
  32'h3e5e44ac /* (11, 20, 21) */,
  32'h3df94537 /* (7, 20, 21) */,
  32'h3db0b965 /* (3, 20, 21) */,
  32'h3db336e0 /* (31, 16, 21) */,
  32'h3de14ffa /* (27, 16, 21) */,
  32'h3e3e5da7 /* (23, 16, 21) */,
  32'h3eb2bd2a /* (19, 16, 21) */,
  32'h3ecca1ac /* (15, 16, 21) */,
  32'h3e84c8e0 /* (11, 16, 21) */,
  32'h3e0d9cf0 /* (7, 16, 21) */,
  32'h3dc1602b /* (3, 16, 21) */,
  32'h3da53628 /* (31, 12, 21) */,
  32'h3dca9d53 /* (27, 12, 21) */,
  32'h3e23781b /* (23, 12, 21) */,
  32'h3e91dfe2 /* (19, 12, 21) */,
  32'h3ea31756 /* (15, 12, 21) */,
  32'h3e5e44ac /* (11, 12, 21) */,
  32'h3df94537 /* (7, 12, 21) */,
  32'h3db0b965 /* (3, 12, 21) */,
  32'h3d513c3d /* (31, 8, 21) */,
  32'h3d77c8fd /* (27, 8, 21) */,
  32'h3dbc4d73 /* (23, 8, 21) */,
  32'h3e1e607d /* (19, 8, 21) */,
  32'h3e2c9c6c /* (15, 8, 21) */,
  32'h3df84bb3 /* (11, 8, 21) */,
  32'h3d941bce /* (7, 8, 21) */,
  32'h3d5d0a38 /* (3, 8, 21) */,
  32'h3d1f5dc3 /* (31, 4, 21) */,
  32'h3d358341 /* (27, 4, 21) */,
  32'h3d81d711 /* (23, 4, 21) */,
  32'h3dcf13a3 /* (19, 4, 21) */,
  32'h3ddcf428 /* (15, 4, 21) */,
  32'h3da66ad4 /* (11, 4, 21) */,
  32'h3d52976b /* (7, 4, 21) */,
  32'h3d25fa09 /* (3, 4, 21) */,
  32'h3d147e90 /* (31, 0, 21) */,
  32'h3d25e815 /* (27, 0, 21) */,
  32'h3d66dac1 /* (23, 0, 21) */,
  32'h3db3fd83 /* (19, 0, 21) */,
  32'h3dbe6d47 /* (15, 0, 21) */,
  32'h3d922642 /* (11, 0, 21) */,
  32'h3d3dcd22 /* (7, 0, 21) */,
  32'h3d198ce9 /* (3, 0, 21) */,
  32'h3d294c4b /* (31, 28, 17) */,
  32'h3d4def9b /* (27, 28, 17) */,
  32'h3da3c1ed /* (23, 28, 17) */,
  32'h3e0ff4ce /* (19, 28, 17) */,
  32'h3e1fe07e /* (15, 28, 17) */,
  32'h3ddcf428 /* (11, 28, 17) */,
  32'h3d7b9f11 /* (7, 28, 17) */,
  32'h3d349293 /* (3, 28, 17) */,
  32'h3d7a003f /* (31, 24, 17) */,
  32'h3d9a5b6b /* (27, 24, 17) */,
  32'h3dfc30a3 /* (23, 24, 17) */,
  32'h3e640ba2 /* (19, 24, 17) */,
  32'h3e803f85 /* (15, 24, 17) */,
  32'h3e2c9c6c /* (11, 24, 17) */,
  32'h3dbf0444 /* (7, 24, 17) */,
  32'h3d8608f0 /* (3, 24, 17) */,
  32'h3ddd43c2 /* (31, 20, 17) */,
  32'h3e0ae903 /* (27, 20, 17) */,
  32'h3e6a25fd /* (23, 20, 17) */,
  32'h3edb3822 /* (19, 20, 17) */,
  32'h3efaa119 /* (15, 20, 17) */,
  32'h3ea31756 /* (11, 20, 17) */,
  32'h3e2e6a71 /* (7, 20, 17) */,
  32'h3deea44d /* (3, 20, 17) */,
  32'h3e02e976 /* (31, 16, 17) */,
  32'h3e26bbbb /* (27, 16, 17) */,
  32'h3e908107 /* (23, 16, 17) */,
  32'h3f0bd969 /* (19, 16, 17) */,
  32'h3f2286f8 /* (15, 16, 17) */,
  32'h3ecca1ac /* (11, 16, 17) */,
  32'h3e540b9b /* (7, 16, 17) */,
  32'h3e0de417 /* (3, 16, 17) */,
  32'h3ddd43c2 /* (31, 12, 17) */,
  32'h3e0ae903 /* (27, 12, 17) */,
  32'h3e6a25fd /* (23, 12, 17) */,
  32'h3edb3822 /* (19, 12, 17) */,
  32'h3efaa119 /* (15, 12, 17) */,
  32'h3ea31756 /* (11, 12, 17) */,
  32'h3e2e6a71 /* (7, 12, 17) */,
  32'h3deea44d /* (3, 12, 17) */,
  32'h3d7a003f /* (31, 8, 17) */,
  32'h3d9a5b6b /* (27, 8, 17) */,
  32'h3dfc30a3 /* (23, 8, 17) */,
  32'h3e640ba2 /* (19, 8, 17) */,
  32'h3e803f85 /* (15, 8, 17) */,
  32'h3e2c9c6c /* (11, 8, 17) */,
  32'h3dbf0444 /* (7, 8, 17) */,
  32'h3d8608f0 /* (3, 8, 17) */,
  32'h3d294c4b /* (31, 4, 17) */,
  32'h3d4def9b /* (27, 4, 17) */,
  32'h3da3c1ed /* (23, 4, 17) */,
  32'h3e0ff4ce /* (19, 4, 17) */,
  32'h3e1fe07e /* (15, 4, 17) */,
  32'h3ddcf428 /* (11, 4, 17) */,
  32'h3d7b9f11 /* (7, 4, 17) */,
  32'h3d349293 /* (3, 4, 17) */,
  32'h3d155505 /* (31, 0, 17) */,
  32'h3d347f0a /* (27, 0, 17) */,
  32'h3d8df2c1 /* (23, 0, 17) */,
  32'h3df6cc6d /* (19, 0, 17) */,
  32'h3e086183 /* (15, 0, 17) */,
  32'h3dbe6d47 /* (11, 0, 17) */,
  32'h3d5b6048 /* (7, 0, 17) */,
  32'h3d1eeabe /* (3, 0, 17) */,
  32'h3d2e802a /* (31, 28, 13) */,
  32'h3d4ea6a0 /* (27, 28, 13) */,
  32'h3d9d0afa /* (23, 28, 13) */,
  32'h3e0415cb /* (19, 28, 13) */,
  32'h3e0ff4ce /* (15, 28, 13) */,
  32'h3dcf13a3 /* (11, 28, 13) */,
  32'h3d770afc /* (7, 28, 13) */,
  32'h3d385879 /* (3, 28, 13) */,
  32'h3d7573b6 /* (31, 24, 13) */,
  32'h3d94d380 /* (27, 24, 13) */,
  32'h3deb6b6d /* (23, 24, 13) */,
  32'h3e4dd3dc /* (19, 24, 13) */,
  32'h3e640ba2 /* (15, 24, 13) */,
  32'h3e1e607d /* (11, 24, 13) */,
  32'h3db56072 /* (7, 24, 13) */,
  32'h3d82c188 /* (3, 24, 13) */,
  32'h3dce8d02 /* (31, 20, 13) */,
  32'h3e00477d /* (27, 20, 13) */,
  32'h3e53dc51 /* (23, 20, 13) */,
  32'h3ec1d890 /* (19, 20, 13) */,
  32'h3edb3822 /* (15, 20, 13) */,
  32'h3e91dfe2 /* (11, 20, 13) */,
  32'h3e1f8cbf /* (7, 20, 13) */,
  32'h3dddef48 /* (3, 20, 13) */,
  32'h3deaafef /* (31, 16, 13) */,
  32'h3e1486b7 /* (27, 16, 13) */,
  32'h3e7e4b9d /* (23, 16, 13) */,
  32'h3ef27895 /* (19, 16, 13) */,
  32'h3f0bd969 /* (15, 16, 13) */,
  32'h3eb2bd2a /* (11, 16, 13) */,
  32'h3e3bd4ee /* (7, 16, 13) */,
  32'h3dfdd31f /* (3, 16, 13) */,
  32'h3dce8d02 /* (31, 12, 13) */,
  32'h3e00477d /* (27, 12, 13) */,
  32'h3e53dc51 /* (23, 12, 13) */,
  32'h3ec1d890 /* (19, 12, 13) */,
  32'h3edb3822 /* (15, 12, 13) */,
  32'h3e91dfe2 /* (11, 12, 13) */,
  32'h3e1f8cbf /* (7, 12, 13) */,
  32'h3dddef48 /* (3, 12, 13) */,
  32'h3d7573b6 /* (31, 8, 13) */,
  32'h3d94d380 /* (27, 8, 13) */,
  32'h3deb6b6d /* (23, 8, 13) */,
  32'h3e4dd3dc /* (19, 8, 13) */,
  32'h3e640ba2 /* (15, 8, 13) */,
  32'h3e1e607d /* (11, 8, 13) */,
  32'h3db56072 /* (7, 8, 13) */,
  32'h3d82c188 /* (3, 8, 13) */,
  32'h3d2e802a /* (31, 4, 13) */,
  32'h3d4ea6a0 /* (27, 4, 13) */,
  32'h3d9d0afa /* (23, 4, 13) */,
  32'h3e0415cb /* (19, 4, 13) */,
  32'h3e0ff4ce /* (15, 4, 13) */,
  32'h3dcf13a3 /* (11, 4, 13) */,
  32'h3d770afc /* (7, 4, 13) */,
  32'h3d385879 /* (3, 4, 13) */,
  32'h3d1d4601 /* (31, 0, 13) */,
  32'h3d384488 /* (27, 0, 13) */,
  32'h3d89a49e /* (23, 0, 13) */,
  32'h3de3e928 /* (19, 0, 13) */,
  32'h3df6cc6d /* (15, 0, 13) */,
  32'h3db3fd83 /* (11, 0, 13) */,
  32'h3d5a6fdd /* (7, 0, 13) */,
  32'h3d258110 /* (3, 0, 13) */,
  32'h3d13f199 /* (31, 28, 9) */,
  32'h3d1ee50b /* (27, 28, 9) */,
  32'h3d51a9d2 /* (23, 28, 9) */,
  32'h3d9d0afa /* (19, 28, 9) */,
  32'h3da3c1ed /* (15, 28, 9) */,
  32'h3d81d711 /* (11, 28, 9) */,
  32'h3d30de15 /* (7, 28, 9) */,
  32'h3d16b5b2 /* (3, 28, 9) */,
  32'h3d2fba80 /* (31, 24, 9) */,
  32'h3d49c96c /* (27, 24, 9) */,
  32'h3d921bde /* (23, 24, 9) */,
  32'h3deb6b6d /* (19, 24, 9) */,
  32'h3dfc30a3 /* (15, 24, 9) */,
  32'h3dbc4d73 /* (11, 24, 9) */,
  32'h3d6b8b35 /* (7, 24, 9) */,
  32'h3d37919e /* (3, 24, 9) */,
  32'h3d803124 /* (31, 20, 9) */,
  32'h3d9af1c2 /* (27, 20, 9) */,
  32'h3df3b4f2 /* (23, 20, 9) */,
  32'h3e53dc51 /* (19, 20, 9) */,
  32'h3e6a25fd /* (15, 20, 9) */,
  32'h3e23781b /* (11, 20, 9) */,
  32'h3dbc51f9 /* (7, 20, 9) */,
  32'h3d886b82 /* (3, 20, 9) */,
  32'h3d8420c9 /* (31, 16, 9) */,
  32'h3da4f2f4 /* (27, 16, 9) */,
  32'h3e0981d7 /* (23, 16, 9) */,
  32'h3e7e4b9d /* (19, 16, 9) */,
  32'h3e908107 /* (15, 16, 9) */,
  32'h3e3e5da7 /* (11, 16, 9) */,
  32'h3dce1075 /* (7, 16, 9) */,
  32'h3d8e3848 /* (3, 16, 9) */,
  32'h3d803124 /* (31, 12, 9) */,
  32'h3d9af1c2 /* (27, 12, 9) */,
  32'h3df3b4f2 /* (23, 12, 9) */,
  32'h3e53dc51 /* (19, 12, 9) */,
  32'h3e6a25fd /* (15, 12, 9) */,
  32'h3e23781b /* (11, 12, 9) */,
  32'h3dbc51f9 /* (7, 12, 9) */,
  32'h3d886b82 /* (3, 12, 9) */,
  32'h3d2fba80 /* (31, 8, 9) */,
  32'h3d49c96c /* (27, 8, 9) */,
  32'h3d921bde /* (23, 8, 9) */,
  32'h3deb6b6d /* (19, 8, 9) */,
  32'h3dfc30a3 /* (15, 8, 9) */,
  32'h3dbc4d73 /* (11, 8, 9) */,
  32'h3d6b8b35 /* (7, 8, 9) */,
  32'h3d37919e /* (3, 8, 9) */,
  32'h3d13f199 /* (31, 4, 9) */,
  32'h3d1ee50b /* (27, 4, 9) */,
  32'h3d51a9d2 /* (23, 4, 9) */,
  32'h3d9d0afa /* (19, 4, 9) */,
  32'h3da3c1ed /* (15, 4, 9) */,
  32'h3d81d711 /* (11, 4, 9) */,
  32'h3d30de15 /* (7, 4, 9) */,
  32'h3d16b5b2 /* (3, 4, 9) */,
  32'h3d11a5c6 /* (31, 0, 9) */,
  32'h3d16a564 /* (27, 0, 9) */,
  32'h3d3dc47d /* (23, 0, 9) */,
  32'h3d89a49e /* (19, 0, 9) */,
  32'h3d8df2c1 /* (15, 0, 9) */,
  32'h3d66dac1 /* (11, 0, 9) */,
  32'h3d23a039 /* (7, 0, 9) */,
  32'h3d1237a7 /* (3, 0, 9) */,
  32'h3d334ee4 /* (31, 28, 5) */,
  32'h3d189061 /* (27, 28, 5) */,
  32'h3d1ee50b /* (23, 28, 5) */,
  32'h3d4ea6a0 /* (19, 28, 5) */,
  32'h3d4def9b /* (15, 28, 5) */,
  32'h3d358341 /* (11, 28, 5) */,
  32'h3d1508af /* (7, 28, 5) */,
  32'h3d25f5ce /* (3, 28, 5) */,
  32'h3d1412fd /* (31, 24, 5) */,
  32'h3d1c4d38 /* (27, 24, 5) */,
  32'h3d49c96c /* (23, 24, 5) */,
  32'h3d94d380 /* (19, 24, 5) */,
  32'h3d9a5b6b /* (15, 24, 5) */,
  32'h3d77c8fd /* (11, 24, 5) */,
  32'h3d2bff3e /* (7, 24, 5) */,
  32'h3d15d660 /* (3, 24, 5) */,
  32'h3d310ad3 /* (31, 20, 5) */,
  32'h3d4f6dfc /* (27, 20, 5) */,
  32'h3d9af1c2 /* (23, 20, 5) */,
  32'h3e00477d /* (19, 20, 5) */,
  32'h3e0ae903 /* (15, 20, 5) */,
  32'h3dca9d53 /* (11, 20, 5) */,
  32'h3d75e4d4 /* (7, 20, 5) */,
  32'h3d3a4ebb /* (3, 20, 5) */,
  32'h3d24852f /* (31, 16, 5) */,
  32'h3d4ab7f7 /* (27, 16, 5) */,
  32'h3da4f2f4 /* (23, 16, 5) */,
  32'h3e1486b7 /* (19, 16, 5) */,
  32'h3e26bbbb /* (15, 16, 5) */,
  32'h3de14ffa /* (11, 16, 5) */,
  32'h3d7a662c /* (7, 16, 5) */,
  32'h3d3046d8 /* (3, 16, 5) */,
  32'h3d310ad3 /* (31, 12, 5) */,
  32'h3d4f6dfc /* (27, 12, 5) */,
  32'h3d9af1c2 /* (23, 12, 5) */,
  32'h3e00477d /* (19, 12, 5) */,
  32'h3e0ae903 /* (15, 12, 5) */,
  32'h3dca9d53 /* (11, 12, 5) */,
  32'h3d75e4d4 /* (7, 12, 5) */,
  32'h3d3a4ebb /* (3, 12, 5) */,
  32'h3d1412fd /* (31, 8, 5) */,
  32'h3d1c4d38 /* (27, 8, 5) */,
  32'h3d49c96c /* (23, 8, 5) */,
  32'h3d94d380 /* (19, 8, 5) */,
  32'h3d9a5b6b /* (15, 8, 5) */,
  32'h3d77c8fd /* (11, 8, 5) */,
  32'h3d2bff3e /* (7, 8, 5) */,
  32'h3d15d660 /* (3, 8, 5) */,
  32'h3d334ee4 /* (31, 4, 5) */,
  32'h3d189061 /* (27, 4, 5) */,
  32'h3d1ee50b /* (23, 4, 5) */,
  32'h3d4ea6a0 /* (19, 4, 5) */,
  32'h3d4def9b /* (15, 4, 5) */,
  32'h3d358341 /* (11, 4, 5) */,
  32'h3d1508af /* (7, 4, 5) */,
  32'h3d25f5ce /* (3, 4, 5) */,
  32'h3d6e9998 /* (31, 0, 5) */,
  32'h3d25e3da /* (27, 0, 5) */,
  32'h3d16a564 /* (23, 0, 5) */,
  32'h3d384488 /* (19, 0, 5) */,
  32'h3d347f0a /* (15, 0, 5) */,
  32'h3d25e815 /* (11, 0, 5) */,
  32'h3d154f7b /* (7, 0, 5) */,
  32'h3d490b0e /* (3, 0, 5) */,
  32'h3d9c757b /* (31, 28, 1) */,
  32'h3d334ee4 /* (27, 28, 1) */,
  32'h3d13f199 /* (23, 28, 1) */,
  32'h3d2e802a /* (19, 28, 1) */,
  32'h3d294c4b /* (15, 28, 1) */,
  32'h3d1f5dc3 /* (11, 28, 1) */,
  32'h3d17ff6b /* (7, 28, 1) */,
  32'h3d6eb36b /* (3, 28, 1) */,
  32'h3d1704d7 /* (31, 24, 1) */,
  32'h3d1412fd /* (27, 24, 1) */,
  32'h3d2fba80 /* (23, 24, 1) */,
  32'h3d7573b6 /* (19, 24, 1) */,
  32'h3d7a003f /* (15, 24, 1) */,
  32'h3d513c3d /* (11, 24, 1) */,
  32'h3d1bb8b6 /* (7, 24, 1) */,
  32'h3d146963 /* (3, 24, 1) */,
  32'h3d1a2df1 /* (31, 20, 1) */,
  32'h3d310ad3 /* (27, 20, 1) */,
  32'h3d803124 /* (23, 20, 1) */,
  32'h3dce8d02 /* (19, 20, 1) */,
  32'h3ddd43c2 /* (15, 20, 1) */,
  32'h3da53628 /* (11, 20, 1) */,
  32'h3d4ea8e5 /* (7, 20, 1) */,
  32'h3d210eee /* (3, 20, 1) */,
  32'h3d067e68 /* (31, 16, 1) */,
  32'h3d24852f /* (27, 16, 1) */,
  32'h3d8420c9 /* (23, 16, 1) */,
  32'h3deaafef /* (19, 16, 1) */,
  32'h3e02e976 /* (15, 16, 1) */,
  32'h3db336e0 /* (11, 16, 1) */,
  32'h3d49f75a /* (7, 16, 1) */,
  32'h3d0fbc59 /* (3, 16, 1) */,
  32'h3d1a2df1 /* (31, 12, 1) */,
  32'h3d310ad3 /* (27, 12, 1) */,
  32'h3d803124 /* (23, 12, 1) */,
  32'h3dce8d02 /* (19, 12, 1) */,
  32'h3ddd43c2 /* (15, 12, 1) */,
  32'h3da53628 /* (11, 12, 1) */,
  32'h3d4ea8e5 /* (7, 12, 1) */,
  32'h3d210eee /* (3, 12, 1) */,
  32'h3d1704d7 /* (31, 8, 1) */,
  32'h3d1412fd /* (27, 8, 1) */,
  32'h3d2fba80 /* (23, 8, 1) */,
  32'h3d7573b6 /* (19, 8, 1) */,
  32'h3d7a003f /* (15, 8, 1) */,
  32'h3d513c3d /* (11, 8, 1) */,
  32'h3d1bb8b6 /* (7, 8, 1) */,
  32'h3d146963 /* (3, 8, 1) */,
  32'h3d9c757b /* (31, 4, 1) */,
  32'h3d334ee4 /* (27, 4, 1) */,
  32'h3d13f199 /* (23, 4, 1) */,
  32'h3d2e802a /* (19, 4, 1) */,
  32'h3d294c4b /* (15, 4, 1) */,
  32'h3d1f5dc3 /* (11, 4, 1) */,
  32'h3d17ff6b /* (7, 4, 1) */,
  32'h3d6eb36b /* (3, 4, 1) */,
  32'h3f10fe39 /* (31, 0, 1) */,
  32'h3d6e9998 /* (27, 0, 1) */,
  32'h3d11a5c6 /* (23, 0, 1) */,
  32'h3d1d4601 /* (19, 0, 1) */,
  32'h3d155505 /* (15, 0, 1) */,
  32'h3d147e90 /* (11, 0, 1) */,
  32'h3d25463b /* (7, 0, 1) */,
  32'h3dff9e3f /* (3, 0, 1) */,
  32'h3d5defd3 /* (30, 28, 29) */,
  32'h3d1b3fff /* (26, 28, 29) */,
  32'h3d1cff11 /* (22, 28, 29) */,
  32'h3d3b1e93 /* (18, 28, 29) */,
  32'h3d3b1e93 /* (14, 28, 29) */,
  32'h3d1cff11 /* (10, 28, 29) */,
  32'h3d1b3fff /* (6, 28, 29) */,
  32'h3d5defd3 /* (2, 28, 29) */,
  32'h3d13e9f7 /* (30, 24, 29) */,
  32'h3d19bf4b /* (26, 24, 29) */,
  32'h3d48bc7e /* (22, 24, 29) */,
  32'h3d880501 /* (18, 24, 29) */,
  32'h3d880501 /* (14, 24, 29) */,
  32'h3d48bc7e /* (10, 24, 29) */,
  32'h3d19bf4b /* (6, 24, 29) */,
  32'h3d13e9f7 /* (2, 24, 29) */,
  32'h3d23d587 /* (30, 20, 29) */,
  32'h3d48406d /* (26, 20, 29) */,
  32'h3d9aff71 /* (22, 20, 29) */,
  32'h3decc5e8 /* (18, 20, 29) */,
  32'h3decc5e8 /* (14, 20, 29) */,
  32'h3d9aff71 /* (10, 20, 29) */,
  32'h3d48406d /* (6, 20, 29) */,
  32'h3d23d587 /* (2, 20, 29) */,
  32'h3d13661d /* (30, 16, 29) */,
  32'h3d41d3ae /* (26, 16, 29) */,
  32'h3da59d10 /* (22, 16, 29) */,
  32'h3e0a27e7 /* (18, 16, 29) */,
  32'h3e0a27e7 /* (14, 16, 29) */,
  32'h3da59d10 /* (10, 16, 29) */,
  32'h3d41d3ae /* (6, 16, 29) */,
  32'h3d13661d /* (2, 16, 29) */,
  32'h3d23d587 /* (30, 12, 29) */,
  32'h3d48406d /* (26, 12, 29) */,
  32'h3d9aff71 /* (22, 12, 29) */,
  32'h3decc5e8 /* (18, 12, 29) */,
  32'h3decc5e8 /* (14, 12, 29) */,
  32'h3d9aff71 /* (10, 12, 29) */,
  32'h3d48406d /* (6, 12, 29) */,
  32'h3d23d587 /* (2, 12, 29) */,
  32'h3d13e9f7 /* (30, 8, 29) */,
  32'h3d19bf4b /* (26, 8, 29) */,
  32'h3d48bc7e /* (22, 8, 29) */,
  32'h3d880501 /* (18, 8, 29) */,
  32'h3d880501 /* (14, 8, 29) */,
  32'h3d48bc7e /* (10, 8, 29) */,
  32'h3d19bf4b /* (6, 8, 29) */,
  32'h3d13e9f7 /* (2, 8, 29) */,
  32'h3d5defd3 /* (30, 4, 29) */,
  32'h3d1b3fff /* (26, 4, 29) */,
  32'h3d1cff11 /* (22, 4, 29) */,
  32'h3d3b1e93 /* (18, 4, 29) */,
  32'h3d3b1e93 /* (14, 4, 29) */,
  32'h3d1cff11 /* (10, 4, 29) */,
  32'h3d1b3fff /* (6, 4, 29) */,
  32'h3d5defd3 /* (2, 4, 29) */,
  32'h3dcbea25 /* (30, 0, 29) */,
  32'h3d2d5b95 /* (26, 0, 29) */,
  32'h3d144f19 /* (22, 0, 29) */,
  32'h3d262b6e /* (18, 0, 29) */,
  32'h3d262b6e /* (14, 0, 29) */,
  32'h3d144f19 /* (10, 0, 29) */,
  32'h3d2d5b95 /* (6, 0, 29) */,
  32'h3dcbea25 /* (2, 0, 29) */,
  32'h3d16c6a3 /* (30, 28, 25) */,
  32'h3d17902e /* (26, 28, 25) */,
  32'h3d404057 /* (22, 28, 25) */,
  32'h3d800deb /* (18, 28, 25) */,
  32'h3d800deb /* (14, 28, 25) */,
  32'h3d404057 /* (10, 28, 25) */,
  32'h3d17902e /* (6, 28, 25) */,
  32'h3d16c6a3 /* (2, 28, 25) */,
  32'h3d1d59b0 /* (30, 24, 25) */,
  32'h3d35cd98 /* (26, 24, 25) */,
  32'h3d83c517 /* (22, 24, 25) */,
  32'h3dbf672f /* (18, 24, 25) */,
  32'h3dbf672f /* (14, 24, 25) */,
  32'h3d83c517 /* (10, 24, 25) */,
  32'h3d35cd98 /* (6, 24, 25) */,
  32'h3d1d59b0 /* (2, 24, 25) */,
  32'h3d530d8e /* (30, 20, 25) */,
  32'h3d859348 /* (26, 20, 25) */,
  32'h3dd85675 /* (22, 20, 25) */,
  32'h3e2baf50 /* (18, 20, 25) */,
  32'h3e2baf50 /* (14, 20, 25) */,
  32'h3dd85675 /* (10, 20, 25) */,
  32'h3d859348 /* (6, 20, 25) */,
  32'h3d530d8e /* (2, 20, 25) */,
  32'h3d4f6a6e /* (30, 16, 25) */,
  32'h3d8a46e7 /* (26, 16, 25) */,
  32'h3df142da /* (22, 16, 25) */,
  32'h3e4d7ce8 /* (18, 16, 25) */,
  32'h3e4d7ce8 /* (14, 16, 25) */,
  32'h3df142da /* (10, 16, 25) */,
  32'h3d8a46e7 /* (6, 16, 25) */,
  32'h3d4f6a6e /* (2, 16, 25) */,
  32'h3d530d8e /* (30, 12, 25) */,
  32'h3d859348 /* (26, 12, 25) */,
  32'h3dd85675 /* (22, 12, 25) */,
  32'h3e2baf50 /* (18, 12, 25) */,
  32'h3e2baf50 /* (14, 12, 25) */,
  32'h3dd85675 /* (10, 12, 25) */,
  32'h3d859348 /* (6, 12, 25) */,
  32'h3d530d8e /* (2, 12, 25) */,
  32'h3d1d59b0 /* (30, 8, 25) */,
  32'h3d35cd98 /* (26, 8, 25) */,
  32'h3d83c517 /* (22, 8, 25) */,
  32'h3dbf672f /* (18, 8, 25) */,
  32'h3dbf672f /* (14, 8, 25) */,
  32'h3d83c517 /* (10, 8, 25) */,
  32'h3d35cd98 /* (6, 8, 25) */,
  32'h3d1d59b0 /* (2, 8, 25) */,
  32'h3d16c6a3 /* (30, 4, 25) */,
  32'h3d17902e /* (26, 4, 25) */,
  32'h3d404057 /* (22, 4, 25) */,
  32'h3d800deb /* (18, 4, 25) */,
  32'h3d800deb /* (14, 4, 25) */,
  32'h3d404057 /* (10, 4, 25) */,
  32'h3d17902e /* (6, 4, 25) */,
  32'h3d16c6a3 /* (2, 4, 25) */,
  32'h3d21b235 /* (30, 0, 25) */,
  32'h3d1459dd /* (26, 0, 25) */,
  32'h3d2f5f5a /* (22, 0, 25) */,
  32'h3d60bf24 /* (18, 0, 25) */,
  32'h3d60bf24 /* (14, 0, 25) */,
  32'h3d2f5f5a /* (10, 0, 25) */,
  32'h3d1459dd /* (6, 0, 25) */,
  32'h3d21b235 /* (2, 0, 25) */,
  32'h3d21c128 /* (30, 28, 21) */,
  32'h3d41fb9f /* (26, 28, 21) */,
  32'h3d92b699 /* (22, 28, 21) */,
  32'h3ddc0819 /* (18, 28, 21) */,
  32'h3ddc0819 /* (14, 28, 21) */,
  32'h3d92b699 /* (10, 28, 21) */,
  32'h3d41fb9f /* (6, 28, 21) */,
  32'h3d21c128 /* (2, 28, 21) */,
  32'h3d558b1c /* (30, 24, 21) */,
  32'h3d865b59 /* (26, 24, 21) */,
  32'h3dd7e578 /* (22, 24, 21) */,
  32'h3e2a27e4 /* (18, 24, 21) */,
  32'h3e2a27e4 /* (14, 24, 21) */,
  32'h3dd7e578 /* (10, 24, 21) */,
  32'h3d865b59 /* (6, 24, 21) */,
  32'h3d558b1c /* (2, 24, 21) */,
  32'h3da96c08 /* (30, 20, 21) */,
  32'h3ddec971 /* (26, 20, 21) */,
  32'h3e3e5baf /* (22, 20, 21) */,
  32'h3e9ecc49 /* (18, 20, 21) */,
  32'h3e9ecc49 /* (14, 20, 21) */,
  32'h3e3e5baf /* (10, 20, 21) */,
  32'h3ddec971 /* (6, 20, 21) */,
  32'h3da96c08 /* (2, 20, 21) */,
  32'h3db86416 /* (30, 16, 21) */,
  32'h3dfa4afe /* (26, 16, 21) */,
  32'h3e60898b /* (22, 16, 21) */,
  32'h3ec4f0a1 /* (18, 16, 21) */,
  32'h3ec4f0a1 /* (14, 16, 21) */,
  32'h3e60898b /* (10, 16, 21) */,
  32'h3dfa4afe /* (6, 16, 21) */,
  32'h3db86416 /* (2, 16, 21) */,
  32'h3da96c08 /* (30, 12, 21) */,
  32'h3ddec971 /* (26, 12, 21) */,
  32'h3e3e5baf /* (22, 12, 21) */,
  32'h3e9ecc49 /* (18, 12, 21) */,
  32'h3e9ecc49 /* (14, 12, 21) */,
  32'h3e3e5baf /* (10, 12, 21) */,
  32'h3ddec971 /* (6, 12, 21) */,
  32'h3da96c08 /* (2, 12, 21) */,
  32'h3d558b1c /* (30, 8, 21) */,
  32'h3d865b59 /* (26, 8, 21) */,
  32'h3dd7e578 /* (22, 8, 21) */,
  32'h3e2a27e4 /* (18, 8, 21) */,
  32'h3e2a27e4 /* (14, 8, 21) */,
  32'h3dd7e578 /* (10, 8, 21) */,
  32'h3d865b59 /* (6, 8, 21) */,
  32'h3d558b1c /* (2, 8, 21) */,
  32'h3d21c128 /* (30, 4, 21) */,
  32'h3d41fb9f /* (26, 4, 21) */,
  32'h3d92b699 /* (22, 4, 21) */,
  32'h3ddc0819 /* (18, 4, 21) */,
  32'h3ddc0819 /* (14, 4, 21) */,
  32'h3d92b699 /* (10, 4, 21) */,
  32'h3d41fb9f /* (6, 4, 21) */,
  32'h3d21c128 /* (2, 4, 21) */,
  32'h3d164ce1 /* (30, 0, 21) */,
  32'h3d3013e2 /* (26, 0, 21) */,
  32'h3d819abc /* (22, 0, 21) */,
  32'h3dbe661f /* (18, 0, 21) */,
  32'h3dbe661f /* (14, 0, 21) */,
  32'h3d819abc /* (10, 0, 21) */,
  32'h3d3013e2 /* (6, 0, 21) */,
  32'h3d164ce1 /* (2, 0, 21) */,
  32'h3d2d6bba /* (30, 28, 17) */,
  32'h3d61b1de /* (26, 28, 17) */,
  32'h3dbdf4f8 /* (22, 28, 17) */,
  32'h3e1c2ca1 /* (18, 28, 17) */,
  32'h3e1c2ca1 /* (14, 28, 17) */,
  32'h3dbdf4f8 /* (10, 28, 17) */,
  32'h3d61b1de /* (6, 28, 17) */,
  32'h3d2d6bba /* (2, 28, 17) */,
  32'h3d804df8 /* (30, 24, 17) */,
  32'h3daa3349 /* (26, 24, 17) */,
  32'h3e135573 /* (22, 24, 17) */,
  32'h3e79034c /* (18, 24, 17) */,
  32'h3e79034c /* (14, 24, 17) */,
  32'h3e135573 /* (10, 24, 17) */,
  32'h3daa3349 /* (6, 24, 17) */,
  32'h3d804df8 /* (2, 24, 17) */,
  32'h3de39dff /* (30, 20, 17) */,
  32'h3e1a3a56 /* (26, 20, 17) */,
  32'h3e89fde5 /* (22, 20, 17) */,
  32'h3ef15f91 /* (18, 20, 17) */,
  32'h3ef15f91 /* (14, 20, 17) */,
  32'h3e89fde5 /* (10, 20, 17) */,
  32'h3e1a3a56 /* (6, 20, 17) */,
  32'h3de39dff /* (2, 20, 17) */,
  32'h3e06ec2e /* (30, 16, 17) */,
  32'h3e3a3d1a /* (26, 16, 17) */,
  32'h3eabb572 /* (22, 16, 17) */,
  32'h3f1b42bd /* (18, 16, 17) */,
  32'h3f1b42bd /* (14, 16, 17) */,
  32'h3eabb572 /* (10, 16, 17) */,
  32'h3e3a3d1a /* (6, 16, 17) */,
  32'h3e06ec2e /* (2, 16, 17) */,
  32'h3de39dff /* (30, 12, 17) */,
  32'h3e1a3a56 /* (26, 12, 17) */,
  32'h3e89fde5 /* (22, 12, 17) */,
  32'h3ef15f91 /* (18, 12, 17) */,
  32'h3ef15f91 /* (14, 12, 17) */,
  32'h3e89fde5 /* (10, 12, 17) */,
  32'h3e1a3a56 /* (6, 12, 17) */,
  32'h3de39dff /* (2, 12, 17) */,
  32'h3d804df8 /* (30, 8, 17) */,
  32'h3daa3349 /* (26, 8, 17) */,
  32'h3e135573 /* (22, 8, 17) */,
  32'h3e79034c /* (18, 8, 17) */,
  32'h3e79034c /* (14, 8, 17) */,
  32'h3e135573 /* (10, 8, 17) */,
  32'h3daa3349 /* (6, 8, 17) */,
  32'h3d804df8 /* (2, 8, 17) */,
  32'h3d2d6bba /* (30, 4, 17) */,
  32'h3d61b1de /* (26, 4, 17) */,
  32'h3dbdf4f8 /* (22, 4, 17) */,
  32'h3e1c2ca1 /* (18, 4, 17) */,
  32'h3e1c2ca1 /* (14, 4, 17) */,
  32'h3dbdf4f8 /* (10, 4, 17) */,
  32'h3d61b1de /* (6, 4, 17) */,
  32'h3d2d6bba /* (2, 4, 17) */,
  32'h3d18d610 /* (30, 0, 17) */,
  32'h3d455011 /* (26, 0, 17) */,
  32'h3da42e1b /* (22, 0, 17) */,
  32'h3e05899d /* (18, 0, 17) */,
  32'h3e05899d /* (14, 0, 17) */,
  32'h3da42e1b /* (10, 0, 17) */,
  32'h3d455011 /* (6, 0, 17) */,
  32'h3d18d610 /* (2, 0, 17) */,
  32'h3d3217f4 /* (30, 28, 13) */,
  32'h3d601ae9 /* (26, 28, 13) */,
  32'h3db40e50 /* (22, 28, 13) */,
  32'h3e0de89e /* (18, 28, 13) */,
  32'h3e0de89e /* (14, 28, 13) */,
  32'h3db40e50 /* (10, 28, 13) */,
  32'h3d601ae9 /* (6, 28, 13) */,
  32'h3d3217f4 /* (2, 28, 13) */,
  32'h3d7b52f8 /* (30, 24, 13) */,
  32'h3da2e7a9 /* (26, 24, 13) */,
  32'h3e085939 /* (22, 24, 13) */,
  32'h3e5f05ce /* (18, 24, 13) */,
  32'h3e5f05ce /* (14, 24, 13) */,
  32'h3e085939 /* (10, 24, 13) */,
  32'h3da2e7a9 /* (6, 24, 13) */,
  32'h3d7b52f8 /* (2, 24, 13) */,
  32'h3dd42d31 /* (30, 20, 13) */,
  32'h3e0dc95f /* (26, 20, 13) */,
  32'h3e7848b5 /* (22, 20, 13) */,
  32'h3ed441df /* (18, 20, 13) */,
  32'h3ed441df /* (14, 20, 13) */,
  32'h3e7848b5 /* (10, 20, 13) */,
  32'h3e0dc95f /* (6, 20, 13) */,
  32'h3dd42d31 /* (2, 20, 13) */,
  32'h3df1ae3d /* (30, 16, 13) */,
  32'h3e2576a9 /* (26, 16, 13) */,
  32'h3e968a40 /* (22, 16, 13) */,
  32'h3f06176f /* (18, 16, 13) */,
  32'h3f06176f /* (14, 16, 13) */,
  32'h3e968a40 /* (10, 16, 13) */,
  32'h3e2576a9 /* (6, 16, 13) */,
  32'h3df1ae3d /* (2, 16, 13) */,
  32'h3dd42d31 /* (30, 12, 13) */,
  32'h3e0dc95f /* (26, 12, 13) */,
  32'h3e7848b5 /* (22, 12, 13) */,
  32'h3ed441df /* (18, 12, 13) */,
  32'h3ed441df /* (14, 12, 13) */,
  32'h3e7848b5 /* (10, 12, 13) */,
  32'h3e0dc95f /* (6, 12, 13) */,
  32'h3dd42d31 /* (2, 12, 13) */,
  32'h3d7b52f8 /* (30, 8, 13) */,
  32'h3da2e7a9 /* (26, 8, 13) */,
  32'h3e085939 /* (22, 8, 13) */,
  32'h3e5f05ce /* (18, 8, 13) */,
  32'h3e5f05ce /* (14, 8, 13) */,
  32'h3e085939 /* (10, 8, 13) */,
  32'h3da2e7a9 /* (6, 8, 13) */,
  32'h3d7b52f8 /* (2, 8, 13) */,
  32'h3d3217f4 /* (30, 4, 13) */,
  32'h3d601ae9 /* (26, 4, 13) */,
  32'h3db40e50 /* (22, 4, 13) */,
  32'h3e0de89e /* (18, 4, 13) */,
  32'h3e0de89e /* (14, 4, 13) */,
  32'h3db40e50 /* (10, 4, 13) */,
  32'h3d601ae9 /* (6, 4, 13) */,
  32'h3d3217f4 /* (2, 4, 13) */,
  32'h3d2045b1 /* (30, 0, 13) */,
  32'h3d4703b2 /* (26, 0, 13) */,
  32'h3d9d248b /* (22, 0, 13) */,
  32'h3df40add /* (18, 0, 13) */,
  32'h3df40add /* (14, 0, 13) */,
  32'h3d9d248b /* (10, 0, 13) */,
  32'h3d4703b2 /* (6, 0, 13) */,
  32'h3d2045b1 /* (2, 0, 13) */,
  32'h3d14de35 /* (30, 28, 9) */,
  32'h3d2657dd /* (26, 28, 9) */,
  32'h3d68b7a2 /* (22, 28, 9) */,
  32'h3da4db8a /* (18, 28, 9) */,
  32'h3da4db8a /* (14, 28, 9) */,
  32'h3d68b7a2 /* (10, 28, 9) */,
  32'h3d2657dd /* (6, 28, 9) */,
  32'h3d14de35 /* (2, 28, 9) */,
  32'h3d3291f6 /* (30, 24, 9) */,
  32'h3d584c0c /* (26, 24, 9) */,
  32'h3da590e9 /* (22, 24, 9) */,
  32'h3dfaaa60 /* (18, 24, 9) */,
  32'h3dfaaa60 /* (14, 24, 9) */,
  32'h3da590e9 /* (10, 24, 9) */,
  32'h3d584c0c /* (6, 24, 9) */,
  32'h3d3291f6 /* (2, 24, 9) */,
  32'h3d833332 /* (30, 20, 9) */,
  32'h3da96159 /* (26, 20, 9) */,
  32'h3e0cf021 /* (22, 20, 9) */,
  32'h3e654448 /* (18, 20, 9) */,
  32'h3e654448 /* (14, 20, 9) */,
  32'h3e0cf021 /* (10, 20, 9) */,
  32'h3da96159 /* (6, 20, 9) */,
  32'h3d833332 /* (2, 20, 9) */,
  32'h3d87d16b /* (30, 16, 9) */,
  32'h3db6b309 /* (26, 16, 9) */,
  32'h3e21930d /* (22, 16, 9) */,
  32'h3e8b9344 /* (18, 16, 9) */,
  32'h3e8b9344 /* (14, 16, 9) */,
  32'h3e21930d /* (10, 16, 9) */,
  32'h3db6b309 /* (6, 16, 9) */,
  32'h3d87d16b /* (2, 16, 9) */,
  32'h3d833332 /* (30, 12, 9) */,
  32'h3da96159 /* (26, 12, 9) */,
  32'h3e0cf021 /* (22, 12, 9) */,
  32'h3e654448 /* (18, 12, 9) */,
  32'h3e654448 /* (14, 12, 9) */,
  32'h3e0cf021 /* (10, 12, 9) */,
  32'h3da96159 /* (6, 12, 9) */,
  32'h3d833332 /* (2, 12, 9) */,
  32'h3d3291f6 /* (30, 8, 9) */,
  32'h3d584c0c /* (26, 8, 9) */,
  32'h3da590e9 /* (22, 8, 9) */,
  32'h3dfaaa60 /* (18, 8, 9) */,
  32'h3dfaaa60 /* (14, 8, 9) */,
  32'h3da590e9 /* (10, 8, 9) */,
  32'h3d584c0c /* (6, 8, 9) */,
  32'h3d3291f6 /* (2, 8, 9) */,
  32'h3d14de35 /* (30, 4, 9) */,
  32'h3d2657dd /* (26, 4, 9) */,
  32'h3d68b7a2 /* (22, 4, 9) */,
  32'h3da4db8a /* (18, 4, 9) */,
  32'h3da4db8a /* (14, 4, 9) */,
  32'h3d68b7a2 /* (10, 4, 9) */,
  32'h3d2657dd /* (6, 4, 9) */,
  32'h3d14de35 /* (2, 4, 9) */,
  32'h3d11b684 /* (30, 0, 9) */,
  32'h3d1bc36a /* (26, 0, 9) */,
  32'h3d50a575 /* (22, 0, 9) */,
  32'h3d8fa52c /* (18, 0, 9) */,
  32'h3d8fa52c /* (14, 0, 9) */,
  32'h3d50a575 /* (10, 0, 9) */,
  32'h3d1bc36a /* (6, 0, 9) */,
  32'h3d11b684 /* (2, 0, 9) */,
  32'h3d2d8e0e /* (30, 28, 5) */,
  32'h3d153e19 /* (26, 28, 5) */,
  32'h3d28e3b2 /* (22, 28, 5) */,
  32'h3d53bb31 /* (18, 28, 5) */,
  32'h3d53bb31 /* (14, 28, 5) */,
  32'h3d28e3b2 /* (10, 28, 5) */,
  32'h3d153e19 /* (6, 28, 5) */,
  32'h3d2d8e0e /* (2, 28, 5) */,
  32'h3d149b5c /* (30, 24, 5) */,
  32'h3d22af34 /* (26, 24, 5) */,
  32'h3d5ef675 /* (22, 24, 5) */,
  32'h3d9bc970 /* (18, 24, 5) */,
  32'h3d9bc970 /* (14, 24, 5) */,
  32'h3d5ef675 /* (10, 24, 5) */,
  32'h3d22af34 /* (6, 24, 5) */,
  32'h3d149b5c /* (2, 24, 5) */,
  32'h3d346b02 /* (30, 20, 5) */,
  32'h3d6007ad /* (26, 20, 5) */,
  32'h3db0e528 /* (22, 20, 5) */,
  32'h3e095be4 /* (18, 20, 5) */,
  32'h3e095be4 /* (14, 20, 5) */,
  32'h3db0e528 /* (10, 20, 5) */,
  32'h3d6007ad /* (6, 20, 5) */,
  32'h3d346b02 /* (2, 20, 5) */,
  32'h3d28d1e5 /* (30, 16, 5) */,
  32'h3d5f53fb /* (26, 16, 5) */,
  32'h3dc0863e /* (22, 16, 5) */,
  32'h3e2205a1 /* (18, 16, 5) */,
  32'h3e2205a1 /* (14, 16, 5) */,
  32'h3dc0863e /* (10, 16, 5) */,
  32'h3d5f53fb /* (6, 16, 5) */,
  32'h3d28d1e5 /* (2, 16, 5) */,
  32'h3d346b02 /* (30, 12, 5) */,
  32'h3d6007ad /* (26, 12, 5) */,
  32'h3db0e528 /* (22, 12, 5) */,
  32'h3e095be4 /* (18, 12, 5) */,
  32'h3e095be4 /* (14, 12, 5) */,
  32'h3db0e528 /* (10, 12, 5) */,
  32'h3d6007ad /* (6, 12, 5) */,
  32'h3d346b02 /* (2, 12, 5) */,
  32'h3d149b5c /* (30, 8, 5) */,
  32'h3d22af34 /* (26, 8, 5) */,
  32'h3d5ef675 /* (22, 8, 5) */,
  32'h3d9bc970 /* (18, 8, 5) */,
  32'h3d9bc970 /* (14, 8, 5) */,
  32'h3d5ef675 /* (10, 8, 5) */,
  32'h3d22af34 /* (6, 8, 5) */,
  32'h3d149b5c /* (2, 8, 5) */,
  32'h3d2d8e0e /* (30, 4, 5) */,
  32'h3d153e19 /* (26, 4, 5) */,
  32'h3d28e3b2 /* (22, 4, 5) */,
  32'h3d53bb31 /* (18, 4, 5) */,
  32'h3d53bb31 /* (14, 4, 5) */,
  32'h3d28e3b2 /* (10, 4, 5) */,
  32'h3d153e19 /* (6, 4, 5) */,
  32'h3d2d8e0e /* (2, 4, 5) */,
  32'h3d5dd7d1 /* (30, 0, 5) */,
  32'h3d1b2f33 /* (26, 0, 5) */,
  32'h3d1cee15 /* (22, 0, 5) */,
  32'h3d3b0a55 /* (18, 0, 5) */,
  32'h3d3b0a55 /* (14, 0, 5) */,
  32'h3d1cee15 /* (10, 0, 5) */,
  32'h3d1b2f33 /* (6, 0, 5) */,
  32'h3d5dd7d1 /* (2, 0, 5) */,
  32'h3d8b1391 /* (30, 28, 1) */,
  32'h3d222a9c /* (26, 28, 1) */,
  32'h3d1839e3 /* (22, 28, 1) */,
  32'h3d303352 /* (18, 28, 1) */,
  32'h3d303352 /* (14, 28, 1) */,
  32'h3d1839e3 /* (10, 28, 1) */,
  32'h3d222a9c /* (6, 28, 1) */,
  32'h3d8b1391 /* (2, 28, 1) */,
  32'h3d15ce12 /* (30, 24, 1) */,
  32'h3d169650 /* (26, 24, 1) */,
  32'h3d3f0366 /* (22, 24, 1) */,
  32'h3d7e759f /* (18, 24, 1) */,
  32'h3d7e759f /* (14, 24, 1) */,
  32'h3d3f0366 /* (10, 24, 1) */,
  32'h3d169650 /* (6, 24, 1) */,
  32'h3d15ce12 /* (2, 24, 1) */,
  32'h3d1cac31 /* (30, 20, 1) */,
  32'h3d3dc5f0 /* (26, 20, 1) */,
  32'h3d91435f /* (22, 20, 1) */,
  32'h3ddbed5a /* (18, 20, 1) */,
  32'h3ddbed5a /* (14, 20, 1) */,
  32'h3d91435f /* (10, 20, 1) */,
  32'h3d3dc5f0 /* (6, 20, 1) */,
  32'h3d1cac31 /* (2, 20, 1) */,
  32'h3d09dfab /* (30, 16, 1) */,
  32'h3d34b66a /* (26, 16, 1) */,
  32'h3d99ac24 /* (22, 16, 1) */,
  32'h3dff32bb /* (18, 16, 1) */,
  32'h3dff32bb /* (14, 16, 1) */,
  32'h3d99ac24 /* (10, 16, 1) */,
  32'h3d34b66a /* (6, 16, 1) */,
  32'h3d09dfab /* (2, 16, 1) */,
  32'h3d1cac31 /* (30, 12, 1) */,
  32'h3d3dc5f0 /* (26, 12, 1) */,
  32'h3d91435f /* (22, 12, 1) */,
  32'h3ddbed5a /* (18, 12, 1) */,
  32'h3ddbed5a /* (14, 12, 1) */,
  32'h3d91435f /* (10, 12, 1) */,
  32'h3d3dc5f0 /* (6, 12, 1) */,
  32'h3d1cac31 /* (2, 12, 1) */,
  32'h3d15ce12 /* (30, 8, 1) */,
  32'h3d169650 /* (26, 8, 1) */,
  32'h3d3f0366 /* (22, 8, 1) */,
  32'h3d7e759f /* (18, 8, 1) */,
  32'h3d7e759f /* (14, 8, 1) */,
  32'h3d3f0366 /* (10, 8, 1) */,
  32'h3d169650 /* (6, 8, 1) */,
  32'h3d15ce12 /* (2, 8, 1) */,
  32'h3d8b1391 /* (30, 4, 1) */,
  32'h3d222a9c /* (26, 4, 1) */,
  32'h3d1839e3 /* (22, 4, 1) */,
  32'h3d303352 /* (18, 4, 1) */,
  32'h3d303352 /* (14, 4, 1) */,
  32'h3d1839e3 /* (10, 4, 1) */,
  32'h3d222a9c /* (6, 4, 1) */,
  32'h3d8b1391 /* (2, 4, 1) */,
  32'h3e709592 /* (30, 0, 1) */,
  32'h3d3f59b8 /* (26, 0, 1) */,
  32'h3d1142bb /* (22, 0, 1) */,
  32'h3d1ceee6 /* (18, 0, 1) */,
  32'h3d1ceee6 /* (14, 0, 1) */,
  32'h3d1142bb /* (10, 0, 1) */,
  32'h3d3f59b8 /* (6, 0, 1) */,
  32'h3e709592 /* (2, 0, 1) */,
  32'h3d4920d0 /* (29, 28, 29) */,
  32'h3d155fa4 /* (25, 28, 29) */,
  32'h3d25fa09 /* (21, 28, 29) */,
  32'h3d349293 /* (17, 28, 29) */,
  32'h3d385879 /* (13, 28, 29) */,
  32'h3d16b5b2 /* (9, 28, 29) */,
  32'h3d25f5ce /* (5, 28, 29) */,
  32'h3d6eb36b /* (1, 28, 29) */,
  32'h3d1392fe /* (29, 24, 29) */,
  32'h3d2054cd /* (25, 24, 29) */,
  32'h3d5d0a38 /* (21, 24, 29) */,
  32'h3d8608f0 /* (17, 24, 29) */,
  32'h3d82c188 /* (13, 24, 29) */,
  32'h3d37919e /* (9, 24, 29) */,
  32'h3d15d660 /* (5, 24, 29) */,
  32'h3d146963 /* (1, 24, 29) */,
  32'h3d28b308 /* (29, 20, 29) */,
  32'h3d5ab0e1 /* (25, 20, 29) */,
  32'h3db0b965 /* (21, 20, 29) */,
  32'h3deea44d /* (17, 20, 29) */,
  32'h3dddef48 /* (13, 20, 29) */,
  32'h3d886b82 /* (9, 20, 29) */,
  32'h3d3a4ebb /* (5, 20, 29) */,
  32'h3d210eee /* (1, 20, 29) */,
  32'h3d19c07a /* (29, 16, 29) */,
  32'h3d58de26 /* (25, 16, 29) */,
  32'h3dc1602b /* (21, 16, 29) */,
  32'h3e0de417 /* (17, 16, 29) */,
  32'h3dfdd31f /* (13, 16, 29) */,
  32'h3d8e3848 /* (9, 16, 29) */,
  32'h3d3046d8 /* (5, 16, 29) */,
  32'h3d0fbc59 /* (1, 16, 29) */,
  32'h3d28b308 /* (29, 12, 29) */,
  32'h3d5ab0e1 /* (25, 12, 29) */,
  32'h3db0b965 /* (21, 12, 29) */,
  32'h3deea44d /* (17, 12, 29) */,
  32'h3dddef48 /* (13, 12, 29) */,
  32'h3d886b82 /* (9, 12, 29) */,
  32'h3d3a4ebb /* (5, 12, 29) */,
  32'h3d210eee /* (1, 12, 29) */,
  32'h3d1392fe /* (29, 8, 29) */,
  32'h3d2054cd /* (25, 8, 29) */,
  32'h3d5d0a38 /* (21, 8, 29) */,
  32'h3d8608f0 /* (17, 8, 29) */,
  32'h3d82c188 /* (13, 8, 29) */,
  32'h3d37919e /* (9, 8, 29) */,
  32'h3d15d660 /* (5, 8, 29) */,
  32'h3d146963 /* (1, 8, 29) */,
  32'h3d4920d0 /* (29, 4, 29) */,
  32'h3d155fa4 /* (25, 4, 29) */,
  32'h3d25fa09 /* (21, 4, 29) */,
  32'h3d349293 /* (17, 4, 29) */,
  32'h3d385879 /* (13, 4, 29) */,
  32'h3d16b5b2 /* (9, 4, 29) */,
  32'h3d25f5ce /* (5, 4, 29) */,
  32'h3d6eb36b /* (1, 4, 29) */,
  32'h3d9c797c /* (29, 0, 29) */,
  32'h3d1cfd70 /* (25, 0, 29) */,
  32'h3d198ce9 /* (21, 0, 29) */,
  32'h3d1eeabe /* (17, 0, 29) */,
  32'h3d258110 /* (13, 0, 29) */,
  32'h3d1237a7 /* (9, 0, 29) */,
  32'h3d490b0e /* (5, 0, 29) */,
  32'h3dff9e3f /* (1, 0, 29) */,
  32'h3d155fa4 /* (29, 28, 25) */,
  32'h3d1cbb18 /* (25, 28, 25) */,
  32'h3d52976b /* (21, 28, 25) */,
  32'h3d7b9f11 /* (17, 28, 25) */,
  32'h3d770afc /* (13, 28, 25) */,
  32'h3d30de15 /* (9, 28, 25) */,
  32'h3d1508af /* (5, 28, 25) */,
  32'h3d17ff6b /* (1, 28, 25) */,
  32'h3d2054cd /* (29, 24, 25) */,
  32'h3d432bf1 /* (25, 24, 25) */,
  32'h3d941bce /* (21, 24, 25) */,
  32'h3dbf0444 /* (17, 24, 25) */,
  32'h3db56072 /* (13, 24, 25) */,
  32'h3d6b8b35 /* (9, 24, 25) */,
  32'h3d2bff3e /* (5, 24, 25) */,
  32'h3d1bb8b6 /* (1, 24, 25) */,
  32'h3d5ab0e1 /* (29, 20, 25) */,
  32'h3d938890 /* (25, 20, 25) */,
  32'h3df94537 /* (21, 20, 25) */,
  32'h3e2e6a71 /* (17, 20, 25) */,
  32'h3e1f8cbf /* (13, 20, 25) */,
  32'h3dbc51f9 /* (9, 20, 25) */,
  32'h3d75e4d4 /* (5, 20, 25) */,
  32'h3d4ea8e5 /* (1, 20, 25) */,
  32'h3d58de26 /* (29, 16, 25) */,
  32'h3d9b7830 /* (25, 16, 25) */,
  32'h3e0d9cf0 /* (21, 16, 25) */,
  32'h3e540b9b /* (17, 16, 25) */,
  32'h3e3bd4ee /* (13, 16, 25) */,
  32'h3dce1075 /* (9, 16, 25) */,
  32'h3d7a662c /* (5, 16, 25) */,
  32'h3d49f75a /* (1, 16, 25) */,
  32'h3d5ab0e1 /* (29, 12, 25) */,
  32'h3d938890 /* (25, 12, 25) */,
  32'h3df94537 /* (21, 12, 25) */,
  32'h3e2e6a71 /* (17, 12, 25) */,
  32'h3e1f8cbf /* (13, 12, 25) */,
  32'h3dbc51f9 /* (9, 12, 25) */,
  32'h3d75e4d4 /* (5, 12, 25) */,
  32'h3d4ea8e5 /* (1, 12, 25) */,
  32'h3d2054cd /* (29, 8, 25) */,
  32'h3d432bf1 /* (25, 8, 25) */,
  32'h3d941bce /* (21, 8, 25) */,
  32'h3dbf0444 /* (17, 8, 25) */,
  32'h3db56072 /* (13, 8, 25) */,
  32'h3d6b8b35 /* (9, 8, 25) */,
  32'h3d2bff3e /* (5, 8, 25) */,
  32'h3d1bb8b6 /* (1, 8, 25) */,
  32'h3d155fa4 /* (29, 4, 25) */,
  32'h3d1cbb18 /* (25, 4, 25) */,
  32'h3d52976b /* (21, 4, 25) */,
  32'h3d7b9f11 /* (17, 4, 25) */,
  32'h3d770afc /* (13, 4, 25) */,
  32'h3d30de15 /* (9, 4, 25) */,
  32'h3d1508af /* (5, 4, 25) */,
  32'h3d17ff6b /* (1, 4, 25) */,
  32'h3d1cfd70 /* (29, 0, 25) */,
  32'h3d162f74 /* (25, 0, 25) */,
  32'h3d3dcd22 /* (21, 0, 25) */,
  32'h3d5b6048 /* (17, 0, 25) */,
  32'h3d5a6fdd /* (13, 0, 25) */,
  32'h3d23a039 /* (9, 0, 25) */,
  32'h3d154f7b /* (5, 0, 25) */,
  32'h3d25463b /* (1, 0, 25) */,
  32'h3d25fa09 /* (29, 28, 21) */,
  32'h3d52976b /* (25, 28, 21) */,
  32'h3da66ad4 /* (21, 28, 21) */,
  32'h3ddcf428 /* (17, 28, 21) */,
  32'h3dcf13a3 /* (13, 28, 21) */,
  32'h3d81d711 /* (9, 28, 21) */,
  32'h3d358341 /* (5, 28, 21) */,
  32'h3d1f5dc3 /* (1, 28, 21) */,
  32'h3d5d0a38 /* (29, 24, 21) */,
  32'h3d941bce /* (25, 24, 21) */,
  32'h3df84bb3 /* (21, 24, 21) */,
  32'h3e2c9c6c /* (17, 24, 21) */,
  32'h3e1e607d /* (13, 24, 21) */,
  32'h3dbc4d73 /* (9, 24, 21) */,
  32'h3d77c8fd /* (5, 24, 21) */,
  32'h3d513c3d /* (1, 24, 21) */,
  32'h3db0b965 /* (29, 20, 21) */,
  32'h3df94537 /* (25, 20, 21) */,
  32'h3e5e44ac /* (21, 20, 21) */,
  32'h3ea31756 /* (17, 20, 21) */,
  32'h3e91dfe2 /* (13, 20, 21) */,
  32'h3e23781b /* (9, 20, 21) */,
  32'h3dca9d53 /* (5, 20, 21) */,
  32'h3da53628 /* (1, 20, 21) */,
  32'h3dc1602b /* (29, 16, 21) */,
  32'h3e0d9cf0 /* (25, 16, 21) */,
  32'h3e84c8e0 /* (21, 16, 21) */,
  32'h3ecca1ac /* (17, 16, 21) */,
  32'h3eb2bd2a /* (13, 16, 21) */,
  32'h3e3e5da7 /* (9, 16, 21) */,
  32'h3de14ffa /* (5, 16, 21) */,
  32'h3db336e0 /* (1, 16, 21) */,
  32'h3db0b965 /* (29, 12, 21) */,
  32'h3df94537 /* (25, 12, 21) */,
  32'h3e5e44ac /* (21, 12, 21) */,
  32'h3ea31756 /* (17, 12, 21) */,
  32'h3e91dfe2 /* (13, 12, 21) */,
  32'h3e23781b /* (9, 12, 21) */,
  32'h3dca9d53 /* (5, 12, 21) */,
  32'h3da53628 /* (1, 12, 21) */,
  32'h3d5d0a38 /* (29, 8, 21) */,
  32'h3d941bce /* (25, 8, 21) */,
  32'h3df84bb3 /* (21, 8, 21) */,
  32'h3e2c9c6c /* (17, 8, 21) */,
  32'h3e1e607d /* (13, 8, 21) */,
  32'h3dbc4d73 /* (9, 8, 21) */,
  32'h3d77c8fd /* (5, 8, 21) */,
  32'h3d513c3d /* (1, 8, 21) */,
  32'h3d25fa09 /* (29, 4, 21) */,
  32'h3d52976b /* (25, 4, 21) */,
  32'h3da66ad4 /* (21, 4, 21) */,
  32'h3ddcf428 /* (17, 4, 21) */,
  32'h3dcf13a3 /* (13, 4, 21) */,
  32'h3d81d711 /* (9, 4, 21) */,
  32'h3d358341 /* (5, 4, 21) */,
  32'h3d1f5dc3 /* (1, 4, 21) */,
  32'h3d198ce9 /* (29, 0, 21) */,
  32'h3d3dcd22 /* (25, 0, 21) */,
  32'h3d922642 /* (21, 0, 21) */,
  32'h3dbe6d47 /* (17, 0, 21) */,
  32'h3db3fd83 /* (13, 0, 21) */,
  32'h3d66dac1 /* (9, 0, 21) */,
  32'h3d25e815 /* (5, 0, 21) */,
  32'h3d147e90 /* (1, 0, 21) */,
  32'h3d349293 /* (29, 28, 17) */,
  32'h3d7b9f11 /* (25, 28, 17) */,
  32'h3ddcf428 /* (21, 28, 17) */,
  32'h3e1fe07e /* (17, 28, 17) */,
  32'h3e0ff4ce /* (13, 28, 17) */,
  32'h3da3c1ed /* (9, 28, 17) */,
  32'h3d4def9b /* (5, 28, 17) */,
  32'h3d294c4b /* (1, 28, 17) */,
  32'h3d8608f0 /* (29, 24, 17) */,
  32'h3dbf0444 /* (25, 24, 17) */,
  32'h3e2c9c6c /* (21, 24, 17) */,
  32'h3e803f85 /* (17, 24, 17) */,
  32'h3e640ba2 /* (13, 24, 17) */,
  32'h3dfc30a3 /* (9, 24, 17) */,
  32'h3d9a5b6b /* (5, 24, 17) */,
  32'h3d7a003f /* (1, 24, 17) */,
  32'h3deea44d /* (29, 20, 17) */,
  32'h3e2e6a71 /* (25, 20, 17) */,
  32'h3ea31756 /* (21, 20, 17) */,
  32'h3efaa119 /* (17, 20, 17) */,
  32'h3edb3822 /* (13, 20, 17) */,
  32'h3e6a25fd /* (9, 20, 17) */,
  32'h3e0ae903 /* (5, 20, 17) */,
  32'h3ddd43c2 /* (1, 20, 17) */,
  32'h3e0de417 /* (29, 16, 17) */,
  32'h3e540b9b /* (25, 16, 17) */,
  32'h3ecca1ac /* (21, 16, 17) */,
  32'h3f2286f8 /* (17, 16, 17) */,
  32'h3f0bd969 /* (13, 16, 17) */,
  32'h3e908107 /* (9, 16, 17) */,
  32'h3e26bbbb /* (5, 16, 17) */,
  32'h3e02e976 /* (1, 16, 17) */,
  32'h3deea44d /* (29, 12, 17) */,
  32'h3e2e6a71 /* (25, 12, 17) */,
  32'h3ea31756 /* (21, 12, 17) */,
  32'h3efaa119 /* (17, 12, 17) */,
  32'h3edb3822 /* (13, 12, 17) */,
  32'h3e6a25fd /* (9, 12, 17) */,
  32'h3e0ae903 /* (5, 12, 17) */,
  32'h3ddd43c2 /* (1, 12, 17) */,
  32'h3d8608f0 /* (29, 8, 17) */,
  32'h3dbf0444 /* (25, 8, 17) */,
  32'h3e2c9c6c /* (21, 8, 17) */,
  32'h3e803f85 /* (17, 8, 17) */,
  32'h3e640ba2 /* (13, 8, 17) */,
  32'h3dfc30a3 /* (9, 8, 17) */,
  32'h3d9a5b6b /* (5, 8, 17) */,
  32'h3d7a003f /* (1, 8, 17) */,
  32'h3d349293 /* (29, 4, 17) */,
  32'h3d7b9f11 /* (25, 4, 17) */,
  32'h3ddcf428 /* (21, 4, 17) */,
  32'h3e1fe07e /* (17, 4, 17) */,
  32'h3e0ff4ce /* (13, 4, 17) */,
  32'h3da3c1ed /* (9, 4, 17) */,
  32'h3d4def9b /* (5, 4, 17) */,
  32'h3d294c4b /* (1, 4, 17) */,
  32'h3d1eeabe /* (29, 0, 17) */,
  32'h3d5b6048 /* (25, 0, 17) */,
  32'h3dbe6d47 /* (21, 0, 17) */,
  32'h3e086183 /* (17, 0, 17) */,
  32'h3df6cc6d /* (13, 0, 17) */,
  32'h3d8df2c1 /* (9, 0, 17) */,
  32'h3d347f0a /* (5, 0, 17) */,
  32'h3d155505 /* (1, 0, 17) */,
  32'h3d385879 /* (29, 28, 13) */,
  32'h3d770afc /* (25, 28, 13) */,
  32'h3dcf13a3 /* (21, 28, 13) */,
  32'h3e0ff4ce /* (17, 28, 13) */,
  32'h3e0415cb /* (13, 28, 13) */,
  32'h3d9d0afa /* (9, 28, 13) */,
  32'h3d4ea6a0 /* (5, 28, 13) */,
  32'h3d2e802a /* (1, 28, 13) */,
  32'h3d82c188 /* (29, 24, 13) */,
  32'h3db56072 /* (25, 24, 13) */,
  32'h3e1e607d /* (21, 24, 13) */,
  32'h3e640ba2 /* (17, 24, 13) */,
  32'h3e4dd3dc /* (13, 24, 13) */,
  32'h3deb6b6d /* (9, 24, 13) */,
  32'h3d94d380 /* (5, 24, 13) */,
  32'h3d7573b6 /* (1, 24, 13) */,
  32'h3dddef48 /* (29, 20, 13) */,
  32'h3e1f8cbf /* (25, 20, 13) */,
  32'h3e91dfe2 /* (21, 20, 13) */,
  32'h3edb3822 /* (17, 20, 13) */,
  32'h3ec1d890 /* (13, 20, 13) */,
  32'h3e53dc51 /* (9, 20, 13) */,
  32'h3e00477d /* (5, 20, 13) */,
  32'h3dce8d02 /* (1, 20, 13) */,
  32'h3dfdd31f /* (29, 16, 13) */,
  32'h3e3bd4ee /* (25, 16, 13) */,
  32'h3eb2bd2a /* (21, 16, 13) */,
  32'h3f0bd969 /* (17, 16, 13) */,
  32'h3ef27895 /* (13, 16, 13) */,
  32'h3e7e4b9d /* (9, 16, 13) */,
  32'h3e1486b7 /* (5, 16, 13) */,
  32'h3deaafef /* (1, 16, 13) */,
  32'h3dddef48 /* (29, 12, 13) */,
  32'h3e1f8cbf /* (25, 12, 13) */,
  32'h3e91dfe2 /* (21, 12, 13) */,
  32'h3edb3822 /* (17, 12, 13) */,
  32'h3ec1d890 /* (13, 12, 13) */,
  32'h3e53dc51 /* (9, 12, 13) */,
  32'h3e00477d /* (5, 12, 13) */,
  32'h3dce8d02 /* (1, 12, 13) */,
  32'h3d82c188 /* (29, 8, 13) */,
  32'h3db56072 /* (25, 8, 13) */,
  32'h3e1e607d /* (21, 8, 13) */,
  32'h3e640ba2 /* (17, 8, 13) */,
  32'h3e4dd3dc /* (13, 8, 13) */,
  32'h3deb6b6d /* (9, 8, 13) */,
  32'h3d94d380 /* (5, 8, 13) */,
  32'h3d7573b6 /* (1, 8, 13) */,
  32'h3d385879 /* (29, 4, 13) */,
  32'h3d770afc /* (25, 4, 13) */,
  32'h3dcf13a3 /* (21, 4, 13) */,
  32'h3e0ff4ce /* (17, 4, 13) */,
  32'h3e0415cb /* (13, 4, 13) */,
  32'h3d9d0afa /* (9, 4, 13) */,
  32'h3d4ea6a0 /* (5, 4, 13) */,
  32'h3d2e802a /* (1, 4, 13) */,
  32'h3d258110 /* (29, 0, 13) */,
  32'h3d5a6fdd /* (25, 0, 13) */,
  32'h3db3fd83 /* (21, 0, 13) */,
  32'h3df6cc6d /* (17, 0, 13) */,
  32'h3de3e928 /* (13, 0, 13) */,
  32'h3d89a49e /* (9, 0, 13) */,
  32'h3d384488 /* (5, 0, 13) */,
  32'h3d1d4601 /* (1, 0, 13) */,
  32'h3d16b5b2 /* (29, 28, 9) */,
  32'h3d30de15 /* (25, 28, 9) */,
  32'h3d81d711 /* (21, 28, 9) */,
  32'h3da3c1ed /* (17, 28, 9) */,
  32'h3d9d0afa /* (13, 28, 9) */,
  32'h3d51a9d2 /* (9, 28, 9) */,
  32'h3d1ee50b /* (5, 28, 9) */,
  32'h3d13f199 /* (1, 28, 9) */,
  32'h3d37919e /* (29, 24, 9) */,
  32'h3d6b8b35 /* (25, 24, 9) */,
  32'h3dbc4d73 /* (21, 24, 9) */,
  32'h3dfc30a3 /* (17, 24, 9) */,
  32'h3deb6b6d /* (13, 24, 9) */,
  32'h3d921bde /* (9, 24, 9) */,
  32'h3d49c96c /* (5, 24, 9) */,
  32'h3d2fba80 /* (1, 24, 9) */,
  32'h3d886b82 /* (29, 20, 9) */,
  32'h3dbc51f9 /* (25, 20, 9) */,
  32'h3e23781b /* (21, 20, 9) */,
  32'h3e6a25fd /* (17, 20, 9) */,
  32'h3e53dc51 /* (13, 20, 9) */,
  32'h3df3b4f2 /* (9, 20, 9) */,
  32'h3d9af1c2 /* (5, 20, 9) */,
  32'h3d803124 /* (1, 20, 9) */,
  32'h3d8e3848 /* (29, 16, 9) */,
  32'h3dce1075 /* (25, 16, 9) */,
  32'h3e3e5da7 /* (21, 16, 9) */,
  32'h3e908107 /* (17, 16, 9) */,
  32'h3e7e4b9d /* (13, 16, 9) */,
  32'h3e0981d7 /* (9, 16, 9) */,
  32'h3da4f2f4 /* (5, 16, 9) */,
  32'h3d8420c9 /* (1, 16, 9) */,
  32'h3d886b82 /* (29, 12, 9) */,
  32'h3dbc51f9 /* (25, 12, 9) */,
  32'h3e23781b /* (21, 12, 9) */,
  32'h3e6a25fd /* (17, 12, 9) */,
  32'h3e53dc51 /* (13, 12, 9) */,
  32'h3df3b4f2 /* (9, 12, 9) */,
  32'h3d9af1c2 /* (5, 12, 9) */,
  32'h3d803124 /* (1, 12, 9) */,
  32'h3d37919e /* (29, 8, 9) */,
  32'h3d6b8b35 /* (25, 8, 9) */,
  32'h3dbc4d73 /* (21, 8, 9) */,
  32'h3dfc30a3 /* (17, 8, 9) */,
  32'h3deb6b6d /* (13, 8, 9) */,
  32'h3d921bde /* (9, 8, 9) */,
  32'h3d49c96c /* (5, 8, 9) */,
  32'h3d2fba80 /* (1, 8, 9) */,
  32'h3d16b5b2 /* (29, 4, 9) */,
  32'h3d30de15 /* (25, 4, 9) */,
  32'h3d81d711 /* (21, 4, 9) */,
  32'h3da3c1ed /* (17, 4, 9) */,
  32'h3d9d0afa /* (13, 4, 9) */,
  32'h3d51a9d2 /* (9, 4, 9) */,
  32'h3d1ee50b /* (5, 4, 9) */,
  32'h3d13f199 /* (1, 4, 9) */,
  32'h3d1237a7 /* (29, 0, 9) */,
  32'h3d23a039 /* (25, 0, 9) */,
  32'h3d66dac1 /* (21, 0, 9) */,
  32'h3d8df2c1 /* (17, 0, 9) */,
  32'h3d89a49e /* (13, 0, 9) */,
  32'h3d3dc47d /* (9, 0, 9) */,
  32'h3d16a564 /* (5, 0, 9) */,
  32'h3d11a5c6 /* (1, 0, 9) */,
  32'h3d25f5ce /* (29, 28, 5) */,
  32'h3d1508af /* (25, 28, 5) */,
  32'h3d358341 /* (21, 28, 5) */,
  32'h3d4def9b /* (17, 28, 5) */,
  32'h3d4ea6a0 /* (13, 28, 5) */,
  32'h3d1ee50b /* (9, 28, 5) */,
  32'h3d189061 /* (5, 28, 5) */,
  32'h3d334ee4 /* (1, 28, 5) */,
  32'h3d15d660 /* (29, 24, 5) */,
  32'h3d2bff3e /* (25, 24, 5) */,
  32'h3d77c8fd /* (21, 24, 5) */,
  32'h3d9a5b6b /* (17, 24, 5) */,
  32'h3d94d380 /* (13, 24, 5) */,
  32'h3d49c96c /* (9, 24, 5) */,
  32'h3d1c4d38 /* (5, 24, 5) */,
  32'h3d1412fd /* (1, 24, 5) */,
  32'h3d3a4ebb /* (29, 20, 5) */,
  32'h3d75e4d4 /* (25, 20, 5) */,
  32'h3dca9d53 /* (21, 20, 5) */,
  32'h3e0ae903 /* (17, 20, 5) */,
  32'h3e00477d /* (13, 20, 5) */,
  32'h3d9af1c2 /* (9, 20, 5) */,
  32'h3d4f6dfc /* (5, 20, 5) */,
  32'h3d310ad3 /* (1, 20, 5) */,
  32'h3d3046d8 /* (29, 16, 5) */,
  32'h3d7a662c /* (25, 16, 5) */,
  32'h3de14ffa /* (21, 16, 5) */,
  32'h3e26bbbb /* (17, 16, 5) */,
  32'h3e1486b7 /* (13, 16, 5) */,
  32'h3da4f2f4 /* (9, 16, 5) */,
  32'h3d4ab7f7 /* (5, 16, 5) */,
  32'h3d24852f /* (1, 16, 5) */,
  32'h3d3a4ebb /* (29, 12, 5) */,
  32'h3d75e4d4 /* (25, 12, 5) */,
  32'h3dca9d53 /* (21, 12, 5) */,
  32'h3e0ae903 /* (17, 12, 5) */,
  32'h3e00477d /* (13, 12, 5) */,
  32'h3d9af1c2 /* (9, 12, 5) */,
  32'h3d4f6dfc /* (5, 12, 5) */,
  32'h3d310ad3 /* (1, 12, 5) */,
  32'h3d15d660 /* (29, 8, 5) */,
  32'h3d2bff3e /* (25, 8, 5) */,
  32'h3d77c8fd /* (21, 8, 5) */,
  32'h3d9a5b6b /* (17, 8, 5) */,
  32'h3d94d380 /* (13, 8, 5) */,
  32'h3d49c96c /* (9, 8, 5) */,
  32'h3d1c4d38 /* (5, 8, 5) */,
  32'h3d1412fd /* (1, 8, 5) */,
  32'h3d25f5ce /* (29, 4, 5) */,
  32'h3d1508af /* (25, 4, 5) */,
  32'h3d358341 /* (21, 4, 5) */,
  32'h3d4def9b /* (17, 4, 5) */,
  32'h3d4ea6a0 /* (13, 4, 5) */,
  32'h3d1ee50b /* (9, 4, 5) */,
  32'h3d189061 /* (5, 4, 5) */,
  32'h3d334ee4 /* (1, 4, 5) */,
  32'h3d490b0e /* (29, 0, 5) */,
  32'h3d154f7b /* (25, 0, 5) */,
  32'h3d25e815 /* (21, 0, 5) */,
  32'h3d347f0a /* (17, 0, 5) */,
  32'h3d384488 /* (13, 0, 5) */,
  32'h3d16a564 /* (9, 0, 5) */,
  32'h3d25e3da /* (5, 0, 5) */,
  32'h3d6e9998 /* (1, 0, 5) */,
  32'h3d6eb36b /* (29, 28, 1) */,
  32'h3d17ff6b /* (25, 28, 1) */,
  32'h3d1f5dc3 /* (21, 28, 1) */,
  32'h3d294c4b /* (17, 28, 1) */,
  32'h3d2e802a /* (13, 28, 1) */,
  32'h3d13f199 /* (9, 28, 1) */,
  32'h3d334ee4 /* (5, 28, 1) */,
  32'h3d9c757b /* (1, 28, 1) */,
  32'h3d146963 /* (29, 24, 1) */,
  32'h3d1bb8b6 /* (25, 24, 1) */,
  32'h3d513c3d /* (21, 24, 1) */,
  32'h3d7a003f /* (17, 24, 1) */,
  32'h3d7573b6 /* (13, 24, 1) */,
  32'h3d2fba80 /* (9, 24, 1) */,
  32'h3d1412fd /* (5, 24, 1) */,
  32'h3d1704d7 /* (1, 24, 1) */,
  32'h3d210eee /* (29, 20, 1) */,
  32'h3d4ea8e5 /* (25, 20, 1) */,
  32'h3da53628 /* (21, 20, 1) */,
  32'h3ddd43c2 /* (17, 20, 1) */,
  32'h3dce8d02 /* (13, 20, 1) */,
  32'h3d803124 /* (9, 20, 1) */,
  32'h3d310ad3 /* (5, 20, 1) */,
  32'h3d1a2df1 /* (1, 20, 1) */,
  32'h3d0fbc59 /* (29, 16, 1) */,
  32'h3d49f75a /* (25, 16, 1) */,
  32'h3db336e0 /* (21, 16, 1) */,
  32'h3e02e976 /* (17, 16, 1) */,
  32'h3deaafef /* (13, 16, 1) */,
  32'h3d8420c9 /* (9, 16, 1) */,
  32'h3d24852f /* (5, 16, 1) */,
  32'h3d067e68 /* (1, 16, 1) */,
  32'h3d210eee /* (29, 12, 1) */,
  32'h3d4ea8e5 /* (25, 12, 1) */,
  32'h3da53628 /* (21, 12, 1) */,
  32'h3ddd43c2 /* (17, 12, 1) */,
  32'h3dce8d02 /* (13, 12, 1) */,
  32'h3d803124 /* (9, 12, 1) */,
  32'h3d310ad3 /* (5, 12, 1) */,
  32'h3d1a2df1 /* (1, 12, 1) */,
  32'h3d146963 /* (29, 8, 1) */,
  32'h3d1bb8b6 /* (25, 8, 1) */,
  32'h3d513c3d /* (21, 8, 1) */,
  32'h3d7a003f /* (17, 8, 1) */,
  32'h3d7573b6 /* (13, 8, 1) */,
  32'h3d2fba80 /* (9, 8, 1) */,
  32'h3d1412fd /* (5, 8, 1) */,
  32'h3d1704d7 /* (1, 8, 1) */,
  32'h3d6eb36b /* (29, 4, 1) */,
  32'h3d17ff6b /* (25, 4, 1) */,
  32'h3d1f5dc3 /* (21, 4, 1) */,
  32'h3d294c4b /* (17, 4, 1) */,
  32'h3d2e802a /* (13, 4, 1) */,
  32'h3d13f199 /* (9, 4, 1) */,
  32'h3d334ee4 /* (5, 4, 1) */,
  32'h3d9c757b /* (1, 4, 1) */,
  32'h3dff9e3f /* (29, 0, 1) */,
  32'h3d25463b /* (25, 0, 1) */,
  32'h3d147e90 /* (21, 0, 1) */,
  32'h3d155505 /* (17, 0, 1) */,
  32'h3d1d4601 /* (13, 0, 1) */,
  32'h3d11a5c6 /* (9, 0, 1) */,
  32'h3d6e9998 /* (5, 0, 1) */,
  32'h3f10fe39 /* (1, 0, 1) */,
  32'h3d358b49 /* (28, 28, 29) */,
  32'h3d13fed6 /* (24, 28, 29) */,
  32'h3d30047a /* (20, 28, 29) */,
  32'h3d232f37 /* (16, 28, 29) */,
  32'h3d30047a /* (12, 28, 29) */,
  32'h3d13fed6 /* (8, 28, 29) */,
  32'h3d358b49 /* (4, 28, 29) */,
  32'h3d7541a2 /* (0, 28, 29) */,
  32'h3d13fed6 /* (28, 24, 29) */,
  32'h3d2a2238 /* (24, 24, 29) */,
  32'h3d729483 /* (20, 24, 29) */,
  32'h3d76a38f /* (16, 24, 29) */,
  32'h3d729483 /* (12, 24, 29) */,
  32'h3d2a2238 /* (8, 24, 29) */,
  32'h3d13fed6 /* (4, 24, 29) */,
  32'h3d14a194 /* (0, 24, 29) */,
  32'h3d30047a /* (28, 20, 29) */,
  32'h3d729483 /* (24, 20, 29) */,
  32'h3dc823b1 /* (20, 20, 29) */,
  32'h3de007f6 /* (16, 20, 29) */,
  32'h3dc823b1 /* (12, 20, 29) */,
  32'h3d729483 /* (8, 20, 29) */,
  32'h3d30047a /* (4, 20, 29) */,
  32'h3d202826 /* (0, 20, 29) */,
  32'h3d232f37 /* (28, 16, 29) */,
  32'h3d76a38f /* (24, 16, 29) */,
  32'h3de007f6 /* (20, 16, 29) */,
  32'h3e078d5a /* (16, 16, 29) */,
  32'h3de007f6 /* (12, 16, 29) */,
  32'h3d76a38f /* (8, 16, 29) */,
  32'h3d232f37 /* (4, 16, 29) */,
  32'h3d0e89f8 /* (0, 16, 29) */,
  32'h3d30047a /* (28, 12, 29) */,
  32'h3d729483 /* (24, 12, 29) */,
  32'h3dc823b1 /* (20, 12, 29) */,
  32'h3de007f6 /* (16, 12, 29) */,
  32'h3dc823b1 /* (12, 12, 29) */,
  32'h3d729483 /* (8, 12, 29) */,
  32'h3d30047a /* (4, 12, 29) */,
  32'h3d202826 /* (0, 12, 29) */,
  32'h3d13fed6 /* (28, 8, 29) */,
  32'h3d2a2238 /* (24, 8, 29) */,
  32'h3d729483 /* (20, 8, 29) */,
  32'h3d76a38f /* (16, 8, 29) */,
  32'h3d729483 /* (12, 8, 29) */,
  32'h3d2a2238 /* (8, 8, 29) */,
  32'h3d13fed6 /* (4, 8, 29) */,
  32'h3d14a194 /* (0, 8, 29) */,
  32'h3d358b49 /* (28, 4, 29) */,
  32'h3d13fed6 /* (24, 4, 29) */,
  32'h3d30047a /* (20, 4, 29) */,
  32'h3d232f37 /* (16, 4, 29) */,
  32'h3d30047a /* (12, 4, 29) */,
  32'h3d13fed6 /* (8, 4, 29) */,
  32'h3d358b49 /* (4, 4, 29) */,
  32'h3d7541a2 /* (0, 4, 29) */,
  32'h3d7541a2 /* (28, 0, 29) */,
  32'h3d14a194 /* (24, 0, 29) */,
  32'h3d202826 /* (20, 0, 29) */,
  32'h3d0e89f8 /* (16, 0, 29) */,
  32'h3d202826 /* (12, 0, 29) */,
  32'h3d14a194 /* (8, 0, 29) */,
  32'h3d7541a2 /* (4, 0, 29) */,
  32'h3e0c4c59 /* (0, 0, 29) */,
  32'h3d148979 /* (28, 28, 25) */,
  32'h3d250b86 /* (24, 28, 25) */,
  32'h3d66108f /* (20, 28, 25) */,
  32'h3d66e7bc /* (16, 28, 25) */,
  32'h3d66108f /* (12, 28, 25) */,
  32'h3d250b86 /* (8, 28, 25) */,
  32'h3d148979 /* (4, 28, 25) */,
  32'h3d1879c9 /* (0, 28, 25) */,
  32'h3d250b86 /* (28, 24, 25) */,
  32'h3d54dbd1 /* (24, 24, 25) */,
  32'h3da58a7f /* (20, 24, 25) */,
  32'h3db1ba44 /* (16, 24, 25) */,
  32'h3da58a7f /* (12, 24, 25) */,
  32'h3d54dbd1 /* (8, 24, 25) */,
  32'h3d250b86 /* (4, 24, 25) */,
  32'h3d1b34b2 /* (0, 24, 25) */,
  32'h3d66108f /* (28, 20, 25) */,
  32'h3da58a7f /* (24, 20, 25) */,
  32'h3e0e8e1e /* (20, 20, 25) */,
  32'h3e24eefd /* (16, 20, 25) */,
  32'h3e0e8e1e /* (12, 20, 25) */,
  32'h3da58a7f /* (8, 20, 25) */,
  32'h3d66108f /* (4, 20, 25) */,
  32'h3d4d39f8 /* (0, 20, 25) */,
  32'h3d66e7bc /* (28, 16, 25) */,
  32'h3db1ba44 /* (24, 16, 25) */,
  32'h3e24eefd /* (20, 16, 25) */,
  32'h3e4b7c7a /* (16, 16, 25) */,
  32'h3e24eefd /* (12, 16, 25) */,
  32'h3db1ba44 /* (8, 16, 25) */,
  32'h3d66e7bc /* (4, 16, 25) */,
  32'h3d482f92 /* (0, 16, 25) */,
  32'h3d66108f /* (28, 12, 25) */,
  32'h3da58a7f /* (24, 12, 25) */,
  32'h3e0e8e1e /* (20, 12, 25) */,
  32'h3e24eefd /* (16, 12, 25) */,
  32'h3e0e8e1e /* (12, 12, 25) */,
  32'h3da58a7f /* (8, 12, 25) */,
  32'h3d66108f /* (4, 12, 25) */,
  32'h3d4d39f8 /* (0, 12, 25) */,
  32'h3d250b86 /* (28, 8, 25) */,
  32'h3d54dbd1 /* (24, 8, 25) */,
  32'h3da58a7f /* (20, 8, 25) */,
  32'h3db1ba44 /* (16, 8, 25) */,
  32'h3da58a7f /* (12, 8, 25) */,
  32'h3d54dbd1 /* (8, 8, 25) */,
  32'h3d250b86 /* (4, 8, 25) */,
  32'h3d1b34b2 /* (0, 8, 25) */,
  32'h3d148979 /* (28, 4, 25) */,
  32'h3d250b86 /* (24, 4, 25) */,
  32'h3d66108f /* (20, 4, 25) */,
  32'h3d66e7bc /* (16, 4, 25) */,
  32'h3d66108f /* (12, 4, 25) */,
  32'h3d250b86 /* (8, 4, 25) */,
  32'h3d148979 /* (4, 4, 25) */,
  32'h3d1879c9 /* (0, 4, 25) */,
  32'h3d1879c9 /* (28, 0, 25) */,
  32'h3d1b34b2 /* (24, 0, 25) */,
  32'h3d4d39f8 /* (20, 0, 25) */,
  32'h3d482f92 /* (16, 0, 25) */,
  32'h3d4d39f8 /* (12, 0, 25) */,
  32'h3d1b34b2 /* (8, 0, 25) */,
  32'h3d1879c9 /* (4, 0, 25) */,
  32'h3d269d45 /* (0, 0, 25) */,
  32'h3d2c64eb /* (28, 28, 21) */,
  32'h3d683712 /* (24, 28, 21) */,
  32'h3dbb90ec /* (20, 28, 21) */,
  32'h3dcebbc1 /* (16, 28, 21) */,
  32'h3dbb90ec /* (12, 28, 21) */,
  32'h3d683712 /* (8, 28, 21) */,
  32'h3d2c64eb /* (4, 28, 21) */,
  32'h3d1e982c /* (0, 28, 21) */,
  32'h3d683712 /* (28, 24, 21) */,
  32'h3da5dafd /* (24, 24, 21) */,
  32'h3e0dbead /* (20, 24, 21) */,
  32'h3e2301df /* (16, 24, 21) */,
  32'h3e0dbead /* (12, 24, 21) */,
  32'h3da5dafd /* (8, 24, 21) */,
  32'h3d683712 /* (4, 24, 21) */,
  32'h3d4fd499 /* (0, 24, 21) */,
  32'h3dbb90ec /* (28, 20, 21) */,
  32'h3e0dbead /* (24, 20, 21) */,
  32'h3e80c082 /* (20, 20, 21) */,
  32'h3e9bce24 /* (16, 20, 21) */,
  32'h3e80c082 /* (12, 20, 21) */,
  32'h3e0dbead /* (8, 20, 21) */,
  32'h3dbb90ec /* (4, 20, 21) */,
  32'h3da3d600 /* (0, 20, 21) */,
  32'h3dcebbc1 /* (28, 16, 21) */,
  32'h3e2301df /* (24, 16, 21) */,
  32'h3e9bce24 /* (20, 16, 21) */,
  32'h3ec5ad99 /* (16, 16, 21) */,
  32'h3e9bce24 /* (12, 16, 21) */,
  32'h3e2301df /* (8, 16, 21) */,
  32'h3dcebbc1 /* (4, 16, 21) */,
  32'h3db1860e /* (0, 16, 21) */,
  32'h3dbb90ec /* (28, 12, 21) */,
  32'h3e0dbead /* (24, 12, 21) */,
  32'h3e80c082 /* (20, 12, 21) */,
  32'h3e9bce24 /* (16, 12, 21) */,
  32'h3e80c082 /* (12, 12, 21) */,
  32'h3e0dbead /* (8, 12, 21) */,
  32'h3dbb90ec /* (4, 12, 21) */,
  32'h3da3d600 /* (0, 12, 21) */,
  32'h3d683712 /* (28, 8, 21) */,
  32'h3da5dafd /* (24, 8, 21) */,
  32'h3e0dbead /* (20, 8, 21) */,
  32'h3e2301df /* (16, 8, 21) */,
  32'h3e0dbead /* (12, 8, 21) */,
  32'h3da5dafd /* (8, 8, 21) */,
  32'h3d683712 /* (4, 8, 21) */,
  32'h3d4fd499 /* (0, 8, 21) */,
  32'h3d2c64eb /* (28, 4, 21) */,
  32'h3d683712 /* (24, 4, 21) */,
  32'h3dbb90ec /* (20, 4, 21) */,
  32'h3dcebbc1 /* (16, 4, 21) */,
  32'h3dbb90ec /* (12, 4, 21) */,
  32'h3d683712 /* (8, 4, 21) */,
  32'h3d2c64eb /* (4, 4, 21) */,
  32'h3d1e982c /* (0, 4, 21) */,
  32'h3d1e982c /* (28, 0, 21) */,
  32'h3d4fd499 /* (24, 0, 21) */,
  32'h3da3d600 /* (20, 0, 21) */,
  32'h3db1860e /* (16, 0, 21) */,
  32'h3da3d600 /* (12, 0, 21) */,
  32'h3d4fd499 /* (8, 0, 21) */,
  32'h3d1e982c /* (4, 0, 21) */,
  32'h3d13eab3 /* (0, 0, 21) */,
  32'h3d3f317e /* (28, 28, 17) */,
  32'h3d8e8b3a /* (24, 28, 17) */,
  32'h3dff07bf /* (20, 28, 17) */,
  32'h3e18449a /* (16, 28, 17) */,
  32'h3dff07bf /* (12, 28, 17) */,
  32'h3d8e8b3a /* (8, 28, 17) */,
  32'h3d3f317e /* (4, 28, 17) */,
  32'h3d27f384 /* (0, 28, 17) */,
  32'h3d8e8b3a /* (28, 24, 17) */,
  32'h3dd9f1d0 /* (24, 24, 17) */,
  32'h3e48a298 /* (20, 24, 17) */,
  32'h3e75b861 /* (16, 24, 17) */,
  32'h3e48a298 /* (12, 24, 17) */,
  32'h3dd9f1d0 /* (8, 24, 17) */,
  32'h3d8e8b3a /* (4, 24, 17) */,
  32'h3d77d78b /* (0, 24, 17) */,
  32'h3dff07bf /* (28, 20, 17) */,
  32'h3e48a298 /* (24, 20, 17) */,
  32'h3ebf3a63 /* (20, 20, 17) */,
  32'h3ef1f40b /* (16, 20, 17) */,
  32'h3ebf3a63 /* (12, 20, 17) */,
  32'h3e48a298 /* (8, 20, 17) */,
  32'h3dff07bf /* (4, 20, 17) */,
  32'h3ddb309a /* (0, 20, 17) */,
  32'h3e18449a /* (28, 16, 17) */,
  32'h3e75b861 /* (24, 16, 17) */,
  32'h3ef1f40b /* (20, 16, 17) */,
  32'h3f1e253a /* (16, 16, 17) */,
  32'h3ef1f40b /* (12, 16, 17) */,
  32'h3e75b861 /* (8, 16, 17) */,
  32'h3e18449a /* (4, 16, 17) */,
  32'h3e019a4f /* (0, 16, 17) */,
  32'h3dff07bf /* (28, 12, 17) */,
  32'h3e48a298 /* (24, 12, 17) */,
  32'h3ebf3a63 /* (20, 12, 17) */,
  32'h3ef1f40b /* (16, 12, 17) */,
  32'h3ebf3a63 /* (12, 12, 17) */,
  32'h3e48a298 /* (8, 12, 17) */,
  32'h3dff07bf /* (4, 12, 17) */,
  32'h3ddb309a /* (0, 12, 17) */,
  32'h3d8e8b3a /* (28, 8, 17) */,
  32'h3dd9f1d0 /* (24, 8, 17) */,
  32'h3e48a298 /* (20, 8, 17) */,
  32'h3e75b861 /* (16, 8, 17) */,
  32'h3e48a298 /* (12, 8, 17) */,
  32'h3dd9f1d0 /* (8, 8, 17) */,
  32'h3d8e8b3a /* (4, 8, 17) */,
  32'h3d77d78b /* (0, 8, 17) */,
  32'h3d3f317e /* (28, 4, 17) */,
  32'h3d8e8b3a /* (24, 4, 17) */,
  32'h3dff07bf /* (20, 4, 17) */,
  32'h3e18449a /* (16, 4, 17) */,
  32'h3dff07bf /* (12, 4, 17) */,
  32'h3d8e8b3a /* (8, 4, 17) */,
  32'h3d3f317e /* (4, 4, 17) */,
  32'h3d27f384 /* (0, 4, 17) */,
  32'h3d27f384 /* (28, 0, 17) */,
  32'h3d77d78b /* (24, 0, 17) */,
  32'h3ddb309a /* (20, 0, 17) */,
  32'h3e019a4f /* (16, 0, 17) */,
  32'h3ddb309a /* (12, 0, 17) */,
  32'h3d77d78b /* (8, 0, 17) */,
  32'h3d27f384 /* (4, 0, 17) */,
  32'h3d14300c /* (0, 0, 17) */,
  32'h3d41aa67 /* (28, 28, 13) */,
  32'h3d8a5278 /* (24, 28, 13) */,
  32'h3dec6d9f /* (20, 28, 13) */,
  32'h3e07f264 /* (16, 28, 13) */,
  32'h3dec6d9f /* (12, 28, 13) */,
  32'h3d8a5278 /* (8, 28, 13) */,
  32'h3d41aa67 /* (4, 28, 13) */,
  32'h3d2d543a /* (0, 28, 13) */,
  32'h3d8a5278 /* (28, 24, 13) */,
  32'h3dcd36cb /* (24, 24, 13) */,
  32'h3e368e5b /* (20, 24, 13) */,
  32'h3e58f4b1 /* (16, 24, 13) */,
  32'h3e368e5b /* (12, 24, 13) */,
  32'h3dcd36cb /* (8, 24, 13) */,
  32'h3d8a5278 /* (4, 24, 13) */,
  32'h3d7388b1 /* (0, 24, 13) */,
  32'h3dec6d9f /* (28, 20, 13) */,
  32'h3e368e5b /* (24, 20, 13) */,
  32'h3eaa0eb2 /* (20, 20, 13) */,
  32'h3ed28b29 /* (16, 20, 13) */,
  32'h3eaa0eb2 /* (12, 20, 13) */,
  32'h3e368e5b /* (8, 20, 13) */,
  32'h3dec6d9f /* (4, 20, 13) */,
  32'h3dccb681 /* (0, 20, 13) */,
  32'h3e07f264 /* (28, 16, 13) */,
  32'h3e58f4b1 /* (24, 16, 13) */,
  32'h3ed28b29 /* (20, 16, 13) */,
  32'h3f079668 /* (16, 16, 13) */,
  32'h3ed28b29 /* (12, 16, 13) */,
  32'h3e58f4b1 /* (8, 16, 13) */,
  32'h3e07f264 /* (4, 16, 13) */,
  32'h3de8675d /* (0, 16, 13) */,
  32'h3dec6d9f /* (28, 12, 13) */,
  32'h3e368e5b /* (24, 12, 13) */,
  32'h3eaa0eb2 /* (20, 12, 13) */,
  32'h3ed28b29 /* (16, 12, 13) */,
  32'h3eaa0eb2 /* (12, 12, 13) */,
  32'h3e368e5b /* (8, 12, 13) */,
  32'h3dec6d9f /* (4, 12, 13) */,
  32'h3dccb681 /* (0, 12, 13) */,
  32'h3d8a5278 /* (28, 8, 13) */,
  32'h3dcd36cb /* (24, 8, 13) */,
  32'h3e368e5b /* (20, 8, 13) */,
  32'h3e58f4b1 /* (16, 8, 13) */,
  32'h3e368e5b /* (12, 8, 13) */,
  32'h3dcd36cb /* (8, 8, 13) */,
  32'h3d8a5278 /* (4, 8, 13) */,
  32'h3d7388b1 /* (0, 8, 13) */,
  32'h3d41aa67 /* (28, 4, 13) */,
  32'h3d8a5278 /* (24, 4, 13) */,
  32'h3dec6d9f /* (20, 4, 13) */,
  32'h3e07f264 /* (16, 4, 13) */,
  32'h3dec6d9f /* (12, 4, 13) */,
  32'h3d8a5278 /* (8, 4, 13) */,
  32'h3d41aa67 /* (4, 4, 13) */,
  32'h3d2d543a /* (0, 4, 13) */,
  32'h3d2d543a /* (28, 0, 13) */,
  32'h3d7388b1 /* (24, 0, 13) */,
  32'h3dccb681 /* (20, 0, 13) */,
  32'h3de8675d /* (16, 0, 13) */,
  32'h3dccb681 /* (12, 0, 13) */,
  32'h3d7388b1 /* (8, 0, 13) */,
  32'h3d2d543a /* (4, 0, 13) */,
  32'h3d1c4c09 /* (0, 0, 13) */,
  32'h3d19e157 /* (28, 28, 9) */,
  32'h3d3f1eea /* (24, 28, 9) */,
  32'h3d902ce0 /* (20, 28, 9) */,
  32'h3d97bb42 /* (16, 28, 9) */,
  32'h3d902ce0 /* (12, 28, 9) */,
  32'h3d3f1eea /* (8, 28, 9) */,
  32'h3d19e157 /* (4, 28, 9) */,
  32'h3d13aacb /* (0, 28, 9) */,
  32'h3d3f1eea /* (28, 24, 9) */,
  32'h3d824402 /* (24, 24, 9) */,
  32'h3dd4c19e /* (20, 24, 9) */,
  32'h3dec5cc9 /* (16, 24, 9) */,
  32'h3dd4c19e /* (12, 24, 9) */,
  32'h3d824402 /* (8, 24, 9) */,
  32'h3d3f1eea /* (4, 24, 9) */,
  32'h3d2eceba /* (0, 24, 9) */,
  32'h3d902ce0 /* (28, 20, 9) */,
  32'h3dd4c19e /* (24, 20, 9) */,
  32'h3e3c290c /* (20, 20, 9) */,
  32'h3e5e82df /* (16, 20, 9) */,
  32'h3e3c290c /* (12, 20, 9) */,
  32'h3dd4c19e /* (8, 20, 9) */,
  32'h3d902ce0 /* (4, 20, 9) */,
  32'h3d7e6b4b /* (0, 20, 9) */,
  32'h3d97bb42 /* (28, 16, 9) */,
  32'h3dec5cc9 /* (24, 16, 9) */,
  32'h3e5e82df /* (20, 16, 9) */,
  32'h3e8b1bdf /* (16, 16, 9) */,
  32'h3e5e82df /* (12, 16, 9) */,
  32'h3dec5cc9 /* (8, 16, 9) */,
  32'h3d97bb42 /* (4, 16, 9) */,
  32'h3d82ec35 /* (0, 16, 9) */,
  32'h3d902ce0 /* (28, 12, 9) */,
  32'h3dd4c19e /* (24, 12, 9) */,
  32'h3e3c290c /* (20, 12, 9) */,
  32'h3e5e82df /* (16, 12, 9) */,
  32'h3e3c290c /* (12, 12, 9) */,
  32'h3dd4c19e /* (8, 12, 9) */,
  32'h3d902ce0 /* (4, 12, 9) */,
  32'h3d7e6b4b /* (0, 12, 9) */,
  32'h3d3f1eea /* (28, 8, 9) */,
  32'h3d824402 /* (24, 8, 9) */,
  32'h3dd4c19e /* (20, 8, 9) */,
  32'h3dec5cc9 /* (16, 8, 9) */,
  32'h3dd4c19e /* (12, 8, 9) */,
  32'h3d824402 /* (8, 8, 9) */,
  32'h3d3f1eea /* (4, 8, 9) */,
  32'h3d2eceba /* (0, 8, 9) */,
  32'h3d19e157 /* (28, 4, 9) */,
  32'h3d3f1eea /* (24, 4, 9) */,
  32'h3d902ce0 /* (20, 4, 9) */,
  32'h3d97bb42 /* (16, 4, 9) */,
  32'h3d902ce0 /* (12, 4, 9) */,
  32'h3d3f1eea /* (8, 4, 9) */,
  32'h3d19e157 /* (4, 4, 9) */,
  32'h3d13aacb /* (0, 4, 9) */,
  32'h3d13aacb /* (28, 0, 9) */,
  32'h3d2eceba /* (24, 0, 9) */,
  32'h3d7e6b4b /* (20, 0, 9) */,
  32'h3d82ec35 /* (16, 0, 9) */,
  32'h3d7e6b4b /* (12, 0, 9) */,
  32'h3d2eceba /* (8, 0, 9) */,
  32'h3d13aacb /* (4, 0, 9) */,
  32'h3d11ab15 /* (0, 0, 9) */,
  32'h3d1e7527 /* (28, 28, 5) */,
  32'h3d183845 /* (24, 28, 5) */,
  32'h3d431db1 /* (20, 28, 5) */,
  32'h3d3b5943 /* (16, 28, 5) */,
  32'h3d431db1 /* (12, 28, 5) */,
  32'h3d183845 /* (8, 28, 5) */,
  32'h3d1e7527 /* (4, 28, 5) */,
  32'h3d3577a5 /* (0, 28, 5) */,
  32'h3d183845 /* (28, 24, 5) */,
  32'h3d38dbff /* (24, 24, 5) */,
  32'h3d89129f /* (20, 24, 5) */,
  32'h3d8eb3bf /* (16, 24, 5) */,
  32'h3d89129f /* (12, 24, 5) */,
  32'h3d38dbff /* (8, 24, 5) */,
  32'h3d183845 /* (4, 24, 5) */,
  32'h3d13eed3 /* (0, 24, 5) */,
  32'h3d431db1 /* (28, 20, 5) */,
  32'h3d89129f /* (24, 20, 5) */,
  32'h3de671da /* (20, 20, 5) */,
  32'h3e02cee2 /* (16, 20, 5) */,
  32'h3de671da /* (12, 20, 5) */,
  32'h3d89129f /* (8, 20, 5) */,
  32'h3d431db1 /* (4, 20, 5) */,
  32'h3d2ff16f /* (0, 20, 5) */,
  32'h3d3b5943 /* (28, 16, 5) */,
  32'h3d8eb3bf /* (24, 16, 5) */,
  32'h3e02cee2 /* (20, 16, 5) */,
  32'h3e1f95bf /* (16, 16, 5) */,
  32'h3e02cee2 /* (12, 16, 5) */,
  32'h3d8eb3bf /* (8, 16, 5) */,
  32'h3d3b5943 /* (4, 16, 5) */,
  32'h3d231d8f /* (0, 16, 5) */,
  32'h3d431db1 /* (28, 12, 5) */,
  32'h3d89129f /* (24, 12, 5) */,
  32'h3de671da /* (20, 12, 5) */,
  32'h3e02cee2 /* (16, 12, 5) */,
  32'h3de671da /* (12, 12, 5) */,
  32'h3d89129f /* (8, 12, 5) */,
  32'h3d431db1 /* (4, 12, 5) */,
  32'h3d2ff16f /* (0, 12, 5) */,
  32'h3d183845 /* (28, 8, 5) */,
  32'h3d38dbff /* (24, 8, 5) */,
  32'h3d89129f /* (20, 8, 5) */,
  32'h3d8eb3bf /* (16, 8, 5) */,
  32'h3d89129f /* (12, 8, 5) */,
  32'h3d38dbff /* (8, 8, 5) */,
  32'h3d183845 /* (4, 8, 5) */,
  32'h3d13eed3 /* (0, 8, 5) */,
  32'h3d1e7527 /* (28, 4, 5) */,
  32'h3d183845 /* (24, 4, 5) */,
  32'h3d431db1 /* (20, 4, 5) */,
  32'h3d3b5943 /* (16, 4, 5) */,
  32'h3d431db1 /* (12, 4, 5) */,
  32'h3d183845 /* (8, 4, 5) */,
  32'h3d1e7527 /* (4, 4, 5) */,
  32'h3d3577a5 /* (0, 4, 5) */,
  32'h3d3577a5 /* (28, 0, 5) */,
  32'h3d13eed3 /* (24, 0, 5) */,
  32'h3d2ff16f /* (20, 0, 5) */,
  32'h3d231d8f /* (16, 0, 5) */,
  32'h3d2ff16f /* (12, 0, 5) */,
  32'h3d13eed3 /* (8, 0, 5) */,
  32'h3d3577a5 /* (4, 0, 5) */,
  32'h3d75271a /* (0, 0, 5) */,
  32'h3d4cb45d /* (28, 28, 1) */,
  32'h3d139499 /* (24, 28, 1) */,
  32'h3d27af27 /* (20, 28, 1) */,
  32'h3d18708b /* (16, 28, 1) */,
  32'h3d27af27 /* (12, 28, 1) */,
  32'h3d139499 /* (8, 28, 1) */,
  32'h3d4cb45d /* (4, 28, 1) */,
  32'h3da3aa58 /* (0, 28, 1) */,
  32'h3d139499 /* (28, 24, 1) */,
  32'h3d23fb6f /* (24, 24, 1) */,
  32'h3d649547 /* (20, 24, 1) */,
  32'h3d656b11 /* (16, 24, 1) */,
  32'h3d649547 /* (12, 24, 1) */,
  32'h3d23fb6f /* (8, 24, 1) */,
  32'h3d139499 /* (4, 24, 1) */,
  32'h3d177e6a /* (0, 24, 1) */,
  32'h3d27af27 /* (28, 20, 1) */,
  32'h3d649547 /* (24, 20, 1) */,
  32'h3dbaaaa9 /* (20, 20, 1) */,
  32'h3dcf60c6 /* (16, 20, 1) */,
  32'h3dbaaaa9 /* (12, 20, 1) */,
  32'h3d649547 /* (8, 20, 1) */,
  32'h3d27af27 /* (4, 20, 1) */,
  32'h3d195f14 /* (0, 20, 1) */,
  32'h3d18708b /* (28, 16, 1) */,
  32'h3d656b11 /* (24, 16, 1) */,
  32'h3dcf60c6 /* (20, 16, 1) */,
  32'h3df9e164 /* (16, 16, 1) */,
  32'h3dcf60c6 /* (12, 16, 1) */,
  32'h3d656b11 /* (8, 16, 1) */,
  32'h3d18708b /* (4, 16, 1) */,
  32'h3d0563b9 /* (0, 16, 1) */,
  32'h3d27af27 /* (28, 12, 1) */,
  32'h3d649547 /* (24, 12, 1) */,
  32'h3dbaaaa9 /* (20, 12, 1) */,
  32'h3dcf60c6 /* (16, 12, 1) */,
  32'h3dbaaaa9 /* (12, 12, 1) */,
  32'h3d649547 /* (8, 12, 1) */,
  32'h3d27af27 /* (4, 12, 1) */,
  32'h3d195f14 /* (0, 12, 1) */,
  32'h3d139499 /* (28, 8, 1) */,
  32'h3d23fb6f /* (24, 8, 1) */,
  32'h3d649547 /* (20, 8, 1) */,
  32'h3d656b11 /* (16, 8, 1) */,
  32'h3d649547 /* (12, 8, 1) */,
  32'h3d23fb6f /* (8, 8, 1) */,
  32'h3d139499 /* (4, 8, 1) */,
  32'h3d177e6a /* (0, 8, 1) */,
  32'h3d4cb45d /* (28, 4, 1) */,
  32'h3d139499 /* (24, 4, 1) */,
  32'h3d27af27 /* (20, 4, 1) */,
  32'h3d18708b /* (16, 4, 1) */,
  32'h3d27af27 /* (12, 4, 1) */,
  32'h3d139499 /* (8, 4, 1) */,
  32'h3d4cb45d /* (4, 4, 1) */,
  32'h3da3aa58 /* (0, 4, 1) */,
  32'h3da3aa58 /* (28, 0, 1) */,
  32'h3d177e6a /* (24, 0, 1) */,
  32'h3d195f14 /* (20, 0, 1) */,
  32'h3d0563b9 /* (16, 0, 1) */,
  32'h3d195f14 /* (12, 0, 1) */,
  32'h3d177e6a /* (8, 0, 1) */,
  32'h3da3aa58 /* (4, 0, 1) */,
  32'h3f8f3ec8 /* (0, 0, 1) */,
  32'h3d9c757b /* (31, 31, 28) */,
  32'h3d334ee4 /* (27, 31, 28) */,
  32'h3d13f199 /* (23, 31, 28) */,
  32'h3d2e802a /* (19, 31, 28) */,
  32'h3d294c4b /* (15, 31, 28) */,
  32'h3d1f5dc3 /* (11, 31, 28) */,
  32'h3d17ff6b /* (7, 31, 28) */,
  32'h3d6eb36b /* (3, 31, 28) */,
  32'h3d334ee4 /* (31, 27, 28) */,
  32'h3d189061 /* (27, 27, 28) */,
  32'h3d1ee50b /* (23, 27, 28) */,
  32'h3d4ea6a0 /* (19, 27, 28) */,
  32'h3d4def9b /* (15, 27, 28) */,
  32'h3d358341 /* (11, 27, 28) */,
  32'h3d1508af /* (7, 27, 28) */,
  32'h3d25f5ce /* (3, 27, 28) */,
  32'h3d13f199 /* (31, 23, 28) */,
  32'h3d1ee50b /* (27, 23, 28) */,
  32'h3d51a9d2 /* (23, 23, 28) */,
  32'h3d9d0afa /* (19, 23, 28) */,
  32'h3da3c1ed /* (15, 23, 28) */,
  32'h3d81d711 /* (11, 23, 28) */,
  32'h3d30de15 /* (7, 23, 28) */,
  32'h3d16b5b2 /* (3, 23, 28) */,
  32'h3d2e802a /* (31, 19, 28) */,
  32'h3d4ea6a0 /* (27, 19, 28) */,
  32'h3d9d0afa /* (23, 19, 28) */,
  32'h3e0415cb /* (19, 19, 28) */,
  32'h3e0ff4ce /* (15, 19, 28) */,
  32'h3dcf13a3 /* (11, 19, 28) */,
  32'h3d770afc /* (7, 19, 28) */,
  32'h3d385879 /* (3, 19, 28) */,
  32'h3d294c4b /* (31, 15, 28) */,
  32'h3d4def9b /* (27, 15, 28) */,
  32'h3da3c1ed /* (23, 15, 28) */,
  32'h3e0ff4ce /* (19, 15, 28) */,
  32'h3e1fe07e /* (15, 15, 28) */,
  32'h3ddcf428 /* (11, 15, 28) */,
  32'h3d7b9f11 /* (7, 15, 28) */,
  32'h3d349293 /* (3, 15, 28) */,
  32'h3d1f5dc3 /* (31, 11, 28) */,
  32'h3d358341 /* (27, 11, 28) */,
  32'h3d81d711 /* (23, 11, 28) */,
  32'h3dcf13a3 /* (19, 11, 28) */,
  32'h3ddcf428 /* (15, 11, 28) */,
  32'h3da66ad4 /* (11, 11, 28) */,
  32'h3d52976b /* (7, 11, 28) */,
  32'h3d25fa09 /* (3, 11, 28) */,
  32'h3d17ff6b /* (31, 7, 28) */,
  32'h3d1508af /* (27, 7, 28) */,
  32'h3d30de15 /* (23, 7, 28) */,
  32'h3d770afc /* (19, 7, 28) */,
  32'h3d7b9f11 /* (15, 7, 28) */,
  32'h3d52976b /* (11, 7, 28) */,
  32'h3d1cbb18 /* (7, 7, 28) */,
  32'h3d155fa4 /* (3, 7, 28) */,
  32'h3d6eb36b /* (31, 3, 28) */,
  32'h3d25f5ce /* (27, 3, 28) */,
  32'h3d16b5b2 /* (23, 3, 28) */,
  32'h3d385879 /* (19, 3, 28) */,
  32'h3d349293 /* (15, 3, 28) */,
  32'h3d25fa09 /* (11, 3, 28) */,
  32'h3d155fa4 /* (7, 3, 28) */,
  32'h3d4920d0 /* (3, 3, 28) */,
  32'h3d1704d7 /* (31, 31, 24) */,
  32'h3d1412fd /* (27, 31, 24) */,
  32'h3d2fba80 /* (23, 31, 24) */,
  32'h3d7573b6 /* (19, 31, 24) */,
  32'h3d7a003f /* (15, 31, 24) */,
  32'h3d513c3d /* (11, 31, 24) */,
  32'h3d1bb8b6 /* (7, 31, 24) */,
  32'h3d146963 /* (3, 31, 24) */,
  32'h3d1412fd /* (31, 27, 24) */,
  32'h3d1c4d38 /* (27, 27, 24) */,
  32'h3d49c96c /* (23, 27, 24) */,
  32'h3d94d380 /* (19, 27, 24) */,
  32'h3d9a5b6b /* (15, 27, 24) */,
  32'h3d77c8fd /* (11, 27, 24) */,
  32'h3d2bff3e /* (7, 27, 24) */,
  32'h3d15d660 /* (3, 27, 24) */,
  32'h3d2fba80 /* (31, 23, 24) */,
  32'h3d49c96c /* (27, 23, 24) */,
  32'h3d921bde /* (23, 23, 24) */,
  32'h3deb6b6d /* (19, 23, 24) */,
  32'h3dfc30a3 /* (15, 23, 24) */,
  32'h3dbc4d73 /* (11, 23, 24) */,
  32'h3d6b8b35 /* (7, 23, 24) */,
  32'h3d37919e /* (3, 23, 24) */,
  32'h3d7573b6 /* (31, 19, 24) */,
  32'h3d94d380 /* (27, 19, 24) */,
  32'h3deb6b6d /* (23, 19, 24) */,
  32'h3e4dd3dc /* (19, 19, 24) */,
  32'h3e640ba2 /* (15, 19, 24) */,
  32'h3e1e607d /* (11, 19, 24) */,
  32'h3db56072 /* (7, 19, 24) */,
  32'h3d82c188 /* (3, 19, 24) */,
  32'h3d7a003f /* (31, 15, 24) */,
  32'h3d9a5b6b /* (27, 15, 24) */,
  32'h3dfc30a3 /* (23, 15, 24) */,
  32'h3e640ba2 /* (19, 15, 24) */,
  32'h3e803f85 /* (15, 15, 24) */,
  32'h3e2c9c6c /* (11, 15, 24) */,
  32'h3dbf0444 /* (7, 15, 24) */,
  32'h3d8608f0 /* (3, 15, 24) */,
  32'h3d513c3d /* (31, 11, 24) */,
  32'h3d77c8fd /* (27, 11, 24) */,
  32'h3dbc4d73 /* (23, 11, 24) */,
  32'h3e1e607d /* (19, 11, 24) */,
  32'h3e2c9c6c /* (15, 11, 24) */,
  32'h3df84bb3 /* (11, 11, 24) */,
  32'h3d941bce /* (7, 11, 24) */,
  32'h3d5d0a38 /* (3, 11, 24) */,
  32'h3d1bb8b6 /* (31, 7, 24) */,
  32'h3d2bff3e /* (27, 7, 24) */,
  32'h3d6b8b35 /* (23, 7, 24) */,
  32'h3db56072 /* (19, 7, 24) */,
  32'h3dbf0444 /* (15, 7, 24) */,
  32'h3d941bce /* (11, 7, 24) */,
  32'h3d432bf1 /* (7, 7, 24) */,
  32'h3d2054cd /* (3, 7, 24) */,
  32'h3d146963 /* (31, 3, 24) */,
  32'h3d15d660 /* (27, 3, 24) */,
  32'h3d37919e /* (23, 3, 24) */,
  32'h3d82c188 /* (19, 3, 24) */,
  32'h3d8608f0 /* (15, 3, 24) */,
  32'h3d5d0a38 /* (11, 3, 24) */,
  32'h3d2054cd /* (7, 3, 24) */,
  32'h3d1392fe /* (3, 3, 24) */,
  32'h3d1a2df1 /* (31, 31, 20) */,
  32'h3d310ad3 /* (27, 31, 20) */,
  32'h3d803124 /* (23, 31, 20) */,
  32'h3dce8d02 /* (19, 31, 20) */,
  32'h3ddd43c2 /* (15, 31, 20) */,
  32'h3da53628 /* (11, 31, 20) */,
  32'h3d4ea8e5 /* (7, 31, 20) */,
  32'h3d210eee /* (3, 31, 20) */,
  32'h3d310ad3 /* (31, 27, 20) */,
  32'h3d4f6dfc /* (27, 27, 20) */,
  32'h3d9af1c2 /* (23, 27, 20) */,
  32'h3e00477d /* (19, 27, 20) */,
  32'h3e0ae903 /* (15, 27, 20) */,
  32'h3dca9d53 /* (11, 27, 20) */,
  32'h3d75e4d4 /* (7, 27, 20) */,
  32'h3d3a4ebb /* (3, 27, 20) */,
  32'h3d803124 /* (31, 23, 20) */,
  32'h3d9af1c2 /* (27, 23, 20) */,
  32'h3df3b4f2 /* (23, 23, 20) */,
  32'h3e53dc51 /* (19, 23, 20) */,
  32'h3e6a25fd /* (15, 23, 20) */,
  32'h3e23781b /* (11, 23, 20) */,
  32'h3dbc51f9 /* (7, 23, 20) */,
  32'h3d886b82 /* (3, 23, 20) */,
  32'h3dce8d02 /* (31, 19, 20) */,
  32'h3e00477d /* (27, 19, 20) */,
  32'h3e53dc51 /* (23, 19, 20) */,
  32'h3ec1d890 /* (19, 19, 20) */,
  32'h3edb3822 /* (15, 19, 20) */,
  32'h3e91dfe2 /* (11, 19, 20) */,
  32'h3e1f8cbf /* (7, 19, 20) */,
  32'h3dddef48 /* (3, 19, 20) */,
  32'h3ddd43c2 /* (31, 15, 20) */,
  32'h3e0ae903 /* (27, 15, 20) */,
  32'h3e6a25fd /* (23, 15, 20) */,
  32'h3edb3822 /* (19, 15, 20) */,
  32'h3efaa119 /* (15, 15, 20) */,
  32'h3ea31756 /* (11, 15, 20) */,
  32'h3e2e6a71 /* (7, 15, 20) */,
  32'h3deea44d /* (3, 15, 20) */,
  32'h3da53628 /* (31, 11, 20) */,
  32'h3dca9d53 /* (27, 11, 20) */,
  32'h3e23781b /* (23, 11, 20) */,
  32'h3e91dfe2 /* (19, 11, 20) */,
  32'h3ea31756 /* (15, 11, 20) */,
  32'h3e5e44ac /* (11, 11, 20) */,
  32'h3df94537 /* (7, 11, 20) */,
  32'h3db0b965 /* (3, 11, 20) */,
  32'h3d4ea8e5 /* (31, 7, 20) */,
  32'h3d75e4d4 /* (27, 7, 20) */,
  32'h3dbc51f9 /* (23, 7, 20) */,
  32'h3e1f8cbf /* (19, 7, 20) */,
  32'h3e2e6a71 /* (15, 7, 20) */,
  32'h3df94537 /* (11, 7, 20) */,
  32'h3d938890 /* (7, 7, 20) */,
  32'h3d5ab0e1 /* (3, 7, 20) */,
  32'h3d210eee /* (31, 3, 20) */,
  32'h3d3a4ebb /* (27, 3, 20) */,
  32'h3d886b82 /* (23, 3, 20) */,
  32'h3dddef48 /* (19, 3, 20) */,
  32'h3deea44d /* (15, 3, 20) */,
  32'h3db0b965 /* (11, 3, 20) */,
  32'h3d5ab0e1 /* (7, 3, 20) */,
  32'h3d28b308 /* (3, 3, 20) */,
  32'h3d067e68 /* (31, 31, 16) */,
  32'h3d24852f /* (27, 31, 16) */,
  32'h3d8420c9 /* (23, 31, 16) */,
  32'h3deaafef /* (19, 31, 16) */,
  32'h3e02e976 /* (15, 31, 16) */,
  32'h3db336e0 /* (11, 31, 16) */,
  32'h3d49f75a /* (7, 31, 16) */,
  32'h3d0fbc59 /* (3, 31, 16) */,
  32'h3d24852f /* (31, 27, 16) */,
  32'h3d4ab7f7 /* (27, 27, 16) */,
  32'h3da4f2f4 /* (23, 27, 16) */,
  32'h3e1486b7 /* (19, 27, 16) */,
  32'h3e26bbbb /* (15, 27, 16) */,
  32'h3de14ffa /* (11, 27, 16) */,
  32'h3d7a662c /* (7, 27, 16) */,
  32'h3d3046d8 /* (3, 27, 16) */,
  32'h3d8420c9 /* (31, 23, 16) */,
  32'h3da4f2f4 /* (27, 23, 16) */,
  32'h3e0981d7 /* (23, 23, 16) */,
  32'h3e7e4b9d /* (19, 23, 16) */,
  32'h3e908107 /* (15, 23, 16) */,
  32'h3e3e5da7 /* (11, 23, 16) */,
  32'h3dce1075 /* (7, 23, 16) */,
  32'h3d8e3848 /* (3, 23, 16) */,
  32'h3deaafef /* (31, 19, 16) */,
  32'h3e1486b7 /* (27, 19, 16) */,
  32'h3e7e4b9d /* (23, 19, 16) */,
  32'h3ef27895 /* (19, 19, 16) */,
  32'h3f0bd969 /* (15, 19, 16) */,
  32'h3eb2bd2a /* (11, 19, 16) */,
  32'h3e3bd4ee /* (7, 19, 16) */,
  32'h3dfdd31f /* (3, 19, 16) */,
  32'h3e02e976 /* (31, 15, 16) */,
  32'h3e26bbbb /* (27, 15, 16) */,
  32'h3e908107 /* (23, 15, 16) */,
  32'h3f0bd969 /* (19, 15, 16) */,
  32'h3f2286f8 /* (15, 15, 16) */,
  32'h3ecca1ac /* (11, 15, 16) */,
  32'h3e540b9b /* (7, 15, 16) */,
  32'h3e0de417 /* (3, 15, 16) */,
  32'h3db336e0 /* (31, 11, 16) */,
  32'h3de14ffa /* (27, 11, 16) */,
  32'h3e3e5da7 /* (23, 11, 16) */,
  32'h3eb2bd2a /* (19, 11, 16) */,
  32'h3ecca1ac /* (15, 11, 16) */,
  32'h3e84c8e0 /* (11, 11, 16) */,
  32'h3e0d9cf0 /* (7, 11, 16) */,
  32'h3dc1602b /* (3, 11, 16) */,
  32'h3d49f75a /* (31, 7, 16) */,
  32'h3d7a662c /* (27, 7, 16) */,
  32'h3dce1075 /* (23, 7, 16) */,
  32'h3e3bd4ee /* (19, 7, 16) */,
  32'h3e540b9b /* (15, 7, 16) */,
  32'h3e0d9cf0 /* (11, 7, 16) */,
  32'h3d9b7830 /* (7, 7, 16) */,
  32'h3d58de26 /* (3, 7, 16) */,
  32'h3d0fbc59 /* (31, 3, 16) */,
  32'h3d3046d8 /* (27, 3, 16) */,
  32'h3d8e3848 /* (23, 3, 16) */,
  32'h3dfdd31f /* (19, 3, 16) */,
  32'h3e0de417 /* (15, 3, 16) */,
  32'h3dc1602b /* (11, 3, 16) */,
  32'h3d58de26 /* (7, 3, 16) */,
  32'h3d19c07a /* (3, 3, 16) */,
  32'h3d1a2df1 /* (31, 31, 12) */,
  32'h3d310ad3 /* (27, 31, 12) */,
  32'h3d803124 /* (23, 31, 12) */,
  32'h3dce8d02 /* (19, 31, 12) */,
  32'h3ddd43c2 /* (15, 31, 12) */,
  32'h3da53628 /* (11, 31, 12) */,
  32'h3d4ea8e5 /* (7, 31, 12) */,
  32'h3d210eee /* (3, 31, 12) */,
  32'h3d310ad3 /* (31, 27, 12) */,
  32'h3d4f6dfc /* (27, 27, 12) */,
  32'h3d9af1c2 /* (23, 27, 12) */,
  32'h3e00477d /* (19, 27, 12) */,
  32'h3e0ae903 /* (15, 27, 12) */,
  32'h3dca9d53 /* (11, 27, 12) */,
  32'h3d75e4d4 /* (7, 27, 12) */,
  32'h3d3a4ebb /* (3, 27, 12) */,
  32'h3d803124 /* (31, 23, 12) */,
  32'h3d9af1c2 /* (27, 23, 12) */,
  32'h3df3b4f2 /* (23, 23, 12) */,
  32'h3e53dc51 /* (19, 23, 12) */,
  32'h3e6a25fd /* (15, 23, 12) */,
  32'h3e23781b /* (11, 23, 12) */,
  32'h3dbc51f9 /* (7, 23, 12) */,
  32'h3d886b82 /* (3, 23, 12) */,
  32'h3dce8d02 /* (31, 19, 12) */,
  32'h3e00477d /* (27, 19, 12) */,
  32'h3e53dc51 /* (23, 19, 12) */,
  32'h3ec1d890 /* (19, 19, 12) */,
  32'h3edb3822 /* (15, 19, 12) */,
  32'h3e91dfe2 /* (11, 19, 12) */,
  32'h3e1f8cbf /* (7, 19, 12) */,
  32'h3dddef48 /* (3, 19, 12) */,
  32'h3ddd43c2 /* (31, 15, 12) */,
  32'h3e0ae903 /* (27, 15, 12) */,
  32'h3e6a25fd /* (23, 15, 12) */,
  32'h3edb3822 /* (19, 15, 12) */,
  32'h3efaa119 /* (15, 15, 12) */,
  32'h3ea31756 /* (11, 15, 12) */,
  32'h3e2e6a71 /* (7, 15, 12) */,
  32'h3deea44d /* (3, 15, 12) */,
  32'h3da53628 /* (31, 11, 12) */,
  32'h3dca9d53 /* (27, 11, 12) */,
  32'h3e23781b /* (23, 11, 12) */,
  32'h3e91dfe2 /* (19, 11, 12) */,
  32'h3ea31756 /* (15, 11, 12) */,
  32'h3e5e44ac /* (11, 11, 12) */,
  32'h3df94537 /* (7, 11, 12) */,
  32'h3db0b965 /* (3, 11, 12) */,
  32'h3d4ea8e5 /* (31, 7, 12) */,
  32'h3d75e4d4 /* (27, 7, 12) */,
  32'h3dbc51f9 /* (23, 7, 12) */,
  32'h3e1f8cbf /* (19, 7, 12) */,
  32'h3e2e6a71 /* (15, 7, 12) */,
  32'h3df94537 /* (11, 7, 12) */,
  32'h3d938890 /* (7, 7, 12) */,
  32'h3d5ab0e1 /* (3, 7, 12) */,
  32'h3d210eee /* (31, 3, 12) */,
  32'h3d3a4ebb /* (27, 3, 12) */,
  32'h3d886b82 /* (23, 3, 12) */,
  32'h3dddef48 /* (19, 3, 12) */,
  32'h3deea44d /* (15, 3, 12) */,
  32'h3db0b965 /* (11, 3, 12) */,
  32'h3d5ab0e1 /* (7, 3, 12) */,
  32'h3d28b308 /* (3, 3, 12) */,
  32'h3d1704d7 /* (31, 31, 8) */,
  32'h3d1412fd /* (27, 31, 8) */,
  32'h3d2fba80 /* (23, 31, 8) */,
  32'h3d7573b6 /* (19, 31, 8) */,
  32'h3d7a003f /* (15, 31, 8) */,
  32'h3d513c3d /* (11, 31, 8) */,
  32'h3d1bb8b6 /* (7, 31, 8) */,
  32'h3d146963 /* (3, 31, 8) */,
  32'h3d1412fd /* (31, 27, 8) */,
  32'h3d1c4d38 /* (27, 27, 8) */,
  32'h3d49c96c /* (23, 27, 8) */,
  32'h3d94d380 /* (19, 27, 8) */,
  32'h3d9a5b6b /* (15, 27, 8) */,
  32'h3d77c8fd /* (11, 27, 8) */,
  32'h3d2bff3e /* (7, 27, 8) */,
  32'h3d15d660 /* (3, 27, 8) */,
  32'h3d2fba80 /* (31, 23, 8) */,
  32'h3d49c96c /* (27, 23, 8) */,
  32'h3d921bde /* (23, 23, 8) */,
  32'h3deb6b6d /* (19, 23, 8) */,
  32'h3dfc30a3 /* (15, 23, 8) */,
  32'h3dbc4d73 /* (11, 23, 8) */,
  32'h3d6b8b35 /* (7, 23, 8) */,
  32'h3d37919e /* (3, 23, 8) */,
  32'h3d7573b6 /* (31, 19, 8) */,
  32'h3d94d380 /* (27, 19, 8) */,
  32'h3deb6b6d /* (23, 19, 8) */,
  32'h3e4dd3dc /* (19, 19, 8) */,
  32'h3e640ba2 /* (15, 19, 8) */,
  32'h3e1e607d /* (11, 19, 8) */,
  32'h3db56072 /* (7, 19, 8) */,
  32'h3d82c188 /* (3, 19, 8) */,
  32'h3d7a003f /* (31, 15, 8) */,
  32'h3d9a5b6b /* (27, 15, 8) */,
  32'h3dfc30a3 /* (23, 15, 8) */,
  32'h3e640ba2 /* (19, 15, 8) */,
  32'h3e803f85 /* (15, 15, 8) */,
  32'h3e2c9c6c /* (11, 15, 8) */,
  32'h3dbf0444 /* (7, 15, 8) */,
  32'h3d8608f0 /* (3, 15, 8) */,
  32'h3d513c3d /* (31, 11, 8) */,
  32'h3d77c8fd /* (27, 11, 8) */,
  32'h3dbc4d73 /* (23, 11, 8) */,
  32'h3e1e607d /* (19, 11, 8) */,
  32'h3e2c9c6c /* (15, 11, 8) */,
  32'h3df84bb3 /* (11, 11, 8) */,
  32'h3d941bce /* (7, 11, 8) */,
  32'h3d5d0a38 /* (3, 11, 8) */,
  32'h3d1bb8b6 /* (31, 7, 8) */,
  32'h3d2bff3e /* (27, 7, 8) */,
  32'h3d6b8b35 /* (23, 7, 8) */,
  32'h3db56072 /* (19, 7, 8) */,
  32'h3dbf0444 /* (15, 7, 8) */,
  32'h3d941bce /* (11, 7, 8) */,
  32'h3d432bf1 /* (7, 7, 8) */,
  32'h3d2054cd /* (3, 7, 8) */,
  32'h3d146963 /* (31, 3, 8) */,
  32'h3d15d660 /* (27, 3, 8) */,
  32'h3d37919e /* (23, 3, 8) */,
  32'h3d82c188 /* (19, 3, 8) */,
  32'h3d8608f0 /* (15, 3, 8) */,
  32'h3d5d0a38 /* (11, 3, 8) */,
  32'h3d2054cd /* (7, 3, 8) */,
  32'h3d1392fe /* (3, 3, 8) */,
  32'h3d9c757b /* (31, 31, 4) */,
  32'h3d334ee4 /* (27, 31, 4) */,
  32'h3d13f199 /* (23, 31, 4) */,
  32'h3d2e802a /* (19, 31, 4) */,
  32'h3d294c4b /* (15, 31, 4) */,
  32'h3d1f5dc3 /* (11, 31, 4) */,
  32'h3d17ff6b /* (7, 31, 4) */,
  32'h3d6eb36b /* (3, 31, 4) */,
  32'h3d334ee4 /* (31, 27, 4) */,
  32'h3d189061 /* (27, 27, 4) */,
  32'h3d1ee50b /* (23, 27, 4) */,
  32'h3d4ea6a0 /* (19, 27, 4) */,
  32'h3d4def9b /* (15, 27, 4) */,
  32'h3d358341 /* (11, 27, 4) */,
  32'h3d1508af /* (7, 27, 4) */,
  32'h3d25f5ce /* (3, 27, 4) */,
  32'h3d13f199 /* (31, 23, 4) */,
  32'h3d1ee50b /* (27, 23, 4) */,
  32'h3d51a9d2 /* (23, 23, 4) */,
  32'h3d9d0afa /* (19, 23, 4) */,
  32'h3da3c1ed /* (15, 23, 4) */,
  32'h3d81d711 /* (11, 23, 4) */,
  32'h3d30de15 /* (7, 23, 4) */,
  32'h3d16b5b2 /* (3, 23, 4) */,
  32'h3d2e802a /* (31, 19, 4) */,
  32'h3d4ea6a0 /* (27, 19, 4) */,
  32'h3d9d0afa /* (23, 19, 4) */,
  32'h3e0415cb /* (19, 19, 4) */,
  32'h3e0ff4ce /* (15, 19, 4) */,
  32'h3dcf13a3 /* (11, 19, 4) */,
  32'h3d770afc /* (7, 19, 4) */,
  32'h3d385879 /* (3, 19, 4) */,
  32'h3d294c4b /* (31, 15, 4) */,
  32'h3d4def9b /* (27, 15, 4) */,
  32'h3da3c1ed /* (23, 15, 4) */,
  32'h3e0ff4ce /* (19, 15, 4) */,
  32'h3e1fe07e /* (15, 15, 4) */,
  32'h3ddcf428 /* (11, 15, 4) */,
  32'h3d7b9f11 /* (7, 15, 4) */,
  32'h3d349293 /* (3, 15, 4) */,
  32'h3d1f5dc3 /* (31, 11, 4) */,
  32'h3d358341 /* (27, 11, 4) */,
  32'h3d81d711 /* (23, 11, 4) */,
  32'h3dcf13a3 /* (19, 11, 4) */,
  32'h3ddcf428 /* (15, 11, 4) */,
  32'h3da66ad4 /* (11, 11, 4) */,
  32'h3d52976b /* (7, 11, 4) */,
  32'h3d25fa09 /* (3, 11, 4) */,
  32'h3d17ff6b /* (31, 7, 4) */,
  32'h3d1508af /* (27, 7, 4) */,
  32'h3d30de15 /* (23, 7, 4) */,
  32'h3d770afc /* (19, 7, 4) */,
  32'h3d7b9f11 /* (15, 7, 4) */,
  32'h3d52976b /* (11, 7, 4) */,
  32'h3d1cbb18 /* (7, 7, 4) */,
  32'h3d155fa4 /* (3, 7, 4) */,
  32'h3d6eb36b /* (31, 3, 4) */,
  32'h3d25f5ce /* (27, 3, 4) */,
  32'h3d16b5b2 /* (23, 3, 4) */,
  32'h3d385879 /* (19, 3, 4) */,
  32'h3d349293 /* (15, 3, 4) */,
  32'h3d25fa09 /* (11, 3, 4) */,
  32'h3d155fa4 /* (7, 3, 4) */,
  32'h3d4920d0 /* (3, 3, 4) */,
  32'h3f10fe39 /* (31, 31, 0) */,
  32'h3d6e9998 /* (27, 31, 0) */,
  32'h3d11a5c6 /* (23, 31, 0) */,
  32'h3d1d4601 /* (19, 31, 0) */,
  32'h3d155505 /* (15, 31, 0) */,
  32'h3d147e90 /* (11, 31, 0) */,
  32'h3d25463b /* (7, 31, 0) */,
  32'h3dff9e3f /* (3, 31, 0) */,
  32'h3d6e9998 /* (31, 27, 0) */,
  32'h3d25e3da /* (27, 27, 0) */,
  32'h3d16a564 /* (23, 27, 0) */,
  32'h3d384488 /* (19, 27, 0) */,
  32'h3d347f0a /* (15, 27, 0) */,
  32'h3d25e815 /* (11, 27, 0) */,
  32'h3d154f7b /* (7, 27, 0) */,
  32'h3d490b0e /* (3, 27, 0) */,
  32'h3d11a5c6 /* (31, 23, 0) */,
  32'h3d16a564 /* (27, 23, 0) */,
  32'h3d3dc47d /* (23, 23, 0) */,
  32'h3d89a49e /* (19, 23, 0) */,
  32'h3d8df2c1 /* (15, 23, 0) */,
  32'h3d66dac1 /* (11, 23, 0) */,
  32'h3d23a039 /* (7, 23, 0) */,
  32'h3d1237a7 /* (3, 23, 0) */,
  32'h3d1d4601 /* (31, 19, 0) */,
  32'h3d384488 /* (27, 19, 0) */,
  32'h3d89a49e /* (23, 19, 0) */,
  32'h3de3e928 /* (19, 19, 0) */,
  32'h3df6cc6d /* (15, 19, 0) */,
  32'h3db3fd83 /* (11, 19, 0) */,
  32'h3d5a6fdd /* (7, 19, 0) */,
  32'h3d258110 /* (3, 19, 0) */,
  32'h3d155505 /* (31, 15, 0) */,
  32'h3d347f0a /* (27, 15, 0) */,
  32'h3d8df2c1 /* (23, 15, 0) */,
  32'h3df6cc6d /* (19, 15, 0) */,
  32'h3e086183 /* (15, 15, 0) */,
  32'h3dbe6d47 /* (11, 15, 0) */,
  32'h3d5b6048 /* (7, 15, 0) */,
  32'h3d1eeabe /* (3, 15, 0) */,
  32'h3d147e90 /* (31, 11, 0) */,
  32'h3d25e815 /* (27, 11, 0) */,
  32'h3d66dac1 /* (23, 11, 0) */,
  32'h3db3fd83 /* (19, 11, 0) */,
  32'h3dbe6d47 /* (15, 11, 0) */,
  32'h3d922642 /* (11, 11, 0) */,
  32'h3d3dcd22 /* (7, 11, 0) */,
  32'h3d198ce9 /* (3, 11, 0) */,
  32'h3d25463b /* (31, 7, 0) */,
  32'h3d154f7b /* (27, 7, 0) */,
  32'h3d23a039 /* (23, 7, 0) */,
  32'h3d5a6fdd /* (19, 7, 0) */,
  32'h3d5b6048 /* (15, 7, 0) */,
  32'h3d3dcd22 /* (11, 7, 0) */,
  32'h3d162f74 /* (7, 7, 0) */,
  32'h3d1cfd70 /* (3, 7, 0) */,
  32'h3dff9e3f /* (31, 3, 0) */,
  32'h3d490b0e /* (27, 3, 0) */,
  32'h3d1237a7 /* (23, 3, 0) */,
  32'h3d258110 /* (19, 3, 0) */,
  32'h3d1eeabe /* (15, 3, 0) */,
  32'h3d198ce9 /* (11, 3, 0) */,
  32'h3d1cfd70 /* (7, 3, 0) */,
  32'h3d9c797c /* (3, 3, 0) */,
  32'h3d8b1391 /* (30, 31, 28) */,
  32'h3d222a9c /* (26, 31, 28) */,
  32'h3d1839e3 /* (22, 31, 28) */,
  32'h3d303352 /* (18, 31, 28) */,
  32'h3d303352 /* (14, 31, 28) */,
  32'h3d1839e3 /* (10, 31, 28) */,
  32'h3d222a9c /* (6, 31, 28) */,
  32'h3d8b1391 /* (2, 31, 28) */,
  32'h3d2d8e0e /* (30, 27, 28) */,
  32'h3d153e19 /* (26, 27, 28) */,
  32'h3d28e3b2 /* (22, 27, 28) */,
  32'h3d53bb31 /* (18, 27, 28) */,
  32'h3d53bb31 /* (14, 27, 28) */,
  32'h3d28e3b2 /* (10, 27, 28) */,
  32'h3d153e19 /* (6, 27, 28) */,
  32'h3d2d8e0e /* (2, 27, 28) */,
  32'h3d14de35 /* (30, 23, 28) */,
  32'h3d2657dd /* (26, 23, 28) */,
  32'h3d68b7a2 /* (22, 23, 28) */,
  32'h3da4db8a /* (18, 23, 28) */,
  32'h3da4db8a /* (14, 23, 28) */,
  32'h3d68b7a2 /* (10, 23, 28) */,
  32'h3d2657dd /* (6, 23, 28) */,
  32'h3d14de35 /* (2, 23, 28) */,
  32'h3d3217f4 /* (30, 19, 28) */,
  32'h3d601ae9 /* (26, 19, 28) */,
  32'h3db40e50 /* (22, 19, 28) */,
  32'h3e0de89e /* (18, 19, 28) */,
  32'h3e0de89e /* (14, 19, 28) */,
  32'h3db40e50 /* (10, 19, 28) */,
  32'h3d601ae9 /* (6, 19, 28) */,
  32'h3d3217f4 /* (2, 19, 28) */,
  32'h3d2d6bba /* (30, 15, 28) */,
  32'h3d61b1de /* (26, 15, 28) */,
  32'h3dbdf4f8 /* (22, 15, 28) */,
  32'h3e1c2ca1 /* (18, 15, 28) */,
  32'h3e1c2ca1 /* (14, 15, 28) */,
  32'h3dbdf4f8 /* (10, 15, 28) */,
  32'h3d61b1de /* (6, 15, 28) */,
  32'h3d2d6bba /* (2, 15, 28) */,
  32'h3d21c128 /* (30, 11, 28) */,
  32'h3d41fb9f /* (26, 11, 28) */,
  32'h3d92b699 /* (22, 11, 28) */,
  32'h3ddc0819 /* (18, 11, 28) */,
  32'h3ddc0819 /* (14, 11, 28) */,
  32'h3d92b699 /* (10, 11, 28) */,
  32'h3d41fb9f /* (6, 11, 28) */,
  32'h3d21c128 /* (2, 11, 28) */,
  32'h3d16c6a3 /* (30, 7, 28) */,
  32'h3d17902e /* (26, 7, 28) */,
  32'h3d404057 /* (22, 7, 28) */,
  32'h3d800deb /* (18, 7, 28) */,
  32'h3d800deb /* (14, 7, 28) */,
  32'h3d404057 /* (10, 7, 28) */,
  32'h3d17902e /* (6, 7, 28) */,
  32'h3d16c6a3 /* (2, 7, 28) */,
  32'h3d5defd3 /* (30, 3, 28) */,
  32'h3d1b3fff /* (26, 3, 28) */,
  32'h3d1cff11 /* (22, 3, 28) */,
  32'h3d3b1e93 /* (18, 3, 28) */,
  32'h3d3b1e93 /* (14, 3, 28) */,
  32'h3d1cff11 /* (10, 3, 28) */,
  32'h3d1b3fff /* (6, 3, 28) */,
  32'h3d5defd3 /* (2, 3, 28) */,
  32'h3d15ce12 /* (30, 31, 24) */,
  32'h3d169650 /* (26, 31, 24) */,
  32'h3d3f0366 /* (22, 31, 24) */,
  32'h3d7e759f /* (18, 31, 24) */,
  32'h3d7e759f /* (14, 31, 24) */,
  32'h3d3f0366 /* (10, 31, 24) */,
  32'h3d169650 /* (6, 31, 24) */,
  32'h3d15ce12 /* (2, 31, 24) */,
  32'h3d149b5c /* (30, 27, 24) */,
  32'h3d22af34 /* (26, 27, 24) */,
  32'h3d5ef675 /* (22, 27, 24) */,
  32'h3d9bc970 /* (18, 27, 24) */,
  32'h3d9bc970 /* (14, 27, 24) */,
  32'h3d5ef675 /* (10, 27, 24) */,
  32'h3d22af34 /* (6, 27, 24) */,
  32'h3d149b5c /* (2, 27, 24) */,
  32'h3d3291f6 /* (30, 23, 24) */,
  32'h3d584c0c /* (26, 23, 24) */,
  32'h3da590e9 /* (22, 23, 24) */,
  32'h3dfaaa60 /* (18, 23, 24) */,
  32'h3dfaaa60 /* (14, 23, 24) */,
  32'h3da590e9 /* (10, 23, 24) */,
  32'h3d584c0c /* (6, 23, 24) */,
  32'h3d3291f6 /* (2, 23, 24) */,
  32'h3d7b52f8 /* (30, 19, 24) */,
  32'h3da2e7a9 /* (26, 19, 24) */,
  32'h3e085939 /* (22, 19, 24) */,
  32'h3e5f05ce /* (18, 19, 24) */,
  32'h3e5f05ce /* (14, 19, 24) */,
  32'h3e085939 /* (10, 19, 24) */,
  32'h3da2e7a9 /* (6, 19, 24) */,
  32'h3d7b52f8 /* (2, 19, 24) */,
  32'h3d804df8 /* (30, 15, 24) */,
  32'h3daa3349 /* (26, 15, 24) */,
  32'h3e135573 /* (22, 15, 24) */,
  32'h3e79034c /* (18, 15, 24) */,
  32'h3e79034c /* (14, 15, 24) */,
  32'h3e135573 /* (10, 15, 24) */,
  32'h3daa3349 /* (6, 15, 24) */,
  32'h3d804df8 /* (2, 15, 24) */,
  32'h3d558b1c /* (30, 11, 24) */,
  32'h3d865b59 /* (26, 11, 24) */,
  32'h3dd7e578 /* (22, 11, 24) */,
  32'h3e2a27e4 /* (18, 11, 24) */,
  32'h3e2a27e4 /* (14, 11, 24) */,
  32'h3dd7e578 /* (10, 11, 24) */,
  32'h3d865b59 /* (6, 11, 24) */,
  32'h3d558b1c /* (2, 11, 24) */,
  32'h3d1d59b0 /* (30, 7, 24) */,
  32'h3d35cd98 /* (26, 7, 24) */,
  32'h3d83c517 /* (22, 7, 24) */,
  32'h3dbf672f /* (18, 7, 24) */,
  32'h3dbf672f /* (14, 7, 24) */,
  32'h3d83c517 /* (10, 7, 24) */,
  32'h3d35cd98 /* (6, 7, 24) */,
  32'h3d1d59b0 /* (2, 7, 24) */,
  32'h3d13e9f7 /* (30, 3, 24) */,
  32'h3d19bf4b /* (26, 3, 24) */,
  32'h3d48bc7e /* (22, 3, 24) */,
  32'h3d880501 /* (18, 3, 24) */,
  32'h3d880501 /* (14, 3, 24) */,
  32'h3d48bc7e /* (10, 3, 24) */,
  32'h3d19bf4b /* (6, 3, 24) */,
  32'h3d13e9f7 /* (2, 3, 24) */,
  32'h3d1cac31 /* (30, 31, 20) */,
  32'h3d3dc5f0 /* (26, 31, 20) */,
  32'h3d91435f /* (22, 31, 20) */,
  32'h3ddbed5a /* (18, 31, 20) */,
  32'h3ddbed5a /* (14, 31, 20) */,
  32'h3d91435f /* (10, 31, 20) */,
  32'h3d3dc5f0 /* (6, 31, 20) */,
  32'h3d1cac31 /* (2, 31, 20) */,
  32'h3d346b02 /* (30, 27, 20) */,
  32'h3d6007ad /* (26, 27, 20) */,
  32'h3db0e528 /* (22, 27, 20) */,
  32'h3e095be4 /* (18, 27, 20) */,
  32'h3e095be4 /* (14, 27, 20) */,
  32'h3db0e528 /* (10, 27, 20) */,
  32'h3d6007ad /* (6, 27, 20) */,
  32'h3d346b02 /* (2, 27, 20) */,
  32'h3d833332 /* (30, 23, 20) */,
  32'h3da96159 /* (26, 23, 20) */,
  32'h3e0cf021 /* (22, 23, 20) */,
  32'h3e654448 /* (18, 23, 20) */,
  32'h3e654448 /* (14, 23, 20) */,
  32'h3e0cf021 /* (10, 23, 20) */,
  32'h3da96159 /* (6, 23, 20) */,
  32'h3d833332 /* (2, 23, 20) */,
  32'h3dd42d31 /* (30, 19, 20) */,
  32'h3e0dc95f /* (26, 19, 20) */,
  32'h3e7848b5 /* (22, 19, 20) */,
  32'h3ed441df /* (18, 19, 20) */,
  32'h3ed441df /* (14, 19, 20) */,
  32'h3e7848b5 /* (10, 19, 20) */,
  32'h3e0dc95f /* (6, 19, 20) */,
  32'h3dd42d31 /* (2, 19, 20) */,
  32'h3de39dff /* (30, 15, 20) */,
  32'h3e1a3a56 /* (26, 15, 20) */,
  32'h3e89fde5 /* (22, 15, 20) */,
  32'h3ef15f91 /* (18, 15, 20) */,
  32'h3ef15f91 /* (14, 15, 20) */,
  32'h3e89fde5 /* (10, 15, 20) */,
  32'h3e1a3a56 /* (6, 15, 20) */,
  32'h3de39dff /* (2, 15, 20) */,
  32'h3da96c08 /* (30, 11, 20) */,
  32'h3ddec971 /* (26, 11, 20) */,
  32'h3e3e5baf /* (22, 11, 20) */,
  32'h3e9ecc49 /* (18, 11, 20) */,
  32'h3e9ecc49 /* (14, 11, 20) */,
  32'h3e3e5baf /* (10, 11, 20) */,
  32'h3ddec971 /* (6, 11, 20) */,
  32'h3da96c08 /* (2, 11, 20) */,
  32'h3d530d8e /* (30, 7, 20) */,
  32'h3d859348 /* (26, 7, 20) */,
  32'h3dd85675 /* (22, 7, 20) */,
  32'h3e2baf50 /* (18, 7, 20) */,
  32'h3e2baf50 /* (14, 7, 20) */,
  32'h3dd85675 /* (10, 7, 20) */,
  32'h3d859348 /* (6, 7, 20) */,
  32'h3d530d8e /* (2, 7, 20) */,
  32'h3d23d587 /* (30, 3, 20) */,
  32'h3d48406d /* (26, 3, 20) */,
  32'h3d9aff71 /* (22, 3, 20) */,
  32'h3decc5e8 /* (18, 3, 20) */,
  32'h3decc5e8 /* (14, 3, 20) */,
  32'h3d9aff71 /* (10, 3, 20) */,
  32'h3d48406d /* (6, 3, 20) */,
  32'h3d23d587 /* (2, 3, 20) */,
  32'h3d09dfab /* (30, 31, 16) */,
  32'h3d34b66a /* (26, 31, 16) */,
  32'h3d99ac24 /* (22, 31, 16) */,
  32'h3dff32bb /* (18, 31, 16) */,
  32'h3dff32bb /* (14, 31, 16) */,
  32'h3d99ac24 /* (10, 31, 16) */,
  32'h3d34b66a /* (6, 31, 16) */,
  32'h3d09dfab /* (2, 31, 16) */,
  32'h3d28d1e5 /* (30, 27, 16) */,
  32'h3d5f53fb /* (26, 27, 16) */,
  32'h3dc0863e /* (22, 27, 16) */,
  32'h3e2205a1 /* (18, 27, 16) */,
  32'h3e2205a1 /* (14, 27, 16) */,
  32'h3dc0863e /* (10, 27, 16) */,
  32'h3d5f53fb /* (6, 27, 16) */,
  32'h3d28d1e5 /* (2, 27, 16) */,
  32'h3d87d16b /* (30, 23, 16) */,
  32'h3db6b309 /* (26, 23, 16) */,
  32'h3e21930d /* (22, 23, 16) */,
  32'h3e8b9344 /* (18, 23, 16) */,
  32'h3e8b9344 /* (14, 23, 16) */,
  32'h3e21930d /* (10, 23, 16) */,
  32'h3db6b309 /* (6, 23, 16) */,
  32'h3d87d16b /* (2, 23, 16) */,
  32'h3df1ae3d /* (30, 19, 16) */,
  32'h3e2576a9 /* (26, 19, 16) */,
  32'h3e968a40 /* (22, 19, 16) */,
  32'h3f06176f /* (18, 19, 16) */,
  32'h3f06176f /* (14, 19, 16) */,
  32'h3e968a40 /* (10, 19, 16) */,
  32'h3e2576a9 /* (6, 19, 16) */,
  32'h3df1ae3d /* (2, 19, 16) */,
  32'h3e06ec2e /* (30, 15, 16) */,
  32'h3e3a3d1a /* (26, 15, 16) */,
  32'h3eabb572 /* (22, 15, 16) */,
  32'h3f1b42bd /* (18, 15, 16) */,
  32'h3f1b42bd /* (14, 15, 16) */,
  32'h3eabb572 /* (10, 15, 16) */,
  32'h3e3a3d1a /* (6, 15, 16) */,
  32'h3e06ec2e /* (2, 15, 16) */,
  32'h3db86416 /* (30, 11, 16) */,
  32'h3dfa4afe /* (26, 11, 16) */,
  32'h3e60898b /* (22, 11, 16) */,
  32'h3ec4f0a1 /* (18, 11, 16) */,
  32'h3ec4f0a1 /* (14, 11, 16) */,
  32'h3e60898b /* (10, 11, 16) */,
  32'h3dfa4afe /* (6, 11, 16) */,
  32'h3db86416 /* (2, 11, 16) */,
  32'h3d4f6a6e /* (30, 7, 16) */,
  32'h3d8a46e7 /* (26, 7, 16) */,
  32'h3df142da /* (22, 7, 16) */,
  32'h3e4d7ce8 /* (18, 7, 16) */,
  32'h3e4d7ce8 /* (14, 7, 16) */,
  32'h3df142da /* (10, 7, 16) */,
  32'h3d8a46e7 /* (6, 7, 16) */,
  32'h3d4f6a6e /* (2, 7, 16) */,
  32'h3d13661d /* (30, 3, 16) */,
  32'h3d41d3ae /* (26, 3, 16) */,
  32'h3da59d10 /* (22, 3, 16) */,
  32'h3e0a27e7 /* (18, 3, 16) */,
  32'h3e0a27e7 /* (14, 3, 16) */,
  32'h3da59d10 /* (10, 3, 16) */,
  32'h3d41d3ae /* (6, 3, 16) */,
  32'h3d13661d /* (2, 3, 16) */,
  32'h3d1cac31 /* (30, 31, 12) */,
  32'h3d3dc5f0 /* (26, 31, 12) */,
  32'h3d91435f /* (22, 31, 12) */,
  32'h3ddbed5a /* (18, 31, 12) */,
  32'h3ddbed5a /* (14, 31, 12) */,
  32'h3d91435f /* (10, 31, 12) */,
  32'h3d3dc5f0 /* (6, 31, 12) */,
  32'h3d1cac31 /* (2, 31, 12) */,
  32'h3d346b02 /* (30, 27, 12) */,
  32'h3d6007ad /* (26, 27, 12) */,
  32'h3db0e528 /* (22, 27, 12) */,
  32'h3e095be4 /* (18, 27, 12) */,
  32'h3e095be4 /* (14, 27, 12) */,
  32'h3db0e528 /* (10, 27, 12) */,
  32'h3d6007ad /* (6, 27, 12) */,
  32'h3d346b02 /* (2, 27, 12) */,
  32'h3d833332 /* (30, 23, 12) */,
  32'h3da96159 /* (26, 23, 12) */,
  32'h3e0cf021 /* (22, 23, 12) */,
  32'h3e654448 /* (18, 23, 12) */,
  32'h3e654448 /* (14, 23, 12) */,
  32'h3e0cf021 /* (10, 23, 12) */,
  32'h3da96159 /* (6, 23, 12) */,
  32'h3d833332 /* (2, 23, 12) */,
  32'h3dd42d31 /* (30, 19, 12) */,
  32'h3e0dc95f /* (26, 19, 12) */,
  32'h3e7848b5 /* (22, 19, 12) */,
  32'h3ed441df /* (18, 19, 12) */,
  32'h3ed441df /* (14, 19, 12) */,
  32'h3e7848b5 /* (10, 19, 12) */,
  32'h3e0dc95f /* (6, 19, 12) */,
  32'h3dd42d31 /* (2, 19, 12) */,
  32'h3de39dff /* (30, 15, 12) */,
  32'h3e1a3a56 /* (26, 15, 12) */,
  32'h3e89fde5 /* (22, 15, 12) */,
  32'h3ef15f91 /* (18, 15, 12) */,
  32'h3ef15f91 /* (14, 15, 12) */,
  32'h3e89fde5 /* (10, 15, 12) */,
  32'h3e1a3a56 /* (6, 15, 12) */,
  32'h3de39dff /* (2, 15, 12) */,
  32'h3da96c08 /* (30, 11, 12) */,
  32'h3ddec971 /* (26, 11, 12) */,
  32'h3e3e5baf /* (22, 11, 12) */,
  32'h3e9ecc49 /* (18, 11, 12) */,
  32'h3e9ecc49 /* (14, 11, 12) */,
  32'h3e3e5baf /* (10, 11, 12) */,
  32'h3ddec971 /* (6, 11, 12) */,
  32'h3da96c08 /* (2, 11, 12) */,
  32'h3d530d8e /* (30, 7, 12) */,
  32'h3d859348 /* (26, 7, 12) */,
  32'h3dd85675 /* (22, 7, 12) */,
  32'h3e2baf50 /* (18, 7, 12) */,
  32'h3e2baf50 /* (14, 7, 12) */,
  32'h3dd85675 /* (10, 7, 12) */,
  32'h3d859348 /* (6, 7, 12) */,
  32'h3d530d8e /* (2, 7, 12) */,
  32'h3d23d587 /* (30, 3, 12) */,
  32'h3d48406d /* (26, 3, 12) */,
  32'h3d9aff71 /* (22, 3, 12) */,
  32'h3decc5e8 /* (18, 3, 12) */,
  32'h3decc5e8 /* (14, 3, 12) */,
  32'h3d9aff71 /* (10, 3, 12) */,
  32'h3d48406d /* (6, 3, 12) */,
  32'h3d23d587 /* (2, 3, 12) */,
  32'h3d15ce12 /* (30, 31, 8) */,
  32'h3d169650 /* (26, 31, 8) */,
  32'h3d3f0366 /* (22, 31, 8) */,
  32'h3d7e759f /* (18, 31, 8) */,
  32'h3d7e759f /* (14, 31, 8) */,
  32'h3d3f0366 /* (10, 31, 8) */,
  32'h3d169650 /* (6, 31, 8) */,
  32'h3d15ce12 /* (2, 31, 8) */,
  32'h3d149b5c /* (30, 27, 8) */,
  32'h3d22af34 /* (26, 27, 8) */,
  32'h3d5ef675 /* (22, 27, 8) */,
  32'h3d9bc970 /* (18, 27, 8) */,
  32'h3d9bc970 /* (14, 27, 8) */,
  32'h3d5ef675 /* (10, 27, 8) */,
  32'h3d22af34 /* (6, 27, 8) */,
  32'h3d149b5c /* (2, 27, 8) */,
  32'h3d3291f6 /* (30, 23, 8) */,
  32'h3d584c0c /* (26, 23, 8) */,
  32'h3da590e9 /* (22, 23, 8) */,
  32'h3dfaaa60 /* (18, 23, 8) */,
  32'h3dfaaa60 /* (14, 23, 8) */,
  32'h3da590e9 /* (10, 23, 8) */,
  32'h3d584c0c /* (6, 23, 8) */,
  32'h3d3291f6 /* (2, 23, 8) */,
  32'h3d7b52f8 /* (30, 19, 8) */,
  32'h3da2e7a9 /* (26, 19, 8) */,
  32'h3e085939 /* (22, 19, 8) */,
  32'h3e5f05ce /* (18, 19, 8) */,
  32'h3e5f05ce /* (14, 19, 8) */,
  32'h3e085939 /* (10, 19, 8) */,
  32'h3da2e7a9 /* (6, 19, 8) */,
  32'h3d7b52f8 /* (2, 19, 8) */,
  32'h3d804df8 /* (30, 15, 8) */,
  32'h3daa3349 /* (26, 15, 8) */,
  32'h3e135573 /* (22, 15, 8) */,
  32'h3e79034c /* (18, 15, 8) */,
  32'h3e79034c /* (14, 15, 8) */,
  32'h3e135573 /* (10, 15, 8) */,
  32'h3daa3349 /* (6, 15, 8) */,
  32'h3d804df8 /* (2, 15, 8) */,
  32'h3d558b1c /* (30, 11, 8) */,
  32'h3d865b59 /* (26, 11, 8) */,
  32'h3dd7e578 /* (22, 11, 8) */,
  32'h3e2a27e4 /* (18, 11, 8) */,
  32'h3e2a27e4 /* (14, 11, 8) */,
  32'h3dd7e578 /* (10, 11, 8) */,
  32'h3d865b59 /* (6, 11, 8) */,
  32'h3d558b1c /* (2, 11, 8) */,
  32'h3d1d59b0 /* (30, 7, 8) */,
  32'h3d35cd98 /* (26, 7, 8) */,
  32'h3d83c517 /* (22, 7, 8) */,
  32'h3dbf672f /* (18, 7, 8) */,
  32'h3dbf672f /* (14, 7, 8) */,
  32'h3d83c517 /* (10, 7, 8) */,
  32'h3d35cd98 /* (6, 7, 8) */,
  32'h3d1d59b0 /* (2, 7, 8) */,
  32'h3d13e9f7 /* (30, 3, 8) */,
  32'h3d19bf4b /* (26, 3, 8) */,
  32'h3d48bc7e /* (22, 3, 8) */,
  32'h3d880501 /* (18, 3, 8) */,
  32'h3d880501 /* (14, 3, 8) */,
  32'h3d48bc7e /* (10, 3, 8) */,
  32'h3d19bf4b /* (6, 3, 8) */,
  32'h3d13e9f7 /* (2, 3, 8) */,
  32'h3d8b1391 /* (30, 31, 4) */,
  32'h3d222a9c /* (26, 31, 4) */,
  32'h3d1839e3 /* (22, 31, 4) */,
  32'h3d303352 /* (18, 31, 4) */,
  32'h3d303352 /* (14, 31, 4) */,
  32'h3d1839e3 /* (10, 31, 4) */,
  32'h3d222a9c /* (6, 31, 4) */,
  32'h3d8b1391 /* (2, 31, 4) */,
  32'h3d2d8e0e /* (30, 27, 4) */,
  32'h3d153e19 /* (26, 27, 4) */,
  32'h3d28e3b2 /* (22, 27, 4) */,
  32'h3d53bb31 /* (18, 27, 4) */,
  32'h3d53bb31 /* (14, 27, 4) */,
  32'h3d28e3b2 /* (10, 27, 4) */,
  32'h3d153e19 /* (6, 27, 4) */,
  32'h3d2d8e0e /* (2, 27, 4) */,
  32'h3d14de35 /* (30, 23, 4) */,
  32'h3d2657dd /* (26, 23, 4) */,
  32'h3d68b7a2 /* (22, 23, 4) */,
  32'h3da4db8a /* (18, 23, 4) */,
  32'h3da4db8a /* (14, 23, 4) */,
  32'h3d68b7a2 /* (10, 23, 4) */,
  32'h3d2657dd /* (6, 23, 4) */,
  32'h3d14de35 /* (2, 23, 4) */,
  32'h3d3217f4 /* (30, 19, 4) */,
  32'h3d601ae9 /* (26, 19, 4) */,
  32'h3db40e50 /* (22, 19, 4) */,
  32'h3e0de89e /* (18, 19, 4) */,
  32'h3e0de89e /* (14, 19, 4) */,
  32'h3db40e50 /* (10, 19, 4) */,
  32'h3d601ae9 /* (6, 19, 4) */,
  32'h3d3217f4 /* (2, 19, 4) */,
  32'h3d2d6bba /* (30, 15, 4) */,
  32'h3d61b1de /* (26, 15, 4) */,
  32'h3dbdf4f8 /* (22, 15, 4) */,
  32'h3e1c2ca1 /* (18, 15, 4) */,
  32'h3e1c2ca1 /* (14, 15, 4) */,
  32'h3dbdf4f8 /* (10, 15, 4) */,
  32'h3d61b1de /* (6, 15, 4) */,
  32'h3d2d6bba /* (2, 15, 4) */,
  32'h3d21c128 /* (30, 11, 4) */,
  32'h3d41fb9f /* (26, 11, 4) */,
  32'h3d92b699 /* (22, 11, 4) */,
  32'h3ddc0819 /* (18, 11, 4) */,
  32'h3ddc0819 /* (14, 11, 4) */,
  32'h3d92b699 /* (10, 11, 4) */,
  32'h3d41fb9f /* (6, 11, 4) */,
  32'h3d21c128 /* (2, 11, 4) */,
  32'h3d16c6a3 /* (30, 7, 4) */,
  32'h3d17902e /* (26, 7, 4) */,
  32'h3d404057 /* (22, 7, 4) */,
  32'h3d800deb /* (18, 7, 4) */,
  32'h3d800deb /* (14, 7, 4) */,
  32'h3d404057 /* (10, 7, 4) */,
  32'h3d17902e /* (6, 7, 4) */,
  32'h3d16c6a3 /* (2, 7, 4) */,
  32'h3d5defd3 /* (30, 3, 4) */,
  32'h3d1b3fff /* (26, 3, 4) */,
  32'h3d1cff11 /* (22, 3, 4) */,
  32'h3d3b1e93 /* (18, 3, 4) */,
  32'h3d3b1e93 /* (14, 3, 4) */,
  32'h3d1cff11 /* (10, 3, 4) */,
  32'h3d1b3fff /* (6, 3, 4) */,
  32'h3d5defd3 /* (2, 3, 4) */,
  32'h3e709592 /* (30, 31, 0) */,
  32'h3d3f59b8 /* (26, 31, 0) */,
  32'h3d1142bb /* (22, 31, 0) */,
  32'h3d1ceee6 /* (18, 31, 0) */,
  32'h3d1ceee6 /* (14, 31, 0) */,
  32'h3d1142bb /* (10, 31, 0) */,
  32'h3d3f59b8 /* (6, 31, 0) */,
  32'h3e709592 /* (2, 31, 0) */,
  32'h3d5dd7d1 /* (30, 27, 0) */,
  32'h3d1b2f33 /* (26, 27, 0) */,
  32'h3d1cee15 /* (22, 27, 0) */,
  32'h3d3b0a55 /* (18, 27, 0) */,
  32'h3d3b0a55 /* (14, 27, 0) */,
  32'h3d1cee15 /* (10, 27, 0) */,
  32'h3d1b2f33 /* (6, 27, 0) */,
  32'h3d5dd7d1 /* (2, 27, 0) */,
  32'h3d11b684 /* (30, 23, 0) */,
  32'h3d1bc36a /* (26, 23, 0) */,
  32'h3d50a575 /* (22, 23, 0) */,
  32'h3d8fa52c /* (18, 23, 0) */,
  32'h3d8fa52c /* (14, 23, 0) */,
  32'h3d50a575 /* (10, 23, 0) */,
  32'h3d1bc36a /* (6, 23, 0) */,
  32'h3d11b684 /* (2, 23, 0) */,
  32'h3d2045b1 /* (30, 19, 0) */,
  32'h3d4703b2 /* (26, 19, 0) */,
  32'h3d9d248b /* (22, 19, 0) */,
  32'h3df40add /* (18, 19, 0) */,
  32'h3df40add /* (14, 19, 0) */,
  32'h3d9d248b /* (10, 19, 0) */,
  32'h3d4703b2 /* (6, 19, 0) */,
  32'h3d2045b1 /* (2, 19, 0) */,
  32'h3d18d610 /* (30, 15, 0) */,
  32'h3d455011 /* (26, 15, 0) */,
  32'h3da42e1b /* (22, 15, 0) */,
  32'h3e05899d /* (18, 15, 0) */,
  32'h3e05899d /* (14, 15, 0) */,
  32'h3da42e1b /* (10, 15, 0) */,
  32'h3d455011 /* (6, 15, 0) */,
  32'h3d18d610 /* (2, 15, 0) */,
  32'h3d164ce1 /* (30, 11, 0) */,
  32'h3d3013e2 /* (26, 11, 0) */,
  32'h3d819abc /* (22, 11, 0) */,
  32'h3dbe661f /* (18, 11, 0) */,
  32'h3dbe661f /* (14, 11, 0) */,
  32'h3d819abc /* (10, 11, 0) */,
  32'h3d3013e2 /* (6, 11, 0) */,
  32'h3d164ce1 /* (2, 11, 0) */,
  32'h3d21b235 /* (30, 7, 0) */,
  32'h3d1459dd /* (26, 7, 0) */,
  32'h3d2f5f5a /* (22, 7, 0) */,
  32'h3d60bf24 /* (18, 7, 0) */,
  32'h3d60bf24 /* (14, 7, 0) */,
  32'h3d2f5f5a /* (10, 7, 0) */,
  32'h3d1459dd /* (6, 7, 0) */,
  32'h3d21b235 /* (2, 7, 0) */,
  32'h3dcbea25 /* (30, 3, 0) */,
  32'h3d2d5b95 /* (26, 3, 0) */,
  32'h3d144f19 /* (22, 3, 0) */,
  32'h3d262b6e /* (18, 3, 0) */,
  32'h3d262b6e /* (14, 3, 0) */,
  32'h3d144f19 /* (10, 3, 0) */,
  32'h3d2d5b95 /* (6, 3, 0) */,
  32'h3dcbea25 /* (2, 3, 0) */,
  32'h3d6eb36b /* (29, 31, 28) */,
  32'h3d17ff6b /* (25, 31, 28) */,
  32'h3d1f5dc3 /* (21, 31, 28) */,
  32'h3d294c4b /* (17, 31, 28) */,
  32'h3d2e802a /* (13, 31, 28) */,
  32'h3d13f199 /* (9, 31, 28) */,
  32'h3d334ee4 /* (5, 31, 28) */,
  32'h3d9c757b /* (1, 31, 28) */,
  32'h3d25f5ce /* (29, 27, 28) */,
  32'h3d1508af /* (25, 27, 28) */,
  32'h3d358341 /* (21, 27, 28) */,
  32'h3d4def9b /* (17, 27, 28) */,
  32'h3d4ea6a0 /* (13, 27, 28) */,
  32'h3d1ee50b /* (9, 27, 28) */,
  32'h3d189061 /* (5, 27, 28) */,
  32'h3d334ee4 /* (1, 27, 28) */,
  32'h3d16b5b2 /* (29, 23, 28) */,
  32'h3d30de15 /* (25, 23, 28) */,
  32'h3d81d711 /* (21, 23, 28) */,
  32'h3da3c1ed /* (17, 23, 28) */,
  32'h3d9d0afa /* (13, 23, 28) */,
  32'h3d51a9d2 /* (9, 23, 28) */,
  32'h3d1ee50b /* (5, 23, 28) */,
  32'h3d13f199 /* (1, 23, 28) */,
  32'h3d385879 /* (29, 19, 28) */,
  32'h3d770afc /* (25, 19, 28) */,
  32'h3dcf13a3 /* (21, 19, 28) */,
  32'h3e0ff4ce /* (17, 19, 28) */,
  32'h3e0415cb /* (13, 19, 28) */,
  32'h3d9d0afa /* (9, 19, 28) */,
  32'h3d4ea6a0 /* (5, 19, 28) */,
  32'h3d2e802a /* (1, 19, 28) */,
  32'h3d349293 /* (29, 15, 28) */,
  32'h3d7b9f11 /* (25, 15, 28) */,
  32'h3ddcf428 /* (21, 15, 28) */,
  32'h3e1fe07e /* (17, 15, 28) */,
  32'h3e0ff4ce /* (13, 15, 28) */,
  32'h3da3c1ed /* (9, 15, 28) */,
  32'h3d4def9b /* (5, 15, 28) */,
  32'h3d294c4b /* (1, 15, 28) */,
  32'h3d25fa09 /* (29, 11, 28) */,
  32'h3d52976b /* (25, 11, 28) */,
  32'h3da66ad4 /* (21, 11, 28) */,
  32'h3ddcf428 /* (17, 11, 28) */,
  32'h3dcf13a3 /* (13, 11, 28) */,
  32'h3d81d711 /* (9, 11, 28) */,
  32'h3d358341 /* (5, 11, 28) */,
  32'h3d1f5dc3 /* (1, 11, 28) */,
  32'h3d155fa4 /* (29, 7, 28) */,
  32'h3d1cbb18 /* (25, 7, 28) */,
  32'h3d52976b /* (21, 7, 28) */,
  32'h3d7b9f11 /* (17, 7, 28) */,
  32'h3d770afc /* (13, 7, 28) */,
  32'h3d30de15 /* (9, 7, 28) */,
  32'h3d1508af /* (5, 7, 28) */,
  32'h3d17ff6b /* (1, 7, 28) */,
  32'h3d4920d0 /* (29, 3, 28) */,
  32'h3d155fa4 /* (25, 3, 28) */,
  32'h3d25fa09 /* (21, 3, 28) */,
  32'h3d349293 /* (17, 3, 28) */,
  32'h3d385879 /* (13, 3, 28) */,
  32'h3d16b5b2 /* (9, 3, 28) */,
  32'h3d25f5ce /* (5, 3, 28) */,
  32'h3d6eb36b /* (1, 3, 28) */,
  32'h3d146963 /* (29, 31, 24) */,
  32'h3d1bb8b6 /* (25, 31, 24) */,
  32'h3d513c3d /* (21, 31, 24) */,
  32'h3d7a003f /* (17, 31, 24) */,
  32'h3d7573b6 /* (13, 31, 24) */,
  32'h3d2fba80 /* (9, 31, 24) */,
  32'h3d1412fd /* (5, 31, 24) */,
  32'h3d1704d7 /* (1, 31, 24) */,
  32'h3d15d660 /* (29, 27, 24) */,
  32'h3d2bff3e /* (25, 27, 24) */,
  32'h3d77c8fd /* (21, 27, 24) */,
  32'h3d9a5b6b /* (17, 27, 24) */,
  32'h3d94d380 /* (13, 27, 24) */,
  32'h3d49c96c /* (9, 27, 24) */,
  32'h3d1c4d38 /* (5, 27, 24) */,
  32'h3d1412fd /* (1, 27, 24) */,
  32'h3d37919e /* (29, 23, 24) */,
  32'h3d6b8b35 /* (25, 23, 24) */,
  32'h3dbc4d73 /* (21, 23, 24) */,
  32'h3dfc30a3 /* (17, 23, 24) */,
  32'h3deb6b6d /* (13, 23, 24) */,
  32'h3d921bde /* (9, 23, 24) */,
  32'h3d49c96c /* (5, 23, 24) */,
  32'h3d2fba80 /* (1, 23, 24) */,
  32'h3d82c188 /* (29, 19, 24) */,
  32'h3db56072 /* (25, 19, 24) */,
  32'h3e1e607d /* (21, 19, 24) */,
  32'h3e640ba2 /* (17, 19, 24) */,
  32'h3e4dd3dc /* (13, 19, 24) */,
  32'h3deb6b6d /* (9, 19, 24) */,
  32'h3d94d380 /* (5, 19, 24) */,
  32'h3d7573b6 /* (1, 19, 24) */,
  32'h3d8608f0 /* (29, 15, 24) */,
  32'h3dbf0444 /* (25, 15, 24) */,
  32'h3e2c9c6c /* (21, 15, 24) */,
  32'h3e803f85 /* (17, 15, 24) */,
  32'h3e640ba2 /* (13, 15, 24) */,
  32'h3dfc30a3 /* (9, 15, 24) */,
  32'h3d9a5b6b /* (5, 15, 24) */,
  32'h3d7a003f /* (1, 15, 24) */,
  32'h3d5d0a38 /* (29, 11, 24) */,
  32'h3d941bce /* (25, 11, 24) */,
  32'h3df84bb3 /* (21, 11, 24) */,
  32'h3e2c9c6c /* (17, 11, 24) */,
  32'h3e1e607d /* (13, 11, 24) */,
  32'h3dbc4d73 /* (9, 11, 24) */,
  32'h3d77c8fd /* (5, 11, 24) */,
  32'h3d513c3d /* (1, 11, 24) */,
  32'h3d2054cd /* (29, 7, 24) */,
  32'h3d432bf1 /* (25, 7, 24) */,
  32'h3d941bce /* (21, 7, 24) */,
  32'h3dbf0444 /* (17, 7, 24) */,
  32'h3db56072 /* (13, 7, 24) */,
  32'h3d6b8b35 /* (9, 7, 24) */,
  32'h3d2bff3e /* (5, 7, 24) */,
  32'h3d1bb8b6 /* (1, 7, 24) */,
  32'h3d1392fe /* (29, 3, 24) */,
  32'h3d2054cd /* (25, 3, 24) */,
  32'h3d5d0a38 /* (21, 3, 24) */,
  32'h3d8608f0 /* (17, 3, 24) */,
  32'h3d82c188 /* (13, 3, 24) */,
  32'h3d37919e /* (9, 3, 24) */,
  32'h3d15d660 /* (5, 3, 24) */,
  32'h3d146963 /* (1, 3, 24) */,
  32'h3d210eee /* (29, 31, 20) */,
  32'h3d4ea8e5 /* (25, 31, 20) */,
  32'h3da53628 /* (21, 31, 20) */,
  32'h3ddd43c2 /* (17, 31, 20) */,
  32'h3dce8d02 /* (13, 31, 20) */,
  32'h3d803124 /* (9, 31, 20) */,
  32'h3d310ad3 /* (5, 31, 20) */,
  32'h3d1a2df1 /* (1, 31, 20) */,
  32'h3d3a4ebb /* (29, 27, 20) */,
  32'h3d75e4d4 /* (25, 27, 20) */,
  32'h3dca9d53 /* (21, 27, 20) */,
  32'h3e0ae903 /* (17, 27, 20) */,
  32'h3e00477d /* (13, 27, 20) */,
  32'h3d9af1c2 /* (9, 27, 20) */,
  32'h3d4f6dfc /* (5, 27, 20) */,
  32'h3d310ad3 /* (1, 27, 20) */,
  32'h3d886b82 /* (29, 23, 20) */,
  32'h3dbc51f9 /* (25, 23, 20) */,
  32'h3e23781b /* (21, 23, 20) */,
  32'h3e6a25fd /* (17, 23, 20) */,
  32'h3e53dc51 /* (13, 23, 20) */,
  32'h3df3b4f2 /* (9, 23, 20) */,
  32'h3d9af1c2 /* (5, 23, 20) */,
  32'h3d803124 /* (1, 23, 20) */,
  32'h3dddef48 /* (29, 19, 20) */,
  32'h3e1f8cbf /* (25, 19, 20) */,
  32'h3e91dfe2 /* (21, 19, 20) */,
  32'h3edb3822 /* (17, 19, 20) */,
  32'h3ec1d890 /* (13, 19, 20) */,
  32'h3e53dc51 /* (9, 19, 20) */,
  32'h3e00477d /* (5, 19, 20) */,
  32'h3dce8d02 /* (1, 19, 20) */,
  32'h3deea44d /* (29, 15, 20) */,
  32'h3e2e6a71 /* (25, 15, 20) */,
  32'h3ea31756 /* (21, 15, 20) */,
  32'h3efaa119 /* (17, 15, 20) */,
  32'h3edb3822 /* (13, 15, 20) */,
  32'h3e6a25fd /* (9, 15, 20) */,
  32'h3e0ae903 /* (5, 15, 20) */,
  32'h3ddd43c2 /* (1, 15, 20) */,
  32'h3db0b965 /* (29, 11, 20) */,
  32'h3df94537 /* (25, 11, 20) */,
  32'h3e5e44ac /* (21, 11, 20) */,
  32'h3ea31756 /* (17, 11, 20) */,
  32'h3e91dfe2 /* (13, 11, 20) */,
  32'h3e23781b /* (9, 11, 20) */,
  32'h3dca9d53 /* (5, 11, 20) */,
  32'h3da53628 /* (1, 11, 20) */,
  32'h3d5ab0e1 /* (29, 7, 20) */,
  32'h3d938890 /* (25, 7, 20) */,
  32'h3df94537 /* (21, 7, 20) */,
  32'h3e2e6a71 /* (17, 7, 20) */,
  32'h3e1f8cbf /* (13, 7, 20) */,
  32'h3dbc51f9 /* (9, 7, 20) */,
  32'h3d75e4d4 /* (5, 7, 20) */,
  32'h3d4ea8e5 /* (1, 7, 20) */,
  32'h3d28b308 /* (29, 3, 20) */,
  32'h3d5ab0e1 /* (25, 3, 20) */,
  32'h3db0b965 /* (21, 3, 20) */,
  32'h3deea44d /* (17, 3, 20) */,
  32'h3dddef48 /* (13, 3, 20) */,
  32'h3d886b82 /* (9, 3, 20) */,
  32'h3d3a4ebb /* (5, 3, 20) */,
  32'h3d210eee /* (1, 3, 20) */,
  32'h3d0fbc59 /* (29, 31, 16) */,
  32'h3d49f75a /* (25, 31, 16) */,
  32'h3db336e0 /* (21, 31, 16) */,
  32'h3e02e976 /* (17, 31, 16) */,
  32'h3deaafef /* (13, 31, 16) */,
  32'h3d8420c9 /* (9, 31, 16) */,
  32'h3d24852f /* (5, 31, 16) */,
  32'h3d067e68 /* (1, 31, 16) */,
  32'h3d3046d8 /* (29, 27, 16) */,
  32'h3d7a662c /* (25, 27, 16) */,
  32'h3de14ffa /* (21, 27, 16) */,
  32'h3e26bbbb /* (17, 27, 16) */,
  32'h3e1486b7 /* (13, 27, 16) */,
  32'h3da4f2f4 /* (9, 27, 16) */,
  32'h3d4ab7f7 /* (5, 27, 16) */,
  32'h3d24852f /* (1, 27, 16) */,
  32'h3d8e3848 /* (29, 23, 16) */,
  32'h3dce1075 /* (25, 23, 16) */,
  32'h3e3e5da7 /* (21, 23, 16) */,
  32'h3e908107 /* (17, 23, 16) */,
  32'h3e7e4b9d /* (13, 23, 16) */,
  32'h3e0981d7 /* (9, 23, 16) */,
  32'h3da4f2f4 /* (5, 23, 16) */,
  32'h3d8420c9 /* (1, 23, 16) */,
  32'h3dfdd31f /* (29, 19, 16) */,
  32'h3e3bd4ee /* (25, 19, 16) */,
  32'h3eb2bd2a /* (21, 19, 16) */,
  32'h3f0bd969 /* (17, 19, 16) */,
  32'h3ef27895 /* (13, 19, 16) */,
  32'h3e7e4b9d /* (9, 19, 16) */,
  32'h3e1486b7 /* (5, 19, 16) */,
  32'h3deaafef /* (1, 19, 16) */,
  32'h3e0de417 /* (29, 15, 16) */,
  32'h3e540b9b /* (25, 15, 16) */,
  32'h3ecca1ac /* (21, 15, 16) */,
  32'h3f2286f8 /* (17, 15, 16) */,
  32'h3f0bd969 /* (13, 15, 16) */,
  32'h3e908107 /* (9, 15, 16) */,
  32'h3e26bbbb /* (5, 15, 16) */,
  32'h3e02e976 /* (1, 15, 16) */,
  32'h3dc1602b /* (29, 11, 16) */,
  32'h3e0d9cf0 /* (25, 11, 16) */,
  32'h3e84c8e0 /* (21, 11, 16) */,
  32'h3ecca1ac /* (17, 11, 16) */,
  32'h3eb2bd2a /* (13, 11, 16) */,
  32'h3e3e5da7 /* (9, 11, 16) */,
  32'h3de14ffa /* (5, 11, 16) */,
  32'h3db336e0 /* (1, 11, 16) */,
  32'h3d58de26 /* (29, 7, 16) */,
  32'h3d9b7830 /* (25, 7, 16) */,
  32'h3e0d9cf0 /* (21, 7, 16) */,
  32'h3e540b9b /* (17, 7, 16) */,
  32'h3e3bd4ee /* (13, 7, 16) */,
  32'h3dce1075 /* (9, 7, 16) */,
  32'h3d7a662c /* (5, 7, 16) */,
  32'h3d49f75a /* (1, 7, 16) */,
  32'h3d19c07a /* (29, 3, 16) */,
  32'h3d58de26 /* (25, 3, 16) */,
  32'h3dc1602b /* (21, 3, 16) */,
  32'h3e0de417 /* (17, 3, 16) */,
  32'h3dfdd31f /* (13, 3, 16) */,
  32'h3d8e3848 /* (9, 3, 16) */,
  32'h3d3046d8 /* (5, 3, 16) */,
  32'h3d0fbc59 /* (1, 3, 16) */,
  32'h3d210eee /* (29, 31, 12) */,
  32'h3d4ea8e5 /* (25, 31, 12) */,
  32'h3da53628 /* (21, 31, 12) */,
  32'h3ddd43c2 /* (17, 31, 12) */,
  32'h3dce8d02 /* (13, 31, 12) */,
  32'h3d803124 /* (9, 31, 12) */,
  32'h3d310ad3 /* (5, 31, 12) */,
  32'h3d1a2df1 /* (1, 31, 12) */,
  32'h3d3a4ebb /* (29, 27, 12) */,
  32'h3d75e4d4 /* (25, 27, 12) */,
  32'h3dca9d53 /* (21, 27, 12) */,
  32'h3e0ae903 /* (17, 27, 12) */,
  32'h3e00477d /* (13, 27, 12) */,
  32'h3d9af1c2 /* (9, 27, 12) */,
  32'h3d4f6dfc /* (5, 27, 12) */,
  32'h3d310ad3 /* (1, 27, 12) */,
  32'h3d886b82 /* (29, 23, 12) */,
  32'h3dbc51f9 /* (25, 23, 12) */,
  32'h3e23781b /* (21, 23, 12) */,
  32'h3e6a25fd /* (17, 23, 12) */,
  32'h3e53dc51 /* (13, 23, 12) */,
  32'h3df3b4f2 /* (9, 23, 12) */,
  32'h3d9af1c2 /* (5, 23, 12) */,
  32'h3d803124 /* (1, 23, 12) */,
  32'h3dddef48 /* (29, 19, 12) */,
  32'h3e1f8cbf /* (25, 19, 12) */,
  32'h3e91dfe2 /* (21, 19, 12) */,
  32'h3edb3822 /* (17, 19, 12) */,
  32'h3ec1d890 /* (13, 19, 12) */,
  32'h3e53dc51 /* (9, 19, 12) */,
  32'h3e00477d /* (5, 19, 12) */,
  32'h3dce8d02 /* (1, 19, 12) */,
  32'h3deea44d /* (29, 15, 12) */,
  32'h3e2e6a71 /* (25, 15, 12) */,
  32'h3ea31756 /* (21, 15, 12) */,
  32'h3efaa119 /* (17, 15, 12) */,
  32'h3edb3822 /* (13, 15, 12) */,
  32'h3e6a25fd /* (9, 15, 12) */,
  32'h3e0ae903 /* (5, 15, 12) */,
  32'h3ddd43c2 /* (1, 15, 12) */,
  32'h3db0b965 /* (29, 11, 12) */,
  32'h3df94537 /* (25, 11, 12) */,
  32'h3e5e44ac /* (21, 11, 12) */,
  32'h3ea31756 /* (17, 11, 12) */,
  32'h3e91dfe2 /* (13, 11, 12) */,
  32'h3e23781b /* (9, 11, 12) */,
  32'h3dca9d53 /* (5, 11, 12) */,
  32'h3da53628 /* (1, 11, 12) */,
  32'h3d5ab0e1 /* (29, 7, 12) */,
  32'h3d938890 /* (25, 7, 12) */,
  32'h3df94537 /* (21, 7, 12) */,
  32'h3e2e6a71 /* (17, 7, 12) */,
  32'h3e1f8cbf /* (13, 7, 12) */,
  32'h3dbc51f9 /* (9, 7, 12) */,
  32'h3d75e4d4 /* (5, 7, 12) */,
  32'h3d4ea8e5 /* (1, 7, 12) */,
  32'h3d28b308 /* (29, 3, 12) */,
  32'h3d5ab0e1 /* (25, 3, 12) */,
  32'h3db0b965 /* (21, 3, 12) */,
  32'h3deea44d /* (17, 3, 12) */,
  32'h3dddef48 /* (13, 3, 12) */,
  32'h3d886b82 /* (9, 3, 12) */,
  32'h3d3a4ebb /* (5, 3, 12) */,
  32'h3d210eee /* (1, 3, 12) */,
  32'h3d146963 /* (29, 31, 8) */,
  32'h3d1bb8b6 /* (25, 31, 8) */,
  32'h3d513c3d /* (21, 31, 8) */,
  32'h3d7a003f /* (17, 31, 8) */,
  32'h3d7573b6 /* (13, 31, 8) */,
  32'h3d2fba80 /* (9, 31, 8) */,
  32'h3d1412fd /* (5, 31, 8) */,
  32'h3d1704d7 /* (1, 31, 8) */,
  32'h3d15d660 /* (29, 27, 8) */,
  32'h3d2bff3e /* (25, 27, 8) */,
  32'h3d77c8fd /* (21, 27, 8) */,
  32'h3d9a5b6b /* (17, 27, 8) */,
  32'h3d94d380 /* (13, 27, 8) */,
  32'h3d49c96c /* (9, 27, 8) */,
  32'h3d1c4d38 /* (5, 27, 8) */,
  32'h3d1412fd /* (1, 27, 8) */,
  32'h3d37919e /* (29, 23, 8) */,
  32'h3d6b8b35 /* (25, 23, 8) */,
  32'h3dbc4d73 /* (21, 23, 8) */,
  32'h3dfc30a3 /* (17, 23, 8) */,
  32'h3deb6b6d /* (13, 23, 8) */,
  32'h3d921bde /* (9, 23, 8) */,
  32'h3d49c96c /* (5, 23, 8) */,
  32'h3d2fba80 /* (1, 23, 8) */,
  32'h3d82c188 /* (29, 19, 8) */,
  32'h3db56072 /* (25, 19, 8) */,
  32'h3e1e607d /* (21, 19, 8) */,
  32'h3e640ba2 /* (17, 19, 8) */,
  32'h3e4dd3dc /* (13, 19, 8) */,
  32'h3deb6b6d /* (9, 19, 8) */,
  32'h3d94d380 /* (5, 19, 8) */,
  32'h3d7573b6 /* (1, 19, 8) */,
  32'h3d8608f0 /* (29, 15, 8) */,
  32'h3dbf0444 /* (25, 15, 8) */,
  32'h3e2c9c6c /* (21, 15, 8) */,
  32'h3e803f85 /* (17, 15, 8) */,
  32'h3e640ba2 /* (13, 15, 8) */,
  32'h3dfc30a3 /* (9, 15, 8) */,
  32'h3d9a5b6b /* (5, 15, 8) */,
  32'h3d7a003f /* (1, 15, 8) */,
  32'h3d5d0a38 /* (29, 11, 8) */,
  32'h3d941bce /* (25, 11, 8) */,
  32'h3df84bb3 /* (21, 11, 8) */,
  32'h3e2c9c6c /* (17, 11, 8) */,
  32'h3e1e607d /* (13, 11, 8) */,
  32'h3dbc4d73 /* (9, 11, 8) */,
  32'h3d77c8fd /* (5, 11, 8) */,
  32'h3d513c3d /* (1, 11, 8) */,
  32'h3d2054cd /* (29, 7, 8) */,
  32'h3d432bf1 /* (25, 7, 8) */,
  32'h3d941bce /* (21, 7, 8) */,
  32'h3dbf0444 /* (17, 7, 8) */,
  32'h3db56072 /* (13, 7, 8) */,
  32'h3d6b8b35 /* (9, 7, 8) */,
  32'h3d2bff3e /* (5, 7, 8) */,
  32'h3d1bb8b6 /* (1, 7, 8) */,
  32'h3d1392fe /* (29, 3, 8) */,
  32'h3d2054cd /* (25, 3, 8) */,
  32'h3d5d0a38 /* (21, 3, 8) */,
  32'h3d8608f0 /* (17, 3, 8) */,
  32'h3d82c188 /* (13, 3, 8) */,
  32'h3d37919e /* (9, 3, 8) */,
  32'h3d15d660 /* (5, 3, 8) */,
  32'h3d146963 /* (1, 3, 8) */,
  32'h3d6eb36b /* (29, 31, 4) */,
  32'h3d17ff6b /* (25, 31, 4) */,
  32'h3d1f5dc3 /* (21, 31, 4) */,
  32'h3d294c4b /* (17, 31, 4) */,
  32'h3d2e802a /* (13, 31, 4) */,
  32'h3d13f199 /* (9, 31, 4) */,
  32'h3d334ee4 /* (5, 31, 4) */,
  32'h3d9c757b /* (1, 31, 4) */,
  32'h3d25f5ce /* (29, 27, 4) */,
  32'h3d1508af /* (25, 27, 4) */,
  32'h3d358341 /* (21, 27, 4) */,
  32'h3d4def9b /* (17, 27, 4) */,
  32'h3d4ea6a0 /* (13, 27, 4) */,
  32'h3d1ee50b /* (9, 27, 4) */,
  32'h3d189061 /* (5, 27, 4) */,
  32'h3d334ee4 /* (1, 27, 4) */,
  32'h3d16b5b2 /* (29, 23, 4) */,
  32'h3d30de15 /* (25, 23, 4) */,
  32'h3d81d711 /* (21, 23, 4) */,
  32'h3da3c1ed /* (17, 23, 4) */,
  32'h3d9d0afa /* (13, 23, 4) */,
  32'h3d51a9d2 /* (9, 23, 4) */,
  32'h3d1ee50b /* (5, 23, 4) */,
  32'h3d13f199 /* (1, 23, 4) */,
  32'h3d385879 /* (29, 19, 4) */,
  32'h3d770afc /* (25, 19, 4) */,
  32'h3dcf13a3 /* (21, 19, 4) */,
  32'h3e0ff4ce /* (17, 19, 4) */,
  32'h3e0415cb /* (13, 19, 4) */,
  32'h3d9d0afa /* (9, 19, 4) */,
  32'h3d4ea6a0 /* (5, 19, 4) */,
  32'h3d2e802a /* (1, 19, 4) */,
  32'h3d349293 /* (29, 15, 4) */,
  32'h3d7b9f11 /* (25, 15, 4) */,
  32'h3ddcf428 /* (21, 15, 4) */,
  32'h3e1fe07e /* (17, 15, 4) */,
  32'h3e0ff4ce /* (13, 15, 4) */,
  32'h3da3c1ed /* (9, 15, 4) */,
  32'h3d4def9b /* (5, 15, 4) */,
  32'h3d294c4b /* (1, 15, 4) */,
  32'h3d25fa09 /* (29, 11, 4) */,
  32'h3d52976b /* (25, 11, 4) */,
  32'h3da66ad4 /* (21, 11, 4) */,
  32'h3ddcf428 /* (17, 11, 4) */,
  32'h3dcf13a3 /* (13, 11, 4) */,
  32'h3d81d711 /* (9, 11, 4) */,
  32'h3d358341 /* (5, 11, 4) */,
  32'h3d1f5dc3 /* (1, 11, 4) */,
  32'h3d155fa4 /* (29, 7, 4) */,
  32'h3d1cbb18 /* (25, 7, 4) */,
  32'h3d52976b /* (21, 7, 4) */,
  32'h3d7b9f11 /* (17, 7, 4) */,
  32'h3d770afc /* (13, 7, 4) */,
  32'h3d30de15 /* (9, 7, 4) */,
  32'h3d1508af /* (5, 7, 4) */,
  32'h3d17ff6b /* (1, 7, 4) */,
  32'h3d4920d0 /* (29, 3, 4) */,
  32'h3d155fa4 /* (25, 3, 4) */,
  32'h3d25fa09 /* (21, 3, 4) */,
  32'h3d349293 /* (17, 3, 4) */,
  32'h3d385879 /* (13, 3, 4) */,
  32'h3d16b5b2 /* (9, 3, 4) */,
  32'h3d25f5ce /* (5, 3, 4) */,
  32'h3d6eb36b /* (1, 3, 4) */,
  32'h3dff9e3f /* (29, 31, 0) */,
  32'h3d25463b /* (25, 31, 0) */,
  32'h3d147e90 /* (21, 31, 0) */,
  32'h3d155505 /* (17, 31, 0) */,
  32'h3d1d4601 /* (13, 31, 0) */,
  32'h3d11a5c6 /* (9, 31, 0) */,
  32'h3d6e9998 /* (5, 31, 0) */,
  32'h3f10fe39 /* (1, 31, 0) */,
  32'h3d490b0e /* (29, 27, 0) */,
  32'h3d154f7b /* (25, 27, 0) */,
  32'h3d25e815 /* (21, 27, 0) */,
  32'h3d347f0a /* (17, 27, 0) */,
  32'h3d384488 /* (13, 27, 0) */,
  32'h3d16a564 /* (9, 27, 0) */,
  32'h3d25e3da /* (5, 27, 0) */,
  32'h3d6e9998 /* (1, 27, 0) */,
  32'h3d1237a7 /* (29, 23, 0) */,
  32'h3d23a039 /* (25, 23, 0) */,
  32'h3d66dac1 /* (21, 23, 0) */,
  32'h3d8df2c1 /* (17, 23, 0) */,
  32'h3d89a49e /* (13, 23, 0) */,
  32'h3d3dc47d /* (9, 23, 0) */,
  32'h3d16a564 /* (5, 23, 0) */,
  32'h3d11a5c6 /* (1, 23, 0) */,
  32'h3d258110 /* (29, 19, 0) */,
  32'h3d5a6fdd /* (25, 19, 0) */,
  32'h3db3fd83 /* (21, 19, 0) */,
  32'h3df6cc6d /* (17, 19, 0) */,
  32'h3de3e928 /* (13, 19, 0) */,
  32'h3d89a49e /* (9, 19, 0) */,
  32'h3d384488 /* (5, 19, 0) */,
  32'h3d1d4601 /* (1, 19, 0) */,
  32'h3d1eeabe /* (29, 15, 0) */,
  32'h3d5b6048 /* (25, 15, 0) */,
  32'h3dbe6d47 /* (21, 15, 0) */,
  32'h3e086183 /* (17, 15, 0) */,
  32'h3df6cc6d /* (13, 15, 0) */,
  32'h3d8df2c1 /* (9, 15, 0) */,
  32'h3d347f0a /* (5, 15, 0) */,
  32'h3d155505 /* (1, 15, 0) */,
  32'h3d198ce9 /* (29, 11, 0) */,
  32'h3d3dcd22 /* (25, 11, 0) */,
  32'h3d922642 /* (21, 11, 0) */,
  32'h3dbe6d47 /* (17, 11, 0) */,
  32'h3db3fd83 /* (13, 11, 0) */,
  32'h3d66dac1 /* (9, 11, 0) */,
  32'h3d25e815 /* (5, 11, 0) */,
  32'h3d147e90 /* (1, 11, 0) */,
  32'h3d1cfd70 /* (29, 7, 0) */,
  32'h3d162f74 /* (25, 7, 0) */,
  32'h3d3dcd22 /* (21, 7, 0) */,
  32'h3d5b6048 /* (17, 7, 0) */,
  32'h3d5a6fdd /* (13, 7, 0) */,
  32'h3d23a039 /* (9, 7, 0) */,
  32'h3d154f7b /* (5, 7, 0) */,
  32'h3d25463b /* (1, 7, 0) */,
  32'h3d9c797c /* (29, 3, 0) */,
  32'h3d1cfd70 /* (25, 3, 0) */,
  32'h3d198ce9 /* (21, 3, 0) */,
  32'h3d1eeabe /* (17, 3, 0) */,
  32'h3d258110 /* (13, 3, 0) */,
  32'h3d1237a7 /* (9, 3, 0) */,
  32'h3d490b0e /* (5, 3, 0) */,
  32'h3dff9e3f /* (1, 3, 0) */,
  32'h3d4cb45d /* (28, 31, 28) */,
  32'h3d139499 /* (24, 31, 28) */,
  32'h3d27af27 /* (20, 31, 28) */,
  32'h3d18708b /* (16, 31, 28) */,
  32'h3d27af27 /* (12, 31, 28) */,
  32'h3d139499 /* (8, 31, 28) */,
  32'h3d4cb45d /* (4, 31, 28) */,
  32'h3da3aa58 /* (0, 31, 28) */,
  32'h3d1e7527 /* (28, 27, 28) */,
  32'h3d183845 /* (24, 27, 28) */,
  32'h3d431db1 /* (20, 27, 28) */,
  32'h3d3b5943 /* (16, 27, 28) */,
  32'h3d431db1 /* (12, 27, 28) */,
  32'h3d183845 /* (8, 27, 28) */,
  32'h3d1e7527 /* (4, 27, 28) */,
  32'h3d3577a5 /* (0, 27, 28) */,
  32'h3d19e157 /* (28, 23, 28) */,
  32'h3d3f1eea /* (24, 23, 28) */,
  32'h3d902ce0 /* (20, 23, 28) */,
  32'h3d97bb42 /* (16, 23, 28) */,
  32'h3d902ce0 /* (12, 23, 28) */,
  32'h3d3f1eea /* (8, 23, 28) */,
  32'h3d19e157 /* (4, 23, 28) */,
  32'h3d13aacb /* (0, 23, 28) */,
  32'h3d41aa67 /* (28, 19, 28) */,
  32'h3d8a5278 /* (24, 19, 28) */,
  32'h3dec6d9f /* (20, 19, 28) */,
  32'h3e07f264 /* (16, 19, 28) */,
  32'h3dec6d9f /* (12, 19, 28) */,
  32'h3d8a5278 /* (8, 19, 28) */,
  32'h3d41aa67 /* (4, 19, 28) */,
  32'h3d2d543a /* (0, 19, 28) */,
  32'h3d3f317e /* (28, 15, 28) */,
  32'h3d8e8b3a /* (24, 15, 28) */,
  32'h3dff07bf /* (20, 15, 28) */,
  32'h3e18449a /* (16, 15, 28) */,
  32'h3dff07bf /* (12, 15, 28) */,
  32'h3d8e8b3a /* (8, 15, 28) */,
  32'h3d3f317e /* (4, 15, 28) */,
  32'h3d27f384 /* (0, 15, 28) */,
  32'h3d2c64eb /* (28, 11, 28) */,
  32'h3d683712 /* (24, 11, 28) */,
  32'h3dbb90ec /* (20, 11, 28) */,
  32'h3dcebbc1 /* (16, 11, 28) */,
  32'h3dbb90ec /* (12, 11, 28) */,
  32'h3d683712 /* (8, 11, 28) */,
  32'h3d2c64eb /* (4, 11, 28) */,
  32'h3d1e982c /* (0, 11, 28) */,
  32'h3d148979 /* (28, 7, 28) */,
  32'h3d250b86 /* (24, 7, 28) */,
  32'h3d66108f /* (20, 7, 28) */,
  32'h3d66e7bc /* (16, 7, 28) */,
  32'h3d66108f /* (12, 7, 28) */,
  32'h3d250b86 /* (8, 7, 28) */,
  32'h3d148979 /* (4, 7, 28) */,
  32'h3d1879c9 /* (0, 7, 28) */,
  32'h3d358b49 /* (28, 3, 28) */,
  32'h3d13fed6 /* (24, 3, 28) */,
  32'h3d30047a /* (20, 3, 28) */,
  32'h3d232f37 /* (16, 3, 28) */,
  32'h3d30047a /* (12, 3, 28) */,
  32'h3d13fed6 /* (8, 3, 28) */,
  32'h3d358b49 /* (4, 3, 28) */,
  32'h3d7541a2 /* (0, 3, 28) */,
  32'h3d139499 /* (28, 31, 24) */,
  32'h3d23fb6f /* (24, 31, 24) */,
  32'h3d649547 /* (20, 31, 24) */,
  32'h3d656b11 /* (16, 31, 24) */,
  32'h3d649547 /* (12, 31, 24) */,
  32'h3d23fb6f /* (8, 31, 24) */,
  32'h3d139499 /* (4, 31, 24) */,
  32'h3d177e6a /* (0, 31, 24) */,
  32'h3d183845 /* (28, 27, 24) */,
  32'h3d38dbff /* (24, 27, 24) */,
  32'h3d89129f /* (20, 27, 24) */,
  32'h3d8eb3bf /* (16, 27, 24) */,
  32'h3d89129f /* (12, 27, 24) */,
  32'h3d38dbff /* (8, 27, 24) */,
  32'h3d183845 /* (4, 27, 24) */,
  32'h3d13eed3 /* (0, 27, 24) */,
  32'h3d3f1eea /* (28, 23, 24) */,
  32'h3d824402 /* (24, 23, 24) */,
  32'h3dd4c19e /* (20, 23, 24) */,
  32'h3dec5cc9 /* (16, 23, 24) */,
  32'h3dd4c19e /* (12, 23, 24) */,
  32'h3d824402 /* (8, 23, 24) */,
  32'h3d3f1eea /* (4, 23, 24) */,
  32'h3d2eceba /* (0, 23, 24) */,
  32'h3d8a5278 /* (28, 19, 24) */,
  32'h3dcd36cb /* (24, 19, 24) */,
  32'h3e368e5b /* (20, 19, 24) */,
  32'h3e58f4b1 /* (16, 19, 24) */,
  32'h3e368e5b /* (12, 19, 24) */,
  32'h3dcd36cb /* (8, 19, 24) */,
  32'h3d8a5278 /* (4, 19, 24) */,
  32'h3d7388b1 /* (0, 19, 24) */,
  32'h3d8e8b3a /* (28, 15, 24) */,
  32'h3dd9f1d0 /* (24, 15, 24) */,
  32'h3e48a298 /* (20, 15, 24) */,
  32'h3e75b861 /* (16, 15, 24) */,
  32'h3e48a298 /* (12, 15, 24) */,
  32'h3dd9f1d0 /* (8, 15, 24) */,
  32'h3d8e8b3a /* (4, 15, 24) */,
  32'h3d77d78b /* (0, 15, 24) */,
  32'h3d683712 /* (28, 11, 24) */,
  32'h3da5dafd /* (24, 11, 24) */,
  32'h3e0dbead /* (20, 11, 24) */,
  32'h3e2301df /* (16, 11, 24) */,
  32'h3e0dbead /* (12, 11, 24) */,
  32'h3da5dafd /* (8, 11, 24) */,
  32'h3d683712 /* (4, 11, 24) */,
  32'h3d4fd499 /* (0, 11, 24) */,
  32'h3d250b86 /* (28, 7, 24) */,
  32'h3d54dbd1 /* (24, 7, 24) */,
  32'h3da58a7f /* (20, 7, 24) */,
  32'h3db1ba44 /* (16, 7, 24) */,
  32'h3da58a7f /* (12, 7, 24) */,
  32'h3d54dbd1 /* (8, 7, 24) */,
  32'h3d250b86 /* (4, 7, 24) */,
  32'h3d1b34b2 /* (0, 7, 24) */,
  32'h3d13fed6 /* (28, 3, 24) */,
  32'h3d2a2238 /* (24, 3, 24) */,
  32'h3d729483 /* (20, 3, 24) */,
  32'h3d76a38f /* (16, 3, 24) */,
  32'h3d729483 /* (12, 3, 24) */,
  32'h3d2a2238 /* (8, 3, 24) */,
  32'h3d13fed6 /* (4, 3, 24) */,
  32'h3d14a194 /* (0, 3, 24) */,
  32'h3d27af27 /* (28, 31, 20) */,
  32'h3d649547 /* (24, 31, 20) */,
  32'h3dbaaaa9 /* (20, 31, 20) */,
  32'h3dcf60c6 /* (16, 31, 20) */,
  32'h3dbaaaa9 /* (12, 31, 20) */,
  32'h3d649547 /* (8, 31, 20) */,
  32'h3d27af27 /* (4, 31, 20) */,
  32'h3d195f14 /* (0, 31, 20) */,
  32'h3d431db1 /* (28, 27, 20) */,
  32'h3d89129f /* (24, 27, 20) */,
  32'h3de671da /* (20, 27, 20) */,
  32'h3e02cee2 /* (16, 27, 20) */,
  32'h3de671da /* (12, 27, 20) */,
  32'h3d89129f /* (8, 27, 20) */,
  32'h3d431db1 /* (4, 27, 20) */,
  32'h3d2ff16f /* (0, 27, 20) */,
  32'h3d902ce0 /* (28, 23, 20) */,
  32'h3dd4c19e /* (24, 23, 20) */,
  32'h3e3c290c /* (20, 23, 20) */,
  32'h3e5e82df /* (16, 23, 20) */,
  32'h3e3c290c /* (12, 23, 20) */,
  32'h3dd4c19e /* (8, 23, 20) */,
  32'h3d902ce0 /* (4, 23, 20) */,
  32'h3d7e6b4b /* (0, 23, 20) */,
  32'h3dec6d9f /* (28, 19, 20) */,
  32'h3e368e5b /* (24, 19, 20) */,
  32'h3eaa0eb2 /* (20, 19, 20) */,
  32'h3ed28b29 /* (16, 19, 20) */,
  32'h3eaa0eb2 /* (12, 19, 20) */,
  32'h3e368e5b /* (8, 19, 20) */,
  32'h3dec6d9f /* (4, 19, 20) */,
  32'h3dccb681 /* (0, 19, 20) */,
  32'h3dff07bf /* (28, 15, 20) */,
  32'h3e48a298 /* (24, 15, 20) */,
  32'h3ebf3a63 /* (20, 15, 20) */,
  32'h3ef1f40b /* (16, 15, 20) */,
  32'h3ebf3a63 /* (12, 15, 20) */,
  32'h3e48a298 /* (8, 15, 20) */,
  32'h3dff07bf /* (4, 15, 20) */,
  32'h3ddb309a /* (0, 15, 20) */,
  32'h3dbb90ec /* (28, 11, 20) */,
  32'h3e0dbead /* (24, 11, 20) */,
  32'h3e80c082 /* (20, 11, 20) */,
  32'h3e9bce24 /* (16, 11, 20) */,
  32'h3e80c082 /* (12, 11, 20) */,
  32'h3e0dbead /* (8, 11, 20) */,
  32'h3dbb90ec /* (4, 11, 20) */,
  32'h3da3d600 /* (0, 11, 20) */,
  32'h3d66108f /* (28, 7, 20) */,
  32'h3da58a7f /* (24, 7, 20) */,
  32'h3e0e8e1e /* (20, 7, 20) */,
  32'h3e24eefd /* (16, 7, 20) */,
  32'h3e0e8e1e /* (12, 7, 20) */,
  32'h3da58a7f /* (8, 7, 20) */,
  32'h3d66108f /* (4, 7, 20) */,
  32'h3d4d39f8 /* (0, 7, 20) */,
  32'h3d30047a /* (28, 3, 20) */,
  32'h3d729483 /* (24, 3, 20) */,
  32'h3dc823b1 /* (20, 3, 20) */,
  32'h3de007f6 /* (16, 3, 20) */,
  32'h3dc823b1 /* (12, 3, 20) */,
  32'h3d729483 /* (8, 3, 20) */,
  32'h3d30047a /* (4, 3, 20) */,
  32'h3d202826 /* (0, 3, 20) */,
  32'h3d18708b /* (28, 31, 16) */,
  32'h3d656b11 /* (24, 31, 16) */,
  32'h3dcf60c6 /* (20, 31, 16) */,
  32'h3df9e164 /* (16, 31, 16) */,
  32'h3dcf60c6 /* (12, 31, 16) */,
  32'h3d656b11 /* (8, 31, 16) */,
  32'h3d18708b /* (4, 31, 16) */,
  32'h3d0563b9 /* (0, 31, 16) */,
  32'h3d3b5943 /* (28, 27, 16) */,
  32'h3d8eb3bf /* (24, 27, 16) */,
  32'h3e02cee2 /* (20, 27, 16) */,
  32'h3e1f95bf /* (16, 27, 16) */,
  32'h3e02cee2 /* (12, 27, 16) */,
  32'h3d8eb3bf /* (8, 27, 16) */,
  32'h3d3b5943 /* (4, 27, 16) */,
  32'h3d231d8f /* (0, 27, 16) */,
  32'h3d97bb42 /* (28, 23, 16) */,
  32'h3dec5cc9 /* (24, 23, 16) */,
  32'h3e5e82df /* (20, 23, 16) */,
  32'h3e8b1bdf /* (16, 23, 16) */,
  32'h3e5e82df /* (12, 23, 16) */,
  32'h3dec5cc9 /* (8, 23, 16) */,
  32'h3d97bb42 /* (4, 23, 16) */,
  32'h3d82ec35 /* (0, 23, 16) */,
  32'h3e07f264 /* (28, 19, 16) */,
  32'h3e58f4b1 /* (24, 19, 16) */,
  32'h3ed28b29 /* (20, 19, 16) */,
  32'h3f079668 /* (16, 19, 16) */,
  32'h3ed28b29 /* (12, 19, 16) */,
  32'h3e58f4b1 /* (8, 19, 16) */,
  32'h3e07f264 /* (4, 19, 16) */,
  32'h3de8675d /* (0, 19, 16) */,
  32'h3e18449a /* (28, 15, 16) */,
  32'h3e75b861 /* (24, 15, 16) */,
  32'h3ef1f40b /* (20, 15, 16) */,
  32'h3f1e253a /* (16, 15, 16) */,
  32'h3ef1f40b /* (12, 15, 16) */,
  32'h3e75b861 /* (8, 15, 16) */,
  32'h3e18449a /* (4, 15, 16) */,
  32'h3e019a4f /* (0, 15, 16) */,
  32'h3dcebbc1 /* (28, 11, 16) */,
  32'h3e2301df /* (24, 11, 16) */,
  32'h3e9bce24 /* (20, 11, 16) */,
  32'h3ec5ad99 /* (16, 11, 16) */,
  32'h3e9bce24 /* (12, 11, 16) */,
  32'h3e2301df /* (8, 11, 16) */,
  32'h3dcebbc1 /* (4, 11, 16) */,
  32'h3db1860e /* (0, 11, 16) */,
  32'h3d66e7bc /* (28, 7, 16) */,
  32'h3db1ba44 /* (24, 7, 16) */,
  32'h3e24eefd /* (20, 7, 16) */,
  32'h3e4b7c7a /* (16, 7, 16) */,
  32'h3e24eefd /* (12, 7, 16) */,
  32'h3db1ba44 /* (8, 7, 16) */,
  32'h3d66e7bc /* (4, 7, 16) */,
  32'h3d482f92 /* (0, 7, 16) */,
  32'h3d232f37 /* (28, 3, 16) */,
  32'h3d76a38f /* (24, 3, 16) */,
  32'h3de007f6 /* (20, 3, 16) */,
  32'h3e078d5a /* (16, 3, 16) */,
  32'h3de007f6 /* (12, 3, 16) */,
  32'h3d76a38f /* (8, 3, 16) */,
  32'h3d232f37 /* (4, 3, 16) */,
  32'h3d0e89f8 /* (0, 3, 16) */,
  32'h3d27af27 /* (28, 31, 12) */,
  32'h3d649547 /* (24, 31, 12) */,
  32'h3dbaaaa9 /* (20, 31, 12) */,
  32'h3dcf60c6 /* (16, 31, 12) */,
  32'h3dbaaaa9 /* (12, 31, 12) */,
  32'h3d649547 /* (8, 31, 12) */,
  32'h3d27af27 /* (4, 31, 12) */,
  32'h3d195f14 /* (0, 31, 12) */,
  32'h3d431db1 /* (28, 27, 12) */,
  32'h3d89129f /* (24, 27, 12) */,
  32'h3de671da /* (20, 27, 12) */,
  32'h3e02cee2 /* (16, 27, 12) */,
  32'h3de671da /* (12, 27, 12) */,
  32'h3d89129f /* (8, 27, 12) */,
  32'h3d431db1 /* (4, 27, 12) */,
  32'h3d2ff16f /* (0, 27, 12) */,
  32'h3d902ce0 /* (28, 23, 12) */,
  32'h3dd4c19e /* (24, 23, 12) */,
  32'h3e3c290c /* (20, 23, 12) */,
  32'h3e5e82df /* (16, 23, 12) */,
  32'h3e3c290c /* (12, 23, 12) */,
  32'h3dd4c19e /* (8, 23, 12) */,
  32'h3d902ce0 /* (4, 23, 12) */,
  32'h3d7e6b4b /* (0, 23, 12) */,
  32'h3dec6d9f /* (28, 19, 12) */,
  32'h3e368e5b /* (24, 19, 12) */,
  32'h3eaa0eb2 /* (20, 19, 12) */,
  32'h3ed28b29 /* (16, 19, 12) */,
  32'h3eaa0eb2 /* (12, 19, 12) */,
  32'h3e368e5b /* (8, 19, 12) */,
  32'h3dec6d9f /* (4, 19, 12) */,
  32'h3dccb681 /* (0, 19, 12) */,
  32'h3dff07bf /* (28, 15, 12) */,
  32'h3e48a298 /* (24, 15, 12) */,
  32'h3ebf3a63 /* (20, 15, 12) */,
  32'h3ef1f40b /* (16, 15, 12) */,
  32'h3ebf3a63 /* (12, 15, 12) */,
  32'h3e48a298 /* (8, 15, 12) */,
  32'h3dff07bf /* (4, 15, 12) */,
  32'h3ddb309a /* (0, 15, 12) */,
  32'h3dbb90ec /* (28, 11, 12) */,
  32'h3e0dbead /* (24, 11, 12) */,
  32'h3e80c082 /* (20, 11, 12) */,
  32'h3e9bce24 /* (16, 11, 12) */,
  32'h3e80c082 /* (12, 11, 12) */,
  32'h3e0dbead /* (8, 11, 12) */,
  32'h3dbb90ec /* (4, 11, 12) */,
  32'h3da3d600 /* (0, 11, 12) */,
  32'h3d66108f /* (28, 7, 12) */,
  32'h3da58a7f /* (24, 7, 12) */,
  32'h3e0e8e1e /* (20, 7, 12) */,
  32'h3e24eefd /* (16, 7, 12) */,
  32'h3e0e8e1e /* (12, 7, 12) */,
  32'h3da58a7f /* (8, 7, 12) */,
  32'h3d66108f /* (4, 7, 12) */,
  32'h3d4d39f8 /* (0, 7, 12) */,
  32'h3d30047a /* (28, 3, 12) */,
  32'h3d729483 /* (24, 3, 12) */,
  32'h3dc823b1 /* (20, 3, 12) */,
  32'h3de007f6 /* (16, 3, 12) */,
  32'h3dc823b1 /* (12, 3, 12) */,
  32'h3d729483 /* (8, 3, 12) */,
  32'h3d30047a /* (4, 3, 12) */,
  32'h3d202826 /* (0, 3, 12) */,
  32'h3d139499 /* (28, 31, 8) */,
  32'h3d23fb6f /* (24, 31, 8) */,
  32'h3d649547 /* (20, 31, 8) */,
  32'h3d656b11 /* (16, 31, 8) */,
  32'h3d649547 /* (12, 31, 8) */,
  32'h3d23fb6f /* (8, 31, 8) */,
  32'h3d139499 /* (4, 31, 8) */,
  32'h3d177e6a /* (0, 31, 8) */,
  32'h3d183845 /* (28, 27, 8) */,
  32'h3d38dbff /* (24, 27, 8) */,
  32'h3d89129f /* (20, 27, 8) */,
  32'h3d8eb3bf /* (16, 27, 8) */,
  32'h3d89129f /* (12, 27, 8) */,
  32'h3d38dbff /* (8, 27, 8) */,
  32'h3d183845 /* (4, 27, 8) */,
  32'h3d13eed3 /* (0, 27, 8) */,
  32'h3d3f1eea /* (28, 23, 8) */,
  32'h3d824402 /* (24, 23, 8) */,
  32'h3dd4c19e /* (20, 23, 8) */,
  32'h3dec5cc9 /* (16, 23, 8) */,
  32'h3dd4c19e /* (12, 23, 8) */,
  32'h3d824402 /* (8, 23, 8) */,
  32'h3d3f1eea /* (4, 23, 8) */,
  32'h3d2eceba /* (0, 23, 8) */,
  32'h3d8a5278 /* (28, 19, 8) */,
  32'h3dcd36cb /* (24, 19, 8) */,
  32'h3e368e5b /* (20, 19, 8) */,
  32'h3e58f4b1 /* (16, 19, 8) */,
  32'h3e368e5b /* (12, 19, 8) */,
  32'h3dcd36cb /* (8, 19, 8) */,
  32'h3d8a5278 /* (4, 19, 8) */,
  32'h3d7388b1 /* (0, 19, 8) */,
  32'h3d8e8b3a /* (28, 15, 8) */,
  32'h3dd9f1d0 /* (24, 15, 8) */,
  32'h3e48a298 /* (20, 15, 8) */,
  32'h3e75b861 /* (16, 15, 8) */,
  32'h3e48a298 /* (12, 15, 8) */,
  32'h3dd9f1d0 /* (8, 15, 8) */,
  32'h3d8e8b3a /* (4, 15, 8) */,
  32'h3d77d78b /* (0, 15, 8) */,
  32'h3d683712 /* (28, 11, 8) */,
  32'h3da5dafd /* (24, 11, 8) */,
  32'h3e0dbead /* (20, 11, 8) */,
  32'h3e2301df /* (16, 11, 8) */,
  32'h3e0dbead /* (12, 11, 8) */,
  32'h3da5dafd /* (8, 11, 8) */,
  32'h3d683712 /* (4, 11, 8) */,
  32'h3d4fd499 /* (0, 11, 8) */,
  32'h3d250b86 /* (28, 7, 8) */,
  32'h3d54dbd1 /* (24, 7, 8) */,
  32'h3da58a7f /* (20, 7, 8) */,
  32'h3db1ba44 /* (16, 7, 8) */,
  32'h3da58a7f /* (12, 7, 8) */,
  32'h3d54dbd1 /* (8, 7, 8) */,
  32'h3d250b86 /* (4, 7, 8) */,
  32'h3d1b34b2 /* (0, 7, 8) */,
  32'h3d13fed6 /* (28, 3, 8) */,
  32'h3d2a2238 /* (24, 3, 8) */,
  32'h3d729483 /* (20, 3, 8) */,
  32'h3d76a38f /* (16, 3, 8) */,
  32'h3d729483 /* (12, 3, 8) */,
  32'h3d2a2238 /* (8, 3, 8) */,
  32'h3d13fed6 /* (4, 3, 8) */,
  32'h3d14a194 /* (0, 3, 8) */,
  32'h3d4cb45d /* (28, 31, 4) */,
  32'h3d139499 /* (24, 31, 4) */,
  32'h3d27af27 /* (20, 31, 4) */,
  32'h3d18708b /* (16, 31, 4) */,
  32'h3d27af27 /* (12, 31, 4) */,
  32'h3d139499 /* (8, 31, 4) */,
  32'h3d4cb45d /* (4, 31, 4) */,
  32'h3da3aa58 /* (0, 31, 4) */,
  32'h3d1e7527 /* (28, 27, 4) */,
  32'h3d183845 /* (24, 27, 4) */,
  32'h3d431db1 /* (20, 27, 4) */,
  32'h3d3b5943 /* (16, 27, 4) */,
  32'h3d431db1 /* (12, 27, 4) */,
  32'h3d183845 /* (8, 27, 4) */,
  32'h3d1e7527 /* (4, 27, 4) */,
  32'h3d3577a5 /* (0, 27, 4) */,
  32'h3d19e157 /* (28, 23, 4) */,
  32'h3d3f1eea /* (24, 23, 4) */,
  32'h3d902ce0 /* (20, 23, 4) */,
  32'h3d97bb42 /* (16, 23, 4) */,
  32'h3d902ce0 /* (12, 23, 4) */,
  32'h3d3f1eea /* (8, 23, 4) */,
  32'h3d19e157 /* (4, 23, 4) */,
  32'h3d13aacb /* (0, 23, 4) */,
  32'h3d41aa67 /* (28, 19, 4) */,
  32'h3d8a5278 /* (24, 19, 4) */,
  32'h3dec6d9f /* (20, 19, 4) */,
  32'h3e07f264 /* (16, 19, 4) */,
  32'h3dec6d9f /* (12, 19, 4) */,
  32'h3d8a5278 /* (8, 19, 4) */,
  32'h3d41aa67 /* (4, 19, 4) */,
  32'h3d2d543a /* (0, 19, 4) */,
  32'h3d3f317e /* (28, 15, 4) */,
  32'h3d8e8b3a /* (24, 15, 4) */,
  32'h3dff07bf /* (20, 15, 4) */,
  32'h3e18449a /* (16, 15, 4) */,
  32'h3dff07bf /* (12, 15, 4) */,
  32'h3d8e8b3a /* (8, 15, 4) */,
  32'h3d3f317e /* (4, 15, 4) */,
  32'h3d27f384 /* (0, 15, 4) */,
  32'h3d2c64eb /* (28, 11, 4) */,
  32'h3d683712 /* (24, 11, 4) */,
  32'h3dbb90ec /* (20, 11, 4) */,
  32'h3dcebbc1 /* (16, 11, 4) */,
  32'h3dbb90ec /* (12, 11, 4) */,
  32'h3d683712 /* (8, 11, 4) */,
  32'h3d2c64eb /* (4, 11, 4) */,
  32'h3d1e982c /* (0, 11, 4) */,
  32'h3d148979 /* (28, 7, 4) */,
  32'h3d250b86 /* (24, 7, 4) */,
  32'h3d66108f /* (20, 7, 4) */,
  32'h3d66e7bc /* (16, 7, 4) */,
  32'h3d66108f /* (12, 7, 4) */,
  32'h3d250b86 /* (8, 7, 4) */,
  32'h3d148979 /* (4, 7, 4) */,
  32'h3d1879c9 /* (0, 7, 4) */,
  32'h3d358b49 /* (28, 3, 4) */,
  32'h3d13fed6 /* (24, 3, 4) */,
  32'h3d30047a /* (20, 3, 4) */,
  32'h3d232f37 /* (16, 3, 4) */,
  32'h3d30047a /* (12, 3, 4) */,
  32'h3d13fed6 /* (8, 3, 4) */,
  32'h3d358b49 /* (4, 3, 4) */,
  32'h3d7541a2 /* (0, 3, 4) */,
  32'h3da3aa58 /* (28, 31, 0) */,
  32'h3d177e6a /* (24, 31, 0) */,
  32'h3d195f14 /* (20, 31, 0) */,
  32'h3d0563b9 /* (16, 31, 0) */,
  32'h3d195f14 /* (12, 31, 0) */,
  32'h3d177e6a /* (8, 31, 0) */,
  32'h3da3aa58 /* (4, 31, 0) */,
  32'h3f8f3ec8 /* (0, 31, 0) */,
  32'h3d3577a5 /* (28, 27, 0) */,
  32'h3d13eed3 /* (24, 27, 0) */,
  32'h3d2ff16f /* (20, 27, 0) */,
  32'h3d231d8f /* (16, 27, 0) */,
  32'h3d2ff16f /* (12, 27, 0) */,
  32'h3d13eed3 /* (8, 27, 0) */,
  32'h3d3577a5 /* (4, 27, 0) */,
  32'h3d75271a /* (0, 27, 0) */,
  32'h3d13aacb /* (28, 23, 0) */,
  32'h3d2eceba /* (24, 23, 0) */,
  32'h3d7e6b4b /* (20, 23, 0) */,
  32'h3d82ec35 /* (16, 23, 0) */,
  32'h3d7e6b4b /* (12, 23, 0) */,
  32'h3d2eceba /* (8, 23, 0) */,
  32'h3d13aacb /* (4, 23, 0) */,
  32'h3d11ab15 /* (0, 23, 0) */,
  32'h3d2d543a /* (28, 19, 0) */,
  32'h3d7388b1 /* (24, 19, 0) */,
  32'h3dccb681 /* (20, 19, 0) */,
  32'h3de8675d /* (16, 19, 0) */,
  32'h3dccb681 /* (12, 19, 0) */,
  32'h3d7388b1 /* (8, 19, 0) */,
  32'h3d2d543a /* (4, 19, 0) */,
  32'h3d1c4c09 /* (0, 19, 0) */,
  32'h3d27f384 /* (28, 15, 0) */,
  32'h3d77d78b /* (24, 15, 0) */,
  32'h3ddb309a /* (20, 15, 0) */,
  32'h3e019a4f /* (16, 15, 0) */,
  32'h3ddb309a /* (12, 15, 0) */,
  32'h3d77d78b /* (8, 15, 0) */,
  32'h3d27f384 /* (4, 15, 0) */,
  32'h3d14300c /* (0, 15, 0) */,
  32'h3d1e982c /* (28, 11, 0) */,
  32'h3d4fd499 /* (24, 11, 0) */,
  32'h3da3d600 /* (20, 11, 0) */,
  32'h3db1860e /* (16, 11, 0) */,
  32'h3da3d600 /* (12, 11, 0) */,
  32'h3d4fd499 /* (8, 11, 0) */,
  32'h3d1e982c /* (4, 11, 0) */,
  32'h3d13eab3 /* (0, 11, 0) */,
  32'h3d1879c9 /* (28, 7, 0) */,
  32'h3d1b34b2 /* (24, 7, 0) */,
  32'h3d4d39f8 /* (20, 7, 0) */,
  32'h3d482f92 /* (16, 7, 0) */,
  32'h3d4d39f8 /* (12, 7, 0) */,
  32'h3d1b34b2 /* (8, 7, 0) */,
  32'h3d1879c9 /* (4, 7, 0) */,
  32'h3d269d45 /* (0, 7, 0) */,
  32'h3d7541a2 /* (28, 3, 0) */,
  32'h3d14a194 /* (24, 3, 0) */,
  32'h3d202826 /* (20, 3, 0) */,
  32'h3d0e89f8 /* (16, 3, 0) */,
  32'h3d202826 /* (12, 3, 0) */,
  32'h3d14a194 /* (8, 3, 0) */,
  32'h3d7541a2 /* (4, 3, 0) */,
  32'h3e0c4c59 /* (0, 3, 0) */,
  32'h3d8b1391 /* (31, 30, 28) */,
  32'h3d2d8e0e /* (27, 30, 28) */,
  32'h3d14de35 /* (23, 30, 28) */,
  32'h3d3217f4 /* (19, 30, 28) */,
  32'h3d2d6bba /* (15, 30, 28) */,
  32'h3d21c128 /* (11, 30, 28) */,
  32'h3d16c6a3 /* (7, 30, 28) */,
  32'h3d5defd3 /* (3, 30, 28) */,
  32'h3d222a9c /* (31, 26, 28) */,
  32'h3d153e19 /* (27, 26, 28) */,
  32'h3d2657dd /* (23, 26, 28) */,
  32'h3d601ae9 /* (19, 26, 28) */,
  32'h3d61b1de /* (15, 26, 28) */,
  32'h3d41fb9f /* (11, 26, 28) */,
  32'h3d17902e /* (7, 26, 28) */,
  32'h3d1b3fff /* (3, 26, 28) */,
  32'h3d1839e3 /* (31, 22, 28) */,
  32'h3d28e3b2 /* (27, 22, 28) */,
  32'h3d68b7a2 /* (23, 22, 28) */,
  32'h3db40e50 /* (19, 22, 28) */,
  32'h3dbdf4f8 /* (15, 22, 28) */,
  32'h3d92b699 /* (11, 22, 28) */,
  32'h3d404057 /* (7, 22, 28) */,
  32'h3d1cff11 /* (3, 22, 28) */,
  32'h3d303352 /* (31, 18, 28) */,
  32'h3d53bb31 /* (27, 18, 28) */,
  32'h3da4db8a /* (23, 18, 28) */,
  32'h3e0de89e /* (19, 18, 28) */,
  32'h3e1c2ca1 /* (15, 18, 28) */,
  32'h3ddc0819 /* (11, 18, 28) */,
  32'h3d800deb /* (7, 18, 28) */,
  32'h3d3b1e93 /* (3, 18, 28) */,
  32'h3d303352 /* (31, 14, 28) */,
  32'h3d53bb31 /* (27, 14, 28) */,
  32'h3da4db8a /* (23, 14, 28) */,
  32'h3e0de89e /* (19, 14, 28) */,
  32'h3e1c2ca1 /* (15, 14, 28) */,
  32'h3ddc0819 /* (11, 14, 28) */,
  32'h3d800deb /* (7, 14, 28) */,
  32'h3d3b1e93 /* (3, 14, 28) */,
  32'h3d1839e3 /* (31, 10, 28) */,
  32'h3d28e3b2 /* (27, 10, 28) */,
  32'h3d68b7a2 /* (23, 10, 28) */,
  32'h3db40e50 /* (19, 10, 28) */,
  32'h3dbdf4f8 /* (15, 10, 28) */,
  32'h3d92b699 /* (11, 10, 28) */,
  32'h3d404057 /* (7, 10, 28) */,
  32'h3d1cff11 /* (3, 10, 28) */,
  32'h3d222a9c /* (31, 6, 28) */,
  32'h3d153e19 /* (27, 6, 28) */,
  32'h3d2657dd /* (23, 6, 28) */,
  32'h3d601ae9 /* (19, 6, 28) */,
  32'h3d61b1de /* (15, 6, 28) */,
  32'h3d41fb9f /* (11, 6, 28) */,
  32'h3d17902e /* (7, 6, 28) */,
  32'h3d1b3fff /* (3, 6, 28) */,
  32'h3d8b1391 /* (31, 2, 28) */,
  32'h3d2d8e0e /* (27, 2, 28) */,
  32'h3d14de35 /* (23, 2, 28) */,
  32'h3d3217f4 /* (19, 2, 28) */,
  32'h3d2d6bba /* (15, 2, 28) */,
  32'h3d21c128 /* (11, 2, 28) */,
  32'h3d16c6a3 /* (7, 2, 28) */,
  32'h3d5defd3 /* (3, 2, 28) */,
  32'h3d15ce12 /* (31, 30, 24) */,
  32'h3d149b5c /* (27, 30, 24) */,
  32'h3d3291f6 /* (23, 30, 24) */,
  32'h3d7b52f8 /* (19, 30, 24) */,
  32'h3d804df8 /* (15, 30, 24) */,
  32'h3d558b1c /* (11, 30, 24) */,
  32'h3d1d59b0 /* (7, 30, 24) */,
  32'h3d13e9f7 /* (3, 30, 24) */,
  32'h3d169650 /* (31, 26, 24) */,
  32'h3d22af34 /* (27, 26, 24) */,
  32'h3d584c0c /* (23, 26, 24) */,
  32'h3da2e7a9 /* (19, 26, 24) */,
  32'h3daa3349 /* (15, 26, 24) */,
  32'h3d865b59 /* (11, 26, 24) */,
  32'h3d35cd98 /* (7, 26, 24) */,
  32'h3d19bf4b /* (3, 26, 24) */,
  32'h3d3f0366 /* (31, 22, 24) */,
  32'h3d5ef675 /* (27, 22, 24) */,
  32'h3da590e9 /* (23, 22, 24) */,
  32'h3e085939 /* (19, 22, 24) */,
  32'h3e135573 /* (15, 22, 24) */,
  32'h3dd7e578 /* (11, 22, 24) */,
  32'h3d83c517 /* (7, 22, 24) */,
  32'h3d48bc7e /* (3, 22, 24) */,
  32'h3d7e759f /* (31, 18, 24) */,
  32'h3d9bc970 /* (27, 18, 24) */,
  32'h3dfaaa60 /* (23, 18, 24) */,
  32'h3e5f05ce /* (19, 18, 24) */,
  32'h3e79034c /* (15, 18, 24) */,
  32'h3e2a27e4 /* (11, 18, 24) */,
  32'h3dbf672f /* (7, 18, 24) */,
  32'h3d880501 /* (3, 18, 24) */,
  32'h3d7e759f /* (31, 14, 24) */,
  32'h3d9bc970 /* (27, 14, 24) */,
  32'h3dfaaa60 /* (23, 14, 24) */,
  32'h3e5f05ce /* (19, 14, 24) */,
  32'h3e79034c /* (15, 14, 24) */,
  32'h3e2a27e4 /* (11, 14, 24) */,
  32'h3dbf672f /* (7, 14, 24) */,
  32'h3d880501 /* (3, 14, 24) */,
  32'h3d3f0366 /* (31, 10, 24) */,
  32'h3d5ef675 /* (27, 10, 24) */,
  32'h3da590e9 /* (23, 10, 24) */,
  32'h3e085939 /* (19, 10, 24) */,
  32'h3e135573 /* (15, 10, 24) */,
  32'h3dd7e578 /* (11, 10, 24) */,
  32'h3d83c517 /* (7, 10, 24) */,
  32'h3d48bc7e /* (3, 10, 24) */,
  32'h3d169650 /* (31, 6, 24) */,
  32'h3d22af34 /* (27, 6, 24) */,
  32'h3d584c0c /* (23, 6, 24) */,
  32'h3da2e7a9 /* (19, 6, 24) */,
  32'h3daa3349 /* (15, 6, 24) */,
  32'h3d865b59 /* (11, 6, 24) */,
  32'h3d35cd98 /* (7, 6, 24) */,
  32'h3d19bf4b /* (3, 6, 24) */,
  32'h3d15ce12 /* (31, 2, 24) */,
  32'h3d149b5c /* (27, 2, 24) */,
  32'h3d3291f6 /* (23, 2, 24) */,
  32'h3d7b52f8 /* (19, 2, 24) */,
  32'h3d804df8 /* (15, 2, 24) */,
  32'h3d558b1c /* (11, 2, 24) */,
  32'h3d1d59b0 /* (7, 2, 24) */,
  32'h3d13e9f7 /* (3, 2, 24) */,
  32'h3d1cac31 /* (31, 30, 20) */,
  32'h3d346b02 /* (27, 30, 20) */,
  32'h3d833332 /* (23, 30, 20) */,
  32'h3dd42d31 /* (19, 30, 20) */,
  32'h3de39dff /* (15, 30, 20) */,
  32'h3da96c08 /* (11, 30, 20) */,
  32'h3d530d8e /* (7, 30, 20) */,
  32'h3d23d587 /* (3, 30, 20) */,
  32'h3d3dc5f0 /* (31, 26, 20) */,
  32'h3d6007ad /* (27, 26, 20) */,
  32'h3da96159 /* (23, 26, 20) */,
  32'h3e0dc95f /* (19, 26, 20) */,
  32'h3e1a3a56 /* (15, 26, 20) */,
  32'h3ddec971 /* (11, 26, 20) */,
  32'h3d859348 /* (7, 26, 20) */,
  32'h3d48406d /* (3, 26, 20) */,
  32'h3d91435f /* (31, 22, 20) */,
  32'h3db0e528 /* (27, 22, 20) */,
  32'h3e0cf021 /* (23, 22, 20) */,
  32'h3e7848b5 /* (19, 22, 20) */,
  32'h3e89fde5 /* (15, 22, 20) */,
  32'h3e3e5baf /* (11, 22, 20) */,
  32'h3dd85675 /* (7, 22, 20) */,
  32'h3d9aff71 /* (3, 22, 20) */,
  32'h3ddbed5a /* (31, 18, 20) */,
  32'h3e095be4 /* (27, 18, 20) */,
  32'h3e654448 /* (23, 18, 20) */,
  32'h3ed441df /* (19, 18, 20) */,
  32'h3ef15f91 /* (15, 18, 20) */,
  32'h3e9ecc49 /* (11, 18, 20) */,
  32'h3e2baf50 /* (7, 18, 20) */,
  32'h3decc5e8 /* (3, 18, 20) */,
  32'h3ddbed5a /* (31, 14, 20) */,
  32'h3e095be4 /* (27, 14, 20) */,
  32'h3e654448 /* (23, 14, 20) */,
  32'h3ed441df /* (19, 14, 20) */,
  32'h3ef15f91 /* (15, 14, 20) */,
  32'h3e9ecc49 /* (11, 14, 20) */,
  32'h3e2baf50 /* (7, 14, 20) */,
  32'h3decc5e8 /* (3, 14, 20) */,
  32'h3d91435f /* (31, 10, 20) */,
  32'h3db0e528 /* (27, 10, 20) */,
  32'h3e0cf021 /* (23, 10, 20) */,
  32'h3e7848b5 /* (19, 10, 20) */,
  32'h3e89fde5 /* (15, 10, 20) */,
  32'h3e3e5baf /* (11, 10, 20) */,
  32'h3dd85675 /* (7, 10, 20) */,
  32'h3d9aff71 /* (3, 10, 20) */,
  32'h3d3dc5f0 /* (31, 6, 20) */,
  32'h3d6007ad /* (27, 6, 20) */,
  32'h3da96159 /* (23, 6, 20) */,
  32'h3e0dc95f /* (19, 6, 20) */,
  32'h3e1a3a56 /* (15, 6, 20) */,
  32'h3ddec971 /* (11, 6, 20) */,
  32'h3d859348 /* (7, 6, 20) */,
  32'h3d48406d /* (3, 6, 20) */,
  32'h3d1cac31 /* (31, 2, 20) */,
  32'h3d346b02 /* (27, 2, 20) */,
  32'h3d833332 /* (23, 2, 20) */,
  32'h3dd42d31 /* (19, 2, 20) */,
  32'h3de39dff /* (15, 2, 20) */,
  32'h3da96c08 /* (11, 2, 20) */,
  32'h3d530d8e /* (7, 2, 20) */,
  32'h3d23d587 /* (3, 2, 20) */,
  32'h3d09dfab /* (31, 30, 16) */,
  32'h3d28d1e5 /* (27, 30, 16) */,
  32'h3d87d16b /* (23, 30, 16) */,
  32'h3df1ae3d /* (19, 30, 16) */,
  32'h3e06ec2e /* (15, 30, 16) */,
  32'h3db86416 /* (11, 30, 16) */,
  32'h3d4f6a6e /* (7, 30, 16) */,
  32'h3d13661d /* (3, 30, 16) */,
  32'h3d34b66a /* (31, 26, 16) */,
  32'h3d5f53fb /* (27, 26, 16) */,
  32'h3db6b309 /* (23, 26, 16) */,
  32'h3e2576a9 /* (19, 26, 16) */,
  32'h3e3a3d1a /* (15, 26, 16) */,
  32'h3dfa4afe /* (11, 26, 16) */,
  32'h3d8a46e7 /* (7, 26, 16) */,
  32'h3d41d3ae /* (3, 26, 16) */,
  32'h3d99ac24 /* (31, 22, 16) */,
  32'h3dc0863e /* (27, 22, 16) */,
  32'h3e21930d /* (23, 22, 16) */,
  32'h3e968a40 /* (19, 22, 16) */,
  32'h3eabb572 /* (15, 22, 16) */,
  32'h3e60898b /* (11, 22, 16) */,
  32'h3df142da /* (7, 22, 16) */,
  32'h3da59d10 /* (3, 22, 16) */,
  32'h3dff32bb /* (31, 18, 16) */,
  32'h3e2205a1 /* (27, 18, 16) */,
  32'h3e8b9344 /* (23, 18, 16) */,
  32'h3f06176f /* (19, 18, 16) */,
  32'h3f1b42bd /* (15, 18, 16) */,
  32'h3ec4f0a1 /* (11, 18, 16) */,
  32'h3e4d7ce8 /* (7, 18, 16) */,
  32'h3e0a27e7 /* (3, 18, 16) */,
  32'h3dff32bb /* (31, 14, 16) */,
  32'h3e2205a1 /* (27, 14, 16) */,
  32'h3e8b9344 /* (23, 14, 16) */,
  32'h3f06176f /* (19, 14, 16) */,
  32'h3f1b42bd /* (15, 14, 16) */,
  32'h3ec4f0a1 /* (11, 14, 16) */,
  32'h3e4d7ce8 /* (7, 14, 16) */,
  32'h3e0a27e7 /* (3, 14, 16) */,
  32'h3d99ac24 /* (31, 10, 16) */,
  32'h3dc0863e /* (27, 10, 16) */,
  32'h3e21930d /* (23, 10, 16) */,
  32'h3e968a40 /* (19, 10, 16) */,
  32'h3eabb572 /* (15, 10, 16) */,
  32'h3e60898b /* (11, 10, 16) */,
  32'h3df142da /* (7, 10, 16) */,
  32'h3da59d10 /* (3, 10, 16) */,
  32'h3d34b66a /* (31, 6, 16) */,
  32'h3d5f53fb /* (27, 6, 16) */,
  32'h3db6b309 /* (23, 6, 16) */,
  32'h3e2576a9 /* (19, 6, 16) */,
  32'h3e3a3d1a /* (15, 6, 16) */,
  32'h3dfa4afe /* (11, 6, 16) */,
  32'h3d8a46e7 /* (7, 6, 16) */,
  32'h3d41d3ae /* (3, 6, 16) */,
  32'h3d09dfab /* (31, 2, 16) */,
  32'h3d28d1e5 /* (27, 2, 16) */,
  32'h3d87d16b /* (23, 2, 16) */,
  32'h3df1ae3d /* (19, 2, 16) */,
  32'h3e06ec2e /* (15, 2, 16) */,
  32'h3db86416 /* (11, 2, 16) */,
  32'h3d4f6a6e /* (7, 2, 16) */,
  32'h3d13661d /* (3, 2, 16) */,
  32'h3d1cac31 /* (31, 30, 12) */,
  32'h3d346b02 /* (27, 30, 12) */,
  32'h3d833332 /* (23, 30, 12) */,
  32'h3dd42d31 /* (19, 30, 12) */,
  32'h3de39dff /* (15, 30, 12) */,
  32'h3da96c08 /* (11, 30, 12) */,
  32'h3d530d8e /* (7, 30, 12) */,
  32'h3d23d587 /* (3, 30, 12) */,
  32'h3d3dc5f0 /* (31, 26, 12) */,
  32'h3d6007ad /* (27, 26, 12) */,
  32'h3da96159 /* (23, 26, 12) */,
  32'h3e0dc95f /* (19, 26, 12) */,
  32'h3e1a3a56 /* (15, 26, 12) */,
  32'h3ddec971 /* (11, 26, 12) */,
  32'h3d859348 /* (7, 26, 12) */,
  32'h3d48406d /* (3, 26, 12) */,
  32'h3d91435f /* (31, 22, 12) */,
  32'h3db0e528 /* (27, 22, 12) */,
  32'h3e0cf021 /* (23, 22, 12) */,
  32'h3e7848b5 /* (19, 22, 12) */,
  32'h3e89fde5 /* (15, 22, 12) */,
  32'h3e3e5baf /* (11, 22, 12) */,
  32'h3dd85675 /* (7, 22, 12) */,
  32'h3d9aff71 /* (3, 22, 12) */,
  32'h3ddbed5a /* (31, 18, 12) */,
  32'h3e095be4 /* (27, 18, 12) */,
  32'h3e654448 /* (23, 18, 12) */,
  32'h3ed441df /* (19, 18, 12) */,
  32'h3ef15f91 /* (15, 18, 12) */,
  32'h3e9ecc49 /* (11, 18, 12) */,
  32'h3e2baf50 /* (7, 18, 12) */,
  32'h3decc5e8 /* (3, 18, 12) */,
  32'h3ddbed5a /* (31, 14, 12) */,
  32'h3e095be4 /* (27, 14, 12) */,
  32'h3e654448 /* (23, 14, 12) */,
  32'h3ed441df /* (19, 14, 12) */,
  32'h3ef15f91 /* (15, 14, 12) */,
  32'h3e9ecc49 /* (11, 14, 12) */,
  32'h3e2baf50 /* (7, 14, 12) */,
  32'h3decc5e8 /* (3, 14, 12) */,
  32'h3d91435f /* (31, 10, 12) */,
  32'h3db0e528 /* (27, 10, 12) */,
  32'h3e0cf021 /* (23, 10, 12) */,
  32'h3e7848b5 /* (19, 10, 12) */,
  32'h3e89fde5 /* (15, 10, 12) */,
  32'h3e3e5baf /* (11, 10, 12) */,
  32'h3dd85675 /* (7, 10, 12) */,
  32'h3d9aff71 /* (3, 10, 12) */,
  32'h3d3dc5f0 /* (31, 6, 12) */,
  32'h3d6007ad /* (27, 6, 12) */,
  32'h3da96159 /* (23, 6, 12) */,
  32'h3e0dc95f /* (19, 6, 12) */,
  32'h3e1a3a56 /* (15, 6, 12) */,
  32'h3ddec971 /* (11, 6, 12) */,
  32'h3d859348 /* (7, 6, 12) */,
  32'h3d48406d /* (3, 6, 12) */,
  32'h3d1cac31 /* (31, 2, 12) */,
  32'h3d346b02 /* (27, 2, 12) */,
  32'h3d833332 /* (23, 2, 12) */,
  32'h3dd42d31 /* (19, 2, 12) */,
  32'h3de39dff /* (15, 2, 12) */,
  32'h3da96c08 /* (11, 2, 12) */,
  32'h3d530d8e /* (7, 2, 12) */,
  32'h3d23d587 /* (3, 2, 12) */,
  32'h3d15ce12 /* (31, 30, 8) */,
  32'h3d149b5c /* (27, 30, 8) */,
  32'h3d3291f6 /* (23, 30, 8) */,
  32'h3d7b52f8 /* (19, 30, 8) */,
  32'h3d804df8 /* (15, 30, 8) */,
  32'h3d558b1c /* (11, 30, 8) */,
  32'h3d1d59b0 /* (7, 30, 8) */,
  32'h3d13e9f7 /* (3, 30, 8) */,
  32'h3d169650 /* (31, 26, 8) */,
  32'h3d22af34 /* (27, 26, 8) */,
  32'h3d584c0c /* (23, 26, 8) */,
  32'h3da2e7a9 /* (19, 26, 8) */,
  32'h3daa3349 /* (15, 26, 8) */,
  32'h3d865b59 /* (11, 26, 8) */,
  32'h3d35cd98 /* (7, 26, 8) */,
  32'h3d19bf4b /* (3, 26, 8) */,
  32'h3d3f0366 /* (31, 22, 8) */,
  32'h3d5ef675 /* (27, 22, 8) */,
  32'h3da590e9 /* (23, 22, 8) */,
  32'h3e085939 /* (19, 22, 8) */,
  32'h3e135573 /* (15, 22, 8) */,
  32'h3dd7e578 /* (11, 22, 8) */,
  32'h3d83c517 /* (7, 22, 8) */,
  32'h3d48bc7e /* (3, 22, 8) */,
  32'h3d7e759f /* (31, 18, 8) */,
  32'h3d9bc970 /* (27, 18, 8) */,
  32'h3dfaaa60 /* (23, 18, 8) */,
  32'h3e5f05ce /* (19, 18, 8) */,
  32'h3e79034c /* (15, 18, 8) */,
  32'h3e2a27e4 /* (11, 18, 8) */,
  32'h3dbf672f /* (7, 18, 8) */,
  32'h3d880501 /* (3, 18, 8) */,
  32'h3d7e759f /* (31, 14, 8) */,
  32'h3d9bc970 /* (27, 14, 8) */,
  32'h3dfaaa60 /* (23, 14, 8) */,
  32'h3e5f05ce /* (19, 14, 8) */,
  32'h3e79034c /* (15, 14, 8) */,
  32'h3e2a27e4 /* (11, 14, 8) */,
  32'h3dbf672f /* (7, 14, 8) */,
  32'h3d880501 /* (3, 14, 8) */,
  32'h3d3f0366 /* (31, 10, 8) */,
  32'h3d5ef675 /* (27, 10, 8) */,
  32'h3da590e9 /* (23, 10, 8) */,
  32'h3e085939 /* (19, 10, 8) */,
  32'h3e135573 /* (15, 10, 8) */,
  32'h3dd7e578 /* (11, 10, 8) */,
  32'h3d83c517 /* (7, 10, 8) */,
  32'h3d48bc7e /* (3, 10, 8) */,
  32'h3d169650 /* (31, 6, 8) */,
  32'h3d22af34 /* (27, 6, 8) */,
  32'h3d584c0c /* (23, 6, 8) */,
  32'h3da2e7a9 /* (19, 6, 8) */,
  32'h3daa3349 /* (15, 6, 8) */,
  32'h3d865b59 /* (11, 6, 8) */,
  32'h3d35cd98 /* (7, 6, 8) */,
  32'h3d19bf4b /* (3, 6, 8) */,
  32'h3d15ce12 /* (31, 2, 8) */,
  32'h3d149b5c /* (27, 2, 8) */,
  32'h3d3291f6 /* (23, 2, 8) */,
  32'h3d7b52f8 /* (19, 2, 8) */,
  32'h3d804df8 /* (15, 2, 8) */,
  32'h3d558b1c /* (11, 2, 8) */,
  32'h3d1d59b0 /* (7, 2, 8) */,
  32'h3d13e9f7 /* (3, 2, 8) */,
  32'h3d8b1391 /* (31, 30, 4) */,
  32'h3d2d8e0e /* (27, 30, 4) */,
  32'h3d14de35 /* (23, 30, 4) */,
  32'h3d3217f4 /* (19, 30, 4) */,
  32'h3d2d6bba /* (15, 30, 4) */,
  32'h3d21c128 /* (11, 30, 4) */,
  32'h3d16c6a3 /* (7, 30, 4) */,
  32'h3d5defd3 /* (3, 30, 4) */,
  32'h3d222a9c /* (31, 26, 4) */,
  32'h3d153e19 /* (27, 26, 4) */,
  32'h3d2657dd /* (23, 26, 4) */,
  32'h3d601ae9 /* (19, 26, 4) */,
  32'h3d61b1de /* (15, 26, 4) */,
  32'h3d41fb9f /* (11, 26, 4) */,
  32'h3d17902e /* (7, 26, 4) */,
  32'h3d1b3fff /* (3, 26, 4) */,
  32'h3d1839e3 /* (31, 22, 4) */,
  32'h3d28e3b2 /* (27, 22, 4) */,
  32'h3d68b7a2 /* (23, 22, 4) */,
  32'h3db40e50 /* (19, 22, 4) */,
  32'h3dbdf4f8 /* (15, 22, 4) */,
  32'h3d92b699 /* (11, 22, 4) */,
  32'h3d404057 /* (7, 22, 4) */,
  32'h3d1cff11 /* (3, 22, 4) */,
  32'h3d303352 /* (31, 18, 4) */,
  32'h3d53bb31 /* (27, 18, 4) */,
  32'h3da4db8a /* (23, 18, 4) */,
  32'h3e0de89e /* (19, 18, 4) */,
  32'h3e1c2ca1 /* (15, 18, 4) */,
  32'h3ddc0819 /* (11, 18, 4) */,
  32'h3d800deb /* (7, 18, 4) */,
  32'h3d3b1e93 /* (3, 18, 4) */,
  32'h3d303352 /* (31, 14, 4) */,
  32'h3d53bb31 /* (27, 14, 4) */,
  32'h3da4db8a /* (23, 14, 4) */,
  32'h3e0de89e /* (19, 14, 4) */,
  32'h3e1c2ca1 /* (15, 14, 4) */,
  32'h3ddc0819 /* (11, 14, 4) */,
  32'h3d800deb /* (7, 14, 4) */,
  32'h3d3b1e93 /* (3, 14, 4) */,
  32'h3d1839e3 /* (31, 10, 4) */,
  32'h3d28e3b2 /* (27, 10, 4) */,
  32'h3d68b7a2 /* (23, 10, 4) */,
  32'h3db40e50 /* (19, 10, 4) */,
  32'h3dbdf4f8 /* (15, 10, 4) */,
  32'h3d92b699 /* (11, 10, 4) */,
  32'h3d404057 /* (7, 10, 4) */,
  32'h3d1cff11 /* (3, 10, 4) */,
  32'h3d222a9c /* (31, 6, 4) */,
  32'h3d153e19 /* (27, 6, 4) */,
  32'h3d2657dd /* (23, 6, 4) */,
  32'h3d601ae9 /* (19, 6, 4) */,
  32'h3d61b1de /* (15, 6, 4) */,
  32'h3d41fb9f /* (11, 6, 4) */,
  32'h3d17902e /* (7, 6, 4) */,
  32'h3d1b3fff /* (3, 6, 4) */,
  32'h3d8b1391 /* (31, 2, 4) */,
  32'h3d2d8e0e /* (27, 2, 4) */,
  32'h3d14de35 /* (23, 2, 4) */,
  32'h3d3217f4 /* (19, 2, 4) */,
  32'h3d2d6bba /* (15, 2, 4) */,
  32'h3d21c128 /* (11, 2, 4) */,
  32'h3d16c6a3 /* (7, 2, 4) */,
  32'h3d5defd3 /* (3, 2, 4) */,
  32'h3e709592 /* (31, 30, 0) */,
  32'h3d5dd7d1 /* (27, 30, 0) */,
  32'h3d11b684 /* (23, 30, 0) */,
  32'h3d2045b1 /* (19, 30, 0) */,
  32'h3d18d610 /* (15, 30, 0) */,
  32'h3d164ce1 /* (11, 30, 0) */,
  32'h3d21b235 /* (7, 30, 0) */,
  32'h3dcbea25 /* (3, 30, 0) */,
  32'h3d3f59b8 /* (31, 26, 0) */,
  32'h3d1b2f33 /* (27, 26, 0) */,
  32'h3d1bc36a /* (23, 26, 0) */,
  32'h3d4703b2 /* (19, 26, 0) */,
  32'h3d455011 /* (15, 26, 0) */,
  32'h3d3013e2 /* (11, 26, 0) */,
  32'h3d1459dd /* (7, 26, 0) */,
  32'h3d2d5b95 /* (3, 26, 0) */,
  32'h3d1142bb /* (31, 22, 0) */,
  32'h3d1cee15 /* (27, 22, 0) */,
  32'h3d50a575 /* (23, 22, 0) */,
  32'h3d9d248b /* (19, 22, 0) */,
  32'h3da42e1b /* (15, 22, 0) */,
  32'h3d819abc /* (11, 22, 0) */,
  32'h3d2f5f5a /* (7, 22, 0) */,
  32'h3d144f19 /* (3, 22, 0) */,
  32'h3d1ceee6 /* (31, 18, 0) */,
  32'h3d3b0a55 /* (27, 18, 0) */,
  32'h3d8fa52c /* (23, 18, 0) */,
  32'h3df40add /* (19, 18, 0) */,
  32'h3e05899d /* (15, 18, 0) */,
  32'h3dbe661f /* (11, 18, 0) */,
  32'h3d60bf24 /* (7, 18, 0) */,
  32'h3d262b6e /* (3, 18, 0) */,
  32'h3d1ceee6 /* (31, 14, 0) */,
  32'h3d3b0a55 /* (27, 14, 0) */,
  32'h3d8fa52c /* (23, 14, 0) */,
  32'h3df40add /* (19, 14, 0) */,
  32'h3e05899d /* (15, 14, 0) */,
  32'h3dbe661f /* (11, 14, 0) */,
  32'h3d60bf24 /* (7, 14, 0) */,
  32'h3d262b6e /* (3, 14, 0) */,
  32'h3d1142bb /* (31, 10, 0) */,
  32'h3d1cee15 /* (27, 10, 0) */,
  32'h3d50a575 /* (23, 10, 0) */,
  32'h3d9d248b /* (19, 10, 0) */,
  32'h3da42e1b /* (15, 10, 0) */,
  32'h3d819abc /* (11, 10, 0) */,
  32'h3d2f5f5a /* (7, 10, 0) */,
  32'h3d144f19 /* (3, 10, 0) */,
  32'h3d3f59b8 /* (31, 6, 0) */,
  32'h3d1b2f33 /* (27, 6, 0) */,
  32'h3d1bc36a /* (23, 6, 0) */,
  32'h3d4703b2 /* (19, 6, 0) */,
  32'h3d455011 /* (15, 6, 0) */,
  32'h3d3013e2 /* (11, 6, 0) */,
  32'h3d1459dd /* (7, 6, 0) */,
  32'h3d2d5b95 /* (3, 6, 0) */,
  32'h3e709592 /* (31, 2, 0) */,
  32'h3d5dd7d1 /* (27, 2, 0) */,
  32'h3d11b684 /* (23, 2, 0) */,
  32'h3d2045b1 /* (19, 2, 0) */,
  32'h3d18d610 /* (15, 2, 0) */,
  32'h3d164ce1 /* (11, 2, 0) */,
  32'h3d21b235 /* (7, 2, 0) */,
  32'h3dcbea25 /* (3, 2, 0) */,
  32'h3d7c66bd /* (30, 30, 28) */,
  32'h3d1f2a5d /* (26, 30, 28) */,
  32'h3d19eb69 /* (22, 30, 28) */,
  32'h3d3430e1 /* (18, 30, 28) */,
  32'h3d3430e1 /* (14, 30, 28) */,
  32'h3d19eb69 /* (10, 30, 28) */,
  32'h3d1f2a5d /* (6, 30, 28) */,
  32'h3d7c66bd /* (2, 30, 28) */,
  32'h3d1f2a5d /* (30, 26, 28) */,
  32'h3d1508f6 /* (26, 26, 28) */,
  32'h3d32cc97 /* (22, 26, 28) */,
  32'h3d66ec8b /* (18, 26, 28) */,
  32'h3d66ec8b /* (14, 26, 28) */,
  32'h3d32cc97 /* (10, 26, 28) */,
  32'h3d1508f6 /* (6, 26, 28) */,
  32'h3d1f2a5d /* (2, 26, 28) */,
  32'h3d19eb69 /* (30, 22, 28) */,
  32'h3d32cc97 /* (26, 22, 28) */,
  32'h3d825da2 /* (22, 22, 28) */,
  32'h3dbe2f24 /* (18, 22, 28) */,
  32'h3dbe2f24 /* (14, 22, 28) */,
  32'h3d825da2 /* (10, 22, 28) */,
  32'h3d32cc97 /* (6, 22, 28) */,
  32'h3d19eb69 /* (2, 22, 28) */,
  32'h3d3430e1 /* (30, 18, 28) */,
  32'h3d66ec8b /* (26, 18, 28) */,
  32'h3dbe2f24 /* (22, 18, 28) */,
  32'h3e193b79 /* (18, 18, 28) */,
  32'h3e193b79 /* (14, 18, 28) */,
  32'h3dbe2f24 /* (10, 18, 28) */,
  32'h3d66ec8b /* (6, 18, 28) */,
  32'h3d3430e1 /* (2, 18, 28) */,
  32'h3d3430e1 /* (30, 14, 28) */,
  32'h3d66ec8b /* (26, 14, 28) */,
  32'h3dbe2f24 /* (22, 14, 28) */,
  32'h3e193b79 /* (18, 14, 28) */,
  32'h3e193b79 /* (14, 14, 28) */,
  32'h3dbe2f24 /* (10, 14, 28) */,
  32'h3d66ec8b /* (6, 14, 28) */,
  32'h3d3430e1 /* (2, 14, 28) */,
  32'h3d19eb69 /* (30, 10, 28) */,
  32'h3d32cc97 /* (26, 10, 28) */,
  32'h3d825da2 /* (22, 10, 28) */,
  32'h3dbe2f24 /* (18, 10, 28) */,
  32'h3dbe2f24 /* (14, 10, 28) */,
  32'h3d825da2 /* (10, 10, 28) */,
  32'h3d32cc97 /* (6, 10, 28) */,
  32'h3d19eb69 /* (2, 10, 28) */,
  32'h3d1f2a5d /* (30, 6, 28) */,
  32'h3d1508f6 /* (26, 6, 28) */,
  32'h3d32cc97 /* (22, 6, 28) */,
  32'h3d66ec8b /* (18, 6, 28) */,
  32'h3d66ec8b /* (14, 6, 28) */,
  32'h3d32cc97 /* (10, 6, 28) */,
  32'h3d1508f6 /* (6, 6, 28) */,
  32'h3d1f2a5d /* (2, 6, 28) */,
  32'h3d7c66bd /* (30, 2, 28) */,
  32'h3d1f2a5d /* (26, 2, 28) */,
  32'h3d19eb69 /* (22, 2, 28) */,
  32'h3d3430e1 /* (18, 2, 28) */,
  32'h3d3430e1 /* (14, 2, 28) */,
  32'h3d19eb69 /* (10, 2, 28) */,
  32'h3d1f2a5d /* (6, 2, 28) */,
  32'h3d7c66bd /* (2, 2, 28) */,
  32'h3d14e1d9 /* (30, 30, 24) */,
  32'h3d17a967 /* (26, 30, 24) */,
  32'h3d428d9a /* (22, 30, 24) */,
  32'h3d8271c0 /* (18, 30, 24) */,
  32'h3d8271c0 /* (14, 30, 24) */,
  32'h3d428d9a /* (10, 30, 24) */,
  32'h3d17a967 /* (6, 30, 24) */,
  32'h3d14e1d9 /* (2, 30, 24) */,
  32'h3d17a967 /* (30, 26, 24) */,
  32'h3d2aa638 /* (26, 26, 24) */,
  32'h3d7076ff /* (22, 26, 24) */,
  32'h3dab2ff1 /* (18, 26, 24) */,
  32'h3dab2ff1 /* (14, 26, 24) */,
  32'h3d7076ff /* (10, 26, 24) */,
  32'h3d2aa638 /* (6, 26, 24) */,
  32'h3d17a967 /* (2, 26, 24) */,
  32'h3d428d9a /* (30, 22, 24) */,
  32'h3d7076ff /* (26, 22, 24) */,
  32'h3dbcbfdf /* (22, 22, 24) */,
  32'h3e11d65f /* (18, 22, 24) */,
  32'h3e11d65f /* (14, 22, 24) */,
  32'h3dbcbfdf /* (10, 22, 24) */,
  32'h3d7076ff /* (6, 22, 24) */,
  32'h3d428d9a /* (2, 22, 24) */,
  32'h3d8271c0 /* (30, 18, 24) */,
  32'h3dab2ff1 /* (26, 18, 24) */,
  32'h3e11d65f /* (22, 18, 24) */,
  32'h3e729d82 /* (18, 18, 24) */,
  32'h3e729d82 /* (14, 18, 24) */,
  32'h3e11d65f /* (10, 18, 24) */,
  32'h3dab2ff1 /* (6, 18, 24) */,
  32'h3d8271c0 /* (2, 18, 24) */,
  32'h3d8271c0 /* (30, 14, 24) */,
  32'h3dab2ff1 /* (26, 14, 24) */,
  32'h3e11d65f /* (22, 14, 24) */,
  32'h3e729d82 /* (18, 14, 24) */,
  32'h3e729d82 /* (14, 14, 24) */,
  32'h3e11d65f /* (10, 14, 24) */,
  32'h3dab2ff1 /* (6, 14, 24) */,
  32'h3d8271c0 /* (2, 14, 24) */,
  32'h3d428d9a /* (30, 10, 24) */,
  32'h3d7076ff /* (26, 10, 24) */,
  32'h3dbcbfdf /* (22, 10, 24) */,
  32'h3e11d65f /* (18, 10, 24) */,
  32'h3e11d65f /* (14, 10, 24) */,
  32'h3dbcbfdf /* (10, 10, 24) */,
  32'h3d7076ff /* (6, 10, 24) */,
  32'h3d428d9a /* (2, 10, 24) */,
  32'h3d17a967 /* (30, 6, 24) */,
  32'h3d2aa638 /* (26, 6, 24) */,
  32'h3d7076ff /* (22, 6, 24) */,
  32'h3dab2ff1 /* (18, 6, 24) */,
  32'h3dab2ff1 /* (14, 6, 24) */,
  32'h3d7076ff /* (10, 6, 24) */,
  32'h3d2aa638 /* (6, 6, 24) */,
  32'h3d17a967 /* (2, 6, 24) */,
  32'h3d14e1d9 /* (30, 2, 24) */,
  32'h3d17a967 /* (26, 2, 24) */,
  32'h3d428d9a /* (22, 2, 24) */,
  32'h3d8271c0 /* (18, 2, 24) */,
  32'h3d8271c0 /* (14, 2, 24) */,
  32'h3d428d9a /* (10, 2, 24) */,
  32'h3d17a967 /* (6, 2, 24) */,
  32'h3d14e1d9 /* (2, 2, 24) */,
  32'h3d1f454c /* (30, 30, 20) */,
  32'h3d41987e /* (26, 30, 20) */,
  32'h3d94d2ae /* (22, 30, 20) */,
  32'h3de2162b /* (18, 30, 20) */,
  32'h3de2162b /* (14, 30, 20) */,
  32'h3d94d2ae /* (10, 30, 20) */,
  32'h3d41987e /* (6, 30, 20) */,
  32'h3d1f454c /* (2, 30, 20) */,
  32'h3d41987e /* (30, 26, 20) */,
  32'h3d72a853 /* (26, 26, 20) */,
  32'h3dc1f419 /* (22, 26, 20) */,
  32'h3e182d5a /* (18, 26, 20) */,
  32'h3e182d5a /* (14, 26, 20) */,
  32'h3dc1f419 /* (10, 26, 20) */,
  32'h3d72a853 /* (6, 26, 20) */,
  32'h3d41987e /* (2, 26, 20) */,
  32'h3d94d2ae /* (30, 22, 20) */,
  32'h3dc1f419 /* (26, 22, 20) */,
  32'h3e239217 /* (22, 22, 20) */,
  32'h3e86bd25 /* (18, 22, 20) */,
  32'h3e86bd25 /* (14, 22, 20) */,
  32'h3e239217 /* (10, 22, 20) */,
  32'h3dc1f419 /* (6, 22, 20) */,
  32'h3d94d2ae /* (2, 22, 20) */,
  32'h3de2162b /* (30, 18, 20) */,
  32'h3e182d5a /* (26, 18, 20) */,
  32'h3e86bd25 /* (22, 18, 20) */,
  32'h3ee912bc /* (18, 18, 20) */,
  32'h3ee912bc /* (14, 18, 20) */,
  32'h3e86bd25 /* (10, 18, 20) */,
  32'h3e182d5a /* (6, 18, 20) */,
  32'h3de2162b /* (2, 18, 20) */,
  32'h3de2162b /* (30, 14, 20) */,
  32'h3e182d5a /* (26, 14, 20) */,
  32'h3e86bd25 /* (22, 14, 20) */,
  32'h3ee912bc /* (18, 14, 20) */,
  32'h3ee912bc /* (14, 14, 20) */,
  32'h3e86bd25 /* (10, 14, 20) */,
  32'h3e182d5a /* (6, 14, 20) */,
  32'h3de2162b /* (2, 14, 20) */,
  32'h3d94d2ae /* (30, 10, 20) */,
  32'h3dc1f419 /* (26, 10, 20) */,
  32'h3e239217 /* (22, 10, 20) */,
  32'h3e86bd25 /* (18, 10, 20) */,
  32'h3e86bd25 /* (14, 10, 20) */,
  32'h3e239217 /* (10, 10, 20) */,
  32'h3dc1f419 /* (6, 10, 20) */,
  32'h3d94d2ae /* (2, 10, 20) */,
  32'h3d41987e /* (30, 6, 20) */,
  32'h3d72a853 /* (26, 6, 20) */,
  32'h3dc1f419 /* (22, 6, 20) */,
  32'h3e182d5a /* (18, 6, 20) */,
  32'h3e182d5a /* (14, 6, 20) */,
  32'h3dc1f419 /* (10, 6, 20) */,
  32'h3d72a853 /* (6, 6, 20) */,
  32'h3d41987e /* (2, 6, 20) */,
  32'h3d1f454c /* (30, 2, 20) */,
  32'h3d41987e /* (26, 2, 20) */,
  32'h3d94d2ae /* (22, 2, 20) */,
  32'h3de2162b /* (18, 2, 20) */,
  32'h3de2162b /* (14, 2, 20) */,
  32'h3d94d2ae /* (10, 2, 20) */,
  32'h3d41987e /* (6, 2, 20) */,
  32'h3d1f454c /* (2, 2, 20) */,
  32'h3d0d5b74 /* (30, 30, 16) */,
  32'h3d39823a /* (26, 30, 16) */,
  32'h3d9e09be /* (22, 30, 16) */,
  32'h3e0374c7 /* (18, 30, 16) */,
  32'h3e0374c7 /* (14, 30, 16) */,
  32'h3d9e09be /* (10, 30, 16) */,
  32'h3d39823a /* (6, 30, 16) */,
  32'h3d0d5b74 /* (2, 30, 16) */,
  32'h3d39823a /* (30, 26, 16) */,
  32'h3d765452 /* (26, 26, 16) */,
  32'h3dd58e62 /* (22, 26, 16) */,
  32'h3e34be0d /* (18, 26, 16) */,
  32'h3e34be0d /* (14, 26, 16) */,
  32'h3dd58e62 /* (10, 26, 16) */,
  32'h3d765452 /* (6, 26, 16) */,
  32'h3d39823a /* (2, 26, 16) */,
  32'h3d9e09be /* (30, 22, 16) */,
  32'h3dd58e62 /* (26, 22, 16) */,
  32'h3e3e36ae /* (22, 22, 16) */,
  32'h3ea58eba /* (18, 22, 16) */,
  32'h3ea58eba /* (14, 22, 16) */,
  32'h3e3e36ae /* (10, 22, 16) */,
  32'h3dd58e62 /* (6, 22, 16) */,
  32'h3d9e09be /* (2, 22, 16) */,
  32'h3e0374c7 /* (30, 18, 16) */,
  32'h3e34be0d /* (26, 18, 16) */,
  32'h3ea58eba /* (22, 18, 16) */,
  32'h3f14977b /* (18, 18, 16) */,
  32'h3f14977b /* (14, 18, 16) */,
  32'h3ea58eba /* (10, 18, 16) */,
  32'h3e34be0d /* (6, 18, 16) */,
  32'h3e0374c7 /* (2, 18, 16) */,
  32'h3e0374c7 /* (30, 14, 16) */,
  32'h3e34be0d /* (26, 14, 16) */,
  32'h3ea58eba /* (22, 14, 16) */,
  32'h3f14977b /* (18, 14, 16) */,
  32'h3f14977b /* (14, 14, 16) */,
  32'h3ea58eba /* (10, 14, 16) */,
  32'h3e34be0d /* (6, 14, 16) */,
  32'h3e0374c7 /* (2, 14, 16) */,
  32'h3d9e09be /* (30, 10, 16) */,
  32'h3dd58e62 /* (26, 10, 16) */,
  32'h3e3e36ae /* (22, 10, 16) */,
  32'h3ea58eba /* (18, 10, 16) */,
  32'h3ea58eba /* (14, 10, 16) */,
  32'h3e3e36ae /* (10, 10, 16) */,
  32'h3dd58e62 /* (6, 10, 16) */,
  32'h3d9e09be /* (2, 10, 16) */,
  32'h3d39823a /* (30, 6, 16) */,
  32'h3d765452 /* (26, 6, 16) */,
  32'h3dd58e62 /* (22, 6, 16) */,
  32'h3e34be0d /* (18, 6, 16) */,
  32'h3e34be0d /* (14, 6, 16) */,
  32'h3dd58e62 /* (10, 6, 16) */,
  32'h3d765452 /* (6, 6, 16) */,
  32'h3d39823a /* (2, 6, 16) */,
  32'h3d0d5b74 /* (30, 2, 16) */,
  32'h3d39823a /* (26, 2, 16) */,
  32'h3d9e09be /* (22, 2, 16) */,
  32'h3e0374c7 /* (18, 2, 16) */,
  32'h3e0374c7 /* (14, 2, 16) */,
  32'h3d9e09be /* (10, 2, 16) */,
  32'h3d39823a /* (6, 2, 16) */,
  32'h3d0d5b74 /* (2, 2, 16) */,
  32'h3d1f454c /* (30, 30, 12) */,
  32'h3d41987e /* (26, 30, 12) */,
  32'h3d94d2ae /* (22, 30, 12) */,
  32'h3de2162b /* (18, 30, 12) */,
  32'h3de2162b /* (14, 30, 12) */,
  32'h3d94d2ae /* (10, 30, 12) */,
  32'h3d41987e /* (6, 30, 12) */,
  32'h3d1f454c /* (2, 30, 12) */,
  32'h3d41987e /* (30, 26, 12) */,
  32'h3d72a853 /* (26, 26, 12) */,
  32'h3dc1f419 /* (22, 26, 12) */,
  32'h3e182d5a /* (18, 26, 12) */,
  32'h3e182d5a /* (14, 26, 12) */,
  32'h3dc1f419 /* (10, 26, 12) */,
  32'h3d72a853 /* (6, 26, 12) */,
  32'h3d41987e /* (2, 26, 12) */,
  32'h3d94d2ae /* (30, 22, 12) */,
  32'h3dc1f419 /* (26, 22, 12) */,
  32'h3e239217 /* (22, 22, 12) */,
  32'h3e86bd25 /* (18, 22, 12) */,
  32'h3e86bd25 /* (14, 22, 12) */,
  32'h3e239217 /* (10, 22, 12) */,
  32'h3dc1f419 /* (6, 22, 12) */,
  32'h3d94d2ae /* (2, 22, 12) */,
  32'h3de2162b /* (30, 18, 12) */,
  32'h3e182d5a /* (26, 18, 12) */,
  32'h3e86bd25 /* (22, 18, 12) */,
  32'h3ee912bc /* (18, 18, 12) */,
  32'h3ee912bc /* (14, 18, 12) */,
  32'h3e86bd25 /* (10, 18, 12) */,
  32'h3e182d5a /* (6, 18, 12) */,
  32'h3de2162b /* (2, 18, 12) */,
  32'h3de2162b /* (30, 14, 12) */,
  32'h3e182d5a /* (26, 14, 12) */,
  32'h3e86bd25 /* (22, 14, 12) */,
  32'h3ee912bc /* (18, 14, 12) */,
  32'h3ee912bc /* (14, 14, 12) */,
  32'h3e86bd25 /* (10, 14, 12) */,
  32'h3e182d5a /* (6, 14, 12) */,
  32'h3de2162b /* (2, 14, 12) */,
  32'h3d94d2ae /* (30, 10, 12) */,
  32'h3dc1f419 /* (26, 10, 12) */,
  32'h3e239217 /* (22, 10, 12) */,
  32'h3e86bd25 /* (18, 10, 12) */,
  32'h3e86bd25 /* (14, 10, 12) */,
  32'h3e239217 /* (10, 10, 12) */,
  32'h3dc1f419 /* (6, 10, 12) */,
  32'h3d94d2ae /* (2, 10, 12) */,
  32'h3d41987e /* (30, 6, 12) */,
  32'h3d72a853 /* (26, 6, 12) */,
  32'h3dc1f419 /* (22, 6, 12) */,
  32'h3e182d5a /* (18, 6, 12) */,
  32'h3e182d5a /* (14, 6, 12) */,
  32'h3dc1f419 /* (10, 6, 12) */,
  32'h3d72a853 /* (6, 6, 12) */,
  32'h3d41987e /* (2, 6, 12) */,
  32'h3d1f454c /* (30, 2, 12) */,
  32'h3d41987e /* (26, 2, 12) */,
  32'h3d94d2ae /* (22, 2, 12) */,
  32'h3de2162b /* (18, 2, 12) */,
  32'h3de2162b /* (14, 2, 12) */,
  32'h3d94d2ae /* (10, 2, 12) */,
  32'h3d41987e /* (6, 2, 12) */,
  32'h3d1f454c /* (2, 2, 12) */,
  32'h3d14e1d9 /* (30, 30, 8) */,
  32'h3d17a967 /* (26, 30, 8) */,
  32'h3d428d9a /* (22, 30, 8) */,
  32'h3d8271c0 /* (18, 30, 8) */,
  32'h3d8271c0 /* (14, 30, 8) */,
  32'h3d428d9a /* (10, 30, 8) */,
  32'h3d17a967 /* (6, 30, 8) */,
  32'h3d14e1d9 /* (2, 30, 8) */,
  32'h3d17a967 /* (30, 26, 8) */,
  32'h3d2aa638 /* (26, 26, 8) */,
  32'h3d7076ff /* (22, 26, 8) */,
  32'h3dab2ff1 /* (18, 26, 8) */,
  32'h3dab2ff1 /* (14, 26, 8) */,
  32'h3d7076ff /* (10, 26, 8) */,
  32'h3d2aa638 /* (6, 26, 8) */,
  32'h3d17a967 /* (2, 26, 8) */,
  32'h3d428d9a /* (30, 22, 8) */,
  32'h3d7076ff /* (26, 22, 8) */,
  32'h3dbcbfdf /* (22, 22, 8) */,
  32'h3e11d65f /* (18, 22, 8) */,
  32'h3e11d65f /* (14, 22, 8) */,
  32'h3dbcbfdf /* (10, 22, 8) */,
  32'h3d7076ff /* (6, 22, 8) */,
  32'h3d428d9a /* (2, 22, 8) */,
  32'h3d8271c0 /* (30, 18, 8) */,
  32'h3dab2ff1 /* (26, 18, 8) */,
  32'h3e11d65f /* (22, 18, 8) */,
  32'h3e729d82 /* (18, 18, 8) */,
  32'h3e729d82 /* (14, 18, 8) */,
  32'h3e11d65f /* (10, 18, 8) */,
  32'h3dab2ff1 /* (6, 18, 8) */,
  32'h3d8271c0 /* (2, 18, 8) */,
  32'h3d8271c0 /* (30, 14, 8) */,
  32'h3dab2ff1 /* (26, 14, 8) */,
  32'h3e11d65f /* (22, 14, 8) */,
  32'h3e729d82 /* (18, 14, 8) */,
  32'h3e729d82 /* (14, 14, 8) */,
  32'h3e11d65f /* (10, 14, 8) */,
  32'h3dab2ff1 /* (6, 14, 8) */,
  32'h3d8271c0 /* (2, 14, 8) */,
  32'h3d428d9a /* (30, 10, 8) */,
  32'h3d7076ff /* (26, 10, 8) */,
  32'h3dbcbfdf /* (22, 10, 8) */,
  32'h3e11d65f /* (18, 10, 8) */,
  32'h3e11d65f /* (14, 10, 8) */,
  32'h3dbcbfdf /* (10, 10, 8) */,
  32'h3d7076ff /* (6, 10, 8) */,
  32'h3d428d9a /* (2, 10, 8) */,
  32'h3d17a967 /* (30, 6, 8) */,
  32'h3d2aa638 /* (26, 6, 8) */,
  32'h3d7076ff /* (22, 6, 8) */,
  32'h3dab2ff1 /* (18, 6, 8) */,
  32'h3dab2ff1 /* (14, 6, 8) */,
  32'h3d7076ff /* (10, 6, 8) */,
  32'h3d2aa638 /* (6, 6, 8) */,
  32'h3d17a967 /* (2, 6, 8) */,
  32'h3d14e1d9 /* (30, 2, 8) */,
  32'h3d17a967 /* (26, 2, 8) */,
  32'h3d428d9a /* (22, 2, 8) */,
  32'h3d8271c0 /* (18, 2, 8) */,
  32'h3d8271c0 /* (14, 2, 8) */,
  32'h3d428d9a /* (10, 2, 8) */,
  32'h3d17a967 /* (6, 2, 8) */,
  32'h3d14e1d9 /* (2, 2, 8) */,
  32'h3d7c66bd /* (30, 30, 4) */,
  32'h3d1f2a5d /* (26, 30, 4) */,
  32'h3d19eb69 /* (22, 30, 4) */,
  32'h3d3430e1 /* (18, 30, 4) */,
  32'h3d3430e1 /* (14, 30, 4) */,
  32'h3d19eb69 /* (10, 30, 4) */,
  32'h3d1f2a5d /* (6, 30, 4) */,
  32'h3d7c66bd /* (2, 30, 4) */,
  32'h3d1f2a5d /* (30, 26, 4) */,
  32'h3d1508f6 /* (26, 26, 4) */,
  32'h3d32cc97 /* (22, 26, 4) */,
  32'h3d66ec8b /* (18, 26, 4) */,
  32'h3d66ec8b /* (14, 26, 4) */,
  32'h3d32cc97 /* (10, 26, 4) */,
  32'h3d1508f6 /* (6, 26, 4) */,
  32'h3d1f2a5d /* (2, 26, 4) */,
  32'h3d19eb69 /* (30, 22, 4) */,
  32'h3d32cc97 /* (26, 22, 4) */,
  32'h3d825da2 /* (22, 22, 4) */,
  32'h3dbe2f24 /* (18, 22, 4) */,
  32'h3dbe2f24 /* (14, 22, 4) */,
  32'h3d825da2 /* (10, 22, 4) */,
  32'h3d32cc97 /* (6, 22, 4) */,
  32'h3d19eb69 /* (2, 22, 4) */,
  32'h3d3430e1 /* (30, 18, 4) */,
  32'h3d66ec8b /* (26, 18, 4) */,
  32'h3dbe2f24 /* (22, 18, 4) */,
  32'h3e193b79 /* (18, 18, 4) */,
  32'h3e193b79 /* (14, 18, 4) */,
  32'h3dbe2f24 /* (10, 18, 4) */,
  32'h3d66ec8b /* (6, 18, 4) */,
  32'h3d3430e1 /* (2, 18, 4) */,
  32'h3d3430e1 /* (30, 14, 4) */,
  32'h3d66ec8b /* (26, 14, 4) */,
  32'h3dbe2f24 /* (22, 14, 4) */,
  32'h3e193b79 /* (18, 14, 4) */,
  32'h3e193b79 /* (14, 14, 4) */,
  32'h3dbe2f24 /* (10, 14, 4) */,
  32'h3d66ec8b /* (6, 14, 4) */,
  32'h3d3430e1 /* (2, 14, 4) */,
  32'h3d19eb69 /* (30, 10, 4) */,
  32'h3d32cc97 /* (26, 10, 4) */,
  32'h3d825da2 /* (22, 10, 4) */,
  32'h3dbe2f24 /* (18, 10, 4) */,
  32'h3dbe2f24 /* (14, 10, 4) */,
  32'h3d825da2 /* (10, 10, 4) */,
  32'h3d32cc97 /* (6, 10, 4) */,
  32'h3d19eb69 /* (2, 10, 4) */,
  32'h3d1f2a5d /* (30, 6, 4) */,
  32'h3d1508f6 /* (26, 6, 4) */,
  32'h3d32cc97 /* (22, 6, 4) */,
  32'h3d66ec8b /* (18, 6, 4) */,
  32'h3d66ec8b /* (14, 6, 4) */,
  32'h3d32cc97 /* (10, 6, 4) */,
  32'h3d1508f6 /* (6, 6, 4) */,
  32'h3d1f2a5d /* (2, 6, 4) */,
  32'h3d7c66bd /* (30, 2, 4) */,
  32'h3d1f2a5d /* (26, 2, 4) */,
  32'h3d19eb69 /* (22, 2, 4) */,
  32'h3d3430e1 /* (18, 2, 4) */,
  32'h3d3430e1 /* (14, 2, 4) */,
  32'h3d19eb69 /* (10, 2, 4) */,
  32'h3d1f2a5d /* (6, 2, 4) */,
  32'h3d7c66bd /* (2, 2, 4) */,
  32'h3e1befb2 /* (30, 30, 0) */,
  32'h3d378ea1 /* (26, 30, 0) */,
  32'h3d124c17 /* (22, 30, 0) */,
  32'h3d204e75 /* (18, 30, 0) */,
  32'h3d204e75 /* (14, 30, 0) */,
  32'h3d124c17 /* (10, 30, 0) */,
  32'h3d378ea1 /* (6, 30, 0) */,
  32'h3e1befb2 /* (2, 30, 0) */,
  32'h3d378ea1 /* (30, 26, 0) */,
  32'h3d160c85 /* (26, 26, 0) */,
  32'h3d249cf9 /* (22, 26, 0) */,
  32'h3d4b578e /* (18, 26, 0) */,
  32'h3d4b578e /* (14, 26, 0) */,
  32'h3d249cf9 /* (10, 26, 0) */,
  32'h3d160c85 /* (6, 26, 0) */,
  32'h3d378ea1 /* (2, 26, 0) */,
  32'h3d124c17 /* (30, 22, 0) */,
  32'h3d249cf9 /* (26, 22, 0) */,
  32'h3d67f590 /* (22, 22, 0) */,
  32'h3da521d3 /* (18, 22, 0) */,
  32'h3da521d3 /* (14, 22, 0) */,
  32'h3d67f590 /* (10, 22, 0) */,
  32'h3d249cf9 /* (6, 22, 0) */,
  32'h3d124c17 /* (2, 22, 0) */,
  32'h3d204e75 /* (30, 18, 0) */,
  32'h3d4b578e /* (26, 18, 0) */,
  32'h3da521d3 /* (22, 18, 0) */,
  32'h3e036079 /* (18, 18, 0) */,
  32'h3e036079 /* (14, 18, 0) */,
  32'h3da521d3 /* (10, 18, 0) */,
  32'h3d4b578e /* (6, 18, 0) */,
  32'h3d204e75 /* (2, 18, 0) */,
  32'h3d204e75 /* (30, 14, 0) */,
  32'h3d4b578e /* (26, 14, 0) */,
  32'h3da521d3 /* (22, 14, 0) */,
  32'h3e036079 /* (18, 14, 0) */,
  32'h3e036079 /* (14, 14, 0) */,
  32'h3da521d3 /* (10, 14, 0) */,
  32'h3d4b578e /* (6, 14, 0) */,
  32'h3d204e75 /* (2, 14, 0) */,
  32'h3d124c17 /* (30, 10, 0) */,
  32'h3d249cf9 /* (26, 10, 0) */,
  32'h3d67f590 /* (22, 10, 0) */,
  32'h3da521d3 /* (18, 10, 0) */,
  32'h3da521d3 /* (14, 10, 0) */,
  32'h3d67f590 /* (10, 10, 0) */,
  32'h3d249cf9 /* (6, 10, 0) */,
  32'h3d124c17 /* (2, 10, 0) */,
  32'h3d378ea1 /* (30, 6, 0) */,
  32'h3d160c85 /* (26, 6, 0) */,
  32'h3d249cf9 /* (22, 6, 0) */,
  32'h3d4b578e /* (18, 6, 0) */,
  32'h3d4b578e /* (14, 6, 0) */,
  32'h3d249cf9 /* (10, 6, 0) */,
  32'h3d160c85 /* (6, 6, 0) */,
  32'h3d378ea1 /* (2, 6, 0) */,
  32'h3e1befb2 /* (30, 2, 0) */,
  32'h3d378ea1 /* (26, 2, 0) */,
  32'h3d124c17 /* (22, 2, 0) */,
  32'h3d204e75 /* (18, 2, 0) */,
  32'h3d204e75 /* (14, 2, 0) */,
  32'h3d124c17 /* (10, 2, 0) */,
  32'h3d378ea1 /* (6, 2, 0) */,
  32'h3e1befb2 /* (2, 2, 0) */,
  32'h3d5defd3 /* (29, 30, 28) */,
  32'h3d16c6a3 /* (25, 30, 28) */,
  32'h3d21c128 /* (21, 30, 28) */,
  32'h3d2d6bba /* (17, 30, 28) */,
  32'h3d3217f4 /* (13, 30, 28) */,
  32'h3d14de35 /* (9, 30, 28) */,
  32'h3d2d8e0e /* (5, 30, 28) */,
  32'h3d8b1391 /* (1, 30, 28) */,
  32'h3d1b3fff /* (29, 26, 28) */,
  32'h3d17902e /* (25, 26, 28) */,
  32'h3d41fb9f /* (21, 26, 28) */,
  32'h3d61b1de /* (17, 26, 28) */,
  32'h3d601ae9 /* (13, 26, 28) */,
  32'h3d2657dd /* (9, 26, 28) */,
  32'h3d153e19 /* (5, 26, 28) */,
  32'h3d222a9c /* (1, 26, 28) */,
  32'h3d1cff11 /* (29, 22, 28) */,
  32'h3d404057 /* (25, 22, 28) */,
  32'h3d92b699 /* (21, 22, 28) */,
  32'h3dbdf4f8 /* (17, 22, 28) */,
  32'h3db40e50 /* (13, 22, 28) */,
  32'h3d68b7a2 /* (9, 22, 28) */,
  32'h3d28e3b2 /* (5, 22, 28) */,
  32'h3d1839e3 /* (1, 22, 28) */,
  32'h3d3b1e93 /* (29, 18, 28) */,
  32'h3d800deb /* (25, 18, 28) */,
  32'h3ddc0819 /* (21, 18, 28) */,
  32'h3e1c2ca1 /* (17, 18, 28) */,
  32'h3e0de89e /* (13, 18, 28) */,
  32'h3da4db8a /* (9, 18, 28) */,
  32'h3d53bb31 /* (5, 18, 28) */,
  32'h3d303352 /* (1, 18, 28) */,
  32'h3d3b1e93 /* (29, 14, 28) */,
  32'h3d800deb /* (25, 14, 28) */,
  32'h3ddc0819 /* (21, 14, 28) */,
  32'h3e1c2ca1 /* (17, 14, 28) */,
  32'h3e0de89e /* (13, 14, 28) */,
  32'h3da4db8a /* (9, 14, 28) */,
  32'h3d53bb31 /* (5, 14, 28) */,
  32'h3d303352 /* (1, 14, 28) */,
  32'h3d1cff11 /* (29, 10, 28) */,
  32'h3d404057 /* (25, 10, 28) */,
  32'h3d92b699 /* (21, 10, 28) */,
  32'h3dbdf4f8 /* (17, 10, 28) */,
  32'h3db40e50 /* (13, 10, 28) */,
  32'h3d68b7a2 /* (9, 10, 28) */,
  32'h3d28e3b2 /* (5, 10, 28) */,
  32'h3d1839e3 /* (1, 10, 28) */,
  32'h3d1b3fff /* (29, 6, 28) */,
  32'h3d17902e /* (25, 6, 28) */,
  32'h3d41fb9f /* (21, 6, 28) */,
  32'h3d61b1de /* (17, 6, 28) */,
  32'h3d601ae9 /* (13, 6, 28) */,
  32'h3d2657dd /* (9, 6, 28) */,
  32'h3d153e19 /* (5, 6, 28) */,
  32'h3d222a9c /* (1, 6, 28) */,
  32'h3d5defd3 /* (29, 2, 28) */,
  32'h3d16c6a3 /* (25, 2, 28) */,
  32'h3d21c128 /* (21, 2, 28) */,
  32'h3d2d6bba /* (17, 2, 28) */,
  32'h3d3217f4 /* (13, 2, 28) */,
  32'h3d14de35 /* (9, 2, 28) */,
  32'h3d2d8e0e /* (5, 2, 28) */,
  32'h3d8b1391 /* (1, 2, 28) */,
  32'h3d13e9f7 /* (29, 30, 24) */,
  32'h3d1d59b0 /* (25, 30, 24) */,
  32'h3d558b1c /* (21, 30, 24) */,
  32'h3d804df8 /* (17, 30, 24) */,
  32'h3d7b52f8 /* (13, 30, 24) */,
  32'h3d3291f6 /* (9, 30, 24) */,
  32'h3d149b5c /* (5, 30, 24) */,
  32'h3d15ce12 /* (1, 30, 24) */,
  32'h3d19bf4b /* (29, 26, 24) */,
  32'h3d35cd98 /* (25, 26, 24) */,
  32'h3d865b59 /* (21, 26, 24) */,
  32'h3daa3349 /* (17, 26, 24) */,
  32'h3da2e7a9 /* (13, 26, 24) */,
  32'h3d584c0c /* (9, 26, 24) */,
  32'h3d22af34 /* (5, 26, 24) */,
  32'h3d169650 /* (1, 26, 24) */,
  32'h3d48bc7e /* (29, 22, 24) */,
  32'h3d83c517 /* (25, 22, 24) */,
  32'h3dd7e578 /* (21, 22, 24) */,
  32'h3e135573 /* (17, 22, 24) */,
  32'h3e085939 /* (13, 22, 24) */,
  32'h3da590e9 /* (9, 22, 24) */,
  32'h3d5ef675 /* (5, 22, 24) */,
  32'h3d3f0366 /* (1, 22, 24) */,
  32'h3d880501 /* (29, 18, 24) */,
  32'h3dbf672f /* (25, 18, 24) */,
  32'h3e2a27e4 /* (21, 18, 24) */,
  32'h3e79034c /* (17, 18, 24) */,
  32'h3e5f05ce /* (13, 18, 24) */,
  32'h3dfaaa60 /* (9, 18, 24) */,
  32'h3d9bc970 /* (5, 18, 24) */,
  32'h3d7e759f /* (1, 18, 24) */,
  32'h3d880501 /* (29, 14, 24) */,
  32'h3dbf672f /* (25, 14, 24) */,
  32'h3e2a27e4 /* (21, 14, 24) */,
  32'h3e79034c /* (17, 14, 24) */,
  32'h3e5f05ce /* (13, 14, 24) */,
  32'h3dfaaa60 /* (9, 14, 24) */,
  32'h3d9bc970 /* (5, 14, 24) */,
  32'h3d7e759f /* (1, 14, 24) */,
  32'h3d48bc7e /* (29, 10, 24) */,
  32'h3d83c517 /* (25, 10, 24) */,
  32'h3dd7e578 /* (21, 10, 24) */,
  32'h3e135573 /* (17, 10, 24) */,
  32'h3e085939 /* (13, 10, 24) */,
  32'h3da590e9 /* (9, 10, 24) */,
  32'h3d5ef675 /* (5, 10, 24) */,
  32'h3d3f0366 /* (1, 10, 24) */,
  32'h3d19bf4b /* (29, 6, 24) */,
  32'h3d35cd98 /* (25, 6, 24) */,
  32'h3d865b59 /* (21, 6, 24) */,
  32'h3daa3349 /* (17, 6, 24) */,
  32'h3da2e7a9 /* (13, 6, 24) */,
  32'h3d584c0c /* (9, 6, 24) */,
  32'h3d22af34 /* (5, 6, 24) */,
  32'h3d169650 /* (1, 6, 24) */,
  32'h3d13e9f7 /* (29, 2, 24) */,
  32'h3d1d59b0 /* (25, 2, 24) */,
  32'h3d558b1c /* (21, 2, 24) */,
  32'h3d804df8 /* (17, 2, 24) */,
  32'h3d7b52f8 /* (13, 2, 24) */,
  32'h3d3291f6 /* (9, 2, 24) */,
  32'h3d149b5c /* (5, 2, 24) */,
  32'h3d15ce12 /* (1, 2, 24) */,
  32'h3d23d587 /* (29, 30, 20) */,
  32'h3d530d8e /* (25, 30, 20) */,
  32'h3da96c08 /* (21, 30, 20) */,
  32'h3de39dff /* (17, 30, 20) */,
  32'h3dd42d31 /* (13, 30, 20) */,
  32'h3d833332 /* (9, 30, 20) */,
  32'h3d346b02 /* (5, 30, 20) */,
  32'h3d1cac31 /* (1, 30, 20) */,
  32'h3d48406d /* (29, 26, 20) */,
  32'h3d859348 /* (25, 26, 20) */,
  32'h3ddec971 /* (21, 26, 20) */,
  32'h3e1a3a56 /* (17, 26, 20) */,
  32'h3e0dc95f /* (13, 26, 20) */,
  32'h3da96159 /* (9, 26, 20) */,
  32'h3d6007ad /* (5, 26, 20) */,
  32'h3d3dc5f0 /* (1, 26, 20) */,
  32'h3d9aff71 /* (29, 22, 20) */,
  32'h3dd85675 /* (25, 22, 20) */,
  32'h3e3e5baf /* (21, 22, 20) */,
  32'h3e89fde5 /* (17, 22, 20) */,
  32'h3e7848b5 /* (13, 22, 20) */,
  32'h3e0cf021 /* (9, 22, 20) */,
  32'h3db0e528 /* (5, 22, 20) */,
  32'h3d91435f /* (1, 22, 20) */,
  32'h3decc5e8 /* (29, 18, 20) */,
  32'h3e2baf50 /* (25, 18, 20) */,
  32'h3e9ecc49 /* (21, 18, 20) */,
  32'h3ef15f91 /* (17, 18, 20) */,
  32'h3ed441df /* (13, 18, 20) */,
  32'h3e654448 /* (9, 18, 20) */,
  32'h3e095be4 /* (5, 18, 20) */,
  32'h3ddbed5a /* (1, 18, 20) */,
  32'h3decc5e8 /* (29, 14, 20) */,
  32'h3e2baf50 /* (25, 14, 20) */,
  32'h3e9ecc49 /* (21, 14, 20) */,
  32'h3ef15f91 /* (17, 14, 20) */,
  32'h3ed441df /* (13, 14, 20) */,
  32'h3e654448 /* (9, 14, 20) */,
  32'h3e095be4 /* (5, 14, 20) */,
  32'h3ddbed5a /* (1, 14, 20) */,
  32'h3d9aff71 /* (29, 10, 20) */,
  32'h3dd85675 /* (25, 10, 20) */,
  32'h3e3e5baf /* (21, 10, 20) */,
  32'h3e89fde5 /* (17, 10, 20) */,
  32'h3e7848b5 /* (13, 10, 20) */,
  32'h3e0cf021 /* (9, 10, 20) */,
  32'h3db0e528 /* (5, 10, 20) */,
  32'h3d91435f /* (1, 10, 20) */,
  32'h3d48406d /* (29, 6, 20) */,
  32'h3d859348 /* (25, 6, 20) */,
  32'h3ddec971 /* (21, 6, 20) */,
  32'h3e1a3a56 /* (17, 6, 20) */,
  32'h3e0dc95f /* (13, 6, 20) */,
  32'h3da96159 /* (9, 6, 20) */,
  32'h3d6007ad /* (5, 6, 20) */,
  32'h3d3dc5f0 /* (1, 6, 20) */,
  32'h3d23d587 /* (29, 2, 20) */,
  32'h3d530d8e /* (25, 2, 20) */,
  32'h3da96c08 /* (21, 2, 20) */,
  32'h3de39dff /* (17, 2, 20) */,
  32'h3dd42d31 /* (13, 2, 20) */,
  32'h3d833332 /* (9, 2, 20) */,
  32'h3d346b02 /* (5, 2, 20) */,
  32'h3d1cac31 /* (1, 2, 20) */,
  32'h3d13661d /* (29, 30, 16) */,
  32'h3d4f6a6e /* (25, 30, 16) */,
  32'h3db86416 /* (21, 30, 16) */,
  32'h3e06ec2e /* (17, 30, 16) */,
  32'h3df1ae3d /* (13, 30, 16) */,
  32'h3d87d16b /* (9, 30, 16) */,
  32'h3d28d1e5 /* (5, 30, 16) */,
  32'h3d09dfab /* (1, 30, 16) */,
  32'h3d41d3ae /* (29, 26, 16) */,
  32'h3d8a46e7 /* (25, 26, 16) */,
  32'h3dfa4afe /* (21, 26, 16) */,
  32'h3e3a3d1a /* (17, 26, 16) */,
  32'h3e2576a9 /* (13, 26, 16) */,
  32'h3db6b309 /* (9, 26, 16) */,
  32'h3d5f53fb /* (5, 26, 16) */,
  32'h3d34b66a /* (1, 26, 16) */,
  32'h3da59d10 /* (29, 22, 16) */,
  32'h3df142da /* (25, 22, 16) */,
  32'h3e60898b /* (21, 22, 16) */,
  32'h3eabb572 /* (17, 22, 16) */,
  32'h3e968a40 /* (13, 22, 16) */,
  32'h3e21930d /* (9, 22, 16) */,
  32'h3dc0863e /* (5, 22, 16) */,
  32'h3d99ac24 /* (1, 22, 16) */,
  32'h3e0a27e7 /* (29, 18, 16) */,
  32'h3e4d7ce8 /* (25, 18, 16) */,
  32'h3ec4f0a1 /* (21, 18, 16) */,
  32'h3f1b42bd /* (17, 18, 16) */,
  32'h3f06176f /* (13, 18, 16) */,
  32'h3e8b9344 /* (9, 18, 16) */,
  32'h3e2205a1 /* (5, 18, 16) */,
  32'h3dff32bb /* (1, 18, 16) */,
  32'h3e0a27e7 /* (29, 14, 16) */,
  32'h3e4d7ce8 /* (25, 14, 16) */,
  32'h3ec4f0a1 /* (21, 14, 16) */,
  32'h3f1b42bd /* (17, 14, 16) */,
  32'h3f06176f /* (13, 14, 16) */,
  32'h3e8b9344 /* (9, 14, 16) */,
  32'h3e2205a1 /* (5, 14, 16) */,
  32'h3dff32bb /* (1, 14, 16) */,
  32'h3da59d10 /* (29, 10, 16) */,
  32'h3df142da /* (25, 10, 16) */,
  32'h3e60898b /* (21, 10, 16) */,
  32'h3eabb572 /* (17, 10, 16) */,
  32'h3e968a40 /* (13, 10, 16) */,
  32'h3e21930d /* (9, 10, 16) */,
  32'h3dc0863e /* (5, 10, 16) */,
  32'h3d99ac24 /* (1, 10, 16) */,
  32'h3d41d3ae /* (29, 6, 16) */,
  32'h3d8a46e7 /* (25, 6, 16) */,
  32'h3dfa4afe /* (21, 6, 16) */,
  32'h3e3a3d1a /* (17, 6, 16) */,
  32'h3e2576a9 /* (13, 6, 16) */,
  32'h3db6b309 /* (9, 6, 16) */,
  32'h3d5f53fb /* (5, 6, 16) */,
  32'h3d34b66a /* (1, 6, 16) */,
  32'h3d13661d /* (29, 2, 16) */,
  32'h3d4f6a6e /* (25, 2, 16) */,
  32'h3db86416 /* (21, 2, 16) */,
  32'h3e06ec2e /* (17, 2, 16) */,
  32'h3df1ae3d /* (13, 2, 16) */,
  32'h3d87d16b /* (9, 2, 16) */,
  32'h3d28d1e5 /* (5, 2, 16) */,
  32'h3d09dfab /* (1, 2, 16) */,
  32'h3d23d587 /* (29, 30, 12) */,
  32'h3d530d8e /* (25, 30, 12) */,
  32'h3da96c08 /* (21, 30, 12) */,
  32'h3de39dff /* (17, 30, 12) */,
  32'h3dd42d31 /* (13, 30, 12) */,
  32'h3d833332 /* (9, 30, 12) */,
  32'h3d346b02 /* (5, 30, 12) */,
  32'h3d1cac31 /* (1, 30, 12) */,
  32'h3d48406d /* (29, 26, 12) */,
  32'h3d859348 /* (25, 26, 12) */,
  32'h3ddec971 /* (21, 26, 12) */,
  32'h3e1a3a56 /* (17, 26, 12) */,
  32'h3e0dc95f /* (13, 26, 12) */,
  32'h3da96159 /* (9, 26, 12) */,
  32'h3d6007ad /* (5, 26, 12) */,
  32'h3d3dc5f0 /* (1, 26, 12) */,
  32'h3d9aff71 /* (29, 22, 12) */,
  32'h3dd85675 /* (25, 22, 12) */,
  32'h3e3e5baf /* (21, 22, 12) */,
  32'h3e89fde5 /* (17, 22, 12) */,
  32'h3e7848b5 /* (13, 22, 12) */,
  32'h3e0cf021 /* (9, 22, 12) */,
  32'h3db0e528 /* (5, 22, 12) */,
  32'h3d91435f /* (1, 22, 12) */,
  32'h3decc5e8 /* (29, 18, 12) */,
  32'h3e2baf50 /* (25, 18, 12) */,
  32'h3e9ecc49 /* (21, 18, 12) */,
  32'h3ef15f91 /* (17, 18, 12) */,
  32'h3ed441df /* (13, 18, 12) */,
  32'h3e654448 /* (9, 18, 12) */,
  32'h3e095be4 /* (5, 18, 12) */,
  32'h3ddbed5a /* (1, 18, 12) */,
  32'h3decc5e8 /* (29, 14, 12) */,
  32'h3e2baf50 /* (25, 14, 12) */,
  32'h3e9ecc49 /* (21, 14, 12) */,
  32'h3ef15f91 /* (17, 14, 12) */,
  32'h3ed441df /* (13, 14, 12) */,
  32'h3e654448 /* (9, 14, 12) */,
  32'h3e095be4 /* (5, 14, 12) */,
  32'h3ddbed5a /* (1, 14, 12) */,
  32'h3d9aff71 /* (29, 10, 12) */,
  32'h3dd85675 /* (25, 10, 12) */,
  32'h3e3e5baf /* (21, 10, 12) */,
  32'h3e89fde5 /* (17, 10, 12) */,
  32'h3e7848b5 /* (13, 10, 12) */,
  32'h3e0cf021 /* (9, 10, 12) */,
  32'h3db0e528 /* (5, 10, 12) */,
  32'h3d91435f /* (1, 10, 12) */,
  32'h3d48406d /* (29, 6, 12) */,
  32'h3d859348 /* (25, 6, 12) */,
  32'h3ddec971 /* (21, 6, 12) */,
  32'h3e1a3a56 /* (17, 6, 12) */,
  32'h3e0dc95f /* (13, 6, 12) */,
  32'h3da96159 /* (9, 6, 12) */,
  32'h3d6007ad /* (5, 6, 12) */,
  32'h3d3dc5f0 /* (1, 6, 12) */,
  32'h3d23d587 /* (29, 2, 12) */,
  32'h3d530d8e /* (25, 2, 12) */,
  32'h3da96c08 /* (21, 2, 12) */,
  32'h3de39dff /* (17, 2, 12) */,
  32'h3dd42d31 /* (13, 2, 12) */,
  32'h3d833332 /* (9, 2, 12) */,
  32'h3d346b02 /* (5, 2, 12) */,
  32'h3d1cac31 /* (1, 2, 12) */,
  32'h3d13e9f7 /* (29, 30, 8) */,
  32'h3d1d59b0 /* (25, 30, 8) */,
  32'h3d558b1c /* (21, 30, 8) */,
  32'h3d804df8 /* (17, 30, 8) */,
  32'h3d7b52f8 /* (13, 30, 8) */,
  32'h3d3291f6 /* (9, 30, 8) */,
  32'h3d149b5c /* (5, 30, 8) */,
  32'h3d15ce12 /* (1, 30, 8) */,
  32'h3d19bf4b /* (29, 26, 8) */,
  32'h3d35cd98 /* (25, 26, 8) */,
  32'h3d865b59 /* (21, 26, 8) */,
  32'h3daa3349 /* (17, 26, 8) */,
  32'h3da2e7a9 /* (13, 26, 8) */,
  32'h3d584c0c /* (9, 26, 8) */,
  32'h3d22af34 /* (5, 26, 8) */,
  32'h3d169650 /* (1, 26, 8) */,
  32'h3d48bc7e /* (29, 22, 8) */,
  32'h3d83c517 /* (25, 22, 8) */,
  32'h3dd7e578 /* (21, 22, 8) */,
  32'h3e135573 /* (17, 22, 8) */,
  32'h3e085939 /* (13, 22, 8) */,
  32'h3da590e9 /* (9, 22, 8) */,
  32'h3d5ef675 /* (5, 22, 8) */,
  32'h3d3f0366 /* (1, 22, 8) */,
  32'h3d880501 /* (29, 18, 8) */,
  32'h3dbf672f /* (25, 18, 8) */,
  32'h3e2a27e4 /* (21, 18, 8) */,
  32'h3e79034c /* (17, 18, 8) */,
  32'h3e5f05ce /* (13, 18, 8) */,
  32'h3dfaaa60 /* (9, 18, 8) */,
  32'h3d9bc970 /* (5, 18, 8) */,
  32'h3d7e759f /* (1, 18, 8) */,
  32'h3d880501 /* (29, 14, 8) */,
  32'h3dbf672f /* (25, 14, 8) */,
  32'h3e2a27e4 /* (21, 14, 8) */,
  32'h3e79034c /* (17, 14, 8) */,
  32'h3e5f05ce /* (13, 14, 8) */,
  32'h3dfaaa60 /* (9, 14, 8) */,
  32'h3d9bc970 /* (5, 14, 8) */,
  32'h3d7e759f /* (1, 14, 8) */,
  32'h3d48bc7e /* (29, 10, 8) */,
  32'h3d83c517 /* (25, 10, 8) */,
  32'h3dd7e578 /* (21, 10, 8) */,
  32'h3e135573 /* (17, 10, 8) */,
  32'h3e085939 /* (13, 10, 8) */,
  32'h3da590e9 /* (9, 10, 8) */,
  32'h3d5ef675 /* (5, 10, 8) */,
  32'h3d3f0366 /* (1, 10, 8) */,
  32'h3d19bf4b /* (29, 6, 8) */,
  32'h3d35cd98 /* (25, 6, 8) */,
  32'h3d865b59 /* (21, 6, 8) */,
  32'h3daa3349 /* (17, 6, 8) */,
  32'h3da2e7a9 /* (13, 6, 8) */,
  32'h3d584c0c /* (9, 6, 8) */,
  32'h3d22af34 /* (5, 6, 8) */,
  32'h3d169650 /* (1, 6, 8) */,
  32'h3d13e9f7 /* (29, 2, 8) */,
  32'h3d1d59b0 /* (25, 2, 8) */,
  32'h3d558b1c /* (21, 2, 8) */,
  32'h3d804df8 /* (17, 2, 8) */,
  32'h3d7b52f8 /* (13, 2, 8) */,
  32'h3d3291f6 /* (9, 2, 8) */,
  32'h3d149b5c /* (5, 2, 8) */,
  32'h3d15ce12 /* (1, 2, 8) */,
  32'h3d5defd3 /* (29, 30, 4) */,
  32'h3d16c6a3 /* (25, 30, 4) */,
  32'h3d21c128 /* (21, 30, 4) */,
  32'h3d2d6bba /* (17, 30, 4) */,
  32'h3d3217f4 /* (13, 30, 4) */,
  32'h3d14de35 /* (9, 30, 4) */,
  32'h3d2d8e0e /* (5, 30, 4) */,
  32'h3d8b1391 /* (1, 30, 4) */,
  32'h3d1b3fff /* (29, 26, 4) */,
  32'h3d17902e /* (25, 26, 4) */,
  32'h3d41fb9f /* (21, 26, 4) */,
  32'h3d61b1de /* (17, 26, 4) */,
  32'h3d601ae9 /* (13, 26, 4) */,
  32'h3d2657dd /* (9, 26, 4) */,
  32'h3d153e19 /* (5, 26, 4) */,
  32'h3d222a9c /* (1, 26, 4) */,
  32'h3d1cff11 /* (29, 22, 4) */,
  32'h3d404057 /* (25, 22, 4) */,
  32'h3d92b699 /* (21, 22, 4) */,
  32'h3dbdf4f8 /* (17, 22, 4) */,
  32'h3db40e50 /* (13, 22, 4) */,
  32'h3d68b7a2 /* (9, 22, 4) */,
  32'h3d28e3b2 /* (5, 22, 4) */,
  32'h3d1839e3 /* (1, 22, 4) */,
  32'h3d3b1e93 /* (29, 18, 4) */,
  32'h3d800deb /* (25, 18, 4) */,
  32'h3ddc0819 /* (21, 18, 4) */,
  32'h3e1c2ca1 /* (17, 18, 4) */,
  32'h3e0de89e /* (13, 18, 4) */,
  32'h3da4db8a /* (9, 18, 4) */,
  32'h3d53bb31 /* (5, 18, 4) */,
  32'h3d303352 /* (1, 18, 4) */,
  32'h3d3b1e93 /* (29, 14, 4) */,
  32'h3d800deb /* (25, 14, 4) */,
  32'h3ddc0819 /* (21, 14, 4) */,
  32'h3e1c2ca1 /* (17, 14, 4) */,
  32'h3e0de89e /* (13, 14, 4) */,
  32'h3da4db8a /* (9, 14, 4) */,
  32'h3d53bb31 /* (5, 14, 4) */,
  32'h3d303352 /* (1, 14, 4) */,
  32'h3d1cff11 /* (29, 10, 4) */,
  32'h3d404057 /* (25, 10, 4) */,
  32'h3d92b699 /* (21, 10, 4) */,
  32'h3dbdf4f8 /* (17, 10, 4) */,
  32'h3db40e50 /* (13, 10, 4) */,
  32'h3d68b7a2 /* (9, 10, 4) */,
  32'h3d28e3b2 /* (5, 10, 4) */,
  32'h3d1839e3 /* (1, 10, 4) */,
  32'h3d1b3fff /* (29, 6, 4) */,
  32'h3d17902e /* (25, 6, 4) */,
  32'h3d41fb9f /* (21, 6, 4) */,
  32'h3d61b1de /* (17, 6, 4) */,
  32'h3d601ae9 /* (13, 6, 4) */,
  32'h3d2657dd /* (9, 6, 4) */,
  32'h3d153e19 /* (5, 6, 4) */,
  32'h3d222a9c /* (1, 6, 4) */,
  32'h3d5defd3 /* (29, 2, 4) */,
  32'h3d16c6a3 /* (25, 2, 4) */,
  32'h3d21c128 /* (21, 2, 4) */,
  32'h3d2d6bba /* (17, 2, 4) */,
  32'h3d3217f4 /* (13, 2, 4) */,
  32'h3d14de35 /* (9, 2, 4) */,
  32'h3d2d8e0e /* (5, 2, 4) */,
  32'h3d8b1391 /* (1, 2, 4) */,
  32'h3dcbea25 /* (29, 30, 0) */,
  32'h3d21b235 /* (25, 30, 0) */,
  32'h3d164ce1 /* (21, 30, 0) */,
  32'h3d18d610 /* (17, 30, 0) */,
  32'h3d2045b1 /* (13, 30, 0) */,
  32'h3d11b684 /* (9, 30, 0) */,
  32'h3d5dd7d1 /* (5, 30, 0) */,
  32'h3e709592 /* (1, 30, 0) */,
  32'h3d2d5b95 /* (29, 26, 0) */,
  32'h3d1459dd /* (25, 26, 0) */,
  32'h3d3013e2 /* (21, 26, 0) */,
  32'h3d455011 /* (17, 26, 0) */,
  32'h3d4703b2 /* (13, 26, 0) */,
  32'h3d1bc36a /* (9, 26, 0) */,
  32'h3d1b2f33 /* (5, 26, 0) */,
  32'h3d3f59b8 /* (1, 26, 0) */,
  32'h3d144f19 /* (29, 22, 0) */,
  32'h3d2f5f5a /* (25, 22, 0) */,
  32'h3d819abc /* (21, 22, 0) */,
  32'h3da42e1b /* (17, 22, 0) */,
  32'h3d9d248b /* (13, 22, 0) */,
  32'h3d50a575 /* (9, 22, 0) */,
  32'h3d1cee15 /* (5, 22, 0) */,
  32'h3d1142bb /* (1, 22, 0) */,
  32'h3d262b6e /* (29, 18, 0) */,
  32'h3d60bf24 /* (25, 18, 0) */,
  32'h3dbe661f /* (21, 18, 0) */,
  32'h3e05899d /* (17, 18, 0) */,
  32'h3df40add /* (13, 18, 0) */,
  32'h3d8fa52c /* (9, 18, 0) */,
  32'h3d3b0a55 /* (5, 18, 0) */,
  32'h3d1ceee6 /* (1, 18, 0) */,
  32'h3d262b6e /* (29, 14, 0) */,
  32'h3d60bf24 /* (25, 14, 0) */,
  32'h3dbe661f /* (21, 14, 0) */,
  32'h3e05899d /* (17, 14, 0) */,
  32'h3df40add /* (13, 14, 0) */,
  32'h3d8fa52c /* (9, 14, 0) */,
  32'h3d3b0a55 /* (5, 14, 0) */,
  32'h3d1ceee6 /* (1, 14, 0) */,
  32'h3d144f19 /* (29, 10, 0) */,
  32'h3d2f5f5a /* (25, 10, 0) */,
  32'h3d819abc /* (21, 10, 0) */,
  32'h3da42e1b /* (17, 10, 0) */,
  32'h3d9d248b /* (13, 10, 0) */,
  32'h3d50a575 /* (9, 10, 0) */,
  32'h3d1cee15 /* (5, 10, 0) */,
  32'h3d1142bb /* (1, 10, 0) */,
  32'h3d2d5b95 /* (29, 6, 0) */,
  32'h3d1459dd /* (25, 6, 0) */,
  32'h3d3013e2 /* (21, 6, 0) */,
  32'h3d455011 /* (17, 6, 0) */,
  32'h3d4703b2 /* (13, 6, 0) */,
  32'h3d1bc36a /* (9, 6, 0) */,
  32'h3d1b2f33 /* (5, 6, 0) */,
  32'h3d3f59b8 /* (1, 6, 0) */,
  32'h3dcbea25 /* (29, 2, 0) */,
  32'h3d21b235 /* (25, 2, 0) */,
  32'h3d164ce1 /* (21, 2, 0) */,
  32'h3d18d610 /* (17, 2, 0) */,
  32'h3d2045b1 /* (13, 2, 0) */,
  32'h3d11b684 /* (9, 2, 0) */,
  32'h3d5dd7d1 /* (5, 2, 0) */,
  32'h3e709592 /* (1, 2, 0) */,
  32'h3d429928 /* (28, 30, 28) */,
  32'h3d139519 /* (24, 30, 28) */,
  32'h3d2ab74a /* (20, 30, 28) */,
  32'h3d1c5e8a /* (16, 30, 28) */,
  32'h3d2ab74a /* (12, 30, 28) */,
  32'h3d139519 /* (8, 30, 28) */,
  32'h3d429928 /* (4, 30, 28) */,
  32'h3d90451b /* (0, 30, 28) */,
  32'h3d1796af /* (28, 26, 28) */,
  32'h3d1d3fef /* (24, 26, 28) */,
  32'h3d522ea6 /* (20, 26, 28) */,
  32'h3d4e2dc2 /* (16, 26, 28) */,
  32'h3d522ea6 /* (12, 26, 28) */,
  32'h3d1d3fef /* (8, 26, 28) */,
  32'h3d1796af /* (4, 26, 28) */,
  32'h3d234ae8 /* (0, 26, 28) */,
  32'h3d21d2a4 /* (28, 22, 28) */,
  32'h3d51ff4c /* (24, 22, 28) */,
  32'h3da42ada /* (20, 22, 28) */,
  32'h3db0df4f /* (16, 22, 28) */,
  32'h3da42ada /* (12, 22, 28) */,
  32'h3d51ff4c /* (8, 22, 28) */,
  32'h3d21d2a4 /* (4, 22, 28) */,
  32'h3d17b006 /* (0, 22, 28) */,
  32'h3d456b70 /* (28, 18, 28) */,
  32'h3d904c26 /* (24, 18, 28) */,
  32'h3dfca6c8 /* (20, 18, 28) */,
  32'h3e1420e4 /* (16, 18, 28) */,
  32'h3dfca6c8 /* (12, 18, 28) */,
  32'h3d904c26 /* (8, 18, 28) */,
  32'h3d456b70 /* (4, 18, 28) */,
  32'h3d2ee5c8 /* (0, 18, 28) */,
  32'h3d456b70 /* (28, 14, 28) */,
  32'h3d904c26 /* (24, 14, 28) */,
  32'h3dfca6c8 /* (20, 14, 28) */,
  32'h3e1420e4 /* (16, 14, 28) */,
  32'h3dfca6c8 /* (12, 14, 28) */,
  32'h3d904c26 /* (8, 14, 28) */,
  32'h3d456b70 /* (4, 14, 28) */,
  32'h3d2ee5c8 /* (0, 14, 28) */,
  32'h3d21d2a4 /* (28, 10, 28) */,
  32'h3d51ff4c /* (24, 10, 28) */,
  32'h3da42ada /* (20, 10, 28) */,
  32'h3db0df4f /* (16, 10, 28) */,
  32'h3da42ada /* (12, 10, 28) */,
  32'h3d51ff4c /* (8, 10, 28) */,
  32'h3d21d2a4 /* (4, 10, 28) */,
  32'h3d17b006 /* (0, 10, 28) */,
  32'h3d1796af /* (28, 6, 28) */,
  32'h3d1d3fef /* (24, 6, 28) */,
  32'h3d522ea6 /* (20, 6, 28) */,
  32'h3d4e2dc2 /* (16, 6, 28) */,
  32'h3d522ea6 /* (12, 6, 28) */,
  32'h3d1d3fef /* (8, 6, 28) */,
  32'h3d1796af /* (4, 6, 28) */,
  32'h3d234ae8 /* (0, 6, 28) */,
  32'h3d429928 /* (28, 2, 28) */,
  32'h3d139519 /* (24, 2, 28) */,
  32'h3d2ab74a /* (20, 2, 28) */,
  32'h3d1c5e8a /* (16, 2, 28) */,
  32'h3d2ab74a /* (12, 2, 28) */,
  32'h3d139519 /* (8, 2, 28) */,
  32'h3d429928 /* (4, 2, 28) */,
  32'h3d90451b /* (0, 2, 28) */,
  32'h3d139519 /* (28, 30, 24) */,
  32'h3d263161 /* (24, 30, 24) */,
  32'h3d69b2a3 /* (20, 30, 24) */,
  32'h3d6bb726 /* (16, 30, 24) */,
  32'h3d69b2a3 /* (12, 30, 24) */,
  32'h3d263161 /* (8, 30, 24) */,
  32'h3d139519 /* (4, 30, 24) */,
  32'h3d162cf4 /* (0, 30, 24) */,
  32'h3d1d3fef /* (28, 26, 24) */,
  32'h3d44d2c5 /* (24, 26, 24) */,
  32'h3d95625b /* (20, 26, 24) */,
  32'h3d9dd43f /* (16, 26, 24) */,
  32'h3d95625b /* (12, 26, 24) */,
  32'h3d44d2c5 /* (8, 26, 24) */,
  32'h3d1d3fef /* (4, 26, 24) */,
  32'h3d164277 /* (0, 26, 24) */,
  32'h3d51ff4c /* (28, 22, 24) */,
  32'h3d92b00e /* (24, 22, 24) */,
  32'h3df53c17 /* (20, 22, 24) */,
  32'h3e0a9c46 /* (16, 22, 24) */,
  32'h3df53c17 /* (12, 22, 24) */,
  32'h3d92b00e /* (8, 22, 24) */,
  32'h3d51ff4c /* (4, 22, 24) */,
  32'h3d3ddc84 /* (0, 22, 24) */,
  32'h3d904c26 /* (28, 18, 24) */,
  32'h3dd9849b /* (24, 18, 24) */,
  32'h3e44fc23 /* (20, 18, 24) */,
  32'h3e6dbe20 /* (16, 18, 24) */,
  32'h3e44fc23 /* (12, 18, 24) */,
  32'h3dd9849b /* (8, 18, 24) */,
  32'h3d904c26 /* (4, 18, 24) */,
  32'h3d7c5be6 /* (0, 18, 24) */,
  32'h3d904c26 /* (28, 14, 24) */,
  32'h3dd9849b /* (24, 14, 24) */,
  32'h3e44fc23 /* (20, 14, 24) */,
  32'h3e6dbe20 /* (16, 14, 24) */,
  32'h3e44fc23 /* (12, 14, 24) */,
  32'h3dd9849b /* (8, 14, 24) */,
  32'h3d904c26 /* (4, 14, 24) */,
  32'h3d7c5be6 /* (0, 14, 24) */,
  32'h3d51ff4c /* (28, 10, 24) */,
  32'h3d92b00e /* (24, 10, 24) */,
  32'h3df53c17 /* (20, 10, 24) */,
  32'h3e0a9c46 /* (16, 10, 24) */,
  32'h3df53c17 /* (12, 10, 24) */,
  32'h3d92b00e /* (8, 10, 24) */,
  32'h3d51ff4c /* (4, 10, 24) */,
  32'h3d3ddc84 /* (0, 10, 24) */,
  32'h3d1d3fef /* (28, 6, 24) */,
  32'h3d44d2c5 /* (24, 6, 24) */,
  32'h3d95625b /* (20, 6, 24) */,
  32'h3d9dd43f /* (16, 6, 24) */,
  32'h3d95625b /* (12, 6, 24) */,
  32'h3d44d2c5 /* (8, 6, 24) */,
  32'h3d1d3fef /* (4, 6, 24) */,
  32'h3d164277 /* (0, 6, 24) */,
  32'h3d139519 /* (28, 2, 24) */,
  32'h3d263161 /* (24, 2, 24) */,
  32'h3d69b2a3 /* (20, 2, 24) */,
  32'h3d6bb726 /* (16, 2, 24) */,
  32'h3d69b2a3 /* (12, 2, 24) */,
  32'h3d263161 /* (8, 2, 24) */,
  32'h3d139519 /* (4, 2, 24) */,
  32'h3d162cf4 /* (0, 2, 24) */,
  32'h3d2ab74a /* (28, 30, 20) */,
  32'h3d69b2a3 /* (24, 30, 20) */,
  32'h3dbf980c /* (20, 30, 20) */,
  32'h3dd576ed /* (16, 30, 20) */,
  32'h3dbf980c /* (12, 30, 20) */,
  32'h3d69b2a3 /* (8, 30, 20) */,
  32'h3d2ab74a /* (4, 30, 20) */,
  32'h3d1bd472 /* (0, 30, 20) */,
  32'h3d522ea6 /* (28, 26, 20) */,
  32'h3d95625b /* (24, 26, 20) */,
  32'h3dfe11f4 /* (20, 26, 20) */,
  32'h3e11854b /* (16, 26, 20) */,
  32'h3dfe11f4 /* (12, 26, 20) */,
  32'h3d95625b /* (8, 26, 20) */,
  32'h3d522ea6 /* (4, 26, 20) */,
  32'h3d3c86f4 /* (0, 26, 20) */,
  32'h3da42ada /* (28, 22, 20) */,
  32'h3df53c17 /* (24, 22, 20) */,
  32'h3e5bd2f1 /* (20, 22, 20) */,
  32'h3e837a14 /* (16, 22, 20) */,
  32'h3e5bd2f1 /* (12, 22, 20) */,
  32'h3df53c17 /* (8, 22, 20) */,
  32'h3da42ada /* (4, 22, 20) */,
  32'h3d9019ab /* (0, 22, 20) */,
  32'h3dfca6c8 /* (28, 18, 20) */,
  32'h3e44fc23 /* (24, 18, 20) */,
  32'h3eb9abaa /* (20, 18, 20) */,
  32'h3ee86d0e /* (16, 18, 20) */,
  32'h3eb9abaa /* (12, 18, 20) */,
  32'h3e44fc23 /* (8, 18, 20) */,
  32'h3dfca6c8 /* (4, 18, 20) */,
  32'h3dd9ea44 /* (0, 18, 20) */,
  32'h3dfca6c8 /* (28, 14, 20) */,
  32'h3e44fc23 /* (24, 14, 20) */,
  32'h3eb9abaa /* (20, 14, 20) */,
  32'h3ee86d0e /* (16, 14, 20) */,
  32'h3eb9abaa /* (12, 14, 20) */,
  32'h3e44fc23 /* (8, 14, 20) */,
  32'h3dfca6c8 /* (4, 14, 20) */,
  32'h3dd9ea44 /* (0, 14, 20) */,
  32'h3da42ada /* (28, 10, 20) */,
  32'h3df53c17 /* (24, 10, 20) */,
  32'h3e5bd2f1 /* (20, 10, 20) */,
  32'h3e837a14 /* (16, 10, 20) */,
  32'h3e5bd2f1 /* (12, 10, 20) */,
  32'h3df53c17 /* (8, 10, 20) */,
  32'h3da42ada /* (4, 10, 20) */,
  32'h3d9019ab /* (0, 10, 20) */,
  32'h3d522ea6 /* (28, 6, 20) */,
  32'h3d95625b /* (24, 6, 20) */,
  32'h3dfe11f4 /* (20, 6, 20) */,
  32'h3e11854b /* (16, 6, 20) */,
  32'h3dfe11f4 /* (12, 6, 20) */,
  32'h3d95625b /* (8, 6, 20) */,
  32'h3d522ea6 /* (4, 6, 20) */,
  32'h3d3c86f4 /* (0, 6, 20) */,
  32'h3d2ab74a /* (28, 2, 20) */,
  32'h3d69b2a3 /* (24, 2, 20) */,
  32'h3dbf980c /* (20, 2, 20) */,
  32'h3dd576ed /* (16, 2, 20) */,
  32'h3dbf980c /* (12, 2, 20) */,
  32'h3d69b2a3 /* (8, 2, 20) */,
  32'h3d2ab74a /* (4, 2, 20) */,
  32'h3d1bd472 /* (0, 2, 20) */,
  32'h3d1c5e8a /* (28, 30, 16) */,
  32'h3d6bb726 /* (24, 30, 16) */,
  32'h3dd576ed /* (20, 30, 16) */,
  32'h3e00d0e8 /* (16, 30, 16) */,
  32'h3dd576ed /* (12, 30, 16) */,
  32'h3d6bb726 /* (8, 30, 16) */,
  32'h3d1c5e8a /* (4, 30, 16) */,
  32'h3d08bc50 /* (0, 30, 16) */,
  32'h3d4e2dc2 /* (28, 26, 16) */,
  32'h3d9dd43f /* (24, 26, 16) */,
  32'h3e11854b /* (20, 26, 16) */,
  32'h3e327927 /* (16, 26, 16) */,
  32'h3e11854b /* (12, 26, 16) */,
  32'h3d9dd43f /* (8, 26, 16) */,
  32'h3d4e2dc2 /* (4, 26, 16) */,
  32'h3d332545 /* (0, 26, 16) */,
  32'h3db0df4f /* (28, 22, 16) */,
  32'h3e0a9c46 /* (24, 22, 16) */,
  32'h3e837a14 /* (20, 22, 16) */,
  32'h3ea594bb /* (16, 22, 16) */,
  32'h3e837a14 /* (12, 22, 16) */,
  32'h3e0a9c46 /* (8, 22, 16) */,
  32'h3db0df4f /* (4, 22, 16) */,
  32'h3d983f17 /* (0, 22, 16) */,
  32'h3e1420e4 /* (28, 18, 16) */,
  32'h3e6dbe20 /* (24, 18, 16) */,
  32'h3ee86d0e /* (20, 18, 16) */,
  32'h3f16cd97 /* (16, 18, 16) */,
  32'h3ee86d0e /* (12, 18, 16) */,
  32'h3e6dbe20 /* (8, 18, 16) */,
  32'h3e1420e4 /* (4, 18, 16) */,
  32'h3dfcae00 /* (0, 18, 16) */,
  32'h3e1420e4 /* (28, 14, 16) */,
  32'h3e6dbe20 /* (24, 14, 16) */,
  32'h3ee86d0e /* (20, 14, 16) */,
  32'h3f16cd97 /* (16, 14, 16) */,
  32'h3ee86d0e /* (12, 14, 16) */,
  32'h3e6dbe20 /* (8, 14, 16) */,
  32'h3e1420e4 /* (4, 14, 16) */,
  32'h3dfcae00 /* (0, 14, 16) */,
  32'h3db0df4f /* (28, 10, 16) */,
  32'h3e0a9c46 /* (24, 10, 16) */,
  32'h3e837a14 /* (20, 10, 16) */,
  32'h3ea594bb /* (16, 10, 16) */,
  32'h3e837a14 /* (12, 10, 16) */,
  32'h3e0a9c46 /* (8, 10, 16) */,
  32'h3db0df4f /* (4, 10, 16) */,
  32'h3d983f17 /* (0, 10, 16) */,
  32'h3d4e2dc2 /* (28, 6, 16) */,
  32'h3d9dd43f /* (24, 6, 16) */,
  32'h3e11854b /* (20, 6, 16) */,
  32'h3e327927 /* (16, 6, 16) */,
  32'h3e11854b /* (12, 6, 16) */,
  32'h3d9dd43f /* (8, 6, 16) */,
  32'h3d4e2dc2 /* (4, 6, 16) */,
  32'h3d332545 /* (0, 6, 16) */,
  32'h3d1c5e8a /* (28, 2, 16) */,
  32'h3d6bb726 /* (24, 2, 16) */,
  32'h3dd576ed /* (20, 2, 16) */,
  32'h3e00d0e8 /* (16, 2, 16) */,
  32'h3dd576ed /* (12, 2, 16) */,
  32'h3d6bb726 /* (8, 2, 16) */,
  32'h3d1c5e8a /* (4, 2, 16) */,
  32'h3d08bc50 /* (0, 2, 16) */,
  32'h3d2ab74a /* (28, 30, 12) */,
  32'h3d69b2a3 /* (24, 30, 12) */,
  32'h3dbf980c /* (20, 30, 12) */,
  32'h3dd576ed /* (16, 30, 12) */,
  32'h3dbf980c /* (12, 30, 12) */,
  32'h3d69b2a3 /* (8, 30, 12) */,
  32'h3d2ab74a /* (4, 30, 12) */,
  32'h3d1bd472 /* (0, 30, 12) */,
  32'h3d522ea6 /* (28, 26, 12) */,
  32'h3d95625b /* (24, 26, 12) */,
  32'h3dfe11f4 /* (20, 26, 12) */,
  32'h3e11854b /* (16, 26, 12) */,
  32'h3dfe11f4 /* (12, 26, 12) */,
  32'h3d95625b /* (8, 26, 12) */,
  32'h3d522ea6 /* (4, 26, 12) */,
  32'h3d3c86f4 /* (0, 26, 12) */,
  32'h3da42ada /* (28, 22, 12) */,
  32'h3df53c17 /* (24, 22, 12) */,
  32'h3e5bd2f1 /* (20, 22, 12) */,
  32'h3e837a14 /* (16, 22, 12) */,
  32'h3e5bd2f1 /* (12, 22, 12) */,
  32'h3df53c17 /* (8, 22, 12) */,
  32'h3da42ada /* (4, 22, 12) */,
  32'h3d9019ab /* (0, 22, 12) */,
  32'h3dfca6c8 /* (28, 18, 12) */,
  32'h3e44fc23 /* (24, 18, 12) */,
  32'h3eb9abaa /* (20, 18, 12) */,
  32'h3ee86d0e /* (16, 18, 12) */,
  32'h3eb9abaa /* (12, 18, 12) */,
  32'h3e44fc23 /* (8, 18, 12) */,
  32'h3dfca6c8 /* (4, 18, 12) */,
  32'h3dd9ea44 /* (0, 18, 12) */,
  32'h3dfca6c8 /* (28, 14, 12) */,
  32'h3e44fc23 /* (24, 14, 12) */,
  32'h3eb9abaa /* (20, 14, 12) */,
  32'h3ee86d0e /* (16, 14, 12) */,
  32'h3eb9abaa /* (12, 14, 12) */,
  32'h3e44fc23 /* (8, 14, 12) */,
  32'h3dfca6c8 /* (4, 14, 12) */,
  32'h3dd9ea44 /* (0, 14, 12) */,
  32'h3da42ada /* (28, 10, 12) */,
  32'h3df53c17 /* (24, 10, 12) */,
  32'h3e5bd2f1 /* (20, 10, 12) */,
  32'h3e837a14 /* (16, 10, 12) */,
  32'h3e5bd2f1 /* (12, 10, 12) */,
  32'h3df53c17 /* (8, 10, 12) */,
  32'h3da42ada /* (4, 10, 12) */,
  32'h3d9019ab /* (0, 10, 12) */,
  32'h3d522ea6 /* (28, 6, 12) */,
  32'h3d95625b /* (24, 6, 12) */,
  32'h3dfe11f4 /* (20, 6, 12) */,
  32'h3e11854b /* (16, 6, 12) */,
  32'h3dfe11f4 /* (12, 6, 12) */,
  32'h3d95625b /* (8, 6, 12) */,
  32'h3d522ea6 /* (4, 6, 12) */,
  32'h3d3c86f4 /* (0, 6, 12) */,
  32'h3d2ab74a /* (28, 2, 12) */,
  32'h3d69b2a3 /* (24, 2, 12) */,
  32'h3dbf980c /* (20, 2, 12) */,
  32'h3dd576ed /* (16, 2, 12) */,
  32'h3dbf980c /* (12, 2, 12) */,
  32'h3d69b2a3 /* (8, 2, 12) */,
  32'h3d2ab74a /* (4, 2, 12) */,
  32'h3d1bd472 /* (0, 2, 12) */,
  32'h3d139519 /* (28, 30, 8) */,
  32'h3d263161 /* (24, 30, 8) */,
  32'h3d69b2a3 /* (20, 30, 8) */,
  32'h3d6bb726 /* (16, 30, 8) */,
  32'h3d69b2a3 /* (12, 30, 8) */,
  32'h3d263161 /* (8, 30, 8) */,
  32'h3d139519 /* (4, 30, 8) */,
  32'h3d162cf4 /* (0, 30, 8) */,
  32'h3d1d3fef /* (28, 26, 8) */,
  32'h3d44d2c5 /* (24, 26, 8) */,
  32'h3d95625b /* (20, 26, 8) */,
  32'h3d9dd43f /* (16, 26, 8) */,
  32'h3d95625b /* (12, 26, 8) */,
  32'h3d44d2c5 /* (8, 26, 8) */,
  32'h3d1d3fef /* (4, 26, 8) */,
  32'h3d164277 /* (0, 26, 8) */,
  32'h3d51ff4c /* (28, 22, 8) */,
  32'h3d92b00e /* (24, 22, 8) */,
  32'h3df53c17 /* (20, 22, 8) */,
  32'h3e0a9c46 /* (16, 22, 8) */,
  32'h3df53c17 /* (12, 22, 8) */,
  32'h3d92b00e /* (8, 22, 8) */,
  32'h3d51ff4c /* (4, 22, 8) */,
  32'h3d3ddc84 /* (0, 22, 8) */,
  32'h3d904c26 /* (28, 18, 8) */,
  32'h3dd9849b /* (24, 18, 8) */,
  32'h3e44fc23 /* (20, 18, 8) */,
  32'h3e6dbe20 /* (16, 18, 8) */,
  32'h3e44fc23 /* (12, 18, 8) */,
  32'h3dd9849b /* (8, 18, 8) */,
  32'h3d904c26 /* (4, 18, 8) */,
  32'h3d7c5be6 /* (0, 18, 8) */,
  32'h3d904c26 /* (28, 14, 8) */,
  32'h3dd9849b /* (24, 14, 8) */,
  32'h3e44fc23 /* (20, 14, 8) */,
  32'h3e6dbe20 /* (16, 14, 8) */,
  32'h3e44fc23 /* (12, 14, 8) */,
  32'h3dd9849b /* (8, 14, 8) */,
  32'h3d904c26 /* (4, 14, 8) */,
  32'h3d7c5be6 /* (0, 14, 8) */,
  32'h3d51ff4c /* (28, 10, 8) */,
  32'h3d92b00e /* (24, 10, 8) */,
  32'h3df53c17 /* (20, 10, 8) */,
  32'h3e0a9c46 /* (16, 10, 8) */,
  32'h3df53c17 /* (12, 10, 8) */,
  32'h3d92b00e /* (8, 10, 8) */,
  32'h3d51ff4c /* (4, 10, 8) */,
  32'h3d3ddc84 /* (0, 10, 8) */,
  32'h3d1d3fef /* (28, 6, 8) */,
  32'h3d44d2c5 /* (24, 6, 8) */,
  32'h3d95625b /* (20, 6, 8) */,
  32'h3d9dd43f /* (16, 6, 8) */,
  32'h3d95625b /* (12, 6, 8) */,
  32'h3d44d2c5 /* (8, 6, 8) */,
  32'h3d1d3fef /* (4, 6, 8) */,
  32'h3d164277 /* (0, 6, 8) */,
  32'h3d139519 /* (28, 2, 8) */,
  32'h3d263161 /* (24, 2, 8) */,
  32'h3d69b2a3 /* (20, 2, 8) */,
  32'h3d6bb726 /* (16, 2, 8) */,
  32'h3d69b2a3 /* (12, 2, 8) */,
  32'h3d263161 /* (8, 2, 8) */,
  32'h3d139519 /* (4, 2, 8) */,
  32'h3d162cf4 /* (0, 2, 8) */,
  32'h3d429928 /* (28, 30, 4) */,
  32'h3d139519 /* (24, 30, 4) */,
  32'h3d2ab74a /* (20, 30, 4) */,
  32'h3d1c5e8a /* (16, 30, 4) */,
  32'h3d2ab74a /* (12, 30, 4) */,
  32'h3d139519 /* (8, 30, 4) */,
  32'h3d429928 /* (4, 30, 4) */,
  32'h3d90451b /* (0, 30, 4) */,
  32'h3d1796af /* (28, 26, 4) */,
  32'h3d1d3fef /* (24, 26, 4) */,
  32'h3d522ea6 /* (20, 26, 4) */,
  32'h3d4e2dc2 /* (16, 26, 4) */,
  32'h3d522ea6 /* (12, 26, 4) */,
  32'h3d1d3fef /* (8, 26, 4) */,
  32'h3d1796af /* (4, 26, 4) */,
  32'h3d234ae8 /* (0, 26, 4) */,
  32'h3d21d2a4 /* (28, 22, 4) */,
  32'h3d51ff4c /* (24, 22, 4) */,
  32'h3da42ada /* (20, 22, 4) */,
  32'h3db0df4f /* (16, 22, 4) */,
  32'h3da42ada /* (12, 22, 4) */,
  32'h3d51ff4c /* (8, 22, 4) */,
  32'h3d21d2a4 /* (4, 22, 4) */,
  32'h3d17b006 /* (0, 22, 4) */,
  32'h3d456b70 /* (28, 18, 4) */,
  32'h3d904c26 /* (24, 18, 4) */,
  32'h3dfca6c8 /* (20, 18, 4) */,
  32'h3e1420e4 /* (16, 18, 4) */,
  32'h3dfca6c8 /* (12, 18, 4) */,
  32'h3d904c26 /* (8, 18, 4) */,
  32'h3d456b70 /* (4, 18, 4) */,
  32'h3d2ee5c8 /* (0, 18, 4) */,
  32'h3d456b70 /* (28, 14, 4) */,
  32'h3d904c26 /* (24, 14, 4) */,
  32'h3dfca6c8 /* (20, 14, 4) */,
  32'h3e1420e4 /* (16, 14, 4) */,
  32'h3dfca6c8 /* (12, 14, 4) */,
  32'h3d904c26 /* (8, 14, 4) */,
  32'h3d456b70 /* (4, 14, 4) */,
  32'h3d2ee5c8 /* (0, 14, 4) */,
  32'h3d21d2a4 /* (28, 10, 4) */,
  32'h3d51ff4c /* (24, 10, 4) */,
  32'h3da42ada /* (20, 10, 4) */,
  32'h3db0df4f /* (16, 10, 4) */,
  32'h3da42ada /* (12, 10, 4) */,
  32'h3d51ff4c /* (8, 10, 4) */,
  32'h3d21d2a4 /* (4, 10, 4) */,
  32'h3d17b006 /* (0, 10, 4) */,
  32'h3d1796af /* (28, 6, 4) */,
  32'h3d1d3fef /* (24, 6, 4) */,
  32'h3d522ea6 /* (20, 6, 4) */,
  32'h3d4e2dc2 /* (16, 6, 4) */,
  32'h3d522ea6 /* (12, 6, 4) */,
  32'h3d1d3fef /* (8, 6, 4) */,
  32'h3d1796af /* (4, 6, 4) */,
  32'h3d234ae8 /* (0, 6, 4) */,
  32'h3d429928 /* (28, 2, 4) */,
  32'h3d139519 /* (24, 2, 4) */,
  32'h3d2ab74a /* (20, 2, 4) */,
  32'h3d1c5e8a /* (16, 2, 4) */,
  32'h3d2ab74a /* (12, 2, 4) */,
  32'h3d139519 /* (8, 2, 4) */,
  32'h3d429928 /* (4, 2, 4) */,
  32'h3d90451b /* (0, 2, 4) */,
  32'h3d90451b /* (28, 30, 0) */,
  32'h3d162cf4 /* (24, 30, 0) */,
  32'h3d1bd472 /* (20, 30, 0) */,
  32'h3d08bc50 /* (16, 30, 0) */,
  32'h3d1bd472 /* (12, 30, 0) */,
  32'h3d162cf4 /* (8, 30, 0) */,
  32'h3d90451b /* (4, 30, 0) */,
  32'h3e948d77 /* (0, 30, 0) */,
  32'h3d234ae8 /* (28, 26, 0) */,
  32'h3d164277 /* (24, 26, 0) */,
  32'h3d3c86f4 /* (20, 26, 0) */,
  32'h3d332545 /* (16, 26, 0) */,
  32'h3d3c86f4 /* (12, 26, 0) */,
  32'h3d164277 /* (8, 26, 0) */,
  32'h3d234ae8 /* (4, 26, 0) */,
  32'h3d424b89 /* (0, 26, 0) */,
  32'h3d17b006 /* (28, 22, 0) */,
  32'h3d3ddc84 /* (24, 22, 0) */,
  32'h3d9019ab /* (20, 22, 0) */,
  32'h3d983f17 /* (16, 22, 0) */,
  32'h3d9019ab /* (12, 22, 0) */,
  32'h3d3ddc84 /* (8, 22, 0) */,
  32'h3d17b006 /* (4, 22, 0) */,
  32'h3d10f1da /* (0, 22, 0) */,
  32'h3d2ee5c8 /* (28, 18, 0) */,
  32'h3d7c5be6 /* (24, 18, 0) */,
  32'h3dd9ea44 /* (20, 18, 0) */,
  32'h3dfcae00 /* (16, 18, 0) */,
  32'h3dd9ea44 /* (12, 18, 0) */,
  32'h3d7c5be6 /* (8, 18, 0) */,
  32'h3d2ee5c8 /* (4, 18, 0) */,
  32'h3d1bd51d /* (0, 18, 0) */,
  32'h3d2ee5c8 /* (28, 14, 0) */,
  32'h3d7c5be6 /* (24, 14, 0) */,
  32'h3dd9ea44 /* (20, 14, 0) */,
  32'h3dfcae00 /* (16, 14, 0) */,
  32'h3dd9ea44 /* (12, 14, 0) */,
  32'h3d7c5be6 /* (8, 14, 0) */,
  32'h3d2ee5c8 /* (4, 14, 0) */,
  32'h3d1bd51d /* (0, 14, 0) */,
  32'h3d17b006 /* (28, 10, 0) */,
  32'h3d3ddc84 /* (24, 10, 0) */,
  32'h3d9019ab /* (20, 10, 0) */,
  32'h3d983f17 /* (16, 10, 0) */,
  32'h3d9019ab /* (12, 10, 0) */,
  32'h3d3ddc84 /* (8, 10, 0) */,
  32'h3d17b006 /* (4, 10, 0) */,
  32'h3d10f1da /* (0, 10, 0) */,
  32'h3d234ae8 /* (28, 6, 0) */,
  32'h3d164277 /* (24, 6, 0) */,
  32'h3d3c86f4 /* (20, 6, 0) */,
  32'h3d332545 /* (16, 6, 0) */,
  32'h3d3c86f4 /* (12, 6, 0) */,
  32'h3d164277 /* (8, 6, 0) */,
  32'h3d234ae8 /* (4, 6, 0) */,
  32'h3d424b89 /* (0, 6, 0) */,
  32'h3d90451b /* (28, 2, 0) */,
  32'h3d162cf4 /* (24, 2, 0) */,
  32'h3d1bd472 /* (20, 2, 0) */,
  32'h3d08bc50 /* (16, 2, 0) */,
  32'h3d1bd472 /* (12, 2, 0) */,
  32'h3d162cf4 /* (8, 2, 0) */,
  32'h3d90451b /* (4, 2, 0) */,
  32'h3e948d77 /* (0, 2, 0) */,
  32'h3d6eb36b /* (31, 29, 28) */,
  32'h3d25f5ce /* (27, 29, 28) */,
  32'h3d16b5b2 /* (23, 29, 28) */,
  32'h3d385879 /* (19, 29, 28) */,
  32'h3d349293 /* (15, 29, 28) */,
  32'h3d25fa09 /* (11, 29, 28) */,
  32'h3d155fa4 /* (7, 29, 28) */,
  32'h3d4920d0 /* (3, 29, 28) */,
  32'h3d17ff6b /* (31, 25, 28) */,
  32'h3d1508af /* (27, 25, 28) */,
  32'h3d30de15 /* (23, 25, 28) */,
  32'h3d770afc /* (19, 25, 28) */,
  32'h3d7b9f11 /* (15, 25, 28) */,
  32'h3d52976b /* (11, 25, 28) */,
  32'h3d1cbb18 /* (7, 25, 28) */,
  32'h3d155fa4 /* (3, 25, 28) */,
  32'h3d1f5dc3 /* (31, 21, 28) */,
  32'h3d358341 /* (27, 21, 28) */,
  32'h3d81d711 /* (23, 21, 28) */,
  32'h3dcf13a3 /* (19, 21, 28) */,
  32'h3ddcf428 /* (15, 21, 28) */,
  32'h3da66ad4 /* (11, 21, 28) */,
  32'h3d52976b /* (7, 21, 28) */,
  32'h3d25fa09 /* (3, 21, 28) */,
  32'h3d294c4b /* (31, 17, 28) */,
  32'h3d4def9b /* (27, 17, 28) */,
  32'h3da3c1ed /* (23, 17, 28) */,
  32'h3e0ff4ce /* (19, 17, 28) */,
  32'h3e1fe07e /* (15, 17, 28) */,
  32'h3ddcf428 /* (11, 17, 28) */,
  32'h3d7b9f11 /* (7, 17, 28) */,
  32'h3d349293 /* (3, 17, 28) */,
  32'h3d2e802a /* (31, 13, 28) */,
  32'h3d4ea6a0 /* (27, 13, 28) */,
  32'h3d9d0afa /* (23, 13, 28) */,
  32'h3e0415cb /* (19, 13, 28) */,
  32'h3e0ff4ce /* (15, 13, 28) */,
  32'h3dcf13a3 /* (11, 13, 28) */,
  32'h3d770afc /* (7, 13, 28) */,
  32'h3d385879 /* (3, 13, 28) */,
  32'h3d13f199 /* (31, 9, 28) */,
  32'h3d1ee50b /* (27, 9, 28) */,
  32'h3d51a9d2 /* (23, 9, 28) */,
  32'h3d9d0afa /* (19, 9, 28) */,
  32'h3da3c1ed /* (15, 9, 28) */,
  32'h3d81d711 /* (11, 9, 28) */,
  32'h3d30de15 /* (7, 9, 28) */,
  32'h3d16b5b2 /* (3, 9, 28) */,
  32'h3d334ee4 /* (31, 5, 28) */,
  32'h3d189061 /* (27, 5, 28) */,
  32'h3d1ee50b /* (23, 5, 28) */,
  32'h3d4ea6a0 /* (19, 5, 28) */,
  32'h3d4def9b /* (15, 5, 28) */,
  32'h3d358341 /* (11, 5, 28) */,
  32'h3d1508af /* (7, 5, 28) */,
  32'h3d25f5ce /* (3, 5, 28) */,
  32'h3d9c757b /* (31, 1, 28) */,
  32'h3d334ee4 /* (27, 1, 28) */,
  32'h3d13f199 /* (23, 1, 28) */,
  32'h3d2e802a /* (19, 1, 28) */,
  32'h3d294c4b /* (15, 1, 28) */,
  32'h3d1f5dc3 /* (11, 1, 28) */,
  32'h3d17ff6b /* (7, 1, 28) */,
  32'h3d6eb36b /* (3, 1, 28) */,
  32'h3d146963 /* (31, 29, 24) */,
  32'h3d15d660 /* (27, 29, 24) */,
  32'h3d37919e /* (23, 29, 24) */,
  32'h3d82c188 /* (19, 29, 24) */,
  32'h3d8608f0 /* (15, 29, 24) */,
  32'h3d5d0a38 /* (11, 29, 24) */,
  32'h3d2054cd /* (7, 29, 24) */,
  32'h3d1392fe /* (3, 29, 24) */,
  32'h3d1bb8b6 /* (31, 25, 24) */,
  32'h3d2bff3e /* (27, 25, 24) */,
  32'h3d6b8b35 /* (23, 25, 24) */,
  32'h3db56072 /* (19, 25, 24) */,
  32'h3dbf0444 /* (15, 25, 24) */,
  32'h3d941bce /* (11, 25, 24) */,
  32'h3d432bf1 /* (7, 25, 24) */,
  32'h3d2054cd /* (3, 25, 24) */,
  32'h3d513c3d /* (31, 21, 24) */,
  32'h3d77c8fd /* (27, 21, 24) */,
  32'h3dbc4d73 /* (23, 21, 24) */,
  32'h3e1e607d /* (19, 21, 24) */,
  32'h3e2c9c6c /* (15, 21, 24) */,
  32'h3df84bb3 /* (11, 21, 24) */,
  32'h3d941bce /* (7, 21, 24) */,
  32'h3d5d0a38 /* (3, 21, 24) */,
  32'h3d7a003f /* (31, 17, 24) */,
  32'h3d9a5b6b /* (27, 17, 24) */,
  32'h3dfc30a3 /* (23, 17, 24) */,
  32'h3e640ba2 /* (19, 17, 24) */,
  32'h3e803f85 /* (15, 17, 24) */,
  32'h3e2c9c6c /* (11, 17, 24) */,
  32'h3dbf0444 /* (7, 17, 24) */,
  32'h3d8608f0 /* (3, 17, 24) */,
  32'h3d7573b6 /* (31, 13, 24) */,
  32'h3d94d380 /* (27, 13, 24) */,
  32'h3deb6b6d /* (23, 13, 24) */,
  32'h3e4dd3dc /* (19, 13, 24) */,
  32'h3e640ba2 /* (15, 13, 24) */,
  32'h3e1e607d /* (11, 13, 24) */,
  32'h3db56072 /* (7, 13, 24) */,
  32'h3d82c188 /* (3, 13, 24) */,
  32'h3d2fba80 /* (31, 9, 24) */,
  32'h3d49c96c /* (27, 9, 24) */,
  32'h3d921bde /* (23, 9, 24) */,
  32'h3deb6b6d /* (19, 9, 24) */,
  32'h3dfc30a3 /* (15, 9, 24) */,
  32'h3dbc4d73 /* (11, 9, 24) */,
  32'h3d6b8b35 /* (7, 9, 24) */,
  32'h3d37919e /* (3, 9, 24) */,
  32'h3d1412fd /* (31, 5, 24) */,
  32'h3d1c4d38 /* (27, 5, 24) */,
  32'h3d49c96c /* (23, 5, 24) */,
  32'h3d94d380 /* (19, 5, 24) */,
  32'h3d9a5b6b /* (15, 5, 24) */,
  32'h3d77c8fd /* (11, 5, 24) */,
  32'h3d2bff3e /* (7, 5, 24) */,
  32'h3d15d660 /* (3, 5, 24) */,
  32'h3d1704d7 /* (31, 1, 24) */,
  32'h3d1412fd /* (27, 1, 24) */,
  32'h3d2fba80 /* (23, 1, 24) */,
  32'h3d7573b6 /* (19, 1, 24) */,
  32'h3d7a003f /* (15, 1, 24) */,
  32'h3d513c3d /* (11, 1, 24) */,
  32'h3d1bb8b6 /* (7, 1, 24) */,
  32'h3d146963 /* (3, 1, 24) */,
  32'h3d210eee /* (31, 29, 20) */,
  32'h3d3a4ebb /* (27, 29, 20) */,
  32'h3d886b82 /* (23, 29, 20) */,
  32'h3dddef48 /* (19, 29, 20) */,
  32'h3deea44d /* (15, 29, 20) */,
  32'h3db0b965 /* (11, 29, 20) */,
  32'h3d5ab0e1 /* (7, 29, 20) */,
  32'h3d28b308 /* (3, 29, 20) */,
  32'h3d4ea8e5 /* (31, 25, 20) */,
  32'h3d75e4d4 /* (27, 25, 20) */,
  32'h3dbc51f9 /* (23, 25, 20) */,
  32'h3e1f8cbf /* (19, 25, 20) */,
  32'h3e2e6a71 /* (15, 25, 20) */,
  32'h3df94537 /* (11, 25, 20) */,
  32'h3d938890 /* (7, 25, 20) */,
  32'h3d5ab0e1 /* (3, 25, 20) */,
  32'h3da53628 /* (31, 21, 20) */,
  32'h3dca9d53 /* (27, 21, 20) */,
  32'h3e23781b /* (23, 21, 20) */,
  32'h3e91dfe2 /* (19, 21, 20) */,
  32'h3ea31756 /* (15, 21, 20) */,
  32'h3e5e44ac /* (11, 21, 20) */,
  32'h3df94537 /* (7, 21, 20) */,
  32'h3db0b965 /* (3, 21, 20) */,
  32'h3ddd43c2 /* (31, 17, 20) */,
  32'h3e0ae903 /* (27, 17, 20) */,
  32'h3e6a25fd /* (23, 17, 20) */,
  32'h3edb3822 /* (19, 17, 20) */,
  32'h3efaa119 /* (15, 17, 20) */,
  32'h3ea31756 /* (11, 17, 20) */,
  32'h3e2e6a71 /* (7, 17, 20) */,
  32'h3deea44d /* (3, 17, 20) */,
  32'h3dce8d02 /* (31, 13, 20) */,
  32'h3e00477d /* (27, 13, 20) */,
  32'h3e53dc51 /* (23, 13, 20) */,
  32'h3ec1d890 /* (19, 13, 20) */,
  32'h3edb3822 /* (15, 13, 20) */,
  32'h3e91dfe2 /* (11, 13, 20) */,
  32'h3e1f8cbf /* (7, 13, 20) */,
  32'h3dddef48 /* (3, 13, 20) */,
  32'h3d803124 /* (31, 9, 20) */,
  32'h3d9af1c2 /* (27, 9, 20) */,
  32'h3df3b4f2 /* (23, 9, 20) */,
  32'h3e53dc51 /* (19, 9, 20) */,
  32'h3e6a25fd /* (15, 9, 20) */,
  32'h3e23781b /* (11, 9, 20) */,
  32'h3dbc51f9 /* (7, 9, 20) */,
  32'h3d886b82 /* (3, 9, 20) */,
  32'h3d310ad3 /* (31, 5, 20) */,
  32'h3d4f6dfc /* (27, 5, 20) */,
  32'h3d9af1c2 /* (23, 5, 20) */,
  32'h3e00477d /* (19, 5, 20) */,
  32'h3e0ae903 /* (15, 5, 20) */,
  32'h3dca9d53 /* (11, 5, 20) */,
  32'h3d75e4d4 /* (7, 5, 20) */,
  32'h3d3a4ebb /* (3, 5, 20) */,
  32'h3d1a2df1 /* (31, 1, 20) */,
  32'h3d310ad3 /* (27, 1, 20) */,
  32'h3d803124 /* (23, 1, 20) */,
  32'h3dce8d02 /* (19, 1, 20) */,
  32'h3ddd43c2 /* (15, 1, 20) */,
  32'h3da53628 /* (11, 1, 20) */,
  32'h3d4ea8e5 /* (7, 1, 20) */,
  32'h3d210eee /* (3, 1, 20) */,
  32'h3d0fbc59 /* (31, 29, 16) */,
  32'h3d3046d8 /* (27, 29, 16) */,
  32'h3d8e3848 /* (23, 29, 16) */,
  32'h3dfdd31f /* (19, 29, 16) */,
  32'h3e0de417 /* (15, 29, 16) */,
  32'h3dc1602b /* (11, 29, 16) */,
  32'h3d58de26 /* (7, 29, 16) */,
  32'h3d19c07a /* (3, 29, 16) */,
  32'h3d49f75a /* (31, 25, 16) */,
  32'h3d7a662c /* (27, 25, 16) */,
  32'h3dce1075 /* (23, 25, 16) */,
  32'h3e3bd4ee /* (19, 25, 16) */,
  32'h3e540b9b /* (15, 25, 16) */,
  32'h3e0d9cf0 /* (11, 25, 16) */,
  32'h3d9b7830 /* (7, 25, 16) */,
  32'h3d58de26 /* (3, 25, 16) */,
  32'h3db336e0 /* (31, 21, 16) */,
  32'h3de14ffa /* (27, 21, 16) */,
  32'h3e3e5da7 /* (23, 21, 16) */,
  32'h3eb2bd2a /* (19, 21, 16) */,
  32'h3ecca1ac /* (15, 21, 16) */,
  32'h3e84c8e0 /* (11, 21, 16) */,
  32'h3e0d9cf0 /* (7, 21, 16) */,
  32'h3dc1602b /* (3, 21, 16) */,
  32'h3e02e976 /* (31, 17, 16) */,
  32'h3e26bbbb /* (27, 17, 16) */,
  32'h3e908107 /* (23, 17, 16) */,
  32'h3f0bd969 /* (19, 17, 16) */,
  32'h3f2286f8 /* (15, 17, 16) */,
  32'h3ecca1ac /* (11, 17, 16) */,
  32'h3e540b9b /* (7, 17, 16) */,
  32'h3e0de417 /* (3, 17, 16) */,
  32'h3deaafef /* (31, 13, 16) */,
  32'h3e1486b7 /* (27, 13, 16) */,
  32'h3e7e4b9d /* (23, 13, 16) */,
  32'h3ef27895 /* (19, 13, 16) */,
  32'h3f0bd969 /* (15, 13, 16) */,
  32'h3eb2bd2a /* (11, 13, 16) */,
  32'h3e3bd4ee /* (7, 13, 16) */,
  32'h3dfdd31f /* (3, 13, 16) */,
  32'h3d8420c9 /* (31, 9, 16) */,
  32'h3da4f2f4 /* (27, 9, 16) */,
  32'h3e0981d7 /* (23, 9, 16) */,
  32'h3e7e4b9d /* (19, 9, 16) */,
  32'h3e908107 /* (15, 9, 16) */,
  32'h3e3e5da7 /* (11, 9, 16) */,
  32'h3dce1075 /* (7, 9, 16) */,
  32'h3d8e3848 /* (3, 9, 16) */,
  32'h3d24852f /* (31, 5, 16) */,
  32'h3d4ab7f7 /* (27, 5, 16) */,
  32'h3da4f2f4 /* (23, 5, 16) */,
  32'h3e1486b7 /* (19, 5, 16) */,
  32'h3e26bbbb /* (15, 5, 16) */,
  32'h3de14ffa /* (11, 5, 16) */,
  32'h3d7a662c /* (7, 5, 16) */,
  32'h3d3046d8 /* (3, 5, 16) */,
  32'h3d067e68 /* (31, 1, 16) */,
  32'h3d24852f /* (27, 1, 16) */,
  32'h3d8420c9 /* (23, 1, 16) */,
  32'h3deaafef /* (19, 1, 16) */,
  32'h3e02e976 /* (15, 1, 16) */,
  32'h3db336e0 /* (11, 1, 16) */,
  32'h3d49f75a /* (7, 1, 16) */,
  32'h3d0fbc59 /* (3, 1, 16) */,
  32'h3d210eee /* (31, 29, 12) */,
  32'h3d3a4ebb /* (27, 29, 12) */,
  32'h3d886b82 /* (23, 29, 12) */,
  32'h3dddef48 /* (19, 29, 12) */,
  32'h3deea44d /* (15, 29, 12) */,
  32'h3db0b965 /* (11, 29, 12) */,
  32'h3d5ab0e1 /* (7, 29, 12) */,
  32'h3d28b308 /* (3, 29, 12) */,
  32'h3d4ea8e5 /* (31, 25, 12) */,
  32'h3d75e4d4 /* (27, 25, 12) */,
  32'h3dbc51f9 /* (23, 25, 12) */,
  32'h3e1f8cbf /* (19, 25, 12) */,
  32'h3e2e6a71 /* (15, 25, 12) */,
  32'h3df94537 /* (11, 25, 12) */,
  32'h3d938890 /* (7, 25, 12) */,
  32'h3d5ab0e1 /* (3, 25, 12) */,
  32'h3da53628 /* (31, 21, 12) */,
  32'h3dca9d53 /* (27, 21, 12) */,
  32'h3e23781b /* (23, 21, 12) */,
  32'h3e91dfe2 /* (19, 21, 12) */,
  32'h3ea31756 /* (15, 21, 12) */,
  32'h3e5e44ac /* (11, 21, 12) */,
  32'h3df94537 /* (7, 21, 12) */,
  32'h3db0b965 /* (3, 21, 12) */,
  32'h3ddd43c2 /* (31, 17, 12) */,
  32'h3e0ae903 /* (27, 17, 12) */,
  32'h3e6a25fd /* (23, 17, 12) */,
  32'h3edb3822 /* (19, 17, 12) */,
  32'h3efaa119 /* (15, 17, 12) */,
  32'h3ea31756 /* (11, 17, 12) */,
  32'h3e2e6a71 /* (7, 17, 12) */,
  32'h3deea44d /* (3, 17, 12) */,
  32'h3dce8d02 /* (31, 13, 12) */,
  32'h3e00477d /* (27, 13, 12) */,
  32'h3e53dc51 /* (23, 13, 12) */,
  32'h3ec1d890 /* (19, 13, 12) */,
  32'h3edb3822 /* (15, 13, 12) */,
  32'h3e91dfe2 /* (11, 13, 12) */,
  32'h3e1f8cbf /* (7, 13, 12) */,
  32'h3dddef48 /* (3, 13, 12) */,
  32'h3d803124 /* (31, 9, 12) */,
  32'h3d9af1c2 /* (27, 9, 12) */,
  32'h3df3b4f2 /* (23, 9, 12) */,
  32'h3e53dc51 /* (19, 9, 12) */,
  32'h3e6a25fd /* (15, 9, 12) */,
  32'h3e23781b /* (11, 9, 12) */,
  32'h3dbc51f9 /* (7, 9, 12) */,
  32'h3d886b82 /* (3, 9, 12) */,
  32'h3d310ad3 /* (31, 5, 12) */,
  32'h3d4f6dfc /* (27, 5, 12) */,
  32'h3d9af1c2 /* (23, 5, 12) */,
  32'h3e00477d /* (19, 5, 12) */,
  32'h3e0ae903 /* (15, 5, 12) */,
  32'h3dca9d53 /* (11, 5, 12) */,
  32'h3d75e4d4 /* (7, 5, 12) */,
  32'h3d3a4ebb /* (3, 5, 12) */,
  32'h3d1a2df1 /* (31, 1, 12) */,
  32'h3d310ad3 /* (27, 1, 12) */,
  32'h3d803124 /* (23, 1, 12) */,
  32'h3dce8d02 /* (19, 1, 12) */,
  32'h3ddd43c2 /* (15, 1, 12) */,
  32'h3da53628 /* (11, 1, 12) */,
  32'h3d4ea8e5 /* (7, 1, 12) */,
  32'h3d210eee /* (3, 1, 12) */,
  32'h3d146963 /* (31, 29, 8) */,
  32'h3d15d660 /* (27, 29, 8) */,
  32'h3d37919e /* (23, 29, 8) */,
  32'h3d82c188 /* (19, 29, 8) */,
  32'h3d8608f0 /* (15, 29, 8) */,
  32'h3d5d0a38 /* (11, 29, 8) */,
  32'h3d2054cd /* (7, 29, 8) */,
  32'h3d1392fe /* (3, 29, 8) */,
  32'h3d1bb8b6 /* (31, 25, 8) */,
  32'h3d2bff3e /* (27, 25, 8) */,
  32'h3d6b8b35 /* (23, 25, 8) */,
  32'h3db56072 /* (19, 25, 8) */,
  32'h3dbf0444 /* (15, 25, 8) */,
  32'h3d941bce /* (11, 25, 8) */,
  32'h3d432bf1 /* (7, 25, 8) */,
  32'h3d2054cd /* (3, 25, 8) */,
  32'h3d513c3d /* (31, 21, 8) */,
  32'h3d77c8fd /* (27, 21, 8) */,
  32'h3dbc4d73 /* (23, 21, 8) */,
  32'h3e1e607d /* (19, 21, 8) */,
  32'h3e2c9c6c /* (15, 21, 8) */,
  32'h3df84bb3 /* (11, 21, 8) */,
  32'h3d941bce /* (7, 21, 8) */,
  32'h3d5d0a38 /* (3, 21, 8) */,
  32'h3d7a003f /* (31, 17, 8) */,
  32'h3d9a5b6b /* (27, 17, 8) */,
  32'h3dfc30a3 /* (23, 17, 8) */,
  32'h3e640ba2 /* (19, 17, 8) */,
  32'h3e803f85 /* (15, 17, 8) */,
  32'h3e2c9c6c /* (11, 17, 8) */,
  32'h3dbf0444 /* (7, 17, 8) */,
  32'h3d8608f0 /* (3, 17, 8) */,
  32'h3d7573b6 /* (31, 13, 8) */,
  32'h3d94d380 /* (27, 13, 8) */,
  32'h3deb6b6d /* (23, 13, 8) */,
  32'h3e4dd3dc /* (19, 13, 8) */,
  32'h3e640ba2 /* (15, 13, 8) */,
  32'h3e1e607d /* (11, 13, 8) */,
  32'h3db56072 /* (7, 13, 8) */,
  32'h3d82c188 /* (3, 13, 8) */,
  32'h3d2fba80 /* (31, 9, 8) */,
  32'h3d49c96c /* (27, 9, 8) */,
  32'h3d921bde /* (23, 9, 8) */,
  32'h3deb6b6d /* (19, 9, 8) */,
  32'h3dfc30a3 /* (15, 9, 8) */,
  32'h3dbc4d73 /* (11, 9, 8) */,
  32'h3d6b8b35 /* (7, 9, 8) */,
  32'h3d37919e /* (3, 9, 8) */,
  32'h3d1412fd /* (31, 5, 8) */,
  32'h3d1c4d38 /* (27, 5, 8) */,
  32'h3d49c96c /* (23, 5, 8) */,
  32'h3d94d380 /* (19, 5, 8) */,
  32'h3d9a5b6b /* (15, 5, 8) */,
  32'h3d77c8fd /* (11, 5, 8) */,
  32'h3d2bff3e /* (7, 5, 8) */,
  32'h3d15d660 /* (3, 5, 8) */,
  32'h3d1704d7 /* (31, 1, 8) */,
  32'h3d1412fd /* (27, 1, 8) */,
  32'h3d2fba80 /* (23, 1, 8) */,
  32'h3d7573b6 /* (19, 1, 8) */,
  32'h3d7a003f /* (15, 1, 8) */,
  32'h3d513c3d /* (11, 1, 8) */,
  32'h3d1bb8b6 /* (7, 1, 8) */,
  32'h3d146963 /* (3, 1, 8) */,
  32'h3d6eb36b /* (31, 29, 4) */,
  32'h3d25f5ce /* (27, 29, 4) */,
  32'h3d16b5b2 /* (23, 29, 4) */,
  32'h3d385879 /* (19, 29, 4) */,
  32'h3d349293 /* (15, 29, 4) */,
  32'h3d25fa09 /* (11, 29, 4) */,
  32'h3d155fa4 /* (7, 29, 4) */,
  32'h3d4920d0 /* (3, 29, 4) */,
  32'h3d17ff6b /* (31, 25, 4) */,
  32'h3d1508af /* (27, 25, 4) */,
  32'h3d30de15 /* (23, 25, 4) */,
  32'h3d770afc /* (19, 25, 4) */,
  32'h3d7b9f11 /* (15, 25, 4) */,
  32'h3d52976b /* (11, 25, 4) */,
  32'h3d1cbb18 /* (7, 25, 4) */,
  32'h3d155fa4 /* (3, 25, 4) */,
  32'h3d1f5dc3 /* (31, 21, 4) */,
  32'h3d358341 /* (27, 21, 4) */,
  32'h3d81d711 /* (23, 21, 4) */,
  32'h3dcf13a3 /* (19, 21, 4) */,
  32'h3ddcf428 /* (15, 21, 4) */,
  32'h3da66ad4 /* (11, 21, 4) */,
  32'h3d52976b /* (7, 21, 4) */,
  32'h3d25fa09 /* (3, 21, 4) */,
  32'h3d294c4b /* (31, 17, 4) */,
  32'h3d4def9b /* (27, 17, 4) */,
  32'h3da3c1ed /* (23, 17, 4) */,
  32'h3e0ff4ce /* (19, 17, 4) */,
  32'h3e1fe07e /* (15, 17, 4) */,
  32'h3ddcf428 /* (11, 17, 4) */,
  32'h3d7b9f11 /* (7, 17, 4) */,
  32'h3d349293 /* (3, 17, 4) */,
  32'h3d2e802a /* (31, 13, 4) */,
  32'h3d4ea6a0 /* (27, 13, 4) */,
  32'h3d9d0afa /* (23, 13, 4) */,
  32'h3e0415cb /* (19, 13, 4) */,
  32'h3e0ff4ce /* (15, 13, 4) */,
  32'h3dcf13a3 /* (11, 13, 4) */,
  32'h3d770afc /* (7, 13, 4) */,
  32'h3d385879 /* (3, 13, 4) */,
  32'h3d13f199 /* (31, 9, 4) */,
  32'h3d1ee50b /* (27, 9, 4) */,
  32'h3d51a9d2 /* (23, 9, 4) */,
  32'h3d9d0afa /* (19, 9, 4) */,
  32'h3da3c1ed /* (15, 9, 4) */,
  32'h3d81d711 /* (11, 9, 4) */,
  32'h3d30de15 /* (7, 9, 4) */,
  32'h3d16b5b2 /* (3, 9, 4) */,
  32'h3d334ee4 /* (31, 5, 4) */,
  32'h3d189061 /* (27, 5, 4) */,
  32'h3d1ee50b /* (23, 5, 4) */,
  32'h3d4ea6a0 /* (19, 5, 4) */,
  32'h3d4def9b /* (15, 5, 4) */,
  32'h3d358341 /* (11, 5, 4) */,
  32'h3d1508af /* (7, 5, 4) */,
  32'h3d25f5ce /* (3, 5, 4) */,
  32'h3d9c757b /* (31, 1, 4) */,
  32'h3d334ee4 /* (27, 1, 4) */,
  32'h3d13f199 /* (23, 1, 4) */,
  32'h3d2e802a /* (19, 1, 4) */,
  32'h3d294c4b /* (15, 1, 4) */,
  32'h3d1f5dc3 /* (11, 1, 4) */,
  32'h3d17ff6b /* (7, 1, 4) */,
  32'h3d6eb36b /* (3, 1, 4) */,
  32'h3dff9e3f /* (31, 29, 0) */,
  32'h3d490b0e /* (27, 29, 0) */,
  32'h3d1237a7 /* (23, 29, 0) */,
  32'h3d258110 /* (19, 29, 0) */,
  32'h3d1eeabe /* (15, 29, 0) */,
  32'h3d198ce9 /* (11, 29, 0) */,
  32'h3d1cfd70 /* (7, 29, 0) */,
  32'h3d9c797c /* (3, 29, 0) */,
  32'h3d25463b /* (31, 25, 0) */,
  32'h3d154f7b /* (27, 25, 0) */,
  32'h3d23a039 /* (23, 25, 0) */,
  32'h3d5a6fdd /* (19, 25, 0) */,
  32'h3d5b6048 /* (15, 25, 0) */,
  32'h3d3dcd22 /* (11, 25, 0) */,
  32'h3d162f74 /* (7, 25, 0) */,
  32'h3d1cfd70 /* (3, 25, 0) */,
  32'h3d147e90 /* (31, 21, 0) */,
  32'h3d25e815 /* (27, 21, 0) */,
  32'h3d66dac1 /* (23, 21, 0) */,
  32'h3db3fd83 /* (19, 21, 0) */,
  32'h3dbe6d47 /* (15, 21, 0) */,
  32'h3d922642 /* (11, 21, 0) */,
  32'h3d3dcd22 /* (7, 21, 0) */,
  32'h3d198ce9 /* (3, 21, 0) */,
  32'h3d155505 /* (31, 17, 0) */,
  32'h3d347f0a /* (27, 17, 0) */,
  32'h3d8df2c1 /* (23, 17, 0) */,
  32'h3df6cc6d /* (19, 17, 0) */,
  32'h3e086183 /* (15, 17, 0) */,
  32'h3dbe6d47 /* (11, 17, 0) */,
  32'h3d5b6048 /* (7, 17, 0) */,
  32'h3d1eeabe /* (3, 17, 0) */,
  32'h3d1d4601 /* (31, 13, 0) */,
  32'h3d384488 /* (27, 13, 0) */,
  32'h3d89a49e /* (23, 13, 0) */,
  32'h3de3e928 /* (19, 13, 0) */,
  32'h3df6cc6d /* (15, 13, 0) */,
  32'h3db3fd83 /* (11, 13, 0) */,
  32'h3d5a6fdd /* (7, 13, 0) */,
  32'h3d258110 /* (3, 13, 0) */,
  32'h3d11a5c6 /* (31, 9, 0) */,
  32'h3d16a564 /* (27, 9, 0) */,
  32'h3d3dc47d /* (23, 9, 0) */,
  32'h3d89a49e /* (19, 9, 0) */,
  32'h3d8df2c1 /* (15, 9, 0) */,
  32'h3d66dac1 /* (11, 9, 0) */,
  32'h3d23a039 /* (7, 9, 0) */,
  32'h3d1237a7 /* (3, 9, 0) */,
  32'h3d6e9998 /* (31, 5, 0) */,
  32'h3d25e3da /* (27, 5, 0) */,
  32'h3d16a564 /* (23, 5, 0) */,
  32'h3d384488 /* (19, 5, 0) */,
  32'h3d347f0a /* (15, 5, 0) */,
  32'h3d25e815 /* (11, 5, 0) */,
  32'h3d154f7b /* (7, 5, 0) */,
  32'h3d490b0e /* (3, 5, 0) */,
  32'h3f10fe39 /* (31, 1, 0) */,
  32'h3d6e9998 /* (27, 1, 0) */,
  32'h3d11a5c6 /* (23, 1, 0) */,
  32'h3d1d4601 /* (19, 1, 0) */,
  32'h3d155505 /* (15, 1, 0) */,
  32'h3d147e90 /* (11, 1, 0) */,
  32'h3d25463b /* (7, 1, 0) */,
  32'h3dff9e3f /* (3, 1, 0) */,
  32'h3d5defd3 /* (30, 29, 28) */,
  32'h3d1b3fff /* (26, 29, 28) */,
  32'h3d1cff11 /* (22, 29, 28) */,
  32'h3d3b1e93 /* (18, 29, 28) */,
  32'h3d3b1e93 /* (14, 29, 28) */,
  32'h3d1cff11 /* (10, 29, 28) */,
  32'h3d1b3fff /* (6, 29, 28) */,
  32'h3d5defd3 /* (2, 29, 28) */,
  32'h3d16c6a3 /* (30, 25, 28) */,
  32'h3d17902e /* (26, 25, 28) */,
  32'h3d404057 /* (22, 25, 28) */,
  32'h3d800deb /* (18, 25, 28) */,
  32'h3d800deb /* (14, 25, 28) */,
  32'h3d404057 /* (10, 25, 28) */,
  32'h3d17902e /* (6, 25, 28) */,
  32'h3d16c6a3 /* (2, 25, 28) */,
  32'h3d21c128 /* (30, 21, 28) */,
  32'h3d41fb9f /* (26, 21, 28) */,
  32'h3d92b699 /* (22, 21, 28) */,
  32'h3ddc0819 /* (18, 21, 28) */,
  32'h3ddc0819 /* (14, 21, 28) */,
  32'h3d92b699 /* (10, 21, 28) */,
  32'h3d41fb9f /* (6, 21, 28) */,
  32'h3d21c128 /* (2, 21, 28) */,
  32'h3d2d6bba /* (30, 17, 28) */,
  32'h3d61b1de /* (26, 17, 28) */,
  32'h3dbdf4f8 /* (22, 17, 28) */,
  32'h3e1c2ca1 /* (18, 17, 28) */,
  32'h3e1c2ca1 /* (14, 17, 28) */,
  32'h3dbdf4f8 /* (10, 17, 28) */,
  32'h3d61b1de /* (6, 17, 28) */,
  32'h3d2d6bba /* (2, 17, 28) */,
  32'h3d3217f4 /* (30, 13, 28) */,
  32'h3d601ae9 /* (26, 13, 28) */,
  32'h3db40e50 /* (22, 13, 28) */,
  32'h3e0de89e /* (18, 13, 28) */,
  32'h3e0de89e /* (14, 13, 28) */,
  32'h3db40e50 /* (10, 13, 28) */,
  32'h3d601ae9 /* (6, 13, 28) */,
  32'h3d3217f4 /* (2, 13, 28) */,
  32'h3d14de35 /* (30, 9, 28) */,
  32'h3d2657dd /* (26, 9, 28) */,
  32'h3d68b7a2 /* (22, 9, 28) */,
  32'h3da4db8a /* (18, 9, 28) */,
  32'h3da4db8a /* (14, 9, 28) */,
  32'h3d68b7a2 /* (10, 9, 28) */,
  32'h3d2657dd /* (6, 9, 28) */,
  32'h3d14de35 /* (2, 9, 28) */,
  32'h3d2d8e0e /* (30, 5, 28) */,
  32'h3d153e19 /* (26, 5, 28) */,
  32'h3d28e3b2 /* (22, 5, 28) */,
  32'h3d53bb31 /* (18, 5, 28) */,
  32'h3d53bb31 /* (14, 5, 28) */,
  32'h3d28e3b2 /* (10, 5, 28) */,
  32'h3d153e19 /* (6, 5, 28) */,
  32'h3d2d8e0e /* (2, 5, 28) */,
  32'h3d8b1391 /* (30, 1, 28) */,
  32'h3d222a9c /* (26, 1, 28) */,
  32'h3d1839e3 /* (22, 1, 28) */,
  32'h3d303352 /* (18, 1, 28) */,
  32'h3d303352 /* (14, 1, 28) */,
  32'h3d1839e3 /* (10, 1, 28) */,
  32'h3d222a9c /* (6, 1, 28) */,
  32'h3d8b1391 /* (2, 1, 28) */,
  32'h3d13e9f7 /* (30, 29, 24) */,
  32'h3d19bf4b /* (26, 29, 24) */,
  32'h3d48bc7e /* (22, 29, 24) */,
  32'h3d880501 /* (18, 29, 24) */,
  32'h3d880501 /* (14, 29, 24) */,
  32'h3d48bc7e /* (10, 29, 24) */,
  32'h3d19bf4b /* (6, 29, 24) */,
  32'h3d13e9f7 /* (2, 29, 24) */,
  32'h3d1d59b0 /* (30, 25, 24) */,
  32'h3d35cd98 /* (26, 25, 24) */,
  32'h3d83c517 /* (22, 25, 24) */,
  32'h3dbf672f /* (18, 25, 24) */,
  32'h3dbf672f /* (14, 25, 24) */,
  32'h3d83c517 /* (10, 25, 24) */,
  32'h3d35cd98 /* (6, 25, 24) */,
  32'h3d1d59b0 /* (2, 25, 24) */,
  32'h3d558b1c /* (30, 21, 24) */,
  32'h3d865b59 /* (26, 21, 24) */,
  32'h3dd7e578 /* (22, 21, 24) */,
  32'h3e2a27e4 /* (18, 21, 24) */,
  32'h3e2a27e4 /* (14, 21, 24) */,
  32'h3dd7e578 /* (10, 21, 24) */,
  32'h3d865b59 /* (6, 21, 24) */,
  32'h3d558b1c /* (2, 21, 24) */,
  32'h3d804df8 /* (30, 17, 24) */,
  32'h3daa3349 /* (26, 17, 24) */,
  32'h3e135573 /* (22, 17, 24) */,
  32'h3e79034c /* (18, 17, 24) */,
  32'h3e79034c /* (14, 17, 24) */,
  32'h3e135573 /* (10, 17, 24) */,
  32'h3daa3349 /* (6, 17, 24) */,
  32'h3d804df8 /* (2, 17, 24) */,
  32'h3d7b52f8 /* (30, 13, 24) */,
  32'h3da2e7a9 /* (26, 13, 24) */,
  32'h3e085939 /* (22, 13, 24) */,
  32'h3e5f05ce /* (18, 13, 24) */,
  32'h3e5f05ce /* (14, 13, 24) */,
  32'h3e085939 /* (10, 13, 24) */,
  32'h3da2e7a9 /* (6, 13, 24) */,
  32'h3d7b52f8 /* (2, 13, 24) */,
  32'h3d3291f6 /* (30, 9, 24) */,
  32'h3d584c0c /* (26, 9, 24) */,
  32'h3da590e9 /* (22, 9, 24) */,
  32'h3dfaaa60 /* (18, 9, 24) */,
  32'h3dfaaa60 /* (14, 9, 24) */,
  32'h3da590e9 /* (10, 9, 24) */,
  32'h3d584c0c /* (6, 9, 24) */,
  32'h3d3291f6 /* (2, 9, 24) */,
  32'h3d149b5c /* (30, 5, 24) */,
  32'h3d22af34 /* (26, 5, 24) */,
  32'h3d5ef675 /* (22, 5, 24) */,
  32'h3d9bc970 /* (18, 5, 24) */,
  32'h3d9bc970 /* (14, 5, 24) */,
  32'h3d5ef675 /* (10, 5, 24) */,
  32'h3d22af34 /* (6, 5, 24) */,
  32'h3d149b5c /* (2, 5, 24) */,
  32'h3d15ce12 /* (30, 1, 24) */,
  32'h3d169650 /* (26, 1, 24) */,
  32'h3d3f0366 /* (22, 1, 24) */,
  32'h3d7e759f /* (18, 1, 24) */,
  32'h3d7e759f /* (14, 1, 24) */,
  32'h3d3f0366 /* (10, 1, 24) */,
  32'h3d169650 /* (6, 1, 24) */,
  32'h3d15ce12 /* (2, 1, 24) */,
  32'h3d23d587 /* (30, 29, 20) */,
  32'h3d48406d /* (26, 29, 20) */,
  32'h3d9aff71 /* (22, 29, 20) */,
  32'h3decc5e8 /* (18, 29, 20) */,
  32'h3decc5e8 /* (14, 29, 20) */,
  32'h3d9aff71 /* (10, 29, 20) */,
  32'h3d48406d /* (6, 29, 20) */,
  32'h3d23d587 /* (2, 29, 20) */,
  32'h3d530d8e /* (30, 25, 20) */,
  32'h3d859348 /* (26, 25, 20) */,
  32'h3dd85675 /* (22, 25, 20) */,
  32'h3e2baf50 /* (18, 25, 20) */,
  32'h3e2baf50 /* (14, 25, 20) */,
  32'h3dd85675 /* (10, 25, 20) */,
  32'h3d859348 /* (6, 25, 20) */,
  32'h3d530d8e /* (2, 25, 20) */,
  32'h3da96c08 /* (30, 21, 20) */,
  32'h3ddec971 /* (26, 21, 20) */,
  32'h3e3e5baf /* (22, 21, 20) */,
  32'h3e9ecc49 /* (18, 21, 20) */,
  32'h3e9ecc49 /* (14, 21, 20) */,
  32'h3e3e5baf /* (10, 21, 20) */,
  32'h3ddec971 /* (6, 21, 20) */,
  32'h3da96c08 /* (2, 21, 20) */,
  32'h3de39dff /* (30, 17, 20) */,
  32'h3e1a3a56 /* (26, 17, 20) */,
  32'h3e89fde5 /* (22, 17, 20) */,
  32'h3ef15f91 /* (18, 17, 20) */,
  32'h3ef15f91 /* (14, 17, 20) */,
  32'h3e89fde5 /* (10, 17, 20) */,
  32'h3e1a3a56 /* (6, 17, 20) */,
  32'h3de39dff /* (2, 17, 20) */,
  32'h3dd42d31 /* (30, 13, 20) */,
  32'h3e0dc95f /* (26, 13, 20) */,
  32'h3e7848b5 /* (22, 13, 20) */,
  32'h3ed441df /* (18, 13, 20) */,
  32'h3ed441df /* (14, 13, 20) */,
  32'h3e7848b5 /* (10, 13, 20) */,
  32'h3e0dc95f /* (6, 13, 20) */,
  32'h3dd42d31 /* (2, 13, 20) */,
  32'h3d833332 /* (30, 9, 20) */,
  32'h3da96159 /* (26, 9, 20) */,
  32'h3e0cf021 /* (22, 9, 20) */,
  32'h3e654448 /* (18, 9, 20) */,
  32'h3e654448 /* (14, 9, 20) */,
  32'h3e0cf021 /* (10, 9, 20) */,
  32'h3da96159 /* (6, 9, 20) */,
  32'h3d833332 /* (2, 9, 20) */,
  32'h3d346b02 /* (30, 5, 20) */,
  32'h3d6007ad /* (26, 5, 20) */,
  32'h3db0e528 /* (22, 5, 20) */,
  32'h3e095be4 /* (18, 5, 20) */,
  32'h3e095be4 /* (14, 5, 20) */,
  32'h3db0e528 /* (10, 5, 20) */,
  32'h3d6007ad /* (6, 5, 20) */,
  32'h3d346b02 /* (2, 5, 20) */,
  32'h3d1cac31 /* (30, 1, 20) */,
  32'h3d3dc5f0 /* (26, 1, 20) */,
  32'h3d91435f /* (22, 1, 20) */,
  32'h3ddbed5a /* (18, 1, 20) */,
  32'h3ddbed5a /* (14, 1, 20) */,
  32'h3d91435f /* (10, 1, 20) */,
  32'h3d3dc5f0 /* (6, 1, 20) */,
  32'h3d1cac31 /* (2, 1, 20) */,
  32'h3d13661d /* (30, 29, 16) */,
  32'h3d41d3ae /* (26, 29, 16) */,
  32'h3da59d10 /* (22, 29, 16) */,
  32'h3e0a27e7 /* (18, 29, 16) */,
  32'h3e0a27e7 /* (14, 29, 16) */,
  32'h3da59d10 /* (10, 29, 16) */,
  32'h3d41d3ae /* (6, 29, 16) */,
  32'h3d13661d /* (2, 29, 16) */,
  32'h3d4f6a6e /* (30, 25, 16) */,
  32'h3d8a46e7 /* (26, 25, 16) */,
  32'h3df142da /* (22, 25, 16) */,
  32'h3e4d7ce8 /* (18, 25, 16) */,
  32'h3e4d7ce8 /* (14, 25, 16) */,
  32'h3df142da /* (10, 25, 16) */,
  32'h3d8a46e7 /* (6, 25, 16) */,
  32'h3d4f6a6e /* (2, 25, 16) */,
  32'h3db86416 /* (30, 21, 16) */,
  32'h3dfa4afe /* (26, 21, 16) */,
  32'h3e60898b /* (22, 21, 16) */,
  32'h3ec4f0a1 /* (18, 21, 16) */,
  32'h3ec4f0a1 /* (14, 21, 16) */,
  32'h3e60898b /* (10, 21, 16) */,
  32'h3dfa4afe /* (6, 21, 16) */,
  32'h3db86416 /* (2, 21, 16) */,
  32'h3e06ec2e /* (30, 17, 16) */,
  32'h3e3a3d1a /* (26, 17, 16) */,
  32'h3eabb572 /* (22, 17, 16) */,
  32'h3f1b42bd /* (18, 17, 16) */,
  32'h3f1b42bd /* (14, 17, 16) */,
  32'h3eabb572 /* (10, 17, 16) */,
  32'h3e3a3d1a /* (6, 17, 16) */,
  32'h3e06ec2e /* (2, 17, 16) */,
  32'h3df1ae3d /* (30, 13, 16) */,
  32'h3e2576a9 /* (26, 13, 16) */,
  32'h3e968a40 /* (22, 13, 16) */,
  32'h3f06176f /* (18, 13, 16) */,
  32'h3f06176f /* (14, 13, 16) */,
  32'h3e968a40 /* (10, 13, 16) */,
  32'h3e2576a9 /* (6, 13, 16) */,
  32'h3df1ae3d /* (2, 13, 16) */,
  32'h3d87d16b /* (30, 9, 16) */,
  32'h3db6b309 /* (26, 9, 16) */,
  32'h3e21930d /* (22, 9, 16) */,
  32'h3e8b9344 /* (18, 9, 16) */,
  32'h3e8b9344 /* (14, 9, 16) */,
  32'h3e21930d /* (10, 9, 16) */,
  32'h3db6b309 /* (6, 9, 16) */,
  32'h3d87d16b /* (2, 9, 16) */,
  32'h3d28d1e5 /* (30, 5, 16) */,
  32'h3d5f53fb /* (26, 5, 16) */,
  32'h3dc0863e /* (22, 5, 16) */,
  32'h3e2205a1 /* (18, 5, 16) */,
  32'h3e2205a1 /* (14, 5, 16) */,
  32'h3dc0863e /* (10, 5, 16) */,
  32'h3d5f53fb /* (6, 5, 16) */,
  32'h3d28d1e5 /* (2, 5, 16) */,
  32'h3d09dfab /* (30, 1, 16) */,
  32'h3d34b66a /* (26, 1, 16) */,
  32'h3d99ac24 /* (22, 1, 16) */,
  32'h3dff32bb /* (18, 1, 16) */,
  32'h3dff32bb /* (14, 1, 16) */,
  32'h3d99ac24 /* (10, 1, 16) */,
  32'h3d34b66a /* (6, 1, 16) */,
  32'h3d09dfab /* (2, 1, 16) */,
  32'h3d23d587 /* (30, 29, 12) */,
  32'h3d48406d /* (26, 29, 12) */,
  32'h3d9aff71 /* (22, 29, 12) */,
  32'h3decc5e8 /* (18, 29, 12) */,
  32'h3decc5e8 /* (14, 29, 12) */,
  32'h3d9aff71 /* (10, 29, 12) */,
  32'h3d48406d /* (6, 29, 12) */,
  32'h3d23d587 /* (2, 29, 12) */,
  32'h3d530d8e /* (30, 25, 12) */,
  32'h3d859348 /* (26, 25, 12) */,
  32'h3dd85675 /* (22, 25, 12) */,
  32'h3e2baf50 /* (18, 25, 12) */,
  32'h3e2baf50 /* (14, 25, 12) */,
  32'h3dd85675 /* (10, 25, 12) */,
  32'h3d859348 /* (6, 25, 12) */,
  32'h3d530d8e /* (2, 25, 12) */,
  32'h3da96c08 /* (30, 21, 12) */,
  32'h3ddec971 /* (26, 21, 12) */,
  32'h3e3e5baf /* (22, 21, 12) */,
  32'h3e9ecc49 /* (18, 21, 12) */,
  32'h3e9ecc49 /* (14, 21, 12) */,
  32'h3e3e5baf /* (10, 21, 12) */,
  32'h3ddec971 /* (6, 21, 12) */,
  32'h3da96c08 /* (2, 21, 12) */,
  32'h3de39dff /* (30, 17, 12) */,
  32'h3e1a3a56 /* (26, 17, 12) */,
  32'h3e89fde5 /* (22, 17, 12) */,
  32'h3ef15f91 /* (18, 17, 12) */,
  32'h3ef15f91 /* (14, 17, 12) */,
  32'h3e89fde5 /* (10, 17, 12) */,
  32'h3e1a3a56 /* (6, 17, 12) */,
  32'h3de39dff /* (2, 17, 12) */,
  32'h3dd42d31 /* (30, 13, 12) */,
  32'h3e0dc95f /* (26, 13, 12) */,
  32'h3e7848b5 /* (22, 13, 12) */,
  32'h3ed441df /* (18, 13, 12) */,
  32'h3ed441df /* (14, 13, 12) */,
  32'h3e7848b5 /* (10, 13, 12) */,
  32'h3e0dc95f /* (6, 13, 12) */,
  32'h3dd42d31 /* (2, 13, 12) */,
  32'h3d833332 /* (30, 9, 12) */,
  32'h3da96159 /* (26, 9, 12) */,
  32'h3e0cf021 /* (22, 9, 12) */,
  32'h3e654448 /* (18, 9, 12) */,
  32'h3e654448 /* (14, 9, 12) */,
  32'h3e0cf021 /* (10, 9, 12) */,
  32'h3da96159 /* (6, 9, 12) */,
  32'h3d833332 /* (2, 9, 12) */,
  32'h3d346b02 /* (30, 5, 12) */,
  32'h3d6007ad /* (26, 5, 12) */,
  32'h3db0e528 /* (22, 5, 12) */,
  32'h3e095be4 /* (18, 5, 12) */,
  32'h3e095be4 /* (14, 5, 12) */,
  32'h3db0e528 /* (10, 5, 12) */,
  32'h3d6007ad /* (6, 5, 12) */,
  32'h3d346b02 /* (2, 5, 12) */,
  32'h3d1cac31 /* (30, 1, 12) */,
  32'h3d3dc5f0 /* (26, 1, 12) */,
  32'h3d91435f /* (22, 1, 12) */,
  32'h3ddbed5a /* (18, 1, 12) */,
  32'h3ddbed5a /* (14, 1, 12) */,
  32'h3d91435f /* (10, 1, 12) */,
  32'h3d3dc5f0 /* (6, 1, 12) */,
  32'h3d1cac31 /* (2, 1, 12) */,
  32'h3d13e9f7 /* (30, 29, 8) */,
  32'h3d19bf4b /* (26, 29, 8) */,
  32'h3d48bc7e /* (22, 29, 8) */,
  32'h3d880501 /* (18, 29, 8) */,
  32'h3d880501 /* (14, 29, 8) */,
  32'h3d48bc7e /* (10, 29, 8) */,
  32'h3d19bf4b /* (6, 29, 8) */,
  32'h3d13e9f7 /* (2, 29, 8) */,
  32'h3d1d59b0 /* (30, 25, 8) */,
  32'h3d35cd98 /* (26, 25, 8) */,
  32'h3d83c517 /* (22, 25, 8) */,
  32'h3dbf672f /* (18, 25, 8) */,
  32'h3dbf672f /* (14, 25, 8) */,
  32'h3d83c517 /* (10, 25, 8) */,
  32'h3d35cd98 /* (6, 25, 8) */,
  32'h3d1d59b0 /* (2, 25, 8) */,
  32'h3d558b1c /* (30, 21, 8) */,
  32'h3d865b59 /* (26, 21, 8) */,
  32'h3dd7e578 /* (22, 21, 8) */,
  32'h3e2a27e4 /* (18, 21, 8) */,
  32'h3e2a27e4 /* (14, 21, 8) */,
  32'h3dd7e578 /* (10, 21, 8) */,
  32'h3d865b59 /* (6, 21, 8) */,
  32'h3d558b1c /* (2, 21, 8) */,
  32'h3d804df8 /* (30, 17, 8) */,
  32'h3daa3349 /* (26, 17, 8) */,
  32'h3e135573 /* (22, 17, 8) */,
  32'h3e79034c /* (18, 17, 8) */,
  32'h3e79034c /* (14, 17, 8) */,
  32'h3e135573 /* (10, 17, 8) */,
  32'h3daa3349 /* (6, 17, 8) */,
  32'h3d804df8 /* (2, 17, 8) */,
  32'h3d7b52f8 /* (30, 13, 8) */,
  32'h3da2e7a9 /* (26, 13, 8) */,
  32'h3e085939 /* (22, 13, 8) */,
  32'h3e5f05ce /* (18, 13, 8) */,
  32'h3e5f05ce /* (14, 13, 8) */,
  32'h3e085939 /* (10, 13, 8) */,
  32'h3da2e7a9 /* (6, 13, 8) */,
  32'h3d7b52f8 /* (2, 13, 8) */,
  32'h3d3291f6 /* (30, 9, 8) */,
  32'h3d584c0c /* (26, 9, 8) */,
  32'h3da590e9 /* (22, 9, 8) */,
  32'h3dfaaa60 /* (18, 9, 8) */,
  32'h3dfaaa60 /* (14, 9, 8) */,
  32'h3da590e9 /* (10, 9, 8) */,
  32'h3d584c0c /* (6, 9, 8) */,
  32'h3d3291f6 /* (2, 9, 8) */,
  32'h3d149b5c /* (30, 5, 8) */,
  32'h3d22af34 /* (26, 5, 8) */,
  32'h3d5ef675 /* (22, 5, 8) */,
  32'h3d9bc970 /* (18, 5, 8) */,
  32'h3d9bc970 /* (14, 5, 8) */,
  32'h3d5ef675 /* (10, 5, 8) */,
  32'h3d22af34 /* (6, 5, 8) */,
  32'h3d149b5c /* (2, 5, 8) */,
  32'h3d15ce12 /* (30, 1, 8) */,
  32'h3d169650 /* (26, 1, 8) */,
  32'h3d3f0366 /* (22, 1, 8) */,
  32'h3d7e759f /* (18, 1, 8) */,
  32'h3d7e759f /* (14, 1, 8) */,
  32'h3d3f0366 /* (10, 1, 8) */,
  32'h3d169650 /* (6, 1, 8) */,
  32'h3d15ce12 /* (2, 1, 8) */,
  32'h3d5defd3 /* (30, 29, 4) */,
  32'h3d1b3fff /* (26, 29, 4) */,
  32'h3d1cff11 /* (22, 29, 4) */,
  32'h3d3b1e93 /* (18, 29, 4) */,
  32'h3d3b1e93 /* (14, 29, 4) */,
  32'h3d1cff11 /* (10, 29, 4) */,
  32'h3d1b3fff /* (6, 29, 4) */,
  32'h3d5defd3 /* (2, 29, 4) */,
  32'h3d16c6a3 /* (30, 25, 4) */,
  32'h3d17902e /* (26, 25, 4) */,
  32'h3d404057 /* (22, 25, 4) */,
  32'h3d800deb /* (18, 25, 4) */,
  32'h3d800deb /* (14, 25, 4) */,
  32'h3d404057 /* (10, 25, 4) */,
  32'h3d17902e /* (6, 25, 4) */,
  32'h3d16c6a3 /* (2, 25, 4) */,
  32'h3d21c128 /* (30, 21, 4) */,
  32'h3d41fb9f /* (26, 21, 4) */,
  32'h3d92b699 /* (22, 21, 4) */,
  32'h3ddc0819 /* (18, 21, 4) */,
  32'h3ddc0819 /* (14, 21, 4) */,
  32'h3d92b699 /* (10, 21, 4) */,
  32'h3d41fb9f /* (6, 21, 4) */,
  32'h3d21c128 /* (2, 21, 4) */,
  32'h3d2d6bba /* (30, 17, 4) */,
  32'h3d61b1de /* (26, 17, 4) */,
  32'h3dbdf4f8 /* (22, 17, 4) */,
  32'h3e1c2ca1 /* (18, 17, 4) */,
  32'h3e1c2ca1 /* (14, 17, 4) */,
  32'h3dbdf4f8 /* (10, 17, 4) */,
  32'h3d61b1de /* (6, 17, 4) */,
  32'h3d2d6bba /* (2, 17, 4) */,
  32'h3d3217f4 /* (30, 13, 4) */,
  32'h3d601ae9 /* (26, 13, 4) */,
  32'h3db40e50 /* (22, 13, 4) */,
  32'h3e0de89e /* (18, 13, 4) */,
  32'h3e0de89e /* (14, 13, 4) */,
  32'h3db40e50 /* (10, 13, 4) */,
  32'h3d601ae9 /* (6, 13, 4) */,
  32'h3d3217f4 /* (2, 13, 4) */,
  32'h3d14de35 /* (30, 9, 4) */,
  32'h3d2657dd /* (26, 9, 4) */,
  32'h3d68b7a2 /* (22, 9, 4) */,
  32'h3da4db8a /* (18, 9, 4) */,
  32'h3da4db8a /* (14, 9, 4) */,
  32'h3d68b7a2 /* (10, 9, 4) */,
  32'h3d2657dd /* (6, 9, 4) */,
  32'h3d14de35 /* (2, 9, 4) */,
  32'h3d2d8e0e /* (30, 5, 4) */,
  32'h3d153e19 /* (26, 5, 4) */,
  32'h3d28e3b2 /* (22, 5, 4) */,
  32'h3d53bb31 /* (18, 5, 4) */,
  32'h3d53bb31 /* (14, 5, 4) */,
  32'h3d28e3b2 /* (10, 5, 4) */,
  32'h3d153e19 /* (6, 5, 4) */,
  32'h3d2d8e0e /* (2, 5, 4) */,
  32'h3d8b1391 /* (30, 1, 4) */,
  32'h3d222a9c /* (26, 1, 4) */,
  32'h3d1839e3 /* (22, 1, 4) */,
  32'h3d303352 /* (18, 1, 4) */,
  32'h3d303352 /* (14, 1, 4) */,
  32'h3d1839e3 /* (10, 1, 4) */,
  32'h3d222a9c /* (6, 1, 4) */,
  32'h3d8b1391 /* (2, 1, 4) */,
  32'h3dcbea25 /* (30, 29, 0) */,
  32'h3d2d5b95 /* (26, 29, 0) */,
  32'h3d144f19 /* (22, 29, 0) */,
  32'h3d262b6e /* (18, 29, 0) */,
  32'h3d262b6e /* (14, 29, 0) */,
  32'h3d144f19 /* (10, 29, 0) */,
  32'h3d2d5b95 /* (6, 29, 0) */,
  32'h3dcbea25 /* (2, 29, 0) */,
  32'h3d21b235 /* (30, 25, 0) */,
  32'h3d1459dd /* (26, 25, 0) */,
  32'h3d2f5f5a /* (22, 25, 0) */,
  32'h3d60bf24 /* (18, 25, 0) */,
  32'h3d60bf24 /* (14, 25, 0) */,
  32'h3d2f5f5a /* (10, 25, 0) */,
  32'h3d1459dd /* (6, 25, 0) */,
  32'h3d21b235 /* (2, 25, 0) */,
  32'h3d164ce1 /* (30, 21, 0) */,
  32'h3d3013e2 /* (26, 21, 0) */,
  32'h3d819abc /* (22, 21, 0) */,
  32'h3dbe661f /* (18, 21, 0) */,
  32'h3dbe661f /* (14, 21, 0) */,
  32'h3d819abc /* (10, 21, 0) */,
  32'h3d3013e2 /* (6, 21, 0) */,
  32'h3d164ce1 /* (2, 21, 0) */,
  32'h3d18d610 /* (30, 17, 0) */,
  32'h3d455011 /* (26, 17, 0) */,
  32'h3da42e1b /* (22, 17, 0) */,
  32'h3e05899d /* (18, 17, 0) */,
  32'h3e05899d /* (14, 17, 0) */,
  32'h3da42e1b /* (10, 17, 0) */,
  32'h3d455011 /* (6, 17, 0) */,
  32'h3d18d610 /* (2, 17, 0) */,
  32'h3d2045b1 /* (30, 13, 0) */,
  32'h3d4703b2 /* (26, 13, 0) */,
  32'h3d9d248b /* (22, 13, 0) */,
  32'h3df40add /* (18, 13, 0) */,
  32'h3df40add /* (14, 13, 0) */,
  32'h3d9d248b /* (10, 13, 0) */,
  32'h3d4703b2 /* (6, 13, 0) */,
  32'h3d2045b1 /* (2, 13, 0) */,
  32'h3d11b684 /* (30, 9, 0) */,
  32'h3d1bc36a /* (26, 9, 0) */,
  32'h3d50a575 /* (22, 9, 0) */,
  32'h3d8fa52c /* (18, 9, 0) */,
  32'h3d8fa52c /* (14, 9, 0) */,
  32'h3d50a575 /* (10, 9, 0) */,
  32'h3d1bc36a /* (6, 9, 0) */,
  32'h3d11b684 /* (2, 9, 0) */,
  32'h3d5dd7d1 /* (30, 5, 0) */,
  32'h3d1b2f33 /* (26, 5, 0) */,
  32'h3d1cee15 /* (22, 5, 0) */,
  32'h3d3b0a55 /* (18, 5, 0) */,
  32'h3d3b0a55 /* (14, 5, 0) */,
  32'h3d1cee15 /* (10, 5, 0) */,
  32'h3d1b2f33 /* (6, 5, 0) */,
  32'h3d5dd7d1 /* (2, 5, 0) */,
  32'h3e709592 /* (30, 1, 0) */,
  32'h3d3f59b8 /* (26, 1, 0) */,
  32'h3d1142bb /* (22, 1, 0) */,
  32'h3d1ceee6 /* (18, 1, 0) */,
  32'h3d1ceee6 /* (14, 1, 0) */,
  32'h3d1142bb /* (10, 1, 0) */,
  32'h3d3f59b8 /* (6, 1, 0) */,
  32'h3e709592 /* (2, 1, 0) */,
  32'h3d4920d0 /* (29, 29, 28) */,
  32'h3d155fa4 /* (25, 29, 28) */,
  32'h3d25fa09 /* (21, 29, 28) */,
  32'h3d349293 /* (17, 29, 28) */,
  32'h3d385879 /* (13, 29, 28) */,
  32'h3d16b5b2 /* (9, 29, 28) */,
  32'h3d25f5ce /* (5, 29, 28) */,
  32'h3d6eb36b /* (1, 29, 28) */,
  32'h3d155fa4 /* (29, 25, 28) */,
  32'h3d1cbb18 /* (25, 25, 28) */,
  32'h3d52976b /* (21, 25, 28) */,
  32'h3d7b9f11 /* (17, 25, 28) */,
  32'h3d770afc /* (13, 25, 28) */,
  32'h3d30de15 /* (9, 25, 28) */,
  32'h3d1508af /* (5, 25, 28) */,
  32'h3d17ff6b /* (1, 25, 28) */,
  32'h3d25fa09 /* (29, 21, 28) */,
  32'h3d52976b /* (25, 21, 28) */,
  32'h3da66ad4 /* (21, 21, 28) */,
  32'h3ddcf428 /* (17, 21, 28) */,
  32'h3dcf13a3 /* (13, 21, 28) */,
  32'h3d81d711 /* (9, 21, 28) */,
  32'h3d358341 /* (5, 21, 28) */,
  32'h3d1f5dc3 /* (1, 21, 28) */,
  32'h3d349293 /* (29, 17, 28) */,
  32'h3d7b9f11 /* (25, 17, 28) */,
  32'h3ddcf428 /* (21, 17, 28) */,
  32'h3e1fe07e /* (17, 17, 28) */,
  32'h3e0ff4ce /* (13, 17, 28) */,
  32'h3da3c1ed /* (9, 17, 28) */,
  32'h3d4def9b /* (5, 17, 28) */,
  32'h3d294c4b /* (1, 17, 28) */,
  32'h3d385879 /* (29, 13, 28) */,
  32'h3d770afc /* (25, 13, 28) */,
  32'h3dcf13a3 /* (21, 13, 28) */,
  32'h3e0ff4ce /* (17, 13, 28) */,
  32'h3e0415cb /* (13, 13, 28) */,
  32'h3d9d0afa /* (9, 13, 28) */,
  32'h3d4ea6a0 /* (5, 13, 28) */,
  32'h3d2e802a /* (1, 13, 28) */,
  32'h3d16b5b2 /* (29, 9, 28) */,
  32'h3d30de15 /* (25, 9, 28) */,
  32'h3d81d711 /* (21, 9, 28) */,
  32'h3da3c1ed /* (17, 9, 28) */,
  32'h3d9d0afa /* (13, 9, 28) */,
  32'h3d51a9d2 /* (9, 9, 28) */,
  32'h3d1ee50b /* (5, 9, 28) */,
  32'h3d13f199 /* (1, 9, 28) */,
  32'h3d25f5ce /* (29, 5, 28) */,
  32'h3d1508af /* (25, 5, 28) */,
  32'h3d358341 /* (21, 5, 28) */,
  32'h3d4def9b /* (17, 5, 28) */,
  32'h3d4ea6a0 /* (13, 5, 28) */,
  32'h3d1ee50b /* (9, 5, 28) */,
  32'h3d189061 /* (5, 5, 28) */,
  32'h3d334ee4 /* (1, 5, 28) */,
  32'h3d6eb36b /* (29, 1, 28) */,
  32'h3d17ff6b /* (25, 1, 28) */,
  32'h3d1f5dc3 /* (21, 1, 28) */,
  32'h3d294c4b /* (17, 1, 28) */,
  32'h3d2e802a /* (13, 1, 28) */,
  32'h3d13f199 /* (9, 1, 28) */,
  32'h3d334ee4 /* (5, 1, 28) */,
  32'h3d9c757b /* (1, 1, 28) */,
  32'h3d1392fe /* (29, 29, 24) */,
  32'h3d2054cd /* (25, 29, 24) */,
  32'h3d5d0a38 /* (21, 29, 24) */,
  32'h3d8608f0 /* (17, 29, 24) */,
  32'h3d82c188 /* (13, 29, 24) */,
  32'h3d37919e /* (9, 29, 24) */,
  32'h3d15d660 /* (5, 29, 24) */,
  32'h3d146963 /* (1, 29, 24) */,
  32'h3d2054cd /* (29, 25, 24) */,
  32'h3d432bf1 /* (25, 25, 24) */,
  32'h3d941bce /* (21, 25, 24) */,
  32'h3dbf0444 /* (17, 25, 24) */,
  32'h3db56072 /* (13, 25, 24) */,
  32'h3d6b8b35 /* (9, 25, 24) */,
  32'h3d2bff3e /* (5, 25, 24) */,
  32'h3d1bb8b6 /* (1, 25, 24) */,
  32'h3d5d0a38 /* (29, 21, 24) */,
  32'h3d941bce /* (25, 21, 24) */,
  32'h3df84bb3 /* (21, 21, 24) */,
  32'h3e2c9c6c /* (17, 21, 24) */,
  32'h3e1e607d /* (13, 21, 24) */,
  32'h3dbc4d73 /* (9, 21, 24) */,
  32'h3d77c8fd /* (5, 21, 24) */,
  32'h3d513c3d /* (1, 21, 24) */,
  32'h3d8608f0 /* (29, 17, 24) */,
  32'h3dbf0444 /* (25, 17, 24) */,
  32'h3e2c9c6c /* (21, 17, 24) */,
  32'h3e803f85 /* (17, 17, 24) */,
  32'h3e640ba2 /* (13, 17, 24) */,
  32'h3dfc30a3 /* (9, 17, 24) */,
  32'h3d9a5b6b /* (5, 17, 24) */,
  32'h3d7a003f /* (1, 17, 24) */,
  32'h3d82c188 /* (29, 13, 24) */,
  32'h3db56072 /* (25, 13, 24) */,
  32'h3e1e607d /* (21, 13, 24) */,
  32'h3e640ba2 /* (17, 13, 24) */,
  32'h3e4dd3dc /* (13, 13, 24) */,
  32'h3deb6b6d /* (9, 13, 24) */,
  32'h3d94d380 /* (5, 13, 24) */,
  32'h3d7573b6 /* (1, 13, 24) */,
  32'h3d37919e /* (29, 9, 24) */,
  32'h3d6b8b35 /* (25, 9, 24) */,
  32'h3dbc4d73 /* (21, 9, 24) */,
  32'h3dfc30a3 /* (17, 9, 24) */,
  32'h3deb6b6d /* (13, 9, 24) */,
  32'h3d921bde /* (9, 9, 24) */,
  32'h3d49c96c /* (5, 9, 24) */,
  32'h3d2fba80 /* (1, 9, 24) */,
  32'h3d15d660 /* (29, 5, 24) */,
  32'h3d2bff3e /* (25, 5, 24) */,
  32'h3d77c8fd /* (21, 5, 24) */,
  32'h3d9a5b6b /* (17, 5, 24) */,
  32'h3d94d380 /* (13, 5, 24) */,
  32'h3d49c96c /* (9, 5, 24) */,
  32'h3d1c4d38 /* (5, 5, 24) */,
  32'h3d1412fd /* (1, 5, 24) */,
  32'h3d146963 /* (29, 1, 24) */,
  32'h3d1bb8b6 /* (25, 1, 24) */,
  32'h3d513c3d /* (21, 1, 24) */,
  32'h3d7a003f /* (17, 1, 24) */,
  32'h3d7573b6 /* (13, 1, 24) */,
  32'h3d2fba80 /* (9, 1, 24) */,
  32'h3d1412fd /* (5, 1, 24) */,
  32'h3d1704d7 /* (1, 1, 24) */,
  32'h3d28b308 /* (29, 29, 20) */,
  32'h3d5ab0e1 /* (25, 29, 20) */,
  32'h3db0b965 /* (21, 29, 20) */,
  32'h3deea44d /* (17, 29, 20) */,
  32'h3dddef48 /* (13, 29, 20) */,
  32'h3d886b82 /* (9, 29, 20) */,
  32'h3d3a4ebb /* (5, 29, 20) */,
  32'h3d210eee /* (1, 29, 20) */,
  32'h3d5ab0e1 /* (29, 25, 20) */,
  32'h3d938890 /* (25, 25, 20) */,
  32'h3df94537 /* (21, 25, 20) */,
  32'h3e2e6a71 /* (17, 25, 20) */,
  32'h3e1f8cbf /* (13, 25, 20) */,
  32'h3dbc51f9 /* (9, 25, 20) */,
  32'h3d75e4d4 /* (5, 25, 20) */,
  32'h3d4ea8e5 /* (1, 25, 20) */,
  32'h3db0b965 /* (29, 21, 20) */,
  32'h3df94537 /* (25, 21, 20) */,
  32'h3e5e44ac /* (21, 21, 20) */,
  32'h3ea31756 /* (17, 21, 20) */,
  32'h3e91dfe2 /* (13, 21, 20) */,
  32'h3e23781b /* (9, 21, 20) */,
  32'h3dca9d53 /* (5, 21, 20) */,
  32'h3da53628 /* (1, 21, 20) */,
  32'h3deea44d /* (29, 17, 20) */,
  32'h3e2e6a71 /* (25, 17, 20) */,
  32'h3ea31756 /* (21, 17, 20) */,
  32'h3efaa119 /* (17, 17, 20) */,
  32'h3edb3822 /* (13, 17, 20) */,
  32'h3e6a25fd /* (9, 17, 20) */,
  32'h3e0ae903 /* (5, 17, 20) */,
  32'h3ddd43c2 /* (1, 17, 20) */,
  32'h3dddef48 /* (29, 13, 20) */,
  32'h3e1f8cbf /* (25, 13, 20) */,
  32'h3e91dfe2 /* (21, 13, 20) */,
  32'h3edb3822 /* (17, 13, 20) */,
  32'h3ec1d890 /* (13, 13, 20) */,
  32'h3e53dc51 /* (9, 13, 20) */,
  32'h3e00477d /* (5, 13, 20) */,
  32'h3dce8d02 /* (1, 13, 20) */,
  32'h3d886b82 /* (29, 9, 20) */,
  32'h3dbc51f9 /* (25, 9, 20) */,
  32'h3e23781b /* (21, 9, 20) */,
  32'h3e6a25fd /* (17, 9, 20) */,
  32'h3e53dc51 /* (13, 9, 20) */,
  32'h3df3b4f2 /* (9, 9, 20) */,
  32'h3d9af1c2 /* (5, 9, 20) */,
  32'h3d803124 /* (1, 9, 20) */,
  32'h3d3a4ebb /* (29, 5, 20) */,
  32'h3d75e4d4 /* (25, 5, 20) */,
  32'h3dca9d53 /* (21, 5, 20) */,
  32'h3e0ae903 /* (17, 5, 20) */,
  32'h3e00477d /* (13, 5, 20) */,
  32'h3d9af1c2 /* (9, 5, 20) */,
  32'h3d4f6dfc /* (5, 5, 20) */,
  32'h3d310ad3 /* (1, 5, 20) */,
  32'h3d210eee /* (29, 1, 20) */,
  32'h3d4ea8e5 /* (25, 1, 20) */,
  32'h3da53628 /* (21, 1, 20) */,
  32'h3ddd43c2 /* (17, 1, 20) */,
  32'h3dce8d02 /* (13, 1, 20) */,
  32'h3d803124 /* (9, 1, 20) */,
  32'h3d310ad3 /* (5, 1, 20) */,
  32'h3d1a2df1 /* (1, 1, 20) */,
  32'h3d19c07a /* (29, 29, 16) */,
  32'h3d58de26 /* (25, 29, 16) */,
  32'h3dc1602b /* (21, 29, 16) */,
  32'h3e0de417 /* (17, 29, 16) */,
  32'h3dfdd31f /* (13, 29, 16) */,
  32'h3d8e3848 /* (9, 29, 16) */,
  32'h3d3046d8 /* (5, 29, 16) */,
  32'h3d0fbc59 /* (1, 29, 16) */,
  32'h3d58de26 /* (29, 25, 16) */,
  32'h3d9b7830 /* (25, 25, 16) */,
  32'h3e0d9cf0 /* (21, 25, 16) */,
  32'h3e540b9b /* (17, 25, 16) */,
  32'h3e3bd4ee /* (13, 25, 16) */,
  32'h3dce1075 /* (9, 25, 16) */,
  32'h3d7a662c /* (5, 25, 16) */,
  32'h3d49f75a /* (1, 25, 16) */,
  32'h3dc1602b /* (29, 21, 16) */,
  32'h3e0d9cf0 /* (25, 21, 16) */,
  32'h3e84c8e0 /* (21, 21, 16) */,
  32'h3ecca1ac /* (17, 21, 16) */,
  32'h3eb2bd2a /* (13, 21, 16) */,
  32'h3e3e5da7 /* (9, 21, 16) */,
  32'h3de14ffa /* (5, 21, 16) */,
  32'h3db336e0 /* (1, 21, 16) */,
  32'h3e0de417 /* (29, 17, 16) */,
  32'h3e540b9b /* (25, 17, 16) */,
  32'h3ecca1ac /* (21, 17, 16) */,
  32'h3f2286f8 /* (17, 17, 16) */,
  32'h3f0bd969 /* (13, 17, 16) */,
  32'h3e908107 /* (9, 17, 16) */,
  32'h3e26bbbb /* (5, 17, 16) */,
  32'h3e02e976 /* (1, 17, 16) */,
  32'h3dfdd31f /* (29, 13, 16) */,
  32'h3e3bd4ee /* (25, 13, 16) */,
  32'h3eb2bd2a /* (21, 13, 16) */,
  32'h3f0bd969 /* (17, 13, 16) */,
  32'h3ef27895 /* (13, 13, 16) */,
  32'h3e7e4b9d /* (9, 13, 16) */,
  32'h3e1486b7 /* (5, 13, 16) */,
  32'h3deaafef /* (1, 13, 16) */,
  32'h3d8e3848 /* (29, 9, 16) */,
  32'h3dce1075 /* (25, 9, 16) */,
  32'h3e3e5da7 /* (21, 9, 16) */,
  32'h3e908107 /* (17, 9, 16) */,
  32'h3e7e4b9d /* (13, 9, 16) */,
  32'h3e0981d7 /* (9, 9, 16) */,
  32'h3da4f2f4 /* (5, 9, 16) */,
  32'h3d8420c9 /* (1, 9, 16) */,
  32'h3d3046d8 /* (29, 5, 16) */,
  32'h3d7a662c /* (25, 5, 16) */,
  32'h3de14ffa /* (21, 5, 16) */,
  32'h3e26bbbb /* (17, 5, 16) */,
  32'h3e1486b7 /* (13, 5, 16) */,
  32'h3da4f2f4 /* (9, 5, 16) */,
  32'h3d4ab7f7 /* (5, 5, 16) */,
  32'h3d24852f /* (1, 5, 16) */,
  32'h3d0fbc59 /* (29, 1, 16) */,
  32'h3d49f75a /* (25, 1, 16) */,
  32'h3db336e0 /* (21, 1, 16) */,
  32'h3e02e976 /* (17, 1, 16) */,
  32'h3deaafef /* (13, 1, 16) */,
  32'h3d8420c9 /* (9, 1, 16) */,
  32'h3d24852f /* (5, 1, 16) */,
  32'h3d067e68 /* (1, 1, 16) */,
  32'h3d28b308 /* (29, 29, 12) */,
  32'h3d5ab0e1 /* (25, 29, 12) */,
  32'h3db0b965 /* (21, 29, 12) */,
  32'h3deea44d /* (17, 29, 12) */,
  32'h3dddef48 /* (13, 29, 12) */,
  32'h3d886b82 /* (9, 29, 12) */,
  32'h3d3a4ebb /* (5, 29, 12) */,
  32'h3d210eee /* (1, 29, 12) */,
  32'h3d5ab0e1 /* (29, 25, 12) */,
  32'h3d938890 /* (25, 25, 12) */,
  32'h3df94537 /* (21, 25, 12) */,
  32'h3e2e6a71 /* (17, 25, 12) */,
  32'h3e1f8cbf /* (13, 25, 12) */,
  32'h3dbc51f9 /* (9, 25, 12) */,
  32'h3d75e4d4 /* (5, 25, 12) */,
  32'h3d4ea8e5 /* (1, 25, 12) */,
  32'h3db0b965 /* (29, 21, 12) */,
  32'h3df94537 /* (25, 21, 12) */,
  32'h3e5e44ac /* (21, 21, 12) */,
  32'h3ea31756 /* (17, 21, 12) */,
  32'h3e91dfe2 /* (13, 21, 12) */,
  32'h3e23781b /* (9, 21, 12) */,
  32'h3dca9d53 /* (5, 21, 12) */,
  32'h3da53628 /* (1, 21, 12) */,
  32'h3deea44d /* (29, 17, 12) */,
  32'h3e2e6a71 /* (25, 17, 12) */,
  32'h3ea31756 /* (21, 17, 12) */,
  32'h3efaa119 /* (17, 17, 12) */,
  32'h3edb3822 /* (13, 17, 12) */,
  32'h3e6a25fd /* (9, 17, 12) */,
  32'h3e0ae903 /* (5, 17, 12) */,
  32'h3ddd43c2 /* (1, 17, 12) */,
  32'h3dddef48 /* (29, 13, 12) */,
  32'h3e1f8cbf /* (25, 13, 12) */,
  32'h3e91dfe2 /* (21, 13, 12) */,
  32'h3edb3822 /* (17, 13, 12) */,
  32'h3ec1d890 /* (13, 13, 12) */,
  32'h3e53dc51 /* (9, 13, 12) */,
  32'h3e00477d /* (5, 13, 12) */,
  32'h3dce8d02 /* (1, 13, 12) */,
  32'h3d886b82 /* (29, 9, 12) */,
  32'h3dbc51f9 /* (25, 9, 12) */,
  32'h3e23781b /* (21, 9, 12) */,
  32'h3e6a25fd /* (17, 9, 12) */,
  32'h3e53dc51 /* (13, 9, 12) */,
  32'h3df3b4f2 /* (9, 9, 12) */,
  32'h3d9af1c2 /* (5, 9, 12) */,
  32'h3d803124 /* (1, 9, 12) */,
  32'h3d3a4ebb /* (29, 5, 12) */,
  32'h3d75e4d4 /* (25, 5, 12) */,
  32'h3dca9d53 /* (21, 5, 12) */,
  32'h3e0ae903 /* (17, 5, 12) */,
  32'h3e00477d /* (13, 5, 12) */,
  32'h3d9af1c2 /* (9, 5, 12) */,
  32'h3d4f6dfc /* (5, 5, 12) */,
  32'h3d310ad3 /* (1, 5, 12) */,
  32'h3d210eee /* (29, 1, 12) */,
  32'h3d4ea8e5 /* (25, 1, 12) */,
  32'h3da53628 /* (21, 1, 12) */,
  32'h3ddd43c2 /* (17, 1, 12) */,
  32'h3dce8d02 /* (13, 1, 12) */,
  32'h3d803124 /* (9, 1, 12) */,
  32'h3d310ad3 /* (5, 1, 12) */,
  32'h3d1a2df1 /* (1, 1, 12) */,
  32'h3d1392fe /* (29, 29, 8) */,
  32'h3d2054cd /* (25, 29, 8) */,
  32'h3d5d0a38 /* (21, 29, 8) */,
  32'h3d8608f0 /* (17, 29, 8) */,
  32'h3d82c188 /* (13, 29, 8) */,
  32'h3d37919e /* (9, 29, 8) */,
  32'h3d15d660 /* (5, 29, 8) */,
  32'h3d146963 /* (1, 29, 8) */,
  32'h3d2054cd /* (29, 25, 8) */,
  32'h3d432bf1 /* (25, 25, 8) */,
  32'h3d941bce /* (21, 25, 8) */,
  32'h3dbf0444 /* (17, 25, 8) */,
  32'h3db56072 /* (13, 25, 8) */,
  32'h3d6b8b35 /* (9, 25, 8) */,
  32'h3d2bff3e /* (5, 25, 8) */,
  32'h3d1bb8b6 /* (1, 25, 8) */,
  32'h3d5d0a38 /* (29, 21, 8) */,
  32'h3d941bce /* (25, 21, 8) */,
  32'h3df84bb3 /* (21, 21, 8) */,
  32'h3e2c9c6c /* (17, 21, 8) */,
  32'h3e1e607d /* (13, 21, 8) */,
  32'h3dbc4d73 /* (9, 21, 8) */,
  32'h3d77c8fd /* (5, 21, 8) */,
  32'h3d513c3d /* (1, 21, 8) */,
  32'h3d8608f0 /* (29, 17, 8) */,
  32'h3dbf0444 /* (25, 17, 8) */,
  32'h3e2c9c6c /* (21, 17, 8) */,
  32'h3e803f85 /* (17, 17, 8) */,
  32'h3e640ba2 /* (13, 17, 8) */,
  32'h3dfc30a3 /* (9, 17, 8) */,
  32'h3d9a5b6b /* (5, 17, 8) */,
  32'h3d7a003f /* (1, 17, 8) */,
  32'h3d82c188 /* (29, 13, 8) */,
  32'h3db56072 /* (25, 13, 8) */,
  32'h3e1e607d /* (21, 13, 8) */,
  32'h3e640ba2 /* (17, 13, 8) */,
  32'h3e4dd3dc /* (13, 13, 8) */,
  32'h3deb6b6d /* (9, 13, 8) */,
  32'h3d94d380 /* (5, 13, 8) */,
  32'h3d7573b6 /* (1, 13, 8) */,
  32'h3d37919e /* (29, 9, 8) */,
  32'h3d6b8b35 /* (25, 9, 8) */,
  32'h3dbc4d73 /* (21, 9, 8) */,
  32'h3dfc30a3 /* (17, 9, 8) */,
  32'h3deb6b6d /* (13, 9, 8) */,
  32'h3d921bde /* (9, 9, 8) */,
  32'h3d49c96c /* (5, 9, 8) */,
  32'h3d2fba80 /* (1, 9, 8) */,
  32'h3d15d660 /* (29, 5, 8) */,
  32'h3d2bff3e /* (25, 5, 8) */,
  32'h3d77c8fd /* (21, 5, 8) */,
  32'h3d9a5b6b /* (17, 5, 8) */,
  32'h3d94d380 /* (13, 5, 8) */,
  32'h3d49c96c /* (9, 5, 8) */,
  32'h3d1c4d38 /* (5, 5, 8) */,
  32'h3d1412fd /* (1, 5, 8) */,
  32'h3d146963 /* (29, 1, 8) */,
  32'h3d1bb8b6 /* (25, 1, 8) */,
  32'h3d513c3d /* (21, 1, 8) */,
  32'h3d7a003f /* (17, 1, 8) */,
  32'h3d7573b6 /* (13, 1, 8) */,
  32'h3d2fba80 /* (9, 1, 8) */,
  32'h3d1412fd /* (5, 1, 8) */,
  32'h3d1704d7 /* (1, 1, 8) */,
  32'h3d4920d0 /* (29, 29, 4) */,
  32'h3d155fa4 /* (25, 29, 4) */,
  32'h3d25fa09 /* (21, 29, 4) */,
  32'h3d349293 /* (17, 29, 4) */,
  32'h3d385879 /* (13, 29, 4) */,
  32'h3d16b5b2 /* (9, 29, 4) */,
  32'h3d25f5ce /* (5, 29, 4) */,
  32'h3d6eb36b /* (1, 29, 4) */,
  32'h3d155fa4 /* (29, 25, 4) */,
  32'h3d1cbb18 /* (25, 25, 4) */,
  32'h3d52976b /* (21, 25, 4) */,
  32'h3d7b9f11 /* (17, 25, 4) */,
  32'h3d770afc /* (13, 25, 4) */,
  32'h3d30de15 /* (9, 25, 4) */,
  32'h3d1508af /* (5, 25, 4) */,
  32'h3d17ff6b /* (1, 25, 4) */,
  32'h3d25fa09 /* (29, 21, 4) */,
  32'h3d52976b /* (25, 21, 4) */,
  32'h3da66ad4 /* (21, 21, 4) */,
  32'h3ddcf428 /* (17, 21, 4) */,
  32'h3dcf13a3 /* (13, 21, 4) */,
  32'h3d81d711 /* (9, 21, 4) */,
  32'h3d358341 /* (5, 21, 4) */,
  32'h3d1f5dc3 /* (1, 21, 4) */,
  32'h3d349293 /* (29, 17, 4) */,
  32'h3d7b9f11 /* (25, 17, 4) */,
  32'h3ddcf428 /* (21, 17, 4) */,
  32'h3e1fe07e /* (17, 17, 4) */,
  32'h3e0ff4ce /* (13, 17, 4) */,
  32'h3da3c1ed /* (9, 17, 4) */,
  32'h3d4def9b /* (5, 17, 4) */,
  32'h3d294c4b /* (1, 17, 4) */,
  32'h3d385879 /* (29, 13, 4) */,
  32'h3d770afc /* (25, 13, 4) */,
  32'h3dcf13a3 /* (21, 13, 4) */,
  32'h3e0ff4ce /* (17, 13, 4) */,
  32'h3e0415cb /* (13, 13, 4) */,
  32'h3d9d0afa /* (9, 13, 4) */,
  32'h3d4ea6a0 /* (5, 13, 4) */,
  32'h3d2e802a /* (1, 13, 4) */,
  32'h3d16b5b2 /* (29, 9, 4) */,
  32'h3d30de15 /* (25, 9, 4) */,
  32'h3d81d711 /* (21, 9, 4) */,
  32'h3da3c1ed /* (17, 9, 4) */,
  32'h3d9d0afa /* (13, 9, 4) */,
  32'h3d51a9d2 /* (9, 9, 4) */,
  32'h3d1ee50b /* (5, 9, 4) */,
  32'h3d13f199 /* (1, 9, 4) */,
  32'h3d25f5ce /* (29, 5, 4) */,
  32'h3d1508af /* (25, 5, 4) */,
  32'h3d358341 /* (21, 5, 4) */,
  32'h3d4def9b /* (17, 5, 4) */,
  32'h3d4ea6a0 /* (13, 5, 4) */,
  32'h3d1ee50b /* (9, 5, 4) */,
  32'h3d189061 /* (5, 5, 4) */,
  32'h3d334ee4 /* (1, 5, 4) */,
  32'h3d6eb36b /* (29, 1, 4) */,
  32'h3d17ff6b /* (25, 1, 4) */,
  32'h3d1f5dc3 /* (21, 1, 4) */,
  32'h3d294c4b /* (17, 1, 4) */,
  32'h3d2e802a /* (13, 1, 4) */,
  32'h3d13f199 /* (9, 1, 4) */,
  32'h3d334ee4 /* (5, 1, 4) */,
  32'h3d9c757b /* (1, 1, 4) */,
  32'h3d9c797c /* (29, 29, 0) */,
  32'h3d1cfd70 /* (25, 29, 0) */,
  32'h3d198ce9 /* (21, 29, 0) */,
  32'h3d1eeabe /* (17, 29, 0) */,
  32'h3d258110 /* (13, 29, 0) */,
  32'h3d1237a7 /* (9, 29, 0) */,
  32'h3d490b0e /* (5, 29, 0) */,
  32'h3dff9e3f /* (1, 29, 0) */,
  32'h3d1cfd70 /* (29, 25, 0) */,
  32'h3d162f74 /* (25, 25, 0) */,
  32'h3d3dcd22 /* (21, 25, 0) */,
  32'h3d5b6048 /* (17, 25, 0) */,
  32'h3d5a6fdd /* (13, 25, 0) */,
  32'h3d23a039 /* (9, 25, 0) */,
  32'h3d154f7b /* (5, 25, 0) */,
  32'h3d25463b /* (1, 25, 0) */,
  32'h3d198ce9 /* (29, 21, 0) */,
  32'h3d3dcd22 /* (25, 21, 0) */,
  32'h3d922642 /* (21, 21, 0) */,
  32'h3dbe6d47 /* (17, 21, 0) */,
  32'h3db3fd83 /* (13, 21, 0) */,
  32'h3d66dac1 /* (9, 21, 0) */,
  32'h3d25e815 /* (5, 21, 0) */,
  32'h3d147e90 /* (1, 21, 0) */,
  32'h3d1eeabe /* (29, 17, 0) */,
  32'h3d5b6048 /* (25, 17, 0) */,
  32'h3dbe6d47 /* (21, 17, 0) */,
  32'h3e086183 /* (17, 17, 0) */,
  32'h3df6cc6d /* (13, 17, 0) */,
  32'h3d8df2c1 /* (9, 17, 0) */,
  32'h3d347f0a /* (5, 17, 0) */,
  32'h3d155505 /* (1, 17, 0) */,
  32'h3d258110 /* (29, 13, 0) */,
  32'h3d5a6fdd /* (25, 13, 0) */,
  32'h3db3fd83 /* (21, 13, 0) */,
  32'h3df6cc6d /* (17, 13, 0) */,
  32'h3de3e928 /* (13, 13, 0) */,
  32'h3d89a49e /* (9, 13, 0) */,
  32'h3d384488 /* (5, 13, 0) */,
  32'h3d1d4601 /* (1, 13, 0) */,
  32'h3d1237a7 /* (29, 9, 0) */,
  32'h3d23a039 /* (25, 9, 0) */,
  32'h3d66dac1 /* (21, 9, 0) */,
  32'h3d8df2c1 /* (17, 9, 0) */,
  32'h3d89a49e /* (13, 9, 0) */,
  32'h3d3dc47d /* (9, 9, 0) */,
  32'h3d16a564 /* (5, 9, 0) */,
  32'h3d11a5c6 /* (1, 9, 0) */,
  32'h3d490b0e /* (29, 5, 0) */,
  32'h3d154f7b /* (25, 5, 0) */,
  32'h3d25e815 /* (21, 5, 0) */,
  32'h3d347f0a /* (17, 5, 0) */,
  32'h3d384488 /* (13, 5, 0) */,
  32'h3d16a564 /* (9, 5, 0) */,
  32'h3d25e3da /* (5, 5, 0) */,
  32'h3d6e9998 /* (1, 5, 0) */,
  32'h3dff9e3f /* (29, 1, 0) */,
  32'h3d25463b /* (25, 1, 0) */,
  32'h3d147e90 /* (21, 1, 0) */,
  32'h3d155505 /* (17, 1, 0) */,
  32'h3d1d4601 /* (13, 1, 0) */,
  32'h3d11a5c6 /* (9, 1, 0) */,
  32'h3d6e9998 /* (5, 1, 0) */,
  32'h3f10fe39 /* (1, 1, 0) */,
  32'h3d358b49 /* (28, 29, 28) */,
  32'h3d13fed6 /* (24, 29, 28) */,
  32'h3d30047a /* (20, 29, 28) */,
  32'h3d232f37 /* (16, 29, 28) */,
  32'h3d30047a /* (12, 29, 28) */,
  32'h3d13fed6 /* (8, 29, 28) */,
  32'h3d358b49 /* (4, 29, 28) */,
  32'h3d7541a2 /* (0, 29, 28) */,
  32'h3d148979 /* (28, 25, 28) */,
  32'h3d250b86 /* (24, 25, 28) */,
  32'h3d66108f /* (20, 25, 28) */,
  32'h3d66e7bc /* (16, 25, 28) */,
  32'h3d66108f /* (12, 25, 28) */,
  32'h3d250b86 /* (8, 25, 28) */,
  32'h3d148979 /* (4, 25, 28) */,
  32'h3d1879c9 /* (0, 25, 28) */,
  32'h3d2c64eb /* (28, 21, 28) */,
  32'h3d683712 /* (24, 21, 28) */,
  32'h3dbb90ec /* (20, 21, 28) */,
  32'h3dcebbc1 /* (16, 21, 28) */,
  32'h3dbb90ec /* (12, 21, 28) */,
  32'h3d683712 /* (8, 21, 28) */,
  32'h3d2c64eb /* (4, 21, 28) */,
  32'h3d1e982c /* (0, 21, 28) */,
  32'h3d3f317e /* (28, 17, 28) */,
  32'h3d8e8b3a /* (24, 17, 28) */,
  32'h3dff07bf /* (20, 17, 28) */,
  32'h3e18449a /* (16, 17, 28) */,
  32'h3dff07bf /* (12, 17, 28) */,
  32'h3d8e8b3a /* (8, 17, 28) */,
  32'h3d3f317e /* (4, 17, 28) */,
  32'h3d27f384 /* (0, 17, 28) */,
  32'h3d41aa67 /* (28, 13, 28) */,
  32'h3d8a5278 /* (24, 13, 28) */,
  32'h3dec6d9f /* (20, 13, 28) */,
  32'h3e07f264 /* (16, 13, 28) */,
  32'h3dec6d9f /* (12, 13, 28) */,
  32'h3d8a5278 /* (8, 13, 28) */,
  32'h3d41aa67 /* (4, 13, 28) */,
  32'h3d2d543a /* (0, 13, 28) */,
  32'h3d19e157 /* (28, 9, 28) */,
  32'h3d3f1eea /* (24, 9, 28) */,
  32'h3d902ce0 /* (20, 9, 28) */,
  32'h3d97bb42 /* (16, 9, 28) */,
  32'h3d902ce0 /* (12, 9, 28) */,
  32'h3d3f1eea /* (8, 9, 28) */,
  32'h3d19e157 /* (4, 9, 28) */,
  32'h3d13aacb /* (0, 9, 28) */,
  32'h3d1e7527 /* (28, 5, 28) */,
  32'h3d183845 /* (24, 5, 28) */,
  32'h3d431db1 /* (20, 5, 28) */,
  32'h3d3b5943 /* (16, 5, 28) */,
  32'h3d431db1 /* (12, 5, 28) */,
  32'h3d183845 /* (8, 5, 28) */,
  32'h3d1e7527 /* (4, 5, 28) */,
  32'h3d3577a5 /* (0, 5, 28) */,
  32'h3d4cb45d /* (28, 1, 28) */,
  32'h3d139499 /* (24, 1, 28) */,
  32'h3d27af27 /* (20, 1, 28) */,
  32'h3d18708b /* (16, 1, 28) */,
  32'h3d27af27 /* (12, 1, 28) */,
  32'h3d139499 /* (8, 1, 28) */,
  32'h3d4cb45d /* (4, 1, 28) */,
  32'h3da3aa58 /* (0, 1, 28) */,
  32'h3d13fed6 /* (28, 29, 24) */,
  32'h3d2a2238 /* (24, 29, 24) */,
  32'h3d729483 /* (20, 29, 24) */,
  32'h3d76a38f /* (16, 29, 24) */,
  32'h3d729483 /* (12, 29, 24) */,
  32'h3d2a2238 /* (8, 29, 24) */,
  32'h3d13fed6 /* (4, 29, 24) */,
  32'h3d14a194 /* (0, 29, 24) */,
  32'h3d250b86 /* (28, 25, 24) */,
  32'h3d54dbd1 /* (24, 25, 24) */,
  32'h3da58a7f /* (20, 25, 24) */,
  32'h3db1ba44 /* (16, 25, 24) */,
  32'h3da58a7f /* (12, 25, 24) */,
  32'h3d54dbd1 /* (8, 25, 24) */,
  32'h3d250b86 /* (4, 25, 24) */,
  32'h3d1b34b2 /* (0, 25, 24) */,
  32'h3d683712 /* (28, 21, 24) */,
  32'h3da5dafd /* (24, 21, 24) */,
  32'h3e0dbead /* (20, 21, 24) */,
  32'h3e2301df /* (16, 21, 24) */,
  32'h3e0dbead /* (12, 21, 24) */,
  32'h3da5dafd /* (8, 21, 24) */,
  32'h3d683712 /* (4, 21, 24) */,
  32'h3d4fd499 /* (0, 21, 24) */,
  32'h3d8e8b3a /* (28, 17, 24) */,
  32'h3dd9f1d0 /* (24, 17, 24) */,
  32'h3e48a298 /* (20, 17, 24) */,
  32'h3e75b861 /* (16, 17, 24) */,
  32'h3e48a298 /* (12, 17, 24) */,
  32'h3dd9f1d0 /* (8, 17, 24) */,
  32'h3d8e8b3a /* (4, 17, 24) */,
  32'h3d77d78b /* (0, 17, 24) */,
  32'h3d8a5278 /* (28, 13, 24) */,
  32'h3dcd36cb /* (24, 13, 24) */,
  32'h3e368e5b /* (20, 13, 24) */,
  32'h3e58f4b1 /* (16, 13, 24) */,
  32'h3e368e5b /* (12, 13, 24) */,
  32'h3dcd36cb /* (8, 13, 24) */,
  32'h3d8a5278 /* (4, 13, 24) */,
  32'h3d7388b1 /* (0, 13, 24) */,
  32'h3d3f1eea /* (28, 9, 24) */,
  32'h3d824402 /* (24, 9, 24) */,
  32'h3dd4c19e /* (20, 9, 24) */,
  32'h3dec5cc9 /* (16, 9, 24) */,
  32'h3dd4c19e /* (12, 9, 24) */,
  32'h3d824402 /* (8, 9, 24) */,
  32'h3d3f1eea /* (4, 9, 24) */,
  32'h3d2eceba /* (0, 9, 24) */,
  32'h3d183845 /* (28, 5, 24) */,
  32'h3d38dbff /* (24, 5, 24) */,
  32'h3d89129f /* (20, 5, 24) */,
  32'h3d8eb3bf /* (16, 5, 24) */,
  32'h3d89129f /* (12, 5, 24) */,
  32'h3d38dbff /* (8, 5, 24) */,
  32'h3d183845 /* (4, 5, 24) */,
  32'h3d13eed3 /* (0, 5, 24) */,
  32'h3d139499 /* (28, 1, 24) */,
  32'h3d23fb6f /* (24, 1, 24) */,
  32'h3d649547 /* (20, 1, 24) */,
  32'h3d656b11 /* (16, 1, 24) */,
  32'h3d649547 /* (12, 1, 24) */,
  32'h3d23fb6f /* (8, 1, 24) */,
  32'h3d139499 /* (4, 1, 24) */,
  32'h3d177e6a /* (0, 1, 24) */,
  32'h3d30047a /* (28, 29, 20) */,
  32'h3d729483 /* (24, 29, 20) */,
  32'h3dc823b1 /* (20, 29, 20) */,
  32'h3de007f6 /* (16, 29, 20) */,
  32'h3dc823b1 /* (12, 29, 20) */,
  32'h3d729483 /* (8, 29, 20) */,
  32'h3d30047a /* (4, 29, 20) */,
  32'h3d202826 /* (0, 29, 20) */,
  32'h3d66108f /* (28, 25, 20) */,
  32'h3da58a7f /* (24, 25, 20) */,
  32'h3e0e8e1e /* (20, 25, 20) */,
  32'h3e24eefd /* (16, 25, 20) */,
  32'h3e0e8e1e /* (12, 25, 20) */,
  32'h3da58a7f /* (8, 25, 20) */,
  32'h3d66108f /* (4, 25, 20) */,
  32'h3d4d39f8 /* (0, 25, 20) */,
  32'h3dbb90ec /* (28, 21, 20) */,
  32'h3e0dbead /* (24, 21, 20) */,
  32'h3e80c082 /* (20, 21, 20) */,
  32'h3e9bce24 /* (16, 21, 20) */,
  32'h3e80c082 /* (12, 21, 20) */,
  32'h3e0dbead /* (8, 21, 20) */,
  32'h3dbb90ec /* (4, 21, 20) */,
  32'h3da3d600 /* (0, 21, 20) */,
  32'h3dff07bf /* (28, 17, 20) */,
  32'h3e48a298 /* (24, 17, 20) */,
  32'h3ebf3a63 /* (20, 17, 20) */,
  32'h3ef1f40b /* (16, 17, 20) */,
  32'h3ebf3a63 /* (12, 17, 20) */,
  32'h3e48a298 /* (8, 17, 20) */,
  32'h3dff07bf /* (4, 17, 20) */,
  32'h3ddb309a /* (0, 17, 20) */,
  32'h3dec6d9f /* (28, 13, 20) */,
  32'h3e368e5b /* (24, 13, 20) */,
  32'h3eaa0eb2 /* (20, 13, 20) */,
  32'h3ed28b29 /* (16, 13, 20) */,
  32'h3eaa0eb2 /* (12, 13, 20) */,
  32'h3e368e5b /* (8, 13, 20) */,
  32'h3dec6d9f /* (4, 13, 20) */,
  32'h3dccb681 /* (0, 13, 20) */,
  32'h3d902ce0 /* (28, 9, 20) */,
  32'h3dd4c19e /* (24, 9, 20) */,
  32'h3e3c290c /* (20, 9, 20) */,
  32'h3e5e82df /* (16, 9, 20) */,
  32'h3e3c290c /* (12, 9, 20) */,
  32'h3dd4c19e /* (8, 9, 20) */,
  32'h3d902ce0 /* (4, 9, 20) */,
  32'h3d7e6b4b /* (0, 9, 20) */,
  32'h3d431db1 /* (28, 5, 20) */,
  32'h3d89129f /* (24, 5, 20) */,
  32'h3de671da /* (20, 5, 20) */,
  32'h3e02cee2 /* (16, 5, 20) */,
  32'h3de671da /* (12, 5, 20) */,
  32'h3d89129f /* (8, 5, 20) */,
  32'h3d431db1 /* (4, 5, 20) */,
  32'h3d2ff16f /* (0, 5, 20) */,
  32'h3d27af27 /* (28, 1, 20) */,
  32'h3d649547 /* (24, 1, 20) */,
  32'h3dbaaaa9 /* (20, 1, 20) */,
  32'h3dcf60c6 /* (16, 1, 20) */,
  32'h3dbaaaa9 /* (12, 1, 20) */,
  32'h3d649547 /* (8, 1, 20) */,
  32'h3d27af27 /* (4, 1, 20) */,
  32'h3d195f14 /* (0, 1, 20) */,
  32'h3d232f37 /* (28, 29, 16) */,
  32'h3d76a38f /* (24, 29, 16) */,
  32'h3de007f6 /* (20, 29, 16) */,
  32'h3e078d5a /* (16, 29, 16) */,
  32'h3de007f6 /* (12, 29, 16) */,
  32'h3d76a38f /* (8, 29, 16) */,
  32'h3d232f37 /* (4, 29, 16) */,
  32'h3d0e89f8 /* (0, 29, 16) */,
  32'h3d66e7bc /* (28, 25, 16) */,
  32'h3db1ba44 /* (24, 25, 16) */,
  32'h3e24eefd /* (20, 25, 16) */,
  32'h3e4b7c7a /* (16, 25, 16) */,
  32'h3e24eefd /* (12, 25, 16) */,
  32'h3db1ba44 /* (8, 25, 16) */,
  32'h3d66e7bc /* (4, 25, 16) */,
  32'h3d482f92 /* (0, 25, 16) */,
  32'h3dcebbc1 /* (28, 21, 16) */,
  32'h3e2301df /* (24, 21, 16) */,
  32'h3e9bce24 /* (20, 21, 16) */,
  32'h3ec5ad99 /* (16, 21, 16) */,
  32'h3e9bce24 /* (12, 21, 16) */,
  32'h3e2301df /* (8, 21, 16) */,
  32'h3dcebbc1 /* (4, 21, 16) */,
  32'h3db1860e /* (0, 21, 16) */,
  32'h3e18449a /* (28, 17, 16) */,
  32'h3e75b861 /* (24, 17, 16) */,
  32'h3ef1f40b /* (20, 17, 16) */,
  32'h3f1e253a /* (16, 17, 16) */,
  32'h3ef1f40b /* (12, 17, 16) */,
  32'h3e75b861 /* (8, 17, 16) */,
  32'h3e18449a /* (4, 17, 16) */,
  32'h3e019a4f /* (0, 17, 16) */,
  32'h3e07f264 /* (28, 13, 16) */,
  32'h3e58f4b1 /* (24, 13, 16) */,
  32'h3ed28b29 /* (20, 13, 16) */,
  32'h3f079668 /* (16, 13, 16) */,
  32'h3ed28b29 /* (12, 13, 16) */,
  32'h3e58f4b1 /* (8, 13, 16) */,
  32'h3e07f264 /* (4, 13, 16) */,
  32'h3de8675d /* (0, 13, 16) */,
  32'h3d97bb42 /* (28, 9, 16) */,
  32'h3dec5cc9 /* (24, 9, 16) */,
  32'h3e5e82df /* (20, 9, 16) */,
  32'h3e8b1bdf /* (16, 9, 16) */,
  32'h3e5e82df /* (12, 9, 16) */,
  32'h3dec5cc9 /* (8, 9, 16) */,
  32'h3d97bb42 /* (4, 9, 16) */,
  32'h3d82ec35 /* (0, 9, 16) */,
  32'h3d3b5943 /* (28, 5, 16) */,
  32'h3d8eb3bf /* (24, 5, 16) */,
  32'h3e02cee2 /* (20, 5, 16) */,
  32'h3e1f95bf /* (16, 5, 16) */,
  32'h3e02cee2 /* (12, 5, 16) */,
  32'h3d8eb3bf /* (8, 5, 16) */,
  32'h3d3b5943 /* (4, 5, 16) */,
  32'h3d231d8f /* (0, 5, 16) */,
  32'h3d18708b /* (28, 1, 16) */,
  32'h3d656b11 /* (24, 1, 16) */,
  32'h3dcf60c6 /* (20, 1, 16) */,
  32'h3df9e164 /* (16, 1, 16) */,
  32'h3dcf60c6 /* (12, 1, 16) */,
  32'h3d656b11 /* (8, 1, 16) */,
  32'h3d18708b /* (4, 1, 16) */,
  32'h3d0563b9 /* (0, 1, 16) */,
  32'h3d30047a /* (28, 29, 12) */,
  32'h3d729483 /* (24, 29, 12) */,
  32'h3dc823b1 /* (20, 29, 12) */,
  32'h3de007f6 /* (16, 29, 12) */,
  32'h3dc823b1 /* (12, 29, 12) */,
  32'h3d729483 /* (8, 29, 12) */,
  32'h3d30047a /* (4, 29, 12) */,
  32'h3d202826 /* (0, 29, 12) */,
  32'h3d66108f /* (28, 25, 12) */,
  32'h3da58a7f /* (24, 25, 12) */,
  32'h3e0e8e1e /* (20, 25, 12) */,
  32'h3e24eefd /* (16, 25, 12) */,
  32'h3e0e8e1e /* (12, 25, 12) */,
  32'h3da58a7f /* (8, 25, 12) */,
  32'h3d66108f /* (4, 25, 12) */,
  32'h3d4d39f8 /* (0, 25, 12) */,
  32'h3dbb90ec /* (28, 21, 12) */,
  32'h3e0dbead /* (24, 21, 12) */,
  32'h3e80c082 /* (20, 21, 12) */,
  32'h3e9bce24 /* (16, 21, 12) */,
  32'h3e80c082 /* (12, 21, 12) */,
  32'h3e0dbead /* (8, 21, 12) */,
  32'h3dbb90ec /* (4, 21, 12) */,
  32'h3da3d600 /* (0, 21, 12) */,
  32'h3dff07bf /* (28, 17, 12) */,
  32'h3e48a298 /* (24, 17, 12) */,
  32'h3ebf3a63 /* (20, 17, 12) */,
  32'h3ef1f40b /* (16, 17, 12) */,
  32'h3ebf3a63 /* (12, 17, 12) */,
  32'h3e48a298 /* (8, 17, 12) */,
  32'h3dff07bf /* (4, 17, 12) */,
  32'h3ddb309a /* (0, 17, 12) */,
  32'h3dec6d9f /* (28, 13, 12) */,
  32'h3e368e5b /* (24, 13, 12) */,
  32'h3eaa0eb2 /* (20, 13, 12) */,
  32'h3ed28b29 /* (16, 13, 12) */,
  32'h3eaa0eb2 /* (12, 13, 12) */,
  32'h3e368e5b /* (8, 13, 12) */,
  32'h3dec6d9f /* (4, 13, 12) */,
  32'h3dccb681 /* (0, 13, 12) */,
  32'h3d902ce0 /* (28, 9, 12) */,
  32'h3dd4c19e /* (24, 9, 12) */,
  32'h3e3c290c /* (20, 9, 12) */,
  32'h3e5e82df /* (16, 9, 12) */,
  32'h3e3c290c /* (12, 9, 12) */,
  32'h3dd4c19e /* (8, 9, 12) */,
  32'h3d902ce0 /* (4, 9, 12) */,
  32'h3d7e6b4b /* (0, 9, 12) */,
  32'h3d431db1 /* (28, 5, 12) */,
  32'h3d89129f /* (24, 5, 12) */,
  32'h3de671da /* (20, 5, 12) */,
  32'h3e02cee2 /* (16, 5, 12) */,
  32'h3de671da /* (12, 5, 12) */,
  32'h3d89129f /* (8, 5, 12) */,
  32'h3d431db1 /* (4, 5, 12) */,
  32'h3d2ff16f /* (0, 5, 12) */,
  32'h3d27af27 /* (28, 1, 12) */,
  32'h3d649547 /* (24, 1, 12) */,
  32'h3dbaaaa9 /* (20, 1, 12) */,
  32'h3dcf60c6 /* (16, 1, 12) */,
  32'h3dbaaaa9 /* (12, 1, 12) */,
  32'h3d649547 /* (8, 1, 12) */,
  32'h3d27af27 /* (4, 1, 12) */,
  32'h3d195f14 /* (0, 1, 12) */,
  32'h3d13fed6 /* (28, 29, 8) */,
  32'h3d2a2238 /* (24, 29, 8) */,
  32'h3d729483 /* (20, 29, 8) */,
  32'h3d76a38f /* (16, 29, 8) */,
  32'h3d729483 /* (12, 29, 8) */,
  32'h3d2a2238 /* (8, 29, 8) */,
  32'h3d13fed6 /* (4, 29, 8) */,
  32'h3d14a194 /* (0, 29, 8) */,
  32'h3d250b86 /* (28, 25, 8) */,
  32'h3d54dbd1 /* (24, 25, 8) */,
  32'h3da58a7f /* (20, 25, 8) */,
  32'h3db1ba44 /* (16, 25, 8) */,
  32'h3da58a7f /* (12, 25, 8) */,
  32'h3d54dbd1 /* (8, 25, 8) */,
  32'h3d250b86 /* (4, 25, 8) */,
  32'h3d1b34b2 /* (0, 25, 8) */,
  32'h3d683712 /* (28, 21, 8) */,
  32'h3da5dafd /* (24, 21, 8) */,
  32'h3e0dbead /* (20, 21, 8) */,
  32'h3e2301df /* (16, 21, 8) */,
  32'h3e0dbead /* (12, 21, 8) */,
  32'h3da5dafd /* (8, 21, 8) */,
  32'h3d683712 /* (4, 21, 8) */,
  32'h3d4fd499 /* (0, 21, 8) */,
  32'h3d8e8b3a /* (28, 17, 8) */,
  32'h3dd9f1d0 /* (24, 17, 8) */,
  32'h3e48a298 /* (20, 17, 8) */,
  32'h3e75b861 /* (16, 17, 8) */,
  32'h3e48a298 /* (12, 17, 8) */,
  32'h3dd9f1d0 /* (8, 17, 8) */,
  32'h3d8e8b3a /* (4, 17, 8) */,
  32'h3d77d78b /* (0, 17, 8) */,
  32'h3d8a5278 /* (28, 13, 8) */,
  32'h3dcd36cb /* (24, 13, 8) */,
  32'h3e368e5b /* (20, 13, 8) */,
  32'h3e58f4b1 /* (16, 13, 8) */,
  32'h3e368e5b /* (12, 13, 8) */,
  32'h3dcd36cb /* (8, 13, 8) */,
  32'h3d8a5278 /* (4, 13, 8) */,
  32'h3d7388b1 /* (0, 13, 8) */,
  32'h3d3f1eea /* (28, 9, 8) */,
  32'h3d824402 /* (24, 9, 8) */,
  32'h3dd4c19e /* (20, 9, 8) */,
  32'h3dec5cc9 /* (16, 9, 8) */,
  32'h3dd4c19e /* (12, 9, 8) */,
  32'h3d824402 /* (8, 9, 8) */,
  32'h3d3f1eea /* (4, 9, 8) */,
  32'h3d2eceba /* (0, 9, 8) */,
  32'h3d183845 /* (28, 5, 8) */,
  32'h3d38dbff /* (24, 5, 8) */,
  32'h3d89129f /* (20, 5, 8) */,
  32'h3d8eb3bf /* (16, 5, 8) */,
  32'h3d89129f /* (12, 5, 8) */,
  32'h3d38dbff /* (8, 5, 8) */,
  32'h3d183845 /* (4, 5, 8) */,
  32'h3d13eed3 /* (0, 5, 8) */,
  32'h3d139499 /* (28, 1, 8) */,
  32'h3d23fb6f /* (24, 1, 8) */,
  32'h3d649547 /* (20, 1, 8) */,
  32'h3d656b11 /* (16, 1, 8) */,
  32'h3d649547 /* (12, 1, 8) */,
  32'h3d23fb6f /* (8, 1, 8) */,
  32'h3d139499 /* (4, 1, 8) */,
  32'h3d177e6a /* (0, 1, 8) */,
  32'h3d358b49 /* (28, 29, 4) */,
  32'h3d13fed6 /* (24, 29, 4) */,
  32'h3d30047a /* (20, 29, 4) */,
  32'h3d232f37 /* (16, 29, 4) */,
  32'h3d30047a /* (12, 29, 4) */,
  32'h3d13fed6 /* (8, 29, 4) */,
  32'h3d358b49 /* (4, 29, 4) */,
  32'h3d7541a2 /* (0, 29, 4) */,
  32'h3d148979 /* (28, 25, 4) */,
  32'h3d250b86 /* (24, 25, 4) */,
  32'h3d66108f /* (20, 25, 4) */,
  32'h3d66e7bc /* (16, 25, 4) */,
  32'h3d66108f /* (12, 25, 4) */,
  32'h3d250b86 /* (8, 25, 4) */,
  32'h3d148979 /* (4, 25, 4) */,
  32'h3d1879c9 /* (0, 25, 4) */,
  32'h3d2c64eb /* (28, 21, 4) */,
  32'h3d683712 /* (24, 21, 4) */,
  32'h3dbb90ec /* (20, 21, 4) */,
  32'h3dcebbc1 /* (16, 21, 4) */,
  32'h3dbb90ec /* (12, 21, 4) */,
  32'h3d683712 /* (8, 21, 4) */,
  32'h3d2c64eb /* (4, 21, 4) */,
  32'h3d1e982c /* (0, 21, 4) */,
  32'h3d3f317e /* (28, 17, 4) */,
  32'h3d8e8b3a /* (24, 17, 4) */,
  32'h3dff07bf /* (20, 17, 4) */,
  32'h3e18449a /* (16, 17, 4) */,
  32'h3dff07bf /* (12, 17, 4) */,
  32'h3d8e8b3a /* (8, 17, 4) */,
  32'h3d3f317e /* (4, 17, 4) */,
  32'h3d27f384 /* (0, 17, 4) */,
  32'h3d41aa67 /* (28, 13, 4) */,
  32'h3d8a5278 /* (24, 13, 4) */,
  32'h3dec6d9f /* (20, 13, 4) */,
  32'h3e07f264 /* (16, 13, 4) */,
  32'h3dec6d9f /* (12, 13, 4) */,
  32'h3d8a5278 /* (8, 13, 4) */,
  32'h3d41aa67 /* (4, 13, 4) */,
  32'h3d2d543a /* (0, 13, 4) */,
  32'h3d19e157 /* (28, 9, 4) */,
  32'h3d3f1eea /* (24, 9, 4) */,
  32'h3d902ce0 /* (20, 9, 4) */,
  32'h3d97bb42 /* (16, 9, 4) */,
  32'h3d902ce0 /* (12, 9, 4) */,
  32'h3d3f1eea /* (8, 9, 4) */,
  32'h3d19e157 /* (4, 9, 4) */,
  32'h3d13aacb /* (0, 9, 4) */,
  32'h3d1e7527 /* (28, 5, 4) */,
  32'h3d183845 /* (24, 5, 4) */,
  32'h3d431db1 /* (20, 5, 4) */,
  32'h3d3b5943 /* (16, 5, 4) */,
  32'h3d431db1 /* (12, 5, 4) */,
  32'h3d183845 /* (8, 5, 4) */,
  32'h3d1e7527 /* (4, 5, 4) */,
  32'h3d3577a5 /* (0, 5, 4) */,
  32'h3d4cb45d /* (28, 1, 4) */,
  32'h3d139499 /* (24, 1, 4) */,
  32'h3d27af27 /* (20, 1, 4) */,
  32'h3d18708b /* (16, 1, 4) */,
  32'h3d27af27 /* (12, 1, 4) */,
  32'h3d139499 /* (8, 1, 4) */,
  32'h3d4cb45d /* (4, 1, 4) */,
  32'h3da3aa58 /* (0, 1, 4) */,
  32'h3d7541a2 /* (28, 29, 0) */,
  32'h3d14a194 /* (24, 29, 0) */,
  32'h3d202826 /* (20, 29, 0) */,
  32'h3d0e89f8 /* (16, 29, 0) */,
  32'h3d202826 /* (12, 29, 0) */,
  32'h3d14a194 /* (8, 29, 0) */,
  32'h3d7541a2 /* (4, 29, 0) */,
  32'h3e0c4c59 /* (0, 29, 0) */,
  32'h3d1879c9 /* (28, 25, 0) */,
  32'h3d1b34b2 /* (24, 25, 0) */,
  32'h3d4d39f8 /* (20, 25, 0) */,
  32'h3d482f92 /* (16, 25, 0) */,
  32'h3d4d39f8 /* (12, 25, 0) */,
  32'h3d1b34b2 /* (8, 25, 0) */,
  32'h3d1879c9 /* (4, 25, 0) */,
  32'h3d269d45 /* (0, 25, 0) */,
  32'h3d1e982c /* (28, 21, 0) */,
  32'h3d4fd499 /* (24, 21, 0) */,
  32'h3da3d600 /* (20, 21, 0) */,
  32'h3db1860e /* (16, 21, 0) */,
  32'h3da3d600 /* (12, 21, 0) */,
  32'h3d4fd499 /* (8, 21, 0) */,
  32'h3d1e982c /* (4, 21, 0) */,
  32'h3d13eab3 /* (0, 21, 0) */,
  32'h3d27f384 /* (28, 17, 0) */,
  32'h3d77d78b /* (24, 17, 0) */,
  32'h3ddb309a /* (20, 17, 0) */,
  32'h3e019a4f /* (16, 17, 0) */,
  32'h3ddb309a /* (12, 17, 0) */,
  32'h3d77d78b /* (8, 17, 0) */,
  32'h3d27f384 /* (4, 17, 0) */,
  32'h3d14300c /* (0, 17, 0) */,
  32'h3d2d543a /* (28, 13, 0) */,
  32'h3d7388b1 /* (24, 13, 0) */,
  32'h3dccb681 /* (20, 13, 0) */,
  32'h3de8675d /* (16, 13, 0) */,
  32'h3dccb681 /* (12, 13, 0) */,
  32'h3d7388b1 /* (8, 13, 0) */,
  32'h3d2d543a /* (4, 13, 0) */,
  32'h3d1c4c09 /* (0, 13, 0) */,
  32'h3d13aacb /* (28, 9, 0) */,
  32'h3d2eceba /* (24, 9, 0) */,
  32'h3d7e6b4b /* (20, 9, 0) */,
  32'h3d82ec35 /* (16, 9, 0) */,
  32'h3d7e6b4b /* (12, 9, 0) */,
  32'h3d2eceba /* (8, 9, 0) */,
  32'h3d13aacb /* (4, 9, 0) */,
  32'h3d11ab15 /* (0, 9, 0) */,
  32'h3d3577a5 /* (28, 5, 0) */,
  32'h3d13eed3 /* (24, 5, 0) */,
  32'h3d2ff16f /* (20, 5, 0) */,
  32'h3d231d8f /* (16, 5, 0) */,
  32'h3d2ff16f /* (12, 5, 0) */,
  32'h3d13eed3 /* (8, 5, 0) */,
  32'h3d3577a5 /* (4, 5, 0) */,
  32'h3d75271a /* (0, 5, 0) */,
  32'h3da3aa58 /* (28, 1, 0) */,
  32'h3d177e6a /* (24, 1, 0) */,
  32'h3d195f14 /* (20, 1, 0) */,
  32'h3d0563b9 /* (16, 1, 0) */,
  32'h3d195f14 /* (12, 1, 0) */,
  32'h3d177e6a /* (8, 1, 0) */,
  32'h3da3aa58 /* (4, 1, 0) */,
  32'h3f8f3ec8 /* (0, 1, 0) */,
  32'h3d4cb45d /* (31, 28, 28) */,
  32'h3d1e7527 /* (27, 28, 28) */,
  32'h3d19e157 /* (23, 28, 28) */,
  32'h3d41aa67 /* (19, 28, 28) */,
  32'h3d3f317e /* (15, 28, 28) */,
  32'h3d2c64eb /* (11, 28, 28) */,
  32'h3d148979 /* (7, 28, 28) */,
  32'h3d358b49 /* (3, 28, 28) */,
  32'h3d139499 /* (31, 24, 28) */,
  32'h3d183845 /* (27, 24, 28) */,
  32'h3d3f1eea /* (23, 24, 28) */,
  32'h3d8a5278 /* (19, 24, 28) */,
  32'h3d8e8b3a /* (15, 24, 28) */,
  32'h3d683712 /* (11, 24, 28) */,
  32'h3d250b86 /* (7, 24, 28) */,
  32'h3d13fed6 /* (3, 24, 28) */,
  32'h3d27af27 /* (31, 20, 28) */,
  32'h3d431db1 /* (27, 20, 28) */,
  32'h3d902ce0 /* (23, 20, 28) */,
  32'h3dec6d9f /* (19, 20, 28) */,
  32'h3dff07bf /* (15, 20, 28) */,
  32'h3dbb90ec /* (11, 20, 28) */,
  32'h3d66108f /* (7, 20, 28) */,
  32'h3d30047a /* (3, 20, 28) */,
  32'h3d18708b /* (31, 16, 28) */,
  32'h3d3b5943 /* (27, 16, 28) */,
  32'h3d97bb42 /* (23, 16, 28) */,
  32'h3e07f264 /* (19, 16, 28) */,
  32'h3e18449a /* (15, 16, 28) */,
  32'h3dcebbc1 /* (11, 16, 28) */,
  32'h3d66e7bc /* (7, 16, 28) */,
  32'h3d232f37 /* (3, 16, 28) */,
  32'h3d27af27 /* (31, 12, 28) */,
  32'h3d431db1 /* (27, 12, 28) */,
  32'h3d902ce0 /* (23, 12, 28) */,
  32'h3dec6d9f /* (19, 12, 28) */,
  32'h3dff07bf /* (15, 12, 28) */,
  32'h3dbb90ec /* (11, 12, 28) */,
  32'h3d66108f /* (7, 12, 28) */,
  32'h3d30047a /* (3, 12, 28) */,
  32'h3d139499 /* (31, 8, 28) */,
  32'h3d183845 /* (27, 8, 28) */,
  32'h3d3f1eea /* (23, 8, 28) */,
  32'h3d8a5278 /* (19, 8, 28) */,
  32'h3d8e8b3a /* (15, 8, 28) */,
  32'h3d683712 /* (11, 8, 28) */,
  32'h3d250b86 /* (7, 8, 28) */,
  32'h3d13fed6 /* (3, 8, 28) */,
  32'h3d4cb45d /* (31, 4, 28) */,
  32'h3d1e7527 /* (27, 4, 28) */,
  32'h3d19e157 /* (23, 4, 28) */,
  32'h3d41aa67 /* (19, 4, 28) */,
  32'h3d3f317e /* (15, 4, 28) */,
  32'h3d2c64eb /* (11, 4, 28) */,
  32'h3d148979 /* (7, 4, 28) */,
  32'h3d358b49 /* (3, 4, 28) */,
  32'h3da3aa58 /* (31, 0, 28) */,
  32'h3d3577a5 /* (27, 0, 28) */,
  32'h3d13aacb /* (23, 0, 28) */,
  32'h3d2d543a /* (19, 0, 28) */,
  32'h3d27f384 /* (15, 0, 28) */,
  32'h3d1e982c /* (11, 0, 28) */,
  32'h3d1879c9 /* (7, 0, 28) */,
  32'h3d7541a2 /* (3, 0, 28) */,
  32'h3d139499 /* (31, 28, 24) */,
  32'h3d183845 /* (27, 28, 24) */,
  32'h3d3f1eea /* (23, 28, 24) */,
  32'h3d8a5278 /* (19, 28, 24) */,
  32'h3d8e8b3a /* (15, 28, 24) */,
  32'h3d683712 /* (11, 28, 24) */,
  32'h3d250b86 /* (7, 28, 24) */,
  32'h3d13fed6 /* (3, 28, 24) */,
  32'h3d23fb6f /* (31, 24, 24) */,
  32'h3d38dbff /* (27, 24, 24) */,
  32'h3d824402 /* (23, 24, 24) */,
  32'h3dcd36cb /* (19, 24, 24) */,
  32'h3dd9f1d0 /* (15, 24, 24) */,
  32'h3da5dafd /* (11, 24, 24) */,
  32'h3d54dbd1 /* (7, 24, 24) */,
  32'h3d2a2238 /* (3, 24, 24) */,
  32'h3d649547 /* (31, 20, 24) */,
  32'h3d89129f /* (27, 20, 24) */,
  32'h3dd4c19e /* (23, 20, 24) */,
  32'h3e368e5b /* (19, 20, 24) */,
  32'h3e48a298 /* (15, 20, 24) */,
  32'h3e0dbead /* (11, 20, 24) */,
  32'h3da58a7f /* (7, 20, 24) */,
  32'h3d729483 /* (3, 20, 24) */,
  32'h3d656b11 /* (31, 16, 24) */,
  32'h3d8eb3bf /* (27, 16, 24) */,
  32'h3dec5cc9 /* (23, 16, 24) */,
  32'h3e58f4b1 /* (19, 16, 24) */,
  32'h3e75b861 /* (15, 16, 24) */,
  32'h3e2301df /* (11, 16, 24) */,
  32'h3db1ba44 /* (7, 16, 24) */,
  32'h3d76a38f /* (3, 16, 24) */,
  32'h3d649547 /* (31, 12, 24) */,
  32'h3d89129f /* (27, 12, 24) */,
  32'h3dd4c19e /* (23, 12, 24) */,
  32'h3e368e5b /* (19, 12, 24) */,
  32'h3e48a298 /* (15, 12, 24) */,
  32'h3e0dbead /* (11, 12, 24) */,
  32'h3da58a7f /* (7, 12, 24) */,
  32'h3d729483 /* (3, 12, 24) */,
  32'h3d23fb6f /* (31, 8, 24) */,
  32'h3d38dbff /* (27, 8, 24) */,
  32'h3d824402 /* (23, 8, 24) */,
  32'h3dcd36cb /* (19, 8, 24) */,
  32'h3dd9f1d0 /* (15, 8, 24) */,
  32'h3da5dafd /* (11, 8, 24) */,
  32'h3d54dbd1 /* (7, 8, 24) */,
  32'h3d2a2238 /* (3, 8, 24) */,
  32'h3d139499 /* (31, 4, 24) */,
  32'h3d183845 /* (27, 4, 24) */,
  32'h3d3f1eea /* (23, 4, 24) */,
  32'h3d8a5278 /* (19, 4, 24) */,
  32'h3d8e8b3a /* (15, 4, 24) */,
  32'h3d683712 /* (11, 4, 24) */,
  32'h3d250b86 /* (7, 4, 24) */,
  32'h3d13fed6 /* (3, 4, 24) */,
  32'h3d177e6a /* (31, 0, 24) */,
  32'h3d13eed3 /* (27, 0, 24) */,
  32'h3d2eceba /* (23, 0, 24) */,
  32'h3d7388b1 /* (19, 0, 24) */,
  32'h3d77d78b /* (15, 0, 24) */,
  32'h3d4fd499 /* (11, 0, 24) */,
  32'h3d1b34b2 /* (7, 0, 24) */,
  32'h3d14a194 /* (3, 0, 24) */,
  32'h3d27af27 /* (31, 28, 20) */,
  32'h3d431db1 /* (27, 28, 20) */,
  32'h3d902ce0 /* (23, 28, 20) */,
  32'h3dec6d9f /* (19, 28, 20) */,
  32'h3dff07bf /* (15, 28, 20) */,
  32'h3dbb90ec /* (11, 28, 20) */,
  32'h3d66108f /* (7, 28, 20) */,
  32'h3d30047a /* (3, 28, 20) */,
  32'h3d649547 /* (31, 24, 20) */,
  32'h3d89129f /* (27, 24, 20) */,
  32'h3dd4c19e /* (23, 24, 20) */,
  32'h3e368e5b /* (19, 24, 20) */,
  32'h3e48a298 /* (15, 24, 20) */,
  32'h3e0dbead /* (11, 24, 20) */,
  32'h3da58a7f /* (7, 24, 20) */,
  32'h3d729483 /* (3, 24, 20) */,
  32'h3dbaaaa9 /* (31, 20, 20) */,
  32'h3de671da /* (27, 20, 20) */,
  32'h3e3c290c /* (23, 20, 20) */,
  32'h3eaa0eb2 /* (19, 20, 20) */,
  32'h3ebf3a63 /* (15, 20, 20) */,
  32'h3e80c082 /* (11, 20, 20) */,
  32'h3e0e8e1e /* (7, 20, 20) */,
  32'h3dc823b1 /* (3, 20, 20) */,
  32'h3dcf60c6 /* (31, 16, 20) */,
  32'h3e02cee2 /* (27, 16, 20) */,
  32'h3e5e82df /* (23, 16, 20) */,
  32'h3ed28b29 /* (19, 16, 20) */,
  32'h3ef1f40b /* (15, 16, 20) */,
  32'h3e9bce24 /* (11, 16, 20) */,
  32'h3e24eefd /* (7, 16, 20) */,
  32'h3de007f6 /* (3, 16, 20) */,
  32'h3dbaaaa9 /* (31, 12, 20) */,
  32'h3de671da /* (27, 12, 20) */,
  32'h3e3c290c /* (23, 12, 20) */,
  32'h3eaa0eb2 /* (19, 12, 20) */,
  32'h3ebf3a63 /* (15, 12, 20) */,
  32'h3e80c082 /* (11, 12, 20) */,
  32'h3e0e8e1e /* (7, 12, 20) */,
  32'h3dc823b1 /* (3, 12, 20) */,
  32'h3d649547 /* (31, 8, 20) */,
  32'h3d89129f /* (27, 8, 20) */,
  32'h3dd4c19e /* (23, 8, 20) */,
  32'h3e368e5b /* (19, 8, 20) */,
  32'h3e48a298 /* (15, 8, 20) */,
  32'h3e0dbead /* (11, 8, 20) */,
  32'h3da58a7f /* (7, 8, 20) */,
  32'h3d729483 /* (3, 8, 20) */,
  32'h3d27af27 /* (31, 4, 20) */,
  32'h3d431db1 /* (27, 4, 20) */,
  32'h3d902ce0 /* (23, 4, 20) */,
  32'h3dec6d9f /* (19, 4, 20) */,
  32'h3dff07bf /* (15, 4, 20) */,
  32'h3dbb90ec /* (11, 4, 20) */,
  32'h3d66108f /* (7, 4, 20) */,
  32'h3d30047a /* (3, 4, 20) */,
  32'h3d195f14 /* (31, 0, 20) */,
  32'h3d2ff16f /* (27, 0, 20) */,
  32'h3d7e6b4b /* (23, 0, 20) */,
  32'h3dccb681 /* (19, 0, 20) */,
  32'h3ddb309a /* (15, 0, 20) */,
  32'h3da3d600 /* (11, 0, 20) */,
  32'h3d4d39f8 /* (7, 0, 20) */,
  32'h3d202826 /* (3, 0, 20) */,
  32'h3d18708b /* (31, 28, 16) */,
  32'h3d3b5943 /* (27, 28, 16) */,
  32'h3d97bb42 /* (23, 28, 16) */,
  32'h3e07f264 /* (19, 28, 16) */,
  32'h3e18449a /* (15, 28, 16) */,
  32'h3dcebbc1 /* (11, 28, 16) */,
  32'h3d66e7bc /* (7, 28, 16) */,
  32'h3d232f37 /* (3, 28, 16) */,
  32'h3d656b11 /* (31, 24, 16) */,
  32'h3d8eb3bf /* (27, 24, 16) */,
  32'h3dec5cc9 /* (23, 24, 16) */,
  32'h3e58f4b1 /* (19, 24, 16) */,
  32'h3e75b861 /* (15, 24, 16) */,
  32'h3e2301df /* (11, 24, 16) */,
  32'h3db1ba44 /* (7, 24, 16) */,
  32'h3d76a38f /* (3, 24, 16) */,
  32'h3dcf60c6 /* (31, 20, 16) */,
  32'h3e02cee2 /* (27, 20, 16) */,
  32'h3e5e82df /* (23, 20, 16) */,
  32'h3ed28b29 /* (19, 20, 16) */,
  32'h3ef1f40b /* (15, 20, 16) */,
  32'h3e9bce24 /* (11, 20, 16) */,
  32'h3e24eefd /* (7, 20, 16) */,
  32'h3de007f6 /* (3, 20, 16) */,
  32'h3df9e164 /* (31, 16, 16) */,
  32'h3e1f95bf /* (27, 16, 16) */,
  32'h3e8b1bdf /* (23, 16, 16) */,
  32'h3f079668 /* (19, 16, 16) */,
  32'h3f1e253a /* (15, 16, 16) */,
  32'h3ec5ad99 /* (11, 16, 16) */,
  32'h3e4b7c7a /* (7, 16, 16) */,
  32'h3e078d5a /* (3, 16, 16) */,
  32'h3dcf60c6 /* (31, 12, 16) */,
  32'h3e02cee2 /* (27, 12, 16) */,
  32'h3e5e82df /* (23, 12, 16) */,
  32'h3ed28b29 /* (19, 12, 16) */,
  32'h3ef1f40b /* (15, 12, 16) */,
  32'h3e9bce24 /* (11, 12, 16) */,
  32'h3e24eefd /* (7, 12, 16) */,
  32'h3de007f6 /* (3, 12, 16) */,
  32'h3d656b11 /* (31, 8, 16) */,
  32'h3d8eb3bf /* (27, 8, 16) */,
  32'h3dec5cc9 /* (23, 8, 16) */,
  32'h3e58f4b1 /* (19, 8, 16) */,
  32'h3e75b861 /* (15, 8, 16) */,
  32'h3e2301df /* (11, 8, 16) */,
  32'h3db1ba44 /* (7, 8, 16) */,
  32'h3d76a38f /* (3, 8, 16) */,
  32'h3d18708b /* (31, 4, 16) */,
  32'h3d3b5943 /* (27, 4, 16) */,
  32'h3d97bb42 /* (23, 4, 16) */,
  32'h3e07f264 /* (19, 4, 16) */,
  32'h3e18449a /* (15, 4, 16) */,
  32'h3dcebbc1 /* (11, 4, 16) */,
  32'h3d66e7bc /* (7, 4, 16) */,
  32'h3d232f37 /* (3, 4, 16) */,
  32'h3d0563b9 /* (31, 0, 16) */,
  32'h3d231d8f /* (27, 0, 16) */,
  32'h3d82ec35 /* (23, 0, 16) */,
  32'h3de8675d /* (19, 0, 16) */,
  32'h3e019a4f /* (15, 0, 16) */,
  32'h3db1860e /* (11, 0, 16) */,
  32'h3d482f92 /* (7, 0, 16) */,
  32'h3d0e89f8 /* (3, 0, 16) */,
  32'h3d27af27 /* (31, 28, 12) */,
  32'h3d431db1 /* (27, 28, 12) */,
  32'h3d902ce0 /* (23, 28, 12) */,
  32'h3dec6d9f /* (19, 28, 12) */,
  32'h3dff07bf /* (15, 28, 12) */,
  32'h3dbb90ec /* (11, 28, 12) */,
  32'h3d66108f /* (7, 28, 12) */,
  32'h3d30047a /* (3, 28, 12) */,
  32'h3d649547 /* (31, 24, 12) */,
  32'h3d89129f /* (27, 24, 12) */,
  32'h3dd4c19e /* (23, 24, 12) */,
  32'h3e368e5b /* (19, 24, 12) */,
  32'h3e48a298 /* (15, 24, 12) */,
  32'h3e0dbead /* (11, 24, 12) */,
  32'h3da58a7f /* (7, 24, 12) */,
  32'h3d729483 /* (3, 24, 12) */,
  32'h3dbaaaa9 /* (31, 20, 12) */,
  32'h3de671da /* (27, 20, 12) */,
  32'h3e3c290c /* (23, 20, 12) */,
  32'h3eaa0eb2 /* (19, 20, 12) */,
  32'h3ebf3a63 /* (15, 20, 12) */,
  32'h3e80c082 /* (11, 20, 12) */,
  32'h3e0e8e1e /* (7, 20, 12) */,
  32'h3dc823b1 /* (3, 20, 12) */,
  32'h3dcf60c6 /* (31, 16, 12) */,
  32'h3e02cee2 /* (27, 16, 12) */,
  32'h3e5e82df /* (23, 16, 12) */,
  32'h3ed28b29 /* (19, 16, 12) */,
  32'h3ef1f40b /* (15, 16, 12) */,
  32'h3e9bce24 /* (11, 16, 12) */,
  32'h3e24eefd /* (7, 16, 12) */,
  32'h3de007f6 /* (3, 16, 12) */,
  32'h3dbaaaa9 /* (31, 12, 12) */,
  32'h3de671da /* (27, 12, 12) */,
  32'h3e3c290c /* (23, 12, 12) */,
  32'h3eaa0eb2 /* (19, 12, 12) */,
  32'h3ebf3a63 /* (15, 12, 12) */,
  32'h3e80c082 /* (11, 12, 12) */,
  32'h3e0e8e1e /* (7, 12, 12) */,
  32'h3dc823b1 /* (3, 12, 12) */,
  32'h3d649547 /* (31, 8, 12) */,
  32'h3d89129f /* (27, 8, 12) */,
  32'h3dd4c19e /* (23, 8, 12) */,
  32'h3e368e5b /* (19, 8, 12) */,
  32'h3e48a298 /* (15, 8, 12) */,
  32'h3e0dbead /* (11, 8, 12) */,
  32'h3da58a7f /* (7, 8, 12) */,
  32'h3d729483 /* (3, 8, 12) */,
  32'h3d27af27 /* (31, 4, 12) */,
  32'h3d431db1 /* (27, 4, 12) */,
  32'h3d902ce0 /* (23, 4, 12) */,
  32'h3dec6d9f /* (19, 4, 12) */,
  32'h3dff07bf /* (15, 4, 12) */,
  32'h3dbb90ec /* (11, 4, 12) */,
  32'h3d66108f /* (7, 4, 12) */,
  32'h3d30047a /* (3, 4, 12) */,
  32'h3d195f14 /* (31, 0, 12) */,
  32'h3d2ff16f /* (27, 0, 12) */,
  32'h3d7e6b4b /* (23, 0, 12) */,
  32'h3dccb681 /* (19, 0, 12) */,
  32'h3ddb309a /* (15, 0, 12) */,
  32'h3da3d600 /* (11, 0, 12) */,
  32'h3d4d39f8 /* (7, 0, 12) */,
  32'h3d202826 /* (3, 0, 12) */,
  32'h3d139499 /* (31, 28, 8) */,
  32'h3d183845 /* (27, 28, 8) */,
  32'h3d3f1eea /* (23, 28, 8) */,
  32'h3d8a5278 /* (19, 28, 8) */,
  32'h3d8e8b3a /* (15, 28, 8) */,
  32'h3d683712 /* (11, 28, 8) */,
  32'h3d250b86 /* (7, 28, 8) */,
  32'h3d13fed6 /* (3, 28, 8) */,
  32'h3d23fb6f /* (31, 24, 8) */,
  32'h3d38dbff /* (27, 24, 8) */,
  32'h3d824402 /* (23, 24, 8) */,
  32'h3dcd36cb /* (19, 24, 8) */,
  32'h3dd9f1d0 /* (15, 24, 8) */,
  32'h3da5dafd /* (11, 24, 8) */,
  32'h3d54dbd1 /* (7, 24, 8) */,
  32'h3d2a2238 /* (3, 24, 8) */,
  32'h3d649547 /* (31, 20, 8) */,
  32'h3d89129f /* (27, 20, 8) */,
  32'h3dd4c19e /* (23, 20, 8) */,
  32'h3e368e5b /* (19, 20, 8) */,
  32'h3e48a298 /* (15, 20, 8) */,
  32'h3e0dbead /* (11, 20, 8) */,
  32'h3da58a7f /* (7, 20, 8) */,
  32'h3d729483 /* (3, 20, 8) */,
  32'h3d656b11 /* (31, 16, 8) */,
  32'h3d8eb3bf /* (27, 16, 8) */,
  32'h3dec5cc9 /* (23, 16, 8) */,
  32'h3e58f4b1 /* (19, 16, 8) */,
  32'h3e75b861 /* (15, 16, 8) */,
  32'h3e2301df /* (11, 16, 8) */,
  32'h3db1ba44 /* (7, 16, 8) */,
  32'h3d76a38f /* (3, 16, 8) */,
  32'h3d649547 /* (31, 12, 8) */,
  32'h3d89129f /* (27, 12, 8) */,
  32'h3dd4c19e /* (23, 12, 8) */,
  32'h3e368e5b /* (19, 12, 8) */,
  32'h3e48a298 /* (15, 12, 8) */,
  32'h3e0dbead /* (11, 12, 8) */,
  32'h3da58a7f /* (7, 12, 8) */,
  32'h3d729483 /* (3, 12, 8) */,
  32'h3d23fb6f /* (31, 8, 8) */,
  32'h3d38dbff /* (27, 8, 8) */,
  32'h3d824402 /* (23, 8, 8) */,
  32'h3dcd36cb /* (19, 8, 8) */,
  32'h3dd9f1d0 /* (15, 8, 8) */,
  32'h3da5dafd /* (11, 8, 8) */,
  32'h3d54dbd1 /* (7, 8, 8) */,
  32'h3d2a2238 /* (3, 8, 8) */,
  32'h3d139499 /* (31, 4, 8) */,
  32'h3d183845 /* (27, 4, 8) */,
  32'h3d3f1eea /* (23, 4, 8) */,
  32'h3d8a5278 /* (19, 4, 8) */,
  32'h3d8e8b3a /* (15, 4, 8) */,
  32'h3d683712 /* (11, 4, 8) */,
  32'h3d250b86 /* (7, 4, 8) */,
  32'h3d13fed6 /* (3, 4, 8) */,
  32'h3d177e6a /* (31, 0, 8) */,
  32'h3d13eed3 /* (27, 0, 8) */,
  32'h3d2eceba /* (23, 0, 8) */,
  32'h3d7388b1 /* (19, 0, 8) */,
  32'h3d77d78b /* (15, 0, 8) */,
  32'h3d4fd499 /* (11, 0, 8) */,
  32'h3d1b34b2 /* (7, 0, 8) */,
  32'h3d14a194 /* (3, 0, 8) */,
  32'h3d4cb45d /* (31, 28, 4) */,
  32'h3d1e7527 /* (27, 28, 4) */,
  32'h3d19e157 /* (23, 28, 4) */,
  32'h3d41aa67 /* (19, 28, 4) */,
  32'h3d3f317e /* (15, 28, 4) */,
  32'h3d2c64eb /* (11, 28, 4) */,
  32'h3d148979 /* (7, 28, 4) */,
  32'h3d358b49 /* (3, 28, 4) */,
  32'h3d139499 /* (31, 24, 4) */,
  32'h3d183845 /* (27, 24, 4) */,
  32'h3d3f1eea /* (23, 24, 4) */,
  32'h3d8a5278 /* (19, 24, 4) */,
  32'h3d8e8b3a /* (15, 24, 4) */,
  32'h3d683712 /* (11, 24, 4) */,
  32'h3d250b86 /* (7, 24, 4) */,
  32'h3d13fed6 /* (3, 24, 4) */,
  32'h3d27af27 /* (31, 20, 4) */,
  32'h3d431db1 /* (27, 20, 4) */,
  32'h3d902ce0 /* (23, 20, 4) */,
  32'h3dec6d9f /* (19, 20, 4) */,
  32'h3dff07bf /* (15, 20, 4) */,
  32'h3dbb90ec /* (11, 20, 4) */,
  32'h3d66108f /* (7, 20, 4) */,
  32'h3d30047a /* (3, 20, 4) */,
  32'h3d18708b /* (31, 16, 4) */,
  32'h3d3b5943 /* (27, 16, 4) */,
  32'h3d97bb42 /* (23, 16, 4) */,
  32'h3e07f264 /* (19, 16, 4) */,
  32'h3e18449a /* (15, 16, 4) */,
  32'h3dcebbc1 /* (11, 16, 4) */,
  32'h3d66e7bc /* (7, 16, 4) */,
  32'h3d232f37 /* (3, 16, 4) */,
  32'h3d27af27 /* (31, 12, 4) */,
  32'h3d431db1 /* (27, 12, 4) */,
  32'h3d902ce0 /* (23, 12, 4) */,
  32'h3dec6d9f /* (19, 12, 4) */,
  32'h3dff07bf /* (15, 12, 4) */,
  32'h3dbb90ec /* (11, 12, 4) */,
  32'h3d66108f /* (7, 12, 4) */,
  32'h3d30047a /* (3, 12, 4) */,
  32'h3d139499 /* (31, 8, 4) */,
  32'h3d183845 /* (27, 8, 4) */,
  32'h3d3f1eea /* (23, 8, 4) */,
  32'h3d8a5278 /* (19, 8, 4) */,
  32'h3d8e8b3a /* (15, 8, 4) */,
  32'h3d683712 /* (11, 8, 4) */,
  32'h3d250b86 /* (7, 8, 4) */,
  32'h3d13fed6 /* (3, 8, 4) */,
  32'h3d4cb45d /* (31, 4, 4) */,
  32'h3d1e7527 /* (27, 4, 4) */,
  32'h3d19e157 /* (23, 4, 4) */,
  32'h3d41aa67 /* (19, 4, 4) */,
  32'h3d3f317e /* (15, 4, 4) */,
  32'h3d2c64eb /* (11, 4, 4) */,
  32'h3d148979 /* (7, 4, 4) */,
  32'h3d358b49 /* (3, 4, 4) */,
  32'h3da3aa58 /* (31, 0, 4) */,
  32'h3d3577a5 /* (27, 0, 4) */,
  32'h3d13aacb /* (23, 0, 4) */,
  32'h3d2d543a /* (19, 0, 4) */,
  32'h3d27f384 /* (15, 0, 4) */,
  32'h3d1e982c /* (11, 0, 4) */,
  32'h3d1879c9 /* (7, 0, 4) */,
  32'h3d7541a2 /* (3, 0, 4) */,
  32'h3da3aa58 /* (31, 28, 0) */,
  32'h3d3577a5 /* (27, 28, 0) */,
  32'h3d13aacb /* (23, 28, 0) */,
  32'h3d2d543a /* (19, 28, 0) */,
  32'h3d27f384 /* (15, 28, 0) */,
  32'h3d1e982c /* (11, 28, 0) */,
  32'h3d1879c9 /* (7, 28, 0) */,
  32'h3d7541a2 /* (3, 28, 0) */,
  32'h3d177e6a /* (31, 24, 0) */,
  32'h3d13eed3 /* (27, 24, 0) */,
  32'h3d2eceba /* (23, 24, 0) */,
  32'h3d7388b1 /* (19, 24, 0) */,
  32'h3d77d78b /* (15, 24, 0) */,
  32'h3d4fd499 /* (11, 24, 0) */,
  32'h3d1b34b2 /* (7, 24, 0) */,
  32'h3d14a194 /* (3, 24, 0) */,
  32'h3d195f14 /* (31, 20, 0) */,
  32'h3d2ff16f /* (27, 20, 0) */,
  32'h3d7e6b4b /* (23, 20, 0) */,
  32'h3dccb681 /* (19, 20, 0) */,
  32'h3ddb309a /* (15, 20, 0) */,
  32'h3da3d600 /* (11, 20, 0) */,
  32'h3d4d39f8 /* (7, 20, 0) */,
  32'h3d202826 /* (3, 20, 0) */,
  32'h3d0563b9 /* (31, 16, 0) */,
  32'h3d231d8f /* (27, 16, 0) */,
  32'h3d82ec35 /* (23, 16, 0) */,
  32'h3de8675d /* (19, 16, 0) */,
  32'h3e019a4f /* (15, 16, 0) */,
  32'h3db1860e /* (11, 16, 0) */,
  32'h3d482f92 /* (7, 16, 0) */,
  32'h3d0e89f8 /* (3, 16, 0) */,
  32'h3d195f14 /* (31, 12, 0) */,
  32'h3d2ff16f /* (27, 12, 0) */,
  32'h3d7e6b4b /* (23, 12, 0) */,
  32'h3dccb681 /* (19, 12, 0) */,
  32'h3ddb309a /* (15, 12, 0) */,
  32'h3da3d600 /* (11, 12, 0) */,
  32'h3d4d39f8 /* (7, 12, 0) */,
  32'h3d202826 /* (3, 12, 0) */,
  32'h3d177e6a /* (31, 8, 0) */,
  32'h3d13eed3 /* (27, 8, 0) */,
  32'h3d2eceba /* (23, 8, 0) */,
  32'h3d7388b1 /* (19, 8, 0) */,
  32'h3d77d78b /* (15, 8, 0) */,
  32'h3d4fd499 /* (11, 8, 0) */,
  32'h3d1b34b2 /* (7, 8, 0) */,
  32'h3d14a194 /* (3, 8, 0) */,
  32'h3da3aa58 /* (31, 4, 0) */,
  32'h3d3577a5 /* (27, 4, 0) */,
  32'h3d13aacb /* (23, 4, 0) */,
  32'h3d2d543a /* (19, 4, 0) */,
  32'h3d27f384 /* (15, 4, 0) */,
  32'h3d1e982c /* (11, 4, 0) */,
  32'h3d1879c9 /* (7, 4, 0) */,
  32'h3d7541a2 /* (3, 4, 0) */,
  32'h3f8f3ec8 /* (31, 0, 0) */,
  32'h3d75271a /* (27, 0, 0) */,
  32'h3d11ab15 /* (23, 0, 0) */,
  32'h3d1c4c09 /* (19, 0, 0) */,
  32'h3d14300c /* (15, 0, 0) */,
  32'h3d13eab3 /* (11, 0, 0) */,
  32'h3d269d45 /* (7, 0, 0) */,
  32'h3e0c4c59 /* (3, 0, 0) */,
  32'h3d429928 /* (30, 28, 28) */,
  32'h3d1796af /* (26, 28, 28) */,
  32'h3d21d2a4 /* (22, 28, 28) */,
  32'h3d456b70 /* (18, 28, 28) */,
  32'h3d456b70 /* (14, 28, 28) */,
  32'h3d21d2a4 /* (10, 28, 28) */,
  32'h3d1796af /* (6, 28, 28) */,
  32'h3d429928 /* (2, 28, 28) */,
  32'h3d139519 /* (30, 24, 28) */,
  32'h3d1d3fef /* (26, 24, 28) */,
  32'h3d51ff4c /* (22, 24, 28) */,
  32'h3d904c26 /* (18, 24, 28) */,
  32'h3d904c26 /* (14, 24, 28) */,
  32'h3d51ff4c /* (10, 24, 28) */,
  32'h3d1d3fef /* (6, 24, 28) */,
  32'h3d139519 /* (2, 24, 28) */,
  32'h3d2ab74a /* (30, 20, 28) */,
  32'h3d522ea6 /* (26, 20, 28) */,
  32'h3da42ada /* (22, 20, 28) */,
  32'h3dfca6c8 /* (18, 20, 28) */,
  32'h3dfca6c8 /* (14, 20, 28) */,
  32'h3da42ada /* (10, 20, 28) */,
  32'h3d522ea6 /* (6, 20, 28) */,
  32'h3d2ab74a /* (2, 20, 28) */,
  32'h3d1c5e8a /* (30, 16, 28) */,
  32'h3d4e2dc2 /* (26, 16, 28) */,
  32'h3db0df4f /* (22, 16, 28) */,
  32'h3e1420e4 /* (18, 16, 28) */,
  32'h3e1420e4 /* (14, 16, 28) */,
  32'h3db0df4f /* (10, 16, 28) */,
  32'h3d4e2dc2 /* (6, 16, 28) */,
  32'h3d1c5e8a /* (2, 16, 28) */,
  32'h3d2ab74a /* (30, 12, 28) */,
  32'h3d522ea6 /* (26, 12, 28) */,
  32'h3da42ada /* (22, 12, 28) */,
  32'h3dfca6c8 /* (18, 12, 28) */,
  32'h3dfca6c8 /* (14, 12, 28) */,
  32'h3da42ada /* (10, 12, 28) */,
  32'h3d522ea6 /* (6, 12, 28) */,
  32'h3d2ab74a /* (2, 12, 28) */,
  32'h3d139519 /* (30, 8, 28) */,
  32'h3d1d3fef /* (26, 8, 28) */,
  32'h3d51ff4c /* (22, 8, 28) */,
  32'h3d904c26 /* (18, 8, 28) */,
  32'h3d904c26 /* (14, 8, 28) */,
  32'h3d51ff4c /* (10, 8, 28) */,
  32'h3d1d3fef /* (6, 8, 28) */,
  32'h3d139519 /* (2, 8, 28) */,
  32'h3d429928 /* (30, 4, 28) */,
  32'h3d1796af /* (26, 4, 28) */,
  32'h3d21d2a4 /* (22, 4, 28) */,
  32'h3d456b70 /* (18, 4, 28) */,
  32'h3d456b70 /* (14, 4, 28) */,
  32'h3d21d2a4 /* (10, 4, 28) */,
  32'h3d1796af /* (6, 4, 28) */,
  32'h3d429928 /* (2, 4, 28) */,
  32'h3d90451b /* (30, 0, 28) */,
  32'h3d234ae8 /* (26, 0, 28) */,
  32'h3d17b006 /* (22, 0, 28) */,
  32'h3d2ee5c8 /* (18, 0, 28) */,
  32'h3d2ee5c8 /* (14, 0, 28) */,
  32'h3d17b006 /* (10, 0, 28) */,
  32'h3d234ae8 /* (6, 0, 28) */,
  32'h3d90451b /* (2, 0, 28) */,
  32'h3d139519 /* (30, 28, 24) */,
  32'h3d1d3fef /* (26, 28, 24) */,
  32'h3d51ff4c /* (22, 28, 24) */,
  32'h3d904c26 /* (18, 28, 24) */,
  32'h3d904c26 /* (14, 28, 24) */,
  32'h3d51ff4c /* (10, 28, 24) */,
  32'h3d1d3fef /* (6, 28, 24) */,
  32'h3d139519 /* (2, 28, 24) */,
  32'h3d263161 /* (30, 24, 24) */,
  32'h3d44d2c5 /* (26, 24, 24) */,
  32'h3d92b00e /* (22, 24, 24) */,
  32'h3dd9849b /* (18, 24, 24) */,
  32'h3dd9849b /* (14, 24, 24) */,
  32'h3d92b00e /* (10, 24, 24) */,
  32'h3d44d2c5 /* (6, 24, 24) */,
  32'h3d263161 /* (2, 24, 24) */,
  32'h3d69b2a3 /* (30, 20, 24) */,
  32'h3d95625b /* (26, 20, 24) */,
  32'h3df53c17 /* (22, 20, 24) */,
  32'h3e44fc23 /* (18, 20, 24) */,
  32'h3e44fc23 /* (14, 20, 24) */,
  32'h3df53c17 /* (10, 20, 24) */,
  32'h3d95625b /* (6, 20, 24) */,
  32'h3d69b2a3 /* (2, 20, 24) */,
  32'h3d6bb726 /* (30, 16, 24) */,
  32'h3d9dd43f /* (26, 16, 24) */,
  32'h3e0a9c46 /* (22, 16, 24) */,
  32'h3e6dbe20 /* (18, 16, 24) */,
  32'h3e6dbe20 /* (14, 16, 24) */,
  32'h3e0a9c46 /* (10, 16, 24) */,
  32'h3d9dd43f /* (6, 16, 24) */,
  32'h3d6bb726 /* (2, 16, 24) */,
  32'h3d69b2a3 /* (30, 12, 24) */,
  32'h3d95625b /* (26, 12, 24) */,
  32'h3df53c17 /* (22, 12, 24) */,
  32'h3e44fc23 /* (18, 12, 24) */,
  32'h3e44fc23 /* (14, 12, 24) */,
  32'h3df53c17 /* (10, 12, 24) */,
  32'h3d95625b /* (6, 12, 24) */,
  32'h3d69b2a3 /* (2, 12, 24) */,
  32'h3d263161 /* (30, 8, 24) */,
  32'h3d44d2c5 /* (26, 8, 24) */,
  32'h3d92b00e /* (22, 8, 24) */,
  32'h3dd9849b /* (18, 8, 24) */,
  32'h3dd9849b /* (14, 8, 24) */,
  32'h3d92b00e /* (10, 8, 24) */,
  32'h3d44d2c5 /* (6, 8, 24) */,
  32'h3d263161 /* (2, 8, 24) */,
  32'h3d139519 /* (30, 4, 24) */,
  32'h3d1d3fef /* (26, 4, 24) */,
  32'h3d51ff4c /* (22, 4, 24) */,
  32'h3d904c26 /* (18, 4, 24) */,
  32'h3d904c26 /* (14, 4, 24) */,
  32'h3d51ff4c /* (10, 4, 24) */,
  32'h3d1d3fef /* (6, 4, 24) */,
  32'h3d139519 /* (2, 4, 24) */,
  32'h3d162cf4 /* (30, 0, 24) */,
  32'h3d164277 /* (26, 0, 24) */,
  32'h3d3ddc84 /* (22, 0, 24) */,
  32'h3d7c5be6 /* (18, 0, 24) */,
  32'h3d7c5be6 /* (14, 0, 24) */,
  32'h3d3ddc84 /* (10, 0, 24) */,
  32'h3d164277 /* (6, 0, 24) */,
  32'h3d162cf4 /* (2, 0, 24) */,
  32'h3d2ab74a /* (30, 28, 20) */,
  32'h3d522ea6 /* (26, 28, 20) */,
  32'h3da42ada /* (22, 28, 20) */,
  32'h3dfca6c8 /* (18, 28, 20) */,
  32'h3dfca6c8 /* (14, 28, 20) */,
  32'h3da42ada /* (10, 28, 20) */,
  32'h3d522ea6 /* (6, 28, 20) */,
  32'h3d2ab74a /* (2, 28, 20) */,
  32'h3d69b2a3 /* (30, 24, 20) */,
  32'h3d95625b /* (26, 24, 20) */,
  32'h3df53c17 /* (22, 24, 20) */,
  32'h3e44fc23 /* (18, 24, 20) */,
  32'h3e44fc23 /* (14, 24, 20) */,
  32'h3df53c17 /* (10, 24, 20) */,
  32'h3d95625b /* (6, 24, 20) */,
  32'h3d69b2a3 /* (2, 24, 20) */,
  32'h3dbf980c /* (30, 20, 20) */,
  32'h3dfe11f4 /* (26, 20, 20) */,
  32'h3e5bd2f1 /* (22, 20, 20) */,
  32'h3eb9abaa /* (18, 20, 20) */,
  32'h3eb9abaa /* (14, 20, 20) */,
  32'h3e5bd2f1 /* (10, 20, 20) */,
  32'h3dfe11f4 /* (6, 20, 20) */,
  32'h3dbf980c /* (2, 20, 20) */,
  32'h3dd576ed /* (30, 16, 20) */,
  32'h3e11854b /* (26, 16, 20) */,
  32'h3e837a14 /* (22, 16, 20) */,
  32'h3ee86d0e /* (18, 16, 20) */,
  32'h3ee86d0e /* (14, 16, 20) */,
  32'h3e837a14 /* (10, 16, 20) */,
  32'h3e11854b /* (6, 16, 20) */,
  32'h3dd576ed /* (2, 16, 20) */,
  32'h3dbf980c /* (30, 12, 20) */,
  32'h3dfe11f4 /* (26, 12, 20) */,
  32'h3e5bd2f1 /* (22, 12, 20) */,
  32'h3eb9abaa /* (18, 12, 20) */,
  32'h3eb9abaa /* (14, 12, 20) */,
  32'h3e5bd2f1 /* (10, 12, 20) */,
  32'h3dfe11f4 /* (6, 12, 20) */,
  32'h3dbf980c /* (2, 12, 20) */,
  32'h3d69b2a3 /* (30, 8, 20) */,
  32'h3d95625b /* (26, 8, 20) */,
  32'h3df53c17 /* (22, 8, 20) */,
  32'h3e44fc23 /* (18, 8, 20) */,
  32'h3e44fc23 /* (14, 8, 20) */,
  32'h3df53c17 /* (10, 8, 20) */,
  32'h3d95625b /* (6, 8, 20) */,
  32'h3d69b2a3 /* (2, 8, 20) */,
  32'h3d2ab74a /* (30, 4, 20) */,
  32'h3d522ea6 /* (26, 4, 20) */,
  32'h3da42ada /* (22, 4, 20) */,
  32'h3dfca6c8 /* (18, 4, 20) */,
  32'h3dfca6c8 /* (14, 4, 20) */,
  32'h3da42ada /* (10, 4, 20) */,
  32'h3d522ea6 /* (6, 4, 20) */,
  32'h3d2ab74a /* (2, 4, 20) */,
  32'h3d1bd472 /* (30, 0, 20) */,
  32'h3d3c86f4 /* (26, 0, 20) */,
  32'h3d9019ab /* (22, 0, 20) */,
  32'h3dd9ea44 /* (18, 0, 20) */,
  32'h3dd9ea44 /* (14, 0, 20) */,
  32'h3d9019ab /* (10, 0, 20) */,
  32'h3d3c86f4 /* (6, 0, 20) */,
  32'h3d1bd472 /* (2, 0, 20) */,
  32'h3d1c5e8a /* (30, 28, 16) */,
  32'h3d4e2dc2 /* (26, 28, 16) */,
  32'h3db0df4f /* (22, 28, 16) */,
  32'h3e1420e4 /* (18, 28, 16) */,
  32'h3e1420e4 /* (14, 28, 16) */,
  32'h3db0df4f /* (10, 28, 16) */,
  32'h3d4e2dc2 /* (6, 28, 16) */,
  32'h3d1c5e8a /* (2, 28, 16) */,
  32'h3d6bb726 /* (30, 24, 16) */,
  32'h3d9dd43f /* (26, 24, 16) */,
  32'h3e0a9c46 /* (22, 24, 16) */,
  32'h3e6dbe20 /* (18, 24, 16) */,
  32'h3e6dbe20 /* (14, 24, 16) */,
  32'h3e0a9c46 /* (10, 24, 16) */,
  32'h3d9dd43f /* (6, 24, 16) */,
  32'h3d6bb726 /* (2, 24, 16) */,
  32'h3dd576ed /* (30, 20, 16) */,
  32'h3e11854b /* (26, 20, 16) */,
  32'h3e837a14 /* (22, 20, 16) */,
  32'h3ee86d0e /* (18, 20, 16) */,
  32'h3ee86d0e /* (14, 20, 16) */,
  32'h3e837a14 /* (10, 20, 16) */,
  32'h3e11854b /* (6, 20, 16) */,
  32'h3dd576ed /* (2, 20, 16) */,
  32'h3e00d0e8 /* (30, 16, 16) */,
  32'h3e327927 /* (26, 16, 16) */,
  32'h3ea594bb /* (22, 16, 16) */,
  32'h3f16cd97 /* (18, 16, 16) */,
  32'h3f16cd97 /* (14, 16, 16) */,
  32'h3ea594bb /* (10, 16, 16) */,
  32'h3e327927 /* (6, 16, 16) */,
  32'h3e00d0e8 /* (2, 16, 16) */,
  32'h3dd576ed /* (30, 12, 16) */,
  32'h3e11854b /* (26, 12, 16) */,
  32'h3e837a14 /* (22, 12, 16) */,
  32'h3ee86d0e /* (18, 12, 16) */,
  32'h3ee86d0e /* (14, 12, 16) */,
  32'h3e837a14 /* (10, 12, 16) */,
  32'h3e11854b /* (6, 12, 16) */,
  32'h3dd576ed /* (2, 12, 16) */,
  32'h3d6bb726 /* (30, 8, 16) */,
  32'h3d9dd43f /* (26, 8, 16) */,
  32'h3e0a9c46 /* (22, 8, 16) */,
  32'h3e6dbe20 /* (18, 8, 16) */,
  32'h3e6dbe20 /* (14, 8, 16) */,
  32'h3e0a9c46 /* (10, 8, 16) */,
  32'h3d9dd43f /* (6, 8, 16) */,
  32'h3d6bb726 /* (2, 8, 16) */,
  32'h3d1c5e8a /* (30, 4, 16) */,
  32'h3d4e2dc2 /* (26, 4, 16) */,
  32'h3db0df4f /* (22, 4, 16) */,
  32'h3e1420e4 /* (18, 4, 16) */,
  32'h3e1420e4 /* (14, 4, 16) */,
  32'h3db0df4f /* (10, 4, 16) */,
  32'h3d4e2dc2 /* (6, 4, 16) */,
  32'h3d1c5e8a /* (2, 4, 16) */,
  32'h3d08bc50 /* (30, 0, 16) */,
  32'h3d332545 /* (26, 0, 16) */,
  32'h3d983f17 /* (22, 0, 16) */,
  32'h3dfcae00 /* (18, 0, 16) */,
  32'h3dfcae00 /* (14, 0, 16) */,
  32'h3d983f17 /* (10, 0, 16) */,
  32'h3d332545 /* (6, 0, 16) */,
  32'h3d08bc50 /* (2, 0, 16) */,
  32'h3d2ab74a /* (30, 28, 12) */,
  32'h3d522ea6 /* (26, 28, 12) */,
  32'h3da42ada /* (22, 28, 12) */,
  32'h3dfca6c8 /* (18, 28, 12) */,
  32'h3dfca6c8 /* (14, 28, 12) */,
  32'h3da42ada /* (10, 28, 12) */,
  32'h3d522ea6 /* (6, 28, 12) */,
  32'h3d2ab74a /* (2, 28, 12) */,
  32'h3d69b2a3 /* (30, 24, 12) */,
  32'h3d95625b /* (26, 24, 12) */,
  32'h3df53c17 /* (22, 24, 12) */,
  32'h3e44fc23 /* (18, 24, 12) */,
  32'h3e44fc23 /* (14, 24, 12) */,
  32'h3df53c17 /* (10, 24, 12) */,
  32'h3d95625b /* (6, 24, 12) */,
  32'h3d69b2a3 /* (2, 24, 12) */,
  32'h3dbf980c /* (30, 20, 12) */,
  32'h3dfe11f4 /* (26, 20, 12) */,
  32'h3e5bd2f1 /* (22, 20, 12) */,
  32'h3eb9abaa /* (18, 20, 12) */,
  32'h3eb9abaa /* (14, 20, 12) */,
  32'h3e5bd2f1 /* (10, 20, 12) */,
  32'h3dfe11f4 /* (6, 20, 12) */,
  32'h3dbf980c /* (2, 20, 12) */,
  32'h3dd576ed /* (30, 16, 12) */,
  32'h3e11854b /* (26, 16, 12) */,
  32'h3e837a14 /* (22, 16, 12) */,
  32'h3ee86d0e /* (18, 16, 12) */,
  32'h3ee86d0e /* (14, 16, 12) */,
  32'h3e837a14 /* (10, 16, 12) */,
  32'h3e11854b /* (6, 16, 12) */,
  32'h3dd576ed /* (2, 16, 12) */,
  32'h3dbf980c /* (30, 12, 12) */,
  32'h3dfe11f4 /* (26, 12, 12) */,
  32'h3e5bd2f1 /* (22, 12, 12) */,
  32'h3eb9abaa /* (18, 12, 12) */,
  32'h3eb9abaa /* (14, 12, 12) */,
  32'h3e5bd2f1 /* (10, 12, 12) */,
  32'h3dfe11f4 /* (6, 12, 12) */,
  32'h3dbf980c /* (2, 12, 12) */,
  32'h3d69b2a3 /* (30, 8, 12) */,
  32'h3d95625b /* (26, 8, 12) */,
  32'h3df53c17 /* (22, 8, 12) */,
  32'h3e44fc23 /* (18, 8, 12) */,
  32'h3e44fc23 /* (14, 8, 12) */,
  32'h3df53c17 /* (10, 8, 12) */,
  32'h3d95625b /* (6, 8, 12) */,
  32'h3d69b2a3 /* (2, 8, 12) */,
  32'h3d2ab74a /* (30, 4, 12) */,
  32'h3d522ea6 /* (26, 4, 12) */,
  32'h3da42ada /* (22, 4, 12) */,
  32'h3dfca6c8 /* (18, 4, 12) */,
  32'h3dfca6c8 /* (14, 4, 12) */,
  32'h3da42ada /* (10, 4, 12) */,
  32'h3d522ea6 /* (6, 4, 12) */,
  32'h3d2ab74a /* (2, 4, 12) */,
  32'h3d1bd472 /* (30, 0, 12) */,
  32'h3d3c86f4 /* (26, 0, 12) */,
  32'h3d9019ab /* (22, 0, 12) */,
  32'h3dd9ea44 /* (18, 0, 12) */,
  32'h3dd9ea44 /* (14, 0, 12) */,
  32'h3d9019ab /* (10, 0, 12) */,
  32'h3d3c86f4 /* (6, 0, 12) */,
  32'h3d1bd472 /* (2, 0, 12) */,
  32'h3d139519 /* (30, 28, 8) */,
  32'h3d1d3fef /* (26, 28, 8) */,
  32'h3d51ff4c /* (22, 28, 8) */,
  32'h3d904c26 /* (18, 28, 8) */,
  32'h3d904c26 /* (14, 28, 8) */,
  32'h3d51ff4c /* (10, 28, 8) */,
  32'h3d1d3fef /* (6, 28, 8) */,
  32'h3d139519 /* (2, 28, 8) */,
  32'h3d263161 /* (30, 24, 8) */,
  32'h3d44d2c5 /* (26, 24, 8) */,
  32'h3d92b00e /* (22, 24, 8) */,
  32'h3dd9849b /* (18, 24, 8) */,
  32'h3dd9849b /* (14, 24, 8) */,
  32'h3d92b00e /* (10, 24, 8) */,
  32'h3d44d2c5 /* (6, 24, 8) */,
  32'h3d263161 /* (2, 24, 8) */,
  32'h3d69b2a3 /* (30, 20, 8) */,
  32'h3d95625b /* (26, 20, 8) */,
  32'h3df53c17 /* (22, 20, 8) */,
  32'h3e44fc23 /* (18, 20, 8) */,
  32'h3e44fc23 /* (14, 20, 8) */,
  32'h3df53c17 /* (10, 20, 8) */,
  32'h3d95625b /* (6, 20, 8) */,
  32'h3d69b2a3 /* (2, 20, 8) */,
  32'h3d6bb726 /* (30, 16, 8) */,
  32'h3d9dd43f /* (26, 16, 8) */,
  32'h3e0a9c46 /* (22, 16, 8) */,
  32'h3e6dbe20 /* (18, 16, 8) */,
  32'h3e6dbe20 /* (14, 16, 8) */,
  32'h3e0a9c46 /* (10, 16, 8) */,
  32'h3d9dd43f /* (6, 16, 8) */,
  32'h3d6bb726 /* (2, 16, 8) */,
  32'h3d69b2a3 /* (30, 12, 8) */,
  32'h3d95625b /* (26, 12, 8) */,
  32'h3df53c17 /* (22, 12, 8) */,
  32'h3e44fc23 /* (18, 12, 8) */,
  32'h3e44fc23 /* (14, 12, 8) */,
  32'h3df53c17 /* (10, 12, 8) */,
  32'h3d95625b /* (6, 12, 8) */,
  32'h3d69b2a3 /* (2, 12, 8) */,
  32'h3d263161 /* (30, 8, 8) */,
  32'h3d44d2c5 /* (26, 8, 8) */,
  32'h3d92b00e /* (22, 8, 8) */,
  32'h3dd9849b /* (18, 8, 8) */,
  32'h3dd9849b /* (14, 8, 8) */,
  32'h3d92b00e /* (10, 8, 8) */,
  32'h3d44d2c5 /* (6, 8, 8) */,
  32'h3d263161 /* (2, 8, 8) */,
  32'h3d139519 /* (30, 4, 8) */,
  32'h3d1d3fef /* (26, 4, 8) */,
  32'h3d51ff4c /* (22, 4, 8) */,
  32'h3d904c26 /* (18, 4, 8) */,
  32'h3d904c26 /* (14, 4, 8) */,
  32'h3d51ff4c /* (10, 4, 8) */,
  32'h3d1d3fef /* (6, 4, 8) */,
  32'h3d139519 /* (2, 4, 8) */,
  32'h3d162cf4 /* (30, 0, 8) */,
  32'h3d164277 /* (26, 0, 8) */,
  32'h3d3ddc84 /* (22, 0, 8) */,
  32'h3d7c5be6 /* (18, 0, 8) */,
  32'h3d7c5be6 /* (14, 0, 8) */,
  32'h3d3ddc84 /* (10, 0, 8) */,
  32'h3d164277 /* (6, 0, 8) */,
  32'h3d162cf4 /* (2, 0, 8) */,
  32'h3d429928 /* (30, 28, 4) */,
  32'h3d1796af /* (26, 28, 4) */,
  32'h3d21d2a4 /* (22, 28, 4) */,
  32'h3d456b70 /* (18, 28, 4) */,
  32'h3d456b70 /* (14, 28, 4) */,
  32'h3d21d2a4 /* (10, 28, 4) */,
  32'h3d1796af /* (6, 28, 4) */,
  32'h3d429928 /* (2, 28, 4) */,
  32'h3d139519 /* (30, 24, 4) */,
  32'h3d1d3fef /* (26, 24, 4) */,
  32'h3d51ff4c /* (22, 24, 4) */,
  32'h3d904c26 /* (18, 24, 4) */,
  32'h3d904c26 /* (14, 24, 4) */,
  32'h3d51ff4c /* (10, 24, 4) */,
  32'h3d1d3fef /* (6, 24, 4) */,
  32'h3d139519 /* (2, 24, 4) */,
  32'h3d2ab74a /* (30, 20, 4) */,
  32'h3d522ea6 /* (26, 20, 4) */,
  32'h3da42ada /* (22, 20, 4) */,
  32'h3dfca6c8 /* (18, 20, 4) */,
  32'h3dfca6c8 /* (14, 20, 4) */,
  32'h3da42ada /* (10, 20, 4) */,
  32'h3d522ea6 /* (6, 20, 4) */,
  32'h3d2ab74a /* (2, 20, 4) */,
  32'h3d1c5e8a /* (30, 16, 4) */,
  32'h3d4e2dc2 /* (26, 16, 4) */,
  32'h3db0df4f /* (22, 16, 4) */,
  32'h3e1420e4 /* (18, 16, 4) */,
  32'h3e1420e4 /* (14, 16, 4) */,
  32'h3db0df4f /* (10, 16, 4) */,
  32'h3d4e2dc2 /* (6, 16, 4) */,
  32'h3d1c5e8a /* (2, 16, 4) */,
  32'h3d2ab74a /* (30, 12, 4) */,
  32'h3d522ea6 /* (26, 12, 4) */,
  32'h3da42ada /* (22, 12, 4) */,
  32'h3dfca6c8 /* (18, 12, 4) */,
  32'h3dfca6c8 /* (14, 12, 4) */,
  32'h3da42ada /* (10, 12, 4) */,
  32'h3d522ea6 /* (6, 12, 4) */,
  32'h3d2ab74a /* (2, 12, 4) */,
  32'h3d139519 /* (30, 8, 4) */,
  32'h3d1d3fef /* (26, 8, 4) */,
  32'h3d51ff4c /* (22, 8, 4) */,
  32'h3d904c26 /* (18, 8, 4) */,
  32'h3d904c26 /* (14, 8, 4) */,
  32'h3d51ff4c /* (10, 8, 4) */,
  32'h3d1d3fef /* (6, 8, 4) */,
  32'h3d139519 /* (2, 8, 4) */,
  32'h3d429928 /* (30, 4, 4) */,
  32'h3d1796af /* (26, 4, 4) */,
  32'h3d21d2a4 /* (22, 4, 4) */,
  32'h3d456b70 /* (18, 4, 4) */,
  32'h3d456b70 /* (14, 4, 4) */,
  32'h3d21d2a4 /* (10, 4, 4) */,
  32'h3d1796af /* (6, 4, 4) */,
  32'h3d429928 /* (2, 4, 4) */,
  32'h3d90451b /* (30, 0, 4) */,
  32'h3d234ae8 /* (26, 0, 4) */,
  32'h3d17b006 /* (22, 0, 4) */,
  32'h3d2ee5c8 /* (18, 0, 4) */,
  32'h3d2ee5c8 /* (14, 0, 4) */,
  32'h3d17b006 /* (10, 0, 4) */,
  32'h3d234ae8 /* (6, 0, 4) */,
  32'h3d90451b /* (2, 0, 4) */,
  32'h3d90451b /* (30, 28, 0) */,
  32'h3d234ae8 /* (26, 28, 0) */,
  32'h3d17b006 /* (22, 28, 0) */,
  32'h3d2ee5c8 /* (18, 28, 0) */,
  32'h3d2ee5c8 /* (14, 28, 0) */,
  32'h3d17b006 /* (10, 28, 0) */,
  32'h3d234ae8 /* (6, 28, 0) */,
  32'h3d90451b /* (2, 28, 0) */,
  32'h3d162cf4 /* (30, 24, 0) */,
  32'h3d164277 /* (26, 24, 0) */,
  32'h3d3ddc84 /* (22, 24, 0) */,
  32'h3d7c5be6 /* (18, 24, 0) */,
  32'h3d7c5be6 /* (14, 24, 0) */,
  32'h3d3ddc84 /* (10, 24, 0) */,
  32'h3d164277 /* (6, 24, 0) */,
  32'h3d162cf4 /* (2, 24, 0) */,
  32'h3d1bd472 /* (30, 20, 0) */,
  32'h3d3c86f4 /* (26, 20, 0) */,
  32'h3d9019ab /* (22, 20, 0) */,
  32'h3dd9ea44 /* (18, 20, 0) */,
  32'h3dd9ea44 /* (14, 20, 0) */,
  32'h3d9019ab /* (10, 20, 0) */,
  32'h3d3c86f4 /* (6, 20, 0) */,
  32'h3d1bd472 /* (2, 20, 0) */,
  32'h3d08bc50 /* (30, 16, 0) */,
  32'h3d332545 /* (26, 16, 0) */,
  32'h3d983f17 /* (22, 16, 0) */,
  32'h3dfcae00 /* (18, 16, 0) */,
  32'h3dfcae00 /* (14, 16, 0) */,
  32'h3d983f17 /* (10, 16, 0) */,
  32'h3d332545 /* (6, 16, 0) */,
  32'h3d08bc50 /* (2, 16, 0) */,
  32'h3d1bd472 /* (30, 12, 0) */,
  32'h3d3c86f4 /* (26, 12, 0) */,
  32'h3d9019ab /* (22, 12, 0) */,
  32'h3dd9ea44 /* (18, 12, 0) */,
  32'h3dd9ea44 /* (14, 12, 0) */,
  32'h3d9019ab /* (10, 12, 0) */,
  32'h3d3c86f4 /* (6, 12, 0) */,
  32'h3d1bd472 /* (2, 12, 0) */,
  32'h3d162cf4 /* (30, 8, 0) */,
  32'h3d164277 /* (26, 8, 0) */,
  32'h3d3ddc84 /* (22, 8, 0) */,
  32'h3d7c5be6 /* (18, 8, 0) */,
  32'h3d7c5be6 /* (14, 8, 0) */,
  32'h3d3ddc84 /* (10, 8, 0) */,
  32'h3d164277 /* (6, 8, 0) */,
  32'h3d162cf4 /* (2, 8, 0) */,
  32'h3d90451b /* (30, 4, 0) */,
  32'h3d234ae8 /* (26, 4, 0) */,
  32'h3d17b006 /* (22, 4, 0) */,
  32'h3d2ee5c8 /* (18, 4, 0) */,
  32'h3d2ee5c8 /* (14, 4, 0) */,
  32'h3d17b006 /* (10, 4, 0) */,
  32'h3d234ae8 /* (6, 4, 0) */,
  32'h3d90451b /* (2, 4, 0) */,
  32'h3e948d77 /* (30, 0, 0) */,
  32'h3d424b89 /* (26, 0, 0) */,
  32'h3d10f1da /* (22, 0, 0) */,
  32'h3d1bd51d /* (18, 0, 0) */,
  32'h3d1bd51d /* (14, 0, 0) */,
  32'h3d10f1da /* (10, 0, 0) */,
  32'h3d424b89 /* (6, 0, 0) */,
  32'h3e948d77 /* (2, 0, 0) */,
  32'h3d358b49 /* (29, 28, 28) */,
  32'h3d148979 /* (25, 28, 28) */,
  32'h3d2c64eb /* (21, 28, 28) */,
  32'h3d3f317e /* (17, 28, 28) */,
  32'h3d41aa67 /* (13, 28, 28) */,
  32'h3d19e157 /* (9, 28, 28) */,
  32'h3d1e7527 /* (5, 28, 28) */,
  32'h3d4cb45d /* (1, 28, 28) */,
  32'h3d13fed6 /* (29, 24, 28) */,
  32'h3d250b86 /* (25, 24, 28) */,
  32'h3d683712 /* (21, 24, 28) */,
  32'h3d8e8b3a /* (17, 24, 28) */,
  32'h3d8a5278 /* (13, 24, 28) */,
  32'h3d3f1eea /* (9, 24, 28) */,
  32'h3d183845 /* (5, 24, 28) */,
  32'h3d139499 /* (1, 24, 28) */,
  32'h3d30047a /* (29, 20, 28) */,
  32'h3d66108f /* (25, 20, 28) */,
  32'h3dbb90ec /* (21, 20, 28) */,
  32'h3dff07bf /* (17, 20, 28) */,
  32'h3dec6d9f /* (13, 20, 28) */,
  32'h3d902ce0 /* (9, 20, 28) */,
  32'h3d431db1 /* (5, 20, 28) */,
  32'h3d27af27 /* (1, 20, 28) */,
  32'h3d232f37 /* (29, 16, 28) */,
  32'h3d66e7bc /* (25, 16, 28) */,
  32'h3dcebbc1 /* (21, 16, 28) */,
  32'h3e18449a /* (17, 16, 28) */,
  32'h3e07f264 /* (13, 16, 28) */,
  32'h3d97bb42 /* (9, 16, 28) */,
  32'h3d3b5943 /* (5, 16, 28) */,
  32'h3d18708b /* (1, 16, 28) */,
  32'h3d30047a /* (29, 12, 28) */,
  32'h3d66108f /* (25, 12, 28) */,
  32'h3dbb90ec /* (21, 12, 28) */,
  32'h3dff07bf /* (17, 12, 28) */,
  32'h3dec6d9f /* (13, 12, 28) */,
  32'h3d902ce0 /* (9, 12, 28) */,
  32'h3d431db1 /* (5, 12, 28) */,
  32'h3d27af27 /* (1, 12, 28) */,
  32'h3d13fed6 /* (29, 8, 28) */,
  32'h3d250b86 /* (25, 8, 28) */,
  32'h3d683712 /* (21, 8, 28) */,
  32'h3d8e8b3a /* (17, 8, 28) */,
  32'h3d8a5278 /* (13, 8, 28) */,
  32'h3d3f1eea /* (9, 8, 28) */,
  32'h3d183845 /* (5, 8, 28) */,
  32'h3d139499 /* (1, 8, 28) */,
  32'h3d358b49 /* (29, 4, 28) */,
  32'h3d148979 /* (25, 4, 28) */,
  32'h3d2c64eb /* (21, 4, 28) */,
  32'h3d3f317e /* (17, 4, 28) */,
  32'h3d41aa67 /* (13, 4, 28) */,
  32'h3d19e157 /* (9, 4, 28) */,
  32'h3d1e7527 /* (5, 4, 28) */,
  32'h3d4cb45d /* (1, 4, 28) */,
  32'h3d7541a2 /* (29, 0, 28) */,
  32'h3d1879c9 /* (25, 0, 28) */,
  32'h3d1e982c /* (21, 0, 28) */,
  32'h3d27f384 /* (17, 0, 28) */,
  32'h3d2d543a /* (13, 0, 28) */,
  32'h3d13aacb /* (9, 0, 28) */,
  32'h3d3577a5 /* (5, 0, 28) */,
  32'h3da3aa58 /* (1, 0, 28) */,
  32'h3d13fed6 /* (29, 28, 24) */,
  32'h3d250b86 /* (25, 28, 24) */,
  32'h3d683712 /* (21, 28, 24) */,
  32'h3d8e8b3a /* (17, 28, 24) */,
  32'h3d8a5278 /* (13, 28, 24) */,
  32'h3d3f1eea /* (9, 28, 24) */,
  32'h3d183845 /* (5, 28, 24) */,
  32'h3d139499 /* (1, 28, 24) */,
  32'h3d2a2238 /* (29, 24, 24) */,
  32'h3d54dbd1 /* (25, 24, 24) */,
  32'h3da5dafd /* (21, 24, 24) */,
  32'h3dd9f1d0 /* (17, 24, 24) */,
  32'h3dcd36cb /* (13, 24, 24) */,
  32'h3d824402 /* (9, 24, 24) */,
  32'h3d38dbff /* (5, 24, 24) */,
  32'h3d23fb6f /* (1, 24, 24) */,
  32'h3d729483 /* (29, 20, 24) */,
  32'h3da58a7f /* (25, 20, 24) */,
  32'h3e0dbead /* (21, 20, 24) */,
  32'h3e48a298 /* (17, 20, 24) */,
  32'h3e368e5b /* (13, 20, 24) */,
  32'h3dd4c19e /* (9, 20, 24) */,
  32'h3d89129f /* (5, 20, 24) */,
  32'h3d649547 /* (1, 20, 24) */,
  32'h3d76a38f /* (29, 16, 24) */,
  32'h3db1ba44 /* (25, 16, 24) */,
  32'h3e2301df /* (21, 16, 24) */,
  32'h3e75b861 /* (17, 16, 24) */,
  32'h3e58f4b1 /* (13, 16, 24) */,
  32'h3dec5cc9 /* (9, 16, 24) */,
  32'h3d8eb3bf /* (5, 16, 24) */,
  32'h3d656b11 /* (1, 16, 24) */,
  32'h3d729483 /* (29, 12, 24) */,
  32'h3da58a7f /* (25, 12, 24) */,
  32'h3e0dbead /* (21, 12, 24) */,
  32'h3e48a298 /* (17, 12, 24) */,
  32'h3e368e5b /* (13, 12, 24) */,
  32'h3dd4c19e /* (9, 12, 24) */,
  32'h3d89129f /* (5, 12, 24) */,
  32'h3d649547 /* (1, 12, 24) */,
  32'h3d2a2238 /* (29, 8, 24) */,
  32'h3d54dbd1 /* (25, 8, 24) */,
  32'h3da5dafd /* (21, 8, 24) */,
  32'h3dd9f1d0 /* (17, 8, 24) */,
  32'h3dcd36cb /* (13, 8, 24) */,
  32'h3d824402 /* (9, 8, 24) */,
  32'h3d38dbff /* (5, 8, 24) */,
  32'h3d23fb6f /* (1, 8, 24) */,
  32'h3d13fed6 /* (29, 4, 24) */,
  32'h3d250b86 /* (25, 4, 24) */,
  32'h3d683712 /* (21, 4, 24) */,
  32'h3d8e8b3a /* (17, 4, 24) */,
  32'h3d8a5278 /* (13, 4, 24) */,
  32'h3d3f1eea /* (9, 4, 24) */,
  32'h3d183845 /* (5, 4, 24) */,
  32'h3d139499 /* (1, 4, 24) */,
  32'h3d14a194 /* (29, 0, 24) */,
  32'h3d1b34b2 /* (25, 0, 24) */,
  32'h3d4fd499 /* (21, 0, 24) */,
  32'h3d77d78b /* (17, 0, 24) */,
  32'h3d7388b1 /* (13, 0, 24) */,
  32'h3d2eceba /* (9, 0, 24) */,
  32'h3d13eed3 /* (5, 0, 24) */,
  32'h3d177e6a /* (1, 0, 24) */,
  32'h3d30047a /* (29, 28, 20) */,
  32'h3d66108f /* (25, 28, 20) */,
  32'h3dbb90ec /* (21, 28, 20) */,
  32'h3dff07bf /* (17, 28, 20) */,
  32'h3dec6d9f /* (13, 28, 20) */,
  32'h3d902ce0 /* (9, 28, 20) */,
  32'h3d431db1 /* (5, 28, 20) */,
  32'h3d27af27 /* (1, 28, 20) */,
  32'h3d729483 /* (29, 24, 20) */,
  32'h3da58a7f /* (25, 24, 20) */,
  32'h3e0dbead /* (21, 24, 20) */,
  32'h3e48a298 /* (17, 24, 20) */,
  32'h3e368e5b /* (13, 24, 20) */,
  32'h3dd4c19e /* (9, 24, 20) */,
  32'h3d89129f /* (5, 24, 20) */,
  32'h3d649547 /* (1, 24, 20) */,
  32'h3dc823b1 /* (29, 20, 20) */,
  32'h3e0e8e1e /* (25, 20, 20) */,
  32'h3e80c082 /* (21, 20, 20) */,
  32'h3ebf3a63 /* (17, 20, 20) */,
  32'h3eaa0eb2 /* (13, 20, 20) */,
  32'h3e3c290c /* (9, 20, 20) */,
  32'h3de671da /* (5, 20, 20) */,
  32'h3dbaaaa9 /* (1, 20, 20) */,
  32'h3de007f6 /* (29, 16, 20) */,
  32'h3e24eefd /* (25, 16, 20) */,
  32'h3e9bce24 /* (21, 16, 20) */,
  32'h3ef1f40b /* (17, 16, 20) */,
  32'h3ed28b29 /* (13, 16, 20) */,
  32'h3e5e82df /* (9, 16, 20) */,
  32'h3e02cee2 /* (5, 16, 20) */,
  32'h3dcf60c6 /* (1, 16, 20) */,
  32'h3dc823b1 /* (29, 12, 20) */,
  32'h3e0e8e1e /* (25, 12, 20) */,
  32'h3e80c082 /* (21, 12, 20) */,
  32'h3ebf3a63 /* (17, 12, 20) */,
  32'h3eaa0eb2 /* (13, 12, 20) */,
  32'h3e3c290c /* (9, 12, 20) */,
  32'h3de671da /* (5, 12, 20) */,
  32'h3dbaaaa9 /* (1, 12, 20) */,
  32'h3d729483 /* (29, 8, 20) */,
  32'h3da58a7f /* (25, 8, 20) */,
  32'h3e0dbead /* (21, 8, 20) */,
  32'h3e48a298 /* (17, 8, 20) */,
  32'h3e368e5b /* (13, 8, 20) */,
  32'h3dd4c19e /* (9, 8, 20) */,
  32'h3d89129f /* (5, 8, 20) */,
  32'h3d649547 /* (1, 8, 20) */,
  32'h3d30047a /* (29, 4, 20) */,
  32'h3d66108f /* (25, 4, 20) */,
  32'h3dbb90ec /* (21, 4, 20) */,
  32'h3dff07bf /* (17, 4, 20) */,
  32'h3dec6d9f /* (13, 4, 20) */,
  32'h3d902ce0 /* (9, 4, 20) */,
  32'h3d431db1 /* (5, 4, 20) */,
  32'h3d27af27 /* (1, 4, 20) */,
  32'h3d202826 /* (29, 0, 20) */,
  32'h3d4d39f8 /* (25, 0, 20) */,
  32'h3da3d600 /* (21, 0, 20) */,
  32'h3ddb309a /* (17, 0, 20) */,
  32'h3dccb681 /* (13, 0, 20) */,
  32'h3d7e6b4b /* (9, 0, 20) */,
  32'h3d2ff16f /* (5, 0, 20) */,
  32'h3d195f14 /* (1, 0, 20) */,
  32'h3d232f37 /* (29, 28, 16) */,
  32'h3d66e7bc /* (25, 28, 16) */,
  32'h3dcebbc1 /* (21, 28, 16) */,
  32'h3e18449a /* (17, 28, 16) */,
  32'h3e07f264 /* (13, 28, 16) */,
  32'h3d97bb42 /* (9, 28, 16) */,
  32'h3d3b5943 /* (5, 28, 16) */,
  32'h3d18708b /* (1, 28, 16) */,
  32'h3d76a38f /* (29, 24, 16) */,
  32'h3db1ba44 /* (25, 24, 16) */,
  32'h3e2301df /* (21, 24, 16) */,
  32'h3e75b861 /* (17, 24, 16) */,
  32'h3e58f4b1 /* (13, 24, 16) */,
  32'h3dec5cc9 /* (9, 24, 16) */,
  32'h3d8eb3bf /* (5, 24, 16) */,
  32'h3d656b11 /* (1, 24, 16) */,
  32'h3de007f6 /* (29, 20, 16) */,
  32'h3e24eefd /* (25, 20, 16) */,
  32'h3e9bce24 /* (21, 20, 16) */,
  32'h3ef1f40b /* (17, 20, 16) */,
  32'h3ed28b29 /* (13, 20, 16) */,
  32'h3e5e82df /* (9, 20, 16) */,
  32'h3e02cee2 /* (5, 20, 16) */,
  32'h3dcf60c6 /* (1, 20, 16) */,
  32'h3e078d5a /* (29, 16, 16) */,
  32'h3e4b7c7a /* (25, 16, 16) */,
  32'h3ec5ad99 /* (21, 16, 16) */,
  32'h3f1e253a /* (17, 16, 16) */,
  32'h3f079668 /* (13, 16, 16) */,
  32'h3e8b1bdf /* (9, 16, 16) */,
  32'h3e1f95bf /* (5, 16, 16) */,
  32'h3df9e164 /* (1, 16, 16) */,
  32'h3de007f6 /* (29, 12, 16) */,
  32'h3e24eefd /* (25, 12, 16) */,
  32'h3e9bce24 /* (21, 12, 16) */,
  32'h3ef1f40b /* (17, 12, 16) */,
  32'h3ed28b29 /* (13, 12, 16) */,
  32'h3e5e82df /* (9, 12, 16) */,
  32'h3e02cee2 /* (5, 12, 16) */,
  32'h3dcf60c6 /* (1, 12, 16) */,
  32'h3d76a38f /* (29, 8, 16) */,
  32'h3db1ba44 /* (25, 8, 16) */,
  32'h3e2301df /* (21, 8, 16) */,
  32'h3e75b861 /* (17, 8, 16) */,
  32'h3e58f4b1 /* (13, 8, 16) */,
  32'h3dec5cc9 /* (9, 8, 16) */,
  32'h3d8eb3bf /* (5, 8, 16) */,
  32'h3d656b11 /* (1, 8, 16) */,
  32'h3d232f37 /* (29, 4, 16) */,
  32'h3d66e7bc /* (25, 4, 16) */,
  32'h3dcebbc1 /* (21, 4, 16) */,
  32'h3e18449a /* (17, 4, 16) */,
  32'h3e07f264 /* (13, 4, 16) */,
  32'h3d97bb42 /* (9, 4, 16) */,
  32'h3d3b5943 /* (5, 4, 16) */,
  32'h3d18708b /* (1, 4, 16) */,
  32'h3d0e89f8 /* (29, 0, 16) */,
  32'h3d482f92 /* (25, 0, 16) */,
  32'h3db1860e /* (21, 0, 16) */,
  32'h3e019a4f /* (17, 0, 16) */,
  32'h3de8675d /* (13, 0, 16) */,
  32'h3d82ec35 /* (9, 0, 16) */,
  32'h3d231d8f /* (5, 0, 16) */,
  32'h3d0563b9 /* (1, 0, 16) */,
  32'h3d30047a /* (29, 28, 12) */,
  32'h3d66108f /* (25, 28, 12) */,
  32'h3dbb90ec /* (21, 28, 12) */,
  32'h3dff07bf /* (17, 28, 12) */,
  32'h3dec6d9f /* (13, 28, 12) */,
  32'h3d902ce0 /* (9, 28, 12) */,
  32'h3d431db1 /* (5, 28, 12) */,
  32'h3d27af27 /* (1, 28, 12) */,
  32'h3d729483 /* (29, 24, 12) */,
  32'h3da58a7f /* (25, 24, 12) */,
  32'h3e0dbead /* (21, 24, 12) */,
  32'h3e48a298 /* (17, 24, 12) */,
  32'h3e368e5b /* (13, 24, 12) */,
  32'h3dd4c19e /* (9, 24, 12) */,
  32'h3d89129f /* (5, 24, 12) */,
  32'h3d649547 /* (1, 24, 12) */,
  32'h3dc823b1 /* (29, 20, 12) */,
  32'h3e0e8e1e /* (25, 20, 12) */,
  32'h3e80c082 /* (21, 20, 12) */,
  32'h3ebf3a63 /* (17, 20, 12) */,
  32'h3eaa0eb2 /* (13, 20, 12) */,
  32'h3e3c290c /* (9, 20, 12) */,
  32'h3de671da /* (5, 20, 12) */,
  32'h3dbaaaa9 /* (1, 20, 12) */,
  32'h3de007f6 /* (29, 16, 12) */,
  32'h3e24eefd /* (25, 16, 12) */,
  32'h3e9bce24 /* (21, 16, 12) */,
  32'h3ef1f40b /* (17, 16, 12) */,
  32'h3ed28b29 /* (13, 16, 12) */,
  32'h3e5e82df /* (9, 16, 12) */,
  32'h3e02cee2 /* (5, 16, 12) */,
  32'h3dcf60c6 /* (1, 16, 12) */,
  32'h3dc823b1 /* (29, 12, 12) */,
  32'h3e0e8e1e /* (25, 12, 12) */,
  32'h3e80c082 /* (21, 12, 12) */,
  32'h3ebf3a63 /* (17, 12, 12) */,
  32'h3eaa0eb2 /* (13, 12, 12) */,
  32'h3e3c290c /* (9, 12, 12) */,
  32'h3de671da /* (5, 12, 12) */,
  32'h3dbaaaa9 /* (1, 12, 12) */,
  32'h3d729483 /* (29, 8, 12) */,
  32'h3da58a7f /* (25, 8, 12) */,
  32'h3e0dbead /* (21, 8, 12) */,
  32'h3e48a298 /* (17, 8, 12) */,
  32'h3e368e5b /* (13, 8, 12) */,
  32'h3dd4c19e /* (9, 8, 12) */,
  32'h3d89129f /* (5, 8, 12) */,
  32'h3d649547 /* (1, 8, 12) */,
  32'h3d30047a /* (29, 4, 12) */,
  32'h3d66108f /* (25, 4, 12) */,
  32'h3dbb90ec /* (21, 4, 12) */,
  32'h3dff07bf /* (17, 4, 12) */,
  32'h3dec6d9f /* (13, 4, 12) */,
  32'h3d902ce0 /* (9, 4, 12) */,
  32'h3d431db1 /* (5, 4, 12) */,
  32'h3d27af27 /* (1, 4, 12) */,
  32'h3d202826 /* (29, 0, 12) */,
  32'h3d4d39f8 /* (25, 0, 12) */,
  32'h3da3d600 /* (21, 0, 12) */,
  32'h3ddb309a /* (17, 0, 12) */,
  32'h3dccb681 /* (13, 0, 12) */,
  32'h3d7e6b4b /* (9, 0, 12) */,
  32'h3d2ff16f /* (5, 0, 12) */,
  32'h3d195f14 /* (1, 0, 12) */,
  32'h3d13fed6 /* (29, 28, 8) */,
  32'h3d250b86 /* (25, 28, 8) */,
  32'h3d683712 /* (21, 28, 8) */,
  32'h3d8e8b3a /* (17, 28, 8) */,
  32'h3d8a5278 /* (13, 28, 8) */,
  32'h3d3f1eea /* (9, 28, 8) */,
  32'h3d183845 /* (5, 28, 8) */,
  32'h3d139499 /* (1, 28, 8) */,
  32'h3d2a2238 /* (29, 24, 8) */,
  32'h3d54dbd1 /* (25, 24, 8) */,
  32'h3da5dafd /* (21, 24, 8) */,
  32'h3dd9f1d0 /* (17, 24, 8) */,
  32'h3dcd36cb /* (13, 24, 8) */,
  32'h3d824402 /* (9, 24, 8) */,
  32'h3d38dbff /* (5, 24, 8) */,
  32'h3d23fb6f /* (1, 24, 8) */,
  32'h3d729483 /* (29, 20, 8) */,
  32'h3da58a7f /* (25, 20, 8) */,
  32'h3e0dbead /* (21, 20, 8) */,
  32'h3e48a298 /* (17, 20, 8) */,
  32'h3e368e5b /* (13, 20, 8) */,
  32'h3dd4c19e /* (9, 20, 8) */,
  32'h3d89129f /* (5, 20, 8) */,
  32'h3d649547 /* (1, 20, 8) */,
  32'h3d76a38f /* (29, 16, 8) */,
  32'h3db1ba44 /* (25, 16, 8) */,
  32'h3e2301df /* (21, 16, 8) */,
  32'h3e75b861 /* (17, 16, 8) */,
  32'h3e58f4b1 /* (13, 16, 8) */,
  32'h3dec5cc9 /* (9, 16, 8) */,
  32'h3d8eb3bf /* (5, 16, 8) */,
  32'h3d656b11 /* (1, 16, 8) */,
  32'h3d729483 /* (29, 12, 8) */,
  32'h3da58a7f /* (25, 12, 8) */,
  32'h3e0dbead /* (21, 12, 8) */,
  32'h3e48a298 /* (17, 12, 8) */,
  32'h3e368e5b /* (13, 12, 8) */,
  32'h3dd4c19e /* (9, 12, 8) */,
  32'h3d89129f /* (5, 12, 8) */,
  32'h3d649547 /* (1, 12, 8) */,
  32'h3d2a2238 /* (29, 8, 8) */,
  32'h3d54dbd1 /* (25, 8, 8) */,
  32'h3da5dafd /* (21, 8, 8) */,
  32'h3dd9f1d0 /* (17, 8, 8) */,
  32'h3dcd36cb /* (13, 8, 8) */,
  32'h3d824402 /* (9, 8, 8) */,
  32'h3d38dbff /* (5, 8, 8) */,
  32'h3d23fb6f /* (1, 8, 8) */,
  32'h3d13fed6 /* (29, 4, 8) */,
  32'h3d250b86 /* (25, 4, 8) */,
  32'h3d683712 /* (21, 4, 8) */,
  32'h3d8e8b3a /* (17, 4, 8) */,
  32'h3d8a5278 /* (13, 4, 8) */,
  32'h3d3f1eea /* (9, 4, 8) */,
  32'h3d183845 /* (5, 4, 8) */,
  32'h3d139499 /* (1, 4, 8) */,
  32'h3d14a194 /* (29, 0, 8) */,
  32'h3d1b34b2 /* (25, 0, 8) */,
  32'h3d4fd499 /* (21, 0, 8) */,
  32'h3d77d78b /* (17, 0, 8) */,
  32'h3d7388b1 /* (13, 0, 8) */,
  32'h3d2eceba /* (9, 0, 8) */,
  32'h3d13eed3 /* (5, 0, 8) */,
  32'h3d177e6a /* (1, 0, 8) */,
  32'h3d358b49 /* (29, 28, 4) */,
  32'h3d148979 /* (25, 28, 4) */,
  32'h3d2c64eb /* (21, 28, 4) */,
  32'h3d3f317e /* (17, 28, 4) */,
  32'h3d41aa67 /* (13, 28, 4) */,
  32'h3d19e157 /* (9, 28, 4) */,
  32'h3d1e7527 /* (5, 28, 4) */,
  32'h3d4cb45d /* (1, 28, 4) */,
  32'h3d13fed6 /* (29, 24, 4) */,
  32'h3d250b86 /* (25, 24, 4) */,
  32'h3d683712 /* (21, 24, 4) */,
  32'h3d8e8b3a /* (17, 24, 4) */,
  32'h3d8a5278 /* (13, 24, 4) */,
  32'h3d3f1eea /* (9, 24, 4) */,
  32'h3d183845 /* (5, 24, 4) */,
  32'h3d139499 /* (1, 24, 4) */,
  32'h3d30047a /* (29, 20, 4) */,
  32'h3d66108f /* (25, 20, 4) */,
  32'h3dbb90ec /* (21, 20, 4) */,
  32'h3dff07bf /* (17, 20, 4) */,
  32'h3dec6d9f /* (13, 20, 4) */,
  32'h3d902ce0 /* (9, 20, 4) */,
  32'h3d431db1 /* (5, 20, 4) */,
  32'h3d27af27 /* (1, 20, 4) */,
  32'h3d232f37 /* (29, 16, 4) */,
  32'h3d66e7bc /* (25, 16, 4) */,
  32'h3dcebbc1 /* (21, 16, 4) */,
  32'h3e18449a /* (17, 16, 4) */,
  32'h3e07f264 /* (13, 16, 4) */,
  32'h3d97bb42 /* (9, 16, 4) */,
  32'h3d3b5943 /* (5, 16, 4) */,
  32'h3d18708b /* (1, 16, 4) */,
  32'h3d30047a /* (29, 12, 4) */,
  32'h3d66108f /* (25, 12, 4) */,
  32'h3dbb90ec /* (21, 12, 4) */,
  32'h3dff07bf /* (17, 12, 4) */,
  32'h3dec6d9f /* (13, 12, 4) */,
  32'h3d902ce0 /* (9, 12, 4) */,
  32'h3d431db1 /* (5, 12, 4) */,
  32'h3d27af27 /* (1, 12, 4) */,
  32'h3d13fed6 /* (29, 8, 4) */,
  32'h3d250b86 /* (25, 8, 4) */,
  32'h3d683712 /* (21, 8, 4) */,
  32'h3d8e8b3a /* (17, 8, 4) */,
  32'h3d8a5278 /* (13, 8, 4) */,
  32'h3d3f1eea /* (9, 8, 4) */,
  32'h3d183845 /* (5, 8, 4) */,
  32'h3d139499 /* (1, 8, 4) */,
  32'h3d358b49 /* (29, 4, 4) */,
  32'h3d148979 /* (25, 4, 4) */,
  32'h3d2c64eb /* (21, 4, 4) */,
  32'h3d3f317e /* (17, 4, 4) */,
  32'h3d41aa67 /* (13, 4, 4) */,
  32'h3d19e157 /* (9, 4, 4) */,
  32'h3d1e7527 /* (5, 4, 4) */,
  32'h3d4cb45d /* (1, 4, 4) */,
  32'h3d7541a2 /* (29, 0, 4) */,
  32'h3d1879c9 /* (25, 0, 4) */,
  32'h3d1e982c /* (21, 0, 4) */,
  32'h3d27f384 /* (17, 0, 4) */,
  32'h3d2d543a /* (13, 0, 4) */,
  32'h3d13aacb /* (9, 0, 4) */,
  32'h3d3577a5 /* (5, 0, 4) */,
  32'h3da3aa58 /* (1, 0, 4) */,
  32'h3d7541a2 /* (29, 28, 0) */,
  32'h3d1879c9 /* (25, 28, 0) */,
  32'h3d1e982c /* (21, 28, 0) */,
  32'h3d27f384 /* (17, 28, 0) */,
  32'h3d2d543a /* (13, 28, 0) */,
  32'h3d13aacb /* (9, 28, 0) */,
  32'h3d3577a5 /* (5, 28, 0) */,
  32'h3da3aa58 /* (1, 28, 0) */,
  32'h3d14a194 /* (29, 24, 0) */,
  32'h3d1b34b2 /* (25, 24, 0) */,
  32'h3d4fd499 /* (21, 24, 0) */,
  32'h3d77d78b /* (17, 24, 0) */,
  32'h3d7388b1 /* (13, 24, 0) */,
  32'h3d2eceba /* (9, 24, 0) */,
  32'h3d13eed3 /* (5, 24, 0) */,
  32'h3d177e6a /* (1, 24, 0) */,
  32'h3d202826 /* (29, 20, 0) */,
  32'h3d4d39f8 /* (25, 20, 0) */,
  32'h3da3d600 /* (21, 20, 0) */,
  32'h3ddb309a /* (17, 20, 0) */,
  32'h3dccb681 /* (13, 20, 0) */,
  32'h3d7e6b4b /* (9, 20, 0) */,
  32'h3d2ff16f /* (5, 20, 0) */,
  32'h3d195f14 /* (1, 20, 0) */,
  32'h3d0e89f8 /* (29, 16, 0) */,
  32'h3d482f92 /* (25, 16, 0) */,
  32'h3db1860e /* (21, 16, 0) */,
  32'h3e019a4f /* (17, 16, 0) */,
  32'h3de8675d /* (13, 16, 0) */,
  32'h3d82ec35 /* (9, 16, 0) */,
  32'h3d231d8f /* (5, 16, 0) */,
  32'h3d0563b9 /* (1, 16, 0) */,
  32'h3d202826 /* (29, 12, 0) */,
  32'h3d4d39f8 /* (25, 12, 0) */,
  32'h3da3d600 /* (21, 12, 0) */,
  32'h3ddb309a /* (17, 12, 0) */,
  32'h3dccb681 /* (13, 12, 0) */,
  32'h3d7e6b4b /* (9, 12, 0) */,
  32'h3d2ff16f /* (5, 12, 0) */,
  32'h3d195f14 /* (1, 12, 0) */,
  32'h3d14a194 /* (29, 8, 0) */,
  32'h3d1b34b2 /* (25, 8, 0) */,
  32'h3d4fd499 /* (21, 8, 0) */,
  32'h3d77d78b /* (17, 8, 0) */,
  32'h3d7388b1 /* (13, 8, 0) */,
  32'h3d2eceba /* (9, 8, 0) */,
  32'h3d13eed3 /* (5, 8, 0) */,
  32'h3d177e6a /* (1, 8, 0) */,
  32'h3d7541a2 /* (29, 4, 0) */,
  32'h3d1879c9 /* (25, 4, 0) */,
  32'h3d1e982c /* (21, 4, 0) */,
  32'h3d27f384 /* (17, 4, 0) */,
  32'h3d2d543a /* (13, 4, 0) */,
  32'h3d13aacb /* (9, 4, 0) */,
  32'h3d3577a5 /* (5, 4, 0) */,
  32'h3da3aa58 /* (1, 4, 0) */,
  32'h3e0c4c59 /* (29, 0, 0) */,
  32'h3d269d45 /* (25, 0, 0) */,
  32'h3d13eab3 /* (21, 0, 0) */,
  32'h3d14300c /* (17, 0, 0) */,
  32'h3d1c4c09 /* (13, 0, 0) */,
  32'h3d11ab15 /* (9, 0, 0) */,
  32'h3d75271a /* (5, 0, 0) */,
  32'h3f8f3ec8 /* (1, 0, 0) */,
  32'h3d28c974 /* (28, 28, 28) */,
  32'h3d15577e /* (24, 28, 28) */,
  32'h3d37f7fd /* (20, 28, 28) */,
  32'h3d2d4da1 /* (16, 28, 28) */,
  32'h3d37f7fd /* (12, 28, 28) */,
  32'h3d15577e /* (8, 28, 28) */,
  32'h3d28c974 /* (4, 28, 28) */,
  32'h3d508e8d /* (0, 28, 28) */,
  32'h3d15577e /* (28, 24, 28) */,
  32'h3d302eb0 /* (24, 24, 28) */,
  32'h3d7fc9dc /* (20, 24, 28) */,
  32'h3d836eb0 /* (16, 24, 28) */,
  32'h3d7fc9dc /* (12, 24, 28) */,
  32'h3d302eb0 /* (8, 24, 28) */,
  32'h3d15577e /* (4, 24, 28) */,
  32'h3d139fbd /* (0, 24, 28) */,
  32'h3d37f7fd /* (28, 20, 28) */,
  32'h3d7fc9dc /* (24, 20, 28) */,
  32'h3dd4d413 /* (20, 20, 28) */,
  32'h3defbf1f /* (16, 20, 28) */,
  32'h3dd4d413 /* (12, 20, 28) */,
  32'h3d7fc9dc /* (8, 20, 28) */,
  32'h3d37f7fd /* (4, 20, 28) */,
  32'h3d26b2c0 /* (0, 20, 28) */,
  32'h3d2d4da1 /* (28, 16, 28) */,
  32'h3d836eb0 /* (24, 16, 28) */,
  32'h3defbf1f /* (20, 16, 28) */,
  32'h3e11966c /* (16, 16, 28) */,
  32'h3defbf1f /* (12, 16, 28) */,
  32'h3d836eb0 /* (8, 16, 28) */,
  32'h3d2d4da1 /* (4, 16, 28) */,
  32'h3d1727de /* (0, 16, 28) */,
  32'h3d37f7fd /* (28, 12, 28) */,
  32'h3d7fc9dc /* (24, 12, 28) */,
  32'h3dd4d413 /* (20, 12, 28) */,
  32'h3defbf1f /* (16, 12, 28) */,
  32'h3dd4d413 /* (12, 12, 28) */,
  32'h3d7fc9dc /* (8, 12, 28) */,
  32'h3d37f7fd /* (4, 12, 28) */,
  32'h3d26b2c0 /* (0, 12, 28) */,
  32'h3d15577e /* (28, 8, 28) */,
  32'h3d302eb0 /* (24, 8, 28) */,
  32'h3d7fc9dc /* (20, 8, 28) */,
  32'h3d836eb0 /* (16, 8, 28) */,
  32'h3d7fc9dc /* (12, 8, 28) */,
  32'h3d302eb0 /* (8, 8, 28) */,
  32'h3d15577e /* (4, 8, 28) */,
  32'h3d139fbd /* (0, 8, 28) */,
  32'h3d28c974 /* (28, 4, 28) */,
  32'h3d15577e /* (24, 4, 28) */,
  32'h3d37f7fd /* (20, 4, 28) */,
  32'h3d2d4da1 /* (16, 4, 28) */,
  32'h3d37f7fd /* (12, 4, 28) */,
  32'h3d15577e /* (8, 4, 28) */,
  32'h3d28c974 /* (4, 4, 28) */,
  32'h3d508e8d /* (0, 4, 28) */,
  32'h3d508e8d /* (28, 0, 28) */,
  32'h3d139fbd /* (24, 0, 28) */,
  32'h3d26b2c0 /* (20, 0, 28) */,
  32'h3d1727de /* (16, 0, 28) */,
  32'h3d26b2c0 /* (12, 0, 28) */,
  32'h3d139fbd /* (8, 0, 28) */,
  32'h3d508e8d /* (4, 0, 28) */,
  32'h3dabcc5c /* (0, 0, 28) */,
  32'h3d15577e /* (28, 28, 24) */,
  32'h3d302eb0 /* (24, 28, 24) */,
  32'h3d7fc9dc /* (20, 28, 24) */,
  32'h3d836eb0 /* (16, 28, 24) */,
  32'h3d7fc9dc /* (12, 28, 24) */,
  32'h3d302eb0 /* (8, 28, 24) */,
  32'h3d15577e /* (4, 28, 24) */,
  32'h3d139fbd /* (0, 28, 24) */,
  32'h3d302eb0 /* (28, 24, 24) */,
  32'h3d69d3eb /* (24, 24, 24) */,
  32'h3dba61a5 /* (20, 24, 24) */,
  32'h3dcb8235 /* (16, 24, 24) */,
  32'h3dba61a5 /* (12, 24, 24) */,
  32'h3d69d3eb /* (8, 24, 24) */,
  32'h3d302eb0 /* (4, 24, 24) */,
  32'h3d234568 /* (0, 24, 24) */,
  32'h3d7fc9dc /* (28, 20, 24) */,
  32'h3dba61a5 /* (24, 20, 24) */,
  32'h3e22a180 /* (20, 20, 24) */,
  32'h3e3e2eae /* (16, 20, 24) */,
  32'h3e22a180 /* (12, 20, 24) */,
  32'h3dba61a5 /* (8, 20, 24) */,
  32'h3d7fc9dc /* (4, 20, 24) */,
  32'h3d62e9d3 /* (0, 20, 24) */,
  32'h3d836eb0 /* (28, 16, 24) */,
  32'h3dcb8235 /* (24, 16, 24) */,
  32'h3e3e2eae /* (20, 16, 24) */,
  32'h3e6c2939 /* (16, 16, 24) */,
  32'h3e3e2eae /* (12, 16, 24) */,
  32'h3dcb8235 /* (8, 16, 24) */,
  32'h3d836eb0 /* (4, 16, 24) */,
  32'h3d635c6b /* (0, 16, 24) */,
  32'h3d7fc9dc /* (28, 12, 24) */,
  32'h3dba61a5 /* (24, 12, 24) */,
  32'h3e22a180 /* (20, 12, 24) */,
  32'h3e3e2eae /* (16, 12, 24) */,
  32'h3e22a180 /* (12, 12, 24) */,
  32'h3dba61a5 /* (8, 12, 24) */,
  32'h3d7fc9dc /* (4, 12, 24) */,
  32'h3d62e9d3 /* (0, 12, 24) */,
  32'h3d302eb0 /* (28, 8, 24) */,
  32'h3d69d3eb /* (24, 8, 24) */,
  32'h3dba61a5 /* (20, 8, 24) */,
  32'h3dcb8235 /* (16, 8, 24) */,
  32'h3dba61a5 /* (12, 8, 24) */,
  32'h3d69d3eb /* (8, 8, 24) */,
  32'h3d302eb0 /* (4, 8, 24) */,
  32'h3d234568 /* (0, 8, 24) */,
  32'h3d15577e /* (28, 4, 24) */,
  32'h3d302eb0 /* (24, 4, 24) */,
  32'h3d7fc9dc /* (20, 4, 24) */,
  32'h3d836eb0 /* (16, 4, 24) */,
  32'h3d7fc9dc /* (12, 4, 24) */,
  32'h3d302eb0 /* (8, 4, 24) */,
  32'h3d15577e /* (4, 4, 24) */,
  32'h3d139fbd /* (0, 4, 24) */,
  32'h3d139fbd /* (28, 0, 24) */,
  32'h3d234568 /* (24, 0, 24) */,
  32'h3d62e9d3 /* (20, 0, 24) */,
  32'h3d635c6b /* (16, 0, 24) */,
  32'h3d62e9d3 /* (12, 0, 24) */,
  32'h3d234568 /* (8, 0, 24) */,
  32'h3d139fbd /* (4, 0, 24) */,
  32'h3d180196 /* (0, 0, 24) */,
  32'h3d37f7fd /* (28, 28, 20) */,
  32'h3d7fc9dc /* (24, 28, 20) */,
  32'h3dd4d413 /* (20, 28, 20) */,
  32'h3defbf1f /* (16, 28, 20) */,
  32'h3dd4d413 /* (12, 28, 20) */,
  32'h3d7fc9dc /* (8, 28, 20) */,
  32'h3d37f7fd /* (4, 28, 20) */,
  32'h3d26b2c0 /* (0, 28, 20) */,
  32'h3d7fc9dc /* (28, 24, 20) */,
  32'h3dba61a5 /* (24, 24, 20) */,
  32'h3e22a180 /* (20, 24, 20) */,
  32'h3e3e2eae /* (16, 24, 20) */,
  32'h3e22a180 /* (12, 24, 20) */,
  32'h3dba61a5 /* (8, 24, 20) */,
  32'h3d7fc9dc /* (4, 24, 20) */,
  32'h3d62e9d3 /* (0, 24, 20) */,
  32'h3dd4d413 /* (28, 20, 20) */,
  32'h3e22a180 /* (24, 20, 20) */,
  32'h3e95a2cf /* (20, 20, 20) */,
  32'h3eb72c7f /* (16, 20, 20) */,
  32'h3e95a2cf /* (12, 20, 20) */,
  32'h3e22a180 /* (8, 20, 20) */,
  32'h3dd4d413 /* (4, 20, 20) */,
  32'h3db90e8b /* (0, 20, 20) */,
  32'h3defbf1f /* (28, 16, 20) */,
  32'h3e3e2eae /* (24, 16, 20) */,
  32'h3eb72c7f /* (20, 16, 20) */,
  32'h3eea2758 /* (16, 16, 20) */,
  32'h3eb72c7f /* (12, 16, 20) */,
  32'h3e3e2eae /* (8, 16, 20) */,
  32'h3defbf1f /* (4, 16, 20) */,
  32'h3dcd63f0 /* (0, 16, 20) */,
  32'h3dd4d413 /* (28, 12, 20) */,
  32'h3e22a180 /* (24, 12, 20) */,
  32'h3e95a2cf /* (20, 12, 20) */,
  32'h3eb72c7f /* (16, 12, 20) */,
  32'h3e95a2cf /* (12, 12, 20) */,
  32'h3e22a180 /* (8, 12, 20) */,
  32'h3dd4d413 /* (4, 12, 20) */,
  32'h3db90e8b /* (0, 12, 20) */,
  32'h3d7fc9dc /* (28, 8, 20) */,
  32'h3dba61a5 /* (24, 8, 20) */,
  32'h3e22a180 /* (20, 8, 20) */,
  32'h3e3e2eae /* (16, 8, 20) */,
  32'h3e22a180 /* (12, 8, 20) */,
  32'h3dba61a5 /* (8, 8, 20) */,
  32'h3d7fc9dc /* (4, 8, 20) */,
  32'h3d62e9d3 /* (0, 8, 20) */,
  32'h3d37f7fd /* (28, 4, 20) */,
  32'h3d7fc9dc /* (24, 4, 20) */,
  32'h3dd4d413 /* (20, 4, 20) */,
  32'h3defbf1f /* (16, 4, 20) */,
  32'h3dd4d413 /* (12, 4, 20) */,
  32'h3d7fc9dc /* (8, 4, 20) */,
  32'h3d37f7fd /* (4, 4, 20) */,
  32'h3d26b2c0 /* (0, 4, 20) */,
  32'h3d26b2c0 /* (28, 0, 20) */,
  32'h3d62e9d3 /* (24, 0, 20) */,
  32'h3db90e8b /* (20, 0, 20) */,
  32'h3dcd63f0 /* (16, 0, 20) */,
  32'h3db90e8b /* (12, 0, 20) */,
  32'h3d62e9d3 /* (8, 0, 20) */,
  32'h3d26b2c0 /* (4, 0, 20) */,
  32'h3d189328 /* (0, 0, 20) */,
  32'h3d2d4da1 /* (28, 28, 16) */,
  32'h3d836eb0 /* (24, 28, 16) */,
  32'h3defbf1f /* (20, 28, 16) */,
  32'h3e11966c /* (16, 28, 16) */,
  32'h3defbf1f /* (12, 28, 16) */,
  32'h3d836eb0 /* (8, 28, 16) */,
  32'h3d2d4da1 /* (4, 28, 16) */,
  32'h3d1727de /* (0, 28, 16) */,
  32'h3d836eb0 /* (28, 24, 16) */,
  32'h3dcb8235 /* (24, 24, 16) */,
  32'h3e3e2eae /* (20, 24, 16) */,
  32'h3e6c2939 /* (16, 24, 16) */,
  32'h3e3e2eae /* (12, 24, 16) */,
  32'h3dcb8235 /* (8, 24, 16) */,
  32'h3d836eb0 /* (4, 24, 16) */,
  32'h3d635c6b /* (0, 24, 16) */,
  32'h3defbf1f /* (28, 20, 16) */,
  32'h3e3e2eae /* (24, 20, 16) */,
  32'h3eb72c7f /* (20, 20, 16) */,
  32'h3eea2758 /* (16, 20, 16) */,
  32'h3eb72c7f /* (12, 20, 16) */,
  32'h3e3e2eae /* (8, 20, 16) */,
  32'h3defbf1f /* (4, 20, 16) */,
  32'h3dcd63f0 /* (0, 20, 16) */,
  32'h3e11966c /* (28, 16, 16) */,
  32'h3e6c2939 /* (24, 16, 16) */,
  32'h3eea2758 /* (20, 16, 16) */,
  32'h3f1a278c /* (16, 16, 16) */,
  32'h3eea2758 /* (12, 16, 16) */,
  32'h3e6c2939 /* (8, 16, 16) */,
  32'h3e11966c /* (4, 16, 16) */,
  32'h3df759b6 /* (0, 16, 16) */,
  32'h3defbf1f /* (28, 12, 16) */,
  32'h3e3e2eae /* (24, 12, 16) */,
  32'h3eb72c7f /* (20, 12, 16) */,
  32'h3eea2758 /* (16, 12, 16) */,
  32'h3eb72c7f /* (12, 12, 16) */,
  32'h3e3e2eae /* (8, 12, 16) */,
  32'h3defbf1f /* (4, 12, 16) */,
  32'h3dcd63f0 /* (0, 12, 16) */,
  32'h3d836eb0 /* (28, 8, 16) */,
  32'h3dcb8235 /* (24, 8, 16) */,
  32'h3e3e2eae /* (20, 8, 16) */,
  32'h3e6c2939 /* (16, 8, 16) */,
  32'h3e3e2eae /* (12, 8, 16) */,
  32'h3dcb8235 /* (8, 8, 16) */,
  32'h3d836eb0 /* (4, 8, 16) */,
  32'h3d635c6b /* (0, 8, 16) */,
  32'h3d2d4da1 /* (28, 4, 16) */,
  32'h3d836eb0 /* (24, 4, 16) */,
  32'h3defbf1f /* (20, 4, 16) */,
  32'h3e11966c /* (16, 4, 16) */,
  32'h3defbf1f /* (12, 4, 16) */,
  32'h3d836eb0 /* (8, 4, 16) */,
  32'h3d2d4da1 /* (4, 4, 16) */,
  32'h3d1727de /* (0, 4, 16) */,
  32'h3d1727de /* (28, 0, 16) */,
  32'h3d635c6b /* (24, 0, 16) */,
  32'h3dcd63f0 /* (20, 0, 16) */,
  32'h3df759b6 /* (16, 0, 16) */,
  32'h3dcd63f0 /* (12, 0, 16) */,
  32'h3d635c6b /* (8, 0, 16) */,
  32'h3d1727de /* (4, 0, 16) */,
  32'h3d044bdf /* (0, 0, 16) */,
  32'h3d37f7fd /* (28, 28, 12) */,
  32'h3d7fc9dc /* (24, 28, 12) */,
  32'h3dd4d413 /* (20, 28, 12) */,
  32'h3defbf1f /* (16, 28, 12) */,
  32'h3dd4d413 /* (12, 28, 12) */,
  32'h3d7fc9dc /* (8, 28, 12) */,
  32'h3d37f7fd /* (4, 28, 12) */,
  32'h3d26b2c0 /* (0, 28, 12) */,
  32'h3d7fc9dc /* (28, 24, 12) */,
  32'h3dba61a5 /* (24, 24, 12) */,
  32'h3e22a180 /* (20, 24, 12) */,
  32'h3e3e2eae /* (16, 24, 12) */,
  32'h3e22a180 /* (12, 24, 12) */,
  32'h3dba61a5 /* (8, 24, 12) */,
  32'h3d7fc9dc /* (4, 24, 12) */,
  32'h3d62e9d3 /* (0, 24, 12) */,
  32'h3dd4d413 /* (28, 20, 12) */,
  32'h3e22a180 /* (24, 20, 12) */,
  32'h3e95a2cf /* (20, 20, 12) */,
  32'h3eb72c7f /* (16, 20, 12) */,
  32'h3e95a2cf /* (12, 20, 12) */,
  32'h3e22a180 /* (8, 20, 12) */,
  32'h3dd4d413 /* (4, 20, 12) */,
  32'h3db90e8b /* (0, 20, 12) */,
  32'h3defbf1f /* (28, 16, 12) */,
  32'h3e3e2eae /* (24, 16, 12) */,
  32'h3eb72c7f /* (20, 16, 12) */,
  32'h3eea2758 /* (16, 16, 12) */,
  32'h3eb72c7f /* (12, 16, 12) */,
  32'h3e3e2eae /* (8, 16, 12) */,
  32'h3defbf1f /* (4, 16, 12) */,
  32'h3dcd63f0 /* (0, 16, 12) */,
  32'h3dd4d413 /* (28, 12, 12) */,
  32'h3e22a180 /* (24, 12, 12) */,
  32'h3e95a2cf /* (20, 12, 12) */,
  32'h3eb72c7f /* (16, 12, 12) */,
  32'h3e95a2cf /* (12, 12, 12) */,
  32'h3e22a180 /* (8, 12, 12) */,
  32'h3dd4d413 /* (4, 12, 12) */,
  32'h3db90e8b /* (0, 12, 12) */,
  32'h3d7fc9dc /* (28, 8, 12) */,
  32'h3dba61a5 /* (24, 8, 12) */,
  32'h3e22a180 /* (20, 8, 12) */,
  32'h3e3e2eae /* (16, 8, 12) */,
  32'h3e22a180 /* (12, 8, 12) */,
  32'h3dba61a5 /* (8, 8, 12) */,
  32'h3d7fc9dc /* (4, 8, 12) */,
  32'h3d62e9d3 /* (0, 8, 12) */,
  32'h3d37f7fd /* (28, 4, 12) */,
  32'h3d7fc9dc /* (24, 4, 12) */,
  32'h3dd4d413 /* (20, 4, 12) */,
  32'h3defbf1f /* (16, 4, 12) */,
  32'h3dd4d413 /* (12, 4, 12) */,
  32'h3d7fc9dc /* (8, 4, 12) */,
  32'h3d37f7fd /* (4, 4, 12) */,
  32'h3d26b2c0 /* (0, 4, 12) */,
  32'h3d26b2c0 /* (28, 0, 12) */,
  32'h3d62e9d3 /* (24, 0, 12) */,
  32'h3db90e8b /* (20, 0, 12) */,
  32'h3dcd63f0 /* (16, 0, 12) */,
  32'h3db90e8b /* (12, 0, 12) */,
  32'h3d62e9d3 /* (8, 0, 12) */,
  32'h3d26b2c0 /* (4, 0, 12) */,
  32'h3d189328 /* (0, 0, 12) */,
  32'h3d15577e /* (28, 28, 8) */,
  32'h3d302eb0 /* (24, 28, 8) */,
  32'h3d7fc9dc /* (20, 28, 8) */,
  32'h3d836eb0 /* (16, 28, 8) */,
  32'h3d7fc9dc /* (12, 28, 8) */,
  32'h3d302eb0 /* (8, 28, 8) */,
  32'h3d15577e /* (4, 28, 8) */,
  32'h3d139fbd /* (0, 28, 8) */,
  32'h3d302eb0 /* (28, 24, 8) */,
  32'h3d69d3eb /* (24, 24, 8) */,
  32'h3dba61a5 /* (20, 24, 8) */,
  32'h3dcb8235 /* (16, 24, 8) */,
  32'h3dba61a5 /* (12, 24, 8) */,
  32'h3d69d3eb /* (8, 24, 8) */,
  32'h3d302eb0 /* (4, 24, 8) */,
  32'h3d234568 /* (0, 24, 8) */,
  32'h3d7fc9dc /* (28, 20, 8) */,
  32'h3dba61a5 /* (24, 20, 8) */,
  32'h3e22a180 /* (20, 20, 8) */,
  32'h3e3e2eae /* (16, 20, 8) */,
  32'h3e22a180 /* (12, 20, 8) */,
  32'h3dba61a5 /* (8, 20, 8) */,
  32'h3d7fc9dc /* (4, 20, 8) */,
  32'h3d62e9d3 /* (0, 20, 8) */,
  32'h3d836eb0 /* (28, 16, 8) */,
  32'h3dcb8235 /* (24, 16, 8) */,
  32'h3e3e2eae /* (20, 16, 8) */,
  32'h3e6c2939 /* (16, 16, 8) */,
  32'h3e3e2eae /* (12, 16, 8) */,
  32'h3dcb8235 /* (8, 16, 8) */,
  32'h3d836eb0 /* (4, 16, 8) */,
  32'h3d635c6b /* (0, 16, 8) */,
  32'h3d7fc9dc /* (28, 12, 8) */,
  32'h3dba61a5 /* (24, 12, 8) */,
  32'h3e22a180 /* (20, 12, 8) */,
  32'h3e3e2eae /* (16, 12, 8) */,
  32'h3e22a180 /* (12, 12, 8) */,
  32'h3dba61a5 /* (8, 12, 8) */,
  32'h3d7fc9dc /* (4, 12, 8) */,
  32'h3d62e9d3 /* (0, 12, 8) */,
  32'h3d302eb0 /* (28, 8, 8) */,
  32'h3d69d3eb /* (24, 8, 8) */,
  32'h3dba61a5 /* (20, 8, 8) */,
  32'h3dcb8235 /* (16, 8, 8) */,
  32'h3dba61a5 /* (12, 8, 8) */,
  32'h3d69d3eb /* (8, 8, 8) */,
  32'h3d302eb0 /* (4, 8, 8) */,
  32'h3d234568 /* (0, 8, 8) */,
  32'h3d15577e /* (28, 4, 8) */,
  32'h3d302eb0 /* (24, 4, 8) */,
  32'h3d7fc9dc /* (20, 4, 8) */,
  32'h3d836eb0 /* (16, 4, 8) */,
  32'h3d7fc9dc /* (12, 4, 8) */,
  32'h3d302eb0 /* (8, 4, 8) */,
  32'h3d15577e /* (4, 4, 8) */,
  32'h3d139fbd /* (0, 4, 8) */,
  32'h3d139fbd /* (28, 0, 8) */,
  32'h3d234568 /* (24, 0, 8) */,
  32'h3d62e9d3 /* (20, 0, 8) */,
  32'h3d635c6b /* (16, 0, 8) */,
  32'h3d62e9d3 /* (12, 0, 8) */,
  32'h3d234568 /* (8, 0, 8) */,
  32'h3d139fbd /* (4, 0, 8) */,
  32'h3d180196 /* (0, 0, 8) */,
  32'h3d28c974 /* (28, 28, 4) */,
  32'h3d15577e /* (24, 28, 4) */,
  32'h3d37f7fd /* (20, 28, 4) */,
  32'h3d2d4da1 /* (16, 28, 4) */,
  32'h3d37f7fd /* (12, 28, 4) */,
  32'h3d15577e /* (8, 28, 4) */,
  32'h3d28c974 /* (4, 28, 4) */,
  32'h3d508e8d /* (0, 28, 4) */,
  32'h3d15577e /* (28, 24, 4) */,
  32'h3d302eb0 /* (24, 24, 4) */,
  32'h3d7fc9dc /* (20, 24, 4) */,
  32'h3d836eb0 /* (16, 24, 4) */,
  32'h3d7fc9dc /* (12, 24, 4) */,
  32'h3d302eb0 /* (8, 24, 4) */,
  32'h3d15577e /* (4, 24, 4) */,
  32'h3d139fbd /* (0, 24, 4) */,
  32'h3d37f7fd /* (28, 20, 4) */,
  32'h3d7fc9dc /* (24, 20, 4) */,
  32'h3dd4d413 /* (20, 20, 4) */,
  32'h3defbf1f /* (16, 20, 4) */,
  32'h3dd4d413 /* (12, 20, 4) */,
  32'h3d7fc9dc /* (8, 20, 4) */,
  32'h3d37f7fd /* (4, 20, 4) */,
  32'h3d26b2c0 /* (0, 20, 4) */,
  32'h3d2d4da1 /* (28, 16, 4) */,
  32'h3d836eb0 /* (24, 16, 4) */,
  32'h3defbf1f /* (20, 16, 4) */,
  32'h3e11966c /* (16, 16, 4) */,
  32'h3defbf1f /* (12, 16, 4) */,
  32'h3d836eb0 /* (8, 16, 4) */,
  32'h3d2d4da1 /* (4, 16, 4) */,
  32'h3d1727de /* (0, 16, 4) */,
  32'h3d37f7fd /* (28, 12, 4) */,
  32'h3d7fc9dc /* (24, 12, 4) */,
  32'h3dd4d413 /* (20, 12, 4) */,
  32'h3defbf1f /* (16, 12, 4) */,
  32'h3dd4d413 /* (12, 12, 4) */,
  32'h3d7fc9dc /* (8, 12, 4) */,
  32'h3d37f7fd /* (4, 12, 4) */,
  32'h3d26b2c0 /* (0, 12, 4) */,
  32'h3d15577e /* (28, 8, 4) */,
  32'h3d302eb0 /* (24, 8, 4) */,
  32'h3d7fc9dc /* (20, 8, 4) */,
  32'h3d836eb0 /* (16, 8, 4) */,
  32'h3d7fc9dc /* (12, 8, 4) */,
  32'h3d302eb0 /* (8, 8, 4) */,
  32'h3d15577e /* (4, 8, 4) */,
  32'h3d139fbd /* (0, 8, 4) */,
  32'h3d28c974 /* (28, 4, 4) */,
  32'h3d15577e /* (24, 4, 4) */,
  32'h3d37f7fd /* (20, 4, 4) */,
  32'h3d2d4da1 /* (16, 4, 4) */,
  32'h3d37f7fd /* (12, 4, 4) */,
  32'h3d15577e /* (8, 4, 4) */,
  32'h3d28c974 /* (4, 4, 4) */,
  32'h3d508e8d /* (0, 4, 4) */,
  32'h3d508e8d /* (28, 0, 4) */,
  32'h3d139fbd /* (24, 0, 4) */,
  32'h3d26b2c0 /* (20, 0, 4) */,
  32'h3d1727de /* (16, 0, 4) */,
  32'h3d26b2c0 /* (12, 0, 4) */,
  32'h3d139fbd /* (8, 0, 4) */,
  32'h3d508e8d /* (4, 0, 4) */,
  32'h3dabcc5c /* (0, 0, 4) */,
  32'h3d508e8d /* (28, 28, 0) */,
  32'h3d139fbd /* (24, 28, 0) */,
  32'h3d26b2c0 /* (20, 28, 0) */,
  32'h3d1727de /* (16, 28, 0) */,
  32'h3d26b2c0 /* (12, 28, 0) */,
  32'h3d139fbd /* (8, 28, 0) */,
  32'h3d508e8d /* (4, 28, 0) */,
  32'h3dabcc5c /* (0, 28, 0) */,
  32'h3d139fbd /* (28, 24, 0) */,
  32'h3d234568 /* (24, 24, 0) */,
  32'h3d62e9d3 /* (20, 24, 0) */,
  32'h3d635c6b /* (16, 24, 0) */,
  32'h3d62e9d3 /* (12, 24, 0) */,
  32'h3d234568 /* (8, 24, 0) */,
  32'h3d139fbd /* (4, 24, 0) */,
  32'h3d180196 /* (0, 24, 0) */,
  32'h3d26b2c0 /* (28, 20, 0) */,
  32'h3d62e9d3 /* (24, 20, 0) */,
  32'h3db90e8b /* (20, 20, 0) */,
  32'h3dcd63f0 /* (16, 20, 0) */,
  32'h3db90e8b /* (12, 20, 0) */,
  32'h3d62e9d3 /* (8, 20, 0) */,
  32'h3d26b2c0 /* (4, 20, 0) */,
  32'h3d189328 /* (0, 20, 0) */,
  32'h3d1727de /* (28, 16, 0) */,
  32'h3d635c6b /* (24, 16, 0) */,
  32'h3dcd63f0 /* (20, 16, 0) */,
  32'h3df759b6 /* (16, 16, 0) */,
  32'h3dcd63f0 /* (12, 16, 0) */,
  32'h3d635c6b /* (8, 16, 0) */,
  32'h3d1727de /* (4, 16, 0) */,
  32'h3d044bdf /* (0, 16, 0) */,
  32'h3d26b2c0 /* (28, 12, 0) */,
  32'h3d62e9d3 /* (24, 12, 0) */,
  32'h3db90e8b /* (20, 12, 0) */,
  32'h3dcd63f0 /* (16, 12, 0) */,
  32'h3db90e8b /* (12, 12, 0) */,
  32'h3d62e9d3 /* (8, 12, 0) */,
  32'h3d26b2c0 /* (4, 12, 0) */,
  32'h3d189328 /* (0, 12, 0) */,
  32'h3d139fbd /* (28, 8, 0) */,
  32'h3d234568 /* (24, 8, 0) */,
  32'h3d62e9d3 /* (20, 8, 0) */,
  32'h3d635c6b /* (16, 8, 0) */,
  32'h3d62e9d3 /* (12, 8, 0) */,
  32'h3d234568 /* (8, 8, 0) */,
  32'h3d139fbd /* (4, 8, 0) */,
  32'h3d180196 /* (0, 8, 0) */,
  32'h3d508e8d /* (28, 4, 0) */,
  32'h3d139fbd /* (24, 4, 0) */,
  32'h3d26b2c0 /* (20, 4, 0) */,
  32'h3d1727de /* (16, 4, 0) */,
  32'h3d26b2c0 /* (12, 4, 0) */,
  32'h3d139fbd /* (8, 4, 0) */,
  32'h3d508e8d /* (4, 4, 0) */,
  32'h3dabcc5c /* (0, 4, 0) */,
  32'h3dabcc5c /* (28, 0, 0) */,
  32'h3d180196 /* (24, 0, 0) */,
  32'h3d189328 /* (20, 0, 0) */,
  32'h3d044bdf /* (16, 0, 0) */,
  32'h3d189328 /* (12, 0, 0) */,
  32'h3d180196 /* (8, 0, 0) */,
  32'h3dabcc5c /* (4, 0, 0) */,
  32'h3f800000 /* (0, 0, 0) */};
