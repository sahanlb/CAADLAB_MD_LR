-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
txfmGZ+C+Z4r/dHhJHsOr6jvnuJee1citAowoKkWwsEYRpTxRTRYGIXvW6B/CtM5
xhX7G/AVxuDatttrsqF237UhlE0tHYG2AdWA47NRCuhDm4Djb69pX8+Fe9B7/Gs2
lpY0hhBmmu34vPFEW3EIhDlylxd3WE/VcZk2fkgpwDM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5648)
`protect data_block
alfuXNMoNL5ZB8DYsyUg7eNF5CicEcPpd60vcHjneiPg9MAzUkB/khtMsCzjDS2x
ad6LaOkBQez5jJDFTux+sSABrmxGmgsxy9IIqZ5mer/qNgda4v04xcBMQQr9emi0
xKEqKDZpuTmuaCwEtFdFA9nFY4fVUnaGK21IZEAJVPSXS2XTY1LlTsh42RhNE/2C
BNxhLF5vNX2PMFd3Ec40kA6aw7xdXzYyouq8WMignMHcGOSip588x6cxuupgO2hk
pS0H6MQ69VkGgu/FFIEeelA06MG/zjEtWbVk8hG7s5Gg5Q4/5Z7LqII+lst5K+JT
lNtFd9dTJhjuPMDzwAnh7IlHgH9lHeS3qYeXfoLaUg0w0sF94fS/nMdGEn5rCbpA
q+cpj4CVIKqz1f3qkw4PIzOAnmY0NKku79dkHXpOdSIZVU+XHLlRicCus5n905TP
SvwdqyZz2hYwD6q4Cry5NAI3TkA5sJxFTdJiGeNbPUbsgvkOWBRt5f3OWWQdtoL3
ZqZVTkGzxOlXimr8GDLX9fBNdp203gDYsv+Q4v8HOAuNg1LHoTqtD+yAx5cAdVdg
z9S9ZkwmoljpwWFbXSvmHLMbfgP4QJgOpNAKixIfqSKoX+l5Sm37fVJ3OoSo0Rwv
nUTQGZePczVpKua1BFO49bYgrsFJqr/TBf93Bi5GZa+PQuEVKuL4tZVZ8gXbHyyx
tb7T1ymtAyI6RBbH9OYWYir+MB40CRrbUlM17WUG+Wp1kijVDgmGrATO72MGcc3R
9NoYWjbwWGvwmzqS9i5A5Ou2zcHGx8L4tkqFqn4MK1bfO7H0xKW30deLtaatfI6P
tdX2NWeJaki5Ps10vMNlzVl/t1fKAJ+LR1E7x1/SOzjJkkrxosu2rzozUgDAJEop
jw3DC3gF2ZhuZUYpL+FNTz6tjYKAqPr9Or6GLVRAXrcVVRg8YeMfmFcvuT8EieO8
eQKH4T1OBZG1BEeegPQnNW9DHAhBgOmCNv94x4JJe1RcBkCXgRzgeQ+/3IQBDPcv
DHBxJJG7iEtiv3G+7bUngClTq9/NxQV1WDOQYBC2D9JfnJWV2mCDFkrXQSgsV/E5
4S0Q7AwIhux9CEJgnZqQ2LNO55aSDL92gD2Z+tVwSwlQBan/z3i4bpwlb2YZT9Ol
X2gNvukPXgi9v1zHf47Y1nWO5m9eJSREVlzcz9aYJZIm6A1I+KWzuo9V8K3SvvuJ
6xYgmhbA9kxPh+u3Cj7cGCCcZ03JGlW7JXhntMJ2erwL6clgGiRcXuk0k1t/ymK2
+hNBsJMJf1F1KCfqylqnAOvtHcOQS20PTXdr4CPoDsFxVRwzoe4AiAredt/vkNdg
JIGBD+dOGeiI8TkqpcdquVi+uR/inKVPu5dMe3jKltEL07pJhyJjoGLGGDKKIFaK
Hzu+vnQPTWBUcxoNG1njUxvw8izq6JfZUM0zC8GpBW7Am5lETTCo77MTzI9RXO2z
LKocxoWcfF0Z1qP8vUVcY+x0dOiyqgmXcZg+zMsJ5NcxQByfLxgb/cUirWNflvuD
hqwDcHQqJKSee0iGcIXpHMlOHL/8d8+703QFP0+kaaAxAlLrwG9l+emjmGn9aAc5
ZGyQ2yYsineNRTMsxNEntP7PWy6DQeBUrqgCyeQvJMSKHRPlQCa/c7QYoH3/eCTR
5JbD2l/edkzAYR7q6d6ClelhZalCVPhwr4yC8YltLIFzF58CMimoLLXmSy4YCJyj
C2Fiy5KQBsQ/C3Q7PyBnBjVjnzs1SnNs3lt7h/Hvuyy4HdtVcfbdfasnqXzYRAwR
n7RFrVZAezIdJ7AMoPenudNWNXFYM9j1tFXSyh2Pvke6WJjuFNmhb6kGvCXqBGGK
G9aSjvp4cuKx80pS5mpe9sKx/yEBB2jOtV6oLNzY8i/qj75qyx7DPzHo8bFHQK5g
a7hSdavhYKKqBl57PYSImA0RVGlOBPEY1LhdqQ+V/n1KL82stKeODFGPCXaY1D5c
2f3wXIrchGII7Dp2+4nnY77wLGN107OAMT+izGd/TzA+PVlM9haMEamiN66IyGSj
KKEFHzezAKLXIz6EqeJBmQb5JCxde/UIj6k1ZryhEPg0i4bhR+wMyzgMiPT6GcyT
p6/eaSxIWhzdQcGCh4GoW31rRz4gcgmVMJRt5Yma6XZR6gr5W9tr3/SsmyaC22Hj
Pql0iMaEDDF7OLJuYdVAdTFUTrOfqlfrtvJiA9jrDFWAlp8z6dYI6cdL80F65SZC
PomIZly0gUp/VMSnyLrz2Ln6/TyKx3TNhgtEMaZJEsiPIbpazkf+1XpJl3uAKwp8
ZTyTsLiWaAfYQokFyL1pK2Ej+TfhAUcw3rjxoYe2b+HrMZFWIHYI9I3+piEsACgF
xilyM0Bi4BU+mfIhhSGHwzXQkLAfPHRE+rCMJ0sYWg9tfq8xocfHHvOsQbleJohr
kqjZmpAp90FGh+0KY7Mt2pM2KoC47V5gSrgPg3Bh5ef+auoODWPA2n920aKcjTL6
J7CspSa+1KrF2T5rlR4w1pM2mFymKmVEy1I0y7xV0+NfunoXGGTDQqsFxkLlm1BY
ccAKG94O8Ns3L6ThPnOJRTDTjVNEp/4BNf3Hcl2/ZJepqW5d2ByoV0cAkVp5VBU9
YXAKR66LbNX+4BNxXRztJr7Z8C0G25t3dmPJHUhNHPDwaqXXKTcRxndNUbsVXHpI
5nXZA9/xECUrrSWtP4p6xfErkeBJq/i0ZSZWku/PwRVvx1OF1wOzHQXk9kLW2pJJ
OSaxmrLzTAeDCFBfPLrOb1bDgMWEpAP0dH0lUqpUQqZ5E6wq6Ihgj4jTVS8iyUZw
gZWwmV7QjI31syiW+QETZNcZgSSrjA/5BGKrWp6G3s4V5WOF0k8tLVwNApIUGcGW
L+7CMZaFGMRrnq9zccnzPvMRMkc/tTc0EbukUIDngiJy3VQt/HIcWJcHAlx4eNGh
0bbzHZS3FeC1xZfIH9k666Iyh9jbsEMpZEX8xXEVOVFWJHCbIsK6nSfJOCj9JQmo
/IJhvETWyMXbCzOJ3VA3kGJg3GM/zsMt7XZxNag02PWfTlchy8h89Tvqe9wP+YTw
zR/rT+lSh0SQNwefPrVjvkzqm9wzJi6sP2JD5o/sw1KNaMrZoy1xjbzIrybmeXPJ
lAt3pkh65uTJM98hxfG9lZ7p4Y8uQyRgzguQzD/b96TC3SfsJDu78mxrdb5iRvVY
N/VFOG/e/Ybk28Tj8bL2DoEBi4RGy8Bp96nHA3BVv8NcisEP/0bl9hkj617m4hlv
zfr7EEcdot1G4zx5LIn+IJNSUbVjF6rYNEC3NWzu42DlsrrrZntLL1mGDjTpjH6A
OB+NN8ATMThMeA1c22CFhtNCXxfCe5IwlCRXaZpwne9YaYAXHp/V72oKzu/BBPiZ
eb3g7dzmylz5aswQhIKjW1pvLiNTSoUXwFgdD1PDcR/khTytWXA9lswjvXbSWFQi
fb/EJPdRULGMI78urhQctWd3Gep44vF8IgdNPmWtB4D9m8R8OxHrS6e6JvqvwARm
uF40ES0/eT0PbU93Sl+VosSm8fWiAwCyuP5xl6x54dJTylx+ZG4xJXjUOFkxMzfH
7YOm8s6HDizsncveV1OcaawYNf172L8/7MnLPdcCWI9i/Mp+Sc2swUhgTmzO2Uwx
3mv7r0EoFjrBNGjJ2uys7UU8LPKwx1mu7psu9gJTIKEKx0iKyJq6dLBP0+5Pu82m
L5apIqogo5CF/WoMaF/I3FWeyIs0tGEELseDXARI+JLh0e7jSPn7FNIyf8Ph6XO9
x7OzQvz22gPvO5Zvenb4Ytf2K4WMmXmHm2iBhOgaXo8U0iFQn92VJmJipzhLJZZ/
iEpYCPxeaGe8aDA4o9vV/gie3FzHQ1+YQ7YOVsAKmZOvTFbUP3PfHihXoEni84D2
jHlpA3EC45aL0MtrtdTNYBW5LmgS9UYxU1UsRT2Vw451qfdgst5fP+6Rv3b39uCu
6Zxcsyn1iTfl0kFZBJpVeOLqhVNv8WCen3UJ2DkHz/U3aE5uB+U6CFKgpZblOenX
21DsVFfwNUX8BqIaASFzGbC7ff2i9v2aNNOU2qPtfTzOkKvG80N6RRbUjpBWCHT2
yzIcBaMR3UwKjFiB/cfGwQLtSO99mm4rEBeNVcC1Uhq0Ah5pe3enZ1408a+JFO4w
384BTy+dEjYZPNKzhrHjEXbFS2JTXcrJTWOKcfUlm37N6vTS5980+Bduzwauy3Zr
y2F9SlKCgPva890/hRnLCaWQ45fNuQdv5/gMDxmb+2RU7FJXMD+aY/x7/h5k/McS
V3JcUvXkpZJ/xZGsz1Y9iJkm482uKQZs182kr7lwVpE//SdK9IsyeVJErutQL7wx
7owW/R9ewcbOjbP/M2tw9NrqYDgGA1oMJO7ne331bMiCMSdmnX5n7yvaAtcDe45S
xvReN8QA/JcHXWzwmzVjLSD4wiTh/zP/oV2lX+Jh1CLbAgZvYWp7D1VgNcmgGa+T
qm9dpB3dmVGX4offnmvxL5gPDPM2VbZqVkvTiayz436uOxtnWebfiHJdhox96ix9
oHVFOSV2qbLTtlpM3hHGlpbY9zqsh+vuOm8LadTAmUU+FQrZLdk0fmlKMuzBiNJE
GMVmFrsNRohbjd2FWIlhEjFeTju2iHGl56+Ej+3eYewWwtGo1sJLQEXONVGDJ2Rt
J9rZ63+MTj6t/UFNve4BujRrq3gXBkY6oTdEnnnG8M2uPGMH+fd6PxwZWZoyCTnw
k+yXHy1ilmJXdPCsdI9GUZjdb0QAZ4h+RfFO0cRKp+mMuOKMhDPcGM7oSwS6uWz/
bIMbLkx0+imc4ArXAuAFTYZ6ei6Su5uMxnaJky6uKfEFPgggHCLaekB4afGXTrTE
ivPsZbkvGC/nQE6OqfNXanmNBSEFpQFlkE5Bm3XekSwOPrMxD9iKe7uJuO/m9WCC
Zqi4DU0GibduLyr1t37avDXHzvd+QIZuud1Go6DqMZ2BXqFG4glMHpp/3DNZFrPj
Ft9hFlPiUmgh/qnbRgwJYKpUlCtczwxwplF4irkZ/iTrIS909Q7A0ssMOZGcKzvh
9r1xQn0E/aoK3AphFg+ly2x2PN+tmfYRouBSSvty5qOY2xlIufBo3LXutP7CMLoP
R32uLjBibUn4+92FJuPMCdk8B/4dR7nGTIB829hHVYruHPKCidLklBAMLe11K8G5
4jvz2YjIjWOqO81Zo7PDBl68wIlpvw5qoMiUgITxVKlc8ROB1fJr1+KgzIcAZT81
KJIcrqr+/14jR/nr1cUDfq/2QNMNqihTmPjQOuON8FJPCbUylxczuP0BsxM/gfp9
vmAvfk4ZbAt7AB5sCvQOpfELXhXjzMvZn5bfBSiVdgn/tIRliUgvvWfyNKy578zX
9CPIYxUjRb525cE1xI5EvyKYJtuvzBqRqbMiI42q4Jjw2+tEISiLU8pcOOFengxT
XBu3jSweHSxLwDP+VRgi136qObaidtAAy4X49IEvTxyY+EMLI/CsZkrT+/eD6+uq
vRUvDHDtTqw8uQ0yE9cEsefCFk1MQ5MuzrK+gsnMM83Dc8OB8NF7iVi4rCtPRWOE
58kOl4FrRdWsI9DpC5WvmDb7mIKzlh8vW/zRcft6djU16WF/KR1WWajxxVyaWkZ3
8Z0nmsS/lOxI51QhkFSfzAuFeipH/kAHuitGttaDN+xg14B9vwABkJVPH60uyFBo
8e8H87hfgxj7hMHmou06sd+Kng4YCT3UJYUea0cxaQiGaelKFMlWKV86hNtUL3Lp
oYtc+YBfjtWLKzUOptjN2eqT8ATF7FWhQGJxQVyTWwvoq5kSkwUqzXh33ZE50ZxC
0T7YKuCXJmbWRKInbNTzA6Yv37utSjvPlu19C21d+MBlDosmdT1MvBSy4w/gUT95
Oml5Q7C8L15YDc61dgUecayrQ99uvbAHglmVU8u69grFuAU2hLwCdA4z9FpS5QjZ
rASOUqA331qSz1cxVFNttC1rEI6EGE8vOfS+muy7kNM7YVdSem/am5SIgyp7TIsy
2MRF9LUaptZ+teEds2M2TpkIJd0HOGMVmvQRiGR5YGEdiu8Yf4WqXqD4Ka6i8pyZ
WN+mcys0ygfBT04x6K8JEbW4S77sPn05bVPvJSe5onMyqDOx4RbmfgE+Vo2Hetyb
hH4OzFaMEI4n2Rl6ZG5kc48ZUbtur4Y+dv04qjRo6/6jS9CGLbcMCkLatyqX2p5I
8lcspqd0lB601fcsLDSqd4fAXeuwzS+tbpuWwJWlu/urWjgkvy+87w9n3lB4NQcl
5H8Xh5uZDfCO77m+p0vNzPXCpaYyF1Rl/Ld3CuhN2HNJZbK1FWv6bQnbxz2xwTQI
F0JT06KmUxn6X+AFetEmdJ0A+vk7lIoCJ06TbjDt103zD30jdiii1C7+6dZLu0TD
3GVGC1Im/0ZEz7ZKbr8YDc8l5b1Gr3fSpgOGb1dRmbydvfD7sVf4OGhrCCIgeCiX
HnD+hJKKjUcpubmplOIzatygf2eMbyPZ11WZ32YriKUa4tnqyyEBWdvdIk1gE1cC
StC9xhxHuw+14AHAvkdIl1QNnNzCJaxmSVv6yvXcYZiHjYkUwi3CK1KVUattdU17
/iKoxEpEqq9nRs+/B3teSkgZbJ8uesaSri9dK+oOa0MZ13MljU0dT2hymjqPh/HJ
EU8xVA6ir7WU2ZM/BN3aC1eyEcEG1IX4Xidz1yxKtDibBh+jJ6ZodfH5y16ypBEi
x7msej2xVziyWMEnDJYtDSrlnrVRaLN7V7KewqCLu5do0iTP2hq2YRouIc46pckx
gbehEfyyVskLNlXlW77aOdXsR4nYNNuP3XWuR8wza5ef6AOmugaO8usfTZXgXRC3
i23ZQeBW2bsHg4Cu/shhb/TCehHuZCnx5kzSte2VL+CtXIdm0PIS4kePK2xCWpqw
TL88gWLUwmNfY3ZHomncYsqGMTymOEg1RjIFUAq/JxzKRzrWmrBOjSJFwf1iuw9V
gYKCo3GSkoJjJMc1opxQ9VYGprMUa9ZgiMGyRzn3wSHNOp5Ekd5yuSw1oCwBbE5+
LvblNXlxg2447w2JAoluyUn7q4PIRnBax97mOjoK6+SWAI6OonzLuh+DDfW5vE/N
sjWaz8WST6AT3GeK4GR6kiMiM2baUlqoVQ33u2v0JF/5FRr/FJLHChsU8gbKwtUI
JxBKrRvTR27pjepYOI31lim8jSKEfEQIQq17kGFFpjyIySSsy1uVVs+V/TgeJsqM
y4T+f6aSPcQJiKrxJEHjKHHglCpE48W4//76eZd/iEVTpev1CdUB5Srz4fJ20LGB
SUjLNkCftglEYNHhgg0d+UIUATFYdu5eigH62iabBZIYSvj/TXrO0qDsb3fQoIXX
2lla3VgTAb1hyr/FdXae7agmnkYP87AcKUoSLe4oPeI86YR4+vDUAoGe2QhB51uA
TQPOqbrOdQPVYaUWtKeir4U4xmW7wjKOud+b31p21hBKp53F6umFYIX9p3U1fm28
pjJ4VOLbi+D8w2CRdRvcshzJA5F9U+9+4t2mtXLv7FQ=
`protect end_protected
