localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTX_CHK = {
  {32'h3f3e33ba, 32'h40406ff4} /* (31, 31, 31) {real, imag} */,
  {32'h3df0f9d4, 32'h40f3cc9e} /* (31, 31, 30) {real, imag} */,
  {32'hbe930cb6, 32'h40c28aa6} /* (31, 31, 29) {real, imag} */,
  {32'hbf3aa0a1, 32'h408a903e} /* (31, 31, 28) {real, imag} */,
  {32'h3da09cb4, 32'h4089860d} /* (31, 31, 27) {real, imag} */,
  {32'hbe03f53e, 32'h40a25dba} /* (31, 31, 26) {real, imag} */,
  {32'h4018811e, 32'h408b8e38} /* (31, 31, 25) {real, imag} */,
  {32'hbed25468, 32'h40a37598} /* (31, 31, 24) {real, imag} */,
  {32'hbf8f21b5, 32'h40a48d23} /* (31, 31, 23) {real, imag} */,
  {32'hbf5c8ddd, 32'h40d2a772} /* (31, 31, 22) {real, imag} */,
  {32'h3f60a13c, 32'h402eff23} /* (31, 31, 21) {real, imag} */,
  {32'h3fa1f960, 32'hc05c68f2} /* (31, 31, 20) {real, imag} */,
  {32'h3fb7bf2e, 32'hc0675295} /* (31, 31, 19) {real, imag} */,
  {32'hbe7cb3c4, 32'hc0824455} /* (31, 31, 18) {real, imag} */,
  {32'h3e8919da, 32'hc0474011} /* (31, 31, 17) {real, imag} */,
  {32'hbe508a40, 32'hc0b2d2b2} /* (31, 31, 16) {real, imag} */,
  {32'h3f7df615, 32'hc0beb4d2} /* (31, 31, 15) {real, imag} */,
  {32'h3f6a5189, 32'hc08d614f} /* (31, 31, 14) {real, imag} */,
  {32'h3fb4254a, 32'hc086056e} /* (31, 31, 13) {real, imag} */,
  {32'hbef07825, 32'hc0922bbe} /* (31, 31, 12) {real, imag} */,
  {32'h3ebb1666, 32'hc03ae851} /* (31, 31, 11) {real, imag} */,
  {32'h3d6c1b4c, 32'h408647cc} /* (31, 31, 10) {real, imag} */,
  {32'h3f3f4f88, 32'h4036def2} /* (31, 31, 9) {real, imag} */,
  {32'h401dae88, 32'h406702fd} /* (31, 31, 8) {real, imag} */,
  {32'h3f65fc5a, 32'h40826525} /* (31, 31, 7) {real, imag} */,
  {32'hbfdf4916, 32'h408f9dfd} /* (31, 31, 6) {real, imag} */,
  {32'hbd618a90, 32'h4093e12f} /* (31, 31, 5) {real, imag} */,
  {32'h3edf7962, 32'h405b6c55} /* (31, 31, 4) {real, imag} */,
  {32'h3f2036d2, 32'h402acd4c} /* (31, 31, 3) {real, imag} */,
  {32'h3d01148c, 32'h3fd78983} /* (31, 31, 2) {real, imag} */,
  {32'h3f45a380, 32'h407e3bdc} /* (31, 31, 1) {real, imag} */,
  {32'h3f338ca5, 32'h4020666a} /* (31, 31, 0) {real, imag} */,
  {32'h3f8d8e6a, 32'h4091158a} /* (31, 30, 31) {real, imag} */,
  {32'h403c8724, 32'h41299a68} /* (31, 30, 30) {real, imag} */,
  {32'h4099d85c, 32'h411dd9f7} /* (31, 30, 29) {real, imag} */,
  {32'h40064a5e, 32'h40de3687} /* (31, 30, 28) {real, imag} */,
  {32'h4030b5c6, 32'h409c984a} /* (31, 30, 27) {real, imag} */,
  {32'h3f3ff99e, 32'h40a421e6} /* (31, 30, 26) {real, imag} */,
  {32'h3f6694fc, 32'h40d209dd} /* (31, 30, 25) {real, imag} */,
  {32'h3e6152cd, 32'h411fb032} /* (31, 30, 24) {real, imag} */,
  {32'h3f8c2a69, 32'h40f24654} /* (31, 30, 23) {real, imag} */,
  {32'h3e9aa86e, 32'h411f393e} /* (31, 30, 22) {real, imag} */,
  {32'h401fbec6, 32'h405a5ef2} /* (31, 30, 21) {real, imag} */,
  {32'hbebe9b8e, 32'hc1171088} /* (31, 30, 20) {real, imag} */,
  {32'hbf9033c6, 32'hc10006e9} /* (31, 30, 19) {real, imag} */,
  {32'hbfa51a8a, 32'hc11a2e18} /* (31, 30, 18) {real, imag} */,
  {32'hbf08c376, 32'hc0d4fb80} /* (31, 30, 17) {real, imag} */,
  {32'hbf5e4760, 32'hc1199259} /* (31, 30, 16) {real, imag} */,
  {32'hbfacd556, 32'hc114fa20} /* (31, 30, 15) {real, imag} */,
  {32'hc090f5c8, 32'hc10ed162} /* (31, 30, 14) {real, imag} */,
  {32'hc07135ae, 32'hc1049922} /* (31, 30, 13) {real, imag} */,
  {32'hbfb0b31e, 32'hc0df1bd8} /* (31, 30, 12) {real, imag} */,
  {32'hbfaa849c, 32'hc08745be} /* (31, 30, 11) {real, imag} */,
  {32'hc0627ba0, 32'h4096b352} /* (31, 30, 10) {real, imag} */,
  {32'h3e1d8cf2, 32'h409ffdca} /* (31, 30, 9) {real, imag} */,
  {32'h404a156a, 32'h41082ec6} /* (31, 30, 8) {real, imag} */,
  {32'h3fc58f4b, 32'h40e1fb70} /* (31, 30, 7) {real, imag} */,
  {32'hc016c686, 32'h40b3456b} /* (31, 30, 6) {real, imag} */,
  {32'hbfbe3c6e, 32'h40f8dbff} /* (31, 30, 5) {real, imag} */,
  {32'h3fb080d4, 32'h40cf08b4} /* (31, 30, 4) {real, imag} */,
  {32'h4029ab14, 32'h40b9f85c} /* (31, 30, 3) {real, imag} */,
  {32'h3fca2fa0, 32'h40d2f373} /* (31, 30, 2) {real, imag} */,
  {32'h3ff7440c, 32'h410a2035} /* (31, 30, 1) {real, imag} */,
  {32'h3f80fb6e, 32'h4080f559} /* (31, 30, 0) {real, imag} */,
  {32'h3fe26e4e, 32'h40a1a97a} /* (31, 29, 31) {real, imag} */,
  {32'h400e7512, 32'h411d636e} /* (31, 29, 30) {real, imag} */,
  {32'h3ff23e4d, 32'h40c08b68} /* (31, 29, 29) {real, imag} */,
  {32'h3fe52446, 32'h40a0dd0a} /* (31, 29, 28) {real, imag} */,
  {32'h3ee5d564, 32'h409fceba} /* (31, 29, 27) {real, imag} */,
  {32'hbfd9e8f8, 32'h40c34258} /* (31, 29, 26) {real, imag} */,
  {32'h3ea06c74, 32'h40d5e27c} /* (31, 29, 25) {real, imag} */,
  {32'h402e894c, 32'h40cf07ba} /* (31, 29, 24) {real, imag} */,
  {32'h3fa7ba30, 32'h40c518de} /* (31, 29, 23) {real, imag} */,
  {32'hbf80e7e5, 32'h4106ca24} /* (31, 29, 22) {real, imag} */,
  {32'hbff032b0, 32'h40a9426b} /* (31, 29, 21) {real, imag} */,
  {32'hc0ac7af6, 32'hc102ace9} /* (31, 29, 20) {real, imag} */,
  {32'hbfb1637b, 32'hc0f568ee} /* (31, 29, 19) {real, imag} */,
  {32'hc028bbca, 32'hc1189014} /* (31, 29, 18) {real, imag} */,
  {32'hc05b5cc9, 32'hc0c049cc} /* (31, 29, 17) {real, imag} */,
  {32'hbfb1a6ad, 32'hc0b0a810} /* (31, 29, 16) {real, imag} */,
  {32'hbfe8500a, 32'hc0fbf634} /* (31, 29, 15) {real, imag} */,
  {32'hc08de528, 32'hc0e26604} /* (31, 29, 14) {real, imag} */,
  {32'hc0b22285, 32'hc0e85e0f} /* (31, 29, 13) {real, imag} */,
  {32'hc00f2632, 32'hc0cc3302} /* (31, 29, 12) {real, imag} */,
  {32'hc02bc2b6, 32'hc0933b41} /* (31, 29, 11) {real, imag} */,
  {32'hc0a78254, 32'h3f9b741e} /* (31, 29, 10) {real, imag} */,
  {32'hbee0b086, 32'h408b8a6c} /* (31, 29, 9) {real, imag} */,
  {32'h408b2f2e, 32'h41218358} /* (31, 29, 8) {real, imag} */,
  {32'h3fc69bb2, 32'h4112e0c7} /* (31, 29, 7) {real, imag} */,
  {32'hbeda995b, 32'h40a87132} /* (31, 29, 6) {real, imag} */,
  {32'hc0023d00, 32'h40963c0a} /* (31, 29, 5) {real, imag} */,
  {32'hbef64539, 32'h406159ae} /* (31, 29, 4) {real, imag} */,
  {32'h401b25c3, 32'h40c4c8d8} /* (31, 29, 3) {real, imag} */,
  {32'h3ff46b51, 32'h410f2413} /* (31, 29, 2) {real, imag} */,
  {32'h3ed9a390, 32'h413f422c} /* (31, 29, 1) {real, imag} */,
  {32'h3fad3bb1, 32'h4092e6aa} /* (31, 29, 0) {real, imag} */,
  {32'h3fe6fd5a, 32'h40ae522a} /* (31, 28, 31) {real, imag} */,
  {32'h3f804398, 32'h41061616} /* (31, 28, 30) {real, imag} */,
  {32'hbe106590, 32'h40cbd3fd} /* (31, 28, 29) {real, imag} */,
  {32'h3fa4163f, 32'h40c2e2f5} /* (31, 28, 28) {real, imag} */,
  {32'hbf46b255, 32'h40b7b5f2} /* (31, 28, 27) {real, imag} */,
  {32'hbf8078fe, 32'h40ce4218} /* (31, 28, 26) {real, imag} */,
  {32'h4066aeeb, 32'h41116fcc} /* (31, 28, 25) {real, imag} */,
  {32'h40baf834, 32'h41253f2e} /* (31, 28, 24) {real, imag} */,
  {32'h3f60cd8a, 32'h412bd523} /* (31, 28, 23) {real, imag} */,
  {32'hc005db3d, 32'h412279cf} /* (31, 28, 22) {real, imag} */,
  {32'hbee260b2, 32'h40c8926e} /* (31, 28, 21) {real, imag} */,
  {32'hbfbad340, 32'hc07c24c3} /* (31, 28, 20) {real, imag} */,
  {32'hbe2b2f11, 32'hc0c90ddf} /* (31, 28, 19) {real, imag} */,
  {32'hc0094472, 32'hc132ae34} /* (31, 28, 18) {real, imag} */,
  {32'hbf4d0dbf, 32'hc10f0788} /* (31, 28, 17) {real, imag} */,
  {32'hbd1df618, 32'hc107abea} /* (31, 28, 16) {real, imag} */,
  {32'hc068b29c, 32'hc124d76f} /* (31, 28, 15) {real, imag} */,
  {32'hc09c91ab, 32'hc1059ce8} /* (31, 28, 14) {real, imag} */,
  {32'hc080ba32, 32'hc0ac4f79} /* (31, 28, 13) {real, imag} */,
  {32'hbfb9fa06, 32'hc0ee52e0} /* (31, 28, 12) {real, imag} */,
  {32'hc00c5b4e, 32'hc0f07383} /* (31, 28, 11) {real, imag} */,
  {32'hbec9143e, 32'h3fd2f5b0} /* (31, 28, 10) {real, imag} */,
  {32'h3fd79bee, 32'h40c53143} /* (31, 28, 9) {real, imag} */,
  {32'h3fbe7681, 32'h40ec81b8} /* (31, 28, 8) {real, imag} */,
  {32'h3faf62e8, 32'h40ea3220} /* (31, 28, 7) {real, imag} */,
  {32'h4010d493, 32'h40e1f2b9} /* (31, 28, 6) {real, imag} */,
  {32'hbec3bb45, 32'h4108eeec} /* (31, 28, 5) {real, imag} */,
  {32'h3dc39caa, 32'h411e3d1e} /* (31, 28, 4) {real, imag} */,
  {32'h401456f4, 32'h4112ed8e} /* (31, 28, 3) {real, imag} */,
  {32'h404d5afa, 32'h41003eab} /* (31, 28, 2) {real, imag} */,
  {32'h4001fa5b, 32'h4114890f} /* (31, 28, 1) {real, imag} */,
  {32'h3f936de9, 32'h40895519} /* (31, 28, 0) {real, imag} */,
  {32'h40286a18, 32'h40aa60b7} /* (31, 27, 31) {real, imag} */,
  {32'hbf2805a4, 32'h410b2b08} /* (31, 27, 30) {real, imag} */,
  {32'hc01f7092, 32'h41191bfe} /* (31, 27, 29) {real, imag} */,
  {32'hbf04da33, 32'h40e968cb} /* (31, 27, 28) {real, imag} */,
  {32'h3f2bc5ca, 32'h40f568d0} /* (31, 27, 27) {real, imag} */,
  {32'h3faa2744, 32'h4128ef7c} /* (31, 27, 26) {real, imag} */,
  {32'h3ed9972b, 32'h412c8f1b} /* (31, 27, 25) {real, imag} */,
  {32'h400d96b7, 32'h4133cd78} /* (31, 27, 24) {real, imag} */,
  {32'hbead19a1, 32'h41367e68} /* (31, 27, 23) {real, imag} */,
  {32'hbfff158a, 32'h4100a812} /* (31, 27, 22) {real, imag} */,
  {32'h3f8ca4ae, 32'h404b712c} /* (31, 27, 21) {real, imag} */,
  {32'h4003c7bc, 32'hc07a8483} /* (31, 27, 20) {real, imag} */,
  {32'h401b7c2c, 32'hc0e34cdd} /* (31, 27, 19) {real, imag} */,
  {32'hbea8b4a0, 32'hc115ee26} /* (31, 27, 18) {real, imag} */,
  {32'hbedd594c, 32'hc118890b} /* (31, 27, 17) {real, imag} */,
  {32'hbed91f6a, 32'hc12b0334} /* (31, 27, 16) {real, imag} */,
  {32'hbf826200, 32'hc114ed43} /* (31, 27, 15) {real, imag} */,
  {32'hc05ed63c, 32'hc106ade9} /* (31, 27, 14) {real, imag} */,
  {32'hc04a02ce, 32'hc0d1fbfa} /* (31, 27, 13) {real, imag} */,
  {32'h3f3310b0, 32'hc0e5ad19} /* (31, 27, 12) {real, imag} */,
  {32'h40157cdd, 32'hc10a392f} /* (31, 27, 11) {real, imag} */,
  {32'h402ccc1c, 32'h3f83751d} /* (31, 27, 10) {real, imag} */,
  {32'h409102a7, 32'h4119d613} /* (31, 27, 9) {real, imag} */,
  {32'h40745090, 32'h410d646b} /* (31, 27, 8) {real, imag} */,
  {32'h406fb87c, 32'h41003f7c} /* (31, 27, 7) {real, imag} */,
  {32'h3fe5a972, 32'h41096692} /* (31, 27, 6) {real, imag} */,
  {32'h401424a0, 32'h413c9936} /* (31, 27, 5) {real, imag} */,
  {32'h40587ff3, 32'h416180d3} /* (31, 27, 4) {real, imag} */,
  {32'h40064d51, 32'h4111e618} /* (31, 27, 3) {real, imag} */,
  {32'h3faf2f84, 32'h40ca4951} /* (31, 27, 2) {real, imag} */,
  {32'h3fee6d36, 32'h40f5f82e} /* (31, 27, 1) {real, imag} */,
  {32'h3ea1c760, 32'h40b04fe7} /* (31, 27, 0) {real, imag} */,
  {32'h3fe30119, 32'h4073f22c} /* (31, 26, 31) {real, imag} */,
  {32'hbf8cd09c, 32'h4103f50d} /* (31, 26, 30) {real, imag} */,
  {32'hc059e721, 32'h41499391} /* (31, 26, 29) {real, imag} */,
  {32'hbfc535eb, 32'h41320b80} /* (31, 26, 28) {real, imag} */,
  {32'h400cf535, 32'h411c55db} /* (31, 26, 27) {real, imag} */,
  {32'h4002fbf6, 32'h4140a36b} /* (31, 26, 26) {real, imag} */,
  {32'hbff7c4e7, 32'h41491e84} /* (31, 26, 25) {real, imag} */,
  {32'h40090f22, 32'h41072ed2} /* (31, 26, 24) {real, imag} */,
  {32'h3f0c9cac, 32'h40dc41b8} /* (31, 26, 23) {real, imag} */,
  {32'hbef6efd7, 32'h40efac28} /* (31, 26, 22) {real, imag} */,
  {32'h3f7b8df8, 32'h408444e8} /* (31, 26, 21) {real, imag} */,
  {32'h3f410203, 32'hc04f2f8c} /* (31, 26, 20) {real, imag} */,
  {32'h3f230e8c, 32'hc10aa014} /* (31, 26, 19) {real, imag} */,
  {32'hbea7fdd7, 32'hc0eabbbc} /* (31, 26, 18) {real, imag} */,
  {32'h3f2e3908, 32'hc0f826b4} /* (31, 26, 17) {real, imag} */,
  {32'h3f87fffa, 32'hc11b68e2} /* (31, 26, 16) {real, imag} */,
  {32'hbfd7368d, 32'hc0b8fa7d} /* (31, 26, 15) {real, imag} */,
  {32'hc04041df, 32'hc0f38238} /* (31, 26, 14) {real, imag} */,
  {32'hc077a4e1, 32'hc10f47ec} /* (31, 26, 13) {real, imag} */,
  {32'hbf514abe, 32'hc0c3c0d6} /* (31, 26, 12) {real, imag} */,
  {32'h3d205250, 32'hc09062ce} /* (31, 26, 11) {real, imag} */,
  {32'h3fbf4df1, 32'h40bfd2f3} /* (31, 26, 10) {real, imag} */,
  {32'h40070209, 32'h414d53f1} /* (31, 26, 9) {real, imag} */,
  {32'h406ec56d, 32'h4129f7bd} /* (31, 26, 8) {real, imag} */,
  {32'h40176ae6, 32'h412826e2} /* (31, 26, 7) {real, imag} */,
  {32'h3f77631c, 32'h40f5ba39} /* (31, 26, 6) {real, imag} */,
  {32'h400c50c8, 32'h40d9145d} /* (31, 26, 5) {real, imag} */,
  {32'h400fca36, 32'h4112443a} /* (31, 26, 4) {real, imag} */,
  {32'h3f4a9f86, 32'h40edd56d} /* (31, 26, 3) {real, imag} */,
  {32'h3ef35f05, 32'h40e9466f} /* (31, 26, 2) {real, imag} */,
  {32'h401453e3, 32'h4116a864} /* (31, 26, 1) {real, imag} */,
  {32'h3fa4d427, 32'h40b85ea7} /* (31, 26, 0) {real, imag} */,
  {32'h3fb3afb5, 32'h40a0f3b0} /* (31, 25, 31) {real, imag} */,
  {32'h3f29415f, 32'h410eb610} /* (31, 25, 30) {real, imag} */,
  {32'hbfd3151e, 32'h4129e9fa} /* (31, 25, 29) {real, imag} */,
  {32'hc02b4110, 32'h412f22a7} /* (31, 25, 28) {real, imag} */,
  {32'h400da622, 32'h410d41f6} /* (31, 25, 27) {real, imag} */,
  {32'h404c428e, 32'h410c05b6} /* (31, 25, 26) {real, imag} */,
  {32'hc028fca2, 32'h412779e4} /* (31, 25, 25) {real, imag} */,
  {32'hbfa815c2, 32'h40f313d6} /* (31, 25, 24) {real, imag} */,
  {32'h3f8ee2fa, 32'h40a41b1f} /* (31, 25, 23) {real, imag} */,
  {32'h3f475121, 32'h40ced002} /* (31, 25, 22) {real, imag} */,
  {32'h3ecc40bc, 32'h40853b64} /* (31, 25, 21) {real, imag} */,
  {32'hbf17f57c, 32'hc0a24d44} /* (31, 25, 20) {real, imag} */,
  {32'hbe1c7110, 32'hc12130e0} /* (31, 25, 19) {real, imag} */,
  {32'h3fa4aff6, 32'hc10dae24} /* (31, 25, 18) {real, imag} */,
  {32'h3fd9d589, 32'hc12070b6} /* (31, 25, 17) {real, imag} */,
  {32'h40522e7c, 32'hc11d6f3a} /* (31, 25, 16) {real, imag} */,
  {32'hbf7a0346, 32'hc0985339} /* (31, 25, 15) {real, imag} */,
  {32'hc07e2e62, 32'hc0f26b04} /* (31, 25, 14) {real, imag} */,
  {32'hc037e23e, 32'hc13148dc} /* (31, 25, 13) {real, imag} */,
  {32'hc031c6b6, 32'hc0ffa739} /* (31, 25, 12) {real, imag} */,
  {32'hbfc71602, 32'hc017da24} /* (31, 25, 11) {real, imag} */,
  {32'h3ff3892e, 32'h41079c7c} /* (31, 25, 10) {real, imag} */,
  {32'hbf9ea37e, 32'h414937d3} /* (31, 25, 9) {real, imag} */,
  {32'hbed686b4, 32'h410d218a} /* (31, 25, 8) {real, imag} */,
  {32'h3f2933b6, 32'h4101504f} /* (31, 25, 7) {real, imag} */,
  {32'h3f2fe4bc, 32'h40e8161a} /* (31, 25, 6) {real, imag} */,
  {32'h3e7779d4, 32'h40d70052} /* (31, 25, 5) {real, imag} */,
  {32'hbf3ac76a, 32'h4102c86c} /* (31, 25, 4) {real, imag} */,
  {32'hbec234b6, 32'h410c669d} /* (31, 25, 3) {real, imag} */,
  {32'h3efca8ef, 32'h410a7408} /* (31, 25, 2) {real, imag} */,
  {32'hbf2f815f, 32'h4116a046} /* (31, 25, 1) {real, imag} */,
  {32'hbfb6842b, 32'h408c47e6} /* (31, 25, 0) {real, imag} */,
  {32'h3dd67418, 32'h40722b44} /* (31, 24, 31) {real, imag} */,
  {32'h3fe028ee, 32'h40dc5ef8} /* (31, 24, 30) {real, imag} */,
  {32'hbf475944, 32'h40b2648e} /* (31, 24, 29) {real, imag} */,
  {32'hc00f14e6, 32'h410aa046} /* (31, 24, 28) {real, imag} */,
  {32'h3fe27fc2, 32'h40ddbf10} /* (31, 24, 27) {real, imag} */,
  {32'h402c91ed, 32'h40901bbe} /* (31, 24, 26) {real, imag} */,
  {32'hbd86acf4, 32'h40e486e2} /* (31, 24, 25) {real, imag} */,
  {32'h3e0e781c, 32'h40e11f44} /* (31, 24, 24) {real, imag} */,
  {32'h4063baab, 32'h40c4401d} /* (31, 24, 23) {real, imag} */,
  {32'h40266d6c, 32'h40f67ec0} /* (31, 24, 22) {real, imag} */,
  {32'h400a372d, 32'h40836a4e} /* (31, 24, 21) {real, imag} */,
  {32'hbcd3afe0, 32'hc0df4f65} /* (31, 24, 20) {real, imag} */,
  {32'hbfdceb0e, 32'hc10bc4c6} /* (31, 24, 19) {real, imag} */,
  {32'h3f1244e4, 32'hc0dd5787} /* (31, 24, 18) {real, imag} */,
  {32'h3e9e62a3, 32'hc10fbd9a} /* (31, 24, 17) {real, imag} */,
  {32'hbde2d010, 32'hc10cbcca} /* (31, 24, 16) {real, imag} */,
  {32'hbf668b19, 32'hc0f14e5e} /* (31, 24, 15) {real, imag} */,
  {32'hc013e0bd, 32'hc0e7a852} /* (31, 24, 14) {real, imag} */,
  {32'h3f11ad4d, 32'hc1187580} /* (31, 24, 13) {real, imag} */,
  {32'hbf2fd0c3, 32'hc1006caa} /* (31, 24, 12) {real, imag} */,
  {32'h3fad57e9, 32'hc0286abd} /* (31, 24, 11) {real, imag} */,
  {32'h3fdd1c04, 32'h40e86704} /* (31, 24, 10) {real, imag} */,
  {32'hbe55182c, 32'h412569ee} /* (31, 24, 9) {real, imag} */,
  {32'h40244481, 32'h4105d348} /* (31, 24, 8) {real, imag} */,
  {32'h4028aaf6, 32'h4111a38d} /* (31, 24, 7) {real, imag} */,
  {32'h4048ef0c, 32'h40fb8250} /* (31, 24, 6) {real, imag} */,
  {32'h3f4b4015, 32'h40e12a4c} /* (31, 24, 5) {real, imag} */,
  {32'hbf2c3f15, 32'h41130e00} /* (31, 24, 4) {real, imag} */,
  {32'h3ff37078, 32'h41306de2} /* (31, 24, 3) {real, imag} */,
  {32'h404693f6, 32'h410f8a3e} /* (31, 24, 2) {real, imag} */,
  {32'h3e4bb654, 32'h40d71c0d} /* (31, 24, 1) {real, imag} */,
  {32'hbff3ae2c, 32'h405576da} /* (31, 24, 0) {real, imag} */,
  {32'hbec471f2, 32'h403bbac5} /* (31, 23, 31) {real, imag} */,
  {32'hbf147dcc, 32'h40f6b335} /* (31, 23, 30) {real, imag} */,
  {32'hbfc8a022, 32'h4101e6f4} /* (31, 23, 29) {real, imag} */,
  {32'h3d493200, 32'h41079497} /* (31, 23, 28) {real, imag} */,
  {32'h3facf260, 32'h40c46d18} /* (31, 23, 27) {real, imag} */,
  {32'h3ff54f94, 32'h40b26ead} /* (31, 23, 26) {real, imag} */,
  {32'h3f9df6cf, 32'h40e431c6} /* (31, 23, 25) {real, imag} */,
  {32'h3fe33bf2, 32'h40f3fadc} /* (31, 23, 24) {real, imag} */,
  {32'h40b8ab12, 32'h4126443e} /* (31, 23, 23) {real, imag} */,
  {32'h409d96bf, 32'h410d42c5} /* (31, 23, 22) {real, imag} */,
  {32'h40811e26, 32'h4056f11d} /* (31, 23, 21) {real, imag} */,
  {32'h3fc62e26, 32'hc1011642} /* (31, 23, 20) {real, imag} */,
  {32'hbfb8f2cc, 32'hc10fedd0} /* (31, 23, 19) {real, imag} */,
  {32'hbf17f75e, 32'hc0c6bf84} /* (31, 23, 18) {real, imag} */,
  {32'h3ff67d20, 32'hc0ec893e} /* (31, 23, 17) {real, imag} */,
  {32'hbf949112, 32'hc0f5b4c8} /* (31, 23, 16) {real, imag} */,
  {32'hbfbdd10a, 32'hc0f2f51d} /* (31, 23, 15) {real, imag} */,
  {32'hbf83f461, 32'hc0fc531c} /* (31, 23, 14) {real, imag} */,
  {32'h3f9d0328, 32'hc1150166} /* (31, 23, 13) {real, imag} */,
  {32'h3f9eb3db, 32'hc1111d97} /* (31, 23, 12) {real, imag} */,
  {32'h40886c1c, 32'hc08d00ec} /* (31, 23, 11) {real, imag} */,
  {32'h404e5136, 32'h4060b16e} /* (31, 23, 10) {real, imag} */,
  {32'hbd831ce6, 32'h40cfddd2} /* (31, 23, 9) {real, imag} */,
  {32'h3fc80c4e, 32'h40c8808e} /* (31, 23, 8) {real, imag} */,
  {32'h3ff255ae, 32'h410a3dbb} /* (31, 23, 7) {real, imag} */,
  {32'h401a8308, 32'h411c2082} /* (31, 23, 6) {real, imag} */,
  {32'h3f019c4e, 32'h4133358a} /* (31, 23, 5) {real, imag} */,
  {32'h3f2a80b3, 32'h4130d0ce} /* (31, 23, 4) {real, imag} */,
  {32'h4019bbc0, 32'h41017669} /* (31, 23, 3) {real, imag} */,
  {32'h406266e3, 32'h40be9750} /* (31, 23, 2) {real, imag} */,
  {32'h3f1572c3, 32'h40e390cc} /* (31, 23, 1) {real, imag} */,
  {32'h3d32fd78, 32'h40736f1b} /* (31, 23, 0) {real, imag} */,
  {32'hbf6c5cb2, 32'h406b597c} /* (31, 22, 31) {real, imag} */,
  {32'hbfbe93b6, 32'h40ed9135} /* (31, 22, 30) {real, imag} */,
  {32'hbfee9fd0, 32'h411700b4} /* (31, 22, 29) {real, imag} */,
  {32'hc009e994, 32'h411c5ea0} /* (31, 22, 28) {real, imag} */,
  {32'hbfb6b14b, 32'h40fc6490} /* (31, 22, 27) {real, imag} */,
  {32'hbe10791b, 32'h40d61af4} /* (31, 22, 26) {real, imag} */,
  {32'hbe05d6c2, 32'h40d0daa5} /* (31, 22, 25) {real, imag} */,
  {32'hbf18c4d6, 32'h40eb0308} /* (31, 22, 24) {real, imag} */,
  {32'h403113a2, 32'h413c0223} /* (31, 22, 23) {real, imag} */,
  {32'h408fe4cb, 32'h41252c56} /* (31, 22, 22) {real, imag} */,
  {32'h40105a0e, 32'h405362c4} /* (31, 22, 21) {real, imag} */,
  {32'h3f8d2c52, 32'hc0d178aa} /* (31, 22, 20) {real, imag} */,
  {32'hbdc26ad4, 32'hc11fec44} /* (31, 22, 19) {real, imag} */,
  {32'h3f124189, 32'hc1237056} /* (31, 22, 18) {real, imag} */,
  {32'h3ec0b9a3, 32'hc102fe6e} /* (31, 22, 17) {real, imag} */,
  {32'hbfd32efe, 32'hc1052ca9} /* (31, 22, 16) {real, imag} */,
  {32'hc02522f8, 32'hc0ead6ac} /* (31, 22, 15) {real, imag} */,
  {32'hbf233b02, 32'hc11222c0} /* (31, 22, 14) {real, imag} */,
  {32'h3f4da032, 32'hc12f7e86} /* (31, 22, 13) {real, imag} */,
  {32'h3fe47fde, 32'hc15383fd} /* (31, 22, 12) {real, imag} */,
  {32'h402b081f, 32'hc113c8f2} /* (31, 22, 11) {real, imag} */,
  {32'h40105e8e, 32'h40131490} /* (31, 22, 10) {real, imag} */,
  {32'hbea4caa8, 32'h4103da72} /* (31, 22, 9) {real, imag} */,
  {32'hbe940136, 32'h4101c844} /* (31, 22, 8) {real, imag} */,
  {32'h400ce6f2, 32'h410f25e5} /* (31, 22, 7) {real, imag} */,
  {32'h3fd8e1e6, 32'h4100ca11} /* (31, 22, 6) {real, imag} */,
  {32'hbee49a24, 32'h410cced8} /* (31, 22, 5) {real, imag} */,
  {32'h4037cbc7, 32'h40d49660} /* (31, 22, 4) {real, imag} */,
  {32'h406879cc, 32'h40cfb8a4} /* (31, 22, 3) {real, imag} */,
  {32'h3fe71258, 32'h40de7304} /* (31, 22, 2) {real, imag} */,
  {32'h403e8ae0, 32'h40f68604} /* (31, 22, 1) {real, imag} */,
  {32'h3fc39e77, 32'h4078ced0} /* (31, 22, 0) {real, imag} */,
  {32'hbf7c4bd1, 32'h40189a02} /* (31, 21, 31) {real, imag} */,
  {32'h3fe9cd3b, 32'h40bb32a6} /* (31, 21, 30) {real, imag} */,
  {32'h4036796c, 32'h40c98723} /* (31, 21, 29) {real, imag} */,
  {32'hbf0b57ee, 32'h40de8062} /* (31, 21, 28) {real, imag} */,
  {32'h3def6460, 32'h40a49d54} /* (31, 21, 27) {real, imag} */,
  {32'h3fd630ca, 32'h401d3d96} /* (31, 21, 26) {real, imag} */,
  {32'h40048cc1, 32'h40ac2ac2} /* (31, 21, 25) {real, imag} */,
  {32'hbf597418, 32'h408885c4} /* (31, 21, 24) {real, imag} */,
  {32'hbe9c2c22, 32'h408075ec} /* (31, 21, 23) {real, imag} */,
  {32'hbfe15c09, 32'h40713c00} /* (31, 21, 22) {real, imag} */,
  {32'hbfde3f4e, 32'h400377e6} /* (31, 21, 21) {real, imag} */,
  {32'h3ee7a064, 32'hc0050ec0} /* (31, 21, 20) {real, imag} */,
  {32'h3e76fed1, 32'hc08ab9e4} /* (31, 21, 19) {real, imag} */,
  {32'h3fdcf0a8, 32'hc0aed4dc} /* (31, 21, 18) {real, imag} */,
  {32'h3d98c6dc, 32'hc08644de} /* (31, 21, 17) {real, imag} */,
  {32'hbf95bc5a, 32'hc002f5d7} /* (31, 21, 16) {real, imag} */,
  {32'hc07f9749, 32'hc000c370} /* (31, 21, 15) {real, imag} */,
  {32'hbfcc9002, 32'hc0ab3c8f} /* (31, 21, 14) {real, imag} */,
  {32'h3fad6ef6, 32'hc0e4b98e} /* (31, 21, 13) {real, imag} */,
  {32'hbe7cbbf9, 32'hc0deef85} /* (31, 21, 12) {real, imag} */,
  {32'h3fd8aa5a, 32'hc022c329} /* (31, 21, 11) {real, imag} */,
  {32'h405da10a, 32'h408e0e8e} /* (31, 21, 10) {real, imag} */,
  {32'hbec3376d, 32'h40998e0f} /* (31, 21, 9) {real, imag} */,
  {32'hbfe13e80, 32'h40c1e174} /* (31, 21, 8) {real, imag} */,
  {32'h3f0b2724, 32'h40aace6a} /* (31, 21, 7) {real, imag} */,
  {32'h3f9b0220, 32'h3f525b27} /* (31, 21, 6) {real, imag} */,
  {32'hbf8abd1f, 32'h401d9d17} /* (31, 21, 5) {real, imag} */,
  {32'hbed2fa79, 32'h3ffa6cd0} /* (31, 21, 4) {real, imag} */,
  {32'hbe6e9655, 32'h3fcce369} /* (31, 21, 3) {real, imag} */,
  {32'h3f904190, 32'h405ce936} /* (31, 21, 2) {real, imag} */,
  {32'h3fc491aa, 32'h406ef1c6} /* (31, 21, 1) {real, imag} */,
  {32'hbf3fd7a2, 32'h3f85104c} /* (31, 21, 0) {real, imag} */,
  {32'hbed8ea6c, 32'hc066c033} /* (31, 20, 31) {real, imag} */,
  {32'h3ff4c8bc, 32'hc0d20571} /* (31, 20, 30) {real, imag} */,
  {32'h40886c0a, 32'hc0bd4076} /* (31, 20, 29) {real, imag} */,
  {32'h407861e4, 32'hc03e0628} /* (31, 20, 28) {real, imag} */,
  {32'h3fa76193, 32'hc0a6a2ae} /* (31, 20, 27) {real, imag} */,
  {32'hbd5a4bd8, 32'hc0e47666} /* (31, 20, 26) {real, imag} */,
  {32'h406a6eaa, 32'hc04685e2} /* (31, 20, 25) {real, imag} */,
  {32'hbf84349e, 32'hc08b0e90} /* (31, 20, 24) {real, imag} */,
  {32'hbe468b90, 32'hc10f451c} /* (31, 20, 23) {real, imag} */,
  {32'h3ef9500e, 32'hc113cc44} /* (31, 20, 22) {real, imag} */,
  {32'hbdd276e0, 32'hc07d41a0} /* (31, 20, 21) {real, imag} */,
  {32'hbd7dae18, 32'h4083bd05} /* (31, 20, 20) {real, imag} */,
  {32'hbf89045e, 32'h40c56495} /* (31, 20, 19) {real, imag} */,
  {32'h3e11b292, 32'h409ceb59} /* (31, 20, 18) {real, imag} */,
  {32'h3e253054, 32'h40feede6} /* (31, 20, 17) {real, imag} */,
  {32'hbe2f243e, 32'h40f199a2} /* (31, 20, 16) {real, imag} */,
  {32'hc0403cc8, 32'h40c78932} /* (31, 20, 15) {real, imag} */,
  {32'hbfe32829, 32'h40938362} /* (31, 20, 14) {real, imag} */,
  {32'h403f2aed, 32'h409919b5} /* (31, 20, 13) {real, imag} */,
  {32'h3f53d00d, 32'h40b78a2a} /* (31, 20, 12) {real, imag} */,
  {32'h3fbd33c8, 32'h40e99769} /* (31, 20, 11) {real, imag} */,
  {32'h40383e6c, 32'hbe527498} /* (31, 20, 10) {real, imag} */,
  {32'hbfcb085c, 32'hc0d769b6} /* (31, 20, 9) {real, imag} */,
  {32'hc085760d, 32'hc0d0e030} /* (31, 20, 8) {real, imag} */,
  {32'hbf3afd98, 32'hc0ba4b7a} /* (31, 20, 7) {real, imag} */,
  {32'hbf8a2605, 32'hc0de58f8} /* (31, 20, 6) {real, imag} */,
  {32'hbefa2e36, 32'hc073e354} /* (31, 20, 5) {real, imag} */,
  {32'hc00f44b8, 32'hc0c8a28c} /* (31, 20, 4) {real, imag} */,
  {32'hc06b81ee, 32'hc0f2d848} /* (31, 20, 3) {real, imag} */,
  {32'hbefd424e, 32'hc09afaac} /* (31, 20, 2) {real, imag} */,
  {32'h3f5cb598, 32'hc0d70775} /* (31, 20, 1) {real, imag} */,
  {32'hbef3cbc8, 32'hc096a236} /* (31, 20, 0) {real, imag} */,
  {32'hbc9630d0, 32'hc07bb8d5} /* (31, 19, 31) {real, imag} */,
  {32'h3fe37603, 32'hc1056942} /* (31, 19, 30) {real, imag} */,
  {32'h3f4c7f9b, 32'hc10c3afc} /* (31, 19, 29) {real, imag} */,
  {32'h3f205430, 32'hc0dcca6c} /* (31, 19, 28) {real, imag} */,
  {32'h3f5e1696, 32'hc1049d56} /* (31, 19, 27) {real, imag} */,
  {32'h3da60492, 32'hc11b5dde} /* (31, 19, 26) {real, imag} */,
  {32'h3f378110, 32'hc0eb990b} /* (31, 19, 25) {real, imag} */,
  {32'hc01e067a, 32'hc10ccb1c} /* (31, 19, 24) {real, imag} */,
  {32'hc05eeb97, 32'hc136d108} /* (31, 19, 23) {real, imag} */,
  {32'hbf9966bc, 32'hc13269a9} /* (31, 19, 22) {real, imag} */,
  {32'hbf47a643, 32'hc0ae22b4} /* (31, 19, 21) {real, imag} */,
  {32'hbe4c2715, 32'h40c0486b} /* (31, 19, 20) {real, imag} */,
  {32'h3f8349da, 32'h40f856de} /* (31, 19, 19) {real, imag} */,
  {32'h3eeb1b06, 32'h40ece5dc} /* (31, 19, 18) {real, imag} */,
  {32'h3e09bc06, 32'h41103b0c} /* (31, 19, 17) {real, imag} */,
  {32'h3fa45ca1, 32'h411986dc} /* (31, 19, 16) {real, imag} */,
  {32'h3f8b2704, 32'h4112a94b} /* (31, 19, 15) {real, imag} */,
  {32'h3fabc60f, 32'h410e1498} /* (31, 19, 14) {real, imag} */,
  {32'h403a4484, 32'h410e77a2} /* (31, 19, 13) {real, imag} */,
  {32'h3ed7a569, 32'h410ef5bc} /* (31, 19, 12) {real, imag} */,
  {32'h3fdad3c3, 32'h40b0b13e} /* (31, 19, 11) {real, imag} */,
  {32'h4054c45e, 32'hc0704152} /* (31, 19, 10) {real, imag} */,
  {32'hc00c6e47, 32'hc0fd2a72} /* (31, 19, 9) {real, imag} */,
  {32'hc0937f48, 32'hc1022e58} /* (31, 19, 8) {real, imag} */,
  {32'h3fc572c2, 32'hc0f0e1a0} /* (31, 19, 7) {real, imag} */,
  {32'hbeb39ba6, 32'hc0de984f} /* (31, 19, 6) {real, imag} */,
  {32'hbea370c8, 32'hc0a76244} /* (31, 19, 5) {real, imag} */,
  {32'hbf2b83ce, 32'hc0dce896} /* (31, 19, 4) {real, imag} */,
  {32'hbfe6ecbe, 32'hc0e06f20} /* (31, 19, 3) {real, imag} */,
  {32'hc08ec1f2, 32'hc0fce337} /* (31, 19, 2) {real, imag} */,
  {32'hc07f57f8, 32'hc109dcd8} /* (31, 19, 1) {real, imag} */,
  {32'hc01b893c, 32'hc096076c} /* (31, 19, 0) {real, imag} */,
  {32'hc02e05aa, 32'hc0d7d3ec} /* (31, 18, 31) {real, imag} */,
  {32'hbfc7771e, 32'hc12e4310} /* (31, 18, 30) {real, imag} */,
  {32'hbfcfc400, 32'hc10eab25} /* (31, 18, 29) {real, imag} */,
  {32'hbf2d763a, 32'hc0ef3e53} /* (31, 18, 28) {real, imag} */,
  {32'hbfb23210, 32'hc0f24569} /* (31, 18, 27) {real, imag} */,
  {32'h3ed55cc6, 32'hc0bdb049} /* (31, 18, 26) {real, imag} */,
  {32'hbfff5f19, 32'hc1045102} /* (31, 18, 25) {real, imag} */,
  {32'hc05da901, 32'hc142c301} /* (31, 18, 24) {real, imag} */,
  {32'hc0493b3a, 32'hc11a03d0} /* (31, 18, 23) {real, imag} */,
  {32'hbf1c67e2, 32'hc0bce0bb} /* (31, 18, 22) {real, imag} */,
  {32'hbfd8c593, 32'hc0477bb8} /* (31, 18, 21) {real, imag} */,
  {32'hbf90236e, 32'h40df4f71} /* (31, 18, 20) {real, imag} */,
  {32'h400e0674, 32'h410d33e7} /* (31, 18, 19) {real, imag} */,
  {32'h404a4b4c, 32'h40f7513e} /* (31, 18, 18) {real, imag} */,
  {32'h402b95f7, 32'h410ca71d} /* (31, 18, 17) {real, imag} */,
  {32'h407daee9, 32'h4113aacb} /* (31, 18, 16) {real, imag} */,
  {32'h40588684, 32'h41181e53} /* (31, 18, 15) {real, imag} */,
  {32'h3fda4666, 32'h41098ac7} /* (31, 18, 14) {real, imag} */,
  {32'hbee001f8, 32'h4104bf3b} /* (31, 18, 13) {real, imag} */,
  {32'hbe7d4ccc, 32'h410873a7} /* (31, 18, 12) {real, imag} */,
  {32'hbdbf4df8, 32'h407874e0} /* (31, 18, 11) {real, imag} */,
  {32'hbf5dec64, 32'hc09c5292} /* (31, 18, 10) {real, imag} */,
  {32'hc09c6032, 32'hc0e14d00} /* (31, 18, 9) {real, imag} */,
  {32'hc04da3f3, 32'hc10a0147} /* (31, 18, 8) {real, imag} */,
  {32'h3fc7be50, 32'hc1073c52} /* (31, 18, 7) {real, imag} */,
  {32'h3fd52d02, 32'hc0e56285} /* (31, 18, 6) {real, imag} */,
  {32'h3fb098c0, 32'hc0b5fa17} /* (31, 18, 5) {real, imag} */,
  {32'hbffa2733, 32'hc0bb3274} /* (31, 18, 4) {real, imag} */,
  {32'hbf10115c, 32'hc0da00dc} /* (31, 18, 3) {real, imag} */,
  {32'hc0134c64, 32'hc11133ea} /* (31, 18, 2) {real, imag} */,
  {32'hc09237c4, 32'hc11ef9f2} /* (31, 18, 1) {real, imag} */,
  {32'hc0842470, 32'hc0d73eb0} /* (31, 18, 0) {real, imag} */,
  {32'hc04165c6, 32'hc0a0467a} /* (31, 17, 31) {real, imag} */,
  {32'hc060d77a, 32'hc1088456} /* (31, 17, 30) {real, imag} */,
  {32'hc02bf998, 32'hc1118fb8} /* (31, 17, 29) {real, imag} */,
  {32'hbffc724a, 32'hc11a50f0} /* (31, 17, 28) {real, imag} */,
  {32'hbf42c016, 32'hc111402b} /* (31, 17, 27) {real, imag} */,
  {32'h3f76793a, 32'hc0c13cfd} /* (31, 17, 26) {real, imag} */,
  {32'hbfca35c0, 32'hc106ebaa} /* (31, 17, 25) {real, imag} */,
  {32'hc07d9fd3, 32'hc1560c62} /* (31, 17, 24) {real, imag} */,
  {32'hbf1127e1, 32'hc1360f7a} /* (31, 17, 23) {real, imag} */,
  {32'h3fb59523, 32'hc0f2f5d8} /* (31, 17, 22) {real, imag} */,
  {32'hc027c148, 32'hbf9223f4} /* (31, 17, 21) {real, imag} */,
  {32'hbd2937f8, 32'h40e02cb0} /* (31, 17, 20) {real, imag} */,
  {32'h3fa59d10, 32'h410ed796} /* (31, 17, 19) {real, imag} */,
  {32'h3fbb5b02, 32'h4108b9b1} /* (31, 17, 18) {real, imag} */,
  {32'h3ff522f3, 32'h40d13328} /* (31, 17, 17) {real, imag} */,
  {32'h401c6164, 32'h40e436f7} /* (31, 17, 16) {real, imag} */,
  {32'h401bd18a, 32'h410fc79b} /* (31, 17, 15) {real, imag} */,
  {32'h4081b80a, 32'h41070308} /* (31, 17, 14) {real, imag} */,
  {32'h3f3a66b2, 32'h4109a9d6} /* (31, 17, 13) {real, imag} */,
  {32'h3feedef1, 32'h4126204a} /* (31, 17, 12) {real, imag} */,
  {32'h4014a9d6, 32'h409a7202} /* (31, 17, 11) {real, imag} */,
  {32'h3f5dc6c2, 32'hc08a7cd3} /* (31, 17, 10) {real, imag} */,
  {32'hc0155ab7, 32'hc10b81f2} /* (31, 17, 9) {real, imag} */,
  {32'hc04ebca3, 32'hc10b3a62} /* (31, 17, 8) {real, imag} */,
  {32'h3eb761f2, 32'hc1129218} /* (31, 17, 7) {real, imag} */,
  {32'h4097bc86, 32'hc1274ca6} /* (31, 17, 6) {real, imag} */,
  {32'h401aaf5c, 32'hc107c71e} /* (31, 17, 5) {real, imag} */,
  {32'hbf907c2c, 32'hc106dc6e} /* (31, 17, 4) {real, imag} */,
  {32'hbf417ad5, 32'hc116b366} /* (31, 17, 3) {real, imag} */,
  {32'hc030958c, 32'hc1127ed8} /* (31, 17, 2) {real, imag} */,
  {32'hc065a9b6, 32'hc1143c0c} /* (31, 17, 1) {real, imag} */,
  {32'hbffe9d73, 32'hc0c6f233} /* (31, 17, 0) {real, imag} */,
  {32'hbf7a5aaa, 32'hc0921fdc} /* (31, 16, 31) {real, imag} */,
  {32'hbff52826, 32'hc1270204} /* (31, 16, 30) {real, imag} */,
  {32'hc0409d46, 32'hc113d9e2} /* (31, 16, 29) {real, imag} */,
  {32'hc00f2c4c, 32'hc11ad5be} /* (31, 16, 28) {real, imag} */,
  {32'hbfac1d2f, 32'hc10fe8da} /* (31, 16, 27) {real, imag} */,
  {32'h3d6db3b0, 32'hc0dd3190} /* (31, 16, 26) {real, imag} */,
  {32'hbf78c02e, 32'hc0fe75fe} /* (31, 16, 25) {real, imag} */,
  {32'hc05802f7, 32'hc1293d70} /* (31, 16, 24) {real, imag} */,
  {32'h3f58b67a, 32'hc12b7ec6} /* (31, 16, 23) {real, imag} */,
  {32'h406aad8c, 32'hc1129095} /* (31, 16, 22) {real, imag} */,
  {32'h3edd5f60, 32'h3e93ca03} /* (31, 16, 21) {real, imag} */,
  {32'h4023c096, 32'h4107dafa} /* (31, 16, 20) {real, imag} */,
  {32'h402bdaf6, 32'h4115cd5e} /* (31, 16, 19) {real, imag} */,
  {32'h3f60c905, 32'h4119b166} /* (31, 16, 18) {real, imag} */,
  {32'h3e056dda, 32'h40fb6ccb} /* (31, 16, 17) {real, imag} */,
  {32'hbecef594, 32'h40dfead1} /* (31, 16, 16) {real, imag} */,
  {32'h3fa2878e, 32'h40dd9b53} /* (31, 16, 15) {real, imag} */,
  {32'h403eb18e, 32'h4121c4c8} /* (31, 16, 14) {real, imag} */,
  {32'h40172034, 32'h412c2200} /* (31, 16, 13) {real, imag} */,
  {32'h400d3368, 32'h41146def} /* (31, 16, 12) {real, imag} */,
  {32'h3f0889ac, 32'h40b2d5ad} /* (31, 16, 11) {real, imag} */,
  {32'hbfb556fb, 32'hc04e6c68} /* (31, 16, 10) {real, imag} */,
  {32'hbfadb7ad, 32'hc10c525c} /* (31, 16, 9) {real, imag} */,
  {32'hbfc6b589, 32'hc0d83e4b} /* (31, 16, 8) {real, imag} */,
  {32'h3f8dbefe, 32'hc0f82cce} /* (31, 16, 7) {real, imag} */,
  {32'h3fefbc3b, 32'hc10b4106} /* (31, 16, 6) {real, imag} */,
  {32'hbf1dce0d, 32'hc0df07f2} /* (31, 16, 5) {real, imag} */,
  {32'hc012db1f, 32'hc104d541} /* (31, 16, 4) {real, imag} */,
  {32'hbfda21cf, 32'hc12a455b} /* (31, 16, 3) {real, imag} */,
  {32'hbfe8ac0c, 32'hc128af99} /* (31, 16, 2) {real, imag} */,
  {32'hc031fef1, 32'hc1165ca4} /* (31, 16, 1) {real, imag} */,
  {32'h3ee91d0c, 32'hc087d8d1} /* (31, 16, 0) {real, imag} */,
  {32'hbd19c1b0, 32'hc0890dca} /* (31, 15, 31) {real, imag} */,
  {32'hbfa56b4a, 32'hc11bfe10} /* (31, 15, 30) {real, imag} */,
  {32'hbf957958, 32'hc117d5aa} /* (31, 15, 29) {real, imag} */,
  {32'h3eb9fda3, 32'hc1275287} /* (31, 15, 28) {real, imag} */,
  {32'hbb86f240, 32'hc11bb30a} /* (31, 15, 27) {real, imag} */,
  {32'hbefed505, 32'hc117b846} /* (31, 15, 26) {real, imag} */,
  {32'hbfd9f66c, 32'hc105983e} /* (31, 15, 25) {real, imag} */,
  {32'hbf818f1a, 32'hc111d680} /* (31, 15, 24) {real, imag} */,
  {32'h401c40ad, 32'hc11f98ec} /* (31, 15, 23) {real, imag} */,
  {32'h3eb8ec8f, 32'hc08dd8d0} /* (31, 15, 22) {real, imag} */,
  {32'hbfcaa4a8, 32'h401a12ef} /* (31, 15, 21) {real, imag} */,
  {32'h3fa8eb14, 32'h4117e0bf} /* (31, 15, 20) {real, imag} */,
  {32'h4037f2a8, 32'h411848be} /* (31, 15, 19) {real, imag} */,
  {32'h3fa32266, 32'h411be3b0} /* (31, 15, 18) {real, imag} */,
  {32'h3eb40f39, 32'h412d92f6} /* (31, 15, 17) {real, imag} */,
  {32'h3fc652d4, 32'h412757ec} /* (31, 15, 16) {real, imag} */,
  {32'h400ca3d6, 32'h40d78a16} /* (31, 15, 15) {real, imag} */,
  {32'h3fccb0b6, 32'h40f4397a} /* (31, 15, 14) {real, imag} */,
  {32'h3e645052, 32'h40f79099} /* (31, 15, 13) {real, imag} */,
  {32'h3d7dc440, 32'h4109623e} /* (31, 15, 12) {real, imag} */,
  {32'h3f3be06f, 32'h40e29e0a} /* (31, 15, 11) {real, imag} */,
  {32'hc0443a75, 32'hbf69b30c} /* (31, 15, 10) {real, imag} */,
  {32'hc047ca22, 32'hc0be3c86} /* (31, 15, 9) {real, imag} */,
  {32'hc0350eda, 32'hc0eed412} /* (31, 15, 8) {real, imag} */,
  {32'hc002bccc, 32'hc107e1f7} /* (31, 15, 7) {real, imag} */,
  {32'h3f24d2ab, 32'hc0e165ce} /* (31, 15, 6) {real, imag} */,
  {32'hbfb43ff0, 32'hc093353b} /* (31, 15, 5) {real, imag} */,
  {32'hc041c6c8, 32'hc11a84fc} /* (31, 15, 4) {real, imag} */,
  {32'hc0850986, 32'hc13fa0b4} /* (31, 15, 3) {real, imag} */,
  {32'hbebca06a, 32'hc13a2cc4} /* (31, 15, 2) {real, imag} */,
  {32'h3eecd992, 32'hc12ab2d8} /* (31, 15, 1) {real, imag} */,
  {32'h4008da78, 32'hc0bff4ea} /* (31, 15, 0) {real, imag} */,
  {32'h3f28feae, 32'hc061de68} /* (31, 14, 31) {real, imag} */,
  {32'hbf10f828, 32'hc0eabbc5} /* (31, 14, 30) {real, imag} */,
  {32'hbeb062c6, 32'hc0ee178b} /* (31, 14, 29) {real, imag} */,
  {32'h3fd641c0, 32'hc1103554} /* (31, 14, 28) {real, imag} */,
  {32'h4022f844, 32'hc11738cf} /* (31, 14, 27) {real, imag} */,
  {32'h3f37dd46, 32'hc11aa0f4} /* (31, 14, 26) {real, imag} */,
  {32'hc01a65f6, 32'hc115cd2a} /* (31, 14, 25) {real, imag} */,
  {32'hc08410ba, 32'hc10657b0} /* (31, 14, 24) {real, imag} */,
  {32'hbfdf4b53, 32'hc1223cf4} /* (31, 14, 23) {real, imag} */,
  {32'hc05aed4f, 32'hc0cd0939} /* (31, 14, 22) {real, imag} */,
  {32'hbf4e51a6, 32'hc0108f1b} /* (31, 14, 21) {real, imag} */,
  {32'h3ff6c0dd, 32'h40a9566a} /* (31, 14, 20) {real, imag} */,
  {32'h400e223b, 32'h40b38851} /* (31, 14, 19) {real, imag} */,
  {32'hbef0f788, 32'h40ae98c4} /* (31, 14, 18) {real, imag} */,
  {32'hc041aff3, 32'h40d993bd} /* (31, 14, 17) {real, imag} */,
  {32'h3f299fc0, 32'h40f547ee} /* (31, 14, 16) {real, imag} */,
  {32'h3fdfe74a, 32'h40e74d17} /* (31, 14, 15) {real, imag} */,
  {32'h4003bb65, 32'h40fc7bc9} /* (31, 14, 14) {real, imag} */,
  {32'hbed3bbda, 32'h410c748a} /* (31, 14, 13) {real, imag} */,
  {32'h3f12d1e7, 32'h410b8ef0} /* (31, 14, 12) {real, imag} */,
  {32'h3de40668, 32'h40fcff2c} /* (31, 14, 11) {real, imag} */,
  {32'hbfc3feb3, 32'hbf971177} /* (31, 14, 10) {real, imag} */,
  {32'hc04a731e, 32'hc0dc35cf} /* (31, 14, 9) {real, imag} */,
  {32'hc02d8f33, 32'hc108eb47} /* (31, 14, 8) {real, imag} */,
  {32'hbe15e6f0, 32'hc1267d56} /* (31, 14, 7) {real, imag} */,
  {32'h4005c1e4, 32'hc1042dc8} /* (31, 14, 6) {real, imag} */,
  {32'hbeb40918, 32'hc0ce37f4} /* (31, 14, 5) {real, imag} */,
  {32'hbefc74d8, 32'hc11d2347} /* (31, 14, 4) {real, imag} */,
  {32'hbfaa32b5, 32'hc105ef56} /* (31, 14, 3) {real, imag} */,
  {32'hbcad1260, 32'hc0ff93b4} /* (31, 14, 2) {real, imag} */,
  {32'h40298d1e, 32'hc13adda3} /* (31, 14, 1) {real, imag} */,
  {32'h405292ca, 32'hc0fc16d0} /* (31, 14, 0) {real, imag} */,
  {32'hbf20e0f0, 32'hc0821875} /* (31, 13, 31) {real, imag} */,
  {32'h3f07f2dc, 32'hc108984d} /* (31, 13, 30) {real, imag} */,
  {32'h3f952d84, 32'hc0d588c8} /* (31, 13, 29) {real, imag} */,
  {32'h4000db60, 32'hc117d4b2} /* (31, 13, 28) {real, imag} */,
  {32'h3fca6a8a, 32'hc11ddd7a} /* (31, 13, 27) {real, imag} */,
  {32'hbebb15f8, 32'hc0cd96a6} /* (31, 13, 26) {real, imag} */,
  {32'hbfac1539, 32'hc0bf48a5} /* (31, 13, 25) {real, imag} */,
  {32'hc0147e7e, 32'hc10be176} /* (31, 13, 24) {real, imag} */,
  {32'hbed43dfd, 32'hc131faee} /* (31, 13, 23) {real, imag} */,
  {32'hbe542db4, 32'hc116dde6} /* (31, 13, 22) {real, imag} */,
  {32'hbf15e04a, 32'hc05cfb9f} /* (31, 13, 21) {real, imag} */,
  {32'hbe8b2d31, 32'h409273e5} /* (31, 13, 20) {real, imag} */,
  {32'hbe9e2841, 32'h40df469a} /* (31, 13, 19) {real, imag} */,
  {32'hbfc3a9a0, 32'h40b3318c} /* (31, 13, 18) {real, imag} */,
  {32'hbfd6f9e6, 32'h40b331a8} /* (31, 13, 17) {real, imag} */,
  {32'hbf4d8127, 32'h40d97f05} /* (31, 13, 16) {real, imag} */,
  {32'h3fe62839, 32'h40ffab5b} /* (31, 13, 15) {real, imag} */,
  {32'h400d7a6d, 32'h40d916be} /* (31, 13, 14) {real, imag} */,
  {32'h40154680, 32'h4105298b} /* (31, 13, 13) {real, imag} */,
  {32'h3f3f9810, 32'h410b659c} /* (31, 13, 12) {real, imag} */,
  {32'hbf8b6178, 32'h40fe9376} /* (31, 13, 11) {real, imag} */,
  {32'hc01aba80, 32'hc07f618f} /* (31, 13, 10) {real, imag} */,
  {32'hc0b6b01a, 32'hc12c065b} /* (31, 13, 9) {real, imag} */,
  {32'hc0cae482, 32'hc10c086c} /* (31, 13, 8) {real, imag} */,
  {32'hbe814249, 32'hc116fb9c} /* (31, 13, 7) {real, imag} */,
  {32'h3f520e64, 32'hc1206a44} /* (31, 13, 6) {real, imag} */,
  {32'hc004e79f, 32'hc12dd538} /* (31, 13, 5) {real, imag} */,
  {32'hc02f15f2, 32'hc128e182} /* (31, 13, 4) {real, imag} */,
  {32'hc0539854, 32'hc0fadf48} /* (31, 13, 3) {real, imag} */,
  {32'hbf08759e, 32'hc081938a} /* (31, 13, 2) {real, imag} */,
  {32'h3ff495f3, 32'hc0eab581} /* (31, 13, 1) {real, imag} */,
  {32'h3fe6ed38, 32'hc0ba5245} /* (31, 13, 0) {real, imag} */,
  {32'hbf3fe50a, 32'hc09f9b2b} /* (31, 12, 31) {real, imag} */,
  {32'h3fa3f1e2, 32'hc11259cf} /* (31, 12, 30) {real, imag} */,
  {32'h40621f46, 32'hc0eca033} /* (31, 12, 29) {real, imag} */,
  {32'h3fe4b9b4, 32'hc1193717} /* (31, 12, 28) {real, imag} */,
  {32'hc062fdda, 32'hc10aef92} /* (31, 12, 27) {real, imag} */,
  {32'hc0a49f72, 32'hc0edb72b} /* (31, 12, 26) {real, imag} */,
  {32'hc0021522, 32'hc0c2e610} /* (31, 12, 25) {real, imag} */,
  {32'h3ffdee3a, 32'hc11d279a} /* (31, 12, 24) {real, imag} */,
  {32'h3e87a363, 32'hc12eb661} /* (31, 12, 23) {real, imag} */,
  {32'hc033a2ca, 32'hc1008246} /* (31, 12, 22) {real, imag} */,
  {32'hc03d812c, 32'hc06885c2} /* (31, 12, 21) {real, imag} */,
  {32'hbfdf26b8, 32'h40c4e545} /* (31, 12, 20) {real, imag} */,
  {32'hbdc47dec, 32'h41183002} /* (31, 12, 19) {real, imag} */,
  {32'h3e30a54a, 32'h410630f4} /* (31, 12, 18) {real, imag} */,
  {32'hbdd92cfc, 32'h411ba262} /* (31, 12, 17) {real, imag} */,
  {32'h3dd3a6b4, 32'h411f7072} /* (31, 12, 16) {real, imag} */,
  {32'h403a7d75, 32'h4111a9e0} /* (31, 12, 15) {real, imag} */,
  {32'h408616af, 32'h40d174df} /* (31, 12, 14) {real, imag} */,
  {32'h4072c05e, 32'h40fd651b} /* (31, 12, 13) {real, imag} */,
  {32'h3ed5f730, 32'h4134dc68} /* (31, 12, 12) {real, imag} */,
  {32'hbf81c814, 32'h40d4b932} /* (31, 12, 11) {real, imag} */,
  {32'hbf6ee4f4, 32'hc0efd7de} /* (31, 12, 10) {real, imag} */,
  {32'hc05cf7bb, 32'hc135f8b8} /* (31, 12, 9) {real, imag} */,
  {32'hc094bdd4, 32'hc10ed303} /* (31, 12, 8) {real, imag} */,
  {32'hbf7633db, 32'hc10e799e} /* (31, 12, 7) {real, imag} */,
  {32'hbf1baeef, 32'hc1240bac} /* (31, 12, 6) {real, imag} */,
  {32'hbfa79fc0, 32'hc11b9be8} /* (31, 12, 5) {real, imag} */,
  {32'hbf8d1397, 32'hc0ec5399} /* (31, 12, 4) {real, imag} */,
  {32'hc0069d0e, 32'hc0a187d2} /* (31, 12, 3) {real, imag} */,
  {32'hbfc67b62, 32'hc05f943c} /* (31, 12, 2) {real, imag} */,
  {32'hbf163cf4, 32'hc0500ec0} /* (31, 12, 1) {real, imag} */,
  {32'hbee26648, 32'hc0143ec8} /* (31, 12, 0) {real, imag} */,
  {32'hbf20baa1, 32'hc027db46} /* (31, 11, 31) {real, imag} */,
  {32'hbfc0e177, 32'hc0bc74d6} /* (31, 11, 30) {real, imag} */,
  {32'h3db7341e, 32'hc0951eff} /* (31, 11, 29) {real, imag} */,
  {32'hbebe8073, 32'hc0c7fc07} /* (31, 11, 28) {real, imag} */,
  {32'hbfea5576, 32'hc0d4d02c} /* (31, 11, 27) {real, imag} */,
  {32'hbfda9fde, 32'hc0e19714} /* (31, 11, 26) {real, imag} */,
  {32'hc005d541, 32'hc0cd2d56} /* (31, 11, 25) {real, imag} */,
  {32'h3fc10c3b, 32'hc126fbbc} /* (31, 11, 24) {real, imag} */,
  {32'h4002fcf8, 32'hc10cee31} /* (31, 11, 23) {real, imag} */,
  {32'hc04c228b, 32'hc0cb10c4} /* (31, 11, 22) {real, imag} */,
  {32'hc0169eaa, 32'hbfc384ee} /* (31, 11, 21) {real, imag} */,
  {32'hbe29b734, 32'h40a13f68} /* (31, 11, 20) {real, imag} */,
  {32'h3e2fbe7c, 32'h40a3d17c} /* (31, 11, 19) {real, imag} */,
  {32'hbdeb72f8, 32'h406a36ab} /* (31, 11, 18) {real, imag} */,
  {32'hbe4e2150, 32'h40a3f6dc} /* (31, 11, 17) {real, imag} */,
  {32'h3ec7fbac, 32'h40c358cc} /* (31, 11, 16) {real, imag} */,
  {32'h3f2983e0, 32'h40992c89} /* (31, 11, 15) {real, imag} */,
  {32'h3fb78725, 32'h409e1e6d} /* (31, 11, 14) {real, imag} */,
  {32'hbe063a0c, 32'h40af94b9} /* (31, 11, 13) {real, imag} */,
  {32'hc02e197a, 32'h40fd8164} /* (31, 11, 12) {real, imag} */,
  {32'hc07edc3f, 32'h40a62986} /* (31, 11, 11) {real, imag} */,
  {32'hbfaedca6, 32'hc076f4e9} /* (31, 11, 10) {real, imag} */,
  {32'hbfa75016, 32'hc0d275df} /* (31, 11, 9) {real, imag} */,
  {32'hbf663456, 32'hc10863da} /* (31, 11, 8) {real, imag} */,
  {32'h3fb5c943, 32'hc112fb07} /* (31, 11, 7) {real, imag} */,
  {32'hbf1a50ea, 32'hc1111db4} /* (31, 11, 6) {real, imag} */,
  {32'hc03d2eba, 32'hc0c3a51f} /* (31, 11, 5) {real, imag} */,
  {32'h3f9f0ea7, 32'hc0960568} /* (31, 11, 4) {real, imag} */,
  {32'hc01065a4, 32'hc00e7c6b} /* (31, 11, 3) {real, imag} */,
  {32'hc09bc2ca, 32'hc0be0f4d} /* (31, 11, 2) {real, imag} */,
  {32'hc013b5bb, 32'hc09fb3d5} /* (31, 11, 1) {real, imag} */,
  {32'hbf3118e4, 32'hbfdc0b74} /* (31, 11, 0) {real, imag} */,
  {32'h3f843d40, 32'h40069f0e} /* (31, 10, 31) {real, imag} */,
  {32'hbe3d032f, 32'h4084fd73} /* (31, 10, 30) {real, imag} */,
  {32'hc01613f4, 32'h40e67c36} /* (31, 10, 29) {real, imag} */,
  {32'hbfcf2840, 32'h40be9a84} /* (31, 10, 28) {real, imag} */,
  {32'h3feef866, 32'h40ad64e1} /* (31, 10, 27) {real, imag} */,
  {32'h3ef844be, 32'h3feff1dc} /* (31, 10, 26) {real, imag} */,
  {32'h3fc2bbbb, 32'h3fa5d730} /* (31, 10, 25) {real, imag} */,
  {32'h4037e6eb, 32'h3e324d15} /* (31, 10, 24) {real, imag} */,
  {32'h408e39c4, 32'h406f3758} /* (31, 10, 23) {real, imag} */,
  {32'h3e1187ac, 32'h40959077} /* (31, 10, 22) {real, imag} */,
  {32'hbfcee815, 32'h408a685e} /* (31, 10, 21) {real, imag} */,
  {32'hbf5804b3, 32'hbf4316f2} /* (31, 10, 20) {real, imag} */,
  {32'h3f3c6314, 32'hc094a474} /* (31, 10, 19) {real, imag} */,
  {32'h3ea907a6, 32'hc0cb15e5} /* (31, 10, 18) {real, imag} */,
  {32'hc001d244, 32'hc08e8a75} /* (31, 10, 17) {real, imag} */,
  {32'hbf6039f8, 32'hc0f17913} /* (31, 10, 16) {real, imag} */,
  {32'hc06de258, 32'hc0c12574} /* (31, 10, 15) {real, imag} */,
  {32'hc00f7250, 32'hc031eaa6} /* (31, 10, 14) {real, imag} */,
  {32'hbff1f4d7, 32'hc035bfcb} /* (31, 10, 13) {real, imag} */,
  {32'hc042b2ec, 32'hc05699fa} /* (31, 10, 12) {real, imag} */,
  {32'hbe499ef2, 32'hc02aa641} /* (31, 10, 11) {real, imag} */,
  {32'h3fa0e8fa, 32'hbf413653} /* (31, 10, 10) {real, imag} */,
  {32'h4002db33, 32'h401cfb4c} /* (31, 10, 9) {real, imag} */,
  {32'h3f286e0d, 32'h3faaeef5} /* (31, 10, 8) {real, imag} */,
  {32'h3fef621c, 32'h3fbf19fe} /* (31, 10, 7) {real, imag} */,
  {32'h3ffbeb9e, 32'h40137c6c} /* (31, 10, 6) {real, imag} */,
  {32'hbeb14d5c, 32'h409e82d6} /* (31, 10, 5) {real, imag} */,
  {32'h40217930, 32'h409dc264} /* (31, 10, 4) {real, imag} */,
  {32'hbfb96968, 32'h40c26433} /* (31, 10, 3) {real, imag} */,
  {32'hc03e3f00, 32'h3f400d3a} /* (31, 10, 2) {real, imag} */,
  {32'hc002995c, 32'h40063c94} /* (31, 10, 1) {real, imag} */,
  {32'hbcbd1688, 32'h401c0571} /* (31, 10, 0) {real, imag} */,
  {32'h3fdfc816, 32'h403ce72d} /* (31, 9, 31) {real, imag} */,
  {32'h4050d0f0, 32'h40b4caac} /* (31, 9, 30) {real, imag} */,
  {32'h3fbe5b68, 32'h411293d5} /* (31, 9, 29) {real, imag} */,
  {32'hbf33d006, 32'h4129b5a3} /* (31, 9, 28) {real, imag} */,
  {32'h3fbd2496, 32'h41408898} /* (31, 9, 27) {real, imag} */,
  {32'hbd9c17cc, 32'h410d5694} /* (31, 9, 26) {real, imag} */,
  {32'h3fd3980a, 32'h40f1bf3f} /* (31, 9, 25) {real, imag} */,
  {32'h3fa2cb2c, 32'h4101a3bb} /* (31, 9, 24) {real, imag} */,
  {32'h3fea7170, 32'h410dd6c4} /* (31, 9, 23) {real, imag} */,
  {32'h3fdb4699, 32'h40eeb038} /* (31, 9, 22) {real, imag} */,
  {32'hbf03999a, 32'h40bfef7d} /* (31, 9, 21) {real, imag} */,
  {32'hc0077152, 32'hc03c8507} /* (31, 9, 20) {real, imag} */,
  {32'hbe8f7a25, 32'hc0bea81a} /* (31, 9, 19) {real, imag} */,
  {32'hbf5e1bba, 32'hc11cb8fa} /* (31, 9, 18) {real, imag} */,
  {32'hc0972cc4, 32'hc1120f44} /* (31, 9, 17) {real, imag} */,
  {32'hc08bd0bc, 32'hc1227f9c} /* (31, 9, 16) {real, imag} */,
  {32'hc082e936, 32'hc112c55c} /* (31, 9, 15) {real, imag} */,
  {32'hc02e7350, 32'hc117892b} /* (31, 9, 14) {real, imag} */,
  {32'hbf98745d, 32'hc103e816} /* (31, 9, 13) {real, imag} */,
  {32'h3f43de2d, 32'hc0b8a6c2} /* (31, 9, 12) {real, imag} */,
  {32'h402cf976, 32'hc09a5275} /* (31, 9, 11) {real, imag} */,
  {32'h4001081c, 32'h3fad21f4} /* (31, 9, 10) {real, imag} */,
  {32'h408144f9, 32'h40bab180} /* (31, 9, 9) {real, imag} */,
  {32'h3ff0a9a0, 32'h410db0f2} /* (31, 9, 8) {real, imag} */,
  {32'h402770ad, 32'h412d8f0a} /* (31, 9, 7) {real, imag} */,
  {32'h3ff77dde, 32'h410e7b98} /* (31, 9, 6) {real, imag} */,
  {32'h3fd34f43, 32'h41062826} /* (31, 9, 5) {real, imag} */,
  {32'h404acd6c, 32'h40e69190} /* (31, 9, 4) {real, imag} */,
  {32'hbf1fa756, 32'h41045453} /* (31, 9, 3) {real, imag} */,
  {32'hc008b703, 32'h40be14c8} /* (31, 9, 2) {real, imag} */,
  {32'h3f73b32e, 32'h40eec5d1} /* (31, 9, 1) {real, imag} */,
  {32'h3ffdbf93, 32'h40a34e83} /* (31, 9, 0) {real, imag} */,
  {32'h4027cd70, 32'h4038bf84} /* (31, 8, 31) {real, imag} */,
  {32'h405c52f6, 32'h40aefd8f} /* (31, 8, 30) {real, imag} */,
  {32'h405b55b9, 32'h4119d27e} /* (31, 8, 29) {real, imag} */,
  {32'hbe2daeda, 32'h411887ac} /* (31, 8, 28) {real, imag} */,
  {32'h3f1b811b, 32'h411718e2} /* (31, 8, 27) {real, imag} */,
  {32'h3f84a788, 32'h411150d2} /* (31, 8, 26) {real, imag} */,
  {32'h3f35a4e5, 32'h40f639eb} /* (31, 8, 25) {real, imag} */,
  {32'hc02531ea, 32'h4130ed38} /* (31, 8, 24) {real, imag} */,
  {32'h3d77d3d8, 32'h4130ba5b} /* (31, 8, 23) {real, imag} */,
  {32'h3fdb96bd, 32'h410bc3a4} /* (31, 8, 22) {real, imag} */,
  {32'h3f982473, 32'h4095df1f} /* (31, 8, 21) {real, imag} */,
  {32'hbf1bc038, 32'hc08d9e5c} /* (31, 8, 20) {real, imag} */,
  {32'hbf298b52, 32'hc09617bb} /* (31, 8, 19) {real, imag} */,
  {32'hbfa12b4c, 32'hc0be806e} /* (31, 8, 18) {real, imag} */,
  {32'hc0345bec, 32'hc0e9dcf4} /* (31, 8, 17) {real, imag} */,
  {32'hc01f5393, 32'hc1020708} /* (31, 8, 16) {real, imag} */,
  {32'hbf1a0160, 32'hc12386b8} /* (31, 8, 15) {real, imag} */,
  {32'hc08dab9e, 32'hc113baf7} /* (31, 8, 14) {real, imag} */,
  {32'hc097d45d, 32'hc0fce002} /* (31, 8, 13) {real, imag} */,
  {32'hbff9171a, 32'hc0b57cf9} /* (31, 8, 12) {real, imag} */,
  {32'hbfc1dc15, 32'hc0a58d4c} /* (31, 8, 11) {real, imag} */,
  {32'hbfba5338, 32'h3fa65716} /* (31, 8, 10) {real, imag} */,
  {32'h3f350172, 32'h40826c68} /* (31, 8, 9) {real, imag} */,
  {32'hbec8a572, 32'h41119ac8} /* (31, 8, 8) {real, imag} */,
  {32'hbeb152bb, 32'h41335012} /* (31, 8, 7) {real, imag} */,
  {32'hbe78b661, 32'h4112e9d0} /* (31, 8, 6) {real, imag} */,
  {32'h3e98b813, 32'h40ea2b75} /* (31, 8, 5) {real, imag} */,
  {32'h4005d022, 32'h40b5fc8a} /* (31, 8, 4) {real, imag} */,
  {32'h3fc76e66, 32'h40c265c5} /* (31, 8, 3) {real, imag} */,
  {32'h3f6f2e06, 32'h41023619} /* (31, 8, 2) {real, imag} */,
  {32'h403c7b13, 32'h4101336f} /* (31, 8, 1) {real, imag} */,
  {32'h405afba6, 32'h408339b8} /* (31, 8, 0) {real, imag} */,
  {32'h40708508, 32'h40912fd6} /* (31, 7, 31) {real, imag} */,
  {32'h407bd172, 32'h41014d50} /* (31, 7, 30) {real, imag} */,
  {32'h3f74b5d5, 32'h4130b132} /* (31, 7, 29) {real, imag} */,
  {32'hbfd22eed, 32'h410dc78c} /* (31, 7, 28) {real, imag} */,
  {32'hbf3e3fa4, 32'h40dbf53a} /* (31, 7, 27) {real, imag} */,
  {32'hbf2958d6, 32'h40a948de} /* (31, 7, 26) {real, imag} */,
  {32'h404554f8, 32'h40ae2e47} /* (31, 7, 25) {real, imag} */,
  {32'h3e835d62, 32'h4106c0da} /* (31, 7, 24) {real, imag} */,
  {32'h3fc40c41, 32'h412183df} /* (31, 7, 23) {real, imag} */,
  {32'h3f8463e2, 32'h4140a466} /* (31, 7, 22) {real, imag} */,
  {32'h4052ed34, 32'h40cdc551} /* (31, 7, 21) {real, imag} */,
  {32'h4046737f, 32'hc0ac01a3} /* (31, 7, 20) {real, imag} */,
  {32'hbfe0080a, 32'hc0f09e44} /* (31, 7, 19) {real, imag} */,
  {32'hbf9810cf, 32'hc0e12830} /* (31, 7, 18) {real, imag} */,
  {32'hbefa420c, 32'hc0bdd6d2} /* (31, 7, 17) {real, imag} */,
  {32'h3ef70f4d, 32'hc0ff00b0} /* (31, 7, 16) {real, imag} */,
  {32'h3fb1deb0, 32'hc11c1faa} /* (31, 7, 15) {real, imag} */,
  {32'hbee8e36c, 32'hc10eaa6c} /* (31, 7, 14) {real, imag} */,
  {32'hc00caf5c, 32'hc1089bd8} /* (31, 7, 13) {real, imag} */,
  {32'hbf902b00, 32'hc115dccc} /* (31, 7, 12) {real, imag} */,
  {32'hc086abbc, 32'hc0c3ac6c} /* (31, 7, 11) {real, imag} */,
  {32'hbfec6974, 32'h4032def3} /* (31, 7, 10) {real, imag} */,
  {32'h3ff8d2ce, 32'h40cfcc14} /* (31, 7, 9) {real, imag} */,
  {32'h3fc13a96, 32'h4146d839} /* (31, 7, 8) {real, imag} */,
  {32'hbff76513, 32'h412308bd} /* (31, 7, 7) {real, imag} */,
  {32'hbe17a84a, 32'h4107c88a} /* (31, 7, 6) {real, imag} */,
  {32'h3f936704, 32'h410082c6} /* (31, 7, 5) {real, imag} */,
  {32'hbdcd8728, 32'h40f57e3c} /* (31, 7, 4) {real, imag} */,
  {32'h3f192e3e, 32'h40ff0e87} /* (31, 7, 3) {real, imag} */,
  {32'h402b813f, 32'h41225155} /* (31, 7, 2) {real, imag} */,
  {32'h3f8e8706, 32'h410a5a69} /* (31, 7, 1) {real, imag} */,
  {32'h3fbe68c6, 32'h4056ae7a} /* (31, 7, 0) {real, imag} */,
  {32'h4022da9c, 32'h4071531d} /* (31, 6, 31) {real, imag} */,
  {32'h40858d79, 32'h40b30a10} /* (31, 6, 30) {real, imag} */,
  {32'h403cda72, 32'h40a85978} /* (31, 6, 29) {real, imag} */,
  {32'hbfaa41f7, 32'h40fe21d4} /* (31, 6, 28) {real, imag} */,
  {32'hc02f5306, 32'h40e3b088} /* (31, 6, 27) {real, imag} */,
  {32'hbfc92da8, 32'h40ade30a} /* (31, 6, 26) {real, imag} */,
  {32'h4047cfee, 32'h40b2d036} /* (31, 6, 25) {real, imag} */,
  {32'h3fe0ff50, 32'h40fc36c4} /* (31, 6, 24) {real, imag} */,
  {32'h4001fcf9, 32'h410dbc8b} /* (31, 6, 23) {real, imag} */,
  {32'h401cced0, 32'h412156eb} /* (31, 6, 22) {real, imag} */,
  {32'h400c3eb0, 32'h40c09188} /* (31, 6, 21) {real, imag} */,
  {32'h3f01108c, 32'hc0a4cf48} /* (31, 6, 20) {real, imag} */,
  {32'hc0157938, 32'hc0d9989a} /* (31, 6, 19) {real, imag} */,
  {32'hbfbaa637, 32'hc10b42ac} /* (31, 6, 18) {real, imag} */,
  {32'hbf8d2f14, 32'hc0ea42f3} /* (31, 6, 17) {real, imag} */,
  {32'hbf1bdf41, 32'hc10b8f82} /* (31, 6, 16) {real, imag} */,
  {32'hc0321f02, 32'hc12446ae} /* (31, 6, 15) {real, imag} */,
  {32'hbf8fd547, 32'hc118385c} /* (31, 6, 14) {real, imag} */,
  {32'hbff34b9f, 32'hc10c337a} /* (31, 6, 13) {real, imag} */,
  {32'h3f40d9f9, 32'hc12b8bee} /* (31, 6, 12) {real, imag} */,
  {32'hbfb59126, 32'hc0b92f58} /* (31, 6, 11) {real, imag} */,
  {32'h3f7d7424, 32'h4007c224} /* (31, 6, 10) {real, imag} */,
  {32'h404ce793, 32'h409f818e} /* (31, 6, 9) {real, imag} */,
  {32'hbe8dc1c5, 32'h4120a8f8} /* (31, 6, 8) {real, imag} */,
  {32'hbefb9ee4, 32'h40d88214} /* (31, 6, 7) {real, imag} */,
  {32'h3f930089, 32'h410c0fc8} /* (31, 6, 6) {real, imag} */,
  {32'h401346b8, 32'h411b1547} /* (31, 6, 5) {real, imag} */,
  {32'h3fa43282, 32'h4100d77b} /* (31, 6, 4) {real, imag} */,
  {32'h3fe83424, 32'h411389c0} /* (31, 6, 3) {real, imag} */,
  {32'h4040378a, 32'h4115583c} /* (31, 6, 2) {real, imag} */,
  {32'h40000662, 32'h4116bed8} /* (31, 6, 1) {real, imag} */,
  {32'h3f1ff264, 32'h4094184c} /* (31, 6, 0) {real, imag} */,
  {32'h3f8db188, 32'h40b7c7e2} /* (31, 5, 31) {real, imag} */,
  {32'h40050c3c, 32'h40f31b98} /* (31, 5, 30) {real, imag} */,
  {32'h40753cfe, 32'h40e6b6a8} /* (31, 5, 29) {real, imag} */,
  {32'h3f0d2537, 32'h410822e0} /* (31, 5, 28) {real, imag} */,
  {32'hc03f3724, 32'h412583b5} /* (31, 5, 27) {real, imag} */,
  {32'hbf6404a3, 32'h40eb24b6} /* (31, 5, 26) {real, imag} */,
  {32'h3f675e98, 32'h40bd16c9} /* (31, 5, 25) {real, imag} */,
  {32'h3f86e3e8, 32'h40b8f815} /* (31, 5, 24) {real, imag} */,
  {32'h3f787e7e, 32'h41093498} /* (31, 5, 23) {real, imag} */,
  {32'h3fe87647, 32'h41137a34} /* (31, 5, 22) {real, imag} */,
  {32'h40420d02, 32'h40b71014} /* (31, 5, 21) {real, imag} */,
  {32'h3fe6604e, 32'h4014bc2a} /* (31, 5, 20) {real, imag} */,
  {32'h3f90193f, 32'h4024cf2e} /* (31, 5, 19) {real, imag} */,
  {32'hbdcc6988, 32'h40136a7a} /* (31, 5, 18) {real, imag} */,
  {32'hc053aee9, 32'h40384229} /* (31, 5, 17) {real, imag} */,
  {32'hc04c73f4, 32'hbf8c9c87} /* (31, 5, 16) {real, imag} */,
  {32'hc0250978, 32'hc1170d00} /* (31, 5, 15) {real, imag} */,
  {32'hc004a2ba, 32'hc11e14c1} /* (31, 5, 14) {real, imag} */,
  {32'hc01c9d95, 32'hc0b01c80} /* (31, 5, 13) {real, imag} */,
  {32'h4013d11d, 32'hc0eca9bc} /* (31, 5, 12) {real, imag} */,
  {32'hbf8f7a9c, 32'hc1123310} /* (31, 5, 11) {real, imag} */,
  {32'hbf627a67, 32'hc090ffb9} /* (31, 5, 10) {real, imag} */,
  {32'h3f6a5728, 32'hc04e84d5} /* (31, 5, 9) {real, imag} */,
  {32'hbfbd5a0c, 32'hc083561f} /* (31, 5, 8) {real, imag} */,
  {32'hbe100d90, 32'hc056fdc4} /* (31, 5, 7) {real, imag} */,
  {32'hbf9d5b8d, 32'hbec1473c} /* (31, 5, 6) {real, imag} */,
  {32'h401672b5, 32'h40e0e1f4} /* (31, 5, 5) {real, imag} */,
  {32'h406ad54c, 32'h40ed65b0} /* (31, 5, 4) {real, imag} */,
  {32'h403c6bfe, 32'h41290389} /* (31, 5, 3) {real, imag} */,
  {32'h40130c42, 32'h41187565} /* (31, 5, 2) {real, imag} */,
  {32'h3faab43e, 32'h41261c37} /* (31, 5, 1) {real, imag} */,
  {32'h3f686682, 32'h40a4408e} /* (31, 5, 0) {real, imag} */,
  {32'hbf9885d4, 32'h40a65d5c} /* (31, 4, 31) {real, imag} */,
  {32'hbfcd4fe0, 32'h410eb819} /* (31, 4, 30) {real, imag} */,
  {32'hbf47b3ed, 32'h40e45f0e} /* (31, 4, 29) {real, imag} */,
  {32'hbf9c797b, 32'h40ca7cf2} /* (31, 4, 28) {real, imag} */,
  {32'hc02efdb1, 32'h4133e12f} /* (31, 4, 27) {real, imag} */,
  {32'hc0258eae, 32'h410f112c} /* (31, 4, 26) {real, imag} */,
  {32'hc0499fa8, 32'h4101c264} /* (31, 4, 25) {real, imag} */,
  {32'hc0009dda, 32'h41022be2} /* (31, 4, 24) {real, imag} */,
  {32'hbfab6683, 32'h41138249} /* (31, 4, 23) {real, imag} */,
  {32'hc00f2a79, 32'h4127090a} /* (31, 4, 22) {real, imag} */,
  {32'h3f06f58a, 32'h4115de73} /* (31, 4, 21) {real, imag} */,
  {32'h40036d71, 32'h412987a1} /* (31, 4, 20) {real, imag} */,
  {32'h3fd4096a, 32'h411324ca} /* (31, 4, 19) {real, imag} */,
  {32'h3f8b623c, 32'h410f64fe} /* (31, 4, 18) {real, imag} */,
  {32'hbe2f509c, 32'h411c898a} /* (31, 4, 17) {real, imag} */,
  {32'hbfc75118, 32'h408ee8fe} /* (31, 4, 16) {real, imag} */,
  {32'hbe822c00, 32'hc105f316} /* (31, 4, 15) {real, imag} */,
  {32'hc00dd65e, 32'hc0e85edc} /* (31, 4, 14) {real, imag} */,
  {32'hbfa1a482, 32'hc096b1cf} /* (31, 4, 13) {real, imag} */,
  {32'h3e875943, 32'hc0ff5804} /* (31, 4, 12) {real, imag} */,
  {32'hc0218d48, 32'hc113684d} /* (31, 4, 11) {real, imag} */,
  {32'hc02bd995, 32'hc0c97328} /* (31, 4, 10) {real, imag} */,
  {32'hbf1ff08a, 32'hc1049600} /* (31, 4, 9) {real, imag} */,
  {32'hbfd3cb65, 32'hc13d2652} /* (31, 4, 8) {real, imag} */,
  {32'hbf24343d, 32'hc1170ee6} /* (31, 4, 7) {real, imag} */,
  {32'hbf279aae, 32'hc0efb04f} /* (31, 4, 6) {real, imag} */,
  {32'h4071972f, 32'h3f5135b2} /* (31, 4, 5) {real, imag} */,
  {32'h40a1b5ae, 32'h40cd6fe8} /* (31, 4, 4) {real, imag} */,
  {32'h3fbf7a2e, 32'h41071afb} /* (31, 4, 3) {real, imag} */,
  {32'hbe0464aa, 32'h40e5cba6} /* (31, 4, 2) {real, imag} */,
  {32'hbf882409, 32'h410ecf96} /* (31, 4, 1) {real, imag} */,
  {32'h3e8a3045, 32'h40a70a44} /* (31, 4, 0) {real, imag} */,
  {32'hbfb7bf67, 32'h408dbf94} /* (31, 3, 31) {real, imag} */,
  {32'h3fdab86c, 32'h40f87aea} /* (31, 3, 30) {real, imag} */,
  {32'h3cfa8e10, 32'h40fa002d} /* (31, 3, 29) {real, imag} */,
  {32'hc00af643, 32'h40e940a2} /* (31, 3, 28) {real, imag} */,
  {32'hbead4cc9, 32'h4108d6f8} /* (31, 3, 27) {real, imag} */,
  {32'h3eaf6e02, 32'h40da27de} /* (31, 3, 26) {real, imag} */,
  {32'hbf82af02, 32'h411694d8} /* (31, 3, 25) {real, imag} */,
  {32'hc03c64ee, 32'h4146cc10} /* (31, 3, 24) {real, imag} */,
  {32'hbf90dd96, 32'h41253761} /* (31, 3, 23) {real, imag} */,
  {32'h3e92a0dc, 32'h411f129a} /* (31, 3, 22) {real, imag} */,
  {32'h3fb2bc49, 32'h411c0a3a} /* (31, 3, 21) {real, imag} */,
  {32'h3fb1d09a, 32'h410ff323} /* (31, 3, 20) {real, imag} */,
  {32'h3b3b3c00, 32'h40ebb832} /* (31, 3, 19) {real, imag} */,
  {32'h3f709766, 32'h40e7f70a} /* (31, 3, 18) {real, imag} */,
  {32'h3ffee701, 32'h40fb44f4} /* (31, 3, 17) {real, imag} */,
  {32'hbfa030ab, 32'h406ec0d4} /* (31, 3, 16) {real, imag} */,
  {32'hbf51425e, 32'hc0e08a05} /* (31, 3, 15) {real, imag} */,
  {32'hbff78a00, 32'hc1086eb8} /* (31, 3, 14) {real, imag} */,
  {32'hbf9c8e1d, 32'hc1078a48} /* (31, 3, 13) {real, imag} */,
  {32'hc015e8b0, 32'hc11fcdc0} /* (31, 3, 12) {real, imag} */,
  {32'hbf87dfe7, 32'hc128ab93} /* (31, 3, 11) {real, imag} */,
  {32'hbff15dfa, 32'hc0d76f1d} /* (31, 3, 10) {real, imag} */,
  {32'hc0159a3f, 32'hc10c2102} /* (31, 3, 9) {real, imag} */,
  {32'hc02a3af4, 32'hc142e808} /* (31, 3, 8) {real, imag} */,
  {32'hc02e094e, 32'hc16ccb7a} /* (31, 3, 7) {real, imag} */,
  {32'hc01c3205, 32'hc12fb5b8} /* (31, 3, 6) {real, imag} */,
  {32'hbff0c5e0, 32'h3ff32004} /* (31, 3, 5) {real, imag} */,
  {32'hbf4e47b3, 32'h41310fda} /* (31, 3, 4) {real, imag} */,
  {32'hbf6ffa00, 32'h40fe504c} /* (31, 3, 3) {real, imag} */,
  {32'h402a3362, 32'h40f366ce} /* (31, 3, 2) {real, imag} */,
  {32'h3ff67885, 32'h411bacd5} /* (31, 3, 1) {real, imag} */,
  {32'hbd85e9c4, 32'h40c5bf04} /* (31, 3, 0) {real, imag} */,
  {32'hbeb84a55, 32'h40600214} /* (31, 2, 31) {real, imag} */,
  {32'h401842e7, 32'h40ded0a8} /* (31, 2, 30) {real, imag} */,
  {32'h3e2833b8, 32'h410bd75f} /* (31, 2, 29) {real, imag} */,
  {32'hc033876e, 32'h410f4b8e} /* (31, 2, 28) {real, imag} */,
  {32'h3d1e25a8, 32'h40f986ca} /* (31, 2, 27) {real, imag} */,
  {32'h3fda5011, 32'h40cd1912} /* (31, 2, 26) {real, imag} */,
  {32'hbc6422a0, 32'h4115f4b4} /* (31, 2, 25) {real, imag} */,
  {32'h3e63c7f8, 32'h4139c046} /* (31, 2, 24) {real, imag} */,
  {32'h3fc2db00, 32'h4131d8a7} /* (31, 2, 23) {real, imag} */,
  {32'h407cbfe9, 32'h410b46e6} /* (31, 2, 22) {real, imag} */,
  {32'h401bbd52, 32'h40d572be} /* (31, 2, 21) {real, imag} */,
  {32'hbf28974a, 32'h40e75a1f} /* (31, 2, 20) {real, imag} */,
  {32'hbeebe65a, 32'h4121b5a0} /* (31, 2, 19) {real, imag} */,
  {32'h400628c1, 32'h412c440a} /* (31, 2, 18) {real, imag} */,
  {32'h401c2ceb, 32'h410aa99a} /* (31, 2, 17) {real, imag} */,
  {32'hbf74836b, 32'h40ca84da} /* (31, 2, 16) {real, imag} */,
  {32'hbee18916, 32'hbffeda6b} /* (31, 2, 15) {real, imag} */,
  {32'h3e8e8ae2, 32'hc0f60b56} /* (31, 2, 14) {real, imag} */,
  {32'h3f11caa8, 32'hc10b4dd7} /* (31, 2, 13) {real, imag} */,
  {32'h3f142b2f, 32'hc0f9967f} /* (31, 2, 12) {real, imag} */,
  {32'h3f4f152f, 32'hc0e78a94} /* (31, 2, 11) {real, imag} */,
  {32'hbfa3d9ec, 32'hc0d4dcca} /* (31, 2, 10) {real, imag} */,
  {32'hbfc9124c, 32'hc0e5f85a} /* (31, 2, 9) {real, imag} */,
  {32'hc0012881, 32'hc1151f37} /* (31, 2, 8) {real, imag} */,
  {32'hbfcdec8a, 32'hc13f1d7c} /* (31, 2, 7) {real, imag} */,
  {32'hbf5d1549, 32'hc1257ca0} /* (31, 2, 6) {real, imag} */,
  {32'hc086fb92, 32'h40328fc8} /* (31, 2, 5) {real, imag} */,
  {32'hc0896375, 32'h41210cd6} /* (31, 2, 4) {real, imag} */,
  {32'hbf3646a1, 32'h41043156} /* (31, 2, 3) {real, imag} */,
  {32'h3fe08413, 32'h4131a6db} /* (31, 2, 2) {real, imag} */,
  {32'h3e8a2987, 32'h41069f5a} /* (31, 2, 1) {real, imag} */,
  {32'hbf7646d3, 32'h404d5ee4} /* (31, 2, 0) {real, imag} */,
  {32'h3e1f8b68, 32'h3fca4872} /* (31, 1, 31) {real, imag} */,
  {32'h3ed4f557, 32'h409446f2} /* (31, 1, 30) {real, imag} */,
  {32'h3f4ece2a, 32'h410f7e00} /* (31, 1, 29) {real, imag} */,
  {32'h3f0b788a, 32'h41397801} /* (31, 1, 28) {real, imag} */,
  {32'h3ed30fc5, 32'h4131c037} /* (31, 1, 27) {real, imag} */,
  {32'h3f03dd47, 32'h41046014} /* (31, 1, 26) {real, imag} */,
  {32'h3fb1ad2f, 32'h40ea3142} /* (31, 1, 25) {real, imag} */,
  {32'h40411f24, 32'h4105c18d} /* (31, 1, 24) {real, imag} */,
  {32'h401bb2b6, 32'h40ed940c} /* (31, 1, 23) {real, imag} */,
  {32'h405bbbf5, 32'h40228dba} /* (31, 1, 22) {real, imag} */,
  {32'h3fdf5cb9, 32'h409e115c} /* (31, 1, 21) {real, imag} */,
  {32'hbe79f0d7, 32'h40de606b} /* (31, 1, 20) {real, imag} */,
  {32'h3f813268, 32'h40ff4e5c} /* (31, 1, 19) {real, imag} */,
  {32'h4082c4b4, 32'h41129040} /* (31, 1, 18) {real, imag} */,
  {32'h40b3154e, 32'h410a6673} /* (31, 1, 17) {real, imag} */,
  {32'h3eeebcc1, 32'h40bf84e2} /* (31, 1, 16) {real, imag} */,
  {32'hbf8f69d1, 32'hc009e19e} /* (31, 1, 15) {real, imag} */,
  {32'h3f63b0a4, 32'hc0ca0202} /* (31, 1, 14) {real, imag} */,
  {32'h40202784, 32'hc0ce2cc9} /* (31, 1, 13) {real, imag} */,
  {32'hbe6d0dac, 32'hc0ed7988} /* (31, 1, 12) {real, imag} */,
  {32'hbf773530, 32'hc0f08e75} /* (31, 1, 11) {real, imag} */,
  {32'h3f318ef8, 32'hc0cbc8fa} /* (31, 1, 10) {real, imag} */,
  {32'h3e84aeb8, 32'hc0d61749} /* (31, 1, 9) {real, imag} */,
  {32'h3e488e20, 32'hc11b58fc} /* (31, 1, 8) {real, imag} */,
  {32'h4066fd9c, 32'hc0fd4aa9} /* (31, 1, 7) {real, imag} */,
  {32'h4059bf28, 32'hc0b7ee34} /* (31, 1, 6) {real, imag} */,
  {32'hc0067c51, 32'h3d68abd0} /* (31, 1, 5) {real, imag} */,
  {32'hbf745343, 32'h4086e9ea} /* (31, 1, 4) {real, imag} */,
  {32'h401e0858, 32'h40e09d4f} /* (31, 1, 3) {real, imag} */,
  {32'h40125fe1, 32'h40dbf98e} /* (31, 1, 2) {real, imag} */,
  {32'hbf2434da, 32'h40babb36} /* (31, 1, 1) {real, imag} */,
  {32'hbeeb5f14, 32'h40041de9} /* (31, 1, 0) {real, imag} */,
  {32'h3f2253fa, 32'h4009cb42} /* (31, 0, 31) {real, imag} */,
  {32'h3e8c7019, 32'h40524b3d} /* (31, 0, 30) {real, imag} */,
  {32'hbef5413c, 32'h4052dc8f} /* (31, 0, 29) {real, imag} */,
  {32'hbf2f94a6, 32'h40befcbc} /* (31, 0, 28) {real, imag} */,
  {32'hbecc3bff, 32'h41241210} /* (31, 0, 27) {real, imag} */,
  {32'h3ead008f, 32'h4107f058} /* (31, 0, 26) {real, imag} */,
  {32'h4008d35f, 32'h4081d6cd} /* (31, 0, 25) {real, imag} */,
  {32'h3f9923f6, 32'h40698ac6} /* (31, 0, 24) {real, imag} */,
  {32'hbfbd361e, 32'h40134fc0} /* (31, 0, 23) {real, imag} */,
  {32'h3f9fa477, 32'h3f24c766} /* (31, 0, 22) {real, imag} */,
  {32'h40289836, 32'h4006b68b} /* (31, 0, 21) {real, imag} */,
  {32'h3ffef21d, 32'h403b2764} /* (31, 0, 20) {real, imag} */,
  {32'h3f4b26fc, 32'h40164ba4} /* (31, 0, 19) {real, imag} */,
  {32'h3f6712d3, 32'h403624eb} /* (31, 0, 18) {real, imag} */,
  {32'h4031c478, 32'h408b793c} /* (31, 0, 17) {real, imag} */,
  {32'hbe439c74, 32'h400c26c5} /* (31, 0, 16) {real, imag} */,
  {32'hbfa5ff47, 32'hc01d95f6} /* (31, 0, 15) {real, imag} */,
  {32'h3f8a8e13, 32'hc08ea482} /* (31, 0, 14) {real, imag} */,
  {32'h3fa7cc36, 32'hc0474116} /* (31, 0, 13) {real, imag} */,
  {32'hc00eb34c, 32'hc08e16da} /* (31, 0, 12) {real, imag} */,
  {32'hc01b622c, 32'hc0b30860} /* (31, 0, 11) {real, imag} */,
  {32'h3f1fb5f8, 32'hc080bf6c} /* (31, 0, 10) {real, imag} */,
  {32'h3e9d2039, 32'hc0971bca} /* (31, 0, 9) {real, imag} */,
  {32'h3e8ee750, 32'hc0c83518} /* (31, 0, 8) {real, imag} */,
  {32'h3fbb5e17, 32'hc04e868e} /* (31, 0, 7) {real, imag} */,
  {32'h401e2ce4, 32'hbec7268f} /* (31, 0, 6) {real, imag} */,
  {32'h3de617a0, 32'h3cd6fd38} /* (31, 0, 5) {real, imag} */,
  {32'hbd3bdd64, 32'h3f9b5364} /* (31, 0, 4) {real, imag} */,
  {32'hbf4821e7, 32'h408ad53b} /* (31, 0, 3) {real, imag} */,
  {32'hbf1584c2, 32'h40590231} /* (31, 0, 2) {real, imag} */,
  {32'h3e00f1b0, 32'h4089d1b8} /* (31, 0, 1) {real, imag} */,
  {32'h3e3903ca, 32'h401235b4} /* (31, 0, 0) {real, imag} */,
  {32'h3d01967e, 32'hc06484f2} /* (30, 31, 31) {real, imag} */,
  {32'h3f571cc3, 32'hc0c5fae4} /* (30, 31, 30) {real, imag} */,
  {32'hbfcc8416, 32'hc0d66968} /* (30, 31, 29) {real, imag} */,
  {32'hc06914d1, 32'hc1002642} /* (30, 31, 28) {real, imag} */,
  {32'hc035e531, 32'hc1232dcb} /* (30, 31, 27) {real, imag} */,
  {32'hbfab88b7, 32'hc130cc3c} /* (30, 31, 26) {real, imag} */,
  {32'hbff75967, 32'hc116bc59} /* (30, 31, 25) {real, imag} */,
  {32'hbfedaf13, 32'hc111b4b6} /* (30, 31, 24) {real, imag} */,
  {32'hc01bc83f, 32'hc0f37ce0} /* (30, 31, 23) {real, imag} */,
  {32'hc01f56fc, 32'hc0fee966} /* (30, 31, 22) {real, imag} */,
  {32'hc00dbc31, 32'hc0668e8a} /* (30, 31, 21) {real, imag} */,
  {32'h3e40eda6, 32'h404ebf0d} /* (30, 31, 20) {real, imag} */,
  {32'h3f0a4e8f, 32'h4096e0a9} /* (30, 31, 19) {real, imag} */,
  {32'hbf85b1b8, 32'h4092b51a} /* (30, 31, 18) {real, imag} */,
  {32'hbf30783a, 32'h409218d5} /* (30, 31, 17) {real, imag} */,
  {32'h3fa5e0a8, 32'h40bfe476} /* (30, 31, 16) {real, imag} */,
  {32'h3fb6a424, 32'h410171d2} /* (30, 31, 15) {real, imag} */,
  {32'h40271418, 32'h41156335} /* (30, 31, 14) {real, imag} */,
  {32'h3fa26cd6, 32'h41380c3f} /* (30, 31, 13) {real, imag} */,
  {32'h3f96b9ce, 32'h4102e7fc} /* (30, 31, 12) {real, imag} */,
  {32'h3fdd53ae, 32'h40c5f0bb} /* (30, 31, 11) {real, imag} */,
  {32'hc0244d94, 32'hbfe2cc68} /* (30, 31, 10) {real, imag} */,
  {32'hbf625198, 32'hc0f997be} /* (30, 31, 9) {real, imag} */,
  {32'hbfdb148c, 32'hc0e5fcc8} /* (30, 31, 8) {real, imag} */,
  {32'hc086896d, 32'hc0bd8844} /* (30, 31, 7) {real, imag} */,
  {32'hbfc4a4ce, 32'hc104697e} /* (30, 31, 6) {real, imag} */,
  {32'hbfb5f2a3, 32'hc1173129} /* (30, 31, 5) {real, imag} */,
  {32'hbfa11c2e, 32'hc1024bf7} /* (30, 31, 4) {real, imag} */,
  {32'hc006f431, 32'hc0ea75a3} /* (30, 31, 3) {real, imag} */,
  {32'hc0119f1d, 32'hc1262d3e} /* (30, 31, 2) {real, imag} */,
  {32'hbfb78eb0, 32'hc0f4f4b9} /* (30, 31, 1) {real, imag} */,
  {32'hbfb3e2eb, 32'hc07c73d8} /* (30, 31, 0) {real, imag} */,
  {32'hbff97500, 32'hc0f2f2b5} /* (30, 30, 31) {real, imag} */,
  {32'hc02cc1c3, 32'hc12f9ede} /* (30, 30, 30) {real, imag} */,
  {32'hc0add34c, 32'hc11cfb2c} /* (30, 30, 29) {real, imag} */,
  {32'hc0eb2d76, 32'hc159af2a} /* (30, 30, 28) {real, imag} */,
  {32'hc0b53924, 32'hc17678fb} /* (30, 30, 27) {real, imag} */,
  {32'hbffcbee2, 32'hc17dcb0b} /* (30, 30, 26) {real, imag} */,
  {32'h3f956ad0, 32'hc18bf9c8} /* (30, 30, 25) {real, imag} */,
  {32'h3f091831, 32'hc1836d46} /* (30, 30, 24) {real, imag} */,
  {32'hbf5dc9e5, 32'hc173635f} /* (30, 30, 23) {real, imag} */,
  {32'hc0383bd8, 32'hc16fac52} /* (30, 30, 22) {real, imag} */,
  {32'hbfe496ab, 32'hc0dcf8da} /* (30, 30, 21) {real, imag} */,
  {32'h4059d509, 32'h40dd545a} /* (30, 30, 20) {real, imag} */,
  {32'h407a7f15, 32'h4130790e} /* (30, 30, 19) {real, imag} */,
  {32'hbf2031c4, 32'h413f5978} /* (30, 30, 18) {real, imag} */,
  {32'h3e51746e, 32'h41472484} /* (30, 30, 17) {real, imag} */,
  {32'h403704b5, 32'h4150356a} /* (30, 30, 16) {real, imag} */,
  {32'h40484edc, 32'h4161a592} /* (30, 30, 15) {real, imag} */,
  {32'h40670428, 32'h41803eee} /* (30, 30, 14) {real, imag} */,
  {32'h3fa0da62, 32'h418af233} /* (30, 30, 13) {real, imag} */,
  {32'h3efd8fea, 32'h417dcbf4} /* (30, 30, 12) {real, imag} */,
  {32'h3f877cf4, 32'h4117c0e8} /* (30, 30, 11) {real, imag} */,
  {32'hc04ffd9d, 32'hc0cad558} /* (30, 30, 10) {real, imag} */,
  {32'hbfca73b4, 32'hc17fc247} /* (30, 30, 9) {real, imag} */,
  {32'hc03be682, 32'hc148d753} /* (30, 30, 8) {real, imag} */,
  {32'hc0d0378c, 32'hc13df1b8} /* (30, 30, 7) {real, imag} */,
  {32'hc03a25f4, 32'hc1784a83} /* (30, 30, 6) {real, imag} */,
  {32'hc02ebc94, 32'hc176ac4c} /* (30, 30, 5) {real, imag} */,
  {32'hc0c4c026, 32'hc185bdf2} /* (30, 30, 4) {real, imag} */,
  {32'hc08ae32b, 32'hc15df9e8} /* (30, 30, 3) {real, imag} */,
  {32'hc0d8f1e8, 32'hc14eeb80} /* (30, 30, 2) {real, imag} */,
  {32'hbf16643d, 32'hc120e0b6} /* (30, 30, 1) {real, imag} */,
  {32'h3f566ce9, 32'hc0b0a7ec} /* (30, 30, 0) {real, imag} */,
  {32'hc08fa42d, 32'hc12704b7} /* (30, 29, 31) {real, imag} */,
  {32'hc08a9e6d, 32'hc1887bfa} /* (30, 29, 30) {real, imag} */,
  {32'hc07fb06b, 32'hc150b0bf} /* (30, 29, 29) {real, imag} */,
  {32'hc08f8282, 32'hc14279fa} /* (30, 29, 28) {real, imag} */,
  {32'hc00b76cc, 32'hc144be26} /* (30, 29, 27) {real, imag} */,
  {32'hbf28eefd, 32'hc15bbc2e} /* (30, 29, 26) {real, imag} */,
  {32'h3fb4a9aa, 32'hc1912eef} /* (30, 29, 25) {real, imag} */,
  {32'hc0398dcb, 32'hc185e91c} /* (30, 29, 24) {real, imag} */,
  {32'hc03ee124, 32'hc18944f8} /* (30, 29, 23) {real, imag} */,
  {32'hc010471b, 32'hc166f80e} /* (30, 29, 22) {real, imag} */,
  {32'hbf015566, 32'hc0763bb8} /* (30, 29, 21) {real, imag} */,
  {32'h40906642, 32'h4147e176} /* (30, 29, 20) {real, imag} */,
  {32'h40759a4c, 32'h4182d0d4} /* (30, 29, 19) {real, imag} */,
  {32'h4017e9a0, 32'h41743d3f} /* (30, 29, 18) {real, imag} */,
  {32'h4025c351, 32'h4182e302} /* (30, 29, 17) {real, imag} */,
  {32'h4058be03, 32'h4189af5e} /* (30, 29, 16) {real, imag} */,
  {32'h408b1f7e, 32'h4174035e} /* (30, 29, 15) {real, imag} */,
  {32'h4066c90a, 32'h416d87ef} /* (30, 29, 14) {real, imag} */,
  {32'h40909910, 32'h416cdc6a} /* (30, 29, 13) {real, imag} */,
  {32'h40756f2a, 32'h417cfc76} /* (30, 29, 12) {real, imag} */,
  {32'h4050d7a4, 32'h41128a2b} /* (30, 29, 11) {real, imag} */,
  {32'hc02eccb9, 32'hc0beb67b} /* (30, 29, 10) {real, imag} */,
  {32'hc0918eb0, 32'hc1662d39} /* (30, 29, 9) {real, imag} */,
  {32'hc099aa87, 32'hc13e4b4a} /* (30, 29, 8) {real, imag} */,
  {32'hc083fbe0, 32'hc138436f} /* (30, 29, 7) {real, imag} */,
  {32'hc0745f33, 32'hc156363c} /* (30, 29, 6) {real, imag} */,
  {32'hc0860080, 32'hc1687ecc} /* (30, 29, 5) {real, imag} */,
  {32'hc109ff19, 32'hc18b6154} /* (30, 29, 4) {real, imag} */,
  {32'hc0e327d4, 32'hc16af390} /* (30, 29, 3) {real, imag} */,
  {32'hc0a120cf, 32'hc130babc} /* (30, 29, 2) {real, imag} */,
  {32'hbf63b60d, 32'hc136758f} /* (30, 29, 1) {real, imag} */,
  {32'hbfb07cd1, 32'hc0ed4158} /* (30, 29, 0) {real, imag} */,
  {32'hc062570a, 32'hc0f60d90} /* (30, 28, 31) {real, imag} */,
  {32'hc02e7abc, 32'hc183801b} /* (30, 28, 30) {real, imag} */,
  {32'hbf7df1c6, 32'hc179a8d8} /* (30, 28, 29) {real, imag} */,
  {32'hc02fe32d, 32'hc16d36ce} /* (30, 28, 28) {real, imag} */,
  {32'hbfa78496, 32'hc17401ad} /* (30, 28, 27) {real, imag} */,
  {32'h3ea5f1a9, 32'hc16f687a} /* (30, 28, 26) {real, imag} */,
  {32'hbf16715e, 32'hc17687e8} /* (30, 28, 25) {real, imag} */,
  {32'hc0ba2ace, 32'hc184789d} /* (30, 28, 24) {real, imag} */,
  {32'hc0ae36c0, 32'hc186c194} /* (30, 28, 23) {real, imag} */,
  {32'hbfd4e9c1, 32'hc16f07ce} /* (30, 28, 22) {real, imag} */,
  {32'h3fb40d97, 32'hc0a6bc74} /* (30, 28, 21) {real, imag} */,
  {32'h40306d4d, 32'h414c80a3} /* (30, 28, 20) {real, imag} */,
  {32'h4012cc22, 32'h418bdbd6} /* (30, 28, 19) {real, imag} */,
  {32'h404bf77e, 32'h416bc2b4} /* (30, 28, 18) {real, imag} */,
  {32'h4058f32e, 32'h4168ae62} /* (30, 28, 17) {real, imag} */,
  {32'h40599de7, 32'h41882094} /* (30, 28, 16) {real, imag} */,
  {32'h409fec38, 32'h41807ed9} /* (30, 28, 15) {real, imag} */,
  {32'h40a35f5e, 32'h414a690b} /* (30, 28, 14) {real, imag} */,
  {32'h40baff0f, 32'h41433171} /* (30, 28, 13) {real, imag} */,
  {32'h40862042, 32'h416e5923} /* (30, 28, 12) {real, imag} */,
  {32'h4024afe2, 32'h413254ac} /* (30, 28, 11) {real, imag} */,
  {32'hbff6cca6, 32'hc06c8f43} /* (30, 28, 10) {real, imag} */,
  {32'hc06385d0, 32'hc178d51a} /* (30, 28, 9) {real, imag} */,
  {32'hbfa7377a, 32'hc180bc54} /* (30, 28, 8) {real, imag} */,
  {32'hc0478616, 32'hc1604f44} /* (30, 28, 7) {real, imag} */,
  {32'hc03dff8c, 32'hc16a1b2c} /* (30, 28, 6) {real, imag} */,
  {32'hc07323b7, 32'hc16d1e73} /* (30, 28, 5) {real, imag} */,
  {32'hc0d6b6ea, 32'hc16cac17} /* (30, 28, 4) {real, imag} */,
  {32'hc0b50d72, 32'hc14389c3} /* (30, 28, 3) {real, imag} */,
  {32'hc08ac776, 32'hc1479271} /* (30, 28, 2) {real, imag} */,
  {32'hc008a0bf, 32'hc14dda9a} /* (30, 28, 1) {real, imag} */,
  {32'hbf986316, 32'hc112f82d} /* (30, 28, 0) {real, imag} */,
  {32'hc04c1ee4, 32'hc0f6dd73} /* (30, 27, 31) {real, imag} */,
  {32'hc01f0f72, 32'hc17f78c6} /* (30, 27, 30) {real, imag} */,
  {32'hc0492120, 32'hc183b549} /* (30, 27, 29) {real, imag} */,
  {32'hc030266c, 32'hc184bcdc} /* (30, 27, 28) {real, imag} */,
  {32'hbe3151c8, 32'hc18ca6e4} /* (30, 27, 27) {real, imag} */,
  {32'h3f1c0601, 32'hc17e9f0c} /* (30, 27, 26) {real, imag} */,
  {32'hbf81189f, 32'hc17f9b12} /* (30, 27, 25) {real, imag} */,
  {32'hc0968457, 32'hc182acd8} /* (30, 27, 24) {real, imag} */,
  {32'hc1055670, 32'hc17ac879} /* (30, 27, 23) {real, imag} */,
  {32'hc03b7457, 32'hc16e2e40} /* (30, 27, 22) {real, imag} */,
  {32'h4038bf7c, 32'hc0e7fc3e} /* (30, 27, 21) {real, imag} */,
  {32'h40adb724, 32'h410cddc8} /* (30, 27, 20) {real, imag} */,
  {32'h4093ace4, 32'h4163c620} /* (30, 27, 19) {real, imag} */,
  {32'h4046d3a5, 32'h416b9b61} /* (30, 27, 18) {real, imag} */,
  {32'h40a8e5b8, 32'h4166ee20} /* (30, 27, 17) {real, imag} */,
  {32'h4088d543, 32'h416020e3} /* (30, 27, 16) {real, imag} */,
  {32'h4089a02b, 32'h41879417} /* (30, 27, 15) {real, imag} */,
  {32'h40a83880, 32'h415eb8a2} /* (30, 27, 14) {real, imag} */,
  {32'h408159af, 32'h413ad5fe} /* (30, 27, 13) {real, imag} */,
  {32'h406caec0, 32'h414d2f4f} /* (30, 27, 12) {real, imag} */,
  {32'h3fdb74d9, 32'h413fb2f6} /* (30, 27, 11) {real, imag} */,
  {32'hbd1873a0, 32'hc0b27098} /* (30, 27, 10) {real, imag} */,
  {32'h3f1552fe, 32'hc1812fdc} /* (30, 27, 9) {real, imag} */,
  {32'hbfb5a81a, 32'hc183682e} /* (30, 27, 8) {real, imag} */,
  {32'hc0a1668d, 32'hc179d131} /* (30, 27, 7) {real, imag} */,
  {32'hc0266652, 32'hc18c6e24} /* (30, 27, 6) {real, imag} */,
  {32'hc082f97c, 32'hc18f7ef6} /* (30, 27, 5) {real, imag} */,
  {32'hc0acfd90, 32'hc171eed2} /* (30, 27, 4) {real, imag} */,
  {32'hbf84d202, 32'hc15f33e4} /* (30, 27, 3) {real, imag} */,
  {32'hc0381f15, 32'hc1696f32} /* (30, 27, 2) {real, imag} */,
  {32'hc09ef037, 32'hc1557ef2} /* (30, 27, 1) {real, imag} */,
  {32'hc02f7741, 32'hc114bc07} /* (30, 27, 0) {real, imag} */,
  {32'hc0597787, 32'hc0d22497} /* (30, 26, 31) {real, imag} */,
  {32'hc0577822, 32'hc14d3ae4} /* (30, 26, 30) {real, imag} */,
  {32'hc042d31a, 32'hc15f004d} /* (30, 26, 29) {real, imag} */,
  {32'hbfd72f06, 32'hc14e9584} /* (30, 26, 28) {real, imag} */,
  {32'h3f413b22, 32'hc158091a} /* (30, 26, 27) {real, imag} */,
  {32'hbf2e56ce, 32'hc1651f9c} /* (30, 26, 26) {real, imag} */,
  {32'hc02d2e70, 32'hc18f994d} /* (30, 26, 25) {real, imag} */,
  {32'hc048e3ee, 32'hc193844f} /* (30, 26, 24) {real, imag} */,
  {32'hc08004a5, 32'hc17cf510} /* (30, 26, 23) {real, imag} */,
  {32'hc0370346, 32'hc15f445a} /* (30, 26, 22) {real, imag} */,
  {32'h3fc9d830, 32'hc0a81412} /* (30, 26, 21) {real, imag} */,
  {32'h4096eb5e, 32'h411c04ce} /* (30, 26, 20) {real, imag} */,
  {32'h40803979, 32'h41482370} /* (30, 26, 19) {real, imag} */,
  {32'h3ec027ca, 32'h415b9c7c} /* (30, 26, 18) {real, imag} */,
  {32'h4056eab4, 32'h416815da} /* (30, 26, 17) {real, imag} */,
  {32'h4048e249, 32'h416a0b57} /* (30, 26, 16) {real, imag} */,
  {32'h404d3e7f, 32'h418c4606} /* (30, 26, 15) {real, imag} */,
  {32'h40a78b48, 32'h417e13b6} /* (30, 26, 14) {real, imag} */,
  {32'h40788fea, 32'h41595f06} /* (30, 26, 13) {real, imag} */,
  {32'h40104e11, 32'h41725806} /* (30, 26, 12) {real, imag} */,
  {32'h4013fd9a, 32'h41274984} /* (30, 26, 11) {real, imag} */,
  {32'h3ebe3786, 32'hc087eda8} /* (30, 26, 10) {real, imag} */,
  {32'hc086f1ab, 32'hc16d2ff0} /* (30, 26, 9) {real, imag} */,
  {32'hc0a95b3a, 32'hc1881d28} /* (30, 26, 8) {real, imag} */,
  {32'hc019d0e2, 32'hc15a7c25} /* (30, 26, 7) {real, imag} */,
  {32'hbf8b5922, 32'hc14ad9c2} /* (30, 26, 6) {real, imag} */,
  {32'hc087d0c0, 32'hc1553276} /* (30, 26, 5) {real, imag} */,
  {32'hc095c716, 32'hc1419e8d} /* (30, 26, 4) {real, imag} */,
  {32'hbf32cd1b, 32'hc15c6620} /* (30, 26, 3) {real, imag} */,
  {32'hc06d9aea, 32'hc17ef46f} /* (30, 26, 2) {real, imag} */,
  {32'hc0c4fc10, 32'hc15818dd} /* (30, 26, 1) {real, imag} */,
  {32'hc059fd4f, 32'hc10c9b3a} /* (30, 26, 0) {real, imag} */,
  {32'hc008c0ca, 32'hc0f945dc} /* (30, 25, 31) {real, imag} */,
  {32'hc0103faf, 32'hc14fcb81} /* (30, 25, 30) {real, imag} */,
  {32'hbffa9420, 32'hc1673317} /* (30, 25, 29) {real, imag} */,
  {32'hc031f468, 32'hc16a0e09} /* (30, 25, 28) {real, imag} */,
  {32'hbf431873, 32'hc17bc2e8} /* (30, 25, 27) {real, imag} */,
  {32'hc00e9591, 32'hc17bb100} /* (30, 25, 26) {real, imag} */,
  {32'hc0156ab6, 32'hc19aab18} /* (30, 25, 25) {real, imag} */,
  {32'hbf99551f, 32'hc187b78e} /* (30, 25, 24) {real, imag} */,
  {32'hbfe2f5fd, 32'hc164064d} /* (30, 25, 23) {real, imag} */,
  {32'hbfe307b1, 32'hc186d0c8} /* (30, 25, 22) {real, imag} */,
  {32'h3d344cb8, 32'hc0fb1c0f} /* (30, 25, 21) {real, imag} */,
  {32'h405db358, 32'h414aab16} /* (30, 25, 20) {real, imag} */,
  {32'h40abc648, 32'h416dda26} /* (30, 25, 19) {real, imag} */,
  {32'h3fbbfe65, 32'h416a55ed} /* (30, 25, 18) {real, imag} */,
  {32'h3fc7af9b, 32'h41787799} /* (30, 25, 17) {real, imag} */,
  {32'h3fe2cccf, 32'h416c4e5a} /* (30, 25, 16) {real, imag} */,
  {32'h405bdc97, 32'h41800671} /* (30, 25, 15) {real, imag} */,
  {32'h3f808440, 32'h418179ee} /* (30, 25, 14) {real, imag} */,
  {32'hbf78214f, 32'h4169c6d2} /* (30, 25, 13) {real, imag} */,
  {32'h4011058e, 32'h41745a83} /* (30, 25, 12) {real, imag} */,
  {32'h40b743fa, 32'h413a6962} /* (30, 25, 11) {real, imag} */,
  {32'h3f8e91a0, 32'hc09b8f27} /* (30, 25, 10) {real, imag} */,
  {32'hc0b62fa0, 32'hc185442c} /* (30, 25, 9) {real, imag} */,
  {32'hc08c087c, 32'hc1a65d98} /* (30, 25, 8) {real, imag} */,
  {32'hc0598fbc, 32'hc16e6062} /* (30, 25, 7) {real, imag} */,
  {32'hc01e9f24, 32'hc14e868a} /* (30, 25, 6) {real, imag} */,
  {32'hc02d8a1a, 32'hc1735ebc} /* (30, 25, 5) {real, imag} */,
  {32'hc050325f, 32'hc1674787} /* (30, 25, 4) {real, imag} */,
  {32'hc01aed4e, 32'hc14f58c6} /* (30, 25, 3) {real, imag} */,
  {32'hc0869e79, 32'hc181abc0} /* (30, 25, 2) {real, imag} */,
  {32'hc0c77a0a, 32'hc14e992a} /* (30, 25, 1) {real, imag} */,
  {32'hc0330ce2, 32'hc0fd2c58} /* (30, 25, 0) {real, imag} */,
  {32'hbff96bc3, 32'hc0c5f43a} /* (30, 24, 31) {real, imag} */,
  {32'hc00e3698, 32'hc13f4091} /* (30, 24, 30) {real, imag} */,
  {32'h3f621614, 32'hc15866ec} /* (30, 24, 29) {real, imag} */,
  {32'hbffaf4dd, 32'hc1601451} /* (30, 24, 28) {real, imag} */,
  {32'hc0a7fdb2, 32'hc176b026} /* (30, 24, 27) {real, imag} */,
  {32'hc0b81b27, 32'hc16bd699} /* (30, 24, 26) {real, imag} */,
  {32'hc0504354, 32'hc17e1b6c} /* (30, 24, 25) {real, imag} */,
  {32'hc0419962, 32'hc1711b77} /* (30, 24, 24) {real, imag} */,
  {32'hc013c6ac, 32'hc160c720} /* (30, 24, 23) {real, imag} */,
  {32'hbf85dcbe, 32'hc174543f} /* (30, 24, 22) {real, imag} */,
  {32'h3f63c68b, 32'hc0b0eb6e} /* (30, 24, 21) {real, imag} */,
  {32'h40d815fe, 32'h416ce95a} /* (30, 24, 20) {real, imag} */,
  {32'h40cab6ba, 32'h41828528} /* (30, 24, 19) {real, imag} */,
  {32'h400ffc6e, 32'h417778f9} /* (30, 24, 18) {real, imag} */,
  {32'h3fb48675, 32'h41734ff8} /* (30, 24, 17) {real, imag} */,
  {32'hbec8c092, 32'h41811c12} /* (30, 24, 16) {real, imag} */,
  {32'h3fd6c809, 32'h4185474e} /* (30, 24, 15) {real, imag} */,
  {32'hbf4587ce, 32'h4183df40} /* (30, 24, 14) {real, imag} */,
  {32'h3f967bdb, 32'h4153994e} /* (30, 24, 13) {real, imag} */,
  {32'h40b7138c, 32'h4172fe7a} /* (30, 24, 12) {real, imag} */,
  {32'h4062733b, 32'h4155b8f2} /* (30, 24, 11) {real, imag} */,
  {32'hc0ae1b33, 32'hc0ce1a20} /* (30, 24, 10) {real, imag} */,
  {32'hc0d84288, 32'hc19c959a} /* (30, 24, 9) {real, imag} */,
  {32'hc040964a, 32'hc1b513a0} /* (30, 24, 8) {real, imag} */,
  {32'hc03d13ec, 32'hc19397ca} /* (30, 24, 7) {real, imag} */,
  {32'hc0339986, 32'hc17699d1} /* (30, 24, 6) {real, imag} */,
  {32'hc00beac7, 32'hc13e3e3c} /* (30, 24, 5) {real, imag} */,
  {32'hc016dbfa, 32'hc1300aa9} /* (30, 24, 4) {real, imag} */,
  {32'hc02cbefe, 32'hc166473f} /* (30, 24, 3) {real, imag} */,
  {32'hc0ae24fe, 32'hc1827d6e} /* (30, 24, 2) {real, imag} */,
  {32'hc0a8f2ac, 32'hc14261c2} /* (30, 24, 1) {real, imag} */,
  {32'hc00a6af2, 32'hc0d2d48e} /* (30, 24, 0) {real, imag} */,
  {32'hbf99b3c2, 32'hc0c5b6e7} /* (30, 23, 31) {real, imag} */,
  {32'hbfcf2aff, 32'hc14f4ecd} /* (30, 23, 30) {real, imag} */,
  {32'hbbdf1680, 32'hc1649f21} /* (30, 23, 29) {real, imag} */,
  {32'hc01c65e3, 32'hc16d10a7} /* (30, 23, 28) {real, imag} */,
  {32'hc0bd678e, 32'hc170a1e8} /* (30, 23, 27) {real, imag} */,
  {32'hc09a6115, 32'hc151c546} /* (30, 23, 26) {real, imag} */,
  {32'hbfdf426b, 32'hc12b6ba2} /* (30, 23, 25) {real, imag} */,
  {32'hc024db88, 32'hc14de7e0} /* (30, 23, 24) {real, imag} */,
  {32'hbfa98bc6, 32'hc181a5d2} /* (30, 23, 23) {real, imag} */,
  {32'hbe33991c, 32'hc176c391} /* (30, 23, 22) {real, imag} */,
  {32'hbf50d3e6, 32'hc0d6eb04} /* (30, 23, 21) {real, imag} */,
  {32'h408d1869, 32'h4154bf02} /* (30, 23, 20) {real, imag} */,
  {32'h4082711f, 32'h418bd736} /* (30, 23, 19) {real, imag} */,
  {32'h3fc8525d, 32'h41929d8b} /* (30, 23, 18) {real, imag} */,
  {32'h3f894077, 32'h4172267c} /* (30, 23, 17) {real, imag} */,
  {32'hbdc07718, 32'h416be15c} /* (30, 23, 16) {real, imag} */,
  {32'hbfa29050, 32'h414b28ef} /* (30, 23, 15) {real, imag} */,
  {32'hbe8e5856, 32'h416be773} /* (30, 23, 14) {real, imag} */,
  {32'h408447e8, 32'h4151091a} /* (30, 23, 13) {real, imag} */,
  {32'h409d1556, 32'h415dd9c0} /* (30, 23, 12) {real, imag} */,
  {32'h406891da, 32'h41415546} /* (30, 23, 11) {real, imag} */,
  {32'hc07228ea, 32'hc0af59be} /* (30, 23, 10) {real, imag} */,
  {32'hc09db60f, 32'hc179ca1a} /* (30, 23, 9) {real, imag} */,
  {32'hc07dc1b6, 32'hc18e0b05} /* (30, 23, 8) {real, imag} */,
  {32'hc031d48e, 32'hc189ffee} /* (30, 23, 7) {real, imag} */,
  {32'hbff50aad, 32'hc15f198d} /* (30, 23, 6) {real, imag} */,
  {32'h3ebace82, 32'hc15048a8} /* (30, 23, 5) {real, imag} */,
  {32'hbef7bfec, 32'hc14d5724} /* (30, 23, 4) {real, imag} */,
  {32'hbff42819, 32'hc181a1ac} /* (30, 23, 3) {real, imag} */,
  {32'hc08c60d6, 32'hc16feaee} /* (30, 23, 2) {real, imag} */,
  {32'hc0291170, 32'hc15e3d20} /* (30, 23, 1) {real, imag} */,
  {32'h3f4c755c, 32'hc0e4e965} /* (30, 23, 0) {real, imag} */,
  {32'hbe664b64, 32'hc1011560} /* (30, 22, 31) {real, imag} */,
  {32'hbedfb97e, 32'hc1881d72} /* (30, 22, 30) {real, imag} */,
  {32'hbf909aa7, 32'hc18b5d39} /* (30, 22, 29) {real, imag} */,
  {32'hc05db881, 32'hc17d350e} /* (30, 22, 28) {real, imag} */,
  {32'hc0c79db0, 32'hc145b610} /* (30, 22, 27) {real, imag} */,
  {32'hc0b5ed42, 32'hc130743c} /* (30, 22, 26) {real, imag} */,
  {32'hc07460d8, 32'hc1086ebe} /* (30, 22, 25) {real, imag} */,
  {32'hbfdc6d6a, 32'hc13f3eac} /* (30, 22, 24) {real, imag} */,
  {32'hbfb204a2, 32'hc180301b} /* (30, 22, 23) {real, imag} */,
  {32'hbf77aba6, 32'hc161b7d2} /* (30, 22, 22) {real, imag} */,
  {32'hc042607a, 32'hc0b549b4} /* (30, 22, 21) {real, imag} */,
  {32'h3fd5d75c, 32'h414ab91f} /* (30, 22, 20) {real, imag} */,
  {32'h3fc2f339, 32'h4181c484} /* (30, 22, 19) {real, imag} */,
  {32'hbf6ba41c, 32'h416e80b2} /* (30, 22, 18) {real, imag} */,
  {32'h3f8664f8, 32'h414e6e33} /* (30, 22, 17) {real, imag} */,
  {32'h3f3263be, 32'h414b334e} /* (30, 22, 16) {real, imag} */,
  {32'h3e6388c8, 32'h4116b692} /* (30, 22, 15) {real, imag} */,
  {32'h4078ed4a, 32'h414c8c9f} /* (30, 22, 14) {real, imag} */,
  {32'h4078ffa8, 32'h416ca544} /* (30, 22, 13) {real, imag} */,
  {32'h3f975a96, 32'h4148b194} /* (30, 22, 12) {real, imag} */,
  {32'h3e6432f8, 32'h411cd6e9} /* (30, 22, 11) {real, imag} */,
  {32'hc050a57a, 32'hc0acaf4a} /* (30, 22, 10) {real, imag} */,
  {32'hc0543203, 32'hc15a7c82} /* (30, 22, 9) {real, imag} */,
  {32'hc0593bc6, 32'hc168eb24} /* (30, 22, 8) {real, imag} */,
  {32'hc030b0f4, 32'hc16ff3de} /* (30, 22, 7) {real, imag} */,
  {32'hc015d188, 32'hc145733c} /* (30, 22, 6) {real, imag} */,
  {32'hbd7b0130, 32'hc14ae50d} /* (30, 22, 5) {real, imag} */,
  {32'h3faf658c, 32'hc1687224} /* (30, 22, 4) {real, imag} */,
  {32'hbffceab1, 32'hc179b170} /* (30, 22, 3) {real, imag} */,
  {32'hc083dbe7, 32'hc18bc943} /* (30, 22, 2) {real, imag} */,
  {32'hc00c3e33, 32'hc192fc22} /* (30, 22, 1) {real, imag} */,
  {32'hbeccc8f5, 32'hc11f83fe} /* (30, 22, 0) {real, imag} */,
  {32'hbf908741, 32'hc084b31c} /* (30, 21, 31) {real, imag} */,
  {32'hbf9f9087, 32'hc0ccf566} /* (30, 21, 30) {real, imag} */,
  {32'hbea55982, 32'hc0d101ae} /* (30, 21, 29) {real, imag} */,
  {32'hc03cf67f, 32'hc0a14d9d} /* (30, 21, 28) {real, imag} */,
  {32'hc0ac3783, 32'hc052459d} /* (30, 21, 27) {real, imag} */,
  {32'hc0952e2f, 32'hc08b7560} /* (30, 21, 26) {real, imag} */,
  {32'hc008434e, 32'hbf15193c} /* (30, 21, 25) {real, imag} */,
  {32'hbf2dc041, 32'hc05cae9e} /* (30, 21, 24) {real, imag} */,
  {32'hbed0d976, 32'hc089e9ec} /* (30, 21, 23) {real, imag} */,
  {32'hbf8fc93e, 32'hc0a19827} /* (30, 21, 22) {real, imag} */,
  {32'hc04741b1, 32'hc0900ad0} /* (30, 21, 21) {real, imag} */,
  {32'h40010dbc, 32'h3fe86169} /* (30, 21, 20) {real, imag} */,
  {32'h402e0886, 32'h40f0c79a} /* (30, 21, 19) {real, imag} */,
  {32'hbf91531c, 32'h4097eeca} /* (30, 21, 18) {real, imag} */,
  {32'hbf62a262, 32'h40729006} /* (30, 21, 17) {real, imag} */,
  {32'hbec3d879, 32'h40833532} /* (30, 21, 16) {real, imag} */,
  {32'h3f8914b4, 32'h4091c06a} /* (30, 21, 15) {real, imag} */,
  {32'hbe1d126c, 32'h40f3c040} /* (30, 21, 14) {real, imag} */,
  {32'hbff18174, 32'h40c6c987} /* (30, 21, 13) {real, imag} */,
  {32'hc0338ab0, 32'h407e1a66} /* (30, 21, 12) {real, imag} */,
  {32'h3f536a0a, 32'h4097ef96} /* (30, 21, 11) {real, imag} */,
  {32'hbf23f6b6, 32'hc01444d2} /* (30, 21, 10) {real, imag} */,
  {32'hbf0f2ed6, 32'hc0dcab18} /* (30, 21, 9) {real, imag} */,
  {32'hbe833504, 32'hc08e9da6} /* (30, 21, 8) {real, imag} */,
  {32'h3f070205, 32'hc09d6582} /* (30, 21, 7) {real, imag} */,
  {32'hbfb19111, 32'hc0824589} /* (30, 21, 6) {real, imag} */,
  {32'hbeb90d37, 32'hc03fecff} /* (30, 21, 5) {real, imag} */,
  {32'h40021654, 32'hc0efd75e} /* (30, 21, 4) {real, imag} */,
  {32'hbfa04006, 32'hc0e046ac} /* (30, 21, 3) {real, imag} */,
  {32'hc0827c18, 32'hc0d70af2} /* (30, 21, 2) {real, imag} */,
  {32'hbfecc51a, 32'hc107c4fb} /* (30, 21, 1) {real, imag} */,
  {32'hbf815597, 32'hc0a475cc} /* (30, 21, 0) {real, imag} */,
  {32'h3e36e7ea, 32'h40ca08e6} /* (30, 20, 31) {real, imag} */,
  {32'h3f8d8ba4, 32'h4150bf8a} /* (30, 20, 30) {real, imag} */,
  {32'hbece3a24, 32'h41436925} /* (30, 20, 29) {real, imag} */,
  {32'hbfa1c225, 32'h416a96a6} /* (30, 20, 28) {real, imag} */,
  {32'hc047e75c, 32'h414debcc} /* (30, 20, 27) {real, imag} */,
  {32'hc0365f14, 32'h41024d8a} /* (30, 20, 26) {real, imag} */,
  {32'h40353848, 32'h416a7aaf} /* (30, 20, 25) {real, imag} */,
  {32'h400a30fc, 32'h417fce40} /* (30, 20, 24) {real, imag} */,
  {32'hbd97b7b0, 32'h41372cd8} /* (30, 20, 23) {real, imag} */,
  {32'h3f3629be, 32'h4127246d} /* (30, 20, 22) {real, imag} */,
  {32'hbfc8a0c4, 32'h4032c8ec} /* (30, 20, 21) {real, imag} */,
  {32'hbf8fed04, 32'hc10b3c12} /* (30, 20, 20) {real, imag} */,
  {32'h3da85340, 32'hc1003e74} /* (30, 20, 19) {real, imag} */,
  {32'hbf9304aa, 32'hc119bbc2} /* (30, 20, 18) {real, imag} */,
  {32'hbe8722da, 32'hc144120c} /* (30, 20, 17) {real, imag} */,
  {32'hbf251f1e, 32'hc13cbd86} /* (30, 20, 16) {real, imag} */,
  {32'hbfb3941f, 32'hc11f38f2} /* (30, 20, 15) {real, imag} */,
  {32'hc0559ec0, 32'hc11599f5} /* (30, 20, 14) {real, imag} */,
  {32'hc0400bc2, 32'hc1432304} /* (30, 20, 13) {real, imag} */,
  {32'hc089fb10, 32'hc144dab2} /* (30, 20, 12) {real, imag} */,
  {32'hbf194392, 32'hc1011956} /* (30, 20, 11) {real, imag} */,
  {32'h3f8f3142, 32'h40a181d7} /* (30, 20, 10) {real, imag} */,
  {32'h3ffb5890, 32'h41044714} /* (30, 20, 9) {real, imag} */,
  {32'h40454258, 32'h41003b87} /* (30, 20, 8) {real, imag} */,
  {32'h402d7ef0, 32'h41262899} /* (30, 20, 7) {real, imag} */,
  {32'h3d99fb08, 32'h414cc296} /* (30, 20, 6) {real, imag} */,
  {32'h3fd3f01c, 32'h4179d006} /* (30, 20, 5) {real, imag} */,
  {32'h3fc2b674, 32'h411f88ba} /* (30, 20, 4) {real, imag} */,
  {32'h400aa68d, 32'h412224e4} /* (30, 20, 3) {real, imag} */,
  {32'h402bc168, 32'h4159d878} /* (30, 20, 2) {real, imag} */,
  {32'h3fd6a2c8, 32'h41160dd2} /* (30, 20, 1) {real, imag} */,
  {32'hbf08c9fc, 32'h4069bdf6} /* (30, 20, 0) {real, imag} */,
  {32'h3f89c3c0, 32'h4101939e} /* (30, 19, 31) {real, imag} */,
  {32'h400e03d8, 32'h41714ef3} /* (30, 19, 30) {real, imag} */,
  {32'h3ffe87fb, 32'h416684e3} /* (30, 19, 29) {real, imag} */,
  {32'h3fa1354c, 32'h418024fc} /* (30, 19, 28) {real, imag} */,
  {32'hbf347415, 32'h4170dcde} /* (30, 19, 27) {real, imag} */,
  {32'h3f492915, 32'h413261fe} /* (30, 19, 26) {real, imag} */,
  {32'h4087cc45, 32'h4153ef83} /* (30, 19, 25) {real, imag} */,
  {32'h40c8bde2, 32'h418965a8} /* (30, 19, 24) {real, imag} */,
  {32'h404f0c54, 32'h416f58b9} /* (30, 19, 23) {real, imag} */,
  {32'h404dd98e, 32'h415fb9ad} /* (30, 19, 22) {real, imag} */,
  {32'h3f5f82ad, 32'h408a0d4e} /* (30, 19, 21) {real, imag} */,
  {32'hc05ddf86, 32'hc14a3092} /* (30, 19, 20) {real, imag} */,
  {32'hc026097c, 32'hc15a799a} /* (30, 19, 19) {real, imag} */,
  {32'hbef65a27, 32'hc14d5e90} /* (30, 19, 18) {real, imag} */,
  {32'hc021fa2f, 32'hc15191c7} /* (30, 19, 17) {real, imag} */,
  {32'hc077508a, 32'hc181d836} /* (30, 19, 16) {real, imag} */,
  {32'hc0a74bba, 32'hc197e2fc} /* (30, 19, 15) {real, imag} */,
  {32'hc08307e0, 32'hc170174e} /* (30, 19, 14) {real, imag} */,
  {32'hbf4f46ad, 32'hc1736589} /* (30, 19, 13) {real, imag} */,
  {32'h3e568d6c, 32'hc17c5194} /* (30, 19, 12) {real, imag} */,
  {32'hbfb0ce62, 32'hc15aeb46} /* (30, 19, 11) {real, imag} */,
  {32'hbdcb70e8, 32'h4073c605} /* (30, 19, 10) {real, imag} */,
  {32'h3fe16f16, 32'h414fba21} /* (30, 19, 9) {real, imag} */,
  {32'h4092e571, 32'h413267da} /* (30, 19, 8) {real, imag} */,
  {32'h3fd9debe, 32'h41693aad} /* (30, 19, 7) {real, imag} */,
  {32'hbfad3ff2, 32'h413d0892} /* (30, 19, 6) {real, imag} */,
  {32'h40372dd4, 32'h4174a9ba} /* (30, 19, 5) {real, imag} */,
  {32'h407e83a6, 32'h4179e1c2} /* (30, 19, 4) {real, imag} */,
  {32'h40a2e9be, 32'h414ace70} /* (30, 19, 3) {real, imag} */,
  {32'h40c20f1e, 32'h41704afd} /* (30, 19, 2) {real, imag} */,
  {32'h40a1dfbe, 32'h4163832c} /* (30, 19, 1) {real, imag} */,
  {32'h400e5635, 32'h4102e9fd} /* (30, 19, 0) {real, imag} */,
  {32'h3fa5a41c, 32'h410501aa} /* (30, 18, 31) {real, imag} */,
  {32'h40814c8c, 32'h4172b0be} /* (30, 18, 30) {real, imag} */,
  {32'h4024b6ae, 32'h416cbab6} /* (30, 18, 29) {real, imag} */,
  {32'h40266029, 32'h41722c34} /* (30, 18, 28) {real, imag} */,
  {32'h407dcd86, 32'h415017c6} /* (30, 18, 27) {real, imag} */,
  {32'h40922adb, 32'h41426b3e} /* (30, 18, 26) {real, imag} */,
  {32'h40a40cb2, 32'h413ee2da} /* (30, 18, 25) {real, imag} */,
  {32'h41190b2c, 32'h416356c6} /* (30, 18, 24) {real, imag} */,
  {32'h40c2fc05, 32'h418047e0} /* (30, 18, 23) {real, imag} */,
  {32'h4005ec80, 32'h416354fa} /* (30, 18, 22) {real, imag} */,
  {32'hbeb018db, 32'h40fadd75} /* (30, 18, 21) {real, imag} */,
  {32'hc073d2ee, 32'hc1013cf8} /* (30, 18, 20) {real, imag} */,
  {32'hbfbfeece, 32'hc152e299} /* (30, 18, 19) {real, imag} */,
  {32'hbdcbdbd8, 32'hc16f3f34} /* (30, 18, 18) {real, imag} */,
  {32'hc09f2374, 32'hc145ce40} /* (30, 18, 17) {real, imag} */,
  {32'hc0b7a824, 32'hc166b24e} /* (30, 18, 16) {real, imag} */,
  {32'hc0aca078, 32'hc17b1dc9} /* (30, 18, 15) {real, imag} */,
  {32'hc0852ae8, 32'hc159a55c} /* (30, 18, 14) {real, imag} */,
  {32'hc062f5e6, 32'hc16cadb4} /* (30, 18, 13) {real, imag} */,
  {32'hbff2b08f, 32'hc17693db} /* (30, 18, 12) {real, imag} */,
  {32'hbff0ab29, 32'hc16dd0b0} /* (30, 18, 11) {real, imag} */,
  {32'h3fcb31ec, 32'h40918978} /* (30, 18, 10) {real, imag} */,
  {32'h400dc286, 32'h415a929f} /* (30, 18, 9) {real, imag} */,
  {32'h4056c8f2, 32'h41663c58} /* (30, 18, 8) {real, imag} */,
  {32'h3ffd7706, 32'h4180cee0} /* (30, 18, 7) {real, imag} */,
  {32'h3e6e1524, 32'h41705960} /* (30, 18, 6) {real, imag} */,
  {32'h3ff2937e, 32'h4184bb00} /* (30, 18, 5) {real, imag} */,
  {32'h40b3f756, 32'h417a704e} /* (30, 18, 4) {real, imag} */,
  {32'h40c5b7b4, 32'h41472763} /* (30, 18, 3) {real, imag} */,
  {32'h408704aa, 32'h41449405} /* (30, 18, 2) {real, imag} */,
  {32'h4026e35c, 32'h416e585a} /* (30, 18, 1) {real, imag} */,
  {32'h402c61de, 32'h4121d978} /* (30, 18, 0) {real, imag} */,
  {32'h40248ce2, 32'h40d929f2} /* (30, 17, 31) {real, imag} */,
  {32'h40c7ac8c, 32'h4166da44} /* (30, 17, 30) {real, imag} */,
  {32'h408dcdb4, 32'h4177a93a} /* (30, 17, 29) {real, imag} */,
  {32'h408bb4cd, 32'h4182159c} /* (30, 17, 28) {real, imag} */,
  {32'h4083947e, 32'h4181bc46} /* (30, 17, 27) {real, imag} */,
  {32'h405bc536, 32'h4157e101} /* (30, 17, 26) {real, imag} */,
  {32'h40837c7a, 32'h414fad3a} /* (30, 17, 25) {real, imag} */,
  {32'h40c38844, 32'h4160dae1} /* (30, 17, 24) {real, imag} */,
  {32'h4089882e, 32'h41950560} /* (30, 17, 23) {real, imag} */,
  {32'h4022a194, 32'h4173139d} /* (30, 17, 22) {real, imag} */,
  {32'h3ea8ff22, 32'h40e6dbd4} /* (30, 17, 21) {real, imag} */,
  {32'hbfb1765e, 32'hc1039cd4} /* (30, 17, 20) {real, imag} */,
  {32'hbf36ef18, 32'hc167e81c} /* (30, 17, 19) {real, imag} */,
  {32'hbfa53181, 32'hc18445c7} /* (30, 17, 18) {real, imag} */,
  {32'hc0947edc, 32'hc180a4d6} /* (30, 17, 17) {real, imag} */,
  {32'hc098db82, 32'hc16d57a6} /* (30, 17, 16) {real, imag} */,
  {32'hc07982a1, 32'hc155e8ec} /* (30, 17, 15) {real, imag} */,
  {32'hc0507893, 32'hc1458740} /* (30, 17, 14) {real, imag} */,
  {32'hc04647c0, 32'hc12eeefa} /* (30, 17, 13) {real, imag} */,
  {32'hbff1a5c1, 32'hc152ddf5} /* (30, 17, 12) {real, imag} */,
  {32'h3e87ed8c, 32'hc139f290} /* (30, 17, 11) {real, imag} */,
  {32'h4097d742, 32'h40c4ef6c} /* (30, 17, 10) {real, imag} */,
  {32'h40913a58, 32'h4141e8ca} /* (30, 17, 9) {real, imag} */,
  {32'h40730958, 32'h4162d3f4} /* (30, 17, 8) {real, imag} */,
  {32'h3fdc9c43, 32'h414a3b46} /* (30, 17, 7) {real, imag} */,
  {32'h40305274, 32'h417fedb2} /* (30, 17, 6) {real, imag} */,
  {32'h3fce0918, 32'h418631ae} /* (30, 17, 5) {real, imag} */,
  {32'h405b41b4, 32'h418aaa95} /* (30, 17, 4) {real, imag} */,
  {32'h40bc7e0a, 32'h4181bfe0} /* (30, 17, 3) {real, imag} */,
  {32'h407f6122, 32'h417ca7c6} /* (30, 17, 2) {real, imag} */,
  {32'hbf21b2a8, 32'h416a4c1e} /* (30, 17, 1) {real, imag} */,
  {32'h3e614880, 32'h40ff8926} /* (30, 17, 0) {real, imag} */,
  {32'h3f7c2d8c, 32'h40fcb814} /* (30, 16, 31) {real, imag} */,
  {32'h407702ad, 32'h4175ea4c} /* (30, 16, 30) {real, imag} */,
  {32'h40810b34, 32'h4160bd5a} /* (30, 16, 29) {real, imag} */,
  {32'h40c5ac54, 32'h41502a26} /* (30, 16, 28) {real, imag} */,
  {32'h40c06b03, 32'h4179dd76} /* (30, 16, 27) {real, imag} */,
  {32'h4036de60, 32'h416d4cfe} /* (30, 16, 26) {real, imag} */,
  {32'h400c4e65, 32'h41817538} /* (30, 16, 25) {real, imag} */,
  {32'h3f919e17, 32'h4187970c} /* (30, 16, 24) {real, imag} */,
  {32'h3eb64abe, 32'h4190ac72} /* (30, 16, 23) {real, imag} */,
  {32'h401befb1, 32'h41681114} /* (30, 16, 22) {real, imag} */,
  {32'h3fce5eec, 32'h407747fd} /* (30, 16, 21) {real, imag} */,
  {32'hbf7b9aa6, 32'hc1601302} /* (30, 16, 20) {real, imag} */,
  {32'hc00ed286, 32'hc1861d00} /* (30, 16, 19) {real, imag} */,
  {32'hc0480112, 32'hc179eaa7} /* (30, 16, 18) {real, imag} */,
  {32'hc09eaddb, 32'hc17b662e} /* (30, 16, 17) {real, imag} */,
  {32'hc09831da, 32'hc183e67a} /* (30, 16, 16) {real, imag} */,
  {32'hc0bdb1ce, 32'hc16f0c4e} /* (30, 16, 15) {real, imag} */,
  {32'hc0927377, 32'hc13e02de} /* (30, 16, 14) {real, imag} */,
  {32'hc0777918, 32'hc163cc96} /* (30, 16, 13) {real, imag} */,
  {32'hbfe48bed, 32'hc1812aa5} /* (30, 16, 12) {real, imag} */,
  {32'h3eb407aa, 32'hc138dacd} /* (30, 16, 11) {real, imag} */,
  {32'h407e1018, 32'h40c771c2} /* (30, 16, 10) {real, imag} */,
  {32'h40b8dc94, 32'h4163d402} /* (30, 16, 9) {real, imag} */,
  {32'h40c5c3b8, 32'h41693a3c} /* (30, 16, 8) {real, imag} */,
  {32'h40129c5b, 32'h414863e4} /* (30, 16, 7) {real, imag} */,
  {32'hbf4872ac, 32'h413eb3ec} /* (30, 16, 6) {real, imag} */,
  {32'hbfcdfb54, 32'h415bfd55} /* (30, 16, 5) {real, imag} */,
  {32'hbe611498, 32'h4164ffac} /* (30, 16, 4) {real, imag} */,
  {32'h40828ce3, 32'h4172c833} /* (30, 16, 3) {real, imag} */,
  {32'h4092307a, 32'h415bab00} /* (30, 16, 2) {real, imag} */,
  {32'h401b47ec, 32'h4156d3b2} /* (30, 16, 1) {real, imag} */,
  {32'h3eb0b51b, 32'h40f9a560} /* (30, 16, 0) {real, imag} */,
  {32'h3f6df2ed, 32'h4114d7a6} /* (30, 15, 31) {real, imag} */,
  {32'h4036884a, 32'h418c1504} /* (30, 15, 30) {real, imag} */,
  {32'h4072cd34, 32'h41858f04} /* (30, 15, 29) {real, imag} */,
  {32'h4069061e, 32'h41603b09} /* (30, 15, 28) {real, imag} */,
  {32'h40973be0, 32'h415f2bca} /* (30, 15, 27) {real, imag} */,
  {32'h4083aef2, 32'h4183b880} /* (30, 15, 26) {real, imag} */,
  {32'h40751733, 32'h4178aec2} /* (30, 15, 25) {real, imag} */,
  {32'h4034e0ac, 32'h415f051a} /* (30, 15, 24) {real, imag} */,
  {32'hbdd3c05c, 32'h41787658} /* (30, 15, 23) {real, imag} */,
  {32'h40880f95, 32'h416fb11b} /* (30, 15, 22) {real, imag} */,
  {32'h401ba26c, 32'h407aafe0} /* (30, 15, 21) {real, imag} */,
  {32'hc013894c, 32'hc138d42b} /* (30, 15, 20) {real, imag} */,
  {32'hbfbafdd9, 32'hc150d61c} /* (30, 15, 19) {real, imag} */,
  {32'hc0089aae, 32'hc14c0378} /* (30, 15, 18) {real, imag} */,
  {32'hc06f5296, 32'hc144a71c} /* (30, 15, 17) {real, imag} */,
  {32'hc055b716, 32'hc154e291} /* (30, 15, 16) {real, imag} */,
  {32'hc05ab234, 32'hc172efd0} /* (30, 15, 15) {real, imag} */,
  {32'hc043a42e, 32'hc1437a6f} /* (30, 15, 14) {real, imag} */,
  {32'hc079482c, 32'hc17e6541} /* (30, 15, 13) {real, imag} */,
  {32'hc0718df9, 32'hc191cb4a} /* (30, 15, 12) {real, imag} */,
  {32'hbffb4c58, 32'hc15f6e78} /* (30, 15, 11) {real, imag} */,
  {32'h403e79be, 32'h40ad9adc} /* (30, 15, 10) {real, imag} */,
  {32'h40b7e82b, 32'h416bea90} /* (30, 15, 9) {real, imag} */,
  {32'h40b60bbe, 32'h4181cdae} /* (30, 15, 8) {real, imag} */,
  {32'h40a7dea2, 32'h418bf8f3} /* (30, 15, 7) {real, imag} */,
  {32'h3fcc2f29, 32'h415ed9e4} /* (30, 15, 6) {real, imag} */,
  {32'hbe054b14, 32'h4166313f} /* (30, 15, 5) {real, imag} */,
  {32'h404f8163, 32'h41698046} /* (30, 15, 4) {real, imag} */,
  {32'h40a36b83, 32'h416b87a4} /* (30, 15, 3) {real, imag} */,
  {32'h40d59c49, 32'h414cdf3d} /* (30, 15, 2) {real, imag} */,
  {32'h40b3d0a8, 32'h416e9026} /* (30, 15, 1) {real, imag} */,
  {32'h3fe8591a, 32'h4115ed41} /* (30, 15, 0) {real, imag} */,
  {32'h3f2e44b8, 32'h410ccc4a} /* (30, 14, 31) {real, imag} */,
  {32'h40045784, 32'h4184a7c2} /* (30, 14, 30) {real, imag} */,
  {32'h3fdba09b, 32'h418e7b40} /* (30, 14, 29) {real, imag} */,
  {32'h40080326, 32'h41834504} /* (30, 14, 28) {real, imag} */,
  {32'h406aa9b8, 32'h415e4ce4} /* (30, 14, 27) {real, imag} */,
  {32'h408a549e, 32'h41569b14} /* (30, 14, 26) {real, imag} */,
  {32'h40891db7, 32'h4147824e} /* (30, 14, 25) {real, imag} */,
  {32'h3f81df8e, 32'h414c4068} /* (30, 14, 24) {real, imag} */,
  {32'h3f1a00a8, 32'h416132a4} /* (30, 14, 23) {real, imag} */,
  {32'h40aa0708, 32'h4186f8d2} /* (30, 14, 22) {real, imag} */,
  {32'h4069b2c2, 32'h40f22889} /* (30, 14, 21) {real, imag} */,
  {32'hbfeffc48, 32'hc12ba3e5} /* (30, 14, 20) {real, imag} */,
  {32'hc067685c, 32'hc151e210} /* (30, 14, 19) {real, imag} */,
  {32'hc0413113, 32'hc146cb30} /* (30, 14, 18) {real, imag} */,
  {32'hbfadba1b, 32'hc157617f} /* (30, 14, 17) {real, imag} */,
  {32'hbe407ed2, 32'hc15c0017} /* (30, 14, 16) {real, imag} */,
  {32'hbf825958, 32'hc1759822} /* (30, 14, 15) {real, imag} */,
  {32'hc09baae3, 32'hc159ac36} /* (30, 14, 14) {real, imag} */,
  {32'hc0a0cb84, 32'hc159cd9f} /* (30, 14, 13) {real, imag} */,
  {32'hc04dac30, 32'hc168f73c} /* (30, 14, 12) {real, imag} */,
  {32'hbf03ff20, 32'hc1438bdd} /* (30, 14, 11) {real, imag} */,
  {32'h4051db1e, 32'h4039987c} /* (30, 14, 10) {real, imag} */,
  {32'h40a3c585, 32'h4161c732} /* (30, 14, 9) {real, imag} */,
  {32'h4049b4ff, 32'h41886413} /* (30, 14, 8) {real, imag} */,
  {32'h403b4157, 32'h4184963a} /* (30, 14, 7) {real, imag} */,
  {32'h3fb9d12a, 32'h414d94cc} /* (30, 14, 6) {real, imag} */,
  {32'h3d7d6c00, 32'h4137ceb8} /* (30, 14, 5) {real, imag} */,
  {32'h3fbbdefb, 32'h412f265c} /* (30, 14, 4) {real, imag} */,
  {32'h40832c30, 32'h4141c34d} /* (30, 14, 3) {real, imag} */,
  {32'h40d1915e, 32'h41529554} /* (30, 14, 2) {real, imag} */,
  {32'h409c5a0e, 32'h41885cfe} /* (30, 14, 1) {real, imag} */,
  {32'h3edf19b8, 32'h41324645} /* (30, 14, 0) {real, imag} */,
  {32'h3f7230b0, 32'h4107254e} /* (30, 13, 31) {real, imag} */,
  {32'h404a2108, 32'h417f7f5c} /* (30, 13, 30) {real, imag} */,
  {32'h408e5b3c, 32'h418bd9a4} /* (30, 13, 29) {real, imag} */,
  {32'h4032ad42, 32'h418fb20c} /* (30, 13, 28) {real, imag} */,
  {32'h3f1be061, 32'h415ec1e2} /* (30, 13, 27) {real, imag} */,
  {32'h407be294, 32'h413d5c26} /* (30, 13, 26) {real, imag} */,
  {32'h40a7fcdb, 32'h413a4b45} /* (30, 13, 25) {real, imag} */,
  {32'h3f9519e2, 32'h414d8f06} /* (30, 13, 24) {real, imag} */,
  {32'h3e0cb07c, 32'h41450bb4} /* (30, 13, 23) {real, imag} */,
  {32'h4027dcce, 32'h41891bf4} /* (30, 13, 22) {real, imag} */,
  {32'h3e22f6b0, 32'h4116bf44} /* (30, 13, 21) {real, imag} */,
  {32'hc04bcfd2, 32'hc1297bc2} /* (30, 13, 20) {real, imag} */,
  {32'hc0054a34, 32'hc18774f8} /* (30, 13, 19) {real, imag} */,
  {32'hc0100e5c, 32'hc16cff8a} /* (30, 13, 18) {real, imag} */,
  {32'hc043ccb0, 32'hc172c18e} /* (30, 13, 17) {real, imag} */,
  {32'hc041f0ef, 32'hc1485542} /* (30, 13, 16) {real, imag} */,
  {32'hbfd1108f, 32'hc132762e} /* (30, 13, 15) {real, imag} */,
  {32'hc03ec7bf, 32'hc15bda37} /* (30, 13, 14) {real, imag} */,
  {32'hc03f66d0, 32'hc15505fa} /* (30, 13, 13) {real, imag} */,
  {32'hbfdc1127, 32'hc145e167} /* (30, 13, 12) {real, imag} */,
  {32'hbf9b7a30, 32'hc12b2d48} /* (30, 13, 11) {real, imag} */,
  {32'h3ffd092c, 32'h40848cf6} /* (30, 13, 10) {real, imag} */,
  {32'h40a067e0, 32'h41475582} /* (30, 13, 9) {real, imag} */,
  {32'h4014f1c8, 32'h41862f5e} /* (30, 13, 8) {real, imag} */,
  {32'h4006b3fc, 32'h4183adfe} /* (30, 13, 7) {real, imag} */,
  {32'h3e8346f4, 32'h4143fc1b} /* (30, 13, 6) {real, imag} */,
  {32'hbe1ab5d4, 32'h412ec3b0} /* (30, 13, 5) {real, imag} */,
  {32'hbed16703, 32'h410d597c} /* (30, 13, 4) {real, imag} */,
  {32'h408f5434, 32'h412d37e0} /* (30, 13, 3) {real, imag} */,
  {32'h40c2bf2d, 32'h414d20a5} /* (30, 13, 2) {real, imag} */,
  {32'h408673f7, 32'h4184ef24} /* (30, 13, 1) {real, imag} */,
  {32'h3f5c4113, 32'h4130b131} /* (30, 13, 0) {real, imag} */,
  {32'hbe777d66, 32'h40eee60e} /* (30, 12, 31) {real, imag} */,
  {32'h3faf8b52, 32'h415e1a63} /* (30, 12, 30) {real, imag} */,
  {32'h4079a5bf, 32'h4163fce6} /* (30, 12, 29) {real, imag} */,
  {32'h40583f1b, 32'h41809afb} /* (30, 12, 28) {real, imag} */,
  {32'h3fd6a3ee, 32'h4162ee44} /* (30, 12, 27) {real, imag} */,
  {32'h4050e364, 32'h412883b4} /* (30, 12, 26) {real, imag} */,
  {32'h40c444ac, 32'h41258680} /* (30, 12, 25) {real, imag} */,
  {32'h409ec35d, 32'h414bc10e} /* (30, 12, 24) {real, imag} */,
  {32'h4041d396, 32'h4167d02c} /* (30, 12, 23) {real, imag} */,
  {32'h3fbd3f7e, 32'h4190366e} /* (30, 12, 22) {real, imag} */,
  {32'h4018452c, 32'h41006618} /* (30, 12, 21) {real, imag} */,
  {32'hbf475efa, 32'hc123411c} /* (30, 12, 20) {real, imag} */,
  {32'h3faa49dc, 32'hc19c9c8a} /* (30, 12, 19) {real, imag} */,
  {32'h403d405c, 32'hc1861e3a} /* (30, 12, 18) {real, imag} */,
  {32'hbeb2c9e8, 32'hc187b7ec} /* (30, 12, 17) {real, imag} */,
  {32'hc06e02c8, 32'hc16e0364} /* (30, 12, 16) {real, imag} */,
  {32'hc08dd4d7, 32'hc137356e} /* (30, 12, 15) {real, imag} */,
  {32'hc085a03e, 32'hc1683f1c} /* (30, 12, 14) {real, imag} */,
  {32'hbf9e9ace, 32'hc156373a} /* (30, 12, 13) {real, imag} */,
  {32'h3e69f514, 32'hc1303cd1} /* (30, 12, 12) {real, imag} */,
  {32'h3fcf2f5a, 32'hc111f349} /* (30, 12, 11) {real, imag} */,
  {32'hbde92edc, 32'h40eb70a4} /* (30, 12, 10) {real, imag} */,
  {32'h402734b4, 32'h414ec5fe} /* (30, 12, 9) {real, imag} */,
  {32'h3f3cf854, 32'h4162eaef} /* (30, 12, 8) {real, imag} */,
  {32'h4062e213, 32'h418054e0} /* (30, 12, 7) {real, imag} */,
  {32'h408950fe, 32'h41670ac4} /* (30, 12, 6) {real, imag} */,
  {32'h402bbbd0, 32'h415416eb} /* (30, 12, 5) {real, imag} */,
  {32'h40106ac1, 32'h4142474e} /* (30, 12, 4) {real, imag} */,
  {32'h403e7cf2, 32'h4174083c} /* (30, 12, 3) {real, imag} */,
  {32'h400f836c, 32'h4170f980} /* (30, 12, 2) {real, imag} */,
  {32'h40110265, 32'h418b031e} /* (30, 12, 1) {real, imag} */,
  {32'h3f9177ae, 32'h41097857} /* (30, 12, 0) {real, imag} */,
  {32'h3e5eee54, 32'h4095946a} /* (30, 11, 31) {real, imag} */,
  {32'h3ee96381, 32'h410c50a8} /* (30, 11, 30) {real, imag} */,
  {32'h3fde0ba0, 32'h410c3f93} /* (30, 11, 29) {real, imag} */,
  {32'h3fd489d4, 32'h414d8e01} /* (30, 11, 28) {real, imag} */,
  {32'h3fadbb6c, 32'h412b531c} /* (30, 11, 27) {real, imag} */,
  {32'hbf518947, 32'h410c4d49} /* (30, 11, 26) {real, imag} */,
  {32'h3fd0443a, 32'h410b1500} /* (30, 11, 25) {real, imag} */,
  {32'h3fdddfee, 32'h411fd9ec} /* (30, 11, 24) {real, imag} */,
  {32'hbfa47d48, 32'h41365fce} /* (30, 11, 23) {real, imag} */,
  {32'hbfabfee8, 32'h4135757c} /* (30, 11, 22) {real, imag} */,
  {32'h406f449a, 32'h40550988} /* (30, 11, 21) {real, imag} */,
  {32'h3e967070, 32'hc0e9d56c} /* (30, 11, 20) {real, imag} */,
  {32'h3e311f45, 32'hc14983bd} /* (30, 11, 19) {real, imag} */,
  {32'h3f76c4c3, 32'hc1437e86} /* (30, 11, 18) {real, imag} */,
  {32'h3fa7230a, 32'hc1702826} /* (30, 11, 17) {real, imag} */,
  {32'hc02b0c6a, 32'hc145d38d} /* (30, 11, 16) {real, imag} */,
  {32'hc09dc27e, 32'hc1256b5c} /* (30, 11, 15) {real, imag} */,
  {32'hc083f2ce, 32'hc140f63a} /* (30, 11, 14) {real, imag} */,
  {32'hc01a5e88, 32'hc140413e} /* (30, 11, 13) {real, imag} */,
  {32'hbfe8c569, 32'hc1202157} /* (30, 11, 12) {real, imag} */,
  {32'h3f0b5df5, 32'hc0bac488} /* (30, 11, 11) {real, imag} */,
  {32'h3f2370b1, 32'h41084442} /* (30, 11, 10) {real, imag} */,
  {32'h3f615a6f, 32'h4131839b} /* (30, 11, 9) {real, imag} */,
  {32'h3f9c303c, 32'h411e3a32} /* (30, 11, 8) {real, imag} */,
  {32'hbe5b2dda, 32'h414207d2} /* (30, 11, 7) {real, imag} */,
  {32'h408f0f0a, 32'h41483840} /* (30, 11, 6) {real, imag} */,
  {32'h40aa971f, 32'h4106830f} /* (30, 11, 5) {real, imag} */,
  {32'h402e15e9, 32'h4102ec99} /* (30, 11, 4) {real, imag} */,
  {32'h3fe80430, 32'h41378e16} /* (30, 11, 3) {real, imag} */,
  {32'h4039670c, 32'h4127817a} /* (30, 11, 2) {real, imag} */,
  {32'h4054e744, 32'h41383d49} /* (30, 11, 1) {real, imag} */,
  {32'h3f65b1e5, 32'h40c086d3} /* (30, 11, 0) {real, imag} */,
  {32'hbd6ce0f4, 32'hc0bc47ec} /* (30, 10, 31) {real, imag} */,
  {32'h3dd04e50, 32'hc0e4bcec} /* (30, 10, 30) {real, imag} */,
  {32'h3fd2bf4f, 32'hc0ed4cae} /* (30, 10, 29) {real, imag} */,
  {32'hbf816082, 32'hc0e14596} /* (30, 10, 28) {real, imag} */,
  {32'hc0629b4b, 32'hc1084f32} /* (30, 10, 27) {real, imag} */,
  {32'hc076035f, 32'hc0d9335a} /* (30, 10, 26) {real, imag} */,
  {32'hc016b34b, 32'hc0b8da0a} /* (30, 10, 25) {real, imag} */,
  {32'hc058ee37, 32'hc0f8ffc1} /* (30, 10, 24) {real, imag} */,
  {32'hc08bbbc8, 32'hc0dbd30d} /* (30, 10, 23) {real, imag} */,
  {32'hc02591a7, 32'hc1050b4d} /* (30, 10, 22) {real, imag} */,
  {32'hbf8602ef, 32'hc099445a} /* (30, 10, 21) {real, imag} */,
  {32'hbef103af, 32'h40950036} /* (30, 10, 20) {real, imag} */,
  {32'h3f9756f0, 32'h40e36416} /* (30, 10, 19) {real, imag} */,
  {32'h400d5dbe, 32'h40a9a037} /* (30, 10, 18) {real, imag} */,
  {32'h3fe795b8, 32'h404ccd0a} /* (30, 10, 17) {real, imag} */,
  {32'h3f8cd445, 32'h40c1ba76} /* (30, 10, 16) {real, imag} */,
  {32'hbf91b779, 32'h40d4e461} /* (30, 10, 15) {real, imag} */,
  {32'hbeb9e4f6, 32'h407189a4} /* (30, 10, 14) {real, imag} */,
  {32'h3f76ad58, 32'h4067c845} /* (30, 10, 13) {real, imag} */,
  {32'h3fdc2cbe, 32'h40e4dbb6} /* (30, 10, 12) {real, imag} */,
  {32'h401b9282, 32'h40d78261} /* (30, 10, 11) {real, imag} */,
  {32'h3f334d67, 32'h3eca6a65} /* (30, 10, 10) {real, imag} */,
  {32'hc000f4cd, 32'hc0b4495a} /* (30, 10, 9) {real, imag} */,
  {32'hbfa3cf0f, 32'hc0ae12c2} /* (30, 10, 8) {real, imag} */,
  {32'hc0baa72c, 32'hc0d6461b} /* (30, 10, 7) {real, imag} */,
  {32'hbf85b150, 32'hc0fe01d1} /* (30, 10, 6) {real, imag} */,
  {32'hbf6c6867, 32'hc117857b} /* (30, 10, 5) {real, imag} */,
  {32'hbb09b800, 32'hc119ef8a} /* (30, 10, 4) {real, imag} */,
  {32'h40459a6a, 32'hc0cf786c} /* (30, 10, 3) {real, imag} */,
  {32'h3fe8ac23, 32'hc0e331e6} /* (30, 10, 2) {real, imag} */,
  {32'hbebbf837, 32'hc0f0147a} /* (30, 10, 1) {real, imag} */,
  {32'hbfcdabb4, 32'hc0c83a28} /* (30, 10, 0) {real, imag} */,
  {32'hc0254c98, 32'hc10c36b4} /* (30, 9, 31) {real, imag} */,
  {32'hc055f853, 32'hc165e18a} /* (30, 9, 30) {real, imag} */,
  {32'hbf59642c, 32'hc1806803} /* (30, 9, 29) {real, imag} */,
  {32'hc01a0926, 32'hc18debe0} /* (30, 9, 28) {real, imag} */,
  {32'hc03473d5, 32'hc16c75eb} /* (30, 9, 27) {real, imag} */,
  {32'hbfa881b4, 32'hc15b6a70} /* (30, 9, 26) {real, imag} */,
  {32'hc0338633, 32'hc140c15a} /* (30, 9, 25) {real, imag} */,
  {32'hc00f0674, 32'hc1739bd6} /* (30, 9, 24) {real, imag} */,
  {32'hc086cf16, 32'hc14e38d4} /* (30, 9, 23) {real, imag} */,
  {32'hc0a67042, 32'hc15c31f6} /* (30, 9, 22) {real, imag} */,
  {32'hc0307e90, 32'hc10ec7ac} /* (30, 9, 21) {real, imag} */,
  {32'hbeb9ecb0, 32'h40f17206} /* (30, 9, 20) {real, imag} */,
  {32'h404325bb, 32'h41491124} /* (30, 9, 19) {real, imag} */,
  {32'h40283b6e, 32'h415dbd00} /* (30, 9, 18) {real, imag} */,
  {32'h405086ea, 32'h415f022e} /* (30, 9, 17) {real, imag} */,
  {32'h40918270, 32'h41863786} /* (30, 9, 16) {real, imag} */,
  {32'h407b73f8, 32'h4197f9e5} /* (30, 9, 15) {real, imag} */,
  {32'h3fea1e35, 32'h415d5ae2} /* (30, 9, 14) {real, imag} */,
  {32'h4058b657, 32'h412ec9ba} /* (30, 9, 13) {real, imag} */,
  {32'h406460e6, 32'h41783314} /* (30, 9, 12) {real, imag} */,
  {32'h40257886, 32'h413f68c8} /* (30, 9, 11) {real, imag} */,
  {32'hbee81c51, 32'hc0c0bcee} /* (30, 9, 10) {real, imag} */,
  {32'hc02617ac, 32'hc17a4a8a} /* (30, 9, 9) {real, imag} */,
  {32'hc031d668, 32'hc1541c9f} /* (30, 9, 8) {real, imag} */,
  {32'hc0991bec, 32'hc1413ba8} /* (30, 9, 7) {real, imag} */,
  {32'hbfab6dd5, 32'hc1596413} /* (30, 9, 6) {real, imag} */,
  {32'hc0260c18, 32'hc16a5b05} /* (30, 9, 5) {real, imag} */,
  {32'hbfba99db, 32'hc181c03c} /* (30, 9, 4) {real, imag} */,
  {32'h3f7a21c5, 32'hc1741581} /* (30, 9, 3) {real, imag} */,
  {32'hbf7047f4, 32'hc14dcea1} /* (30, 9, 2) {real, imag} */,
  {32'hbfec943e, 32'hc150720d} /* (30, 9, 1) {real, imag} */,
  {32'hc010b2bb, 32'hc10e086b} /* (30, 9, 0) {real, imag} */,
  {32'hc05be5bb, 32'hc1000b0e} /* (30, 8, 31) {real, imag} */,
  {32'hc040bfb1, 32'hc15a4770} /* (30, 8, 30) {real, imag} */,
  {32'hbff7fce6, 32'hc1790fc2} /* (30, 8, 29) {real, imag} */,
  {32'hbfcabbe1, 32'hc178df1a} /* (30, 8, 28) {real, imag} */,
  {32'hc022a408, 32'hc17958a8} /* (30, 8, 27) {real, imag} */,
  {32'hbff25a4f, 32'hc18980db} /* (30, 8, 26) {real, imag} */,
  {32'hbd735550, 32'hc15c9464} /* (30, 8, 25) {real, imag} */,
  {32'h3dc1ac48, 32'hc167d216} /* (30, 8, 24) {real, imag} */,
  {32'hc09956fc, 32'hc152896d} /* (30, 8, 23) {real, imag} */,
  {32'hc09388b6, 32'hc165d60d} /* (30, 8, 22) {real, imag} */,
  {32'h3edba324, 32'hc100fd68} /* (30, 8, 21) {real, imag} */,
  {32'hbeb9f780, 32'h41064036} /* (30, 8, 20) {real, imag} */,
  {32'h40087b96, 32'h4155f265} /* (30, 8, 19) {real, imag} */,
  {32'h403cea72, 32'h417052ae} /* (30, 8, 18) {real, imag} */,
  {32'h40893214, 32'h4158f286} /* (30, 8, 17) {real, imag} */,
  {32'h40c0f56e, 32'h4159bf23} /* (30, 8, 16) {real, imag} */,
  {32'h4079008b, 32'h419a2c71} /* (30, 8, 15) {real, imag} */,
  {32'h4052b547, 32'h417b2e80} /* (30, 8, 14) {real, imag} */,
  {32'h3fd9774a, 32'h41150dc6} /* (30, 8, 13) {real, imag} */,
  {32'hbda93f24, 32'h416312cc} /* (30, 8, 12) {real, imag} */,
  {32'hbe4ce4a8, 32'h41541082} /* (30, 8, 11) {real, imag} */,
  {32'hc0837890, 32'hc0bd6183} /* (30, 8, 10) {real, imag} */,
  {32'hc08c04a6, 32'hc171190b} /* (30, 8, 9) {real, imag} */,
  {32'hc022e856, 32'hc14f2f86} /* (30, 8, 8) {real, imag} */,
  {32'hbf873892, 32'hc13a8d5c} /* (30, 8, 7) {real, imag} */,
  {32'h3e4fd640, 32'hc165bc08} /* (30, 8, 6) {real, imag} */,
  {32'hc008059a, 32'hc16217f5} /* (30, 8, 5) {real, imag} */,
  {32'hc093fea0, 32'hc165e434} /* (30, 8, 4) {real, imag} */,
  {32'hc012d35d, 32'hc16119d0} /* (30, 8, 3) {real, imag} */,
  {32'hc01d5a19, 32'hc151828d} /* (30, 8, 2) {real, imag} */,
  {32'hc02a57cc, 32'hc14d8cf0} /* (30, 8, 1) {real, imag} */,
  {32'hc05e6fa0, 32'hc0cfb576} /* (30, 8, 0) {real, imag} */,
  {32'hc0353c1a, 32'hc0f38f3d} /* (30, 7, 31) {real, imag} */,
  {32'hc0345b08, 32'hc13fa5b9} /* (30, 7, 30) {real, imag} */,
  {32'hc0286922, 32'hc15b2d8a} /* (30, 7, 29) {real, imag} */,
  {32'hbf71d983, 32'hc1435194} /* (30, 7, 28) {real, imag} */,
  {32'hc04135ca, 32'hc161c90e} /* (30, 7, 27) {real, imag} */,
  {32'hc0795b88, 32'hc18c8cca} /* (30, 7, 26) {real, imag} */,
  {32'hc003891c, 32'hc18f69e6} /* (30, 7, 25) {real, imag} */,
  {32'hc05623f9, 32'hc1898c53} /* (30, 7, 24) {real, imag} */,
  {32'hc0725166, 32'hc14a8ca3} /* (30, 7, 23) {real, imag} */,
  {32'hc065d886, 32'hc159823a} /* (30, 7, 22) {real, imag} */,
  {32'hc072ad98, 32'hc109f6be} /* (30, 7, 21) {real, imag} */,
  {32'hc02754a4, 32'h412e9ab1} /* (30, 7, 20) {real, imag} */,
  {32'h3fa35d6d, 32'h41718477} /* (30, 7, 19) {real, imag} */,
  {32'h409a2e72, 32'h4175247f} /* (30, 7, 18) {real, imag} */,
  {32'h40b79a3a, 32'h41844084} /* (30, 7, 17) {real, imag} */,
  {32'h40af33e0, 32'h41698897} /* (30, 7, 16) {real, imag} */,
  {32'h40c4f368, 32'h417bb7f9} /* (30, 7, 15) {real, imag} */,
  {32'h40c373fb, 32'h41676f5f} /* (30, 7, 14) {real, imag} */,
  {32'h408f0756, 32'h41196658} /* (30, 7, 13) {real, imag} */,
  {32'h406e733e, 32'h415b6c08} /* (30, 7, 12) {real, imag} */,
  {32'h404b71b0, 32'h413f5ea7} /* (30, 7, 11) {real, imag} */,
  {32'hc0171887, 32'hc0b29a24} /* (30, 7, 10) {real, imag} */,
  {32'hc0a1a356, 32'hc138ed86} /* (30, 7, 9) {real, imag} */,
  {32'hc04f7fa0, 32'hc13fe5b8} /* (30, 7, 8) {real, imag} */,
  {32'hbfc9fad6, 32'hc1689ef8} /* (30, 7, 7) {real, imag} */,
  {32'hc00ef2a4, 32'hc1806acc} /* (30, 7, 6) {real, imag} */,
  {32'hbff03aa7, 32'hc18a161f} /* (30, 7, 5) {real, imag} */,
  {32'hc0ad888c, 32'hc192d084} /* (30, 7, 4) {real, imag} */,
  {32'hc0829f18, 32'hc1821926} /* (30, 7, 3) {real, imag} */,
  {32'hc016433a, 32'hc16de660} /* (30, 7, 2) {real, imag} */,
  {32'hc0377c56, 32'hc1446287} /* (30, 7, 1) {real, imag} */,
  {32'hbffd5208, 32'hc0b240bb} /* (30, 7, 0) {real, imag} */,
  {32'hbf9ba987, 32'hc0d1c411} /* (30, 6, 31) {real, imag} */,
  {32'hc059d930, 32'hc102fe34} /* (30, 6, 30) {real, imag} */,
  {32'hc08646b6, 32'hc15375fa} /* (30, 6, 29) {real, imag} */,
  {32'hc01601f9, 32'hc13f12f1} /* (30, 6, 28) {real, imag} */,
  {32'hc0754b05, 32'hc14c6112} /* (30, 6, 27) {real, imag} */,
  {32'hc0c96764, 32'hc17943c6} /* (30, 6, 26) {real, imag} */,
  {32'hc0b31774, 32'hc186c383} /* (30, 6, 25) {real, imag} */,
  {32'hc0979de8, 32'hc159e994} /* (30, 6, 24) {real, imag} */,
  {32'hc019fd9c, 32'hc122edd1} /* (30, 6, 23) {real, imag} */,
  {32'hc053e515, 32'hc13c0afa} /* (30, 6, 22) {real, imag} */,
  {32'hc076f21d, 32'hc12d8eae} /* (30, 6, 21) {real, imag} */,
  {32'h401467aa, 32'h40a362ec} /* (30, 6, 20) {real, imag} */,
  {32'h405d4dec, 32'h41262b18} /* (30, 6, 19) {real, imag} */,
  {32'h400d403b, 32'h41564b0a} /* (30, 6, 18) {real, imag} */,
  {32'h4011959d, 32'h41545a84} /* (30, 6, 17) {real, imag} */,
  {32'h408f3d67, 32'h4163087a} /* (30, 6, 16) {real, imag} */,
  {32'h40a0c56e, 32'h416789fa} /* (30, 6, 15) {real, imag} */,
  {32'h406db0ee, 32'h418b3ade} /* (30, 6, 14) {real, imag} */,
  {32'h406fe94a, 32'h41761d52} /* (30, 6, 13) {real, imag} */,
  {32'h4085f678, 32'h4169169a} /* (30, 6, 12) {real, imag} */,
  {32'h4070c070, 32'h41314468} /* (30, 6, 11) {real, imag} */,
  {32'hbf3a5ea9, 32'hc02395b9} /* (30, 6, 10) {real, imag} */,
  {32'hc087e63c, 32'hc126223f} /* (30, 6, 9) {real, imag} */,
  {32'hc0769526, 32'hc13c3408} /* (30, 6, 8) {real, imag} */,
  {32'hbfaafb90, 32'hc13d6f79} /* (30, 6, 7) {real, imag} */,
  {32'hc003a184, 32'hc1540f97} /* (30, 6, 6) {real, imag} */,
  {32'hc0a04c7c, 32'hc142345d} /* (30, 6, 5) {real, imag} */,
  {32'hc085cdbc, 32'hc16d8a42} /* (30, 6, 4) {real, imag} */,
  {32'hc04c9e71, 32'hc170da3e} /* (30, 6, 3) {real, imag} */,
  {32'hc0a0c842, 32'hc160d6b2} /* (30, 6, 2) {real, imag} */,
  {32'hc038d7be, 32'hc1520940} /* (30, 6, 1) {real, imag} */,
  {32'hbf46790c, 32'hc0e0a89c} /* (30, 6, 0) {real, imag} */,
  {32'hbfd88a78, 32'hc0bcf6be} /* (30, 5, 31) {real, imag} */,
  {32'hbf53b20a, 32'hc140703d} /* (30, 5, 30) {real, imag} */,
  {32'hc0163ee6, 32'hc18b33c4} /* (30, 5, 29) {real, imag} */,
  {32'hbfe799a3, 32'hc1705050} /* (30, 5, 28) {real, imag} */,
  {32'hc093f1f5, 32'hc183193e} /* (30, 5, 27) {real, imag} */,
  {32'hc09cd44e, 32'hc184dc7a} /* (30, 5, 26) {real, imag} */,
  {32'hc07d52d4, 32'hc17b9a4d} /* (30, 5, 25) {real, imag} */,
  {32'hbfdcd53b, 32'hc1720bb1} /* (30, 5, 24) {real, imag} */,
  {32'hc09f6272, 32'hc14f0a34} /* (30, 5, 23) {real, imag} */,
  {32'hc0ace72a, 32'hc149de0d} /* (30, 5, 22) {real, imag} */,
  {32'hc005b348, 32'hc164b32a} /* (30, 5, 21) {real, imag} */,
  {32'hbf17e261, 32'hc11fea44} /* (30, 5, 20) {real, imag} */,
  {32'hbfa40210, 32'hc0900374} /* (30, 5, 19) {real, imag} */,
  {32'hbfb2748f, 32'hbffac7e8} /* (30, 5, 18) {real, imag} */,
  {32'hc035e0fa, 32'hc0960959} /* (30, 5, 17) {real, imag} */,
  {32'hbd16cfe8, 32'h3efe768e} /* (30, 5, 16) {real, imag} */,
  {32'h3fb6c016, 32'h410e0306} /* (30, 5, 15) {real, imag} */,
  {32'h4007e0be, 32'h4160fc60} /* (30, 5, 14) {real, imag} */,
  {32'h402e1f86, 32'h41540993} /* (30, 5, 13) {real, imag} */,
  {32'h40898652, 32'h4163fab1} /* (30, 5, 12) {real, imag} */,
  {32'h40632818, 32'h4181d21b} /* (30, 5, 11) {real, imag} */,
  {32'hbfc269fa, 32'h411cf982} /* (30, 5, 10) {real, imag} */,
  {32'hbf78d2c7, 32'h4032aab0} /* (30, 5, 9) {real, imag} */,
  {32'hbf4af91a, 32'h4063137f} /* (30, 5, 8) {real, imag} */,
  {32'hbfbc1048, 32'h40b9a1a7} /* (30, 5, 7) {real, imag} */,
  {32'hbd33c4d8, 32'h401bebfc} /* (30, 5, 6) {real, imag} */,
  {32'hbfc64b67, 32'hc0cc2f81} /* (30, 5, 5) {real, imag} */,
  {32'hbffc1679, 32'hc14570bb} /* (30, 5, 4) {real, imag} */,
  {32'hbfbd31f8, 32'hc176c134} /* (30, 5, 3) {real, imag} */,
  {32'hc0a5d6b2, 32'hc15f64be} /* (30, 5, 2) {real, imag} */,
  {32'hc0b5f0d3, 32'hc14dd6bc} /* (30, 5, 1) {real, imag} */,
  {32'hc019788d, 32'hc0ee8942} /* (30, 5, 0) {real, imag} */,
  {32'hc0227103, 32'hc0dfaf08} /* (30, 4, 31) {real, imag} */,
  {32'hc064d6c6, 32'hc166acfa} /* (30, 4, 30) {real, imag} */,
  {32'hc05bce11, 32'hc1906d3e} /* (30, 4, 29) {real, imag} */,
  {32'hbfe561a5, 32'hc181f9ca} /* (30, 4, 28) {real, imag} */,
  {32'hc0482d6e, 32'hc17e9be9} /* (30, 4, 27) {real, imag} */,
  {32'hc00be1bb, 32'hc156b2d8} /* (30, 4, 26) {real, imag} */,
  {32'hbf08e2c8, 32'hc1439a2e} /* (30, 4, 25) {real, imag} */,
  {32'h3f4b6805, 32'hc17985a6} /* (30, 4, 24) {real, imag} */,
  {32'hc040d33a, 32'hc17699d4} /* (30, 4, 23) {real, imag} */,
  {32'hc081ee9b, 32'hc16fe47b} /* (30, 4, 22) {real, imag} */,
  {32'hc04d5bbd, 32'hc19479b8} /* (30, 4, 21) {real, imag} */,
  {32'hc0670d08, 32'hc1906ed2} /* (30, 4, 20) {real, imag} */,
  {32'hc03eea3d, 32'hc15e9d1a} /* (30, 4, 19) {real, imag} */,
  {32'hc023bc0e, 32'hc1569dac} /* (30, 4, 18) {real, imag} */,
  {32'hc0997415, 32'hc17152c4} /* (30, 4, 17) {real, imag} */,
  {32'hc00db662, 32'hc120451d} /* (30, 4, 16) {real, imag} */,
  {32'h40110925, 32'h40b4c20a} /* (30, 4, 15) {real, imag} */,
  {32'h4045345a, 32'h4136a7db} /* (30, 4, 14) {real, imag} */,
  {32'h3fadc388, 32'h413d57cc} /* (30, 4, 13) {real, imag} */,
  {32'h409568c3, 32'h4127c508} /* (30, 4, 12) {real, imag} */,
  {32'h40804d1c, 32'h4165b6ab} /* (30, 4, 11) {real, imag} */,
  {32'hbe716550, 32'h4180b914} /* (30, 4, 10) {real, imag} */,
  {32'h3fbf8557, 32'h41683f2a} /* (30, 4, 9) {real, imag} */,
  {32'h40334b90, 32'h41777614} /* (30, 4, 8) {real, imag} */,
  {32'h3fba6b75, 32'h4165fac8} /* (30, 4, 7) {real, imag} */,
  {32'h401f3834, 32'h413b1850} /* (30, 4, 6) {real, imag} */,
  {32'hbeafa313, 32'hc0bad6a4} /* (30, 4, 5) {real, imag} */,
  {32'hc0320b2e, 32'hc15bb8f6} /* (30, 4, 4) {real, imag} */,
  {32'hc0342d5a, 32'hc17e626e} /* (30, 4, 3) {real, imag} */,
  {32'hc0515c0b, 32'hc1752ff9} /* (30, 4, 2) {real, imag} */,
  {32'hc0bbb685, 32'hc12cf854} /* (30, 4, 1) {real, imag} */,
  {32'hc0353f81, 32'hc0ba6936} /* (30, 4, 0) {real, imag} */,
  {32'h3ded73f0, 32'hc0f6dcef} /* (30, 3, 31) {real, imag} */,
  {32'hc094dde2, 32'hc186d9c6} /* (30, 3, 30) {real, imag} */,
  {32'hc06bdae6, 32'hc18f2a68} /* (30, 3, 29) {real, imag} */,
  {32'h3e953541, 32'hc17ce517} /* (30, 3, 28) {real, imag} */,
  {32'h3ed1eb4c, 32'hc1623a4d} /* (30, 3, 27) {real, imag} */,
  {32'hbfb3b025, 32'hc138bccd} /* (30, 3, 26) {real, imag} */,
  {32'hc0815b91, 32'hc13629b8} /* (30, 3, 25) {real, imag} */,
  {32'hc089f202, 32'hc17286f4} /* (30, 3, 24) {real, imag} */,
  {32'hc04023fc, 32'hc17c9c14} /* (30, 3, 23) {real, imag} */,
  {32'hc02a4cc0, 32'hc18176e1} /* (30, 3, 22) {real, imag} */,
  {32'hc04ce9a6, 32'hc1752e62} /* (30, 3, 21) {real, imag} */,
  {32'hc02de4ae, 32'hc1736ac6} /* (30, 3, 20) {real, imag} */,
  {32'hc0c4e470, 32'hc16967be} /* (30, 3, 19) {real, imag} */,
  {32'hc0d1a4f9, 32'hc17aca91} /* (30, 3, 18) {real, imag} */,
  {32'hc0696006, 32'hc1803bf0} /* (30, 3, 17) {real, imag} */,
  {32'hbf030670, 32'hc125b570} /* (30, 3, 16) {real, imag} */,
  {32'h3fbcdd00, 32'h410038dc} /* (30, 3, 15) {real, imag} */,
  {32'h3f94120a, 32'h414c3c06} /* (30, 3, 14) {real, imag} */,
  {32'h3fbad72b, 32'h415f1470} /* (30, 3, 13) {real, imag} */,
  {32'h404623d2, 32'h4154a672} /* (30, 3, 12) {real, imag} */,
  {32'h4062228e, 32'h4168e039} /* (30, 3, 11) {real, imag} */,
  {32'h3ffbe354, 32'h41749ff0} /* (30, 3, 10) {real, imag} */,
  {32'h4070880c, 32'h416193f7} /* (30, 3, 9) {real, imag} */,
  {32'h40a311bd, 32'h415c5243} /* (30, 3, 8) {real, imag} */,
  {32'h4040ae40, 32'h41578a6c} /* (30, 3, 7) {real, imag} */,
  {32'h40602a44, 32'h415558db} /* (30, 3, 6) {real, imag} */,
  {32'hbf45ddb6, 32'hc089abd0} /* (30, 3, 5) {real, imag} */,
  {32'h3d904a30, 32'hc15ef3c0} /* (30, 3, 4) {real, imag} */,
  {32'hbf9e2abc, 32'hc17e4387} /* (30, 3, 3) {real, imag} */,
  {32'hbfb17a7b, 32'hc1907018} /* (30, 3, 2) {real, imag} */,
  {32'hc055d48e, 32'hc15b2b54} /* (30, 3, 1) {real, imag} */,
  {32'hbf289ee2, 32'hc0b3dd52} /* (30, 3, 0) {real, imag} */,
  {32'hbf82607a, 32'hc0ff89c0} /* (30, 2, 31) {real, imag} */,
  {32'hc01ab8a3, 32'hc1852ef1} /* (30, 2, 30) {real, imag} */,
  {32'hbfeadd8a, 32'hc180b616} /* (30, 2, 29) {real, imag} */,
  {32'hbf52ed5c, 32'hc172671e} /* (30, 2, 28) {real, imag} */,
  {32'hbf80c270, 32'hc15eb8cb} /* (30, 2, 27) {real, imag} */,
  {32'hc00e4d78, 32'hc153d746} /* (30, 2, 26) {real, imag} */,
  {32'hc0cd6eaa, 32'hc1632b34} /* (30, 2, 25) {real, imag} */,
  {32'hc098f1cd, 32'hc17d3946} /* (30, 2, 24) {real, imag} */,
  {32'hc034ce82, 32'hc1800f8a} /* (30, 2, 23) {real, imag} */,
  {32'hc0480fa2, 32'hc13c795e} /* (30, 2, 22) {real, imag} */,
  {32'hc01d2590, 32'hc13b0f04} /* (30, 2, 21) {real, imag} */,
  {32'hc03c5d51, 32'hc17038ad} /* (30, 2, 20) {real, imag} */,
  {32'hc0c8385f, 32'hc1841b06} /* (30, 2, 19) {real, imag} */,
  {32'hc11c4fba, 32'hc16b6cda} /* (30, 2, 18) {real, imag} */,
  {32'hc0fb8c0c, 32'hc16b0750} /* (30, 2, 17) {real, imag} */,
  {32'hbfd8833b, 32'hc108a8f8} /* (30, 2, 16) {real, imag} */,
  {32'h3f9837ea, 32'h41148f80} /* (30, 2, 15) {real, imag} */,
  {32'h3ff75afc, 32'h414fc892} /* (30, 2, 14) {real, imag} */,
  {32'h407a43d0, 32'h41653e5f} /* (30, 2, 13) {real, imag} */,
  {32'h3fe8f713, 32'h4166c89e} /* (30, 2, 12) {real, imag} */,
  {32'h4083e4b7, 32'h41522277} /* (30, 2, 11) {real, imag} */,
  {32'h4099567e, 32'h415fc42a} /* (30, 2, 10) {real, imag} */,
  {32'h40890d95, 32'h417c8b68} /* (30, 2, 9) {real, imag} */,
  {32'h40b5170a, 32'h41599fac} /* (30, 2, 8) {real, imag} */,
  {32'h4030c3a6, 32'h4151b358} /* (30, 2, 7) {real, imag} */,
  {32'h3fc74f40, 32'h4171c01e} /* (30, 2, 6) {real, imag} */,
  {32'hc02d9c68, 32'hbf99459a} /* (30, 2, 5) {real, imag} */,
  {32'hc040acc4, 32'hc167ed73} /* (30, 2, 4) {real, imag} */,
  {32'hc017a68e, 32'hc17e892b} /* (30, 2, 3) {real, imag} */,
  {32'hc05b05a2, 32'hc188b10a} /* (30, 2, 2) {real, imag} */,
  {32'hc0b5af07, 32'hc170bdc6} /* (30, 2, 1) {real, imag} */,
  {32'hc044c696, 32'hc0c38da2} /* (30, 2, 0) {real, imag} */,
  {32'hc017d2a5, 32'hc0c994e8} /* (30, 1, 31) {real, imag} */,
  {32'hc048b23a, 32'hc13dedc5} /* (30, 1, 30) {real, imag} */,
  {32'hc065dc5b, 32'hc15ee71e} /* (30, 1, 29) {real, imag} */,
  {32'hc02463da, 32'hc1554bf5} /* (30, 1, 28) {real, imag} */,
  {32'hbfc6107b, 32'hc171bd89} /* (30, 1, 27) {real, imag} */,
  {32'hbf6c20d5, 32'hc15ad129} /* (30, 1, 26) {real, imag} */,
  {32'hc08a87fa, 32'hc15adeaa} /* (30, 1, 25) {real, imag} */,
  {32'hc08b522c, 32'hc174b13c} /* (30, 1, 24) {real, imag} */,
  {32'hc008a0f8, 32'hc183c354} /* (30, 1, 23) {real, imag} */,
  {32'hbf684378, 32'hc15020e8} /* (30, 1, 22) {real, imag} */,
  {32'hbf126e63, 32'hc1395606} /* (30, 1, 21) {real, imag} */,
  {32'hc015de9e, 32'hc15fe496} /* (30, 1, 20) {real, imag} */,
  {32'hc0706d43, 32'hc1788ffb} /* (30, 1, 19) {real, imag} */,
  {32'hc10eb30e, 32'hc18da710} /* (30, 1, 18) {real, imag} */,
  {32'hc0a42dfa, 32'hc18a329f} /* (30, 1, 17) {real, imag} */,
  {32'hbfd5a4a8, 32'hc0f3d5f1} /* (30, 1, 16) {real, imag} */,
  {32'h3f4c58e8, 32'h41179a4c} /* (30, 1, 15) {real, imag} */,
  {32'h4017cc2b, 32'h416b9cf8} /* (30, 1, 14) {real, imag} */,
  {32'h40c1755a, 32'h417c8a3b} /* (30, 1, 13) {real, imag} */,
  {32'h40a256b4, 32'h4176052e} /* (30, 1, 12) {real, imag} */,
  {32'h4053fe52, 32'h414fdfed} /* (30, 1, 11) {real, imag} */,
  {32'h40210d5a, 32'h41794304} /* (30, 1, 10) {real, imag} */,
  {32'h40268b5c, 32'h41847a92} /* (30, 1, 9) {real, imag} */,
  {32'h400fd340, 32'h4165bf40} /* (30, 1, 8) {real, imag} */,
  {32'h4041cb22, 32'h417422a4} /* (30, 1, 7) {real, imag} */,
  {32'h401b28e8, 32'h41884e3e} /* (30, 1, 6) {real, imag} */,
  {32'hbf886cee, 32'hbf921506} /* (30, 1, 5) {real, imag} */,
  {32'hc0b5b47e, 32'hc1673e26} /* (30, 1, 4) {real, imag} */,
  {32'hc0889218, 32'hc16fcc1f} /* (30, 1, 3) {real, imag} */,
  {32'hc01646e6, 32'hc15c1128} /* (30, 1, 2) {real, imag} */,
  {32'hc0a594f1, 32'hc14b82df} /* (30, 1, 1) {real, imag} */,
  {32'hc08665e8, 32'hc0d59646} /* (30, 1, 0) {real, imag} */,
  {32'hc01ea9c2, 32'hc05573a2} /* (30, 0, 31) {real, imag} */,
  {32'hc01017e8, 32'hc0b2bdf4} /* (30, 0, 30) {real, imag} */,
  {32'hbfec5a25, 32'hc0ed2504} /* (30, 0, 29) {real, imag} */,
  {32'hbf9c33eb, 32'hc0f6f3e9} /* (30, 0, 28) {real, imag} */,
  {32'hbf8ce83c, 32'hc106f129} /* (30, 0, 27) {real, imag} */,
  {32'h3ef73516, 32'hc10d1a9e} /* (30, 0, 26) {real, imag} */,
  {32'hbfd28671, 32'hc0d6e410} /* (30, 0, 25) {real, imag} */,
  {32'hc03fc071, 32'hc0e20e80} /* (30, 0, 24) {real, imag} */,
  {32'hbfdaa77d, 32'hc11d2d1c} /* (30, 0, 23) {real, imag} */,
  {32'hbff02ee3, 32'hc1013334} /* (30, 0, 22) {real, imag} */,
  {32'hbffb61cc, 32'hc0c2936a} /* (30, 0, 21) {real, imag} */,
  {32'hbfb90842, 32'hc0f8398e} /* (30, 0, 20) {real, imag} */,
  {32'hc00b4cc0, 32'hc10067e1} /* (30, 0, 19) {real, imag} */,
  {32'hc08b0743, 32'hc11d988a} /* (30, 0, 18) {real, imag} */,
  {32'hbf971482, 32'hc117f687} /* (30, 0, 17) {real, imag} */,
  {32'hbec1e074, 32'hc00c2d24} /* (30, 0, 16) {real, imag} */,
  {32'hbd891488, 32'h40c63af6} /* (30, 0, 15) {real, imag} */,
  {32'h3ee15476, 32'h410fc311} /* (30, 0, 14) {real, imag} */,
  {32'h40024147, 32'h41298237} /* (30, 0, 13) {real, imag} */,
  {32'h4061874e, 32'h4111df22} /* (30, 0, 12) {real, imag} */,
  {32'h4051bad4, 32'h410111a5} /* (30, 0, 11) {real, imag} */,
  {32'h3fc0e5b0, 32'h40f09574} /* (30, 0, 10) {real, imag} */,
  {32'h4008a9a3, 32'h40bd340a} /* (30, 0, 9) {real, imag} */,
  {32'h3f304bbe, 32'h40cda0eb} /* (30, 0, 8) {real, imag} */,
  {32'h403a82fe, 32'h410c8e4e} /* (30, 0, 7) {real, imag} */,
  {32'h4046b414, 32'h410e26f4} /* (30, 0, 6) {real, imag} */,
  {32'h3f0bd734, 32'hbfdb67e6} /* (30, 0, 5) {real, imag} */,
  {32'hbfd6a6b1, 32'hc0ebe3c6} /* (30, 0, 4) {real, imag} */,
  {32'hc022fbb1, 32'hc0fb4586} /* (30, 0, 3) {real, imag} */,
  {32'hbf5c161f, 32'hc0d9dc42} /* (30, 0, 2) {real, imag} */,
  {32'hbfdb09f6, 32'hc0ec5f82} /* (30, 0, 1) {real, imag} */,
  {32'hc01e342c, 32'hc0bde6ae} /* (30, 0, 0) {real, imag} */,
  {32'hbf23fc40, 32'h3e9e3f56} /* (29, 31, 31) {real, imag} */,
  {32'hbf986902, 32'h3d7bed00} /* (29, 31, 30) {real, imag} */,
  {32'hbf9489ba, 32'hc023d0f0} /* (29, 31, 29) {real, imag} */,
  {32'hc03c8b61, 32'hc05b652e} /* (29, 31, 28) {real, imag} */,
  {32'hbfe7cba2, 32'hc0703c0d} /* (29, 31, 27) {real, imag} */,
  {32'hbf74ef53, 32'hbffd8d3b} /* (29, 31, 26) {real, imag} */,
  {32'hbf38be58, 32'hc083a241} /* (29, 31, 25) {real, imag} */,
  {32'h3ef0fc4a, 32'hc08e397a} /* (29, 31, 24) {real, imag} */,
  {32'h3f094a32, 32'hc05db876} /* (29, 31, 23) {real, imag} */,
  {32'h3f37bb82, 32'hc0853850} /* (29, 31, 22) {real, imag} */,
  {32'h3f8dfa78, 32'hc03fc80a} /* (29, 31, 21) {real, imag} */,
  {32'h4006992a, 32'h403ad95e} /* (29, 31, 20) {real, imag} */,
  {32'h3e2c0e0f, 32'h40321a18} /* (29, 31, 19) {real, imag} */,
  {32'hbd0d90c0, 32'h3e75d1ec} /* (29, 31, 18) {real, imag} */,
  {32'h3f0cf424, 32'h3d904708} /* (29, 31, 17) {real, imag} */,
  {32'h3fa80d52, 32'h4020ca93} /* (29, 31, 16) {real, imag} */,
  {32'h3f76770f, 32'h4010e2c0} /* (29, 31, 15) {real, imag} */,
  {32'h401901b9, 32'h4086ffb0} /* (29, 31, 14) {real, imag} */,
  {32'h3ec7c43c, 32'h40b4ce6a} /* (29, 31, 13) {real, imag} */,
  {32'h3f0bdd0f, 32'h4096f3d4} /* (29, 31, 12) {real, imag} */,
  {32'h3f2b0a28, 32'h4000717a} /* (29, 31, 11) {real, imag} */,
  {32'h3e1eb758, 32'hc08d694a} /* (29, 31, 10) {real, imag} */,
  {32'h3d319ca0, 32'hc08e51f2} /* (29, 31, 9) {real, imag} */,
  {32'h3edf2d4d, 32'hc0817d77} /* (29, 31, 8) {real, imag} */,
  {32'h3cfb3ac0, 32'hc073c158} /* (29, 31, 7) {real, imag} */,
  {32'hbe696f4e, 32'hc0039ab4} /* (29, 31, 6) {real, imag} */,
  {32'hbf3abd8f, 32'hbf915aba} /* (29, 31, 5) {real, imag} */,
  {32'h3eafefbb, 32'hc02309d5} /* (29, 31, 4) {real, imag} */,
  {32'h3f84013e, 32'hc01e9cc4} /* (29, 31, 3) {real, imag} */,
  {32'hbf5f2439, 32'hc02b9034} /* (29, 31, 2) {real, imag} */,
  {32'hc02cd63c, 32'hc08b170b} /* (29, 31, 1) {real, imag} */,
  {32'hbf064877, 32'hbfa31383} /* (29, 31, 0) {real, imag} */,
  {32'hbfb544ce, 32'hbf0a03d8} /* (29, 30, 31) {real, imag} */,
  {32'hbee7308c, 32'hbfcae33a} /* (29, 30, 30) {real, imag} */,
  {32'hbf5d86be, 32'hc05a15a9} /* (29, 30, 29) {real, imag} */,
  {32'hc0a2ad46, 32'hc0d9177b} /* (29, 30, 28) {real, imag} */,
  {32'hc0571a76, 32'hc0c5f076} /* (29, 30, 27) {real, imag} */,
  {32'hbf294ad3, 32'hc0741462} /* (29, 30, 26) {real, imag} */,
  {32'hc01073da, 32'hc0cc82a0} /* (29, 30, 25) {real, imag} */,
  {32'hbff8cc74, 32'hc0c13f58} /* (29, 30, 24) {real, imag} */,
  {32'hc043d842, 32'hc09bd6d8} /* (29, 30, 23) {real, imag} */,
  {32'hc01c5278, 32'hc0b6761d} /* (29, 30, 22) {real, imag} */,
  {32'h3c8bd518, 32'hc08bbe38} /* (29, 30, 21) {real, imag} */,
  {32'h407a3a1f, 32'h40a2724b} /* (29, 30, 20) {real, imag} */,
  {32'h3fbe7a91, 32'h408deadf} /* (29, 30, 19) {real, imag} */,
  {32'h3f798c5c, 32'h402ec78a} /* (29, 30, 18) {real, imag} */,
  {32'h3fdac6e0, 32'h40560ca5} /* (29, 30, 17) {real, imag} */,
  {32'h40551773, 32'h40b59719} /* (29, 30, 16) {real, imag} */,
  {32'hbece87d9, 32'h408b6ad6} /* (29, 30, 15) {real, imag} */,
  {32'h406b03d7, 32'h409e8dc0} /* (29, 30, 14) {real, imag} */,
  {32'h3f9ddd02, 32'h40db20af} /* (29, 30, 13) {real, imag} */,
  {32'h3f9161e8, 32'h4101e577} /* (29, 30, 12) {real, imag} */,
  {32'h401cc9c0, 32'h40cadcf4} /* (29, 30, 11) {real, imag} */,
  {32'h3f948c3c, 32'hc0696537} /* (29, 30, 10) {real, imag} */,
  {32'h3efb69e8, 32'hc0bb95b0} /* (29, 30, 9) {real, imag} */,
  {32'h3f8754d2, 32'hc0bd9eb8} /* (29, 30, 8) {real, imag} */,
  {32'h3f5b06be, 32'hc0bfb12c} /* (29, 30, 7) {real, imag} */,
  {32'h3eb852ac, 32'hc06f5754} /* (29, 30, 6) {real, imag} */,
  {32'hbf646352, 32'hc093d86f} /* (29, 30, 5) {real, imag} */,
  {32'h3f6cc4df, 32'hc0cd1018} /* (29, 30, 4) {real, imag} */,
  {32'hbf05ecf7, 32'hc0b8dbce} /* (29, 30, 3) {real, imag} */,
  {32'hc000c539, 32'hc0bfc374} /* (29, 30, 2) {real, imag} */,
  {32'hc0612333, 32'hc0b74cf3} /* (29, 30, 1) {real, imag} */,
  {32'hbfea4ead, 32'hbff1631d} /* (29, 30, 0) {real, imag} */,
  {32'hc02def62, 32'hc01d336b} /* (29, 29, 31) {real, imag} */,
  {32'h3eb79030, 32'hc0a5f7f0} /* (29, 29, 30) {real, imag} */,
  {32'h3fc38429, 32'hc0b7ea9c} /* (29, 29, 29) {real, imag} */,
  {32'hc09edc68, 32'hc0af1d68} /* (29, 29, 28) {real, imag} */,
  {32'hc064871a, 32'hc0ad6af9} /* (29, 29, 27) {real, imag} */,
  {32'h3eacc596, 32'hc0c71a10} /* (29, 29, 26) {real, imag} */,
  {32'hbf82a415, 32'hc0f94aee} /* (29, 29, 25) {real, imag} */,
  {32'hbfc57e52, 32'hc0b9e780} /* (29, 29, 24) {real, imag} */,
  {32'hbf5d3aa8, 32'hc0492a25} /* (29, 29, 23) {real, imag} */,
  {32'hbfc5a17d, 32'hc0a7f4f8} /* (29, 29, 22) {real, imag} */,
  {32'hbff68f01, 32'hc08262c3} /* (29, 29, 21) {real, imag} */,
  {32'h403551fc, 32'h40cb400c} /* (29, 29, 20) {real, imag} */,
  {32'h4087edda, 32'h40f6616e} /* (29, 29, 19) {real, imag} */,
  {32'h406cc163, 32'h40b90aa1} /* (29, 29, 18) {real, imag} */,
  {32'h3fba669a, 32'h409d776d} /* (29, 29, 17) {real, imag} */,
  {32'h3ffa4dbe, 32'h4097cfca} /* (29, 29, 16) {real, imag} */,
  {32'hbf8706ae, 32'h40b3faae} /* (29, 29, 15) {real, imag} */,
  {32'h402c73e8, 32'h40c3fef0} /* (29, 29, 14) {real, imag} */,
  {32'h3f68f91b, 32'h4093d4bd} /* (29, 29, 13) {real, imag} */,
  {32'h3f7541cc, 32'h40f24cd8} /* (29, 29, 12) {real, imag} */,
  {32'h3ff78d4b, 32'h40cd30e4} /* (29, 29, 11) {real, imag} */,
  {32'hbf6e20ec, 32'hc03bb69e} /* (29, 29, 10) {real, imag} */,
  {32'hc033defa, 32'hc0ae6c4e} /* (29, 29, 9) {real, imag} */,
  {32'hbfd8b5be, 32'hc0b76ff5} /* (29, 29, 8) {real, imag} */,
  {32'hbefa651c, 32'hc0ae6494} /* (29, 29, 7) {real, imag} */,
  {32'h3b387400, 32'hc01edf16} /* (29, 29, 6) {real, imag} */,
  {32'hc06e3917, 32'hc0431da6} /* (29, 29, 5) {real, imag} */,
  {32'hbfb8470e, 32'hc0c8a480} /* (29, 29, 4) {real, imag} */,
  {32'h3f0bcb7a, 32'hc0f55459} /* (29, 29, 3) {real, imag} */,
  {32'hbf0bd209, 32'hc0de12c5} /* (29, 29, 2) {real, imag} */,
  {32'hbf6b584c, 32'hc0222eec} /* (29, 29, 1) {real, imag} */,
  {32'hbfbc23d4, 32'h3eb79dd4} /* (29, 29, 0) {real, imag} */,
  {32'hbfde23e8, 32'hc07d8172} /* (29, 28, 31) {real, imag} */,
  {32'h3f44b39e, 32'hc0f2f644} /* (29, 28, 30) {real, imag} */,
  {32'h3f0f2800, 32'hc0e6bd12} /* (29, 28, 29) {real, imag} */,
  {32'hc0901b98, 32'hc0309942} /* (29, 28, 28) {real, imag} */,
  {32'hbfaf7cb6, 32'hc0874a9a} /* (29, 28, 27) {real, imag} */,
  {32'h3faa1aec, 32'hc0d8e472} /* (29, 28, 26) {real, imag} */,
  {32'h3f5724f2, 32'hc09828fb} /* (29, 28, 25) {real, imag} */,
  {32'hbf628b81, 32'hc0202446} /* (29, 28, 24) {real, imag} */,
  {32'hbf9efbf2, 32'hc039880a} /* (29, 28, 23) {real, imag} */,
  {32'hc08b3c32, 32'hc0d54f00} /* (29, 28, 22) {real, imag} */,
  {32'hc0c08e16, 32'hc0869d4b} /* (29, 28, 21) {real, imag} */,
  {32'h3fef62e9, 32'h40a59976} /* (29, 28, 20) {real, imag} */,
  {32'h40b8348d, 32'h4108fce5} /* (29, 28, 19) {real, imag} */,
  {32'h40049d60, 32'h40a4f019} /* (29, 28, 18) {real, imag} */,
  {32'h3f45f52a, 32'h404df096} /* (29, 28, 17) {real, imag} */,
  {32'h3fd474ef, 32'h404f392f} /* (29, 28, 16) {real, imag} */,
  {32'h3f851f82, 32'h40a1456c} /* (29, 28, 15) {real, imag} */,
  {32'h3fb2704c, 32'h40c64dac} /* (29, 28, 14) {real, imag} */,
  {32'h3e9965ba, 32'h40ad9486} /* (29, 28, 13) {real, imag} */,
  {32'h3eff8202, 32'h40c0500f} /* (29, 28, 12) {real, imag} */,
  {32'hbe8beb17, 32'h40a1f3dd} /* (29, 28, 11) {real, imag} */,
  {32'hc0a4daf1, 32'hc0834e07} /* (29, 28, 10) {real, imag} */,
  {32'hc0b94788, 32'hc0f1d89a} /* (29, 28, 9) {real, imag} */,
  {32'hc0a4e688, 32'hc10319ca} /* (29, 28, 8) {real, imag} */,
  {32'hc05485d9, 32'hc0f251f5} /* (29, 28, 7) {real, imag} */,
  {32'hbf942c08, 32'hbff2889a} /* (29, 28, 6) {real, imag} */,
  {32'hc07991f3, 32'hc041c93e} /* (29, 28, 5) {real, imag} */,
  {32'hbf70caa1, 32'hc0ea0ae4} /* (29, 28, 4) {real, imag} */,
  {32'h3ede7f90, 32'hc11ed1dc} /* (29, 28, 3) {real, imag} */,
  {32'h3e1ae764, 32'hc0d1891d} /* (29, 28, 2) {real, imag} */,
  {32'h3fe790f2, 32'hc00d925f} /* (29, 28, 1) {real, imag} */,
  {32'hbfc6f680, 32'hbf81d8f0} /* (29, 28, 0) {real, imag} */,
  {32'h3e7515c0, 32'hbffeaeb5} /* (29, 27, 31) {real, imag} */,
  {32'h3f203383, 32'hc0372341} /* (29, 27, 30) {real, imag} */,
  {32'hbeb1a052, 32'hc056a084} /* (29, 27, 29) {real, imag} */,
  {32'hc085e5da, 32'hc0325fd3} /* (29, 27, 28) {real, imag} */,
  {32'hbf95c87f, 32'hc0ddeae0} /* (29, 27, 27) {real, imag} */,
  {32'h3fd567a4, 32'hc1219ab9} /* (29, 27, 26) {real, imag} */,
  {32'h40286f50, 32'hc0cc28ac} /* (29, 27, 25) {real, imag} */,
  {32'h3f1e7969, 32'hc0a17f90} /* (29, 27, 24) {real, imag} */,
  {32'hbf39f02c, 32'hc0840a53} /* (29, 27, 23) {real, imag} */,
  {32'hc026ca4a, 32'hc08fb5f6} /* (29, 27, 22) {real, imag} */,
  {32'hc0af1a89, 32'hc023bc00} /* (29, 27, 21) {real, imag} */,
  {32'hbeb568d8, 32'h40ad9c68} /* (29, 27, 20) {real, imag} */,
  {32'h3faf7631, 32'h4105feac} /* (29, 27, 19) {real, imag} */,
  {32'h3f83720a, 32'h40dfa610} /* (29, 27, 18) {real, imag} */,
  {32'h40184354, 32'h408d83c0} /* (29, 27, 17) {real, imag} */,
  {32'h3f122cae, 32'h40890d88} /* (29, 27, 16) {real, imag} */,
  {32'hbf8bce37, 32'h40559b8f} /* (29, 27, 15) {real, imag} */,
  {32'hbed32a52, 32'h404e5475} /* (29, 27, 14) {real, imag} */,
  {32'h3fe47c68, 32'h40f53bf4} /* (29, 27, 13) {real, imag} */,
  {32'h3fe668ad, 32'h40bde93c} /* (29, 27, 12) {real, imag} */,
  {32'hbf37daff, 32'h409fe602} /* (29, 27, 11) {real, imag} */,
  {32'hc05d752e, 32'hc065fd16} /* (29, 27, 10) {real, imag} */,
  {32'hc01ec614, 32'hc1000dfa} /* (29, 27, 9) {real, imag} */,
  {32'hc06e4d5e, 32'hc0c0a397} /* (29, 27, 8) {real, imag} */,
  {32'hc01be1e9, 32'hc0c1d964} /* (29, 27, 7) {real, imag} */,
  {32'hbfdd9e1a, 32'hc008d24a} /* (29, 27, 6) {real, imag} */,
  {32'hc07a72ed, 32'hc091dd0a} /* (29, 27, 5) {real, imag} */,
  {32'hbd046d78, 32'hc1036f99} /* (29, 27, 4) {real, imag} */,
  {32'hbf768735, 32'hc11ef222} /* (29, 27, 3) {real, imag} */,
  {32'hc01a895e, 32'hc0d645ae} /* (29, 27, 2) {real, imag} */,
  {32'h3f22de14, 32'hc066f10e} /* (29, 27, 1) {real, imag} */,
  {32'h3e9bf91b, 32'hc018a690} /* (29, 27, 0) {real, imag} */,
  {32'hbceb5dd0, 32'hc00457b9} /* (29, 26, 31) {real, imag} */,
  {32'h3dc4dc20, 32'hc05ebd8d} /* (29, 26, 30) {real, imag} */,
  {32'h3cf4c940, 32'hc0c8cb48} /* (29, 26, 29) {real, imag} */,
  {32'hc01d38c2, 32'hc08f6f5c} /* (29, 26, 28) {real, imag} */,
  {32'hc00f8aa4, 32'hc0ce955a} /* (29, 26, 27) {real, imag} */,
  {32'hbfccb0e0, 32'hc0fc4f95} /* (29, 26, 26) {real, imag} */,
  {32'h3ffdc514, 32'hc0b2aae2} /* (29, 26, 25) {real, imag} */,
  {32'h3f43085e, 32'hc1021434} /* (29, 26, 24) {real, imag} */,
  {32'hc02c0808, 32'hc0a9b795} /* (29, 26, 23) {real, imag} */,
  {32'hc0343645, 32'hc0578528} /* (29, 26, 22) {real, imag} */,
  {32'hbfd25ef6, 32'hbfd1bad5} /* (29, 26, 21) {real, imag} */,
  {32'h3f908fe6, 32'h40c8b6b0} /* (29, 26, 20) {real, imag} */,
  {32'h40199b31, 32'h40e15986} /* (29, 26, 19) {real, imag} */,
  {32'h4081173d, 32'h40d9e55a} /* (29, 26, 18) {real, imag} */,
  {32'h408616ed, 32'h40bdf192} /* (29, 26, 17) {real, imag} */,
  {32'h3e0b9268, 32'h4090789e} /* (29, 26, 16) {real, imag} */,
  {32'hbfac4c58, 32'h40a81742} /* (29, 26, 15) {real, imag} */,
  {32'h3f93c0f1, 32'h409652df} /* (29, 26, 14) {real, imag} */,
  {32'h406a1186, 32'h40845b7a} /* (29, 26, 13) {real, imag} */,
  {32'h40612a9b, 32'h40672fe2} /* (29, 26, 12) {real, imag} */,
  {32'h4046d639, 32'h403d0f46} /* (29, 26, 11) {real, imag} */,
  {32'hbf178a45, 32'hbfaa64f0} /* (29, 26, 10) {real, imag} */,
  {32'hc0219b78, 32'hc0ed009f} /* (29, 26, 9) {real, imag} */,
  {32'hbf6a3b5a, 32'hc0597766} /* (29, 26, 8) {real, imag} */,
  {32'hbef6141c, 32'hbfe9268a} /* (29, 26, 7) {real, imag} */,
  {32'hbfde61f7, 32'hbff90f3e} /* (29, 26, 6) {real, imag} */,
  {32'hbf620598, 32'hc049275a} /* (29, 26, 5) {real, imag} */,
  {32'hbf67a844, 32'hc0956d2a} /* (29, 26, 4) {real, imag} */,
  {32'hbfdc7822, 32'hc09c3c6f} /* (29, 26, 3) {real, imag} */,
  {32'hbf3d4e36, 32'hc08bb40f} /* (29, 26, 2) {real, imag} */,
  {32'hbf2aa87c, 32'hc04c6ad2} /* (29, 26, 1) {real, imag} */,
  {32'h3eeabc78, 32'hc0182784} /* (29, 26, 0) {real, imag} */,
  {32'hbfaf1b18, 32'hc07d9958} /* (29, 25, 31) {real, imag} */,
  {32'hbf3eda1c, 32'hc0ea79e0} /* (29, 25, 30) {real, imag} */,
  {32'hbe50191c, 32'hc0d56060} /* (29, 25, 29) {real, imag} */,
  {32'hbcd91310, 32'hc09d67ce} /* (29, 25, 28) {real, imag} */,
  {32'hc007c7da, 32'hc09bb400} /* (29, 25, 27) {real, imag} */,
  {32'hc003e261, 32'hc0c410a1} /* (29, 25, 26) {real, imag} */,
  {32'h3ffc8561, 32'hc0ca16a4} /* (29, 25, 25) {real, imag} */,
  {32'h3e3d7fa8, 32'hc0d7a09d} /* (29, 25, 24) {real, imag} */,
  {32'hc0458c02, 32'hc0a85d4b} /* (29, 25, 23) {real, imag} */,
  {32'hc0326a71, 32'hc0563d19} /* (29, 25, 22) {real, imag} */,
  {32'hbfc55014, 32'h3fcbc695} /* (29, 25, 21) {real, imag} */,
  {32'hbf4df390, 32'h40d2f698} /* (29, 25, 20) {real, imag} */,
  {32'h3fed69ac, 32'h4092dd1a} /* (29, 25, 19) {real, imag} */,
  {32'h4080ec14, 32'h40be22f5} /* (29, 25, 18) {real, imag} */,
  {32'hbf2732c2, 32'h40c11eda} /* (29, 25, 17) {real, imag} */,
  {32'hbf97bebe, 32'h4073f4ec} /* (29, 25, 16) {real, imag} */,
  {32'h40201f26, 32'h40eb703e} /* (29, 25, 15) {real, imag} */,
  {32'h40a32925, 32'h411ee4d0} /* (29, 25, 14) {real, imag} */,
  {32'h3feb7421, 32'h401dc00c} /* (29, 25, 13) {real, imag} */,
  {32'h3f72cb7d, 32'h3fcbd431} /* (29, 25, 12) {real, imag} */,
  {32'h3dea0cf5, 32'h40306052} /* (29, 25, 11) {real, imag} */,
  {32'hbfc5b5c0, 32'hc013c836} /* (29, 25, 10) {real, imag} */,
  {32'hc04b058a, 32'hc0d3851c} /* (29, 25, 9) {real, imag} */,
  {32'hc04a840c, 32'hc0b052f4} /* (29, 25, 8) {real, imag} */,
  {32'hbff3f80a, 32'hc0929998} /* (29, 25, 7) {real, imag} */,
  {32'hbfdc859a, 32'hc0a36bbe} /* (29, 25, 6) {real, imag} */,
  {32'h3e8d8eea, 32'hc0f9ec00} /* (29, 25, 5) {real, imag} */,
  {32'h3e99b21c, 32'hc0fe0274} /* (29, 25, 4) {real, imag} */,
  {32'h3edb95f5, 32'hc0946513} /* (29, 25, 3) {real, imag} */,
  {32'h3f0c61bc, 32'hc02cebf0} /* (29, 25, 2) {real, imag} */,
  {32'hbfb568c6, 32'hbf107271} /* (29, 25, 1) {real, imag} */,
  {32'hbf407f32, 32'hc0259504} /* (29, 25, 0) {real, imag} */,
  {32'hbecfa7da, 32'hc06b466e} /* (29, 24, 31) {real, imag} */,
  {32'hbf84d274, 32'hc10d8ece} /* (29, 24, 30) {real, imag} */,
  {32'h3e08c794, 32'hc0a8356b} /* (29, 24, 29) {real, imag} */,
  {32'h3ef19bc0, 32'hc0a679d4} /* (29, 24, 28) {real, imag} */,
  {32'hc0148564, 32'hc0bb1b7e} /* (29, 24, 27) {real, imag} */,
  {32'h3e163950, 32'hc0fe03d0} /* (29, 24, 26) {real, imag} */,
  {32'h3fa38c62, 32'hc1117cb7} /* (29, 24, 25) {real, imag} */,
  {32'hbffe1d74, 32'hc06ce2ab} /* (29, 24, 24) {real, imag} */,
  {32'hc083eecb, 32'hc07e125a} /* (29, 24, 23) {real, imag} */,
  {32'hc0318fee, 32'hc0802488} /* (29, 24, 22) {real, imag} */,
  {32'hc059f07f, 32'hbec92274} /* (29, 24, 21) {real, imag} */,
  {32'hc03d11fe, 32'h409ed97c} /* (29, 24, 20) {real, imag} */,
  {32'h3f3c392d, 32'h4099d75a} /* (29, 24, 19) {real, imag} */,
  {32'h40293788, 32'h40bea5ea} /* (29, 24, 18) {real, imag} */,
  {32'hbed1ddac, 32'h408c15cc} /* (29, 24, 17) {real, imag} */,
  {32'h4041cd07, 32'h40774f7c} /* (29, 24, 16) {real, imag} */,
  {32'h409e5f72, 32'h40fc1686} /* (29, 24, 15) {real, imag} */,
  {32'h40c1a9c1, 32'h411e1afe} /* (29, 24, 14) {real, imag} */,
  {32'h3f65d0cc, 32'h40601c00} /* (29, 24, 13) {real, imag} */,
  {32'hbeaf6ac8, 32'h3fcf5082} /* (29, 24, 12) {real, imag} */,
  {32'h3ef0458a, 32'h3f98d3b2} /* (29, 24, 11) {real, imag} */,
  {32'h3f075db3, 32'hc0a18718} /* (29, 24, 10) {real, imag} */,
  {32'hbf1c25bb, 32'hc0bdd440} /* (29, 24, 9) {real, imag} */,
  {32'hc08c2a00, 32'hc0ac2238} /* (29, 24, 8) {real, imag} */,
  {32'hbff4186e, 32'hc0c750fa} /* (29, 24, 7) {real, imag} */,
  {32'hbfb07c76, 32'hc0dbc094} /* (29, 24, 6) {real, imag} */,
  {32'h3c1ba2c0, 32'hc0e97b70} /* (29, 24, 5) {real, imag} */,
  {32'h3f3874e0, 32'hc09d7ad9} /* (29, 24, 4) {real, imag} */,
  {32'h3ef25373, 32'hc0d4302c} /* (29, 24, 3) {real, imag} */,
  {32'h3ffc1394, 32'hc0e82fdf} /* (29, 24, 2) {real, imag} */,
  {32'h3f02eb5a, 32'hc081d758} /* (29, 24, 1) {real, imag} */,
  {32'h3ebf2cda, 32'hc03add63} /* (29, 24, 0) {real, imag} */,
  {32'hbf69442f, 32'hc08132f6} /* (29, 23, 31) {real, imag} */,
  {32'hc030dce4, 32'hc0c4ecd6} /* (29, 23, 30) {real, imag} */,
  {32'hbfcaaf24, 32'hc0bd589c} /* (29, 23, 29) {real, imag} */,
  {32'hbf22389d, 32'hc0a69e34} /* (29, 23, 28) {real, imag} */,
  {32'hc04413cf, 32'hc1070e10} /* (29, 23, 27) {real, imag} */,
  {32'hbfaada2a, 32'hc10c4b3c} /* (29, 23, 26) {real, imag} */,
  {32'hbd93c438, 32'hc0db12a7} /* (29, 23, 25) {real, imag} */,
  {32'hbfd6898c, 32'hc0085fd0} /* (29, 23, 24) {real, imag} */,
  {32'hc005dcba, 32'hc083cca2} /* (29, 23, 23) {real, imag} */,
  {32'hc006e09c, 32'hc0a25fc1} /* (29, 23, 22) {real, imag} */,
  {32'hc063a0e8, 32'hbfd41efe} /* (29, 23, 21) {real, imag} */,
  {32'hc022e8de, 32'h40750465} /* (29, 23, 20) {real, imag} */,
  {32'hbf01dd62, 32'h40b54a40} /* (29, 23, 19) {real, imag} */,
  {32'hbf005f81, 32'h40cccd82} /* (29, 23, 18) {real, imag} */,
  {32'hbe480b5c, 32'h40aa0abe} /* (29, 23, 17) {real, imag} */,
  {32'h4032d2fc, 32'h4004819a} /* (29, 23, 16) {real, imag} */,
  {32'h3d8b6708, 32'h408d148e} /* (29, 23, 15) {real, imag} */,
  {32'h3fb63798, 32'h40fe4697} /* (29, 23, 14) {real, imag} */,
  {32'h3fb63d7a, 32'h4079dbd4} /* (29, 23, 13) {real, imag} */,
  {32'h401de69e, 32'h3fc44fba} /* (29, 23, 12) {real, imag} */,
  {32'h3f568fc0, 32'h406e2ee9} /* (29, 23, 11) {real, imag} */,
  {32'hbe06b5ee, 32'hbfc7fd36} /* (29, 23, 10) {real, imag} */,
  {32'h3fe89e28, 32'hc0b151ac} /* (29, 23, 9) {real, imag} */,
  {32'hbfefe5e8, 32'hc0cdc9a5} /* (29, 23, 8) {real, imag} */,
  {32'hc0137507, 32'hc0fcf237} /* (29, 23, 7) {real, imag} */,
  {32'h3f30e700, 32'hc0bb2d28} /* (29, 23, 6) {real, imag} */,
  {32'hbed9377a, 32'hc0a8e7a5} /* (29, 23, 5) {real, imag} */,
  {32'hbf6c3daa, 32'hc0838c8a} /* (29, 23, 4) {real, imag} */,
  {32'h3ed46497, 32'hc0c5bb74} /* (29, 23, 3) {real, imag} */,
  {32'h401e4263, 32'hc0ce9a8c} /* (29, 23, 2) {real, imag} */,
  {32'h40082e3b, 32'hc0c8ed6f} /* (29, 23, 1) {real, imag} */,
  {32'h3fc12d42, 32'hc08f58a4} /* (29, 23, 0) {real, imag} */,
  {32'hbf60637c, 32'hc013a220} /* (29, 22, 31) {real, imag} */,
  {32'hbf2b9c69, 32'hc082ccc8} /* (29, 22, 30) {real, imag} */,
  {32'hbff8a947, 32'hc0bef31b} /* (29, 22, 29) {real, imag} */,
  {32'hc05b74e0, 32'hc0742bb2} /* (29, 22, 28) {real, imag} */,
  {32'hc0a66d03, 32'hc0b3e254} /* (29, 22, 27) {real, imag} */,
  {32'hc006bc85, 32'hc0c0e5b2} /* (29, 22, 26) {real, imag} */,
  {32'hbde416b8, 32'hc0bd3c61} /* (29, 22, 25) {real, imag} */,
  {32'h3e6be200, 32'hc0add610} /* (29, 22, 24) {real, imag} */,
  {32'h3ea35d9f, 32'hc0b853b7} /* (29, 22, 23) {real, imag} */,
  {32'hbf201a46, 32'hc099e864} /* (29, 22, 22) {real, imag} */,
  {32'hbf19cc94, 32'hc07dc18a} /* (29, 22, 21) {real, imag} */,
  {32'hbe249e96, 32'h407c17ce} /* (29, 22, 20) {real, imag} */,
  {32'hbf93f0e0, 32'h40e59640} /* (29, 22, 19) {real, imag} */,
  {32'hc0136e42, 32'h40bc1b2e} /* (29, 22, 18) {real, imag} */,
  {32'hbfc94d88, 32'h4081d5f2} /* (29, 22, 17) {real, imag} */,
  {32'h3ffdad48, 32'h403d4d4e} /* (29, 22, 16) {real, imag} */,
  {32'h3eda28df, 32'h406d4526} /* (29, 22, 15) {real, imag} */,
  {32'hbf00d638, 32'h40ee6f89} /* (29, 22, 14) {real, imag} */,
  {32'h40011dfe, 32'h40c854c8} /* (29, 22, 13) {real, imag} */,
  {32'h404f3072, 32'h403cdc2e} /* (29, 22, 12) {real, imag} */,
  {32'h3ea74c55, 32'h3fd8564e} /* (29, 22, 11) {real, imag} */,
  {32'hbfe446b9, 32'hc03c29e0} /* (29, 22, 10) {real, imag} */,
  {32'h3eaf3140, 32'hc08af502} /* (29, 22, 9) {real, imag} */,
  {32'hbff8f87a, 32'hc07e2c2a} /* (29, 22, 8) {real, imag} */,
  {32'hc0215e9e, 32'hc0b8bb97} /* (29, 22, 7) {real, imag} */,
  {32'hbf7b5874, 32'hc0b7d416} /* (29, 22, 6) {real, imag} */,
  {32'hbf999740, 32'hc0e511f6} /* (29, 22, 5) {real, imag} */,
  {32'hbf8d275e, 32'hc0a8b746} /* (29, 22, 4) {real, imag} */,
  {32'hbecbcee4, 32'hc0f68bfe} /* (29, 22, 3) {real, imag} */,
  {32'h3ffdb84e, 32'hc0a9abae} /* (29, 22, 2) {real, imag} */,
  {32'h3eabb3f5, 32'hc0195e2a} /* (29, 22, 1) {real, imag} */,
  {32'hbd8a282e, 32'hc0196510} /* (29, 22, 0) {real, imag} */,
  {32'hbf638c8f, 32'hbe9c2771} /* (29, 21, 31) {real, imag} */,
  {32'hbec2c233, 32'hbf2102f0} /* (29, 21, 30) {real, imag} */,
  {32'hbe0623f0, 32'hbfac584d} /* (29, 21, 29) {real, imag} */,
  {32'hc0134002, 32'hc00e4c96} /* (29, 21, 28) {real, imag} */,
  {32'hbf801725, 32'hc0218ee3} /* (29, 21, 27) {real, imag} */,
  {32'h40236db2, 32'hbfd5f0b8} /* (29, 21, 26) {real, imag} */,
  {32'h3fa2c210, 32'hc0045f50} /* (29, 21, 25) {real, imag} */,
  {32'hbe1f9e4c, 32'hbf7f50ae} /* (29, 21, 24) {real, imag} */,
  {32'hbd4350d4, 32'hbfa42e6c} /* (29, 21, 23) {real, imag} */,
  {32'hbf351d7b, 32'h3ee3a63a} /* (29, 21, 22) {real, imag} */,
  {32'h3e7a7991, 32'hc007db9d} /* (29, 21, 21) {real, imag} */,
  {32'hbff667ef, 32'h40288880} /* (29, 21, 20) {real, imag} */,
  {32'hc07c1d8a, 32'h40599368} /* (29, 21, 19) {real, imag} */,
  {32'hc002a86d, 32'h404aac98} /* (29, 21, 18) {real, imag} */,
  {32'hc0019fb6, 32'h4061f3c4} /* (29, 21, 17) {real, imag} */,
  {32'h3feb3220, 32'h40493bda} /* (29, 21, 16) {real, imag} */,
  {32'h3f8a307c, 32'h400c5a8c} /* (29, 21, 15) {real, imag} */,
  {32'hbf4d894e, 32'h408d7af2} /* (29, 21, 14) {real, imag} */,
  {32'h3fd7f5cd, 32'h40379ba7} /* (29, 21, 13) {real, imag} */,
  {32'h4079c864, 32'h3fbcdeae} /* (29, 21, 12) {real, imag} */,
  {32'h3f9468ab, 32'hbeb4e695} /* (29, 21, 11) {real, imag} */,
  {32'hc04a70d0, 32'hc02c9dea} /* (29, 21, 10) {real, imag} */,
  {32'h3e7972c2, 32'hbff3c444} /* (29, 21, 9) {real, imag} */,
  {32'h3e30d28c, 32'hbf5e4f79} /* (29, 21, 8) {real, imag} */,
  {32'hc021b1e4, 32'hbf4bcb25} /* (29, 21, 7) {real, imag} */,
  {32'hc018c56b, 32'hbfae4ed4} /* (29, 21, 6) {real, imag} */,
  {32'hbee90c91, 32'hc035d740} /* (29, 21, 5) {real, imag} */,
  {32'hbe9c9d84, 32'hc0357de7} /* (29, 21, 4) {real, imag} */,
  {32'h3ee258f9, 32'hc08b5126} /* (29, 21, 3) {real, imag} */,
  {32'h3f17bece, 32'hc00ec0c6} /* (29, 21, 2) {real, imag} */,
  {32'hc0091ee3, 32'hbddc529c} /* (29, 21, 1) {real, imag} */,
  {32'hc0057da2, 32'hbe367b26} /* (29, 21, 0) {real, imag} */,
  {32'hbf14b2bc, 32'h402d7bdc} /* (29, 20, 31) {real, imag} */,
  {32'hbfcf166a, 32'h40a373ea} /* (29, 20, 30) {real, imag} */,
  {32'h402447a6, 32'h40c433ce} /* (29, 20, 29) {real, imag} */,
  {32'h40235fdc, 32'h40646992} /* (29, 20, 28) {real, imag} */,
  {32'h40926ac2, 32'h4063a1f6} /* (29, 20, 27) {real, imag} */,
  {32'h409a51cd, 32'h40aff5ec} /* (29, 20, 26) {real, imag} */,
  {32'h40a8f873, 32'h40f91b59} /* (29, 20, 25) {real, imag} */,
  {32'h3f762dd8, 32'h41158cc2} /* (29, 20, 24) {real, imag} */,
  {32'hbf824351, 32'h40f9b904} /* (29, 20, 23) {real, imag} */,
  {32'h3e11132e, 32'h40a5687a} /* (29, 20, 22) {real, imag} */,
  {32'hbd5b9b20, 32'h3fff5a47} /* (29, 20, 21) {real, imag} */,
  {32'hbfd41847, 32'hc043f9aa} /* (29, 20, 20) {real, imag} */,
  {32'hc0901cb9, 32'hc08862ce} /* (29, 20, 19) {real, imag} */,
  {32'hc09c67d9, 32'hc04efeb6} /* (29, 20, 18) {real, imag} */,
  {32'hc09a26d6, 32'hc06cfeb0} /* (29, 20, 17) {real, imag} */,
  {32'hc0037637, 32'hc04aa1a1} /* (29, 20, 16) {real, imag} */,
  {32'hbfe1d432, 32'hc064f980} /* (29, 20, 15) {real, imag} */,
  {32'hbfe89bc0, 32'hc07007aa} /* (29, 20, 14) {real, imag} */,
  {32'hbea523e7, 32'hc0ab1c44} /* (29, 20, 13) {real, imag} */,
  {32'h40212432, 32'hc035a3cd} /* (29, 20, 12) {real, imag} */,
  {32'hbe8c20ce, 32'hbf0fc6ee} /* (29, 20, 11) {real, imag} */,
  {32'hc00e02f1, 32'h3e0a5984} /* (29, 20, 10) {real, imag} */,
  {32'h3ec845bf, 32'h4052377f} /* (29, 20, 9) {real, imag} */,
  {32'hbde4a018, 32'h409842e3} /* (29, 20, 8) {real, imag} */,
  {32'hbfcbb702, 32'h40bb399e} /* (29, 20, 7) {real, imag} */,
  {32'h3c967a40, 32'h40d0f33c} /* (29, 20, 6) {real, imag} */,
  {32'h3fa78757, 32'h40a2da33} /* (29, 20, 5) {real, imag} */,
  {32'h4010469a, 32'h40c3c12b} /* (29, 20, 4) {real, imag} */,
  {32'h40278782, 32'h40979f28} /* (29, 20, 3) {real, imag} */,
  {32'h3fda2fe3, 32'h404c49be} /* (29, 20, 2) {real, imag} */,
  {32'hbfcef41c, 32'h408c92a8} /* (29, 20, 1) {real, imag} */,
  {32'hbfe6505b, 32'h3f8f4962} /* (29, 20, 0) {real, imag} */,
  {32'h3f2be11c, 32'h40b182bc} /* (29, 19, 31) {real, imag} */,
  {32'hbfca5dfe, 32'h40c0d088} /* (29, 19, 30) {real, imag} */,
  {32'h3fde29d7, 32'h4079b290} /* (29, 19, 29) {real, imag} */,
  {32'h3ffeb5a3, 32'h4087e267} /* (29, 19, 28) {real, imag} */,
  {32'h40956758, 32'h4086d96a} /* (29, 19, 27) {real, imag} */,
  {32'h40041548, 32'h40bba6a6} /* (29, 19, 26) {real, imag} */,
  {32'h40541987, 32'h40d1ddaa} /* (29, 19, 25) {real, imag} */,
  {32'h40372f08, 32'h40c1e542} /* (29, 19, 24) {real, imag} */,
  {32'h3fe0b42c, 32'h40d7632e} /* (29, 19, 23) {real, imag} */,
  {32'h3f694bb1, 32'h40e38736} /* (29, 19, 22) {real, imag} */,
  {32'hbf83d3e1, 32'h40183be2} /* (29, 19, 21) {real, imag} */,
  {32'hbf3ef815, 32'hc08ca3ea} /* (29, 19, 20) {real, imag} */,
  {32'hbff7b877, 32'hc06d5010} /* (29, 19, 19) {real, imag} */,
  {32'hc0806fa6, 32'hc0a6b9fc} /* (29, 19, 18) {real, imag} */,
  {32'hc0715701, 32'hc0e0334a} /* (29, 19, 17) {real, imag} */,
  {32'hc0385063, 32'hc08e93c4} /* (29, 19, 16) {real, imag} */,
  {32'hbf9e94b0, 32'hc05c283e} /* (29, 19, 15) {real, imag} */,
  {32'hc01936b4, 32'hc0b7712d} /* (29, 19, 14) {real, imag} */,
  {32'hc087197e, 32'hc0fd2aae} /* (29, 19, 13) {real, imag} */,
  {32'hc01434d1, 32'hc0c38558} /* (29, 19, 12) {real, imag} */,
  {32'hbf4de5db, 32'hc039efd4} /* (29, 19, 11) {real, imag} */,
  {32'hc020fc66, 32'h404c437c} /* (29, 19, 10) {real, imag} */,
  {32'hc040649e, 32'h40c59909} /* (29, 19, 9) {real, imag} */,
  {32'hbf777267, 32'h41011f99} /* (29, 19, 8) {real, imag} */,
  {32'hbf859eb4, 32'h40d58af7} /* (29, 19, 7) {real, imag} */,
  {32'h3f3050bc, 32'h40b8972e} /* (29, 19, 6) {real, imag} */,
  {32'h3fad9290, 32'h40d64199} /* (29, 19, 5) {real, imag} */,
  {32'h400eafd9, 32'h40d0dd1b} /* (29, 19, 4) {real, imag} */,
  {32'h4053f36a, 32'h40cc6d56} /* (29, 19, 3) {real, imag} */,
  {32'h404d1b97, 32'h40964aaf} /* (29, 19, 2) {real, imag} */,
  {32'hbead93a2, 32'h4096c350} /* (29, 19, 1) {real, imag} */,
  {32'h3e6db6f6, 32'h40088f29} /* (29, 19, 0) {real, imag} */,
  {32'hbfa291cf, 32'h40cdc03e} /* (29, 18, 31) {real, imag} */,
  {32'hbe3d9f90, 32'h40e2ea12} /* (29, 18, 30) {real, imag} */,
  {32'h3f28ac68, 32'h407408a4} /* (29, 18, 29) {real, imag} */,
  {32'hbf0f346c, 32'h40984229} /* (29, 18, 28) {real, imag} */,
  {32'h40052839, 32'h40b468fe} /* (29, 18, 27) {real, imag} */,
  {32'h3faf4a5e, 32'h40bb6a34} /* (29, 18, 26) {real, imag} */,
  {32'h4042e15a, 32'h408d321b} /* (29, 18, 25) {real, imag} */,
  {32'h403565d8, 32'h409d934e} /* (29, 18, 24) {real, imag} */,
  {32'h403a854e, 32'h408a5c54} /* (29, 18, 23) {real, imag} */,
  {32'h40039e74, 32'h40a301e7} /* (29, 18, 22) {real, imag} */,
  {32'hbfc30d8f, 32'h4009ce51} /* (29, 18, 21) {real, imag} */,
  {32'h3ee1c54a, 32'hc0d7f2e8} /* (29, 18, 20) {real, imag} */,
  {32'hbfa50815, 32'hc0ab65fe} /* (29, 18, 19) {real, imag} */,
  {32'hc09ca92f, 32'hc0aee8a7} /* (29, 18, 18) {real, imag} */,
  {32'hc089188e, 32'hc0c80b48} /* (29, 18, 17) {real, imag} */,
  {32'hc07dabda, 32'hc0564dd3} /* (29, 18, 16) {real, imag} */,
  {32'hc012a05b, 32'hc0a353ba} /* (29, 18, 15) {real, imag} */,
  {32'hc042b0aa, 32'hc105da74} /* (29, 18, 14) {real, imag} */,
  {32'hc03b30aa, 32'hc106b9a8} /* (29, 18, 13) {real, imag} */,
  {32'hc0015ce6, 32'hc0e3b5d5} /* (29, 18, 12) {real, imag} */,
  {32'hbf47dcf2, 32'hc09258f6} /* (29, 18, 11) {real, imag} */,
  {32'hc026fcc2, 32'h40278d26} /* (29, 18, 10) {real, imag} */,
  {32'hc0344b7f, 32'h40bafd5c} /* (29, 18, 9) {real, imag} */,
  {32'h3f01c9e9, 32'h40e2f7e0} /* (29, 18, 8) {real, imag} */,
  {32'h3f1e3130, 32'h40de18ac} /* (29, 18, 7) {real, imag} */,
  {32'h3fa2f134, 32'h40901cc7} /* (29, 18, 6) {real, imag} */,
  {32'h3fe321b8, 32'h40669469} /* (29, 18, 5) {real, imag} */,
  {32'h3f28383c, 32'h4088e7d4} /* (29, 18, 4) {real, imag} */,
  {32'h3fd89e92, 32'h40c03108} /* (29, 18, 3) {real, imag} */,
  {32'h3f790fa4, 32'h40c406ae} /* (29, 18, 2) {real, imag} */,
  {32'h3e83e67c, 32'h40a12cf4} /* (29, 18, 1) {real, imag} */,
  {32'h3fbc0a6c, 32'h401c9cea} /* (29, 18, 0) {real, imag} */,
  {32'h3f23b8bc, 32'h40dd3ca5} /* (29, 17, 31) {real, imag} */,
  {32'h4018d5e6, 32'h411ccde4} /* (29, 17, 30) {real, imag} */,
  {32'h400efc42, 32'h40c2cf16} /* (29, 17, 29) {real, imag} */,
  {32'h3f205307, 32'h40bb637f} /* (29, 17, 28) {real, imag} */,
  {32'h3fa5de4f, 32'h40a774ca} /* (29, 17, 27) {real, imag} */,
  {32'h3f6715d2, 32'h409de2e4} /* (29, 17, 26) {real, imag} */,
  {32'h4087c0a6, 32'h40b9c3a2} /* (29, 17, 25) {real, imag} */,
  {32'h4009c262, 32'h40cf8898} /* (29, 17, 24) {real, imag} */,
  {32'h4018cc7c, 32'h40b83e3c} /* (29, 17, 23) {real, imag} */,
  {32'h3fab1069, 32'h4070b69e} /* (29, 17, 22) {real, imag} */,
  {32'hbf53dc68, 32'h401b20cb} /* (29, 17, 21) {real, imag} */,
  {32'h3fd670fe, 32'hc0a16e69} /* (29, 17, 20) {real, imag} */,
  {32'hbfb10ae3, 32'hc07d69be} /* (29, 17, 19) {real, imag} */,
  {32'hc090db56, 32'hc092231a} /* (29, 17, 18) {real, imag} */,
  {32'hc09dcecf, 32'hc0eeddca} /* (29, 17, 17) {real, imag} */,
  {32'hc040d146, 32'hc06d50ce} /* (29, 17, 16) {real, imag} */,
  {32'hbffbc713, 32'hc0a52148} /* (29, 17, 15) {real, imag} */,
  {32'hbfa54d35, 32'hc105e5c0} /* (29, 17, 14) {real, imag} */,
  {32'hbecb3b8c, 32'hc0dcba60} /* (29, 17, 13) {real, imag} */,
  {32'hbfab47ac, 32'hc094aec1} /* (29, 17, 12) {real, imag} */,
  {32'hbf973e32, 32'hc09df11e} /* (29, 17, 11) {real, imag} */,
  {32'hc065c9da, 32'hbe482854} /* (29, 17, 10) {real, imag} */,
  {32'hbf9ad68e, 32'h408ed0d2} /* (29, 17, 9) {real, imag} */,
  {32'hbfa47677, 32'h4098691e} /* (29, 17, 8) {real, imag} */,
  {32'h3e1e1b8e, 32'h40aabaee} /* (29, 17, 7) {real, imag} */,
  {32'h403a25b4, 32'h40bce1b4} /* (29, 17, 6) {real, imag} */,
  {32'h4035454b, 32'h403ba606} /* (29, 17, 5) {real, imag} */,
  {32'h3ed19a60, 32'h406b00d3} /* (29, 17, 4) {real, imag} */,
  {32'hc004a79a, 32'h40ded42d} /* (29, 17, 3) {real, imag} */,
  {32'h3f034cf4, 32'h40b4cff5} /* (29, 17, 2) {real, imag} */,
  {32'h4029dc37, 32'h4066eef5} /* (29, 17, 1) {real, imag} */,
  {32'h3f737831, 32'h402d1a14} /* (29, 17, 0) {real, imag} */,
  {32'h3f867462, 32'h408ab702} /* (29, 16, 31) {real, imag} */,
  {32'h403a6aaa, 32'h4115bd52} /* (29, 16, 30) {real, imag} */,
  {32'h40054f77, 32'h40bd5767} /* (29, 16, 29) {real, imag} */,
  {32'hbea2741c, 32'h40936682} /* (29, 16, 28) {real, imag} */,
  {32'h3fac9137, 32'h3fdf44e5} /* (29, 16, 27) {real, imag} */,
  {32'h3ff72225, 32'h3f899d8e} /* (29, 16, 26) {real, imag} */,
  {32'h409205e2, 32'h409d0b40} /* (29, 16, 25) {real, imag} */,
  {32'h3f937ac8, 32'h409148c0} /* (29, 16, 24) {real, imag} */,
  {32'h3f3524fd, 32'h40a45d7a} /* (29, 16, 23) {real, imag} */,
  {32'h405848dc, 32'h409180de} /* (29, 16, 22) {real, imag} */,
  {32'h3f22b54b, 32'h400f2258} /* (29, 16, 21) {real, imag} */,
  {32'hbfe44120, 32'hc065ae04} /* (29, 16, 20) {real, imag} */,
  {32'hbfd5a360, 32'hc08e5d4e} /* (29, 16, 19) {real, imag} */,
  {32'hc0262495, 32'hc073c0de} /* (29, 16, 18) {real, imag} */,
  {32'hbfd949e2, 32'hc09d6b12} /* (29, 16, 17) {real, imag} */,
  {32'h3f9445f9, 32'hc0cdf196} /* (29, 16, 16) {real, imag} */,
  {32'hbf3a1ce7, 32'hc0d7c7d4} /* (29, 16, 15) {real, imag} */,
  {32'hbf1bc8ed, 32'hc0971f26} /* (29, 16, 14) {real, imag} */,
  {32'h3eafc692, 32'hc0867266} /* (29, 16, 13) {real, imag} */,
  {32'h3f1fb225, 32'hc07466fc} /* (29, 16, 12) {real, imag} */,
  {32'hc010419e, 32'hc023c8fe} /* (29, 16, 11) {real, imag} */,
  {32'hc0851f68, 32'h3fe31309} /* (29, 16, 10) {real, imag} */,
  {32'h3f310be0, 32'h407ad4d4} /* (29, 16, 9) {real, imag} */,
  {32'h3efd83c0, 32'h408d90f8} /* (29, 16, 8) {real, imag} */,
  {32'h3fa0dcd4, 32'h40b1420c} /* (29, 16, 7) {real, imag} */,
  {32'h40283e8a, 32'h40fad32e} /* (29, 16, 6) {real, imag} */,
  {32'h40310a9e, 32'h40a9f578} /* (29, 16, 5) {real, imag} */,
  {32'h3fe3ec54, 32'h40c672f0} /* (29, 16, 4) {real, imag} */,
  {32'hbe65b428, 32'h40f6739c} /* (29, 16, 3) {real, imag} */,
  {32'h3fc85017, 32'h410c1f8e} /* (29, 16, 2) {real, imag} */,
  {32'h4054b614, 32'h40f1116c} /* (29, 16, 1) {real, imag} */,
  {32'h3f0da093, 32'h4091a7f6} /* (29, 16, 0) {real, imag} */,
  {32'h3ffd5b98, 32'h40512254} /* (29, 15, 31) {real, imag} */,
  {32'h4053879f, 32'h40d9da49} /* (29, 15, 30) {real, imag} */,
  {32'h403429b9, 32'h409a8462} /* (29, 15, 29) {real, imag} */,
  {32'h3f89f639, 32'h4087800c} /* (29, 15, 28) {real, imag} */,
  {32'h3fe34a12, 32'h4046ae4e} /* (29, 15, 27) {real, imag} */,
  {32'h40782f17, 32'h3fbc108f} /* (29, 15, 26) {real, imag} */,
  {32'h40d85be7, 32'h405e2ae5} /* (29, 15, 25) {real, imag} */,
  {32'h3fe49ae6, 32'h40831c69} /* (29, 15, 24) {real, imag} */,
  {32'h3f01eb9c, 32'h405b6949} /* (29, 15, 23) {real, imag} */,
  {32'h40682d4d, 32'h402d6a8c} /* (29, 15, 22) {real, imag} */,
  {32'h3f903327, 32'hbfc05654} /* (29, 15, 21) {real, imag} */,
  {32'hc07b5097, 32'hc0c6ea7a} /* (29, 15, 20) {real, imag} */,
  {32'hc04ad2e3, 32'hc03569af} /* (29, 15, 19) {real, imag} */,
  {32'hbf1ec740, 32'hc0285b5a} /* (29, 15, 18) {real, imag} */,
  {32'hbd6c36c8, 32'hc07f7248} /* (29, 15, 17) {real, imag} */,
  {32'hc01b681c, 32'hc0be5368} /* (29, 15, 16) {real, imag} */,
  {32'hbf58e613, 32'hc09eb10e} /* (29, 15, 15) {real, imag} */,
  {32'h3e1409bd, 32'hc08ca6c8} /* (29, 15, 14) {real, imag} */,
  {32'hbf972830, 32'hc0c6f1f6} /* (29, 15, 13) {real, imag} */,
  {32'hc031d010, 32'hc0ae6c77} /* (29, 15, 12) {real, imag} */,
  {32'hc0a0834c, 32'hbe96af30} /* (29, 15, 11) {real, imag} */,
  {32'hc07b16ec, 32'h4045a54f} /* (29, 15, 10) {real, imag} */,
  {32'hbfb063fc, 32'h4088f22e} /* (29, 15, 9) {real, imag} */,
  {32'h3ed26e10, 32'h40a3acb9} /* (29, 15, 8) {real, imag} */,
  {32'h40046604, 32'h40b309f0} /* (29, 15, 7) {real, imag} */,
  {32'h402e2f1c, 32'h404ae68d} /* (29, 15, 6) {real, imag} */,
  {32'h4086028c, 32'h407f4f0c} /* (29, 15, 5) {real, imag} */,
  {32'h403d3ff0, 32'h40a4d9c7} /* (29, 15, 4) {real, imag} */,
  {32'h4072c38b, 32'h40ba0a7a} /* (29, 15, 3) {real, imag} */,
  {32'h4095257e, 32'h40cdc506} /* (29, 15, 2) {real, imag} */,
  {32'h40355430, 32'h409fb21c} /* (29, 15, 1) {real, imag} */,
  {32'hbef22ba7, 32'h3fd0d544} /* (29, 15, 0) {real, imag} */,
  {32'h3f9f7290, 32'h4090d176} /* (29, 14, 31) {real, imag} */,
  {32'h405509f2, 32'h40c66895} /* (29, 14, 30) {real, imag} */,
  {32'h407dc35e, 32'h404adb77} /* (29, 14, 29) {real, imag} */,
  {32'h40666b09, 32'h403dd1c0} /* (29, 14, 28) {real, imag} */,
  {32'h400ce2e8, 32'h408d2511} /* (29, 14, 27) {real, imag} */,
  {32'h408352d6, 32'h40954fb2} /* (29, 14, 26) {real, imag} */,
  {32'h40f1dd86, 32'h40a873a0} /* (29, 14, 25) {real, imag} */,
  {32'h40c94e50, 32'h40bb5326} /* (29, 14, 24) {real, imag} */,
  {32'h40a6b5d2, 32'h40d9b15c} /* (29, 14, 23) {real, imag} */,
  {32'h404de288, 32'h40b40ca1} /* (29, 14, 22) {real, imag} */,
  {32'hbf837c8a, 32'h3f2d7c33} /* (29, 14, 21) {real, imag} */,
  {32'hbffd3d83, 32'hc08772d3} /* (29, 14, 20) {real, imag} */,
  {32'hbef01cf8, 32'hc029f946} /* (29, 14, 19) {real, imag} */,
  {32'hbfc81883, 32'hc0545dd8} /* (29, 14, 18) {real, imag} */,
  {32'hc0044bc1, 32'hc0948ca6} /* (29, 14, 17) {real, imag} */,
  {32'hc03aad95, 32'hc0b0ed78} /* (29, 14, 16) {real, imag} */,
  {32'hbff89288, 32'hc03c1138} /* (29, 14, 15) {real, imag} */,
  {32'hbe5114d8, 32'hc0215408} /* (29, 14, 14) {real, imag} */,
  {32'hbff51b5a, 32'hc0c272ac} /* (29, 14, 13) {real, imag} */,
  {32'hc04d93ce, 32'hc09e2144} /* (29, 14, 12) {real, imag} */,
  {32'hc03da8fc, 32'hc036ea74} /* (29, 14, 11) {real, imag} */,
  {32'h3f228186, 32'h40448403} /* (29, 14, 10) {real, imag} */,
  {32'h3fbafa33, 32'h41077e24} /* (29, 14, 9) {real, imag} */,
  {32'h3ff979b3, 32'h4115c190} /* (29, 14, 8) {real, imag} */,
  {32'h4045b407, 32'h40c0f325} /* (29, 14, 7) {real, imag} */,
  {32'h3fe75410, 32'h400b64b0} /* (29, 14, 6) {real, imag} */,
  {32'h40579a54, 32'h40d08ba2} /* (29, 14, 5) {real, imag} */,
  {32'h402adbeb, 32'h40a3cefa} /* (29, 14, 4) {real, imag} */,
  {32'h404834b8, 32'h40bbbc88} /* (29, 14, 3) {real, imag} */,
  {32'h40a160dc, 32'h40476944} /* (29, 14, 2) {real, imag} */,
  {32'h401ebbd1, 32'h40037266} /* (29, 14, 1) {real, imag} */,
  {32'hbfa57640, 32'h3fe3618e} /* (29, 14, 0) {real, imag} */,
  {32'h3edbefe3, 32'h40876fb1} /* (29, 13, 31) {real, imag} */,
  {32'h400420c8, 32'h409099a0} /* (29, 13, 30) {real, imag} */,
  {32'h405acdb6, 32'h40c1ac32} /* (29, 13, 29) {real, imag} */,
  {32'h3fc2a08e, 32'h40dbb699} /* (29, 13, 28) {real, imag} */,
  {32'h40080788, 32'h40be333f} /* (29, 13, 27) {real, imag} */,
  {32'h401cacaa, 32'h40d83d82} /* (29, 13, 26) {real, imag} */,
  {32'h40287188, 32'h40d7d249} /* (29, 13, 25) {real, imag} */,
  {32'h406bea3c, 32'h41015b30} /* (29, 13, 24) {real, imag} */,
  {32'h40466922, 32'h410dd926} /* (29, 13, 23) {real, imag} */,
  {32'h402c9498, 32'h40fbd961} /* (29, 13, 22) {real, imag} */,
  {32'hbc2dc600, 32'h3fd4f1d0} /* (29, 13, 21) {real, imag} */,
  {32'hbf29f668, 32'hc0af83a0} /* (29, 13, 20) {real, imag} */,
  {32'hbf922a1a, 32'hc0c585f0} /* (29, 13, 19) {real, imag} */,
  {32'hc0157600, 32'hc0b45812} /* (29, 13, 18) {real, imag} */,
  {32'hbfd7c7bf, 32'hc0c697bd} /* (29, 13, 17) {real, imag} */,
  {32'hbfbe94be, 32'hc0de6bec} /* (29, 13, 16) {real, imag} */,
  {32'h3f240703, 32'hc058f851} /* (29, 13, 15) {real, imag} */,
  {32'h3f11ba20, 32'hbf137f9d} /* (29, 13, 14) {real, imag} */,
  {32'hc01a585d, 32'hc0683492} /* (29, 13, 13) {real, imag} */,
  {32'hc068471e, 32'hc0bee69a} /* (29, 13, 12) {real, imag} */,
  {32'hc066d065, 32'hc0af6c56} /* (29, 13, 11) {real, imag} */,
  {32'h3f45b14a, 32'h4082dc9e} /* (29, 13, 10) {real, imag} */,
  {32'h408c1990, 32'h4117753c} /* (29, 13, 9) {real, imag} */,
  {32'h403be916, 32'h40edbbef} /* (29, 13, 8) {real, imag} */,
  {32'h4077300d, 32'h40882d2a} /* (29, 13, 7) {real, imag} */,
  {32'h3fb579c3, 32'h409dfbeb} /* (29, 13, 6) {real, imag} */,
  {32'h3fc5d83c, 32'h41113100} /* (29, 13, 5) {real, imag} */,
  {32'h3f9b1a28, 32'h40cf0daa} /* (29, 13, 4) {real, imag} */,
  {32'h3f8822e8, 32'h40be0823} /* (29, 13, 3) {real, imag} */,
  {32'h3fdac35f, 32'h4067182c} /* (29, 13, 2) {real, imag} */,
  {32'h3fa6fc35, 32'h409d2ca0} /* (29, 13, 1) {real, imag} */,
  {32'hbe8b88a5, 32'h407c1950} /* (29, 13, 0) {real, imag} */,
  {32'hbf32d99e, 32'h3fe255f2} /* (29, 12, 31) {real, imag} */,
  {32'hbee9fcc4, 32'h405ab1ec} /* (29, 12, 30) {real, imag} */,
  {32'hbf0c2ace, 32'h4092950a} /* (29, 12, 29) {real, imag} */,
  {32'h3fb1c7b8, 32'h411152c4} /* (29, 12, 28) {real, imag} */,
  {32'h4023d1b8, 32'h411df772} /* (29, 12, 27) {real, imag} */,
  {32'h40209c82, 32'h40f2567e} /* (29, 12, 26) {real, imag} */,
  {32'h3fe97ef0, 32'h4104d0b4} /* (29, 12, 25) {real, imag} */,
  {32'h3fb27715, 32'h411d57c4} /* (29, 12, 24) {real, imag} */,
  {32'h402310bf, 32'h40d53659} /* (29, 12, 23) {real, imag} */,
  {32'h402978c8, 32'h408e8612} /* (29, 12, 22) {real, imag} */,
  {32'hbf9b3170, 32'h3ec10af2} /* (29, 12, 21) {real, imag} */,
  {32'hbfb8051a, 32'hc0b65841} /* (29, 12, 20) {real, imag} */,
  {32'h3f58ec9d, 32'hc0d3eba4} /* (29, 12, 19) {real, imag} */,
  {32'hc004d0b0, 32'hc0cb7691} /* (29, 12, 18) {real, imag} */,
  {32'hc059442a, 32'hc0b8fb3a} /* (29, 12, 17) {real, imag} */,
  {32'h3f9113ad, 32'hc0bc1d0a} /* (29, 12, 16) {real, imag} */,
  {32'h404174d0, 32'hc087defc} /* (29, 12, 15) {real, imag} */,
  {32'hbc4aa870, 32'hc005bb47} /* (29, 12, 14) {real, imag} */,
  {32'hc089a2c7, 32'hbfe0bfd4} /* (29, 12, 13) {real, imag} */,
  {32'hc08b59fb, 32'hc08b6f4d} /* (29, 12, 12) {real, imag} */,
  {32'hc0991358, 32'hc08e0b2d} /* (29, 12, 11) {real, imag} */,
  {32'hbfd67e20, 32'h40657e66} /* (29, 12, 10) {real, imag} */,
  {32'h3f81e89e, 32'h40d4d477} /* (29, 12, 9) {real, imag} */,
  {32'h4034f774, 32'h40a783b8} /* (29, 12, 8) {real, imag} */,
  {32'h40000254, 32'h40923f3e} /* (29, 12, 7) {real, imag} */,
  {32'h3e99dbd6, 32'h40f68f40} /* (29, 12, 6) {real, imag} */,
  {32'h3fa212c5, 32'h40ecbb74} /* (29, 12, 5) {real, imag} */,
  {32'h3eea2ed6, 32'h40b33296} /* (29, 12, 4) {real, imag} */,
  {32'h3ed54984, 32'h409f2878} /* (29, 12, 3) {real, imag} */,
  {32'h3ee0f9ce, 32'h40d61b4e} /* (29, 12, 2) {real, imag} */,
  {32'h3f644a5a, 32'h41185e24} /* (29, 12, 1) {real, imag} */,
  {32'hbf73334f, 32'h40bd00b7} /* (29, 12, 0) {real, imag} */,
  {32'hbf6a6f29, 32'h40108b0c} /* (29, 11, 31) {real, imag} */,
  {32'hbfe96428, 32'h4068be15} /* (29, 11, 30) {real, imag} */,
  {32'h3febc604, 32'h404435de} /* (29, 11, 29) {real, imag} */,
  {32'h400fe54e, 32'h40b4d082} /* (29, 11, 28) {real, imag} */,
  {32'h40027764, 32'h410884a3} /* (29, 11, 27) {real, imag} */,
  {32'h40673494, 32'h40a9eae0} /* (29, 11, 26) {real, imag} */,
  {32'h401341cc, 32'h40cb0d6e} /* (29, 11, 25) {real, imag} */,
  {32'h3f647fba, 32'h40e21f3e} /* (29, 11, 24) {real, imag} */,
  {32'h3f9656d0, 32'h4028dc46} /* (29, 11, 23) {real, imag} */,
  {32'hbe167e58, 32'h408bda4e} /* (29, 11, 22) {real, imag} */,
  {32'hc075dbbc, 32'h3fcf5fae} /* (29, 11, 21) {real, imag} */,
  {32'hc03a36e6, 32'hc01add60} /* (29, 11, 20) {real, imag} */,
  {32'h4015a686, 32'hc09e6aaa} /* (29, 11, 19) {real, imag} */,
  {32'h3d8e005c, 32'hc09ff11f} /* (29, 11, 18) {real, imag} */,
  {32'hc024f3f2, 32'hc03b8694} /* (29, 11, 17) {real, imag} */,
  {32'h3fcfe389, 32'hc070609c} /* (29, 11, 16) {real, imag} */,
  {32'h3f17e0c0, 32'hc0a99bb1} /* (29, 11, 15) {real, imag} */,
  {32'hbf7b1dca, 32'hc0834a47} /* (29, 11, 14) {real, imag} */,
  {32'hbf960516, 32'hc08ad824} /* (29, 11, 13) {real, imag} */,
  {32'hbfe36012, 32'hc08d834c} /* (29, 11, 12) {real, imag} */,
  {32'hbfe11412, 32'hc084e4fb} /* (29, 11, 11) {real, imag} */,
  {32'h3f302583, 32'h3f849ffe} /* (29, 11, 10) {real, imag} */,
  {32'h3eb94eaa, 32'h40a1d45c} /* (29, 11, 9) {real, imag} */,
  {32'h3fa1c922, 32'h40b0ad3c} /* (29, 11, 8) {real, imag} */,
  {32'h3fec4ec9, 32'h40ce01c0} /* (29, 11, 7) {real, imag} */,
  {32'h3fee3e2e, 32'h40b24c0e} /* (29, 11, 6) {real, imag} */,
  {32'h3f844d8c, 32'h408c349f} /* (29, 11, 5) {real, imag} */,
  {32'hbb88c780, 32'h402e830c} /* (29, 11, 4) {real, imag} */,
  {32'hbe21961a, 32'h4076c964} /* (29, 11, 3) {real, imag} */,
  {32'h3f24382e, 32'h40b254fa} /* (29, 11, 2) {real, imag} */,
  {32'hbf5a3840, 32'h40c288c8} /* (29, 11, 1) {real, imag} */,
  {32'hbf9e2e9a, 32'h407169c9} /* (29, 11, 0) {real, imag} */,
  {32'hbc2bdfa0, 32'hbf3b55de} /* (29, 10, 31) {real, imag} */,
  {32'hbf99d21c, 32'hbf1f6742} /* (29, 10, 30) {real, imag} */,
  {32'h3f659762, 32'h3ecdc93a} /* (29, 10, 29) {real, imag} */,
  {32'h3d9f3718, 32'h3d790510} /* (29, 10, 28) {real, imag} */,
  {32'hbfa3401a, 32'hbfa1f6b8} /* (29, 10, 27) {real, imag} */,
  {32'h3ea206a0, 32'hbf9f3838} /* (29, 10, 26) {real, imag} */,
  {32'h3fd91645, 32'hbff8286a} /* (29, 10, 25) {real, imag} */,
  {32'h3d98a490, 32'hbf422630} /* (29, 10, 24) {real, imag} */,
  {32'hbfb7cd60, 32'hc09da647} /* (29, 10, 23) {real, imag} */,
  {32'hc04c8029, 32'hc031bc1c} /* (29, 10, 22) {real, imag} */,
  {32'hbf34a51c, 32'hc0493dc7} /* (29, 10, 21) {real, imag} */,
  {32'h3feb2830, 32'h3f665a07} /* (29, 10, 20) {real, imag} */,
  {32'h3ff4f516, 32'h402ba6a8} /* (29, 10, 19) {real, imag} */,
  {32'h3f6b7a73, 32'h3fe84883} /* (29, 10, 18) {real, imag} */,
  {32'h40249b7e, 32'h40b567d8} /* (29, 10, 17) {real, imag} */,
  {32'h3f6dbafe, 32'h407e26ee} /* (29, 10, 16) {real, imag} */,
  {32'hc0332004, 32'h3f6fd99e} /* (29, 10, 15) {real, imag} */,
  {32'hbf17b9fe, 32'h3f8fc9f6} /* (29, 10, 14) {real, imag} */,
  {32'hbd47c7ba, 32'h3ed1f63a} /* (29, 10, 13) {real, imag} */,
  {32'h3f281464, 32'h400cf29c} /* (29, 10, 12) {real, imag} */,
  {32'h3faa88af, 32'h3fdb9ae4} /* (29, 10, 11) {real, imag} */,
  {32'h3f985f19, 32'hbecb7a4a} /* (29, 10, 10) {real, imag} */,
  {32'hbefd1332, 32'h3a4f3a00} /* (29, 10, 9) {real, imag} */,
  {32'hbe9487d7, 32'hbfaf55b8} /* (29, 10, 8) {real, imag} */,
  {32'h3f8f5f50, 32'hbfce7413} /* (29, 10, 7) {real, imag} */,
  {32'h3f4fd752, 32'hc016b3d7} /* (29, 10, 6) {real, imag} */,
  {32'h3e77de34, 32'hbf3a61df} /* (29, 10, 5) {real, imag} */,
  {32'h3f0889c4, 32'hc0728d2b} /* (29, 10, 4) {real, imag} */,
  {32'hc000fbe4, 32'hc08a31dd} /* (29, 10, 3) {real, imag} */,
  {32'hc000e00a, 32'hbf68e017} /* (29, 10, 2) {real, imag} */,
  {32'hbfffa6d4, 32'hbfadb452} /* (29, 10, 1) {real, imag} */,
  {32'hbf89ed43, 32'hbffde762} /* (29, 10, 0) {real, imag} */,
  {32'hbff440fc, 32'hc0c3e124} /* (29, 9, 31) {real, imag} */,
  {32'hc02c520c, 32'hc0fa84b4} /* (29, 9, 30) {real, imag} */,
  {32'hbff92a26, 32'hc0d72a14} /* (29, 9, 29) {real, imag} */,
  {32'hbe9ee5bb, 32'hc062f9fc} /* (29, 9, 28) {real, imag} */,
  {32'hbdb78ff0, 32'hc0948044} /* (29, 9, 27) {real, imag} */,
  {32'hbfcbc558, 32'hc06c311e} /* (29, 9, 26) {real, imag} */,
  {32'hbf9fbe38, 32'hc0a70491} /* (29, 9, 25) {real, imag} */,
  {32'hbfd97819, 32'hc09a169e} /* (29, 9, 24) {real, imag} */,
  {32'hc052be3c, 32'hc0e9939a} /* (29, 9, 23) {real, imag} */,
  {32'hc0982956, 32'hc0e4591c} /* (29, 9, 22) {real, imag} */,
  {32'hc054bf7a, 32'hc073b006} /* (29, 9, 21) {real, imag} */,
  {32'h40263b42, 32'h3fb10eee} /* (29, 9, 20) {real, imag} */,
  {32'h4020c176, 32'h40acbec9} /* (29, 9, 19) {real, imag} */,
  {32'h3f2bf702, 32'h406eee5c} /* (29, 9, 18) {real, imag} */,
  {32'h3fb3d29b, 32'h40ac6642} /* (29, 9, 17) {real, imag} */,
  {32'hbfdc5136, 32'h40baeff1} /* (29, 9, 16) {real, imag} */,
  {32'hbf6916b7, 32'h405c072c} /* (29, 9, 15) {real, imag} */,
  {32'h3dde2a98, 32'h4019cb29} /* (29, 9, 14) {real, imag} */,
  {32'h3fa968eb, 32'h40b20b45} /* (29, 9, 13) {real, imag} */,
  {32'h3f8b22d8, 32'h4111f0a3} /* (29, 9, 12) {real, imag} */,
  {32'h3fca34d3, 32'h40c1be30} /* (29, 9, 11) {real, imag} */,
  {32'hbc7d7120, 32'h3f3e4c40} /* (29, 9, 10) {real, imag} */,
  {32'hbf88d5cd, 32'hbfcf2878} /* (29, 9, 9) {real, imag} */,
  {32'hbed039b2, 32'hc098be91} /* (29, 9, 8) {real, imag} */,
  {32'hbfffab2e, 32'hc0b014b3} /* (29, 9, 7) {real, imag} */,
  {32'hc045ba3e, 32'hc05ee25b} /* (29, 9, 6) {real, imag} */,
  {32'h3d5379b0, 32'hc03a723e} /* (29, 9, 5) {real, imag} */,
  {32'hc000ab3a, 32'hc0982774} /* (29, 9, 4) {real, imag} */,
  {32'hc074b346, 32'hc1140d3c} /* (29, 9, 3) {real, imag} */,
  {32'hc07476fc, 32'hc0e1d47a} /* (29, 9, 2) {real, imag} */,
  {32'hc03d1121, 32'hc08ad423} /* (29, 9, 1) {real, imag} */,
  {32'hbfc6a05a, 32'hc039aa2e} /* (29, 9, 0) {real, imag} */,
  {32'hc00cfa62, 32'hc070dd73} /* (29, 8, 31) {real, imag} */,
  {32'hc07d1817, 32'hc0ae174c} /* (29, 8, 30) {real, imag} */,
  {32'hc013257e, 32'hc0f660cd} /* (29, 8, 29) {real, imag} */,
  {32'h3fb26afc, 32'hc063ae25} /* (29, 8, 28) {real, imag} */,
  {32'h402d0d2f, 32'hc08bf33d} /* (29, 8, 27) {real, imag} */,
  {32'h3f6bba6c, 32'hc0b8fca5} /* (29, 8, 26) {real, imag} */,
  {32'h3edb7348, 32'hc0aa2508} /* (29, 8, 25) {real, imag} */,
  {32'hbff4da6e, 32'hc0ab0901} /* (29, 8, 24) {real, imag} */,
  {32'hc05f3722, 32'hc0da8135} /* (29, 8, 23) {real, imag} */,
  {32'hc0d29a70, 32'hc0d7c1f0} /* (29, 8, 22) {real, imag} */,
  {32'hc08f07f1, 32'hbf4bf242} /* (29, 8, 21) {real, imag} */,
  {32'h3f8796d0, 32'h4060a864} /* (29, 8, 20) {real, imag} */,
  {32'h401818dc, 32'h40a73a4d} /* (29, 8, 19) {real, imag} */,
  {32'h3fc1f52f, 32'h40d14b4a} /* (29, 8, 18) {real, imag} */,
  {32'h3f1d9ad5, 32'h40dd9599} /* (29, 8, 17) {real, imag} */,
  {32'hbf5a2850, 32'h40a3907f} /* (29, 8, 16) {real, imag} */,
  {32'h3fd2bfea, 32'h405b163a} /* (29, 8, 15) {real, imag} */,
  {32'h40673d3c, 32'h4091902e} /* (29, 8, 14) {real, imag} */,
  {32'h406b34ea, 32'h40ced7f1} /* (29, 8, 13) {real, imag} */,
  {32'h3f54558e, 32'h41136d05} /* (29, 8, 12) {real, imag} */,
  {32'h400c33f2, 32'h40a53e11} /* (29, 8, 11) {real, imag} */,
  {32'h3f5c07df, 32'hbf4e6fd5} /* (29, 8, 10) {real, imag} */,
  {32'hbee8655a, 32'hc0695e66} /* (29, 8, 9) {real, imag} */,
  {32'hbf7a45da, 32'hc0d68e46} /* (29, 8, 8) {real, imag} */,
  {32'hbfffd0b7, 32'hc0cfddfb} /* (29, 8, 7) {real, imag} */,
  {32'hc0075820, 32'hc0868211} /* (29, 8, 6) {real, imag} */,
  {32'h3f908306, 32'hc0421943} /* (29, 8, 5) {real, imag} */,
  {32'hbf16025d, 32'hc0bf037e} /* (29, 8, 4) {real, imag} */,
  {32'hc0631b0a, 32'hc0eb0f26} /* (29, 8, 3) {real, imag} */,
  {32'hc073c2ac, 32'hc0c3a29c} /* (29, 8, 2) {real, imag} */,
  {32'hbf8cc938, 32'hc0b15390} /* (29, 8, 1) {real, imag} */,
  {32'h3fe1591e, 32'hc01d5970} /* (29, 8, 0) {real, imag} */,
  {32'hbfaba2e2, 32'hbf69882e} /* (29, 7, 31) {real, imag} */,
  {32'hc04d5930, 32'hc0542640} /* (29, 7, 30) {real, imag} */,
  {32'hbd5a4c30, 32'hc0e37dee} /* (29, 7, 29) {real, imag} */,
  {32'h3fc1f19e, 32'hc0edf586} /* (29, 7, 28) {real, imag} */,
  {32'h3f88de0a, 32'hc0c5563a} /* (29, 7, 27) {real, imag} */,
  {32'hbfab0d0d, 32'hc0baa85e} /* (29, 7, 26) {real, imag} */,
  {32'hbff2fc19, 32'hc0a77a79} /* (29, 7, 25) {real, imag} */,
  {32'hc0202a42, 32'hc0d3a3b4} /* (29, 7, 24) {real, imag} */,
  {32'hc06105cf, 32'hc0c4c2d3} /* (29, 7, 23) {real, imag} */,
  {32'hc082652c, 32'hc05dabe0} /* (29, 7, 22) {real, imag} */,
  {32'hbf835650, 32'h40033ec8} /* (29, 7, 21) {real, imag} */,
  {32'h40133d5e, 32'h40c6712a} /* (29, 7, 20) {real, imag} */,
  {32'h40569c8b, 32'h4085c39d} /* (29, 7, 19) {real, imag} */,
  {32'h3e3b9408, 32'h406831b7} /* (29, 7, 18) {real, imag} */,
  {32'h3f8e0a0c, 32'h40e3dacf} /* (29, 7, 17) {real, imag} */,
  {32'h4007f3c7, 32'h40d002a6} /* (29, 7, 16) {real, imag} */,
  {32'h4073cc74, 32'h409964ca} /* (29, 7, 15) {real, imag} */,
  {32'h40941af9, 32'h40c38676} /* (29, 7, 14) {real, imag} */,
  {32'h40778623, 32'h40b76cf3} /* (29, 7, 13) {real, imag} */,
  {32'hbf8466d0, 32'h4089e83e} /* (29, 7, 12) {real, imag} */,
  {32'hc06bec38, 32'h4023e113} /* (29, 7, 11) {real, imag} */,
  {32'hbea46b22, 32'hc0187458} /* (29, 7, 10) {real, imag} */,
  {32'h3dfcb200, 32'hc0c6ebc5} /* (29, 7, 9) {real, imag} */,
  {32'hbf882ca8, 32'hc0d3f2bc} /* (29, 7, 8) {real, imag} */,
  {32'h3f94fad5, 32'hc057a684} /* (29, 7, 7) {real, imag} */,
  {32'h3f2a977a, 32'hc050ea5c} /* (29, 7, 6) {real, imag} */,
  {32'hc01f2868, 32'hc0b8b79b} /* (29, 7, 5) {real, imag} */,
  {32'hbe46bb9c, 32'hc0db7c7c} /* (29, 7, 4) {real, imag} */,
  {32'hbfca062b, 32'hc1017026} /* (29, 7, 3) {real, imag} */,
  {32'hc0a02c1c, 32'hc0ed7df0} /* (29, 7, 2) {real, imag} */,
  {32'hc002561e, 32'hc0c000c6} /* (29, 7, 1) {real, imag} */,
  {32'hbd0e6618, 32'hc012529f} /* (29, 7, 0) {real, imag} */,
  {32'hbef0f380, 32'hc00f07b8} /* (29, 6, 31) {real, imag} */,
  {32'hbf9b25d2, 32'hc0774eed} /* (29, 6, 30) {real, imag} */,
  {32'h3fc5750e, 32'hc0ea971d} /* (29, 6, 29) {real, imag} */,
  {32'h3eb3c5be, 32'hc0fb6f46} /* (29, 6, 28) {real, imag} */,
  {32'hc07f6577, 32'hc0bace02} /* (29, 6, 27) {real, imag} */,
  {32'hc08df2e4, 32'hc0b4c673} /* (29, 6, 26) {real, imag} */,
  {32'hc04cefbe, 32'hc08fc8b8} /* (29, 6, 25) {real, imag} */,
  {32'hbf557ffc, 32'hc0c36dce} /* (29, 6, 24) {real, imag} */,
  {32'hbfd74202, 32'hc0b2bf3e} /* (29, 6, 23) {real, imag} */,
  {32'hc08f804c, 32'hc056d0ac} /* (29, 6, 22) {real, imag} */,
  {32'hbf866d14, 32'hbf147aa4} /* (29, 6, 21) {real, imag} */,
  {32'h40869b38, 32'h405cce8a} /* (29, 6, 20) {real, imag} */,
  {32'h4059c510, 32'h400baec0} /* (29, 6, 19) {real, imag} */,
  {32'h3d82735c, 32'h400255b0} /* (29, 6, 18) {real, imag} */,
  {32'hbe4cfbca, 32'h4090f409} /* (29, 6, 17) {real, imag} */,
  {32'h3e3440cc, 32'h40baa8c4} /* (29, 6, 16) {real, imag} */,
  {32'h405aef0d, 32'h40c06559} /* (29, 6, 15) {real, imag} */,
  {32'h3ff8891c, 32'h40c83b19} /* (29, 6, 14) {real, imag} */,
  {32'h4032b8b0, 32'h40c17014} /* (29, 6, 13) {real, imag} */,
  {32'h3fb5728b, 32'h40c10400} /* (29, 6, 12) {real, imag} */,
  {32'hbfec3f0a, 32'h40b479fd} /* (29, 6, 11) {real, imag} */,
  {32'hc05f5166, 32'hc00b3b53} /* (29, 6, 10) {real, imag} */,
  {32'hc0906dd6, 32'hc0980e14} /* (29, 6, 9) {real, imag} */,
  {32'hc06319a8, 32'hc047457e} /* (29, 6, 8) {real, imag} */,
  {32'h3fbdae13, 32'hc0876fde} /* (29, 6, 7) {real, imag} */,
  {32'hbde35a54, 32'hc0bc6bbe} /* (29, 6, 6) {real, imag} */,
  {32'hc08d0c1a, 32'hc0f2c7eb} /* (29, 6, 5) {real, imag} */,
  {32'hc0156b48, 32'hc089875f} /* (29, 6, 4) {real, imag} */,
  {32'h3ed983fa, 32'hc075f7c9} /* (29, 6, 3) {real, imag} */,
  {32'h3c72d580, 32'hc0b81c46} /* (29, 6, 2) {real, imag} */,
  {32'h3f74b34c, 32'hc0b88e2e} /* (29, 6, 1) {real, imag} */,
  {32'hbe84322a, 32'hc05abd48} /* (29, 6, 0) {real, imag} */,
  {32'hc0409ec8, 32'hc088cc55} /* (29, 5, 31) {real, imag} */,
  {32'hc05025d5, 32'hc06b08ca} /* (29, 5, 30) {real, imag} */,
  {32'hbe390230, 32'hc0a100d2} /* (29, 5, 29) {real, imag} */,
  {32'hbfa04f53, 32'hc0f0e0fc} /* (29, 5, 28) {real, imag} */,
  {32'hc05492cc, 32'hc0cc4bfe} /* (29, 5, 27) {real, imag} */,
  {32'hc00a4f3e, 32'hc10c1f89} /* (29, 5, 26) {real, imag} */,
  {32'hbfb6a9d3, 32'hc10a4273} /* (29, 5, 25) {real, imag} */,
  {32'hc044435a, 32'hc0d44398} /* (29, 5, 24) {real, imag} */,
  {32'hbfa5e8eb, 32'hc0c81f12} /* (29, 5, 23) {real, imag} */,
  {32'hc0248e56, 32'hc0c9ab02} /* (29, 5, 22) {real, imag} */,
  {32'hbf9c1336, 32'hc0bbf53a} /* (29, 5, 21) {real, imag} */,
  {32'h3fdb65bd, 32'hc0a20cad} /* (29, 5, 20) {real, imag} */,
  {32'h4023c2e7, 32'hc05953ba} /* (29, 5, 19) {real, imag} */,
  {32'h40104467, 32'hbfc2dfb0} /* (29, 5, 18) {real, imag} */,
  {32'h3f166a8a, 32'hc0286461} /* (29, 5, 17) {real, imag} */,
  {32'hbfa8fc38, 32'hbfcacd0a} /* (29, 5, 16) {real, imag} */,
  {32'h3faa3188, 32'h409180df} /* (29, 5, 15) {real, imag} */,
  {32'h401708c4, 32'h4091b1f6} /* (29, 5, 14) {real, imag} */,
  {32'h40474bba, 32'h40c792f1} /* (29, 5, 13) {real, imag} */,
  {32'h3fa862fc, 32'h40ff8a1e} /* (29, 5, 12) {real, imag} */,
  {32'h40387b80, 32'h40e10c44} /* (29, 5, 11) {real, imag} */,
  {32'h3fd751f8, 32'h3fdd477a} /* (29, 5, 10) {real, imag} */,
  {32'hbf766ec2, 32'h3ea5bbe8} /* (29, 5, 9) {real, imag} */,
  {32'h3fa36036, 32'h3f1c378e} /* (29, 5, 8) {real, imag} */,
  {32'h3ff4ef0d, 32'hbf8aa11a} /* (29, 5, 7) {real, imag} */,
  {32'h3f1d2e04, 32'hbf93f626} /* (29, 5, 6) {real, imag} */,
  {32'hc0169a8e, 32'hc09a39f4} /* (29, 5, 5) {real, imag} */,
  {32'hc0423246, 32'hc0881f33} /* (29, 5, 4) {real, imag} */,
  {32'hbf9fc77d, 32'hc03e2292} /* (29, 5, 3) {real, imag} */,
  {32'h3fa826c7, 32'hc0873b66} /* (29, 5, 2) {real, imag} */,
  {32'h3f82cf17, 32'hc0e4408f} /* (29, 5, 1) {real, imag} */,
  {32'hbf7ba3b4, 32'hc0b1b16f} /* (29, 5, 0) {real, imag} */,
  {32'hc020a680, 32'hc060e288} /* (29, 4, 31) {real, imag} */,
  {32'hc005d34a, 32'hc095073c} /* (29, 4, 30) {real, imag} */,
  {32'h3f51a2bc, 32'hc0825e46} /* (29, 4, 29) {real, imag} */,
  {32'hbf94c211, 32'hc0fc21db} /* (29, 4, 28) {real, imag} */,
  {32'hc01e2685, 32'hc113d960} /* (29, 4, 27) {real, imag} */,
  {32'hc0207459, 32'hc0fe1e6e} /* (29, 4, 26) {real, imag} */,
  {32'hbf9f894d, 32'hc0d16aa4} /* (29, 4, 25) {real, imag} */,
  {32'hc091ce93, 32'hc0bb837c} /* (29, 4, 24) {real, imag} */,
  {32'hc001b111, 32'hc087a940} /* (29, 4, 23) {real, imag} */,
  {32'hbf264955, 32'hc0129e66} /* (29, 4, 22) {real, imag} */,
  {32'h3eb4b4d2, 32'hbfe723b9} /* (29, 4, 21) {real, imag} */,
  {32'hbf676bdb, 32'hc0c63d8c} /* (29, 4, 20) {real, imag} */,
  {32'hbe45bbfe, 32'hc0bfd534} /* (29, 4, 19) {real, imag} */,
  {32'hba8e4100, 32'hc092e091} /* (29, 4, 18) {real, imag} */,
  {32'h3f4e0678, 32'hc0acdccb} /* (29, 4, 17) {real, imag} */,
  {32'hbf5c34f9, 32'hc04dff78} /* (29, 4, 16) {real, imag} */,
  {32'h3fcc3c1e, 32'h40cae614} /* (29, 4, 15) {real, imag} */,
  {32'h4076be20, 32'h404939f4} /* (29, 4, 14) {real, imag} */,
  {32'h4015fb5c, 32'h408b02c0} /* (29, 4, 13) {real, imag} */,
  {32'hbe0ffdd8, 32'h40dd6402} /* (29, 4, 12) {real, imag} */,
  {32'h3e77d3a0, 32'h40cad47b} /* (29, 4, 11) {real, imag} */,
  {32'h4032df9c, 32'h40a1968e} /* (29, 4, 10) {real, imag} */,
  {32'h403b5299, 32'h3f9acb90} /* (29, 4, 9) {real, imag} */,
  {32'h4003a506, 32'h40095675} /* (29, 4, 8) {real, imag} */,
  {32'h404892da, 32'h403750b1} /* (29, 4, 7) {real, imag} */,
  {32'h3fe7c51f, 32'h409d037a} /* (29, 4, 6) {real, imag} */,
  {32'hc031df10, 32'h3ee7f9c9} /* (29, 4, 5) {real, imag} */,
  {32'hbfa1f2e4, 32'hc02db69e} /* (29, 4, 4) {real, imag} */,
  {32'hc04f9281, 32'hc095f957} /* (29, 4, 3) {real, imag} */,
  {32'hc029ec14, 32'hc09d413e} /* (29, 4, 2) {real, imag} */,
  {32'hbfe825ee, 32'hc0bb5e0c} /* (29, 4, 1) {real, imag} */,
  {32'hbfb34724, 32'hc086589d} /* (29, 4, 0) {real, imag} */,
  {32'hc0176bd6, 32'hc00db347} /* (29, 3, 31) {real, imag} */,
  {32'hc036a821, 32'hc0ccb838} /* (29, 3, 30) {real, imag} */,
  {32'h3fdef498, 32'hc0f92023} /* (29, 3, 29) {real, imag} */,
  {32'hbfbec5e8, 32'hc1089daa} /* (29, 3, 28) {real, imag} */,
  {32'hc08182a9, 32'hc102f916} /* (29, 3, 27) {real, imag} */,
  {32'hc043fd00, 32'hc0d5fbd3} /* (29, 3, 26) {real, imag} */,
  {32'hc00f8b9b, 32'hc0b8651f} /* (29, 3, 25) {real, imag} */,
  {32'hc004b038, 32'hc0b277c4} /* (29, 3, 24) {real, imag} */,
  {32'hbfceb00c, 32'hc01ac16f} /* (29, 3, 23) {real, imag} */,
  {32'hbfa0302e, 32'hbeaeb4d6} /* (29, 3, 22) {real, imag} */,
  {32'hbf73dc22, 32'hc04a115d} /* (29, 3, 21) {real, imag} */,
  {32'hc011a93f, 32'hc0aa748b} /* (29, 3, 20) {real, imag} */,
  {32'hc0267a0f, 32'hc09a2a5c} /* (29, 3, 19) {real, imag} */,
  {32'hc02dc48d, 32'hc071e2c0} /* (29, 3, 18) {real, imag} */,
  {32'hc00ddcea, 32'hc0aef9cb} /* (29, 3, 17) {real, imag} */,
  {32'hc009ae40, 32'hc09a1f7d} /* (29, 3, 16) {real, imag} */,
  {32'hbf3cc29a, 32'h401b6bea} /* (29, 3, 15) {real, imag} */,
  {32'h3fec06b4, 32'h40963dee} /* (29, 3, 14) {real, imag} */,
  {32'h3ff764e4, 32'h40c87840} /* (29, 3, 13) {real, imag} */,
  {32'h3ed86a66, 32'h40dd206f} /* (29, 3, 12) {real, imag} */,
  {32'hbfe6cf48, 32'h40c2919e} /* (29, 3, 11) {real, imag} */,
  {32'h3e926560, 32'h40ccafd2} /* (29, 3, 10) {real, imag} */,
  {32'h3fb4f755, 32'h3fdf2b2a} /* (29, 3, 9) {real, imag} */,
  {32'hbfc1217a, 32'h402bbf0c} /* (29, 3, 8) {real, imag} */,
  {32'h3f4ce0d2, 32'h40e3d674} /* (29, 3, 7) {real, imag} */,
  {32'h3f7a8397, 32'h4101d836} /* (29, 3, 6) {real, imag} */,
  {32'hc0417429, 32'h404b9a48} /* (29, 3, 5) {real, imag} */,
  {32'hbf939c9b, 32'hbff6ba1c} /* (29, 3, 4) {real, imag} */,
  {32'hc0ab3be8, 32'hc0dcf364} /* (29, 3, 3) {real, imag} */,
  {32'hc091924d, 32'hc0f47d6e} /* (29, 3, 2) {real, imag} */,
  {32'hc0311a24, 32'hc0d0f5ef} /* (29, 3, 1) {real, imag} */,
  {32'hc00c633e, 32'hc072fef0} /* (29, 3, 0) {real, imag} */,
  {32'hc0447305, 32'hc017e3ac} /* (29, 2, 31) {real, imag} */,
  {32'hc0b7f99b, 32'hc09e9d2f} /* (29, 2, 30) {real, imag} */,
  {32'hbff1bd5f, 32'hc0fb14ac} /* (29, 2, 29) {real, imag} */,
  {32'hbf8a097a, 32'hc0fb2db2} /* (29, 2, 28) {real, imag} */,
  {32'hbffb72d4, 32'hc0c835d1} /* (29, 2, 27) {real, imag} */,
  {32'hbf132d95, 32'hc0cd8666} /* (29, 2, 26) {real, imag} */,
  {32'hbfd1f94f, 32'hc0cd054a} /* (29, 2, 25) {real, imag} */,
  {32'hc0356a8b, 32'hc0801a82} /* (29, 2, 24) {real, imag} */,
  {32'hc035e6e6, 32'hbf94e2a2} /* (29, 2, 23) {real, imag} */,
  {32'hc0b5b828, 32'hc0841513} /* (29, 2, 22) {real, imag} */,
  {32'hc08b5da0, 32'hc10b427e} /* (29, 2, 21) {real, imag} */,
  {32'hbfa4f828, 32'hc113543c} /* (29, 2, 20) {real, imag} */,
  {32'hbf327ba6, 32'hc0e1b94a} /* (29, 2, 19) {real, imag} */,
  {32'h3f9b5b16, 32'hc0835031} /* (29, 2, 18) {real, imag} */,
  {32'hc016e6d1, 32'hc0cb0f92} /* (29, 2, 17) {real, imag} */,
  {32'hc0bf7418, 32'hc018a166} /* (29, 2, 16) {real, imag} */,
  {32'hc05e9d17, 32'h4071dff3} /* (29, 2, 15) {real, imag} */,
  {32'h3f33f07a, 32'h409efd54} /* (29, 2, 14) {real, imag} */,
  {32'h3f5fb81d, 32'h40927e8a} /* (29, 2, 13) {real, imag} */,
  {32'hbf957517, 32'h40ca1687} /* (29, 2, 12) {real, imag} */,
  {32'h3ec94c34, 32'h40f50460} /* (29, 2, 11) {real, imag} */,
  {32'h3fa22ed2, 32'h4106fcdc} /* (29, 2, 10) {real, imag} */,
  {32'h3fcc2107, 32'h410e4d94} /* (29, 2, 9) {real, imag} */,
  {32'hbefe1e76, 32'h4098f0cf} /* (29, 2, 8) {real, imag} */,
  {32'hbff2ffea, 32'h40e5c952} /* (29, 2, 7) {real, imag} */,
  {32'h3f85b46a, 32'h41219c84} /* (29, 2, 6) {real, imag} */,
  {32'h3f3524c8, 32'h3f9db1e9} /* (29, 2, 5) {real, imag} */,
  {32'h3db4ddc8, 32'hc08c22c3} /* (29, 2, 4) {real, imag} */,
  {32'hc079fa98, 32'hc0ad9b03} /* (29, 2, 3) {real, imag} */,
  {32'hc09705bc, 32'hc0732f24} /* (29, 2, 2) {real, imag} */,
  {32'hc067d582, 32'hc0a745da} /* (29, 2, 1) {real, imag} */,
  {32'hc017bfce, 32'hc08ced7a} /* (29, 2, 0) {real, imag} */,
  {32'hbf9df608, 32'hbff9d01c} /* (29, 1, 31) {real, imag} */,
  {32'hc015264d, 32'hc048b739} /* (29, 1, 30) {real, imag} */,
  {32'hbfbdb12c, 32'hc076e5df} /* (29, 1, 29) {real, imag} */,
  {32'h3e5bafda, 32'hc092f1ee} /* (29, 1, 28) {real, imag} */,
  {32'hbf5affa0, 32'hc0bb7be4} /* (29, 1, 27) {real, imag} */,
  {32'hbf140ebe, 32'hc0c86882} /* (29, 1, 26) {real, imag} */,
  {32'hbfa2b647, 32'hc0d4a30b} /* (29, 1, 25) {real, imag} */,
  {32'hbfbe9011, 32'hc08fed5e} /* (29, 1, 24) {real, imag} */,
  {32'hc067c494, 32'hc00c36a2} /* (29, 1, 23) {real, imag} */,
  {32'hc06d1cbc, 32'hc083213c} /* (29, 1, 22) {real, imag} */,
  {32'hbf939799, 32'hc0e4bc8e} /* (29, 1, 21) {real, imag} */,
  {32'hbf3f83f2, 32'hc089e6c2} /* (29, 1, 20) {real, imag} */,
  {32'hbe0ec798, 32'hc0a33d8e} /* (29, 1, 19) {real, imag} */,
  {32'h3fadf332, 32'hc0b148bc} /* (29, 1, 18) {real, imag} */,
  {32'hc0143646, 32'hc0bfec40} /* (29, 1, 17) {real, imag} */,
  {32'hc08f6d25, 32'hc06827f2} /* (29, 1, 16) {real, imag} */,
  {32'hbfdbe7e5, 32'h3fdb2fac} /* (29, 1, 15) {real, imag} */,
  {32'hbf0661fb, 32'h4079355b} /* (29, 1, 14) {real, imag} */,
  {32'h3eed5d84, 32'h409bc014} /* (29, 1, 13) {real, imag} */,
  {32'h3febdcc2, 32'h40d112a8} /* (29, 1, 12) {real, imag} */,
  {32'h403b4306, 32'h410cc7a0} /* (29, 1, 11) {real, imag} */,
  {32'h40126db3, 32'h40db73a4} /* (29, 1, 10) {real, imag} */,
  {32'h409dd165, 32'h410d4d0a} /* (29, 1, 9) {real, imag} */,
  {32'h405e45ee, 32'h40d1ee00} /* (29, 1, 8) {real, imag} */,
  {32'h3f5c9f08, 32'h40c5c8a8} /* (29, 1, 7) {real, imag} */,
  {32'h4079cc94, 32'h40ca592f} /* (29, 1, 6) {real, imag} */,
  {32'h40313855, 32'hbf2d8496} /* (29, 1, 5) {real, imag} */,
  {32'hbfb0ce43, 32'hc0b09469} /* (29, 1, 4) {real, imag} */,
  {32'hc081cf32, 32'hc0ad8334} /* (29, 1, 3) {real, imag} */,
  {32'hc055396a, 32'hc0299013} /* (29, 1, 2) {real, imag} */,
  {32'hbf95143e, 32'hc04c8fea} /* (29, 1, 1) {real, imag} */,
  {32'hbe913799, 32'hc0286d07} /* (29, 1, 0) {real, imag} */,
  {32'hbf25587e, 32'hbf755ab3} /* (29, 0, 31) {real, imag} */,
  {32'hbfd90625, 32'hc0039709} /* (29, 0, 30) {real, imag} */,
  {32'hbf294938, 32'hc0310656} /* (29, 0, 29) {real, imag} */,
  {32'h3ee2f69b, 32'hbf993268} /* (29, 0, 28) {real, imag} */,
  {32'hbfce76a9, 32'hc01a830c} /* (29, 0, 27) {real, imag} */,
  {32'hbfdcdc88, 32'hc04a3fd8} /* (29, 0, 26) {real, imag} */,
  {32'hbe9194d2, 32'hc056ce43} /* (29, 0, 25) {real, imag} */,
  {32'h3f8926a2, 32'hc040f377} /* (29, 0, 24) {real, imag} */,
  {32'hbf398d3f, 32'hc01e98ef} /* (29, 0, 23) {real, imag} */,
  {32'h3c84dcc0, 32'hc00e36b7} /* (29, 0, 22) {real, imag} */,
  {32'h3f47b63e, 32'hbfce6d69} /* (29, 0, 21) {real, imag} */,
  {32'hc00952cb, 32'hbd8a98dc} /* (29, 0, 20) {real, imag} */,
  {32'hbfbca118, 32'hc000e4ca} /* (29, 0, 19) {real, imag} */,
  {32'hbf14cd99, 32'hc07354a8} /* (29, 0, 18) {real, imag} */,
  {32'hbfe994a8, 32'hc040bc88} /* (29, 0, 17) {real, imag} */,
  {32'hbf932fba, 32'hc007a172} /* (29, 0, 16) {real, imag} */,
  {32'h3f98dd81, 32'hbd9e1ec4} /* (29, 0, 15) {real, imag} */,
  {32'h3e29a290, 32'h406092da} /* (29, 0, 14) {real, imag} */,
  {32'h3efda7f6, 32'h40a99562} /* (29, 0, 13) {real, imag} */,
  {32'h40080915, 32'h408ac17c} /* (29, 0, 12) {real, imag} */,
  {32'h3fc7be93, 32'h401edb8a} /* (29, 0, 11) {real, imag} */,
  {32'h3f7f7c20, 32'h3f1830a2} /* (29, 0, 10) {real, imag} */,
  {32'h40119950, 32'h404137b4} /* (29, 0, 9) {real, imag} */,
  {32'h3fc88348, 32'h40453b65} /* (29, 0, 8) {real, imag} */,
  {32'h3fa82e97, 32'h40543dcb} /* (29, 0, 7) {real, imag} */,
  {32'h3ff9e7d7, 32'h4031e8f8} /* (29, 0, 6) {real, imag} */,
  {32'h3f4b4e2a, 32'hbf9996fb} /* (29, 0, 5) {real, imag} */,
  {32'hbd8b9742, 32'hc0537325} /* (29, 0, 4) {real, imag} */,
  {32'hbf69412a, 32'hc07f6a44} /* (29, 0, 3) {real, imag} */,
  {32'hbf7d2994, 32'hc071d448} /* (29, 0, 2) {real, imag} */,
  {32'hbf1bf15a, 32'hc00ee712} /* (29, 0, 1) {real, imag} */,
  {32'hbeb9f424, 32'hbef83b38} /* (29, 0, 0) {real, imag} */,
  {32'hbb2a1380, 32'hbfe55793} /* (28, 31, 31) {real, imag} */,
  {32'hbf90e643, 32'hc08b3cbe} /* (28, 31, 30) {real, imag} */,
  {32'hbff18948, 32'hc09a93bb} /* (28, 31, 29) {real, imag} */,
  {32'hc0111137, 32'hc0940d86} /* (28, 31, 28) {real, imag} */,
  {32'hbf8b6595, 32'hc04f7456} /* (28, 31, 27) {real, imag} */,
  {32'hbee810ca, 32'hc0492ab4} /* (28, 31, 26) {real, imag} */,
  {32'hbe184ac0, 32'hc070082b} /* (28, 31, 25) {real, imag} */,
  {32'hbeedb80c, 32'hc01c1d48} /* (28, 31, 24) {real, imag} */,
  {32'hbfa55d48, 32'hc01de1e0} /* (28, 31, 23) {real, imag} */,
  {32'hbfe326f3, 32'hbfdd8fb0} /* (28, 31, 22) {real, imag} */,
  {32'hbf24f4e7, 32'hc008b007} /* (28, 31, 21) {real, imag} */,
  {32'h3f460b86, 32'h3e333028} /* (28, 31, 20) {real, imag} */,
  {32'h3dcc10e6, 32'h40138e36} /* (28, 31, 19) {real, imag} */,
  {32'hbc029b18, 32'h40514078} /* (28, 31, 18) {real, imag} */,
  {32'hbce60810, 32'h40674750} /* (28, 31, 17) {real, imag} */,
  {32'hbf46230e, 32'h3f51c62e} /* (28, 31, 16) {real, imag} */,
  {32'hbed6b442, 32'h3fef3ef9} /* (28, 31, 15) {real, imag} */,
  {32'h3f6feee3, 32'h40703adc} /* (28, 31, 14) {real, imag} */,
  {32'h3e56eaca, 32'h3fd0d051} /* (28, 31, 13) {real, imag} */,
  {32'h3f1245c8, 32'h3fee9fb4} /* (28, 31, 12) {real, imag} */,
  {32'h3fc36aca, 32'h40425026} /* (28, 31, 11) {real, imag} */,
  {32'h3dd57516, 32'hbe4ae007} /* (28, 31, 10) {real, imag} */,
  {32'hbfef6c3a, 32'hc0274b40} /* (28, 31, 9) {real, imag} */,
  {32'hbf03cca6, 32'hbff60e7e} /* (28, 31, 8) {real, imag} */,
  {32'h3f4574ff, 32'hc0109768} /* (28, 31, 7) {real, imag} */,
  {32'h3ea04386, 32'hc0126892} /* (28, 31, 6) {real, imag} */,
  {32'hbfedc90c, 32'hc04fab11} /* (28, 31, 5) {real, imag} */,
  {32'hc0308aea, 32'hbfedadf2} /* (28, 31, 4) {real, imag} */,
  {32'hbf8a19d3, 32'hc03aaa7f} /* (28, 31, 3) {real, imag} */,
  {32'hbfbb08b9, 32'hc063a80d} /* (28, 31, 2) {real, imag} */,
  {32'hbeb3282a, 32'hc083d19b} /* (28, 31, 1) {real, imag} */,
  {32'h3db72ce0, 32'hbf86f732} /* (28, 31, 0) {real, imag} */,
  {32'hbdc034c8, 32'hc013bd4e} /* (28, 30, 31) {real, imag} */,
  {32'hbf07a3f6, 32'hc0b6c985} /* (28, 30, 30) {real, imag} */,
  {32'hc0156a5f, 32'hc0d50de8} /* (28, 30, 29) {real, imag} */,
  {32'hc025f80f, 32'hc0b662d6} /* (28, 30, 28) {real, imag} */,
  {32'hbf747d9c, 32'hc0a59a7a} /* (28, 30, 27) {real, imag} */,
  {32'hbe4f82f4, 32'hc0dd9762} /* (28, 30, 26) {real, imag} */,
  {32'hc00b6af0, 32'hc0baa496} /* (28, 30, 25) {real, imag} */,
  {32'hc010b3b6, 32'hc096e4a4} /* (28, 30, 24) {real, imag} */,
  {32'hc019ad80, 32'hc0983df3} /* (28, 30, 23) {real, imag} */,
  {32'hbf88fb76, 32'hc0aaba8b} /* (28, 30, 22) {real, imag} */,
  {32'h3e254958, 32'hc05e82f6} /* (28, 30, 21) {real, imag} */,
  {32'h4004878d, 32'h4094def8} /* (28, 30, 20) {real, imag} */,
  {32'h3e808c24, 32'h40bf083a} /* (28, 30, 19) {real, imag} */,
  {32'h3e9d3cb0, 32'h40d878d1} /* (28, 30, 18) {real, imag} */,
  {32'h3faa11d6, 32'h40eb3d2c} /* (28, 30, 17) {real, imag} */,
  {32'h3ea3113b, 32'h40a6342b} /* (28, 30, 16) {real, imag} */,
  {32'h3f19b7d0, 32'h40d5dc40} /* (28, 30, 15) {real, imag} */,
  {32'h4010b6e4, 32'h40f5aba5} /* (28, 30, 14) {real, imag} */,
  {32'h3e50516b, 32'h40a43b5d} /* (28, 30, 13) {real, imag} */,
  {32'h3f0cdaa8, 32'h407b3916} /* (28, 30, 12) {real, imag} */,
  {32'h3fd0ca79, 32'h409960eb} /* (28, 30, 11) {real, imag} */,
  {32'hbf92456a, 32'h3f78f616} /* (28, 30, 10) {real, imag} */,
  {32'hc0a974a2, 32'hc0992024} /* (28, 30, 9) {real, imag} */,
  {32'hc068fea2, 32'hc095a244} /* (28, 30, 8) {real, imag} */,
  {32'hc0048eaa, 32'hc096d4fe} /* (28, 30, 7) {real, imag} */,
  {32'hbfbbe76c, 32'hc0b281d4} /* (28, 30, 6) {real, imag} */,
  {32'hbf8e0f6a, 32'hc05749f6} /* (28, 30, 5) {real, imag} */,
  {32'hc0889d88, 32'hc085f3b7} /* (28, 30, 4) {real, imag} */,
  {32'hc0ae5a0d, 32'hc0aed984} /* (28, 30, 3) {real, imag} */,
  {32'hc040e772, 32'hc0c292fa} /* (28, 30, 2) {real, imag} */,
  {32'h40043288, 32'hc0cc3f6e} /* (28, 30, 1) {real, imag} */,
  {32'h3f005c94, 32'hc0509a90} /* (28, 30, 0) {real, imag} */,
  {32'hbf47c2ec, 32'hbfeade69} /* (28, 29, 31) {real, imag} */,
  {32'hc02496a6, 32'hc086ec38} /* (28, 29, 30) {real, imag} */,
  {32'hc087ba82, 32'hc0ab6893} /* (28, 29, 29) {real, imag} */,
  {32'hc046d46c, 32'hc05a19ae} /* (28, 29, 28) {real, imag} */,
  {32'hbfdf22df, 32'hc0634daf} /* (28, 29, 27) {real, imag} */,
  {32'hbfce3c82, 32'hc0b0fad6} /* (28, 29, 26) {real, imag} */,
  {32'hc02e0596, 32'hc08d2941} /* (28, 29, 25) {real, imag} */,
  {32'hc03cba01, 32'hc0c41a2c} /* (28, 29, 24) {real, imag} */,
  {32'hc06161b6, 32'hc0a8e8e4} /* (28, 29, 23) {real, imag} */,
  {32'hbf09144d, 32'hc0c2fb5e} /* (28, 29, 22) {real, imag} */,
  {32'hbfbf2ab7, 32'hc0011eac} /* (28, 29, 21) {real, imag} */,
  {32'h3f1c87fe, 32'h41085f15} /* (28, 29, 20) {real, imag} */,
  {32'h3fd82dce, 32'h40a3368a} /* (28, 29, 19) {real, imag} */,
  {32'h401c927a, 32'h4089cba2} /* (28, 29, 18) {real, imag} */,
  {32'h40396f4a, 32'h40dc199a} /* (28, 29, 17) {real, imag} */,
  {32'h3fdeb468, 32'h40cfdbfe} /* (28, 29, 16) {real, imag} */,
  {32'h3fc702f2, 32'h408fdfaa} /* (28, 29, 15) {real, imag} */,
  {32'h408e720c, 32'h40ce3d04} /* (28, 29, 14) {real, imag} */,
  {32'h40360b6c, 32'h40aedb02} /* (28, 29, 13) {real, imag} */,
  {32'h3f9bbc5d, 32'h403e5fe8} /* (28, 29, 12) {real, imag} */,
  {32'hbbdd3200, 32'h404eed4a} /* (28, 29, 11) {real, imag} */,
  {32'hbf6a4468, 32'hbf80b78a} /* (28, 29, 10) {real, imag} */,
  {32'hc0601efb, 32'hc0903ba1} /* (28, 29, 9) {real, imag} */,
  {32'hc09175f2, 32'hc0aeb010} /* (28, 29, 8) {real, imag} */,
  {32'hc08eb3ea, 32'hc0a18ea4} /* (28, 29, 7) {real, imag} */,
  {32'hc05a39ec, 32'hc084bd91} /* (28, 29, 6) {real, imag} */,
  {32'hbfbb9a0d, 32'hc0a210f5} /* (28, 29, 5) {real, imag} */,
  {32'hbfb0814f, 32'hc0ba5900} /* (28, 29, 4) {real, imag} */,
  {32'hc09cb02c, 32'hc0c1b964} /* (28, 29, 3) {real, imag} */,
  {32'hc093d571, 32'hc08d877d} /* (28, 29, 2) {real, imag} */,
  {32'hbf164c1d, 32'hc08f6657} /* (28, 29, 1) {real, imag} */,
  {32'hbd86e7c4, 32'hc064c9fa} /* (28, 29, 0) {real, imag} */,
  {32'hc016c7e0, 32'hbf25b102} /* (28, 28, 31) {real, imag} */,
  {32'hc0ab7c2b, 32'hc085a30a} /* (28, 28, 30) {real, imag} */,
  {32'hc0a61fc4, 32'hc0e85491} /* (28, 28, 29) {real, imag} */,
  {32'hbfa71630, 32'hc0ca9aea} /* (28, 28, 28) {real, imag} */,
  {32'hc02e86b9, 32'hc065476b} /* (28, 28, 27) {real, imag} */,
  {32'hc078dbec, 32'hc0b20909} /* (28, 28, 26) {real, imag} */,
  {32'hbfc18f70, 32'hc0a0f07a} /* (28, 28, 25) {real, imag} */,
  {32'hbf4a4dd7, 32'hc0988319} /* (28, 28, 24) {real, imag} */,
  {32'hc007a982, 32'hc06897b5} /* (28, 28, 23) {real, imag} */,
  {32'hbf610d54, 32'hc0987f84} /* (28, 28, 22) {real, imag} */,
  {32'hc08a8d4b, 32'hc06010b9} /* (28, 28, 21) {real, imag} */,
  {32'hbea3f1e3, 32'h409dde1f} /* (28, 28, 20) {real, imag} */,
  {32'h408a37d7, 32'h405b1728} /* (28, 28, 19) {real, imag} */,
  {32'h40e01572, 32'h40848f96} /* (28, 28, 18) {real, imag} */,
  {32'h40a69e65, 32'h40ba0cd5} /* (28, 28, 17) {real, imag} */,
  {32'h403efab7, 32'h40447d1b} /* (28, 28, 16) {real, imag} */,
  {32'h40274cd4, 32'hbf8e8b4d} /* (28, 28, 15) {real, imag} */,
  {32'h40488b07, 32'h4073afa8} /* (28, 28, 14) {real, imag} */,
  {32'h4050fc47, 32'h405bd2ae} /* (28, 28, 13) {real, imag} */,
  {32'h40291dc4, 32'h40031ab8} /* (28, 28, 12) {real, imag} */,
  {32'hbdc27239, 32'h405088d4} /* (28, 28, 11) {real, imag} */,
  {32'hc0426f54, 32'hc05bfde2} /* (28, 28, 10) {real, imag} */,
  {32'hc0743e51, 32'hc095fc97} /* (28, 28, 9) {real, imag} */,
  {32'hbfee131e, 32'hc0967b94} /* (28, 28, 8) {real, imag} */,
  {32'hc054cec0, 32'hc0a61689} /* (28, 28, 7) {real, imag} */,
  {32'hc07ca72c, 32'hc0192f76} /* (28, 28, 6) {real, imag} */,
  {32'hc053d66a, 32'hc0655256} /* (28, 28, 5) {real, imag} */,
  {32'hc01aa901, 32'hc0782550} /* (28, 28, 4) {real, imag} */,
  {32'hc056480b, 32'hc08f1f36} /* (28, 28, 3) {real, imag} */,
  {32'hc0a09c37, 32'hc026859a} /* (28, 28, 2) {real, imag} */,
  {32'hc055a9f9, 32'hbfcd5630} /* (28, 28, 1) {real, imag} */,
  {32'hbf9f8c05, 32'hbf9fa1f4} /* (28, 28, 0) {real, imag} */,
  {32'hbf169ff6, 32'hc008b328} /* (28, 27, 31) {real, imag} */,
  {32'hc09cbe4e, 32'hc0a9d4a4} /* (28, 27, 30) {real, imag} */,
  {32'hc0caa516, 32'hc09921f5} /* (28, 27, 29) {real, imag} */,
  {32'hc025eef4, 32'hc01de5d0} /* (28, 27, 28) {real, imag} */,
  {32'hc0628fe0, 32'h3d132b08} /* (28, 27, 27) {real, imag} */,
  {32'hc06a927a, 32'hc08ce195} /* (28, 27, 26) {real, imag} */,
  {32'hbea2df6d, 32'hc0c4c861} /* (28, 27, 25) {real, imag} */,
  {32'h3feab81e, 32'hc06061a2} /* (28, 27, 24) {real, imag} */,
  {32'h3e0caf6f, 32'hc032e1c7} /* (28, 27, 23) {real, imag} */,
  {32'hc028eed8, 32'hc0aaccda} /* (28, 27, 22) {real, imag} */,
  {32'hc02c8fcc, 32'hc0d207ff} /* (28, 27, 21) {real, imag} */,
  {32'hbdcd27b0, 32'h400c4e4e} /* (28, 27, 20) {real, imag} */,
  {32'h40803974, 32'h4086525b} /* (28, 27, 19) {real, imag} */,
  {32'h40e95260, 32'h407b7c08} /* (28, 27, 18) {real, imag} */,
  {32'h40574d74, 32'h4047c8e4} /* (28, 27, 17) {real, imag} */,
  {32'h400fbcc6, 32'h403fb99c} /* (28, 27, 16) {real, imag} */,
  {32'h3f0c9959, 32'h3fbd191e} /* (28, 27, 15) {real, imag} */,
  {32'h3eb15fb4, 32'h40946206} /* (28, 27, 14) {real, imag} */,
  {32'hbe92c52a, 32'h40aa950a} /* (28, 27, 13) {real, imag} */,
  {32'h3fa519f4, 32'h404ce1a0} /* (28, 27, 12) {real, imag} */,
  {32'h3feae9ca, 32'h4073678e} /* (28, 27, 11) {real, imag} */,
  {32'hbeb0378c, 32'hc088142a} /* (28, 27, 10) {real, imag} */,
  {32'hc081bfd1, 32'hc0c23e38} /* (28, 27, 9) {real, imag} */,
  {32'hc03fe1e6, 32'hc09307cc} /* (28, 27, 8) {real, imag} */,
  {32'hc040192a, 32'hc09e8c84} /* (28, 27, 7) {real, imag} */,
  {32'hc03d3ca2, 32'hc099bb48} /* (28, 27, 6) {real, imag} */,
  {32'hc007f916, 32'hc0913fd5} /* (28, 27, 5) {real, imag} */,
  {32'hc030c9cf, 32'hc0356a6a} /* (28, 27, 4) {real, imag} */,
  {32'hc0800b18, 32'hc06a34f1} /* (28, 27, 3) {real, imag} */,
  {32'hc03ce924, 32'hc05c81e2} /* (28, 27, 2) {real, imag} */,
  {32'hbfac887f, 32'hc0008524} /* (28, 27, 1) {real, imag} */,
  {32'hbe566e50, 32'h3f43e9b6} /* (28, 27, 0) {real, imag} */,
  {32'hbfd5c54c, 32'hbfebb8d8} /* (28, 26, 31) {real, imag} */,
  {32'hc097cb72, 32'hc0756506} /* (28, 26, 30) {real, imag} */,
  {32'hc06bd624, 32'hc0902e08} /* (28, 26, 29) {real, imag} */,
  {32'hbeb9e438, 32'hc0950e7a} /* (28, 26, 28) {real, imag} */,
  {32'hc04c131f, 32'hc05af4a0} /* (28, 26, 27) {real, imag} */,
  {32'hc086f3be, 32'hc0928714} /* (28, 26, 26) {real, imag} */,
  {32'hbfeaa5c6, 32'hc0908790} /* (28, 26, 25) {real, imag} */,
  {32'h3fd56e5f, 32'hbf62958b} /* (28, 26, 24) {real, imag} */,
  {32'h3f46e86a, 32'hc012815d} /* (28, 26, 23) {real, imag} */,
  {32'hbfc93e91, 32'hc06cf66e} /* (28, 26, 22) {real, imag} */,
  {32'hbdf04118, 32'hc06c533c} /* (28, 26, 21) {real, imag} */,
  {32'h3f7fad97, 32'h404fb3a2} /* (28, 26, 20) {real, imag} */,
  {32'h3fb08e5a, 32'h405ab486} /* (28, 26, 19) {real, imag} */,
  {32'h4033323a, 32'h40140fb6} /* (28, 26, 18) {real, imag} */,
  {32'h3fce4922, 32'h3fd2c397} /* (28, 26, 17) {real, imag} */,
  {32'h40437fd0, 32'h4095fbca} /* (28, 26, 16) {real, imag} */,
  {32'hbd59a328, 32'h406e9d5a} /* (28, 26, 15) {real, imag} */,
  {32'hbfb23083, 32'h40a7d15c} /* (28, 26, 14) {real, imag} */,
  {32'hbfdc182e, 32'h40babf64} /* (28, 26, 13) {real, imag} */,
  {32'hbe23c0f3, 32'h40970b3c} /* (28, 26, 12) {real, imag} */,
  {32'h3fe8af80, 32'h40696bc0} /* (28, 26, 11) {real, imag} */,
  {32'h3f713c70, 32'hbfbcd5bd} /* (28, 26, 10) {real, imag} */,
  {32'hc0807cf0, 32'hc04a415a} /* (28, 26, 9) {real, imag} */,
  {32'hc074fb93, 32'hc0bad20f} /* (28, 26, 8) {real, imag} */,
  {32'hbf98a13c, 32'hc0bf9a9e} /* (28, 26, 7) {real, imag} */,
  {32'hbfdd403a, 32'hc0bab092} /* (28, 26, 6) {real, imag} */,
  {32'hbfbea09f, 32'hc0b68e2c} /* (28, 26, 5) {real, imag} */,
  {32'hbfbd60a2, 32'hc041086a} /* (28, 26, 4) {real, imag} */,
  {32'hc0391268, 32'hc08961f5} /* (28, 26, 3) {real, imag} */,
  {32'hbff74f58, 32'hc09e7692} /* (28, 26, 2) {real, imag} */,
  {32'hbfe1cc50, 32'hc0a33945} /* (28, 26, 1) {real, imag} */,
  {32'hbf817817, 32'hbfe02d97} /* (28, 26, 0) {real, imag} */,
  {32'hbfeea039, 32'hc0715f54} /* (28, 25, 31) {real, imag} */,
  {32'hc0932852, 32'hc0c9f1be} /* (28, 25, 30) {real, imag} */,
  {32'hc0959131, 32'hc0664a66} /* (28, 25, 29) {real, imag} */,
  {32'h3ed68204, 32'hc07cdc56} /* (28, 25, 28) {real, imag} */,
  {32'hbe245276, 32'hc101a504} /* (28, 25, 27) {real, imag} */,
  {32'hbf016e98, 32'hc1125cb6} /* (28, 25, 26) {real, imag} */,
  {32'hc06117c8, 32'hc0abaf5f} /* (28, 25, 25) {real, imag} */,
  {32'hc00c791c, 32'hc038bf4f} /* (28, 25, 24) {real, imag} */,
  {32'hbe860814, 32'hc082ef2e} /* (28, 25, 23) {real, imag} */,
  {32'h3ee53bd4, 32'hc0a5300d} /* (28, 25, 22) {real, imag} */,
  {32'h401eb90b, 32'hbfe43bed} /* (28, 25, 21) {real, imag} */,
  {32'h4064b7f4, 32'h4100116a} /* (28, 25, 20) {real, imag} */,
  {32'h3f5cced5, 32'h4100324b} /* (28, 25, 19) {real, imag} */,
  {32'h3f0e2af6, 32'h40593e39} /* (28, 25, 18) {real, imag} */,
  {32'h3fda8bce, 32'h3fc881fb} /* (28, 25, 17) {real, imag} */,
  {32'h407f1270, 32'h4084330a} /* (28, 25, 16) {real, imag} */,
  {32'h3f29b61f, 32'h40902648} /* (28, 25, 15) {real, imag} */,
  {32'hbf3204ac, 32'h40ca1779} /* (28, 25, 14) {real, imag} */,
  {32'h3ec98a7a, 32'h41045d61} /* (28, 25, 13) {real, imag} */,
  {32'h3f1401e6, 32'h40ebbc4f} /* (28, 25, 12) {real, imag} */,
  {32'h3e81a4ed, 32'h4068939b} /* (28, 25, 11) {real, imag} */,
  {32'hbf84696c, 32'hbfc04698} /* (28, 25, 10) {real, imag} */,
  {32'hc0a4b30a, 32'hc0977de6} /* (28, 25, 9) {real, imag} */,
  {32'hc07508df, 32'hc0b65d29} /* (28, 25, 8) {real, imag} */,
  {32'hbeab72f6, 32'hc0a0578a} /* (28, 25, 7) {real, imag} */,
  {32'hbe0b4f58, 32'hc063840e} /* (28, 25, 6) {real, imag} */,
  {32'hbf25cbaa, 32'hc08c64da} /* (28, 25, 5) {real, imag} */,
  {32'hc02883ba, 32'hc02846ce} /* (28, 25, 4) {real, imag} */,
  {32'hc033c344, 32'hc04c9c8d} /* (28, 25, 3) {real, imag} */,
  {32'hbead1c86, 32'hc06e262e} /* (28, 25, 2) {real, imag} */,
  {32'hbfa1bd32, 32'hc0f280d4} /* (28, 25, 1) {real, imag} */,
  {32'hbf8f893a, 32'hc08a629e} /* (28, 25, 0) {real, imag} */,
  {32'hbf6fe70a, 32'hc0b03064} /* (28, 24, 31) {real, imag} */,
  {32'hbf2921ef, 32'hc0c7ec20} /* (28, 24, 30) {real, imag} */,
  {32'hbfab73b4, 32'hc06c7136} /* (28, 24, 29) {real, imag} */,
  {32'h3edf5b6e, 32'hc09685ca} /* (28, 24, 28) {real, imag} */,
  {32'hbfc7b1ba, 32'hc026c2f8} /* (28, 24, 27) {real, imag} */,
  {32'hc0377e28, 32'hc0d686ab} /* (28, 24, 26) {real, imag} */,
  {32'hc091dd84, 32'hc0ef1046} /* (28, 24, 25) {real, imag} */,
  {32'hc05f876d, 32'hc0d0375b} /* (28, 24, 24) {real, imag} */,
  {32'hbf24dfac, 32'hc0eaa6ec} /* (28, 24, 23) {real, imag} */,
  {32'hbf96c9e6, 32'hc1011bd1} /* (28, 24, 22) {real, imag} */,
  {32'hbf9ea10f, 32'hc039f105} /* (28, 24, 21) {real, imag} */,
  {32'h3fce41ec, 32'h40becf6b} /* (28, 24, 20) {real, imag} */,
  {32'h3eea9b16, 32'h409a42f4} /* (28, 24, 19) {real, imag} */,
  {32'h3fbb76a7, 32'h4054aff6} /* (28, 24, 18) {real, imag} */,
  {32'h4080c10f, 32'h40a3bda8} /* (28, 24, 17) {real, imag} */,
  {32'h401dacf0, 32'h409a09d2} /* (28, 24, 16) {real, imag} */,
  {32'hbd28e638, 32'h405a4ca3} /* (28, 24, 15) {real, imag} */,
  {32'h404c733e, 32'h40e83cb6} /* (28, 24, 14) {real, imag} */,
  {32'h4037bbe3, 32'h410625d3} /* (28, 24, 13) {real, imag} */,
  {32'h3f7c02a8, 32'h4060e198} /* (28, 24, 12) {real, imag} */,
  {32'h3e23f470, 32'h3ff20748} /* (28, 24, 11) {real, imag} */,
  {32'hbfea4ac2, 32'hc0418c38} /* (28, 24, 10) {real, imag} */,
  {32'hc082fd76, 32'hc0c5936e} /* (28, 24, 9) {real, imag} */,
  {32'hc095ff48, 32'hc09ee504} /* (28, 24, 8) {real, imag} */,
  {32'hc03aeeec, 32'hc057d958} /* (28, 24, 7) {real, imag} */,
  {32'hbd833ff0, 32'hc0442b3a} /* (28, 24, 6) {real, imag} */,
  {32'hbf11c679, 32'hc0c1b09f} /* (28, 24, 5) {real, imag} */,
  {32'hbfd37f0e, 32'hc0a8905e} /* (28, 24, 4) {real, imag} */,
  {32'hc023cb79, 32'hc0ae6df0} /* (28, 24, 3) {real, imag} */,
  {32'hbf13da50, 32'hc09d0a9c} /* (28, 24, 2) {real, imag} */,
  {32'hbf824eb2, 32'hc0ecc0f4} /* (28, 24, 1) {real, imag} */,
  {32'hbf49ef68, 32'hc0936584} /* (28, 24, 0) {real, imag} */,
  {32'hbf856529, 32'hc08d8594} /* (28, 23, 31) {real, imag} */,
  {32'hbf257b7e, 32'hc0b29cd6} /* (28, 23, 30) {real, imag} */,
  {32'hbf134114, 32'hc0b242e9} /* (28, 23, 29) {real, imag} */,
  {32'hbf2baf05, 32'hc09ef4c8} /* (28, 23, 28) {real, imag} */,
  {32'hc04fd332, 32'hc01e6eb1} /* (28, 23, 27) {real, imag} */,
  {32'hc0bcc9ca, 32'hc0a4bf30} /* (28, 23, 26) {real, imag} */,
  {32'hc0466fb0, 32'hc0c99a8e} /* (28, 23, 25) {real, imag} */,
  {32'hbe99fae7, 32'hc0a0108e} /* (28, 23, 24) {real, imag} */,
  {32'hbfdaa9a2, 32'hc0b685ae} /* (28, 23, 23) {real, imag} */,
  {32'hc01057ed, 32'hc0d906ca} /* (28, 23, 22) {real, imag} */,
  {32'hbe46fd90, 32'hc04700da} /* (28, 23, 21) {real, imag} */,
  {32'h40157965, 32'h403f5b5a} /* (28, 23, 20) {real, imag} */,
  {32'h3f750364, 32'h4007953c} /* (28, 23, 19) {real, imag} */,
  {32'h402d4c63, 32'h402fd7e0} /* (28, 23, 18) {real, imag} */,
  {32'h4027655c, 32'h40a85842} /* (28, 23, 17) {real, imag} */,
  {32'h3f9e9bee, 32'h40c1e3fb} /* (28, 23, 16) {real, imag} */,
  {32'h40026fb4, 32'h40b81080} /* (28, 23, 15) {real, imag} */,
  {32'h402209a2, 32'h40e4d275} /* (28, 23, 14) {real, imag} */,
  {32'h3f2be564, 32'h40d8c63d} /* (28, 23, 13) {real, imag} */,
  {32'h3f31c713, 32'h40533152} /* (28, 23, 12) {real, imag} */,
  {32'h3fb3247c, 32'h401bfeb2} /* (28, 23, 11) {real, imag} */,
  {32'h3f877d8a, 32'hbf819d98} /* (28, 23, 10) {real, imag} */,
  {32'h3c866b70, 32'hc08a86cd} /* (28, 23, 9) {real, imag} */,
  {32'hc023eb7f, 32'hc08e00da} /* (28, 23, 8) {real, imag} */,
  {32'hbf9c9340, 32'hc00bf10b} /* (28, 23, 7) {real, imag} */,
  {32'hbe76d970, 32'hc0513e52} /* (28, 23, 6) {real, imag} */,
  {32'hbf4beec5, 32'hc0ee7801} /* (28, 23, 5) {real, imag} */,
  {32'hbebd4834, 32'hc09da75c} /* (28, 23, 4) {real, imag} */,
  {32'h3feaea31, 32'hc06b0a30} /* (28, 23, 3) {real, imag} */,
  {32'hbe9a50d9, 32'hc0b10610} /* (28, 23, 2) {real, imag} */,
  {32'hbff43eba, 32'hc0b5def8} /* (28, 23, 1) {real, imag} */,
  {32'hbfad80cd, 32'hc0519d5b} /* (28, 23, 0) {real, imag} */,
  {32'hc04f5c96, 32'hc0630b19} /* (28, 22, 31) {real, imag} */,
  {32'hbfbf13a2, 32'hc0788804} /* (28, 22, 30) {real, imag} */,
  {32'hbf35d336, 32'hc09c72ea} /* (28, 22, 29) {real, imag} */,
  {32'hc007d5d8, 32'hc0d48d26} /* (28, 22, 28) {real, imag} */,
  {32'hbfcc8be0, 32'hc10085a0} /* (28, 22, 27) {real, imag} */,
  {32'hc0308f7a, 32'hc0ad62e5} /* (28, 22, 26) {real, imag} */,
  {32'hbf8e92c8, 32'hc0421cef} /* (28, 22, 25) {real, imag} */,
  {32'hbe85756e, 32'hc0959b15} /* (28, 22, 24) {real, imag} */,
  {32'hbf837aa1, 32'hc0e5b0ac} /* (28, 22, 23) {real, imag} */,
  {32'hc05b26a7, 32'hc0dcda19} /* (28, 22, 22) {real, imag} */,
  {32'h3f2fe722, 32'hc053de04} /* (28, 22, 21) {real, imag} */,
  {32'h4071e552, 32'hbf15256a} /* (28, 22, 20) {real, imag} */,
  {32'h3f9c7d00, 32'hbf185e81} /* (28, 22, 19) {real, imag} */,
  {32'h3fd75238, 32'h3fdfcaa8} /* (28, 22, 18) {real, imag} */,
  {32'h3f9314ac, 32'h40c519e7} /* (28, 22, 17) {real, imag} */,
  {32'h3fd433fd, 32'h40d0f9ae} /* (28, 22, 16) {real, imag} */,
  {32'h3fc57ba9, 32'h40c17e48} /* (28, 22, 15) {real, imag} */,
  {32'hbb4733c0, 32'h40c3b0f6} /* (28, 22, 14) {real, imag} */,
  {32'h3ff40b98, 32'h40ac474d} /* (28, 22, 13) {real, imag} */,
  {32'h404ce806, 32'h40bf7bc2} /* (28, 22, 12) {real, imag} */,
  {32'h407bcae6, 32'h40913555} /* (28, 22, 11) {real, imag} */,
  {32'h404d96d0, 32'hc0010cec} /* (28, 22, 10) {real, imag} */,
  {32'hbecf8556, 32'hc0ff9e2a} /* (28, 22, 9) {real, imag} */,
  {32'hbfc8b5ed, 32'hc113ccfc} /* (28, 22, 8) {real, imag} */,
  {32'hbfe97b96, 32'hc0cab56b} /* (28, 22, 7) {real, imag} */,
  {32'hbf52bac6, 32'hc070eea1} /* (28, 22, 6) {real, imag} */,
  {32'hbef83099, 32'hc0e3c8fc} /* (28, 22, 5) {real, imag} */,
  {32'hbeecec14, 32'hc09cf7db} /* (28, 22, 4) {real, imag} */,
  {32'h3f56f27c, 32'hbfbc6ef2} /* (28, 22, 3) {real, imag} */,
  {32'hbe98295a, 32'hc0977c84} /* (28, 22, 2) {real, imag} */,
  {32'hbf95ccb2, 32'hc072bfe8} /* (28, 22, 1) {real, imag} */,
  {32'hc00fae0a, 32'hbffad31e} /* (28, 22, 0) {real, imag} */,
  {32'hbf86d980, 32'hc026f694} /* (28, 21, 31) {real, imag} */,
  {32'hbf2e52ff, 32'hc0858314} /* (28, 21, 30) {real, imag} */,
  {32'hc0199b30, 32'hbfdb6894} /* (28, 21, 29) {real, imag} */,
  {32'hc05817fe, 32'hc0578f66} /* (28, 21, 28) {real, imag} */,
  {32'hbf8ab0bc, 32'hc0d58741} /* (28, 21, 27) {real, imag} */,
  {32'h3fcccf00, 32'hc05159dc} /* (28, 21, 26) {real, imag} */,
  {32'hbe807315, 32'hbfb9d74c} /* (28, 21, 25) {real, imag} */,
  {32'hc051f121, 32'hc057cd55} /* (28, 21, 24) {real, imag} */,
  {32'h3f516faf, 32'hc08b8716} /* (28, 21, 23) {real, imag} */,
  {32'hbe0c3ff1, 32'hc0113750} /* (28, 21, 22) {real, imag} */,
  {32'hbf20065e, 32'h3f40e47c} /* (28, 21, 21) {real, imag} */,
  {32'hbe3c72af, 32'hbf781422} /* (28, 21, 20) {real, imag} */,
  {32'hbfb34cd4, 32'hbf4306ca} /* (28, 21, 19) {real, imag} */,
  {32'hbe9527c0, 32'h400ca6b6} /* (28, 21, 18) {real, imag} */,
  {32'h3f07751a, 32'h409c8d9c} /* (28, 21, 17) {real, imag} */,
  {32'h3fe89a26, 32'h409f54f0} /* (28, 21, 16) {real, imag} */,
  {32'h3f3fe40e, 32'h402bbe4a} /* (28, 21, 15) {real, imag} */,
  {32'hbf5c44a5, 32'h3fbb9d47} /* (28, 21, 14) {real, imag} */,
  {32'h3f8d7080, 32'h3fae431c} /* (28, 21, 13) {real, imag} */,
  {32'h3fda3c8c, 32'h3ebd6096} /* (28, 21, 12) {real, imag} */,
  {32'h3dfeab74, 32'h3b862fc0} /* (28, 21, 11) {real, imag} */,
  {32'hbee60ea4, 32'hbfbd814d} /* (28, 21, 10) {real, imag} */,
  {32'hbfda77f2, 32'hc104b877} /* (28, 21, 9) {real, imag} */,
  {32'hc00a23b7, 32'hc102e422} /* (28, 21, 8) {real, imag} */,
  {32'hbfce30c7, 32'hc089764b} /* (28, 21, 7) {real, imag} */,
  {32'hbed94aa3, 32'h3f7c2a1f} /* (28, 21, 6) {real, imag} */,
  {32'hbfa85e3c, 32'h3f34f66d} /* (28, 21, 5) {real, imag} */,
  {32'hbfacddda, 32'hbfeef9dc} /* (28, 21, 4) {real, imag} */,
  {32'hbf8b2bd6, 32'hbf44af87} /* (28, 21, 3) {real, imag} */,
  {32'hbe02090e, 32'hbef73d12} /* (28, 21, 2) {real, imag} */,
  {32'hbd1d5630, 32'hbf88c5aa} /* (28, 21, 1) {real, imag} */,
  {32'hbf4242ea, 32'hbd221440} /* (28, 21, 0) {real, imag} */,
  {32'h3f195046, 32'h3f484645} /* (28, 20, 31) {real, imag} */,
  {32'h3e9346e2, 32'hbf85a9fd} /* (28, 20, 30) {real, imag} */,
  {32'hbf122617, 32'h404a9985} /* (28, 20, 29) {real, imag} */,
  {32'hbf6f7e65, 32'h40bb60f4} /* (28, 20, 28) {real, imag} */,
  {32'hc00543ad, 32'h407549b2} /* (28, 20, 27) {real, imag} */,
  {32'h3fa01c37, 32'h40299cac} /* (28, 20, 26) {real, imag} */,
  {32'h40169192, 32'h403c928d} /* (28, 20, 25) {real, imag} */,
  {32'h3eef75a2, 32'h4070a94a} /* (28, 20, 24) {real, imag} */,
  {32'h3ff24446, 32'h40bc48f0} /* (28, 20, 23) {real, imag} */,
  {32'h40815946, 32'h40b2fbac} /* (28, 20, 22) {real, imag} */,
  {32'h3f18fdc5, 32'h400d48df} /* (28, 20, 21) {real, imag} */,
  {32'hc005cdfd, 32'hc02ae7c6} /* (28, 20, 20) {real, imag} */,
  {32'hc07ddc20, 32'hbfe6fb64} /* (28, 20, 19) {real, imag} */,
  {32'hc06ba4bf, 32'hbfe094ad} /* (28, 20, 18) {real, imag} */,
  {32'hbfec15ea, 32'h3e794bf4} /* (28, 20, 17) {real, imag} */,
  {32'hc008f951, 32'h3f3f44ff} /* (28, 20, 16) {real, imag} */,
  {32'hc0240404, 32'hc0847555} /* (28, 20, 15) {real, imag} */,
  {32'hbf8c0851, 32'hc0cc8308} /* (28, 20, 14) {real, imag} */,
  {32'h3f820389, 32'hc09b94f6} /* (28, 20, 13) {real, imag} */,
  {32'h3f17410f, 32'hc0d2bb36} /* (28, 20, 12) {real, imag} */,
  {32'hbfb6134f, 32'hc0a8d832} /* (28, 20, 11) {real, imag} */,
  {32'hc008d79f, 32'h3e6eaab7} /* (28, 20, 10) {real, imag} */,
  {32'h3f940372, 32'hbe22c148} /* (28, 20, 9) {real, imag} */,
  {32'h3fb9f7cb, 32'h40529b25} /* (28, 20, 8) {real, imag} */,
  {32'h3eb95997, 32'h40a9431e} /* (28, 20, 7) {real, imag} */,
  {32'h3f001623, 32'h40b1bc02} /* (28, 20, 6) {real, imag} */,
  {32'h3f0f8a65, 32'h40491458} /* (28, 20, 5) {real, imag} */,
  {32'h3f8d12ca, 32'h40510e5c} /* (28, 20, 4) {real, imag} */,
  {32'h3fb2834f, 32'h4085aeb2} /* (28, 20, 3) {real, imag} */,
  {32'h40358db0, 32'h40a3ab8c} /* (28, 20, 2) {real, imag} */,
  {32'h3fe12170, 32'h4076e4b9} /* (28, 20, 1) {real, imag} */,
  {32'h3f4b62a3, 32'h4048607a} /* (28, 20, 0) {real, imag} */,
  {32'h3fd8f79d, 32'h3ffca8ad} /* (28, 19, 31) {real, imag} */,
  {32'h402b927d, 32'h3fc47ab4} /* (28, 19, 30) {real, imag} */,
  {32'h3fd26972, 32'h404d1f44} /* (28, 19, 29) {real, imag} */,
  {32'hc0114250, 32'h40b9cd5c} /* (28, 19, 28) {real, imag} */,
  {32'hbe41540e, 32'h40ccac62} /* (28, 19, 27) {real, imag} */,
  {32'h3f92ff1c, 32'h40a86a4e} /* (28, 19, 26) {real, imag} */,
  {32'h3e9f85ae, 32'h40edb42a} /* (28, 19, 25) {real, imag} */,
  {32'h3e922ae7, 32'h40ef8a1e} /* (28, 19, 24) {real, imag} */,
  {32'h402a8cb7, 32'h40e6680d} /* (28, 19, 23) {real, imag} */,
  {32'h409b5e3c, 32'h40bcd85f} /* (28, 19, 22) {real, imag} */,
  {32'h405e5822, 32'h3faa3b94} /* (28, 19, 21) {real, imag} */,
  {32'h3f225fb6, 32'hc0ac6ca1} /* (28, 19, 20) {real, imag} */,
  {32'hbf8a1ed8, 32'hc0d6bcdc} /* (28, 19, 19) {real, imag} */,
  {32'hbfa246ba, 32'hc0fc0577} /* (28, 19, 18) {real, imag} */,
  {32'h3fb4f2d8, 32'hc0a84ee5} /* (28, 19, 17) {real, imag} */,
  {32'h3ef61188, 32'hbefdfc43} /* (28, 19, 16) {real, imag} */,
  {32'hbe3e73d8, 32'hc02fa427} /* (28, 19, 15) {real, imag} */,
  {32'h3f8d4f65, 32'hc07eaf27} /* (28, 19, 14) {real, imag} */,
  {32'h400194ed, 32'hc0952e8a} /* (28, 19, 13) {real, imag} */,
  {32'h3e43d0a8, 32'hc0ecd1ee} /* (28, 19, 12) {real, imag} */,
  {32'hbfc1436e, 32'hc0b9dc85} /* (28, 19, 11) {real, imag} */,
  {32'hbe2d29c4, 32'h40060f48} /* (28, 19, 10) {real, imag} */,
  {32'h3f365377, 32'h40a835ba} /* (28, 19, 9) {real, imag} */,
  {32'hbe4172ea, 32'h4104071c} /* (28, 19, 8) {real, imag} */,
  {32'h3fc3e328, 32'h40f85663} /* (28, 19, 7) {real, imag} */,
  {32'h3fedbc78, 32'h40093458} /* (28, 19, 6) {real, imag} */,
  {32'h408d83c8, 32'h3e55b1d0} /* (28, 19, 5) {real, imag} */,
  {32'h401cf4aa, 32'h407f3e7a} /* (28, 19, 4) {real, imag} */,
  {32'h3e0340aa, 32'h409bb1c1} /* (28, 19, 3) {real, imag} */,
  {32'h40476878, 32'h409983d2} /* (28, 19, 2) {real, imag} */,
  {32'h4021157a, 32'h40e62c16} /* (28, 19, 1) {real, imag} */,
  {32'h3fe43afd, 32'h40a2221b} /* (28, 19, 0) {real, imag} */,
  {32'h3f8f60c8, 32'h407ee72b} /* (28, 18, 31) {real, imag} */,
  {32'h401597a8, 32'h408dc00e} /* (28, 18, 30) {real, imag} */,
  {32'h403e7efe, 32'h3fc16ac4} /* (28, 18, 29) {real, imag} */,
  {32'h3f959319, 32'h3fadb0a4} /* (28, 18, 28) {real, imag} */,
  {32'h40636dcc, 32'h408d502c} /* (28, 18, 27) {real, imag} */,
  {32'h4045450d, 32'h40aacbcb} /* (28, 18, 26) {real, imag} */,
  {32'h3f742d54, 32'h409fb03b} /* (28, 18, 25) {real, imag} */,
  {32'h3fc8d634, 32'h40ac40c8} /* (28, 18, 24) {real, imag} */,
  {32'h403c5948, 32'h408d025e} /* (28, 18, 23) {real, imag} */,
  {32'h4099ee2e, 32'h40742e95} /* (28, 18, 22) {real, imag} */,
  {32'h409d3f51, 32'h3dc9c858} /* (28, 18, 21) {real, imag} */,
  {32'h3fda04a6, 32'hc0cb9846} /* (28, 18, 20) {real, imag} */,
  {32'hbfff6f9c, 32'hc0dc69ac} /* (28, 18, 19) {real, imag} */,
  {32'hc059d9fa, 32'hc0e4b872} /* (28, 18, 18) {real, imag} */,
  {32'h3f804285, 32'hc0efed22} /* (28, 18, 17) {real, imag} */,
  {32'h4089780f, 32'hc014a00c} /* (28, 18, 16) {real, imag} */,
  {32'h4019b0ac, 32'hbfaccb05} /* (28, 18, 15) {real, imag} */,
  {32'h3e5ba62a, 32'hc066c0bc} /* (28, 18, 14) {real, imag} */,
  {32'hbf867339, 32'hc0aded96} /* (28, 18, 13) {real, imag} */,
  {32'h3f956954, 32'hc0ba0d74} /* (28, 18, 12) {real, imag} */,
  {32'hbe8e8470, 32'hc09f22f4} /* (28, 18, 11) {real, imag} */,
  {32'h3ff72bfc, 32'h406a1f90} /* (28, 18, 10) {real, imag} */,
  {32'h40303042, 32'h4105f7fe} /* (28, 18, 9) {real, imag} */,
  {32'h3c0d4558, 32'h40dc7d48} /* (28, 18, 8) {real, imag} */,
  {32'h3fa4e7a2, 32'h4092a322} /* (28, 18, 7) {real, imag} */,
  {32'h3ff88099, 32'h3f8f8be9} /* (28, 18, 6) {real, imag} */,
  {32'h3ffc2836, 32'h3ea030f0} /* (28, 18, 5) {real, imag} */,
  {32'h3f74c3b0, 32'h4061ffee} /* (28, 18, 4) {real, imag} */,
  {32'h3e5d8734, 32'h40775aae} /* (28, 18, 3) {real, imag} */,
  {32'h4031b714, 32'h408972b1} /* (28, 18, 2) {real, imag} */,
  {32'h3f23ce58, 32'h40971cb3} /* (28, 18, 1) {real, imag} */,
  {32'h3e6edea8, 32'h4094d72c} /* (28, 18, 0) {real, imag} */,
  {32'h3f06d937, 32'h406c9fa4} /* (28, 17, 31) {real, imag} */,
  {32'h3f137066, 32'h40cdc758} /* (28, 17, 30) {real, imag} */,
  {32'h403df83c, 32'h40900445} /* (28, 17, 29) {real, imag} */,
  {32'h4098c18a, 32'h40234d47} /* (28, 17, 28) {real, imag} */,
  {32'h4020c2f2, 32'h40c8c232} /* (28, 17, 27) {real, imag} */,
  {32'h3fa81de1, 32'h40c5c5c7} /* (28, 17, 26) {real, imag} */,
  {32'h402180fc, 32'h405b752a} /* (28, 17, 25) {real, imag} */,
  {32'h4077620a, 32'h402b90e1} /* (28, 17, 24) {real, imag} */,
  {32'h4098f478, 32'h404605bd} /* (28, 17, 23) {real, imag} */,
  {32'h40946642, 32'h40adb354} /* (28, 17, 22) {real, imag} */,
  {32'h40a1e6ac, 32'h3e38d06a} /* (28, 17, 21) {real, imag} */,
  {32'h3f8f7544, 32'hc0b04e16} /* (28, 17, 20) {real, imag} */,
  {32'hbf7718fc, 32'hc06cafb7} /* (28, 17, 19) {real, imag} */,
  {32'hc0189e97, 32'hbfaabdbe} /* (28, 17, 18) {real, imag} */,
  {32'hc024bf76, 32'hc0ad03fc} /* (28, 17, 17) {real, imag} */,
  {32'h3f127b28, 32'hc0b3a1a8} /* (28, 17, 16) {real, imag} */,
  {32'hbf2694f3, 32'hc08504ed} /* (28, 17, 15) {real, imag} */,
  {32'hc0866a12, 32'hc04010ff} /* (28, 17, 14) {real, imag} */,
  {32'hc06a99e2, 32'hc0556404} /* (28, 17, 13) {real, imag} */,
  {32'hc026733c, 32'hc086c80f} /* (28, 17, 12) {real, imag} */,
  {32'hbf5646bc, 32'hc000e5a0} /* (28, 17, 11) {real, imag} */,
  {32'h3f980bfa, 32'h40bb046c} /* (28, 17, 10) {real, imag} */,
  {32'h40224060, 32'h40dd5b91} /* (28, 17, 9) {real, imag} */,
  {32'h3fdcc6ad, 32'h40951a4a} /* (28, 17, 8) {real, imag} */,
  {32'h405c5578, 32'h40aca6ca} /* (28, 17, 7) {real, imag} */,
  {32'h4010473e, 32'h40cfb23c} /* (28, 17, 6) {real, imag} */,
  {32'hc0337f36, 32'h408358da} /* (28, 17, 5) {real, imag} */,
  {32'hbf984851, 32'h40863d52} /* (28, 17, 4) {real, imag} */,
  {32'h3e854cb2, 32'h3fd15608} /* (28, 17, 3) {real, imag} */,
  {32'hbffc3f47, 32'hbf0935f7} /* (28, 17, 2) {real, imag} */,
  {32'hc00a2801, 32'h3fd5516c} /* (28, 17, 1) {real, imag} */,
  {32'h3f0a5755, 32'h405d71fc} /* (28, 17, 0) {real, imag} */,
  {32'hbf101bea, 32'h40022428} /* (28, 16, 31) {real, imag} */,
  {32'h3da94208, 32'h40a01d1a} /* (28, 16, 30) {real, imag} */,
  {32'h40340356, 32'h40bb55f2} /* (28, 16, 29) {real, imag} */,
  {32'h4067fe3b, 32'h4059a41a} /* (28, 16, 28) {real, imag} */,
  {32'h3fdcb534, 32'h40a2431e} /* (28, 16, 27) {real, imag} */,
  {32'h3ede4ca4, 32'h408d8f76} /* (28, 16, 26) {real, imag} */,
  {32'h3f8ac3bd, 32'h4075dc87} /* (28, 16, 25) {real, imag} */,
  {32'h403ab86f, 32'h40bd5cd0} /* (28, 16, 24) {real, imag} */,
  {32'h4083f552, 32'h4082db37} /* (28, 16, 23) {real, imag} */,
  {32'h405ed41c, 32'h40c52915} /* (28, 16, 22) {real, imag} */,
  {32'h4004d860, 32'h4035a2c9} /* (28, 16, 21) {real, imag} */,
  {32'hbf6e7eac, 32'hc0ab0fd5} /* (28, 16, 20) {real, imag} */,
  {32'hbf659db8, 32'hc0c37966} /* (28, 16, 19) {real, imag} */,
  {32'h3f7a54ea, 32'hc05e4636} /* (28, 16, 18) {real, imag} */,
  {32'hbffd56bc, 32'hc0c7da92} /* (28, 16, 17) {real, imag} */,
  {32'hc013760e, 32'hc0c4291a} /* (28, 16, 16) {real, imag} */,
  {32'hbf3729b1, 32'hc0d7f1fa} /* (28, 16, 15) {real, imag} */,
  {32'hc03ecbd2, 32'hc09eacbe} /* (28, 16, 14) {real, imag} */,
  {32'hc0460af2, 32'hc08cd396} /* (28, 16, 13) {real, imag} */,
  {32'hc0941c2a, 32'hc093b986} /* (28, 16, 12) {real, imag} */,
  {32'hbfb900a4, 32'hc0212c86} /* (28, 16, 11) {real, imag} */,
  {32'h3f8947e2, 32'h40743fd6} /* (28, 16, 10) {real, imag} */,
  {32'h4023c67c, 32'h40a5627e} /* (28, 16, 9) {real, imag} */,
  {32'h3feae2b6, 32'h40a923f6} /* (28, 16, 8) {real, imag} */,
  {32'h4056827e, 32'h41099040} /* (28, 16, 7) {real, imag} */,
  {32'h4021b516, 32'h41103d3a} /* (28, 16, 6) {real, imag} */,
  {32'h3d373cbc, 32'h40a05c77} /* (28, 16, 5) {real, imag} */,
  {32'h3faea607, 32'h403f10f3} /* (28, 16, 4) {real, imag} */,
  {32'h3f575fb4, 32'h403c448d} /* (28, 16, 3) {real, imag} */,
  {32'hbf8a6e31, 32'h406c0fa4} /* (28, 16, 2) {real, imag} */,
  {32'h3f99f5d8, 32'h40b6aa04} /* (28, 16, 1) {real, imag} */,
  {32'h3fc841d0, 32'h40706166} /* (28, 16, 0) {real, imag} */,
  {32'hbf9f3f0b, 32'h3ff0f968} /* (28, 15, 31) {real, imag} */,
  {32'hbf84d7f7, 32'h40382a5d} /* (28, 15, 30) {real, imag} */,
  {32'h3f8709b8, 32'h408fd70c} /* (28, 15, 29) {real, imag} */,
  {32'h4016c760, 32'h40ae988c} /* (28, 15, 28) {real, imag} */,
  {32'h3fe16804, 32'h40a1dbe7} /* (28, 15, 27) {real, imag} */,
  {32'h3d88419c, 32'h4066415a} /* (28, 15, 26) {real, imag} */,
  {32'hbfd46514, 32'h405d0c36} /* (28, 15, 25) {real, imag} */,
  {32'hbf2d20ba, 32'h40972c15} /* (28, 15, 24) {real, imag} */,
  {32'h3f48a65f, 32'h40aee574} /* (28, 15, 23) {real, imag} */,
  {32'h3f010900, 32'h40d570e2} /* (28, 15, 22) {real, imag} */,
  {32'hbedd8aeb, 32'h40a7c5ed} /* (28, 15, 21) {real, imag} */,
  {32'hbfa4a130, 32'hbfbcebce} /* (28, 15, 20) {real, imag} */,
  {32'hbf9eb5ab, 32'hc0d12f7a} /* (28, 15, 19) {real, imag} */,
  {32'h3f32437a, 32'hc0a5d2a0} /* (28, 15, 18) {real, imag} */,
  {32'hbefdac28, 32'hc0bf4332} /* (28, 15, 17) {real, imag} */,
  {32'hbfe89059, 32'hc0d92264} /* (28, 15, 16) {real, imag} */,
  {32'hbf3d4459, 32'hc0ceb5dc} /* (28, 15, 15) {real, imag} */,
  {32'hbf739b16, 32'hc0e84ad4} /* (28, 15, 14) {real, imag} */,
  {32'h3f2448c3, 32'hc094ce2a} /* (28, 15, 13) {real, imag} */,
  {32'hbfe48c60, 32'hc03a167a} /* (28, 15, 12) {real, imag} */,
  {32'hbf0ae2b8, 32'hc017fafa} /* (28, 15, 11) {real, imag} */,
  {32'h3fdd1d46, 32'h404f35dc} /* (28, 15, 10) {real, imag} */,
  {32'h40032ec6, 32'h409b6288} /* (28, 15, 9) {real, imag} */,
  {32'h3fd9eacc, 32'h409ba0e2} /* (28, 15, 8) {real, imag} */,
  {32'h4039b959, 32'h40fbd5ef} /* (28, 15, 7) {real, imag} */,
  {32'h406e9acc, 32'h40d4e2f2} /* (28, 15, 6) {real, imag} */,
  {32'h4004932e, 32'h408bbaeb} /* (28, 15, 5) {real, imag} */,
  {32'h4013a4f3, 32'h400b2602} /* (28, 15, 4) {real, imag} */,
  {32'h3fe3d24c, 32'h4058c6b5} /* (28, 15, 3) {real, imag} */,
  {32'h3f9dfc81, 32'h40c99c92} /* (28, 15, 2) {real, imag} */,
  {32'h3fce52cf, 32'h40d4468d} /* (28, 15, 1) {real, imag} */,
  {32'h3feac00c, 32'h40551500} /* (28, 15, 0) {real, imag} */,
  {32'h3f18cd8b, 32'h3ff14911} /* (28, 14, 31) {real, imag} */,
  {32'h3fd611f8, 32'h401ac97c} /* (28, 14, 30) {real, imag} */,
  {32'h3fd4676e, 32'h40b52a2e} /* (28, 14, 29) {real, imag} */,
  {32'hbf8c15f8, 32'h40d185f8} /* (28, 14, 28) {real, imag} */,
  {32'hbe8d56f2, 32'h4091e0e5} /* (28, 14, 27) {real, imag} */,
  {32'hbe3cd9e4, 32'h4031ff92} /* (28, 14, 26) {real, imag} */,
  {32'hbfb0a2ae, 32'h4020f3b6} /* (28, 14, 25) {real, imag} */,
  {32'h4028858d, 32'h40606eae} /* (28, 14, 24) {real, imag} */,
  {32'h408480bf, 32'h408cbb6e} /* (28, 14, 23) {real, imag} */,
  {32'h3f1b1f58, 32'h40c15e56} /* (28, 14, 22) {real, imag} */,
  {32'hbff27688, 32'h406039b2} /* (28, 14, 21) {real, imag} */,
  {32'hbea45f68, 32'hc03d8e24} /* (28, 14, 20) {real, imag} */,
  {32'hc08224f8, 32'hc0b29e1c} /* (28, 14, 19) {real, imag} */,
  {32'hc04c5584, 32'hc094774e} /* (28, 14, 18) {real, imag} */,
  {32'hbf2bb8b0, 32'hc099c866} /* (28, 14, 17) {real, imag} */,
  {32'hbfa55495, 32'hc0fd4fa7} /* (28, 14, 16) {real, imag} */,
  {32'hbf3795ec, 32'hc0d72160} /* (28, 14, 15) {real, imag} */,
  {32'hc02e12c6, 32'hc0ef9bad} /* (28, 14, 14) {real, imag} */,
  {32'hbfa73d30, 32'hc0a334ae} /* (28, 14, 13) {real, imag} */,
  {32'hc01a8eac, 32'hbfdbb394} /* (28, 14, 12) {real, imag} */,
  {32'hbfa04b10, 32'hbf9acbc0} /* (28, 14, 11) {real, imag} */,
  {32'h3fc63c73, 32'h40913361} /* (28, 14, 10) {real, imag} */,
  {32'h3ec4d3ea, 32'h40b00efe} /* (28, 14, 9) {real, imag} */,
  {32'hbe0a9ac4, 32'h4081a47f} /* (28, 14, 8) {real, imag} */,
  {32'h3fc53bd4, 32'h409a530e} /* (28, 14, 7) {real, imag} */,
  {32'h3fc3a150, 32'h40acac57} /* (28, 14, 6) {real, imag} */,
  {32'h3fb86d70, 32'h40944764} /* (28, 14, 5) {real, imag} */,
  {32'h4065beef, 32'h406f9877} /* (28, 14, 4) {real, imag} */,
  {32'h409f44c4, 32'h40d637c6} /* (28, 14, 3) {real, imag} */,
  {32'h403bffea, 32'h40f42494} /* (28, 14, 2) {real, imag} */,
  {32'h3f944ca2, 32'h406f3bfc} /* (28, 14, 1) {real, imag} */,
  {32'h3fd2909a, 32'h3f34bd1e} /* (28, 14, 0) {real, imag} */,
  {32'h4016d642, 32'h3fef3c45} /* (28, 13, 31) {real, imag} */,
  {32'h40719df4, 32'h40b777d6} /* (28, 13, 30) {real, imag} */,
  {32'h405b031e, 32'h40dba3dc} /* (28, 13, 29) {real, imag} */,
  {32'h3ff2a66a, 32'h40e11c2b} /* (28, 13, 28) {real, imag} */,
  {32'h3ecf4a78, 32'h40a8dcca} /* (28, 13, 27) {real, imag} */,
  {32'hbe50d8b8, 32'h4064030b} /* (28, 13, 26) {real, imag} */,
  {32'h404edbb2, 32'h40ae1bde} /* (28, 13, 25) {real, imag} */,
  {32'h4083c9c6, 32'h40f2e9a4} /* (28, 13, 24) {real, imag} */,
  {32'h4017007a, 32'h409ee4ac} /* (28, 13, 23) {real, imag} */,
  {32'hbf9788c2, 32'h4073e05b} /* (28, 13, 22) {real, imag} */,
  {32'hbfd73af2, 32'h4023f1b9} /* (28, 13, 21) {real, imag} */,
  {32'h3f386c74, 32'hc047b682} /* (28, 13, 20) {real, imag} */,
  {32'hc039c226, 32'hc07be793} /* (28, 13, 19) {real, imag} */,
  {32'hc09fde33, 32'hbf8d8c0b} /* (28, 13, 18) {real, imag} */,
  {32'hc01a81aa, 32'hc09e8817} /* (28, 13, 17) {real, imag} */,
  {32'hbffaa4a5, 32'hc1062e90} /* (28, 13, 16) {real, imag} */,
  {32'hbfafc154, 32'hc100dc1f} /* (28, 13, 15) {real, imag} */,
  {32'hbf2a9c16, 32'hc0f8ce13} /* (28, 13, 14) {real, imag} */,
  {32'h3f603c69, 32'hc0919955} /* (28, 13, 13) {real, imag} */,
  {32'hbfdd997c, 32'hc02c5656} /* (28, 13, 12) {real, imag} */,
  {32'hc00aec5c, 32'hbf319418} /* (28, 13, 11) {real, imag} */,
  {32'h3fec85a8, 32'h40886c58} /* (28, 13, 10) {real, imag} */,
  {32'h3fdcc792, 32'h40aaafd8} /* (28, 13, 9) {real, imag} */,
  {32'h3ff65524, 32'h40a27734} /* (28, 13, 8) {real, imag} */,
  {32'h40577191, 32'h409ea676} /* (28, 13, 7) {real, imag} */,
  {32'h3f9aa62a, 32'h40a0f17c} /* (28, 13, 6) {real, imag} */,
  {32'h3f5317ca, 32'h40af46eb} /* (28, 13, 5) {real, imag} */,
  {32'h404f824e, 32'h40b0957e} /* (28, 13, 4) {real, imag} */,
  {32'h40a6c779, 32'h40ff7f2a} /* (28, 13, 3) {real, imag} */,
  {32'h4020d361, 32'h40d1b175} /* (28, 13, 2) {real, imag} */,
  {32'hbd35bcd0, 32'h4051011c} /* (28, 13, 1) {real, imag} */,
  {32'hbe89e5fe, 32'h3fc78322} /* (28, 13, 0) {real, imag} */,
  {32'h40778010, 32'h3fdf719d} /* (28, 12, 31) {real, imag} */,
  {32'h408e5bb6, 32'h40bc539a} /* (28, 12, 30) {real, imag} */,
  {32'h403bd002, 32'h40e3bf1b} /* (28, 12, 29) {real, imag} */,
  {32'h4056f851, 32'h40ccef86} /* (28, 12, 28) {real, imag} */,
  {32'h400893b8, 32'h40baff12} /* (28, 12, 27) {real, imag} */,
  {32'h4021622d, 32'h40a3d2f0} /* (28, 12, 26) {real, imag} */,
  {32'h406e88b3, 32'h40e89c98} /* (28, 12, 25) {real, imag} */,
  {32'h4085a2f8, 32'h40f8ad7f} /* (28, 12, 24) {real, imag} */,
  {32'h4010eb3f, 32'h40a454b1} /* (28, 12, 23) {real, imag} */,
  {32'h3f0ed524, 32'h4080be71} /* (28, 12, 22) {real, imag} */,
  {32'h3fb563ed, 32'h4052c9c9} /* (28, 12, 21) {real, imag} */,
  {32'hbf010075, 32'hc054ba3c} /* (28, 12, 20) {real, imag} */,
  {32'hc0bf76db, 32'hc0aeff4e} /* (28, 12, 19) {real, imag} */,
  {32'hc0f55e8d, 32'hc0333e07} /* (28, 12, 18) {real, imag} */,
  {32'hc095bb62, 32'hc0b1656c} /* (28, 12, 17) {real, imag} */,
  {32'hc0860537, 32'hc0e55258} /* (28, 12, 16) {real, imag} */,
  {32'hc015f434, 32'hc0d854c0} /* (28, 12, 15) {real, imag} */,
  {32'h3f5c4630, 32'hc0abe1b4} /* (28, 12, 14) {real, imag} */,
  {32'h3fbd3641, 32'hc0ad4589} /* (28, 12, 13) {real, imag} */,
  {32'hbfdefc0f, 32'hc104e4c2} /* (28, 12, 12) {real, imag} */,
  {32'hc06a044c, 32'hc0c1be48} /* (28, 12, 11) {real, imag} */,
  {32'h3e839cf3, 32'h3e8fc052} /* (28, 12, 10) {real, imag} */,
  {32'h3fa470b2, 32'h40881fda} /* (28, 12, 9) {real, imag} */,
  {32'h40050388, 32'h40b6beb6} /* (28, 12, 8) {real, imag} */,
  {32'h404b334e, 32'h40aa04d5} /* (28, 12, 7) {real, imag} */,
  {32'h408f687c, 32'h40a2f794} /* (28, 12, 6) {real, imag} */,
  {32'h40912b0e, 32'h4067530e} /* (28, 12, 5) {real, imag} */,
  {32'h400bae76, 32'h4053c7a0} /* (28, 12, 4) {real, imag} */,
  {32'h407e6900, 32'h40c8ce92} /* (28, 12, 3) {real, imag} */,
  {32'h40b5f4c0, 32'h40be396a} /* (28, 12, 2) {real, imag} */,
  {32'h408c5f0c, 32'h40c05424} /* (28, 12, 1) {real, imag} */,
  {32'h3feeb9ec, 32'h408571ff} /* (28, 12, 0) {real, imag} */,
  {32'h401a521e, 32'h3f67dde6} /* (28, 11, 31) {real, imag} */,
  {32'h3ff04cfe, 32'h40736f2e} /* (28, 11, 30) {real, imag} */,
  {32'h3f148a53, 32'h40c74b76} /* (28, 11, 29) {real, imag} */,
  {32'h3f81bfb6, 32'h40923f32} /* (28, 11, 28) {real, imag} */,
  {32'h3efbb496, 32'h40567b8a} /* (28, 11, 27) {real, imag} */,
  {32'h3fec483d, 32'h402430fe} /* (28, 11, 26) {real, imag} */,
  {32'h3fdcf1ff, 32'h406934c8} /* (28, 11, 25) {real, imag} */,
  {32'h407612c1, 32'h403bbe8e} /* (28, 11, 24) {real, imag} */,
  {32'h402a2504, 32'h4099a0c0} /* (28, 11, 23) {real, imag} */,
  {32'h3f83c14b, 32'h40839d42} /* (28, 11, 22) {real, imag} */,
  {32'h401fdf5e, 32'h40a073b9} /* (28, 11, 21) {real, imag} */,
  {32'h3eeb1def, 32'hbf353671} /* (28, 11, 20) {real, imag} */,
  {32'hc01c48b0, 32'hc0820673} /* (28, 11, 19) {real, imag} */,
  {32'hc0637e7a, 32'hc09b8a28} /* (28, 11, 18) {real, imag} */,
  {32'hc08853f8, 32'hc0caf940} /* (28, 11, 17) {real, imag} */,
  {32'hc07274f0, 32'hc09885b6} /* (28, 11, 16) {real, imag} */,
  {32'hc017aa97, 32'hc026fa15} /* (28, 11, 15) {real, imag} */,
  {32'hbecc037e, 32'hc09cffcc} /* (28, 11, 14) {real, imag} */,
  {32'hbf133b60, 32'hc094955f} /* (28, 11, 13) {real, imag} */,
  {32'hbfa8c687, 32'hc09c878e} /* (28, 11, 12) {real, imag} */,
  {32'hc007f51f, 32'hc0a7f78a} /* (28, 11, 11) {real, imag} */,
  {32'hc03abdc8, 32'h3fc482d9} /* (28, 11, 10) {real, imag} */,
  {32'h3fc2fc36, 32'h40ec2e51} /* (28, 11, 9) {real, imag} */,
  {32'h40662ca4, 32'h40babfd8} /* (28, 11, 8) {real, imag} */,
  {32'h409a633d, 32'h40b039ac} /* (28, 11, 7) {real, imag} */,
  {32'h40c36b7e, 32'h40de74fe} /* (28, 11, 6) {real, imag} */,
  {32'h40808802, 32'h40c13ad0} /* (28, 11, 5) {real, imag} */,
  {32'h402cf1a6, 32'h40729936} /* (28, 11, 4) {real, imag} */,
  {32'h4045b3fa, 32'h406a92d1} /* (28, 11, 3) {real, imag} */,
  {32'h404af6e1, 32'h404cf7ae} /* (28, 11, 2) {real, imag} */,
  {32'h3f59df00, 32'h4081e1bb} /* (28, 11, 1) {real, imag} */,
  {32'h3fd0cca4, 32'h404b0e41} /* (28, 11, 0) {real, imag} */,
  {32'hbfd253cc, 32'hc06992a8} /* (28, 10, 31) {real, imag} */,
  {32'hc04026b5, 32'hc045ec32} /* (28, 10, 30) {real, imag} */,
  {32'hbfe14e06, 32'hbff80f44} /* (28, 10, 29) {real, imag} */,
  {32'hbfb4734c, 32'hc074382c} /* (28, 10, 28) {real, imag} */,
  {32'hc02759be, 32'hc07a4fd4} /* (28, 10, 27) {real, imag} */,
  {32'hbf9d2de9, 32'hc0955d22} /* (28, 10, 26) {real, imag} */,
  {32'hbf7904e5, 32'hc08691b8} /* (28, 10, 25) {real, imag} */,
  {32'hbe2c4758, 32'hc0770484} /* (28, 10, 24) {real, imag} */,
  {32'h3d90c036, 32'hbea3a29c} /* (28, 10, 23) {real, imag} */,
  {32'hbf19fdb9, 32'hbf1d72f6} /* (28, 10, 22) {real, imag} */,
  {32'h3ee3877b, 32'h4069a158} /* (28, 10, 21) {real, imag} */,
  {32'h403d49c2, 32'h408a062a} /* (28, 10, 20) {real, imag} */,
  {32'h3fb0712a, 32'h3f0598b2} /* (28, 10, 19) {real, imag} */,
  {32'h400b8880, 32'h3e082ea0} /* (28, 10, 18) {real, imag} */,
  {32'h401893b4, 32'h3fab98a1} /* (28, 10, 17) {real, imag} */,
  {32'hbf988c53, 32'h401d228d} /* (28, 10, 16) {real, imag} */,
  {32'hbff8a099, 32'h40941a4e} /* (28, 10, 15) {real, imag} */,
  {32'hbe2e9128, 32'h3ff0b422} /* (28, 10, 14) {real, imag} */,
  {32'h3f5cb248, 32'h401483c2} /* (28, 10, 13) {real, imag} */,
  {32'h3fa8b28d, 32'h4020caeb} /* (28, 10, 12) {real, imag} */,
  {32'h3ef2911e, 32'h3fc0ba04} /* (28, 10, 11) {real, imag} */,
  {32'hbf5ab3e8, 32'h3f3662bb} /* (28, 10, 10) {real, imag} */,
  {32'h3fa55964, 32'h3e3d2630} /* (28, 10, 9) {real, imag} */,
  {32'h3f8725a7, 32'hc025d318} /* (28, 10, 8) {real, imag} */,
  {32'h3e439e80, 32'hbf0c95db} /* (28, 10, 7) {real, imag} */,
  {32'h3fcde138, 32'h40009fea} /* (28, 10, 6) {real, imag} */,
  {32'h3ec1486e, 32'hbe5b1e45} /* (28, 10, 5) {real, imag} */,
  {32'hbda8b564, 32'hbf73a9bd} /* (28, 10, 4) {real, imag} */,
  {32'h3ea090f6, 32'hc05a4f4d} /* (28, 10, 3) {real, imag} */,
  {32'h3e132a39, 32'hc0ba6621} /* (28, 10, 2) {real, imag} */,
  {32'hc05b5ac2, 32'hc0a87b95} /* (28, 10, 1) {real, imag} */,
  {32'hbf95c5ec, 32'hc065f720} /* (28, 10, 0) {real, imag} */,
  {32'hc01f841f, 32'hc080deb8} /* (28, 9, 31) {real, imag} */,
  {32'hc04ebc12, 32'hc0c3880a} /* (28, 9, 30) {real, imag} */,
  {32'hc02a7d45, 32'hc0098cb3} /* (28, 9, 29) {real, imag} */,
  {32'hc01f90c4, 32'hc08f29c2} /* (28, 9, 28) {real, imag} */,
  {32'hc076f58c, 32'hc0c5ebe3} /* (28, 9, 27) {real, imag} */,
  {32'hc02d0d02, 32'hc0f6e8fe} /* (28, 9, 26) {real, imag} */,
  {32'hc014d262, 32'hc0dbc6d2} /* (28, 9, 25) {real, imag} */,
  {32'hc03b90bc, 32'hc0b5f12e} /* (28, 9, 24) {real, imag} */,
  {32'hbfae09ab, 32'hc083a901} /* (28, 9, 23) {real, imag} */,
  {32'hbff19077, 32'hc0d84cc0} /* (28, 9, 22) {real, imag} */,
  {32'hbf28c779, 32'hc0221f25} /* (28, 9, 21) {real, imag} */,
  {32'h3fb8f130, 32'h4095211b} /* (28, 9, 20) {real, imag} */,
  {32'h3ff5bcd3, 32'h406a4895} /* (28, 9, 19) {real, imag} */,
  {32'h3f00cfe6, 32'h40710180} /* (28, 9, 18) {real, imag} */,
  {32'h401ec09f, 32'h40bd3bdd} /* (28, 9, 17) {real, imag} */,
  {32'h4029a758, 32'h40939c66} /* (28, 9, 16) {real, imag} */,
  {32'h3e82f99e, 32'h40c5868e} /* (28, 9, 15) {real, imag} */,
  {32'h401e9476, 32'h40cfcd12} /* (28, 9, 14) {real, imag} */,
  {32'h3f828f39, 32'h40378679} /* (28, 9, 13) {real, imag} */,
  {32'h3fd47c1e, 32'h4088db5c} /* (28, 9, 12) {real, imag} */,
  {32'h3f95e725, 32'h4080c478} /* (28, 9, 11) {real, imag} */,
  {32'hc023cf39, 32'hbf75e2aa} /* (28, 9, 10) {real, imag} */,
  {32'hbf954d6d, 32'hc03cc59d} /* (28, 9, 9) {real, imag} */,
  {32'hbfa38906, 32'hc049caeb} /* (28, 9, 8) {real, imag} */,
  {32'hc0218fa6, 32'hc05f1c5c} /* (28, 9, 7) {real, imag} */,
  {32'h3f524a0b, 32'hbffad769} /* (28, 9, 6) {real, imag} */,
  {32'hbfc2095c, 32'hc0ce8d55} /* (28, 9, 5) {real, imag} */,
  {32'hbee025fc, 32'hc0d4fb5c} /* (28, 9, 4) {real, imag} */,
  {32'hbf936917, 32'hc0d6a489} /* (28, 9, 3) {real, imag} */,
  {32'hbf846d03, 32'hc1058f28} /* (28, 9, 2) {real, imag} */,
  {32'hc018e616, 32'hc10219df} /* (28, 9, 1) {real, imag} */,
  {32'hbfce068f, 32'hc0aa5884} /* (28, 9, 0) {real, imag} */,
  {32'hbfc050c5, 32'hc093f578} /* (28, 8, 31) {real, imag} */,
  {32'hbefac69c, 32'hc0d503da} /* (28, 8, 30) {real, imag} */,
  {32'hbf2b1128, 32'hc03cad75} /* (28, 8, 29) {real, imag} */,
  {32'hbeebb18e, 32'hc057cc29} /* (28, 8, 28) {real, imag} */,
  {32'hbf5f271f, 32'hc0387652} /* (28, 8, 27) {real, imag} */,
  {32'hbf0897c2, 32'hc09369aa} /* (28, 8, 26) {real, imag} */,
  {32'hbf5603fe, 32'hc062e252} /* (28, 8, 25) {real, imag} */,
  {32'hc02c75e6, 32'hc0757320} /* (28, 8, 24) {real, imag} */,
  {32'hc0099894, 32'hc075a6d7} /* (28, 8, 23) {real, imag} */,
  {32'hbf9acfa2, 32'hc09db6fa} /* (28, 8, 22) {real, imag} */,
  {32'hbf933457, 32'hc009fb9b} /* (28, 8, 21) {real, imag} */,
  {32'hbf9f3d6e, 32'h408b1fc2} /* (28, 8, 20) {real, imag} */,
  {32'hbd0f901a, 32'h40a84f4c} /* (28, 8, 19) {real, imag} */,
  {32'hbf6a76d7, 32'h4046af56} /* (28, 8, 18) {real, imag} */,
  {32'h3f890413, 32'h403e98d8} /* (28, 8, 17) {real, imag} */,
  {32'h40931506, 32'h40891a27} /* (28, 8, 16) {real, imag} */,
  {32'h3f99eb77, 32'h40750af2} /* (28, 8, 15) {real, imag} */,
  {32'h4036d118, 32'h40c9129a} /* (28, 8, 14) {real, imag} */,
  {32'h405a77e2, 32'h4092548b} /* (28, 8, 13) {real, imag} */,
  {32'h4025f046, 32'h40949d3c} /* (28, 8, 12) {real, imag} */,
  {32'h3fb0d1a9, 32'h3fee243a} /* (28, 8, 11) {real, imag} */,
  {32'h3c366ac0, 32'hc08b06d5} /* (28, 8, 10) {real, imag} */,
  {32'h3d8397f4, 32'hc084a422} /* (28, 8, 9) {real, imag} */,
  {32'hbf7a1625, 32'hbffc3934} /* (28, 8, 8) {real, imag} */,
  {32'hc01beeeb, 32'hc033599e} /* (28, 8, 7) {real, imag} */,
  {32'h3f15e495, 32'hc056fb1e} /* (28, 8, 6) {real, imag} */,
  {32'hc016f64a, 32'hc09a4960} /* (28, 8, 5) {real, imag} */,
  {32'hbeed48ca, 32'hc09ac014} /* (28, 8, 4) {real, imag} */,
  {32'hbe73f4d4, 32'hc0ea9d78} /* (28, 8, 3) {real, imag} */,
  {32'hc07f31c2, 32'hc0f148be} /* (28, 8, 2) {real, imag} */,
  {32'hc08467eb, 32'hc0d35e12} /* (28, 8, 1) {real, imag} */,
  {32'hbffb33aa, 32'hc0aff3f1} /* (28, 8, 0) {real, imag} */,
  {32'hbf4ae59c, 32'hc094e537} /* (28, 7, 31) {real, imag} */,
  {32'hbf46e7d8, 32'hc0c72c3f} /* (28, 7, 30) {real, imag} */,
  {32'h3ff9704c, 32'hc09d198c} /* (28, 7, 29) {real, imag} */,
  {32'hbd191c60, 32'hc0a002bb} /* (28, 7, 28) {real, imag} */,
  {32'hbfcb51f0, 32'hc04040dd} /* (28, 7, 27) {real, imag} */,
  {32'hbfdb155d, 32'hc080a250} /* (28, 7, 26) {real, imag} */,
  {32'hc00384eb, 32'hc06d93c4} /* (28, 7, 25) {real, imag} */,
  {32'hbfb374b9, 32'hc0b98f68} /* (28, 7, 24) {real, imag} */,
  {32'hc06e0fc4, 32'hc0965484} /* (28, 7, 23) {real, imag} */,
  {32'hbfe98c6c, 32'hc0a130b3} /* (28, 7, 22) {real, imag} */,
  {32'hbf36e7c8, 32'hbfcfad43} /* (28, 7, 21) {real, imag} */,
  {32'h3f9287e6, 32'h40d785f3} /* (28, 7, 20) {real, imag} */,
  {32'h3f6ffb62, 32'h40ac7c92} /* (28, 7, 19) {real, imag} */,
  {32'hbe8ebc52, 32'h4082749b} /* (28, 7, 18) {real, imag} */,
  {32'h3e1ea2f6, 32'h40815a46} /* (28, 7, 17) {real, imag} */,
  {32'h3db56784, 32'h4067816c} /* (28, 7, 16) {real, imag} */,
  {32'hbf73e91e, 32'h40b4050b} /* (28, 7, 15) {real, imag} */,
  {32'h3fd0e542, 32'h40e0a67c} /* (28, 7, 14) {real, imag} */,
  {32'h405c7f26, 32'h409a5a86} /* (28, 7, 13) {real, imag} */,
  {32'h3fb56270, 32'h40940c91} /* (28, 7, 12) {real, imag} */,
  {32'h3f081141, 32'h3ff8ffa7} /* (28, 7, 11) {real, imag} */,
  {32'h3f0c664d, 32'hc0b17481} /* (28, 7, 10) {real, imag} */,
  {32'hbfe2cd8e, 32'hc0d3416b} /* (28, 7, 9) {real, imag} */,
  {32'hbfb3e6cc, 32'hc0b3a5f5} /* (28, 7, 8) {real, imag} */,
  {32'hbf92179c, 32'hc08df42a} /* (28, 7, 7) {real, imag} */,
  {32'hbfe9332b, 32'hc07e273a} /* (28, 7, 6) {real, imag} */,
  {32'hc01fc5a6, 32'hc09f9fd6} /* (28, 7, 5) {real, imag} */,
  {32'hc02ae63a, 32'hc09bc6ec} /* (28, 7, 4) {real, imag} */,
  {32'hbfc4d5c6, 32'hc0bc0c6a} /* (28, 7, 3) {real, imag} */,
  {32'hc0c2a92a, 32'hc0e2916a} /* (28, 7, 2) {real, imag} */,
  {32'hc08f1fb6, 32'hc0b807f0} /* (28, 7, 1) {real, imag} */,
  {32'h3d81c520, 32'hc041c7f0} /* (28, 7, 0) {real, imag} */,
  {32'hbf2f1181, 32'hc03ece16} /* (28, 6, 31) {real, imag} */,
  {32'hbfb6f213, 32'hc0e8d8c8} /* (28, 6, 30) {real, imag} */,
  {32'hbe5ceb64, 32'hc0be8afd} /* (28, 6, 29) {real, imag} */,
  {32'hbfd3d302, 32'hc04c4732} /* (28, 6, 28) {real, imag} */,
  {32'hc00bfd08, 32'hc0218c98} /* (28, 6, 27) {real, imag} */,
  {32'hc06d842a, 32'hc0634524} /* (28, 6, 26) {real, imag} */,
  {32'hc08b096c, 32'hc0b890f4} /* (28, 6, 25) {real, imag} */,
  {32'hbfde7c87, 32'hc0e434a0} /* (28, 6, 24) {real, imag} */,
  {32'hc0538da0, 32'hc085250b} /* (28, 6, 23) {real, imag} */,
  {32'hc0881583, 32'hc0a0349a} /* (28, 6, 22) {real, imag} */,
  {32'hc088575f, 32'hc01829b4} /* (28, 6, 21) {real, imag} */,
  {32'h400108b4, 32'h40cd7fe8} /* (28, 6, 20) {real, imag} */,
  {32'h3fc036b5, 32'h409cf15e} /* (28, 6, 19) {real, imag} */,
  {32'h3ffcea60, 32'h4046759a} /* (28, 6, 18) {real, imag} */,
  {32'h3f6db947, 32'h40c2b57c} /* (28, 6, 17) {real, imag} */,
  {32'h3f802ece, 32'h40845a54} /* (28, 6, 16) {real, imag} */,
  {32'h3d8317d4, 32'h4098047e} /* (28, 6, 15) {real, imag} */,
  {32'h3f238b2c, 32'h409784eb} /* (28, 6, 14) {real, imag} */,
  {32'h4015b0b0, 32'h3fe5e003} /* (28, 6, 13) {real, imag} */,
  {32'h3ff6f9d6, 32'h40a64b95} /* (28, 6, 12) {real, imag} */,
  {32'h3fe5194b, 32'h4077e18f} /* (28, 6, 11) {real, imag} */,
  {32'hbf304632, 32'hbfc073e8} /* (28, 6, 10) {real, imag} */,
  {32'hc0934811, 32'hc0a9f355} /* (28, 6, 9) {real, imag} */,
  {32'hc03c965b, 32'hc09b61de} /* (28, 6, 8) {real, imag} */,
  {32'hc0391d0d, 32'hc05b098d} /* (28, 6, 7) {real, imag} */,
  {32'hbf472c43, 32'hc0a718d2} /* (28, 6, 6) {real, imag} */,
  {32'hbf21b40f, 32'hc0d09c47} /* (28, 6, 5) {real, imag} */,
  {32'hc059ba83, 32'hc0db4b56} /* (28, 6, 4) {real, imag} */,
  {32'hbfe31331, 32'hc0ab9bf2} /* (28, 6, 3) {real, imag} */,
  {32'hbfdd3520, 32'hc0dec746} /* (28, 6, 2) {real, imag} */,
  {32'hc012af6c, 32'hc0999654} /* (28, 6, 1) {real, imag} */,
  {32'hbf311dbc, 32'hbf1e1072} /* (28, 6, 0) {real, imag} */,
  {32'hbfee2cb9, 32'hc0ac44b8} /* (28, 5, 31) {real, imag} */,
  {32'hc093431a, 32'hc0c3729c} /* (28, 5, 30) {real, imag} */,
  {32'hc06f1dfc, 32'hc0b988e0} /* (28, 5, 29) {real, imag} */,
  {32'hc02d6b6f, 32'hc0a7d448} /* (28, 5, 28) {real, imag} */,
  {32'hbfe6404c, 32'hc0155981} /* (28, 5, 27) {real, imag} */,
  {32'hbfcea652, 32'hbfb8affa} /* (28, 5, 26) {real, imag} */,
  {32'hc0093ded, 32'hc062bb9e} /* (28, 5, 25) {real, imag} */,
  {32'hbe4d4134, 32'hc0c8a45e} /* (28, 5, 24) {real, imag} */,
  {32'hc0189aaf, 32'hc0a11d3f} /* (28, 5, 23) {real, imag} */,
  {32'hc07e2ed7, 32'hc0983ddc} /* (28, 5, 22) {real, imag} */,
  {32'hc0c693ec, 32'hc0132f6f} /* (28, 5, 21) {real, imag} */,
  {32'hbfb5f994, 32'h3f8ccbc9} /* (28, 5, 20) {real, imag} */,
  {32'hbf511a96, 32'h3e8a4b47} /* (28, 5, 19) {real, imag} */,
  {32'hc0085c8c, 32'hbf953a78} /* (28, 5, 18) {real, imag} */,
  {32'hc017029c, 32'h3f93e58f} /* (28, 5, 17) {real, imag} */,
  {32'hbfa76626, 32'h3e4a7d5b} /* (28, 5, 16) {real, imag} */,
  {32'h3e88a274, 32'h40340a48} /* (28, 5, 15) {real, imag} */,
  {32'h3ece4391, 32'h40248f94} /* (28, 5, 14) {real, imag} */,
  {32'h3f4ba5ea, 32'h4040d5ea} /* (28, 5, 13) {real, imag} */,
  {32'hbf48846b, 32'h40b86a6e} /* (28, 5, 12) {real, imag} */,
  {32'h3fcbd78d, 32'h40a5689c} /* (28, 5, 11) {real, imag} */,
  {32'hbe8bceb8, 32'h40973b0e} /* (28, 5, 10) {real, imag} */,
  {32'hbe8ee5c5, 32'h40545a52} /* (28, 5, 9) {real, imag} */,
  {32'hbefbe734, 32'h40457438} /* (28, 5, 8) {real, imag} */,
  {32'hbf98ba52, 32'h3fdfa18e} /* (28, 5, 7) {real, imag} */,
  {32'hbce5cd20, 32'hc011c794} /* (28, 5, 6) {real, imag} */,
  {32'hbf6870a7, 32'hc097d7fa} /* (28, 5, 5) {real, imag} */,
  {32'hbfcb260f, 32'hc10affe6} /* (28, 5, 4) {real, imag} */,
  {32'hc055e617, 32'hc0946546} /* (28, 5, 3) {real, imag} */,
  {32'hc0574e8c, 32'hc0935e27} /* (28, 5, 2) {real, imag} */,
  {32'hbfe896b8, 32'hc0786222} /* (28, 5, 1) {real, imag} */,
  {32'hbf75e182, 32'hbfb3a299} /* (28, 5, 0) {real, imag} */,
  {32'hbf8575bd, 32'hc090793c} /* (28, 4, 31) {real, imag} */,
  {32'hc08e548e, 32'hc0ac5ad0} /* (28, 4, 30) {real, imag} */,
  {32'hc085cdd2, 32'hc0afae46} /* (28, 4, 29) {real, imag} */,
  {32'hbf9d1158, 32'hc0a47174} /* (28, 4, 28) {real, imag} */,
  {32'h3f1acf57, 32'hc0906be8} /* (28, 4, 27) {real, imag} */,
  {32'h3f429b82, 32'hc04724bc} /* (28, 4, 26) {real, imag} */,
  {32'hbf5fcdd4, 32'hc00877f3} /* (28, 4, 25) {real, imag} */,
  {32'h3f98c703, 32'hc085f451} /* (28, 4, 24) {real, imag} */,
  {32'hbf6d1495, 32'hc0be2ca0} /* (28, 4, 23) {real, imag} */,
  {32'hc02ff7e0, 32'hc0ac022a} /* (28, 4, 22) {real, imag} */,
  {32'hc08f6ac5, 32'hc0b1144c} /* (28, 4, 21) {real, imag} */,
  {32'hc0b89366, 32'hc0a29934} /* (28, 4, 20) {real, imag} */,
  {32'hc033b29c, 32'hc085235f} /* (28, 4, 19) {real, imag} */,
  {32'hc05dec88, 32'hc0a1fbca} /* (28, 4, 18) {real, imag} */,
  {32'hc0be9192, 32'hc099f629} /* (28, 4, 17) {real, imag} */,
  {32'hc0a83a98, 32'hc00a9385} /* (28, 4, 16) {real, imag} */,
  {32'h3ec0b611, 32'h409c2768} /* (28, 4, 15) {real, imag} */,
  {32'h3ff7004b, 32'h40a07a92} /* (28, 4, 14) {real, imag} */,
  {32'h3e1d5a7e, 32'h4061803f} /* (28, 4, 13) {real, imag} */,
  {32'hbfccd680, 32'h409db210} /* (28, 4, 12) {real, imag} */,
  {32'h3e9c54ce, 32'h40db5718} /* (28, 4, 11) {real, imag} */,
  {32'h400450cc, 32'h41004f7c} /* (28, 4, 10) {real, imag} */,
  {32'h403bfe3c, 32'h40f0a5f1} /* (28, 4, 9) {real, imag} */,
  {32'h402bf483, 32'h40e6fefa} /* (28, 4, 8) {real, imag} */,
  {32'h4000bc2e, 32'h40b2ab3c} /* (28, 4, 7) {real, imag} */,
  {32'h3f57a28e, 32'h403a296a} /* (28, 4, 6) {real, imag} */,
  {32'hbfe992d2, 32'h3e230d44} /* (28, 4, 5) {real, imag} */,
  {32'hc0679d2e, 32'hc09bb19e} /* (28, 4, 4) {real, imag} */,
  {32'hbfbf6c12, 32'hc072e4c2} /* (28, 4, 3) {real, imag} */,
  {32'hc0371a3e, 32'hc016929a} /* (28, 4, 2) {real, imag} */,
  {32'hbeb3de0e, 32'hc0924226} /* (28, 4, 1) {real, imag} */,
  {32'h3ea11006, 32'hc018b3ec} /* (28, 4, 0) {real, imag} */,
  {32'hbe69b537, 32'hc04b7258} /* (28, 3, 31) {real, imag} */,
  {32'hc034eaa8, 32'hc0717a28} /* (28, 3, 30) {real, imag} */,
  {32'hc0813f5f, 32'hc050fcd2} /* (28, 3, 29) {real, imag} */,
  {32'hc084aaee, 32'hbfe95426} /* (28, 3, 28) {real, imag} */,
  {32'hc06dc496, 32'hc0ae48f1} /* (28, 3, 27) {real, imag} */,
  {32'hbee55cd8, 32'hc0b61a6c} /* (28, 3, 26) {real, imag} */,
  {32'hbf542c2d, 32'hc081c89e} /* (28, 3, 25) {real, imag} */,
  {32'hbe25fee7, 32'hc0addac8} /* (28, 3, 24) {real, imag} */,
  {32'hbee55a2b, 32'hc09ca7df} /* (28, 3, 23) {real, imag} */,
  {32'hc0077fb6, 32'hc0d6f37c} /* (28, 3, 22) {real, imag} */,
  {32'hbfecaef2, 32'hc0a282f0} /* (28, 3, 21) {real, imag} */,
  {32'hc01ff259, 32'hc096ccd2} /* (28, 3, 20) {real, imag} */,
  {32'hbf5f8408, 32'hc09c9f6a} /* (28, 3, 19) {real, imag} */,
  {32'hc07b46b7, 32'hc0ba6a2e} /* (28, 3, 18) {real, imag} */,
  {32'hc081f5d4, 32'hc0993e5a} /* (28, 3, 17) {real, imag} */,
  {32'hc0132f04, 32'hc007f1e8} /* (28, 3, 16) {real, imag} */,
  {32'h3fa4a7d6, 32'h4047cb5c} /* (28, 3, 15) {real, imag} */,
  {32'h4030309c, 32'h40a976f3} /* (28, 3, 14) {real, imag} */,
  {32'h4023165f, 32'h40aac019} /* (28, 3, 13) {real, imag} */,
  {32'h3f3fa6bc, 32'h40e77eb3} /* (28, 3, 12) {real, imag} */,
  {32'h4042a3de, 32'h40ff9648} /* (28, 3, 11) {real, imag} */,
  {32'h405a5c58, 32'h40d2ba78} /* (28, 3, 10) {real, imag} */,
  {32'h3fdb0d44, 32'h40cb6684} /* (28, 3, 9) {real, imag} */,
  {32'h3fdaa7b0, 32'h40c0215e} /* (28, 3, 8) {real, imag} */,
  {32'hbfe32990, 32'h40affb44} /* (28, 3, 7) {real, imag} */,
  {32'h3f10b5a2, 32'h4081226f} /* (28, 3, 6) {real, imag} */,
  {32'hbf8055ee, 32'hbf61e053} /* (28, 3, 5) {real, imag} */,
  {32'hc06f9419, 32'hc0a36c6f} /* (28, 3, 4) {real, imag} */,
  {32'h4018015c, 32'hc07777aa} /* (28, 3, 3) {real, imag} */,
  {32'hbe32d42a, 32'h3ec3974c} /* (28, 3, 2) {real, imag} */,
  {32'h3fd01547, 32'hbffbb3c0} /* (28, 3, 1) {real, imag} */,
  {32'hbec1d89d, 32'hbff7c3d2} /* (28, 3, 0) {real, imag} */,
  {32'hbf816a42, 32'hc03330d7} /* (28, 2, 31) {real, imag} */,
  {32'hbfb79e36, 32'hc0c3a1f4} /* (28, 2, 30) {real, imag} */,
  {32'hc0146bf6, 32'hc07a6ca6} /* (28, 2, 29) {real, imag} */,
  {32'hc066f9a6, 32'hc0833f3a} /* (28, 2, 28) {real, imag} */,
  {32'hc062084c, 32'hc0ab7326} /* (28, 2, 27) {real, imag} */,
  {32'hc022f3aa, 32'hc0a73f12} /* (28, 2, 26) {real, imag} */,
  {32'hc014bbdf, 32'hc06c047a} /* (28, 2, 25) {real, imag} */,
  {32'hc0211f55, 32'hc042ffc8} /* (28, 2, 24) {real, imag} */,
  {32'hbf1ffb40, 32'hc018a3ae} /* (28, 2, 23) {real, imag} */,
  {32'hbfe2c754, 32'hc0b0f66e} /* (28, 2, 22) {real, imag} */,
  {32'hbff9eb4b, 32'hc09ce697} /* (28, 2, 21) {real, imag} */,
  {32'hbf8d40a5, 32'hc093ada9} /* (28, 2, 20) {real, imag} */,
  {32'hbfb7b439, 32'hc0a0b937} /* (28, 2, 19) {real, imag} */,
  {32'hc09627f8, 32'hc0fd3d5e} /* (28, 2, 18) {real, imag} */,
  {32'hc04cac32, 32'hc0aa0a7f} /* (28, 2, 17) {real, imag} */,
  {32'hbfa4a6f6, 32'hbfc38de4} /* (28, 2, 16) {real, imag} */,
  {32'h3f96d335, 32'h404e902a} /* (28, 2, 15) {real, imag} */,
  {32'h4061350d, 32'h404a0ca2} /* (28, 2, 14) {real, imag} */,
  {32'h40b728fc, 32'h409edadb} /* (28, 2, 13) {real, imag} */,
  {32'h4046cfe2, 32'h40ae9708} /* (28, 2, 12) {real, imag} */,
  {32'h4070458a, 32'h40bc8e14} /* (28, 2, 11) {real, imag} */,
  {32'h4093a0fe, 32'h40b00e82} /* (28, 2, 10) {real, imag} */,
  {32'h403b4ce8, 32'h40bed87e} /* (28, 2, 9) {real, imag} */,
  {32'h400e5b6b, 32'h406a7a67} /* (28, 2, 8) {real, imag} */,
  {32'hbf0f33a2, 32'h40b18e08} /* (28, 2, 7) {real, imag} */,
  {32'h3faf2393, 32'h408e5d1c} /* (28, 2, 6) {real, imag} */,
  {32'h3ed6ef1c, 32'hc02822f5} /* (28, 2, 5) {real, imag} */,
  {32'hc02374a1, 32'hc0d22542} /* (28, 2, 4) {real, imag} */,
  {32'h3f3f7885, 32'hc0c7602b} /* (28, 2, 3) {real, imag} */,
  {32'hbe4ef712, 32'hc022d2d4} /* (28, 2, 2) {real, imag} */,
  {32'hbcb96ef8, 32'hc04586b4} /* (28, 2, 1) {real, imag} */,
  {32'hbfab4f36, 32'hc0091a4e} /* (28, 2, 0) {real, imag} */,
  {32'hc0057caf, 32'hbffcc127} /* (28, 1, 31) {real, imag} */,
  {32'hc025cfda, 32'hc078d922} /* (28, 1, 30) {real, imag} */,
  {32'hbfc3ae48, 32'hc0390198} /* (28, 1, 29) {real, imag} */,
  {32'hbfad28b8, 32'hc07158ae} /* (28, 1, 28) {real, imag} */,
  {32'hbfbbca7b, 32'hbfff0e14} /* (28, 1, 27) {real, imag} */,
  {32'hbfc36b72, 32'hbfc7ea62} /* (28, 1, 26) {real, imag} */,
  {32'hbf0a45f0, 32'hc0198c48} /* (28, 1, 25) {real, imag} */,
  {32'hbfd61b0a, 32'hbff5951b} /* (28, 1, 24) {real, imag} */,
  {32'hc013c9c1, 32'hc002fccf} /* (28, 1, 23) {real, imag} */,
  {32'hc03a2e55, 32'hc05f97b7} /* (28, 1, 22) {real, imag} */,
  {32'hc00b724c, 32'hc09903d4} /* (28, 1, 21) {real, imag} */,
  {32'hbf9602dc, 32'hc059f9fa} /* (28, 1, 20) {real, imag} */,
  {32'hc0633efe, 32'hc06f0a98} /* (28, 1, 19) {real, imag} */,
  {32'hc09b0667, 32'hc0c0d0f9} /* (28, 1, 18) {real, imag} */,
  {32'hc0441ec2, 32'hc08eba62} /* (28, 1, 17) {real, imag} */,
  {32'hc05d8ca6, 32'hbf9648b1} /* (28, 1, 16) {real, imag} */,
  {32'h3fa2c447, 32'h400dfb39} /* (28, 1, 15) {real, imag} */,
  {32'h4087bf1a, 32'h3fd8aa9c} /* (28, 1, 14) {real, imag} */,
  {32'h40a31a76, 32'h403801c6} /* (28, 1, 13) {real, imag} */,
  {32'h4094b97a, 32'h407278a6} /* (28, 1, 12) {real, imag} */,
  {32'h40325418, 32'h40d97ff9} /* (28, 1, 11) {real, imag} */,
  {32'h3f337f6a, 32'h40c36918} /* (28, 1, 10) {real, imag} */,
  {32'h3ee010b7, 32'h4098c4a5} /* (28, 1, 9) {real, imag} */,
  {32'h406410ae, 32'h40734d26} /* (28, 1, 8) {real, imag} */,
  {32'h400bcd64, 32'h408fc52c} /* (28, 1, 7) {real, imag} */,
  {32'hbe37ae58, 32'h40a334a4} /* (28, 1, 6) {real, imag} */,
  {32'hc002db93, 32'hbde5a610} /* (28, 1, 5) {real, imag} */,
  {32'hbfcac572, 32'hc091921d} /* (28, 1, 4) {real, imag} */,
  {32'h3e9d205f, 32'hc0aa292d} /* (28, 1, 3) {real, imag} */,
  {32'hbf7d133e, 32'hc080ce41} /* (28, 1, 2) {real, imag} */,
  {32'hbfc0aaa5, 32'hc057c38c} /* (28, 1, 1) {real, imag} */,
  {32'hbfff3f60, 32'hbf9820c2} /* (28, 1, 0) {real, imag} */,
  {32'hbf2022f7, 32'hc016a72e} /* (28, 0, 31) {real, imag} */,
  {32'hc00aa408, 32'hbfd4c7f4} /* (28, 0, 30) {real, imag} */,
  {32'hc006bc70, 32'hbfbff62e} /* (28, 0, 29) {real, imag} */,
  {32'hbf9fda7d, 32'hc00eb574} /* (28, 0, 28) {real, imag} */,
  {32'hbfdc0bbc, 32'hbf93220c} /* (28, 0, 27) {real, imag} */,
  {32'hbfa5d875, 32'hbebf8ca9} /* (28, 0, 26) {real, imag} */,
  {32'h3e941138, 32'hbfbfddb2} /* (28, 0, 25) {real, imag} */,
  {32'hbfaa8dcc, 32'hbf95e9bf} /* (28, 0, 24) {real, imag} */,
  {32'hc04339e4, 32'hc018f072} /* (28, 0, 23) {real, imag} */,
  {32'hc0437bb4, 32'hc02bdb96} /* (28, 0, 22) {real, imag} */,
  {32'hc00b4ae0, 32'hc0752c79} /* (28, 0, 21) {real, imag} */,
  {32'hbfcfcb12, 32'hc003fce7} /* (28, 0, 20) {real, imag} */,
  {32'hc03729c4, 32'hbf94a770} /* (28, 0, 19) {real, imag} */,
  {32'hc01d8a8c, 32'hbfd0cade} /* (28, 0, 18) {real, imag} */,
  {32'hbf1ae02d, 32'hbfc718f6} /* (28, 0, 17) {real, imag} */,
  {32'hbf85f9a8, 32'hbec6649a} /* (28, 0, 16) {real, imag} */,
  {32'h3f33aafe, 32'h3fd36aee} /* (28, 0, 15) {real, imag} */,
  {32'h3faab354, 32'h402dc358} /* (28, 0, 14) {real, imag} */,
  {32'hbeeef802, 32'h4055550c} /* (28, 0, 13) {real, imag} */,
  {32'h3f458595, 32'h403d2462} /* (28, 0, 12) {real, imag} */,
  {32'h3f5c8b1e, 32'h40741187} /* (28, 0, 11) {real, imag} */,
  {32'hbf83d288, 32'h4064803e} /* (28, 0, 10) {real, imag} */,
  {32'hc025a006, 32'h402951b5} /* (28, 0, 9) {real, imag} */,
  {32'h3f51d1f0, 32'h401aa48c} /* (28, 0, 8) {real, imag} */,
  {32'h3fc180dc, 32'h404eb7cd} /* (28, 0, 7) {real, imag} */,
  {32'h3f9a3c56, 32'h4077031a} /* (28, 0, 6) {real, imag} */,
  {32'hbf327cfe, 32'hbd379986} /* (28, 0, 5) {real, imag} */,
  {32'hbf46a603, 32'hbfed28e4} /* (28, 0, 4) {real, imag} */,
  {32'hbee01b5e, 32'hc07553cf} /* (28, 0, 3) {real, imag} */,
  {32'hbfea9794, 32'hc070801a} /* (28, 0, 2) {real, imag} */,
  {32'hbeed8c88, 32'hc00f4184} /* (28, 0, 1) {real, imag} */,
  {32'hbd127990, 32'hbf25bdbc} /* (28, 0, 0) {real, imag} */,
  {32'h3f86cc84, 32'h3ec18892} /* (27, 31, 31) {real, imag} */,
  {32'h3fdf1535, 32'h3ee77387} /* (27, 31, 30) {real, imag} */,
  {32'hbe061118, 32'h401076e4} /* (27, 31, 29) {real, imag} */,
  {32'h3e4449ec, 32'h3fcf2648} /* (27, 31, 28) {real, imag} */,
  {32'h400272b3, 32'h401c52d6} /* (27, 31, 27) {real, imag} */,
  {32'h402e0a5a, 32'h405accf5} /* (27, 31, 26) {real, imag} */,
  {32'h40192240, 32'h40025582} /* (27, 31, 25) {real, imag} */,
  {32'h400943aa, 32'h3fc65a0d} /* (27, 31, 24) {real, imag} */,
  {32'h3e80fc19, 32'h3f785c01} /* (27, 31, 23) {real, imag} */,
  {32'hbeafc95d, 32'h3fb0e738} /* (27, 31, 22) {real, imag} */,
  {32'hbfcb4d89, 32'hbf516cfb} /* (27, 31, 21) {real, imag} */,
  {32'hc00ff9dc, 32'hbf9f0c16} /* (27, 31, 20) {real, imag} */,
  {32'hbfc41404, 32'h3e40b88d} /* (27, 31, 19) {real, imag} */,
  {32'h3d16c210, 32'hbf4e7b24} /* (27, 31, 18) {real, imag} */,
  {32'hbf30c22c, 32'hc0238b02} /* (27, 31, 17) {real, imag} */,
  {32'h3ecf103f, 32'h3dbd2790} /* (27, 31, 16) {real, imag} */,
  {32'h3f1ae8e8, 32'h3e76c586} /* (27, 31, 15) {real, imag} */,
  {32'hbf7f3012, 32'hbd795850} /* (27, 31, 14) {real, imag} */,
  {32'h3e117bcf, 32'hbfdb5c0c} /* (27, 31, 13) {real, imag} */,
  {32'h3f48669c, 32'hc015dac6} /* (27, 31, 12) {real, imag} */,
  {32'hbe0062b2, 32'hbf99349c} /* (27, 31, 11) {real, imag} */,
  {32'h3fb7ee3c, 32'h3f478444} /* (27, 31, 10) {real, imag} */,
  {32'h3f647396, 32'h3f04af19} /* (27, 31, 9) {real, imag} */,
  {32'hbe846a9c, 32'h3f3fee78} /* (27, 31, 8) {real, imag} */,
  {32'h3ec1a468, 32'h3e9cf84a} /* (27, 31, 7) {real, imag} */,
  {32'h3e92bae4, 32'h3fc9d1da} /* (27, 31, 6) {real, imag} */,
  {32'h3e46a7e2, 32'h4013c3cd} /* (27, 31, 5) {real, imag} */,
  {32'hbf10964a, 32'h3ff121ec} /* (27, 31, 4) {real, imag} */,
  {32'h3d5d36c0, 32'h401f142d} /* (27, 31, 3) {real, imag} */,
  {32'h3e58e068, 32'h3fb91aad} /* (27, 31, 2) {real, imag} */,
  {32'hbec240d6, 32'h3fc422f1} /* (27, 31, 1) {real, imag} */,
  {32'h3f186bc4, 32'hbd8533d6} /* (27, 31, 0) {real, imag} */,
  {32'h3f84cf59, 32'h3f0e53aa} /* (27, 30, 31) {real, imag} */,
  {32'h403ef993, 32'h3fdfa33c} /* (27, 30, 30) {real, imag} */,
  {32'h3fc3f0b0, 32'h40603b9a} /* (27, 30, 29) {real, imag} */,
  {32'h3f76e93e, 32'h4008fe3c} /* (27, 30, 28) {real, imag} */,
  {32'h3fc7d8d8, 32'h407db2b7} /* (27, 30, 27) {real, imag} */,
  {32'h3f4f42b5, 32'h409bb444} /* (27, 30, 26) {real, imag} */,
  {32'h3fcb3439, 32'h4056957e} /* (27, 30, 25) {real, imag} */,
  {32'h3ff34eec, 32'h402c00f8} /* (27, 30, 24) {real, imag} */,
  {32'h40185fcd, 32'h4021d02c} /* (27, 30, 23) {real, imag} */,
  {32'h4047c284, 32'h3fe1f5e0} /* (27, 30, 22) {real, imag} */,
  {32'hbf2d82d2, 32'hbf4b33ce} /* (27, 30, 21) {real, imag} */,
  {32'hc08e1466, 32'hc0695309} /* (27, 30, 20) {real, imag} */,
  {32'hc0b3e85e, 32'hbfbe79b5} /* (27, 30, 19) {real, imag} */,
  {32'hbfaae44a, 32'hc036ecee} /* (27, 30, 18) {real, imag} */,
  {32'hbef71f6e, 32'hc0953d31} /* (27, 30, 17) {real, imag} */,
  {32'h3f72d973, 32'hc056221a} /* (27, 30, 16) {real, imag} */,
  {32'hbf7ec28f, 32'hbffafb1e} /* (27, 30, 15) {real, imag} */,
  {32'hbf9133e2, 32'hbf3bc508} /* (27, 30, 14) {real, imag} */,
  {32'hbd1c2910, 32'hbfe4e679} /* (27, 30, 13) {real, imag} */,
  {32'hbf51f00d, 32'hc081ff34} /* (27, 30, 12) {real, imag} */,
  {32'hbfda083e, 32'hc06bdefe} /* (27, 30, 11) {real, imag} */,
  {32'h401726ff, 32'h3ebe7211} /* (27, 30, 10) {real, imag} */,
  {32'h400a81f4, 32'h3ffd28a0} /* (27, 30, 9) {real, imag} */,
  {32'hbec4d87c, 32'h400afbf8} /* (27, 30, 8) {real, imag} */,
  {32'h3f1581db, 32'h3fec728a} /* (27, 30, 7) {real, imag} */,
  {32'h3fd99ea3, 32'h404d6876} /* (27, 30, 6) {real, imag} */,
  {32'h3e6ac088, 32'h408a3f40} /* (27, 30, 5) {real, imag} */,
  {32'h3ea2e182, 32'h4010faf4} /* (27, 30, 4) {real, imag} */,
  {32'hbea90298, 32'h3fee4112} /* (27, 30, 3) {real, imag} */,
  {32'h402b34f2, 32'h3ee70914} /* (27, 30, 2) {real, imag} */,
  {32'h3d264f70, 32'h40074ee2} /* (27, 30, 1) {real, imag} */,
  {32'hbf5523e6, 32'h3f897266} /* (27, 30, 0) {real, imag} */,
  {32'h3eac693a, 32'h3fb690a5} /* (27, 29, 31) {real, imag} */,
  {32'h403013f3, 32'h40469abe} /* (27, 29, 30) {real, imag} */,
  {32'h40139ecc, 32'h403b58cc} /* (27, 29, 29) {real, imag} */,
  {32'h3fb49807, 32'h40269228} /* (27, 29, 28) {real, imag} */,
  {32'h3fe2c84f, 32'h40686954} /* (27, 29, 27) {real, imag} */,
  {32'hbf78120f, 32'h4035d4ad} /* (27, 29, 26) {real, imag} */,
  {32'h3d8c4a38, 32'h4064729d} /* (27, 29, 25) {real, imag} */,
  {32'h3f483d04, 32'h401497dc} /* (27, 29, 24) {real, imag} */,
  {32'h400b5a68, 32'h3f901336} /* (27, 29, 23) {real, imag} */,
  {32'h3f963edf, 32'hbeea6be8} /* (27, 29, 22) {real, imag} */,
  {32'hbe1cca98, 32'h3fd19d8c} /* (27, 29, 21) {real, imag} */,
  {32'hbff7ec54, 32'hbf256b10} /* (27, 29, 20) {real, imag} */,
  {32'hc0c807c5, 32'h3e4917c0} /* (27, 29, 19) {real, imag} */,
  {32'hc077175b, 32'hbf0bf190} /* (27, 29, 18) {real, imag} */,
  {32'hc07f163e, 32'hc03e8162} /* (27, 29, 17) {real, imag} */,
  {32'hc05c6a56, 32'hc0963db2} /* (27, 29, 16) {real, imag} */,
  {32'hbfe81e9c, 32'hc08881bb} /* (27, 29, 15) {real, imag} */,
  {32'h3fcdfa14, 32'hc005201e} /* (27, 29, 14) {real, imag} */,
  {32'hbe68e174, 32'hbee8178a} /* (27, 29, 13) {real, imag} */,
  {32'hc0592792, 32'hc0012244} /* (27, 29, 12) {real, imag} */,
  {32'hc04ae31e, 32'hbffaecaf} /* (27, 29, 11) {real, imag} */,
  {32'h3f5a3e72, 32'h3f9c822c} /* (27, 29, 10) {real, imag} */,
  {32'h408c797d, 32'h3fdc052d} /* (27, 29, 9) {real, imag} */,
  {32'h4017080c, 32'h403076fc} /* (27, 29, 8) {real, imag} */,
  {32'h3f8944ba, 32'h404fb234} /* (27, 29, 7) {real, imag} */,
  {32'h40402ec6, 32'h3ff71c51} /* (27, 29, 6) {real, imag} */,
  {32'h404a4d4e, 32'h4070715c} /* (27, 29, 5) {real, imag} */,
  {32'h3ffa049e, 32'h40007e30} /* (27, 29, 4) {real, imag} */,
  {32'hbe76a1d6, 32'h400d697d} /* (27, 29, 3) {real, imag} */,
  {32'h4084f2d5, 32'h3fb76f5c} /* (27, 29, 2) {real, imag} */,
  {32'h40774c0b, 32'h4012e410} /* (27, 29, 1) {real, imag} */,
  {32'h3f3bfebc, 32'h4018f62d} /* (27, 29, 0) {real, imag} */,
  {32'h3f617fca, 32'h3fbb3e70} /* (27, 28, 31) {real, imag} */,
  {32'h3fcaca16, 32'h40264b7d} /* (27, 28, 30) {real, imag} */,
  {32'h3f172494, 32'h3f2d0948} /* (27, 28, 29) {real, imag} */,
  {32'h3fed6410, 32'h3fbfcb25} /* (27, 28, 28) {real, imag} */,
  {32'h4052ee49, 32'h3fa9f988} /* (27, 28, 27) {real, imag} */,
  {32'hbfd264b4, 32'h3f5f834a} /* (27, 28, 26) {real, imag} */,
  {32'hbfce88dd, 32'h3ff114db} /* (27, 28, 25) {real, imag} */,
  {32'hbe3c6f24, 32'h406968d9} /* (27, 28, 24) {real, imag} */,
  {32'h3f44635e, 32'h3fc67ffd} /* (27, 28, 23) {real, imag} */,
  {32'hbfabd2dd, 32'hbe1fcad4} /* (27, 28, 22) {real, imag} */,
  {32'hbfb48f46, 32'h40263ea8} /* (27, 28, 21) {real, imag} */,
  {32'hbfb2e1f1, 32'h400bc9fa} /* (27, 28, 20) {real, imag} */,
  {32'hc00b04c0, 32'h3f848c65} /* (27, 28, 19) {real, imag} */,
  {32'hc02add5e, 32'hbf2466e0} /* (27, 28, 18) {real, imag} */,
  {32'hc02068b6, 32'hc00a1dc2} /* (27, 28, 17) {real, imag} */,
  {32'hc062d24b, 32'hc0525abb} /* (27, 28, 16) {real, imag} */,
  {32'hc05bf708, 32'hc03643f4} /* (27, 28, 15) {real, imag} */,
  {32'hbf75b00e, 32'hbffa04ba} /* (27, 28, 14) {real, imag} */,
  {32'hbfc31d9c, 32'hbfb88b75} /* (27, 28, 13) {real, imag} */,
  {32'hbfeae1b2, 32'hbfb7da6a} /* (27, 28, 12) {real, imag} */,
  {32'hbfc9528b, 32'hc0898ff2} /* (27, 28, 11) {real, imag} */,
  {32'hbf48390c, 32'h3f39d560} /* (27, 28, 10) {real, imag} */,
  {32'h401bb740, 32'h408636b8} /* (27, 28, 9) {real, imag} */,
  {32'h401b073e, 32'h40524066} /* (27, 28, 8) {real, imag} */,
  {32'h3ff5b338, 32'h400b2f2f} /* (27, 28, 7) {real, imag} */,
  {32'h403877ea, 32'h3fe976f3} /* (27, 28, 6) {real, imag} */,
  {32'h401057ce, 32'h40559e44} /* (27, 28, 5) {real, imag} */,
  {32'h3f68ac31, 32'h3f9133e2} /* (27, 28, 4) {real, imag} */,
  {32'h3fe66992, 32'h404547ac} /* (27, 28, 3) {real, imag} */,
  {32'h40853d8c, 32'h4044ef97} /* (27, 28, 2) {real, imag} */,
  {32'h3feaa412, 32'h3fe7bd43} /* (27, 28, 1) {real, imag} */,
  {32'hbe56d964, 32'h3fb0f1cc} /* (27, 28, 0) {real, imag} */,
  {32'h3f7b3a48, 32'h3f6c4fd9} /* (27, 27, 31) {real, imag} */,
  {32'h3f16a2c1, 32'h3faefa26} /* (27, 27, 30) {real, imag} */,
  {32'hbfe71616, 32'hbf82894f} /* (27, 27, 29) {real, imag} */,
  {32'h40163643, 32'h3edb9452} /* (27, 27, 28) {real, imag} */,
  {32'h406a91b2, 32'hbd0596e0} /* (27, 27, 27) {real, imag} */,
  {32'hbf5a5545, 32'h400f00c0} /* (27, 27, 26) {real, imag} */,
  {32'hc06ac3c8, 32'h408fcddc} /* (27, 27, 25) {real, imag} */,
  {32'hbeb959ee, 32'h408b3c8a} /* (27, 27, 24) {real, imag} */,
  {32'h3fe1e5a8, 32'h3f81f666} /* (27, 27, 23) {real, imag} */,
  {32'h4012a858, 32'h3f8c68d0} /* (27, 27, 22) {real, imag} */,
  {32'hbde9f658, 32'h408b4374} /* (27, 27, 21) {real, imag} */,
  {32'hbf5e20b8, 32'h3f8cf9cc} /* (27, 27, 20) {real, imag} */,
  {32'hbf7034a0, 32'hbec8a6a4} /* (27, 27, 19) {real, imag} */,
  {32'hc05ac066, 32'hc04d423a} /* (27, 27, 18) {real, imag} */,
  {32'hbfe1e0fe, 32'hc080ad29} /* (27, 27, 17) {real, imag} */,
  {32'h3f25248e, 32'hc06f8716} /* (27, 27, 16) {real, imag} */,
  {32'hc015c8a5, 32'hbfe63150} /* (27, 27, 15) {real, imag} */,
  {32'hbf6964c5, 32'h3be30a80} /* (27, 27, 14) {real, imag} */,
  {32'hbfdcb2f4, 32'hbf90b8b6} /* (27, 27, 13) {real, imag} */,
  {32'hc05790d0, 32'hc0449b74} /* (27, 27, 12) {real, imag} */,
  {32'hc01ed7d3, 32'hc0a2e0d2} /* (27, 27, 11) {real, imag} */,
  {32'h3c7ee200, 32'h3fca3089} /* (27, 27, 10) {real, imag} */,
  {32'hbfabe7f8, 32'h409d59cc} /* (27, 27, 9) {real, imag} */,
  {32'h3f7e882e, 32'h401038d8} /* (27, 27, 8) {real, imag} */,
  {32'h3f9ed8a5, 32'h3fe2430b} /* (27, 27, 7) {real, imag} */,
  {32'h3fd24db8, 32'h3fa1bd2c} /* (27, 27, 6) {real, imag} */,
  {32'hbf42fa43, 32'h408011a2} /* (27, 27, 5) {real, imag} */,
  {32'hbf68ab9a, 32'h408a0eb0} /* (27, 27, 4) {real, imag} */,
  {32'h3fe5767e, 32'h40531c10} /* (27, 27, 3) {real, imag} */,
  {32'h401cb186, 32'h3f7bdf4b} /* (27, 27, 2) {real, imag} */,
  {32'h3fe465d5, 32'h3f993498} /* (27, 27, 1) {real, imag} */,
  {32'h3f86490c, 32'h3f84c6a6} /* (27, 27, 0) {real, imag} */,
  {32'hbdd2ddba, 32'h3f13bff3} /* (27, 26, 31) {real, imag} */,
  {32'hbf05eca5, 32'hbf10cc74} /* (27, 26, 30) {real, imag} */,
  {32'hc01b01ae, 32'hbe35e1cc} /* (27, 26, 29) {real, imag} */,
  {32'hbc8b8d40, 32'h3fa20009} /* (27, 26, 28) {real, imag} */,
  {32'h403404e4, 32'hbef7dccc} /* (27, 26, 27) {real, imag} */,
  {32'h403f66f5, 32'h40897228} /* (27, 26, 26) {real, imag} */,
  {32'h3f7fdb84, 32'h408bb020} /* (27, 26, 25) {real, imag} */,
  {32'h3ffd8e05, 32'h3f645638} /* (27, 26, 24) {real, imag} */,
  {32'h404cc058, 32'h3f350f48} /* (27, 26, 23) {real, imag} */,
  {32'h401c9db9, 32'h3f9d531c} /* (27, 26, 22) {real, imag} */,
  {32'hbfb22e0c, 32'h403d8ae0} /* (27, 26, 21) {real, imag} */,
  {32'hbfadc356, 32'hbf48670e} /* (27, 26, 20) {real, imag} */,
  {32'hbded7c98, 32'hbff3ec7e} /* (27, 26, 19) {real, imag} */,
  {32'hbf9d4ea8, 32'hc08433c2} /* (27, 26, 18) {real, imag} */,
  {32'hbfd31cbb, 32'hc0602168} /* (27, 26, 17) {real, imag} */,
  {32'h3f32119e, 32'hc05948c0} /* (27, 26, 16) {real, imag} */,
  {32'hbfb57610, 32'hc017422f} /* (27, 26, 15) {real, imag} */,
  {32'hc00a2265, 32'hc004edc6} /* (27, 26, 14) {real, imag} */,
  {32'hbfcf7d2c, 32'hbfb2f8fa} /* (27, 26, 13) {real, imag} */,
  {32'hc01f66b2, 32'hbf36209d} /* (27, 26, 12) {real, imag} */,
  {32'hc023c0d3, 32'hbead35ac} /* (27, 26, 11) {real, imag} */,
  {32'h3e04fb38, 32'h402354b9} /* (27, 26, 10) {real, imag} */,
  {32'h3e706dd8, 32'h3f962cc4} /* (27, 26, 9) {real, imag} */,
  {32'hbe3ec0e2, 32'h3ff0647c} /* (27, 26, 8) {real, imag} */,
  {32'h3e84f96a, 32'h40069af8} /* (27, 26, 7) {real, imag} */,
  {32'h3f88b21e, 32'h3f45c97c} /* (27, 26, 6) {real, imag} */,
  {32'h3eff166c, 32'h40791ec7} /* (27, 26, 5) {real, imag} */,
  {32'hbc2b3f00, 32'h40863e82} /* (27, 26, 4) {real, imag} */,
  {32'hbf5a82a3, 32'h3fd7da05} /* (27, 26, 3) {real, imag} */,
  {32'h3f3515cc, 32'h3e57b9d0} /* (27, 26, 2) {real, imag} */,
  {32'h3cb14c80, 32'h3e60c904} /* (27, 26, 1) {real, imag} */,
  {32'hbfb05ca9, 32'h3f22527a} /* (27, 26, 0) {real, imag} */,
  {32'hbea50bbe, 32'h3fdad0b0} /* (27, 25, 31) {real, imag} */,
  {32'h3ed8299e, 32'h401df9ae} /* (27, 25, 30) {real, imag} */,
  {32'h3e291f1c, 32'h40405598} /* (27, 25, 29) {real, imag} */,
  {32'h3ebaf7a8, 32'h40233f50} /* (27, 25, 28) {real, imag} */,
  {32'h3fe35c29, 32'h3fc49e83} /* (27, 25, 27) {real, imag} */,
  {32'h401661bc, 32'h40179c18} /* (27, 25, 26) {real, imag} */,
  {32'h4033b69a, 32'h3fa5d505} /* (27, 25, 25) {real, imag} */,
  {32'h4099294c, 32'h3fe92160} /* (27, 25, 24) {real, imag} */,
  {32'h4065d8e1, 32'h40708824} /* (27, 25, 23) {real, imag} */,
  {32'h403252f2, 32'h3fd297c3} /* (27, 25, 22) {real, imag} */,
  {32'h3ef8cc02, 32'h3fe430b1} /* (27, 25, 21) {real, imag} */,
  {32'h3ecf66f0, 32'hc03dbfe2} /* (27, 25, 20) {real, imag} */,
  {32'hbede3cb6, 32'hc08650cd} /* (27, 25, 19) {real, imag} */,
  {32'hbf73c6bc, 32'hbe67f078} /* (27, 25, 18) {real, imag} */,
  {32'hc06de39c, 32'h3f9f934b} /* (27, 25, 17) {real, imag} */,
  {32'hc03a45dd, 32'h3f102759} /* (27, 25, 16) {real, imag} */,
  {32'hc00ad25a, 32'hbfe32046} /* (27, 25, 15) {real, imag} */,
  {32'hbf20b0be, 32'hc0447947} /* (27, 25, 14) {real, imag} */,
  {32'hbf187ffb, 32'hc04ff002} /* (27, 25, 13) {real, imag} */,
  {32'hc0536004, 32'hbf1afee6} /* (27, 25, 12) {real, imag} */,
  {32'hc0804fb3, 32'h3f892b52} /* (27, 25, 11) {real, imag} */,
  {32'h3f1e9a15, 32'h403a9ab2} /* (27, 25, 10) {real, imag} */,
  {32'h3e297358, 32'h3fa22f7e} /* (27, 25, 9) {real, imag} */,
  {32'hbff52631, 32'h407e4d78} /* (27, 25, 8) {real, imag} */,
  {32'hbfc7c368, 32'h400ad3f1} /* (27, 25, 7) {real, imag} */,
  {32'h3e0cc50a, 32'hbe9079ce} /* (27, 25, 6) {real, imag} */,
  {32'h3ffa22d5, 32'h3f61c766} /* (27, 25, 5) {real, imag} */,
  {32'h3c5fb040, 32'h402ce42f} /* (27, 25, 4) {real, imag} */,
  {32'h3f2a00b6, 32'h4007b8f2} /* (27, 25, 3) {real, imag} */,
  {32'h40121e04, 32'h3f71582e} /* (27, 25, 2) {real, imag} */,
  {32'h3d5a7c00, 32'h4028b508} /* (27, 25, 1) {real, imag} */,
  {32'hbff4e120, 32'h3fc0696e} /* (27, 25, 0) {real, imag} */,
  {32'h3f9e26fc, 32'h3faa045e} /* (27, 24, 31) {real, imag} */,
  {32'h40324540, 32'h3fda1b0c} /* (27, 24, 30) {real, imag} */,
  {32'h40894b38, 32'h402d4d2c} /* (27, 24, 29) {real, imag} */,
  {32'h409c6304, 32'h40a3fd18} /* (27, 24, 28) {real, imag} */,
  {32'h40853ceb, 32'h409bfb37} /* (27, 24, 27) {real, imag} */,
  {32'h4025f578, 32'h4033106b} /* (27, 24, 26) {real, imag} */,
  {32'h401a6100, 32'h3fd5aa58} /* (27, 24, 25) {real, imag} */,
  {32'h4062e0c8, 32'h403606c8} /* (27, 24, 24) {real, imag} */,
  {32'h4004a277, 32'h40915d39} /* (27, 24, 23) {real, imag} */,
  {32'h408224ae, 32'h405779ac} /* (27, 24, 22) {real, imag} */,
  {32'h401338b7, 32'h40206b7e} /* (27, 24, 21) {real, imag} */,
  {32'h4037f372, 32'hbe7cd9ac} /* (27, 24, 20) {real, imag} */,
  {32'h3e778f74, 32'hc021a59a} /* (27, 24, 19) {real, imag} */,
  {32'hbfe8aec6, 32'h3f91f51a} /* (27, 24, 18) {real, imag} */,
  {32'hc0ceaeea, 32'h3ff8ec70} /* (27, 24, 17) {real, imag} */,
  {32'hc0cdd1cc, 32'hbf1dfd22} /* (27, 24, 16) {real, imag} */,
  {32'hc001fdbf, 32'hc0966f56} /* (27, 24, 15) {real, imag} */,
  {32'hbedb4bc8, 32'hc09c51cc} /* (27, 24, 14) {real, imag} */,
  {32'hc06f6c90, 32'hc08a9f2a} /* (27, 24, 13) {real, imag} */,
  {32'hc0cc2a86, 32'hbfecc373} /* (27, 24, 12) {real, imag} */,
  {32'hc054c62e, 32'hc001efea} /* (27, 24, 11) {real, imag} */,
  {32'hbec5ac72, 32'h3f9de423} /* (27, 24, 10) {real, imag} */,
  {32'h3de6bbf0, 32'h40538ce9} /* (27, 24, 9) {real, imag} */,
  {32'hbfbdf01b, 32'h40b205be} /* (27, 24, 8) {real, imag} */,
  {32'hbfe27e3d, 32'h401d7590} /* (27, 24, 7) {real, imag} */,
  {32'hbfd5290a, 32'hbeb95e05} /* (27, 24, 6) {real, imag} */,
  {32'h3f1c528a, 32'hbfcd81ee} /* (27, 24, 5) {real, imag} */,
  {32'hbf58b49a, 32'h3f1d88a0} /* (27, 24, 4) {real, imag} */,
  {32'h3e6aec5e, 32'h3f94ad00} /* (27, 24, 3) {real, imag} */,
  {32'h3f8ae594, 32'h3f890978} /* (27, 24, 2) {real, imag} */,
  {32'h3f874a58, 32'h4059e61c} /* (27, 24, 1) {real, imag} */,
  {32'h3c8847f0, 32'h3fa93d4c} /* (27, 24, 0) {real, imag} */,
  {32'h40064b23, 32'h3f39e86e} /* (27, 23, 31) {real, imag} */,
  {32'h408c7ee6, 32'h3f66ddaa} /* (27, 23, 30) {real, imag} */,
  {32'h40475b7a, 32'h40393d30} /* (27, 23, 29) {real, imag} */,
  {32'h40529a1d, 32'h40c003db} /* (27, 23, 28) {real, imag} */,
  {32'h40ae55d3, 32'h40b725ba} /* (27, 23, 27) {real, imag} */,
  {32'h404b6b4c, 32'h404a17bc} /* (27, 23, 26) {real, imag} */,
  {32'h40084dca, 32'h3fb459fb} /* (27, 23, 25) {real, imag} */,
  {32'h3f881d44, 32'h402e06a1} /* (27, 23, 24) {real, imag} */,
  {32'h401e604b, 32'h408ce065} /* (27, 23, 23) {real, imag} */,
  {32'h40119e70, 32'h408b3d0d} /* (27, 23, 22) {real, imag} */,
  {32'hbf26c9b8, 32'h3f3866fb} /* (27, 23, 21) {real, imag} */,
  {32'h3f19816c, 32'hbf1847c8} /* (27, 23, 20) {real, imag} */,
  {32'h40027994, 32'hbf9f5d29} /* (27, 23, 19) {real, imag} */,
  {32'h3f679f60, 32'hc0134334} /* (27, 23, 18) {real, imag} */,
  {32'hc03fd97e, 32'hc051ad1a} /* (27, 23, 17) {real, imag} */,
  {32'hc028893e, 32'hc0321930} /* (27, 23, 16) {real, imag} */,
  {32'hbf2e1a33, 32'hc0a53cb6} /* (27, 23, 15) {real, imag} */,
  {32'hc04ca205, 32'hc0abdc34} /* (27, 23, 14) {real, imag} */,
  {32'hc0a18c83, 32'hc081bd93} /* (27, 23, 13) {real, imag} */,
  {32'hc06f949a, 32'hc0679e6a} /* (27, 23, 12) {real, imag} */,
  {32'hbf5340e3, 32'hbf44e1b2} /* (27, 23, 11) {real, imag} */,
  {32'hbf4a020c, 32'h4017c142} /* (27, 23, 10) {real, imag} */,
  {32'hbe8c3c52, 32'h407d8856} /* (27, 23, 9) {real, imag} */,
  {32'h3fce7fe9, 32'h40ad3b93} /* (27, 23, 8) {real, imag} */,
  {32'h3ebfcf5e, 32'h40835c7e} /* (27, 23, 7) {real, imag} */,
  {32'hbfa346b3, 32'h40461a3e} /* (27, 23, 6) {real, imag} */,
  {32'hbf5e54e9, 32'h403e9627} /* (27, 23, 5) {real, imag} */,
  {32'hc00cefaf, 32'hbda93270} /* (27, 23, 4) {real, imag} */,
  {32'h3e0c81a2, 32'hbe207404} /* (27, 23, 3) {real, imag} */,
  {32'h3f4e81df, 32'h3fb9f427} /* (27, 23, 2) {real, imag} */,
  {32'h3e518e70, 32'hbe8c7bbe} /* (27, 23, 1) {real, imag} */,
  {32'h3f8577e5, 32'hbe1d6988} /* (27, 23, 0) {real, imag} */,
  {32'h3fbe1450, 32'h4032c3e6} /* (27, 22, 31) {real, imag} */,
  {32'h402357ba, 32'h4076e3da} /* (27, 22, 30) {real, imag} */,
  {32'h3fa8f815, 32'h40bd2944} /* (27, 22, 29) {real, imag} */,
  {32'h3f7865aa, 32'h40a09120} /* (27, 22, 28) {real, imag} */,
  {32'h40364efb, 32'h407775be} /* (27, 22, 27) {real, imag} */,
  {32'h3fb9fe74, 32'h40476152} /* (27, 22, 26) {real, imag} */,
  {32'h3fb75e98, 32'h3fa09e06} /* (27, 22, 25) {real, imag} */,
  {32'h3f6c822a, 32'h40269e8c} /* (27, 22, 24) {real, imag} */,
  {32'h40481868, 32'h404d140b} /* (27, 22, 23) {real, imag} */,
  {32'h403a02a2, 32'h4049f1e1} /* (27, 22, 22) {real, imag} */,
  {32'hbef73f8c, 32'h3e46df52} /* (27, 22, 21) {real, imag} */,
  {32'hc00119be, 32'hbf59672c} /* (27, 22, 20) {real, imag} */,
  {32'hbf3ebde0, 32'hc005428c} /* (27, 22, 19) {real, imag} */,
  {32'hbe356b48, 32'hc0781bea} /* (27, 22, 18) {real, imag} */,
  {32'hc00b200b, 32'hc06bd553} /* (27, 22, 17) {real, imag} */,
  {32'hbe975bc6, 32'hbf9589a0} /* (27, 22, 16) {real, imag} */,
  {32'h3ef852cd, 32'hbfafae8a} /* (27, 22, 15) {real, imag} */,
  {32'hbfabdfbb, 32'hbfcd873b} /* (27, 22, 14) {real, imag} */,
  {32'hbf5e04f2, 32'hbec9e12a} /* (27, 22, 13) {real, imag} */,
  {32'hc009a80b, 32'h3f15f522} /* (27, 22, 12) {real, imag} */,
  {32'hbfad9bc8, 32'h3fb63c12} /* (27, 22, 11) {real, imag} */,
  {32'h3ec6d3a8, 32'h402cdeaa} /* (27, 22, 10) {real, imag} */,
  {32'h4023f948, 32'h3fd04b04} /* (27, 22, 9) {real, imag} */,
  {32'h409ba3a3, 32'h406b1e3e} /* (27, 22, 8) {real, imag} */,
  {32'h404138e8, 32'h40631773} /* (27, 22, 7) {real, imag} */,
  {32'h3ffdd81f, 32'h4051df24} /* (27, 22, 6) {real, imag} */,
  {32'h3f590478, 32'h406c9183} /* (27, 22, 5) {real, imag} */,
  {32'hbf82ba8e, 32'h3f33b62f} /* (27, 22, 4) {real, imag} */,
  {32'h3d1c3d30, 32'h3f41d6ed} /* (27, 22, 3) {real, imag} */,
  {32'hbf023496, 32'h3f25a06e} /* (27, 22, 2) {real, imag} */,
  {32'h3ee1f0a4, 32'hbf26daa6} /* (27, 22, 1) {real, imag} */,
  {32'h3f748112, 32'h3f423fb0} /* (27, 22, 0) {real, imag} */,
  {32'hbfa417f5, 32'h3f859949} /* (27, 21, 31) {real, imag} */,
  {32'hbf8ce5e8, 32'h4022b9f6} /* (27, 21, 30) {real, imag} */,
  {32'h3ef65c7a, 32'h406357ec} /* (27, 21, 29) {real, imag} */,
  {32'h3fb8c68a, 32'hbef9b606} /* (27, 21, 28) {real, imag} */,
  {32'h4012a3ec, 32'h401831ee} /* (27, 21, 27) {real, imag} */,
  {32'h3f5b9422, 32'h3febe71c} /* (27, 21, 26) {real, imag} */,
  {32'hbf8ba480, 32'h3eec1d1b} /* (27, 21, 25) {real, imag} */,
  {32'hbf995bd6, 32'h3f5b9ce8} /* (27, 21, 24) {real, imag} */,
  {32'h3e8dab0b, 32'h3f2284e4} /* (27, 21, 23) {real, imag} */,
  {32'h3fc7282c, 32'h3ff0abd8} /* (27, 21, 22) {real, imag} */,
  {32'h3e07a1c8, 32'h4005a818} /* (27, 21, 21) {real, imag} */,
  {32'hbf6190a8, 32'hbe073d18} /* (27, 21, 20) {real, imag} */,
  {32'hbf9463c9, 32'hc00558cb} /* (27, 21, 19) {real, imag} */,
  {32'h3efa5824, 32'hbf8ad3a3} /* (27, 21, 18) {real, imag} */,
  {32'hbf9b7078, 32'h3a8b6a00} /* (27, 21, 17) {real, imag} */,
  {32'hbf09fa4d, 32'h3f5318ea} /* (27, 21, 16) {real, imag} */,
  {32'h3f19a8a0, 32'hbdf89c78} /* (27, 21, 15) {real, imag} */,
  {32'h3f88b9ba, 32'hbf7d8e3a} /* (27, 21, 14) {real, imag} */,
  {32'h3f95a7f1, 32'h3f6939f8} /* (27, 21, 13) {real, imag} */,
  {32'h3f0142cc, 32'h3e8166f0} /* (27, 21, 12) {real, imag} */,
  {32'hbf190370, 32'h3ec59360} /* (27, 21, 11) {real, imag} */,
  {32'hbfbfaf15, 32'h3f3c2926} /* (27, 21, 10) {real, imag} */,
  {32'hbe7333c6, 32'h4001624d} /* (27, 21, 9) {real, imag} */,
  {32'h409267e3, 32'h3fa20f76} /* (27, 21, 8) {real, imag} */,
  {32'h3ff9ee27, 32'h3fc6d0f0} /* (27, 21, 7) {real, imag} */,
  {32'h4031e47b, 32'h3f90c6a0} /* (27, 21, 6) {real, imag} */,
  {32'h3fea4cd6, 32'hbeb8a38c} /* (27, 21, 5) {real, imag} */,
  {32'h3f727290, 32'h3e8f52ee} /* (27, 21, 4) {real, imag} */,
  {32'h4046c22c, 32'h3fff36e3} /* (27, 21, 3) {real, imag} */,
  {32'h3faecdff, 32'hbfb707e5} /* (27, 21, 2) {real, imag} */,
  {32'h3f70d256, 32'hbfea2d10} /* (27, 21, 1) {real, imag} */,
  {32'h3f35a54c, 32'h3eaf68be} /* (27, 21, 0) {real, imag} */,
  {32'hc005738a, 32'hbfdd2c67} /* (27, 20, 31) {real, imag} */,
  {32'hc0509a6c, 32'hbf78c875} /* (27, 20, 30) {real, imag} */,
  {32'hbff0eeef, 32'h3f1f7a7e} /* (27, 20, 29) {real, imag} */,
  {32'hbda99b78, 32'hc0340606} /* (27, 20, 28) {real, imag} */,
  {32'h3f49a0f2, 32'hc0068338} /* (27, 20, 27) {real, imag} */,
  {32'hbf8ad6ce, 32'hc0369dfb} /* (27, 20, 26) {real, imag} */,
  {32'hc05f89b7, 32'hbf73980e} /* (27, 20, 25) {real, imag} */,
  {32'hbff07ae6, 32'h3ee0d208} /* (27, 20, 24) {real, imag} */,
  {32'hbff575db, 32'hc03a52d2} /* (27, 20, 23) {real, imag} */,
  {32'hbe89f4d8, 32'hbfa16870} /* (27, 20, 22) {real, imag} */,
  {32'h3f2fe53e, 32'h3ef003dc} /* (27, 20, 21) {real, imag} */,
  {32'h3f0d0244, 32'h40033f3f} /* (27, 20, 20) {real, imag} */,
  {32'h3e28bee8, 32'h3e9123ba} /* (27, 20, 19) {real, imag} */,
  {32'h4056b254, 32'h3ebd7fdc} /* (27, 20, 18) {real, imag} */,
  {32'h405cb2f8, 32'h3f0450c1} /* (27, 20, 17) {real, imag} */,
  {32'h3f867684, 32'h40271159} /* (27, 20, 16) {real, imag} */,
  {32'hc0163712, 32'h3eaee06f} /* (27, 20, 15) {real, imag} */,
  {32'hbf929415, 32'h3f7051e3} /* (27, 20, 14) {real, imag} */,
  {32'hbed5fdb6, 32'h3facb945} /* (27, 20, 13) {real, imag} */,
  {32'h3f652dc3, 32'h3f8742e9} /* (27, 20, 12) {real, imag} */,
  {32'hbff8a86a, 32'h3fbe3521} /* (27, 20, 11) {real, imag} */,
  {32'hc08ed6b8, 32'hc0011ad9} /* (27, 20, 10) {real, imag} */,
  {32'hc059d288, 32'hbfba0c3c} /* (27, 20, 9) {real, imag} */,
  {32'h3f8577ba, 32'hc04b2da6} /* (27, 20, 8) {real, imag} */,
  {32'hbf8c3b9d, 32'hc023c44c} /* (27, 20, 7) {real, imag} */,
  {32'hbf129df8, 32'hbfa4dfe0} /* (27, 20, 6) {real, imag} */,
  {32'hbfe04136, 32'hc02e4475} /* (27, 20, 5) {real, imag} */,
  {32'hbff70ed4, 32'hbf998cbe} /* (27, 20, 4) {real, imag} */,
  {32'hbecc63b8, 32'h3ecf7d98} /* (27, 20, 3) {real, imag} */,
  {32'h3dc33938, 32'hc03ee305} /* (27, 20, 2) {real, imag} */,
  {32'h3f4ebf28, 32'hc0897aef} /* (27, 20, 1) {real, imag} */,
  {32'hbe1886f6, 32'hc00a84e2} /* (27, 20, 0) {real, imag} */,
  {32'h3fbb4fb1, 32'hbf769471} /* (27, 19, 31) {real, imag} */,
  {32'h3fbb565f, 32'hbf8ba292} /* (27, 19, 30) {real, imag} */,
  {32'h3f3b7331, 32'h3f010fa9} /* (27, 19, 29) {real, imag} */,
  {32'h3eced446, 32'hbf333b48} /* (27, 19, 28) {real, imag} */,
  {32'h3dec14b8, 32'hc0312b0f} /* (27, 19, 27) {real, imag} */,
  {32'hbf8a2f38, 32'hc01969dc} /* (27, 19, 26) {real, imag} */,
  {32'hc012c232, 32'h3df75020} /* (27, 19, 25) {real, imag} */,
  {32'hbfe2b922, 32'h3e722c30} /* (27, 19, 24) {real, imag} */,
  {32'hc045706a, 32'hbff525cd} /* (27, 19, 23) {real, imag} */,
  {32'hbfc06eea, 32'hc007cac6} /* (27, 19, 22) {real, imag} */,
  {32'hbd5d6be4, 32'h3e6d8418} /* (27, 19, 21) {real, imag} */,
  {32'h3f8b50ee, 32'h405b5527} /* (27, 19, 20) {real, imag} */,
  {32'h4023c4d4, 32'h4066beb8} /* (27, 19, 19) {real, imag} */,
  {32'h40638130, 32'hbe27bbb8} /* (27, 19, 18) {real, imag} */,
  {32'h402f2ce1, 32'h3f100b96} /* (27, 19, 17) {real, imag} */,
  {32'h3ff05b23, 32'h400f2f0a} /* (27, 19, 16) {real, imag} */,
  {32'h3fa251ed, 32'h3efc2062} /* (27, 19, 15) {real, imag} */,
  {32'h3f339bb8, 32'h40001416} /* (27, 19, 14) {real, imag} */,
  {32'h3faa6bad, 32'h3faeff5d} /* (27, 19, 13) {real, imag} */,
  {32'h3ff5ca72, 32'h3d5eb330} /* (27, 19, 12) {real, imag} */,
  {32'h3ef4a9f2, 32'h3fc93916} /* (27, 19, 11) {real, imag} */,
  {32'hc02d2ff4, 32'hbe1e77d0} /* (27, 19, 10) {real, imag} */,
  {32'hbf2904d7, 32'hc024ef1a} /* (27, 19, 9) {real, imag} */,
  {32'h3f7bc0e8, 32'hc080257c} /* (27, 19, 8) {real, imag} */,
  {32'h3ee6d872, 32'hc05cf702} /* (27, 19, 7) {real, imag} */,
  {32'hbe387130, 32'hc02ed1ce} /* (27, 19, 6) {real, imag} */,
  {32'hc019b1b2, 32'hc05d4a46} /* (27, 19, 5) {real, imag} */,
  {32'hc00699f0, 32'hc0327d44} /* (27, 19, 4) {real, imag} */,
  {32'hc00f8d08, 32'hbf344ca6} /* (27, 19, 3) {real, imag} */,
  {32'hbf4d258d, 32'hbfd2445f} /* (27, 19, 2) {real, imag} */,
  {32'h3e386d1c, 32'hbfdda522} /* (27, 19, 1) {real, imag} */,
  {32'h3f4de2d8, 32'hbf158f0c} /* (27, 19, 0) {real, imag} */,
  {32'h3fe88a7c, 32'hc00b44a8} /* (27, 18, 31) {real, imag} */,
  {32'h3f796d52, 32'hc06dd126} /* (27, 18, 30) {real, imag} */,
  {32'hbfaf6c12, 32'hbfdce0da} /* (27, 18, 29) {real, imag} */,
  {32'hbf464d60, 32'h3f4ba29a} /* (27, 18, 28) {real, imag} */,
  {32'h3e92acd8, 32'h3ef036fa} /* (27, 18, 27) {real, imag} */,
  {32'hbe8635e4, 32'h3eac63e6} /* (27, 18, 26) {real, imag} */,
  {32'hbf41e133, 32'hbfe44e5d} /* (27, 18, 25) {real, imag} */,
  {32'hc0698f6d, 32'hc0455029} /* (27, 18, 24) {real, imag} */,
  {32'hc059551a, 32'hc076ba20} /* (27, 18, 23) {real, imag} */,
  {32'hbf4bd4f2, 32'hc0820970} /* (27, 18, 22) {real, imag} */,
  {32'hbeac6eeb, 32'hbfbeac36} /* (27, 18, 21) {real, imag} */,
  {32'h40032110, 32'h400dd637} /* (27, 18, 20) {real, imag} */,
  {32'h404eb98c, 32'h4032ad68} /* (27, 18, 19) {real, imag} */,
  {32'h4019e04b, 32'hbf290432} /* (27, 18, 18) {real, imag} */,
  {32'h403dceba, 32'h3fcce1df} /* (27, 18, 17) {real, imag} */,
  {32'h3f707793, 32'h403db9bb} /* (27, 18, 16) {real, imag} */,
  {32'h4016ed38, 32'h3fb51203} /* (27, 18, 15) {real, imag} */,
  {32'h403db41a, 32'h405a29dc} /* (27, 18, 14) {real, imag} */,
  {32'h3fe9d642, 32'h403a1522} /* (27, 18, 13) {real, imag} */,
  {32'h3cfabac0, 32'h3f3341f2} /* (27, 18, 12) {real, imag} */,
  {32'h405e3b33, 32'h3fe0db91} /* (27, 18, 11) {real, imag} */,
  {32'h3fce40ca, 32'h3e18a498} /* (27, 18, 10) {real, imag} */,
  {32'hbf796e74, 32'hc00e9cad} /* (27, 18, 9) {real, imag} */,
  {32'hbfa0d485, 32'hc0044d00} /* (27, 18, 8) {real, imag} */,
  {32'h3f94e65a, 32'hbeae6540} /* (27, 18, 7) {real, imag} */,
  {32'hbe2f1e68, 32'hc0817894} /* (27, 18, 6) {real, imag} */,
  {32'hbf3cbfd6, 32'hc0730970} /* (27, 18, 5) {real, imag} */,
  {32'hbfb02bd0, 32'hc03bbba2} /* (27, 18, 4) {real, imag} */,
  {32'hbf488698, 32'hc02f7dbe} /* (27, 18, 3) {real, imag} */,
  {32'hbe0eb2e8, 32'hbecf281d} /* (27, 18, 2) {real, imag} */,
  {32'hbe7d41b0, 32'hc0404ac0} /* (27, 18, 1) {real, imag} */,
  {32'h4012ac98, 32'hc0057180} /* (27, 18, 0) {real, imag} */,
  {32'hbf446644, 32'hc0465cb0} /* (27, 17, 31) {real, imag} */,
  {32'hbf03de94, 32'hc0cb6b4c} /* (27, 17, 30) {real, imag} */,
  {32'hbf330a48, 32'hc06061d5} /* (27, 17, 29) {real, imag} */,
  {32'h3f8f1b4a, 32'hbeb49618} /* (27, 17, 28) {real, imag} */,
  {32'h405e7b89, 32'hbfd8f43e} /* (27, 17, 27) {real, imag} */,
  {32'h40387b07, 32'hbf03272b} /* (27, 17, 26) {real, imag} */,
  {32'hbf10248c, 32'hc06072ec} /* (27, 17, 25) {real, imag} */,
  {32'hc03fe108, 32'hc0a8b77e} /* (27, 17, 24) {real, imag} */,
  {32'hbfd9bdf4, 32'hc0b297fc} /* (27, 17, 23) {real, imag} */,
  {32'hbf923a3c, 32'hc0311d7e} /* (27, 17, 22) {real, imag} */,
  {32'h3f004ebe, 32'hbf7bf433} /* (27, 17, 21) {real, imag} */,
  {32'h40452bb7, 32'h3f577e59} /* (27, 17, 20) {real, imag} */,
  {32'h4059a834, 32'h3f843a5f} /* (27, 17, 19) {real, imag} */,
  {32'h4032a0c8, 32'hbf9d1bf9} /* (27, 17, 18) {real, imag} */,
  {32'h402ea3dc, 32'h3f098c1c} /* (27, 17, 17) {real, imag} */,
  {32'h400e8728, 32'h3f834455} /* (27, 17, 16) {real, imag} */,
  {32'h4075f217, 32'h3f5334fc} /* (27, 17, 15) {real, imag} */,
  {32'h40592463, 32'h3ef18da8} /* (27, 17, 14) {real, imag} */,
  {32'h402625c5, 32'h3e4018d4} /* (27, 17, 13) {real, imag} */,
  {32'h4018711e, 32'h3f882328} /* (27, 17, 12) {real, imag} */,
  {32'h401d0750, 32'h3ee486da} /* (27, 17, 11) {real, imag} */,
  {32'h3f8dc9aa, 32'hc009aceb} /* (27, 17, 10) {real, imag} */,
  {32'hbfda1290, 32'hc023919c} /* (27, 17, 9) {real, imag} */,
  {32'hbe1c8ef0, 32'hc0445b01} /* (27, 17, 8) {real, imag} */,
  {32'h3f9f7d73, 32'hbfc18fea} /* (27, 17, 7) {real, imag} */,
  {32'h3f97b6d1, 32'hc006126e} /* (27, 17, 6) {real, imag} */,
  {32'hc009e36e, 32'hc02d1cc5} /* (27, 17, 5) {real, imag} */,
  {32'hc03c95e0, 32'hc0186d14} /* (27, 17, 4) {real, imag} */,
  {32'hbf980918, 32'hc0295c2b} /* (27, 17, 3) {real, imag} */,
  {32'h3f437e26, 32'hc01fd304} /* (27, 17, 2) {real, imag} */,
  {32'hbf13ff0c, 32'hc007d9c0} /* (27, 17, 1) {real, imag} */,
  {32'hbec7ada7, 32'hc0033e7e} /* (27, 17, 0) {real, imag} */,
  {32'hbf53f77d, 32'hbf905cdc} /* (27, 16, 31) {real, imag} */,
  {32'h3d86e010, 32'hc08da47a} /* (27, 16, 30) {real, imag} */,
  {32'hbea62352, 32'hc0690f5b} /* (27, 16, 29) {real, imag} */,
  {32'h4057071b, 32'hbff755cd} /* (27, 16, 28) {real, imag} */,
  {32'h403b80fc, 32'hc072ad82} /* (27, 16, 27) {real, imag} */,
  {32'h3ef3df2a, 32'hc01a3369} /* (27, 16, 26) {real, imag} */,
  {32'hbf54f634, 32'hc07eafb1} /* (27, 16, 25) {real, imag} */,
  {32'hbf4db1d2, 32'hc072e79a} /* (27, 16, 24) {real, imag} */,
  {32'hc023e7ec, 32'hc0ba1ad0} /* (27, 16, 23) {real, imag} */,
  {32'hc08ea251, 32'hc08493a2} /* (27, 16, 22) {real, imag} */,
  {32'h3e4ab06c, 32'hbfc08314} /* (27, 16, 21) {real, imag} */,
  {32'h406720cb, 32'hbdc651d0} /* (27, 16, 20) {real, imag} */,
  {32'h406fca26, 32'h3f87d4c8} /* (27, 16, 19) {real, imag} */,
  {32'h40750b28, 32'h400a58ec} /* (27, 16, 18) {real, imag} */,
  {32'h4027d8be, 32'h40582f33} /* (27, 16, 17) {real, imag} */,
  {32'h4015ee10, 32'h40603913} /* (27, 16, 16) {real, imag} */,
  {32'h403b4954, 32'h4029133e} /* (27, 16, 15) {real, imag} */,
  {32'h3fab35ab, 32'hbe8130cc} /* (27, 16, 14) {real, imag} */,
  {32'h40059482, 32'h3f715223} /* (27, 16, 13) {real, imag} */,
  {32'h408c51ca, 32'h406dfdcc} /* (27, 16, 12) {real, imag} */,
  {32'h40223ac0, 32'h403c5606} /* (27, 16, 11) {real, imag} */,
  {32'h400db6ac, 32'h3f6cbcb5} /* (27, 16, 10) {real, imag} */,
  {32'h3f9065c4, 32'hbe979d3c} /* (27, 16, 9) {real, imag} */,
  {32'h40255cae, 32'hc0597a33} /* (27, 16, 8) {real, imag} */,
  {32'h3ff6890a, 32'hc07819f9} /* (27, 16, 7) {real, imag} */,
  {32'h40559ac4, 32'hc021ab18} /* (27, 16, 6) {real, imag} */,
  {32'hbf116cc8, 32'hc01d01b8} /* (27, 16, 5) {real, imag} */,
  {32'hbfd38f38, 32'hc020ae06} /* (27, 16, 4) {real, imag} */,
  {32'hbff0af78, 32'h3d407a40} /* (27, 16, 3) {real, imag} */,
  {32'hc001399a, 32'hbff54de2} /* (27, 16, 2) {real, imag} */,
  {32'hc03cbf06, 32'hbfe9caf9} /* (27, 16, 1) {real, imag} */,
  {32'hc01599e5, 32'hbf038e1b} /* (27, 16, 0) {real, imag} */,
  {32'h3e90d4a0, 32'hbf6686b1} /* (27, 15, 31) {real, imag} */,
  {32'h3f18dafe, 32'hc0050d3b} /* (27, 15, 30) {real, imag} */,
  {32'hc00cc3e6, 32'hc02388d7} /* (27, 15, 29) {real, imag} */,
  {32'hc00c511b, 32'hbff7402e} /* (27, 15, 28) {real, imag} */,
  {32'hc05b390e, 32'hc09a9335} /* (27, 15, 27) {real, imag} */,
  {32'hbfcd4f2e, 32'hc0a1e643} /* (27, 15, 26) {real, imag} */,
  {32'hbfb53348, 32'hc02de67a} /* (27, 15, 25) {real, imag} */,
  {32'h3f2a482d, 32'hc03b8f75} /* (27, 15, 24) {real, imag} */,
  {32'hc053374e, 32'hc0d12b50} /* (27, 15, 23) {real, imag} */,
  {32'hc0a4c4e5, 32'hc0d4f11e} /* (27, 15, 22) {real, imag} */,
  {32'hbf870453, 32'hc0232ecc} /* (27, 15, 21) {real, imag} */,
  {32'h4023209e, 32'hbf56e7aa} /* (27, 15, 20) {real, imag} */,
  {32'h3f482a42, 32'h3f7b340d} /* (27, 15, 19) {real, imag} */,
  {32'hbea3b68e, 32'h405473d9} /* (27, 15, 18) {real, imag} */,
  {32'h3ecfca9b, 32'h408b1283} /* (27, 15, 17) {real, imag} */,
  {32'h3f053c2c, 32'h4088fa60} /* (27, 15, 16) {real, imag} */,
  {32'hbf10526a, 32'h4053386a} /* (27, 15, 15) {real, imag} */,
  {32'hbf90ca0e, 32'h4018f6b0} /* (27, 15, 14) {real, imag} */,
  {32'hbecef88e, 32'h409267a6} /* (27, 15, 13) {real, imag} */,
  {32'h3e3dfa5c, 32'h408be1ab} /* (27, 15, 12) {real, imag} */,
  {32'h3d4cafc0, 32'h4051aeb7} /* (27, 15, 11) {real, imag} */,
  {32'h3d409bc0, 32'hbea94dc4} /* (27, 15, 10) {real, imag} */,
  {32'hbe7c6070, 32'hbfd515b1} /* (27, 15, 9) {real, imag} */,
  {32'h3f8a1fa8, 32'hbfffaf7e} /* (27, 15, 8) {real, imag} */,
  {32'h3f41da06, 32'hc02bbbec} /* (27, 15, 7) {real, imag} */,
  {32'h3faccaaa, 32'hc04917a7} /* (27, 15, 6) {real, imag} */,
  {32'h3fef859e, 32'hbf89d848} /* (27, 15, 5) {real, imag} */,
  {32'hbe6b2dc4, 32'h3f0b332c} /* (27, 15, 4) {real, imag} */,
  {32'hc02e6464, 32'h3edc6ea0} /* (27, 15, 3) {real, imag} */,
  {32'hc072b1c9, 32'hbf56cf68} /* (27, 15, 2) {real, imag} */,
  {32'hc088c7fe, 32'hbfe6b1cb} /* (27, 15, 1) {real, imag} */,
  {32'hc04bb62c, 32'hbfccaf35} /* (27, 15, 0) {real, imag} */,
  {32'hbf657fe2, 32'hbee28506} /* (27, 14, 31) {real, imag} */,
  {32'hbf409042, 32'h3f8bff6c} /* (27, 14, 30) {real, imag} */,
  {32'hbffccc18, 32'hbf85fd66} /* (27, 14, 29) {real, imag} */,
  {32'hc014f7a0, 32'hc0707842} /* (27, 14, 28) {real, imag} */,
  {32'hc0498304, 32'hc086dc13} /* (27, 14, 27) {real, imag} */,
  {32'hbfa4f4f1, 32'hbfea5e8d} /* (27, 14, 26) {real, imag} */,
  {32'hbe576e20, 32'hbfb0f818} /* (27, 14, 25) {real, imag} */,
  {32'h3ea315ae, 32'hbff84344} /* (27, 14, 24) {real, imag} */,
  {32'hc07ed662, 32'hc0998f6a} /* (27, 14, 23) {real, imag} */,
  {32'hc086026c, 32'hc09d3e6c} /* (27, 14, 22) {real, imag} */,
  {32'hbed32604, 32'hbfc5e22e} /* (27, 14, 21) {real, imag} */,
  {32'h3fb24982, 32'h3ec63c70} /* (27, 14, 20) {real, imag} */,
  {32'h3f810e03, 32'h40312a82} /* (27, 14, 19) {real, imag} */,
  {32'hbf4358be, 32'h405e69fb} /* (27, 14, 18) {real, imag} */,
  {32'hbff7c78e, 32'h4065c2ce} /* (27, 14, 17) {real, imag} */,
  {32'hbe90f1a6, 32'h402c5b10} /* (27, 14, 16) {real, imag} */,
  {32'hbf06b22f, 32'h3fc59d6a} /* (27, 14, 15) {real, imag} */,
  {32'hc01a4480, 32'h3ff7ac9a} /* (27, 14, 14) {real, imag} */,
  {32'hbfe4a077, 32'h407d9c84} /* (27, 14, 13) {real, imag} */,
  {32'hbf5c8970, 32'h3f999af9} /* (27, 14, 12) {real, imag} */,
  {32'hbfa346f1, 32'h3f23be34} /* (27, 14, 11) {real, imag} */,
  {32'hc082f4df, 32'hbe4d236c} /* (27, 14, 10) {real, imag} */,
  {32'hc001dfa6, 32'hc0225830} /* (27, 14, 9) {real, imag} */,
  {32'hbf8ac0cd, 32'hbfdb4ab2} /* (27, 14, 8) {real, imag} */,
  {32'hc0632cb0, 32'hc013cc22} /* (27, 14, 7) {real, imag} */,
  {32'hbfe9d608, 32'hbfa2217a} /* (27, 14, 6) {real, imag} */,
  {32'h3ea7d384, 32'h3f0213d0} /* (27, 14, 5) {real, imag} */,
  {32'hbfc3f4aa, 32'hbf25a1d7} /* (27, 14, 4) {real, imag} */,
  {32'hbfdc4cd5, 32'hbf2aeb74} /* (27, 14, 3) {real, imag} */,
  {32'hc031a250, 32'hbe2559dc} /* (27, 14, 2) {real, imag} */,
  {32'hc084228f, 32'hbfbcf976} /* (27, 14, 1) {real, imag} */,
  {32'hc05ea6ad, 32'hbf3c7d7d} /* (27, 14, 0) {real, imag} */,
  {32'hbf9a4d9b, 32'hbc7cbce0} /* (27, 13, 31) {real, imag} */,
  {32'hc01e0336, 32'h3f891e5a} /* (27, 13, 30) {real, imag} */,
  {32'hc05aabe4, 32'hbee63f98} /* (27, 13, 29) {real, imag} */,
  {32'hbfb97817, 32'hc0248ca0} /* (27, 13, 28) {real, imag} */,
  {32'hbf1902a8, 32'hbfc9db73} /* (27, 13, 27) {real, imag} */,
  {32'hbf23fb22, 32'h3eb3f918} /* (27, 13, 26) {real, imag} */,
  {32'hbee57b84, 32'h3e270410} /* (27, 13, 25) {real, imag} */,
  {32'hbfeb6cc6, 32'h3e88c408} /* (27, 13, 24) {real, imag} */,
  {32'hc0210c00, 32'hbee2c3a0} /* (27, 13, 23) {real, imag} */,
  {32'hc0707a3e, 32'hbf698f56} /* (27, 13, 22) {real, imag} */,
  {32'hbfc23e05, 32'hbfd99f2a} /* (27, 13, 21) {real, imag} */,
  {32'h3efc557c, 32'h3fefe0be} /* (27, 13, 20) {real, imag} */,
  {32'h3fda560f, 32'h40079492} /* (27, 13, 19) {real, imag} */,
  {32'h3f80d20b, 32'h404a245c} /* (27, 13, 18) {real, imag} */,
  {32'h3d8822c0, 32'h403ec888} /* (27, 13, 17) {real, imag} */,
  {32'hbfa1664a, 32'h3f6d09f0} /* (27, 13, 16) {real, imag} */,
  {32'hbf427134, 32'h3fa2e816} /* (27, 13, 15) {real, imag} */,
  {32'hbfa5526f, 32'h3fbea2b1} /* (27, 13, 14) {real, imag} */,
  {32'hbfc25eac, 32'h4009a635} /* (27, 13, 13) {real, imag} */,
  {32'hbf30a732, 32'h3f9cdb18} /* (27, 13, 12) {real, imag} */,
  {32'h3e9f50d2, 32'hbef35bc0} /* (27, 13, 11) {real, imag} */,
  {32'hc0126ece, 32'hc00e2688} /* (27, 13, 10) {real, imag} */,
  {32'hc02f00aa, 32'hc020652e} /* (27, 13, 9) {real, imag} */,
  {32'hbf53a7bc, 32'hbd194a10} /* (27, 13, 8) {real, imag} */,
  {32'hc05b3a57, 32'hc0144e05} /* (27, 13, 7) {real, imag} */,
  {32'hc0176532, 32'hc0083495} /* (27, 13, 6) {real, imag} */,
  {32'hbe04c35e, 32'hbecc6840} /* (27, 13, 5) {real, imag} */,
  {32'hbf455ed5, 32'hbf6bed12} /* (27, 13, 4) {real, imag} */,
  {32'hbfd9f92c, 32'hc0077a71} /* (27, 13, 3) {real, imag} */,
  {32'hc0352ffa, 32'hbfbd4e08} /* (27, 13, 2) {real, imag} */,
  {32'hc05a6a38, 32'hbece06e4} /* (27, 13, 1) {real, imag} */,
  {32'hbf6dd414, 32'hbf0fab08} /* (27, 13, 0) {real, imag} */,
  {32'hbf5ca718, 32'h3cf85c60} /* (27, 12, 31) {real, imag} */,
  {32'hbfaecb5e, 32'hc0011c2c} /* (27, 12, 30) {real, imag} */,
  {32'hc09b5b24, 32'hc05c64d9} /* (27, 12, 29) {real, imag} */,
  {32'hc077e169, 32'hc07fd708} /* (27, 12, 28) {real, imag} */,
  {32'hbf35fb86, 32'hc003e6a6} /* (27, 12, 27) {real, imag} */,
  {32'hbf77a4ce, 32'hc04d256e} /* (27, 12, 26) {real, imag} */,
  {32'hc0325b6c, 32'hc07cb926} /* (27, 12, 25) {real, imag} */,
  {32'hc07fa9f3, 32'h3e333b24} /* (27, 12, 24) {real, imag} */,
  {32'hc007bcc2, 32'h4023f987} /* (27, 12, 23) {real, imag} */,
  {32'hbfdd7493, 32'h3f315fca} /* (27, 12, 22) {real, imag} */,
  {32'h3f65c185, 32'h3f89f2d5} /* (27, 12, 21) {real, imag} */,
  {32'h3f85d2d0, 32'h40494517} /* (27, 12, 20) {real, imag} */,
  {32'h3f07f3c2, 32'h40657be0} /* (27, 12, 19) {real, imag} */,
  {32'h3fc20064, 32'h402550e6} /* (27, 12, 18) {real, imag} */,
  {32'h3ecdf280, 32'h4031a804} /* (27, 12, 17) {real, imag} */,
  {32'hbe885e2f, 32'h3f5ffd18} /* (27, 12, 16) {real, imag} */,
  {32'h3fa9afd8, 32'h400fc2a0} /* (27, 12, 15) {real, imag} */,
  {32'hbf62b597, 32'h3e845612} /* (27, 12, 14) {real, imag} */,
  {32'hbf56c4a9, 32'h3fa18e78} /* (27, 12, 13) {real, imag} */,
  {32'h4007f2cc, 32'h3feabd96} /* (27, 12, 12) {real, imag} */,
  {32'h3fc8f960, 32'h4026b8d2} /* (27, 12, 11) {real, imag} */,
  {32'hbf3d9ea4, 32'hbfc4002c} /* (27, 12, 10) {real, imag} */,
  {32'hbfc424e5, 32'hc01f0bb9} /* (27, 12, 9) {real, imag} */,
  {32'hbf86498d, 32'hbf8f24cc} /* (27, 12, 8) {real, imag} */,
  {32'hbfe93eb3, 32'hbfdafba3} /* (27, 12, 7) {real, imag} */,
  {32'hc07253ff, 32'hbfdb3cfd} /* (27, 12, 6) {real, imag} */,
  {32'hc00fadc6, 32'hbebb955a} /* (27, 12, 5) {real, imag} */,
  {32'hbf6854d0, 32'h3cabce60} /* (27, 12, 4) {real, imag} */,
  {32'hbfea8ac6, 32'hc01ef62c} /* (27, 12, 3) {real, imag} */,
  {32'hc01e4354, 32'hc0351a5e} /* (27, 12, 2) {real, imag} */,
  {32'hc0183a94, 32'hc00aceb9} /* (27, 12, 1) {real, imag} */,
  {32'hbe8c0139, 32'hbf62d5f7} /* (27, 12, 0) {real, imag} */,
  {32'h3e2a4df8, 32'h3fb14ce4} /* (27, 11, 31) {real, imag} */,
  {32'hbf8178f4, 32'hbe2c6b60} /* (27, 11, 30) {real, imag} */,
  {32'hc0620fc2, 32'hbfd4309f} /* (27, 11, 29) {real, imag} */,
  {32'hc02b2d63, 32'hc05ec191} /* (27, 11, 28) {real, imag} */,
  {32'hbf7d8d83, 32'hbfd4325c} /* (27, 11, 27) {real, imag} */,
  {32'hbfe1123f, 32'hc071f1b5} /* (27, 11, 26) {real, imag} */,
  {32'hbf9d7efa, 32'hc073d0a4} /* (27, 11, 25) {real, imag} */,
  {32'hbf26f034, 32'hbf32e83a} /* (27, 11, 24) {real, imag} */,
  {32'hbca33c00, 32'hbf8bf648} /* (27, 11, 23) {real, imag} */,
  {32'h3ea488d1, 32'hbfab6a0c} /* (27, 11, 22) {real, imag} */,
  {32'h3f94d79c, 32'h3dbdf9e8} /* (27, 11, 21) {real, imag} */,
  {32'h400805e8, 32'h3f675a99} /* (27, 11, 20) {real, imag} */,
  {32'h3f943084, 32'h3fddaa43} /* (27, 11, 19) {real, imag} */,
  {32'hbe1795ca, 32'h40008b3a} /* (27, 11, 18) {real, imag} */,
  {32'hbf159bea, 32'h40070207} /* (27, 11, 17) {real, imag} */,
  {32'h3f7a05be, 32'hbf211bb9} /* (27, 11, 16) {real, imag} */,
  {32'h3faf0478, 32'h3f63ec98} /* (27, 11, 15) {real, imag} */,
  {32'hbf568694, 32'h3f09d171} /* (27, 11, 14) {real, imag} */,
  {32'hbeddf32c, 32'h402451d5} /* (27, 11, 13) {real, imag} */,
  {32'h404a1a9c, 32'h3f186d7a} /* (27, 11, 12) {real, imag} */,
  {32'h4012ed98, 32'h3e1cfd38} /* (27, 11, 11) {real, imag} */,
  {32'hbfa0cced, 32'hbfa041ea} /* (27, 11, 10) {real, imag} */,
  {32'hc0915c95, 32'hbf2bee3d} /* (27, 11, 9) {real, imag} */,
  {32'hc06a6ed8, 32'hbf079964} /* (27, 11, 8) {real, imag} */,
  {32'hbf4aef1a, 32'hbfb5c122} /* (27, 11, 7) {real, imag} */,
  {32'hc0686e7b, 32'hbfc3e3c3} /* (27, 11, 6) {real, imag} */,
  {32'hc0a3df53, 32'hbf86813e} /* (27, 11, 5) {real, imag} */,
  {32'hc05f7946, 32'h3fdf17e4} /* (27, 11, 4) {real, imag} */,
  {32'hbfb4a5ad, 32'h3fdabaed} /* (27, 11, 3) {real, imag} */,
  {32'h3e362754, 32'hc0168150} /* (27, 11, 2) {real, imag} */,
  {32'hbfa83912, 32'hc09e8267} /* (27, 11, 1) {real, imag} */,
  {32'hbfa5cc70, 32'hbfb60756} /* (27, 11, 0) {real, imag} */,
  {32'h3fff1d42, 32'h3fc3c34a} /* (27, 10, 31) {real, imag} */,
  {32'h3fb352a7, 32'h400685ce} /* (27, 10, 30) {real, imag} */,
  {32'hbf363150, 32'h407bf4ba} /* (27, 10, 29) {real, imag} */,
  {32'h3eab7364, 32'h3feaff6e} /* (27, 10, 28) {real, imag} */,
  {32'hbf5f86c0, 32'h3f74be41} /* (27, 10, 27) {real, imag} */,
  {32'hbf95f683, 32'hbed323dd} /* (27, 10, 26) {real, imag} */,
  {32'hbfb7bd86, 32'hbeee0d30} /* (27, 10, 25) {real, imag} */,
  {32'h3eb05932, 32'h3fc3ecca} /* (27, 10, 24) {real, imag} */,
  {32'h3f4cc386, 32'h3f9fa0ea} /* (27, 10, 23) {real, imag} */,
  {32'hbf884e50, 32'h3ffdf89a} /* (27, 10, 22) {real, imag} */,
  {32'h38390000, 32'h3fcf814c} /* (27, 10, 21) {real, imag} */,
  {32'h3f846a13, 32'hbe818338} /* (27, 10, 20) {real, imag} */,
  {32'h3f41ef02, 32'hbff77068} /* (27, 10, 19) {real, imag} */,
  {32'hbf2ba190, 32'hbf9b5b86} /* (27, 10, 18) {real, imag} */,
  {32'hbf3f1bbf, 32'hc00e30ba} /* (27, 10, 17) {real, imag} */,
  {32'hbf6a34da, 32'hc023a703} /* (27, 10, 16) {real, imag} */,
  {32'hbe81f0c2, 32'hc0246ac6} /* (27, 10, 15) {real, imag} */,
  {32'h3dc98654, 32'hbfef8038} /* (27, 10, 14) {real, imag} */,
  {32'hbf7fd2e2, 32'hbf14f2da} /* (27, 10, 13) {real, imag} */,
  {32'hbe5e2ba5, 32'hc04702d8} /* (27, 10, 12) {real, imag} */,
  {32'hc0169799, 32'hc08b1fe6} /* (27, 10, 11) {real, imag} */,
  {32'hbf653144, 32'h3f0f24ac} /* (27, 10, 10) {real, imag} */,
  {32'hc0183e08, 32'h3f8db5d2} /* (27, 10, 9) {real, imag} */,
  {32'hbf2acced, 32'h3fb46482} /* (27, 10, 8) {real, imag} */,
  {32'h3f91c5b8, 32'h3edef88c} /* (27, 10, 7) {real, imag} */,
  {32'hbfdd1f58, 32'h3f76bc62} /* (27, 10, 6) {real, imag} */,
  {32'hc040bd78, 32'h3dff65c0} /* (27, 10, 5) {real, imag} */,
  {32'hbed8cda8, 32'h40004d32} /* (27, 10, 4) {real, imag} */,
  {32'h3fb03af4, 32'h40628870} /* (27, 10, 3) {real, imag} */,
  {32'h3f89f141, 32'h3fdfff96} /* (27, 10, 2) {real, imag} */,
  {32'h3f4ee5f0, 32'h3dec6528} /* (27, 10, 1) {real, imag} */,
  {32'h3eb82210, 32'h3fc0e50c} /* (27, 10, 0) {real, imag} */,
  {32'h3fd6917e, 32'h3fba1e0c} /* (27, 9, 31) {real, imag} */,
  {32'h40385302, 32'h4033cd8c} /* (27, 9, 30) {real, imag} */,
  {32'hbf1fdc26, 32'h408ef262} /* (27, 9, 29) {real, imag} */,
  {32'hbfd3c30a, 32'h40656c52} /* (27, 9, 28) {real, imag} */,
  {32'hbe36a130, 32'h40307e18} /* (27, 9, 27) {real, imag} */,
  {32'h3ed064ea, 32'h3fbfc08e} /* (27, 9, 26) {real, imag} */,
  {32'h3e260864, 32'h400f08f5} /* (27, 9, 25) {real, imag} */,
  {32'h3fd7d0af, 32'h4089fc4e} /* (27, 9, 24) {real, imag} */,
  {32'h3fcccbed, 32'h3f7ac47c} /* (27, 9, 23) {real, imag} */,
  {32'h3ff77d28, 32'h40090ba4} /* (27, 9, 22) {real, imag} */,
  {32'h40263963, 32'h3ff990dc} /* (27, 9, 21) {real, imag} */,
  {32'h3db09e60, 32'hbe9ceb20} /* (27, 9, 20) {real, imag} */,
  {32'hbf452f04, 32'hbffdffca} /* (27, 9, 19) {real, imag} */,
  {32'hbfd2b4e7, 32'hc0bc5480} /* (27, 9, 18) {real, imag} */,
  {32'hc01b3299, 32'hc0ade52e} /* (27, 9, 17) {real, imag} */,
  {32'hc019138e, 32'hc03b3ac6} /* (27, 9, 16) {real, imag} */,
  {32'h3eaac192, 32'hc083f90d} /* (27, 9, 15) {real, imag} */,
  {32'hbf08fc20, 32'hc0720c08} /* (27, 9, 14) {real, imag} */,
  {32'hc0340618, 32'hc09e98ea} /* (27, 9, 13) {real, imag} */,
  {32'hbf836a70, 32'hc0402102} /* (27, 9, 12) {real, imag} */,
  {32'hbf31bf9a, 32'hbf5ce314} /* (27, 9, 11) {real, imag} */,
  {32'hbe2d0710, 32'h400b3088} /* (27, 9, 10) {real, imag} */,
  {32'hbe1c5d64, 32'h401032df} /* (27, 9, 9) {real, imag} */,
  {32'h407a7cec, 32'h400105ca} /* (27, 9, 8) {real, imag} */,
  {32'h40477198, 32'h3d470ee0} /* (27, 9, 7) {real, imag} */,
  {32'h3e14dddc, 32'h3fd4e5e6} /* (27, 9, 6) {real, imag} */,
  {32'h3e9eadaa, 32'h401ca331} /* (27, 9, 5) {real, imag} */,
  {32'h3ef0c3dc, 32'h3fd51801} /* (27, 9, 4) {real, imag} */,
  {32'h3f9593b3, 32'h3fba09d1} /* (27, 9, 3) {real, imag} */,
  {32'h402960e6, 32'h4034e680} /* (27, 9, 2) {real, imag} */,
  {32'h40063670, 32'h405967c0} /* (27, 9, 1) {real, imag} */,
  {32'h3e4d3d20, 32'h402a7c15} /* (27, 9, 0) {real, imag} */,
  {32'h3fbe5ebb, 32'h3fe15aef} /* (27, 8, 31) {real, imag} */,
  {32'h40125754, 32'h3fed7b18} /* (27, 8, 30) {real, imag} */,
  {32'hc0384e8f, 32'h40795c30} /* (27, 8, 29) {real, imag} */,
  {32'hbf0f9fdd, 32'h4079746d} /* (27, 8, 28) {real, imag} */,
  {32'h3e229b78, 32'h40167e07} /* (27, 8, 27) {real, imag} */,
  {32'h3f08f944, 32'h3fded139} /* (27, 8, 26) {real, imag} */,
  {32'h3e58dc97, 32'h403288f7} /* (27, 8, 25) {real, imag} */,
  {32'h40371e84, 32'h40122ecb} /* (27, 8, 24) {real, imag} */,
  {32'h3fef3067, 32'hbe39aaf0} /* (27, 8, 23) {real, imag} */,
  {32'hbaee0c00, 32'h4028240a} /* (27, 8, 22) {real, imag} */,
  {32'hbf50fc2a, 32'hbe7dd6e0} /* (27, 8, 21) {real, imag} */,
  {32'hbf60e8b5, 32'hbf826c56} /* (27, 8, 20) {real, imag} */,
  {32'hc004a49e, 32'hbf990010} /* (27, 8, 19) {real, imag} */,
  {32'hc002da67, 32'hc0a25daa} /* (27, 8, 18) {real, imag} */,
  {32'hc01f4fb8, 32'hc05ee326} /* (27, 8, 17) {real, imag} */,
  {32'hc0667012, 32'hc066fa2a} /* (27, 8, 16) {real, imag} */,
  {32'hbfdd6a8a, 32'hc061c06e} /* (27, 8, 15) {real, imag} */,
  {32'h3eacf902, 32'hbf11fda2} /* (27, 8, 14) {real, imag} */,
  {32'hbf6b9dba, 32'hc0837c86} /* (27, 8, 13) {real, imag} */,
  {32'hbff05e1d, 32'hc073b0bf} /* (27, 8, 12) {real, imag} */,
  {32'h3f66b7dc, 32'hc0352d39} /* (27, 8, 11) {real, imag} */,
  {32'h3fc2595a, 32'h3f699778} /* (27, 8, 10) {real, imag} */,
  {32'h4020e12c, 32'h3feda017} /* (27, 8, 9) {real, imag} */,
  {32'h409720b0, 32'h40328cf0} /* (27, 8, 8) {real, imag} */,
  {32'h4024cd42, 32'h40473ee2} /* (27, 8, 7) {real, imag} */,
  {32'hbe3c0fa4, 32'h40b84690} /* (27, 8, 6) {real, imag} */,
  {32'h400171ac, 32'h40a5a14a} /* (27, 8, 5) {real, imag} */,
  {32'h40005d37, 32'h40126cc4} /* (27, 8, 4) {real, imag} */,
  {32'h3fd1f30d, 32'h3f4db8f4} /* (27, 8, 3) {real, imag} */,
  {32'h3fa4c52c, 32'h3feb5dfc} /* (27, 8, 2) {real, imag} */,
  {32'h3e7bc294, 32'h4022bc0c} /* (27, 8, 1) {real, imag} */,
  {32'hbee21331, 32'h402ee007} /* (27, 8, 0) {real, imag} */,
  {32'h3f71460a, 32'h3f2d94d8} /* (27, 7, 31) {real, imag} */,
  {32'h3fa9b1a4, 32'h400e12b6} /* (27, 7, 30) {real, imag} */,
  {32'hc048988b, 32'h400c80be} /* (27, 7, 29) {real, imag} */,
  {32'hbf8d46ce, 32'h3ff1a5f8} /* (27, 7, 28) {real, imag} */,
  {32'h3fcd3620, 32'h3fd8dba7} /* (27, 7, 27) {real, imag} */,
  {32'h400b8532, 32'h3f7219d6} /* (27, 7, 26) {real, imag} */,
  {32'hbed910c8, 32'h403b3b0c} /* (27, 7, 25) {real, imag} */,
  {32'h3f1a9f26, 32'h4067830d} /* (27, 7, 24) {real, imag} */,
  {32'h401a2e0c, 32'h403400bc} /* (27, 7, 23) {real, imag} */,
  {32'h3fc51d8b, 32'h4045f23a} /* (27, 7, 22) {real, imag} */,
  {32'hc00c30dc, 32'h3f571c4d} /* (27, 7, 21) {real, imag} */,
  {32'hc0090901, 32'hc0109917} /* (27, 7, 20) {real, imag} */,
  {32'hbcb7f000, 32'hc06684d0} /* (27, 7, 19) {real, imag} */,
  {32'hbf062611, 32'hc0966009} /* (27, 7, 18) {real, imag} */,
  {32'hc04fe8c1, 32'hc0a7e684} /* (27, 7, 17) {real, imag} */,
  {32'hc03d4d73, 32'hc0264d18} /* (27, 7, 16) {real, imag} */,
  {32'hbf8710f8, 32'hbf988b5c} /* (27, 7, 15) {real, imag} */,
  {32'hbf98656f, 32'h3eefb5d4} /* (27, 7, 14) {real, imag} */,
  {32'hbfe8b1e6, 32'hc0207fd0} /* (27, 7, 13) {real, imag} */,
  {32'hbfc125b7, 32'hc013189b} /* (27, 7, 12) {real, imag} */,
  {32'hc0457f56, 32'hc0889118} /* (27, 7, 11) {real, imag} */,
  {32'h3f6910fc, 32'h3f1d8fa4} /* (27, 7, 10) {real, imag} */,
  {32'h400c9a66, 32'h404c4748} /* (27, 7, 9) {real, imag} */,
  {32'h3fce6f04, 32'h4091f98a} /* (27, 7, 8) {real, imag} */,
  {32'h3eba6e73, 32'h3fa94294} /* (27, 7, 7) {real, imag} */,
  {32'h3f7c0ee5, 32'h4043d01d} /* (27, 7, 6) {real, imag} */,
  {32'h3e982430, 32'h405140ca} /* (27, 7, 5) {real, imag} */,
  {32'h3fe8c095, 32'h3fbe9a43} /* (27, 7, 4) {real, imag} */,
  {32'h401f7eff, 32'hbfacacc9} /* (27, 7, 3) {real, imag} */,
  {32'h3ec43580, 32'hbfde82aa} /* (27, 7, 2) {real, imag} */,
  {32'hbf92bef4, 32'h3fd8e47c} /* (27, 7, 1) {real, imag} */,
  {32'hbd057ae0, 32'h401e2092} /* (27, 7, 0) {real, imag} */,
  {32'hbe4da3d6, 32'hbcb2fbb0} /* (27, 6, 31) {real, imag} */,
  {32'h3f0f9c30, 32'h4006c30f} /* (27, 6, 30) {real, imag} */,
  {32'h3f8b3142, 32'h407a41a2} /* (27, 6, 29) {real, imag} */,
  {32'h3fa4c70a, 32'h3fa20c29} /* (27, 6, 28) {real, imag} */,
  {32'h407f0e84, 32'h3e8a958c} /* (27, 6, 27) {real, imag} */,
  {32'h40398812, 32'h400f0a67} /* (27, 6, 26) {real, imag} */,
  {32'h3fb64a27, 32'h405217c0} /* (27, 6, 25) {real, imag} */,
  {32'hbf1cf722, 32'h404afc71} /* (27, 6, 24) {real, imag} */,
  {32'h3e14e8dc, 32'h40748d60} /* (27, 6, 23) {real, imag} */,
  {32'h3fd7adfc, 32'h408dd33b} /* (27, 6, 22) {real, imag} */,
  {32'hbef58e78, 32'h404af78c} /* (27, 6, 21) {real, imag} */,
  {32'hc004aef2, 32'h3ef34cda} /* (27, 6, 20) {real, imag} */,
  {32'hbf93629e, 32'hc04ac6e8} /* (27, 6, 19) {real, imag} */,
  {32'hbf1cf8b6, 32'hc050dc91} /* (27, 6, 18) {real, imag} */,
  {32'hc02867b1, 32'hc01c8c4b} /* (27, 6, 17) {real, imag} */,
  {32'hbf959bdc, 32'hbd9376c0} /* (27, 6, 16) {real, imag} */,
  {32'h3e829736, 32'hbf49112f} /* (27, 6, 15) {real, imag} */,
  {32'hbea56f96, 32'hc00a7da4} /* (27, 6, 14) {real, imag} */,
  {32'hc0094f1b, 32'hc04b3b10} /* (27, 6, 13) {real, imag} */,
  {32'hbdb42508, 32'hbf9fc3bd} /* (27, 6, 12) {real, imag} */,
  {32'hc02723d8, 32'hbf99942d} /* (27, 6, 11) {real, imag} */,
  {32'hbdc371f8, 32'h3f120737} /* (27, 6, 10) {real, imag} */,
  {32'h400cedca, 32'h3fbe9bb7} /* (27, 6, 9) {real, imag} */,
  {32'h40461ec9, 32'h3fa5b1e1} /* (27, 6, 8) {real, imag} */,
  {32'h3fb8499b, 32'hbe02d7b8} /* (27, 6, 7) {real, imag} */,
  {32'h4025067e, 32'h3fcbdc64} /* (27, 6, 6) {real, imag} */,
  {32'hbf85d34e, 32'h404ddd92} /* (27, 6, 5) {real, imag} */,
  {32'hbe91231e, 32'h4085a002} /* (27, 6, 4) {real, imag} */,
  {32'h3f2d27ee, 32'h3fd3f724} /* (27, 6, 3) {real, imag} */,
  {32'h401c033a, 32'h3fa433e4} /* (27, 6, 2) {real, imag} */,
  {32'h400a72dd, 32'h404dba13} /* (27, 6, 1) {real, imag} */,
  {32'h3f8da5f8, 32'h4000f5ca} /* (27, 6, 0) {real, imag} */,
  {32'h3ed1455e, 32'hbcc34ea0} /* (27, 5, 31) {real, imag} */,
  {32'hbda8a308, 32'h3f93038a} /* (27, 5, 30) {real, imag} */,
  {32'h3fd636d9, 32'h406bdaa4} /* (27, 5, 29) {real, imag} */,
  {32'h3fef4fb3, 32'h407f27d4} /* (27, 5, 28) {real, imag} */,
  {32'h403c7e11, 32'h3f965e66} /* (27, 5, 27) {real, imag} */,
  {32'h401b1563, 32'h3c290ec0} /* (27, 5, 26) {real, imag} */,
  {32'h400274f8, 32'h40573922} /* (27, 5, 25) {real, imag} */,
  {32'h3eb169b4, 32'h40650529} /* (27, 5, 24) {real, imag} */,
  {32'hbeb9eb18, 32'h40060b54} /* (27, 5, 23) {real, imag} */,
  {32'hbea45154, 32'h408b28fc} /* (27, 5, 22) {real, imag} */,
  {32'h3f408ea0, 32'h4093a6d2} /* (27, 5, 21) {real, imag} */,
  {32'hbf1418be, 32'h409d5e26} /* (27, 5, 20) {real, imag} */,
  {32'hbf9142ae, 32'h40044c1e} /* (27, 5, 19) {real, imag} */,
  {32'hbf7adb04, 32'h3ce434e0} /* (27, 5, 18) {real, imag} */,
  {32'hbe993f11, 32'h3f416d15} /* (27, 5, 17) {real, imag} */,
  {32'h3fc1f95c, 32'hbf4455b8} /* (27, 5, 16) {real, imag} */,
  {32'hbfa53e68, 32'hbfed65ba} /* (27, 5, 15) {real, imag} */,
  {32'hc089f20c, 32'hc0762eed} /* (27, 5, 14) {real, imag} */,
  {32'hc044637a, 32'hc006c9d0} /* (27, 5, 13) {real, imag} */,
  {32'h3e2262a0, 32'hbf1b2fec} /* (27, 5, 12) {real, imag} */,
  {32'h3f4488f5, 32'h3f42766c} /* (27, 5, 11) {real, imag} */,
  {32'hbf8bfe4a, 32'hbfb8ec45} /* (27, 5, 10) {real, imag} */,
  {32'hbf758334, 32'hbf3be7be} /* (27, 5, 9) {real, imag} */,
  {32'hbff93f81, 32'hbf7765e6} /* (27, 5, 8) {real, imag} */,
  {32'hc00a282a, 32'hbf224ce5} /* (27, 5, 7) {real, imag} */,
  {32'hbfe9cac6, 32'h3ee7bb7e} /* (27, 5, 6) {real, imag} */,
  {32'hc00c9a2e, 32'h40588c3f} /* (27, 5, 5) {real, imag} */,
  {32'hbeef24ca, 32'h400c9977} /* (27, 5, 4) {real, imag} */,
  {32'h3f3a3f3e, 32'h3f283d62} /* (27, 5, 3) {real, imag} */,
  {32'h3f7f6148, 32'h3fe36d9e} /* (27, 5, 2) {real, imag} */,
  {32'h3d47df10, 32'h4054d7a4} /* (27, 5, 1) {real, imag} */,
  {32'h3f2033ad, 32'h401d060c} /* (27, 5, 0) {real, imag} */,
  {32'h3f18c680, 32'h3f4a1d45} /* (27, 4, 31) {real, imag} */,
  {32'h4022e5f8, 32'h40219400} /* (27, 4, 30) {real, imag} */,
  {32'h3fc52fcb, 32'h4066772f} /* (27, 4, 29) {real, imag} */,
  {32'h3f0a3f3e, 32'h4093ba69} /* (27, 4, 28) {real, imag} */,
  {32'h3f98b6e2, 32'h3faa5788} /* (27, 4, 27) {real, imag} */,
  {32'h40298ee1, 32'hc0434833} /* (27, 4, 26) {real, imag} */,
  {32'h4036a730, 32'hbff96190} /* (27, 4, 25) {real, imag} */,
  {32'h3f43d3e7, 32'h401c5be8} /* (27, 4, 24) {real, imag} */,
  {32'h3fac1bf6, 32'h406865f1} /* (27, 4, 23) {real, imag} */,
  {32'h3fc202c0, 32'h40a11ebb} /* (27, 4, 22) {real, imag} */,
  {32'h400bb3c2, 32'h40affbfc} /* (27, 4, 21) {real, imag} */,
  {32'h3fdbd92d, 32'h402d8bac} /* (27, 4, 20) {real, imag} */,
  {32'hbebd045d, 32'h3fdafaa4} /* (27, 4, 19) {real, imag} */,
  {32'h3ed4b624, 32'h4008c4f2} /* (27, 4, 18) {real, imag} */,
  {32'h3f132a63, 32'h40107b40} /* (27, 4, 17) {real, imag} */,
  {32'h400b4958, 32'h3f01fe40} /* (27, 4, 16) {real, imag} */,
  {32'hbf4d1a18, 32'hbec99c56} /* (27, 4, 15) {real, imag} */,
  {32'hc097baa9, 32'hbf604f30} /* (27, 4, 14) {real, imag} */,
  {32'hc055cd6c, 32'hbfc91f68} /* (27, 4, 13) {real, imag} */,
  {32'hbf9ce882, 32'hbfb77687} /* (27, 4, 12) {real, imag} */,
  {32'h3efdd552, 32'h3d21bcf0} /* (27, 4, 11) {real, imag} */,
  {32'hc01addae, 32'h3f0b14c8} /* (27, 4, 10) {real, imag} */,
  {32'hc0612674, 32'hbfb52539} /* (27, 4, 9) {real, imag} */,
  {32'hc04ac067, 32'hbfca405d} /* (27, 4, 8) {real, imag} */,
  {32'hbff152a2, 32'hbed18e0e} /* (27, 4, 7) {real, imag} */,
  {32'hc0700ab3, 32'hbfa43262} /* (27, 4, 6) {real, imag} */,
  {32'hc0193114, 32'h402a7e14} /* (27, 4, 5) {real, imag} */,
  {32'h3f679882, 32'h4098e85e} /* (27, 4, 4) {real, imag} */,
  {32'h3ff75ee3, 32'h404a812b} /* (27, 4, 3) {real, imag} */,
  {32'h3f9d9032, 32'h3fb14c3c} /* (27, 4, 2) {real, imag} */,
  {32'h3fc9a178, 32'h3ed27ff1} /* (27, 4, 1) {real, imag} */,
  {32'h3fa46c53, 32'h3e7a8e7e} /* (27, 4, 0) {real, imag} */,
  {32'h3ff9e249, 32'h3fa8f971} /* (27, 3, 31) {real, imag} */,
  {32'h40a7d4dc, 32'h3fc1657f} /* (27, 3, 30) {real, imag} */,
  {32'h4032a0cd, 32'h3f915aa4} /* (27, 3, 29) {real, imag} */,
  {32'h3fd33b48, 32'h406c610e} /* (27, 3, 28) {real, imag} */,
  {32'h4004a288, 32'h4040b55f} /* (27, 3, 27) {real, imag} */,
  {32'h3ff872cb, 32'h3e6a4d90} /* (27, 3, 26) {real, imag} */,
  {32'h4042fc02, 32'hbfd76853} /* (27, 3, 25) {real, imag} */,
  {32'h3fd53ea8, 32'h3f8ff66b} /* (27, 3, 24) {real, imag} */,
  {32'h3f909b94, 32'h3fd8c1ff} /* (27, 3, 23) {real, imag} */,
  {32'h3fe946a3, 32'h4029a855} /* (27, 3, 22) {real, imag} */,
  {32'h3fac9610, 32'h402c6056} /* (27, 3, 21) {real, imag} */,
  {32'hbf79c520, 32'h3fc13282} /* (27, 3, 20) {real, imag} */,
  {32'hbfba1c1b, 32'h40201bc2} /* (27, 3, 19) {real, imag} */,
  {32'h4049d2de, 32'h40a49ca2} /* (27, 3, 18) {real, imag} */,
  {32'h3fa26937, 32'h3fe7fadf} /* (27, 3, 17) {real, imag} */,
  {32'h3fb7a111, 32'h40213197} /* (27, 3, 16) {real, imag} */,
  {32'hbf59bc4c, 32'hbeaabf7a} /* (27, 3, 15) {real, imag} */,
  {32'hc09353c7, 32'hbed6673a} /* (27, 3, 14) {real, imag} */,
  {32'hc03ac4fd, 32'hc089c132} /* (27, 3, 13) {real, imag} */,
  {32'hbf83d2e0, 32'hc05d44c0} /* (27, 3, 12) {real, imag} */,
  {32'hbfb6ccd8, 32'hbf22a140} /* (27, 3, 11) {real, imag} */,
  {32'hc03c3c2c, 32'h3f0c552d} /* (27, 3, 10) {real, imag} */,
  {32'hbff6a01b, 32'hc01d23a1} /* (27, 3, 9) {real, imag} */,
  {32'hbec10c9e, 32'hbfa657e3} /* (27, 3, 8) {real, imag} */,
  {32'h3f9c2c41, 32'h3e3c2000} /* (27, 3, 7) {real, imag} */,
  {32'hc01a8732, 32'hbe41fabc} /* (27, 3, 6) {real, imag} */,
  {32'h3d88ec90, 32'h401db864} /* (27, 3, 5) {real, imag} */,
  {32'h400d272b, 32'h4099d501} /* (27, 3, 4) {real, imag} */,
  {32'h4023502a, 32'h4097c59b} /* (27, 3, 3) {real, imag} */,
  {32'h4013ea19, 32'h400853ca} /* (27, 3, 2) {real, imag} */,
  {32'h3f22139f, 32'h3f89e719} /* (27, 3, 1) {real, imag} */,
  {32'h3f3dbcff, 32'h3fd3b6b4} /* (27, 3, 0) {real, imag} */,
  {32'h3f5885b3, 32'h3f142448} /* (27, 2, 31) {real, imag} */,
  {32'h3fe38d45, 32'h3fa1ebce} /* (27, 2, 30) {real, imag} */,
  {32'h4053636e, 32'hbe623976} /* (27, 2, 29) {real, imag} */,
  {32'h3fe3ef70, 32'h3f4ed799} /* (27, 2, 28) {real, imag} */,
  {32'h40076cd9, 32'h403ecb4e} /* (27, 2, 27) {real, imag} */,
  {32'h4088fd81, 32'h40499588} /* (27, 2, 26) {real, imag} */,
  {32'h408420d2, 32'h3f1c8f70} /* (27, 2, 25) {real, imag} */,
  {32'h3fff1ae9, 32'h40024e78} /* (27, 2, 24) {real, imag} */,
  {32'hbf53a4ec, 32'h4014a4ba} /* (27, 2, 23) {real, imag} */,
  {32'h3f8953ae, 32'h40236e9c} /* (27, 2, 22) {real, imag} */,
  {32'h4086014b, 32'h4019d7c5} /* (27, 2, 21) {real, imag} */,
  {32'h402da5ea, 32'h3ff05191} /* (27, 2, 20) {real, imag} */,
  {32'h3f96894a, 32'h40ab63be} /* (27, 2, 19) {real, imag} */,
  {32'h4021a4f8, 32'h40cc2772} /* (27, 2, 18) {real, imag} */,
  {32'h3fcf4cca, 32'h40c07053} /* (27, 2, 17) {real, imag} */,
  {32'h4015f1e0, 32'h40a55ad5} /* (27, 2, 16) {real, imag} */,
  {32'h3ef69545, 32'hbeee41d8} /* (27, 2, 15) {real, imag} */,
  {32'hc02e8321, 32'h3de6a60c} /* (27, 2, 14) {real, imag} */,
  {32'hbfc16c1e, 32'hc010beaa} /* (27, 2, 13) {real, imag} */,
  {32'hbf9f4cb5, 32'hc05b875d} /* (27, 2, 12) {real, imag} */,
  {32'hbfa0da0e, 32'hc01116ec} /* (27, 2, 11) {real, imag} */,
  {32'h3ed8fff4, 32'hc0139bf7} /* (27, 2, 10) {real, imag} */,
  {32'h3f6a59db, 32'hc095b350} /* (27, 2, 9) {real, imag} */,
  {32'hbf998b22, 32'hc02bb511} /* (27, 2, 8) {real, imag} */,
  {32'h3e51fc54, 32'hbf884678} /* (27, 2, 7) {real, imag} */,
  {32'hbe32c23c, 32'hbf1557c2} /* (27, 2, 6) {real, imag} */,
  {32'h3f7d31bb, 32'h4028ff6e} /* (27, 2, 5) {real, imag} */,
  {32'h3fba47a8, 32'h40235d3a} /* (27, 2, 4) {real, imag} */,
  {32'h3fc85d95, 32'h404db895} /* (27, 2, 3) {real, imag} */,
  {32'h4088bfb6, 32'h4051cb9a} /* (27, 2, 2) {real, imag} */,
  {32'h4017c5a1, 32'h3fbb0b08} /* (27, 2, 1) {real, imag} */,
  {32'h3f8d95fc, 32'h3fb1d088} /* (27, 2, 0) {real, imag} */,
  {32'hbe0b1848, 32'h3efb366f} /* (27, 1, 31) {real, imag} */,
  {32'h3ef76a22, 32'h3fd663e2} /* (27, 1, 30) {real, imag} */,
  {32'h3f7953a1, 32'h40002ba2} /* (27, 1, 29) {real, imag} */,
  {32'hbf063a34, 32'h3f55dc5c} /* (27, 1, 28) {real, imag} */,
  {32'h3fcf9f20, 32'h401ca0f3} /* (27, 1, 27) {real, imag} */,
  {32'h405317b4, 32'h4013bcfc} /* (27, 1, 26) {real, imag} */,
  {32'h40403348, 32'h4029b606} /* (27, 1, 25) {real, imag} */,
  {32'h3f9b0e19, 32'h3f83d3b6} /* (27, 1, 24) {real, imag} */,
  {32'hbea1b6ae, 32'h3fa3687c} /* (27, 1, 23) {real, imag} */,
  {32'h3e67ad98, 32'h405cd8cf} /* (27, 1, 22) {real, imag} */,
  {32'h3fe201cd, 32'h406e0f86} /* (27, 1, 21) {real, imag} */,
  {32'h4076d79d, 32'h400313ea} /* (27, 1, 20) {real, imag} */,
  {32'h3f761ff8, 32'h40b373c7} /* (27, 1, 19) {real, imag} */,
  {32'h3d416ce0, 32'h40d4023c} /* (27, 1, 18) {real, imag} */,
  {32'hbecfa014, 32'h40f4e042} /* (27, 1, 17) {real, imag} */,
  {32'h3fcb36ef, 32'h40a4a253} /* (27, 1, 16) {real, imag} */,
  {32'h3f76139d, 32'h3eb044ec} /* (27, 1, 15) {real, imag} */,
  {32'hbf942c57, 32'hbfcd815c} /* (27, 1, 14) {real, imag} */,
  {32'hbf944889, 32'hbfbf6c09} /* (27, 1, 13) {real, imag} */,
  {32'hbf129211, 32'hbffe6bbd} /* (27, 1, 12) {real, imag} */,
  {32'h3f992399, 32'hc04999e7} /* (27, 1, 11) {real, imag} */,
  {32'hbee82508, 32'hc067dcb8} /* (27, 1, 10) {real, imag} */,
  {32'hbe883eb8, 32'hc0af76db} /* (27, 1, 9) {real, imag} */,
  {32'hc00b9933, 32'hc0a4b02b} /* (27, 1, 8) {real, imag} */,
  {32'hc008e69a, 32'hc01383ff} /* (27, 1, 7) {real, imag} */,
  {32'hc0165d50, 32'h3f18734e} /* (27, 1, 6) {real, imag} */,
  {32'h3f8b2fd9, 32'h3f81a75c} /* (27, 1, 5) {real, imag} */,
  {32'h3f886ffd, 32'hbee514b5} /* (27, 1, 4) {real, imag} */,
  {32'hbf133b1b, 32'h3ff24b90} /* (27, 1, 3) {real, imag} */,
  {32'h3eafc7ea, 32'h405af4e4} /* (27, 1, 2) {real, imag} */,
  {32'h3ff2cbe3, 32'h3fba1748} /* (27, 1, 1) {real, imag} */,
  {32'h3fca0c38, 32'h3e8825e8} /* (27, 1, 0) {real, imag} */,
  {32'h3c77c3f0, 32'h3dd56508} /* (27, 0, 31) {real, imag} */,
  {32'h3f498e21, 32'h3f0a4718} /* (27, 0, 30) {real, imag} */,
  {32'h3effb5af, 32'h40011877} /* (27, 0, 29) {real, imag} */,
  {32'hbf223992, 32'h3e8ad38e} /* (27, 0, 28) {real, imag} */,
  {32'h3ff15a78, 32'h3ef80e34} /* (27, 0, 27) {real, imag} */,
  {32'h4060b48a, 32'h3f9d709a} /* (27, 0, 26) {real, imag} */,
  {32'h3ffcf6cd, 32'h3f91b86a} /* (27, 0, 25) {real, imag} */,
  {32'h3f9668a8, 32'h3efc3847} /* (27, 0, 24) {real, imag} */,
  {32'h3f96d8f6, 32'hbf0b4476} /* (27, 0, 23) {real, imag} */,
  {32'h3f31989a, 32'h3f489870} /* (27, 0, 22) {real, imag} */,
  {32'h3f107932, 32'h3fc10338} /* (27, 0, 21) {real, imag} */,
  {32'h407fd350, 32'h3f8dea08} /* (27, 0, 20) {real, imag} */,
  {32'h40172c40, 32'h4010b356} /* (27, 0, 19) {real, imag} */,
  {32'h3fcf79c4, 32'h40382734} /* (27, 0, 18) {real, imag} */,
  {32'h3ef7ff18, 32'h3fcd7986} /* (27, 0, 17) {real, imag} */,
  {32'hbf54d43a, 32'h3f6cc9e1} /* (27, 0, 16) {real, imag} */,
  {32'hbf1d52a0, 32'h3e00e47b} /* (27, 0, 15) {real, imag} */,
  {32'hbfbfa2d6, 32'hbfad490e} /* (27, 0, 14) {real, imag} */,
  {32'hbe791d0c, 32'hbfb93300} /* (27, 0, 13) {real, imag} */,
  {32'hbc2864e0, 32'hc00c0678} /* (27, 0, 12) {real, imag} */,
  {32'h3e485812, 32'hbffb04aa} /* (27, 0, 11) {real, imag} */,
  {32'hbfabd68d, 32'hbf97babd} /* (27, 0, 10) {real, imag} */,
  {32'hbf39993b, 32'hbfc89ba0} /* (27, 0, 9) {real, imag} */,
  {32'hbec6cb85, 32'hc046b0ca} /* (27, 0, 8) {real, imag} */,
  {32'hbf658b20, 32'hbfc939a3} /* (27, 0, 7) {real, imag} */,
  {32'hbff1a2b8, 32'h3eda0001} /* (27, 0, 6) {real, imag} */,
  {32'hbd58bcc0, 32'hbf3dd043} /* (27, 0, 5) {real, imag} */,
  {32'h3ed89e86, 32'hbef07906} /* (27, 0, 4) {real, imag} */,
  {32'h3e2538a8, 32'h3fc6a460} /* (27, 0, 3) {real, imag} */,
  {32'hbfebcc72, 32'h3fce4cb0} /* (27, 0, 2) {real, imag} */,
  {32'hbf239bac, 32'hbcf018c0} /* (27, 0, 1) {real, imag} */,
  {32'h3fac9f5c, 32'hbf946464} /* (27, 0, 0) {real, imag} */,
  {32'h3eb8ed12, 32'h3eafd44d} /* (26, 31, 31) {real, imag} */,
  {32'h3f1f0261, 32'hbe7a1fa0} /* (26, 31, 30) {real, imag} */,
  {32'hbf39ba04, 32'hbfc854b0} /* (26, 31, 29) {real, imag} */,
  {32'h3f3c28c2, 32'hbe8f6842} /* (26, 31, 28) {real, imag} */,
  {32'h40411b32, 32'h3f223875} /* (26, 31, 27) {real, imag} */,
  {32'h3fb1dd32, 32'h40282e34} /* (26, 31, 26) {real, imag} */,
  {32'h3f17ad3a, 32'h3f4183bb} /* (26, 31, 25) {real, imag} */,
  {32'hbf2e28be, 32'hbf8a685a} /* (26, 31, 24) {real, imag} */,
  {32'h3da1db08, 32'hbcd7fd20} /* (26, 31, 23) {real, imag} */,
  {32'hbf2b29da, 32'hbfe38665} /* (26, 31, 22) {real, imag} */,
  {32'hbf0f29a9, 32'hc021feb9} /* (26, 31, 21) {real, imag} */,
  {32'hc01a9a83, 32'hbec1c3f1} /* (26, 31, 20) {real, imag} */,
  {32'hc014360e, 32'hbfe36b9f} /* (26, 31, 19) {real, imag} */,
  {32'hbf640bfc, 32'hbfeaf9c5} /* (26, 31, 18) {real, imag} */,
  {32'hbf8802a5, 32'h3d8ab4a0} /* (26, 31, 17) {real, imag} */,
  {32'hbf539d04, 32'h3f2703fe} /* (26, 31, 16) {real, imag} */,
  {32'hbf915c2e, 32'h3ffc1407} /* (26, 31, 15) {real, imag} */,
  {32'hbfb94b35, 32'h3fcc79fb} /* (26, 31, 14) {real, imag} */,
  {32'hbfa26463, 32'h3e8c92f0} /* (26, 31, 13) {real, imag} */,
  {32'hbd8278c0, 32'h3d0242e0} /* (26, 31, 12) {real, imag} */,
  {32'hbec7de23, 32'h3f229546} /* (26, 31, 11) {real, imag} */,
  {32'h3f723f84, 32'h401141ba} /* (26, 31, 10) {real, imag} */,
  {32'h3f7eace8, 32'h3eeacf04} /* (26, 31, 9) {real, imag} */,
  {32'h3fcd1d5f, 32'hbf8ca9b2} /* (26, 31, 8) {real, imag} */,
  {32'hbf40fb5e, 32'h3ef54444} /* (26, 31, 7) {real, imag} */,
  {32'h3f36fdbd, 32'h3c12aa80} /* (26, 31, 6) {real, imag} */,
  {32'h3f9d1f9e, 32'h3e89a1b4} /* (26, 31, 5) {real, imag} */,
  {32'hbe06e804, 32'h3fe55ae2} /* (26, 31, 4) {real, imag} */,
  {32'h3f403b5f, 32'h3fbda512} /* (26, 31, 3) {real, imag} */,
  {32'h40422443, 32'h3f0790c1} /* (26, 31, 2) {real, imag} */,
  {32'h40368687, 32'h3d1ac280} /* (26, 31, 1) {real, imag} */,
  {32'h3ff823fb, 32'hbe524754} /* (26, 31, 0) {real, imag} */,
  {32'h3f53d6c4, 32'h3f02b434} /* (26, 30, 31) {real, imag} */,
  {32'h3ff07be2, 32'hbe19cc40} /* (26, 30, 30) {real, imag} */,
  {32'hbf1b04ce, 32'hc00cb18c} /* (26, 30, 29) {real, imag} */,
  {32'h3eafd1dc, 32'hbf00e864} /* (26, 30, 28) {real, imag} */,
  {32'h40460ee6, 32'h3f36e17e} /* (26, 30, 27) {real, imag} */,
  {32'h401aedaa, 32'h40165540} /* (26, 30, 26) {real, imag} */,
  {32'hbf36faec, 32'h3f67edac} /* (26, 30, 25) {real, imag} */,
  {32'hbf820cdc, 32'hbfbd55da} /* (26, 30, 24) {real, imag} */,
  {32'hbf2c724c, 32'h3fa9cc66} /* (26, 30, 23) {real, imag} */,
  {32'hbfcee29f, 32'hbe97bfb8} /* (26, 30, 22) {real, imag} */,
  {32'hbe7ee898, 32'hc0793ec1} /* (26, 30, 21) {real, imag} */,
  {32'hbd0f5e00, 32'hc007de78} /* (26, 30, 20) {real, imag} */,
  {32'hbf3389d3, 32'hc0363e8f} /* (26, 30, 19) {real, imag} */,
  {32'hbeeae7e6, 32'hc04a6128} /* (26, 30, 18) {real, imag} */,
  {32'hbfa6dab1, 32'hbfcd4105} /* (26, 30, 17) {real, imag} */,
  {32'hbf6da475, 32'hbec20cba} /* (26, 30, 16) {real, imag} */,
  {32'hbe3e7d1c, 32'hbbab4700} /* (26, 30, 15) {real, imag} */,
  {32'hbff6adf8, 32'hbf918d4d} /* (26, 30, 14) {real, imag} */,
  {32'hbf432c20, 32'h3f1f0616} /* (26, 30, 13) {real, imag} */,
  {32'hbf49baab, 32'h4009c74e} /* (26, 30, 12) {real, imag} */,
  {32'hbfc3c1d9, 32'h3f4b7660} /* (26, 30, 11) {real, imag} */,
  {32'h3e424ea4, 32'h3fa75274} /* (26, 30, 10) {real, imag} */,
  {32'hbed17bee, 32'h3f0ff126} /* (26, 30, 9) {real, imag} */,
  {32'h3f87b600, 32'hbf5085c2} /* (26, 30, 8) {real, imag} */,
  {32'h3fd56919, 32'h3fc79813} /* (26, 30, 7) {real, imag} */,
  {32'h3ec175c0, 32'h3fd352e5} /* (26, 30, 6) {real, imag} */,
  {32'hbeff6108, 32'h3ea7c080} /* (26, 30, 5) {real, imag} */,
  {32'h3f0625ca, 32'h3ff99898} /* (26, 30, 4) {real, imag} */,
  {32'h3fd1c968, 32'h4018cb4a} /* (26, 30, 3) {real, imag} */,
  {32'h3fe3d8a6, 32'h3f5f5530} /* (26, 30, 2) {real, imag} */,
  {32'hbf879fae, 32'hbeb40b58} /* (26, 30, 1) {real, imag} */,
  {32'hbf7479e0, 32'hbffcc0ac} /* (26, 30, 0) {real, imag} */,
  {32'h3f258f1e, 32'hbe4db7dc} /* (26, 29, 31) {real, imag} */,
  {32'h3e91ac6c, 32'h3eb5ef50} /* (26, 29, 30) {real, imag} */,
  {32'hbf3a2dd6, 32'hbdf6b610} /* (26, 29, 29) {real, imag} */,
  {32'h3fbf73a2, 32'hbe94f58c} /* (26, 29, 28) {real, imag} */,
  {32'h402ef59b, 32'hbe20baec} /* (26, 29, 27) {real, imag} */,
  {32'h3fd82dac, 32'h4010824a} /* (26, 29, 26) {real, imag} */,
  {32'hbd4a2210, 32'h3feccc6a} /* (26, 29, 25) {real, imag} */,
  {32'h3fda64de, 32'hbfba0b9e} /* (26, 29, 24) {real, imag} */,
  {32'hbf81a156, 32'h3f4dda1c} /* (26, 29, 23) {real, imag} */,
  {32'hbeb35b82, 32'hbdc1a8c0} /* (26, 29, 22) {real, imag} */,
  {32'h3f8db77a, 32'hbfea45a8} /* (26, 29, 21) {real, imag} */,
  {32'h3fb995fc, 32'hc06e444a} /* (26, 29, 20) {real, imag} */,
  {32'hbe2f5924, 32'hc0296a64} /* (26, 29, 19) {real, imag} */,
  {32'hbf2c4174, 32'hbfac4ad1} /* (26, 29, 18) {real, imag} */,
  {32'h3fb0ce7e, 32'hbf5678ef} /* (26, 29, 17) {real, imag} */,
  {32'h3fba8f14, 32'h400d16ec} /* (26, 29, 16) {real, imag} */,
  {32'h401e72fa, 32'h40007709} /* (26, 29, 15) {real, imag} */,
  {32'h403f8adc, 32'hbfafd9f4} /* (26, 29, 14) {real, imag} */,
  {32'h4014fabc, 32'hbf0fba90} /* (26, 29, 13) {real, imag} */,
  {32'hbef34fae, 32'h3edcb68c} /* (26, 29, 12) {real, imag} */,
  {32'hbf3cc61c, 32'h3f25540e} /* (26, 29, 11) {real, imag} */,
  {32'h3e88cdd4, 32'h3f9de02a} /* (26, 29, 10) {real, imag} */,
  {32'hbf97f64b, 32'h3f46646a} /* (26, 29, 9) {real, imag} */,
  {32'h3f8aec04, 32'hbe5439a8} /* (26, 29, 8) {real, imag} */,
  {32'h40525093, 32'h4006f804} /* (26, 29, 7) {real, imag} */,
  {32'hbf3d7286, 32'h400e1940} /* (26, 29, 6) {real, imag} */,
  {32'hc00e9236, 32'hbf5de2cf} /* (26, 29, 5) {real, imag} */,
  {32'h3dc4e7a0, 32'hbf6c5e0a} /* (26, 29, 4) {real, imag} */,
  {32'h3f83e598, 32'h3f4462fa} /* (26, 29, 3) {real, imag} */,
  {32'hbfe570d2, 32'h3ed9ed38} /* (26, 29, 2) {real, imag} */,
  {32'hc04ba56d, 32'hbef74d6a} /* (26, 29, 1) {real, imag} */,
  {32'hbf3b00a3, 32'hbfbafe72} /* (26, 29, 0) {real, imag} */,
  {32'h3ec67e6c, 32'hc0203788} /* (26, 28, 31) {real, imag} */,
  {32'hbfa10bdc, 32'hbf20461a} /* (26, 28, 30) {real, imag} */,
  {32'hbf1bb9a8, 32'h3f9e18f8} /* (26, 28, 29) {real, imag} */,
  {32'h400e78d6, 32'h3fb10c9c} /* (26, 28, 28) {real, imag} */,
  {32'h40353528, 32'hbc226300} /* (26, 28, 27) {real, imag} */,
  {32'h3fb89bf8, 32'h3f8325d7} /* (26, 28, 26) {real, imag} */,
  {32'hbeffb00c, 32'h3d81d240} /* (26, 28, 25) {real, imag} */,
  {32'h402c20b6, 32'hbf48f1d0} /* (26, 28, 24) {real, imag} */,
  {32'h3fad650c, 32'h3c544f80} /* (26, 28, 23) {real, imag} */,
  {32'h3ff21cd8, 32'hbf95ed7f} /* (26, 28, 22) {real, imag} */,
  {32'h3fb512ba, 32'h3eec4af2} /* (26, 28, 21) {real, imag} */,
  {32'hc054925c, 32'hbf149c81} /* (26, 28, 20) {real, imag} */,
  {32'hc0271f66, 32'h3d296000} /* (26, 28, 19) {real, imag} */,
  {32'hbe0bbfcc, 32'hbf83d3b4} /* (26, 28, 18) {real, imag} */,
  {32'hbf2130cd, 32'hbf8bbff5} /* (26, 28, 17) {real, imag} */,
  {32'hc00da723, 32'h4019e9f2} /* (26, 28, 16) {real, imag} */,
  {32'h3d0c3340, 32'h40353e62} /* (26, 28, 15) {real, imag} */,
  {32'h401fc758, 32'h3f1a58d2} /* (26, 28, 14) {real, imag} */,
  {32'h401f99cc, 32'hbf47259e} /* (26, 28, 13) {real, imag} */,
  {32'h3f494c2a, 32'hc00142c0} /* (26, 28, 12) {real, imag} */,
  {32'h400e0966, 32'hbf4283d1} /* (26, 28, 11) {real, imag} */,
  {32'h4021f100, 32'hbf9ab006} /* (26, 28, 10) {real, imag} */,
  {32'hbee0487c, 32'h3fc29abe} /* (26, 28, 9) {real, imag} */,
  {32'hbf9c4bfa, 32'h3f4f6a7c} /* (26, 28, 8) {real, imag} */,
  {32'hbe424c50, 32'h3f23bbfa} /* (26, 28, 7) {real, imag} */,
  {32'hbf48184c, 32'h3f12922e} /* (26, 28, 6) {real, imag} */,
  {32'hbf5aa14f, 32'h3f44abe0} /* (26, 28, 5) {real, imag} */,
  {32'h3f4d9178, 32'h3f875932} /* (26, 28, 4) {real, imag} */,
  {32'h3f547080, 32'h3f55adc2} /* (26, 28, 3) {real, imag} */,
  {32'h3eec14a6, 32'h3f2366cc} /* (26, 28, 2) {real, imag} */,
  {32'h3f79ae2f, 32'hbe85034e} /* (26, 28, 1) {real, imag} */,
  {32'h3f07555a, 32'hbf3fd885} /* (26, 28, 0) {real, imag} */,
  {32'hbeb6c85e, 32'hbf301fb5} /* (26, 27, 31) {real, imag} */,
  {32'hbfaabd13, 32'hbf38880c} /* (26, 27, 30) {real, imag} */,
  {32'hbf4e94ad, 32'h3ff33082} /* (26, 27, 29) {real, imag} */,
  {32'hbfb41334, 32'h407a471c} /* (26, 27, 28) {real, imag} */,
  {32'h3e9fef52, 32'h3f475cea} /* (26, 27, 27) {real, imag} */,
  {32'h405f5621, 32'hbffa907d} /* (26, 27, 26) {real, imag} */,
  {32'h3fe22904, 32'hc01513ef} /* (26, 27, 25) {real, imag} */,
  {32'hbed6bff8, 32'h4004c36b} /* (26, 27, 24) {real, imag} */,
  {32'h3f7ad5b4, 32'h3f669c92} /* (26, 27, 23) {real, imag} */,
  {32'h3f55707d, 32'h3f1252bf} /* (26, 27, 22) {real, imag} */,
  {32'h3f7c7c10, 32'h3f11a9c5} /* (26, 27, 21) {real, imag} */,
  {32'hbfb3d9ba, 32'h3eafd170} /* (26, 27, 20) {real, imag} */,
  {32'hc02ead05, 32'hbf0cf096} /* (26, 27, 19) {real, imag} */,
  {32'hc0069107, 32'hbfd4735c} /* (26, 27, 18) {real, imag} */,
  {32'hc017aa0b, 32'h3f8b8f7d} /* (26, 27, 17) {real, imag} */,
  {32'hc001465e, 32'h3f641c35} /* (26, 27, 16) {real, imag} */,
  {32'h3dff66d0, 32'hbf7d95e2} /* (26, 27, 15) {real, imag} */,
  {32'h3f1a650e, 32'h3f54379a} /* (26, 27, 14) {real, imag} */,
  {32'h3f07fe3e, 32'h3fa06012} /* (26, 27, 13) {real, imag} */,
  {32'hbd8ec9c8, 32'hc0034e2e} /* (26, 27, 12) {real, imag} */,
  {32'h3fffd3f0, 32'hbeb263aa} /* (26, 27, 11) {real, imag} */,
  {32'h3fd0ea1a, 32'hbf056220} /* (26, 27, 10) {real, imag} */,
  {32'hbfe3aed1, 32'h3fd2a02c} /* (26, 27, 9) {real, imag} */,
  {32'hc05cd75c, 32'h3f68dd14} /* (26, 27, 8) {real, imag} */,
  {32'hc03ab422, 32'hbeead05c} /* (26, 27, 7) {real, imag} */,
  {32'hbebc3016, 32'h3e404138} /* (26, 27, 6) {real, imag} */,
  {32'h3f7be7f8, 32'hbf0a1d35} /* (26, 27, 5) {real, imag} */,
  {32'h3f196656, 32'hbf494bec} /* (26, 27, 4) {real, imag} */,
  {32'h3f035b5b, 32'hbe1c2038} /* (26, 27, 3) {real, imag} */,
  {32'h3f4efadc, 32'hbfb15e8c} /* (26, 27, 2) {real, imag} */,
  {32'h3efd4e2c, 32'h3f2680a6} /* (26, 27, 1) {real, imag} */,
  {32'hbf97c180, 32'h3f8c0d30} /* (26, 27, 0) {real, imag} */,
  {32'hbeecd59e, 32'h3ed393fa} /* (26, 26, 31) {real, imag} */,
  {32'hbfb8c3cb, 32'h3e11917c} /* (26, 26, 30) {real, imag} */,
  {32'hbf951d1a, 32'h3fccc106} /* (26, 26, 29) {real, imag} */,
  {32'hbfacd871, 32'h401f294d} /* (26, 26, 28) {real, imag} */,
  {32'hbcbe0438, 32'h3faaf29c} /* (26, 26, 27) {real, imag} */,
  {32'h3f959911, 32'hbe88808c} /* (26, 26, 26) {real, imag} */,
  {32'h3f19eafe, 32'hbefb783c} /* (26, 26, 25) {real, imag} */,
  {32'hbff87bb2, 32'h3fcc83d4} /* (26, 26, 24) {real, imag} */,
  {32'hbe942e72, 32'h3ff5789d} /* (26, 26, 23) {real, imag} */,
  {32'h3c2db580, 32'h3faaf530} /* (26, 26, 22) {real, imag} */,
  {32'hbede3b16, 32'h3f285add} /* (26, 26, 21) {real, imag} */,
  {32'hbeb7c714, 32'h3ece062e} /* (26, 26, 20) {real, imag} */,
  {32'hbd5e17c0, 32'hbe0a2e58} /* (26, 26, 19) {real, imag} */,
  {32'hbfd35895, 32'hc019f8a4} /* (26, 26, 18) {real, imag} */,
  {32'hc03db6dc, 32'h3f503bf5} /* (26, 26, 17) {real, imag} */,
  {32'hbe9efa02, 32'h3ea8f856} /* (26, 26, 16) {real, imag} */,
  {32'hbf3d5a35, 32'hc04fc2d0} /* (26, 26, 15) {real, imag} */,
  {32'hbf3e2c50, 32'hbfca7dbf} /* (26, 26, 14) {real, imag} */,
  {32'hbe95a5f0, 32'hbe9e30e4} /* (26, 26, 13) {real, imag} */,
  {32'hbf2d6318, 32'hbeab90b6} /* (26, 26, 12) {real, imag} */,
  {32'h3f1e326e, 32'h3f47ee6d} /* (26, 26, 11) {real, imag} */,
  {32'hbf8ef085, 32'h3f443e3b} /* (26, 26, 10) {real, imag} */,
  {32'hbfe18672, 32'h3fcec66b} /* (26, 26, 9) {real, imag} */,
  {32'hbf9aee5c, 32'h40130914} /* (26, 26, 8) {real, imag} */,
  {32'hbfde002b, 32'hbf96eddb} /* (26, 26, 7) {real, imag} */,
  {32'hbfd06acc, 32'hc0353361} /* (26, 26, 6) {real, imag} */,
  {32'h3f4d0a98, 32'hbf9dee2a} /* (26, 26, 5) {real, imag} */,
  {32'hbfb488f8, 32'hc009c9ab} /* (26, 26, 4) {real, imag} */,
  {32'hc007bd18, 32'hc0782adc} /* (26, 26, 3) {real, imag} */,
  {32'hbf34919a, 32'hc08d2880} /* (26, 26, 2) {real, imag} */,
  {32'hbf94e038, 32'hbf6e6828} /* (26, 26, 1) {real, imag} */,
  {32'hbf95d82c, 32'h3f1e956e} /* (26, 26, 0) {real, imag} */,
  {32'hbfb9cd65, 32'h3f8dc7e8} /* (26, 25, 31) {real, imag} */,
  {32'hc009b8ce, 32'h3ef28876} /* (26, 25, 30) {real, imag} */,
  {32'hbfc09ebe, 32'h3eec9cc6} /* (26, 25, 29) {real, imag} */,
  {32'hbf40a07c, 32'h3fa9519c} /* (26, 25, 28) {real, imag} */,
  {32'h3f4e0d22, 32'h401ba548} /* (26, 25, 27) {real, imag} */,
  {32'h3ef6ba7e, 32'h3ff6ce00} /* (26, 25, 26) {real, imag} */,
  {32'h3dc5b4e0, 32'h400855cf} /* (26, 25, 25) {real, imag} */,
  {32'hbfc2662a, 32'h3f752d1c} /* (26, 25, 24) {real, imag} */,
  {32'hbf4407aa, 32'h3fc1059c} /* (26, 25, 23) {real, imag} */,
  {32'hbf8bad89, 32'h401aace2} /* (26, 25, 22) {real, imag} */,
  {32'hbfe1cf11, 32'h3f8767b0} /* (26, 25, 21) {real, imag} */,
  {32'h3e90302c, 32'h3f311826} /* (26, 25, 20) {real, imag} */,
  {32'h400c355c, 32'h4003175f} /* (26, 25, 19) {real, imag} */,
  {32'hbe5830e0, 32'hbf3e8776} /* (26, 25, 18) {real, imag} */,
  {32'hc022e036, 32'h3f303456} /* (26, 25, 17) {real, imag} */,
  {32'h3ff8d0db, 32'h3f808a14} /* (26, 25, 16) {real, imag} */,
  {32'h3ffec784, 32'hbed40a5a} /* (26, 25, 15) {real, imag} */,
  {32'h3fdd8fa8, 32'hbf50b738} /* (26, 25, 14) {real, imag} */,
  {32'h403b6078, 32'hbf5b8e02} /* (26, 25, 13) {real, imag} */,
  {32'h3e32b5a0, 32'hbdec4f70} /* (26, 25, 12) {real, imag} */,
  {32'h3f562d46, 32'hbde22590} /* (26, 25, 11) {real, imag} */,
  {32'hbf88a8da, 32'hbfca1418} /* (26, 25, 10) {real, imag} */,
  {32'hbff1ecc7, 32'hbd38ee20} /* (26, 25, 9) {real, imag} */,
  {32'h3f599ccc, 32'h40263375} /* (26, 25, 8) {real, imag} */,
  {32'h3fc607e9, 32'hbf8587d1} /* (26, 25, 7) {real, imag} */,
  {32'h3e386414, 32'hc034b730} /* (26, 25, 6) {real, imag} */,
  {32'h3e05b464, 32'hc0198208} /* (26, 25, 5) {real, imag} */,
  {32'hbfa5c849, 32'hc0170fde} /* (26, 25, 4) {real, imag} */,
  {32'hc00b0613, 32'hc05ba6cc} /* (26, 25, 3) {real, imag} */,
  {32'hbf396e18, 32'hbfac6e7b} /* (26, 25, 2) {real, imag} */,
  {32'hbf24bed2, 32'hc020a5d9} /* (26, 25, 1) {real, imag} */,
  {32'hbf27ac52, 32'hbf0d140c} /* (26, 25, 0) {real, imag} */,
  {32'hbfcf9ba5, 32'hbfb2cd24} /* (26, 24, 31) {real, imag} */,
  {32'hbe454338, 32'hbfdff0a9} /* (26, 24, 30) {real, imag} */,
  {32'h3f90c89d, 32'hbf8fdb06} /* (26, 24, 29) {real, imag} */,
  {32'h3f9f0c6e, 32'hbe1f3058} /* (26, 24, 28) {real, imag} */,
  {32'h3fc7b9c9, 32'h3fce0003} /* (26, 24, 27) {real, imag} */,
  {32'hbf1a2a10, 32'h40007ffa} /* (26, 24, 26) {real, imag} */,
  {32'h3da91e28, 32'h40985f9f} /* (26, 24, 25) {real, imag} */,
  {32'hbc47a840, 32'h402f0b02} /* (26, 24, 24) {real, imag} */,
  {32'h3f8af200, 32'h3fdb4228} /* (26, 24, 23) {real, imag} */,
  {32'hbfdcb314, 32'h3f07884e} /* (26, 24, 22) {real, imag} */,
  {32'hbffd7104, 32'h3ff4c4e4} /* (26, 24, 21) {real, imag} */,
  {32'hbe0d1118, 32'h3fd27bd8} /* (26, 24, 20) {real, imag} */,
  {32'h3ff86ad9, 32'h3f3e9734} /* (26, 24, 19) {real, imag} */,
  {32'h3f8306e7, 32'hbfc41db6} /* (26, 24, 18) {real, imag} */,
  {32'hbfaf3526, 32'h3f271a52} /* (26, 24, 17) {real, imag} */,
  {32'h40193f26, 32'hbefad2d4} /* (26, 24, 16) {real, imag} */,
  {32'h3ffa5fbc, 32'hc02f2ad3} /* (26, 24, 15) {real, imag} */,
  {32'h3fc5b277, 32'hc04121c9} /* (26, 24, 14) {real, imag} */,
  {32'h40d16606, 32'hbfade0ef} /* (26, 24, 13) {real, imag} */,
  {32'h40205827, 32'h3ec283d4} /* (26, 24, 12) {real, imag} */,
  {32'h4002050f, 32'hbdd0c5e8} /* (26, 24, 11) {real, imag} */,
  {32'h3ffb290d, 32'hc04cdd32} /* (26, 24, 10) {real, imag} */,
  {32'h3e55cb10, 32'h3ea9052c} /* (26, 24, 9) {real, imag} */,
  {32'h3e6b4fa8, 32'h3fa9ebb8} /* (26, 24, 8) {real, imag} */,
  {32'h3f22dae7, 32'hc0001fee} /* (26, 24, 7) {real, imag} */,
  {32'hbeb8b406, 32'hbeadf734} /* (26, 24, 6) {real, imag} */,
  {32'hbfbe590b, 32'hbf89d837} /* (26, 24, 5) {real, imag} */,
  {32'hbfa841a4, 32'hbf0716b7} /* (26, 24, 4) {real, imag} */,
  {32'hbf0af1a1, 32'hbfdb0f1b} /* (26, 24, 3) {real, imag} */,
  {32'hbf01fc54, 32'hbe8aaa18} /* (26, 24, 2) {real, imag} */,
  {32'h3f41c800, 32'hbe393eec} /* (26, 24, 1) {real, imag} */,
  {32'h3f16de4c, 32'h3e88d377} /* (26, 24, 0) {real, imag} */,
  {32'hbf1df689, 32'h3dac3240} /* (26, 23, 31) {real, imag} */,
  {32'hbdbdc5f0, 32'h3f314bb4} /* (26, 23, 30) {real, imag} */,
  {32'h3f37343a, 32'hbd8235f8} /* (26, 23, 29) {real, imag} */,
  {32'h3e574540, 32'h3e074c20} /* (26, 23, 28) {real, imag} */,
  {32'h3fedd428, 32'h4057e526} /* (26, 23, 27) {real, imag} */,
  {32'hbea8ab64, 32'h405dd35a} /* (26, 23, 26) {real, imag} */,
  {32'h3f3d401e, 32'h406076b1} /* (26, 23, 25) {real, imag} */,
  {32'h400754e7, 32'h404fc388} /* (26, 23, 24) {real, imag} */,
  {32'h3dd3f3e0, 32'h402292a9} /* (26, 23, 23) {real, imag} */,
  {32'h3ef9d2e4, 32'h3feb2d86} /* (26, 23, 22) {real, imag} */,
  {32'h3eedaea3, 32'h400bbbda} /* (26, 23, 21) {real, imag} */,
  {32'h3e81871c, 32'h3fa402f7} /* (26, 23, 20) {real, imag} */,
  {32'hbfc57397, 32'h3c3b9880} /* (26, 23, 19) {real, imag} */,
  {32'hbfc39a53, 32'hbf8fd005} /* (26, 23, 18) {real, imag} */,
  {32'hc0417b1e, 32'h3fcd107a} /* (26, 23, 17) {real, imag} */,
  {32'h3f43f8af, 32'h3d3ad480} /* (26, 23, 16) {real, imag} */,
  {32'h3fbc575e, 32'hc025ff94} /* (26, 23, 15) {real, imag} */,
  {32'hbec55bae, 32'hc046c4b2} /* (26, 23, 14) {real, imag} */,
  {32'h406f73be, 32'hbf6c20b6} /* (26, 23, 13) {real, imag} */,
  {32'h3fac416d, 32'h3f06cc0e} /* (26, 23, 12) {real, imag} */,
  {32'h3f1a5811, 32'h3f287798} /* (26, 23, 11) {real, imag} */,
  {32'h403c80e3, 32'hbf31b7fd} /* (26, 23, 10) {real, imag} */,
  {32'h40001812, 32'h3ef6965c} /* (26, 23, 9) {real, imag} */,
  {32'hbdf488f8, 32'hbd458a70} /* (26, 23, 8) {real, imag} */,
  {32'hbe4ca6c4, 32'hbfa2f991} /* (26, 23, 7) {real, imag} */,
  {32'hbf2b9986, 32'h3fc8d5a3} /* (26, 23, 6) {real, imag} */,
  {32'hc0370b69, 32'h3f646f2b} /* (26, 23, 5) {real, imag} */,
  {32'hbfe1fcf0, 32'hbe4aacd8} /* (26, 23, 4) {real, imag} */,
  {32'hbf0928a8, 32'hbef7eb2c} /* (26, 23, 3) {real, imag} */,
  {32'h3e8d02dc, 32'hbf8ca284} /* (26, 23, 2) {real, imag} */,
  {32'h3ff5578a, 32'h3e5b8d90} /* (26, 23, 1) {real, imag} */,
  {32'h3f84aabd, 32'h3dd380a8} /* (26, 23, 0) {real, imag} */,
  {32'h3dae3c20, 32'h3dcc81d8} /* (26, 22, 31) {real, imag} */,
  {32'h3f6a6249, 32'h3fd7dd47} /* (26, 22, 30) {real, imag} */,
  {32'h3f230010, 32'h3fa6f478} /* (26, 22, 29) {real, imag} */,
  {32'h3fc4a038, 32'h3f629200} /* (26, 22, 28) {real, imag} */,
  {32'h40443c77, 32'h40430430} /* (26, 22, 27) {real, imag} */,
  {32'h4008bd74, 32'h405a11a8} /* (26, 22, 26) {real, imag} */,
  {32'hbf11738e, 32'h3feda1e2} /* (26, 22, 25) {real, imag} */,
  {32'hbf48f87a, 32'h4000ab6d} /* (26, 22, 24) {real, imag} */,
  {32'hbfa97b06, 32'h3fc4b56e} /* (26, 22, 23) {real, imag} */,
  {32'hbf8e7dba, 32'h3dccb568} /* (26, 22, 22) {real, imag} */,
  {32'hbf588a53, 32'hbfe47342} /* (26, 22, 21) {real, imag} */,
  {32'hbdef8408, 32'hbf200846} /* (26, 22, 20) {real, imag} */,
  {32'hc02b0ff6, 32'h3e840f00} /* (26, 22, 19) {real, imag} */,
  {32'hbfea38ca, 32'h3d60f7c0} /* (26, 22, 18) {real, imag} */,
  {32'hc03762ed, 32'h3fd620b2} /* (26, 22, 17) {real, imag} */,
  {32'hbfe7ad64, 32'h40054b13} /* (26, 22, 16) {real, imag} */,
  {32'h3ec17f0a, 32'h3eb6a20e} /* (26, 22, 15) {real, imag} */,
  {32'hbfebda4a, 32'hbf49cd8a} /* (26, 22, 14) {real, imag} */,
  {32'hbf1385fc, 32'hbff75a70} /* (26, 22, 13) {real, imag} */,
  {32'h3f71abcb, 32'hc024288b} /* (26, 22, 12) {real, imag} */,
  {32'h4007d7f7, 32'hbfd92914} /* (26, 22, 11) {real, imag} */,
  {32'h4011036f, 32'hbdf4a598} /* (26, 22, 10) {real, imag} */,
  {32'h4023808f, 32'h40106c78} /* (26, 22, 9) {real, imag} */,
  {32'h3fb9324e, 32'h3f85c4e7} /* (26, 22, 8) {real, imag} */,
  {32'h3ef3b7ca, 32'h401a64be} /* (26, 22, 7) {real, imag} */,
  {32'h3cbcac00, 32'h3fca8354} /* (26, 22, 6) {real, imag} */,
  {32'hbfdb9ed0, 32'hbe837190} /* (26, 22, 5) {real, imag} */,
  {32'hc0038781, 32'hbf563c82} /* (26, 22, 4) {real, imag} */,
  {32'hbf8b32f9, 32'h3ed01a70} /* (26, 22, 3) {real, imag} */,
  {32'hbecb4b40, 32'hbf9e7de6} /* (26, 22, 2) {real, imag} */,
  {32'h3fa8660a, 32'h3f7690e4} /* (26, 22, 1) {real, imag} */,
  {32'h4028fbf2, 32'hbe55db0c} /* (26, 22, 0) {real, imag} */,
  {32'hbed10dbe, 32'hbf9e27bf} /* (26, 21, 31) {real, imag} */,
  {32'h3f9158ad, 32'hbfdf7204} /* (26, 21, 30) {real, imag} */,
  {32'h3fb4f2fe, 32'h3f82e369} /* (26, 21, 29) {real, imag} */,
  {32'h4005528c, 32'h3fb3dc84} /* (26, 21, 28) {real, imag} */,
  {32'h40249ea5, 32'h3fe5d972} /* (26, 21, 27) {real, imag} */,
  {32'h3fe4b485, 32'h4018d902} /* (26, 21, 26) {real, imag} */,
  {32'hbf07080e, 32'h3f892300} /* (26, 21, 25) {real, imag} */,
  {32'hbf6af5fe, 32'h3f1a0f90} /* (26, 21, 24) {real, imag} */,
  {32'hbf44e6bc, 32'hbf19ff8c} /* (26, 21, 23) {real, imag} */,
  {32'hbf2d8fef, 32'hc05f51fc} /* (26, 21, 22) {real, imag} */,
  {32'hbdc60c30, 32'hc0a7cd40} /* (26, 21, 21) {real, imag} */,
  {32'h3ef10fa4, 32'hbf006d5e} /* (26, 21, 20) {real, imag} */,
  {32'h3fc3870f, 32'h3fe5964a} /* (26, 21, 19) {real, imag} */,
  {32'h3e1ddbc4, 32'h40139316} /* (26, 21, 18) {real, imag} */,
  {32'hc00f1a82, 32'h3f9af7b1} /* (26, 21, 17) {real, imag} */,
  {32'hc031540e, 32'h3ee4b87e} /* (26, 21, 16) {real, imag} */,
  {32'h3fbab2bc, 32'hbed996a8} /* (26, 21, 15) {real, imag} */,
  {32'h3cb1fe00, 32'hbf257cad} /* (26, 21, 14) {real, imag} */,
  {32'hbff9ad44, 32'hbede5cd2} /* (26, 21, 13) {real, imag} */,
  {32'hbed53cc0, 32'hbf539673} /* (26, 21, 12) {real, imag} */,
  {32'h3fba3935, 32'hbf41eba1} /* (26, 21, 11) {real, imag} */,
  {32'h3f3ea733, 32'h3fd39faa} /* (26, 21, 10) {real, imag} */,
  {32'h3f48cc38, 32'h4028ae4b} /* (26, 21, 9) {real, imag} */,
  {32'h3e120d50, 32'h3f974da3} /* (26, 21, 8) {real, imag} */,
  {32'hbf1b665a, 32'h3fc311f5} /* (26, 21, 7) {real, imag} */,
  {32'h3ffd53fe, 32'hbf6010d2} /* (26, 21, 6) {real, imag} */,
  {32'h3fadc4b6, 32'hc010cb4d} /* (26, 21, 5) {real, imag} */,
  {32'h3f88094f, 32'hbfff2021} /* (26, 21, 4) {real, imag} */,
  {32'h3f4ea6fd, 32'hbf04f016} /* (26, 21, 3) {real, imag} */,
  {32'h3ec7494c, 32'hc0057e97} /* (26, 21, 2) {real, imag} */,
  {32'hbf1aecbc, 32'hbe5f7a4c} /* (26, 21, 1) {real, imag} */,
  {32'hbd47a920, 32'hbf2b3498} /* (26, 21, 0) {real, imag} */,
  {32'h3df9f644, 32'hbfd0a96e} /* (26, 20, 31) {real, imag} */,
  {32'h3ff202c7, 32'hc00b1c16} /* (26, 20, 30) {real, imag} */,
  {32'h4015ae20, 32'hbf2624b8} /* (26, 20, 29) {real, imag} */,
  {32'h3f93e160, 32'hbf93d694} /* (26, 20, 28) {real, imag} */,
  {32'h3ed04264, 32'hbeb522d8} /* (26, 20, 27) {real, imag} */,
  {32'h3e0c82c4, 32'h3f506de6} /* (26, 20, 26) {real, imag} */,
  {32'hbf859dfd, 32'h3f1685d3} /* (26, 20, 25) {real, imag} */,
  {32'hbe1622a8, 32'h3fa616eb} /* (26, 20, 24) {real, imag} */,
  {32'hbfac9548, 32'hbfea805a} /* (26, 20, 23) {real, imag} */,
  {32'hbf6756c4, 32'hc0755e80} /* (26, 20, 22) {real, imag} */,
  {32'h3ed9d2f2, 32'hc0451008} /* (26, 20, 21) {real, imag} */,
  {32'h3fb90996, 32'hbf814171} /* (26, 20, 20) {real, imag} */,
  {32'h3fb9002c, 32'h3ffd31c7} /* (26, 20, 19) {real, imag} */,
  {32'hbcd88128, 32'h4074a9b9} /* (26, 20, 18) {real, imag} */,
  {32'hc007ea2a, 32'h402f2f82} /* (26, 20, 17) {real, imag} */,
  {32'h3c44ca20, 32'hbf6a60c0} /* (26, 20, 16) {real, imag} */,
  {32'h40286915, 32'h3df96810} /* (26, 20, 15) {real, imag} */,
  {32'h3f88c29f, 32'h3e87e1ee} /* (26, 20, 14) {real, imag} */,
  {32'hbfa80fb0, 32'hbf438213} /* (26, 20, 13) {real, imag} */,
  {32'h3f12068a, 32'h3c2bd6c0} /* (26, 20, 12) {real, imag} */,
  {32'h3f01d76e, 32'hbf57eab2} /* (26, 20, 11) {real, imag} */,
  {32'hbf91a355, 32'hbf9092ff} /* (26, 20, 10) {real, imag} */,
  {32'h3f8f8344, 32'h3f28b93e} /* (26, 20, 9) {real, imag} */,
  {32'h3fb4f664, 32'h3f93cb3f} /* (26, 20, 8) {real, imag} */,
  {32'h3eaeec4c, 32'h3fcf5328} /* (26, 20, 7) {real, imag} */,
  {32'h4002c7fa, 32'hbe3cdfd0} /* (26, 20, 6) {real, imag} */,
  {32'h3f9b853e, 32'hbfd994f0} /* (26, 20, 5) {real, imag} */,
  {32'h402e3532, 32'hbe79cc90} /* (26, 20, 4) {real, imag} */,
  {32'h40381cae, 32'h3f4515e3} /* (26, 20, 3) {real, imag} */,
  {32'h3ff62b0a, 32'hbfe15cbc} /* (26, 20, 2) {real, imag} */,
  {32'hbf8d692d, 32'hbf5e750a} /* (26, 20, 1) {real, imag} */,
  {32'hbfc4a533, 32'h3e6713b3} /* (26, 20, 0) {real, imag} */,
  {32'hbdbda960, 32'h3dcbc080} /* (26, 19, 31) {real, imag} */,
  {32'hbdc01418, 32'hbf346124} /* (26, 19, 30) {real, imag} */,
  {32'h3f1a4bba, 32'hbf9cc31e} /* (26, 19, 29) {real, imag} */,
  {32'hbf3d13b9, 32'hbfebf3a6} /* (26, 19, 28) {real, imag} */,
  {32'hbf3c507d, 32'h3e7ede70} /* (26, 19, 27) {real, imag} */,
  {32'hbf1cee66, 32'hbf18681b} /* (26, 19, 26) {real, imag} */,
  {32'hc057da16, 32'hbe9c9db4} /* (26, 19, 25) {real, imag} */,
  {32'hc083b8b2, 32'h3e0c0bd8} /* (26, 19, 24) {real, imag} */,
  {32'hbe08f4e8, 32'hbf08ed3a} /* (26, 19, 23) {real, imag} */,
  {32'h3ef8bd92, 32'hbf2faae2} /* (26, 19, 22) {real, imag} */,
  {32'h3e98648e, 32'hbf0a85d7} /* (26, 19, 21) {real, imag} */,
  {32'h3fc89290, 32'h3faf6505} /* (26, 19, 20) {real, imag} */,
  {32'hbde60300, 32'h3fd81ac8} /* (26, 19, 19) {real, imag} */,
  {32'h3ee4d21c, 32'h40256536} /* (26, 19, 18) {real, imag} */,
  {32'h3d587a70, 32'h40886b42} /* (26, 19, 17) {real, imag} */,
  {32'hbd7b75e0, 32'h3f43cca7} /* (26, 19, 16) {real, imag} */,
  {32'h3f5997e4, 32'h3fb1cfe4} /* (26, 19, 15) {real, imag} */,
  {32'hc0042d35, 32'h3e2aaa00} /* (26, 19, 14) {real, imag} */,
  {32'hc010c0a1, 32'hbfe893be} /* (26, 19, 13) {real, imag} */,
  {32'hbe7eb91c, 32'hc008ad50} /* (26, 19, 12) {real, imag} */,
  {32'hbfa7b388, 32'hc0508f39} /* (26, 19, 11) {real, imag} */,
  {32'hbf8de790, 32'hc0644528} /* (26, 19, 10) {real, imag} */,
  {32'h40177949, 32'hbee6f1e8} /* (26, 19, 9) {real, imag} */,
  {32'h401465a3, 32'h3ff51f78} /* (26, 19, 8) {real, imag} */,
  {32'h3fdfe1f5, 32'h406cbf86} /* (26, 19, 7) {real, imag} */,
  {32'h402bb444, 32'h4038e3e4} /* (26, 19, 6) {real, imag} */,
  {32'h3ea9017e, 32'hbdd51a80} /* (26, 19, 5) {real, imag} */,
  {32'h3e87f780, 32'h3ffdb377} /* (26, 19, 4) {real, imag} */,
  {32'h4010cbd5, 32'h4046a437} /* (26, 19, 3) {real, imag} */,
  {32'h3f8d4f6f, 32'hbe11fc78} /* (26, 19, 2) {real, imag} */,
  {32'hbe326df8, 32'hbe7b6170} /* (26, 19, 1) {real, imag} */,
  {32'hbfb28940, 32'hbed6681a} /* (26, 19, 0) {real, imag} */,
  {32'h3f723f73, 32'h3f65ea5e} /* (26, 18, 31) {real, imag} */,
  {32'hbf7214c4, 32'h3e517aa0} /* (26, 18, 30) {real, imag} */,
  {32'hbf0507ee, 32'hbfbba18a} /* (26, 18, 29) {real, imag} */,
  {32'hbf8d6f09, 32'hbf86fa5c} /* (26, 18, 28) {real, imag} */,
  {32'h3f4875e6, 32'hbf9cb64e} /* (26, 18, 27) {real, imag} */,
  {32'h3f8c30e5, 32'hc019d864} /* (26, 18, 26) {real, imag} */,
  {32'hc01e5736, 32'hbfbacb79} /* (26, 18, 25) {real, imag} */,
  {32'hbfc906d8, 32'hc04168cb} /* (26, 18, 24) {real, imag} */,
  {32'h40261ec0, 32'hbfccd071} /* (26, 18, 23) {real, imag} */,
  {32'h3f04fe0a, 32'hbff1e895} /* (26, 18, 22) {real, imag} */,
  {32'hbf4875cf, 32'hc08095ce} /* (26, 18, 21) {real, imag} */,
  {32'h400dabd0, 32'hc0033dd7} /* (26, 18, 20) {real, imag} */,
  {32'hbd575fb0, 32'hbfe7c308} /* (26, 18, 19) {real, imag} */,
  {32'h3e8081c3, 32'h3f6fa56f} /* (26, 18, 18) {real, imag} */,
  {32'h3f1e88fe, 32'h4060d21c} /* (26, 18, 17) {real, imag} */,
  {32'hc01ab4ea, 32'h4014bc3e} /* (26, 18, 16) {real, imag} */,
  {32'hbea2eff0, 32'h3ffdc744} /* (26, 18, 15) {real, imag} */,
  {32'hbfa80ca8, 32'h3fb32e29} /* (26, 18, 14) {real, imag} */,
  {32'hbf71686a, 32'hbf541f1a} /* (26, 18, 13) {real, imag} */,
  {32'h3edc7be6, 32'hc04d6b8e} /* (26, 18, 12) {real, imag} */,
  {32'h3e5adc18, 32'hc0597d3c} /* (26, 18, 11) {real, imag} */,
  {32'h3ea8b47a, 32'hbe6293b8} /* (26, 18, 10) {real, imag} */,
  {32'h3f9fc2d0, 32'h3ffd3e8a} /* (26, 18, 9) {real, imag} */,
  {32'h3f1bf54c, 32'h40456718} /* (26, 18, 8) {real, imag} */,
  {32'hbf82d8d0, 32'h40852c60} /* (26, 18, 7) {real, imag} */,
  {32'h3f7c5894, 32'h3ed022c0} /* (26, 18, 6) {real, imag} */,
  {32'h3fa0479e, 32'hc037ed97} /* (26, 18, 5) {real, imag} */,
  {32'h3fe81c7a, 32'hbfeaa674} /* (26, 18, 4) {real, imag} */,
  {32'h4026e9ac, 32'h3b82b200} /* (26, 18, 3) {real, imag} */,
  {32'h400fbf03, 32'hbee00da6} /* (26, 18, 2) {real, imag} */,
  {32'h40688041, 32'h3e730350} /* (26, 18, 1) {real, imag} */,
  {32'h3f42e974, 32'hbd446fa0} /* (26, 18, 0) {real, imag} */,
  {32'h3fc2240c, 32'h40102ae7} /* (26, 17, 31) {real, imag} */,
  {32'h400c5854, 32'h3eeca2e8} /* (26, 17, 30) {real, imag} */,
  {32'h3f3f7755, 32'hbfc085b0} /* (26, 17, 29) {real, imag} */,
  {32'h3f470846, 32'hbfe61771} /* (26, 17, 28) {real, imag} */,
  {32'h3f30f11e, 32'hc0347fb7} /* (26, 17, 27) {real, imag} */,
  {32'h3faa0660, 32'hc0873c6b} /* (26, 17, 26) {real, imag} */,
  {32'h3f520e4e, 32'hc028688c} /* (26, 17, 25) {real, imag} */,
  {32'h403922a3, 32'hc021927a} /* (26, 17, 24) {real, imag} */,
  {32'h402a8c96, 32'hbf34eb88} /* (26, 17, 23) {real, imag} */,
  {32'h3fc0e128, 32'h3e8f4d1e} /* (26, 17, 22) {real, imag} */,
  {32'hbe7845d4, 32'hc00f4b70} /* (26, 17, 21) {real, imag} */,
  {32'h3ff62f60, 32'hc04953f4} /* (26, 17, 20) {real, imag} */,
  {32'h3f55183a, 32'hc009da60} /* (26, 17, 19) {real, imag} */,
  {32'h3f2b530c, 32'hbfc0023a} /* (26, 17, 18) {real, imag} */,
  {32'h3f31b71a, 32'hbf75c74e} /* (26, 17, 17) {real, imag} */,
  {32'h3f3bbf84, 32'h3fc1ecec} /* (26, 17, 16) {real, imag} */,
  {32'h3f3e83ec, 32'h4037edf3} /* (26, 17, 15) {real, imag} */,
  {32'h3f55d8e6, 32'h3ffe83e2} /* (26, 17, 14) {real, imag} */,
  {32'h3e97f5ee, 32'hbe049674} /* (26, 17, 13) {real, imag} */,
  {32'h3ed55ab0, 32'hbfea6098} /* (26, 17, 12) {real, imag} */,
  {32'h3f8aa296, 32'hbf84e4fc} /* (26, 17, 11) {real, imag} */,
  {32'h3fb20069, 32'h40232005} /* (26, 17, 10) {real, imag} */,
  {32'h400078c0, 32'h40a32772} /* (26, 17, 9) {real, imag} */,
  {32'h4056ec0b, 32'h406cb6d9} /* (26, 17, 8) {real, imag} */,
  {32'hbde8ddd0, 32'h3e106e20} /* (26, 17, 7) {real, imag} */,
  {32'hbefbf430, 32'h3d34b8e0} /* (26, 17, 6) {real, imag} */,
  {32'h3fc4cb26, 32'hbfb2df84} /* (26, 17, 5) {real, imag} */,
  {32'h3fcfd877, 32'hc086b098} /* (26, 17, 4) {real, imag} */,
  {32'h3f2e46c4, 32'hc0743790} /* (26, 17, 3) {real, imag} */,
  {32'h3ecce480, 32'hbf55265a} /* (26, 17, 2) {real, imag} */,
  {32'h4051a6d2, 32'h3f4119b6} /* (26, 17, 1) {real, imag} */,
  {32'h3de14d30, 32'h400b9a04} /* (26, 17, 0) {real, imag} */,
  {32'hbef15470, 32'h3cd7cc60} /* (26, 16, 31) {real, imag} */,
  {32'h3e2120dc, 32'hbcb90a00} /* (26, 16, 30) {real, imag} */,
  {32'h3eb91d34, 32'hbe289054} /* (26, 16, 29) {real, imag} */,
  {32'h3fdc3677, 32'hc0412236} /* (26, 16, 28) {real, imag} */,
  {32'h3f22233e, 32'hbf81f9c8} /* (26, 16, 27) {real, imag} */,
  {32'hbe95fa2c, 32'hbfc3fa93} /* (26, 16, 26) {real, imag} */,
  {32'hbe950a68, 32'hc02e5dbf} /* (26, 16, 25) {real, imag} */,
  {32'h3fc42384, 32'hbf3f8d76} /* (26, 16, 24) {real, imag} */,
  {32'h401aeb7a, 32'h3f926868} /* (26, 16, 23) {real, imag} */,
  {32'h4013f1a2, 32'h400638d2} /* (26, 16, 22) {real, imag} */,
  {32'h3efbe088, 32'hbedc513a} /* (26, 16, 21) {real, imag} */,
  {32'h3fea5019, 32'hbf9d4d94} /* (26, 16, 20) {real, imag} */,
  {32'h3f8fea62, 32'hbfec0b9f} /* (26, 16, 19) {real, imag} */,
  {32'hbe62d538, 32'hc01ff778} /* (26, 16, 18) {real, imag} */,
  {32'hbfeb9283, 32'hbf26cc5c} /* (26, 16, 17) {real, imag} */,
  {32'hbe8b2cc8, 32'h3fa8badd} /* (26, 16, 16) {real, imag} */,
  {32'hbf49fa8a, 32'h3ffa8579} /* (26, 16, 15) {real, imag} */,
  {32'h3e1c26f8, 32'h3f99db78} /* (26, 16, 14) {real, imag} */,
  {32'h3f5c0ef2, 32'h3eb13ae4} /* (26, 16, 13) {real, imag} */,
  {32'hbed3fe58, 32'hbf855f2b} /* (26, 16, 12) {real, imag} */,
  {32'hbe97423a, 32'h3f9fc6fc} /* (26, 16, 11) {real, imag} */,
  {32'hbf1297e5, 32'h403454ac} /* (26, 16, 10) {real, imag} */,
  {32'h3e4752c0, 32'h407d2a15} /* (26, 16, 9) {real, imag} */,
  {32'h3f205c10, 32'h3fd5f677} /* (26, 16, 8) {real, imag} */,
  {32'hbf6ce1a4, 32'hbfd176a6} /* (26, 16, 7) {real, imag} */,
  {32'h3f38048e, 32'hbffd9283} /* (26, 16, 6) {real, imag} */,
  {32'h3fb8cdec, 32'hbfbe0411} /* (26, 16, 5) {real, imag} */,
  {32'h3e732fe0, 32'hc041aed2} /* (26, 16, 4) {real, imag} */,
  {32'hbfc4b3ca, 32'hc02cd37a} /* (26, 16, 3) {real, imag} */,
  {32'hbfd8c784, 32'hbea719ec} /* (26, 16, 2) {real, imag} */,
  {32'h3ebd0898, 32'hbf8ae200} /* (26, 16, 1) {real, imag} */,
  {32'hbf6b9bb0, 32'hbfdef3bc} /* (26, 16, 0) {real, imag} */,
  {32'hbebb5991, 32'hbf3536a1} /* (26, 15, 31) {real, imag} */,
  {32'h3e3ff114, 32'h3eb0c0b8} /* (26, 15, 30) {real, imag} */,
  {32'h3fdc7953, 32'h3f303ee1} /* (26, 15, 29) {real, imag} */,
  {32'h3f986494, 32'hc04de3e4} /* (26, 15, 28) {real, imag} */,
  {32'hbf1e444e, 32'hbe206480} /* (26, 15, 27) {real, imag} */,
  {32'hbfe5ea31, 32'hbe481188} /* (26, 15, 26) {real, imag} */,
  {32'hbfa49401, 32'hc011074a} /* (26, 15, 25) {real, imag} */,
  {32'hbfe1d576, 32'hbfc1b99e} /* (26, 15, 24) {real, imag} */,
  {32'hbd4e5b60, 32'hbfb8b388} /* (26, 15, 23) {real, imag} */,
  {32'hbf0f2f06, 32'hbf100b50} /* (26, 15, 22) {real, imag} */,
  {32'hbecc3416, 32'hbf6d28fe} /* (26, 15, 21) {real, imag} */,
  {32'h3ec890db, 32'h3f15dffe} /* (26, 15, 20) {real, imag} */,
  {32'h3f874163, 32'h3e32c9fc} /* (26, 15, 19) {real, imag} */,
  {32'hbecde4c4, 32'hbfeffc10} /* (26, 15, 18) {real, imag} */,
  {32'hbff0cad2, 32'h3d9654c0} /* (26, 15, 17) {real, imag} */,
  {32'hbf6e8787, 32'h3ee91260} /* (26, 15, 16) {real, imag} */,
  {32'hbfdecd56, 32'h402bdbfc} /* (26, 15, 15) {real, imag} */,
  {32'hbfa71072, 32'h3f88650b} /* (26, 15, 14) {real, imag} */,
  {32'hc00639da, 32'h3f7c2515} /* (26, 15, 13) {real, imag} */,
  {32'hc0571beb, 32'hbf3c2b38} /* (26, 15, 12) {real, imag} */,
  {32'hbfc9e875, 32'hbee9a57c} /* (26, 15, 11) {real, imag} */,
  {32'hbfd84718, 32'h3fd7fedd} /* (26, 15, 10) {real, imag} */,
  {32'hbf104042, 32'h3fcf5ac0} /* (26, 15, 9) {real, imag} */,
  {32'hbfe6cda7, 32'h3fb11aae} /* (26, 15, 8) {real, imag} */,
  {32'hbf5f657c, 32'hbf2962a8} /* (26, 15, 7) {real, imag} */,
  {32'h3fddcf3a, 32'hbf573d76} /* (26, 15, 6) {real, imag} */,
  {32'h3f2a46ac, 32'h3ef03bac} /* (26, 15, 5) {real, imag} */,
  {32'h3e5f638c, 32'h3f424f08} /* (26, 15, 4) {real, imag} */,
  {32'hbfaf0036, 32'h3cfbe5c0} /* (26, 15, 3) {real, imag} */,
  {32'hbf881f37, 32'h3f52df08} /* (26, 15, 2) {real, imag} */,
  {32'h3f02a8f0, 32'hbfde1d3d} /* (26, 15, 1) {real, imag} */,
  {32'hbf235db0, 32'hbff37094} /* (26, 15, 0) {real, imag} */,
  {32'hbf4612dc, 32'h3d1a5400} /* (26, 14, 31) {real, imag} */,
  {32'hbee814a0, 32'h3ff5dd15} /* (26, 14, 30) {real, imag} */,
  {32'h3f057b54, 32'h40298865} /* (26, 14, 29) {real, imag} */,
  {32'hbfd2637a, 32'hbe77e5b8} /* (26, 14, 28) {real, imag} */,
  {32'h3d98d1f0, 32'h3ed1b35c} /* (26, 14, 27) {real, imag} */,
  {32'hbfa98e4d, 32'h3f05a485} /* (26, 14, 26) {real, imag} */,
  {32'hbffc6df6, 32'h3f106053} /* (26, 14, 25) {real, imag} */,
  {32'hc04b3c62, 32'hbfae8ec2} /* (26, 14, 24) {real, imag} */,
  {32'hc024147a, 32'hbff08563} /* (26, 14, 23) {real, imag} */,
  {32'hc0008dc8, 32'hbd1dcb20} /* (26, 14, 22) {real, imag} */,
  {32'hc05c79f0, 32'hbe73f9f4} /* (26, 14, 21) {real, imag} */,
  {32'hbfa892ce, 32'h3f18d173} /* (26, 14, 20) {real, imag} */,
  {32'h3fa57250, 32'hbf946862} /* (26, 14, 19) {real, imag} */,
  {32'h3fba5690, 32'hc00b3169} /* (26, 14, 18) {real, imag} */,
  {32'hbd29d3d0, 32'hbd613e20} /* (26, 14, 17) {real, imag} */,
  {32'h3f25b88e, 32'h3ffcc9ea} /* (26, 14, 16) {real, imag} */,
  {32'h3dd180e8, 32'h403cec38} /* (26, 14, 15) {real, imag} */,
  {32'h3f3a9d08, 32'h3e116404} /* (26, 14, 14) {real, imag} */,
  {32'hbf9de086, 32'h3e83af60} /* (26, 14, 13) {real, imag} */,
  {32'hbfc0437d, 32'h3eddbc50} /* (26, 14, 12) {real, imag} */,
  {32'hbfc3542a, 32'hbebcc6a8} /* (26, 14, 11) {real, imag} */,
  {32'hc005c333, 32'h3fbb53bb} /* (26, 14, 10) {real, imag} */,
  {32'hbf6f6d96, 32'h3f80abef} /* (26, 14, 9) {real, imag} */,
  {32'hbf64a192, 32'h3e8b4c2c} /* (26, 14, 8) {real, imag} */,
  {32'hbe57f1ec, 32'hc01a9fb0} /* (26, 14, 7) {real, imag} */,
  {32'hbeede1a4, 32'hbf953806} /* (26, 14, 6) {real, imag} */,
  {32'h3e31ebc9, 32'h3f4ecc3a} /* (26, 14, 5) {real, imag} */,
  {32'h3f88cf29, 32'h3f692aac} /* (26, 14, 4) {real, imag} */,
  {32'h3eed582e, 32'h3fa6d66a} /* (26, 14, 3) {real, imag} */,
  {32'hbf40f5a4, 32'h3f7ee122} /* (26, 14, 2) {real, imag} */,
  {32'h3d098880, 32'hc020a262} /* (26, 14, 1) {real, imag} */,
  {32'h3e9a6f5e, 32'hbf04e4b8} /* (26, 14, 0) {real, imag} */,
  {32'hbf8c238e, 32'hbf41ba8f} /* (26, 13, 31) {real, imag} */,
  {32'hc0117cf7, 32'hbf1d62fc} /* (26, 13, 30) {real, imag} */,
  {32'hbf4e4235, 32'h3f78f3e6} /* (26, 13, 29) {real, imag} */,
  {32'hbfb18f64, 32'hbf78aae6} /* (26, 13, 28) {real, imag} */,
  {32'h40145366, 32'hbfe58ff4} /* (26, 13, 27) {real, imag} */,
  {32'h3f8f172e, 32'h3f77ffee} /* (26, 13, 26) {real, imag} */,
  {32'hbfd5a220, 32'h3f1a44f9} /* (26, 13, 25) {real, imag} */,
  {32'hc03b12b6, 32'hbef1a8f0} /* (26, 13, 24) {real, imag} */,
  {32'hc06d2ba5, 32'h3ed5317c} /* (26, 13, 23) {real, imag} */,
  {32'h3e50df10, 32'h3ee6563c} /* (26, 13, 22) {real, imag} */,
  {32'hbff2f282, 32'hbeb25c32} /* (26, 13, 21) {real, imag} */,
  {32'hc0304186, 32'h3f4e3752} /* (26, 13, 20) {real, imag} */,
  {32'hc016563b, 32'hbf8846ec} /* (26, 13, 19) {real, imag} */,
  {32'hbf856847, 32'hbf1cf69f} /* (26, 13, 18) {real, imag} */,
  {32'h3f711f90, 32'h3ea647e0} /* (26, 13, 17) {real, imag} */,
  {32'h3f0a39c3, 32'h3f129d94} /* (26, 13, 16) {real, imag} */,
  {32'h3de2fba8, 32'h400f6adb} /* (26, 13, 15) {real, imag} */,
  {32'h3faa10bc, 32'h3fe9ba2e} /* (26, 13, 14) {real, imag} */,
  {32'h3fadecde, 32'h3f6f084e} /* (26, 13, 13) {real, imag} */,
  {32'hbf84ece2, 32'h3e683898} /* (26, 13, 12) {real, imag} */,
  {32'hc02eab8e, 32'h3e09a6a8} /* (26, 13, 11) {real, imag} */,
  {32'hc00871c7, 32'hbf13d2d2} /* (26, 13, 10) {real, imag} */,
  {32'h3e648530, 32'hbf5a982a} /* (26, 13, 9) {real, imag} */,
  {32'h3fd16e6a, 32'h40290810} /* (26, 13, 8) {real, imag} */,
  {32'hbe4f2698, 32'h4026ccf6} /* (26, 13, 7) {real, imag} */,
  {32'hc00b554e, 32'h3fae5513} /* (26, 13, 6) {real, imag} */,
  {32'h3f30d40a, 32'h3f7e74ff} /* (26, 13, 5) {real, imag} */,
  {32'h4011847f, 32'hbe97f093} /* (26, 13, 4) {real, imag} */,
  {32'h3f8c689e, 32'h3f4dab68} /* (26, 13, 3) {real, imag} */,
  {32'h3fb7f518, 32'hbfe2fefe} /* (26, 13, 2) {real, imag} */,
  {32'h3f710ec0, 32'hbff6715b} /* (26, 13, 1) {real, imag} */,
  {32'h3e16aa00, 32'h3f45236d} /* (26, 13, 0) {real, imag} */,
  {32'hbf98d850, 32'h3f1d2216} /* (26, 12, 31) {real, imag} */,
  {32'hc00bd6de, 32'hbf4e3eeb} /* (26, 12, 30) {real, imag} */,
  {32'h3f3af68c, 32'h3df4af68} /* (26, 12, 29) {real, imag} */,
  {32'h40298b25, 32'hbff672da} /* (26, 12, 28) {real, imag} */,
  {32'h404c19da, 32'hbfd28e1e} /* (26, 12, 27) {real, imag} */,
  {32'h3d794710, 32'h3f75857a} /* (26, 12, 26) {real, imag} */,
  {32'hbeca6734, 32'hbeb432a8} /* (26, 12, 25) {real, imag} */,
  {32'hbf1888b4, 32'hbe03a8d0} /* (26, 12, 24) {real, imag} */,
  {32'hbfd8b7d2, 32'h4013912e} /* (26, 12, 23) {real, imag} */,
  {32'h3f0bc792, 32'h400be16c} /* (26, 12, 22) {real, imag} */,
  {32'h3f17abd2, 32'hbf5350c1} /* (26, 12, 21) {real, imag} */,
  {32'hc02014a8, 32'hbebb172c} /* (26, 12, 20) {real, imag} */,
  {32'hc0a29628, 32'hbfc735c6} /* (26, 12, 19) {real, imag} */,
  {32'hbf3b67f3, 32'h3edfaa44} /* (26, 12, 18) {real, imag} */,
  {32'h404df554, 32'hbf8e3955} /* (26, 12, 17) {real, imag} */,
  {32'h3ffadaf7, 32'hc02700dd} /* (26, 12, 16) {real, imag} */,
  {32'h3f9f7783, 32'h3efb23de} /* (26, 12, 15) {real, imag} */,
  {32'h3f9ec309, 32'h402106f4} /* (26, 12, 14) {real, imag} */,
  {32'h401d6497, 32'h3fc6fe88} /* (26, 12, 13) {real, imag} */,
  {32'h3f3f1554, 32'hc01aa1da} /* (26, 12, 12) {real, imag} */,
  {32'hbf74aaec, 32'hc0145e37} /* (26, 12, 11) {real, imag} */,
  {32'hbf5052da, 32'hbfdc2cec} /* (26, 12, 10) {real, imag} */,
  {32'h3d387b90, 32'hbf6b74aa} /* (26, 12, 9) {real, imag} */,
  {32'hbf9d9f8b, 32'h40208e13} /* (26, 12, 8) {real, imag} */,
  {32'hbf27590a, 32'h3ffe63ec} /* (26, 12, 7) {real, imag} */,
  {32'hbfd58922, 32'hbe492c94} /* (26, 12, 6) {real, imag} */,
  {32'h3e3b67c8, 32'hbcf7d700} /* (26, 12, 5) {real, imag} */,
  {32'h3f920dac, 32'h3e2bf854} /* (26, 12, 4) {real, imag} */,
  {32'h3cd55a60, 32'h3fcc4157} /* (26, 12, 3) {real, imag} */,
  {32'h3fe61dfd, 32'hbfb1ac14} /* (26, 12, 2) {real, imag} */,
  {32'h3f2d5014, 32'hbf86bcfa} /* (26, 12, 1) {real, imag} */,
  {32'hbea7d01c, 32'h3fa40d82} /* (26, 12, 0) {real, imag} */,
  {32'hbf156432, 32'hbfa1f1ca} /* (26, 11, 31) {real, imag} */,
  {32'hbf730a94, 32'hc00f755e} /* (26, 11, 30) {real, imag} */,
  {32'h3e5f4324, 32'h3f7cc184} /* (26, 11, 29) {real, imag} */,
  {32'h3fc7e691, 32'h3db5a010} /* (26, 11, 28) {real, imag} */,
  {32'h3fea9341, 32'hbf9a0e4b} /* (26, 11, 27) {real, imag} */,
  {32'h3e08530e, 32'hbec2453e} /* (26, 11, 26) {real, imag} */,
  {32'hbf2fad8f, 32'h3e5f7738} /* (26, 11, 25) {real, imag} */,
  {32'hbcf701e0, 32'hbe54a9a0} /* (26, 11, 24) {real, imag} */,
  {32'hbf1d916c, 32'h3f309454} /* (26, 11, 23) {real, imag} */,
  {32'h3e55ff88, 32'hbf032c19} /* (26, 11, 22) {real, imag} */,
  {32'h40145a68, 32'hbf22c028} /* (26, 11, 21) {real, imag} */,
  {32'h40097c14, 32'hc011bbf2} /* (26, 11, 20) {real, imag} */,
  {32'h3e9543f9, 32'hbfd2082b} /* (26, 11, 19) {real, imag} */,
  {32'h3ff886a8, 32'h3f800e07} /* (26, 11, 18) {real, imag} */,
  {32'h3fa2ec10, 32'hbfb88038} /* (26, 11, 17) {real, imag} */,
  {32'h3ed813c8, 32'hc099278b} /* (26, 11, 16) {real, imag} */,
  {32'h3fd84c51, 32'hc02fd49f} /* (26, 11, 15) {real, imag} */,
  {32'h40213a92, 32'hbecf921a} /* (26, 11, 14) {real, imag} */,
  {32'h3f93862a, 32'h3fbeee44} /* (26, 11, 13) {real, imag} */,
  {32'h3f198fd4, 32'hbffddcad} /* (26, 11, 12) {real, imag} */,
  {32'hbed3199e, 32'hc06dc2af} /* (26, 11, 11) {real, imag} */,
  {32'h3f1cabfd, 32'hc076594c} /* (26, 11, 10) {real, imag} */,
  {32'h3f033fdd, 32'hc01a340d} /* (26, 11, 9) {real, imag} */,
  {32'hbd729520, 32'hbc2f5940} /* (26, 11, 8) {real, imag} */,
  {32'hbdaba424, 32'hc00ab998} /* (26, 11, 7) {real, imag} */,
  {32'h3f2cbc96, 32'hc0643945} /* (26, 11, 6) {real, imag} */,
  {32'h3fdf6a1e, 32'hbfb86f6a} /* (26, 11, 5) {real, imag} */,
  {32'hbeaea53a, 32'h3cc15460} /* (26, 11, 4) {real, imag} */,
  {32'hbfc45519, 32'hbd997538} /* (26, 11, 3) {real, imag} */,
  {32'hbf1387c9, 32'hbfd5f21e} /* (26, 11, 2) {real, imag} */,
  {32'h402ed45e, 32'hbff51aa9} /* (26, 11, 1) {real, imag} */,
  {32'h4016cc51, 32'hbfa87d8b} /* (26, 11, 0) {real, imag} */,
  {32'hbebd7422, 32'hbfd3b4f3} /* (26, 10, 31) {real, imag} */,
  {32'h3f1d7750, 32'hc040f412} /* (26, 10, 30) {real, imag} */,
  {32'hbf619e12, 32'hbfd9ea17} /* (26, 10, 29) {real, imag} */,
  {32'hbf5d6b78, 32'h4018bc7d} /* (26, 10, 28) {real, imag} */,
  {32'hbff688f8, 32'h400d097a} /* (26, 10, 27) {real, imag} */,
  {32'h3f8a6039, 32'hbf0fddf3} /* (26, 10, 26) {real, imag} */,
  {32'h3efbfc46, 32'h3fef834e} /* (26, 10, 25) {real, imag} */,
  {32'h3fae1ce2, 32'h40542866} /* (26, 10, 24) {real, imag} */,
  {32'h4010eb29, 32'h3f9fb11a} /* (26, 10, 23) {real, imag} */,
  {32'h3fda16c6, 32'hbe9391fc} /* (26, 10, 22) {real, imag} */,
  {32'h3fa71975, 32'hbe79cae6} /* (26, 10, 21) {real, imag} */,
  {32'h405f24dc, 32'hc046ab84} /* (26, 10, 20) {real, imag} */,
  {32'h3f6ebc98, 32'hbfe45e6e} /* (26, 10, 19) {real, imag} */,
  {32'h3f06458c, 32'h3f18abd6} /* (26, 10, 18) {real, imag} */,
  {32'hbfd310dd, 32'hc029460c} /* (26, 10, 17) {real, imag} */,
  {32'hbf03d07e, 32'hc0852fe9} /* (26, 10, 16) {real, imag} */,
  {32'hbe3b5fbc, 32'hbdb16398} /* (26, 10, 15) {real, imag} */,
  {32'h3e3fd894, 32'h3faa664c} /* (26, 10, 14) {real, imag} */,
  {32'h3e38d43c, 32'h40715d70} /* (26, 10, 13) {real, imag} */,
  {32'hbe61e768, 32'hbd906828} /* (26, 10, 12) {real, imag} */,
  {32'hbfd9d8c7, 32'hc06082df} /* (26, 10, 11) {real, imag} */,
  {32'hbf7e6357, 32'hc0009dfa} /* (26, 10, 10) {real, imag} */,
  {32'h3f169b92, 32'hbd37d300} /* (26, 10, 9) {real, imag} */,
  {32'h40149d06, 32'h3e087335} /* (26, 10, 8) {real, imag} */,
  {32'h4005ce0c, 32'hc01b56da} /* (26, 10, 7) {real, imag} */,
  {32'h4062d1a6, 32'hbfe816f9} /* (26, 10, 6) {real, imag} */,
  {32'h3fcebddd, 32'hbf69ce9d} /* (26, 10, 5) {real, imag} */,
  {32'h3f0f9237, 32'hbfbf86b2} /* (26, 10, 4) {real, imag} */,
  {32'h3c790d40, 32'hbfb817ce} /* (26, 10, 3) {real, imag} */,
  {32'hbfbcbbfe, 32'hbfef2718} /* (26, 10, 2) {real, imag} */,
  {32'h402f6d06, 32'hbfa37415} /* (26, 10, 1) {real, imag} */,
  {32'h401c590b, 32'hbedd3bae} /* (26, 10, 0) {real, imag} */,
  {32'h3f83aba3, 32'hbf1211b0} /* (26, 9, 31) {real, imag} */,
  {32'h3f6097b5, 32'hbfb01ada} /* (26, 9, 30) {real, imag} */,
  {32'hbf3135e8, 32'hbf0e36da} /* (26, 9, 29) {real, imag} */,
  {32'h3f88d3c6, 32'h3eefd6dc} /* (26, 9, 28) {real, imag} */,
  {32'h3ea702aa, 32'h3f4c9939} /* (26, 9, 27) {real, imag} */,
  {32'h40045dd4, 32'hbf5855a1} /* (26, 9, 26) {real, imag} */,
  {32'h3f37cf57, 32'h3f4fe79b} /* (26, 9, 25) {real, imag} */,
  {32'h3f045818, 32'h3faa83bc} /* (26, 9, 24) {real, imag} */,
  {32'h400a0b5b, 32'h40079cd3} /* (26, 9, 23) {real, imag} */,
  {32'h3fab7c5b, 32'h3efbe81c} /* (26, 9, 22) {real, imag} */,
  {32'hbe8be266, 32'hbe46e948} /* (26, 9, 21) {real, imag} */,
  {32'h3f896ad5, 32'hc047d9be} /* (26, 9, 20) {real, imag} */,
  {32'hbece811a, 32'hbf6621e2} /* (26, 9, 19) {real, imag} */,
  {32'h3f3fb592, 32'h3ecbc87a} /* (26, 9, 18) {real, imag} */,
  {32'hbee08e12, 32'hc0133b4c} /* (26, 9, 17) {real, imag} */,
  {32'h3f13c444, 32'hbff87a87} /* (26, 9, 16) {real, imag} */,
  {32'hbf29f3f6, 32'h3ffc2c4c} /* (26, 9, 15) {real, imag} */,
  {32'h3ed46814, 32'h3f87a1c6} /* (26, 9, 14) {real, imag} */,
  {32'h3f8d276a, 32'h3fe72e0e} /* (26, 9, 13) {real, imag} */,
  {32'hbd481510, 32'h3d736e40} /* (26, 9, 12) {real, imag} */,
  {32'h3e39b4d8, 32'hbf94df86} /* (26, 9, 11) {real, imag} */,
  {32'h3f675ef4, 32'hbe0203f8} /* (26, 9, 10) {real, imag} */,
  {32'h4022b74b, 32'h3f8f4f7a} /* (26, 9, 9) {real, imag} */,
  {32'h3fe6e470, 32'h40015910} /* (26, 9, 8) {real, imag} */,
  {32'h3ef6b904, 32'hbddbf420} /* (26, 9, 7) {real, imag} */,
  {32'h401d1794, 32'hbfa2ad8a} /* (26, 9, 6) {real, imag} */,
  {32'hc0030a2c, 32'hc02b3e4c} /* (26, 9, 5) {real, imag} */,
  {32'hbf19b191, 32'hc03312ba} /* (26, 9, 4) {real, imag} */,
  {32'h3fae010e, 32'hc0192fa0} /* (26, 9, 3) {real, imag} */,
  {32'hbed27235, 32'hc003c0e5} /* (26, 9, 2) {real, imag} */,
  {32'h3f1698e3, 32'hbf1de93c} /* (26, 9, 1) {real, imag} */,
  {32'h3e1ed1b4, 32'h3e9e3398} /* (26, 9, 0) {real, imag} */,
  {32'hbf1b1690, 32'hbf5cd652} /* (26, 8, 31) {real, imag} */,
  {32'hbe03dfa8, 32'hbfaea5e2} /* (26, 8, 30) {real, imag} */,
  {32'h3fad3ea0, 32'hbe029ae0} /* (26, 8, 29) {real, imag} */,
  {32'h402ade29, 32'hbf013056} /* (26, 8, 28) {real, imag} */,
  {32'h40775728, 32'hbfe1f80e} /* (26, 8, 27) {real, imag} */,
  {32'h3ff45410, 32'hbe3765b8} /* (26, 8, 26) {real, imag} */,
  {32'hbf3de9e1, 32'hbef0f164} /* (26, 8, 25) {real, imag} */,
  {32'hbfc7fede, 32'hbfa009e6} /* (26, 8, 24) {real, imag} */,
  {32'hbf235f38, 32'hbde01fa0} /* (26, 8, 23) {real, imag} */,
  {32'hbe254424, 32'h3fc25a36} /* (26, 8, 22) {real, imag} */,
  {32'h3cb10fe0, 32'h3f6acea6} /* (26, 8, 21) {real, imag} */,
  {32'h3f1ca228, 32'hbf9681fa} /* (26, 8, 20) {real, imag} */,
  {32'h3fa084e0, 32'hc017cdfc} /* (26, 8, 19) {real, imag} */,
  {32'h3d99d4a0, 32'hbfd4bf9c} /* (26, 8, 18) {real, imag} */,
  {32'h3f5d4aa1, 32'hbf89f81c} /* (26, 8, 17) {real, imag} */,
  {32'h3e470408, 32'h3dafee50} /* (26, 8, 16) {real, imag} */,
  {32'hbe02ea40, 32'hbfc12ba6} /* (26, 8, 15) {real, imag} */,
  {32'h4051da5f, 32'hbdfba548} /* (26, 8, 14) {real, imag} */,
  {32'h3faf90ee, 32'h3ff9c3ce} /* (26, 8, 13) {real, imag} */,
  {32'hbf938f3c, 32'h4060e6e2} /* (26, 8, 12) {real, imag} */,
  {32'hbd9836e8, 32'h3f62b63f} /* (26, 8, 11) {real, imag} */,
  {32'h3f9959f8, 32'hbeb1fb2c} /* (26, 8, 10) {real, imag} */,
  {32'h401332a2, 32'hbff8292a} /* (26, 8, 9) {real, imag} */,
  {32'h40599234, 32'hbea2ebce} /* (26, 8, 8) {real, imag} */,
  {32'h4050c55e, 32'hc00cc6b5} /* (26, 8, 7) {real, imag} */,
  {32'h3ff3afe7, 32'hc0456b71} /* (26, 8, 6) {real, imag} */,
  {32'hc0132a50, 32'hc02f039b} /* (26, 8, 5) {real, imag} */,
  {32'hbf9d104b, 32'hc00babbc} /* (26, 8, 4) {real, imag} */,
  {32'h3fdc1c36, 32'hbffdcfa2} /* (26, 8, 3) {real, imag} */,
  {32'hbfa0441a, 32'hc0013b4c} /* (26, 8, 2) {real, imag} */,
  {32'hbf532533, 32'h3f8884e0} /* (26, 8, 1) {real, imag} */,
  {32'h3edadfa6, 32'h3fe2120e} /* (26, 8, 0) {real, imag} */,
  {32'h3e837eec, 32'hbfc62576} /* (26, 7, 31) {real, imag} */,
  {32'hbfa580f0, 32'hbf174018} /* (26, 7, 30) {real, imag} */,
  {32'h3d2a73c0, 32'hbf5f960a} /* (26, 7, 29) {real, imag} */,
  {32'h3fc79dd7, 32'hbf5aafdf} /* (26, 7, 28) {real, imag} */,
  {32'h4047c7cc, 32'hbf2ebbbf} /* (26, 7, 27) {real, imag} */,
  {32'h4006dc46, 32'hbf836e04} /* (26, 7, 26) {real, imag} */,
  {32'hbdcd92c0, 32'hbf8f14aa} /* (26, 7, 25) {real, imag} */,
  {32'h3c8aba40, 32'h3ed7eabc} /* (26, 7, 24) {real, imag} */,
  {32'h3d9928d0, 32'hc02c4c39} /* (26, 7, 23) {real, imag} */,
  {32'hbe476a28, 32'hbefd85f4} /* (26, 7, 22) {real, imag} */,
  {32'h3ff948b8, 32'h3ff895dd} /* (26, 7, 21) {real, imag} */,
  {32'h3fcd29c0, 32'h3e615e9c} /* (26, 7, 20) {real, imag} */,
  {32'h40368d35, 32'hc08ebf56} /* (26, 7, 19) {real, imag} */,
  {32'h3f94300c, 32'hbfefa77a} /* (26, 7, 18) {real, imag} */,
  {32'h3e582b90, 32'hbf258b34} /* (26, 7, 17) {real, imag} */,
  {32'hbf16097a, 32'hbf874f29} /* (26, 7, 16) {real, imag} */,
  {32'hbf19b58c, 32'hc0220a82} /* (26, 7, 15) {real, imag} */,
  {32'h3fdcfbd4, 32'hbf9e0cea} /* (26, 7, 14) {real, imag} */,
  {32'h3fe10bbc, 32'h3f56490e} /* (26, 7, 13) {real, imag} */,
  {32'h3ebbaa9a, 32'h3f9aaa9d} /* (26, 7, 12) {real, imag} */,
  {32'h3fac9a57, 32'h3eaa5ed2} /* (26, 7, 11) {real, imag} */,
  {32'hbd916cf0, 32'hc0286dfb} /* (26, 7, 10) {real, imag} */,
  {32'h3ea13420, 32'hc0852c73} /* (26, 7, 9) {real, imag} */,
  {32'h3fb2aeca, 32'hbf9a2e31} /* (26, 7, 8) {real, imag} */,
  {32'h4023e852, 32'hc05a5a93} /* (26, 7, 7) {real, imag} */,
  {32'h3e83636a, 32'hc090ec44} /* (26, 7, 6) {real, imag} */,
  {32'hbf59e2fe, 32'hbffae81a} /* (26, 7, 5) {real, imag} */,
  {32'hbf56d9cc, 32'h3f6db777} /* (26, 7, 4) {real, imag} */,
  {32'h3f1fbc23, 32'hbf0e6f58} /* (26, 7, 3) {real, imag} */,
  {32'hbf96143a, 32'hbfad052b} /* (26, 7, 2) {real, imag} */,
  {32'hbe6d926c, 32'hbfc3a9df} /* (26, 7, 1) {real, imag} */,
  {32'h3f8039e4, 32'hbf8bd933} /* (26, 7, 0) {real, imag} */,
  {32'h3e756870, 32'hbed0aa88} /* (26, 6, 31) {real, imag} */,
  {32'h3ebda694, 32'h3d8e9f38} /* (26, 6, 30) {real, imag} */,
  {32'hbf27065e, 32'h3ee55db4} /* (26, 6, 29) {real, imag} */,
  {32'hbf537536, 32'h3ed077c6} /* (26, 6, 28) {real, imag} */,
  {32'h3f43e10c, 32'h3fcd576e} /* (26, 6, 27) {real, imag} */,
  {32'h3fe0cc50, 32'hbeb53034} /* (26, 6, 26) {real, imag} */,
  {32'h3f99a10d, 32'hbf660d92} /* (26, 6, 25) {real, imag} */,
  {32'h3f89204c, 32'hbfcea037} /* (26, 6, 24) {real, imag} */,
  {32'h3f438c03, 32'hc070bc50} /* (26, 6, 23) {real, imag} */,
  {32'hbdd0ad18, 32'hc020309c} /* (26, 6, 22) {real, imag} */,
  {32'h3f959ed5, 32'hbfaaf5f8} /* (26, 6, 21) {real, imag} */,
  {32'h3ff3ca49, 32'h3f2c3120} /* (26, 6, 20) {real, imag} */,
  {32'h400c91ca, 32'hbfc54760} /* (26, 6, 19) {real, imag} */,
  {32'h3e4e5ec8, 32'hbfa4f2d0} /* (26, 6, 18) {real, imag} */,
  {32'hbedadf10, 32'h3f77d0cb} /* (26, 6, 17) {real, imag} */,
  {32'h3f7fb6d2, 32'hbf4e96e2} /* (26, 6, 16) {real, imag} */,
  {32'h40033092, 32'hbf3358c8} /* (26, 6, 15) {real, imag} */,
  {32'h3f7da980, 32'hbfbbe416} /* (26, 6, 14) {real, imag} */,
  {32'h3f781329, 32'hbf34910b} /* (26, 6, 13) {real, imag} */,
  {32'hbf2635cd, 32'h3d4f19d0} /* (26, 6, 12) {real, imag} */,
  {32'h3fb4df81, 32'h3f349ebd} /* (26, 6, 11) {real, imag} */,
  {32'h3fffbf39, 32'hbf877a67} /* (26, 6, 10) {real, imag} */,
  {32'hbedf9db4, 32'hc04ea182} /* (26, 6, 9) {real, imag} */,
  {32'h3fd4215e, 32'hbee3e7a6} /* (26, 6, 8) {real, imag} */,
  {32'h403c46e2, 32'hc00e8fc0} /* (26, 6, 7) {real, imag} */,
  {32'h3f63a0ce, 32'hbfe7f4bc} /* (26, 6, 6) {real, imag} */,
  {32'h3f8ad952, 32'h3d4c4db0} /* (26, 6, 5) {real, imag} */,
  {32'h3ec6aab4, 32'h3fcc8c78} /* (26, 6, 4) {real, imag} */,
  {32'h3ec1d5e6, 32'hbe0e85c4} /* (26, 6, 3) {real, imag} */,
  {32'h3f25b8b2, 32'h3e189ff8} /* (26, 6, 2) {real, imag} */,
  {32'h3fcc1236, 32'hbd518700} /* (26, 6, 1) {real, imag} */,
  {32'h3f86c974, 32'hbf9f6fb9} /* (26, 6, 0) {real, imag} */,
  {32'h3e9c441c, 32'hbef58270} /* (26, 5, 31) {real, imag} */,
  {32'hbe7ea4fc, 32'hbee38b92} /* (26, 5, 30) {real, imag} */,
  {32'hbf5cf1c2, 32'h3e8d9da0} /* (26, 5, 29) {real, imag} */,
  {32'hbff14e4e, 32'hbf6d9aa6} /* (26, 5, 28) {real, imag} */,
  {32'hbefb5bac, 32'h40010788} /* (26, 5, 27) {real, imag} */,
  {32'hbd086cc0, 32'h3eb63172} /* (26, 5, 26) {real, imag} */,
  {32'h3f8e64ec, 32'h3fb46f7d} /* (26, 5, 25) {real, imag} */,
  {32'h3f95ecd4, 32'h3f286a42} /* (26, 5, 24) {real, imag} */,
  {32'h3f5fe954, 32'hbf3d99cc} /* (26, 5, 23) {real, imag} */,
  {32'hbfd53a05, 32'hc02b8a5e} /* (26, 5, 22) {real, imag} */,
  {32'hc06d6ddc, 32'hbfa778a0} /* (26, 5, 21) {real, imag} */,
  {32'hc01bd3b8, 32'hbf2eff9e} /* (26, 5, 20) {real, imag} */,
  {32'h3e5aac04, 32'hbebb2a7e} /* (26, 5, 19) {real, imag} */,
  {32'h3fb570a9, 32'h3f9e491e} /* (26, 5, 18) {real, imag} */,
  {32'hbfc3daae, 32'h3fe84e5e} /* (26, 5, 17) {real, imag} */,
  {32'hbfbebf69, 32'hbffc5285} /* (26, 5, 16) {real, imag} */,
  {32'h3f3241c2, 32'hbfefe0c9} /* (26, 5, 15) {real, imag} */,
  {32'h400c4ca2, 32'hc01cf5e0} /* (26, 5, 14) {real, imag} */,
  {32'h3f453aef, 32'hbf503bf2} /* (26, 5, 13) {real, imag} */,
  {32'hbf9983c2, 32'hbe842848} /* (26, 5, 12) {real, imag} */,
  {32'hbf8bd8a4, 32'h3f8252b6} /* (26, 5, 11) {real, imag} */,
  {32'h3f989bbe, 32'h3f897732} /* (26, 5, 10) {real, imag} */,
  {32'h40290a04, 32'hbd205b18} /* (26, 5, 9) {real, imag} */,
  {32'h4037c756, 32'hbf8a5578} /* (26, 5, 8) {real, imag} */,
  {32'h402195e4, 32'hc05cbeeb} /* (26, 5, 7) {real, imag} */,
  {32'h3b711c00, 32'hc01c7e30} /* (26, 5, 6) {real, imag} */,
  {32'hbf39cd18, 32'hbd2a8440} /* (26, 5, 5) {real, imag} */,
  {32'hbf339d51, 32'h3dfb8430} /* (26, 5, 4) {real, imag} */,
  {32'hbf6facbf, 32'h3f08a71c} /* (26, 5, 3) {real, imag} */,
  {32'hbfc476ad, 32'h3eed3ff4} /* (26, 5, 2) {real, imag} */,
  {32'hbe7e6e88, 32'h3f90109a} /* (26, 5, 1) {real, imag} */,
  {32'hbf613a34, 32'hbf346ea6} /* (26, 5, 0) {real, imag} */,
  {32'h3f81cff4, 32'hbf55485f} /* (26, 4, 31) {real, imag} */,
  {32'h40016dfc, 32'hbfc1fde4} /* (26, 4, 30) {real, imag} */,
  {32'h3f3e57a3, 32'hbeb860c0} /* (26, 4, 29) {real, imag} */,
  {32'hbfa2dfbb, 32'hbe03f660} /* (26, 4, 28) {real, imag} */,
  {32'hc004f95c, 32'hbfa3c21d} /* (26, 4, 27) {real, imag} */,
  {32'hbf411f53, 32'hc0785c09} /* (26, 4, 26) {real, imag} */,
  {32'hbd966314, 32'hc00b54d6} /* (26, 4, 25) {real, imag} */,
  {32'hbf1bba5f, 32'h3f688270} /* (26, 4, 24) {real, imag} */,
  {32'h3f83063e, 32'h3fd8e372} /* (26, 4, 23) {real, imag} */,
  {32'h3f8f1904, 32'hbfd55830} /* (26, 4, 22) {real, imag} */,
  {32'hbfb5348c, 32'hbf1818c4} /* (26, 4, 21) {real, imag} */,
  {32'hc016539c, 32'hbf82dc7c} /* (26, 4, 20) {real, imag} */,
  {32'hbf6201e6, 32'h3fa9543b} /* (26, 4, 19) {real, imag} */,
  {32'h3f0371b9, 32'h409b09bc} /* (26, 4, 18) {real, imag} */,
  {32'h3f1e8c2a, 32'h401c1732} /* (26, 4, 17) {real, imag} */,
  {32'hbf8b30cd, 32'h3de7c220} /* (26, 4, 16) {real, imag} */,
  {32'hc0036b89, 32'hbfcfc9bc} /* (26, 4, 15) {real, imag} */,
  {32'h3fb115d2, 32'hc05589e6} /* (26, 4, 14) {real, imag} */,
  {32'hbd0d0d70, 32'hc0029086} /* (26, 4, 13) {real, imag} */,
  {32'hbf38639e, 32'hbe94bc0c} /* (26, 4, 12) {real, imag} */,
  {32'hbe8de412, 32'h3f9b86ce} /* (26, 4, 11) {real, imag} */,
  {32'h3f0b8d0a, 32'h3f8da1b1} /* (26, 4, 10) {real, imag} */,
  {32'h3fdb79e2, 32'h3fdf2635} /* (26, 4, 9) {real, imag} */,
  {32'hbf4b6cbe, 32'hbfada844} /* (26, 4, 8) {real, imag} */,
  {32'hbe8c35a8, 32'hbfedb118} /* (26, 4, 7) {real, imag} */,
  {32'hbe9eeb7a, 32'hc01768e7} /* (26, 4, 6) {real, imag} */,
  {32'h3f4f66d0, 32'hc0024ba0} /* (26, 4, 5) {real, imag} */,
  {32'h3e7ee268, 32'hbfb0b6f9} /* (26, 4, 4) {real, imag} */,
  {32'hc00ab8fa, 32'hbda90ee0} /* (26, 4, 3) {real, imag} */,
  {32'hc02556a2, 32'h3f0abfa0} /* (26, 4, 2) {real, imag} */,
  {32'h3ee48794, 32'h3d9d2800} /* (26, 4, 1) {real, imag} */,
  {32'hbf0a84d3, 32'hbf751d13} /* (26, 4, 0) {real, imag} */,
  {32'hbe9c5ab0, 32'hbf947c88} /* (26, 3, 31) {real, imag} */,
  {32'h3fa679a2, 32'hc010b770} /* (26, 3, 30) {real, imag} */,
  {32'h3fabb16f, 32'h3f67c4e2} /* (26, 3, 29) {real, imag} */,
  {32'h3fa66b21, 32'h3ff21b34} /* (26, 3, 28) {real, imag} */,
  {32'hbfc50bda, 32'hbf7ae8f0} /* (26, 3, 27) {real, imag} */,
  {32'hc0072554, 32'hc05a4ca2} /* (26, 3, 26) {real, imag} */,
  {32'hbf9a1c68, 32'hc02073a5} /* (26, 3, 25) {real, imag} */,
  {32'hc003588d, 32'h3ec5bfa6} /* (26, 3, 24) {real, imag} */,
  {32'hbe74ca08, 32'h3edfc52e} /* (26, 3, 23) {real, imag} */,
  {32'h3fc4e584, 32'hbf6d5018} /* (26, 3, 22) {real, imag} */,
  {32'hbe9f117e, 32'hbe97b70c} /* (26, 3, 21) {real, imag} */,
  {32'h3fae32ef, 32'h3f3eda2a} /* (26, 3, 20) {real, imag} */,
  {32'h40143319, 32'h3e99462c} /* (26, 3, 19) {real, imag} */,
  {32'hbfe33621, 32'hbe8a88ac} /* (26, 3, 18) {real, imag} */,
  {32'hbf13ca1e, 32'h3fb4efb4} /* (26, 3, 17) {real, imag} */,
  {32'h3f87f8c2, 32'h400c5539} /* (26, 3, 16) {real, imag} */,
  {32'hbebe78f1, 32'h3fff26a2} /* (26, 3, 15) {real, imag} */,
  {32'h3ec280f6, 32'h3f244460} /* (26, 3, 14) {real, imag} */,
  {32'hc000af84, 32'hbd5537a0} /* (26, 3, 13) {real, imag} */,
  {32'hbef812c0, 32'h3fbbd5cb} /* (26, 3, 12) {real, imag} */,
  {32'h3fb02355, 32'h405620ae} /* (26, 3, 11) {real, imag} */,
  {32'hbf2cd5a6, 32'h40080708} /* (26, 3, 10) {real, imag} */,
  {32'hbf27f3d0, 32'h3d97d198} /* (26, 3, 9) {real, imag} */,
  {32'hbfe38bf1, 32'hbf6eefc2} /* (26, 3, 8) {real, imag} */,
  {32'h3e1a4ba0, 32'hc0248e4b} /* (26, 3, 7) {real, imag} */,
  {32'hbf2f19bd, 32'hc078063e} /* (26, 3, 6) {real, imag} */,
  {32'hbdd56e14, 32'hc07da054} /* (26, 3, 5) {real, imag} */,
  {32'h3f29a2f2, 32'hc01d8390} /* (26, 3, 4) {real, imag} */,
  {32'hbf76e542, 32'hbf81669c} /* (26, 3, 3) {real, imag} */,
  {32'h3de505dc, 32'hbe8039c4} /* (26, 3, 2) {real, imag} */,
  {32'h4007806b, 32'h3e360d80} /* (26, 3, 1) {real, imag} */,
  {32'h3f41b860, 32'hbf8bce09} /* (26, 3, 0) {real, imag} */,
  {32'hbf1edfea, 32'hbf1c2741} /* (26, 2, 31) {real, imag} */,
  {32'h3f5f4a93, 32'hbf8fee7e} /* (26, 2, 30) {real, imag} */,
  {32'hbf59e182, 32'h3df48630} /* (26, 2, 29) {real, imag} */,
  {32'hbea75850, 32'h3ffc28c3} /* (26, 2, 28) {real, imag} */,
  {32'h3f0b298c, 32'h3faaf4b5} /* (26, 2, 27) {real, imag} */,
  {32'hc0397f8c, 32'hbfa34728} /* (26, 2, 26) {real, imag} */,
  {32'hc00a91ad, 32'hbf2b82c8} /* (26, 2, 25) {real, imag} */,
  {32'hbfe12932, 32'h3f6f69db} /* (26, 2, 24) {real, imag} */,
  {32'h3c86dc40, 32'h402bff32} /* (26, 2, 23) {real, imag} */,
  {32'h3f9238c8, 32'h3fbbf398} /* (26, 2, 22) {real, imag} */,
  {32'h3fa535a2, 32'h4009520b} /* (26, 2, 21) {real, imag} */,
  {32'h4085f3a6, 32'h407300c0} /* (26, 2, 20) {real, imag} */,
  {32'h409a547c, 32'hbec688d0} /* (26, 2, 19) {real, imag} */,
  {32'h3f9b80da, 32'hc01e139d} /* (26, 2, 18) {real, imag} */,
  {32'h3f10778a, 32'hc041ed86} /* (26, 2, 17) {real, imag} */,
  {32'h3faa767a, 32'hbf56fc64} /* (26, 2, 16) {real, imag} */,
  {32'hbf1855bc, 32'h3f2a25ee} /* (26, 2, 15) {real, imag} */,
  {32'hbd78c3c0, 32'h3fbc94da} /* (26, 2, 14) {real, imag} */,
  {32'hbe9619e0, 32'h4019f3bf} /* (26, 2, 13) {real, imag} */,
  {32'hbf56adef, 32'h3f5fe2a2} /* (26, 2, 12) {real, imag} */,
  {32'hbec819dc, 32'h40698906} /* (26, 2, 11) {real, imag} */,
  {32'hbf5fb3f4, 32'h3eed2824} /* (26, 2, 10) {real, imag} */,
  {32'h3f188d26, 32'hbf599c68} /* (26, 2, 9) {real, imag} */,
  {32'hbe00b360, 32'hbe9086a4} /* (26, 2, 8) {real, imag} */,
  {32'hbd375030, 32'hbfbc7c1a} /* (26, 2, 7) {real, imag} */,
  {32'hbf84d459, 32'hbfa8aae3} /* (26, 2, 6) {real, imag} */,
  {32'hc0109e0a, 32'hc032f131} /* (26, 2, 5) {real, imag} */,
  {32'hbfb47204, 32'hbf0447d0} /* (26, 2, 4) {real, imag} */,
  {32'h3f7cfc2b, 32'hbf099087} /* (26, 2, 3) {real, imag} */,
  {32'h3f8acfda, 32'hbf5ac0b0} /* (26, 2, 2) {real, imag} */,
  {32'h3f46ba52, 32'h3f0260a6} /* (26, 2, 1) {real, imag} */,
  {32'hbea6b6e4, 32'h3ed0d324} /* (26, 2, 0) {real, imag} */,
  {32'h3f8b66c6, 32'hbca28600} /* (26, 1, 31) {real, imag} */,
  {32'h40030aca, 32'hbe764c08} /* (26, 1, 30) {real, imag} */,
  {32'h3f66a61b, 32'h3ec4a988} /* (26, 1, 29) {real, imag} */,
  {32'h3e62ce40, 32'h3fd89acf} /* (26, 1, 28) {real, imag} */,
  {32'h3fc0973a, 32'h3f7e988e} /* (26, 1, 27) {real, imag} */,
  {32'hbfdb18bc, 32'hbfaa59bd} /* (26, 1, 26) {real, imag} */,
  {32'hc00aed21, 32'hbfe7db67} /* (26, 1, 25) {real, imag} */,
  {32'hbfa788e4, 32'hbe0ca958} /* (26, 1, 24) {real, imag} */,
  {32'hbe65ae48, 32'h405ba102} /* (26, 1, 23) {real, imag} */,
  {32'hbf67ac4f, 32'h3f9836a6} /* (26, 1, 22) {real, imag} */,
  {32'hba2a4400, 32'h4099634d} /* (26, 1, 21) {real, imag} */,
  {32'h3eabce68, 32'h402b739a} /* (26, 1, 20) {real, imag} */,
  {32'h3ffe7c8c, 32'hbf5df26c} /* (26, 1, 19) {real, imag} */,
  {32'h3f651da8, 32'hbd87d760} /* (26, 1, 18) {real, imag} */,
  {32'hbf0d38ae, 32'hbfb7a6ce} /* (26, 1, 17) {real, imag} */,
  {32'hbf53db6a, 32'h3d877c68} /* (26, 1, 16) {real, imag} */,
  {32'hbfc8480c, 32'h3f1b8473} /* (26, 1, 15) {real, imag} */,
  {32'h3fa2af52, 32'h4029cde9} /* (26, 1, 14) {real, imag} */,
  {32'h3f9174c0, 32'h40644110} /* (26, 1, 13) {real, imag} */,
  {32'h3f5342d0, 32'h3f8d1db8} /* (26, 1, 12) {real, imag} */,
  {32'h3e005e50, 32'h3fdd6fc0} /* (26, 1, 11) {real, imag} */,
  {32'hbefafa6e, 32'hbece91cc} /* (26, 1, 10) {real, imag} */,
  {32'h3f57b870, 32'hbf7463a0} /* (26, 1, 9) {real, imag} */,
  {32'h3f3bdfa8, 32'h3f5e98ba} /* (26, 1, 8) {real, imag} */,
  {32'hbf71c51e, 32'hbe145b68} /* (26, 1, 7) {real, imag} */,
  {32'hbfb223ca, 32'h3f305602} /* (26, 1, 6) {real, imag} */,
  {32'hc023b622, 32'hbf2d58bc} /* (26, 1, 5) {real, imag} */,
  {32'hbfcd5595, 32'hbe637068} /* (26, 1, 4) {real, imag} */,
  {32'hbf24ac61, 32'h3f4222aa} /* (26, 1, 3) {real, imag} */,
  {32'hbef80bf7, 32'hbf967d27} /* (26, 1, 2) {real, imag} */,
  {32'h3fefa6fa, 32'h3f8ce932} /* (26, 1, 1) {real, imag} */,
  {32'h3f0936d1, 32'h3fe27d22} /* (26, 1, 0) {real, imag} */,
  {32'h3fab7342, 32'hbf12af5f} /* (26, 0, 31) {real, imag} */,
  {32'h3fd0d210, 32'hbede6772} /* (26, 0, 30) {real, imag} */,
  {32'h3fb08fcb, 32'h3ed05c10} /* (26, 0, 29) {real, imag} */,
  {32'h3fe72478, 32'h3f3d70e8} /* (26, 0, 28) {real, imag} */,
  {32'h3f60b7fb, 32'h3e906b6a} /* (26, 0, 27) {real, imag} */,
  {32'hbfe268dc, 32'hbf23faeb} /* (26, 0, 26) {real, imag} */,
  {32'hbf37043c, 32'hbe6973ba} /* (26, 0, 25) {real, imag} */,
  {32'hbe44f1a0, 32'hbe4b97b4} /* (26, 0, 24) {real, imag} */,
  {32'h3cf343c0, 32'h3d7e8fa0} /* (26, 0, 23) {real, imag} */,
  {32'hbf8ac449, 32'hbf18bbd2} /* (26, 0, 22) {real, imag} */,
  {32'hbf2a2be6, 32'h3fe584a3} /* (26, 0, 21) {real, imag} */,
  {32'hbfdd4f1e, 32'h3f567398} /* (26, 0, 20) {real, imag} */,
  {32'hbe4815e0, 32'h3e8b972e} /* (26, 0, 19) {real, imag} */,
  {32'hbf2349be, 32'h3d1db850} /* (26, 0, 18) {real, imag} */,
  {32'hbfcf0b44, 32'h3f1e355b} /* (26, 0, 17) {real, imag} */,
  {32'hbfc9ab66, 32'h3ebe88c2} /* (26, 0, 16) {real, imag} */,
  {32'hbf4b9ace, 32'h3e797ec8} /* (26, 0, 15) {real, imag} */,
  {32'h400413e3, 32'h3ff0236e} /* (26, 0, 14) {real, imag} */,
  {32'h3fba0535, 32'h3fb8d942} /* (26, 0, 13) {real, imag} */,
  {32'h3ff7b938, 32'hbf84bb18} /* (26, 0, 12) {real, imag} */,
  {32'h400ed162, 32'h3e201a20} /* (26, 0, 11) {real, imag} */,
  {32'h3fc9e64f, 32'h3fbffd6e} /* (26, 0, 10) {real, imag} */,
  {32'h3edca77e, 32'h3e6c1190} /* (26, 0, 9) {real, imag} */,
  {32'hbf1c15dc, 32'h3fa7a0be} /* (26, 0, 8) {real, imag} */,
  {32'hbfff8945, 32'h3f8347b4} /* (26, 0, 7) {real, imag} */,
  {32'hc01f47ef, 32'h3f25f69e} /* (26, 0, 6) {real, imag} */,
  {32'hbf6f4e72, 32'h3f7e00a5} /* (26, 0, 5) {real, imag} */,
  {32'hbe79acf0, 32'h3f532ece} /* (26, 0, 4) {real, imag} */,
  {32'h3eb4b83a, 32'h3f903a80} /* (26, 0, 3) {real, imag} */,
  {32'h3f7e7832, 32'hbf307c09} /* (26, 0, 2) {real, imag} */,
  {32'h3ffcf58c, 32'h3edd6140} /* (26, 0, 1) {real, imag} */,
  {32'h3f44131e, 32'h3f8be2da} /* (26, 0, 0) {real, imag} */,
  {32'hbf8f6ba8, 32'hbe8e2108} /* (25, 31, 31) {real, imag} */,
  {32'hbf839c43, 32'hbf5197d2} /* (25, 31, 30) {real, imag} */,
  {32'hbfe2b12b, 32'hbd1e6080} /* (25, 31, 29) {real, imag} */,
  {32'hbf029e6e, 32'hbe7fa802} /* (25, 31, 28) {real, imag} */,
  {32'hbd206838, 32'hbf886002} /* (25, 31, 27) {real, imag} */,
  {32'hbfa4d401, 32'hbf5885d8} /* (25, 31, 26) {real, imag} */,
  {32'h3a179c00, 32'h3f0e26d0} /* (25, 31, 25) {real, imag} */,
  {32'h3f7b91f8, 32'h3fe109c0} /* (25, 31, 24) {real, imag} */,
  {32'h3fb5811e, 32'h3f8b1ce0} /* (25, 31, 23) {real, imag} */,
  {32'h3f991b21, 32'h3ea66a03} /* (25, 31, 22) {real, imag} */,
  {32'h3f96b794, 32'h3f153dea} /* (25, 31, 21) {real, imag} */,
  {32'h3fa30cc1, 32'h3fae2479} /* (25, 31, 20) {real, imag} */,
  {32'hbd8be810, 32'h3f760419} /* (25, 31, 19) {real, imag} */,
  {32'h3dbb40a4, 32'h3f3e043e} /* (25, 31, 18) {real, imag} */,
  {32'h3ef74bc8, 32'hbf3fe5fa} /* (25, 31, 17) {real, imag} */,
  {32'h3f40902e, 32'hbe13c1be} /* (25, 31, 16) {real, imag} */,
  {32'h3e2f5f03, 32'hbf45cf06} /* (25, 31, 15) {real, imag} */,
  {32'hbfc07db2, 32'hbe32990f} /* (25, 31, 14) {real, imag} */,
  {32'hbfff7603, 32'hbfafb13a} /* (25, 31, 13) {real, imag} */,
  {32'h3ed0239c, 32'hc0147afe} /* (25, 31, 12) {real, imag} */,
  {32'h3fefa61a, 32'hbfd65368} /* (25, 31, 11) {real, imag} */,
  {32'hbe0d0bc7, 32'hc001268e} /* (25, 31, 10) {real, imag} */,
  {32'h3e1d0d3c, 32'h3ce0da90} /* (25, 31, 9) {real, imag} */,
  {32'h3f6398a5, 32'h3f62cd50} /* (25, 31, 8) {real, imag} */,
  {32'h400f4538, 32'h3e95e618} /* (25, 31, 7) {real, imag} */,
  {32'h3d897a70, 32'hbf00549a} /* (25, 31, 6) {real, imag} */,
  {32'hbe54c9c8, 32'hc03022d1} /* (25, 31, 5) {real, imag} */,
  {32'hbecd2d9f, 32'hbfd424ee} /* (25, 31, 4) {real, imag} */,
  {32'hbfade374, 32'h3f0d0bd7} /* (25, 31, 3) {real, imag} */,
  {32'hbe79bc77, 32'h3eafa922} /* (25, 31, 2) {real, imag} */,
  {32'h3f464511, 32'h3f9a84c6} /* (25, 31, 1) {real, imag} */,
  {32'hbf84740a, 32'h3f32b4c0} /* (25, 31, 0) {real, imag} */,
  {32'hbfc86320, 32'h3f8914d7} /* (25, 30, 31) {real, imag} */,
  {32'hbfd0da86, 32'h3f9b3c08} /* (25, 30, 30) {real, imag} */,
  {32'hbfac0794, 32'h3f934f94} /* (25, 30, 29) {real, imag} */,
  {32'h3f81ff44, 32'h3eefa6ed} /* (25, 30, 28) {real, imag} */,
  {32'h3face322, 32'hbf9fc338} /* (25, 30, 27) {real, imag} */,
  {32'hbf3d221e, 32'h3e9ded64} /* (25, 30, 26) {real, imag} */,
  {32'h3eb89214, 32'h3f42b2e0} /* (25, 30, 25) {real, imag} */,
  {32'h3e748ed8, 32'h4029f24e} /* (25, 30, 24) {real, imag} */,
  {32'hbce451d0, 32'h3f4587d4} /* (25, 30, 23) {real, imag} */,
  {32'h3d8ebe02, 32'hbfba42cc} /* (25, 30, 22) {real, imag} */,
  {32'hbf0caa55, 32'hbd18d308} /* (25, 30, 21) {real, imag} */,
  {32'hbd295f30, 32'h3f421f60} /* (25, 30, 20) {real, imag} */,
  {32'hc018912a, 32'h3e7f5d94} /* (25, 30, 19) {real, imag} */,
  {32'hc0097128, 32'h3f32e9d9} /* (25, 30, 18) {real, imag} */,
  {32'h3fb186bd, 32'hbdd6dd32} /* (25, 30, 17) {real, imag} */,
  {32'h3f6349ba, 32'h3f9a5b7d} /* (25, 30, 16) {real, imag} */,
  {32'hbfd2080b, 32'h3e9a8c0c} /* (25, 30, 15) {real, imag} */,
  {32'hbff03075, 32'hbf6315c4} /* (25, 30, 14) {real, imag} */,
  {32'hbfcd0672, 32'hc01d3506} /* (25, 30, 13) {real, imag} */,
  {32'hbe5606ac, 32'hc0771ee5} /* (25, 30, 12) {real, imag} */,
  {32'h3facd87e, 32'hbf4a06fc} /* (25, 30, 11) {real, imag} */,
  {32'h3f14cf43, 32'hbe2a4b58} /* (25, 30, 10) {real, imag} */,
  {32'h3ef7e768, 32'h3fac9967} /* (25, 30, 9) {real, imag} */,
  {32'h3eda22ca, 32'h3fec78ea} /* (25, 30, 8) {real, imag} */,
  {32'h402a4eea, 32'h3e4acfc0} /* (25, 30, 7) {real, imag} */,
  {32'hbf90025d, 32'hbfb1f7d0} /* (25, 30, 6) {real, imag} */,
  {32'hc03cffe2, 32'hc02e11b7} /* (25, 30, 5) {real, imag} */,
  {32'hbffa6b44, 32'hc0122946} /* (25, 30, 4) {real, imag} */,
  {32'hbfa8c09c, 32'hbf274deb} /* (25, 30, 3) {real, imag} */,
  {32'h3d80ba10, 32'h3f393a7a} /* (25, 30, 2) {real, imag} */,
  {32'h3e03663c, 32'h405c00c2} /* (25, 30, 1) {real, imag} */,
  {32'hbf86022d, 32'h400a5e52} /* (25, 30, 0) {real, imag} */,
  {32'hbf3d74ad, 32'h3f66aaac} /* (25, 29, 31) {real, imag} */,
  {32'hbf38b68a, 32'h3f495aa8} /* (25, 29, 30) {real, imag} */,
  {32'hbf9282d3, 32'h3e5a53a8} /* (25, 29, 29) {real, imag} */,
  {32'h3fe03a80, 32'h400cf7fe} /* (25, 29, 28) {real, imag} */,
  {32'h406c079e, 32'h3fbb034f} /* (25, 29, 27) {real, imag} */,
  {32'h3fa5bee0, 32'hbd9552a8} /* (25, 29, 26) {real, imag} */,
  {32'h3f22aec6, 32'h3e650fc8} /* (25, 29, 25) {real, imag} */,
  {32'h3b86d500, 32'h3feb9a32} /* (25, 29, 24) {real, imag} */,
  {32'hbfb53e62, 32'h3ee230b7} /* (25, 29, 23) {real, imag} */,
  {32'hbe288ea8, 32'hbf54355c} /* (25, 29, 22) {real, imag} */,
  {32'hbf8c519f, 32'h3fe5e506} /* (25, 29, 21) {real, imag} */,
  {32'hbff4fe24, 32'h3f8fe0ae} /* (25, 29, 20) {real, imag} */,
  {32'hc078936d, 32'hbfcba601} /* (25, 29, 19) {real, imag} */,
  {32'hc0550d76, 32'hbd3153d0} /* (25, 29, 18) {real, imag} */,
  {32'h3f0ff873, 32'hbf2853a7} /* (25, 29, 17) {real, imag} */,
  {32'h3f3de902, 32'hbdca16c0} /* (25, 29, 16) {real, imag} */,
  {32'hbfbe4430, 32'hbd717d10} /* (25, 29, 15) {real, imag} */,
  {32'hbd974360, 32'hbe00b920} /* (25, 29, 14) {real, imag} */,
  {32'h3f9f1336, 32'hbe28dd58} /* (25, 29, 13) {real, imag} */,
  {32'hbf1375ae, 32'hbffe276e} /* (25, 29, 12) {real, imag} */,
  {32'hbf41c8ca, 32'h3efc2a7a} /* (25, 29, 11) {real, imag} */,
  {32'hbc40b880, 32'h40033830} /* (25, 29, 10) {real, imag} */,
  {32'hbecdd678, 32'h3fa05eba} /* (25, 29, 9) {real, imag} */,
  {32'hbf4bff80, 32'h3ffda430} /* (25, 29, 8) {real, imag} */,
  {32'hbeafd484, 32'h3f6ff917} /* (25, 29, 7) {real, imag} */,
  {32'hc032de7c, 32'hbf1addbc} /* (25, 29, 6) {real, imag} */,
  {32'hc0821e54, 32'hbf598410} /* (25, 29, 5) {real, imag} */,
  {32'hbf83e00c, 32'hbede1872} /* (25, 29, 4) {real, imag} */,
  {32'h3f1f618c, 32'hc01048ac} /* (25, 29, 3) {real, imag} */,
  {32'h3fa45796, 32'hc0407793} /* (25, 29, 2) {real, imag} */,
  {32'h3ed8e06e, 32'h3f1a445d} /* (25, 29, 1) {real, imag} */,
  {32'hbfde07a0, 32'h3fde0056} /* (25, 29, 0) {real, imag} */,
  {32'h3e5a24e6, 32'hbf7c42f0} /* (25, 28, 31) {real, imag} */,
  {32'hbf9551e3, 32'hc0069222} /* (25, 28, 30) {real, imag} */,
  {32'hc0629421, 32'hbf4ea468} /* (25, 28, 29) {real, imag} */,
  {32'h3ef0c24b, 32'h3fadb1b1} /* (25, 28, 28) {real, imag} */,
  {32'h4065801f, 32'h3fdf23e4} /* (25, 28, 27) {real, imag} */,
  {32'h3d945982, 32'hbfc45960} /* (25, 28, 26) {real, imag} */,
  {32'hbf2ae3da, 32'h3df81130} /* (25, 28, 25) {real, imag} */,
  {32'h3f71bbb0, 32'h3f1712d5} /* (25, 28, 24) {real, imag} */,
  {32'h3f82d485, 32'h3f135252} /* (25, 28, 23) {real, imag} */,
  {32'h400b0378, 32'h40482ab5} /* (25, 28, 22) {real, imag} */,
  {32'h3ff201d8, 32'h4006fd4a} /* (25, 28, 21) {real, imag} */,
  {32'h3f819a94, 32'h3fbefd65} /* (25, 28, 20) {real, imag} */,
  {32'hbfbbcf98, 32'hbec17c40} /* (25, 28, 19) {real, imag} */,
  {32'hc0047c7e, 32'hbe359c28} /* (25, 28, 18) {real, imag} */,
  {32'hbf6cce08, 32'hbf931f60} /* (25, 28, 17) {real, imag} */,
  {32'hbf9003a9, 32'h3f7ae97c} /* (25, 28, 16) {real, imag} */,
  {32'hbf7135a0, 32'h3f719681} /* (25, 28, 15) {real, imag} */,
  {32'hbf0b083c, 32'h3d950da0} /* (25, 28, 14) {real, imag} */,
  {32'h3f9eb4fe, 32'h3f9020b9} /* (25, 28, 13) {real, imag} */,
  {32'hbf6d2f02, 32'hbdf066e8} /* (25, 28, 12) {real, imag} */,
  {32'hbf779898, 32'h3f51b8c3} /* (25, 28, 11) {real, imag} */,
  {32'h4005f14a, 32'h403df1eb} /* (25, 28, 10) {real, imag} */,
  {32'h40532fd2, 32'h402a5d27} /* (25, 28, 9) {real, imag} */,
  {32'h3e850d13, 32'h3fab7aac} /* (25, 28, 8) {real, imag} */,
  {32'hbf777b89, 32'h3f97a525} /* (25, 28, 7) {real, imag} */,
  {32'hc0012220, 32'h3f3faf16} /* (25, 28, 6) {real, imag} */,
  {32'h3e975f24, 32'h3f53cfa6} /* (25, 28, 5) {real, imag} */,
  {32'h3fac2dd3, 32'h3fdf7c02} /* (25, 28, 4) {real, imag} */,
  {32'h3f605b49, 32'h3fcaa59b} /* (25, 28, 3) {real, imag} */,
  {32'h3f134f17, 32'hbf88d41e} /* (25, 28, 2) {real, imag} */,
  {32'h3f5aa6cc, 32'hbf9bb667} /* (25, 28, 1) {real, imag} */,
  {32'hbe977dc4, 32'hbf63fd4e} /* (25, 28, 0) {real, imag} */,
  {32'hbfeb98bc, 32'hbef5f246} /* (25, 27, 31) {real, imag} */,
  {32'hbfdb3f62, 32'hbf8f481b} /* (25, 27, 30) {real, imag} */,
  {32'hbde312b8, 32'hbe98bc14} /* (25, 27, 29) {real, imag} */,
  {32'h3f9086b8, 32'hbfbb3382} /* (25, 27, 28) {real, imag} */,
  {32'h3fb0428b, 32'h3d463ea0} /* (25, 27, 27) {real, imag} */,
  {32'hbfa814a6, 32'hbe38c514} /* (25, 27, 26) {real, imag} */,
  {32'hbf8cebf0, 32'h3bfa33c0} /* (25, 27, 25) {real, imag} */,
  {32'h3f0d8315, 32'h3fa22daf} /* (25, 27, 24) {real, imag} */,
  {32'h3f149380, 32'h3f27e572} /* (25, 27, 23) {real, imag} */,
  {32'h4007fe44, 32'h408876a9} /* (25, 27, 22) {real, imag} */,
  {32'h3ff7925b, 32'h3fe4385b} /* (25, 27, 21) {real, imag} */,
  {32'h3f42475a, 32'hbfb4e3b2} /* (25, 27, 20) {real, imag} */,
  {32'h3ebf1698, 32'hbfba7a60} /* (25, 27, 19) {real, imag} */,
  {32'h3f1652e0, 32'hbde47da8} /* (25, 27, 18) {real, imag} */,
  {32'h3e644b38, 32'h3de233d0} /* (25, 27, 17) {real, imag} */,
  {32'hbf453acc, 32'h3e851210} /* (25, 27, 16) {real, imag} */,
  {32'h3f2d5300, 32'h40017102} /* (25, 27, 15) {real, imag} */,
  {32'h400a425a, 32'hbe0a6e70} /* (25, 27, 14) {real, imag} */,
  {32'h3fa55b4f, 32'hbfb8e2a6} /* (25, 27, 13) {real, imag} */,
  {32'hbf5c92ca, 32'h3c8fede0} /* (25, 27, 12) {real, imag} */,
  {32'hbfd939b2, 32'hbdf808b0} /* (25, 27, 11) {real, imag} */,
  {32'h3ee5eed0, 32'h4000ffeb} /* (25, 27, 10) {real, imag} */,
  {32'h40225cb4, 32'h401b1a3a} /* (25, 27, 9) {real, imag} */,
  {32'h3f55b975, 32'h3fe01d07} /* (25, 27, 8) {real, imag} */,
  {32'h3fa60c43, 32'h40230300} /* (25, 27, 7) {real, imag} */,
  {32'h3f7c45d5, 32'h402f001a} /* (25, 27, 6) {real, imag} */,
  {32'h3fbe5702, 32'h403f9f3b} /* (25, 27, 5) {real, imag} */,
  {32'h3e03a588, 32'h3fe63392} /* (25, 27, 4) {real, imag} */,
  {32'h3eb1869a, 32'h3f088731} /* (25, 27, 3) {real, imag} */,
  {32'h4035152a, 32'h3e8d9931} /* (25, 27, 2) {real, imag} */,
  {32'h3f9706db, 32'h3f1c29b5} /* (25, 27, 1) {real, imag} */,
  {32'hbf87e43b, 32'hbebd82b8} /* (25, 27, 0) {real, imag} */,
  {32'hbf8271a4, 32'hbf96b2bb} /* (25, 26, 31) {real, imag} */,
  {32'hbf5679a6, 32'hbf3730cd} /* (25, 26, 30) {real, imag} */,
  {32'hbe1d76f4, 32'h3e901a9e} /* (25, 26, 29) {real, imag} */,
  {32'h3f411830, 32'hbf53308c} /* (25, 26, 28) {real, imag} */,
  {32'hbd178af0, 32'h3ee1e65c} /* (25, 26, 27) {real, imag} */,
  {32'hbfc45029, 32'hbe3020cc} /* (25, 26, 26) {real, imag} */,
  {32'hbee54b74, 32'hbf959280} /* (25, 26, 25) {real, imag} */,
  {32'h3f179d58, 32'h3fe104bc} /* (25, 26, 24) {real, imag} */,
  {32'hbf89b26c, 32'h3e966fbf} /* (25, 26, 23) {real, imag} */,
  {32'hbe8a5ef3, 32'h3f9d5690} /* (25, 26, 22) {real, imag} */,
  {32'hbea0b800, 32'h3f5b647e} /* (25, 26, 21) {real, imag} */,
  {32'hc00db592, 32'hbf9b5fda} /* (25, 26, 20) {real, imag} */,
  {32'hbf12a808, 32'hbf0f6d68} /* (25, 26, 19) {real, imag} */,
  {32'hbfa24e13, 32'h3ebb5960} /* (25, 26, 18) {real, imag} */,
  {32'hbf87a9c6, 32'hbfb58c38} /* (25, 26, 17) {real, imag} */,
  {32'hbf5fbcf2, 32'hbfea6cfa} /* (25, 26, 16) {real, imag} */,
  {32'h3fccb344, 32'h402abc9c} /* (25, 26, 15) {real, imag} */,
  {32'h404628e2, 32'h3fbaea29} /* (25, 26, 14) {real, imag} */,
  {32'h3eed8266, 32'hbfd0d444} /* (25, 26, 13) {real, imag} */,
  {32'hbf5e8892, 32'hbed1edf2} /* (25, 26, 12) {real, imag} */,
  {32'hbf710c32, 32'h3eac8464} /* (25, 26, 11) {real, imag} */,
  {32'hbf3230d7, 32'h402f9670} /* (25, 26, 10) {real, imag} */,
  {32'h3f64287c, 32'h3fff974e} /* (25, 26, 9) {real, imag} */,
  {32'h3faa3b2c, 32'h3f94966c} /* (25, 26, 8) {real, imag} */,
  {32'h4024933a, 32'h3fd45c72} /* (25, 26, 7) {real, imag} */,
  {32'h4048e5f0, 32'h4003df4e} /* (25, 26, 6) {real, imag} */,
  {32'h3f96a463, 32'h40245661} /* (25, 26, 5) {real, imag} */,
  {32'hbfd135e7, 32'h3f9cc0a0} /* (25, 26, 4) {real, imag} */,
  {32'hbf94779e, 32'h3f0ef7d1} /* (25, 26, 3) {real, imag} */,
  {32'h3feac6ef, 32'h3f540d4c} /* (25, 26, 2) {real, imag} */,
  {32'h3f433e32, 32'h3fb17250} /* (25, 26, 1) {real, imag} */,
  {32'hbf8ea2ac, 32'h3dddff34} /* (25, 26, 0) {real, imag} */,
  {32'h3eae0817, 32'hbf673c9c} /* (25, 25, 31) {real, imag} */,
  {32'hbf6559c6, 32'hbfd3a1de} /* (25, 25, 30) {real, imag} */,
  {32'hbf6f8814, 32'hbfb9f079} /* (25, 25, 29) {real, imag} */,
  {32'h3ea5bf12, 32'h3f150aa0} /* (25, 25, 28) {real, imag} */,
  {32'hbf5c4538, 32'h3f24d1cb} /* (25, 25, 27) {real, imag} */,
  {32'hc02806ae, 32'h3f6be99a} /* (25, 25, 26) {real, imag} */,
  {32'hbfd4d6e4, 32'hbf90a8a2} /* (25, 25, 25) {real, imag} */,
  {32'h3f248f71, 32'h3f1d6cec} /* (25, 25, 24) {real, imag} */,
  {32'h3c22d040, 32'h3fda53ca} /* (25, 25, 23) {real, imag} */,
  {32'h3e2df1d8, 32'h3f965320} /* (25, 25, 22) {real, imag} */,
  {32'hc0083f15, 32'h3fb56e96} /* (25, 25, 21) {real, imag} */,
  {32'hbee5e020, 32'h3fb87af1} /* (25, 25, 20) {real, imag} */,
  {32'h401196df, 32'h3e5f4d4c} /* (25, 25, 19) {real, imag} */,
  {32'hbe132932, 32'h3e496fb8} /* (25, 25, 18) {real, imag} */,
  {32'h3fb1d3a8, 32'hbf7d2f3a} /* (25, 25, 17) {real, imag} */,
  {32'h3fadf4a0, 32'hc036ccab} /* (25, 25, 16) {real, imag} */,
  {32'h3ea31978, 32'h3dc0448c} /* (25, 25, 15) {real, imag} */,
  {32'h3dde6c78, 32'h4005c2b2} /* (25, 25, 14) {real, imag} */,
  {32'hbf3b9950, 32'h3f75dd89} /* (25, 25, 13) {real, imag} */,
  {32'hbf550070, 32'hbf76c0e6} /* (25, 25, 12) {real, imag} */,
  {32'hbf5d5dba, 32'h3f671d05} /* (25, 25, 11) {real, imag} */,
  {32'hbf580836, 32'h4031d176} /* (25, 25, 10) {real, imag} */,
  {32'hbe2b0f78, 32'h3efc55ca} /* (25, 25, 9) {real, imag} */,
  {32'hbfd2d146, 32'hbf40bac4} /* (25, 25, 8) {real, imag} */,
  {32'hbebee08a, 32'hbe85fef7} /* (25, 25, 7) {real, imag} */,
  {32'h4046216e, 32'h40022b38} /* (25, 25, 6) {real, imag} */,
  {32'h400e8301, 32'h402f77cb} /* (25, 25, 5) {real, imag} */,
  {32'hbf9bff70, 32'h3f24b117} /* (25, 25, 4) {real, imag} */,
  {32'hbf8c2c25, 32'h3e68993a} /* (25, 25, 3) {real, imag} */,
  {32'hbf3d3af6, 32'h3fc26885} /* (25, 25, 2) {real, imag} */,
  {32'h3f72d158, 32'h3fb97679} /* (25, 25, 1) {real, imag} */,
  {32'h3fb18062, 32'hbf3eecf1} /* (25, 25, 0) {real, imag} */,
  {32'h3e32f0f1, 32'hbea2eb0c} /* (25, 24, 31) {real, imag} */,
  {32'hbe830478, 32'h3e92ae9b} /* (25, 24, 30) {real, imag} */,
  {32'hbfd5426b, 32'hbe2d43c0} /* (25, 24, 29) {real, imag} */,
  {32'hbfb1b37f, 32'h4014ead8} /* (25, 24, 28) {real, imag} */,
  {32'hbfa7de1c, 32'h3f984618} /* (25, 24, 27) {real, imag} */,
  {32'hbf747451, 32'hbec0989a} /* (25, 24, 26) {real, imag} */,
  {32'hbf485845, 32'hbe5a0176} /* (25, 24, 25) {real, imag} */,
  {32'h3f95ef69, 32'hbf135375} /* (25, 24, 24) {real, imag} */,
  {32'h3fb96a6a, 32'h3f2d6d62} /* (25, 24, 23) {real, imag} */,
  {32'h3dea4e10, 32'h3f80e666} /* (25, 24, 22) {real, imag} */,
  {32'hbedff3c9, 32'h3efc782a} /* (25, 24, 21) {real, imag} */,
  {32'h40162fbe, 32'hbf5479ff} /* (25, 24, 20) {real, imag} */,
  {32'h3fef54e3, 32'hbff741b1} /* (25, 24, 19) {real, imag} */,
  {32'h3fb64789, 32'hbf8486a0} /* (25, 24, 18) {real, imag} */,
  {32'h4065eb98, 32'hbf826482} /* (25, 24, 17) {real, imag} */,
  {32'h3fb5d904, 32'hbfb66eee} /* (25, 24, 16) {real, imag} */,
  {32'hbfadf8ec, 32'hbf0c40f0} /* (25, 24, 15) {real, imag} */,
  {32'hbf938944, 32'h3f5dad46} /* (25, 24, 14) {real, imag} */,
  {32'hbf3095f0, 32'h3fa3a8c3} /* (25, 24, 13) {real, imag} */,
  {32'hc0863dbc, 32'h3f4e183d} /* (25, 24, 12) {real, imag} */,
  {32'hc02edfea, 32'h3f19f6b7} /* (25, 24, 11) {real, imag} */,
  {32'h3f96d64a, 32'h3f396b44} /* (25, 24, 10) {real, imag} */,
  {32'h3f7f82db, 32'hbfbe6ba4} /* (25, 24, 9) {real, imag} */,
  {32'hbf3eea9d, 32'h3da885a0} /* (25, 24, 8) {real, imag} */,
  {32'hbf2d4110, 32'h3fd533e6} /* (25, 24, 7) {real, imag} */,
  {32'h3ff1d04a, 32'h40284914} /* (25, 24, 6) {real, imag} */,
  {32'h3fdb9ac0, 32'h3fe70aa0} /* (25, 24, 5) {real, imag} */,
  {32'h3f1dd20e, 32'h3f19abce} /* (25, 24, 4) {real, imag} */,
  {32'hbdb45430, 32'h3f949132} /* (25, 24, 3) {real, imag} */,
  {32'hbf46711f, 32'h3fe215c4} /* (25, 24, 2) {real, imag} */,
  {32'h402decef, 32'h3f6c09c6} /* (25, 24, 1) {real, imag} */,
  {32'h3fd59f2e, 32'hbe943bde} /* (25, 24, 0) {real, imag} */,
  {32'hbf78a0db, 32'h3ee09a7e} /* (25, 23, 31) {real, imag} */,
  {32'hbf173140, 32'h3eed7677} /* (25, 23, 30) {real, imag} */,
  {32'h3efb5014, 32'h3fb19657} /* (25, 23, 29) {real, imag} */,
  {32'hbe057e40, 32'h400eae75} /* (25, 23, 28) {real, imag} */,
  {32'h3d6c3dc8, 32'h3f4afbb6} /* (25, 23, 27) {real, imag} */,
  {32'h3f9841e6, 32'h3f8d9c0a} /* (25, 23, 26) {real, imag} */,
  {32'h3f0f4760, 32'h3f95f9c8} /* (25, 23, 25) {real, imag} */,
  {32'h3f84e5bc, 32'hbf29e91c} /* (25, 23, 24) {real, imag} */,
  {32'h3fa4a017, 32'hc0192aa2} /* (25, 23, 23) {real, imag} */,
  {32'h3ec5e244, 32'hbfd46b80} /* (25, 23, 22) {real, imag} */,
  {32'h3f945588, 32'hbf640990} /* (25, 23, 21) {real, imag} */,
  {32'h3d169620, 32'hbfa36fb9} /* (25, 23, 20) {real, imag} */,
  {32'h3f81877a, 32'hbe026a36} /* (25, 23, 19) {real, imag} */,
  {32'h3ffeb2c0, 32'hbefb522d} /* (25, 23, 18) {real, imag} */,
  {32'h401040af, 32'hbfe23fc2} /* (25, 23, 17) {real, imag} */,
  {32'h3f5b814f, 32'hbf4a09c2} /* (25, 23, 16) {real, imag} */,
  {32'hbfde2f6f, 32'h3ec475a4} /* (25, 23, 15) {real, imag} */,
  {32'hbf888d71, 32'h401d96d8} /* (25, 23, 14) {real, imag} */,
  {32'hbf87ba68, 32'h3fef7971} /* (25, 23, 13) {real, imag} */,
  {32'hbff404d2, 32'h3f959064} /* (25, 23, 12) {real, imag} */,
  {32'hbfa08bfe, 32'h3f7de26c} /* (25, 23, 11) {real, imag} */,
  {32'h3fd7f2cf, 32'hbea2538c} /* (25, 23, 10) {real, imag} */,
  {32'h3ff268eb, 32'h3e2e519f} /* (25, 23, 9) {real, imag} */,
  {32'h3f18c320, 32'h3f6b0fee} /* (25, 23, 8) {real, imag} */,
  {32'hbf474aba, 32'h3f8577c1} /* (25, 23, 7) {real, imag} */,
  {32'h3f17520c, 32'h3fea58a1} /* (25, 23, 6) {real, imag} */,
  {32'h3fd41ece, 32'h3ff09530} /* (25, 23, 5) {real, imag} */,
  {32'hbe81ff28, 32'h3f8d6552} /* (25, 23, 4) {real, imag} */,
  {32'hbed6a758, 32'h400b9490} /* (25, 23, 3) {real, imag} */,
  {32'h3f16657d, 32'hbf233aea} /* (25, 23, 2) {real, imag} */,
  {32'h4034314c, 32'hbfde341d} /* (25, 23, 1) {real, imag} */,
  {32'h3f407d46, 32'hbf26c838} /* (25, 23, 0) {real, imag} */,
  {32'h3fb79b7d, 32'h3e9c2dcf} /* (25, 22, 31) {real, imag} */,
  {32'h40044032, 32'h3fb75af6} /* (25, 22, 30) {real, imag} */,
  {32'h400330c4, 32'h3e191e20} /* (25, 22, 29) {real, imag} */,
  {32'hbe8a2994, 32'h3f92143a} /* (25, 22, 28) {real, imag} */,
  {32'hbf064bb8, 32'h3f9d5864} /* (25, 22, 27) {real, imag} */,
  {32'h3f92a61a, 32'h3f3f10ce} /* (25, 22, 26) {real, imag} */,
  {32'h3e9dc692, 32'h3c6a3100} /* (25, 22, 25) {real, imag} */,
  {32'h3eca997b, 32'hbeabbb56} /* (25, 22, 24) {real, imag} */,
  {32'hbfac1ebc, 32'hbf2dea52} /* (25, 22, 23) {real, imag} */,
  {32'hbfd9f5f3, 32'hbffa2848} /* (25, 22, 22) {real, imag} */,
  {32'h3efcaeec, 32'hbe868811} /* (25, 22, 21) {real, imag} */,
  {32'h3e648d48, 32'h3f05329f} /* (25, 22, 20) {real, imag} */,
  {32'h3f86d549, 32'h4053ab83} /* (25, 22, 19) {real, imag} */,
  {32'hbd845508, 32'h3f9eb66f} /* (25, 22, 18) {real, imag} */,
  {32'h3fd87ada, 32'hbf06411e} /* (25, 22, 17) {real, imag} */,
  {32'h40225285, 32'h3ee6583a} /* (25, 22, 16) {real, imag} */,
  {32'hbee0885c, 32'hbf5918fe} /* (25, 22, 15) {real, imag} */,
  {32'hbfd67223, 32'h3f7a4cfa} /* (25, 22, 14) {real, imag} */,
  {32'hbffa01d7, 32'h3fddc95a} /* (25, 22, 13) {real, imag} */,
  {32'h3f56c312, 32'h3fb46c18} /* (25, 22, 12) {real, imag} */,
  {32'h3f8350d6, 32'h3dbaf130} /* (25, 22, 11) {real, imag} */,
  {32'h3df4843c, 32'hbfbb5dc6} /* (25, 22, 10) {real, imag} */,
  {32'h3c8c4140, 32'hc018dc78} /* (25, 22, 9) {real, imag} */,
  {32'h3f20379e, 32'hbf52fce8} /* (25, 22, 8) {real, imag} */,
  {32'h3e2f2668, 32'hbfc3deed} /* (25, 22, 7) {real, imag} */,
  {32'h3d8398f8, 32'h3f8aa682} /* (25, 22, 6) {real, imag} */,
  {32'h3ff2b544, 32'h3fef11d5} /* (25, 22, 5) {real, imag} */,
  {32'h3f9f4452, 32'h3e1f418c} /* (25, 22, 4) {real, imag} */,
  {32'h4012a1a6, 32'hbf4d81dc} /* (25, 22, 3) {real, imag} */,
  {32'h3fc62a98, 32'hbfbe6c8c} /* (25, 22, 2) {real, imag} */,
  {32'h3f40abb6, 32'hbe4027e8} /* (25, 22, 1) {real, imag} */,
  {32'h3e940b43, 32'hbf2844d5} /* (25, 22, 0) {real, imag} */,
  {32'h3f7704f1, 32'hbf7f7e55} /* (25, 21, 31) {real, imag} */,
  {32'hbc68e3e0, 32'h3f34cca6} /* (25, 21, 30) {real, imag} */,
  {32'hbfb5601e, 32'h3f2f10ba} /* (25, 21, 29) {real, imag} */,
  {32'hc045af35, 32'h3f766773} /* (25, 21, 28) {real, imag} */,
  {32'hbf8f2b34, 32'h40248de5} /* (25, 21, 27) {real, imag} */,
  {32'hbe966e08, 32'h3fc04564} /* (25, 21, 26) {real, imag} */,
  {32'hbfb908d4, 32'hbf02fddd} /* (25, 21, 25) {real, imag} */,
  {32'h3e023c74, 32'hbdb45410} /* (25, 21, 24) {real, imag} */,
  {32'h3ea31f15, 32'h3f8c3a7f} /* (25, 21, 23) {real, imag} */,
  {32'h3e28df90, 32'h3fa5d5ec} /* (25, 21, 22) {real, imag} */,
  {32'h3ec6d2d7, 32'h3fbe8fff} /* (25, 21, 21) {real, imag} */,
  {32'h3ffa4ab0, 32'hbf2c8c09} /* (25, 21, 20) {real, imag} */,
  {32'h3ffb3b9c, 32'h3f5f1250} /* (25, 21, 19) {real, imag} */,
  {32'h3fad7c34, 32'h3f58d5e6} /* (25, 21, 18) {real, imag} */,
  {32'h3f9e8ad8, 32'h3e93a452} /* (25, 21, 17) {real, imag} */,
  {32'h3eaea62a, 32'h3f52b81f} /* (25, 21, 16) {real, imag} */,
  {32'hbe46df90, 32'hbd129c88} /* (25, 21, 15) {real, imag} */,
  {32'h3f0d37a6, 32'h3f1d17ff} /* (25, 21, 14) {real, imag} */,
  {32'h3fbabc8e, 32'hbe231d98} /* (25, 21, 13) {real, imag} */,
  {32'h3f61b892, 32'h3e85c28c} /* (25, 21, 12) {real, imag} */,
  {32'hbda45be0, 32'hbcfd1240} /* (25, 21, 11) {real, imag} */,
  {32'h3e9a07e6, 32'hbfbedee2} /* (25, 21, 10) {real, imag} */,
  {32'h403ac5e1, 32'hc03b4f77} /* (25, 21, 9) {real, imag} */,
  {32'h401f3784, 32'hbfd12052} /* (25, 21, 8) {real, imag} */,
  {32'hbed8b152, 32'hbfc66819} /* (25, 21, 7) {real, imag} */,
  {32'hbfaf6e34, 32'hbdba2e3c} /* (25, 21, 6) {real, imag} */,
  {32'h3f5958c5, 32'hbef528f5} /* (25, 21, 5) {real, imag} */,
  {32'h3f329604, 32'hbf40f4bc} /* (25, 21, 4) {real, imag} */,
  {32'h4003a2fa, 32'hbf9956d4} /* (25, 21, 3) {real, imag} */,
  {32'h3f0b2238, 32'hbfb208b9} /* (25, 21, 2) {real, imag} */,
  {32'hbe8ae62b, 32'h3fab5e90} /* (25, 21, 1) {real, imag} */,
  {32'hbd5f0488, 32'h3f6df0fe} /* (25, 21, 0) {real, imag} */,
  {32'h3ec222f2, 32'hbe814846} /* (25, 20, 31) {real, imag} */,
  {32'h3f2d28d4, 32'h3f4b0ffe} /* (25, 20, 30) {real, imag} */,
  {32'hbfaf6f0a, 32'h3f3c8b9a} /* (25, 20, 29) {real, imag} */,
  {32'hc033b117, 32'h3eeb0f86} /* (25, 20, 28) {real, imag} */,
  {32'hbfc05aca, 32'h3fe53bd4} /* (25, 20, 27) {real, imag} */,
  {32'hbf81afae, 32'h3f91f7f2} /* (25, 20, 26) {real, imag} */,
  {32'hbfab99ff, 32'hc00c4c82} /* (25, 20, 25) {real, imag} */,
  {32'h3fbc662b, 32'hbfedfc05} /* (25, 20, 24) {real, imag} */,
  {32'h401ac61a, 32'h3f966456} /* (25, 20, 23) {real, imag} */,
  {32'h3f852a74, 32'h40505892} /* (25, 20, 22) {real, imag} */,
  {32'h3ed077a8, 32'h407287af} /* (25, 20, 21) {real, imag} */,
  {32'h3ff5bde2, 32'h3fd7fe67} /* (25, 20, 20) {real, imag} */,
  {32'h3f9108dd, 32'hbeb84738} /* (25, 20, 19) {real, imag} */,
  {32'h3f3ef7b0, 32'hbf45c61e} /* (25, 20, 18) {real, imag} */,
  {32'hbeb3e832, 32'hbed1ee4c} /* (25, 20, 17) {real, imag} */,
  {32'h3e924a30, 32'h3f97f314} /* (25, 20, 16) {real, imag} */,
  {32'h3f674a81, 32'h3eaa48fa} /* (25, 20, 15) {real, imag} */,
  {32'h3fe8b48e, 32'h3fa969f5} /* (25, 20, 14) {real, imag} */,
  {32'h3fb0d3c4, 32'h3ebc009e} /* (25, 20, 13) {real, imag} */,
  {32'h3f4eda6e, 32'h3f0e40d8} /* (25, 20, 12) {real, imag} */,
  {32'h401a3857, 32'hbee4d320} /* (25, 20, 11) {real, imag} */,
  {32'h403ed83b, 32'hbfb9b1f4} /* (25, 20, 10) {real, imag} */,
  {32'h4054ccb9, 32'hbe8cd5d4} /* (25, 20, 9) {real, imag} */,
  {32'h400af2fa, 32'hbe84ff60} /* (25, 20, 8) {real, imag} */,
  {32'h3ed64a30, 32'h3de49c50} /* (25, 20, 7) {real, imag} */,
  {32'hbe85441e, 32'h3f52c06c} /* (25, 20, 6) {real, imag} */,
  {32'h3f1bc1b7, 32'hbf891c49} /* (25, 20, 5) {real, imag} */,
  {32'h3f689508, 32'hbe89a6ea} /* (25, 20, 4) {real, imag} */,
  {32'h3f828be0, 32'h3e841184} /* (25, 20, 3) {real, imag} */,
  {32'hbf5b6649, 32'h3f0d8fa1} /* (25, 20, 2) {real, imag} */,
  {32'h3e3fac8c, 32'h3f8289b3} /* (25, 20, 1) {real, imag} */,
  {32'hbdc37548, 32'h3f93f738} /* (25, 20, 0) {real, imag} */,
  {32'hbe0327d6, 32'hbeaeb760} /* (25, 19, 31) {real, imag} */,
  {32'h3fc6bf03, 32'hbd899b40} /* (25, 19, 30) {real, imag} */,
  {32'hbe0926d8, 32'hbed454da} /* (25, 19, 29) {real, imag} */,
  {32'hbf94f579, 32'h3e68239c} /* (25, 19, 28) {real, imag} */,
  {32'hc01ee5f7, 32'h3ed7437e} /* (25, 19, 27) {real, imag} */,
  {32'hbfd76a66, 32'h3f040031} /* (25, 19, 26) {real, imag} */,
  {32'hbe1c66f6, 32'hbfe8c48c} /* (25, 19, 25) {real, imag} */,
  {32'hbebd5839, 32'hbf4b04b0} /* (25, 19, 24) {real, imag} */,
  {32'hbfab45f9, 32'h3fce82e7} /* (25, 19, 23) {real, imag} */,
  {32'hbf2aec00, 32'h3fa7a7da} /* (25, 19, 22) {real, imag} */,
  {32'h3e241f80, 32'h404571ca} /* (25, 19, 21) {real, imag} */,
  {32'h3f499a6c, 32'h3f4831e5} /* (25, 19, 20) {real, imag} */,
  {32'h3f2de360, 32'hbfc010ed} /* (25, 19, 19) {real, imag} */,
  {32'h3f0f90a7, 32'hbfc76e4c} /* (25, 19, 18) {real, imag} */,
  {32'hbfa3449a, 32'h3f737270} /* (25, 19, 17) {real, imag} */,
  {32'h3e98b592, 32'h3ebc3571} /* (25, 19, 16) {real, imag} */,
  {32'h3f944889, 32'hbe1e1e26} /* (25, 19, 15) {real, imag} */,
  {32'h3f96cd84, 32'h3f2649e8} /* (25, 19, 14) {real, imag} */,
  {32'h3f1ff8c3, 32'h3f7df400} /* (25, 19, 13) {real, imag} */,
  {32'h3f166947, 32'h3fdc71d4} /* (25, 19, 12) {real, imag} */,
  {32'h3f5db09f, 32'hbf0531fe} /* (25, 19, 11) {real, imag} */,
  {32'h3e8f6176, 32'h3f2ea5ad} /* (25, 19, 10) {real, imag} */,
  {32'h3fd78390, 32'h404aedd5} /* (25, 19, 9) {real, imag} */,
  {32'h3fbdf997, 32'h3ff47783} /* (25, 19, 8) {real, imag} */,
  {32'h3f93e592, 32'h3fb2fbb4} /* (25, 19, 7) {real, imag} */,
  {32'h3e7a9cd8, 32'h3f900f4e} /* (25, 19, 6) {real, imag} */,
  {32'h3f387c69, 32'hbf5034ec} /* (25, 19, 5) {real, imag} */,
  {32'h404ddeb4, 32'hbe5468f6} /* (25, 19, 4) {real, imag} */,
  {32'h3f138393, 32'h3ff78acc} /* (25, 19, 3) {real, imag} */,
  {32'hbfad7c7e, 32'h3f93ae00} /* (25, 19, 2) {real, imag} */,
  {32'h3f316a51, 32'h3ef0a88a} /* (25, 19, 1) {real, imag} */,
  {32'h3e0c5e08, 32'hbedcfe07} /* (25, 19, 0) {real, imag} */,
  {32'h3f591882, 32'h3d9eac40} /* (25, 18, 31) {real, imag} */,
  {32'h401f86bb, 32'hbdaf22a4} /* (25, 18, 30) {real, imag} */,
  {32'h3f552fc8, 32'hbfa1b477} /* (25, 18, 29) {real, imag} */,
  {32'hbebf60f4, 32'hc02c19f8} /* (25, 18, 28) {real, imag} */,
  {32'hc029a9bd, 32'hbf99d8b2} /* (25, 18, 27) {real, imag} */,
  {32'hc04b5265, 32'hbf13d1d1} /* (25, 18, 26) {real, imag} */,
  {32'hbff91306, 32'h3e7b1ca4} /* (25, 18, 25) {real, imag} */,
  {32'hc044cf5c, 32'h3fb87e2b} /* (25, 18, 24) {real, imag} */,
  {32'hc049fa00, 32'h3fa51650} /* (25, 18, 23) {real, imag} */,
  {32'hbf858d7b, 32'h3f0d1ee4} /* (25, 18, 22) {real, imag} */,
  {32'h3dd732f0, 32'h3fa4f357} /* (25, 18, 21) {real, imag} */,
  {32'h3e1d2358, 32'h3e64d230} /* (25, 18, 20) {real, imag} */,
  {32'hbf237c08, 32'h3cdd5a50} /* (25, 18, 19) {real, imag} */,
  {32'h3ed19d68, 32'h3f9b72d2} /* (25, 18, 18) {real, imag} */,
  {32'h3e2b97b0, 32'h3e4e926e} /* (25, 18, 17) {real, imag} */,
  {32'h40051237, 32'hbd7d7640} /* (25, 18, 16) {real, imag} */,
  {32'h3f9d29e2, 32'h3f70d016} /* (25, 18, 15) {real, imag} */,
  {32'hbf83620e, 32'hbe88fc74} /* (25, 18, 14) {real, imag} */,
  {32'h3e362948, 32'h3fd23ae8} /* (25, 18, 13) {real, imag} */,
  {32'hbf0d9780, 32'h40059b16} /* (25, 18, 12) {real, imag} */,
  {32'hbf4d9680, 32'h3facf886} /* (25, 18, 11) {real, imag} */,
  {32'h3f02a132, 32'h4010a3ef} /* (25, 18, 10) {real, imag} */,
  {32'h3fc627c8, 32'hbe694508} /* (25, 18, 9) {real, imag} */,
  {32'h3ecc4778, 32'hc0092811} /* (25, 18, 8) {real, imag} */,
  {32'h3fb46214, 32'hbfca458e} /* (25, 18, 7) {real, imag} */,
  {32'hbea992e2, 32'hbf2c3ee2} /* (25, 18, 6) {real, imag} */,
  {32'hbf995c68, 32'hbe4b4350} /* (25, 18, 5) {real, imag} */,
  {32'h3f39d7a2, 32'hbda2c700} /* (25, 18, 4) {real, imag} */,
  {32'h3f4dbd54, 32'h3f797c72} /* (25, 18, 3) {real, imag} */,
  {32'hbf45d323, 32'hbed38b6c} /* (25, 18, 2) {real, imag} */,
  {32'hbf003dde, 32'hbda9a9e0} /* (25, 18, 1) {real, imag} */,
  {32'hbeb20614, 32'h3edbd9f6} /* (25, 18, 0) {real, imag} */,
  {32'h3fac5102, 32'h3f78a39c} /* (25, 17, 31) {real, imag} */,
  {32'h3fc2ef7c, 32'h3f06695a} /* (25, 17, 30) {real, imag} */,
  {32'hbfa75b46, 32'hbd0b24b0} /* (25, 17, 29) {real, imag} */,
  {32'hbf6cb1a1, 32'hbf030276} /* (25, 17, 28) {real, imag} */,
  {32'hc01ab8f5, 32'hbf1087d8} /* (25, 17, 27) {real, imag} */,
  {32'hc068d566, 32'hc0390f91} /* (25, 17, 26) {real, imag} */,
  {32'hc039c38e, 32'hbfb90d3c} /* (25, 17, 25) {real, imag} */,
  {32'hc064b788, 32'h3e2d3ad0} /* (25, 17, 24) {real, imag} */,
  {32'hc045d406, 32'h3f05241e} /* (25, 17, 23) {real, imag} */,
  {32'hbfe44125, 32'h3ef39964} /* (25, 17, 22) {real, imag} */,
  {32'hbec8f662, 32'hbfc6a2ea} /* (25, 17, 21) {real, imag} */,
  {32'h3edda1be, 32'h3d995bdc} /* (25, 17, 20) {real, imag} */,
  {32'h3dc45f6a, 32'h40214f6b} /* (25, 17, 19) {real, imag} */,
  {32'h3ee82634, 32'h405ef112} /* (25, 17, 18) {real, imag} */,
  {32'h3fa54513, 32'h3fb54a43} /* (25, 17, 17) {real, imag} */,
  {32'h3fcafccd, 32'hbbf2d580} /* (25, 17, 16) {real, imag} */,
  {32'hbfb3edf2, 32'h3f17213a} /* (25, 17, 15) {real, imag} */,
  {32'hbf278b24, 32'h3fb2d56c} /* (25, 17, 14) {real, imag} */,
  {32'h3e1815b8, 32'h402899c0} /* (25, 17, 13) {real, imag} */,
  {32'hc05729df, 32'h401cbda8} /* (25, 17, 12) {real, imag} */,
  {32'hbfcee157, 32'h3e8fe206} /* (25, 17, 11) {real, imag} */,
  {32'h3f53d424, 32'hc012f904} /* (25, 17, 10) {real, imag} */,
  {32'h3e5030f0, 32'hc025f8f9} /* (25, 17, 9) {real, imag} */,
  {32'hbf628548, 32'hbfd98a48} /* (25, 17, 8) {real, imag} */,
  {32'hbf77b0ee, 32'hc0438266} /* (25, 17, 7) {real, imag} */,
  {32'hbfa16202, 32'hbf985e95} /* (25, 17, 6) {real, imag} */,
  {32'hbfd32582, 32'hbf5f93ee} /* (25, 17, 5) {real, imag} */,
  {32'hbd14c9e8, 32'hbf141444} /* (25, 17, 4) {real, imag} */,
  {32'h3fc9f370, 32'hbd499990} /* (25, 17, 3) {real, imag} */,
  {32'h3e6704ca, 32'hbeff71ea} /* (25, 17, 2) {real, imag} */,
  {32'hbf09aebc, 32'h3efec35c} /* (25, 17, 1) {real, imag} */,
  {32'h3dd1f0a0, 32'h3f886876} /* (25, 17, 0) {real, imag} */,
  {32'hbee2895d, 32'h3fa77912} /* (25, 16, 31) {real, imag} */,
  {32'h3d92f3a0, 32'hbf2bbb46} /* (25, 16, 30) {real, imag} */,
  {32'h3e9716ac, 32'hbe90bc58} /* (25, 16, 29) {real, imag} */,
  {32'hbf944950, 32'h3d8ff4c0} /* (25, 16, 28) {real, imag} */,
  {32'h3f3788a0, 32'hbfc25461} /* (25, 16, 27) {real, imag} */,
  {32'h3e06f830, 32'hc022b70f} /* (25, 16, 26) {real, imag} */,
  {32'h3f48862a, 32'hbfa44fd3} /* (25, 16, 25) {real, imag} */,
  {32'h3f9e63df, 32'hbf357a39} /* (25, 16, 24) {real, imag} */,
  {32'hbf1f6200, 32'hbdb122c0} /* (25, 16, 23) {real, imag} */,
  {32'hbef7a89c, 32'h3f8241c1} /* (25, 16, 22) {real, imag} */,
  {32'hbd247e40, 32'hbf80c6da} /* (25, 16, 21) {real, imag} */,
  {32'h3eeeed98, 32'hbe9f9f60} /* (25, 16, 20) {real, imag} */,
  {32'hbcdfd2c0, 32'h401341d2} /* (25, 16, 19) {real, imag} */,
  {32'hbdf21af8, 32'h404b908d} /* (25, 16, 18) {real, imag} */,
  {32'h3fcfb7c4, 32'h3fc6aac2} /* (25, 16, 17) {real, imag} */,
  {32'h3e2817fc, 32'h3f5af5f4} /* (25, 16, 16) {real, imag} */,
  {32'hbfab79df, 32'h3f9a4ce4} /* (25, 16, 15) {real, imag} */,
  {32'h3f37f543, 32'h3f9c3e24} /* (25, 16, 14) {real, imag} */,
  {32'h3e98a534, 32'h400c6d12} /* (25, 16, 13) {real, imag} */,
  {32'hbf14a69a, 32'hbf0d827f} /* (25, 16, 12) {real, imag} */,
  {32'h3ff15dfa, 32'hbd7c5d20} /* (25, 16, 11) {real, imag} */,
  {32'h3fdc8e32, 32'hbf3ef707} /* (25, 16, 10) {real, imag} */,
  {32'h403543d5, 32'hbfd35924} /* (25, 16, 9) {real, imag} */,
  {32'h3f85b580, 32'hc04fde76} /* (25, 16, 8) {real, imag} */,
  {32'hbe534aa6, 32'hc03e0bf2} /* (25, 16, 7) {real, imag} */,
  {32'hbfa32644, 32'h3f1e2b96} /* (25, 16, 6) {real, imag} */,
  {32'hbfa87286, 32'h3e4ca8f8} /* (25, 16, 5) {real, imag} */,
  {32'hbf3d466a, 32'hbe612b72} /* (25, 16, 4) {real, imag} */,
  {32'hbf6ac45c, 32'hbf4b7490} /* (25, 16, 3) {real, imag} */,
  {32'hbf271e44, 32'hbfa46ef5} /* (25, 16, 2) {real, imag} */,
  {32'h3fa2e2df, 32'hbf3f08a4} /* (25, 16, 1) {real, imag} */,
  {32'hbea15e60, 32'h3f145322} /* (25, 16, 0) {real, imag} */,
  {32'hbfa9a0b4, 32'h4012969f} /* (25, 15, 31) {real, imag} */,
  {32'hbf56f7c4, 32'h3dd99160} /* (25, 15, 30) {real, imag} */,
  {32'h3f9002fb, 32'h3fc9dd81} /* (25, 15, 29) {real, imag} */,
  {32'h3ef68dd0, 32'h3fb0c0f0} /* (25, 15, 28) {real, imag} */,
  {32'h3ff538d2, 32'hbf85e233} /* (25, 15, 27) {real, imag} */,
  {32'h3fd05509, 32'hc003787b} /* (25, 15, 26) {real, imag} */,
  {32'h3fc78926, 32'hc027a9c8} /* (25, 15, 25) {real, imag} */,
  {32'h3fe980a4, 32'hbfcefad2} /* (25, 15, 24) {real, imag} */,
  {32'hbf8cfbe7, 32'hbfaab764} /* (25, 15, 23) {real, imag} */,
  {32'hbff64801, 32'h3f0f9100} /* (25, 15, 22) {real, imag} */,
  {32'hbfc23ca1, 32'h3ff7fc55} /* (25, 15, 21) {real, imag} */,
  {32'h3f31d427, 32'h40007d3e} /* (25, 15, 20) {real, imag} */,
  {32'h3fb785ed, 32'h3f2b784c} /* (25, 15, 19) {real, imag} */,
  {32'hbd3c1930, 32'h4024a97e} /* (25, 15, 18) {real, imag} */,
  {32'h3fabb40b, 32'h3fd8d066} /* (25, 15, 17) {real, imag} */,
  {32'h3eef0810, 32'h3fefec56} /* (25, 15, 16) {real, imag} */,
  {32'hbfa943c2, 32'h3f6f4f3e} /* (25, 15, 15) {real, imag} */,
  {32'hbfc8f92c, 32'h3eb2916c} /* (25, 15, 14) {real, imag} */,
  {32'hc0475cf4, 32'h3eab1bc7} /* (25, 15, 13) {real, imag} */,
  {32'hbfdcb3f5, 32'h3f419356} /* (25, 15, 12) {real, imag} */,
  {32'h3fc7e146, 32'h3f89f907} /* (25, 15, 11) {real, imag} */,
  {32'h3f6b5fed, 32'hbfa37d5a} /* (25, 15, 10) {real, imag} */,
  {32'h4009a1fb, 32'hc02844ba} /* (25, 15, 9) {real, imag} */,
  {32'h3fc4ebd4, 32'hc01ad136} /* (25, 15, 8) {real, imag} */,
  {32'h3fa1ec3b, 32'hbf6b8f30} /* (25, 15, 7) {real, imag} */,
  {32'h3e85d850, 32'h3f73b258} /* (25, 15, 6) {real, imag} */,
  {32'hbef140ae, 32'h3e87b553} /* (25, 15, 5) {real, imag} */,
  {32'hbededae8, 32'hbef62720} /* (25, 15, 4) {real, imag} */,
  {32'hbfa07f51, 32'hbfa7c76e} /* (25, 15, 3) {real, imag} */,
  {32'hbf555668, 32'hbfb2fc7a} /* (25, 15, 2) {real, imag} */,
  {32'h3ff8cd47, 32'hbf56d6aa} /* (25, 15, 1) {real, imag} */,
  {32'h3f61fb3a, 32'h3da27180} /* (25, 15, 0) {real, imag} */,
  {32'h3ed7daac, 32'h3f03f862} /* (25, 14, 31) {real, imag} */,
  {32'h3e8ad90e, 32'hbe4eed48} /* (25, 14, 30) {real, imag} */,
  {32'h3ed68232, 32'hc0074a5d} /* (25, 14, 29) {real, imag} */,
  {32'h3f371491, 32'hbec28e6f} /* (25, 14, 28) {real, imag} */,
  {32'hbf80558a, 32'h3f418346} /* (25, 14, 27) {real, imag} */,
  {32'h3e72f064, 32'hbf9a747e} /* (25, 14, 26) {real, imag} */,
  {32'h3fa3d306, 32'hc007e594} /* (25, 14, 25) {real, imag} */,
  {32'h3fe13bc6, 32'hbfac1123} /* (25, 14, 24) {real, imag} */,
  {32'h3f5d19f6, 32'hbf37fe08} /* (25, 14, 23) {real, imag} */,
  {32'h3f6607e2, 32'hbf3437bc} /* (25, 14, 22) {real, imag} */,
  {32'h3f277d26, 32'hbf167704} /* (25, 14, 21) {real, imag} */,
  {32'hbf291b7c, 32'h3ee952bc} /* (25, 14, 20) {real, imag} */,
  {32'h3f708766, 32'h3f322ba5} /* (25, 14, 19) {real, imag} */,
  {32'hbe64743c, 32'h3ffe0b3c} /* (25, 14, 18) {real, imag} */,
  {32'hbf30454f, 32'h3f195d74} /* (25, 14, 17) {real, imag} */,
  {32'h3f74a05b, 32'h3fa06f82} /* (25, 14, 16) {real, imag} */,
  {32'hbfbfe443, 32'h3f5a705f} /* (25, 14, 15) {real, imag} */,
  {32'hbfcaa908, 32'h3f7dcf16} /* (25, 14, 14) {real, imag} */,
  {32'h3eb767b6, 32'h3f9a7e3c} /* (25, 14, 13) {real, imag} */,
  {32'h3f109198, 32'h400bb12c} /* (25, 14, 12) {real, imag} */,
  {32'h3f931382, 32'h3f9d8624} /* (25, 14, 11) {real, imag} */,
  {32'h3ee0e6b9, 32'hbfdff212} /* (25, 14, 10) {real, imag} */,
  {32'h3fbd4cc6, 32'hbfe50055} /* (25, 14, 9) {real, imag} */,
  {32'h3fc56750, 32'h3f52a536} /* (25, 14, 8) {real, imag} */,
  {32'h400b3749, 32'h3df53f50} /* (25, 14, 7) {real, imag} */,
  {32'h3fc59064, 32'hbe32f4ce} /* (25, 14, 6) {real, imag} */,
  {32'h3f1714f6, 32'h3f432c5c} /* (25, 14, 5) {real, imag} */,
  {32'hbcbe86c8, 32'hbebf2dd9} /* (25, 14, 4) {real, imag} */,
  {32'hbf40e5d6, 32'hbff34a10} /* (25, 14, 3) {real, imag} */,
  {32'hbfe3a70e, 32'hbfea2489} /* (25, 14, 2) {real, imag} */,
  {32'hbf31ea8a, 32'hc013bf20} /* (25, 14, 1) {real, imag} */,
  {32'h3fddfd76, 32'hbfcd4a2a} /* (25, 14, 0) {real, imag} */,
  {32'h3ee55966, 32'hbedc98bc} /* (25, 13, 31) {real, imag} */,
  {32'hbf1ce290, 32'hbd089358} /* (25, 13, 30) {real, imag} */,
  {32'hbf2fd704, 32'hbf0dc15b} /* (25, 13, 29) {real, imag} */,
  {32'h3f3ff07c, 32'h3f2be2e6} /* (25, 13, 28) {real, imag} */,
  {32'hbe851e2a, 32'h3fcbec6c} /* (25, 13, 27) {real, imag} */,
  {32'hbea37e10, 32'hbeaba59e} /* (25, 13, 26) {real, imag} */,
  {32'h3f27a74b, 32'hc0042f6a} /* (25, 13, 25) {real, imag} */,
  {32'h3f36e286, 32'hbf202168} /* (25, 13, 24) {real, imag} */,
  {32'h3fbe2006, 32'h3f6cf9da} /* (25, 13, 23) {real, imag} */,
  {32'h4038a7e8, 32'hbf3a45ba} /* (25, 13, 22) {real, imag} */,
  {32'h404f1cae, 32'hbf58825a} /* (25, 13, 21) {real, imag} */,
  {32'hbf7a976c, 32'hbf77c6b2} /* (25, 13, 20) {real, imag} */,
  {32'hc01b9520, 32'h3fe76fba} /* (25, 13, 19) {real, imag} */,
  {32'hbfff794f, 32'h3f9fe219} /* (25, 13, 18) {real, imag} */,
  {32'hc0236762, 32'hbd685b00} /* (25, 13, 17) {real, imag} */,
  {32'hbfc1dc93, 32'h3f1c8eb6} /* (25, 13, 16) {real, imag} */,
  {32'hbf5533c8, 32'hbe646be0} /* (25, 13, 15) {real, imag} */,
  {32'h3e96916d, 32'hbedd9dea} /* (25, 13, 14) {real, imag} */,
  {32'h3f8f5795, 32'h3e0ca5be} /* (25, 13, 13) {real, imag} */,
  {32'h3f78db26, 32'h3f2584b0} /* (25, 13, 12) {real, imag} */,
  {32'h3fd40add, 32'hbf7ec947} /* (25, 13, 11) {real, imag} */,
  {32'h3df88b98, 32'hc035b3e6} /* (25, 13, 10) {real, imag} */,
  {32'h3e16b5c0, 32'hbfc908ef} /* (25, 13, 9) {real, imag} */,
  {32'hbe9c5454, 32'h3e761ff8} /* (25, 13, 8) {real, imag} */,
  {32'hbf083280, 32'hbeca2e70} /* (25, 13, 7) {real, imag} */,
  {32'h3fcb547c, 32'hbe1f7d57} /* (25, 13, 6) {real, imag} */,
  {32'h3fcd3a80, 32'h4003538c} /* (25, 13, 5) {real, imag} */,
  {32'hbf16ee16, 32'h3e1fd95c} /* (25, 13, 4) {real, imag} */,
  {32'hbf87f790, 32'hc003ddfe} /* (25, 13, 3) {real, imag} */,
  {32'hbfab7ae7, 32'hbfbd97c0} /* (25, 13, 2) {real, imag} */,
  {32'hbf965c7c, 32'hc0174bb0} /* (25, 13, 1) {real, imag} */,
  {32'h3ecc3b68, 32'hbfdbb972} /* (25, 13, 0) {real, imag} */,
  {32'hbf56da6a, 32'hbf828d10} /* (25, 12, 31) {real, imag} */,
  {32'hc04cc0c0, 32'hbf5e2992} /* (25, 12, 30) {real, imag} */,
  {32'hc0098099, 32'hbeac049e} /* (25, 12, 29) {real, imag} */,
  {32'h3ebd68ac, 32'h40011d48} /* (25, 12, 28) {real, imag} */,
  {32'h3f2169aa, 32'h3fa32672} /* (25, 12, 27) {real, imag} */,
  {32'hbed5440c, 32'h3e98f15c} /* (25, 12, 26) {real, imag} */,
  {32'hbeaabbd8, 32'hbf2ceb6b} /* (25, 12, 25) {real, imag} */,
  {32'hbf96172d, 32'hc0055066} /* (25, 12, 24) {real, imag} */,
  {32'h3d268d50, 32'hbf8f2bdd} /* (25, 12, 23) {real, imag} */,
  {32'h3f3d96cc, 32'hbfc91971} /* (25, 12, 22) {real, imag} */,
  {32'h4027585c, 32'hbf8bc75c} /* (25, 12, 21) {real, imag} */,
  {32'h3fa03c78, 32'h3de1a4b8} /* (25, 12, 20) {real, imag} */,
  {32'hbf484d8e, 32'h4012e7a6} /* (25, 12, 19) {real, imag} */,
  {32'hbeae0928, 32'h3f8f9a32} /* (25, 12, 18) {real, imag} */,
  {32'hc015c328, 32'hbf050404} /* (25, 12, 17) {real, imag} */,
  {32'hc00731eb, 32'h3f87ba5c} /* (25, 12, 16) {real, imag} */,
  {32'h3f4a85d2, 32'hbf925ec7} /* (25, 12, 15) {real, imag} */,
  {32'h3f4e329c, 32'hbe9c25cc} /* (25, 12, 14) {real, imag} */,
  {32'hbf9ea922, 32'h3f6907e6} /* (25, 12, 13) {real, imag} */,
  {32'hbf234118, 32'h3fdffef9} /* (25, 12, 12) {real, imag} */,
  {32'h3f1458e0, 32'hbf9a65ce} /* (25, 12, 11) {real, imag} */,
  {32'hbf3ceb42, 32'hbfa75602} /* (25, 12, 10) {real, imag} */,
  {32'hbf7c7308, 32'h3f7ae16f} /* (25, 12, 9) {real, imag} */,
  {32'h3ea4060c, 32'hbe1c76a0} /* (25, 12, 8) {real, imag} */,
  {32'hbe8e3a34, 32'hbefe8912} /* (25, 12, 7) {real, imag} */,
  {32'h3f907e9b, 32'h3fbd80e8} /* (25, 12, 6) {real, imag} */,
  {32'h4035651b, 32'h3fb44f30} /* (25, 12, 5) {real, imag} */,
  {32'h3ea901d8, 32'hbe871dcf} /* (25, 12, 4) {real, imag} */,
  {32'hbf0b35d1, 32'h3f370c25} /* (25, 12, 3) {real, imag} */,
  {32'hbf7aa316, 32'hbf0e5f57} /* (25, 12, 2) {real, imag} */,
  {32'hbf637af1, 32'hc02023c7} /* (25, 12, 1) {real, imag} */,
  {32'hbeb40b53, 32'hbf994033} /* (25, 12, 0) {real, imag} */,
  {32'hbf71e8cf, 32'hbf040cae} /* (25, 11, 31) {real, imag} */,
  {32'hbfbc1ff2, 32'h3f456cc1} /* (25, 11, 30) {real, imag} */,
  {32'hbfa7ec9f, 32'hbeb8fb16} /* (25, 11, 29) {real, imag} */,
  {32'hbf09db34, 32'h3f8906d2} /* (25, 11, 28) {real, imag} */,
  {32'hbf2f3602, 32'hbd83bb88} /* (25, 11, 27) {real, imag} */,
  {32'h3d3773e0, 32'hbf638189} /* (25, 11, 26) {real, imag} */,
  {32'h3f952231, 32'h3de32b38} /* (25, 11, 25) {real, imag} */,
  {32'hbf3bf695, 32'h3f17e9de} /* (25, 11, 24) {real, imag} */,
  {32'hbe6fff60, 32'hbfaeaa2e} /* (25, 11, 23) {real, imag} */,
  {32'h3fae3351, 32'hbedad5a8} /* (25, 11, 22) {real, imag} */,
  {32'h3f07973e, 32'hbfeaf2f6} /* (25, 11, 21) {real, imag} */,
  {32'hbd968490, 32'hbf8cb838} /* (25, 11, 20) {real, imag} */,
  {32'hbf051f95, 32'h402ac1b0} /* (25, 11, 19) {real, imag} */,
  {32'h3ea80958, 32'h40128a41} /* (25, 11, 18) {real, imag} */,
  {32'hbf2966ff, 32'hbf80877b} /* (25, 11, 17) {real, imag} */,
  {32'hbf8a80fc, 32'h40433ec0} /* (25, 11, 16) {real, imag} */,
  {32'h3deff4e4, 32'h3fe8403c} /* (25, 11, 15) {real, imag} */,
  {32'hbfda3e4f, 32'h3f2c367e} /* (25, 11, 14) {real, imag} */,
  {32'hc00f0bf5, 32'h3f5cb702} /* (25, 11, 13) {real, imag} */,
  {32'hbf1f032e, 32'hbe5a1fe8} /* (25, 11, 12) {real, imag} */,
  {32'h3bb40400, 32'hbe518c18} /* (25, 11, 11) {real, imag} */,
  {32'hbf71eaff, 32'hbfa31589} /* (25, 11, 10) {real, imag} */,
  {32'hbfd980a2, 32'h3c2e7100} /* (25, 11, 9) {real, imag} */,
  {32'hc01a3db8, 32'hbf9abfd2} /* (25, 11, 8) {real, imag} */,
  {32'hc0349e4f, 32'hbf8851e0} /* (25, 11, 7) {real, imag} */,
  {32'hc00e7c50, 32'h3fef984e} /* (25, 11, 6) {real, imag} */,
  {32'h3ebc39e4, 32'hbd1cc900} /* (25, 11, 5) {real, imag} */,
  {32'hbd1bdca8, 32'hc0206ce0} /* (25, 11, 4) {real, imag} */,
  {32'h3f350007, 32'hbfad0cb4} /* (25, 11, 3) {real, imag} */,
  {32'h3e8ab62c, 32'hbfce46ce} /* (25, 11, 2) {real, imag} */,
  {32'h3e946711, 32'hc001e8a2} /* (25, 11, 1) {real, imag} */,
  {32'hbeaae442, 32'hbf15cfe3} /* (25, 11, 0) {real, imag} */,
  {32'h3dbcef4e, 32'hbf085bbd} /* (25, 10, 31) {real, imag} */,
  {32'hbf0276e9, 32'h3f878be8} /* (25, 10, 30) {real, imag} */,
  {32'h3fd07793, 32'h4086ff07} /* (25, 10, 29) {real, imag} */,
  {32'hbf4ddc0a, 32'h3fa03486} /* (25, 10, 28) {real, imag} */,
  {32'hbff1146b, 32'hbdbd4c98} /* (25, 10, 27) {real, imag} */,
  {32'h3fe505a6, 32'hbe8ca096} /* (25, 10, 26) {real, imag} */,
  {32'h3f175ea2, 32'h3f156912} /* (25, 10, 25) {real, imag} */,
  {32'hbf03d49a, 32'h3fac3210} /* (25, 10, 24) {real, imag} */,
  {32'hbfa63862, 32'hbe272b18} /* (25, 10, 23) {real, imag} */,
  {32'h3fb9cac4, 32'h4010e3b8} /* (25, 10, 22) {real, imag} */,
  {32'hbfb6fcd7, 32'h3fa32840} /* (25, 10, 21) {real, imag} */,
  {32'hbff7b1c0, 32'hbfecfe11} /* (25, 10, 20) {real, imag} */,
  {32'hbf6fcc3e, 32'h3f57bda4} /* (25, 10, 19) {real, imag} */,
  {32'hc01095ee, 32'h40190108} /* (25, 10, 18) {real, imag} */,
  {32'hbed67a14, 32'hbf61d735} /* (25, 10, 17) {real, imag} */,
  {32'h3ec6d5ca, 32'h3fed0042} /* (25, 10, 16) {real, imag} */,
  {32'hbe772338, 32'h40752d7e} /* (25, 10, 15) {real, imag} */,
  {32'hbfac447d, 32'h4017b5d8} /* (25, 10, 14) {real, imag} */,
  {32'hbe47fec0, 32'h3ed9df44} /* (25, 10, 13) {real, imag} */,
  {32'h3e525988, 32'hc026fae4} /* (25, 10, 12) {real, imag} */,
  {32'hbf2cf9c4, 32'hbf9ef54e} /* (25, 10, 11) {real, imag} */,
  {32'hc029f9f6, 32'hbf532651} /* (25, 10, 10) {real, imag} */,
  {32'hc00d8558, 32'hbf74b200} /* (25, 10, 9) {real, imag} */,
  {32'hbf9abbea, 32'hbffc684c} /* (25, 10, 8) {real, imag} */,
  {32'hc0832a93, 32'h3eb83d40} /* (25, 10, 7) {real, imag} */,
  {32'hc03cc236, 32'h3f79f9f5} /* (25, 10, 6) {real, imag} */,
  {32'hbf85884e, 32'h3f980344} /* (25, 10, 5) {real, imag} */,
  {32'hbf131bec, 32'h3e83d3a4} /* (25, 10, 4) {real, imag} */,
  {32'h3fb8b905, 32'hbf52c829} /* (25, 10, 3) {real, imag} */,
  {32'h3f701ce2, 32'hbf380373} /* (25, 10, 2) {real, imag} */,
  {32'h3f269a5c, 32'hbf72a5da} /* (25, 10, 1) {real, imag} */,
  {32'h3d072554, 32'h3e935976} /* (25, 10, 0) {real, imag} */,
  {32'h3ea6e190, 32'hbf4e4785} /* (25, 9, 31) {real, imag} */,
  {32'hbfd2d0b2, 32'h3fbc4530} /* (25, 9, 30) {real, imag} */,
  {32'hbf3d0200, 32'h4084d786} /* (25, 9, 29) {real, imag} */,
  {32'hbfdeba38, 32'h3fee691f} /* (25, 9, 28) {real, imag} */,
  {32'hbe38ea84, 32'h3f8c6eed} /* (25, 9, 27) {real, imag} */,
  {32'h3f4c96e8, 32'hbe8f261d} /* (25, 9, 26) {real, imag} */,
  {32'hbf4b359c, 32'hbff165dd} /* (25, 9, 25) {real, imag} */,
  {32'hbf897122, 32'hc01a19e8} /* (25, 9, 24) {real, imag} */,
  {32'hbf9939e4, 32'h3f85592c} /* (25, 9, 23) {real, imag} */,
  {32'h3f3178a6, 32'h402f8dec} /* (25, 9, 22) {real, imag} */,
  {32'h3ec1f42e, 32'h3f53df04} /* (25, 9, 21) {real, imag} */,
  {32'hbfb237e4, 32'hbff27060} /* (25, 9, 20) {real, imag} */,
  {32'hc03d5650, 32'h3e24f2a8} /* (25, 9, 19) {real, imag} */,
  {32'hbffc59c4, 32'h3ecc4434} /* (25, 9, 18) {real, imag} */,
  {32'h3dbb4e50, 32'hbf2b6422} /* (25, 9, 17) {real, imag} */,
  {32'h3f4e2e9a, 32'h3f500bc0} /* (25, 9, 16) {real, imag} */,
  {32'h3f492c93, 32'h40434cae} /* (25, 9, 15) {real, imag} */,
  {32'hbf9668f2, 32'h406a2816} /* (25, 9, 14) {real, imag} */,
  {32'hbd6d20e0, 32'h403e5f33} /* (25, 9, 13) {real, imag} */,
  {32'h3f6488ea, 32'hbe360ce8} /* (25, 9, 12) {real, imag} */,
  {32'h3ecb6bde, 32'hbfd5729e} /* (25, 9, 11) {real, imag} */,
  {32'hbeb4e35c, 32'hbfc0768d} /* (25, 9, 10) {real, imag} */,
  {32'hbe9c5d70, 32'hbf1ccfba} /* (25, 9, 9) {real, imag} */,
  {32'hbf8b6ef6, 32'hbf676122} /* (25, 9, 8) {real, imag} */,
  {32'hc03eb8bc, 32'h3f56aa80} /* (25, 9, 7) {real, imag} */,
  {32'hbebba2b0, 32'h3f69bde0} /* (25, 9, 6) {real, imag} */,
  {32'h3f8d6848, 32'h3ebbbe99} /* (25, 9, 5) {real, imag} */,
  {32'h3f7fcff4, 32'h403010ec} /* (25, 9, 4) {real, imag} */,
  {32'h3f96e160, 32'h4029f073} /* (25, 9, 3) {real, imag} */,
  {32'hbd78ae80, 32'h3ca57780} /* (25, 9, 2) {real, imag} */,
  {32'hbf81b1e4, 32'hbea8a7c3} /* (25, 9, 1) {real, imag} */,
  {32'hbea73632, 32'h3e3a3a98} /* (25, 9, 0) {real, imag} */,
  {32'h3f0b0e56, 32'hbf7abf84} /* (25, 8, 31) {real, imag} */,
  {32'hbfd0ec63, 32'h3ff66896} /* (25, 8, 30) {real, imag} */,
  {32'hbd666b80, 32'h3fd19dc8} /* (25, 8, 29) {real, imag} */,
  {32'hc000122a, 32'h3e359a42} /* (25, 8, 28) {real, imag} */,
  {32'hc001737a, 32'h3f88a9a4} /* (25, 8, 27) {real, imag} */,
  {32'hbf82054e, 32'h3f812153} /* (25, 8, 26) {real, imag} */,
  {32'hbe3e172f, 32'hc00458e8} /* (25, 8, 25) {real, imag} */,
  {32'hbf164ba8, 32'hc085dde6} /* (25, 8, 24) {real, imag} */,
  {32'hbed3a1d8, 32'hbe3c5af8} /* (25, 8, 23) {real, imag} */,
  {32'h3f942633, 32'hbe869308} /* (25, 8, 22) {real, imag} */,
  {32'h3feb7d23, 32'h3f670090} /* (25, 8, 21) {real, imag} */,
  {32'h3f9a50e8, 32'h400cdb71} /* (25, 8, 20) {real, imag} */,
  {32'hbffe02ff, 32'h3f969f5b} /* (25, 8, 19) {real, imag} */,
  {32'hbe91847f, 32'hbf7e56f6} /* (25, 8, 18) {real, imag} */,
  {32'hbd88aa78, 32'h3f065b96} /* (25, 8, 17) {real, imag} */,
  {32'hbf611d04, 32'h3ff14604} /* (25, 8, 16) {real, imag} */,
  {32'h3ebc1994, 32'h405b1157} /* (25, 8, 15) {real, imag} */,
  {32'hbf925db5, 32'h40121aa6} /* (25, 8, 14) {real, imag} */,
  {32'hbfa07e10, 32'h3fad31e0} /* (25, 8, 13) {real, imag} */,
  {32'h3fea8b6f, 32'h3ec67b58} /* (25, 8, 12) {real, imag} */,
  {32'h3ef09620, 32'h3f7190e0} /* (25, 8, 11) {real, imag} */,
  {32'h3f34fb1c, 32'hbb975000} /* (25, 8, 10) {real, imag} */,
  {32'h3ff84add, 32'h3e04adb0} /* (25, 8, 9) {real, imag} */,
  {32'h3e874ec8, 32'h3f6421f0} /* (25, 8, 8) {real, imag} */,
  {32'h3f9ed4af, 32'hbffd7bd0} /* (25, 8, 7) {real, imag} */,
  {32'h3fd9b75e, 32'hbf0f952f} /* (25, 8, 6) {real, imag} */,
  {32'h3fcd75fd, 32'h3faf85f9} /* (25, 8, 5) {real, imag} */,
  {32'hbf0add29, 32'h3fe1e01d} /* (25, 8, 4) {real, imag} */,
  {32'hbf54cb78, 32'h402f13a8} /* (25, 8, 3) {real, imag} */,
  {32'h3eb3e2ec, 32'h3fb5ce5f} /* (25, 8, 2) {real, imag} */,
  {32'h3f945147, 32'h3f3d0a6c} /* (25, 8, 1) {real, imag} */,
  {32'h3ed68cec, 32'h3d040660} /* (25, 8, 0) {real, imag} */,
  {32'hbf3f1ae3, 32'h3f4abea3} /* (25, 7, 31) {real, imag} */,
  {32'hbf17b6ab, 32'h3fe6977a} /* (25, 7, 30) {real, imag} */,
  {32'h403ae15b, 32'h3fa115a3} /* (25, 7, 29) {real, imag} */,
  {32'h3fffd40b, 32'hbe3eaaf4} /* (25, 7, 28) {real, imag} */,
  {32'hbeb5b9fe, 32'h3f0d0913} /* (25, 7, 27) {real, imag} */,
  {32'hbe7deaf4, 32'h403bdbad} /* (25, 7, 26) {real, imag} */,
  {32'hbf0573ba, 32'h3d55dea0} /* (25, 7, 25) {real, imag} */,
  {32'hbe8f6e32, 32'hc037efd4} /* (25, 7, 24) {real, imag} */,
  {32'h3f92ccb5, 32'hbf77d34c} /* (25, 7, 23) {real, imag} */,
  {32'h3fd74811, 32'hbf9859a6} /* (25, 7, 22) {real, imag} */,
  {32'hbe010878, 32'h40074730} /* (25, 7, 21) {real, imag} */,
  {32'hbf2d603c, 32'h409d8d02} /* (25, 7, 20) {real, imag} */,
  {32'h3eed0e46, 32'h3fb67800} /* (25, 7, 19) {real, imag} */,
  {32'h3ffebe02, 32'hbfaa457c} /* (25, 7, 18) {real, imag} */,
  {32'h3e909bea, 32'h3f1e42a6} /* (25, 7, 17) {real, imag} */,
  {32'h3fdccdd1, 32'h3fc06252} /* (25, 7, 16) {real, imag} */,
  {32'h3f8706ce, 32'h3ffa4b62} /* (25, 7, 15) {real, imag} */,
  {32'hbf637307, 32'hbbdebd80} /* (25, 7, 14) {real, imag} */,
  {32'hbfd537df, 32'hbf2312b2} /* (25, 7, 13) {real, imag} */,
  {32'h3f804050, 32'h3d094a00} /* (25, 7, 12) {real, imag} */,
  {32'h3fa2927e, 32'h4002a6e7} /* (25, 7, 11) {real, imag} */,
  {32'hbf24cb62, 32'h3ebaa43c} /* (25, 7, 10) {real, imag} */,
  {32'h3f9b8a3e, 32'hbfb6c00c} /* (25, 7, 9) {real, imag} */,
  {32'hbe4aee3a, 32'hbe3af180} /* (25, 7, 8) {real, imag} */,
  {32'h3ffe4621, 32'hc006ae57} /* (25, 7, 7) {real, imag} */,
  {32'hbf24d720, 32'h3e250b94} /* (25, 7, 6) {real, imag} */,
  {32'h3ef01e34, 32'h3fe8d295} /* (25, 7, 5) {real, imag} */,
  {32'h3f30ccdc, 32'h3eb60f5b} /* (25, 7, 4) {real, imag} */,
  {32'h3d904410, 32'h400ce86b} /* (25, 7, 3) {real, imag} */,
  {32'h3fbd03fe, 32'h3f5f5880} /* (25, 7, 2) {real, imag} */,
  {32'h4035e1e6, 32'hbf963df0} /* (25, 7, 1) {real, imag} */,
  {32'h3f516d8c, 32'hbf6191fc} /* (25, 7, 0) {real, imag} */,
  {32'hbe057844, 32'h3f8882fc} /* (25, 6, 31) {real, imag} */,
  {32'hbf71ed84, 32'h40196b2b} /* (25, 6, 30) {real, imag} */,
  {32'hbf3d8851, 32'h3ed4151c} /* (25, 6, 29) {real, imag} */,
  {32'h400a4a16, 32'hbf728c62} /* (25, 6, 28) {real, imag} */,
  {32'h402031de, 32'h3fa4caf4} /* (25, 6, 27) {real, imag} */,
  {32'h3c5ff040, 32'h3fd5a010} /* (25, 6, 26) {real, imag} */,
  {32'h3da27bb0, 32'h3d904ba0} /* (25, 6, 25) {real, imag} */,
  {32'hbeb4d0a0, 32'hbec6e5e5} /* (25, 6, 24) {real, imag} */,
  {32'h3f89a74c, 32'hbf121aa6} /* (25, 6, 23) {real, imag} */,
  {32'h3f5418bc, 32'hbfbba6a2} /* (25, 6, 22) {real, imag} */,
  {32'h3df46050, 32'h3de104b8} /* (25, 6, 21) {real, imag} */,
  {32'h3ea07079, 32'h401eca8e} /* (25, 6, 20) {real, imag} */,
  {32'hbf364e3b, 32'h3f916f95} /* (25, 6, 19) {real, imag} */,
  {32'h3f0bc0ea, 32'hbf8cb9a3} /* (25, 6, 18) {real, imag} */,
  {32'h4011d40c, 32'hbec97d29} /* (25, 6, 17) {real, imag} */,
  {32'h40045af8, 32'h3f4e08b4} /* (25, 6, 16) {real, imag} */,
  {32'hbe8223fe, 32'hbea234a7} /* (25, 6, 15) {real, imag} */,
  {32'hbe8b005b, 32'h3f566a6d} /* (25, 6, 14) {real, imag} */,
  {32'hc02a5c51, 32'h3fdfeaf0} /* (25, 6, 13) {real, imag} */,
  {32'hbf068f07, 32'h3ed32bb0} /* (25, 6, 12) {real, imag} */,
  {32'h3fef8c1b, 32'h3f3441c8} /* (25, 6, 11) {real, imag} */,
  {32'h3fbbb156, 32'h3f55f3d3} /* (25, 6, 10) {real, imag} */,
  {32'h3f5fceb5, 32'hbf00345e} /* (25, 6, 9) {real, imag} */,
  {32'hc02ee8a2, 32'hbfc4c265} /* (25, 6, 8) {real, imag} */,
  {32'hbf648dce, 32'hc00e447e} /* (25, 6, 7) {real, imag} */,
  {32'hbe1d85f0, 32'h3f7f3ad3} /* (25, 6, 6) {real, imag} */,
  {32'h3faa76fd, 32'h4014e267} /* (25, 6, 5) {real, imag} */,
  {32'h3fe4ac41, 32'h404bec94} /* (25, 6, 4) {real, imag} */,
  {32'h3fb0354f, 32'h4008fc75} /* (25, 6, 3) {real, imag} */,
  {32'hbe6c8290, 32'h3f399906} /* (25, 6, 2) {real, imag} */,
  {32'h3f347812, 32'h3c4eb700} /* (25, 6, 1) {real, imag} */,
  {32'h3b14bb80, 32'h3ed861e8} /* (25, 6, 0) {real, imag} */,
  {32'h3ee7e750, 32'hbef01a2e} /* (25, 5, 31) {real, imag} */,
  {32'h3f1d4b9a, 32'h3f58c622} /* (25, 5, 30) {real, imag} */,
  {32'hbfcfa360, 32'hbf429e50} /* (25, 5, 29) {real, imag} */,
  {32'hbf94e611, 32'hbf3dfa67} /* (25, 5, 28) {real, imag} */,
  {32'h3f31eb80, 32'h3ffd91c7} /* (25, 5, 27) {real, imag} */,
  {32'h3fa6cd10, 32'h3fb8576f} /* (25, 5, 26) {real, imag} */,
  {32'h3e7edc70, 32'h40067f35} /* (25, 5, 25) {real, imag} */,
  {32'hbf8465a4, 32'h3ff98907} /* (25, 5, 24) {real, imag} */,
  {32'hc004d290, 32'h3e5fc024} /* (25, 5, 23) {real, imag} */,
  {32'hbebd6270, 32'hbf08ba56} /* (25, 5, 22) {real, imag} */,
  {32'h3fe25224, 32'h3ee9cf88} /* (25, 5, 21) {real, imag} */,
  {32'h3f494f61, 32'h4016868a} /* (25, 5, 20) {real, imag} */,
  {32'hc0490780, 32'h3f7f80be} /* (25, 5, 19) {real, imag} */,
  {32'hc0270934, 32'hbfd580fe} /* (25, 5, 18) {real, imag} */,
  {32'hbecff6a2, 32'hc004dd40} /* (25, 5, 17) {real, imag} */,
  {32'hbe3ebf3e, 32'h3f972e88} /* (25, 5, 16) {real, imag} */,
  {32'hbeb8ab4a, 32'h3f1fad74} /* (25, 5, 15) {real, imag} */,
  {32'hbe124b14, 32'hbd985ea8} /* (25, 5, 14) {real, imag} */,
  {32'hc013d509, 32'h3ee21b90} /* (25, 5, 13) {real, imag} */,
  {32'hbf40ed50, 32'h3df91b18} /* (25, 5, 12) {real, imag} */,
  {32'h3f097bf1, 32'hbff6eb0b} /* (25, 5, 11) {real, imag} */,
  {32'h3d918490, 32'hbf92c842} /* (25, 5, 10) {real, imag} */,
  {32'hbf8d64c6, 32'h3ca84300} /* (25, 5, 9) {real, imag} */,
  {32'hc04ff316, 32'hbfbd3c02} /* (25, 5, 8) {real, imag} */,
  {32'hbffe6458, 32'hc025fb16} /* (25, 5, 7) {real, imag} */,
  {32'h3fa9868b, 32'h3f507be5} /* (25, 5, 6) {real, imag} */,
  {32'h4027e931, 32'h3f89c314} /* (25, 5, 5) {real, imag} */,
  {32'h3ef7df34, 32'h403b87a6} /* (25, 5, 4) {real, imag} */,
  {32'h3fdc4aac, 32'h3fc9d738} /* (25, 5, 3) {real, imag} */,
  {32'h3e3c6488, 32'h3f3a2fe8} /* (25, 5, 2) {real, imag} */,
  {32'hbf525f28, 32'hbfc55e0e} /* (25, 5, 1) {real, imag} */,
  {32'h3f335052, 32'hbf44b006} /* (25, 5, 0) {real, imag} */,
  {32'h3f036484, 32'hbfaae32c} /* (25, 4, 31) {real, imag} */,
  {32'h3e843d50, 32'hbf24abc2} /* (25, 4, 30) {real, imag} */,
  {32'hbc4c66c0, 32'h3f9af1f6} /* (25, 4, 29) {real, imag} */,
  {32'hbf26a128, 32'h3fc6ff81} /* (25, 4, 28) {real, imag} */,
  {32'h3fee5f78, 32'h3e912116} /* (25, 4, 27) {real, imag} */,
  {32'h3f7c6d9a, 32'hbebe6300} /* (25, 4, 26) {real, imag} */,
  {32'hbf83e2e6, 32'h3ec64d50} /* (25, 4, 25) {real, imag} */,
  {32'hbdb04938, 32'h3eda57a9} /* (25, 4, 24) {real, imag} */,
  {32'hbfc235ea, 32'h3d8d7100} /* (25, 4, 23) {real, imag} */,
  {32'hbfabfb46, 32'hbfcd28dc} /* (25, 4, 22) {real, imag} */,
  {32'hbf6c5239, 32'hbfc6a57e} /* (25, 4, 21) {real, imag} */,
  {32'h3ed30140, 32'h3ec5fcf8} /* (25, 4, 20) {real, imag} */,
  {32'hc031fba9, 32'h3e275406} /* (25, 4, 19) {real, imag} */,
  {32'hc044e03c, 32'hbee7f6e8} /* (25, 4, 18) {real, imag} */,
  {32'hbf7683ce, 32'hbe29df70} /* (25, 4, 17) {real, imag} */,
  {32'h3f4049c2, 32'hbf9bee90} /* (25, 4, 16) {real, imag} */,
  {32'h3f84b6cf, 32'hc033f9d6} /* (25, 4, 15) {real, imag} */,
  {32'h3ea2087c, 32'hc00f49af} /* (25, 4, 14) {real, imag} */,
  {32'hbfdae6c0, 32'hc002a88a} /* (25, 4, 13) {real, imag} */,
  {32'hbf8b4e30, 32'h3de48422} /* (25, 4, 12) {real, imag} */,
  {32'hbee9186e, 32'hbfd36037} /* (25, 4, 11) {real, imag} */,
  {32'hbedb104a, 32'h3ed1e7c4} /* (25, 4, 10) {real, imag} */,
  {32'hbf2a8b7e, 32'h3f83e0ce} /* (25, 4, 9) {real, imag} */,
  {32'hc0133e2d, 32'hc020a836} /* (25, 4, 8) {real, imag} */,
  {32'hc0082ed2, 32'hc00ee874} /* (25, 4, 7) {real, imag} */,
  {32'hbf9a96d2, 32'hbeafb481} /* (25, 4, 6) {real, imag} */,
  {32'hbe2aa7f0, 32'hbfe0a974} /* (25, 4, 5) {real, imag} */,
  {32'hbf8c2b29, 32'h3f9ae7bc} /* (25, 4, 4) {real, imag} */,
  {32'hbf16e942, 32'h3f52471f} /* (25, 4, 3) {real, imag} */,
  {32'h3f6eefeb, 32'hbea789b8} /* (25, 4, 2) {real, imag} */,
  {32'hbef3b1e2, 32'hbf0b7532} /* (25, 4, 1) {real, imag} */,
  {32'h3f9da22e, 32'h3dab31d8} /* (25, 4, 0) {real, imag} */,
  {32'h3ea6b3d8, 32'hbecf45a7} /* (25, 3, 31) {real, imag} */,
  {32'h3f5e45ff, 32'h3ee74000} /* (25, 3, 30) {real, imag} */,
  {32'h3f906779, 32'h3fea1179} /* (25, 3, 29) {real, imag} */,
  {32'h3ffe079f, 32'h401e3428} /* (25, 3, 28) {real, imag} */,
  {32'h40867072, 32'h3f4d42fe} /* (25, 3, 27) {real, imag} */,
  {32'h3fa8916a, 32'hbf8c24b6} /* (25, 3, 26) {real, imag} */,
  {32'hbdba8fb0, 32'hbf5913b5} /* (25, 3, 25) {real, imag} */,
  {32'h3f99f02a, 32'hc014f98f} /* (25, 3, 24) {real, imag} */,
  {32'hbf67eada, 32'hbfaa03fa} /* (25, 3, 23) {real, imag} */,
  {32'hbfebcade, 32'hbfa31f1c} /* (25, 3, 22) {real, imag} */,
  {32'h3f24186c, 32'hbf8f205a} /* (25, 3, 21) {real, imag} */,
  {32'h4024fec6, 32'hbf616a14} /* (25, 3, 20) {real, imag} */,
  {32'hbddc5998, 32'hc003e618} /* (25, 3, 19) {real, imag} */,
  {32'hc004f228, 32'h3fbc9ddf} /* (25, 3, 18) {real, imag} */,
  {32'h3ece5088, 32'h4001b6e8} /* (25, 3, 17) {real, imag} */,
  {32'h3fa6f2e6, 32'hbea7a875} /* (25, 3, 16) {real, imag} */,
  {32'h3f39846e, 32'hc0783dee} /* (25, 3, 15) {real, imag} */,
  {32'h3faf4291, 32'hc088a319} /* (25, 3, 14) {real, imag} */,
  {32'hbf4bd963, 32'hbf09d3ba} /* (25, 3, 13) {real, imag} */,
  {32'hbf237f4c, 32'h3fce2cec} /* (25, 3, 12) {real, imag} */,
  {32'hc000889a, 32'hbf165add} /* (25, 3, 11) {real, imag} */,
  {32'hbf38c3d5, 32'h3f17ef3e} /* (25, 3, 10) {real, imag} */,
  {32'hbf958a5d, 32'h3fb35d14} /* (25, 3, 9) {real, imag} */,
  {32'hbfadacba, 32'hbf86f743} /* (25, 3, 8) {real, imag} */,
  {32'hbf874efc, 32'h3eb0c2ec} /* (25, 3, 7) {real, imag} */,
  {32'h3e51e4e0, 32'hbf11fd61} /* (25, 3, 6) {real, imag} */,
  {32'h3f64dea1, 32'hc046ee91} /* (25, 3, 5) {real, imag} */,
  {32'hbf44cfec, 32'h3e267f10} /* (25, 3, 4) {real, imag} */,
  {32'hbf8f0385, 32'h3fba6d5d} /* (25, 3, 3) {real, imag} */,
  {32'hbf8c1708, 32'hbea85cec} /* (25, 3, 2) {real, imag} */,
  {32'h3fd395c5, 32'hbefa3420} /* (25, 3, 1) {real, imag} */,
  {32'h3fc35abd, 32'h3ed0eba0} /* (25, 3, 0) {real, imag} */,
  {32'hbf4e6a75, 32'h3e4702ee} /* (25, 2, 31) {real, imag} */,
  {32'h3e97e542, 32'h3f684344} /* (25, 2, 30) {real, imag} */,
  {32'h3e081caa, 32'h3f8101ca} /* (25, 2, 29) {real, imag} */,
  {32'h3f134ed9, 32'h3ef3d4d6} /* (25, 2, 28) {real, imag} */,
  {32'h3fe451b3, 32'hbf4d1504} /* (25, 2, 27) {real, imag} */,
  {32'h3dafeeb0, 32'hbfe8a074} /* (25, 2, 26) {real, imag} */,
  {32'h3f0eeefc, 32'hbfc55d90} /* (25, 2, 25) {real, imag} */,
  {32'h4019c1e8, 32'hc0423fa3} /* (25, 2, 24) {real, imag} */,
  {32'hbf9205bc, 32'hbfd2696e} /* (25, 2, 23) {real, imag} */,
  {32'hbfa8ca9e, 32'h3e8df8dc} /* (25, 2, 22) {real, imag} */,
  {32'h3fc037f5, 32'h3f844cfe} /* (25, 2, 21) {real, imag} */,
  {32'h3fbf1d47, 32'h3d97f7d4} /* (25, 2, 20) {real, imag} */,
  {32'h3ea83b3b, 32'hbfc8ebb8} /* (25, 2, 19) {real, imag} */,
  {32'hbfce007e, 32'h3f7d155e} /* (25, 2, 18) {real, imag} */,
  {32'hbeafd307, 32'h3f8dd544} /* (25, 2, 17) {real, imag} */,
  {32'hbf6e7ebe, 32'hbf1d5ce0} /* (25, 2, 16) {real, imag} */,
  {32'hc020584a, 32'hc037a6d0} /* (25, 2, 15) {real, imag} */,
  {32'hbf86f7e2, 32'hc05bbe0f} /* (25, 2, 14) {real, imag} */,
  {32'hbf48b442, 32'h3f74a392} /* (25, 2, 13) {real, imag} */,
  {32'hbed6c818, 32'h4015c5d5} /* (25, 2, 12) {real, imag} */,
  {32'hbec529c8, 32'h3ea46598} /* (25, 2, 11) {real, imag} */,
  {32'hc0145114, 32'h3dd12768} /* (25, 2, 10) {real, imag} */,
  {32'hc0659e2e, 32'h3fe4e40e} /* (25, 2, 9) {real, imag} */,
  {32'hbd2db750, 32'h3f31ed38} /* (25, 2, 8) {real, imag} */,
  {32'h3edc3ae0, 32'h3f804e1b} /* (25, 2, 7) {real, imag} */,
  {32'h3f919348, 32'h3fbbf67e} /* (25, 2, 6) {real, imag} */,
  {32'h3f8a8eba, 32'hc001366c} /* (25, 2, 5) {real, imag} */,
  {32'hbf046330, 32'hc034baab} /* (25, 2, 4) {real, imag} */,
  {32'h3d5d2da0, 32'hbfd7cf47} /* (25, 2, 3) {real, imag} */,
  {32'h3e8a51fe, 32'hbf76add2} /* (25, 2, 2) {real, imag} */,
  {32'h3f149fd7, 32'hbfd52142} /* (25, 2, 1) {real, imag} */,
  {32'hbefb606c, 32'hbf7646d3} /* (25, 2, 0) {real, imag} */,
  {32'hbee3eacf, 32'hbf219ae4} /* (25, 1, 31) {real, imag} */,
  {32'h3ee77ea4, 32'h3d91440c} /* (25, 1, 30) {real, imag} */,
  {32'h3ebae542, 32'h3ffc3201} /* (25, 1, 29) {real, imag} */,
  {32'h3fdf95a4, 32'h3fa308b8} /* (25, 1, 28) {real, imag} */,
  {32'h3f1cf6d8, 32'hbf0a349d} /* (25, 1, 27) {real, imag} */,
  {32'hbf6d26dc, 32'hbf872f64} /* (25, 1, 26) {real, imag} */,
  {32'hbe60c8d8, 32'hbf2ae6fe} /* (25, 1, 25) {real, imag} */,
  {32'h3fe1cc28, 32'hbfa26b7c} /* (25, 1, 24) {real, imag} */,
  {32'hbc9601a0, 32'h3e2405b0} /* (25, 1, 23) {real, imag} */,
  {32'h3f8567fb, 32'h400fda00} /* (25, 1, 22) {real, imag} */,
  {32'h3f8a39d2, 32'h4016e08e} /* (25, 1, 21) {real, imag} */,
  {32'hbe86f49e, 32'h3f7d2ebe} /* (25, 1, 20) {real, imag} */,
  {32'h3f1c1efd, 32'hbf16a2fd} /* (25, 1, 19) {real, imag} */,
  {32'hbfe67871, 32'h3e9652c8} /* (25, 1, 18) {real, imag} */,
  {32'hbfd239ca, 32'h3ea07b2c} /* (25, 1, 17) {real, imag} */,
  {32'h3e318fc8, 32'h3eecf2eb} /* (25, 1, 16) {real, imag} */,
  {32'hbe85b3ae, 32'h3e91038a} /* (25, 1, 15) {real, imag} */,
  {32'hbe8dc553, 32'hbf5ff5f4} /* (25, 1, 14) {real, imag} */,
  {32'hbfee67f9, 32'hc015832d} /* (25, 1, 13) {real, imag} */,
  {32'hbfe979eb, 32'hbf2a629c} /* (25, 1, 12) {real, imag} */,
  {32'h3e53c854, 32'h3f1301a8} /* (25, 1, 11) {real, imag} */,
  {32'hc01dce47, 32'h3e873b8a} /* (25, 1, 10) {real, imag} */,
  {32'hc0284bac, 32'h401277fc} /* (25, 1, 9) {real, imag} */,
  {32'h3f727250, 32'h3feebd90} /* (25, 1, 8) {real, imag} */,
  {32'h3fbc31af, 32'h3f63d29a} /* (25, 1, 7) {real, imag} */,
  {32'h3eac26d0, 32'h3f8c49a8} /* (25, 1, 6) {real, imag} */,
  {32'h3f0b2831, 32'hbfb4671b} /* (25, 1, 5) {real, imag} */,
  {32'hbe3e9988, 32'hc05a8bce} /* (25, 1, 4) {real, imag} */,
  {32'hbfd4ea4e, 32'hc021149c} /* (25, 1, 3) {real, imag} */,
  {32'h3f05931a, 32'hbea3ff92} /* (25, 1, 2) {real, imag} */,
  {32'h3f2f0e72, 32'hbf8baef6} /* (25, 1, 1) {real, imag} */,
  {32'h3e788d04, 32'hc0049185} /* (25, 1, 0) {real, imag} */,
  {32'hbf76eca2, 32'hbf1a9764} /* (25, 0, 31) {real, imag} */,
  {32'hbeff48d0, 32'hbd557c08} /* (25, 0, 30) {real, imag} */,
  {32'hbf702360, 32'h3fd2d172} /* (25, 0, 29) {real, imag} */,
  {32'h3f3ef1e6, 32'h3f973008} /* (25, 0, 28) {real, imag} */,
  {32'h3e1f62ec, 32'h3f1f0c04} /* (25, 0, 27) {real, imag} */,
  {32'hbf9adecb, 32'hbebd8352} /* (25, 0, 26) {real, imag} */,
  {32'hbe8c0b94, 32'hbc952180} /* (25, 0, 25) {real, imag} */,
  {32'h3fab9e82, 32'hbe962dbe} /* (25, 0, 24) {real, imag} */,
  {32'h3f20ad12, 32'hbc776c20} /* (25, 0, 23) {real, imag} */,
  {32'h3f957e54, 32'h3f2163be} /* (25, 0, 22) {real, imag} */,
  {32'h3e97d5d0, 32'h3f7e2464} /* (25, 0, 21) {real, imag} */,
  {32'hbef1a132, 32'h3f4092e1} /* (25, 0, 20) {real, imag} */,
  {32'hbde8b260, 32'hbf915024} /* (25, 0, 19) {real, imag} */,
  {32'hbd9d435a, 32'hbf1ad1a9} /* (25, 0, 18) {real, imag} */,
  {32'hbf25d009, 32'h3e0d4878} /* (25, 0, 17) {real, imag} */,
  {32'h3e2ffbb0, 32'h3f9a9129} /* (25, 0, 16) {real, imag} */,
  {32'h3f30431c, 32'h3f454ee2} /* (25, 0, 15) {real, imag} */,
  {32'h3fdcfe79, 32'h3e904fe0} /* (25, 0, 14) {real, imag} */,
  {32'hbf3862c8, 32'hc027f8e0} /* (25, 0, 13) {real, imag} */,
  {32'hbfb1eaa0, 32'hbff4ce91} /* (25, 0, 12) {real, imag} */,
  {32'hbf903dac, 32'hbf195238} /* (25, 0, 11) {real, imag} */,
  {32'hbfcea005, 32'h3faf75b2} /* (25, 0, 10) {real, imag} */,
  {32'hbf6101e6, 32'h3f4f9054} /* (25, 0, 9) {real, imag} */,
  {32'h3f330295, 32'h3f424038} /* (25, 0, 8) {real, imag} */,
  {32'h3f05c102, 32'h3e8c1926} /* (25, 0, 7) {real, imag} */,
  {32'hbfa660ef, 32'hbec5ac5b} /* (25, 0, 6) {real, imag} */,
  {32'hbe54d64e, 32'hbf7159b1} /* (25, 0, 5) {real, imag} */,
  {32'h3eeb5784, 32'hbf853738} /* (25, 0, 4) {real, imag} */,
  {32'hbf906bfa, 32'hbe5922e9} /* (25, 0, 3) {real, imag} */,
  {32'hbea86ada, 32'h3f86a56c} /* (25, 0, 2) {real, imag} */,
  {32'h3ddbf910, 32'hbcaa3080} /* (25, 0, 1) {real, imag} */,
  {32'hbddc8db4, 32'hbfb21a1a} /* (25, 0, 0) {real, imag} */,
  {32'hbf53abfe, 32'hbe2fa19c} /* (24, 31, 31) {real, imag} */,
  {32'hbfae7ae0, 32'h3ee1e9ea} /* (24, 31, 30) {real, imag} */,
  {32'hbffe45e2, 32'h3f0cd25a} /* (24, 31, 29) {real, imag} */,
  {32'hc0084a97, 32'hbfadacab} /* (24, 31, 28) {real, imag} */,
  {32'hbfab89b6, 32'hbf0d89cb} /* (24, 31, 27) {real, imag} */,
  {32'hbdd74d38, 32'h3f464f0e} /* (24, 31, 26) {real, imag} */,
  {32'hc00b75ce, 32'hbfb12704} /* (24, 31, 25) {real, imag} */,
  {32'hc03f9031, 32'hbf2f5886} /* (24, 31, 24) {real, imag} */,
  {32'hbffb9831, 32'hbfceff88} /* (24, 31, 23) {real, imag} */,
  {32'hbfb1e41f, 32'hbfc9a143} /* (24, 31, 22) {real, imag} */,
  {32'hbe5c6731, 32'hbf4af048} /* (24, 31, 21) {real, imag} */,
  {32'h3f5a23e2, 32'h3f66a744} /* (24, 31, 20) {real, imag} */,
  {32'h3f8aac40, 32'h3f9bce02} /* (24, 31, 19) {real, imag} */,
  {32'h3f0ea902, 32'h3edc20a6} /* (24, 31, 18) {real, imag} */,
  {32'h3e10cf8a, 32'h3ee40574} /* (24, 31, 17) {real, imag} */,
  {32'h3f1fbc13, 32'h3f42c2b8} /* (24, 31, 16) {real, imag} */,
  {32'hbf0546d8, 32'h3fe3b630} /* (24, 31, 15) {real, imag} */,
  {32'h3f85fe5d, 32'h3fa569a6} /* (24, 31, 14) {real, imag} */,
  {32'h3ff3eeac, 32'h3fdd24b6} /* (24, 31, 13) {real, imag} */,
  {32'h3f7e5ec8, 32'h40002a66} /* (24, 31, 12) {real, imag} */,
  {32'h3f9de393, 32'h4018d738} /* (24, 31, 11) {real, imag} */,
  {32'h3f413b9d, 32'h3f50afbb} /* (24, 31, 10) {real, imag} */,
  {32'h3fc64d3a, 32'hbe4756ea} /* (24, 31, 9) {real, imag} */,
  {32'h3e4eb1a0, 32'hbeccc150} /* (24, 31, 8) {real, imag} */,
  {32'h3ee88ff0, 32'hc0016d47} /* (24, 31, 7) {real, imag} */,
  {32'hbf5c7e77, 32'hbfe44b48} /* (24, 31, 6) {real, imag} */,
  {32'hc002f4c6, 32'hbffb7e3d} /* (24, 31, 5) {real, imag} */,
  {32'hbf0b0010, 32'hbfea50e6} /* (24, 31, 4) {real, imag} */,
  {32'hbefc5662, 32'hbfd047e3} /* (24, 31, 3) {real, imag} */,
  {32'h3f3c028d, 32'hc04cc009} /* (24, 31, 2) {real, imag} */,
  {32'hbf3f0720, 32'hbff86a3e} /* (24, 31, 1) {real, imag} */,
  {32'hc0170cf9, 32'hbe496c0e} /* (24, 31, 0) {real, imag} */,
  {32'hbfda2124, 32'hbee5b8ef} /* (24, 30, 31) {real, imag} */,
  {32'hc0457104, 32'h3f874822} /* (24, 30, 30) {real, imag} */,
  {32'hc055c0a4, 32'h3f093e8e} /* (24, 30, 29) {real, imag} */,
  {32'hc0295e30, 32'hc02569f2} /* (24, 30, 28) {real, imag} */,
  {32'hc00e09d4, 32'h3ee4b1c8} /* (24, 30, 27) {real, imag} */,
  {32'hbfc2f25e, 32'h3fe5259a} /* (24, 30, 26) {real, imag} */,
  {32'hc01a8e77, 32'hbf990209} /* (24, 30, 25) {real, imag} */,
  {32'hc05cbc4f, 32'hbf0cbae0} /* (24, 30, 24) {real, imag} */,
  {32'hc03b4795, 32'hc0029d99} /* (24, 30, 23) {real, imag} */,
  {32'hbf29049f, 32'hc034a9c0} /* (24, 30, 22) {real, imag} */,
  {32'h3ee1090e, 32'hbdb35398} /* (24, 30, 21) {real, imag} */,
  {32'h3f051d2a, 32'h402039d6} /* (24, 30, 20) {real, imag} */,
  {32'h3f0155af, 32'h4042c433} /* (24, 30, 19) {real, imag} */,
  {32'h4008c014, 32'h3fdfebbe} /* (24, 30, 18) {real, imag} */,
  {32'h400c68e6, 32'h3fd58abf} /* (24, 30, 17) {real, imag} */,
  {32'h3fca4bcc, 32'h403160ff} /* (24, 30, 16) {real, imag} */,
  {32'h3fd41a5a, 32'h40574ca6} /* (24, 30, 15) {real, imag} */,
  {32'h405fe2a6, 32'h404ee3f4} /* (24, 30, 14) {real, imag} */,
  {32'h4038c278, 32'h4043d46e} /* (24, 30, 13) {real, imag} */,
  {32'h400fcf1f, 32'h4024dfd0} /* (24, 30, 12) {real, imag} */,
  {32'h4027ca66, 32'h3f87016a} /* (24, 30, 11) {real, imag} */,
  {32'h3f8aaa63, 32'hbf2bdcba} /* (24, 30, 10) {real, imag} */,
  {32'h3f83f54e, 32'h3d558750} /* (24, 30, 9) {real, imag} */,
  {32'hbf5c3150, 32'hbf2de8de} /* (24, 30, 8) {real, imag} */,
  {32'hbfb70d25, 32'hc0010fe1} /* (24, 30, 7) {real, imag} */,
  {32'hc009babe, 32'hc05327a0} /* (24, 30, 6) {real, imag} */,
  {32'hc01b64a0, 32'hc0a70a93} /* (24, 30, 5) {real, imag} */,
  {32'hbfa5fcb5, 32'hc04b3d8a} /* (24, 30, 4) {real, imag} */,
  {32'hbfd8e2ec, 32'hbf96427e} /* (24, 30, 3) {real, imag} */,
  {32'hbe65cc48, 32'hc05fed59} /* (24, 30, 2) {real, imag} */,
  {32'hbfe783a6, 32'hc0159413} /* (24, 30, 1) {real, imag} */,
  {32'hc0444253, 32'hbf7fa3c4} /* (24, 30, 0) {real, imag} */,
  {32'hc01aee8d, 32'h3f0c5460} /* (24, 29, 31) {real, imag} */,
  {32'hc04259fa, 32'hbf500c03} /* (24, 29, 30) {real, imag} */,
  {32'hc023c67e, 32'hc03529b3} /* (24, 29, 29) {real, imag} */,
  {32'hbfdb9e09, 32'hc047aea2} /* (24, 29, 28) {real, imag} */,
  {32'hbfe3461f, 32'hbfae807c} /* (24, 29, 27) {real, imag} */,
  {32'hbf88ec2d, 32'hbf4d389e} /* (24, 29, 26) {real, imag} */,
  {32'hbe0e3758, 32'hbf967eba} /* (24, 29, 25) {real, imag} */,
  {32'hbffe1922, 32'hbe8f03e2} /* (24, 29, 24) {real, imag} */,
  {32'hc004da7b, 32'hbfae5942} /* (24, 29, 23) {real, imag} */,
  {32'h3f2a3fcd, 32'hc04031b9} /* (24, 29, 22) {real, imag} */,
  {32'h3fdb2c03, 32'hbf79b57e} /* (24, 29, 21) {real, imag} */,
  {32'h3ebb33aa, 32'h3ffc6a27} /* (24, 29, 20) {real, imag} */,
  {32'hc00ff469, 32'h3ff53587} /* (24, 29, 19) {real, imag} */,
  {32'h3e8b354a, 32'h3feb489a} /* (24, 29, 18) {real, imag} */,
  {32'h400e2188, 32'h3f8fff74} /* (24, 29, 17) {real, imag} */,
  {32'h3fc19f20, 32'h3fe05037} /* (24, 29, 16) {real, imag} */,
  {32'h400d96c0, 32'h3fd50394} /* (24, 29, 15) {real, imag} */,
  {32'h40233310, 32'h3febb05a} /* (24, 29, 14) {real, imag} */,
  {32'h3fe27c3b, 32'h3fe5c8ef} /* (24, 29, 13) {real, imag} */,
  {32'h40226380, 32'h3fcc1970} /* (24, 29, 12) {real, imag} */,
  {32'h406e6899, 32'h3ed0ecb4} /* (24, 29, 11) {real, imag} */,
  {32'h3eb65080, 32'hbfff9863} /* (24, 29, 10) {real, imag} */,
  {32'hc030d09b, 32'hc024ec95} /* (24, 29, 9) {real, imag} */,
  {32'hc03c675f, 32'hc00f7c85} /* (24, 29, 8) {real, imag} */,
  {32'hc002823a, 32'hbfd0fec4} /* (24, 29, 7) {real, imag} */,
  {32'hbfea15b6, 32'hc040dfc5} /* (24, 29, 6) {real, imag} */,
  {32'hc0033ee9, 32'hc09d45cc} /* (24, 29, 5) {real, imag} */,
  {32'hbf144b7e, 32'hc08bf74e} /* (24, 29, 4) {real, imag} */,
  {32'hbee7d2b8, 32'hc02a474c} /* (24, 29, 3) {real, imag} */,
  {32'h3ec522ac, 32'hc051ab44} /* (24, 29, 2) {real, imag} */,
  {32'hbfff86c6, 32'hbfb3dd57} /* (24, 29, 1) {real, imag} */,
  {32'hc053dcf2, 32'hbfa61bf2} /* (24, 29, 0) {real, imag} */,
  {32'hc0118782, 32'hbe780d4a} /* (24, 28, 31) {real, imag} */,
  {32'hc0169cb8, 32'hc03a2dfc} /* (24, 28, 30) {real, imag} */,
  {32'hbfd02f8e, 32'hc0597ad3} /* (24, 28, 29) {real, imag} */,
  {32'hbf753ed4, 32'hc00f406d} /* (24, 28, 28) {real, imag} */,
  {32'hbfd568bb, 32'hc00028a5} /* (24, 28, 27) {real, imag} */,
  {32'hbf3c9fb2, 32'hc05eea43} /* (24, 28, 26) {real, imag} */,
  {32'h3f2df2b0, 32'hbff5a3ba} /* (24, 28, 25) {real, imag} */,
  {32'hc00e0838, 32'h3d79f780} /* (24, 28, 24) {real, imag} */,
  {32'hbfd660b3, 32'hc044d5d2} /* (24, 28, 23) {real, imag} */,
  {32'h3ef1a1b5, 32'hc03ebdc2} /* (24, 28, 22) {real, imag} */,
  {32'h3faf77da, 32'hc00ac3b6} /* (24, 28, 21) {real, imag} */,
  {32'h3f314c66, 32'h3fb559a6} /* (24, 28, 20) {real, imag} */,
  {32'hbfc0f097, 32'h40102176} /* (24, 28, 19) {real, imag} */,
  {32'hbcadd760, 32'h402aa3c6} /* (24, 28, 18) {real, imag} */,
  {32'h3e836358, 32'h3fbca286} /* (24, 28, 17) {real, imag} */,
  {32'h3f672d06, 32'h3ef57e54} /* (24, 28, 16) {real, imag} */,
  {32'h401a783a, 32'hbd452bc8} /* (24, 28, 15) {real, imag} */,
  {32'h3f8d3b07, 32'h3de322f4} /* (24, 28, 14) {real, imag} */,
  {32'h3fb19bce, 32'h3f19d3ac} /* (24, 28, 13) {real, imag} */,
  {32'h3f8970c7, 32'h3fed2a86} /* (24, 28, 12) {real, imag} */,
  {32'h4042fdd2, 32'h3fa390bc} /* (24, 28, 11) {real, imag} */,
  {32'h3e76a73c, 32'hbeac68c8} /* (24, 28, 10) {real, imag} */,
  {32'hc0285fd9, 32'hc02881dc} /* (24, 28, 9) {real, imag} */,
  {32'hc00fadf6, 32'hc0014144} /* (24, 28, 8) {real, imag} */,
  {32'hbf0a2556, 32'hbfd5a65e} /* (24, 28, 7) {real, imag} */,
  {32'hbfdac50d, 32'hc023c928} /* (24, 28, 6) {real, imag} */,
  {32'hbfa3fbd5, 32'hc05a56c0} /* (24, 28, 5) {real, imag} */,
  {32'hbe120c7c, 32'hc05225b6} /* (24, 28, 4) {real, imag} */,
  {32'hbfc26d00, 32'hc01236de} /* (24, 28, 3) {real, imag} */,
  {32'hbf22d3bb, 32'hc0265668} /* (24, 28, 2) {real, imag} */,
  {32'hc0484cde, 32'hc017d4f1} /* (24, 28, 1) {real, imag} */,
  {32'hc056af14, 32'hc0091770} /* (24, 28, 0) {real, imag} */,
  {32'hbfd1e2a0, 32'hbf96453e} /* (24, 27, 31) {real, imag} */,
  {32'hbfc82fdf, 32'hc0304ddc} /* (24, 27, 30) {real, imag} */,
  {32'hc00a8a52, 32'hc02e26ee} /* (24, 27, 29) {real, imag} */,
  {32'hbfb47c25, 32'hc0373c9d} /* (24, 27, 28) {real, imag} */,
  {32'hc014702c, 32'hbfed2ec0} /* (24, 27, 27) {real, imag} */,
  {32'hc0241d20, 32'hc022786f} /* (24, 27, 26) {real, imag} */,
  {32'hbf9f190a, 32'hbf1d78a0} /* (24, 27, 25) {real, imag} */,
  {32'hc08940ac, 32'hbfbb608b} /* (24, 27, 24) {real, imag} */,
  {32'hc081aa2a, 32'hc082889f} /* (24, 27, 23) {real, imag} */,
  {32'hc0349d5a, 32'hc06dddb4} /* (24, 27, 22) {real, imag} */,
  {32'hbf44569e, 32'hc063ec97} /* (24, 27, 21) {real, imag} */,
  {32'h3f88c502, 32'h3fc36b07} /* (24, 27, 20) {real, imag} */,
  {32'h3f0b2151, 32'h401ec115} /* (24, 27, 19) {real, imag} */,
  {32'h3ff62378, 32'h405d9556} /* (24, 27, 18) {real, imag} */,
  {32'h3f390b49, 32'h4068fb1a} /* (24, 27, 17) {real, imag} */,
  {32'hbeb0fc80, 32'h4048b79a} /* (24, 27, 16) {real, imag} */,
  {32'h3fea3b9b, 32'h3ff32fde} /* (24, 27, 15) {real, imag} */,
  {32'h3f557cde, 32'h3f3a8da8} /* (24, 27, 14) {real, imag} */,
  {32'h3fc81176, 32'h3bb73900} /* (24, 27, 13) {real, imag} */,
  {32'h3f9fd4ad, 32'h3f9c956c} /* (24, 27, 12) {real, imag} */,
  {32'h40512108, 32'h403e886a} /* (24, 27, 11) {real, imag} */,
  {32'h3ea4837a, 32'h3edf2fc6} /* (24, 27, 10) {real, imag} */,
  {32'hbdcc1b30, 32'hbf98570c} /* (24, 27, 9) {real, imag} */,
  {32'h3db36f70, 32'hbf8f39e8} /* (24, 27, 8) {real, imag} */,
  {32'h3d77cca0, 32'hbf627dd2} /* (24, 27, 7) {real, imag} */,
  {32'hbfdf5128, 32'hbfcab63a} /* (24, 27, 6) {real, imag} */,
  {32'h3d298740, 32'hc01fcea8} /* (24, 27, 5) {real, imag} */,
  {32'h3eeffaf6, 32'hc033df8c} /* (24, 27, 4) {real, imag} */,
  {32'hbfbe3726, 32'hbfe1efac} /* (24, 27, 3) {real, imag} */,
  {32'hbfa83402, 32'hc03a1d93} /* (24, 27, 2) {real, imag} */,
  {32'hbfafa9cc, 32'hc01cbc85} /* (24, 27, 1) {real, imag} */,
  {32'hbfcef8c6, 32'hc0070e32} /* (24, 27, 0) {real, imag} */,
  {32'hbe43ab4a, 32'hbf431e1d} /* (24, 26, 31) {real, imag} */,
  {32'hc00ddd0f, 32'hc027d2e4} /* (24, 26, 30) {real, imag} */,
  {32'hc06c6440, 32'hbfceda60} /* (24, 26, 29) {real, imag} */,
  {32'hbfdadbcc, 32'hbf2a9e10} /* (24, 26, 28) {real, imag} */,
  {32'hc00c1818, 32'hbfc87126} /* (24, 26, 27) {real, imag} */,
  {32'hc0126a6d, 32'hbf008b48} /* (24, 26, 26) {real, imag} */,
  {32'hc00a64b0, 32'hbeba0d4c} /* (24, 26, 25) {real, imag} */,
  {32'hc03e7cb4, 32'hbffc7afa} /* (24, 26, 24) {real, imag} */,
  {32'hbfe3145f, 32'hbfd4c85a} /* (24, 26, 23) {real, imag} */,
  {32'hbfa36dbd, 32'hc0154034} /* (24, 26, 22) {real, imag} */,
  {32'hbecde314, 32'hc05ae1f2} /* (24, 26, 21) {real, imag} */,
  {32'h3fdace00, 32'hbc038980} /* (24, 26, 20) {real, imag} */,
  {32'h400a460a, 32'h3fcd71a3} /* (24, 26, 19) {real, imag} */,
  {32'h402e4b99, 32'h40119d2c} /* (24, 26, 18) {real, imag} */,
  {32'h40160cd0, 32'h404b6220} /* (24, 26, 17) {real, imag} */,
  {32'h3efa613c, 32'h408a8f46} /* (24, 26, 16) {real, imag} */,
  {32'h40254bfa, 32'h40207975} /* (24, 26, 15) {real, imag} */,
  {32'h3ffdfce1, 32'h402544ff} /* (24, 26, 14) {real, imag} */,
  {32'h3fe5422a, 32'h3fb1f496} /* (24, 26, 13) {real, imag} */,
  {32'h400da916, 32'h3fe2b244} /* (24, 26, 12) {real, imag} */,
  {32'h3f8c3ab7, 32'h4036a9b6} /* (24, 26, 11) {real, imag} */,
  {32'hbf6f12a4, 32'hbff12cfe} /* (24, 26, 10) {real, imag} */,
  {32'hbea3b134, 32'hc03f74da} /* (24, 26, 9) {real, imag} */,
  {32'h3e8d91f8, 32'hbf8f36b8} /* (24, 26, 8) {real, imag} */,
  {32'hc021025c, 32'hbebbcfde} /* (24, 26, 7) {real, imag} */,
  {32'hc0510b33, 32'hbe5c9e0c} /* (24, 26, 6) {real, imag} */,
  {32'hc00ba79a, 32'hbee4bcb8} /* (24, 26, 5) {real, imag} */,
  {32'hbf125260, 32'hbf9fb6c8} /* (24, 26, 4) {real, imag} */,
  {32'hbfe51bd1, 32'hc02850b3} /* (24, 26, 3) {real, imag} */,
  {32'hc0066968, 32'hc0226d84} /* (24, 26, 2) {real, imag} */,
  {32'h3e8e5aa8, 32'hc00c0da6} /* (24, 26, 1) {real, imag} */,
  {32'hbe6b8fac, 32'hc00379a6} /* (24, 26, 0) {real, imag} */,
  {32'hbf26097c, 32'hbf327680} /* (24, 25, 31) {real, imag} */,
  {32'hc03c4246, 32'hbfceb2f9} /* (24, 25, 30) {real, imag} */,
  {32'hc09b2253, 32'hbf308c99} /* (24, 25, 29) {real, imag} */,
  {32'hc031a9f8, 32'h3e8609f8} /* (24, 25, 28) {real, imag} */,
  {32'hbfaed643, 32'hbfddae73} /* (24, 25, 27) {real, imag} */,
  {32'hbf9d01d0, 32'hbf575ec2} /* (24, 25, 26) {real, imag} */,
  {32'hc0062ff4, 32'h3d498ec0} /* (24, 25, 25) {real, imag} */,
  {32'hbf60ac63, 32'hbffc196f} /* (24, 25, 24) {real, imag} */,
  {32'hbefc9ae4, 32'hbf8cfdb4} /* (24, 25, 23) {real, imag} */,
  {32'hbf84651e, 32'hc0003681} /* (24, 25, 22) {real, imag} */,
  {32'hbf3b8c36, 32'h3ca17300} /* (24, 25, 21) {real, imag} */,
  {32'h3fa4c49a, 32'h40151dde} /* (24, 25, 20) {real, imag} */,
  {32'h3fe819f4, 32'h4003ff42} /* (24, 25, 19) {real, imag} */,
  {32'h403120ac, 32'h3fc3767c} /* (24, 25, 18) {real, imag} */,
  {32'h408ea604, 32'h4013803c} /* (24, 25, 17) {real, imag} */,
  {32'h402fd70c, 32'h406a8e2c} /* (24, 25, 16) {real, imag} */,
  {32'h4030d0ae, 32'h402e4a70} /* (24, 25, 15) {real, imag} */,
  {32'h405763ac, 32'h3fbfb3ec} /* (24, 25, 14) {real, imag} */,
  {32'h405f9232, 32'hbec24bc0} /* (24, 25, 13) {real, imag} */,
  {32'h401db3aa, 32'h40471986} /* (24, 25, 12) {real, imag} */,
  {32'hbe0d3d80, 32'h40189904} /* (24, 25, 11) {real, imag} */,
  {32'hc0000842, 32'hbfb6d9a8} /* (24, 25, 10) {real, imag} */,
  {32'hc03a5114, 32'hc026398c} /* (24, 25, 9) {real, imag} */,
  {32'hc02da418, 32'hc059662a} /* (24, 25, 8) {real, imag} */,
  {32'hc041a3de, 32'hbfdb8700} /* (24, 25, 7) {real, imag} */,
  {32'hc0471d92, 32'hbd5b9180} /* (24, 25, 6) {real, imag} */,
  {32'hc086ccaa, 32'hbdbdc010} /* (24, 25, 5) {real, imag} */,
  {32'hc057a03f, 32'hbf05847a} /* (24, 25, 4) {real, imag} */,
  {32'hc0634b2a, 32'hc01e8595} /* (24, 25, 3) {real, imag} */,
  {32'hc032af7f, 32'hc0124b2e} /* (24, 25, 2) {real, imag} */,
  {32'hbf769a58, 32'hbfde8c8a} /* (24, 25, 1) {real, imag} */,
  {32'hbebdd9e0, 32'hbfb77d4a} /* (24, 25, 0) {real, imag} */,
  {32'hbf9f1f34, 32'hbef0ce6c} /* (24, 24, 31) {real, imag} */,
  {32'hbfc89390, 32'hbfd60bed} /* (24, 24, 30) {real, imag} */,
  {32'hc0223903, 32'hc0274f7f} /* (24, 24, 29) {real, imag} */,
  {32'hbfb21cda, 32'hbfd41534} /* (24, 24, 28) {real, imag} */,
  {32'h3d0c1120, 32'hc0388058} /* (24, 24, 27) {real, imag} */,
  {32'h3ed3b276, 32'hc00f5587} /* (24, 24, 26) {real, imag} */,
  {32'h3eded40a, 32'h3f013758} /* (24, 24, 25) {real, imag} */,
  {32'hc0030696, 32'hbf96e3cf} /* (24, 24, 24) {real, imag} */,
  {32'hc01bae08, 32'hbfed7d65} /* (24, 24, 23) {real, imag} */,
  {32'hbf8f21b5, 32'hc04bc561} /* (24, 24, 22) {real, imag} */,
  {32'hbf43ea80, 32'h3ed10628} /* (24, 24, 21) {real, imag} */,
  {32'h3ffc1a77, 32'h4085511a} /* (24, 24, 20) {real, imag} */,
  {32'h3f1f73ba, 32'h404b14c7} /* (24, 24, 19) {real, imag} */,
  {32'h3f8c92b3, 32'h3fea8485} /* (24, 24, 18) {real, imag} */,
  {32'h405ec67e, 32'h4001a1c0} /* (24, 24, 17) {real, imag} */,
  {32'h4050bb58, 32'h3fbe5441} /* (24, 24, 16) {real, imag} */,
  {32'h3f351053, 32'h3fcc623d} /* (24, 24, 15) {real, imag} */,
  {32'h4010ab94, 32'hbed9bfcc} /* (24, 24, 14) {real, imag} */,
  {32'h4026a5fc, 32'h3f166118} /* (24, 24, 13) {real, imag} */,
  {32'h406bb1a2, 32'h3f579ace} /* (24, 24, 12) {real, imag} */,
  {32'h40186232, 32'h3f28bbb8} /* (24, 24, 11) {real, imag} */,
  {32'hbf434244, 32'hbf7be8dc} /* (24, 24, 10) {real, imag} */,
  {32'hc04a2d9e, 32'hc0474ed7} /* (24, 24, 9) {real, imag} */,
  {32'hc0898078, 32'hbfdb37f7} /* (24, 24, 8) {real, imag} */,
  {32'hbf8bc0b8, 32'hbf2764fc} /* (24, 24, 7) {real, imag} */,
  {32'hbf9ece8c, 32'hbfb84ff6} /* (24, 24, 6) {real, imag} */,
  {32'hc005d076, 32'hbf827514} /* (24, 24, 5) {real, imag} */,
  {32'hbf83bfa6, 32'hbf288ae5} /* (24, 24, 4) {real, imag} */,
  {32'hc06cb4ca, 32'hbfe10704} /* (24, 24, 3) {real, imag} */,
  {32'hc091de66, 32'hc0229112} /* (24, 24, 2) {real, imag} */,
  {32'hc013bb9e, 32'hc004186c} /* (24, 24, 1) {real, imag} */,
  {32'hbfdaec92, 32'hbf33309b} /* (24, 24, 0) {real, imag} */,
  {32'hbfa603c7, 32'hbd75a500} /* (24, 23, 31) {real, imag} */,
  {32'hbd2a1f20, 32'hc018fb26} /* (24, 23, 30) {real, imag} */,
  {32'h3f65981c, 32'hc09e195c} /* (24, 23, 29) {real, imag} */,
  {32'hbea4c694, 32'hc05e2116} /* (24, 23, 28) {real, imag} */,
  {32'hbf51f6f4, 32'hc06a23fa} /* (24, 23, 27) {real, imag} */,
  {32'hbf72ce74, 32'hc0292778} /* (24, 23, 26) {real, imag} */,
  {32'hbf2a4682, 32'hbf2a07e3} /* (24, 23, 25) {real, imag} */,
  {32'hbffe303c, 32'h3e870d76} /* (24, 23, 24) {real, imag} */,
  {32'hc008c420, 32'hbf966de5} /* (24, 23, 23) {real, imag} */,
  {32'hc01ca0a2, 32'hbfcf408d} /* (24, 23, 22) {real, imag} */,
  {32'hbf383eb2, 32'h3f1f8cb9} /* (24, 23, 21) {real, imag} */,
  {32'h404c6448, 32'h4032777a} /* (24, 23, 20) {real, imag} */,
  {32'h40052754, 32'h3fd1f706} /* (24, 23, 19) {real, imag} */,
  {32'h401184bf, 32'h3e9c8622} /* (24, 23, 18) {real, imag} */,
  {32'h4023c6a4, 32'h4000123e} /* (24, 23, 17) {real, imag} */,
  {32'h3ffc654b, 32'h40234509} /* (24, 23, 16) {real, imag} */,
  {32'h3ecce3ec, 32'h401bc7ae} /* (24, 23, 15) {real, imag} */,
  {32'h40087ed0, 32'h3eed90e0} /* (24, 23, 14) {real, imag} */,
  {32'h4029c90a, 32'h3f958f9d} /* (24, 23, 13) {real, imag} */,
  {32'h400b50f6, 32'h3ef5932e} /* (24, 23, 12) {real, imag} */,
  {32'h3f8abf63, 32'h3d6eab90} /* (24, 23, 11) {real, imag} */,
  {32'hc01b9180, 32'hbfd808ff} /* (24, 23, 10) {real, imag} */,
  {32'hc03d7405, 32'hc07b722c} /* (24, 23, 9) {real, imag} */,
  {32'hc08e25da, 32'hbfe83b1a} /* (24, 23, 8) {real, imag} */,
  {32'hbf86418c, 32'hbfa6186a} /* (24, 23, 7) {real, imag} */,
  {32'hbfbeee80, 32'hc007bcb9} /* (24, 23, 6) {real, imag} */,
  {32'hbfccda96, 32'hc02a1319} /* (24, 23, 5) {real, imag} */,
  {32'h3d273440, 32'hbfe9606c} /* (24, 23, 4) {real, imag} */,
  {32'hbede4314, 32'hbf994940} /* (24, 23, 3) {real, imag} */,
  {32'hc012ab0c, 32'hbff80db9} /* (24, 23, 2) {real, imag} */,
  {32'hc053ae26, 32'hc0128207} /* (24, 23, 1) {real, imag} */,
  {32'hc0290bea, 32'hbfa0be16} /* (24, 23, 0) {real, imag} */,
  {32'hbf6cb19d, 32'hbfca3825} /* (24, 22, 31) {real, imag} */,
  {32'hbcf1a5c0, 32'hbfb77e34} /* (24, 22, 30) {real, imag} */,
  {32'hbe4637c4, 32'hbf6b53c6} /* (24, 22, 29) {real, imag} */,
  {32'hbfb30b9c, 32'hc019bf42} /* (24, 22, 28) {real, imag} */,
  {32'hbf895000, 32'hc01b5084} /* (24, 22, 27) {real, imag} */,
  {32'hc0287db9, 32'hbecb9570} /* (24, 22, 26) {real, imag} */,
  {32'hc0710e9a, 32'hbf48d27b} /* (24, 22, 25) {real, imag} */,
  {32'hc0366066, 32'hbeddee62} /* (24, 22, 24) {real, imag} */,
  {32'hc03c4c72, 32'hbf987504} /* (24, 22, 23) {real, imag} */,
  {32'hc04c2576, 32'hbfee1a88} /* (24, 22, 22) {real, imag} */,
  {32'h3e8346aa, 32'hbf09cd94} /* (24, 22, 21) {real, imag} */,
  {32'h40735bc6, 32'h3ff5c93b} /* (24, 22, 20) {real, imag} */,
  {32'h408ab9c3, 32'h4033b629} /* (24, 22, 19) {real, imag} */,
  {32'h400b3f54, 32'h3fa3323a} /* (24, 22, 18) {real, imag} */,
  {32'h3fbbaf50, 32'h3ff13b0c} /* (24, 22, 17) {real, imag} */,
  {32'h3ee015f2, 32'h408dd978} /* (24, 22, 16) {real, imag} */,
  {32'h3ffc70d4, 32'h40557e76} /* (24, 22, 15) {real, imag} */,
  {32'h404425ea, 32'h3f824568} /* (24, 22, 14) {real, imag} */,
  {32'h4076f892, 32'h3fe935c3} /* (24, 22, 13) {real, imag} */,
  {32'h3f967a8f, 32'h4048a4b4} /* (24, 22, 12) {real, imag} */,
  {32'h3f289662, 32'h4016f8d5} /* (24, 22, 11) {real, imag} */,
  {32'hbfe6d5b4, 32'hbfbb6627} /* (24, 22, 10) {real, imag} */,
  {32'hc03e85a5, 32'hc046cd3f} /* (24, 22, 9) {real, imag} */,
  {32'hc06128f7, 32'hc06afe66} /* (24, 22, 8) {real, imag} */,
  {32'hc029e028, 32'hbfd77921} /* (24, 22, 7) {real, imag} */,
  {32'hc075eaa8, 32'hc01166b9} /* (24, 22, 6) {real, imag} */,
  {32'hc043bb24, 32'hc00918dd} /* (24, 22, 5) {real, imag} */,
  {32'hc00cd918, 32'hc00ab2fa} /* (24, 22, 4) {real, imag} */,
  {32'hbfad91b4, 32'hbff313a9} /* (24, 22, 3) {real, imag} */,
  {32'hc025592c, 32'hbf3d3946} /* (24, 22, 2) {real, imag} */,
  {32'hc03d5b0e, 32'hbfb5f617} /* (24, 22, 1) {real, imag} */,
  {32'hbfe42941, 32'hbff84c7c} /* (24, 22, 0) {real, imag} */,
  {32'h3f192a4c, 32'hc007fcf3} /* (24, 21, 31) {real, imag} */,
  {32'hbe2b1aca, 32'hc0113857} /* (24, 21, 30) {real, imag} */,
  {32'hbf8a26aa, 32'hbedde5b2} /* (24, 21, 29) {real, imag} */,
  {32'hbfa1639f, 32'hc02b6ec0} /* (24, 21, 28) {real, imag} */,
  {32'hbf41722e, 32'hc065f7c4} /* (24, 21, 27) {real, imag} */,
  {32'hbfabe012, 32'hc0165123} /* (24, 21, 26) {real, imag} */,
  {32'hbfb4c298, 32'hbf7d4e00} /* (24, 21, 25) {real, imag} */,
  {32'hbf82e7a1, 32'h3f19c0e4} /* (24, 21, 24) {real, imag} */,
  {32'hbf7d4512, 32'hbea2d26a} /* (24, 21, 23) {real, imag} */,
  {32'hbf4c1225, 32'h3f2c9017} /* (24, 21, 22) {real, imag} */,
  {32'h3fb57cd3, 32'h3f79792c} /* (24, 21, 21) {real, imag} */,
  {32'hbe851faa, 32'h400d1962} /* (24, 21, 20) {real, imag} */,
  {32'hbb944ac0, 32'h3fb027f2} /* (24, 21, 19) {real, imag} */,
  {32'h3e666e80, 32'hbb956180} /* (24, 21, 18) {real, imag} */,
  {32'h3ece6b32, 32'hbf467e76} /* (24, 21, 17) {real, imag} */,
  {32'hbeaecdb4, 32'h3ed084fa} /* (24, 21, 16) {real, imag} */,
  {32'h3fb56476, 32'h3f5c6d02} /* (24, 21, 15) {real, imag} */,
  {32'h401dcfb0, 32'h3ef6e3fa} /* (24, 21, 14) {real, imag} */,
  {32'h3ff07350, 32'h3fb43bd2} /* (24, 21, 13) {real, imag} */,
  {32'h3dd6e1a0, 32'h405e3c28} /* (24, 21, 12) {real, imag} */,
  {32'hbf662b40, 32'h4008295e} /* (24, 21, 11) {real, imag} */,
  {32'hbef9fe4b, 32'h3d055948} /* (24, 21, 10) {real, imag} */,
  {32'hc00bed34, 32'hbfbc2528} /* (24, 21, 9) {real, imag} */,
  {32'hbfc2d176, 32'hbece589c} /* (24, 21, 8) {real, imag} */,
  {32'hbfeab9ea, 32'hbee5dd75} /* (24, 21, 7) {real, imag} */,
  {32'hc0817128, 32'hbfc1eb11} /* (24, 21, 6) {real, imag} */,
  {32'hc023fa59, 32'h3efae98a} /* (24, 21, 5) {real, imag} */,
  {32'hc002c59e, 32'hbdeedf50} /* (24, 21, 4) {real, imag} */,
  {32'hbfd37376, 32'hbeebfa28} /* (24, 21, 3) {real, imag} */,
  {32'hbf584d54, 32'h3f9208be} /* (24, 21, 2) {real, imag} */,
  {32'hbc198d80, 32'hbf811ece} /* (24, 21, 1) {real, imag} */,
  {32'hbf24dad4, 32'hbf65f520} /* (24, 21, 0) {real, imag} */,
  {32'h3fbb0387, 32'hbf8d1a84} /* (24, 20, 31) {real, imag} */,
  {32'h3f3334a0, 32'h3da9bc90} /* (24, 20, 30) {real, imag} */,
  {32'h3f915946, 32'h3f966ece} /* (24, 20, 29) {real, imag} */,
  {32'hbf071d58, 32'hbf86ff4e} /* (24, 20, 28) {real, imag} */,
  {32'hbc3cc700, 32'hbfeb42da} /* (24, 20, 27) {real, imag} */,
  {32'h400e504a, 32'hc017cffd} /* (24, 20, 26) {real, imag} */,
  {32'h40159e86, 32'hbd782680} /* (24, 20, 25) {real, imag} */,
  {32'h40112b94, 32'h400cfe19} /* (24, 20, 24) {real, imag} */,
  {32'h400acfb8, 32'h3ffbdb7f} /* (24, 20, 23) {real, imag} */,
  {32'h3ff21ed4, 32'h408140a8} /* (24, 20, 22) {real, imag} */,
  {32'h400e89bb, 32'h40590254} /* (24, 20, 21) {real, imag} */,
  {32'hbfa4a2e4, 32'h402c26ef} /* (24, 20, 20) {real, imag} */,
  {32'hbffb8f27, 32'h3f09f438} /* (24, 20, 19) {real, imag} */,
  {32'hbf14e90e, 32'hbff9fbe2} /* (24, 20, 18) {real, imag} */,
  {32'hbf4849db, 32'hc0309a47} /* (24, 20, 17) {real, imag} */,
  {32'hc01366f3, 32'hc05a83bf} /* (24, 20, 16) {real, imag} */,
  {32'hbfca909d, 32'hc05bcba4} /* (24, 20, 15) {real, imag} */,
  {32'hbee5dbcb, 32'hc0142636} /* (24, 20, 14) {real, imag} */,
  {32'hbf3c9b93, 32'hbf8eb2ce} /* (24, 20, 13) {real, imag} */,
  {32'hbf7c7ce5, 32'h3f5671c6} /* (24, 20, 12) {real, imag} */,
  {32'hbf50e62a, 32'h3df06c60} /* (24, 20, 11) {real, imag} */,
  {32'h3f9501ee, 32'h3f7da7d8} /* (24, 20, 10) {real, imag} */,
  {32'hbe6a3920, 32'h3fb27cb8} /* (24, 20, 9) {real, imag} */,
  {32'hbecfc20a, 32'h3f9a90d3} /* (24, 20, 8) {real, imag} */,
  {32'h3f52f954, 32'h3efc5e62} /* (24, 20, 7) {real, imag} */,
  {32'h3fa18f54, 32'h400664ea} /* (24, 20, 6) {real, imag} */,
  {32'h3e009c90, 32'h401e7f84} /* (24, 20, 5) {real, imag} */,
  {32'h3deedff8, 32'h3fe1532e} /* (24, 20, 4) {real, imag} */,
  {32'h3fa7260f, 32'h3f8a3751} /* (24, 20, 3) {real, imag} */,
  {32'h3f442d46, 32'h3fcb4702} /* (24, 20, 2) {real, imag} */,
  {32'h4001cf46, 32'h3fa62014} /* (24, 20, 1) {real, imag} */,
  {32'h3fcda652, 32'h3f389a89} /* (24, 20, 0) {real, imag} */,
  {32'h3f472eb4, 32'hbede304c} /* (24, 19, 31) {real, imag} */,
  {32'h3ffe46ef, 32'h3f3ecd41} /* (24, 19, 30) {real, imag} */,
  {32'h402edf5c, 32'h3f59ffa8} /* (24, 19, 29) {real, imag} */,
  {32'h3e94702c, 32'h3ce992c0} /* (24, 19, 28) {real, imag} */,
  {32'h3f458dc1, 32'h3f753bbe} /* (24, 19, 27) {real, imag} */,
  {32'h3febc7a1, 32'h40002af8} /* (24, 19, 26) {real, imag} */,
  {32'h3fcceac6, 32'h3ff911e0} /* (24, 19, 25) {real, imag} */,
  {32'h401f1bc0, 32'h3fc66b80} /* (24, 19, 24) {real, imag} */,
  {32'h4046ef40, 32'h40364ca9} /* (24, 19, 23) {real, imag} */,
  {32'h40586cba, 32'h4024dae9} /* (24, 19, 22) {real, imag} */,
  {32'h402e6326, 32'h3fc1c319} /* (24, 19, 21) {real, imag} */,
  {32'h3f4c68c1, 32'h3fb5d1e1} /* (24, 19, 20) {real, imag} */,
  {32'hbfebef17, 32'h3f737aa9} /* (24, 19, 19) {real, imag} */,
  {32'hbfe89754, 32'hbfaa8b1c} /* (24, 19, 18) {real, imag} */,
  {32'hc03f4516, 32'hc04f3385} /* (24, 19, 17) {real, imag} */,
  {32'hc0646340, 32'hc08a2f60} /* (24, 19, 16) {real, imag} */,
  {32'hc02be56e, 32'hc0a842e2} /* (24, 19, 15) {real, imag} */,
  {32'hbfce11e6, 32'hc0583aee} /* (24, 19, 14) {real, imag} */,
  {32'hbf877872, 32'hc0483d30} /* (24, 19, 13) {real, imag} */,
  {32'hc00cb08e, 32'hbf90c8f3} /* (24, 19, 12) {real, imag} */,
  {32'hc0127bcc, 32'h3eb257e0} /* (24, 19, 11) {real, imag} */,
  {32'h3f7f3ba0, 32'h3fe58341} /* (24, 19, 10) {real, imag} */,
  {32'h3eac64a8, 32'h3fc9c229} /* (24, 19, 9) {real, imag} */,
  {32'hbf11e529, 32'h3e81c3e8} /* (24, 19, 8) {real, imag} */,
  {32'h3f3d65cf, 32'hbf5a5f84} /* (24, 19, 7) {real, imag} */,
  {32'h3fe12e96, 32'h3f8a50f0} /* (24, 19, 6) {real, imag} */,
  {32'h3fb302d3, 32'h3f7d4f39} /* (24, 19, 5) {real, imag} */,
  {32'h401efe2a, 32'h3fe95713} /* (24, 19, 4) {real, imag} */,
  {32'h3faa1d24, 32'h40395ad5} /* (24, 19, 3) {real, imag} */,
  {32'hbf0a9a04, 32'h4001f870} /* (24, 19, 2) {real, imag} */,
  {32'h401ddc20, 32'h3f319c40} /* (24, 19, 1) {real, imag} */,
  {32'h3fec42f4, 32'hbde893d0} /* (24, 19, 0) {real, imag} */,
  {32'h3f0d929c, 32'h3f2527d4} /* (24, 18, 31) {real, imag} */,
  {32'h3ea94c1c, 32'h3fb1ee29} /* (24, 18, 30) {real, imag} */,
  {32'hbd10be00, 32'h3fc090ed} /* (24, 18, 29) {real, imag} */,
  {32'h3e3f85aa, 32'h3fc42553} /* (24, 18, 28) {real, imag} */,
  {32'h3f837958, 32'h4020cf72} /* (24, 18, 27) {real, imag} */,
  {32'h3e78bcd8, 32'h4014773e} /* (24, 18, 26) {real, imag} */,
  {32'h3ef8958c, 32'h3fdd6a52} /* (24, 18, 25) {real, imag} */,
  {32'h406d8dd2, 32'h3e936024} /* (24, 18, 24) {real, imag} */,
  {32'h3fce7c08, 32'h40170e36} /* (24, 18, 23) {real, imag} */,
  {32'h3fa11014, 32'h3fec940e} /* (24, 18, 22) {real, imag} */,
  {32'h4030189e, 32'hbfac2285} /* (24, 18, 21) {real, imag} */,
  {32'h3edaa36e, 32'h3fb5a752} /* (24, 18, 20) {real, imag} */,
  {32'hbfc68f5a, 32'h3ed1fe64} /* (24, 18, 19) {real, imag} */,
  {32'hbece286c, 32'hbfb94988} /* (24, 18, 18) {real, imag} */,
  {32'hc05b19ab, 32'hc05047d1} /* (24, 18, 17) {real, imag} */,
  {32'hc02c2cb7, 32'hc02c4176} /* (24, 18, 16) {real, imag} */,
  {32'hc012a841, 32'hc013cf91} /* (24, 18, 15) {real, imag} */,
  {32'hbf9d138e, 32'hbfa2ae92} /* (24, 18, 14) {real, imag} */,
  {32'hbf7e5dd8, 32'hc0111b62} /* (24, 18, 13) {real, imag} */,
  {32'hbf4ba73f, 32'hbd37f3d0} /* (24, 18, 12) {real, imag} */,
  {32'hbfb99ff3, 32'h3f6d1c9d} /* (24, 18, 11) {real, imag} */,
  {32'h4015b803, 32'h3f109e1b} /* (24, 18, 10) {real, imag} */,
  {32'h3fdbc64d, 32'h3f178c22} /* (24, 18, 9) {real, imag} */,
  {32'h3f14f499, 32'h3fac21b8} /* (24, 18, 8) {real, imag} */,
  {32'h3f426eee, 32'h404cc86f} /* (24, 18, 7) {real, imag} */,
  {32'h4012f465, 32'h407d8850} /* (24, 18, 6) {real, imag} */,
  {32'h405e62d1, 32'h3fce0c86} /* (24, 18, 5) {real, imag} */,
  {32'h4070957c, 32'hbf1fbbc6} /* (24, 18, 4) {real, imag} */,
  {32'h3ffbfe46, 32'h3f887961} /* (24, 18, 3) {real, imag} */,
  {32'hbf4f577a, 32'h401c9248} /* (24, 18, 2) {real, imag} */,
  {32'h40135098, 32'h3f0d1c2d} /* (24, 18, 1) {real, imag} */,
  {32'h401274ea, 32'hbf879d46} /* (24, 18, 0) {real, imag} */,
  {32'h3f550cda, 32'hbed465ae} /* (24, 17, 31) {real, imag} */,
  {32'hbf03c1cc, 32'h3f102b78} /* (24, 17, 30) {real, imag} */,
  {32'hbfc15ea5, 32'h3ed01c90} /* (24, 17, 29) {real, imag} */,
  {32'h3c8bf200, 32'h3ec6089a} /* (24, 17, 28) {real, imag} */,
  {32'h40071424, 32'h3fc62591} /* (24, 17, 27) {real, imag} */,
  {32'h3fbc5da1, 32'h3f9da03b} /* (24, 17, 26) {real, imag} */,
  {32'h4028afe6, 32'h40432088} /* (24, 17, 25) {real, imag} */,
  {32'h40495904, 32'h40152b9e} /* (24, 17, 24) {real, imag} */,
  {32'hbf9044b9, 32'h4039e5ca} /* (24, 17, 23) {real, imag} */,
  {32'h3fdd40ae, 32'h3ffc5d1e} /* (24, 17, 22) {real, imag} */,
  {32'h4055c3a4, 32'h3f6b4244} /* (24, 17, 21) {real, imag} */,
  {32'hbe81addc, 32'h3f95d64c} /* (24, 17, 20) {real, imag} */,
  {32'hbff9a458, 32'hbffb96a3} /* (24, 17, 19) {real, imag} */,
  {32'hbf966340, 32'hc080510e} /* (24, 17, 18) {real, imag} */,
  {32'hc024b22c, 32'hc048c814} /* (24, 17, 17) {real, imag} */,
  {32'hc03c0316, 32'hbf057412} /* (24, 17, 16) {real, imag} */,
  {32'hc066fa88, 32'hbe36fe60} /* (24, 17, 15) {real, imag} */,
  {32'hc0467a48, 32'hbfb25e39} /* (24, 17, 14) {real, imag} */,
  {32'hbfe3a2a6, 32'hc0294086} /* (24, 17, 13) {real, imag} */,
  {32'hbf878f43, 32'hbfc683b5} /* (24, 17, 12) {real, imag} */,
  {32'hbfc8e971, 32'h3eb18f5c} /* (24, 17, 11) {real, imag} */,
  {32'h4050e823, 32'h405b8dd3} /* (24, 17, 10) {real, imag} */,
  {32'h403d4a6b, 32'h400d8286} /* (24, 17, 9) {real, imag} */,
  {32'h3f23675c, 32'h3fd2c556} /* (24, 17, 8) {real, imag} */,
  {32'h3ecf2cf2, 32'h40499ee7} /* (24, 17, 7) {real, imag} */,
  {32'h3fca6ec1, 32'h408e491c} /* (24, 17, 6) {real, imag} */,
  {32'h4080e41c, 32'h404800aa} /* (24, 17, 5) {real, imag} */,
  {32'h402fbc78, 32'h3f574382} /* (24, 17, 4) {real, imag} */,
  {32'h3f6aac10, 32'h40229ee0} /* (24, 17, 3) {real, imag} */,
  {32'h3ffd9650, 32'h405dc63a} /* (24, 17, 2) {real, imag} */,
  {32'h406fbdeb, 32'h40140f37} /* (24, 17, 1) {real, imag} */,
  {32'h401b617e, 32'h3e85ee08} /* (24, 17, 0) {real, imag} */,
  {32'h3d2aba20, 32'h3e391dbc} /* (24, 16, 31) {real, imag} */,
  {32'hbdefd530, 32'h3f484c5b} /* (24, 16, 30) {real, imag} */,
  {32'h3fca8cf3, 32'h3fb2015d} /* (24, 16, 29) {real, imag} */,
  {32'h3f7e60ab, 32'h3fad0237} /* (24, 16, 28) {real, imag} */,
  {32'h403f1a06, 32'h3f0e60a7} /* (24, 16, 27) {real, imag} */,
  {32'h3f7e632a, 32'h4011c2a0} /* (24, 16, 26) {real, imag} */,
  {32'h3f8e5ad4, 32'h4045d01e} /* (24, 16, 25) {real, imag} */,
  {32'h3fb9feac, 32'h3fd3706e} /* (24, 16, 24) {real, imag} */,
  {32'hbe03d54c, 32'h401650e8} /* (24, 16, 23) {real, imag} */,
  {32'h4006a772, 32'h40096410} /* (24, 16, 22) {real, imag} */,
  {32'h3fb9f30a, 32'h3fc52de0} /* (24, 16, 21) {real, imag} */,
  {32'hbe5292f0, 32'h3f5c1c97} /* (24, 16, 20) {real, imag} */,
  {32'hc01d4e98, 32'hc025ef0e} /* (24, 16, 19) {real, imag} */,
  {32'hbf257b53, 32'hc0164501} /* (24, 16, 18) {real, imag} */,
  {32'hbf868a00, 32'hbf280162} /* (24, 16, 17) {real, imag} */,
  {32'hc03e7f05, 32'h3f008212} /* (24, 16, 16) {real, imag} */,
  {32'hc04b4340, 32'h3ee1d428} /* (24, 16, 15) {real, imag} */,
  {32'hc06c4866, 32'hbfe0a58a} /* (24, 16, 14) {real, imag} */,
  {32'hc03eca37, 32'hc04c91d8} /* (24, 16, 13) {real, imag} */,
  {32'hc06d6552, 32'hc0203290} /* (24, 16, 12) {real, imag} */,
  {32'hc00ddd5c, 32'hbf012fa0} /* (24, 16, 11) {real, imag} */,
  {32'h3ff6f2f8, 32'h40525d22} /* (24, 16, 10) {real, imag} */,
  {32'h401663ea, 32'h403d17e1} /* (24, 16, 9) {real, imag} */,
  {32'h3ffc8c41, 32'h400a9d06} /* (24, 16, 8) {real, imag} */,
  {32'h3ff0ff14, 32'h405d3610} /* (24, 16, 7) {real, imag} */,
  {32'h3f77c1ac, 32'h40b7c6ce} /* (24, 16, 6) {real, imag} */,
  {32'h403d3d4c, 32'h406a9e28} /* (24, 16, 5) {real, imag} */,
  {32'h40166dce, 32'h400d5ae2} /* (24, 16, 4) {real, imag} */,
  {32'h4005e4ea, 32'h3fda93a6} /* (24, 16, 3) {real, imag} */,
  {32'h409fcbf8, 32'h3fe2e62c} /* (24, 16, 2) {real, imag} */,
  {32'h40424c5b, 32'h403e4ce0} /* (24, 16, 1) {real, imag} */,
  {32'h3f9638dc, 32'h400c7a43} /* (24, 16, 0) {real, imag} */,
  {32'h3ea1fee2, 32'h3f60a4fd} /* (24, 15, 31) {real, imag} */,
  {32'h40079e42, 32'h40023428} /* (24, 15, 30) {real, imag} */,
  {32'h40792916, 32'h405fd0b0} /* (24, 15, 29) {real, imag} */,
  {32'h40129747, 32'h40302756} /* (24, 15, 28) {real, imag} */,
  {32'h40389a07, 32'h3fc2aadf} /* (24, 15, 27) {real, imag} */,
  {32'h3f8206d2, 32'h40415238} /* (24, 15, 26) {real, imag} */,
  {32'h3f0a2028, 32'h40314342} /* (24, 15, 25) {real, imag} */,
  {32'hbfb51689, 32'h3f1c9cbb} /* (24, 15, 24) {real, imag} */,
  {32'h3fc28ead, 32'h3f43b62a} /* (24, 15, 23) {real, imag} */,
  {32'h4020812c, 32'h3fac925a} /* (24, 15, 22) {real, imag} */,
  {32'h3f26f538, 32'h3ef12188} /* (24, 15, 21) {real, imag} */,
  {32'hbf9e35cc, 32'h3ec8c992} /* (24, 15, 20) {real, imag} */,
  {32'hc0296e24, 32'hbf853953} /* (24, 15, 19) {real, imag} */,
  {32'h3f01480b, 32'hbf98a9a1} /* (24, 15, 18) {real, imag} */,
  {32'h3fcdee00, 32'hbfa53c21} /* (24, 15, 17) {real, imag} */,
  {32'hc000dfae, 32'hbf8140bf} /* (24, 15, 16) {real, imag} */,
  {32'hc058c865, 32'hbfbb662b} /* (24, 15, 15) {real, imag} */,
  {32'hc049ab4e, 32'hbfb9b99b} /* (24, 15, 14) {real, imag} */,
  {32'hc02465c0, 32'hc0321b74} /* (24, 15, 13) {real, imag} */,
  {32'hbfe5ed86, 32'hc0033502} /* (24, 15, 12) {real, imag} */,
  {32'hbe16c150, 32'hbf9587f8} /* (24, 15, 11) {real, imag} */,
  {32'h3fffa1d5, 32'h3ffc36a0} /* (24, 15, 10) {real, imag} */,
  {32'h402b1e80, 32'h4080e82e} /* (24, 15, 9) {real, imag} */,
  {32'h3f92b804, 32'h3f8ef401} /* (24, 15, 8) {real, imag} */,
  {32'h3ee8fa48, 32'h3eb6a368} /* (24, 15, 7) {real, imag} */,
  {32'h3fd26ddc, 32'h401605f0} /* (24, 15, 6) {real, imag} */,
  {32'h4078a8c5, 32'h40249826} /* (24, 15, 5) {real, imag} */,
  {32'h401fc872, 32'h407630f8} /* (24, 15, 4) {real, imag} */,
  {32'h4071a139, 32'h3fee5b58} /* (24, 15, 3) {real, imag} */,
  {32'h40b8b2f0, 32'h3fd10475} /* (24, 15, 2) {real, imag} */,
  {32'h4018c947, 32'h40655f61} /* (24, 15, 1) {real, imag} */,
  {32'hbc949be0, 32'h3f3716a2} /* (24, 15, 0) {real, imag} */,
  {32'h3f42d5d8, 32'h3f7c4e8a} /* (24, 14, 31) {real, imag} */,
  {32'h3ff2f50e, 32'h407a4872} /* (24, 14, 30) {real, imag} */,
  {32'h4043ec25, 32'h40b80fde} /* (24, 14, 29) {real, imag} */,
  {32'h404a5f03, 32'h406a98b2} /* (24, 14, 28) {real, imag} */,
  {32'h401e01cf, 32'h40631799} /* (24, 14, 27) {real, imag} */,
  {32'h3ee046ac, 32'h407f5108} /* (24, 14, 26) {real, imag} */,
  {32'h3f8e1a83, 32'h4052e1ac} /* (24, 14, 25) {real, imag} */,
  {32'h3f4aaf18, 32'hbf2d0964} /* (24, 14, 24) {real, imag} */,
  {32'h3ff61fc7, 32'hbeb7b048} /* (24, 14, 23) {real, imag} */,
  {32'h3f4d856c, 32'h3fafc050} /* (24, 14, 22) {real, imag} */,
  {32'hbd09f490, 32'h3fc6e1c0} /* (24, 14, 21) {real, imag} */,
  {32'hc0296a11, 32'hbe3047a0} /* (24, 14, 20) {real, imag} */,
  {32'hc01a6d02, 32'hc01b5df4} /* (24, 14, 19) {real, imag} */,
  {32'hbe4ee388, 32'hc05fbf78} /* (24, 14, 18) {real, imag} */,
  {32'hbf0621f8, 32'hc03a4cf8} /* (24, 14, 17) {real, imag} */,
  {32'hbfcd0e82, 32'hbf9a7f62} /* (24, 14, 16) {real, imag} */,
  {32'hbffe2876, 32'hc0272b0a} /* (24, 14, 15) {real, imag} */,
  {32'hbf71b7fc, 32'hbffe24ae} /* (24, 14, 14) {real, imag} */,
  {32'hbf85bbdc, 32'hc0349d82} /* (24, 14, 13) {real, imag} */,
  {32'hbf1b9233, 32'hc0448604} /* (24, 14, 12) {real, imag} */,
  {32'hbe3fe4f0, 32'hbfde4db1} /* (24, 14, 11) {real, imag} */,
  {32'h3fe1920b, 32'h3df01b8c} /* (24, 14, 10) {real, imag} */,
  {32'h3fedfe54, 32'h3fd27c9e} /* (24, 14, 9) {real, imag} */,
  {32'h3ddbeb38, 32'h3fca51d6} /* (24, 14, 8) {real, imag} */,
  {32'hbd851318, 32'h3fecf4b2} /* (24, 14, 7) {real, imag} */,
  {32'h40199e7d, 32'h3f9eb2fb} /* (24, 14, 6) {real, imag} */,
  {32'h409f99e7, 32'h3f96a133} /* (24, 14, 5) {real, imag} */,
  {32'h405e64be, 32'h402f8947} /* (24, 14, 4) {real, imag} */,
  {32'h400fdc76, 32'h3fb78f4c} /* (24, 14, 3) {real, imag} */,
  {32'h3f493394, 32'h4013b9e4} /* (24, 14, 2) {real, imag} */,
  {32'hbf2d41b2, 32'h4043ef4a} /* (24, 14, 1) {real, imag} */,
  {32'hbf8bc9a6, 32'hbef40ae9} /* (24, 14, 0) {real, imag} */,
  {32'h3e125e98, 32'h3fa9c622} /* (24, 13, 31) {real, imag} */,
  {32'h3e66ba5c, 32'h4047e717} /* (24, 13, 30) {real, imag} */,
  {32'h3f55bfe4, 32'h405fe2ba} /* (24, 13, 29) {real, imag} */,
  {32'h3fc77d9c, 32'h401763d8} /* (24, 13, 28) {real, imag} */,
  {32'h40774740, 32'h40836a73} /* (24, 13, 27) {real, imag} */,
  {32'h4005dcf9, 32'h40879b2c} /* (24, 13, 26) {real, imag} */,
  {32'h3fd6f842, 32'h403c1e33} /* (24, 13, 25) {real, imag} */,
  {32'h4062e27e, 32'h3ee16bbc} /* (24, 13, 24) {real, imag} */,
  {32'h401f6c7e, 32'h3fed872e} /* (24, 13, 23) {real, imag} */,
  {32'h3ebf8baa, 32'h4088236a} /* (24, 13, 22) {real, imag} */,
  {32'h3f80551b, 32'h4015ed22} /* (24, 13, 21) {real, imag} */,
  {32'hc006070e, 32'h3eddc5c2} /* (24, 13, 20) {real, imag} */,
  {32'hc0241084, 32'hc0038140} /* (24, 13, 19) {real, imag} */,
  {32'hbfd8f870, 32'hc0710cb0} /* (24, 13, 18) {real, imag} */,
  {32'hbf8deec4, 32'hc040ece9} /* (24, 13, 17) {real, imag} */,
  {32'h3eaedff4, 32'hc0805316} /* (24, 13, 16) {real, imag} */,
  {32'h3e32d778, 32'hc0476776} /* (24, 13, 15) {real, imag} */,
  {32'h3f7967d3, 32'hbfed3de6} /* (24, 13, 14) {real, imag} */,
  {32'hbfe64bbe, 32'hbb8ed180} /* (24, 13, 13) {real, imag} */,
  {32'hbfedabd1, 32'hbf7efcbb} /* (24, 13, 12) {real, imag} */,
  {32'hbfc6e250, 32'hbfd3370e} /* (24, 13, 11) {real, imag} */,
  {32'hbe5236ec, 32'h3eafa781} /* (24, 13, 10) {real, imag} */,
  {32'h3f8a2938, 32'h40043c91} /* (24, 13, 9) {real, imag} */,
  {32'h3ffe9ac7, 32'h40319b00} /* (24, 13, 8) {real, imag} */,
  {32'h4066e5d6, 32'h3fde31f2} /* (24, 13, 7) {real, imag} */,
  {32'h405d3ac2, 32'h4014fd16} /* (24, 13, 6) {real, imag} */,
  {32'h40286ffc, 32'h3ffe1d46} /* (24, 13, 5) {real, imag} */,
  {32'h40683378, 32'h40251810} /* (24, 13, 4) {real, imag} */,
  {32'h4060a390, 32'h3fed1e3b} /* (24, 13, 3) {real, imag} */,
  {32'h3eeedf60, 32'h403a70bc} /* (24, 13, 2) {real, imag} */,
  {32'h3d905840, 32'h3fc9c2b8} /* (24, 13, 1) {real, imag} */,
  {32'hbdf19b00, 32'h3f01e73f} /* (24, 13, 0) {real, imag} */,
  {32'h3f30e725, 32'h40011c2c} /* (24, 12, 31) {real, imag} */,
  {32'h3faa9ce7, 32'h3ff43e04} /* (24, 12, 30) {real, imag} */,
  {32'h3f405386, 32'h3f86c499} /* (24, 12, 29) {real, imag} */,
  {32'hbf67b75c, 32'h3f88145a} /* (24, 12, 28) {real, imag} */,
  {32'h3fcbdf9b, 32'h3fe4ac86} /* (24, 12, 27) {real, imag} */,
  {32'h4028326e, 32'h40020680} /* (24, 12, 26) {real, imag} */,
  {32'h3ff93417, 32'h4076634a} /* (24, 12, 25) {real, imag} */,
  {32'h402a9670, 32'h40626580} /* (24, 12, 24) {real, imag} */,
  {32'h3fd80655, 32'h408a9b33} /* (24, 12, 23) {real, imag} */,
  {32'h401f903c, 32'h40935b13} /* (24, 12, 22) {real, imag} */,
  {32'h4061fdfc, 32'h3fd09ff0} /* (24, 12, 21) {real, imag} */,
  {32'h3e945e2e, 32'hbbc22f00} /* (24, 12, 20) {real, imag} */,
  {32'hc00895ca, 32'hbec2fd78} /* (24, 12, 19) {real, imag} */,
  {32'hc0083d6b, 32'hc0147b36} /* (24, 12, 18) {real, imag} */,
  {32'hc00266a8, 32'hc0341daa} /* (24, 12, 17) {real, imag} */,
  {32'hbf51ee04, 32'hc0559df2} /* (24, 12, 16) {real, imag} */,
  {32'hbf67fecc, 32'hbffa6384} /* (24, 12, 15) {real, imag} */,
  {32'hbed50a88, 32'hc0002d01} /* (24, 12, 14) {real, imag} */,
  {32'hc022f4ee, 32'h3cbf48e0} /* (24, 12, 13) {real, imag} */,
  {32'hbff67c90, 32'hbe849d28} /* (24, 12, 12) {real, imag} */,
  {32'h3eb48870, 32'hbf5bc556} /* (24, 12, 11) {real, imag} */,
  {32'h3faed33a, 32'h40145a06} /* (24, 12, 10) {real, imag} */,
  {32'h3fd921be, 32'h400364ee} /* (24, 12, 9) {real, imag} */,
  {32'h40299991, 32'h3ff6a152} /* (24, 12, 8) {real, imag} */,
  {32'h400a4f7b, 32'h3f8715d4} /* (24, 12, 7) {real, imag} */,
  {32'h3fc6fd31, 32'h400d7ee4} /* (24, 12, 6) {real, imag} */,
  {32'h3f194286, 32'h4031bd0a} /* (24, 12, 5) {real, imag} */,
  {32'h4021f3f2, 32'h403e90e4} /* (24, 12, 4) {real, imag} */,
  {32'h3fceeaa1, 32'h3f886f30} /* (24, 12, 3) {real, imag} */,
  {32'h3fdfb464, 32'h3f52b928} /* (24, 12, 2) {real, imag} */,
  {32'h3fec5a98, 32'h3f8192c9} /* (24, 12, 1) {real, imag} */,
  {32'h3f7e03c5, 32'h3f8fdc82} /* (24, 12, 0) {real, imag} */,
  {32'h3bab4200, 32'h3fd79722} /* (24, 11, 31) {real, imag} */,
  {32'h3f926dd8, 32'h3fc2f820} /* (24, 11, 30) {real, imag} */,
  {32'h40371931, 32'h3f86c480} /* (24, 11, 29) {real, imag} */,
  {32'h400b1bf2, 32'h3afd5800} /* (24, 11, 28) {real, imag} */,
  {32'h3ff9b382, 32'hbef44294} /* (24, 11, 27) {real, imag} */,
  {32'h402b4dce, 32'h3e6c5640} /* (24, 11, 26) {real, imag} */,
  {32'h3ff69f20, 32'h40563b15} /* (24, 11, 25) {real, imag} */,
  {32'h3efd28e2, 32'h404663b6} /* (24, 11, 24) {real, imag} */,
  {32'h3f81c942, 32'h408b8e35} /* (24, 11, 23) {real, imag} */,
  {32'h402a6b5a, 32'h40871c47} /* (24, 11, 22) {real, imag} */,
  {32'h401f703a, 32'hbeaa71a4} /* (24, 11, 21) {real, imag} */,
  {32'hbed37b6c, 32'hbf93e50e} /* (24, 11, 20) {real, imag} */,
  {32'hbfe35caa, 32'h3e13a91c} /* (24, 11, 19) {real, imag} */,
  {32'hc04d9881, 32'hc0138ea0} /* (24, 11, 18) {real, imag} */,
  {32'hc084c2af, 32'hc02cd2ae} /* (24, 11, 17) {real, imag} */,
  {32'hc011ba02, 32'hc040440c} /* (24, 11, 16) {real, imag} */,
  {32'hbfe0672e, 32'hbfeffb46} /* (24, 11, 15) {real, imag} */,
  {32'hbbeb9c80, 32'hbfa94e60} /* (24, 11, 14) {real, imag} */,
  {32'h3ee2dad4, 32'h3e4cf1f4} /* (24, 11, 13) {real, imag} */,
  {32'hbea2ce6d, 32'hbfaf044e} /* (24, 11, 12) {real, imag} */,
  {32'h3f0250d5, 32'hc002400e} /* (24, 11, 11) {real, imag} */,
  {32'h3f22bae1, 32'h3f11e448} /* (24, 11, 10) {real, imag} */,
  {32'h3f8d79e6, 32'h3f122e74} /* (24, 11, 9) {real, imag} */,
  {32'h3eafb5b0, 32'h40038ac4} /* (24, 11, 8) {real, imag} */,
  {32'hbf45d808, 32'h3fd757fc} /* (24, 11, 7) {real, imag} */,
  {32'h3f48b6ea, 32'h3fb7ba70} /* (24, 11, 6) {real, imag} */,
  {32'h3f1cd990, 32'h4076cfa7} /* (24, 11, 5) {real, imag} */,
  {32'h3e903ea8, 32'h401142eb} /* (24, 11, 4) {real, imag} */,
  {32'h3f957454, 32'hbd7f47b0} /* (24, 11, 3) {real, imag} */,
  {32'h3f27e993, 32'hbe9c5fce} /* (24, 11, 2) {real, imag} */,
  {32'hbdc95e58, 32'h4016f962} /* (24, 11, 1) {real, imag} */,
  {32'hbe4af45c, 32'h3ff5afc9} /* (24, 11, 0) {real, imag} */,
  {32'hbf5ade30, 32'h3f5dfa30} /* (24, 10, 31) {real, imag} */,
  {32'hbfce97f7, 32'h3f154d00} /* (24, 10, 30) {real, imag} */,
  {32'hbf98c817, 32'h3e8e0ba6} /* (24, 10, 29) {real, imag} */,
  {32'hbdde2d30, 32'h3ecd1302} /* (24, 10, 28) {real, imag} */,
  {32'hbf9d8ffa, 32'hbefc3498} /* (24, 10, 27) {real, imag} */,
  {32'hbfb6d8e0, 32'hbfc00ab1} /* (24, 10, 26) {real, imag} */,
  {32'h3e202e80, 32'hbf88e666} /* (24, 10, 25) {real, imag} */,
  {32'hbe3fab04, 32'h3fc9f762} /* (24, 10, 24) {real, imag} */,
  {32'hbf7575b1, 32'h40289f0e} /* (24, 10, 23) {real, imag} */,
  {32'hbf857610, 32'hbea0adae} /* (24, 10, 22) {real, imag} */,
  {32'hbf67790c, 32'hc0785870} /* (24, 10, 21) {real, imag} */,
  {32'hbdec76a0, 32'hbea65db0} /* (24, 10, 20) {real, imag} */,
  {32'h3fc6a52f, 32'h400afe52} /* (24, 10, 19) {real, imag} */,
  {32'hbefcc588, 32'hbfcbe24b} /* (24, 10, 18) {real, imag} */,
  {32'hbf681bc4, 32'hbe7a8e18} /* (24, 10, 17) {real, imag} */,
  {32'h3fba3a39, 32'h3ecd2406} /* (24, 10, 16) {real, imag} */,
  {32'h3ffabc42, 32'h3fa2661f} /* (24, 10, 15) {real, imag} */,
  {32'h3fc931e4, 32'h3e8594e9} /* (24, 10, 14) {real, imag} */,
  {32'h3f1c0996, 32'h3fee0d6c} /* (24, 10, 13) {real, imag} */,
  {32'h3f28f448, 32'hbeac4ba6} /* (24, 10, 12) {real, imag} */,
  {32'hbf009212, 32'h3f2363c6} /* (24, 10, 11) {real, imag} */,
  {32'hbe6ab3cc, 32'hbf239800} /* (24, 10, 10) {real, imag} */,
  {32'hbf8eae55, 32'hc05b2a05} /* (24, 10, 9) {real, imag} */,
  {32'hc0017c80, 32'hc0272fb7} /* (24, 10, 8) {real, imag} */,
  {32'hc04029c9, 32'hc0088d1c} /* (24, 10, 7) {real, imag} */,
  {32'hbffadb42, 32'hbfb1a245} /* (24, 10, 6) {real, imag} */,
  {32'hbf1e90ff, 32'h3e726d00} /* (24, 10, 5) {real, imag} */,
  {32'hbfb8b534, 32'h3f3a77de} /* (24, 10, 4) {real, imag} */,
  {32'hbfe30a22, 32'h3f99c7f8} /* (24, 10, 3) {real, imag} */,
  {32'hc00f46ea, 32'hbfa13f50} /* (24, 10, 2) {real, imag} */,
  {32'hbf8f116c, 32'hbfd18ea0} /* (24, 10, 1) {real, imag} */,
  {32'hbf533350, 32'hbea7a952} /* (24, 10, 0) {real, imag} */,
  {32'h3d9c4128, 32'hbfa5c0c2} /* (24, 9, 31) {real, imag} */,
  {32'hc001dc16, 32'hbf10c832} /* (24, 9, 30) {real, imag} */,
  {32'hc0265af9, 32'h3caabe80} /* (24, 9, 29) {real, imag} */,
  {32'hc01abbc7, 32'h3e7ff190} /* (24, 9, 28) {real, imag} */,
  {32'hc0848f46, 32'hbf4a28fb} /* (24, 9, 27) {real, imag} */,
  {32'hc0450942, 32'hc0164118} /* (24, 9, 26) {real, imag} */,
  {32'hbdce2358, 32'hc012603a} /* (24, 9, 25) {real, imag} */,
  {32'hbeb1d9d8, 32'hbeb11464} /* (24, 9, 24) {real, imag} */,
  {32'hc014786e, 32'hbe041d00} /* (24, 9, 23) {real, imag} */,
  {32'hc03774fc, 32'hc065a411} /* (24, 9, 22) {real, imag} */,
  {32'hc0000426, 32'hc080bf08} /* (24, 9, 21) {real, imag} */,
  {32'h3fa7a90e, 32'h3f432c90} /* (24, 9, 20) {real, imag} */,
  {32'h40299260, 32'h4026f6da} /* (24, 9, 19) {real, imag} */,
  {32'h3fd75553, 32'hbec7c3da} /* (24, 9, 18) {real, imag} */,
  {32'h3fde3f4f, 32'hbec9642a} /* (24, 9, 17) {real, imag} */,
  {32'h4047865e, 32'h3fa58fdf} /* (24, 9, 16) {real, imag} */,
  {32'h4027a8e8, 32'h3ff24afe} /* (24, 9, 15) {real, imag} */,
  {32'h4009283e, 32'hbedf1200} /* (24, 9, 14) {real, imag} */,
  {32'hbef4af40, 32'h3f6eb45c} /* (24, 9, 13) {real, imag} */,
  {32'h3fcb2eb6, 32'hbfdae580} /* (24, 9, 12) {real, imag} */,
  {32'h3fbda60e, 32'h3f34c9c3} /* (24, 9, 11) {real, imag} */,
  {32'h3e941183, 32'h3f51f754} /* (24, 9, 10) {real, imag} */,
  {32'hbf9b1c0e, 32'hc02e374a} /* (24, 9, 9) {real, imag} */,
  {32'hc040784e, 32'hc08a3750} /* (24, 9, 8) {real, imag} */,
  {32'hc06384bd, 32'hc06283a4} /* (24, 9, 7) {real, imag} */,
  {32'hc003bc94, 32'hbff30a9e} /* (24, 9, 6) {real, imag} */,
  {32'hbfa45eb7, 32'hbfb12a46} /* (24, 9, 5) {real, imag} */,
  {32'hbeb2e716, 32'hbf914973} /* (24, 9, 4) {real, imag} */,
  {32'hbfed8272, 32'hbe559048} /* (24, 9, 3) {real, imag} */,
  {32'hc04ac0ff, 32'hc01a7df4} /* (24, 9, 2) {real, imag} */,
  {32'hbfea47c2, 32'hc0539c46} /* (24, 9, 1) {real, imag} */,
  {32'hbeff1ce8, 32'hbff6e7e4} /* (24, 9, 0) {real, imag} */,
  {32'h3f669044, 32'hbc9ad070} /* (24, 8, 31) {real, imag} */,
  {32'h3e4a7e9a, 32'hbf5fdb60} /* (24, 8, 30) {real, imag} */,
  {32'hbf20d376, 32'hbfbce18c} /* (24, 8, 29) {real, imag} */,
  {32'hbecb38de, 32'hbfd745a8} /* (24, 8, 28) {real, imag} */,
  {32'hbfd097e7, 32'hbf80b27d} /* (24, 8, 27) {real, imag} */,
  {32'hbfd174b4, 32'hc01d2b2a} /* (24, 8, 26) {real, imag} */,
  {32'hbf35f0c0, 32'hc081e25a} /* (24, 8, 25) {real, imag} */,
  {32'h3f7a41bc, 32'hbf89e0b0} /* (24, 8, 24) {real, imag} */,
  {32'hbf845c45, 32'hbf83b85e} /* (24, 8, 23) {real, imag} */,
  {32'hc0429d8c, 32'hc0827548} /* (24, 8, 22) {real, imag} */,
  {32'hbf1397ad, 32'hc00ef4c6} /* (24, 8, 21) {real, imag} */,
  {32'h3fae22a6, 32'h3f5d3c46} /* (24, 8, 20) {real, imag} */,
  {32'h3fece4c2, 32'h3fbedc8c} /* (24, 8, 19) {real, imag} */,
  {32'h3ed8975c, 32'h40108263} /* (24, 8, 18) {real, imag} */,
  {32'h3f86cc18, 32'h401b2aec} /* (24, 8, 17) {real, imag} */,
  {32'h4068480f, 32'h40508222} /* (24, 8, 16) {real, imag} */,
  {32'h4041954e, 32'h401bcced} /* (24, 8, 15) {real, imag} */,
  {32'h4038cca2, 32'h3d36d380} /* (24, 8, 14) {real, imag} */,
  {32'h40456649, 32'hbe7fe214} /* (24, 8, 13) {real, imag} */,
  {32'h40840a10, 32'hbf2fe880} /* (24, 8, 12) {real, imag} */,
  {32'h40449c99, 32'h3f6bfaf7} /* (24, 8, 11) {real, imag} */,
  {32'h3fcdcba4, 32'h3f698e62} /* (24, 8, 10) {real, imag} */,
  {32'h3eb1078d, 32'hbf62e16a} /* (24, 8, 9) {real, imag} */,
  {32'hbfc8b6d0, 32'hbf984370} /* (24, 8, 8) {real, imag} */,
  {32'hc080497e, 32'hbf14cdbb} /* (24, 8, 7) {real, imag} */,
  {32'hc06455a1, 32'hbfabe074} /* (24, 8, 6) {real, imag} */,
  {32'hbffeae86, 32'hc03f7df0} /* (24, 8, 5) {real, imag} */,
  {32'hbf8aa352, 32'hbfd1019a} /* (24, 8, 4) {real, imag} */,
  {32'hc0054324, 32'h3f2a9ec0} /* (24, 8, 3) {real, imag} */,
  {32'hc0625d86, 32'hbfc13b4a} /* (24, 8, 2) {real, imag} */,
  {32'hc084397b, 32'hc0065452} /* (24, 8, 1) {real, imag} */,
  {32'hbfc2681a, 32'hbf8d05ed} /* (24, 8, 0) {real, imag} */,
  {32'hbfbed5c6, 32'hc01a0f72} /* (24, 7, 31) {real, imag} */,
  {32'hbea369f8, 32'hc0880462} /* (24, 7, 30) {real, imag} */,
  {32'h3ee75ca0, 32'hc052aaf1} /* (24, 7, 29) {real, imag} */,
  {32'hbd20fa20, 32'hbfd01215} /* (24, 7, 28) {real, imag} */,
  {32'hbf05f7b0, 32'hbfc12591} /* (24, 7, 27) {real, imag} */,
  {32'hbfb1e9cb, 32'hbfb5dc84} /* (24, 7, 26) {real, imag} */,
  {32'h3ea8acf0, 32'hc07acdd4} /* (24, 7, 25) {real, imag} */,
  {32'hbe8f666c, 32'hc00fb37e} /* (24, 7, 24) {real, imag} */,
  {32'hc00987c4, 32'hbf960c82} /* (24, 7, 23) {real, imag} */,
  {32'hc043b0c3, 32'hc0071a17} /* (24, 7, 22) {real, imag} */,
  {32'h3f5f81b2, 32'hbf993822} /* (24, 7, 21) {real, imag} */,
  {32'h3f703f54, 32'h3fdf3762} /* (24, 7, 20) {real, imag} */,
  {32'hbe189554, 32'h3f71f348} /* (24, 7, 19) {real, imag} */,
  {32'hbe8e41a4, 32'h4026ac5c} /* (24, 7, 18) {real, imag} */,
  {32'h3fa52e26, 32'h3f87db17} /* (24, 7, 17) {real, imag} */,
  {32'h3fe13c2f, 32'h40237a5a} /* (24, 7, 16) {real, imag} */,
  {32'h3e877432, 32'h402387a4} /* (24, 7, 15) {real, imag} */,
  {32'h403a94e4, 32'h3f8c9748} /* (24, 7, 14) {real, imag} */,
  {32'h4053a9c6, 32'h3f915e89} /* (24, 7, 13) {real, imag} */,
  {32'h403d51b5, 32'h3fc24f26} /* (24, 7, 12) {real, imag} */,
  {32'h4028d191, 32'h3ebcecee} /* (24, 7, 11) {real, imag} */,
  {32'h3df390a0, 32'hbf140fca} /* (24, 7, 10) {real, imag} */,
  {32'hbd92ef80, 32'hbfa5e870} /* (24, 7, 9) {real, imag} */,
  {32'hbe4f3008, 32'hc00c3b5b} /* (24, 7, 8) {real, imag} */,
  {32'hc02b6e83, 32'hbff6d92c} /* (24, 7, 7) {real, imag} */,
  {32'hc06f2e54, 32'hc027707a} /* (24, 7, 6) {real, imag} */,
  {32'hc0177d4c, 32'hc083e535} /* (24, 7, 5) {real, imag} */,
  {32'hc0177bda, 32'hc05950e2} /* (24, 7, 4) {real, imag} */,
  {32'hc01a86f3, 32'hbf968aa2} /* (24, 7, 3) {real, imag} */,
  {32'hc03194a2, 32'hbf9a75f2} /* (24, 7, 2) {real, imag} */,
  {32'hc01c78e8, 32'hc003ea64} /* (24, 7, 1) {real, imag} */,
  {32'hbf9c8944, 32'hbf862350} /* (24, 7, 0) {real, imag} */,
  {32'hbfaff50b, 32'hc0175aa8} /* (24, 6, 31) {real, imag} */,
  {32'hbe7eb44c, 32'hc03772eb} /* (24, 6, 30) {real, imag} */,
  {32'hc00deff0, 32'hbfddfe4b} /* (24, 6, 29) {real, imag} */,
  {32'hbfe8c92a, 32'hc003e238} /* (24, 6, 28) {real, imag} */,
  {32'hbf6a349e, 32'hc010a3f5} /* (24, 6, 27) {real, imag} */,
  {32'hbeb0bbe4, 32'hc0476c22} /* (24, 6, 26) {real, imag} */,
  {32'h3e50c120, 32'hc05fd8e5} /* (24, 6, 25) {real, imag} */,
  {32'hc002d2b0, 32'hbfff40f4} /* (24, 6, 24) {real, imag} */,
  {32'hc010fd56, 32'h3e816524} /* (24, 6, 23) {real, imag} */,
  {32'hc00f0234, 32'hbf836ca3} /* (24, 6, 22) {real, imag} */,
  {32'hbf2e0bce, 32'hc00aac50} /* (24, 6, 21) {real, imag} */,
  {32'h3f5cc01f, 32'h4023c868} /* (24, 6, 20) {real, imag} */,
  {32'h3e34d124, 32'h3fbb37ff} /* (24, 6, 19) {real, imag} */,
  {32'h3fa89d0e, 32'h40189f94} /* (24, 6, 18) {real, imag} */,
  {32'h3fbfe70a, 32'h401a5ef3} /* (24, 6, 17) {real, imag} */,
  {32'h3f138bac, 32'h3fd475d4} /* (24, 6, 16) {real, imag} */,
  {32'h3f51b5db, 32'h3fa1b158} /* (24, 6, 15) {real, imag} */,
  {32'h40060b86, 32'h400b3148} /* (24, 6, 14) {real, imag} */,
  {32'h3f6a4e68, 32'h4037203e} /* (24, 6, 13) {real, imag} */,
  {32'h3f15ef3d, 32'h3fe6daba} /* (24, 6, 12) {real, imag} */,
  {32'h3f7bcea4, 32'h3e8d2ee0} /* (24, 6, 11) {real, imag} */,
  {32'hc018696c, 32'hbf937aa8} /* (24, 6, 10) {real, imag} */,
  {32'hc03d135a, 32'hc05630f0} /* (24, 6, 9) {real, imag} */,
  {32'hbfe1bfc4, 32'hc0828042} /* (24, 6, 8) {real, imag} */,
  {32'hc02f3d4e, 32'hbfec862c} /* (24, 6, 7) {real, imag} */,
  {32'hc051ed30, 32'hbfb187bd} /* (24, 6, 6) {real, imag} */,
  {32'hbff7f187, 32'hbfcbf671} /* (24, 6, 5) {real, imag} */,
  {32'hbff27b9f, 32'hc06cdaee} /* (24, 6, 4) {real, imag} */,
  {32'hbf9f2d34, 32'hc03f1dbc} /* (24, 6, 3) {real, imag} */,
  {32'hbf80f6b0, 32'hbff6c60f} /* (24, 6, 2) {real, imag} */,
  {32'hc045d915, 32'hc01e8f2b} /* (24, 6, 1) {real, imag} */,
  {32'hbfe7b605, 32'hbf5cfca7} /* (24, 6, 0) {real, imag} */,
  {32'h3d0a11a0, 32'hbf0abe2c} /* (24, 5, 31) {real, imag} */,
  {32'hbf4c7f56, 32'hbfa500d8} /* (24, 5, 30) {real, imag} */,
  {32'hc01db64a, 32'hbfccc286} /* (24, 5, 29) {real, imag} */,
  {32'hc030f21e, 32'hc068c3b8} /* (24, 5, 28) {real, imag} */,
  {32'hbff0a988, 32'hc0248105} /* (24, 5, 27) {real, imag} */,
  {32'hbfe325d2, 32'hc01f3b2c} /* (24, 5, 26) {real, imag} */,
  {32'hbd1c81f0, 32'hc04dc922} /* (24, 5, 25) {real, imag} */,
  {32'hbf9acb02, 32'hbf97ef26} /* (24, 5, 24) {real, imag} */,
  {32'hbf94653e, 32'hbefe27ae} /* (24, 5, 23) {real, imag} */,
  {32'hbfa19bca, 32'hbff32dd0} /* (24, 5, 22) {real, imag} */,
  {32'hc04cd078, 32'hc00360b8} /* (24, 5, 21) {real, imag} */,
  {32'hbfb30e06, 32'hbe5b6e98} /* (24, 5, 20) {real, imag} */,
  {32'h3f565680, 32'hbfa79ac4} /* (24, 5, 19) {real, imag} */,
  {32'h400ef0d6, 32'hbe902e36} /* (24, 5, 18) {real, imag} */,
  {32'hbe4745e8, 32'h3fc081be} /* (24, 5, 17) {real, imag} */,
  {32'h3efb8796, 32'h3f8b5d12} /* (24, 5, 16) {real, imag} */,
  {32'h402b174f, 32'h3fb46558} /* (24, 5, 15) {real, imag} */,
  {32'h40633654, 32'h402f75e3} /* (24, 5, 14) {real, imag} */,
  {32'h3fb2615c, 32'h400271ce} /* (24, 5, 13) {real, imag} */,
  {32'h3fb5eb26, 32'h3f26809c} /* (24, 5, 12) {real, imag} */,
  {32'h3f897058, 32'h3e146fb0} /* (24, 5, 11) {real, imag} */,
  {32'hbf8c8aa4, 32'hbf953e88} /* (24, 5, 10) {real, imag} */,
  {32'h3e1e4916, 32'hbff3695a} /* (24, 5, 9) {real, imag} */,
  {32'h3fcf4e8c, 32'hbebdc0bf} /* (24, 5, 8) {real, imag} */,
  {32'h3fa0b0af, 32'h3fc97426} /* (24, 5, 7) {real, imag} */,
  {32'h3e3b2940, 32'h3d2170f4} /* (24, 5, 6) {real, imag} */,
  {32'hbd6c1a20, 32'h3dd5afa0} /* (24, 5, 5) {real, imag} */,
  {32'hbf684f31, 32'hc018d4e8} /* (24, 5, 4) {real, imag} */,
  {32'hbffa1032, 32'hc0176292} /* (24, 5, 3) {real, imag} */,
  {32'hbfd46578, 32'hc0208856} /* (24, 5, 2) {real, imag} */,
  {32'hc02bdd69, 32'hc02006ce} /* (24, 5, 1) {real, imag} */,
  {32'hbefe3a12, 32'hbdb2eae0} /* (24, 5, 0) {real, imag} */,
  {32'h3eae0f00, 32'h3f526000} /* (24, 4, 31) {real, imag} */,
  {32'h3f8f41e0, 32'hbe4a8528} /* (24, 4, 30) {real, imag} */,
  {32'hbf4fdcd0, 32'hbdf93cb0} /* (24, 4, 29) {real, imag} */,
  {32'hc0632608, 32'hbfd59451} /* (24, 4, 28) {real, imag} */,
  {32'hbf5205ea, 32'hbf894189} /* (24, 4, 27) {real, imag} */,
  {32'hbfe5f033, 32'hbee1a866} /* (24, 4, 26) {real, imag} */,
  {32'hbfcce55c, 32'hbfcf07d1} /* (24, 4, 25) {real, imag} */,
  {32'hc0222063, 32'hbfcfeef3} /* (24, 4, 24) {real, imag} */,
  {32'hbf7671f1, 32'hbfa020df} /* (24, 4, 23) {real, imag} */,
  {32'hbff65d0e, 32'hbf8d3cd9} /* (24, 4, 22) {real, imag} */,
  {32'hc03aa674, 32'hbfbffc78} /* (24, 4, 21) {real, imag} */,
  {32'hc0519392, 32'hbf9f4242} /* (24, 4, 20) {real, imag} */,
  {32'hbf9cf1c6, 32'hc00a9791} /* (24, 4, 19) {real, imag} */,
  {32'hbee49210, 32'hc01351e2} /* (24, 4, 18) {real, imag} */,
  {32'hbf8c7203, 32'hc04dad4c} /* (24, 4, 17) {real, imag} */,
  {32'hbf488cdd, 32'hc03a69b2} /* (24, 4, 16) {real, imag} */,
  {32'h400700e2, 32'hbd0d1d00} /* (24, 4, 15) {real, imag} */,
  {32'h40846746, 32'h3f800cd3} /* (24, 4, 14) {real, imag} */,
  {32'h4017bb2c, 32'h3ebec31c} /* (24, 4, 13) {real, imag} */,
  {32'h3fa3e270, 32'hbfa001d4} /* (24, 4, 12) {real, imag} */,
  {32'h3f29a758, 32'h3f6477af} /* (24, 4, 11) {real, imag} */,
  {32'h3e587bb8, 32'hbe563e78} /* (24, 4, 10) {real, imag} */,
  {32'h4005e1c9, 32'h3ee56be4} /* (24, 4, 9) {real, imag} */,
  {32'h4058895b, 32'h401dd169} /* (24, 4, 8) {real, imag} */,
  {32'h40262b84, 32'h40200932} /* (24, 4, 7) {real, imag} */,
  {32'h3fcca50e, 32'h3ebfc7cc} /* (24, 4, 6) {real, imag} */,
  {32'hbf1c86cf, 32'hbf201f34} /* (24, 4, 5) {real, imag} */,
  {32'hc004ecb0, 32'hbfb50104} /* (24, 4, 4) {real, imag} */,
  {32'hc03b9b54, 32'hc04157fd} /* (24, 4, 3) {real, imag} */,
  {32'hc0431a20, 32'hc0271f8c} /* (24, 4, 2) {real, imag} */,
  {32'hc04d0d32, 32'hc00228f2} /* (24, 4, 1) {real, imag} */,
  {32'hbfdcbcc7, 32'hbebee4ee} /* (24, 4, 0) {real, imag} */,
  {32'hbf816eac, 32'hbf3485a4} /* (24, 3, 31) {real, imag} */,
  {32'hbe448f4c, 32'hc01cd738} /* (24, 3, 30) {real, imag} */,
  {32'hbdcc3d00, 32'hc0261ec0} /* (24, 3, 29) {real, imag} */,
  {32'hc021aa7e, 32'hc0697d90} /* (24, 3, 28) {real, imag} */,
  {32'hbf65f7dc, 32'hc03239aa} /* (24, 3, 27) {real, imag} */,
  {32'hbfa3f9ec, 32'hbf91c07a} /* (24, 3, 26) {real, imag} */,
  {32'hbfdceb5c, 32'hbf01309e} /* (24, 3, 25) {real, imag} */,
  {32'hc07620a0, 32'hbfdfb38b} /* (24, 3, 24) {real, imag} */,
  {32'hbf094c81, 32'hc0170c94} /* (24, 3, 23) {real, imag} */,
  {32'hc02e3220, 32'hbfc24ea5} /* (24, 3, 22) {real, imag} */,
  {32'hc0691798, 32'hc02333c3} /* (24, 3, 21) {real, imag} */,
  {32'hc0481fdb, 32'hbfa2d9d6} /* (24, 3, 20) {real, imag} */,
  {32'hc00a9982, 32'hc02801c4} /* (24, 3, 19) {real, imag} */,
  {32'hc0768ca2, 32'hc0452ed4} /* (24, 3, 18) {real, imag} */,
  {32'hc01f30fc, 32'hc03c983b} /* (24, 3, 17) {real, imag} */,
  {32'hbf2ceed6, 32'hc0036265} /* (24, 3, 16) {real, imag} */,
  {32'h3fc79254, 32'h400d6c13} /* (24, 3, 15) {real, imag} */,
  {32'h40413332, 32'h3ff758bf} /* (24, 3, 14) {real, imag} */,
  {32'h401d10d6, 32'h403b13a5} /* (24, 3, 13) {real, imag} */,
  {32'h40061982, 32'h3ed9eb50} /* (24, 3, 12) {real, imag} */,
  {32'h3fbe0145, 32'h3eb40542} /* (24, 3, 11) {real, imag} */,
  {32'h3faa4921, 32'h3f843f64} /* (24, 3, 10) {real, imag} */,
  {32'h3fd66e41, 32'h3f416bc4} /* (24, 3, 9) {real, imag} */,
  {32'h401ad6cc, 32'h3fe42d44} /* (24, 3, 8) {real, imag} */,
  {32'h3ff3ff1b, 32'h4027514c} /* (24, 3, 7) {real, imag} */,
  {32'h3f24c7fa, 32'h3f57197f} /* (24, 3, 6) {real, imag} */,
  {32'h3e5631fa, 32'hbfde5e86} /* (24, 3, 5) {real, imag} */,
  {32'hbf934e2a, 32'hc0039cda} /* (24, 3, 4) {real, imag} */,
  {32'hbfcdd4da, 32'hc065754a} /* (24, 3, 3) {real, imag} */,
  {32'hbff31b5e, 32'hc03d4d01} /* (24, 3, 2) {real, imag} */,
  {32'hbfd148d5, 32'hc0039fc1} /* (24, 3, 1) {real, imag} */,
  {32'hbfe7b66d, 32'hbeba50e4} /* (24, 3, 0) {real, imag} */,
  {32'hbec07f68, 32'hbe72fbf4} /* (24, 2, 31) {real, imag} */,
  {32'hbf6858a5, 32'hbfeda0ce} /* (24, 2, 30) {real, imag} */,
  {32'hbd9a4248, 32'hc00b249a} /* (24, 2, 29) {real, imag} */,
  {32'hc01ac10a, 32'hc069fe3b} /* (24, 2, 28) {real, imag} */,
  {32'hc01ed8d0, 32'hc01e17a0} /* (24, 2, 27) {real, imag} */,
  {32'hc009ae5c, 32'hbf53e40e} /* (24, 2, 26) {real, imag} */,
  {32'hbf3991b9, 32'h3e54f2a2} /* (24, 2, 25) {real, imag} */,
  {32'hbf35348c, 32'h3dc86650} /* (24, 2, 24) {real, imag} */,
  {32'h3f57f39c, 32'hbfab3a95} /* (24, 2, 23) {real, imag} */,
  {32'hc0131bcb, 32'hbe2585fc} /* (24, 2, 22) {real, imag} */,
  {32'hc0670370, 32'hc0478fad} /* (24, 2, 21) {real, imag} */,
  {32'hbf79f4a4, 32'hc01b4cb6} /* (24, 2, 20) {real, imag} */,
  {32'hbfa7ac31, 32'hc00c6ec0} /* (24, 2, 19) {real, imag} */,
  {32'hc04770cb, 32'hc03dd3b4} /* (24, 2, 18) {real, imag} */,
  {32'hc05abda5, 32'hbfd25ac7} /* (24, 2, 17) {real, imag} */,
  {32'hbc27d600, 32'h3e4ff738} /* (24, 2, 16) {real, imag} */,
  {32'h3ff05c26, 32'h4086faa7} /* (24, 2, 15) {real, imag} */,
  {32'h3f63e449, 32'h403e453e} /* (24, 2, 14) {real, imag} */,
  {32'h3f7c3904, 32'h408efd4f} /* (24, 2, 13) {real, imag} */,
  {32'h407591a6, 32'h4075c2a9} /* (24, 2, 12) {real, imag} */,
  {32'h40584641, 32'h4045e47a} /* (24, 2, 11) {real, imag} */,
  {32'h3fe60f87, 32'h3ff1d5ef} /* (24, 2, 10) {real, imag} */,
  {32'hbf020194, 32'h3fc64d94} /* (24, 2, 9) {real, imag} */,
  {32'h3f2a70a1, 32'h40028d2e} /* (24, 2, 8) {real, imag} */,
  {32'h4002b65b, 32'h3ff3fc4c} /* (24, 2, 7) {real, imag} */,
  {32'h3ff408c8, 32'h3ffefe3a} /* (24, 2, 6) {real, imag} */,
  {32'h404b7fcc, 32'hbe95d24f} /* (24, 2, 5) {real, imag} */,
  {32'h3f5b8353, 32'hc06308ab} /* (24, 2, 4) {real, imag} */,
  {32'hc0011e86, 32'hc0608bb9} /* (24, 2, 3) {real, imag} */,
  {32'hbf0b2d24, 32'hc0435087} /* (24, 2, 2) {real, imag} */,
  {32'h3ff061c8, 32'hc07a799e} /* (24, 2, 1) {real, imag} */,
  {32'hbdbd6834, 32'hc004aaca} /* (24, 2, 0) {real, imag} */,
  {32'h3fca2a1c, 32'hbf5db2e5} /* (24, 1, 31) {real, imag} */,
  {32'hbf12c9fc, 32'hc0194de2} /* (24, 1, 30) {real, imag} */,
  {32'hc016bccb, 32'hbfb09c1f} /* (24, 1, 29) {real, imag} */,
  {32'hc095f85c, 32'hc00dbaa2} /* (24, 1, 28) {real, imag} */,
  {32'hc082c7f6, 32'hc014fda8} /* (24, 1, 27) {real, imag} */,
  {32'hbfa68913, 32'hbfee4244} /* (24, 1, 26) {real, imag} */,
  {32'hbe9097d8, 32'hbfc52690} /* (24, 1, 25) {real, imag} */,
  {32'hbe5925a8, 32'hbf1d72de} /* (24, 1, 24) {real, imag} */,
  {32'h3f91ed2e, 32'hc01d676a} /* (24, 1, 23) {real, imag} */,
  {32'hbf94e9a7, 32'hc029a8c4} /* (24, 1, 22) {real, imag} */,
  {32'hbfd0e044, 32'hc0407348} /* (24, 1, 21) {real, imag} */,
  {32'h3e4587ec, 32'hc0370448} /* (24, 1, 20) {real, imag} */,
  {32'hbf18246e, 32'hc0477676} /* (24, 1, 19) {real, imag} */,
  {32'hbf88d695, 32'hc082e22e} /* (24, 1, 18) {real, imag} */,
  {32'hbfd14bc4, 32'hbfb97bb8} /* (24, 1, 17) {real, imag} */,
  {32'h3faf407e, 32'hbe6147c0} /* (24, 1, 16) {real, imag} */,
  {32'h40024234, 32'h4027f180} /* (24, 1, 15) {real, imag} */,
  {32'h3e0f1bd0, 32'h40635072} /* (24, 1, 14) {real, imag} */,
  {32'h3f9c2e3e, 32'h3fa86206} /* (24, 1, 13) {real, imag} */,
  {32'h40084a76, 32'h3fdd2060} /* (24, 1, 12) {real, imag} */,
  {32'h40714cde, 32'h402acbfd} /* (24, 1, 11) {real, imag} */,
  {32'h4045adfb, 32'h40427c67} /* (24, 1, 10) {real, imag} */,
  {32'h3f08aab1, 32'h4009e869} /* (24, 1, 9) {real, imag} */,
  {32'h3f9ff604, 32'h40107666} /* (24, 1, 8) {real, imag} */,
  {32'h40109026, 32'h3e953226} /* (24, 1, 7) {real, imag} */,
  {32'h4032f410, 32'hbe14cf18} /* (24, 1, 6) {real, imag} */,
  {32'hbe1668b6, 32'hbe9b3fec} /* (24, 1, 5) {real, imag} */,
  {32'hbfed39f6, 32'hc0430626} /* (24, 1, 4) {real, imag} */,
  {32'hc00b5bf7, 32'hbff2e35c} /* (24, 1, 3) {real, imag} */,
  {32'h3f26437c, 32'hbffb601d} /* (24, 1, 2) {real, imag} */,
  {32'h401eaa64, 32'hbfd4be5c} /* (24, 1, 1) {real, imag} */,
  {32'h3fb71b68, 32'hbf880617} /* (24, 1, 0) {real, imag} */,
  {32'h3d8f6c84, 32'hbe98a277} /* (24, 0, 31) {real, imag} */,
  {32'hbf8b63d6, 32'hbe0c79a6} /* (24, 0, 30) {real, imag} */,
  {32'hc02514bf, 32'h3e209f2e} /* (24, 0, 29) {real, imag} */,
  {32'hc0690db2, 32'hbf4015c0} /* (24, 0, 28) {real, imag} */,
  {32'hc072fd0c, 32'hbff106ae} /* (24, 0, 27) {real, imag} */,
  {32'hbf74348e, 32'hbfd4f560} /* (24, 0, 26) {real, imag} */,
  {32'hbf1bf4e5, 32'hbf224366} /* (24, 0, 25) {real, imag} */,
  {32'hbe7c37a0, 32'h3f5b9d5c} /* (24, 0, 24) {real, imag} */,
  {32'h3dbe8808, 32'hbff7aa26} /* (24, 0, 23) {real, imag} */,
  {32'hbf29548a, 32'hc03f9f0b} /* (24, 0, 22) {real, imag} */,
  {32'hbf1d04ed, 32'hbf648ce6} /* (24, 0, 21) {real, imag} */,
  {32'h3d7b6b20, 32'hbee14873} /* (24, 0, 20) {real, imag} */,
  {32'hbda93d40, 32'hbfdb2e6a} /* (24, 0, 19) {real, imag} */,
  {32'hbead3ab0, 32'hbff0c93e} /* (24, 0, 18) {real, imag} */,
  {32'hbed222d4, 32'hbf3d953e} /* (24, 0, 17) {real, imag} */,
  {32'h3f6539bc, 32'hbf349962} /* (24, 0, 16) {real, imag} */,
  {32'h3f4f84d8, 32'h3f359b88} /* (24, 0, 15) {real, imag} */,
  {32'h3f7225e6, 32'h4010dbe6} /* (24, 0, 14) {real, imag} */,
  {32'h400ce0a2, 32'h3f40171b} /* (24, 0, 13) {real, imag} */,
  {32'h3f2b14ee, 32'h3fab367a} /* (24, 0, 12) {real, imag} */,
  {32'h3fa75646, 32'h3ff2a6ce} /* (24, 0, 11) {real, imag} */,
  {32'h3f64ec04, 32'h3faa04c6} /* (24, 0, 10) {real, imag} */,
  {32'h3f39ad56, 32'hbf04b7aa} /* (24, 0, 9) {real, imag} */,
  {32'h3fcabc94, 32'hbdd4f8f8} /* (24, 0, 8) {real, imag} */,
  {32'h4011c5bb, 32'hbf39e498} /* (24, 0, 7) {real, imag} */,
  {32'h3f9c02ea, 32'hbfd5c74a} /* (24, 0, 6) {real, imag} */,
  {32'hbfb7f67e, 32'hbf0dc23c} /* (24, 0, 5) {real, imag} */,
  {32'hbffc3fba, 32'hbf85b6d5} /* (24, 0, 4) {real, imag} */,
  {32'hbf9ae831, 32'hbf31b52e} /* (24, 0, 3) {real, imag} */,
  {32'h3f5639ce, 32'hc0013f58} /* (24, 0, 2) {real, imag} */,
  {32'h3fa4e7f8, 32'hbf464a7e} /* (24, 0, 1) {real, imag} */,
  {32'hbb4a6b00, 32'h3e8a287c} /* (24, 0, 0) {real, imag} */,
  {32'hbe7092c4, 32'hbf6a6604} /* (23, 31, 31) {real, imag} */,
  {32'hbe5fd6b8, 32'hbf4702fa} /* (23, 31, 30) {real, imag} */,
  {32'hbfa39d41, 32'h3e6e1240} /* (23, 31, 29) {real, imag} */,
  {32'hbfbd719b, 32'hbf2150a0} /* (23, 31, 28) {real, imag} */,
  {32'hbf142c60, 32'hbde10f28} /* (23, 31, 27) {real, imag} */,
  {32'hbf110686, 32'hbfbd8744} /* (23, 31, 26) {real, imag} */,
  {32'hbfdf8496, 32'hbf8de650} /* (23, 31, 25) {real, imag} */,
  {32'hbf40c672, 32'hbf922778} /* (23, 31, 24) {real, imag} */,
  {32'h3f3e6a90, 32'hbf4a340d} /* (23, 31, 23) {real, imag} */,
  {32'h3f90e59f, 32'hbe33412a} /* (23, 31, 22) {real, imag} */,
  {32'hbe8d4c0e, 32'hbe86ba05} /* (23, 31, 21) {real, imag} */,
  {32'hbe044f48, 32'hbec631f4} /* (23, 31, 20) {real, imag} */,
  {32'h3f842e11, 32'hbe4cf80c} /* (23, 31, 19) {real, imag} */,
  {32'hbd4ee2b8, 32'h3f7e1a4a} /* (23, 31, 18) {real, imag} */,
  {32'hbf88859c, 32'hbde63fd4} /* (23, 31, 17) {real, imag} */,
  {32'hbf87c6b9, 32'hbeacefbf} /* (23, 31, 16) {real, imag} */,
  {32'hbe6f663d, 32'h3f0586c2} /* (23, 31, 15) {real, imag} */,
  {32'h3ffae518, 32'hbe7a763f} /* (23, 31, 14) {real, imag} */,
  {32'h402efd1a, 32'h3ece33ac} /* (23, 31, 13) {real, imag} */,
  {32'hbe133f88, 32'h3f1d9482} /* (23, 31, 12) {real, imag} */,
  {32'hbf494d9d, 32'hbe956d22} /* (23, 31, 11) {real, imag} */,
  {32'h3de3d142, 32'h3f789394} /* (23, 31, 10) {real, imag} */,
  {32'hbdbb6ea8, 32'hbe99585f} /* (23, 31, 9) {real, imag} */,
  {32'hbe7c5ac4, 32'hbf3fc72a} /* (23, 31, 8) {real, imag} */,
  {32'h3f14e32c, 32'h3eab773c} /* (23, 31, 7) {real, imag} */,
  {32'h3e82dfd4, 32'h3f80c95f} /* (23, 31, 6) {real, imag} */,
  {32'h3e31ce08, 32'h3d6f6740} /* (23, 31, 5) {real, imag} */,
  {32'h3ecb4805, 32'hbec2c3ca} /* (23, 31, 4) {real, imag} */,
  {32'h3eaec606, 32'h3f38562f} /* (23, 31, 3) {real, imag} */,
  {32'h3ecd62c0, 32'h3fa1a424} /* (23, 31, 2) {real, imag} */,
  {32'hbdc2c0c8, 32'hbd8ccc60} /* (23, 31, 1) {real, imag} */,
  {32'hbdf32578, 32'hbe264500} /* (23, 31, 0) {real, imag} */,
  {32'hc000638a, 32'hbf274a96} /* (23, 30, 31) {real, imag} */,
  {32'hc010bc27, 32'hbe2b3300} /* (23, 30, 30) {real, imag} */,
  {32'hc0150320, 32'hbf8dfe70} /* (23, 30, 29) {real, imag} */,
  {32'hbf7381d3, 32'hbf2605ee} /* (23, 30, 28) {real, imag} */,
  {32'hbf2e3744, 32'h3e850e55} /* (23, 30, 27) {real, imag} */,
  {32'hbf059d62, 32'hc03415b0} /* (23, 30, 26) {real, imag} */,
  {32'hbfb09127, 32'hbfd6d360} /* (23, 30, 25) {real, imag} */,
  {32'hbfa7c3e5, 32'hbfbefa79} /* (23, 30, 24) {real, imag} */,
  {32'hbeb90205, 32'hbfa98ba4} /* (23, 30, 23) {real, imag} */,
  {32'hbf0fd620, 32'hbdbe3888} /* (23, 30, 22) {real, imag} */,
  {32'hbfa37c2a, 32'h3f828d1c} /* (23, 30, 21) {real, imag} */,
  {32'hbf0dc5bb, 32'h3f9e15f0} /* (23, 30, 20) {real, imag} */,
  {32'h3f68006c, 32'hbebd8876} /* (23, 30, 19) {real, imag} */,
  {32'hbf91c4ec, 32'h3f5100d1} /* (23, 30, 18) {real, imag} */,
  {32'hc023a514, 32'h3f07cf0a} /* (23, 30, 17) {real, imag} */,
  {32'hbfa8bc75, 32'h3f39bc2a} /* (23, 30, 16) {real, imag} */,
  {32'h3e821a94, 32'h40114e4c} /* (23, 30, 15) {real, imag} */,
  {32'h3ffa4f49, 32'h4003d32c} /* (23, 30, 14) {real, imag} */,
  {32'h4082cd22, 32'h3f9e6541} /* (23, 30, 13) {real, imag} */,
  {32'h3fa6df40, 32'h3e62eef0} /* (23, 30, 12) {real, imag} */,
  {32'hbf38ef5b, 32'h3eef8fc0} /* (23, 30, 11) {real, imag} */,
  {32'hbf46b2b5, 32'h4004df88} /* (23, 30, 10) {real, imag} */,
  {32'h3cfaab80, 32'hbf1ce2c0} /* (23, 30, 9) {real, imag} */,
  {32'hbdf67358, 32'hbf89155a} /* (23, 30, 8) {real, imag} */,
  {32'hbf010538, 32'hbefab2d0} /* (23, 30, 7) {real, imag} */,
  {32'h3bc2ad00, 32'h3fb9097c} /* (23, 30, 6) {real, imag} */,
  {32'h3e7bda58, 32'h3f75bfe3} /* (23, 30, 5) {real, imag} */,
  {32'h3ec5bce0, 32'hbf03c940} /* (23, 30, 4) {real, imag} */,
  {32'hbee1fbf2, 32'h3eb851aa} /* (23, 30, 3) {real, imag} */,
  {32'h3ec69da4, 32'h3fc09181} /* (23, 30, 2) {real, imag} */,
  {32'hbf517785, 32'h3f16c33e} /* (23, 30, 1) {real, imag} */,
  {32'hbf701ffa, 32'hbe1c4158} /* (23, 30, 0) {real, imag} */,
  {32'hc00ff6df, 32'h3f963fc8} /* (23, 29, 31) {real, imag} */,
  {32'hc0841a06, 32'h3fcd5444} /* (23, 29, 30) {real, imag} */,
  {32'hc00de1da, 32'hbfd8a175} /* (23, 29, 29) {real, imag} */,
  {32'h3bc20d80, 32'hbe1188a8} /* (23, 29, 28) {real, imag} */,
  {32'hbef7fafc, 32'h3f452bae} /* (23, 29, 27) {real, imag} */,
  {32'h3e30d530, 32'hbfdc0a16} /* (23, 29, 26) {real, imag} */,
  {32'hbf5ddab2, 32'hbf36ff7a} /* (23, 29, 25) {real, imag} */,
  {32'hbfb1a325, 32'hbd949ae0} /* (23, 29, 24) {real, imag} */,
  {32'hbf56620c, 32'hbf546df4} /* (23, 29, 23) {real, imag} */,
  {32'hbfe9dd49, 32'hbe971218} /* (23, 29, 22) {real, imag} */,
  {32'hc035c9e4, 32'h3f0c1258} /* (23, 29, 21) {real, imag} */,
  {32'hbfd327b8, 32'h3f2aeef4} /* (23, 29, 20) {real, imag} */,
  {32'h3eaea4d8, 32'h3e9544dc} /* (23, 29, 19) {real, imag} */,
  {32'hbebd2134, 32'h3e4dbaec} /* (23, 29, 18) {real, imag} */,
  {32'hbf4a3535, 32'h3f0bbc59} /* (23, 29, 17) {real, imag} */,
  {32'h3fb7a025, 32'h3f0f3db4} /* (23, 29, 16) {real, imag} */,
  {32'h3fa67c64, 32'h3fbeee2c} /* (23, 29, 15) {real, imag} */,
  {32'hbc3a0200, 32'h3f80acda} /* (23, 29, 14) {real, imag} */,
  {32'h3f83f574, 32'hbf15f02a} /* (23, 29, 13) {real, imag} */,
  {32'h3fd1d833, 32'hbf820b72} /* (23, 29, 12) {real, imag} */,
  {32'h3f926043, 32'hbea7090e} /* (23, 29, 11) {real, imag} */,
  {32'hbf3a3632, 32'hbf39515c} /* (23, 29, 10) {real, imag} */,
  {32'hbf77b6f4, 32'hbfd7275a} /* (23, 29, 9) {real, imag} */,
  {32'hbfac0ab8, 32'hbfaf1e20} /* (23, 29, 8) {real, imag} */,
  {32'hbf938a5d, 32'hbf893902} /* (23, 29, 7) {real, imag} */,
  {32'h3f183722, 32'hbf4c5dd0} /* (23, 29, 6) {real, imag} */,
  {32'hbd4bae40, 32'hbfcb9db6} /* (23, 29, 5) {real, imag} */,
  {32'hbf6e3dfd, 32'hc018cb0e} /* (23, 29, 4) {real, imag} */,
  {32'hbfe4dc36, 32'hbf1bdad0} /* (23, 29, 3) {real, imag} */,
  {32'h3f21a174, 32'hbf0b7d34} /* (23, 29, 2) {real, imag} */,
  {32'h3e3ee79c, 32'hbfdc7b2e} /* (23, 29, 1) {real, imag} */,
  {32'hbe250e0c, 32'hbe90babe} /* (23, 29, 0) {real, imag} */,
  {32'hbf18d1e2, 32'h3f5b6938} /* (23, 28, 31) {real, imag} */,
  {32'hc03d35fe, 32'h3f7c415a} /* (23, 28, 30) {real, imag} */,
  {32'hc0024bb9, 32'hbfc1d88c} /* (23, 28, 29) {real, imag} */,
  {32'hbe4d4f5a, 32'hbf59fd32} /* (23, 28, 28) {real, imag} */,
  {32'hbfa90712, 32'h3ed8f160} /* (23, 28, 27) {real, imag} */,
  {32'hbe2b8ebf, 32'hbeb7b6c8} /* (23, 28, 26) {real, imag} */,
  {32'hbf5366fa, 32'hbf9de8f9} /* (23, 28, 25) {real, imag} */,
  {32'hbf9d6bcc, 32'hc00dafbd} /* (23, 28, 24) {real, imag} */,
  {32'hbf17bc56, 32'h3e1f9bc8} /* (23, 28, 23) {real, imag} */,
  {32'hbf11529b, 32'h3f26f6ec} /* (23, 28, 22) {real, imag} */,
  {32'hbfc34192, 32'h3fbc84e8} /* (23, 28, 21) {real, imag} */,
  {32'h3d27bf90, 32'h40041b40} /* (23, 28, 20) {real, imag} */,
  {32'h3ffd3ad2, 32'h3fbd1cce} /* (23, 28, 19) {real, imag} */,
  {32'h3fae1c98, 32'h3f8aff53} /* (23, 28, 18) {real, imag} */,
  {32'h3ec43730, 32'h3e4807fe} /* (23, 28, 17) {real, imag} */,
  {32'h3f1e4ce2, 32'hbbd60c00} /* (23, 28, 16) {real, imag} */,
  {32'h3f5b3e88, 32'h3df26748} /* (23, 28, 15) {real, imag} */,
  {32'hbe397430, 32'h3e5949f0} /* (23, 28, 14) {real, imag} */,
  {32'hbc8f3ee0, 32'hbf58e8a6} /* (23, 28, 13) {real, imag} */,
  {32'h3fd71f73, 32'hbea643ba} /* (23, 28, 12) {real, imag} */,
  {32'h3fd99a0c, 32'h3e674a2c} /* (23, 28, 11) {real, imag} */,
  {32'hbff80dd0, 32'hbf621ba0} /* (23, 28, 10) {real, imag} */,
  {32'hbf84aac3, 32'hbfccc1d2} /* (23, 28, 9) {real, imag} */,
  {32'hbdd58cb4, 32'hbb9e2000} /* (23, 28, 8) {real, imag} */,
  {32'h3f3a9433, 32'hbe93a19c} /* (23, 28, 7) {real, imag} */,
  {32'hbf4bc91e, 32'hbf8deb55} /* (23, 28, 6) {real, imag} */,
  {32'hc020c2ce, 32'hc036e358} /* (23, 28, 5) {real, imag} */,
  {32'hbf90a9a5, 32'hbf7e64ef} /* (23, 28, 4) {real, imag} */,
  {32'hbf13d80f, 32'hbf9c5c2b} /* (23, 28, 3) {real, imag} */,
  {32'hbdf12a88, 32'hbf9adb10} /* (23, 28, 2) {real, imag} */,
  {32'hbfb33380, 32'hbf46dbf6} /* (23, 28, 1) {real, imag} */,
  {32'hbfba2c36, 32'h3eb6a63c} /* (23, 28, 0) {real, imag} */,
  {32'hbea77dbe, 32'h3f80c0c2} /* (23, 27, 31) {real, imag} */,
  {32'hbe8525a0, 32'hbde5af30} /* (23, 27, 30) {real, imag} */,
  {32'h3e06fc24, 32'hc0182332} /* (23, 27, 29) {real, imag} */,
  {32'hbe6889d4, 32'hc00fed79} /* (23, 27, 28) {real, imag} */,
  {32'hbfbed93b, 32'hbf98315f} /* (23, 27, 27) {real, imag} */,
  {32'hc0131271, 32'h3f40bf9b} /* (23, 27, 26) {real, imag} */,
  {32'hc0144376, 32'hbf71f308} /* (23, 27, 25) {real, imag} */,
  {32'h3d124750, 32'hbffed9fd} /* (23, 27, 24) {real, imag} */,
  {32'hbe3bf222, 32'h3fb8c161} /* (23, 27, 23) {real, imag} */,
  {32'hbfa7e78a, 32'hbd620a00} /* (23, 27, 22) {real, imag} */,
  {32'hbf93c107, 32'h3fb3e421} /* (23, 27, 21) {real, imag} */,
  {32'hbec8659c, 32'h40159d6d} /* (23, 27, 20) {real, imag} */,
  {32'h3e997df8, 32'hbd908e60} /* (23, 27, 19) {real, imag} */,
  {32'h4012771a, 32'h3e6a476c} /* (23, 27, 18) {real, imag} */,
  {32'h3fc4af6f, 32'h3c5a9c80} /* (23, 27, 17) {real, imag} */,
  {32'hbe45c550, 32'h3f612e90} /* (23, 27, 16) {real, imag} */,
  {32'h3fd1cf88, 32'h3ea2547c} /* (23, 27, 15) {real, imag} */,
  {32'h3ee3be7c, 32'hbde610a0} /* (23, 27, 14) {real, imag} */,
  {32'h3f0dd752, 32'hbe1a4dd4} /* (23, 27, 13) {real, imag} */,
  {32'h3f531672, 32'h3eb45d06} /* (23, 27, 12) {real, imag} */,
  {32'hbe376dac, 32'h3fb6758b} /* (23, 27, 11) {real, imag} */,
  {32'hbfff42c0, 32'h3f9123f8} /* (23, 27, 10) {real, imag} */,
  {32'hbfadf66b, 32'hbf813a20} /* (23, 27, 9) {real, imag} */,
  {32'hbfb595ca, 32'hbe9a55c4} /* (23, 27, 8) {real, imag} */,
  {32'h3ee701ec, 32'h3e06af38} /* (23, 27, 7) {real, imag} */,
  {32'hbf7fcb3b, 32'h3ed5ba44} /* (23, 27, 6) {real, imag} */,
  {32'hbfe359e2, 32'hbfb8f8f2} /* (23, 27, 5) {real, imag} */,
  {32'hbf822043, 32'hbc527900} /* (23, 27, 4) {real, imag} */,
  {32'hbef6fa96, 32'h3cedf820} /* (23, 27, 3) {real, imag} */,
  {32'hbe269b40, 32'h3ec57c91} /* (23, 27, 2) {real, imag} */,
  {32'hc03eecd4, 32'h3e133d24} /* (23, 27, 1) {real, imag} */,
  {32'hbfe175f1, 32'hbe1fb280} /* (23, 27, 0) {real, imag} */,
  {32'hbf5b144b, 32'hbe8cd704} /* (23, 26, 31) {real, imag} */,
  {32'hbfe11ed1, 32'hbeca42ba} /* (23, 26, 30) {real, imag} */,
  {32'hbf3de09d, 32'hbfed3f4c} /* (23, 26, 29) {real, imag} */,
  {32'h3fc75b38, 32'hbf710bac} /* (23, 26, 28) {real, imag} */,
  {32'h3ee6e7f2, 32'h3de557b0} /* (23, 26, 27) {real, imag} */,
  {32'hc0195010, 32'hbe12d6ac} /* (23, 26, 26) {real, imag} */,
  {32'hc018a612, 32'hbf881330} /* (23, 26, 25) {real, imag} */,
  {32'hbf8c6f10, 32'hbfb63390} /* (23, 26, 24) {real, imag} */,
  {32'hbeb68d90, 32'h3e1ef3ae} /* (23, 26, 23) {real, imag} */,
  {32'hbf203116, 32'hbff10e0c} /* (23, 26, 22) {real, imag} */,
  {32'hbfa77294, 32'hbfcc41ed} /* (23, 26, 21) {real, imag} */,
  {32'hbf08acb6, 32'hbf7a68a3} /* (23, 26, 20) {real, imag} */,
  {32'h3f9f1288, 32'hbf1b54b8} /* (23, 26, 19) {real, imag} */,
  {32'h3fcc5d0b, 32'h3f7880d4} /* (23, 26, 18) {real, imag} */,
  {32'h3ea3afb7, 32'h3f023a2f} /* (23, 26, 17) {real, imag} */,
  {32'h3e33b438, 32'h3f43bd99} /* (23, 26, 16) {real, imag} */,
  {32'h3f9f85ce, 32'hbeaacc88} /* (23, 26, 15) {real, imag} */,
  {32'h3f10b342, 32'hbfe4e9cf} /* (23, 26, 14) {real, imag} */,
  {32'h3f1c8703, 32'hbd809fa0} /* (23, 26, 13) {real, imag} */,
  {32'h3f3e812c, 32'h3ed5d966} /* (23, 26, 12) {real, imag} */,
  {32'h3f757c72, 32'h3f1a04d2} /* (23, 26, 11) {real, imag} */,
  {32'hbf656f5b, 32'h3f7b0796} /* (23, 26, 10) {real, imag} */,
  {32'hc0415f8b, 32'hbfd93efe} /* (23, 26, 9) {real, imag} */,
  {32'hc0196320, 32'hbfd5d550} /* (23, 26, 8) {real, imag} */,
  {32'hbed87440, 32'hbdbae168} /* (23, 26, 7) {real, imag} */,
  {32'hbf81f60c, 32'hbebc5e3a} /* (23, 26, 6) {real, imag} */,
  {32'hc011b4b2, 32'hbf9c7f4c} /* (23, 26, 5) {real, imag} */,
  {32'hbfd409f7, 32'h3e5963c0} /* (23, 26, 4) {real, imag} */,
  {32'hbf83d48c, 32'h3f82c30a} /* (23, 26, 3) {real, imag} */,
  {32'hbf985573, 32'hbe869440} /* (23, 26, 2) {real, imag} */,
  {32'hbfe95bdf, 32'hbfc7d06c} /* (23, 26, 1) {real, imag} */,
  {32'h3e9e3bb8, 32'hbeb415f3} /* (23, 26, 0) {real, imag} */,
  {32'hbe3cf7c2, 32'hbfce30f4} /* (23, 25, 31) {real, imag} */,
  {32'hbf933863, 32'hbfaeba12} /* (23, 25, 30) {real, imag} */,
  {32'hbfd18d76, 32'hbebe0ce4} /* (23, 25, 29) {real, imag} */,
  {32'hbe735b9c, 32'h3fc61194} /* (23, 25, 28) {real, imag} */,
  {32'hbf3501a0, 32'h3f1531d7} /* (23, 25, 27) {real, imag} */,
  {32'hc00d46ec, 32'hbfa6129b} /* (23, 25, 26) {real, imag} */,
  {32'h3c560400, 32'hbf8afe26} /* (23, 25, 25) {real, imag} */,
  {32'hbc9e20e0, 32'hc00214f6} /* (23, 25, 24) {real, imag} */,
  {32'h3f9811b2, 32'hc01bb173} /* (23, 25, 23) {real, imag} */,
  {32'h3fc5bf81, 32'hc02e53ee} /* (23, 25, 22) {real, imag} */,
  {32'hbea4cc96, 32'hc01a2c8a} /* (23, 25, 21) {real, imag} */,
  {32'h3fbd5ab4, 32'h3de57110} /* (23, 25, 20) {real, imag} */,
  {32'h3feb9952, 32'h3f8125ce} /* (23, 25, 19) {real, imag} */,
  {32'h3f3cca70, 32'h3dbd97b0} /* (23, 25, 18) {real, imag} */,
  {32'hbe847d28, 32'h3ee2b51c} /* (23, 25, 17) {real, imag} */,
  {32'h3f894d80, 32'h3ec5e7b0} /* (23, 25, 16) {real, imag} */,
  {32'h3f84f6aa, 32'hbf1dc7b6} /* (23, 25, 15) {real, imag} */,
  {32'h3e1ceb3c, 32'hbfba0190} /* (23, 25, 14) {real, imag} */,
  {32'hbe020700, 32'h3dd57f88} /* (23, 25, 13) {real, imag} */,
  {32'h3e1a3130, 32'h3f44a2da} /* (23, 25, 12) {real, imag} */,
  {32'h3ebd28f7, 32'hbe1d331c} /* (23, 25, 11) {real, imag} */,
  {32'hbfa3204f, 32'hbed4d3d4} /* (23, 25, 10) {real, imag} */,
  {32'hc024d0f2, 32'hbf913e82} /* (23, 25, 9) {real, imag} */,
  {32'hc022cc3f, 32'hc0095c2f} /* (23, 25, 8) {real, imag} */,
  {32'hbf09938d, 32'hbec53637} /* (23, 25, 7) {real, imag} */,
  {32'hbe8e6840, 32'hbe95e3cc} /* (23, 25, 6) {real, imag} */,
  {32'hc00f1ab7, 32'hbfc4985a} /* (23, 25, 5) {real, imag} */,
  {32'hbfcedde4, 32'h3e3d47cc} /* (23, 25, 4) {real, imag} */,
  {32'hbe901054, 32'h3f349956} /* (23, 25, 3) {real, imag} */,
  {32'hbf32fdf6, 32'hbe7ca398} /* (23, 25, 2) {real, imag} */,
  {32'hbfbc00bc, 32'hbf57df52} /* (23, 25, 1) {real, imag} */,
  {32'hbf0d6274, 32'h3d6f5510} /* (23, 25, 0) {real, imag} */,
  {32'h3dd98002, 32'hbf2fceba} /* (23, 24, 31) {real, imag} */,
  {32'hc01363e1, 32'hbf7c8ebe} /* (23, 24, 30) {real, imag} */,
  {32'hc03abea4, 32'hbf5f4660} /* (23, 24, 29) {real, imag} */,
  {32'hbf2e9a2e, 32'h3f3d1ba8} /* (23, 24, 28) {real, imag} */,
  {32'h3fcd4eb6, 32'hbf7078f9} /* (23, 24, 27) {real, imag} */,
  {32'hbf649da9, 32'hbf26cc5d} /* (23, 24, 26) {real, imag} */,
  {32'h3f40da37, 32'hbe3e66a6} /* (23, 24, 25) {real, imag} */,
  {32'h3fac3b4d, 32'hbf97b012} /* (23, 24, 24) {real, imag} */,
  {32'h400b5806, 32'hc01bce7c} /* (23, 24, 23) {real, imag} */,
  {32'h3fa6c2a9, 32'hbfcec392} /* (23, 24, 22) {real, imag} */,
  {32'hbec83429, 32'hbf6608b9} /* (23, 24, 21) {real, imag} */,
  {32'h3fafc3ec, 32'h3f1c5db1} /* (23, 24, 20) {real, imag} */,
  {32'h3fc4fe21, 32'h3f75a262} /* (23, 24, 19) {real, imag} */,
  {32'hbf2c7abe, 32'h3f311270} /* (23, 24, 18) {real, imag} */,
  {32'hc01b8e28, 32'h3f13ef4c} /* (23, 24, 17) {real, imag} */,
  {32'h3da8f428, 32'h3fa27fe8} /* (23, 24, 16) {real, imag} */,
  {32'h3f7b25b1, 32'h3fba7e78} /* (23, 24, 15) {real, imag} */,
  {32'h3eca540f, 32'h3fa41b21} /* (23, 24, 14) {real, imag} */,
  {32'hbba54c00, 32'h3f4ed846} /* (23, 24, 13) {real, imag} */,
  {32'h3ef04b68, 32'h3f5ccfdd} /* (23, 24, 12) {real, imag} */,
  {32'h3f5fbf88, 32'h3f64c86d} /* (23, 24, 11) {real, imag} */,
  {32'hbf913dba, 32'hbf0a7d54} /* (23, 24, 10) {real, imag} */,
  {32'h3ea7d256, 32'hbe827b40} /* (23, 24, 9) {real, imag} */,
  {32'h3de0e258, 32'hc00e1a41} /* (23, 24, 8) {real, imag} */,
  {32'h3f945d04, 32'hbed34000} /* (23, 24, 7) {real, imag} */,
  {32'h3f62a4ac, 32'h3f34b55a} /* (23, 24, 6) {real, imag} */,
  {32'hbd693000, 32'hbfa1ebc6} /* (23, 24, 5) {real, imag} */,
  {32'h3d2839e0, 32'hbf17ba7e} /* (23, 24, 4) {real, imag} */,
  {32'h3fdbba41, 32'h3fe282b6} /* (23, 24, 3) {real, imag} */,
  {32'h3f5c6f5d, 32'h3f56af58} /* (23, 24, 2) {real, imag} */,
  {32'hbf97fd6a, 32'h3f58ac1a} /* (23, 24, 1) {real, imag} */,
  {32'hbfa07ba2, 32'hbe0c4674} /* (23, 24, 0) {real, imag} */,
  {32'hbb9b2480, 32'hbf57acc5} /* (23, 23, 31) {real, imag} */,
  {32'hc0314a51, 32'hbf6db760} /* (23, 23, 30) {real, imag} */,
  {32'hc0331164, 32'h3e746688} /* (23, 23, 29) {real, imag} */,
  {32'hbfe726de, 32'hbed39cea} /* (23, 23, 28) {real, imag} */,
  {32'h3f0afdc4, 32'hbfacf223} /* (23, 23, 27) {real, imag} */,
  {32'h3f88c74e, 32'hbfbb4d82} /* (23, 23, 26) {real, imag} */,
  {32'h3f3b334c, 32'hbfde8eac} /* (23, 23, 25) {real, imag} */,
  {32'h3e4fa6fc, 32'hc0152209} /* (23, 23, 24) {real, imag} */,
  {32'hbf474b1a, 32'hc03492b2} /* (23, 23, 23) {real, imag} */,
  {32'hbf201cb6, 32'hbfe9f990} /* (23, 23, 22) {real, imag} */,
  {32'h3fd26a36, 32'hbf398134} /* (23, 23, 21) {real, imag} */,
  {32'h3f94fce1, 32'h3f6596b2} /* (23, 23, 20) {real, imag} */,
  {32'hbfa7a7e0, 32'h3f8777d9} /* (23, 23, 19) {real, imag} */,
  {32'hbfe900c4, 32'h3fb29535} /* (23, 23, 18) {real, imag} */,
  {32'hbfbc0fee, 32'h3fcbffee} /* (23, 23, 17) {real, imag} */,
  {32'hbe8d9bea, 32'h3fc854f7} /* (23, 23, 16) {real, imag} */,
  {32'h3f120b66, 32'h3fff6bdb} /* (23, 23, 15) {real, imag} */,
  {32'h3f26565e, 32'h3f52ab96} /* (23, 23, 14) {real, imag} */,
  {32'h3e5dbf9c, 32'hbfa053d9} /* (23, 23, 13) {real, imag} */,
  {32'h3f1b9a45, 32'hbf5a0560} /* (23, 23, 12) {real, imag} */,
  {32'h3f8d477a, 32'h3f1acd20} /* (23, 23, 11) {real, imag} */,
  {32'hbebb5bb4, 32'hbdc6d170} /* (23, 23, 10) {real, imag} */,
  {32'h3fb26581, 32'hbef409f0} /* (23, 23, 9) {real, imag} */,
  {32'h3f878f4e, 32'hbff3dcc3} /* (23, 23, 8) {real, imag} */,
  {32'h3ecc952c, 32'hbf216d56} /* (23, 23, 7) {real, imag} */,
  {32'h3f9e8efa, 32'hbf508306} /* (23, 23, 6) {real, imag} */,
  {32'h3f94ae4e, 32'h3eb5bec0} /* (23, 23, 5) {real, imag} */,
  {32'hbfabd5ce, 32'hbdf435a4} /* (23, 23, 4) {real, imag} */,
  {32'hbfa98592, 32'h3ed8691c} /* (23, 23, 3) {real, imag} */,
  {32'hbf39cac9, 32'h3e8d6cfc} /* (23, 23, 2) {real, imag} */,
  {32'hbe4e4da8, 32'hbd877110} /* (23, 23, 1) {real, imag} */,
  {32'hbf0ba168, 32'hbfabb84d} /* (23, 23, 0) {real, imag} */,
  {32'hbe7be3f8, 32'h3e3c6eae} /* (23, 22, 31) {real, imag} */,
  {32'hbfeea250, 32'hbf030e74} /* (23, 22, 30) {real, imag} */,
  {32'hbf369e6e, 32'h3e136760} /* (23, 22, 29) {real, imag} */,
  {32'hbf9543cd, 32'hc01409d1} /* (23, 22, 28) {real, imag} */,
  {32'hbe93d7af, 32'hc026396a} /* (23, 22, 27) {real, imag} */,
  {32'hbdea8288, 32'hbff4ffe3} /* (23, 22, 26) {real, imag} */,
  {32'h3f38490d, 32'hbfd57e80} /* (23, 22, 25) {real, imag} */,
  {32'h3e9c3c03, 32'hbf92b3e8} /* (23, 22, 24) {real, imag} */,
  {32'hc0033c8c, 32'hbfc1f909} /* (23, 22, 23) {real, imag} */,
  {32'hbd9d0370, 32'hbf95cf60} /* (23, 22, 22) {real, imag} */,
  {32'h40049768, 32'hbf1f6042} /* (23, 22, 21) {real, imag} */,
  {32'h3f5c7f72, 32'h3f853cca} /* (23, 22, 20) {real, imag} */,
  {32'hbfd337af, 32'h3f2a24fc} /* (23, 22, 19) {real, imag} */,
  {32'h3f3e72bf, 32'h3f5f7f96} /* (23, 22, 18) {real, imag} */,
  {32'h400981c5, 32'h3f31a8be} /* (23, 22, 17) {real, imag} */,
  {32'hbec19378, 32'h3f00476d} /* (23, 22, 16) {real, imag} */,
  {32'h3e699658, 32'h3f31749a} /* (23, 22, 15) {real, imag} */,
  {32'hbf1ae3c2, 32'hbec2ed3b} /* (23, 22, 14) {real, imag} */,
  {32'h3edb6864, 32'hbfbe1fde} /* (23, 22, 13) {real, imag} */,
  {32'h3fa5ac99, 32'hbfd61b38} /* (23, 22, 12) {real, imag} */,
  {32'h3dfd9b20, 32'hbf013e5a} /* (23, 22, 11) {real, imag} */,
  {32'hbf061cce, 32'h3c1dbb40} /* (23, 22, 10) {real, imag} */,
  {32'h3ea68484, 32'hbfc63a52} /* (23, 22, 9) {real, imag} */,
  {32'h402bc15c, 32'hbfaa5efc} /* (23, 22, 8) {real, imag} */,
  {32'hbe1d8878, 32'hbdfcf050} /* (23, 22, 7) {real, imag} */,
  {32'hbecf0892, 32'hbf9d1c04} /* (23, 22, 6) {real, imag} */,
  {32'hbfa3cd40, 32'h3e590458} /* (23, 22, 5) {real, imag} */,
  {32'hc000b585, 32'h3f3d4b6b} /* (23, 22, 4) {real, imag} */,
  {32'hc01189c6, 32'h3f4d9210} /* (23, 22, 3) {real, imag} */,
  {32'hbf8d2e12, 32'h3e8e0de8} /* (23, 22, 2) {real, imag} */,
  {32'h3e2abb18, 32'h3e84838c} /* (23, 22, 1) {real, imag} */,
  {32'h3e5ee3d6, 32'hbf14231b} /* (23, 22, 0) {real, imag} */,
  {32'h3dcb7498, 32'hbc66f840} /* (23, 21, 31) {real, imag} */,
  {32'hbe8b7f37, 32'hbea4ec9d} /* (23, 21, 30) {real, imag} */,
  {32'h3ff54dbe, 32'hbf593bfe} /* (23, 21, 29) {real, imag} */,
  {32'h3fb490fa, 32'hbfe8fed6} /* (23, 21, 28) {real, imag} */,
  {32'h3ef68a67, 32'hc01a0d77} /* (23, 21, 27) {real, imag} */,
  {32'hbfdb051e, 32'hc014d22a} /* (23, 21, 26) {real, imag} */,
  {32'h3ef79bde, 32'hbfbb4d8c} /* (23, 21, 25) {real, imag} */,
  {32'h3f80ed5c, 32'hbf5c50c2} /* (23, 21, 24) {real, imag} */,
  {32'hbefed22b, 32'hbfc94da1} /* (23, 21, 23) {real, imag} */,
  {32'h3fa38847, 32'hbf949a40} /* (23, 21, 22) {real, imag} */,
  {32'h3fa9aa6f, 32'hbf839cc5} /* (23, 21, 21) {real, imag} */,
  {32'h3f9b275a, 32'hbe2a4154} /* (23, 21, 20) {real, imag} */,
  {32'h3e1c7bc4, 32'hbf32dc12} /* (23, 21, 19) {real, imag} */,
  {32'hbf17dd5c, 32'hbedfd9f0} /* (23, 21, 18) {real, imag} */,
  {32'h3f9c25d6, 32'hbf348521} /* (23, 21, 17) {real, imag} */,
  {32'h3ed69336, 32'hc0067598} /* (23, 21, 16) {real, imag} */,
  {32'hbdeedde0, 32'hbf3d6dea} /* (23, 21, 15) {real, imag} */,
  {32'hc00b7bf0, 32'hbf6abd4b} /* (23, 21, 14) {real, imag} */,
  {32'h3f17e6dc, 32'hbf917247} /* (23, 21, 13) {real, imag} */,
  {32'h400615d2, 32'hbe1cc227} /* (23, 21, 12) {real, imag} */,
  {32'h3f93012f, 32'h3f13b565} /* (23, 21, 11) {real, imag} */,
  {32'hbf9a35ea, 32'h3ebd0de6} /* (23, 21, 10) {real, imag} */,
  {32'hbff62f12, 32'hc010f021} /* (23, 21, 9) {real, imag} */,
  {32'h3f8191ad, 32'hc03741ef} /* (23, 21, 8) {real, imag} */,
  {32'h3ec26816, 32'hbf99b049} /* (23, 21, 7) {real, imag} */,
  {32'hbeb79e4e, 32'hbf544f8a} /* (23, 21, 6) {real, imag} */,
  {32'hbfa12447, 32'hbf886cd9} /* (23, 21, 5) {real, imag} */,
  {32'h3e81c779, 32'h3f36a96c} /* (23, 21, 4) {real, imag} */,
  {32'hbed73586, 32'h3fe41004} /* (23, 21, 3) {real, imag} */,
  {32'hbfa6bdc0, 32'h3f0b6292} /* (23, 21, 2) {real, imag} */,
  {32'hbed8b88b, 32'hbe0958f0} /* (23, 21, 1) {real, imag} */,
  {32'h3f44178a, 32'hbebd40dc} /* (23, 21, 0) {real, imag} */,
  {32'h3e619da4, 32'h3f6186d3} /* (23, 20, 31) {real, imag} */,
  {32'hbf6227b4, 32'h3e103346} /* (23, 20, 30) {real, imag} */,
  {32'h3f55a71c, 32'h3e4f5b68} /* (23, 20, 29) {real, imag} */,
  {32'h3f61e31f, 32'h3fbbfc52} /* (23, 20, 28) {real, imag} */,
  {32'h3fa76bae, 32'hbda1c388} /* (23, 20, 27) {real, imag} */,
  {32'hbd4d2a00, 32'hbfac30fa} /* (23, 20, 26) {real, imag} */,
  {32'h3ef35b70, 32'h3ed1a014} /* (23, 20, 25) {real, imag} */,
  {32'h3f93bce7, 32'h3fa9ef0d} /* (23, 20, 24) {real, imag} */,
  {32'h3f2e8ba6, 32'h3f7f6eac} /* (23, 20, 23) {real, imag} */,
  {32'hbea0c3ba, 32'hbeb28050} /* (23, 20, 22) {real, imag} */,
  {32'h3df55fc0, 32'hbf4440b4} /* (23, 20, 21) {real, imag} */,
  {32'h3eccc3a8, 32'hbed215b4} /* (23, 20, 20) {real, imag} */,
  {32'h3fda58cf, 32'hbfdc7ae8} /* (23, 20, 19) {real, imag} */,
  {32'hbf09cb76, 32'hc00319a6} /* (23, 20, 18) {real, imag} */,
  {32'hbf2a4ee5, 32'hbed04bfc} /* (23, 20, 17) {real, imag} */,
  {32'h3f41eb58, 32'hbfbf937c} /* (23, 20, 16) {real, imag} */,
  {32'hbf790b53, 32'hbf53e22b} /* (23, 20, 15) {real, imag} */,
  {32'hbff0899e, 32'hbf51620e} /* (23, 20, 14) {real, imag} */,
  {32'hbeeeed47, 32'hbf6aab39} /* (23, 20, 13) {real, imag} */,
  {32'h3ee3bf34, 32'hbec00c38} /* (23, 20, 12) {real, imag} */,
  {32'h3fcd4406, 32'h3f2dcbe4} /* (23, 20, 11) {real, imag} */,
  {32'h3eb4ac48, 32'h3f1f0070} /* (23, 20, 10) {real, imag} */,
  {32'hbebc7ea8, 32'hbff01a97} /* (23, 20, 9) {real, imag} */,
  {32'h3f96a434, 32'h3f00d8bc} /* (23, 20, 8) {real, imag} */,
  {32'h40185dca, 32'h3f69e73a} /* (23, 20, 7) {real, imag} */,
  {32'h3f1f0d05, 32'hbf22e990} /* (23, 20, 6) {real, imag} */,
  {32'hbf03b229, 32'hbfeaaa8b} /* (23, 20, 5) {real, imag} */,
  {32'h40126759, 32'hbead5292} /* (23, 20, 4) {real, imag} */,
  {32'h3f4e0224, 32'h400399e6} /* (23, 20, 3) {real, imag} */,
  {32'hbfc4a0aa, 32'h401181a4} /* (23, 20, 2) {real, imag} */,
  {32'hbf5e0061, 32'h3fa77e55} /* (23, 20, 1) {real, imag} */,
  {32'h3f5e9c95, 32'h3f5f917c} /* (23, 20, 0) {real, imag} */,
  {32'hbe17b3ce, 32'h3fea7a84} /* (23, 19, 31) {real, imag} */,
  {32'h3e885714, 32'h3f9203ee} /* (23, 19, 30) {real, imag} */,
  {32'h3f333d62, 32'hbf8ae1bc} /* (23, 19, 29) {real, imag} */,
  {32'hbef8ce7c, 32'h3f77cfdf} /* (23, 19, 28) {real, imag} */,
  {32'h3eec9318, 32'h3fbac2e6} /* (23, 19, 27) {real, imag} */,
  {32'h3f14f559, 32'h3d048510} /* (23, 19, 26) {real, imag} */,
  {32'h3f58a6aa, 32'h3d9dd900} /* (23, 19, 25) {real, imag} */,
  {32'h3f908d86, 32'h4001dfea} /* (23, 19, 24) {real, imag} */,
  {32'hbe24b8a8, 32'h4004bd9e} /* (23, 19, 23) {real, imag} */,
  {32'hc00105aa, 32'h3f9fa25e} /* (23, 19, 22) {real, imag} */,
  {32'hbd5b8800, 32'h3ef55b54} /* (23, 19, 21) {real, imag} */,
  {32'hbe3b9338, 32'h3f7fe115} /* (23, 19, 20) {real, imag} */,
  {32'h3fb234bc, 32'hbf47789a} /* (23, 19, 19) {real, imag} */,
  {32'h3e7bfe4c, 32'hbfde67e0} /* (23, 19, 18) {real, imag} */,
  {32'hbf2d96d0, 32'hbf810204} /* (23, 19, 17) {real, imag} */,
  {32'h3f3c2169, 32'hbf5dc8c0} /* (23, 19, 16) {real, imag} */,
  {32'hbecea625, 32'h3e8df80d} /* (23, 19, 15) {real, imag} */,
  {32'hbf6e855c, 32'hbe105082} /* (23, 19, 14) {real, imag} */,
  {32'hbf14ab0d, 32'hbe9e1391} /* (23, 19, 13) {real, imag} */,
  {32'hbfdc5f56, 32'hbf85886c} /* (23, 19, 12) {real, imag} */,
  {32'hbf6fd08d, 32'h3eb222bc} /* (23, 19, 11) {real, imag} */,
  {32'h3ea7c92a, 32'hbf901d6a} /* (23, 19, 10) {real, imag} */,
  {32'h3fa8eb68, 32'hc0209fc7} /* (23, 19, 9) {real, imag} */,
  {32'h40182cbe, 32'h3e7c6ea8} /* (23, 19, 8) {real, imag} */,
  {32'h4053146f, 32'h3fb5a884} /* (23, 19, 7) {real, imag} */,
  {32'h3fe0cd09, 32'h3ecf4e7a} /* (23, 19, 6) {real, imag} */,
  {32'h3ea76292, 32'h3f41891e} /* (23, 19, 5) {real, imag} */,
  {32'h3f4926a6, 32'h3ed2afe5} /* (23, 19, 4) {real, imag} */,
  {32'h3f9a9746, 32'h3f98c440} /* (23, 19, 3) {real, imag} */,
  {32'hbe2a9e3c, 32'h3f35e45f} /* (23, 19, 2) {real, imag} */,
  {32'hbfcf38c4, 32'h3f4da4f5} /* (23, 19, 1) {real, imag} */,
  {32'hbf8d568e, 32'h3fa76c57} /* (23, 19, 0) {real, imag} */,
  {32'h3f55a572, 32'h3f77edc8} /* (23, 18, 31) {real, imag} */,
  {32'h3f2e38fc, 32'h3f33be1c} /* (23, 18, 30) {real, imag} */,
  {32'h3f59aac8, 32'hc00a7616} /* (23, 18, 29) {real, imag} */,
  {32'h3e917174, 32'hbfd3dbb3} /* (23, 18, 28) {real, imag} */,
  {32'h3d211b80, 32'hbe146204} /* (23, 18, 27) {real, imag} */,
  {32'hbefe60f8, 32'h3ea6998e} /* (23, 18, 26) {real, imag} */,
  {32'hbd117740, 32'h3f87d990} /* (23, 18, 25) {real, imag} */,
  {32'h3fc35e27, 32'h4003a050} /* (23, 18, 24) {real, imag} */,
  {32'h3e309378, 32'hbf2f42a8} /* (23, 18, 23) {real, imag} */,
  {32'hbfde22b1, 32'hbf55a610} /* (23, 18, 22) {real, imag} */,
  {32'hbfc26b2c, 32'hbe671ce8} /* (23, 18, 21) {real, imag} */,
  {32'hbf5795c6, 32'h3f805700} /* (23, 18, 20) {real, imag} */,
  {32'h3f567150, 32'h3f297c6a} /* (23, 18, 19) {real, imag} */,
  {32'h3e66f2a0, 32'h3f993d5a} /* (23, 18, 18) {real, imag} */,
  {32'hbebb8f58, 32'h3f2604fc} /* (23, 18, 17) {real, imag} */,
  {32'h3f8b6b82, 32'hbfe5ca5a} /* (23, 18, 16) {real, imag} */,
  {32'h3dcbe360, 32'hbf7fb3aa} /* (23, 18, 15) {real, imag} */,
  {32'hbeddf2e6, 32'hbfd87a85} /* (23, 18, 14) {real, imag} */,
  {32'hbfe777df, 32'hc0585b86} /* (23, 18, 13) {real, imag} */,
  {32'hc042d884, 32'hc00e7b1e} /* (23, 18, 12) {real, imag} */,
  {32'hc02ea6e8, 32'hbeae5fb6} /* (23, 18, 11) {real, imag} */,
  {32'hbf9822ce, 32'hbfd0503e} /* (23, 18, 10) {real, imag} */,
  {32'h3fc332c4, 32'hbf7ff242} /* (23, 18, 9) {real, imag} */,
  {32'h3ff9892a, 32'h3f9698ca} /* (23, 18, 8) {real, imag} */,
  {32'h3fc4eeb0, 32'h40138b0d} /* (23, 18, 7) {real, imag} */,
  {32'h3f94557a, 32'h401e0220} /* (23, 18, 6) {real, imag} */,
  {32'hbd93c4e0, 32'h400c0e82} /* (23, 18, 5) {real, imag} */,
  {32'hbf52501e, 32'h3faccbfd} /* (23, 18, 4) {real, imag} */,
  {32'h3efcf6f0, 32'hbf0d28ae} /* (23, 18, 3) {real, imag} */,
  {32'h3f289045, 32'hbf8d1c43} /* (23, 18, 2) {real, imag} */,
  {32'hc010969e, 32'hbed32c98} /* (23, 18, 1) {real, imag} */,
  {32'hc01be1d2, 32'hbea7c69a} /* (23, 18, 0) {real, imag} */,
  {32'h3dfba898, 32'hbeb7aa40} /* (23, 17, 31) {real, imag} */,
  {32'h3f92078c, 32'hbf882eab} /* (23, 17, 30) {real, imag} */,
  {32'h402278a4, 32'hbefa73a6} /* (23, 17, 29) {real, imag} */,
  {32'h4022a5d5, 32'hbffc88c3} /* (23, 17, 28) {real, imag} */,
  {32'h3f998c9e, 32'hbf680c48} /* (23, 17, 27) {real, imag} */,
  {32'hbef1820c, 32'h3f86ea06} /* (23, 17, 26) {real, imag} */,
  {32'hbf7f33f2, 32'h401b459a} /* (23, 17, 25) {real, imag} */,
  {32'h3f924e17, 32'h3fc30ab6} /* (23, 17, 24) {real, imag} */,
  {32'h3f6f7d18, 32'h3e7468d8} /* (23, 17, 23) {real, imag} */,
  {32'hbf951849, 32'h3f80319f} /* (23, 17, 22) {real, imag} */,
  {32'hc002dbbd, 32'hbe9fd770} /* (23, 17, 21) {real, imag} */,
  {32'hc014469a, 32'hbf1fe3e8} /* (23, 17, 20) {real, imag} */,
  {32'hbed53966, 32'hbf11e6f5} /* (23, 17, 19) {real, imag} */,
  {32'h3f301932, 32'hbd67a500} /* (23, 17, 18) {real, imag} */,
  {32'hbf7b8456, 32'h3f56c116} /* (23, 17, 17) {real, imag} */,
  {32'hbdf88810, 32'hbe89d73e} /* (23, 17, 16) {real, imag} */,
  {32'h3eb66d96, 32'hbf2ef9a6} /* (23, 17, 15) {real, imag} */,
  {32'h3f6d6220, 32'hbf35da58} /* (23, 17, 14) {real, imag} */,
  {32'hbfa17d5d, 32'hc018a46c} /* (23, 17, 13) {real, imag} */,
  {32'hc00f998d, 32'hc066c3c0} /* (23, 17, 12) {real, imag} */,
  {32'hbfdc1f47, 32'hbfeca30e} /* (23, 17, 11) {real, imag} */,
  {32'h3e987e68, 32'h3e85a894} /* (23, 17, 10) {real, imag} */,
  {32'h3fad46c0, 32'h4004d55d} /* (23, 17, 9) {real, imag} */,
  {32'h3ec7be78, 32'h40141810} /* (23, 17, 8) {real, imag} */,
  {32'h3e3bcb06, 32'h40354e7e} /* (23, 17, 7) {real, imag} */,
  {32'hbeb92b78, 32'h4080024c} /* (23, 17, 6) {real, imag} */,
  {32'h3eaa9ebe, 32'h3f9d6fad} /* (23, 17, 5) {real, imag} */,
  {32'hbec4f97d, 32'hbe92a8c9} /* (23, 17, 4) {real, imag} */,
  {32'hbb7bd000, 32'hbfbef7b4} /* (23, 17, 3) {real, imag} */,
  {32'h3ee98bc5, 32'hbea2263a} /* (23, 17, 2) {real, imag} */,
  {32'hbfa863ba, 32'hbe563ec8} /* (23, 17, 1) {real, imag} */,
  {32'hbfb61712, 32'hbf84f17c} /* (23, 17, 0) {real, imag} */,
  {32'h3dbf003c, 32'hbfc98f82} /* (23, 16, 31) {real, imag} */,
  {32'h40076c81, 32'hbfe41b2f} /* (23, 16, 30) {real, imag} */,
  {32'h4048aa28, 32'h3f8dd590} /* (23, 16, 29) {real, imag} */,
  {32'h3f7dcce8, 32'h3f9c65c0} /* (23, 16, 28) {real, imag} */,
  {32'hbde012bc, 32'h3f7e3bee} /* (23, 16, 27) {real, imag} */,
  {32'h3f3cdacc, 32'h3fdb28f6} /* (23, 16, 26) {real, imag} */,
  {32'h3ecf4da4, 32'h3feebae1} /* (23, 16, 25) {real, imag} */,
  {32'h3d8897f0, 32'h3f1d25e7} /* (23, 16, 24) {real, imag} */,
  {32'h3ce87df0, 32'h40153304} /* (23, 16, 23) {real, imag} */,
  {32'hbdf98b30, 32'h401abcd6} /* (23, 16, 22) {real, imag} */,
  {32'hbf55166c, 32'h3ed070e2} /* (23, 16, 21) {real, imag} */,
  {32'hc000b2b4, 32'hbd657400} /* (23, 16, 20) {real, imag} */,
  {32'hbfe12499, 32'h3f12c3da} /* (23, 16, 19) {real, imag} */,
  {32'hbe0a9e1c, 32'hbf2e9b3c} /* (23, 16, 18) {real, imag} */,
  {32'h3ef35250, 32'hbf9caee6} /* (23, 16, 17) {real, imag} */,
  {32'h3f2e7963, 32'hbfd236ae} /* (23, 16, 16) {real, imag} */,
  {32'hbf5870a6, 32'hbfa2417a} /* (23, 16, 15) {real, imag} */,
  {32'hbee8197a, 32'h3f1dc990} /* (23, 16, 14) {real, imag} */,
  {32'hc01442f4, 32'h3f9361f4} /* (23, 16, 13) {real, imag} */,
  {32'hc0269b82, 32'hbf19417f} /* (23, 16, 12) {real, imag} */,
  {32'h3e17ac40, 32'hc002168c} /* (23, 16, 11) {real, imag} */,
  {32'h3f9f38ea, 32'hbf173a95} /* (23, 16, 10) {real, imag} */,
  {32'h3f9943aa, 32'h3fbd0efa} /* (23, 16, 9) {real, imag} */,
  {32'hbf17e280, 32'h400d4b5a} /* (23, 16, 8) {real, imag} */,
  {32'hbce2af30, 32'h4039cbea} /* (23, 16, 7) {real, imag} */,
  {32'h3fb6ca36, 32'h403d8e8a} /* (23, 16, 6) {real, imag} */,
  {32'h3f8feaac, 32'hbeacc34c} /* (23, 16, 5) {real, imag} */,
  {32'h3fa57aa9, 32'hbf2bc0ac} /* (23, 16, 4) {real, imag} */,
  {32'h3f943e36, 32'hc007f5c8} /* (23, 16, 3) {real, imag} */,
  {32'hbf1ffc5c, 32'hbf2a6292} /* (23, 16, 2) {real, imag} */,
  {32'h3f450ef2, 32'h3f353e24} /* (23, 16, 1) {real, imag} */,
  {32'h3f754d30, 32'hbf3f21ce} /* (23, 16, 0) {real, imag} */,
  {32'h3e0d1d0c, 32'hbf87d2aa} /* (23, 15, 31) {real, imag} */,
  {32'h3f4d0d44, 32'hbf91484a} /* (23, 15, 30) {real, imag} */,
  {32'h3f8c1687, 32'h3f6290f6} /* (23, 15, 29) {real, imag} */,
  {32'h3f86f330, 32'h4036053e} /* (23, 15, 28) {real, imag} */,
  {32'h3e678cd0, 32'h400e35a6} /* (23, 15, 27) {real, imag} */,
  {32'hbf16517e, 32'h3faca61e} /* (23, 15, 26) {real, imag} */,
  {32'h3f76349c, 32'h3ebadf9c} /* (23, 15, 25) {real, imag} */,
  {32'hbe7e8164, 32'h3fd54622} /* (23, 15, 24) {real, imag} */,
  {32'hbf097bb6, 32'h4066305c} /* (23, 15, 23) {real, imag} */,
  {32'h3f72c1ce, 32'h4009b36e} /* (23, 15, 22) {real, imag} */,
  {32'h401c8ce8, 32'h3e525268} /* (23, 15, 21) {real, imag} */,
  {32'h3f84bbcc, 32'hbf8aaa1a} /* (23, 15, 20) {real, imag} */,
  {32'hbe840eac, 32'hbf949ee2} /* (23, 15, 19) {real, imag} */,
  {32'hbf1fc523, 32'hbf4c2cca} /* (23, 15, 18) {real, imag} */,
  {32'h3ee52e4c, 32'hbf987bc6} /* (23, 15, 17) {real, imag} */,
  {32'h3f8a54fc, 32'hbf9cc526} /* (23, 15, 16) {real, imag} */,
  {32'hbe42c4a0, 32'hbfaf6b93} /* (23, 15, 15) {real, imag} */,
  {32'hbf48a430, 32'h3de69870} /* (23, 15, 14) {real, imag} */,
  {32'hbf429092, 32'hbe460032} /* (23, 15, 13) {real, imag} */,
  {32'hbfa0af4d, 32'h3e8c0a74} /* (23, 15, 12) {real, imag} */,
  {32'hbf2dc800, 32'hbfb06d29} /* (23, 15, 11) {real, imag} */,
  {32'h3f5697c5, 32'hbfde3032} /* (23, 15, 10) {real, imag} */,
  {32'h3e054630, 32'h3ec7bed4} /* (23, 15, 9) {real, imag} */,
  {32'hbf8f6d82, 32'h3ff94714} /* (23, 15, 8) {real, imag} */,
  {32'hbf8aad03, 32'h3fbd95a2} /* (23, 15, 7) {real, imag} */,
  {32'h3e993eb0, 32'h3faf54b6} /* (23, 15, 6) {real, imag} */,
  {32'h3f1b6f5b, 32'hbf61a9ba} /* (23, 15, 5) {real, imag} */,
  {32'h3fd7b25e, 32'h3e01e920} /* (23, 15, 4) {real, imag} */,
  {32'h3f104706, 32'hbfb12fde} /* (23, 15, 3) {real, imag} */,
  {32'hbf01d0c0, 32'hbecb5d26} /* (23, 15, 2) {real, imag} */,
  {32'h3fc55dcb, 32'h403eb2b0} /* (23, 15, 1) {real, imag} */,
  {32'h3fe2683b, 32'h3efd23e8} /* (23, 15, 0) {real, imag} */,
  {32'h3ecd21e0, 32'hbe20d218} /* (23, 14, 31) {real, imag} */,
  {32'h3f1bcdc7, 32'hbeded44c} /* (23, 14, 30) {real, imag} */,
  {32'hbe3c79bb, 32'hbf787228} /* (23, 14, 29) {real, imag} */,
  {32'h3f981aa8, 32'h3ec62d71} /* (23, 14, 28) {real, imag} */,
  {32'h3ffd15be, 32'h3f2d59be} /* (23, 14, 27) {real, imag} */,
  {32'h3fc34538, 32'h3e91000a} /* (23, 14, 26) {real, imag} */,
  {32'h3fc0ae3e, 32'hbd64a500} /* (23, 14, 25) {real, imag} */,
  {32'hbf658cb5, 32'h3f3f8f5e} /* (23, 14, 24) {real, imag} */,
  {32'hbef04b85, 32'h3ef2e131} /* (23, 14, 23) {real, imag} */,
  {32'h3f929dcf, 32'hbfb6b74e} /* (23, 14, 22) {real, imag} */,
  {32'h3fb0181b, 32'hc03fbb5d} /* (23, 14, 21) {real, imag} */,
  {32'h3fdccb1e, 32'hbff8b6e5} /* (23, 14, 20) {real, imag} */,
  {32'h3fdb61fd, 32'hb875c000} /* (23, 14, 19) {real, imag} */,
  {32'hbeecf41e, 32'hbdd8ea40} /* (23, 14, 18) {real, imag} */,
  {32'h3e856892, 32'hbfa224fe} /* (23, 14, 17) {real, imag} */,
  {32'h3bed6580, 32'hbf942d46} /* (23, 14, 16) {real, imag} */,
  {32'hbf149fd2, 32'hbfa74770} /* (23, 14, 15) {real, imag} */,
  {32'h3d3ac340, 32'hbeed0c94} /* (23, 14, 14) {real, imag} */,
  {32'h3efabc46, 32'hbfbd64fe} /* (23, 14, 13) {real, imag} */,
  {32'h3e5ec9c0, 32'h3f2c8146} /* (23, 14, 12) {real, imag} */,
  {32'hbea45688, 32'h3f86df2c} /* (23, 14, 11) {real, imag} */,
  {32'h3eeff4c7, 32'h3f9e246a} /* (23, 14, 10) {real, imag} */,
  {32'hbed26f10, 32'h3f5001c6} /* (23, 14, 9) {real, imag} */,
  {32'hbf48aa4d, 32'h3df5f2f4} /* (23, 14, 8) {real, imag} */,
  {32'h3f5992b4, 32'h3dd2e550} /* (23, 14, 7) {real, imag} */,
  {32'h3ecbd3c0, 32'hbe08baee} /* (23, 14, 6) {real, imag} */,
  {32'h3f87580d, 32'hbf4b20b4} /* (23, 14, 5) {real, imag} */,
  {32'h3f049962, 32'h3e4e1cae} /* (23, 14, 4) {real, imag} */,
  {32'hbfbff6d1, 32'h3d99ca60} /* (23, 14, 3) {real, imag} */,
  {32'h3f126d97, 32'hbf93ffd1} /* (23, 14, 2) {real, imag} */,
  {32'h40082d60, 32'h3e518420} /* (23, 14, 1) {real, imag} */,
  {32'h3fad86a0, 32'h3d67ccb0} /* (23, 14, 0) {real, imag} */,
  {32'h3ec5737e, 32'hbec3bb3c} /* (23, 13, 31) {real, imag} */,
  {32'h3f024f28, 32'hbedf09a3} /* (23, 13, 30) {real, imag} */,
  {32'hbf379b88, 32'hbeaa1cbe} /* (23, 13, 29) {real, imag} */,
  {32'hbeba4d48, 32'hbe786eaa} /* (23, 13, 28) {real, imag} */,
  {32'h3eccb8d6, 32'h3f8ddc78} /* (23, 13, 27) {real, imag} */,
  {32'hbe123c70, 32'h3f7266f9} /* (23, 13, 26) {real, imag} */,
  {32'h3f066cbb, 32'hbd907b20} /* (23, 13, 25) {real, imag} */,
  {32'h3efe5b7c, 32'hbfa00838} /* (23, 13, 24) {real, imag} */,
  {32'h3f0def3c, 32'hc00bcbe6} /* (23, 13, 23) {real, imag} */,
  {32'h3f97180f, 32'hc028a6dc} /* (23, 13, 22) {real, imag} */,
  {32'h3f2306ce, 32'hc018c1d0} /* (23, 13, 21) {real, imag} */,
  {32'h3fc21184, 32'hc04f6486} /* (23, 13, 20) {real, imag} */,
  {32'h3fb423d9, 32'hbf926b66} /* (23, 13, 19) {real, imag} */,
  {32'h3f33d9ba, 32'hbe9069fc} /* (23, 13, 18) {real, imag} */,
  {32'h3abdf400, 32'hc0003746} /* (23, 13, 17) {real, imag} */,
  {32'hbf45211a, 32'hbfb72ead} /* (23, 13, 16) {real, imag} */,
  {32'hbda67c7c, 32'hbf5cbf28} /* (23, 13, 15) {real, imag} */,
  {32'h3e54aaba, 32'hbd4f36d0} /* (23, 13, 14) {real, imag} */,
  {32'h3fbe7e3b, 32'hbf6015b4} /* (23, 13, 13) {real, imag} */,
  {32'h3fb6970f, 32'h3e8667c0} /* (23, 13, 12) {real, imag} */,
  {32'h3e3f7308, 32'h3f82b27c} /* (23, 13, 11) {real, imag} */,
  {32'h3f82f87e, 32'h3fcef621} /* (23, 13, 10) {real, imag} */,
  {32'h3ce37b00, 32'h4016982a} /* (23, 13, 9) {real, imag} */,
  {32'h3e6ea888, 32'h3ebf90ec} /* (23, 13, 8) {real, imag} */,
  {32'h4066eaac, 32'h3fbfb7f0} /* (23, 13, 7) {real, imag} */,
  {32'h3f99639c, 32'hbd2bc7dc} /* (23, 13, 6) {real, imag} */,
  {32'h3fc4e7c4, 32'hbf8c9d05} /* (23, 13, 5) {real, imag} */,
  {32'h3fe22e11, 32'hbf8dfa44} /* (23, 13, 4) {real, imag} */,
  {32'h3f1b32b0, 32'h3eb75fa8} /* (23, 13, 3) {real, imag} */,
  {32'h3f9caded, 32'hbf140558} /* (23, 13, 2) {real, imag} */,
  {32'h3fdf550c, 32'hbfa95916} /* (23, 13, 1) {real, imag} */,
  {32'h3f9249a4, 32'hbe589f24} /* (23, 13, 0) {real, imag} */,
  {32'h3fa23c3b, 32'hbdab7420} /* (23, 12, 31) {real, imag} */,
  {32'h3f557768, 32'h3f68f2da} /* (23, 12, 30) {real, imag} */,
  {32'hbf8e6fa2, 32'h3fc1c6f2} /* (23, 12, 29) {real, imag} */,
  {32'hbf752812, 32'h3f8e84ff} /* (23, 12, 28) {real, imag} */,
  {32'hbf0fabae, 32'h3ea86538} /* (23, 12, 27) {real, imag} */,
  {32'hbf9ca0f1, 32'h3fda8ba7} /* (23, 12, 26) {real, imag} */,
  {32'h3dc0fa80, 32'hbf18df33} /* (23, 12, 25) {real, imag} */,
  {32'h3f08b186, 32'hbf001cb6} /* (23, 12, 24) {real, imag} */,
  {32'h3f150ebd, 32'h3fe32d3f} /* (23, 12, 23) {real, imag} */,
  {32'h3fc7e58a, 32'h3fb3ccf3} /* (23, 12, 22) {real, imag} */,
  {32'hbea6e1f8, 32'h3f8cbaa0} /* (23, 12, 21) {real, imag} */,
  {32'h3eced6a6, 32'hbf822546} /* (23, 12, 20) {real, imag} */,
  {32'h3f31c9de, 32'hbfe6549d} /* (23, 12, 19) {real, imag} */,
  {32'h3f204ff4, 32'h3e4534c0} /* (23, 12, 18) {real, imag} */,
  {32'hbc446280, 32'hbfb1c2a2} /* (23, 12, 17) {real, imag} */,
  {32'hbf48aa14, 32'h3ee57300} /* (23, 12, 16) {real, imag} */,
  {32'h3e5b2888, 32'h3fcb1db5} /* (23, 12, 15) {real, imag} */,
  {32'hbe3d5930, 32'hbe145718} /* (23, 12, 14) {real, imag} */,
  {32'h3fb97758, 32'hbf884c6d} /* (23, 12, 13) {real, imag} */,
  {32'h3ff21250, 32'hbff73cb5} /* (23, 12, 12) {real, imag} */,
  {32'h3ec31498, 32'hbd7a3440} /* (23, 12, 11) {real, imag} */,
  {32'h4003760e, 32'h3f27573d} /* (23, 12, 10) {real, imag} */,
  {32'h3f95dd70, 32'hbef2ba02} /* (23, 12, 9) {real, imag} */,
  {32'hbe22f2d8, 32'hbf3520f0} /* (23, 12, 8) {real, imag} */,
  {32'h40270a56, 32'h3f9d0af2} /* (23, 12, 7) {real, imag} */,
  {32'h40109458, 32'h3f77c310} /* (23, 12, 6) {real, imag} */,
  {32'h40069107, 32'h3ef4ab82} /* (23, 12, 5) {real, imag} */,
  {32'h3f8366c6, 32'hbeedc1d7} /* (23, 12, 4) {real, imag} */,
  {32'hbe3fbf34, 32'hbf8dd542} /* (23, 12, 3) {real, imag} */,
  {32'hbfcf3bc9, 32'hbf3cdc77} /* (23, 12, 2) {real, imag} */,
  {32'hbf5e9403, 32'hbfb79692} /* (23, 12, 1) {real, imag} */,
  {32'h3e9733fd, 32'hbe943874} /* (23, 12, 0) {real, imag} */,
  {32'hbd911e38, 32'hbc941a80} /* (23, 11, 31) {real, imag} */,
  {32'hbf5e98a4, 32'hbe1a179c} /* (23, 11, 30) {real, imag} */,
  {32'hbfb61d2b, 32'h3cd27898} /* (23, 11, 29) {real, imag} */,
  {32'hbfa10f62, 32'h3f91fa42} /* (23, 11, 28) {real, imag} */,
  {32'hc00c2bae, 32'h3f7df227} /* (23, 11, 27) {real, imag} */,
  {32'hbff0b211, 32'h3fc9b9e0} /* (23, 11, 26) {real, imag} */,
  {32'hbe4f2c0a, 32'hbe9f25b2} /* (23, 11, 25) {real, imag} */,
  {32'h3df0dc18, 32'hbf1e4802} /* (23, 11, 24) {real, imag} */,
  {32'h3da7bb40, 32'h3e64e6ac} /* (23, 11, 23) {real, imag} */,
  {32'h3f9f7e65, 32'h3fdba72c} /* (23, 11, 22) {real, imag} */,
  {32'hbf0bffb2, 32'h3fa9df96} /* (23, 11, 21) {real, imag} */,
  {32'hbf843dc7, 32'h3f221f27} /* (23, 11, 20) {real, imag} */,
  {32'h3f38de53, 32'h3f5cc52a} /* (23, 11, 19) {real, imag} */,
  {32'hbf898b4d, 32'hbc245700} /* (23, 11, 18) {real, imag} */,
  {32'hbff6fcac, 32'hc00aa00a} /* (23, 11, 17) {real, imag} */,
  {32'h3d7b7770, 32'h3f9066e4} /* (23, 11, 16) {real, imag} */,
  {32'h3e033b02, 32'h3f5e5684} /* (23, 11, 15) {real, imag} */,
  {32'hbfa5e907, 32'hc020c0ec} /* (23, 11, 14) {real, imag} */,
  {32'h3f90e368, 32'hc02dba98} /* (23, 11, 13) {real, imag} */,
  {32'h40331ca2, 32'hc014372c} /* (23, 11, 12) {real, imag} */,
  {32'h3f96ac68, 32'h3eb4d0f4} /* (23, 11, 11) {real, imag} */,
  {32'h3fe20aa4, 32'h3f679c66} /* (23, 11, 10) {real, imag} */,
  {32'h3fd1dcbe, 32'hc025ada3} /* (23, 11, 9) {real, imag} */,
  {32'hbd4d38a0, 32'hbf8416be} /* (23, 11, 8) {real, imag} */,
  {32'h3f5c84a8, 32'hbe9bb48e} /* (23, 11, 7) {real, imag} */,
  {32'h3f8cb68f, 32'hbdd3a840} /* (23, 11, 6) {real, imag} */,
  {32'h3fb93dcd, 32'h3e1d74c0} /* (23, 11, 5) {real, imag} */,
  {32'h3d42bdd8, 32'h3f13e48e} /* (23, 11, 4) {real, imag} */,
  {32'hbe237afc, 32'hbef92bde} /* (23, 11, 3) {real, imag} */,
  {32'h3e8b944c, 32'hbed7fe08} /* (23, 11, 2) {real, imag} */,
  {32'h3ece6311, 32'hbf7e36f6} /* (23, 11, 1) {real, imag} */,
  {32'hbeb03ca2, 32'hbea180aa} /* (23, 11, 0) {real, imag} */,
  {32'h3d868afe, 32'hbf8871ca} /* (23, 10, 31) {real, imag} */,
  {32'hbfab76da, 32'hbe21e3e4} /* (23, 10, 30) {real, imag} */,
  {32'hbf892121, 32'hbf44ddb8} /* (23, 10, 29) {real, imag} */,
  {32'hbf8c5e8f, 32'hbf24f2f4} /* (23, 10, 28) {real, imag} */,
  {32'hc010d618, 32'h3f8bcd60} /* (23, 10, 27) {real, imag} */,
  {32'hbfd57668, 32'h3f8aeb20} /* (23, 10, 26) {real, imag} */,
  {32'hbf84f6a1, 32'hbfa63364} /* (23, 10, 25) {real, imag} */,
  {32'hbe3e15cf, 32'hc03b49c8} /* (23, 10, 24) {real, imag} */,
  {32'hbebd6174, 32'hc0284d40} /* (23, 10, 23) {real, imag} */,
  {32'h3eb465aa, 32'hbedbe9c0} /* (23, 10, 22) {real, imag} */,
  {32'h3f482e9a, 32'hbfa43926} /* (23, 10, 21) {real, imag} */,
  {32'h3f1af997, 32'h3fa482c7} /* (23, 10, 20) {real, imag} */,
  {32'h3ed270cf, 32'h4040a3b3} /* (23, 10, 19) {real, imag} */,
  {32'hbfa2cd55, 32'h3ee66ed4} /* (23, 10, 18) {real, imag} */,
  {32'hc00b290a, 32'hbf837aee} /* (23, 10, 17) {real, imag} */,
  {32'hbf793473, 32'h3f8abef4} /* (23, 10, 16) {real, imag} */,
  {32'hbfec87db, 32'h3e1d0a08} /* (23, 10, 15) {real, imag} */,
  {32'hbef4dd7c, 32'hbfc65ae2} /* (23, 10, 14) {real, imag} */,
  {32'h3f29cfad, 32'hc00368d2} /* (23, 10, 13) {real, imag} */,
  {32'h3fba6180, 32'hbf12c936} /* (23, 10, 12) {real, imag} */,
  {32'h3febc550, 32'h3fdbba3c} /* (23, 10, 11) {real, imag} */,
  {32'h3f46c331, 32'hbf0157bf} /* (23, 10, 10) {real, imag} */,
  {32'hbeb9a1fc, 32'hc0293968} /* (23, 10, 9) {real, imag} */,
  {32'hbf9c5110, 32'hbf5a3eb8} /* (23, 10, 8) {real, imag} */,
  {32'hbf9f428b, 32'hbfec2bfe} /* (23, 10, 7) {real, imag} */,
  {32'hbf796d32, 32'hbf5721db} /* (23, 10, 6) {real, imag} */,
  {32'hbf8e6684, 32'hbf017cb4} /* (23, 10, 5) {real, imag} */,
  {32'hbf55e854, 32'h3e1637e8} /* (23, 10, 4) {real, imag} */,
  {32'h3fa8496b, 32'h3fc45a7c} /* (23, 10, 3) {real, imag} */,
  {32'h40404cee, 32'h3f8b5240} /* (23, 10, 2) {real, imag} */,
  {32'h3f83fb27, 32'h3f7ddbf8} /* (23, 10, 1) {real, imag} */,
  {32'hbf0277df, 32'h3f8e76c6} /* (23, 10, 0) {real, imag} */,
  {32'h3f81c7f7, 32'hbf2f54f5} /* (23, 9, 31) {real, imag} */,
  {32'h3e9c791e, 32'hbf3bfb3f} /* (23, 9, 30) {real, imag} */,
  {32'hbecb7e60, 32'hbdb63c40} /* (23, 9, 29) {real, imag} */,
  {32'hbf27b678, 32'hbf0907aa} /* (23, 9, 28) {real, imag} */,
  {32'hbf818760, 32'hbf23a226} /* (23, 9, 27) {real, imag} */,
  {32'hbf402404, 32'h3ddfbd4c} /* (23, 9, 26) {real, imag} */,
  {32'h3e7e1650, 32'hc0089f2e} /* (23, 9, 25) {real, imag} */,
  {32'h3e63970c, 32'hc045e570} /* (23, 9, 24) {real, imag} */,
  {32'h3f3de571, 32'hc022eda2} /* (23, 9, 23) {real, imag} */,
  {32'h3fd67d13, 32'hc01f655e} /* (23, 9, 22) {real, imag} */,
  {32'h3f5ceb73, 32'hbff13456} /* (23, 9, 21) {real, imag} */,
  {32'h3f87cb32, 32'h3fc1d47e} /* (23, 9, 20) {real, imag} */,
  {32'h3e1a92b0, 32'h4000e6f8} /* (23, 9, 19) {real, imag} */,
  {32'h3e6cc290, 32'h401d5cb2} /* (23, 9, 18) {real, imag} */,
  {32'hbe2f9f38, 32'h4032d80a} /* (23, 9, 17) {real, imag} */,
  {32'h3d774ca0, 32'h3fee9134} /* (23, 9, 16) {real, imag} */,
  {32'hbffd2d78, 32'hbe7b1680} /* (23, 9, 15) {real, imag} */,
  {32'h3fbf0b22, 32'hbfc53423} /* (23, 9, 14) {real, imag} */,
  {32'h3fdd933d, 32'hc01a84d5} /* (23, 9, 13) {real, imag} */,
  {32'h3fbb65e3, 32'hbf898329} /* (23, 9, 12) {real, imag} */,
  {32'h3fca5a08, 32'h4003f5d7} /* (23, 9, 11) {real, imag} */,
  {32'h3f933fcf, 32'hbf8816f5} /* (23, 9, 10) {real, imag} */,
  {32'hbf120564, 32'hc034ef24} /* (23, 9, 9) {real, imag} */,
  {32'hbf1df328, 32'hbfb6713d} /* (23, 9, 8) {real, imag} */,
  {32'hbf4ca7c8, 32'hc0046b04} /* (23, 9, 7) {real, imag} */,
  {32'hbfa36ee4, 32'h3f848de4} /* (23, 9, 6) {real, imag} */,
  {32'hbfeeb54c, 32'h3e9fe661} /* (23, 9, 5) {real, imag} */,
  {32'hbf784078, 32'hbf2f0690} /* (23, 9, 4) {real, imag} */,
  {32'h3fc6ee2e, 32'hbeed7998} /* (23, 9, 3) {real, imag} */,
  {32'h400097d9, 32'hbfb90464} /* (23, 9, 2) {real, imag} */,
  {32'hbe8c3390, 32'hbe91d37b} /* (23, 9, 1) {real, imag} */,
  {32'h3cf7d3e0, 32'hbbcfe100} /* (23, 9, 0) {real, imag} */,
  {32'h3f8d2f7d, 32'h3ecfd9b4} /* (23, 8, 31) {real, imag} */,
  {32'h3f81cbbd, 32'h3d6d4e10} /* (23, 8, 30) {real, imag} */,
  {32'hbfc02bac, 32'h3de19e00} /* (23, 8, 29) {real, imag} */,
  {32'hc0188486, 32'h3e671a22} /* (23, 8, 28) {real, imag} */,
  {32'hbf64ee88, 32'hbece00e8} /* (23, 8, 27) {real, imag} */,
  {32'hbe3572ec, 32'h3ea5002c} /* (23, 8, 26) {real, imag} */,
  {32'h3e341521, 32'hbfdd99d8} /* (23, 8, 25) {real, imag} */,
  {32'h3e1cad00, 32'hc01f2daa} /* (23, 8, 24) {real, imag} */,
  {32'h3fa62682, 32'hbf6b95e6} /* (23, 8, 23) {real, imag} */,
  {32'h40088a7a, 32'hbfacd0ac} /* (23, 8, 22) {real, imag} */,
  {32'h3f0645ea, 32'h3f6a0a10} /* (23, 8, 21) {real, imag} */,
  {32'h3f8abc1a, 32'h40064fdf} /* (23, 8, 20) {real, imag} */,
  {32'hbe43cd88, 32'h3f8519d5} /* (23, 8, 19) {real, imag} */,
  {32'h3e9eac19, 32'h3fe4ed0b} /* (23, 8, 18) {real, imag} */,
  {32'h3edb3542, 32'h402b7344} /* (23, 8, 17) {real, imag} */,
  {32'h3f95dd80, 32'h3e6dc9b0} /* (23, 8, 16) {real, imag} */,
  {32'h3fd61d7d, 32'hbfa6503e} /* (23, 8, 15) {real, imag} */,
  {32'h40012e36, 32'hbfa9b4ba} /* (23, 8, 14) {real, imag} */,
  {32'h3fc5872e, 32'hbfb2113e} /* (23, 8, 13) {real, imag} */,
  {32'h402a67ea, 32'hbfc2fcb3} /* (23, 8, 12) {real, imag} */,
  {32'h3fb5da74, 32'h3fdba218} /* (23, 8, 11) {real, imag} */,
  {32'h3f0a04f2, 32'h3ecd5538} /* (23, 8, 10) {real, imag} */,
  {32'hbea961fc, 32'hbf8d2b54} /* (23, 8, 9) {real, imag} */,
  {32'hbee61e38, 32'hbd142200} /* (23, 8, 8) {real, imag} */,
  {32'hbe776a46, 32'hc00f8d60} /* (23, 8, 7) {real, imag} */,
  {32'hbf589d71, 32'h3eb3d1a2} /* (23, 8, 6) {real, imag} */,
  {32'hbf28db6a, 32'h3e858624} /* (23, 8, 5) {real, imag} */,
  {32'hbecf533a, 32'h3e3176c8} /* (23, 8, 4) {real, imag} */,
  {32'h3f635b7c, 32'hbf1a9174} /* (23, 8, 3) {real, imag} */,
  {32'h3f5b90a6, 32'hc01dad1a} /* (23, 8, 2) {real, imag} */,
  {32'h3f75966a, 32'hbf73891c} /* (23, 8, 1) {real, imag} */,
  {32'h3f8f261b, 32'hbf082e02} /* (23, 8, 0) {real, imag} */,
  {32'h3f575e1f, 32'hbd9eef48} /* (23, 7, 31) {real, imag} */,
  {32'h3f999d82, 32'h3f4f80c4} /* (23, 7, 30) {real, imag} */,
  {32'hbebd9488, 32'h3f901d7f} /* (23, 7, 29) {real, imag} */,
  {32'hbfed9cf5, 32'hbdb75428} /* (23, 7, 28) {real, imag} */,
  {32'hbcd449d8, 32'hbe54fd13} /* (23, 7, 27) {real, imag} */,
  {32'h3ebeb83e, 32'hbea36328} /* (23, 7, 26) {real, imag} */,
  {32'h3e6dff58, 32'hc01e44ea} /* (23, 7, 25) {real, imag} */,
  {32'h3ff60ed0, 32'hc00c0420} /* (23, 7, 24) {real, imag} */,
  {32'h3e3f7e28, 32'h3d904a20} /* (23, 7, 23) {real, imag} */,
  {32'h3f42f122, 32'hbfa34ab2} /* (23, 7, 22) {real, imag} */,
  {32'h3f0e230a, 32'h3e48ff60} /* (23, 7, 21) {real, imag} */,
  {32'h3e996850, 32'h3fc7e818} /* (23, 7, 20) {real, imag} */,
  {32'hbdd744a8, 32'hbeae5cbe} /* (23, 7, 19) {real, imag} */,
  {32'h3f35c454, 32'h3e0a9380} /* (23, 7, 18) {real, imag} */,
  {32'h3f2227d5, 32'h3fe9bcf5} /* (23, 7, 17) {real, imag} */,
  {32'h3ddd3c10, 32'hbe8928c0} /* (23, 7, 16) {real, imag} */,
  {32'h3fd76d52, 32'h3f96284a} /* (23, 7, 15) {real, imag} */,
  {32'h3fcf5f08, 32'h3f8f8f44} /* (23, 7, 14) {real, imag} */,
  {32'h3fbcbe71, 32'h3eceb1fd} /* (23, 7, 13) {real, imag} */,
  {32'h40209d7c, 32'hbf36fdc0} /* (23, 7, 12) {real, imag} */,
  {32'h3fbbaa86, 32'h3fa6be38} /* (23, 7, 11) {real, imag} */,
  {32'h3f04625e, 32'h3fb7f2ef} /* (23, 7, 10) {real, imag} */,
  {32'h3da977c8, 32'h3fd83258} /* (23, 7, 9) {real, imag} */,
  {32'h3e6259a6, 32'h3fb4ee04} /* (23, 7, 8) {real, imag} */,
  {32'h3df8c350, 32'hbff13eee} /* (23, 7, 7) {real, imag} */,
  {32'hbdd29e84, 32'hbfdbab22} /* (23, 7, 6) {real, imag} */,
  {32'hbfed0bc5, 32'hbf721c82} /* (23, 7, 5) {real, imag} */,
  {32'hbf3ac94c, 32'hbe0f60ba} /* (23, 7, 4) {real, imag} */,
  {32'h3fa1b391, 32'h3f661374} /* (23, 7, 3) {real, imag} */,
  {32'hbf182cfd, 32'hbf619ee8} /* (23, 7, 2) {real, imag} */,
  {32'hbeff9bcc, 32'hbe8b99f8} /* (23, 7, 1) {real, imag} */,
  {32'h3e8851b4, 32'h3e4ab788} /* (23, 7, 0) {real, imag} */,
  {32'h3f5cdc5b, 32'hbef71858} /* (23, 6, 31) {real, imag} */,
  {32'h3f56ce70, 32'h3f4c7ef0} /* (23, 6, 30) {real, imag} */,
  {32'h3e95a0be, 32'h3cdd7e40} /* (23, 6, 29) {real, imag} */,
  {32'h3e580a00, 32'hbed51464} /* (23, 6, 28) {real, imag} */,
  {32'h3ffdbb07, 32'hbe441950} /* (23, 6, 27) {real, imag} */,
  {32'h3feb3344, 32'hbf6c8dcf} /* (23, 6, 26) {real, imag} */,
  {32'hbfb85e19, 32'hbfa96f0a} /* (23, 6, 25) {real, imag} */,
  {32'hbf6c1ec0, 32'h3e8eca5b} /* (23, 6, 24) {real, imag} */,
  {32'hbf660a68, 32'h3f8d4bad} /* (23, 6, 23) {real, imag} */,
  {32'hbf2efd64, 32'hbfc47d32} /* (23, 6, 22) {real, imag} */,
  {32'hbf6a7d5a, 32'hbf823952} /* (23, 6, 21) {real, imag} */,
  {32'hbf48b698, 32'h3f7e6860} /* (23, 6, 20) {real, imag} */,
  {32'hbe1f909c, 32'hbec59a7c} /* (23, 6, 19) {real, imag} */,
  {32'h3f8965dd, 32'h3e210a78} /* (23, 6, 18) {real, imag} */,
  {32'h3f364372, 32'h3f0aab6c} /* (23, 6, 17) {real, imag} */,
  {32'hbf58ce54, 32'hbfcd6e76} /* (23, 6, 16) {real, imag} */,
  {32'h3f1a0811, 32'hbedf6337} /* (23, 6, 15) {real, imag} */,
  {32'h3f64aefa, 32'h3e89099a} /* (23, 6, 14) {real, imag} */,
  {32'h3f334894, 32'h3e818df0} /* (23, 6, 13) {real, imag} */,
  {32'hbf3f0f5f, 32'h3dd4a480} /* (23, 6, 12) {real, imag} */,
  {32'hbfc0b339, 32'h3e49e7f0} /* (23, 6, 11) {real, imag} */,
  {32'hbf8717a6, 32'h3f227795} /* (23, 6, 10) {real, imag} */,
  {32'hbf3b92ff, 32'h3faba607} /* (23, 6, 9) {real, imag} */,
  {32'h3facb9c5, 32'h3ff12a53} /* (23, 6, 8) {real, imag} */,
  {32'h3e2c9186, 32'hbf51007a} /* (23, 6, 7) {real, imag} */,
  {32'hc0020d70, 32'hc02e8ad7} /* (23, 6, 6) {real, imag} */,
  {32'hc02e1d10, 32'hc0149c4b} /* (23, 6, 5) {real, imag} */,
  {32'h3ef4ab9c, 32'hc005c05a} /* (23, 6, 4) {real, imag} */,
  {32'h3f0dda9e, 32'hbf280a3c} /* (23, 6, 3) {real, imag} */,
  {32'hbf7ec21c, 32'h3f6ffb4e} /* (23, 6, 2) {real, imag} */,
  {32'h3f0ee8c2, 32'hbe80bc18} /* (23, 6, 1) {real, imag} */,
  {32'h3f49c3f8, 32'hbea0eeb8} /* (23, 6, 0) {real, imag} */,
  {32'h3e17bf40, 32'hbf4e8baf} /* (23, 5, 31) {real, imag} */,
  {32'h3e984a1c, 32'hbe13f5fa} /* (23, 5, 30) {real, imag} */,
  {32'hbf23dd1c, 32'h3e2f73f0} /* (23, 5, 29) {real, imag} */,
  {32'hbf7fcdee, 32'hbf25ebf7} /* (23, 5, 28) {real, imag} */,
  {32'h3f6810a0, 32'hbecd7564} /* (23, 5, 27) {real, imag} */,
  {32'h3df1ec88, 32'hbf6feb4a} /* (23, 5, 26) {real, imag} */,
  {32'hbfd0fce2, 32'hbf8a2300} /* (23, 5, 25) {real, imag} */,
  {32'hbf6cdb41, 32'hbe0d4d28} /* (23, 5, 24) {real, imag} */,
  {32'hbedf50c4, 32'hbf803b08} /* (23, 5, 23) {real, imag} */,
  {32'hbe8c2c70, 32'hbfe9c667} /* (23, 5, 22) {real, imag} */,
  {32'hbf8ffee0, 32'hbe6b7330} /* (23, 5, 21) {real, imag} */,
  {32'hbff27c16, 32'h3fc445ff} /* (23, 5, 20) {real, imag} */,
  {32'hbf761fc2, 32'h3ec79cf0} /* (23, 5, 19) {real, imag} */,
  {32'h3e4abc58, 32'hbe981928} /* (23, 5, 18) {real, imag} */,
  {32'hbfa66ef6, 32'hbfb5855f} /* (23, 5, 17) {real, imag} */,
  {32'hbeae398d, 32'hc03c42d0} /* (23, 5, 16) {real, imag} */,
  {32'h3ece5776, 32'hc031e159} /* (23, 5, 15) {real, imag} */,
  {32'hbe1760b4, 32'hbf3f9ab5} /* (23, 5, 14) {real, imag} */,
  {32'hbde756a0, 32'hbf4ae5a8} /* (23, 5, 13) {real, imag} */,
  {32'hbf9645a0, 32'h3e144b1c} /* (23, 5, 12) {real, imag} */,
  {32'hbfb45c06, 32'hbe395dc8} /* (23, 5, 11) {real, imag} */,
  {32'hbf44a07c, 32'h3d7379d0} /* (23, 5, 10) {real, imag} */,
  {32'hbf9c45e0, 32'h3f9fb46c} /* (23, 5, 9) {real, imag} */,
  {32'h3f6a17f6, 32'h400509a8} /* (23, 5, 8) {real, imag} */,
  {32'h3f885820, 32'h3f4060eb} /* (23, 5, 7) {real, imag} */,
  {32'hc00c16ac, 32'hbf90049b} /* (23, 5, 6) {real, imag} */,
  {32'hc0106d4b, 32'hbf7ac281} /* (23, 5, 5) {real, imag} */,
  {32'h3f1f5aba, 32'hbdf969f0} /* (23, 5, 4) {real, imag} */,
  {32'h3e74bec0, 32'hbf606488} /* (23, 5, 3) {real, imag} */,
  {32'h3edfc624, 32'hbf8377d8} /* (23, 5, 2) {real, imag} */,
  {32'h3e9d33ff, 32'hbe02fd50} /* (23, 5, 1) {real, imag} */,
  {32'hbe29a19a, 32'h3f7337da} /* (23, 5, 0) {real, imag} */,
  {32'h3f86acbe, 32'hbf88e580} /* (23, 4, 31) {real, imag} */,
  {32'h40017544, 32'h3e79ed16} /* (23, 4, 30) {real, imag} */,
  {32'h3e807222, 32'hbf010f9b} /* (23, 4, 29) {real, imag} */,
  {32'hbfd856e8, 32'hc0032dbe} /* (23, 4, 28) {real, imag} */,
  {32'hbfb90146, 32'hbf452e25} /* (23, 4, 27) {real, imag} */,
  {32'hbe6bd256, 32'h3ef1f2c0} /* (23, 4, 26) {real, imag} */,
  {32'h3ec00a78, 32'hbcb54380} /* (23, 4, 25) {real, imag} */,
  {32'h3d539410, 32'hbfa3f720} /* (23, 4, 24) {real, imag} */,
  {32'hbfa0a426, 32'hbfd42da6} /* (23, 4, 23) {real, imag} */,
  {32'hbf179e13, 32'hbd8485b8} /* (23, 4, 22) {real, imag} */,
  {32'h3e5fdc7c, 32'h3f969fc6} /* (23, 4, 21) {real, imag} */,
  {32'hbe2efb60, 32'h3febb4fe} /* (23, 4, 20) {real, imag} */,
  {32'hbf8d80c6, 32'h3e5ead26} /* (23, 4, 19) {real, imag} */,
  {32'h3e10a508, 32'hbe8429d8} /* (23, 4, 18) {real, imag} */,
  {32'hbd98e0b0, 32'hbfa5ad42} /* (23, 4, 17) {real, imag} */,
  {32'h3f807843, 32'hbfcd43dc} /* (23, 4, 16) {real, imag} */,
  {32'h3fd523cf, 32'hbfaf874c} /* (23, 4, 15) {real, imag} */,
  {32'h3fc53003, 32'hbeaea340} /* (23, 4, 14) {real, imag} */,
  {32'h3f95869e, 32'hbe9d9236} /* (23, 4, 13) {real, imag} */,
  {32'h3fcff4c4, 32'h3eb64290} /* (23, 4, 12) {real, imag} */,
  {32'h3fa18048, 32'h3f870ead} /* (23, 4, 11) {real, imag} */,
  {32'h3f865ed8, 32'h3f268f3e} /* (23, 4, 10) {real, imag} */,
  {32'hbf038cb2, 32'h3f0a351c} /* (23, 4, 9) {real, imag} */,
  {32'hbf370b3c, 32'h3f1dbd06} /* (23, 4, 8) {real, imag} */,
  {32'h3eb35c2e, 32'h3f0016ae} /* (23, 4, 7) {real, imag} */,
  {32'hbecacc78, 32'h3ec21417} /* (23, 4, 6) {real, imag} */,
  {32'hc00f68ef, 32'h3e0df43c} /* (23, 4, 5) {real, imag} */,
  {32'hbfd72227, 32'hbe5dfad0} /* (23, 4, 4) {real, imag} */,
  {32'h3ef273ac, 32'hbfab8ca4} /* (23, 4, 3) {real, imag} */,
  {32'h3f6e7b2b, 32'hbfe11264} /* (23, 4, 2) {real, imag} */,
  {32'hbf30ed41, 32'hbfce2cbd} /* (23, 4, 1) {real, imag} */,
  {32'hbf0a3034, 32'hbf294b11} /* (23, 4, 0) {real, imag} */,
  {32'h3f8fe1bc, 32'hbf02fe2a} /* (23, 3, 31) {real, imag} */,
  {32'h3eda690e, 32'h3fd30d90} /* (23, 3, 30) {real, imag} */,
  {32'hbe99a623, 32'h3fa5c9af} /* (23, 3, 29) {real, imag} */,
  {32'hbf9d5007, 32'hc02bcdf0} /* (23, 3, 28) {real, imag} */,
  {32'hbfc29076, 32'hc0037cac} /* (23, 3, 27) {real, imag} */,
  {32'hbf0f3f8b, 32'h3e416ed0} /* (23, 3, 26) {real, imag} */,
  {32'hbfcdbc2f, 32'hbe93dcca} /* (23, 3, 25) {real, imag} */,
  {32'hbf8c2f9e, 32'hc00d8d7d} /* (23, 3, 24) {real, imag} */,
  {32'hbfad60a5, 32'hc04af5ef} /* (23, 3, 23) {real, imag} */,
  {32'hbfc30f92, 32'hbf2151d8} /* (23, 3, 22) {real, imag} */,
  {32'hbf0e7854, 32'h3ec166f7} /* (23, 3, 21) {real, imag} */,
  {32'h3db83190, 32'h3efda097} /* (23, 3, 20) {real, imag} */,
  {32'hbe948bfe, 32'hbd3acc00} /* (23, 3, 19) {real, imag} */,
  {32'h3f4ca30a, 32'h3f315702} /* (23, 3, 18) {real, imag} */,
  {32'hbd94e8c0, 32'hbf19b534} /* (23, 3, 17) {real, imag} */,
  {32'h3ebd5480, 32'hbf1d668e} /* (23, 3, 16) {real, imag} */,
  {32'h3f33de0e, 32'hbf9a2ff9} /* (23, 3, 15) {real, imag} */,
  {32'h3f3d6772, 32'h3def2b40} /* (23, 3, 14) {real, imag} */,
  {32'h3fa8727e, 32'hbeef92d4} /* (23, 3, 13) {real, imag} */,
  {32'h40396c82, 32'hbf897b30} /* (23, 3, 12) {real, imag} */,
  {32'h40285c72, 32'h3fd6ebc6} /* (23, 3, 11) {real, imag} */,
  {32'h3fb6e96e, 32'h3fc6b2bd} /* (23, 3, 10) {real, imag} */,
  {32'hbceec3c0, 32'h3edeee22} /* (23, 3, 9) {real, imag} */,
  {32'hbe678790, 32'h3e834683} /* (23, 3, 8) {real, imag} */,
  {32'h3f3960c9, 32'h3f3732a6} /* (23, 3, 7) {real, imag} */,
  {32'h3f546cb8, 32'hbd428790} /* (23, 3, 6) {real, imag} */,
  {32'hbee5c86a, 32'h3fb61a3e} /* (23, 3, 5) {real, imag} */,
  {32'hbfe9122a, 32'h3ef2ce48} /* (23, 3, 4) {real, imag} */,
  {32'h3ec98f13, 32'hc009cc38} /* (23, 3, 3) {real, imag} */,
  {32'h3e000c40, 32'hc02fb804} /* (23, 3, 2) {real, imag} */,
  {32'hc0184b5e, 32'hbfe82858} /* (23, 3, 1) {real, imag} */,
  {32'hbf2bdf0e, 32'hbfdbc580} /* (23, 3, 0) {real, imag} */,
  {32'hbe0727f4, 32'h3e0900fe} /* (23, 2, 31) {real, imag} */,
  {32'hbfbc9fba, 32'h3f6dcdc4} /* (23, 2, 30) {real, imag} */,
  {32'hbf1f7b46, 32'h3e8a57e0} /* (23, 2, 29) {real, imag} */,
  {32'h3e6e9ea4, 32'hbfec2c8e} /* (23, 2, 28) {real, imag} */,
  {32'hbf63ab96, 32'hbfc60932} /* (23, 2, 27) {real, imag} */,
  {32'hbf05a08e, 32'h3ee554e0} /* (23, 2, 26) {real, imag} */,
  {32'hbfa613f2, 32'h3f06125c} /* (23, 2, 25) {real, imag} */,
  {32'hbfae6947, 32'hbed50998} /* (23, 2, 24) {real, imag} */,
  {32'h3e1dab3c, 32'hbfe6750e} /* (23, 2, 23) {real, imag} */,
  {32'h3f38f381, 32'hbfdc07cb} /* (23, 2, 22) {real, imag} */,
  {32'h3f02459a, 32'hbe2fb77c} /* (23, 2, 21) {real, imag} */,
  {32'h3e081048, 32'h3e875fc5} /* (23, 2, 20) {real, imag} */,
  {32'hbe04a60a, 32'hbdb214c8} /* (23, 2, 19) {real, imag} */,
  {32'h3f4e2955, 32'h3f875303} /* (23, 2, 18) {real, imag} */,
  {32'h3e1f6832, 32'h3eda4222} /* (23, 2, 17) {real, imag} */,
  {32'hbf8f3355, 32'hbe1894a0} /* (23, 2, 16) {real, imag} */,
  {32'hbd7cfb80, 32'h3ec897d4} /* (23, 2, 15) {real, imag} */,
  {32'hbec43ec0, 32'h3ee657d8} /* (23, 2, 14) {real, imag} */,
  {32'hbf99438d, 32'hbee6437b} /* (23, 2, 13) {real, imag} */,
  {32'h3f7319a0, 32'hbf3b6099} /* (23, 2, 12) {real, imag} */,
  {32'h3fc937d8, 32'hbf18d384} /* (23, 2, 11) {real, imag} */,
  {32'h3fb766ef, 32'h3e1ef5b4} /* (23, 2, 10) {real, imag} */,
  {32'h3dc198d0, 32'h3f8d408e} /* (23, 2, 9) {real, imag} */,
  {32'h3f9bdb22, 32'h3fd6bf5c} /* (23, 2, 8) {real, imag} */,
  {32'h4000e204, 32'h3f9a4b7b} /* (23, 2, 7) {real, imag} */,
  {32'h3fdfad48, 32'hbf42d0b0} /* (23, 2, 6) {real, imag} */,
  {32'hbf80442e, 32'h3eeaa640} /* (23, 2, 5) {real, imag} */,
  {32'hbf0ab8b8, 32'h3fa657aa} /* (23, 2, 4) {real, imag} */,
  {32'h40024096, 32'hbfdab899} /* (23, 2, 3) {real, imag} */,
  {32'hbe83a872, 32'hc02329ae} /* (23, 2, 2) {real, imag} */,
  {32'hbf536b61, 32'hbffe6c4e} /* (23, 2, 1) {real, imag} */,
  {32'h3ef18f36, 32'hbfc7cb10} /* (23, 2, 0) {real, imag} */,
  {32'hbf8ff3b4, 32'hbe97a4c0} /* (23, 1, 31) {real, imag} */,
  {32'hbfd9589b, 32'hbe22b67a} /* (23, 1, 30) {real, imag} */,
  {32'hbf356497, 32'hbebee2e4} /* (23, 1, 29) {real, imag} */,
  {32'h3f994710, 32'hbe2d2c9c} /* (23, 1, 28) {real, imag} */,
  {32'hbd82e0fc, 32'h3f6c0e83} /* (23, 1, 27) {real, imag} */,
  {32'hbcfd7070, 32'h3fb11ef6} /* (23, 1, 26) {real, imag} */,
  {32'hbfbef23b, 32'h3f7a3906} /* (23, 1, 25) {real, imag} */,
  {32'hbf2f9bcf, 32'h3f6a6c64} /* (23, 1, 24) {real, imag} */,
  {32'hbe16c6f4, 32'hbf00777c} /* (23, 1, 23) {real, imag} */,
  {32'hbe2f9e88, 32'hbfbdb0a5} /* (23, 1, 22) {real, imag} */,
  {32'hbf82df42, 32'hbd8d1590} /* (23, 1, 21) {real, imag} */,
  {32'hbf3ce6f3, 32'h3fbe0609} /* (23, 1, 20) {real, imag} */,
  {32'hbf2970d3, 32'h3f24415b} /* (23, 1, 19) {real, imag} */,
  {32'h3e610848, 32'hbedc2118} /* (23, 1, 18) {real, imag} */,
  {32'hbff6d1b2, 32'hbf66e632} /* (23, 1, 17) {real, imag} */,
  {32'hc03a376e, 32'hbf5467da} /* (23, 1, 16) {real, imag} */,
  {32'hbf369605, 32'hbfadd1dc} /* (23, 1, 15) {real, imag} */,
  {32'h3edafa9d, 32'hbfbf23d0} /* (23, 1, 14) {real, imag} */,
  {32'hbf264146, 32'h3f2efacf} /* (23, 1, 13) {real, imag} */,
  {32'hbfb1e61d, 32'hbcdd8900} /* (23, 1, 12) {real, imag} */,
  {32'hbe8b058e, 32'h3caa5480} /* (23, 1, 11) {real, imag} */,
  {32'h3f1014ec, 32'h3f63b6fd} /* (23, 1, 10) {real, imag} */,
  {32'h3e857b9c, 32'h3f40e8c0} /* (23, 1, 9) {real, imag} */,
  {32'h3fb6611c, 32'h3f9094d8} /* (23, 1, 8) {real, imag} */,
  {32'h401c873e, 32'h3f0c0a7a} /* (23, 1, 7) {real, imag} */,
  {32'h40071087, 32'hbfc88fb8} /* (23, 1, 6) {real, imag} */,
  {32'hbf3f69fb, 32'hbf91cd0b} /* (23, 1, 5) {real, imag} */,
  {32'hbe65b558, 32'h3ef9cc50} /* (23, 1, 4) {real, imag} */,
  {32'h3eebf23e, 32'hbf15938c} /* (23, 1, 3) {real, imag} */,
  {32'hbfd387b3, 32'hbef22022} /* (23, 1, 2) {real, imag} */,
  {32'hbf2b1fe0, 32'hbecef488} /* (23, 1, 1) {real, imag} */,
  {32'h3e9898de, 32'hbf19a47d} /* (23, 1, 0) {real, imag} */,
  {32'hbeea2a49, 32'hbf317aa0} /* (23, 0, 31) {real, imag} */,
  {32'hbf097b26, 32'h3eac8147} /* (23, 0, 30) {real, imag} */,
  {32'hbf0527c2, 32'h3f6e6183} /* (23, 0, 29) {real, imag} */,
  {32'h3d768120, 32'h3f070ae0} /* (23, 0, 28) {real, imag} */,
  {32'h3e1903ac, 32'h3e6b4912} /* (23, 0, 27) {real, imag} */,
  {32'hbf127556, 32'h3cec32e0} /* (23, 0, 26) {real, imag} */,
  {32'hbf48dffa, 32'h3e50bc70} /* (23, 0, 25) {real, imag} */,
  {32'hbe84baa8, 32'h3f5c1d35} /* (23, 0, 24) {real, imag} */,
  {32'hbe81fbd8, 32'h3e44ea7a} /* (23, 0, 23) {real, imag} */,
  {32'hbf50e0b2, 32'hbf04c526} /* (23, 0, 22) {real, imag} */,
  {32'hbfc8329e, 32'hbe890908} /* (23, 0, 21) {real, imag} */,
  {32'hbf640eeb, 32'h3e86880a} /* (23, 0, 20) {real, imag} */,
  {32'h3e4f9658, 32'h3f1ad854} /* (23, 0, 19) {real, imag} */,
  {32'h3e0d346b, 32'h3e92d57a} /* (23, 0, 18) {real, imag} */,
  {32'hbfe0bbee, 32'h3eba251c} /* (23, 0, 17) {real, imag} */,
  {32'hbfa3b486, 32'h3e32d448} /* (23, 0, 16) {real, imag} */,
  {32'hbe42c2c6, 32'hbef5f19c} /* (23, 0, 15) {real, imag} */,
  {32'h3f1e8fc6, 32'hbfa7f1fe} /* (23, 0, 14) {real, imag} */,
  {32'h3f8020f3, 32'hbdc08180} /* (23, 0, 13) {real, imag} */,
  {32'hbf54e3d8, 32'h3e8a28bc} /* (23, 0, 12) {real, imag} */,
  {32'hbeed88ae, 32'h3dbf9d5c} /* (23, 0, 11) {real, imag} */,
  {32'h3effe34c, 32'hbd857b28} /* (23, 0, 10) {real, imag} */,
  {32'h3eae5d61, 32'hbf80fd95} /* (23, 0, 9) {real, imag} */,
  {32'h3f4659b1, 32'hbf288530} /* (23, 0, 8) {real, imag} */,
  {32'h3fe2941b, 32'hbe83888e} /* (23, 0, 7) {real, imag} */,
  {32'h3f8eba0f, 32'hbf38852c} /* (23, 0, 6) {real, imag} */,
  {32'h3ec57a8b, 32'hbf114b8f} /* (23, 0, 5) {real, imag} */,
  {32'hbf1768f6, 32'hbd814498} /* (23, 0, 4) {real, imag} */,
  {32'hbee5823a, 32'h3efbb9ec} /* (23, 0, 3) {real, imag} */,
  {32'hbf1dba37, 32'h3f6ac649} /* (23, 0, 2) {real, imag} */,
  {32'hbe8d1f54, 32'hbf1d44a4} /* (23, 0, 1) {real, imag} */,
  {32'h3eef2767, 32'hbf1c906d} /* (23, 0, 0) {real, imag} */,
  {32'hbe06886c, 32'h3e1b216a} /* (22, 31, 31) {real, imag} */,
  {32'h3ef93112, 32'h3c886a00} /* (22, 31, 30) {real, imag} */,
  {32'hbe99ce58, 32'h3eb05162} /* (22, 31, 29) {real, imag} */,
  {32'hbf611ba6, 32'hbe797814} /* (22, 31, 28) {real, imag} */,
  {32'hbeefa240, 32'hbe7d66ac} /* (22, 31, 27) {real, imag} */,
  {32'hbf12839c, 32'hbf741a86} /* (22, 31, 26) {real, imag} */,
  {32'hbf9c745f, 32'hbefe16ca} /* (22, 31, 25) {real, imag} */,
  {32'hbf789da6, 32'hbefa42c8} /* (22, 31, 24) {real, imag} */,
  {32'hbf847a88, 32'hbf837aa0} /* (22, 31, 23) {real, imag} */,
  {32'hbef754d4, 32'hbfa6e567} /* (22, 31, 22) {real, imag} */,
  {32'hbe505964, 32'hbf73c30c} /* (22, 31, 21) {real, imag} */,
  {32'hbe00c620, 32'hbdf5bb64} /* (22, 31, 20) {real, imag} */,
  {32'hbd3bfb60, 32'h3ebc4d64} /* (22, 31, 19) {real, imag} */,
  {32'h3eb273c8, 32'h3e9292dc} /* (22, 31, 18) {real, imag} */,
  {32'h3f3b357a, 32'h3f8d39cb} /* (22, 31, 17) {real, imag} */,
  {32'h3e7839fe, 32'h3e3cccfa} /* (22, 31, 16) {real, imag} */,
  {32'h3d87ec28, 32'h3e984f04} /* (22, 31, 15) {real, imag} */,
  {32'h3f339e7e, 32'h3f227036} /* (22, 31, 14) {real, imag} */,
  {32'h3f559fa2, 32'h3e352a40} /* (22, 31, 13) {real, imag} */,
  {32'h3f9d65da, 32'h3e8852ec} /* (22, 31, 12) {real, imag} */,
  {32'h3faff7df, 32'hbee4d16d} /* (22, 31, 11) {real, imag} */,
  {32'hbe997360, 32'hbf61945e} /* (22, 31, 10) {real, imag} */,
  {32'hbe0c6520, 32'hbeb3c514} /* (22, 31, 9) {real, imag} */,
  {32'hbf0fe6c2, 32'hbf205aa8} /* (22, 31, 8) {real, imag} */,
  {32'h3ed077b4, 32'hbe801264} /* (22, 31, 7) {real, imag} */,
  {32'h3f94eb54, 32'hbea6a28c} /* (22, 31, 6) {real, imag} */,
  {32'hbeb467c8, 32'hbf8e7ee7} /* (22, 31, 5) {real, imag} */,
  {32'hbf8cfba8, 32'hbf92d2c2} /* (22, 31, 4) {real, imag} */,
  {32'hbf0063d1, 32'hbed0e05a} /* (22, 31, 3) {real, imag} */,
  {32'hbf50b148, 32'h3f4de2d9} /* (22, 31, 2) {real, imag} */,
  {32'hbecdad80, 32'h401498da} /* (22, 31, 1) {real, imag} */,
  {32'hbec4eddc, 32'h3f8afc8c} /* (22, 31, 0) {real, imag} */,
  {32'h3edd3e28, 32'h3ddd8a24} /* (22, 30, 31) {real, imag} */,
  {32'h3fd16a9e, 32'hbe0b0960} /* (22, 30, 30) {real, imag} */,
  {32'h3f852e3f, 32'h3de1f0b0} /* (22, 30, 29) {real, imag} */,
  {32'hbf17e49a, 32'hbf270d34} /* (22, 30, 28) {real, imag} */,
  {32'hbfb4c563, 32'hbf66e4ea} /* (22, 30, 27) {real, imag} */,
  {32'hbfc63e3c, 32'h3ea858f0} /* (22, 30, 26) {real, imag} */,
  {32'hbfe88b86, 32'h3e7298f0} /* (22, 30, 25) {real, imag} */,
  {32'hc047964e, 32'hbeb09d58} /* (22, 30, 24) {real, imag} */,
  {32'hc015fb71, 32'hbf277254} /* (22, 30, 23) {real, imag} */,
  {32'h3f609d12, 32'hbfed428a} /* (22, 30, 22) {real, imag} */,
  {32'hbfa217cb, 32'hbfcacc7e} /* (22, 30, 21) {real, imag} */,
  {32'hbfe8f804, 32'hbf870119} /* (22, 30, 20) {real, imag} */,
  {32'h3e1556f4, 32'hbd3c5bc0} /* (22, 30, 19) {real, imag} */,
  {32'h3f93c5f2, 32'h3f06130e} /* (22, 30, 18) {real, imag} */,
  {32'h3f4c1956, 32'h3f9bb6fb} /* (22, 30, 17) {real, imag} */,
  {32'h3f8e0ace, 32'h3f920fb6} /* (22, 30, 16) {real, imag} */,
  {32'h3f126311, 32'h3dabb250} /* (22, 30, 15) {real, imag} */,
  {32'h3e514be0, 32'hbf4e509a} /* (22, 30, 14) {real, imag} */,
  {32'h3f688750, 32'hbfc7ef71} /* (22, 30, 13) {real, imag} */,
  {32'h3fde2d3a, 32'hbf3e63ae} /* (22, 30, 12) {real, imag} */,
  {32'h3f306906, 32'hbf1163e0} /* (22, 30, 11) {real, imag} */,
  {32'hbf614853, 32'hbf852e9c} /* (22, 30, 10) {real, imag} */,
  {32'hbf398d37, 32'hbe947534} /* (22, 30, 9) {real, imag} */,
  {32'hbfa359a4, 32'hbf76999a} /* (22, 30, 8) {real, imag} */,
  {32'hbf73ea2e, 32'hbfd144fd} /* (22, 30, 7) {real, imag} */,
  {32'h3ffb32cc, 32'hbf17b33e} /* (22, 30, 6) {real, imag} */,
  {32'hbf445854, 32'hbfbe9728} /* (22, 30, 5) {real, imag} */,
  {32'hbfeb435f, 32'hbf8b089c} /* (22, 30, 4) {real, imag} */,
  {32'hbf5889f7, 32'hbf933029} /* (22, 30, 3) {real, imag} */,
  {32'hbf1d97ac, 32'h3f7d8398} /* (22, 30, 2) {real, imag} */,
  {32'hbf24d2c3, 32'h3fee1e86} /* (22, 30, 1) {real, imag} */,
  {32'hbee37778, 32'h3e5d74f0} /* (22, 30, 0) {real, imag} */,
  {32'h3fb8809b, 32'hbea70f8e} /* (22, 29, 31) {real, imag} */,
  {32'h401f9980, 32'hbed61f70} /* (22, 29, 30) {real, imag} */,
  {32'h3f83a23d, 32'hbee81044} /* (22, 29, 29) {real, imag} */,
  {32'hbfbeaab2, 32'hbf5ada36} /* (22, 29, 28) {real, imag} */,
  {32'hbf9a4190, 32'h3ef575ba} /* (22, 29, 27) {real, imag} */,
  {32'h3f436938, 32'h3ebfab90} /* (22, 29, 26) {real, imag} */,
  {32'hbefd67a2, 32'hbf646a3d} /* (22, 29, 25) {real, imag} */,
  {32'hc012ac41, 32'hbf95d396} /* (22, 29, 24) {real, imag} */,
  {32'hbfebf0f6, 32'hbfef190e} /* (22, 29, 23) {real, imag} */,
  {32'h3e49cabc, 32'hc045d098} /* (22, 29, 22) {real, imag} */,
  {32'hbec9adef, 32'hbf92a250} /* (22, 29, 21) {real, imag} */,
  {32'h3e73c884, 32'hbfb91b80} /* (22, 29, 20) {real, imag} */,
  {32'h3fb859f0, 32'hbf48b7da} /* (22, 29, 19) {real, imag} */,
  {32'h3fc1b03a, 32'hbf93ed11} /* (22, 29, 18) {real, imag} */,
  {32'h3f82ac2e, 32'h3ece8542} /* (22, 29, 17) {real, imag} */,
  {32'h3f694858, 32'h3f9f3438} /* (22, 29, 16) {real, imag} */,
  {32'h3de68ec0, 32'h3f25f7a4} /* (22, 29, 15) {real, imag} */,
  {32'h3ee42570, 32'h3e0ddbc0} /* (22, 29, 14) {real, imag} */,
  {32'h3ec48820, 32'hbdca5100} /* (22, 29, 13) {real, imag} */,
  {32'h3fd71a6c, 32'hbf9957f5} /* (22, 29, 12) {real, imag} */,
  {32'h3fed428e, 32'hbf19ee4a} /* (22, 29, 11) {real, imag} */,
  {32'h3f6acd6a, 32'h3e382fbc} /* (22, 29, 10) {real, imag} */,
  {32'h3e34b4e8, 32'h3e7f6c28} /* (22, 29, 9) {real, imag} */,
  {32'hbf3a3f98, 32'hbfa45be1} /* (22, 29, 8) {real, imag} */,
  {32'h3e150e10, 32'hbff4aefc} /* (22, 29, 7) {real, imag} */,
  {32'h3f9b6ad9, 32'hbf506c28} /* (22, 29, 6) {real, imag} */,
  {32'hbe937510, 32'hbf20850f} /* (22, 29, 5) {real, imag} */,
  {32'hbea9bb98, 32'hbf9415c5} /* (22, 29, 4) {real, imag} */,
  {32'hbf2268a0, 32'h3e85f264} /* (22, 29, 3) {real, imag} */,
  {32'hbfaf6f56, 32'h3fa124aa} /* (22, 29, 2) {real, imag} */,
  {32'hbfd5227e, 32'h3f7fd55b} /* (22, 29, 1) {real, imag} */,
  {32'hbe6c70ac, 32'hbe52cf34} /* (22, 29, 0) {real, imag} */,
  {32'h3f1f909e, 32'hbf4c2f68} /* (22, 28, 31) {real, imag} */,
  {32'h3e96f8cf, 32'hbf9c986d} /* (22, 28, 30) {real, imag} */,
  {32'hbee7acc0, 32'hbf1dff07} /* (22, 28, 29) {real, imag} */,
  {32'hbf275e7f, 32'h3f268ac8} /* (22, 28, 28) {real, imag} */,
  {32'hbe7690e0, 32'h3fe8ef56} /* (22, 28, 27) {real, imag} */,
  {32'hbedad990, 32'h3eea505c} /* (22, 28, 26) {real, imag} */,
  {32'hbf99627b, 32'hbf88cd2c} /* (22, 28, 25) {real, imag} */,
  {32'hbf5ba63a, 32'hbfb56748} /* (22, 28, 24) {real, imag} */,
  {32'hbf006ad8, 32'hc0046836} /* (22, 28, 23) {real, imag} */,
  {32'h3f3d09b8, 32'hbfe1399f} /* (22, 28, 22) {real, imag} */,
  {32'h3f4b4cd4, 32'h3ebd5aba} /* (22, 28, 21) {real, imag} */,
  {32'h4010f6da, 32'h3f516e3f} /* (22, 28, 20) {real, imag} */,
  {32'h3fcc3be0, 32'h3ea04480} /* (22, 28, 19) {real, imag} */,
  {32'h3f88e23a, 32'hbff49758} /* (22, 28, 18) {real, imag} */,
  {32'h3ed25d06, 32'hbf18335a} /* (22, 28, 17) {real, imag} */,
  {32'h3ec47426, 32'hbd582280} /* (22, 28, 16) {real, imag} */,
  {32'hbf18c8dc, 32'h3c61ed80} /* (22, 28, 15) {real, imag} */,
  {32'h3f5abc90, 32'hbe8e4aec} /* (22, 28, 14) {real, imag} */,
  {32'h3f0803e0, 32'h3e4bfae8} /* (22, 28, 13) {real, imag} */,
  {32'hbda5baf0, 32'h3f20f286} /* (22, 28, 12) {real, imag} */,
  {32'h3ca79840, 32'h3f0c25bf} /* (22, 28, 11) {real, imag} */,
  {32'h3efe5b6c, 32'hbf522319} /* (22, 28, 10) {real, imag} */,
  {32'h3db97810, 32'hbea4c878} /* (22, 28, 9) {real, imag} */,
  {32'h3c0db6c0, 32'hbfd9640a} /* (22, 28, 8) {real, imag} */,
  {32'h404d3c63, 32'hbe5b1658} /* (22, 28, 7) {real, imag} */,
  {32'h3fa9121a, 32'h3ef9716c} /* (22, 28, 6) {real, imag} */,
  {32'h3dd259c8, 32'h3efa16d0} /* (22, 28, 5) {real, imag} */,
  {32'h3ec91960, 32'hbf3c0e3c} /* (22, 28, 4) {real, imag} */,
  {32'hbea29130, 32'hbf255f8e} /* (22, 28, 3) {real, imag} */,
  {32'hbfcc0cae, 32'hbe4ac490} /* (22, 28, 2) {real, imag} */,
  {32'hbf35c139, 32'h3eeb1602} /* (22, 28, 1) {real, imag} */,
  {32'h3f98e359, 32'h3efb63a6} /* (22, 28, 0) {real, imag} */,
  {32'hbdf44ff8, 32'hbf2ef359} /* (22, 27, 31) {real, imag} */,
  {32'hbf8e84e3, 32'hc03a2bdf} /* (22, 27, 30) {real, imag} */,
  {32'hbf6a909d, 32'hc0067089} /* (22, 27, 29) {real, imag} */,
  {32'hbc9c1220, 32'hbee3650c} /* (22, 27, 28) {real, imag} */,
  {32'h3fa541b4, 32'h4004ea2a} /* (22, 27, 27) {real, imag} */,
  {32'hbe6be170, 32'h3fd6d6b7} /* (22, 27, 26) {real, imag} */,
  {32'hbe153520, 32'hbda37360} /* (22, 27, 25) {real, imag} */,
  {32'h3f9ecbe6, 32'hbebf9ae8} /* (22, 27, 24) {real, imag} */,
  {32'h3eebcf88, 32'hbf68fb2e} /* (22, 27, 23) {real, imag} */,
  {32'h3f641a3d, 32'hbf076c61} /* (22, 27, 22) {real, imag} */,
  {32'hbcf96b80, 32'hbed971be} /* (22, 27, 21) {real, imag} */,
  {32'h3edbd4d8, 32'h3f8a585e} /* (22, 27, 20) {real, imag} */,
  {32'h3dc1b8a0, 32'h3ef9e774} /* (22, 27, 19) {real, imag} */,
  {32'hbd4dd740, 32'h3e89949e} /* (22, 27, 18) {real, imag} */,
  {32'h3e990828, 32'hbe9b425c} /* (22, 27, 17) {real, imag} */,
  {32'h3e19e080, 32'h3e887a0a} /* (22, 27, 16) {real, imag} */,
  {32'h3e846b74, 32'h3f30505e} /* (22, 27, 15) {real, imag} */,
  {32'h3f72d356, 32'hbf48c316} /* (22, 27, 14) {real, imag} */,
  {32'hbed25ac4, 32'hbf15f1ac} /* (22, 27, 13) {real, imag} */,
  {32'hbf979700, 32'h3f588c10} /* (22, 27, 12) {real, imag} */,
  {32'hbd1ea500, 32'h3ec36796} /* (22, 27, 11) {real, imag} */,
  {32'h3d4ea480, 32'hbf0e9e38} /* (22, 27, 10) {real, imag} */,
  {32'hbfed75c1, 32'h3f3ee720} /* (22, 27, 9) {real, imag} */,
  {32'hbf709700, 32'hbec0bbf8} /* (22, 27, 8) {real, imag} */,
  {32'h3f843c95, 32'hbe46a438} /* (22, 27, 7) {real, imag} */,
  {32'h3f0eb9a5, 32'hbeed0f24} /* (22, 27, 6) {real, imag} */,
  {32'h3eb442f0, 32'hbe8868aa} /* (22, 27, 5) {real, imag} */,
  {32'hbf5f5a5a, 32'h3f83711a} /* (22, 27, 4) {real, imag} */,
  {32'h3f04e633, 32'h3e976c84} /* (22, 27, 3) {real, imag} */,
  {32'h3f0bbb24, 32'hbf5683a0} /* (22, 27, 2) {real, imag} */,
  {32'h3e035998, 32'hbd94ec50} /* (22, 27, 1) {real, imag} */,
  {32'h3f685101, 32'h3f1ccce7} /* (22, 27, 0) {real, imag} */,
  {32'hbecbb616, 32'hbf2b311b} /* (22, 26, 31) {real, imag} */,
  {32'hbf4a587e, 32'hbfc79628} /* (22, 26, 30) {real, imag} */,
  {32'hbebb36b6, 32'hbeec42a8} /* (22, 26, 29) {real, imag} */,
  {32'hbf8cf255, 32'hbeaee868} /* (22, 26, 28) {real, imag} */,
  {32'hbe72e107, 32'h3f505ba8} /* (22, 26, 27) {real, imag} */,
  {32'h3ebb9964, 32'hbee9fb0c} /* (22, 26, 26) {real, imag} */,
  {32'h3f08590e, 32'h3f1f0752} /* (22, 26, 25) {real, imag} */,
  {32'h3f4e292c, 32'h3f46d9d8} /* (22, 26, 24) {real, imag} */,
  {32'hbef45232, 32'hbf77a346} /* (22, 26, 23) {real, imag} */,
  {32'hbf2d3ba2, 32'hbfc0d0a8} /* (22, 26, 22) {real, imag} */,
  {32'h3e1d99a4, 32'hbf9da56c} /* (22, 26, 21) {real, imag} */,
  {32'h3e9d2b4c, 32'h3da5c3f8} /* (22, 26, 20) {real, imag} */,
  {32'hbebcfc38, 32'h3e567608} /* (22, 26, 19) {real, imag} */,
  {32'hbc930040, 32'h3f90cb90} /* (22, 26, 18) {real, imag} */,
  {32'h3ec1da6c, 32'h3f103fe5} /* (22, 26, 17) {real, imag} */,
  {32'hbebda5b2, 32'hbd9966e8} /* (22, 26, 16) {real, imag} */,
  {32'h3fb33b76, 32'h3eeacbe0} /* (22, 26, 15) {real, imag} */,
  {32'h3f924d74, 32'hbf7055b6} /* (22, 26, 14) {real, imag} */,
  {32'h3ec9aac0, 32'hbf94a731} /* (22, 26, 13) {real, imag} */,
  {32'hbf595f28, 32'hbfb59f32} /* (22, 26, 12) {real, imag} */,
  {32'h3fc79aeb, 32'h3d4291d0} /* (22, 26, 11) {real, imag} */,
  {32'h3fc5b0a1, 32'hbf8f165d} /* (22, 26, 10) {real, imag} */,
  {32'hbf874572, 32'hbf4427ca} /* (22, 26, 9) {real, imag} */,
  {32'hbff2bd54, 32'hbf07f09e} /* (22, 26, 8) {real, imag} */,
  {32'hbf930daf, 32'h3f1667d2} /* (22, 26, 7) {real, imag} */,
  {32'hbef3bd80, 32'h3c214300} /* (22, 26, 6) {real, imag} */,
  {32'h3ee056e0, 32'h3ef0b7ea} /* (22, 26, 5) {real, imag} */,
  {32'hbe8d140e, 32'h3e59d4f4} /* (22, 26, 4) {real, imag} */,
  {32'h3e4c6b44, 32'h3df6ef30} /* (22, 26, 3) {real, imag} */,
  {32'hbf8d08c9, 32'hbecde140} /* (22, 26, 2) {real, imag} */,
  {32'hbfe26b88, 32'hbf342e20} /* (22, 26, 1) {real, imag} */,
  {32'hbeeb8d12, 32'hbea47bdc} /* (22, 26, 0) {real, imag} */,
  {32'h3d1e58e0, 32'hbf41d3a4} /* (22, 25, 31) {real, imag} */,
  {32'hbfa3c328, 32'hbfd49c16} /* (22, 25, 30) {real, imag} */,
  {32'hbead19b8, 32'hbec1a88a} /* (22, 25, 29) {real, imag} */,
  {32'hbf980262, 32'hbf445d09} /* (22, 25, 28) {real, imag} */,
  {32'hbf2d106e, 32'h3f931818} /* (22, 25, 27) {real, imag} */,
  {32'h3f3166ef, 32'h3ed4c310} /* (22, 25, 26) {real, imag} */,
  {32'h3f4703fc, 32'hbd3b3540} /* (22, 25, 25) {real, imag} */,
  {32'hbe4c294c, 32'h3f9462be} /* (22, 25, 24) {real, imag} */,
  {32'hbfe45471, 32'h3e269b84} /* (22, 25, 23) {real, imag} */,
  {32'hbfebfc01, 32'hbf2f9418} /* (22, 25, 22) {real, imag} */,
  {32'h3f1a9b12, 32'hbe0f0e5e} /* (22, 25, 21) {real, imag} */,
  {32'h3f7ee846, 32'h3f49ef0e} /* (22, 25, 20) {real, imag} */,
  {32'h3f1af6f0, 32'hbf3d66dc} /* (22, 25, 19) {real, imag} */,
  {32'h3f156310, 32'hbe7734f8} /* (22, 25, 18) {real, imag} */,
  {32'h3f648860, 32'hbe1784c8} /* (22, 25, 17) {real, imag} */,
  {32'h3f902d8f, 32'hbe50fac0} /* (22, 25, 16) {real, imag} */,
  {32'h3f49b838, 32'hbeb92dca} /* (22, 25, 15) {real, imag} */,
  {32'h3e92e780, 32'hc0165adc} /* (22, 25, 14) {real, imag} */,
  {32'h3f8b8cf0, 32'hbf868485} /* (22, 25, 13) {real, imag} */,
  {32'h3f0d7d80, 32'hbface843} /* (22, 25, 12) {real, imag} */,
  {32'hbedf1774, 32'hbd87a890} /* (22, 25, 11) {real, imag} */,
  {32'h3e8d5029, 32'hbfa231e4} /* (22, 25, 10) {real, imag} */,
  {32'hbf223ece, 32'hbf5ac092} /* (22, 25, 9) {real, imag} */,
  {32'hbfca3bba, 32'h3f06cf34} /* (22, 25, 8) {real, imag} */,
  {32'hbf9647e7, 32'h3f30836e} /* (22, 25, 7) {real, imag} */,
  {32'hbf1ab5eb, 32'hbf5eb4c6} /* (22, 25, 6) {real, imag} */,
  {32'hbec8d0de, 32'hbf947c34} /* (22, 25, 5) {real, imag} */,
  {32'hbf0c824a, 32'hbe77ba88} /* (22, 25, 4) {real, imag} */,
  {32'hbeecac98, 32'hbe973034} /* (22, 25, 3) {real, imag} */,
  {32'hbfafe65c, 32'hbf81c7fb} /* (22, 25, 2) {real, imag} */,
  {32'hbfebd7e9, 32'hbfcc4652} /* (22, 25, 1) {real, imag} */,
  {32'h3ee0010c, 32'hbf927d66} /* (22, 25, 0) {real, imag} */,
  {32'hbf56a6da, 32'h3d1440f0} /* (22, 24, 31) {real, imag} */,
  {32'hc0164842, 32'hbfd81505} /* (22, 24, 30) {real, imag} */,
  {32'hbfc6a3df, 32'hbf405b6c} /* (22, 24, 29) {real, imag} */,
  {32'hc02252a5, 32'hbe37f718} /* (22, 24, 28) {real, imag} */,
  {32'hbfc290eb, 32'h3996b000} /* (22, 24, 27) {real, imag} */,
  {32'h3f5d9910, 32'hbe814edc} /* (22, 24, 26) {real, imag} */,
  {32'h3f1a7e4d, 32'h3ec67df0} /* (22, 24, 25) {real, imag} */,
  {32'hbe17c304, 32'h3f18b7a6} /* (22, 24, 24) {real, imag} */,
  {32'hc035813a, 32'h3e9bacd0} /* (22, 24, 23) {real, imag} */,
  {32'hc0142716, 32'h3f91d10b} /* (22, 24, 22) {real, imag} */,
  {32'hbdb45368, 32'h3cd2bb20} /* (22, 24, 21) {real, imag} */,
  {32'hbe02a358, 32'h3ec8f850} /* (22, 24, 20) {real, imag} */,
  {32'h3f4d0602, 32'hbf46f9d4} /* (22, 24, 19) {real, imag} */,
  {32'h3f94556f, 32'hbff26b7a} /* (22, 24, 18) {real, imag} */,
  {32'h3f6d7993, 32'hbf261f9e} /* (22, 24, 17) {real, imag} */,
  {32'h3f0e5720, 32'h3e99953c} /* (22, 24, 16) {real, imag} */,
  {32'h3fe0568c, 32'h3f647acd} /* (22, 24, 15) {real, imag} */,
  {32'h4019dc94, 32'h3f32eb34} /* (22, 24, 14) {real, imag} */,
  {32'h3e2cbe70, 32'hbf60fdc6} /* (22, 24, 13) {real, imag} */,
  {32'h3e624310, 32'hbf9ff6cb} /* (22, 24, 12) {real, imag} */,
  {32'hbf87eec2, 32'hbdc777e8} /* (22, 24, 11) {real, imag} */,
  {32'hbe9538bc, 32'hbfa3eb7b} /* (22, 24, 10) {real, imag} */,
  {32'hbfad9db6, 32'hbefa0954} /* (22, 24, 9) {real, imag} */,
  {32'hc01131d2, 32'hbebbbc00} /* (22, 24, 8) {real, imag} */,
  {32'hbf514009, 32'h3e5090f8} /* (22, 24, 7) {real, imag} */,
  {32'hbf81b2d6, 32'hbf6a8b62} /* (22, 24, 6) {real, imag} */,
  {32'hbfc7dc5b, 32'hbfeafe0f} /* (22, 24, 5) {real, imag} */,
  {32'hbfacaa44, 32'hbe598bbc} /* (22, 24, 4) {real, imag} */,
  {32'hbf97b080, 32'h3f1e5aea} /* (22, 24, 3) {real, imag} */,
  {32'hbe6652f0, 32'h3b8a0a00} /* (22, 24, 2) {real, imag} */,
  {32'hbf58dcc8, 32'hbf46daf3} /* (22, 24, 1) {real, imag} */,
  {32'h3e50c4b0, 32'hbf3768ac} /* (22, 24, 0) {real, imag} */,
  {32'hbfa9fef4, 32'hbf4d3024} /* (22, 23, 31) {real, imag} */,
  {32'hc044c9e2, 32'hc003088d} /* (22, 23, 30) {real, imag} */,
  {32'hc00d9832, 32'hbfaa8a18} /* (22, 23, 29) {real, imag} */,
  {32'hc03e48a6, 32'hbf5dfcc0} /* (22, 23, 28) {real, imag} */,
  {32'hc0091c52, 32'hbf900890} /* (22, 23, 27) {real, imag} */,
  {32'hbe3d13c8, 32'hbf5f09d2} /* (22, 23, 26) {real, imag} */,
  {32'hbea44fc4, 32'hbf014a4c} /* (22, 23, 25) {real, imag} */,
  {32'hbfa9dd9e, 32'hbf02b750} /* (22, 23, 24) {real, imag} */,
  {32'hc058cef1, 32'hbd97f7a0} /* (22, 23, 23) {real, imag} */,
  {32'hc0197bc4, 32'h400f73ef} /* (22, 23, 22) {real, imag} */,
  {32'hbf5c72e6, 32'hbee53b2a} /* (22, 23, 21) {real, imag} */,
  {32'hbdcede10, 32'hbf812ef9} /* (22, 23, 20) {real, imag} */,
  {32'h3f6a1d92, 32'h3e129888} /* (22, 23, 19) {real, imag} */,
  {32'h3df8c850, 32'hbf0954ba} /* (22, 23, 18) {real, imag} */,
  {32'hbee920b4, 32'hbf1a7524} /* (22, 23, 17) {real, imag} */,
  {32'h3ef4cafe, 32'h3f2d65b0} /* (22, 23, 16) {real, imag} */,
  {32'h3ff1e3f2, 32'h3fc33d4c} /* (22, 23, 15) {real, imag} */,
  {32'h400f218e, 32'h3f980fc3} /* (22, 23, 14) {real, imag} */,
  {32'h3ef9a410, 32'hbefda02c} /* (22, 23, 13) {real, imag} */,
  {32'h3e4a8be8, 32'hbe9388b4} /* (22, 23, 12) {real, imag} */,
  {32'hbf0f2367, 32'h3f6f9e20} /* (22, 23, 11) {real, imag} */,
  {32'hbfc2b7fe, 32'hbdce5e28} /* (22, 23, 10) {real, imag} */,
  {32'hc00916b0, 32'hbf8101c1} /* (22, 23, 9) {real, imag} */,
  {32'hbf2ba7ef, 32'hbf6c9157} /* (22, 23, 8) {real, imag} */,
  {32'hbe497f44, 32'h3e9b484c} /* (22, 23, 7) {real, imag} */,
  {32'hbf4dd74e, 32'h3f79c25e} /* (22, 23, 6) {real, imag} */,
  {32'hc0086b9f, 32'h3f1aaf9b} /* (22, 23, 5) {real, imag} */,
  {32'hbfce58e8, 32'h3db856d0} /* (22, 23, 4) {real, imag} */,
  {32'hbfa6b4b4, 32'h3f707142} /* (22, 23, 3) {real, imag} */,
  {32'hbd83c350, 32'h3ff98b00} /* (22, 23, 2) {real, imag} */,
  {32'h3e8dc888, 32'h3f86ce76} /* (22, 23, 1) {real, imag} */,
  {32'hbf284cca, 32'h3ef92e82} /* (22, 23, 0) {real, imag} */,
  {32'h3d4c8b40, 32'hbeebd32a} /* (22, 22, 31) {real, imag} */,
  {32'hc01deb2e, 32'hbf55c2aa} /* (22, 22, 30) {real, imag} */,
  {32'hc01f5fe0, 32'hbed91d80} /* (22, 22, 29) {real, imag} */,
  {32'hbfa99528, 32'hbf0bb888} /* (22, 22, 28) {real, imag} */,
  {32'hbf98e766, 32'h3bcd0800} /* (22, 22, 27) {real, imag} */,
  {32'hbedf92d0, 32'hbec41320} /* (22, 22, 26) {real, imag} */,
  {32'hbebc9524, 32'hbfc484e0} /* (22, 22, 25) {real, imag} */,
  {32'hbf37255a, 32'hbfa76eb2} /* (22, 22, 24) {real, imag} */,
  {32'hbfb56d7e, 32'hbf764b54} /* (22, 22, 23) {real, imag} */,
  {32'hbf70774c, 32'h3ed3af1a} /* (22, 22, 22) {real, imag} */,
  {32'hbe7dbf7c, 32'h3dad48e8} /* (22, 22, 21) {real, imag} */,
  {32'hbfa07ec0, 32'hbe948acc} /* (22, 22, 20) {real, imag} */,
  {32'hbfab0bc4, 32'h3e4c48c0} /* (22, 22, 19) {real, imag} */,
  {32'hbf14e724, 32'h3f9d6056} /* (22, 22, 18) {real, imag} */,
  {32'h3f005174, 32'h3f998bce} /* (22, 22, 17) {real, imag} */,
  {32'h3fbb75e4, 32'h3f87ef86} /* (22, 22, 16) {real, imag} */,
  {32'h3f431675, 32'h3f7d4867} /* (22, 22, 15) {real, imag} */,
  {32'h3ed310c6, 32'h3f568786} /* (22, 22, 14) {real, imag} */,
  {32'h3f507b84, 32'hbf2d7608} /* (22, 22, 13) {real, imag} */,
  {32'h3ea76366, 32'h3f73cc5d} /* (22, 22, 12) {real, imag} */,
  {32'h3ebd5f98, 32'h3fddcdd8} /* (22, 22, 11) {real, imag} */,
  {32'hbfd360d8, 32'h3e4b33c4} /* (22, 22, 10) {real, imag} */,
  {32'hc02944fd, 32'hbfa74439} /* (22, 22, 9) {real, imag} */,
  {32'hbe69a034, 32'h3eaa85fc} /* (22, 22, 8) {real, imag} */,
  {32'hbc9cde60, 32'h400b5ecc} /* (22, 22, 7) {real, imag} */,
  {32'hbe2b7ce0, 32'h3fc4ccf0} /* (22, 22, 6) {real, imag} */,
  {32'hbf35dfa8, 32'h3fa425e8} /* (22, 22, 5) {real, imag} */,
  {32'hbf7d0e44, 32'hbf5d51fa} /* (22, 22, 4) {real, imag} */,
  {32'hbe915f04, 32'h3e33e8c0} /* (22, 22, 3) {real, imag} */,
  {32'h3e7be680, 32'h3fc2f93a} /* (22, 22, 2) {real, imag} */,
  {32'hbf2092db, 32'h3ef10308} /* (22, 22, 1) {real, imag} */,
  {32'hbe3d6798, 32'h3f06718d} /* (22, 22, 0) {real, imag} */,
  {32'h3ea0735a, 32'h3f5b24b2} /* (22, 21, 31) {real, imag} */,
  {32'hbd2927a0, 32'h3f5d12e0} /* (22, 21, 30) {real, imag} */,
  {32'hbf0d99eb, 32'hbfb9ba0d} /* (22, 21, 29) {real, imag} */,
  {32'hbfbed6dc, 32'hc0136fe1} /* (22, 21, 28) {real, imag} */,
  {32'hbf669370, 32'h3f11529f} /* (22, 21, 27) {real, imag} */,
  {32'hbe8233f4, 32'h3d97aac0} /* (22, 21, 26) {real, imag} */,
  {32'hbe355117, 32'hbf5f8a6d} /* (22, 21, 25) {real, imag} */,
  {32'h3f036f7a, 32'hbfd03c66} /* (22, 21, 24) {real, imag} */,
  {32'hbdac18b4, 32'hbf610e98} /* (22, 21, 23) {real, imag} */,
  {32'h3eff2ffa, 32'hbf3229fe} /* (22, 21, 22) {real, imag} */,
  {32'h3f21d382, 32'h3dba4da0} /* (22, 21, 21) {real, imag} */,
  {32'hbfc1dced, 32'hbee37baf} /* (22, 21, 20) {real, imag} */,
  {32'hbfebc42b, 32'h3cff5860} /* (22, 21, 19) {real, imag} */,
  {32'h3dc78d88, 32'h3fe29f2b} /* (22, 21, 18) {real, imag} */,
  {32'h3fa55cbe, 32'h3f72576e} /* (22, 21, 17) {real, imag} */,
  {32'h3fc020f4, 32'h3cf0f9d8} /* (22, 21, 16) {real, imag} */,
  {32'h3e670c14, 32'h3f25d8f8} /* (22, 21, 15) {real, imag} */,
  {32'h3f83cf5e, 32'h3fd8a398} /* (22, 21, 14) {real, imag} */,
  {32'h3fa8d5bc, 32'h3dde59b8} /* (22, 21, 13) {real, imag} */,
  {32'h3ecf7090, 32'hbf10ef77} /* (22, 21, 12) {real, imag} */,
  {32'hbf3835a2, 32'h3f59c77d} /* (22, 21, 11) {real, imag} */,
  {32'hc007438e, 32'h3ebff4b2} /* (22, 21, 10) {real, imag} */,
  {32'hc04303b1, 32'h400ca805} /* (22, 21, 9) {real, imag} */,
  {32'hbf148758, 32'h3fd747cb} /* (22, 21, 8) {real, imag} */,
  {32'h3d483548, 32'h3f87d91d} /* (22, 21, 7) {real, imag} */,
  {32'hbf931908, 32'hbec32be4} /* (22, 21, 6) {real, imag} */,
  {32'hbf36e444, 32'h3ecc6198} /* (22, 21, 5) {real, imag} */,
  {32'hbeb4b103, 32'hbf60c6a6} /* (22, 21, 4) {real, imag} */,
  {32'hbfda9306, 32'h3e6ed3e6} /* (22, 21, 3) {real, imag} */,
  {32'hbe87a9b4, 32'h3f4bfad5} /* (22, 21, 2) {real, imag} */,
  {32'hbd3e3c00, 32'h3f15101d} /* (22, 21, 1) {real, imag} */,
  {32'h3f63de9a, 32'h3e4706f0} /* (22, 21, 0) {real, imag} */,
  {32'h3f26760c, 32'h400825fb} /* (22, 20, 31) {real, imag} */,
  {32'h3fbcf81f, 32'h406239f0} /* (22, 20, 30) {real, imag} */,
  {32'h3f8f5c59, 32'hbda13880} /* (22, 20, 29) {real, imag} */,
  {32'h3f270318, 32'hbfc569e0} /* (22, 20, 28) {real, imag} */,
  {32'h3f4393ea, 32'hbecb6ee8} /* (22, 20, 27) {real, imag} */,
  {32'h3fa100ea, 32'h3f021576} /* (22, 20, 26) {real, imag} */,
  {32'h3fbacd9f, 32'h3f93de2a} /* (22, 20, 25) {real, imag} */,
  {32'h401764d8, 32'hbbe3e900} /* (22, 20, 24) {real, imag} */,
  {32'h3f261099, 32'h3f471d95} /* (22, 20, 23) {real, imag} */,
  {32'hbe8fe1c8, 32'h3e2e2bf8} /* (22, 20, 22) {real, imag} */,
  {32'h3ee63206, 32'h3f55777c} /* (22, 20, 21) {real, imag} */,
  {32'hbf066cd8, 32'hbf44186a} /* (22, 20, 20) {real, imag} */,
  {32'hbf461fd0, 32'hbf650566} /* (22, 20, 19) {real, imag} */,
  {32'h3e5eb7bb, 32'h3f86b28a} /* (22, 20, 18) {real, imag} */,
  {32'h3f8524a3, 32'h3ee61330} /* (22, 20, 17) {real, imag} */,
  {32'h3f193698, 32'hbeee5d60} /* (22, 20, 16) {real, imag} */,
  {32'h3e6f0780, 32'hbecc7dbc} /* (22, 20, 15) {real, imag} */,
  {32'h40057b86, 32'h3f8351f8} /* (22, 20, 14) {real, imag} */,
  {32'h3db6aa80, 32'hbcf4ea60} /* (22, 20, 13) {real, imag} */,
  {32'hbfe4c767, 32'hbf824616} /* (22, 20, 12) {real, imag} */,
  {32'hbf8dc085, 32'hbe14eda8} /* (22, 20, 11) {real, imag} */,
  {32'hbfb2d6db, 32'hbe36fbc8} /* (22, 20, 10) {real, imag} */,
  {32'hbfa5b6c4, 32'h40051850} /* (22, 20, 9) {real, imag} */,
  {32'h3f25b9b0, 32'h3f1f71b6} /* (22, 20, 8) {real, imag} */,
  {32'h3f85cc03, 32'hbf774947} /* (22, 20, 7) {real, imag} */,
  {32'hbe11c344, 32'hbf1a4a1c} /* (22, 20, 6) {real, imag} */,
  {32'hbe4c47cc, 32'h3dd76db8} /* (22, 20, 5) {real, imag} */,
  {32'h3e63e2a0, 32'hbf882a12} /* (22, 20, 4) {real, imag} */,
  {32'hbf5bf39e, 32'hbf95be26} /* (22, 20, 3) {real, imag} */,
  {32'hbf3cc69c, 32'hbf17d470} /* (22, 20, 2) {real, imag} */,
  {32'hbea9d054, 32'h3e5e1108} /* (22, 20, 1) {real, imag} */,
  {32'h3f3bf9f2, 32'hbe2a23cd} /* (22, 20, 0) {real, imag} */,
  {32'h3e54bcb0, 32'h3fa3884e} /* (22, 19, 31) {real, imag} */,
  {32'h3e602354, 32'h40253987} /* (22, 19, 30) {real, imag} */,
  {32'hbf2a7abe, 32'h3ec0d8e8} /* (22, 19, 29) {real, imag} */,
  {32'h3e8d49be, 32'hbfb9ebf2} /* (22, 19, 28) {real, imag} */,
  {32'h3fc29046, 32'hbf9ffec2} /* (22, 19, 27) {real, imag} */,
  {32'h400c2744, 32'h3d43cdd0} /* (22, 19, 26) {real, imag} */,
  {32'h3fffd988, 32'h3fa508cf} /* (22, 19, 25) {real, imag} */,
  {32'h3fabc5d6, 32'h3f498c76} /* (22, 19, 24) {real, imag} */,
  {32'hbef98cc4, 32'h401dfbe8} /* (22, 19, 23) {real, imag} */,
  {32'hbf7fe88f, 32'h3f685756} /* (22, 19, 22) {real, imag} */,
  {32'hbe9d090e, 32'h3fce439e} /* (22, 19, 21) {real, imag} */,
  {32'hbf82a4e4, 32'h3eddac54} /* (22, 19, 20) {real, imag} */,
  {32'hbf361148, 32'hbfb03dd4} /* (22, 19, 19) {real, imag} */,
  {32'h3f1f709e, 32'hbed4a394} /* (22, 19, 18) {real, imag} */,
  {32'h3fd7e628, 32'h3ef1ed50} /* (22, 19, 17) {real, imag} */,
  {32'h3f9dbf05, 32'hbf05b5a9} /* (22, 19, 16) {real, imag} */,
  {32'hbe4cde70, 32'hbf73e6c8} /* (22, 19, 15) {real, imag} */,
  {32'h3f01247c, 32'hbf520690} /* (22, 19, 14) {real, imag} */,
  {32'hbfcbf0b6, 32'hbeb823f8} /* (22, 19, 13) {real, imag} */,
  {32'hbfd58ca0, 32'h3f9f6a7f} /* (22, 19, 12) {real, imag} */,
  {32'hbf9d2410, 32'h3f19b4b4} /* (22, 19, 11) {real, imag} */,
  {32'hbf0866cc, 32'hbe41ddd8} /* (22, 19, 10) {real, imag} */,
  {32'h3fa14502, 32'h3ee31d48} /* (22, 19, 9) {real, imag} */,
  {32'h3f742874, 32'hbf8b46b8} /* (22, 19, 8) {real, imag} */,
  {32'h3fa768dd, 32'hc013b8ce} /* (22, 19, 7) {real, imag} */,
  {32'h3f0d93f8, 32'hbec91f94} /* (22, 19, 6) {real, imag} */,
  {32'h3e53099c, 32'h3fcf70d8} /* (22, 19, 5) {real, imag} */,
  {32'h40035504, 32'h3f873217} /* (22, 19, 4) {real, imag} */,
  {32'h3fd7f02a, 32'h3e41ab50} /* (22, 19, 3) {real, imag} */,
  {32'hbf0c7f7a, 32'hbec85fbc} /* (22, 19, 2) {real, imag} */,
  {32'hbe3909d8, 32'h3fec228a} /* (22, 19, 1) {real, imag} */,
  {32'h3f798217, 32'h40160f61} /* (22, 19, 0) {real, imag} */,
  {32'h3f80b34a, 32'h3e8e0e64} /* (22, 18, 31) {real, imag} */,
  {32'h3f0b1b3c, 32'h3f608920} /* (22, 18, 30) {real, imag} */,
  {32'hbf89de7b, 32'h40017357} /* (22, 18, 29) {real, imag} */,
  {32'hbf99efd5, 32'h3eb79c9e} /* (22, 18, 28) {real, imag} */,
  {32'hbe69e828, 32'hbf667f2c} /* (22, 18, 27) {real, imag} */,
  {32'h3fbc3001, 32'hbf56d31a} /* (22, 18, 26) {real, imag} */,
  {32'h3f99c23c, 32'hbf100c82} /* (22, 18, 25) {real, imag} */,
  {32'h3fad1020, 32'h3e601350} /* (22, 18, 24) {real, imag} */,
  {32'h3e99615c, 32'h40149db0} /* (22, 18, 23) {real, imag} */,
  {32'hbf0e95d6, 32'h3fdbde1b} /* (22, 18, 22) {real, imag} */,
  {32'hbf5e73e7, 32'h4007e474} /* (22, 18, 21) {real, imag} */,
  {32'hbfd6114f, 32'hbf8bb4c0} /* (22, 18, 20) {real, imag} */,
  {32'hbf3f2f83, 32'hc02055f4} /* (22, 18, 19) {real, imag} */,
  {32'hbf4cd54e, 32'hbf8c27e8} /* (22, 18, 18) {real, imag} */,
  {32'h3eb7d36c, 32'h3f7baf68} /* (22, 18, 17) {real, imag} */,
  {32'h3f59d128, 32'h3ebdeb40} /* (22, 18, 16) {real, imag} */,
  {32'hbe32c8c0, 32'h3e824dc0} /* (22, 18, 15) {real, imag} */,
  {32'hbee0dea0, 32'hbf1f3416} /* (22, 18, 14) {real, imag} */,
  {32'hc02a4f98, 32'hbf8f3a8d} /* (22, 18, 13) {real, imag} */,
  {32'hc01a01cb, 32'h3f958daf} /* (22, 18, 12) {real, imag} */,
  {32'hbf9c70f9, 32'h3fec9b70} /* (22, 18, 11) {real, imag} */,
  {32'h3e41da04, 32'h4018e500} /* (22, 18, 10) {real, imag} */,
  {32'h3dea0b00, 32'h3fc84dfe} /* (22, 18, 9) {real, imag} */,
  {32'h3e7f85b0, 32'hbf389a02} /* (22, 18, 8) {real, imag} */,
  {32'h400b986a, 32'hbff3669a} /* (22, 18, 7) {real, imag} */,
  {32'h3ffda25a, 32'hbeff5350} /* (22, 18, 6) {real, imag} */,
  {32'h3f5213ec, 32'h3f962f8e} /* (22, 18, 5) {real, imag} */,
  {32'h3fa71ed2, 32'h3f6b1f18} /* (22, 18, 4) {real, imag} */,
  {32'h3f1a97b8, 32'h3f5a881c} /* (22, 18, 3) {real, imag} */,
  {32'hbe5bc2b0, 32'h3f917d22} /* (22, 18, 2) {real, imag} */,
  {32'hbc782d00, 32'h3fd8f0ce} /* (22, 18, 1) {real, imag} */,
  {32'h3e9bbd38, 32'h400b6d6e} /* (22, 18, 0) {real, imag} */,
  {32'h3f9496ca, 32'h3f3ab17c} /* (22, 17, 31) {real, imag} */,
  {32'h3f6f78ba, 32'h3f9a1c92} /* (22, 17, 30) {real, imag} */,
  {32'h3eb2af2a, 32'h3ff15b0c} /* (22, 17, 29) {real, imag} */,
  {32'h3e5c2bd8, 32'h3ff15baf} /* (22, 17, 28) {real, imag} */,
  {32'hbf0f1472, 32'h3e6a8fd0} /* (22, 17, 27) {real, imag} */,
  {32'hbd0aa270, 32'h3f940b99} /* (22, 17, 26) {real, imag} */,
  {32'h3f487e16, 32'hbc2bc080} /* (22, 17, 25) {real, imag} */,
  {32'h3f36cecc, 32'hbf57f5a0} /* (22, 17, 24) {real, imag} */,
  {32'hbda4e440, 32'h3e847d90} /* (22, 17, 23) {real, imag} */,
  {32'hbf06eb61, 32'h3dd583f8} /* (22, 17, 22) {real, imag} */,
  {32'hbfaa10d4, 32'hbf39351e} /* (22, 17, 21) {real, imag} */,
  {32'hc0279436, 32'hc00665e2} /* (22, 17, 20) {real, imag} */,
  {32'hbf8f0983, 32'hbf5f3ba0} /* (22, 17, 19) {real, imag} */,
  {32'hbfbfe706, 32'h3edb4768} /* (22, 17, 18) {real, imag} */,
  {32'h3e3725e8, 32'h3f6173e2} /* (22, 17, 17) {real, imag} */,
  {32'hbea01768, 32'hbf7570b0} /* (22, 17, 16) {real, imag} */,
  {32'hbc3a9900, 32'hbf243744} /* (22, 17, 15) {real, imag} */,
  {32'hbe808634, 32'h3f559824} /* (22, 17, 14) {real, imag} */,
  {32'hbf9b05f8, 32'h3e7e7a6c} /* (22, 17, 13) {real, imag} */,
  {32'hbf129cf0, 32'h3efed450} /* (22, 17, 12) {real, imag} */,
  {32'hbf755733, 32'h3f8aff3c} /* (22, 17, 11) {real, imag} */,
  {32'h3f35054e, 32'h400068ef} /* (22, 17, 10) {real, imag} */,
  {32'h3f382e90, 32'h400f116d} /* (22, 17, 9) {real, imag} */,
  {32'h3f76c4a4, 32'h3f09e9b4} /* (22, 17, 8) {real, imag} */,
  {32'h3fe155cf, 32'hbf7a9d08} /* (22, 17, 7) {real, imag} */,
  {32'h3fcdcdec, 32'hbf719182} /* (22, 17, 6) {real, imag} */,
  {32'h3f92518e, 32'h3f8eaa20} /* (22, 17, 5) {real, imag} */,
  {32'h4015d934, 32'h3f418aac} /* (22, 17, 4) {real, imag} */,
  {32'h3f50a084, 32'h3d6feb00} /* (22, 17, 3) {real, imag} */,
  {32'hbf2acf60, 32'hbee48a74} /* (22, 17, 2) {real, imag} */,
  {32'hbfad54d5, 32'h3f8193fb} /* (22, 17, 1) {real, imag} */,
  {32'hbea97e24, 32'h3f4dde4a} /* (22, 17, 0) {real, imag} */,
  {32'h3f6b83f0, 32'hbc8a76a0} /* (22, 16, 31) {real, imag} */,
  {32'h3fb2e144, 32'h3f1f5108} /* (22, 16, 30) {real, imag} */,
  {32'h3fbe11bd, 32'h3f9a718a} /* (22, 16, 29) {real, imag} */,
  {32'h3f836dd3, 32'h3ee1c500} /* (22, 16, 28) {real, imag} */,
  {32'hbbd8f500, 32'h3f0e6040} /* (22, 16, 27) {real, imag} */,
  {32'hbdf69d30, 32'h3fbd2201} /* (22, 16, 26) {real, imag} */,
  {32'h3f8008a6, 32'h3f083b64} /* (22, 16, 25) {real, imag} */,
  {32'h3f9a86d4, 32'hbfadff0b} /* (22, 16, 24) {real, imag} */,
  {32'h3ea47480, 32'hbf472d40} /* (22, 16, 23) {real, imag} */,
  {32'hbf8f3444, 32'hbdfef040} /* (22, 16, 22) {real, imag} */,
  {32'hc00c0669, 32'h3f0d20f1} /* (22, 16, 21) {real, imag} */,
  {32'hbfdd3463, 32'h3ebdcf20} /* (22, 16, 20) {real, imag} */,
  {32'hbfa30386, 32'h3f46a8ba} /* (22, 16, 19) {real, imag} */,
  {32'hc007312c, 32'h3f1e8000} /* (22, 16, 18) {real, imag} */,
  {32'hc0011bd4, 32'hbd38aa40} /* (22, 16, 17) {real, imag} */,
  {32'hbf1a7c44, 32'hbf425d06} /* (22, 16, 16) {real, imag} */,
  {32'h3eabb02c, 32'hbca758c0} /* (22, 16, 15) {real, imag} */,
  {32'hbe7e14a8, 32'h3ed98620} /* (22, 16, 14) {real, imag} */,
  {32'hbfaea407, 32'hbf98614f} /* (22, 16, 13) {real, imag} */,
  {32'hbf2b08bc, 32'hbf512456} /* (22, 16, 12) {real, imag} */,
  {32'hbfcd14a2, 32'h3ed4c580} /* (22, 16, 11) {real, imag} */,
  {32'h3f633c33, 32'h3ee860a4} /* (22, 16, 10) {real, imag} */,
  {32'h3ff65334, 32'h4003c44f} /* (22, 16, 9) {real, imag} */,
  {32'h3f82a738, 32'h3fb70d5f} /* (22, 16, 8) {real, imag} */,
  {32'h3fc64182, 32'h3e00bf14} /* (22, 16, 7) {real, imag} */,
  {32'h3fcd83ef, 32'hbf16398e} /* (22, 16, 6) {real, imag} */,
  {32'h3f711628, 32'h3f45af2e} /* (22, 16, 5) {real, imag} */,
  {32'h3ff74f30, 32'h3f0855da} /* (22, 16, 4) {real, imag} */,
  {32'h3fcf4af2, 32'hbf8213c1} /* (22, 16, 3) {real, imag} */,
  {32'hbe4d2d20, 32'hbfb8ccaf} /* (22, 16, 2) {real, imag} */,
  {32'hc00d6f9f, 32'h3f254b07} /* (22, 16, 1) {real, imag} */,
  {32'hbf48f42c, 32'h3f856f32} /* (22, 16, 0) {real, imag} */,
  {32'h3f06af20, 32'hbc685640} /* (22, 15, 31) {real, imag} */,
  {32'h3fa9515a, 32'h3e8f81b8} /* (22, 15, 30) {real, imag} */,
  {32'h3f9c6d37, 32'h3da64008} /* (22, 15, 29) {real, imag} */,
  {32'h3f94b8e4, 32'hbf35d84a} /* (22, 15, 28) {real, imag} */,
  {32'h3f1239f2, 32'h3f0a7578} /* (22, 15, 27) {real, imag} */,
  {32'h3f3d76c6, 32'h3f733fde} /* (22, 15, 26) {real, imag} */,
  {32'h3e5eff78, 32'h3f82d898} /* (22, 15, 25) {real, imag} */,
  {32'h3fcbcce2, 32'h3ea9d596} /* (22, 15, 24) {real, imag} */,
  {32'h400547c2, 32'hbf35bb00} /* (22, 15, 23) {real, imag} */,
  {32'h3f82afd1, 32'hbf7d34e8} /* (22, 15, 22) {real, imag} */,
  {32'hbf88b92c, 32'h3ecfed6c} /* (22, 15, 21) {real, imag} */,
  {32'hbf96f709, 32'hbf4b8bda} /* (22, 15, 20) {real, imag} */,
  {32'hbfff760d, 32'hbf529a29} /* (22, 15, 19) {real, imag} */,
  {32'hc00bff80, 32'hbf800160} /* (22, 15, 18) {real, imag} */,
  {32'hbfdb1342, 32'hbee4d390} /* (22, 15, 17) {real, imag} */,
  {32'hbed46f6e, 32'h3edee960} /* (22, 15, 16) {real, imag} */,
  {32'hbf126d14, 32'h3f6b955e} /* (22, 15, 15) {real, imag} */,
  {32'hbd17bdb0, 32'h3f38d06e} /* (22, 15, 14) {real, imag} */,
  {32'h3f0f82b1, 32'hc019bfeb} /* (22, 15, 13) {real, imag} */,
  {32'h3f441f14, 32'hc009c916} /* (22, 15, 12) {real, imag} */,
  {32'hbf5e821a, 32'h3df2cd90} /* (22, 15, 11) {real, imag} */,
  {32'h3eb1ff80, 32'h3f4221ee} /* (22, 15, 10) {real, imag} */,
  {32'h3f82b307, 32'h3ef6cd80} /* (22, 15, 9) {real, imag} */,
  {32'h3f1b759a, 32'hbec120a6} /* (22, 15, 8) {real, imag} */,
  {32'h3f958a5a, 32'hbeedfc70} /* (22, 15, 7) {real, imag} */,
  {32'h4007836f, 32'h3f59c1da} /* (22, 15, 6) {real, imag} */,
  {32'h400d182b, 32'h3cb659c0} /* (22, 15, 5) {real, imag} */,
  {32'h3f983b82, 32'hbe4ba0e0} /* (22, 15, 4) {real, imag} */,
  {32'h3f54dd24, 32'h3e16c718} /* (22, 15, 3) {real, imag} */,
  {32'hbee4779c, 32'h3e0e80e0} /* (22, 15, 2) {real, imag} */,
  {32'hc01ddd3a, 32'h3e0ebad8} /* (22, 15, 1) {real, imag} */,
  {32'hbf83ae6c, 32'h3f18fc31} /* (22, 15, 0) {real, imag} */,
  {32'h3e8e3578, 32'h3df71ec0} /* (22, 14, 31) {real, imag} */,
  {32'h3fbeacb0, 32'hbf32d496} /* (22, 14, 30) {real, imag} */,
  {32'h3ee16868, 32'h3e65d790} /* (22, 14, 29) {real, imag} */,
  {32'h3f0ca06c, 32'h3f59615a} /* (22, 14, 28) {real, imag} */,
  {32'h3efba1dc, 32'h3fa0997b} /* (22, 14, 27) {real, imag} */,
  {32'h3f0815a6, 32'h3fa8f012} /* (22, 14, 26) {real, imag} */,
  {32'h3e959db8, 32'h3f959042} /* (22, 14, 25) {real, imag} */,
  {32'h3f9b43e7, 32'h3fa9fa66} /* (22, 14, 24) {real, imag} */,
  {32'h3fe23835, 32'h3e671468} /* (22, 14, 23) {real, imag} */,
  {32'h4003679a, 32'hbecd6704} /* (22, 14, 22) {real, imag} */,
  {32'h3f79bc8e, 32'hbe907962} /* (22, 14, 21) {real, imag} */,
  {32'hbf92831e, 32'hbf8e61e6} /* (22, 14, 20) {real, imag} */,
  {32'hbf888980, 32'hbf5b98f4} /* (22, 14, 19) {real, imag} */,
  {32'hbf9bbfd4, 32'hbf7586c4} /* (22, 14, 18) {real, imag} */,
  {32'hbe3b7514, 32'hbf1c654a} /* (22, 14, 17) {real, imag} */,
  {32'hbe15dfca, 32'h3fe1176a} /* (22, 14, 16) {real, imag} */,
  {32'hbf1ccd13, 32'h3f3ea842} /* (22, 14, 15) {real, imag} */,
  {32'h3fc73504, 32'hbedddb8e} /* (22, 14, 14) {real, imag} */,
  {32'h3fa7c63a, 32'hbfca4a48} /* (22, 14, 13) {real, imag} */,
  {32'hbf1044e2, 32'hbfa8f454} /* (22, 14, 12) {real, imag} */,
  {32'hbf18707c, 32'h3f1e04e4} /* (22, 14, 11) {real, imag} */,
  {32'hbf53f0c1, 32'h3f486c8a} /* (22, 14, 10) {real, imag} */,
  {32'hbf0d6a2e, 32'h3da2f870} /* (22, 14, 9) {real, imag} */,
  {32'h3edd670c, 32'hbd3afda0} /* (22, 14, 8) {real, imag} */,
  {32'h3f8fd342, 32'h3f392ab1} /* (22, 14, 7) {real, imag} */,
  {32'h3f29404e, 32'h3f0da995} /* (22, 14, 6) {real, imag} */,
  {32'h3e187b49, 32'hbfa6b173} /* (22, 14, 5) {real, imag} */,
  {32'h3f4f3b52, 32'hbf9fd48a} /* (22, 14, 4) {real, imag} */,
  {32'h3f09a0f7, 32'hbf6ca7d4} /* (22, 14, 3) {real, imag} */,
  {32'hbfa29402, 32'hbde737b0} /* (22, 14, 2) {real, imag} */,
  {32'hbfb33548, 32'hbda272c0} /* (22, 14, 1) {real, imag} */,
  {32'hbf36e159, 32'hbd9d5700} /* (22, 14, 0) {real, imag} */,
  {32'h3f6c349c, 32'hbe86d49e} /* (22, 13, 31) {real, imag} */,
  {32'h40074597, 32'hbfb5e566} /* (22, 13, 30) {real, imag} */,
  {32'hbf20fe05, 32'h3d981970} /* (22, 13, 29) {real, imag} */,
  {32'hbfa07024, 32'hbf221da6} /* (22, 13, 28) {real, imag} */,
  {32'hbf4604aa, 32'h3e463b3c} /* (22, 13, 27) {real, imag} */,
  {32'hbc35eb40, 32'h3f603bb6} /* (22, 13, 26) {real, imag} */,
  {32'h3f5f4ca8, 32'h3d935888} /* (22, 13, 25) {real, imag} */,
  {32'h3e4640c0, 32'h3f2deb48} /* (22, 13, 24) {real, imag} */,
  {32'h3f2dcd1c, 32'h3e6be418} /* (22, 13, 23) {real, imag} */,
  {32'h3f3dcf74, 32'h3ef0e1bc} /* (22, 13, 22) {real, imag} */,
  {32'h3f859d7a, 32'h3f179d5f} /* (22, 13, 21) {real, imag} */,
  {32'hbf3ff868, 32'h3e53e548} /* (22, 13, 20) {real, imag} */,
  {32'h3f12615c, 32'h3d05b800} /* (22, 13, 19) {real, imag} */,
  {32'h3f98b8fd, 32'hbf32e567} /* (22, 13, 18) {real, imag} */,
  {32'hbf51e9c8, 32'hbf143fc0} /* (22, 13, 17) {real, imag} */,
  {32'hbf9aa566, 32'h3fc0365a} /* (22, 13, 16) {real, imag} */,
  {32'hbf2cf6bb, 32'h3f35d454} /* (22, 13, 15) {real, imag} */,
  {32'h3ef62e9e, 32'hbf8b92a6} /* (22, 13, 14) {real, imag} */,
  {32'h3dc11c20, 32'hc0133d70} /* (22, 13, 13) {real, imag} */,
  {32'hbf4c4a6c, 32'hbf9623d9} /* (22, 13, 12) {real, imag} */,
  {32'hbdfad0b0, 32'h3f83c599} /* (22, 13, 11) {real, imag} */,
  {32'hbf3da80c, 32'h3feb4ae5} /* (22, 13, 10) {real, imag} */,
  {32'hbf3f1644, 32'h40148e12} /* (22, 13, 9) {real, imag} */,
  {32'hbee805b8, 32'h3f87e5f0} /* (22, 13, 8) {real, imag} */,
  {32'h3f5323aa, 32'h3de685c0} /* (22, 13, 7) {real, imag} */,
  {32'h3f9c92c0, 32'hbfa2f889} /* (22, 13, 6) {real, imag} */,
  {32'hbe3c2a58, 32'hc018fc7a} /* (22, 13, 5) {real, imag} */,
  {32'h3e5887b0, 32'hbf29bbba} /* (22, 13, 4) {real, imag} */,
  {32'h3e2a4270, 32'hbe3711e0} /* (22, 13, 3) {real, imag} */,
  {32'hbf176078, 32'h3f90244e} /* (22, 13, 2) {real, imag} */,
  {32'hbed778e0, 32'h3e07fb28} /* (22, 13, 1) {real, imag} */,
  {32'hbebb5af0, 32'h3f46a265} /* (22, 13, 0) {real, imag} */,
  {32'h3e4ddc1c, 32'h3f7eb3ca} /* (22, 12, 31) {real, imag} */,
  {32'h3f404f6f, 32'h3fae5d4a} /* (22, 12, 30) {real, imag} */,
  {32'hbd487240, 32'h3ec7854a} /* (22, 12, 29) {real, imag} */,
  {32'hbe9d04a8, 32'hbf98dde2} /* (22, 12, 28) {real, imag} */,
  {32'hbe1d1ca8, 32'h3e84f286} /* (22, 12, 27) {real, imag} */,
  {32'h3f549a29, 32'h3ff47691} /* (22, 12, 26) {real, imag} */,
  {32'h3f223996, 32'hbeb15348} /* (22, 12, 25) {real, imag} */,
  {32'h3e86ba78, 32'h3ea69fa8} /* (22, 12, 24) {real, imag} */,
  {32'h3f1dd3db, 32'h3f9852d5} /* (22, 12, 23) {real, imag} */,
  {32'h3fe68ff1, 32'h3fc75faf} /* (22, 12, 22) {real, imag} */,
  {32'h3fb43c4d, 32'h3f3fc413} /* (22, 12, 21) {real, imag} */,
  {32'h3f29dbac, 32'hbdd7bd70} /* (22, 12, 20) {real, imag} */,
  {32'h3ff6c6c4, 32'h3ecaee68} /* (22, 12, 19) {real, imag} */,
  {32'h3f174f65, 32'h3f163272} /* (22, 12, 18) {real, imag} */,
  {32'hbf91c941, 32'hbf363d7a} /* (22, 12, 17) {real, imag} */,
  {32'hbf841f05, 32'hbf4b8b3c} /* (22, 12, 16) {real, imag} */,
  {32'hbeb098c4, 32'h3e98af2e} /* (22, 12, 15) {real, imag} */,
  {32'hbf12055e, 32'hbe89ea74} /* (22, 12, 14) {real, imag} */,
  {32'hbf67b895, 32'hbf9b20bc} /* (22, 12, 13) {real, imag} */,
  {32'hbc88b170, 32'hbf99bb70} /* (22, 12, 12) {real, imag} */,
  {32'h3f9b08c6, 32'h3f0ac547} /* (22, 12, 11) {real, imag} */,
  {32'h3e8480a3, 32'h3ff4a352} /* (22, 12, 10) {real, imag} */,
  {32'hbe166dbc, 32'h4047a3ea} /* (22, 12, 9) {real, imag} */,
  {32'hbf03cc96, 32'h3ff50b62} /* (22, 12, 8) {real, imag} */,
  {32'h3d907470, 32'hbf0b31d8} /* (22, 12, 7) {real, imag} */,
  {32'h3f368dfc, 32'hbf9890be} /* (22, 12, 6) {real, imag} */,
  {32'hbe7c4df8, 32'hbf1fc508} /* (22, 12, 5) {real, imag} */,
  {32'h3e964e32, 32'h3f75b995} /* (22, 12, 4) {real, imag} */,
  {32'h3e7812ac, 32'h3fd1d86f} /* (22, 12, 3) {real, imag} */,
  {32'hbf26b9f6, 32'h3fbabe14} /* (22, 12, 2) {real, imag} */,
  {32'hbfb0aeaa, 32'h3d869060} /* (22, 12, 1) {real, imag} */,
  {32'hbf852a93, 32'h3f4af29c} /* (22, 12, 0) {real, imag} */,
  {32'hbf22759e, 32'h3dd5cdc8} /* (22, 11, 31) {real, imag} */,
  {32'hbcd23f70, 32'h3fa119e2} /* (22, 11, 30) {real, imag} */,
  {32'h3fa12b94, 32'h3f095d90} /* (22, 11, 29) {real, imag} */,
  {32'h3f7e333a, 32'h3f0187ba} /* (22, 11, 28) {real, imag} */,
  {32'h3e9967a4, 32'h3ff7da49} /* (22, 11, 27) {real, imag} */,
  {32'hbebd60a9, 32'h3f8500a4} /* (22, 11, 26) {real, imag} */,
  {32'hbd6ff570, 32'hbf2974f2} /* (22, 11, 25) {real, imag} */,
  {32'h3fc401f8, 32'h3f9f3210} /* (22, 11, 24) {real, imag} */,
  {32'h3e3d8aae, 32'h403b76a9} /* (22, 11, 23) {real, imag} */,
  {32'h3e8ab784, 32'h3f105f1f} /* (22, 11, 22) {real, imag} */,
  {32'hbe842074, 32'h3ea05508} /* (22, 11, 21) {real, imag} */,
  {32'hbf740300, 32'h3ef77a92} /* (22, 11, 20) {real, imag} */,
  {32'hbe6418ae, 32'h3f013ec2} /* (22, 11, 19) {real, imag} */,
  {32'h3f2b1cf8, 32'h3ea6137c} /* (22, 11, 18) {real, imag} */,
  {32'hbe318fbc, 32'hbde5b240} /* (22, 11, 17) {real, imag} */,
  {32'hbf04fea4, 32'h3eada4d0} /* (22, 11, 16) {real, imag} */,
  {32'hbee02b0c, 32'h3e76db10} /* (22, 11, 15) {real, imag} */,
  {32'hbf985104, 32'hbe19fd74} /* (22, 11, 14) {real, imag} */,
  {32'hbf7772f4, 32'h3ce0e300} /* (22, 11, 13) {real, imag} */,
  {32'hbf8aba5a, 32'hbf0d7242} /* (22, 11, 12) {real, imag} */,
  {32'h3eac7e7a, 32'h3ef60f38} /* (22, 11, 11) {real, imag} */,
  {32'h3f026dfd, 32'h3fc7f308} /* (22, 11, 10) {real, imag} */,
  {32'h3f118ced, 32'h3fae4636} /* (22, 11, 9) {real, imag} */,
  {32'h3fc1e3f7, 32'h3e31e74c} /* (22, 11, 8) {real, imag} */,
  {32'hbf51b514, 32'hbf5d3960} /* (22, 11, 7) {real, imag} */,
  {32'hbfb9fbd9, 32'h3e34b870} /* (22, 11, 6) {real, imag} */,
  {32'hbda796e0, 32'h3f9e6858} /* (22, 11, 5) {real, imag} */,
  {32'h3ede18f6, 32'h3f430987} /* (22, 11, 4) {real, imag} */,
  {32'h3ebd44cc, 32'hbf0fed8f} /* (22, 11, 3) {real, imag} */,
  {32'hbfad0a3c, 32'h3e826da8} /* (22, 11, 2) {real, imag} */,
  {32'hc00465ca, 32'h3d4b1b60} /* (22, 11, 1) {real, imag} */,
  {32'hbf876466, 32'hbf134da2} /* (22, 11, 0) {real, imag} */,
  {32'hbef68852, 32'h3dd39a10} /* (22, 10, 31) {real, imag} */,
  {32'hbedfb1e0, 32'h3f11cfc0} /* (22, 10, 30) {real, imag} */,
  {32'h3f47733e, 32'h3f5d7e12} /* (22, 10, 29) {real, imag} */,
  {32'h3f7c0094, 32'h3eb41f28} /* (22, 10, 28) {real, imag} */,
  {32'h3e85c6b8, 32'h3dade4c0} /* (22, 10, 27) {real, imag} */,
  {32'hbf1a60ee, 32'h3f6bbb95} /* (22, 10, 26) {real, imag} */,
  {32'h3e752afc, 32'h3f86b5e2} /* (22, 10, 25) {real, imag} */,
  {32'h3eeeb17e, 32'h3fc922e4} /* (22, 10, 24) {real, imag} */,
  {32'hc02c8517, 32'h3f791b18} /* (22, 10, 23) {real, imag} */,
  {32'hc03524c3, 32'hbf981191} /* (22, 10, 22) {real, imag} */,
  {32'hc0164a3e, 32'h3decb554} /* (22, 10, 21) {real, imag} */,
  {32'hbfe3bb2f, 32'h3fcdb09d} /* (22, 10, 20) {real, imag} */,
  {32'h3e125720, 32'h3eebd780} /* (22, 10, 19) {real, imag} */,
  {32'h3ffb145e, 32'hbf5a16ba} /* (22, 10, 18) {real, imag} */,
  {32'h3fa3ea71, 32'hbfbc14c0} /* (22, 10, 17) {real, imag} */,
  {32'h3e9c18c4, 32'hbed6ab54} /* (22, 10, 16) {real, imag} */,
  {32'h3d4cc64e, 32'h3f015ef1} /* (22, 10, 15) {real, imag} */,
  {32'hbf8dba52, 32'hbea38d80} /* (22, 10, 14) {real, imag} */,
  {32'hbf3fa0c8, 32'h3e19a1f8} /* (22, 10, 13) {real, imag} */,
  {32'hbfb76067, 32'hbf0271bd} /* (22, 10, 12) {real, imag} */,
  {32'hbf1a3166, 32'hbf7ebb14} /* (22, 10, 11) {real, imag} */,
  {32'h3f017e31, 32'h3cb83100} /* (22, 10, 10) {real, imag} */,
  {32'hbeddfa8c, 32'hbf30e86c} /* (22, 10, 9) {real, imag} */,
  {32'hbf6acf62, 32'hbeff401e} /* (22, 10, 8) {real, imag} */,
  {32'hbf8152a2, 32'hbecb8024} /* (22, 10, 7) {real, imag} */,
  {32'hbeb607f4, 32'h3f203b62} /* (22, 10, 6) {real, imag} */,
  {32'h3e7a08d8, 32'hbd2c15d0} /* (22, 10, 5) {real, imag} */,
  {32'h3edc6f8e, 32'h3f978e60} /* (22, 10, 4) {real, imag} */,
  {32'h3e239414, 32'hbe960aea} /* (22, 10, 3) {real, imag} */,
  {32'hbebf7a80, 32'hbf4291a0} /* (22, 10, 2) {real, imag} */,
  {32'h3e993fb0, 32'h40007a14} /* (22, 10, 1) {real, imag} */,
  {32'h3f51b440, 32'h3f80d1d8} /* (22, 10, 0) {real, imag} */,
  {32'h3ec77b6c, 32'hbed4a1d0} /* (22, 9, 31) {real, imag} */,
  {32'hbcb7dc60, 32'h3e103e30} /* (22, 9, 30) {real, imag} */,
  {32'hbde5d0c0, 32'h3f47e2de} /* (22, 9, 29) {real, imag} */,
  {32'h3ceca1a0, 32'h3e94ee5c} /* (22, 9, 28) {real, imag} */,
  {32'h3e8dd18a, 32'hbf153f37} /* (22, 9, 27) {real, imag} */,
  {32'hbb796e00, 32'h3e82ed9e} /* (22, 9, 26) {real, imag} */,
  {32'h3f4adaf7, 32'h3f7a6fcb} /* (22, 9, 25) {real, imag} */,
  {32'h3fa26768, 32'h3e8c86c0} /* (22, 9, 24) {real, imag} */,
  {32'hbfd0759a, 32'hbfb29cea} /* (22, 9, 23) {real, imag} */,
  {32'hc00e5f12, 32'hbff0af69} /* (22, 9, 22) {real, imag} */,
  {32'hbfbbe01c, 32'hbf06a0ba} /* (22, 9, 21) {real, imag} */,
  {32'hbfa993f3, 32'h3fca6047} /* (22, 9, 20) {real, imag} */,
  {32'h3f1eb253, 32'h3e4af998} /* (22, 9, 19) {real, imag} */,
  {32'h3fdb2d41, 32'hbf983dd2} /* (22, 9, 18) {real, imag} */,
  {32'h3f89ee3c, 32'hbf82e0e7} /* (22, 9, 17) {real, imag} */,
  {32'hbf10b2cc, 32'hbfcad4db} /* (22, 9, 16) {real, imag} */,
  {32'h3f2a09fa, 32'h3d11ba80} /* (22, 9, 15) {real, imag} */,
  {32'h3f1d6832, 32'h3e4d0a30} /* (22, 9, 14) {real, imag} */,
  {32'h3f462d94, 32'hbe3045f4} /* (22, 9, 13) {real, imag} */,
  {32'h3ed75f9e, 32'hbedfcb88} /* (22, 9, 12) {real, imag} */,
  {32'hbf90f469, 32'hbf959ea6} /* (22, 9, 11) {real, imag} */,
  {32'hbfb68760, 32'hbf5283ae} /* (22, 9, 10) {real, imag} */,
  {32'hbfd7c1c6, 32'hbf7f12a5} /* (22, 9, 9) {real, imag} */,
  {32'hbf0728a0, 32'hbeb1d0bc} /* (22, 9, 8) {real, imag} */,
  {32'h3edf09a4, 32'h3e844178} /* (22, 9, 7) {real, imag} */,
  {32'h3e5a5768, 32'h3f3a8f44} /* (22, 9, 6) {real, imag} */,
  {32'h3e826dd4, 32'h3e61b918} /* (22, 9, 5) {real, imag} */,
  {32'h3f709b5f, 32'h3fdc527d} /* (22, 9, 4) {real, imag} */,
  {32'h3f9f5412, 32'h3ff59971} /* (22, 9, 3) {real, imag} */,
  {32'h3f9c1527, 32'h3f8281a6} /* (22, 9, 2) {real, imag} */,
  {32'hbf06e59d, 32'h403d03ef} /* (22, 9, 1) {real, imag} */,
  {32'hbf2b3467, 32'h3fe2d34a} /* (22, 9, 0) {real, imag} */,
  {32'h3f26b710, 32'hbea13794} /* (22, 8, 31) {real, imag} */,
  {32'h3fa99ecf, 32'h3ece0618} /* (22, 8, 30) {real, imag} */,
  {32'hbe5b0d80, 32'h3eb49e10} /* (22, 8, 29) {real, imag} */,
  {32'h3d3dc140, 32'h3e8ace74} /* (22, 8, 28) {real, imag} */,
  {32'hbed32064, 32'hbf41955c} /* (22, 8, 27) {real, imag} */,
  {32'hbfc694a8, 32'hbf97761f} /* (22, 8, 26) {real, imag} */,
  {32'hbf19bdf1, 32'h3e8d598c} /* (22, 8, 25) {real, imag} */,
  {32'hbfbcf396, 32'hbf5b214c} /* (22, 8, 24) {real, imag} */,
  {32'hbfc0b798, 32'hbf8c5896} /* (22, 8, 23) {real, imag} */,
  {32'hbfa7adbc, 32'hbf5f876c} /* (22, 8, 22) {real, imag} */,
  {32'hbf15a22d, 32'hbfe40fd1} /* (22, 8, 21) {real, imag} */,
  {32'hbf0584a0, 32'hbe9e218a} /* (22, 8, 20) {real, imag} */,
  {32'h3f3e6d98, 32'hbfa322b8} /* (22, 8, 19) {real, imag} */,
  {32'h3fc98606, 32'hc00f22bc} /* (22, 8, 18) {real, imag} */,
  {32'h3f2ed381, 32'hbf8a0ae8} /* (22, 8, 17) {real, imag} */,
  {32'hbf3d965e, 32'h3f11a482} /* (22, 8, 16) {real, imag} */,
  {32'h3f92d498, 32'h3fb1855a} /* (22, 8, 15) {real, imag} */,
  {32'h3fd04e02, 32'hbe9491f2} /* (22, 8, 14) {real, imag} */,
  {32'h3f9b351e, 32'h3f180a84} /* (22, 8, 13) {real, imag} */,
  {32'h3f911d4c, 32'h3f9c4944} /* (22, 8, 12) {real, imag} */,
  {32'hbf8feac6, 32'hbfb7bcf0} /* (22, 8, 11) {real, imag} */,
  {32'hc012306e, 32'hbf810557} /* (22, 8, 10) {real, imag} */,
  {32'hbf393f4e, 32'h3f22276c} /* (22, 8, 9) {real, imag} */,
  {32'h3f6cb9b0, 32'hbe89b9ee} /* (22, 8, 8) {real, imag} */,
  {32'h3fb80eac, 32'h3f007964} /* (22, 8, 7) {real, imag} */,
  {32'h3e63ebd8, 32'h3f66854c} /* (22, 8, 6) {real, imag} */,
  {32'hbdddbab0, 32'h3f3710d4} /* (22, 8, 5) {real, imag} */,
  {32'h3fc797c1, 32'hbeccf0d4} /* (22, 8, 4) {real, imag} */,
  {32'h3f9c45be, 32'h3fa19b1e} /* (22, 8, 3) {real, imag} */,
  {32'h3fe0c39a, 32'h3fe65ff7} /* (22, 8, 2) {real, imag} */,
  {32'hbf3317b3, 32'h3fd81cb0} /* (22, 8, 1) {real, imag} */,
  {32'hbfd745f6, 32'h3f304cb8} /* (22, 8, 0) {real, imag} */,
  {32'hbc54f180, 32'hbea7601a} /* (22, 7, 31) {real, imag} */,
  {32'h3fbc2b14, 32'h3ed6b200} /* (22, 7, 30) {real, imag} */,
  {32'h3e89aa88, 32'h3f4d6c06} /* (22, 7, 29) {real, imag} */,
  {32'hbfce2325, 32'h3f208b41} /* (22, 7, 28) {real, imag} */,
  {32'hbf83887b, 32'h3e8271a2} /* (22, 7, 27) {real, imag} */,
  {32'hbf320f76, 32'hbefc35b0} /* (22, 7, 26) {real, imag} */,
  {32'hbe988710, 32'h3f921cf6} /* (22, 7, 25) {real, imag} */,
  {32'h3ede1ff4, 32'h3f2cc06e} /* (22, 7, 24) {real, imag} */,
  {32'h3dbb7cd0, 32'hbeeb7e88} /* (22, 7, 23) {real, imag} */,
  {32'hbf48bd3a, 32'h3dfa3a70} /* (22, 7, 22) {real, imag} */,
  {32'hbf1c294f, 32'h3e19aa18} /* (22, 7, 21) {real, imag} */,
  {32'hbf541860, 32'hbdadb888} /* (22, 7, 20) {real, imag} */,
  {32'h3eebeca8, 32'h3eed4ab4} /* (22, 7, 19) {real, imag} */,
  {32'h3ed0cea2, 32'hbf8e93ce} /* (22, 7, 18) {real, imag} */,
  {32'h3f2c1ae4, 32'hbf3c5374} /* (22, 7, 17) {real, imag} */,
  {32'hbf97a87d, 32'h3f5dce26} /* (22, 7, 16) {real, imag} */,
  {32'hbe956798, 32'h400f5c2e} /* (22, 7, 15) {real, imag} */,
  {32'h400a4b4e, 32'h3f84fa4e} /* (22, 7, 14) {real, imag} */,
  {32'h3f931744, 32'h3fbb0467} /* (22, 7, 13) {real, imag} */,
  {32'hbf25543b, 32'h40106c46} /* (22, 7, 12) {real, imag} */,
  {32'hbe93dc74, 32'hbf51802f} /* (22, 7, 11) {real, imag} */,
  {32'hbf9a61f3, 32'hbf1bbbe4} /* (22, 7, 10) {real, imag} */,
  {32'hbf6203f8, 32'h3f11310a} /* (22, 7, 9) {real, imag} */,
  {32'hbf5488bb, 32'hbdd36210} /* (22, 7, 8) {real, imag} */,
  {32'hbf854184, 32'h3f916b3a} /* (22, 7, 7) {real, imag} */,
  {32'hbe09d36c, 32'h3f6a362e} /* (22, 7, 6) {real, imag} */,
  {32'hbefc83fc, 32'hbcb02480} /* (22, 7, 5) {real, imag} */,
  {32'h3f81492a, 32'hbfc48344} /* (22, 7, 4) {real, imag} */,
  {32'h3eae66f6, 32'h3e4cd5c0} /* (22, 7, 3) {real, imag} */,
  {32'hbf131474, 32'h3edd9a14} /* (22, 7, 2) {real, imag} */,
  {32'h3e643a34, 32'h3fa8c5ed} /* (22, 7, 1) {real, imag} */,
  {32'hbebe25e8, 32'h3f5289ee} /* (22, 7, 0) {real, imag} */,
  {32'h3f11f4d4, 32'hbca92f80} /* (22, 6, 31) {real, imag} */,
  {32'h3f3a3622, 32'h3f49d127} /* (22, 6, 30) {real, imag} */,
  {32'h3f7286fa, 32'h3b7f9a00} /* (22, 6, 29) {real, imag} */,
  {32'hbf3ab2b6, 32'h3e941776} /* (22, 6, 28) {real, imag} */,
  {32'hbed66518, 32'h3fb19032} /* (22, 6, 27) {real, imag} */,
  {32'hbf1495d0, 32'h3f06c3d6} /* (22, 6, 26) {real, imag} */,
  {32'h3e25b428, 32'h3fb4c35f} /* (22, 6, 25) {real, imag} */,
  {32'h3f05c060, 32'h3d09d920} /* (22, 6, 24) {real, imag} */,
  {32'h3f64ae53, 32'hbf575a50} /* (22, 6, 23) {real, imag} */,
  {32'h3d1800d0, 32'hbed695f0} /* (22, 6, 22) {real, imag} */,
  {32'h3f5bd042, 32'hbadff000} /* (22, 6, 21) {real, imag} */,
  {32'h3f571206, 32'hbe99a130} /* (22, 6, 20) {real, imag} */,
  {32'h3fa61d55, 32'h3f2b0cd0} /* (22, 6, 19) {real, imag} */,
  {32'h3f83e7a5, 32'h3e7bec7c} /* (22, 6, 18) {real, imag} */,
  {32'h3fb4a464, 32'h3e8070e6} /* (22, 6, 17) {real, imag} */,
  {32'hbee6605c, 32'h3f94f943} /* (22, 6, 16) {real, imag} */,
  {32'hbe839a9c, 32'h3f34a8d8} /* (22, 6, 15) {real, imag} */,
  {32'h40050340, 32'h3e290ed0} /* (22, 6, 14) {real, imag} */,
  {32'h3e4d04e4, 32'h3f58ee3d} /* (22, 6, 13) {real, imag} */,
  {32'hbf7862ad, 32'h3f5004a5} /* (22, 6, 12) {real, imag} */,
  {32'h3ebbc644, 32'hbf7f4203} /* (22, 6, 11) {real, imag} */,
  {32'h3dc402f0, 32'hbf53c19e} /* (22, 6, 10) {real, imag} */,
  {32'hbfbf5055, 32'hbf3ffba2} /* (22, 6, 9) {real, imag} */,
  {32'hbfb1da66, 32'hbf1661f3} /* (22, 6, 8) {real, imag} */,
  {32'hbfc857cc, 32'hbf4ea0b6} /* (22, 6, 7) {real, imag} */,
  {32'hbf9d4ac9, 32'hbf995898} /* (22, 6, 6) {real, imag} */,
  {32'h3eb0f958, 32'hbfd07b96} /* (22, 6, 5) {real, imag} */,
  {32'h3f66487a, 32'hbff4e378} /* (22, 6, 4) {real, imag} */,
  {32'h3ea88f46, 32'h3d983378} /* (22, 6, 3) {real, imag} */,
  {32'hbf3810ae, 32'h4007ab00} /* (22, 6, 2) {real, imag} */,
  {32'hbf6b1d54, 32'h401862bc} /* (22, 6, 1) {real, imag} */,
  {32'h3bb77e00, 32'h3f4df206} /* (22, 6, 0) {real, imag} */,
  {32'h3dda31b0, 32'hbf23a69c} /* (22, 5, 31) {real, imag} */,
  {32'hbfa63a9c, 32'hbd1b9090} /* (22, 5, 30) {real, imag} */,
  {32'hbf3ff222, 32'hbf4c2400} /* (22, 5, 29) {real, imag} */,
  {32'hbff2a052, 32'hbf060c2e} /* (22, 5, 28) {real, imag} */,
  {32'hbf9bedc7, 32'hbdd52790} /* (22, 5, 27) {real, imag} */,
  {32'hbc759700, 32'hbfbccb5c} /* (22, 5, 26) {real, imag} */,
  {32'h3eee947e, 32'hbe1ceb38} /* (22, 5, 25) {real, imag} */,
  {32'hbfedb6cc, 32'hbfb7fa1f} /* (22, 5, 24) {real, imag} */,
  {32'hbf08303c, 32'hbff7a97a} /* (22, 5, 23) {real, imag} */,
  {32'h3e8fca4c, 32'hbe2cc428} /* (22, 5, 22) {real, imag} */,
  {32'h402abdb8, 32'h3caeabe0} /* (22, 5, 21) {real, imag} */,
  {32'h3fcdb06c, 32'hbf550cee} /* (22, 5, 20) {real, imag} */,
  {32'h3facae82, 32'hbdbe5b36} /* (22, 5, 19) {real, imag} */,
  {32'h3f09e23e, 32'h3e98be1b} /* (22, 5, 18) {real, imag} */,
  {32'h3fead6ec, 32'h3e66aefc} /* (22, 5, 17) {real, imag} */,
  {32'h3c1aab80, 32'h3ed89adc} /* (22, 5, 16) {real, imag} */,
  {32'hbf8a4069, 32'hbf9aa06d} /* (22, 5, 15) {real, imag} */,
  {32'h3fb9e670, 32'hbf92c419} /* (22, 5, 14) {real, imag} */,
  {32'hbe9d00e2, 32'hbf230a32} /* (22, 5, 13) {real, imag} */,
  {32'hbfc3f4b2, 32'hbf113164} /* (22, 5, 12) {real, imag} */,
  {32'hbeead350, 32'h3ebf1f18} /* (22, 5, 11) {real, imag} */,
  {32'h3f9647da, 32'hbec1ba9e} /* (22, 5, 10) {real, imag} */,
  {32'h3f0ed9c0, 32'h3da49984} /* (22, 5, 9) {real, imag} */,
  {32'h3f11c3e2, 32'h3e5faa64} /* (22, 5, 8) {real, imag} */,
  {32'hbe3d5260, 32'hbebc9290} /* (22, 5, 7) {real, imag} */,
  {32'h3f4c66ed, 32'hbfa92a3d} /* (22, 5, 6) {real, imag} */,
  {32'hbd419580, 32'hbf64b8d4} /* (22, 5, 5) {real, imag} */,
  {32'h3e7fc81c, 32'hbfd564a1} /* (22, 5, 4) {real, imag} */,
  {32'hbf2e35af, 32'hbeded8f8} /* (22, 5, 3) {real, imag} */,
  {32'hbfefa419, 32'h4015dd84} /* (22, 5, 2) {real, imag} */,
  {32'hbf8e3469, 32'h400785bb} /* (22, 5, 1) {real, imag} */,
  {32'h3e598a20, 32'h3dd4b0b4} /* (22, 5, 0) {real, imag} */,
  {32'h3dabbd00, 32'hbed3830e} /* (22, 4, 31) {real, imag} */,
  {32'hbf670e29, 32'hbdb00980} /* (22, 4, 30) {real, imag} */,
  {32'hbfce6e22, 32'hbf8093e8} /* (22, 4, 29) {real, imag} */,
  {32'hc0288538, 32'hbf8fa86c} /* (22, 4, 28) {real, imag} */,
  {32'hbfd395cc, 32'hbdd9e010} /* (22, 4, 27) {real, imag} */,
  {32'h3f8dc1ea, 32'hbe7d5290} /* (22, 4, 26) {real, imag} */,
  {32'h3f54d6ee, 32'hbe6af7e8} /* (22, 4, 25) {real, imag} */,
  {32'hbee22dee, 32'hbfb764d8} /* (22, 4, 24) {real, imag} */,
  {32'hbf2bbe6c, 32'hbec844f8} /* (22, 4, 23) {real, imag} */,
  {32'hbe817b60, 32'h3fa8963c} /* (22, 4, 22) {real, imag} */,
  {32'h4006408e, 32'h401bf06f} /* (22, 4, 21) {real, imag} */,
  {32'h3f616f90, 32'h3efaadb0} /* (22, 4, 20) {real, imag} */,
  {32'h3ea1bda4, 32'hbe4e9328} /* (22, 4, 19) {real, imag} */,
  {32'h3f7119b1, 32'hbd334fc0} /* (22, 4, 18) {real, imag} */,
  {32'h3e912594, 32'h3eacee20} /* (22, 4, 17) {real, imag} */,
  {32'hbfba62d9, 32'h3fa43882} /* (22, 4, 16) {real, imag} */,
  {32'hbfa5c83e, 32'h3f1b69e7} /* (22, 4, 15) {real, imag} */,
  {32'h3e2d7bf0, 32'h3f52ef96} /* (22, 4, 14) {real, imag} */,
  {32'h3f704db9, 32'h3f527ae2} /* (22, 4, 13) {real, imag} */,
  {32'h3e6dccc8, 32'hbe1350d8} /* (22, 4, 12) {real, imag} */,
  {32'h3f819e00, 32'h3ba50980} /* (22, 4, 11) {real, imag} */,
  {32'h3f233e3a, 32'hbf0f3976} /* (22, 4, 10) {real, imag} */,
  {32'h3fd673d2, 32'hbf153ca6} /* (22, 4, 9) {real, imag} */,
  {32'h402c24ee, 32'h3f48aef1} /* (22, 4, 8) {real, imag} */,
  {32'h3e235810, 32'h3fbf0670} /* (22, 4, 7) {real, imag} */,
  {32'h3f3cf35b, 32'h3faed8ba} /* (22, 4, 6) {real, imag} */,
  {32'hbe773120, 32'h3f5c1462} /* (22, 4, 5) {real, imag} */,
  {32'hbeae1cfc, 32'hbf95c8b9} /* (22, 4, 4) {real, imag} */,
  {32'hbf200388, 32'hbf5eaed4} /* (22, 4, 3) {real, imag} */,
  {32'hbe7ec5a0, 32'h3c724800} /* (22, 4, 2) {real, imag} */,
  {32'h3f248802, 32'hbef55000} /* (22, 4, 1) {real, imag} */,
  {32'h3f2a72f5, 32'hbf5e2c53} /* (22, 4, 0) {real, imag} */,
  {32'hbeacf858, 32'hbef51b40} /* (22, 3, 31) {real, imag} */,
  {32'hbf5c5da4, 32'hbf81f464} /* (22, 3, 30) {real, imag} */,
  {32'hc009dd28, 32'hbfefd1ab} /* (22, 3, 29) {real, imag} */,
  {32'hbf583c5e, 32'hbf6c7c37} /* (22, 3, 28) {real, imag} */,
  {32'hbf925496, 32'h3f7c3518} /* (22, 3, 27) {real, imag} */,
  {32'hbf9966e4, 32'h3f009ee2} /* (22, 3, 26) {real, imag} */,
  {32'hbf9b1058, 32'hbeddb1a8} /* (22, 3, 25) {real, imag} */,
  {32'hbe55a750, 32'hbf06db85} /* (22, 3, 24) {real, imag} */,
  {32'hbfa81a81, 32'h3e1f7c9c} /* (22, 3, 23) {real, imag} */,
  {32'hbf838d7c, 32'h3f4899d0} /* (22, 3, 22) {real, imag} */,
  {32'hbd85def8, 32'h401970f8} /* (22, 3, 21) {real, imag} */,
  {32'hbfa1e2d1, 32'h3e518be8} /* (22, 3, 20) {real, imag} */,
  {32'hbf5a6bfc, 32'hbfb91649} /* (22, 3, 19) {real, imag} */,
  {32'h3e723eb8, 32'hc02278bc} /* (22, 3, 18) {real, imag} */,
  {32'h3ec49f74, 32'hbf536240} /* (22, 3, 17) {real, imag} */,
  {32'hbee3aaa8, 32'h3e410150} /* (22, 3, 16) {real, imag} */,
  {32'hbe3c0f22, 32'h40089e5f} /* (22, 3, 15) {real, imag} */,
  {32'hbf26ae35, 32'h4008e944} /* (22, 3, 14) {real, imag} */,
  {32'h3f45c336, 32'h3f77011e} /* (22, 3, 13) {real, imag} */,
  {32'h3fd94dd0, 32'h3f0c6716} /* (22, 3, 12) {real, imag} */,
  {32'h3f1f42ca, 32'h3d86d3b0} /* (22, 3, 11) {real, imag} */,
  {32'h3f6a5c7a, 32'h3f6a97a2} /* (22, 3, 10) {real, imag} */,
  {32'h3f291af0, 32'h3f63d523} /* (22, 3, 9) {real, imag} */,
  {32'h3faa6b83, 32'h3bbe3b00} /* (22, 3, 8) {real, imag} */,
  {32'h3f494c48, 32'hbe6c5d50} /* (22, 3, 7) {real, imag} */,
  {32'h3fc62da6, 32'h3f9e9aa3} /* (22, 3, 6) {real, imag} */,
  {32'h3e8f2f5b, 32'h3f824d25} /* (22, 3, 5) {real, imag} */,
  {32'hbf19779e, 32'hbd9ec4f0} /* (22, 3, 4) {real, imag} */,
  {32'hbeb76044, 32'hbd325980} /* (22, 3, 3) {real, imag} */,
  {32'hbf14ecdc, 32'h3f3eaf1e} /* (22, 3, 2) {real, imag} */,
  {32'h3ade3800, 32'hbf0170e0} /* (22, 3, 1) {real, imag} */,
  {32'h3ec30688, 32'hbf5a3af6} /* (22, 3, 0) {real, imag} */,
  {32'hbf05ee4e, 32'hbf1d86b1} /* (22, 2, 31) {real, imag} */,
  {32'hbf71762d, 32'hbd9f1fe0} /* (22, 2, 30) {real, imag} */,
  {32'hbf244812, 32'h3d1e4060} /* (22, 2, 29) {real, imag} */,
  {32'hbd476a00, 32'hbf089b8a} /* (22, 2, 28) {real, imag} */,
  {32'hbe5e5e30, 32'hbf5c4776} /* (22, 2, 27) {real, imag} */,
  {32'hbf20dc36, 32'hbf7a17d0} /* (22, 2, 26) {real, imag} */,
  {32'h3e935108, 32'hbfc45b3c} /* (22, 2, 25) {real, imag} */,
  {32'hbddae8a0, 32'hbfcebbb6} /* (22, 2, 24) {real, imag} */,
  {32'hbfa138cf, 32'hbf145f80} /* (22, 2, 23) {real, imag} */,
  {32'h3e21fe00, 32'hbe74d9bc} /* (22, 2, 22) {real, imag} */,
  {32'h3f4496a4, 32'h400efc95} /* (22, 2, 21) {real, imag} */,
  {32'hbd83a020, 32'h3ef558c0} /* (22, 2, 20) {real, imag} */,
  {32'h3e279500, 32'hbf0c2b58} /* (22, 2, 19) {real, imag} */,
  {32'h3f9eecfa, 32'hc001f343} /* (22, 2, 18) {real, imag} */,
  {32'h3f80478d, 32'hbface948} /* (22, 2, 17) {real, imag} */,
  {32'h3f0efe85, 32'hbff6b654} /* (22, 2, 16) {real, imag} */,
  {32'h3f734a8c, 32'h3e84befc} /* (22, 2, 15) {real, imag} */,
  {32'h3ee5f5a8, 32'h3f9644da} /* (22, 2, 14) {real, imag} */,
  {32'h3e5b7480, 32'h401763f1} /* (22, 2, 13) {real, imag} */,
  {32'h3f259ad9, 32'h3f8dea09} /* (22, 2, 12) {real, imag} */,
  {32'hbe0ca7b8, 32'h3c31c480} /* (22, 2, 11) {real, imag} */,
  {32'h3f51ab5c, 32'h3f7ec7fa} /* (22, 2, 10) {real, imag} */,
  {32'h3fd597bb, 32'h3dc6aa40} /* (22, 2, 9) {real, imag} */,
  {32'h3f4cf798, 32'hbf81f829} /* (22, 2, 8) {real, imag} */,
  {32'h3f66462d, 32'hbfa263c6} /* (22, 2, 7) {real, imag} */,
  {32'h40006778, 32'h3e831b14} /* (22, 2, 6) {real, imag} */,
  {32'h3f2616b4, 32'hbe44b870} /* (22, 2, 5) {real, imag} */,
  {32'hbd6c1700, 32'hbf1a9fb8} /* (22, 2, 4) {real, imag} */,
  {32'hbf9b574a, 32'hbe1f2adc} /* (22, 2, 3) {real, imag} */,
  {32'hbfe5cb1e, 32'h3f425448} /* (22, 2, 2) {real, imag} */,
  {32'hbe80a05c, 32'h3d807ab0} /* (22, 2, 1) {real, imag} */,
  {32'h3ef99e8c, 32'hbf7c6a8e} /* (22, 2, 0) {real, imag} */,
  {32'hbecb41e8, 32'hbd0c3340} /* (22, 1, 31) {real, imag} */,
  {32'hbfbb6524, 32'h3f28ba26} /* (22, 1, 30) {real, imag} */,
  {32'hbf77ac35, 32'h3f2b934c} /* (22, 1, 29) {real, imag} */,
  {32'hbf37e950, 32'h3f02f17e} /* (22, 1, 28) {real, imag} */,
  {32'h3dfd02e0, 32'hbf0d1caa} /* (22, 1, 27) {real, imag} */,
  {32'h3ec4e11e, 32'h3f3040ee} /* (22, 1, 26) {real, imag} */,
  {32'hbe985fd8, 32'h3e87b6f4} /* (22, 1, 25) {real, imag} */,
  {32'hbf482348, 32'hbfafaf33} /* (22, 1, 24) {real, imag} */,
  {32'h3e81539c, 32'hc0019ff2} /* (22, 1, 23) {real, imag} */,
  {32'hbdb0c778, 32'hbe8d9a06} /* (22, 1, 22) {real, imag} */,
  {32'h3e551abc, 32'h3fc0ccf4} /* (22, 1, 21) {real, imag} */,
  {32'h3fa987c2, 32'h3f720816} /* (22, 1, 20) {real, imag} */,
  {32'h3f5585c8, 32'h3ef2ba08} /* (22, 1, 19) {real, imag} */,
  {32'h3fe6ae4c, 32'hbf47d9ec} /* (22, 1, 18) {real, imag} */,
  {32'h3f849cc9, 32'hbeddd1ba} /* (22, 1, 17) {real, imag} */,
  {32'hbf135e6e, 32'hbf5ab1d7} /* (22, 1, 16) {real, imag} */,
  {32'h3eb55fde, 32'h3dc38d18} /* (22, 1, 15) {real, imag} */,
  {32'h3eb5a838, 32'h3fc0262a} /* (22, 1, 14) {real, imag} */,
  {32'hbfa6bbdc, 32'h40224760} /* (22, 1, 13) {real, imag} */,
  {32'hbf2d6b40, 32'h3f818ac4} /* (22, 1, 12) {real, imag} */,
  {32'hbf55b784, 32'hbf46ae70} /* (22, 1, 11) {real, imag} */,
  {32'h3daf4d48, 32'hbcbf9cc0} /* (22, 1, 10) {real, imag} */,
  {32'h3fd9f11c, 32'h3f79acd8} /* (22, 1, 9) {real, imag} */,
  {32'h4033b35c, 32'h3ed1f3b4} /* (22, 1, 8) {real, imag} */,
  {32'h3fec0585, 32'h3f102b86} /* (22, 1, 7) {real, imag} */,
  {32'h3f953466, 32'h3f3c0372} /* (22, 1, 6) {real, imag} */,
  {32'h3fbb206c, 32'hbf82535b} /* (22, 1, 5) {real, imag} */,
  {32'h3fa5821f, 32'hbfc21db5} /* (22, 1, 4) {real, imag} */,
  {32'hbe7d7464, 32'h3ef50784} /* (22, 1, 3) {real, imag} */,
  {32'hbed6eb27, 32'h3fcbb2d1} /* (22, 1, 2) {real, imag} */,
  {32'hbeef66e6, 32'h3f1f844d} /* (22, 1, 1) {real, imag} */,
  {32'hbefe8de6, 32'hbdd0c8c0} /* (22, 1, 0) {real, imag} */,
  {32'h3e43bc7c, 32'h3e405bfc} /* (22, 0, 31) {real, imag} */,
  {32'hbec3235e, 32'h3ea03d36} /* (22, 0, 30) {real, imag} */,
  {32'hbf932f3b, 32'h3e8d05f0} /* (22, 0, 29) {real, imag} */,
  {32'hbf2d9b50, 32'h3e9a62b0} /* (22, 0, 28) {real, imag} */,
  {32'h3ed1b1b6, 32'h3ebd24ca} /* (22, 0, 27) {real, imag} */,
  {32'hbe2f8aa0, 32'h3f581b7d} /* (22, 0, 26) {real, imag} */,
  {32'hbfbdda10, 32'hbe27b36a} /* (22, 0, 25) {real, imag} */,
  {32'hbfc39a24, 32'hbfa79822} /* (22, 0, 24) {real, imag} */,
  {32'h3dd486f0, 32'hc01c57ee} /* (22, 0, 23) {real, imag} */,
  {32'hbf3dab2a, 32'hbf3a46c6} /* (22, 0, 22) {real, imag} */,
  {32'h3d910034, 32'hbda6bde0} /* (22, 0, 21) {real, imag} */,
  {32'h3fd579ec, 32'h3ef1fff0} /* (22, 0, 20) {real, imag} */,
  {32'h3ec5e580, 32'h3ebb336e} /* (22, 0, 19) {real, imag} */,
  {32'h3f211942, 32'h3f4b0ddd} /* (22, 0, 18) {real, imag} */,
  {32'h3f60dd5c, 32'h3f8f6462} /* (22, 0, 17) {real, imag} */,
  {32'hbf42b574, 32'h3d615b84} /* (22, 0, 16) {real, imag} */,
  {32'h3ed1663d, 32'h3f869221} /* (22, 0, 15) {real, imag} */,
  {32'h3fbf31fa, 32'h3fa35cd6} /* (22, 0, 14) {real, imag} */,
  {32'hbee925ec, 32'h3f4f0a64} /* (22, 0, 13) {real, imag} */,
  {32'hbf6b74e9, 32'h3e604bac} /* (22, 0, 12) {real, imag} */,
  {32'hbe7c1140, 32'hbdaf3f40} /* (22, 0, 11) {real, imag} */,
  {32'hbe3c47e8, 32'h3e09e56c} /* (22, 0, 10) {real, imag} */,
  {32'h3f207bf3, 32'h3f1d51bc} /* (22, 0, 9) {real, imag} */,
  {32'h400271d4, 32'h3ec218d0} /* (22, 0, 8) {real, imag} */,
  {32'h3fd56fbb, 32'hbcf67400} /* (22, 0, 7) {real, imag} */,
  {32'h3f743424, 32'hbea47924} /* (22, 0, 6) {real, imag} */,
  {32'h3f7c4c76, 32'hbf751019} /* (22, 0, 5) {real, imag} */,
  {32'h3f622764, 32'hbf88afbd} /* (22, 0, 4) {real, imag} */,
  {32'hbe979f46, 32'h3e15c85c} /* (22, 0, 3) {real, imag} */,
  {32'hbe482338, 32'h3f4d17b7} /* (22, 0, 2) {real, imag} */,
  {32'h3d0bb540, 32'h3fab0aa6} /* (22, 0, 1) {real, imag} */,
  {32'h3e5a14a6, 32'h3eb894c0} /* (22, 0, 0) {real, imag} */,
  {32'h3ee45ab2, 32'h3e8936a6} /* (21, 31, 31) {real, imag} */,
  {32'h3e8e9cac, 32'h3f173560} /* (21, 31, 30) {real, imag} */,
  {32'hbee079ac, 32'hbe4de958} /* (21, 31, 29) {real, imag} */,
  {32'hbeb8fd02, 32'hbf439618} /* (21, 31, 28) {real, imag} */,
  {32'h3eb3fba8, 32'hbfd2f65c} /* (21, 31, 27) {real, imag} */,
  {32'h3e1b6a38, 32'hbf72d37c} /* (21, 31, 26) {real, imag} */,
  {32'hbf25ad96, 32'h3e96a1e8} /* (21, 31, 25) {real, imag} */,
  {32'h3f26a079, 32'hbdf2ed50} /* (21, 31, 24) {real, imag} */,
  {32'h3ec7c1a1, 32'h3f32f827} /* (21, 31, 23) {real, imag} */,
  {32'h3e302226, 32'h3e769e50} /* (21, 31, 22) {real, imag} */,
  {32'hbeadcf8c, 32'hbe592114} /* (21, 31, 21) {real, imag} */,
  {32'hbef994a8, 32'hbf36dc53} /* (21, 31, 20) {real, imag} */,
  {32'hbf02ec64, 32'hbeef592e} /* (21, 31, 19) {real, imag} */,
  {32'hbf15bbdd, 32'h3e1de9f8} /* (21, 31, 18) {real, imag} */,
  {32'hbed98b07, 32'h3e3008b8} /* (21, 31, 17) {real, imag} */,
  {32'hbe920715, 32'hbe787330} /* (21, 31, 16) {real, imag} */,
  {32'h3e0b9170, 32'hbd051246} /* (21, 31, 15) {real, imag} */,
  {32'h3e46c07e, 32'hbd4de050} /* (21, 31, 14) {real, imag} */,
  {32'hbe968b28, 32'hbfc3a1d4} /* (21, 31, 13) {real, imag} */,
  {32'hbef87b80, 32'hbfc613d4} /* (21, 31, 12) {real, imag} */,
  {32'h3e2915ee, 32'hbc858460} /* (21, 31, 11) {real, imag} */,
  {32'h3f2afa57, 32'hbf354702} /* (21, 31, 10) {real, imag} */,
  {32'h3db02f00, 32'hbdec6648} /* (21, 31, 9) {real, imag} */,
  {32'h3d532920, 32'h3e07ee2e} /* (21, 31, 8) {real, imag} */,
  {32'h3ec11dc0, 32'h3e179ddc} /* (21, 31, 7) {real, imag} */,
  {32'h3ee8b938, 32'h3f35a900} /* (21, 31, 6) {real, imag} */,
  {32'h3f4c918e, 32'h3f405ec5} /* (21, 31, 5) {real, imag} */,
  {32'h3dbcff0c, 32'h3f4a931c} /* (21, 31, 4) {real, imag} */,
  {32'h3f218dce, 32'h3f0d5cf0} /* (21, 31, 3) {real, imag} */,
  {32'h3f6d74f2, 32'h3f796c86} /* (21, 31, 2) {real, imag} */,
  {32'h3fa3058c, 32'h3f9f9275} /* (21, 31, 1) {real, imag} */,
  {32'h3fa11899, 32'h3d74efb4} /* (21, 31, 0) {real, imag} */,
  {32'hbd95a150, 32'hbe9964ad} /* (21, 30, 31) {real, imag} */,
  {32'h3f6e7b04, 32'h3f772adc} /* (21, 30, 30) {real, imag} */,
  {32'h3e8084c0, 32'h3fa57734} /* (21, 30, 29) {real, imag} */,
  {32'h3ce10540, 32'h3e96b160} /* (21, 30, 28) {real, imag} */,
  {32'h3f5c04d8, 32'hbfa44d9a} /* (21, 30, 27) {real, imag} */,
  {32'h3f9a62e2, 32'hbfa159d2} /* (21, 30, 26) {real, imag} */,
  {32'hbeaf43f4, 32'h3f0a9096} /* (21, 30, 25) {real, imag} */,
  {32'h3e9fc3e0, 32'h3f87fdf0} /* (21, 30, 24) {real, imag} */,
  {32'h3f19681b, 32'h3ff98378} /* (21, 30, 23) {real, imag} */,
  {32'h3e0db840, 32'h3fb71e36} /* (21, 30, 22) {real, imag} */,
  {32'hbed42814, 32'hbe13f7fa} /* (21, 30, 21) {real, imag} */,
  {32'hbf16afec, 32'hbfc5e5ea} /* (21, 30, 20) {real, imag} */,
  {32'h3ed9c9b8, 32'hbf6553ea} /* (21, 30, 19) {real, imag} */,
  {32'h3e05e064, 32'h3c89b4c0} /* (21, 30, 18) {real, imag} */,
  {32'hbf8f2f3e, 32'h3dd25640} /* (21, 30, 17) {real, imag} */,
  {32'hbe7ce174, 32'hbf605f18} /* (21, 30, 16) {real, imag} */,
  {32'hbeb20a0a, 32'hbd67a600} /* (21, 30, 15) {real, imag} */,
  {32'hbf2343ed, 32'hbe726970} /* (21, 30, 14) {real, imag} */,
  {32'hbeeea3fa, 32'hbfe8f199} /* (21, 30, 13) {real, imag} */,
  {32'h3e26024c, 32'hbfa3993a} /* (21, 30, 12) {real, imag} */,
  {32'h3f939a80, 32'h3f78a0b0} /* (21, 30, 11) {real, imag} */,
  {32'h3fa4bab2, 32'h3efe11c1} /* (21, 30, 10) {real, imag} */,
  {32'hbdfecbb0, 32'h3ea90070} /* (21, 30, 9) {real, imag} */,
  {32'hbec86df4, 32'h3f397df8} /* (21, 30, 8) {real, imag} */,
  {32'h3f8220f4, 32'h3dc8f0e0} /* (21, 30, 7) {real, imag} */,
  {32'h3f6186a2, 32'h3f51d9e8} /* (21, 30, 6) {real, imag} */,
  {32'h3fa00103, 32'h3fcf96e4} /* (21, 30, 5) {real, imag} */,
  {32'h3e39cc25, 32'h3fb602a5} /* (21, 30, 4) {real, imag} */,
  {32'h3ed04a18, 32'h3f5ccfad} /* (21, 30, 3) {real, imag} */,
  {32'h3f386d50, 32'h3fbbd2ad} /* (21, 30, 2) {real, imag} */,
  {32'h3ffd6ebc, 32'h3f969c81} /* (21, 30, 1) {real, imag} */,
  {32'h3ff70deb, 32'h3e9c2aca} /* (21, 30, 0) {real, imag} */,
  {32'h3e8082ee, 32'hbf983ccf} /* (21, 29, 31) {real, imag} */,
  {32'h3f8711fe, 32'hbdf6ffb0} /* (21, 29, 30) {real, imag} */,
  {32'h3e1891b8, 32'h3fb0e621} /* (21, 29, 29) {real, imag} */,
  {32'h3f48f2c6, 32'h3fc622f0} /* (21, 29, 28) {real, imag} */,
  {32'h3fc69619, 32'h3fddb2e9} /* (21, 29, 27) {real, imag} */,
  {32'h3ee79fc2, 32'h3f9fd406} /* (21, 29, 26) {real, imag} */,
  {32'hbf8db9fa, 32'h3fccfb96} /* (21, 29, 25) {real, imag} */,
  {32'h3f8bb6ea, 32'h4015971e} /* (21, 29, 24) {real, imag} */,
  {32'h4033e720, 32'h3fdf2600} /* (21, 29, 23) {real, imag} */,
  {32'h3fa0e10d, 32'h3ffb8452} /* (21, 29, 22) {real, imag} */,
  {32'h3f36cf72, 32'h3fdec9d2} /* (21, 29, 21) {real, imag} */,
  {32'hbdbb9ff8, 32'h3e335380} /* (21, 29, 20) {real, imag} */,
  {32'h3f39c7f0, 32'hbf0093b0} /* (21, 29, 19) {real, imag} */,
  {32'hbeaf6ee8, 32'h3e5b2460} /* (21, 29, 18) {real, imag} */,
  {32'hbf69503a, 32'h3e7649c8} /* (21, 29, 17) {real, imag} */,
  {32'hbf02ed78, 32'hbf0d99d4} /* (21, 29, 16) {real, imag} */,
  {32'hbf99ed94, 32'hbeed0634} /* (21, 29, 15) {real, imag} */,
  {32'hc00e6094, 32'hbf232408} /* (21, 29, 14) {real, imag} */,
  {32'hbff43262, 32'hbf3b1af1} /* (21, 29, 13) {real, imag} */,
  {32'h3dd371c0, 32'h3f0afc96} /* (21, 29, 12) {real, imag} */,
  {32'h3f8cad34, 32'h3f8e26dd} /* (21, 29, 11) {real, imag} */,
  {32'h3fb5cc9f, 32'h3d32d090} /* (21, 29, 10) {real, imag} */,
  {32'h3f700bb8, 32'h3f29ec0e} /* (21, 29, 9) {real, imag} */,
  {32'h3f86b129, 32'h3f53a6a2} /* (21, 29, 8) {real, imag} */,
  {32'h3f82eeb2, 32'h3f26a014} /* (21, 29, 7) {real, imag} */,
  {32'h3fd1a26d, 32'h3facfce9} /* (21, 29, 6) {real, imag} */,
  {32'h3fc7c7db, 32'h3fa3cda4} /* (21, 29, 5) {real, imag} */,
  {32'h3ec69448, 32'h3f2d33c0} /* (21, 29, 4) {real, imag} */,
  {32'hbc8480b0, 32'h3ee3ad08} /* (21, 29, 3) {real, imag} */,
  {32'h3e13d660, 32'h3f0d33a1} /* (21, 29, 2) {real, imag} */,
  {32'h3f9d7eb2, 32'hbf123fe2} /* (21, 29, 1) {real, imag} */,
  {32'h3f381d4e, 32'hbf4c9438} /* (21, 29, 0) {real, imag} */,
  {32'h3f18d2ae, 32'h3ebe2b5a} /* (21, 28, 31) {real, imag} */,
  {32'h3fc5e3d2, 32'h3fbd48ae} /* (21, 28, 30) {real, imag} */,
  {32'h3f11c2a8, 32'h3fac67f8} /* (21, 28, 29) {real, imag} */,
  {32'h3eabf93e, 32'h3f9b7eff} /* (21, 28, 28) {real, imag} */,
  {32'h3fb7536e, 32'h4003c887} /* (21, 28, 27) {real, imag} */,
  {32'h3f71aa41, 32'h3faa6d69} /* (21, 28, 26) {real, imag} */,
  {32'h3f14362e, 32'h3fb3aad5} /* (21, 28, 25) {real, imag} */,
  {32'h3ffbc480, 32'h40168567} /* (21, 28, 24) {real, imag} */,
  {32'h403b3f82, 32'h3fa9911b} /* (21, 28, 23) {real, imag} */,
  {32'h3fe20faf, 32'h3eb7c7b6} /* (21, 28, 22) {real, imag} */,
  {32'h3f055d50, 32'hbe785980} /* (21, 28, 21) {real, imag} */,
  {32'hbfd70469, 32'hbec97024} /* (21, 28, 20) {real, imag} */,
  {32'hbf82edff, 32'hbf192bb6} /* (21, 28, 19) {real, imag} */,
  {32'hc008f4ae, 32'hbf52150c} /* (21, 28, 18) {real, imag} */,
  {32'hbf618b99, 32'hbf2687b2} /* (21, 28, 17) {real, imag} */,
  {32'hbf24908c, 32'hbd9ecaa0} /* (21, 28, 16) {real, imag} */,
  {32'hbfae7ab9, 32'hbe1f0ae8} /* (21, 28, 15) {real, imag} */,
  {32'hbfa437e5, 32'h3e1ca394} /* (21, 28, 14) {real, imag} */,
  {32'hc001e644, 32'hbea640ac} /* (21, 28, 13) {real, imag} */,
  {32'hbdbf7838, 32'h3e9b664a} /* (21, 28, 12) {real, imag} */,
  {32'h3f20e36a, 32'h3f84a656} /* (21, 28, 11) {real, imag} */,
  {32'h3fc28e14, 32'hbeaf78e8} /* (21, 28, 10) {real, imag} */,
  {32'h400efa56, 32'h3e6b53b0} /* (21, 28, 9) {real, imag} */,
  {32'h40148e14, 32'h3f776fc6} /* (21, 28, 8) {real, imag} */,
  {32'h3f7f0278, 32'h3fa1dde6} /* (21, 28, 7) {real, imag} */,
  {32'h3fc404d0, 32'h3f82a731} /* (21, 28, 6) {real, imag} */,
  {32'h3f2e072e, 32'h3fe8cbe1} /* (21, 28, 5) {real, imag} */,
  {32'h3ee0bc1a, 32'h3f15d824} /* (21, 28, 4) {real, imag} */,
  {32'h3f6f0ffc, 32'h3e95ad84} /* (21, 28, 3) {real, imag} */,
  {32'h3ee9d1d8, 32'hbd30e0c0} /* (21, 28, 2) {real, imag} */,
  {32'h3f9d4284, 32'hbf3715d2} /* (21, 28, 1) {real, imag} */,
  {32'h3f7b836d, 32'hbf5de384} /* (21, 28, 0) {real, imag} */,
  {32'hbde5e940, 32'h3f617af3} /* (21, 27, 31) {real, imag} */,
  {32'h3e375584, 32'h3fc3469a} /* (21, 27, 30) {real, imag} */,
  {32'hbeefd996, 32'h3f40eafa} /* (21, 27, 29) {real, imag} */,
  {32'h3e048780, 32'h3f96b61a} /* (21, 27, 28) {real, imag} */,
  {32'h3f004ef8, 32'h402aa90a} /* (21, 27, 27) {real, imag} */,
  {32'h3e1b4a0c, 32'h3f06e286} /* (21, 27, 26) {real, imag} */,
  {32'h4006a890, 32'h3f65ad54} /* (21, 27, 25) {real, imag} */,
  {32'h40022b4e, 32'h3fc4eef2} /* (21, 27, 24) {real, imag} */,
  {32'h3f043e3d, 32'h3d99e808} /* (21, 27, 23) {real, imag} */,
  {32'hb96fa000, 32'hbed3b442} /* (21, 27, 22) {real, imag} */,
  {32'hbe100574, 32'hbee2e944} /* (21, 27, 21) {real, imag} */,
  {32'hc03caab7, 32'hbf96167c} /* (21, 27, 20) {real, imag} */,
  {32'hc03709b7, 32'hbf83d387} /* (21, 27, 19) {real, imag} */,
  {32'hbff6313b, 32'hbf6007b6} /* (21, 27, 18) {real, imag} */,
  {32'hbef16480, 32'hbfb95b90} /* (21, 27, 17) {real, imag} */,
  {32'hbf190a0a, 32'hbf9d5a98} /* (21, 27, 16) {real, imag} */,
  {32'hbfc14ad2, 32'hbf661717} /* (21, 27, 15) {real, imag} */,
  {32'hbf749827, 32'h3f20bd6d} /* (21, 27, 14) {real, imag} */,
  {32'hbf42024c, 32'hbf3e1cdb} /* (21, 27, 13) {real, imag} */,
  {32'hbe211440, 32'hbf1f3c54} /* (21, 27, 12) {real, imag} */,
  {32'h3f18b91d, 32'hbce8cf80} /* (21, 27, 11) {real, imag} */,
  {32'h3f3f320c, 32'h3e337548} /* (21, 27, 10) {real, imag} */,
  {32'h3fdee510, 32'h3f8f4461} /* (21, 27, 9) {real, imag} */,
  {32'h40171e96, 32'h3d9ae770} /* (21, 27, 8) {real, imag} */,
  {32'h3fabe143, 32'h3f3d1526} /* (21, 27, 7) {real, imag} */,
  {32'h3ff9c2f8, 32'h3f5d9545} /* (21, 27, 6) {real, imag} */,
  {32'h3f3b9f73, 32'h3fcf5473} /* (21, 27, 5) {real, imag} */,
  {32'hbdacc2ac, 32'h3e9317a8} /* (21, 27, 4) {real, imag} */,
  {32'h3f80cb62, 32'h3f78b7f2} /* (21, 27, 3) {real, imag} */,
  {32'h3f03b86e, 32'h3f0c2b87} /* (21, 27, 2) {real, imag} */,
  {32'h3f8bd1a7, 32'hbe1b1bac} /* (21, 27, 1) {real, imag} */,
  {32'h3f82109c, 32'h3e6cf8d0} /* (21, 27, 0) {real, imag} */,
  {32'hbe68a545, 32'h3f0a7cf3} /* (21, 26, 31) {real, imag} */,
  {32'hbc98cda0, 32'h3f0ab17e} /* (21, 26, 30) {real, imag} */,
  {32'h3ea6e394, 32'h3fa23c9a} /* (21, 26, 29) {real, imag} */,
  {32'h3fc1b45d, 32'h3ff15f35} /* (21, 26, 28) {real, imag} */,
  {32'h3e294f88, 32'h3f3002f2} /* (21, 26, 27) {real, imag} */,
  {32'hbf89090e, 32'hbf12bdb4} /* (21, 26, 26) {real, imag} */,
  {32'h3ebe8b58, 32'h3e0959b0} /* (21, 26, 25) {real, imag} */,
  {32'h3f89d005, 32'hbf0b0858} /* (21, 26, 24) {real, imag} */,
  {32'hbee664bc, 32'hbee8b401} /* (21, 26, 23) {real, imag} */,
  {32'hbf60eed8, 32'h3f2aa017} /* (21, 26, 22) {real, imag} */,
  {32'h3e927f4a, 32'h3b94c300} /* (21, 26, 21) {real, imag} */,
  {32'hbf803992, 32'hbfbdde43} /* (21, 26, 20) {real, imag} */,
  {32'hbf393fa7, 32'hbf30feac} /* (21, 26, 19) {real, imag} */,
  {32'hbeab8cd8, 32'hbf1362e2} /* (21, 26, 18) {real, imag} */,
  {32'hbf5f2076, 32'hbf7b7786} /* (21, 26, 17) {real, imag} */,
  {32'h3e3e40c8, 32'h3de9ccb0} /* (21, 26, 16) {real, imag} */,
  {32'h3ec58c1c, 32'hbf232f8f} /* (21, 26, 15) {real, imag} */,
  {32'hbf4057c5, 32'hbe6efac8} /* (21, 26, 14) {real, imag} */,
  {32'hbf77ee08, 32'hbf589418} /* (21, 26, 13) {real, imag} */,
  {32'h3d9fd970, 32'hbf96ef60} /* (21, 26, 12) {real, imag} */,
  {32'h3d7cf100, 32'hbf30a2d2} /* (21, 26, 11) {real, imag} */,
  {32'h3c83bbac, 32'h3f15bf5d} /* (21, 26, 10) {real, imag} */,
  {32'h3fc00e23, 32'h3f83800c} /* (21, 26, 9) {real, imag} */,
  {32'h3f0155b6, 32'hbe21dcc0} /* (21, 26, 8) {real, imag} */,
  {32'hbe312e13, 32'h3e427ff4} /* (21, 26, 7) {real, imag} */,
  {32'h3f84890a, 32'h3f70ff14} /* (21, 26, 6) {real, imag} */,
  {32'h3f0c6992, 32'hbea41468} /* (21, 26, 5) {real, imag} */,
  {32'h3f3f4550, 32'hbfab62db} /* (21, 26, 4) {real, imag} */,
  {32'h3f551129, 32'h3f0cbd06} /* (21, 26, 3) {real, imag} */,
  {32'h3f179328, 32'h3f54fe7c} /* (21, 26, 2) {real, imag} */,
  {32'h3f905488, 32'h3e0e9db4} /* (21, 26, 1) {real, imag} */,
  {32'h3ee04ef4, 32'h3ee4fe28} /* (21, 26, 0) {real, imag} */,
  {32'h3f1345e9, 32'h3f46bf10} /* (21, 25, 31) {real, imag} */,
  {32'h3f5adc6f, 32'h3fd7345c} /* (21, 25, 30) {real, imag} */,
  {32'h3f3a4a47, 32'h3f676a74} /* (21, 25, 29) {real, imag} */,
  {32'h3f60c138, 32'h3e8ba794} /* (21, 25, 28) {real, imag} */,
  {32'h3e77bfd8, 32'hbf350b3a} /* (21, 25, 27) {real, imag} */,
  {32'h3cb9cd80, 32'hbf228160} /* (21, 25, 26) {real, imag} */,
  {32'h3f4bd0a0, 32'hbe87275c} /* (21, 25, 25) {real, imag} */,
  {32'h3fd10f49, 32'h3e54bea0} /* (21, 25, 24) {real, imag} */,
  {32'h3f70e3cc, 32'h3e9e2150} /* (21, 25, 23) {real, imag} */,
  {32'h3eb1f56c, 32'h3f06313a} /* (21, 25, 22) {real, imag} */,
  {32'h3e81515a, 32'hbda20670} /* (21, 25, 21) {real, imag} */,
  {32'hbecbc510, 32'hbf132394} /* (21, 25, 20) {real, imag} */,
  {32'h3f1e9691, 32'h3f99a2ff} /* (21, 25, 19) {real, imag} */,
  {32'hbf152d2c, 32'h3f08de1e} /* (21, 25, 18) {real, imag} */,
  {32'hbf844669, 32'hbe788528} /* (21, 25, 17) {real, imag} */,
  {32'h3abf2800, 32'hbea09b26} /* (21, 25, 16) {real, imag} */,
  {32'hbe81803c, 32'hbf3a3170} /* (21, 25, 15) {real, imag} */,
  {32'h3ec57fb4, 32'hbfa5d3da} /* (21, 25, 14) {real, imag} */,
  {32'hbe8c2b34, 32'hbf8fa748} /* (21, 25, 13) {real, imag} */,
  {32'h3f842e48, 32'hbf5c9dca} /* (21, 25, 12) {real, imag} */,
  {32'hbede9610, 32'hbf99d17e} /* (21, 25, 11) {real, imag} */,
  {32'h3c061e40, 32'h3ef0b660} /* (21, 25, 10) {real, imag} */,
  {32'h3f9f0067, 32'h3ec4add0} /* (21, 25, 9) {real, imag} */,
  {32'hbdb17690, 32'h3e570120} /* (21, 25, 8) {real, imag} */,
  {32'hbf06fcb0, 32'h3dd34b60} /* (21, 25, 7) {real, imag} */,
  {32'h3f2e605e, 32'h3fc8c380} /* (21, 25, 6) {real, imag} */,
  {32'h3ecb9f1c, 32'hbf8598c9} /* (21, 25, 5) {real, imag} */,
  {32'h3f8851fc, 32'hc0127ca1} /* (21, 25, 4) {real, imag} */,
  {32'h3f4639b6, 32'h3d8b9df0} /* (21, 25, 3) {real, imag} */,
  {32'h3f9a02d4, 32'h3fcd7f15} /* (21, 25, 2) {real, imag} */,
  {32'h401fbd90, 32'h3e4aa3e0} /* (21, 25, 1) {real, imag} */,
  {32'h3f91523e, 32'h3d2599f0} /* (21, 25, 0) {real, imag} */,
  {32'h3fa67ca4, 32'h3f132782} /* (21, 24, 31) {real, imag} */,
  {32'h3f97dda3, 32'h3fb6c9d8} /* (21, 24, 30) {real, imag} */,
  {32'h3e9c15e4, 32'h3fbb6601} /* (21, 24, 29) {real, imag} */,
  {32'hbf58dab4, 32'h3d1473c0} /* (21, 24, 28) {real, imag} */,
  {32'h3e215d60, 32'h3ec83870} /* (21, 24, 27) {real, imag} */,
  {32'h3f126848, 32'h3e325c10} /* (21, 24, 26) {real, imag} */,
  {32'h3faeadb4, 32'h3d24d880} /* (21, 24, 25) {real, imag} */,
  {32'h4000bc82, 32'hbf02c9c0} /* (21, 24, 24) {real, imag} */,
  {32'h3fc45684, 32'h3f7c32e8} /* (21, 24, 23) {real, imag} */,
  {32'h3e8c4bf0, 32'h3fa0cf5b} /* (21, 24, 22) {real, imag} */,
  {32'hbf1a5884, 32'h3e84ac00} /* (21, 24, 21) {real, imag} */,
  {32'hbf65bb9a, 32'hbeff481e} /* (21, 24, 20) {real, imag} */,
  {32'hbfd36352, 32'h3f91f7fa} /* (21, 24, 19) {real, imag} */,
  {32'hbfec64ec, 32'h3fbc0e1e} /* (21, 24, 18) {real, imag} */,
  {32'hbf8dbd60, 32'h3ef0ce1e} /* (21, 24, 17) {real, imag} */,
  {32'hbf762ecc, 32'hbe5ae55a} /* (21, 24, 16) {real, imag} */,
  {32'hbf7304f4, 32'hbe23f730} /* (21, 24, 15) {real, imag} */,
  {32'h3f8a83ae, 32'hbd55c8c0} /* (21, 24, 14) {real, imag} */,
  {32'h401189fa, 32'hbd4d3d00} /* (21, 24, 13) {real, imag} */,
  {32'h3f59fbc4, 32'hbedfbb34} /* (21, 24, 12) {real, imag} */,
  {32'hbeee1d70, 32'hbfbaafac} /* (21, 24, 11) {real, imag} */,
  {32'h3fd8014c, 32'hbec1ca27} /* (21, 24, 10) {real, imag} */,
  {32'h3fd0bcad, 32'h3e982ca8} /* (21, 24, 9) {real, imag} */,
  {32'h3f2dcc4e, 32'h3f1c3590} /* (21, 24, 8) {real, imag} */,
  {32'h3dd78430, 32'h3e877564} /* (21, 24, 7) {real, imag} */,
  {32'h3e6983e0, 32'h3f8c7cdb} /* (21, 24, 6) {real, imag} */,
  {32'h3f9c7e87, 32'h3db3c388} /* (21, 24, 5) {real, imag} */,
  {32'h3f3532d2, 32'hbf3c5b6c} /* (21, 24, 4) {real, imag} */,
  {32'h3e3ec69e, 32'h3e4c5560} /* (21, 24, 3) {real, imag} */,
  {32'h3f82b2a4, 32'h3fd0d5b0} /* (21, 24, 2) {real, imag} */,
  {32'h3fe53c14, 32'h3ecc4d20} /* (21, 24, 1) {real, imag} */,
  {32'h3ed787c1, 32'h3f5397b0} /* (21, 24, 0) {real, imag} */,
  {32'h3faceb92, 32'h3dd6e47c} /* (21, 23, 31) {real, imag} */,
  {32'h3f96fbd0, 32'hbe2d1998} /* (21, 23, 30) {real, imag} */,
  {32'h3f6210ea, 32'h3f86b4e5} /* (21, 23, 29) {real, imag} */,
  {32'hbf50b56c, 32'h3f14fa88} /* (21, 23, 28) {real, imag} */,
  {32'hbe8b0030, 32'h3f2564c4} /* (21, 23, 27) {real, imag} */,
  {32'h3eaa2f50, 32'h3b76e600} /* (21, 23, 26) {real, imag} */,
  {32'h3f71a21c, 32'h3f5e0862} /* (21, 23, 25) {real, imag} */,
  {32'h3fda666c, 32'h3df7a4e0} /* (21, 23, 24) {real, imag} */,
  {32'h40577841, 32'h3fc74540} /* (21, 23, 23) {real, imag} */,
  {32'h3fcead30, 32'h3fca1793} /* (21, 23, 22) {real, imag} */,
  {32'hbe2f6c49, 32'h3f056cb5} /* (21, 23, 21) {real, imag} */,
  {32'hbf432e30, 32'h3ea58eef} /* (21, 23, 20) {real, imag} */,
  {32'hbfadaba9, 32'hbea814c4} /* (21, 23, 19) {real, imag} */,
  {32'hc02a972e, 32'hbe1579b8} /* (21, 23, 18) {real, imag} */,
  {32'hbffd8d35, 32'hbe3de3c0} /* (21, 23, 17) {real, imag} */,
  {32'hbfa5e570, 32'h3eb528f4} /* (21, 23, 16) {real, imag} */,
  {32'hbe2a3dac, 32'hbe9e9f68} /* (21, 23, 15) {real, imag} */,
  {32'h3eecef58, 32'hbf119960} /* (21, 23, 14) {real, imag} */,
  {32'h3fd6c2fc, 32'hbe9f30dc} /* (21, 23, 13) {real, imag} */,
  {32'h3f5171d6, 32'hbe29b8c8} /* (21, 23, 12) {real, imag} */,
  {32'h3e405b54, 32'hbf206f68} /* (21, 23, 11) {real, imag} */,
  {32'h3fbd29d4, 32'hbe15dee8} /* (21, 23, 10) {real, imag} */,
  {32'h3f52745b, 32'h3c59fd80} /* (21, 23, 9) {real, imag} */,
  {32'h3f79acfe, 32'h3f0fe7d8} /* (21, 23, 8) {real, imag} */,
  {32'hbd03d110, 32'h3f16067c} /* (21, 23, 7) {real, imag} */,
  {32'h3e282d78, 32'h3fd0bcc7} /* (21, 23, 6) {real, imag} */,
  {32'h3f9a61f8, 32'h3fa05566} /* (21, 23, 5) {real, imag} */,
  {32'h3e133410, 32'h3f8a9c5d} /* (21, 23, 4) {real, imag} */,
  {32'hbf6b79f8, 32'h3eaafdce} /* (21, 23, 3) {real, imag} */,
  {32'h3def7f78, 32'h3f36e522} /* (21, 23, 2) {real, imag} */,
  {32'h3fcb5515, 32'h3e0567d4} /* (21, 23, 1) {real, imag} */,
  {32'h3ec325a4, 32'h3f178316} /* (21, 23, 0) {real, imag} */,
  {32'h3fcce4fc, 32'h3ea65964} /* (21, 22, 31) {real, imag} */,
  {32'h3fb3b8eb, 32'h3db27870} /* (21, 22, 30) {real, imag} */,
  {32'h3fb99459, 32'hbe433a50} /* (21, 22, 29) {real, imag} */,
  {32'h3f47dd66, 32'h3e23ab40} /* (21, 22, 28) {real, imag} */,
  {32'h3e03a4f0, 32'hbe3f2cb8} /* (21, 22, 27) {real, imag} */,
  {32'h3f587cb8, 32'h3dcf7f90} /* (21, 22, 26) {real, imag} */,
  {32'h3fd9bfa0, 32'h3fa7e778} /* (21, 22, 25) {real, imag} */,
  {32'h3ffba29d, 32'h3eaa0d8c} /* (21, 22, 24) {real, imag} */,
  {32'h40496b06, 32'hbe89d508} /* (21, 22, 23) {real, imag} */,
  {32'h3fe626fc, 32'h3eb668d8} /* (21, 22, 22) {real, imag} */,
  {32'h3f6100fe, 32'h3ed2ceb1} /* (21, 22, 21) {real, imag} */,
  {32'hbfc820eb, 32'h3e02863e} /* (21, 22, 20) {real, imag} */,
  {32'hbefbcc00, 32'hbea8287c} /* (21, 22, 19) {real, imag} */,
  {32'hbf91b451, 32'hbf9c3dd4} /* (21, 22, 18) {real, imag} */,
  {32'hbfc6cdf2, 32'hbf4b0ee4} /* (21, 22, 17) {real, imag} */,
  {32'hbf559ef5, 32'hbd4d3110} /* (21, 22, 16) {real, imag} */,
  {32'hbeafd4db, 32'hbeb6f1de} /* (21, 22, 15) {real, imag} */,
  {32'hbd9d9170, 32'hbf30615e} /* (21, 22, 14) {real, imag} */,
  {32'h3e4e3b06, 32'hbf9d2450} /* (21, 22, 13) {real, imag} */,
  {32'h3e1112b0, 32'hbfdab089} /* (21, 22, 12) {real, imag} */,
  {32'hbdfc4c90, 32'hbfbe3186} /* (21, 22, 11) {real, imag} */,
  {32'h3fdf5e94, 32'hbe000220} /* (21, 22, 10) {real, imag} */,
  {32'h400297f8, 32'h3f6a45c0} /* (21, 22, 9) {real, imag} */,
  {32'h400dadfc, 32'h3f30bf58} /* (21, 22, 8) {real, imag} */,
  {32'h3f86a564, 32'h3f6d24a4} /* (21, 22, 7) {real, imag} */,
  {32'h3fdcdc31, 32'h3f982c68} /* (21, 22, 6) {real, imag} */,
  {32'h3f6a74ac, 32'h3f881b12} /* (21, 22, 5) {real, imag} */,
  {32'hbe7fda14, 32'h3f75398b} /* (21, 22, 4) {real, imag} */,
  {32'h3ea17e86, 32'h3f3c8fc1} /* (21, 22, 3) {real, imag} */,
  {32'h3f7dee7a, 32'h3f7384be} /* (21, 22, 2) {real, imag} */,
  {32'h40114c2a, 32'hbf4e87c2} /* (21, 22, 1) {real, imag} */,
  {32'h3f9a4f77, 32'h3cc41c40} /* (21, 22, 0) {real, imag} */,
  {32'h3f87a975, 32'h3eaffae1} /* (21, 21, 31) {real, imag} */,
  {32'h3f1cdc3c, 32'h3f2638f2} /* (21, 21, 30) {real, imag} */,
  {32'h3ee8a174, 32'hbefcb194} /* (21, 21, 29) {real, imag} */,
  {32'h3de38ff8, 32'hbce070e0} /* (21, 21, 28) {real, imag} */,
  {32'hbe247b88, 32'h3fda1dd5} /* (21, 21, 27) {real, imag} */,
  {32'h3fa02c6d, 32'h3fb37248} /* (21, 21, 26) {real, imag} */,
  {32'h4002c543, 32'h3f650d20} /* (21, 21, 25) {real, imag} */,
  {32'h3f8d6338, 32'hbdc6cb00} /* (21, 21, 24) {real, imag} */,
  {32'h3e1f1f16, 32'hbdb6bb00} /* (21, 21, 23) {real, imag} */,
  {32'h3e9b892c, 32'h3e6af7d0} /* (21, 21, 22) {real, imag} */,
  {32'h3f09145a, 32'hbebb2c14} /* (21, 21, 21) {real, imag} */,
  {32'hbfec933a, 32'hbfcc17bd} /* (21, 21, 20) {real, imag} */,
  {32'hbf771f16, 32'hbe4af56c} /* (21, 21, 19) {real, imag} */,
  {32'h3f864db0, 32'h3c0c4480} /* (21, 21, 18) {real, imag} */,
  {32'h3dd67f78, 32'hbf35fec7} /* (21, 21, 17) {real, imag} */,
  {32'hbea5794a, 32'hbf031de4} /* (21, 21, 16) {real, imag} */,
  {32'hbfa2c641, 32'hbf290b54} /* (21, 21, 15) {real, imag} */,
  {32'hbee44bf6, 32'hbea13b1c} /* (21, 21, 14) {real, imag} */,
  {32'hbf01a914, 32'hbf2ba7e2} /* (21, 21, 13) {real, imag} */,
  {32'hbe8fb300, 32'hbfef6acc} /* (21, 21, 12) {real, imag} */,
  {32'h3c422c00, 32'hbfc7560e} /* (21, 21, 11) {real, imag} */,
  {32'h3f92a70f, 32'h3f11c620} /* (21, 21, 10) {real, imag} */,
  {32'h3f92bdeb, 32'h3ffdfb8b} /* (21, 21, 9) {real, imag} */,
  {32'h4009f972, 32'h3fc1ca5a} /* (21, 21, 8) {real, imag} */,
  {32'h4027874a, 32'h3fb63e4c} /* (21, 21, 7) {real, imag} */,
  {32'h40260421, 32'h3e33d2e4} /* (21, 21, 6) {real, imag} */,
  {32'h3f579d6c, 32'hbe221064} /* (21, 21, 5) {real, imag} */,
  {32'hbf225a50, 32'h3de0bf2a} /* (21, 21, 4) {real, imag} */,
  {32'h3eab3164, 32'hbeaeb784} /* (21, 21, 3) {real, imag} */,
  {32'h3f6acf72, 32'h3fc2d853} /* (21, 21, 2) {real, imag} */,
  {32'h3f2aeb52, 32'hbe1eec0c} /* (21, 21, 1) {real, imag} */,
  {32'h3e0f08ba, 32'h3e6a23bc} /* (21, 21, 0) {real, imag} */,
  {32'hbe3d2fa0, 32'hbe68a498} /* (21, 20, 31) {real, imag} */,
  {32'hbeccb75c, 32'hbef9f412} /* (21, 20, 30) {real, imag} */,
  {32'hbf8d4813, 32'hbeff7d5c} /* (21, 20, 29) {real, imag} */,
  {32'hbfd4f8f6, 32'hbf7e41f2} /* (21, 20, 28) {real, imag} */,
  {32'hbf9bb97f, 32'h3e7d5388} /* (21, 20, 27) {real, imag} */,
  {32'h3e633c54, 32'h3f7ff91d} /* (21, 20, 26) {real, imag} */,
  {32'h3f2e7214, 32'h3eb697dc} /* (21, 20, 25) {real, imag} */,
  {32'h3e652620, 32'hbf151a8c} /* (21, 20, 24) {real, imag} */,
  {32'hbeb34504, 32'hbf295c14} /* (21, 20, 23) {real, imag} */,
  {32'hbeb4bd10, 32'hbf90c010} /* (21, 20, 22) {real, imag} */,
  {32'h3df3cc84, 32'hbfa82d5b} /* (21, 20, 21) {real, imag} */,
  {32'hbec00b28, 32'hbf935d4a} /* (21, 20, 20) {real, imag} */,
  {32'hbf02c086, 32'hbe792f84} /* (21, 20, 19) {real, imag} */,
  {32'h3f49d97e, 32'hbf025e36} /* (21, 20, 18) {real, imag} */,
  {32'h3f89fbd8, 32'hbf255695} /* (21, 20, 17) {real, imag} */,
  {32'h3f8c2ed4, 32'hbe854c58} /* (21, 20, 16) {real, imag} */,
  {32'h3d863370, 32'hbedbbef1} /* (21, 20, 15) {real, imag} */,
  {32'hbf07bd2a, 32'h3f1e693f} /* (21, 20, 14) {real, imag} */,
  {32'h3e97ad82, 32'hbdf868b0} /* (21, 20, 13) {real, imag} */,
  {32'h3f7e3011, 32'hbe839078} /* (21, 20, 12) {real, imag} */,
  {32'h3e03a6d0, 32'hbf9392df} /* (21, 20, 11) {real, imag} */,
  {32'hbf9ab332, 32'hbf44c651} /* (21, 20, 10) {real, imag} */,
  {32'hbf7d448e, 32'h3dec78e0} /* (21, 20, 9) {real, imag} */,
  {32'h3fc2077c, 32'h3f8a5c74} /* (21, 20, 8) {real, imag} */,
  {32'h3fdc42e7, 32'h3f09e57a} /* (21, 20, 7) {real, imag} */,
  {32'h3eca8a57, 32'hbfbe8e4a} /* (21, 20, 6) {real, imag} */,
  {32'hbefe5790, 32'hbf2ea9dc} /* (21, 20, 5) {real, imag} */,
  {32'hbf2be5b4, 32'h3ef929ea} /* (21, 20, 4) {real, imag} */,
  {32'hbf81f476, 32'hbe410d00} /* (21, 20, 3) {real, imag} */,
  {32'hbf520ee7, 32'h3fca6e4e} /* (21, 20, 2) {real, imag} */,
  {32'hbf25a020, 32'hbebdf39c} /* (21, 20, 1) {real, imag} */,
  {32'hbea53689, 32'hbf007b18} /* (21, 20, 0) {real, imag} */,
  {32'hbe98f63c, 32'hbed34a0a} /* (21, 19, 31) {real, imag} */,
  {32'h3f2ddc9a, 32'hbea70f42} /* (21, 19, 30) {real, imag} */,
  {32'h3da28068, 32'hbd36f894} /* (21, 19, 29) {real, imag} */,
  {32'hbf6eeb01, 32'hbfa17bc6} /* (21, 19, 28) {real, imag} */,
  {32'hbfdd8c2e, 32'hbfac05de} /* (21, 19, 27) {real, imag} */,
  {32'hbf3fb6af, 32'h3f26df76} /* (21, 19, 26) {real, imag} */,
  {32'h3e7b4180, 32'h3f2ed360} /* (21, 19, 25) {real, imag} */,
  {32'h3e7d42d0, 32'hbf7e5b4c} /* (21, 19, 24) {real, imag} */,
  {32'hbdde0000, 32'hbffb7dd3} /* (21, 19, 23) {real, imag} */,
  {32'hbfc76b1e, 32'hbfd55635} /* (21, 19, 22) {real, imag} */,
  {32'hbe2f4171, 32'hbf6d20be} /* (21, 19, 21) {real, imag} */,
  {32'h3fa9dcc6, 32'hbfa55872} /* (21, 19, 20) {real, imag} */,
  {32'h3f5e6c93, 32'hbf16b110} /* (21, 19, 19) {real, imag} */,
  {32'hbde6b380, 32'h3eb9ed74} /* (21, 19, 18) {real, imag} */,
  {32'h3e15a990, 32'hbc22ba80} /* (21, 19, 17) {real, imag} */,
  {32'h3fcf9ab5, 32'h3f3b2bfe} /* (21, 19, 16) {real, imag} */,
  {32'h3f4b3c7e, 32'h3f5ae05f} /* (21, 19, 15) {real, imag} */,
  {32'hbd5f4e40, 32'h3fadf1dd} /* (21, 19, 14) {real, imag} */,
  {32'h3f69a2ae, 32'hbddf1830} /* (21, 19, 13) {real, imag} */,
  {32'h3f96861a, 32'h3d0f5d70} /* (21, 19, 12) {real, imag} */,
  {32'hbf048e9f, 32'h3cf22d00} /* (21, 19, 11) {real, imag} */,
  {32'hbff1e4a0, 32'hbf3ca662} /* (21, 19, 10) {real, imag} */,
  {32'hbf721c4b, 32'hbda27cb0} /* (21, 19, 9) {real, imag} */,
  {32'h3f948024, 32'h3f349fec} /* (21, 19, 8) {real, imag} */,
  {32'h3dcb03a8, 32'h3f414a98} /* (21, 19, 7) {real, imag} */,
  {32'hbeff4a78, 32'h3dc69330} /* (21, 19, 6) {real, imag} */,
  {32'hbf139da8, 32'hbefc6b3c} /* (21, 19, 5) {real, imag} */,
  {32'hbf9cf210, 32'hbe9c3104} /* (21, 19, 4) {real, imag} */,
  {32'hbf536c88, 32'h3f7e425a} /* (21, 19, 3) {real, imag} */,
  {32'h3d824e58, 32'h3ef5fc54} /* (21, 19, 2) {real, imag} */,
  {32'h3e296cbc, 32'hbf4d2fc5} /* (21, 19, 1) {real, imag} */,
  {32'hbe34658e, 32'hbe773000} /* (21, 19, 0) {real, imag} */,
  {32'hbf856abc, 32'h3ed2c5e4} /* (21, 18, 31) {real, imag} */,
  {32'h3f2f4212, 32'h3d7c9f20} /* (21, 18, 30) {real, imag} */,
  {32'h3f96073e, 32'hbf5a6c24} /* (21, 18, 29) {real, imag} */,
  {32'hbe281a50, 32'hbfa578d1} /* (21, 18, 28) {real, imag} */,
  {32'hbfc5ae56, 32'hbf60f0d3} /* (21, 18, 27) {real, imag} */,
  {32'hbf9ce98d, 32'h3eb481f6} /* (21, 18, 26) {real, imag} */,
  {32'hbf96a18c, 32'h3f2a339a} /* (21, 18, 25) {real, imag} */,
  {32'hbf0842bc, 32'hbef18428} /* (21, 18, 24) {real, imag} */,
  {32'hbefa8e44, 32'h3ef6db44} /* (21, 18, 23) {real, imag} */,
  {32'hbee340f4, 32'h3f0d01c6} /* (21, 18, 22) {real, imag} */,
  {32'h3ed16321, 32'hbec62ca2} /* (21, 18, 21) {real, imag} */,
  {32'h3f4a77bc, 32'hbf88f8fa} /* (21, 18, 20) {real, imag} */,
  {32'h3f7b6948, 32'hbe637398} /* (21, 18, 19) {real, imag} */,
  {32'h3f72f084, 32'h3fb7960b} /* (21, 18, 18) {real, imag} */,
  {32'h3f62bf52, 32'h3ff40bed} /* (21, 18, 17) {real, imag} */,
  {32'h3ff08a62, 32'h3fdf19be} /* (21, 18, 16) {real, imag} */,
  {32'h3f88e78f, 32'h3edf5f04} /* (21, 18, 15) {real, imag} */,
  {32'hbe3ca1c8, 32'h3f4df9d2} /* (21, 18, 14) {real, imag} */,
  {32'hbe6a7300, 32'h3ec1d110} /* (21, 18, 13) {real, imag} */,
  {32'hbf749346, 32'h3f88a311} /* (21, 18, 12) {real, imag} */,
  {32'hbfbf05e2, 32'h4008358a} /* (21, 18, 11) {real, imag} */,
  {32'hbf9fae80, 32'hbeeba364} /* (21, 18, 10) {real, imag} */,
  {32'hbfa92baa, 32'hbffc7b46} /* (21, 18, 9) {real, imag} */,
  {32'h3f9c0c71, 32'hbfc6d94b} /* (21, 18, 8) {real, imag} */,
  {32'h3ed97740, 32'hbf0e7028} /* (21, 18, 7) {real, imag} */,
  {32'h3e5f4510, 32'hbf0ae552} /* (21, 18, 6) {real, imag} */,
  {32'h3f49259c, 32'hbf68c160} /* (21, 18, 5) {real, imag} */,
  {32'hbec1ac70, 32'hbf6b64c8} /* (21, 18, 4) {real, imag} */,
  {32'hbda42be4, 32'hbdda7600} /* (21, 18, 3) {real, imag} */,
  {32'h3e3d6b88, 32'hbe8171c5} /* (21, 18, 2) {real, imag} */,
  {32'h3ee56060, 32'h3dd423c0} /* (21, 18, 1) {real, imag} */,
  {32'hbf4d54d9, 32'h3eb44cea} /* (21, 18, 0) {real, imag} */,
  {32'hbf0d3cfc, 32'hbb662e00} /* (21, 17, 31) {real, imag} */,
  {32'hbda74fa0, 32'hbe3fc0c0} /* (21, 17, 30) {real, imag} */,
  {32'h3e95e070, 32'hbf942c86} /* (21, 17, 29) {real, imag} */,
  {32'hbf964bb6, 32'hbf37f33c} /* (21, 17, 28) {real, imag} */,
  {32'hbfc5f6c6, 32'h3eb6e7f6} /* (21, 17, 27) {real, imag} */,
  {32'hbf3db134, 32'h3e428d44} /* (21, 17, 26) {real, imag} */,
  {32'hbfb10616, 32'hbf514990} /* (21, 17, 25) {real, imag} */,
  {32'hbf7a8e4a, 32'hbfbc9b65} /* (21, 17, 24) {real, imag} */,
  {32'hbf918d48, 32'h3f89c57a} /* (21, 17, 23) {real, imag} */,
  {32'hbf825daa, 32'hbd363180} /* (21, 17, 22) {real, imag} */,
  {32'hbf6ec854, 32'hbf0ea081} /* (21, 17, 21) {real, imag} */,
  {32'hbea57d38, 32'hbf693a45} /* (21, 17, 20) {real, imag} */,
  {32'h3f39448e, 32'hbd9ded00} /* (21, 17, 19) {real, imag} */,
  {32'h3f70e8b0, 32'h3fb9e099} /* (21, 17, 18) {real, imag} */,
  {32'h3fddddec, 32'h4027eba7} /* (21, 17, 17) {real, imag} */,
  {32'h3ff96320, 32'h3fcaad4d} /* (21, 17, 16) {real, imag} */,
  {32'h3f7d6c94, 32'h3f01f028} /* (21, 17, 15) {real, imag} */,
  {32'h3deaa4a0, 32'hbc854f00} /* (21, 17, 14) {real, imag} */,
  {32'h3e89fb38, 32'h3ec826c2} /* (21, 17, 13) {real, imag} */,
  {32'hbe68d928, 32'h3f88afea} /* (21, 17, 12) {real, imag} */,
  {32'hbfb91304, 32'h3fcd681e} /* (21, 17, 11) {real, imag} */,
  {32'hbf8e3142, 32'hbf8df2bc} /* (21, 17, 10) {real, imag} */,
  {32'hbf20365c, 32'hc02c1fd8} /* (21, 17, 9) {real, imag} */,
  {32'hbeece6d8, 32'hc0212367} /* (21, 17, 8) {real, imag} */,
  {32'hbf311fc6, 32'hbfd5ec2e} /* (21, 17, 7) {real, imag} */,
  {32'hbed77a6c, 32'hbf8b1134} /* (21, 17, 6) {real, imag} */,
  {32'hbede22c0, 32'h3de123a0} /* (21, 17, 5) {real, imag} */,
  {32'hbf22c7fe, 32'h3e10afd8} /* (21, 17, 4) {real, imag} */,
  {32'hbee84ffe, 32'h3f041b60} /* (21, 17, 3) {real, imag} */,
  {32'hbd8fcd8c, 32'h3e0b9d28} /* (21, 17, 2) {real, imag} */,
  {32'h3f4ad2b0, 32'h3f8406d3} /* (21, 17, 1) {real, imag} */,
  {32'hbe92991f, 32'h3f0441ac} /* (21, 17, 0) {real, imag} */,
  {32'hbf0d6fe9, 32'hbf1898ac} /* (21, 16, 31) {real, imag} */,
  {32'h3e1d7a68, 32'h3e548450} /* (21, 16, 30) {real, imag} */,
  {32'h3ed1f346, 32'hbef21ad8} /* (21, 16, 29) {real, imag} */,
  {32'hbf64c1bc, 32'hbf60e366} /* (21, 16, 28) {real, imag} */,
  {32'hbf8d153d, 32'hbeaef7cc} /* (21, 16, 27) {real, imag} */,
  {32'hbf3cb7c1, 32'hbf9389a6} /* (21, 16, 26) {real, imag} */,
  {32'hbf3efc54, 32'hc02e4d47} /* (21, 16, 25) {real, imag} */,
  {32'hbf02d75a, 32'hc0141596} /* (21, 16, 24) {real, imag} */,
  {32'hbf784cbe, 32'hbee8c208} /* (21, 16, 23) {real, imag} */,
  {32'hbfcbc7f0, 32'hbf31c594} /* (21, 16, 22) {real, imag} */,
  {32'hbfa610a2, 32'h3f6af25f} /* (21, 16, 21) {real, imag} */,
  {32'h3dfd0260, 32'hbebe5210} /* (21, 16, 20) {real, imag} */,
  {32'h3f98f3a8, 32'h3ee62812} /* (21, 16, 19) {real, imag} */,
  {32'h3f98b995, 32'h3fb9ad9d} /* (21, 16, 18) {real, imag} */,
  {32'hbd7df000, 32'h3fc1a1d6} /* (21, 16, 17) {real, imag} */,
  {32'h3f62e052, 32'h3f73a18c} /* (21, 16, 16) {real, imag} */,
  {32'h3f8e7631, 32'hbe2400a8} /* (21, 16, 15) {real, imag} */,
  {32'h3f207e92, 32'hbfa9ad4a} /* (21, 16, 14) {real, imag} */,
  {32'hbf510c45, 32'hbebd20d6} /* (21, 16, 13) {real, imag} */,
  {32'hbef3d4c0, 32'h3d85a410} /* (21, 16, 12) {real, imag} */,
  {32'hbe1d2248, 32'h3e2cfba8} /* (21, 16, 11) {real, imag} */,
  {32'h3d1dbf00, 32'hbf8f5342} /* (21, 16, 10) {real, imag} */,
  {32'h3f7d788f, 32'hbf65ba8a} /* (21, 16, 9) {real, imag} */,
  {32'hbfa14451, 32'hbdb11420} /* (21, 16, 8) {real, imag} */,
  {32'hc01e778b, 32'hbf2c0ac4} /* (21, 16, 7) {real, imag} */,
  {32'hbfa5b085, 32'hbfd39097} /* (21, 16, 6) {real, imag} */,
  {32'hbeee9fc0, 32'hbd7d8b60} /* (21, 16, 5) {real, imag} */,
  {32'hbf92e0f4, 32'h3ec34e50} /* (21, 16, 4) {real, imag} */,
  {32'hbffb7b56, 32'h3e34c3f0} /* (21, 16, 3) {real, imag} */,
  {32'hbea107b4, 32'h3ea8f010} /* (21, 16, 2) {real, imag} */,
  {32'h3ef3e7a0, 32'h3f6fcb1e} /* (21, 16, 1) {real, imag} */,
  {32'h3e0cff70, 32'h3d8bd618} /* (21, 16, 0) {real, imag} */,
  {32'h3c158880, 32'hbf177831} /* (21, 15, 31) {real, imag} */,
  {32'hbf46104e, 32'h3fa3ba6c} /* (21, 15, 30) {real, imag} */,
  {32'hbebe1d3c, 32'h3f1d7a14} /* (21, 15, 29) {real, imag} */,
  {32'hbfa15958, 32'hbfb65358} /* (21, 15, 28) {real, imag} */,
  {32'hbf5df988, 32'hbfbe860b} /* (21, 15, 27) {real, imag} */,
  {32'hbf1139fb, 32'hbf947115} /* (21, 15, 26) {real, imag} */,
  {32'hbfc18f78, 32'hbfb673f4} /* (21, 15, 25) {real, imag} */,
  {32'hbf838953, 32'hbf9c5d1e} /* (21, 15, 24) {real, imag} */,
  {32'hbf5f99f0, 32'h3ed87068} /* (21, 15, 23) {real, imag} */,
  {32'hbf9630ab, 32'hbe8cd9a8} /* (21, 15, 22) {real, imag} */,
  {32'hbead98c4, 32'h3dad42d0} /* (21, 15, 21) {real, imag} */,
  {32'h3f1c0a89, 32'hbe062958} /* (21, 15, 20) {real, imag} */,
  {32'h3f78ce7c, 32'h3f9b9bf2} /* (21, 15, 19) {real, imag} */,
  {32'h3c5ac7d0, 32'h3ff5f50a} /* (21, 15, 18) {real, imag} */,
  {32'hbf37e48e, 32'h3fd24357} /* (21, 15, 17) {real, imag} */,
  {32'h3f9c13dc, 32'h3f219e0e} /* (21, 15, 16) {real, imag} */,
  {32'h3fb7a58d, 32'hbf1a911a} /* (21, 15, 15) {real, imag} */,
  {32'h3fc9dca6, 32'hbfa0507b} /* (21, 15, 14) {real, imag} */,
  {32'hbee42f16, 32'hbe787f30} /* (21, 15, 13) {real, imag} */,
  {32'hbfd88eac, 32'hbe5bbf20} /* (21, 15, 12) {real, imag} */,
  {32'hbf0be7f4, 32'hbe8b6670} /* (21, 15, 11) {real, imag} */,
  {32'hbf33727c, 32'hbf62f3d8} /* (21, 15, 10) {real, imag} */,
  {32'hbe5ad368, 32'hbfe39af7} /* (21, 15, 9) {real, imag} */,
  {32'hbfea583c, 32'hbf024444} /* (21, 15, 8) {real, imag} */,
  {32'hc0323e1e, 32'h3f3552f4} /* (21, 15, 7) {real, imag} */,
  {32'hbf83e326, 32'hbdeb1360} /* (21, 15, 6) {real, imag} */,
  {32'h3ec0c8fe, 32'hbeb31a56} /* (21, 15, 5) {real, imag} */,
  {32'h3e602a0c, 32'hbdad7dc4} /* (21, 15, 4) {real, imag} */,
  {32'hbf066974, 32'hbe6756a0} /* (21, 15, 3) {real, imag} */,
  {32'h3d219cc0, 32'h3d161900} /* (21, 15, 2) {real, imag} */,
  {32'h3f4ddd04, 32'h3f44922a} /* (21, 15, 1) {real, imag} */,
  {32'h3ec1635c, 32'h3e8fb5f4} /* (21, 15, 0) {real, imag} */,
  {32'hbfb1886b, 32'hbdf80438} /* (21, 14, 31) {real, imag} */,
  {32'hc0380748, 32'h3f218ab8} /* (21, 14, 30) {real, imag} */,
  {32'hc01193fe, 32'hbe05b7f8} /* (21, 14, 29) {real, imag} */,
  {32'hbfe6d475, 32'hbfd57cf0} /* (21, 14, 28) {real, imag} */,
  {32'hc011826c, 32'hbf990d8d} /* (21, 14, 27) {real, imag} */,
  {32'hc013834e, 32'hbe6f87d8} /* (21, 14, 26) {real, imag} */,
  {32'hc02547f4, 32'hbf72ca48} /* (21, 14, 25) {real, imag} */,
  {32'hbfd6f038, 32'hbfa68e3c} /* (21, 14, 24) {real, imag} */,
  {32'hbfcd1bd4, 32'hbef2f0c8} /* (21, 14, 23) {real, imag} */,
  {32'hc00bc0aa, 32'h3f31e754} /* (21, 14, 22) {real, imag} */,
  {32'hbf291a0e, 32'h3f441b05} /* (21, 14, 21) {real, imag} */,
  {32'h3faac95c, 32'h3f459824} /* (21, 14, 20) {real, imag} */,
  {32'h3eda13c4, 32'h3f48998d} /* (21, 14, 19) {real, imag} */,
  {32'hbd557220, 32'h3f318294} /* (21, 14, 18) {real, imag} */,
  {32'h3f2551e9, 32'h3dbd2270} /* (21, 14, 17) {real, imag} */,
  {32'h3faf45c2, 32'h3f178480} /* (21, 14, 16) {real, imag} */,
  {32'h3fd5590c, 32'hbd191ef0} /* (21, 14, 15) {real, imag} */,
  {32'h4012e6cc, 32'h3e34aca0} /* (21, 14, 14) {real, imag} */,
  {32'h3fda6de5, 32'h3e3d78e8} /* (21, 14, 13) {real, imag} */,
  {32'h3f233a4c, 32'hbef4407c} /* (21, 14, 12) {real, imag} */,
  {32'h3f751832, 32'hbf2dc0a8} /* (21, 14, 11) {real, imag} */,
  {32'hbf895d4c, 32'hbfcc6c8c} /* (21, 14, 10) {real, imag} */,
  {32'hbf4158e8, 32'hc00a81ec} /* (21, 14, 9) {real, imag} */,
  {32'hbe5af508, 32'hbf6f336c} /* (21, 14, 8) {real, imag} */,
  {32'hbfd5ba59, 32'hbf3a5b52} /* (21, 14, 7) {real, imag} */,
  {32'hbfaa876c, 32'hbbfc8980} /* (21, 14, 6) {real, imag} */,
  {32'h3e72f188, 32'h3f24f264} /* (21, 14, 5) {real, imag} */,
  {32'h3f777d5d, 32'h3d823008} /* (21, 14, 4) {real, imag} */,
  {32'h3e36c180, 32'h3de96a80} /* (21, 14, 3) {real, imag} */,
  {32'hbdded1b0, 32'h3f6eebdf} /* (21, 14, 2) {real, imag} */,
  {32'h3faa8ec1, 32'h3f9261b0} /* (21, 14, 1) {real, imag} */,
  {32'h3f1f631c, 32'h3f0a168b} /* (21, 14, 0) {real, imag} */,
  {32'hbfb86ee9, 32'hbf0f93ca} /* (21, 13, 31) {real, imag} */,
  {32'hc038ad5a, 32'hbf29ca1d} /* (21, 13, 30) {real, imag} */,
  {32'hc0115d06, 32'hbff9d01a} /* (21, 13, 29) {real, imag} */,
  {32'hc0156a74, 32'hc00549b8} /* (21, 13, 28) {real, imag} */,
  {32'hbfeeafca, 32'hbf211466} /* (21, 13, 27) {real, imag} */,
  {32'hbfdc6ceb, 32'h3e801f68} /* (21, 13, 26) {real, imag} */,
  {32'hc021db20, 32'hbf712a18} /* (21, 13, 25) {real, imag} */,
  {32'hc006ae8e, 32'hbfeb63b8} /* (21, 13, 24) {real, imag} */,
  {32'hbfa44994, 32'hc00bc588} /* (21, 13, 23) {real, imag} */,
  {32'hc004219e, 32'hbfa8ca05} /* (21, 13, 22) {real, imag} */,
  {32'hbff47825, 32'hbf4c7755} /* (21, 13, 21) {real, imag} */,
  {32'h3fcd35b9, 32'hbf2807e4} /* (21, 13, 20) {real, imag} */,
  {32'h3fb73bf3, 32'hbfa260e0} /* (21, 13, 19) {real, imag} */,
  {32'h3fe3c7d5, 32'hbf0d0790} /* (21, 13, 18) {real, imag} */,
  {32'h3fccfd1e, 32'hbec1bf20} /* (21, 13, 17) {real, imag} */,
  {32'h3fa90e94, 32'hbc8784f0} /* (21, 13, 16) {real, imag} */,
  {32'h3efc97b4, 32'hbe63385c} /* (21, 13, 15) {real, imag} */,
  {32'h3f694f62, 32'h3f2d4b8e} /* (21, 13, 14) {real, imag} */,
  {32'h3fea5e68, 32'h3e8e0e48} /* (21, 13, 13) {real, imag} */,
  {32'h3fd2fea1, 32'hbf236023} /* (21, 13, 12) {real, imag} */,
  {32'h3f79e9dd, 32'hbf6c7158} /* (21, 13, 11) {real, imag} */,
  {32'hc00685ee, 32'hbfe76258} /* (21, 13, 10) {real, imag} */,
  {32'hbf0b2a1a, 32'hc0131e60} /* (21, 13, 9) {real, imag} */,
  {32'hbc253e00, 32'hbf23647d} /* (21, 13, 8) {real, imag} */,
  {32'hbf990f62, 32'hbfc752a0} /* (21, 13, 7) {real, imag} */,
  {32'hbf8b3d00, 32'hbf347b1f} /* (21, 13, 6) {real, imag} */,
  {32'hbd50b5f8, 32'h3e06fb40} /* (21, 13, 5) {real, imag} */,
  {32'hbe155564, 32'hbf8fa79f} /* (21, 13, 4) {real, imag} */,
  {32'hbfa0a71a, 32'hbea300b0} /* (21, 13, 3) {real, imag} */,
  {32'hbf9ba868, 32'h3fa6f1be} /* (21, 13, 2) {real, imag} */,
  {32'h3f6caf40, 32'h3fd45193} /* (21, 13, 1) {real, imag} */,
  {32'h3e8ab4a7, 32'h3e908e80} /* (21, 13, 0) {real, imag} */,
  {32'hbde5bbac, 32'hbfd88ec4} /* (21, 12, 31) {real, imag} */,
  {32'hbeb6883a, 32'hbfc5ca9a} /* (21, 12, 30) {real, imag} */,
  {32'hbeefc2d0, 32'hbfed7ade} /* (21, 12, 29) {real, imag} */,
  {32'hbf98aba6, 32'hbf9925b1} /* (21, 12, 28) {real, imag} */,
  {32'hbfeb10c7, 32'h3e2435f8} /* (21, 12, 27) {real, imag} */,
  {32'hbf05f9a2, 32'h3ec806a0} /* (21, 12, 26) {real, imag} */,
  {32'hbf95b6d0, 32'hbfe6acbd} /* (21, 12, 25) {real, imag} */,
  {32'hbff6ff1a, 32'hbeeeba4e} /* (21, 12, 24) {real, imag} */,
  {32'hbff6b3d5, 32'hbeb30988} /* (21, 12, 23) {real, imag} */,
  {32'hbf72f062, 32'hbf5c0230} /* (21, 12, 22) {real, imag} */,
  {32'hbfbaa88e, 32'hbf3f4c28} /* (21, 12, 21) {real, imag} */,
  {32'h3f5f3b68, 32'hbebee290} /* (21, 12, 20) {real, imag} */,
  {32'h401c42ec, 32'hbec55f10} /* (21, 12, 19) {real, imag} */,
  {32'h4025713e, 32'hbf418192} /* (21, 12, 18) {real, imag} */,
  {32'h40100a27, 32'hbf234bde} /* (21, 12, 17) {real, imag} */,
  {32'h3f465d78, 32'hbe1730b0} /* (21, 12, 16) {real, imag} */,
  {32'h3e47dd00, 32'hbe114488} /* (21, 12, 15) {real, imag} */,
  {32'h3f67603b, 32'h3edb81b6} /* (21, 12, 14) {real, imag} */,
  {32'h3f9bb39e, 32'h3ea2433a} /* (21, 12, 13) {real, imag} */,
  {32'h4003bbb8, 32'h3f186410} /* (21, 12, 12) {real, imag} */,
  {32'hbe3bb8e0, 32'h3e541998} /* (21, 12, 11) {real, imag} */,
  {32'hbfefb90c, 32'hbe479bc0} /* (21, 12, 10) {real, imag} */,
  {32'hbef5562c, 32'hbf9b2d6e} /* (21, 12, 9) {real, imag} */,
  {32'hbf311c82, 32'hbf53dd53} /* (21, 12, 8) {real, imag} */,
  {32'hbf001bf2, 32'hbf8918d5} /* (21, 12, 7) {real, imag} */,
  {32'hbf85b482, 32'hbf24ba66} /* (21, 12, 6) {real, imag} */,
  {32'hbf48a028, 32'hbed62622} /* (21, 12, 5) {real, imag} */,
  {32'hbeeffaf8, 32'hbf297765} /* (21, 12, 4) {real, imag} */,
  {32'hbf82b2de, 32'hbf7d8d5a} /* (21, 12, 3) {real, imag} */,
  {32'hc004ea22, 32'hbf155e4a} /* (21, 12, 2) {real, imag} */,
  {32'hbf3203b2, 32'h3f726f0c} /* (21, 12, 1) {real, imag} */,
  {32'h3e974e87, 32'hbd4f4230} /* (21, 12, 0) {real, imag} */,
  {32'h3ec52b9c, 32'hbe618014} /* (21, 11, 31) {real, imag} */,
  {32'h3ea41945, 32'hbe63ca98} /* (21, 11, 30) {real, imag} */,
  {32'h3e03a688, 32'hbf32db32} /* (21, 11, 29) {real, imag} */,
  {32'h3d67b940, 32'hbf7b9d8c} /* (21, 11, 28) {real, imag} */,
  {32'hbe6cbecc, 32'hbe72af94} /* (21, 11, 27) {real, imag} */,
  {32'hbeac55f4, 32'h3f2a7384} /* (21, 11, 26) {real, imag} */,
  {32'h3ec78a85, 32'hbf5cf492} /* (21, 11, 25) {real, imag} */,
  {32'hbf3bd5cc, 32'h3f8acf31} /* (21, 11, 24) {real, imag} */,
  {32'hc00786f4, 32'h3eda7928} /* (21, 11, 23) {real, imag} */,
  {32'hbf6c96de, 32'hbe727764} /* (21, 11, 22) {real, imag} */,
  {32'hbf23ef2c, 32'hbecc63e6} /* (21, 11, 21) {real, imag} */,
  {32'h3e82a7fc, 32'h3ed63aba} /* (21, 11, 20) {real, imag} */,
  {32'h3e6b21fc, 32'h3f669d8e} /* (21, 11, 19) {real, imag} */,
  {32'h3f655732, 32'h3f6c5654} /* (21, 11, 18) {real, imag} */,
  {32'h3f2e9ae6, 32'h3ebbfe90} /* (21, 11, 17) {real, imag} */,
  {32'hbedacf3b, 32'h3cbc5460} /* (21, 11, 16) {real, imag} */,
  {32'hbcae1520, 32'h3eaa81f8} /* (21, 11, 15) {real, imag} */,
  {32'h3f713ea8, 32'h3f8430f4} /* (21, 11, 14) {real, imag} */,
  {32'h3f93f519, 32'h3f8ef65c} /* (21, 11, 13) {real, imag} */,
  {32'h3f1ba632, 32'h3fa5cb5a} /* (21, 11, 12) {real, imag} */,
  {32'hbf6aff44, 32'h3f91cf73} /* (21, 11, 11) {real, imag} */,
  {32'hbf4aed3e, 32'h3cceede0} /* (21, 11, 10) {real, imag} */,
  {32'hbeab75d0, 32'hbff876e6} /* (21, 11, 9) {real, imag} */,
  {32'hbff54d2d, 32'hbfdb949e} /* (21, 11, 8) {real, imag} */,
  {32'hbfd025b7, 32'h3eb96640} /* (21, 11, 7) {real, imag} */,
  {32'hbf441204, 32'h3ff78d7d} /* (21, 11, 6) {real, imag} */,
  {32'hbf2fd878, 32'h3f9eb0b0} /* (21, 11, 5) {real, imag} */,
  {32'hbf411828, 32'hbf156bd0} /* (21, 11, 4) {real, imag} */,
  {32'hbf0d46be, 32'hbf58c49e} /* (21, 11, 3) {real, imag} */,
  {32'hbf4c422b, 32'h3f09331a} /* (21, 11, 2) {real, imag} */,
  {32'hbf9f2d5e, 32'hbe86cb60} /* (21, 11, 1) {real, imag} */,
  {32'hbf141088, 32'hbf1cded5} /* (21, 11, 0) {real, imag} */,
  {32'h3da3d280, 32'h3f4f4be5} /* (21, 10, 31) {real, imag} */,
  {32'h3e76cd70, 32'h3eb16642} /* (21, 10, 30) {real, imag} */,
  {32'h3fced138, 32'hbd6fef80} /* (21, 10, 29) {real, imag} */,
  {32'h4011b2ee, 32'hbeb4d7fa} /* (21, 10, 28) {real, imag} */,
  {32'h402bdc70, 32'hbf996d7e} /* (21, 10, 27) {real, imag} */,
  {32'h3fa56595, 32'h3e9dbd93} /* (21, 10, 26) {real, imag} */,
  {32'h3fdd44a4, 32'hbdbb1960} /* (21, 10, 25) {real, imag} */,
  {32'h3ed9a810, 32'hbef66f28} /* (21, 10, 24) {real, imag} */,
  {32'hbf73dcae, 32'hbfd91044} /* (21, 10, 23) {real, imag} */,
  {32'hbee7daca, 32'hbf4d2f1c} /* (21, 10, 22) {real, imag} */,
  {32'h3da6bc70, 32'hbf4cdf89} /* (21, 10, 21) {real, imag} */,
  {32'hbf4447da, 32'hbea13ca4} /* (21, 10, 20) {real, imag} */,
  {32'hc004bc0c, 32'hbe0c0500} /* (21, 10, 19) {real, imag} */,
  {32'hbfa13742, 32'h3f7bb4a4} /* (21, 10, 18) {real, imag} */,
  {32'hbf86d956, 32'h3ef1f93e} /* (21, 10, 17) {real, imag} */,
  {32'h3e717dc2, 32'hbfb1987e} /* (21, 10, 16) {real, imag} */,
  {32'hbf08724b, 32'hbf0d4d54} /* (21, 10, 15) {real, imag} */,
  {32'h3db126e4, 32'h3f88587a} /* (21, 10, 14) {real, imag} */,
  {32'h3e5ca94e, 32'h3f5cbcfe} /* (21, 10, 13) {real, imag} */,
  {32'hbd0ab5b4, 32'h3e934a1c} /* (21, 10, 12) {real, imag} */,
  {32'hbf30fc48, 32'hbf2de48c} /* (21, 10, 11) {real, imag} */,
  {32'hbf999ee0, 32'hbfac39fb} /* (21, 10, 10) {real, imag} */,
  {32'hbe9bf5a8, 32'hc000ede3} /* (21, 10, 9) {real, imag} */,
  {32'hbf93194e, 32'hbfa53168} /* (21, 10, 8) {real, imag} */,
  {32'hbfb690fe, 32'h3f3226f8} /* (21, 10, 7) {real, imag} */,
  {32'hbf4c3f97, 32'h4053f624} /* (21, 10, 6) {real, imag} */,
  {32'h3c26c000, 32'h40333dc2} /* (21, 10, 5) {real, imag} */,
  {32'h3f00aa70, 32'h3d5eed50} /* (21, 10, 4) {real, imag} */,
  {32'h3ce508a0, 32'h3e065060} /* (21, 10, 3) {real, imag} */,
  {32'h3eddfa84, 32'h4005383f} /* (21, 10, 2) {real, imag} */,
  {32'h3fbf0f12, 32'h3f64decf} /* (21, 10, 1) {real, imag} */,
  {32'h3fa2abc6, 32'h3ecf4f48} /* (21, 10, 0) {real, imag} */,
  {32'h3e9494ae, 32'h3faf200a} /* (21, 9, 31) {real, imag} */,
  {32'h3fe0e293, 32'h3f475e06} /* (21, 9, 30) {real, imag} */,
  {32'h4020f3b4, 32'hbf84c8b9} /* (21, 9, 29) {real, imag} */,
  {32'h3fedd5c6, 32'hbd154c60} /* (21, 9, 28) {real, imag} */,
  {32'h40076847, 32'hbe237a58} /* (21, 9, 27) {real, imag} */,
  {32'h3fb83da0, 32'hbf03e707} /* (21, 9, 26) {real, imag} */,
  {32'h3eb61aba, 32'hbec8dd70} /* (21, 9, 25) {real, imag} */,
  {32'h3ee3a084, 32'hbf3f20be} /* (21, 9, 24) {real, imag} */,
  {32'h3fc31b69, 32'hbfa5e4b2} /* (21, 9, 23) {real, imag} */,
  {32'h3e132280, 32'h3f11bee6} /* (21, 9, 22) {real, imag} */,
  {32'hbd2b1f40, 32'h3eb619e8} /* (21, 9, 21) {real, imag} */,
  {32'hbfdbc11c, 32'hbf1b69c8} /* (21, 9, 20) {real, imag} */,
  {32'hbfc5491e, 32'hbebd0c98} /* (21, 9, 19) {real, imag} */,
  {32'hbf790226, 32'h3ebc4c68} /* (21, 9, 18) {real, imag} */,
  {32'hbf5a672c, 32'hbe95b440} /* (21, 9, 17) {real, imag} */,
  {32'hbd2245a0, 32'hbfc3bae3} /* (21, 9, 16) {real, imag} */,
  {32'hc0038232, 32'hbfcb5464} /* (21, 9, 15) {real, imag} */,
  {32'hbf679ce6, 32'hbe9c85f0} /* (21, 9, 14) {real, imag} */,
  {32'hbf6a4016, 32'h3e41d300} /* (21, 9, 13) {real, imag} */,
  {32'hbef418e2, 32'h3e557368} /* (21, 9, 12) {real, imag} */,
  {32'hbf73e5ea, 32'hbf0ec174} /* (21, 9, 11) {real, imag} */,
  {32'hbfacaecc, 32'hbf8a67cc} /* (21, 9, 10) {real, imag} */,
  {32'hbf83cf46, 32'hbfe7bf9a} /* (21, 9, 9) {real, imag} */,
  {32'hbf8a9a40, 32'hbfaefe3c} /* (21, 9, 8) {real, imag} */,
  {32'hbf11f570, 32'hbf1a90ae} /* (21, 9, 7) {real, imag} */,
  {32'h3ec62096, 32'h3f8eafd8} /* (21, 9, 6) {real, imag} */,
  {32'h3edb198a, 32'h3fcdc4ee} /* (21, 9, 5) {real, imag} */,
  {32'h3f8350eb, 32'hbf024aba} /* (21, 9, 4) {real, imag} */,
  {32'h3f87df4f, 32'h3e9bc164} /* (21, 9, 3) {real, imag} */,
  {32'h3fbfe1df, 32'h3e1e89a0} /* (21, 9, 2) {real, imag} */,
  {32'h3fbbac79, 32'h3eef18e8} /* (21, 9, 1) {real, imag} */,
  {32'h3f614b2c, 32'h3f524e04} /* (21, 9, 0) {real, imag} */,
  {32'h3ee56df0, 32'h3f444a1e} /* (21, 8, 31) {real, imag} */,
  {32'h40112784, 32'h3fb73de4} /* (21, 8, 30) {real, imag} */,
  {32'h3fe7ff26, 32'h3e0cdd88} /* (21, 8, 29) {real, imag} */,
  {32'hbde55568, 32'h3e61f830} /* (21, 8, 28) {real, imag} */,
  {32'hbf23a4da, 32'h3f726a63} /* (21, 8, 27) {real, imag} */,
  {32'hbef8a899, 32'h3ea0f51c} /* (21, 8, 26) {real, imag} */,
  {32'h3e5dbde7, 32'hbdbed2a0} /* (21, 8, 25) {real, imag} */,
  {32'h3fce47e7, 32'h3d8eb5e0} /* (21, 8, 24) {real, imag} */,
  {32'h3fff9e99, 32'h3f24d148} /* (21, 8, 23) {real, imag} */,
  {32'h3f9a7d99, 32'h3fc5cc4b} /* (21, 8, 22) {real, imag} */,
  {32'h3f9f7b15, 32'h3fb620be} /* (21, 8, 21) {real, imag} */,
  {32'hbede5072, 32'hbf1c44bb} /* (21, 8, 20) {real, imag} */,
  {32'hbf475b76, 32'hbf81ff68} /* (21, 8, 19) {real, imag} */,
  {32'hbf39c51c, 32'hbedb7d20} /* (21, 8, 18) {real, imag} */,
  {32'hbfc86574, 32'hbe81b4f0} /* (21, 8, 17) {real, imag} */,
  {32'hbf79468e, 32'hbfc22c83} /* (21, 8, 16) {real, imag} */,
  {32'hbf9367e0, 32'hbfc83e70} /* (21, 8, 15) {real, imag} */,
  {32'hbfe07ba0, 32'hbf640966} /* (21, 8, 14) {real, imag} */,
  {32'hbf9a0a51, 32'h3d4536c0} /* (21, 8, 13) {real, imag} */,
  {32'h3f2a642e, 32'hbf56ac84} /* (21, 8, 12) {real, imag} */,
  {32'h3e7b7570, 32'hbf3bada8} /* (21, 8, 11) {real, imag} */,
  {32'h3f07edc3, 32'hbef9df28} /* (21, 8, 10) {real, imag} */,
  {32'hbef32a74, 32'h3ebe3f1c} /* (21, 8, 9) {real, imag} */,
  {32'hbf514986, 32'h3ea2ad04} /* (21, 8, 8) {real, imag} */,
  {32'hbf120134, 32'h3f4314ce} /* (21, 8, 7) {real, imag} */,
  {32'h3fb7d404, 32'h3f29fa64} /* (21, 8, 6) {real, imag} */,
  {32'h3fb2280d, 32'h3f358bf4} /* (21, 8, 5) {real, imag} */,
  {32'h3f91cb16, 32'h3fcff1ed} /* (21, 8, 4) {real, imag} */,
  {32'hbdd3d230, 32'h3fb02b48} /* (21, 8, 3) {real, imag} */,
  {32'h3ed05c30, 32'hbfa0d328} /* (21, 8, 2) {real, imag} */,
  {32'h3f640465, 32'hbf0bb4f6} /* (21, 8, 1) {real, imag} */,
  {32'h3e9daadd, 32'h3f704e0c} /* (21, 8, 0) {real, imag} */,
  {32'hbe805a35, 32'h3f031c5e} /* (21, 7, 31) {real, imag} */,
  {32'h3f611200, 32'h3f91225a} /* (21, 7, 30) {real, imag} */,
  {32'h3ef5a438, 32'h3fd5443f} /* (21, 7, 29) {real, imag} */,
  {32'hbf3ff870, 32'h3fe7d074} /* (21, 7, 28) {real, imag} */,
  {32'hbf88a77a, 32'h3f2c8d32} /* (21, 7, 27) {real, imag} */,
  {32'h3d67d060, 32'hbf66bada} /* (21, 7, 26) {real, imag} */,
  {32'h3fb8ea90, 32'hbea8f108} /* (21, 7, 25) {real, imag} */,
  {32'h3f8bf6d1, 32'h3f2c48cc} /* (21, 7, 24) {real, imag} */,
  {32'h3f051b76, 32'h3fc574f9} /* (21, 7, 23) {real, imag} */,
  {32'h3fb7f5fd, 32'h3f988ee7} /* (21, 7, 22) {real, imag} */,
  {32'h4026fbd0, 32'h3f725f17} /* (21, 7, 21) {real, imag} */,
  {32'h3fbb6894, 32'h3e101bb0} /* (21, 7, 20) {real, imag} */,
  {32'h3e9a1720, 32'hbf029746} /* (21, 7, 19) {real, imag} */,
  {32'hbf40d6e7, 32'h3e807db0} /* (21, 7, 18) {real, imag} */,
  {32'hbfbec4d2, 32'h3ea2a800} /* (21, 7, 17) {real, imag} */,
  {32'hbf74d784, 32'hbe9be720} /* (21, 7, 16) {real, imag} */,
  {32'hbf695d64, 32'h3eeb9bd6} /* (21, 7, 15) {real, imag} */,
  {32'hbfd5e427, 32'h3ef6827c} /* (21, 7, 14) {real, imag} */,
  {32'hc013ff91, 32'h3f396417} /* (21, 7, 13) {real, imag} */,
  {32'h3dc9e540, 32'hbf854b26} /* (21, 7, 12) {real, imag} */,
  {32'h3f275ac0, 32'hbf6e9228} /* (21, 7, 11) {real, imag} */,
  {32'h3f45169c, 32'h3ed4cac9} /* (21, 7, 10) {real, imag} */,
  {32'h3e8bfe6c, 32'h3f2b2346} /* (21, 7, 9) {real, imag} */,
  {32'h3e03187c, 32'h3d936f80} /* (21, 7, 8) {real, imag} */,
  {32'hbf8d5c39, 32'h3eafa0e4} /* (21, 7, 7) {real, imag} */,
  {32'h3f0a0c51, 32'h3f0708d4} /* (21, 7, 6) {real, imag} */,
  {32'h40067bef, 32'h3f9e303b} /* (21, 7, 5) {real, imag} */,
  {32'h3fef917f, 32'h3ff72593} /* (21, 7, 4) {real, imag} */,
  {32'hbf2143b4, 32'h3fa3d01f} /* (21, 7, 3) {real, imag} */,
  {32'h3f03ec70, 32'hbd237d30} /* (21, 7, 2) {real, imag} */,
  {32'h3f1a780c, 32'h3f87d910} /* (21, 7, 1) {real, imag} */,
  {32'h3eb3756e, 32'h3f366a2d} /* (21, 7, 0) {real, imag} */,
  {32'hbf294acc, 32'h3f52225a} /* (21, 6, 31) {real, imag} */,
  {32'hbcab6500, 32'h3fd500ea} /* (21, 6, 30) {real, imag} */,
  {32'h3f200d91, 32'h3fd1b04b} /* (21, 6, 29) {real, imag} */,
  {32'hbece8b06, 32'h3ff1c67b} /* (21, 6, 28) {real, imag} */,
  {32'hbf8479af, 32'h3ef1fff4} /* (21, 6, 27) {real, imag} */,
  {32'h3f732e72, 32'hbfd2330e} /* (21, 6, 26) {real, imag} */,
  {32'h3f48ba0e, 32'hbea301fc} /* (21, 6, 25) {real, imag} */,
  {32'h3d922590, 32'h3fb6dd76} /* (21, 6, 24) {real, imag} */,
  {32'h3e184b4c, 32'h3f22b2b8} /* (21, 6, 23) {real, imag} */,
  {32'hbded47d8, 32'hbe2a8ca0} /* (21, 6, 22) {real, imag} */,
  {32'h3f9fec16, 32'hbdcee290} /* (21, 6, 21) {real, imag} */,
  {32'h3f547396, 32'h3f420bcb} /* (21, 6, 20) {real, imag} */,
  {32'h3ef2fef2, 32'h3f31a74e} /* (21, 6, 19) {real, imag} */,
  {32'hbf1bd37a, 32'h3fdd687a} /* (21, 6, 18) {real, imag} */,
  {32'hbf827d02, 32'h3fbd134e} /* (21, 6, 17) {real, imag} */,
  {32'hbfb5fcc0, 32'h3ed53240} /* (21, 6, 16) {real, imag} */,
  {32'hbfadee94, 32'h3f8e6d5e} /* (21, 6, 15) {real, imag} */,
  {32'hbf627093, 32'h3f6ba929} /* (21, 6, 14) {real, imag} */,
  {32'hbfba142e, 32'h3fbfe378} /* (21, 6, 13) {real, imag} */,
  {32'hbf8d0920, 32'hbf44db4e} /* (21, 6, 12) {real, imag} */,
  {32'hbecd3844, 32'hbfc7209b} /* (21, 6, 11) {real, imag} */,
  {32'hbe13933c, 32'h3f435069} /* (21, 6, 10) {real, imag} */,
  {32'h3e939900, 32'h3f794726} /* (21, 6, 9) {real, imag} */,
  {32'h3ebc5e30, 32'hbf99f92b} /* (21, 6, 8) {real, imag} */,
  {32'hbedbd5bc, 32'hbf4eb41e} /* (21, 6, 7) {real, imag} */,
  {32'h3d170de0, 32'h3e9720e0} /* (21, 6, 6) {real, imag} */,
  {32'h3fb4a856, 32'h3fda3125} /* (21, 6, 5) {real, imag} */,
  {32'h3f8a7ab4, 32'h3f421754} /* (21, 6, 4) {real, imag} */,
  {32'h3dd14880, 32'hbf0a3af8} /* (21, 6, 3) {real, imag} */,
  {32'h3eff34a4, 32'hbe2bed90} /* (21, 6, 2) {real, imag} */,
  {32'h3f4f8fc8, 32'h3f724164} /* (21, 6, 1) {real, imag} */,
  {32'h3d7a7880, 32'h3edd9d54} /* (21, 6, 0) {real, imag} */,
  {32'h3ededf56, 32'h3f86b1f6} /* (21, 5, 31) {real, imag} */,
  {32'h3fa571ba, 32'h3fcb553a} /* (21, 5, 30) {real, imag} */,
  {32'h3f6082d2, 32'h3f187200} /* (21, 5, 29) {real, imag} */,
  {32'h3eab959c, 32'h3f882878} /* (21, 5, 28) {real, imag} */,
  {32'hbeb617b8, 32'h3c8bed80} /* (21, 5, 27) {real, imag} */,
  {32'h3f03f4a4, 32'hbf9327d6} /* (21, 5, 26) {real, imag} */,
  {32'h3d13a560, 32'h3f256fea} /* (21, 5, 25) {real, imag} */,
  {32'h3efd5074, 32'h3fa5546a} /* (21, 5, 24) {real, imag} */,
  {32'h3f56c8e4, 32'hbf016a76} /* (21, 5, 23) {real, imag} */,
  {32'h3f02e556, 32'hbfc1929d} /* (21, 5, 22) {real, imag} */,
  {32'h3f8c38b0, 32'hbf9ead0e} /* (21, 5, 21) {real, imag} */,
  {32'h3ec5cf84, 32'h3f34ec94} /* (21, 5, 20) {real, imag} */,
  {32'hbeae48d6, 32'hbd9bfa50} /* (21, 5, 19) {real, imag} */,
  {32'h3e7e0178, 32'h3e2d7f3c} /* (21, 5, 18) {real, imag} */,
  {32'h3ee6f485, 32'h3f235851} /* (21, 5, 17) {real, imag} */,
  {32'h3c8fbae0, 32'h3f90db24} /* (21, 5, 16) {real, imag} */,
  {32'hbfa19ec6, 32'h3f01291d} /* (21, 5, 15) {real, imag} */,
  {32'hbf82324e, 32'h3f4236fc} /* (21, 5, 14) {real, imag} */,
  {32'hbf336fe4, 32'h3fa3b10a} /* (21, 5, 13) {real, imag} */,
  {32'hc002e267, 32'hbf9b61a8} /* (21, 5, 12) {real, imag} */,
  {32'hc0204ce8, 32'hbf982d10} /* (21, 5, 11) {real, imag} */,
  {32'hbfb001d8, 32'h3fa6b5d3} /* (21, 5, 10) {real, imag} */,
  {32'hbf90e79a, 32'h3fc80771} /* (21, 5, 9) {real, imag} */,
  {32'hbf91fd65, 32'hbf5b4758} /* (21, 5, 8) {real, imag} */,
  {32'hbfa5b522, 32'hbf4402c5} /* (21, 5, 7) {real, imag} */,
  {32'hbfd1f866, 32'h3f6d09d5} /* (21, 5, 6) {real, imag} */,
  {32'hbe311958, 32'h3fdabad6} /* (21, 5, 5) {real, imag} */,
  {32'h3f8a228c, 32'h3f92bf7c} /* (21, 5, 4) {real, imag} */,
  {32'h3fdeedf9, 32'hbef3dc8b} /* (21, 5, 3) {real, imag} */,
  {32'h3fdff17a, 32'hbe563464} /* (21, 5, 2) {real, imag} */,
  {32'h3fd5616e, 32'hbd374ea0} /* (21, 5, 1) {real, imag} */,
  {32'h3f8122f4, 32'h3e300138} /* (21, 5, 0) {real, imag} */,
  {32'h3eed1088, 32'h3fbcbda8} /* (21, 4, 31) {real, imag} */,
  {32'h3efe1460, 32'h401b3268} /* (21, 4, 30) {real, imag} */,
  {32'h3f965bf9, 32'h3faa137a} /* (21, 4, 29) {real, imag} */,
  {32'h3f0f997a, 32'h3f46ff1a} /* (21, 4, 28) {real, imag} */,
  {32'h3fb7cd82, 32'h3fa7fefc} /* (21, 4, 27) {real, imag} */,
  {32'h3f8e5afe, 32'h3f6fc814} /* (21, 4, 26) {real, imag} */,
  {32'h3f0fc0b8, 32'h3f2095b4} /* (21, 4, 25) {real, imag} */,
  {32'h3e35e23c, 32'h3f00e882} /* (21, 4, 24) {real, imag} */,
  {32'hbd734e10, 32'hbeb21018} /* (21, 4, 23) {real, imag} */,
  {32'hbc849420, 32'hbf6a1c08} /* (21, 4, 22) {real, imag} */,
  {32'h3fd5f3dd, 32'hbf55b920} /* (21, 4, 21) {real, imag} */,
  {32'h402a77a0, 32'hbd7553e0} /* (21, 4, 20) {real, imag} */,
  {32'h3f81e119, 32'hbf85f908} /* (21, 4, 19) {real, imag} */,
  {32'h3f9be7fc, 32'hbf034d46} /* (21, 4, 18) {real, imag} */,
  {32'h3f36c00b, 32'hbecef42c} /* (21, 4, 17) {real, imag} */,
  {32'h3fccecdd, 32'h3d6d4180} /* (21, 4, 16) {real, imag} */,
  {32'h3daec1e4, 32'hbed5f256} /* (21, 4, 15) {real, imag} */,
  {32'hbfcdec19, 32'hbe85d748} /* (21, 4, 14) {real, imag} */,
  {32'hbf07c152, 32'hbe095454} /* (21, 4, 13) {real, imag} */,
  {32'hbfa9cd82, 32'hbf8b5dcf} /* (21, 4, 12) {real, imag} */,
  {32'hc0083ca8, 32'hbfc19fc4} /* (21, 4, 11) {real, imag} */,
  {32'hbf8e9795, 32'hbbbe1fc0} /* (21, 4, 10) {real, imag} */,
  {32'hbfee0ccb, 32'h3eda334d} /* (21, 4, 9) {real, imag} */,
  {32'hc007a7a5, 32'hbfd2ab8b} /* (21, 4, 8) {real, imag} */,
  {32'hbfd6252a, 32'hbf9d7c30} /* (21, 4, 7) {real, imag} */,
  {32'hc020abf3, 32'hbc54b3c0} /* (21, 4, 6) {real, imag} */,
  {32'hbeb68144, 32'h3f60c67a} /* (21, 4, 5) {real, imag} */,
  {32'h401501da, 32'h3f8ffe62} /* (21, 4, 4) {real, imag} */,
  {32'h3fdc3d95, 32'hbe9539c8} /* (21, 4, 3) {real, imag} */,
  {32'h3fcf2988, 32'hbfa89bb4} /* (21, 4, 2) {real, imag} */,
  {32'h3fad65b4, 32'hbf6087bc} /* (21, 4, 1) {real, imag} */,
  {32'h3f99211d, 32'h3f0110a4} /* (21, 4, 0) {real, imag} */,
  {32'h3eb8ccac, 32'h3f028a6a} /* (21, 3, 31) {real, imag} */,
  {32'h3f029ec4, 32'h3ff60055} /* (21, 3, 30) {real, imag} */,
  {32'h3f28f9d4, 32'h3fb383f2} /* (21, 3, 29) {real, imag} */,
  {32'h3ef53428, 32'h3dc32f70} /* (21, 3, 28) {real, imag} */,
  {32'h3f93f131, 32'h3f2bf704} /* (21, 3, 27) {real, imag} */,
  {32'h3ebcf694, 32'h3fc58b62} /* (21, 3, 26) {real, imag} */,
  {32'h3ead9504, 32'h3f7f52aa} /* (21, 3, 25) {real, imag} */,
  {32'hbf0c73bf, 32'h3f6357b6} /* (21, 3, 24) {real, imag} */,
  {32'h3f3cc993, 32'h3ec6f95c} /* (21, 3, 23) {real, imag} */,
  {32'h3f871d0d, 32'h3e1ff580} /* (21, 3, 22) {real, imag} */,
  {32'h3ed475b6, 32'h3f58ce61} /* (21, 3, 21) {real, imag} */,
  {32'h3fc3ae62, 32'h3f873ea2} /* (21, 3, 20) {real, imag} */,
  {32'h3fc718e1, 32'hbf175fbe} /* (21, 3, 19) {real, imag} */,
  {32'h3fae6b57, 32'hbe9595e8} /* (21, 3, 18) {real, imag} */,
  {32'h3f86b62b, 32'h3ddee2e0} /* (21, 3, 17) {real, imag} */,
  {32'h3fb6540d, 32'h3d8ddf60} /* (21, 3, 16) {real, imag} */,
  {32'h3fb4e27a, 32'hbf3fed0f} /* (21, 3, 15) {real, imag} */,
  {32'hbe98be80, 32'hbebc1792} /* (21, 3, 14) {real, imag} */,
  {32'hbe035890, 32'h3f882cb6} /* (21, 3, 13) {real, imag} */,
  {32'h3e7356d2, 32'hbeb1acb0} /* (21, 3, 12) {real, imag} */,
  {32'hbec7065e, 32'hc04627c4} /* (21, 3, 11) {real, imag} */,
  {32'hbf838738, 32'hbf296aab} /* (21, 3, 10) {real, imag} */,
  {32'hbfd415dd, 32'hbe914320} /* (21, 3, 9) {real, imag} */,
  {32'hbff2463c, 32'hbfc93341} /* (21, 3, 8) {real, imag} */,
  {32'hbfab509b, 32'hc007e54d} /* (21, 3, 7) {real, imag} */,
  {32'hbfd691e0, 32'h3e907502} /* (21, 3, 6) {real, imag} */,
  {32'h3f7f71ee, 32'h400ded3a} /* (21, 3, 5) {real, imag} */,
  {32'h3fecf8ba, 32'h3ff2a490} /* (21, 3, 4) {real, imag} */,
  {32'h3f3569b8, 32'h3f5a21b8} /* (21, 3, 3) {real, imag} */,
  {32'hbe084940, 32'h3ec4fe68} /* (21, 3, 2) {real, imag} */,
  {32'hbd4d9d10, 32'hbbc0b300} /* (21, 3, 1) {real, imag} */,
  {32'h3e3dd004, 32'h3f6c53af} /* (21, 3, 0) {real, imag} */,
  {32'h3fc97986, 32'hbef78db0} /* (21, 2, 31) {real, imag} */,
  {32'h400fd198, 32'h3e63ec30} /* (21, 2, 30) {real, imag} */,
  {32'h3c128400, 32'h3f93ac1f} /* (21, 2, 29) {real, imag} */,
  {32'h3f450b70, 32'h3f5e23b1} /* (21, 2, 28) {real, imag} */,
  {32'hbe9c6a00, 32'h3f020146} /* (21, 2, 27) {real, imag} */,
  {32'hbf824b40, 32'h3faebe4b} /* (21, 2, 26) {real, imag} */,
  {32'h3f8918aa, 32'h3fabc074} /* (21, 2, 25) {real, imag} */,
  {32'h3f9eb7b7, 32'h3f519638} /* (21, 2, 24) {real, imag} */,
  {32'h3fdf6082, 32'h3e893fe0} /* (21, 2, 23) {real, imag} */,
  {32'h3f9c58fe, 32'h3f87848d} /* (21, 2, 22) {real, imag} */,
  {32'h3e4010a0, 32'h3f76ecc4} /* (21, 2, 21) {real, imag} */,
  {32'h3f0c232a, 32'h3f9d3729} /* (21, 2, 20) {real, imag} */,
  {32'h3f804a16, 32'h3f50750c} /* (21, 2, 19) {real, imag} */,
  {32'h4008bf0c, 32'h400147e4} /* (21, 2, 18) {real, imag} */,
  {32'h4039b907, 32'h401b020e} /* (21, 2, 17) {real, imag} */,
  {32'h3f349eae, 32'h3f66c438} /* (21, 2, 16) {real, imag} */,
  {32'h3f954adf, 32'hbf32e94c} /* (21, 2, 15) {real, imag} */,
  {32'h3f90e2b6, 32'hbf860903} /* (21, 2, 14) {real, imag} */,
  {32'hbed4eea2, 32'h3f2e1092} /* (21, 2, 13) {real, imag} */,
  {32'hbf79b15e, 32'hbe6e8810} /* (21, 2, 12) {real, imag} */,
  {32'h3e1ebbf0, 32'hc02aaaa4} /* (21, 2, 11) {real, imag} */,
  {32'h3df59af0, 32'h3f1c0f43} /* (21, 2, 10) {real, imag} */,
  {32'hbf9ecdfc, 32'h3f87a40e} /* (21, 2, 9) {real, imag} */,
  {32'hbfd13872, 32'hbe7ed890} /* (21, 2, 8) {real, imag} */,
  {32'hbf4c46f7, 32'hbf10b210} /* (21, 2, 7) {real, imag} */,
  {32'hbf331587, 32'h3f7496f2} /* (21, 2, 6) {real, imag} */,
  {32'h3ea5ade2, 32'h3fdbfabb} /* (21, 2, 5) {real, imag} */,
  {32'h3fcd1ab0, 32'h3f4dfaba} /* (21, 2, 4) {real, imag} */,
  {32'h3fe72109, 32'hbb67a400} /* (21, 2, 3) {real, imag} */,
  {32'h3fb1b06d, 32'hbd6986e0} /* (21, 2, 2) {real, imag} */,
  {32'h3fa77178, 32'h3ef06930} /* (21, 2, 1) {real, imag} */,
  {32'h3f158dc0, 32'h3f855308} /* (21, 2, 0) {real, imag} */,
  {32'h3f8d755a, 32'h3f267d22} /* (21, 1, 31) {real, imag} */,
  {32'h3f9322b4, 32'h3e45973c} /* (21, 1, 30) {real, imag} */,
  {32'hbf11749f, 32'hbf7bafc8} /* (21, 1, 29) {real, imag} */,
  {32'h3f0b83ec, 32'hbe9aeee4} /* (21, 1, 28) {real, imag} */,
  {32'hbee76160, 32'h3d9d3500} /* (21, 1, 27) {real, imag} */,
  {32'hbd626580, 32'h3f458ad6} /* (21, 1, 26) {real, imag} */,
  {32'h3fd3f231, 32'h3f415f5a} /* (21, 1, 25) {real, imag} */,
  {32'h4007c814, 32'hbfaead02} /* (21, 1, 24) {real, imag} */,
  {32'h3fd0c93c, 32'hbf94a5d2} /* (21, 1, 23) {real, imag} */,
  {32'h3faabf9e, 32'h3f778504} /* (21, 1, 22) {real, imag} */,
  {32'h3ee6c0ec, 32'h3f073098} /* (21, 1, 21) {real, imag} */,
  {32'h3ee21bb8, 32'h3eda2350} /* (21, 1, 20) {real, imag} */,
  {32'h3ea6ecc0, 32'h3f45dcc8} /* (21, 1, 19) {real, imag} */,
  {32'h3f961c11, 32'h40251429} /* (21, 1, 18) {real, imag} */,
  {32'h4013a26e, 32'h40517adc} /* (21, 1, 17) {real, imag} */,
  {32'h3e9481dc, 32'h3ec218b0} /* (21, 1, 16) {real, imag} */,
  {32'hbe9e9dd2, 32'hbfb6922f} /* (21, 1, 15) {real, imag} */,
  {32'hbf7f7a8a, 32'hbf8116a4} /* (21, 1, 14) {real, imag} */,
  {32'hbf716f06, 32'h3f0879be} /* (21, 1, 13) {real, imag} */,
  {32'hbef01db2, 32'hbea805ec} /* (21, 1, 12) {real, imag} */,
  {32'h3e5da128, 32'hbfe9287a} /* (21, 1, 11) {real, imag} */,
  {32'h3e0a5f30, 32'h3dda77c0} /* (21, 1, 10) {real, imag} */,
  {32'hbf50aed4, 32'h3dec3640} /* (21, 1, 9) {real, imag} */,
  {32'hbf1cabc4, 32'hbfa6ea5c} /* (21, 1, 8) {real, imag} */,
  {32'hbe72fe08, 32'hbe4a7ed0} /* (21, 1, 7) {real, imag} */,
  {32'h3e43e4f8, 32'hbf27634e} /* (21, 1, 6) {real, imag} */,
  {32'h3e9a1cf7, 32'hbf2f5d91} /* (21, 1, 5) {real, imag} */,
  {32'h4013c52e, 32'hbd92f774} /* (21, 1, 4) {real, imag} */,
  {32'h4004c956, 32'hbf3228ef} /* (21, 1, 3) {real, imag} */,
  {32'h3f9a5ca4, 32'hbf3b5e1a} /* (21, 1, 2) {real, imag} */,
  {32'h3f41c0a2, 32'h3f99678c} /* (21, 1, 1) {real, imag} */,
  {32'h3f5812b7, 32'h3fcc6d88} /* (21, 1, 0) {real, imag} */,
  {32'h3e8ac790, 32'h3f2d71c9} /* (21, 0, 31) {real, imag} */,
  {32'h3db8a338, 32'hbdf347ec} /* (21, 0, 30) {real, imag} */,
  {32'hbf4719e8, 32'hbfd36387} /* (21, 0, 29) {real, imag} */,
  {32'hbec729bc, 32'hbf592af3} /* (21, 0, 28) {real, imag} */,
  {32'hbeca1d9a, 32'hbf27f0fe} /* (21, 0, 27) {real, imag} */,
  {32'h3e0453e8, 32'h3d56d720} /* (21, 0, 26) {real, imag} */,
  {32'h3f41a332, 32'h3e28e518} /* (21, 0, 25) {real, imag} */,
  {32'h3fb196c2, 32'hbf808d29} /* (21, 0, 24) {real, imag} */,
  {32'h3fe3d1d2, 32'hbf1165c8} /* (21, 0, 23) {real, imag} */,
  {32'h3fb1b883, 32'h3ec84b68} /* (21, 0, 22) {real, imag} */,
  {32'h3ebb3563, 32'h3eb6c160} /* (21, 0, 21) {real, imag} */,
  {32'h3e6fd400, 32'hbdfe8980} /* (21, 0, 20) {real, imag} */,
  {32'hbe8d1bc4, 32'hbe8edb8c} /* (21, 0, 19) {real, imag} */,
  {32'hbe781594, 32'h3f81947c} /* (21, 0, 18) {real, imag} */,
  {32'h3d7bb9e0, 32'h3f866d84} /* (21, 0, 17) {real, imag} */,
  {32'h3e1c3fb8, 32'hbefa97ea} /* (21, 0, 16) {real, imag} */,
  {32'h3e8c4c54, 32'hbf00282b} /* (21, 0, 15) {real, imag} */,
  {32'hbf1368cb, 32'hbd0ae6d0} /* (21, 0, 14) {real, imag} */,
  {32'hbf556cd3, 32'h3c1cc940} /* (21, 0, 13) {real, imag} */,
  {32'hbeff9b27, 32'hbf0c4bb0} /* (21, 0, 12) {real, imag} */,
  {32'hbec6eb97, 32'hbf0d53fd} /* (21, 0, 11) {real, imag} */,
  {32'hbeeb33b0, 32'h3c8b9340} /* (21, 0, 10) {real, imag} */,
  {32'hbec551fa, 32'h3e5395d4} /* (21, 0, 9) {real, imag} */,
  {32'h3ec9ac2f, 32'h3dd91380} /* (21, 0, 8) {real, imag} */,
  {32'hbf0ff754, 32'h3f3b389a} /* (21, 0, 7) {real, imag} */,
  {32'hbe7a0374, 32'hbe6ec70e} /* (21, 0, 6) {real, imag} */,
  {32'h3fd1eb48, 32'hbe971e4a} /* (21, 0, 5) {real, imag} */,
  {32'h40068ab7, 32'h3e6d6485} /* (21, 0, 4) {real, imag} */,
  {32'h3f99c879, 32'h3ca58ca0} /* (21, 0, 3) {real, imag} */,
  {32'h3f7db2cc, 32'hbe2c34ec} /* (21, 0, 2) {real, imag} */,
  {32'h3f5e1580, 32'h3e5c2920} /* (21, 0, 1) {real, imag} */,
  {32'h3f164d6d, 32'h3eff3c86} /* (21, 0, 0) {real, imag} */,
  {32'hbea9e695, 32'h3e6f9b68} /* (20, 31, 31) {real, imag} */,
  {32'hbe910638, 32'hbe3d1720} /* (20, 31, 30) {real, imag} */,
  {32'hbf1680c0, 32'hbebe7240} /* (20, 31, 29) {real, imag} */,
  {32'hbf2d9604, 32'hbefa8178} /* (20, 31, 28) {real, imag} */,
  {32'hbf7ae8e6, 32'hbdd7d300} /* (20, 31, 27) {real, imag} */,
  {32'h3e836b14, 32'h3f6c9446} /* (20, 31, 26) {real, imag} */,
  {32'h3fa0f739, 32'h3f956bae} /* (20, 31, 25) {real, imag} */,
  {32'h3f8e2b03, 32'h3cb378c0} /* (20, 31, 24) {real, imag} */,
  {32'hbcae3d80, 32'hbf5bbcb6} /* (20, 31, 23) {real, imag} */,
  {32'hbefc9004, 32'hbebd1818} /* (20, 31, 22) {real, imag} */,
  {32'h3e161c31, 32'h3dd4aae0} /* (20, 31, 21) {real, imag} */,
  {32'hbe307026, 32'h3f041eba} /* (20, 31, 20) {real, imag} */,
  {32'h3e40cf6d, 32'h3ef99428} /* (20, 31, 19) {real, imag} */,
  {32'hbe5d9112, 32'h3f0c4bbe} /* (20, 31, 18) {real, imag} */,
  {32'hbf14202a, 32'hbe9416dc} /* (20, 31, 17) {real, imag} */,
  {32'hbf79aedc, 32'hbe323b7a} /* (20, 31, 16) {real, imag} */,
  {32'hbee85e5a, 32'h3dc71b30} /* (20, 31, 15) {real, imag} */,
  {32'h3ef149d2, 32'hbe5c5ef0} /* (20, 31, 14) {real, imag} */,
  {32'hbe913dba, 32'hbec6bd6c} /* (20, 31, 13) {real, imag} */,
  {32'h3f04d154, 32'h3e311f70} /* (20, 31, 12) {real, imag} */,
  {32'h3e63f78c, 32'hbe086860} /* (20, 31, 11) {real, imag} */,
  {32'h3e49b825, 32'h3eb39fb8} /* (20, 31, 10) {real, imag} */,
  {32'hbd7205e0, 32'h3ef781f8} /* (20, 31, 9) {real, imag} */,
  {32'hbf72ce5a, 32'h3ea06ba8} /* (20, 31, 8) {real, imag} */,
  {32'hbf61e8ed, 32'hbefbb536} /* (20, 31, 7) {real, imag} */,
  {32'hbea0bfac, 32'hbf05410f} /* (20, 31, 6) {real, imag} */,
  {32'h3e8da598, 32'hbf1be4c4} /* (20, 31, 5) {real, imag} */,
  {32'h3e2e4728, 32'hbdd2af58} /* (20, 31, 4) {real, imag} */,
  {32'hbf65cd10, 32'h3ee603d8} /* (20, 31, 3) {real, imag} */,
  {32'hbfa2c183, 32'h3eadd3c8} /* (20, 31, 2) {real, imag} */,
  {32'hbe95dbc0, 32'hbf44e696} /* (20, 31, 1) {real, imag} */,
  {32'h3e20c92c, 32'hbe6f4700} /* (20, 31, 0) {real, imag} */,
  {32'h3e2b92b0, 32'h3f1208f8} /* (20, 30, 31) {real, imag} */,
  {32'h3da3e300, 32'h3f512438} /* (20, 30, 30) {real, imag} */,
  {32'hbde75ce0, 32'h3f3953ac} /* (20, 30, 29) {real, imag} */,
  {32'hbd92b8c0, 32'hbe83dc90} /* (20, 30, 28) {real, imag} */,
  {32'hbf88983c, 32'h3eaaf4d8} /* (20, 30, 27) {real, imag} */,
  {32'h3e8987d6, 32'h3fef51a8} /* (20, 30, 26) {real, imag} */,
  {32'h3fde443d, 32'h3fb732d8} /* (20, 30, 25) {real, imag} */,
  {32'h3fdb9e9a, 32'h3e890888} /* (20, 30, 24) {real, imag} */,
  {32'h3e217078, 32'hbf80e888} /* (20, 30, 23) {real, imag} */,
  {32'hbf157b78, 32'hbec1ce00} /* (20, 30, 22) {real, imag} */,
  {32'h3f5d14de, 32'hbe25f8c0} /* (20, 30, 21) {real, imag} */,
  {32'h3edf509e, 32'h3f503f78} /* (20, 30, 20) {real, imag} */,
  {32'h3eaddb58, 32'h3ea20f88} /* (20, 30, 19) {real, imag} */,
  {32'hbd974b2e, 32'h3cfbab00} /* (20, 30, 18) {real, imag} */,
  {32'hbc8076a0, 32'h3de27960} /* (20, 30, 17) {real, imag} */,
  {32'hbf22b5a2, 32'h3f130180} /* (20, 30, 16) {real, imag} */,
  {32'hbf10c1fe, 32'hbec01138} /* (20, 30, 15) {real, imag} */,
  {32'h3e15e158, 32'hbfe8a7f4} /* (20, 30, 14) {real, imag} */,
  {32'hbe45747f, 32'hbf98613d} /* (20, 30, 13) {real, imag} */,
  {32'h3f5a307c, 32'hbe8f1db0} /* (20, 30, 12) {real, imag} */,
  {32'h3ec0060c, 32'hbe8d6fe0} /* (20, 30, 11) {real, imag} */,
  {32'h3f69a261, 32'h3ecd548d} /* (20, 30, 10) {real, imag} */,
  {32'h3e819f20, 32'hbdb15ae0} /* (20, 30, 9) {real, imag} */,
  {32'hbf651cd0, 32'hbfa2c9e0} /* (20, 30, 8) {real, imag} */,
  {32'hbf8a1ddd, 32'hbfe389e1} /* (20, 30, 7) {real, imag} */,
  {32'hbe4dc264, 32'hbfd3e57e} /* (20, 30, 6) {real, imag} */,
  {32'hbddb6140, 32'hbf96e9b4} /* (20, 30, 5) {real, imag} */,
  {32'hbe8f79ac, 32'hbda33540} /* (20, 30, 4) {real, imag} */,
  {32'hbf4fb8d8, 32'h3d233040} /* (20, 30, 3) {real, imag} */,
  {32'hbf9ea86d, 32'hbea5e7a0} /* (20, 30, 2) {real, imag} */,
  {32'h3ea0de94, 32'hbedfc538} /* (20, 30, 1) {real, imag} */,
  {32'h3f20382e, 32'h3e9de794} /* (20, 30, 0) {real, imag} */,
  {32'h3f06605e, 32'hbe3456a8} /* (20, 29, 31) {real, imag} */,
  {32'h3e7590b8, 32'h3f94dd3c} /* (20, 29, 30) {real, imag} */,
  {32'hbeca0f84, 32'h3fd189eb} /* (20, 29, 29) {real, imag} */,
  {32'hbf9a3e50, 32'h3e653380} /* (20, 29, 28) {real, imag} */,
  {32'hbf210892, 32'hbe1226a0} /* (20, 29, 27) {real, imag} */,
  {32'h3f2463c8, 32'h3ee73988} /* (20, 29, 26) {real, imag} */,
  {32'h3f11f2f2, 32'h3f6a7362} /* (20, 29, 25) {real, imag} */,
  {32'h3f33140c, 32'h3f5ddb74} /* (20, 29, 24) {real, imag} */,
  {32'h3d860390, 32'hbe9bdfb8} /* (20, 29, 23) {real, imag} */,
  {32'h3ef5d8c6, 32'hbf57ee90} /* (20, 29, 22) {real, imag} */,
  {32'h3fe9304b, 32'hbf016e74} /* (20, 29, 21) {real, imag} */,
  {32'h3fb1a026, 32'h3fa3f600} /* (20, 29, 20) {real, imag} */,
  {32'h3f89ba36, 32'h3f352474} /* (20, 29, 19) {real, imag} */,
  {32'h3ef60132, 32'h3bc3d200} /* (20, 29, 18) {real, imag} */,
  {32'hbc9df500, 32'h3f249564} /* (20, 29, 17) {real, imag} */,
  {32'h3ee3664a, 32'h3bd5be00} /* (20, 29, 16) {real, imag} */,
  {32'h3e8e14fa, 32'h3d5db900} /* (20, 29, 15) {real, imag} */,
  {32'h3ee2f1a0, 32'hbecab4a0} /* (20, 29, 14) {real, imag} */,
  {32'h3f2800f6, 32'hbcd3bc00} /* (20, 29, 13) {real, imag} */,
  {32'h3fcbc7b7, 32'h3f20eef8} /* (20, 29, 12) {real, imag} */,
  {32'h3f80d36f, 32'h3ee036fc} /* (20, 29, 11) {real, imag} */,
  {32'h3fb59e1c, 32'hbefd2b82} /* (20, 29, 10) {real, imag} */,
  {32'h3f3f07dc, 32'hbf1babb0} /* (20, 29, 9) {real, imag} */,
  {32'h3ece9af8, 32'hbf9befa0} /* (20, 29, 8) {real, imag} */,
  {32'hbf788c54, 32'hbfabf3d2} /* (20, 29, 7) {real, imag} */,
  {32'hbf9be379, 32'hbf57ffee} /* (20, 29, 6) {real, imag} */,
  {32'hbf3f901e, 32'hbf9935c8} /* (20, 29, 5) {real, imag} */,
  {32'hbf22602e, 32'hbe25da90} /* (20, 29, 4) {real, imag} */,
  {32'hbfccc134, 32'h3e363c10} /* (20, 29, 3) {real, imag} */,
  {32'hbf49433e, 32'hbf7e215a} /* (20, 29, 2) {real, imag} */,
  {32'h3f0c9a27, 32'hbf544ec6} /* (20, 29, 1) {real, imag} */,
  {32'h3f255ac6, 32'hbed51b0c} /* (20, 29, 0) {real, imag} */,
  {32'hbe5defa8, 32'hbdba2384} /* (20, 28, 31) {real, imag} */,
  {32'hbe28e640, 32'h3f810032} /* (20, 28, 30) {real, imag} */,
  {32'hbf2c6330, 32'h3f5c2378} /* (20, 28, 29) {real, imag} */,
  {32'hbfd0af34, 32'hbf25e12c} /* (20, 28, 28) {real, imag} */,
  {32'hbe84ee90, 32'hbf135ebc} /* (20, 28, 27) {real, imag} */,
  {32'h3e35c788, 32'h3ec16bd0} /* (20, 28, 26) {real, imag} */,
  {32'h3f024590, 32'h3e9ccaa8} /* (20, 28, 25) {real, imag} */,
  {32'h3cb31f60, 32'hbda76540} /* (20, 28, 24) {real, imag} */,
  {32'hbf4d7ede, 32'hbe34c020} /* (20, 28, 23) {real, imag} */,
  {32'hbefe0908, 32'hbf196ef0} /* (20, 28, 22) {real, imag} */,
  {32'h3f813959, 32'hbf1ac8a4} /* (20, 28, 21) {real, imag} */,
  {32'h3f9091e8, 32'h3ef3a650} /* (20, 28, 20) {real, imag} */,
  {32'h3f6f666a, 32'h3ef1d234} /* (20, 28, 19) {real, imag} */,
  {32'h3ee4a708, 32'hbe8fe9e8} /* (20, 28, 18) {real, imag} */,
  {32'h3e539920, 32'hbf4a1ea0} /* (20, 28, 17) {real, imag} */,
  {32'h3f2b669c, 32'hbf022ab8} /* (20, 28, 16) {real, imag} */,
  {32'h3eb72d64, 32'h3f39e6e2} /* (20, 28, 15) {real, imag} */,
  {32'h3e072ad0, 32'hbea1509c} /* (20, 28, 14) {real, imag} */,
  {32'h3ec5d548, 32'h3dbda850} /* (20, 28, 13) {real, imag} */,
  {32'h3f8c902b, 32'h3eef2044} /* (20, 28, 12) {real, imag} */,
  {32'h3dd936d9, 32'hbf255ef6} /* (20, 28, 11) {real, imag} */,
  {32'hbe7f5050, 32'hbc3c6c00} /* (20, 28, 10) {real, imag} */,
  {32'h3d36e440, 32'h3fab0c87} /* (20, 28, 9) {real, imag} */,
  {32'h3f447798, 32'h3f7333f4} /* (20, 28, 8) {real, imag} */,
  {32'hbe272da8, 32'h3cba8500} /* (20, 28, 7) {real, imag} */,
  {32'hbef04a70, 32'h3dd51320} /* (20, 28, 6) {real, imag} */,
  {32'h3ddb3b30, 32'hbe920974} /* (20, 28, 5) {real, imag} */,
  {32'hbf08ceec, 32'h3ea05314} /* (20, 28, 4) {real, imag} */,
  {32'hbfced17a, 32'h3fa4821f} /* (20, 28, 3) {real, imag} */,
  {32'h3d586880, 32'h3f1115e2} /* (20, 28, 2) {real, imag} */,
  {32'hbdca22c0, 32'hbf78b8f0} /* (20, 28, 1) {real, imag} */,
  {32'hbe860913, 32'hbf806796} /* (20, 28, 0) {real, imag} */,
  {32'hbdb35d2c, 32'h3d4a32e0} /* (20, 27, 31) {real, imag} */,
  {32'h3dbf2480, 32'h3f765da0} /* (20, 27, 30) {real, imag} */,
  {32'h3e1d5e50, 32'h3f04d628} /* (20, 27, 29) {real, imag} */,
  {32'h3f0863b2, 32'hbe628268} /* (20, 27, 28) {real, imag} */,
  {32'h3efc39dc, 32'hbf0867e0} /* (20, 27, 27) {real, imag} */,
  {32'hbe6b4550, 32'h3f273710} /* (20, 27, 26) {real, imag} */,
  {32'hbeb0f567, 32'h3d09d780} /* (20, 27, 25) {real, imag} */,
  {32'hbf064090, 32'hbd853050} /* (20, 27, 24) {real, imag} */,
  {32'h3e83a05c, 32'hbed28f90} /* (20, 27, 23) {real, imag} */,
  {32'h3d596a00, 32'hbeae02a8} /* (20, 27, 22) {real, imag} */,
  {32'h3ef73d84, 32'hbd9de840} /* (20, 27, 21) {real, imag} */,
  {32'h3f4237ee, 32'h3f32cc5a} /* (20, 27, 20) {real, imag} */,
  {32'hbe5f3dd0, 32'h3f17c366} /* (20, 27, 19) {real, imag} */,
  {32'hbf7626f0, 32'h3eb4aabc} /* (20, 27, 18) {real, imag} */,
  {32'hbf6a9358, 32'h3f72af46} /* (20, 27, 17) {real, imag} */,
  {32'hbd9534b0, 32'h3eeaf778} /* (20, 27, 16) {real, imag} */,
  {32'hbcb203a0, 32'h3f97651e} /* (20, 27, 15) {real, imag} */,
  {32'hbea23d8c, 32'hbee03230} /* (20, 27, 14) {real, imag} */,
  {32'h3b870880, 32'hbf1b8eec} /* (20, 27, 13) {real, imag} */,
  {32'h3ec1a6e9, 32'hbecb4c50} /* (20, 27, 12) {real, imag} */,
  {32'hbe8bc558, 32'hbfe249c5} /* (20, 27, 11) {real, imag} */,
  {32'hbe826d54, 32'hbf1ba740} /* (20, 27, 10) {real, imag} */,
  {32'h3f21f38e, 32'hbebcc0f8} /* (20, 27, 9) {real, imag} */,
  {32'h3f7292b8, 32'h3e47c450} /* (20, 27, 8) {real, imag} */,
  {32'h3f6474d0, 32'h3f684e04} /* (20, 27, 7) {real, imag} */,
  {32'h3dda6ef0, 32'h3f845e22} /* (20, 27, 6) {real, imag} */,
  {32'hbe117500, 32'hbda81fc0} /* (20, 27, 5) {real, imag} */,
  {32'h3f0e154c, 32'hbe764b38} /* (20, 27, 4) {real, imag} */,
  {32'h3eecd5b8, 32'h3e7643f0} /* (20, 27, 3) {real, imag} */,
  {32'h3e8ac608, 32'h3f9d9aad} /* (20, 27, 2) {real, imag} */,
  {32'hbf234a02, 32'hbd2639a0} /* (20, 27, 1) {real, imag} */,
  {32'hbf0869aa, 32'hbf02339a} /* (20, 27, 0) {real, imag} */,
  {32'h3e3b6d04, 32'h3f17f480} /* (20, 26, 31) {real, imag} */,
  {32'h3e7ef6f0, 32'h3f975ca1} /* (20, 26, 30) {real, imag} */,
  {32'h3f30514e, 32'h3e35e7d0} /* (20, 26, 29) {real, imag} */,
  {32'h3f45f342, 32'h3f5d2864} /* (20, 26, 28) {real, imag} */,
  {32'hbed5a130, 32'h3f380f52} /* (20, 26, 27) {real, imag} */,
  {32'hbe2292c0, 32'h3e523230} /* (20, 26, 26) {real, imag} */,
  {32'hbeae5f40, 32'h3d957da0} /* (20, 26, 25) {real, imag} */,
  {32'hbf844be5, 32'h3f20a9e5} /* (20, 26, 24) {real, imag} */,
  {32'h3f087f76, 32'hbf1479d0} /* (20, 26, 23) {real, imag} */,
  {32'hbc08f380, 32'hbf3af7ea} /* (20, 26, 22) {real, imag} */,
  {32'hbf8aeeea, 32'h3edf2d64} /* (20, 26, 21) {real, imag} */,
  {32'h3ececc42, 32'h3e777f18} /* (20, 26, 20) {real, imag} */,
  {32'h3f3c00f0, 32'hbdf07370} /* (20, 26, 19) {real, imag} */,
  {32'h3e471aa8, 32'h3e6255e0} /* (20, 26, 18) {real, imag} */,
  {32'h3eca38e2, 32'h3f8f210d} /* (20, 26, 17) {real, imag} */,
  {32'h3f2d9408, 32'h3f3d569e} /* (20, 26, 16) {real, imag} */,
  {32'hbe33edee, 32'h3e811da8} /* (20, 26, 15) {real, imag} */,
  {32'hbf08a59a, 32'hbf2da52c} /* (20, 26, 14) {real, imag} */,
  {32'hbdeb1e68, 32'hbf280684} /* (20, 26, 13) {real, imag} */,
  {32'h3ca54b18, 32'hbf4e3c0e} /* (20, 26, 12) {real, imag} */,
  {32'hbeda1d30, 32'hbf624952} /* (20, 26, 11) {real, imag} */,
  {32'hbde7b3ac, 32'hbdd3b150} /* (20, 26, 10) {real, imag} */,
  {32'hbeed7060, 32'hbfc40704} /* (20, 26, 9) {real, imag} */,
  {32'h3dd29420, 32'hbf5481f0} /* (20, 26, 8) {real, imag} */,
  {32'h3f61d61d, 32'h3f5e60fc} /* (20, 26, 7) {real, imag} */,
  {32'h3dc22428, 32'h3fac1606} /* (20, 26, 6) {real, imag} */,
  {32'h3d4603a0, 32'hbe066500} /* (20, 26, 5) {real, imag} */,
  {32'h3f4b38fd, 32'hbe9ea0d0} /* (20, 26, 4) {real, imag} */,
  {32'h3c8d50c0, 32'h3e98af64} /* (20, 26, 3) {real, imag} */,
  {32'hbea53f4a, 32'h3f3b1650} /* (20, 26, 2) {real, imag} */,
  {32'hbf86b1a8, 32'h3f2a5990} /* (20, 26, 1) {real, imag} */,
  {32'hbf60d0a8, 32'h3e27f3c8} /* (20, 26, 0) {real, imag} */,
  {32'h3e2a8e48, 32'h3ecf4ab0} /* (20, 25, 31) {real, imag} */,
  {32'h3e906320, 32'h3fadc49a} /* (20, 25, 30) {real, imag} */,
  {32'hbda66600, 32'hbe4f7788} /* (20, 25, 29) {real, imag} */,
  {32'hbe0d8d40, 32'h3f2367de} /* (20, 25, 28) {real, imag} */,
  {32'hbe33423a, 32'h3f7e4dc4} /* (20, 25, 27) {real, imag} */,
  {32'hbdb302d0, 32'h3ef7a010} /* (20, 25, 26) {real, imag} */,
  {32'h3e268838, 32'h3e6d3ea0} /* (20, 25, 25) {real, imag} */,
  {32'hbeefc5c4, 32'h3e87b490} /* (20, 25, 24) {real, imag} */,
  {32'hbe373e68, 32'hbf79fa3c} /* (20, 25, 23) {real, imag} */,
  {32'hbf1f0aa6, 32'hbf87a1b4} /* (20, 25, 22) {real, imag} */,
  {32'hbf8485c8, 32'h3f008ede} /* (20, 25, 21) {real, imag} */,
  {32'hbec431f0, 32'hbf203170} /* (20, 25, 20) {real, imag} */,
  {32'h3f653f87, 32'hbfa4f928} /* (20, 25, 19) {real, imag} */,
  {32'h3f69c3e2, 32'hbe7512d0} /* (20, 25, 18) {real, imag} */,
  {32'h40004fe8, 32'hbe8f317c} /* (20, 25, 17) {real, imag} */,
  {32'h3fcce1e9, 32'hbd92da20} /* (20, 25, 16) {real, imag} */,
  {32'h3e93cabe, 32'h3d37f040} /* (20, 25, 15) {real, imag} */,
  {32'hbf3a8794, 32'hbe27b2a0} /* (20, 25, 14) {real, imag} */,
  {32'hbf3b1a83, 32'h3e37d640} /* (20, 25, 13) {real, imag} */,
  {32'h3d95dc14, 32'hbf77dad8} /* (20, 25, 12) {real, imag} */,
  {32'h3cca9eac, 32'hbefdaf28} /* (20, 25, 11) {real, imag} */,
  {32'h3e5cabcc, 32'h3d99cbe8} /* (20, 25, 10) {real, imag} */,
  {32'hbf4096dc, 32'hbf955dd5} /* (20, 25, 9) {real, imag} */,
  {32'hbed57248, 32'hbfd3eb34} /* (20, 25, 8) {real, imag} */,
  {32'h3f3e44fb, 32'h3da32e60} /* (20, 25, 7) {real, imag} */,
  {32'h3f6395de, 32'h3e9b60f4} /* (20, 25, 6) {real, imag} */,
  {32'h3d4b79e0, 32'h3e894af0} /* (20, 25, 5) {real, imag} */,
  {32'h3c89a640, 32'h3e9eb818} /* (20, 25, 4) {real, imag} */,
  {32'hbf5a3933, 32'h3fc000c6} /* (20, 25, 3) {real, imag} */,
  {32'hbfb46da6, 32'h3fb7580f} /* (20, 25, 2) {real, imag} */,
  {32'hbfc6832e, 32'hbeb7c2a8} /* (20, 25, 1) {real, imag} */,
  {32'hbf8eac30, 32'hbf38a7b6} /* (20, 25, 0) {real, imag} */,
  {32'h3e8529af, 32'h3f0df180} /* (20, 24, 31) {real, imag} */,
  {32'h3e57e21c, 32'h3e178dd0} /* (20, 24, 30) {real, imag} */,
  {32'h3e96072c, 32'hbed06ea0} /* (20, 24, 29) {real, imag} */,
  {32'h3f6e1f51, 32'hbd9bbd60} /* (20, 24, 28) {real, imag} */,
  {32'h3f686687, 32'hbdb213d0} /* (20, 24, 27) {real, imag} */,
  {32'h3f3eb7ee, 32'hbe6a3260} /* (20, 24, 26) {real, imag} */,
  {32'h3efa89b8, 32'hbfecac96} /* (20, 24, 25) {real, imag} */,
  {32'hbf1f000c, 32'hbfa17840} /* (20, 24, 24) {real, imag} */,
  {32'hbfb090c6, 32'hbf499120} /* (20, 24, 23) {real, imag} */,
  {32'hbf382329, 32'hbf3f8e10} /* (20, 24, 22) {real, imag} */,
  {32'hbebb4af5, 32'hbd3aac00} /* (20, 24, 21) {real, imag} */,
  {32'hbfc3ef16, 32'hbf110b18} /* (20, 24, 20) {real, imag} */,
  {32'hbfb8e2bc, 32'hbf9cce8f} /* (20, 24, 19) {real, imag} */,
  {32'hbf9e6281, 32'hbb77e800} /* (20, 24, 18) {real, imag} */,
  {32'hbeb70cb4, 32'h3c4edd00} /* (20, 24, 17) {real, imag} */,
  {32'h3f8fe5be, 32'hbe0d8ec0} /* (20, 24, 16) {real, imag} */,
  {32'h3ea83a93, 32'h3f11ad6c} /* (20, 24, 15) {real, imag} */,
  {32'h3cf6b5c0, 32'h3f9a6406} /* (20, 24, 14) {real, imag} */,
  {32'hbea83890, 32'h3f969066} /* (20, 24, 13) {real, imag} */,
  {32'h3f49c5da, 32'h3f224c98} /* (20, 24, 12) {real, imag} */,
  {32'h40107bce, 32'hbd6cf710} /* (20, 24, 11) {real, imag} */,
  {32'h3fdb79fe, 32'hbea3b01c} /* (20, 24, 10) {real, imag} */,
  {32'h3e37bec0, 32'hbf6084e0} /* (20, 24, 9) {real, imag} */,
  {32'h3d972520, 32'hbfba9d29} /* (20, 24, 8) {real, imag} */,
  {32'h3f6471ae, 32'hbe81df14} /* (20, 24, 7) {real, imag} */,
  {32'h3faf8e0a, 32'hbde6ac30} /* (20, 24, 6) {real, imag} */,
  {32'hbf236253, 32'h3f8f6c48} /* (20, 24, 5) {real, imag} */,
  {32'h3e0e7484, 32'h3fde2711} /* (20, 24, 4) {real, imag} */,
  {32'h3d0ec140, 32'h3fce16a0} /* (20, 24, 3) {real, imag} */,
  {32'hbf56db44, 32'h3f85eac4} /* (20, 24, 2) {real, imag} */,
  {32'h3da28898, 32'h3ea19b00} /* (20, 24, 1) {real, imag} */,
  {32'h3da0bab4, 32'hbea26c58} /* (20, 24, 0) {real, imag} */,
  {32'h3f11ad72, 32'h3f673700} /* (20, 23, 31) {real, imag} */,
  {32'hbe84cc84, 32'h3e45fa80} /* (20, 23, 30) {real, imag} */,
  {32'hbebff398, 32'hbeaaf910} /* (20, 23, 29) {real, imag} */,
  {32'h3f25d0f9, 32'hbee24ec8} /* (20, 23, 28) {real, imag} */,
  {32'hbd8282b0, 32'hbf2112dc} /* (20, 23, 27) {real, imag} */,
  {32'hbeb5ac48, 32'hbf9a0946} /* (20, 23, 26) {real, imag} */,
  {32'h3f7f53ba, 32'hbfc7a21e} /* (20, 23, 25) {real, imag} */,
  {32'hbeb56e9d, 32'hbe3b11f0} /* (20, 23, 24) {real, imag} */,
  {32'hc011b652, 32'h3ee85600} /* (20, 23, 23) {real, imag} */,
  {32'hbffdfe72, 32'h3d2f1580} /* (20, 23, 22) {real, imag} */,
  {32'hbf6d9608, 32'h3e158588} /* (20, 23, 21) {real, imag} */,
  {32'hbfd753fe, 32'h3e9091c4} /* (20, 23, 20) {real, imag} */,
  {32'hbfed72d0, 32'hbd3bd7e0} /* (20, 23, 19) {real, imag} */,
  {32'hbfa06754, 32'h3d9a37d0} /* (20, 23, 18) {real, imag} */,
  {32'hbfa98db2, 32'hbfb1dc59} /* (20, 23, 17) {real, imag} */,
  {32'h3ea2dc0e, 32'hbf99b920} /* (20, 23, 16) {real, imag} */,
  {32'h3d9851d0, 32'hbeeeae80} /* (20, 23, 15) {real, imag} */,
  {32'hbdcf0730, 32'h3e50ebe0} /* (20, 23, 14) {real, imag} */,
  {32'hbe7cde98, 32'h3f8390c4} /* (20, 23, 13) {real, imag} */,
  {32'h3f227e25, 32'h3fc62b5b} /* (20, 23, 12) {real, imag} */,
  {32'h3f9501c2, 32'h3f9a1c19} /* (20, 23, 11) {real, imag} */,
  {32'h3f93d5e2, 32'h3f518d93} /* (20, 23, 10) {real, imag} */,
  {32'h3f6d33ae, 32'h3e857eb0} /* (20, 23, 9) {real, imag} */,
  {32'h3f856dea, 32'hbea272a0} /* (20, 23, 8) {real, imag} */,
  {32'h3f5a81ff, 32'hbf9f7f6c} /* (20, 23, 7) {real, imag} */,
  {32'h3f1004da, 32'hbfb94d47} /* (20, 23, 6) {real, imag} */,
  {32'hbf52d75b, 32'hbedfbc70} /* (20, 23, 5) {real, imag} */,
  {32'h3eb5c8ec, 32'h3f1f937c} /* (20, 23, 4) {real, imag} */,
  {32'h3ef74b3c, 32'hbbc24b00} /* (20, 23, 3) {real, imag} */,
  {32'hbf2acfcc, 32'hbd1ca240} /* (20, 23, 2) {real, imag} */,
  {32'h3df40920, 32'h3f58c9c4} /* (20, 23, 1) {real, imag} */,
  {32'h3f13a59a, 32'h3fa6feda} /* (20, 23, 0) {real, imag} */,
  {32'hbc960740, 32'hbe2e5e10} /* (20, 22, 31) {real, imag} */,
  {32'hbf9ad9c8, 32'hbeac7450} /* (20, 22, 30) {real, imag} */,
  {32'hbf9f02f6, 32'h3edb0638} /* (20, 22, 29) {real, imag} */,
  {32'hbf3a463a, 32'hbea42518} /* (20, 22, 28) {real, imag} */,
  {32'hbf9b6696, 32'hbef19170} /* (20, 22, 27) {real, imag} */,
  {32'hbf31320a, 32'hbf816cb4} /* (20, 22, 26) {real, imag} */,
  {32'h3ebdd398, 32'hbf63bce8} /* (20, 22, 25) {real, imag} */,
  {32'hbe567d23, 32'h3eb61050} /* (20, 22, 24) {real, imag} */,
  {32'hbff6db2f, 32'h3f4ea100} /* (20, 22, 23) {real, imag} */,
  {32'hbff6481e, 32'h3eced280} /* (20, 22, 22) {real, imag} */,
  {32'hbedbd6f8, 32'h3f2aa010} /* (20, 22, 21) {real, imag} */,
  {32'hbf41440e, 32'h3f338706} /* (20, 22, 20) {real, imag} */,
  {32'hbf604d58, 32'hbe65d4dc} /* (20, 22, 19) {real, imag} */,
  {32'hbf87ab9c, 32'hbfd2d622} /* (20, 22, 18) {real, imag} */,
  {32'hbf3fb003, 32'hbfad27e0} /* (20, 22, 17) {real, imag} */,
  {32'h3f39c7e6, 32'hbf90a1f6} /* (20, 22, 16) {real, imag} */,
  {32'hbdd2aab0, 32'hbf8ba12a} /* (20, 22, 15) {real, imag} */,
  {32'hbecbb15c, 32'h3e24b130} /* (20, 22, 14) {real, imag} */,
  {32'h3ed996d0, 32'h3f90334c} /* (20, 22, 13) {real, imag} */,
  {32'h3e95eb34, 32'h3f4f97c0} /* (20, 22, 12) {real, imag} */,
  {32'hbd9196b0, 32'h3f89b9f4} /* (20, 22, 11) {real, imag} */,
  {32'h3f0f7f22, 32'h3f547327} /* (20, 22, 10) {real, imag} */,
  {32'h3db2d1b8, 32'hbdc5dca0} /* (20, 22, 9) {real, imag} */,
  {32'hbed7168c, 32'h3ecce910} /* (20, 22, 8) {real, imag} */,
  {32'h3e4b90c0, 32'hbf8330f4} /* (20, 22, 7) {real, imag} */,
  {32'h3ea126ac, 32'hbf3edeac} /* (20, 22, 6) {real, imag} */,
  {32'h3dd729a4, 32'hbeca58c8} /* (20, 22, 5) {real, imag} */,
  {32'hbf15ca1c, 32'h3df291c0} /* (20, 22, 4) {real, imag} */,
  {32'hbf00c2bc, 32'h3a333400} /* (20, 22, 3) {real, imag} */,
  {32'hbfba8a16, 32'hbf668c9c} /* (20, 22, 2) {real, imag} */,
  {32'hbebd9261, 32'h3f2014b2} /* (20, 22, 1) {real, imag} */,
  {32'h3e8085e4, 32'h3f879822} /* (20, 22, 0) {real, imag} */,
  {32'h3efa261e, 32'hbe1b2528} /* (20, 21, 31) {real, imag} */,
  {32'h3e512e18, 32'hbf4896f6} /* (20, 21, 30) {real, imag} */,
  {32'h3eab043c, 32'h3ebbe212} /* (20, 21, 29) {real, imag} */,
  {32'hbe8b675c, 32'h3f023dfc} /* (20, 21, 28) {real, imag} */,
  {32'hbf331a7f, 32'h3ef08e70} /* (20, 21, 27) {real, imag} */,
  {32'hbf5c74a4, 32'h3ea0cd14} /* (20, 21, 26) {real, imag} */,
  {32'hbf8fe2e0, 32'h3f4bd2c9} /* (20, 21, 25) {real, imag} */,
  {32'hbe971bf0, 32'h3d22fcc0} /* (20, 21, 24) {real, imag} */,
  {32'hbf26f337, 32'hbf396f5a} /* (20, 21, 23) {real, imag} */,
  {32'hbf0127c0, 32'hbe1f5fe8} /* (20, 21, 22) {real, imag} */,
  {32'hbf30ef62, 32'h3ec70b70} /* (20, 21, 21) {real, imag} */,
  {32'hbdf003b2, 32'h3c96dd10} /* (20, 21, 20) {real, imag} */,
  {32'hbe0b02ec, 32'hbf0b0738} /* (20, 21, 19) {real, imag} */,
  {32'hbf4c6b80, 32'hbfa3ee51} /* (20, 21, 18) {real, imag} */,
  {32'hbf186cae, 32'h3cd52480} /* (20, 21, 17) {real, imag} */,
  {32'h3e99019e, 32'hbf0380cc} /* (20, 21, 16) {real, imag} */,
  {32'hbf02049c, 32'hbddcbd60} /* (20, 21, 15) {real, imag} */,
  {32'hbf89c946, 32'h3f3dbbea} /* (20, 21, 14) {real, imag} */,
  {32'hbdbf99b8, 32'h3f54dce7} /* (20, 21, 13) {real, imag} */,
  {32'h3ea8e692, 32'h3f82642c} /* (20, 21, 12) {real, imag} */,
  {32'hbe8353c5, 32'h3f2d6ce0} /* (20, 21, 11) {real, imag} */,
  {32'hbdef36c8, 32'hbebcd224} /* (20, 21, 10) {real, imag} */,
  {32'h3f4bcf4c, 32'hbfa4efce} /* (20, 21, 9) {real, imag} */,
  {32'h3eec3056, 32'hbe2ccb60} /* (20, 21, 8) {real, imag} */,
  {32'h3f141922, 32'hbee98b74} /* (20, 21, 7) {real, imag} */,
  {32'hbe0819f2, 32'h3f3141df} /* (20, 21, 6) {real, imag} */,
  {32'h3c1a6dc0, 32'h3f250e89} /* (20, 21, 5) {real, imag} */,
  {32'hbea10166, 32'h3f2d0c97} /* (20, 21, 4) {real, imag} */,
  {32'hbe8b1c4a, 32'h3f747fed} /* (20, 21, 3) {real, imag} */,
  {32'hbf2b0b50, 32'h3f2d9f5b} /* (20, 21, 2) {real, imag} */,
  {32'h3e8606f6, 32'h3faf05b8} /* (20, 21, 1) {real, imag} */,
  {32'h3f1c8ea8, 32'h3f2f7f42} /* (20, 21, 0) {real, imag} */,
  {32'hbe8bb0fb, 32'h3eb692be} /* (20, 20, 31) {real, imag} */,
  {32'hbed1cada, 32'hbdb0ebac} /* (20, 20, 30) {real, imag} */,
  {32'hbd727a10, 32'h3e54c470} /* (20, 20, 29) {real, imag} */,
  {32'hbf49f623, 32'h3dee1ae0} /* (20, 20, 28) {real, imag} */,
  {32'hbf03d9b8, 32'h3f91f829} /* (20, 20, 27) {real, imag} */,
  {32'hbe412730, 32'h3f1f9a9c} /* (20, 20, 26) {real, imag} */,
  {32'hbe0f0b48, 32'hbd4eb780} /* (20, 20, 25) {real, imag} */,
  {32'h3fa340b4, 32'hbeae7cb0} /* (20, 20, 24) {real, imag} */,
  {32'h3fa64d42, 32'h3e05afb0} /* (20, 20, 23) {real, imag} */,
  {32'h3f01ed26, 32'h3ea990e0} /* (20, 20, 22) {real, imag} */,
  {32'hbf5a8329, 32'h3e854730} /* (20, 20, 21) {real, imag} */,
  {32'hbf991c67, 32'hbdc72cd0} /* (20, 20, 20) {real, imag} */,
  {32'hbe7d3c00, 32'hbf5e0da4} /* (20, 20, 19) {real, imag} */,
  {32'h3f460d4c, 32'hbe84faf4} /* (20, 20, 18) {real, imag} */,
  {32'h3f12a719, 32'h3fd3dbf8} /* (20, 20, 17) {real, imag} */,
  {32'h3f8bb36a, 32'h3f2b6fdf} /* (20, 20, 16) {real, imag} */,
  {32'h3e822b74, 32'hbe13a6c0} /* (20, 20, 15) {real, imag} */,
  {32'hbf02b46a, 32'h3ea08688} /* (20, 20, 14) {real, imag} */,
  {32'hbf829ced, 32'h3e99df48} /* (20, 20, 13) {real, imag} */,
  {32'hbf956996, 32'hbd960420} /* (20, 20, 12) {real, imag} */,
  {32'hbf950749, 32'h3efb7a58} /* (20, 20, 11) {real, imag} */,
  {32'hbf2b0ff3, 32'hbe12d7e9} /* (20, 20, 10) {real, imag} */,
  {32'h3f624818, 32'hbfae6023} /* (20, 20, 9) {real, imag} */,
  {32'h3f306b92, 32'hbfa58ad6} /* (20, 20, 8) {real, imag} */,
  {32'h3ec2de59, 32'hbf2d32c0} /* (20, 20, 7) {real, imag} */,
  {32'hbe33c83c, 32'h3f656298} /* (20, 20, 6) {real, imag} */,
  {32'h3ebca397, 32'h3fa8661c} /* (20, 20, 5) {real, imag} */,
  {32'h3f138bf8, 32'h3e92398c} /* (20, 20, 4) {real, imag} */,
  {32'h3ed6b075, 32'h3f07ce0c} /* (20, 20, 3) {real, imag} */,
  {32'h3e8f5c48, 32'h3f2d0090} /* (20, 20, 2) {real, imag} */,
  {32'h3f11dee1, 32'h3f41f364} /* (20, 20, 1) {real, imag} */,
  {32'h3f0486a7, 32'h3f39541e} /* (20, 20, 0) {real, imag} */,
  {32'hbef1887c, 32'h3d67cee0} /* (20, 19, 31) {real, imag} */,
  {32'hbeba53b8, 32'hbf211785} /* (20, 19, 30) {real, imag} */,
  {32'hbf8f1a84, 32'h3da7edf0} /* (20, 19, 29) {real, imag} */,
  {32'hbedf965e, 32'h3e8fe3e0} /* (20, 19, 28) {real, imag} */,
  {32'h3e80630b, 32'h3f7a8acc} /* (20, 19, 27) {real, imag} */,
  {32'h3f895b0e, 32'hbe1c83d0} /* (20, 19, 26) {real, imag} */,
  {32'h3f17d8d9, 32'hbe86cf78} /* (20, 19, 25) {real, imag} */,
  {32'h3f54a47c, 32'hbfa3f842} /* (20, 19, 24) {real, imag} */,
  {32'h3f064908, 32'h3e3d9fa0} /* (20, 19, 23) {real, imag} */,
  {32'h3edbf1b8, 32'h3f226e38} /* (20, 19, 22) {real, imag} */,
  {32'h3ebdcf14, 32'h3ed43168} /* (20, 19, 21) {real, imag} */,
  {32'hbe9c6a49, 32'h3f2a7528} /* (20, 19, 20) {real, imag} */,
  {32'hbe6cbc44, 32'hbe013a70} /* (20, 19, 19) {real, imag} */,
  {32'h3dd9a958, 32'h3eef6190} /* (20, 19, 18) {real, imag} */,
  {32'h3f0e5b8a, 32'h3f757c68} /* (20, 19, 17) {real, imag} */,
  {32'hbe7b4f80, 32'hbef9c30b} /* (20, 19, 16) {real, imag} */,
  {32'hbf102058, 32'hbef8d2b0} /* (20, 19, 15) {real, imag} */,
  {32'hbef18b34, 32'hbe293f30} /* (20, 19, 14) {real, imag} */,
  {32'hbf293914, 32'h3c47f600} /* (20, 19, 13) {real, imag} */,
  {32'hbf86cdac, 32'hbf8c8d36} /* (20, 19, 12) {real, imag} */,
  {32'hbed79bc6, 32'hbef678b0} /* (20, 19, 11) {real, imag} */,
  {32'h3fa17b04, 32'h3d581e20} /* (20, 19, 10) {real, imag} */,
  {32'h3f936ec0, 32'hbe624730} /* (20, 19, 9) {real, imag} */,
  {32'h3ea4a4c9, 32'hbe4ba960} /* (20, 19, 8) {real, imag} */,
  {32'hbc5f4980, 32'hbec0d5d0} /* (20, 19, 7) {real, imag} */,
  {32'h3efe8bb0, 32'hbf1dcc86} /* (20, 19, 6) {real, imag} */,
  {32'h3f67f2ac, 32'h3eae6d80} /* (20, 19, 5) {real, imag} */,
  {32'h3eb8c1fc, 32'h3f95f2f5} /* (20, 19, 4) {real, imag} */,
  {32'hbf3f1de2, 32'h3f745158} /* (20, 19, 3) {real, imag} */,
  {32'h3e025fa0, 32'h3dff1160} /* (20, 19, 2) {real, imag} */,
  {32'h3f92611c, 32'h3f07cee0} /* (20, 19, 1) {real, imag} */,
  {32'h3ea7114c, 32'h3fce2c5c} /* (20, 19, 0) {real, imag} */,
  {32'h3df72a28, 32'hbf11d844} /* (20, 18, 31) {real, imag} */,
  {32'hbe8290b4, 32'hbf2500d2} /* (20, 18, 30) {real, imag} */,
  {32'hbea96ef4, 32'hbf8a8c64} /* (20, 18, 29) {real, imag} */,
  {32'h3e006368, 32'hbe184d64} /* (20, 18, 28) {real, imag} */,
  {32'hbe523bf8, 32'h3f051960} /* (20, 18, 27) {real, imag} */,
  {32'h3f7453bc, 32'h3e462180} /* (20, 18, 26) {real, imag} */,
  {32'h3fa5e158, 32'h3dcaeac0} /* (20, 18, 25) {real, imag} */,
  {32'h3f104568, 32'h3e9c4658} /* (20, 18, 24) {real, imag} */,
  {32'hbf38847a, 32'h3f32ddac} /* (20, 18, 23) {real, imag} */,
  {32'hbcc0de80, 32'h3f6d5214} /* (20, 18, 22) {real, imag} */,
  {32'h3f9dd9c5, 32'h3f37a7a7} /* (20, 18, 21) {real, imag} */,
  {32'h3e3c6824, 32'h3f79573c} /* (20, 18, 20) {real, imag} */,
  {32'h3ef207c6, 32'h3f982712} /* (20, 18, 19) {real, imag} */,
  {32'hbfd34804, 32'h3f07ba60} /* (20, 18, 18) {real, imag} */,
  {32'hc0051faa, 32'h3b79e400} /* (20, 18, 17) {real, imag} */,
  {32'hbf569918, 32'hbe97ba4c} /* (20, 18, 16) {real, imag} */,
  {32'hbef508ca, 32'hbf5f60be} /* (20, 18, 15) {real, imag} */,
  {32'hbf4281bc, 32'hbf050c7a} /* (20, 18, 14) {real, imag} */,
  {32'hbf9793e1, 32'h3f2c558c} /* (20, 18, 13) {real, imag} */,
  {32'hbfbea8d2, 32'hbe93d6c8} /* (20, 18, 12) {real, imag} */,
  {32'hbf603970, 32'hbf7a2ba2} /* (20, 18, 11) {real, imag} */,
  {32'h3e810032, 32'h3e668b98} /* (20, 18, 10) {real, imag} */,
  {32'h3f4a9ed9, 32'h3fb018a4} /* (20, 18, 9) {real, imag} */,
  {32'h3d9e08e5, 32'h3fb99e52} /* (20, 18, 8) {real, imag} */,
  {32'hbe3a3184, 32'h3f47943c} /* (20, 18, 7) {real, imag} */,
  {32'hbee47fe4, 32'hbdf2aff0} /* (20, 18, 6) {real, imag} */,
  {32'hbea89d88, 32'hbec05190} /* (20, 18, 5) {real, imag} */,
  {32'hbeeb0f38, 32'h3f24b908} /* (20, 18, 4) {real, imag} */,
  {32'hbf6ab60d, 32'h3fa60ae9} /* (20, 18, 3) {real, imag} */,
  {32'hbf30fea0, 32'h3fa8dc20} /* (20, 18, 2) {real, imag} */,
  {32'h3eb13c78, 32'h3d481900} /* (20, 18, 1) {real, imag} */,
  {32'h3e0f5de8, 32'h3f8d071b} /* (20, 18, 0) {real, imag} */,
  {32'h3b9cdc00, 32'hbe471030} /* (20, 17, 31) {real, imag} */,
  {32'hbf2346d6, 32'hbdaa8c20} /* (20, 17, 30) {real, imag} */,
  {32'hbef254c4, 32'hbec6e9f0} /* (20, 17, 29) {real, imag} */,
  {32'h3e723cc0, 32'h3dc64940} /* (20, 17, 28) {real, imag} */,
  {32'h3f31c8f8, 32'h3f4fc030} /* (20, 17, 27) {real, imag} */,
  {32'h3f6f3eda, 32'h3f94f400} /* (20, 17, 26) {real, imag} */,
  {32'h3fbd26e0, 32'h3f720d1e} /* (20, 17, 25) {real, imag} */,
  {32'h3ed57774, 32'h3f65bdec} /* (20, 17, 24) {real, imag} */,
  {32'hbfa404e0, 32'h3f221740} /* (20, 17, 23) {real, imag} */,
  {32'hbe82b2e8, 32'h3fc10f20} /* (20, 17, 22) {real, imag} */,
  {32'h3f379850, 32'h3f512982} /* (20, 17, 21) {real, imag} */,
  {32'hbf4c547d, 32'h3fc14193} /* (20, 17, 20) {real, imag} */,
  {32'hbdfbd480, 32'h3f884a9a} /* (20, 17, 19) {real, imag} */,
  {32'hbfa17c9e, 32'h3e445ab0} /* (20, 17, 18) {real, imag} */,
  {32'hbfb24340, 32'h3f1bb950} /* (20, 17, 17) {real, imag} */,
  {32'h3dcafe14, 32'hbece4fe8} /* (20, 17, 16) {real, imag} */,
  {32'hbef83fe3, 32'hbf7a144e} /* (20, 17, 15) {real, imag} */,
  {32'hbf5a4d4c, 32'h3c79f100} /* (20, 17, 14) {real, imag} */,
  {32'hbf45ee72, 32'h3f8b9297} /* (20, 17, 13) {real, imag} */,
  {32'hbf7f467a, 32'h3bf50400} /* (20, 17, 12) {real, imag} */,
  {32'hbe985521, 32'hbea73abc} /* (20, 17, 11) {real, imag} */,
  {32'h3e8159c7, 32'h3f1d0e88} /* (20, 17, 10) {real, imag} */,
  {32'hbd5db060, 32'h3faadfdc} /* (20, 17, 9) {real, imag} */,
  {32'hbf88fc75, 32'h400cbbd0} /* (20, 17, 8) {real, imag} */,
  {32'hbf838e10, 32'h3f82bb00} /* (20, 17, 7) {real, imag} */,
  {32'hbfccd122, 32'hbdc4adc0} /* (20, 17, 6) {real, imag} */,
  {32'hbfa58280, 32'hbf422bbc} /* (20, 17, 5) {real, imag} */,
  {32'hbf2d6074, 32'hbe10a330} /* (20, 17, 4) {real, imag} */,
  {32'hbf9e539e, 32'hbdc52cd8} /* (20, 17, 3) {real, imag} */,
  {32'hbfb6bfc5, 32'hbd917a08} /* (20, 17, 2) {real, imag} */,
  {32'h3e412fd0, 32'hbeb28a7e} /* (20, 17, 1) {real, imag} */,
  {32'h3f973030, 32'h3e91e9ec} /* (20, 17, 0) {real, imag} */,
  {32'h3b72a700, 32'hbde2cbd0} /* (20, 16, 31) {real, imag} */,
  {32'hbd7acbd0, 32'hbee8a518} /* (20, 16, 30) {real, imag} */,
  {32'hbf29b98e, 32'hbf19fb8c} /* (20, 16, 29) {real, imag} */,
  {32'h3e40d340, 32'h3e339720} /* (20, 16, 28) {real, imag} */,
  {32'h3e969eb8, 32'h3f2aa064} /* (20, 16, 27) {real, imag} */,
  {32'h3f2ffa62, 32'h3ecdb980} /* (20, 16, 26) {real, imag} */,
  {32'h3f86781f, 32'h3f89ab3a} /* (20, 16, 25) {real, imag} */,
  {32'h3f6faff7, 32'hbf1d9814} /* (20, 16, 24) {real, imag} */,
  {32'hbde455e0, 32'hbf64870a} /* (20, 16, 23) {real, imag} */,
  {32'h3ea16f94, 32'h3f1d9b78} /* (20, 16, 22) {real, imag} */,
  {32'hbe08ead8, 32'h3e6f7d90} /* (20, 16, 21) {real, imag} */,
  {32'hbf8b7786, 32'h3f6c1f68} /* (20, 16, 20) {real, imag} */,
  {32'hbf1e6a18, 32'h3e0494e0} /* (20, 16, 19) {real, imag} */,
  {32'hbf0e135c, 32'hbf6a3b6e} /* (20, 16, 18) {real, imag} */,
  {32'hbe9d34f0, 32'hbeb74af8} /* (20, 16, 17) {real, imag} */,
  {32'hbda04780, 32'hbce7aa00} /* (20, 16, 16) {real, imag} */,
  {32'h3d6b3650, 32'h3f09b9fc} /* (20, 16, 15) {real, imag} */,
  {32'hbf3c9cea, 32'h3ee63528} /* (20, 16, 14) {real, imag} */,
  {32'hbeb55364, 32'hbf148834} /* (20, 16, 13) {real, imag} */,
  {32'hbe4ca970, 32'hbf5c9392} /* (20, 16, 12) {real, imag} */,
  {32'h3ee61858, 32'hbf99bc93} /* (20, 16, 11) {real, imag} */,
  {32'h3f0817b9, 32'hbf88e7fb} /* (20, 16, 10) {real, imag} */,
  {32'hbe50dc88, 32'h3f08ba7c} /* (20, 16, 9) {real, imag} */,
  {32'hbf66199c, 32'h3f01db6c} /* (20, 16, 8) {real, imag} */,
  {32'hbe8cfa9c, 32'h3df91740} /* (20, 16, 7) {real, imag} */,
  {32'hbeca3508, 32'h3f35c988} /* (20, 16, 6) {real, imag} */,
  {32'hbe9174b0, 32'hbf8b494b} /* (20, 16, 5) {real, imag} */,
  {32'hbf4feb2a, 32'hbfa82cb2} /* (20, 16, 4) {real, imag} */,
  {32'hbfe3a294, 32'hbfc448ee} /* (20, 16, 3) {real, imag} */,
  {32'hbfa69adf, 32'hbfad1e29} /* (20, 16, 2) {real, imag} */,
  {32'h3d37a290, 32'hbf3ec1ec} /* (20, 16, 1) {real, imag} */,
  {32'h3e10e0d4, 32'hbe9ede30} /* (20, 16, 0) {real, imag} */,
  {32'hbeedb1ac, 32'h3e2853bc} /* (20, 15, 31) {real, imag} */,
  {32'hbf9accbb, 32'hbd1af540} /* (20, 15, 30) {real, imag} */,
  {32'hc0004f74, 32'h3e8247a0} /* (20, 15, 29) {real, imag} */,
  {32'hbd0ae780, 32'hbd7764c0} /* (20, 15, 28) {real, imag} */,
  {32'h3f34168d, 32'hbe35a460} /* (20, 15, 27) {real, imag} */,
  {32'h3f71ed4c, 32'h3d2b6ae0} /* (20, 15, 26) {real, imag} */,
  {32'h3fb6c48e, 32'h3f10fbee} /* (20, 15, 25) {real, imag} */,
  {32'h3f61fb46, 32'hbef3a3d0} /* (20, 15, 24) {real, imag} */,
  {32'h3f2c2285, 32'hbf58e1e0} /* (20, 15, 23) {real, imag} */,
  {32'h3e64a349, 32'hbc95db80} /* (20, 15, 22) {real, imag} */,
  {32'hbf0176bd, 32'hbacb6000} /* (20, 15, 21) {real, imag} */,
  {32'h3e0241ec, 32'h3d1d41c0} /* (20, 15, 20) {real, imag} */,
  {32'hbdea9550, 32'hbe9ab3f0} /* (20, 15, 19) {real, imag} */,
  {32'hbdedd39c, 32'hbef07920} /* (20, 15, 18) {real, imag} */,
  {32'h3ed5aee8, 32'hbd0d1280} /* (20, 15, 17) {real, imag} */,
  {32'hbcc42080, 32'h3e826a98} /* (20, 15, 16) {real, imag} */,
  {32'hbeb8feda, 32'h3f736b60} /* (20, 15, 15) {real, imag} */,
  {32'hbf0f512a, 32'h3f4c828c} /* (20, 15, 14) {real, imag} */,
  {32'hbe85cc4e, 32'hbdc36c60} /* (20, 15, 13) {real, imag} */,
  {32'hbd145fc0, 32'hbf8a483f} /* (20, 15, 12) {real, imag} */,
  {32'h3ec762a5, 32'hbf6e01be} /* (20, 15, 11) {real, imag} */,
  {32'hbdf79000, 32'h3a1ff800} /* (20, 15, 10) {real, imag} */,
  {32'hbefdc188, 32'h3f8a4d6d} /* (20, 15, 9) {real, imag} */,
  {32'hbf7e4414, 32'h3e9fa768} /* (20, 15, 8) {real, imag} */,
  {32'hbf61e6ac, 32'hbda08c40} /* (20, 15, 7) {real, imag} */,
  {32'h3df133b0, 32'h3e7b43d0} /* (20, 15, 6) {real, imag} */,
  {32'h3ed16d0c, 32'hbdb95e80} /* (20, 15, 5) {real, imag} */,
  {32'hbea9e310, 32'hbd31d300} /* (20, 15, 4) {real, imag} */,
  {32'hbf6f637c, 32'hbf19d63c} /* (20, 15, 3) {real, imag} */,
  {32'hbeee966c, 32'hbecd5408} /* (20, 15, 2) {real, imag} */,
  {32'h3f06fce2, 32'hbeb3f520} /* (20, 15, 1) {real, imag} */,
  {32'hbd9aa9f8, 32'hbdf6a530} /* (20, 15, 0) {real, imag} */,
  {32'hbf05521f, 32'hbf1c0f5a} /* (20, 14, 31) {real, imag} */,
  {32'hbf84bc28, 32'hbf56a0a0} /* (20, 14, 30) {real, imag} */,
  {32'hbf83e0ae, 32'h3ec1bf08} /* (20, 14, 29) {real, imag} */,
  {32'hbe2a8140, 32'h3ee1ad50} /* (20, 14, 28) {real, imag} */,
  {32'h3f47a44f, 32'hbe814450} /* (20, 14, 27) {real, imag} */,
  {32'h3f896c2c, 32'h3e845f0c} /* (20, 14, 26) {real, imag} */,
  {32'h3f8ee150, 32'h3f988e36} /* (20, 14, 25) {real, imag} */,
  {32'h3f0057d8, 32'h3eabbfc4} /* (20, 14, 24) {real, imag} */,
  {32'h3f0b8aa2, 32'hbebafe60} /* (20, 14, 23) {real, imag} */,
  {32'h3cc75750, 32'hbd1a10c0} /* (20, 14, 22) {real, imag} */,
  {32'hbedf2550, 32'hbe3c8f80} /* (20, 14, 21) {real, imag} */,
  {32'hbf895496, 32'h3e6617c8} /* (20, 14, 20) {real, imag} */,
  {32'hbf15cf8c, 32'hbf9e7ef2} /* (20, 14, 19) {real, imag} */,
  {32'hbeca3f1c, 32'hbf6d91d0} /* (20, 14, 18) {real, imag} */,
  {32'hbee0ad17, 32'hbda7d4a0} /* (20, 14, 17) {real, imag} */,
  {32'hbf32406e, 32'hbea54b70} /* (20, 14, 16) {real, imag} */,
  {32'hbf1b4a7a, 32'h3c3cff00} /* (20, 14, 15) {real, imag} */,
  {32'h3e81573c, 32'h3fa6f88c} /* (20, 14, 14) {real, imag} */,
  {32'hbe479368, 32'h3f9bb455} /* (20, 14, 13) {real, imag} */,
  {32'h3ee30caa, 32'h3e2b5084} /* (20, 14, 12) {real, imag} */,
  {32'hbeb63430, 32'h3e294b1c} /* (20, 14, 11) {real, imag} */,
  {32'hbfa56863, 32'hbeb876d0} /* (20, 14, 10) {real, imag} */,
  {32'hbf880dc2, 32'hbc19f100} /* (20, 14, 9) {real, imag} */,
  {32'hbf3aa0b3, 32'hbdaa0880} /* (20, 14, 8) {real, imag} */,
  {32'hbf77fcfd, 32'hbed8f0f8} /* (20, 14, 7) {real, imag} */,
  {32'hbd535430, 32'hbcb51f00} /* (20, 14, 6) {real, imag} */,
  {32'h3f37a934, 32'h3ef78040} /* (20, 14, 5) {real, imag} */,
  {32'h3e5182b0, 32'h3ec81028} /* (20, 14, 4) {real, imag} */,
  {32'hbe091f30, 32'hbe4822c0} /* (20, 14, 3) {real, imag} */,
  {32'h39faf000, 32'hbe0d6170} /* (20, 14, 2) {real, imag} */,
  {32'h3e64a51c, 32'h3f028a10} /* (20, 14, 1) {real, imag} */,
  {32'hbe8eea86, 32'h3f678df6} /* (20, 14, 0) {real, imag} */,
  {32'hbdc34b10, 32'hbf2f2e32} /* (20, 13, 31) {real, imag} */,
  {32'h3ee281cc, 32'hbf3550a0} /* (20, 13, 30) {real, imag} */,
  {32'h3f3b5f00, 32'h3e0a8af0} /* (20, 13, 29) {real, imag} */,
  {32'h3ea57768, 32'hbecd93c0} /* (20, 13, 28) {real, imag} */,
  {32'hbe5e93f0, 32'hbf857950} /* (20, 13, 27) {real, imag} */,
  {32'h3ef63cec, 32'h3ec71fe8} /* (20, 13, 26) {real, imag} */,
  {32'h3f171bf6, 32'h3fb6ec7e} /* (20, 13, 25) {real, imag} */,
  {32'h3edf9470, 32'h3e865290} /* (20, 13, 24) {real, imag} */,
  {32'h3ee69c8c, 32'hbf1b3e44} /* (20, 13, 23) {real, imag} */,
  {32'hbef21a76, 32'h3c459100} /* (20, 13, 22) {real, imag} */,
  {32'hbfc8f42e, 32'h3e210bf0} /* (20, 13, 21) {real, imag} */,
  {32'hc0089c75, 32'h3f7bca12} /* (20, 13, 20) {real, imag} */,
  {32'hbf447382, 32'hbf91b82a} /* (20, 13, 19) {real, imag} */,
  {32'hbf9c73f7, 32'hbf0dc0f0} /* (20, 13, 18) {real, imag} */,
  {32'h3e3696a8, 32'h3ec0bdf0} /* (20, 13, 17) {real, imag} */,
  {32'h3f4c098e, 32'hbeb453b0} /* (20, 13, 16) {real, imag} */,
  {32'hbe7105bc, 32'h3e2bb930} /* (20, 13, 15) {real, imag} */,
  {32'hbf56aa88, 32'h3f982dc4} /* (20, 13, 14) {real, imag} */,
  {32'hbebc59fa, 32'h3fcf6ab4} /* (20, 13, 13) {real, imag} */,
  {32'h3f1a8e88, 32'h3ed255a8} /* (20, 13, 12) {real, imag} */,
  {32'hbc294a80, 32'hbe9d9dc8} /* (20, 13, 11) {real, imag} */,
  {32'hbf61a911, 32'hbf06f034} /* (20, 13, 10) {real, imag} */,
  {32'hbf32a6cd, 32'hbc0c8700} /* (20, 13, 9) {real, imag} */,
  {32'hbe87e198, 32'h3fa21a0e} /* (20, 13, 8) {real, imag} */,
  {32'hbdefdf20, 32'h3e8da008} /* (20, 13, 7) {real, imag} */,
  {32'hbe903bfc, 32'hbeb46d60} /* (20, 13, 6) {real, imag} */,
  {32'h3e1ddd28, 32'h3eef9f70} /* (20, 13, 5) {real, imag} */,
  {32'hbd9d5d30, 32'hbd4baac0} /* (20, 13, 4) {real, imag} */,
  {32'h3dc20a00, 32'hbe8fc520} /* (20, 13, 3) {real, imag} */,
  {32'h3dfb3680, 32'h3f7813e8} /* (20, 13, 2) {real, imag} */,
  {32'h3f519f9d, 32'h3f8538c8} /* (20, 13, 1) {real, imag} */,
  {32'hbbc241a0, 32'h3f1afbf7} /* (20, 13, 0) {real, imag} */,
  {32'hbd1164e0, 32'hbeb3553c} /* (20, 12, 31) {real, imag} */,
  {32'h3f605f76, 32'hbda5d4a0} /* (20, 12, 30) {real, imag} */,
  {32'h3f163772, 32'h3d238a80} /* (20, 12, 29) {real, imag} */,
  {32'hbe1c0be0, 32'hbe748680} /* (20, 12, 28) {real, imag} */,
  {32'h3ec86c94, 32'hbe6ecc70} /* (20, 12, 27) {real, imag} */,
  {32'h3f18399c, 32'h3eb6aef8} /* (20, 12, 26) {real, imag} */,
  {32'h3f260904, 32'h3f3af234} /* (20, 12, 25) {real, imag} */,
  {32'h3ebb79a0, 32'h3f7265f8} /* (20, 12, 24) {real, imag} */,
  {32'hbe645f90, 32'h3f1d3868} /* (20, 12, 23) {real, imag} */,
  {32'hbf4f8e24, 32'hbe1ad398} /* (20, 12, 22) {real, imag} */,
  {32'hbf17f93a, 32'hbe83d368} /* (20, 12, 21) {real, imag} */,
  {32'hbee15fba, 32'hbf3a4e36} /* (20, 12, 20) {real, imag} */,
  {32'h3de79500, 32'hbfc77e2a} /* (20, 12, 19) {real, imag} */,
  {32'hbf3ea5b8, 32'hbeb0bdb8} /* (20, 12, 18) {real, imag} */,
  {32'hbe883768, 32'h3eacdc78} /* (20, 12, 17) {real, imag} */,
  {32'h3b5a1800, 32'hbf35c12c} /* (20, 12, 16) {real, imag} */,
  {32'h3d6a4720, 32'hbd90f4e0} /* (20, 12, 15) {real, imag} */,
  {32'hbf69d1c8, 32'h3fcbf8b2} /* (20, 12, 14) {real, imag} */,
  {32'hbeb262a0, 32'h3fe6bb03} /* (20, 12, 13) {real, imag} */,
  {32'h3e869fec, 32'h3e830490} /* (20, 12, 12) {real, imag} */,
  {32'h3f3a619a, 32'hbf49d380} /* (20, 12, 11) {real, imag} */,
  {32'h3dc25c85, 32'h3e3e965b} /* (20, 12, 10) {real, imag} */,
  {32'hbee02d84, 32'h3f1a09c4} /* (20, 12, 9) {real, imag} */,
  {32'h3ec75844, 32'h3fb9c3dc} /* (20, 12, 8) {real, imag} */,
  {32'h3ed01c04, 32'h3f808cd4} /* (20, 12, 7) {real, imag} */,
  {32'h3f6bbfb0, 32'h3f0db7fc} /* (20, 12, 6) {real, imag} */,
  {32'h3f262052, 32'h3f5f5258} /* (20, 12, 5) {real, imag} */,
  {32'hbe34fe90, 32'hbf57459e} /* (20, 12, 4) {real, imag} */,
  {32'hbf196366, 32'hbefcdc68} /* (20, 12, 3) {real, imag} */,
  {32'hbf02f7f0, 32'h3ec6ddb8} /* (20, 12, 2) {real, imag} */,
  {32'h3f9b9b07, 32'h3f874cf2} /* (20, 12, 1) {real, imag} */,
  {32'h3f16c28b, 32'h3d76e000} /* (20, 12, 0) {real, imag} */,
  {32'h3c29b600, 32'hbec96b3c} /* (20, 11, 31) {real, imag} */,
  {32'h3f2a8ee8, 32'hbf4bbfa6} /* (20, 11, 30) {real, imag} */,
  {32'hbf11f24b, 32'hbf9ee1b6} /* (20, 11, 29) {real, imag} */,
  {32'hbfda9ab8, 32'hbf579e84} /* (20, 11, 28) {real, imag} */,
  {32'hbf34be19, 32'h3e9d6230} /* (20, 11, 27) {real, imag} */,
  {32'hbef87fac, 32'hbd8a8330} /* (20, 11, 26) {real, imag} */,
  {32'hbe976d8c, 32'hbfba526b} /* (20, 11, 25) {real, imag} */,
  {32'hbf1d68bc, 32'hbf5d6412} /* (20, 11, 24) {real, imag} */,
  {32'hbd2e8c60, 32'h3ef6ebb8} /* (20, 11, 23) {real, imag} */,
  {32'h3f76adb9, 32'hbf08c6ec} /* (20, 11, 22) {real, imag} */,
  {32'h3ed2bd98, 32'hbeb70c90} /* (20, 11, 21) {real, imag} */,
  {32'hbf18519a, 32'hbf652bfd} /* (20, 11, 20) {real, imag} */,
  {32'hbf706f18, 32'hbfc23874} /* (20, 11, 19) {real, imag} */,
  {32'h3e0a44c8, 32'hc00acbd5} /* (20, 11, 18) {real, imag} */,
  {32'h3e808d18, 32'hbf3c75d4} /* (20, 11, 17) {real, imag} */,
  {32'h3f1761f8, 32'hbdae7700} /* (20, 11, 16) {real, imag} */,
  {32'h3ee600fa, 32'hbe951348} /* (20, 11, 15) {real, imag} */,
  {32'hbf1385fb, 32'h3fb3367a} /* (20, 11, 14) {real, imag} */,
  {32'h3c8a4470, 32'h3f8575e3} /* (20, 11, 13) {real, imag} */,
  {32'h3fa4edd9, 32'hbf3054dc} /* (20, 11, 12) {real, imag} */,
  {32'h3f9136bc, 32'hbf6833e4} /* (20, 11, 11) {real, imag} */,
  {32'h3ef5de44, 32'hbd9a2450} /* (20, 11, 10) {real, imag} */,
  {32'hbe2553d8, 32'hbea8d210} /* (20, 11, 9) {real, imag} */,
  {32'h3f110a58, 32'h3eaf2e68} /* (20, 11, 8) {real, imag} */,
  {32'h3f5e03d6, 32'h3eefc0a0} /* (20, 11, 7) {real, imag} */,
  {32'h3f909546, 32'h3f1738a0} /* (20, 11, 6) {real, imag} */,
  {32'h3fa4f1e8, 32'h3f44d94c} /* (20, 11, 5) {real, imag} */,
  {32'h3f016566, 32'hbf6141d8} /* (20, 11, 4) {real, imag} */,
  {32'hbfa2a888, 32'h3ebcabf8} /* (20, 11, 3) {real, imag} */,
  {32'hbf521714, 32'h3edab7e0} /* (20, 11, 2) {real, imag} */,
  {32'h3e1328ee, 32'h3f154840} /* (20, 11, 1) {real, imag} */,
  {32'h3ec32df2, 32'h3edd9640} /* (20, 11, 0) {real, imag} */,
  {32'hbe9e19f0, 32'hbf4fdf78} /* (20, 10, 31) {real, imag} */,
  {32'h3d3c2a80, 32'hbfd713f0} /* (20, 10, 30) {real, imag} */,
  {32'h3f19f584, 32'hbf778aa0} /* (20, 10, 29) {real, imag} */,
  {32'hbcd69760, 32'hbf016b06} /* (20, 10, 28) {real, imag} */,
  {32'hbe783968, 32'h3e1fbc60} /* (20, 10, 27) {real, imag} */,
  {32'hbec15c48, 32'hbee3b638} /* (20, 10, 26) {real, imag} */,
  {32'hbf8d98c9, 32'hbf4d6ca2} /* (20, 10, 25) {real, imag} */,
  {32'hc0008426, 32'hbf731afa} /* (20, 10, 24) {real, imag} */,
  {32'hbd24e9eb, 32'h3f314ff8} /* (20, 10, 23) {real, imag} */,
  {32'h3d319170, 32'h3fb34b53} /* (20, 10, 22) {real, imag} */,
  {32'hbe50bf46, 32'h3f7b3b7a} /* (20, 10, 21) {real, imag} */,
  {32'h3e598e48, 32'hbd96dc20} /* (20, 10, 20) {real, imag} */,
  {32'hbb54d500, 32'hbe060513} /* (20, 10, 19) {real, imag} */,
  {32'h3e02c638, 32'hbf96e8f8} /* (20, 10, 18) {real, imag} */,
  {32'h3ee1ac3c, 32'hbf876f5b} /* (20, 10, 17) {real, imag} */,
  {32'h3fd882fd, 32'h3e625170} /* (20, 10, 16) {real, imag} */,
  {32'h40088bb0, 32'h3f2f0404} /* (20, 10, 15) {real, imag} */,
  {32'h3f8682bb, 32'h3e6b2244} /* (20, 10, 14) {real, imag} */,
  {32'h3e20e510, 32'hbf67ddca} /* (20, 10, 13) {real, imag} */,
  {32'h3f145e22, 32'h3d82c780} /* (20, 10, 12) {real, imag} */,
  {32'h3dcc18d8, 32'h3eb926c2} /* (20, 10, 11) {real, imag} */,
  {32'hbeac60df, 32'h3f39536f} /* (20, 10, 10) {real, imag} */,
  {32'hbf08c954, 32'hbd1a934e} /* (20, 10, 9) {real, imag} */,
  {32'h3e4633ca, 32'h3ed11ab8} /* (20, 10, 8) {real, imag} */,
  {32'h3f67f430, 32'h3f5dee05} /* (20, 10, 7) {real, imag} */,
  {32'h3f367234, 32'h3f5df5b2} /* (20, 10, 6) {real, imag} */,
  {32'hbef6ad92, 32'h3eb7651e} /* (20, 10, 5) {real, imag} */,
  {32'h3f0853da, 32'h3f05d9df} /* (20, 10, 4) {real, imag} */,
  {32'h3e83537a, 32'h3f2527bc} /* (20, 10, 3) {real, imag} */,
  {32'h3ee02ccc, 32'h3c51a400} /* (20, 10, 2) {real, imag} */,
  {32'h3e35b1c0, 32'h3f64c2b0} /* (20, 10, 1) {real, imag} */,
  {32'h3e1fd57c, 32'h3e04a418} /* (20, 10, 0) {real, imag} */,
  {32'hbf0568c5, 32'hbf5de200} /* (20, 9, 31) {real, imag} */,
  {32'hbebe4a14, 32'hbdadc2a0} /* (20, 9, 30) {real, imag} */,
  {32'h3f700afd, 32'h3f446089} /* (20, 9, 29) {real, imag} */,
  {32'h3f082f7b, 32'hbd191940} /* (20, 9, 28) {real, imag} */,
  {32'hbe18fa78, 32'h3f1e9388} /* (20, 9, 27) {real, imag} */,
  {32'hbecbb42c, 32'h3f014a3c} /* (20, 9, 26) {real, imag} */,
  {32'hbf767667, 32'h3f6a6d4c} /* (20, 9, 25) {real, imag} */,
  {32'hbfc056f4, 32'hbe0e1230} /* (20, 9, 24) {real, imag} */,
  {32'hbf5551a2, 32'h3e7b15a0} /* (20, 9, 23) {real, imag} */,
  {32'hbf652c7a, 32'h3f3ced58} /* (20, 9, 22) {real, imag} */,
  {32'hbea91f22, 32'h3f86838e} /* (20, 9, 21) {real, imag} */,
  {32'hbe82b8ae, 32'hbdce8300} /* (20, 9, 20) {real, imag} */,
  {32'hbe9fc69c, 32'h3e1b0240} /* (20, 9, 19) {real, imag} */,
  {32'h3f2a4ada, 32'h3e7790f8} /* (20, 9, 18) {real, imag} */,
  {32'h400fee29, 32'hbed579f0} /* (20, 9, 17) {real, imag} */,
  {32'h3fda1a18, 32'hbe494cf0} /* (20, 9, 16) {real, imag} */,
  {32'h3f412831, 32'h3f8271fe} /* (20, 9, 15) {real, imag} */,
  {32'hbed29af0, 32'h3f31f4b0} /* (20, 9, 14) {real, imag} */,
  {32'hbf6b1242, 32'hbe9a4f18} /* (20, 9, 13) {real, imag} */,
  {32'h3debc168, 32'h3f5f7e50} /* (20, 9, 12) {real, imag} */,
  {32'h3f4c6f3e, 32'h3eeffe88} /* (20, 9, 11) {real, imag} */,
  {32'h3e0db190, 32'h3ea3dd43} /* (20, 9, 10) {real, imag} */,
  {32'hbe711cc8, 32'hbe97bb90} /* (20, 9, 9) {real, imag} */,
  {32'h3ef47840, 32'h3ef23b18} /* (20, 9, 8) {real, imag} */,
  {32'h3f5310db, 32'h3e6b0898} /* (20, 9, 7) {real, imag} */,
  {32'hbee4e38e, 32'h3de93a70} /* (20, 9, 6) {real, imag} */,
  {32'hbe4c341c, 32'h3e06a0a0} /* (20, 9, 5) {real, imag} */,
  {32'hbc5be910, 32'hbec49da8} /* (20, 9, 4) {real, imag} */,
  {32'hbe2c8d18, 32'hbd30a080} /* (20, 9, 3) {real, imag} */,
  {32'h3e82365c, 32'h3e8946a0} /* (20, 9, 2) {real, imag} */,
  {32'hbc519e80, 32'hbf1ab7d4} /* (20, 9, 1) {real, imag} */,
  {32'h3f0c3d56, 32'hbf2e3b48} /* (20, 9, 0) {real, imag} */,
  {32'h3d000660, 32'h3e161540} /* (20, 8, 31) {real, imag} */,
  {32'hbe06aee5, 32'h3f4b51b0} /* (20, 8, 30) {real, imag} */,
  {32'h3e8dfee7, 32'h3fd91536} /* (20, 8, 29) {real, imag} */,
  {32'h3c6861d0, 32'h3fcdd4be} /* (20, 8, 28) {real, imag} */,
  {32'h3e172e9c, 32'h3f2bf742} /* (20, 8, 27) {real, imag} */,
  {32'hbdf2dce4, 32'h3f47fb7e} /* (20, 8, 26) {real, imag} */,
  {32'hbf127406, 32'h3fafd663} /* (20, 8, 25) {real, imag} */,
  {32'hbf870c94, 32'hbd5707a0} /* (20, 8, 24) {real, imag} */,
  {32'hbe9ac844, 32'hbf351ff4} /* (20, 8, 23) {real, imag} */,
  {32'h3e40731c, 32'h3f05065c} /* (20, 8, 22) {real, imag} */,
  {32'hbd746d20, 32'h3f06ae43} /* (20, 8, 21) {real, imag} */,
  {32'h3e6b1784, 32'h3d5b9780} /* (20, 8, 20) {real, imag} */,
  {32'hbd53cd86, 32'h3f1ef450} /* (20, 8, 19) {real, imag} */,
  {32'h3f92ed4c, 32'h3f361306} /* (20, 8, 18) {real, imag} */,
  {32'h3fdebd91, 32'hbea48b38} /* (20, 8, 17) {real, imag} */,
  {32'hbe8dfd58, 32'hbfb78730} /* (20, 8, 16) {real, imag} */,
  {32'hbf8502b9, 32'hbf08f98a} /* (20, 8, 15) {real, imag} */,
  {32'hbf6d4c0a, 32'h3f686b5c} /* (20, 8, 14) {real, imag} */,
  {32'hbf043dd6, 32'h3f1a12c0} /* (20, 8, 13) {real, imag} */,
  {32'h3ea83ecc, 32'h3f15d6c8} /* (20, 8, 12) {real, imag} */,
  {32'h3f35d12a, 32'h3e3c1960} /* (20, 8, 11) {real, imag} */,
  {32'hbf3ff211, 32'hbf46bbf0} /* (20, 8, 10) {real, imag} */,
  {32'hbeec2c0b, 32'hbf7e075e} /* (20, 8, 9) {real, imag} */,
  {32'h3f41b99d, 32'hbdc24878} /* (20, 8, 8) {real, imag} */,
  {32'hbeee83ca, 32'hbe124f88} /* (20, 8, 7) {real, imag} */,
  {32'hbf1f02db, 32'h3ea00304} /* (20, 8, 6) {real, imag} */,
  {32'h3f8ed522, 32'h3e3436a0} /* (20, 8, 5) {real, imag} */,
  {32'h3fced698, 32'hbfa55156} /* (20, 8, 4) {real, imag} */,
  {32'h3f6414e1, 32'h3e2f9440} /* (20, 8, 3) {real, imag} */,
  {32'h3eb97934, 32'hbee98080} /* (20, 8, 2) {real, imag} */,
  {32'hbecb2b90, 32'hbfae6ce8} /* (20, 8, 1) {real, imag} */,
  {32'h3d604450, 32'hbe60fd20} /* (20, 8, 0) {real, imag} */,
  {32'hbf818f55, 32'hbe7cc020} /* (20, 7, 31) {real, imag} */,
  {32'hbf5fb938, 32'hbf8db374} /* (20, 7, 30) {real, imag} */,
  {32'hbd06d940, 32'hbd8387a0} /* (20, 7, 29) {real, imag} */,
  {32'h3e3973a0, 32'h3f560338} /* (20, 7, 28) {real, imag} */,
  {32'h3f2282c8, 32'h3f4bafb4} /* (20, 7, 27) {real, imag} */,
  {32'h3eb2a5b4, 32'h3f78bc80} /* (20, 7, 26) {real, imag} */,
  {32'hbeff4f48, 32'h3fcf9faf} /* (20, 7, 25) {real, imag} */,
  {32'hbf750382, 32'h3f21f76c} /* (20, 7, 24) {real, imag} */,
  {32'h3f35b5fa, 32'hbf930628} /* (20, 7, 23) {real, imag} */,
  {32'h3ed55736, 32'hbf67d258} /* (20, 7, 22) {real, imag} */,
  {32'hbefc9b7b, 32'h3c25ed00} /* (20, 7, 21) {real, imag} */,
  {32'h3f1dae64, 32'h3d031900} /* (20, 7, 20) {real, imag} */,
  {32'hbea3cf18, 32'h3f0aecc4} /* (20, 7, 19) {real, imag} */,
  {32'hbf0f8323, 32'h3e9fb590} /* (20, 7, 18) {real, imag} */,
  {32'hbe384496, 32'hbdce8b60} /* (20, 7, 17) {real, imag} */,
  {32'hbf439124, 32'hbf56687e} /* (20, 7, 16) {real, imag} */,
  {32'hbf38588c, 32'hbf60fe58} /* (20, 7, 15) {real, imag} */,
  {32'hbe95ec7e, 32'h3eb05ab8} /* (20, 7, 14) {real, imag} */,
  {32'h3da53320, 32'h3e60b940} /* (20, 7, 13) {real, imag} */,
  {32'h3eea69c6, 32'h3e418b60} /* (20, 7, 12) {real, imag} */,
  {32'h3e9d8f93, 32'h3e7fc3f8} /* (20, 7, 11) {real, imag} */,
  {32'hbf88a9c8, 32'hbf32f628} /* (20, 7, 10) {real, imag} */,
  {32'hbee3a656, 32'hbe0947a0} /* (20, 7, 9) {real, imag} */,
  {32'h3e0c2974, 32'hbec76410} /* (20, 7, 8) {real, imag} */,
  {32'h3cc0e620, 32'hbe2d4b40} /* (20, 7, 7) {real, imag} */,
  {32'h3ac8ac00, 32'h3f975464} /* (20, 7, 6) {real, imag} */,
  {32'h3f292f6a, 32'h3f101e20} /* (20, 7, 5) {real, imag} */,
  {32'h3f29f22e, 32'hbf97f41c} /* (20, 7, 4) {real, imag} */,
  {32'h3f1365c5, 32'hbf245330} /* (20, 7, 3) {real, imag} */,
  {32'h3f446be0, 32'hbd3acd40} /* (20, 7, 2) {real, imag} */,
  {32'hbf0ddb12, 32'h3d083740} /* (20, 7, 1) {real, imag} */,
  {32'hbf39e755, 32'h3f0c804c} /* (20, 7, 0) {real, imag} */,
  {32'h3d3a9c90, 32'hbeecc3ec} /* (20, 6, 31) {real, imag} */,
  {32'h3ec6d9e0, 32'hbf6b4170} /* (20, 6, 30) {real, imag} */,
  {32'h3ec1dcca, 32'hbdc2dbc0} /* (20, 6, 29) {real, imag} */,
  {32'hbea9b6f0, 32'hbe642130} /* (20, 6, 28) {real, imag} */,
  {32'h3de89710, 32'h3f16091e} /* (20, 6, 27) {real, imag} */,
  {32'hbedf4f54, 32'h3e24b7f8} /* (20, 6, 26) {real, imag} */,
  {32'hbed24f20, 32'hbdfea120} /* (20, 6, 25) {real, imag} */,
  {32'hbf6ac8ee, 32'h3e722870} /* (20, 6, 24) {real, imag} */,
  {32'hbf8039f1, 32'h3c8ecd00} /* (20, 6, 23) {real, imag} */,
  {32'hbf862f64, 32'hbf65d304} /* (20, 6, 22) {real, imag} */,
  {32'hbec6c654, 32'hbf3e190a} /* (20, 6, 21) {real, imag} */,
  {32'h3f0d9caf, 32'h3efd2d58} /* (20, 6, 20) {real, imag} */,
  {32'h3ed30308, 32'hbe97a0d8} /* (20, 6, 19) {real, imag} */,
  {32'hbdff2a60, 32'hbf8b513d} /* (20, 6, 18) {real, imag} */,
  {32'hbe826946, 32'hbe75e910} /* (20, 6, 17) {real, imag} */,
  {32'hbf2c48cb, 32'h3ee19370} /* (20, 6, 16) {real, imag} */,
  {32'hbf1dbd7c, 32'hbe1ddd30} /* (20, 6, 15) {real, imag} */,
  {32'h3eaa3f34, 32'hbf63ec16} /* (20, 6, 14) {real, imag} */,
  {32'hbf0a0b64, 32'hbf5fa9be} /* (20, 6, 13) {real, imag} */,
  {32'hbfbf3f40, 32'hbf75c0c0} /* (20, 6, 12) {real, imag} */,
  {32'hbe7f05b8, 32'hbef2f398} /* (20, 6, 11) {real, imag} */,
  {32'h3f1d8c36, 32'hbf46e208} /* (20, 6, 10) {real, imag} */,
  {32'h3f436280, 32'hbe977320} /* (20, 6, 9) {real, imag} */,
  {32'hbe211170, 32'h3ed6d4c8} /* (20, 6, 8) {real, imag} */,
  {32'h3e05a3e0, 32'h3fbf028a} /* (20, 6, 7) {real, imag} */,
  {32'hbed73d62, 32'h3fa9dbda} /* (20, 6, 6) {real, imag} */,
  {32'hbf0918dd, 32'h3f137808} /* (20, 6, 5) {real, imag} */,
  {32'h3ea34e80, 32'hbefe3c88} /* (20, 6, 4) {real, imag} */,
  {32'hbf304eb6, 32'h3db62fe0} /* (20, 6, 3) {real, imag} */,
  {32'hbfb4887c, 32'h3f3066a4} /* (20, 6, 2) {real, imag} */,
  {32'hbfbeeddc, 32'h3eb58aa8} /* (20, 6, 1) {real, imag} */,
  {32'hbe92e4c0, 32'h3ee80b2d} /* (20, 6, 0) {real, imag} */,
  {32'h3e1d5188, 32'h3de58280} /* (20, 5, 31) {real, imag} */,
  {32'h3e312dd0, 32'hbf8dd0fe} /* (20, 5, 30) {real, imag} */,
  {32'h3e5d0160, 32'hbf356a24} /* (20, 5, 29) {real, imag} */,
  {32'hbfaf1a02, 32'hbf204204} /* (20, 5, 28) {real, imag} */,
  {32'hbe809ff0, 32'hbec9bd68} /* (20, 5, 27) {real, imag} */,
  {32'h3f0b85a1, 32'h3e9dd3b6} /* (20, 5, 26) {real, imag} */,
  {32'h3f764d7f, 32'h3ca55e00} /* (20, 5, 25) {real, imag} */,
  {32'hbedf504e, 32'hbba12200} /* (20, 5, 24) {real, imag} */,
  {32'hbf68ff3d, 32'h3f3044d0} /* (20, 5, 23) {real, imag} */,
  {32'h3f1631fc, 32'h3e579930} /* (20, 5, 22) {real, imag} */,
  {32'h3e3d59c0, 32'hbfb43912} /* (20, 5, 21) {real, imag} */,
  {32'h3ec2445e, 32'h3f0a7368} /* (20, 5, 20) {real, imag} */,
  {32'h3f7d2454, 32'h3eee5f7d} /* (20, 5, 19) {real, imag} */,
  {32'hbf176a76, 32'hbf0b926c} /* (20, 5, 18) {real, imag} */,
  {32'hbf2c83bd, 32'hbf5fe219} /* (20, 5, 17) {real, imag} */,
  {32'hbd67fad0, 32'h3e6069d7} /* (20, 5, 16) {real, imag} */,
  {32'h3ea26ada, 32'h3acb9c00} /* (20, 5, 15) {real, imag} */,
  {32'h3ee721d7, 32'hbf37e5e9} /* (20, 5, 14) {real, imag} */,
  {32'hbe00489e, 32'hbf001752} /* (20, 5, 13) {real, imag} */,
  {32'hbe5b1cf0, 32'h3b925000} /* (20, 5, 12) {real, imag} */,
  {32'h3e8c9034, 32'h3f093ed0} /* (20, 5, 11) {real, imag} */,
  {32'h4013aba2, 32'hbd88e3e0} /* (20, 5, 10) {real, imag} */,
  {32'h3f83c1c2, 32'hbf86b403} /* (20, 5, 9) {real, imag} */,
  {32'h3cb07660, 32'hbf0b5316} /* (20, 5, 8) {real, imag} */,
  {32'hbe7d4af4, 32'h3f913c50} /* (20, 5, 7) {real, imag} */,
  {32'hbfa8f162, 32'h3fc1e55f} /* (20, 5, 6) {real, imag} */,
  {32'hbe4c3454, 32'hbee794d8} /* (20, 5, 5) {real, imag} */,
  {32'h3e5dbd30, 32'hbf2a4f88} /* (20, 5, 4) {real, imag} */,
  {32'hbf313bb4, 32'h3f7248a0} /* (20, 5, 3) {real, imag} */,
  {32'hbfabc56f, 32'hbc8edb00} /* (20, 5, 2) {real, imag} */,
  {32'hbefe25ee, 32'hbf3d4fca} /* (20, 5, 1) {real, imag} */,
  {32'h3ec76440, 32'h3f182672} /* (20, 5, 0) {real, imag} */,
  {32'hbf21a6cd, 32'h3e5e4fc0} /* (20, 4, 31) {real, imag} */,
  {32'hbf4291b2, 32'h397dc000} /* (20, 4, 30) {real, imag} */,
  {32'hbe6d4a20, 32'hbd9a69c0} /* (20, 4, 29) {real, imag} */,
  {32'hbec355af, 32'hbf20c3c4} /* (20, 4, 28) {real, imag} */,
  {32'hbee9c816, 32'hbf8372e0} /* (20, 4, 27) {real, imag} */,
  {32'hbeccd9f8, 32'h3e1fc8b0} /* (20, 4, 26) {real, imag} */,
  {32'h3fa49f7a, 32'h3f3b1574} /* (20, 4, 25) {real, imag} */,
  {32'h3f62fa42, 32'h3f3021d2} /* (20, 4, 24) {real, imag} */,
  {32'h3f219e77, 32'h3eddd778} /* (20, 4, 23) {real, imag} */,
  {32'h3f6b3888, 32'h3f160e44} /* (20, 4, 22) {real, imag} */,
  {32'h3de3fa00, 32'hbf016754} /* (20, 4, 21) {real, imag} */,
  {32'h3e5ac110, 32'h3f5cd2c8} /* (20, 4, 20) {real, imag} */,
  {32'hbe63b748, 32'h3f63f958} /* (20, 4, 19) {real, imag} */,
  {32'hbf864ad1, 32'hbe878b90} /* (20, 4, 18) {real, imag} */,
  {32'hbe241e20, 32'hbf48fd78} /* (20, 4, 17) {real, imag} */,
  {32'h3ec1b800, 32'h3e164df0} /* (20, 4, 16) {real, imag} */,
  {32'h3f3e8d14, 32'h3e7508d0} /* (20, 4, 15) {real, imag} */,
  {32'h3f4c2076, 32'h3eeb7e60} /* (20, 4, 14) {real, imag} */,
  {32'h3e82935d, 32'hbe047510} /* (20, 4, 13) {real, imag} */,
  {32'h3f1eaff8, 32'hbf2cdc78} /* (20, 4, 12) {real, imag} */,
  {32'h3ede1b8a, 32'h3e90d848} /* (20, 4, 11) {real, imag} */,
  {32'h3f5c1086, 32'hbe474d90} /* (20, 4, 10) {real, imag} */,
  {32'hbdf97f10, 32'hbe5ad120} /* (20, 4, 9) {real, imag} */,
  {32'hbf9510e2, 32'h3f28d03c} /* (20, 4, 8) {real, imag} */,
  {32'hbf308a92, 32'h3e814448} /* (20, 4, 7) {real, imag} */,
  {32'h3ef38895, 32'h3eaaad74} /* (20, 4, 6) {real, imag} */,
  {32'h3fb162b0, 32'hbf3c91d1} /* (20, 4, 5) {real, imag} */,
  {32'h3fa3c0dd, 32'hbf3953a0} /* (20, 4, 4) {real, imag} */,
  {32'h3e4dd4cc, 32'h3f708aba} /* (20, 4, 3) {real, imag} */,
  {32'hbf2d3b48, 32'hbe79c750} /* (20, 4, 2) {real, imag} */,
  {32'hbec403fa, 32'hbed72318} /* (20, 4, 1) {real, imag} */,
  {32'h3d801320, 32'h3cd45ac0} /* (20, 4, 0) {real, imag} */,
  {32'hbebce9f0, 32'h3f7cddee} /* (20, 3, 31) {real, imag} */,
  {32'hbebf69ec, 32'h3ef8b5dc} /* (20, 3, 30) {real, imag} */,
  {32'h3e5f1280, 32'h3da0e970} /* (20, 3, 29) {real, imag} */,
  {32'h3e5c8b80, 32'hbed07488} /* (20, 3, 28) {real, imag} */,
  {32'hbeb65a5c, 32'hbee787f0} /* (20, 3, 27) {real, imag} */,
  {32'hbe8cc378, 32'hbec85a00} /* (20, 3, 26) {real, imag} */,
  {32'h3ef93446, 32'h3ea517e0} /* (20, 3, 25) {real, imag} */,
  {32'h3e9b9e50, 32'hbeb518e8} /* (20, 3, 24) {real, imag} */,
  {32'hbf1619dc, 32'hbf00c518} /* (20, 3, 23) {real, imag} */,
  {32'hbf6aa2d4, 32'h3f17ff28} /* (20, 3, 22) {real, imag} */,
  {32'hbb50a400, 32'h3eb6f938} /* (20, 3, 21) {real, imag} */,
  {32'h3ee79ee0, 32'h3e3f2e80} /* (20, 3, 20) {real, imag} */,
  {32'h3f2228b6, 32'h3dc0e2a0} /* (20, 3, 19) {real, imag} */,
  {32'h3d3f88c0, 32'hbf663f4c} /* (20, 3, 18) {real, imag} */,
  {32'h3d81ac40, 32'hbe07f1c0} /* (20, 3, 17) {real, imag} */,
  {32'hbe38f088, 32'h3f34f43d} /* (20, 3, 16) {real, imag} */,
  {32'h3ea676be, 32'h3e146a08} /* (20, 3, 15) {real, imag} */,
  {32'h3eca73a4, 32'h3fb3fd67} /* (20, 3, 14) {real, imag} */,
  {32'hbee67e08, 32'h3f96212c} /* (20, 3, 13) {real, imag} */,
  {32'hbcc9d180, 32'hbfa22394} /* (20, 3, 12) {real, imag} */,
  {32'hbf57b41e, 32'hbdf975a0} /* (20, 3, 11) {real, imag} */,
  {32'hbf6010a2, 32'h3f8ee702} /* (20, 3, 10) {real, imag} */,
  {32'hbf295baf, 32'h3fabff22} /* (20, 3, 9) {real, imag} */,
  {32'hbec24d20, 32'h3fbdeae6} /* (20, 3, 8) {real, imag} */,
  {32'hbdae7400, 32'h3dd29680} /* (20, 3, 7) {real, imag} */,
  {32'h3dfddaec, 32'hbf26851a} /* (20, 3, 6) {real, imag} */,
  {32'h3f098824, 32'hbfbe81b6} /* (20, 3, 5) {real, imag} */,
  {32'h3f527e74, 32'hbff36fe1} /* (20, 3, 4) {real, imag} */,
  {32'h3eaf7bd4, 32'hbf5ddb10} /* (20, 3, 3) {real, imag} */,
  {32'hbf3bffd2, 32'hbef6634c} /* (20, 3, 2) {real, imag} */,
  {32'hbf397252, 32'h3e589bfc} /* (20, 3, 1) {real, imag} */,
  {32'h3e13bc26, 32'h3e363a34} /* (20, 3, 0) {real, imag} */,
  {32'hbcbd3810, 32'h3e182ff0} /* (20, 2, 31) {real, imag} */,
  {32'h3e82e1de, 32'hbf6b79c4} /* (20, 2, 30) {real, imag} */,
  {32'h3fba9806, 32'hbf7e3660} /* (20, 2, 29) {real, imag} */,
  {32'h3ffc756c, 32'h3da175e0} /* (20, 2, 28) {real, imag} */,
  {32'h3f3deeb0, 32'h3dd0f700} /* (20, 2, 27) {real, imag} */,
  {32'h3f07017c, 32'hbe53d4d0} /* (20, 2, 26) {real, imag} */,
  {32'hbf59db14, 32'h3f39a93a} /* (20, 2, 25) {real, imag} */,
  {32'hbf412775, 32'h3f08a4ee} /* (20, 2, 24) {real, imag} */,
  {32'hbf1e29c4, 32'hbeb1d9e4} /* (20, 2, 23) {real, imag} */,
  {32'hbf17f207, 32'h3f82337e} /* (20, 2, 22) {real, imag} */,
  {32'h3f1a7862, 32'h3fc597c1} /* (20, 2, 21) {real, imag} */,
  {32'h3edb2815, 32'h3f663460} /* (20, 2, 20) {real, imag} */,
  {32'hbe1d6e98, 32'h3efe4a30} /* (20, 2, 19) {real, imag} */,
  {32'hbed876a8, 32'hbf90fd8e} /* (20, 2, 18) {real, imag} */,
  {32'hbd3ba4c0, 32'hbeffe000} /* (20, 2, 17) {real, imag} */,
  {32'h3d0bf890, 32'h3ef6dd40} /* (20, 2, 16) {real, imag} */,
  {32'hbdaa2c10, 32'h3e17a008} /* (20, 2, 15) {real, imag} */,
  {32'hbf128f74, 32'h40119dd8} /* (20, 2, 14) {real, imag} */,
  {32'hbf27fd38, 32'h3f8a6fb8} /* (20, 2, 13) {real, imag} */,
  {32'hbee2ebc4, 32'hbedc55b8} /* (20, 2, 12) {real, imag} */,
  {32'hbf18512e, 32'h3e552350} /* (20, 2, 11) {real, imag} */,
  {32'h3e2b96a0, 32'h3f38ddfc} /* (20, 2, 10) {real, imag} */,
  {32'h3f1cc16e, 32'h3f51eb28} /* (20, 2, 9) {real, imag} */,
  {32'h3ea98746, 32'h3f53bcec} /* (20, 2, 8) {real, imag} */,
  {32'h3ee762a8, 32'h3ea6fad0} /* (20, 2, 7) {real, imag} */,
  {32'hbf1b7c26, 32'hbdac87e0} /* (20, 2, 6) {real, imag} */,
  {32'h3f660cc6, 32'hbe482950} /* (20, 2, 5) {real, imag} */,
  {32'h3fa2bb68, 32'hbf83b8d8} /* (20, 2, 4) {real, imag} */,
  {32'h3f1c1a27, 32'hbe436060} /* (20, 2, 3) {real, imag} */,
  {32'hbdbfd6dd, 32'hba941400} /* (20, 2, 2) {real, imag} */,
  {32'h3e8a5700, 32'hbdbfb7d0} /* (20, 2, 1) {real, imag} */,
  {32'h3ea8e26a, 32'hbe135f50} /* (20, 2, 0) {real, imag} */,
  {32'hbcfd5380, 32'h3f1c4a8a} /* (20, 1, 31) {real, imag} */,
  {32'h3f01a9a2, 32'h3ea45cb0} /* (20, 1, 30) {real, imag} */,
  {32'h3f908e82, 32'h3c1d2580} /* (20, 1, 29) {real, imag} */,
  {32'h3fa07772, 32'h3db97a40} /* (20, 1, 28) {real, imag} */,
  {32'h3f7d1216, 32'h3f2fc4ff} /* (20, 1, 27) {real, imag} */,
  {32'h3f0cdddc, 32'hbe055be0} /* (20, 1, 26) {real, imag} */,
  {32'hbed5a468, 32'h3f3b11f2} /* (20, 1, 25) {real, imag} */,
  {32'hbe34de50, 32'h3f19ca46} /* (20, 1, 24) {real, imag} */,
  {32'h3e5d6570, 32'hbef36c88} /* (20, 1, 23) {real, imag} */,
  {32'hbf8cd6ae, 32'h3f4d09cc} /* (20, 1, 22) {real, imag} */,
  {32'hbf379d67, 32'h3ef1b668} /* (20, 1, 21) {real, imag} */,
  {32'h3e7cd8f2, 32'hbf08c326} /* (20, 1, 20) {real, imag} */,
  {32'hbeb147a8, 32'h3e181b18} /* (20, 1, 19) {real, imag} */,
  {32'hbf272818, 32'hbe1b61e0} /* (20, 1, 18) {real, imag} */,
  {32'hbf1094e2, 32'hbf9c466a} /* (20, 1, 17) {real, imag} */,
  {32'h3e4d5f20, 32'hbf219b82} /* (20, 1, 16) {real, imag} */,
  {32'h3ef5de05, 32'h3f071423} /* (20, 1, 15) {real, imag} */,
  {32'hbeb72cd8, 32'h4003d204} /* (20, 1, 14) {real, imag} */,
  {32'hbf4f96fc, 32'h3ea53d38} /* (20, 1, 13) {real, imag} */,
  {32'hbf0eb604, 32'hbf4b9140} /* (20, 1, 12) {real, imag} */,
  {32'h3f3d8578, 32'hbea328e0} /* (20, 1, 11) {real, imag} */,
  {32'h3fe4f827, 32'h3f07c8f0} /* (20, 1, 10) {real, imag} */,
  {32'h3f0d07cf, 32'hbe6f5b80} /* (20, 1, 9) {real, imag} */,
  {32'h3de988f0, 32'hbf0fcc32} /* (20, 1, 8) {real, imag} */,
  {32'h3e0cfc88, 32'h3f26f9fa} /* (20, 1, 7) {real, imag} */,
  {32'hbe4d8680, 32'h3f4f2440} /* (20, 1, 6) {real, imag} */,
  {32'h3fdddb24, 32'h3f5d8a53} /* (20, 1, 5) {real, imag} */,
  {32'h3fd59a80, 32'hbf33329a} /* (20, 1, 4) {real, imag} */,
  {32'hbc2379e0, 32'hbf528048} /* (20, 1, 3) {real, imag} */,
  {32'hbf04eaf6, 32'hbe857904} /* (20, 1, 2) {real, imag} */,
  {32'hbca05280, 32'hbe637648} /* (20, 1, 1) {real, imag} */,
  {32'h3e30a084, 32'h3e0a9c14} /* (20, 1, 0) {real, imag} */,
  {32'hbf1d3d21, 32'h3ecafc4c} /* (20, 0, 31) {real, imag} */,
  {32'hbe8639bc, 32'h3e7fad70} /* (20, 0, 30) {real, imag} */,
  {32'h3ece1524, 32'hbe868a5e} /* (20, 0, 29) {real, imag} */,
  {32'h3ebb5e1c, 32'h3dab4d40} /* (20, 0, 28) {real, imag} */,
  {32'h3f00b9f8, 32'h3f959728} /* (20, 0, 27) {real, imag} */,
  {32'h3e572198, 32'h3e0b18be} /* (20, 0, 26) {real, imag} */,
  {32'h3e412248, 32'h3f27caa4} /* (20, 0, 25) {real, imag} */,
  {32'h3ef6aeb4, 32'h3f2f6c60} /* (20, 0, 24) {real, imag} */,
  {32'h3eb3f2cc, 32'hbdcfb2d0} /* (20, 0, 23) {real, imag} */,
  {32'hbef07e90, 32'h3e124fa8} /* (20, 0, 22) {real, imag} */,
  {32'hbf080cf6, 32'h3d480cc0} /* (20, 0, 21) {real, imag} */,
  {32'hbe2d106c, 32'hbf59ec78} /* (20, 0, 20) {real, imag} */,
  {32'h3d9aabb0, 32'hbeeb37fa} /* (20, 0, 19) {real, imag} */,
  {32'h3f10c336, 32'h3e1b3598} /* (20, 0, 18) {real, imag} */,
  {32'h3e266b6f, 32'hbf4eef93} /* (20, 0, 17) {real, imag} */,
  {32'hbf0ab20c, 32'hbf13af55} /* (20, 0, 16) {real, imag} */,
  {32'h3eaa510c, 32'hbe04d84c} /* (20, 0, 15) {real, imag} */,
  {32'h3f1cd000, 32'h3f11783e} /* (20, 0, 14) {real, imag} */,
  {32'hbd9b83c0, 32'hbe707678} /* (20, 0, 13) {real, imag} */,
  {32'h3efc5402, 32'hbf117430} /* (20, 0, 12) {real, imag} */,
  {32'h3f8118d3, 32'h3df27260} /* (20, 0, 11) {real, imag} */,
  {32'h3f01d284, 32'h3f36f7ca} /* (20, 0, 10) {real, imag} */,
  {32'h3dcb5600, 32'h3ef41328} /* (20, 0, 9) {real, imag} */,
  {32'hbeafa064, 32'hbeeb2bf4} /* (20, 0, 8) {real, imag} */,
  {32'hbf0948d7, 32'h3e53a1a0} /* (20, 0, 7) {real, imag} */,
  {32'hbef2e922, 32'h3eee896c} /* (20, 0, 6) {real, imag} */,
  {32'h3f1fbf32, 32'h3e56a6ae} /* (20, 0, 5) {real, imag} */,
  {32'h3ea5954e, 32'h3e51ae40} /* (20, 0, 4) {real, imag} */,
  {32'hbce4ac98, 32'hbf152214} /* (20, 0, 3) {real, imag} */,
  {32'h3e711d70, 32'hbef4e530} /* (20, 0, 2) {real, imag} */,
  {32'h3f128a50, 32'hbeda6ea0} /* (20, 0, 1) {real, imag} */,
  {32'h3eb1a2c0, 32'hbe60fec6} /* (20, 0, 0) {real, imag} */,
  {32'h3e288860, 32'h3ecfdf3e} /* (19, 31, 31) {real, imag} */,
  {32'h3f4ae69f, 32'h3f3215ed} /* (19, 31, 30) {real, imag} */,
  {32'h3da954a8, 32'hbe783818} /* (19, 31, 29) {real, imag} */,
  {32'hbc2d4300, 32'h3c569780} /* (19, 31, 28) {real, imag} */,
  {32'hbe6bebb0, 32'h3f3026ec} /* (19, 31, 27) {real, imag} */,
  {32'hbf1cd991, 32'h3e7029f8} /* (19, 31, 26) {real, imag} */,
  {32'hbea47ac8, 32'h3e67ed60} /* (19, 31, 25) {real, imag} */,
  {32'hbf206883, 32'hbe2e6fc0} /* (19, 31, 24) {real, imag} */,
  {32'h3eae0bfe, 32'hbee3adac} /* (19, 31, 23) {real, imag} */,
  {32'h3f6cf37a, 32'h3bfdb000} /* (19, 31, 22) {real, imag} */,
  {32'h3db02fe0, 32'h3f0a2ec2} /* (19, 31, 21) {real, imag} */,
  {32'h3dcebf90, 32'h3ddf3bf0} /* (19, 31, 20) {real, imag} */,
  {32'hbd74b18c, 32'hbd5c9b60} /* (19, 31, 19) {real, imag} */,
  {32'h3eaf3a10, 32'h3e5d45fc} /* (19, 31, 18) {real, imag} */,
  {32'h3f5700c8, 32'hbf1ea2ed} /* (19, 31, 17) {real, imag} */,
  {32'h3f01b799, 32'hbf86901e} /* (19, 31, 16) {real, imag} */,
  {32'h3f1891f5, 32'hbf352eca} /* (19, 31, 15) {real, imag} */,
  {32'hbae76800, 32'h3e9c3ae0} /* (19, 31, 14) {real, imag} */,
  {32'hbf46bb72, 32'hbda075a0} /* (19, 31, 13) {real, imag} */,
  {32'hbf3cfaeb, 32'hbd34c1c0} /* (19, 31, 12) {real, imag} */,
  {32'hbeb4d99b, 32'h3efdb714} /* (19, 31, 11) {real, imag} */,
  {32'hbe19a4b0, 32'h3f6add80} /* (19, 31, 10) {real, imag} */,
  {32'h3ea278e8, 32'h3e2076f0} /* (19, 31, 9) {real, imag} */,
  {32'h3f1581a6, 32'hbeda184c} /* (19, 31, 8) {real, imag} */,
  {32'h3f214e0a, 32'hbe204f28} /* (19, 31, 7) {real, imag} */,
  {32'h3f371758, 32'h3ef0d4ec} /* (19, 31, 6) {real, imag} */,
  {32'hbefac8ea, 32'h3f610355} /* (19, 31, 5) {real, imag} */,
  {32'hbf70dc12, 32'h3f32e1f0} /* (19, 31, 4) {real, imag} */,
  {32'hbed17aa0, 32'hbf0419be} /* (19, 31, 3) {real, imag} */,
  {32'hbe2d986c, 32'hbe435cb8} /* (19, 31, 2) {real, imag} */,
  {32'h3e588610, 32'h3e8520e0} /* (19, 31, 1) {real, imag} */,
  {32'hbec62546, 32'h3ca5a200} /* (19, 31, 0) {real, imag} */,
  {32'hbe3bab40, 32'h3f0c2d20} /* (19, 30, 31) {real, imag} */,
  {32'h3f194366, 32'h3f0b4d5c} /* (19, 30, 30) {real, imag} */,
  {32'hbe5d4208, 32'hbf447a84} /* (19, 30, 29) {real, imag} */,
  {32'h3e1a1af0, 32'hbf14fdc8} /* (19, 30, 28) {real, imag} */,
  {32'h3e59df80, 32'hbf33666c} /* (19, 30, 27) {real, imag} */,
  {32'hbf61c235, 32'hbea50d4c} /* (19, 30, 26) {real, imag} */,
  {32'hbfb1da41, 32'h3eab5600} /* (19, 30, 25) {real, imag} */,
  {32'hc00d09cc, 32'hbf305e34} /* (19, 30, 24) {real, imag} */,
  {32'hbdfd7b70, 32'hbf455ed8} /* (19, 30, 23) {real, imag} */,
  {32'h3f55ef43, 32'h3f2f7f18} /* (19, 30, 22) {real, imag} */,
  {32'h3de19a2e, 32'h3ec979f8} /* (19, 30, 21) {real, imag} */,
  {32'h3e8d1448, 32'hbe0ade80} /* (19, 30, 20) {real, imag} */,
  {32'hbe0dca88, 32'hbe2b7200} /* (19, 30, 19) {real, imag} */,
  {32'h3efeb474, 32'h3ec9a8c8} /* (19, 30, 18) {real, imag} */,
  {32'h3fe525d4, 32'hbe97e370} /* (19, 30, 17) {real, imag} */,
  {32'h3f7020f4, 32'hbec23f10} /* (19, 30, 16) {real, imag} */,
  {32'h3f8e6b4c, 32'h3e3aad30} /* (19, 30, 15) {real, imag} */,
  {32'h3f5af094, 32'h3d01c840} /* (19, 30, 14) {real, imag} */,
  {32'hbe8ae272, 32'hbea66eb0} /* (19, 30, 13) {real, imag} */,
  {32'hbf66d3c3, 32'h3e9e7f38} /* (19, 30, 12) {real, imag} */,
  {32'hbf928df4, 32'h3f90eb22} /* (19, 30, 11) {real, imag} */,
  {32'hbfbb8f3c, 32'h3f56bccc} /* (19, 30, 10) {real, imag} */,
  {32'h3f4c72ee, 32'hbd88a220} /* (19, 30, 9) {real, imag} */,
  {32'h3fe415fa, 32'hbe619330} /* (19, 30, 8) {real, imag} */,
  {32'h3ee0a639, 32'h3e7f5610} /* (19, 30, 7) {real, imag} */,
  {32'hbf0018e8, 32'h3ed5918c} /* (19, 30, 6) {real, imag} */,
  {32'hbf9188dd, 32'h3fa6baa1} /* (19, 30, 5) {real, imag} */,
  {32'hbf871a60, 32'hbc930c00} /* (19, 30, 4) {real, imag} */,
  {32'h3c4434c0, 32'hbf62ae98} /* (19, 30, 3) {real, imag} */,
  {32'h3f0e6eef, 32'h3f12c110} /* (19, 30, 2) {real, imag} */,
  {32'h3fb4e40e, 32'h3f86a0e4} /* (19, 30, 1) {real, imag} */,
  {32'h3ef3d9e4, 32'h3dfa06b0} /* (19, 30, 0) {real, imag} */,
  {32'hbe80a7e0, 32'hbd8a8ce0} /* (19, 29, 31) {real, imag} */,
  {32'h3e0d5640, 32'hbc1ffd00} /* (19, 29, 30) {real, imag} */,
  {32'hbf15aede, 32'h3ec4d580} /* (19, 29, 29) {real, imag} */,
  {32'hbe901c00, 32'hbe8065f8} /* (19, 29, 28) {real, imag} */,
  {32'hbe0bd620, 32'hbf8cec3c} /* (19, 29, 27) {real, imag} */,
  {32'hbfa108d0, 32'hbef4ce68} /* (19, 29, 26) {real, imag} */,
  {32'hbf8c50d7, 32'hbf16de5c} /* (19, 29, 25) {real, imag} */,
  {32'hbf55ad63, 32'hbe9338f0} /* (19, 29, 24) {real, imag} */,
  {32'h3e0a440e, 32'h3dbf20e0} /* (19, 29, 23) {real, imag} */,
  {32'hbf06cc6e, 32'h3f8d5f42} /* (19, 29, 22) {real, imag} */,
  {32'hbf01074e, 32'hbea4faa4} /* (19, 29, 21) {real, imag} */,
  {32'hbf207a06, 32'hbf7b97c0} /* (19, 29, 20) {real, imag} */,
  {32'hbf2642a2, 32'hbf7b6eac} /* (19, 29, 19) {real, imag} */,
  {32'hbec2f8a8, 32'hbe7526c0} /* (19, 29, 18) {real, imag} */,
  {32'h3f232268, 32'hbe9aec20} /* (19, 29, 17) {real, imag} */,
  {32'h3ef5827a, 32'hbf03d2f8} /* (19, 29, 16) {real, imag} */,
  {32'h3f221197, 32'h3f243e14} /* (19, 29, 15) {real, imag} */,
  {32'h3f1140d0, 32'h3eaa6e90} /* (19, 29, 14) {real, imag} */,
  {32'h3f11e119, 32'hbd494180} /* (19, 29, 13) {real, imag} */,
  {32'h3e690c8e, 32'h3f37d574} /* (19, 29, 12) {real, imag} */,
  {32'hbf06a49e, 32'h3f83077a} /* (19, 29, 11) {real, imag} */,
  {32'hbf8f1f92, 32'h3f5ffa98} /* (19, 29, 10) {real, imag} */,
  {32'h3e82c5dc, 32'h3eeb4ba0} /* (19, 29, 9) {real, imag} */,
  {32'h3f7ebfe1, 32'h3d392a80} /* (19, 29, 8) {real, imag} */,
  {32'h3f2ee626, 32'hbe0d60c0} /* (19, 29, 7) {real, imag} */,
  {32'hbeff8e90, 32'hbe5ec508} /* (19, 29, 6) {real, imag} */,
  {32'hbd952ca0, 32'h3e92609c} /* (19, 29, 5) {real, imag} */,
  {32'h3f19c554, 32'hbf3da9dc} /* (19, 29, 4) {real, imag} */,
  {32'h3fc6bb35, 32'hbf460268} /* (19, 29, 3) {real, imag} */,
  {32'h3f03a9d5, 32'h3f8b51cc} /* (19, 29, 2) {real, imag} */,
  {32'h3f7043a8, 32'h3fa3aecc} /* (19, 29, 1) {real, imag} */,
  {32'h3f2a2c9b, 32'h3edc9edc} /* (19, 29, 0) {real, imag} */,
  {32'h3e7df464, 32'hbeac1354} /* (19, 28, 31) {real, imag} */,
  {32'h3e9f38f4, 32'hbd5e94c0} /* (19, 28, 30) {real, imag} */,
  {32'h3eaaaa57, 32'h3f1ead7c} /* (19, 28, 29) {real, imag} */,
  {32'hbebecd58, 32'hbe246be8} /* (19, 28, 28) {real, imag} */,
  {32'hbe0bab00, 32'hbe8d1e78} /* (19, 28, 27) {real, imag} */,
  {32'h3e1bf8ac, 32'h3f811f54} /* (19, 28, 26) {real, imag} */,
  {32'h3e0d2528, 32'hbd1eac80} /* (19, 28, 25) {real, imag} */,
  {32'h3eacaf5e, 32'h3e2688c0} /* (19, 28, 24) {real, imag} */,
  {32'hbed0952e, 32'h3f250df6} /* (19, 28, 23) {real, imag} */,
  {32'hbfe15730, 32'h3f3e9bdc} /* (19, 28, 22) {real, imag} */,
  {32'hbf4eed00, 32'hbf28e2d8} /* (19, 28, 21) {real, imag} */,
  {32'h3daf9e10, 32'hbfe6e0d8} /* (19, 28, 20) {real, imag} */,
  {32'hbca43700, 32'hbfd05240} /* (19, 28, 19) {real, imag} */,
  {32'h3dfe4730, 32'hbf1674b8} /* (19, 28, 18) {real, imag} */,
  {32'h3f3a72f6, 32'hbecdf760} /* (19, 28, 17) {real, imag} */,
  {32'h3f8e7b91, 32'hbf10c09c} /* (19, 28, 16) {real, imag} */,
  {32'h3fa7506e, 32'h3eed5578} /* (19, 28, 15) {real, imag} */,
  {32'h3efe019c, 32'h3b2ac400} /* (19, 28, 14) {real, imag} */,
  {32'h3e8571a2, 32'hbdff9ae0} /* (19, 28, 13) {real, imag} */,
  {32'h3e9482ca, 32'h3f6bf748} /* (19, 28, 12) {real, imag} */,
  {32'h3eefddfd, 32'h3f2e6f78} /* (19, 28, 11) {real, imag} */,
  {32'h3e89a190, 32'h3f317f9a} /* (19, 28, 10) {real, imag} */,
  {32'h3ec11658, 32'h3f1f300c} /* (19, 28, 9) {real, imag} */,
  {32'hbf19eb5c, 32'hbd838600} /* (19, 28, 8) {real, imag} */,
  {32'h3c844780, 32'hbf784f18} /* (19, 28, 7) {real, imag} */,
  {32'hbddd3688, 32'hbf2565cc} /* (19, 28, 6) {real, imag} */,
  {32'hbea3df98, 32'hbe9d40b8} /* (19, 28, 5) {real, imag} */,
  {32'h3e55b69c, 32'h3ed61600} /* (19, 28, 4) {real, imag} */,
  {32'h3ea755cc, 32'h3e1e3f60} /* (19, 28, 3) {real, imag} */,
  {32'hbf083b55, 32'h3f444f30} /* (19, 28, 2) {real, imag} */,
  {32'h3e6a06a0, 32'h3e6de030} /* (19, 28, 1) {real, imag} */,
  {32'h3f232169, 32'hbe69bdea} /* (19, 28, 0) {real, imag} */,
  {32'h3e899f90, 32'h3f2aa406} /* (19, 27, 31) {real, imag} */,
  {32'h3f5f7513, 32'h3e2d4010} /* (19, 27, 30) {real, imag} */,
  {32'h3fb29bb6, 32'hbece7470} /* (19, 27, 29) {real, imag} */,
  {32'h3ea1109c, 32'hbf8dcd28} /* (19, 27, 28) {real, imag} */,
  {32'h3ed36adc, 32'hbf3fee74} /* (19, 27, 27) {real, imag} */,
  {32'h3f22d300, 32'h3f81a658} /* (19, 27, 26) {real, imag} */,
  {32'h3d8df830, 32'h3efc1bc0} /* (19, 27, 25) {real, imag} */,
  {32'hbece6e1e, 32'h3e248280} /* (19, 27, 24) {real, imag} */,
  {32'hbfc8637c, 32'h3f1364a0} /* (19, 27, 23) {real, imag} */,
  {32'hbfce9203, 32'h3ed0e640} /* (19, 27, 22) {real, imag} */,
  {32'hbf0c7ff8, 32'h3e910dc0} /* (19, 27, 21) {real, imag} */,
  {32'hbd8409c0, 32'hbdbe0620} /* (19, 27, 20) {real, imag} */,
  {32'hbebcc13c, 32'hbd3c0e00} /* (19, 27, 19) {real, imag} */,
  {32'h3eae25b2, 32'hbe2328c0} /* (19, 27, 18) {real, imag} */,
  {32'h3f16c676, 32'hbf8721eb} /* (19, 27, 17) {real, imag} */,
  {32'h3ea1cd8c, 32'hbf5fc56c} /* (19, 27, 16) {real, imag} */,
  {32'hbddb0680, 32'hbf2974cc} /* (19, 27, 15) {real, imag} */,
  {32'hbcdd7de0, 32'hbeb73d28} /* (19, 27, 14) {real, imag} */,
  {32'h3f1214bd, 32'hbf24cb20} /* (19, 27, 13) {real, imag} */,
  {32'h3e4e4658, 32'hbe159980} /* (19, 27, 12) {real, imag} */,
  {32'h3f266139, 32'h3f24a06c} /* (19, 27, 11) {real, imag} */,
  {32'h3f1dee1a, 32'h3f7fd4f0} /* (19, 27, 10) {real, imag} */,
  {32'h3f90b571, 32'h3f87341c} /* (19, 27, 9) {real, imag} */,
  {32'hbf10e390, 32'h3e675660} /* (19, 27, 8) {real, imag} */,
  {32'hbf836196, 32'hbea6fed8} /* (19, 27, 7) {real, imag} */,
  {32'hbf0f670c, 32'hbf634337} /* (19, 27, 6) {real, imag} */,
  {32'hbf33c3ac, 32'hbef654e0} /* (19, 27, 5) {real, imag} */,
  {32'hbf50a5b8, 32'h3ec43920} /* (19, 27, 4) {real, imag} */,
  {32'hbf055b19, 32'hbf257a38} /* (19, 27, 3) {real, imag} */,
  {32'hbdd0b5d0, 32'h3e093b30} /* (19, 27, 2) {real, imag} */,
  {32'h3e57bd5a, 32'h3e08d7e8} /* (19, 27, 1) {real, imag} */,
  {32'h3ecf8ff1, 32'h3ec9197e} /* (19, 27, 0) {real, imag} */,
  {32'h3eacdad8, 32'h3f314cd3} /* (19, 26, 31) {real, imag} */,
  {32'h3f40753a, 32'h3ed4cbe8} /* (19, 26, 30) {real, imag} */,
  {32'h3f092ccc, 32'hbf945296} /* (19, 26, 29) {real, imag} */,
  {32'h3e007910, 32'hbfb34287} /* (19, 26, 28) {real, imag} */,
  {32'h3fb03d5a, 32'hbf2a60e4} /* (19, 26, 27) {real, imag} */,
  {32'h3f8f7260, 32'h3ecee6b0} /* (19, 26, 26) {real, imag} */,
  {32'h3f333378, 32'h3e7d2560} /* (19, 26, 25) {real, imag} */,
  {32'h3e00d8f8, 32'hbf391d88} /* (19, 26, 24) {real, imag} */,
  {32'hbf99db85, 32'hbd2e2c80} /* (19, 26, 23) {real, imag} */,
  {32'hbf8effe8, 32'h3d2e4e20} /* (19, 26, 22) {real, imag} */,
  {32'hbe16650c, 32'h3d0ad3a0} /* (19, 26, 21) {real, imag} */,
  {32'h3ef79f39, 32'h3eb14d90} /* (19, 26, 20) {real, imag} */,
  {32'h3f014ccc, 32'h3f1cb4c0} /* (19, 26, 19) {real, imag} */,
  {32'h3f859a3b, 32'h3e9bf080} /* (19, 26, 18) {real, imag} */,
  {32'hbdd53f00, 32'hbf810bd0} /* (19, 26, 17) {real, imag} */,
  {32'hbe0c2528, 32'h3c9c2080} /* (19, 26, 16) {real, imag} */,
  {32'h3ecd0a6a, 32'h3ee26b20} /* (19, 26, 15) {real, imag} */,
  {32'h3f5f8b36, 32'hbd83efc0} /* (19, 26, 14) {real, imag} */,
  {32'h3ef9170c, 32'hbf985996} /* (19, 26, 13) {real, imag} */,
  {32'h3e258150, 32'hbf574ac6} /* (19, 26, 12) {real, imag} */,
  {32'h3f1064f8, 32'h3eb9a6e8} /* (19, 26, 11) {real, imag} */,
  {32'h3eb2a971, 32'h3f4fadc8} /* (19, 26, 10) {real, imag} */,
  {32'h3f3d852a, 32'h3f406948} /* (19, 26, 9) {real, imag} */,
  {32'hbdf5a850, 32'h3f213450} /* (19, 26, 8) {real, imag} */,
  {32'hbee66e44, 32'h3f12107d} /* (19, 26, 7) {real, imag} */,
  {32'hbf46779a, 32'hbd22f800} /* (19, 26, 6) {real, imag} */,
  {32'hbf967844, 32'h3e133288} /* (19, 26, 5) {real, imag} */,
  {32'hbeb2a700, 32'h3ed02cc8} /* (19, 26, 4) {real, imag} */,
  {32'h3eb9081a, 32'hbe8588f0} /* (19, 26, 3) {real, imag} */,
  {32'h3f99a3fd, 32'hbe571760} /* (19, 26, 2) {real, imag} */,
  {32'h3f70ef82, 32'hbe042e70} /* (19, 26, 1) {real, imag} */,
  {32'h3e8c3748, 32'h3d399620} /* (19, 26, 0) {real, imag} */,
  {32'h3ee60144, 32'h3e7f75e0} /* (19, 25, 31) {real, imag} */,
  {32'hbe707698, 32'h3f0df18c} /* (19, 25, 30) {real, imag} */,
  {32'hbed3add6, 32'hbe3a53b0} /* (19, 25, 29) {real, imag} */,
  {32'h3b7a1380, 32'hbf9bb0be} /* (19, 25, 28) {real, imag} */,
  {32'h3fb117ae, 32'hbf41f49c} /* (19, 25, 27) {real, imag} */,
  {32'h3fca7fc7, 32'h3e494f20} /* (19, 25, 26) {real, imag} */,
  {32'h3f698c0e, 32'h3f278998} /* (19, 25, 25) {real, imag} */,
  {32'h3ef0a3d4, 32'hbeb54310} /* (19, 25, 24) {real, imag} */,
  {32'h3b45b800, 32'h3e1d2500} /* (19, 25, 23) {real, imag} */,
  {32'hbed4ce08, 32'h3efeaa20} /* (19, 25, 22) {real, imag} */,
  {32'h3f151d37, 32'h3f0e838e} /* (19, 25, 21) {real, imag} */,
  {32'h3eacca28, 32'h3f536280} /* (19, 25, 20) {real, imag} */,
  {32'hbe78460c, 32'h3f120db4} /* (19, 25, 19) {real, imag} */,
  {32'h3f98b0f8, 32'h3ed901b0} /* (19, 25, 18) {real, imag} */,
  {32'h3fbf07d9, 32'hbeb9b600} /* (19, 25, 17) {real, imag} */,
  {32'h3f37dc95, 32'h3ec76c14} /* (19, 25, 16) {real, imag} */,
  {32'h3d06c920, 32'h3f41be20} /* (19, 25, 15) {real, imag} */,
  {32'hbee18af0, 32'h3ef5fe80} /* (19, 25, 14) {real, imag} */,
  {32'hbe6323d8, 32'hbf124290} /* (19, 25, 13) {real, imag} */,
  {32'h3f07e1f3, 32'h3f5f55ce} /* (19, 25, 12) {real, imag} */,
  {32'h3e007706, 32'h3f653748} /* (19, 25, 11) {real, imag} */,
  {32'hbee83392, 32'h3e30a848} /* (19, 25, 10) {real, imag} */,
  {32'hbeda5d08, 32'hbf0b8f4c} /* (19, 25, 9) {real, imag} */,
  {32'hbee9a754, 32'h3e839178} /* (19, 25, 8) {real, imag} */,
  {32'hbeeec1fa, 32'h3cc2f080} /* (19, 25, 7) {real, imag} */,
  {32'hbf522bdc, 32'hbef9ab88} /* (19, 25, 6) {real, imag} */,
  {32'hbfa1188e, 32'h3f9ef8a0} /* (19, 25, 5) {real, imag} */,
  {32'hbb0ecc00, 32'h3f699b3c} /* (19, 25, 4) {real, imag} */,
  {32'hbe28a0f6, 32'hbda437c0} /* (19, 25, 3) {real, imag} */,
  {32'h3f083f9a, 32'hbe1963d0} /* (19, 25, 2) {real, imag} */,
  {32'h3f1d4883, 32'h3ee9e3fe} /* (19, 25, 1) {real, imag} */,
  {32'hbdac1274, 32'h3f459eb2} /* (19, 25, 0) {real, imag} */,
  {32'h3e7fced4, 32'hbd8b5940} /* (19, 24, 31) {real, imag} */,
  {32'hbf39cf8b, 32'h3ec21380} /* (19, 24, 30) {real, imag} */,
  {32'hbe702f24, 32'h3f34df48} /* (19, 24, 29) {real, imag} */,
  {32'h3e104a70, 32'hbda7ba40} /* (19, 24, 28) {real, imag} */,
  {32'hbd17ef60, 32'hbe58ce80} /* (19, 24, 27) {real, imag} */,
  {32'h3f469994, 32'h3ecb08b8} /* (19, 24, 26) {real, imag} */,
  {32'h3e82c368, 32'hbe842b20} /* (19, 24, 25) {real, imag} */,
  {32'h3f0c99b8, 32'hbee19048} /* (19, 24, 24) {real, imag} */,
  {32'h3f859505, 32'h3e59c2a8} /* (19, 24, 23) {real, imag} */,
  {32'h3e978940, 32'h3e922718} /* (19, 24, 22) {real, imag} */,
  {32'h3f33508c, 32'h3f7c8aaa} /* (19, 24, 21) {real, imag} */,
  {32'hbf106dc6, 32'h3f31d6c0} /* (19, 24, 20) {real, imag} */,
  {32'hbf4cab4d, 32'hbef0a9e0} /* (19, 24, 19) {real, imag} */,
  {32'hbe2b3a68, 32'hbf20dcec} /* (19, 24, 18) {real, imag} */,
  {32'h3f90c519, 32'hbe89d1a0} /* (19, 24, 17) {real, imag} */,
  {32'h3e8144f8, 32'hbe709380} /* (19, 24, 16) {real, imag} */,
  {32'hbf49d194, 32'hbe8beeb8} /* (19, 24, 15) {real, imag} */,
  {32'hbf9a74f8, 32'h3eb881b0} /* (19, 24, 14) {real, imag} */,
  {32'hbdffe110, 32'h3dd64ad0} /* (19, 24, 13) {real, imag} */,
  {32'h3d899b20, 32'h3fb021fc} /* (19, 24, 12) {real, imag} */,
  {32'hbfaae1a2, 32'h3f759cdc} /* (19, 24, 11) {real, imag} */,
  {32'hbf97c3e0, 32'h3efee750} /* (19, 24, 10) {real, imag} */,
  {32'hbf043a29, 32'hbf2f0250} /* (19, 24, 9) {real, imag} */,
  {32'hbf2ed3f6, 32'hbea883e0} /* (19, 24, 8) {real, imag} */,
  {32'hbe650ca4, 32'hbe17bc80} /* (19, 24, 7) {real, imag} */,
  {32'hbe1f2ba0, 32'hbf5f2ffc} /* (19, 24, 6) {real, imag} */,
  {32'hbea6fac6, 32'h3f390e10} /* (19, 24, 5) {real, imag} */,
  {32'hbdddb3c8, 32'h3edfef50} /* (19, 24, 4) {real, imag} */,
  {32'hbf34e182, 32'hbe535540} /* (19, 24, 3) {real, imag} */,
  {32'h3ea090d2, 32'h3e76b4e0} /* (19, 24, 2) {real, imag} */,
  {32'h3f613710, 32'h3f8f2e98} /* (19, 24, 1) {real, imag} */,
  {32'h3efc374e, 32'h3f60653c} /* (19, 24, 0) {real, imag} */,
  {32'h3eb438ba, 32'h3f041234} /* (19, 23, 31) {real, imag} */,
  {32'h3e1b7230, 32'h3fbe08f2} /* (19, 23, 30) {real, imag} */,
  {32'h3d878ae8, 32'h3f8fa2ba} /* (19, 23, 29) {real, imag} */,
  {32'h3ca9a6e0, 32'hbdd31180} /* (19, 23, 28) {real, imag} */,
  {32'hbe3a5a10, 32'hbf31eb88} /* (19, 23, 27) {real, imag} */,
  {32'h3e0123c4, 32'hbeba6a40} /* (19, 23, 26) {real, imag} */,
  {32'h3f2e13c3, 32'hbf0d3cb8} /* (19, 23, 25) {real, imag} */,
  {32'h3f9e8d24, 32'h3d81f940} /* (19, 23, 24) {real, imag} */,
  {32'h3ed36d7c, 32'h3e22cbd0} /* (19, 23, 23) {real, imag} */,
  {32'hbe653c40, 32'h3f11ead8} /* (19, 23, 22) {real, imag} */,
  {32'h3e51be60, 32'h3fb10cb2} /* (19, 23, 21) {real, imag} */,
  {32'hbf4250fa, 32'h3e604b30} /* (19, 23, 20) {real, imag} */,
  {32'hbda025d0, 32'hbf29b3e4} /* (19, 23, 19) {real, imag} */,
  {32'hbf113e9f, 32'hbeca9a28} /* (19, 23, 18) {real, imag} */,
  {32'hbea72862, 32'h3e8166a8} /* (19, 23, 17) {real, imag} */,
  {32'hbee85d30, 32'h3deab390} /* (19, 23, 16) {real, imag} */,
  {32'hbf39452f, 32'hbec65ef0} /* (19, 23, 15) {real, imag} */,
  {32'hbf068885, 32'h3d85afc0} /* (19, 23, 14) {real, imag} */,
  {32'hbebac07a, 32'h3f044d42} /* (19, 23, 13) {real, imag} */,
  {32'hbf0eb86c, 32'h3f55cd91} /* (19, 23, 12) {real, imag} */,
  {32'hbf91b74b, 32'h3cf2ee80} /* (19, 23, 11) {real, imag} */,
  {32'hbe716cce, 32'hbd75f0c0} /* (19, 23, 10) {real, imag} */,
  {32'hbdb7e468, 32'h3f0ee810} /* (19, 23, 9) {real, imag} */,
  {32'hbdfe5918, 32'h3e6acc60} /* (19, 23, 8) {real, imag} */,
  {32'h3e5b3dd0, 32'h3f60c388} /* (19, 23, 7) {real, imag} */,
  {32'h3e6593de, 32'hbe084d40} /* (19, 23, 6) {real, imag} */,
  {32'h3f56ce23, 32'h3ec14780} /* (19, 23, 5) {real, imag} */,
  {32'h3e805af4, 32'h3c6b5b00} /* (19, 23, 4) {real, imag} */,
  {32'hbf75d882, 32'hbeee85b8} /* (19, 23, 3) {real, imag} */,
  {32'hbf858e72, 32'h3e68f840} /* (19, 23, 2) {real, imag} */,
  {32'hbebfe0c6, 32'h3f8475cc} /* (19, 23, 1) {real, imag} */,
  {32'h3e38a7a4, 32'h3f25227c} /* (19, 23, 0) {real, imag} */,
  {32'h3e94bd58, 32'h3e955384} /* (19, 22, 31) {real, imag} */,
  {32'hbd5a6cb0, 32'h3fb84f09} /* (19, 22, 30) {real, imag} */,
  {32'hbf0cf06e, 32'h3f95958c} /* (19, 22, 29) {real, imag} */,
  {32'hbebfa31c, 32'hbf1b5908} /* (19, 22, 28) {real, imag} */,
  {32'h3dc7d080, 32'hbf39b594} /* (19, 22, 27) {real, imag} */,
  {32'h3e81d93a, 32'hbf0949d4} /* (19, 22, 26) {real, imag} */,
  {32'h3e500774, 32'hbf2d7e78} /* (19, 22, 25) {real, imag} */,
  {32'h3db7b8c0, 32'hbd7decc0} /* (19, 22, 24) {real, imag} */,
  {32'hbf1e9558, 32'hbe6b6e20} /* (19, 22, 23) {real, imag} */,
  {32'hbf1cd056, 32'h3e618d10} /* (19, 22, 22) {real, imag} */,
  {32'hbee4bb99, 32'h3f9df7d3} /* (19, 22, 21) {real, imag} */,
  {32'hbf03f5ea, 32'h3f1c808a} /* (19, 22, 20) {real, imag} */,
  {32'h3ede2907, 32'hbf38b8a4} /* (19, 22, 19) {real, imag} */,
  {32'hbd026940, 32'h3cb05b80} /* (19, 22, 18) {real, imag} */,
  {32'hbf6514b1, 32'h3ecdbc98} /* (19, 22, 17) {real, imag} */,
  {32'hbfa711b4, 32'h3dcc5c40} /* (19, 22, 16) {real, imag} */,
  {32'hbf551866, 32'hbee82314} /* (19, 22, 15) {real, imag} */,
  {32'hbf6f6f44, 32'hbef74760} /* (19, 22, 14) {real, imag} */,
  {32'hbf6b7958, 32'h3e6929c0} /* (19, 22, 13) {real, imag} */,
  {32'hbee91070, 32'h3f6648e6} /* (19, 22, 12) {real, imag} */,
  {32'h3ea534e7, 32'hbcf18e60} /* (19, 22, 11) {real, imag} */,
  {32'hbe23bf08, 32'h3d4ac920} /* (19, 22, 10) {real, imag} */,
  {32'hbf65fdc4, 32'h3d760b40} /* (19, 22, 9) {real, imag} */,
  {32'hbf04ca55, 32'hbf43d218} /* (19, 22, 8) {real, imag} */,
  {32'hbde91ff0, 32'hbdaf1980} /* (19, 22, 7) {real, imag} */,
  {32'hbeb20e38, 32'hbdf790e0} /* (19, 22, 6) {real, imag} */,
  {32'h3f087ff7, 32'hbf63ac9c} /* (19, 22, 5) {real, imag} */,
  {32'h3ef3c0dc, 32'hbef47ab8} /* (19, 22, 4) {real, imag} */,
  {32'h3ed5f2b8, 32'hbf254770} /* (19, 22, 3) {real, imag} */,
  {32'hbee21490, 32'hbf8ed530} /* (19, 22, 2) {real, imag} */,
  {32'hbece4a45, 32'hbc9b5ec0} /* (19, 22, 1) {real, imag} */,
  {32'h3b1675c0, 32'h3f05daf6} /* (19, 22, 0) {real, imag} */,
  {32'h3e7f7edc, 32'hbf473bf0} /* (19, 21, 31) {real, imag} */,
  {32'hbe411bc6, 32'hbf19e1ec} /* (19, 21, 30) {real, imag} */,
  {32'hbf7bce70, 32'h3f5bb43d} /* (19, 21, 29) {real, imag} */,
  {32'hbf9a10e4, 32'hbe9a65ec} /* (19, 21, 28) {real, imag} */,
  {32'hbd9a55f0, 32'hbf3dde84} /* (19, 21, 27) {real, imag} */,
  {32'h3f0fb85e, 32'hbc8be6e0} /* (19, 21, 26) {real, imag} */,
  {32'hbf245982, 32'hbef367b4} /* (19, 21, 25) {real, imag} */,
  {32'hbf60db53, 32'hbcd6bcc0} /* (19, 21, 24) {real, imag} */,
  {32'hbea40ca8, 32'hbe5049f8} /* (19, 21, 23) {real, imag} */,
  {32'h3e7bbea4, 32'hbf505393} /* (19, 21, 22) {real, imag} */,
  {32'hbc85af78, 32'h3e10dba0} /* (19, 21, 21) {real, imag} */,
  {32'h3d19b220, 32'h3f2b1654} /* (19, 21, 20) {real, imag} */,
  {32'h3eb4c600, 32'hbeabf1f4} /* (19, 21, 19) {real, imag} */,
  {32'h3e1d53a4, 32'h3d9a9dc0} /* (19, 21, 18) {real, imag} */,
  {32'h3f059460, 32'h3dced5d0} /* (19, 21, 17) {real, imag} */,
  {32'hbe9e45c2, 32'hbf65d268} /* (19, 21, 16) {real, imag} */,
  {32'hbf0dea14, 32'h3da8afd0} /* (19, 21, 15) {real, imag} */,
  {32'hbf1cf42c, 32'h3e51e330} /* (19, 21, 14) {real, imag} */,
  {32'hbefb176c, 32'hbd4ebbc0} /* (19, 21, 13) {real, imag} */,
  {32'hbdeb9810, 32'hbc885320} /* (19, 21, 12) {real, imag} */,
  {32'h3f8d6d41, 32'hbebb7df7} /* (19, 21, 11) {real, imag} */,
  {32'h3e793d80, 32'hbf582481} /* (19, 21, 10) {real, imag} */,
  {32'hbe21b5de, 32'hbfc4b99c} /* (19, 21, 9) {real, imag} */,
  {32'h3d1c7310, 32'hbfcec69e} /* (19, 21, 8) {real, imag} */,
  {32'hbd96a4c0, 32'hbf3e81b7} /* (19, 21, 7) {real, imag} */,
  {32'hbea11b10, 32'hbe37d334} /* (19, 21, 6) {real, imag} */,
  {32'h3e07f0da, 32'hbf4f3940} /* (19, 21, 5) {real, imag} */,
  {32'hbeff576c, 32'hbf05c22c} /* (19, 21, 4) {real, imag} */,
  {32'h3e746ae6, 32'hbe10e990} /* (19, 21, 3) {real, imag} */,
  {32'hbeb06acd, 32'hbfc3f369} /* (19, 21, 2) {real, imag} */,
  {32'hbf17293c, 32'hbf20661a} /* (19, 21, 1) {real, imag} */,
  {32'h3d8e2410, 32'h3c1fd368} /* (19, 21, 0) {real, imag} */,
  {32'h3e20b250, 32'hbd52e680} /* (19, 20, 31) {real, imag} */,
  {32'h3e9030ce, 32'hbefdfd28} /* (19, 20, 30) {real, imag} */,
  {32'hbebd022c, 32'h3f66e4e4} /* (19, 20, 29) {real, imag} */,
  {32'hbf5fdb86, 32'hbe434da0} /* (19, 20, 28) {real, imag} */,
  {32'h3ed94e68, 32'hbfa0fdec} /* (19, 20, 27) {real, imag} */,
  {32'h3e167cc0, 32'hbeddbcd0} /* (19, 20, 26) {real, imag} */,
  {32'hbe62e660, 32'hbd562e80} /* (19, 20, 25) {real, imag} */,
  {32'hbf4207c8, 32'hbf066da8} /* (19, 20, 24) {real, imag} */,
  {32'hbfb3e023, 32'h3e722080} /* (19, 20, 23) {real, imag} */,
  {32'hbef8df4f, 32'h3eb7b140} /* (19, 20, 22) {real, imag} */,
  {32'h3f27156c, 32'hbd8a5490} /* (19, 20, 21) {real, imag} */,
  {32'h3e9d84d4, 32'h3e52e128} /* (19, 20, 20) {real, imag} */,
  {32'h3ee8dcd0, 32'h3e676f30} /* (19, 20, 19) {real, imag} */,
  {32'h3ee83c30, 32'hbca3c480} /* (19, 20, 18) {real, imag} */,
  {32'h3fc031ce, 32'h3f010260} /* (19, 20, 17) {real, imag} */,
  {32'h3f23662b, 32'hbf1a0bd4} /* (19, 20, 16) {real, imag} */,
  {32'hbeb59340, 32'h3e516660} /* (19, 20, 15) {real, imag} */,
  {32'hbf34acdd, 32'h3f3e1e68} /* (19, 20, 14) {real, imag} */,
  {32'hbe82309d, 32'h3f8b53aa} /* (19, 20, 13) {real, imag} */,
  {32'h3ee46b34, 32'h3f0aa4f4} /* (19, 20, 12) {real, imag} */,
  {32'h3f785a2f, 32'hbea2eb20} /* (19, 20, 11) {real, imag} */,
  {32'h3fa3b374, 32'hbea4a362} /* (19, 20, 10) {real, imag} */,
  {32'h3dc26de4, 32'hbefdc2c0} /* (19, 20, 9) {real, imag} */,
  {32'hbebb2692, 32'hbee443b0} /* (19, 20, 8) {real, imag} */,
  {32'h3f1f0e04, 32'h3f0a0254} /* (19, 20, 7) {real, imag} */,
  {32'h3f99833f, 32'hbd429d00} /* (19, 20, 6) {real, imag} */,
  {32'h3f88a3cb, 32'hbf93a897} /* (19, 20, 5) {real, imag} */,
  {32'hbedc189c, 32'hbf58c5a8} /* (19, 20, 4) {real, imag} */,
  {32'hbfb7c143, 32'h3f149a00} /* (19, 20, 3) {real, imag} */,
  {32'hbf6d27f2, 32'hbeee674c} /* (19, 20, 2) {real, imag} */,
  {32'hbd9f9148, 32'hbe516430} /* (19, 20, 1) {real, imag} */,
  {32'hbd367200, 32'hbd882220} /* (19, 20, 0) {real, imag} */,
  {32'hbea1b07d, 32'h3f599d60} /* (19, 19, 31) {real, imag} */,
  {32'hbcff21a0, 32'h3e3df900} /* (19, 19, 30) {real, imag} */,
  {32'h3eb26814, 32'h3d97f070} /* (19, 19, 29) {real, imag} */,
  {32'h3d12c720, 32'hbf5ec8aa} /* (19, 19, 28) {real, imag} */,
  {32'h3f73f254, 32'hbf60adbc} /* (19, 19, 27) {real, imag} */,
  {32'h3f251b12, 32'hbf007a3c} /* (19, 19, 26) {real, imag} */,
  {32'h3f30434c, 32'hbf24aa8c} /* (19, 19, 25) {real, imag} */,
  {32'h3ee7559c, 32'hbf4f1198} /* (19, 19, 24) {real, imag} */,
  {32'hbf2fb280, 32'h3f5cca94} /* (19, 19, 23) {real, imag} */,
  {32'hbf6dd55b, 32'h3fa0a908} /* (19, 19, 22) {real, imag} */,
  {32'hbd44b980, 32'hbf026b0d} /* (19, 19, 21) {real, imag} */,
  {32'h3ddfbb30, 32'h3bdac800} /* (19, 19, 20) {real, imag} */,
  {32'hbd84ab70, 32'h3fc266ff} /* (19, 19, 19) {real, imag} */,
  {32'hbc7b0980, 32'h3f573004} /* (19, 19, 18) {real, imag} */,
  {32'h3f6f019c, 32'h3e9cee20} /* (19, 19, 17) {real, imag} */,
  {32'hbe1f5cf0, 32'hbe920e40} /* (19, 19, 16) {real, imag} */,
  {32'hbf1a081b, 32'h3e4ba888} /* (19, 19, 15) {real, imag} */,
  {32'hbe07e568, 32'hbedea670} /* (19, 19, 14) {real, imag} */,
  {32'h3f10d7ec, 32'hbe25acc0} /* (19, 19, 13) {real, imag} */,
  {32'h3ecd77a6, 32'hbe2a7310} /* (19, 19, 12) {real, imag} */,
  {32'h3eb8a862, 32'hbf81f915} /* (19, 19, 11) {real, imag} */,
  {32'h3f6b76da, 32'hbeba0170} /* (19, 19, 10) {real, imag} */,
  {32'h3e28cd38, 32'h3e19d9e0} /* (19, 19, 9) {real, imag} */,
  {32'hbf040f41, 32'h3f233c10} /* (19, 19, 8) {real, imag} */,
  {32'hbcd401c0, 32'h3f5830a8} /* (19, 19, 7) {real, imag} */,
  {32'h3da85d40, 32'hbe10d980} /* (19, 19, 6) {real, imag} */,
  {32'h3d93c3c8, 32'hbe0578a0} /* (19, 19, 5) {real, imag} */,
  {32'hbd1cb440, 32'hbdacc7c0} /* (19, 19, 4) {real, imag} */,
  {32'hbf4510b8, 32'hbecaa828} /* (19, 19, 3) {real, imag} */,
  {32'hbf93375a, 32'hbf188a08} /* (19, 19, 2) {real, imag} */,
  {32'hbea19a32, 32'h3ecae0d0} /* (19, 19, 1) {real, imag} */,
  {32'hbe2282a2, 32'h3e078670} /* (19, 19, 0) {real, imag} */,
  {32'hbf21601a, 32'h3e91e040} /* (19, 18, 31) {real, imag} */,
  {32'hbf2c81e0, 32'hbebef210} /* (19, 18, 30) {real, imag} */,
  {32'h3e52c318, 32'hbe19f900} /* (19, 18, 29) {real, imag} */,
  {32'hbe1289de, 32'h3d854b40} /* (19, 18, 28) {real, imag} */,
  {32'hbeb05ab8, 32'h3ed25638} /* (19, 18, 27) {real, imag} */,
  {32'h3e76aab4, 32'h3e8fecb0} /* (19, 18, 26) {real, imag} */,
  {32'h3f01351e, 32'hbf296a0a} /* (19, 18, 25) {real, imag} */,
  {32'h3ed64b60, 32'h3f0f1114} /* (19, 18, 24) {real, imag} */,
  {32'h3d6c55c0, 32'h3fa7726a} /* (19, 18, 23) {real, imag} */,
  {32'hbf17bd5c, 32'h3ec88240} /* (19, 18, 22) {real, imag} */,
  {32'hbe52ae48, 32'hbe092130} /* (19, 18, 21) {real, imag} */,
  {32'hbf37af21, 32'h3e25b6c0} /* (19, 18, 20) {real, imag} */,
  {32'hbf902feb, 32'h3fa6d32a} /* (19, 18, 19) {real, imag} */,
  {32'h3da71240, 32'h3eb04dc0} /* (19, 18, 18) {real, imag} */,
  {32'h3f020486, 32'hbed640a8} /* (19, 18, 17) {real, imag} */,
  {32'hbf18bb30, 32'hbf34dc84} /* (19, 18, 16) {real, imag} */,
  {32'hbf15a9cc, 32'hbf3cb270} /* (19, 18, 15) {real, imag} */,
  {32'hbdb4b2a0, 32'hbfaf141c} /* (19, 18, 14) {real, imag} */,
  {32'h3f2e96f6, 32'hbfb5ea80} /* (19, 18, 13) {real, imag} */,
  {32'h3ebbf424, 32'hbf1bc4b8} /* (19, 18, 12) {real, imag} */,
  {32'hbcdcd8c0, 32'hbf091eb4} /* (19, 18, 11) {real, imag} */,
  {32'hbf6fd7a0, 32'hbfa56f69} /* (19, 18, 10) {real, imag} */,
  {32'hbf48dc9c, 32'hbe781170} /* (19, 18, 9) {real, imag} */,
  {32'hbe9327ee, 32'h3cb4bc00} /* (19, 18, 8) {real, imag} */,
  {32'hbf361a6c, 32'hbf2b5abc} /* (19, 18, 7) {real, imag} */,
  {32'hbf8d674a, 32'hbe986330} /* (19, 18, 6) {real, imag} */,
  {32'hbf31fc3c, 32'h3e2b7c30} /* (19, 18, 5) {real, imag} */,
  {32'hbd685cc0, 32'hbdd7ed80} /* (19, 18, 4) {real, imag} */,
  {32'hbe5e36f0, 32'hbe4b3010} /* (19, 18, 3) {real, imag} */,
  {32'h3c145be0, 32'hbefcc980} /* (19, 18, 2) {real, imag} */,
  {32'h3ee30eac, 32'h3eedf158} /* (19, 18, 1) {real, imag} */,
  {32'hbe2dd8c8, 32'h3e96423c} /* (19, 18, 0) {real, imag} */,
  {32'hbf03c664, 32'h3eabe990} /* (19, 17, 31) {real, imag} */,
  {32'hbf560eb6, 32'hbe2120a0} /* (19, 17, 30) {real, imag} */,
  {32'hbf12b85c, 32'hbf1316d4} /* (19, 17, 29) {real, imag} */,
  {32'hbf7d7cb9, 32'h3fa0a584} /* (19, 17, 28) {real, imag} */,
  {32'hbfa04029, 32'h3f55785c} /* (19, 17, 27) {real, imag} */,
  {32'h3e26e2e0, 32'h3f1287b0} /* (19, 17, 26) {real, imag} */,
  {32'h3f14c46a, 32'h3f2a9884} /* (19, 17, 25) {real, imag} */,
  {32'h3ebff0e0, 32'h3f3e2e70} /* (19, 17, 24) {real, imag} */,
  {32'h3f0cfba1, 32'h3e887108} /* (19, 17, 23) {real, imag} */,
  {32'hbf2abf76, 32'hbec3fad0} /* (19, 17, 22) {real, imag} */,
  {32'hbf775228, 32'h3dde2c20} /* (19, 17, 21) {real, imag} */,
  {32'hbdb83518, 32'hbea75f00} /* (19, 17, 20) {real, imag} */,
  {32'hbe768720, 32'h3e982b14} /* (19, 17, 19) {real, imag} */,
  {32'hbd8f4be0, 32'h3d42a2c0} /* (19, 17, 18) {real, imag} */,
  {32'h3f11b9a0, 32'hbe3915b0} /* (19, 17, 17) {real, imag} */,
  {32'hbe020210, 32'hbec60d10} /* (19, 17, 16) {real, imag} */,
  {32'hbd3cb5a0, 32'hbf8ed58e} /* (19, 17, 15) {real, imag} */,
  {32'h3e8fb214, 32'hbfb202ac} /* (19, 17, 14) {real, imag} */,
  {32'h3ed41e58, 32'hbf4ba504} /* (19, 17, 13) {real, imag} */,
  {32'h3e92dec8, 32'hbe1eade0} /* (19, 17, 12) {real, imag} */,
  {32'h3f42ab7c, 32'h3d5217c0} /* (19, 17, 11) {real, imag} */,
  {32'hbf19b296, 32'hbf3e14ed} /* (19, 17, 10) {real, imag} */,
  {32'hbedc9860, 32'hbd6dbf00} /* (19, 17, 9) {real, imag} */,
  {32'h3ea360bc, 32'h3e366a60} /* (19, 17, 8) {real, imag} */,
  {32'h3e220736, 32'hbf484b2c} /* (19, 17, 7) {real, imag} */,
  {32'hbf66f76e, 32'hbf46132c} /* (19, 17, 6) {real, imag} */,
  {32'hbec32508, 32'hbe93f9c0} /* (19, 17, 5) {real, imag} */,
  {32'h3e8b4aa8, 32'hbf1cce3c} /* (19, 17, 4) {real, imag} */,
  {32'h3ece6f46, 32'hbe852ab0} /* (19, 17, 3) {real, imag} */,
  {32'h3ea67f31, 32'h3db2be80} /* (19, 17, 2) {real, imag} */,
  {32'h3f093b40, 32'hbc62d000} /* (19, 17, 1) {real, imag} */,
  {32'h3d094460, 32'hbd850a70} /* (19, 17, 0) {real, imag} */,
  {32'h3f144b7a, 32'h3c735400} /* (19, 16, 31) {real, imag} */,
  {32'h3dac8eb0, 32'h3e6f5c80} /* (19, 16, 30) {real, imag} */,
  {32'hbf3e9aab, 32'h3ea7e5f0} /* (19, 16, 29) {real, imag} */,
  {32'hbf1e59c0, 32'h3f5d6886} /* (19, 16, 28) {real, imag} */,
  {32'hbf8591f1, 32'h3f56a0ce} /* (19, 16, 27) {real, imag} */,
  {32'hbf49aaee, 32'h3e074148} /* (19, 16, 26) {real, imag} */,
  {32'hbe945658, 32'h3efbfc28} /* (19, 16, 25) {real, imag} */,
  {32'hbebe37a9, 32'h3cf3b080} /* (19, 16, 24) {real, imag} */,
  {32'h3e84d292, 32'h3ec37638} /* (19, 16, 23) {real, imag} */,
  {32'hbed5b7d0, 32'h3efcf3a8} /* (19, 16, 22) {real, imag} */,
  {32'hbce06ae0, 32'h3ea959ae} /* (19, 16, 21) {real, imag} */,
  {32'h3fc388b4, 32'h3f0ff998} /* (19, 16, 20) {real, imag} */,
  {32'h3fd07504, 32'h3f8fd684} /* (19, 16, 19) {real, imag} */,
  {32'h3f882086, 32'h3e9dd34c} /* (19, 16, 18) {real, imag} */,
  {32'h3e04152c, 32'hbeb1b898} /* (19, 16, 17) {real, imag} */,
  {32'hbfa9a6fb, 32'hbf853878} /* (19, 16, 16) {real, imag} */,
  {32'hbf400869, 32'hbeffa500} /* (19, 16, 15) {real, imag} */,
  {32'h3f64e8f5, 32'hbf509250} /* (19, 16, 14) {real, imag} */,
  {32'hbe05ec7c, 32'hbb037400} /* (19, 16, 13) {real, imag} */,
  {32'hbfa06a94, 32'h3e9f216c} /* (19, 16, 12) {real, imag} */,
  {32'hbec3dd16, 32'h3f3858e3} /* (19, 16, 11) {real, imag} */,
  {32'hbef43d90, 32'h3da099a0} /* (19, 16, 10) {real, imag} */,
  {32'h3f1ea4d6, 32'hbe0ff880} /* (19, 16, 9) {real, imag} */,
  {32'h3faebd1c, 32'h3e044ed0} /* (19, 16, 8) {real, imag} */,
  {32'h3f5a7e70, 32'hbdc80d00} /* (19, 16, 7) {real, imag} */,
  {32'h3e01d550, 32'h3e1f50f0} /* (19, 16, 6) {real, imag} */,
  {32'h3f090740, 32'hbd9aa460} /* (19, 16, 5) {real, imag} */,
  {32'h3f848ac8, 32'hbd6a4740} /* (19, 16, 4) {real, imag} */,
  {32'h3f9fa327, 32'h3dbad060} /* (19, 16, 3) {real, imag} */,
  {32'h3ef37bbc, 32'h3e7cf760} /* (19, 16, 2) {real, imag} */,
  {32'hb9a1f000, 32'h3ee1c678} /* (19, 16, 1) {real, imag} */,
  {32'h3eb445f6, 32'h3f134ffc} /* (19, 16, 0) {real, imag} */,
  {32'h3f2052d1, 32'h3dcfd680} /* (19, 15, 31) {real, imag} */,
  {32'h3f926682, 32'h3ceb0d00} /* (19, 15, 30) {real, imag} */,
  {32'h3ea56cf8, 32'h3e877060} /* (19, 15, 29) {real, imag} */,
  {32'hbfac5555, 32'hbd38a400} /* (19, 15, 28) {real, imag} */,
  {32'hbfa1f686, 32'h3fb4098b} /* (19, 15, 27) {real, imag} */,
  {32'hbfe38e9a, 32'h3f383f5a} /* (19, 15, 26) {real, imag} */,
  {32'hbfd43eb4, 32'hbe346a10} /* (19, 15, 25) {real, imag} */,
  {32'hbf3b39f5, 32'hbe5c2c78} /* (19, 15, 24) {real, imag} */,
  {32'h3f279f94, 32'h3f05454c} /* (19, 15, 23) {real, imag} */,
  {32'hbec311c8, 32'h3fd51d77} /* (19, 15, 22) {real, imag} */,
  {32'hbe09a2d2, 32'h3f80c87e} /* (19, 15, 21) {real, imag} */,
  {32'h3f8ecd86, 32'h3efdbe20} /* (19, 15, 20) {real, imag} */,
  {32'h3fa1d0a2, 32'h3f836fba} /* (19, 15, 19) {real, imag} */,
  {32'h3ff1c4e4, 32'h3f3e160f} /* (19, 15, 18) {real, imag} */,
  {32'h3f198ed4, 32'h3dceccf0} /* (19, 15, 17) {real, imag} */,
  {32'hbf81233a, 32'hbf7128a0} /* (19, 15, 16) {real, imag} */,
  {32'hbf5ea5b5, 32'hbf384b30} /* (19, 15, 15) {real, imag} */,
  {32'h3e9d1f34, 32'hbed94c50} /* (19, 15, 14) {real, imag} */,
  {32'hbf155c83, 32'hbeb73a78} /* (19, 15, 13) {real, imag} */,
  {32'hc0114714, 32'hbef899d0} /* (19, 15, 12) {real, imag} */,
  {32'hbfd47323, 32'h3f13a884} /* (19, 15, 11) {real, imag} */,
  {32'hbf26c340, 32'hbeb35348} /* (19, 15, 10) {real, imag} */,
  {32'h3e8ba0d2, 32'hbf5c1c9c} /* (19, 15, 9) {real, imag} */,
  {32'h3f002cf2, 32'hbf8a5ddc} /* (19, 15, 8) {real, imag} */,
  {32'h3e947038, 32'hbc571800} /* (19, 15, 7) {real, imag} */,
  {32'h3ecdd330, 32'h3f479c6c} /* (19, 15, 6) {real, imag} */,
  {32'h3ed11028, 32'h3f6832c6} /* (19, 15, 5) {real, imag} */,
  {32'h3f31d8a8, 32'h3ef0d530} /* (19, 15, 4) {real, imag} */,
  {32'h3fe48e32, 32'h3eabc288} /* (19, 15, 3) {real, imag} */,
  {32'h3fcbd886, 32'h3e4efc70} /* (19, 15, 2) {real, imag} */,
  {32'hbf162136, 32'h3eb961e8} /* (19, 15, 1) {real, imag} */,
  {32'hbec9727d, 32'h3f56cac4} /* (19, 15, 0) {real, imag} */,
  {32'hbea206e3, 32'h3f2a30d2} /* (19, 14, 31) {real, imag} */,
  {32'h3ef4f000, 32'h3f524de8} /* (19, 14, 30) {real, imag} */,
  {32'h3e8fe020, 32'hbe0a1250} /* (19, 14, 29) {real, imag} */,
  {32'hbf6cf894, 32'hbf16f64a} /* (19, 14, 28) {real, imag} */,
  {32'hbf5af660, 32'h3f97071b} /* (19, 14, 27) {real, imag} */,
  {32'hbef3fc98, 32'hbcb21200} /* (19, 14, 26) {real, imag} */,
  {32'hbf705db4, 32'hbf64d808} /* (19, 14, 25) {real, imag} */,
  {32'hbf11347c, 32'hbe007eb0} /* (19, 14, 24) {real, imag} */,
  {32'h3f7097a0, 32'h3eb62998} /* (19, 14, 23) {real, imag} */,
  {32'h3f0a39b8, 32'h3fb816ec} /* (19, 14, 22) {real, imag} */,
  {32'h3c25b400, 32'h3fac28b2} /* (19, 14, 21) {real, imag} */,
  {32'hbee783cc, 32'h3e873dd4} /* (19, 14, 20) {real, imag} */,
  {32'h3e70f040, 32'h3f2eceda} /* (19, 14, 19) {real, imag} */,
  {32'h3f6a486a, 32'h3e3bccd8} /* (19, 14, 18) {real, imag} */,
  {32'h3e553a64, 32'hbe800268} /* (19, 14, 17) {real, imag} */,
  {32'hbf24f4cc, 32'hbe923198} /* (19, 14, 16) {real, imag} */,
  {32'hbe462090, 32'hbe194700} /* (19, 14, 15) {real, imag} */,
  {32'h3c9c2940, 32'hbeb26a1c} /* (19, 14, 14) {real, imag} */,
  {32'hbf3b1569, 32'hbf32d5ec} /* (19, 14, 13) {real, imag} */,
  {32'hbf847f95, 32'hbf8843ea} /* (19, 14, 12) {real, imag} */,
  {32'h3f0a9878, 32'hbda60260} /* (19, 14, 11) {real, imag} */,
  {32'h3f7850fa, 32'hbe689c30} /* (19, 14, 10) {real, imag} */,
  {32'h3eca2694, 32'h3d251f80} /* (19, 14, 9) {real, imag} */,
  {32'hbed6cae4, 32'hbd827300} /* (19, 14, 8) {real, imag} */,
  {32'hbf6fbffc, 32'h3e363aa0} /* (19, 14, 7) {real, imag} */,
  {32'hbed76c66, 32'h3ea9bbc0} /* (19, 14, 6) {real, imag} */,
  {32'hbf49ca52, 32'h3f12d484} /* (19, 14, 5) {real, imag} */,
  {32'hbed789d8, 32'h3d3e0540} /* (19, 14, 4) {real, imag} */,
  {32'h3f4e7fd6, 32'h3c8f6080} /* (19, 14, 3) {real, imag} */,
  {32'h3f97a45e, 32'hbdbd6530} /* (19, 14, 2) {real, imag} */,
  {32'hbf6dd810, 32'h3e2c1558} /* (19, 14, 1) {real, imag} */,
  {32'hbf4b6a11, 32'h3e2fc010} /* (19, 14, 0) {real, imag} */,
  {32'h3d87afc4, 32'h3f3a8cb8} /* (19, 13, 31) {real, imag} */,
  {32'h3f348fbe, 32'h3f615e74} /* (19, 13, 30) {real, imag} */,
  {32'h3e96f880, 32'h3f06ae18} /* (19, 13, 29) {real, imag} */,
  {32'h3e645880, 32'h3ed50670} /* (19, 13, 28) {real, imag} */,
  {32'hbf936816, 32'h3d208a80} /* (19, 13, 27) {real, imag} */,
  {32'hbe962464, 32'hbf4473a4} /* (19, 13, 26) {real, imag} */,
  {32'h3d8287f0, 32'hbec0fc30} /* (19, 13, 25) {real, imag} */,
  {32'hbf1eea42, 32'h3dacc000} /* (19, 13, 24) {real, imag} */,
  {32'hbe981760, 32'h3ebd6830} /* (19, 13, 23) {real, imag} */,
  {32'h3ed49f40, 32'h3f6ea7b8} /* (19, 13, 22) {real, imag} */,
  {32'h3ee3b618, 32'h3eb1e802} /* (19, 13, 21) {real, imag} */,
  {32'hbf3c9f70, 32'hbe040940} /* (19, 13, 20) {real, imag} */,
  {32'h3e13c41c, 32'hbcdb9100} /* (19, 13, 19) {real, imag} */,
  {32'hbd84de80, 32'hbeae6a40} /* (19, 13, 18) {real, imag} */,
  {32'hbec142d4, 32'hbf7db728} /* (19, 13, 17) {real, imag} */,
  {32'hbee18a48, 32'hbf5e8e6c} /* (19, 13, 16) {real, imag} */,
  {32'hbf09a105, 32'h3f92ba9e} /* (19, 13, 15) {real, imag} */,
  {32'h3e114ddc, 32'h3f27960b} /* (19, 13, 14) {real, imag} */,
  {32'hbeb544f8, 32'hbeb103e0} /* (19, 13, 13) {real, imag} */,
  {32'hbbde8800, 32'hbf7b4340} /* (19, 13, 12) {real, imag} */,
  {32'h3fbe0da6, 32'hbea735f8} /* (19, 13, 11) {real, imag} */,
  {32'h3fce669f, 32'hbeb98200} /* (19, 13, 10) {real, imag} */,
  {32'h3f8ee8b6, 32'h3f20e5c8} /* (19, 13, 9) {real, imag} */,
  {32'h3edae4ec, 32'h3f31b0b8} /* (19, 13, 8) {real, imag} */,
  {32'hbe180e10, 32'h3ecfa80c} /* (19, 13, 7) {real, imag} */,
  {32'h3db67390, 32'hbea1fd00} /* (19, 13, 6) {real, imag} */,
  {32'hbf43ac4c, 32'hbe2e8aa0} /* (19, 13, 5) {real, imag} */,
  {32'hbf7ae65f, 32'h3e00f8c0} /* (19, 13, 4) {real, imag} */,
  {32'hbf0e6cb4, 32'h3f09ed88} /* (19, 13, 3) {real, imag} */,
  {32'h3e8aee38, 32'h3f528aca} /* (19, 13, 2) {real, imag} */,
  {32'hbea22fa3, 32'h3faf18f0} /* (19, 13, 1) {real, imag} */,
  {32'hbf3a2a2e, 32'h3eb14a90} /* (19, 13, 0) {real, imag} */,
  {32'h3eac5533, 32'h3f88820e} /* (19, 12, 31) {real, imag} */,
  {32'h3f58ad5a, 32'h3f8c3104} /* (19, 12, 30) {real, imag} */,
  {32'h3e9e51ec, 32'h3eb2cc28} /* (19, 12, 29) {real, imag} */,
  {32'hbdbf30d8, 32'h3f225340} /* (19, 12, 28) {real, imag} */,
  {32'hbf73a8b4, 32'h3ef88b40} /* (19, 12, 27) {real, imag} */,
  {32'hbf0432ae, 32'hbf3393b0} /* (19, 12, 26) {real, imag} */,
  {32'hbe43e0c0, 32'hbf6522c8} /* (19, 12, 25) {real, imag} */,
  {32'hbf38935e, 32'hbe9976d0} /* (19, 12, 24) {real, imag} */,
  {32'hbf4b5af5, 32'hbf21c468} /* (19, 12, 23) {real, imag} */,
  {32'hbf3ee2f9, 32'hbdb7c480} /* (19, 12, 22) {real, imag} */,
  {32'h3dd2daf8, 32'h3e4ec43c} /* (19, 12, 21) {real, imag} */,
  {32'hbef554d9, 32'h3ea5f1f0} /* (19, 12, 20) {real, imag} */,
  {32'hbebe9afa, 32'h3e9353d8} /* (19, 12, 19) {real, imag} */,
  {32'h3d74c020, 32'hbf14a8d8} /* (19, 12, 18) {real, imag} */,
  {32'h3efb1b88, 32'hbf207940} /* (19, 12, 17) {real, imag} */,
  {32'hbe81bea3, 32'hbe025f80} /* (19, 12, 16) {real, imag} */,
  {32'hbebd1740, 32'h3f8fa776} /* (19, 12, 15) {real, imag} */,
  {32'h3e11e5f7, 32'h3e238714} /* (19, 12, 14) {real, imag} */,
  {32'hbd431300, 32'hbebaa658} /* (19, 12, 13) {real, imag} */,
  {32'hbee28d74, 32'hbdbfb740} /* (19, 12, 12) {real, imag} */,
  {32'h3f8e1ff6, 32'hbf0cbc6e} /* (19, 12, 11) {real, imag} */,
  {32'h3eada028, 32'hbea8d8c4} /* (19, 12, 10) {real, imag} */,
  {32'hbea0009a, 32'h3f1819d8} /* (19, 12, 9) {real, imag} */,
  {32'h3f6b4e45, 32'h3e9023c8} /* (19, 12, 8) {real, imag} */,
  {32'h3edf26c0, 32'h3f88eee9} /* (19, 12, 7) {real, imag} */,
  {32'hbf059dcb, 32'h3f55e640} /* (19, 12, 6) {real, imag} */,
  {32'hbed45370, 32'hbe27b7c0} /* (19, 12, 5) {real, imag} */,
  {32'hbe20ccdc, 32'hbed21fa0} /* (19, 12, 4) {real, imag} */,
  {32'h3f4157b6, 32'hbf09ab50} /* (19, 12, 3) {real, imag} */,
  {32'h3fa22d3a, 32'h3f02b93c} /* (19, 12, 2) {real, imag} */,
  {32'h3f92acdd, 32'h3fda25d4} /* (19, 12, 1) {real, imag} */,
  {32'hbf09dca9, 32'h3f1f12f8} /* (19, 12, 0) {real, imag} */,
  {32'hbe96423e, 32'h3e1ba500} /* (19, 11, 31) {real, imag} */,
  {32'h3b618d00, 32'h3f1a1b44} /* (19, 11, 30) {real, imag} */,
  {32'h3ec0a216, 32'h3cac25c0} /* (19, 11, 29) {real, imag} */,
  {32'hbeffd746, 32'h3e3c6f70} /* (19, 11, 28) {real, imag} */,
  {32'hbd812578, 32'h3f5063c0} /* (19, 11, 27) {real, imag} */,
  {32'h3e676ec0, 32'h3d4d3640} /* (19, 11, 26) {real, imag} */,
  {32'hbd8ad010, 32'hbf3aed4c} /* (19, 11, 25) {real, imag} */,
  {32'h3d8e5ff4, 32'hbe606430} /* (19, 11, 24) {real, imag} */,
  {32'hbf338383, 32'hbeb04c8c} /* (19, 11, 23) {real, imag} */,
  {32'hbf8a5d03, 32'hbe866d58} /* (19, 11, 22) {real, imag} */,
  {32'hbe8e0420, 32'h3f1f8670} /* (19, 11, 21) {real, imag} */,
  {32'h3d7e2e60, 32'hbd8fce00} /* (19, 11, 20) {real, imag} */,
  {32'h3e9b42c4, 32'hbab28000} /* (19, 11, 19) {real, imag} */,
  {32'h3f002000, 32'hbe322320} /* (19, 11, 18) {real, imag} */,
  {32'hbebdcb48, 32'hbd226ca0} /* (19, 11, 17) {real, imag} */,
  {32'hbf7eab7e, 32'h3f910e79} /* (19, 11, 16) {real, imag} */,
  {32'h3f54ff8a, 32'h3f8478ac} /* (19, 11, 15) {real, imag} */,
  {32'h3fc8b817, 32'h3edb0ee4} /* (19, 11, 14) {real, imag} */,
  {32'h38f70000, 32'h3f03dc0c} /* (19, 11, 13) {real, imag} */,
  {32'hbf94dcde, 32'hbe4c7a70} /* (19, 11, 12) {real, imag} */,
  {32'h3e121b60, 32'h3e612838} /* (19, 11, 11) {real, imag} */,
  {32'hbefadeae, 32'h3e1fe170} /* (19, 11, 10) {real, imag} */,
  {32'hbf181e69, 32'hbe0c46c0} /* (19, 11, 9) {real, imag} */,
  {32'h3f889c7a, 32'hbe980b78} /* (19, 11, 8) {real, imag} */,
  {32'h3f8bf963, 32'h3ef47020} /* (19, 11, 7) {real, imag} */,
  {32'hbf719428, 32'hbf2b7fac} /* (19, 11, 6) {real, imag} */,
  {32'hbd2cbb30, 32'hbfc2100b} /* (19, 11, 5) {real, imag} */,
  {32'h3f1ce9cb, 32'hbf16bc78} /* (19, 11, 4) {real, imag} */,
  {32'h3f7ac96e, 32'hbed704ac} /* (19, 11, 3) {real, imag} */,
  {32'h3eefc6f0, 32'h3bce5600} /* (19, 11, 2) {real, imag} */,
  {32'h3f13f796, 32'h3eb28450} /* (19, 11, 1) {real, imag} */,
  {32'hbee6b447, 32'hbecdc8a8} /* (19, 11, 0) {real, imag} */,
  {32'hbf7969bc, 32'h3e8a9017} /* (19, 10, 31) {real, imag} */,
  {32'hbf9f6460, 32'h3edc34e8} /* (19, 10, 30) {real, imag} */,
  {32'hbef26537, 32'hbf296fcd} /* (19, 10, 29) {real, imag} */,
  {32'hbe734234, 32'hbe4c3084} /* (19, 10, 28) {real, imag} */,
  {32'h3edb5909, 32'hbf310473} /* (19, 10, 27) {real, imag} */,
  {32'h3ecca832, 32'h3da3f360} /* (19, 10, 26) {real, imag} */,
  {32'hbf3d1346, 32'h3f0583e8} /* (19, 10, 25) {real, imag} */,
  {32'hbf31e209, 32'h3e70547a} /* (19, 10, 24) {real, imag} */,
  {32'hbed8e0e8, 32'h3e5d7520} /* (19, 10, 23) {real, imag} */,
  {32'hbf268664, 32'h3e22e038} /* (19, 10, 22) {real, imag} */,
  {32'hbf888ac3, 32'h3ed057f8} /* (19, 10, 21) {real, imag} */,
  {32'hbe849870, 32'hbefb6ade} /* (19, 10, 20) {real, imag} */,
  {32'h3ec91a6e, 32'hbed790c0} /* (19, 10, 19) {real, imag} */,
  {32'h3f8f78b2, 32'h3fab290f} /* (19, 10, 18) {real, imag} */,
  {32'h3f8b3794, 32'h3fc188f6} /* (19, 10, 17) {real, imag} */,
  {32'hbf1608f0, 32'h3f8f5b1c} /* (19, 10, 16) {real, imag} */,
  {32'h3eb006f8, 32'hbd0b6308} /* (19, 10, 15) {real, imag} */,
  {32'h3fac69a9, 32'h3db0a168} /* (19, 10, 14) {real, imag} */,
  {32'h3e09bc92, 32'h3f2deb45} /* (19, 10, 13) {real, imag} */,
  {32'hbf06d8a8, 32'hbe737504} /* (19, 10, 12) {real, imag} */,
  {32'hbcf72040, 32'h3e79a3f4} /* (19, 10, 11) {real, imag} */,
  {32'h3e85e8b7, 32'h3e0de904} /* (19, 10, 10) {real, imag} */,
  {32'h3e0856f4, 32'h3ed58fdd} /* (19, 10, 9) {real, imag} */,
  {32'h3f8e895e, 32'h3f2a5fc4} /* (19, 10, 8) {real, imag} */,
  {32'h3fa97452, 32'h3f6dc8ea} /* (19, 10, 7) {real, imag} */,
  {32'hbe42a6e6, 32'hbf2b96c5} /* (19, 10, 6) {real, imag} */,
  {32'h3ee229de, 32'hbfe5ef80} /* (19, 10, 5) {real, imag} */,
  {32'h3f0647c0, 32'hbf41fc74} /* (19, 10, 4) {real, imag} */,
  {32'h3ed4dc22, 32'h3e828150} /* (19, 10, 3) {real, imag} */,
  {32'hbf447e5d, 32'hbeba7f9a} /* (19, 10, 2) {real, imag} */,
  {32'hbf223a7c, 32'hbf6a46af} /* (19, 10, 1) {real, imag} */,
  {32'hbf26cada, 32'hbf328530} /* (19, 10, 0) {real, imag} */,
  {32'hbf87a870, 32'h3e881720} /* (19, 9, 31) {real, imag} */,
  {32'hbfb617a1, 32'hbeb5f618} /* (19, 9, 30) {real, imag} */,
  {32'h3e9b8ed0, 32'hbf834142} /* (19, 9, 29) {real, imag} */,
  {32'h3f579e2e, 32'hbede43e0} /* (19, 9, 28) {real, imag} */,
  {32'hbeec68f4, 32'hbe896b40} /* (19, 9, 27) {real, imag} */,
  {32'hbf0d735d, 32'hbda45560} /* (19, 9, 26) {real, imag} */,
  {32'hbd5530f0, 32'h3d79af80} /* (19, 9, 25) {real, imag} */,
  {32'hbdd741b0, 32'hbeda13a0} /* (19, 9, 24) {real, imag} */,
  {32'h3f2900ca, 32'hbdcb49e0} /* (19, 9, 23) {real, imag} */,
  {32'h3db77f40, 32'hbf1f4100} /* (19, 9, 22) {real, imag} */,
  {32'hbf738f2e, 32'hbef992ac} /* (19, 9, 21) {real, imag} */,
  {32'hbf6fb136, 32'hbf52ebe4} /* (19, 9, 20) {real, imag} */,
  {32'hbf522788, 32'hbe67f6c0} /* (19, 9, 19) {real, imag} */,
  {32'h3f5494e2, 32'h3fc24b39} /* (19, 9, 18) {real, imag} */,
  {32'h3f96d2e5, 32'h3f6a7d44} /* (19, 9, 17) {real, imag} */,
  {32'hbe0420c0, 32'hbec4e470} /* (19, 9, 16) {real, imag} */,
  {32'hbf3e8c0b, 32'hbeedc9f0} /* (19, 9, 15) {real, imag} */,
  {32'h3eb290d2, 32'hbed3fd56} /* (19, 9, 14) {real, imag} */,
  {32'h3ee6a014, 32'h3ebf1730} /* (19, 9, 13) {real, imag} */,
  {32'h3ef85376, 32'h3f58cac0} /* (19, 9, 12) {real, imag} */,
  {32'h3ed1cf6c, 32'h3e46a950} /* (19, 9, 11) {real, imag} */,
  {32'h3f3552d8, 32'hbe1c6b00} /* (19, 9, 10) {real, imag} */,
  {32'h3fb567ef, 32'h3ef06a86} /* (19, 9, 9) {real, imag} */,
  {32'h3f5bb6e3, 32'hbe7d6ca0} /* (19, 9, 8) {real, imag} */,
  {32'h3dd9e7b8, 32'h3eb57b90} /* (19, 9, 7) {real, imag} */,
  {32'h3e85317c, 32'h3d473780} /* (19, 9, 6) {real, imag} */,
  {32'h3f3915bf, 32'hbf07670a} /* (19, 9, 5) {real, imag} */,
  {32'hbdf930b0, 32'hbe8c5d18} /* (19, 9, 4) {real, imag} */,
  {32'hbe648c38, 32'h3f0547e8} /* (19, 9, 3) {real, imag} */,
  {32'hbeee3a30, 32'h3cb48380} /* (19, 9, 2) {real, imag} */,
  {32'hbf5a9098, 32'hbf56945a} /* (19, 9, 1) {real, imag} */,
  {32'hbf0b710f, 32'hbe9ce8a0} /* (19, 9, 0) {real, imag} */,
  {32'hbf7893e6, 32'h3f1afcd4} /* (19, 8, 31) {real, imag} */,
  {32'hbf51ab84, 32'h3e9cdb88} /* (19, 8, 30) {real, imag} */,
  {32'h3f7b6bce, 32'hbf05d948} /* (19, 8, 29) {real, imag} */,
  {32'h3ed71b26, 32'hbf8ce4c2} /* (19, 8, 28) {real, imag} */,
  {32'hbeddf6e8, 32'h3e208e60} /* (19, 8, 27) {real, imag} */,
  {32'hbf3f7236, 32'h3e9a8330} /* (19, 8, 26) {real, imag} */,
  {32'hbe9bc580, 32'hbeb1f7b8} /* (19, 8, 25) {real, imag} */,
  {32'hbe761010, 32'hbebeee50} /* (19, 8, 24) {real, imag} */,
  {32'h3db41dd0, 32'hbf4f3938} /* (19, 8, 23) {real, imag} */,
  {32'h3f306fc0, 32'hbf8733de} /* (19, 8, 22) {real, imag} */,
  {32'h3f0da988, 32'hbda8b990} /* (19, 8, 21) {real, imag} */,
  {32'hbc6e0740, 32'hbd1afd00} /* (19, 8, 20) {real, imag} */,
  {32'hbf14bce9, 32'hbe9cd910} /* (19, 8, 19) {real, imag} */,
  {32'h3d54f9a0, 32'hbd15bcc0} /* (19, 8, 18) {real, imag} */,
  {32'h3f071d8d, 32'hbf039188} /* (19, 8, 17) {real, imag} */,
  {32'h3d92bb00, 32'hbf66f428} /* (19, 8, 16) {real, imag} */,
  {32'hbea1b10e, 32'hbe3529e0} /* (19, 8, 15) {real, imag} */,
  {32'h3d64bb80, 32'hbf0f0ec0} /* (19, 8, 14) {real, imag} */,
  {32'hbe7bf978, 32'hbed974f0} /* (19, 8, 13) {real, imag} */,
  {32'hbf10b5ee, 32'hbeb6e660} /* (19, 8, 12) {real, imag} */,
  {32'hbf4b1f86, 32'hbf258ac8} /* (19, 8, 11) {real, imag} */,
  {32'hbdeb0a18, 32'hbea63e72} /* (19, 8, 10) {real, imag} */,
  {32'h3e8a3a18, 32'h3e7f6968} /* (19, 8, 9) {real, imag} */,
  {32'hbcd14b40, 32'hbeb911a8} /* (19, 8, 8) {real, imag} */,
  {32'hbe7b1e38, 32'hbcc49900} /* (19, 8, 7) {real, imag} */,
  {32'hbc568f80, 32'h3ea66b40} /* (19, 8, 6) {real, imag} */,
  {32'h3e1893a0, 32'hbf012964} /* (19, 8, 5) {real, imag} */,
  {32'h3e1f6cbc, 32'hbee2b2d8} /* (19, 8, 4) {real, imag} */,
  {32'hbe5e91b0, 32'h3eeb9ea0} /* (19, 8, 3) {real, imag} */,
  {32'hbf061a92, 32'h3e99fe70} /* (19, 8, 2) {real, imag} */,
  {32'hbf1e401f, 32'hbed3bdc8} /* (19, 8, 1) {real, imag} */,
  {32'hbe659a78, 32'h3ba79500} /* (19, 8, 0) {real, imag} */,
  {32'hbe2abfdc, 32'h3f38d5b2} /* (19, 7, 31) {real, imag} */,
  {32'hbe4813a8, 32'h3e88d1dc} /* (19, 7, 30) {real, imag} */,
  {32'h3e17a20c, 32'h3ead3648} /* (19, 7, 29) {real, imag} */,
  {32'hbe418894, 32'hbf426764} /* (19, 7, 28) {real, imag} */,
  {32'hbde90858, 32'hbeb09a00} /* (19, 7, 27) {real, imag} */,
  {32'hbc009980, 32'hbe396fc0} /* (19, 7, 26) {real, imag} */,
  {32'h3c124a80, 32'h3e287c60} /* (19, 7, 25) {real, imag} */,
  {32'hbf50a65a, 32'h3fa337be} /* (19, 7, 24) {real, imag} */,
  {32'hbf468a4c, 32'hbdd2c9c0} /* (19, 7, 23) {real, imag} */,
  {32'h3e998598, 32'h3d32a320} /* (19, 7, 22) {real, imag} */,
  {32'h3f0447e9, 32'h3ec8fb5e} /* (19, 7, 21) {real, imag} */,
  {32'h3f89a928, 32'hbe963aa8} /* (19, 7, 20) {real, imag} */,
  {32'h3e515490, 32'h3e3f5ee8} /* (19, 7, 19) {real, imag} */,
  {32'hbe8581e4, 32'h3e2f0d70} /* (19, 7, 18) {real, imag} */,
  {32'h3e00b524, 32'hbd75cc80} /* (19, 7, 17) {real, imag} */,
  {32'hbf139d55, 32'hbdbf05e0} /* (19, 7, 16) {real, imag} */,
  {32'hbf1b75f2, 32'hbe8e1ea0} /* (19, 7, 15) {real, imag} */,
  {32'hbf6da79a, 32'hbeb99aa8} /* (19, 7, 14) {real, imag} */,
  {32'hbf01744c, 32'hbedf8d80} /* (19, 7, 13) {real, imag} */,
  {32'h3ef35ff2, 32'hbf709fb4} /* (19, 7, 12) {real, imag} */,
  {32'hbde0dc40, 32'hbf708de4} /* (19, 7, 11) {real, imag} */,
  {32'hbeeecbd0, 32'hbf94f7c8} /* (19, 7, 10) {real, imag} */,
  {32'hbf10a0b0, 32'hbf33a268} /* (19, 7, 9) {real, imag} */,
  {32'h3e9b867a, 32'h3e27add0} /* (19, 7, 8) {real, imag} */,
  {32'hbeb8f2e7, 32'h3f567652} /* (19, 7, 7) {real, imag} */,
  {32'hbf1d72f4, 32'h3f2f23ae} /* (19, 7, 6) {real, imag} */,
  {32'hbef506bc, 32'hbe0ab2e0} /* (19, 7, 5) {real, imag} */,
  {32'h3e759294, 32'hbe749c10} /* (19, 7, 4) {real, imag} */,
  {32'hbe8e3f24, 32'h3ee69690} /* (19, 7, 3) {real, imag} */,
  {32'hbe6ded90, 32'h3da52e00} /* (19, 7, 2) {real, imag} */,
  {32'h3e0f52d8, 32'hbeaab838} /* (19, 7, 1) {real, imag} */,
  {32'hbcccdcb0, 32'h3ef8aa18} /* (19, 7, 0) {real, imag} */,
  {32'hbf2bbdde, 32'hbcf89540} /* (19, 6, 31) {real, imag} */,
  {32'hbee5e5b8, 32'hbe46c1b0} /* (19, 6, 30) {real, imag} */,
  {32'hbf76f487, 32'h3e7cf620} /* (19, 6, 29) {real, imag} */,
  {32'hbfc57708, 32'h3e829758} /* (19, 6, 28) {real, imag} */,
  {32'hbf9640a2, 32'h3dcd3780} /* (19, 6, 27) {real, imag} */,
  {32'h3ed11f18, 32'h3df72380} /* (19, 6, 26) {real, imag} */,
  {32'h3f24bb54, 32'h3eeba8b8} /* (19, 6, 25) {real, imag} */,
  {32'hbf262344, 32'h3f95dbf2} /* (19, 6, 24) {real, imag} */,
  {32'hbf5406dc, 32'hbe3af4b0} /* (19, 6, 23) {real, imag} */,
  {32'h3ead9148, 32'hbdf49e70} /* (19, 6, 22) {real, imag} */,
  {32'h3fa0e386, 32'h3eb5bc6d} /* (19, 6, 21) {real, imag} */,
  {32'h3f95b15c, 32'h3d9a8090} /* (19, 6, 20) {real, imag} */,
  {32'hbcd89dc0, 32'hbe852ccc} /* (19, 6, 19) {real, imag} */,
  {32'h3d396d48, 32'hbea73b24} /* (19, 6, 18) {real, imag} */,
  {32'hbd1c9a58, 32'hbe409580} /* (19, 6, 17) {real, imag} */,
  {32'hbf53df21, 32'h3ed3b910} /* (19, 6, 16) {real, imag} */,
  {32'hbf01038c, 32'h3ef7b7d0} /* (19, 6, 15) {real, imag} */,
  {32'hbf2ccc31, 32'hbe51c340} /* (19, 6, 14) {real, imag} */,
  {32'hbefe24d0, 32'h3e1b59b0} /* (19, 6, 13) {real, imag} */,
  {32'h3f9b64cd, 32'hbe3c6bf0} /* (19, 6, 12) {real, imag} */,
  {32'h3f756b93, 32'h3f18be88} /* (19, 6, 11) {real, imag} */,
  {32'hbcf59100, 32'hbd3ac740} /* (19, 6, 10) {real, imag} */,
  {32'hbe446830, 32'h3e0c7230} /* (19, 6, 9) {real, imag} */,
  {32'hbebbeb68, 32'h3f3ba492} /* (19, 6, 8) {real, imag} */,
  {32'hbf8b7fdb, 32'h3f919041} /* (19, 6, 7) {real, imag} */,
  {32'hbf31967a, 32'h3f2efa9c} /* (19, 6, 6) {real, imag} */,
  {32'hbe601ff0, 32'hbf2215c8} /* (19, 6, 5) {real, imag} */,
  {32'hbf2ee0df, 32'hbec5dfe0} /* (19, 6, 4) {real, imag} */,
  {32'h3eeb2d02, 32'hbda93020} /* (19, 6, 3) {real, imag} */,
  {32'h3fcb9c4d, 32'hbe899d60} /* (19, 6, 2) {real, imag} */,
  {32'h3f900988, 32'hbf985a42} /* (19, 6, 1) {real, imag} */,
  {32'h3da5d2e8, 32'hbe972e6c} /* (19, 6, 0) {real, imag} */,
  {32'hbf978b34, 32'h3edb59b4} /* (19, 5, 31) {real, imag} */,
  {32'hbed212b8, 32'h3e90d34c} /* (19, 5, 30) {real, imag} */,
  {32'hbf1494c8, 32'hbe52e0b0} /* (19, 5, 29) {real, imag} */,
  {32'hbfa8dc4b, 32'hbddc8220} /* (19, 5, 28) {real, imag} */,
  {32'hbf482918, 32'h3f3e0420} /* (19, 5, 27) {real, imag} */,
  {32'h3f91690c, 32'h3d4db700} /* (19, 5, 26) {real, imag} */,
  {32'h3f692ee6, 32'h3ef60e60} /* (19, 5, 25) {real, imag} */,
  {32'hbe805e74, 32'h3f272cc0} /* (19, 5, 24) {real, imag} */,
  {32'hbe3fd3a8, 32'hbf1986ec} /* (19, 5, 23) {real, imag} */,
  {32'h3e848a78, 32'hbf3b86d4} /* (19, 5, 22) {real, imag} */,
  {32'h3f3b2749, 32'h3e68cd50} /* (19, 5, 21) {real, imag} */,
  {32'h3e2b0238, 32'h3d7d8600} /* (19, 5, 20) {real, imag} */,
  {32'hbf91aaa6, 32'hbe54fde8} /* (19, 5, 19) {real, imag} */,
  {32'hbeb6a6a6, 32'h3eeee3e2} /* (19, 5, 18) {real, imag} */,
  {32'hbe484420, 32'h3e854730} /* (19, 5, 17) {real, imag} */,
  {32'hbeca0381, 32'h3f5d70f5} /* (19, 5, 16) {real, imag} */,
  {32'hbd9802c8, 32'h3e77cda0} /* (19, 5, 15) {real, imag} */,
  {32'h3e8e7de0, 32'hbeba2a00} /* (19, 5, 14) {real, imag} */,
  {32'hbec275bc, 32'h3ed55db0} /* (19, 5, 13) {real, imag} */,
  {32'hbeb420f8, 32'hbd567100} /* (19, 5, 12) {real, imag} */,
  {32'h3f3dac9e, 32'h3e33ef40} /* (19, 5, 11) {real, imag} */,
  {32'h3ef3aaf8, 32'hbe616354} /* (19, 5, 10) {real, imag} */,
  {32'hbd8c4a64, 32'h3e159ff0} /* (19, 5, 9) {real, imag} */,
  {32'h3c0c1e40, 32'hbf08b43a} /* (19, 5, 8) {real, imag} */,
  {32'hbecb0edc, 32'hbe8a68aa} /* (19, 5, 7) {real, imag} */,
  {32'h3e1d008a, 32'hbf100f77} /* (19, 5, 6) {real, imag} */,
  {32'h3ee143b0, 32'h3d83ff80} /* (19, 5, 5) {real, imag} */,
  {32'h3ec40464, 32'h3ea51e30} /* (19, 5, 4) {real, imag} */,
  {32'h3ef2ffb4, 32'hbf0201c6} /* (19, 5, 3) {real, imag} */,
  {32'h3fcf92e3, 32'hbf325374} /* (19, 5, 2) {real, imag} */,
  {32'h3f4bbce8, 32'hbf83ec84} /* (19, 5, 1) {real, imag} */,
  {32'hbe82ee3d, 32'hbd43e680} /* (19, 5, 0) {real, imag} */,
  {32'hbf91f375, 32'h3e84df84} /* (19, 4, 31) {real, imag} */,
  {32'hbee4c450, 32'hbda683a0} /* (19, 4, 30) {real, imag} */,
  {32'hbe5617d8, 32'hbe7b01f0} /* (19, 4, 29) {real, imag} */,
  {32'hbf0d66a6, 32'h3d1e1380} /* (19, 4, 28) {real, imag} */,
  {32'hbf118eab, 32'hbe671080} /* (19, 4, 27) {real, imag} */,
  {32'h3e429910, 32'hbf2966b0} /* (19, 4, 26) {real, imag} */,
  {32'h3f143be2, 32'hbea43a08} /* (19, 4, 25) {real, imag} */,
  {32'h3f37b048, 32'h3ea888e8} /* (19, 4, 24) {real, imag} */,
  {32'h3eaab6f8, 32'hbea73ad8} /* (19, 4, 23) {real, imag} */,
  {32'hbf1ed2b1, 32'h3dc92a20} /* (19, 4, 22) {real, imag} */,
  {32'h3dedc628, 32'h3f96e647} /* (19, 4, 21) {real, imag} */,
  {32'h3f0e608b, 32'h3d8a1280} /* (19, 4, 20) {real, imag} */,
  {32'hbef6c60b, 32'hbec63418} /* (19, 4, 19) {real, imag} */,
  {32'hbeaf1eb3, 32'h3ee85a10} /* (19, 4, 18) {real, imag} */,
  {32'hbd4ccea8, 32'h3fa35848} /* (19, 4, 17) {real, imag} */,
  {32'hbe3f8bec, 32'h3fce0ead} /* (19, 4, 16) {real, imag} */,
  {32'h3ef4f1a2, 32'hbede8f20} /* (19, 4, 15) {real, imag} */,
  {32'h3f81d833, 32'hbf62f90e} /* (19, 4, 14) {real, imag} */,
  {32'hbe271048, 32'hbd430a40} /* (19, 4, 13) {real, imag} */,
  {32'hbe55cac8, 32'hbeb0c950} /* (19, 4, 12) {real, imag} */,
  {32'h3e8a7844, 32'hbe83b8a0} /* (19, 4, 11) {real, imag} */,
  {32'h3f2ad366, 32'hbe69d650} /* (19, 4, 10) {real, imag} */,
  {32'h3f9b9dc2, 32'hbf5fb50c} /* (19, 4, 9) {real, imag} */,
  {32'h3fd55504, 32'hbfc53aed} /* (19, 4, 8) {real, imag} */,
  {32'h3f66ad40, 32'hbec3fb28} /* (19, 4, 7) {real, imag} */,
  {32'h3f0a35aa, 32'h3e1aeca0} /* (19, 4, 6) {real, imag} */,
  {32'hbe704b70, 32'h3e9a6df7} /* (19, 4, 5) {real, imag} */,
  {32'h3ea6ce9e, 32'h3e3286f8} /* (19, 4, 4) {real, imag} */,
  {32'h3fb0a432, 32'hbca5b900} /* (19, 4, 3) {real, imag} */,
  {32'h3fa873ef, 32'hbe907438} /* (19, 4, 2) {real, imag} */,
  {32'h3f0cdbd7, 32'h3e0b2b10} /* (19, 4, 1) {real, imag} */,
  {32'hbe21ef60, 32'h3e9efd54} /* (19, 4, 0) {real, imag} */,
  {32'hbedaff8c, 32'hbef979a0} /* (19, 3, 31) {real, imag} */,
  {32'hbe0c16b0, 32'hbf337e04} /* (19, 3, 30) {real, imag} */,
  {32'hbe6c7914, 32'hbd4a7d80} /* (19, 3, 29) {real, imag} */,
  {32'hbf6eb755, 32'h3f3e39c8} /* (19, 3, 28) {real, imag} */,
  {32'hbfc43634, 32'h3e5b8ee0} /* (19, 3, 27) {real, imag} */,
  {32'hbf5c5cbe, 32'h3ec0f450} /* (19, 3, 26) {real, imag} */,
  {32'hbf214bac, 32'hbd0d9880} /* (19, 3, 25) {real, imag} */,
  {32'h3d7a7240, 32'h3ecf11c0} /* (19, 3, 24) {real, imag} */,
  {32'h3ce69460, 32'hbe171d40} /* (19, 3, 23) {real, imag} */,
  {32'hbdfd9ce0, 32'hbc5889c0} /* (19, 3, 22) {real, imag} */,
  {32'h3ef2bcbb, 32'h3ef5a488} /* (19, 3, 21) {real, imag} */,
  {32'h3d8d68a0, 32'hbe841cd0} /* (19, 3, 20) {real, imag} */,
  {32'h3e2b2270, 32'hbe5736b0} /* (19, 3, 19) {real, imag} */,
  {32'hbd859fe0, 32'hbf5fd0ce} /* (19, 3, 18) {real, imag} */,
  {32'hbc559880, 32'h3e0b0380} /* (19, 3, 17) {real, imag} */,
  {32'hbf28e226, 32'hbe7ffb80} /* (19, 3, 16) {real, imag} */,
  {32'hbea6a77d, 32'hbf90110b} /* (19, 3, 15) {real, imag} */,
  {32'h3f164f27, 32'hbfc78472} /* (19, 3, 14) {real, imag} */,
  {32'h3f6c8c4f, 32'hbfa82216} /* (19, 3, 13) {real, imag} */,
  {32'h3f8d4602, 32'hbfc62084} /* (19, 3, 12) {real, imag} */,
  {32'h3f8b8ec0, 32'hbf25d454} /* (19, 3, 11) {real, imag} */,
  {32'h3f9c8b5b, 32'hbd849660} /* (19, 3, 10) {real, imag} */,
  {32'h3fb0dabf, 32'hbfa744e4} /* (19, 3, 9) {real, imag} */,
  {32'h3f51bbfb, 32'hbfbd2d98} /* (19, 3, 8) {real, imag} */,
  {32'hbec2650d, 32'hbe661350} /* (19, 3, 7) {real, imag} */,
  {32'hbde8e9f8, 32'h3f0bf340} /* (19, 3, 6) {real, imag} */,
  {32'hbe6fc290, 32'h3d2638e0} /* (19, 3, 5) {real, imag} */,
  {32'h3e352088, 32'h3e2c13bc} /* (19, 3, 4) {real, imag} */,
  {32'h3f102f70, 32'h3dac9e00} /* (19, 3, 3) {real, imag} */,
  {32'h3e2c4160, 32'h3dbae180} /* (19, 3, 2) {real, imag} */,
  {32'hbe793c88, 32'h3e55dba0} /* (19, 3, 1) {real, imag} */,
  {32'hbdbb6490, 32'hbe900f10} /* (19, 3, 0) {real, imag} */,
  {32'hbe9d3118, 32'hbf918558} /* (19, 2, 31) {real, imag} */,
  {32'hbec687e0, 32'hbf7e1918} /* (19, 2, 30) {real, imag} */,
  {32'hbeb3c5e4, 32'hbdc1c860} /* (19, 2, 29) {real, imag} */,
  {32'hbd0eade0, 32'hbe8c8368} /* (19, 2, 28) {real, imag} */,
  {32'hbf51a895, 32'h3dd0b1c0} /* (19, 2, 27) {real, imag} */,
  {32'hbe1796f4, 32'h3f6b020c} /* (19, 2, 26) {real, imag} */,
  {32'hbe0b6368, 32'hbe80b4b0} /* (19, 2, 25) {real, imag} */,
  {32'hbf3895a4, 32'hbc1cf300} /* (19, 2, 24) {real, imag} */,
  {32'hbef0c7e0, 32'h3e5758bc} /* (19, 2, 23) {real, imag} */,
  {32'h3d87dec0, 32'hbf256496} /* (19, 2, 22) {real, imag} */,
  {32'h3f246efc, 32'hbf0befc8} /* (19, 2, 21) {real, imag} */,
  {32'hbdf7e920, 32'hbd327b00} /* (19, 2, 20) {real, imag} */,
  {32'h3f322976, 32'h3f39bd38} /* (19, 2, 19) {real, imag} */,
  {32'hbdd988e8, 32'hbe5a69f8} /* (19, 2, 18) {real, imag} */,
  {32'hbf1c1364, 32'hbed70848} /* (19, 2, 17) {real, imag} */,
  {32'h3e3ceb00, 32'hbf84370e} /* (19, 2, 16) {real, imag} */,
  {32'h3ecf0888, 32'hbfc7d622} /* (19, 2, 15) {real, imag} */,
  {32'hbcfe0890, 32'hbfdfc1da} /* (19, 2, 14) {real, imag} */,
  {32'hbc11ebc0, 32'hbf4b0a26} /* (19, 2, 13) {real, imag} */,
  {32'h3e465fe0, 32'hbf594458} /* (19, 2, 12) {real, imag} */,
  {32'h3f60c146, 32'hbf2832dc} /* (19, 2, 11) {real, imag} */,
  {32'h3edf0ada, 32'hbf5fb9d8} /* (19, 2, 10) {real, imag} */,
  {32'h3e234950, 32'hbfd92ed0} /* (19, 2, 9) {real, imag} */,
  {32'hbec4f496, 32'hbfafbde4} /* (19, 2, 8) {real, imag} */,
  {32'hbdf8e920, 32'hbee8c7e0} /* (19, 2, 7) {real, imag} */,
  {32'h3ea742ba, 32'h3fa815bc} /* (19, 2, 6) {real, imag} */,
  {32'hbce2a200, 32'h3f7fdbb6} /* (19, 2, 5) {real, imag} */,
  {32'h3ed86b56, 32'hbdf989c0} /* (19, 2, 4) {real, imag} */,
  {32'h3e7f8fb8, 32'h3edae120} /* (19, 2, 3) {real, imag} */,
  {32'h3edbce08, 32'h3f8b8e33} /* (19, 2, 2) {real, imag} */,
  {32'h3f2f5ad2, 32'h3f420fac} /* (19, 2, 1) {real, imag} */,
  {32'h3e1aa728, 32'hbf028624} /* (19, 2, 0) {real, imag} */,
  {32'h3d1f49a0, 32'hbf3dd3f8} /* (19, 1, 31) {real, imag} */,
  {32'h3eb6b0e2, 32'hbf9c084e} /* (19, 1, 30) {real, imag} */,
  {32'h3f2b2f3b, 32'h3c626300} /* (19, 1, 29) {real, imag} */,
  {32'h3ecbd0b1, 32'hbf112b34} /* (19, 1, 28) {real, imag} */,
  {32'hbf3e8e88, 32'hbe6ded80} /* (19, 1, 27) {real, imag} */,
  {32'hbf7dd1b2, 32'h3f06cfb8} /* (19, 1, 26) {real, imag} */,
  {32'hbec8b594, 32'hbe5d8860} /* (19, 1, 25) {real, imag} */,
  {32'hbc366200, 32'hbf0d3d60} /* (19, 1, 24) {real, imag} */,
  {32'h3f1a21d0, 32'h3f6846fe} /* (19, 1, 23) {real, imag} */,
  {32'h3f346400, 32'h3f068f48} /* (19, 1, 22) {real, imag} */,
  {32'h3f3daf1e, 32'hbecb6160} /* (19, 1, 21) {real, imag} */,
  {32'h3e6ed478, 32'hbeaa2f28} /* (19, 1, 20) {real, imag} */,
  {32'h3f2edb2a, 32'h3eafae98} /* (19, 1, 19) {real, imag} */,
  {32'hbe24f750, 32'hbde51760} /* (19, 1, 18) {real, imag} */,
  {32'hbf80bdff, 32'hbe81bec0} /* (19, 1, 17) {real, imag} */,
  {32'hbd193d80, 32'hbf544eb6} /* (19, 1, 16) {real, imag} */,
  {32'h3e12a718, 32'hbf9034fe} /* (19, 1, 15) {real, imag} */,
  {32'hbf429d45, 32'hbf65a7a4} /* (19, 1, 14) {real, imag} */,
  {32'hbfc4dedd, 32'hbed9b4d8} /* (19, 1, 13) {real, imag} */,
  {32'hbf591555, 32'h3e70a870} /* (19, 1, 12) {real, imag} */,
  {32'h3dc977d0, 32'h3ed66f00} /* (19, 1, 11) {real, imag} */,
  {32'h3e8f8c18, 32'hbef5b998} /* (19, 1, 10) {real, imag} */,
  {32'h3e40f620, 32'hbf441008} /* (19, 1, 9) {real, imag} */,
  {32'hbe02e360, 32'h3eecfb38} /* (19, 1, 8) {real, imag} */,
  {32'h3f416bda, 32'hbe427710} /* (19, 1, 7) {real, imag} */,
  {32'h3efd76dc, 32'hbdda7440} /* (19, 1, 6) {real, imag} */,
  {32'hbf6c11d3, 32'h3f25ab40} /* (19, 1, 5) {real, imag} */,
  {32'h3d6c5860, 32'h3dd05d40} /* (19, 1, 4) {real, imag} */,
  {32'h3f4eccec, 32'hbe21bf10} /* (19, 1, 3) {real, imag} */,
  {32'h3f51d546, 32'h3e7fbff0} /* (19, 1, 2) {real, imag} */,
  {32'h3f3b23ce, 32'h3efaf10c} /* (19, 1, 1) {real, imag} */,
  {32'h3e2eaff2, 32'hbd849da0} /* (19, 1, 0) {real, imag} */,
  {32'h3d41f408, 32'h3d679090} /* (19, 0, 31) {real, imag} */,
  {32'h3ef2597c, 32'hbec07288} /* (19, 0, 30) {real, imag} */,
  {32'h3edb83af, 32'h3e8d00dc} /* (19, 0, 29) {real, imag} */,
  {32'h3d1055a0, 32'h3ef076dc} /* (19, 0, 28) {real, imag} */,
  {32'hbf491476, 32'h3f34f092} /* (19, 0, 27) {real, imag} */,
  {32'hbf4ab3af, 32'h3f2e4e5e} /* (19, 0, 26) {real, imag} */,
  {32'hbea9fe6e, 32'h3f1ab484} /* (19, 0, 25) {real, imag} */,
  {32'h3f07c6b0, 32'h3efc9818} /* (19, 0, 24) {real, imag} */,
  {32'h3f9cc678, 32'h3f185a0d} /* (19, 0, 23) {real, imag} */,
  {32'h3f92fb65, 32'h3f153080} /* (19, 0, 22) {real, imag} */,
  {32'h3ea4e284, 32'h3e495eb8} /* (19, 0, 21) {real, imag} */,
  {32'hbe062a80, 32'hbdbf24b4} /* (19, 0, 20) {real, imag} */,
  {32'h3cd995e0, 32'h3e867134} /* (19, 0, 19) {real, imag} */,
  {32'h3e7e1bdc, 32'hbe6a1e00} /* (19, 0, 18) {real, imag} */,
  {32'h3d0ba230, 32'hbdc23280} /* (19, 0, 17) {real, imag} */,
  {32'h3bd19100, 32'hbeca805e} /* (19, 0, 16) {real, imag} */,
  {32'h3cb30540, 32'hbed34720} /* (19, 0, 15) {real, imag} */,
  {32'hbf35e58a, 32'hbd08b180} /* (19, 0, 14) {real, imag} */,
  {32'hbf86d84a, 32'h3ddf4cc0} /* (19, 0, 13) {real, imag} */,
  {32'h3e190690, 32'h3ec83788} /* (19, 0, 12) {real, imag} */,
  {32'h3d7378e0, 32'h3e6e6b60} /* (19, 0, 11) {real, imag} */,
  {32'h3b116980, 32'h3d0aa398} /* (19, 0, 10) {real, imag} */,
  {32'hbd2e5060, 32'h3e6205c8} /* (19, 0, 9) {real, imag} */,
  {32'h3e98c5f0, 32'h3f2bd6fc} /* (19, 0, 8) {real, imag} */,
  {32'h3f0c7e2e, 32'hbe5957d0} /* (19, 0, 7) {real, imag} */,
  {32'h3ecddb4c, 32'hbf486f2d} /* (19, 0, 6) {real, imag} */,
  {32'hbeb1248c, 32'h3ece2e21} /* (19, 0, 5) {real, imag} */,
  {32'hbe118cdf, 32'h3f50e20c} /* (19, 0, 4) {real, imag} */,
  {32'h3f43a64e, 32'hbe235460} /* (19, 0, 3) {real, imag} */,
  {32'h3eb1a8cd, 32'hbe10d4b8} /* (19, 0, 2) {real, imag} */,
  {32'hbcc7bf30, 32'h3ec63724} /* (19, 0, 1) {real, imag} */,
  {32'hbec86414, 32'h3f0c8208} /* (19, 0, 0) {real, imag} */,
  {32'hbe358a0c, 32'hbd08aae0} /* (18, 31, 31) {real, imag} */,
  {32'hbf2f9e5d, 32'hbf0116d8} /* (18, 31, 30) {real, imag} */,
  {32'hbf3f4cd3, 32'hbe467100} /* (18, 31, 29) {real, imag} */,
  {32'hbf1d620c, 32'hbda4d400} /* (18, 31, 28) {real, imag} */,
  {32'hbe903168, 32'hbe269f40} /* (18, 31, 27) {real, imag} */,
  {32'hbe446cc8, 32'h3e036ea0} /* (18, 31, 26) {real, imag} */,
  {32'h3e3aadc8, 32'h3e6d8040} /* (18, 31, 25) {real, imag} */,
  {32'h3ed1fd04, 32'h3e597fe0} /* (18, 31, 24) {real, imag} */,
  {32'hbe473990, 32'hbeceb5b8} /* (18, 31, 23) {real, imag} */,
  {32'hbe146f98, 32'hbe9b1a80} /* (18, 31, 22) {real, imag} */,
  {32'h3f1aa943, 32'h3d0ddf00} /* (18, 31, 21) {real, imag} */,
  {32'h3f50012e, 32'hbf030cf0} /* (18, 31, 20) {real, imag} */,
  {32'hbd1c50e0, 32'hbe871450} /* (18, 31, 19) {real, imag} */,
  {32'hbeb44aa5, 32'h3e3837d0} /* (18, 31, 18) {real, imag} */,
  {32'h3e436452, 32'h3e46ec20} /* (18, 31, 17) {real, imag} */,
  {32'h3e99f1f7, 32'h3e078800} /* (18, 31, 16) {real, imag} */,
  {32'h3eeabdea, 32'h3e8394b0} /* (18, 31, 15) {real, imag} */,
  {32'h3f242754, 32'h3f13ba30} /* (18, 31, 14) {real, imag} */,
  {32'h3e9e68b8, 32'h3e52adc0} /* (18, 31, 13) {real, imag} */,
  {32'hbefa6fa0, 32'h3ec8d2b8} /* (18, 31, 12) {real, imag} */,
  {32'hbe7ec214, 32'h3f869c74} /* (18, 31, 11) {real, imag} */,
  {32'h3e82fd64, 32'h3e362d14} /* (18, 31, 10) {real, imag} */,
  {32'hbee8c7d0, 32'hbedf0800} /* (18, 31, 9) {real, imag} */,
  {32'hbf300884, 32'h3e6eeb40} /* (18, 31, 8) {real, imag} */,
  {32'hbeb20770, 32'h3ef7e6b8} /* (18, 31, 7) {real, imag} */,
  {32'hbf13de40, 32'hbdf5a9c0} /* (18, 31, 6) {real, imag} */,
  {32'hbf3a0baa, 32'hbe911f60} /* (18, 31, 5) {real, imag} */,
  {32'hbf07379e, 32'hbec789c8} /* (18, 31, 4) {real, imag} */,
  {32'hbf7b3ca5, 32'hbf205648} /* (18, 31, 3) {real, imag} */,
  {32'hbecd5432, 32'hbf056da8} /* (18, 31, 2) {real, imag} */,
  {32'hbf0a681d, 32'h3dea9c40} /* (18, 31, 1) {real, imag} */,
  {32'hbe94894c, 32'h3cdd5180} /* (18, 31, 0) {real, imag} */,
  {32'hbf4baa78, 32'h3f386958} /* (18, 30, 31) {real, imag} */,
  {32'hbf85ddc2, 32'h3f87dab0} /* (18, 30, 30) {real, imag} */,
  {32'hbef999c0, 32'h3f1fdee8} /* (18, 30, 29) {real, imag} */,
  {32'hbf5f1614, 32'h3e5b2e60} /* (18, 30, 28) {real, imag} */,
  {32'hbf7ca7f0, 32'h3e6024c0} /* (18, 30, 27) {real, imag} */,
  {32'hbedcb0d2, 32'h3e9a97a0} /* (18, 30, 26) {real, imag} */,
  {32'h3cf44b20, 32'h3d468300} /* (18, 30, 25) {real, imag} */,
  {32'h3e7071c4, 32'h3f205e40} /* (18, 30, 24) {real, imag} */,
  {32'h3cceeb60, 32'hbeae55e0} /* (18, 30, 23) {real, imag} */,
  {32'hbec3c5fc, 32'hbefc65d0} /* (18, 30, 22) {real, imag} */,
  {32'h3ec984f4, 32'h3efa0248} /* (18, 30, 21) {real, imag} */,
  {32'h3f26b704, 32'h3e96f608} /* (18, 30, 20) {real, imag} */,
  {32'h3e9c46f8, 32'hbeae07b0} /* (18, 30, 19) {real, imag} */,
  {32'hbe54dda0, 32'hbcfa1800} /* (18, 30, 18) {real, imag} */,
  {32'h3ea9002f, 32'h3cbe4b00} /* (18, 30, 17) {real, imag} */,
  {32'h3ecd97e8, 32'hbb0bd800} /* (18, 30, 16) {real, imag} */,
  {32'h3eb7686c, 32'h3ea66180} /* (18, 30, 15) {real, imag} */,
  {32'h3f1b2c1e, 32'h3f7686f0} /* (18, 30, 14) {real, imag} */,
  {32'hbd994540, 32'h3e789b80} /* (18, 30, 13) {real, imag} */,
  {32'hbf2e6ee7, 32'h3e376700} /* (18, 30, 12) {real, imag} */,
  {32'h3e6f1e00, 32'h3f67eeb8} /* (18, 30, 11) {real, imag} */,
  {32'h3efa75e8, 32'h3ed72340} /* (18, 30, 10) {real, imag} */,
  {32'hbea7fcf6, 32'hbf6b5ff0} /* (18, 30, 9) {real, imag} */,
  {32'hbefb0bf4, 32'h3ebf52a0} /* (18, 30, 8) {real, imag} */,
  {32'hbce50e00, 32'h3f567b58} /* (18, 30, 7) {real, imag} */,
  {32'hbf372e8a, 32'hbee43ae0} /* (18, 30, 6) {real, imag} */,
  {32'hbf6832c0, 32'hbe8f95a0} /* (18, 30, 5) {real, imag} */,
  {32'hbecba320, 32'hbd8e8700} /* (18, 30, 4) {real, imag} */,
  {32'hbe15b9e0, 32'hbf086080} /* (18, 30, 3) {real, imag} */,
  {32'hbf13de94, 32'hbea97780} /* (18, 30, 2) {real, imag} */,
  {32'hbf28ba0d, 32'h3e85ec40} /* (18, 30, 1) {real, imag} */,
  {32'hbd39f060, 32'h3f13b710} /* (18, 30, 0) {real, imag} */,
  {32'hbf6d4d08, 32'hbdcf0380} /* (18, 29, 31) {real, imag} */,
  {32'hbf1dcd28, 32'h3e510540} /* (18, 29, 30) {real, imag} */,
  {32'h3f1be1f4, 32'h3e48b480} /* (18, 29, 29) {real, imag} */,
  {32'h3c189500, 32'h3ed5fd40} /* (18, 29, 28) {real, imag} */,
  {32'hbf943470, 32'h3ef57690} /* (18, 29, 27) {real, imag} */,
  {32'hbfb8a09a, 32'h3f1df280} /* (18, 29, 26) {real, imag} */,
  {32'hbf54470b, 32'h3d864f00} /* (18, 29, 25) {real, imag} */,
  {32'hbf2b19c4, 32'h3e2a4200} /* (18, 29, 24) {real, imag} */,
  {32'hbef70fc0, 32'hbf2dc5f0} /* (18, 29, 23) {real, imag} */,
  {32'hbe8d0ca8, 32'hbed9e330} /* (18, 29, 22) {real, imag} */,
  {32'hbe3980be, 32'h3e8723fc} /* (18, 29, 21) {real, imag} */,
  {32'h3d9f46c0, 32'h3e62ea80} /* (18, 29, 20) {real, imag} */,
  {32'h3dbdd4d0, 32'hbf229070} /* (18, 29, 19) {real, imag} */,
  {32'h3f69cca2, 32'h3eb40ce0} /* (18, 29, 18) {real, imag} */,
  {32'h3f0e9734, 32'h3eb61b60} /* (18, 29, 17) {real, imag} */,
  {32'hbd3811c0, 32'hbf17dbd0} /* (18, 29, 16) {real, imag} */,
  {32'hbe11c030, 32'h3e887a30} /* (18, 29, 15) {real, imag} */,
  {32'h3e228f00, 32'h3f946e68} /* (18, 29, 14) {real, imag} */,
  {32'hbd014000, 32'h3f384ec0} /* (18, 29, 13) {real, imag} */,
  {32'hbe2ffea0, 32'h3ef1b950} /* (18, 29, 12) {real, imag} */,
  {32'h3f744746, 32'hbe8432e0} /* (18, 29, 11) {real, imag} */,
  {32'h3e915638, 32'hbe478da0} /* (18, 29, 10) {real, imag} */,
  {32'hbf0f99b2, 32'hbfaa4a30} /* (18, 29, 9) {real, imag} */,
  {32'hbebe4850, 32'hbebf9000} /* (18, 29, 8) {real, imag} */,
  {32'hbec26d78, 32'h3f20c6d0} /* (18, 29, 7) {real, imag} */,
  {32'hbf1f6d84, 32'hbdf46f00} /* (18, 29, 6) {real, imag} */,
  {32'hbe38b720, 32'hbec853b0} /* (18, 29, 5) {real, imag} */,
  {32'h3e4e9540, 32'hbed5fec0} /* (18, 29, 4) {real, imag} */,
  {32'h3f40c99c, 32'hbe2ad0a0} /* (18, 29, 3) {real, imag} */,
  {32'hbf043c88, 32'h3dba1000} /* (18, 29, 2) {real, imag} */,
  {32'hbef6d81e, 32'h3e92c460} /* (18, 29, 1) {real, imag} */,
  {32'hbc52a300, 32'h3f31611c} /* (18, 29, 0) {real, imag} */,
  {32'hbe772718, 32'hbf0b3fa4} /* (18, 28, 31) {real, imag} */,
  {32'h3e3f6fc8, 32'hbf1aa380} /* (18, 28, 30) {real, imag} */,
  {32'h3fbbb5dd, 32'h3e6f5d00} /* (18, 28, 29) {real, imag} */,
  {32'h3c97d580, 32'h3f139f68} /* (18, 28, 28) {real, imag} */,
  {32'hbf846fa2, 32'hbd0f2700} /* (18, 28, 27) {real, imag} */,
  {32'hbf87b06c, 32'h3eacec40} /* (18, 28, 26) {real, imag} */,
  {32'hbf876313, 32'hbc51b600} /* (18, 28, 25) {real, imag} */,
  {32'hbf463950, 32'h3e755280} /* (18, 28, 24) {real, imag} */,
  {32'hbf6c9630, 32'hbedfb880} /* (18, 28, 23) {real, imag} */,
  {32'hbee909fc, 32'hbeebe400} /* (18, 28, 22) {real, imag} */,
  {32'hbf11abc0, 32'hbf17f630} /* (18, 28, 21) {real, imag} */,
  {32'hbde410e0, 32'hbda1f680} /* (18, 28, 20) {real, imag} */,
  {32'hbe2d2a80, 32'hbedaf6e0} /* (18, 28, 19) {real, imag} */,
  {32'h3f3f3560, 32'hbe90e280} /* (18, 28, 18) {real, imag} */,
  {32'hbea8acbc, 32'hbd81b180} /* (18, 28, 17) {real, imag} */,
  {32'hbec96038, 32'hbee211e0} /* (18, 28, 16) {real, imag} */,
  {32'h3e8b3be0, 32'hbcde4c00} /* (18, 28, 15) {real, imag} */,
  {32'h3f558260, 32'h3f035230} /* (18, 28, 14) {real, imag} */,
  {32'h3f2a7018, 32'h3f0f9c50} /* (18, 28, 13) {real, imag} */,
  {32'h3f41438e, 32'h3ed5d160} /* (18, 28, 12) {real, imag} */,
  {32'h3e9b200c, 32'hbf0615e0} /* (18, 28, 11) {real, imag} */,
  {32'hbe296380, 32'hbee7b0a8} /* (18, 28, 10) {real, imag} */,
  {32'hbedb2764, 32'hbea5c940} /* (18, 28, 9) {real, imag} */,
  {32'hbf781a5c, 32'hbe4fc8e0} /* (18, 28, 8) {real, imag} */,
  {32'hbf1ed412, 32'h3e80ad40} /* (18, 28, 7) {real, imag} */,
  {32'hbf379b86, 32'h3ee89100} /* (18, 28, 6) {real, imag} */,
  {32'hbf01b6dc, 32'hbd87b280} /* (18, 28, 5) {real, imag} */,
  {32'hbddaecc0, 32'h3f251810} /* (18, 28, 4) {real, imag} */,
  {32'h3cb17e80, 32'hbe7dd540} /* (18, 28, 3) {real, imag} */,
  {32'hbed377b0, 32'hbe2f4d80} /* (18, 28, 2) {real, imag} */,
  {32'hbf053aa5, 32'h3e60e080} /* (18, 28, 1) {real, imag} */,
  {32'hbeed5626, 32'h3d87bc80} /* (18, 28, 0) {real, imag} */,
  {32'h3e339fa0, 32'hbede6670} /* (18, 27, 31) {real, imag} */,
  {32'h3eeea1c4, 32'hbedb2c10} /* (18, 27, 30) {real, imag} */,
  {32'h3f9b10e8, 32'hbd30f600} /* (18, 27, 29) {real, imag} */,
  {32'hbf78b712, 32'h3f3fec90} /* (18, 27, 28) {real, imag} */,
  {32'hc01045e8, 32'h3e86eda0} /* (18, 27, 27) {real, imag} */,
  {32'hbfaa7cea, 32'hbec8a5c0} /* (18, 27, 26) {real, imag} */,
  {32'hbf42fa6e, 32'hbfa5b754} /* (18, 27, 25) {real, imag} */,
  {32'hbf669a68, 32'hbf3e68d0} /* (18, 27, 24) {real, imag} */,
  {32'hbf2e8368, 32'hbfc2a2b8} /* (18, 27, 23) {real, imag} */,
  {32'hbf433664, 32'hbf808da0} /* (18, 27, 22) {real, imag} */,
  {32'hbf4f9972, 32'hbd83be80} /* (18, 27, 21) {real, imag} */,
  {32'hbe9c64a8, 32'h3da7a340} /* (18, 27, 20) {real, imag} */,
  {32'h3d8c57a0, 32'h3c441200} /* (18, 27, 19) {real, imag} */,
  {32'h3f307cb4, 32'hbe9cc420} /* (18, 27, 18) {real, imag} */,
  {32'h3ee57928, 32'hbea14180} /* (18, 27, 17) {real, imag} */,
  {32'h3e7c36e0, 32'hbf1fcc50} /* (18, 27, 16) {real, imag} */,
  {32'h3f890d75, 32'hbea99440} /* (18, 27, 15) {real, imag} */,
  {32'h3f3cefd0, 32'hbf0c47c8} /* (18, 27, 14) {real, imag} */,
  {32'h3cb8df00, 32'h3da161c0} /* (18, 27, 13) {real, imag} */,
  {32'hbebd18a0, 32'hbdb72f80} /* (18, 27, 12) {real, imag} */,
  {32'hbf927a27, 32'hbf293040} /* (18, 27, 11) {real, imag} */,
  {32'hbf4e3be2, 32'hbe81e178} /* (18, 27, 10) {real, imag} */,
  {32'hbe0bf188, 32'h3f36a760} /* (18, 27, 9) {real, imag} */,
  {32'hbe5e3fec, 32'h3ea2ad80} /* (18, 27, 8) {real, imag} */,
  {32'hbe9b1970, 32'h3d607600} /* (18, 27, 7) {real, imag} */,
  {32'hbead4ca4, 32'h3dc75f80} /* (18, 27, 6) {real, imag} */,
  {32'hbec11b48, 32'h3f045bd0} /* (18, 27, 5) {real, imag} */,
  {32'hbec7dc58, 32'h3ec91b30} /* (18, 27, 4) {real, imag} */,
  {32'hbf29f0d7, 32'hbe97da70} /* (18, 27, 3) {real, imag} */,
  {32'hbed633c8, 32'h3ed48640} /* (18, 27, 2) {real, imag} */,
  {32'hbe5898a0, 32'h3edec670} /* (18, 27, 1) {real, imag} */,
  {32'hbf3b0f04, 32'h3d040100} /* (18, 27, 0) {real, imag} */,
  {32'hbebd6768, 32'hbed1db30} /* (18, 26, 31) {real, imag} */,
  {32'hbe988694, 32'hbf5be578} /* (18, 26, 30) {real, imag} */,
  {32'h3e4bd520, 32'hbf855058} /* (18, 26, 29) {real, imag} */,
  {32'hbedcb8ee, 32'hbd32c400} /* (18, 26, 28) {real, imag} */,
  {32'hbfa19bf7, 32'hbed5b4b0} /* (18, 26, 27) {real, imag} */,
  {32'hbf838169, 32'hbf829c28} /* (18, 26, 26) {real, imag} */,
  {32'hbf1f44a4, 32'hbf07bfa0} /* (18, 26, 25) {real, imag} */,
  {32'hbf06bfa8, 32'hbf4eaaa0} /* (18, 26, 24) {real, imag} */,
  {32'hbf0a795a, 32'hbf75ff80} /* (18, 26, 23) {real, imag} */,
  {32'hbe83d7cc, 32'hbd6ba480} /* (18, 26, 22) {real, imag} */,
  {32'h3e5e8cec, 32'h3e9d7260} /* (18, 26, 21) {real, imag} */,
  {32'h3f3e914c, 32'hbc9f6b00} /* (18, 26, 20) {real, imag} */,
  {32'h3f613b2a, 32'h3e513900} /* (18, 26, 19) {real, imag} */,
  {32'h3fd8bf16, 32'h3f3464a8} /* (18, 26, 18) {real, imag} */,
  {32'h3f9d18d0, 32'h3e9f3780} /* (18, 26, 17) {real, imag} */,
  {32'h3ee5c098, 32'hbf11feb0} /* (18, 26, 16) {real, imag} */,
  {32'h3f2f5d5c, 32'h3ee34e60} /* (18, 26, 15) {real, imag} */,
  {32'h3ed42908, 32'hbed6e240} /* (18, 26, 14) {real, imag} */,
  {32'h3dd7eff0, 32'hbdc6e640} /* (18, 26, 13) {real, imag} */,
  {32'h3de54c20, 32'hbe7a06a0} /* (18, 26, 12) {real, imag} */,
  {32'h3d8ae950, 32'hbf500c78} /* (18, 26, 11) {real, imag} */,
  {32'hbe7e42e4, 32'hbea62ed8} /* (18, 26, 10) {real, imag} */,
  {32'hbefc32f4, 32'hbbd95000} /* (18, 26, 9) {real, imag} */,
  {32'hbecbf860, 32'h3d78cc00} /* (18, 26, 8) {real, imag} */,
  {32'hbf6d3394, 32'hbe9a1ba0} /* (18, 26, 7) {real, imag} */,
  {32'hbe301f70, 32'h3bf6f400} /* (18, 26, 6) {real, imag} */,
  {32'hbd6939c0, 32'hbe042580} /* (18, 26, 5) {real, imag} */,
  {32'h3e3e21a0, 32'hbe8a76e0} /* (18, 26, 4) {real, imag} */,
  {32'h3d996948, 32'h3d67f480} /* (18, 26, 3) {real, imag} */,
  {32'hbf1d2006, 32'h3f0c6b70} /* (18, 26, 2) {real, imag} */,
  {32'h3e0af280, 32'h3e62a2c0} /* (18, 26, 1) {real, imag} */,
  {32'h3dae1960, 32'hbdec6880} /* (18, 26, 0) {real, imag} */,
  {32'hbe991058, 32'hba8d1800} /* (18, 25, 31) {real, imag} */,
  {32'h3d94f560, 32'hbf3df430} /* (18, 25, 30) {real, imag} */,
  {32'h3cd854a0, 32'hbf4ad790} /* (18, 25, 29) {real, imag} */,
  {32'h3e03c380, 32'hbe1c9340} /* (18, 25, 28) {real, imag} */,
  {32'hbedcb2ea, 32'hbea2d0f0} /* (18, 25, 27) {real, imag} */,
  {32'hbf1dc185, 32'hbf934e80} /* (18, 25, 26) {real, imag} */,
  {32'hbee5cb6e, 32'hbdf20980} /* (18, 25, 25) {real, imag} */,
  {32'hbe9f9150, 32'hbefa6540} /* (18, 25, 24) {real, imag} */,
  {32'hbe0212a0, 32'hbe88d220} /* (18, 25, 23) {real, imag} */,
  {32'hbeeb6984, 32'h3f08f250} /* (18, 25, 22) {real, imag} */,
  {32'hbdd40a1c, 32'h3e4c54a0} /* (18, 25, 21) {real, imag} */,
  {32'h3ee31a68, 32'hbec35e10} /* (18, 25, 20) {real, imag} */,
  {32'h3f4b43a0, 32'h3e31f980} /* (18, 25, 19) {real, imag} */,
  {32'h3f9b762f, 32'h3f80d1e8} /* (18, 25, 18) {real, imag} */,
  {32'h3f0cefca, 32'h3f354270} /* (18, 25, 17) {real, imag} */,
  {32'h3f147ed6, 32'h3c147800} /* (18, 25, 16) {real, imag} */,
  {32'h3f5c8c44, 32'h3f636ca0} /* (18, 25, 15) {real, imag} */,
  {32'h3f73b650, 32'h3f17a680} /* (18, 25, 14) {real, imag} */,
  {32'h3fa4080e, 32'h3ec9b2c0} /* (18, 25, 13) {real, imag} */,
  {32'h3f3cef6e, 32'h3ee50d20} /* (18, 25, 12) {real, imag} */,
  {32'h3e36b700, 32'hbccced00} /* (18, 25, 11) {real, imag} */,
  {32'hbf2fc462, 32'hbe26ad40} /* (18, 25, 10) {real, imag} */,
  {32'hbf7233f0, 32'hbf94571c} /* (18, 25, 9) {real, imag} */,
  {32'hbf3be3f8, 32'hbf0b9590} /* (18, 25, 8) {real, imag} */,
  {32'hbf758a22, 32'hbe929f10} /* (18, 25, 7) {real, imag} */,
  {32'hbe9131ec, 32'h3f155b88} /* (18, 25, 6) {real, imag} */,
  {32'hbe527520, 32'h3eb8bf80} /* (18, 25, 5) {real, imag} */,
  {32'h3e34a360, 32'hbf13daf0} /* (18, 25, 4) {real, imag} */,
  {32'hbdb57af0, 32'hbf279680} /* (18, 25, 3) {real, imag} */,
  {32'hbf822aa3, 32'hbecd3a20} /* (18, 25, 2) {real, imag} */,
  {32'hbf0fdb54, 32'hbe159ce0} /* (18, 25, 1) {real, imag} */,
  {32'hbe9a4fe4, 32'h3de4d2a0} /* (18, 25, 0) {real, imag} */,
  {32'h3d420940, 32'h3d0c6300} /* (18, 24, 31) {real, imag} */,
  {32'h3ef9c928, 32'hbe4f4140} /* (18, 24, 30) {real, imag} */,
  {32'hbe7781d0, 32'h3ee6f8c0} /* (18, 24, 29) {real, imag} */,
  {32'hbf121cd6, 32'h3dc8af00} /* (18, 24, 28) {real, imag} */,
  {32'hbf9d2b98, 32'hbe0b2e20} /* (18, 24, 27) {real, imag} */,
  {32'hbf8148fc, 32'hbeb46e60} /* (18, 24, 26) {real, imag} */,
  {32'hbf1ae8ce, 32'h3dd79200} /* (18, 24, 25) {real, imag} */,
  {32'hbf2ad64e, 32'hbf048510} /* (18, 24, 24) {real, imag} */,
  {32'h3d69d480, 32'hbfa15ed0} /* (18, 24, 23) {real, imag} */,
  {32'hbf2eea88, 32'hbc5df400} /* (18, 24, 22) {real, imag} */,
  {32'hbf259117, 32'hbd32d240} /* (18, 24, 21) {real, imag} */,
  {32'hbf3618d4, 32'hbdccb400} /* (18, 24, 20) {real, imag} */,
  {32'h3f0915fc, 32'h3f4e6970} /* (18, 24, 19) {real, imag} */,
  {32'h3f3931c2, 32'h3fc7f178} /* (18, 24, 18) {real, imag} */,
  {32'h3f64ed9e, 32'h3f010118} /* (18, 24, 17) {real, imag} */,
  {32'h3f5e62a3, 32'h3c8aa600} /* (18, 24, 16) {real, imag} */,
  {32'hbdb092a0, 32'h3e51a780} /* (18, 24, 15) {real, imag} */,
  {32'h3f10102a, 32'h3f1bed10} /* (18, 24, 14) {real, imag} */,
  {32'h3f3e7a9a, 32'h3ef2d900} /* (18, 24, 13) {real, imag} */,
  {32'h3f833c18, 32'h3f748580} /* (18, 24, 12) {real, imag} */,
  {32'h3e6990d0, 32'h3ed9b9b0} /* (18, 24, 11) {real, imag} */,
  {32'hbf40db78, 32'hbed59ff8} /* (18, 24, 10) {real, imag} */,
  {32'hbf1f23b4, 32'hbf5327d0} /* (18, 24, 9) {real, imag} */,
  {32'h3efaa124, 32'hbf2d4740} /* (18, 24, 8) {real, imag} */,
  {32'hbecf8684, 32'hbea7a1e0} /* (18, 24, 7) {real, imag} */,
  {32'hbf22b6ea, 32'hbde6d080} /* (18, 24, 6) {real, imag} */,
  {32'hbee28390, 32'hbedcc390} /* (18, 24, 5) {real, imag} */,
  {32'hbcb52100, 32'hbed9d360} /* (18, 24, 4) {real, imag} */,
  {32'h3d505440, 32'hbe6f5340} /* (18, 24, 3) {real, imag} */,
  {32'hbfa5ab06, 32'h3e180c40} /* (18, 24, 2) {real, imag} */,
  {32'hbfafe866, 32'h3f675d80} /* (18, 24, 1) {real, imag} */,
  {32'hbf0ac25e, 32'h3f0f440c} /* (18, 24, 0) {real, imag} */,
  {32'hbe89ee12, 32'hbf5b3488} /* (18, 23, 31) {real, imag} */,
  {32'hbefe02ec, 32'hbee15020} /* (18, 23, 30) {real, imag} */,
  {32'hbf2d3f77, 32'h3deb3480} /* (18, 23, 29) {real, imag} */,
  {32'hbf1b9334, 32'h3d5b1700} /* (18, 23, 28) {real, imag} */,
  {32'hbf0dd5bc, 32'h3db8d500} /* (18, 23, 27) {real, imag} */,
  {32'hbf899e2d, 32'hbe9502d0} /* (18, 23, 26) {real, imag} */,
  {32'hbf5724ce, 32'h3e988fe0} /* (18, 23, 25) {real, imag} */,
  {32'hbf32706f, 32'hbccc0d00} /* (18, 23, 24) {real, imag} */,
  {32'hbc06f980, 32'hbf3d9b10} /* (18, 23, 23) {real, imag} */,
  {32'hbf2d2959, 32'hbeb0a6e0} /* (18, 23, 22) {real, imag} */,
  {32'hbf413d2a, 32'hbd7cdfc0} /* (18, 23, 21) {real, imag} */,
  {32'h3ecd52f0, 32'hbdb28a40} /* (18, 23, 20) {real, imag} */,
  {32'h3f6fe27a, 32'h3def0400} /* (18, 23, 19) {real, imag} */,
  {32'h3f566c96, 32'h3f44c7e0} /* (18, 23, 18) {real, imag} */,
  {32'h3fcea78f, 32'h3d3a4c00} /* (18, 23, 17) {real, imag} */,
  {32'h3fca72de, 32'h3e1fc860} /* (18, 23, 16) {real, imag} */,
  {32'h3ec8ecb0, 32'h3efb90e0} /* (18, 23, 15) {real, imag} */,
  {32'h3c3b2640, 32'h3e95ccc0} /* (18, 23, 14) {real, imag} */,
  {32'h3e321178, 32'h3ee04cf0} /* (18, 23, 13) {real, imag} */,
  {32'h3f9e4901, 32'h3f6cb138} /* (18, 23, 12) {real, imag} */,
  {32'hbdc49480, 32'h3e34e980} /* (18, 23, 11) {real, imag} */,
  {32'hbf93e224, 32'hbef25970} /* (18, 23, 10) {real, imag} */,
  {32'hbf695948, 32'h3dcbf840} /* (18, 23, 9) {real, imag} */,
  {32'h3f019508, 32'hbeb11440} /* (18, 23, 8) {real, imag} */,
  {32'hbe40a0a8, 32'hbf08d050} /* (18, 23, 7) {real, imag} */,
  {32'hbdc19270, 32'hbf302e10} /* (18, 23, 6) {real, imag} */,
  {32'h3c407ac0, 32'hbf8e70b4} /* (18, 23, 5) {real, imag} */,
  {32'hbf1246a2, 32'hbf695330} /* (18, 23, 4) {real, imag} */,
  {32'hbeeec85c, 32'hbf017be0} /* (18, 23, 3) {real, imag} */,
  {32'hbf37841c, 32'h3de67e00} /* (18, 23, 2) {real, imag} */,
  {32'hbef462a4, 32'h3f8c55b4} /* (18, 23, 1) {real, imag} */,
  {32'hbc8d0fb0, 32'h3e7b4aa0} /* (18, 23, 0) {real, imag} */,
  {32'hbf63616f, 32'hbe928ef0} /* (18, 22, 31) {real, imag} */,
  {32'hbf2d9843, 32'h3ed95100} /* (18, 22, 30) {real, imag} */,
  {32'hbe0691d8, 32'h3de7a300} /* (18, 22, 29) {real, imag} */,
  {32'h3e59e790, 32'hbee3e8c0} /* (18, 22, 28) {real, imag} */,
  {32'h3efcde00, 32'hbeb493f0} /* (18, 22, 27) {real, imag} */,
  {32'hbdc95ee0, 32'hbf16d1f8} /* (18, 22, 26) {real, imag} */,
  {32'hbed6439c, 32'h3eaadd50} /* (18, 22, 25) {real, imag} */,
  {32'hbf92f798, 32'h3e166700} /* (18, 22, 24) {real, imag} */,
  {32'hbef8428a, 32'h3ed3d2b0} /* (18, 22, 23) {real, imag} */,
  {32'hbeca71c8, 32'h3ed2cec0} /* (18, 22, 22) {real, imag} */,
  {32'hbf796bb8, 32'hbd85f0a0} /* (18, 22, 21) {real, imag} */,
  {32'h3e82ef06, 32'h3d51fb00} /* (18, 22, 20) {real, imag} */,
  {32'h3fa5d495, 32'hbe95f3f0} /* (18, 22, 19) {real, imag} */,
  {32'h3f850a2a, 32'hbce1ee00} /* (18, 22, 18) {real, imag} */,
  {32'h3f889b48, 32'hbe94e1e0} /* (18, 22, 17) {real, imag} */,
  {32'h3f9d1f90, 32'h3e7a1e20} /* (18, 22, 16) {real, imag} */,
  {32'h3f282fcc, 32'hbb752000} /* (18, 22, 15) {real, imag} */,
  {32'h3f34e526, 32'hbf2787b0} /* (18, 22, 14) {real, imag} */,
  {32'h3f2e11f0, 32'h3d69e200} /* (18, 22, 13) {real, imag} */,
  {32'h3e71b028, 32'hbec949c0} /* (18, 22, 12) {real, imag} */,
  {32'hbde38cc0, 32'hbe2867c0} /* (18, 22, 11) {real, imag} */,
  {32'hbf31e752, 32'h3e945aa0} /* (18, 22, 10) {real, imag} */,
  {32'hbf2c439c, 32'h3efca820} /* (18, 22, 9) {real, imag} */,
  {32'hbecd228c, 32'h3eba3980} /* (18, 22, 8) {real, imag} */,
  {32'hbf28a748, 32'h3dd8d400} /* (18, 22, 7) {real, imag} */,
  {32'hbf193747, 32'hbe0ce880} /* (18, 22, 6) {real, imag} */,
  {32'hbe9b991e, 32'hbe42e840} /* (18, 22, 5) {real, imag} */,
  {32'hbf173d8c, 32'h3c5c0a00} /* (18, 22, 4) {real, imag} */,
  {32'hbf999c5d, 32'hbeaef450} /* (18, 22, 3) {real, imag} */,
  {32'hbf338db8, 32'hbf4d5780} /* (18, 22, 2) {real, imag} */,
  {32'hbea1d4a8, 32'hbe1463c0} /* (18, 22, 1) {real, imag} */,
  {32'hbedb3249, 32'hbe560de0} /* (18, 22, 0) {real, imag} */,
  {32'hbf1b3004, 32'h3e84231c} /* (18, 21, 31) {real, imag} */,
  {32'hbf6b91ae, 32'h3f30128c} /* (18, 21, 30) {real, imag} */,
  {32'hbf3a8099, 32'h3ef06408} /* (18, 21, 29) {real, imag} */,
  {32'hbf0cc7fc, 32'hbef9bd80} /* (18, 21, 28) {real, imag} */,
  {32'h3dfa1e40, 32'hbf56eb14} /* (18, 21, 27) {real, imag} */,
  {32'h3f15e298, 32'hbee80ed8} /* (18, 21, 26) {real, imag} */,
  {32'h3e74aa88, 32'hbe053632} /* (18, 21, 25) {real, imag} */,
  {32'hbe960594, 32'hbe253968} /* (18, 21, 24) {real, imag} */,
  {32'h3effc094, 32'h3ee6b740} /* (18, 21, 23) {real, imag} */,
  {32'hbf040c6a, 32'h3ee18ff0} /* (18, 21, 22) {real, imag} */,
  {32'hbf96991e, 32'hbe8e1550} /* (18, 21, 21) {real, imag} */,
  {32'hbf32daaa, 32'hbf207f9e} /* (18, 21, 20) {real, imag} */,
  {32'h3ddf4f00, 32'hbf028f00} /* (18, 21, 19) {real, imag} */,
  {32'h3f522507, 32'h3ce39180} /* (18, 21, 18) {real, imag} */,
  {32'h3f8ff9b3, 32'hbf2f89ca} /* (18, 21, 17) {real, imag} */,
  {32'h3ea1ecab, 32'hbca65000} /* (18, 21, 16) {real, imag} */,
  {32'hbe5394d4, 32'h3e944e40} /* (18, 21, 15) {real, imag} */,
  {32'h3f58a677, 32'hbef439a0} /* (18, 21, 14) {real, imag} */,
  {32'h39c7f800, 32'hbef842b0} /* (18, 21, 13) {real, imag} */,
  {32'hbf60ace9, 32'hbfb324e4} /* (18, 21, 12) {real, imag} */,
  {32'h3e015c78, 32'hbf1ac0f0} /* (18, 21, 11) {real, imag} */,
  {32'hbd2beab8, 32'h3ec177fc} /* (18, 21, 10) {real, imag} */,
  {32'hbea0d75c, 32'h3d51abc0} /* (18, 21, 9) {real, imag} */,
  {32'hbea7af7c, 32'hbe2e6b10} /* (18, 21, 8) {real, imag} */,
  {32'hbf41de3b, 32'h3f291b14} /* (18, 21, 7) {real, imag} */,
  {32'hbf64edca, 32'h3eec6264} /* (18, 21, 6) {real, imag} */,
  {32'hbef995c7, 32'h3e2871b0} /* (18, 21, 5) {real, imag} */,
  {32'h3ea99e94, 32'h3f57fcf0} /* (18, 21, 4) {real, imag} */,
  {32'hbd0a22b0, 32'h3ebc7758} /* (18, 21, 3) {real, imag} */,
  {32'hbdbbe100, 32'h3e5e4480} /* (18, 21, 2) {real, imag} */,
  {32'hbf150309, 32'h3eb65720} /* (18, 21, 1) {real, imag} */,
  {32'hbef81c9c, 32'hbd3a6500} /* (18, 21, 0) {real, imag} */,
  {32'hbe6e1d76, 32'hbe7841b0} /* (18, 20, 31) {real, imag} */,
  {32'h3d536640, 32'hbee758b0} /* (18, 20, 30) {real, imag} */,
  {32'hbebd7814, 32'h3ea0dca0} /* (18, 20, 29) {real, imag} */,
  {32'hbed5157c, 32'hbc9c0c00} /* (18, 20, 28) {real, imag} */,
  {32'h3ef900c4, 32'hbf06aa60} /* (18, 20, 27) {real, imag} */,
  {32'h3eedbbec, 32'hbf63cce8} /* (18, 20, 26) {real, imag} */,
  {32'h3f4062ce, 32'hbe4152c0} /* (18, 20, 25) {real, imag} */,
  {32'h3f27287c, 32'hbe245780} /* (18, 20, 24) {real, imag} */,
  {32'h3f702378, 32'hbf3d1160} /* (18, 20, 23) {real, imag} */,
  {32'hbf02e9e6, 32'hbf6ace50} /* (18, 20, 22) {real, imag} */,
  {32'hbf66f5cc, 32'hbec8d41c} /* (18, 20, 21) {real, imag} */,
  {32'hbf839c96, 32'hbedd2a00} /* (18, 20, 20) {real, imag} */,
  {32'hbf9f457a, 32'hbecf7030} /* (18, 20, 19) {real, imag} */,
  {32'h3ee79b46, 32'hbf288f28} /* (18, 20, 18) {real, imag} */,
  {32'h3e906e3a, 32'hbf877dc8} /* (18, 20, 17) {real, imag} */,
  {32'hbf46423e, 32'hbf02f2b0} /* (18, 20, 16) {real, imag} */,
  {32'hbf2149be, 32'h3e3abfa0} /* (18, 20, 15) {real, imag} */,
  {32'hbc834640, 32'h3db34980} /* (18, 20, 14) {real, imag} */,
  {32'hbecb7fb0, 32'hbee016d0} /* (18, 20, 13) {real, imag} */,
  {32'hbed50840, 32'hbf883570} /* (18, 20, 12) {real, imag} */,
  {32'hbcad80c0, 32'h3eabe4c8} /* (18, 20, 11) {real, imag} */,
  {32'h3e137bb0, 32'h3fa7cb8b} /* (18, 20, 10) {real, imag} */,
  {32'h3e186760, 32'h3c46b200} /* (18, 20, 9) {real, imag} */,
  {32'h3e93884c, 32'hbf396a6c} /* (18, 20, 8) {real, imag} */,
  {32'h3e7f8a48, 32'h3d9ae380} /* (18, 20, 7) {real, imag} */,
  {32'h3f0fc7a1, 32'h3e6d8880} /* (18, 20, 6) {real, imag} */,
  {32'h3f8e5980, 32'h3e298520} /* (18, 20, 5) {real, imag} */,
  {32'h3fa3b9ec, 32'h3eeb1990} /* (18, 20, 4) {real, imag} */,
  {32'h3f83a2d8, 32'h3f9407a0} /* (18, 20, 3) {real, imag} */,
  {32'h3f31cab0, 32'h3f9fce0c} /* (18, 20, 2) {real, imag} */,
  {32'h3eb08170, 32'h3f29fdd8} /* (18, 20, 1) {real, imag} */,
  {32'h3e8a3bd8, 32'hbe5669a0} /* (18, 20, 0) {real, imag} */,
  {32'h3f0122eb, 32'h3a136000} /* (18, 19, 31) {real, imag} */,
  {32'h3f7f7800, 32'hbeb1d620} /* (18, 19, 30) {real, imag} */,
  {32'h3f739ce6, 32'h3f5eedf0} /* (18, 19, 29) {real, imag} */,
  {32'h3f9a5edc, 32'h3eb65420} /* (18, 19, 28) {real, imag} */,
  {32'h3f52dcbb, 32'hbe683a80} /* (18, 19, 27) {real, imag} */,
  {32'h3ee30d76, 32'hbebd8280} /* (18, 19, 26) {real, imag} */,
  {32'h3f51f38a, 32'h3ed4f960} /* (18, 19, 25) {real, imag} */,
  {32'h3f19c3c0, 32'h3ec32500} /* (18, 19, 24) {real, imag} */,
  {32'h3f34edf4, 32'hbe3926c0} /* (18, 19, 23) {real, imag} */,
  {32'h3e8f7a3c, 32'hbf20c390} /* (18, 19, 22) {real, imag} */,
  {32'hbef2a33a, 32'hbf774cb0} /* (18, 19, 21) {real, imag} */,
  {32'hbf72e26a, 32'hbf7d9cc8} /* (18, 19, 20) {real, imag} */,
  {32'hbfadfbb8, 32'hbf093d60} /* (18, 19, 19) {real, imag} */,
  {32'hbe5ed82e, 32'hbf1faf78} /* (18, 19, 18) {real, imag} */,
  {32'hbdddfde0, 32'hbf43d310} /* (18, 19, 17) {real, imag} */,
  {32'hbf0b1898, 32'hbf18e4c8} /* (18, 19, 16) {real, imag} */,
  {32'hbe242a70, 32'hbf0b4640} /* (18, 19, 15) {real, imag} */,
  {32'hbdf42800, 32'hbe45efc0} /* (18, 19, 14) {real, imag} */,
  {32'hbef5336a, 32'hbeca3aa0} /* (18, 19, 13) {real, imag} */,
  {32'h3d31cdf0, 32'hbf76c5a0} /* (18, 19, 12) {real, imag} */,
  {32'h3e25af74, 32'h3ee31190} /* (18, 19, 11) {real, imag} */,
  {32'h3e4ada1c, 32'h3f2dcdec} /* (18, 19, 10) {real, imag} */,
  {32'h3f1c52bc, 32'hbee33c20} /* (18, 19, 9) {real, imag} */,
  {32'h3e25cf60, 32'hbe70afa0} /* (18, 19, 8) {real, imag} */,
  {32'h3e9894b0, 32'hbeb86500} /* (18, 19, 7) {real, imag} */,
  {32'h3e40349c, 32'hbedf8600} /* (18, 19, 6) {real, imag} */,
  {32'h3f5125f8, 32'hbe823540} /* (18, 19, 5) {real, imag} */,
  {32'h3f7fb76a, 32'hbea025b0} /* (18, 19, 4) {real, imag} */,
  {32'h3f1217c4, 32'h3f36b238} /* (18, 19, 3) {real, imag} */,
  {32'h3fa21718, 32'h3f9a8348} /* (18, 19, 2) {real, imag} */,
  {32'h3fa0ce7e, 32'h3dff01c0} /* (18, 19, 1) {real, imag} */,
  {32'h3f0cfb8b, 32'hbf2c627c} /* (18, 19, 0) {real, imag} */,
  {32'h3ebdbd06, 32'hbd616080} /* (18, 18, 31) {real, imag} */,
  {32'h3f48a584, 32'hbf0d2f20} /* (18, 18, 30) {real, imag} */,
  {32'h3ebe9154, 32'h3eda1f50} /* (18, 18, 29) {real, imag} */,
  {32'h3f4cb151, 32'hbddbbe00} /* (18, 18, 28) {real, imag} */,
  {32'h3f563a78, 32'hbf638708} /* (18, 18, 27) {real, imag} */,
  {32'h3f30563a, 32'h3e2f6700} /* (18, 18, 26) {real, imag} */,
  {32'h3f1b7be0, 32'h3f91ad38} /* (18, 18, 25) {real, imag} */,
  {32'h3fa54f60, 32'h3fa49974} /* (18, 18, 24) {real, imag} */,
  {32'h3ff01d04, 32'h3f3fc310} /* (18, 18, 23) {real, imag} */,
  {32'h3f4e218e, 32'hbe7ae3a0} /* (18, 18, 22) {real, imag} */,
  {32'hbeae4d41, 32'hbfd9c0ec} /* (18, 18, 21) {real, imag} */,
  {32'hbf4cf5d6, 32'hbf7e3b08} /* (18, 18, 20) {real, imag} */,
  {32'hbfbb08b6, 32'hbf46f3d0} /* (18, 18, 19) {real, imag} */,
  {32'hbffad278, 32'hbf6e8588} /* (18, 18, 18) {real, imag} */,
  {32'hbf7eb224, 32'hbf780f20} /* (18, 18, 17) {real, imag} */,
  {32'hbeeb51e8, 32'hbf067cf8} /* (18, 18, 16) {real, imag} */,
  {32'hbef75e30, 32'hbe9a2520} /* (18, 18, 15) {real, imag} */,
  {32'hbe7a0848, 32'h3dcea540} /* (18, 18, 14) {real, imag} */,
  {32'hbf145aee, 32'hbea109c0} /* (18, 18, 13) {real, imag} */,
  {32'hbf2b1dda, 32'hbe1533c0} /* (18, 18, 12) {real, imag} */,
  {32'h3e98269c, 32'h3f50a758} /* (18, 18, 11) {real, imag} */,
  {32'h3c5fc2c0, 32'h3f04424c} /* (18, 18, 10) {real, imag} */,
  {32'h3daa2b30, 32'hbefd5960} /* (18, 18, 9) {real, imag} */,
  {32'h3f71fc8e, 32'hbe66b200} /* (18, 18, 8) {real, imag} */,
  {32'h3f92cf26, 32'hbb8e0000} /* (18, 18, 7) {real, imag} */,
  {32'h3f26a651, 32'h3e816e80} /* (18, 18, 6) {real, imag} */,
  {32'h3e54e0ec, 32'h3d8ef080} /* (18, 18, 5) {real, imag} */,
  {32'h3e999350, 32'h3d4e1580} /* (18, 18, 4) {real, imag} */,
  {32'h3ebaeef0, 32'h3edb8e20} /* (18, 18, 3) {real, imag} */,
  {32'h3f8f9af8, 32'h3e714d40} /* (18, 18, 2) {real, imag} */,
  {32'h3f9bbe10, 32'hbeb25f40} /* (18, 18, 1) {real, imag} */,
  {32'h3eaa526c, 32'hbf2942b8} /* (18, 18, 0) {real, imag} */,
  {32'h3de8b450, 32'hbee73d40} /* (18, 17, 31) {real, imag} */,
  {32'h3e423210, 32'hbe98fd30} /* (18, 17, 30) {real, imag} */,
  {32'h3ebecd58, 32'h3e299400} /* (18, 17, 29) {real, imag} */,
  {32'h3f482fba, 32'hbea663b0} /* (18, 17, 28) {real, imag} */,
  {32'h3f5a28ac, 32'hbf242178} /* (18, 17, 27) {real, imag} */,
  {32'h3f468de6, 32'h3d377900} /* (18, 17, 26) {real, imag} */,
  {32'h3f394772, 32'h3eaa28f0} /* (18, 17, 25) {real, imag} */,
  {32'h3f4a0228, 32'h3f25a8f0} /* (18, 17, 24) {real, imag} */,
  {32'h3f23f34c, 32'h3f0a2cb0} /* (18, 17, 23) {real, imag} */,
  {32'h3f8c1620, 32'h3f01a140} /* (18, 17, 22) {real, imag} */,
  {32'h3f2fdd29, 32'hbe066200} /* (18, 17, 21) {real, imag} */,
  {32'hbe3e9c50, 32'h3a032000} /* (18, 17, 20) {real, imag} */,
  {32'h3e6dd3da, 32'hbde02d00} /* (18, 17, 19) {real, imag} */,
  {32'hbfa1955d, 32'hbf321280} /* (18, 17, 18) {real, imag} */,
  {32'hbffbc3ef, 32'hbfe34d54} /* (18, 17, 17) {real, imag} */,
  {32'hbf97a146, 32'hbf1d21a0} /* (18, 17, 16) {real, imag} */,
  {32'hbfa40a22, 32'hbc515a00} /* (18, 17, 15) {real, imag} */,
  {32'hbf9de5f2, 32'h3f049aa8} /* (18, 17, 14) {real, imag} */,
  {32'hbeba39f0, 32'h3e24d600} /* (18, 17, 13) {real, imag} */,
  {32'hbf033892, 32'h3f2e7950} /* (18, 17, 12) {real, imag} */,
  {32'h3dd02880, 32'h3f22a950} /* (18, 17, 11) {real, imag} */,
  {32'hbd42eb40, 32'h3e677e80} /* (18, 17, 10) {real, imag} */,
  {32'h3f31cae0, 32'h3cff8500} /* (18, 17, 9) {real, imag} */,
  {32'h3fb3d558, 32'h3e9211b0} /* (18, 17, 8) {real, imag} */,
  {32'h3faddb8b, 32'h3eb51d00} /* (18, 17, 7) {real, imag} */,
  {32'h3f689a92, 32'h3f0b3dd8} /* (18, 17, 6) {real, imag} */,
  {32'hbea44400, 32'h3d8a3780} /* (18, 17, 5) {real, imag} */,
  {32'hbed67bfc, 32'h3e1dd200} /* (18, 17, 4) {real, imag} */,
  {32'h3eced3f8, 32'h3d70e800} /* (18, 17, 3) {real, imag} */,
  {32'h3f14b166, 32'hbd773400} /* (18, 17, 2) {real, imag} */,
  {32'h3f7ad82c, 32'h3d296500} /* (18, 17, 1) {real, imag} */,
  {32'h3f13aa84, 32'hbf009eac} /* (18, 17, 0) {real, imag} */,
  {32'h3ee3880c, 32'hbed57f48} /* (18, 16, 31) {real, imag} */,
  {32'h3e6f4290, 32'hbebf4030} /* (18, 16, 30) {real, imag} */,
  {32'h3f11e964, 32'hbe3518e0} /* (18, 16, 29) {real, imag} */,
  {32'h3f608954, 32'h3e9304c0} /* (18, 16, 28) {real, imag} */,
  {32'h3fb68ebc, 32'h3e905210} /* (18, 16, 27) {real, imag} */,
  {32'h3f93b5c1, 32'hbdd99640} /* (18, 16, 26) {real, imag} */,
  {32'h3f05e5d7, 32'hbded2d80} /* (18, 16, 25) {real, imag} */,
  {32'hbd994bf0, 32'hbeade9a0} /* (18, 16, 24) {real, imag} */,
  {32'hbe65b4a4, 32'hbedee680} /* (18, 16, 23) {real, imag} */,
  {32'h3f03be0c, 32'h3de82e80} /* (18, 16, 22) {real, imag} */,
  {32'h3ed501e8, 32'h3f2c1a84} /* (18, 16, 21) {real, imag} */,
  {32'hbe2ff178, 32'h3ea6fdc0} /* (18, 16, 20) {real, imag} */,
  {32'h3f64d22d, 32'h3f233410} /* (18, 16, 19) {real, imag} */,
  {32'h3cf10cc0, 32'h3efe7020} /* (18, 16, 18) {real, imag} */,
  {32'hbf4101d0, 32'hbea03240} /* (18, 16, 17) {real, imag} */,
  {32'hbf84b2cb, 32'hbdf9de80} /* (18, 16, 16) {real, imag} */,
  {32'hbfb93280, 32'hbf991110} /* (18, 16, 15) {real, imag} */,
  {32'hbfe414ac, 32'hbeb5dc00} /* (18, 16, 14) {real, imag} */,
  {32'hbf71a592, 32'hbe809a50} /* (18, 16, 13) {real, imag} */,
  {32'hbf87f8b7, 32'h3f032838} /* (18, 16, 12) {real, imag} */,
  {32'h3e145a04, 32'h3f24b970} /* (18, 16, 11) {real, imag} */,
  {32'h3d0643a0, 32'h3f4ef214} /* (18, 16, 10) {real, imag} */,
  {32'h3f6c8b7c, 32'h3fb48670} /* (18, 16, 9) {real, imag} */,
  {32'h4001da3c, 32'h3f3e50a8} /* (18, 16, 8) {real, imag} */,
  {32'h3fb3a2e2, 32'h3f28efb8} /* (18, 16, 7) {real, imag} */,
  {32'h3f526c78, 32'h3e8b0770} /* (18, 16, 6) {real, imag} */,
  {32'h3e1d66ec, 32'h3db46a00} /* (18, 16, 5) {real, imag} */,
  {32'h3ede16ec, 32'hbd55c600} /* (18, 16, 4) {real, imag} */,
  {32'h3f830925, 32'hbe4beec0} /* (18, 16, 3) {real, imag} */,
  {32'h3fd237df, 32'h3dff5400} /* (18, 16, 2) {real, imag} */,
  {32'h3fbee468, 32'h3f82ed00} /* (18, 16, 1) {real, imag} */,
  {32'h3f1e0d1e, 32'hbd1ad800} /* (18, 16, 0) {real, imag} */,
  {32'h3f8b96c4, 32'hbe591b80} /* (18, 15, 31) {real, imag} */,
  {32'h3f0ca140, 32'hbf0de050} /* (18, 15, 30) {real, imag} */,
  {32'h3f362d90, 32'hbf3e4950} /* (18, 15, 29) {real, imag} */,
  {32'h3ec90014, 32'hbedd6a20} /* (18, 15, 28) {real, imag} */,
  {32'h3e40a170, 32'h3eeef5d0} /* (18, 15, 27) {real, imag} */,
  {32'h3ecf2f3c, 32'h3f273db0} /* (18, 15, 26) {real, imag} */,
  {32'h3e46b250, 32'h3edf3c00} /* (18, 15, 25) {real, imag} */,
  {32'hbec698e0, 32'hbe574ee0} /* (18, 15, 24) {real, imag} */,
  {32'hbf350aba, 32'hbecce330} /* (18, 15, 23) {real, imag} */,
  {32'hbf062c52, 32'hbf134450} /* (18, 15, 22) {real, imag} */,
  {32'hbe8f9020, 32'hbe8202dc} /* (18, 15, 21) {real, imag} */,
  {32'hbe952a14, 32'hbeb4f0a0} /* (18, 15, 20) {real, imag} */,
  {32'h3f1c2136, 32'h3e6038e0} /* (18, 15, 19) {real, imag} */,
  {32'hbf182292, 32'h3dce5340} /* (18, 15, 18) {real, imag} */,
  {32'hbf50fd82, 32'h3eeb2700} /* (18, 15, 17) {real, imag} */,
  {32'hbf56ba78, 32'h3ee4d220} /* (18, 15, 16) {real, imag} */,
  {32'hbfa74087, 32'hbf3ac578} /* (18, 15, 15) {real, imag} */,
  {32'hbfed2385, 32'hbedb0ea0} /* (18, 15, 14) {real, imag} */,
  {32'hbfbaaa18, 32'hbe24b1c0} /* (18, 15, 13) {real, imag} */,
  {32'hbf4ebcdc, 32'h3e75eac0} /* (18, 15, 12) {real, imag} */,
  {32'h3e436ecc, 32'h3ee61b60} /* (18, 15, 11) {real, imag} */,
  {32'h3d6a1500, 32'h3f8fae28} /* (18, 15, 10) {real, imag} */,
  {32'h3efd1110, 32'h3fe17664} /* (18, 15, 9) {real, imag} */,
  {32'h3f8ee368, 32'h3e8f9950} /* (18, 15, 8) {real, imag} */,
  {32'h3fcca86e, 32'h3f022ee0} /* (18, 15, 7) {real, imag} */,
  {32'h3ee0bd3c, 32'h3ed56270} /* (18, 15, 6) {real, imag} */,
  {32'h3d5972f0, 32'h3dd41d80} /* (18, 15, 5) {real, imag} */,
  {32'h3f8167ce, 32'hbe367580} /* (18, 15, 4) {real, imag} */,
  {32'h3f5be158, 32'hbf131fd8} /* (18, 15, 3) {real, imag} */,
  {32'h3f8d5194, 32'h3c8fa400} /* (18, 15, 2) {real, imag} */,
  {32'h3f8c452e, 32'h3efe9090} /* (18, 15, 1) {real, imag} */,
  {32'h3f331603, 32'hbe30b1c0} /* (18, 15, 0) {real, imag} */,
  {32'h3e8417a8, 32'hbf111f80} /* (18, 14, 31) {real, imag} */,
  {32'hbe187e10, 32'h3ee1d580} /* (18, 14, 30) {real, imag} */,
  {32'h3f61aeee, 32'h3f0e0ab0} /* (18, 14, 29) {real, imag} */,
  {32'h3f08e206, 32'h3eb29160} /* (18, 14, 28) {real, imag} */,
  {32'hbe17c5f0, 32'h3f01e368} /* (18, 14, 27) {real, imag} */,
  {32'h3eaf1548, 32'h3e522900} /* (18, 14, 26) {real, imag} */,
  {32'h3f377fb8, 32'h3da6cc40} /* (18, 14, 25) {real, imag} */,
  {32'h3e9bae4e, 32'h3df6f6c0} /* (18, 14, 24) {real, imag} */,
  {32'hbe30e4ce, 32'h3e2aff60} /* (18, 14, 23) {real, imag} */,
  {32'h3e006b90, 32'h3c452000} /* (18, 14, 22) {real, imag} */,
  {32'h3b87ab00, 32'hbe287660} /* (18, 14, 21) {real, imag} */,
  {32'hbf0e9e1f, 32'hbf16a190} /* (18, 14, 20) {real, imag} */,
  {32'hbe1de160, 32'hbf805f7c} /* (18, 14, 19) {real, imag} */,
  {32'hbef89fa8, 32'hbee9c0c0} /* (18, 14, 18) {real, imag} */,
  {32'hbf6a412a, 32'hbd882d80} /* (18, 14, 17) {real, imag} */,
  {32'hbecfd63d, 32'h3d43f700} /* (18, 14, 16) {real, imag} */,
  {32'hbd8391e8, 32'hbc76d200} /* (18, 14, 15) {real, imag} */,
  {32'hbf215798, 32'h3d0bfa00} /* (18, 14, 14) {real, imag} */,
  {32'hbd9a0e20, 32'h3d945980} /* (18, 14, 13) {real, imag} */,
  {32'h3e8abf54, 32'hbe9a6bb0} /* (18, 14, 12) {real, imag} */,
  {32'hbef018b0, 32'hbe5b6540} /* (18, 14, 11) {real, imag} */,
  {32'h3d973970, 32'h3f083c46} /* (18, 14, 10) {real, imag} */,
  {32'h3ee7e110, 32'h3f087f48} /* (18, 14, 9) {real, imag} */,
  {32'h3f21ea98, 32'hbe180580} /* (18, 14, 8) {real, imag} */,
  {32'h3fa6a27e, 32'hbe7c1700} /* (18, 14, 7) {real, imag} */,
  {32'h3f95bed2, 32'hbe253b20} /* (18, 14, 6) {real, imag} */,
  {32'h3f410e10, 32'hbe24c360} /* (18, 14, 5) {real, imag} */,
  {32'h3e94f6a4, 32'h3e647180} /* (18, 14, 4) {real, imag} */,
  {32'h3e6d9fd0, 32'h3e924ea0} /* (18, 14, 3) {real, imag} */,
  {32'h3f367bb4, 32'h3de0a400} /* (18, 14, 2) {real, imag} */,
  {32'h3f7bb75c, 32'hbf73d6d0} /* (18, 14, 1) {real, imag} */,
  {32'h3f6bdafc, 32'hbf7369d0} /* (18, 14, 0) {real, imag} */,
  {32'hbdec1b14, 32'hbe109c80} /* (18, 13, 31) {real, imag} */,
  {32'h3dfda2b0, 32'h3ea6b110} /* (18, 13, 30) {real, imag} */,
  {32'h3f3cf31e, 32'h3f3af6f0} /* (18, 13, 29) {real, imag} */,
  {32'h3ec447e4, 32'h3f66ad60} /* (18, 13, 28) {real, imag} */,
  {32'h3f29275f, 32'h3e8475c0} /* (18, 13, 27) {real, imag} */,
  {32'h3f60ea5e, 32'h3e196900} /* (18, 13, 26) {real, imag} */,
  {32'h3f873e10, 32'h3f0363b0} /* (18, 13, 25) {real, imag} */,
  {32'h3fb234fa, 32'h3d26b780} /* (18, 13, 24) {real, imag} */,
  {32'h3f72c19b, 32'h3e26f560} /* (18, 13, 23) {real, imag} */,
  {32'h3fcb2879, 32'h3f0ffac0} /* (18, 13, 22) {real, imag} */,
  {32'h3ec1639c, 32'h3f4e0780} /* (18, 13, 21) {real, imag} */,
  {32'hbf72f776, 32'h3e34b220} /* (18, 13, 20) {real, imag} */,
  {32'hbdc57240, 32'hbf80b5b8} /* (18, 13, 19) {real, imag} */,
  {32'h3dcb6170, 32'hbf3ba920} /* (18, 13, 18) {real, imag} */,
  {32'hbe18ade0, 32'hbf473740} /* (18, 13, 17) {real, imag} */,
  {32'hbea6de88, 32'hbf3b3b18} /* (18, 13, 16) {real, imag} */,
  {32'hbe6152b0, 32'hbe8b5850} /* (18, 13, 15) {real, imag} */,
  {32'hbf0e7b9c, 32'hbe2ad5c0} /* (18, 13, 14) {real, imag} */,
  {32'hbf7438f6, 32'hbf376bc8} /* (18, 13, 13) {real, imag} */,
  {32'hbf95dbd9, 32'hbf410c10} /* (18, 13, 12) {real, imag} */,
  {32'hbf5299e4, 32'hbeebde80} /* (18, 13, 11) {real, imag} */,
  {32'hbd9b5678, 32'h3e660d28} /* (18, 13, 10) {real, imag} */,
  {32'hbe97eb18, 32'h3dfccd80} /* (18, 13, 9) {real, imag} */,
  {32'h3e42afa8, 32'h3ea5cd60} /* (18, 13, 8) {real, imag} */,
  {32'h3fc48c07, 32'h3e8ff080} /* (18, 13, 7) {real, imag} */,
  {32'h3ff373e7, 32'hbe2ccbc0} /* (18, 13, 6) {real, imag} */,
  {32'h3f517039, 32'hbf499b78} /* (18, 13, 5) {real, imag} */,
  {32'h3e8d30ef, 32'hbf3bcc30} /* (18, 13, 4) {real, imag} */,
  {32'h3e4903d0, 32'hbf1f1058} /* (18, 13, 3) {real, imag} */,
  {32'h3f38f3e8, 32'hbf452190} /* (18, 13, 2) {real, imag} */,
  {32'h3f849c9d, 32'hbfb6e124} /* (18, 13, 1) {real, imag} */,
  {32'h3eb74e72, 32'hbf8424c8} /* (18, 13, 0) {real, imag} */,
  {32'h3eedc40f, 32'hbe54c550} /* (18, 12, 31) {real, imag} */,
  {32'h3f18de82, 32'hbe9df420} /* (18, 12, 30) {real, imag} */,
  {32'h3efcb8f8, 32'h3e8fb240} /* (18, 12, 29) {real, imag} */,
  {32'h3f67201c, 32'h3eda8c70} /* (18, 12, 28) {real, imag} */,
  {32'h3f94f100, 32'h3d3e9780} /* (18, 12, 27) {real, imag} */,
  {32'h3f5ee432, 32'hbe720e00} /* (18, 12, 26) {real, imag} */,
  {32'h3eff1e18, 32'h3e863dd0} /* (18, 12, 25) {real, imag} */,
  {32'h3e4795c0, 32'hbe9d2dd0} /* (18, 12, 24) {real, imag} */,
  {32'h3d3194a0, 32'hbe1dd920} /* (18, 12, 23) {real, imag} */,
  {32'h3e848440, 32'h3f2a1980} /* (18, 12, 22) {real, imag} */,
  {32'h3e8af8e4, 32'h3f3be740} /* (18, 12, 21) {real, imag} */,
  {32'hbf31025e, 32'h3e2a6900} /* (18, 12, 20) {real, imag} */,
  {32'hbed78120, 32'hbee85580} /* (18, 12, 19) {real, imag} */,
  {32'hbecc6164, 32'hbebbed00} /* (18, 12, 18) {real, imag} */,
  {32'hbf3419e0, 32'hbf95c864} /* (18, 12, 17) {real, imag} */,
  {32'hbf6b9e80, 32'hbf8430a0} /* (18, 12, 16) {real, imag} */,
  {32'hbea0e670, 32'hbda65300} /* (18, 12, 15) {real, imag} */,
  {32'hbf246dce, 32'hbee8d870} /* (18, 12, 14) {real, imag} */,
  {32'hbf88dfb2, 32'hbf1ad0b8} /* (18, 12, 13) {real, imag} */,
  {32'hbfdb64a2, 32'hbf283770} /* (18, 12, 12) {real, imag} */,
  {32'hbfdeb992, 32'hbed0a7a0} /* (18, 12, 11) {real, imag} */,
  {32'hbed7c3af, 32'hbe7a3800} /* (18, 12, 10) {real, imag} */,
  {32'h3ee315d4, 32'hbd83c240} /* (18, 12, 9) {real, imag} */,
  {32'h3fc14016, 32'h3e5a3940} /* (18, 12, 8) {real, imag} */,
  {32'h3fb5900a, 32'hbef7a300} /* (18, 12, 7) {real, imag} */,
  {32'h3f9b73f2, 32'hbf116440} /* (18, 12, 6) {real, imag} */,
  {32'h3fa082ef, 32'hbf6c8320} /* (18, 12, 5) {real, imag} */,
  {32'h3f707d23, 32'hbfc137f4} /* (18, 12, 4) {real, imag} */,
  {32'h3efaab0c, 32'hbfca34e0} /* (18, 12, 3) {real, imag} */,
  {32'h3fa141ce, 32'hbf144db0} /* (18, 12, 2) {real, imag} */,
  {32'h3f9b703e, 32'hbdcaf280} /* (18, 12, 1) {real, imag} */,
  {32'h3f0c345d, 32'hbe4a7ac0} /* (18, 12, 0) {real, imag} */,
  {32'h3ebc4c68, 32'h3e23e840} /* (18, 11, 31) {real, imag} */,
  {32'h3ed860bd, 32'h3f28fc40} /* (18, 11, 30) {real, imag} */,
  {32'h3f72e278, 32'h3f050010} /* (18, 11, 29) {real, imag} */,
  {32'h4011fa0f, 32'hbe091ac0} /* (18, 11, 28) {real, imag} */,
  {32'h3faa50aa, 32'hbc0c8a00} /* (18, 11, 27) {real, imag} */,
  {32'hbe3fc614, 32'hbe0d6ec0} /* (18, 11, 26) {real, imag} */,
  {32'hbefd8ea0, 32'h3f30d1f8} /* (18, 11, 25) {real, imag} */,
  {32'hbe99a3be, 32'h3ea61b80} /* (18, 11, 24) {real, imag} */,
  {32'hbf0c43f9, 32'hbebcbcf0} /* (18, 11, 23) {real, imag} */,
  {32'hbebb5f8a, 32'h3cd39800} /* (18, 11, 22) {real, imag} */,
  {32'hbe37ab18, 32'h3f196544} /* (18, 11, 21) {real, imag} */,
  {32'hbe7d0ad8, 32'h3f3f6b10} /* (18, 11, 20) {real, imag} */,
  {32'hbe57b1cb, 32'h3dccad80} /* (18, 11, 19) {real, imag} */,
  {32'hbf78dce1, 32'hbde0a6c0} /* (18, 11, 18) {real, imag} */,
  {32'hbf830942, 32'hbf7359c8} /* (18, 11, 17) {real, imag} */,
  {32'hbefc0b0c, 32'hbf0644b0} /* (18, 11, 16) {real, imag} */,
  {32'h3e9ba9f8, 32'h3e971dd0} /* (18, 11, 15) {real, imag} */,
  {32'hbec25ef8, 32'hbd33e780} /* (18, 11, 14) {real, imag} */,
  {32'hbf09b0da, 32'hbf3fa9f8} /* (18, 11, 13) {real, imag} */,
  {32'hbf02f96e, 32'hbe877fa0} /* (18, 11, 12) {real, imag} */,
  {32'hbfcbed02, 32'h3e9f0bc8} /* (18, 11, 11) {real, imag} */,
  {32'hbf1acac7, 32'hbea93b90} /* (18, 11, 10) {real, imag} */,
  {32'h3ee44a16, 32'hbec17e40} /* (18, 11, 9) {real, imag} */,
  {32'h3f597fa7, 32'h3ced0700} /* (18, 11, 8) {real, imag} */,
  {32'h3f4251a0, 32'hbe5280c0} /* (18, 11, 7) {real, imag} */,
  {32'h3fc29652, 32'hbee29a70} /* (18, 11, 6) {real, imag} */,
  {32'h3fcc617d, 32'hbef91548} /* (18, 11, 5) {real, imag} */,
  {32'h3f864a3a, 32'hbd0fa900} /* (18, 11, 4) {real, imag} */,
  {32'h3ecdcf32, 32'hbd905100} /* (18, 11, 3) {real, imag} */,
  {32'h3f9d03a8, 32'h3eb8e5b0} /* (18, 11, 2) {real, imag} */,
  {32'h3f36492e, 32'h3f08c9b0} /* (18, 11, 1) {real, imag} */,
  {32'h3f030e0d, 32'h3e1a3ea0} /* (18, 11, 0) {real, imag} */,
  {32'hbe331e8d, 32'hbe51cd70} /* (18, 10, 31) {real, imag} */,
  {32'hbe092c00, 32'h3e160a10} /* (18, 10, 30) {real, imag} */,
  {32'h3efc289c, 32'hbd83d980} /* (18, 10, 29) {real, imag} */,
  {32'h3e484c74, 32'hbf7bf720} /* (18, 10, 28) {real, imag} */,
  {32'hbf2762a4, 32'hbf0fb568} /* (18, 10, 27) {real, imag} */,
  {32'hbf612414, 32'h3f190ec4} /* (18, 10, 26) {real, imag} */,
  {32'hbf41918d, 32'h3f7c3f7c} /* (18, 10, 25) {real, imag} */,
  {32'hbe86cb98, 32'h3f44fbe8} /* (18, 10, 24) {real, imag} */,
  {32'hbf9fb85d, 32'h3e95f950} /* (18, 10, 23) {real, imag} */,
  {32'hbf816d8a, 32'hbf6b0ff0} /* (18, 10, 22) {real, imag} */,
  {32'hbecf519d, 32'hbeac2840} /* (18, 10, 21) {real, imag} */,
  {32'hbe25d8a2, 32'h3f651b94} /* (18, 10, 20) {real, imag} */,
  {32'h3f0798a0, 32'h3f326410} /* (18, 10, 19) {real, imag} */,
  {32'h3dc3ae50, 32'hbdd66700} /* (18, 10, 18) {real, imag} */,
  {32'h3e665ed0, 32'hbf2de91a} /* (18, 10, 17) {real, imag} */,
  {32'hbdaf0bd0, 32'h3df75e80} /* (18, 10, 16) {real, imag} */,
  {32'h3f8a19e3, 32'h3e926190} /* (18, 10, 15) {real, imag} */,
  {32'h3e388b1b, 32'hbf0a1c58} /* (18, 10, 14) {real, imag} */,
  {32'hbeb2266f, 32'hbf9a12aa} /* (18, 10, 13) {real, imag} */,
  {32'hbe8ba1d2, 32'h3e3e0980} /* (18, 10, 12) {real, imag} */,
  {32'hbddb8de0, 32'h3e5494c0} /* (18, 10, 11) {real, imag} */,
  {32'hbf14a2a9, 32'hbd885c7c} /* (18, 10, 10) {real, imag} */,
  {32'hbf6c8744, 32'hbdf110a0} /* (18, 10, 9) {real, imag} */,
  {32'hbf59787d, 32'h3f56c214} /* (18, 10, 8) {real, imag} */,
  {32'hbf064424, 32'h3defabc0} /* (18, 10, 7) {real, imag} */,
  {32'h3e163060, 32'hbead0dd0} /* (18, 10, 6) {real, imag} */,
  {32'hbf049155, 32'h3e389940} /* (18, 10, 5) {real, imag} */,
  {32'hbf8012e6, 32'h3f42dad8} /* (18, 10, 4) {real, imag} */,
  {32'hbe9028b0, 32'h3f3c373c} /* (18, 10, 3) {real, imag} */,
  {32'h3ecc7ebc, 32'h3f7557a0} /* (18, 10, 2) {real, imag} */,
  {32'hbf46b85c, 32'h3f8fde48} /* (18, 10, 1) {real, imag} */,
  {32'hbeada406, 32'h3e813af8} /* (18, 10, 0) {real, imag} */,
  {32'hbf11d8bc, 32'h3e95acc0} /* (18, 9, 31) {real, imag} */,
  {32'hbf3b0764, 32'hbf12fae8} /* (18, 9, 30) {real, imag} */,
  {32'hbf6a80e8, 32'hbf8d8e90} /* (18, 9, 29) {real, imag} */,
  {32'hbf8e933b, 32'hbf391b90} /* (18, 9, 28) {real, imag} */,
  {32'hbfa84a9e, 32'hbe937d20} /* (18, 9, 27) {real, imag} */,
  {32'hbf77094d, 32'h3f7a8690} /* (18, 9, 26) {real, imag} */,
  {32'hbf66a3f3, 32'h3fbee49c} /* (18, 9, 25) {real, imag} */,
  {32'hbf056c58, 32'h3fbc6b00} /* (18, 9, 24) {real, imag} */,
  {32'hbf4e0654, 32'hbec573c0} /* (18, 9, 23) {real, imag} */,
  {32'hbfb66c11, 32'hbf6a9bc8} /* (18, 9, 22) {real, imag} */,
  {32'h3e6057a8, 32'h3f329840} /* (18, 9, 21) {real, imag} */,
  {32'h3f14234f, 32'h3f9da62a} /* (18, 9, 20) {real, imag} */,
  {32'h3f4968dc, 32'h3b937000} /* (18, 9, 19) {real, imag} */,
  {32'h3ec9cf54, 32'hbf9e22a4} /* (18, 9, 18) {real, imag} */,
  {32'h3da20850, 32'hbeaba7d0} /* (18, 9, 17) {real, imag} */,
  {32'h3c7f0900, 32'h3f034150} /* (18, 9, 16) {real, imag} */,
  {32'h3fa6bf10, 32'h3f9c1c50} /* (18, 9, 15) {real, imag} */,
  {32'h3f66d48a, 32'h3e66c420} /* (18, 9, 14) {real, imag} */,
  {32'h3f17668c, 32'hbefb6890} /* (18, 9, 13) {real, imag} */,
  {32'h3ec46eb0, 32'h3f35b0e0} /* (18, 9, 12) {real, imag} */,
  {32'h3f86317d, 32'h3f2c8660} /* (18, 9, 11) {real, imag} */,
  {32'h3af7df00, 32'h3cdafb80} /* (18, 9, 10) {real, imag} */,
  {32'hbfd994a4, 32'h3ec7b200} /* (18, 9, 9) {real, imag} */,
  {32'hc00f4c7e, 32'h3f2d45f0} /* (18, 9, 8) {real, imag} */,
  {32'hbfb7ca1f, 32'hbe584840} /* (18, 9, 7) {real, imag} */,
  {32'hbf946a01, 32'hbf2f9750} /* (18, 9, 6) {real, imag} */,
  {32'hbfd2198f, 32'hbe5df140} /* (18, 9, 5) {real, imag} */,
  {32'hc002f816, 32'h3e356540} /* (18, 9, 4) {real, imag} */,
  {32'hbf0e8b9f, 32'h3f084c50} /* (18, 9, 3) {real, imag} */,
  {32'h3ea76303, 32'h3f8cce18} /* (18, 9, 2) {real, imag} */,
  {32'h3da89e90, 32'h3fd70278} /* (18, 9, 1) {real, imag} */,
  {32'hbeca5726, 32'h3f3f5870} /* (18, 9, 0) {real, imag} */,
  {32'hbf215224, 32'h3eb72c80} /* (18, 8, 31) {real, imag} */,
  {32'hbf97cf96, 32'hbf3516d8} /* (18, 8, 30) {real, imag} */,
  {32'hbfb7f406, 32'hbf2f31b8} /* (18, 8, 29) {real, imag} */,
  {32'hbf649b2e, 32'hbd87d980} /* (18, 8, 28) {real, imag} */,
  {32'hbf95e94a, 32'hbf10a340} /* (18, 8, 27) {real, imag} */,
  {32'hbf8a1b29, 32'h3f169b20} /* (18, 8, 26) {real, imag} */,
  {32'hbed53ea2, 32'h3f884814} /* (18, 8, 25) {real, imag} */,
  {32'hbd386870, 32'h3fb3a59c} /* (18, 8, 24) {real, imag} */,
  {32'hbdaf2e00, 32'h3e083c40} /* (18, 8, 23) {real, imag} */,
  {32'hbf116ba0, 32'hbee3dc20} /* (18, 8, 22) {real, imag} */,
  {32'hbf12e51e, 32'h3ec8dec0} /* (18, 8, 21) {real, imag} */,
  {32'h3f0bb8ba, 32'h3f060be8} /* (18, 8, 20) {real, imag} */,
  {32'h3fa682d0, 32'h3dd68680} /* (18, 8, 19) {real, imag} */,
  {32'h3f403398, 32'hbf59e300} /* (18, 8, 18) {real, imag} */,
  {32'h3e6efc50, 32'hbf015aa0} /* (18, 8, 17) {real, imag} */,
  {32'h3efed3c0, 32'hbd7f7100} /* (18, 8, 16) {real, imag} */,
  {32'h3fa3644e, 32'h3e272280} /* (18, 8, 15) {real, imag} */,
  {32'h3f6bebc4, 32'hbf01e1c0} /* (18, 8, 14) {real, imag} */,
  {32'h3f3219c3, 32'hbf2e2da0} /* (18, 8, 13) {real, imag} */,
  {32'h3f224808, 32'h3e5d5be0} /* (18, 8, 12) {real, imag} */,
  {32'h3fc8705c, 32'h3f331c88} /* (18, 8, 11) {real, imag} */,
  {32'h3ecece48, 32'h3d7b6800} /* (18, 8, 10) {real, imag} */,
  {32'hbfc7786a, 32'h3eb270e0} /* (18, 8, 9) {real, imag} */,
  {32'hbfae8f16, 32'h3e2a79e0} /* (18, 8, 8) {real, imag} */,
  {32'hbf468ffc, 32'hbcfff100} /* (18, 8, 7) {real, imag} */,
  {32'hbfbf3e68, 32'hbedc2250} /* (18, 8, 6) {real, imag} */,
  {32'hbf5ffb32, 32'hbe7ff2c0} /* (18, 8, 5) {real, imag} */,
  {32'hbfa9f729, 32'h3d406a00} /* (18, 8, 4) {real, imag} */,
  {32'hbf5d85cc, 32'hbe056c20} /* (18, 8, 3) {real, imag} */,
  {32'h3ed342f0, 32'h3ed51aa0} /* (18, 8, 2) {real, imag} */,
  {32'hbe5fc940, 32'h3f94ce3c} /* (18, 8, 1) {real, imag} */,
  {32'hbfb3ae6f, 32'h3f2d224c} /* (18, 8, 0) {real, imag} */,
  {32'hbe88a400, 32'hbf131558} /* (18, 7, 31) {real, imag} */,
  {32'hbf3201f0, 32'hbf00a6b0} /* (18, 7, 30) {real, imag} */,
  {32'hbfc46779, 32'h3c49d000} /* (18, 7, 29) {real, imag} */,
  {32'hbf426395, 32'hbe1009a0} /* (18, 7, 28) {real, imag} */,
  {32'hbf267dee, 32'hbf0d8ed8} /* (18, 7, 27) {real, imag} */,
  {32'hbf19efb0, 32'h3e349700} /* (18, 7, 26) {real, imag} */,
  {32'hbefed7cc, 32'h3f21cec0} /* (18, 7, 25) {real, imag} */,
  {32'hbe8b26a0, 32'h3f59a8a0} /* (18, 7, 24) {real, imag} */,
  {32'hbe529328, 32'h3ec71be0} /* (18, 7, 23) {real, imag} */,
  {32'hbda0cba0, 32'hbe3c2d60} /* (18, 7, 22) {real, imag} */,
  {32'hbe96b680, 32'hbf30e4d8} /* (18, 7, 21) {real, imag} */,
  {32'h3f177ce2, 32'hbef291a0} /* (18, 7, 20) {real, imag} */,
  {32'h3f72cf9e, 32'h3d01af00} /* (18, 7, 19) {real, imag} */,
  {32'h3f26dc90, 32'h3ec0eca0} /* (18, 7, 18) {real, imag} */,
  {32'h3eb07b48, 32'h3de71d80} /* (18, 7, 17) {real, imag} */,
  {32'h3f83d278, 32'hbdb40680} /* (18, 7, 16) {real, imag} */,
  {32'h3fa23606, 32'hbf9174d8} /* (18, 7, 15) {real, imag} */,
  {32'h3f2d4ca8, 32'hbf0b0f40} /* (18, 7, 14) {real, imag} */,
  {32'h3eb47df8, 32'hbe12e860} /* (18, 7, 13) {real, imag} */,
  {32'h3e42e678, 32'hbf158480} /* (18, 7, 12) {real, imag} */,
  {32'h3f9308c0, 32'hbec77760} /* (18, 7, 11) {real, imag} */,
  {32'hbdb34520, 32'hbeae6990} /* (18, 7, 10) {real, imag} */,
  {32'hbf29242c, 32'hbf3a3678} /* (18, 7, 9) {real, imag} */,
  {32'hbf4434a6, 32'h3d6c4580} /* (18, 7, 8) {real, imag} */,
  {32'hbf420311, 32'hbe791f60} /* (18, 7, 7) {real, imag} */,
  {32'hbfa481d9, 32'hbf259478} /* (18, 7, 6) {real, imag} */,
  {32'hbf0aa23e, 32'hbeee55c0} /* (18, 7, 5) {real, imag} */,
  {32'hbf6f8614, 32'h3eca20c0} /* (18, 7, 4) {real, imag} */,
  {32'hbebe6828, 32'h3e93a520} /* (18, 7, 3) {real, imag} */,
  {32'h3e067f90, 32'h3deb8000} /* (18, 7, 2) {real, imag} */,
  {32'hbf8090f8, 32'h3f289910} /* (18, 7, 1) {real, imag} */,
  {32'hbf88da0c, 32'h3e8e1af0} /* (18, 7, 0) {real, imag} */,
  {32'hbf473c46, 32'hbeb46160} /* (18, 6, 31) {real, imag} */,
  {32'hbee4bbec, 32'hbeb9d4b0} /* (18, 6, 30) {real, imag} */,
  {32'hbf05bf5e, 32'h3edfa040} /* (18, 6, 29) {real, imag} */,
  {32'hbf292db7, 32'h3e9225e0} /* (18, 6, 28) {real, imag} */,
  {32'hbf0e774c, 32'h3ee84200} /* (18, 6, 27) {real, imag} */,
  {32'hbef65320, 32'h3f23d598} /* (18, 6, 26) {real, imag} */,
  {32'hbed100a0, 32'h3f4d2660} /* (18, 6, 25) {real, imag} */,
  {32'hbe707530, 32'h3ed53f40} /* (18, 6, 24) {real, imag} */,
  {32'hbe4c0500, 32'h3f5879b0} /* (18, 6, 23) {real, imag} */,
  {32'hbd704fc0, 32'h3f024638} /* (18, 6, 22) {real, imag} */,
  {32'hbe909738, 32'hbe713800} /* (18, 6, 21) {real, imag} */,
  {32'hbe817014, 32'h3dcd78a0} /* (18, 6, 20) {real, imag} */,
  {32'h3f13bc52, 32'h3e97b510} /* (18, 6, 19) {real, imag} */,
  {32'h3f824bec, 32'h3f992350} /* (18, 6, 18) {real, imag} */,
  {32'h3f7ac2fd, 32'h3e4e01a0} /* (18, 6, 17) {real, imag} */,
  {32'h3f62303a, 32'hbe1a0f00} /* (18, 6, 16) {real, imag} */,
  {32'h3eae0860, 32'hbe90e000} /* (18, 6, 15) {real, imag} */,
  {32'h3ed3a0f0, 32'h3db22680} /* (18, 6, 14) {real, imag} */,
  {32'h3f381e70, 32'hbde21fc0} /* (18, 6, 13) {real, imag} */,
  {32'h3f4eacec, 32'hbf6ce8a8} /* (18, 6, 12) {real, imag} */,
  {32'h3f4c1cb0, 32'hbec6ce50} /* (18, 6, 11) {real, imag} */,
  {32'h3d3dd9b0, 32'hbf1394e0} /* (18, 6, 10) {real, imag} */,
  {32'h3f4dfc56, 32'hbf2a7400} /* (18, 6, 9) {real, imag} */,
  {32'h3f56efbe, 32'h3e01a980} /* (18, 6, 8) {real, imag} */,
  {32'hbdbf8628, 32'hbf828c98} /* (18, 6, 7) {real, imag} */,
  {32'hbf6bbc48, 32'hbfef5548} /* (18, 6, 6) {real, imag} */,
  {32'hbf5783b4, 32'hbfa3a9e8} /* (18, 6, 5) {real, imag} */,
  {32'hbf9353f2, 32'h3ecdd640} /* (18, 6, 4) {real, imag} */,
  {32'hbee3ba78, 32'h3f924764} /* (18, 6, 3) {real, imag} */,
  {32'hbe6dd000, 32'hbc906c00} /* (18, 6, 2) {real, imag} */,
  {32'h3da4bc80, 32'hbf3a93e8} /* (18, 6, 1) {real, imag} */,
  {32'hbdb78ba0, 32'hbea44588} /* (18, 6, 0) {real, imag} */,
  {32'hbf432a44, 32'hbf322964} /* (18, 5, 31) {real, imag} */,
  {32'hbf081dc0, 32'hbf036d50} /* (18, 5, 30) {real, imag} */,
  {32'hbf4ba796, 32'h3eb41aa0} /* (18, 5, 29) {real, imag} */,
  {32'hbfa988e9, 32'h3f2ddd00} /* (18, 5, 28) {real, imag} */,
  {32'hbf980963, 32'h3fa5e7b8} /* (18, 5, 27) {real, imag} */,
  {32'hbf63674c, 32'h3f999c88} /* (18, 5, 26) {real, imag} */,
  {32'hbf0a40fa, 32'h3f70ebf0} /* (18, 5, 25) {real, imag} */,
  {32'hbf26ad62, 32'h3f447ab0} /* (18, 5, 24) {real, imag} */,
  {32'hbf5b663c, 32'h3f790de0} /* (18, 5, 23) {real, imag} */,
  {32'hbf07ee50, 32'h3dc3af00} /* (18, 5, 22) {real, imag} */,
  {32'hbf401143, 32'h3d7c8a80} /* (18, 5, 21) {real, imag} */,
  {32'hbf99f51a, 32'h3d9ab4c0} /* (18, 5, 20) {real, imag} */,
  {32'hbe95f652, 32'h3d7ce780} /* (18, 5, 19) {real, imag} */,
  {32'h3f236356, 32'h3e6ffe60} /* (18, 5, 18) {real, imag} */,
  {32'h3ef2c294, 32'hbe529020} /* (18, 5, 17) {real, imag} */,
  {32'hbb840040, 32'h3b2aa000} /* (18, 5, 16) {real, imag} */,
  {32'h3d4f2400, 32'h3e4b64a0} /* (18, 5, 15) {real, imag} */,
  {32'h3e88971c, 32'h3f6e9708} /* (18, 5, 14) {real, imag} */,
  {32'h3f3044b2, 32'hbee83520} /* (18, 5, 13) {real, imag} */,
  {32'h3f292f80, 32'hbf26a5f0} /* (18, 5, 12) {real, imag} */,
  {32'h3ec5fc90, 32'h3db29400} /* (18, 5, 11) {real, imag} */,
  {32'h3d7a3520, 32'h3ecfa290} /* (18, 5, 10) {real, imag} */,
  {32'h3f1b1119, 32'h3e989130} /* (18, 5, 9) {real, imag} */,
  {32'h3fa8275f, 32'h3f042c54} /* (18, 5, 8) {real, imag} */,
  {32'h3f1e733b, 32'hbf511b88} /* (18, 5, 7) {real, imag} */,
  {32'h3ec11d49, 32'hbfb6d13d} /* (18, 5, 6) {real, imag} */,
  {32'hbde3e310, 32'hbf1da228} /* (18, 5, 5) {real, imag} */,
  {32'hbf874383, 32'hbeeb02e0} /* (18, 5, 4) {real, imag} */,
  {32'hbeac9132, 32'h3ef19b80} /* (18, 5, 3) {real, imag} */,
  {32'hbe05f300, 32'hbe83e040} /* (18, 5, 2) {real, imag} */,
  {32'hbf480648, 32'hbf293060} /* (18, 5, 1) {real, imag} */,
  {32'hbed918c0, 32'hbeebe500} /* (18, 5, 0) {real, imag} */,
  {32'hbea299a8, 32'hbe961218} /* (18, 4, 31) {real, imag} */,
  {32'hbebeebc0, 32'h3f104380} /* (18, 4, 30) {real, imag} */,
  {32'hbee1a798, 32'h3f3071f0} /* (18, 4, 29) {real, imag} */,
  {32'hbf58b962, 32'h3f3febb0} /* (18, 4, 28) {real, imag} */,
  {32'hbf148d46, 32'h3f815d28} /* (18, 4, 27) {real, imag} */,
  {32'hbf555ad5, 32'h3f23dcc0} /* (18, 4, 26) {real, imag} */,
  {32'hbf592d0c, 32'h3e8bc3c0} /* (18, 4, 25) {real, imag} */,
  {32'hbf9abb86, 32'h3e86a240} /* (18, 4, 24) {real, imag} */,
  {32'hbe715378, 32'h3e810c00} /* (18, 4, 23) {real, imag} */,
  {32'hbec7a140, 32'h3e1d3840} /* (18, 4, 22) {real, imag} */,
  {32'hbf712a44, 32'h3e594f00} /* (18, 4, 21) {real, imag} */,
  {32'hbfbd6e28, 32'hbf9351e8} /* (18, 4, 20) {real, imag} */,
  {32'hbf417868, 32'hbfbaef54} /* (18, 4, 19) {real, imag} */,
  {32'hbd8e77c0, 32'hbf8bc860} /* (18, 4, 18) {real, imag} */,
  {32'hbe691360, 32'hbf70b020} /* (18, 4, 17) {real, imag} */,
  {32'hbf3dc18e, 32'hbe973860} /* (18, 4, 16) {real, imag} */,
  {32'h3e768790, 32'h3e87e9d8} /* (18, 4, 15) {real, imag} */,
  {32'h3f367492, 32'h3f8dafb8} /* (18, 4, 14) {real, imag} */,
  {32'h3e43fbac, 32'h3e8e9a80} /* (18, 4, 13) {real, imag} */,
  {32'h3e039f20, 32'h3d72de80} /* (18, 4, 12) {real, imag} */,
  {32'h3f1bccdc, 32'h3e948660} /* (18, 4, 11) {real, imag} */,
  {32'h3e760920, 32'h3e9328a0} /* (18, 4, 10) {real, imag} */,
  {32'hbc40ef80, 32'hbdd856c0} /* (18, 4, 9) {real, imag} */,
  {32'h3ea16b2c, 32'h3b21e000} /* (18, 4, 8) {real, imag} */,
  {32'h3fa37061, 32'h3d988b40} /* (18, 4, 7) {real, imag} */,
  {32'h3fdd3158, 32'hbead0d00} /* (18, 4, 6) {real, imag} */,
  {32'h3ecc9c65, 32'hbed2e348} /* (18, 4, 5) {real, imag} */,
  {32'hbf822fde, 32'hbf066ea8} /* (18, 4, 4) {real, imag} */,
  {32'hbf186628, 32'hbe53b500} /* (18, 4, 3) {real, imag} */,
  {32'hbf00d8e4, 32'h3df64980} /* (18, 4, 2) {real, imag} */,
  {32'hbf5e09a8, 32'hbd1bcc00} /* (18, 4, 1) {real, imag} */,
  {32'hbef7da58, 32'hbd83ee20} /* (18, 4, 0) {real, imag} */,
  {32'hbf3b4f1e, 32'h3e4d1660} /* (18, 3, 31) {real, imag} */,
  {32'hbf27249c, 32'h3e259680} /* (18, 3, 30) {real, imag} */,
  {32'h3e68b470, 32'hbecd8420} /* (18, 3, 29) {real, imag} */,
  {32'hbec32853, 32'hbe2febc0} /* (18, 3, 28) {real, imag} */,
  {32'h3e9b701c, 32'h3dd74d80} /* (18, 3, 27) {real, imag} */,
  {32'hbe45f8b8, 32'h3cd67a00} /* (18, 3, 26) {real, imag} */,
  {32'hbf547da8, 32'hbe28dce0} /* (18, 3, 25) {real, imag} */,
  {32'hbfae719c, 32'hbf5a7b40} /* (18, 3, 24) {real, imag} */,
  {32'hbe9f51f4, 32'hbea0e310} /* (18, 3, 23) {real, imag} */,
  {32'hbf010888, 32'h3e8d3040} /* (18, 3, 22) {real, imag} */,
  {32'hbe80652c, 32'h3ecbef50} /* (18, 3, 21) {real, imag} */,
  {32'hbf20566c, 32'h3d8122c0} /* (18, 3, 20) {real, imag} */,
  {32'hbf3cc404, 32'hbf9620a0} /* (18, 3, 19) {real, imag} */,
  {32'hbe2e7ee0, 32'hbf90c898} /* (18, 3, 18) {real, imag} */,
  {32'hbf024608, 32'hbef6c6c0} /* (18, 3, 17) {real, imag} */,
  {32'hbf9afd14, 32'h3e9c9b90} /* (18, 3, 16) {real, imag} */,
  {32'hbe15904c, 32'h3e8cfbe8} /* (18, 3, 15) {real, imag} */,
  {32'h3fa707a2, 32'h3f0ab7e8} /* (18, 3, 14) {real, imag} */,
  {32'h3eae3524, 32'h3f1e86a0} /* (18, 3, 13) {real, imag} */,
  {32'h3c2ed180, 32'h3e97ce40} /* (18, 3, 12) {real, imag} */,
  {32'h3ed1e888, 32'h3f8601c8} /* (18, 3, 11) {real, imag} */,
  {32'h3ae9f800, 32'h3ebe1080} /* (18, 3, 10) {real, imag} */,
  {32'hbdca3530, 32'hbdcba380} /* (18, 3, 9) {real, imag} */,
  {32'hbe87da70, 32'hbe7dcf40} /* (18, 3, 8) {real, imag} */,
  {32'h3edfe940, 32'hbecd4bc0} /* (18, 3, 7) {real, imag} */,
  {32'h3fad27ff, 32'hbf8b04e8} /* (18, 3, 6) {real, imag} */,
  {32'h3f1fbfee, 32'hbef10f04} /* (18, 3, 5) {real, imag} */,
  {32'hbf3f50e6, 32'h3e9b9890} /* (18, 3, 4) {real, imag} */,
  {32'hbf55f488, 32'h3f8c1d68} /* (18, 3, 3) {real, imag} */,
  {32'hbe60ba68, 32'h3fcc69f8} /* (18, 3, 2) {real, imag} */,
  {32'hbeaecb80, 32'h3f112340} /* (18, 3, 1) {real, imag} */,
  {32'hbeed84b4, 32'hbe5611c0} /* (18, 3, 0) {real, imag} */,
  {32'hbe570e5c, 32'h3df18c80} /* (18, 2, 31) {real, imag} */,
  {32'hbcc6ed80, 32'hbce28400} /* (18, 2, 30) {real, imag} */,
  {32'h3c089800, 32'hbf796030} /* (18, 2, 29) {real, imag} */,
  {32'hbf71c5a8, 32'hbf65a628} /* (18, 2, 28) {real, imag} */,
  {32'hbf8399ca, 32'hbea880a0} /* (18, 2, 27) {real, imag} */,
  {32'hbf4a0863, 32'hbda12140} /* (18, 2, 26) {real, imag} */,
  {32'hbf421fbc, 32'hbe4dc3a0} /* (18, 2, 25) {real, imag} */,
  {32'hbf9acf68, 32'hbe9d5ec0} /* (18, 2, 24) {real, imag} */,
  {32'hbf8a3f0a, 32'hbe56b040} /* (18, 2, 23) {real, imag} */,
  {32'hbfa103b4, 32'hbf66dd60} /* (18, 2, 22) {real, imag} */,
  {32'hbf46b0ea, 32'hbe979100} /* (18, 2, 21) {real, imag} */,
  {32'hbf753f00, 32'h3f2b6e10} /* (18, 2, 20) {real, imag} */,
  {32'hbf00e1e8, 32'hbe4b03c0} /* (18, 2, 19) {real, imag} */,
  {32'h3ef49580, 32'hbf5ce078} /* (18, 2, 18) {real, imag} */,
  {32'hbe03ca90, 32'hbf8850fc} /* (18, 2, 17) {real, imag} */,
  {32'hbf9f5e01, 32'hbe999210} /* (18, 2, 16) {real, imag} */,
  {32'h3bb23a00, 32'hbf147598} /* (18, 2, 15) {real, imag} */,
  {32'h3fcd6cf4, 32'hbd11c980} /* (18, 2, 14) {real, imag} */,
  {32'h3f42b08a, 32'hbe6791c0} /* (18, 2, 13) {real, imag} */,
  {32'h3f28d25a, 32'hbebac600} /* (18, 2, 12) {real, imag} */,
  {32'h3f54e7d6, 32'h3f81e1e8} /* (18, 2, 11) {real, imag} */,
  {32'h3eb55af8, 32'h3ee39c50} /* (18, 2, 10) {real, imag} */,
  {32'h3e8b8d50, 32'hbe8f00f0} /* (18, 2, 9) {real, imag} */,
  {32'h3eab63e0, 32'hbf21ce58} /* (18, 2, 8) {real, imag} */,
  {32'h3ea6e950, 32'hbee76d80} /* (18, 2, 7) {real, imag} */,
  {32'h3f17fd14, 32'hbee1c220} /* (18, 2, 6) {real, imag} */,
  {32'hbf58e496, 32'hbf58c6e9} /* (18, 2, 5) {real, imag} */,
  {32'hbf102578, 32'h3eb309a0} /* (18, 2, 4) {real, imag} */,
  {32'hbf378c91, 32'h3fc2f348} /* (18, 2, 3) {real, imag} */,
  {32'hbeb58770, 32'h3eff1aa0} /* (18, 2, 2) {real, imag} */,
  {32'h3eabe5f0, 32'h3e11f1e0} /* (18, 2, 1) {real, imag} */,
  {32'hbe0806d8, 32'hbe81ee88} /* (18, 2, 0) {real, imag} */,
  {32'h3e9df970, 32'hbe02bdf0} /* (18, 1, 31) {real, imag} */,
  {32'h3e611310, 32'hbe28b740} /* (18, 1, 30) {real, imag} */,
  {32'h3e74d9d0, 32'hbf418878} /* (18, 1, 29) {real, imag} */,
  {32'hbf4b4386, 32'hbf57ab50} /* (18, 1, 28) {real, imag} */,
  {32'hbfbef6f5, 32'hbf98b7c8} /* (18, 1, 27) {real, imag} */,
  {32'hbf7a24b1, 32'hbf591ad0} /* (18, 1, 26) {real, imag} */,
  {32'hbe9a0e98, 32'hbea9e100} /* (18, 1, 25) {real, imag} */,
  {32'hbf836eaf, 32'h3eca6770} /* (18, 1, 24) {real, imag} */,
  {32'hbf4ca9be, 32'hbe76b140} /* (18, 1, 23) {real, imag} */,
  {32'hbeeea0ac, 32'hbfa48b6c} /* (18, 1, 22) {real, imag} */,
  {32'hbf0c4477, 32'hbf6d4d90} /* (18, 1, 21) {real, imag} */,
  {32'hbf68a752, 32'hbe9196b0} /* (18, 1, 20) {real, imag} */,
  {32'h3eae3578, 32'hbd430c00} /* (18, 1, 19) {real, imag} */,
  {32'h3f9feff0, 32'hbe5e6fc0} /* (18, 1, 18) {real, imag} */,
  {32'h3f27d180, 32'hbeeede40} /* (18, 1, 17) {real, imag} */,
  {32'hbeb20d56, 32'hbf200538} /* (18, 1, 16) {real, imag} */,
  {32'h3f1eff62, 32'hbf8508ac} /* (18, 1, 15) {real, imag} */,
  {32'h3f86825a, 32'hbf733178} /* (18, 1, 14) {real, imag} */,
  {32'h3ea78fc8, 32'hbf57b9b0} /* (18, 1, 13) {real, imag} */,
  {32'h3f7dfce0, 32'h3ef497d0} /* (18, 1, 12) {real, imag} */,
  {32'h3e9f8b80, 32'h3fbfa868} /* (18, 1, 11) {real, imag} */,
  {32'h3eeff43c, 32'h3e6df100} /* (18, 1, 10) {real, imag} */,
  {32'h3f29fa98, 32'hbf1672c0} /* (18, 1, 9) {real, imag} */,
  {32'h3eca1ed4, 32'hbc03f000} /* (18, 1, 8) {real, imag} */,
  {32'h3eb018a8, 32'h3e4a9f00} /* (18, 1, 7) {real, imag} */,
  {32'h3fc2cb1f, 32'hbe456540} /* (18, 1, 6) {real, imag} */,
  {32'h3d826a08, 32'hbf23baf9} /* (18, 1, 5) {real, imag} */,
  {32'h3e091c00, 32'h3f56fc78} /* (18, 1, 4) {real, imag} */,
  {32'hbe46ffb0, 32'h3f019f30} /* (18, 1, 3) {real, imag} */,
  {32'hbe83433c, 32'hbf2c9cd8} /* (18, 1, 2) {real, imag} */,
  {32'h3f085270, 32'hbf6d09d0} /* (18, 1, 1) {real, imag} */,
  {32'h3ef4c168, 32'hbed16760} /* (18, 1, 0) {real, imag} */,
  {32'h3ee3e2a0, 32'hbeb1e70c} /* (18, 0, 31) {real, imag} */,
  {32'hbe119240, 32'hbe6b9c70} /* (18, 0, 30) {real, imag} */,
  {32'hbec821a4, 32'hbd970320} /* (18, 0, 29) {real, imag} */,
  {32'hbec90634, 32'hbdc568c0} /* (18, 0, 28) {real, imag} */,
  {32'hbf5316d6, 32'hbf4b118c} /* (18, 0, 27) {real, imag} */,
  {32'hbec46a6e, 32'hbec30010} /* (18, 0, 26) {real, imag} */,
  {32'hbde4cb30, 32'hbdd2a380} /* (18, 0, 25) {real, imag} */,
  {32'hbf6ae3fc, 32'h3c33d900} /* (18, 0, 24) {real, imag} */,
  {32'hbf0bed7a, 32'hbdc8cac0} /* (18, 0, 23) {real, imag} */,
  {32'hbddf77b0, 32'hbeaa1540} /* (18, 0, 22) {real, imag} */,
  {32'hbec3900a, 32'hbeb17460} /* (18, 0, 21) {real, imag} */,
  {32'hbede7c46, 32'hbea3bec0} /* (18, 0, 20) {real, imag} */,
  {32'h3e710768, 32'hbeae2098} /* (18, 0, 19) {real, imag} */,
  {32'h3e531960, 32'hbeeb0b90} /* (18, 0, 18) {real, imag} */,
  {32'hbe1c096c, 32'hbe96b160} /* (18, 0, 17) {real, imag} */,
  {32'h3e2da850, 32'hbed54a24} /* (18, 0, 16) {real, imag} */,
  {32'h3f517eba, 32'hbf266d20} /* (18, 0, 15) {real, imag} */,
  {32'h3ee4a9ae, 32'hbf307270} /* (18, 0, 14) {real, imag} */,
  {32'h3ec8c67e, 32'hbe9dcca0} /* (18, 0, 13) {real, imag} */,
  {32'h3eaf07a0, 32'h3e4d4e00} /* (18, 0, 12) {real, imag} */,
  {32'hbe14fbe8, 32'h3f4ac70c} /* (18, 0, 11) {real, imag} */,
  {32'h3f1572fb, 32'h3f15ee60} /* (18, 0, 10) {real, imag} */,
  {32'h3e08f010, 32'h3d1cc140} /* (18, 0, 9) {real, imag} */,
  {32'hbe3e11f8, 32'h3e2f5e60} /* (18, 0, 8) {real, imag} */,
  {32'h3e3bcf00, 32'hbdd05d00} /* (18, 0, 7) {real, imag} */,
  {32'h3f96357f, 32'hbe673d60} /* (18, 0, 6) {real, imag} */,
  {32'h3e0122c6, 32'hbe9d1076} /* (18, 0, 5) {real, imag} */,
  {32'hbee4d374, 32'h3e7d2e90} /* (18, 0, 4) {real, imag} */,
  {32'hbed26a28, 32'hbe9f80f8} /* (18, 0, 3) {real, imag} */,
  {32'hbf12d10d, 32'hbf1efa4c} /* (18, 0, 2) {real, imag} */,
  {32'hbe40f47c, 32'hbebc4100} /* (18, 0, 1) {real, imag} */,
  {32'h3e980288, 32'hbe058140} /* (18, 0, 0) {real, imag} */,
  {32'h3e2729d2, 32'h3e6560e0} /* (17, 31, 31) {real, imag} */,
  {32'h3eb8c64d, 32'h3dc1ffc0} /* (17, 31, 30) {real, imag} */,
  {32'h3f0728d1, 32'hbea432f8} /* (17, 31, 29) {real, imag} */,
  {32'h3e9e435a, 32'hbf58f5b0} /* (17, 31, 28) {real, imag} */,
  {32'h3e56299a, 32'hbe715ca0} /* (17, 31, 27) {real, imag} */,
  {32'h3e76cdea, 32'h3f045f84} /* (17, 31, 26) {real, imag} */,
  {32'h3e9001c4, 32'hbe487b30} /* (17, 31, 25) {real, imag} */,
  {32'h3d817120, 32'hbe3827c0} /* (17, 31, 24) {real, imag} */,
  {32'h3f1eb7be, 32'hbd8428c0} /* (17, 31, 23) {real, imag} */,
  {32'h3f12515b, 32'hbf34fee0} /* (17, 31, 22) {real, imag} */,
  {32'h3d9fb2fc, 32'hbed5c568} /* (17, 31, 21) {real, imag} */,
  {32'hbdf72b80, 32'hbf344d26} /* (17, 31, 20) {real, imag} */,
  {32'h3e4c9abc, 32'hbd247d00} /* (17, 31, 19) {real, imag} */,
  {32'hbdf53020, 32'hbe29eef8} /* (17, 31, 18) {real, imag} */,
  {32'hbe549749, 32'hbf3489b8} /* (17, 31, 17) {real, imag} */,
  {32'hbf097ff7, 32'hbe08a460} /* (17, 31, 16) {real, imag} */,
  {32'hbd8ef9f8, 32'hbe952928} /* (17, 31, 15) {real, imag} */,
  {32'hbe04856c, 32'hbe6d51e0} /* (17, 31, 14) {real, imag} */,
  {32'hbed9903e, 32'hbf547a74} /* (17, 31, 13) {real, imag} */,
  {32'hbf03553e, 32'hbf34992a} /* (17, 31, 12) {real, imag} */,
  {32'hbec967c6, 32'hbe979d88} /* (17, 31, 11) {real, imag} */,
  {32'hbe3fdb49, 32'hbe2c71e0} /* (17, 31, 10) {real, imag} */,
  {32'hbd6b4e18, 32'hbea8e704} /* (17, 31, 9) {real, imag} */,
  {32'h3f0bd69d, 32'hbf0e6edc} /* (17, 31, 8) {real, imag} */,
  {32'hbe705dc8, 32'h3f4a36d8} /* (17, 31, 7) {real, imag} */,
  {32'h3e0f58c4, 32'h3ef41c50} /* (17, 31, 6) {real, imag} */,
  {32'h3f4ca65f, 32'h3e41cba0} /* (17, 31, 5) {real, imag} */,
  {32'h3f277a67, 32'hbe1e3650} /* (17, 31, 4) {real, imag} */,
  {32'h3f55db1a, 32'hbe6eefc0} /* (17, 31, 3) {real, imag} */,
  {32'h3dab4c4e, 32'hbd6d7800} /* (17, 31, 2) {real, imag} */,
  {32'h3d7e4940, 32'h3e20a700} /* (17, 31, 1) {real, imag} */,
  {32'h3ee38eea, 32'h3ebe8e0c} /* (17, 31, 0) {real, imag} */,
  {32'h3e0f2c4c, 32'hbdb82de0} /* (17, 30, 31) {real, imag} */,
  {32'h3dd0c530, 32'hbeb51c30} /* (17, 30, 30) {real, imag} */,
  {32'h3f67fa14, 32'hbf07bb10} /* (17, 30, 29) {real, imag} */,
  {32'h3f272664, 32'hbfab042c} /* (17, 30, 28) {real, imag} */,
  {32'h3f21859a, 32'hbf02818c} /* (17, 30, 27) {real, imag} */,
  {32'h3e0f952a, 32'h3e74f400} /* (17, 30, 26) {real, imag} */,
  {32'h3d868c1c, 32'hbebfba70} /* (17, 30, 25) {real, imag} */,
  {32'h3dc7905a, 32'h3efa3d80} /* (17, 30, 24) {real, imag} */,
  {32'h3e960de4, 32'h3efaf560} /* (17, 30, 23) {real, imag} */,
  {32'h3f3f3e59, 32'hbf912a8c} /* (17, 30, 22) {real, imag} */,
  {32'h3e815bf4, 32'hbf2a9998} /* (17, 30, 21) {real, imag} */,
  {32'h3d8af1c6, 32'hbe644e80} /* (17, 30, 20) {real, imag} */,
  {32'h3f57c03a, 32'h3e70fc00} /* (17, 30, 19) {real, imag} */,
  {32'h3e93adf6, 32'h3d0cc600} /* (17, 30, 18) {real, imag} */,
  {32'hbec84ef6, 32'hbf5d0fa4} /* (17, 30, 17) {real, imag} */,
  {32'hbea8e087, 32'hbeca8880} /* (17, 30, 16) {real, imag} */,
  {32'h3d35b0f0, 32'hbe61f0e0} /* (17, 30, 15) {real, imag} */,
  {32'hbd24aac0, 32'h3a6fa000} /* (17, 30, 14) {real, imag} */,
  {32'hbe9d7f14, 32'hbf3248dc} /* (17, 30, 13) {real, imag} */,
  {32'hbf443d0d, 32'hbf146c10} /* (17, 30, 12) {real, imag} */,
  {32'hbef2c3fe, 32'hbf1e36ae} /* (17, 30, 11) {real, imag} */,
  {32'h3d191760, 32'hbeeaa688} /* (17, 30, 10) {real, imag} */,
  {32'h3f08e918, 32'hbec72cf8} /* (17, 30, 9) {real, imag} */,
  {32'h3eba66e0, 32'hbf7862c8} /* (17, 30, 8) {real, imag} */,
  {32'h3def15f0, 32'h3edc5298} /* (17, 30, 7) {real, imag} */,
  {32'h3f8f0353, 32'h3f311498} /* (17, 30, 6) {real, imag} */,
  {32'h3f8371c6, 32'h3e0e0ea0} /* (17, 30, 5) {real, imag} */,
  {32'h3f904a84, 32'h3e281060} /* (17, 30, 4) {real, imag} */,
  {32'h3f3f7bf1, 32'hbe91db58} /* (17, 30, 3) {real, imag} */,
  {32'hbf0e514c, 32'h3db08500} /* (17, 30, 2) {real, imag} */,
  {32'hbeb723de, 32'hbc19c400} /* (17, 30, 1) {real, imag} */,
  {32'h3e65df52, 32'h3e929234} /* (17, 30, 0) {real, imag} */,
  {32'hbefd999e, 32'h3e5d1b00} /* (17, 29, 31) {real, imag} */,
  {32'hbce06500, 32'hbed8c150} /* (17, 29, 30) {real, imag} */,
  {32'h3f06356a, 32'hbf47a050} /* (17, 29, 29) {real, imag} */,
  {32'h3eda9c28, 32'hbe88fa08} /* (17, 29, 28) {real, imag} */,
  {32'h3f1edba2, 32'hbeefbc18} /* (17, 29, 27) {real, imag} */,
  {32'h3d29f3f0, 32'hbec8eed8} /* (17, 29, 26) {real, imag} */,
  {32'h3e6547c8, 32'h3cafaf80} /* (17, 29, 25) {real, imag} */,
  {32'hbe590700, 32'h3f04de30} /* (17, 29, 24) {real, imag} */,
  {32'hbbfcae00, 32'h3d5ba3c0} /* (17, 29, 23) {real, imag} */,
  {32'h3f6db1b6, 32'hbf1acc74} /* (17, 29, 22) {real, imag} */,
  {32'h3f68448c, 32'hbed21590} /* (17, 29, 21) {real, imag} */,
  {32'h3f77b094, 32'hbe5b5cb0} /* (17, 29, 20) {real, imag} */,
  {32'h3f361796, 32'hbb6d2000} /* (17, 29, 19) {real, imag} */,
  {32'h3f9221c3, 32'hbe957190} /* (17, 29, 18) {real, imag} */,
  {32'h3ed7fd78, 32'hbf3ca5ac} /* (17, 29, 17) {real, imag} */,
  {32'hbdbe50d0, 32'hbf38dffc} /* (17, 29, 16) {real, imag} */,
  {32'hbf0a06b3, 32'hbf2db084} /* (17, 29, 15) {real, imag} */,
  {32'hbe598200, 32'hbc4a1c00} /* (17, 29, 14) {real, imag} */,
  {32'h3eb39750, 32'hbc4f3200} /* (17, 29, 13) {real, imag} */,
  {32'hbf5faf80, 32'hbe3d3d90} /* (17, 29, 12) {real, imag} */,
  {32'hbf756b3a, 32'hbe926730} /* (17, 29, 11) {real, imag} */,
  {32'hbec09660, 32'hbe532ea4} /* (17, 29, 10) {real, imag} */,
  {32'h3e9289a6, 32'hbda201a0} /* (17, 29, 9) {real, imag} */,
  {32'hbd881820, 32'hbf0b64c8} /* (17, 29, 8) {real, imag} */,
  {32'h3d9160b8, 32'hbeb2e260} /* (17, 29, 7) {real, imag} */,
  {32'h3f563f16, 32'hbd098700} /* (17, 29, 6) {real, imag} */,
  {32'h3f1b0b33, 32'h3d8f1420} /* (17, 29, 5) {real, imag} */,
  {32'h3f40ddda, 32'hbe3e63c0} /* (17, 29, 4) {real, imag} */,
  {32'h3eb1e108, 32'hbd8790a0} /* (17, 29, 3) {real, imag} */,
  {32'hbf052816, 32'h3f31a690} /* (17, 29, 2) {real, imag} */,
  {32'hbef5a36c, 32'hbe63f000} /* (17, 29, 1) {real, imag} */,
  {32'hbec177d8, 32'hbec07840} /* (17, 29, 0) {real, imag} */,
  {32'hbedafbc8, 32'h3ef1ae18} /* (17, 28, 31) {real, imag} */,
  {32'hbeb8b6b8, 32'hbf00aa08} /* (17, 28, 30) {real, imag} */,
  {32'hbc63a100, 32'hbf17cee8} /* (17, 28, 29) {real, imag} */,
  {32'h3cc143c0, 32'h3f2f12d8} /* (17, 28, 28) {real, imag} */,
  {32'h3f161107, 32'h3d946ae0} /* (17, 28, 27) {real, imag} */,
  {32'h3ed6e5b0, 32'hbf88929a} /* (17, 28, 26) {real, imag} */,
  {32'h3f7d58d4, 32'hbd2fc680} /* (17, 28, 25) {real, imag} */,
  {32'h3f4de884, 32'h3dc42100} /* (17, 28, 24) {real, imag} */,
  {32'h3f61bba2, 32'hbe8a2360} /* (17, 28, 23) {real, imag} */,
  {32'h3f825be6, 32'h3c400c00} /* (17, 28, 22) {real, imag} */,
  {32'h3f68fdf7, 32'hbec65748} /* (17, 28, 21) {real, imag} */,
  {32'h3f8106d6, 32'hbf356e6c} /* (17, 28, 20) {real, imag} */,
  {32'h3f187358, 32'hbe8efb10} /* (17, 28, 19) {real, imag} */,
  {32'h3f559ea2, 32'hbecca7b0} /* (17, 28, 18) {real, imag} */,
  {32'h3f318cfd, 32'hbf033eb0} /* (17, 28, 17) {real, imag} */,
  {32'h3e0cf18a, 32'hbeb8ddb0} /* (17, 28, 16) {real, imag} */,
  {32'hbf6fa6a0, 32'hbf0bc090} /* (17, 28, 15) {real, imag} */,
  {32'hbf2b96b0, 32'hbc87e500} /* (17, 28, 14) {real, imag} */,
  {32'hbdba5e30, 32'h3f158ff8} /* (17, 28, 13) {real, imag} */,
  {32'hbf44c7a3, 32'h3f413bac} /* (17, 28, 12) {real, imag} */,
  {32'hbee99cce, 32'h3f02e188} /* (17, 28, 11) {real, imag} */,
  {32'hbe2f4d28, 32'h3e5dff2c} /* (17, 28, 10) {real, imag} */,
  {32'hbeeae198, 32'hbd4a7b80} /* (17, 28, 9) {real, imag} */,
  {32'h3d60f220, 32'h3da927a0} /* (17, 28, 8) {real, imag} */,
  {32'h3e744b54, 32'h3e967848} /* (17, 28, 7) {real, imag} */,
  {32'h3e8e8730, 32'h3dc262c0} /* (17, 28, 6) {real, imag} */,
  {32'h3e92d20d, 32'hbe9e8e40} /* (17, 28, 5) {real, imag} */,
  {32'h3d158974, 32'hbf0432e8} /* (17, 28, 4) {real, imag} */,
  {32'h3e260478, 32'h3e992440} /* (17, 28, 3) {real, imag} */,
  {32'hbed32aec, 32'h3e8fd5a0} /* (17, 28, 2) {real, imag} */,
  {32'hbe565cc0, 32'hbeaa7260} /* (17, 28, 1) {real, imag} */,
  {32'hbe0d27a0, 32'hbe983850} /* (17, 28, 0) {real, imag} */,
  {32'hbe895b70, 32'hbdc4c740} /* (17, 27, 31) {real, imag} */,
  {32'hbf3b7648, 32'hbf0421b8} /* (17, 27, 30) {real, imag} */,
  {32'h3e3dae78, 32'hbee4bb10} /* (17, 27, 29) {real, imag} */,
  {32'h3e5e6e8d, 32'h3ebe0430} /* (17, 27, 28) {real, imag} */,
  {32'hbea0cb63, 32'h3dc0bc60} /* (17, 27, 27) {real, imag} */,
  {32'hbe2e9ffc, 32'hbf309328} /* (17, 27, 26) {real, imag} */,
  {32'h3f09cb34, 32'h3e3219c0} /* (17, 27, 25) {real, imag} */,
  {32'h3f10059c, 32'hbebf2ef0} /* (17, 27, 24) {real, imag} */,
  {32'h3efa8c57, 32'hbf0e9df8} /* (17, 27, 23) {real, imag} */,
  {32'h3d9be758, 32'h3e15b730} /* (17, 27, 22) {real, imag} */,
  {32'hbaf7f600, 32'hbe3300d0} /* (17, 27, 21) {real, imag} */,
  {32'h3c9a4040, 32'hbf0dc0c4} /* (17, 27, 20) {real, imag} */,
  {32'h3d369f20, 32'h3e20aaa0} /* (17, 27, 19) {real, imag} */,
  {32'h3ee3bfb4, 32'h3e78f6e0} /* (17, 27, 18) {real, imag} */,
  {32'h3f52fe1a, 32'h3eea6fe0} /* (17, 27, 17) {real, imag} */,
  {32'h3e6df2f4, 32'h3e0edd00} /* (17, 27, 16) {real, imag} */,
  {32'hbf06652d, 32'hbed48c60} /* (17, 27, 15) {real, imag} */,
  {32'hbebb64f0, 32'h3eeb20e0} /* (17, 27, 14) {real, imag} */,
  {32'hbf2dce68, 32'h3f79dbfc} /* (17, 27, 13) {real, imag} */,
  {32'hbec4dfa0, 32'h3f6cdbe8} /* (17, 27, 12) {real, imag} */,
  {32'h3f000e54, 32'h3f3edb3c} /* (17, 27, 11) {real, imag} */,
  {32'h3f046412, 32'h3eeefb6b} /* (17, 27, 10) {real, imag} */,
  {32'h3d163980, 32'h3e437440} /* (17, 27, 9) {real, imag} */,
  {32'h3b674600, 32'h3ec77c60} /* (17, 27, 8) {real, imag} */,
  {32'h3e989780, 32'h3fa99a14} /* (17, 27, 7) {real, imag} */,
  {32'hbf0e414f, 32'h3f3ca7cc} /* (17, 27, 6) {real, imag} */,
  {32'h3e85cf70, 32'hbf14bcc8} /* (17, 27, 5) {real, imag} */,
  {32'h3f2b8004, 32'hbf441850} /* (17, 27, 4) {real, imag} */,
  {32'h3ec78b26, 32'h3e91d870} /* (17, 27, 3) {real, imag} */,
  {32'hbdea6d00, 32'h3eb39620} /* (17, 27, 2) {real, imag} */,
  {32'h3ea9d206, 32'hbf0e52d4} /* (17, 27, 1) {real, imag} */,
  {32'h3e56e200, 32'hbeced3b0} /* (17, 27, 0) {real, imag} */,
  {32'h3e4247c8, 32'h3de23bf0} /* (17, 26, 31) {real, imag} */,
  {32'h3d0c2950, 32'h3f165360} /* (17, 26, 30) {real, imag} */,
  {32'h3ee37918, 32'h3ec47a60} /* (17, 26, 29) {real, imag} */,
  {32'hbdd2d570, 32'h3f3ee9c8} /* (17, 26, 28) {real, imag} */,
  {32'hbf2aaeef, 32'h3f509b50} /* (17, 26, 27) {real, imag} */,
  {32'hbe63d268, 32'h3eb464e0} /* (17, 26, 26) {real, imag} */,
  {32'hbda5f570, 32'h3e2512e0} /* (17, 26, 25) {real, imag} */,
  {32'hbe8d40a0, 32'h3e1ba600} /* (17, 26, 24) {real, imag} */,
  {32'hbbdc5780, 32'h3e93d978} /* (17, 26, 23) {real, imag} */,
  {32'h3cecbd50, 32'hbddbd3e0} /* (17, 26, 22) {real, imag} */,
  {32'hbcec9b10, 32'h3d519180} /* (17, 26, 21) {real, imag} */,
  {32'hbed4d5e6, 32'h3ec871ac} /* (17, 26, 20) {real, imag} */,
  {32'hbe495f0e, 32'h3ed1ceb0} /* (17, 26, 19) {real, imag} */,
  {32'hbe585dce, 32'h3f3d3570} /* (17, 26, 18) {real, imag} */,
  {32'hbd8e001c, 32'h3f26a22c} /* (17, 26, 17) {real, imag} */,
  {32'h3e272afc, 32'h3c72ea00} /* (17, 26, 16) {real, imag} */,
  {32'h3f103402, 32'hbc739a00} /* (17, 26, 15) {real, imag} */,
  {32'h3f71d048, 32'h3ebb55d8} /* (17, 26, 14) {real, imag} */,
  {32'h3f0a429c, 32'h3ef57eb0} /* (17, 26, 13) {real, imag} */,
  {32'h3d2e3488, 32'h3f2123a0} /* (17, 26, 12) {real, imag} */,
  {32'h3e8912d2, 32'h3f0ff546} /* (17, 26, 11) {real, imag} */,
  {32'h3e97c778, 32'hbe69f5a0} /* (17, 26, 10) {real, imag} */,
  {32'h3c0c7f00, 32'hbe54ad40} /* (17, 26, 9) {real, imag} */,
  {32'hbe253c90, 32'h3e3b1840} /* (17, 26, 8) {real, imag} */,
  {32'h3c10d600, 32'h3eba9030} /* (17, 26, 7) {real, imag} */,
  {32'hbe89955c, 32'h3ec500f0} /* (17, 26, 6) {real, imag} */,
  {32'h3f2f2dfe, 32'h3e0dde20} /* (17, 26, 5) {real, imag} */,
  {32'h3f43f30e, 32'hbe92b360} /* (17, 26, 4) {real, imag} */,
  {32'h3f04cef6, 32'hbcf53900} /* (17, 26, 3) {real, imag} */,
  {32'h3ef03bcd, 32'hbd9440c0} /* (17, 26, 2) {real, imag} */,
  {32'h3ebb7ad2, 32'hbede22b0} /* (17, 26, 1) {real, imag} */,
  {32'h3ea7d35b, 32'h3cb2ed00} /* (17, 26, 0) {real, imag} */,
  {32'h3ed5c26b, 32'h3f277be0} /* (17, 25, 31) {real, imag} */,
  {32'h3c980d20, 32'h3f12c520} /* (17, 25, 30) {real, imag} */,
  {32'h3f230bcf, 32'h3ee436c0} /* (17, 25, 29) {real, imag} */,
  {32'h3eaff3d0, 32'h3f010830} /* (17, 25, 28) {real, imag} */,
  {32'h3e219400, 32'h3f45ebf8} /* (17, 25, 27) {real, imag} */,
  {32'h3e6968d0, 32'h3ee263c0} /* (17, 25, 26) {real, imag} */,
  {32'hbe7ef1e0, 32'h3ecbd1c0} /* (17, 25, 25) {real, imag} */,
  {32'hbdd3b908, 32'h3eef26a0} /* (17, 25, 24) {real, imag} */,
  {32'h3e989a1e, 32'h3f5d2e78} /* (17, 25, 23) {real, imag} */,
  {32'hbeb89c12, 32'h3f1a694c} /* (17, 25, 22) {real, imag} */,
  {32'hbd3e1900, 32'h3f00d292} /* (17, 25, 21) {real, imag} */,
  {32'hbeb80a41, 32'h3f691274} /* (17, 25, 20) {real, imag} */,
  {32'hbe949454, 32'h3f4d5ec0} /* (17, 25, 19) {real, imag} */,
  {32'hbd8fbc88, 32'h3e849690} /* (17, 25, 18) {real, imag} */,
  {32'hbe2ded18, 32'h3f322e78} /* (17, 25, 17) {real, imag} */,
  {32'h3e9a2c34, 32'hbcb78d00} /* (17, 25, 16) {real, imag} */,
  {32'h3f30462e, 32'h3e4ff480} /* (17, 25, 15) {real, imag} */,
  {32'h3f16f9f0, 32'h3d030180} /* (17, 25, 14) {real, imag} */,
  {32'h3e8fd0e0, 32'hbf823964} /* (17, 25, 13) {real, imag} */,
  {32'hbe372cd0, 32'hbea8aab0} /* (17, 25, 12) {real, imag} */,
  {32'h3eb413e2, 32'hbd9f9210} /* (17, 25, 11) {real, imag} */,
  {32'h3e777f80, 32'h3efec400} /* (17, 25, 10) {real, imag} */,
  {32'hbd74e410, 32'h3f110eb0} /* (17, 25, 9) {real, imag} */,
  {32'hbd49e300, 32'h3e0d9f80} /* (17, 25, 8) {real, imag} */,
  {32'hbe3ceb72, 32'hbdb266e0} /* (17, 25, 7) {real, imag} */,
  {32'hbe820de8, 32'h3ecb6988} /* (17, 25, 6) {real, imag} */,
  {32'h3e8d0b02, 32'h3f93ccb0} /* (17, 25, 5) {real, imag} */,
  {32'h3f17477c, 32'h3f49d0c0} /* (17, 25, 4) {real, imag} */,
  {32'h3e3621b0, 32'h3f66339c} /* (17, 25, 3) {real, imag} */,
  {32'hbf0951c0, 32'h3e964a50} /* (17, 25, 2) {real, imag} */,
  {32'hbd902e70, 32'hbd477b80} /* (17, 25, 1) {real, imag} */,
  {32'h3ec56c2c, 32'h3e7df340} /* (17, 25, 0) {real, imag} */,
  {32'h3ea70323, 32'h3f3e0582} /* (17, 24, 31) {real, imag} */,
  {32'h3df6a508, 32'h3f32b4a4} /* (17, 24, 30) {real, imag} */,
  {32'h3e5473d0, 32'hbde58300} /* (17, 24, 29) {real, imag} */,
  {32'h3db318f0, 32'hbf7b1b80} /* (17, 24, 28) {real, imag} */,
  {32'hbddbc938, 32'hbe9f0f98} /* (17, 24, 27) {real, imag} */,
  {32'hbed98478, 32'hbe9d0c38} /* (17, 24, 26) {real, imag} */,
  {32'h3cd95e90, 32'hbd3aae00} /* (17, 24, 25) {real, imag} */,
  {32'h3f4c5659, 32'h3ee90c30} /* (17, 24, 24) {real, imag} */,
  {32'h3e0cb5e0, 32'h3f2c76a8} /* (17, 24, 23) {real, imag} */,
  {32'hbf464928, 32'h3ec39c60} /* (17, 24, 22) {real, imag} */,
  {32'hbe4f88e0, 32'hbd1ce7c0} /* (17, 24, 21) {real, imag} */,
  {32'h3d844438, 32'h3ef12950} /* (17, 24, 20) {real, imag} */,
  {32'h3d3bb7c0, 32'h3f499ba0} /* (17, 24, 19) {real, imag} */,
  {32'h3f557ad0, 32'hbf08b228} /* (17, 24, 18) {real, imag} */,
  {32'h3e8ec385, 32'h3d41bb80} /* (17, 24, 17) {real, imag} */,
  {32'h3e587408, 32'hbe48b540} /* (17, 24, 16) {real, imag} */,
  {32'h3d5cbdb0, 32'hbebaedf8} /* (17, 24, 15) {real, imag} */,
  {32'hbec98bd6, 32'hbf2d42b0} /* (17, 24, 14) {real, imag} */,
  {32'hbe89fdf0, 32'hbfee57f4} /* (17, 24, 13) {real, imag} */,
  {32'hbe0272d4, 32'hbf957d7e} /* (17, 24, 12) {real, imag} */,
  {32'h3e0b6838, 32'h3e602530} /* (17, 24, 11) {real, imag} */,
  {32'h3e21f524, 32'h3f7bb7c4} /* (17, 24, 10) {real, imag} */,
  {32'h3d8f6cc8, 32'h3f820b34} /* (17, 24, 9) {real, imag} */,
  {32'h3e543cb0, 32'hbe6c7a00} /* (17, 24, 8) {real, imag} */,
  {32'hbe602a48, 32'h3e1bc140} /* (17, 24, 7) {real, imag} */,
  {32'hbf30c3d2, 32'h3e98baf8} /* (17, 24, 6) {real, imag} */,
  {32'h3daceb58, 32'h3f34b7e0} /* (17, 24, 5) {real, imag} */,
  {32'h3f04aca7, 32'h3f031ef0} /* (17, 24, 4) {real, imag} */,
  {32'h3f17f46b, 32'h3ecc9640} /* (17, 24, 3) {real, imag} */,
  {32'hbe864dc0, 32'h3da9b540} /* (17, 24, 2) {real, imag} */,
  {32'hbf8633e8, 32'h3ef12610} /* (17, 24, 1) {real, imag} */,
  {32'hbe710bc0, 32'hbd1c9d00} /* (17, 24, 0) {real, imag} */,
  {32'h3e899e02, 32'h3f36c6d4} /* (17, 23, 31) {real, imag} */,
  {32'hbd8533bc, 32'h3f203658} /* (17, 23, 30) {real, imag} */,
  {32'hbecd1fa2, 32'h3c107400} /* (17, 23, 29) {real, imag} */,
  {32'hbda21180, 32'hbe638540} /* (17, 23, 28) {real, imag} */,
  {32'h3db23960, 32'hbe2d2d10} /* (17, 23, 27) {real, imag} */,
  {32'hbe82ed72, 32'hbe4c5780} /* (17, 23, 26) {real, imag} */,
  {32'hbdf101d0, 32'h3e1188d0} /* (17, 23, 25) {real, imag} */,
  {32'h3f173f3c, 32'h3ed636f8} /* (17, 23, 24) {real, imag} */,
  {32'hbf015880, 32'h3efbfb80} /* (17, 23, 23) {real, imag} */,
  {32'hbf78414a, 32'hbe01b640} /* (17, 23, 22) {real, imag} */,
  {32'h3ddddf90, 32'h3d0c9b40} /* (17, 23, 21) {real, imag} */,
  {32'h3e80069e, 32'hbd9be240} /* (17, 23, 20) {real, imag} */,
  {32'h3f0410f1, 32'h3e538680} /* (17, 23, 19) {real, imag} */,
  {32'h3fd75c33, 32'hbf0dfec8} /* (17, 23, 18) {real, imag} */,
  {32'h3f2478e7, 32'hbf60d0d0} /* (17, 23, 17) {real, imag} */,
  {32'hbf0814f2, 32'hbf882768} /* (17, 23, 16) {real, imag} */,
  {32'hbefcf591, 32'hbf54f298} /* (17, 23, 15) {real, imag} */,
  {32'hbdb69af0, 32'hbe09d090} /* (17, 23, 14) {real, imag} */,
  {32'hbeac34d6, 32'hbd423580} /* (17, 23, 13) {real, imag} */,
  {32'hbf2d607a, 32'h3d835d80} /* (17, 23, 12) {real, imag} */,
  {32'hbec8e740, 32'h3e10e980} /* (17, 23, 11) {real, imag} */,
  {32'hbe3f7730, 32'h3eb306c0} /* (17, 23, 10) {real, imag} */,
  {32'hbe83612a, 32'h3e9bc880} /* (17, 23, 9) {real, imag} */,
  {32'h3e603ab0, 32'h3d871e80} /* (17, 23, 8) {real, imag} */,
  {32'h3e250100, 32'hbdf9c180} /* (17, 23, 7) {real, imag} */,
  {32'hbf5be1c2, 32'h3e1f0000} /* (17, 23, 6) {real, imag} */,
  {32'hbe5cb710, 32'h3efb8e80} /* (17, 23, 5) {real, imag} */,
  {32'hbdd3c790, 32'h3eedadc0} /* (17, 23, 4) {real, imag} */,
  {32'h3e8108a4, 32'hbedb9d78} /* (17, 23, 3) {real, imag} */,
  {32'hbb47c000, 32'hbf51faf4} /* (17, 23, 2) {real, imag} */,
  {32'hbf4a8429, 32'h3e1fda90} /* (17, 23, 1) {real, imag} */,
  {32'hbeff275d, 32'h3eb5f548} /* (17, 23, 0) {real, imag} */,
  {32'h3f0e032a, 32'h3ef1cbbc} /* (17, 22, 31) {real, imag} */,
  {32'h3f0a515c, 32'h3f61a978} /* (17, 22, 30) {real, imag} */,
  {32'h3f1f9f60, 32'h3ec3cd70} /* (17, 22, 29) {real, imag} */,
  {32'h3f9b4db9, 32'hbce4fb00} /* (17, 22, 28) {real, imag} */,
  {32'h3f4180ea, 32'hbf1d7440} /* (17, 22, 27) {real, imag} */,
  {32'h3ea09522, 32'hbf555890} /* (17, 22, 26) {real, imag} */,
  {32'h3e08195a, 32'hbe6553e0} /* (17, 22, 25) {real, imag} */,
  {32'h3e56edce, 32'h3e122500} /* (17, 22, 24) {real, imag} */,
  {32'hbf3f2342, 32'h3db35f80} /* (17, 22, 23) {real, imag} */,
  {32'hbf6e4dd6, 32'h3ce5b500} /* (17, 22, 22) {real, imag} */,
  {32'hbea8ddfc, 32'h3e8db420} /* (17, 22, 21) {real, imag} */,
  {32'h3dd55288, 32'hbe562a00} /* (17, 22, 20) {real, imag} */,
  {32'hbda7d694, 32'hbe252e00} /* (17, 22, 19) {real, imag} */,
  {32'h3efa7542, 32'hbe9bdd90} /* (17, 22, 18) {real, imag} */,
  {32'hbe0a372e, 32'hbe289680} /* (17, 22, 17) {real, imag} */,
  {32'hbf7de92d, 32'hbf592440} /* (17, 22, 16) {real, imag} */,
  {32'hbf15b57e, 32'hbf0eb62c} /* (17, 22, 15) {real, imag} */,
  {32'h3e1bcd3e, 32'h3ee63a40} /* (17, 22, 14) {real, imag} */,
  {32'h3ec60a53, 32'h3f5cef78} /* (17, 22, 13) {real, imag} */,
  {32'h3de24e08, 32'h3f6c14b0} /* (17, 22, 12) {real, imag} */,
  {32'hbe200580, 32'h3ee57640} /* (17, 22, 11) {real, imag} */,
  {32'hbf1b6860, 32'h3d979b70} /* (17, 22, 10) {real, imag} */,
  {32'hbe1632a0, 32'hbcce9100} /* (17, 22, 9) {real, imag} */,
  {32'hbde60088, 32'h3f41da98} /* (17, 22, 8) {real, imag} */,
  {32'h3ebb5610, 32'h3ce2d200} /* (17, 22, 7) {real, imag} */,
  {32'h3e601474, 32'hbe98ccf8} /* (17, 22, 6) {real, imag} */,
  {32'h3ca2c980, 32'h3e930ef0} /* (17, 22, 5) {real, imag} */,
  {32'hbe11bcd0, 32'h3f6c00f8} /* (17, 22, 4) {real, imag} */,
  {32'hbe8b82fc, 32'h3e050840} /* (17, 22, 3) {real, imag} */,
  {32'hbf67b6a8, 32'hbf03b4d0} /* (17, 22, 2) {real, imag} */,
  {32'hbf4d96ce, 32'hbe2c83c0} /* (17, 22, 1) {real, imag} */,
  {32'hbf3df622, 32'h3e84c0c0} /* (17, 22, 0) {real, imag} */,
  {32'h3e667c84, 32'h3f05cfaa} /* (17, 21, 31) {real, imag} */,
  {32'h3e99a12c, 32'h3eca1040} /* (17, 21, 30) {real, imag} */,
  {32'h3ee1d994, 32'h3e612ec0} /* (17, 21, 29) {real, imag} */,
  {32'h3f8d0c00, 32'hbd56adc0} /* (17, 21, 28) {real, imag} */,
  {32'h3f4bef1d, 32'hbecd3d80} /* (17, 21, 27) {real, imag} */,
  {32'h3f13c1fc, 32'hbecdff60} /* (17, 21, 26) {real, imag} */,
  {32'h3f39f995, 32'hbf0426e0} /* (17, 21, 25) {real, imag} */,
  {32'h3ef49410, 32'h3a1ed000} /* (17, 21, 24) {real, imag} */,
  {32'hbe81449e, 32'h3d098fc0} /* (17, 21, 23) {real, imag} */,
  {32'hbf3133c6, 32'h3cf27300} /* (17, 21, 22) {real, imag} */,
  {32'hbddcd488, 32'hbc473800} /* (17, 21, 21) {real, imag} */,
  {32'h3eb643c4, 32'hbed7edf4} /* (17, 21, 20) {real, imag} */,
  {32'hbe3466b1, 32'hbd115080} /* (17, 21, 19) {real, imag} */,
  {32'hbd7c3ad0, 32'hbf3c74c0} /* (17, 21, 18) {real, imag} */,
  {32'hbe19d85e, 32'hbee5d860} /* (17, 21, 17) {real, imag} */,
  {32'hbea5215e, 32'h3f044cb5} /* (17, 21, 16) {real, imag} */,
  {32'hbec76588, 32'hbd796600} /* (17, 21, 15) {real, imag} */,
  {32'hbe5e21c4, 32'h3db375c0} /* (17, 21, 14) {real, imag} */,
  {32'h3ea01c3e, 32'h3eeed7d0} /* (17, 21, 13) {real, imag} */,
  {32'h3e2621c9, 32'h3ee52190} /* (17, 21, 12) {real, imag} */,
  {32'hbcbc71e0, 32'hbe008eb0} /* (17, 21, 11) {real, imag} */,
  {32'hbecb15d0, 32'hbeb50d90} /* (17, 21, 10) {real, imag} */,
  {32'h3dc6162c, 32'hbd0be900} /* (17, 21, 9) {real, imag} */,
  {32'hbe9e1f7e, 32'h3e8101a8} /* (17, 21, 8) {real, imag} */,
  {32'hbd286480, 32'h3f0dca70} /* (17, 21, 7) {real, imag} */,
  {32'h3f94b570, 32'hbef1c932} /* (17, 21, 6) {real, imag} */,
  {32'h3f98c73b, 32'h3dee8700} /* (17, 21, 5) {real, imag} */,
  {32'h3f3faebc, 32'h3f05de3c} /* (17, 21, 4) {real, imag} */,
  {32'hbeb42b22, 32'h3e771e10} /* (17, 21, 3) {real, imag} */,
  {32'hbf19fe21, 32'h3eda65d4} /* (17, 21, 2) {real, imag} */,
  {32'hbec323a0, 32'h3f390b86} /* (17, 21, 1) {real, imag} */,
  {32'hbe32d572, 32'h3f452ead} /* (17, 21, 0) {real, imag} */,
  {32'h3deb4780, 32'h3f1f8fe4} /* (17, 20, 31) {real, imag} */,
  {32'h3dcbcc80, 32'h3ee422b0} /* (17, 20, 30) {real, imag} */,
  {32'h3eaad2f4, 32'hbdc3e8e0} /* (17, 20, 29) {real, imag} */,
  {32'h3fb9d3d4, 32'hbe3080d8} /* (17, 20, 28) {real, imag} */,
  {32'h3f36022a, 32'hbe879e80} /* (17, 20, 27) {real, imag} */,
  {32'h3eec670b, 32'hbdadeca0} /* (17, 20, 26) {real, imag} */,
  {32'h3ed61930, 32'hbe7bd888} /* (17, 20, 25) {real, imag} */,
  {32'h3dd51cbc, 32'hbe996e80} /* (17, 20, 24) {real, imag} */,
  {32'hbdfe7e10, 32'h3ea78870} /* (17, 20, 23) {real, imag} */,
  {32'hbeaad1b2, 32'h3efa1530} /* (17, 20, 22) {real, imag} */,
  {32'hbe572950, 32'hbea02f1c} /* (17, 20, 21) {real, imag} */,
  {32'h3e2cb86e, 32'hbf45f600} /* (17, 20, 20) {real, imag} */,
  {32'h3e9a3320, 32'hbf1c3f88} /* (17, 20, 19) {real, imag} */,
  {32'hbd20f2da, 32'hbf84effc} /* (17, 20, 18) {real, imag} */,
  {32'hbe57d9fc, 32'hbf423070} /* (17, 20, 17) {real, imag} */,
  {32'h3f55bb40, 32'h3e6af500} /* (17, 20, 16) {real, imag} */,
  {32'h3eae8970, 32'hbd8a7780} /* (17, 20, 15) {real, imag} */,
  {32'hbf2299ce, 32'hbe99f5b8} /* (17, 20, 14) {real, imag} */,
  {32'hbe00c7b0, 32'hbf0d6648} /* (17, 20, 13) {real, imag} */,
  {32'h3f829efa, 32'h3d12b300} /* (17, 20, 12) {real, imag} */,
  {32'h3f44e65f, 32'h3eb913f0} /* (17, 20, 11) {real, imag} */,
  {32'h3c316f80, 32'h3e449830} /* (17, 20, 10) {real, imag} */,
  {32'h3ebc10a0, 32'h3e067210} /* (17, 20, 9) {real, imag} */,
  {32'h3e02f520, 32'hbece0520} /* (17, 20, 8) {real, imag} */,
  {32'h3dc61494, 32'h3efe83b8} /* (17, 20, 7) {real, imag} */,
  {32'h3f61fc93, 32'hbf2678d0} /* (17, 20, 6) {real, imag} */,
  {32'h3e376a9b, 32'h3dc86cf0} /* (17, 20, 5) {real, imag} */,
  {32'hbe8a824a, 32'h3e65f980} /* (17, 20, 4) {real, imag} */,
  {32'hbdb39310, 32'h3e655e80} /* (17, 20, 3) {real, imag} */,
  {32'hbf0e7799, 32'h3eedd648} /* (17, 20, 2) {real, imag} */,
  {32'hbf0f2a92, 32'h3ea34bb0} /* (17, 20, 1) {real, imag} */,
  {32'h3d302300, 32'h3ecf9848} /* (17, 20, 0) {real, imag} */,
  {32'h3ec24ad3, 32'h3dee9460} /* (17, 19, 31) {real, imag} */,
  {32'h3ee5df54, 32'hbeccfe40} /* (17, 19, 30) {real, imag} */,
  {32'h3e9943ea, 32'hbefc5d30} /* (17, 19, 29) {real, imag} */,
  {32'h3f49f880, 32'hbe5b6340} /* (17, 19, 28) {real, imag} */,
  {32'h3ea3c9a0, 32'hbe3ddf80} /* (17, 19, 27) {real, imag} */,
  {32'h3ec6efb0, 32'h3e3150e0} /* (17, 19, 26) {real, imag} */,
  {32'h3e8dc3e9, 32'h3de52900} /* (17, 19, 25) {real, imag} */,
  {32'hbe031c60, 32'hbe24a900} /* (17, 19, 24) {real, imag} */,
  {32'hbefd43d0, 32'h3e82aac0} /* (17, 19, 23) {real, imag} */,
  {32'hbf4c90fa, 32'h3dcb0380} /* (17, 19, 22) {real, imag} */,
  {32'hbf06332d, 32'hbefc9718} /* (17, 19, 21) {real, imag} */,
  {32'h3e82505a, 32'hbf8e04e0} /* (17, 19, 20) {real, imag} */,
  {32'hbdc0b020, 32'hbf032b20} /* (17, 19, 19) {real, imag} */,
  {32'hbf46f115, 32'hbf40d580} /* (17, 19, 18) {real, imag} */,
  {32'hbe803b4b, 32'hbf449948} /* (17, 19, 17) {real, imag} */,
  {32'h3f6c6916, 32'h3e9c3f10} /* (17, 19, 16) {real, imag} */,
  {32'h3f3618cc, 32'h3e12c340} /* (17, 19, 15) {real, imag} */,
  {32'h3eb0e035, 32'hbeda33f0} /* (17, 19, 14) {real, imag} */,
  {32'h3f0d3a36, 32'hbf866590} /* (17, 19, 13) {real, imag} */,
  {32'h3f5102ce, 32'hbf3be278} /* (17, 19, 12) {real, imag} */,
  {32'h3ee182a4, 32'h3ee8ec20} /* (17, 19, 11) {real, imag} */,
  {32'hbe576e40, 32'h3f0c2cd8} /* (17, 19, 10) {real, imag} */,
  {32'hbe676154, 32'h3ec96940} /* (17, 19, 9) {real, imag} */,
  {32'h3d3aee40, 32'hbe9dbb90} /* (17, 19, 8) {real, imag} */,
  {32'hbe4fade8, 32'hbe33f2b0} /* (17, 19, 7) {real, imag} */,
  {32'hbe0de454, 32'hbf3a8168} /* (17, 19, 6) {real, imag} */,
  {32'hbeb33450, 32'hbe46b910} /* (17, 19, 5) {real, imag} */,
  {32'hbf3029e0, 32'hbea56ca0} /* (17, 19, 4) {real, imag} */,
  {32'hbe234928, 32'hbe8cd918} /* (17, 19, 3) {real, imag} */,
  {32'h3c86f180, 32'h3e15bba0} /* (17, 19, 2) {real, imag} */,
  {32'hbf03dfe8, 32'h3eccfb10} /* (17, 19, 1) {real, imag} */,
  {32'h3ca99ec0, 32'h3c387d00} /* (17, 19, 0) {real, imag} */,
  {32'hbe585688, 32'h3ef6e8c0} /* (17, 18, 31) {real, imag} */,
  {32'hbe98e618, 32'hbe649a40} /* (17, 18, 30) {real, imag} */,
  {32'h3ef02270, 32'hbe6d1f00} /* (17, 18, 29) {real, imag} */,
  {32'h3ead834c, 32'h3eb0bf30} /* (17, 18, 28) {real, imag} */,
  {32'hbeb9e1ca, 32'hbdcfc440} /* (17, 18, 27) {real, imag} */,
  {32'hbef49ce2, 32'h3f0b19c0} /* (17, 18, 26) {real, imag} */,
  {32'h3ea3cc1c, 32'h3e4db800} /* (17, 18, 25) {real, imag} */,
  {32'hb89f0000, 32'h3e364f40} /* (17, 18, 24) {real, imag} */,
  {32'hbf32c25e, 32'hbeed2c40} /* (17, 18, 23) {real, imag} */,
  {32'hbf85fd9e, 32'hbe994290} /* (17, 18, 22) {real, imag} */,
  {32'hbed4d1e4, 32'h3e18e420} /* (17, 18, 21) {real, imag} */,
  {32'h3dd0ba88, 32'hbea88010} /* (17, 18, 20) {real, imag} */,
  {32'hbea4e25c, 32'h3d1c9700} /* (17, 18, 19) {real, imag} */,
  {32'hbf05c5d6, 32'hbf6c4900} /* (17, 18, 18) {real, imag} */,
  {32'h3e84d8a8, 32'hbf203090} /* (17, 18, 17) {real, imag} */,
  {32'h3f02250c, 32'h3c32dc00} /* (17, 18, 16) {real, imag} */,
  {32'h3ecd3dcc, 32'hbe9f7720} /* (17, 18, 15) {real, imag} */,
  {32'h3f60be9c, 32'hbf39a82c} /* (17, 18, 14) {real, imag} */,
  {32'h3f556edc, 32'hbf434010} /* (17, 18, 13) {real, imag} */,
  {32'h3ee6a672, 32'hbf8ae180} /* (17, 18, 12) {real, imag} */,
  {32'h3d018410, 32'h3e931f30} /* (17, 18, 11) {real, imag} */,
  {32'h3e24ca38, 32'h3f58d9a4} /* (17, 18, 10) {real, imag} */,
  {32'hbed6a4d8, 32'h3e434e70} /* (17, 18, 9) {real, imag} */,
  {32'hbf994536, 32'h3ced1a00} /* (17, 18, 8) {real, imag} */,
  {32'hbf8b4c2c, 32'hbea18540} /* (17, 18, 7) {real, imag} */,
  {32'hbd989b68, 32'hbf103ec8} /* (17, 18, 6) {real, imag} */,
  {32'h3e842008, 32'hbf483ce8} /* (17, 18, 5) {real, imag} */,
  {32'h3e434a48, 32'hbf159e34} /* (17, 18, 4) {real, imag} */,
  {32'h3ea81e99, 32'hbc289000} /* (17, 18, 3) {real, imag} */,
  {32'h3f2474bb, 32'hbf18e3d8} /* (17, 18, 2) {real, imag} */,
  {32'h3ecfe668, 32'h3ecb5650} /* (17, 18, 1) {real, imag} */,
  {32'hbe7071c0, 32'h3f2e1b14} /* (17, 18, 0) {real, imag} */,
  {32'hbf991a3b, 32'h3ededa80} /* (17, 17, 31) {real, imag} */,
  {32'hbf56cb8e, 32'h3e19da40} /* (17, 17, 30) {real, imag} */,
  {32'h3d908810, 32'hbe1c3e20} /* (17, 17, 29) {real, imag} */,
  {32'h3e03125c, 32'hbbf0b800} /* (17, 17, 28) {real, imag} */,
  {32'hbe9ea8ec, 32'hbea225a0} /* (17, 17, 27) {real, imag} */,
  {32'hbf5dca6a, 32'h3d7c9780} /* (17, 17, 26) {real, imag} */,
  {32'hbf7b3c03, 32'h3de1edc0} /* (17, 17, 25) {real, imag} */,
  {32'hbf49c924, 32'hbd546180} /* (17, 17, 24) {real, imag} */,
  {32'hbf1ae4f5, 32'hbeab9890} /* (17, 17, 23) {real, imag} */,
  {32'hbf33af62, 32'hbe995cd8} /* (17, 17, 22) {real, imag} */,
  {32'h3e7cffd0, 32'hbdde8428} /* (17, 17, 21) {real, imag} */,
  {32'h3f10e092, 32'h3e00ecf0} /* (17, 17, 20) {real, imag} */,
  {32'h3c3f2980, 32'h3de82580} /* (17, 17, 19) {real, imag} */,
  {32'hbe02638c, 32'hbed710e0} /* (17, 17, 18) {real, imag} */,
  {32'hbee6ea7c, 32'hbe058e40} /* (17, 17, 17) {real, imag} */,
  {32'h3cd65d00, 32'hbee49a30} /* (17, 17, 16) {real, imag} */,
  {32'h3f05b012, 32'hbee96dc0} /* (17, 17, 15) {real, imag} */,
  {32'h3f396aa0, 32'hbe8df5c0} /* (17, 17, 14) {real, imag} */,
  {32'h3ed65e0c, 32'hbf0a80a8} /* (17, 17, 13) {real, imag} */,
  {32'h3f5a99da, 32'hbed3f540} /* (17, 17, 12) {real, imag} */,
  {32'h3f48a3ab, 32'h3f7b5258} /* (17, 17, 11) {real, imag} */,
  {32'h3ee95d7c, 32'h3f9a733c} /* (17, 17, 10) {real, imag} */,
  {32'hbf747fd0, 32'h3f63c568} /* (17, 17, 9) {real, imag} */,
  {32'hbf536bd4, 32'hbd639500} /* (17, 17, 8) {real, imag} */,
  {32'hbe48ecb8, 32'hbe892b50} /* (17, 17, 7) {real, imag} */,
  {32'hbe9b0300, 32'hbe5e3080} /* (17, 17, 6) {real, imag} */,
  {32'h3e87e754, 32'hbf42b364} /* (17, 17, 5) {real, imag} */,
  {32'hbe97dd27, 32'h3c01a400} /* (17, 17, 4) {real, imag} */,
  {32'hbe2c469c, 32'hbef8c3c0} /* (17, 17, 3) {real, imag} */,
  {32'h3f169960, 32'hbf2c4060} /* (17, 17, 2) {real, imag} */,
  {32'h3c40ca80, 32'h3f3d72a0} /* (17, 17, 1) {real, imag} */,
  {32'hbf3b355a, 32'h3f8b29d4} /* (17, 17, 0) {real, imag} */,
  {32'hbf1c4f0a, 32'h3e8c5598} /* (17, 16, 31) {real, imag} */,
  {32'hbf271314, 32'h3e7878e0} /* (17, 16, 30) {real, imag} */,
  {32'hbf0480f0, 32'hbdffaec0} /* (17, 16, 29) {real, imag} */,
  {32'hbec13040, 32'hbf3b2740} /* (17, 16, 28) {real, imag} */,
  {32'hbf0ce2aa, 32'hbeb64670} /* (17, 16, 27) {real, imag} */,
  {32'hbf41b0f7, 32'hbf3989c4} /* (17, 16, 26) {real, imag} */,
  {32'hbf7f9caa, 32'hbf46c52c} /* (17, 16, 25) {real, imag} */,
  {32'hbf358e14, 32'h3df3cb40} /* (17, 16, 24) {real, imag} */,
  {32'h3e29cf66, 32'h3eb7f0c0} /* (17, 16, 23) {real, imag} */,
  {32'hbe800ae8, 32'hbde53d80} /* (17, 16, 22) {real, imag} */,
  {32'h3cf54900, 32'hbec86a01} /* (17, 16, 21) {real, imag} */,
  {32'h3eb4b6c4, 32'hbef96fb0} /* (17, 16, 20) {real, imag} */,
  {32'h3e535278, 32'hbf120b28} /* (17, 16, 19) {real, imag} */,
  {32'h3f150395, 32'hbda37500} /* (17, 16, 18) {real, imag} */,
  {32'h3f3b32be, 32'h3e101aa0} /* (17, 16, 17) {real, imag} */,
  {32'h3f8def93, 32'hbf187c88} /* (17, 16, 16) {real, imag} */,
  {32'h3f1f41c8, 32'hbf110578} /* (17, 16, 15) {real, imag} */,
  {32'hbda93400, 32'hbeddbe40} /* (17, 16, 14) {real, imag} */,
  {32'hbf1d5536, 32'hbf21a3b8} /* (17, 16, 13) {real, imag} */,
  {32'h3f12e45f, 32'h3df41680} /* (17, 16, 12) {real, imag} */,
  {32'h3ef95870, 32'h3f71b198} /* (17, 16, 11) {real, imag} */,
  {32'h3f02d2ae, 32'h3f51d1ea} /* (17, 16, 10) {real, imag} */,
  {32'hbef02bbf, 32'h3f065c28} /* (17, 16, 9) {real, imag} */,
  {32'hbf1cd86e, 32'hbdc683c0} /* (17, 16, 8) {real, imag} */,
  {32'h3aff0800, 32'h3d43ff40} /* (17, 16, 7) {real, imag} */,
  {32'hbd1694a0, 32'hbd43bb00} /* (17, 16, 6) {real, imag} */,
  {32'hbf0c0dd9, 32'hbe347c40} /* (17, 16, 5) {real, imag} */,
  {32'hbf41bf44, 32'h3f1247f0} /* (17, 16, 4) {real, imag} */,
  {32'hbf2033d2, 32'hbe425d40} /* (17, 16, 3) {real, imag} */,
  {32'hbee01220, 32'hbe90b120} /* (17, 16, 2) {real, imag} */,
  {32'hbf5eb25c, 32'h3f9f0a8c} /* (17, 16, 1) {real, imag} */,
  {32'hbf079b7a, 32'h3fa00a64} /* (17, 16, 0) {real, imag} */,
  {32'h3d6abdf0, 32'h3dda6880} /* (17, 15, 31) {real, imag} */,
  {32'hbe6068d0, 32'hbefe72c0} /* (17, 15, 30) {real, imag} */,
  {32'hbf16d3f4, 32'hbf7aa940} /* (17, 15, 29) {real, imag} */,
  {32'hbdeaaab4, 32'hbf6e70f0} /* (17, 15, 28) {real, imag} */,
  {32'hbee05e0b, 32'hbf82b0e4} /* (17, 15, 27) {real, imag} */,
  {32'hbecfbc63, 32'hbf8d9474} /* (17, 15, 26) {real, imag} */,
  {32'hbe9fb010, 32'hbf9844b4} /* (17, 15, 25) {real, imag} */,
  {32'h3e39c98c, 32'h3e619760} /* (17, 15, 24) {real, imag} */,
  {32'h3f40d659, 32'h3d8ee600} /* (17, 15, 23) {real, imag} */,
  {32'hbeb2e665, 32'hbe917f88} /* (17, 15, 22) {real, imag} */,
  {32'hbecff048, 32'hbdf15960} /* (17, 15, 21) {real, imag} */,
  {32'h3bbde500, 32'hbea4ed60} /* (17, 15, 20) {real, imag} */,
  {32'h3f4aba8c, 32'hbf2315a8} /* (17, 15, 19) {real, imag} */,
  {32'h3f806242, 32'h3dd4d180} /* (17, 15, 18) {real, imag} */,
  {32'h3f6b19b8, 32'h3caa2100} /* (17, 15, 17) {real, imag} */,
  {32'h3fabdc7c, 32'hbe2df4a0} /* (17, 15, 16) {real, imag} */,
  {32'h3f29303c, 32'hbe6f6dc0} /* (17, 15, 15) {real, imag} */,
  {32'hbbc47000, 32'hbf39e6cc} /* (17, 15, 14) {real, imag} */,
  {32'h3e5dec06, 32'hbc3a1e00} /* (17, 15, 13) {real, imag} */,
  {32'h3e957c18, 32'h3e4687e0} /* (17, 15, 12) {real, imag} */,
  {32'h3d784aa0, 32'hbe4bc580} /* (17, 15, 11) {real, imag} */,
  {32'h3f19fd44, 32'hbefd94b8} /* (17, 15, 10) {real, imag} */,
  {32'hbebc97ac, 32'hbf1729c0} /* (17, 15, 9) {real, imag} */,
  {32'hbed19120, 32'hbf0248c0} /* (17, 15, 8) {real, imag} */,
  {32'hbe137368, 32'h3f028a70} /* (17, 15, 7) {real, imag} */,
  {32'hbdd2b5c8, 32'h3f31804c} /* (17, 15, 6) {real, imag} */,
  {32'hbf18d484, 32'h3c976900} /* (17, 15, 5) {real, imag} */,
  {32'hbf202358, 32'hbeb89ab0} /* (17, 15, 4) {real, imag} */,
  {32'hbf62f4dc, 32'h3dd520c0} /* (17, 15, 3) {real, imag} */,
  {32'hbf03cccf, 32'h3e5d9b20} /* (17, 15, 2) {real, imag} */,
  {32'hbf455eb1, 32'h3e939e80} /* (17, 15, 1) {real, imag} */,
  {32'hbefb0cb4, 32'h3ec79080} /* (17, 15, 0) {real, imag} */,
  {32'h3ea81773, 32'hbdc52100} /* (17, 14, 31) {real, imag} */,
  {32'h3dac2130, 32'hbf127798} /* (17, 14, 30) {real, imag} */,
  {32'hbd2a2f74, 32'hbfaac034} /* (17, 14, 29) {real, imag} */,
  {32'h3f29dde0, 32'hbf5a72d8} /* (17, 14, 28) {real, imag} */,
  {32'h3e20e598, 32'hbf43c810} /* (17, 14, 27) {real, imag} */,
  {32'hbf7f4484, 32'hbdfdd900} /* (17, 14, 26) {real, imag} */,
  {32'hbf5736f0, 32'hbf29cd38} /* (17, 14, 25) {real, imag} */,
  {32'hbeb1e8c8, 32'hbd781080} /* (17, 14, 24) {real, imag} */,
  {32'hbf109d9a, 32'h3f644c60} /* (17, 14, 23) {real, imag} */,
  {32'hbf1faa0c, 32'h3f93844c} /* (17, 14, 22) {real, imag} */,
  {32'hbeceb720, 32'h3e7a1d10} /* (17, 14, 21) {real, imag} */,
  {32'h3eee9d7c, 32'hbeaac890} /* (17, 14, 20) {real, imag} */,
  {32'h3f834bba, 32'h3dca6440} /* (17, 14, 19) {real, imag} */,
  {32'h3fa039f8, 32'hbe344840} /* (17, 14, 18) {real, imag} */,
  {32'h3ec716d8, 32'hbf2ba2e8} /* (17, 14, 17) {real, imag} */,
  {32'h3ed4e47c, 32'hbd900680} /* (17, 14, 16) {real, imag} */,
  {32'h3efbcbe6, 32'h3eb72df0} /* (17, 14, 15) {real, imag} */,
  {32'h3ee76d80, 32'h3e3eb3a0} /* (17, 14, 14) {real, imag} */,
  {32'h3fb64e10, 32'h3f0d3188} /* (17, 14, 13) {real, imag} */,
  {32'h3f333d81, 32'h3eaf8710} /* (17, 14, 12) {real, imag} */,
  {32'h3d28e550, 32'hbf1d99b4} /* (17, 14, 11) {real, imag} */,
  {32'hbd8a0d90, 32'hbe3c7ce8} /* (17, 14, 10) {real, imag} */,
  {32'hbf1e9f1a, 32'h3e222b60} /* (17, 14, 9) {real, imag} */,
  {32'hbe805318, 32'hbe55d9c0} /* (17, 14, 8) {real, imag} */,
  {32'h3ed410dc, 32'h3e814320} /* (17, 14, 7) {real, imag} */,
  {32'hbd664620, 32'h3f3e1d5c} /* (17, 14, 6) {real, imag} */,
  {32'h3d5d903c, 32'hbdc06460} /* (17, 14, 5) {real, imag} */,
  {32'h3eb69d86, 32'hbf07c7f0} /* (17, 14, 4) {real, imag} */,
  {32'h3e2e2d98, 32'hbdbb7ec0} /* (17, 14, 3) {real, imag} */,
  {32'h3e0616c4, 32'hbe9788c0} /* (17, 14, 2) {real, imag} */,
  {32'h3e10cf78, 32'hbec262e0} /* (17, 14, 1) {real, imag} */,
  {32'hbdd956f0, 32'h3e8ba940} /* (17, 14, 0) {real, imag} */,
  {32'h3ea23b14, 32'hbdee34b0} /* (17, 13, 31) {real, imag} */,
  {32'h3e9e3be9, 32'hbe90c320} /* (17, 13, 30) {real, imag} */,
  {32'hbd16dd30, 32'hbf36aeb0} /* (17, 13, 29) {real, imag} */,
  {32'h3f22d9a0, 32'hbd29fb80} /* (17, 13, 28) {real, imag} */,
  {32'h3d300ce0, 32'h3e8419c0} /* (17, 13, 27) {real, imag} */,
  {32'hbf8df90e, 32'h3d148d40} /* (17, 13, 26) {real, imag} */,
  {32'hbf7d953e, 32'hbed45770} /* (17, 13, 25) {real, imag} */,
  {32'hbf0b7d76, 32'hbd843b00} /* (17, 13, 24) {real, imag} */,
  {32'hbf316f74, 32'h3e9bc350} /* (17, 13, 23) {real, imag} */,
  {32'h3ea4c6ce, 32'h3f01f4e0} /* (17, 13, 22) {real, imag} */,
  {32'h3d1753e0, 32'h3f02067c} /* (17, 13, 21) {real, imag} */,
  {32'h3f38f7e8, 32'h3d82f4c0} /* (17, 13, 20) {real, imag} */,
  {32'h3f3fe360, 32'h3dcc5400} /* (17, 13, 19) {real, imag} */,
  {32'h3e731b90, 32'hbe6ea0f0} /* (17, 13, 18) {real, imag} */,
  {32'h3ed3ecba, 32'hbf2b5844} /* (17, 13, 17) {real, imag} */,
  {32'h3f206e35, 32'hbf0791f8} /* (17, 13, 16) {real, imag} */,
  {32'h3ef8b5c4, 32'h3e81d690} /* (17, 13, 15) {real, imag} */,
  {32'h3e8dc3fe, 32'h3e8aa0d0} /* (17, 13, 14) {real, imag} */,
  {32'h3e519368, 32'hbd7fe000} /* (17, 13, 13) {real, imag} */,
  {32'h3efbc068, 32'hbf1420a8} /* (17, 13, 12) {real, imag} */,
  {32'h3e854772, 32'hbf802a0e} /* (17, 13, 11) {real, imag} */,
  {32'hbea21280, 32'hbe48de90} /* (17, 13, 10) {real, imag} */,
  {32'hbe64b680, 32'h3e22f740} /* (17, 13, 9) {real, imag} */,
  {32'h3ea956c0, 32'h3ec06ff0} /* (17, 13, 8) {real, imag} */,
  {32'h3e5cc0f2, 32'h3f03e2e8} /* (17, 13, 7) {real, imag} */,
  {32'hbe910c44, 32'h3eb818f0} /* (17, 13, 6) {real, imag} */,
  {32'hbebe8238, 32'h3de70b00} /* (17, 13, 5) {real, imag} */,
  {32'hbec9338c, 32'hbc810300} /* (17, 13, 4) {real, imag} */,
  {32'hbf07c446, 32'h3f1b74d0} /* (17, 13, 3) {real, imag} */,
  {32'h3e1495ee, 32'h3ec7aa48} /* (17, 13, 2) {real, imag} */,
  {32'h3e775e08, 32'h3bef4400} /* (17, 13, 1) {real, imag} */,
  {32'hbc362300, 32'hbebe0690} /* (17, 13, 0) {real, imag} */,
  {32'h3e675958, 32'h3cd64900} /* (17, 12, 31) {real, imag} */,
  {32'h3eab34ea, 32'hbed74be0} /* (17, 12, 30) {real, imag} */,
  {32'hbe457900, 32'hbf1fdff8} /* (17, 12, 29) {real, imag} */,
  {32'h3ec60568, 32'h3e91e360} /* (17, 12, 28) {real, imag} */,
  {32'h3d89ee90, 32'h3f7c661c} /* (17, 12, 27) {real, imag} */,
  {32'hbddc28e0, 32'h3ecba3b0} /* (17, 12, 26) {real, imag} */,
  {32'hbd0217a0, 32'hbf08258c} /* (17, 12, 25) {real, imag} */,
  {32'h3dbbda00, 32'hbd000780} /* (17, 12, 24) {real, imag} */,
  {32'hbecf3fdf, 32'h3dab3b80} /* (17, 12, 23) {real, imag} */,
  {32'h3f1cb42e, 32'hbed204c8} /* (17, 12, 22) {real, imag} */,
  {32'h3e4da818, 32'h3ee072bc} /* (17, 12, 21) {real, imag} */,
  {32'h3f5f8a09, 32'h3eb646d0} /* (17, 12, 20) {real, imag} */,
  {32'h3f81dddd, 32'hbeef4690} /* (17, 12, 19) {real, imag} */,
  {32'h3e01553e, 32'hbe5214e0} /* (17, 12, 18) {real, imag} */,
  {32'hbe1abf02, 32'hbe4f79a0} /* (17, 12, 17) {real, imag} */,
  {32'h3ee242a3, 32'hbeb27940} /* (17, 12, 16) {real, imag} */,
  {32'h3e2e3ea0, 32'h3e0c1400} /* (17, 12, 15) {real, imag} */,
  {32'hbea82010, 32'h3e121e20} /* (17, 12, 14) {real, imag} */,
  {32'hbe93a8b0, 32'hbe9c0750} /* (17, 12, 13) {real, imag} */,
  {32'h3eaa60d0, 32'h3de4cb00} /* (17, 12, 12) {real, imag} */,
  {32'h3eb97ec6, 32'hbc6a0300} /* (17, 12, 11) {real, imag} */,
  {32'hbe1efb20, 32'hbeceabd8} /* (17, 12, 10) {real, imag} */,
  {32'h3e1507f0, 32'hbe1919a0} /* (17, 12, 9) {real, imag} */,
  {32'hbdad61a0, 32'h3efd9fe0} /* (17, 12, 8) {real, imag} */,
  {32'hbe88b3b2, 32'h3e7fd240} /* (17, 12, 7) {real, imag} */,
  {32'hbebd40fa, 32'hbd15da00} /* (17, 12, 6) {real, imag} */,
  {32'hbf25653f, 32'h3d165c80} /* (17, 12, 5) {real, imag} */,
  {32'hbf9578d1, 32'hbdb4b9c0} /* (17, 12, 4) {real, imag} */,
  {32'hbfae8320, 32'h3edf3840} /* (17, 12, 3) {real, imag} */,
  {32'hbd855a68, 32'h3ead655c} /* (17, 12, 2) {real, imag} */,
  {32'h3e2f43f0, 32'h3e829be0} /* (17, 12, 1) {real, imag} */,
  {32'hbe78c7ec, 32'hbda3a6e0} /* (17, 12, 0) {real, imag} */,
  {32'hbda04188, 32'hbe55ae38} /* (17, 11, 31) {real, imag} */,
  {32'h3daa43e0, 32'hbf2929dc} /* (17, 11, 30) {real, imag} */,
  {32'h3d2f3804, 32'hbf103480} /* (17, 11, 29) {real, imag} */,
  {32'hbd0a01b8, 32'h3e61e4e0} /* (17, 11, 28) {real, imag} */,
  {32'hbeb688ae, 32'h3f997866} /* (17, 11, 27) {real, imag} */,
  {32'h3da8e038, 32'h3f66d37c} /* (17, 11, 26) {real, imag} */,
  {32'h3ea6f5d8, 32'hbf0fae10} /* (17, 11, 25) {real, imag} */,
  {32'hbebb5364, 32'hbc80f000} /* (17, 11, 24) {real, imag} */,
  {32'hbf937060, 32'h3eee4260} /* (17, 11, 23) {real, imag} */,
  {32'h3ec698f0, 32'h3e5f0b50} /* (17, 11, 22) {real, imag} */,
  {32'h3f6536c2, 32'h3e03ff34} /* (17, 11, 21) {real, imag} */,
  {32'h3fa74998, 32'h3e3dc5f0} /* (17, 11, 20) {real, imag} */,
  {32'h3f6a6377, 32'hbea1ce58} /* (17, 11, 19) {real, imag} */,
  {32'hbe9c78e2, 32'hbf27cc74} /* (17, 11, 18) {real, imag} */,
  {32'hbef76828, 32'hbe50a390} /* (17, 11, 17) {real, imag} */,
  {32'h3e87368c, 32'h3e82dc98} /* (17, 11, 16) {real, imag} */,
  {32'h3e942339, 32'hbc9eb700} /* (17, 11, 15) {real, imag} */,
  {32'hbe88546c, 32'hbd829ac0} /* (17, 11, 14) {real, imag} */,
  {32'hbedd806e, 32'h3d6a9380} /* (17, 11, 13) {real, imag} */,
  {32'h3d50ca40, 32'h3f09bc7c} /* (17, 11, 12) {real, imag} */,
  {32'h3ea565a8, 32'h3ec35078} /* (17, 11, 11) {real, imag} */,
  {32'h3e9a82be, 32'h3e084f90} /* (17, 11, 10) {real, imag} */,
  {32'h3e62356c, 32'h3f6b2f98} /* (17, 11, 9) {real, imag} */,
  {32'hbf8c3f48, 32'h3f864b0c} /* (17, 11, 8) {real, imag} */,
  {32'hbf2c83ba, 32'h3eb830e0} /* (17, 11, 7) {real, imag} */,
  {32'hbf3e6116, 32'hbe4f6f20} /* (17, 11, 6) {real, imag} */,
  {32'hbf1301b6, 32'hbdcb5d40} /* (17, 11, 5) {real, imag} */,
  {32'hbf1c6afa, 32'hbe8a5460} /* (17, 11, 4) {real, imag} */,
  {32'hbf46eb29, 32'hbeade128} /* (17, 11, 3) {real, imag} */,
  {32'hbeb69fa8, 32'h3e8bd120} /* (17, 11, 2) {real, imag} */,
  {32'h3d0c0900, 32'h3f0550a8} /* (17, 11, 1) {real, imag} */,
  {32'hbdb344d0, 32'h3cec3620} /* (17, 11, 0) {real, imag} */,
  {32'hbdc05fc8, 32'h3eb5a520} /* (17, 10, 31) {real, imag} */,
  {32'h3e14a79f, 32'hbe9982c0} /* (17, 10, 30) {real, imag} */,
  {32'hbf36d843, 32'hbe39bc70} /* (17, 10, 29) {real, imag} */,
  {32'hbec2fd26, 32'h3d1eb700} /* (17, 10, 28) {real, imag} */,
  {32'hbe3661d0, 32'h3ec53330} /* (17, 10, 27) {real, imag} */,
  {32'hbe966c06, 32'h3ea2d318} /* (17, 10, 26) {real, imag} */,
  {32'hbd9d5d70, 32'hbdee78b8} /* (17, 10, 25) {real, imag} */,
  {32'hbd0e9540, 32'hbd1d2b6c} /* (17, 10, 24) {real, imag} */,
  {32'hbf33c8a0, 32'h3f417218} /* (17, 10, 23) {real, imag} */,
  {32'h3f22b9fb, 32'h3f6605a8} /* (17, 10, 22) {real, imag} */,
  {32'h3f763166, 32'hbe837680} /* (17, 10, 21) {real, imag} */,
  {32'h3fa9ff1c, 32'h3c894af0} /* (17, 10, 20) {real, imag} */,
  {32'h3ddab6b4, 32'h3f5102a4} /* (17, 10, 19) {real, imag} */,
  {32'hbf2eaaff, 32'hbe7f8b60} /* (17, 10, 18) {real, imag} */,
  {32'hbe5f74c0, 32'hbf405348} /* (17, 10, 17) {real, imag} */,
  {32'hbd66e7c0, 32'hbee97d50} /* (17, 10, 16) {real, imag} */,
  {32'h3f156356, 32'hbf268064} /* (17, 10, 15) {real, imag} */,
  {32'hbcd30b00, 32'hbf24e11c} /* (17, 10, 14) {real, imag} */,
  {32'hbcbf9dc0, 32'h3e020c00} /* (17, 10, 13) {real, imag} */,
  {32'h3e83f33c, 32'hbebf3960} /* (17, 10, 12) {real, imag} */,
  {32'h3c8d2670, 32'h3d962e80} /* (17, 10, 11) {real, imag} */,
  {32'h3e924696, 32'h3f4cf58b} /* (17, 10, 10) {real, imag} */,
  {32'h3f11012c, 32'h3f3b7a96} /* (17, 10, 9) {real, imag} */,
  {32'hbf408bd1, 32'h3e725428} /* (17, 10, 8) {real, imag} */,
  {32'hbe4e3bf0, 32'hbda43ac0} /* (17, 10, 7) {real, imag} */,
  {32'h3dda1d68, 32'hbe1714b8} /* (17, 10, 6) {real, imag} */,
  {32'hbd7c461c, 32'h3d8b1b80} /* (17, 10, 5) {real, imag} */,
  {32'hbe887e88, 32'hbf0308ec} /* (17, 10, 4) {real, imag} */,
  {32'hbf2b2500, 32'hbeefcf50} /* (17, 10, 3) {real, imag} */,
  {32'hbf747efa, 32'h3be9adc0} /* (17, 10, 2) {real, imag} */,
  {32'hbf4b9958, 32'h3f1b3697} /* (17, 10, 1) {real, imag} */,
  {32'hbeb0882e, 32'h3ef6f01a} /* (17, 10, 0) {real, imag} */,
  {32'hbeae9aaa, 32'h3e567df0} /* (17, 9, 31) {real, imag} */,
  {32'h3dde07c0, 32'h3d61fa00} /* (17, 9, 30) {real, imag} */,
  {32'hbf1cfa28, 32'h3e0eeb40} /* (17, 9, 29) {real, imag} */,
  {32'hbec143bf, 32'hbce3d200} /* (17, 9, 28) {real, imag} */,
  {32'h3ef594fe, 32'hbe51fd60} /* (17, 9, 27) {real, imag} */,
  {32'hbe618c12, 32'hbc9ba400} /* (17, 9, 26) {real, imag} */,
  {32'hbe7074f0, 32'h3eeac950} /* (17, 9, 25) {real, imag} */,
  {32'h3ce680e0, 32'h3e2157c0} /* (17, 9, 24) {real, imag} */,
  {32'h3cf5c8c0, 32'h3eb8eaf0} /* (17, 9, 23) {real, imag} */,
  {32'h3d451f20, 32'h3eebb3c8} /* (17, 9, 22) {real, imag} */,
  {32'h3e8b2497, 32'h3c8c9700} /* (17, 9, 21) {real, imag} */,
  {32'h3f3dbb77, 32'hbe8d0990} /* (17, 9, 20) {real, imag} */,
  {32'h3e47123a, 32'h3f8214b2} /* (17, 9, 19) {real, imag} */,
  {32'hbeb5e034, 32'h3e4fa620} /* (17, 9, 18) {real, imag} */,
  {32'hbf31088c, 32'hbf4d1ce0} /* (17, 9, 17) {real, imag} */,
  {32'hbef82088, 32'hbebcf1f0} /* (17, 9, 16) {real, imag} */,
  {32'hbc157d00, 32'hbeb0bbc0} /* (17, 9, 15) {real, imag} */,
  {32'hbf255116, 32'hbe7c3b40} /* (17, 9, 14) {real, imag} */,
  {32'hbdcbb970, 32'h3e3be900} /* (17, 9, 13) {real, imag} */,
  {32'hbe88f52e, 32'hbd159b40} /* (17, 9, 12) {real, imag} */,
  {32'hbf001538, 32'h3f0709b0} /* (17, 9, 11) {real, imag} */,
  {32'h3e49d7b8, 32'h3f5922f7} /* (17, 9, 10) {real, imag} */,
  {32'h3f24e006, 32'h3da96d00} /* (17, 9, 9) {real, imag} */,
  {32'h3e94cff8, 32'hbf14c738} /* (17, 9, 8) {real, imag} */,
  {32'h3e09da90, 32'hbed509f0} /* (17, 9, 7) {real, imag} */,
  {32'h3ebd6b38, 32'hbd4ebe80} /* (17, 9, 6) {real, imag} */,
  {32'h3f3c41ba, 32'h3ee07270} /* (17, 9, 5) {real, imag} */,
  {32'h3e4d3328, 32'hbda4fa80} /* (17, 9, 4) {real, imag} */,
  {32'hbd45c458, 32'hbf0b68d0} /* (17, 9, 3) {real, imag} */,
  {32'h3db01a60, 32'h3e5e5800} /* (17, 9, 2) {real, imag} */,
  {32'h3db95b94, 32'hbd1ad080} /* (17, 9, 1) {real, imag} */,
  {32'h3e08fca8, 32'hbd604c80} /* (17, 9, 0) {real, imag} */,
  {32'hbf21fa4e, 32'h3e2c2248} /* (17, 8, 31) {real, imag} */,
  {32'hbf002872, 32'h3e511560} /* (17, 8, 30) {real, imag} */,
  {32'hbe686f70, 32'hbe052a60} /* (17, 8, 29) {real, imag} */,
  {32'h3d2e5168, 32'h3e5af2e0} /* (17, 8, 28) {real, imag} */,
  {32'h3eadad6e, 32'h3e665e80} /* (17, 8, 27) {real, imag} */,
  {32'h3e8c76b6, 32'hbe816fe0} /* (17, 8, 26) {real, imag} */,
  {32'h3de15f98, 32'hbf17e158} /* (17, 8, 25) {real, imag} */,
  {32'hbf1501ee, 32'hbf3237e0} /* (17, 8, 24) {real, imag} */,
  {32'hbe988bdb, 32'h3dc85a80} /* (17, 8, 23) {real, imag} */,
  {32'hbd21eca0, 32'hbd780800} /* (17, 8, 22) {real, imag} */,
  {32'h3ee3de29, 32'hbf07f618} /* (17, 8, 21) {real, imag} */,
  {32'h3e8caf88, 32'hbe92ba28} /* (17, 8, 20) {real, imag} */,
  {32'hbd8b8760, 32'h3ed4d2f0} /* (17, 8, 19) {real, imag} */,
  {32'hbed804a1, 32'hbeac4be0} /* (17, 8, 18) {real, imag} */,
  {32'hbf7113ce, 32'hbf1f8914} /* (17, 8, 17) {real, imag} */,
  {32'hbe8f8850, 32'hbe603ce0} /* (17, 8, 16) {real, imag} */,
  {32'hbdb70ccc, 32'h3bab0400} /* (17, 8, 15) {real, imag} */,
  {32'hbf518300, 32'h3eae9440} /* (17, 8, 14) {real, imag} */,
  {32'hbedf63d0, 32'h3ac0a000} /* (17, 8, 13) {real, imag} */,
  {32'hbf595d7f, 32'hbf0092e8} /* (17, 8, 12) {real, imag} */,
  {32'hbf291dfe, 32'h3e3cad20} /* (17, 8, 11) {real, imag} */,
  {32'h3ededc6a, 32'h3e3d9680} /* (17, 8, 10) {real, imag} */,
  {32'h3ecc2d54, 32'hbe981d28} /* (17, 8, 9) {real, imag} */,
  {32'h3d34c7f0, 32'hbe8be0b0} /* (17, 8, 8) {real, imag} */,
  {32'h3c41f0a0, 32'hbe5797a0} /* (17, 8, 7) {real, imag} */,
  {32'h3f063b12, 32'hbf1de4b8} /* (17, 8, 6) {real, imag} */,
  {32'h3f2dda32, 32'h3bc6b400} /* (17, 8, 5) {real, imag} */,
  {32'h3eb07b60, 32'h3ca53e80} /* (17, 8, 4) {real, imag} */,
  {32'h3e6a9380, 32'hbe352520} /* (17, 8, 3) {real, imag} */,
  {32'h3f290f06, 32'h3e765010} /* (17, 8, 2) {real, imag} */,
  {32'h3f078fcc, 32'h3d9f07a0} /* (17, 8, 1) {real, imag} */,
  {32'h3f0cdfcc, 32'hbe1b3db0} /* (17, 8, 0) {real, imag} */,
  {32'hbf078332, 32'h3e613b30} /* (17, 7, 31) {real, imag} */,
  {32'hbf4d4740, 32'h3cd1ee00} /* (17, 7, 30) {real, imag} */,
  {32'hbf197733, 32'hbf0bf218} /* (17, 7, 29) {real, imag} */,
  {32'h3ecf600c, 32'hbebacb50} /* (17, 7, 28) {real, imag} */,
  {32'h3dffc3b0, 32'h3dbaf520} /* (17, 7, 27) {real, imag} */,
  {32'h3ee278e4, 32'h3e40de90} /* (17, 7, 26) {real, imag} */,
  {32'h3f83410f, 32'hbee4ac90} /* (17, 7, 25) {real, imag} */,
  {32'h3e1b34c4, 32'hbe12de20} /* (17, 7, 24) {real, imag} */,
  {32'h3e494748, 32'h3f106460} /* (17, 7, 23) {real, imag} */,
  {32'h3f4dae99, 32'h3ea07240} /* (17, 7, 22) {real, imag} */,
  {32'h3f2700a6, 32'hbebfc220} /* (17, 7, 21) {real, imag} */,
  {32'hbeda4328, 32'h3dea3ac0} /* (17, 7, 20) {real, imag} */,
  {32'hbf3c0cdd, 32'h3eef2a88} /* (17, 7, 19) {real, imag} */,
  {32'hbe5b90b2, 32'hbe4617f0} /* (17, 7, 18) {real, imag} */,
  {32'hbf4dd990, 32'hbe4026c0} /* (17, 7, 17) {real, imag} */,
  {32'hbe90b46d, 32'h3d7ca000} /* (17, 7, 16) {real, imag} */,
  {32'h3ec51f42, 32'hbd52cd80} /* (17, 7, 15) {real, imag} */,
  {32'h3f39b4e0, 32'hbe628680} /* (17, 7, 14) {real, imag} */,
  {32'hbd9ddee0, 32'h3c88cb00} /* (17, 7, 13) {real, imag} */,
  {32'hbf76cc60, 32'hbc037e00} /* (17, 7, 12) {real, imag} */,
  {32'hbf403662, 32'hbed084a0} /* (17, 7, 11) {real, imag} */,
  {32'h3eafbc30, 32'hbea78cc8} /* (17, 7, 10) {real, imag} */,
  {32'h3f3b5c73, 32'hbe25d2d0} /* (17, 7, 9) {real, imag} */,
  {32'hbe57d2a0, 32'h3dd6b980} /* (17, 7, 8) {real, imag} */,
  {32'hbe39dc78, 32'h3f144d30} /* (17, 7, 7) {real, imag} */,
  {32'h3e99a9cf, 32'h3da5bd00} /* (17, 7, 6) {real, imag} */,
  {32'h3f6c2d68, 32'hbe890f10} /* (17, 7, 5) {real, imag} */,
  {32'h3f634d3c, 32'h3ea616b8} /* (17, 7, 4) {real, imag} */,
  {32'h3f132cce, 32'hbe85f590} /* (17, 7, 3) {real, imag} */,
  {32'h3f0e8ec4, 32'h3d314300} /* (17, 7, 2) {real, imag} */,
  {32'h3ed2c195, 32'hbe30c680} /* (17, 7, 1) {real, imag} */,
  {32'h3ec4bc4e, 32'hbedd9230} /* (17, 7, 0) {real, imag} */,
  {32'hbe92c41c, 32'h3cc56700} /* (17, 6, 31) {real, imag} */,
  {32'hbe7114a8, 32'hbbbc4800} /* (17, 6, 30) {real, imag} */,
  {32'hbedb33e0, 32'hbe9fb8b8} /* (17, 6, 29) {real, imag} */,
  {32'hbe0d1b48, 32'hbe99f8f8} /* (17, 6, 28) {real, imag} */,
  {32'hbeaa5f9c, 32'hbe54f840} /* (17, 6, 27) {real, imag} */,
  {32'h3e3b0194, 32'hbcadd380} /* (17, 6, 26) {real, imag} */,
  {32'h3edb4cdc, 32'h3e116310} /* (17, 6, 25) {real, imag} */,
  {32'h3cd4d600, 32'h3e60cfc0} /* (17, 6, 24) {real, imag} */,
  {32'h3f616014, 32'h3da5f600} /* (17, 6, 23) {real, imag} */,
  {32'h3f6db643, 32'h3de92980} /* (17, 6, 22) {real, imag} */,
  {32'h3f1a67cd, 32'h3d1c0d00} /* (17, 6, 21) {real, imag} */,
  {32'hbec32297, 32'h3bf0f000} /* (17, 6, 20) {real, imag} */,
  {32'hbf3970e0, 32'h3e5aef30} /* (17, 6, 19) {real, imag} */,
  {32'hbd7926e0, 32'hbf15e9d8} /* (17, 6, 18) {real, imag} */,
  {32'hbe21708e, 32'hbf85b914} /* (17, 6, 17) {real, imag} */,
  {32'hbe531308, 32'hbebbac30} /* (17, 6, 16) {real, imag} */,
  {32'hbdb65e80, 32'h3e1f3200} /* (17, 6, 15) {real, imag} */,
  {32'h3f638a82, 32'hbdfbfa40} /* (17, 6, 14) {real, imag} */,
  {32'h3ebacd94, 32'hbea34500} /* (17, 6, 13) {real, imag} */,
  {32'hbf136527, 32'hbe46c900} /* (17, 6, 12) {real, imag} */,
  {32'hbefa2cda, 32'hbf4682b4} /* (17, 6, 11) {real, imag} */,
  {32'h3dbf75c0, 32'hbf2b4490} /* (17, 6, 10) {real, imag} */,
  {32'h3ebfba08, 32'hbe199240} /* (17, 6, 9) {real, imag} */,
  {32'hbeb3f465, 32'h3ef49290} /* (17, 6, 8) {real, imag} */,
  {32'hbf0fd1be, 32'hbe3c9e00} /* (17, 6, 7) {real, imag} */,
  {32'hbecb3dd9, 32'hbe2b75e0} /* (17, 6, 6) {real, imag} */,
  {32'h3df2ad10, 32'h3ea39160} /* (17, 6, 5) {real, imag} */,
  {32'h3eb9b730, 32'h3ed08948} /* (17, 6, 4) {real, imag} */,
  {32'h3e9811d8, 32'hbec35b60} /* (17, 6, 3) {real, imag} */,
  {32'h3e400cc8, 32'hbf087f20} /* (17, 6, 2) {real, imag} */,
  {32'hbe83a684, 32'hbedb3cb0} /* (17, 6, 1) {real, imag} */,
  {32'h3de58ba4, 32'hbed09cc8} /* (17, 6, 0) {real, imag} */,
  {32'hbec3f13a, 32'hbdb4cd40} /* (17, 5, 31) {real, imag} */,
  {32'h3dab7360, 32'hbdd69780} /* (17, 5, 30) {real, imag} */,
  {32'hbe430898, 32'hbe0652c0} /* (17, 5, 29) {real, imag} */,
  {32'hbefe5356, 32'hbebeea10} /* (17, 5, 28) {real, imag} */,
  {32'hbf1c754e, 32'hbb8c8000} /* (17, 5, 27) {real, imag} */,
  {32'h3ea51ad2, 32'hbe3ecdb0} /* (17, 5, 26) {real, imag} */,
  {32'hbea3d233, 32'hbef261b0} /* (17, 5, 25) {real, imag} */,
  {32'hbe8f0a8a, 32'h3eb52f30} /* (17, 5, 24) {real, imag} */,
  {32'h3f1a24b0, 32'h3e7341e0} /* (17, 5, 23) {real, imag} */,
  {32'h3eaf3fe4, 32'hbe44b860} /* (17, 5, 22) {real, imag} */,
  {32'hbeaee19c, 32'hbc154900} /* (17, 5, 21) {real, imag} */,
  {32'hbe9b04ae, 32'hbf02ebc4} /* (17, 5, 20) {real, imag} */,
  {32'h3d11eb40, 32'hbed0c8d4} /* (17, 5, 19) {real, imag} */,
  {32'h3d527770, 32'hbf277ece} /* (17, 5, 18) {real, imag} */,
  {32'hbd91cf80, 32'hbf67bce5} /* (17, 5, 17) {real, imag} */,
  {32'hbf1841ce, 32'hbe2fec28} /* (17, 5, 16) {real, imag} */,
  {32'hbe8fc720, 32'h3e9835b0} /* (17, 5, 15) {real, imag} */,
  {32'h3e97866e, 32'hbd9e9e80} /* (17, 5, 14) {real, imag} */,
  {32'h3da26ee0, 32'hbedc80d8} /* (17, 5, 13) {real, imag} */,
  {32'hbee2f898, 32'hbedf30e0} /* (17, 5, 12) {real, imag} */,
  {32'hbeec33f4, 32'hbed3c5f0} /* (17, 5, 11) {real, imag} */,
  {32'hbf025a67, 32'hbe3dd220} /* (17, 5, 10) {real, imag} */,
  {32'h3ead1318, 32'hbec57048} /* (17, 5, 9) {real, imag} */,
  {32'hbdfef7e8, 32'hbe016868} /* (17, 5, 8) {real, imag} */,
  {32'hbf8a8997, 32'hbf9089e7} /* (17, 5, 7) {real, imag} */,
  {32'hbf4bec45, 32'hbee89dc8} /* (17, 5, 6) {real, imag} */,
  {32'hbead5788, 32'h3f9eb0c6} /* (17, 5, 5) {real, imag} */,
  {32'hbd902330, 32'h3f53cb80} /* (17, 5, 4) {real, imag} */,
  {32'h3f5253c0, 32'h3d3c9100} /* (17, 5, 3) {real, imag} */,
  {32'h3ecc1f2c, 32'hbbe23800} /* (17, 5, 2) {real, imag} */,
  {32'hbd49c380, 32'h3f2fdd70} /* (17, 5, 1) {real, imag} */,
  {32'hbdab8e14, 32'h3e2a4230} /* (17, 5, 0) {real, imag} */,
  {32'hbefea862, 32'h3ddab440} /* (17, 4, 31) {real, imag} */,
  {32'hbeb02d6e, 32'h3f22b8f0} /* (17, 4, 30) {real, imag} */,
  {32'h3e5a3194, 32'h3eaf7de8} /* (17, 4, 29) {real, imag} */,
  {32'hbebf4913, 32'hbf0897b0} /* (17, 4, 28) {real, imag} */,
  {32'hbf26efe4, 32'hbea2fe80} /* (17, 4, 27) {real, imag} */,
  {32'hbe12f858, 32'h3d650000} /* (17, 4, 26) {real, imag} */,
  {32'hbe41d588, 32'h3ebfe0b0} /* (17, 4, 25) {real, imag} */,
  {32'hbde0dd40, 32'h3f757d88} /* (17, 4, 24) {real, imag} */,
  {32'h3e09fc78, 32'h3f70a8b0} /* (17, 4, 23) {real, imag} */,
  {32'h3ee5e7aa, 32'h3bfb1000} /* (17, 4, 22) {real, imag} */,
  {32'hbea02210, 32'h3d330f00} /* (17, 4, 21) {real, imag} */,
  {32'hbe707d10, 32'hbe751440} /* (17, 4, 20) {real, imag} */,
  {32'h3e8c24d8, 32'h3d973e00} /* (17, 4, 19) {real, imag} */,
  {32'hbdf12bb8, 32'hbde95840} /* (17, 4, 18) {real, imag} */,
  {32'hbeca8e52, 32'hbcfb1000} /* (17, 4, 17) {real, imag} */,
  {32'hbe6ff924, 32'h3f77335c} /* (17, 4, 16) {real, imag} */,
  {32'h3e9109f8, 32'h3f217d20} /* (17, 4, 15) {real, imag} */,
  {32'h3f1da52c, 32'hbe03c870} /* (17, 4, 14) {real, imag} */,
  {32'h3dc357e0, 32'hbeb7e3d0} /* (17, 4, 13) {real, imag} */,
  {32'hbf514cd2, 32'h3dfca320} /* (17, 4, 12) {real, imag} */,
  {32'hbf070472, 32'hbe6a6440} /* (17, 4, 11) {real, imag} */,
  {32'hbea9adb8, 32'h3dde3c00} /* (17, 4, 10) {real, imag} */,
  {32'hbf2ea7aa, 32'h3ed37770} /* (17, 4, 9) {real, imag} */,
  {32'hbf6e4056, 32'h3e41d1e0} /* (17, 4, 8) {real, imag} */,
  {32'hbf6ed3f1, 32'hbf144818} /* (17, 4, 7) {real, imag} */,
  {32'hbf3a0cc6, 32'hbf666fe8} /* (17, 4, 6) {real, imag} */,
  {32'hbe1a2b10, 32'h3d163ca8} /* (17, 4, 5) {real, imag} */,
  {32'h3e3044c0, 32'h3ed72d60} /* (17, 4, 4) {real, imag} */,
  {32'h3f91eab2, 32'h3ec62560} /* (17, 4, 3) {real, imag} */,
  {32'h3ebdaa41, 32'h3e706790} /* (17, 4, 2) {real, imag} */,
  {32'hbe499a22, 32'hbdabf440} /* (17, 4, 1) {real, imag} */,
  {32'hbe3d2076, 32'h3e1f44b0} /* (17, 4, 0) {real, imag} */,
  {32'hbe996cf4, 32'h3ed34ca0} /* (17, 3, 31) {real, imag} */,
  {32'hbeb3d50e, 32'h3f7ec5cc} /* (17, 3, 30) {real, imag} */,
  {32'h3f135038, 32'h3e4b1460} /* (17, 3, 29) {real, imag} */,
  {32'h3f207d8c, 32'hbde3ce80} /* (17, 3, 28) {real, imag} */,
  {32'h3ec88999, 32'h3e993430} /* (17, 3, 27) {real, imag} */,
  {32'h3f2cdef1, 32'h3f507940} /* (17, 3, 26) {real, imag} */,
  {32'h3ece0492, 32'h3c4a1000} /* (17, 3, 25) {real, imag} */,
  {32'h3e825f24, 32'hbebbc630} /* (17, 3, 24) {real, imag} */,
  {32'h3dfceab8, 32'hbe9c8ea0} /* (17, 3, 23) {real, imag} */,
  {32'h3f19b2c2, 32'hbe38f200} /* (17, 3, 22) {real, imag} */,
  {32'h3f0c8a3e, 32'hbef41300} /* (17, 3, 21) {real, imag} */,
  {32'hbe082ae4, 32'hbe56d700} /* (17, 3, 20) {real, imag} */,
  {32'hbf3a7fae, 32'h3da83200} /* (17, 3, 19) {real, imag} */,
  {32'hbf87eff9, 32'h3e804c88} /* (17, 3, 18) {real, imag} */,
  {32'hbf2c9002, 32'h3e784600} /* (17, 3, 17) {real, imag} */,
  {32'h3e0f34a8, 32'h3f504c32} /* (17, 3, 16) {real, imag} */,
  {32'h3e0a64aa, 32'hbc226a00} /* (17, 3, 15) {real, imag} */,
  {32'h3e96bbf8, 32'hbe9ffb60} /* (17, 3, 14) {real, imag} */,
  {32'h3d7242a0, 32'hbeb3f590} /* (17, 3, 13) {real, imag} */,
  {32'hbf748516, 32'h3ed155d0} /* (17, 3, 12) {real, imag} */,
  {32'hbe501fc0, 32'hbefda320} /* (17, 3, 11) {real, imag} */,
  {32'hbecb4caa, 32'hbe098420} /* (17, 3, 10) {real, imag} */,
  {32'hbf8a942e, 32'h3e9164c0} /* (17, 3, 9) {real, imag} */,
  {32'hbd848cd0, 32'hbe5f6a00} /* (17, 3, 8) {real, imag} */,
  {32'h3e84d114, 32'hbf980c2c} /* (17, 3, 7) {real, imag} */,
  {32'hbd3a36c0, 32'hbfba10e4} /* (17, 3, 6) {real, imag} */,
  {32'h3f3f6109, 32'hbf7c438d} /* (17, 3, 5) {real, imag} */,
  {32'h3f1d3255, 32'h3de731c0} /* (17, 3, 4) {real, imag} */,
  {32'h3f2b52ec, 32'h3f768b2c} /* (17, 3, 3) {real, imag} */,
  {32'h3f261002, 32'h3f6c1924} /* (17, 3, 2) {real, imag} */,
  {32'h3e9cdee4, 32'h3e486b40} /* (17, 3, 1) {real, imag} */,
  {32'h3e56e522, 32'h3ed0bfc8} /* (17, 3, 0) {real, imag} */,
  {32'hbed9029f, 32'h3acb1c00} /* (17, 2, 31) {real, imag} */,
  {32'h3dff1320, 32'h3e4650c0} /* (17, 2, 30) {real, imag} */,
  {32'h3f7f2676, 32'h3eb9a1a0} /* (17, 2, 29) {real, imag} */,
  {32'h3fd3f55c, 32'h3e992140} /* (17, 2, 28) {real, imag} */,
  {32'h3f5ff9b6, 32'h3e9f0360} /* (17, 2, 27) {real, imag} */,
  {32'h3f11678e, 32'h3f674ffc} /* (17, 2, 26) {real, imag} */,
  {32'h3f021986, 32'hbe9da510} /* (17, 2, 25) {real, imag} */,
  {32'h3f8515c3, 32'hbe8e3750} /* (17, 2, 24) {real, imag} */,
  {32'h3ed7e2b2, 32'hbf2cfb10} /* (17, 2, 23) {real, imag} */,
  {32'h3e566fb0, 32'hbed58d10} /* (17, 2, 22) {real, imag} */,
  {32'h3ec262dc, 32'h3e63b050} /* (17, 2, 21) {real, imag} */,
  {32'hbe1de84a, 32'h3eae61b0} /* (17, 2, 20) {real, imag} */,
  {32'hbf16e58f, 32'hbebcad40} /* (17, 2, 19) {real, imag} */,
  {32'hbfc95664, 32'hbe0f3080} /* (17, 2, 18) {real, imag} */,
  {32'hbf324cac, 32'hbd627880} /* (17, 2, 17) {real, imag} */,
  {32'h3e4b4f2c, 32'h3e4f7ff0} /* (17, 2, 16) {real, imag} */,
  {32'hbe83067e, 32'hbe3a6d68} /* (17, 2, 15) {real, imag} */,
  {32'hbed038aa, 32'hbd6565c0} /* (17, 2, 14) {real, imag} */,
  {32'hbeab02c7, 32'h3d98e880} /* (17, 2, 13) {real, imag} */,
  {32'hbe8cd4fe, 32'h3f238598} /* (17, 2, 12) {real, imag} */,
  {32'h3dc6b028, 32'h3e55d240} /* (17, 2, 11) {real, imag} */,
  {32'hbf57da5f, 32'h3df04400} /* (17, 2, 10) {real, imag} */,
  {32'hbf544b19, 32'hbea0c820} /* (17, 2, 9) {real, imag} */,
  {32'h3e851186, 32'hbdb23e80} /* (17, 2, 8) {real, imag} */,
  {32'h3e4e6e5c, 32'hbf73fd38} /* (17, 2, 7) {real, imag} */,
  {32'h3c5898c0, 32'hbfdb2ff4} /* (17, 2, 6) {real, imag} */,
  {32'h3f7e5e44, 32'hbf5ca278} /* (17, 2, 5) {real, imag} */,
  {32'h3ee98f20, 32'h3efc3870} /* (17, 2, 4) {real, imag} */,
  {32'hbe777c3c, 32'h3f287e90} /* (17, 2, 3) {real, imag} */,
  {32'h3f13cc12, 32'h3e96df20} /* (17, 2, 2) {real, imag} */,
  {32'h3ebc62c7, 32'hbed88988} /* (17, 2, 1) {real, imag} */,
  {32'h3e3dcce4, 32'hbe9130dc} /* (17, 2, 0) {real, imag} */,
  {32'hbf1ad656, 32'hbec91510} /* (17, 1, 31) {real, imag} */,
  {32'hbe586a2e, 32'hbd4cf940} /* (17, 1, 30) {real, imag} */,
  {32'h3ca06840, 32'h3f0e8620} /* (17, 1, 29) {real, imag} */,
  {32'h3e9ba038, 32'h3f29ff50} /* (17, 1, 28) {real, imag} */,
  {32'hbe17262e, 32'h3e173ac0} /* (17, 1, 27) {real, imag} */,
  {32'hbe5fb1c0, 32'hbeba8f58} /* (17, 1, 26) {real, imag} */,
  {32'hbe5d4e18, 32'hbf6a1cf4} /* (17, 1, 25) {real, imag} */,
  {32'h3cc0fdc0, 32'h3d693100} /* (17, 1, 24) {real, imag} */,
  {32'hbdd9dac0, 32'h3ed21de8} /* (17, 1, 23) {real, imag} */,
  {32'h3daab8c0, 32'hbe2e5b88} /* (17, 1, 22) {real, imag} */,
  {32'h3e0c4708, 32'h3e3f8100} /* (17, 1, 21) {real, imag} */,
  {32'hbe3853d7, 32'h3f0ccac8} /* (17, 1, 20) {real, imag} */,
  {32'hbe205fd4, 32'hbe886a00} /* (17, 1, 19) {real, imag} */,
  {32'hbf6968b0, 32'hbf177358} /* (17, 1, 18) {real, imag} */,
  {32'hbdf77a60, 32'h3ef97a60} /* (17, 1, 17) {real, imag} */,
  {32'hbe1c8142, 32'h3f663810} /* (17, 1, 16) {real, imag} */,
  {32'hbe54216a, 32'hbb3c6200} /* (17, 1, 15) {real, imag} */,
  {32'h3eecb161, 32'h3ec51640} /* (17, 1, 14) {real, imag} */,
  {32'h3d80a4f0, 32'h3f0e5c48} /* (17, 1, 13) {real, imag} */,
  {32'hbe167ecc, 32'h3f259750} /* (17, 1, 12) {real, imag} */,
  {32'hbea34ec4, 32'h3ef80570} /* (17, 1, 11) {real, imag} */,
  {32'hbf05ed52, 32'hbf0b5838} /* (17, 1, 10) {real, imag} */,
  {32'hbe08ff58, 32'hbee41390} /* (17, 1, 9) {real, imag} */,
  {32'h3ede188c, 32'h3e9b7170} /* (17, 1, 8) {real, imag} */,
  {32'h3cc791c0, 32'hbdd50ec0} /* (17, 1, 7) {real, imag} */,
  {32'hbe33cdb8, 32'hbf7ea39c} /* (17, 1, 6) {real, imag} */,
  {32'hbe18d9d4, 32'hbeed5e6c} /* (17, 1, 5) {real, imag} */,
  {32'hbe146774, 32'h3f0cb2f0} /* (17, 1, 4) {real, imag} */,
  {32'hbea8ecf4, 32'h3da8f7c0} /* (17, 1, 3) {real, imag} */,
  {32'h3ea4082e, 32'hbf1aac0c} /* (17, 1, 2) {real, imag} */,
  {32'h3e75e692, 32'hbf4e6264} /* (17, 1, 1) {real, imag} */,
  {32'hbb927d00, 32'hbf2c22bb} /* (17, 1, 0) {real, imag} */,
  {32'hbe8e0127, 32'h3e180230} /* (17, 0, 31) {real, imag} */,
  {32'hbed1d47d, 32'hbdf08ca0} /* (17, 0, 30) {real, imag} */,
  {32'hbf1f8cc0, 32'hbec8d9e8} /* (17, 0, 29) {real, imag} */,
  {32'hbe60fa38, 32'hbde139a0} /* (17, 0, 28) {real, imag} */,
  {32'hbe919bc5, 32'hbed1f6d0} /* (17, 0, 27) {real, imag} */,
  {32'hbd83cc74, 32'hbee79af0} /* (17, 0, 26) {real, imag} */,
  {32'h3bb6ca00, 32'hbf0c4590} /* (17, 0, 25) {real, imag} */,
  {32'hbe90c1e3, 32'h3e2dfca8} /* (17, 0, 24) {real, imag} */,
  {32'hbea8f684, 32'h3f1ee9b2} /* (17, 0, 23) {real, imag} */,
  {32'h3e13a2f8, 32'hbd77d9b8} /* (17, 0, 22) {real, imag} */,
  {32'h3e85ddc4, 32'h3da8e480} /* (17, 0, 21) {real, imag} */,
  {32'hbdce49b0, 32'h3f190886} /* (17, 0, 20) {real, imag} */,
  {32'hbd1941a8, 32'h3e917060} /* (17, 0, 19) {real, imag} */,
  {32'hbe18637c, 32'hbe87fea8} /* (17, 0, 18) {real, imag} */,
  {32'h3e656fd0, 32'h3ee33840} /* (17, 0, 17) {real, imag} */,
  {32'hbe396768, 32'h3e9093e8} /* (17, 0, 16) {real, imag} */,
  {32'hbe6ad578, 32'hbe91ff10} /* (17, 0, 15) {real, imag} */,
  {32'h3e627c98, 32'h3e7a1500} /* (17, 0, 14) {real, imag} */,
  {32'h3e741fbc, 32'hbe1e9f60} /* (17, 0, 13) {real, imag} */,
  {32'hbe32b268, 32'hbe3b3f70} /* (17, 0, 12) {real, imag} */,
  {32'hbf30a782, 32'hbe048940} /* (17, 0, 11) {real, imag} */,
  {32'hbeb93976, 32'hbf1ffedc} /* (17, 0, 10) {real, imag} */,
  {32'hbdf56baf, 32'hbed53a38} /* (17, 0, 9) {real, imag} */,
  {32'h3e49b1c1, 32'h3e1d30b0} /* (17, 0, 8) {real, imag} */,
  {32'hbe75bcf8, 32'hbdb353b0} /* (17, 0, 7) {real, imag} */,
  {32'h3e1bb980, 32'hbf00f06c} /* (17, 0, 6) {real, imag} */,
  {32'hbe053c44, 32'hbe9d1d7a} /* (17, 0, 5) {real, imag} */,
  {32'hbec2740a, 32'hbd5dd430} /* (17, 0, 4) {real, imag} */,
  {32'h3c866da0, 32'hbe9b68b0} /* (17, 0, 3) {real, imag} */,
  {32'h3ed856e4, 32'hbe9fea38} /* (17, 0, 2) {real, imag} */,
  {32'h3f2a4788, 32'hbded3820} /* (17, 0, 1) {real, imag} */,
  {32'h3f047024, 32'hbe72aac0} /* (17, 0, 0) {real, imag} */,
  {32'h3e1bef3c, 32'h00000000} /* (16, 31, 31) {real, imag} */,
  {32'hbf28c52b, 32'h00000000} /* (16, 31, 30) {real, imag} */,
  {32'hbf9be408, 32'h00000000} /* (16, 31, 29) {real, imag} */,
  {32'hbeb9a5a2, 32'h00000000} /* (16, 31, 28) {real, imag} */,
  {32'hbcc0bb20, 32'h00000000} /* (16, 31, 27) {real, imag} */,
  {32'h3e853d8a, 32'h00000000} /* (16, 31, 26) {real, imag} */,
  {32'h3e129550, 32'h00000000} /* (16, 31, 25) {real, imag} */,
  {32'hbcedcfc0, 32'h00000000} /* (16, 31, 24) {real, imag} */,
  {32'hbee1817e, 32'h00000000} /* (16, 31, 23) {real, imag} */,
  {32'h3e9817a8, 32'h00000000} /* (16, 31, 22) {real, imag} */,
  {32'h3f13c640, 32'h00000000} /* (16, 31, 21) {real, imag} */,
  {32'h3e600108, 32'h00000000} /* (16, 31, 20) {real, imag} */,
  {32'hbc8a8100, 32'h00000000} /* (16, 31, 19) {real, imag} */,
  {32'hbeb05524, 32'h00000000} /* (16, 31, 18) {real, imag} */,
  {32'hbdcfb160, 32'h00000000} /* (16, 31, 17) {real, imag} */,
  {32'hbed368f8, 32'h00000000} /* (16, 31, 16) {real, imag} */,
  {32'hbeeba0d7, 32'h00000000} /* (16, 31, 15) {real, imag} */,
  {32'hbc885fe0, 32'h00000000} /* (16, 31, 14) {real, imag} */,
  {32'h3f51e654, 32'h00000000} /* (16, 31, 13) {real, imag} */,
  {32'h3f935368, 32'h00000000} /* (16, 31, 12) {real, imag} */,
  {32'h3cad2d60, 32'h00000000} /* (16, 31, 11) {real, imag} */,
  {32'hbf27ae91, 32'h00000000} /* (16, 31, 10) {real, imag} */,
  {32'hbf18448a, 32'h00000000} /* (16, 31, 9) {real, imag} */,
  {32'hbf92f876, 32'h00000000} /* (16, 31, 8) {real, imag} */,
  {32'hbf56415e, 32'h00000000} /* (16, 31, 7) {real, imag} */,
  {32'hbf6b08e5, 32'h00000000} /* (16, 31, 6) {real, imag} */,
  {32'hbf9f20de, 32'h00000000} /* (16, 31, 5) {real, imag} */,
  {32'hbe5ef024, 32'h00000000} /* (16, 31, 4) {real, imag} */,
  {32'h3eaec902, 32'h00000000} /* (16, 31, 3) {real, imag} */,
  {32'h3e85edfe, 32'h00000000} /* (16, 31, 2) {real, imag} */,
  {32'h3f33e594, 32'h00000000} /* (16, 31, 1) {real, imag} */,
  {32'h3eb80524, 32'h00000000} /* (16, 31, 0) {real, imag} */,
  {32'h3e4af7a6, 32'h00000000} /* (16, 30, 31) {real, imag} */,
  {32'h3e66d78c, 32'h00000000} /* (16, 30, 30) {real, imag} */,
  {32'hbf7bdb5a, 32'h00000000} /* (16, 30, 29) {real, imag} */,
  {32'hbf2cc240, 32'h00000000} /* (16, 30, 28) {real, imag} */,
  {32'hbe2664d8, 32'h00000000} /* (16, 30, 27) {real, imag} */,
  {32'h3f5e986f, 32'h00000000} /* (16, 30, 26) {real, imag} */,
  {32'hbe952518, 32'h00000000} /* (16, 30, 25) {real, imag} */,
  {32'hbe438410, 32'h00000000} /* (16, 30, 24) {real, imag} */,
  {32'hbdc49580, 32'h00000000} /* (16, 30, 23) {real, imag} */,
  {32'h3e8acd6e, 32'h00000000} /* (16, 30, 22) {real, imag} */,
  {32'h3f403620, 32'h00000000} /* (16, 30, 21) {real, imag} */,
  {32'h3f36fbbb, 32'h00000000} /* (16, 30, 20) {real, imag} */,
  {32'h3e34ac5c, 32'h00000000} /* (16, 30, 19) {real, imag} */,
  {32'hbf01aa76, 32'h00000000} /* (16, 30, 18) {real, imag} */,
  {32'hbc93d440, 32'h00000000} /* (16, 30, 17) {real, imag} */,
  {32'hbdb87f88, 32'h00000000} /* (16, 30, 16) {real, imag} */,
  {32'h3e243e74, 32'h00000000} /* (16, 30, 15) {real, imag} */,
  {32'h3f0cc2c8, 32'h00000000} /* (16, 30, 14) {real, imag} */,
  {32'h3f5b625e, 32'h00000000} /* (16, 30, 13) {real, imag} */,
  {32'h3f38c3e8, 32'h00000000} /* (16, 30, 12) {real, imag} */,
  {32'hbeb669fa, 32'h00000000} /* (16, 30, 11) {real, imag} */,
  {32'hbe0782d0, 32'h00000000} /* (16, 30, 10) {real, imag} */,
  {32'hbe16ed5c, 32'h00000000} /* (16, 30, 9) {real, imag} */,
  {32'hbf87fc27, 32'h00000000} /* (16, 30, 8) {real, imag} */,
  {32'hbf547d46, 32'h00000000} /* (16, 30, 7) {real, imag} */,
  {32'hbf15459a, 32'h00000000} /* (16, 30, 6) {real, imag} */,
  {32'hbf730056, 32'h00000000} /* (16, 30, 5) {real, imag} */,
  {32'hbeef7978, 32'h00000000} /* (16, 30, 4) {real, imag} */,
  {32'hbd671990, 32'h00000000} /* (16, 30, 3) {real, imag} */,
  {32'hbe6b6a88, 32'h00000000} /* (16, 30, 2) {real, imag} */,
  {32'h3f4cfca0, 32'h00000000} /* (16, 30, 1) {real, imag} */,
  {32'h3e3ea5d0, 32'h00000000} /* (16, 30, 0) {real, imag} */,
  {32'h3f0839f0, 32'h00000000} /* (16, 29, 31) {real, imag} */,
  {32'h3f812b2c, 32'h00000000} /* (16, 29, 30) {real, imag} */,
  {32'hbea342a8, 32'h00000000} /* (16, 29, 29) {real, imag} */,
  {32'h3de56030, 32'h00000000} /* (16, 29, 28) {real, imag} */,
  {32'h3f34d742, 32'h00000000} /* (16, 29, 27) {real, imag} */,
  {32'h3ee2d1e8, 32'h00000000} /* (16, 29, 26) {real, imag} */,
  {32'hbee3e2b8, 32'h00000000} /* (16, 29, 25) {real, imag} */,
  {32'hbf40bbf4, 32'h00000000} /* (16, 29, 24) {real, imag} */,
  {32'hbda1a4d8, 32'h00000000} /* (16, 29, 23) {real, imag} */,
  {32'hbe2a7eec, 32'h00000000} /* (16, 29, 22) {real, imag} */,
  {32'hbdeeaf80, 32'h00000000} /* (16, 29, 21) {real, imag} */,
  {32'hbd482550, 32'h00000000} /* (16, 29, 20) {real, imag} */,
  {32'hbf0355a6, 32'h00000000} /* (16, 29, 19) {real, imag} */,
  {32'hbf90fd68, 32'h00000000} /* (16, 29, 18) {real, imag} */,
  {32'hbd7e4d00, 32'h00000000} /* (16, 29, 17) {real, imag} */,
  {32'h3f1a5e76, 32'h00000000} /* (16, 29, 16) {real, imag} */,
  {32'h3fc1483e, 32'h00000000} /* (16, 29, 15) {real, imag} */,
  {32'h3fa73b5e, 32'h00000000} /* (16, 29, 14) {real, imag} */,
  {32'h3edbcff0, 32'h00000000} /* (16, 29, 13) {real, imag} */,
  {32'hbece5088, 32'h00000000} /* (16, 29, 12) {real, imag} */,
  {32'hbed265c4, 32'h00000000} /* (16, 29, 11) {real, imag} */,
  {32'h3edcf6d4, 32'h00000000} /* (16, 29, 10) {real, imag} */,
  {32'h3e918bf0, 32'h00000000} /* (16, 29, 9) {real, imag} */,
  {32'hbe7d8ebc, 32'h00000000} /* (16, 29, 8) {real, imag} */,
  {32'hbda81320, 32'h00000000} /* (16, 29, 7) {real, imag} */,
  {32'h3ea7d038, 32'h00000000} /* (16, 29, 6) {real, imag} */,
  {32'h3f00eab4, 32'h00000000} /* (16, 29, 5) {real, imag} */,
  {32'h3ea8c530, 32'h00000000} /* (16, 29, 4) {real, imag} */,
  {32'hbeb50f6c, 32'h00000000} /* (16, 29, 3) {real, imag} */,
  {32'hbf36b544, 32'h00000000} /* (16, 29, 2) {real, imag} */,
  {32'hbcf385e0, 32'h00000000} /* (16, 29, 1) {real, imag} */,
  {32'hbe16e6b8, 32'h00000000} /* (16, 29, 0) {real, imag} */,
  {32'h3d134548, 32'h00000000} /* (16, 28, 31) {real, imag} */,
  {32'h3fa2d38e, 32'h00000000} /* (16, 28, 30) {real, imag} */,
  {32'h3f55b250, 32'h00000000} /* (16, 28, 29) {real, imag} */,
  {32'h3f3a2608, 32'h00000000} /* (16, 28, 28) {real, imag} */,
  {32'h3fb60483, 32'h00000000} /* (16, 28, 27) {real, imag} */,
  {32'h3e457be8, 32'h00000000} /* (16, 28, 26) {real, imag} */,
  {32'hbe5cab10, 32'h00000000} /* (16, 28, 25) {real, imag} */,
  {32'hbe03e860, 32'h00000000} /* (16, 28, 24) {real, imag} */,
  {32'hbda8f590, 32'h00000000} /* (16, 28, 23) {real, imag} */,
  {32'hbebd9974, 32'h00000000} /* (16, 28, 22) {real, imag} */,
  {32'h3d27f070, 32'h00000000} /* (16, 28, 21) {real, imag} */,
  {32'hbebfd9ec, 32'h00000000} /* (16, 28, 20) {real, imag} */,
  {32'hbf888393, 32'h00000000} /* (16, 28, 19) {real, imag} */,
  {32'hbf96b52a, 32'h00000000} /* (16, 28, 18) {real, imag} */,
  {32'hbf54e708, 32'h00000000} /* (16, 28, 17) {real, imag} */,
  {32'hbea297c8, 32'h00000000} /* (16, 28, 16) {real, imag} */,
  {32'h3f2cf968, 32'h00000000} /* (16, 28, 15) {real, imag} */,
  {32'hbed75da8, 32'h00000000} /* (16, 28, 14) {real, imag} */,
  {32'hbf27f690, 32'h00000000} /* (16, 28, 13) {real, imag} */,
  {32'hbf4739fc, 32'h00000000} /* (16, 28, 12) {real, imag} */,
  {32'hbe35b300, 32'h00000000} /* (16, 28, 11) {real, imag} */,
  {32'hbe88efd8, 32'h00000000} /* (16, 28, 10) {real, imag} */,
  {32'hbf2ce98c, 32'h00000000} /* (16, 28, 9) {real, imag} */,
  {32'hbeef5dd8, 32'h00000000} /* (16, 28, 8) {real, imag} */,
  {32'h3e8bed94, 32'h00000000} /* (16, 28, 7) {real, imag} */,
  {32'h3f980b79, 32'h00000000} /* (16, 28, 6) {real, imag} */,
  {32'h3f0d4938, 32'h00000000} /* (16, 28, 5) {real, imag} */,
  {32'h3f9000d8, 32'h00000000} /* (16, 28, 4) {real, imag} */,
  {32'h3f0b8828, 32'h00000000} /* (16, 28, 3) {real, imag} */,
  {32'h3f38c59b, 32'h00000000} /* (16, 28, 2) {real, imag} */,
  {32'h3eef7a4c, 32'h00000000} /* (16, 28, 1) {real, imag} */,
  {32'hbc57fe00, 32'h00000000} /* (16, 28, 0) {real, imag} */,
  {32'h3f1bea98, 32'h00000000} /* (16, 27, 31) {real, imag} */,
  {32'h3fe9c1b3, 32'h00000000} /* (16, 27, 30) {real, imag} */,
  {32'h400d1f82, 32'h00000000} /* (16, 27, 29) {real, imag} */,
  {32'h3f82148b, 32'h00000000} /* (16, 27, 28) {real, imag} */,
  {32'h3f7984c3, 32'h00000000} /* (16, 27, 27) {real, imag} */,
  {32'hbf4a306e, 32'h00000000} /* (16, 27, 26) {real, imag} */,
  {32'hbf90e3c0, 32'h00000000} /* (16, 27, 25) {real, imag} */,
  {32'h3f3e2c7e, 32'h00000000} /* (16, 27, 24) {real, imag} */,
  {32'h3fc5bb54, 32'h00000000} /* (16, 27, 23) {real, imag} */,
  {32'h3f946afb, 32'h00000000} /* (16, 27, 22) {real, imag} */,
  {32'h3f486fe4, 32'h00000000} /* (16, 27, 21) {real, imag} */,
  {32'h3f04433e, 32'h00000000} /* (16, 27, 20) {real, imag} */,
  {32'hbf4e6877, 32'h00000000} /* (16, 27, 19) {real, imag} */,
  {32'hbf98e86b, 32'h00000000} /* (16, 27, 18) {real, imag} */,
  {32'hbf59fb1d, 32'h00000000} /* (16, 27, 17) {real, imag} */,
  {32'hbe019a90, 32'h00000000} /* (16, 27, 16) {real, imag} */,
  {32'h3e6dacc8, 32'h00000000} /* (16, 27, 15) {real, imag} */,
  {32'hbf75af7c, 32'h00000000} /* (16, 27, 14) {real, imag} */,
  {32'hbf278646, 32'h00000000} /* (16, 27, 13) {real, imag} */,
  {32'h3e857348, 32'h00000000} /* (16, 27, 12) {real, imag} */,
  {32'hba25c000, 32'h00000000} /* (16, 27, 11) {real, imag} */,
  {32'hbe4c1de8, 32'h00000000} /* (16, 27, 10) {real, imag} */,
  {32'hbd820990, 32'h00000000} /* (16, 27, 9) {real, imag} */,
  {32'h3e870130, 32'h00000000} /* (16, 27, 8) {real, imag} */,
  {32'h3e569528, 32'h00000000} /* (16, 27, 7) {real, imag} */,
  {32'h3ec85a18, 32'h00000000} /* (16, 27, 6) {real, imag} */,
  {32'h3ed916bc, 32'h00000000} /* (16, 27, 5) {real, imag} */,
  {32'h3f6d030b, 32'h00000000} /* (16, 27, 4) {real, imag} */,
  {32'h3f0c8380, 32'h00000000} /* (16, 27, 3) {real, imag} */,
  {32'h3fb00296, 32'h00000000} /* (16, 27, 2) {real, imag} */,
  {32'h3f370644, 32'h00000000} /* (16, 27, 1) {real, imag} */,
  {32'h3ec290ba, 32'h00000000} /* (16, 27, 0) {real, imag} */,
  {32'h3e45a7b4, 32'h00000000} /* (16, 26, 31) {real, imag} */,
  {32'h3e34cc48, 32'h00000000} /* (16, 26, 30) {real, imag} */,
  {32'h3eaa42dc, 32'h00000000} /* (16, 26, 29) {real, imag} */,
  {32'hbde26f78, 32'h00000000} /* (16, 26, 28) {real, imag} */,
  {32'h3e98cad4, 32'h00000000} /* (16, 26, 27) {real, imag} */,
  {32'hbf7dc6e4, 32'h00000000} /* (16, 26, 26) {real, imag} */,
  {32'hbf2faf2c, 32'h00000000} /* (16, 26, 25) {real, imag} */,
  {32'h3e0b6f70, 32'h00000000} /* (16, 26, 24) {real, imag} */,
  {32'hbe210940, 32'h00000000} /* (16, 26, 23) {real, imag} */,
  {32'h3d99f2f0, 32'h00000000} /* (16, 26, 22) {real, imag} */,
  {32'hbeca57a8, 32'h00000000} /* (16, 26, 21) {real, imag} */,
  {32'h3e225140, 32'h00000000} /* (16, 26, 20) {real, imag} */,
  {32'hbe88ed90, 32'h00000000} /* (16, 26, 19) {real, imag} */,
  {32'hbf174e82, 32'h00000000} /* (16, 26, 18) {real, imag} */,
  {32'hbe9f9278, 32'h00000000} /* (16, 26, 17) {real, imag} */,
  {32'h3f07e2d8, 32'h00000000} /* (16, 26, 16) {real, imag} */,
  {32'h3eabc5a8, 32'h00000000} /* (16, 26, 15) {real, imag} */,
  {32'hbedb663c, 32'h00000000} /* (16, 26, 14) {real, imag} */,
  {32'hbebbfb22, 32'h00000000} /* (16, 26, 13) {real, imag} */,
  {32'h3f4a6ff5, 32'h00000000} /* (16, 26, 12) {real, imag} */,
  {32'hbd6a12e0, 32'h00000000} /* (16, 26, 11) {real, imag} */,
  {32'h3e802888, 32'h00000000} /* (16, 26, 10) {real, imag} */,
  {32'h3f9b9f8f, 32'h00000000} /* (16, 26, 9) {real, imag} */,
  {32'h3fcf7286, 32'h00000000} /* (16, 26, 8) {real, imag} */,
  {32'h3f07c5cc, 32'h00000000} /* (16, 26, 7) {real, imag} */,
  {32'hbe897d1e, 32'h00000000} /* (16, 26, 6) {real, imag} */,
  {32'h3e2a94f8, 32'h00000000} /* (16, 26, 5) {real, imag} */,
  {32'h3dbec5f0, 32'h00000000} /* (16, 26, 4) {real, imag} */,
  {32'hbed7e28c, 32'h00000000} /* (16, 26, 3) {real, imag} */,
  {32'h3ef58b28, 32'h00000000} /* (16, 26, 2) {real, imag} */,
  {32'h3e634eb8, 32'h00000000} /* (16, 26, 1) {real, imag} */,
  {32'h3e900b48, 32'h00000000} /* (16, 26, 0) {real, imag} */,
  {32'h3ec394fd, 32'h00000000} /* (16, 25, 31) {real, imag} */,
  {32'h3ecc9910, 32'h00000000} /* (16, 25, 30) {real, imag} */,
  {32'hbef5d536, 32'h00000000} /* (16, 25, 29) {real, imag} */,
  {32'hbcd6e000, 32'h00000000} /* (16, 25, 28) {real, imag} */,
  {32'h3eef62b8, 32'h00000000} /* (16, 25, 27) {real, imag} */,
  {32'hbed0f3b4, 32'h00000000} /* (16, 25, 26) {real, imag} */,
  {32'hbeaa798c, 32'h00000000} /* (16, 25, 25) {real, imag} */,
  {32'hbe875122, 32'h00000000} /* (16, 25, 24) {real, imag} */,
  {32'hbf4cd690, 32'h00000000} /* (16, 25, 23) {real, imag} */,
  {32'h3e4c0930, 32'h00000000} /* (16, 25, 22) {real, imag} */,
  {32'hbd7229c0, 32'h00000000} /* (16, 25, 21) {real, imag} */,
  {32'hbdd63e60, 32'h00000000} /* (16, 25, 20) {real, imag} */,
  {32'h3d8b6100, 32'h00000000} /* (16, 25, 19) {real, imag} */,
  {32'hbe9e6afe, 32'h00000000} /* (16, 25, 18) {real, imag} */,
  {32'hbf2f4990, 32'h00000000} /* (16, 25, 17) {real, imag} */,
  {32'hbe385ac0, 32'h00000000} /* (16, 25, 16) {real, imag} */,
  {32'hbf45e168, 32'h00000000} /* (16, 25, 15) {real, imag} */,
  {32'hbf7571c8, 32'h00000000} /* (16, 25, 14) {real, imag} */,
  {32'hbe915100, 32'h00000000} /* (16, 25, 13) {real, imag} */,
  {32'h3e26e410, 32'h00000000} /* (16, 25, 12) {real, imag} */,
  {32'h3f340fe2, 32'h00000000} /* (16, 25, 11) {real, imag} */,
  {32'h3f7af34e, 32'h00000000} /* (16, 25, 10) {real, imag} */,
  {32'h3e6d3300, 32'h00000000} /* (16, 25, 9) {real, imag} */,
  {32'hbf6c1c24, 32'h00000000} /* (16, 25, 8) {real, imag} */,
  {32'hbf46908f, 32'h00000000} /* (16, 25, 7) {real, imag} */,
  {32'hbf940aa4, 32'h00000000} /* (16, 25, 6) {real, imag} */,
  {32'hbf7c7d70, 32'h00000000} /* (16, 25, 5) {real, imag} */,
  {32'hbf2d49ca, 32'h00000000} /* (16, 25, 4) {real, imag} */,
  {32'hbef2cb06, 32'h00000000} /* (16, 25, 3) {real, imag} */,
  {32'h3f1d3bf4, 32'h00000000} /* (16, 25, 2) {real, imag} */,
  {32'h3f118084, 32'h00000000} /* (16, 25, 1) {real, imag} */,
  {32'h3d5911c0, 32'h00000000} /* (16, 25, 0) {real, imag} */,
  {32'h3ecaa584, 32'h00000000} /* (16, 24, 31) {real, imag} */,
  {32'hbd013020, 32'h00000000} /* (16, 24, 30) {real, imag} */,
  {32'h3ef59528, 32'h00000000} /* (16, 24, 29) {real, imag} */,
  {32'h3fae72c6, 32'h00000000} /* (16, 24, 28) {real, imag} */,
  {32'h3f788a16, 32'h00000000} /* (16, 24, 27) {real, imag} */,
  {32'hbdd9fea8, 32'h00000000} /* (16, 24, 26) {real, imag} */,
  {32'hbf232f23, 32'h00000000} /* (16, 24, 25) {real, imag} */,
  {32'hbf82e9f7, 32'h00000000} /* (16, 24, 24) {real, imag} */,
  {32'hbf1ffaa4, 32'h00000000} /* (16, 24, 23) {real, imag} */,
  {32'h3ec21a04, 32'h00000000} /* (16, 24, 22) {real, imag} */,
  {32'hbf0a664c, 32'h00000000} /* (16, 24, 21) {real, imag} */,
  {32'hbf51ac8e, 32'h00000000} /* (16, 24, 20) {real, imag} */,
  {32'hbe82a784, 32'h00000000} /* (16, 24, 19) {real, imag} */,
  {32'h3e19a6d0, 32'h00000000} /* (16, 24, 18) {real, imag} */,
  {32'hbd076100, 32'h00000000} /* (16, 24, 17) {real, imag} */,
  {32'h3eb78a48, 32'h00000000} /* (16, 24, 16) {real, imag} */,
  {32'hbe9567d6, 32'h00000000} /* (16, 24, 15) {real, imag} */,
  {32'hbfa5f6c4, 32'h00000000} /* (16, 24, 14) {real, imag} */,
  {32'h3e507358, 32'h00000000} /* (16, 24, 13) {real, imag} */,
  {32'hbea4a390, 32'h00000000} /* (16, 24, 12) {real, imag} */,
  {32'hbe7d88d0, 32'h00000000} /* (16, 24, 11) {real, imag} */,
  {32'hbdd82ae0, 32'h00000000} /* (16, 24, 10) {real, imag} */,
  {32'hbebcb718, 32'h00000000} /* (16, 24, 9) {real, imag} */,
  {32'hbf5a2e66, 32'h00000000} /* (16, 24, 8) {real, imag} */,
  {32'hbec70b10, 32'h00000000} /* (16, 24, 7) {real, imag} */,
  {32'hbf8559c0, 32'h00000000} /* (16, 24, 6) {real, imag} */,
  {32'hbf19529e, 32'h00000000} /* (16, 24, 5) {real, imag} */,
  {32'hbea99960, 32'h00000000} /* (16, 24, 4) {real, imag} */,
  {32'hbe256e28, 32'h00000000} /* (16, 24, 3) {real, imag} */,
  {32'h3f0d2294, 32'h00000000} /* (16, 24, 2) {real, imag} */,
  {32'h3ef7b5d0, 32'h00000000} /* (16, 24, 1) {real, imag} */,
  {32'h3eae7968, 32'h00000000} /* (16, 24, 0) {real, imag} */,
  {32'h3f07c984, 32'h00000000} /* (16, 23, 31) {real, imag} */,
  {32'h3ed6b6a0, 32'h00000000} /* (16, 23, 30) {real, imag} */,
  {32'h3ef91810, 32'h00000000} /* (16, 23, 29) {real, imag} */,
  {32'h3f122074, 32'h00000000} /* (16, 23, 28) {real, imag} */,
  {32'h3dd409e0, 32'h00000000} /* (16, 23, 27) {real, imag} */,
  {32'h3e60ccb0, 32'h00000000} /* (16, 23, 26) {real, imag} */,
  {32'h3ee31f8c, 32'h00000000} /* (16, 23, 25) {real, imag} */,
  {32'hbf78d28d, 32'h00000000} /* (16, 23, 24) {real, imag} */,
  {32'hbf768f5a, 32'h00000000} /* (16, 23, 23) {real, imag} */,
  {32'h3e8da8cc, 32'h00000000} /* (16, 23, 22) {real, imag} */,
  {32'hbe6d20b8, 32'h00000000} /* (16, 23, 21) {real, imag} */,
  {32'hbe7bced8, 32'h00000000} /* (16, 23, 20) {real, imag} */,
  {32'h3e0f84d0, 32'h00000000} /* (16, 23, 19) {real, imag} */,
  {32'hbe1e7f1c, 32'h00000000} /* (16, 23, 18) {real, imag} */,
  {32'h3e262350, 32'h00000000} /* (16, 23, 17) {real, imag} */,
  {32'h3ec2a5e4, 32'h00000000} /* (16, 23, 16) {real, imag} */,
  {32'h3ea60fac, 32'h00000000} /* (16, 23, 15) {real, imag} */,
  {32'hbecf6874, 32'h00000000} /* (16, 23, 14) {real, imag} */,
  {32'hbd61f500, 32'h00000000} /* (16, 23, 13) {real, imag} */,
  {32'hbe422544, 32'h00000000} /* (16, 23, 12) {real, imag} */,
  {32'hbf0655da, 32'h00000000} /* (16, 23, 11) {real, imag} */,
  {32'hbf17268c, 32'h00000000} /* (16, 23, 10) {real, imag} */,
  {32'hbf2cc82c, 32'h00000000} /* (16, 23, 9) {real, imag} */,
  {32'hbf949d10, 32'h00000000} /* (16, 23, 8) {real, imag} */,
  {32'hbf558508, 32'h00000000} /* (16, 23, 7) {real, imag} */,
  {32'hbf172683, 32'h00000000} /* (16, 23, 6) {real, imag} */,
  {32'h3d540900, 32'h00000000} /* (16, 23, 5) {real, imag} */,
  {32'h3e924c30, 32'h00000000} /* (16, 23, 4) {real, imag} */,
  {32'h3f11a3d3, 32'h00000000} /* (16, 23, 3) {real, imag} */,
  {32'h3da98a90, 32'h00000000} /* (16, 23, 2) {real, imag} */,
  {32'hbf51977c, 32'h00000000} /* (16, 23, 1) {real, imag} */,
  {32'h3d26ea20, 32'h00000000} /* (16, 23, 0) {real, imag} */,
  {32'h3e77916c, 32'h00000000} /* (16, 22, 31) {real, imag} */,
  {32'h3f3a5246, 32'h00000000} /* (16, 22, 30) {real, imag} */,
  {32'hbf14cdbb, 32'h00000000} /* (16, 22, 29) {real, imag} */,
  {32'hbf94fb85, 32'h00000000} /* (16, 22, 28) {real, imag} */,
  {32'hbf05c172, 32'h00000000} /* (16, 22, 27) {real, imag} */,
  {32'h3edc8030, 32'h00000000} /* (16, 22, 26) {real, imag} */,
  {32'h3e61f46c, 32'h00000000} /* (16, 22, 25) {real, imag} */,
  {32'hbf911b5a, 32'h00000000} /* (16, 22, 24) {real, imag} */,
  {32'hbf400520, 32'h00000000} /* (16, 22, 23) {real, imag} */,
  {32'h3e97cbd0, 32'h00000000} /* (16, 22, 22) {real, imag} */,
  {32'hbd279550, 32'h00000000} /* (16, 22, 21) {real, imag} */,
  {32'h3e9a8414, 32'h00000000} /* (16, 22, 20) {real, imag} */,
  {32'h3f4e8ee8, 32'h00000000} /* (16, 22, 19) {real, imag} */,
  {32'h3d5ebb20, 32'h00000000} /* (16, 22, 18) {real, imag} */,
  {32'h3ee806d6, 32'h00000000} /* (16, 22, 17) {real, imag} */,
  {32'h3f662ea9, 32'h00000000} /* (16, 22, 16) {real, imag} */,
  {32'h3ec328c8, 32'h00000000} /* (16, 22, 15) {real, imag} */,
  {32'h3e4abd8c, 32'h00000000} /* (16, 22, 14) {real, imag} */,
  {32'h3f0ff81e, 32'h00000000} /* (16, 22, 13) {real, imag} */,
  {32'h3f79ff32, 32'h00000000} /* (16, 22, 12) {real, imag} */,
  {32'h3e00a398, 32'h00000000} /* (16, 22, 11) {real, imag} */,
  {32'h3e23b1ac, 32'h00000000} /* (16, 22, 10) {real, imag} */,
  {32'hbecafbd0, 32'h00000000} /* (16, 22, 9) {real, imag} */,
  {32'hbedb1adc, 32'h00000000} /* (16, 22, 8) {real, imag} */,
  {32'hbefe6714, 32'h00000000} /* (16, 22, 7) {real, imag} */,
  {32'hbec96be8, 32'h00000000} /* (16, 22, 6) {real, imag} */,
  {32'h3ee0e9d0, 32'h00000000} /* (16, 22, 5) {real, imag} */,
  {32'h3f2345a5, 32'h00000000} /* (16, 22, 4) {real, imag} */,
  {32'h3f5448fe, 32'h00000000} /* (16, 22, 3) {real, imag} */,
  {32'h3e9d6eb0, 32'h00000000} /* (16, 22, 2) {real, imag} */,
  {32'hbf3b9bbc, 32'h00000000} /* (16, 22, 1) {real, imag} */,
  {32'hbf01073a, 32'h00000000} /* (16, 22, 0) {real, imag} */,
  {32'hbdfe69e0, 32'h00000000} /* (16, 21, 31) {real, imag} */,
  {32'hbea729d5, 32'h00000000} /* (16, 21, 30) {real, imag} */,
  {32'hbfb4750c, 32'h00000000} /* (16, 21, 29) {real, imag} */,
  {32'hbfb3728c, 32'h00000000} /* (16, 21, 28) {real, imag} */,
  {32'hbf345a82, 32'h00000000} /* (16, 21, 27) {real, imag} */,
  {32'hbf0135ec, 32'h00000000} /* (16, 21, 26) {real, imag} */,
  {32'hbdc73000, 32'h00000000} /* (16, 21, 25) {real, imag} */,
  {32'hbf5783da, 32'h00000000} /* (16, 21, 24) {real, imag} */,
  {32'hbd294510, 32'h00000000} /* (16, 21, 23) {real, imag} */,
  {32'h3e8fc4f0, 32'h00000000} /* (16, 21, 22) {real, imag} */,
  {32'hbf17ff84, 32'h00000000} /* (16, 21, 21) {real, imag} */,
  {32'hbe826a14, 32'h00000000} /* (16, 21, 20) {real, imag} */,
  {32'h3f1e0dd1, 32'h00000000} /* (16, 21, 19) {real, imag} */,
  {32'h3f168f0c, 32'h00000000} /* (16, 21, 18) {real, imag} */,
  {32'h3f4c7bdf, 32'h00000000} /* (16, 21, 17) {real, imag} */,
  {32'h3f7fb553, 32'h00000000} /* (16, 21, 16) {real, imag} */,
  {32'h3e98e389, 32'h00000000} /* (16, 21, 15) {real, imag} */,
  {32'hbe32e610, 32'h00000000} /* (16, 21, 14) {real, imag} */,
  {32'h3f019510, 32'h00000000} /* (16, 21, 13) {real, imag} */,
  {32'h3eac78e8, 32'h00000000} /* (16, 21, 12) {real, imag} */,
  {32'hbde9df40, 32'h00000000} /* (16, 21, 11) {real, imag} */,
  {32'h3e21d8dc, 32'h00000000} /* (16, 21, 10) {real, imag} */,
  {32'h3f253e90, 32'h00000000} /* (16, 21, 9) {real, imag} */,
  {32'h3f561901, 32'h00000000} /* (16, 21, 8) {real, imag} */,
  {32'hbf33135a, 32'h00000000} /* (16, 21, 7) {real, imag} */,
  {32'h3bba5e00, 32'h00000000} /* (16, 21, 6) {real, imag} */,
  {32'h3dc22188, 32'h00000000} /* (16, 21, 5) {real, imag} */,
  {32'hbe75dce0, 32'h00000000} /* (16, 21, 4) {real, imag} */,
  {32'hbd9dfcf8, 32'h00000000} /* (16, 21, 3) {real, imag} */,
  {32'h3e455310, 32'h00000000} /* (16, 21, 2) {real, imag} */,
  {32'hbcbcc8c0, 32'h00000000} /* (16, 21, 1) {real, imag} */,
  {32'hbe9363f0, 32'h00000000} /* (16, 21, 0) {real, imag} */,
  {32'hbd9f1e10, 32'h00000000} /* (16, 20, 31) {real, imag} */,
  {32'h3da47fe0, 32'h00000000} /* (16, 20, 30) {real, imag} */,
  {32'h3ebfda76, 32'h00000000} /* (16, 20, 29) {real, imag} */,
  {32'h3e297a94, 32'h00000000} /* (16, 20, 28) {real, imag} */,
  {32'hbf1a0454, 32'h00000000} /* (16, 20, 27) {real, imag} */,
  {32'hbee36802, 32'h00000000} /* (16, 20, 26) {real, imag} */,
  {32'hbee45500, 32'h00000000} /* (16, 20, 25) {real, imag} */,
  {32'hbe401a48, 32'h00000000} /* (16, 20, 24) {real, imag} */,
  {32'h3ef43564, 32'h00000000} /* (16, 20, 23) {real, imag} */,
  {32'h3e093250, 32'h00000000} /* (16, 20, 22) {real, imag} */,
  {32'hbd2a3a80, 32'h00000000} /* (16, 20, 21) {real, imag} */,
  {32'hbda037e0, 32'h00000000} /* (16, 20, 20) {real, imag} */,
  {32'h3e3c0ef8, 32'h00000000} /* (16, 20, 19) {real, imag} */,
  {32'hbe81e884, 32'h00000000} /* (16, 20, 18) {real, imag} */,
  {32'h3e583cd4, 32'h00000000} /* (16, 20, 17) {real, imag} */,
  {32'h3ef91f20, 32'h00000000} /* (16, 20, 16) {real, imag} */,
  {32'h3e513738, 32'h00000000} /* (16, 20, 15) {real, imag} */,
  {32'hbf085d60, 32'h00000000} /* (16, 20, 14) {real, imag} */,
  {32'hbe0a4c44, 32'h00000000} /* (16, 20, 13) {real, imag} */,
  {32'hbee8bbde, 32'h00000000} /* (16, 20, 12) {real, imag} */,
  {32'hbf3365ec, 32'h00000000} /* (16, 20, 11) {real, imag} */,
  {32'hbf42e9a2, 32'h00000000} /* (16, 20, 10) {real, imag} */,
  {32'h3f34d134, 32'h00000000} /* (16, 20, 9) {real, imag} */,
  {32'h3e128be8, 32'h00000000} /* (16, 20, 8) {real, imag} */,
  {32'hbfaa592c, 32'h00000000} /* (16, 20, 7) {real, imag} */,
  {32'hbe4377ac, 32'h00000000} /* (16, 20, 6) {real, imag} */,
  {32'hbee0f590, 32'h00000000} /* (16, 20, 5) {real, imag} */,
  {32'hbecdadae, 32'h00000000} /* (16, 20, 4) {real, imag} */,
  {32'h3ebc1008, 32'h00000000} /* (16, 20, 3) {real, imag} */,
  {32'h3f7741d6, 32'h00000000} /* (16, 20, 2) {real, imag} */,
  {32'hbe140a30, 32'h00000000} /* (16, 20, 1) {real, imag} */,
  {32'hbed36ad2, 32'h00000000} /* (16, 20, 0) {real, imag} */,
  {32'h3deebdf0, 32'h00000000} /* (16, 19, 31) {real, imag} */,
  {32'h3ec55e54, 32'h00000000} /* (16, 19, 30) {real, imag} */,
  {32'h3f2d0776, 32'h00000000} /* (16, 19, 29) {real, imag} */,
  {32'h3e9bcd88, 32'h00000000} /* (16, 19, 28) {real, imag} */,
  {32'hbf1259d1, 32'h00000000} /* (16, 19, 27) {real, imag} */,
  {32'hbf21fc55, 32'h00000000} /* (16, 19, 26) {real, imag} */,
  {32'hbf2aab44, 32'h00000000} /* (16, 19, 25) {real, imag} */,
  {32'h3d808540, 32'h00000000} /* (16, 19, 24) {real, imag} */,
  {32'h3f142124, 32'h00000000} /* (16, 19, 23) {real, imag} */,
  {32'h3eccdcd4, 32'h00000000} /* (16, 19, 22) {real, imag} */,
  {32'h3d36a3c0, 32'h00000000} /* (16, 19, 21) {real, imag} */,
  {32'hbd45cc28, 32'h00000000} /* (16, 19, 20) {real, imag} */,
  {32'hbd104950, 32'h00000000} /* (16, 19, 19) {real, imag} */,
  {32'hbf24fcdc, 32'h00000000} /* (16, 19, 18) {real, imag} */,
  {32'hbf7aa3ca, 32'h00000000} /* (16, 19, 17) {real, imag} */,
  {32'hbf5470de, 32'h00000000} /* (16, 19, 16) {real, imag} */,
  {32'hbf6e4288, 32'h00000000} /* (16, 19, 15) {real, imag} */,
  {32'hbf6cf8d4, 32'h00000000} /* (16, 19, 14) {real, imag} */,
  {32'hbf47dc06, 32'h00000000} /* (16, 19, 13) {real, imag} */,
  {32'hbe7ef158, 32'h00000000} /* (16, 19, 12) {real, imag} */,
  {32'hbe6865c8, 32'h00000000} /* (16, 19, 11) {real, imag} */,
  {32'h3f4c5352, 32'h00000000} /* (16, 19, 10) {real, imag} */,
  {32'h3f82982f, 32'h00000000} /* (16, 19, 9) {real, imag} */,
  {32'h3f5d5634, 32'h00000000} /* (16, 19, 8) {real, imag} */,
  {32'hbd831300, 32'h00000000} /* (16, 19, 7) {real, imag} */,
  {32'h3ebdcf20, 32'h00000000} /* (16, 19, 6) {real, imag} */,
  {32'hbe090a94, 32'h00000000} /* (16, 19, 5) {real, imag} */,
  {32'hbeb54384, 32'h00000000} /* (16, 19, 4) {real, imag} */,
  {32'h3e76f9d0, 32'h00000000} /* (16, 19, 3) {real, imag} */,
  {32'h3ec6e504, 32'h00000000} /* (16, 19, 2) {real, imag} */,
  {32'hbf0b5786, 32'h00000000} /* (16, 19, 1) {real, imag} */,
  {32'hbf79d07a, 32'h00000000} /* (16, 19, 0) {real, imag} */,
  {32'h3fa04229, 32'h00000000} /* (16, 18, 31) {real, imag} */,
  {32'h3fd5fe4e, 32'h00000000} /* (16, 18, 30) {real, imag} */,
  {32'h3f7c917e, 32'h00000000} /* (16, 18, 29) {real, imag} */,
  {32'h3e747e3a, 32'h00000000} /* (16, 18, 28) {real, imag} */,
  {32'hbf1408aa, 32'h00000000} /* (16, 18, 27) {real, imag} */,
  {32'hbf1672de, 32'h00000000} /* (16, 18, 26) {real, imag} */,
  {32'hbf028f52, 32'h00000000} /* (16, 18, 25) {real, imag} */,
  {32'h3dec3c40, 32'h00000000} /* (16, 18, 24) {real, imag} */,
  {32'h3f3c8520, 32'h00000000} /* (16, 18, 23) {real, imag} */,
  {32'h3ee5b368, 32'h00000000} /* (16, 18, 22) {real, imag} */,
  {32'h3f21a4a6, 32'h00000000} /* (16, 18, 21) {real, imag} */,
  {32'h3dce6b98, 32'h00000000} /* (16, 18, 20) {real, imag} */,
  {32'hbe82454e, 32'h00000000} /* (16, 18, 19) {real, imag} */,
  {32'hbe5dbfb8, 32'h00000000} /* (16, 18, 18) {real, imag} */,
  {32'hbf9184f4, 32'h00000000} /* (16, 18, 17) {real, imag} */,
  {32'hbf4cf42a, 32'h00000000} /* (16, 18, 16) {real, imag} */,
  {32'hbe14ad54, 32'h00000000} /* (16, 18, 15) {real, imag} */,
  {32'hbcca4500, 32'h00000000} /* (16, 18, 14) {real, imag} */,
  {32'hbf78649c, 32'h00000000} /* (16, 18, 13) {real, imag} */,
  {32'hbf4336ea, 32'h00000000} /* (16, 18, 12) {real, imag} */,
  {32'hbd873d58, 32'h00000000} /* (16, 18, 11) {real, imag} */,
  {32'h3e18225c, 32'h00000000} /* (16, 18, 10) {real, imag} */,
  {32'h3ede0980, 32'h00000000} /* (16, 18, 9) {real, imag} */,
  {32'hbea780a6, 32'h00000000} /* (16, 18, 8) {real, imag} */,
  {32'hbf05e246, 32'h00000000} /* (16, 18, 7) {real, imag} */,
  {32'h3f581e3e, 32'h00000000} /* (16, 18, 6) {real, imag} */,
  {32'h3ed6ef24, 32'h00000000} /* (16, 18, 5) {real, imag} */,
  {32'hbf0e3cc0, 32'h00000000} /* (16, 18, 4) {real, imag} */,
  {32'hbf86d5e6, 32'h00000000} /* (16, 18, 3) {real, imag} */,
  {32'hbf25de30, 32'h00000000} /* (16, 18, 2) {real, imag} */,
  {32'h3dde9120, 32'h00000000} /* (16, 18, 1) {real, imag} */,
  {32'h3db52520, 32'h00000000} /* (16, 18, 0) {real, imag} */,
  {32'h3f921b6a, 32'h00000000} /* (16, 17, 31) {real, imag} */,
  {32'h3f868ada, 32'h00000000} /* (16, 17, 30) {real, imag} */,
  {32'h3f0cec7a, 32'h00000000} /* (16, 17, 29) {real, imag} */,
  {32'hbe7a43bc, 32'h00000000} /* (16, 17, 28) {real, imag} */,
  {32'hbeffa174, 32'h00000000} /* (16, 17, 27) {real, imag} */,
  {32'hbf186480, 32'h00000000} /* (16, 17, 26) {real, imag} */,
  {32'hbf9171f5, 32'h00000000} /* (16, 17, 25) {real, imag} */,
  {32'h3dd85690, 32'h00000000} /* (16, 17, 24) {real, imag} */,
  {32'hbe004dd8, 32'h00000000} /* (16, 17, 23) {real, imag} */,
  {32'h3d666fc0, 32'h00000000} /* (16, 17, 22) {real, imag} */,
  {32'h3f10e3ee, 32'h00000000} /* (16, 17, 21) {real, imag} */,
  {32'hbe8eedaa, 32'h00000000} /* (16, 17, 20) {real, imag} */,
  {32'hbf746ac7, 32'h00000000} /* (16, 17, 19) {real, imag} */,
  {32'h3bc36100, 32'h00000000} /* (16, 17, 18) {real, imag} */,
  {32'hbf2d2a62, 32'h00000000} /* (16, 17, 17) {real, imag} */,
  {32'hbd83c4c0, 32'h00000000} /* (16, 17, 16) {real, imag} */,
  {32'hbef0a42c, 32'h00000000} /* (16, 17, 15) {real, imag} */,
  {32'hbe9b09f8, 32'h00000000} /* (16, 17, 14) {real, imag} */,
  {32'hbde34d68, 32'h00000000} /* (16, 17, 13) {real, imag} */,
  {32'hbf3d2f78, 32'h00000000} /* (16, 17, 12) {real, imag} */,
  {32'hbea050f8, 32'h00000000} /* (16, 17, 11) {real, imag} */,
  {32'hbf193dc0, 32'h00000000} /* (16, 17, 10) {real, imag} */,
  {32'h3f4ae9ce, 32'h00000000} /* (16, 17, 9) {real, imag} */,
  {32'hbd918ac0, 32'h00000000} /* (16, 17, 8) {real, imag} */,
  {32'hbf24a5bb, 32'h00000000} /* (16, 17, 7) {real, imag} */,
  {32'h3ed2f74c, 32'h00000000} /* (16, 17, 6) {real, imag} */,
  {32'h3dc9aef0, 32'h00000000} /* (16, 17, 5) {real, imag} */,
  {32'h3c40dfc0, 32'h00000000} /* (16, 17, 4) {real, imag} */,
  {32'h3eaea120, 32'h00000000} /* (16, 17, 3) {real, imag} */,
  {32'hbe1c47e0, 32'h00000000} /* (16, 17, 2) {real, imag} */,
  {32'h3e9541e0, 32'h00000000} /* (16, 17, 1) {real, imag} */,
  {32'h3f3b5094, 32'h00000000} /* (16, 17, 0) {real, imag} */,
  {32'h3e93a094, 32'h00000000} /* (16, 16, 31) {real, imag} */,
  {32'h3e944664, 32'h00000000} /* (16, 16, 30) {real, imag} */,
  {32'h3f131124, 32'h00000000} /* (16, 16, 29) {real, imag} */,
  {32'h3f1aace3, 32'h00000000} /* (16, 16, 28) {real, imag} */,
  {32'h3f4498a2, 32'h00000000} /* (16, 16, 27) {real, imag} */,
  {32'h3eb91c3c, 32'h00000000} /* (16, 16, 26) {real, imag} */,
  {32'h3bd73280, 32'h00000000} /* (16, 16, 25) {real, imag} */,
  {32'h3e15fd80, 32'h00000000} /* (16, 16, 24) {real, imag} */,
  {32'hbf3293a9, 32'h00000000} /* (16, 16, 23) {real, imag} */,
  {32'hbdc2cb80, 32'h00000000} /* (16, 16, 22) {real, imag} */,
  {32'h3e9e49d8, 32'h00000000} /* (16, 16, 21) {real, imag} */,
  {32'hbed9ad32, 32'h00000000} /* (16, 16, 20) {real, imag} */,
  {32'hbf43d0ca, 32'h00000000} /* (16, 16, 19) {real, imag} */,
  {32'hbd5bdb00, 32'h00000000} /* (16, 16, 18) {real, imag} */,
  {32'hbe255cb4, 32'h00000000} /* (16, 16, 17) {real, imag} */,
  {32'h3ec69944, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'h3ef742f0, 32'h00000000} /* (16, 16, 15) {real, imag} */,
  {32'h3f1e8ca2, 32'h00000000} /* (16, 16, 14) {real, imag} */,
  {32'h3f982a3e, 32'h00000000} /* (16, 16, 13) {real, imag} */,
  {32'hbed76690, 32'h00000000} /* (16, 16, 12) {real, imag} */,
  {32'hbea5c720, 32'h00000000} /* (16, 16, 11) {real, imag} */,
  {32'h3d1ea890, 32'h00000000} /* (16, 16, 10) {real, imag} */,
  {32'h3f0e7164, 32'h00000000} /* (16, 16, 9) {real, imag} */,
  {32'h3f2f0692, 32'h00000000} /* (16, 16, 8) {real, imag} */,
  {32'hbe9e6620, 32'h00000000} /* (16, 16, 7) {real, imag} */,
  {32'hbec27d90, 32'h00000000} /* (16, 16, 6) {real, imag} */,
  {32'hbec40f18, 32'h00000000} /* (16, 16, 5) {real, imag} */,
  {32'hbf50a908, 32'h00000000} /* (16, 16, 4) {real, imag} */,
  {32'h3f2b9dae, 32'h00000000} /* (16, 16, 3) {real, imag} */,
  {32'hbe280ea0, 32'h00000000} /* (16, 16, 2) {real, imag} */,
  {32'hbf16e38e, 32'h00000000} /* (16, 16, 1) {real, imag} */,
  {32'h3de969b0, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'hbe4b61a8, 32'h00000000} /* (16, 15, 31) {real, imag} */,
  {32'hbf208630, 32'h00000000} /* (16, 15, 30) {real, imag} */,
  {32'h3ecbbb38, 32'h00000000} /* (16, 15, 29) {real, imag} */,
  {32'h3f97ef48, 32'h00000000} /* (16, 15, 28) {real, imag} */,
  {32'h3f2601e2, 32'h00000000} /* (16, 15, 27) {real, imag} */,
  {32'h3e40a4be, 32'h00000000} /* (16, 15, 26) {real, imag} */,
  {32'hbeda1c98, 32'h00000000} /* (16, 15, 25) {real, imag} */,
  {32'hbf3fccb5, 32'h00000000} /* (16, 15, 24) {real, imag} */,
  {32'hbfb07dac, 32'h00000000} /* (16, 15, 23) {real, imag} */,
  {32'hbe5fe204, 32'h00000000} /* (16, 15, 22) {real, imag} */,
  {32'h3ed2e378, 32'h00000000} /* (16, 15, 21) {real, imag} */,
  {32'h3ed0c82c, 32'h00000000} /* (16, 15, 20) {real, imag} */,
  {32'hbe9bbafc, 32'h00000000} /* (16, 15, 19) {real, imag} */,
  {32'hbd4b71a0, 32'h00000000} /* (16, 15, 18) {real, imag} */,
  {32'hbf0ed86a, 32'h00000000} /* (16, 15, 17) {real, imag} */,
  {32'hbe861c60, 32'h00000000} /* (16, 15, 16) {real, imag} */,
  {32'hbde4a990, 32'h00000000} /* (16, 15, 15) {real, imag} */,
  {32'hbe99c514, 32'h00000000} /* (16, 15, 14) {real, imag} */,
  {32'h3df32cd0, 32'h00000000} /* (16, 15, 13) {real, imag} */,
  {32'hbf2c2af4, 32'h00000000} /* (16, 15, 12) {real, imag} */,
  {32'hbf4a0584, 32'h00000000} /* (16, 15, 11) {real, imag} */,
  {32'hbee28672, 32'h00000000} /* (16, 15, 10) {real, imag} */,
  {32'hbef40730, 32'h00000000} /* (16, 15, 9) {real, imag} */,
  {32'hbf2742d2, 32'h00000000} /* (16, 15, 8) {real, imag} */,
  {32'hbec9a550, 32'h00000000} /* (16, 15, 7) {real, imag} */,
  {32'hbf990d78, 32'h00000000} /* (16, 15, 6) {real, imag} */,
  {32'hbfb2209b, 32'h00000000} /* (16, 15, 5) {real, imag} */,
  {32'hbf5bfa2c, 32'h00000000} /* (16, 15, 4) {real, imag} */,
  {32'hbe001580, 32'h00000000} /* (16, 15, 3) {real, imag} */,
  {32'hbeb4b9cc, 32'h00000000} /* (16, 15, 2) {real, imag} */,
  {32'hbe871b20, 32'h00000000} /* (16, 15, 1) {real, imag} */,
  {32'hbec7bbfc, 32'h00000000} /* (16, 15, 0) {real, imag} */,
  {32'h3f1bcfc6, 32'h00000000} /* (16, 14, 31) {real, imag} */,
  {32'h3caea480, 32'h00000000} /* (16, 14, 30) {real, imag} */,
  {32'h3cde2280, 32'h00000000} /* (16, 14, 29) {real, imag} */,
  {32'h3d28abe0, 32'h00000000} /* (16, 14, 28) {real, imag} */,
  {32'hbe124b24, 32'h00000000} /* (16, 14, 27) {real, imag} */,
  {32'h3f07a372, 32'h00000000} /* (16, 14, 26) {real, imag} */,
  {32'h3debfac0, 32'h00000000} /* (16, 14, 25) {real, imag} */,
  {32'hbecf8f60, 32'h00000000} /* (16, 14, 24) {real, imag} */,
  {32'h3e3264c8, 32'h00000000} /* (16, 14, 23) {real, imag} */,
  {32'h3eb612c8, 32'h00000000} /* (16, 14, 22) {real, imag} */,
  {32'h3e364520, 32'h00000000} /* (16, 14, 21) {real, imag} */,
  {32'h3f166636, 32'h00000000} /* (16, 14, 20) {real, imag} */,
  {32'h3eb35780, 32'h00000000} /* (16, 14, 19) {real, imag} */,
  {32'h3eb57650, 32'h00000000} /* (16, 14, 18) {real, imag} */,
  {32'h3f48c57e, 32'h00000000} /* (16, 14, 17) {real, imag} */,
  {32'h3f4762fc, 32'h00000000} /* (16, 14, 16) {real, imag} */,
  {32'h3de0c910, 32'h00000000} /* (16, 14, 15) {real, imag} */,
  {32'hbef445c0, 32'h00000000} /* (16, 14, 14) {real, imag} */,
  {32'hbe5f8204, 32'h00000000} /* (16, 14, 13) {real, imag} */,
  {32'hbf6d508d, 32'h00000000} /* (16, 14, 12) {real, imag} */,
  {32'h3d3627e0, 32'h00000000} /* (16, 14, 11) {real, imag} */,
  {32'h3d718e80, 32'h00000000} /* (16, 14, 10) {real, imag} */,
  {32'hbd1db810, 32'h00000000} /* (16, 14, 9) {real, imag} */,
  {32'hbe62605c, 32'h00000000} /* (16, 14, 8) {real, imag} */,
  {32'hbf02ede8, 32'h00000000} /* (16, 14, 7) {real, imag} */,
  {32'hbf905207, 32'h00000000} /* (16, 14, 6) {real, imag} */,
  {32'hbf413386, 32'h00000000} /* (16, 14, 5) {real, imag} */,
  {32'hbe85c128, 32'h00000000} /* (16, 14, 4) {real, imag} */,
  {32'h3e7957c0, 32'h00000000} /* (16, 14, 3) {real, imag} */,
  {32'hbe02be18, 32'h00000000} /* (16, 14, 2) {real, imag} */,
  {32'hbe18f948, 32'h00000000} /* (16, 14, 1) {real, imag} */,
  {32'hbda30e08, 32'h00000000} /* (16, 14, 0) {real, imag} */,
  {32'h3f279846, 32'h00000000} /* (16, 13, 31) {real, imag} */,
  {32'h3e5c87b0, 32'h00000000} /* (16, 13, 30) {real, imag} */,
  {32'hbe6d8b50, 32'h00000000} /* (16, 13, 29) {real, imag} */,
  {32'hbf32b1c0, 32'h00000000} /* (16, 13, 28) {real, imag} */,
  {32'hbf17370a, 32'h00000000} /* (16, 13, 27) {real, imag} */,
  {32'h3f221f10, 32'h00000000} /* (16, 13, 26) {real, imag} */,
  {32'h3f052958, 32'h00000000} /* (16, 13, 25) {real, imag} */,
  {32'hbdd565c0, 32'h00000000} /* (16, 13, 24) {real, imag} */,
  {32'h3ee2b792, 32'h00000000} /* (16, 13, 23) {real, imag} */,
  {32'hbf598f54, 32'h00000000} /* (16, 13, 22) {real, imag} */,
  {32'hbecc4260, 32'h00000000} /* (16, 13, 21) {real, imag} */,
  {32'h3f9a7048, 32'h00000000} /* (16, 13, 20) {real, imag} */,
  {32'hbd7c4180, 32'h00000000} /* (16, 13, 19) {real, imag} */,
  {32'h3d1c31e0, 32'h00000000} /* (16, 13, 18) {real, imag} */,
  {32'h3fe0686a, 32'h00000000} /* (16, 13, 17) {real, imag} */,
  {32'h3fc922f5, 32'h00000000} /* (16, 13, 16) {real, imag} */,
  {32'h3f69d408, 32'h00000000} /* (16, 13, 15) {real, imag} */,
  {32'hbda8c580, 32'h00000000} /* (16, 13, 14) {real, imag} */,
  {32'h3efa02b0, 32'h00000000} /* (16, 13, 13) {real, imag} */,
  {32'h3ea96b2e, 32'h00000000} /* (16, 13, 12) {real, imag} */,
  {32'h3f1bf3d5, 32'h00000000} /* (16, 13, 11) {real, imag} */,
  {32'h3d8b7a8c, 32'h00000000} /* (16, 13, 10) {real, imag} */,
  {32'hbdd1b260, 32'h00000000} /* (16, 13, 9) {real, imag} */,
  {32'h3e1d29c0, 32'h00000000} /* (16, 13, 8) {real, imag} */,
  {32'hbf13b534, 32'h00000000} /* (16, 13, 7) {real, imag} */,
  {32'hbee08610, 32'h00000000} /* (16, 13, 6) {real, imag} */,
  {32'hbe0d7ea4, 32'h00000000} /* (16, 13, 5) {real, imag} */,
  {32'hbd4be7a0, 32'h00000000} /* (16, 13, 4) {real, imag} */,
  {32'h3eda181c, 32'h00000000} /* (16, 13, 3) {real, imag} */,
  {32'hbf07aa80, 32'h00000000} /* (16, 13, 2) {real, imag} */,
  {32'hbf5d82a0, 32'h00000000} /* (16, 13, 1) {real, imag} */,
  {32'h3e8bda6a, 32'h00000000} /* (16, 13, 0) {real, imag} */,
  {32'hbd0addd0, 32'h00000000} /* (16, 12, 31) {real, imag} */,
  {32'hbf133632, 32'h00000000} /* (16, 12, 30) {real, imag} */,
  {32'hbf03bd10, 32'h00000000} /* (16, 12, 29) {real, imag} */,
  {32'h3ed2603a, 32'h00000000} /* (16, 12, 28) {real, imag} */,
  {32'h3f48b2ca, 32'h00000000} /* (16, 12, 27) {real, imag} */,
  {32'hbd2bc030, 32'h00000000} /* (16, 12, 26) {real, imag} */,
  {32'hbe219fe0, 32'h00000000} /* (16, 12, 25) {real, imag} */,
  {32'hbedd1e7c, 32'h00000000} /* (16, 12, 24) {real, imag} */,
  {32'hbd984ad0, 32'h00000000} /* (16, 12, 23) {real, imag} */,
  {32'hbf8c8f4c, 32'h00000000} /* (16, 12, 22) {real, imag} */,
  {32'hbf2f3710, 32'h00000000} /* (16, 12, 21) {real, imag} */,
  {32'h3f1ee54b, 32'h00000000} /* (16, 12, 20) {real, imag} */,
  {32'hbeefd0c8, 32'h00000000} /* (16, 12, 19) {real, imag} */,
  {32'h3e3da7cc, 32'h00000000} /* (16, 12, 18) {real, imag} */,
  {32'h40048332, 32'h00000000} /* (16, 12, 17) {real, imag} */,
  {32'h3f8aa4d0, 32'h00000000} /* (16, 12, 16) {real, imag} */,
  {32'h3e9c42d0, 32'h00000000} /* (16, 12, 15) {real, imag} */,
  {32'h3db42ec0, 32'h00000000} /* (16, 12, 14) {real, imag} */,
  {32'h3f419b21, 32'h00000000} /* (16, 12, 13) {real, imag} */,
  {32'hbe930568, 32'h00000000} /* (16, 12, 12) {real, imag} */,
  {32'hbf000952, 32'h00000000} /* (16, 12, 11) {real, imag} */,
  {32'hbe33e770, 32'h00000000} /* (16, 12, 10) {real, imag} */,
  {32'hbe97a40a, 32'h00000000} /* (16, 12, 9) {real, imag} */,
  {32'h3e90a5a0, 32'h00000000} /* (16, 12, 8) {real, imag} */,
  {32'h3e7c74c0, 32'h00000000} /* (16, 12, 7) {real, imag} */,
  {32'h3e9590c4, 32'h00000000} /* (16, 12, 6) {real, imag} */,
  {32'hbe27f1a0, 32'h00000000} /* (16, 12, 5) {real, imag} */,
  {32'hbf1d5e62, 32'h00000000} /* (16, 12, 4) {real, imag} */,
  {32'hbf716185, 32'h00000000} /* (16, 12, 3) {real, imag} */,
  {32'hbf52ca34, 32'h00000000} /* (16, 12, 2) {real, imag} */,
  {32'hbf5d61ae, 32'h00000000} /* (16, 12, 1) {real, imag} */,
  {32'h3e88c280, 32'h00000000} /* (16, 12, 0) {real, imag} */,
  {32'h3d6dd0c0, 32'h00000000} /* (16, 11, 31) {real, imag} */,
  {32'h3e5ed860, 32'h00000000} /* (16, 11, 30) {real, imag} */,
  {32'hbf42fc4d, 32'h00000000} /* (16, 11, 29) {real, imag} */,
  {32'hbedb676e, 32'h00000000} /* (16, 11, 28) {real, imag} */,
  {32'h3f11c97b, 32'h00000000} /* (16, 11, 27) {real, imag} */,
  {32'hbebde35c, 32'h00000000} /* (16, 11, 26) {real, imag} */,
  {32'hbf4ea814, 32'h00000000} /* (16, 11, 25) {real, imag} */,
  {32'hbcfdd3e0, 32'h00000000} /* (16, 11, 24) {real, imag} */,
  {32'h3f6644f6, 32'h00000000} /* (16, 11, 23) {real, imag} */,
  {32'hbcf5ee00, 32'h00000000} /* (16, 11, 22) {real, imag} */,
  {32'hbedcc160, 32'h00000000} /* (16, 11, 21) {real, imag} */,
  {32'hbf2d42e6, 32'h00000000} /* (16, 11, 20) {real, imag} */,
  {32'hbe2d3ce0, 32'h00000000} /* (16, 11, 19) {real, imag} */,
  {32'hbf42408e, 32'h00000000} /* (16, 11, 18) {real, imag} */,
  {32'h3e9c6588, 32'h00000000} /* (16, 11, 17) {real, imag} */,
  {32'h3ef3abb0, 32'h00000000} /* (16, 11, 16) {real, imag} */,
  {32'h3e97e422, 32'h00000000} /* (16, 11, 15) {real, imag} */,
  {32'hbf0eb042, 32'h00000000} /* (16, 11, 14) {real, imag} */,
  {32'h3e47709c, 32'h00000000} /* (16, 11, 13) {real, imag} */,
  {32'hbda60344, 32'h00000000} /* (16, 11, 12) {real, imag} */,
  {32'hbdf01ee8, 32'h00000000} /* (16, 11, 11) {real, imag} */,
  {32'hbd9f6098, 32'h00000000} /* (16, 11, 10) {real, imag} */,
  {32'hbea350c2, 32'h00000000} /* (16, 11, 9) {real, imag} */,
  {32'h3f958f49, 32'h00000000} /* (16, 11, 8) {real, imag} */,
  {32'h3f8f95c8, 32'h00000000} /* (16, 11, 7) {real, imag} */,
  {32'h3ece401a, 32'h00000000} /* (16, 11, 6) {real, imag} */,
  {32'hbf546f24, 32'h00000000} /* (16, 11, 5) {real, imag} */,
  {32'hbee53c98, 32'h00000000} /* (16, 11, 4) {real, imag} */,
  {32'h3e962ab2, 32'h00000000} /* (16, 11, 3) {real, imag} */,
  {32'hbf0ae694, 32'h00000000} /* (16, 11, 2) {real, imag} */,
  {32'hbf3e1b41, 32'h00000000} /* (16, 11, 1) {real, imag} */,
  {32'hbe0213d8, 32'h00000000} /* (16, 11, 0) {real, imag} */,
  {32'hbf106acc, 32'h00000000} /* (16, 10, 31) {real, imag} */,
  {32'hbf04687c, 32'h00000000} /* (16, 10, 30) {real, imag} */,
  {32'h3d0fc840, 32'h00000000} /* (16, 10, 29) {real, imag} */,
  {32'hbed244e4, 32'h00000000} /* (16, 10, 28) {real, imag} */,
  {32'h3e1308a0, 32'h00000000} /* (16, 10, 27) {real, imag} */,
  {32'h3dcf2730, 32'h00000000} /* (16, 10, 26) {real, imag} */,
  {32'h3cf92160, 32'h00000000} /* (16, 10, 25) {real, imag} */,
  {32'h3f804230, 32'h00000000} /* (16, 10, 24) {real, imag} */,
  {32'h3f862c36, 32'h00000000} /* (16, 10, 23) {real, imag} */,
  {32'hbe252130, 32'h00000000} /* (16, 10, 22) {real, imag} */,
  {32'hbe98f700, 32'h00000000} /* (16, 10, 21) {real, imag} */,
  {32'hbe3bf050, 32'h00000000} /* (16, 10, 20) {real, imag} */,
  {32'h3d895490, 32'h00000000} /* (16, 10, 19) {real, imag} */,
  {32'hbea866dc, 32'h00000000} /* (16, 10, 18) {real, imag} */,
  {32'hbe7bb290, 32'h00000000} /* (16, 10, 17) {real, imag} */,
  {32'h3f2e3c3c, 32'h00000000} /* (16, 10, 16) {real, imag} */,
  {32'h3f815f97, 32'h00000000} /* (16, 10, 15) {real, imag} */,
  {32'hbf23fe37, 32'h00000000} /* (16, 10, 14) {real, imag} */,
  {32'hbe2dd1d2, 32'h00000000} /* (16, 10, 13) {real, imag} */,
  {32'h3eb2d73a, 32'h00000000} /* (16, 10, 12) {real, imag} */,
  {32'h3e1718f0, 32'h00000000} /* (16, 10, 11) {real, imag} */,
  {32'hbedbced8, 32'h00000000} /* (16, 10, 10) {real, imag} */,
  {32'hbec41454, 32'h00000000} /* (16, 10, 9) {real, imag} */,
  {32'h3ea98454, 32'h00000000} /* (16, 10, 8) {real, imag} */,
  {32'hbf0d4554, 32'h00000000} /* (16, 10, 7) {real, imag} */,
  {32'h3ccf1800, 32'h00000000} /* (16, 10, 6) {real, imag} */,
  {32'hbe1b35a0, 32'h00000000} /* (16, 10, 5) {real, imag} */,
  {32'h3e48dff8, 32'h00000000} /* (16, 10, 4) {real, imag} */,
  {32'h3ed6dfd0, 32'h00000000} /* (16, 10, 3) {real, imag} */,
  {32'h3d92c840, 32'h00000000} /* (16, 10, 2) {real, imag} */,
  {32'h3e2a6368, 32'h00000000} /* (16, 10, 1) {real, imag} */,
  {32'hbcc5ade0, 32'h00000000} /* (16, 10, 0) {real, imag} */,
  {32'hbe92594a, 32'h00000000} /* (16, 9, 31) {real, imag} */,
  {32'h3c09f500, 32'h00000000} /* (16, 9, 30) {real, imag} */,
  {32'h3d8658b0, 32'h00000000} /* (16, 9, 29) {real, imag} */,
  {32'hbea8f168, 32'h00000000} /* (16, 9, 28) {real, imag} */,
  {32'h3e7ceba4, 32'h00000000} /* (16, 9, 27) {real, imag} */,
  {32'h3f0eb1fe, 32'h00000000} /* (16, 9, 26) {real, imag} */,
  {32'h3f06390a, 32'h00000000} /* (16, 9, 25) {real, imag} */,
  {32'h3f47d412, 32'h00000000} /* (16, 9, 24) {real, imag} */,
  {32'h3d951b78, 32'h00000000} /* (16, 9, 23) {real, imag} */,
  {32'hbe74b450, 32'h00000000} /* (16, 9, 22) {real, imag} */,
  {32'h3f0b5597, 32'h00000000} /* (16, 9, 21) {real, imag} */,
  {32'hbef2cd80, 32'h00000000} /* (16, 9, 20) {real, imag} */,
  {32'hbf5cb7b1, 32'h00000000} /* (16, 9, 19) {real, imag} */,
  {32'h3cdc31c0, 32'h00000000} /* (16, 9, 18) {real, imag} */,
  {32'hbf2b82af, 32'h00000000} /* (16, 9, 17) {real, imag} */,
  {32'hbec63788, 32'h00000000} /* (16, 9, 16) {real, imag} */,
  {32'hbeb583c8, 32'h00000000} /* (16, 9, 15) {real, imag} */,
  {32'hbf3ab9e0, 32'h00000000} /* (16, 9, 14) {real, imag} */,
  {32'h3e258f90, 32'h00000000} /* (16, 9, 13) {real, imag} */,
  {32'h3eb335e6, 32'h00000000} /* (16, 9, 12) {real, imag} */,
  {32'h3db17680, 32'h00000000} /* (16, 9, 11) {real, imag} */,
  {32'h3f06cc00, 32'h00000000} /* (16, 9, 10) {real, imag} */,
  {32'h3f519998, 32'h00000000} /* (16, 9, 9) {real, imag} */,
  {32'h3f3d94e4, 32'h00000000} /* (16, 9, 8) {real, imag} */,
  {32'h3d55b840, 32'h00000000} /* (16, 9, 7) {real, imag} */,
  {32'h3d6a5590, 32'h00000000} /* (16, 9, 6) {real, imag} */,
  {32'h3e906e4c, 32'h00000000} /* (16, 9, 5) {real, imag} */,
  {32'hbe8d0a72, 32'h00000000} /* (16, 9, 4) {real, imag} */,
  {32'hbe6245a8, 32'h00000000} /* (16, 9, 3) {real, imag} */,
  {32'h3e993530, 32'h00000000} /* (16, 9, 2) {real, imag} */,
  {32'hbe840e84, 32'h00000000} /* (16, 9, 1) {real, imag} */,
  {32'hbf3f13d0, 32'h00000000} /* (16, 9, 0) {real, imag} */,
  {32'h3ec10e69, 32'h00000000} /* (16, 8, 31) {real, imag} */,
  {32'hbdfdfccc, 32'h00000000} /* (16, 8, 30) {real, imag} */,
  {32'hbe69c078, 32'h00000000} /* (16, 8, 29) {real, imag} */,
  {32'hbe278f40, 32'h00000000} /* (16, 8, 28) {real, imag} */,
  {32'h3e531000, 32'h00000000} /* (16, 8, 27) {real, imag} */,
  {32'h3db40bc8, 32'h00000000} /* (16, 8, 26) {real, imag} */,
  {32'h3e3f02b0, 32'h00000000} /* (16, 8, 25) {real, imag} */,
  {32'h3fb35d6e, 32'h00000000} /* (16, 8, 24) {real, imag} */,
  {32'h3eadba7c, 32'h00000000} /* (16, 8, 23) {real, imag} */,
  {32'hbf1b670c, 32'h00000000} /* (16, 8, 22) {real, imag} */,
  {32'hbec9b456, 32'h00000000} /* (16, 8, 21) {real, imag} */,
  {32'hbf0eee47, 32'h00000000} /* (16, 8, 20) {real, imag} */,
  {32'hbeaf20e8, 32'h00000000} /* (16, 8, 19) {real, imag} */,
  {32'hbebc5ef2, 32'h00000000} /* (16, 8, 18) {real, imag} */,
  {32'hbf55c7c3, 32'h00000000} /* (16, 8, 17) {real, imag} */,
  {32'hbf8409f5, 32'h00000000} /* (16, 8, 16) {real, imag} */,
  {32'hbf936103, 32'h00000000} /* (16, 8, 15) {real, imag} */,
  {32'hbf4a5620, 32'h00000000} /* (16, 8, 14) {real, imag} */,
  {32'hbea1e000, 32'h00000000} /* (16, 8, 13) {real, imag} */,
  {32'hbef1cb70, 32'h00000000} /* (16, 8, 12) {real, imag} */,
  {32'hbe2715b4, 32'h00000000} /* (16, 8, 11) {real, imag} */,
  {32'h3fd861f0, 32'h00000000} /* (16, 8, 10) {real, imag} */,
  {32'h3f884d22, 32'h00000000} /* (16, 8, 9) {real, imag} */,
  {32'h3d81aef0, 32'h00000000} /* (16, 8, 8) {real, imag} */,
  {32'h3eae79c8, 32'h00000000} /* (16, 8, 7) {real, imag} */,
  {32'hbe259010, 32'h00000000} /* (16, 8, 6) {real, imag} */,
  {32'hbd7cec40, 32'h00000000} /* (16, 8, 5) {real, imag} */,
  {32'hbec687fc, 32'h00000000} /* (16, 8, 4) {real, imag} */,
  {32'h3e97dde8, 32'h00000000} /* (16, 8, 3) {real, imag} */,
  {32'h3ee70aee, 32'h00000000} /* (16, 8, 2) {real, imag} */,
  {32'h3d549fc0, 32'h00000000} /* (16, 8, 1) {real, imag} */,
  {32'hbe8b2eac, 32'h00000000} /* (16, 8, 0) {real, imag} */,
  {32'h3ed1483a, 32'h00000000} /* (16, 7, 31) {real, imag} */,
  {32'hbe522260, 32'h00000000} /* (16, 7, 30) {real, imag} */,
  {32'h3ee571d0, 32'h00000000} /* (16, 7, 29) {real, imag} */,
  {32'h3ea2d150, 32'h00000000} /* (16, 7, 28) {real, imag} */,
  {32'h3eb94d54, 32'h00000000} /* (16, 7, 27) {real, imag} */,
  {32'h3e3cc7e0, 32'h00000000} /* (16, 7, 26) {real, imag} */,
  {32'h3d89d5c0, 32'h00000000} /* (16, 7, 25) {real, imag} */,
  {32'h3f2313fa, 32'h00000000} /* (16, 7, 24) {real, imag} */,
  {32'h3f1e718a, 32'h00000000} /* (16, 7, 23) {real, imag} */,
  {32'h3e83d9f0, 32'h00000000} /* (16, 7, 22) {real, imag} */,
  {32'hbd28c2c0, 32'h00000000} /* (16, 7, 21) {real, imag} */,
  {32'h3da72528, 32'h00000000} /* (16, 7, 20) {real, imag} */,
  {32'h3ecbed56, 32'h00000000} /* (16, 7, 19) {real, imag} */,
  {32'hbf320e7c, 32'h00000000} /* (16, 7, 18) {real, imag} */,
  {32'hbf86e3ab, 32'h00000000} /* (16, 7, 17) {real, imag} */,
  {32'hbfe7661f, 32'h00000000} /* (16, 7, 16) {real, imag} */,
  {32'hbfa6404a, 32'h00000000} /* (16, 7, 15) {real, imag} */,
  {32'hbe290a98, 32'h00000000} /* (16, 7, 14) {real, imag} */,
  {32'h3df2d220, 32'h00000000} /* (16, 7, 13) {real, imag} */,
  {32'h3d814138, 32'h00000000} /* (16, 7, 12) {real, imag} */,
  {32'h3e3636b0, 32'h00000000} /* (16, 7, 11) {real, imag} */,
  {32'h3f76508c, 32'h00000000} /* (16, 7, 10) {real, imag} */,
  {32'h3f7cbbcc, 32'h00000000} /* (16, 7, 9) {real, imag} */,
  {32'h3ee1afb8, 32'h00000000} /* (16, 7, 8) {real, imag} */,
  {32'hbe2347d0, 32'h00000000} /* (16, 7, 7) {real, imag} */,
  {32'hbe5e4ee0, 32'h00000000} /* (16, 7, 6) {real, imag} */,
  {32'hbe401cd8, 32'h00000000} /* (16, 7, 5) {real, imag} */,
  {32'h3f5132b0, 32'h00000000} /* (16, 7, 4) {real, imag} */,
  {32'h3f8da834, 32'h00000000} /* (16, 7, 3) {real, imag} */,
  {32'h3f5d02f2, 32'h00000000} /* (16, 7, 2) {real, imag} */,
  {32'h3f0ffd44, 32'h00000000} /* (16, 7, 1) {real, imag} */,
  {32'h3ec0feb8, 32'h00000000} /* (16, 7, 0) {real, imag} */,
  {32'h3c511b80, 32'h00000000} /* (16, 6, 31) {real, imag} */,
  {32'hbefd5f26, 32'h00000000} /* (16, 6, 30) {real, imag} */,
  {32'hbe57c360, 32'h00000000} /* (16, 6, 29) {real, imag} */,
  {32'hbf252fb6, 32'h00000000} /* (16, 6, 28) {real, imag} */,
  {32'hbefe40d4, 32'h00000000} /* (16, 6, 27) {real, imag} */,
  {32'hbc475580, 32'h00000000} /* (16, 6, 26) {real, imag} */,
  {32'h3eff0828, 32'h00000000} /* (16, 6, 25) {real, imag} */,
  {32'h3db428a0, 32'h00000000} /* (16, 6, 24) {real, imag} */,
  {32'hbecb8c44, 32'h00000000} /* (16, 6, 23) {real, imag} */,
  {32'hbe4639a0, 32'h00000000} /* (16, 6, 22) {real, imag} */,
  {32'h3efbc222, 32'h00000000} /* (16, 6, 21) {real, imag} */,
  {32'h3e967082, 32'h00000000} /* (16, 6, 20) {real, imag} */,
  {32'h3f1731db, 32'h00000000} /* (16, 6, 19) {real, imag} */,
  {32'h3f089fba, 32'h00000000} /* (16, 6, 18) {real, imag} */,
  {32'h3d7e1d10, 32'h00000000} /* (16, 6, 17) {real, imag} */,
  {32'hbf69f2b1, 32'h00000000} /* (16, 6, 16) {real, imag} */,
  {32'hbf5676c9, 32'h00000000} /* (16, 6, 15) {real, imag} */,
  {32'hbfb72c08, 32'h00000000} /* (16, 6, 14) {real, imag} */,
  {32'hbda14670, 32'h00000000} /* (16, 6, 13) {real, imag} */,
  {32'h3f44f9b0, 32'h00000000} /* (16, 6, 12) {real, imag} */,
  {32'h3e43fa70, 32'h00000000} /* (16, 6, 11) {real, imag} */,
  {32'h3f395948, 32'h00000000} /* (16, 6, 10) {real, imag} */,
  {32'h3f6e2b18, 32'h00000000} /* (16, 6, 9) {real, imag} */,
  {32'hbec64104, 32'h00000000} /* (16, 6, 8) {real, imag} */,
  {32'hbf4139ea, 32'h00000000} /* (16, 6, 7) {real, imag} */,
  {32'hbe543440, 32'h00000000} /* (16, 6, 6) {real, imag} */,
  {32'h3e2e00e0, 32'h00000000} /* (16, 6, 5) {real, imag} */,
  {32'h3f9156cc, 32'h00000000} /* (16, 6, 4) {real, imag} */,
  {32'h3fb01cd6, 32'h00000000} /* (16, 6, 3) {real, imag} */,
  {32'h3f3204b3, 32'h00000000} /* (16, 6, 2) {real, imag} */,
  {32'hbeb88440, 32'h00000000} /* (16, 6, 1) {real, imag} */,
  {32'h3c993fa0, 32'h00000000} /* (16, 6, 0) {real, imag} */,
  {32'hbdaabab0, 32'h00000000} /* (16, 5, 31) {real, imag} */,
  {32'hbf177310, 32'h00000000} /* (16, 5, 30) {real, imag} */,
  {32'hbf249274, 32'h00000000} /* (16, 5, 29) {real, imag} */,
  {32'hbf14f1f2, 32'h00000000} /* (16, 5, 28) {real, imag} */,
  {32'hbfafad56, 32'h00000000} /* (16, 5, 27) {real, imag} */,
  {32'hbfa1488b, 32'h00000000} /* (16, 5, 26) {real, imag} */,
  {32'hbe9f8260, 32'h00000000} /* (16, 5, 25) {real, imag} */,
  {32'h3e0cf570, 32'h00000000} /* (16, 5, 24) {real, imag} */,
  {32'hbf38289b, 32'h00000000} /* (16, 5, 23) {real, imag} */,
  {32'hbf068524, 32'h00000000} /* (16, 5, 22) {real, imag} */,
  {32'h3f2183b8, 32'h00000000} /* (16, 5, 21) {real, imag} */,
  {32'h3f041bc6, 32'h00000000} /* (16, 5, 20) {real, imag} */,
  {32'h3f27c369, 32'h00000000} /* (16, 5, 19) {real, imag} */,
  {32'h3f02059a, 32'h00000000} /* (16, 5, 18) {real, imag} */,
  {32'h3d982448, 32'h00000000} /* (16, 5, 17) {real, imag} */,
  {32'hbeee0a62, 32'h00000000} /* (16, 5, 16) {real, imag} */,
  {32'hbeca1608, 32'h00000000} /* (16, 5, 15) {real, imag} */,
  {32'hbed2a2e8, 32'h00000000} /* (16, 5, 14) {real, imag} */,
  {32'h3dc2e388, 32'h00000000} /* (16, 5, 13) {real, imag} */,
  {32'h3f5c6328, 32'h00000000} /* (16, 5, 12) {real, imag} */,
  {32'h3e9c64f8, 32'h00000000} /* (16, 5, 11) {real, imag} */,
  {32'hbdd443d8, 32'h00000000} /* (16, 5, 10) {real, imag} */,
  {32'h3e2cb076, 32'h00000000} /* (16, 5, 9) {real, imag} */,
  {32'hbe9610e0, 32'h00000000} /* (16, 5, 8) {real, imag} */,
  {32'hbc4a1cc0, 32'h00000000} /* (16, 5, 7) {real, imag} */,
  {32'hbf060455, 32'h00000000} /* (16, 5, 6) {real, imag} */,
  {32'h3e9c5b44, 32'h00000000} /* (16, 5, 5) {real, imag} */,
  {32'hbebc587e, 32'h00000000} /* (16, 5, 4) {real, imag} */,
  {32'hbf485e66, 32'h00000000} /* (16, 5, 3) {real, imag} */,
  {32'h3ee8bcf0, 32'h00000000} /* (16, 5, 2) {real, imag} */,
  {32'h3deddab0, 32'h00000000} /* (16, 5, 1) {real, imag} */,
  {32'hbcf76620, 32'h00000000} /* (16, 5, 0) {real, imag} */,
  {32'h3d66e460, 32'h00000000} /* (16, 4, 31) {real, imag} */,
  {32'hbe2dda20, 32'h00000000} /* (16, 4, 30) {real, imag} */,
  {32'hbf61cdc0, 32'h00000000} /* (16, 4, 29) {real, imag} */,
  {32'hbe928ea0, 32'h00000000} /* (16, 4, 28) {real, imag} */,
  {32'h3f0e0e30, 32'h00000000} /* (16, 4, 27) {real, imag} */,
  {32'h3e39a968, 32'h00000000} /* (16, 4, 26) {real, imag} */,
  {32'hbdd00a80, 32'h00000000} /* (16, 4, 25) {real, imag} */,
  {32'hbeabde80, 32'h00000000} /* (16, 4, 24) {real, imag} */,
  {32'hbf57af93, 32'h00000000} /* (16, 4, 23) {real, imag} */,
  {32'hbf31e6bc, 32'h00000000} /* (16, 4, 22) {real, imag} */,
  {32'hbea44cb0, 32'h00000000} /* (16, 4, 21) {real, imag} */,
  {32'hbf4889f6, 32'h00000000} /* (16, 4, 20) {real, imag} */,
  {32'hbde88790, 32'h00000000} /* (16, 4, 19) {real, imag} */,
  {32'h3d41b580, 32'h00000000} /* (16, 4, 18) {real, imag} */,
  {32'hbf078c0a, 32'h00000000} /* (16, 4, 17) {real, imag} */,
  {32'hbf353b88, 32'h00000000} /* (16, 4, 16) {real, imag} */,
  {32'h3e1ecea0, 32'h00000000} /* (16, 4, 15) {real, imag} */,
  {32'h3ee89cbc, 32'h00000000} /* (16, 4, 14) {real, imag} */,
  {32'h3f68f00a, 32'h00000000} /* (16, 4, 13) {real, imag} */,
  {32'h3f9143ee, 32'h00000000} /* (16, 4, 12) {real, imag} */,
  {32'h3fddac06, 32'h00000000} /* (16, 4, 11) {real, imag} */,
  {32'h3e944620, 32'h00000000} /* (16, 4, 10) {real, imag} */,
  {32'h3df17c70, 32'h00000000} /* (16, 4, 9) {real, imag} */,
  {32'h3f41b520, 32'h00000000} /* (16, 4, 8) {real, imag} */,
  {32'h3ed97510, 32'h00000000} /* (16, 4, 7) {real, imag} */,
  {32'h3df2abe0, 32'h00000000} /* (16, 4, 6) {real, imag} */,
  {32'h3f2e7398, 32'h00000000} /* (16, 4, 5) {real, imag} */,
  {32'hbe91b68a, 32'h00000000} /* (16, 4, 4) {real, imag} */,
  {32'hbf584656, 32'h00000000} /* (16, 4, 3) {real, imag} */,
  {32'h3ee1f2bc, 32'h00000000} /* (16, 4, 2) {real, imag} */,
  {32'h3df0e270, 32'h00000000} /* (16, 4, 1) {real, imag} */,
  {32'hbf51155e, 32'h00000000} /* (16, 4, 0) {real, imag} */,
  {32'h3f397dcb, 32'h00000000} /* (16, 3, 31) {real, imag} */,
  {32'h3f57b7bb, 32'h00000000} /* (16, 3, 30) {real, imag} */,
  {32'h3e3d9c58, 32'h00000000} /* (16, 3, 29) {real, imag} */,
  {32'h3f0e0fde, 32'h00000000} /* (16, 3, 28) {real, imag} */,
  {32'h3f3a83dc, 32'h00000000} /* (16, 3, 27) {real, imag} */,
  {32'h3d5a77b0, 32'h00000000} /* (16, 3, 26) {real, imag} */,
  {32'h3d314e50, 32'h00000000} /* (16, 3, 25) {real, imag} */,
  {32'h3f085828, 32'h00000000} /* (16, 3, 24) {real, imag} */,
  {32'h3e83aa50, 32'h00000000} /* (16, 3, 23) {real, imag} */,
  {32'h3e8c3700, 32'h00000000} /* (16, 3, 22) {real, imag} */,
  {32'hbede4d18, 32'h00000000} /* (16, 3, 21) {real, imag} */,
  {32'hbed53308, 32'h00000000} /* (16, 3, 20) {real, imag} */,
  {32'h3ee18374, 32'h00000000} /* (16, 3, 19) {real, imag} */,
  {32'h3f21171e, 32'h00000000} /* (16, 3, 18) {real, imag} */,
  {32'hbf201762, 32'h00000000} /* (16, 3, 17) {real, imag} */,
  {32'hbe507af0, 32'h00000000} /* (16, 3, 16) {real, imag} */,
  {32'h3e1f0230, 32'h00000000} /* (16, 3, 15) {real, imag} */,
  {32'h3ea3aa54, 32'h00000000} /* (16, 3, 14) {real, imag} */,
  {32'h3f33d344, 32'h00000000} /* (16, 3, 13) {real, imag} */,
  {32'h3eb2969c, 32'h00000000} /* (16, 3, 12) {real, imag} */,
  {32'h3f8ff25e, 32'h00000000} /* (16, 3, 11) {real, imag} */,
  {32'h3eb850f4, 32'h00000000} /* (16, 3, 10) {real, imag} */,
  {32'hbdc7aa30, 32'h00000000} /* (16, 3, 9) {real, imag} */,
  {32'hbe237470, 32'h00000000} /* (16, 3, 8) {real, imag} */,
  {32'h3d02aa00, 32'h00000000} /* (16, 3, 7) {real, imag} */,
  {32'h3edc89a2, 32'h00000000} /* (16, 3, 6) {real, imag} */,
  {32'h3f78f51c, 32'h00000000} /* (16, 3, 5) {real, imag} */,
  {32'h3e993cce, 32'h00000000} /* (16, 3, 4) {real, imag} */,
  {32'h3d83fde8, 32'h00000000} /* (16, 3, 3) {real, imag} */,
  {32'h3f332da4, 32'h00000000} /* (16, 3, 2) {real, imag} */,
  {32'h3e025408, 32'h00000000} /* (16, 3, 1) {real, imag} */,
  {32'hbdca0c60, 32'h00000000} /* (16, 3, 0) {real, imag} */,
  {32'h3e1e7544, 32'h00000000} /* (16, 2, 31) {real, imag} */,
  {32'hbd75df40, 32'h00000000} /* (16, 2, 30) {real, imag} */,
  {32'hbdb683a8, 32'h00000000} /* (16, 2, 29) {real, imag} */,
  {32'h3e3edc90, 32'h00000000} /* (16, 2, 28) {real, imag} */,
  {32'hbed39e00, 32'h00000000} /* (16, 2, 27) {real, imag} */,
  {32'hbf3901c4, 32'h00000000} /* (16, 2, 26) {real, imag} */,
  {32'h3f197b70, 32'h00000000} /* (16, 2, 25) {real, imag} */,
  {32'h3f9d01ac, 32'h00000000} /* (16, 2, 24) {real, imag} */,
  {32'h3fa770a5, 32'h00000000} /* (16, 2, 23) {real, imag} */,
  {32'h3f43eaa3, 32'h00000000} /* (16, 2, 22) {real, imag} */,
  {32'hbf857249, 32'h00000000} /* (16, 2, 21) {real, imag} */,
  {32'hbf60275a, 32'h00000000} /* (16, 2, 20) {real, imag} */,
  {32'hbf488380, 32'h00000000} /* (16, 2, 19) {real, imag} */,
  {32'h3edb62f8, 32'h00000000} /* (16, 2, 18) {real, imag} */,
  {32'hbd697720, 32'h00000000} /* (16, 2, 17) {real, imag} */,
  {32'hbc87c5c0, 32'h00000000} /* (16, 2, 16) {real, imag} */,
  {32'h3e5513f4, 32'h00000000} /* (16, 2, 15) {real, imag} */,
  {32'hbf07627b, 32'h00000000} /* (16, 2, 14) {real, imag} */,
  {32'hbf3dd64c, 32'h00000000} /* (16, 2, 13) {real, imag} */,
  {32'h3cc7a940, 32'h00000000} /* (16, 2, 12) {real, imag} */,
  {32'h3ebb6e98, 32'h00000000} /* (16, 2, 11) {real, imag} */,
  {32'h3daf7fe0, 32'h00000000} /* (16, 2, 10) {real, imag} */,
  {32'hbede2878, 32'h00000000} /* (16, 2, 9) {real, imag} */,
  {32'h3db4cec8, 32'h00000000} /* (16, 2, 8) {real, imag} */,
  {32'h3e4d50d4, 32'h00000000} /* (16, 2, 7) {real, imag} */,
  {32'h3be95200, 32'h00000000} /* (16, 2, 6) {real, imag} */,
  {32'h3f370b16, 32'h00000000} /* (16, 2, 5) {real, imag} */,
  {32'h3f4ef193, 32'h00000000} /* (16, 2, 4) {real, imag} */,
  {32'h3f59f426, 32'h00000000} /* (16, 2, 3) {real, imag} */,
  {32'h3ec96d08, 32'h00000000} /* (16, 2, 2) {real, imag} */,
  {32'hbe623588, 32'h00000000} /* (16, 2, 1) {real, imag} */,
  {32'h3d9e2750, 32'h00000000} /* (16, 2, 0) {real, imag} */,
  {32'hbf049718, 32'h00000000} /* (16, 1, 31) {real, imag} */,
  {32'hbf3cd6ea, 32'h00000000} /* (16, 1, 30) {real, imag} */,
  {32'hbf0c10ea, 32'h00000000} /* (16, 1, 29) {real, imag} */,
  {32'hbf64988a, 32'h00000000} /* (16, 1, 28) {real, imag} */,
  {32'h3c9a9500, 32'h00000000} /* (16, 1, 27) {real, imag} */,
  {32'h3f3de246, 32'h00000000} /* (16, 1, 26) {real, imag} */,
  {32'h3f4d9500, 32'h00000000} /* (16, 1, 25) {real, imag} */,
  {32'h3f191e48, 32'h00000000} /* (16, 1, 24) {real, imag} */,
  {32'h3d12e2d0, 32'h00000000} /* (16, 1, 23) {real, imag} */,
  {32'hbe15b700, 32'h00000000} /* (16, 1, 22) {real, imag} */,
  {32'hbdfe9698, 32'h00000000} /* (16, 1, 21) {real, imag} */,
  {32'hbec45a10, 32'h00000000} /* (16, 1, 20) {real, imag} */,
  {32'hbf8490b6, 32'h00000000} /* (16, 1, 19) {real, imag} */,
  {32'h3e4fa658, 32'h00000000} /* (16, 1, 18) {real, imag} */,
  {32'h3f38f9c8, 32'h00000000} /* (16, 1, 17) {real, imag} */,
  {32'h3f2c5b6c, 32'h00000000} /* (16, 1, 16) {real, imag} */,
  {32'h3dce91e8, 32'h00000000} /* (16, 1, 15) {real, imag} */,
  {32'hbf4f176a, 32'h00000000} /* (16, 1, 14) {real, imag} */,
  {32'hbf2586bd, 32'h00000000} /* (16, 1, 13) {real, imag} */,
  {32'h3f3ee9f1, 32'h00000000} /* (16, 1, 12) {real, imag} */,
  {32'h3f8a0b38, 32'h00000000} /* (16, 1, 11) {real, imag} */,
  {32'h3c9e7800, 32'h00000000} /* (16, 1, 10) {real, imag} */,
  {32'h3f049e35, 32'h00000000} /* (16, 1, 9) {real, imag} */,
  {32'h3f63b43a, 32'h00000000} /* (16, 1, 8) {real, imag} */,
  {32'h3f029fa5, 32'h00000000} /* (16, 1, 7) {real, imag} */,
  {32'h3f3d8a28, 32'h00000000} /* (16, 1, 6) {real, imag} */,
  {32'h3f398f3e, 32'h00000000} /* (16, 1, 5) {real, imag} */,
  {32'h3f550438, 32'h00000000} /* (16, 1, 4) {real, imag} */,
  {32'h3f40b4f4, 32'h00000000} /* (16, 1, 3) {real, imag} */,
  {32'hbed80d44, 32'h00000000} /* (16, 1, 2) {real, imag} */,
  {32'hbfb12564, 32'h00000000} /* (16, 1, 1) {real, imag} */,
  {32'hbfac10e4, 32'h00000000} /* (16, 1, 0) {real, imag} */,
  {32'hbdbb67f8, 32'h00000000} /* (16, 0, 31) {real, imag} */,
  {32'hbf05e48c, 32'h00000000} /* (16, 0, 30) {real, imag} */,
  {32'hbf2e3f30, 32'h00000000} /* (16, 0, 29) {real, imag} */,
  {32'hbeb9dabc, 32'h00000000} /* (16, 0, 28) {real, imag} */,
  {32'h3f63f765, 32'h00000000} /* (16, 0, 27) {real, imag} */,
  {32'h3f60b3ee, 32'h00000000} /* (16, 0, 26) {real, imag} */,
  {32'h3ef9bbc5, 32'h00000000} /* (16, 0, 25) {real, imag} */,
  {32'h3e4a8c58, 32'h00000000} /* (16, 0, 24) {real, imag} */,
  {32'hbef443e4, 32'h00000000} /* (16, 0, 23) {real, imag} */,
  {32'hbe365cc0, 32'h00000000} /* (16, 0, 22) {real, imag} */,
  {32'h3f3e3a96, 32'h00000000} /* (16, 0, 21) {real, imag} */,
  {32'h3f15b440, 32'h00000000} /* (16, 0, 20) {real, imag} */,
  {32'h3e3f4cb8, 32'h00000000} /* (16, 0, 19) {real, imag} */,
  {32'h3edd30a8, 32'h00000000} /* (16, 0, 18) {real, imag} */,
  {32'h3f06ccc6, 32'h00000000} /* (16, 0, 17) {real, imag} */,
  {32'h3e490216, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h3dbfcac4, 32'h00000000} /* (16, 0, 15) {real, imag} */,
  {32'hbd0fd500, 32'h00000000} /* (16, 0, 14) {real, imag} */,
  {32'h3e93b1ec, 32'h00000000} /* (16, 0, 13) {real, imag} */,
  {32'h3f50a87b, 32'h00000000} /* (16, 0, 12) {real, imag} */,
  {32'h3f30b428, 32'h00000000} /* (16, 0, 11) {real, imag} */,
  {32'hbe0fbb22, 32'h00000000} /* (16, 0, 10) {real, imag} */,
  {32'h3ec04561, 32'h00000000} /* (16, 0, 9) {real, imag} */,
  {32'h3e008830, 32'h00000000} /* (16, 0, 8) {real, imag} */,
  {32'hbe4be9e8, 32'h00000000} /* (16, 0, 7) {real, imag} */,
  {32'h3e8a886c, 32'h00000000} /* (16, 0, 6) {real, imag} */,
  {32'h3e84c07e, 32'h00000000} /* (16, 0, 5) {real, imag} */,
  {32'h3efc3b44, 32'h00000000} /* (16, 0, 4) {real, imag} */,
  {32'h3f06a742, 32'h00000000} /* (16, 0, 3) {real, imag} */,
  {32'hbf0cfac0, 32'h00000000} /* (16, 0, 2) {real, imag} */,
  {32'hbfb6545f, 32'h00000000} /* (16, 0, 1) {real, imag} */,
  {32'hbfb30e59, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h3e2729d2, 32'hbe6560e0} /* (15, 31, 31) {real, imag} */,
  {32'h3eb8c64d, 32'hbdc1ffc0} /* (15, 31, 30) {real, imag} */,
  {32'h3f0728d1, 32'h3ea432f8} /* (15, 31, 29) {real, imag} */,
  {32'h3e9e435a, 32'h3f58f5b0} /* (15, 31, 28) {real, imag} */,
  {32'h3e56299a, 32'h3e715ca0} /* (15, 31, 27) {real, imag} */,
  {32'h3e76cdea, 32'hbf045f84} /* (15, 31, 26) {real, imag} */,
  {32'h3e9001c4, 32'h3e487b30} /* (15, 31, 25) {real, imag} */,
  {32'h3d817120, 32'h3e3827c0} /* (15, 31, 24) {real, imag} */,
  {32'h3f1eb7be, 32'h3d8428c0} /* (15, 31, 23) {real, imag} */,
  {32'h3f12515b, 32'h3f34fee0} /* (15, 31, 22) {real, imag} */,
  {32'h3d9fb2fc, 32'h3ed5c568} /* (15, 31, 21) {real, imag} */,
  {32'hbdf72b80, 32'h3f344d26} /* (15, 31, 20) {real, imag} */,
  {32'h3e4c9abc, 32'h3d247d00} /* (15, 31, 19) {real, imag} */,
  {32'hbdf53020, 32'h3e29eef8} /* (15, 31, 18) {real, imag} */,
  {32'hbe549749, 32'h3f3489b8} /* (15, 31, 17) {real, imag} */,
  {32'hbf097ff7, 32'h3e08a460} /* (15, 31, 16) {real, imag} */,
  {32'hbd8ef9f8, 32'h3e952928} /* (15, 31, 15) {real, imag} */,
  {32'hbe04856c, 32'h3e6d51e0} /* (15, 31, 14) {real, imag} */,
  {32'hbed9903e, 32'h3f547a74} /* (15, 31, 13) {real, imag} */,
  {32'hbf03553e, 32'h3f34992a} /* (15, 31, 12) {real, imag} */,
  {32'hbec967c6, 32'h3e979d88} /* (15, 31, 11) {real, imag} */,
  {32'hbe3fdb49, 32'h3e2c71e0} /* (15, 31, 10) {real, imag} */,
  {32'hbd6b4e18, 32'h3ea8e704} /* (15, 31, 9) {real, imag} */,
  {32'h3f0bd69d, 32'h3f0e6edc} /* (15, 31, 8) {real, imag} */,
  {32'hbe705dc8, 32'hbf4a36d8} /* (15, 31, 7) {real, imag} */,
  {32'h3e0f58c4, 32'hbef41c50} /* (15, 31, 6) {real, imag} */,
  {32'h3f4ca65f, 32'hbe41cba0} /* (15, 31, 5) {real, imag} */,
  {32'h3f277a67, 32'h3e1e3650} /* (15, 31, 4) {real, imag} */,
  {32'h3f55db1a, 32'h3e6eefc0} /* (15, 31, 3) {real, imag} */,
  {32'h3dab4c4e, 32'h3d6d7800} /* (15, 31, 2) {real, imag} */,
  {32'h3d7e4940, 32'hbe20a700} /* (15, 31, 1) {real, imag} */,
  {32'h3ee38eea, 32'hbebe8e0c} /* (15, 31, 0) {real, imag} */,
  {32'h3e0f2c4c, 32'h3db82de0} /* (15, 30, 31) {real, imag} */,
  {32'h3dd0c530, 32'h3eb51c30} /* (15, 30, 30) {real, imag} */,
  {32'h3f67fa14, 32'h3f07bb10} /* (15, 30, 29) {real, imag} */,
  {32'h3f272664, 32'h3fab042c} /* (15, 30, 28) {real, imag} */,
  {32'h3f21859a, 32'h3f02818c} /* (15, 30, 27) {real, imag} */,
  {32'h3e0f952a, 32'hbe74f400} /* (15, 30, 26) {real, imag} */,
  {32'h3d868c1c, 32'h3ebfba70} /* (15, 30, 25) {real, imag} */,
  {32'h3dc7905a, 32'hbefa3d80} /* (15, 30, 24) {real, imag} */,
  {32'h3e960de4, 32'hbefaf560} /* (15, 30, 23) {real, imag} */,
  {32'h3f3f3e59, 32'h3f912a8c} /* (15, 30, 22) {real, imag} */,
  {32'h3e815bf4, 32'h3f2a9998} /* (15, 30, 21) {real, imag} */,
  {32'h3d8af1c6, 32'h3e644e80} /* (15, 30, 20) {real, imag} */,
  {32'h3f57c03a, 32'hbe70fc00} /* (15, 30, 19) {real, imag} */,
  {32'h3e93adf6, 32'hbd0cc600} /* (15, 30, 18) {real, imag} */,
  {32'hbec84ef6, 32'h3f5d0fa4} /* (15, 30, 17) {real, imag} */,
  {32'hbea8e087, 32'h3eca8880} /* (15, 30, 16) {real, imag} */,
  {32'h3d35b0f0, 32'h3e61f0e0} /* (15, 30, 15) {real, imag} */,
  {32'hbd24aac0, 32'hba6fa000} /* (15, 30, 14) {real, imag} */,
  {32'hbe9d7f14, 32'h3f3248dc} /* (15, 30, 13) {real, imag} */,
  {32'hbf443d0d, 32'h3f146c10} /* (15, 30, 12) {real, imag} */,
  {32'hbef2c3fe, 32'h3f1e36ae} /* (15, 30, 11) {real, imag} */,
  {32'h3d191760, 32'h3eeaa688} /* (15, 30, 10) {real, imag} */,
  {32'h3f08e918, 32'h3ec72cf8} /* (15, 30, 9) {real, imag} */,
  {32'h3eba66e0, 32'h3f7862c8} /* (15, 30, 8) {real, imag} */,
  {32'h3def15f0, 32'hbedc5298} /* (15, 30, 7) {real, imag} */,
  {32'h3f8f0353, 32'hbf311498} /* (15, 30, 6) {real, imag} */,
  {32'h3f8371c6, 32'hbe0e0ea0} /* (15, 30, 5) {real, imag} */,
  {32'h3f904a84, 32'hbe281060} /* (15, 30, 4) {real, imag} */,
  {32'h3f3f7bf1, 32'h3e91db58} /* (15, 30, 3) {real, imag} */,
  {32'hbf0e514c, 32'hbdb08500} /* (15, 30, 2) {real, imag} */,
  {32'hbeb723de, 32'h3c19c400} /* (15, 30, 1) {real, imag} */,
  {32'h3e65df52, 32'hbe929234} /* (15, 30, 0) {real, imag} */,
  {32'hbefd999e, 32'hbe5d1b00} /* (15, 29, 31) {real, imag} */,
  {32'hbce06500, 32'h3ed8c150} /* (15, 29, 30) {real, imag} */,
  {32'h3f06356a, 32'h3f47a050} /* (15, 29, 29) {real, imag} */,
  {32'h3eda9c28, 32'h3e88fa08} /* (15, 29, 28) {real, imag} */,
  {32'h3f1edba2, 32'h3eefbc18} /* (15, 29, 27) {real, imag} */,
  {32'h3d29f3f0, 32'h3ec8eed8} /* (15, 29, 26) {real, imag} */,
  {32'h3e6547c8, 32'hbcafaf80} /* (15, 29, 25) {real, imag} */,
  {32'hbe590700, 32'hbf04de30} /* (15, 29, 24) {real, imag} */,
  {32'hbbfcae00, 32'hbd5ba3c0} /* (15, 29, 23) {real, imag} */,
  {32'h3f6db1b6, 32'h3f1acc74} /* (15, 29, 22) {real, imag} */,
  {32'h3f68448c, 32'h3ed21590} /* (15, 29, 21) {real, imag} */,
  {32'h3f77b094, 32'h3e5b5cb0} /* (15, 29, 20) {real, imag} */,
  {32'h3f361796, 32'h3b6d2000} /* (15, 29, 19) {real, imag} */,
  {32'h3f9221c3, 32'h3e957190} /* (15, 29, 18) {real, imag} */,
  {32'h3ed7fd78, 32'h3f3ca5ac} /* (15, 29, 17) {real, imag} */,
  {32'hbdbe50d0, 32'h3f38dffc} /* (15, 29, 16) {real, imag} */,
  {32'hbf0a06b3, 32'h3f2db084} /* (15, 29, 15) {real, imag} */,
  {32'hbe598200, 32'h3c4a1c00} /* (15, 29, 14) {real, imag} */,
  {32'h3eb39750, 32'h3c4f3200} /* (15, 29, 13) {real, imag} */,
  {32'hbf5faf80, 32'h3e3d3d90} /* (15, 29, 12) {real, imag} */,
  {32'hbf756b3a, 32'h3e926730} /* (15, 29, 11) {real, imag} */,
  {32'hbec09660, 32'h3e532ea4} /* (15, 29, 10) {real, imag} */,
  {32'h3e9289a6, 32'h3da201a0} /* (15, 29, 9) {real, imag} */,
  {32'hbd881820, 32'h3f0b64c8} /* (15, 29, 8) {real, imag} */,
  {32'h3d9160b8, 32'h3eb2e260} /* (15, 29, 7) {real, imag} */,
  {32'h3f563f16, 32'h3d098700} /* (15, 29, 6) {real, imag} */,
  {32'h3f1b0b33, 32'hbd8f1420} /* (15, 29, 5) {real, imag} */,
  {32'h3f40ddda, 32'h3e3e63c0} /* (15, 29, 4) {real, imag} */,
  {32'h3eb1e108, 32'h3d8790a0} /* (15, 29, 3) {real, imag} */,
  {32'hbf052816, 32'hbf31a690} /* (15, 29, 2) {real, imag} */,
  {32'hbef5a36c, 32'h3e63f000} /* (15, 29, 1) {real, imag} */,
  {32'hbec177d8, 32'h3ec07840} /* (15, 29, 0) {real, imag} */,
  {32'hbedafbc8, 32'hbef1ae18} /* (15, 28, 31) {real, imag} */,
  {32'hbeb8b6b8, 32'h3f00aa08} /* (15, 28, 30) {real, imag} */,
  {32'hbc63a100, 32'h3f17cee8} /* (15, 28, 29) {real, imag} */,
  {32'h3cc143c0, 32'hbf2f12d8} /* (15, 28, 28) {real, imag} */,
  {32'h3f161107, 32'hbd946ae0} /* (15, 28, 27) {real, imag} */,
  {32'h3ed6e5b0, 32'h3f88929a} /* (15, 28, 26) {real, imag} */,
  {32'h3f7d58d4, 32'h3d2fc680} /* (15, 28, 25) {real, imag} */,
  {32'h3f4de884, 32'hbdc42100} /* (15, 28, 24) {real, imag} */,
  {32'h3f61bba2, 32'h3e8a2360} /* (15, 28, 23) {real, imag} */,
  {32'h3f825be6, 32'hbc400c00} /* (15, 28, 22) {real, imag} */,
  {32'h3f68fdf7, 32'h3ec65748} /* (15, 28, 21) {real, imag} */,
  {32'h3f8106d6, 32'h3f356e6c} /* (15, 28, 20) {real, imag} */,
  {32'h3f187358, 32'h3e8efb10} /* (15, 28, 19) {real, imag} */,
  {32'h3f559ea2, 32'h3ecca7b0} /* (15, 28, 18) {real, imag} */,
  {32'h3f318cfd, 32'h3f033eb0} /* (15, 28, 17) {real, imag} */,
  {32'h3e0cf18a, 32'h3eb8ddb0} /* (15, 28, 16) {real, imag} */,
  {32'hbf6fa6a0, 32'h3f0bc090} /* (15, 28, 15) {real, imag} */,
  {32'hbf2b96b0, 32'h3c87e500} /* (15, 28, 14) {real, imag} */,
  {32'hbdba5e30, 32'hbf158ff8} /* (15, 28, 13) {real, imag} */,
  {32'hbf44c7a3, 32'hbf413bac} /* (15, 28, 12) {real, imag} */,
  {32'hbee99cce, 32'hbf02e188} /* (15, 28, 11) {real, imag} */,
  {32'hbe2f4d28, 32'hbe5dff2c} /* (15, 28, 10) {real, imag} */,
  {32'hbeeae198, 32'h3d4a7b80} /* (15, 28, 9) {real, imag} */,
  {32'h3d60f220, 32'hbda927a0} /* (15, 28, 8) {real, imag} */,
  {32'h3e744b54, 32'hbe967848} /* (15, 28, 7) {real, imag} */,
  {32'h3e8e8730, 32'hbdc262c0} /* (15, 28, 6) {real, imag} */,
  {32'h3e92d20d, 32'h3e9e8e40} /* (15, 28, 5) {real, imag} */,
  {32'h3d158974, 32'h3f0432e8} /* (15, 28, 4) {real, imag} */,
  {32'h3e260478, 32'hbe992440} /* (15, 28, 3) {real, imag} */,
  {32'hbed32aec, 32'hbe8fd5a0} /* (15, 28, 2) {real, imag} */,
  {32'hbe565cc0, 32'h3eaa7260} /* (15, 28, 1) {real, imag} */,
  {32'hbe0d27a0, 32'h3e983850} /* (15, 28, 0) {real, imag} */,
  {32'hbe895b70, 32'h3dc4c740} /* (15, 27, 31) {real, imag} */,
  {32'hbf3b7648, 32'h3f0421b8} /* (15, 27, 30) {real, imag} */,
  {32'h3e3dae78, 32'h3ee4bb10} /* (15, 27, 29) {real, imag} */,
  {32'h3e5e6e8d, 32'hbebe0430} /* (15, 27, 28) {real, imag} */,
  {32'hbea0cb63, 32'hbdc0bc60} /* (15, 27, 27) {real, imag} */,
  {32'hbe2e9ffc, 32'h3f309328} /* (15, 27, 26) {real, imag} */,
  {32'h3f09cb34, 32'hbe3219c0} /* (15, 27, 25) {real, imag} */,
  {32'h3f10059c, 32'h3ebf2ef0} /* (15, 27, 24) {real, imag} */,
  {32'h3efa8c57, 32'h3f0e9df8} /* (15, 27, 23) {real, imag} */,
  {32'h3d9be758, 32'hbe15b730} /* (15, 27, 22) {real, imag} */,
  {32'hbaf7f600, 32'h3e3300d0} /* (15, 27, 21) {real, imag} */,
  {32'h3c9a4040, 32'h3f0dc0c4} /* (15, 27, 20) {real, imag} */,
  {32'h3d369f20, 32'hbe20aaa0} /* (15, 27, 19) {real, imag} */,
  {32'h3ee3bfb4, 32'hbe78f6e0} /* (15, 27, 18) {real, imag} */,
  {32'h3f52fe1a, 32'hbeea6fe0} /* (15, 27, 17) {real, imag} */,
  {32'h3e6df2f4, 32'hbe0edd00} /* (15, 27, 16) {real, imag} */,
  {32'hbf06652d, 32'h3ed48c60} /* (15, 27, 15) {real, imag} */,
  {32'hbebb64f0, 32'hbeeb20e0} /* (15, 27, 14) {real, imag} */,
  {32'hbf2dce68, 32'hbf79dbfc} /* (15, 27, 13) {real, imag} */,
  {32'hbec4dfa0, 32'hbf6cdbe8} /* (15, 27, 12) {real, imag} */,
  {32'h3f000e54, 32'hbf3edb3c} /* (15, 27, 11) {real, imag} */,
  {32'h3f046412, 32'hbeeefb6b} /* (15, 27, 10) {real, imag} */,
  {32'h3d163980, 32'hbe437440} /* (15, 27, 9) {real, imag} */,
  {32'h3b674600, 32'hbec77c60} /* (15, 27, 8) {real, imag} */,
  {32'h3e989780, 32'hbfa99a14} /* (15, 27, 7) {real, imag} */,
  {32'hbf0e414f, 32'hbf3ca7cc} /* (15, 27, 6) {real, imag} */,
  {32'h3e85cf70, 32'h3f14bcc8} /* (15, 27, 5) {real, imag} */,
  {32'h3f2b8004, 32'h3f441850} /* (15, 27, 4) {real, imag} */,
  {32'h3ec78b26, 32'hbe91d870} /* (15, 27, 3) {real, imag} */,
  {32'hbdea6d00, 32'hbeb39620} /* (15, 27, 2) {real, imag} */,
  {32'h3ea9d206, 32'h3f0e52d4} /* (15, 27, 1) {real, imag} */,
  {32'h3e56e200, 32'h3eced3b0} /* (15, 27, 0) {real, imag} */,
  {32'h3e4247c8, 32'hbde23bf0} /* (15, 26, 31) {real, imag} */,
  {32'h3d0c2950, 32'hbf165360} /* (15, 26, 30) {real, imag} */,
  {32'h3ee37918, 32'hbec47a60} /* (15, 26, 29) {real, imag} */,
  {32'hbdd2d570, 32'hbf3ee9c8} /* (15, 26, 28) {real, imag} */,
  {32'hbf2aaeef, 32'hbf509b50} /* (15, 26, 27) {real, imag} */,
  {32'hbe63d268, 32'hbeb464e0} /* (15, 26, 26) {real, imag} */,
  {32'hbda5f570, 32'hbe2512e0} /* (15, 26, 25) {real, imag} */,
  {32'hbe8d40a0, 32'hbe1ba600} /* (15, 26, 24) {real, imag} */,
  {32'hbbdc5780, 32'hbe93d978} /* (15, 26, 23) {real, imag} */,
  {32'h3cecbd50, 32'h3ddbd3e0} /* (15, 26, 22) {real, imag} */,
  {32'hbcec9b10, 32'hbd519180} /* (15, 26, 21) {real, imag} */,
  {32'hbed4d5e6, 32'hbec871ac} /* (15, 26, 20) {real, imag} */,
  {32'hbe495f0e, 32'hbed1ceb0} /* (15, 26, 19) {real, imag} */,
  {32'hbe585dce, 32'hbf3d3570} /* (15, 26, 18) {real, imag} */,
  {32'hbd8e001c, 32'hbf26a22c} /* (15, 26, 17) {real, imag} */,
  {32'h3e272afc, 32'hbc72ea00} /* (15, 26, 16) {real, imag} */,
  {32'h3f103402, 32'h3c739a00} /* (15, 26, 15) {real, imag} */,
  {32'h3f71d048, 32'hbebb55d8} /* (15, 26, 14) {real, imag} */,
  {32'h3f0a429c, 32'hbef57eb0} /* (15, 26, 13) {real, imag} */,
  {32'h3d2e3488, 32'hbf2123a0} /* (15, 26, 12) {real, imag} */,
  {32'h3e8912d2, 32'hbf0ff546} /* (15, 26, 11) {real, imag} */,
  {32'h3e97c778, 32'h3e69f5a0} /* (15, 26, 10) {real, imag} */,
  {32'h3c0c7f00, 32'h3e54ad40} /* (15, 26, 9) {real, imag} */,
  {32'hbe253c90, 32'hbe3b1840} /* (15, 26, 8) {real, imag} */,
  {32'h3c10d600, 32'hbeba9030} /* (15, 26, 7) {real, imag} */,
  {32'hbe89955c, 32'hbec500f0} /* (15, 26, 6) {real, imag} */,
  {32'h3f2f2dfe, 32'hbe0dde20} /* (15, 26, 5) {real, imag} */,
  {32'h3f43f30e, 32'h3e92b360} /* (15, 26, 4) {real, imag} */,
  {32'h3f04cef6, 32'h3cf53900} /* (15, 26, 3) {real, imag} */,
  {32'h3ef03bcd, 32'h3d9440c0} /* (15, 26, 2) {real, imag} */,
  {32'h3ebb7ad2, 32'h3ede22b0} /* (15, 26, 1) {real, imag} */,
  {32'h3ea7d35b, 32'hbcb2ed00} /* (15, 26, 0) {real, imag} */,
  {32'h3ed5c26b, 32'hbf277be0} /* (15, 25, 31) {real, imag} */,
  {32'h3c980d20, 32'hbf12c520} /* (15, 25, 30) {real, imag} */,
  {32'h3f230bcf, 32'hbee436c0} /* (15, 25, 29) {real, imag} */,
  {32'h3eaff3d0, 32'hbf010830} /* (15, 25, 28) {real, imag} */,
  {32'h3e219400, 32'hbf45ebf8} /* (15, 25, 27) {real, imag} */,
  {32'h3e6968d0, 32'hbee263c0} /* (15, 25, 26) {real, imag} */,
  {32'hbe7ef1e0, 32'hbecbd1c0} /* (15, 25, 25) {real, imag} */,
  {32'hbdd3b908, 32'hbeef26a0} /* (15, 25, 24) {real, imag} */,
  {32'h3e989a1e, 32'hbf5d2e78} /* (15, 25, 23) {real, imag} */,
  {32'hbeb89c12, 32'hbf1a694c} /* (15, 25, 22) {real, imag} */,
  {32'hbd3e1900, 32'hbf00d292} /* (15, 25, 21) {real, imag} */,
  {32'hbeb80a41, 32'hbf691274} /* (15, 25, 20) {real, imag} */,
  {32'hbe949454, 32'hbf4d5ec0} /* (15, 25, 19) {real, imag} */,
  {32'hbd8fbc88, 32'hbe849690} /* (15, 25, 18) {real, imag} */,
  {32'hbe2ded18, 32'hbf322e78} /* (15, 25, 17) {real, imag} */,
  {32'h3e9a2c34, 32'h3cb78d00} /* (15, 25, 16) {real, imag} */,
  {32'h3f30462e, 32'hbe4ff480} /* (15, 25, 15) {real, imag} */,
  {32'h3f16f9f0, 32'hbd030180} /* (15, 25, 14) {real, imag} */,
  {32'h3e8fd0e0, 32'h3f823964} /* (15, 25, 13) {real, imag} */,
  {32'hbe372cd0, 32'h3ea8aab0} /* (15, 25, 12) {real, imag} */,
  {32'h3eb413e2, 32'h3d9f9210} /* (15, 25, 11) {real, imag} */,
  {32'h3e777f80, 32'hbefec400} /* (15, 25, 10) {real, imag} */,
  {32'hbd74e410, 32'hbf110eb0} /* (15, 25, 9) {real, imag} */,
  {32'hbd49e300, 32'hbe0d9f80} /* (15, 25, 8) {real, imag} */,
  {32'hbe3ceb72, 32'h3db266e0} /* (15, 25, 7) {real, imag} */,
  {32'hbe820de8, 32'hbecb6988} /* (15, 25, 6) {real, imag} */,
  {32'h3e8d0b02, 32'hbf93ccb0} /* (15, 25, 5) {real, imag} */,
  {32'h3f17477c, 32'hbf49d0c0} /* (15, 25, 4) {real, imag} */,
  {32'h3e3621b0, 32'hbf66339c} /* (15, 25, 3) {real, imag} */,
  {32'hbf0951c0, 32'hbe964a50} /* (15, 25, 2) {real, imag} */,
  {32'hbd902e70, 32'h3d477b80} /* (15, 25, 1) {real, imag} */,
  {32'h3ec56c2c, 32'hbe7df340} /* (15, 25, 0) {real, imag} */,
  {32'h3ea70323, 32'hbf3e0582} /* (15, 24, 31) {real, imag} */,
  {32'h3df6a508, 32'hbf32b4a4} /* (15, 24, 30) {real, imag} */,
  {32'h3e5473d0, 32'h3de58300} /* (15, 24, 29) {real, imag} */,
  {32'h3db318f0, 32'h3f7b1b80} /* (15, 24, 28) {real, imag} */,
  {32'hbddbc938, 32'h3e9f0f98} /* (15, 24, 27) {real, imag} */,
  {32'hbed98478, 32'h3e9d0c38} /* (15, 24, 26) {real, imag} */,
  {32'h3cd95e90, 32'h3d3aae00} /* (15, 24, 25) {real, imag} */,
  {32'h3f4c5659, 32'hbee90c30} /* (15, 24, 24) {real, imag} */,
  {32'h3e0cb5e0, 32'hbf2c76a8} /* (15, 24, 23) {real, imag} */,
  {32'hbf464928, 32'hbec39c60} /* (15, 24, 22) {real, imag} */,
  {32'hbe4f88e0, 32'h3d1ce7c0} /* (15, 24, 21) {real, imag} */,
  {32'h3d844438, 32'hbef12950} /* (15, 24, 20) {real, imag} */,
  {32'h3d3bb7c0, 32'hbf499ba0} /* (15, 24, 19) {real, imag} */,
  {32'h3f557ad0, 32'h3f08b228} /* (15, 24, 18) {real, imag} */,
  {32'h3e8ec385, 32'hbd41bb80} /* (15, 24, 17) {real, imag} */,
  {32'h3e587408, 32'h3e48b540} /* (15, 24, 16) {real, imag} */,
  {32'h3d5cbdb0, 32'h3ebaedf8} /* (15, 24, 15) {real, imag} */,
  {32'hbec98bd6, 32'h3f2d42b0} /* (15, 24, 14) {real, imag} */,
  {32'hbe89fdf0, 32'h3fee57f4} /* (15, 24, 13) {real, imag} */,
  {32'hbe0272d4, 32'h3f957d7e} /* (15, 24, 12) {real, imag} */,
  {32'h3e0b6838, 32'hbe602530} /* (15, 24, 11) {real, imag} */,
  {32'h3e21f524, 32'hbf7bb7c4} /* (15, 24, 10) {real, imag} */,
  {32'h3d8f6cc8, 32'hbf820b34} /* (15, 24, 9) {real, imag} */,
  {32'h3e543cb0, 32'h3e6c7a00} /* (15, 24, 8) {real, imag} */,
  {32'hbe602a48, 32'hbe1bc140} /* (15, 24, 7) {real, imag} */,
  {32'hbf30c3d2, 32'hbe98baf8} /* (15, 24, 6) {real, imag} */,
  {32'h3daceb58, 32'hbf34b7e0} /* (15, 24, 5) {real, imag} */,
  {32'h3f04aca7, 32'hbf031ef0} /* (15, 24, 4) {real, imag} */,
  {32'h3f17f46b, 32'hbecc9640} /* (15, 24, 3) {real, imag} */,
  {32'hbe864dc0, 32'hbda9b540} /* (15, 24, 2) {real, imag} */,
  {32'hbf8633e8, 32'hbef12610} /* (15, 24, 1) {real, imag} */,
  {32'hbe710bc0, 32'h3d1c9d00} /* (15, 24, 0) {real, imag} */,
  {32'h3e899e02, 32'hbf36c6d4} /* (15, 23, 31) {real, imag} */,
  {32'hbd8533bc, 32'hbf203658} /* (15, 23, 30) {real, imag} */,
  {32'hbecd1fa2, 32'hbc107400} /* (15, 23, 29) {real, imag} */,
  {32'hbda21180, 32'h3e638540} /* (15, 23, 28) {real, imag} */,
  {32'h3db23960, 32'h3e2d2d10} /* (15, 23, 27) {real, imag} */,
  {32'hbe82ed72, 32'h3e4c5780} /* (15, 23, 26) {real, imag} */,
  {32'hbdf101d0, 32'hbe1188d0} /* (15, 23, 25) {real, imag} */,
  {32'h3f173f3c, 32'hbed636f8} /* (15, 23, 24) {real, imag} */,
  {32'hbf015880, 32'hbefbfb80} /* (15, 23, 23) {real, imag} */,
  {32'hbf78414a, 32'h3e01b640} /* (15, 23, 22) {real, imag} */,
  {32'h3ddddf90, 32'hbd0c9b40} /* (15, 23, 21) {real, imag} */,
  {32'h3e80069e, 32'h3d9be240} /* (15, 23, 20) {real, imag} */,
  {32'h3f0410f1, 32'hbe538680} /* (15, 23, 19) {real, imag} */,
  {32'h3fd75c33, 32'h3f0dfec8} /* (15, 23, 18) {real, imag} */,
  {32'h3f2478e7, 32'h3f60d0d0} /* (15, 23, 17) {real, imag} */,
  {32'hbf0814f2, 32'h3f882768} /* (15, 23, 16) {real, imag} */,
  {32'hbefcf591, 32'h3f54f298} /* (15, 23, 15) {real, imag} */,
  {32'hbdb69af0, 32'h3e09d090} /* (15, 23, 14) {real, imag} */,
  {32'hbeac34d6, 32'h3d423580} /* (15, 23, 13) {real, imag} */,
  {32'hbf2d607a, 32'hbd835d80} /* (15, 23, 12) {real, imag} */,
  {32'hbec8e740, 32'hbe10e980} /* (15, 23, 11) {real, imag} */,
  {32'hbe3f7730, 32'hbeb306c0} /* (15, 23, 10) {real, imag} */,
  {32'hbe83612a, 32'hbe9bc880} /* (15, 23, 9) {real, imag} */,
  {32'h3e603ab0, 32'hbd871e80} /* (15, 23, 8) {real, imag} */,
  {32'h3e250100, 32'h3df9c180} /* (15, 23, 7) {real, imag} */,
  {32'hbf5be1c2, 32'hbe1f0000} /* (15, 23, 6) {real, imag} */,
  {32'hbe5cb710, 32'hbefb8e80} /* (15, 23, 5) {real, imag} */,
  {32'hbdd3c790, 32'hbeedadc0} /* (15, 23, 4) {real, imag} */,
  {32'h3e8108a4, 32'h3edb9d78} /* (15, 23, 3) {real, imag} */,
  {32'hbb47c000, 32'h3f51faf4} /* (15, 23, 2) {real, imag} */,
  {32'hbf4a8429, 32'hbe1fda90} /* (15, 23, 1) {real, imag} */,
  {32'hbeff275d, 32'hbeb5f548} /* (15, 23, 0) {real, imag} */,
  {32'h3f0e032a, 32'hbef1cbbc} /* (15, 22, 31) {real, imag} */,
  {32'h3f0a515c, 32'hbf61a978} /* (15, 22, 30) {real, imag} */,
  {32'h3f1f9f60, 32'hbec3cd70} /* (15, 22, 29) {real, imag} */,
  {32'h3f9b4db9, 32'h3ce4fb00} /* (15, 22, 28) {real, imag} */,
  {32'h3f4180ea, 32'h3f1d7440} /* (15, 22, 27) {real, imag} */,
  {32'h3ea09522, 32'h3f555890} /* (15, 22, 26) {real, imag} */,
  {32'h3e08195a, 32'h3e6553e0} /* (15, 22, 25) {real, imag} */,
  {32'h3e56edce, 32'hbe122500} /* (15, 22, 24) {real, imag} */,
  {32'hbf3f2342, 32'hbdb35f80} /* (15, 22, 23) {real, imag} */,
  {32'hbf6e4dd6, 32'hbce5b500} /* (15, 22, 22) {real, imag} */,
  {32'hbea8ddfc, 32'hbe8db420} /* (15, 22, 21) {real, imag} */,
  {32'h3dd55288, 32'h3e562a00} /* (15, 22, 20) {real, imag} */,
  {32'hbda7d694, 32'h3e252e00} /* (15, 22, 19) {real, imag} */,
  {32'h3efa7542, 32'h3e9bdd90} /* (15, 22, 18) {real, imag} */,
  {32'hbe0a372e, 32'h3e289680} /* (15, 22, 17) {real, imag} */,
  {32'hbf7de92d, 32'h3f592440} /* (15, 22, 16) {real, imag} */,
  {32'hbf15b57e, 32'h3f0eb62c} /* (15, 22, 15) {real, imag} */,
  {32'h3e1bcd3e, 32'hbee63a40} /* (15, 22, 14) {real, imag} */,
  {32'h3ec60a53, 32'hbf5cef78} /* (15, 22, 13) {real, imag} */,
  {32'h3de24e08, 32'hbf6c14b0} /* (15, 22, 12) {real, imag} */,
  {32'hbe200580, 32'hbee57640} /* (15, 22, 11) {real, imag} */,
  {32'hbf1b6860, 32'hbd979b70} /* (15, 22, 10) {real, imag} */,
  {32'hbe1632a0, 32'h3cce9100} /* (15, 22, 9) {real, imag} */,
  {32'hbde60088, 32'hbf41da98} /* (15, 22, 8) {real, imag} */,
  {32'h3ebb5610, 32'hbce2d200} /* (15, 22, 7) {real, imag} */,
  {32'h3e601474, 32'h3e98ccf8} /* (15, 22, 6) {real, imag} */,
  {32'h3ca2c980, 32'hbe930ef0} /* (15, 22, 5) {real, imag} */,
  {32'hbe11bcd0, 32'hbf6c00f8} /* (15, 22, 4) {real, imag} */,
  {32'hbe8b82fc, 32'hbe050840} /* (15, 22, 3) {real, imag} */,
  {32'hbf67b6a8, 32'h3f03b4d0} /* (15, 22, 2) {real, imag} */,
  {32'hbf4d96ce, 32'h3e2c83c0} /* (15, 22, 1) {real, imag} */,
  {32'hbf3df622, 32'hbe84c0c0} /* (15, 22, 0) {real, imag} */,
  {32'h3e667c84, 32'hbf05cfaa} /* (15, 21, 31) {real, imag} */,
  {32'h3e99a12c, 32'hbeca1040} /* (15, 21, 30) {real, imag} */,
  {32'h3ee1d994, 32'hbe612ec0} /* (15, 21, 29) {real, imag} */,
  {32'h3f8d0c00, 32'h3d56adc0} /* (15, 21, 28) {real, imag} */,
  {32'h3f4bef1d, 32'h3ecd3d80} /* (15, 21, 27) {real, imag} */,
  {32'h3f13c1fc, 32'h3ecdff60} /* (15, 21, 26) {real, imag} */,
  {32'h3f39f995, 32'h3f0426e0} /* (15, 21, 25) {real, imag} */,
  {32'h3ef49410, 32'hba1ed000} /* (15, 21, 24) {real, imag} */,
  {32'hbe81449e, 32'hbd098fc0} /* (15, 21, 23) {real, imag} */,
  {32'hbf3133c6, 32'hbcf27300} /* (15, 21, 22) {real, imag} */,
  {32'hbddcd488, 32'h3c473800} /* (15, 21, 21) {real, imag} */,
  {32'h3eb643c4, 32'h3ed7edf4} /* (15, 21, 20) {real, imag} */,
  {32'hbe3466b1, 32'h3d115080} /* (15, 21, 19) {real, imag} */,
  {32'hbd7c3ad0, 32'h3f3c74c0} /* (15, 21, 18) {real, imag} */,
  {32'hbe19d85e, 32'h3ee5d860} /* (15, 21, 17) {real, imag} */,
  {32'hbea5215e, 32'hbf044cb5} /* (15, 21, 16) {real, imag} */,
  {32'hbec76588, 32'h3d796600} /* (15, 21, 15) {real, imag} */,
  {32'hbe5e21c4, 32'hbdb375c0} /* (15, 21, 14) {real, imag} */,
  {32'h3ea01c3e, 32'hbeeed7d0} /* (15, 21, 13) {real, imag} */,
  {32'h3e2621c9, 32'hbee52190} /* (15, 21, 12) {real, imag} */,
  {32'hbcbc71e0, 32'h3e008eb0} /* (15, 21, 11) {real, imag} */,
  {32'hbecb15d0, 32'h3eb50d90} /* (15, 21, 10) {real, imag} */,
  {32'h3dc6162c, 32'h3d0be900} /* (15, 21, 9) {real, imag} */,
  {32'hbe9e1f7e, 32'hbe8101a8} /* (15, 21, 8) {real, imag} */,
  {32'hbd286480, 32'hbf0dca70} /* (15, 21, 7) {real, imag} */,
  {32'h3f94b570, 32'h3ef1c932} /* (15, 21, 6) {real, imag} */,
  {32'h3f98c73b, 32'hbdee8700} /* (15, 21, 5) {real, imag} */,
  {32'h3f3faebc, 32'hbf05de3c} /* (15, 21, 4) {real, imag} */,
  {32'hbeb42b22, 32'hbe771e10} /* (15, 21, 3) {real, imag} */,
  {32'hbf19fe21, 32'hbeda65d4} /* (15, 21, 2) {real, imag} */,
  {32'hbec323a0, 32'hbf390b86} /* (15, 21, 1) {real, imag} */,
  {32'hbe32d572, 32'hbf452ead} /* (15, 21, 0) {real, imag} */,
  {32'h3deb4780, 32'hbf1f8fe4} /* (15, 20, 31) {real, imag} */,
  {32'h3dcbcc80, 32'hbee422b0} /* (15, 20, 30) {real, imag} */,
  {32'h3eaad2f4, 32'h3dc3e8e0} /* (15, 20, 29) {real, imag} */,
  {32'h3fb9d3d4, 32'h3e3080d8} /* (15, 20, 28) {real, imag} */,
  {32'h3f36022a, 32'h3e879e80} /* (15, 20, 27) {real, imag} */,
  {32'h3eec670b, 32'h3dadeca0} /* (15, 20, 26) {real, imag} */,
  {32'h3ed61930, 32'h3e7bd888} /* (15, 20, 25) {real, imag} */,
  {32'h3dd51cbc, 32'h3e996e80} /* (15, 20, 24) {real, imag} */,
  {32'hbdfe7e10, 32'hbea78870} /* (15, 20, 23) {real, imag} */,
  {32'hbeaad1b2, 32'hbefa1530} /* (15, 20, 22) {real, imag} */,
  {32'hbe572950, 32'h3ea02f1c} /* (15, 20, 21) {real, imag} */,
  {32'h3e2cb86e, 32'h3f45f600} /* (15, 20, 20) {real, imag} */,
  {32'h3e9a3320, 32'h3f1c3f88} /* (15, 20, 19) {real, imag} */,
  {32'hbd20f2da, 32'h3f84effc} /* (15, 20, 18) {real, imag} */,
  {32'hbe57d9fc, 32'h3f423070} /* (15, 20, 17) {real, imag} */,
  {32'h3f55bb40, 32'hbe6af500} /* (15, 20, 16) {real, imag} */,
  {32'h3eae8970, 32'h3d8a7780} /* (15, 20, 15) {real, imag} */,
  {32'hbf2299ce, 32'h3e99f5b8} /* (15, 20, 14) {real, imag} */,
  {32'hbe00c7b0, 32'h3f0d6648} /* (15, 20, 13) {real, imag} */,
  {32'h3f829efa, 32'hbd12b300} /* (15, 20, 12) {real, imag} */,
  {32'h3f44e65f, 32'hbeb913f0} /* (15, 20, 11) {real, imag} */,
  {32'h3c316f80, 32'hbe449830} /* (15, 20, 10) {real, imag} */,
  {32'h3ebc10a0, 32'hbe067210} /* (15, 20, 9) {real, imag} */,
  {32'h3e02f520, 32'h3ece0520} /* (15, 20, 8) {real, imag} */,
  {32'h3dc61494, 32'hbefe83b8} /* (15, 20, 7) {real, imag} */,
  {32'h3f61fc93, 32'h3f2678d0} /* (15, 20, 6) {real, imag} */,
  {32'h3e376a9b, 32'hbdc86cf0} /* (15, 20, 5) {real, imag} */,
  {32'hbe8a824a, 32'hbe65f980} /* (15, 20, 4) {real, imag} */,
  {32'hbdb39310, 32'hbe655e80} /* (15, 20, 3) {real, imag} */,
  {32'hbf0e7799, 32'hbeedd648} /* (15, 20, 2) {real, imag} */,
  {32'hbf0f2a92, 32'hbea34bb0} /* (15, 20, 1) {real, imag} */,
  {32'h3d302300, 32'hbecf9848} /* (15, 20, 0) {real, imag} */,
  {32'h3ec24ad3, 32'hbdee9460} /* (15, 19, 31) {real, imag} */,
  {32'h3ee5df54, 32'h3eccfe40} /* (15, 19, 30) {real, imag} */,
  {32'h3e9943ea, 32'h3efc5d30} /* (15, 19, 29) {real, imag} */,
  {32'h3f49f880, 32'h3e5b6340} /* (15, 19, 28) {real, imag} */,
  {32'h3ea3c9a0, 32'h3e3ddf80} /* (15, 19, 27) {real, imag} */,
  {32'h3ec6efb0, 32'hbe3150e0} /* (15, 19, 26) {real, imag} */,
  {32'h3e8dc3e9, 32'hbde52900} /* (15, 19, 25) {real, imag} */,
  {32'hbe031c60, 32'h3e24a900} /* (15, 19, 24) {real, imag} */,
  {32'hbefd43d0, 32'hbe82aac0} /* (15, 19, 23) {real, imag} */,
  {32'hbf4c90fa, 32'hbdcb0380} /* (15, 19, 22) {real, imag} */,
  {32'hbf06332d, 32'h3efc9718} /* (15, 19, 21) {real, imag} */,
  {32'h3e82505a, 32'h3f8e04e0} /* (15, 19, 20) {real, imag} */,
  {32'hbdc0b020, 32'h3f032b20} /* (15, 19, 19) {real, imag} */,
  {32'hbf46f115, 32'h3f40d580} /* (15, 19, 18) {real, imag} */,
  {32'hbe803b4b, 32'h3f449948} /* (15, 19, 17) {real, imag} */,
  {32'h3f6c6916, 32'hbe9c3f10} /* (15, 19, 16) {real, imag} */,
  {32'h3f3618cc, 32'hbe12c340} /* (15, 19, 15) {real, imag} */,
  {32'h3eb0e035, 32'h3eda33f0} /* (15, 19, 14) {real, imag} */,
  {32'h3f0d3a36, 32'h3f866590} /* (15, 19, 13) {real, imag} */,
  {32'h3f5102ce, 32'h3f3be278} /* (15, 19, 12) {real, imag} */,
  {32'h3ee182a4, 32'hbee8ec20} /* (15, 19, 11) {real, imag} */,
  {32'hbe576e40, 32'hbf0c2cd8} /* (15, 19, 10) {real, imag} */,
  {32'hbe676154, 32'hbec96940} /* (15, 19, 9) {real, imag} */,
  {32'h3d3aee40, 32'h3e9dbb90} /* (15, 19, 8) {real, imag} */,
  {32'hbe4fade8, 32'h3e33f2b0} /* (15, 19, 7) {real, imag} */,
  {32'hbe0de454, 32'h3f3a8168} /* (15, 19, 6) {real, imag} */,
  {32'hbeb33450, 32'h3e46b910} /* (15, 19, 5) {real, imag} */,
  {32'hbf3029e0, 32'h3ea56ca0} /* (15, 19, 4) {real, imag} */,
  {32'hbe234928, 32'h3e8cd918} /* (15, 19, 3) {real, imag} */,
  {32'h3c86f180, 32'hbe15bba0} /* (15, 19, 2) {real, imag} */,
  {32'hbf03dfe8, 32'hbeccfb10} /* (15, 19, 1) {real, imag} */,
  {32'h3ca99ec0, 32'hbc387d00} /* (15, 19, 0) {real, imag} */,
  {32'hbe585688, 32'hbef6e8c0} /* (15, 18, 31) {real, imag} */,
  {32'hbe98e618, 32'h3e649a40} /* (15, 18, 30) {real, imag} */,
  {32'h3ef02270, 32'h3e6d1f00} /* (15, 18, 29) {real, imag} */,
  {32'h3ead834c, 32'hbeb0bf30} /* (15, 18, 28) {real, imag} */,
  {32'hbeb9e1ca, 32'h3dcfc440} /* (15, 18, 27) {real, imag} */,
  {32'hbef49ce2, 32'hbf0b19c0} /* (15, 18, 26) {real, imag} */,
  {32'h3ea3cc1c, 32'hbe4db800} /* (15, 18, 25) {real, imag} */,
  {32'hb89f0000, 32'hbe364f40} /* (15, 18, 24) {real, imag} */,
  {32'hbf32c25e, 32'h3eed2c40} /* (15, 18, 23) {real, imag} */,
  {32'hbf85fd9e, 32'h3e994290} /* (15, 18, 22) {real, imag} */,
  {32'hbed4d1e4, 32'hbe18e420} /* (15, 18, 21) {real, imag} */,
  {32'h3dd0ba88, 32'h3ea88010} /* (15, 18, 20) {real, imag} */,
  {32'hbea4e25c, 32'hbd1c9700} /* (15, 18, 19) {real, imag} */,
  {32'hbf05c5d6, 32'h3f6c4900} /* (15, 18, 18) {real, imag} */,
  {32'h3e84d8a8, 32'h3f203090} /* (15, 18, 17) {real, imag} */,
  {32'h3f02250c, 32'hbc32dc00} /* (15, 18, 16) {real, imag} */,
  {32'h3ecd3dcc, 32'h3e9f7720} /* (15, 18, 15) {real, imag} */,
  {32'h3f60be9c, 32'h3f39a82c} /* (15, 18, 14) {real, imag} */,
  {32'h3f556edc, 32'h3f434010} /* (15, 18, 13) {real, imag} */,
  {32'h3ee6a672, 32'h3f8ae180} /* (15, 18, 12) {real, imag} */,
  {32'h3d018410, 32'hbe931f30} /* (15, 18, 11) {real, imag} */,
  {32'h3e24ca38, 32'hbf58d9a4} /* (15, 18, 10) {real, imag} */,
  {32'hbed6a4d8, 32'hbe434e70} /* (15, 18, 9) {real, imag} */,
  {32'hbf994536, 32'hbced1a00} /* (15, 18, 8) {real, imag} */,
  {32'hbf8b4c2c, 32'h3ea18540} /* (15, 18, 7) {real, imag} */,
  {32'hbd989b68, 32'h3f103ec8} /* (15, 18, 6) {real, imag} */,
  {32'h3e842008, 32'h3f483ce8} /* (15, 18, 5) {real, imag} */,
  {32'h3e434a48, 32'h3f159e34} /* (15, 18, 4) {real, imag} */,
  {32'h3ea81e99, 32'h3c289000} /* (15, 18, 3) {real, imag} */,
  {32'h3f2474bb, 32'h3f18e3d8} /* (15, 18, 2) {real, imag} */,
  {32'h3ecfe668, 32'hbecb5650} /* (15, 18, 1) {real, imag} */,
  {32'hbe7071c0, 32'hbf2e1b14} /* (15, 18, 0) {real, imag} */,
  {32'hbf991a3b, 32'hbededa80} /* (15, 17, 31) {real, imag} */,
  {32'hbf56cb8e, 32'hbe19da40} /* (15, 17, 30) {real, imag} */,
  {32'h3d908810, 32'h3e1c3e20} /* (15, 17, 29) {real, imag} */,
  {32'h3e03125c, 32'h3bf0b800} /* (15, 17, 28) {real, imag} */,
  {32'hbe9ea8ec, 32'h3ea225a0} /* (15, 17, 27) {real, imag} */,
  {32'hbf5dca6a, 32'hbd7c9780} /* (15, 17, 26) {real, imag} */,
  {32'hbf7b3c03, 32'hbde1edc0} /* (15, 17, 25) {real, imag} */,
  {32'hbf49c924, 32'h3d546180} /* (15, 17, 24) {real, imag} */,
  {32'hbf1ae4f5, 32'h3eab9890} /* (15, 17, 23) {real, imag} */,
  {32'hbf33af62, 32'h3e995cd8} /* (15, 17, 22) {real, imag} */,
  {32'h3e7cffd0, 32'h3dde8428} /* (15, 17, 21) {real, imag} */,
  {32'h3f10e092, 32'hbe00ecf0} /* (15, 17, 20) {real, imag} */,
  {32'h3c3f2980, 32'hbde82580} /* (15, 17, 19) {real, imag} */,
  {32'hbe02638c, 32'h3ed710e0} /* (15, 17, 18) {real, imag} */,
  {32'hbee6ea7c, 32'h3e058e40} /* (15, 17, 17) {real, imag} */,
  {32'h3cd65d00, 32'h3ee49a30} /* (15, 17, 16) {real, imag} */,
  {32'h3f05b012, 32'h3ee96dc0} /* (15, 17, 15) {real, imag} */,
  {32'h3f396aa0, 32'h3e8df5c0} /* (15, 17, 14) {real, imag} */,
  {32'h3ed65e0c, 32'h3f0a80a8} /* (15, 17, 13) {real, imag} */,
  {32'h3f5a99da, 32'h3ed3f540} /* (15, 17, 12) {real, imag} */,
  {32'h3f48a3ab, 32'hbf7b5258} /* (15, 17, 11) {real, imag} */,
  {32'h3ee95d7c, 32'hbf9a733c} /* (15, 17, 10) {real, imag} */,
  {32'hbf747fd0, 32'hbf63c568} /* (15, 17, 9) {real, imag} */,
  {32'hbf536bd4, 32'h3d639500} /* (15, 17, 8) {real, imag} */,
  {32'hbe48ecb8, 32'h3e892b50} /* (15, 17, 7) {real, imag} */,
  {32'hbe9b0300, 32'h3e5e3080} /* (15, 17, 6) {real, imag} */,
  {32'h3e87e754, 32'h3f42b364} /* (15, 17, 5) {real, imag} */,
  {32'hbe97dd27, 32'hbc01a400} /* (15, 17, 4) {real, imag} */,
  {32'hbe2c469c, 32'h3ef8c3c0} /* (15, 17, 3) {real, imag} */,
  {32'h3f169960, 32'h3f2c4060} /* (15, 17, 2) {real, imag} */,
  {32'h3c40ca80, 32'hbf3d72a0} /* (15, 17, 1) {real, imag} */,
  {32'hbf3b355a, 32'hbf8b29d4} /* (15, 17, 0) {real, imag} */,
  {32'hbf1c4f0a, 32'hbe8c5598} /* (15, 16, 31) {real, imag} */,
  {32'hbf271314, 32'hbe7878e0} /* (15, 16, 30) {real, imag} */,
  {32'hbf0480f0, 32'h3dffaec0} /* (15, 16, 29) {real, imag} */,
  {32'hbec13040, 32'h3f3b2740} /* (15, 16, 28) {real, imag} */,
  {32'hbf0ce2aa, 32'h3eb64670} /* (15, 16, 27) {real, imag} */,
  {32'hbf41b0f7, 32'h3f3989c4} /* (15, 16, 26) {real, imag} */,
  {32'hbf7f9caa, 32'h3f46c52c} /* (15, 16, 25) {real, imag} */,
  {32'hbf358e14, 32'hbdf3cb40} /* (15, 16, 24) {real, imag} */,
  {32'h3e29cf66, 32'hbeb7f0c0} /* (15, 16, 23) {real, imag} */,
  {32'hbe800ae8, 32'h3de53d80} /* (15, 16, 22) {real, imag} */,
  {32'h3cf54900, 32'h3ec86a01} /* (15, 16, 21) {real, imag} */,
  {32'h3eb4b6c4, 32'h3ef96fb0} /* (15, 16, 20) {real, imag} */,
  {32'h3e535278, 32'h3f120b28} /* (15, 16, 19) {real, imag} */,
  {32'h3f150395, 32'h3da37500} /* (15, 16, 18) {real, imag} */,
  {32'h3f3b32be, 32'hbe101aa0} /* (15, 16, 17) {real, imag} */,
  {32'h3f8def93, 32'h3f187c88} /* (15, 16, 16) {real, imag} */,
  {32'h3f1f41c8, 32'h3f110578} /* (15, 16, 15) {real, imag} */,
  {32'hbda93400, 32'h3eddbe40} /* (15, 16, 14) {real, imag} */,
  {32'hbf1d5536, 32'h3f21a3b8} /* (15, 16, 13) {real, imag} */,
  {32'h3f12e45f, 32'hbdf41680} /* (15, 16, 12) {real, imag} */,
  {32'h3ef95870, 32'hbf71b198} /* (15, 16, 11) {real, imag} */,
  {32'h3f02d2ae, 32'hbf51d1ea} /* (15, 16, 10) {real, imag} */,
  {32'hbef02bbf, 32'hbf065c28} /* (15, 16, 9) {real, imag} */,
  {32'hbf1cd86e, 32'h3dc683c0} /* (15, 16, 8) {real, imag} */,
  {32'h3aff0800, 32'hbd43ff40} /* (15, 16, 7) {real, imag} */,
  {32'hbd1694a0, 32'h3d43bb00} /* (15, 16, 6) {real, imag} */,
  {32'hbf0c0dd9, 32'h3e347c40} /* (15, 16, 5) {real, imag} */,
  {32'hbf41bf44, 32'hbf1247f0} /* (15, 16, 4) {real, imag} */,
  {32'hbf2033d2, 32'h3e425d40} /* (15, 16, 3) {real, imag} */,
  {32'hbee01220, 32'h3e90b120} /* (15, 16, 2) {real, imag} */,
  {32'hbf5eb25c, 32'hbf9f0a8c} /* (15, 16, 1) {real, imag} */,
  {32'hbf079b7a, 32'hbfa00a64} /* (15, 16, 0) {real, imag} */,
  {32'h3d6abdf0, 32'hbdda6880} /* (15, 15, 31) {real, imag} */,
  {32'hbe6068d0, 32'h3efe72c0} /* (15, 15, 30) {real, imag} */,
  {32'hbf16d3f4, 32'h3f7aa940} /* (15, 15, 29) {real, imag} */,
  {32'hbdeaaab4, 32'h3f6e70f0} /* (15, 15, 28) {real, imag} */,
  {32'hbee05e0b, 32'h3f82b0e4} /* (15, 15, 27) {real, imag} */,
  {32'hbecfbc63, 32'h3f8d9474} /* (15, 15, 26) {real, imag} */,
  {32'hbe9fb010, 32'h3f9844b4} /* (15, 15, 25) {real, imag} */,
  {32'h3e39c98c, 32'hbe619760} /* (15, 15, 24) {real, imag} */,
  {32'h3f40d659, 32'hbd8ee600} /* (15, 15, 23) {real, imag} */,
  {32'hbeb2e665, 32'h3e917f88} /* (15, 15, 22) {real, imag} */,
  {32'hbecff048, 32'h3df15960} /* (15, 15, 21) {real, imag} */,
  {32'h3bbde500, 32'h3ea4ed60} /* (15, 15, 20) {real, imag} */,
  {32'h3f4aba8c, 32'h3f2315a8} /* (15, 15, 19) {real, imag} */,
  {32'h3f806242, 32'hbdd4d180} /* (15, 15, 18) {real, imag} */,
  {32'h3f6b19b8, 32'hbcaa2100} /* (15, 15, 17) {real, imag} */,
  {32'h3fabdc7c, 32'h3e2df4a0} /* (15, 15, 16) {real, imag} */,
  {32'h3f29303c, 32'h3e6f6dc0} /* (15, 15, 15) {real, imag} */,
  {32'hbbc47000, 32'h3f39e6cc} /* (15, 15, 14) {real, imag} */,
  {32'h3e5dec06, 32'h3c3a1e00} /* (15, 15, 13) {real, imag} */,
  {32'h3e957c18, 32'hbe4687e0} /* (15, 15, 12) {real, imag} */,
  {32'h3d784aa0, 32'h3e4bc580} /* (15, 15, 11) {real, imag} */,
  {32'h3f19fd44, 32'h3efd94b8} /* (15, 15, 10) {real, imag} */,
  {32'hbebc97ac, 32'h3f1729c0} /* (15, 15, 9) {real, imag} */,
  {32'hbed19120, 32'h3f0248c0} /* (15, 15, 8) {real, imag} */,
  {32'hbe137368, 32'hbf028a70} /* (15, 15, 7) {real, imag} */,
  {32'hbdd2b5c8, 32'hbf31804c} /* (15, 15, 6) {real, imag} */,
  {32'hbf18d484, 32'hbc976900} /* (15, 15, 5) {real, imag} */,
  {32'hbf202358, 32'h3eb89ab0} /* (15, 15, 4) {real, imag} */,
  {32'hbf62f4dc, 32'hbdd520c0} /* (15, 15, 3) {real, imag} */,
  {32'hbf03cccf, 32'hbe5d9b20} /* (15, 15, 2) {real, imag} */,
  {32'hbf455eb1, 32'hbe939e80} /* (15, 15, 1) {real, imag} */,
  {32'hbefb0cb4, 32'hbec79080} /* (15, 15, 0) {real, imag} */,
  {32'h3ea81773, 32'h3dc52100} /* (15, 14, 31) {real, imag} */,
  {32'h3dac2130, 32'h3f127798} /* (15, 14, 30) {real, imag} */,
  {32'hbd2a2f74, 32'h3faac034} /* (15, 14, 29) {real, imag} */,
  {32'h3f29dde0, 32'h3f5a72d8} /* (15, 14, 28) {real, imag} */,
  {32'h3e20e598, 32'h3f43c810} /* (15, 14, 27) {real, imag} */,
  {32'hbf7f4484, 32'h3dfdd900} /* (15, 14, 26) {real, imag} */,
  {32'hbf5736f0, 32'h3f29cd38} /* (15, 14, 25) {real, imag} */,
  {32'hbeb1e8c8, 32'h3d781080} /* (15, 14, 24) {real, imag} */,
  {32'hbf109d9a, 32'hbf644c60} /* (15, 14, 23) {real, imag} */,
  {32'hbf1faa0c, 32'hbf93844c} /* (15, 14, 22) {real, imag} */,
  {32'hbeceb720, 32'hbe7a1d10} /* (15, 14, 21) {real, imag} */,
  {32'h3eee9d7c, 32'h3eaac890} /* (15, 14, 20) {real, imag} */,
  {32'h3f834bba, 32'hbdca6440} /* (15, 14, 19) {real, imag} */,
  {32'h3fa039f8, 32'h3e344840} /* (15, 14, 18) {real, imag} */,
  {32'h3ec716d8, 32'h3f2ba2e8} /* (15, 14, 17) {real, imag} */,
  {32'h3ed4e47c, 32'h3d900680} /* (15, 14, 16) {real, imag} */,
  {32'h3efbcbe6, 32'hbeb72df0} /* (15, 14, 15) {real, imag} */,
  {32'h3ee76d80, 32'hbe3eb3a0} /* (15, 14, 14) {real, imag} */,
  {32'h3fb64e10, 32'hbf0d3188} /* (15, 14, 13) {real, imag} */,
  {32'h3f333d81, 32'hbeaf8710} /* (15, 14, 12) {real, imag} */,
  {32'h3d28e550, 32'h3f1d99b4} /* (15, 14, 11) {real, imag} */,
  {32'hbd8a0d90, 32'h3e3c7ce8} /* (15, 14, 10) {real, imag} */,
  {32'hbf1e9f1a, 32'hbe222b60} /* (15, 14, 9) {real, imag} */,
  {32'hbe805318, 32'h3e55d9c0} /* (15, 14, 8) {real, imag} */,
  {32'h3ed410dc, 32'hbe814320} /* (15, 14, 7) {real, imag} */,
  {32'hbd664620, 32'hbf3e1d5c} /* (15, 14, 6) {real, imag} */,
  {32'h3d5d903c, 32'h3dc06460} /* (15, 14, 5) {real, imag} */,
  {32'h3eb69d86, 32'h3f07c7f0} /* (15, 14, 4) {real, imag} */,
  {32'h3e2e2d98, 32'h3dbb7ec0} /* (15, 14, 3) {real, imag} */,
  {32'h3e0616c4, 32'h3e9788c0} /* (15, 14, 2) {real, imag} */,
  {32'h3e10cf78, 32'h3ec262e0} /* (15, 14, 1) {real, imag} */,
  {32'hbdd956f0, 32'hbe8ba940} /* (15, 14, 0) {real, imag} */,
  {32'h3ea23b14, 32'h3dee34b0} /* (15, 13, 31) {real, imag} */,
  {32'h3e9e3be9, 32'h3e90c320} /* (15, 13, 30) {real, imag} */,
  {32'hbd16dd30, 32'h3f36aeb0} /* (15, 13, 29) {real, imag} */,
  {32'h3f22d9a0, 32'h3d29fb80} /* (15, 13, 28) {real, imag} */,
  {32'h3d300ce0, 32'hbe8419c0} /* (15, 13, 27) {real, imag} */,
  {32'hbf8df90e, 32'hbd148d40} /* (15, 13, 26) {real, imag} */,
  {32'hbf7d953e, 32'h3ed45770} /* (15, 13, 25) {real, imag} */,
  {32'hbf0b7d76, 32'h3d843b00} /* (15, 13, 24) {real, imag} */,
  {32'hbf316f74, 32'hbe9bc350} /* (15, 13, 23) {real, imag} */,
  {32'h3ea4c6ce, 32'hbf01f4e0} /* (15, 13, 22) {real, imag} */,
  {32'h3d1753e0, 32'hbf02067c} /* (15, 13, 21) {real, imag} */,
  {32'h3f38f7e8, 32'hbd82f4c0} /* (15, 13, 20) {real, imag} */,
  {32'h3f3fe360, 32'hbdcc5400} /* (15, 13, 19) {real, imag} */,
  {32'h3e731b90, 32'h3e6ea0f0} /* (15, 13, 18) {real, imag} */,
  {32'h3ed3ecba, 32'h3f2b5844} /* (15, 13, 17) {real, imag} */,
  {32'h3f206e35, 32'h3f0791f8} /* (15, 13, 16) {real, imag} */,
  {32'h3ef8b5c4, 32'hbe81d690} /* (15, 13, 15) {real, imag} */,
  {32'h3e8dc3fe, 32'hbe8aa0d0} /* (15, 13, 14) {real, imag} */,
  {32'h3e519368, 32'h3d7fe000} /* (15, 13, 13) {real, imag} */,
  {32'h3efbc068, 32'h3f1420a8} /* (15, 13, 12) {real, imag} */,
  {32'h3e854772, 32'h3f802a0e} /* (15, 13, 11) {real, imag} */,
  {32'hbea21280, 32'h3e48de90} /* (15, 13, 10) {real, imag} */,
  {32'hbe64b680, 32'hbe22f740} /* (15, 13, 9) {real, imag} */,
  {32'h3ea956c0, 32'hbec06ff0} /* (15, 13, 8) {real, imag} */,
  {32'h3e5cc0f2, 32'hbf03e2e8} /* (15, 13, 7) {real, imag} */,
  {32'hbe910c44, 32'hbeb818f0} /* (15, 13, 6) {real, imag} */,
  {32'hbebe8238, 32'hbde70b00} /* (15, 13, 5) {real, imag} */,
  {32'hbec9338c, 32'h3c810300} /* (15, 13, 4) {real, imag} */,
  {32'hbf07c446, 32'hbf1b74d0} /* (15, 13, 3) {real, imag} */,
  {32'h3e1495ee, 32'hbec7aa48} /* (15, 13, 2) {real, imag} */,
  {32'h3e775e08, 32'hbbef4400} /* (15, 13, 1) {real, imag} */,
  {32'hbc362300, 32'h3ebe0690} /* (15, 13, 0) {real, imag} */,
  {32'h3e675958, 32'hbcd64900} /* (15, 12, 31) {real, imag} */,
  {32'h3eab34ea, 32'h3ed74be0} /* (15, 12, 30) {real, imag} */,
  {32'hbe457900, 32'h3f1fdff8} /* (15, 12, 29) {real, imag} */,
  {32'h3ec60568, 32'hbe91e360} /* (15, 12, 28) {real, imag} */,
  {32'h3d89ee90, 32'hbf7c661c} /* (15, 12, 27) {real, imag} */,
  {32'hbddc28e0, 32'hbecba3b0} /* (15, 12, 26) {real, imag} */,
  {32'hbd0217a0, 32'h3f08258c} /* (15, 12, 25) {real, imag} */,
  {32'h3dbbda00, 32'h3d000780} /* (15, 12, 24) {real, imag} */,
  {32'hbecf3fdf, 32'hbdab3b80} /* (15, 12, 23) {real, imag} */,
  {32'h3f1cb42e, 32'h3ed204c8} /* (15, 12, 22) {real, imag} */,
  {32'h3e4da818, 32'hbee072bc} /* (15, 12, 21) {real, imag} */,
  {32'h3f5f8a09, 32'hbeb646d0} /* (15, 12, 20) {real, imag} */,
  {32'h3f81dddd, 32'h3eef4690} /* (15, 12, 19) {real, imag} */,
  {32'h3e01553e, 32'h3e5214e0} /* (15, 12, 18) {real, imag} */,
  {32'hbe1abf02, 32'h3e4f79a0} /* (15, 12, 17) {real, imag} */,
  {32'h3ee242a3, 32'h3eb27940} /* (15, 12, 16) {real, imag} */,
  {32'h3e2e3ea0, 32'hbe0c1400} /* (15, 12, 15) {real, imag} */,
  {32'hbea82010, 32'hbe121e20} /* (15, 12, 14) {real, imag} */,
  {32'hbe93a8b0, 32'h3e9c0750} /* (15, 12, 13) {real, imag} */,
  {32'h3eaa60d0, 32'hbde4cb00} /* (15, 12, 12) {real, imag} */,
  {32'h3eb97ec6, 32'h3c6a0300} /* (15, 12, 11) {real, imag} */,
  {32'hbe1efb20, 32'h3eceabd8} /* (15, 12, 10) {real, imag} */,
  {32'h3e1507f0, 32'h3e1919a0} /* (15, 12, 9) {real, imag} */,
  {32'hbdad61a0, 32'hbefd9fe0} /* (15, 12, 8) {real, imag} */,
  {32'hbe88b3b2, 32'hbe7fd240} /* (15, 12, 7) {real, imag} */,
  {32'hbebd40fa, 32'h3d15da00} /* (15, 12, 6) {real, imag} */,
  {32'hbf25653f, 32'hbd165c80} /* (15, 12, 5) {real, imag} */,
  {32'hbf9578d1, 32'h3db4b9c0} /* (15, 12, 4) {real, imag} */,
  {32'hbfae8320, 32'hbedf3840} /* (15, 12, 3) {real, imag} */,
  {32'hbd855a68, 32'hbead655c} /* (15, 12, 2) {real, imag} */,
  {32'h3e2f43f0, 32'hbe829be0} /* (15, 12, 1) {real, imag} */,
  {32'hbe78c7ec, 32'h3da3a6e0} /* (15, 12, 0) {real, imag} */,
  {32'hbda04188, 32'h3e55ae38} /* (15, 11, 31) {real, imag} */,
  {32'h3daa43e0, 32'h3f2929dc} /* (15, 11, 30) {real, imag} */,
  {32'h3d2f3804, 32'h3f103480} /* (15, 11, 29) {real, imag} */,
  {32'hbd0a01b8, 32'hbe61e4e0} /* (15, 11, 28) {real, imag} */,
  {32'hbeb688ae, 32'hbf997866} /* (15, 11, 27) {real, imag} */,
  {32'h3da8e038, 32'hbf66d37c} /* (15, 11, 26) {real, imag} */,
  {32'h3ea6f5d8, 32'h3f0fae10} /* (15, 11, 25) {real, imag} */,
  {32'hbebb5364, 32'h3c80f000} /* (15, 11, 24) {real, imag} */,
  {32'hbf937060, 32'hbeee4260} /* (15, 11, 23) {real, imag} */,
  {32'h3ec698f0, 32'hbe5f0b50} /* (15, 11, 22) {real, imag} */,
  {32'h3f6536c2, 32'hbe03ff34} /* (15, 11, 21) {real, imag} */,
  {32'h3fa74998, 32'hbe3dc5f0} /* (15, 11, 20) {real, imag} */,
  {32'h3f6a6377, 32'h3ea1ce58} /* (15, 11, 19) {real, imag} */,
  {32'hbe9c78e2, 32'h3f27cc74} /* (15, 11, 18) {real, imag} */,
  {32'hbef76828, 32'h3e50a390} /* (15, 11, 17) {real, imag} */,
  {32'h3e87368c, 32'hbe82dc98} /* (15, 11, 16) {real, imag} */,
  {32'h3e942339, 32'h3c9eb700} /* (15, 11, 15) {real, imag} */,
  {32'hbe88546c, 32'h3d829ac0} /* (15, 11, 14) {real, imag} */,
  {32'hbedd806e, 32'hbd6a9380} /* (15, 11, 13) {real, imag} */,
  {32'h3d50ca40, 32'hbf09bc7c} /* (15, 11, 12) {real, imag} */,
  {32'h3ea565a8, 32'hbec35078} /* (15, 11, 11) {real, imag} */,
  {32'h3e9a82be, 32'hbe084f90} /* (15, 11, 10) {real, imag} */,
  {32'h3e62356c, 32'hbf6b2f98} /* (15, 11, 9) {real, imag} */,
  {32'hbf8c3f48, 32'hbf864b0c} /* (15, 11, 8) {real, imag} */,
  {32'hbf2c83ba, 32'hbeb830e0} /* (15, 11, 7) {real, imag} */,
  {32'hbf3e6116, 32'h3e4f6f20} /* (15, 11, 6) {real, imag} */,
  {32'hbf1301b6, 32'h3dcb5d40} /* (15, 11, 5) {real, imag} */,
  {32'hbf1c6afa, 32'h3e8a5460} /* (15, 11, 4) {real, imag} */,
  {32'hbf46eb29, 32'h3eade128} /* (15, 11, 3) {real, imag} */,
  {32'hbeb69fa8, 32'hbe8bd120} /* (15, 11, 2) {real, imag} */,
  {32'h3d0c0900, 32'hbf0550a8} /* (15, 11, 1) {real, imag} */,
  {32'hbdb344d0, 32'hbcec3620} /* (15, 11, 0) {real, imag} */,
  {32'hbdc05fc8, 32'hbeb5a520} /* (15, 10, 31) {real, imag} */,
  {32'h3e14a79f, 32'h3e9982c0} /* (15, 10, 30) {real, imag} */,
  {32'hbf36d843, 32'h3e39bc70} /* (15, 10, 29) {real, imag} */,
  {32'hbec2fd26, 32'hbd1eb700} /* (15, 10, 28) {real, imag} */,
  {32'hbe3661d0, 32'hbec53330} /* (15, 10, 27) {real, imag} */,
  {32'hbe966c06, 32'hbea2d318} /* (15, 10, 26) {real, imag} */,
  {32'hbd9d5d70, 32'h3dee78b8} /* (15, 10, 25) {real, imag} */,
  {32'hbd0e9540, 32'h3d1d2b6c} /* (15, 10, 24) {real, imag} */,
  {32'hbf33c8a0, 32'hbf417218} /* (15, 10, 23) {real, imag} */,
  {32'h3f22b9fb, 32'hbf6605a8} /* (15, 10, 22) {real, imag} */,
  {32'h3f763166, 32'h3e837680} /* (15, 10, 21) {real, imag} */,
  {32'h3fa9ff1c, 32'hbc894af0} /* (15, 10, 20) {real, imag} */,
  {32'h3ddab6b4, 32'hbf5102a4} /* (15, 10, 19) {real, imag} */,
  {32'hbf2eaaff, 32'h3e7f8b60} /* (15, 10, 18) {real, imag} */,
  {32'hbe5f74c0, 32'h3f405348} /* (15, 10, 17) {real, imag} */,
  {32'hbd66e7c0, 32'h3ee97d50} /* (15, 10, 16) {real, imag} */,
  {32'h3f156356, 32'h3f268064} /* (15, 10, 15) {real, imag} */,
  {32'hbcd30b00, 32'h3f24e11c} /* (15, 10, 14) {real, imag} */,
  {32'hbcbf9dc0, 32'hbe020c00} /* (15, 10, 13) {real, imag} */,
  {32'h3e83f33c, 32'h3ebf3960} /* (15, 10, 12) {real, imag} */,
  {32'h3c8d2670, 32'hbd962e80} /* (15, 10, 11) {real, imag} */,
  {32'h3e924696, 32'hbf4cf58b} /* (15, 10, 10) {real, imag} */,
  {32'h3f11012c, 32'hbf3b7a96} /* (15, 10, 9) {real, imag} */,
  {32'hbf408bd1, 32'hbe725428} /* (15, 10, 8) {real, imag} */,
  {32'hbe4e3bf0, 32'h3da43ac0} /* (15, 10, 7) {real, imag} */,
  {32'h3dda1d68, 32'h3e1714b8} /* (15, 10, 6) {real, imag} */,
  {32'hbd7c461c, 32'hbd8b1b80} /* (15, 10, 5) {real, imag} */,
  {32'hbe887e88, 32'h3f0308ec} /* (15, 10, 4) {real, imag} */,
  {32'hbf2b2500, 32'h3eefcf50} /* (15, 10, 3) {real, imag} */,
  {32'hbf747efa, 32'hbbe9adc0} /* (15, 10, 2) {real, imag} */,
  {32'hbf4b9958, 32'hbf1b3697} /* (15, 10, 1) {real, imag} */,
  {32'hbeb0882e, 32'hbef6f01a} /* (15, 10, 0) {real, imag} */,
  {32'hbeae9aaa, 32'hbe567df0} /* (15, 9, 31) {real, imag} */,
  {32'h3dde07c0, 32'hbd61fa00} /* (15, 9, 30) {real, imag} */,
  {32'hbf1cfa28, 32'hbe0eeb40} /* (15, 9, 29) {real, imag} */,
  {32'hbec143bf, 32'h3ce3d200} /* (15, 9, 28) {real, imag} */,
  {32'h3ef594fe, 32'h3e51fd60} /* (15, 9, 27) {real, imag} */,
  {32'hbe618c12, 32'h3c9ba400} /* (15, 9, 26) {real, imag} */,
  {32'hbe7074f0, 32'hbeeac950} /* (15, 9, 25) {real, imag} */,
  {32'h3ce680e0, 32'hbe2157c0} /* (15, 9, 24) {real, imag} */,
  {32'h3cf5c8c0, 32'hbeb8eaf0} /* (15, 9, 23) {real, imag} */,
  {32'h3d451f20, 32'hbeebb3c8} /* (15, 9, 22) {real, imag} */,
  {32'h3e8b2497, 32'hbc8c9700} /* (15, 9, 21) {real, imag} */,
  {32'h3f3dbb77, 32'h3e8d0990} /* (15, 9, 20) {real, imag} */,
  {32'h3e47123a, 32'hbf8214b2} /* (15, 9, 19) {real, imag} */,
  {32'hbeb5e034, 32'hbe4fa620} /* (15, 9, 18) {real, imag} */,
  {32'hbf31088c, 32'h3f4d1ce0} /* (15, 9, 17) {real, imag} */,
  {32'hbef82088, 32'h3ebcf1f0} /* (15, 9, 16) {real, imag} */,
  {32'hbc157d00, 32'h3eb0bbc0} /* (15, 9, 15) {real, imag} */,
  {32'hbf255116, 32'h3e7c3b40} /* (15, 9, 14) {real, imag} */,
  {32'hbdcbb970, 32'hbe3be900} /* (15, 9, 13) {real, imag} */,
  {32'hbe88f52e, 32'h3d159b40} /* (15, 9, 12) {real, imag} */,
  {32'hbf001538, 32'hbf0709b0} /* (15, 9, 11) {real, imag} */,
  {32'h3e49d7b8, 32'hbf5922f7} /* (15, 9, 10) {real, imag} */,
  {32'h3f24e006, 32'hbda96d00} /* (15, 9, 9) {real, imag} */,
  {32'h3e94cff8, 32'h3f14c738} /* (15, 9, 8) {real, imag} */,
  {32'h3e09da90, 32'h3ed509f0} /* (15, 9, 7) {real, imag} */,
  {32'h3ebd6b38, 32'h3d4ebe80} /* (15, 9, 6) {real, imag} */,
  {32'h3f3c41ba, 32'hbee07270} /* (15, 9, 5) {real, imag} */,
  {32'h3e4d3328, 32'h3da4fa80} /* (15, 9, 4) {real, imag} */,
  {32'hbd45c458, 32'h3f0b68d0} /* (15, 9, 3) {real, imag} */,
  {32'h3db01a60, 32'hbe5e5800} /* (15, 9, 2) {real, imag} */,
  {32'h3db95b94, 32'h3d1ad080} /* (15, 9, 1) {real, imag} */,
  {32'h3e08fca8, 32'h3d604c80} /* (15, 9, 0) {real, imag} */,
  {32'hbf21fa4e, 32'hbe2c2248} /* (15, 8, 31) {real, imag} */,
  {32'hbf002872, 32'hbe511560} /* (15, 8, 30) {real, imag} */,
  {32'hbe686f70, 32'h3e052a60} /* (15, 8, 29) {real, imag} */,
  {32'h3d2e5168, 32'hbe5af2e0} /* (15, 8, 28) {real, imag} */,
  {32'h3eadad6e, 32'hbe665e80} /* (15, 8, 27) {real, imag} */,
  {32'h3e8c76b6, 32'h3e816fe0} /* (15, 8, 26) {real, imag} */,
  {32'h3de15f98, 32'h3f17e158} /* (15, 8, 25) {real, imag} */,
  {32'hbf1501ee, 32'h3f3237e0} /* (15, 8, 24) {real, imag} */,
  {32'hbe988bdb, 32'hbdc85a80} /* (15, 8, 23) {real, imag} */,
  {32'hbd21eca0, 32'h3d780800} /* (15, 8, 22) {real, imag} */,
  {32'h3ee3de29, 32'h3f07f618} /* (15, 8, 21) {real, imag} */,
  {32'h3e8caf88, 32'h3e92ba28} /* (15, 8, 20) {real, imag} */,
  {32'hbd8b8760, 32'hbed4d2f0} /* (15, 8, 19) {real, imag} */,
  {32'hbed804a1, 32'h3eac4be0} /* (15, 8, 18) {real, imag} */,
  {32'hbf7113ce, 32'h3f1f8914} /* (15, 8, 17) {real, imag} */,
  {32'hbe8f8850, 32'h3e603ce0} /* (15, 8, 16) {real, imag} */,
  {32'hbdb70ccc, 32'hbbab0400} /* (15, 8, 15) {real, imag} */,
  {32'hbf518300, 32'hbeae9440} /* (15, 8, 14) {real, imag} */,
  {32'hbedf63d0, 32'hbac0a000} /* (15, 8, 13) {real, imag} */,
  {32'hbf595d7f, 32'h3f0092e8} /* (15, 8, 12) {real, imag} */,
  {32'hbf291dfe, 32'hbe3cad20} /* (15, 8, 11) {real, imag} */,
  {32'h3ededc6a, 32'hbe3d9680} /* (15, 8, 10) {real, imag} */,
  {32'h3ecc2d54, 32'h3e981d28} /* (15, 8, 9) {real, imag} */,
  {32'h3d34c7f0, 32'h3e8be0b0} /* (15, 8, 8) {real, imag} */,
  {32'h3c41f0a0, 32'h3e5797a0} /* (15, 8, 7) {real, imag} */,
  {32'h3f063b12, 32'h3f1de4b8} /* (15, 8, 6) {real, imag} */,
  {32'h3f2dda32, 32'hbbc6b400} /* (15, 8, 5) {real, imag} */,
  {32'h3eb07b60, 32'hbca53e80} /* (15, 8, 4) {real, imag} */,
  {32'h3e6a9380, 32'h3e352520} /* (15, 8, 3) {real, imag} */,
  {32'h3f290f06, 32'hbe765010} /* (15, 8, 2) {real, imag} */,
  {32'h3f078fcc, 32'hbd9f07a0} /* (15, 8, 1) {real, imag} */,
  {32'h3f0cdfcc, 32'h3e1b3db0} /* (15, 8, 0) {real, imag} */,
  {32'hbf078332, 32'hbe613b30} /* (15, 7, 31) {real, imag} */,
  {32'hbf4d4740, 32'hbcd1ee00} /* (15, 7, 30) {real, imag} */,
  {32'hbf197733, 32'h3f0bf218} /* (15, 7, 29) {real, imag} */,
  {32'h3ecf600c, 32'h3ebacb50} /* (15, 7, 28) {real, imag} */,
  {32'h3dffc3b0, 32'hbdbaf520} /* (15, 7, 27) {real, imag} */,
  {32'h3ee278e4, 32'hbe40de90} /* (15, 7, 26) {real, imag} */,
  {32'h3f83410f, 32'h3ee4ac90} /* (15, 7, 25) {real, imag} */,
  {32'h3e1b34c4, 32'h3e12de20} /* (15, 7, 24) {real, imag} */,
  {32'h3e494748, 32'hbf106460} /* (15, 7, 23) {real, imag} */,
  {32'h3f4dae99, 32'hbea07240} /* (15, 7, 22) {real, imag} */,
  {32'h3f2700a6, 32'h3ebfc220} /* (15, 7, 21) {real, imag} */,
  {32'hbeda4328, 32'hbdea3ac0} /* (15, 7, 20) {real, imag} */,
  {32'hbf3c0cdd, 32'hbeef2a88} /* (15, 7, 19) {real, imag} */,
  {32'hbe5b90b2, 32'h3e4617f0} /* (15, 7, 18) {real, imag} */,
  {32'hbf4dd990, 32'h3e4026c0} /* (15, 7, 17) {real, imag} */,
  {32'hbe90b46d, 32'hbd7ca000} /* (15, 7, 16) {real, imag} */,
  {32'h3ec51f42, 32'h3d52cd80} /* (15, 7, 15) {real, imag} */,
  {32'h3f39b4e0, 32'h3e628680} /* (15, 7, 14) {real, imag} */,
  {32'hbd9ddee0, 32'hbc88cb00} /* (15, 7, 13) {real, imag} */,
  {32'hbf76cc60, 32'h3c037e00} /* (15, 7, 12) {real, imag} */,
  {32'hbf403662, 32'h3ed084a0} /* (15, 7, 11) {real, imag} */,
  {32'h3eafbc30, 32'h3ea78cc8} /* (15, 7, 10) {real, imag} */,
  {32'h3f3b5c73, 32'h3e25d2d0} /* (15, 7, 9) {real, imag} */,
  {32'hbe57d2a0, 32'hbdd6b980} /* (15, 7, 8) {real, imag} */,
  {32'hbe39dc78, 32'hbf144d30} /* (15, 7, 7) {real, imag} */,
  {32'h3e99a9cf, 32'hbda5bd00} /* (15, 7, 6) {real, imag} */,
  {32'h3f6c2d68, 32'h3e890f10} /* (15, 7, 5) {real, imag} */,
  {32'h3f634d3c, 32'hbea616b8} /* (15, 7, 4) {real, imag} */,
  {32'h3f132cce, 32'h3e85f590} /* (15, 7, 3) {real, imag} */,
  {32'h3f0e8ec4, 32'hbd314300} /* (15, 7, 2) {real, imag} */,
  {32'h3ed2c195, 32'h3e30c680} /* (15, 7, 1) {real, imag} */,
  {32'h3ec4bc4e, 32'h3edd9230} /* (15, 7, 0) {real, imag} */,
  {32'hbe92c41c, 32'hbcc56700} /* (15, 6, 31) {real, imag} */,
  {32'hbe7114a8, 32'h3bbc4800} /* (15, 6, 30) {real, imag} */,
  {32'hbedb33e0, 32'h3e9fb8b8} /* (15, 6, 29) {real, imag} */,
  {32'hbe0d1b48, 32'h3e99f8f8} /* (15, 6, 28) {real, imag} */,
  {32'hbeaa5f9c, 32'h3e54f840} /* (15, 6, 27) {real, imag} */,
  {32'h3e3b0194, 32'h3cadd380} /* (15, 6, 26) {real, imag} */,
  {32'h3edb4cdc, 32'hbe116310} /* (15, 6, 25) {real, imag} */,
  {32'h3cd4d600, 32'hbe60cfc0} /* (15, 6, 24) {real, imag} */,
  {32'h3f616014, 32'hbda5f600} /* (15, 6, 23) {real, imag} */,
  {32'h3f6db643, 32'hbde92980} /* (15, 6, 22) {real, imag} */,
  {32'h3f1a67cd, 32'hbd1c0d00} /* (15, 6, 21) {real, imag} */,
  {32'hbec32297, 32'hbbf0f000} /* (15, 6, 20) {real, imag} */,
  {32'hbf3970e0, 32'hbe5aef30} /* (15, 6, 19) {real, imag} */,
  {32'hbd7926e0, 32'h3f15e9d8} /* (15, 6, 18) {real, imag} */,
  {32'hbe21708e, 32'h3f85b914} /* (15, 6, 17) {real, imag} */,
  {32'hbe531308, 32'h3ebbac30} /* (15, 6, 16) {real, imag} */,
  {32'hbdb65e80, 32'hbe1f3200} /* (15, 6, 15) {real, imag} */,
  {32'h3f638a82, 32'h3dfbfa40} /* (15, 6, 14) {real, imag} */,
  {32'h3ebacd94, 32'h3ea34500} /* (15, 6, 13) {real, imag} */,
  {32'hbf136527, 32'h3e46c900} /* (15, 6, 12) {real, imag} */,
  {32'hbefa2cda, 32'h3f4682b4} /* (15, 6, 11) {real, imag} */,
  {32'h3dbf75c0, 32'h3f2b4490} /* (15, 6, 10) {real, imag} */,
  {32'h3ebfba08, 32'h3e199240} /* (15, 6, 9) {real, imag} */,
  {32'hbeb3f465, 32'hbef49290} /* (15, 6, 8) {real, imag} */,
  {32'hbf0fd1be, 32'h3e3c9e00} /* (15, 6, 7) {real, imag} */,
  {32'hbecb3dd9, 32'h3e2b75e0} /* (15, 6, 6) {real, imag} */,
  {32'h3df2ad10, 32'hbea39160} /* (15, 6, 5) {real, imag} */,
  {32'h3eb9b730, 32'hbed08948} /* (15, 6, 4) {real, imag} */,
  {32'h3e9811d8, 32'h3ec35b60} /* (15, 6, 3) {real, imag} */,
  {32'h3e400cc8, 32'h3f087f20} /* (15, 6, 2) {real, imag} */,
  {32'hbe83a684, 32'h3edb3cb0} /* (15, 6, 1) {real, imag} */,
  {32'h3de58ba4, 32'h3ed09cc8} /* (15, 6, 0) {real, imag} */,
  {32'hbec3f13a, 32'h3db4cd40} /* (15, 5, 31) {real, imag} */,
  {32'h3dab7360, 32'h3dd69780} /* (15, 5, 30) {real, imag} */,
  {32'hbe430898, 32'h3e0652c0} /* (15, 5, 29) {real, imag} */,
  {32'hbefe5356, 32'h3ebeea10} /* (15, 5, 28) {real, imag} */,
  {32'hbf1c754e, 32'h3b8c8000} /* (15, 5, 27) {real, imag} */,
  {32'h3ea51ad2, 32'h3e3ecdb0} /* (15, 5, 26) {real, imag} */,
  {32'hbea3d233, 32'h3ef261b0} /* (15, 5, 25) {real, imag} */,
  {32'hbe8f0a8a, 32'hbeb52f30} /* (15, 5, 24) {real, imag} */,
  {32'h3f1a24b0, 32'hbe7341e0} /* (15, 5, 23) {real, imag} */,
  {32'h3eaf3fe4, 32'h3e44b860} /* (15, 5, 22) {real, imag} */,
  {32'hbeaee19c, 32'h3c154900} /* (15, 5, 21) {real, imag} */,
  {32'hbe9b04ae, 32'h3f02ebc4} /* (15, 5, 20) {real, imag} */,
  {32'h3d11eb40, 32'h3ed0c8d4} /* (15, 5, 19) {real, imag} */,
  {32'h3d527770, 32'h3f277ece} /* (15, 5, 18) {real, imag} */,
  {32'hbd91cf80, 32'h3f67bce5} /* (15, 5, 17) {real, imag} */,
  {32'hbf1841ce, 32'h3e2fec28} /* (15, 5, 16) {real, imag} */,
  {32'hbe8fc720, 32'hbe9835b0} /* (15, 5, 15) {real, imag} */,
  {32'h3e97866e, 32'h3d9e9e80} /* (15, 5, 14) {real, imag} */,
  {32'h3da26ee0, 32'h3edc80d8} /* (15, 5, 13) {real, imag} */,
  {32'hbee2f898, 32'h3edf30e0} /* (15, 5, 12) {real, imag} */,
  {32'hbeec33f4, 32'h3ed3c5f0} /* (15, 5, 11) {real, imag} */,
  {32'hbf025a67, 32'h3e3dd220} /* (15, 5, 10) {real, imag} */,
  {32'h3ead1318, 32'h3ec57048} /* (15, 5, 9) {real, imag} */,
  {32'hbdfef7e8, 32'h3e016868} /* (15, 5, 8) {real, imag} */,
  {32'hbf8a8997, 32'h3f9089e7} /* (15, 5, 7) {real, imag} */,
  {32'hbf4bec45, 32'h3ee89dc8} /* (15, 5, 6) {real, imag} */,
  {32'hbead5788, 32'hbf9eb0c6} /* (15, 5, 5) {real, imag} */,
  {32'hbd902330, 32'hbf53cb80} /* (15, 5, 4) {real, imag} */,
  {32'h3f5253c0, 32'hbd3c9100} /* (15, 5, 3) {real, imag} */,
  {32'h3ecc1f2c, 32'h3be23800} /* (15, 5, 2) {real, imag} */,
  {32'hbd49c380, 32'hbf2fdd70} /* (15, 5, 1) {real, imag} */,
  {32'hbdab8e14, 32'hbe2a4230} /* (15, 5, 0) {real, imag} */,
  {32'hbefea862, 32'hbddab440} /* (15, 4, 31) {real, imag} */,
  {32'hbeb02d6e, 32'hbf22b8f0} /* (15, 4, 30) {real, imag} */,
  {32'h3e5a3194, 32'hbeaf7de8} /* (15, 4, 29) {real, imag} */,
  {32'hbebf4913, 32'h3f0897b0} /* (15, 4, 28) {real, imag} */,
  {32'hbf26efe4, 32'h3ea2fe80} /* (15, 4, 27) {real, imag} */,
  {32'hbe12f858, 32'hbd650000} /* (15, 4, 26) {real, imag} */,
  {32'hbe41d588, 32'hbebfe0b0} /* (15, 4, 25) {real, imag} */,
  {32'hbde0dd40, 32'hbf757d88} /* (15, 4, 24) {real, imag} */,
  {32'h3e09fc78, 32'hbf70a8b0} /* (15, 4, 23) {real, imag} */,
  {32'h3ee5e7aa, 32'hbbfb1000} /* (15, 4, 22) {real, imag} */,
  {32'hbea02210, 32'hbd330f00} /* (15, 4, 21) {real, imag} */,
  {32'hbe707d10, 32'h3e751440} /* (15, 4, 20) {real, imag} */,
  {32'h3e8c24d8, 32'hbd973e00} /* (15, 4, 19) {real, imag} */,
  {32'hbdf12bb8, 32'h3de95840} /* (15, 4, 18) {real, imag} */,
  {32'hbeca8e52, 32'h3cfb1000} /* (15, 4, 17) {real, imag} */,
  {32'hbe6ff924, 32'hbf77335c} /* (15, 4, 16) {real, imag} */,
  {32'h3e9109f8, 32'hbf217d20} /* (15, 4, 15) {real, imag} */,
  {32'h3f1da52c, 32'h3e03c870} /* (15, 4, 14) {real, imag} */,
  {32'h3dc357e0, 32'h3eb7e3d0} /* (15, 4, 13) {real, imag} */,
  {32'hbf514cd2, 32'hbdfca320} /* (15, 4, 12) {real, imag} */,
  {32'hbf070472, 32'h3e6a6440} /* (15, 4, 11) {real, imag} */,
  {32'hbea9adb8, 32'hbdde3c00} /* (15, 4, 10) {real, imag} */,
  {32'hbf2ea7aa, 32'hbed37770} /* (15, 4, 9) {real, imag} */,
  {32'hbf6e4056, 32'hbe41d1e0} /* (15, 4, 8) {real, imag} */,
  {32'hbf6ed3f1, 32'h3f144818} /* (15, 4, 7) {real, imag} */,
  {32'hbf3a0cc6, 32'h3f666fe8} /* (15, 4, 6) {real, imag} */,
  {32'hbe1a2b10, 32'hbd163ca8} /* (15, 4, 5) {real, imag} */,
  {32'h3e3044c0, 32'hbed72d60} /* (15, 4, 4) {real, imag} */,
  {32'h3f91eab2, 32'hbec62560} /* (15, 4, 3) {real, imag} */,
  {32'h3ebdaa41, 32'hbe706790} /* (15, 4, 2) {real, imag} */,
  {32'hbe499a22, 32'h3dabf440} /* (15, 4, 1) {real, imag} */,
  {32'hbe3d2076, 32'hbe1f44b0} /* (15, 4, 0) {real, imag} */,
  {32'hbe996cf4, 32'hbed34ca0} /* (15, 3, 31) {real, imag} */,
  {32'hbeb3d50e, 32'hbf7ec5cc} /* (15, 3, 30) {real, imag} */,
  {32'h3f135038, 32'hbe4b1460} /* (15, 3, 29) {real, imag} */,
  {32'h3f207d8c, 32'h3de3ce80} /* (15, 3, 28) {real, imag} */,
  {32'h3ec88999, 32'hbe993430} /* (15, 3, 27) {real, imag} */,
  {32'h3f2cdef1, 32'hbf507940} /* (15, 3, 26) {real, imag} */,
  {32'h3ece0492, 32'hbc4a1000} /* (15, 3, 25) {real, imag} */,
  {32'h3e825f24, 32'h3ebbc630} /* (15, 3, 24) {real, imag} */,
  {32'h3dfceab8, 32'h3e9c8ea0} /* (15, 3, 23) {real, imag} */,
  {32'h3f19b2c2, 32'h3e38f200} /* (15, 3, 22) {real, imag} */,
  {32'h3f0c8a3e, 32'h3ef41300} /* (15, 3, 21) {real, imag} */,
  {32'hbe082ae4, 32'h3e56d700} /* (15, 3, 20) {real, imag} */,
  {32'hbf3a7fae, 32'hbda83200} /* (15, 3, 19) {real, imag} */,
  {32'hbf87eff9, 32'hbe804c88} /* (15, 3, 18) {real, imag} */,
  {32'hbf2c9002, 32'hbe784600} /* (15, 3, 17) {real, imag} */,
  {32'h3e0f34a8, 32'hbf504c32} /* (15, 3, 16) {real, imag} */,
  {32'h3e0a64aa, 32'h3c226a00} /* (15, 3, 15) {real, imag} */,
  {32'h3e96bbf8, 32'h3e9ffb60} /* (15, 3, 14) {real, imag} */,
  {32'h3d7242a0, 32'h3eb3f590} /* (15, 3, 13) {real, imag} */,
  {32'hbf748516, 32'hbed155d0} /* (15, 3, 12) {real, imag} */,
  {32'hbe501fc0, 32'h3efda320} /* (15, 3, 11) {real, imag} */,
  {32'hbecb4caa, 32'h3e098420} /* (15, 3, 10) {real, imag} */,
  {32'hbf8a942e, 32'hbe9164c0} /* (15, 3, 9) {real, imag} */,
  {32'hbd848cd0, 32'h3e5f6a00} /* (15, 3, 8) {real, imag} */,
  {32'h3e84d114, 32'h3f980c2c} /* (15, 3, 7) {real, imag} */,
  {32'hbd3a36c0, 32'h3fba10e4} /* (15, 3, 6) {real, imag} */,
  {32'h3f3f6109, 32'h3f7c438d} /* (15, 3, 5) {real, imag} */,
  {32'h3f1d3255, 32'hbde731c0} /* (15, 3, 4) {real, imag} */,
  {32'h3f2b52ec, 32'hbf768b2c} /* (15, 3, 3) {real, imag} */,
  {32'h3f261002, 32'hbf6c1924} /* (15, 3, 2) {real, imag} */,
  {32'h3e9cdee4, 32'hbe486b40} /* (15, 3, 1) {real, imag} */,
  {32'h3e56e522, 32'hbed0bfc8} /* (15, 3, 0) {real, imag} */,
  {32'hbed9029f, 32'hbacb1c00} /* (15, 2, 31) {real, imag} */,
  {32'h3dff1320, 32'hbe4650c0} /* (15, 2, 30) {real, imag} */,
  {32'h3f7f2676, 32'hbeb9a1a0} /* (15, 2, 29) {real, imag} */,
  {32'h3fd3f55c, 32'hbe992140} /* (15, 2, 28) {real, imag} */,
  {32'h3f5ff9b6, 32'hbe9f0360} /* (15, 2, 27) {real, imag} */,
  {32'h3f11678e, 32'hbf674ffc} /* (15, 2, 26) {real, imag} */,
  {32'h3f021986, 32'h3e9da510} /* (15, 2, 25) {real, imag} */,
  {32'h3f8515c3, 32'h3e8e3750} /* (15, 2, 24) {real, imag} */,
  {32'h3ed7e2b2, 32'h3f2cfb10} /* (15, 2, 23) {real, imag} */,
  {32'h3e566fb0, 32'h3ed58d10} /* (15, 2, 22) {real, imag} */,
  {32'h3ec262dc, 32'hbe63b050} /* (15, 2, 21) {real, imag} */,
  {32'hbe1de84a, 32'hbeae61b0} /* (15, 2, 20) {real, imag} */,
  {32'hbf16e58f, 32'h3ebcad40} /* (15, 2, 19) {real, imag} */,
  {32'hbfc95664, 32'h3e0f3080} /* (15, 2, 18) {real, imag} */,
  {32'hbf324cac, 32'h3d627880} /* (15, 2, 17) {real, imag} */,
  {32'h3e4b4f2c, 32'hbe4f7ff0} /* (15, 2, 16) {real, imag} */,
  {32'hbe83067e, 32'h3e3a6d68} /* (15, 2, 15) {real, imag} */,
  {32'hbed038aa, 32'h3d6565c0} /* (15, 2, 14) {real, imag} */,
  {32'hbeab02c7, 32'hbd98e880} /* (15, 2, 13) {real, imag} */,
  {32'hbe8cd4fe, 32'hbf238598} /* (15, 2, 12) {real, imag} */,
  {32'h3dc6b028, 32'hbe55d240} /* (15, 2, 11) {real, imag} */,
  {32'hbf57da5f, 32'hbdf04400} /* (15, 2, 10) {real, imag} */,
  {32'hbf544b19, 32'h3ea0c820} /* (15, 2, 9) {real, imag} */,
  {32'h3e851186, 32'h3db23e80} /* (15, 2, 8) {real, imag} */,
  {32'h3e4e6e5c, 32'h3f73fd38} /* (15, 2, 7) {real, imag} */,
  {32'h3c5898c0, 32'h3fdb2ff4} /* (15, 2, 6) {real, imag} */,
  {32'h3f7e5e44, 32'h3f5ca278} /* (15, 2, 5) {real, imag} */,
  {32'h3ee98f20, 32'hbefc3870} /* (15, 2, 4) {real, imag} */,
  {32'hbe777c3c, 32'hbf287e90} /* (15, 2, 3) {real, imag} */,
  {32'h3f13cc12, 32'hbe96df20} /* (15, 2, 2) {real, imag} */,
  {32'h3ebc62c7, 32'h3ed88988} /* (15, 2, 1) {real, imag} */,
  {32'h3e3dcce4, 32'h3e9130dc} /* (15, 2, 0) {real, imag} */,
  {32'hbf1ad656, 32'h3ec91510} /* (15, 1, 31) {real, imag} */,
  {32'hbe586a2e, 32'h3d4cf940} /* (15, 1, 30) {real, imag} */,
  {32'h3ca06840, 32'hbf0e8620} /* (15, 1, 29) {real, imag} */,
  {32'h3e9ba038, 32'hbf29ff50} /* (15, 1, 28) {real, imag} */,
  {32'hbe17262e, 32'hbe173ac0} /* (15, 1, 27) {real, imag} */,
  {32'hbe5fb1c0, 32'h3eba8f58} /* (15, 1, 26) {real, imag} */,
  {32'hbe5d4e18, 32'h3f6a1cf4} /* (15, 1, 25) {real, imag} */,
  {32'h3cc0fdc0, 32'hbd693100} /* (15, 1, 24) {real, imag} */,
  {32'hbdd9dac0, 32'hbed21de8} /* (15, 1, 23) {real, imag} */,
  {32'h3daab8c0, 32'h3e2e5b88} /* (15, 1, 22) {real, imag} */,
  {32'h3e0c4708, 32'hbe3f8100} /* (15, 1, 21) {real, imag} */,
  {32'hbe3853d7, 32'hbf0ccac8} /* (15, 1, 20) {real, imag} */,
  {32'hbe205fd4, 32'h3e886a00} /* (15, 1, 19) {real, imag} */,
  {32'hbf6968b0, 32'h3f177358} /* (15, 1, 18) {real, imag} */,
  {32'hbdf77a60, 32'hbef97a60} /* (15, 1, 17) {real, imag} */,
  {32'hbe1c8142, 32'hbf663810} /* (15, 1, 16) {real, imag} */,
  {32'hbe54216a, 32'h3b3c6200} /* (15, 1, 15) {real, imag} */,
  {32'h3eecb161, 32'hbec51640} /* (15, 1, 14) {real, imag} */,
  {32'h3d80a4f0, 32'hbf0e5c48} /* (15, 1, 13) {real, imag} */,
  {32'hbe167ecc, 32'hbf259750} /* (15, 1, 12) {real, imag} */,
  {32'hbea34ec4, 32'hbef80570} /* (15, 1, 11) {real, imag} */,
  {32'hbf05ed52, 32'h3f0b5838} /* (15, 1, 10) {real, imag} */,
  {32'hbe08ff58, 32'h3ee41390} /* (15, 1, 9) {real, imag} */,
  {32'h3ede188c, 32'hbe9b7170} /* (15, 1, 8) {real, imag} */,
  {32'h3cc791c0, 32'h3dd50ec0} /* (15, 1, 7) {real, imag} */,
  {32'hbe33cdb8, 32'h3f7ea39c} /* (15, 1, 6) {real, imag} */,
  {32'hbe18d9d4, 32'h3eed5e6c} /* (15, 1, 5) {real, imag} */,
  {32'hbe146774, 32'hbf0cb2f0} /* (15, 1, 4) {real, imag} */,
  {32'hbea8ecf4, 32'hbda8f7c0} /* (15, 1, 3) {real, imag} */,
  {32'h3ea4082e, 32'h3f1aac0c} /* (15, 1, 2) {real, imag} */,
  {32'h3e75e692, 32'h3f4e6264} /* (15, 1, 1) {real, imag} */,
  {32'hbb927d00, 32'h3f2c22bb} /* (15, 1, 0) {real, imag} */,
  {32'hbe8e0127, 32'hbe180230} /* (15, 0, 31) {real, imag} */,
  {32'hbed1d47d, 32'h3df08ca0} /* (15, 0, 30) {real, imag} */,
  {32'hbf1f8cc0, 32'h3ec8d9e8} /* (15, 0, 29) {real, imag} */,
  {32'hbe60fa38, 32'h3de139a0} /* (15, 0, 28) {real, imag} */,
  {32'hbe919bc5, 32'h3ed1f6d0} /* (15, 0, 27) {real, imag} */,
  {32'hbd83cc74, 32'h3ee79af0} /* (15, 0, 26) {real, imag} */,
  {32'h3bb6ca00, 32'h3f0c4590} /* (15, 0, 25) {real, imag} */,
  {32'hbe90c1e3, 32'hbe2dfca8} /* (15, 0, 24) {real, imag} */,
  {32'hbea8f684, 32'hbf1ee9b2} /* (15, 0, 23) {real, imag} */,
  {32'h3e13a2f8, 32'h3d77d9b8} /* (15, 0, 22) {real, imag} */,
  {32'h3e85ddc4, 32'hbda8e480} /* (15, 0, 21) {real, imag} */,
  {32'hbdce49b0, 32'hbf190886} /* (15, 0, 20) {real, imag} */,
  {32'hbd1941a8, 32'hbe917060} /* (15, 0, 19) {real, imag} */,
  {32'hbe18637c, 32'h3e87fea8} /* (15, 0, 18) {real, imag} */,
  {32'h3e656fd0, 32'hbee33840} /* (15, 0, 17) {real, imag} */,
  {32'hbe396768, 32'hbe9093e8} /* (15, 0, 16) {real, imag} */,
  {32'hbe6ad578, 32'h3e91ff10} /* (15, 0, 15) {real, imag} */,
  {32'h3e627c98, 32'hbe7a1500} /* (15, 0, 14) {real, imag} */,
  {32'h3e741fbc, 32'h3e1e9f60} /* (15, 0, 13) {real, imag} */,
  {32'hbe32b268, 32'h3e3b3f70} /* (15, 0, 12) {real, imag} */,
  {32'hbf30a782, 32'h3e048940} /* (15, 0, 11) {real, imag} */,
  {32'hbeb93976, 32'h3f1ffedc} /* (15, 0, 10) {real, imag} */,
  {32'hbdf56baf, 32'h3ed53a38} /* (15, 0, 9) {real, imag} */,
  {32'h3e49b1c1, 32'hbe1d30b0} /* (15, 0, 8) {real, imag} */,
  {32'hbe75bcf8, 32'h3db353b0} /* (15, 0, 7) {real, imag} */,
  {32'h3e1bb980, 32'h3f00f06c} /* (15, 0, 6) {real, imag} */,
  {32'hbe053c44, 32'h3e9d1d7a} /* (15, 0, 5) {real, imag} */,
  {32'hbec2740a, 32'h3d5dd430} /* (15, 0, 4) {real, imag} */,
  {32'h3c866da0, 32'h3e9b68b0} /* (15, 0, 3) {real, imag} */,
  {32'h3ed856e4, 32'h3e9fea38} /* (15, 0, 2) {real, imag} */,
  {32'h3f2a4788, 32'h3ded3820} /* (15, 0, 1) {real, imag} */,
  {32'h3f047024, 32'h3e72aac0} /* (15, 0, 0) {real, imag} */,
  {32'hbe358a0c, 32'h3d08aae0} /* (14, 31, 31) {real, imag} */,
  {32'hbf2f9e5d, 32'h3f0116d8} /* (14, 31, 30) {real, imag} */,
  {32'hbf3f4cd3, 32'h3e467100} /* (14, 31, 29) {real, imag} */,
  {32'hbf1d620c, 32'h3da4d400} /* (14, 31, 28) {real, imag} */,
  {32'hbe903168, 32'h3e269f40} /* (14, 31, 27) {real, imag} */,
  {32'hbe446cc8, 32'hbe036ea0} /* (14, 31, 26) {real, imag} */,
  {32'h3e3aadc8, 32'hbe6d8040} /* (14, 31, 25) {real, imag} */,
  {32'h3ed1fd04, 32'hbe597fe0} /* (14, 31, 24) {real, imag} */,
  {32'hbe473990, 32'h3eceb5b8} /* (14, 31, 23) {real, imag} */,
  {32'hbe146f98, 32'h3e9b1a80} /* (14, 31, 22) {real, imag} */,
  {32'h3f1aa943, 32'hbd0ddf00} /* (14, 31, 21) {real, imag} */,
  {32'h3f50012e, 32'h3f030cf0} /* (14, 31, 20) {real, imag} */,
  {32'hbd1c50e0, 32'h3e871450} /* (14, 31, 19) {real, imag} */,
  {32'hbeb44aa5, 32'hbe3837d0} /* (14, 31, 18) {real, imag} */,
  {32'h3e436452, 32'hbe46ec20} /* (14, 31, 17) {real, imag} */,
  {32'h3e99f1f7, 32'hbe078800} /* (14, 31, 16) {real, imag} */,
  {32'h3eeabdea, 32'hbe8394b0} /* (14, 31, 15) {real, imag} */,
  {32'h3f242754, 32'hbf13ba30} /* (14, 31, 14) {real, imag} */,
  {32'h3e9e68b8, 32'hbe52adc0} /* (14, 31, 13) {real, imag} */,
  {32'hbefa6fa0, 32'hbec8d2b8} /* (14, 31, 12) {real, imag} */,
  {32'hbe7ec214, 32'hbf869c74} /* (14, 31, 11) {real, imag} */,
  {32'h3e82fd64, 32'hbe362d14} /* (14, 31, 10) {real, imag} */,
  {32'hbee8c7d0, 32'h3edf0800} /* (14, 31, 9) {real, imag} */,
  {32'hbf300884, 32'hbe6eeb40} /* (14, 31, 8) {real, imag} */,
  {32'hbeb20770, 32'hbef7e6b8} /* (14, 31, 7) {real, imag} */,
  {32'hbf13de40, 32'h3df5a9c0} /* (14, 31, 6) {real, imag} */,
  {32'hbf3a0baa, 32'h3e911f60} /* (14, 31, 5) {real, imag} */,
  {32'hbf07379e, 32'h3ec789c8} /* (14, 31, 4) {real, imag} */,
  {32'hbf7b3ca5, 32'h3f205648} /* (14, 31, 3) {real, imag} */,
  {32'hbecd5432, 32'h3f056da8} /* (14, 31, 2) {real, imag} */,
  {32'hbf0a681d, 32'hbdea9c40} /* (14, 31, 1) {real, imag} */,
  {32'hbe94894c, 32'hbcdd5180} /* (14, 31, 0) {real, imag} */,
  {32'hbf4baa78, 32'hbf386958} /* (14, 30, 31) {real, imag} */,
  {32'hbf85ddc2, 32'hbf87dab0} /* (14, 30, 30) {real, imag} */,
  {32'hbef999c0, 32'hbf1fdee8} /* (14, 30, 29) {real, imag} */,
  {32'hbf5f1614, 32'hbe5b2e60} /* (14, 30, 28) {real, imag} */,
  {32'hbf7ca7f0, 32'hbe6024c0} /* (14, 30, 27) {real, imag} */,
  {32'hbedcb0d2, 32'hbe9a97a0} /* (14, 30, 26) {real, imag} */,
  {32'h3cf44b20, 32'hbd468300} /* (14, 30, 25) {real, imag} */,
  {32'h3e7071c4, 32'hbf205e40} /* (14, 30, 24) {real, imag} */,
  {32'h3cceeb60, 32'h3eae55e0} /* (14, 30, 23) {real, imag} */,
  {32'hbec3c5fc, 32'h3efc65d0} /* (14, 30, 22) {real, imag} */,
  {32'h3ec984f4, 32'hbefa0248} /* (14, 30, 21) {real, imag} */,
  {32'h3f26b704, 32'hbe96f608} /* (14, 30, 20) {real, imag} */,
  {32'h3e9c46f8, 32'h3eae07b0} /* (14, 30, 19) {real, imag} */,
  {32'hbe54dda0, 32'h3cfa1800} /* (14, 30, 18) {real, imag} */,
  {32'h3ea9002f, 32'hbcbe4b00} /* (14, 30, 17) {real, imag} */,
  {32'h3ecd97e8, 32'h3b0bd800} /* (14, 30, 16) {real, imag} */,
  {32'h3eb7686c, 32'hbea66180} /* (14, 30, 15) {real, imag} */,
  {32'h3f1b2c1e, 32'hbf7686f0} /* (14, 30, 14) {real, imag} */,
  {32'hbd994540, 32'hbe789b80} /* (14, 30, 13) {real, imag} */,
  {32'hbf2e6ee7, 32'hbe376700} /* (14, 30, 12) {real, imag} */,
  {32'h3e6f1e00, 32'hbf67eeb8} /* (14, 30, 11) {real, imag} */,
  {32'h3efa75e8, 32'hbed72340} /* (14, 30, 10) {real, imag} */,
  {32'hbea7fcf6, 32'h3f6b5ff0} /* (14, 30, 9) {real, imag} */,
  {32'hbefb0bf4, 32'hbebf52a0} /* (14, 30, 8) {real, imag} */,
  {32'hbce50e00, 32'hbf567b58} /* (14, 30, 7) {real, imag} */,
  {32'hbf372e8a, 32'h3ee43ae0} /* (14, 30, 6) {real, imag} */,
  {32'hbf6832c0, 32'h3e8f95a0} /* (14, 30, 5) {real, imag} */,
  {32'hbecba320, 32'h3d8e8700} /* (14, 30, 4) {real, imag} */,
  {32'hbe15b9e0, 32'h3f086080} /* (14, 30, 3) {real, imag} */,
  {32'hbf13de94, 32'h3ea97780} /* (14, 30, 2) {real, imag} */,
  {32'hbf28ba0d, 32'hbe85ec40} /* (14, 30, 1) {real, imag} */,
  {32'hbd39f060, 32'hbf13b710} /* (14, 30, 0) {real, imag} */,
  {32'hbf6d4d08, 32'h3dcf0380} /* (14, 29, 31) {real, imag} */,
  {32'hbf1dcd28, 32'hbe510540} /* (14, 29, 30) {real, imag} */,
  {32'h3f1be1f4, 32'hbe48b480} /* (14, 29, 29) {real, imag} */,
  {32'h3c189500, 32'hbed5fd40} /* (14, 29, 28) {real, imag} */,
  {32'hbf943470, 32'hbef57690} /* (14, 29, 27) {real, imag} */,
  {32'hbfb8a09a, 32'hbf1df280} /* (14, 29, 26) {real, imag} */,
  {32'hbf54470b, 32'hbd864f00} /* (14, 29, 25) {real, imag} */,
  {32'hbf2b19c4, 32'hbe2a4200} /* (14, 29, 24) {real, imag} */,
  {32'hbef70fc0, 32'h3f2dc5f0} /* (14, 29, 23) {real, imag} */,
  {32'hbe8d0ca8, 32'h3ed9e330} /* (14, 29, 22) {real, imag} */,
  {32'hbe3980be, 32'hbe8723fc} /* (14, 29, 21) {real, imag} */,
  {32'h3d9f46c0, 32'hbe62ea80} /* (14, 29, 20) {real, imag} */,
  {32'h3dbdd4d0, 32'h3f229070} /* (14, 29, 19) {real, imag} */,
  {32'h3f69cca2, 32'hbeb40ce0} /* (14, 29, 18) {real, imag} */,
  {32'h3f0e9734, 32'hbeb61b60} /* (14, 29, 17) {real, imag} */,
  {32'hbd3811c0, 32'h3f17dbd0} /* (14, 29, 16) {real, imag} */,
  {32'hbe11c030, 32'hbe887a30} /* (14, 29, 15) {real, imag} */,
  {32'h3e228f00, 32'hbf946e68} /* (14, 29, 14) {real, imag} */,
  {32'hbd014000, 32'hbf384ec0} /* (14, 29, 13) {real, imag} */,
  {32'hbe2ffea0, 32'hbef1b950} /* (14, 29, 12) {real, imag} */,
  {32'h3f744746, 32'h3e8432e0} /* (14, 29, 11) {real, imag} */,
  {32'h3e915638, 32'h3e478da0} /* (14, 29, 10) {real, imag} */,
  {32'hbf0f99b2, 32'h3faa4a30} /* (14, 29, 9) {real, imag} */,
  {32'hbebe4850, 32'h3ebf9000} /* (14, 29, 8) {real, imag} */,
  {32'hbec26d78, 32'hbf20c6d0} /* (14, 29, 7) {real, imag} */,
  {32'hbf1f6d84, 32'h3df46f00} /* (14, 29, 6) {real, imag} */,
  {32'hbe38b720, 32'h3ec853b0} /* (14, 29, 5) {real, imag} */,
  {32'h3e4e9540, 32'h3ed5fec0} /* (14, 29, 4) {real, imag} */,
  {32'h3f40c99c, 32'h3e2ad0a0} /* (14, 29, 3) {real, imag} */,
  {32'hbf043c88, 32'hbdba1000} /* (14, 29, 2) {real, imag} */,
  {32'hbef6d81e, 32'hbe92c460} /* (14, 29, 1) {real, imag} */,
  {32'hbc52a300, 32'hbf31611c} /* (14, 29, 0) {real, imag} */,
  {32'hbe772718, 32'h3f0b3fa4} /* (14, 28, 31) {real, imag} */,
  {32'h3e3f6fc8, 32'h3f1aa380} /* (14, 28, 30) {real, imag} */,
  {32'h3fbbb5dd, 32'hbe6f5d00} /* (14, 28, 29) {real, imag} */,
  {32'h3c97d580, 32'hbf139f68} /* (14, 28, 28) {real, imag} */,
  {32'hbf846fa2, 32'h3d0f2700} /* (14, 28, 27) {real, imag} */,
  {32'hbf87b06c, 32'hbeacec40} /* (14, 28, 26) {real, imag} */,
  {32'hbf876313, 32'h3c51b600} /* (14, 28, 25) {real, imag} */,
  {32'hbf463950, 32'hbe755280} /* (14, 28, 24) {real, imag} */,
  {32'hbf6c9630, 32'h3edfb880} /* (14, 28, 23) {real, imag} */,
  {32'hbee909fc, 32'h3eebe400} /* (14, 28, 22) {real, imag} */,
  {32'hbf11abc0, 32'h3f17f630} /* (14, 28, 21) {real, imag} */,
  {32'hbde410e0, 32'h3da1f680} /* (14, 28, 20) {real, imag} */,
  {32'hbe2d2a80, 32'h3edaf6e0} /* (14, 28, 19) {real, imag} */,
  {32'h3f3f3560, 32'h3e90e280} /* (14, 28, 18) {real, imag} */,
  {32'hbea8acbc, 32'h3d81b180} /* (14, 28, 17) {real, imag} */,
  {32'hbec96038, 32'h3ee211e0} /* (14, 28, 16) {real, imag} */,
  {32'h3e8b3be0, 32'h3cde4c00} /* (14, 28, 15) {real, imag} */,
  {32'h3f558260, 32'hbf035230} /* (14, 28, 14) {real, imag} */,
  {32'h3f2a7018, 32'hbf0f9c50} /* (14, 28, 13) {real, imag} */,
  {32'h3f41438e, 32'hbed5d160} /* (14, 28, 12) {real, imag} */,
  {32'h3e9b200c, 32'h3f0615e0} /* (14, 28, 11) {real, imag} */,
  {32'hbe296380, 32'h3ee7b0a8} /* (14, 28, 10) {real, imag} */,
  {32'hbedb2764, 32'h3ea5c940} /* (14, 28, 9) {real, imag} */,
  {32'hbf781a5c, 32'h3e4fc8e0} /* (14, 28, 8) {real, imag} */,
  {32'hbf1ed412, 32'hbe80ad40} /* (14, 28, 7) {real, imag} */,
  {32'hbf379b86, 32'hbee89100} /* (14, 28, 6) {real, imag} */,
  {32'hbf01b6dc, 32'h3d87b280} /* (14, 28, 5) {real, imag} */,
  {32'hbddaecc0, 32'hbf251810} /* (14, 28, 4) {real, imag} */,
  {32'h3cb17e80, 32'h3e7dd540} /* (14, 28, 3) {real, imag} */,
  {32'hbed377b0, 32'h3e2f4d80} /* (14, 28, 2) {real, imag} */,
  {32'hbf053aa5, 32'hbe60e080} /* (14, 28, 1) {real, imag} */,
  {32'hbeed5626, 32'hbd87bc80} /* (14, 28, 0) {real, imag} */,
  {32'h3e339fa0, 32'h3ede6670} /* (14, 27, 31) {real, imag} */,
  {32'h3eeea1c4, 32'h3edb2c10} /* (14, 27, 30) {real, imag} */,
  {32'h3f9b10e8, 32'h3d30f600} /* (14, 27, 29) {real, imag} */,
  {32'hbf78b712, 32'hbf3fec90} /* (14, 27, 28) {real, imag} */,
  {32'hc01045e8, 32'hbe86eda0} /* (14, 27, 27) {real, imag} */,
  {32'hbfaa7cea, 32'h3ec8a5c0} /* (14, 27, 26) {real, imag} */,
  {32'hbf42fa6e, 32'h3fa5b754} /* (14, 27, 25) {real, imag} */,
  {32'hbf669a68, 32'h3f3e68d0} /* (14, 27, 24) {real, imag} */,
  {32'hbf2e8368, 32'h3fc2a2b8} /* (14, 27, 23) {real, imag} */,
  {32'hbf433664, 32'h3f808da0} /* (14, 27, 22) {real, imag} */,
  {32'hbf4f9972, 32'h3d83be80} /* (14, 27, 21) {real, imag} */,
  {32'hbe9c64a8, 32'hbda7a340} /* (14, 27, 20) {real, imag} */,
  {32'h3d8c57a0, 32'hbc441200} /* (14, 27, 19) {real, imag} */,
  {32'h3f307cb4, 32'h3e9cc420} /* (14, 27, 18) {real, imag} */,
  {32'h3ee57928, 32'h3ea14180} /* (14, 27, 17) {real, imag} */,
  {32'h3e7c36e0, 32'h3f1fcc50} /* (14, 27, 16) {real, imag} */,
  {32'h3f890d75, 32'h3ea99440} /* (14, 27, 15) {real, imag} */,
  {32'h3f3cefd0, 32'h3f0c47c8} /* (14, 27, 14) {real, imag} */,
  {32'h3cb8df00, 32'hbda161c0} /* (14, 27, 13) {real, imag} */,
  {32'hbebd18a0, 32'h3db72f80} /* (14, 27, 12) {real, imag} */,
  {32'hbf927a27, 32'h3f293040} /* (14, 27, 11) {real, imag} */,
  {32'hbf4e3be2, 32'h3e81e178} /* (14, 27, 10) {real, imag} */,
  {32'hbe0bf188, 32'hbf36a760} /* (14, 27, 9) {real, imag} */,
  {32'hbe5e3fec, 32'hbea2ad80} /* (14, 27, 8) {real, imag} */,
  {32'hbe9b1970, 32'hbd607600} /* (14, 27, 7) {real, imag} */,
  {32'hbead4ca4, 32'hbdc75f80} /* (14, 27, 6) {real, imag} */,
  {32'hbec11b48, 32'hbf045bd0} /* (14, 27, 5) {real, imag} */,
  {32'hbec7dc58, 32'hbec91b30} /* (14, 27, 4) {real, imag} */,
  {32'hbf29f0d7, 32'h3e97da70} /* (14, 27, 3) {real, imag} */,
  {32'hbed633c8, 32'hbed48640} /* (14, 27, 2) {real, imag} */,
  {32'hbe5898a0, 32'hbedec670} /* (14, 27, 1) {real, imag} */,
  {32'hbf3b0f04, 32'hbd040100} /* (14, 27, 0) {real, imag} */,
  {32'hbebd6768, 32'h3ed1db30} /* (14, 26, 31) {real, imag} */,
  {32'hbe988694, 32'h3f5be578} /* (14, 26, 30) {real, imag} */,
  {32'h3e4bd520, 32'h3f855058} /* (14, 26, 29) {real, imag} */,
  {32'hbedcb8ee, 32'h3d32c400} /* (14, 26, 28) {real, imag} */,
  {32'hbfa19bf7, 32'h3ed5b4b0} /* (14, 26, 27) {real, imag} */,
  {32'hbf838169, 32'h3f829c28} /* (14, 26, 26) {real, imag} */,
  {32'hbf1f44a4, 32'h3f07bfa0} /* (14, 26, 25) {real, imag} */,
  {32'hbf06bfa8, 32'h3f4eaaa0} /* (14, 26, 24) {real, imag} */,
  {32'hbf0a795a, 32'h3f75ff80} /* (14, 26, 23) {real, imag} */,
  {32'hbe83d7cc, 32'h3d6ba480} /* (14, 26, 22) {real, imag} */,
  {32'h3e5e8cec, 32'hbe9d7260} /* (14, 26, 21) {real, imag} */,
  {32'h3f3e914c, 32'h3c9f6b00} /* (14, 26, 20) {real, imag} */,
  {32'h3f613b2a, 32'hbe513900} /* (14, 26, 19) {real, imag} */,
  {32'h3fd8bf16, 32'hbf3464a8} /* (14, 26, 18) {real, imag} */,
  {32'h3f9d18d0, 32'hbe9f3780} /* (14, 26, 17) {real, imag} */,
  {32'h3ee5c098, 32'h3f11feb0} /* (14, 26, 16) {real, imag} */,
  {32'h3f2f5d5c, 32'hbee34e60} /* (14, 26, 15) {real, imag} */,
  {32'h3ed42908, 32'h3ed6e240} /* (14, 26, 14) {real, imag} */,
  {32'h3dd7eff0, 32'h3dc6e640} /* (14, 26, 13) {real, imag} */,
  {32'h3de54c20, 32'h3e7a06a0} /* (14, 26, 12) {real, imag} */,
  {32'h3d8ae950, 32'h3f500c78} /* (14, 26, 11) {real, imag} */,
  {32'hbe7e42e4, 32'h3ea62ed8} /* (14, 26, 10) {real, imag} */,
  {32'hbefc32f4, 32'h3bd95000} /* (14, 26, 9) {real, imag} */,
  {32'hbecbf860, 32'hbd78cc00} /* (14, 26, 8) {real, imag} */,
  {32'hbf6d3394, 32'h3e9a1ba0} /* (14, 26, 7) {real, imag} */,
  {32'hbe301f70, 32'hbbf6f400} /* (14, 26, 6) {real, imag} */,
  {32'hbd6939c0, 32'h3e042580} /* (14, 26, 5) {real, imag} */,
  {32'h3e3e21a0, 32'h3e8a76e0} /* (14, 26, 4) {real, imag} */,
  {32'h3d996948, 32'hbd67f480} /* (14, 26, 3) {real, imag} */,
  {32'hbf1d2006, 32'hbf0c6b70} /* (14, 26, 2) {real, imag} */,
  {32'h3e0af280, 32'hbe62a2c0} /* (14, 26, 1) {real, imag} */,
  {32'h3dae1960, 32'h3dec6880} /* (14, 26, 0) {real, imag} */,
  {32'hbe991058, 32'h3a8d1800} /* (14, 25, 31) {real, imag} */,
  {32'h3d94f560, 32'h3f3df430} /* (14, 25, 30) {real, imag} */,
  {32'h3cd854a0, 32'h3f4ad790} /* (14, 25, 29) {real, imag} */,
  {32'h3e03c380, 32'h3e1c9340} /* (14, 25, 28) {real, imag} */,
  {32'hbedcb2ea, 32'h3ea2d0f0} /* (14, 25, 27) {real, imag} */,
  {32'hbf1dc185, 32'h3f934e80} /* (14, 25, 26) {real, imag} */,
  {32'hbee5cb6e, 32'h3df20980} /* (14, 25, 25) {real, imag} */,
  {32'hbe9f9150, 32'h3efa6540} /* (14, 25, 24) {real, imag} */,
  {32'hbe0212a0, 32'h3e88d220} /* (14, 25, 23) {real, imag} */,
  {32'hbeeb6984, 32'hbf08f250} /* (14, 25, 22) {real, imag} */,
  {32'hbdd40a1c, 32'hbe4c54a0} /* (14, 25, 21) {real, imag} */,
  {32'h3ee31a68, 32'h3ec35e10} /* (14, 25, 20) {real, imag} */,
  {32'h3f4b43a0, 32'hbe31f980} /* (14, 25, 19) {real, imag} */,
  {32'h3f9b762f, 32'hbf80d1e8} /* (14, 25, 18) {real, imag} */,
  {32'h3f0cefca, 32'hbf354270} /* (14, 25, 17) {real, imag} */,
  {32'h3f147ed6, 32'hbc147800} /* (14, 25, 16) {real, imag} */,
  {32'h3f5c8c44, 32'hbf636ca0} /* (14, 25, 15) {real, imag} */,
  {32'h3f73b650, 32'hbf17a680} /* (14, 25, 14) {real, imag} */,
  {32'h3fa4080e, 32'hbec9b2c0} /* (14, 25, 13) {real, imag} */,
  {32'h3f3cef6e, 32'hbee50d20} /* (14, 25, 12) {real, imag} */,
  {32'h3e36b700, 32'h3ccced00} /* (14, 25, 11) {real, imag} */,
  {32'hbf2fc462, 32'h3e26ad40} /* (14, 25, 10) {real, imag} */,
  {32'hbf7233f0, 32'h3f94571c} /* (14, 25, 9) {real, imag} */,
  {32'hbf3be3f8, 32'h3f0b9590} /* (14, 25, 8) {real, imag} */,
  {32'hbf758a22, 32'h3e929f10} /* (14, 25, 7) {real, imag} */,
  {32'hbe9131ec, 32'hbf155b88} /* (14, 25, 6) {real, imag} */,
  {32'hbe527520, 32'hbeb8bf80} /* (14, 25, 5) {real, imag} */,
  {32'h3e34a360, 32'h3f13daf0} /* (14, 25, 4) {real, imag} */,
  {32'hbdb57af0, 32'h3f279680} /* (14, 25, 3) {real, imag} */,
  {32'hbf822aa3, 32'h3ecd3a20} /* (14, 25, 2) {real, imag} */,
  {32'hbf0fdb54, 32'h3e159ce0} /* (14, 25, 1) {real, imag} */,
  {32'hbe9a4fe4, 32'hbde4d2a0} /* (14, 25, 0) {real, imag} */,
  {32'h3d420940, 32'hbd0c6300} /* (14, 24, 31) {real, imag} */,
  {32'h3ef9c928, 32'h3e4f4140} /* (14, 24, 30) {real, imag} */,
  {32'hbe7781d0, 32'hbee6f8c0} /* (14, 24, 29) {real, imag} */,
  {32'hbf121cd6, 32'hbdc8af00} /* (14, 24, 28) {real, imag} */,
  {32'hbf9d2b98, 32'h3e0b2e20} /* (14, 24, 27) {real, imag} */,
  {32'hbf8148fc, 32'h3eb46e60} /* (14, 24, 26) {real, imag} */,
  {32'hbf1ae8ce, 32'hbdd79200} /* (14, 24, 25) {real, imag} */,
  {32'hbf2ad64e, 32'h3f048510} /* (14, 24, 24) {real, imag} */,
  {32'h3d69d480, 32'h3fa15ed0} /* (14, 24, 23) {real, imag} */,
  {32'hbf2eea88, 32'h3c5df400} /* (14, 24, 22) {real, imag} */,
  {32'hbf259117, 32'h3d32d240} /* (14, 24, 21) {real, imag} */,
  {32'hbf3618d4, 32'h3dccb400} /* (14, 24, 20) {real, imag} */,
  {32'h3f0915fc, 32'hbf4e6970} /* (14, 24, 19) {real, imag} */,
  {32'h3f3931c2, 32'hbfc7f178} /* (14, 24, 18) {real, imag} */,
  {32'h3f64ed9e, 32'hbf010118} /* (14, 24, 17) {real, imag} */,
  {32'h3f5e62a3, 32'hbc8aa600} /* (14, 24, 16) {real, imag} */,
  {32'hbdb092a0, 32'hbe51a780} /* (14, 24, 15) {real, imag} */,
  {32'h3f10102a, 32'hbf1bed10} /* (14, 24, 14) {real, imag} */,
  {32'h3f3e7a9a, 32'hbef2d900} /* (14, 24, 13) {real, imag} */,
  {32'h3f833c18, 32'hbf748580} /* (14, 24, 12) {real, imag} */,
  {32'h3e6990d0, 32'hbed9b9b0} /* (14, 24, 11) {real, imag} */,
  {32'hbf40db78, 32'h3ed59ff8} /* (14, 24, 10) {real, imag} */,
  {32'hbf1f23b4, 32'h3f5327d0} /* (14, 24, 9) {real, imag} */,
  {32'h3efaa124, 32'h3f2d4740} /* (14, 24, 8) {real, imag} */,
  {32'hbecf8684, 32'h3ea7a1e0} /* (14, 24, 7) {real, imag} */,
  {32'hbf22b6ea, 32'h3de6d080} /* (14, 24, 6) {real, imag} */,
  {32'hbee28390, 32'h3edcc390} /* (14, 24, 5) {real, imag} */,
  {32'hbcb52100, 32'h3ed9d360} /* (14, 24, 4) {real, imag} */,
  {32'h3d505440, 32'h3e6f5340} /* (14, 24, 3) {real, imag} */,
  {32'hbfa5ab06, 32'hbe180c40} /* (14, 24, 2) {real, imag} */,
  {32'hbfafe866, 32'hbf675d80} /* (14, 24, 1) {real, imag} */,
  {32'hbf0ac25e, 32'hbf0f440c} /* (14, 24, 0) {real, imag} */,
  {32'hbe89ee12, 32'h3f5b3488} /* (14, 23, 31) {real, imag} */,
  {32'hbefe02ec, 32'h3ee15020} /* (14, 23, 30) {real, imag} */,
  {32'hbf2d3f77, 32'hbdeb3480} /* (14, 23, 29) {real, imag} */,
  {32'hbf1b9334, 32'hbd5b1700} /* (14, 23, 28) {real, imag} */,
  {32'hbf0dd5bc, 32'hbdb8d500} /* (14, 23, 27) {real, imag} */,
  {32'hbf899e2d, 32'h3e9502d0} /* (14, 23, 26) {real, imag} */,
  {32'hbf5724ce, 32'hbe988fe0} /* (14, 23, 25) {real, imag} */,
  {32'hbf32706f, 32'h3ccc0d00} /* (14, 23, 24) {real, imag} */,
  {32'hbc06f980, 32'h3f3d9b10} /* (14, 23, 23) {real, imag} */,
  {32'hbf2d2959, 32'h3eb0a6e0} /* (14, 23, 22) {real, imag} */,
  {32'hbf413d2a, 32'h3d7cdfc0} /* (14, 23, 21) {real, imag} */,
  {32'h3ecd52f0, 32'h3db28a40} /* (14, 23, 20) {real, imag} */,
  {32'h3f6fe27a, 32'hbdef0400} /* (14, 23, 19) {real, imag} */,
  {32'h3f566c96, 32'hbf44c7e0} /* (14, 23, 18) {real, imag} */,
  {32'h3fcea78f, 32'hbd3a4c00} /* (14, 23, 17) {real, imag} */,
  {32'h3fca72de, 32'hbe1fc860} /* (14, 23, 16) {real, imag} */,
  {32'h3ec8ecb0, 32'hbefb90e0} /* (14, 23, 15) {real, imag} */,
  {32'h3c3b2640, 32'hbe95ccc0} /* (14, 23, 14) {real, imag} */,
  {32'h3e321178, 32'hbee04cf0} /* (14, 23, 13) {real, imag} */,
  {32'h3f9e4901, 32'hbf6cb138} /* (14, 23, 12) {real, imag} */,
  {32'hbdc49480, 32'hbe34e980} /* (14, 23, 11) {real, imag} */,
  {32'hbf93e224, 32'h3ef25970} /* (14, 23, 10) {real, imag} */,
  {32'hbf695948, 32'hbdcbf840} /* (14, 23, 9) {real, imag} */,
  {32'h3f019508, 32'h3eb11440} /* (14, 23, 8) {real, imag} */,
  {32'hbe40a0a8, 32'h3f08d050} /* (14, 23, 7) {real, imag} */,
  {32'hbdc19270, 32'h3f302e10} /* (14, 23, 6) {real, imag} */,
  {32'h3c407ac0, 32'h3f8e70b4} /* (14, 23, 5) {real, imag} */,
  {32'hbf1246a2, 32'h3f695330} /* (14, 23, 4) {real, imag} */,
  {32'hbeeec85c, 32'h3f017be0} /* (14, 23, 3) {real, imag} */,
  {32'hbf37841c, 32'hbde67e00} /* (14, 23, 2) {real, imag} */,
  {32'hbef462a4, 32'hbf8c55b4} /* (14, 23, 1) {real, imag} */,
  {32'hbc8d0fb0, 32'hbe7b4aa0} /* (14, 23, 0) {real, imag} */,
  {32'hbf63616f, 32'h3e928ef0} /* (14, 22, 31) {real, imag} */,
  {32'hbf2d9843, 32'hbed95100} /* (14, 22, 30) {real, imag} */,
  {32'hbe0691d8, 32'hbde7a300} /* (14, 22, 29) {real, imag} */,
  {32'h3e59e790, 32'h3ee3e8c0} /* (14, 22, 28) {real, imag} */,
  {32'h3efcde00, 32'h3eb493f0} /* (14, 22, 27) {real, imag} */,
  {32'hbdc95ee0, 32'h3f16d1f8} /* (14, 22, 26) {real, imag} */,
  {32'hbed6439c, 32'hbeaadd50} /* (14, 22, 25) {real, imag} */,
  {32'hbf92f798, 32'hbe166700} /* (14, 22, 24) {real, imag} */,
  {32'hbef8428a, 32'hbed3d2b0} /* (14, 22, 23) {real, imag} */,
  {32'hbeca71c8, 32'hbed2cec0} /* (14, 22, 22) {real, imag} */,
  {32'hbf796bb8, 32'h3d85f0a0} /* (14, 22, 21) {real, imag} */,
  {32'h3e82ef06, 32'hbd51fb00} /* (14, 22, 20) {real, imag} */,
  {32'h3fa5d495, 32'h3e95f3f0} /* (14, 22, 19) {real, imag} */,
  {32'h3f850a2a, 32'h3ce1ee00} /* (14, 22, 18) {real, imag} */,
  {32'h3f889b48, 32'h3e94e1e0} /* (14, 22, 17) {real, imag} */,
  {32'h3f9d1f90, 32'hbe7a1e20} /* (14, 22, 16) {real, imag} */,
  {32'h3f282fcc, 32'h3b752000} /* (14, 22, 15) {real, imag} */,
  {32'h3f34e526, 32'h3f2787b0} /* (14, 22, 14) {real, imag} */,
  {32'h3f2e11f0, 32'hbd69e200} /* (14, 22, 13) {real, imag} */,
  {32'h3e71b028, 32'h3ec949c0} /* (14, 22, 12) {real, imag} */,
  {32'hbde38cc0, 32'h3e2867c0} /* (14, 22, 11) {real, imag} */,
  {32'hbf31e752, 32'hbe945aa0} /* (14, 22, 10) {real, imag} */,
  {32'hbf2c439c, 32'hbefca820} /* (14, 22, 9) {real, imag} */,
  {32'hbecd228c, 32'hbeba3980} /* (14, 22, 8) {real, imag} */,
  {32'hbf28a748, 32'hbdd8d400} /* (14, 22, 7) {real, imag} */,
  {32'hbf193747, 32'h3e0ce880} /* (14, 22, 6) {real, imag} */,
  {32'hbe9b991e, 32'h3e42e840} /* (14, 22, 5) {real, imag} */,
  {32'hbf173d8c, 32'hbc5c0a00} /* (14, 22, 4) {real, imag} */,
  {32'hbf999c5d, 32'h3eaef450} /* (14, 22, 3) {real, imag} */,
  {32'hbf338db8, 32'h3f4d5780} /* (14, 22, 2) {real, imag} */,
  {32'hbea1d4a8, 32'h3e1463c0} /* (14, 22, 1) {real, imag} */,
  {32'hbedb3249, 32'h3e560de0} /* (14, 22, 0) {real, imag} */,
  {32'hbf1b3004, 32'hbe84231c} /* (14, 21, 31) {real, imag} */,
  {32'hbf6b91ae, 32'hbf30128c} /* (14, 21, 30) {real, imag} */,
  {32'hbf3a8099, 32'hbef06408} /* (14, 21, 29) {real, imag} */,
  {32'hbf0cc7fc, 32'h3ef9bd80} /* (14, 21, 28) {real, imag} */,
  {32'h3dfa1e40, 32'h3f56eb14} /* (14, 21, 27) {real, imag} */,
  {32'h3f15e298, 32'h3ee80ed8} /* (14, 21, 26) {real, imag} */,
  {32'h3e74aa88, 32'h3e053632} /* (14, 21, 25) {real, imag} */,
  {32'hbe960594, 32'h3e253968} /* (14, 21, 24) {real, imag} */,
  {32'h3effc094, 32'hbee6b740} /* (14, 21, 23) {real, imag} */,
  {32'hbf040c6a, 32'hbee18ff0} /* (14, 21, 22) {real, imag} */,
  {32'hbf96991e, 32'h3e8e1550} /* (14, 21, 21) {real, imag} */,
  {32'hbf32daaa, 32'h3f207f9e} /* (14, 21, 20) {real, imag} */,
  {32'h3ddf4f00, 32'h3f028f00} /* (14, 21, 19) {real, imag} */,
  {32'h3f522507, 32'hbce39180} /* (14, 21, 18) {real, imag} */,
  {32'h3f8ff9b3, 32'h3f2f89ca} /* (14, 21, 17) {real, imag} */,
  {32'h3ea1ecab, 32'h3ca65000} /* (14, 21, 16) {real, imag} */,
  {32'hbe5394d4, 32'hbe944e40} /* (14, 21, 15) {real, imag} */,
  {32'h3f58a677, 32'h3ef439a0} /* (14, 21, 14) {real, imag} */,
  {32'h39c7f800, 32'h3ef842b0} /* (14, 21, 13) {real, imag} */,
  {32'hbf60ace9, 32'h3fb324e4} /* (14, 21, 12) {real, imag} */,
  {32'h3e015c78, 32'h3f1ac0f0} /* (14, 21, 11) {real, imag} */,
  {32'hbd2beab8, 32'hbec177fc} /* (14, 21, 10) {real, imag} */,
  {32'hbea0d75c, 32'hbd51abc0} /* (14, 21, 9) {real, imag} */,
  {32'hbea7af7c, 32'h3e2e6b10} /* (14, 21, 8) {real, imag} */,
  {32'hbf41de3b, 32'hbf291b14} /* (14, 21, 7) {real, imag} */,
  {32'hbf64edca, 32'hbeec6264} /* (14, 21, 6) {real, imag} */,
  {32'hbef995c7, 32'hbe2871b0} /* (14, 21, 5) {real, imag} */,
  {32'h3ea99e94, 32'hbf57fcf0} /* (14, 21, 4) {real, imag} */,
  {32'hbd0a22b0, 32'hbebc7758} /* (14, 21, 3) {real, imag} */,
  {32'hbdbbe100, 32'hbe5e4480} /* (14, 21, 2) {real, imag} */,
  {32'hbf150309, 32'hbeb65720} /* (14, 21, 1) {real, imag} */,
  {32'hbef81c9c, 32'h3d3a6500} /* (14, 21, 0) {real, imag} */,
  {32'hbe6e1d76, 32'h3e7841b0} /* (14, 20, 31) {real, imag} */,
  {32'h3d536640, 32'h3ee758b0} /* (14, 20, 30) {real, imag} */,
  {32'hbebd7814, 32'hbea0dca0} /* (14, 20, 29) {real, imag} */,
  {32'hbed5157c, 32'h3c9c0c00} /* (14, 20, 28) {real, imag} */,
  {32'h3ef900c4, 32'h3f06aa60} /* (14, 20, 27) {real, imag} */,
  {32'h3eedbbec, 32'h3f63cce8} /* (14, 20, 26) {real, imag} */,
  {32'h3f4062ce, 32'h3e4152c0} /* (14, 20, 25) {real, imag} */,
  {32'h3f27287c, 32'h3e245780} /* (14, 20, 24) {real, imag} */,
  {32'h3f702378, 32'h3f3d1160} /* (14, 20, 23) {real, imag} */,
  {32'hbf02e9e6, 32'h3f6ace50} /* (14, 20, 22) {real, imag} */,
  {32'hbf66f5cc, 32'h3ec8d41c} /* (14, 20, 21) {real, imag} */,
  {32'hbf839c96, 32'h3edd2a00} /* (14, 20, 20) {real, imag} */,
  {32'hbf9f457a, 32'h3ecf7030} /* (14, 20, 19) {real, imag} */,
  {32'h3ee79b46, 32'h3f288f28} /* (14, 20, 18) {real, imag} */,
  {32'h3e906e3a, 32'h3f877dc8} /* (14, 20, 17) {real, imag} */,
  {32'hbf46423e, 32'h3f02f2b0} /* (14, 20, 16) {real, imag} */,
  {32'hbf2149be, 32'hbe3abfa0} /* (14, 20, 15) {real, imag} */,
  {32'hbc834640, 32'hbdb34980} /* (14, 20, 14) {real, imag} */,
  {32'hbecb7fb0, 32'h3ee016d0} /* (14, 20, 13) {real, imag} */,
  {32'hbed50840, 32'h3f883570} /* (14, 20, 12) {real, imag} */,
  {32'hbcad80c0, 32'hbeabe4c8} /* (14, 20, 11) {real, imag} */,
  {32'h3e137bb0, 32'hbfa7cb8b} /* (14, 20, 10) {real, imag} */,
  {32'h3e186760, 32'hbc46b200} /* (14, 20, 9) {real, imag} */,
  {32'h3e93884c, 32'h3f396a6c} /* (14, 20, 8) {real, imag} */,
  {32'h3e7f8a48, 32'hbd9ae380} /* (14, 20, 7) {real, imag} */,
  {32'h3f0fc7a1, 32'hbe6d8880} /* (14, 20, 6) {real, imag} */,
  {32'h3f8e5980, 32'hbe298520} /* (14, 20, 5) {real, imag} */,
  {32'h3fa3b9ec, 32'hbeeb1990} /* (14, 20, 4) {real, imag} */,
  {32'h3f83a2d8, 32'hbf9407a0} /* (14, 20, 3) {real, imag} */,
  {32'h3f31cab0, 32'hbf9fce0c} /* (14, 20, 2) {real, imag} */,
  {32'h3eb08170, 32'hbf29fdd8} /* (14, 20, 1) {real, imag} */,
  {32'h3e8a3bd8, 32'h3e5669a0} /* (14, 20, 0) {real, imag} */,
  {32'h3f0122eb, 32'hba136000} /* (14, 19, 31) {real, imag} */,
  {32'h3f7f7800, 32'h3eb1d620} /* (14, 19, 30) {real, imag} */,
  {32'h3f739ce6, 32'hbf5eedf0} /* (14, 19, 29) {real, imag} */,
  {32'h3f9a5edc, 32'hbeb65420} /* (14, 19, 28) {real, imag} */,
  {32'h3f52dcbb, 32'h3e683a80} /* (14, 19, 27) {real, imag} */,
  {32'h3ee30d76, 32'h3ebd8280} /* (14, 19, 26) {real, imag} */,
  {32'h3f51f38a, 32'hbed4f960} /* (14, 19, 25) {real, imag} */,
  {32'h3f19c3c0, 32'hbec32500} /* (14, 19, 24) {real, imag} */,
  {32'h3f34edf4, 32'h3e3926c0} /* (14, 19, 23) {real, imag} */,
  {32'h3e8f7a3c, 32'h3f20c390} /* (14, 19, 22) {real, imag} */,
  {32'hbef2a33a, 32'h3f774cb0} /* (14, 19, 21) {real, imag} */,
  {32'hbf72e26a, 32'h3f7d9cc8} /* (14, 19, 20) {real, imag} */,
  {32'hbfadfbb8, 32'h3f093d60} /* (14, 19, 19) {real, imag} */,
  {32'hbe5ed82e, 32'h3f1faf78} /* (14, 19, 18) {real, imag} */,
  {32'hbdddfde0, 32'h3f43d310} /* (14, 19, 17) {real, imag} */,
  {32'hbf0b1898, 32'h3f18e4c8} /* (14, 19, 16) {real, imag} */,
  {32'hbe242a70, 32'h3f0b4640} /* (14, 19, 15) {real, imag} */,
  {32'hbdf42800, 32'h3e45efc0} /* (14, 19, 14) {real, imag} */,
  {32'hbef5336a, 32'h3eca3aa0} /* (14, 19, 13) {real, imag} */,
  {32'h3d31cdf0, 32'h3f76c5a0} /* (14, 19, 12) {real, imag} */,
  {32'h3e25af74, 32'hbee31190} /* (14, 19, 11) {real, imag} */,
  {32'h3e4ada1c, 32'hbf2dcdec} /* (14, 19, 10) {real, imag} */,
  {32'h3f1c52bc, 32'h3ee33c20} /* (14, 19, 9) {real, imag} */,
  {32'h3e25cf60, 32'h3e70afa0} /* (14, 19, 8) {real, imag} */,
  {32'h3e9894b0, 32'h3eb86500} /* (14, 19, 7) {real, imag} */,
  {32'h3e40349c, 32'h3edf8600} /* (14, 19, 6) {real, imag} */,
  {32'h3f5125f8, 32'h3e823540} /* (14, 19, 5) {real, imag} */,
  {32'h3f7fb76a, 32'h3ea025b0} /* (14, 19, 4) {real, imag} */,
  {32'h3f1217c4, 32'hbf36b238} /* (14, 19, 3) {real, imag} */,
  {32'h3fa21718, 32'hbf9a8348} /* (14, 19, 2) {real, imag} */,
  {32'h3fa0ce7e, 32'hbdff01c0} /* (14, 19, 1) {real, imag} */,
  {32'h3f0cfb8b, 32'h3f2c627c} /* (14, 19, 0) {real, imag} */,
  {32'h3ebdbd06, 32'h3d616080} /* (14, 18, 31) {real, imag} */,
  {32'h3f48a584, 32'h3f0d2f20} /* (14, 18, 30) {real, imag} */,
  {32'h3ebe9154, 32'hbeda1f50} /* (14, 18, 29) {real, imag} */,
  {32'h3f4cb151, 32'h3ddbbe00} /* (14, 18, 28) {real, imag} */,
  {32'h3f563a78, 32'h3f638708} /* (14, 18, 27) {real, imag} */,
  {32'h3f30563a, 32'hbe2f6700} /* (14, 18, 26) {real, imag} */,
  {32'h3f1b7be0, 32'hbf91ad38} /* (14, 18, 25) {real, imag} */,
  {32'h3fa54f60, 32'hbfa49974} /* (14, 18, 24) {real, imag} */,
  {32'h3ff01d04, 32'hbf3fc310} /* (14, 18, 23) {real, imag} */,
  {32'h3f4e218e, 32'h3e7ae3a0} /* (14, 18, 22) {real, imag} */,
  {32'hbeae4d41, 32'h3fd9c0ec} /* (14, 18, 21) {real, imag} */,
  {32'hbf4cf5d6, 32'h3f7e3b08} /* (14, 18, 20) {real, imag} */,
  {32'hbfbb08b6, 32'h3f46f3d0} /* (14, 18, 19) {real, imag} */,
  {32'hbffad278, 32'h3f6e8588} /* (14, 18, 18) {real, imag} */,
  {32'hbf7eb224, 32'h3f780f20} /* (14, 18, 17) {real, imag} */,
  {32'hbeeb51e8, 32'h3f067cf8} /* (14, 18, 16) {real, imag} */,
  {32'hbef75e30, 32'h3e9a2520} /* (14, 18, 15) {real, imag} */,
  {32'hbe7a0848, 32'hbdcea540} /* (14, 18, 14) {real, imag} */,
  {32'hbf145aee, 32'h3ea109c0} /* (14, 18, 13) {real, imag} */,
  {32'hbf2b1dda, 32'h3e1533c0} /* (14, 18, 12) {real, imag} */,
  {32'h3e98269c, 32'hbf50a758} /* (14, 18, 11) {real, imag} */,
  {32'h3c5fc2c0, 32'hbf04424c} /* (14, 18, 10) {real, imag} */,
  {32'h3daa2b30, 32'h3efd5960} /* (14, 18, 9) {real, imag} */,
  {32'h3f71fc8e, 32'h3e66b200} /* (14, 18, 8) {real, imag} */,
  {32'h3f92cf26, 32'h3b8e0000} /* (14, 18, 7) {real, imag} */,
  {32'h3f26a651, 32'hbe816e80} /* (14, 18, 6) {real, imag} */,
  {32'h3e54e0ec, 32'hbd8ef080} /* (14, 18, 5) {real, imag} */,
  {32'h3e999350, 32'hbd4e1580} /* (14, 18, 4) {real, imag} */,
  {32'h3ebaeef0, 32'hbedb8e20} /* (14, 18, 3) {real, imag} */,
  {32'h3f8f9af8, 32'hbe714d40} /* (14, 18, 2) {real, imag} */,
  {32'h3f9bbe10, 32'h3eb25f40} /* (14, 18, 1) {real, imag} */,
  {32'h3eaa526c, 32'h3f2942b8} /* (14, 18, 0) {real, imag} */,
  {32'h3de8b450, 32'h3ee73d40} /* (14, 17, 31) {real, imag} */,
  {32'h3e423210, 32'h3e98fd30} /* (14, 17, 30) {real, imag} */,
  {32'h3ebecd58, 32'hbe299400} /* (14, 17, 29) {real, imag} */,
  {32'h3f482fba, 32'h3ea663b0} /* (14, 17, 28) {real, imag} */,
  {32'h3f5a28ac, 32'h3f242178} /* (14, 17, 27) {real, imag} */,
  {32'h3f468de6, 32'hbd377900} /* (14, 17, 26) {real, imag} */,
  {32'h3f394772, 32'hbeaa28f0} /* (14, 17, 25) {real, imag} */,
  {32'h3f4a0228, 32'hbf25a8f0} /* (14, 17, 24) {real, imag} */,
  {32'h3f23f34c, 32'hbf0a2cb0} /* (14, 17, 23) {real, imag} */,
  {32'h3f8c1620, 32'hbf01a140} /* (14, 17, 22) {real, imag} */,
  {32'h3f2fdd29, 32'h3e066200} /* (14, 17, 21) {real, imag} */,
  {32'hbe3e9c50, 32'hba032000} /* (14, 17, 20) {real, imag} */,
  {32'h3e6dd3da, 32'h3de02d00} /* (14, 17, 19) {real, imag} */,
  {32'hbfa1955d, 32'h3f321280} /* (14, 17, 18) {real, imag} */,
  {32'hbffbc3ef, 32'h3fe34d54} /* (14, 17, 17) {real, imag} */,
  {32'hbf97a146, 32'h3f1d21a0} /* (14, 17, 16) {real, imag} */,
  {32'hbfa40a22, 32'h3c515a00} /* (14, 17, 15) {real, imag} */,
  {32'hbf9de5f2, 32'hbf049aa8} /* (14, 17, 14) {real, imag} */,
  {32'hbeba39f0, 32'hbe24d600} /* (14, 17, 13) {real, imag} */,
  {32'hbf033892, 32'hbf2e7950} /* (14, 17, 12) {real, imag} */,
  {32'h3dd02880, 32'hbf22a950} /* (14, 17, 11) {real, imag} */,
  {32'hbd42eb40, 32'hbe677e80} /* (14, 17, 10) {real, imag} */,
  {32'h3f31cae0, 32'hbcff8500} /* (14, 17, 9) {real, imag} */,
  {32'h3fb3d558, 32'hbe9211b0} /* (14, 17, 8) {real, imag} */,
  {32'h3faddb8b, 32'hbeb51d00} /* (14, 17, 7) {real, imag} */,
  {32'h3f689a92, 32'hbf0b3dd8} /* (14, 17, 6) {real, imag} */,
  {32'hbea44400, 32'hbd8a3780} /* (14, 17, 5) {real, imag} */,
  {32'hbed67bfc, 32'hbe1dd200} /* (14, 17, 4) {real, imag} */,
  {32'h3eced3f8, 32'hbd70e800} /* (14, 17, 3) {real, imag} */,
  {32'h3f14b166, 32'h3d773400} /* (14, 17, 2) {real, imag} */,
  {32'h3f7ad82c, 32'hbd296500} /* (14, 17, 1) {real, imag} */,
  {32'h3f13aa84, 32'h3f009eac} /* (14, 17, 0) {real, imag} */,
  {32'h3ee3880c, 32'h3ed57f48} /* (14, 16, 31) {real, imag} */,
  {32'h3e6f4290, 32'h3ebf4030} /* (14, 16, 30) {real, imag} */,
  {32'h3f11e964, 32'h3e3518e0} /* (14, 16, 29) {real, imag} */,
  {32'h3f608954, 32'hbe9304c0} /* (14, 16, 28) {real, imag} */,
  {32'h3fb68ebc, 32'hbe905210} /* (14, 16, 27) {real, imag} */,
  {32'h3f93b5c1, 32'h3dd99640} /* (14, 16, 26) {real, imag} */,
  {32'h3f05e5d7, 32'h3ded2d80} /* (14, 16, 25) {real, imag} */,
  {32'hbd994bf0, 32'h3eade9a0} /* (14, 16, 24) {real, imag} */,
  {32'hbe65b4a4, 32'h3edee680} /* (14, 16, 23) {real, imag} */,
  {32'h3f03be0c, 32'hbde82e80} /* (14, 16, 22) {real, imag} */,
  {32'h3ed501e8, 32'hbf2c1a84} /* (14, 16, 21) {real, imag} */,
  {32'hbe2ff178, 32'hbea6fdc0} /* (14, 16, 20) {real, imag} */,
  {32'h3f64d22d, 32'hbf233410} /* (14, 16, 19) {real, imag} */,
  {32'h3cf10cc0, 32'hbefe7020} /* (14, 16, 18) {real, imag} */,
  {32'hbf4101d0, 32'h3ea03240} /* (14, 16, 17) {real, imag} */,
  {32'hbf84b2cb, 32'h3df9de80} /* (14, 16, 16) {real, imag} */,
  {32'hbfb93280, 32'h3f991110} /* (14, 16, 15) {real, imag} */,
  {32'hbfe414ac, 32'h3eb5dc00} /* (14, 16, 14) {real, imag} */,
  {32'hbf71a592, 32'h3e809a50} /* (14, 16, 13) {real, imag} */,
  {32'hbf87f8b7, 32'hbf032838} /* (14, 16, 12) {real, imag} */,
  {32'h3e145a04, 32'hbf24b970} /* (14, 16, 11) {real, imag} */,
  {32'h3d0643a0, 32'hbf4ef214} /* (14, 16, 10) {real, imag} */,
  {32'h3f6c8b7c, 32'hbfb48670} /* (14, 16, 9) {real, imag} */,
  {32'h4001da3c, 32'hbf3e50a8} /* (14, 16, 8) {real, imag} */,
  {32'h3fb3a2e2, 32'hbf28efb8} /* (14, 16, 7) {real, imag} */,
  {32'h3f526c78, 32'hbe8b0770} /* (14, 16, 6) {real, imag} */,
  {32'h3e1d66ec, 32'hbdb46a00} /* (14, 16, 5) {real, imag} */,
  {32'h3ede16ec, 32'h3d55c600} /* (14, 16, 4) {real, imag} */,
  {32'h3f830925, 32'h3e4beec0} /* (14, 16, 3) {real, imag} */,
  {32'h3fd237df, 32'hbdff5400} /* (14, 16, 2) {real, imag} */,
  {32'h3fbee468, 32'hbf82ed00} /* (14, 16, 1) {real, imag} */,
  {32'h3f1e0d1e, 32'h3d1ad800} /* (14, 16, 0) {real, imag} */,
  {32'h3f8b96c4, 32'h3e591b80} /* (14, 15, 31) {real, imag} */,
  {32'h3f0ca140, 32'h3f0de050} /* (14, 15, 30) {real, imag} */,
  {32'h3f362d90, 32'h3f3e4950} /* (14, 15, 29) {real, imag} */,
  {32'h3ec90014, 32'h3edd6a20} /* (14, 15, 28) {real, imag} */,
  {32'h3e40a170, 32'hbeeef5d0} /* (14, 15, 27) {real, imag} */,
  {32'h3ecf2f3c, 32'hbf273db0} /* (14, 15, 26) {real, imag} */,
  {32'h3e46b250, 32'hbedf3c00} /* (14, 15, 25) {real, imag} */,
  {32'hbec698e0, 32'h3e574ee0} /* (14, 15, 24) {real, imag} */,
  {32'hbf350aba, 32'h3ecce330} /* (14, 15, 23) {real, imag} */,
  {32'hbf062c52, 32'h3f134450} /* (14, 15, 22) {real, imag} */,
  {32'hbe8f9020, 32'h3e8202dc} /* (14, 15, 21) {real, imag} */,
  {32'hbe952a14, 32'h3eb4f0a0} /* (14, 15, 20) {real, imag} */,
  {32'h3f1c2136, 32'hbe6038e0} /* (14, 15, 19) {real, imag} */,
  {32'hbf182292, 32'hbdce5340} /* (14, 15, 18) {real, imag} */,
  {32'hbf50fd82, 32'hbeeb2700} /* (14, 15, 17) {real, imag} */,
  {32'hbf56ba78, 32'hbee4d220} /* (14, 15, 16) {real, imag} */,
  {32'hbfa74087, 32'h3f3ac578} /* (14, 15, 15) {real, imag} */,
  {32'hbfed2385, 32'h3edb0ea0} /* (14, 15, 14) {real, imag} */,
  {32'hbfbaaa18, 32'h3e24b1c0} /* (14, 15, 13) {real, imag} */,
  {32'hbf4ebcdc, 32'hbe75eac0} /* (14, 15, 12) {real, imag} */,
  {32'h3e436ecc, 32'hbee61b60} /* (14, 15, 11) {real, imag} */,
  {32'h3d6a1500, 32'hbf8fae28} /* (14, 15, 10) {real, imag} */,
  {32'h3efd1110, 32'hbfe17664} /* (14, 15, 9) {real, imag} */,
  {32'h3f8ee368, 32'hbe8f9950} /* (14, 15, 8) {real, imag} */,
  {32'h3fcca86e, 32'hbf022ee0} /* (14, 15, 7) {real, imag} */,
  {32'h3ee0bd3c, 32'hbed56270} /* (14, 15, 6) {real, imag} */,
  {32'h3d5972f0, 32'hbdd41d80} /* (14, 15, 5) {real, imag} */,
  {32'h3f8167ce, 32'h3e367580} /* (14, 15, 4) {real, imag} */,
  {32'h3f5be158, 32'h3f131fd8} /* (14, 15, 3) {real, imag} */,
  {32'h3f8d5194, 32'hbc8fa400} /* (14, 15, 2) {real, imag} */,
  {32'h3f8c452e, 32'hbefe9090} /* (14, 15, 1) {real, imag} */,
  {32'h3f331603, 32'h3e30b1c0} /* (14, 15, 0) {real, imag} */,
  {32'h3e8417a8, 32'h3f111f80} /* (14, 14, 31) {real, imag} */,
  {32'hbe187e10, 32'hbee1d580} /* (14, 14, 30) {real, imag} */,
  {32'h3f61aeee, 32'hbf0e0ab0} /* (14, 14, 29) {real, imag} */,
  {32'h3f08e206, 32'hbeb29160} /* (14, 14, 28) {real, imag} */,
  {32'hbe17c5f0, 32'hbf01e368} /* (14, 14, 27) {real, imag} */,
  {32'h3eaf1548, 32'hbe522900} /* (14, 14, 26) {real, imag} */,
  {32'h3f377fb8, 32'hbda6cc40} /* (14, 14, 25) {real, imag} */,
  {32'h3e9bae4e, 32'hbdf6f6c0} /* (14, 14, 24) {real, imag} */,
  {32'hbe30e4ce, 32'hbe2aff60} /* (14, 14, 23) {real, imag} */,
  {32'h3e006b90, 32'hbc452000} /* (14, 14, 22) {real, imag} */,
  {32'h3b87ab00, 32'h3e287660} /* (14, 14, 21) {real, imag} */,
  {32'hbf0e9e1f, 32'h3f16a190} /* (14, 14, 20) {real, imag} */,
  {32'hbe1de160, 32'h3f805f7c} /* (14, 14, 19) {real, imag} */,
  {32'hbef89fa8, 32'h3ee9c0c0} /* (14, 14, 18) {real, imag} */,
  {32'hbf6a412a, 32'h3d882d80} /* (14, 14, 17) {real, imag} */,
  {32'hbecfd63d, 32'hbd43f700} /* (14, 14, 16) {real, imag} */,
  {32'hbd8391e8, 32'h3c76d200} /* (14, 14, 15) {real, imag} */,
  {32'hbf215798, 32'hbd0bfa00} /* (14, 14, 14) {real, imag} */,
  {32'hbd9a0e20, 32'hbd945980} /* (14, 14, 13) {real, imag} */,
  {32'h3e8abf54, 32'h3e9a6bb0} /* (14, 14, 12) {real, imag} */,
  {32'hbef018b0, 32'h3e5b6540} /* (14, 14, 11) {real, imag} */,
  {32'h3d973970, 32'hbf083c46} /* (14, 14, 10) {real, imag} */,
  {32'h3ee7e110, 32'hbf087f48} /* (14, 14, 9) {real, imag} */,
  {32'h3f21ea98, 32'h3e180580} /* (14, 14, 8) {real, imag} */,
  {32'h3fa6a27e, 32'h3e7c1700} /* (14, 14, 7) {real, imag} */,
  {32'h3f95bed2, 32'h3e253b20} /* (14, 14, 6) {real, imag} */,
  {32'h3f410e10, 32'h3e24c360} /* (14, 14, 5) {real, imag} */,
  {32'h3e94f6a4, 32'hbe647180} /* (14, 14, 4) {real, imag} */,
  {32'h3e6d9fd0, 32'hbe924ea0} /* (14, 14, 3) {real, imag} */,
  {32'h3f367bb4, 32'hbde0a400} /* (14, 14, 2) {real, imag} */,
  {32'h3f7bb75c, 32'h3f73d6d0} /* (14, 14, 1) {real, imag} */,
  {32'h3f6bdafc, 32'h3f7369d0} /* (14, 14, 0) {real, imag} */,
  {32'hbdec1b14, 32'h3e109c80} /* (14, 13, 31) {real, imag} */,
  {32'h3dfda2b0, 32'hbea6b110} /* (14, 13, 30) {real, imag} */,
  {32'h3f3cf31e, 32'hbf3af6f0} /* (14, 13, 29) {real, imag} */,
  {32'h3ec447e4, 32'hbf66ad60} /* (14, 13, 28) {real, imag} */,
  {32'h3f29275f, 32'hbe8475c0} /* (14, 13, 27) {real, imag} */,
  {32'h3f60ea5e, 32'hbe196900} /* (14, 13, 26) {real, imag} */,
  {32'h3f873e10, 32'hbf0363b0} /* (14, 13, 25) {real, imag} */,
  {32'h3fb234fa, 32'hbd26b780} /* (14, 13, 24) {real, imag} */,
  {32'h3f72c19b, 32'hbe26f560} /* (14, 13, 23) {real, imag} */,
  {32'h3fcb2879, 32'hbf0ffac0} /* (14, 13, 22) {real, imag} */,
  {32'h3ec1639c, 32'hbf4e0780} /* (14, 13, 21) {real, imag} */,
  {32'hbf72f776, 32'hbe34b220} /* (14, 13, 20) {real, imag} */,
  {32'hbdc57240, 32'h3f80b5b8} /* (14, 13, 19) {real, imag} */,
  {32'h3dcb6170, 32'h3f3ba920} /* (14, 13, 18) {real, imag} */,
  {32'hbe18ade0, 32'h3f473740} /* (14, 13, 17) {real, imag} */,
  {32'hbea6de88, 32'h3f3b3b18} /* (14, 13, 16) {real, imag} */,
  {32'hbe6152b0, 32'h3e8b5850} /* (14, 13, 15) {real, imag} */,
  {32'hbf0e7b9c, 32'h3e2ad5c0} /* (14, 13, 14) {real, imag} */,
  {32'hbf7438f6, 32'h3f376bc8} /* (14, 13, 13) {real, imag} */,
  {32'hbf95dbd9, 32'h3f410c10} /* (14, 13, 12) {real, imag} */,
  {32'hbf5299e4, 32'h3eebde80} /* (14, 13, 11) {real, imag} */,
  {32'hbd9b5678, 32'hbe660d28} /* (14, 13, 10) {real, imag} */,
  {32'hbe97eb18, 32'hbdfccd80} /* (14, 13, 9) {real, imag} */,
  {32'h3e42afa8, 32'hbea5cd60} /* (14, 13, 8) {real, imag} */,
  {32'h3fc48c07, 32'hbe8ff080} /* (14, 13, 7) {real, imag} */,
  {32'h3ff373e7, 32'h3e2ccbc0} /* (14, 13, 6) {real, imag} */,
  {32'h3f517039, 32'h3f499b78} /* (14, 13, 5) {real, imag} */,
  {32'h3e8d30ef, 32'h3f3bcc30} /* (14, 13, 4) {real, imag} */,
  {32'h3e4903d0, 32'h3f1f1058} /* (14, 13, 3) {real, imag} */,
  {32'h3f38f3e8, 32'h3f452190} /* (14, 13, 2) {real, imag} */,
  {32'h3f849c9d, 32'h3fb6e124} /* (14, 13, 1) {real, imag} */,
  {32'h3eb74e72, 32'h3f8424c8} /* (14, 13, 0) {real, imag} */,
  {32'h3eedc40f, 32'h3e54c550} /* (14, 12, 31) {real, imag} */,
  {32'h3f18de82, 32'h3e9df420} /* (14, 12, 30) {real, imag} */,
  {32'h3efcb8f8, 32'hbe8fb240} /* (14, 12, 29) {real, imag} */,
  {32'h3f67201c, 32'hbeda8c70} /* (14, 12, 28) {real, imag} */,
  {32'h3f94f100, 32'hbd3e9780} /* (14, 12, 27) {real, imag} */,
  {32'h3f5ee432, 32'h3e720e00} /* (14, 12, 26) {real, imag} */,
  {32'h3eff1e18, 32'hbe863dd0} /* (14, 12, 25) {real, imag} */,
  {32'h3e4795c0, 32'h3e9d2dd0} /* (14, 12, 24) {real, imag} */,
  {32'h3d3194a0, 32'h3e1dd920} /* (14, 12, 23) {real, imag} */,
  {32'h3e848440, 32'hbf2a1980} /* (14, 12, 22) {real, imag} */,
  {32'h3e8af8e4, 32'hbf3be740} /* (14, 12, 21) {real, imag} */,
  {32'hbf31025e, 32'hbe2a6900} /* (14, 12, 20) {real, imag} */,
  {32'hbed78120, 32'h3ee85580} /* (14, 12, 19) {real, imag} */,
  {32'hbecc6164, 32'h3ebbed00} /* (14, 12, 18) {real, imag} */,
  {32'hbf3419e0, 32'h3f95c864} /* (14, 12, 17) {real, imag} */,
  {32'hbf6b9e80, 32'h3f8430a0} /* (14, 12, 16) {real, imag} */,
  {32'hbea0e670, 32'h3da65300} /* (14, 12, 15) {real, imag} */,
  {32'hbf246dce, 32'h3ee8d870} /* (14, 12, 14) {real, imag} */,
  {32'hbf88dfb2, 32'h3f1ad0b8} /* (14, 12, 13) {real, imag} */,
  {32'hbfdb64a2, 32'h3f283770} /* (14, 12, 12) {real, imag} */,
  {32'hbfdeb992, 32'h3ed0a7a0} /* (14, 12, 11) {real, imag} */,
  {32'hbed7c3af, 32'h3e7a3800} /* (14, 12, 10) {real, imag} */,
  {32'h3ee315d4, 32'h3d83c240} /* (14, 12, 9) {real, imag} */,
  {32'h3fc14016, 32'hbe5a3940} /* (14, 12, 8) {real, imag} */,
  {32'h3fb5900a, 32'h3ef7a300} /* (14, 12, 7) {real, imag} */,
  {32'h3f9b73f2, 32'h3f116440} /* (14, 12, 6) {real, imag} */,
  {32'h3fa082ef, 32'h3f6c8320} /* (14, 12, 5) {real, imag} */,
  {32'h3f707d23, 32'h3fc137f4} /* (14, 12, 4) {real, imag} */,
  {32'h3efaab0c, 32'h3fca34e0} /* (14, 12, 3) {real, imag} */,
  {32'h3fa141ce, 32'h3f144db0} /* (14, 12, 2) {real, imag} */,
  {32'h3f9b703e, 32'h3dcaf280} /* (14, 12, 1) {real, imag} */,
  {32'h3f0c345d, 32'h3e4a7ac0} /* (14, 12, 0) {real, imag} */,
  {32'h3ebc4c68, 32'hbe23e840} /* (14, 11, 31) {real, imag} */,
  {32'h3ed860bd, 32'hbf28fc40} /* (14, 11, 30) {real, imag} */,
  {32'h3f72e278, 32'hbf050010} /* (14, 11, 29) {real, imag} */,
  {32'h4011fa0f, 32'h3e091ac0} /* (14, 11, 28) {real, imag} */,
  {32'h3faa50aa, 32'h3c0c8a00} /* (14, 11, 27) {real, imag} */,
  {32'hbe3fc614, 32'h3e0d6ec0} /* (14, 11, 26) {real, imag} */,
  {32'hbefd8ea0, 32'hbf30d1f8} /* (14, 11, 25) {real, imag} */,
  {32'hbe99a3be, 32'hbea61b80} /* (14, 11, 24) {real, imag} */,
  {32'hbf0c43f9, 32'h3ebcbcf0} /* (14, 11, 23) {real, imag} */,
  {32'hbebb5f8a, 32'hbcd39800} /* (14, 11, 22) {real, imag} */,
  {32'hbe37ab18, 32'hbf196544} /* (14, 11, 21) {real, imag} */,
  {32'hbe7d0ad8, 32'hbf3f6b10} /* (14, 11, 20) {real, imag} */,
  {32'hbe57b1cb, 32'hbdccad80} /* (14, 11, 19) {real, imag} */,
  {32'hbf78dce1, 32'h3de0a6c0} /* (14, 11, 18) {real, imag} */,
  {32'hbf830942, 32'h3f7359c8} /* (14, 11, 17) {real, imag} */,
  {32'hbefc0b0c, 32'h3f0644b0} /* (14, 11, 16) {real, imag} */,
  {32'h3e9ba9f8, 32'hbe971dd0} /* (14, 11, 15) {real, imag} */,
  {32'hbec25ef8, 32'h3d33e780} /* (14, 11, 14) {real, imag} */,
  {32'hbf09b0da, 32'h3f3fa9f8} /* (14, 11, 13) {real, imag} */,
  {32'hbf02f96e, 32'h3e877fa0} /* (14, 11, 12) {real, imag} */,
  {32'hbfcbed02, 32'hbe9f0bc8} /* (14, 11, 11) {real, imag} */,
  {32'hbf1acac7, 32'h3ea93b90} /* (14, 11, 10) {real, imag} */,
  {32'h3ee44a16, 32'h3ec17e40} /* (14, 11, 9) {real, imag} */,
  {32'h3f597fa7, 32'hbced0700} /* (14, 11, 8) {real, imag} */,
  {32'h3f4251a0, 32'h3e5280c0} /* (14, 11, 7) {real, imag} */,
  {32'h3fc29652, 32'h3ee29a70} /* (14, 11, 6) {real, imag} */,
  {32'h3fcc617d, 32'h3ef91548} /* (14, 11, 5) {real, imag} */,
  {32'h3f864a3a, 32'h3d0fa900} /* (14, 11, 4) {real, imag} */,
  {32'h3ecdcf32, 32'h3d905100} /* (14, 11, 3) {real, imag} */,
  {32'h3f9d03a8, 32'hbeb8e5b0} /* (14, 11, 2) {real, imag} */,
  {32'h3f36492e, 32'hbf08c9b0} /* (14, 11, 1) {real, imag} */,
  {32'h3f030e0d, 32'hbe1a3ea0} /* (14, 11, 0) {real, imag} */,
  {32'hbe331e8d, 32'h3e51cd70} /* (14, 10, 31) {real, imag} */,
  {32'hbe092c00, 32'hbe160a10} /* (14, 10, 30) {real, imag} */,
  {32'h3efc289c, 32'h3d83d980} /* (14, 10, 29) {real, imag} */,
  {32'h3e484c74, 32'h3f7bf720} /* (14, 10, 28) {real, imag} */,
  {32'hbf2762a4, 32'h3f0fb568} /* (14, 10, 27) {real, imag} */,
  {32'hbf612414, 32'hbf190ec4} /* (14, 10, 26) {real, imag} */,
  {32'hbf41918d, 32'hbf7c3f7c} /* (14, 10, 25) {real, imag} */,
  {32'hbe86cb98, 32'hbf44fbe8} /* (14, 10, 24) {real, imag} */,
  {32'hbf9fb85d, 32'hbe95f950} /* (14, 10, 23) {real, imag} */,
  {32'hbf816d8a, 32'h3f6b0ff0} /* (14, 10, 22) {real, imag} */,
  {32'hbecf519d, 32'h3eac2840} /* (14, 10, 21) {real, imag} */,
  {32'hbe25d8a2, 32'hbf651b94} /* (14, 10, 20) {real, imag} */,
  {32'h3f0798a0, 32'hbf326410} /* (14, 10, 19) {real, imag} */,
  {32'h3dc3ae50, 32'h3dd66700} /* (14, 10, 18) {real, imag} */,
  {32'h3e665ed0, 32'h3f2de91a} /* (14, 10, 17) {real, imag} */,
  {32'hbdaf0bd0, 32'hbdf75e80} /* (14, 10, 16) {real, imag} */,
  {32'h3f8a19e3, 32'hbe926190} /* (14, 10, 15) {real, imag} */,
  {32'h3e388b1b, 32'h3f0a1c58} /* (14, 10, 14) {real, imag} */,
  {32'hbeb2266f, 32'h3f9a12aa} /* (14, 10, 13) {real, imag} */,
  {32'hbe8ba1d2, 32'hbe3e0980} /* (14, 10, 12) {real, imag} */,
  {32'hbddb8de0, 32'hbe5494c0} /* (14, 10, 11) {real, imag} */,
  {32'hbf14a2a9, 32'h3d885c7c} /* (14, 10, 10) {real, imag} */,
  {32'hbf6c8744, 32'h3df110a0} /* (14, 10, 9) {real, imag} */,
  {32'hbf59787d, 32'hbf56c214} /* (14, 10, 8) {real, imag} */,
  {32'hbf064424, 32'hbdefabc0} /* (14, 10, 7) {real, imag} */,
  {32'h3e163060, 32'h3ead0dd0} /* (14, 10, 6) {real, imag} */,
  {32'hbf049155, 32'hbe389940} /* (14, 10, 5) {real, imag} */,
  {32'hbf8012e6, 32'hbf42dad8} /* (14, 10, 4) {real, imag} */,
  {32'hbe9028b0, 32'hbf3c373c} /* (14, 10, 3) {real, imag} */,
  {32'h3ecc7ebc, 32'hbf7557a0} /* (14, 10, 2) {real, imag} */,
  {32'hbf46b85c, 32'hbf8fde48} /* (14, 10, 1) {real, imag} */,
  {32'hbeada406, 32'hbe813af8} /* (14, 10, 0) {real, imag} */,
  {32'hbf11d8bc, 32'hbe95acc0} /* (14, 9, 31) {real, imag} */,
  {32'hbf3b0764, 32'h3f12fae8} /* (14, 9, 30) {real, imag} */,
  {32'hbf6a80e8, 32'h3f8d8e90} /* (14, 9, 29) {real, imag} */,
  {32'hbf8e933b, 32'h3f391b90} /* (14, 9, 28) {real, imag} */,
  {32'hbfa84a9e, 32'h3e937d20} /* (14, 9, 27) {real, imag} */,
  {32'hbf77094d, 32'hbf7a8690} /* (14, 9, 26) {real, imag} */,
  {32'hbf66a3f3, 32'hbfbee49c} /* (14, 9, 25) {real, imag} */,
  {32'hbf056c58, 32'hbfbc6b00} /* (14, 9, 24) {real, imag} */,
  {32'hbf4e0654, 32'h3ec573c0} /* (14, 9, 23) {real, imag} */,
  {32'hbfb66c11, 32'h3f6a9bc8} /* (14, 9, 22) {real, imag} */,
  {32'h3e6057a8, 32'hbf329840} /* (14, 9, 21) {real, imag} */,
  {32'h3f14234f, 32'hbf9da62a} /* (14, 9, 20) {real, imag} */,
  {32'h3f4968dc, 32'hbb937000} /* (14, 9, 19) {real, imag} */,
  {32'h3ec9cf54, 32'h3f9e22a4} /* (14, 9, 18) {real, imag} */,
  {32'h3da20850, 32'h3eaba7d0} /* (14, 9, 17) {real, imag} */,
  {32'h3c7f0900, 32'hbf034150} /* (14, 9, 16) {real, imag} */,
  {32'h3fa6bf10, 32'hbf9c1c50} /* (14, 9, 15) {real, imag} */,
  {32'h3f66d48a, 32'hbe66c420} /* (14, 9, 14) {real, imag} */,
  {32'h3f17668c, 32'h3efb6890} /* (14, 9, 13) {real, imag} */,
  {32'h3ec46eb0, 32'hbf35b0e0} /* (14, 9, 12) {real, imag} */,
  {32'h3f86317d, 32'hbf2c8660} /* (14, 9, 11) {real, imag} */,
  {32'h3af7df00, 32'hbcdafb80} /* (14, 9, 10) {real, imag} */,
  {32'hbfd994a4, 32'hbec7b200} /* (14, 9, 9) {real, imag} */,
  {32'hc00f4c7e, 32'hbf2d45f0} /* (14, 9, 8) {real, imag} */,
  {32'hbfb7ca1f, 32'h3e584840} /* (14, 9, 7) {real, imag} */,
  {32'hbf946a01, 32'h3f2f9750} /* (14, 9, 6) {real, imag} */,
  {32'hbfd2198f, 32'h3e5df140} /* (14, 9, 5) {real, imag} */,
  {32'hc002f816, 32'hbe356540} /* (14, 9, 4) {real, imag} */,
  {32'hbf0e8b9f, 32'hbf084c50} /* (14, 9, 3) {real, imag} */,
  {32'h3ea76303, 32'hbf8cce18} /* (14, 9, 2) {real, imag} */,
  {32'h3da89e90, 32'hbfd70278} /* (14, 9, 1) {real, imag} */,
  {32'hbeca5726, 32'hbf3f5870} /* (14, 9, 0) {real, imag} */,
  {32'hbf215224, 32'hbeb72c80} /* (14, 8, 31) {real, imag} */,
  {32'hbf97cf96, 32'h3f3516d8} /* (14, 8, 30) {real, imag} */,
  {32'hbfb7f406, 32'h3f2f31b8} /* (14, 8, 29) {real, imag} */,
  {32'hbf649b2e, 32'h3d87d980} /* (14, 8, 28) {real, imag} */,
  {32'hbf95e94a, 32'h3f10a340} /* (14, 8, 27) {real, imag} */,
  {32'hbf8a1b29, 32'hbf169b20} /* (14, 8, 26) {real, imag} */,
  {32'hbed53ea2, 32'hbf884814} /* (14, 8, 25) {real, imag} */,
  {32'hbd386870, 32'hbfb3a59c} /* (14, 8, 24) {real, imag} */,
  {32'hbdaf2e00, 32'hbe083c40} /* (14, 8, 23) {real, imag} */,
  {32'hbf116ba0, 32'h3ee3dc20} /* (14, 8, 22) {real, imag} */,
  {32'hbf12e51e, 32'hbec8dec0} /* (14, 8, 21) {real, imag} */,
  {32'h3f0bb8ba, 32'hbf060be8} /* (14, 8, 20) {real, imag} */,
  {32'h3fa682d0, 32'hbdd68680} /* (14, 8, 19) {real, imag} */,
  {32'h3f403398, 32'h3f59e300} /* (14, 8, 18) {real, imag} */,
  {32'h3e6efc50, 32'h3f015aa0} /* (14, 8, 17) {real, imag} */,
  {32'h3efed3c0, 32'h3d7f7100} /* (14, 8, 16) {real, imag} */,
  {32'h3fa3644e, 32'hbe272280} /* (14, 8, 15) {real, imag} */,
  {32'h3f6bebc4, 32'h3f01e1c0} /* (14, 8, 14) {real, imag} */,
  {32'h3f3219c3, 32'h3f2e2da0} /* (14, 8, 13) {real, imag} */,
  {32'h3f224808, 32'hbe5d5be0} /* (14, 8, 12) {real, imag} */,
  {32'h3fc8705c, 32'hbf331c88} /* (14, 8, 11) {real, imag} */,
  {32'h3ecece48, 32'hbd7b6800} /* (14, 8, 10) {real, imag} */,
  {32'hbfc7786a, 32'hbeb270e0} /* (14, 8, 9) {real, imag} */,
  {32'hbfae8f16, 32'hbe2a79e0} /* (14, 8, 8) {real, imag} */,
  {32'hbf468ffc, 32'h3cfff100} /* (14, 8, 7) {real, imag} */,
  {32'hbfbf3e68, 32'h3edc2250} /* (14, 8, 6) {real, imag} */,
  {32'hbf5ffb32, 32'h3e7ff2c0} /* (14, 8, 5) {real, imag} */,
  {32'hbfa9f729, 32'hbd406a00} /* (14, 8, 4) {real, imag} */,
  {32'hbf5d85cc, 32'h3e056c20} /* (14, 8, 3) {real, imag} */,
  {32'h3ed342f0, 32'hbed51aa0} /* (14, 8, 2) {real, imag} */,
  {32'hbe5fc940, 32'hbf94ce3c} /* (14, 8, 1) {real, imag} */,
  {32'hbfb3ae6f, 32'hbf2d224c} /* (14, 8, 0) {real, imag} */,
  {32'hbe88a400, 32'h3f131558} /* (14, 7, 31) {real, imag} */,
  {32'hbf3201f0, 32'h3f00a6b0} /* (14, 7, 30) {real, imag} */,
  {32'hbfc46779, 32'hbc49d000} /* (14, 7, 29) {real, imag} */,
  {32'hbf426395, 32'h3e1009a0} /* (14, 7, 28) {real, imag} */,
  {32'hbf267dee, 32'h3f0d8ed8} /* (14, 7, 27) {real, imag} */,
  {32'hbf19efb0, 32'hbe349700} /* (14, 7, 26) {real, imag} */,
  {32'hbefed7cc, 32'hbf21cec0} /* (14, 7, 25) {real, imag} */,
  {32'hbe8b26a0, 32'hbf59a8a0} /* (14, 7, 24) {real, imag} */,
  {32'hbe529328, 32'hbec71be0} /* (14, 7, 23) {real, imag} */,
  {32'hbda0cba0, 32'h3e3c2d60} /* (14, 7, 22) {real, imag} */,
  {32'hbe96b680, 32'h3f30e4d8} /* (14, 7, 21) {real, imag} */,
  {32'h3f177ce2, 32'h3ef291a0} /* (14, 7, 20) {real, imag} */,
  {32'h3f72cf9e, 32'hbd01af00} /* (14, 7, 19) {real, imag} */,
  {32'h3f26dc90, 32'hbec0eca0} /* (14, 7, 18) {real, imag} */,
  {32'h3eb07b48, 32'hbde71d80} /* (14, 7, 17) {real, imag} */,
  {32'h3f83d278, 32'h3db40680} /* (14, 7, 16) {real, imag} */,
  {32'h3fa23606, 32'h3f9174d8} /* (14, 7, 15) {real, imag} */,
  {32'h3f2d4ca8, 32'h3f0b0f40} /* (14, 7, 14) {real, imag} */,
  {32'h3eb47df8, 32'h3e12e860} /* (14, 7, 13) {real, imag} */,
  {32'h3e42e678, 32'h3f158480} /* (14, 7, 12) {real, imag} */,
  {32'h3f9308c0, 32'h3ec77760} /* (14, 7, 11) {real, imag} */,
  {32'hbdb34520, 32'h3eae6990} /* (14, 7, 10) {real, imag} */,
  {32'hbf29242c, 32'h3f3a3678} /* (14, 7, 9) {real, imag} */,
  {32'hbf4434a6, 32'hbd6c4580} /* (14, 7, 8) {real, imag} */,
  {32'hbf420311, 32'h3e791f60} /* (14, 7, 7) {real, imag} */,
  {32'hbfa481d9, 32'h3f259478} /* (14, 7, 6) {real, imag} */,
  {32'hbf0aa23e, 32'h3eee55c0} /* (14, 7, 5) {real, imag} */,
  {32'hbf6f8614, 32'hbeca20c0} /* (14, 7, 4) {real, imag} */,
  {32'hbebe6828, 32'hbe93a520} /* (14, 7, 3) {real, imag} */,
  {32'h3e067f90, 32'hbdeb8000} /* (14, 7, 2) {real, imag} */,
  {32'hbf8090f8, 32'hbf289910} /* (14, 7, 1) {real, imag} */,
  {32'hbf88da0c, 32'hbe8e1af0} /* (14, 7, 0) {real, imag} */,
  {32'hbf473c46, 32'h3eb46160} /* (14, 6, 31) {real, imag} */,
  {32'hbee4bbec, 32'h3eb9d4b0} /* (14, 6, 30) {real, imag} */,
  {32'hbf05bf5e, 32'hbedfa040} /* (14, 6, 29) {real, imag} */,
  {32'hbf292db7, 32'hbe9225e0} /* (14, 6, 28) {real, imag} */,
  {32'hbf0e774c, 32'hbee84200} /* (14, 6, 27) {real, imag} */,
  {32'hbef65320, 32'hbf23d598} /* (14, 6, 26) {real, imag} */,
  {32'hbed100a0, 32'hbf4d2660} /* (14, 6, 25) {real, imag} */,
  {32'hbe707530, 32'hbed53f40} /* (14, 6, 24) {real, imag} */,
  {32'hbe4c0500, 32'hbf5879b0} /* (14, 6, 23) {real, imag} */,
  {32'hbd704fc0, 32'hbf024638} /* (14, 6, 22) {real, imag} */,
  {32'hbe909738, 32'h3e713800} /* (14, 6, 21) {real, imag} */,
  {32'hbe817014, 32'hbdcd78a0} /* (14, 6, 20) {real, imag} */,
  {32'h3f13bc52, 32'hbe97b510} /* (14, 6, 19) {real, imag} */,
  {32'h3f824bec, 32'hbf992350} /* (14, 6, 18) {real, imag} */,
  {32'h3f7ac2fd, 32'hbe4e01a0} /* (14, 6, 17) {real, imag} */,
  {32'h3f62303a, 32'h3e1a0f00} /* (14, 6, 16) {real, imag} */,
  {32'h3eae0860, 32'h3e90e000} /* (14, 6, 15) {real, imag} */,
  {32'h3ed3a0f0, 32'hbdb22680} /* (14, 6, 14) {real, imag} */,
  {32'h3f381e70, 32'h3de21fc0} /* (14, 6, 13) {real, imag} */,
  {32'h3f4eacec, 32'h3f6ce8a8} /* (14, 6, 12) {real, imag} */,
  {32'h3f4c1cb0, 32'h3ec6ce50} /* (14, 6, 11) {real, imag} */,
  {32'h3d3dd9b0, 32'h3f1394e0} /* (14, 6, 10) {real, imag} */,
  {32'h3f4dfc56, 32'h3f2a7400} /* (14, 6, 9) {real, imag} */,
  {32'h3f56efbe, 32'hbe01a980} /* (14, 6, 8) {real, imag} */,
  {32'hbdbf8628, 32'h3f828c98} /* (14, 6, 7) {real, imag} */,
  {32'hbf6bbc48, 32'h3fef5548} /* (14, 6, 6) {real, imag} */,
  {32'hbf5783b4, 32'h3fa3a9e8} /* (14, 6, 5) {real, imag} */,
  {32'hbf9353f2, 32'hbecdd640} /* (14, 6, 4) {real, imag} */,
  {32'hbee3ba78, 32'hbf924764} /* (14, 6, 3) {real, imag} */,
  {32'hbe6dd000, 32'h3c906c00} /* (14, 6, 2) {real, imag} */,
  {32'h3da4bc80, 32'h3f3a93e8} /* (14, 6, 1) {real, imag} */,
  {32'hbdb78ba0, 32'h3ea44588} /* (14, 6, 0) {real, imag} */,
  {32'hbf432a44, 32'h3f322964} /* (14, 5, 31) {real, imag} */,
  {32'hbf081dc0, 32'h3f036d50} /* (14, 5, 30) {real, imag} */,
  {32'hbf4ba796, 32'hbeb41aa0} /* (14, 5, 29) {real, imag} */,
  {32'hbfa988e9, 32'hbf2ddd00} /* (14, 5, 28) {real, imag} */,
  {32'hbf980963, 32'hbfa5e7b8} /* (14, 5, 27) {real, imag} */,
  {32'hbf63674c, 32'hbf999c88} /* (14, 5, 26) {real, imag} */,
  {32'hbf0a40fa, 32'hbf70ebf0} /* (14, 5, 25) {real, imag} */,
  {32'hbf26ad62, 32'hbf447ab0} /* (14, 5, 24) {real, imag} */,
  {32'hbf5b663c, 32'hbf790de0} /* (14, 5, 23) {real, imag} */,
  {32'hbf07ee50, 32'hbdc3af00} /* (14, 5, 22) {real, imag} */,
  {32'hbf401143, 32'hbd7c8a80} /* (14, 5, 21) {real, imag} */,
  {32'hbf99f51a, 32'hbd9ab4c0} /* (14, 5, 20) {real, imag} */,
  {32'hbe95f652, 32'hbd7ce780} /* (14, 5, 19) {real, imag} */,
  {32'h3f236356, 32'hbe6ffe60} /* (14, 5, 18) {real, imag} */,
  {32'h3ef2c294, 32'h3e529020} /* (14, 5, 17) {real, imag} */,
  {32'hbb840040, 32'hbb2aa000} /* (14, 5, 16) {real, imag} */,
  {32'h3d4f2400, 32'hbe4b64a0} /* (14, 5, 15) {real, imag} */,
  {32'h3e88971c, 32'hbf6e9708} /* (14, 5, 14) {real, imag} */,
  {32'h3f3044b2, 32'h3ee83520} /* (14, 5, 13) {real, imag} */,
  {32'h3f292f80, 32'h3f26a5f0} /* (14, 5, 12) {real, imag} */,
  {32'h3ec5fc90, 32'hbdb29400} /* (14, 5, 11) {real, imag} */,
  {32'h3d7a3520, 32'hbecfa290} /* (14, 5, 10) {real, imag} */,
  {32'h3f1b1119, 32'hbe989130} /* (14, 5, 9) {real, imag} */,
  {32'h3fa8275f, 32'hbf042c54} /* (14, 5, 8) {real, imag} */,
  {32'h3f1e733b, 32'h3f511b88} /* (14, 5, 7) {real, imag} */,
  {32'h3ec11d49, 32'h3fb6d13d} /* (14, 5, 6) {real, imag} */,
  {32'hbde3e310, 32'h3f1da228} /* (14, 5, 5) {real, imag} */,
  {32'hbf874383, 32'h3eeb02e0} /* (14, 5, 4) {real, imag} */,
  {32'hbeac9132, 32'hbef19b80} /* (14, 5, 3) {real, imag} */,
  {32'hbe05f300, 32'h3e83e040} /* (14, 5, 2) {real, imag} */,
  {32'hbf480648, 32'h3f293060} /* (14, 5, 1) {real, imag} */,
  {32'hbed918c0, 32'h3eebe500} /* (14, 5, 0) {real, imag} */,
  {32'hbea299a8, 32'h3e961218} /* (14, 4, 31) {real, imag} */,
  {32'hbebeebc0, 32'hbf104380} /* (14, 4, 30) {real, imag} */,
  {32'hbee1a798, 32'hbf3071f0} /* (14, 4, 29) {real, imag} */,
  {32'hbf58b962, 32'hbf3febb0} /* (14, 4, 28) {real, imag} */,
  {32'hbf148d46, 32'hbf815d28} /* (14, 4, 27) {real, imag} */,
  {32'hbf555ad5, 32'hbf23dcc0} /* (14, 4, 26) {real, imag} */,
  {32'hbf592d0c, 32'hbe8bc3c0} /* (14, 4, 25) {real, imag} */,
  {32'hbf9abb86, 32'hbe86a240} /* (14, 4, 24) {real, imag} */,
  {32'hbe715378, 32'hbe810c00} /* (14, 4, 23) {real, imag} */,
  {32'hbec7a140, 32'hbe1d3840} /* (14, 4, 22) {real, imag} */,
  {32'hbf712a44, 32'hbe594f00} /* (14, 4, 21) {real, imag} */,
  {32'hbfbd6e28, 32'h3f9351e8} /* (14, 4, 20) {real, imag} */,
  {32'hbf417868, 32'h3fbaef54} /* (14, 4, 19) {real, imag} */,
  {32'hbd8e77c0, 32'h3f8bc860} /* (14, 4, 18) {real, imag} */,
  {32'hbe691360, 32'h3f70b020} /* (14, 4, 17) {real, imag} */,
  {32'hbf3dc18e, 32'h3e973860} /* (14, 4, 16) {real, imag} */,
  {32'h3e768790, 32'hbe87e9d8} /* (14, 4, 15) {real, imag} */,
  {32'h3f367492, 32'hbf8dafb8} /* (14, 4, 14) {real, imag} */,
  {32'h3e43fbac, 32'hbe8e9a80} /* (14, 4, 13) {real, imag} */,
  {32'h3e039f20, 32'hbd72de80} /* (14, 4, 12) {real, imag} */,
  {32'h3f1bccdc, 32'hbe948660} /* (14, 4, 11) {real, imag} */,
  {32'h3e760920, 32'hbe9328a0} /* (14, 4, 10) {real, imag} */,
  {32'hbc40ef80, 32'h3dd856c0} /* (14, 4, 9) {real, imag} */,
  {32'h3ea16b2c, 32'hbb21e000} /* (14, 4, 8) {real, imag} */,
  {32'h3fa37061, 32'hbd988b40} /* (14, 4, 7) {real, imag} */,
  {32'h3fdd3158, 32'h3ead0d00} /* (14, 4, 6) {real, imag} */,
  {32'h3ecc9c65, 32'h3ed2e348} /* (14, 4, 5) {real, imag} */,
  {32'hbf822fde, 32'h3f066ea8} /* (14, 4, 4) {real, imag} */,
  {32'hbf186628, 32'h3e53b500} /* (14, 4, 3) {real, imag} */,
  {32'hbf00d8e4, 32'hbdf64980} /* (14, 4, 2) {real, imag} */,
  {32'hbf5e09a8, 32'h3d1bcc00} /* (14, 4, 1) {real, imag} */,
  {32'hbef7da58, 32'h3d83ee20} /* (14, 4, 0) {real, imag} */,
  {32'hbf3b4f1e, 32'hbe4d1660} /* (14, 3, 31) {real, imag} */,
  {32'hbf27249c, 32'hbe259680} /* (14, 3, 30) {real, imag} */,
  {32'h3e68b470, 32'h3ecd8420} /* (14, 3, 29) {real, imag} */,
  {32'hbec32853, 32'h3e2febc0} /* (14, 3, 28) {real, imag} */,
  {32'h3e9b701c, 32'hbdd74d80} /* (14, 3, 27) {real, imag} */,
  {32'hbe45f8b8, 32'hbcd67a00} /* (14, 3, 26) {real, imag} */,
  {32'hbf547da8, 32'h3e28dce0} /* (14, 3, 25) {real, imag} */,
  {32'hbfae719c, 32'h3f5a7b40} /* (14, 3, 24) {real, imag} */,
  {32'hbe9f51f4, 32'h3ea0e310} /* (14, 3, 23) {real, imag} */,
  {32'hbf010888, 32'hbe8d3040} /* (14, 3, 22) {real, imag} */,
  {32'hbe80652c, 32'hbecbef50} /* (14, 3, 21) {real, imag} */,
  {32'hbf20566c, 32'hbd8122c0} /* (14, 3, 20) {real, imag} */,
  {32'hbf3cc404, 32'h3f9620a0} /* (14, 3, 19) {real, imag} */,
  {32'hbe2e7ee0, 32'h3f90c898} /* (14, 3, 18) {real, imag} */,
  {32'hbf024608, 32'h3ef6c6c0} /* (14, 3, 17) {real, imag} */,
  {32'hbf9afd14, 32'hbe9c9b90} /* (14, 3, 16) {real, imag} */,
  {32'hbe15904c, 32'hbe8cfbe8} /* (14, 3, 15) {real, imag} */,
  {32'h3fa707a2, 32'hbf0ab7e8} /* (14, 3, 14) {real, imag} */,
  {32'h3eae3524, 32'hbf1e86a0} /* (14, 3, 13) {real, imag} */,
  {32'h3c2ed180, 32'hbe97ce40} /* (14, 3, 12) {real, imag} */,
  {32'h3ed1e888, 32'hbf8601c8} /* (14, 3, 11) {real, imag} */,
  {32'h3ae9f800, 32'hbebe1080} /* (14, 3, 10) {real, imag} */,
  {32'hbdca3530, 32'h3dcba380} /* (14, 3, 9) {real, imag} */,
  {32'hbe87da70, 32'h3e7dcf40} /* (14, 3, 8) {real, imag} */,
  {32'h3edfe940, 32'h3ecd4bc0} /* (14, 3, 7) {real, imag} */,
  {32'h3fad27ff, 32'h3f8b04e8} /* (14, 3, 6) {real, imag} */,
  {32'h3f1fbfee, 32'h3ef10f04} /* (14, 3, 5) {real, imag} */,
  {32'hbf3f50e6, 32'hbe9b9890} /* (14, 3, 4) {real, imag} */,
  {32'hbf55f488, 32'hbf8c1d68} /* (14, 3, 3) {real, imag} */,
  {32'hbe60ba68, 32'hbfcc69f8} /* (14, 3, 2) {real, imag} */,
  {32'hbeaecb80, 32'hbf112340} /* (14, 3, 1) {real, imag} */,
  {32'hbeed84b4, 32'h3e5611c0} /* (14, 3, 0) {real, imag} */,
  {32'hbe570e5c, 32'hbdf18c80} /* (14, 2, 31) {real, imag} */,
  {32'hbcc6ed80, 32'h3ce28400} /* (14, 2, 30) {real, imag} */,
  {32'h3c089800, 32'h3f796030} /* (14, 2, 29) {real, imag} */,
  {32'hbf71c5a8, 32'h3f65a628} /* (14, 2, 28) {real, imag} */,
  {32'hbf8399ca, 32'h3ea880a0} /* (14, 2, 27) {real, imag} */,
  {32'hbf4a0863, 32'h3da12140} /* (14, 2, 26) {real, imag} */,
  {32'hbf421fbc, 32'h3e4dc3a0} /* (14, 2, 25) {real, imag} */,
  {32'hbf9acf68, 32'h3e9d5ec0} /* (14, 2, 24) {real, imag} */,
  {32'hbf8a3f0a, 32'h3e56b040} /* (14, 2, 23) {real, imag} */,
  {32'hbfa103b4, 32'h3f66dd60} /* (14, 2, 22) {real, imag} */,
  {32'hbf46b0ea, 32'h3e979100} /* (14, 2, 21) {real, imag} */,
  {32'hbf753f00, 32'hbf2b6e10} /* (14, 2, 20) {real, imag} */,
  {32'hbf00e1e8, 32'h3e4b03c0} /* (14, 2, 19) {real, imag} */,
  {32'h3ef49580, 32'h3f5ce078} /* (14, 2, 18) {real, imag} */,
  {32'hbe03ca90, 32'h3f8850fc} /* (14, 2, 17) {real, imag} */,
  {32'hbf9f5e01, 32'h3e999210} /* (14, 2, 16) {real, imag} */,
  {32'h3bb23a00, 32'h3f147598} /* (14, 2, 15) {real, imag} */,
  {32'h3fcd6cf4, 32'h3d11c980} /* (14, 2, 14) {real, imag} */,
  {32'h3f42b08a, 32'h3e6791c0} /* (14, 2, 13) {real, imag} */,
  {32'h3f28d25a, 32'h3ebac600} /* (14, 2, 12) {real, imag} */,
  {32'h3f54e7d6, 32'hbf81e1e8} /* (14, 2, 11) {real, imag} */,
  {32'h3eb55af8, 32'hbee39c50} /* (14, 2, 10) {real, imag} */,
  {32'h3e8b8d50, 32'h3e8f00f0} /* (14, 2, 9) {real, imag} */,
  {32'h3eab63e0, 32'h3f21ce58} /* (14, 2, 8) {real, imag} */,
  {32'h3ea6e950, 32'h3ee76d80} /* (14, 2, 7) {real, imag} */,
  {32'h3f17fd14, 32'h3ee1c220} /* (14, 2, 6) {real, imag} */,
  {32'hbf58e496, 32'h3f58c6e9} /* (14, 2, 5) {real, imag} */,
  {32'hbf102578, 32'hbeb309a0} /* (14, 2, 4) {real, imag} */,
  {32'hbf378c91, 32'hbfc2f348} /* (14, 2, 3) {real, imag} */,
  {32'hbeb58770, 32'hbeff1aa0} /* (14, 2, 2) {real, imag} */,
  {32'h3eabe5f0, 32'hbe11f1e0} /* (14, 2, 1) {real, imag} */,
  {32'hbe0806d8, 32'h3e81ee88} /* (14, 2, 0) {real, imag} */,
  {32'h3e9df970, 32'h3e02bdf0} /* (14, 1, 31) {real, imag} */,
  {32'h3e611310, 32'h3e28b740} /* (14, 1, 30) {real, imag} */,
  {32'h3e74d9d0, 32'h3f418878} /* (14, 1, 29) {real, imag} */,
  {32'hbf4b4386, 32'h3f57ab50} /* (14, 1, 28) {real, imag} */,
  {32'hbfbef6f5, 32'h3f98b7c8} /* (14, 1, 27) {real, imag} */,
  {32'hbf7a24b1, 32'h3f591ad0} /* (14, 1, 26) {real, imag} */,
  {32'hbe9a0e98, 32'h3ea9e100} /* (14, 1, 25) {real, imag} */,
  {32'hbf836eaf, 32'hbeca6770} /* (14, 1, 24) {real, imag} */,
  {32'hbf4ca9be, 32'h3e76b140} /* (14, 1, 23) {real, imag} */,
  {32'hbeeea0ac, 32'h3fa48b6c} /* (14, 1, 22) {real, imag} */,
  {32'hbf0c4477, 32'h3f6d4d90} /* (14, 1, 21) {real, imag} */,
  {32'hbf68a752, 32'h3e9196b0} /* (14, 1, 20) {real, imag} */,
  {32'h3eae3578, 32'h3d430c00} /* (14, 1, 19) {real, imag} */,
  {32'h3f9feff0, 32'h3e5e6fc0} /* (14, 1, 18) {real, imag} */,
  {32'h3f27d180, 32'h3eeede40} /* (14, 1, 17) {real, imag} */,
  {32'hbeb20d56, 32'h3f200538} /* (14, 1, 16) {real, imag} */,
  {32'h3f1eff62, 32'h3f8508ac} /* (14, 1, 15) {real, imag} */,
  {32'h3f86825a, 32'h3f733178} /* (14, 1, 14) {real, imag} */,
  {32'h3ea78fc8, 32'h3f57b9b0} /* (14, 1, 13) {real, imag} */,
  {32'h3f7dfce0, 32'hbef497d0} /* (14, 1, 12) {real, imag} */,
  {32'h3e9f8b80, 32'hbfbfa868} /* (14, 1, 11) {real, imag} */,
  {32'h3eeff43c, 32'hbe6df100} /* (14, 1, 10) {real, imag} */,
  {32'h3f29fa98, 32'h3f1672c0} /* (14, 1, 9) {real, imag} */,
  {32'h3eca1ed4, 32'h3c03f000} /* (14, 1, 8) {real, imag} */,
  {32'h3eb018a8, 32'hbe4a9f00} /* (14, 1, 7) {real, imag} */,
  {32'h3fc2cb1f, 32'h3e456540} /* (14, 1, 6) {real, imag} */,
  {32'h3d826a08, 32'h3f23baf9} /* (14, 1, 5) {real, imag} */,
  {32'h3e091c00, 32'hbf56fc78} /* (14, 1, 4) {real, imag} */,
  {32'hbe46ffb0, 32'hbf019f30} /* (14, 1, 3) {real, imag} */,
  {32'hbe83433c, 32'h3f2c9cd8} /* (14, 1, 2) {real, imag} */,
  {32'h3f085270, 32'h3f6d09d0} /* (14, 1, 1) {real, imag} */,
  {32'h3ef4c168, 32'h3ed16760} /* (14, 1, 0) {real, imag} */,
  {32'h3ee3e2a0, 32'h3eb1e70c} /* (14, 0, 31) {real, imag} */,
  {32'hbe119240, 32'h3e6b9c70} /* (14, 0, 30) {real, imag} */,
  {32'hbec821a4, 32'h3d970320} /* (14, 0, 29) {real, imag} */,
  {32'hbec90634, 32'h3dc568c0} /* (14, 0, 28) {real, imag} */,
  {32'hbf5316d6, 32'h3f4b118c} /* (14, 0, 27) {real, imag} */,
  {32'hbec46a6e, 32'h3ec30010} /* (14, 0, 26) {real, imag} */,
  {32'hbde4cb30, 32'h3dd2a380} /* (14, 0, 25) {real, imag} */,
  {32'hbf6ae3fc, 32'hbc33d900} /* (14, 0, 24) {real, imag} */,
  {32'hbf0bed7a, 32'h3dc8cac0} /* (14, 0, 23) {real, imag} */,
  {32'hbddf77b0, 32'h3eaa1540} /* (14, 0, 22) {real, imag} */,
  {32'hbec3900a, 32'h3eb17460} /* (14, 0, 21) {real, imag} */,
  {32'hbede7c46, 32'h3ea3bec0} /* (14, 0, 20) {real, imag} */,
  {32'h3e710768, 32'h3eae2098} /* (14, 0, 19) {real, imag} */,
  {32'h3e531960, 32'h3eeb0b90} /* (14, 0, 18) {real, imag} */,
  {32'hbe1c096c, 32'h3e96b160} /* (14, 0, 17) {real, imag} */,
  {32'h3e2da850, 32'h3ed54a24} /* (14, 0, 16) {real, imag} */,
  {32'h3f517eba, 32'h3f266d20} /* (14, 0, 15) {real, imag} */,
  {32'h3ee4a9ae, 32'h3f307270} /* (14, 0, 14) {real, imag} */,
  {32'h3ec8c67e, 32'h3e9dcca0} /* (14, 0, 13) {real, imag} */,
  {32'h3eaf07a0, 32'hbe4d4e00} /* (14, 0, 12) {real, imag} */,
  {32'hbe14fbe8, 32'hbf4ac70c} /* (14, 0, 11) {real, imag} */,
  {32'h3f1572fb, 32'hbf15ee60} /* (14, 0, 10) {real, imag} */,
  {32'h3e08f010, 32'hbd1cc140} /* (14, 0, 9) {real, imag} */,
  {32'hbe3e11f8, 32'hbe2f5e60} /* (14, 0, 8) {real, imag} */,
  {32'h3e3bcf00, 32'h3dd05d00} /* (14, 0, 7) {real, imag} */,
  {32'h3f96357f, 32'h3e673d60} /* (14, 0, 6) {real, imag} */,
  {32'h3e0122c6, 32'h3e9d1076} /* (14, 0, 5) {real, imag} */,
  {32'hbee4d374, 32'hbe7d2e90} /* (14, 0, 4) {real, imag} */,
  {32'hbed26a28, 32'h3e9f80f8} /* (14, 0, 3) {real, imag} */,
  {32'hbf12d10d, 32'h3f1efa4c} /* (14, 0, 2) {real, imag} */,
  {32'hbe40f47c, 32'h3ebc4100} /* (14, 0, 1) {real, imag} */,
  {32'h3e980288, 32'h3e058140} /* (14, 0, 0) {real, imag} */,
  {32'h3e288860, 32'hbecfdf3e} /* (13, 31, 31) {real, imag} */,
  {32'h3f4ae69f, 32'hbf3215ed} /* (13, 31, 30) {real, imag} */,
  {32'h3da954a8, 32'h3e783818} /* (13, 31, 29) {real, imag} */,
  {32'hbc2d4300, 32'hbc569780} /* (13, 31, 28) {real, imag} */,
  {32'hbe6bebb0, 32'hbf3026ec} /* (13, 31, 27) {real, imag} */,
  {32'hbf1cd991, 32'hbe7029f8} /* (13, 31, 26) {real, imag} */,
  {32'hbea47ac8, 32'hbe67ed60} /* (13, 31, 25) {real, imag} */,
  {32'hbf206883, 32'h3e2e6fc0} /* (13, 31, 24) {real, imag} */,
  {32'h3eae0bfe, 32'h3ee3adac} /* (13, 31, 23) {real, imag} */,
  {32'h3f6cf37a, 32'hbbfdb000} /* (13, 31, 22) {real, imag} */,
  {32'h3db02fe0, 32'hbf0a2ec2} /* (13, 31, 21) {real, imag} */,
  {32'h3dcebf90, 32'hbddf3bf0} /* (13, 31, 20) {real, imag} */,
  {32'hbd74b18c, 32'h3d5c9b60} /* (13, 31, 19) {real, imag} */,
  {32'h3eaf3a10, 32'hbe5d45fc} /* (13, 31, 18) {real, imag} */,
  {32'h3f5700c8, 32'h3f1ea2ed} /* (13, 31, 17) {real, imag} */,
  {32'h3f01b799, 32'h3f86901e} /* (13, 31, 16) {real, imag} */,
  {32'h3f1891f5, 32'h3f352eca} /* (13, 31, 15) {real, imag} */,
  {32'hbae76800, 32'hbe9c3ae0} /* (13, 31, 14) {real, imag} */,
  {32'hbf46bb72, 32'h3da075a0} /* (13, 31, 13) {real, imag} */,
  {32'hbf3cfaeb, 32'h3d34c1c0} /* (13, 31, 12) {real, imag} */,
  {32'hbeb4d99b, 32'hbefdb714} /* (13, 31, 11) {real, imag} */,
  {32'hbe19a4b0, 32'hbf6add80} /* (13, 31, 10) {real, imag} */,
  {32'h3ea278e8, 32'hbe2076f0} /* (13, 31, 9) {real, imag} */,
  {32'h3f1581a6, 32'h3eda184c} /* (13, 31, 8) {real, imag} */,
  {32'h3f214e0a, 32'h3e204f28} /* (13, 31, 7) {real, imag} */,
  {32'h3f371758, 32'hbef0d4ec} /* (13, 31, 6) {real, imag} */,
  {32'hbefac8ea, 32'hbf610355} /* (13, 31, 5) {real, imag} */,
  {32'hbf70dc12, 32'hbf32e1f0} /* (13, 31, 4) {real, imag} */,
  {32'hbed17aa0, 32'h3f0419be} /* (13, 31, 3) {real, imag} */,
  {32'hbe2d986c, 32'h3e435cb8} /* (13, 31, 2) {real, imag} */,
  {32'h3e588610, 32'hbe8520e0} /* (13, 31, 1) {real, imag} */,
  {32'hbec62546, 32'hbca5a200} /* (13, 31, 0) {real, imag} */,
  {32'hbe3bab40, 32'hbf0c2d20} /* (13, 30, 31) {real, imag} */,
  {32'h3f194366, 32'hbf0b4d5c} /* (13, 30, 30) {real, imag} */,
  {32'hbe5d4208, 32'h3f447a84} /* (13, 30, 29) {real, imag} */,
  {32'h3e1a1af0, 32'h3f14fdc8} /* (13, 30, 28) {real, imag} */,
  {32'h3e59df80, 32'h3f33666c} /* (13, 30, 27) {real, imag} */,
  {32'hbf61c235, 32'h3ea50d4c} /* (13, 30, 26) {real, imag} */,
  {32'hbfb1da41, 32'hbeab5600} /* (13, 30, 25) {real, imag} */,
  {32'hc00d09cc, 32'h3f305e34} /* (13, 30, 24) {real, imag} */,
  {32'hbdfd7b70, 32'h3f455ed8} /* (13, 30, 23) {real, imag} */,
  {32'h3f55ef43, 32'hbf2f7f18} /* (13, 30, 22) {real, imag} */,
  {32'h3de19a2e, 32'hbec979f8} /* (13, 30, 21) {real, imag} */,
  {32'h3e8d1448, 32'h3e0ade80} /* (13, 30, 20) {real, imag} */,
  {32'hbe0dca88, 32'h3e2b7200} /* (13, 30, 19) {real, imag} */,
  {32'h3efeb474, 32'hbec9a8c8} /* (13, 30, 18) {real, imag} */,
  {32'h3fe525d4, 32'h3e97e370} /* (13, 30, 17) {real, imag} */,
  {32'h3f7020f4, 32'h3ec23f10} /* (13, 30, 16) {real, imag} */,
  {32'h3f8e6b4c, 32'hbe3aad30} /* (13, 30, 15) {real, imag} */,
  {32'h3f5af094, 32'hbd01c840} /* (13, 30, 14) {real, imag} */,
  {32'hbe8ae272, 32'h3ea66eb0} /* (13, 30, 13) {real, imag} */,
  {32'hbf66d3c3, 32'hbe9e7f38} /* (13, 30, 12) {real, imag} */,
  {32'hbf928df4, 32'hbf90eb22} /* (13, 30, 11) {real, imag} */,
  {32'hbfbb8f3c, 32'hbf56bccc} /* (13, 30, 10) {real, imag} */,
  {32'h3f4c72ee, 32'h3d88a220} /* (13, 30, 9) {real, imag} */,
  {32'h3fe415fa, 32'h3e619330} /* (13, 30, 8) {real, imag} */,
  {32'h3ee0a639, 32'hbe7f5610} /* (13, 30, 7) {real, imag} */,
  {32'hbf0018e8, 32'hbed5918c} /* (13, 30, 6) {real, imag} */,
  {32'hbf9188dd, 32'hbfa6baa1} /* (13, 30, 5) {real, imag} */,
  {32'hbf871a60, 32'h3c930c00} /* (13, 30, 4) {real, imag} */,
  {32'h3c4434c0, 32'h3f62ae98} /* (13, 30, 3) {real, imag} */,
  {32'h3f0e6eef, 32'hbf12c110} /* (13, 30, 2) {real, imag} */,
  {32'h3fb4e40e, 32'hbf86a0e4} /* (13, 30, 1) {real, imag} */,
  {32'h3ef3d9e4, 32'hbdfa06b0} /* (13, 30, 0) {real, imag} */,
  {32'hbe80a7e0, 32'h3d8a8ce0} /* (13, 29, 31) {real, imag} */,
  {32'h3e0d5640, 32'h3c1ffd00} /* (13, 29, 30) {real, imag} */,
  {32'hbf15aede, 32'hbec4d580} /* (13, 29, 29) {real, imag} */,
  {32'hbe901c00, 32'h3e8065f8} /* (13, 29, 28) {real, imag} */,
  {32'hbe0bd620, 32'h3f8cec3c} /* (13, 29, 27) {real, imag} */,
  {32'hbfa108d0, 32'h3ef4ce68} /* (13, 29, 26) {real, imag} */,
  {32'hbf8c50d7, 32'h3f16de5c} /* (13, 29, 25) {real, imag} */,
  {32'hbf55ad63, 32'h3e9338f0} /* (13, 29, 24) {real, imag} */,
  {32'h3e0a440e, 32'hbdbf20e0} /* (13, 29, 23) {real, imag} */,
  {32'hbf06cc6e, 32'hbf8d5f42} /* (13, 29, 22) {real, imag} */,
  {32'hbf01074e, 32'h3ea4faa4} /* (13, 29, 21) {real, imag} */,
  {32'hbf207a06, 32'h3f7b97c0} /* (13, 29, 20) {real, imag} */,
  {32'hbf2642a2, 32'h3f7b6eac} /* (13, 29, 19) {real, imag} */,
  {32'hbec2f8a8, 32'h3e7526c0} /* (13, 29, 18) {real, imag} */,
  {32'h3f232268, 32'h3e9aec20} /* (13, 29, 17) {real, imag} */,
  {32'h3ef5827a, 32'h3f03d2f8} /* (13, 29, 16) {real, imag} */,
  {32'h3f221197, 32'hbf243e14} /* (13, 29, 15) {real, imag} */,
  {32'h3f1140d0, 32'hbeaa6e90} /* (13, 29, 14) {real, imag} */,
  {32'h3f11e119, 32'h3d494180} /* (13, 29, 13) {real, imag} */,
  {32'h3e690c8e, 32'hbf37d574} /* (13, 29, 12) {real, imag} */,
  {32'hbf06a49e, 32'hbf83077a} /* (13, 29, 11) {real, imag} */,
  {32'hbf8f1f92, 32'hbf5ffa98} /* (13, 29, 10) {real, imag} */,
  {32'h3e82c5dc, 32'hbeeb4ba0} /* (13, 29, 9) {real, imag} */,
  {32'h3f7ebfe1, 32'hbd392a80} /* (13, 29, 8) {real, imag} */,
  {32'h3f2ee626, 32'h3e0d60c0} /* (13, 29, 7) {real, imag} */,
  {32'hbeff8e90, 32'h3e5ec508} /* (13, 29, 6) {real, imag} */,
  {32'hbd952ca0, 32'hbe92609c} /* (13, 29, 5) {real, imag} */,
  {32'h3f19c554, 32'h3f3da9dc} /* (13, 29, 4) {real, imag} */,
  {32'h3fc6bb35, 32'h3f460268} /* (13, 29, 3) {real, imag} */,
  {32'h3f03a9d5, 32'hbf8b51cc} /* (13, 29, 2) {real, imag} */,
  {32'h3f7043a8, 32'hbfa3aecc} /* (13, 29, 1) {real, imag} */,
  {32'h3f2a2c9b, 32'hbedc9edc} /* (13, 29, 0) {real, imag} */,
  {32'h3e7df464, 32'h3eac1354} /* (13, 28, 31) {real, imag} */,
  {32'h3e9f38f4, 32'h3d5e94c0} /* (13, 28, 30) {real, imag} */,
  {32'h3eaaaa57, 32'hbf1ead7c} /* (13, 28, 29) {real, imag} */,
  {32'hbebecd58, 32'h3e246be8} /* (13, 28, 28) {real, imag} */,
  {32'hbe0bab00, 32'h3e8d1e78} /* (13, 28, 27) {real, imag} */,
  {32'h3e1bf8ac, 32'hbf811f54} /* (13, 28, 26) {real, imag} */,
  {32'h3e0d2528, 32'h3d1eac80} /* (13, 28, 25) {real, imag} */,
  {32'h3eacaf5e, 32'hbe2688c0} /* (13, 28, 24) {real, imag} */,
  {32'hbed0952e, 32'hbf250df6} /* (13, 28, 23) {real, imag} */,
  {32'hbfe15730, 32'hbf3e9bdc} /* (13, 28, 22) {real, imag} */,
  {32'hbf4eed00, 32'h3f28e2d8} /* (13, 28, 21) {real, imag} */,
  {32'h3daf9e10, 32'h3fe6e0d8} /* (13, 28, 20) {real, imag} */,
  {32'hbca43700, 32'h3fd05240} /* (13, 28, 19) {real, imag} */,
  {32'h3dfe4730, 32'h3f1674b8} /* (13, 28, 18) {real, imag} */,
  {32'h3f3a72f6, 32'h3ecdf760} /* (13, 28, 17) {real, imag} */,
  {32'h3f8e7b91, 32'h3f10c09c} /* (13, 28, 16) {real, imag} */,
  {32'h3fa7506e, 32'hbeed5578} /* (13, 28, 15) {real, imag} */,
  {32'h3efe019c, 32'hbb2ac400} /* (13, 28, 14) {real, imag} */,
  {32'h3e8571a2, 32'h3dff9ae0} /* (13, 28, 13) {real, imag} */,
  {32'h3e9482ca, 32'hbf6bf748} /* (13, 28, 12) {real, imag} */,
  {32'h3eefddfd, 32'hbf2e6f78} /* (13, 28, 11) {real, imag} */,
  {32'h3e89a190, 32'hbf317f9a} /* (13, 28, 10) {real, imag} */,
  {32'h3ec11658, 32'hbf1f300c} /* (13, 28, 9) {real, imag} */,
  {32'hbf19eb5c, 32'h3d838600} /* (13, 28, 8) {real, imag} */,
  {32'h3c844780, 32'h3f784f18} /* (13, 28, 7) {real, imag} */,
  {32'hbddd3688, 32'h3f2565cc} /* (13, 28, 6) {real, imag} */,
  {32'hbea3df98, 32'h3e9d40b8} /* (13, 28, 5) {real, imag} */,
  {32'h3e55b69c, 32'hbed61600} /* (13, 28, 4) {real, imag} */,
  {32'h3ea755cc, 32'hbe1e3f60} /* (13, 28, 3) {real, imag} */,
  {32'hbf083b55, 32'hbf444f30} /* (13, 28, 2) {real, imag} */,
  {32'h3e6a06a0, 32'hbe6de030} /* (13, 28, 1) {real, imag} */,
  {32'h3f232169, 32'h3e69bdea} /* (13, 28, 0) {real, imag} */,
  {32'h3e899f90, 32'hbf2aa406} /* (13, 27, 31) {real, imag} */,
  {32'h3f5f7513, 32'hbe2d4010} /* (13, 27, 30) {real, imag} */,
  {32'h3fb29bb6, 32'h3ece7470} /* (13, 27, 29) {real, imag} */,
  {32'h3ea1109c, 32'h3f8dcd28} /* (13, 27, 28) {real, imag} */,
  {32'h3ed36adc, 32'h3f3fee74} /* (13, 27, 27) {real, imag} */,
  {32'h3f22d300, 32'hbf81a658} /* (13, 27, 26) {real, imag} */,
  {32'h3d8df830, 32'hbefc1bc0} /* (13, 27, 25) {real, imag} */,
  {32'hbece6e1e, 32'hbe248280} /* (13, 27, 24) {real, imag} */,
  {32'hbfc8637c, 32'hbf1364a0} /* (13, 27, 23) {real, imag} */,
  {32'hbfce9203, 32'hbed0e640} /* (13, 27, 22) {real, imag} */,
  {32'hbf0c7ff8, 32'hbe910dc0} /* (13, 27, 21) {real, imag} */,
  {32'hbd8409c0, 32'h3dbe0620} /* (13, 27, 20) {real, imag} */,
  {32'hbebcc13c, 32'h3d3c0e00} /* (13, 27, 19) {real, imag} */,
  {32'h3eae25b2, 32'h3e2328c0} /* (13, 27, 18) {real, imag} */,
  {32'h3f16c676, 32'h3f8721eb} /* (13, 27, 17) {real, imag} */,
  {32'h3ea1cd8c, 32'h3f5fc56c} /* (13, 27, 16) {real, imag} */,
  {32'hbddb0680, 32'h3f2974cc} /* (13, 27, 15) {real, imag} */,
  {32'hbcdd7de0, 32'h3eb73d28} /* (13, 27, 14) {real, imag} */,
  {32'h3f1214bd, 32'h3f24cb20} /* (13, 27, 13) {real, imag} */,
  {32'h3e4e4658, 32'h3e159980} /* (13, 27, 12) {real, imag} */,
  {32'h3f266139, 32'hbf24a06c} /* (13, 27, 11) {real, imag} */,
  {32'h3f1dee1a, 32'hbf7fd4f0} /* (13, 27, 10) {real, imag} */,
  {32'h3f90b571, 32'hbf87341c} /* (13, 27, 9) {real, imag} */,
  {32'hbf10e390, 32'hbe675660} /* (13, 27, 8) {real, imag} */,
  {32'hbf836196, 32'h3ea6fed8} /* (13, 27, 7) {real, imag} */,
  {32'hbf0f670c, 32'h3f634337} /* (13, 27, 6) {real, imag} */,
  {32'hbf33c3ac, 32'h3ef654e0} /* (13, 27, 5) {real, imag} */,
  {32'hbf50a5b8, 32'hbec43920} /* (13, 27, 4) {real, imag} */,
  {32'hbf055b19, 32'h3f257a38} /* (13, 27, 3) {real, imag} */,
  {32'hbdd0b5d0, 32'hbe093b30} /* (13, 27, 2) {real, imag} */,
  {32'h3e57bd5a, 32'hbe08d7e8} /* (13, 27, 1) {real, imag} */,
  {32'h3ecf8ff1, 32'hbec9197e} /* (13, 27, 0) {real, imag} */,
  {32'h3eacdad8, 32'hbf314cd3} /* (13, 26, 31) {real, imag} */,
  {32'h3f40753a, 32'hbed4cbe8} /* (13, 26, 30) {real, imag} */,
  {32'h3f092ccc, 32'h3f945296} /* (13, 26, 29) {real, imag} */,
  {32'h3e007910, 32'h3fb34287} /* (13, 26, 28) {real, imag} */,
  {32'h3fb03d5a, 32'h3f2a60e4} /* (13, 26, 27) {real, imag} */,
  {32'h3f8f7260, 32'hbecee6b0} /* (13, 26, 26) {real, imag} */,
  {32'h3f333378, 32'hbe7d2560} /* (13, 26, 25) {real, imag} */,
  {32'h3e00d8f8, 32'h3f391d88} /* (13, 26, 24) {real, imag} */,
  {32'hbf99db85, 32'h3d2e2c80} /* (13, 26, 23) {real, imag} */,
  {32'hbf8effe8, 32'hbd2e4e20} /* (13, 26, 22) {real, imag} */,
  {32'hbe16650c, 32'hbd0ad3a0} /* (13, 26, 21) {real, imag} */,
  {32'h3ef79f39, 32'hbeb14d90} /* (13, 26, 20) {real, imag} */,
  {32'h3f014ccc, 32'hbf1cb4c0} /* (13, 26, 19) {real, imag} */,
  {32'h3f859a3b, 32'hbe9bf080} /* (13, 26, 18) {real, imag} */,
  {32'hbdd53f00, 32'h3f810bd0} /* (13, 26, 17) {real, imag} */,
  {32'hbe0c2528, 32'hbc9c2080} /* (13, 26, 16) {real, imag} */,
  {32'h3ecd0a6a, 32'hbee26b20} /* (13, 26, 15) {real, imag} */,
  {32'h3f5f8b36, 32'h3d83efc0} /* (13, 26, 14) {real, imag} */,
  {32'h3ef9170c, 32'h3f985996} /* (13, 26, 13) {real, imag} */,
  {32'h3e258150, 32'h3f574ac6} /* (13, 26, 12) {real, imag} */,
  {32'h3f1064f8, 32'hbeb9a6e8} /* (13, 26, 11) {real, imag} */,
  {32'h3eb2a971, 32'hbf4fadc8} /* (13, 26, 10) {real, imag} */,
  {32'h3f3d852a, 32'hbf406948} /* (13, 26, 9) {real, imag} */,
  {32'hbdf5a850, 32'hbf213450} /* (13, 26, 8) {real, imag} */,
  {32'hbee66e44, 32'hbf12107d} /* (13, 26, 7) {real, imag} */,
  {32'hbf46779a, 32'h3d22f800} /* (13, 26, 6) {real, imag} */,
  {32'hbf967844, 32'hbe133288} /* (13, 26, 5) {real, imag} */,
  {32'hbeb2a700, 32'hbed02cc8} /* (13, 26, 4) {real, imag} */,
  {32'h3eb9081a, 32'h3e8588f0} /* (13, 26, 3) {real, imag} */,
  {32'h3f99a3fd, 32'h3e571760} /* (13, 26, 2) {real, imag} */,
  {32'h3f70ef82, 32'h3e042e70} /* (13, 26, 1) {real, imag} */,
  {32'h3e8c3748, 32'hbd399620} /* (13, 26, 0) {real, imag} */,
  {32'h3ee60144, 32'hbe7f75e0} /* (13, 25, 31) {real, imag} */,
  {32'hbe707698, 32'hbf0df18c} /* (13, 25, 30) {real, imag} */,
  {32'hbed3add6, 32'h3e3a53b0} /* (13, 25, 29) {real, imag} */,
  {32'h3b7a1380, 32'h3f9bb0be} /* (13, 25, 28) {real, imag} */,
  {32'h3fb117ae, 32'h3f41f49c} /* (13, 25, 27) {real, imag} */,
  {32'h3fca7fc7, 32'hbe494f20} /* (13, 25, 26) {real, imag} */,
  {32'h3f698c0e, 32'hbf278998} /* (13, 25, 25) {real, imag} */,
  {32'h3ef0a3d4, 32'h3eb54310} /* (13, 25, 24) {real, imag} */,
  {32'h3b45b800, 32'hbe1d2500} /* (13, 25, 23) {real, imag} */,
  {32'hbed4ce08, 32'hbefeaa20} /* (13, 25, 22) {real, imag} */,
  {32'h3f151d37, 32'hbf0e838e} /* (13, 25, 21) {real, imag} */,
  {32'h3eacca28, 32'hbf536280} /* (13, 25, 20) {real, imag} */,
  {32'hbe78460c, 32'hbf120db4} /* (13, 25, 19) {real, imag} */,
  {32'h3f98b0f8, 32'hbed901b0} /* (13, 25, 18) {real, imag} */,
  {32'h3fbf07d9, 32'h3eb9b600} /* (13, 25, 17) {real, imag} */,
  {32'h3f37dc95, 32'hbec76c14} /* (13, 25, 16) {real, imag} */,
  {32'h3d06c920, 32'hbf41be20} /* (13, 25, 15) {real, imag} */,
  {32'hbee18af0, 32'hbef5fe80} /* (13, 25, 14) {real, imag} */,
  {32'hbe6323d8, 32'h3f124290} /* (13, 25, 13) {real, imag} */,
  {32'h3f07e1f3, 32'hbf5f55ce} /* (13, 25, 12) {real, imag} */,
  {32'h3e007706, 32'hbf653748} /* (13, 25, 11) {real, imag} */,
  {32'hbee83392, 32'hbe30a848} /* (13, 25, 10) {real, imag} */,
  {32'hbeda5d08, 32'h3f0b8f4c} /* (13, 25, 9) {real, imag} */,
  {32'hbee9a754, 32'hbe839178} /* (13, 25, 8) {real, imag} */,
  {32'hbeeec1fa, 32'hbcc2f080} /* (13, 25, 7) {real, imag} */,
  {32'hbf522bdc, 32'h3ef9ab88} /* (13, 25, 6) {real, imag} */,
  {32'hbfa1188e, 32'hbf9ef8a0} /* (13, 25, 5) {real, imag} */,
  {32'hbb0ecc00, 32'hbf699b3c} /* (13, 25, 4) {real, imag} */,
  {32'hbe28a0f6, 32'h3da437c0} /* (13, 25, 3) {real, imag} */,
  {32'h3f083f9a, 32'h3e1963d0} /* (13, 25, 2) {real, imag} */,
  {32'h3f1d4883, 32'hbee9e3fe} /* (13, 25, 1) {real, imag} */,
  {32'hbdac1274, 32'hbf459eb2} /* (13, 25, 0) {real, imag} */,
  {32'h3e7fced4, 32'h3d8b5940} /* (13, 24, 31) {real, imag} */,
  {32'hbf39cf8b, 32'hbec21380} /* (13, 24, 30) {real, imag} */,
  {32'hbe702f24, 32'hbf34df48} /* (13, 24, 29) {real, imag} */,
  {32'h3e104a70, 32'h3da7ba40} /* (13, 24, 28) {real, imag} */,
  {32'hbd17ef60, 32'h3e58ce80} /* (13, 24, 27) {real, imag} */,
  {32'h3f469994, 32'hbecb08b8} /* (13, 24, 26) {real, imag} */,
  {32'h3e82c368, 32'h3e842b20} /* (13, 24, 25) {real, imag} */,
  {32'h3f0c99b8, 32'h3ee19048} /* (13, 24, 24) {real, imag} */,
  {32'h3f859505, 32'hbe59c2a8} /* (13, 24, 23) {real, imag} */,
  {32'h3e978940, 32'hbe922718} /* (13, 24, 22) {real, imag} */,
  {32'h3f33508c, 32'hbf7c8aaa} /* (13, 24, 21) {real, imag} */,
  {32'hbf106dc6, 32'hbf31d6c0} /* (13, 24, 20) {real, imag} */,
  {32'hbf4cab4d, 32'h3ef0a9e0} /* (13, 24, 19) {real, imag} */,
  {32'hbe2b3a68, 32'h3f20dcec} /* (13, 24, 18) {real, imag} */,
  {32'h3f90c519, 32'h3e89d1a0} /* (13, 24, 17) {real, imag} */,
  {32'h3e8144f8, 32'h3e709380} /* (13, 24, 16) {real, imag} */,
  {32'hbf49d194, 32'h3e8beeb8} /* (13, 24, 15) {real, imag} */,
  {32'hbf9a74f8, 32'hbeb881b0} /* (13, 24, 14) {real, imag} */,
  {32'hbdffe110, 32'hbdd64ad0} /* (13, 24, 13) {real, imag} */,
  {32'h3d899b20, 32'hbfb021fc} /* (13, 24, 12) {real, imag} */,
  {32'hbfaae1a2, 32'hbf759cdc} /* (13, 24, 11) {real, imag} */,
  {32'hbf97c3e0, 32'hbefee750} /* (13, 24, 10) {real, imag} */,
  {32'hbf043a29, 32'h3f2f0250} /* (13, 24, 9) {real, imag} */,
  {32'hbf2ed3f6, 32'h3ea883e0} /* (13, 24, 8) {real, imag} */,
  {32'hbe650ca4, 32'h3e17bc80} /* (13, 24, 7) {real, imag} */,
  {32'hbe1f2ba0, 32'h3f5f2ffc} /* (13, 24, 6) {real, imag} */,
  {32'hbea6fac6, 32'hbf390e10} /* (13, 24, 5) {real, imag} */,
  {32'hbdddb3c8, 32'hbedfef50} /* (13, 24, 4) {real, imag} */,
  {32'hbf34e182, 32'h3e535540} /* (13, 24, 3) {real, imag} */,
  {32'h3ea090d2, 32'hbe76b4e0} /* (13, 24, 2) {real, imag} */,
  {32'h3f613710, 32'hbf8f2e98} /* (13, 24, 1) {real, imag} */,
  {32'h3efc374e, 32'hbf60653c} /* (13, 24, 0) {real, imag} */,
  {32'h3eb438ba, 32'hbf041234} /* (13, 23, 31) {real, imag} */,
  {32'h3e1b7230, 32'hbfbe08f2} /* (13, 23, 30) {real, imag} */,
  {32'h3d878ae8, 32'hbf8fa2ba} /* (13, 23, 29) {real, imag} */,
  {32'h3ca9a6e0, 32'h3dd31180} /* (13, 23, 28) {real, imag} */,
  {32'hbe3a5a10, 32'h3f31eb88} /* (13, 23, 27) {real, imag} */,
  {32'h3e0123c4, 32'h3eba6a40} /* (13, 23, 26) {real, imag} */,
  {32'h3f2e13c3, 32'h3f0d3cb8} /* (13, 23, 25) {real, imag} */,
  {32'h3f9e8d24, 32'hbd81f940} /* (13, 23, 24) {real, imag} */,
  {32'h3ed36d7c, 32'hbe22cbd0} /* (13, 23, 23) {real, imag} */,
  {32'hbe653c40, 32'hbf11ead8} /* (13, 23, 22) {real, imag} */,
  {32'h3e51be60, 32'hbfb10cb2} /* (13, 23, 21) {real, imag} */,
  {32'hbf4250fa, 32'hbe604b30} /* (13, 23, 20) {real, imag} */,
  {32'hbda025d0, 32'h3f29b3e4} /* (13, 23, 19) {real, imag} */,
  {32'hbf113e9f, 32'h3eca9a28} /* (13, 23, 18) {real, imag} */,
  {32'hbea72862, 32'hbe8166a8} /* (13, 23, 17) {real, imag} */,
  {32'hbee85d30, 32'hbdeab390} /* (13, 23, 16) {real, imag} */,
  {32'hbf39452f, 32'h3ec65ef0} /* (13, 23, 15) {real, imag} */,
  {32'hbf068885, 32'hbd85afc0} /* (13, 23, 14) {real, imag} */,
  {32'hbebac07a, 32'hbf044d42} /* (13, 23, 13) {real, imag} */,
  {32'hbf0eb86c, 32'hbf55cd91} /* (13, 23, 12) {real, imag} */,
  {32'hbf91b74b, 32'hbcf2ee80} /* (13, 23, 11) {real, imag} */,
  {32'hbe716cce, 32'h3d75f0c0} /* (13, 23, 10) {real, imag} */,
  {32'hbdb7e468, 32'hbf0ee810} /* (13, 23, 9) {real, imag} */,
  {32'hbdfe5918, 32'hbe6acc60} /* (13, 23, 8) {real, imag} */,
  {32'h3e5b3dd0, 32'hbf60c388} /* (13, 23, 7) {real, imag} */,
  {32'h3e6593de, 32'h3e084d40} /* (13, 23, 6) {real, imag} */,
  {32'h3f56ce23, 32'hbec14780} /* (13, 23, 5) {real, imag} */,
  {32'h3e805af4, 32'hbc6b5b00} /* (13, 23, 4) {real, imag} */,
  {32'hbf75d882, 32'h3eee85b8} /* (13, 23, 3) {real, imag} */,
  {32'hbf858e72, 32'hbe68f840} /* (13, 23, 2) {real, imag} */,
  {32'hbebfe0c6, 32'hbf8475cc} /* (13, 23, 1) {real, imag} */,
  {32'h3e38a7a4, 32'hbf25227c} /* (13, 23, 0) {real, imag} */,
  {32'h3e94bd58, 32'hbe955384} /* (13, 22, 31) {real, imag} */,
  {32'hbd5a6cb0, 32'hbfb84f09} /* (13, 22, 30) {real, imag} */,
  {32'hbf0cf06e, 32'hbf95958c} /* (13, 22, 29) {real, imag} */,
  {32'hbebfa31c, 32'h3f1b5908} /* (13, 22, 28) {real, imag} */,
  {32'h3dc7d080, 32'h3f39b594} /* (13, 22, 27) {real, imag} */,
  {32'h3e81d93a, 32'h3f0949d4} /* (13, 22, 26) {real, imag} */,
  {32'h3e500774, 32'h3f2d7e78} /* (13, 22, 25) {real, imag} */,
  {32'h3db7b8c0, 32'h3d7decc0} /* (13, 22, 24) {real, imag} */,
  {32'hbf1e9558, 32'h3e6b6e20} /* (13, 22, 23) {real, imag} */,
  {32'hbf1cd056, 32'hbe618d10} /* (13, 22, 22) {real, imag} */,
  {32'hbee4bb99, 32'hbf9df7d3} /* (13, 22, 21) {real, imag} */,
  {32'hbf03f5ea, 32'hbf1c808a} /* (13, 22, 20) {real, imag} */,
  {32'h3ede2907, 32'h3f38b8a4} /* (13, 22, 19) {real, imag} */,
  {32'hbd026940, 32'hbcb05b80} /* (13, 22, 18) {real, imag} */,
  {32'hbf6514b1, 32'hbecdbc98} /* (13, 22, 17) {real, imag} */,
  {32'hbfa711b4, 32'hbdcc5c40} /* (13, 22, 16) {real, imag} */,
  {32'hbf551866, 32'h3ee82314} /* (13, 22, 15) {real, imag} */,
  {32'hbf6f6f44, 32'h3ef74760} /* (13, 22, 14) {real, imag} */,
  {32'hbf6b7958, 32'hbe6929c0} /* (13, 22, 13) {real, imag} */,
  {32'hbee91070, 32'hbf6648e6} /* (13, 22, 12) {real, imag} */,
  {32'h3ea534e7, 32'h3cf18e60} /* (13, 22, 11) {real, imag} */,
  {32'hbe23bf08, 32'hbd4ac920} /* (13, 22, 10) {real, imag} */,
  {32'hbf65fdc4, 32'hbd760b40} /* (13, 22, 9) {real, imag} */,
  {32'hbf04ca55, 32'h3f43d218} /* (13, 22, 8) {real, imag} */,
  {32'hbde91ff0, 32'h3daf1980} /* (13, 22, 7) {real, imag} */,
  {32'hbeb20e38, 32'h3df790e0} /* (13, 22, 6) {real, imag} */,
  {32'h3f087ff7, 32'h3f63ac9c} /* (13, 22, 5) {real, imag} */,
  {32'h3ef3c0dc, 32'h3ef47ab8} /* (13, 22, 4) {real, imag} */,
  {32'h3ed5f2b8, 32'h3f254770} /* (13, 22, 3) {real, imag} */,
  {32'hbee21490, 32'h3f8ed530} /* (13, 22, 2) {real, imag} */,
  {32'hbece4a45, 32'h3c9b5ec0} /* (13, 22, 1) {real, imag} */,
  {32'h3b1675c0, 32'hbf05daf6} /* (13, 22, 0) {real, imag} */,
  {32'h3e7f7edc, 32'h3f473bf0} /* (13, 21, 31) {real, imag} */,
  {32'hbe411bc6, 32'h3f19e1ec} /* (13, 21, 30) {real, imag} */,
  {32'hbf7bce70, 32'hbf5bb43d} /* (13, 21, 29) {real, imag} */,
  {32'hbf9a10e4, 32'h3e9a65ec} /* (13, 21, 28) {real, imag} */,
  {32'hbd9a55f0, 32'h3f3dde84} /* (13, 21, 27) {real, imag} */,
  {32'h3f0fb85e, 32'h3c8be6e0} /* (13, 21, 26) {real, imag} */,
  {32'hbf245982, 32'h3ef367b4} /* (13, 21, 25) {real, imag} */,
  {32'hbf60db53, 32'h3cd6bcc0} /* (13, 21, 24) {real, imag} */,
  {32'hbea40ca8, 32'h3e5049f8} /* (13, 21, 23) {real, imag} */,
  {32'h3e7bbea4, 32'h3f505393} /* (13, 21, 22) {real, imag} */,
  {32'hbc85af78, 32'hbe10dba0} /* (13, 21, 21) {real, imag} */,
  {32'h3d19b220, 32'hbf2b1654} /* (13, 21, 20) {real, imag} */,
  {32'h3eb4c600, 32'h3eabf1f4} /* (13, 21, 19) {real, imag} */,
  {32'h3e1d53a4, 32'hbd9a9dc0} /* (13, 21, 18) {real, imag} */,
  {32'h3f059460, 32'hbdced5d0} /* (13, 21, 17) {real, imag} */,
  {32'hbe9e45c2, 32'h3f65d268} /* (13, 21, 16) {real, imag} */,
  {32'hbf0dea14, 32'hbda8afd0} /* (13, 21, 15) {real, imag} */,
  {32'hbf1cf42c, 32'hbe51e330} /* (13, 21, 14) {real, imag} */,
  {32'hbefb176c, 32'h3d4ebbc0} /* (13, 21, 13) {real, imag} */,
  {32'hbdeb9810, 32'h3c885320} /* (13, 21, 12) {real, imag} */,
  {32'h3f8d6d41, 32'h3ebb7df7} /* (13, 21, 11) {real, imag} */,
  {32'h3e793d80, 32'h3f582481} /* (13, 21, 10) {real, imag} */,
  {32'hbe21b5de, 32'h3fc4b99c} /* (13, 21, 9) {real, imag} */,
  {32'h3d1c7310, 32'h3fcec69e} /* (13, 21, 8) {real, imag} */,
  {32'hbd96a4c0, 32'h3f3e81b7} /* (13, 21, 7) {real, imag} */,
  {32'hbea11b10, 32'h3e37d334} /* (13, 21, 6) {real, imag} */,
  {32'h3e07f0da, 32'h3f4f3940} /* (13, 21, 5) {real, imag} */,
  {32'hbeff576c, 32'h3f05c22c} /* (13, 21, 4) {real, imag} */,
  {32'h3e746ae6, 32'h3e10e990} /* (13, 21, 3) {real, imag} */,
  {32'hbeb06acd, 32'h3fc3f369} /* (13, 21, 2) {real, imag} */,
  {32'hbf17293c, 32'h3f20661a} /* (13, 21, 1) {real, imag} */,
  {32'h3d8e2410, 32'hbc1fd368} /* (13, 21, 0) {real, imag} */,
  {32'h3e20b250, 32'h3d52e680} /* (13, 20, 31) {real, imag} */,
  {32'h3e9030ce, 32'h3efdfd28} /* (13, 20, 30) {real, imag} */,
  {32'hbebd022c, 32'hbf66e4e4} /* (13, 20, 29) {real, imag} */,
  {32'hbf5fdb86, 32'h3e434da0} /* (13, 20, 28) {real, imag} */,
  {32'h3ed94e68, 32'h3fa0fdec} /* (13, 20, 27) {real, imag} */,
  {32'h3e167cc0, 32'h3eddbcd0} /* (13, 20, 26) {real, imag} */,
  {32'hbe62e660, 32'h3d562e80} /* (13, 20, 25) {real, imag} */,
  {32'hbf4207c8, 32'h3f066da8} /* (13, 20, 24) {real, imag} */,
  {32'hbfb3e023, 32'hbe722080} /* (13, 20, 23) {real, imag} */,
  {32'hbef8df4f, 32'hbeb7b140} /* (13, 20, 22) {real, imag} */,
  {32'h3f27156c, 32'h3d8a5490} /* (13, 20, 21) {real, imag} */,
  {32'h3e9d84d4, 32'hbe52e128} /* (13, 20, 20) {real, imag} */,
  {32'h3ee8dcd0, 32'hbe676f30} /* (13, 20, 19) {real, imag} */,
  {32'h3ee83c30, 32'h3ca3c480} /* (13, 20, 18) {real, imag} */,
  {32'h3fc031ce, 32'hbf010260} /* (13, 20, 17) {real, imag} */,
  {32'h3f23662b, 32'h3f1a0bd4} /* (13, 20, 16) {real, imag} */,
  {32'hbeb59340, 32'hbe516660} /* (13, 20, 15) {real, imag} */,
  {32'hbf34acdd, 32'hbf3e1e68} /* (13, 20, 14) {real, imag} */,
  {32'hbe82309d, 32'hbf8b53aa} /* (13, 20, 13) {real, imag} */,
  {32'h3ee46b34, 32'hbf0aa4f4} /* (13, 20, 12) {real, imag} */,
  {32'h3f785a2f, 32'h3ea2eb20} /* (13, 20, 11) {real, imag} */,
  {32'h3fa3b374, 32'h3ea4a362} /* (13, 20, 10) {real, imag} */,
  {32'h3dc26de4, 32'h3efdc2c0} /* (13, 20, 9) {real, imag} */,
  {32'hbebb2692, 32'h3ee443b0} /* (13, 20, 8) {real, imag} */,
  {32'h3f1f0e04, 32'hbf0a0254} /* (13, 20, 7) {real, imag} */,
  {32'h3f99833f, 32'h3d429d00} /* (13, 20, 6) {real, imag} */,
  {32'h3f88a3cb, 32'h3f93a897} /* (13, 20, 5) {real, imag} */,
  {32'hbedc189c, 32'h3f58c5a8} /* (13, 20, 4) {real, imag} */,
  {32'hbfb7c143, 32'hbf149a00} /* (13, 20, 3) {real, imag} */,
  {32'hbf6d27f2, 32'h3eee674c} /* (13, 20, 2) {real, imag} */,
  {32'hbd9f9148, 32'h3e516430} /* (13, 20, 1) {real, imag} */,
  {32'hbd367200, 32'h3d882220} /* (13, 20, 0) {real, imag} */,
  {32'hbea1b07d, 32'hbf599d60} /* (13, 19, 31) {real, imag} */,
  {32'hbcff21a0, 32'hbe3df900} /* (13, 19, 30) {real, imag} */,
  {32'h3eb26814, 32'hbd97f070} /* (13, 19, 29) {real, imag} */,
  {32'h3d12c720, 32'h3f5ec8aa} /* (13, 19, 28) {real, imag} */,
  {32'h3f73f254, 32'h3f60adbc} /* (13, 19, 27) {real, imag} */,
  {32'h3f251b12, 32'h3f007a3c} /* (13, 19, 26) {real, imag} */,
  {32'h3f30434c, 32'h3f24aa8c} /* (13, 19, 25) {real, imag} */,
  {32'h3ee7559c, 32'h3f4f1198} /* (13, 19, 24) {real, imag} */,
  {32'hbf2fb280, 32'hbf5cca94} /* (13, 19, 23) {real, imag} */,
  {32'hbf6dd55b, 32'hbfa0a908} /* (13, 19, 22) {real, imag} */,
  {32'hbd44b980, 32'h3f026b0d} /* (13, 19, 21) {real, imag} */,
  {32'h3ddfbb30, 32'hbbdac800} /* (13, 19, 20) {real, imag} */,
  {32'hbd84ab70, 32'hbfc266ff} /* (13, 19, 19) {real, imag} */,
  {32'hbc7b0980, 32'hbf573004} /* (13, 19, 18) {real, imag} */,
  {32'h3f6f019c, 32'hbe9cee20} /* (13, 19, 17) {real, imag} */,
  {32'hbe1f5cf0, 32'h3e920e40} /* (13, 19, 16) {real, imag} */,
  {32'hbf1a081b, 32'hbe4ba888} /* (13, 19, 15) {real, imag} */,
  {32'hbe07e568, 32'h3edea670} /* (13, 19, 14) {real, imag} */,
  {32'h3f10d7ec, 32'h3e25acc0} /* (13, 19, 13) {real, imag} */,
  {32'h3ecd77a6, 32'h3e2a7310} /* (13, 19, 12) {real, imag} */,
  {32'h3eb8a862, 32'h3f81f915} /* (13, 19, 11) {real, imag} */,
  {32'h3f6b76da, 32'h3eba0170} /* (13, 19, 10) {real, imag} */,
  {32'h3e28cd38, 32'hbe19d9e0} /* (13, 19, 9) {real, imag} */,
  {32'hbf040f41, 32'hbf233c10} /* (13, 19, 8) {real, imag} */,
  {32'hbcd401c0, 32'hbf5830a8} /* (13, 19, 7) {real, imag} */,
  {32'h3da85d40, 32'h3e10d980} /* (13, 19, 6) {real, imag} */,
  {32'h3d93c3c8, 32'h3e0578a0} /* (13, 19, 5) {real, imag} */,
  {32'hbd1cb440, 32'h3dacc7c0} /* (13, 19, 4) {real, imag} */,
  {32'hbf4510b8, 32'h3ecaa828} /* (13, 19, 3) {real, imag} */,
  {32'hbf93375a, 32'h3f188a08} /* (13, 19, 2) {real, imag} */,
  {32'hbea19a32, 32'hbecae0d0} /* (13, 19, 1) {real, imag} */,
  {32'hbe2282a2, 32'hbe078670} /* (13, 19, 0) {real, imag} */,
  {32'hbf21601a, 32'hbe91e040} /* (13, 18, 31) {real, imag} */,
  {32'hbf2c81e0, 32'h3ebef210} /* (13, 18, 30) {real, imag} */,
  {32'h3e52c318, 32'h3e19f900} /* (13, 18, 29) {real, imag} */,
  {32'hbe1289de, 32'hbd854b40} /* (13, 18, 28) {real, imag} */,
  {32'hbeb05ab8, 32'hbed25638} /* (13, 18, 27) {real, imag} */,
  {32'h3e76aab4, 32'hbe8fecb0} /* (13, 18, 26) {real, imag} */,
  {32'h3f01351e, 32'h3f296a0a} /* (13, 18, 25) {real, imag} */,
  {32'h3ed64b60, 32'hbf0f1114} /* (13, 18, 24) {real, imag} */,
  {32'h3d6c55c0, 32'hbfa7726a} /* (13, 18, 23) {real, imag} */,
  {32'hbf17bd5c, 32'hbec88240} /* (13, 18, 22) {real, imag} */,
  {32'hbe52ae48, 32'h3e092130} /* (13, 18, 21) {real, imag} */,
  {32'hbf37af21, 32'hbe25b6c0} /* (13, 18, 20) {real, imag} */,
  {32'hbf902feb, 32'hbfa6d32a} /* (13, 18, 19) {real, imag} */,
  {32'h3da71240, 32'hbeb04dc0} /* (13, 18, 18) {real, imag} */,
  {32'h3f020486, 32'h3ed640a8} /* (13, 18, 17) {real, imag} */,
  {32'hbf18bb30, 32'h3f34dc84} /* (13, 18, 16) {real, imag} */,
  {32'hbf15a9cc, 32'h3f3cb270} /* (13, 18, 15) {real, imag} */,
  {32'hbdb4b2a0, 32'h3faf141c} /* (13, 18, 14) {real, imag} */,
  {32'h3f2e96f6, 32'h3fb5ea80} /* (13, 18, 13) {real, imag} */,
  {32'h3ebbf424, 32'h3f1bc4b8} /* (13, 18, 12) {real, imag} */,
  {32'hbcdcd8c0, 32'h3f091eb4} /* (13, 18, 11) {real, imag} */,
  {32'hbf6fd7a0, 32'h3fa56f69} /* (13, 18, 10) {real, imag} */,
  {32'hbf48dc9c, 32'h3e781170} /* (13, 18, 9) {real, imag} */,
  {32'hbe9327ee, 32'hbcb4bc00} /* (13, 18, 8) {real, imag} */,
  {32'hbf361a6c, 32'h3f2b5abc} /* (13, 18, 7) {real, imag} */,
  {32'hbf8d674a, 32'h3e986330} /* (13, 18, 6) {real, imag} */,
  {32'hbf31fc3c, 32'hbe2b7c30} /* (13, 18, 5) {real, imag} */,
  {32'hbd685cc0, 32'h3dd7ed80} /* (13, 18, 4) {real, imag} */,
  {32'hbe5e36f0, 32'h3e4b3010} /* (13, 18, 3) {real, imag} */,
  {32'h3c145be0, 32'h3efcc980} /* (13, 18, 2) {real, imag} */,
  {32'h3ee30eac, 32'hbeedf158} /* (13, 18, 1) {real, imag} */,
  {32'hbe2dd8c8, 32'hbe96423c} /* (13, 18, 0) {real, imag} */,
  {32'hbf03c664, 32'hbeabe990} /* (13, 17, 31) {real, imag} */,
  {32'hbf560eb6, 32'h3e2120a0} /* (13, 17, 30) {real, imag} */,
  {32'hbf12b85c, 32'h3f1316d4} /* (13, 17, 29) {real, imag} */,
  {32'hbf7d7cb9, 32'hbfa0a584} /* (13, 17, 28) {real, imag} */,
  {32'hbfa04029, 32'hbf55785c} /* (13, 17, 27) {real, imag} */,
  {32'h3e26e2e0, 32'hbf1287b0} /* (13, 17, 26) {real, imag} */,
  {32'h3f14c46a, 32'hbf2a9884} /* (13, 17, 25) {real, imag} */,
  {32'h3ebff0e0, 32'hbf3e2e70} /* (13, 17, 24) {real, imag} */,
  {32'h3f0cfba1, 32'hbe887108} /* (13, 17, 23) {real, imag} */,
  {32'hbf2abf76, 32'h3ec3fad0} /* (13, 17, 22) {real, imag} */,
  {32'hbf775228, 32'hbdde2c20} /* (13, 17, 21) {real, imag} */,
  {32'hbdb83518, 32'h3ea75f00} /* (13, 17, 20) {real, imag} */,
  {32'hbe768720, 32'hbe982b14} /* (13, 17, 19) {real, imag} */,
  {32'hbd8f4be0, 32'hbd42a2c0} /* (13, 17, 18) {real, imag} */,
  {32'h3f11b9a0, 32'h3e3915b0} /* (13, 17, 17) {real, imag} */,
  {32'hbe020210, 32'h3ec60d10} /* (13, 17, 16) {real, imag} */,
  {32'hbd3cb5a0, 32'h3f8ed58e} /* (13, 17, 15) {real, imag} */,
  {32'h3e8fb214, 32'h3fb202ac} /* (13, 17, 14) {real, imag} */,
  {32'h3ed41e58, 32'h3f4ba504} /* (13, 17, 13) {real, imag} */,
  {32'h3e92dec8, 32'h3e1eade0} /* (13, 17, 12) {real, imag} */,
  {32'h3f42ab7c, 32'hbd5217c0} /* (13, 17, 11) {real, imag} */,
  {32'hbf19b296, 32'h3f3e14ed} /* (13, 17, 10) {real, imag} */,
  {32'hbedc9860, 32'h3d6dbf00} /* (13, 17, 9) {real, imag} */,
  {32'h3ea360bc, 32'hbe366a60} /* (13, 17, 8) {real, imag} */,
  {32'h3e220736, 32'h3f484b2c} /* (13, 17, 7) {real, imag} */,
  {32'hbf66f76e, 32'h3f46132c} /* (13, 17, 6) {real, imag} */,
  {32'hbec32508, 32'h3e93f9c0} /* (13, 17, 5) {real, imag} */,
  {32'h3e8b4aa8, 32'h3f1cce3c} /* (13, 17, 4) {real, imag} */,
  {32'h3ece6f46, 32'h3e852ab0} /* (13, 17, 3) {real, imag} */,
  {32'h3ea67f31, 32'hbdb2be80} /* (13, 17, 2) {real, imag} */,
  {32'h3f093b40, 32'h3c62d000} /* (13, 17, 1) {real, imag} */,
  {32'h3d094460, 32'h3d850a70} /* (13, 17, 0) {real, imag} */,
  {32'h3f144b7a, 32'hbc735400} /* (13, 16, 31) {real, imag} */,
  {32'h3dac8eb0, 32'hbe6f5c80} /* (13, 16, 30) {real, imag} */,
  {32'hbf3e9aab, 32'hbea7e5f0} /* (13, 16, 29) {real, imag} */,
  {32'hbf1e59c0, 32'hbf5d6886} /* (13, 16, 28) {real, imag} */,
  {32'hbf8591f1, 32'hbf56a0ce} /* (13, 16, 27) {real, imag} */,
  {32'hbf49aaee, 32'hbe074148} /* (13, 16, 26) {real, imag} */,
  {32'hbe945658, 32'hbefbfc28} /* (13, 16, 25) {real, imag} */,
  {32'hbebe37a9, 32'hbcf3b080} /* (13, 16, 24) {real, imag} */,
  {32'h3e84d292, 32'hbec37638} /* (13, 16, 23) {real, imag} */,
  {32'hbed5b7d0, 32'hbefcf3a8} /* (13, 16, 22) {real, imag} */,
  {32'hbce06ae0, 32'hbea959ae} /* (13, 16, 21) {real, imag} */,
  {32'h3fc388b4, 32'hbf0ff998} /* (13, 16, 20) {real, imag} */,
  {32'h3fd07504, 32'hbf8fd684} /* (13, 16, 19) {real, imag} */,
  {32'h3f882086, 32'hbe9dd34c} /* (13, 16, 18) {real, imag} */,
  {32'h3e04152c, 32'h3eb1b898} /* (13, 16, 17) {real, imag} */,
  {32'hbfa9a6fb, 32'h3f853878} /* (13, 16, 16) {real, imag} */,
  {32'hbf400869, 32'h3effa500} /* (13, 16, 15) {real, imag} */,
  {32'h3f64e8f5, 32'h3f509250} /* (13, 16, 14) {real, imag} */,
  {32'hbe05ec7c, 32'h3b037400} /* (13, 16, 13) {real, imag} */,
  {32'hbfa06a94, 32'hbe9f216c} /* (13, 16, 12) {real, imag} */,
  {32'hbec3dd16, 32'hbf3858e3} /* (13, 16, 11) {real, imag} */,
  {32'hbef43d90, 32'hbda099a0} /* (13, 16, 10) {real, imag} */,
  {32'h3f1ea4d6, 32'h3e0ff880} /* (13, 16, 9) {real, imag} */,
  {32'h3faebd1c, 32'hbe044ed0} /* (13, 16, 8) {real, imag} */,
  {32'h3f5a7e70, 32'h3dc80d00} /* (13, 16, 7) {real, imag} */,
  {32'h3e01d550, 32'hbe1f50f0} /* (13, 16, 6) {real, imag} */,
  {32'h3f090740, 32'h3d9aa460} /* (13, 16, 5) {real, imag} */,
  {32'h3f848ac8, 32'h3d6a4740} /* (13, 16, 4) {real, imag} */,
  {32'h3f9fa327, 32'hbdbad060} /* (13, 16, 3) {real, imag} */,
  {32'h3ef37bbc, 32'hbe7cf760} /* (13, 16, 2) {real, imag} */,
  {32'hb9a1f000, 32'hbee1c678} /* (13, 16, 1) {real, imag} */,
  {32'h3eb445f6, 32'hbf134ffc} /* (13, 16, 0) {real, imag} */,
  {32'h3f2052d1, 32'hbdcfd680} /* (13, 15, 31) {real, imag} */,
  {32'h3f926682, 32'hbceb0d00} /* (13, 15, 30) {real, imag} */,
  {32'h3ea56cf8, 32'hbe877060} /* (13, 15, 29) {real, imag} */,
  {32'hbfac5555, 32'h3d38a400} /* (13, 15, 28) {real, imag} */,
  {32'hbfa1f686, 32'hbfb4098b} /* (13, 15, 27) {real, imag} */,
  {32'hbfe38e9a, 32'hbf383f5a} /* (13, 15, 26) {real, imag} */,
  {32'hbfd43eb4, 32'h3e346a10} /* (13, 15, 25) {real, imag} */,
  {32'hbf3b39f5, 32'h3e5c2c78} /* (13, 15, 24) {real, imag} */,
  {32'h3f279f94, 32'hbf05454c} /* (13, 15, 23) {real, imag} */,
  {32'hbec311c8, 32'hbfd51d77} /* (13, 15, 22) {real, imag} */,
  {32'hbe09a2d2, 32'hbf80c87e} /* (13, 15, 21) {real, imag} */,
  {32'h3f8ecd86, 32'hbefdbe20} /* (13, 15, 20) {real, imag} */,
  {32'h3fa1d0a2, 32'hbf836fba} /* (13, 15, 19) {real, imag} */,
  {32'h3ff1c4e4, 32'hbf3e160f} /* (13, 15, 18) {real, imag} */,
  {32'h3f198ed4, 32'hbdceccf0} /* (13, 15, 17) {real, imag} */,
  {32'hbf81233a, 32'h3f7128a0} /* (13, 15, 16) {real, imag} */,
  {32'hbf5ea5b5, 32'h3f384b30} /* (13, 15, 15) {real, imag} */,
  {32'h3e9d1f34, 32'h3ed94c50} /* (13, 15, 14) {real, imag} */,
  {32'hbf155c83, 32'h3eb73a78} /* (13, 15, 13) {real, imag} */,
  {32'hc0114714, 32'h3ef899d0} /* (13, 15, 12) {real, imag} */,
  {32'hbfd47323, 32'hbf13a884} /* (13, 15, 11) {real, imag} */,
  {32'hbf26c340, 32'h3eb35348} /* (13, 15, 10) {real, imag} */,
  {32'h3e8ba0d2, 32'h3f5c1c9c} /* (13, 15, 9) {real, imag} */,
  {32'h3f002cf2, 32'h3f8a5ddc} /* (13, 15, 8) {real, imag} */,
  {32'h3e947038, 32'h3c571800} /* (13, 15, 7) {real, imag} */,
  {32'h3ecdd330, 32'hbf479c6c} /* (13, 15, 6) {real, imag} */,
  {32'h3ed11028, 32'hbf6832c6} /* (13, 15, 5) {real, imag} */,
  {32'h3f31d8a8, 32'hbef0d530} /* (13, 15, 4) {real, imag} */,
  {32'h3fe48e32, 32'hbeabc288} /* (13, 15, 3) {real, imag} */,
  {32'h3fcbd886, 32'hbe4efc70} /* (13, 15, 2) {real, imag} */,
  {32'hbf162136, 32'hbeb961e8} /* (13, 15, 1) {real, imag} */,
  {32'hbec9727d, 32'hbf56cac4} /* (13, 15, 0) {real, imag} */,
  {32'hbea206e3, 32'hbf2a30d2} /* (13, 14, 31) {real, imag} */,
  {32'h3ef4f000, 32'hbf524de8} /* (13, 14, 30) {real, imag} */,
  {32'h3e8fe020, 32'h3e0a1250} /* (13, 14, 29) {real, imag} */,
  {32'hbf6cf894, 32'h3f16f64a} /* (13, 14, 28) {real, imag} */,
  {32'hbf5af660, 32'hbf97071b} /* (13, 14, 27) {real, imag} */,
  {32'hbef3fc98, 32'h3cb21200} /* (13, 14, 26) {real, imag} */,
  {32'hbf705db4, 32'h3f64d808} /* (13, 14, 25) {real, imag} */,
  {32'hbf11347c, 32'h3e007eb0} /* (13, 14, 24) {real, imag} */,
  {32'h3f7097a0, 32'hbeb62998} /* (13, 14, 23) {real, imag} */,
  {32'h3f0a39b8, 32'hbfb816ec} /* (13, 14, 22) {real, imag} */,
  {32'h3c25b400, 32'hbfac28b2} /* (13, 14, 21) {real, imag} */,
  {32'hbee783cc, 32'hbe873dd4} /* (13, 14, 20) {real, imag} */,
  {32'h3e70f040, 32'hbf2eceda} /* (13, 14, 19) {real, imag} */,
  {32'h3f6a486a, 32'hbe3bccd8} /* (13, 14, 18) {real, imag} */,
  {32'h3e553a64, 32'h3e800268} /* (13, 14, 17) {real, imag} */,
  {32'hbf24f4cc, 32'h3e923198} /* (13, 14, 16) {real, imag} */,
  {32'hbe462090, 32'h3e194700} /* (13, 14, 15) {real, imag} */,
  {32'h3c9c2940, 32'h3eb26a1c} /* (13, 14, 14) {real, imag} */,
  {32'hbf3b1569, 32'h3f32d5ec} /* (13, 14, 13) {real, imag} */,
  {32'hbf847f95, 32'h3f8843ea} /* (13, 14, 12) {real, imag} */,
  {32'h3f0a9878, 32'h3da60260} /* (13, 14, 11) {real, imag} */,
  {32'h3f7850fa, 32'h3e689c30} /* (13, 14, 10) {real, imag} */,
  {32'h3eca2694, 32'hbd251f80} /* (13, 14, 9) {real, imag} */,
  {32'hbed6cae4, 32'h3d827300} /* (13, 14, 8) {real, imag} */,
  {32'hbf6fbffc, 32'hbe363aa0} /* (13, 14, 7) {real, imag} */,
  {32'hbed76c66, 32'hbea9bbc0} /* (13, 14, 6) {real, imag} */,
  {32'hbf49ca52, 32'hbf12d484} /* (13, 14, 5) {real, imag} */,
  {32'hbed789d8, 32'hbd3e0540} /* (13, 14, 4) {real, imag} */,
  {32'h3f4e7fd6, 32'hbc8f6080} /* (13, 14, 3) {real, imag} */,
  {32'h3f97a45e, 32'h3dbd6530} /* (13, 14, 2) {real, imag} */,
  {32'hbf6dd810, 32'hbe2c1558} /* (13, 14, 1) {real, imag} */,
  {32'hbf4b6a11, 32'hbe2fc010} /* (13, 14, 0) {real, imag} */,
  {32'h3d87afc4, 32'hbf3a8cb8} /* (13, 13, 31) {real, imag} */,
  {32'h3f348fbe, 32'hbf615e74} /* (13, 13, 30) {real, imag} */,
  {32'h3e96f880, 32'hbf06ae18} /* (13, 13, 29) {real, imag} */,
  {32'h3e645880, 32'hbed50670} /* (13, 13, 28) {real, imag} */,
  {32'hbf936816, 32'hbd208a80} /* (13, 13, 27) {real, imag} */,
  {32'hbe962464, 32'h3f4473a4} /* (13, 13, 26) {real, imag} */,
  {32'h3d8287f0, 32'h3ec0fc30} /* (13, 13, 25) {real, imag} */,
  {32'hbf1eea42, 32'hbdacc000} /* (13, 13, 24) {real, imag} */,
  {32'hbe981760, 32'hbebd6830} /* (13, 13, 23) {real, imag} */,
  {32'h3ed49f40, 32'hbf6ea7b8} /* (13, 13, 22) {real, imag} */,
  {32'h3ee3b618, 32'hbeb1e802} /* (13, 13, 21) {real, imag} */,
  {32'hbf3c9f70, 32'h3e040940} /* (13, 13, 20) {real, imag} */,
  {32'h3e13c41c, 32'h3cdb9100} /* (13, 13, 19) {real, imag} */,
  {32'hbd84de80, 32'h3eae6a40} /* (13, 13, 18) {real, imag} */,
  {32'hbec142d4, 32'h3f7db728} /* (13, 13, 17) {real, imag} */,
  {32'hbee18a48, 32'h3f5e8e6c} /* (13, 13, 16) {real, imag} */,
  {32'hbf09a105, 32'hbf92ba9e} /* (13, 13, 15) {real, imag} */,
  {32'h3e114ddc, 32'hbf27960b} /* (13, 13, 14) {real, imag} */,
  {32'hbeb544f8, 32'h3eb103e0} /* (13, 13, 13) {real, imag} */,
  {32'hbbde8800, 32'h3f7b4340} /* (13, 13, 12) {real, imag} */,
  {32'h3fbe0da6, 32'h3ea735f8} /* (13, 13, 11) {real, imag} */,
  {32'h3fce669f, 32'h3eb98200} /* (13, 13, 10) {real, imag} */,
  {32'h3f8ee8b6, 32'hbf20e5c8} /* (13, 13, 9) {real, imag} */,
  {32'h3edae4ec, 32'hbf31b0b8} /* (13, 13, 8) {real, imag} */,
  {32'hbe180e10, 32'hbecfa80c} /* (13, 13, 7) {real, imag} */,
  {32'h3db67390, 32'h3ea1fd00} /* (13, 13, 6) {real, imag} */,
  {32'hbf43ac4c, 32'h3e2e8aa0} /* (13, 13, 5) {real, imag} */,
  {32'hbf7ae65f, 32'hbe00f8c0} /* (13, 13, 4) {real, imag} */,
  {32'hbf0e6cb4, 32'hbf09ed88} /* (13, 13, 3) {real, imag} */,
  {32'h3e8aee38, 32'hbf528aca} /* (13, 13, 2) {real, imag} */,
  {32'hbea22fa3, 32'hbfaf18f0} /* (13, 13, 1) {real, imag} */,
  {32'hbf3a2a2e, 32'hbeb14a90} /* (13, 13, 0) {real, imag} */,
  {32'h3eac5533, 32'hbf88820e} /* (13, 12, 31) {real, imag} */,
  {32'h3f58ad5a, 32'hbf8c3104} /* (13, 12, 30) {real, imag} */,
  {32'h3e9e51ec, 32'hbeb2cc28} /* (13, 12, 29) {real, imag} */,
  {32'hbdbf30d8, 32'hbf225340} /* (13, 12, 28) {real, imag} */,
  {32'hbf73a8b4, 32'hbef88b40} /* (13, 12, 27) {real, imag} */,
  {32'hbf0432ae, 32'h3f3393b0} /* (13, 12, 26) {real, imag} */,
  {32'hbe43e0c0, 32'h3f6522c8} /* (13, 12, 25) {real, imag} */,
  {32'hbf38935e, 32'h3e9976d0} /* (13, 12, 24) {real, imag} */,
  {32'hbf4b5af5, 32'h3f21c468} /* (13, 12, 23) {real, imag} */,
  {32'hbf3ee2f9, 32'h3db7c480} /* (13, 12, 22) {real, imag} */,
  {32'h3dd2daf8, 32'hbe4ec43c} /* (13, 12, 21) {real, imag} */,
  {32'hbef554d9, 32'hbea5f1f0} /* (13, 12, 20) {real, imag} */,
  {32'hbebe9afa, 32'hbe9353d8} /* (13, 12, 19) {real, imag} */,
  {32'h3d74c020, 32'h3f14a8d8} /* (13, 12, 18) {real, imag} */,
  {32'h3efb1b88, 32'h3f207940} /* (13, 12, 17) {real, imag} */,
  {32'hbe81bea3, 32'h3e025f80} /* (13, 12, 16) {real, imag} */,
  {32'hbebd1740, 32'hbf8fa776} /* (13, 12, 15) {real, imag} */,
  {32'h3e11e5f7, 32'hbe238714} /* (13, 12, 14) {real, imag} */,
  {32'hbd431300, 32'h3ebaa658} /* (13, 12, 13) {real, imag} */,
  {32'hbee28d74, 32'h3dbfb740} /* (13, 12, 12) {real, imag} */,
  {32'h3f8e1ff6, 32'h3f0cbc6e} /* (13, 12, 11) {real, imag} */,
  {32'h3eada028, 32'h3ea8d8c4} /* (13, 12, 10) {real, imag} */,
  {32'hbea0009a, 32'hbf1819d8} /* (13, 12, 9) {real, imag} */,
  {32'h3f6b4e45, 32'hbe9023c8} /* (13, 12, 8) {real, imag} */,
  {32'h3edf26c0, 32'hbf88eee9} /* (13, 12, 7) {real, imag} */,
  {32'hbf059dcb, 32'hbf55e640} /* (13, 12, 6) {real, imag} */,
  {32'hbed45370, 32'h3e27b7c0} /* (13, 12, 5) {real, imag} */,
  {32'hbe20ccdc, 32'h3ed21fa0} /* (13, 12, 4) {real, imag} */,
  {32'h3f4157b6, 32'h3f09ab50} /* (13, 12, 3) {real, imag} */,
  {32'h3fa22d3a, 32'hbf02b93c} /* (13, 12, 2) {real, imag} */,
  {32'h3f92acdd, 32'hbfda25d4} /* (13, 12, 1) {real, imag} */,
  {32'hbf09dca9, 32'hbf1f12f8} /* (13, 12, 0) {real, imag} */,
  {32'hbe96423e, 32'hbe1ba500} /* (13, 11, 31) {real, imag} */,
  {32'h3b618d00, 32'hbf1a1b44} /* (13, 11, 30) {real, imag} */,
  {32'h3ec0a216, 32'hbcac25c0} /* (13, 11, 29) {real, imag} */,
  {32'hbeffd746, 32'hbe3c6f70} /* (13, 11, 28) {real, imag} */,
  {32'hbd812578, 32'hbf5063c0} /* (13, 11, 27) {real, imag} */,
  {32'h3e676ec0, 32'hbd4d3640} /* (13, 11, 26) {real, imag} */,
  {32'hbd8ad010, 32'h3f3aed4c} /* (13, 11, 25) {real, imag} */,
  {32'h3d8e5ff4, 32'h3e606430} /* (13, 11, 24) {real, imag} */,
  {32'hbf338383, 32'h3eb04c8c} /* (13, 11, 23) {real, imag} */,
  {32'hbf8a5d03, 32'h3e866d58} /* (13, 11, 22) {real, imag} */,
  {32'hbe8e0420, 32'hbf1f8670} /* (13, 11, 21) {real, imag} */,
  {32'h3d7e2e60, 32'h3d8fce00} /* (13, 11, 20) {real, imag} */,
  {32'h3e9b42c4, 32'h3ab28000} /* (13, 11, 19) {real, imag} */,
  {32'h3f002000, 32'h3e322320} /* (13, 11, 18) {real, imag} */,
  {32'hbebdcb48, 32'h3d226ca0} /* (13, 11, 17) {real, imag} */,
  {32'hbf7eab7e, 32'hbf910e79} /* (13, 11, 16) {real, imag} */,
  {32'h3f54ff8a, 32'hbf8478ac} /* (13, 11, 15) {real, imag} */,
  {32'h3fc8b817, 32'hbedb0ee4} /* (13, 11, 14) {real, imag} */,
  {32'h38f70000, 32'hbf03dc0c} /* (13, 11, 13) {real, imag} */,
  {32'hbf94dcde, 32'h3e4c7a70} /* (13, 11, 12) {real, imag} */,
  {32'h3e121b60, 32'hbe612838} /* (13, 11, 11) {real, imag} */,
  {32'hbefadeae, 32'hbe1fe170} /* (13, 11, 10) {real, imag} */,
  {32'hbf181e69, 32'h3e0c46c0} /* (13, 11, 9) {real, imag} */,
  {32'h3f889c7a, 32'h3e980b78} /* (13, 11, 8) {real, imag} */,
  {32'h3f8bf963, 32'hbef47020} /* (13, 11, 7) {real, imag} */,
  {32'hbf719428, 32'h3f2b7fac} /* (13, 11, 6) {real, imag} */,
  {32'hbd2cbb30, 32'h3fc2100b} /* (13, 11, 5) {real, imag} */,
  {32'h3f1ce9cb, 32'h3f16bc78} /* (13, 11, 4) {real, imag} */,
  {32'h3f7ac96e, 32'h3ed704ac} /* (13, 11, 3) {real, imag} */,
  {32'h3eefc6f0, 32'hbbce5600} /* (13, 11, 2) {real, imag} */,
  {32'h3f13f796, 32'hbeb28450} /* (13, 11, 1) {real, imag} */,
  {32'hbee6b447, 32'h3ecdc8a8} /* (13, 11, 0) {real, imag} */,
  {32'hbf7969bc, 32'hbe8a9017} /* (13, 10, 31) {real, imag} */,
  {32'hbf9f6460, 32'hbedc34e8} /* (13, 10, 30) {real, imag} */,
  {32'hbef26537, 32'h3f296fcd} /* (13, 10, 29) {real, imag} */,
  {32'hbe734234, 32'h3e4c3084} /* (13, 10, 28) {real, imag} */,
  {32'h3edb5909, 32'h3f310473} /* (13, 10, 27) {real, imag} */,
  {32'h3ecca832, 32'hbda3f360} /* (13, 10, 26) {real, imag} */,
  {32'hbf3d1346, 32'hbf0583e8} /* (13, 10, 25) {real, imag} */,
  {32'hbf31e209, 32'hbe70547a} /* (13, 10, 24) {real, imag} */,
  {32'hbed8e0e8, 32'hbe5d7520} /* (13, 10, 23) {real, imag} */,
  {32'hbf268664, 32'hbe22e038} /* (13, 10, 22) {real, imag} */,
  {32'hbf888ac3, 32'hbed057f8} /* (13, 10, 21) {real, imag} */,
  {32'hbe849870, 32'h3efb6ade} /* (13, 10, 20) {real, imag} */,
  {32'h3ec91a6e, 32'h3ed790c0} /* (13, 10, 19) {real, imag} */,
  {32'h3f8f78b2, 32'hbfab290f} /* (13, 10, 18) {real, imag} */,
  {32'h3f8b3794, 32'hbfc188f6} /* (13, 10, 17) {real, imag} */,
  {32'hbf1608f0, 32'hbf8f5b1c} /* (13, 10, 16) {real, imag} */,
  {32'h3eb006f8, 32'h3d0b6308} /* (13, 10, 15) {real, imag} */,
  {32'h3fac69a9, 32'hbdb0a168} /* (13, 10, 14) {real, imag} */,
  {32'h3e09bc92, 32'hbf2deb45} /* (13, 10, 13) {real, imag} */,
  {32'hbf06d8a8, 32'h3e737504} /* (13, 10, 12) {real, imag} */,
  {32'hbcf72040, 32'hbe79a3f4} /* (13, 10, 11) {real, imag} */,
  {32'h3e85e8b7, 32'hbe0de904} /* (13, 10, 10) {real, imag} */,
  {32'h3e0856f4, 32'hbed58fdd} /* (13, 10, 9) {real, imag} */,
  {32'h3f8e895e, 32'hbf2a5fc4} /* (13, 10, 8) {real, imag} */,
  {32'h3fa97452, 32'hbf6dc8ea} /* (13, 10, 7) {real, imag} */,
  {32'hbe42a6e6, 32'h3f2b96c5} /* (13, 10, 6) {real, imag} */,
  {32'h3ee229de, 32'h3fe5ef80} /* (13, 10, 5) {real, imag} */,
  {32'h3f0647c0, 32'h3f41fc74} /* (13, 10, 4) {real, imag} */,
  {32'h3ed4dc22, 32'hbe828150} /* (13, 10, 3) {real, imag} */,
  {32'hbf447e5d, 32'h3eba7f9a} /* (13, 10, 2) {real, imag} */,
  {32'hbf223a7c, 32'h3f6a46af} /* (13, 10, 1) {real, imag} */,
  {32'hbf26cada, 32'h3f328530} /* (13, 10, 0) {real, imag} */,
  {32'hbf87a870, 32'hbe881720} /* (13, 9, 31) {real, imag} */,
  {32'hbfb617a1, 32'h3eb5f618} /* (13, 9, 30) {real, imag} */,
  {32'h3e9b8ed0, 32'h3f834142} /* (13, 9, 29) {real, imag} */,
  {32'h3f579e2e, 32'h3ede43e0} /* (13, 9, 28) {real, imag} */,
  {32'hbeec68f4, 32'h3e896b40} /* (13, 9, 27) {real, imag} */,
  {32'hbf0d735d, 32'h3da45560} /* (13, 9, 26) {real, imag} */,
  {32'hbd5530f0, 32'hbd79af80} /* (13, 9, 25) {real, imag} */,
  {32'hbdd741b0, 32'h3eda13a0} /* (13, 9, 24) {real, imag} */,
  {32'h3f2900ca, 32'h3dcb49e0} /* (13, 9, 23) {real, imag} */,
  {32'h3db77f40, 32'h3f1f4100} /* (13, 9, 22) {real, imag} */,
  {32'hbf738f2e, 32'h3ef992ac} /* (13, 9, 21) {real, imag} */,
  {32'hbf6fb136, 32'h3f52ebe4} /* (13, 9, 20) {real, imag} */,
  {32'hbf522788, 32'h3e67f6c0} /* (13, 9, 19) {real, imag} */,
  {32'h3f5494e2, 32'hbfc24b39} /* (13, 9, 18) {real, imag} */,
  {32'h3f96d2e5, 32'hbf6a7d44} /* (13, 9, 17) {real, imag} */,
  {32'hbe0420c0, 32'h3ec4e470} /* (13, 9, 16) {real, imag} */,
  {32'hbf3e8c0b, 32'h3eedc9f0} /* (13, 9, 15) {real, imag} */,
  {32'h3eb290d2, 32'h3ed3fd56} /* (13, 9, 14) {real, imag} */,
  {32'h3ee6a014, 32'hbebf1730} /* (13, 9, 13) {real, imag} */,
  {32'h3ef85376, 32'hbf58cac0} /* (13, 9, 12) {real, imag} */,
  {32'h3ed1cf6c, 32'hbe46a950} /* (13, 9, 11) {real, imag} */,
  {32'h3f3552d8, 32'h3e1c6b00} /* (13, 9, 10) {real, imag} */,
  {32'h3fb567ef, 32'hbef06a86} /* (13, 9, 9) {real, imag} */,
  {32'h3f5bb6e3, 32'h3e7d6ca0} /* (13, 9, 8) {real, imag} */,
  {32'h3dd9e7b8, 32'hbeb57b90} /* (13, 9, 7) {real, imag} */,
  {32'h3e85317c, 32'hbd473780} /* (13, 9, 6) {real, imag} */,
  {32'h3f3915bf, 32'h3f07670a} /* (13, 9, 5) {real, imag} */,
  {32'hbdf930b0, 32'h3e8c5d18} /* (13, 9, 4) {real, imag} */,
  {32'hbe648c38, 32'hbf0547e8} /* (13, 9, 3) {real, imag} */,
  {32'hbeee3a30, 32'hbcb48380} /* (13, 9, 2) {real, imag} */,
  {32'hbf5a9098, 32'h3f56945a} /* (13, 9, 1) {real, imag} */,
  {32'hbf0b710f, 32'h3e9ce8a0} /* (13, 9, 0) {real, imag} */,
  {32'hbf7893e6, 32'hbf1afcd4} /* (13, 8, 31) {real, imag} */,
  {32'hbf51ab84, 32'hbe9cdb88} /* (13, 8, 30) {real, imag} */,
  {32'h3f7b6bce, 32'h3f05d948} /* (13, 8, 29) {real, imag} */,
  {32'h3ed71b26, 32'h3f8ce4c2} /* (13, 8, 28) {real, imag} */,
  {32'hbeddf6e8, 32'hbe208e60} /* (13, 8, 27) {real, imag} */,
  {32'hbf3f7236, 32'hbe9a8330} /* (13, 8, 26) {real, imag} */,
  {32'hbe9bc580, 32'h3eb1f7b8} /* (13, 8, 25) {real, imag} */,
  {32'hbe761010, 32'h3ebeee50} /* (13, 8, 24) {real, imag} */,
  {32'h3db41dd0, 32'h3f4f3938} /* (13, 8, 23) {real, imag} */,
  {32'h3f306fc0, 32'h3f8733de} /* (13, 8, 22) {real, imag} */,
  {32'h3f0da988, 32'h3da8b990} /* (13, 8, 21) {real, imag} */,
  {32'hbc6e0740, 32'h3d1afd00} /* (13, 8, 20) {real, imag} */,
  {32'hbf14bce9, 32'h3e9cd910} /* (13, 8, 19) {real, imag} */,
  {32'h3d54f9a0, 32'h3d15bcc0} /* (13, 8, 18) {real, imag} */,
  {32'h3f071d8d, 32'h3f039188} /* (13, 8, 17) {real, imag} */,
  {32'h3d92bb00, 32'h3f66f428} /* (13, 8, 16) {real, imag} */,
  {32'hbea1b10e, 32'h3e3529e0} /* (13, 8, 15) {real, imag} */,
  {32'h3d64bb80, 32'h3f0f0ec0} /* (13, 8, 14) {real, imag} */,
  {32'hbe7bf978, 32'h3ed974f0} /* (13, 8, 13) {real, imag} */,
  {32'hbf10b5ee, 32'h3eb6e660} /* (13, 8, 12) {real, imag} */,
  {32'hbf4b1f86, 32'h3f258ac8} /* (13, 8, 11) {real, imag} */,
  {32'hbdeb0a18, 32'h3ea63e72} /* (13, 8, 10) {real, imag} */,
  {32'h3e8a3a18, 32'hbe7f6968} /* (13, 8, 9) {real, imag} */,
  {32'hbcd14b40, 32'h3eb911a8} /* (13, 8, 8) {real, imag} */,
  {32'hbe7b1e38, 32'h3cc49900} /* (13, 8, 7) {real, imag} */,
  {32'hbc568f80, 32'hbea66b40} /* (13, 8, 6) {real, imag} */,
  {32'h3e1893a0, 32'h3f012964} /* (13, 8, 5) {real, imag} */,
  {32'h3e1f6cbc, 32'h3ee2b2d8} /* (13, 8, 4) {real, imag} */,
  {32'hbe5e91b0, 32'hbeeb9ea0} /* (13, 8, 3) {real, imag} */,
  {32'hbf061a92, 32'hbe99fe70} /* (13, 8, 2) {real, imag} */,
  {32'hbf1e401f, 32'h3ed3bdc8} /* (13, 8, 1) {real, imag} */,
  {32'hbe659a78, 32'hbba79500} /* (13, 8, 0) {real, imag} */,
  {32'hbe2abfdc, 32'hbf38d5b2} /* (13, 7, 31) {real, imag} */,
  {32'hbe4813a8, 32'hbe88d1dc} /* (13, 7, 30) {real, imag} */,
  {32'h3e17a20c, 32'hbead3648} /* (13, 7, 29) {real, imag} */,
  {32'hbe418894, 32'h3f426764} /* (13, 7, 28) {real, imag} */,
  {32'hbde90858, 32'h3eb09a00} /* (13, 7, 27) {real, imag} */,
  {32'hbc009980, 32'h3e396fc0} /* (13, 7, 26) {real, imag} */,
  {32'h3c124a80, 32'hbe287c60} /* (13, 7, 25) {real, imag} */,
  {32'hbf50a65a, 32'hbfa337be} /* (13, 7, 24) {real, imag} */,
  {32'hbf468a4c, 32'h3dd2c9c0} /* (13, 7, 23) {real, imag} */,
  {32'h3e998598, 32'hbd32a320} /* (13, 7, 22) {real, imag} */,
  {32'h3f0447e9, 32'hbec8fb5e} /* (13, 7, 21) {real, imag} */,
  {32'h3f89a928, 32'h3e963aa8} /* (13, 7, 20) {real, imag} */,
  {32'h3e515490, 32'hbe3f5ee8} /* (13, 7, 19) {real, imag} */,
  {32'hbe8581e4, 32'hbe2f0d70} /* (13, 7, 18) {real, imag} */,
  {32'h3e00b524, 32'h3d75cc80} /* (13, 7, 17) {real, imag} */,
  {32'hbf139d55, 32'h3dbf05e0} /* (13, 7, 16) {real, imag} */,
  {32'hbf1b75f2, 32'h3e8e1ea0} /* (13, 7, 15) {real, imag} */,
  {32'hbf6da79a, 32'h3eb99aa8} /* (13, 7, 14) {real, imag} */,
  {32'hbf01744c, 32'h3edf8d80} /* (13, 7, 13) {real, imag} */,
  {32'h3ef35ff2, 32'h3f709fb4} /* (13, 7, 12) {real, imag} */,
  {32'hbde0dc40, 32'h3f708de4} /* (13, 7, 11) {real, imag} */,
  {32'hbeeecbd0, 32'h3f94f7c8} /* (13, 7, 10) {real, imag} */,
  {32'hbf10a0b0, 32'h3f33a268} /* (13, 7, 9) {real, imag} */,
  {32'h3e9b867a, 32'hbe27add0} /* (13, 7, 8) {real, imag} */,
  {32'hbeb8f2e7, 32'hbf567652} /* (13, 7, 7) {real, imag} */,
  {32'hbf1d72f4, 32'hbf2f23ae} /* (13, 7, 6) {real, imag} */,
  {32'hbef506bc, 32'h3e0ab2e0} /* (13, 7, 5) {real, imag} */,
  {32'h3e759294, 32'h3e749c10} /* (13, 7, 4) {real, imag} */,
  {32'hbe8e3f24, 32'hbee69690} /* (13, 7, 3) {real, imag} */,
  {32'hbe6ded90, 32'hbda52e00} /* (13, 7, 2) {real, imag} */,
  {32'h3e0f52d8, 32'h3eaab838} /* (13, 7, 1) {real, imag} */,
  {32'hbcccdcb0, 32'hbef8aa18} /* (13, 7, 0) {real, imag} */,
  {32'hbf2bbdde, 32'h3cf89540} /* (13, 6, 31) {real, imag} */,
  {32'hbee5e5b8, 32'h3e46c1b0} /* (13, 6, 30) {real, imag} */,
  {32'hbf76f487, 32'hbe7cf620} /* (13, 6, 29) {real, imag} */,
  {32'hbfc57708, 32'hbe829758} /* (13, 6, 28) {real, imag} */,
  {32'hbf9640a2, 32'hbdcd3780} /* (13, 6, 27) {real, imag} */,
  {32'h3ed11f18, 32'hbdf72380} /* (13, 6, 26) {real, imag} */,
  {32'h3f24bb54, 32'hbeeba8b8} /* (13, 6, 25) {real, imag} */,
  {32'hbf262344, 32'hbf95dbf2} /* (13, 6, 24) {real, imag} */,
  {32'hbf5406dc, 32'h3e3af4b0} /* (13, 6, 23) {real, imag} */,
  {32'h3ead9148, 32'h3df49e70} /* (13, 6, 22) {real, imag} */,
  {32'h3fa0e386, 32'hbeb5bc6d} /* (13, 6, 21) {real, imag} */,
  {32'h3f95b15c, 32'hbd9a8090} /* (13, 6, 20) {real, imag} */,
  {32'hbcd89dc0, 32'h3e852ccc} /* (13, 6, 19) {real, imag} */,
  {32'h3d396d48, 32'h3ea73b24} /* (13, 6, 18) {real, imag} */,
  {32'hbd1c9a58, 32'h3e409580} /* (13, 6, 17) {real, imag} */,
  {32'hbf53df21, 32'hbed3b910} /* (13, 6, 16) {real, imag} */,
  {32'hbf01038c, 32'hbef7b7d0} /* (13, 6, 15) {real, imag} */,
  {32'hbf2ccc31, 32'h3e51c340} /* (13, 6, 14) {real, imag} */,
  {32'hbefe24d0, 32'hbe1b59b0} /* (13, 6, 13) {real, imag} */,
  {32'h3f9b64cd, 32'h3e3c6bf0} /* (13, 6, 12) {real, imag} */,
  {32'h3f756b93, 32'hbf18be88} /* (13, 6, 11) {real, imag} */,
  {32'hbcf59100, 32'h3d3ac740} /* (13, 6, 10) {real, imag} */,
  {32'hbe446830, 32'hbe0c7230} /* (13, 6, 9) {real, imag} */,
  {32'hbebbeb68, 32'hbf3ba492} /* (13, 6, 8) {real, imag} */,
  {32'hbf8b7fdb, 32'hbf919041} /* (13, 6, 7) {real, imag} */,
  {32'hbf31967a, 32'hbf2efa9c} /* (13, 6, 6) {real, imag} */,
  {32'hbe601ff0, 32'h3f2215c8} /* (13, 6, 5) {real, imag} */,
  {32'hbf2ee0df, 32'h3ec5dfe0} /* (13, 6, 4) {real, imag} */,
  {32'h3eeb2d02, 32'h3da93020} /* (13, 6, 3) {real, imag} */,
  {32'h3fcb9c4d, 32'h3e899d60} /* (13, 6, 2) {real, imag} */,
  {32'h3f900988, 32'h3f985a42} /* (13, 6, 1) {real, imag} */,
  {32'h3da5d2e8, 32'h3e972e6c} /* (13, 6, 0) {real, imag} */,
  {32'hbf978b34, 32'hbedb59b4} /* (13, 5, 31) {real, imag} */,
  {32'hbed212b8, 32'hbe90d34c} /* (13, 5, 30) {real, imag} */,
  {32'hbf1494c8, 32'h3e52e0b0} /* (13, 5, 29) {real, imag} */,
  {32'hbfa8dc4b, 32'h3ddc8220} /* (13, 5, 28) {real, imag} */,
  {32'hbf482918, 32'hbf3e0420} /* (13, 5, 27) {real, imag} */,
  {32'h3f91690c, 32'hbd4db700} /* (13, 5, 26) {real, imag} */,
  {32'h3f692ee6, 32'hbef60e60} /* (13, 5, 25) {real, imag} */,
  {32'hbe805e74, 32'hbf272cc0} /* (13, 5, 24) {real, imag} */,
  {32'hbe3fd3a8, 32'h3f1986ec} /* (13, 5, 23) {real, imag} */,
  {32'h3e848a78, 32'h3f3b86d4} /* (13, 5, 22) {real, imag} */,
  {32'h3f3b2749, 32'hbe68cd50} /* (13, 5, 21) {real, imag} */,
  {32'h3e2b0238, 32'hbd7d8600} /* (13, 5, 20) {real, imag} */,
  {32'hbf91aaa6, 32'h3e54fde8} /* (13, 5, 19) {real, imag} */,
  {32'hbeb6a6a6, 32'hbeeee3e2} /* (13, 5, 18) {real, imag} */,
  {32'hbe484420, 32'hbe854730} /* (13, 5, 17) {real, imag} */,
  {32'hbeca0381, 32'hbf5d70f5} /* (13, 5, 16) {real, imag} */,
  {32'hbd9802c8, 32'hbe77cda0} /* (13, 5, 15) {real, imag} */,
  {32'h3e8e7de0, 32'h3eba2a00} /* (13, 5, 14) {real, imag} */,
  {32'hbec275bc, 32'hbed55db0} /* (13, 5, 13) {real, imag} */,
  {32'hbeb420f8, 32'h3d567100} /* (13, 5, 12) {real, imag} */,
  {32'h3f3dac9e, 32'hbe33ef40} /* (13, 5, 11) {real, imag} */,
  {32'h3ef3aaf8, 32'h3e616354} /* (13, 5, 10) {real, imag} */,
  {32'hbd8c4a64, 32'hbe159ff0} /* (13, 5, 9) {real, imag} */,
  {32'h3c0c1e40, 32'h3f08b43a} /* (13, 5, 8) {real, imag} */,
  {32'hbecb0edc, 32'h3e8a68aa} /* (13, 5, 7) {real, imag} */,
  {32'h3e1d008a, 32'h3f100f77} /* (13, 5, 6) {real, imag} */,
  {32'h3ee143b0, 32'hbd83ff80} /* (13, 5, 5) {real, imag} */,
  {32'h3ec40464, 32'hbea51e30} /* (13, 5, 4) {real, imag} */,
  {32'h3ef2ffb4, 32'h3f0201c6} /* (13, 5, 3) {real, imag} */,
  {32'h3fcf92e3, 32'h3f325374} /* (13, 5, 2) {real, imag} */,
  {32'h3f4bbce8, 32'h3f83ec84} /* (13, 5, 1) {real, imag} */,
  {32'hbe82ee3d, 32'h3d43e680} /* (13, 5, 0) {real, imag} */,
  {32'hbf91f375, 32'hbe84df84} /* (13, 4, 31) {real, imag} */,
  {32'hbee4c450, 32'h3da683a0} /* (13, 4, 30) {real, imag} */,
  {32'hbe5617d8, 32'h3e7b01f0} /* (13, 4, 29) {real, imag} */,
  {32'hbf0d66a6, 32'hbd1e1380} /* (13, 4, 28) {real, imag} */,
  {32'hbf118eab, 32'h3e671080} /* (13, 4, 27) {real, imag} */,
  {32'h3e429910, 32'h3f2966b0} /* (13, 4, 26) {real, imag} */,
  {32'h3f143be2, 32'h3ea43a08} /* (13, 4, 25) {real, imag} */,
  {32'h3f37b048, 32'hbea888e8} /* (13, 4, 24) {real, imag} */,
  {32'h3eaab6f8, 32'h3ea73ad8} /* (13, 4, 23) {real, imag} */,
  {32'hbf1ed2b1, 32'hbdc92a20} /* (13, 4, 22) {real, imag} */,
  {32'h3dedc628, 32'hbf96e647} /* (13, 4, 21) {real, imag} */,
  {32'h3f0e608b, 32'hbd8a1280} /* (13, 4, 20) {real, imag} */,
  {32'hbef6c60b, 32'h3ec63418} /* (13, 4, 19) {real, imag} */,
  {32'hbeaf1eb3, 32'hbee85a10} /* (13, 4, 18) {real, imag} */,
  {32'hbd4ccea8, 32'hbfa35848} /* (13, 4, 17) {real, imag} */,
  {32'hbe3f8bec, 32'hbfce0ead} /* (13, 4, 16) {real, imag} */,
  {32'h3ef4f1a2, 32'h3ede8f20} /* (13, 4, 15) {real, imag} */,
  {32'h3f81d833, 32'h3f62f90e} /* (13, 4, 14) {real, imag} */,
  {32'hbe271048, 32'h3d430a40} /* (13, 4, 13) {real, imag} */,
  {32'hbe55cac8, 32'h3eb0c950} /* (13, 4, 12) {real, imag} */,
  {32'h3e8a7844, 32'h3e83b8a0} /* (13, 4, 11) {real, imag} */,
  {32'h3f2ad366, 32'h3e69d650} /* (13, 4, 10) {real, imag} */,
  {32'h3f9b9dc2, 32'h3f5fb50c} /* (13, 4, 9) {real, imag} */,
  {32'h3fd55504, 32'h3fc53aed} /* (13, 4, 8) {real, imag} */,
  {32'h3f66ad40, 32'h3ec3fb28} /* (13, 4, 7) {real, imag} */,
  {32'h3f0a35aa, 32'hbe1aeca0} /* (13, 4, 6) {real, imag} */,
  {32'hbe704b70, 32'hbe9a6df7} /* (13, 4, 5) {real, imag} */,
  {32'h3ea6ce9e, 32'hbe3286f8} /* (13, 4, 4) {real, imag} */,
  {32'h3fb0a432, 32'h3ca5b900} /* (13, 4, 3) {real, imag} */,
  {32'h3fa873ef, 32'h3e907438} /* (13, 4, 2) {real, imag} */,
  {32'h3f0cdbd7, 32'hbe0b2b10} /* (13, 4, 1) {real, imag} */,
  {32'hbe21ef60, 32'hbe9efd54} /* (13, 4, 0) {real, imag} */,
  {32'hbedaff8c, 32'h3ef979a0} /* (13, 3, 31) {real, imag} */,
  {32'hbe0c16b0, 32'h3f337e04} /* (13, 3, 30) {real, imag} */,
  {32'hbe6c7914, 32'h3d4a7d80} /* (13, 3, 29) {real, imag} */,
  {32'hbf6eb755, 32'hbf3e39c8} /* (13, 3, 28) {real, imag} */,
  {32'hbfc43634, 32'hbe5b8ee0} /* (13, 3, 27) {real, imag} */,
  {32'hbf5c5cbe, 32'hbec0f450} /* (13, 3, 26) {real, imag} */,
  {32'hbf214bac, 32'h3d0d9880} /* (13, 3, 25) {real, imag} */,
  {32'h3d7a7240, 32'hbecf11c0} /* (13, 3, 24) {real, imag} */,
  {32'h3ce69460, 32'h3e171d40} /* (13, 3, 23) {real, imag} */,
  {32'hbdfd9ce0, 32'h3c5889c0} /* (13, 3, 22) {real, imag} */,
  {32'h3ef2bcbb, 32'hbef5a488} /* (13, 3, 21) {real, imag} */,
  {32'h3d8d68a0, 32'h3e841cd0} /* (13, 3, 20) {real, imag} */,
  {32'h3e2b2270, 32'h3e5736b0} /* (13, 3, 19) {real, imag} */,
  {32'hbd859fe0, 32'h3f5fd0ce} /* (13, 3, 18) {real, imag} */,
  {32'hbc559880, 32'hbe0b0380} /* (13, 3, 17) {real, imag} */,
  {32'hbf28e226, 32'h3e7ffb80} /* (13, 3, 16) {real, imag} */,
  {32'hbea6a77d, 32'h3f90110b} /* (13, 3, 15) {real, imag} */,
  {32'h3f164f27, 32'h3fc78472} /* (13, 3, 14) {real, imag} */,
  {32'h3f6c8c4f, 32'h3fa82216} /* (13, 3, 13) {real, imag} */,
  {32'h3f8d4602, 32'h3fc62084} /* (13, 3, 12) {real, imag} */,
  {32'h3f8b8ec0, 32'h3f25d454} /* (13, 3, 11) {real, imag} */,
  {32'h3f9c8b5b, 32'h3d849660} /* (13, 3, 10) {real, imag} */,
  {32'h3fb0dabf, 32'h3fa744e4} /* (13, 3, 9) {real, imag} */,
  {32'h3f51bbfb, 32'h3fbd2d98} /* (13, 3, 8) {real, imag} */,
  {32'hbec2650d, 32'h3e661350} /* (13, 3, 7) {real, imag} */,
  {32'hbde8e9f8, 32'hbf0bf340} /* (13, 3, 6) {real, imag} */,
  {32'hbe6fc290, 32'hbd2638e0} /* (13, 3, 5) {real, imag} */,
  {32'h3e352088, 32'hbe2c13bc} /* (13, 3, 4) {real, imag} */,
  {32'h3f102f70, 32'hbdac9e00} /* (13, 3, 3) {real, imag} */,
  {32'h3e2c4160, 32'hbdbae180} /* (13, 3, 2) {real, imag} */,
  {32'hbe793c88, 32'hbe55dba0} /* (13, 3, 1) {real, imag} */,
  {32'hbdbb6490, 32'h3e900f10} /* (13, 3, 0) {real, imag} */,
  {32'hbe9d3118, 32'h3f918558} /* (13, 2, 31) {real, imag} */,
  {32'hbec687e0, 32'h3f7e1918} /* (13, 2, 30) {real, imag} */,
  {32'hbeb3c5e4, 32'h3dc1c860} /* (13, 2, 29) {real, imag} */,
  {32'hbd0eade0, 32'h3e8c8368} /* (13, 2, 28) {real, imag} */,
  {32'hbf51a895, 32'hbdd0b1c0} /* (13, 2, 27) {real, imag} */,
  {32'hbe1796f4, 32'hbf6b020c} /* (13, 2, 26) {real, imag} */,
  {32'hbe0b6368, 32'h3e80b4b0} /* (13, 2, 25) {real, imag} */,
  {32'hbf3895a4, 32'h3c1cf300} /* (13, 2, 24) {real, imag} */,
  {32'hbef0c7e0, 32'hbe5758bc} /* (13, 2, 23) {real, imag} */,
  {32'h3d87dec0, 32'h3f256496} /* (13, 2, 22) {real, imag} */,
  {32'h3f246efc, 32'h3f0befc8} /* (13, 2, 21) {real, imag} */,
  {32'hbdf7e920, 32'h3d327b00} /* (13, 2, 20) {real, imag} */,
  {32'h3f322976, 32'hbf39bd38} /* (13, 2, 19) {real, imag} */,
  {32'hbdd988e8, 32'h3e5a69f8} /* (13, 2, 18) {real, imag} */,
  {32'hbf1c1364, 32'h3ed70848} /* (13, 2, 17) {real, imag} */,
  {32'h3e3ceb00, 32'h3f84370e} /* (13, 2, 16) {real, imag} */,
  {32'h3ecf0888, 32'h3fc7d622} /* (13, 2, 15) {real, imag} */,
  {32'hbcfe0890, 32'h3fdfc1da} /* (13, 2, 14) {real, imag} */,
  {32'hbc11ebc0, 32'h3f4b0a26} /* (13, 2, 13) {real, imag} */,
  {32'h3e465fe0, 32'h3f594458} /* (13, 2, 12) {real, imag} */,
  {32'h3f60c146, 32'h3f2832dc} /* (13, 2, 11) {real, imag} */,
  {32'h3edf0ada, 32'h3f5fb9d8} /* (13, 2, 10) {real, imag} */,
  {32'h3e234950, 32'h3fd92ed0} /* (13, 2, 9) {real, imag} */,
  {32'hbec4f496, 32'h3fafbde4} /* (13, 2, 8) {real, imag} */,
  {32'hbdf8e920, 32'h3ee8c7e0} /* (13, 2, 7) {real, imag} */,
  {32'h3ea742ba, 32'hbfa815bc} /* (13, 2, 6) {real, imag} */,
  {32'hbce2a200, 32'hbf7fdbb6} /* (13, 2, 5) {real, imag} */,
  {32'h3ed86b56, 32'h3df989c0} /* (13, 2, 4) {real, imag} */,
  {32'h3e7f8fb8, 32'hbedae120} /* (13, 2, 3) {real, imag} */,
  {32'h3edbce08, 32'hbf8b8e33} /* (13, 2, 2) {real, imag} */,
  {32'h3f2f5ad2, 32'hbf420fac} /* (13, 2, 1) {real, imag} */,
  {32'h3e1aa728, 32'h3f028624} /* (13, 2, 0) {real, imag} */,
  {32'h3d1f49a0, 32'h3f3dd3f8} /* (13, 1, 31) {real, imag} */,
  {32'h3eb6b0e2, 32'h3f9c084e} /* (13, 1, 30) {real, imag} */,
  {32'h3f2b2f3b, 32'hbc626300} /* (13, 1, 29) {real, imag} */,
  {32'h3ecbd0b1, 32'h3f112b34} /* (13, 1, 28) {real, imag} */,
  {32'hbf3e8e88, 32'h3e6ded80} /* (13, 1, 27) {real, imag} */,
  {32'hbf7dd1b2, 32'hbf06cfb8} /* (13, 1, 26) {real, imag} */,
  {32'hbec8b594, 32'h3e5d8860} /* (13, 1, 25) {real, imag} */,
  {32'hbc366200, 32'h3f0d3d60} /* (13, 1, 24) {real, imag} */,
  {32'h3f1a21d0, 32'hbf6846fe} /* (13, 1, 23) {real, imag} */,
  {32'h3f346400, 32'hbf068f48} /* (13, 1, 22) {real, imag} */,
  {32'h3f3daf1e, 32'h3ecb6160} /* (13, 1, 21) {real, imag} */,
  {32'h3e6ed478, 32'h3eaa2f28} /* (13, 1, 20) {real, imag} */,
  {32'h3f2edb2a, 32'hbeafae98} /* (13, 1, 19) {real, imag} */,
  {32'hbe24f750, 32'h3de51760} /* (13, 1, 18) {real, imag} */,
  {32'hbf80bdff, 32'h3e81bec0} /* (13, 1, 17) {real, imag} */,
  {32'hbd193d80, 32'h3f544eb6} /* (13, 1, 16) {real, imag} */,
  {32'h3e12a718, 32'h3f9034fe} /* (13, 1, 15) {real, imag} */,
  {32'hbf429d45, 32'h3f65a7a4} /* (13, 1, 14) {real, imag} */,
  {32'hbfc4dedd, 32'h3ed9b4d8} /* (13, 1, 13) {real, imag} */,
  {32'hbf591555, 32'hbe70a870} /* (13, 1, 12) {real, imag} */,
  {32'h3dc977d0, 32'hbed66f00} /* (13, 1, 11) {real, imag} */,
  {32'h3e8f8c18, 32'h3ef5b998} /* (13, 1, 10) {real, imag} */,
  {32'h3e40f620, 32'h3f441008} /* (13, 1, 9) {real, imag} */,
  {32'hbe02e360, 32'hbeecfb38} /* (13, 1, 8) {real, imag} */,
  {32'h3f416bda, 32'h3e427710} /* (13, 1, 7) {real, imag} */,
  {32'h3efd76dc, 32'h3dda7440} /* (13, 1, 6) {real, imag} */,
  {32'hbf6c11d3, 32'hbf25ab40} /* (13, 1, 5) {real, imag} */,
  {32'h3d6c5860, 32'hbdd05d40} /* (13, 1, 4) {real, imag} */,
  {32'h3f4eccec, 32'h3e21bf10} /* (13, 1, 3) {real, imag} */,
  {32'h3f51d546, 32'hbe7fbff0} /* (13, 1, 2) {real, imag} */,
  {32'h3f3b23ce, 32'hbefaf10c} /* (13, 1, 1) {real, imag} */,
  {32'h3e2eaff2, 32'h3d849da0} /* (13, 1, 0) {real, imag} */,
  {32'h3d41f408, 32'hbd679090} /* (13, 0, 31) {real, imag} */,
  {32'h3ef2597c, 32'h3ec07288} /* (13, 0, 30) {real, imag} */,
  {32'h3edb83af, 32'hbe8d00dc} /* (13, 0, 29) {real, imag} */,
  {32'h3d1055a0, 32'hbef076dc} /* (13, 0, 28) {real, imag} */,
  {32'hbf491476, 32'hbf34f092} /* (13, 0, 27) {real, imag} */,
  {32'hbf4ab3af, 32'hbf2e4e5e} /* (13, 0, 26) {real, imag} */,
  {32'hbea9fe6e, 32'hbf1ab484} /* (13, 0, 25) {real, imag} */,
  {32'h3f07c6b0, 32'hbefc9818} /* (13, 0, 24) {real, imag} */,
  {32'h3f9cc678, 32'hbf185a0d} /* (13, 0, 23) {real, imag} */,
  {32'h3f92fb65, 32'hbf153080} /* (13, 0, 22) {real, imag} */,
  {32'h3ea4e284, 32'hbe495eb8} /* (13, 0, 21) {real, imag} */,
  {32'hbe062a80, 32'h3dbf24b4} /* (13, 0, 20) {real, imag} */,
  {32'h3cd995e0, 32'hbe867134} /* (13, 0, 19) {real, imag} */,
  {32'h3e7e1bdc, 32'h3e6a1e00} /* (13, 0, 18) {real, imag} */,
  {32'h3d0ba230, 32'h3dc23280} /* (13, 0, 17) {real, imag} */,
  {32'h3bd19100, 32'h3eca805e} /* (13, 0, 16) {real, imag} */,
  {32'h3cb30540, 32'h3ed34720} /* (13, 0, 15) {real, imag} */,
  {32'hbf35e58a, 32'h3d08b180} /* (13, 0, 14) {real, imag} */,
  {32'hbf86d84a, 32'hbddf4cc0} /* (13, 0, 13) {real, imag} */,
  {32'h3e190690, 32'hbec83788} /* (13, 0, 12) {real, imag} */,
  {32'h3d7378e0, 32'hbe6e6b60} /* (13, 0, 11) {real, imag} */,
  {32'h3b116980, 32'hbd0aa398} /* (13, 0, 10) {real, imag} */,
  {32'hbd2e5060, 32'hbe6205c8} /* (13, 0, 9) {real, imag} */,
  {32'h3e98c5f0, 32'hbf2bd6fc} /* (13, 0, 8) {real, imag} */,
  {32'h3f0c7e2e, 32'h3e5957d0} /* (13, 0, 7) {real, imag} */,
  {32'h3ecddb4c, 32'h3f486f2d} /* (13, 0, 6) {real, imag} */,
  {32'hbeb1248c, 32'hbece2e21} /* (13, 0, 5) {real, imag} */,
  {32'hbe118cdf, 32'hbf50e20c} /* (13, 0, 4) {real, imag} */,
  {32'h3f43a64e, 32'h3e235460} /* (13, 0, 3) {real, imag} */,
  {32'h3eb1a8cd, 32'h3e10d4b8} /* (13, 0, 2) {real, imag} */,
  {32'hbcc7bf30, 32'hbec63724} /* (13, 0, 1) {real, imag} */,
  {32'hbec86414, 32'hbf0c8208} /* (13, 0, 0) {real, imag} */,
  {32'hbea9e695, 32'hbe6f9b68} /* (12, 31, 31) {real, imag} */,
  {32'hbe910638, 32'h3e3d1720} /* (12, 31, 30) {real, imag} */,
  {32'hbf1680c0, 32'h3ebe7240} /* (12, 31, 29) {real, imag} */,
  {32'hbf2d9604, 32'h3efa8178} /* (12, 31, 28) {real, imag} */,
  {32'hbf7ae8e6, 32'h3dd7d300} /* (12, 31, 27) {real, imag} */,
  {32'h3e836b14, 32'hbf6c9446} /* (12, 31, 26) {real, imag} */,
  {32'h3fa0f739, 32'hbf956bae} /* (12, 31, 25) {real, imag} */,
  {32'h3f8e2b03, 32'hbcb378c0} /* (12, 31, 24) {real, imag} */,
  {32'hbcae3d80, 32'h3f5bbcb6} /* (12, 31, 23) {real, imag} */,
  {32'hbefc9004, 32'h3ebd1818} /* (12, 31, 22) {real, imag} */,
  {32'h3e161c31, 32'hbdd4aae0} /* (12, 31, 21) {real, imag} */,
  {32'hbe307026, 32'hbf041eba} /* (12, 31, 20) {real, imag} */,
  {32'h3e40cf6d, 32'hbef99428} /* (12, 31, 19) {real, imag} */,
  {32'hbe5d9112, 32'hbf0c4bbe} /* (12, 31, 18) {real, imag} */,
  {32'hbf14202a, 32'h3e9416dc} /* (12, 31, 17) {real, imag} */,
  {32'hbf79aedc, 32'h3e323b7a} /* (12, 31, 16) {real, imag} */,
  {32'hbee85e5a, 32'hbdc71b30} /* (12, 31, 15) {real, imag} */,
  {32'h3ef149d2, 32'h3e5c5ef0} /* (12, 31, 14) {real, imag} */,
  {32'hbe913dba, 32'h3ec6bd6c} /* (12, 31, 13) {real, imag} */,
  {32'h3f04d154, 32'hbe311f70} /* (12, 31, 12) {real, imag} */,
  {32'h3e63f78c, 32'h3e086860} /* (12, 31, 11) {real, imag} */,
  {32'h3e49b825, 32'hbeb39fb8} /* (12, 31, 10) {real, imag} */,
  {32'hbd7205e0, 32'hbef781f8} /* (12, 31, 9) {real, imag} */,
  {32'hbf72ce5a, 32'hbea06ba8} /* (12, 31, 8) {real, imag} */,
  {32'hbf61e8ed, 32'h3efbb536} /* (12, 31, 7) {real, imag} */,
  {32'hbea0bfac, 32'h3f05410f} /* (12, 31, 6) {real, imag} */,
  {32'h3e8da598, 32'h3f1be4c4} /* (12, 31, 5) {real, imag} */,
  {32'h3e2e4728, 32'h3dd2af58} /* (12, 31, 4) {real, imag} */,
  {32'hbf65cd10, 32'hbee603d8} /* (12, 31, 3) {real, imag} */,
  {32'hbfa2c183, 32'hbeadd3c8} /* (12, 31, 2) {real, imag} */,
  {32'hbe95dbc0, 32'h3f44e696} /* (12, 31, 1) {real, imag} */,
  {32'h3e20c92c, 32'h3e6f4700} /* (12, 31, 0) {real, imag} */,
  {32'h3e2b92b0, 32'hbf1208f8} /* (12, 30, 31) {real, imag} */,
  {32'h3da3e300, 32'hbf512438} /* (12, 30, 30) {real, imag} */,
  {32'hbde75ce0, 32'hbf3953ac} /* (12, 30, 29) {real, imag} */,
  {32'hbd92b8c0, 32'h3e83dc90} /* (12, 30, 28) {real, imag} */,
  {32'hbf88983c, 32'hbeaaf4d8} /* (12, 30, 27) {real, imag} */,
  {32'h3e8987d6, 32'hbfef51a8} /* (12, 30, 26) {real, imag} */,
  {32'h3fde443d, 32'hbfb732d8} /* (12, 30, 25) {real, imag} */,
  {32'h3fdb9e9a, 32'hbe890888} /* (12, 30, 24) {real, imag} */,
  {32'h3e217078, 32'h3f80e888} /* (12, 30, 23) {real, imag} */,
  {32'hbf157b78, 32'h3ec1ce00} /* (12, 30, 22) {real, imag} */,
  {32'h3f5d14de, 32'h3e25f8c0} /* (12, 30, 21) {real, imag} */,
  {32'h3edf509e, 32'hbf503f78} /* (12, 30, 20) {real, imag} */,
  {32'h3eaddb58, 32'hbea20f88} /* (12, 30, 19) {real, imag} */,
  {32'hbd974b2e, 32'hbcfbab00} /* (12, 30, 18) {real, imag} */,
  {32'hbc8076a0, 32'hbde27960} /* (12, 30, 17) {real, imag} */,
  {32'hbf22b5a2, 32'hbf130180} /* (12, 30, 16) {real, imag} */,
  {32'hbf10c1fe, 32'h3ec01138} /* (12, 30, 15) {real, imag} */,
  {32'h3e15e158, 32'h3fe8a7f4} /* (12, 30, 14) {real, imag} */,
  {32'hbe45747f, 32'h3f98613d} /* (12, 30, 13) {real, imag} */,
  {32'h3f5a307c, 32'h3e8f1db0} /* (12, 30, 12) {real, imag} */,
  {32'h3ec0060c, 32'h3e8d6fe0} /* (12, 30, 11) {real, imag} */,
  {32'h3f69a261, 32'hbecd548d} /* (12, 30, 10) {real, imag} */,
  {32'h3e819f20, 32'h3db15ae0} /* (12, 30, 9) {real, imag} */,
  {32'hbf651cd0, 32'h3fa2c9e0} /* (12, 30, 8) {real, imag} */,
  {32'hbf8a1ddd, 32'h3fe389e1} /* (12, 30, 7) {real, imag} */,
  {32'hbe4dc264, 32'h3fd3e57e} /* (12, 30, 6) {real, imag} */,
  {32'hbddb6140, 32'h3f96e9b4} /* (12, 30, 5) {real, imag} */,
  {32'hbe8f79ac, 32'h3da33540} /* (12, 30, 4) {real, imag} */,
  {32'hbf4fb8d8, 32'hbd233040} /* (12, 30, 3) {real, imag} */,
  {32'hbf9ea86d, 32'h3ea5e7a0} /* (12, 30, 2) {real, imag} */,
  {32'h3ea0de94, 32'h3edfc538} /* (12, 30, 1) {real, imag} */,
  {32'h3f20382e, 32'hbe9de794} /* (12, 30, 0) {real, imag} */,
  {32'h3f06605e, 32'h3e3456a8} /* (12, 29, 31) {real, imag} */,
  {32'h3e7590b8, 32'hbf94dd3c} /* (12, 29, 30) {real, imag} */,
  {32'hbeca0f84, 32'hbfd189eb} /* (12, 29, 29) {real, imag} */,
  {32'hbf9a3e50, 32'hbe653380} /* (12, 29, 28) {real, imag} */,
  {32'hbf210892, 32'h3e1226a0} /* (12, 29, 27) {real, imag} */,
  {32'h3f2463c8, 32'hbee73988} /* (12, 29, 26) {real, imag} */,
  {32'h3f11f2f2, 32'hbf6a7362} /* (12, 29, 25) {real, imag} */,
  {32'h3f33140c, 32'hbf5ddb74} /* (12, 29, 24) {real, imag} */,
  {32'h3d860390, 32'h3e9bdfb8} /* (12, 29, 23) {real, imag} */,
  {32'h3ef5d8c6, 32'h3f57ee90} /* (12, 29, 22) {real, imag} */,
  {32'h3fe9304b, 32'h3f016e74} /* (12, 29, 21) {real, imag} */,
  {32'h3fb1a026, 32'hbfa3f600} /* (12, 29, 20) {real, imag} */,
  {32'h3f89ba36, 32'hbf352474} /* (12, 29, 19) {real, imag} */,
  {32'h3ef60132, 32'hbbc3d200} /* (12, 29, 18) {real, imag} */,
  {32'hbc9df500, 32'hbf249564} /* (12, 29, 17) {real, imag} */,
  {32'h3ee3664a, 32'hbbd5be00} /* (12, 29, 16) {real, imag} */,
  {32'h3e8e14fa, 32'hbd5db900} /* (12, 29, 15) {real, imag} */,
  {32'h3ee2f1a0, 32'h3ecab4a0} /* (12, 29, 14) {real, imag} */,
  {32'h3f2800f6, 32'h3cd3bc00} /* (12, 29, 13) {real, imag} */,
  {32'h3fcbc7b7, 32'hbf20eef8} /* (12, 29, 12) {real, imag} */,
  {32'h3f80d36f, 32'hbee036fc} /* (12, 29, 11) {real, imag} */,
  {32'h3fb59e1c, 32'h3efd2b82} /* (12, 29, 10) {real, imag} */,
  {32'h3f3f07dc, 32'h3f1babb0} /* (12, 29, 9) {real, imag} */,
  {32'h3ece9af8, 32'h3f9befa0} /* (12, 29, 8) {real, imag} */,
  {32'hbf788c54, 32'h3fabf3d2} /* (12, 29, 7) {real, imag} */,
  {32'hbf9be379, 32'h3f57ffee} /* (12, 29, 6) {real, imag} */,
  {32'hbf3f901e, 32'h3f9935c8} /* (12, 29, 5) {real, imag} */,
  {32'hbf22602e, 32'h3e25da90} /* (12, 29, 4) {real, imag} */,
  {32'hbfccc134, 32'hbe363c10} /* (12, 29, 3) {real, imag} */,
  {32'hbf49433e, 32'h3f7e215a} /* (12, 29, 2) {real, imag} */,
  {32'h3f0c9a27, 32'h3f544ec6} /* (12, 29, 1) {real, imag} */,
  {32'h3f255ac6, 32'h3ed51b0c} /* (12, 29, 0) {real, imag} */,
  {32'hbe5defa8, 32'h3dba2384} /* (12, 28, 31) {real, imag} */,
  {32'hbe28e640, 32'hbf810032} /* (12, 28, 30) {real, imag} */,
  {32'hbf2c6330, 32'hbf5c2378} /* (12, 28, 29) {real, imag} */,
  {32'hbfd0af34, 32'h3f25e12c} /* (12, 28, 28) {real, imag} */,
  {32'hbe84ee90, 32'h3f135ebc} /* (12, 28, 27) {real, imag} */,
  {32'h3e35c788, 32'hbec16bd0} /* (12, 28, 26) {real, imag} */,
  {32'h3f024590, 32'hbe9ccaa8} /* (12, 28, 25) {real, imag} */,
  {32'h3cb31f60, 32'h3da76540} /* (12, 28, 24) {real, imag} */,
  {32'hbf4d7ede, 32'h3e34c020} /* (12, 28, 23) {real, imag} */,
  {32'hbefe0908, 32'h3f196ef0} /* (12, 28, 22) {real, imag} */,
  {32'h3f813959, 32'h3f1ac8a4} /* (12, 28, 21) {real, imag} */,
  {32'h3f9091e8, 32'hbef3a650} /* (12, 28, 20) {real, imag} */,
  {32'h3f6f666a, 32'hbef1d234} /* (12, 28, 19) {real, imag} */,
  {32'h3ee4a708, 32'h3e8fe9e8} /* (12, 28, 18) {real, imag} */,
  {32'h3e539920, 32'h3f4a1ea0} /* (12, 28, 17) {real, imag} */,
  {32'h3f2b669c, 32'h3f022ab8} /* (12, 28, 16) {real, imag} */,
  {32'h3eb72d64, 32'hbf39e6e2} /* (12, 28, 15) {real, imag} */,
  {32'h3e072ad0, 32'h3ea1509c} /* (12, 28, 14) {real, imag} */,
  {32'h3ec5d548, 32'hbdbda850} /* (12, 28, 13) {real, imag} */,
  {32'h3f8c902b, 32'hbeef2044} /* (12, 28, 12) {real, imag} */,
  {32'h3dd936d9, 32'h3f255ef6} /* (12, 28, 11) {real, imag} */,
  {32'hbe7f5050, 32'h3c3c6c00} /* (12, 28, 10) {real, imag} */,
  {32'h3d36e440, 32'hbfab0c87} /* (12, 28, 9) {real, imag} */,
  {32'h3f447798, 32'hbf7333f4} /* (12, 28, 8) {real, imag} */,
  {32'hbe272da8, 32'hbcba8500} /* (12, 28, 7) {real, imag} */,
  {32'hbef04a70, 32'hbdd51320} /* (12, 28, 6) {real, imag} */,
  {32'h3ddb3b30, 32'h3e920974} /* (12, 28, 5) {real, imag} */,
  {32'hbf08ceec, 32'hbea05314} /* (12, 28, 4) {real, imag} */,
  {32'hbfced17a, 32'hbfa4821f} /* (12, 28, 3) {real, imag} */,
  {32'h3d586880, 32'hbf1115e2} /* (12, 28, 2) {real, imag} */,
  {32'hbdca22c0, 32'h3f78b8f0} /* (12, 28, 1) {real, imag} */,
  {32'hbe860913, 32'h3f806796} /* (12, 28, 0) {real, imag} */,
  {32'hbdb35d2c, 32'hbd4a32e0} /* (12, 27, 31) {real, imag} */,
  {32'h3dbf2480, 32'hbf765da0} /* (12, 27, 30) {real, imag} */,
  {32'h3e1d5e50, 32'hbf04d628} /* (12, 27, 29) {real, imag} */,
  {32'h3f0863b2, 32'h3e628268} /* (12, 27, 28) {real, imag} */,
  {32'h3efc39dc, 32'h3f0867e0} /* (12, 27, 27) {real, imag} */,
  {32'hbe6b4550, 32'hbf273710} /* (12, 27, 26) {real, imag} */,
  {32'hbeb0f567, 32'hbd09d780} /* (12, 27, 25) {real, imag} */,
  {32'hbf064090, 32'h3d853050} /* (12, 27, 24) {real, imag} */,
  {32'h3e83a05c, 32'h3ed28f90} /* (12, 27, 23) {real, imag} */,
  {32'h3d596a00, 32'h3eae02a8} /* (12, 27, 22) {real, imag} */,
  {32'h3ef73d84, 32'h3d9de840} /* (12, 27, 21) {real, imag} */,
  {32'h3f4237ee, 32'hbf32cc5a} /* (12, 27, 20) {real, imag} */,
  {32'hbe5f3dd0, 32'hbf17c366} /* (12, 27, 19) {real, imag} */,
  {32'hbf7626f0, 32'hbeb4aabc} /* (12, 27, 18) {real, imag} */,
  {32'hbf6a9358, 32'hbf72af46} /* (12, 27, 17) {real, imag} */,
  {32'hbd9534b0, 32'hbeeaf778} /* (12, 27, 16) {real, imag} */,
  {32'hbcb203a0, 32'hbf97651e} /* (12, 27, 15) {real, imag} */,
  {32'hbea23d8c, 32'h3ee03230} /* (12, 27, 14) {real, imag} */,
  {32'h3b870880, 32'h3f1b8eec} /* (12, 27, 13) {real, imag} */,
  {32'h3ec1a6e9, 32'h3ecb4c50} /* (12, 27, 12) {real, imag} */,
  {32'hbe8bc558, 32'h3fe249c5} /* (12, 27, 11) {real, imag} */,
  {32'hbe826d54, 32'h3f1ba740} /* (12, 27, 10) {real, imag} */,
  {32'h3f21f38e, 32'h3ebcc0f8} /* (12, 27, 9) {real, imag} */,
  {32'h3f7292b8, 32'hbe47c450} /* (12, 27, 8) {real, imag} */,
  {32'h3f6474d0, 32'hbf684e04} /* (12, 27, 7) {real, imag} */,
  {32'h3dda6ef0, 32'hbf845e22} /* (12, 27, 6) {real, imag} */,
  {32'hbe117500, 32'h3da81fc0} /* (12, 27, 5) {real, imag} */,
  {32'h3f0e154c, 32'h3e764b38} /* (12, 27, 4) {real, imag} */,
  {32'h3eecd5b8, 32'hbe7643f0} /* (12, 27, 3) {real, imag} */,
  {32'h3e8ac608, 32'hbf9d9aad} /* (12, 27, 2) {real, imag} */,
  {32'hbf234a02, 32'h3d2639a0} /* (12, 27, 1) {real, imag} */,
  {32'hbf0869aa, 32'h3f02339a} /* (12, 27, 0) {real, imag} */,
  {32'h3e3b6d04, 32'hbf17f480} /* (12, 26, 31) {real, imag} */,
  {32'h3e7ef6f0, 32'hbf975ca1} /* (12, 26, 30) {real, imag} */,
  {32'h3f30514e, 32'hbe35e7d0} /* (12, 26, 29) {real, imag} */,
  {32'h3f45f342, 32'hbf5d2864} /* (12, 26, 28) {real, imag} */,
  {32'hbed5a130, 32'hbf380f52} /* (12, 26, 27) {real, imag} */,
  {32'hbe2292c0, 32'hbe523230} /* (12, 26, 26) {real, imag} */,
  {32'hbeae5f40, 32'hbd957da0} /* (12, 26, 25) {real, imag} */,
  {32'hbf844be5, 32'hbf20a9e5} /* (12, 26, 24) {real, imag} */,
  {32'h3f087f76, 32'h3f1479d0} /* (12, 26, 23) {real, imag} */,
  {32'hbc08f380, 32'h3f3af7ea} /* (12, 26, 22) {real, imag} */,
  {32'hbf8aeeea, 32'hbedf2d64} /* (12, 26, 21) {real, imag} */,
  {32'h3ececc42, 32'hbe777f18} /* (12, 26, 20) {real, imag} */,
  {32'h3f3c00f0, 32'h3df07370} /* (12, 26, 19) {real, imag} */,
  {32'h3e471aa8, 32'hbe6255e0} /* (12, 26, 18) {real, imag} */,
  {32'h3eca38e2, 32'hbf8f210d} /* (12, 26, 17) {real, imag} */,
  {32'h3f2d9408, 32'hbf3d569e} /* (12, 26, 16) {real, imag} */,
  {32'hbe33edee, 32'hbe811da8} /* (12, 26, 15) {real, imag} */,
  {32'hbf08a59a, 32'h3f2da52c} /* (12, 26, 14) {real, imag} */,
  {32'hbdeb1e68, 32'h3f280684} /* (12, 26, 13) {real, imag} */,
  {32'h3ca54b18, 32'h3f4e3c0e} /* (12, 26, 12) {real, imag} */,
  {32'hbeda1d30, 32'h3f624952} /* (12, 26, 11) {real, imag} */,
  {32'hbde7b3ac, 32'h3dd3b150} /* (12, 26, 10) {real, imag} */,
  {32'hbeed7060, 32'h3fc40704} /* (12, 26, 9) {real, imag} */,
  {32'h3dd29420, 32'h3f5481f0} /* (12, 26, 8) {real, imag} */,
  {32'h3f61d61d, 32'hbf5e60fc} /* (12, 26, 7) {real, imag} */,
  {32'h3dc22428, 32'hbfac1606} /* (12, 26, 6) {real, imag} */,
  {32'h3d4603a0, 32'h3e066500} /* (12, 26, 5) {real, imag} */,
  {32'h3f4b38fd, 32'h3e9ea0d0} /* (12, 26, 4) {real, imag} */,
  {32'h3c8d50c0, 32'hbe98af64} /* (12, 26, 3) {real, imag} */,
  {32'hbea53f4a, 32'hbf3b1650} /* (12, 26, 2) {real, imag} */,
  {32'hbf86b1a8, 32'hbf2a5990} /* (12, 26, 1) {real, imag} */,
  {32'hbf60d0a8, 32'hbe27f3c8} /* (12, 26, 0) {real, imag} */,
  {32'h3e2a8e48, 32'hbecf4ab0} /* (12, 25, 31) {real, imag} */,
  {32'h3e906320, 32'hbfadc49a} /* (12, 25, 30) {real, imag} */,
  {32'hbda66600, 32'h3e4f7788} /* (12, 25, 29) {real, imag} */,
  {32'hbe0d8d40, 32'hbf2367de} /* (12, 25, 28) {real, imag} */,
  {32'hbe33423a, 32'hbf7e4dc4} /* (12, 25, 27) {real, imag} */,
  {32'hbdb302d0, 32'hbef7a010} /* (12, 25, 26) {real, imag} */,
  {32'h3e268838, 32'hbe6d3ea0} /* (12, 25, 25) {real, imag} */,
  {32'hbeefc5c4, 32'hbe87b490} /* (12, 25, 24) {real, imag} */,
  {32'hbe373e68, 32'h3f79fa3c} /* (12, 25, 23) {real, imag} */,
  {32'hbf1f0aa6, 32'h3f87a1b4} /* (12, 25, 22) {real, imag} */,
  {32'hbf8485c8, 32'hbf008ede} /* (12, 25, 21) {real, imag} */,
  {32'hbec431f0, 32'h3f203170} /* (12, 25, 20) {real, imag} */,
  {32'h3f653f87, 32'h3fa4f928} /* (12, 25, 19) {real, imag} */,
  {32'h3f69c3e2, 32'h3e7512d0} /* (12, 25, 18) {real, imag} */,
  {32'h40004fe8, 32'h3e8f317c} /* (12, 25, 17) {real, imag} */,
  {32'h3fcce1e9, 32'h3d92da20} /* (12, 25, 16) {real, imag} */,
  {32'h3e93cabe, 32'hbd37f040} /* (12, 25, 15) {real, imag} */,
  {32'hbf3a8794, 32'h3e27b2a0} /* (12, 25, 14) {real, imag} */,
  {32'hbf3b1a83, 32'hbe37d640} /* (12, 25, 13) {real, imag} */,
  {32'h3d95dc14, 32'h3f77dad8} /* (12, 25, 12) {real, imag} */,
  {32'h3cca9eac, 32'h3efdaf28} /* (12, 25, 11) {real, imag} */,
  {32'h3e5cabcc, 32'hbd99cbe8} /* (12, 25, 10) {real, imag} */,
  {32'hbf4096dc, 32'h3f955dd5} /* (12, 25, 9) {real, imag} */,
  {32'hbed57248, 32'h3fd3eb34} /* (12, 25, 8) {real, imag} */,
  {32'h3f3e44fb, 32'hbda32e60} /* (12, 25, 7) {real, imag} */,
  {32'h3f6395de, 32'hbe9b60f4} /* (12, 25, 6) {real, imag} */,
  {32'h3d4b79e0, 32'hbe894af0} /* (12, 25, 5) {real, imag} */,
  {32'h3c89a640, 32'hbe9eb818} /* (12, 25, 4) {real, imag} */,
  {32'hbf5a3933, 32'hbfc000c6} /* (12, 25, 3) {real, imag} */,
  {32'hbfb46da6, 32'hbfb7580f} /* (12, 25, 2) {real, imag} */,
  {32'hbfc6832e, 32'h3eb7c2a8} /* (12, 25, 1) {real, imag} */,
  {32'hbf8eac30, 32'h3f38a7b6} /* (12, 25, 0) {real, imag} */,
  {32'h3e8529af, 32'hbf0df180} /* (12, 24, 31) {real, imag} */,
  {32'h3e57e21c, 32'hbe178dd0} /* (12, 24, 30) {real, imag} */,
  {32'h3e96072c, 32'h3ed06ea0} /* (12, 24, 29) {real, imag} */,
  {32'h3f6e1f51, 32'h3d9bbd60} /* (12, 24, 28) {real, imag} */,
  {32'h3f686687, 32'h3db213d0} /* (12, 24, 27) {real, imag} */,
  {32'h3f3eb7ee, 32'h3e6a3260} /* (12, 24, 26) {real, imag} */,
  {32'h3efa89b8, 32'h3fecac96} /* (12, 24, 25) {real, imag} */,
  {32'hbf1f000c, 32'h3fa17840} /* (12, 24, 24) {real, imag} */,
  {32'hbfb090c6, 32'h3f499120} /* (12, 24, 23) {real, imag} */,
  {32'hbf382329, 32'h3f3f8e10} /* (12, 24, 22) {real, imag} */,
  {32'hbebb4af5, 32'h3d3aac00} /* (12, 24, 21) {real, imag} */,
  {32'hbfc3ef16, 32'h3f110b18} /* (12, 24, 20) {real, imag} */,
  {32'hbfb8e2bc, 32'h3f9cce8f} /* (12, 24, 19) {real, imag} */,
  {32'hbf9e6281, 32'h3b77e800} /* (12, 24, 18) {real, imag} */,
  {32'hbeb70cb4, 32'hbc4edd00} /* (12, 24, 17) {real, imag} */,
  {32'h3f8fe5be, 32'h3e0d8ec0} /* (12, 24, 16) {real, imag} */,
  {32'h3ea83a93, 32'hbf11ad6c} /* (12, 24, 15) {real, imag} */,
  {32'h3cf6b5c0, 32'hbf9a6406} /* (12, 24, 14) {real, imag} */,
  {32'hbea83890, 32'hbf969066} /* (12, 24, 13) {real, imag} */,
  {32'h3f49c5da, 32'hbf224c98} /* (12, 24, 12) {real, imag} */,
  {32'h40107bce, 32'h3d6cf710} /* (12, 24, 11) {real, imag} */,
  {32'h3fdb79fe, 32'h3ea3b01c} /* (12, 24, 10) {real, imag} */,
  {32'h3e37bec0, 32'h3f6084e0} /* (12, 24, 9) {real, imag} */,
  {32'h3d972520, 32'h3fba9d29} /* (12, 24, 8) {real, imag} */,
  {32'h3f6471ae, 32'h3e81df14} /* (12, 24, 7) {real, imag} */,
  {32'h3faf8e0a, 32'h3de6ac30} /* (12, 24, 6) {real, imag} */,
  {32'hbf236253, 32'hbf8f6c48} /* (12, 24, 5) {real, imag} */,
  {32'h3e0e7484, 32'hbfde2711} /* (12, 24, 4) {real, imag} */,
  {32'h3d0ec140, 32'hbfce16a0} /* (12, 24, 3) {real, imag} */,
  {32'hbf56db44, 32'hbf85eac4} /* (12, 24, 2) {real, imag} */,
  {32'h3da28898, 32'hbea19b00} /* (12, 24, 1) {real, imag} */,
  {32'h3da0bab4, 32'h3ea26c58} /* (12, 24, 0) {real, imag} */,
  {32'h3f11ad72, 32'hbf673700} /* (12, 23, 31) {real, imag} */,
  {32'hbe84cc84, 32'hbe45fa80} /* (12, 23, 30) {real, imag} */,
  {32'hbebff398, 32'h3eaaf910} /* (12, 23, 29) {real, imag} */,
  {32'h3f25d0f9, 32'h3ee24ec8} /* (12, 23, 28) {real, imag} */,
  {32'hbd8282b0, 32'h3f2112dc} /* (12, 23, 27) {real, imag} */,
  {32'hbeb5ac48, 32'h3f9a0946} /* (12, 23, 26) {real, imag} */,
  {32'h3f7f53ba, 32'h3fc7a21e} /* (12, 23, 25) {real, imag} */,
  {32'hbeb56e9d, 32'h3e3b11f0} /* (12, 23, 24) {real, imag} */,
  {32'hc011b652, 32'hbee85600} /* (12, 23, 23) {real, imag} */,
  {32'hbffdfe72, 32'hbd2f1580} /* (12, 23, 22) {real, imag} */,
  {32'hbf6d9608, 32'hbe158588} /* (12, 23, 21) {real, imag} */,
  {32'hbfd753fe, 32'hbe9091c4} /* (12, 23, 20) {real, imag} */,
  {32'hbfed72d0, 32'h3d3bd7e0} /* (12, 23, 19) {real, imag} */,
  {32'hbfa06754, 32'hbd9a37d0} /* (12, 23, 18) {real, imag} */,
  {32'hbfa98db2, 32'h3fb1dc59} /* (12, 23, 17) {real, imag} */,
  {32'h3ea2dc0e, 32'h3f99b920} /* (12, 23, 16) {real, imag} */,
  {32'h3d9851d0, 32'h3eeeae80} /* (12, 23, 15) {real, imag} */,
  {32'hbdcf0730, 32'hbe50ebe0} /* (12, 23, 14) {real, imag} */,
  {32'hbe7cde98, 32'hbf8390c4} /* (12, 23, 13) {real, imag} */,
  {32'h3f227e25, 32'hbfc62b5b} /* (12, 23, 12) {real, imag} */,
  {32'h3f9501c2, 32'hbf9a1c19} /* (12, 23, 11) {real, imag} */,
  {32'h3f93d5e2, 32'hbf518d93} /* (12, 23, 10) {real, imag} */,
  {32'h3f6d33ae, 32'hbe857eb0} /* (12, 23, 9) {real, imag} */,
  {32'h3f856dea, 32'h3ea272a0} /* (12, 23, 8) {real, imag} */,
  {32'h3f5a81ff, 32'h3f9f7f6c} /* (12, 23, 7) {real, imag} */,
  {32'h3f1004da, 32'h3fb94d47} /* (12, 23, 6) {real, imag} */,
  {32'hbf52d75b, 32'h3edfbc70} /* (12, 23, 5) {real, imag} */,
  {32'h3eb5c8ec, 32'hbf1f937c} /* (12, 23, 4) {real, imag} */,
  {32'h3ef74b3c, 32'h3bc24b00} /* (12, 23, 3) {real, imag} */,
  {32'hbf2acfcc, 32'h3d1ca240} /* (12, 23, 2) {real, imag} */,
  {32'h3df40920, 32'hbf58c9c4} /* (12, 23, 1) {real, imag} */,
  {32'h3f13a59a, 32'hbfa6feda} /* (12, 23, 0) {real, imag} */,
  {32'hbc960740, 32'h3e2e5e10} /* (12, 22, 31) {real, imag} */,
  {32'hbf9ad9c8, 32'h3eac7450} /* (12, 22, 30) {real, imag} */,
  {32'hbf9f02f6, 32'hbedb0638} /* (12, 22, 29) {real, imag} */,
  {32'hbf3a463a, 32'h3ea42518} /* (12, 22, 28) {real, imag} */,
  {32'hbf9b6696, 32'h3ef19170} /* (12, 22, 27) {real, imag} */,
  {32'hbf31320a, 32'h3f816cb4} /* (12, 22, 26) {real, imag} */,
  {32'h3ebdd398, 32'h3f63bce8} /* (12, 22, 25) {real, imag} */,
  {32'hbe567d23, 32'hbeb61050} /* (12, 22, 24) {real, imag} */,
  {32'hbff6db2f, 32'hbf4ea100} /* (12, 22, 23) {real, imag} */,
  {32'hbff6481e, 32'hbeced280} /* (12, 22, 22) {real, imag} */,
  {32'hbedbd6f8, 32'hbf2aa010} /* (12, 22, 21) {real, imag} */,
  {32'hbf41440e, 32'hbf338706} /* (12, 22, 20) {real, imag} */,
  {32'hbf604d58, 32'h3e65d4dc} /* (12, 22, 19) {real, imag} */,
  {32'hbf87ab9c, 32'h3fd2d622} /* (12, 22, 18) {real, imag} */,
  {32'hbf3fb003, 32'h3fad27e0} /* (12, 22, 17) {real, imag} */,
  {32'h3f39c7e6, 32'h3f90a1f6} /* (12, 22, 16) {real, imag} */,
  {32'hbdd2aab0, 32'h3f8ba12a} /* (12, 22, 15) {real, imag} */,
  {32'hbecbb15c, 32'hbe24b130} /* (12, 22, 14) {real, imag} */,
  {32'h3ed996d0, 32'hbf90334c} /* (12, 22, 13) {real, imag} */,
  {32'h3e95eb34, 32'hbf4f97c0} /* (12, 22, 12) {real, imag} */,
  {32'hbd9196b0, 32'hbf89b9f4} /* (12, 22, 11) {real, imag} */,
  {32'h3f0f7f22, 32'hbf547327} /* (12, 22, 10) {real, imag} */,
  {32'h3db2d1b8, 32'h3dc5dca0} /* (12, 22, 9) {real, imag} */,
  {32'hbed7168c, 32'hbecce910} /* (12, 22, 8) {real, imag} */,
  {32'h3e4b90c0, 32'h3f8330f4} /* (12, 22, 7) {real, imag} */,
  {32'h3ea126ac, 32'h3f3edeac} /* (12, 22, 6) {real, imag} */,
  {32'h3dd729a4, 32'h3eca58c8} /* (12, 22, 5) {real, imag} */,
  {32'hbf15ca1c, 32'hbdf291c0} /* (12, 22, 4) {real, imag} */,
  {32'hbf00c2bc, 32'hba333400} /* (12, 22, 3) {real, imag} */,
  {32'hbfba8a16, 32'h3f668c9c} /* (12, 22, 2) {real, imag} */,
  {32'hbebd9261, 32'hbf2014b2} /* (12, 22, 1) {real, imag} */,
  {32'h3e8085e4, 32'hbf879822} /* (12, 22, 0) {real, imag} */,
  {32'h3efa261e, 32'h3e1b2528} /* (12, 21, 31) {real, imag} */,
  {32'h3e512e18, 32'h3f4896f6} /* (12, 21, 30) {real, imag} */,
  {32'h3eab043c, 32'hbebbe212} /* (12, 21, 29) {real, imag} */,
  {32'hbe8b675c, 32'hbf023dfc} /* (12, 21, 28) {real, imag} */,
  {32'hbf331a7f, 32'hbef08e70} /* (12, 21, 27) {real, imag} */,
  {32'hbf5c74a4, 32'hbea0cd14} /* (12, 21, 26) {real, imag} */,
  {32'hbf8fe2e0, 32'hbf4bd2c9} /* (12, 21, 25) {real, imag} */,
  {32'hbe971bf0, 32'hbd22fcc0} /* (12, 21, 24) {real, imag} */,
  {32'hbf26f337, 32'h3f396f5a} /* (12, 21, 23) {real, imag} */,
  {32'hbf0127c0, 32'h3e1f5fe8} /* (12, 21, 22) {real, imag} */,
  {32'hbf30ef62, 32'hbec70b70} /* (12, 21, 21) {real, imag} */,
  {32'hbdf003b2, 32'hbc96dd10} /* (12, 21, 20) {real, imag} */,
  {32'hbe0b02ec, 32'h3f0b0738} /* (12, 21, 19) {real, imag} */,
  {32'hbf4c6b80, 32'h3fa3ee51} /* (12, 21, 18) {real, imag} */,
  {32'hbf186cae, 32'hbcd52480} /* (12, 21, 17) {real, imag} */,
  {32'h3e99019e, 32'h3f0380cc} /* (12, 21, 16) {real, imag} */,
  {32'hbf02049c, 32'h3ddcbd60} /* (12, 21, 15) {real, imag} */,
  {32'hbf89c946, 32'hbf3dbbea} /* (12, 21, 14) {real, imag} */,
  {32'hbdbf99b8, 32'hbf54dce7} /* (12, 21, 13) {real, imag} */,
  {32'h3ea8e692, 32'hbf82642c} /* (12, 21, 12) {real, imag} */,
  {32'hbe8353c5, 32'hbf2d6ce0} /* (12, 21, 11) {real, imag} */,
  {32'hbdef36c8, 32'h3ebcd224} /* (12, 21, 10) {real, imag} */,
  {32'h3f4bcf4c, 32'h3fa4efce} /* (12, 21, 9) {real, imag} */,
  {32'h3eec3056, 32'h3e2ccb60} /* (12, 21, 8) {real, imag} */,
  {32'h3f141922, 32'h3ee98b74} /* (12, 21, 7) {real, imag} */,
  {32'hbe0819f2, 32'hbf3141df} /* (12, 21, 6) {real, imag} */,
  {32'h3c1a6dc0, 32'hbf250e89} /* (12, 21, 5) {real, imag} */,
  {32'hbea10166, 32'hbf2d0c97} /* (12, 21, 4) {real, imag} */,
  {32'hbe8b1c4a, 32'hbf747fed} /* (12, 21, 3) {real, imag} */,
  {32'hbf2b0b50, 32'hbf2d9f5b} /* (12, 21, 2) {real, imag} */,
  {32'h3e8606f6, 32'hbfaf05b8} /* (12, 21, 1) {real, imag} */,
  {32'h3f1c8ea8, 32'hbf2f7f42} /* (12, 21, 0) {real, imag} */,
  {32'hbe8bb0fb, 32'hbeb692be} /* (12, 20, 31) {real, imag} */,
  {32'hbed1cada, 32'h3db0ebac} /* (12, 20, 30) {real, imag} */,
  {32'hbd727a10, 32'hbe54c470} /* (12, 20, 29) {real, imag} */,
  {32'hbf49f623, 32'hbdee1ae0} /* (12, 20, 28) {real, imag} */,
  {32'hbf03d9b8, 32'hbf91f829} /* (12, 20, 27) {real, imag} */,
  {32'hbe412730, 32'hbf1f9a9c} /* (12, 20, 26) {real, imag} */,
  {32'hbe0f0b48, 32'h3d4eb780} /* (12, 20, 25) {real, imag} */,
  {32'h3fa340b4, 32'h3eae7cb0} /* (12, 20, 24) {real, imag} */,
  {32'h3fa64d42, 32'hbe05afb0} /* (12, 20, 23) {real, imag} */,
  {32'h3f01ed26, 32'hbea990e0} /* (12, 20, 22) {real, imag} */,
  {32'hbf5a8329, 32'hbe854730} /* (12, 20, 21) {real, imag} */,
  {32'hbf991c67, 32'h3dc72cd0} /* (12, 20, 20) {real, imag} */,
  {32'hbe7d3c00, 32'h3f5e0da4} /* (12, 20, 19) {real, imag} */,
  {32'h3f460d4c, 32'h3e84faf4} /* (12, 20, 18) {real, imag} */,
  {32'h3f12a719, 32'hbfd3dbf8} /* (12, 20, 17) {real, imag} */,
  {32'h3f8bb36a, 32'hbf2b6fdf} /* (12, 20, 16) {real, imag} */,
  {32'h3e822b74, 32'h3e13a6c0} /* (12, 20, 15) {real, imag} */,
  {32'hbf02b46a, 32'hbea08688} /* (12, 20, 14) {real, imag} */,
  {32'hbf829ced, 32'hbe99df48} /* (12, 20, 13) {real, imag} */,
  {32'hbf956996, 32'h3d960420} /* (12, 20, 12) {real, imag} */,
  {32'hbf950749, 32'hbefb7a58} /* (12, 20, 11) {real, imag} */,
  {32'hbf2b0ff3, 32'h3e12d7e9} /* (12, 20, 10) {real, imag} */,
  {32'h3f624818, 32'h3fae6023} /* (12, 20, 9) {real, imag} */,
  {32'h3f306b92, 32'h3fa58ad6} /* (12, 20, 8) {real, imag} */,
  {32'h3ec2de59, 32'h3f2d32c0} /* (12, 20, 7) {real, imag} */,
  {32'hbe33c83c, 32'hbf656298} /* (12, 20, 6) {real, imag} */,
  {32'h3ebca397, 32'hbfa8661c} /* (12, 20, 5) {real, imag} */,
  {32'h3f138bf8, 32'hbe92398c} /* (12, 20, 4) {real, imag} */,
  {32'h3ed6b075, 32'hbf07ce0c} /* (12, 20, 3) {real, imag} */,
  {32'h3e8f5c48, 32'hbf2d0090} /* (12, 20, 2) {real, imag} */,
  {32'h3f11dee1, 32'hbf41f364} /* (12, 20, 1) {real, imag} */,
  {32'h3f0486a7, 32'hbf39541e} /* (12, 20, 0) {real, imag} */,
  {32'hbef1887c, 32'hbd67cee0} /* (12, 19, 31) {real, imag} */,
  {32'hbeba53b8, 32'h3f211785} /* (12, 19, 30) {real, imag} */,
  {32'hbf8f1a84, 32'hbda7edf0} /* (12, 19, 29) {real, imag} */,
  {32'hbedf965e, 32'hbe8fe3e0} /* (12, 19, 28) {real, imag} */,
  {32'h3e80630b, 32'hbf7a8acc} /* (12, 19, 27) {real, imag} */,
  {32'h3f895b0e, 32'h3e1c83d0} /* (12, 19, 26) {real, imag} */,
  {32'h3f17d8d9, 32'h3e86cf78} /* (12, 19, 25) {real, imag} */,
  {32'h3f54a47c, 32'h3fa3f842} /* (12, 19, 24) {real, imag} */,
  {32'h3f064908, 32'hbe3d9fa0} /* (12, 19, 23) {real, imag} */,
  {32'h3edbf1b8, 32'hbf226e38} /* (12, 19, 22) {real, imag} */,
  {32'h3ebdcf14, 32'hbed43168} /* (12, 19, 21) {real, imag} */,
  {32'hbe9c6a49, 32'hbf2a7528} /* (12, 19, 20) {real, imag} */,
  {32'hbe6cbc44, 32'h3e013a70} /* (12, 19, 19) {real, imag} */,
  {32'h3dd9a958, 32'hbeef6190} /* (12, 19, 18) {real, imag} */,
  {32'h3f0e5b8a, 32'hbf757c68} /* (12, 19, 17) {real, imag} */,
  {32'hbe7b4f80, 32'h3ef9c30b} /* (12, 19, 16) {real, imag} */,
  {32'hbf102058, 32'h3ef8d2b0} /* (12, 19, 15) {real, imag} */,
  {32'hbef18b34, 32'h3e293f30} /* (12, 19, 14) {real, imag} */,
  {32'hbf293914, 32'hbc47f600} /* (12, 19, 13) {real, imag} */,
  {32'hbf86cdac, 32'h3f8c8d36} /* (12, 19, 12) {real, imag} */,
  {32'hbed79bc6, 32'h3ef678b0} /* (12, 19, 11) {real, imag} */,
  {32'h3fa17b04, 32'hbd581e20} /* (12, 19, 10) {real, imag} */,
  {32'h3f936ec0, 32'h3e624730} /* (12, 19, 9) {real, imag} */,
  {32'h3ea4a4c9, 32'h3e4ba960} /* (12, 19, 8) {real, imag} */,
  {32'hbc5f4980, 32'h3ec0d5d0} /* (12, 19, 7) {real, imag} */,
  {32'h3efe8bb0, 32'h3f1dcc86} /* (12, 19, 6) {real, imag} */,
  {32'h3f67f2ac, 32'hbeae6d80} /* (12, 19, 5) {real, imag} */,
  {32'h3eb8c1fc, 32'hbf95f2f5} /* (12, 19, 4) {real, imag} */,
  {32'hbf3f1de2, 32'hbf745158} /* (12, 19, 3) {real, imag} */,
  {32'h3e025fa0, 32'hbdff1160} /* (12, 19, 2) {real, imag} */,
  {32'h3f92611c, 32'hbf07cee0} /* (12, 19, 1) {real, imag} */,
  {32'h3ea7114c, 32'hbfce2c5c} /* (12, 19, 0) {real, imag} */,
  {32'h3df72a28, 32'h3f11d844} /* (12, 18, 31) {real, imag} */,
  {32'hbe8290b4, 32'h3f2500d2} /* (12, 18, 30) {real, imag} */,
  {32'hbea96ef4, 32'h3f8a8c64} /* (12, 18, 29) {real, imag} */,
  {32'h3e006368, 32'h3e184d64} /* (12, 18, 28) {real, imag} */,
  {32'hbe523bf8, 32'hbf051960} /* (12, 18, 27) {real, imag} */,
  {32'h3f7453bc, 32'hbe462180} /* (12, 18, 26) {real, imag} */,
  {32'h3fa5e158, 32'hbdcaeac0} /* (12, 18, 25) {real, imag} */,
  {32'h3f104568, 32'hbe9c4658} /* (12, 18, 24) {real, imag} */,
  {32'hbf38847a, 32'hbf32ddac} /* (12, 18, 23) {real, imag} */,
  {32'hbcc0de80, 32'hbf6d5214} /* (12, 18, 22) {real, imag} */,
  {32'h3f9dd9c5, 32'hbf37a7a7} /* (12, 18, 21) {real, imag} */,
  {32'h3e3c6824, 32'hbf79573c} /* (12, 18, 20) {real, imag} */,
  {32'h3ef207c6, 32'hbf982712} /* (12, 18, 19) {real, imag} */,
  {32'hbfd34804, 32'hbf07ba60} /* (12, 18, 18) {real, imag} */,
  {32'hc0051faa, 32'hbb79e400} /* (12, 18, 17) {real, imag} */,
  {32'hbf569918, 32'h3e97ba4c} /* (12, 18, 16) {real, imag} */,
  {32'hbef508ca, 32'h3f5f60be} /* (12, 18, 15) {real, imag} */,
  {32'hbf4281bc, 32'h3f050c7a} /* (12, 18, 14) {real, imag} */,
  {32'hbf9793e1, 32'hbf2c558c} /* (12, 18, 13) {real, imag} */,
  {32'hbfbea8d2, 32'h3e93d6c8} /* (12, 18, 12) {real, imag} */,
  {32'hbf603970, 32'h3f7a2ba2} /* (12, 18, 11) {real, imag} */,
  {32'h3e810032, 32'hbe668b98} /* (12, 18, 10) {real, imag} */,
  {32'h3f4a9ed9, 32'hbfb018a4} /* (12, 18, 9) {real, imag} */,
  {32'h3d9e08e5, 32'hbfb99e52} /* (12, 18, 8) {real, imag} */,
  {32'hbe3a3184, 32'hbf47943c} /* (12, 18, 7) {real, imag} */,
  {32'hbee47fe4, 32'h3df2aff0} /* (12, 18, 6) {real, imag} */,
  {32'hbea89d88, 32'h3ec05190} /* (12, 18, 5) {real, imag} */,
  {32'hbeeb0f38, 32'hbf24b908} /* (12, 18, 4) {real, imag} */,
  {32'hbf6ab60d, 32'hbfa60ae9} /* (12, 18, 3) {real, imag} */,
  {32'hbf30fea0, 32'hbfa8dc20} /* (12, 18, 2) {real, imag} */,
  {32'h3eb13c78, 32'hbd481900} /* (12, 18, 1) {real, imag} */,
  {32'h3e0f5de8, 32'hbf8d071b} /* (12, 18, 0) {real, imag} */,
  {32'h3b9cdc00, 32'h3e471030} /* (12, 17, 31) {real, imag} */,
  {32'hbf2346d6, 32'h3daa8c20} /* (12, 17, 30) {real, imag} */,
  {32'hbef254c4, 32'h3ec6e9f0} /* (12, 17, 29) {real, imag} */,
  {32'h3e723cc0, 32'hbdc64940} /* (12, 17, 28) {real, imag} */,
  {32'h3f31c8f8, 32'hbf4fc030} /* (12, 17, 27) {real, imag} */,
  {32'h3f6f3eda, 32'hbf94f400} /* (12, 17, 26) {real, imag} */,
  {32'h3fbd26e0, 32'hbf720d1e} /* (12, 17, 25) {real, imag} */,
  {32'h3ed57774, 32'hbf65bdec} /* (12, 17, 24) {real, imag} */,
  {32'hbfa404e0, 32'hbf221740} /* (12, 17, 23) {real, imag} */,
  {32'hbe82b2e8, 32'hbfc10f20} /* (12, 17, 22) {real, imag} */,
  {32'h3f379850, 32'hbf512982} /* (12, 17, 21) {real, imag} */,
  {32'hbf4c547d, 32'hbfc14193} /* (12, 17, 20) {real, imag} */,
  {32'hbdfbd480, 32'hbf884a9a} /* (12, 17, 19) {real, imag} */,
  {32'hbfa17c9e, 32'hbe445ab0} /* (12, 17, 18) {real, imag} */,
  {32'hbfb24340, 32'hbf1bb950} /* (12, 17, 17) {real, imag} */,
  {32'h3dcafe14, 32'h3ece4fe8} /* (12, 17, 16) {real, imag} */,
  {32'hbef83fe3, 32'h3f7a144e} /* (12, 17, 15) {real, imag} */,
  {32'hbf5a4d4c, 32'hbc79f100} /* (12, 17, 14) {real, imag} */,
  {32'hbf45ee72, 32'hbf8b9297} /* (12, 17, 13) {real, imag} */,
  {32'hbf7f467a, 32'hbbf50400} /* (12, 17, 12) {real, imag} */,
  {32'hbe985521, 32'h3ea73abc} /* (12, 17, 11) {real, imag} */,
  {32'h3e8159c7, 32'hbf1d0e88} /* (12, 17, 10) {real, imag} */,
  {32'hbd5db060, 32'hbfaadfdc} /* (12, 17, 9) {real, imag} */,
  {32'hbf88fc75, 32'hc00cbbd0} /* (12, 17, 8) {real, imag} */,
  {32'hbf838e10, 32'hbf82bb00} /* (12, 17, 7) {real, imag} */,
  {32'hbfccd122, 32'h3dc4adc0} /* (12, 17, 6) {real, imag} */,
  {32'hbfa58280, 32'h3f422bbc} /* (12, 17, 5) {real, imag} */,
  {32'hbf2d6074, 32'h3e10a330} /* (12, 17, 4) {real, imag} */,
  {32'hbf9e539e, 32'h3dc52cd8} /* (12, 17, 3) {real, imag} */,
  {32'hbfb6bfc5, 32'h3d917a08} /* (12, 17, 2) {real, imag} */,
  {32'h3e412fd0, 32'h3eb28a7e} /* (12, 17, 1) {real, imag} */,
  {32'h3f973030, 32'hbe91e9ec} /* (12, 17, 0) {real, imag} */,
  {32'h3b72a700, 32'h3de2cbd0} /* (12, 16, 31) {real, imag} */,
  {32'hbd7acbd0, 32'h3ee8a518} /* (12, 16, 30) {real, imag} */,
  {32'hbf29b98e, 32'h3f19fb8c} /* (12, 16, 29) {real, imag} */,
  {32'h3e40d340, 32'hbe339720} /* (12, 16, 28) {real, imag} */,
  {32'h3e969eb8, 32'hbf2aa064} /* (12, 16, 27) {real, imag} */,
  {32'h3f2ffa62, 32'hbecdb980} /* (12, 16, 26) {real, imag} */,
  {32'h3f86781f, 32'hbf89ab3a} /* (12, 16, 25) {real, imag} */,
  {32'h3f6faff7, 32'h3f1d9814} /* (12, 16, 24) {real, imag} */,
  {32'hbde455e0, 32'h3f64870a} /* (12, 16, 23) {real, imag} */,
  {32'h3ea16f94, 32'hbf1d9b78} /* (12, 16, 22) {real, imag} */,
  {32'hbe08ead8, 32'hbe6f7d90} /* (12, 16, 21) {real, imag} */,
  {32'hbf8b7786, 32'hbf6c1f68} /* (12, 16, 20) {real, imag} */,
  {32'hbf1e6a18, 32'hbe0494e0} /* (12, 16, 19) {real, imag} */,
  {32'hbf0e135c, 32'h3f6a3b6e} /* (12, 16, 18) {real, imag} */,
  {32'hbe9d34f0, 32'h3eb74af8} /* (12, 16, 17) {real, imag} */,
  {32'hbda04780, 32'h3ce7aa00} /* (12, 16, 16) {real, imag} */,
  {32'h3d6b3650, 32'hbf09b9fc} /* (12, 16, 15) {real, imag} */,
  {32'hbf3c9cea, 32'hbee63528} /* (12, 16, 14) {real, imag} */,
  {32'hbeb55364, 32'h3f148834} /* (12, 16, 13) {real, imag} */,
  {32'hbe4ca970, 32'h3f5c9392} /* (12, 16, 12) {real, imag} */,
  {32'h3ee61858, 32'h3f99bc93} /* (12, 16, 11) {real, imag} */,
  {32'h3f0817b9, 32'h3f88e7fb} /* (12, 16, 10) {real, imag} */,
  {32'hbe50dc88, 32'hbf08ba7c} /* (12, 16, 9) {real, imag} */,
  {32'hbf66199c, 32'hbf01db6c} /* (12, 16, 8) {real, imag} */,
  {32'hbe8cfa9c, 32'hbdf91740} /* (12, 16, 7) {real, imag} */,
  {32'hbeca3508, 32'hbf35c988} /* (12, 16, 6) {real, imag} */,
  {32'hbe9174b0, 32'h3f8b494b} /* (12, 16, 5) {real, imag} */,
  {32'hbf4feb2a, 32'h3fa82cb2} /* (12, 16, 4) {real, imag} */,
  {32'hbfe3a294, 32'h3fc448ee} /* (12, 16, 3) {real, imag} */,
  {32'hbfa69adf, 32'h3fad1e29} /* (12, 16, 2) {real, imag} */,
  {32'h3d37a290, 32'h3f3ec1ec} /* (12, 16, 1) {real, imag} */,
  {32'h3e10e0d4, 32'h3e9ede30} /* (12, 16, 0) {real, imag} */,
  {32'hbeedb1ac, 32'hbe2853bc} /* (12, 15, 31) {real, imag} */,
  {32'hbf9accbb, 32'h3d1af540} /* (12, 15, 30) {real, imag} */,
  {32'hc0004f74, 32'hbe8247a0} /* (12, 15, 29) {real, imag} */,
  {32'hbd0ae780, 32'h3d7764c0} /* (12, 15, 28) {real, imag} */,
  {32'h3f34168d, 32'h3e35a460} /* (12, 15, 27) {real, imag} */,
  {32'h3f71ed4c, 32'hbd2b6ae0} /* (12, 15, 26) {real, imag} */,
  {32'h3fb6c48e, 32'hbf10fbee} /* (12, 15, 25) {real, imag} */,
  {32'h3f61fb46, 32'h3ef3a3d0} /* (12, 15, 24) {real, imag} */,
  {32'h3f2c2285, 32'h3f58e1e0} /* (12, 15, 23) {real, imag} */,
  {32'h3e64a349, 32'h3c95db80} /* (12, 15, 22) {real, imag} */,
  {32'hbf0176bd, 32'h3acb6000} /* (12, 15, 21) {real, imag} */,
  {32'h3e0241ec, 32'hbd1d41c0} /* (12, 15, 20) {real, imag} */,
  {32'hbdea9550, 32'h3e9ab3f0} /* (12, 15, 19) {real, imag} */,
  {32'hbdedd39c, 32'h3ef07920} /* (12, 15, 18) {real, imag} */,
  {32'h3ed5aee8, 32'h3d0d1280} /* (12, 15, 17) {real, imag} */,
  {32'hbcc42080, 32'hbe826a98} /* (12, 15, 16) {real, imag} */,
  {32'hbeb8feda, 32'hbf736b60} /* (12, 15, 15) {real, imag} */,
  {32'hbf0f512a, 32'hbf4c828c} /* (12, 15, 14) {real, imag} */,
  {32'hbe85cc4e, 32'h3dc36c60} /* (12, 15, 13) {real, imag} */,
  {32'hbd145fc0, 32'h3f8a483f} /* (12, 15, 12) {real, imag} */,
  {32'h3ec762a5, 32'h3f6e01be} /* (12, 15, 11) {real, imag} */,
  {32'hbdf79000, 32'hba1ff800} /* (12, 15, 10) {real, imag} */,
  {32'hbefdc188, 32'hbf8a4d6d} /* (12, 15, 9) {real, imag} */,
  {32'hbf7e4414, 32'hbe9fa768} /* (12, 15, 8) {real, imag} */,
  {32'hbf61e6ac, 32'h3da08c40} /* (12, 15, 7) {real, imag} */,
  {32'h3df133b0, 32'hbe7b43d0} /* (12, 15, 6) {real, imag} */,
  {32'h3ed16d0c, 32'h3db95e80} /* (12, 15, 5) {real, imag} */,
  {32'hbea9e310, 32'h3d31d300} /* (12, 15, 4) {real, imag} */,
  {32'hbf6f637c, 32'h3f19d63c} /* (12, 15, 3) {real, imag} */,
  {32'hbeee966c, 32'h3ecd5408} /* (12, 15, 2) {real, imag} */,
  {32'h3f06fce2, 32'h3eb3f520} /* (12, 15, 1) {real, imag} */,
  {32'hbd9aa9f8, 32'h3df6a530} /* (12, 15, 0) {real, imag} */,
  {32'hbf05521f, 32'h3f1c0f5a} /* (12, 14, 31) {real, imag} */,
  {32'hbf84bc28, 32'h3f56a0a0} /* (12, 14, 30) {real, imag} */,
  {32'hbf83e0ae, 32'hbec1bf08} /* (12, 14, 29) {real, imag} */,
  {32'hbe2a8140, 32'hbee1ad50} /* (12, 14, 28) {real, imag} */,
  {32'h3f47a44f, 32'h3e814450} /* (12, 14, 27) {real, imag} */,
  {32'h3f896c2c, 32'hbe845f0c} /* (12, 14, 26) {real, imag} */,
  {32'h3f8ee150, 32'hbf988e36} /* (12, 14, 25) {real, imag} */,
  {32'h3f0057d8, 32'hbeabbfc4} /* (12, 14, 24) {real, imag} */,
  {32'h3f0b8aa2, 32'h3ebafe60} /* (12, 14, 23) {real, imag} */,
  {32'h3cc75750, 32'h3d1a10c0} /* (12, 14, 22) {real, imag} */,
  {32'hbedf2550, 32'h3e3c8f80} /* (12, 14, 21) {real, imag} */,
  {32'hbf895496, 32'hbe6617c8} /* (12, 14, 20) {real, imag} */,
  {32'hbf15cf8c, 32'h3f9e7ef2} /* (12, 14, 19) {real, imag} */,
  {32'hbeca3f1c, 32'h3f6d91d0} /* (12, 14, 18) {real, imag} */,
  {32'hbee0ad17, 32'h3da7d4a0} /* (12, 14, 17) {real, imag} */,
  {32'hbf32406e, 32'h3ea54b70} /* (12, 14, 16) {real, imag} */,
  {32'hbf1b4a7a, 32'hbc3cff00} /* (12, 14, 15) {real, imag} */,
  {32'h3e81573c, 32'hbfa6f88c} /* (12, 14, 14) {real, imag} */,
  {32'hbe479368, 32'hbf9bb455} /* (12, 14, 13) {real, imag} */,
  {32'h3ee30caa, 32'hbe2b5084} /* (12, 14, 12) {real, imag} */,
  {32'hbeb63430, 32'hbe294b1c} /* (12, 14, 11) {real, imag} */,
  {32'hbfa56863, 32'h3eb876d0} /* (12, 14, 10) {real, imag} */,
  {32'hbf880dc2, 32'h3c19f100} /* (12, 14, 9) {real, imag} */,
  {32'hbf3aa0b3, 32'h3daa0880} /* (12, 14, 8) {real, imag} */,
  {32'hbf77fcfd, 32'h3ed8f0f8} /* (12, 14, 7) {real, imag} */,
  {32'hbd535430, 32'h3cb51f00} /* (12, 14, 6) {real, imag} */,
  {32'h3f37a934, 32'hbef78040} /* (12, 14, 5) {real, imag} */,
  {32'h3e5182b0, 32'hbec81028} /* (12, 14, 4) {real, imag} */,
  {32'hbe091f30, 32'h3e4822c0} /* (12, 14, 3) {real, imag} */,
  {32'h39faf000, 32'h3e0d6170} /* (12, 14, 2) {real, imag} */,
  {32'h3e64a51c, 32'hbf028a10} /* (12, 14, 1) {real, imag} */,
  {32'hbe8eea86, 32'hbf678df6} /* (12, 14, 0) {real, imag} */,
  {32'hbdc34b10, 32'h3f2f2e32} /* (12, 13, 31) {real, imag} */,
  {32'h3ee281cc, 32'h3f3550a0} /* (12, 13, 30) {real, imag} */,
  {32'h3f3b5f00, 32'hbe0a8af0} /* (12, 13, 29) {real, imag} */,
  {32'h3ea57768, 32'h3ecd93c0} /* (12, 13, 28) {real, imag} */,
  {32'hbe5e93f0, 32'h3f857950} /* (12, 13, 27) {real, imag} */,
  {32'h3ef63cec, 32'hbec71fe8} /* (12, 13, 26) {real, imag} */,
  {32'h3f171bf6, 32'hbfb6ec7e} /* (12, 13, 25) {real, imag} */,
  {32'h3edf9470, 32'hbe865290} /* (12, 13, 24) {real, imag} */,
  {32'h3ee69c8c, 32'h3f1b3e44} /* (12, 13, 23) {real, imag} */,
  {32'hbef21a76, 32'hbc459100} /* (12, 13, 22) {real, imag} */,
  {32'hbfc8f42e, 32'hbe210bf0} /* (12, 13, 21) {real, imag} */,
  {32'hc0089c75, 32'hbf7bca12} /* (12, 13, 20) {real, imag} */,
  {32'hbf447382, 32'h3f91b82a} /* (12, 13, 19) {real, imag} */,
  {32'hbf9c73f7, 32'h3f0dc0f0} /* (12, 13, 18) {real, imag} */,
  {32'h3e3696a8, 32'hbec0bdf0} /* (12, 13, 17) {real, imag} */,
  {32'h3f4c098e, 32'h3eb453b0} /* (12, 13, 16) {real, imag} */,
  {32'hbe7105bc, 32'hbe2bb930} /* (12, 13, 15) {real, imag} */,
  {32'hbf56aa88, 32'hbf982dc4} /* (12, 13, 14) {real, imag} */,
  {32'hbebc59fa, 32'hbfcf6ab4} /* (12, 13, 13) {real, imag} */,
  {32'h3f1a8e88, 32'hbed255a8} /* (12, 13, 12) {real, imag} */,
  {32'hbc294a80, 32'h3e9d9dc8} /* (12, 13, 11) {real, imag} */,
  {32'hbf61a911, 32'h3f06f034} /* (12, 13, 10) {real, imag} */,
  {32'hbf32a6cd, 32'h3c0c8700} /* (12, 13, 9) {real, imag} */,
  {32'hbe87e198, 32'hbfa21a0e} /* (12, 13, 8) {real, imag} */,
  {32'hbdefdf20, 32'hbe8da008} /* (12, 13, 7) {real, imag} */,
  {32'hbe903bfc, 32'h3eb46d60} /* (12, 13, 6) {real, imag} */,
  {32'h3e1ddd28, 32'hbeef9f70} /* (12, 13, 5) {real, imag} */,
  {32'hbd9d5d30, 32'h3d4baac0} /* (12, 13, 4) {real, imag} */,
  {32'h3dc20a00, 32'h3e8fc520} /* (12, 13, 3) {real, imag} */,
  {32'h3dfb3680, 32'hbf7813e8} /* (12, 13, 2) {real, imag} */,
  {32'h3f519f9d, 32'hbf8538c8} /* (12, 13, 1) {real, imag} */,
  {32'hbbc241a0, 32'hbf1afbf7} /* (12, 13, 0) {real, imag} */,
  {32'hbd1164e0, 32'h3eb3553c} /* (12, 12, 31) {real, imag} */,
  {32'h3f605f76, 32'h3da5d4a0} /* (12, 12, 30) {real, imag} */,
  {32'h3f163772, 32'hbd238a80} /* (12, 12, 29) {real, imag} */,
  {32'hbe1c0be0, 32'h3e748680} /* (12, 12, 28) {real, imag} */,
  {32'h3ec86c94, 32'h3e6ecc70} /* (12, 12, 27) {real, imag} */,
  {32'h3f18399c, 32'hbeb6aef8} /* (12, 12, 26) {real, imag} */,
  {32'h3f260904, 32'hbf3af234} /* (12, 12, 25) {real, imag} */,
  {32'h3ebb79a0, 32'hbf7265f8} /* (12, 12, 24) {real, imag} */,
  {32'hbe645f90, 32'hbf1d3868} /* (12, 12, 23) {real, imag} */,
  {32'hbf4f8e24, 32'h3e1ad398} /* (12, 12, 22) {real, imag} */,
  {32'hbf17f93a, 32'h3e83d368} /* (12, 12, 21) {real, imag} */,
  {32'hbee15fba, 32'h3f3a4e36} /* (12, 12, 20) {real, imag} */,
  {32'h3de79500, 32'h3fc77e2a} /* (12, 12, 19) {real, imag} */,
  {32'hbf3ea5b8, 32'h3eb0bdb8} /* (12, 12, 18) {real, imag} */,
  {32'hbe883768, 32'hbeacdc78} /* (12, 12, 17) {real, imag} */,
  {32'h3b5a1800, 32'h3f35c12c} /* (12, 12, 16) {real, imag} */,
  {32'h3d6a4720, 32'h3d90f4e0} /* (12, 12, 15) {real, imag} */,
  {32'hbf69d1c8, 32'hbfcbf8b2} /* (12, 12, 14) {real, imag} */,
  {32'hbeb262a0, 32'hbfe6bb03} /* (12, 12, 13) {real, imag} */,
  {32'h3e869fec, 32'hbe830490} /* (12, 12, 12) {real, imag} */,
  {32'h3f3a619a, 32'h3f49d380} /* (12, 12, 11) {real, imag} */,
  {32'h3dc25c85, 32'hbe3e965b} /* (12, 12, 10) {real, imag} */,
  {32'hbee02d84, 32'hbf1a09c4} /* (12, 12, 9) {real, imag} */,
  {32'h3ec75844, 32'hbfb9c3dc} /* (12, 12, 8) {real, imag} */,
  {32'h3ed01c04, 32'hbf808cd4} /* (12, 12, 7) {real, imag} */,
  {32'h3f6bbfb0, 32'hbf0db7fc} /* (12, 12, 6) {real, imag} */,
  {32'h3f262052, 32'hbf5f5258} /* (12, 12, 5) {real, imag} */,
  {32'hbe34fe90, 32'h3f57459e} /* (12, 12, 4) {real, imag} */,
  {32'hbf196366, 32'h3efcdc68} /* (12, 12, 3) {real, imag} */,
  {32'hbf02f7f0, 32'hbec6ddb8} /* (12, 12, 2) {real, imag} */,
  {32'h3f9b9b07, 32'hbf874cf2} /* (12, 12, 1) {real, imag} */,
  {32'h3f16c28b, 32'hbd76e000} /* (12, 12, 0) {real, imag} */,
  {32'h3c29b600, 32'h3ec96b3c} /* (12, 11, 31) {real, imag} */,
  {32'h3f2a8ee8, 32'h3f4bbfa6} /* (12, 11, 30) {real, imag} */,
  {32'hbf11f24b, 32'h3f9ee1b6} /* (12, 11, 29) {real, imag} */,
  {32'hbfda9ab8, 32'h3f579e84} /* (12, 11, 28) {real, imag} */,
  {32'hbf34be19, 32'hbe9d6230} /* (12, 11, 27) {real, imag} */,
  {32'hbef87fac, 32'h3d8a8330} /* (12, 11, 26) {real, imag} */,
  {32'hbe976d8c, 32'h3fba526b} /* (12, 11, 25) {real, imag} */,
  {32'hbf1d68bc, 32'h3f5d6412} /* (12, 11, 24) {real, imag} */,
  {32'hbd2e8c60, 32'hbef6ebb8} /* (12, 11, 23) {real, imag} */,
  {32'h3f76adb9, 32'h3f08c6ec} /* (12, 11, 22) {real, imag} */,
  {32'h3ed2bd98, 32'h3eb70c90} /* (12, 11, 21) {real, imag} */,
  {32'hbf18519a, 32'h3f652bfd} /* (12, 11, 20) {real, imag} */,
  {32'hbf706f18, 32'h3fc23874} /* (12, 11, 19) {real, imag} */,
  {32'h3e0a44c8, 32'h400acbd5} /* (12, 11, 18) {real, imag} */,
  {32'h3e808d18, 32'h3f3c75d4} /* (12, 11, 17) {real, imag} */,
  {32'h3f1761f8, 32'h3dae7700} /* (12, 11, 16) {real, imag} */,
  {32'h3ee600fa, 32'h3e951348} /* (12, 11, 15) {real, imag} */,
  {32'hbf1385fb, 32'hbfb3367a} /* (12, 11, 14) {real, imag} */,
  {32'h3c8a4470, 32'hbf8575e3} /* (12, 11, 13) {real, imag} */,
  {32'h3fa4edd9, 32'h3f3054dc} /* (12, 11, 12) {real, imag} */,
  {32'h3f9136bc, 32'h3f6833e4} /* (12, 11, 11) {real, imag} */,
  {32'h3ef5de44, 32'h3d9a2450} /* (12, 11, 10) {real, imag} */,
  {32'hbe2553d8, 32'h3ea8d210} /* (12, 11, 9) {real, imag} */,
  {32'h3f110a58, 32'hbeaf2e68} /* (12, 11, 8) {real, imag} */,
  {32'h3f5e03d6, 32'hbeefc0a0} /* (12, 11, 7) {real, imag} */,
  {32'h3f909546, 32'hbf1738a0} /* (12, 11, 6) {real, imag} */,
  {32'h3fa4f1e8, 32'hbf44d94c} /* (12, 11, 5) {real, imag} */,
  {32'h3f016566, 32'h3f6141d8} /* (12, 11, 4) {real, imag} */,
  {32'hbfa2a888, 32'hbebcabf8} /* (12, 11, 3) {real, imag} */,
  {32'hbf521714, 32'hbedab7e0} /* (12, 11, 2) {real, imag} */,
  {32'h3e1328ee, 32'hbf154840} /* (12, 11, 1) {real, imag} */,
  {32'h3ec32df2, 32'hbedd9640} /* (12, 11, 0) {real, imag} */,
  {32'hbe9e19f0, 32'h3f4fdf78} /* (12, 10, 31) {real, imag} */,
  {32'h3d3c2a80, 32'h3fd713f0} /* (12, 10, 30) {real, imag} */,
  {32'h3f19f584, 32'h3f778aa0} /* (12, 10, 29) {real, imag} */,
  {32'hbcd69760, 32'h3f016b06} /* (12, 10, 28) {real, imag} */,
  {32'hbe783968, 32'hbe1fbc60} /* (12, 10, 27) {real, imag} */,
  {32'hbec15c48, 32'h3ee3b638} /* (12, 10, 26) {real, imag} */,
  {32'hbf8d98c9, 32'h3f4d6ca2} /* (12, 10, 25) {real, imag} */,
  {32'hc0008426, 32'h3f731afa} /* (12, 10, 24) {real, imag} */,
  {32'hbd24e9eb, 32'hbf314ff8} /* (12, 10, 23) {real, imag} */,
  {32'h3d319170, 32'hbfb34b53} /* (12, 10, 22) {real, imag} */,
  {32'hbe50bf46, 32'hbf7b3b7a} /* (12, 10, 21) {real, imag} */,
  {32'h3e598e48, 32'h3d96dc20} /* (12, 10, 20) {real, imag} */,
  {32'hbb54d500, 32'h3e060513} /* (12, 10, 19) {real, imag} */,
  {32'h3e02c638, 32'h3f96e8f8} /* (12, 10, 18) {real, imag} */,
  {32'h3ee1ac3c, 32'h3f876f5b} /* (12, 10, 17) {real, imag} */,
  {32'h3fd882fd, 32'hbe625170} /* (12, 10, 16) {real, imag} */,
  {32'h40088bb0, 32'hbf2f0404} /* (12, 10, 15) {real, imag} */,
  {32'h3f8682bb, 32'hbe6b2244} /* (12, 10, 14) {real, imag} */,
  {32'h3e20e510, 32'h3f67ddca} /* (12, 10, 13) {real, imag} */,
  {32'h3f145e22, 32'hbd82c780} /* (12, 10, 12) {real, imag} */,
  {32'h3dcc18d8, 32'hbeb926c2} /* (12, 10, 11) {real, imag} */,
  {32'hbeac60df, 32'hbf39536f} /* (12, 10, 10) {real, imag} */,
  {32'hbf08c954, 32'h3d1a934e} /* (12, 10, 9) {real, imag} */,
  {32'h3e4633ca, 32'hbed11ab8} /* (12, 10, 8) {real, imag} */,
  {32'h3f67f430, 32'hbf5dee05} /* (12, 10, 7) {real, imag} */,
  {32'h3f367234, 32'hbf5df5b2} /* (12, 10, 6) {real, imag} */,
  {32'hbef6ad92, 32'hbeb7651e} /* (12, 10, 5) {real, imag} */,
  {32'h3f0853da, 32'hbf05d9df} /* (12, 10, 4) {real, imag} */,
  {32'h3e83537a, 32'hbf2527bc} /* (12, 10, 3) {real, imag} */,
  {32'h3ee02ccc, 32'hbc51a400} /* (12, 10, 2) {real, imag} */,
  {32'h3e35b1c0, 32'hbf64c2b0} /* (12, 10, 1) {real, imag} */,
  {32'h3e1fd57c, 32'hbe04a418} /* (12, 10, 0) {real, imag} */,
  {32'hbf0568c5, 32'h3f5de200} /* (12, 9, 31) {real, imag} */,
  {32'hbebe4a14, 32'h3dadc2a0} /* (12, 9, 30) {real, imag} */,
  {32'h3f700afd, 32'hbf446089} /* (12, 9, 29) {real, imag} */,
  {32'h3f082f7b, 32'h3d191940} /* (12, 9, 28) {real, imag} */,
  {32'hbe18fa78, 32'hbf1e9388} /* (12, 9, 27) {real, imag} */,
  {32'hbecbb42c, 32'hbf014a3c} /* (12, 9, 26) {real, imag} */,
  {32'hbf767667, 32'hbf6a6d4c} /* (12, 9, 25) {real, imag} */,
  {32'hbfc056f4, 32'h3e0e1230} /* (12, 9, 24) {real, imag} */,
  {32'hbf5551a2, 32'hbe7b15a0} /* (12, 9, 23) {real, imag} */,
  {32'hbf652c7a, 32'hbf3ced58} /* (12, 9, 22) {real, imag} */,
  {32'hbea91f22, 32'hbf86838e} /* (12, 9, 21) {real, imag} */,
  {32'hbe82b8ae, 32'h3dce8300} /* (12, 9, 20) {real, imag} */,
  {32'hbe9fc69c, 32'hbe1b0240} /* (12, 9, 19) {real, imag} */,
  {32'h3f2a4ada, 32'hbe7790f8} /* (12, 9, 18) {real, imag} */,
  {32'h400fee29, 32'h3ed579f0} /* (12, 9, 17) {real, imag} */,
  {32'h3fda1a18, 32'h3e494cf0} /* (12, 9, 16) {real, imag} */,
  {32'h3f412831, 32'hbf8271fe} /* (12, 9, 15) {real, imag} */,
  {32'hbed29af0, 32'hbf31f4b0} /* (12, 9, 14) {real, imag} */,
  {32'hbf6b1242, 32'h3e9a4f18} /* (12, 9, 13) {real, imag} */,
  {32'h3debc168, 32'hbf5f7e50} /* (12, 9, 12) {real, imag} */,
  {32'h3f4c6f3e, 32'hbeeffe88} /* (12, 9, 11) {real, imag} */,
  {32'h3e0db190, 32'hbea3dd43} /* (12, 9, 10) {real, imag} */,
  {32'hbe711cc8, 32'h3e97bb90} /* (12, 9, 9) {real, imag} */,
  {32'h3ef47840, 32'hbef23b18} /* (12, 9, 8) {real, imag} */,
  {32'h3f5310db, 32'hbe6b0898} /* (12, 9, 7) {real, imag} */,
  {32'hbee4e38e, 32'hbde93a70} /* (12, 9, 6) {real, imag} */,
  {32'hbe4c341c, 32'hbe06a0a0} /* (12, 9, 5) {real, imag} */,
  {32'hbc5be910, 32'h3ec49da8} /* (12, 9, 4) {real, imag} */,
  {32'hbe2c8d18, 32'h3d30a080} /* (12, 9, 3) {real, imag} */,
  {32'h3e82365c, 32'hbe8946a0} /* (12, 9, 2) {real, imag} */,
  {32'hbc519e80, 32'h3f1ab7d4} /* (12, 9, 1) {real, imag} */,
  {32'h3f0c3d56, 32'h3f2e3b48} /* (12, 9, 0) {real, imag} */,
  {32'h3d000660, 32'hbe161540} /* (12, 8, 31) {real, imag} */,
  {32'hbe06aee5, 32'hbf4b51b0} /* (12, 8, 30) {real, imag} */,
  {32'h3e8dfee7, 32'hbfd91536} /* (12, 8, 29) {real, imag} */,
  {32'h3c6861d0, 32'hbfcdd4be} /* (12, 8, 28) {real, imag} */,
  {32'h3e172e9c, 32'hbf2bf742} /* (12, 8, 27) {real, imag} */,
  {32'hbdf2dce4, 32'hbf47fb7e} /* (12, 8, 26) {real, imag} */,
  {32'hbf127406, 32'hbfafd663} /* (12, 8, 25) {real, imag} */,
  {32'hbf870c94, 32'h3d5707a0} /* (12, 8, 24) {real, imag} */,
  {32'hbe9ac844, 32'h3f351ff4} /* (12, 8, 23) {real, imag} */,
  {32'h3e40731c, 32'hbf05065c} /* (12, 8, 22) {real, imag} */,
  {32'hbd746d20, 32'hbf06ae43} /* (12, 8, 21) {real, imag} */,
  {32'h3e6b1784, 32'hbd5b9780} /* (12, 8, 20) {real, imag} */,
  {32'hbd53cd86, 32'hbf1ef450} /* (12, 8, 19) {real, imag} */,
  {32'h3f92ed4c, 32'hbf361306} /* (12, 8, 18) {real, imag} */,
  {32'h3fdebd91, 32'h3ea48b38} /* (12, 8, 17) {real, imag} */,
  {32'hbe8dfd58, 32'h3fb78730} /* (12, 8, 16) {real, imag} */,
  {32'hbf8502b9, 32'h3f08f98a} /* (12, 8, 15) {real, imag} */,
  {32'hbf6d4c0a, 32'hbf686b5c} /* (12, 8, 14) {real, imag} */,
  {32'hbf043dd6, 32'hbf1a12c0} /* (12, 8, 13) {real, imag} */,
  {32'h3ea83ecc, 32'hbf15d6c8} /* (12, 8, 12) {real, imag} */,
  {32'h3f35d12a, 32'hbe3c1960} /* (12, 8, 11) {real, imag} */,
  {32'hbf3ff211, 32'h3f46bbf0} /* (12, 8, 10) {real, imag} */,
  {32'hbeec2c0b, 32'h3f7e075e} /* (12, 8, 9) {real, imag} */,
  {32'h3f41b99d, 32'h3dc24878} /* (12, 8, 8) {real, imag} */,
  {32'hbeee83ca, 32'h3e124f88} /* (12, 8, 7) {real, imag} */,
  {32'hbf1f02db, 32'hbea00304} /* (12, 8, 6) {real, imag} */,
  {32'h3f8ed522, 32'hbe3436a0} /* (12, 8, 5) {real, imag} */,
  {32'h3fced698, 32'h3fa55156} /* (12, 8, 4) {real, imag} */,
  {32'h3f6414e1, 32'hbe2f9440} /* (12, 8, 3) {real, imag} */,
  {32'h3eb97934, 32'h3ee98080} /* (12, 8, 2) {real, imag} */,
  {32'hbecb2b90, 32'h3fae6ce8} /* (12, 8, 1) {real, imag} */,
  {32'h3d604450, 32'h3e60fd20} /* (12, 8, 0) {real, imag} */,
  {32'hbf818f55, 32'h3e7cc020} /* (12, 7, 31) {real, imag} */,
  {32'hbf5fb938, 32'h3f8db374} /* (12, 7, 30) {real, imag} */,
  {32'hbd06d940, 32'h3d8387a0} /* (12, 7, 29) {real, imag} */,
  {32'h3e3973a0, 32'hbf560338} /* (12, 7, 28) {real, imag} */,
  {32'h3f2282c8, 32'hbf4bafb4} /* (12, 7, 27) {real, imag} */,
  {32'h3eb2a5b4, 32'hbf78bc80} /* (12, 7, 26) {real, imag} */,
  {32'hbeff4f48, 32'hbfcf9faf} /* (12, 7, 25) {real, imag} */,
  {32'hbf750382, 32'hbf21f76c} /* (12, 7, 24) {real, imag} */,
  {32'h3f35b5fa, 32'h3f930628} /* (12, 7, 23) {real, imag} */,
  {32'h3ed55736, 32'h3f67d258} /* (12, 7, 22) {real, imag} */,
  {32'hbefc9b7b, 32'hbc25ed00} /* (12, 7, 21) {real, imag} */,
  {32'h3f1dae64, 32'hbd031900} /* (12, 7, 20) {real, imag} */,
  {32'hbea3cf18, 32'hbf0aecc4} /* (12, 7, 19) {real, imag} */,
  {32'hbf0f8323, 32'hbe9fb590} /* (12, 7, 18) {real, imag} */,
  {32'hbe384496, 32'h3dce8b60} /* (12, 7, 17) {real, imag} */,
  {32'hbf439124, 32'h3f56687e} /* (12, 7, 16) {real, imag} */,
  {32'hbf38588c, 32'h3f60fe58} /* (12, 7, 15) {real, imag} */,
  {32'hbe95ec7e, 32'hbeb05ab8} /* (12, 7, 14) {real, imag} */,
  {32'h3da53320, 32'hbe60b940} /* (12, 7, 13) {real, imag} */,
  {32'h3eea69c6, 32'hbe418b60} /* (12, 7, 12) {real, imag} */,
  {32'h3e9d8f93, 32'hbe7fc3f8} /* (12, 7, 11) {real, imag} */,
  {32'hbf88a9c8, 32'h3f32f628} /* (12, 7, 10) {real, imag} */,
  {32'hbee3a656, 32'h3e0947a0} /* (12, 7, 9) {real, imag} */,
  {32'h3e0c2974, 32'h3ec76410} /* (12, 7, 8) {real, imag} */,
  {32'h3cc0e620, 32'h3e2d4b40} /* (12, 7, 7) {real, imag} */,
  {32'h3ac8ac00, 32'hbf975464} /* (12, 7, 6) {real, imag} */,
  {32'h3f292f6a, 32'hbf101e20} /* (12, 7, 5) {real, imag} */,
  {32'h3f29f22e, 32'h3f97f41c} /* (12, 7, 4) {real, imag} */,
  {32'h3f1365c5, 32'h3f245330} /* (12, 7, 3) {real, imag} */,
  {32'h3f446be0, 32'h3d3acd40} /* (12, 7, 2) {real, imag} */,
  {32'hbf0ddb12, 32'hbd083740} /* (12, 7, 1) {real, imag} */,
  {32'hbf39e755, 32'hbf0c804c} /* (12, 7, 0) {real, imag} */,
  {32'h3d3a9c90, 32'h3eecc3ec} /* (12, 6, 31) {real, imag} */,
  {32'h3ec6d9e0, 32'h3f6b4170} /* (12, 6, 30) {real, imag} */,
  {32'h3ec1dcca, 32'h3dc2dbc0} /* (12, 6, 29) {real, imag} */,
  {32'hbea9b6f0, 32'h3e642130} /* (12, 6, 28) {real, imag} */,
  {32'h3de89710, 32'hbf16091e} /* (12, 6, 27) {real, imag} */,
  {32'hbedf4f54, 32'hbe24b7f8} /* (12, 6, 26) {real, imag} */,
  {32'hbed24f20, 32'h3dfea120} /* (12, 6, 25) {real, imag} */,
  {32'hbf6ac8ee, 32'hbe722870} /* (12, 6, 24) {real, imag} */,
  {32'hbf8039f1, 32'hbc8ecd00} /* (12, 6, 23) {real, imag} */,
  {32'hbf862f64, 32'h3f65d304} /* (12, 6, 22) {real, imag} */,
  {32'hbec6c654, 32'h3f3e190a} /* (12, 6, 21) {real, imag} */,
  {32'h3f0d9caf, 32'hbefd2d58} /* (12, 6, 20) {real, imag} */,
  {32'h3ed30308, 32'h3e97a0d8} /* (12, 6, 19) {real, imag} */,
  {32'hbdff2a60, 32'h3f8b513d} /* (12, 6, 18) {real, imag} */,
  {32'hbe826946, 32'h3e75e910} /* (12, 6, 17) {real, imag} */,
  {32'hbf2c48cb, 32'hbee19370} /* (12, 6, 16) {real, imag} */,
  {32'hbf1dbd7c, 32'h3e1ddd30} /* (12, 6, 15) {real, imag} */,
  {32'h3eaa3f34, 32'h3f63ec16} /* (12, 6, 14) {real, imag} */,
  {32'hbf0a0b64, 32'h3f5fa9be} /* (12, 6, 13) {real, imag} */,
  {32'hbfbf3f40, 32'h3f75c0c0} /* (12, 6, 12) {real, imag} */,
  {32'hbe7f05b8, 32'h3ef2f398} /* (12, 6, 11) {real, imag} */,
  {32'h3f1d8c36, 32'h3f46e208} /* (12, 6, 10) {real, imag} */,
  {32'h3f436280, 32'h3e977320} /* (12, 6, 9) {real, imag} */,
  {32'hbe211170, 32'hbed6d4c8} /* (12, 6, 8) {real, imag} */,
  {32'h3e05a3e0, 32'hbfbf028a} /* (12, 6, 7) {real, imag} */,
  {32'hbed73d62, 32'hbfa9dbda} /* (12, 6, 6) {real, imag} */,
  {32'hbf0918dd, 32'hbf137808} /* (12, 6, 5) {real, imag} */,
  {32'h3ea34e80, 32'h3efe3c88} /* (12, 6, 4) {real, imag} */,
  {32'hbf304eb6, 32'hbdb62fe0} /* (12, 6, 3) {real, imag} */,
  {32'hbfb4887c, 32'hbf3066a4} /* (12, 6, 2) {real, imag} */,
  {32'hbfbeeddc, 32'hbeb58aa8} /* (12, 6, 1) {real, imag} */,
  {32'hbe92e4c0, 32'hbee80b2d} /* (12, 6, 0) {real, imag} */,
  {32'h3e1d5188, 32'hbde58280} /* (12, 5, 31) {real, imag} */,
  {32'h3e312dd0, 32'h3f8dd0fe} /* (12, 5, 30) {real, imag} */,
  {32'h3e5d0160, 32'h3f356a24} /* (12, 5, 29) {real, imag} */,
  {32'hbfaf1a02, 32'h3f204204} /* (12, 5, 28) {real, imag} */,
  {32'hbe809ff0, 32'h3ec9bd68} /* (12, 5, 27) {real, imag} */,
  {32'h3f0b85a1, 32'hbe9dd3b6} /* (12, 5, 26) {real, imag} */,
  {32'h3f764d7f, 32'hbca55e00} /* (12, 5, 25) {real, imag} */,
  {32'hbedf504e, 32'h3ba12200} /* (12, 5, 24) {real, imag} */,
  {32'hbf68ff3d, 32'hbf3044d0} /* (12, 5, 23) {real, imag} */,
  {32'h3f1631fc, 32'hbe579930} /* (12, 5, 22) {real, imag} */,
  {32'h3e3d59c0, 32'h3fb43912} /* (12, 5, 21) {real, imag} */,
  {32'h3ec2445e, 32'hbf0a7368} /* (12, 5, 20) {real, imag} */,
  {32'h3f7d2454, 32'hbeee5f7d} /* (12, 5, 19) {real, imag} */,
  {32'hbf176a76, 32'h3f0b926c} /* (12, 5, 18) {real, imag} */,
  {32'hbf2c83bd, 32'h3f5fe219} /* (12, 5, 17) {real, imag} */,
  {32'hbd67fad0, 32'hbe6069d7} /* (12, 5, 16) {real, imag} */,
  {32'h3ea26ada, 32'hbacb9c00} /* (12, 5, 15) {real, imag} */,
  {32'h3ee721d7, 32'h3f37e5e9} /* (12, 5, 14) {real, imag} */,
  {32'hbe00489e, 32'h3f001752} /* (12, 5, 13) {real, imag} */,
  {32'hbe5b1cf0, 32'hbb925000} /* (12, 5, 12) {real, imag} */,
  {32'h3e8c9034, 32'hbf093ed0} /* (12, 5, 11) {real, imag} */,
  {32'h4013aba2, 32'h3d88e3e0} /* (12, 5, 10) {real, imag} */,
  {32'h3f83c1c2, 32'h3f86b403} /* (12, 5, 9) {real, imag} */,
  {32'h3cb07660, 32'h3f0b5316} /* (12, 5, 8) {real, imag} */,
  {32'hbe7d4af4, 32'hbf913c50} /* (12, 5, 7) {real, imag} */,
  {32'hbfa8f162, 32'hbfc1e55f} /* (12, 5, 6) {real, imag} */,
  {32'hbe4c3454, 32'h3ee794d8} /* (12, 5, 5) {real, imag} */,
  {32'h3e5dbd30, 32'h3f2a4f88} /* (12, 5, 4) {real, imag} */,
  {32'hbf313bb4, 32'hbf7248a0} /* (12, 5, 3) {real, imag} */,
  {32'hbfabc56f, 32'h3c8edb00} /* (12, 5, 2) {real, imag} */,
  {32'hbefe25ee, 32'h3f3d4fca} /* (12, 5, 1) {real, imag} */,
  {32'h3ec76440, 32'hbf182672} /* (12, 5, 0) {real, imag} */,
  {32'hbf21a6cd, 32'hbe5e4fc0} /* (12, 4, 31) {real, imag} */,
  {32'hbf4291b2, 32'hb97dc000} /* (12, 4, 30) {real, imag} */,
  {32'hbe6d4a20, 32'h3d9a69c0} /* (12, 4, 29) {real, imag} */,
  {32'hbec355af, 32'h3f20c3c4} /* (12, 4, 28) {real, imag} */,
  {32'hbee9c816, 32'h3f8372e0} /* (12, 4, 27) {real, imag} */,
  {32'hbeccd9f8, 32'hbe1fc8b0} /* (12, 4, 26) {real, imag} */,
  {32'h3fa49f7a, 32'hbf3b1574} /* (12, 4, 25) {real, imag} */,
  {32'h3f62fa42, 32'hbf3021d2} /* (12, 4, 24) {real, imag} */,
  {32'h3f219e77, 32'hbeddd778} /* (12, 4, 23) {real, imag} */,
  {32'h3f6b3888, 32'hbf160e44} /* (12, 4, 22) {real, imag} */,
  {32'h3de3fa00, 32'h3f016754} /* (12, 4, 21) {real, imag} */,
  {32'h3e5ac110, 32'hbf5cd2c8} /* (12, 4, 20) {real, imag} */,
  {32'hbe63b748, 32'hbf63f958} /* (12, 4, 19) {real, imag} */,
  {32'hbf864ad1, 32'h3e878b90} /* (12, 4, 18) {real, imag} */,
  {32'hbe241e20, 32'h3f48fd78} /* (12, 4, 17) {real, imag} */,
  {32'h3ec1b800, 32'hbe164df0} /* (12, 4, 16) {real, imag} */,
  {32'h3f3e8d14, 32'hbe7508d0} /* (12, 4, 15) {real, imag} */,
  {32'h3f4c2076, 32'hbeeb7e60} /* (12, 4, 14) {real, imag} */,
  {32'h3e82935d, 32'h3e047510} /* (12, 4, 13) {real, imag} */,
  {32'h3f1eaff8, 32'h3f2cdc78} /* (12, 4, 12) {real, imag} */,
  {32'h3ede1b8a, 32'hbe90d848} /* (12, 4, 11) {real, imag} */,
  {32'h3f5c1086, 32'h3e474d90} /* (12, 4, 10) {real, imag} */,
  {32'hbdf97f10, 32'h3e5ad120} /* (12, 4, 9) {real, imag} */,
  {32'hbf9510e2, 32'hbf28d03c} /* (12, 4, 8) {real, imag} */,
  {32'hbf308a92, 32'hbe814448} /* (12, 4, 7) {real, imag} */,
  {32'h3ef38895, 32'hbeaaad74} /* (12, 4, 6) {real, imag} */,
  {32'h3fb162b0, 32'h3f3c91d1} /* (12, 4, 5) {real, imag} */,
  {32'h3fa3c0dd, 32'h3f3953a0} /* (12, 4, 4) {real, imag} */,
  {32'h3e4dd4cc, 32'hbf708aba} /* (12, 4, 3) {real, imag} */,
  {32'hbf2d3b48, 32'h3e79c750} /* (12, 4, 2) {real, imag} */,
  {32'hbec403fa, 32'h3ed72318} /* (12, 4, 1) {real, imag} */,
  {32'h3d801320, 32'hbcd45ac0} /* (12, 4, 0) {real, imag} */,
  {32'hbebce9f0, 32'hbf7cddee} /* (12, 3, 31) {real, imag} */,
  {32'hbebf69ec, 32'hbef8b5dc} /* (12, 3, 30) {real, imag} */,
  {32'h3e5f1280, 32'hbda0e970} /* (12, 3, 29) {real, imag} */,
  {32'h3e5c8b80, 32'h3ed07488} /* (12, 3, 28) {real, imag} */,
  {32'hbeb65a5c, 32'h3ee787f0} /* (12, 3, 27) {real, imag} */,
  {32'hbe8cc378, 32'h3ec85a00} /* (12, 3, 26) {real, imag} */,
  {32'h3ef93446, 32'hbea517e0} /* (12, 3, 25) {real, imag} */,
  {32'h3e9b9e50, 32'h3eb518e8} /* (12, 3, 24) {real, imag} */,
  {32'hbf1619dc, 32'h3f00c518} /* (12, 3, 23) {real, imag} */,
  {32'hbf6aa2d4, 32'hbf17ff28} /* (12, 3, 22) {real, imag} */,
  {32'hbb50a400, 32'hbeb6f938} /* (12, 3, 21) {real, imag} */,
  {32'h3ee79ee0, 32'hbe3f2e80} /* (12, 3, 20) {real, imag} */,
  {32'h3f2228b6, 32'hbdc0e2a0} /* (12, 3, 19) {real, imag} */,
  {32'h3d3f88c0, 32'h3f663f4c} /* (12, 3, 18) {real, imag} */,
  {32'h3d81ac40, 32'h3e07f1c0} /* (12, 3, 17) {real, imag} */,
  {32'hbe38f088, 32'hbf34f43d} /* (12, 3, 16) {real, imag} */,
  {32'h3ea676be, 32'hbe146a08} /* (12, 3, 15) {real, imag} */,
  {32'h3eca73a4, 32'hbfb3fd67} /* (12, 3, 14) {real, imag} */,
  {32'hbee67e08, 32'hbf96212c} /* (12, 3, 13) {real, imag} */,
  {32'hbcc9d180, 32'h3fa22394} /* (12, 3, 12) {real, imag} */,
  {32'hbf57b41e, 32'h3df975a0} /* (12, 3, 11) {real, imag} */,
  {32'hbf6010a2, 32'hbf8ee702} /* (12, 3, 10) {real, imag} */,
  {32'hbf295baf, 32'hbfabff22} /* (12, 3, 9) {real, imag} */,
  {32'hbec24d20, 32'hbfbdeae6} /* (12, 3, 8) {real, imag} */,
  {32'hbdae7400, 32'hbdd29680} /* (12, 3, 7) {real, imag} */,
  {32'h3dfddaec, 32'h3f26851a} /* (12, 3, 6) {real, imag} */,
  {32'h3f098824, 32'h3fbe81b6} /* (12, 3, 5) {real, imag} */,
  {32'h3f527e74, 32'h3ff36fe1} /* (12, 3, 4) {real, imag} */,
  {32'h3eaf7bd4, 32'h3f5ddb10} /* (12, 3, 3) {real, imag} */,
  {32'hbf3bffd2, 32'h3ef6634c} /* (12, 3, 2) {real, imag} */,
  {32'hbf397252, 32'hbe589bfc} /* (12, 3, 1) {real, imag} */,
  {32'h3e13bc26, 32'hbe363a34} /* (12, 3, 0) {real, imag} */,
  {32'hbcbd3810, 32'hbe182ff0} /* (12, 2, 31) {real, imag} */,
  {32'h3e82e1de, 32'h3f6b79c4} /* (12, 2, 30) {real, imag} */,
  {32'h3fba9806, 32'h3f7e3660} /* (12, 2, 29) {real, imag} */,
  {32'h3ffc756c, 32'hbda175e0} /* (12, 2, 28) {real, imag} */,
  {32'h3f3deeb0, 32'hbdd0f700} /* (12, 2, 27) {real, imag} */,
  {32'h3f07017c, 32'h3e53d4d0} /* (12, 2, 26) {real, imag} */,
  {32'hbf59db14, 32'hbf39a93a} /* (12, 2, 25) {real, imag} */,
  {32'hbf412775, 32'hbf08a4ee} /* (12, 2, 24) {real, imag} */,
  {32'hbf1e29c4, 32'h3eb1d9e4} /* (12, 2, 23) {real, imag} */,
  {32'hbf17f207, 32'hbf82337e} /* (12, 2, 22) {real, imag} */,
  {32'h3f1a7862, 32'hbfc597c1} /* (12, 2, 21) {real, imag} */,
  {32'h3edb2815, 32'hbf663460} /* (12, 2, 20) {real, imag} */,
  {32'hbe1d6e98, 32'hbefe4a30} /* (12, 2, 19) {real, imag} */,
  {32'hbed876a8, 32'h3f90fd8e} /* (12, 2, 18) {real, imag} */,
  {32'hbd3ba4c0, 32'h3effe000} /* (12, 2, 17) {real, imag} */,
  {32'h3d0bf890, 32'hbef6dd40} /* (12, 2, 16) {real, imag} */,
  {32'hbdaa2c10, 32'hbe17a008} /* (12, 2, 15) {real, imag} */,
  {32'hbf128f74, 32'hc0119dd8} /* (12, 2, 14) {real, imag} */,
  {32'hbf27fd38, 32'hbf8a6fb8} /* (12, 2, 13) {real, imag} */,
  {32'hbee2ebc4, 32'h3edc55b8} /* (12, 2, 12) {real, imag} */,
  {32'hbf18512e, 32'hbe552350} /* (12, 2, 11) {real, imag} */,
  {32'h3e2b96a0, 32'hbf38ddfc} /* (12, 2, 10) {real, imag} */,
  {32'h3f1cc16e, 32'hbf51eb28} /* (12, 2, 9) {real, imag} */,
  {32'h3ea98746, 32'hbf53bcec} /* (12, 2, 8) {real, imag} */,
  {32'h3ee762a8, 32'hbea6fad0} /* (12, 2, 7) {real, imag} */,
  {32'hbf1b7c26, 32'h3dac87e0} /* (12, 2, 6) {real, imag} */,
  {32'h3f660cc6, 32'h3e482950} /* (12, 2, 5) {real, imag} */,
  {32'h3fa2bb68, 32'h3f83b8d8} /* (12, 2, 4) {real, imag} */,
  {32'h3f1c1a27, 32'h3e436060} /* (12, 2, 3) {real, imag} */,
  {32'hbdbfd6dd, 32'h3a941400} /* (12, 2, 2) {real, imag} */,
  {32'h3e8a5700, 32'h3dbfb7d0} /* (12, 2, 1) {real, imag} */,
  {32'h3ea8e26a, 32'h3e135f50} /* (12, 2, 0) {real, imag} */,
  {32'hbcfd5380, 32'hbf1c4a8a} /* (12, 1, 31) {real, imag} */,
  {32'h3f01a9a2, 32'hbea45cb0} /* (12, 1, 30) {real, imag} */,
  {32'h3f908e82, 32'hbc1d2580} /* (12, 1, 29) {real, imag} */,
  {32'h3fa07772, 32'hbdb97a40} /* (12, 1, 28) {real, imag} */,
  {32'h3f7d1216, 32'hbf2fc4ff} /* (12, 1, 27) {real, imag} */,
  {32'h3f0cdddc, 32'h3e055be0} /* (12, 1, 26) {real, imag} */,
  {32'hbed5a468, 32'hbf3b11f2} /* (12, 1, 25) {real, imag} */,
  {32'hbe34de50, 32'hbf19ca46} /* (12, 1, 24) {real, imag} */,
  {32'h3e5d6570, 32'h3ef36c88} /* (12, 1, 23) {real, imag} */,
  {32'hbf8cd6ae, 32'hbf4d09cc} /* (12, 1, 22) {real, imag} */,
  {32'hbf379d67, 32'hbef1b668} /* (12, 1, 21) {real, imag} */,
  {32'h3e7cd8f2, 32'h3f08c326} /* (12, 1, 20) {real, imag} */,
  {32'hbeb147a8, 32'hbe181b18} /* (12, 1, 19) {real, imag} */,
  {32'hbf272818, 32'h3e1b61e0} /* (12, 1, 18) {real, imag} */,
  {32'hbf1094e2, 32'h3f9c466a} /* (12, 1, 17) {real, imag} */,
  {32'h3e4d5f20, 32'h3f219b82} /* (12, 1, 16) {real, imag} */,
  {32'h3ef5de05, 32'hbf071423} /* (12, 1, 15) {real, imag} */,
  {32'hbeb72cd8, 32'hc003d204} /* (12, 1, 14) {real, imag} */,
  {32'hbf4f96fc, 32'hbea53d38} /* (12, 1, 13) {real, imag} */,
  {32'hbf0eb604, 32'h3f4b9140} /* (12, 1, 12) {real, imag} */,
  {32'h3f3d8578, 32'h3ea328e0} /* (12, 1, 11) {real, imag} */,
  {32'h3fe4f827, 32'hbf07c8f0} /* (12, 1, 10) {real, imag} */,
  {32'h3f0d07cf, 32'h3e6f5b80} /* (12, 1, 9) {real, imag} */,
  {32'h3de988f0, 32'h3f0fcc32} /* (12, 1, 8) {real, imag} */,
  {32'h3e0cfc88, 32'hbf26f9fa} /* (12, 1, 7) {real, imag} */,
  {32'hbe4d8680, 32'hbf4f2440} /* (12, 1, 6) {real, imag} */,
  {32'h3fdddb24, 32'hbf5d8a53} /* (12, 1, 5) {real, imag} */,
  {32'h3fd59a80, 32'h3f33329a} /* (12, 1, 4) {real, imag} */,
  {32'hbc2379e0, 32'h3f528048} /* (12, 1, 3) {real, imag} */,
  {32'hbf04eaf6, 32'h3e857904} /* (12, 1, 2) {real, imag} */,
  {32'hbca05280, 32'h3e637648} /* (12, 1, 1) {real, imag} */,
  {32'h3e30a084, 32'hbe0a9c14} /* (12, 1, 0) {real, imag} */,
  {32'hbf1d3d21, 32'hbecafc4c} /* (12, 0, 31) {real, imag} */,
  {32'hbe8639bc, 32'hbe7fad70} /* (12, 0, 30) {real, imag} */,
  {32'h3ece1524, 32'h3e868a5e} /* (12, 0, 29) {real, imag} */,
  {32'h3ebb5e1c, 32'hbdab4d40} /* (12, 0, 28) {real, imag} */,
  {32'h3f00b9f8, 32'hbf959728} /* (12, 0, 27) {real, imag} */,
  {32'h3e572198, 32'hbe0b18be} /* (12, 0, 26) {real, imag} */,
  {32'h3e412248, 32'hbf27caa4} /* (12, 0, 25) {real, imag} */,
  {32'h3ef6aeb4, 32'hbf2f6c60} /* (12, 0, 24) {real, imag} */,
  {32'h3eb3f2cc, 32'h3dcfb2d0} /* (12, 0, 23) {real, imag} */,
  {32'hbef07e90, 32'hbe124fa8} /* (12, 0, 22) {real, imag} */,
  {32'hbf080cf6, 32'hbd480cc0} /* (12, 0, 21) {real, imag} */,
  {32'hbe2d106c, 32'h3f59ec78} /* (12, 0, 20) {real, imag} */,
  {32'h3d9aabb0, 32'h3eeb37fa} /* (12, 0, 19) {real, imag} */,
  {32'h3f10c336, 32'hbe1b3598} /* (12, 0, 18) {real, imag} */,
  {32'h3e266b6f, 32'h3f4eef93} /* (12, 0, 17) {real, imag} */,
  {32'hbf0ab20c, 32'h3f13af55} /* (12, 0, 16) {real, imag} */,
  {32'h3eaa510c, 32'h3e04d84c} /* (12, 0, 15) {real, imag} */,
  {32'h3f1cd000, 32'hbf11783e} /* (12, 0, 14) {real, imag} */,
  {32'hbd9b83c0, 32'h3e707678} /* (12, 0, 13) {real, imag} */,
  {32'h3efc5402, 32'h3f117430} /* (12, 0, 12) {real, imag} */,
  {32'h3f8118d3, 32'hbdf27260} /* (12, 0, 11) {real, imag} */,
  {32'h3f01d284, 32'hbf36f7ca} /* (12, 0, 10) {real, imag} */,
  {32'h3dcb5600, 32'hbef41328} /* (12, 0, 9) {real, imag} */,
  {32'hbeafa064, 32'h3eeb2bf4} /* (12, 0, 8) {real, imag} */,
  {32'hbf0948d7, 32'hbe53a1a0} /* (12, 0, 7) {real, imag} */,
  {32'hbef2e922, 32'hbeee896c} /* (12, 0, 6) {real, imag} */,
  {32'h3f1fbf32, 32'hbe56a6ae} /* (12, 0, 5) {real, imag} */,
  {32'h3ea5954e, 32'hbe51ae40} /* (12, 0, 4) {real, imag} */,
  {32'hbce4ac98, 32'h3f152214} /* (12, 0, 3) {real, imag} */,
  {32'h3e711d70, 32'h3ef4e530} /* (12, 0, 2) {real, imag} */,
  {32'h3f128a50, 32'h3eda6ea0} /* (12, 0, 1) {real, imag} */,
  {32'h3eb1a2c0, 32'h3e60fec6} /* (12, 0, 0) {real, imag} */,
  {32'h3ee45ab2, 32'hbe8936a6} /* (11, 31, 31) {real, imag} */,
  {32'h3e8e9cac, 32'hbf173560} /* (11, 31, 30) {real, imag} */,
  {32'hbee079ac, 32'h3e4de958} /* (11, 31, 29) {real, imag} */,
  {32'hbeb8fd02, 32'h3f439618} /* (11, 31, 28) {real, imag} */,
  {32'h3eb3fba8, 32'h3fd2f65c} /* (11, 31, 27) {real, imag} */,
  {32'h3e1b6a38, 32'h3f72d37c} /* (11, 31, 26) {real, imag} */,
  {32'hbf25ad96, 32'hbe96a1e8} /* (11, 31, 25) {real, imag} */,
  {32'h3f26a079, 32'h3df2ed50} /* (11, 31, 24) {real, imag} */,
  {32'h3ec7c1a1, 32'hbf32f827} /* (11, 31, 23) {real, imag} */,
  {32'h3e302226, 32'hbe769e50} /* (11, 31, 22) {real, imag} */,
  {32'hbeadcf8c, 32'h3e592114} /* (11, 31, 21) {real, imag} */,
  {32'hbef994a8, 32'h3f36dc53} /* (11, 31, 20) {real, imag} */,
  {32'hbf02ec64, 32'h3eef592e} /* (11, 31, 19) {real, imag} */,
  {32'hbf15bbdd, 32'hbe1de9f8} /* (11, 31, 18) {real, imag} */,
  {32'hbed98b07, 32'hbe3008b8} /* (11, 31, 17) {real, imag} */,
  {32'hbe920715, 32'h3e787330} /* (11, 31, 16) {real, imag} */,
  {32'h3e0b9170, 32'h3d051246} /* (11, 31, 15) {real, imag} */,
  {32'h3e46c07e, 32'h3d4de050} /* (11, 31, 14) {real, imag} */,
  {32'hbe968b28, 32'h3fc3a1d4} /* (11, 31, 13) {real, imag} */,
  {32'hbef87b80, 32'h3fc613d4} /* (11, 31, 12) {real, imag} */,
  {32'h3e2915ee, 32'h3c858460} /* (11, 31, 11) {real, imag} */,
  {32'h3f2afa57, 32'h3f354702} /* (11, 31, 10) {real, imag} */,
  {32'h3db02f00, 32'h3dec6648} /* (11, 31, 9) {real, imag} */,
  {32'h3d532920, 32'hbe07ee2e} /* (11, 31, 8) {real, imag} */,
  {32'h3ec11dc0, 32'hbe179ddc} /* (11, 31, 7) {real, imag} */,
  {32'h3ee8b938, 32'hbf35a900} /* (11, 31, 6) {real, imag} */,
  {32'h3f4c918e, 32'hbf405ec5} /* (11, 31, 5) {real, imag} */,
  {32'h3dbcff0c, 32'hbf4a931c} /* (11, 31, 4) {real, imag} */,
  {32'h3f218dce, 32'hbf0d5cf0} /* (11, 31, 3) {real, imag} */,
  {32'h3f6d74f2, 32'hbf796c86} /* (11, 31, 2) {real, imag} */,
  {32'h3fa3058c, 32'hbf9f9275} /* (11, 31, 1) {real, imag} */,
  {32'h3fa11899, 32'hbd74efb4} /* (11, 31, 0) {real, imag} */,
  {32'hbd95a150, 32'h3e9964ad} /* (11, 30, 31) {real, imag} */,
  {32'h3f6e7b04, 32'hbf772adc} /* (11, 30, 30) {real, imag} */,
  {32'h3e8084c0, 32'hbfa57734} /* (11, 30, 29) {real, imag} */,
  {32'h3ce10540, 32'hbe96b160} /* (11, 30, 28) {real, imag} */,
  {32'h3f5c04d8, 32'h3fa44d9a} /* (11, 30, 27) {real, imag} */,
  {32'h3f9a62e2, 32'h3fa159d2} /* (11, 30, 26) {real, imag} */,
  {32'hbeaf43f4, 32'hbf0a9096} /* (11, 30, 25) {real, imag} */,
  {32'h3e9fc3e0, 32'hbf87fdf0} /* (11, 30, 24) {real, imag} */,
  {32'h3f19681b, 32'hbff98378} /* (11, 30, 23) {real, imag} */,
  {32'h3e0db840, 32'hbfb71e36} /* (11, 30, 22) {real, imag} */,
  {32'hbed42814, 32'h3e13f7fa} /* (11, 30, 21) {real, imag} */,
  {32'hbf16afec, 32'h3fc5e5ea} /* (11, 30, 20) {real, imag} */,
  {32'h3ed9c9b8, 32'h3f6553ea} /* (11, 30, 19) {real, imag} */,
  {32'h3e05e064, 32'hbc89b4c0} /* (11, 30, 18) {real, imag} */,
  {32'hbf8f2f3e, 32'hbdd25640} /* (11, 30, 17) {real, imag} */,
  {32'hbe7ce174, 32'h3f605f18} /* (11, 30, 16) {real, imag} */,
  {32'hbeb20a0a, 32'h3d67a600} /* (11, 30, 15) {real, imag} */,
  {32'hbf2343ed, 32'h3e726970} /* (11, 30, 14) {real, imag} */,
  {32'hbeeea3fa, 32'h3fe8f199} /* (11, 30, 13) {real, imag} */,
  {32'h3e26024c, 32'h3fa3993a} /* (11, 30, 12) {real, imag} */,
  {32'h3f939a80, 32'hbf78a0b0} /* (11, 30, 11) {real, imag} */,
  {32'h3fa4bab2, 32'hbefe11c1} /* (11, 30, 10) {real, imag} */,
  {32'hbdfecbb0, 32'hbea90070} /* (11, 30, 9) {real, imag} */,
  {32'hbec86df4, 32'hbf397df8} /* (11, 30, 8) {real, imag} */,
  {32'h3f8220f4, 32'hbdc8f0e0} /* (11, 30, 7) {real, imag} */,
  {32'h3f6186a2, 32'hbf51d9e8} /* (11, 30, 6) {real, imag} */,
  {32'h3fa00103, 32'hbfcf96e4} /* (11, 30, 5) {real, imag} */,
  {32'h3e39cc25, 32'hbfb602a5} /* (11, 30, 4) {real, imag} */,
  {32'h3ed04a18, 32'hbf5ccfad} /* (11, 30, 3) {real, imag} */,
  {32'h3f386d50, 32'hbfbbd2ad} /* (11, 30, 2) {real, imag} */,
  {32'h3ffd6ebc, 32'hbf969c81} /* (11, 30, 1) {real, imag} */,
  {32'h3ff70deb, 32'hbe9c2aca} /* (11, 30, 0) {real, imag} */,
  {32'h3e8082ee, 32'h3f983ccf} /* (11, 29, 31) {real, imag} */,
  {32'h3f8711fe, 32'h3df6ffb0} /* (11, 29, 30) {real, imag} */,
  {32'h3e1891b8, 32'hbfb0e621} /* (11, 29, 29) {real, imag} */,
  {32'h3f48f2c6, 32'hbfc622f0} /* (11, 29, 28) {real, imag} */,
  {32'h3fc69619, 32'hbfddb2e9} /* (11, 29, 27) {real, imag} */,
  {32'h3ee79fc2, 32'hbf9fd406} /* (11, 29, 26) {real, imag} */,
  {32'hbf8db9fa, 32'hbfccfb96} /* (11, 29, 25) {real, imag} */,
  {32'h3f8bb6ea, 32'hc015971e} /* (11, 29, 24) {real, imag} */,
  {32'h4033e720, 32'hbfdf2600} /* (11, 29, 23) {real, imag} */,
  {32'h3fa0e10d, 32'hbffb8452} /* (11, 29, 22) {real, imag} */,
  {32'h3f36cf72, 32'hbfdec9d2} /* (11, 29, 21) {real, imag} */,
  {32'hbdbb9ff8, 32'hbe335380} /* (11, 29, 20) {real, imag} */,
  {32'h3f39c7f0, 32'h3f0093b0} /* (11, 29, 19) {real, imag} */,
  {32'hbeaf6ee8, 32'hbe5b2460} /* (11, 29, 18) {real, imag} */,
  {32'hbf69503a, 32'hbe7649c8} /* (11, 29, 17) {real, imag} */,
  {32'hbf02ed78, 32'h3f0d99d4} /* (11, 29, 16) {real, imag} */,
  {32'hbf99ed94, 32'h3eed0634} /* (11, 29, 15) {real, imag} */,
  {32'hc00e6094, 32'h3f232408} /* (11, 29, 14) {real, imag} */,
  {32'hbff43262, 32'h3f3b1af1} /* (11, 29, 13) {real, imag} */,
  {32'h3dd371c0, 32'hbf0afc96} /* (11, 29, 12) {real, imag} */,
  {32'h3f8cad34, 32'hbf8e26dd} /* (11, 29, 11) {real, imag} */,
  {32'h3fb5cc9f, 32'hbd32d090} /* (11, 29, 10) {real, imag} */,
  {32'h3f700bb8, 32'hbf29ec0e} /* (11, 29, 9) {real, imag} */,
  {32'h3f86b129, 32'hbf53a6a2} /* (11, 29, 8) {real, imag} */,
  {32'h3f82eeb2, 32'hbf26a014} /* (11, 29, 7) {real, imag} */,
  {32'h3fd1a26d, 32'hbfacfce9} /* (11, 29, 6) {real, imag} */,
  {32'h3fc7c7db, 32'hbfa3cda4} /* (11, 29, 5) {real, imag} */,
  {32'h3ec69448, 32'hbf2d33c0} /* (11, 29, 4) {real, imag} */,
  {32'hbc8480b0, 32'hbee3ad08} /* (11, 29, 3) {real, imag} */,
  {32'h3e13d660, 32'hbf0d33a1} /* (11, 29, 2) {real, imag} */,
  {32'h3f9d7eb2, 32'h3f123fe2} /* (11, 29, 1) {real, imag} */,
  {32'h3f381d4e, 32'h3f4c9438} /* (11, 29, 0) {real, imag} */,
  {32'h3f18d2ae, 32'hbebe2b5a} /* (11, 28, 31) {real, imag} */,
  {32'h3fc5e3d2, 32'hbfbd48ae} /* (11, 28, 30) {real, imag} */,
  {32'h3f11c2a8, 32'hbfac67f8} /* (11, 28, 29) {real, imag} */,
  {32'h3eabf93e, 32'hbf9b7eff} /* (11, 28, 28) {real, imag} */,
  {32'h3fb7536e, 32'hc003c887} /* (11, 28, 27) {real, imag} */,
  {32'h3f71aa41, 32'hbfaa6d69} /* (11, 28, 26) {real, imag} */,
  {32'h3f14362e, 32'hbfb3aad5} /* (11, 28, 25) {real, imag} */,
  {32'h3ffbc480, 32'hc0168567} /* (11, 28, 24) {real, imag} */,
  {32'h403b3f82, 32'hbfa9911b} /* (11, 28, 23) {real, imag} */,
  {32'h3fe20faf, 32'hbeb7c7b6} /* (11, 28, 22) {real, imag} */,
  {32'h3f055d50, 32'h3e785980} /* (11, 28, 21) {real, imag} */,
  {32'hbfd70469, 32'h3ec97024} /* (11, 28, 20) {real, imag} */,
  {32'hbf82edff, 32'h3f192bb6} /* (11, 28, 19) {real, imag} */,
  {32'hc008f4ae, 32'h3f52150c} /* (11, 28, 18) {real, imag} */,
  {32'hbf618b99, 32'h3f2687b2} /* (11, 28, 17) {real, imag} */,
  {32'hbf24908c, 32'h3d9ecaa0} /* (11, 28, 16) {real, imag} */,
  {32'hbfae7ab9, 32'h3e1f0ae8} /* (11, 28, 15) {real, imag} */,
  {32'hbfa437e5, 32'hbe1ca394} /* (11, 28, 14) {real, imag} */,
  {32'hc001e644, 32'h3ea640ac} /* (11, 28, 13) {real, imag} */,
  {32'hbdbf7838, 32'hbe9b664a} /* (11, 28, 12) {real, imag} */,
  {32'h3f20e36a, 32'hbf84a656} /* (11, 28, 11) {real, imag} */,
  {32'h3fc28e14, 32'h3eaf78e8} /* (11, 28, 10) {real, imag} */,
  {32'h400efa56, 32'hbe6b53b0} /* (11, 28, 9) {real, imag} */,
  {32'h40148e14, 32'hbf776fc6} /* (11, 28, 8) {real, imag} */,
  {32'h3f7f0278, 32'hbfa1dde6} /* (11, 28, 7) {real, imag} */,
  {32'h3fc404d0, 32'hbf82a731} /* (11, 28, 6) {real, imag} */,
  {32'h3f2e072e, 32'hbfe8cbe1} /* (11, 28, 5) {real, imag} */,
  {32'h3ee0bc1a, 32'hbf15d824} /* (11, 28, 4) {real, imag} */,
  {32'h3f6f0ffc, 32'hbe95ad84} /* (11, 28, 3) {real, imag} */,
  {32'h3ee9d1d8, 32'h3d30e0c0} /* (11, 28, 2) {real, imag} */,
  {32'h3f9d4284, 32'h3f3715d2} /* (11, 28, 1) {real, imag} */,
  {32'h3f7b836d, 32'h3f5de384} /* (11, 28, 0) {real, imag} */,
  {32'hbde5e940, 32'hbf617af3} /* (11, 27, 31) {real, imag} */,
  {32'h3e375584, 32'hbfc3469a} /* (11, 27, 30) {real, imag} */,
  {32'hbeefd996, 32'hbf40eafa} /* (11, 27, 29) {real, imag} */,
  {32'h3e048780, 32'hbf96b61a} /* (11, 27, 28) {real, imag} */,
  {32'h3f004ef8, 32'hc02aa90a} /* (11, 27, 27) {real, imag} */,
  {32'h3e1b4a0c, 32'hbf06e286} /* (11, 27, 26) {real, imag} */,
  {32'h4006a890, 32'hbf65ad54} /* (11, 27, 25) {real, imag} */,
  {32'h40022b4e, 32'hbfc4eef2} /* (11, 27, 24) {real, imag} */,
  {32'h3f043e3d, 32'hbd99e808} /* (11, 27, 23) {real, imag} */,
  {32'hb96fa000, 32'h3ed3b442} /* (11, 27, 22) {real, imag} */,
  {32'hbe100574, 32'h3ee2e944} /* (11, 27, 21) {real, imag} */,
  {32'hc03caab7, 32'h3f96167c} /* (11, 27, 20) {real, imag} */,
  {32'hc03709b7, 32'h3f83d387} /* (11, 27, 19) {real, imag} */,
  {32'hbff6313b, 32'h3f6007b6} /* (11, 27, 18) {real, imag} */,
  {32'hbef16480, 32'h3fb95b90} /* (11, 27, 17) {real, imag} */,
  {32'hbf190a0a, 32'h3f9d5a98} /* (11, 27, 16) {real, imag} */,
  {32'hbfc14ad2, 32'h3f661717} /* (11, 27, 15) {real, imag} */,
  {32'hbf749827, 32'hbf20bd6d} /* (11, 27, 14) {real, imag} */,
  {32'hbf42024c, 32'h3f3e1cdb} /* (11, 27, 13) {real, imag} */,
  {32'hbe211440, 32'h3f1f3c54} /* (11, 27, 12) {real, imag} */,
  {32'h3f18b91d, 32'h3ce8cf80} /* (11, 27, 11) {real, imag} */,
  {32'h3f3f320c, 32'hbe337548} /* (11, 27, 10) {real, imag} */,
  {32'h3fdee510, 32'hbf8f4461} /* (11, 27, 9) {real, imag} */,
  {32'h40171e96, 32'hbd9ae770} /* (11, 27, 8) {real, imag} */,
  {32'h3fabe143, 32'hbf3d1526} /* (11, 27, 7) {real, imag} */,
  {32'h3ff9c2f8, 32'hbf5d9545} /* (11, 27, 6) {real, imag} */,
  {32'h3f3b9f73, 32'hbfcf5473} /* (11, 27, 5) {real, imag} */,
  {32'hbdacc2ac, 32'hbe9317a8} /* (11, 27, 4) {real, imag} */,
  {32'h3f80cb62, 32'hbf78b7f2} /* (11, 27, 3) {real, imag} */,
  {32'h3f03b86e, 32'hbf0c2b87} /* (11, 27, 2) {real, imag} */,
  {32'h3f8bd1a7, 32'h3e1b1bac} /* (11, 27, 1) {real, imag} */,
  {32'h3f82109c, 32'hbe6cf8d0} /* (11, 27, 0) {real, imag} */,
  {32'hbe68a545, 32'hbf0a7cf3} /* (11, 26, 31) {real, imag} */,
  {32'hbc98cda0, 32'hbf0ab17e} /* (11, 26, 30) {real, imag} */,
  {32'h3ea6e394, 32'hbfa23c9a} /* (11, 26, 29) {real, imag} */,
  {32'h3fc1b45d, 32'hbff15f35} /* (11, 26, 28) {real, imag} */,
  {32'h3e294f88, 32'hbf3002f2} /* (11, 26, 27) {real, imag} */,
  {32'hbf89090e, 32'h3f12bdb4} /* (11, 26, 26) {real, imag} */,
  {32'h3ebe8b58, 32'hbe0959b0} /* (11, 26, 25) {real, imag} */,
  {32'h3f89d005, 32'h3f0b0858} /* (11, 26, 24) {real, imag} */,
  {32'hbee664bc, 32'h3ee8b401} /* (11, 26, 23) {real, imag} */,
  {32'hbf60eed8, 32'hbf2aa017} /* (11, 26, 22) {real, imag} */,
  {32'h3e927f4a, 32'hbb94c300} /* (11, 26, 21) {real, imag} */,
  {32'hbf803992, 32'h3fbdde43} /* (11, 26, 20) {real, imag} */,
  {32'hbf393fa7, 32'h3f30feac} /* (11, 26, 19) {real, imag} */,
  {32'hbeab8cd8, 32'h3f1362e2} /* (11, 26, 18) {real, imag} */,
  {32'hbf5f2076, 32'h3f7b7786} /* (11, 26, 17) {real, imag} */,
  {32'h3e3e40c8, 32'hbde9ccb0} /* (11, 26, 16) {real, imag} */,
  {32'h3ec58c1c, 32'h3f232f8f} /* (11, 26, 15) {real, imag} */,
  {32'hbf4057c5, 32'h3e6efac8} /* (11, 26, 14) {real, imag} */,
  {32'hbf77ee08, 32'h3f589418} /* (11, 26, 13) {real, imag} */,
  {32'h3d9fd970, 32'h3f96ef60} /* (11, 26, 12) {real, imag} */,
  {32'h3d7cf100, 32'h3f30a2d2} /* (11, 26, 11) {real, imag} */,
  {32'h3c83bbac, 32'hbf15bf5d} /* (11, 26, 10) {real, imag} */,
  {32'h3fc00e23, 32'hbf83800c} /* (11, 26, 9) {real, imag} */,
  {32'h3f0155b6, 32'h3e21dcc0} /* (11, 26, 8) {real, imag} */,
  {32'hbe312e13, 32'hbe427ff4} /* (11, 26, 7) {real, imag} */,
  {32'h3f84890a, 32'hbf70ff14} /* (11, 26, 6) {real, imag} */,
  {32'h3f0c6992, 32'h3ea41468} /* (11, 26, 5) {real, imag} */,
  {32'h3f3f4550, 32'h3fab62db} /* (11, 26, 4) {real, imag} */,
  {32'h3f551129, 32'hbf0cbd06} /* (11, 26, 3) {real, imag} */,
  {32'h3f179328, 32'hbf54fe7c} /* (11, 26, 2) {real, imag} */,
  {32'h3f905488, 32'hbe0e9db4} /* (11, 26, 1) {real, imag} */,
  {32'h3ee04ef4, 32'hbee4fe28} /* (11, 26, 0) {real, imag} */,
  {32'h3f1345e9, 32'hbf46bf10} /* (11, 25, 31) {real, imag} */,
  {32'h3f5adc6f, 32'hbfd7345c} /* (11, 25, 30) {real, imag} */,
  {32'h3f3a4a47, 32'hbf676a74} /* (11, 25, 29) {real, imag} */,
  {32'h3f60c138, 32'hbe8ba794} /* (11, 25, 28) {real, imag} */,
  {32'h3e77bfd8, 32'h3f350b3a} /* (11, 25, 27) {real, imag} */,
  {32'h3cb9cd80, 32'h3f228160} /* (11, 25, 26) {real, imag} */,
  {32'h3f4bd0a0, 32'h3e87275c} /* (11, 25, 25) {real, imag} */,
  {32'h3fd10f49, 32'hbe54bea0} /* (11, 25, 24) {real, imag} */,
  {32'h3f70e3cc, 32'hbe9e2150} /* (11, 25, 23) {real, imag} */,
  {32'h3eb1f56c, 32'hbf06313a} /* (11, 25, 22) {real, imag} */,
  {32'h3e81515a, 32'h3da20670} /* (11, 25, 21) {real, imag} */,
  {32'hbecbc510, 32'h3f132394} /* (11, 25, 20) {real, imag} */,
  {32'h3f1e9691, 32'hbf99a2ff} /* (11, 25, 19) {real, imag} */,
  {32'hbf152d2c, 32'hbf08de1e} /* (11, 25, 18) {real, imag} */,
  {32'hbf844669, 32'h3e788528} /* (11, 25, 17) {real, imag} */,
  {32'h3abf2800, 32'h3ea09b26} /* (11, 25, 16) {real, imag} */,
  {32'hbe81803c, 32'h3f3a3170} /* (11, 25, 15) {real, imag} */,
  {32'h3ec57fb4, 32'h3fa5d3da} /* (11, 25, 14) {real, imag} */,
  {32'hbe8c2b34, 32'h3f8fa748} /* (11, 25, 13) {real, imag} */,
  {32'h3f842e48, 32'h3f5c9dca} /* (11, 25, 12) {real, imag} */,
  {32'hbede9610, 32'h3f99d17e} /* (11, 25, 11) {real, imag} */,
  {32'h3c061e40, 32'hbef0b660} /* (11, 25, 10) {real, imag} */,
  {32'h3f9f0067, 32'hbec4add0} /* (11, 25, 9) {real, imag} */,
  {32'hbdb17690, 32'hbe570120} /* (11, 25, 8) {real, imag} */,
  {32'hbf06fcb0, 32'hbdd34b60} /* (11, 25, 7) {real, imag} */,
  {32'h3f2e605e, 32'hbfc8c380} /* (11, 25, 6) {real, imag} */,
  {32'h3ecb9f1c, 32'h3f8598c9} /* (11, 25, 5) {real, imag} */,
  {32'h3f8851fc, 32'h40127ca1} /* (11, 25, 4) {real, imag} */,
  {32'h3f4639b6, 32'hbd8b9df0} /* (11, 25, 3) {real, imag} */,
  {32'h3f9a02d4, 32'hbfcd7f15} /* (11, 25, 2) {real, imag} */,
  {32'h401fbd90, 32'hbe4aa3e0} /* (11, 25, 1) {real, imag} */,
  {32'h3f91523e, 32'hbd2599f0} /* (11, 25, 0) {real, imag} */,
  {32'h3fa67ca4, 32'hbf132782} /* (11, 24, 31) {real, imag} */,
  {32'h3f97dda3, 32'hbfb6c9d8} /* (11, 24, 30) {real, imag} */,
  {32'h3e9c15e4, 32'hbfbb6601} /* (11, 24, 29) {real, imag} */,
  {32'hbf58dab4, 32'hbd1473c0} /* (11, 24, 28) {real, imag} */,
  {32'h3e215d60, 32'hbec83870} /* (11, 24, 27) {real, imag} */,
  {32'h3f126848, 32'hbe325c10} /* (11, 24, 26) {real, imag} */,
  {32'h3faeadb4, 32'hbd24d880} /* (11, 24, 25) {real, imag} */,
  {32'h4000bc82, 32'h3f02c9c0} /* (11, 24, 24) {real, imag} */,
  {32'h3fc45684, 32'hbf7c32e8} /* (11, 24, 23) {real, imag} */,
  {32'h3e8c4bf0, 32'hbfa0cf5b} /* (11, 24, 22) {real, imag} */,
  {32'hbf1a5884, 32'hbe84ac00} /* (11, 24, 21) {real, imag} */,
  {32'hbf65bb9a, 32'h3eff481e} /* (11, 24, 20) {real, imag} */,
  {32'hbfd36352, 32'hbf91f7fa} /* (11, 24, 19) {real, imag} */,
  {32'hbfec64ec, 32'hbfbc0e1e} /* (11, 24, 18) {real, imag} */,
  {32'hbf8dbd60, 32'hbef0ce1e} /* (11, 24, 17) {real, imag} */,
  {32'hbf762ecc, 32'h3e5ae55a} /* (11, 24, 16) {real, imag} */,
  {32'hbf7304f4, 32'h3e23f730} /* (11, 24, 15) {real, imag} */,
  {32'h3f8a83ae, 32'h3d55c8c0} /* (11, 24, 14) {real, imag} */,
  {32'h401189fa, 32'h3d4d3d00} /* (11, 24, 13) {real, imag} */,
  {32'h3f59fbc4, 32'h3edfbb34} /* (11, 24, 12) {real, imag} */,
  {32'hbeee1d70, 32'h3fbaafac} /* (11, 24, 11) {real, imag} */,
  {32'h3fd8014c, 32'h3ec1ca27} /* (11, 24, 10) {real, imag} */,
  {32'h3fd0bcad, 32'hbe982ca8} /* (11, 24, 9) {real, imag} */,
  {32'h3f2dcc4e, 32'hbf1c3590} /* (11, 24, 8) {real, imag} */,
  {32'h3dd78430, 32'hbe877564} /* (11, 24, 7) {real, imag} */,
  {32'h3e6983e0, 32'hbf8c7cdb} /* (11, 24, 6) {real, imag} */,
  {32'h3f9c7e87, 32'hbdb3c388} /* (11, 24, 5) {real, imag} */,
  {32'h3f3532d2, 32'h3f3c5b6c} /* (11, 24, 4) {real, imag} */,
  {32'h3e3ec69e, 32'hbe4c5560} /* (11, 24, 3) {real, imag} */,
  {32'h3f82b2a4, 32'hbfd0d5b0} /* (11, 24, 2) {real, imag} */,
  {32'h3fe53c14, 32'hbecc4d20} /* (11, 24, 1) {real, imag} */,
  {32'h3ed787c1, 32'hbf5397b0} /* (11, 24, 0) {real, imag} */,
  {32'h3faceb92, 32'hbdd6e47c} /* (11, 23, 31) {real, imag} */,
  {32'h3f96fbd0, 32'h3e2d1998} /* (11, 23, 30) {real, imag} */,
  {32'h3f6210ea, 32'hbf86b4e5} /* (11, 23, 29) {real, imag} */,
  {32'hbf50b56c, 32'hbf14fa88} /* (11, 23, 28) {real, imag} */,
  {32'hbe8b0030, 32'hbf2564c4} /* (11, 23, 27) {real, imag} */,
  {32'h3eaa2f50, 32'hbb76e600} /* (11, 23, 26) {real, imag} */,
  {32'h3f71a21c, 32'hbf5e0862} /* (11, 23, 25) {real, imag} */,
  {32'h3fda666c, 32'hbdf7a4e0} /* (11, 23, 24) {real, imag} */,
  {32'h40577841, 32'hbfc74540} /* (11, 23, 23) {real, imag} */,
  {32'h3fcead30, 32'hbfca1793} /* (11, 23, 22) {real, imag} */,
  {32'hbe2f6c49, 32'hbf056cb5} /* (11, 23, 21) {real, imag} */,
  {32'hbf432e30, 32'hbea58eef} /* (11, 23, 20) {real, imag} */,
  {32'hbfadaba9, 32'h3ea814c4} /* (11, 23, 19) {real, imag} */,
  {32'hc02a972e, 32'h3e1579b8} /* (11, 23, 18) {real, imag} */,
  {32'hbffd8d35, 32'h3e3de3c0} /* (11, 23, 17) {real, imag} */,
  {32'hbfa5e570, 32'hbeb528f4} /* (11, 23, 16) {real, imag} */,
  {32'hbe2a3dac, 32'h3e9e9f68} /* (11, 23, 15) {real, imag} */,
  {32'h3eecef58, 32'h3f119960} /* (11, 23, 14) {real, imag} */,
  {32'h3fd6c2fc, 32'h3e9f30dc} /* (11, 23, 13) {real, imag} */,
  {32'h3f5171d6, 32'h3e29b8c8} /* (11, 23, 12) {real, imag} */,
  {32'h3e405b54, 32'h3f206f68} /* (11, 23, 11) {real, imag} */,
  {32'h3fbd29d4, 32'h3e15dee8} /* (11, 23, 10) {real, imag} */,
  {32'h3f52745b, 32'hbc59fd80} /* (11, 23, 9) {real, imag} */,
  {32'h3f79acfe, 32'hbf0fe7d8} /* (11, 23, 8) {real, imag} */,
  {32'hbd03d110, 32'hbf16067c} /* (11, 23, 7) {real, imag} */,
  {32'h3e282d78, 32'hbfd0bcc7} /* (11, 23, 6) {real, imag} */,
  {32'h3f9a61f8, 32'hbfa05566} /* (11, 23, 5) {real, imag} */,
  {32'h3e133410, 32'hbf8a9c5d} /* (11, 23, 4) {real, imag} */,
  {32'hbf6b79f8, 32'hbeaafdce} /* (11, 23, 3) {real, imag} */,
  {32'h3def7f78, 32'hbf36e522} /* (11, 23, 2) {real, imag} */,
  {32'h3fcb5515, 32'hbe0567d4} /* (11, 23, 1) {real, imag} */,
  {32'h3ec325a4, 32'hbf178316} /* (11, 23, 0) {real, imag} */,
  {32'h3fcce4fc, 32'hbea65964} /* (11, 22, 31) {real, imag} */,
  {32'h3fb3b8eb, 32'hbdb27870} /* (11, 22, 30) {real, imag} */,
  {32'h3fb99459, 32'h3e433a50} /* (11, 22, 29) {real, imag} */,
  {32'h3f47dd66, 32'hbe23ab40} /* (11, 22, 28) {real, imag} */,
  {32'h3e03a4f0, 32'h3e3f2cb8} /* (11, 22, 27) {real, imag} */,
  {32'h3f587cb8, 32'hbdcf7f90} /* (11, 22, 26) {real, imag} */,
  {32'h3fd9bfa0, 32'hbfa7e778} /* (11, 22, 25) {real, imag} */,
  {32'h3ffba29d, 32'hbeaa0d8c} /* (11, 22, 24) {real, imag} */,
  {32'h40496b06, 32'h3e89d508} /* (11, 22, 23) {real, imag} */,
  {32'h3fe626fc, 32'hbeb668d8} /* (11, 22, 22) {real, imag} */,
  {32'h3f6100fe, 32'hbed2ceb1} /* (11, 22, 21) {real, imag} */,
  {32'hbfc820eb, 32'hbe02863e} /* (11, 22, 20) {real, imag} */,
  {32'hbefbcc00, 32'h3ea8287c} /* (11, 22, 19) {real, imag} */,
  {32'hbf91b451, 32'h3f9c3dd4} /* (11, 22, 18) {real, imag} */,
  {32'hbfc6cdf2, 32'h3f4b0ee4} /* (11, 22, 17) {real, imag} */,
  {32'hbf559ef5, 32'h3d4d3110} /* (11, 22, 16) {real, imag} */,
  {32'hbeafd4db, 32'h3eb6f1de} /* (11, 22, 15) {real, imag} */,
  {32'hbd9d9170, 32'h3f30615e} /* (11, 22, 14) {real, imag} */,
  {32'h3e4e3b06, 32'h3f9d2450} /* (11, 22, 13) {real, imag} */,
  {32'h3e1112b0, 32'h3fdab089} /* (11, 22, 12) {real, imag} */,
  {32'hbdfc4c90, 32'h3fbe3186} /* (11, 22, 11) {real, imag} */,
  {32'h3fdf5e94, 32'h3e000220} /* (11, 22, 10) {real, imag} */,
  {32'h400297f8, 32'hbf6a45c0} /* (11, 22, 9) {real, imag} */,
  {32'h400dadfc, 32'hbf30bf58} /* (11, 22, 8) {real, imag} */,
  {32'h3f86a564, 32'hbf6d24a4} /* (11, 22, 7) {real, imag} */,
  {32'h3fdcdc31, 32'hbf982c68} /* (11, 22, 6) {real, imag} */,
  {32'h3f6a74ac, 32'hbf881b12} /* (11, 22, 5) {real, imag} */,
  {32'hbe7fda14, 32'hbf75398b} /* (11, 22, 4) {real, imag} */,
  {32'h3ea17e86, 32'hbf3c8fc1} /* (11, 22, 3) {real, imag} */,
  {32'h3f7dee7a, 32'hbf7384be} /* (11, 22, 2) {real, imag} */,
  {32'h40114c2a, 32'h3f4e87c2} /* (11, 22, 1) {real, imag} */,
  {32'h3f9a4f77, 32'hbcc41c40} /* (11, 22, 0) {real, imag} */,
  {32'h3f87a975, 32'hbeaffae1} /* (11, 21, 31) {real, imag} */,
  {32'h3f1cdc3c, 32'hbf2638f2} /* (11, 21, 30) {real, imag} */,
  {32'h3ee8a174, 32'h3efcb194} /* (11, 21, 29) {real, imag} */,
  {32'h3de38ff8, 32'h3ce070e0} /* (11, 21, 28) {real, imag} */,
  {32'hbe247b88, 32'hbfda1dd5} /* (11, 21, 27) {real, imag} */,
  {32'h3fa02c6d, 32'hbfb37248} /* (11, 21, 26) {real, imag} */,
  {32'h4002c543, 32'hbf650d20} /* (11, 21, 25) {real, imag} */,
  {32'h3f8d6338, 32'h3dc6cb00} /* (11, 21, 24) {real, imag} */,
  {32'h3e1f1f16, 32'h3db6bb00} /* (11, 21, 23) {real, imag} */,
  {32'h3e9b892c, 32'hbe6af7d0} /* (11, 21, 22) {real, imag} */,
  {32'h3f09145a, 32'h3ebb2c14} /* (11, 21, 21) {real, imag} */,
  {32'hbfec933a, 32'h3fcc17bd} /* (11, 21, 20) {real, imag} */,
  {32'hbf771f16, 32'h3e4af56c} /* (11, 21, 19) {real, imag} */,
  {32'h3f864db0, 32'hbc0c4480} /* (11, 21, 18) {real, imag} */,
  {32'h3dd67f78, 32'h3f35fec7} /* (11, 21, 17) {real, imag} */,
  {32'hbea5794a, 32'h3f031de4} /* (11, 21, 16) {real, imag} */,
  {32'hbfa2c641, 32'h3f290b54} /* (11, 21, 15) {real, imag} */,
  {32'hbee44bf6, 32'h3ea13b1c} /* (11, 21, 14) {real, imag} */,
  {32'hbf01a914, 32'h3f2ba7e2} /* (11, 21, 13) {real, imag} */,
  {32'hbe8fb300, 32'h3fef6acc} /* (11, 21, 12) {real, imag} */,
  {32'h3c422c00, 32'h3fc7560e} /* (11, 21, 11) {real, imag} */,
  {32'h3f92a70f, 32'hbf11c620} /* (11, 21, 10) {real, imag} */,
  {32'h3f92bdeb, 32'hbffdfb8b} /* (11, 21, 9) {real, imag} */,
  {32'h4009f972, 32'hbfc1ca5a} /* (11, 21, 8) {real, imag} */,
  {32'h4027874a, 32'hbfb63e4c} /* (11, 21, 7) {real, imag} */,
  {32'h40260421, 32'hbe33d2e4} /* (11, 21, 6) {real, imag} */,
  {32'h3f579d6c, 32'h3e221064} /* (11, 21, 5) {real, imag} */,
  {32'hbf225a50, 32'hbde0bf2a} /* (11, 21, 4) {real, imag} */,
  {32'h3eab3164, 32'h3eaeb784} /* (11, 21, 3) {real, imag} */,
  {32'h3f6acf72, 32'hbfc2d853} /* (11, 21, 2) {real, imag} */,
  {32'h3f2aeb52, 32'h3e1eec0c} /* (11, 21, 1) {real, imag} */,
  {32'h3e0f08ba, 32'hbe6a23bc} /* (11, 21, 0) {real, imag} */,
  {32'hbe3d2fa0, 32'h3e68a498} /* (11, 20, 31) {real, imag} */,
  {32'hbeccb75c, 32'h3ef9f412} /* (11, 20, 30) {real, imag} */,
  {32'hbf8d4813, 32'h3eff7d5c} /* (11, 20, 29) {real, imag} */,
  {32'hbfd4f8f6, 32'h3f7e41f2} /* (11, 20, 28) {real, imag} */,
  {32'hbf9bb97f, 32'hbe7d5388} /* (11, 20, 27) {real, imag} */,
  {32'h3e633c54, 32'hbf7ff91d} /* (11, 20, 26) {real, imag} */,
  {32'h3f2e7214, 32'hbeb697dc} /* (11, 20, 25) {real, imag} */,
  {32'h3e652620, 32'h3f151a8c} /* (11, 20, 24) {real, imag} */,
  {32'hbeb34504, 32'h3f295c14} /* (11, 20, 23) {real, imag} */,
  {32'hbeb4bd10, 32'h3f90c010} /* (11, 20, 22) {real, imag} */,
  {32'h3df3cc84, 32'h3fa82d5b} /* (11, 20, 21) {real, imag} */,
  {32'hbec00b28, 32'h3f935d4a} /* (11, 20, 20) {real, imag} */,
  {32'hbf02c086, 32'h3e792f84} /* (11, 20, 19) {real, imag} */,
  {32'h3f49d97e, 32'h3f025e36} /* (11, 20, 18) {real, imag} */,
  {32'h3f89fbd8, 32'h3f255695} /* (11, 20, 17) {real, imag} */,
  {32'h3f8c2ed4, 32'h3e854c58} /* (11, 20, 16) {real, imag} */,
  {32'h3d863370, 32'h3edbbef1} /* (11, 20, 15) {real, imag} */,
  {32'hbf07bd2a, 32'hbf1e693f} /* (11, 20, 14) {real, imag} */,
  {32'h3e97ad82, 32'h3df868b0} /* (11, 20, 13) {real, imag} */,
  {32'h3f7e3011, 32'h3e839078} /* (11, 20, 12) {real, imag} */,
  {32'h3e03a6d0, 32'h3f9392df} /* (11, 20, 11) {real, imag} */,
  {32'hbf9ab332, 32'h3f44c651} /* (11, 20, 10) {real, imag} */,
  {32'hbf7d448e, 32'hbdec78e0} /* (11, 20, 9) {real, imag} */,
  {32'h3fc2077c, 32'hbf8a5c74} /* (11, 20, 8) {real, imag} */,
  {32'h3fdc42e7, 32'hbf09e57a} /* (11, 20, 7) {real, imag} */,
  {32'h3eca8a57, 32'h3fbe8e4a} /* (11, 20, 6) {real, imag} */,
  {32'hbefe5790, 32'h3f2ea9dc} /* (11, 20, 5) {real, imag} */,
  {32'hbf2be5b4, 32'hbef929ea} /* (11, 20, 4) {real, imag} */,
  {32'hbf81f476, 32'h3e410d00} /* (11, 20, 3) {real, imag} */,
  {32'hbf520ee7, 32'hbfca6e4e} /* (11, 20, 2) {real, imag} */,
  {32'hbf25a020, 32'h3ebdf39c} /* (11, 20, 1) {real, imag} */,
  {32'hbea53689, 32'h3f007b18} /* (11, 20, 0) {real, imag} */,
  {32'hbe98f63c, 32'h3ed34a0a} /* (11, 19, 31) {real, imag} */,
  {32'h3f2ddc9a, 32'h3ea70f42} /* (11, 19, 30) {real, imag} */,
  {32'h3da28068, 32'h3d36f894} /* (11, 19, 29) {real, imag} */,
  {32'hbf6eeb01, 32'h3fa17bc6} /* (11, 19, 28) {real, imag} */,
  {32'hbfdd8c2e, 32'h3fac05de} /* (11, 19, 27) {real, imag} */,
  {32'hbf3fb6af, 32'hbf26df76} /* (11, 19, 26) {real, imag} */,
  {32'h3e7b4180, 32'hbf2ed360} /* (11, 19, 25) {real, imag} */,
  {32'h3e7d42d0, 32'h3f7e5b4c} /* (11, 19, 24) {real, imag} */,
  {32'hbdde0000, 32'h3ffb7dd3} /* (11, 19, 23) {real, imag} */,
  {32'hbfc76b1e, 32'h3fd55635} /* (11, 19, 22) {real, imag} */,
  {32'hbe2f4171, 32'h3f6d20be} /* (11, 19, 21) {real, imag} */,
  {32'h3fa9dcc6, 32'h3fa55872} /* (11, 19, 20) {real, imag} */,
  {32'h3f5e6c93, 32'h3f16b110} /* (11, 19, 19) {real, imag} */,
  {32'hbde6b380, 32'hbeb9ed74} /* (11, 19, 18) {real, imag} */,
  {32'h3e15a990, 32'h3c22ba80} /* (11, 19, 17) {real, imag} */,
  {32'h3fcf9ab5, 32'hbf3b2bfe} /* (11, 19, 16) {real, imag} */,
  {32'h3f4b3c7e, 32'hbf5ae05f} /* (11, 19, 15) {real, imag} */,
  {32'hbd5f4e40, 32'hbfadf1dd} /* (11, 19, 14) {real, imag} */,
  {32'h3f69a2ae, 32'h3ddf1830} /* (11, 19, 13) {real, imag} */,
  {32'h3f96861a, 32'hbd0f5d70} /* (11, 19, 12) {real, imag} */,
  {32'hbf048e9f, 32'hbcf22d00} /* (11, 19, 11) {real, imag} */,
  {32'hbff1e4a0, 32'h3f3ca662} /* (11, 19, 10) {real, imag} */,
  {32'hbf721c4b, 32'h3da27cb0} /* (11, 19, 9) {real, imag} */,
  {32'h3f948024, 32'hbf349fec} /* (11, 19, 8) {real, imag} */,
  {32'h3dcb03a8, 32'hbf414a98} /* (11, 19, 7) {real, imag} */,
  {32'hbeff4a78, 32'hbdc69330} /* (11, 19, 6) {real, imag} */,
  {32'hbf139da8, 32'h3efc6b3c} /* (11, 19, 5) {real, imag} */,
  {32'hbf9cf210, 32'h3e9c3104} /* (11, 19, 4) {real, imag} */,
  {32'hbf536c88, 32'hbf7e425a} /* (11, 19, 3) {real, imag} */,
  {32'h3d824e58, 32'hbef5fc54} /* (11, 19, 2) {real, imag} */,
  {32'h3e296cbc, 32'h3f4d2fc5} /* (11, 19, 1) {real, imag} */,
  {32'hbe34658e, 32'h3e773000} /* (11, 19, 0) {real, imag} */,
  {32'hbf856abc, 32'hbed2c5e4} /* (11, 18, 31) {real, imag} */,
  {32'h3f2f4212, 32'hbd7c9f20} /* (11, 18, 30) {real, imag} */,
  {32'h3f96073e, 32'h3f5a6c24} /* (11, 18, 29) {real, imag} */,
  {32'hbe281a50, 32'h3fa578d1} /* (11, 18, 28) {real, imag} */,
  {32'hbfc5ae56, 32'h3f60f0d3} /* (11, 18, 27) {real, imag} */,
  {32'hbf9ce98d, 32'hbeb481f6} /* (11, 18, 26) {real, imag} */,
  {32'hbf96a18c, 32'hbf2a339a} /* (11, 18, 25) {real, imag} */,
  {32'hbf0842bc, 32'h3ef18428} /* (11, 18, 24) {real, imag} */,
  {32'hbefa8e44, 32'hbef6db44} /* (11, 18, 23) {real, imag} */,
  {32'hbee340f4, 32'hbf0d01c6} /* (11, 18, 22) {real, imag} */,
  {32'h3ed16321, 32'h3ec62ca2} /* (11, 18, 21) {real, imag} */,
  {32'h3f4a77bc, 32'h3f88f8fa} /* (11, 18, 20) {real, imag} */,
  {32'h3f7b6948, 32'h3e637398} /* (11, 18, 19) {real, imag} */,
  {32'h3f72f084, 32'hbfb7960b} /* (11, 18, 18) {real, imag} */,
  {32'h3f62bf52, 32'hbff40bed} /* (11, 18, 17) {real, imag} */,
  {32'h3ff08a62, 32'hbfdf19be} /* (11, 18, 16) {real, imag} */,
  {32'h3f88e78f, 32'hbedf5f04} /* (11, 18, 15) {real, imag} */,
  {32'hbe3ca1c8, 32'hbf4df9d2} /* (11, 18, 14) {real, imag} */,
  {32'hbe6a7300, 32'hbec1d110} /* (11, 18, 13) {real, imag} */,
  {32'hbf749346, 32'hbf88a311} /* (11, 18, 12) {real, imag} */,
  {32'hbfbf05e2, 32'hc008358a} /* (11, 18, 11) {real, imag} */,
  {32'hbf9fae80, 32'h3eeba364} /* (11, 18, 10) {real, imag} */,
  {32'hbfa92baa, 32'h3ffc7b46} /* (11, 18, 9) {real, imag} */,
  {32'h3f9c0c71, 32'h3fc6d94b} /* (11, 18, 8) {real, imag} */,
  {32'h3ed97740, 32'h3f0e7028} /* (11, 18, 7) {real, imag} */,
  {32'h3e5f4510, 32'h3f0ae552} /* (11, 18, 6) {real, imag} */,
  {32'h3f49259c, 32'h3f68c160} /* (11, 18, 5) {real, imag} */,
  {32'hbec1ac70, 32'h3f6b64c8} /* (11, 18, 4) {real, imag} */,
  {32'hbda42be4, 32'h3dda7600} /* (11, 18, 3) {real, imag} */,
  {32'h3e3d6b88, 32'h3e8171c5} /* (11, 18, 2) {real, imag} */,
  {32'h3ee56060, 32'hbdd423c0} /* (11, 18, 1) {real, imag} */,
  {32'hbf4d54d9, 32'hbeb44cea} /* (11, 18, 0) {real, imag} */,
  {32'hbf0d3cfc, 32'h3b662e00} /* (11, 17, 31) {real, imag} */,
  {32'hbda74fa0, 32'h3e3fc0c0} /* (11, 17, 30) {real, imag} */,
  {32'h3e95e070, 32'h3f942c86} /* (11, 17, 29) {real, imag} */,
  {32'hbf964bb6, 32'h3f37f33c} /* (11, 17, 28) {real, imag} */,
  {32'hbfc5f6c6, 32'hbeb6e7f6} /* (11, 17, 27) {real, imag} */,
  {32'hbf3db134, 32'hbe428d44} /* (11, 17, 26) {real, imag} */,
  {32'hbfb10616, 32'h3f514990} /* (11, 17, 25) {real, imag} */,
  {32'hbf7a8e4a, 32'h3fbc9b65} /* (11, 17, 24) {real, imag} */,
  {32'hbf918d48, 32'hbf89c57a} /* (11, 17, 23) {real, imag} */,
  {32'hbf825daa, 32'h3d363180} /* (11, 17, 22) {real, imag} */,
  {32'hbf6ec854, 32'h3f0ea081} /* (11, 17, 21) {real, imag} */,
  {32'hbea57d38, 32'h3f693a45} /* (11, 17, 20) {real, imag} */,
  {32'h3f39448e, 32'h3d9ded00} /* (11, 17, 19) {real, imag} */,
  {32'h3f70e8b0, 32'hbfb9e099} /* (11, 17, 18) {real, imag} */,
  {32'h3fddddec, 32'hc027eba7} /* (11, 17, 17) {real, imag} */,
  {32'h3ff96320, 32'hbfcaad4d} /* (11, 17, 16) {real, imag} */,
  {32'h3f7d6c94, 32'hbf01f028} /* (11, 17, 15) {real, imag} */,
  {32'h3deaa4a0, 32'h3c854f00} /* (11, 17, 14) {real, imag} */,
  {32'h3e89fb38, 32'hbec826c2} /* (11, 17, 13) {real, imag} */,
  {32'hbe68d928, 32'hbf88afea} /* (11, 17, 12) {real, imag} */,
  {32'hbfb91304, 32'hbfcd681e} /* (11, 17, 11) {real, imag} */,
  {32'hbf8e3142, 32'h3f8df2bc} /* (11, 17, 10) {real, imag} */,
  {32'hbf20365c, 32'h402c1fd8} /* (11, 17, 9) {real, imag} */,
  {32'hbeece6d8, 32'h40212367} /* (11, 17, 8) {real, imag} */,
  {32'hbf311fc6, 32'h3fd5ec2e} /* (11, 17, 7) {real, imag} */,
  {32'hbed77a6c, 32'h3f8b1134} /* (11, 17, 6) {real, imag} */,
  {32'hbede22c0, 32'hbde123a0} /* (11, 17, 5) {real, imag} */,
  {32'hbf22c7fe, 32'hbe10afd8} /* (11, 17, 4) {real, imag} */,
  {32'hbee84ffe, 32'hbf041b60} /* (11, 17, 3) {real, imag} */,
  {32'hbd8fcd8c, 32'hbe0b9d28} /* (11, 17, 2) {real, imag} */,
  {32'h3f4ad2b0, 32'hbf8406d3} /* (11, 17, 1) {real, imag} */,
  {32'hbe92991f, 32'hbf0441ac} /* (11, 17, 0) {real, imag} */,
  {32'hbf0d6fe9, 32'h3f1898ac} /* (11, 16, 31) {real, imag} */,
  {32'h3e1d7a68, 32'hbe548450} /* (11, 16, 30) {real, imag} */,
  {32'h3ed1f346, 32'h3ef21ad8} /* (11, 16, 29) {real, imag} */,
  {32'hbf64c1bc, 32'h3f60e366} /* (11, 16, 28) {real, imag} */,
  {32'hbf8d153d, 32'h3eaef7cc} /* (11, 16, 27) {real, imag} */,
  {32'hbf3cb7c1, 32'h3f9389a6} /* (11, 16, 26) {real, imag} */,
  {32'hbf3efc54, 32'h402e4d47} /* (11, 16, 25) {real, imag} */,
  {32'hbf02d75a, 32'h40141596} /* (11, 16, 24) {real, imag} */,
  {32'hbf784cbe, 32'h3ee8c208} /* (11, 16, 23) {real, imag} */,
  {32'hbfcbc7f0, 32'h3f31c594} /* (11, 16, 22) {real, imag} */,
  {32'hbfa610a2, 32'hbf6af25f} /* (11, 16, 21) {real, imag} */,
  {32'h3dfd0260, 32'h3ebe5210} /* (11, 16, 20) {real, imag} */,
  {32'h3f98f3a8, 32'hbee62812} /* (11, 16, 19) {real, imag} */,
  {32'h3f98b995, 32'hbfb9ad9d} /* (11, 16, 18) {real, imag} */,
  {32'hbd7df000, 32'hbfc1a1d6} /* (11, 16, 17) {real, imag} */,
  {32'h3f62e052, 32'hbf73a18c} /* (11, 16, 16) {real, imag} */,
  {32'h3f8e7631, 32'h3e2400a8} /* (11, 16, 15) {real, imag} */,
  {32'h3f207e92, 32'h3fa9ad4a} /* (11, 16, 14) {real, imag} */,
  {32'hbf510c45, 32'h3ebd20d6} /* (11, 16, 13) {real, imag} */,
  {32'hbef3d4c0, 32'hbd85a410} /* (11, 16, 12) {real, imag} */,
  {32'hbe1d2248, 32'hbe2cfba8} /* (11, 16, 11) {real, imag} */,
  {32'h3d1dbf00, 32'h3f8f5342} /* (11, 16, 10) {real, imag} */,
  {32'h3f7d788f, 32'h3f65ba8a} /* (11, 16, 9) {real, imag} */,
  {32'hbfa14451, 32'h3db11420} /* (11, 16, 8) {real, imag} */,
  {32'hc01e778b, 32'h3f2c0ac4} /* (11, 16, 7) {real, imag} */,
  {32'hbfa5b085, 32'h3fd39097} /* (11, 16, 6) {real, imag} */,
  {32'hbeee9fc0, 32'h3d7d8b60} /* (11, 16, 5) {real, imag} */,
  {32'hbf92e0f4, 32'hbec34e50} /* (11, 16, 4) {real, imag} */,
  {32'hbffb7b56, 32'hbe34c3f0} /* (11, 16, 3) {real, imag} */,
  {32'hbea107b4, 32'hbea8f010} /* (11, 16, 2) {real, imag} */,
  {32'h3ef3e7a0, 32'hbf6fcb1e} /* (11, 16, 1) {real, imag} */,
  {32'h3e0cff70, 32'hbd8bd618} /* (11, 16, 0) {real, imag} */,
  {32'h3c158880, 32'h3f177831} /* (11, 15, 31) {real, imag} */,
  {32'hbf46104e, 32'hbfa3ba6c} /* (11, 15, 30) {real, imag} */,
  {32'hbebe1d3c, 32'hbf1d7a14} /* (11, 15, 29) {real, imag} */,
  {32'hbfa15958, 32'h3fb65358} /* (11, 15, 28) {real, imag} */,
  {32'hbf5df988, 32'h3fbe860b} /* (11, 15, 27) {real, imag} */,
  {32'hbf1139fb, 32'h3f947115} /* (11, 15, 26) {real, imag} */,
  {32'hbfc18f78, 32'h3fb673f4} /* (11, 15, 25) {real, imag} */,
  {32'hbf838953, 32'h3f9c5d1e} /* (11, 15, 24) {real, imag} */,
  {32'hbf5f99f0, 32'hbed87068} /* (11, 15, 23) {real, imag} */,
  {32'hbf9630ab, 32'h3e8cd9a8} /* (11, 15, 22) {real, imag} */,
  {32'hbead98c4, 32'hbdad42d0} /* (11, 15, 21) {real, imag} */,
  {32'h3f1c0a89, 32'h3e062958} /* (11, 15, 20) {real, imag} */,
  {32'h3f78ce7c, 32'hbf9b9bf2} /* (11, 15, 19) {real, imag} */,
  {32'h3c5ac7d0, 32'hbff5f50a} /* (11, 15, 18) {real, imag} */,
  {32'hbf37e48e, 32'hbfd24357} /* (11, 15, 17) {real, imag} */,
  {32'h3f9c13dc, 32'hbf219e0e} /* (11, 15, 16) {real, imag} */,
  {32'h3fb7a58d, 32'h3f1a911a} /* (11, 15, 15) {real, imag} */,
  {32'h3fc9dca6, 32'h3fa0507b} /* (11, 15, 14) {real, imag} */,
  {32'hbee42f16, 32'h3e787f30} /* (11, 15, 13) {real, imag} */,
  {32'hbfd88eac, 32'h3e5bbf20} /* (11, 15, 12) {real, imag} */,
  {32'hbf0be7f4, 32'h3e8b6670} /* (11, 15, 11) {real, imag} */,
  {32'hbf33727c, 32'h3f62f3d8} /* (11, 15, 10) {real, imag} */,
  {32'hbe5ad368, 32'h3fe39af7} /* (11, 15, 9) {real, imag} */,
  {32'hbfea583c, 32'h3f024444} /* (11, 15, 8) {real, imag} */,
  {32'hc0323e1e, 32'hbf3552f4} /* (11, 15, 7) {real, imag} */,
  {32'hbf83e326, 32'h3deb1360} /* (11, 15, 6) {real, imag} */,
  {32'h3ec0c8fe, 32'h3eb31a56} /* (11, 15, 5) {real, imag} */,
  {32'h3e602a0c, 32'h3dad7dc4} /* (11, 15, 4) {real, imag} */,
  {32'hbf066974, 32'h3e6756a0} /* (11, 15, 3) {real, imag} */,
  {32'h3d219cc0, 32'hbd161900} /* (11, 15, 2) {real, imag} */,
  {32'h3f4ddd04, 32'hbf44922a} /* (11, 15, 1) {real, imag} */,
  {32'h3ec1635c, 32'hbe8fb5f4} /* (11, 15, 0) {real, imag} */,
  {32'hbfb1886b, 32'h3df80438} /* (11, 14, 31) {real, imag} */,
  {32'hc0380748, 32'hbf218ab8} /* (11, 14, 30) {real, imag} */,
  {32'hc01193fe, 32'h3e05b7f8} /* (11, 14, 29) {real, imag} */,
  {32'hbfe6d475, 32'h3fd57cf0} /* (11, 14, 28) {real, imag} */,
  {32'hc011826c, 32'h3f990d8d} /* (11, 14, 27) {real, imag} */,
  {32'hc013834e, 32'h3e6f87d8} /* (11, 14, 26) {real, imag} */,
  {32'hc02547f4, 32'h3f72ca48} /* (11, 14, 25) {real, imag} */,
  {32'hbfd6f038, 32'h3fa68e3c} /* (11, 14, 24) {real, imag} */,
  {32'hbfcd1bd4, 32'h3ef2f0c8} /* (11, 14, 23) {real, imag} */,
  {32'hc00bc0aa, 32'hbf31e754} /* (11, 14, 22) {real, imag} */,
  {32'hbf291a0e, 32'hbf441b05} /* (11, 14, 21) {real, imag} */,
  {32'h3faac95c, 32'hbf459824} /* (11, 14, 20) {real, imag} */,
  {32'h3eda13c4, 32'hbf48998d} /* (11, 14, 19) {real, imag} */,
  {32'hbd557220, 32'hbf318294} /* (11, 14, 18) {real, imag} */,
  {32'h3f2551e9, 32'hbdbd2270} /* (11, 14, 17) {real, imag} */,
  {32'h3faf45c2, 32'hbf178480} /* (11, 14, 16) {real, imag} */,
  {32'h3fd5590c, 32'h3d191ef0} /* (11, 14, 15) {real, imag} */,
  {32'h4012e6cc, 32'hbe34aca0} /* (11, 14, 14) {real, imag} */,
  {32'h3fda6de5, 32'hbe3d78e8} /* (11, 14, 13) {real, imag} */,
  {32'h3f233a4c, 32'h3ef4407c} /* (11, 14, 12) {real, imag} */,
  {32'h3f751832, 32'h3f2dc0a8} /* (11, 14, 11) {real, imag} */,
  {32'hbf895d4c, 32'h3fcc6c8c} /* (11, 14, 10) {real, imag} */,
  {32'hbf4158e8, 32'h400a81ec} /* (11, 14, 9) {real, imag} */,
  {32'hbe5af508, 32'h3f6f336c} /* (11, 14, 8) {real, imag} */,
  {32'hbfd5ba59, 32'h3f3a5b52} /* (11, 14, 7) {real, imag} */,
  {32'hbfaa876c, 32'h3bfc8980} /* (11, 14, 6) {real, imag} */,
  {32'h3e72f188, 32'hbf24f264} /* (11, 14, 5) {real, imag} */,
  {32'h3f777d5d, 32'hbd823008} /* (11, 14, 4) {real, imag} */,
  {32'h3e36c180, 32'hbde96a80} /* (11, 14, 3) {real, imag} */,
  {32'hbdded1b0, 32'hbf6eebdf} /* (11, 14, 2) {real, imag} */,
  {32'h3faa8ec1, 32'hbf9261b0} /* (11, 14, 1) {real, imag} */,
  {32'h3f1f631c, 32'hbf0a168b} /* (11, 14, 0) {real, imag} */,
  {32'hbfb86ee9, 32'h3f0f93ca} /* (11, 13, 31) {real, imag} */,
  {32'hc038ad5a, 32'h3f29ca1d} /* (11, 13, 30) {real, imag} */,
  {32'hc0115d06, 32'h3ff9d01a} /* (11, 13, 29) {real, imag} */,
  {32'hc0156a74, 32'h400549b8} /* (11, 13, 28) {real, imag} */,
  {32'hbfeeafca, 32'h3f211466} /* (11, 13, 27) {real, imag} */,
  {32'hbfdc6ceb, 32'hbe801f68} /* (11, 13, 26) {real, imag} */,
  {32'hc021db20, 32'h3f712a18} /* (11, 13, 25) {real, imag} */,
  {32'hc006ae8e, 32'h3feb63b8} /* (11, 13, 24) {real, imag} */,
  {32'hbfa44994, 32'h400bc588} /* (11, 13, 23) {real, imag} */,
  {32'hc004219e, 32'h3fa8ca05} /* (11, 13, 22) {real, imag} */,
  {32'hbff47825, 32'h3f4c7755} /* (11, 13, 21) {real, imag} */,
  {32'h3fcd35b9, 32'h3f2807e4} /* (11, 13, 20) {real, imag} */,
  {32'h3fb73bf3, 32'h3fa260e0} /* (11, 13, 19) {real, imag} */,
  {32'h3fe3c7d5, 32'h3f0d0790} /* (11, 13, 18) {real, imag} */,
  {32'h3fccfd1e, 32'h3ec1bf20} /* (11, 13, 17) {real, imag} */,
  {32'h3fa90e94, 32'h3c8784f0} /* (11, 13, 16) {real, imag} */,
  {32'h3efc97b4, 32'h3e63385c} /* (11, 13, 15) {real, imag} */,
  {32'h3f694f62, 32'hbf2d4b8e} /* (11, 13, 14) {real, imag} */,
  {32'h3fea5e68, 32'hbe8e0e48} /* (11, 13, 13) {real, imag} */,
  {32'h3fd2fea1, 32'h3f236023} /* (11, 13, 12) {real, imag} */,
  {32'h3f79e9dd, 32'h3f6c7158} /* (11, 13, 11) {real, imag} */,
  {32'hc00685ee, 32'h3fe76258} /* (11, 13, 10) {real, imag} */,
  {32'hbf0b2a1a, 32'h40131e60} /* (11, 13, 9) {real, imag} */,
  {32'hbc253e00, 32'h3f23647d} /* (11, 13, 8) {real, imag} */,
  {32'hbf990f62, 32'h3fc752a0} /* (11, 13, 7) {real, imag} */,
  {32'hbf8b3d00, 32'h3f347b1f} /* (11, 13, 6) {real, imag} */,
  {32'hbd50b5f8, 32'hbe06fb40} /* (11, 13, 5) {real, imag} */,
  {32'hbe155564, 32'h3f8fa79f} /* (11, 13, 4) {real, imag} */,
  {32'hbfa0a71a, 32'h3ea300b0} /* (11, 13, 3) {real, imag} */,
  {32'hbf9ba868, 32'hbfa6f1be} /* (11, 13, 2) {real, imag} */,
  {32'h3f6caf40, 32'hbfd45193} /* (11, 13, 1) {real, imag} */,
  {32'h3e8ab4a7, 32'hbe908e80} /* (11, 13, 0) {real, imag} */,
  {32'hbde5bbac, 32'h3fd88ec4} /* (11, 12, 31) {real, imag} */,
  {32'hbeb6883a, 32'h3fc5ca9a} /* (11, 12, 30) {real, imag} */,
  {32'hbeefc2d0, 32'h3fed7ade} /* (11, 12, 29) {real, imag} */,
  {32'hbf98aba6, 32'h3f9925b1} /* (11, 12, 28) {real, imag} */,
  {32'hbfeb10c7, 32'hbe2435f8} /* (11, 12, 27) {real, imag} */,
  {32'hbf05f9a2, 32'hbec806a0} /* (11, 12, 26) {real, imag} */,
  {32'hbf95b6d0, 32'h3fe6acbd} /* (11, 12, 25) {real, imag} */,
  {32'hbff6ff1a, 32'h3eeeba4e} /* (11, 12, 24) {real, imag} */,
  {32'hbff6b3d5, 32'h3eb30988} /* (11, 12, 23) {real, imag} */,
  {32'hbf72f062, 32'h3f5c0230} /* (11, 12, 22) {real, imag} */,
  {32'hbfbaa88e, 32'h3f3f4c28} /* (11, 12, 21) {real, imag} */,
  {32'h3f5f3b68, 32'h3ebee290} /* (11, 12, 20) {real, imag} */,
  {32'h401c42ec, 32'h3ec55f10} /* (11, 12, 19) {real, imag} */,
  {32'h4025713e, 32'h3f418192} /* (11, 12, 18) {real, imag} */,
  {32'h40100a27, 32'h3f234bde} /* (11, 12, 17) {real, imag} */,
  {32'h3f465d78, 32'h3e1730b0} /* (11, 12, 16) {real, imag} */,
  {32'h3e47dd00, 32'h3e114488} /* (11, 12, 15) {real, imag} */,
  {32'h3f67603b, 32'hbedb81b6} /* (11, 12, 14) {real, imag} */,
  {32'h3f9bb39e, 32'hbea2433a} /* (11, 12, 13) {real, imag} */,
  {32'h4003bbb8, 32'hbf186410} /* (11, 12, 12) {real, imag} */,
  {32'hbe3bb8e0, 32'hbe541998} /* (11, 12, 11) {real, imag} */,
  {32'hbfefb90c, 32'h3e479bc0} /* (11, 12, 10) {real, imag} */,
  {32'hbef5562c, 32'h3f9b2d6e} /* (11, 12, 9) {real, imag} */,
  {32'hbf311c82, 32'h3f53dd53} /* (11, 12, 8) {real, imag} */,
  {32'hbf001bf2, 32'h3f8918d5} /* (11, 12, 7) {real, imag} */,
  {32'hbf85b482, 32'h3f24ba66} /* (11, 12, 6) {real, imag} */,
  {32'hbf48a028, 32'h3ed62622} /* (11, 12, 5) {real, imag} */,
  {32'hbeeffaf8, 32'h3f297765} /* (11, 12, 4) {real, imag} */,
  {32'hbf82b2de, 32'h3f7d8d5a} /* (11, 12, 3) {real, imag} */,
  {32'hc004ea22, 32'h3f155e4a} /* (11, 12, 2) {real, imag} */,
  {32'hbf3203b2, 32'hbf726f0c} /* (11, 12, 1) {real, imag} */,
  {32'h3e974e87, 32'h3d4f4230} /* (11, 12, 0) {real, imag} */,
  {32'h3ec52b9c, 32'h3e618014} /* (11, 11, 31) {real, imag} */,
  {32'h3ea41945, 32'h3e63ca98} /* (11, 11, 30) {real, imag} */,
  {32'h3e03a688, 32'h3f32db32} /* (11, 11, 29) {real, imag} */,
  {32'h3d67b940, 32'h3f7b9d8c} /* (11, 11, 28) {real, imag} */,
  {32'hbe6cbecc, 32'h3e72af94} /* (11, 11, 27) {real, imag} */,
  {32'hbeac55f4, 32'hbf2a7384} /* (11, 11, 26) {real, imag} */,
  {32'h3ec78a85, 32'h3f5cf492} /* (11, 11, 25) {real, imag} */,
  {32'hbf3bd5cc, 32'hbf8acf31} /* (11, 11, 24) {real, imag} */,
  {32'hc00786f4, 32'hbeda7928} /* (11, 11, 23) {real, imag} */,
  {32'hbf6c96de, 32'h3e727764} /* (11, 11, 22) {real, imag} */,
  {32'hbf23ef2c, 32'h3ecc63e6} /* (11, 11, 21) {real, imag} */,
  {32'h3e82a7fc, 32'hbed63aba} /* (11, 11, 20) {real, imag} */,
  {32'h3e6b21fc, 32'hbf669d8e} /* (11, 11, 19) {real, imag} */,
  {32'h3f655732, 32'hbf6c5654} /* (11, 11, 18) {real, imag} */,
  {32'h3f2e9ae6, 32'hbebbfe90} /* (11, 11, 17) {real, imag} */,
  {32'hbedacf3b, 32'hbcbc5460} /* (11, 11, 16) {real, imag} */,
  {32'hbcae1520, 32'hbeaa81f8} /* (11, 11, 15) {real, imag} */,
  {32'h3f713ea8, 32'hbf8430f4} /* (11, 11, 14) {real, imag} */,
  {32'h3f93f519, 32'hbf8ef65c} /* (11, 11, 13) {real, imag} */,
  {32'h3f1ba632, 32'hbfa5cb5a} /* (11, 11, 12) {real, imag} */,
  {32'hbf6aff44, 32'hbf91cf73} /* (11, 11, 11) {real, imag} */,
  {32'hbf4aed3e, 32'hbcceede0} /* (11, 11, 10) {real, imag} */,
  {32'hbeab75d0, 32'h3ff876e6} /* (11, 11, 9) {real, imag} */,
  {32'hbff54d2d, 32'h3fdb949e} /* (11, 11, 8) {real, imag} */,
  {32'hbfd025b7, 32'hbeb96640} /* (11, 11, 7) {real, imag} */,
  {32'hbf441204, 32'hbff78d7d} /* (11, 11, 6) {real, imag} */,
  {32'hbf2fd878, 32'hbf9eb0b0} /* (11, 11, 5) {real, imag} */,
  {32'hbf411828, 32'h3f156bd0} /* (11, 11, 4) {real, imag} */,
  {32'hbf0d46be, 32'h3f58c49e} /* (11, 11, 3) {real, imag} */,
  {32'hbf4c422b, 32'hbf09331a} /* (11, 11, 2) {real, imag} */,
  {32'hbf9f2d5e, 32'h3e86cb60} /* (11, 11, 1) {real, imag} */,
  {32'hbf141088, 32'h3f1cded5} /* (11, 11, 0) {real, imag} */,
  {32'h3da3d280, 32'hbf4f4be5} /* (11, 10, 31) {real, imag} */,
  {32'h3e76cd70, 32'hbeb16642} /* (11, 10, 30) {real, imag} */,
  {32'h3fced138, 32'h3d6fef80} /* (11, 10, 29) {real, imag} */,
  {32'h4011b2ee, 32'h3eb4d7fa} /* (11, 10, 28) {real, imag} */,
  {32'h402bdc70, 32'h3f996d7e} /* (11, 10, 27) {real, imag} */,
  {32'h3fa56595, 32'hbe9dbd93} /* (11, 10, 26) {real, imag} */,
  {32'h3fdd44a4, 32'h3dbb1960} /* (11, 10, 25) {real, imag} */,
  {32'h3ed9a810, 32'h3ef66f28} /* (11, 10, 24) {real, imag} */,
  {32'hbf73dcae, 32'h3fd91044} /* (11, 10, 23) {real, imag} */,
  {32'hbee7daca, 32'h3f4d2f1c} /* (11, 10, 22) {real, imag} */,
  {32'h3da6bc70, 32'h3f4cdf89} /* (11, 10, 21) {real, imag} */,
  {32'hbf4447da, 32'h3ea13ca4} /* (11, 10, 20) {real, imag} */,
  {32'hc004bc0c, 32'h3e0c0500} /* (11, 10, 19) {real, imag} */,
  {32'hbfa13742, 32'hbf7bb4a4} /* (11, 10, 18) {real, imag} */,
  {32'hbf86d956, 32'hbef1f93e} /* (11, 10, 17) {real, imag} */,
  {32'h3e717dc2, 32'h3fb1987e} /* (11, 10, 16) {real, imag} */,
  {32'hbf08724b, 32'h3f0d4d54} /* (11, 10, 15) {real, imag} */,
  {32'h3db126e4, 32'hbf88587a} /* (11, 10, 14) {real, imag} */,
  {32'h3e5ca94e, 32'hbf5cbcfe} /* (11, 10, 13) {real, imag} */,
  {32'hbd0ab5b4, 32'hbe934a1c} /* (11, 10, 12) {real, imag} */,
  {32'hbf30fc48, 32'h3f2de48c} /* (11, 10, 11) {real, imag} */,
  {32'hbf999ee0, 32'h3fac39fb} /* (11, 10, 10) {real, imag} */,
  {32'hbe9bf5a8, 32'h4000ede3} /* (11, 10, 9) {real, imag} */,
  {32'hbf93194e, 32'h3fa53168} /* (11, 10, 8) {real, imag} */,
  {32'hbfb690fe, 32'hbf3226f8} /* (11, 10, 7) {real, imag} */,
  {32'hbf4c3f97, 32'hc053f624} /* (11, 10, 6) {real, imag} */,
  {32'h3c26c000, 32'hc0333dc2} /* (11, 10, 5) {real, imag} */,
  {32'h3f00aa70, 32'hbd5eed50} /* (11, 10, 4) {real, imag} */,
  {32'h3ce508a0, 32'hbe065060} /* (11, 10, 3) {real, imag} */,
  {32'h3eddfa84, 32'hc005383f} /* (11, 10, 2) {real, imag} */,
  {32'h3fbf0f12, 32'hbf64decf} /* (11, 10, 1) {real, imag} */,
  {32'h3fa2abc6, 32'hbecf4f48} /* (11, 10, 0) {real, imag} */,
  {32'h3e9494ae, 32'hbfaf200a} /* (11, 9, 31) {real, imag} */,
  {32'h3fe0e293, 32'hbf475e06} /* (11, 9, 30) {real, imag} */,
  {32'h4020f3b4, 32'h3f84c8b9} /* (11, 9, 29) {real, imag} */,
  {32'h3fedd5c6, 32'h3d154c60} /* (11, 9, 28) {real, imag} */,
  {32'h40076847, 32'h3e237a58} /* (11, 9, 27) {real, imag} */,
  {32'h3fb83da0, 32'h3f03e707} /* (11, 9, 26) {real, imag} */,
  {32'h3eb61aba, 32'h3ec8dd70} /* (11, 9, 25) {real, imag} */,
  {32'h3ee3a084, 32'h3f3f20be} /* (11, 9, 24) {real, imag} */,
  {32'h3fc31b69, 32'h3fa5e4b2} /* (11, 9, 23) {real, imag} */,
  {32'h3e132280, 32'hbf11bee6} /* (11, 9, 22) {real, imag} */,
  {32'hbd2b1f40, 32'hbeb619e8} /* (11, 9, 21) {real, imag} */,
  {32'hbfdbc11c, 32'h3f1b69c8} /* (11, 9, 20) {real, imag} */,
  {32'hbfc5491e, 32'h3ebd0c98} /* (11, 9, 19) {real, imag} */,
  {32'hbf790226, 32'hbebc4c68} /* (11, 9, 18) {real, imag} */,
  {32'hbf5a672c, 32'h3e95b440} /* (11, 9, 17) {real, imag} */,
  {32'hbd2245a0, 32'h3fc3bae3} /* (11, 9, 16) {real, imag} */,
  {32'hc0038232, 32'h3fcb5464} /* (11, 9, 15) {real, imag} */,
  {32'hbf679ce6, 32'h3e9c85f0} /* (11, 9, 14) {real, imag} */,
  {32'hbf6a4016, 32'hbe41d300} /* (11, 9, 13) {real, imag} */,
  {32'hbef418e2, 32'hbe557368} /* (11, 9, 12) {real, imag} */,
  {32'hbf73e5ea, 32'h3f0ec174} /* (11, 9, 11) {real, imag} */,
  {32'hbfacaecc, 32'h3f8a67cc} /* (11, 9, 10) {real, imag} */,
  {32'hbf83cf46, 32'h3fe7bf9a} /* (11, 9, 9) {real, imag} */,
  {32'hbf8a9a40, 32'h3faefe3c} /* (11, 9, 8) {real, imag} */,
  {32'hbf11f570, 32'h3f1a90ae} /* (11, 9, 7) {real, imag} */,
  {32'h3ec62096, 32'hbf8eafd8} /* (11, 9, 6) {real, imag} */,
  {32'h3edb198a, 32'hbfcdc4ee} /* (11, 9, 5) {real, imag} */,
  {32'h3f8350eb, 32'h3f024aba} /* (11, 9, 4) {real, imag} */,
  {32'h3f87df4f, 32'hbe9bc164} /* (11, 9, 3) {real, imag} */,
  {32'h3fbfe1df, 32'hbe1e89a0} /* (11, 9, 2) {real, imag} */,
  {32'h3fbbac79, 32'hbeef18e8} /* (11, 9, 1) {real, imag} */,
  {32'h3f614b2c, 32'hbf524e04} /* (11, 9, 0) {real, imag} */,
  {32'h3ee56df0, 32'hbf444a1e} /* (11, 8, 31) {real, imag} */,
  {32'h40112784, 32'hbfb73de4} /* (11, 8, 30) {real, imag} */,
  {32'h3fe7ff26, 32'hbe0cdd88} /* (11, 8, 29) {real, imag} */,
  {32'hbde55568, 32'hbe61f830} /* (11, 8, 28) {real, imag} */,
  {32'hbf23a4da, 32'hbf726a63} /* (11, 8, 27) {real, imag} */,
  {32'hbef8a899, 32'hbea0f51c} /* (11, 8, 26) {real, imag} */,
  {32'h3e5dbde7, 32'h3dbed2a0} /* (11, 8, 25) {real, imag} */,
  {32'h3fce47e7, 32'hbd8eb5e0} /* (11, 8, 24) {real, imag} */,
  {32'h3fff9e99, 32'hbf24d148} /* (11, 8, 23) {real, imag} */,
  {32'h3f9a7d99, 32'hbfc5cc4b} /* (11, 8, 22) {real, imag} */,
  {32'h3f9f7b15, 32'hbfb620be} /* (11, 8, 21) {real, imag} */,
  {32'hbede5072, 32'h3f1c44bb} /* (11, 8, 20) {real, imag} */,
  {32'hbf475b76, 32'h3f81ff68} /* (11, 8, 19) {real, imag} */,
  {32'hbf39c51c, 32'h3edb7d20} /* (11, 8, 18) {real, imag} */,
  {32'hbfc86574, 32'h3e81b4f0} /* (11, 8, 17) {real, imag} */,
  {32'hbf79468e, 32'h3fc22c83} /* (11, 8, 16) {real, imag} */,
  {32'hbf9367e0, 32'h3fc83e70} /* (11, 8, 15) {real, imag} */,
  {32'hbfe07ba0, 32'h3f640966} /* (11, 8, 14) {real, imag} */,
  {32'hbf9a0a51, 32'hbd4536c0} /* (11, 8, 13) {real, imag} */,
  {32'h3f2a642e, 32'h3f56ac84} /* (11, 8, 12) {real, imag} */,
  {32'h3e7b7570, 32'h3f3bada8} /* (11, 8, 11) {real, imag} */,
  {32'h3f07edc3, 32'h3ef9df28} /* (11, 8, 10) {real, imag} */,
  {32'hbef32a74, 32'hbebe3f1c} /* (11, 8, 9) {real, imag} */,
  {32'hbf514986, 32'hbea2ad04} /* (11, 8, 8) {real, imag} */,
  {32'hbf120134, 32'hbf4314ce} /* (11, 8, 7) {real, imag} */,
  {32'h3fb7d404, 32'hbf29fa64} /* (11, 8, 6) {real, imag} */,
  {32'h3fb2280d, 32'hbf358bf4} /* (11, 8, 5) {real, imag} */,
  {32'h3f91cb16, 32'hbfcff1ed} /* (11, 8, 4) {real, imag} */,
  {32'hbdd3d230, 32'hbfb02b48} /* (11, 8, 3) {real, imag} */,
  {32'h3ed05c30, 32'h3fa0d328} /* (11, 8, 2) {real, imag} */,
  {32'h3f640465, 32'h3f0bb4f6} /* (11, 8, 1) {real, imag} */,
  {32'h3e9daadd, 32'hbf704e0c} /* (11, 8, 0) {real, imag} */,
  {32'hbe805a35, 32'hbf031c5e} /* (11, 7, 31) {real, imag} */,
  {32'h3f611200, 32'hbf91225a} /* (11, 7, 30) {real, imag} */,
  {32'h3ef5a438, 32'hbfd5443f} /* (11, 7, 29) {real, imag} */,
  {32'hbf3ff870, 32'hbfe7d074} /* (11, 7, 28) {real, imag} */,
  {32'hbf88a77a, 32'hbf2c8d32} /* (11, 7, 27) {real, imag} */,
  {32'h3d67d060, 32'h3f66bada} /* (11, 7, 26) {real, imag} */,
  {32'h3fb8ea90, 32'h3ea8f108} /* (11, 7, 25) {real, imag} */,
  {32'h3f8bf6d1, 32'hbf2c48cc} /* (11, 7, 24) {real, imag} */,
  {32'h3f051b76, 32'hbfc574f9} /* (11, 7, 23) {real, imag} */,
  {32'h3fb7f5fd, 32'hbf988ee7} /* (11, 7, 22) {real, imag} */,
  {32'h4026fbd0, 32'hbf725f17} /* (11, 7, 21) {real, imag} */,
  {32'h3fbb6894, 32'hbe101bb0} /* (11, 7, 20) {real, imag} */,
  {32'h3e9a1720, 32'h3f029746} /* (11, 7, 19) {real, imag} */,
  {32'hbf40d6e7, 32'hbe807db0} /* (11, 7, 18) {real, imag} */,
  {32'hbfbec4d2, 32'hbea2a800} /* (11, 7, 17) {real, imag} */,
  {32'hbf74d784, 32'h3e9be720} /* (11, 7, 16) {real, imag} */,
  {32'hbf695d64, 32'hbeeb9bd6} /* (11, 7, 15) {real, imag} */,
  {32'hbfd5e427, 32'hbef6827c} /* (11, 7, 14) {real, imag} */,
  {32'hc013ff91, 32'hbf396417} /* (11, 7, 13) {real, imag} */,
  {32'h3dc9e540, 32'h3f854b26} /* (11, 7, 12) {real, imag} */,
  {32'h3f275ac0, 32'h3f6e9228} /* (11, 7, 11) {real, imag} */,
  {32'h3f45169c, 32'hbed4cac9} /* (11, 7, 10) {real, imag} */,
  {32'h3e8bfe6c, 32'hbf2b2346} /* (11, 7, 9) {real, imag} */,
  {32'h3e03187c, 32'hbd936f80} /* (11, 7, 8) {real, imag} */,
  {32'hbf8d5c39, 32'hbeafa0e4} /* (11, 7, 7) {real, imag} */,
  {32'h3f0a0c51, 32'hbf0708d4} /* (11, 7, 6) {real, imag} */,
  {32'h40067bef, 32'hbf9e303b} /* (11, 7, 5) {real, imag} */,
  {32'h3fef917f, 32'hbff72593} /* (11, 7, 4) {real, imag} */,
  {32'hbf2143b4, 32'hbfa3d01f} /* (11, 7, 3) {real, imag} */,
  {32'h3f03ec70, 32'h3d237d30} /* (11, 7, 2) {real, imag} */,
  {32'h3f1a780c, 32'hbf87d910} /* (11, 7, 1) {real, imag} */,
  {32'h3eb3756e, 32'hbf366a2d} /* (11, 7, 0) {real, imag} */,
  {32'hbf294acc, 32'hbf52225a} /* (11, 6, 31) {real, imag} */,
  {32'hbcab6500, 32'hbfd500ea} /* (11, 6, 30) {real, imag} */,
  {32'h3f200d91, 32'hbfd1b04b} /* (11, 6, 29) {real, imag} */,
  {32'hbece8b06, 32'hbff1c67b} /* (11, 6, 28) {real, imag} */,
  {32'hbf8479af, 32'hbef1fff4} /* (11, 6, 27) {real, imag} */,
  {32'h3f732e72, 32'h3fd2330e} /* (11, 6, 26) {real, imag} */,
  {32'h3f48ba0e, 32'h3ea301fc} /* (11, 6, 25) {real, imag} */,
  {32'h3d922590, 32'hbfb6dd76} /* (11, 6, 24) {real, imag} */,
  {32'h3e184b4c, 32'hbf22b2b8} /* (11, 6, 23) {real, imag} */,
  {32'hbded47d8, 32'h3e2a8ca0} /* (11, 6, 22) {real, imag} */,
  {32'h3f9fec16, 32'h3dcee290} /* (11, 6, 21) {real, imag} */,
  {32'h3f547396, 32'hbf420bcb} /* (11, 6, 20) {real, imag} */,
  {32'h3ef2fef2, 32'hbf31a74e} /* (11, 6, 19) {real, imag} */,
  {32'hbf1bd37a, 32'hbfdd687a} /* (11, 6, 18) {real, imag} */,
  {32'hbf827d02, 32'hbfbd134e} /* (11, 6, 17) {real, imag} */,
  {32'hbfb5fcc0, 32'hbed53240} /* (11, 6, 16) {real, imag} */,
  {32'hbfadee94, 32'hbf8e6d5e} /* (11, 6, 15) {real, imag} */,
  {32'hbf627093, 32'hbf6ba929} /* (11, 6, 14) {real, imag} */,
  {32'hbfba142e, 32'hbfbfe378} /* (11, 6, 13) {real, imag} */,
  {32'hbf8d0920, 32'h3f44db4e} /* (11, 6, 12) {real, imag} */,
  {32'hbecd3844, 32'h3fc7209b} /* (11, 6, 11) {real, imag} */,
  {32'hbe13933c, 32'hbf435069} /* (11, 6, 10) {real, imag} */,
  {32'h3e939900, 32'hbf794726} /* (11, 6, 9) {real, imag} */,
  {32'h3ebc5e30, 32'h3f99f92b} /* (11, 6, 8) {real, imag} */,
  {32'hbedbd5bc, 32'h3f4eb41e} /* (11, 6, 7) {real, imag} */,
  {32'h3d170de0, 32'hbe9720e0} /* (11, 6, 6) {real, imag} */,
  {32'h3fb4a856, 32'hbfda3125} /* (11, 6, 5) {real, imag} */,
  {32'h3f8a7ab4, 32'hbf421754} /* (11, 6, 4) {real, imag} */,
  {32'h3dd14880, 32'h3f0a3af8} /* (11, 6, 3) {real, imag} */,
  {32'h3eff34a4, 32'h3e2bed90} /* (11, 6, 2) {real, imag} */,
  {32'h3f4f8fc8, 32'hbf724164} /* (11, 6, 1) {real, imag} */,
  {32'h3d7a7880, 32'hbedd9d54} /* (11, 6, 0) {real, imag} */,
  {32'h3ededf56, 32'hbf86b1f6} /* (11, 5, 31) {real, imag} */,
  {32'h3fa571ba, 32'hbfcb553a} /* (11, 5, 30) {real, imag} */,
  {32'h3f6082d2, 32'hbf187200} /* (11, 5, 29) {real, imag} */,
  {32'h3eab959c, 32'hbf882878} /* (11, 5, 28) {real, imag} */,
  {32'hbeb617b8, 32'hbc8bed80} /* (11, 5, 27) {real, imag} */,
  {32'h3f03f4a4, 32'h3f9327d6} /* (11, 5, 26) {real, imag} */,
  {32'h3d13a560, 32'hbf256fea} /* (11, 5, 25) {real, imag} */,
  {32'h3efd5074, 32'hbfa5546a} /* (11, 5, 24) {real, imag} */,
  {32'h3f56c8e4, 32'h3f016a76} /* (11, 5, 23) {real, imag} */,
  {32'h3f02e556, 32'h3fc1929d} /* (11, 5, 22) {real, imag} */,
  {32'h3f8c38b0, 32'h3f9ead0e} /* (11, 5, 21) {real, imag} */,
  {32'h3ec5cf84, 32'hbf34ec94} /* (11, 5, 20) {real, imag} */,
  {32'hbeae48d6, 32'h3d9bfa50} /* (11, 5, 19) {real, imag} */,
  {32'h3e7e0178, 32'hbe2d7f3c} /* (11, 5, 18) {real, imag} */,
  {32'h3ee6f485, 32'hbf235851} /* (11, 5, 17) {real, imag} */,
  {32'h3c8fbae0, 32'hbf90db24} /* (11, 5, 16) {real, imag} */,
  {32'hbfa19ec6, 32'hbf01291d} /* (11, 5, 15) {real, imag} */,
  {32'hbf82324e, 32'hbf4236fc} /* (11, 5, 14) {real, imag} */,
  {32'hbf336fe4, 32'hbfa3b10a} /* (11, 5, 13) {real, imag} */,
  {32'hc002e267, 32'h3f9b61a8} /* (11, 5, 12) {real, imag} */,
  {32'hc0204ce8, 32'h3f982d10} /* (11, 5, 11) {real, imag} */,
  {32'hbfb001d8, 32'hbfa6b5d3} /* (11, 5, 10) {real, imag} */,
  {32'hbf90e79a, 32'hbfc80771} /* (11, 5, 9) {real, imag} */,
  {32'hbf91fd65, 32'h3f5b4758} /* (11, 5, 8) {real, imag} */,
  {32'hbfa5b522, 32'h3f4402c5} /* (11, 5, 7) {real, imag} */,
  {32'hbfd1f866, 32'hbf6d09d5} /* (11, 5, 6) {real, imag} */,
  {32'hbe311958, 32'hbfdabad6} /* (11, 5, 5) {real, imag} */,
  {32'h3f8a228c, 32'hbf92bf7c} /* (11, 5, 4) {real, imag} */,
  {32'h3fdeedf9, 32'h3ef3dc8b} /* (11, 5, 3) {real, imag} */,
  {32'h3fdff17a, 32'h3e563464} /* (11, 5, 2) {real, imag} */,
  {32'h3fd5616e, 32'h3d374ea0} /* (11, 5, 1) {real, imag} */,
  {32'h3f8122f4, 32'hbe300138} /* (11, 5, 0) {real, imag} */,
  {32'h3eed1088, 32'hbfbcbda8} /* (11, 4, 31) {real, imag} */,
  {32'h3efe1460, 32'hc01b3268} /* (11, 4, 30) {real, imag} */,
  {32'h3f965bf9, 32'hbfaa137a} /* (11, 4, 29) {real, imag} */,
  {32'h3f0f997a, 32'hbf46ff1a} /* (11, 4, 28) {real, imag} */,
  {32'h3fb7cd82, 32'hbfa7fefc} /* (11, 4, 27) {real, imag} */,
  {32'h3f8e5afe, 32'hbf6fc814} /* (11, 4, 26) {real, imag} */,
  {32'h3f0fc0b8, 32'hbf2095b4} /* (11, 4, 25) {real, imag} */,
  {32'h3e35e23c, 32'hbf00e882} /* (11, 4, 24) {real, imag} */,
  {32'hbd734e10, 32'h3eb21018} /* (11, 4, 23) {real, imag} */,
  {32'hbc849420, 32'h3f6a1c08} /* (11, 4, 22) {real, imag} */,
  {32'h3fd5f3dd, 32'h3f55b920} /* (11, 4, 21) {real, imag} */,
  {32'h402a77a0, 32'h3d7553e0} /* (11, 4, 20) {real, imag} */,
  {32'h3f81e119, 32'h3f85f908} /* (11, 4, 19) {real, imag} */,
  {32'h3f9be7fc, 32'h3f034d46} /* (11, 4, 18) {real, imag} */,
  {32'h3f36c00b, 32'h3ecef42c} /* (11, 4, 17) {real, imag} */,
  {32'h3fccecdd, 32'hbd6d4180} /* (11, 4, 16) {real, imag} */,
  {32'h3daec1e4, 32'h3ed5f256} /* (11, 4, 15) {real, imag} */,
  {32'hbfcdec19, 32'h3e85d748} /* (11, 4, 14) {real, imag} */,
  {32'hbf07c152, 32'h3e095454} /* (11, 4, 13) {real, imag} */,
  {32'hbfa9cd82, 32'h3f8b5dcf} /* (11, 4, 12) {real, imag} */,
  {32'hc0083ca8, 32'h3fc19fc4} /* (11, 4, 11) {real, imag} */,
  {32'hbf8e9795, 32'h3bbe1fc0} /* (11, 4, 10) {real, imag} */,
  {32'hbfee0ccb, 32'hbeda334d} /* (11, 4, 9) {real, imag} */,
  {32'hc007a7a5, 32'h3fd2ab8b} /* (11, 4, 8) {real, imag} */,
  {32'hbfd6252a, 32'h3f9d7c30} /* (11, 4, 7) {real, imag} */,
  {32'hc020abf3, 32'h3c54b3c0} /* (11, 4, 6) {real, imag} */,
  {32'hbeb68144, 32'hbf60c67a} /* (11, 4, 5) {real, imag} */,
  {32'h401501da, 32'hbf8ffe62} /* (11, 4, 4) {real, imag} */,
  {32'h3fdc3d95, 32'h3e9539c8} /* (11, 4, 3) {real, imag} */,
  {32'h3fcf2988, 32'h3fa89bb4} /* (11, 4, 2) {real, imag} */,
  {32'h3fad65b4, 32'h3f6087bc} /* (11, 4, 1) {real, imag} */,
  {32'h3f99211d, 32'hbf0110a4} /* (11, 4, 0) {real, imag} */,
  {32'h3eb8ccac, 32'hbf028a6a} /* (11, 3, 31) {real, imag} */,
  {32'h3f029ec4, 32'hbff60055} /* (11, 3, 30) {real, imag} */,
  {32'h3f28f9d4, 32'hbfb383f2} /* (11, 3, 29) {real, imag} */,
  {32'h3ef53428, 32'hbdc32f70} /* (11, 3, 28) {real, imag} */,
  {32'h3f93f131, 32'hbf2bf704} /* (11, 3, 27) {real, imag} */,
  {32'h3ebcf694, 32'hbfc58b62} /* (11, 3, 26) {real, imag} */,
  {32'h3ead9504, 32'hbf7f52aa} /* (11, 3, 25) {real, imag} */,
  {32'hbf0c73bf, 32'hbf6357b6} /* (11, 3, 24) {real, imag} */,
  {32'h3f3cc993, 32'hbec6f95c} /* (11, 3, 23) {real, imag} */,
  {32'h3f871d0d, 32'hbe1ff580} /* (11, 3, 22) {real, imag} */,
  {32'h3ed475b6, 32'hbf58ce61} /* (11, 3, 21) {real, imag} */,
  {32'h3fc3ae62, 32'hbf873ea2} /* (11, 3, 20) {real, imag} */,
  {32'h3fc718e1, 32'h3f175fbe} /* (11, 3, 19) {real, imag} */,
  {32'h3fae6b57, 32'h3e9595e8} /* (11, 3, 18) {real, imag} */,
  {32'h3f86b62b, 32'hbddee2e0} /* (11, 3, 17) {real, imag} */,
  {32'h3fb6540d, 32'hbd8ddf60} /* (11, 3, 16) {real, imag} */,
  {32'h3fb4e27a, 32'h3f3fed0f} /* (11, 3, 15) {real, imag} */,
  {32'hbe98be80, 32'h3ebc1792} /* (11, 3, 14) {real, imag} */,
  {32'hbe035890, 32'hbf882cb6} /* (11, 3, 13) {real, imag} */,
  {32'h3e7356d2, 32'h3eb1acb0} /* (11, 3, 12) {real, imag} */,
  {32'hbec7065e, 32'h404627c4} /* (11, 3, 11) {real, imag} */,
  {32'hbf838738, 32'h3f296aab} /* (11, 3, 10) {real, imag} */,
  {32'hbfd415dd, 32'h3e914320} /* (11, 3, 9) {real, imag} */,
  {32'hbff2463c, 32'h3fc93341} /* (11, 3, 8) {real, imag} */,
  {32'hbfab509b, 32'h4007e54d} /* (11, 3, 7) {real, imag} */,
  {32'hbfd691e0, 32'hbe907502} /* (11, 3, 6) {real, imag} */,
  {32'h3f7f71ee, 32'hc00ded3a} /* (11, 3, 5) {real, imag} */,
  {32'h3fecf8ba, 32'hbff2a490} /* (11, 3, 4) {real, imag} */,
  {32'h3f3569b8, 32'hbf5a21b8} /* (11, 3, 3) {real, imag} */,
  {32'hbe084940, 32'hbec4fe68} /* (11, 3, 2) {real, imag} */,
  {32'hbd4d9d10, 32'h3bc0b300} /* (11, 3, 1) {real, imag} */,
  {32'h3e3dd004, 32'hbf6c53af} /* (11, 3, 0) {real, imag} */,
  {32'h3fc97986, 32'h3ef78db0} /* (11, 2, 31) {real, imag} */,
  {32'h400fd198, 32'hbe63ec30} /* (11, 2, 30) {real, imag} */,
  {32'h3c128400, 32'hbf93ac1f} /* (11, 2, 29) {real, imag} */,
  {32'h3f450b70, 32'hbf5e23b1} /* (11, 2, 28) {real, imag} */,
  {32'hbe9c6a00, 32'hbf020146} /* (11, 2, 27) {real, imag} */,
  {32'hbf824b40, 32'hbfaebe4b} /* (11, 2, 26) {real, imag} */,
  {32'h3f8918aa, 32'hbfabc074} /* (11, 2, 25) {real, imag} */,
  {32'h3f9eb7b7, 32'hbf519638} /* (11, 2, 24) {real, imag} */,
  {32'h3fdf6082, 32'hbe893fe0} /* (11, 2, 23) {real, imag} */,
  {32'h3f9c58fe, 32'hbf87848d} /* (11, 2, 22) {real, imag} */,
  {32'h3e4010a0, 32'hbf76ecc4} /* (11, 2, 21) {real, imag} */,
  {32'h3f0c232a, 32'hbf9d3729} /* (11, 2, 20) {real, imag} */,
  {32'h3f804a16, 32'hbf50750c} /* (11, 2, 19) {real, imag} */,
  {32'h4008bf0c, 32'hc00147e4} /* (11, 2, 18) {real, imag} */,
  {32'h4039b907, 32'hc01b020e} /* (11, 2, 17) {real, imag} */,
  {32'h3f349eae, 32'hbf66c438} /* (11, 2, 16) {real, imag} */,
  {32'h3f954adf, 32'h3f32e94c} /* (11, 2, 15) {real, imag} */,
  {32'h3f90e2b6, 32'h3f860903} /* (11, 2, 14) {real, imag} */,
  {32'hbed4eea2, 32'hbf2e1092} /* (11, 2, 13) {real, imag} */,
  {32'hbf79b15e, 32'h3e6e8810} /* (11, 2, 12) {real, imag} */,
  {32'h3e1ebbf0, 32'h402aaaa4} /* (11, 2, 11) {real, imag} */,
  {32'h3df59af0, 32'hbf1c0f43} /* (11, 2, 10) {real, imag} */,
  {32'hbf9ecdfc, 32'hbf87a40e} /* (11, 2, 9) {real, imag} */,
  {32'hbfd13872, 32'h3e7ed890} /* (11, 2, 8) {real, imag} */,
  {32'hbf4c46f7, 32'h3f10b210} /* (11, 2, 7) {real, imag} */,
  {32'hbf331587, 32'hbf7496f2} /* (11, 2, 6) {real, imag} */,
  {32'h3ea5ade2, 32'hbfdbfabb} /* (11, 2, 5) {real, imag} */,
  {32'h3fcd1ab0, 32'hbf4dfaba} /* (11, 2, 4) {real, imag} */,
  {32'h3fe72109, 32'h3b67a400} /* (11, 2, 3) {real, imag} */,
  {32'h3fb1b06d, 32'h3d6986e0} /* (11, 2, 2) {real, imag} */,
  {32'h3fa77178, 32'hbef06930} /* (11, 2, 1) {real, imag} */,
  {32'h3f158dc0, 32'hbf855308} /* (11, 2, 0) {real, imag} */,
  {32'h3f8d755a, 32'hbf267d22} /* (11, 1, 31) {real, imag} */,
  {32'h3f9322b4, 32'hbe45973c} /* (11, 1, 30) {real, imag} */,
  {32'hbf11749f, 32'h3f7bafc8} /* (11, 1, 29) {real, imag} */,
  {32'h3f0b83ec, 32'h3e9aeee4} /* (11, 1, 28) {real, imag} */,
  {32'hbee76160, 32'hbd9d3500} /* (11, 1, 27) {real, imag} */,
  {32'hbd626580, 32'hbf458ad6} /* (11, 1, 26) {real, imag} */,
  {32'h3fd3f231, 32'hbf415f5a} /* (11, 1, 25) {real, imag} */,
  {32'h4007c814, 32'h3faead02} /* (11, 1, 24) {real, imag} */,
  {32'h3fd0c93c, 32'h3f94a5d2} /* (11, 1, 23) {real, imag} */,
  {32'h3faabf9e, 32'hbf778504} /* (11, 1, 22) {real, imag} */,
  {32'h3ee6c0ec, 32'hbf073098} /* (11, 1, 21) {real, imag} */,
  {32'h3ee21bb8, 32'hbeda2350} /* (11, 1, 20) {real, imag} */,
  {32'h3ea6ecc0, 32'hbf45dcc8} /* (11, 1, 19) {real, imag} */,
  {32'h3f961c11, 32'hc0251429} /* (11, 1, 18) {real, imag} */,
  {32'h4013a26e, 32'hc0517adc} /* (11, 1, 17) {real, imag} */,
  {32'h3e9481dc, 32'hbec218b0} /* (11, 1, 16) {real, imag} */,
  {32'hbe9e9dd2, 32'h3fb6922f} /* (11, 1, 15) {real, imag} */,
  {32'hbf7f7a8a, 32'h3f8116a4} /* (11, 1, 14) {real, imag} */,
  {32'hbf716f06, 32'hbf0879be} /* (11, 1, 13) {real, imag} */,
  {32'hbef01db2, 32'h3ea805ec} /* (11, 1, 12) {real, imag} */,
  {32'h3e5da128, 32'h3fe9287a} /* (11, 1, 11) {real, imag} */,
  {32'h3e0a5f30, 32'hbdda77c0} /* (11, 1, 10) {real, imag} */,
  {32'hbf50aed4, 32'hbdec3640} /* (11, 1, 9) {real, imag} */,
  {32'hbf1cabc4, 32'h3fa6ea5c} /* (11, 1, 8) {real, imag} */,
  {32'hbe72fe08, 32'h3e4a7ed0} /* (11, 1, 7) {real, imag} */,
  {32'h3e43e4f8, 32'h3f27634e} /* (11, 1, 6) {real, imag} */,
  {32'h3e9a1cf7, 32'h3f2f5d91} /* (11, 1, 5) {real, imag} */,
  {32'h4013c52e, 32'h3d92f774} /* (11, 1, 4) {real, imag} */,
  {32'h4004c956, 32'h3f3228ef} /* (11, 1, 3) {real, imag} */,
  {32'h3f9a5ca4, 32'h3f3b5e1a} /* (11, 1, 2) {real, imag} */,
  {32'h3f41c0a2, 32'hbf99678c} /* (11, 1, 1) {real, imag} */,
  {32'h3f5812b7, 32'hbfcc6d88} /* (11, 1, 0) {real, imag} */,
  {32'h3e8ac790, 32'hbf2d71c9} /* (11, 0, 31) {real, imag} */,
  {32'h3db8a338, 32'h3df347ec} /* (11, 0, 30) {real, imag} */,
  {32'hbf4719e8, 32'h3fd36387} /* (11, 0, 29) {real, imag} */,
  {32'hbec729bc, 32'h3f592af3} /* (11, 0, 28) {real, imag} */,
  {32'hbeca1d9a, 32'h3f27f0fe} /* (11, 0, 27) {real, imag} */,
  {32'h3e0453e8, 32'hbd56d720} /* (11, 0, 26) {real, imag} */,
  {32'h3f41a332, 32'hbe28e518} /* (11, 0, 25) {real, imag} */,
  {32'h3fb196c2, 32'h3f808d29} /* (11, 0, 24) {real, imag} */,
  {32'h3fe3d1d2, 32'h3f1165c8} /* (11, 0, 23) {real, imag} */,
  {32'h3fb1b883, 32'hbec84b68} /* (11, 0, 22) {real, imag} */,
  {32'h3ebb3563, 32'hbeb6c160} /* (11, 0, 21) {real, imag} */,
  {32'h3e6fd400, 32'h3dfe8980} /* (11, 0, 20) {real, imag} */,
  {32'hbe8d1bc4, 32'h3e8edb8c} /* (11, 0, 19) {real, imag} */,
  {32'hbe781594, 32'hbf81947c} /* (11, 0, 18) {real, imag} */,
  {32'h3d7bb9e0, 32'hbf866d84} /* (11, 0, 17) {real, imag} */,
  {32'h3e1c3fb8, 32'h3efa97ea} /* (11, 0, 16) {real, imag} */,
  {32'h3e8c4c54, 32'h3f00282b} /* (11, 0, 15) {real, imag} */,
  {32'hbf1368cb, 32'h3d0ae6d0} /* (11, 0, 14) {real, imag} */,
  {32'hbf556cd3, 32'hbc1cc940} /* (11, 0, 13) {real, imag} */,
  {32'hbeff9b27, 32'h3f0c4bb0} /* (11, 0, 12) {real, imag} */,
  {32'hbec6eb97, 32'h3f0d53fd} /* (11, 0, 11) {real, imag} */,
  {32'hbeeb33b0, 32'hbc8b9340} /* (11, 0, 10) {real, imag} */,
  {32'hbec551fa, 32'hbe5395d4} /* (11, 0, 9) {real, imag} */,
  {32'h3ec9ac2f, 32'hbdd91380} /* (11, 0, 8) {real, imag} */,
  {32'hbf0ff754, 32'hbf3b389a} /* (11, 0, 7) {real, imag} */,
  {32'hbe7a0374, 32'h3e6ec70e} /* (11, 0, 6) {real, imag} */,
  {32'h3fd1eb48, 32'h3e971e4a} /* (11, 0, 5) {real, imag} */,
  {32'h40068ab7, 32'hbe6d6485} /* (11, 0, 4) {real, imag} */,
  {32'h3f99c879, 32'hbca58ca0} /* (11, 0, 3) {real, imag} */,
  {32'h3f7db2cc, 32'h3e2c34ec} /* (11, 0, 2) {real, imag} */,
  {32'h3f5e1580, 32'hbe5c2920} /* (11, 0, 1) {real, imag} */,
  {32'h3f164d6d, 32'hbeff3c86} /* (11, 0, 0) {real, imag} */,
  {32'hbe06886c, 32'hbe1b216a} /* (10, 31, 31) {real, imag} */,
  {32'h3ef93112, 32'hbc886a00} /* (10, 31, 30) {real, imag} */,
  {32'hbe99ce58, 32'hbeb05162} /* (10, 31, 29) {real, imag} */,
  {32'hbf611ba6, 32'h3e797814} /* (10, 31, 28) {real, imag} */,
  {32'hbeefa240, 32'h3e7d66ac} /* (10, 31, 27) {real, imag} */,
  {32'hbf12839c, 32'h3f741a86} /* (10, 31, 26) {real, imag} */,
  {32'hbf9c745f, 32'h3efe16ca} /* (10, 31, 25) {real, imag} */,
  {32'hbf789da6, 32'h3efa42c8} /* (10, 31, 24) {real, imag} */,
  {32'hbf847a88, 32'h3f837aa0} /* (10, 31, 23) {real, imag} */,
  {32'hbef754d4, 32'h3fa6e567} /* (10, 31, 22) {real, imag} */,
  {32'hbe505964, 32'h3f73c30c} /* (10, 31, 21) {real, imag} */,
  {32'hbe00c620, 32'h3df5bb64} /* (10, 31, 20) {real, imag} */,
  {32'hbd3bfb60, 32'hbebc4d64} /* (10, 31, 19) {real, imag} */,
  {32'h3eb273c8, 32'hbe9292dc} /* (10, 31, 18) {real, imag} */,
  {32'h3f3b357a, 32'hbf8d39cb} /* (10, 31, 17) {real, imag} */,
  {32'h3e7839fe, 32'hbe3cccfa} /* (10, 31, 16) {real, imag} */,
  {32'h3d87ec28, 32'hbe984f04} /* (10, 31, 15) {real, imag} */,
  {32'h3f339e7e, 32'hbf227036} /* (10, 31, 14) {real, imag} */,
  {32'h3f559fa2, 32'hbe352a40} /* (10, 31, 13) {real, imag} */,
  {32'h3f9d65da, 32'hbe8852ec} /* (10, 31, 12) {real, imag} */,
  {32'h3faff7df, 32'h3ee4d16d} /* (10, 31, 11) {real, imag} */,
  {32'hbe997360, 32'h3f61945e} /* (10, 31, 10) {real, imag} */,
  {32'hbe0c6520, 32'h3eb3c514} /* (10, 31, 9) {real, imag} */,
  {32'hbf0fe6c2, 32'h3f205aa8} /* (10, 31, 8) {real, imag} */,
  {32'h3ed077b4, 32'h3e801264} /* (10, 31, 7) {real, imag} */,
  {32'h3f94eb54, 32'h3ea6a28c} /* (10, 31, 6) {real, imag} */,
  {32'hbeb467c8, 32'h3f8e7ee7} /* (10, 31, 5) {real, imag} */,
  {32'hbf8cfba8, 32'h3f92d2c2} /* (10, 31, 4) {real, imag} */,
  {32'hbf0063d1, 32'h3ed0e05a} /* (10, 31, 3) {real, imag} */,
  {32'hbf50b148, 32'hbf4de2d9} /* (10, 31, 2) {real, imag} */,
  {32'hbecdad80, 32'hc01498da} /* (10, 31, 1) {real, imag} */,
  {32'hbec4eddc, 32'hbf8afc8c} /* (10, 31, 0) {real, imag} */,
  {32'h3edd3e28, 32'hbddd8a24} /* (10, 30, 31) {real, imag} */,
  {32'h3fd16a9e, 32'h3e0b0960} /* (10, 30, 30) {real, imag} */,
  {32'h3f852e3f, 32'hbde1f0b0} /* (10, 30, 29) {real, imag} */,
  {32'hbf17e49a, 32'h3f270d34} /* (10, 30, 28) {real, imag} */,
  {32'hbfb4c563, 32'h3f66e4ea} /* (10, 30, 27) {real, imag} */,
  {32'hbfc63e3c, 32'hbea858f0} /* (10, 30, 26) {real, imag} */,
  {32'hbfe88b86, 32'hbe7298f0} /* (10, 30, 25) {real, imag} */,
  {32'hc047964e, 32'h3eb09d58} /* (10, 30, 24) {real, imag} */,
  {32'hc015fb71, 32'h3f277254} /* (10, 30, 23) {real, imag} */,
  {32'h3f609d12, 32'h3fed428a} /* (10, 30, 22) {real, imag} */,
  {32'hbfa217cb, 32'h3fcacc7e} /* (10, 30, 21) {real, imag} */,
  {32'hbfe8f804, 32'h3f870119} /* (10, 30, 20) {real, imag} */,
  {32'h3e1556f4, 32'h3d3c5bc0} /* (10, 30, 19) {real, imag} */,
  {32'h3f93c5f2, 32'hbf06130e} /* (10, 30, 18) {real, imag} */,
  {32'h3f4c1956, 32'hbf9bb6fb} /* (10, 30, 17) {real, imag} */,
  {32'h3f8e0ace, 32'hbf920fb6} /* (10, 30, 16) {real, imag} */,
  {32'h3f126311, 32'hbdabb250} /* (10, 30, 15) {real, imag} */,
  {32'h3e514be0, 32'h3f4e509a} /* (10, 30, 14) {real, imag} */,
  {32'h3f688750, 32'h3fc7ef71} /* (10, 30, 13) {real, imag} */,
  {32'h3fde2d3a, 32'h3f3e63ae} /* (10, 30, 12) {real, imag} */,
  {32'h3f306906, 32'h3f1163e0} /* (10, 30, 11) {real, imag} */,
  {32'hbf614853, 32'h3f852e9c} /* (10, 30, 10) {real, imag} */,
  {32'hbf398d37, 32'h3e947534} /* (10, 30, 9) {real, imag} */,
  {32'hbfa359a4, 32'h3f76999a} /* (10, 30, 8) {real, imag} */,
  {32'hbf73ea2e, 32'h3fd144fd} /* (10, 30, 7) {real, imag} */,
  {32'h3ffb32cc, 32'h3f17b33e} /* (10, 30, 6) {real, imag} */,
  {32'hbf445854, 32'h3fbe9728} /* (10, 30, 5) {real, imag} */,
  {32'hbfeb435f, 32'h3f8b089c} /* (10, 30, 4) {real, imag} */,
  {32'hbf5889f7, 32'h3f933029} /* (10, 30, 3) {real, imag} */,
  {32'hbf1d97ac, 32'hbf7d8398} /* (10, 30, 2) {real, imag} */,
  {32'hbf24d2c3, 32'hbfee1e86} /* (10, 30, 1) {real, imag} */,
  {32'hbee37778, 32'hbe5d74f0} /* (10, 30, 0) {real, imag} */,
  {32'h3fb8809b, 32'h3ea70f8e} /* (10, 29, 31) {real, imag} */,
  {32'h401f9980, 32'h3ed61f70} /* (10, 29, 30) {real, imag} */,
  {32'h3f83a23d, 32'h3ee81044} /* (10, 29, 29) {real, imag} */,
  {32'hbfbeaab2, 32'h3f5ada36} /* (10, 29, 28) {real, imag} */,
  {32'hbf9a4190, 32'hbef575ba} /* (10, 29, 27) {real, imag} */,
  {32'h3f436938, 32'hbebfab90} /* (10, 29, 26) {real, imag} */,
  {32'hbefd67a2, 32'h3f646a3d} /* (10, 29, 25) {real, imag} */,
  {32'hc012ac41, 32'h3f95d396} /* (10, 29, 24) {real, imag} */,
  {32'hbfebf0f6, 32'h3fef190e} /* (10, 29, 23) {real, imag} */,
  {32'h3e49cabc, 32'h4045d098} /* (10, 29, 22) {real, imag} */,
  {32'hbec9adef, 32'h3f92a250} /* (10, 29, 21) {real, imag} */,
  {32'h3e73c884, 32'h3fb91b80} /* (10, 29, 20) {real, imag} */,
  {32'h3fb859f0, 32'h3f48b7da} /* (10, 29, 19) {real, imag} */,
  {32'h3fc1b03a, 32'h3f93ed11} /* (10, 29, 18) {real, imag} */,
  {32'h3f82ac2e, 32'hbece8542} /* (10, 29, 17) {real, imag} */,
  {32'h3f694858, 32'hbf9f3438} /* (10, 29, 16) {real, imag} */,
  {32'h3de68ec0, 32'hbf25f7a4} /* (10, 29, 15) {real, imag} */,
  {32'h3ee42570, 32'hbe0ddbc0} /* (10, 29, 14) {real, imag} */,
  {32'h3ec48820, 32'h3dca5100} /* (10, 29, 13) {real, imag} */,
  {32'h3fd71a6c, 32'h3f9957f5} /* (10, 29, 12) {real, imag} */,
  {32'h3fed428e, 32'h3f19ee4a} /* (10, 29, 11) {real, imag} */,
  {32'h3f6acd6a, 32'hbe382fbc} /* (10, 29, 10) {real, imag} */,
  {32'h3e34b4e8, 32'hbe7f6c28} /* (10, 29, 9) {real, imag} */,
  {32'hbf3a3f98, 32'h3fa45be1} /* (10, 29, 8) {real, imag} */,
  {32'h3e150e10, 32'h3ff4aefc} /* (10, 29, 7) {real, imag} */,
  {32'h3f9b6ad9, 32'h3f506c28} /* (10, 29, 6) {real, imag} */,
  {32'hbe937510, 32'h3f20850f} /* (10, 29, 5) {real, imag} */,
  {32'hbea9bb98, 32'h3f9415c5} /* (10, 29, 4) {real, imag} */,
  {32'hbf2268a0, 32'hbe85f264} /* (10, 29, 3) {real, imag} */,
  {32'hbfaf6f56, 32'hbfa124aa} /* (10, 29, 2) {real, imag} */,
  {32'hbfd5227e, 32'hbf7fd55b} /* (10, 29, 1) {real, imag} */,
  {32'hbe6c70ac, 32'h3e52cf34} /* (10, 29, 0) {real, imag} */,
  {32'h3f1f909e, 32'h3f4c2f68} /* (10, 28, 31) {real, imag} */,
  {32'h3e96f8cf, 32'h3f9c986d} /* (10, 28, 30) {real, imag} */,
  {32'hbee7acc0, 32'h3f1dff07} /* (10, 28, 29) {real, imag} */,
  {32'hbf275e7f, 32'hbf268ac8} /* (10, 28, 28) {real, imag} */,
  {32'hbe7690e0, 32'hbfe8ef56} /* (10, 28, 27) {real, imag} */,
  {32'hbedad990, 32'hbeea505c} /* (10, 28, 26) {real, imag} */,
  {32'hbf99627b, 32'h3f88cd2c} /* (10, 28, 25) {real, imag} */,
  {32'hbf5ba63a, 32'h3fb56748} /* (10, 28, 24) {real, imag} */,
  {32'hbf006ad8, 32'h40046836} /* (10, 28, 23) {real, imag} */,
  {32'h3f3d09b8, 32'h3fe1399f} /* (10, 28, 22) {real, imag} */,
  {32'h3f4b4cd4, 32'hbebd5aba} /* (10, 28, 21) {real, imag} */,
  {32'h4010f6da, 32'hbf516e3f} /* (10, 28, 20) {real, imag} */,
  {32'h3fcc3be0, 32'hbea04480} /* (10, 28, 19) {real, imag} */,
  {32'h3f88e23a, 32'h3ff49758} /* (10, 28, 18) {real, imag} */,
  {32'h3ed25d06, 32'h3f18335a} /* (10, 28, 17) {real, imag} */,
  {32'h3ec47426, 32'h3d582280} /* (10, 28, 16) {real, imag} */,
  {32'hbf18c8dc, 32'hbc61ed80} /* (10, 28, 15) {real, imag} */,
  {32'h3f5abc90, 32'h3e8e4aec} /* (10, 28, 14) {real, imag} */,
  {32'h3f0803e0, 32'hbe4bfae8} /* (10, 28, 13) {real, imag} */,
  {32'hbda5baf0, 32'hbf20f286} /* (10, 28, 12) {real, imag} */,
  {32'h3ca79840, 32'hbf0c25bf} /* (10, 28, 11) {real, imag} */,
  {32'h3efe5b6c, 32'h3f522319} /* (10, 28, 10) {real, imag} */,
  {32'h3db97810, 32'h3ea4c878} /* (10, 28, 9) {real, imag} */,
  {32'h3c0db6c0, 32'h3fd9640a} /* (10, 28, 8) {real, imag} */,
  {32'h404d3c63, 32'h3e5b1658} /* (10, 28, 7) {real, imag} */,
  {32'h3fa9121a, 32'hbef9716c} /* (10, 28, 6) {real, imag} */,
  {32'h3dd259c8, 32'hbefa16d0} /* (10, 28, 5) {real, imag} */,
  {32'h3ec91960, 32'h3f3c0e3c} /* (10, 28, 4) {real, imag} */,
  {32'hbea29130, 32'h3f255f8e} /* (10, 28, 3) {real, imag} */,
  {32'hbfcc0cae, 32'h3e4ac490} /* (10, 28, 2) {real, imag} */,
  {32'hbf35c139, 32'hbeeb1602} /* (10, 28, 1) {real, imag} */,
  {32'h3f98e359, 32'hbefb63a6} /* (10, 28, 0) {real, imag} */,
  {32'hbdf44ff8, 32'h3f2ef359} /* (10, 27, 31) {real, imag} */,
  {32'hbf8e84e3, 32'h403a2bdf} /* (10, 27, 30) {real, imag} */,
  {32'hbf6a909d, 32'h40067089} /* (10, 27, 29) {real, imag} */,
  {32'hbc9c1220, 32'h3ee3650c} /* (10, 27, 28) {real, imag} */,
  {32'h3fa541b4, 32'hc004ea2a} /* (10, 27, 27) {real, imag} */,
  {32'hbe6be170, 32'hbfd6d6b7} /* (10, 27, 26) {real, imag} */,
  {32'hbe153520, 32'h3da37360} /* (10, 27, 25) {real, imag} */,
  {32'h3f9ecbe6, 32'h3ebf9ae8} /* (10, 27, 24) {real, imag} */,
  {32'h3eebcf88, 32'h3f68fb2e} /* (10, 27, 23) {real, imag} */,
  {32'h3f641a3d, 32'h3f076c61} /* (10, 27, 22) {real, imag} */,
  {32'hbcf96b80, 32'h3ed971be} /* (10, 27, 21) {real, imag} */,
  {32'h3edbd4d8, 32'hbf8a585e} /* (10, 27, 20) {real, imag} */,
  {32'h3dc1b8a0, 32'hbef9e774} /* (10, 27, 19) {real, imag} */,
  {32'hbd4dd740, 32'hbe89949e} /* (10, 27, 18) {real, imag} */,
  {32'h3e990828, 32'h3e9b425c} /* (10, 27, 17) {real, imag} */,
  {32'h3e19e080, 32'hbe887a0a} /* (10, 27, 16) {real, imag} */,
  {32'h3e846b74, 32'hbf30505e} /* (10, 27, 15) {real, imag} */,
  {32'h3f72d356, 32'h3f48c316} /* (10, 27, 14) {real, imag} */,
  {32'hbed25ac4, 32'h3f15f1ac} /* (10, 27, 13) {real, imag} */,
  {32'hbf979700, 32'hbf588c10} /* (10, 27, 12) {real, imag} */,
  {32'hbd1ea500, 32'hbec36796} /* (10, 27, 11) {real, imag} */,
  {32'h3d4ea480, 32'h3f0e9e38} /* (10, 27, 10) {real, imag} */,
  {32'hbfed75c1, 32'hbf3ee720} /* (10, 27, 9) {real, imag} */,
  {32'hbf709700, 32'h3ec0bbf8} /* (10, 27, 8) {real, imag} */,
  {32'h3f843c95, 32'h3e46a438} /* (10, 27, 7) {real, imag} */,
  {32'h3f0eb9a5, 32'h3eed0f24} /* (10, 27, 6) {real, imag} */,
  {32'h3eb442f0, 32'h3e8868aa} /* (10, 27, 5) {real, imag} */,
  {32'hbf5f5a5a, 32'hbf83711a} /* (10, 27, 4) {real, imag} */,
  {32'h3f04e633, 32'hbe976c84} /* (10, 27, 3) {real, imag} */,
  {32'h3f0bbb24, 32'h3f5683a0} /* (10, 27, 2) {real, imag} */,
  {32'h3e035998, 32'h3d94ec50} /* (10, 27, 1) {real, imag} */,
  {32'h3f685101, 32'hbf1ccce7} /* (10, 27, 0) {real, imag} */,
  {32'hbecbb616, 32'h3f2b311b} /* (10, 26, 31) {real, imag} */,
  {32'hbf4a587e, 32'h3fc79628} /* (10, 26, 30) {real, imag} */,
  {32'hbebb36b6, 32'h3eec42a8} /* (10, 26, 29) {real, imag} */,
  {32'hbf8cf255, 32'h3eaee868} /* (10, 26, 28) {real, imag} */,
  {32'hbe72e107, 32'hbf505ba8} /* (10, 26, 27) {real, imag} */,
  {32'h3ebb9964, 32'h3ee9fb0c} /* (10, 26, 26) {real, imag} */,
  {32'h3f08590e, 32'hbf1f0752} /* (10, 26, 25) {real, imag} */,
  {32'h3f4e292c, 32'hbf46d9d8} /* (10, 26, 24) {real, imag} */,
  {32'hbef45232, 32'h3f77a346} /* (10, 26, 23) {real, imag} */,
  {32'hbf2d3ba2, 32'h3fc0d0a8} /* (10, 26, 22) {real, imag} */,
  {32'h3e1d99a4, 32'h3f9da56c} /* (10, 26, 21) {real, imag} */,
  {32'h3e9d2b4c, 32'hbda5c3f8} /* (10, 26, 20) {real, imag} */,
  {32'hbebcfc38, 32'hbe567608} /* (10, 26, 19) {real, imag} */,
  {32'hbc930040, 32'hbf90cb90} /* (10, 26, 18) {real, imag} */,
  {32'h3ec1da6c, 32'hbf103fe5} /* (10, 26, 17) {real, imag} */,
  {32'hbebda5b2, 32'h3d9966e8} /* (10, 26, 16) {real, imag} */,
  {32'h3fb33b76, 32'hbeeacbe0} /* (10, 26, 15) {real, imag} */,
  {32'h3f924d74, 32'h3f7055b6} /* (10, 26, 14) {real, imag} */,
  {32'h3ec9aac0, 32'h3f94a731} /* (10, 26, 13) {real, imag} */,
  {32'hbf595f28, 32'h3fb59f32} /* (10, 26, 12) {real, imag} */,
  {32'h3fc79aeb, 32'hbd4291d0} /* (10, 26, 11) {real, imag} */,
  {32'h3fc5b0a1, 32'h3f8f165d} /* (10, 26, 10) {real, imag} */,
  {32'hbf874572, 32'h3f4427ca} /* (10, 26, 9) {real, imag} */,
  {32'hbff2bd54, 32'h3f07f09e} /* (10, 26, 8) {real, imag} */,
  {32'hbf930daf, 32'hbf1667d2} /* (10, 26, 7) {real, imag} */,
  {32'hbef3bd80, 32'hbc214300} /* (10, 26, 6) {real, imag} */,
  {32'h3ee056e0, 32'hbef0b7ea} /* (10, 26, 5) {real, imag} */,
  {32'hbe8d140e, 32'hbe59d4f4} /* (10, 26, 4) {real, imag} */,
  {32'h3e4c6b44, 32'hbdf6ef30} /* (10, 26, 3) {real, imag} */,
  {32'hbf8d08c9, 32'h3ecde140} /* (10, 26, 2) {real, imag} */,
  {32'hbfe26b88, 32'h3f342e20} /* (10, 26, 1) {real, imag} */,
  {32'hbeeb8d12, 32'h3ea47bdc} /* (10, 26, 0) {real, imag} */,
  {32'h3d1e58e0, 32'h3f41d3a4} /* (10, 25, 31) {real, imag} */,
  {32'hbfa3c328, 32'h3fd49c16} /* (10, 25, 30) {real, imag} */,
  {32'hbead19b8, 32'h3ec1a88a} /* (10, 25, 29) {real, imag} */,
  {32'hbf980262, 32'h3f445d09} /* (10, 25, 28) {real, imag} */,
  {32'hbf2d106e, 32'hbf931818} /* (10, 25, 27) {real, imag} */,
  {32'h3f3166ef, 32'hbed4c310} /* (10, 25, 26) {real, imag} */,
  {32'h3f4703fc, 32'h3d3b3540} /* (10, 25, 25) {real, imag} */,
  {32'hbe4c294c, 32'hbf9462be} /* (10, 25, 24) {real, imag} */,
  {32'hbfe45471, 32'hbe269b84} /* (10, 25, 23) {real, imag} */,
  {32'hbfebfc01, 32'h3f2f9418} /* (10, 25, 22) {real, imag} */,
  {32'h3f1a9b12, 32'h3e0f0e5e} /* (10, 25, 21) {real, imag} */,
  {32'h3f7ee846, 32'hbf49ef0e} /* (10, 25, 20) {real, imag} */,
  {32'h3f1af6f0, 32'h3f3d66dc} /* (10, 25, 19) {real, imag} */,
  {32'h3f156310, 32'h3e7734f8} /* (10, 25, 18) {real, imag} */,
  {32'h3f648860, 32'h3e1784c8} /* (10, 25, 17) {real, imag} */,
  {32'h3f902d8f, 32'h3e50fac0} /* (10, 25, 16) {real, imag} */,
  {32'h3f49b838, 32'h3eb92dca} /* (10, 25, 15) {real, imag} */,
  {32'h3e92e780, 32'h40165adc} /* (10, 25, 14) {real, imag} */,
  {32'h3f8b8cf0, 32'h3f868485} /* (10, 25, 13) {real, imag} */,
  {32'h3f0d7d80, 32'h3face843} /* (10, 25, 12) {real, imag} */,
  {32'hbedf1774, 32'h3d87a890} /* (10, 25, 11) {real, imag} */,
  {32'h3e8d5029, 32'h3fa231e4} /* (10, 25, 10) {real, imag} */,
  {32'hbf223ece, 32'h3f5ac092} /* (10, 25, 9) {real, imag} */,
  {32'hbfca3bba, 32'hbf06cf34} /* (10, 25, 8) {real, imag} */,
  {32'hbf9647e7, 32'hbf30836e} /* (10, 25, 7) {real, imag} */,
  {32'hbf1ab5eb, 32'h3f5eb4c6} /* (10, 25, 6) {real, imag} */,
  {32'hbec8d0de, 32'h3f947c34} /* (10, 25, 5) {real, imag} */,
  {32'hbf0c824a, 32'h3e77ba88} /* (10, 25, 4) {real, imag} */,
  {32'hbeecac98, 32'h3e973034} /* (10, 25, 3) {real, imag} */,
  {32'hbfafe65c, 32'h3f81c7fb} /* (10, 25, 2) {real, imag} */,
  {32'hbfebd7e9, 32'h3fcc4652} /* (10, 25, 1) {real, imag} */,
  {32'h3ee0010c, 32'h3f927d66} /* (10, 25, 0) {real, imag} */,
  {32'hbf56a6da, 32'hbd1440f0} /* (10, 24, 31) {real, imag} */,
  {32'hc0164842, 32'h3fd81505} /* (10, 24, 30) {real, imag} */,
  {32'hbfc6a3df, 32'h3f405b6c} /* (10, 24, 29) {real, imag} */,
  {32'hc02252a5, 32'h3e37f718} /* (10, 24, 28) {real, imag} */,
  {32'hbfc290eb, 32'hb996b000} /* (10, 24, 27) {real, imag} */,
  {32'h3f5d9910, 32'h3e814edc} /* (10, 24, 26) {real, imag} */,
  {32'h3f1a7e4d, 32'hbec67df0} /* (10, 24, 25) {real, imag} */,
  {32'hbe17c304, 32'hbf18b7a6} /* (10, 24, 24) {real, imag} */,
  {32'hc035813a, 32'hbe9bacd0} /* (10, 24, 23) {real, imag} */,
  {32'hc0142716, 32'hbf91d10b} /* (10, 24, 22) {real, imag} */,
  {32'hbdb45368, 32'hbcd2bb20} /* (10, 24, 21) {real, imag} */,
  {32'hbe02a358, 32'hbec8f850} /* (10, 24, 20) {real, imag} */,
  {32'h3f4d0602, 32'h3f46f9d4} /* (10, 24, 19) {real, imag} */,
  {32'h3f94556f, 32'h3ff26b7a} /* (10, 24, 18) {real, imag} */,
  {32'h3f6d7993, 32'h3f261f9e} /* (10, 24, 17) {real, imag} */,
  {32'h3f0e5720, 32'hbe99953c} /* (10, 24, 16) {real, imag} */,
  {32'h3fe0568c, 32'hbf647acd} /* (10, 24, 15) {real, imag} */,
  {32'h4019dc94, 32'hbf32eb34} /* (10, 24, 14) {real, imag} */,
  {32'h3e2cbe70, 32'h3f60fdc6} /* (10, 24, 13) {real, imag} */,
  {32'h3e624310, 32'h3f9ff6cb} /* (10, 24, 12) {real, imag} */,
  {32'hbf87eec2, 32'h3dc777e8} /* (10, 24, 11) {real, imag} */,
  {32'hbe9538bc, 32'h3fa3eb7b} /* (10, 24, 10) {real, imag} */,
  {32'hbfad9db6, 32'h3efa0954} /* (10, 24, 9) {real, imag} */,
  {32'hc01131d2, 32'h3ebbbc00} /* (10, 24, 8) {real, imag} */,
  {32'hbf514009, 32'hbe5090f8} /* (10, 24, 7) {real, imag} */,
  {32'hbf81b2d6, 32'h3f6a8b62} /* (10, 24, 6) {real, imag} */,
  {32'hbfc7dc5b, 32'h3feafe0f} /* (10, 24, 5) {real, imag} */,
  {32'hbfacaa44, 32'h3e598bbc} /* (10, 24, 4) {real, imag} */,
  {32'hbf97b080, 32'hbf1e5aea} /* (10, 24, 3) {real, imag} */,
  {32'hbe6652f0, 32'hbb8a0a00} /* (10, 24, 2) {real, imag} */,
  {32'hbf58dcc8, 32'h3f46daf3} /* (10, 24, 1) {real, imag} */,
  {32'h3e50c4b0, 32'h3f3768ac} /* (10, 24, 0) {real, imag} */,
  {32'hbfa9fef4, 32'h3f4d3024} /* (10, 23, 31) {real, imag} */,
  {32'hc044c9e2, 32'h4003088d} /* (10, 23, 30) {real, imag} */,
  {32'hc00d9832, 32'h3faa8a18} /* (10, 23, 29) {real, imag} */,
  {32'hc03e48a6, 32'h3f5dfcc0} /* (10, 23, 28) {real, imag} */,
  {32'hc0091c52, 32'h3f900890} /* (10, 23, 27) {real, imag} */,
  {32'hbe3d13c8, 32'h3f5f09d2} /* (10, 23, 26) {real, imag} */,
  {32'hbea44fc4, 32'h3f014a4c} /* (10, 23, 25) {real, imag} */,
  {32'hbfa9dd9e, 32'h3f02b750} /* (10, 23, 24) {real, imag} */,
  {32'hc058cef1, 32'h3d97f7a0} /* (10, 23, 23) {real, imag} */,
  {32'hc0197bc4, 32'hc00f73ef} /* (10, 23, 22) {real, imag} */,
  {32'hbf5c72e6, 32'h3ee53b2a} /* (10, 23, 21) {real, imag} */,
  {32'hbdcede10, 32'h3f812ef9} /* (10, 23, 20) {real, imag} */,
  {32'h3f6a1d92, 32'hbe129888} /* (10, 23, 19) {real, imag} */,
  {32'h3df8c850, 32'h3f0954ba} /* (10, 23, 18) {real, imag} */,
  {32'hbee920b4, 32'h3f1a7524} /* (10, 23, 17) {real, imag} */,
  {32'h3ef4cafe, 32'hbf2d65b0} /* (10, 23, 16) {real, imag} */,
  {32'h3ff1e3f2, 32'hbfc33d4c} /* (10, 23, 15) {real, imag} */,
  {32'h400f218e, 32'hbf980fc3} /* (10, 23, 14) {real, imag} */,
  {32'h3ef9a410, 32'h3efda02c} /* (10, 23, 13) {real, imag} */,
  {32'h3e4a8be8, 32'h3e9388b4} /* (10, 23, 12) {real, imag} */,
  {32'hbf0f2367, 32'hbf6f9e20} /* (10, 23, 11) {real, imag} */,
  {32'hbfc2b7fe, 32'h3dce5e28} /* (10, 23, 10) {real, imag} */,
  {32'hc00916b0, 32'h3f8101c1} /* (10, 23, 9) {real, imag} */,
  {32'hbf2ba7ef, 32'h3f6c9157} /* (10, 23, 8) {real, imag} */,
  {32'hbe497f44, 32'hbe9b484c} /* (10, 23, 7) {real, imag} */,
  {32'hbf4dd74e, 32'hbf79c25e} /* (10, 23, 6) {real, imag} */,
  {32'hc0086b9f, 32'hbf1aaf9b} /* (10, 23, 5) {real, imag} */,
  {32'hbfce58e8, 32'hbdb856d0} /* (10, 23, 4) {real, imag} */,
  {32'hbfa6b4b4, 32'hbf707142} /* (10, 23, 3) {real, imag} */,
  {32'hbd83c350, 32'hbff98b00} /* (10, 23, 2) {real, imag} */,
  {32'h3e8dc888, 32'hbf86ce76} /* (10, 23, 1) {real, imag} */,
  {32'hbf284cca, 32'hbef92e82} /* (10, 23, 0) {real, imag} */,
  {32'h3d4c8b40, 32'h3eebd32a} /* (10, 22, 31) {real, imag} */,
  {32'hc01deb2e, 32'h3f55c2aa} /* (10, 22, 30) {real, imag} */,
  {32'hc01f5fe0, 32'h3ed91d80} /* (10, 22, 29) {real, imag} */,
  {32'hbfa99528, 32'h3f0bb888} /* (10, 22, 28) {real, imag} */,
  {32'hbf98e766, 32'hbbcd0800} /* (10, 22, 27) {real, imag} */,
  {32'hbedf92d0, 32'h3ec41320} /* (10, 22, 26) {real, imag} */,
  {32'hbebc9524, 32'h3fc484e0} /* (10, 22, 25) {real, imag} */,
  {32'hbf37255a, 32'h3fa76eb2} /* (10, 22, 24) {real, imag} */,
  {32'hbfb56d7e, 32'h3f764b54} /* (10, 22, 23) {real, imag} */,
  {32'hbf70774c, 32'hbed3af1a} /* (10, 22, 22) {real, imag} */,
  {32'hbe7dbf7c, 32'hbdad48e8} /* (10, 22, 21) {real, imag} */,
  {32'hbfa07ec0, 32'h3e948acc} /* (10, 22, 20) {real, imag} */,
  {32'hbfab0bc4, 32'hbe4c48c0} /* (10, 22, 19) {real, imag} */,
  {32'hbf14e724, 32'hbf9d6056} /* (10, 22, 18) {real, imag} */,
  {32'h3f005174, 32'hbf998bce} /* (10, 22, 17) {real, imag} */,
  {32'h3fbb75e4, 32'hbf87ef86} /* (10, 22, 16) {real, imag} */,
  {32'h3f431675, 32'hbf7d4867} /* (10, 22, 15) {real, imag} */,
  {32'h3ed310c6, 32'hbf568786} /* (10, 22, 14) {real, imag} */,
  {32'h3f507b84, 32'h3f2d7608} /* (10, 22, 13) {real, imag} */,
  {32'h3ea76366, 32'hbf73cc5d} /* (10, 22, 12) {real, imag} */,
  {32'h3ebd5f98, 32'hbfddcdd8} /* (10, 22, 11) {real, imag} */,
  {32'hbfd360d8, 32'hbe4b33c4} /* (10, 22, 10) {real, imag} */,
  {32'hc02944fd, 32'h3fa74439} /* (10, 22, 9) {real, imag} */,
  {32'hbe69a034, 32'hbeaa85fc} /* (10, 22, 8) {real, imag} */,
  {32'hbc9cde60, 32'hc00b5ecc} /* (10, 22, 7) {real, imag} */,
  {32'hbe2b7ce0, 32'hbfc4ccf0} /* (10, 22, 6) {real, imag} */,
  {32'hbf35dfa8, 32'hbfa425e8} /* (10, 22, 5) {real, imag} */,
  {32'hbf7d0e44, 32'h3f5d51fa} /* (10, 22, 4) {real, imag} */,
  {32'hbe915f04, 32'hbe33e8c0} /* (10, 22, 3) {real, imag} */,
  {32'h3e7be680, 32'hbfc2f93a} /* (10, 22, 2) {real, imag} */,
  {32'hbf2092db, 32'hbef10308} /* (10, 22, 1) {real, imag} */,
  {32'hbe3d6798, 32'hbf06718d} /* (10, 22, 0) {real, imag} */,
  {32'h3ea0735a, 32'hbf5b24b2} /* (10, 21, 31) {real, imag} */,
  {32'hbd2927a0, 32'hbf5d12e0} /* (10, 21, 30) {real, imag} */,
  {32'hbf0d99eb, 32'h3fb9ba0d} /* (10, 21, 29) {real, imag} */,
  {32'hbfbed6dc, 32'h40136fe1} /* (10, 21, 28) {real, imag} */,
  {32'hbf669370, 32'hbf11529f} /* (10, 21, 27) {real, imag} */,
  {32'hbe8233f4, 32'hbd97aac0} /* (10, 21, 26) {real, imag} */,
  {32'hbe355117, 32'h3f5f8a6d} /* (10, 21, 25) {real, imag} */,
  {32'h3f036f7a, 32'h3fd03c66} /* (10, 21, 24) {real, imag} */,
  {32'hbdac18b4, 32'h3f610e98} /* (10, 21, 23) {real, imag} */,
  {32'h3eff2ffa, 32'h3f3229fe} /* (10, 21, 22) {real, imag} */,
  {32'h3f21d382, 32'hbdba4da0} /* (10, 21, 21) {real, imag} */,
  {32'hbfc1dced, 32'h3ee37baf} /* (10, 21, 20) {real, imag} */,
  {32'hbfebc42b, 32'hbcff5860} /* (10, 21, 19) {real, imag} */,
  {32'h3dc78d88, 32'hbfe29f2b} /* (10, 21, 18) {real, imag} */,
  {32'h3fa55cbe, 32'hbf72576e} /* (10, 21, 17) {real, imag} */,
  {32'h3fc020f4, 32'hbcf0f9d8} /* (10, 21, 16) {real, imag} */,
  {32'h3e670c14, 32'hbf25d8f8} /* (10, 21, 15) {real, imag} */,
  {32'h3f83cf5e, 32'hbfd8a398} /* (10, 21, 14) {real, imag} */,
  {32'h3fa8d5bc, 32'hbdde59b8} /* (10, 21, 13) {real, imag} */,
  {32'h3ecf7090, 32'h3f10ef77} /* (10, 21, 12) {real, imag} */,
  {32'hbf3835a2, 32'hbf59c77d} /* (10, 21, 11) {real, imag} */,
  {32'hc007438e, 32'hbebff4b2} /* (10, 21, 10) {real, imag} */,
  {32'hc04303b1, 32'hc00ca805} /* (10, 21, 9) {real, imag} */,
  {32'hbf148758, 32'hbfd747cb} /* (10, 21, 8) {real, imag} */,
  {32'h3d483548, 32'hbf87d91d} /* (10, 21, 7) {real, imag} */,
  {32'hbf931908, 32'h3ec32be4} /* (10, 21, 6) {real, imag} */,
  {32'hbf36e444, 32'hbecc6198} /* (10, 21, 5) {real, imag} */,
  {32'hbeb4b103, 32'h3f60c6a6} /* (10, 21, 4) {real, imag} */,
  {32'hbfda9306, 32'hbe6ed3e6} /* (10, 21, 3) {real, imag} */,
  {32'hbe87a9b4, 32'hbf4bfad5} /* (10, 21, 2) {real, imag} */,
  {32'hbd3e3c00, 32'hbf15101d} /* (10, 21, 1) {real, imag} */,
  {32'h3f63de9a, 32'hbe4706f0} /* (10, 21, 0) {real, imag} */,
  {32'h3f26760c, 32'hc00825fb} /* (10, 20, 31) {real, imag} */,
  {32'h3fbcf81f, 32'hc06239f0} /* (10, 20, 30) {real, imag} */,
  {32'h3f8f5c59, 32'h3da13880} /* (10, 20, 29) {real, imag} */,
  {32'h3f270318, 32'h3fc569e0} /* (10, 20, 28) {real, imag} */,
  {32'h3f4393ea, 32'h3ecb6ee8} /* (10, 20, 27) {real, imag} */,
  {32'h3fa100ea, 32'hbf021576} /* (10, 20, 26) {real, imag} */,
  {32'h3fbacd9f, 32'hbf93de2a} /* (10, 20, 25) {real, imag} */,
  {32'h401764d8, 32'h3be3e900} /* (10, 20, 24) {real, imag} */,
  {32'h3f261099, 32'hbf471d95} /* (10, 20, 23) {real, imag} */,
  {32'hbe8fe1c8, 32'hbe2e2bf8} /* (10, 20, 22) {real, imag} */,
  {32'h3ee63206, 32'hbf55777c} /* (10, 20, 21) {real, imag} */,
  {32'hbf066cd8, 32'h3f44186a} /* (10, 20, 20) {real, imag} */,
  {32'hbf461fd0, 32'h3f650566} /* (10, 20, 19) {real, imag} */,
  {32'h3e5eb7bb, 32'hbf86b28a} /* (10, 20, 18) {real, imag} */,
  {32'h3f8524a3, 32'hbee61330} /* (10, 20, 17) {real, imag} */,
  {32'h3f193698, 32'h3eee5d60} /* (10, 20, 16) {real, imag} */,
  {32'h3e6f0780, 32'h3ecc7dbc} /* (10, 20, 15) {real, imag} */,
  {32'h40057b86, 32'hbf8351f8} /* (10, 20, 14) {real, imag} */,
  {32'h3db6aa80, 32'h3cf4ea60} /* (10, 20, 13) {real, imag} */,
  {32'hbfe4c767, 32'h3f824616} /* (10, 20, 12) {real, imag} */,
  {32'hbf8dc085, 32'h3e14eda8} /* (10, 20, 11) {real, imag} */,
  {32'hbfb2d6db, 32'h3e36fbc8} /* (10, 20, 10) {real, imag} */,
  {32'hbfa5b6c4, 32'hc0051850} /* (10, 20, 9) {real, imag} */,
  {32'h3f25b9b0, 32'hbf1f71b6} /* (10, 20, 8) {real, imag} */,
  {32'h3f85cc03, 32'h3f774947} /* (10, 20, 7) {real, imag} */,
  {32'hbe11c344, 32'h3f1a4a1c} /* (10, 20, 6) {real, imag} */,
  {32'hbe4c47cc, 32'hbdd76db8} /* (10, 20, 5) {real, imag} */,
  {32'h3e63e2a0, 32'h3f882a12} /* (10, 20, 4) {real, imag} */,
  {32'hbf5bf39e, 32'h3f95be26} /* (10, 20, 3) {real, imag} */,
  {32'hbf3cc69c, 32'h3f17d470} /* (10, 20, 2) {real, imag} */,
  {32'hbea9d054, 32'hbe5e1108} /* (10, 20, 1) {real, imag} */,
  {32'h3f3bf9f2, 32'h3e2a23cd} /* (10, 20, 0) {real, imag} */,
  {32'h3e54bcb0, 32'hbfa3884e} /* (10, 19, 31) {real, imag} */,
  {32'h3e602354, 32'hc0253987} /* (10, 19, 30) {real, imag} */,
  {32'hbf2a7abe, 32'hbec0d8e8} /* (10, 19, 29) {real, imag} */,
  {32'h3e8d49be, 32'h3fb9ebf2} /* (10, 19, 28) {real, imag} */,
  {32'h3fc29046, 32'h3f9ffec2} /* (10, 19, 27) {real, imag} */,
  {32'h400c2744, 32'hbd43cdd0} /* (10, 19, 26) {real, imag} */,
  {32'h3fffd988, 32'hbfa508cf} /* (10, 19, 25) {real, imag} */,
  {32'h3fabc5d6, 32'hbf498c76} /* (10, 19, 24) {real, imag} */,
  {32'hbef98cc4, 32'hc01dfbe8} /* (10, 19, 23) {real, imag} */,
  {32'hbf7fe88f, 32'hbf685756} /* (10, 19, 22) {real, imag} */,
  {32'hbe9d090e, 32'hbfce439e} /* (10, 19, 21) {real, imag} */,
  {32'hbf82a4e4, 32'hbeddac54} /* (10, 19, 20) {real, imag} */,
  {32'hbf361148, 32'h3fb03dd4} /* (10, 19, 19) {real, imag} */,
  {32'h3f1f709e, 32'h3ed4a394} /* (10, 19, 18) {real, imag} */,
  {32'h3fd7e628, 32'hbef1ed50} /* (10, 19, 17) {real, imag} */,
  {32'h3f9dbf05, 32'h3f05b5a9} /* (10, 19, 16) {real, imag} */,
  {32'hbe4cde70, 32'h3f73e6c8} /* (10, 19, 15) {real, imag} */,
  {32'h3f01247c, 32'h3f520690} /* (10, 19, 14) {real, imag} */,
  {32'hbfcbf0b6, 32'h3eb823f8} /* (10, 19, 13) {real, imag} */,
  {32'hbfd58ca0, 32'hbf9f6a7f} /* (10, 19, 12) {real, imag} */,
  {32'hbf9d2410, 32'hbf19b4b4} /* (10, 19, 11) {real, imag} */,
  {32'hbf0866cc, 32'h3e41ddd8} /* (10, 19, 10) {real, imag} */,
  {32'h3fa14502, 32'hbee31d48} /* (10, 19, 9) {real, imag} */,
  {32'h3f742874, 32'h3f8b46b8} /* (10, 19, 8) {real, imag} */,
  {32'h3fa768dd, 32'h4013b8ce} /* (10, 19, 7) {real, imag} */,
  {32'h3f0d93f8, 32'h3ec91f94} /* (10, 19, 6) {real, imag} */,
  {32'h3e53099c, 32'hbfcf70d8} /* (10, 19, 5) {real, imag} */,
  {32'h40035504, 32'hbf873217} /* (10, 19, 4) {real, imag} */,
  {32'h3fd7f02a, 32'hbe41ab50} /* (10, 19, 3) {real, imag} */,
  {32'hbf0c7f7a, 32'h3ec85fbc} /* (10, 19, 2) {real, imag} */,
  {32'hbe3909d8, 32'hbfec228a} /* (10, 19, 1) {real, imag} */,
  {32'h3f798217, 32'hc0160f61} /* (10, 19, 0) {real, imag} */,
  {32'h3f80b34a, 32'hbe8e0e64} /* (10, 18, 31) {real, imag} */,
  {32'h3f0b1b3c, 32'hbf608920} /* (10, 18, 30) {real, imag} */,
  {32'hbf89de7b, 32'hc0017357} /* (10, 18, 29) {real, imag} */,
  {32'hbf99efd5, 32'hbeb79c9e} /* (10, 18, 28) {real, imag} */,
  {32'hbe69e828, 32'h3f667f2c} /* (10, 18, 27) {real, imag} */,
  {32'h3fbc3001, 32'h3f56d31a} /* (10, 18, 26) {real, imag} */,
  {32'h3f99c23c, 32'h3f100c82} /* (10, 18, 25) {real, imag} */,
  {32'h3fad1020, 32'hbe601350} /* (10, 18, 24) {real, imag} */,
  {32'h3e99615c, 32'hc0149db0} /* (10, 18, 23) {real, imag} */,
  {32'hbf0e95d6, 32'hbfdbde1b} /* (10, 18, 22) {real, imag} */,
  {32'hbf5e73e7, 32'hc007e474} /* (10, 18, 21) {real, imag} */,
  {32'hbfd6114f, 32'h3f8bb4c0} /* (10, 18, 20) {real, imag} */,
  {32'hbf3f2f83, 32'h402055f4} /* (10, 18, 19) {real, imag} */,
  {32'hbf4cd54e, 32'h3f8c27e8} /* (10, 18, 18) {real, imag} */,
  {32'h3eb7d36c, 32'hbf7baf68} /* (10, 18, 17) {real, imag} */,
  {32'h3f59d128, 32'hbebdeb40} /* (10, 18, 16) {real, imag} */,
  {32'hbe32c8c0, 32'hbe824dc0} /* (10, 18, 15) {real, imag} */,
  {32'hbee0dea0, 32'h3f1f3416} /* (10, 18, 14) {real, imag} */,
  {32'hc02a4f98, 32'h3f8f3a8d} /* (10, 18, 13) {real, imag} */,
  {32'hc01a01cb, 32'hbf958daf} /* (10, 18, 12) {real, imag} */,
  {32'hbf9c70f9, 32'hbfec9b70} /* (10, 18, 11) {real, imag} */,
  {32'h3e41da04, 32'hc018e500} /* (10, 18, 10) {real, imag} */,
  {32'h3dea0b00, 32'hbfc84dfe} /* (10, 18, 9) {real, imag} */,
  {32'h3e7f85b0, 32'h3f389a02} /* (10, 18, 8) {real, imag} */,
  {32'h400b986a, 32'h3ff3669a} /* (10, 18, 7) {real, imag} */,
  {32'h3ffda25a, 32'h3eff5350} /* (10, 18, 6) {real, imag} */,
  {32'h3f5213ec, 32'hbf962f8e} /* (10, 18, 5) {real, imag} */,
  {32'h3fa71ed2, 32'hbf6b1f18} /* (10, 18, 4) {real, imag} */,
  {32'h3f1a97b8, 32'hbf5a881c} /* (10, 18, 3) {real, imag} */,
  {32'hbe5bc2b0, 32'hbf917d22} /* (10, 18, 2) {real, imag} */,
  {32'hbc782d00, 32'hbfd8f0ce} /* (10, 18, 1) {real, imag} */,
  {32'h3e9bbd38, 32'hc00b6d6e} /* (10, 18, 0) {real, imag} */,
  {32'h3f9496ca, 32'hbf3ab17c} /* (10, 17, 31) {real, imag} */,
  {32'h3f6f78ba, 32'hbf9a1c92} /* (10, 17, 30) {real, imag} */,
  {32'h3eb2af2a, 32'hbff15b0c} /* (10, 17, 29) {real, imag} */,
  {32'h3e5c2bd8, 32'hbff15baf} /* (10, 17, 28) {real, imag} */,
  {32'hbf0f1472, 32'hbe6a8fd0} /* (10, 17, 27) {real, imag} */,
  {32'hbd0aa270, 32'hbf940b99} /* (10, 17, 26) {real, imag} */,
  {32'h3f487e16, 32'h3c2bc080} /* (10, 17, 25) {real, imag} */,
  {32'h3f36cecc, 32'h3f57f5a0} /* (10, 17, 24) {real, imag} */,
  {32'hbda4e440, 32'hbe847d90} /* (10, 17, 23) {real, imag} */,
  {32'hbf06eb61, 32'hbdd583f8} /* (10, 17, 22) {real, imag} */,
  {32'hbfaa10d4, 32'h3f39351e} /* (10, 17, 21) {real, imag} */,
  {32'hc0279436, 32'h400665e2} /* (10, 17, 20) {real, imag} */,
  {32'hbf8f0983, 32'h3f5f3ba0} /* (10, 17, 19) {real, imag} */,
  {32'hbfbfe706, 32'hbedb4768} /* (10, 17, 18) {real, imag} */,
  {32'h3e3725e8, 32'hbf6173e2} /* (10, 17, 17) {real, imag} */,
  {32'hbea01768, 32'h3f7570b0} /* (10, 17, 16) {real, imag} */,
  {32'hbc3a9900, 32'h3f243744} /* (10, 17, 15) {real, imag} */,
  {32'hbe808634, 32'hbf559824} /* (10, 17, 14) {real, imag} */,
  {32'hbf9b05f8, 32'hbe7e7a6c} /* (10, 17, 13) {real, imag} */,
  {32'hbf129cf0, 32'hbefed450} /* (10, 17, 12) {real, imag} */,
  {32'hbf755733, 32'hbf8aff3c} /* (10, 17, 11) {real, imag} */,
  {32'h3f35054e, 32'hc00068ef} /* (10, 17, 10) {real, imag} */,
  {32'h3f382e90, 32'hc00f116d} /* (10, 17, 9) {real, imag} */,
  {32'h3f76c4a4, 32'hbf09e9b4} /* (10, 17, 8) {real, imag} */,
  {32'h3fe155cf, 32'h3f7a9d08} /* (10, 17, 7) {real, imag} */,
  {32'h3fcdcdec, 32'h3f719182} /* (10, 17, 6) {real, imag} */,
  {32'h3f92518e, 32'hbf8eaa20} /* (10, 17, 5) {real, imag} */,
  {32'h4015d934, 32'hbf418aac} /* (10, 17, 4) {real, imag} */,
  {32'h3f50a084, 32'hbd6feb00} /* (10, 17, 3) {real, imag} */,
  {32'hbf2acf60, 32'h3ee48a74} /* (10, 17, 2) {real, imag} */,
  {32'hbfad54d5, 32'hbf8193fb} /* (10, 17, 1) {real, imag} */,
  {32'hbea97e24, 32'hbf4dde4a} /* (10, 17, 0) {real, imag} */,
  {32'h3f6b83f0, 32'h3c8a76a0} /* (10, 16, 31) {real, imag} */,
  {32'h3fb2e144, 32'hbf1f5108} /* (10, 16, 30) {real, imag} */,
  {32'h3fbe11bd, 32'hbf9a718a} /* (10, 16, 29) {real, imag} */,
  {32'h3f836dd3, 32'hbee1c500} /* (10, 16, 28) {real, imag} */,
  {32'hbbd8f500, 32'hbf0e6040} /* (10, 16, 27) {real, imag} */,
  {32'hbdf69d30, 32'hbfbd2201} /* (10, 16, 26) {real, imag} */,
  {32'h3f8008a6, 32'hbf083b64} /* (10, 16, 25) {real, imag} */,
  {32'h3f9a86d4, 32'h3fadff0b} /* (10, 16, 24) {real, imag} */,
  {32'h3ea47480, 32'h3f472d40} /* (10, 16, 23) {real, imag} */,
  {32'hbf8f3444, 32'h3dfef040} /* (10, 16, 22) {real, imag} */,
  {32'hc00c0669, 32'hbf0d20f1} /* (10, 16, 21) {real, imag} */,
  {32'hbfdd3463, 32'hbebdcf20} /* (10, 16, 20) {real, imag} */,
  {32'hbfa30386, 32'hbf46a8ba} /* (10, 16, 19) {real, imag} */,
  {32'hc007312c, 32'hbf1e8000} /* (10, 16, 18) {real, imag} */,
  {32'hc0011bd4, 32'h3d38aa40} /* (10, 16, 17) {real, imag} */,
  {32'hbf1a7c44, 32'h3f425d06} /* (10, 16, 16) {real, imag} */,
  {32'h3eabb02c, 32'h3ca758c0} /* (10, 16, 15) {real, imag} */,
  {32'hbe7e14a8, 32'hbed98620} /* (10, 16, 14) {real, imag} */,
  {32'hbfaea407, 32'h3f98614f} /* (10, 16, 13) {real, imag} */,
  {32'hbf2b08bc, 32'h3f512456} /* (10, 16, 12) {real, imag} */,
  {32'hbfcd14a2, 32'hbed4c580} /* (10, 16, 11) {real, imag} */,
  {32'h3f633c33, 32'hbee860a4} /* (10, 16, 10) {real, imag} */,
  {32'h3ff65334, 32'hc003c44f} /* (10, 16, 9) {real, imag} */,
  {32'h3f82a738, 32'hbfb70d5f} /* (10, 16, 8) {real, imag} */,
  {32'h3fc64182, 32'hbe00bf14} /* (10, 16, 7) {real, imag} */,
  {32'h3fcd83ef, 32'h3f16398e} /* (10, 16, 6) {real, imag} */,
  {32'h3f711628, 32'hbf45af2e} /* (10, 16, 5) {real, imag} */,
  {32'h3ff74f30, 32'hbf0855da} /* (10, 16, 4) {real, imag} */,
  {32'h3fcf4af2, 32'h3f8213c1} /* (10, 16, 3) {real, imag} */,
  {32'hbe4d2d20, 32'h3fb8ccaf} /* (10, 16, 2) {real, imag} */,
  {32'hc00d6f9f, 32'hbf254b07} /* (10, 16, 1) {real, imag} */,
  {32'hbf48f42c, 32'hbf856f32} /* (10, 16, 0) {real, imag} */,
  {32'h3f06af20, 32'h3c685640} /* (10, 15, 31) {real, imag} */,
  {32'h3fa9515a, 32'hbe8f81b8} /* (10, 15, 30) {real, imag} */,
  {32'h3f9c6d37, 32'hbda64008} /* (10, 15, 29) {real, imag} */,
  {32'h3f94b8e4, 32'h3f35d84a} /* (10, 15, 28) {real, imag} */,
  {32'h3f1239f2, 32'hbf0a7578} /* (10, 15, 27) {real, imag} */,
  {32'h3f3d76c6, 32'hbf733fde} /* (10, 15, 26) {real, imag} */,
  {32'h3e5eff78, 32'hbf82d898} /* (10, 15, 25) {real, imag} */,
  {32'h3fcbcce2, 32'hbea9d596} /* (10, 15, 24) {real, imag} */,
  {32'h400547c2, 32'h3f35bb00} /* (10, 15, 23) {real, imag} */,
  {32'h3f82afd1, 32'h3f7d34e8} /* (10, 15, 22) {real, imag} */,
  {32'hbf88b92c, 32'hbecfed6c} /* (10, 15, 21) {real, imag} */,
  {32'hbf96f709, 32'h3f4b8bda} /* (10, 15, 20) {real, imag} */,
  {32'hbfff760d, 32'h3f529a29} /* (10, 15, 19) {real, imag} */,
  {32'hc00bff80, 32'h3f800160} /* (10, 15, 18) {real, imag} */,
  {32'hbfdb1342, 32'h3ee4d390} /* (10, 15, 17) {real, imag} */,
  {32'hbed46f6e, 32'hbedee960} /* (10, 15, 16) {real, imag} */,
  {32'hbf126d14, 32'hbf6b955e} /* (10, 15, 15) {real, imag} */,
  {32'hbd17bdb0, 32'hbf38d06e} /* (10, 15, 14) {real, imag} */,
  {32'h3f0f82b1, 32'h4019bfeb} /* (10, 15, 13) {real, imag} */,
  {32'h3f441f14, 32'h4009c916} /* (10, 15, 12) {real, imag} */,
  {32'hbf5e821a, 32'hbdf2cd90} /* (10, 15, 11) {real, imag} */,
  {32'h3eb1ff80, 32'hbf4221ee} /* (10, 15, 10) {real, imag} */,
  {32'h3f82b307, 32'hbef6cd80} /* (10, 15, 9) {real, imag} */,
  {32'h3f1b759a, 32'h3ec120a6} /* (10, 15, 8) {real, imag} */,
  {32'h3f958a5a, 32'h3eedfc70} /* (10, 15, 7) {real, imag} */,
  {32'h4007836f, 32'hbf59c1da} /* (10, 15, 6) {real, imag} */,
  {32'h400d182b, 32'hbcb659c0} /* (10, 15, 5) {real, imag} */,
  {32'h3f983b82, 32'h3e4ba0e0} /* (10, 15, 4) {real, imag} */,
  {32'h3f54dd24, 32'hbe16c718} /* (10, 15, 3) {real, imag} */,
  {32'hbee4779c, 32'hbe0e80e0} /* (10, 15, 2) {real, imag} */,
  {32'hc01ddd3a, 32'hbe0ebad8} /* (10, 15, 1) {real, imag} */,
  {32'hbf83ae6c, 32'hbf18fc31} /* (10, 15, 0) {real, imag} */,
  {32'h3e8e3578, 32'hbdf71ec0} /* (10, 14, 31) {real, imag} */,
  {32'h3fbeacb0, 32'h3f32d496} /* (10, 14, 30) {real, imag} */,
  {32'h3ee16868, 32'hbe65d790} /* (10, 14, 29) {real, imag} */,
  {32'h3f0ca06c, 32'hbf59615a} /* (10, 14, 28) {real, imag} */,
  {32'h3efba1dc, 32'hbfa0997b} /* (10, 14, 27) {real, imag} */,
  {32'h3f0815a6, 32'hbfa8f012} /* (10, 14, 26) {real, imag} */,
  {32'h3e959db8, 32'hbf959042} /* (10, 14, 25) {real, imag} */,
  {32'h3f9b43e7, 32'hbfa9fa66} /* (10, 14, 24) {real, imag} */,
  {32'h3fe23835, 32'hbe671468} /* (10, 14, 23) {real, imag} */,
  {32'h4003679a, 32'h3ecd6704} /* (10, 14, 22) {real, imag} */,
  {32'h3f79bc8e, 32'h3e907962} /* (10, 14, 21) {real, imag} */,
  {32'hbf92831e, 32'h3f8e61e6} /* (10, 14, 20) {real, imag} */,
  {32'hbf888980, 32'h3f5b98f4} /* (10, 14, 19) {real, imag} */,
  {32'hbf9bbfd4, 32'h3f7586c4} /* (10, 14, 18) {real, imag} */,
  {32'hbe3b7514, 32'h3f1c654a} /* (10, 14, 17) {real, imag} */,
  {32'hbe15dfca, 32'hbfe1176a} /* (10, 14, 16) {real, imag} */,
  {32'hbf1ccd13, 32'hbf3ea842} /* (10, 14, 15) {real, imag} */,
  {32'h3fc73504, 32'h3edddb8e} /* (10, 14, 14) {real, imag} */,
  {32'h3fa7c63a, 32'h3fca4a48} /* (10, 14, 13) {real, imag} */,
  {32'hbf1044e2, 32'h3fa8f454} /* (10, 14, 12) {real, imag} */,
  {32'hbf18707c, 32'hbf1e04e4} /* (10, 14, 11) {real, imag} */,
  {32'hbf53f0c1, 32'hbf486c8a} /* (10, 14, 10) {real, imag} */,
  {32'hbf0d6a2e, 32'hbda2f870} /* (10, 14, 9) {real, imag} */,
  {32'h3edd670c, 32'h3d3afda0} /* (10, 14, 8) {real, imag} */,
  {32'h3f8fd342, 32'hbf392ab1} /* (10, 14, 7) {real, imag} */,
  {32'h3f29404e, 32'hbf0da995} /* (10, 14, 6) {real, imag} */,
  {32'h3e187b49, 32'h3fa6b173} /* (10, 14, 5) {real, imag} */,
  {32'h3f4f3b52, 32'h3f9fd48a} /* (10, 14, 4) {real, imag} */,
  {32'h3f09a0f7, 32'h3f6ca7d4} /* (10, 14, 3) {real, imag} */,
  {32'hbfa29402, 32'h3de737b0} /* (10, 14, 2) {real, imag} */,
  {32'hbfb33548, 32'h3da272c0} /* (10, 14, 1) {real, imag} */,
  {32'hbf36e159, 32'h3d9d5700} /* (10, 14, 0) {real, imag} */,
  {32'h3f6c349c, 32'h3e86d49e} /* (10, 13, 31) {real, imag} */,
  {32'h40074597, 32'h3fb5e566} /* (10, 13, 30) {real, imag} */,
  {32'hbf20fe05, 32'hbd981970} /* (10, 13, 29) {real, imag} */,
  {32'hbfa07024, 32'h3f221da6} /* (10, 13, 28) {real, imag} */,
  {32'hbf4604aa, 32'hbe463b3c} /* (10, 13, 27) {real, imag} */,
  {32'hbc35eb40, 32'hbf603bb6} /* (10, 13, 26) {real, imag} */,
  {32'h3f5f4ca8, 32'hbd935888} /* (10, 13, 25) {real, imag} */,
  {32'h3e4640c0, 32'hbf2deb48} /* (10, 13, 24) {real, imag} */,
  {32'h3f2dcd1c, 32'hbe6be418} /* (10, 13, 23) {real, imag} */,
  {32'h3f3dcf74, 32'hbef0e1bc} /* (10, 13, 22) {real, imag} */,
  {32'h3f859d7a, 32'hbf179d5f} /* (10, 13, 21) {real, imag} */,
  {32'hbf3ff868, 32'hbe53e548} /* (10, 13, 20) {real, imag} */,
  {32'h3f12615c, 32'hbd05b800} /* (10, 13, 19) {real, imag} */,
  {32'h3f98b8fd, 32'h3f32e567} /* (10, 13, 18) {real, imag} */,
  {32'hbf51e9c8, 32'h3f143fc0} /* (10, 13, 17) {real, imag} */,
  {32'hbf9aa566, 32'hbfc0365a} /* (10, 13, 16) {real, imag} */,
  {32'hbf2cf6bb, 32'hbf35d454} /* (10, 13, 15) {real, imag} */,
  {32'h3ef62e9e, 32'h3f8b92a6} /* (10, 13, 14) {real, imag} */,
  {32'h3dc11c20, 32'h40133d70} /* (10, 13, 13) {real, imag} */,
  {32'hbf4c4a6c, 32'h3f9623d9} /* (10, 13, 12) {real, imag} */,
  {32'hbdfad0b0, 32'hbf83c599} /* (10, 13, 11) {real, imag} */,
  {32'hbf3da80c, 32'hbfeb4ae5} /* (10, 13, 10) {real, imag} */,
  {32'hbf3f1644, 32'hc0148e12} /* (10, 13, 9) {real, imag} */,
  {32'hbee805b8, 32'hbf87e5f0} /* (10, 13, 8) {real, imag} */,
  {32'h3f5323aa, 32'hbde685c0} /* (10, 13, 7) {real, imag} */,
  {32'h3f9c92c0, 32'h3fa2f889} /* (10, 13, 6) {real, imag} */,
  {32'hbe3c2a58, 32'h4018fc7a} /* (10, 13, 5) {real, imag} */,
  {32'h3e5887b0, 32'h3f29bbba} /* (10, 13, 4) {real, imag} */,
  {32'h3e2a4270, 32'h3e3711e0} /* (10, 13, 3) {real, imag} */,
  {32'hbf176078, 32'hbf90244e} /* (10, 13, 2) {real, imag} */,
  {32'hbed778e0, 32'hbe07fb28} /* (10, 13, 1) {real, imag} */,
  {32'hbebb5af0, 32'hbf46a265} /* (10, 13, 0) {real, imag} */,
  {32'h3e4ddc1c, 32'hbf7eb3ca} /* (10, 12, 31) {real, imag} */,
  {32'h3f404f6f, 32'hbfae5d4a} /* (10, 12, 30) {real, imag} */,
  {32'hbd487240, 32'hbec7854a} /* (10, 12, 29) {real, imag} */,
  {32'hbe9d04a8, 32'h3f98dde2} /* (10, 12, 28) {real, imag} */,
  {32'hbe1d1ca8, 32'hbe84f286} /* (10, 12, 27) {real, imag} */,
  {32'h3f549a29, 32'hbff47691} /* (10, 12, 26) {real, imag} */,
  {32'h3f223996, 32'h3eb15348} /* (10, 12, 25) {real, imag} */,
  {32'h3e86ba78, 32'hbea69fa8} /* (10, 12, 24) {real, imag} */,
  {32'h3f1dd3db, 32'hbf9852d5} /* (10, 12, 23) {real, imag} */,
  {32'h3fe68ff1, 32'hbfc75faf} /* (10, 12, 22) {real, imag} */,
  {32'h3fb43c4d, 32'hbf3fc413} /* (10, 12, 21) {real, imag} */,
  {32'h3f29dbac, 32'h3dd7bd70} /* (10, 12, 20) {real, imag} */,
  {32'h3ff6c6c4, 32'hbecaee68} /* (10, 12, 19) {real, imag} */,
  {32'h3f174f65, 32'hbf163272} /* (10, 12, 18) {real, imag} */,
  {32'hbf91c941, 32'h3f363d7a} /* (10, 12, 17) {real, imag} */,
  {32'hbf841f05, 32'h3f4b8b3c} /* (10, 12, 16) {real, imag} */,
  {32'hbeb098c4, 32'hbe98af2e} /* (10, 12, 15) {real, imag} */,
  {32'hbf12055e, 32'h3e89ea74} /* (10, 12, 14) {real, imag} */,
  {32'hbf67b895, 32'h3f9b20bc} /* (10, 12, 13) {real, imag} */,
  {32'hbc88b170, 32'h3f99bb70} /* (10, 12, 12) {real, imag} */,
  {32'h3f9b08c6, 32'hbf0ac547} /* (10, 12, 11) {real, imag} */,
  {32'h3e8480a3, 32'hbff4a352} /* (10, 12, 10) {real, imag} */,
  {32'hbe166dbc, 32'hc047a3ea} /* (10, 12, 9) {real, imag} */,
  {32'hbf03cc96, 32'hbff50b62} /* (10, 12, 8) {real, imag} */,
  {32'h3d907470, 32'h3f0b31d8} /* (10, 12, 7) {real, imag} */,
  {32'h3f368dfc, 32'h3f9890be} /* (10, 12, 6) {real, imag} */,
  {32'hbe7c4df8, 32'h3f1fc508} /* (10, 12, 5) {real, imag} */,
  {32'h3e964e32, 32'hbf75b995} /* (10, 12, 4) {real, imag} */,
  {32'h3e7812ac, 32'hbfd1d86f} /* (10, 12, 3) {real, imag} */,
  {32'hbf26b9f6, 32'hbfbabe14} /* (10, 12, 2) {real, imag} */,
  {32'hbfb0aeaa, 32'hbd869060} /* (10, 12, 1) {real, imag} */,
  {32'hbf852a93, 32'hbf4af29c} /* (10, 12, 0) {real, imag} */,
  {32'hbf22759e, 32'hbdd5cdc8} /* (10, 11, 31) {real, imag} */,
  {32'hbcd23f70, 32'hbfa119e2} /* (10, 11, 30) {real, imag} */,
  {32'h3fa12b94, 32'hbf095d90} /* (10, 11, 29) {real, imag} */,
  {32'h3f7e333a, 32'hbf0187ba} /* (10, 11, 28) {real, imag} */,
  {32'h3e9967a4, 32'hbff7da49} /* (10, 11, 27) {real, imag} */,
  {32'hbebd60a9, 32'hbf8500a4} /* (10, 11, 26) {real, imag} */,
  {32'hbd6ff570, 32'h3f2974f2} /* (10, 11, 25) {real, imag} */,
  {32'h3fc401f8, 32'hbf9f3210} /* (10, 11, 24) {real, imag} */,
  {32'h3e3d8aae, 32'hc03b76a9} /* (10, 11, 23) {real, imag} */,
  {32'h3e8ab784, 32'hbf105f1f} /* (10, 11, 22) {real, imag} */,
  {32'hbe842074, 32'hbea05508} /* (10, 11, 21) {real, imag} */,
  {32'hbf740300, 32'hbef77a92} /* (10, 11, 20) {real, imag} */,
  {32'hbe6418ae, 32'hbf013ec2} /* (10, 11, 19) {real, imag} */,
  {32'h3f2b1cf8, 32'hbea6137c} /* (10, 11, 18) {real, imag} */,
  {32'hbe318fbc, 32'h3de5b240} /* (10, 11, 17) {real, imag} */,
  {32'hbf04fea4, 32'hbeada4d0} /* (10, 11, 16) {real, imag} */,
  {32'hbee02b0c, 32'hbe76db10} /* (10, 11, 15) {real, imag} */,
  {32'hbf985104, 32'h3e19fd74} /* (10, 11, 14) {real, imag} */,
  {32'hbf7772f4, 32'hbce0e300} /* (10, 11, 13) {real, imag} */,
  {32'hbf8aba5a, 32'h3f0d7242} /* (10, 11, 12) {real, imag} */,
  {32'h3eac7e7a, 32'hbef60f38} /* (10, 11, 11) {real, imag} */,
  {32'h3f026dfd, 32'hbfc7f308} /* (10, 11, 10) {real, imag} */,
  {32'h3f118ced, 32'hbfae4636} /* (10, 11, 9) {real, imag} */,
  {32'h3fc1e3f7, 32'hbe31e74c} /* (10, 11, 8) {real, imag} */,
  {32'hbf51b514, 32'h3f5d3960} /* (10, 11, 7) {real, imag} */,
  {32'hbfb9fbd9, 32'hbe34b870} /* (10, 11, 6) {real, imag} */,
  {32'hbda796e0, 32'hbf9e6858} /* (10, 11, 5) {real, imag} */,
  {32'h3ede18f6, 32'hbf430987} /* (10, 11, 4) {real, imag} */,
  {32'h3ebd44cc, 32'h3f0fed8f} /* (10, 11, 3) {real, imag} */,
  {32'hbfad0a3c, 32'hbe826da8} /* (10, 11, 2) {real, imag} */,
  {32'hc00465ca, 32'hbd4b1b60} /* (10, 11, 1) {real, imag} */,
  {32'hbf876466, 32'h3f134da2} /* (10, 11, 0) {real, imag} */,
  {32'hbef68852, 32'hbdd39a10} /* (10, 10, 31) {real, imag} */,
  {32'hbedfb1e0, 32'hbf11cfc0} /* (10, 10, 30) {real, imag} */,
  {32'h3f47733e, 32'hbf5d7e12} /* (10, 10, 29) {real, imag} */,
  {32'h3f7c0094, 32'hbeb41f28} /* (10, 10, 28) {real, imag} */,
  {32'h3e85c6b8, 32'hbdade4c0} /* (10, 10, 27) {real, imag} */,
  {32'hbf1a60ee, 32'hbf6bbb95} /* (10, 10, 26) {real, imag} */,
  {32'h3e752afc, 32'hbf86b5e2} /* (10, 10, 25) {real, imag} */,
  {32'h3eeeb17e, 32'hbfc922e4} /* (10, 10, 24) {real, imag} */,
  {32'hc02c8517, 32'hbf791b18} /* (10, 10, 23) {real, imag} */,
  {32'hc03524c3, 32'h3f981191} /* (10, 10, 22) {real, imag} */,
  {32'hc0164a3e, 32'hbdecb554} /* (10, 10, 21) {real, imag} */,
  {32'hbfe3bb2f, 32'hbfcdb09d} /* (10, 10, 20) {real, imag} */,
  {32'h3e125720, 32'hbeebd780} /* (10, 10, 19) {real, imag} */,
  {32'h3ffb145e, 32'h3f5a16ba} /* (10, 10, 18) {real, imag} */,
  {32'h3fa3ea71, 32'h3fbc14c0} /* (10, 10, 17) {real, imag} */,
  {32'h3e9c18c4, 32'h3ed6ab54} /* (10, 10, 16) {real, imag} */,
  {32'h3d4cc64e, 32'hbf015ef1} /* (10, 10, 15) {real, imag} */,
  {32'hbf8dba52, 32'h3ea38d80} /* (10, 10, 14) {real, imag} */,
  {32'hbf3fa0c8, 32'hbe19a1f8} /* (10, 10, 13) {real, imag} */,
  {32'hbfb76067, 32'h3f0271bd} /* (10, 10, 12) {real, imag} */,
  {32'hbf1a3166, 32'h3f7ebb14} /* (10, 10, 11) {real, imag} */,
  {32'h3f017e31, 32'hbcb83100} /* (10, 10, 10) {real, imag} */,
  {32'hbeddfa8c, 32'h3f30e86c} /* (10, 10, 9) {real, imag} */,
  {32'hbf6acf62, 32'h3eff401e} /* (10, 10, 8) {real, imag} */,
  {32'hbf8152a2, 32'h3ecb8024} /* (10, 10, 7) {real, imag} */,
  {32'hbeb607f4, 32'hbf203b62} /* (10, 10, 6) {real, imag} */,
  {32'h3e7a08d8, 32'h3d2c15d0} /* (10, 10, 5) {real, imag} */,
  {32'h3edc6f8e, 32'hbf978e60} /* (10, 10, 4) {real, imag} */,
  {32'h3e239414, 32'h3e960aea} /* (10, 10, 3) {real, imag} */,
  {32'hbebf7a80, 32'h3f4291a0} /* (10, 10, 2) {real, imag} */,
  {32'h3e993fb0, 32'hc0007a14} /* (10, 10, 1) {real, imag} */,
  {32'h3f51b440, 32'hbf80d1d8} /* (10, 10, 0) {real, imag} */,
  {32'h3ec77b6c, 32'h3ed4a1d0} /* (10, 9, 31) {real, imag} */,
  {32'hbcb7dc60, 32'hbe103e30} /* (10, 9, 30) {real, imag} */,
  {32'hbde5d0c0, 32'hbf47e2de} /* (10, 9, 29) {real, imag} */,
  {32'h3ceca1a0, 32'hbe94ee5c} /* (10, 9, 28) {real, imag} */,
  {32'h3e8dd18a, 32'h3f153f37} /* (10, 9, 27) {real, imag} */,
  {32'hbb796e00, 32'hbe82ed9e} /* (10, 9, 26) {real, imag} */,
  {32'h3f4adaf7, 32'hbf7a6fcb} /* (10, 9, 25) {real, imag} */,
  {32'h3fa26768, 32'hbe8c86c0} /* (10, 9, 24) {real, imag} */,
  {32'hbfd0759a, 32'h3fb29cea} /* (10, 9, 23) {real, imag} */,
  {32'hc00e5f12, 32'h3ff0af69} /* (10, 9, 22) {real, imag} */,
  {32'hbfbbe01c, 32'h3f06a0ba} /* (10, 9, 21) {real, imag} */,
  {32'hbfa993f3, 32'hbfca6047} /* (10, 9, 20) {real, imag} */,
  {32'h3f1eb253, 32'hbe4af998} /* (10, 9, 19) {real, imag} */,
  {32'h3fdb2d41, 32'h3f983dd2} /* (10, 9, 18) {real, imag} */,
  {32'h3f89ee3c, 32'h3f82e0e7} /* (10, 9, 17) {real, imag} */,
  {32'hbf10b2cc, 32'h3fcad4db} /* (10, 9, 16) {real, imag} */,
  {32'h3f2a09fa, 32'hbd11ba80} /* (10, 9, 15) {real, imag} */,
  {32'h3f1d6832, 32'hbe4d0a30} /* (10, 9, 14) {real, imag} */,
  {32'h3f462d94, 32'h3e3045f4} /* (10, 9, 13) {real, imag} */,
  {32'h3ed75f9e, 32'h3edfcb88} /* (10, 9, 12) {real, imag} */,
  {32'hbf90f469, 32'h3f959ea6} /* (10, 9, 11) {real, imag} */,
  {32'hbfb68760, 32'h3f5283ae} /* (10, 9, 10) {real, imag} */,
  {32'hbfd7c1c6, 32'h3f7f12a5} /* (10, 9, 9) {real, imag} */,
  {32'hbf0728a0, 32'h3eb1d0bc} /* (10, 9, 8) {real, imag} */,
  {32'h3edf09a4, 32'hbe844178} /* (10, 9, 7) {real, imag} */,
  {32'h3e5a5768, 32'hbf3a8f44} /* (10, 9, 6) {real, imag} */,
  {32'h3e826dd4, 32'hbe61b918} /* (10, 9, 5) {real, imag} */,
  {32'h3f709b5f, 32'hbfdc527d} /* (10, 9, 4) {real, imag} */,
  {32'h3f9f5412, 32'hbff59971} /* (10, 9, 3) {real, imag} */,
  {32'h3f9c1527, 32'hbf8281a6} /* (10, 9, 2) {real, imag} */,
  {32'hbf06e59d, 32'hc03d03ef} /* (10, 9, 1) {real, imag} */,
  {32'hbf2b3467, 32'hbfe2d34a} /* (10, 9, 0) {real, imag} */,
  {32'h3f26b710, 32'h3ea13794} /* (10, 8, 31) {real, imag} */,
  {32'h3fa99ecf, 32'hbece0618} /* (10, 8, 30) {real, imag} */,
  {32'hbe5b0d80, 32'hbeb49e10} /* (10, 8, 29) {real, imag} */,
  {32'h3d3dc140, 32'hbe8ace74} /* (10, 8, 28) {real, imag} */,
  {32'hbed32064, 32'h3f41955c} /* (10, 8, 27) {real, imag} */,
  {32'hbfc694a8, 32'h3f97761f} /* (10, 8, 26) {real, imag} */,
  {32'hbf19bdf1, 32'hbe8d598c} /* (10, 8, 25) {real, imag} */,
  {32'hbfbcf396, 32'h3f5b214c} /* (10, 8, 24) {real, imag} */,
  {32'hbfc0b798, 32'h3f8c5896} /* (10, 8, 23) {real, imag} */,
  {32'hbfa7adbc, 32'h3f5f876c} /* (10, 8, 22) {real, imag} */,
  {32'hbf15a22d, 32'h3fe40fd1} /* (10, 8, 21) {real, imag} */,
  {32'hbf0584a0, 32'h3e9e218a} /* (10, 8, 20) {real, imag} */,
  {32'h3f3e6d98, 32'h3fa322b8} /* (10, 8, 19) {real, imag} */,
  {32'h3fc98606, 32'h400f22bc} /* (10, 8, 18) {real, imag} */,
  {32'h3f2ed381, 32'h3f8a0ae8} /* (10, 8, 17) {real, imag} */,
  {32'hbf3d965e, 32'hbf11a482} /* (10, 8, 16) {real, imag} */,
  {32'h3f92d498, 32'hbfb1855a} /* (10, 8, 15) {real, imag} */,
  {32'h3fd04e02, 32'h3e9491f2} /* (10, 8, 14) {real, imag} */,
  {32'h3f9b351e, 32'hbf180a84} /* (10, 8, 13) {real, imag} */,
  {32'h3f911d4c, 32'hbf9c4944} /* (10, 8, 12) {real, imag} */,
  {32'hbf8feac6, 32'h3fb7bcf0} /* (10, 8, 11) {real, imag} */,
  {32'hc012306e, 32'h3f810557} /* (10, 8, 10) {real, imag} */,
  {32'hbf393f4e, 32'hbf22276c} /* (10, 8, 9) {real, imag} */,
  {32'h3f6cb9b0, 32'h3e89b9ee} /* (10, 8, 8) {real, imag} */,
  {32'h3fb80eac, 32'hbf007964} /* (10, 8, 7) {real, imag} */,
  {32'h3e63ebd8, 32'hbf66854c} /* (10, 8, 6) {real, imag} */,
  {32'hbdddbab0, 32'hbf3710d4} /* (10, 8, 5) {real, imag} */,
  {32'h3fc797c1, 32'h3eccf0d4} /* (10, 8, 4) {real, imag} */,
  {32'h3f9c45be, 32'hbfa19b1e} /* (10, 8, 3) {real, imag} */,
  {32'h3fe0c39a, 32'hbfe65ff7} /* (10, 8, 2) {real, imag} */,
  {32'hbf3317b3, 32'hbfd81cb0} /* (10, 8, 1) {real, imag} */,
  {32'hbfd745f6, 32'hbf304cb8} /* (10, 8, 0) {real, imag} */,
  {32'hbc54f180, 32'h3ea7601a} /* (10, 7, 31) {real, imag} */,
  {32'h3fbc2b14, 32'hbed6b200} /* (10, 7, 30) {real, imag} */,
  {32'h3e89aa88, 32'hbf4d6c06} /* (10, 7, 29) {real, imag} */,
  {32'hbfce2325, 32'hbf208b41} /* (10, 7, 28) {real, imag} */,
  {32'hbf83887b, 32'hbe8271a2} /* (10, 7, 27) {real, imag} */,
  {32'hbf320f76, 32'h3efc35b0} /* (10, 7, 26) {real, imag} */,
  {32'hbe988710, 32'hbf921cf6} /* (10, 7, 25) {real, imag} */,
  {32'h3ede1ff4, 32'hbf2cc06e} /* (10, 7, 24) {real, imag} */,
  {32'h3dbb7cd0, 32'h3eeb7e88} /* (10, 7, 23) {real, imag} */,
  {32'hbf48bd3a, 32'hbdfa3a70} /* (10, 7, 22) {real, imag} */,
  {32'hbf1c294f, 32'hbe19aa18} /* (10, 7, 21) {real, imag} */,
  {32'hbf541860, 32'h3dadb888} /* (10, 7, 20) {real, imag} */,
  {32'h3eebeca8, 32'hbeed4ab4} /* (10, 7, 19) {real, imag} */,
  {32'h3ed0cea2, 32'h3f8e93ce} /* (10, 7, 18) {real, imag} */,
  {32'h3f2c1ae4, 32'h3f3c5374} /* (10, 7, 17) {real, imag} */,
  {32'hbf97a87d, 32'hbf5dce26} /* (10, 7, 16) {real, imag} */,
  {32'hbe956798, 32'hc00f5c2e} /* (10, 7, 15) {real, imag} */,
  {32'h400a4b4e, 32'hbf84fa4e} /* (10, 7, 14) {real, imag} */,
  {32'h3f931744, 32'hbfbb0467} /* (10, 7, 13) {real, imag} */,
  {32'hbf25543b, 32'hc0106c46} /* (10, 7, 12) {real, imag} */,
  {32'hbe93dc74, 32'h3f51802f} /* (10, 7, 11) {real, imag} */,
  {32'hbf9a61f3, 32'h3f1bbbe4} /* (10, 7, 10) {real, imag} */,
  {32'hbf6203f8, 32'hbf11310a} /* (10, 7, 9) {real, imag} */,
  {32'hbf5488bb, 32'h3dd36210} /* (10, 7, 8) {real, imag} */,
  {32'hbf854184, 32'hbf916b3a} /* (10, 7, 7) {real, imag} */,
  {32'hbe09d36c, 32'hbf6a362e} /* (10, 7, 6) {real, imag} */,
  {32'hbefc83fc, 32'h3cb02480} /* (10, 7, 5) {real, imag} */,
  {32'h3f81492a, 32'h3fc48344} /* (10, 7, 4) {real, imag} */,
  {32'h3eae66f6, 32'hbe4cd5c0} /* (10, 7, 3) {real, imag} */,
  {32'hbf131474, 32'hbedd9a14} /* (10, 7, 2) {real, imag} */,
  {32'h3e643a34, 32'hbfa8c5ed} /* (10, 7, 1) {real, imag} */,
  {32'hbebe25e8, 32'hbf5289ee} /* (10, 7, 0) {real, imag} */,
  {32'h3f11f4d4, 32'h3ca92f80} /* (10, 6, 31) {real, imag} */,
  {32'h3f3a3622, 32'hbf49d127} /* (10, 6, 30) {real, imag} */,
  {32'h3f7286fa, 32'hbb7f9a00} /* (10, 6, 29) {real, imag} */,
  {32'hbf3ab2b6, 32'hbe941776} /* (10, 6, 28) {real, imag} */,
  {32'hbed66518, 32'hbfb19032} /* (10, 6, 27) {real, imag} */,
  {32'hbf1495d0, 32'hbf06c3d6} /* (10, 6, 26) {real, imag} */,
  {32'h3e25b428, 32'hbfb4c35f} /* (10, 6, 25) {real, imag} */,
  {32'h3f05c060, 32'hbd09d920} /* (10, 6, 24) {real, imag} */,
  {32'h3f64ae53, 32'h3f575a50} /* (10, 6, 23) {real, imag} */,
  {32'h3d1800d0, 32'h3ed695f0} /* (10, 6, 22) {real, imag} */,
  {32'h3f5bd042, 32'h3adff000} /* (10, 6, 21) {real, imag} */,
  {32'h3f571206, 32'h3e99a130} /* (10, 6, 20) {real, imag} */,
  {32'h3fa61d55, 32'hbf2b0cd0} /* (10, 6, 19) {real, imag} */,
  {32'h3f83e7a5, 32'hbe7bec7c} /* (10, 6, 18) {real, imag} */,
  {32'h3fb4a464, 32'hbe8070e6} /* (10, 6, 17) {real, imag} */,
  {32'hbee6605c, 32'hbf94f943} /* (10, 6, 16) {real, imag} */,
  {32'hbe839a9c, 32'hbf34a8d8} /* (10, 6, 15) {real, imag} */,
  {32'h40050340, 32'hbe290ed0} /* (10, 6, 14) {real, imag} */,
  {32'h3e4d04e4, 32'hbf58ee3d} /* (10, 6, 13) {real, imag} */,
  {32'hbf7862ad, 32'hbf5004a5} /* (10, 6, 12) {real, imag} */,
  {32'h3ebbc644, 32'h3f7f4203} /* (10, 6, 11) {real, imag} */,
  {32'h3dc402f0, 32'h3f53c19e} /* (10, 6, 10) {real, imag} */,
  {32'hbfbf5055, 32'h3f3ffba2} /* (10, 6, 9) {real, imag} */,
  {32'hbfb1da66, 32'h3f1661f3} /* (10, 6, 8) {real, imag} */,
  {32'hbfc857cc, 32'h3f4ea0b6} /* (10, 6, 7) {real, imag} */,
  {32'hbf9d4ac9, 32'h3f995898} /* (10, 6, 6) {real, imag} */,
  {32'h3eb0f958, 32'h3fd07b96} /* (10, 6, 5) {real, imag} */,
  {32'h3f66487a, 32'h3ff4e378} /* (10, 6, 4) {real, imag} */,
  {32'h3ea88f46, 32'hbd983378} /* (10, 6, 3) {real, imag} */,
  {32'hbf3810ae, 32'hc007ab00} /* (10, 6, 2) {real, imag} */,
  {32'hbf6b1d54, 32'hc01862bc} /* (10, 6, 1) {real, imag} */,
  {32'h3bb77e00, 32'hbf4df206} /* (10, 6, 0) {real, imag} */,
  {32'h3dda31b0, 32'h3f23a69c} /* (10, 5, 31) {real, imag} */,
  {32'hbfa63a9c, 32'h3d1b9090} /* (10, 5, 30) {real, imag} */,
  {32'hbf3ff222, 32'h3f4c2400} /* (10, 5, 29) {real, imag} */,
  {32'hbff2a052, 32'h3f060c2e} /* (10, 5, 28) {real, imag} */,
  {32'hbf9bedc7, 32'h3dd52790} /* (10, 5, 27) {real, imag} */,
  {32'hbc759700, 32'h3fbccb5c} /* (10, 5, 26) {real, imag} */,
  {32'h3eee947e, 32'h3e1ceb38} /* (10, 5, 25) {real, imag} */,
  {32'hbfedb6cc, 32'h3fb7fa1f} /* (10, 5, 24) {real, imag} */,
  {32'hbf08303c, 32'h3ff7a97a} /* (10, 5, 23) {real, imag} */,
  {32'h3e8fca4c, 32'h3e2cc428} /* (10, 5, 22) {real, imag} */,
  {32'h402abdb8, 32'hbcaeabe0} /* (10, 5, 21) {real, imag} */,
  {32'h3fcdb06c, 32'h3f550cee} /* (10, 5, 20) {real, imag} */,
  {32'h3facae82, 32'h3dbe5b36} /* (10, 5, 19) {real, imag} */,
  {32'h3f09e23e, 32'hbe98be1b} /* (10, 5, 18) {real, imag} */,
  {32'h3fead6ec, 32'hbe66aefc} /* (10, 5, 17) {real, imag} */,
  {32'h3c1aab80, 32'hbed89adc} /* (10, 5, 16) {real, imag} */,
  {32'hbf8a4069, 32'h3f9aa06d} /* (10, 5, 15) {real, imag} */,
  {32'h3fb9e670, 32'h3f92c419} /* (10, 5, 14) {real, imag} */,
  {32'hbe9d00e2, 32'h3f230a32} /* (10, 5, 13) {real, imag} */,
  {32'hbfc3f4b2, 32'h3f113164} /* (10, 5, 12) {real, imag} */,
  {32'hbeead350, 32'hbebf1f18} /* (10, 5, 11) {real, imag} */,
  {32'h3f9647da, 32'h3ec1ba9e} /* (10, 5, 10) {real, imag} */,
  {32'h3f0ed9c0, 32'hbda49984} /* (10, 5, 9) {real, imag} */,
  {32'h3f11c3e2, 32'hbe5faa64} /* (10, 5, 8) {real, imag} */,
  {32'hbe3d5260, 32'h3ebc9290} /* (10, 5, 7) {real, imag} */,
  {32'h3f4c66ed, 32'h3fa92a3d} /* (10, 5, 6) {real, imag} */,
  {32'hbd419580, 32'h3f64b8d4} /* (10, 5, 5) {real, imag} */,
  {32'h3e7fc81c, 32'h3fd564a1} /* (10, 5, 4) {real, imag} */,
  {32'hbf2e35af, 32'h3eded8f8} /* (10, 5, 3) {real, imag} */,
  {32'hbfefa419, 32'hc015dd84} /* (10, 5, 2) {real, imag} */,
  {32'hbf8e3469, 32'hc00785bb} /* (10, 5, 1) {real, imag} */,
  {32'h3e598a20, 32'hbdd4b0b4} /* (10, 5, 0) {real, imag} */,
  {32'h3dabbd00, 32'h3ed3830e} /* (10, 4, 31) {real, imag} */,
  {32'hbf670e29, 32'h3db00980} /* (10, 4, 30) {real, imag} */,
  {32'hbfce6e22, 32'h3f8093e8} /* (10, 4, 29) {real, imag} */,
  {32'hc0288538, 32'h3f8fa86c} /* (10, 4, 28) {real, imag} */,
  {32'hbfd395cc, 32'h3dd9e010} /* (10, 4, 27) {real, imag} */,
  {32'h3f8dc1ea, 32'h3e7d5290} /* (10, 4, 26) {real, imag} */,
  {32'h3f54d6ee, 32'h3e6af7e8} /* (10, 4, 25) {real, imag} */,
  {32'hbee22dee, 32'h3fb764d8} /* (10, 4, 24) {real, imag} */,
  {32'hbf2bbe6c, 32'h3ec844f8} /* (10, 4, 23) {real, imag} */,
  {32'hbe817b60, 32'hbfa8963c} /* (10, 4, 22) {real, imag} */,
  {32'h4006408e, 32'hc01bf06f} /* (10, 4, 21) {real, imag} */,
  {32'h3f616f90, 32'hbefaadb0} /* (10, 4, 20) {real, imag} */,
  {32'h3ea1bda4, 32'h3e4e9328} /* (10, 4, 19) {real, imag} */,
  {32'h3f7119b1, 32'h3d334fc0} /* (10, 4, 18) {real, imag} */,
  {32'h3e912594, 32'hbeacee20} /* (10, 4, 17) {real, imag} */,
  {32'hbfba62d9, 32'hbfa43882} /* (10, 4, 16) {real, imag} */,
  {32'hbfa5c83e, 32'hbf1b69e7} /* (10, 4, 15) {real, imag} */,
  {32'h3e2d7bf0, 32'hbf52ef96} /* (10, 4, 14) {real, imag} */,
  {32'h3f704db9, 32'hbf527ae2} /* (10, 4, 13) {real, imag} */,
  {32'h3e6dccc8, 32'h3e1350d8} /* (10, 4, 12) {real, imag} */,
  {32'h3f819e00, 32'hbba50980} /* (10, 4, 11) {real, imag} */,
  {32'h3f233e3a, 32'h3f0f3976} /* (10, 4, 10) {real, imag} */,
  {32'h3fd673d2, 32'h3f153ca6} /* (10, 4, 9) {real, imag} */,
  {32'h402c24ee, 32'hbf48aef1} /* (10, 4, 8) {real, imag} */,
  {32'h3e235810, 32'hbfbf0670} /* (10, 4, 7) {real, imag} */,
  {32'h3f3cf35b, 32'hbfaed8ba} /* (10, 4, 6) {real, imag} */,
  {32'hbe773120, 32'hbf5c1462} /* (10, 4, 5) {real, imag} */,
  {32'hbeae1cfc, 32'h3f95c8b9} /* (10, 4, 4) {real, imag} */,
  {32'hbf200388, 32'h3f5eaed4} /* (10, 4, 3) {real, imag} */,
  {32'hbe7ec5a0, 32'hbc724800} /* (10, 4, 2) {real, imag} */,
  {32'h3f248802, 32'h3ef55000} /* (10, 4, 1) {real, imag} */,
  {32'h3f2a72f5, 32'h3f5e2c53} /* (10, 4, 0) {real, imag} */,
  {32'hbeacf858, 32'h3ef51b40} /* (10, 3, 31) {real, imag} */,
  {32'hbf5c5da4, 32'h3f81f464} /* (10, 3, 30) {real, imag} */,
  {32'hc009dd28, 32'h3fefd1ab} /* (10, 3, 29) {real, imag} */,
  {32'hbf583c5e, 32'h3f6c7c37} /* (10, 3, 28) {real, imag} */,
  {32'hbf925496, 32'hbf7c3518} /* (10, 3, 27) {real, imag} */,
  {32'hbf9966e4, 32'hbf009ee2} /* (10, 3, 26) {real, imag} */,
  {32'hbf9b1058, 32'h3eddb1a8} /* (10, 3, 25) {real, imag} */,
  {32'hbe55a750, 32'h3f06db85} /* (10, 3, 24) {real, imag} */,
  {32'hbfa81a81, 32'hbe1f7c9c} /* (10, 3, 23) {real, imag} */,
  {32'hbf838d7c, 32'hbf4899d0} /* (10, 3, 22) {real, imag} */,
  {32'hbd85def8, 32'hc01970f8} /* (10, 3, 21) {real, imag} */,
  {32'hbfa1e2d1, 32'hbe518be8} /* (10, 3, 20) {real, imag} */,
  {32'hbf5a6bfc, 32'h3fb91649} /* (10, 3, 19) {real, imag} */,
  {32'h3e723eb8, 32'h402278bc} /* (10, 3, 18) {real, imag} */,
  {32'h3ec49f74, 32'h3f536240} /* (10, 3, 17) {real, imag} */,
  {32'hbee3aaa8, 32'hbe410150} /* (10, 3, 16) {real, imag} */,
  {32'hbe3c0f22, 32'hc0089e5f} /* (10, 3, 15) {real, imag} */,
  {32'hbf26ae35, 32'hc008e944} /* (10, 3, 14) {real, imag} */,
  {32'h3f45c336, 32'hbf77011e} /* (10, 3, 13) {real, imag} */,
  {32'h3fd94dd0, 32'hbf0c6716} /* (10, 3, 12) {real, imag} */,
  {32'h3f1f42ca, 32'hbd86d3b0} /* (10, 3, 11) {real, imag} */,
  {32'h3f6a5c7a, 32'hbf6a97a2} /* (10, 3, 10) {real, imag} */,
  {32'h3f291af0, 32'hbf63d523} /* (10, 3, 9) {real, imag} */,
  {32'h3faa6b83, 32'hbbbe3b00} /* (10, 3, 8) {real, imag} */,
  {32'h3f494c48, 32'h3e6c5d50} /* (10, 3, 7) {real, imag} */,
  {32'h3fc62da6, 32'hbf9e9aa3} /* (10, 3, 6) {real, imag} */,
  {32'h3e8f2f5b, 32'hbf824d25} /* (10, 3, 5) {real, imag} */,
  {32'hbf19779e, 32'h3d9ec4f0} /* (10, 3, 4) {real, imag} */,
  {32'hbeb76044, 32'h3d325980} /* (10, 3, 3) {real, imag} */,
  {32'hbf14ecdc, 32'hbf3eaf1e} /* (10, 3, 2) {real, imag} */,
  {32'h3ade3800, 32'h3f0170e0} /* (10, 3, 1) {real, imag} */,
  {32'h3ec30688, 32'h3f5a3af6} /* (10, 3, 0) {real, imag} */,
  {32'hbf05ee4e, 32'h3f1d86b1} /* (10, 2, 31) {real, imag} */,
  {32'hbf71762d, 32'h3d9f1fe0} /* (10, 2, 30) {real, imag} */,
  {32'hbf244812, 32'hbd1e4060} /* (10, 2, 29) {real, imag} */,
  {32'hbd476a00, 32'h3f089b8a} /* (10, 2, 28) {real, imag} */,
  {32'hbe5e5e30, 32'h3f5c4776} /* (10, 2, 27) {real, imag} */,
  {32'hbf20dc36, 32'h3f7a17d0} /* (10, 2, 26) {real, imag} */,
  {32'h3e935108, 32'h3fc45b3c} /* (10, 2, 25) {real, imag} */,
  {32'hbddae8a0, 32'h3fcebbb6} /* (10, 2, 24) {real, imag} */,
  {32'hbfa138cf, 32'h3f145f80} /* (10, 2, 23) {real, imag} */,
  {32'h3e21fe00, 32'h3e74d9bc} /* (10, 2, 22) {real, imag} */,
  {32'h3f4496a4, 32'hc00efc95} /* (10, 2, 21) {real, imag} */,
  {32'hbd83a020, 32'hbef558c0} /* (10, 2, 20) {real, imag} */,
  {32'h3e279500, 32'h3f0c2b58} /* (10, 2, 19) {real, imag} */,
  {32'h3f9eecfa, 32'h4001f343} /* (10, 2, 18) {real, imag} */,
  {32'h3f80478d, 32'h3face948} /* (10, 2, 17) {real, imag} */,
  {32'h3f0efe85, 32'h3ff6b654} /* (10, 2, 16) {real, imag} */,
  {32'h3f734a8c, 32'hbe84befc} /* (10, 2, 15) {real, imag} */,
  {32'h3ee5f5a8, 32'hbf9644da} /* (10, 2, 14) {real, imag} */,
  {32'h3e5b7480, 32'hc01763f1} /* (10, 2, 13) {real, imag} */,
  {32'h3f259ad9, 32'hbf8dea09} /* (10, 2, 12) {real, imag} */,
  {32'hbe0ca7b8, 32'hbc31c480} /* (10, 2, 11) {real, imag} */,
  {32'h3f51ab5c, 32'hbf7ec7fa} /* (10, 2, 10) {real, imag} */,
  {32'h3fd597bb, 32'hbdc6aa40} /* (10, 2, 9) {real, imag} */,
  {32'h3f4cf798, 32'h3f81f829} /* (10, 2, 8) {real, imag} */,
  {32'h3f66462d, 32'h3fa263c6} /* (10, 2, 7) {real, imag} */,
  {32'h40006778, 32'hbe831b14} /* (10, 2, 6) {real, imag} */,
  {32'h3f2616b4, 32'h3e44b870} /* (10, 2, 5) {real, imag} */,
  {32'hbd6c1700, 32'h3f1a9fb8} /* (10, 2, 4) {real, imag} */,
  {32'hbf9b574a, 32'h3e1f2adc} /* (10, 2, 3) {real, imag} */,
  {32'hbfe5cb1e, 32'hbf425448} /* (10, 2, 2) {real, imag} */,
  {32'hbe80a05c, 32'hbd807ab0} /* (10, 2, 1) {real, imag} */,
  {32'h3ef99e8c, 32'h3f7c6a8e} /* (10, 2, 0) {real, imag} */,
  {32'hbecb41e8, 32'h3d0c3340} /* (10, 1, 31) {real, imag} */,
  {32'hbfbb6524, 32'hbf28ba26} /* (10, 1, 30) {real, imag} */,
  {32'hbf77ac35, 32'hbf2b934c} /* (10, 1, 29) {real, imag} */,
  {32'hbf37e950, 32'hbf02f17e} /* (10, 1, 28) {real, imag} */,
  {32'h3dfd02e0, 32'h3f0d1caa} /* (10, 1, 27) {real, imag} */,
  {32'h3ec4e11e, 32'hbf3040ee} /* (10, 1, 26) {real, imag} */,
  {32'hbe985fd8, 32'hbe87b6f4} /* (10, 1, 25) {real, imag} */,
  {32'hbf482348, 32'h3fafaf33} /* (10, 1, 24) {real, imag} */,
  {32'h3e81539c, 32'h40019ff2} /* (10, 1, 23) {real, imag} */,
  {32'hbdb0c778, 32'h3e8d9a06} /* (10, 1, 22) {real, imag} */,
  {32'h3e551abc, 32'hbfc0ccf4} /* (10, 1, 21) {real, imag} */,
  {32'h3fa987c2, 32'hbf720816} /* (10, 1, 20) {real, imag} */,
  {32'h3f5585c8, 32'hbef2ba08} /* (10, 1, 19) {real, imag} */,
  {32'h3fe6ae4c, 32'h3f47d9ec} /* (10, 1, 18) {real, imag} */,
  {32'h3f849cc9, 32'h3eddd1ba} /* (10, 1, 17) {real, imag} */,
  {32'hbf135e6e, 32'h3f5ab1d7} /* (10, 1, 16) {real, imag} */,
  {32'h3eb55fde, 32'hbdc38d18} /* (10, 1, 15) {real, imag} */,
  {32'h3eb5a838, 32'hbfc0262a} /* (10, 1, 14) {real, imag} */,
  {32'hbfa6bbdc, 32'hc0224760} /* (10, 1, 13) {real, imag} */,
  {32'hbf2d6b40, 32'hbf818ac4} /* (10, 1, 12) {real, imag} */,
  {32'hbf55b784, 32'h3f46ae70} /* (10, 1, 11) {real, imag} */,
  {32'h3daf4d48, 32'h3cbf9cc0} /* (10, 1, 10) {real, imag} */,
  {32'h3fd9f11c, 32'hbf79acd8} /* (10, 1, 9) {real, imag} */,
  {32'h4033b35c, 32'hbed1f3b4} /* (10, 1, 8) {real, imag} */,
  {32'h3fec0585, 32'hbf102b86} /* (10, 1, 7) {real, imag} */,
  {32'h3f953466, 32'hbf3c0372} /* (10, 1, 6) {real, imag} */,
  {32'h3fbb206c, 32'h3f82535b} /* (10, 1, 5) {real, imag} */,
  {32'h3fa5821f, 32'h3fc21db5} /* (10, 1, 4) {real, imag} */,
  {32'hbe7d7464, 32'hbef50784} /* (10, 1, 3) {real, imag} */,
  {32'hbed6eb27, 32'hbfcbb2d1} /* (10, 1, 2) {real, imag} */,
  {32'hbeef66e6, 32'hbf1f844d} /* (10, 1, 1) {real, imag} */,
  {32'hbefe8de6, 32'h3dd0c8c0} /* (10, 1, 0) {real, imag} */,
  {32'h3e43bc7c, 32'hbe405bfc} /* (10, 0, 31) {real, imag} */,
  {32'hbec3235e, 32'hbea03d36} /* (10, 0, 30) {real, imag} */,
  {32'hbf932f3b, 32'hbe8d05f0} /* (10, 0, 29) {real, imag} */,
  {32'hbf2d9b50, 32'hbe9a62b0} /* (10, 0, 28) {real, imag} */,
  {32'h3ed1b1b6, 32'hbebd24ca} /* (10, 0, 27) {real, imag} */,
  {32'hbe2f8aa0, 32'hbf581b7d} /* (10, 0, 26) {real, imag} */,
  {32'hbfbdda10, 32'h3e27b36a} /* (10, 0, 25) {real, imag} */,
  {32'hbfc39a24, 32'h3fa79822} /* (10, 0, 24) {real, imag} */,
  {32'h3dd486f0, 32'h401c57ee} /* (10, 0, 23) {real, imag} */,
  {32'hbf3dab2a, 32'h3f3a46c6} /* (10, 0, 22) {real, imag} */,
  {32'h3d910034, 32'h3da6bde0} /* (10, 0, 21) {real, imag} */,
  {32'h3fd579ec, 32'hbef1fff0} /* (10, 0, 20) {real, imag} */,
  {32'h3ec5e580, 32'hbebb336e} /* (10, 0, 19) {real, imag} */,
  {32'h3f211942, 32'hbf4b0ddd} /* (10, 0, 18) {real, imag} */,
  {32'h3f60dd5c, 32'hbf8f6462} /* (10, 0, 17) {real, imag} */,
  {32'hbf42b574, 32'hbd615b84} /* (10, 0, 16) {real, imag} */,
  {32'h3ed1663d, 32'hbf869221} /* (10, 0, 15) {real, imag} */,
  {32'h3fbf31fa, 32'hbfa35cd6} /* (10, 0, 14) {real, imag} */,
  {32'hbee925ec, 32'hbf4f0a64} /* (10, 0, 13) {real, imag} */,
  {32'hbf6b74e9, 32'hbe604bac} /* (10, 0, 12) {real, imag} */,
  {32'hbe7c1140, 32'h3daf3f40} /* (10, 0, 11) {real, imag} */,
  {32'hbe3c47e8, 32'hbe09e56c} /* (10, 0, 10) {real, imag} */,
  {32'h3f207bf3, 32'hbf1d51bc} /* (10, 0, 9) {real, imag} */,
  {32'h400271d4, 32'hbec218d0} /* (10, 0, 8) {real, imag} */,
  {32'h3fd56fbb, 32'h3cf67400} /* (10, 0, 7) {real, imag} */,
  {32'h3f743424, 32'h3ea47924} /* (10, 0, 6) {real, imag} */,
  {32'h3f7c4c76, 32'h3f751019} /* (10, 0, 5) {real, imag} */,
  {32'h3f622764, 32'h3f88afbd} /* (10, 0, 4) {real, imag} */,
  {32'hbe979f46, 32'hbe15c85c} /* (10, 0, 3) {real, imag} */,
  {32'hbe482338, 32'hbf4d17b7} /* (10, 0, 2) {real, imag} */,
  {32'h3d0bb540, 32'hbfab0aa6} /* (10, 0, 1) {real, imag} */,
  {32'h3e5a14a6, 32'hbeb894c0} /* (10, 0, 0) {real, imag} */,
  {32'hbe7092c4, 32'h3f6a6604} /* (9, 31, 31) {real, imag} */,
  {32'hbe5fd6b8, 32'h3f4702fa} /* (9, 31, 30) {real, imag} */,
  {32'hbfa39d41, 32'hbe6e1240} /* (9, 31, 29) {real, imag} */,
  {32'hbfbd719b, 32'h3f2150a0} /* (9, 31, 28) {real, imag} */,
  {32'hbf142c60, 32'h3de10f28} /* (9, 31, 27) {real, imag} */,
  {32'hbf110686, 32'h3fbd8744} /* (9, 31, 26) {real, imag} */,
  {32'hbfdf8496, 32'h3f8de650} /* (9, 31, 25) {real, imag} */,
  {32'hbf40c672, 32'h3f922778} /* (9, 31, 24) {real, imag} */,
  {32'h3f3e6a90, 32'h3f4a340d} /* (9, 31, 23) {real, imag} */,
  {32'h3f90e59f, 32'h3e33412a} /* (9, 31, 22) {real, imag} */,
  {32'hbe8d4c0e, 32'h3e86ba05} /* (9, 31, 21) {real, imag} */,
  {32'hbe044f48, 32'h3ec631f4} /* (9, 31, 20) {real, imag} */,
  {32'h3f842e11, 32'h3e4cf80c} /* (9, 31, 19) {real, imag} */,
  {32'hbd4ee2b8, 32'hbf7e1a4a} /* (9, 31, 18) {real, imag} */,
  {32'hbf88859c, 32'h3de63fd4} /* (9, 31, 17) {real, imag} */,
  {32'hbf87c6b9, 32'h3eacefbf} /* (9, 31, 16) {real, imag} */,
  {32'hbe6f663d, 32'hbf0586c2} /* (9, 31, 15) {real, imag} */,
  {32'h3ffae518, 32'h3e7a763f} /* (9, 31, 14) {real, imag} */,
  {32'h402efd1a, 32'hbece33ac} /* (9, 31, 13) {real, imag} */,
  {32'hbe133f88, 32'hbf1d9482} /* (9, 31, 12) {real, imag} */,
  {32'hbf494d9d, 32'h3e956d22} /* (9, 31, 11) {real, imag} */,
  {32'h3de3d142, 32'hbf789394} /* (9, 31, 10) {real, imag} */,
  {32'hbdbb6ea8, 32'h3e99585f} /* (9, 31, 9) {real, imag} */,
  {32'hbe7c5ac4, 32'h3f3fc72a} /* (9, 31, 8) {real, imag} */,
  {32'h3f14e32c, 32'hbeab773c} /* (9, 31, 7) {real, imag} */,
  {32'h3e82dfd4, 32'hbf80c95f} /* (9, 31, 6) {real, imag} */,
  {32'h3e31ce08, 32'hbd6f6740} /* (9, 31, 5) {real, imag} */,
  {32'h3ecb4805, 32'h3ec2c3ca} /* (9, 31, 4) {real, imag} */,
  {32'h3eaec606, 32'hbf38562f} /* (9, 31, 3) {real, imag} */,
  {32'h3ecd62c0, 32'hbfa1a424} /* (9, 31, 2) {real, imag} */,
  {32'hbdc2c0c8, 32'h3d8ccc60} /* (9, 31, 1) {real, imag} */,
  {32'hbdf32578, 32'h3e264500} /* (9, 31, 0) {real, imag} */,
  {32'hc000638a, 32'h3f274a96} /* (9, 30, 31) {real, imag} */,
  {32'hc010bc27, 32'h3e2b3300} /* (9, 30, 30) {real, imag} */,
  {32'hc0150320, 32'h3f8dfe70} /* (9, 30, 29) {real, imag} */,
  {32'hbf7381d3, 32'h3f2605ee} /* (9, 30, 28) {real, imag} */,
  {32'hbf2e3744, 32'hbe850e55} /* (9, 30, 27) {real, imag} */,
  {32'hbf059d62, 32'h403415b0} /* (9, 30, 26) {real, imag} */,
  {32'hbfb09127, 32'h3fd6d360} /* (9, 30, 25) {real, imag} */,
  {32'hbfa7c3e5, 32'h3fbefa79} /* (9, 30, 24) {real, imag} */,
  {32'hbeb90205, 32'h3fa98ba4} /* (9, 30, 23) {real, imag} */,
  {32'hbf0fd620, 32'h3dbe3888} /* (9, 30, 22) {real, imag} */,
  {32'hbfa37c2a, 32'hbf828d1c} /* (9, 30, 21) {real, imag} */,
  {32'hbf0dc5bb, 32'hbf9e15f0} /* (9, 30, 20) {real, imag} */,
  {32'h3f68006c, 32'h3ebd8876} /* (9, 30, 19) {real, imag} */,
  {32'hbf91c4ec, 32'hbf5100d1} /* (9, 30, 18) {real, imag} */,
  {32'hc023a514, 32'hbf07cf0a} /* (9, 30, 17) {real, imag} */,
  {32'hbfa8bc75, 32'hbf39bc2a} /* (9, 30, 16) {real, imag} */,
  {32'h3e821a94, 32'hc0114e4c} /* (9, 30, 15) {real, imag} */,
  {32'h3ffa4f49, 32'hc003d32c} /* (9, 30, 14) {real, imag} */,
  {32'h4082cd22, 32'hbf9e6541} /* (9, 30, 13) {real, imag} */,
  {32'h3fa6df40, 32'hbe62eef0} /* (9, 30, 12) {real, imag} */,
  {32'hbf38ef5b, 32'hbeef8fc0} /* (9, 30, 11) {real, imag} */,
  {32'hbf46b2b5, 32'hc004df88} /* (9, 30, 10) {real, imag} */,
  {32'h3cfaab80, 32'h3f1ce2c0} /* (9, 30, 9) {real, imag} */,
  {32'hbdf67358, 32'h3f89155a} /* (9, 30, 8) {real, imag} */,
  {32'hbf010538, 32'h3efab2d0} /* (9, 30, 7) {real, imag} */,
  {32'h3bc2ad00, 32'hbfb9097c} /* (9, 30, 6) {real, imag} */,
  {32'h3e7bda58, 32'hbf75bfe3} /* (9, 30, 5) {real, imag} */,
  {32'h3ec5bce0, 32'h3f03c940} /* (9, 30, 4) {real, imag} */,
  {32'hbee1fbf2, 32'hbeb851aa} /* (9, 30, 3) {real, imag} */,
  {32'h3ec69da4, 32'hbfc09181} /* (9, 30, 2) {real, imag} */,
  {32'hbf517785, 32'hbf16c33e} /* (9, 30, 1) {real, imag} */,
  {32'hbf701ffa, 32'h3e1c4158} /* (9, 30, 0) {real, imag} */,
  {32'hc00ff6df, 32'hbf963fc8} /* (9, 29, 31) {real, imag} */,
  {32'hc0841a06, 32'hbfcd5444} /* (9, 29, 30) {real, imag} */,
  {32'hc00de1da, 32'h3fd8a175} /* (9, 29, 29) {real, imag} */,
  {32'h3bc20d80, 32'h3e1188a8} /* (9, 29, 28) {real, imag} */,
  {32'hbef7fafc, 32'hbf452bae} /* (9, 29, 27) {real, imag} */,
  {32'h3e30d530, 32'h3fdc0a16} /* (9, 29, 26) {real, imag} */,
  {32'hbf5ddab2, 32'h3f36ff7a} /* (9, 29, 25) {real, imag} */,
  {32'hbfb1a325, 32'h3d949ae0} /* (9, 29, 24) {real, imag} */,
  {32'hbf56620c, 32'h3f546df4} /* (9, 29, 23) {real, imag} */,
  {32'hbfe9dd49, 32'h3e971218} /* (9, 29, 22) {real, imag} */,
  {32'hc035c9e4, 32'hbf0c1258} /* (9, 29, 21) {real, imag} */,
  {32'hbfd327b8, 32'hbf2aeef4} /* (9, 29, 20) {real, imag} */,
  {32'h3eaea4d8, 32'hbe9544dc} /* (9, 29, 19) {real, imag} */,
  {32'hbebd2134, 32'hbe4dbaec} /* (9, 29, 18) {real, imag} */,
  {32'hbf4a3535, 32'hbf0bbc59} /* (9, 29, 17) {real, imag} */,
  {32'h3fb7a025, 32'hbf0f3db4} /* (9, 29, 16) {real, imag} */,
  {32'h3fa67c64, 32'hbfbeee2c} /* (9, 29, 15) {real, imag} */,
  {32'hbc3a0200, 32'hbf80acda} /* (9, 29, 14) {real, imag} */,
  {32'h3f83f574, 32'h3f15f02a} /* (9, 29, 13) {real, imag} */,
  {32'h3fd1d833, 32'h3f820b72} /* (9, 29, 12) {real, imag} */,
  {32'h3f926043, 32'h3ea7090e} /* (9, 29, 11) {real, imag} */,
  {32'hbf3a3632, 32'h3f39515c} /* (9, 29, 10) {real, imag} */,
  {32'hbf77b6f4, 32'h3fd7275a} /* (9, 29, 9) {real, imag} */,
  {32'hbfac0ab8, 32'h3faf1e20} /* (9, 29, 8) {real, imag} */,
  {32'hbf938a5d, 32'h3f893902} /* (9, 29, 7) {real, imag} */,
  {32'h3f183722, 32'h3f4c5dd0} /* (9, 29, 6) {real, imag} */,
  {32'hbd4bae40, 32'h3fcb9db6} /* (9, 29, 5) {real, imag} */,
  {32'hbf6e3dfd, 32'h4018cb0e} /* (9, 29, 4) {real, imag} */,
  {32'hbfe4dc36, 32'h3f1bdad0} /* (9, 29, 3) {real, imag} */,
  {32'h3f21a174, 32'h3f0b7d34} /* (9, 29, 2) {real, imag} */,
  {32'h3e3ee79c, 32'h3fdc7b2e} /* (9, 29, 1) {real, imag} */,
  {32'hbe250e0c, 32'h3e90babe} /* (9, 29, 0) {real, imag} */,
  {32'hbf18d1e2, 32'hbf5b6938} /* (9, 28, 31) {real, imag} */,
  {32'hc03d35fe, 32'hbf7c415a} /* (9, 28, 30) {real, imag} */,
  {32'hc0024bb9, 32'h3fc1d88c} /* (9, 28, 29) {real, imag} */,
  {32'hbe4d4f5a, 32'h3f59fd32} /* (9, 28, 28) {real, imag} */,
  {32'hbfa90712, 32'hbed8f160} /* (9, 28, 27) {real, imag} */,
  {32'hbe2b8ebf, 32'h3eb7b6c8} /* (9, 28, 26) {real, imag} */,
  {32'hbf5366fa, 32'h3f9de8f9} /* (9, 28, 25) {real, imag} */,
  {32'hbf9d6bcc, 32'h400dafbd} /* (9, 28, 24) {real, imag} */,
  {32'hbf17bc56, 32'hbe1f9bc8} /* (9, 28, 23) {real, imag} */,
  {32'hbf11529b, 32'hbf26f6ec} /* (9, 28, 22) {real, imag} */,
  {32'hbfc34192, 32'hbfbc84e8} /* (9, 28, 21) {real, imag} */,
  {32'h3d27bf90, 32'hc0041b40} /* (9, 28, 20) {real, imag} */,
  {32'h3ffd3ad2, 32'hbfbd1cce} /* (9, 28, 19) {real, imag} */,
  {32'h3fae1c98, 32'hbf8aff53} /* (9, 28, 18) {real, imag} */,
  {32'h3ec43730, 32'hbe4807fe} /* (9, 28, 17) {real, imag} */,
  {32'h3f1e4ce2, 32'h3bd60c00} /* (9, 28, 16) {real, imag} */,
  {32'h3f5b3e88, 32'hbdf26748} /* (9, 28, 15) {real, imag} */,
  {32'hbe397430, 32'hbe5949f0} /* (9, 28, 14) {real, imag} */,
  {32'hbc8f3ee0, 32'h3f58e8a6} /* (9, 28, 13) {real, imag} */,
  {32'h3fd71f73, 32'h3ea643ba} /* (9, 28, 12) {real, imag} */,
  {32'h3fd99a0c, 32'hbe674a2c} /* (9, 28, 11) {real, imag} */,
  {32'hbff80dd0, 32'h3f621ba0} /* (9, 28, 10) {real, imag} */,
  {32'hbf84aac3, 32'h3fccc1d2} /* (9, 28, 9) {real, imag} */,
  {32'hbdd58cb4, 32'h3b9e2000} /* (9, 28, 8) {real, imag} */,
  {32'h3f3a9433, 32'h3e93a19c} /* (9, 28, 7) {real, imag} */,
  {32'hbf4bc91e, 32'h3f8deb55} /* (9, 28, 6) {real, imag} */,
  {32'hc020c2ce, 32'h4036e358} /* (9, 28, 5) {real, imag} */,
  {32'hbf90a9a5, 32'h3f7e64ef} /* (9, 28, 4) {real, imag} */,
  {32'hbf13d80f, 32'h3f9c5c2b} /* (9, 28, 3) {real, imag} */,
  {32'hbdf12a88, 32'h3f9adb10} /* (9, 28, 2) {real, imag} */,
  {32'hbfb33380, 32'h3f46dbf6} /* (9, 28, 1) {real, imag} */,
  {32'hbfba2c36, 32'hbeb6a63c} /* (9, 28, 0) {real, imag} */,
  {32'hbea77dbe, 32'hbf80c0c2} /* (9, 27, 31) {real, imag} */,
  {32'hbe8525a0, 32'h3de5af30} /* (9, 27, 30) {real, imag} */,
  {32'h3e06fc24, 32'h40182332} /* (9, 27, 29) {real, imag} */,
  {32'hbe6889d4, 32'h400fed79} /* (9, 27, 28) {real, imag} */,
  {32'hbfbed93b, 32'h3f98315f} /* (9, 27, 27) {real, imag} */,
  {32'hc0131271, 32'hbf40bf9b} /* (9, 27, 26) {real, imag} */,
  {32'hc0144376, 32'h3f71f308} /* (9, 27, 25) {real, imag} */,
  {32'h3d124750, 32'h3ffed9fd} /* (9, 27, 24) {real, imag} */,
  {32'hbe3bf222, 32'hbfb8c161} /* (9, 27, 23) {real, imag} */,
  {32'hbfa7e78a, 32'h3d620a00} /* (9, 27, 22) {real, imag} */,
  {32'hbf93c107, 32'hbfb3e421} /* (9, 27, 21) {real, imag} */,
  {32'hbec8659c, 32'hc0159d6d} /* (9, 27, 20) {real, imag} */,
  {32'h3e997df8, 32'h3d908e60} /* (9, 27, 19) {real, imag} */,
  {32'h4012771a, 32'hbe6a476c} /* (9, 27, 18) {real, imag} */,
  {32'h3fc4af6f, 32'hbc5a9c80} /* (9, 27, 17) {real, imag} */,
  {32'hbe45c550, 32'hbf612e90} /* (9, 27, 16) {real, imag} */,
  {32'h3fd1cf88, 32'hbea2547c} /* (9, 27, 15) {real, imag} */,
  {32'h3ee3be7c, 32'h3de610a0} /* (9, 27, 14) {real, imag} */,
  {32'h3f0dd752, 32'h3e1a4dd4} /* (9, 27, 13) {real, imag} */,
  {32'h3f531672, 32'hbeb45d06} /* (9, 27, 12) {real, imag} */,
  {32'hbe376dac, 32'hbfb6758b} /* (9, 27, 11) {real, imag} */,
  {32'hbfff42c0, 32'hbf9123f8} /* (9, 27, 10) {real, imag} */,
  {32'hbfadf66b, 32'h3f813a20} /* (9, 27, 9) {real, imag} */,
  {32'hbfb595ca, 32'h3e9a55c4} /* (9, 27, 8) {real, imag} */,
  {32'h3ee701ec, 32'hbe06af38} /* (9, 27, 7) {real, imag} */,
  {32'hbf7fcb3b, 32'hbed5ba44} /* (9, 27, 6) {real, imag} */,
  {32'hbfe359e2, 32'h3fb8f8f2} /* (9, 27, 5) {real, imag} */,
  {32'hbf822043, 32'h3c527900} /* (9, 27, 4) {real, imag} */,
  {32'hbef6fa96, 32'hbcedf820} /* (9, 27, 3) {real, imag} */,
  {32'hbe269b40, 32'hbec57c91} /* (9, 27, 2) {real, imag} */,
  {32'hc03eecd4, 32'hbe133d24} /* (9, 27, 1) {real, imag} */,
  {32'hbfe175f1, 32'h3e1fb280} /* (9, 27, 0) {real, imag} */,
  {32'hbf5b144b, 32'h3e8cd704} /* (9, 26, 31) {real, imag} */,
  {32'hbfe11ed1, 32'h3eca42ba} /* (9, 26, 30) {real, imag} */,
  {32'hbf3de09d, 32'h3fed3f4c} /* (9, 26, 29) {real, imag} */,
  {32'h3fc75b38, 32'h3f710bac} /* (9, 26, 28) {real, imag} */,
  {32'h3ee6e7f2, 32'hbde557b0} /* (9, 26, 27) {real, imag} */,
  {32'hc0195010, 32'h3e12d6ac} /* (9, 26, 26) {real, imag} */,
  {32'hc018a612, 32'h3f881330} /* (9, 26, 25) {real, imag} */,
  {32'hbf8c6f10, 32'h3fb63390} /* (9, 26, 24) {real, imag} */,
  {32'hbeb68d90, 32'hbe1ef3ae} /* (9, 26, 23) {real, imag} */,
  {32'hbf203116, 32'h3ff10e0c} /* (9, 26, 22) {real, imag} */,
  {32'hbfa77294, 32'h3fcc41ed} /* (9, 26, 21) {real, imag} */,
  {32'hbf08acb6, 32'h3f7a68a3} /* (9, 26, 20) {real, imag} */,
  {32'h3f9f1288, 32'h3f1b54b8} /* (9, 26, 19) {real, imag} */,
  {32'h3fcc5d0b, 32'hbf7880d4} /* (9, 26, 18) {real, imag} */,
  {32'h3ea3afb7, 32'hbf023a2f} /* (9, 26, 17) {real, imag} */,
  {32'h3e33b438, 32'hbf43bd99} /* (9, 26, 16) {real, imag} */,
  {32'h3f9f85ce, 32'h3eaacc88} /* (9, 26, 15) {real, imag} */,
  {32'h3f10b342, 32'h3fe4e9cf} /* (9, 26, 14) {real, imag} */,
  {32'h3f1c8703, 32'h3d809fa0} /* (9, 26, 13) {real, imag} */,
  {32'h3f3e812c, 32'hbed5d966} /* (9, 26, 12) {real, imag} */,
  {32'h3f757c72, 32'hbf1a04d2} /* (9, 26, 11) {real, imag} */,
  {32'hbf656f5b, 32'hbf7b0796} /* (9, 26, 10) {real, imag} */,
  {32'hc0415f8b, 32'h3fd93efe} /* (9, 26, 9) {real, imag} */,
  {32'hc0196320, 32'h3fd5d550} /* (9, 26, 8) {real, imag} */,
  {32'hbed87440, 32'h3dbae168} /* (9, 26, 7) {real, imag} */,
  {32'hbf81f60c, 32'h3ebc5e3a} /* (9, 26, 6) {real, imag} */,
  {32'hc011b4b2, 32'h3f9c7f4c} /* (9, 26, 5) {real, imag} */,
  {32'hbfd409f7, 32'hbe5963c0} /* (9, 26, 4) {real, imag} */,
  {32'hbf83d48c, 32'hbf82c30a} /* (9, 26, 3) {real, imag} */,
  {32'hbf985573, 32'h3e869440} /* (9, 26, 2) {real, imag} */,
  {32'hbfe95bdf, 32'h3fc7d06c} /* (9, 26, 1) {real, imag} */,
  {32'h3e9e3bb8, 32'h3eb415f3} /* (9, 26, 0) {real, imag} */,
  {32'hbe3cf7c2, 32'h3fce30f4} /* (9, 25, 31) {real, imag} */,
  {32'hbf933863, 32'h3faeba12} /* (9, 25, 30) {real, imag} */,
  {32'hbfd18d76, 32'h3ebe0ce4} /* (9, 25, 29) {real, imag} */,
  {32'hbe735b9c, 32'hbfc61194} /* (9, 25, 28) {real, imag} */,
  {32'hbf3501a0, 32'hbf1531d7} /* (9, 25, 27) {real, imag} */,
  {32'hc00d46ec, 32'h3fa6129b} /* (9, 25, 26) {real, imag} */,
  {32'h3c560400, 32'h3f8afe26} /* (9, 25, 25) {real, imag} */,
  {32'hbc9e20e0, 32'h400214f6} /* (9, 25, 24) {real, imag} */,
  {32'h3f9811b2, 32'h401bb173} /* (9, 25, 23) {real, imag} */,
  {32'h3fc5bf81, 32'h402e53ee} /* (9, 25, 22) {real, imag} */,
  {32'hbea4cc96, 32'h401a2c8a} /* (9, 25, 21) {real, imag} */,
  {32'h3fbd5ab4, 32'hbde57110} /* (9, 25, 20) {real, imag} */,
  {32'h3feb9952, 32'hbf8125ce} /* (9, 25, 19) {real, imag} */,
  {32'h3f3cca70, 32'hbdbd97b0} /* (9, 25, 18) {real, imag} */,
  {32'hbe847d28, 32'hbee2b51c} /* (9, 25, 17) {real, imag} */,
  {32'h3f894d80, 32'hbec5e7b0} /* (9, 25, 16) {real, imag} */,
  {32'h3f84f6aa, 32'h3f1dc7b6} /* (9, 25, 15) {real, imag} */,
  {32'h3e1ceb3c, 32'h3fba0190} /* (9, 25, 14) {real, imag} */,
  {32'hbe020700, 32'hbdd57f88} /* (9, 25, 13) {real, imag} */,
  {32'h3e1a3130, 32'hbf44a2da} /* (9, 25, 12) {real, imag} */,
  {32'h3ebd28f7, 32'h3e1d331c} /* (9, 25, 11) {real, imag} */,
  {32'hbfa3204f, 32'h3ed4d3d4} /* (9, 25, 10) {real, imag} */,
  {32'hc024d0f2, 32'h3f913e82} /* (9, 25, 9) {real, imag} */,
  {32'hc022cc3f, 32'h40095c2f} /* (9, 25, 8) {real, imag} */,
  {32'hbf09938d, 32'h3ec53637} /* (9, 25, 7) {real, imag} */,
  {32'hbe8e6840, 32'h3e95e3cc} /* (9, 25, 6) {real, imag} */,
  {32'hc00f1ab7, 32'h3fc4985a} /* (9, 25, 5) {real, imag} */,
  {32'hbfcedde4, 32'hbe3d47cc} /* (9, 25, 4) {real, imag} */,
  {32'hbe901054, 32'hbf349956} /* (9, 25, 3) {real, imag} */,
  {32'hbf32fdf6, 32'h3e7ca398} /* (9, 25, 2) {real, imag} */,
  {32'hbfbc00bc, 32'h3f57df52} /* (9, 25, 1) {real, imag} */,
  {32'hbf0d6274, 32'hbd6f5510} /* (9, 25, 0) {real, imag} */,
  {32'h3dd98002, 32'h3f2fceba} /* (9, 24, 31) {real, imag} */,
  {32'hc01363e1, 32'h3f7c8ebe} /* (9, 24, 30) {real, imag} */,
  {32'hc03abea4, 32'h3f5f4660} /* (9, 24, 29) {real, imag} */,
  {32'hbf2e9a2e, 32'hbf3d1ba8} /* (9, 24, 28) {real, imag} */,
  {32'h3fcd4eb6, 32'h3f7078f9} /* (9, 24, 27) {real, imag} */,
  {32'hbf649da9, 32'h3f26cc5d} /* (9, 24, 26) {real, imag} */,
  {32'h3f40da37, 32'h3e3e66a6} /* (9, 24, 25) {real, imag} */,
  {32'h3fac3b4d, 32'h3f97b012} /* (9, 24, 24) {real, imag} */,
  {32'h400b5806, 32'h401bce7c} /* (9, 24, 23) {real, imag} */,
  {32'h3fa6c2a9, 32'h3fcec392} /* (9, 24, 22) {real, imag} */,
  {32'hbec83429, 32'h3f6608b9} /* (9, 24, 21) {real, imag} */,
  {32'h3fafc3ec, 32'hbf1c5db1} /* (9, 24, 20) {real, imag} */,
  {32'h3fc4fe21, 32'hbf75a262} /* (9, 24, 19) {real, imag} */,
  {32'hbf2c7abe, 32'hbf311270} /* (9, 24, 18) {real, imag} */,
  {32'hc01b8e28, 32'hbf13ef4c} /* (9, 24, 17) {real, imag} */,
  {32'h3da8f428, 32'hbfa27fe8} /* (9, 24, 16) {real, imag} */,
  {32'h3f7b25b1, 32'hbfba7e78} /* (9, 24, 15) {real, imag} */,
  {32'h3eca540f, 32'hbfa41b21} /* (9, 24, 14) {real, imag} */,
  {32'hbba54c00, 32'hbf4ed846} /* (9, 24, 13) {real, imag} */,
  {32'h3ef04b68, 32'hbf5ccfdd} /* (9, 24, 12) {real, imag} */,
  {32'h3f5fbf88, 32'hbf64c86d} /* (9, 24, 11) {real, imag} */,
  {32'hbf913dba, 32'h3f0a7d54} /* (9, 24, 10) {real, imag} */,
  {32'h3ea7d256, 32'h3e827b40} /* (9, 24, 9) {real, imag} */,
  {32'h3de0e258, 32'h400e1a41} /* (9, 24, 8) {real, imag} */,
  {32'h3f945d04, 32'h3ed34000} /* (9, 24, 7) {real, imag} */,
  {32'h3f62a4ac, 32'hbf34b55a} /* (9, 24, 6) {real, imag} */,
  {32'hbd693000, 32'h3fa1ebc6} /* (9, 24, 5) {real, imag} */,
  {32'h3d2839e0, 32'h3f17ba7e} /* (9, 24, 4) {real, imag} */,
  {32'h3fdbba41, 32'hbfe282b6} /* (9, 24, 3) {real, imag} */,
  {32'h3f5c6f5d, 32'hbf56af58} /* (9, 24, 2) {real, imag} */,
  {32'hbf97fd6a, 32'hbf58ac1a} /* (9, 24, 1) {real, imag} */,
  {32'hbfa07ba2, 32'h3e0c4674} /* (9, 24, 0) {real, imag} */,
  {32'hbb9b2480, 32'h3f57acc5} /* (9, 23, 31) {real, imag} */,
  {32'hc0314a51, 32'h3f6db760} /* (9, 23, 30) {real, imag} */,
  {32'hc0331164, 32'hbe746688} /* (9, 23, 29) {real, imag} */,
  {32'hbfe726de, 32'h3ed39cea} /* (9, 23, 28) {real, imag} */,
  {32'h3f0afdc4, 32'h3facf223} /* (9, 23, 27) {real, imag} */,
  {32'h3f88c74e, 32'h3fbb4d82} /* (9, 23, 26) {real, imag} */,
  {32'h3f3b334c, 32'h3fde8eac} /* (9, 23, 25) {real, imag} */,
  {32'h3e4fa6fc, 32'h40152209} /* (9, 23, 24) {real, imag} */,
  {32'hbf474b1a, 32'h403492b2} /* (9, 23, 23) {real, imag} */,
  {32'hbf201cb6, 32'h3fe9f990} /* (9, 23, 22) {real, imag} */,
  {32'h3fd26a36, 32'h3f398134} /* (9, 23, 21) {real, imag} */,
  {32'h3f94fce1, 32'hbf6596b2} /* (9, 23, 20) {real, imag} */,
  {32'hbfa7a7e0, 32'hbf8777d9} /* (9, 23, 19) {real, imag} */,
  {32'hbfe900c4, 32'hbfb29535} /* (9, 23, 18) {real, imag} */,
  {32'hbfbc0fee, 32'hbfcbffee} /* (9, 23, 17) {real, imag} */,
  {32'hbe8d9bea, 32'hbfc854f7} /* (9, 23, 16) {real, imag} */,
  {32'h3f120b66, 32'hbfff6bdb} /* (9, 23, 15) {real, imag} */,
  {32'h3f26565e, 32'hbf52ab96} /* (9, 23, 14) {real, imag} */,
  {32'h3e5dbf9c, 32'h3fa053d9} /* (9, 23, 13) {real, imag} */,
  {32'h3f1b9a45, 32'h3f5a0560} /* (9, 23, 12) {real, imag} */,
  {32'h3f8d477a, 32'hbf1acd20} /* (9, 23, 11) {real, imag} */,
  {32'hbebb5bb4, 32'h3dc6d170} /* (9, 23, 10) {real, imag} */,
  {32'h3fb26581, 32'h3ef409f0} /* (9, 23, 9) {real, imag} */,
  {32'h3f878f4e, 32'h3ff3dcc3} /* (9, 23, 8) {real, imag} */,
  {32'h3ecc952c, 32'h3f216d56} /* (9, 23, 7) {real, imag} */,
  {32'h3f9e8efa, 32'h3f508306} /* (9, 23, 6) {real, imag} */,
  {32'h3f94ae4e, 32'hbeb5bec0} /* (9, 23, 5) {real, imag} */,
  {32'hbfabd5ce, 32'h3df435a4} /* (9, 23, 4) {real, imag} */,
  {32'hbfa98592, 32'hbed8691c} /* (9, 23, 3) {real, imag} */,
  {32'hbf39cac9, 32'hbe8d6cfc} /* (9, 23, 2) {real, imag} */,
  {32'hbe4e4da8, 32'h3d877110} /* (9, 23, 1) {real, imag} */,
  {32'hbf0ba168, 32'h3fabb84d} /* (9, 23, 0) {real, imag} */,
  {32'hbe7be3f8, 32'hbe3c6eae} /* (9, 22, 31) {real, imag} */,
  {32'hbfeea250, 32'h3f030e74} /* (9, 22, 30) {real, imag} */,
  {32'hbf369e6e, 32'hbe136760} /* (9, 22, 29) {real, imag} */,
  {32'hbf9543cd, 32'h401409d1} /* (9, 22, 28) {real, imag} */,
  {32'hbe93d7af, 32'h4026396a} /* (9, 22, 27) {real, imag} */,
  {32'hbdea8288, 32'h3ff4ffe3} /* (9, 22, 26) {real, imag} */,
  {32'h3f38490d, 32'h3fd57e80} /* (9, 22, 25) {real, imag} */,
  {32'h3e9c3c03, 32'h3f92b3e8} /* (9, 22, 24) {real, imag} */,
  {32'hc0033c8c, 32'h3fc1f909} /* (9, 22, 23) {real, imag} */,
  {32'hbd9d0370, 32'h3f95cf60} /* (9, 22, 22) {real, imag} */,
  {32'h40049768, 32'h3f1f6042} /* (9, 22, 21) {real, imag} */,
  {32'h3f5c7f72, 32'hbf853cca} /* (9, 22, 20) {real, imag} */,
  {32'hbfd337af, 32'hbf2a24fc} /* (9, 22, 19) {real, imag} */,
  {32'h3f3e72bf, 32'hbf5f7f96} /* (9, 22, 18) {real, imag} */,
  {32'h400981c5, 32'hbf31a8be} /* (9, 22, 17) {real, imag} */,
  {32'hbec19378, 32'hbf00476d} /* (9, 22, 16) {real, imag} */,
  {32'h3e699658, 32'hbf31749a} /* (9, 22, 15) {real, imag} */,
  {32'hbf1ae3c2, 32'h3ec2ed3b} /* (9, 22, 14) {real, imag} */,
  {32'h3edb6864, 32'h3fbe1fde} /* (9, 22, 13) {real, imag} */,
  {32'h3fa5ac99, 32'h3fd61b38} /* (9, 22, 12) {real, imag} */,
  {32'h3dfd9b20, 32'h3f013e5a} /* (9, 22, 11) {real, imag} */,
  {32'hbf061cce, 32'hbc1dbb40} /* (9, 22, 10) {real, imag} */,
  {32'h3ea68484, 32'h3fc63a52} /* (9, 22, 9) {real, imag} */,
  {32'h402bc15c, 32'h3faa5efc} /* (9, 22, 8) {real, imag} */,
  {32'hbe1d8878, 32'h3dfcf050} /* (9, 22, 7) {real, imag} */,
  {32'hbecf0892, 32'h3f9d1c04} /* (9, 22, 6) {real, imag} */,
  {32'hbfa3cd40, 32'hbe590458} /* (9, 22, 5) {real, imag} */,
  {32'hc000b585, 32'hbf3d4b6b} /* (9, 22, 4) {real, imag} */,
  {32'hc01189c6, 32'hbf4d9210} /* (9, 22, 3) {real, imag} */,
  {32'hbf8d2e12, 32'hbe8e0de8} /* (9, 22, 2) {real, imag} */,
  {32'h3e2abb18, 32'hbe84838c} /* (9, 22, 1) {real, imag} */,
  {32'h3e5ee3d6, 32'h3f14231b} /* (9, 22, 0) {real, imag} */,
  {32'h3dcb7498, 32'h3c66f840} /* (9, 21, 31) {real, imag} */,
  {32'hbe8b7f37, 32'h3ea4ec9d} /* (9, 21, 30) {real, imag} */,
  {32'h3ff54dbe, 32'h3f593bfe} /* (9, 21, 29) {real, imag} */,
  {32'h3fb490fa, 32'h3fe8fed6} /* (9, 21, 28) {real, imag} */,
  {32'h3ef68a67, 32'h401a0d77} /* (9, 21, 27) {real, imag} */,
  {32'hbfdb051e, 32'h4014d22a} /* (9, 21, 26) {real, imag} */,
  {32'h3ef79bde, 32'h3fbb4d8c} /* (9, 21, 25) {real, imag} */,
  {32'h3f80ed5c, 32'h3f5c50c2} /* (9, 21, 24) {real, imag} */,
  {32'hbefed22b, 32'h3fc94da1} /* (9, 21, 23) {real, imag} */,
  {32'h3fa38847, 32'h3f949a40} /* (9, 21, 22) {real, imag} */,
  {32'h3fa9aa6f, 32'h3f839cc5} /* (9, 21, 21) {real, imag} */,
  {32'h3f9b275a, 32'h3e2a4154} /* (9, 21, 20) {real, imag} */,
  {32'h3e1c7bc4, 32'h3f32dc12} /* (9, 21, 19) {real, imag} */,
  {32'hbf17dd5c, 32'h3edfd9f0} /* (9, 21, 18) {real, imag} */,
  {32'h3f9c25d6, 32'h3f348521} /* (9, 21, 17) {real, imag} */,
  {32'h3ed69336, 32'h40067598} /* (9, 21, 16) {real, imag} */,
  {32'hbdeedde0, 32'h3f3d6dea} /* (9, 21, 15) {real, imag} */,
  {32'hc00b7bf0, 32'h3f6abd4b} /* (9, 21, 14) {real, imag} */,
  {32'h3f17e6dc, 32'h3f917247} /* (9, 21, 13) {real, imag} */,
  {32'h400615d2, 32'h3e1cc227} /* (9, 21, 12) {real, imag} */,
  {32'h3f93012f, 32'hbf13b565} /* (9, 21, 11) {real, imag} */,
  {32'hbf9a35ea, 32'hbebd0de6} /* (9, 21, 10) {real, imag} */,
  {32'hbff62f12, 32'h4010f021} /* (9, 21, 9) {real, imag} */,
  {32'h3f8191ad, 32'h403741ef} /* (9, 21, 8) {real, imag} */,
  {32'h3ec26816, 32'h3f99b049} /* (9, 21, 7) {real, imag} */,
  {32'hbeb79e4e, 32'h3f544f8a} /* (9, 21, 6) {real, imag} */,
  {32'hbfa12447, 32'h3f886cd9} /* (9, 21, 5) {real, imag} */,
  {32'h3e81c779, 32'hbf36a96c} /* (9, 21, 4) {real, imag} */,
  {32'hbed73586, 32'hbfe41004} /* (9, 21, 3) {real, imag} */,
  {32'hbfa6bdc0, 32'hbf0b6292} /* (9, 21, 2) {real, imag} */,
  {32'hbed8b88b, 32'h3e0958f0} /* (9, 21, 1) {real, imag} */,
  {32'h3f44178a, 32'h3ebd40dc} /* (9, 21, 0) {real, imag} */,
  {32'h3e619da4, 32'hbf6186d3} /* (9, 20, 31) {real, imag} */,
  {32'hbf6227b4, 32'hbe103346} /* (9, 20, 30) {real, imag} */,
  {32'h3f55a71c, 32'hbe4f5b68} /* (9, 20, 29) {real, imag} */,
  {32'h3f61e31f, 32'hbfbbfc52} /* (9, 20, 28) {real, imag} */,
  {32'h3fa76bae, 32'h3da1c388} /* (9, 20, 27) {real, imag} */,
  {32'hbd4d2a00, 32'h3fac30fa} /* (9, 20, 26) {real, imag} */,
  {32'h3ef35b70, 32'hbed1a014} /* (9, 20, 25) {real, imag} */,
  {32'h3f93bce7, 32'hbfa9ef0d} /* (9, 20, 24) {real, imag} */,
  {32'h3f2e8ba6, 32'hbf7f6eac} /* (9, 20, 23) {real, imag} */,
  {32'hbea0c3ba, 32'h3eb28050} /* (9, 20, 22) {real, imag} */,
  {32'h3df55fc0, 32'h3f4440b4} /* (9, 20, 21) {real, imag} */,
  {32'h3eccc3a8, 32'h3ed215b4} /* (9, 20, 20) {real, imag} */,
  {32'h3fda58cf, 32'h3fdc7ae8} /* (9, 20, 19) {real, imag} */,
  {32'hbf09cb76, 32'h400319a6} /* (9, 20, 18) {real, imag} */,
  {32'hbf2a4ee5, 32'h3ed04bfc} /* (9, 20, 17) {real, imag} */,
  {32'h3f41eb58, 32'h3fbf937c} /* (9, 20, 16) {real, imag} */,
  {32'hbf790b53, 32'h3f53e22b} /* (9, 20, 15) {real, imag} */,
  {32'hbff0899e, 32'h3f51620e} /* (9, 20, 14) {real, imag} */,
  {32'hbeeeed47, 32'h3f6aab39} /* (9, 20, 13) {real, imag} */,
  {32'h3ee3bf34, 32'h3ec00c38} /* (9, 20, 12) {real, imag} */,
  {32'h3fcd4406, 32'hbf2dcbe4} /* (9, 20, 11) {real, imag} */,
  {32'h3eb4ac48, 32'hbf1f0070} /* (9, 20, 10) {real, imag} */,
  {32'hbebc7ea8, 32'h3ff01a97} /* (9, 20, 9) {real, imag} */,
  {32'h3f96a434, 32'hbf00d8bc} /* (9, 20, 8) {real, imag} */,
  {32'h40185dca, 32'hbf69e73a} /* (9, 20, 7) {real, imag} */,
  {32'h3f1f0d05, 32'h3f22e990} /* (9, 20, 6) {real, imag} */,
  {32'hbf03b229, 32'h3feaaa8b} /* (9, 20, 5) {real, imag} */,
  {32'h40126759, 32'h3ead5292} /* (9, 20, 4) {real, imag} */,
  {32'h3f4e0224, 32'hc00399e6} /* (9, 20, 3) {real, imag} */,
  {32'hbfc4a0aa, 32'hc01181a4} /* (9, 20, 2) {real, imag} */,
  {32'hbf5e0061, 32'hbfa77e55} /* (9, 20, 1) {real, imag} */,
  {32'h3f5e9c95, 32'hbf5f917c} /* (9, 20, 0) {real, imag} */,
  {32'hbe17b3ce, 32'hbfea7a84} /* (9, 19, 31) {real, imag} */,
  {32'h3e885714, 32'hbf9203ee} /* (9, 19, 30) {real, imag} */,
  {32'h3f333d62, 32'h3f8ae1bc} /* (9, 19, 29) {real, imag} */,
  {32'hbef8ce7c, 32'hbf77cfdf} /* (9, 19, 28) {real, imag} */,
  {32'h3eec9318, 32'hbfbac2e6} /* (9, 19, 27) {real, imag} */,
  {32'h3f14f559, 32'hbd048510} /* (9, 19, 26) {real, imag} */,
  {32'h3f58a6aa, 32'hbd9dd900} /* (9, 19, 25) {real, imag} */,
  {32'h3f908d86, 32'hc001dfea} /* (9, 19, 24) {real, imag} */,
  {32'hbe24b8a8, 32'hc004bd9e} /* (9, 19, 23) {real, imag} */,
  {32'hc00105aa, 32'hbf9fa25e} /* (9, 19, 22) {real, imag} */,
  {32'hbd5b8800, 32'hbef55b54} /* (9, 19, 21) {real, imag} */,
  {32'hbe3b9338, 32'hbf7fe115} /* (9, 19, 20) {real, imag} */,
  {32'h3fb234bc, 32'h3f47789a} /* (9, 19, 19) {real, imag} */,
  {32'h3e7bfe4c, 32'h3fde67e0} /* (9, 19, 18) {real, imag} */,
  {32'hbf2d96d0, 32'h3f810204} /* (9, 19, 17) {real, imag} */,
  {32'h3f3c2169, 32'h3f5dc8c0} /* (9, 19, 16) {real, imag} */,
  {32'hbecea625, 32'hbe8df80d} /* (9, 19, 15) {real, imag} */,
  {32'hbf6e855c, 32'h3e105082} /* (9, 19, 14) {real, imag} */,
  {32'hbf14ab0d, 32'h3e9e1391} /* (9, 19, 13) {real, imag} */,
  {32'hbfdc5f56, 32'h3f85886c} /* (9, 19, 12) {real, imag} */,
  {32'hbf6fd08d, 32'hbeb222bc} /* (9, 19, 11) {real, imag} */,
  {32'h3ea7c92a, 32'h3f901d6a} /* (9, 19, 10) {real, imag} */,
  {32'h3fa8eb68, 32'h40209fc7} /* (9, 19, 9) {real, imag} */,
  {32'h40182cbe, 32'hbe7c6ea8} /* (9, 19, 8) {real, imag} */,
  {32'h4053146f, 32'hbfb5a884} /* (9, 19, 7) {real, imag} */,
  {32'h3fe0cd09, 32'hbecf4e7a} /* (9, 19, 6) {real, imag} */,
  {32'h3ea76292, 32'hbf41891e} /* (9, 19, 5) {real, imag} */,
  {32'h3f4926a6, 32'hbed2afe5} /* (9, 19, 4) {real, imag} */,
  {32'h3f9a9746, 32'hbf98c440} /* (9, 19, 3) {real, imag} */,
  {32'hbe2a9e3c, 32'hbf35e45f} /* (9, 19, 2) {real, imag} */,
  {32'hbfcf38c4, 32'hbf4da4f5} /* (9, 19, 1) {real, imag} */,
  {32'hbf8d568e, 32'hbfa76c57} /* (9, 19, 0) {real, imag} */,
  {32'h3f55a572, 32'hbf77edc8} /* (9, 18, 31) {real, imag} */,
  {32'h3f2e38fc, 32'hbf33be1c} /* (9, 18, 30) {real, imag} */,
  {32'h3f59aac8, 32'h400a7616} /* (9, 18, 29) {real, imag} */,
  {32'h3e917174, 32'h3fd3dbb3} /* (9, 18, 28) {real, imag} */,
  {32'h3d211b80, 32'h3e146204} /* (9, 18, 27) {real, imag} */,
  {32'hbefe60f8, 32'hbea6998e} /* (9, 18, 26) {real, imag} */,
  {32'hbd117740, 32'hbf87d990} /* (9, 18, 25) {real, imag} */,
  {32'h3fc35e27, 32'hc003a050} /* (9, 18, 24) {real, imag} */,
  {32'h3e309378, 32'h3f2f42a8} /* (9, 18, 23) {real, imag} */,
  {32'hbfde22b1, 32'h3f55a610} /* (9, 18, 22) {real, imag} */,
  {32'hbfc26b2c, 32'h3e671ce8} /* (9, 18, 21) {real, imag} */,
  {32'hbf5795c6, 32'hbf805700} /* (9, 18, 20) {real, imag} */,
  {32'h3f567150, 32'hbf297c6a} /* (9, 18, 19) {real, imag} */,
  {32'h3e66f2a0, 32'hbf993d5a} /* (9, 18, 18) {real, imag} */,
  {32'hbebb8f58, 32'hbf2604fc} /* (9, 18, 17) {real, imag} */,
  {32'h3f8b6b82, 32'h3fe5ca5a} /* (9, 18, 16) {real, imag} */,
  {32'h3dcbe360, 32'h3f7fb3aa} /* (9, 18, 15) {real, imag} */,
  {32'hbeddf2e6, 32'h3fd87a85} /* (9, 18, 14) {real, imag} */,
  {32'hbfe777df, 32'h40585b86} /* (9, 18, 13) {real, imag} */,
  {32'hc042d884, 32'h400e7b1e} /* (9, 18, 12) {real, imag} */,
  {32'hc02ea6e8, 32'h3eae5fb6} /* (9, 18, 11) {real, imag} */,
  {32'hbf9822ce, 32'h3fd0503e} /* (9, 18, 10) {real, imag} */,
  {32'h3fc332c4, 32'h3f7ff242} /* (9, 18, 9) {real, imag} */,
  {32'h3ff9892a, 32'hbf9698ca} /* (9, 18, 8) {real, imag} */,
  {32'h3fc4eeb0, 32'hc0138b0d} /* (9, 18, 7) {real, imag} */,
  {32'h3f94557a, 32'hc01e0220} /* (9, 18, 6) {real, imag} */,
  {32'hbd93c4e0, 32'hc00c0e82} /* (9, 18, 5) {real, imag} */,
  {32'hbf52501e, 32'hbfaccbfd} /* (9, 18, 4) {real, imag} */,
  {32'h3efcf6f0, 32'h3f0d28ae} /* (9, 18, 3) {real, imag} */,
  {32'h3f289045, 32'h3f8d1c43} /* (9, 18, 2) {real, imag} */,
  {32'hc010969e, 32'h3ed32c98} /* (9, 18, 1) {real, imag} */,
  {32'hc01be1d2, 32'h3ea7c69a} /* (9, 18, 0) {real, imag} */,
  {32'h3dfba898, 32'h3eb7aa40} /* (9, 17, 31) {real, imag} */,
  {32'h3f92078c, 32'h3f882eab} /* (9, 17, 30) {real, imag} */,
  {32'h402278a4, 32'h3efa73a6} /* (9, 17, 29) {real, imag} */,
  {32'h4022a5d5, 32'h3ffc88c3} /* (9, 17, 28) {real, imag} */,
  {32'h3f998c9e, 32'h3f680c48} /* (9, 17, 27) {real, imag} */,
  {32'hbef1820c, 32'hbf86ea06} /* (9, 17, 26) {real, imag} */,
  {32'hbf7f33f2, 32'hc01b459a} /* (9, 17, 25) {real, imag} */,
  {32'h3f924e17, 32'hbfc30ab6} /* (9, 17, 24) {real, imag} */,
  {32'h3f6f7d18, 32'hbe7468d8} /* (9, 17, 23) {real, imag} */,
  {32'hbf951849, 32'hbf80319f} /* (9, 17, 22) {real, imag} */,
  {32'hc002dbbd, 32'h3e9fd770} /* (9, 17, 21) {real, imag} */,
  {32'hc014469a, 32'h3f1fe3e8} /* (9, 17, 20) {real, imag} */,
  {32'hbed53966, 32'h3f11e6f5} /* (9, 17, 19) {real, imag} */,
  {32'h3f301932, 32'h3d67a500} /* (9, 17, 18) {real, imag} */,
  {32'hbf7b8456, 32'hbf56c116} /* (9, 17, 17) {real, imag} */,
  {32'hbdf88810, 32'h3e89d73e} /* (9, 17, 16) {real, imag} */,
  {32'h3eb66d96, 32'h3f2ef9a6} /* (9, 17, 15) {real, imag} */,
  {32'h3f6d6220, 32'h3f35da58} /* (9, 17, 14) {real, imag} */,
  {32'hbfa17d5d, 32'h4018a46c} /* (9, 17, 13) {real, imag} */,
  {32'hc00f998d, 32'h4066c3c0} /* (9, 17, 12) {real, imag} */,
  {32'hbfdc1f47, 32'h3feca30e} /* (9, 17, 11) {real, imag} */,
  {32'h3e987e68, 32'hbe85a894} /* (9, 17, 10) {real, imag} */,
  {32'h3fad46c0, 32'hc004d55d} /* (9, 17, 9) {real, imag} */,
  {32'h3ec7be78, 32'hc0141810} /* (9, 17, 8) {real, imag} */,
  {32'h3e3bcb06, 32'hc0354e7e} /* (9, 17, 7) {real, imag} */,
  {32'hbeb92b78, 32'hc080024c} /* (9, 17, 6) {real, imag} */,
  {32'h3eaa9ebe, 32'hbf9d6fad} /* (9, 17, 5) {real, imag} */,
  {32'hbec4f97d, 32'h3e92a8c9} /* (9, 17, 4) {real, imag} */,
  {32'hbb7bd000, 32'h3fbef7b4} /* (9, 17, 3) {real, imag} */,
  {32'h3ee98bc5, 32'h3ea2263a} /* (9, 17, 2) {real, imag} */,
  {32'hbfa863ba, 32'h3e563ec8} /* (9, 17, 1) {real, imag} */,
  {32'hbfb61712, 32'h3f84f17c} /* (9, 17, 0) {real, imag} */,
  {32'h3dbf003c, 32'h3fc98f82} /* (9, 16, 31) {real, imag} */,
  {32'h40076c81, 32'h3fe41b2f} /* (9, 16, 30) {real, imag} */,
  {32'h4048aa28, 32'hbf8dd590} /* (9, 16, 29) {real, imag} */,
  {32'h3f7dcce8, 32'hbf9c65c0} /* (9, 16, 28) {real, imag} */,
  {32'hbde012bc, 32'hbf7e3bee} /* (9, 16, 27) {real, imag} */,
  {32'h3f3cdacc, 32'hbfdb28f6} /* (9, 16, 26) {real, imag} */,
  {32'h3ecf4da4, 32'hbfeebae1} /* (9, 16, 25) {real, imag} */,
  {32'h3d8897f0, 32'hbf1d25e7} /* (9, 16, 24) {real, imag} */,
  {32'h3ce87df0, 32'hc0153304} /* (9, 16, 23) {real, imag} */,
  {32'hbdf98b30, 32'hc01abcd6} /* (9, 16, 22) {real, imag} */,
  {32'hbf55166c, 32'hbed070e2} /* (9, 16, 21) {real, imag} */,
  {32'hc000b2b4, 32'h3d657400} /* (9, 16, 20) {real, imag} */,
  {32'hbfe12499, 32'hbf12c3da} /* (9, 16, 19) {real, imag} */,
  {32'hbe0a9e1c, 32'h3f2e9b3c} /* (9, 16, 18) {real, imag} */,
  {32'h3ef35250, 32'h3f9caee6} /* (9, 16, 17) {real, imag} */,
  {32'h3f2e7963, 32'h3fd236ae} /* (9, 16, 16) {real, imag} */,
  {32'hbf5870a6, 32'h3fa2417a} /* (9, 16, 15) {real, imag} */,
  {32'hbee8197a, 32'hbf1dc990} /* (9, 16, 14) {real, imag} */,
  {32'hc01442f4, 32'hbf9361f4} /* (9, 16, 13) {real, imag} */,
  {32'hc0269b82, 32'h3f19417f} /* (9, 16, 12) {real, imag} */,
  {32'h3e17ac40, 32'h4002168c} /* (9, 16, 11) {real, imag} */,
  {32'h3f9f38ea, 32'h3f173a95} /* (9, 16, 10) {real, imag} */,
  {32'h3f9943aa, 32'hbfbd0efa} /* (9, 16, 9) {real, imag} */,
  {32'hbf17e280, 32'hc00d4b5a} /* (9, 16, 8) {real, imag} */,
  {32'hbce2af30, 32'hc039cbea} /* (9, 16, 7) {real, imag} */,
  {32'h3fb6ca36, 32'hc03d8e8a} /* (9, 16, 6) {real, imag} */,
  {32'h3f8feaac, 32'h3eacc34c} /* (9, 16, 5) {real, imag} */,
  {32'h3fa57aa9, 32'h3f2bc0ac} /* (9, 16, 4) {real, imag} */,
  {32'h3f943e36, 32'h4007f5c8} /* (9, 16, 3) {real, imag} */,
  {32'hbf1ffc5c, 32'h3f2a6292} /* (9, 16, 2) {real, imag} */,
  {32'h3f450ef2, 32'hbf353e24} /* (9, 16, 1) {real, imag} */,
  {32'h3f754d30, 32'h3f3f21ce} /* (9, 16, 0) {real, imag} */,
  {32'h3e0d1d0c, 32'h3f87d2aa} /* (9, 15, 31) {real, imag} */,
  {32'h3f4d0d44, 32'h3f91484a} /* (9, 15, 30) {real, imag} */,
  {32'h3f8c1687, 32'hbf6290f6} /* (9, 15, 29) {real, imag} */,
  {32'h3f86f330, 32'hc036053e} /* (9, 15, 28) {real, imag} */,
  {32'h3e678cd0, 32'hc00e35a6} /* (9, 15, 27) {real, imag} */,
  {32'hbf16517e, 32'hbfaca61e} /* (9, 15, 26) {real, imag} */,
  {32'h3f76349c, 32'hbebadf9c} /* (9, 15, 25) {real, imag} */,
  {32'hbe7e8164, 32'hbfd54622} /* (9, 15, 24) {real, imag} */,
  {32'hbf097bb6, 32'hc066305c} /* (9, 15, 23) {real, imag} */,
  {32'h3f72c1ce, 32'hc009b36e} /* (9, 15, 22) {real, imag} */,
  {32'h401c8ce8, 32'hbe525268} /* (9, 15, 21) {real, imag} */,
  {32'h3f84bbcc, 32'h3f8aaa1a} /* (9, 15, 20) {real, imag} */,
  {32'hbe840eac, 32'h3f949ee2} /* (9, 15, 19) {real, imag} */,
  {32'hbf1fc523, 32'h3f4c2cca} /* (9, 15, 18) {real, imag} */,
  {32'h3ee52e4c, 32'h3f987bc6} /* (9, 15, 17) {real, imag} */,
  {32'h3f8a54fc, 32'h3f9cc526} /* (9, 15, 16) {real, imag} */,
  {32'hbe42c4a0, 32'h3faf6b93} /* (9, 15, 15) {real, imag} */,
  {32'hbf48a430, 32'hbde69870} /* (9, 15, 14) {real, imag} */,
  {32'hbf429092, 32'h3e460032} /* (9, 15, 13) {real, imag} */,
  {32'hbfa0af4d, 32'hbe8c0a74} /* (9, 15, 12) {real, imag} */,
  {32'hbf2dc800, 32'h3fb06d29} /* (9, 15, 11) {real, imag} */,
  {32'h3f5697c5, 32'h3fde3032} /* (9, 15, 10) {real, imag} */,
  {32'h3e054630, 32'hbec7bed4} /* (9, 15, 9) {real, imag} */,
  {32'hbf8f6d82, 32'hbff94714} /* (9, 15, 8) {real, imag} */,
  {32'hbf8aad03, 32'hbfbd95a2} /* (9, 15, 7) {real, imag} */,
  {32'h3e993eb0, 32'hbfaf54b6} /* (9, 15, 6) {real, imag} */,
  {32'h3f1b6f5b, 32'h3f61a9ba} /* (9, 15, 5) {real, imag} */,
  {32'h3fd7b25e, 32'hbe01e920} /* (9, 15, 4) {real, imag} */,
  {32'h3f104706, 32'h3fb12fde} /* (9, 15, 3) {real, imag} */,
  {32'hbf01d0c0, 32'h3ecb5d26} /* (9, 15, 2) {real, imag} */,
  {32'h3fc55dcb, 32'hc03eb2b0} /* (9, 15, 1) {real, imag} */,
  {32'h3fe2683b, 32'hbefd23e8} /* (9, 15, 0) {real, imag} */,
  {32'h3ecd21e0, 32'h3e20d218} /* (9, 14, 31) {real, imag} */,
  {32'h3f1bcdc7, 32'h3eded44c} /* (9, 14, 30) {real, imag} */,
  {32'hbe3c79bb, 32'h3f787228} /* (9, 14, 29) {real, imag} */,
  {32'h3f981aa8, 32'hbec62d71} /* (9, 14, 28) {real, imag} */,
  {32'h3ffd15be, 32'hbf2d59be} /* (9, 14, 27) {real, imag} */,
  {32'h3fc34538, 32'hbe91000a} /* (9, 14, 26) {real, imag} */,
  {32'h3fc0ae3e, 32'h3d64a500} /* (9, 14, 25) {real, imag} */,
  {32'hbf658cb5, 32'hbf3f8f5e} /* (9, 14, 24) {real, imag} */,
  {32'hbef04b85, 32'hbef2e131} /* (9, 14, 23) {real, imag} */,
  {32'h3f929dcf, 32'h3fb6b74e} /* (9, 14, 22) {real, imag} */,
  {32'h3fb0181b, 32'h403fbb5d} /* (9, 14, 21) {real, imag} */,
  {32'h3fdccb1e, 32'h3ff8b6e5} /* (9, 14, 20) {real, imag} */,
  {32'h3fdb61fd, 32'h3875c000} /* (9, 14, 19) {real, imag} */,
  {32'hbeecf41e, 32'h3dd8ea40} /* (9, 14, 18) {real, imag} */,
  {32'h3e856892, 32'h3fa224fe} /* (9, 14, 17) {real, imag} */,
  {32'h3bed6580, 32'h3f942d46} /* (9, 14, 16) {real, imag} */,
  {32'hbf149fd2, 32'h3fa74770} /* (9, 14, 15) {real, imag} */,
  {32'h3d3ac340, 32'h3eed0c94} /* (9, 14, 14) {real, imag} */,
  {32'h3efabc46, 32'h3fbd64fe} /* (9, 14, 13) {real, imag} */,
  {32'h3e5ec9c0, 32'hbf2c8146} /* (9, 14, 12) {real, imag} */,
  {32'hbea45688, 32'hbf86df2c} /* (9, 14, 11) {real, imag} */,
  {32'h3eeff4c7, 32'hbf9e246a} /* (9, 14, 10) {real, imag} */,
  {32'hbed26f10, 32'hbf5001c6} /* (9, 14, 9) {real, imag} */,
  {32'hbf48aa4d, 32'hbdf5f2f4} /* (9, 14, 8) {real, imag} */,
  {32'h3f5992b4, 32'hbdd2e550} /* (9, 14, 7) {real, imag} */,
  {32'h3ecbd3c0, 32'h3e08baee} /* (9, 14, 6) {real, imag} */,
  {32'h3f87580d, 32'h3f4b20b4} /* (9, 14, 5) {real, imag} */,
  {32'h3f049962, 32'hbe4e1cae} /* (9, 14, 4) {real, imag} */,
  {32'hbfbff6d1, 32'hbd99ca60} /* (9, 14, 3) {real, imag} */,
  {32'h3f126d97, 32'h3f93ffd1} /* (9, 14, 2) {real, imag} */,
  {32'h40082d60, 32'hbe518420} /* (9, 14, 1) {real, imag} */,
  {32'h3fad86a0, 32'hbd67ccb0} /* (9, 14, 0) {real, imag} */,
  {32'h3ec5737e, 32'h3ec3bb3c} /* (9, 13, 31) {real, imag} */,
  {32'h3f024f28, 32'h3edf09a3} /* (9, 13, 30) {real, imag} */,
  {32'hbf379b88, 32'h3eaa1cbe} /* (9, 13, 29) {real, imag} */,
  {32'hbeba4d48, 32'h3e786eaa} /* (9, 13, 28) {real, imag} */,
  {32'h3eccb8d6, 32'hbf8ddc78} /* (9, 13, 27) {real, imag} */,
  {32'hbe123c70, 32'hbf7266f9} /* (9, 13, 26) {real, imag} */,
  {32'h3f066cbb, 32'h3d907b20} /* (9, 13, 25) {real, imag} */,
  {32'h3efe5b7c, 32'h3fa00838} /* (9, 13, 24) {real, imag} */,
  {32'h3f0def3c, 32'h400bcbe6} /* (9, 13, 23) {real, imag} */,
  {32'h3f97180f, 32'h4028a6dc} /* (9, 13, 22) {real, imag} */,
  {32'h3f2306ce, 32'h4018c1d0} /* (9, 13, 21) {real, imag} */,
  {32'h3fc21184, 32'h404f6486} /* (9, 13, 20) {real, imag} */,
  {32'h3fb423d9, 32'h3f926b66} /* (9, 13, 19) {real, imag} */,
  {32'h3f33d9ba, 32'h3e9069fc} /* (9, 13, 18) {real, imag} */,
  {32'h3abdf400, 32'h40003746} /* (9, 13, 17) {real, imag} */,
  {32'hbf45211a, 32'h3fb72ead} /* (9, 13, 16) {real, imag} */,
  {32'hbda67c7c, 32'h3f5cbf28} /* (9, 13, 15) {real, imag} */,
  {32'h3e54aaba, 32'h3d4f36d0} /* (9, 13, 14) {real, imag} */,
  {32'h3fbe7e3b, 32'h3f6015b4} /* (9, 13, 13) {real, imag} */,
  {32'h3fb6970f, 32'hbe8667c0} /* (9, 13, 12) {real, imag} */,
  {32'h3e3f7308, 32'hbf82b27c} /* (9, 13, 11) {real, imag} */,
  {32'h3f82f87e, 32'hbfcef621} /* (9, 13, 10) {real, imag} */,
  {32'h3ce37b00, 32'hc016982a} /* (9, 13, 9) {real, imag} */,
  {32'h3e6ea888, 32'hbebf90ec} /* (9, 13, 8) {real, imag} */,
  {32'h4066eaac, 32'hbfbfb7f0} /* (9, 13, 7) {real, imag} */,
  {32'h3f99639c, 32'h3d2bc7dc} /* (9, 13, 6) {real, imag} */,
  {32'h3fc4e7c4, 32'h3f8c9d05} /* (9, 13, 5) {real, imag} */,
  {32'h3fe22e11, 32'h3f8dfa44} /* (9, 13, 4) {real, imag} */,
  {32'h3f1b32b0, 32'hbeb75fa8} /* (9, 13, 3) {real, imag} */,
  {32'h3f9caded, 32'h3f140558} /* (9, 13, 2) {real, imag} */,
  {32'h3fdf550c, 32'h3fa95916} /* (9, 13, 1) {real, imag} */,
  {32'h3f9249a4, 32'h3e589f24} /* (9, 13, 0) {real, imag} */,
  {32'h3fa23c3b, 32'h3dab7420} /* (9, 12, 31) {real, imag} */,
  {32'h3f557768, 32'hbf68f2da} /* (9, 12, 30) {real, imag} */,
  {32'hbf8e6fa2, 32'hbfc1c6f2} /* (9, 12, 29) {real, imag} */,
  {32'hbf752812, 32'hbf8e84ff} /* (9, 12, 28) {real, imag} */,
  {32'hbf0fabae, 32'hbea86538} /* (9, 12, 27) {real, imag} */,
  {32'hbf9ca0f1, 32'hbfda8ba7} /* (9, 12, 26) {real, imag} */,
  {32'h3dc0fa80, 32'h3f18df33} /* (9, 12, 25) {real, imag} */,
  {32'h3f08b186, 32'h3f001cb6} /* (9, 12, 24) {real, imag} */,
  {32'h3f150ebd, 32'hbfe32d3f} /* (9, 12, 23) {real, imag} */,
  {32'h3fc7e58a, 32'hbfb3ccf3} /* (9, 12, 22) {real, imag} */,
  {32'hbea6e1f8, 32'hbf8cbaa0} /* (9, 12, 21) {real, imag} */,
  {32'h3eced6a6, 32'h3f822546} /* (9, 12, 20) {real, imag} */,
  {32'h3f31c9de, 32'h3fe6549d} /* (9, 12, 19) {real, imag} */,
  {32'h3f204ff4, 32'hbe4534c0} /* (9, 12, 18) {real, imag} */,
  {32'hbc446280, 32'h3fb1c2a2} /* (9, 12, 17) {real, imag} */,
  {32'hbf48aa14, 32'hbee57300} /* (9, 12, 16) {real, imag} */,
  {32'h3e5b2888, 32'hbfcb1db5} /* (9, 12, 15) {real, imag} */,
  {32'hbe3d5930, 32'h3e145718} /* (9, 12, 14) {real, imag} */,
  {32'h3fb97758, 32'h3f884c6d} /* (9, 12, 13) {real, imag} */,
  {32'h3ff21250, 32'h3ff73cb5} /* (9, 12, 12) {real, imag} */,
  {32'h3ec31498, 32'h3d7a3440} /* (9, 12, 11) {real, imag} */,
  {32'h4003760e, 32'hbf27573d} /* (9, 12, 10) {real, imag} */,
  {32'h3f95dd70, 32'h3ef2ba02} /* (9, 12, 9) {real, imag} */,
  {32'hbe22f2d8, 32'h3f3520f0} /* (9, 12, 8) {real, imag} */,
  {32'h40270a56, 32'hbf9d0af2} /* (9, 12, 7) {real, imag} */,
  {32'h40109458, 32'hbf77c310} /* (9, 12, 6) {real, imag} */,
  {32'h40069107, 32'hbef4ab82} /* (9, 12, 5) {real, imag} */,
  {32'h3f8366c6, 32'h3eedc1d7} /* (9, 12, 4) {real, imag} */,
  {32'hbe3fbf34, 32'h3f8dd542} /* (9, 12, 3) {real, imag} */,
  {32'hbfcf3bc9, 32'h3f3cdc77} /* (9, 12, 2) {real, imag} */,
  {32'hbf5e9403, 32'h3fb79692} /* (9, 12, 1) {real, imag} */,
  {32'h3e9733fd, 32'h3e943874} /* (9, 12, 0) {real, imag} */,
  {32'hbd911e38, 32'h3c941a80} /* (9, 11, 31) {real, imag} */,
  {32'hbf5e98a4, 32'h3e1a179c} /* (9, 11, 30) {real, imag} */,
  {32'hbfb61d2b, 32'hbcd27898} /* (9, 11, 29) {real, imag} */,
  {32'hbfa10f62, 32'hbf91fa42} /* (9, 11, 28) {real, imag} */,
  {32'hc00c2bae, 32'hbf7df227} /* (9, 11, 27) {real, imag} */,
  {32'hbff0b211, 32'hbfc9b9e0} /* (9, 11, 26) {real, imag} */,
  {32'hbe4f2c0a, 32'h3e9f25b2} /* (9, 11, 25) {real, imag} */,
  {32'h3df0dc18, 32'h3f1e4802} /* (9, 11, 24) {real, imag} */,
  {32'h3da7bb40, 32'hbe64e6ac} /* (9, 11, 23) {real, imag} */,
  {32'h3f9f7e65, 32'hbfdba72c} /* (9, 11, 22) {real, imag} */,
  {32'hbf0bffb2, 32'hbfa9df96} /* (9, 11, 21) {real, imag} */,
  {32'hbf843dc7, 32'hbf221f27} /* (9, 11, 20) {real, imag} */,
  {32'h3f38de53, 32'hbf5cc52a} /* (9, 11, 19) {real, imag} */,
  {32'hbf898b4d, 32'h3c245700} /* (9, 11, 18) {real, imag} */,
  {32'hbff6fcac, 32'h400aa00a} /* (9, 11, 17) {real, imag} */,
  {32'h3d7b7770, 32'hbf9066e4} /* (9, 11, 16) {real, imag} */,
  {32'h3e033b02, 32'hbf5e5684} /* (9, 11, 15) {real, imag} */,
  {32'hbfa5e907, 32'h4020c0ec} /* (9, 11, 14) {real, imag} */,
  {32'h3f90e368, 32'h402dba98} /* (9, 11, 13) {real, imag} */,
  {32'h40331ca2, 32'h4014372c} /* (9, 11, 12) {real, imag} */,
  {32'h3f96ac68, 32'hbeb4d0f4} /* (9, 11, 11) {real, imag} */,
  {32'h3fe20aa4, 32'hbf679c66} /* (9, 11, 10) {real, imag} */,
  {32'h3fd1dcbe, 32'h4025ada3} /* (9, 11, 9) {real, imag} */,
  {32'hbd4d38a0, 32'h3f8416be} /* (9, 11, 8) {real, imag} */,
  {32'h3f5c84a8, 32'h3e9bb48e} /* (9, 11, 7) {real, imag} */,
  {32'h3f8cb68f, 32'h3dd3a840} /* (9, 11, 6) {real, imag} */,
  {32'h3fb93dcd, 32'hbe1d74c0} /* (9, 11, 5) {real, imag} */,
  {32'h3d42bdd8, 32'hbf13e48e} /* (9, 11, 4) {real, imag} */,
  {32'hbe237afc, 32'h3ef92bde} /* (9, 11, 3) {real, imag} */,
  {32'h3e8b944c, 32'h3ed7fe08} /* (9, 11, 2) {real, imag} */,
  {32'h3ece6311, 32'h3f7e36f6} /* (9, 11, 1) {real, imag} */,
  {32'hbeb03ca2, 32'h3ea180aa} /* (9, 11, 0) {real, imag} */,
  {32'h3d868afe, 32'h3f8871ca} /* (9, 10, 31) {real, imag} */,
  {32'hbfab76da, 32'h3e21e3e4} /* (9, 10, 30) {real, imag} */,
  {32'hbf892121, 32'h3f44ddb8} /* (9, 10, 29) {real, imag} */,
  {32'hbf8c5e8f, 32'h3f24f2f4} /* (9, 10, 28) {real, imag} */,
  {32'hc010d618, 32'hbf8bcd60} /* (9, 10, 27) {real, imag} */,
  {32'hbfd57668, 32'hbf8aeb20} /* (9, 10, 26) {real, imag} */,
  {32'hbf84f6a1, 32'h3fa63364} /* (9, 10, 25) {real, imag} */,
  {32'hbe3e15cf, 32'h403b49c8} /* (9, 10, 24) {real, imag} */,
  {32'hbebd6174, 32'h40284d40} /* (9, 10, 23) {real, imag} */,
  {32'h3eb465aa, 32'h3edbe9c0} /* (9, 10, 22) {real, imag} */,
  {32'h3f482e9a, 32'h3fa43926} /* (9, 10, 21) {real, imag} */,
  {32'h3f1af997, 32'hbfa482c7} /* (9, 10, 20) {real, imag} */,
  {32'h3ed270cf, 32'hc040a3b3} /* (9, 10, 19) {real, imag} */,
  {32'hbfa2cd55, 32'hbee66ed4} /* (9, 10, 18) {real, imag} */,
  {32'hc00b290a, 32'h3f837aee} /* (9, 10, 17) {real, imag} */,
  {32'hbf793473, 32'hbf8abef4} /* (9, 10, 16) {real, imag} */,
  {32'hbfec87db, 32'hbe1d0a08} /* (9, 10, 15) {real, imag} */,
  {32'hbef4dd7c, 32'h3fc65ae2} /* (9, 10, 14) {real, imag} */,
  {32'h3f29cfad, 32'h400368d2} /* (9, 10, 13) {real, imag} */,
  {32'h3fba6180, 32'h3f12c936} /* (9, 10, 12) {real, imag} */,
  {32'h3febc550, 32'hbfdbba3c} /* (9, 10, 11) {real, imag} */,
  {32'h3f46c331, 32'h3f0157bf} /* (9, 10, 10) {real, imag} */,
  {32'hbeb9a1fc, 32'h40293968} /* (9, 10, 9) {real, imag} */,
  {32'hbf9c5110, 32'h3f5a3eb8} /* (9, 10, 8) {real, imag} */,
  {32'hbf9f428b, 32'h3fec2bfe} /* (9, 10, 7) {real, imag} */,
  {32'hbf796d32, 32'h3f5721db} /* (9, 10, 6) {real, imag} */,
  {32'hbf8e6684, 32'h3f017cb4} /* (9, 10, 5) {real, imag} */,
  {32'hbf55e854, 32'hbe1637e8} /* (9, 10, 4) {real, imag} */,
  {32'h3fa8496b, 32'hbfc45a7c} /* (9, 10, 3) {real, imag} */,
  {32'h40404cee, 32'hbf8b5240} /* (9, 10, 2) {real, imag} */,
  {32'h3f83fb27, 32'hbf7ddbf8} /* (9, 10, 1) {real, imag} */,
  {32'hbf0277df, 32'hbf8e76c6} /* (9, 10, 0) {real, imag} */,
  {32'h3f81c7f7, 32'h3f2f54f5} /* (9, 9, 31) {real, imag} */,
  {32'h3e9c791e, 32'h3f3bfb3f} /* (9, 9, 30) {real, imag} */,
  {32'hbecb7e60, 32'h3db63c40} /* (9, 9, 29) {real, imag} */,
  {32'hbf27b678, 32'h3f0907aa} /* (9, 9, 28) {real, imag} */,
  {32'hbf818760, 32'h3f23a226} /* (9, 9, 27) {real, imag} */,
  {32'hbf402404, 32'hbddfbd4c} /* (9, 9, 26) {real, imag} */,
  {32'h3e7e1650, 32'h40089f2e} /* (9, 9, 25) {real, imag} */,
  {32'h3e63970c, 32'h4045e570} /* (9, 9, 24) {real, imag} */,
  {32'h3f3de571, 32'h4022eda2} /* (9, 9, 23) {real, imag} */,
  {32'h3fd67d13, 32'h401f655e} /* (9, 9, 22) {real, imag} */,
  {32'h3f5ceb73, 32'h3ff13456} /* (9, 9, 21) {real, imag} */,
  {32'h3f87cb32, 32'hbfc1d47e} /* (9, 9, 20) {real, imag} */,
  {32'h3e1a92b0, 32'hc000e6f8} /* (9, 9, 19) {real, imag} */,
  {32'h3e6cc290, 32'hc01d5cb2} /* (9, 9, 18) {real, imag} */,
  {32'hbe2f9f38, 32'hc032d80a} /* (9, 9, 17) {real, imag} */,
  {32'h3d774ca0, 32'hbfee9134} /* (9, 9, 16) {real, imag} */,
  {32'hbffd2d78, 32'h3e7b1680} /* (9, 9, 15) {real, imag} */,
  {32'h3fbf0b22, 32'h3fc53423} /* (9, 9, 14) {real, imag} */,
  {32'h3fdd933d, 32'h401a84d5} /* (9, 9, 13) {real, imag} */,
  {32'h3fbb65e3, 32'h3f898329} /* (9, 9, 12) {real, imag} */,
  {32'h3fca5a08, 32'hc003f5d7} /* (9, 9, 11) {real, imag} */,
  {32'h3f933fcf, 32'h3f8816f5} /* (9, 9, 10) {real, imag} */,
  {32'hbf120564, 32'h4034ef24} /* (9, 9, 9) {real, imag} */,
  {32'hbf1df328, 32'h3fb6713d} /* (9, 9, 8) {real, imag} */,
  {32'hbf4ca7c8, 32'h40046b04} /* (9, 9, 7) {real, imag} */,
  {32'hbfa36ee4, 32'hbf848de4} /* (9, 9, 6) {real, imag} */,
  {32'hbfeeb54c, 32'hbe9fe661} /* (9, 9, 5) {real, imag} */,
  {32'hbf784078, 32'h3f2f0690} /* (9, 9, 4) {real, imag} */,
  {32'h3fc6ee2e, 32'h3eed7998} /* (9, 9, 3) {real, imag} */,
  {32'h400097d9, 32'h3fb90464} /* (9, 9, 2) {real, imag} */,
  {32'hbe8c3390, 32'h3e91d37b} /* (9, 9, 1) {real, imag} */,
  {32'h3cf7d3e0, 32'h3bcfe100} /* (9, 9, 0) {real, imag} */,
  {32'h3f8d2f7d, 32'hbecfd9b4} /* (9, 8, 31) {real, imag} */,
  {32'h3f81cbbd, 32'hbd6d4e10} /* (9, 8, 30) {real, imag} */,
  {32'hbfc02bac, 32'hbde19e00} /* (9, 8, 29) {real, imag} */,
  {32'hc0188486, 32'hbe671a22} /* (9, 8, 28) {real, imag} */,
  {32'hbf64ee88, 32'h3ece00e8} /* (9, 8, 27) {real, imag} */,
  {32'hbe3572ec, 32'hbea5002c} /* (9, 8, 26) {real, imag} */,
  {32'h3e341521, 32'h3fdd99d8} /* (9, 8, 25) {real, imag} */,
  {32'h3e1cad00, 32'h401f2daa} /* (9, 8, 24) {real, imag} */,
  {32'h3fa62682, 32'h3f6b95e6} /* (9, 8, 23) {real, imag} */,
  {32'h40088a7a, 32'h3facd0ac} /* (9, 8, 22) {real, imag} */,
  {32'h3f0645ea, 32'hbf6a0a10} /* (9, 8, 21) {real, imag} */,
  {32'h3f8abc1a, 32'hc0064fdf} /* (9, 8, 20) {real, imag} */,
  {32'hbe43cd88, 32'hbf8519d5} /* (9, 8, 19) {real, imag} */,
  {32'h3e9eac19, 32'hbfe4ed0b} /* (9, 8, 18) {real, imag} */,
  {32'h3edb3542, 32'hc02b7344} /* (9, 8, 17) {real, imag} */,
  {32'h3f95dd80, 32'hbe6dc9b0} /* (9, 8, 16) {real, imag} */,
  {32'h3fd61d7d, 32'h3fa6503e} /* (9, 8, 15) {real, imag} */,
  {32'h40012e36, 32'h3fa9b4ba} /* (9, 8, 14) {real, imag} */,
  {32'h3fc5872e, 32'h3fb2113e} /* (9, 8, 13) {real, imag} */,
  {32'h402a67ea, 32'h3fc2fcb3} /* (9, 8, 12) {real, imag} */,
  {32'h3fb5da74, 32'hbfdba218} /* (9, 8, 11) {real, imag} */,
  {32'h3f0a04f2, 32'hbecd5538} /* (9, 8, 10) {real, imag} */,
  {32'hbea961fc, 32'h3f8d2b54} /* (9, 8, 9) {real, imag} */,
  {32'hbee61e38, 32'h3d142200} /* (9, 8, 8) {real, imag} */,
  {32'hbe776a46, 32'h400f8d60} /* (9, 8, 7) {real, imag} */,
  {32'hbf589d71, 32'hbeb3d1a2} /* (9, 8, 6) {real, imag} */,
  {32'hbf28db6a, 32'hbe858624} /* (9, 8, 5) {real, imag} */,
  {32'hbecf533a, 32'hbe3176c8} /* (9, 8, 4) {real, imag} */,
  {32'h3f635b7c, 32'h3f1a9174} /* (9, 8, 3) {real, imag} */,
  {32'h3f5b90a6, 32'h401dad1a} /* (9, 8, 2) {real, imag} */,
  {32'h3f75966a, 32'h3f73891c} /* (9, 8, 1) {real, imag} */,
  {32'h3f8f261b, 32'h3f082e02} /* (9, 8, 0) {real, imag} */,
  {32'h3f575e1f, 32'h3d9eef48} /* (9, 7, 31) {real, imag} */,
  {32'h3f999d82, 32'hbf4f80c4} /* (9, 7, 30) {real, imag} */,
  {32'hbebd9488, 32'hbf901d7f} /* (9, 7, 29) {real, imag} */,
  {32'hbfed9cf5, 32'h3db75428} /* (9, 7, 28) {real, imag} */,
  {32'hbcd449d8, 32'h3e54fd13} /* (9, 7, 27) {real, imag} */,
  {32'h3ebeb83e, 32'h3ea36328} /* (9, 7, 26) {real, imag} */,
  {32'h3e6dff58, 32'h401e44ea} /* (9, 7, 25) {real, imag} */,
  {32'h3ff60ed0, 32'h400c0420} /* (9, 7, 24) {real, imag} */,
  {32'h3e3f7e28, 32'hbd904a20} /* (9, 7, 23) {real, imag} */,
  {32'h3f42f122, 32'h3fa34ab2} /* (9, 7, 22) {real, imag} */,
  {32'h3f0e230a, 32'hbe48ff60} /* (9, 7, 21) {real, imag} */,
  {32'h3e996850, 32'hbfc7e818} /* (9, 7, 20) {real, imag} */,
  {32'hbdd744a8, 32'h3eae5cbe} /* (9, 7, 19) {real, imag} */,
  {32'h3f35c454, 32'hbe0a9380} /* (9, 7, 18) {real, imag} */,
  {32'h3f2227d5, 32'hbfe9bcf5} /* (9, 7, 17) {real, imag} */,
  {32'h3ddd3c10, 32'h3e8928c0} /* (9, 7, 16) {real, imag} */,
  {32'h3fd76d52, 32'hbf96284a} /* (9, 7, 15) {real, imag} */,
  {32'h3fcf5f08, 32'hbf8f8f44} /* (9, 7, 14) {real, imag} */,
  {32'h3fbcbe71, 32'hbeceb1fd} /* (9, 7, 13) {real, imag} */,
  {32'h40209d7c, 32'h3f36fdc0} /* (9, 7, 12) {real, imag} */,
  {32'h3fbbaa86, 32'hbfa6be38} /* (9, 7, 11) {real, imag} */,
  {32'h3f04625e, 32'hbfb7f2ef} /* (9, 7, 10) {real, imag} */,
  {32'h3da977c8, 32'hbfd83258} /* (9, 7, 9) {real, imag} */,
  {32'h3e6259a6, 32'hbfb4ee04} /* (9, 7, 8) {real, imag} */,
  {32'h3df8c350, 32'h3ff13eee} /* (9, 7, 7) {real, imag} */,
  {32'hbdd29e84, 32'h3fdbab22} /* (9, 7, 6) {real, imag} */,
  {32'hbfed0bc5, 32'h3f721c82} /* (9, 7, 5) {real, imag} */,
  {32'hbf3ac94c, 32'h3e0f60ba} /* (9, 7, 4) {real, imag} */,
  {32'h3fa1b391, 32'hbf661374} /* (9, 7, 3) {real, imag} */,
  {32'hbf182cfd, 32'h3f619ee8} /* (9, 7, 2) {real, imag} */,
  {32'hbeff9bcc, 32'h3e8b99f8} /* (9, 7, 1) {real, imag} */,
  {32'h3e8851b4, 32'hbe4ab788} /* (9, 7, 0) {real, imag} */,
  {32'h3f5cdc5b, 32'h3ef71858} /* (9, 6, 31) {real, imag} */,
  {32'h3f56ce70, 32'hbf4c7ef0} /* (9, 6, 30) {real, imag} */,
  {32'h3e95a0be, 32'hbcdd7e40} /* (9, 6, 29) {real, imag} */,
  {32'h3e580a00, 32'h3ed51464} /* (9, 6, 28) {real, imag} */,
  {32'h3ffdbb07, 32'h3e441950} /* (9, 6, 27) {real, imag} */,
  {32'h3feb3344, 32'h3f6c8dcf} /* (9, 6, 26) {real, imag} */,
  {32'hbfb85e19, 32'h3fa96f0a} /* (9, 6, 25) {real, imag} */,
  {32'hbf6c1ec0, 32'hbe8eca5b} /* (9, 6, 24) {real, imag} */,
  {32'hbf660a68, 32'hbf8d4bad} /* (9, 6, 23) {real, imag} */,
  {32'hbf2efd64, 32'h3fc47d32} /* (9, 6, 22) {real, imag} */,
  {32'hbf6a7d5a, 32'h3f823952} /* (9, 6, 21) {real, imag} */,
  {32'hbf48b698, 32'hbf7e6860} /* (9, 6, 20) {real, imag} */,
  {32'hbe1f909c, 32'h3ec59a7c} /* (9, 6, 19) {real, imag} */,
  {32'h3f8965dd, 32'hbe210a78} /* (9, 6, 18) {real, imag} */,
  {32'h3f364372, 32'hbf0aab6c} /* (9, 6, 17) {real, imag} */,
  {32'hbf58ce54, 32'h3fcd6e76} /* (9, 6, 16) {real, imag} */,
  {32'h3f1a0811, 32'h3edf6337} /* (9, 6, 15) {real, imag} */,
  {32'h3f64aefa, 32'hbe89099a} /* (9, 6, 14) {real, imag} */,
  {32'h3f334894, 32'hbe818df0} /* (9, 6, 13) {real, imag} */,
  {32'hbf3f0f5f, 32'hbdd4a480} /* (9, 6, 12) {real, imag} */,
  {32'hbfc0b339, 32'hbe49e7f0} /* (9, 6, 11) {real, imag} */,
  {32'hbf8717a6, 32'hbf227795} /* (9, 6, 10) {real, imag} */,
  {32'hbf3b92ff, 32'hbfaba607} /* (9, 6, 9) {real, imag} */,
  {32'h3facb9c5, 32'hbff12a53} /* (9, 6, 8) {real, imag} */,
  {32'h3e2c9186, 32'h3f51007a} /* (9, 6, 7) {real, imag} */,
  {32'hc0020d70, 32'h402e8ad7} /* (9, 6, 6) {real, imag} */,
  {32'hc02e1d10, 32'h40149c4b} /* (9, 6, 5) {real, imag} */,
  {32'h3ef4ab9c, 32'h4005c05a} /* (9, 6, 4) {real, imag} */,
  {32'h3f0dda9e, 32'h3f280a3c} /* (9, 6, 3) {real, imag} */,
  {32'hbf7ec21c, 32'hbf6ffb4e} /* (9, 6, 2) {real, imag} */,
  {32'h3f0ee8c2, 32'h3e80bc18} /* (9, 6, 1) {real, imag} */,
  {32'h3f49c3f8, 32'h3ea0eeb8} /* (9, 6, 0) {real, imag} */,
  {32'h3e17bf40, 32'h3f4e8baf} /* (9, 5, 31) {real, imag} */,
  {32'h3e984a1c, 32'h3e13f5fa} /* (9, 5, 30) {real, imag} */,
  {32'hbf23dd1c, 32'hbe2f73f0} /* (9, 5, 29) {real, imag} */,
  {32'hbf7fcdee, 32'h3f25ebf7} /* (9, 5, 28) {real, imag} */,
  {32'h3f6810a0, 32'h3ecd7564} /* (9, 5, 27) {real, imag} */,
  {32'h3df1ec88, 32'h3f6feb4a} /* (9, 5, 26) {real, imag} */,
  {32'hbfd0fce2, 32'h3f8a2300} /* (9, 5, 25) {real, imag} */,
  {32'hbf6cdb41, 32'h3e0d4d28} /* (9, 5, 24) {real, imag} */,
  {32'hbedf50c4, 32'h3f803b08} /* (9, 5, 23) {real, imag} */,
  {32'hbe8c2c70, 32'h3fe9c667} /* (9, 5, 22) {real, imag} */,
  {32'hbf8ffee0, 32'h3e6b7330} /* (9, 5, 21) {real, imag} */,
  {32'hbff27c16, 32'hbfc445ff} /* (9, 5, 20) {real, imag} */,
  {32'hbf761fc2, 32'hbec79cf0} /* (9, 5, 19) {real, imag} */,
  {32'h3e4abc58, 32'h3e981928} /* (9, 5, 18) {real, imag} */,
  {32'hbfa66ef6, 32'h3fb5855f} /* (9, 5, 17) {real, imag} */,
  {32'hbeae398d, 32'h403c42d0} /* (9, 5, 16) {real, imag} */,
  {32'h3ece5776, 32'h4031e159} /* (9, 5, 15) {real, imag} */,
  {32'hbe1760b4, 32'h3f3f9ab5} /* (9, 5, 14) {real, imag} */,
  {32'hbde756a0, 32'h3f4ae5a8} /* (9, 5, 13) {real, imag} */,
  {32'hbf9645a0, 32'hbe144b1c} /* (9, 5, 12) {real, imag} */,
  {32'hbfb45c06, 32'h3e395dc8} /* (9, 5, 11) {real, imag} */,
  {32'hbf44a07c, 32'hbd7379d0} /* (9, 5, 10) {real, imag} */,
  {32'hbf9c45e0, 32'hbf9fb46c} /* (9, 5, 9) {real, imag} */,
  {32'h3f6a17f6, 32'hc00509a8} /* (9, 5, 8) {real, imag} */,
  {32'h3f885820, 32'hbf4060eb} /* (9, 5, 7) {real, imag} */,
  {32'hc00c16ac, 32'h3f90049b} /* (9, 5, 6) {real, imag} */,
  {32'hc0106d4b, 32'h3f7ac281} /* (9, 5, 5) {real, imag} */,
  {32'h3f1f5aba, 32'h3df969f0} /* (9, 5, 4) {real, imag} */,
  {32'h3e74bec0, 32'h3f606488} /* (9, 5, 3) {real, imag} */,
  {32'h3edfc624, 32'h3f8377d8} /* (9, 5, 2) {real, imag} */,
  {32'h3e9d33ff, 32'h3e02fd50} /* (9, 5, 1) {real, imag} */,
  {32'hbe29a19a, 32'hbf7337da} /* (9, 5, 0) {real, imag} */,
  {32'h3f86acbe, 32'h3f88e580} /* (9, 4, 31) {real, imag} */,
  {32'h40017544, 32'hbe79ed16} /* (9, 4, 30) {real, imag} */,
  {32'h3e807222, 32'h3f010f9b} /* (9, 4, 29) {real, imag} */,
  {32'hbfd856e8, 32'h40032dbe} /* (9, 4, 28) {real, imag} */,
  {32'hbfb90146, 32'h3f452e25} /* (9, 4, 27) {real, imag} */,
  {32'hbe6bd256, 32'hbef1f2c0} /* (9, 4, 26) {real, imag} */,
  {32'h3ec00a78, 32'h3cb54380} /* (9, 4, 25) {real, imag} */,
  {32'h3d539410, 32'h3fa3f720} /* (9, 4, 24) {real, imag} */,
  {32'hbfa0a426, 32'h3fd42da6} /* (9, 4, 23) {real, imag} */,
  {32'hbf179e13, 32'h3d8485b8} /* (9, 4, 22) {real, imag} */,
  {32'h3e5fdc7c, 32'hbf969fc6} /* (9, 4, 21) {real, imag} */,
  {32'hbe2efb60, 32'hbfebb4fe} /* (9, 4, 20) {real, imag} */,
  {32'hbf8d80c6, 32'hbe5ead26} /* (9, 4, 19) {real, imag} */,
  {32'h3e10a508, 32'h3e8429d8} /* (9, 4, 18) {real, imag} */,
  {32'hbd98e0b0, 32'h3fa5ad42} /* (9, 4, 17) {real, imag} */,
  {32'h3f807843, 32'h3fcd43dc} /* (9, 4, 16) {real, imag} */,
  {32'h3fd523cf, 32'h3faf874c} /* (9, 4, 15) {real, imag} */,
  {32'h3fc53003, 32'h3eaea340} /* (9, 4, 14) {real, imag} */,
  {32'h3f95869e, 32'h3e9d9236} /* (9, 4, 13) {real, imag} */,
  {32'h3fcff4c4, 32'hbeb64290} /* (9, 4, 12) {real, imag} */,
  {32'h3fa18048, 32'hbf870ead} /* (9, 4, 11) {real, imag} */,
  {32'h3f865ed8, 32'hbf268f3e} /* (9, 4, 10) {real, imag} */,
  {32'hbf038cb2, 32'hbf0a351c} /* (9, 4, 9) {real, imag} */,
  {32'hbf370b3c, 32'hbf1dbd06} /* (9, 4, 8) {real, imag} */,
  {32'h3eb35c2e, 32'hbf0016ae} /* (9, 4, 7) {real, imag} */,
  {32'hbecacc78, 32'hbec21417} /* (9, 4, 6) {real, imag} */,
  {32'hc00f68ef, 32'hbe0df43c} /* (9, 4, 5) {real, imag} */,
  {32'hbfd72227, 32'h3e5dfad0} /* (9, 4, 4) {real, imag} */,
  {32'h3ef273ac, 32'h3fab8ca4} /* (9, 4, 3) {real, imag} */,
  {32'h3f6e7b2b, 32'h3fe11264} /* (9, 4, 2) {real, imag} */,
  {32'hbf30ed41, 32'h3fce2cbd} /* (9, 4, 1) {real, imag} */,
  {32'hbf0a3034, 32'h3f294b11} /* (9, 4, 0) {real, imag} */,
  {32'h3f8fe1bc, 32'h3f02fe2a} /* (9, 3, 31) {real, imag} */,
  {32'h3eda690e, 32'hbfd30d90} /* (9, 3, 30) {real, imag} */,
  {32'hbe99a623, 32'hbfa5c9af} /* (9, 3, 29) {real, imag} */,
  {32'hbf9d5007, 32'h402bcdf0} /* (9, 3, 28) {real, imag} */,
  {32'hbfc29076, 32'h40037cac} /* (9, 3, 27) {real, imag} */,
  {32'hbf0f3f8b, 32'hbe416ed0} /* (9, 3, 26) {real, imag} */,
  {32'hbfcdbc2f, 32'h3e93dcca} /* (9, 3, 25) {real, imag} */,
  {32'hbf8c2f9e, 32'h400d8d7d} /* (9, 3, 24) {real, imag} */,
  {32'hbfad60a5, 32'h404af5ef} /* (9, 3, 23) {real, imag} */,
  {32'hbfc30f92, 32'h3f2151d8} /* (9, 3, 22) {real, imag} */,
  {32'hbf0e7854, 32'hbec166f7} /* (9, 3, 21) {real, imag} */,
  {32'h3db83190, 32'hbefda097} /* (9, 3, 20) {real, imag} */,
  {32'hbe948bfe, 32'h3d3acc00} /* (9, 3, 19) {real, imag} */,
  {32'h3f4ca30a, 32'hbf315702} /* (9, 3, 18) {real, imag} */,
  {32'hbd94e8c0, 32'h3f19b534} /* (9, 3, 17) {real, imag} */,
  {32'h3ebd5480, 32'h3f1d668e} /* (9, 3, 16) {real, imag} */,
  {32'h3f33de0e, 32'h3f9a2ff9} /* (9, 3, 15) {real, imag} */,
  {32'h3f3d6772, 32'hbdef2b40} /* (9, 3, 14) {real, imag} */,
  {32'h3fa8727e, 32'h3eef92d4} /* (9, 3, 13) {real, imag} */,
  {32'h40396c82, 32'h3f897b30} /* (9, 3, 12) {real, imag} */,
  {32'h40285c72, 32'hbfd6ebc6} /* (9, 3, 11) {real, imag} */,
  {32'h3fb6e96e, 32'hbfc6b2bd} /* (9, 3, 10) {real, imag} */,
  {32'hbceec3c0, 32'hbedeee22} /* (9, 3, 9) {real, imag} */,
  {32'hbe678790, 32'hbe834683} /* (9, 3, 8) {real, imag} */,
  {32'h3f3960c9, 32'hbf3732a6} /* (9, 3, 7) {real, imag} */,
  {32'h3f546cb8, 32'h3d428790} /* (9, 3, 6) {real, imag} */,
  {32'hbee5c86a, 32'hbfb61a3e} /* (9, 3, 5) {real, imag} */,
  {32'hbfe9122a, 32'hbef2ce48} /* (9, 3, 4) {real, imag} */,
  {32'h3ec98f13, 32'h4009cc38} /* (9, 3, 3) {real, imag} */,
  {32'h3e000c40, 32'h402fb804} /* (9, 3, 2) {real, imag} */,
  {32'hc0184b5e, 32'h3fe82858} /* (9, 3, 1) {real, imag} */,
  {32'hbf2bdf0e, 32'h3fdbc580} /* (9, 3, 0) {real, imag} */,
  {32'hbe0727f4, 32'hbe0900fe} /* (9, 2, 31) {real, imag} */,
  {32'hbfbc9fba, 32'hbf6dcdc4} /* (9, 2, 30) {real, imag} */,
  {32'hbf1f7b46, 32'hbe8a57e0} /* (9, 2, 29) {real, imag} */,
  {32'h3e6e9ea4, 32'h3fec2c8e} /* (9, 2, 28) {real, imag} */,
  {32'hbf63ab96, 32'h3fc60932} /* (9, 2, 27) {real, imag} */,
  {32'hbf05a08e, 32'hbee554e0} /* (9, 2, 26) {real, imag} */,
  {32'hbfa613f2, 32'hbf06125c} /* (9, 2, 25) {real, imag} */,
  {32'hbfae6947, 32'h3ed50998} /* (9, 2, 24) {real, imag} */,
  {32'h3e1dab3c, 32'h3fe6750e} /* (9, 2, 23) {real, imag} */,
  {32'h3f38f381, 32'h3fdc07cb} /* (9, 2, 22) {real, imag} */,
  {32'h3f02459a, 32'h3e2fb77c} /* (9, 2, 21) {real, imag} */,
  {32'h3e081048, 32'hbe875fc5} /* (9, 2, 20) {real, imag} */,
  {32'hbe04a60a, 32'h3db214c8} /* (9, 2, 19) {real, imag} */,
  {32'h3f4e2955, 32'hbf875303} /* (9, 2, 18) {real, imag} */,
  {32'h3e1f6832, 32'hbeda4222} /* (9, 2, 17) {real, imag} */,
  {32'hbf8f3355, 32'h3e1894a0} /* (9, 2, 16) {real, imag} */,
  {32'hbd7cfb80, 32'hbec897d4} /* (9, 2, 15) {real, imag} */,
  {32'hbec43ec0, 32'hbee657d8} /* (9, 2, 14) {real, imag} */,
  {32'hbf99438d, 32'h3ee6437b} /* (9, 2, 13) {real, imag} */,
  {32'h3f7319a0, 32'h3f3b6099} /* (9, 2, 12) {real, imag} */,
  {32'h3fc937d8, 32'h3f18d384} /* (9, 2, 11) {real, imag} */,
  {32'h3fb766ef, 32'hbe1ef5b4} /* (9, 2, 10) {real, imag} */,
  {32'h3dc198d0, 32'hbf8d408e} /* (9, 2, 9) {real, imag} */,
  {32'h3f9bdb22, 32'hbfd6bf5c} /* (9, 2, 8) {real, imag} */,
  {32'h4000e204, 32'hbf9a4b7b} /* (9, 2, 7) {real, imag} */,
  {32'h3fdfad48, 32'h3f42d0b0} /* (9, 2, 6) {real, imag} */,
  {32'hbf80442e, 32'hbeeaa640} /* (9, 2, 5) {real, imag} */,
  {32'hbf0ab8b8, 32'hbfa657aa} /* (9, 2, 4) {real, imag} */,
  {32'h40024096, 32'h3fdab899} /* (9, 2, 3) {real, imag} */,
  {32'hbe83a872, 32'h402329ae} /* (9, 2, 2) {real, imag} */,
  {32'hbf536b61, 32'h3ffe6c4e} /* (9, 2, 1) {real, imag} */,
  {32'h3ef18f36, 32'h3fc7cb10} /* (9, 2, 0) {real, imag} */,
  {32'hbf8ff3b4, 32'h3e97a4c0} /* (9, 1, 31) {real, imag} */,
  {32'hbfd9589b, 32'h3e22b67a} /* (9, 1, 30) {real, imag} */,
  {32'hbf356497, 32'h3ebee2e4} /* (9, 1, 29) {real, imag} */,
  {32'h3f994710, 32'h3e2d2c9c} /* (9, 1, 28) {real, imag} */,
  {32'hbd82e0fc, 32'hbf6c0e83} /* (9, 1, 27) {real, imag} */,
  {32'hbcfd7070, 32'hbfb11ef6} /* (9, 1, 26) {real, imag} */,
  {32'hbfbef23b, 32'hbf7a3906} /* (9, 1, 25) {real, imag} */,
  {32'hbf2f9bcf, 32'hbf6a6c64} /* (9, 1, 24) {real, imag} */,
  {32'hbe16c6f4, 32'h3f00777c} /* (9, 1, 23) {real, imag} */,
  {32'hbe2f9e88, 32'h3fbdb0a5} /* (9, 1, 22) {real, imag} */,
  {32'hbf82df42, 32'h3d8d1590} /* (9, 1, 21) {real, imag} */,
  {32'hbf3ce6f3, 32'hbfbe0609} /* (9, 1, 20) {real, imag} */,
  {32'hbf2970d3, 32'hbf24415b} /* (9, 1, 19) {real, imag} */,
  {32'h3e610848, 32'h3edc2118} /* (9, 1, 18) {real, imag} */,
  {32'hbff6d1b2, 32'h3f66e632} /* (9, 1, 17) {real, imag} */,
  {32'hc03a376e, 32'h3f5467da} /* (9, 1, 16) {real, imag} */,
  {32'hbf369605, 32'h3fadd1dc} /* (9, 1, 15) {real, imag} */,
  {32'h3edafa9d, 32'h3fbf23d0} /* (9, 1, 14) {real, imag} */,
  {32'hbf264146, 32'hbf2efacf} /* (9, 1, 13) {real, imag} */,
  {32'hbfb1e61d, 32'h3cdd8900} /* (9, 1, 12) {real, imag} */,
  {32'hbe8b058e, 32'hbcaa5480} /* (9, 1, 11) {real, imag} */,
  {32'h3f1014ec, 32'hbf63b6fd} /* (9, 1, 10) {real, imag} */,
  {32'h3e857b9c, 32'hbf40e8c0} /* (9, 1, 9) {real, imag} */,
  {32'h3fb6611c, 32'hbf9094d8} /* (9, 1, 8) {real, imag} */,
  {32'h401c873e, 32'hbf0c0a7a} /* (9, 1, 7) {real, imag} */,
  {32'h40071087, 32'h3fc88fb8} /* (9, 1, 6) {real, imag} */,
  {32'hbf3f69fb, 32'h3f91cd0b} /* (9, 1, 5) {real, imag} */,
  {32'hbe65b558, 32'hbef9cc50} /* (9, 1, 4) {real, imag} */,
  {32'h3eebf23e, 32'h3f15938c} /* (9, 1, 3) {real, imag} */,
  {32'hbfd387b3, 32'h3ef22022} /* (9, 1, 2) {real, imag} */,
  {32'hbf2b1fe0, 32'h3ecef488} /* (9, 1, 1) {real, imag} */,
  {32'h3e9898de, 32'h3f19a47d} /* (9, 1, 0) {real, imag} */,
  {32'hbeea2a49, 32'h3f317aa0} /* (9, 0, 31) {real, imag} */,
  {32'hbf097b26, 32'hbeac8147} /* (9, 0, 30) {real, imag} */,
  {32'hbf0527c2, 32'hbf6e6183} /* (9, 0, 29) {real, imag} */,
  {32'h3d768120, 32'hbf070ae0} /* (9, 0, 28) {real, imag} */,
  {32'h3e1903ac, 32'hbe6b4912} /* (9, 0, 27) {real, imag} */,
  {32'hbf127556, 32'hbcec32e0} /* (9, 0, 26) {real, imag} */,
  {32'hbf48dffa, 32'hbe50bc70} /* (9, 0, 25) {real, imag} */,
  {32'hbe84baa8, 32'hbf5c1d35} /* (9, 0, 24) {real, imag} */,
  {32'hbe81fbd8, 32'hbe44ea7a} /* (9, 0, 23) {real, imag} */,
  {32'hbf50e0b2, 32'h3f04c526} /* (9, 0, 22) {real, imag} */,
  {32'hbfc8329e, 32'h3e890908} /* (9, 0, 21) {real, imag} */,
  {32'hbf640eeb, 32'hbe86880a} /* (9, 0, 20) {real, imag} */,
  {32'h3e4f9658, 32'hbf1ad854} /* (9, 0, 19) {real, imag} */,
  {32'h3e0d346b, 32'hbe92d57a} /* (9, 0, 18) {real, imag} */,
  {32'hbfe0bbee, 32'hbeba251c} /* (9, 0, 17) {real, imag} */,
  {32'hbfa3b486, 32'hbe32d448} /* (9, 0, 16) {real, imag} */,
  {32'hbe42c2c6, 32'h3ef5f19c} /* (9, 0, 15) {real, imag} */,
  {32'h3f1e8fc6, 32'h3fa7f1fe} /* (9, 0, 14) {real, imag} */,
  {32'h3f8020f3, 32'h3dc08180} /* (9, 0, 13) {real, imag} */,
  {32'hbf54e3d8, 32'hbe8a28bc} /* (9, 0, 12) {real, imag} */,
  {32'hbeed88ae, 32'hbdbf9d5c} /* (9, 0, 11) {real, imag} */,
  {32'h3effe34c, 32'h3d857b28} /* (9, 0, 10) {real, imag} */,
  {32'h3eae5d61, 32'h3f80fd95} /* (9, 0, 9) {real, imag} */,
  {32'h3f4659b1, 32'h3f288530} /* (9, 0, 8) {real, imag} */,
  {32'h3fe2941b, 32'h3e83888e} /* (9, 0, 7) {real, imag} */,
  {32'h3f8eba0f, 32'h3f38852c} /* (9, 0, 6) {real, imag} */,
  {32'h3ec57a8b, 32'h3f114b8f} /* (9, 0, 5) {real, imag} */,
  {32'hbf1768f6, 32'h3d814498} /* (9, 0, 4) {real, imag} */,
  {32'hbee5823a, 32'hbefbb9ec} /* (9, 0, 3) {real, imag} */,
  {32'hbf1dba37, 32'hbf6ac649} /* (9, 0, 2) {real, imag} */,
  {32'hbe8d1f54, 32'h3f1d44a4} /* (9, 0, 1) {real, imag} */,
  {32'h3eef2767, 32'h3f1c906d} /* (9, 0, 0) {real, imag} */,
  {32'hbf53abfe, 32'h3e2fa19c} /* (8, 31, 31) {real, imag} */,
  {32'hbfae7ae0, 32'hbee1e9ea} /* (8, 31, 30) {real, imag} */,
  {32'hbffe45e2, 32'hbf0cd25a} /* (8, 31, 29) {real, imag} */,
  {32'hc0084a97, 32'h3fadacab} /* (8, 31, 28) {real, imag} */,
  {32'hbfab89b6, 32'h3f0d89cb} /* (8, 31, 27) {real, imag} */,
  {32'hbdd74d38, 32'hbf464f0e} /* (8, 31, 26) {real, imag} */,
  {32'hc00b75ce, 32'h3fb12704} /* (8, 31, 25) {real, imag} */,
  {32'hc03f9031, 32'h3f2f5886} /* (8, 31, 24) {real, imag} */,
  {32'hbffb9831, 32'h3fceff88} /* (8, 31, 23) {real, imag} */,
  {32'hbfb1e41f, 32'h3fc9a143} /* (8, 31, 22) {real, imag} */,
  {32'hbe5c6731, 32'h3f4af048} /* (8, 31, 21) {real, imag} */,
  {32'h3f5a23e2, 32'hbf66a744} /* (8, 31, 20) {real, imag} */,
  {32'h3f8aac40, 32'hbf9bce02} /* (8, 31, 19) {real, imag} */,
  {32'h3f0ea902, 32'hbedc20a6} /* (8, 31, 18) {real, imag} */,
  {32'h3e10cf8a, 32'hbee40574} /* (8, 31, 17) {real, imag} */,
  {32'h3f1fbc13, 32'hbf42c2b8} /* (8, 31, 16) {real, imag} */,
  {32'hbf0546d8, 32'hbfe3b630} /* (8, 31, 15) {real, imag} */,
  {32'h3f85fe5d, 32'hbfa569a6} /* (8, 31, 14) {real, imag} */,
  {32'h3ff3eeac, 32'hbfdd24b6} /* (8, 31, 13) {real, imag} */,
  {32'h3f7e5ec8, 32'hc0002a66} /* (8, 31, 12) {real, imag} */,
  {32'h3f9de393, 32'hc018d738} /* (8, 31, 11) {real, imag} */,
  {32'h3f413b9d, 32'hbf50afbb} /* (8, 31, 10) {real, imag} */,
  {32'h3fc64d3a, 32'h3e4756ea} /* (8, 31, 9) {real, imag} */,
  {32'h3e4eb1a0, 32'h3eccc150} /* (8, 31, 8) {real, imag} */,
  {32'h3ee88ff0, 32'h40016d47} /* (8, 31, 7) {real, imag} */,
  {32'hbf5c7e77, 32'h3fe44b48} /* (8, 31, 6) {real, imag} */,
  {32'hc002f4c6, 32'h3ffb7e3d} /* (8, 31, 5) {real, imag} */,
  {32'hbf0b0010, 32'h3fea50e6} /* (8, 31, 4) {real, imag} */,
  {32'hbefc5662, 32'h3fd047e3} /* (8, 31, 3) {real, imag} */,
  {32'h3f3c028d, 32'h404cc009} /* (8, 31, 2) {real, imag} */,
  {32'hbf3f0720, 32'h3ff86a3e} /* (8, 31, 1) {real, imag} */,
  {32'hc0170cf9, 32'h3e496c0e} /* (8, 31, 0) {real, imag} */,
  {32'hbfda2124, 32'h3ee5b8ef} /* (8, 30, 31) {real, imag} */,
  {32'hc0457104, 32'hbf874822} /* (8, 30, 30) {real, imag} */,
  {32'hc055c0a4, 32'hbf093e8e} /* (8, 30, 29) {real, imag} */,
  {32'hc0295e30, 32'h402569f2} /* (8, 30, 28) {real, imag} */,
  {32'hc00e09d4, 32'hbee4b1c8} /* (8, 30, 27) {real, imag} */,
  {32'hbfc2f25e, 32'hbfe5259a} /* (8, 30, 26) {real, imag} */,
  {32'hc01a8e77, 32'h3f990209} /* (8, 30, 25) {real, imag} */,
  {32'hc05cbc4f, 32'h3f0cbae0} /* (8, 30, 24) {real, imag} */,
  {32'hc03b4795, 32'h40029d99} /* (8, 30, 23) {real, imag} */,
  {32'hbf29049f, 32'h4034a9c0} /* (8, 30, 22) {real, imag} */,
  {32'h3ee1090e, 32'h3db35398} /* (8, 30, 21) {real, imag} */,
  {32'h3f051d2a, 32'hc02039d6} /* (8, 30, 20) {real, imag} */,
  {32'h3f0155af, 32'hc042c433} /* (8, 30, 19) {real, imag} */,
  {32'h4008c014, 32'hbfdfebbe} /* (8, 30, 18) {real, imag} */,
  {32'h400c68e6, 32'hbfd58abf} /* (8, 30, 17) {real, imag} */,
  {32'h3fca4bcc, 32'hc03160ff} /* (8, 30, 16) {real, imag} */,
  {32'h3fd41a5a, 32'hc0574ca6} /* (8, 30, 15) {real, imag} */,
  {32'h405fe2a6, 32'hc04ee3f4} /* (8, 30, 14) {real, imag} */,
  {32'h4038c278, 32'hc043d46e} /* (8, 30, 13) {real, imag} */,
  {32'h400fcf1f, 32'hc024dfd0} /* (8, 30, 12) {real, imag} */,
  {32'h4027ca66, 32'hbf87016a} /* (8, 30, 11) {real, imag} */,
  {32'h3f8aaa63, 32'h3f2bdcba} /* (8, 30, 10) {real, imag} */,
  {32'h3f83f54e, 32'hbd558750} /* (8, 30, 9) {real, imag} */,
  {32'hbf5c3150, 32'h3f2de8de} /* (8, 30, 8) {real, imag} */,
  {32'hbfb70d25, 32'h40010fe1} /* (8, 30, 7) {real, imag} */,
  {32'hc009babe, 32'h405327a0} /* (8, 30, 6) {real, imag} */,
  {32'hc01b64a0, 32'h40a70a93} /* (8, 30, 5) {real, imag} */,
  {32'hbfa5fcb5, 32'h404b3d8a} /* (8, 30, 4) {real, imag} */,
  {32'hbfd8e2ec, 32'h3f96427e} /* (8, 30, 3) {real, imag} */,
  {32'hbe65cc48, 32'h405fed59} /* (8, 30, 2) {real, imag} */,
  {32'hbfe783a6, 32'h40159413} /* (8, 30, 1) {real, imag} */,
  {32'hc0444253, 32'h3f7fa3c4} /* (8, 30, 0) {real, imag} */,
  {32'hc01aee8d, 32'hbf0c5460} /* (8, 29, 31) {real, imag} */,
  {32'hc04259fa, 32'h3f500c03} /* (8, 29, 30) {real, imag} */,
  {32'hc023c67e, 32'h403529b3} /* (8, 29, 29) {real, imag} */,
  {32'hbfdb9e09, 32'h4047aea2} /* (8, 29, 28) {real, imag} */,
  {32'hbfe3461f, 32'h3fae807c} /* (8, 29, 27) {real, imag} */,
  {32'hbf88ec2d, 32'h3f4d389e} /* (8, 29, 26) {real, imag} */,
  {32'hbe0e3758, 32'h3f967eba} /* (8, 29, 25) {real, imag} */,
  {32'hbffe1922, 32'h3e8f03e2} /* (8, 29, 24) {real, imag} */,
  {32'hc004da7b, 32'h3fae5942} /* (8, 29, 23) {real, imag} */,
  {32'h3f2a3fcd, 32'h404031b9} /* (8, 29, 22) {real, imag} */,
  {32'h3fdb2c03, 32'h3f79b57e} /* (8, 29, 21) {real, imag} */,
  {32'h3ebb33aa, 32'hbffc6a27} /* (8, 29, 20) {real, imag} */,
  {32'hc00ff469, 32'hbff53587} /* (8, 29, 19) {real, imag} */,
  {32'h3e8b354a, 32'hbfeb489a} /* (8, 29, 18) {real, imag} */,
  {32'h400e2188, 32'hbf8fff74} /* (8, 29, 17) {real, imag} */,
  {32'h3fc19f20, 32'hbfe05037} /* (8, 29, 16) {real, imag} */,
  {32'h400d96c0, 32'hbfd50394} /* (8, 29, 15) {real, imag} */,
  {32'h40233310, 32'hbfebb05a} /* (8, 29, 14) {real, imag} */,
  {32'h3fe27c3b, 32'hbfe5c8ef} /* (8, 29, 13) {real, imag} */,
  {32'h40226380, 32'hbfcc1970} /* (8, 29, 12) {real, imag} */,
  {32'h406e6899, 32'hbed0ecb4} /* (8, 29, 11) {real, imag} */,
  {32'h3eb65080, 32'h3fff9863} /* (8, 29, 10) {real, imag} */,
  {32'hc030d09b, 32'h4024ec95} /* (8, 29, 9) {real, imag} */,
  {32'hc03c675f, 32'h400f7c85} /* (8, 29, 8) {real, imag} */,
  {32'hc002823a, 32'h3fd0fec4} /* (8, 29, 7) {real, imag} */,
  {32'hbfea15b6, 32'h4040dfc5} /* (8, 29, 6) {real, imag} */,
  {32'hc0033ee9, 32'h409d45cc} /* (8, 29, 5) {real, imag} */,
  {32'hbf144b7e, 32'h408bf74e} /* (8, 29, 4) {real, imag} */,
  {32'hbee7d2b8, 32'h402a474c} /* (8, 29, 3) {real, imag} */,
  {32'h3ec522ac, 32'h4051ab44} /* (8, 29, 2) {real, imag} */,
  {32'hbfff86c6, 32'h3fb3dd57} /* (8, 29, 1) {real, imag} */,
  {32'hc053dcf2, 32'h3fa61bf2} /* (8, 29, 0) {real, imag} */,
  {32'hc0118782, 32'h3e780d4a} /* (8, 28, 31) {real, imag} */,
  {32'hc0169cb8, 32'h403a2dfc} /* (8, 28, 30) {real, imag} */,
  {32'hbfd02f8e, 32'h40597ad3} /* (8, 28, 29) {real, imag} */,
  {32'hbf753ed4, 32'h400f406d} /* (8, 28, 28) {real, imag} */,
  {32'hbfd568bb, 32'h400028a5} /* (8, 28, 27) {real, imag} */,
  {32'hbf3c9fb2, 32'h405eea43} /* (8, 28, 26) {real, imag} */,
  {32'h3f2df2b0, 32'h3ff5a3ba} /* (8, 28, 25) {real, imag} */,
  {32'hc00e0838, 32'hbd79f780} /* (8, 28, 24) {real, imag} */,
  {32'hbfd660b3, 32'h4044d5d2} /* (8, 28, 23) {real, imag} */,
  {32'h3ef1a1b5, 32'h403ebdc2} /* (8, 28, 22) {real, imag} */,
  {32'h3faf77da, 32'h400ac3b6} /* (8, 28, 21) {real, imag} */,
  {32'h3f314c66, 32'hbfb559a6} /* (8, 28, 20) {real, imag} */,
  {32'hbfc0f097, 32'hc0102176} /* (8, 28, 19) {real, imag} */,
  {32'hbcadd760, 32'hc02aa3c6} /* (8, 28, 18) {real, imag} */,
  {32'h3e836358, 32'hbfbca286} /* (8, 28, 17) {real, imag} */,
  {32'h3f672d06, 32'hbef57e54} /* (8, 28, 16) {real, imag} */,
  {32'h401a783a, 32'h3d452bc8} /* (8, 28, 15) {real, imag} */,
  {32'h3f8d3b07, 32'hbde322f4} /* (8, 28, 14) {real, imag} */,
  {32'h3fb19bce, 32'hbf19d3ac} /* (8, 28, 13) {real, imag} */,
  {32'h3f8970c7, 32'hbfed2a86} /* (8, 28, 12) {real, imag} */,
  {32'h4042fdd2, 32'hbfa390bc} /* (8, 28, 11) {real, imag} */,
  {32'h3e76a73c, 32'h3eac68c8} /* (8, 28, 10) {real, imag} */,
  {32'hc0285fd9, 32'h402881dc} /* (8, 28, 9) {real, imag} */,
  {32'hc00fadf6, 32'h40014144} /* (8, 28, 8) {real, imag} */,
  {32'hbf0a2556, 32'h3fd5a65e} /* (8, 28, 7) {real, imag} */,
  {32'hbfdac50d, 32'h4023c928} /* (8, 28, 6) {real, imag} */,
  {32'hbfa3fbd5, 32'h405a56c0} /* (8, 28, 5) {real, imag} */,
  {32'hbe120c7c, 32'h405225b6} /* (8, 28, 4) {real, imag} */,
  {32'hbfc26d00, 32'h401236de} /* (8, 28, 3) {real, imag} */,
  {32'hbf22d3bb, 32'h40265668} /* (8, 28, 2) {real, imag} */,
  {32'hc0484cde, 32'h4017d4f1} /* (8, 28, 1) {real, imag} */,
  {32'hc056af14, 32'h40091770} /* (8, 28, 0) {real, imag} */,
  {32'hbfd1e2a0, 32'h3f96453e} /* (8, 27, 31) {real, imag} */,
  {32'hbfc82fdf, 32'h40304ddc} /* (8, 27, 30) {real, imag} */,
  {32'hc00a8a52, 32'h402e26ee} /* (8, 27, 29) {real, imag} */,
  {32'hbfb47c25, 32'h40373c9d} /* (8, 27, 28) {real, imag} */,
  {32'hc014702c, 32'h3fed2ec0} /* (8, 27, 27) {real, imag} */,
  {32'hc0241d20, 32'h4022786f} /* (8, 27, 26) {real, imag} */,
  {32'hbf9f190a, 32'h3f1d78a0} /* (8, 27, 25) {real, imag} */,
  {32'hc08940ac, 32'h3fbb608b} /* (8, 27, 24) {real, imag} */,
  {32'hc081aa2a, 32'h4082889f} /* (8, 27, 23) {real, imag} */,
  {32'hc0349d5a, 32'h406dddb4} /* (8, 27, 22) {real, imag} */,
  {32'hbf44569e, 32'h4063ec97} /* (8, 27, 21) {real, imag} */,
  {32'h3f88c502, 32'hbfc36b07} /* (8, 27, 20) {real, imag} */,
  {32'h3f0b2151, 32'hc01ec115} /* (8, 27, 19) {real, imag} */,
  {32'h3ff62378, 32'hc05d9556} /* (8, 27, 18) {real, imag} */,
  {32'h3f390b49, 32'hc068fb1a} /* (8, 27, 17) {real, imag} */,
  {32'hbeb0fc80, 32'hc048b79a} /* (8, 27, 16) {real, imag} */,
  {32'h3fea3b9b, 32'hbff32fde} /* (8, 27, 15) {real, imag} */,
  {32'h3f557cde, 32'hbf3a8da8} /* (8, 27, 14) {real, imag} */,
  {32'h3fc81176, 32'hbbb73900} /* (8, 27, 13) {real, imag} */,
  {32'h3f9fd4ad, 32'hbf9c956c} /* (8, 27, 12) {real, imag} */,
  {32'h40512108, 32'hc03e886a} /* (8, 27, 11) {real, imag} */,
  {32'h3ea4837a, 32'hbedf2fc6} /* (8, 27, 10) {real, imag} */,
  {32'hbdcc1b30, 32'h3f98570c} /* (8, 27, 9) {real, imag} */,
  {32'h3db36f70, 32'h3f8f39e8} /* (8, 27, 8) {real, imag} */,
  {32'h3d77cca0, 32'h3f627dd2} /* (8, 27, 7) {real, imag} */,
  {32'hbfdf5128, 32'h3fcab63a} /* (8, 27, 6) {real, imag} */,
  {32'h3d298740, 32'h401fcea8} /* (8, 27, 5) {real, imag} */,
  {32'h3eeffaf6, 32'h4033df8c} /* (8, 27, 4) {real, imag} */,
  {32'hbfbe3726, 32'h3fe1efac} /* (8, 27, 3) {real, imag} */,
  {32'hbfa83402, 32'h403a1d93} /* (8, 27, 2) {real, imag} */,
  {32'hbfafa9cc, 32'h401cbc85} /* (8, 27, 1) {real, imag} */,
  {32'hbfcef8c6, 32'h40070e32} /* (8, 27, 0) {real, imag} */,
  {32'hbe43ab4a, 32'h3f431e1d} /* (8, 26, 31) {real, imag} */,
  {32'hc00ddd0f, 32'h4027d2e4} /* (8, 26, 30) {real, imag} */,
  {32'hc06c6440, 32'h3fceda60} /* (8, 26, 29) {real, imag} */,
  {32'hbfdadbcc, 32'h3f2a9e10} /* (8, 26, 28) {real, imag} */,
  {32'hc00c1818, 32'h3fc87126} /* (8, 26, 27) {real, imag} */,
  {32'hc0126a6d, 32'h3f008b48} /* (8, 26, 26) {real, imag} */,
  {32'hc00a64b0, 32'h3eba0d4c} /* (8, 26, 25) {real, imag} */,
  {32'hc03e7cb4, 32'h3ffc7afa} /* (8, 26, 24) {real, imag} */,
  {32'hbfe3145f, 32'h3fd4c85a} /* (8, 26, 23) {real, imag} */,
  {32'hbfa36dbd, 32'h40154034} /* (8, 26, 22) {real, imag} */,
  {32'hbecde314, 32'h405ae1f2} /* (8, 26, 21) {real, imag} */,
  {32'h3fdace00, 32'h3c038980} /* (8, 26, 20) {real, imag} */,
  {32'h400a460a, 32'hbfcd71a3} /* (8, 26, 19) {real, imag} */,
  {32'h402e4b99, 32'hc0119d2c} /* (8, 26, 18) {real, imag} */,
  {32'h40160cd0, 32'hc04b6220} /* (8, 26, 17) {real, imag} */,
  {32'h3efa613c, 32'hc08a8f46} /* (8, 26, 16) {real, imag} */,
  {32'h40254bfa, 32'hc0207975} /* (8, 26, 15) {real, imag} */,
  {32'h3ffdfce1, 32'hc02544ff} /* (8, 26, 14) {real, imag} */,
  {32'h3fe5422a, 32'hbfb1f496} /* (8, 26, 13) {real, imag} */,
  {32'h400da916, 32'hbfe2b244} /* (8, 26, 12) {real, imag} */,
  {32'h3f8c3ab7, 32'hc036a9b6} /* (8, 26, 11) {real, imag} */,
  {32'hbf6f12a4, 32'h3ff12cfe} /* (8, 26, 10) {real, imag} */,
  {32'hbea3b134, 32'h403f74da} /* (8, 26, 9) {real, imag} */,
  {32'h3e8d91f8, 32'h3f8f36b8} /* (8, 26, 8) {real, imag} */,
  {32'hc021025c, 32'h3ebbcfde} /* (8, 26, 7) {real, imag} */,
  {32'hc0510b33, 32'h3e5c9e0c} /* (8, 26, 6) {real, imag} */,
  {32'hc00ba79a, 32'h3ee4bcb8} /* (8, 26, 5) {real, imag} */,
  {32'hbf125260, 32'h3f9fb6c8} /* (8, 26, 4) {real, imag} */,
  {32'hbfe51bd1, 32'h402850b3} /* (8, 26, 3) {real, imag} */,
  {32'hc0066968, 32'h40226d84} /* (8, 26, 2) {real, imag} */,
  {32'h3e8e5aa8, 32'h400c0da6} /* (8, 26, 1) {real, imag} */,
  {32'hbe6b8fac, 32'h400379a6} /* (8, 26, 0) {real, imag} */,
  {32'hbf26097c, 32'h3f327680} /* (8, 25, 31) {real, imag} */,
  {32'hc03c4246, 32'h3fceb2f9} /* (8, 25, 30) {real, imag} */,
  {32'hc09b2253, 32'h3f308c99} /* (8, 25, 29) {real, imag} */,
  {32'hc031a9f8, 32'hbe8609f8} /* (8, 25, 28) {real, imag} */,
  {32'hbfaed643, 32'h3fddae73} /* (8, 25, 27) {real, imag} */,
  {32'hbf9d01d0, 32'h3f575ec2} /* (8, 25, 26) {real, imag} */,
  {32'hc0062ff4, 32'hbd498ec0} /* (8, 25, 25) {real, imag} */,
  {32'hbf60ac63, 32'h3ffc196f} /* (8, 25, 24) {real, imag} */,
  {32'hbefc9ae4, 32'h3f8cfdb4} /* (8, 25, 23) {real, imag} */,
  {32'hbf84651e, 32'h40003681} /* (8, 25, 22) {real, imag} */,
  {32'hbf3b8c36, 32'hbca17300} /* (8, 25, 21) {real, imag} */,
  {32'h3fa4c49a, 32'hc0151dde} /* (8, 25, 20) {real, imag} */,
  {32'h3fe819f4, 32'hc003ff42} /* (8, 25, 19) {real, imag} */,
  {32'h403120ac, 32'hbfc3767c} /* (8, 25, 18) {real, imag} */,
  {32'h408ea604, 32'hc013803c} /* (8, 25, 17) {real, imag} */,
  {32'h402fd70c, 32'hc06a8e2c} /* (8, 25, 16) {real, imag} */,
  {32'h4030d0ae, 32'hc02e4a70} /* (8, 25, 15) {real, imag} */,
  {32'h405763ac, 32'hbfbfb3ec} /* (8, 25, 14) {real, imag} */,
  {32'h405f9232, 32'h3ec24bc0} /* (8, 25, 13) {real, imag} */,
  {32'h401db3aa, 32'hc0471986} /* (8, 25, 12) {real, imag} */,
  {32'hbe0d3d80, 32'hc0189904} /* (8, 25, 11) {real, imag} */,
  {32'hc0000842, 32'h3fb6d9a8} /* (8, 25, 10) {real, imag} */,
  {32'hc03a5114, 32'h4026398c} /* (8, 25, 9) {real, imag} */,
  {32'hc02da418, 32'h4059662a} /* (8, 25, 8) {real, imag} */,
  {32'hc041a3de, 32'h3fdb8700} /* (8, 25, 7) {real, imag} */,
  {32'hc0471d92, 32'h3d5b9180} /* (8, 25, 6) {real, imag} */,
  {32'hc086ccaa, 32'h3dbdc010} /* (8, 25, 5) {real, imag} */,
  {32'hc057a03f, 32'h3f05847a} /* (8, 25, 4) {real, imag} */,
  {32'hc0634b2a, 32'h401e8595} /* (8, 25, 3) {real, imag} */,
  {32'hc032af7f, 32'h40124b2e} /* (8, 25, 2) {real, imag} */,
  {32'hbf769a58, 32'h3fde8c8a} /* (8, 25, 1) {real, imag} */,
  {32'hbebdd9e0, 32'h3fb77d4a} /* (8, 25, 0) {real, imag} */,
  {32'hbf9f1f34, 32'h3ef0ce6c} /* (8, 24, 31) {real, imag} */,
  {32'hbfc89390, 32'h3fd60bed} /* (8, 24, 30) {real, imag} */,
  {32'hc0223903, 32'h40274f7f} /* (8, 24, 29) {real, imag} */,
  {32'hbfb21cda, 32'h3fd41534} /* (8, 24, 28) {real, imag} */,
  {32'h3d0c1120, 32'h40388058} /* (8, 24, 27) {real, imag} */,
  {32'h3ed3b276, 32'h400f5587} /* (8, 24, 26) {real, imag} */,
  {32'h3eded40a, 32'hbf013758} /* (8, 24, 25) {real, imag} */,
  {32'hc0030696, 32'h3f96e3cf} /* (8, 24, 24) {real, imag} */,
  {32'hc01bae08, 32'h3fed7d65} /* (8, 24, 23) {real, imag} */,
  {32'hbf8f21b5, 32'h404bc561} /* (8, 24, 22) {real, imag} */,
  {32'hbf43ea80, 32'hbed10628} /* (8, 24, 21) {real, imag} */,
  {32'h3ffc1a77, 32'hc085511a} /* (8, 24, 20) {real, imag} */,
  {32'h3f1f73ba, 32'hc04b14c7} /* (8, 24, 19) {real, imag} */,
  {32'h3f8c92b3, 32'hbfea8485} /* (8, 24, 18) {real, imag} */,
  {32'h405ec67e, 32'hc001a1c0} /* (8, 24, 17) {real, imag} */,
  {32'h4050bb58, 32'hbfbe5441} /* (8, 24, 16) {real, imag} */,
  {32'h3f351053, 32'hbfcc623d} /* (8, 24, 15) {real, imag} */,
  {32'h4010ab94, 32'h3ed9bfcc} /* (8, 24, 14) {real, imag} */,
  {32'h4026a5fc, 32'hbf166118} /* (8, 24, 13) {real, imag} */,
  {32'h406bb1a2, 32'hbf579ace} /* (8, 24, 12) {real, imag} */,
  {32'h40186232, 32'hbf28bbb8} /* (8, 24, 11) {real, imag} */,
  {32'hbf434244, 32'h3f7be8dc} /* (8, 24, 10) {real, imag} */,
  {32'hc04a2d9e, 32'h40474ed7} /* (8, 24, 9) {real, imag} */,
  {32'hc0898078, 32'h3fdb37f7} /* (8, 24, 8) {real, imag} */,
  {32'hbf8bc0b8, 32'h3f2764fc} /* (8, 24, 7) {real, imag} */,
  {32'hbf9ece8c, 32'h3fb84ff6} /* (8, 24, 6) {real, imag} */,
  {32'hc005d076, 32'h3f827514} /* (8, 24, 5) {real, imag} */,
  {32'hbf83bfa6, 32'h3f288ae5} /* (8, 24, 4) {real, imag} */,
  {32'hc06cb4ca, 32'h3fe10704} /* (8, 24, 3) {real, imag} */,
  {32'hc091de66, 32'h40229112} /* (8, 24, 2) {real, imag} */,
  {32'hc013bb9e, 32'h4004186c} /* (8, 24, 1) {real, imag} */,
  {32'hbfdaec92, 32'h3f33309b} /* (8, 24, 0) {real, imag} */,
  {32'hbfa603c7, 32'h3d75a500} /* (8, 23, 31) {real, imag} */,
  {32'hbd2a1f20, 32'h4018fb26} /* (8, 23, 30) {real, imag} */,
  {32'h3f65981c, 32'h409e195c} /* (8, 23, 29) {real, imag} */,
  {32'hbea4c694, 32'h405e2116} /* (8, 23, 28) {real, imag} */,
  {32'hbf51f6f4, 32'h406a23fa} /* (8, 23, 27) {real, imag} */,
  {32'hbf72ce74, 32'h40292778} /* (8, 23, 26) {real, imag} */,
  {32'hbf2a4682, 32'h3f2a07e3} /* (8, 23, 25) {real, imag} */,
  {32'hbffe303c, 32'hbe870d76} /* (8, 23, 24) {real, imag} */,
  {32'hc008c420, 32'h3f966de5} /* (8, 23, 23) {real, imag} */,
  {32'hc01ca0a2, 32'h3fcf408d} /* (8, 23, 22) {real, imag} */,
  {32'hbf383eb2, 32'hbf1f8cb9} /* (8, 23, 21) {real, imag} */,
  {32'h404c6448, 32'hc032777a} /* (8, 23, 20) {real, imag} */,
  {32'h40052754, 32'hbfd1f706} /* (8, 23, 19) {real, imag} */,
  {32'h401184bf, 32'hbe9c8622} /* (8, 23, 18) {real, imag} */,
  {32'h4023c6a4, 32'hc000123e} /* (8, 23, 17) {real, imag} */,
  {32'h3ffc654b, 32'hc0234509} /* (8, 23, 16) {real, imag} */,
  {32'h3ecce3ec, 32'hc01bc7ae} /* (8, 23, 15) {real, imag} */,
  {32'h40087ed0, 32'hbeed90e0} /* (8, 23, 14) {real, imag} */,
  {32'h4029c90a, 32'hbf958f9d} /* (8, 23, 13) {real, imag} */,
  {32'h400b50f6, 32'hbef5932e} /* (8, 23, 12) {real, imag} */,
  {32'h3f8abf63, 32'hbd6eab90} /* (8, 23, 11) {real, imag} */,
  {32'hc01b9180, 32'h3fd808ff} /* (8, 23, 10) {real, imag} */,
  {32'hc03d7405, 32'h407b722c} /* (8, 23, 9) {real, imag} */,
  {32'hc08e25da, 32'h3fe83b1a} /* (8, 23, 8) {real, imag} */,
  {32'hbf86418c, 32'h3fa6186a} /* (8, 23, 7) {real, imag} */,
  {32'hbfbeee80, 32'h4007bcb9} /* (8, 23, 6) {real, imag} */,
  {32'hbfccda96, 32'h402a1319} /* (8, 23, 5) {real, imag} */,
  {32'h3d273440, 32'h3fe9606c} /* (8, 23, 4) {real, imag} */,
  {32'hbede4314, 32'h3f994940} /* (8, 23, 3) {real, imag} */,
  {32'hc012ab0c, 32'h3ff80db9} /* (8, 23, 2) {real, imag} */,
  {32'hc053ae26, 32'h40128207} /* (8, 23, 1) {real, imag} */,
  {32'hc0290bea, 32'h3fa0be16} /* (8, 23, 0) {real, imag} */,
  {32'hbf6cb19d, 32'h3fca3825} /* (8, 22, 31) {real, imag} */,
  {32'hbcf1a5c0, 32'h3fb77e34} /* (8, 22, 30) {real, imag} */,
  {32'hbe4637c4, 32'h3f6b53c6} /* (8, 22, 29) {real, imag} */,
  {32'hbfb30b9c, 32'h4019bf42} /* (8, 22, 28) {real, imag} */,
  {32'hbf895000, 32'h401b5084} /* (8, 22, 27) {real, imag} */,
  {32'hc0287db9, 32'h3ecb9570} /* (8, 22, 26) {real, imag} */,
  {32'hc0710e9a, 32'h3f48d27b} /* (8, 22, 25) {real, imag} */,
  {32'hc0366066, 32'h3eddee62} /* (8, 22, 24) {real, imag} */,
  {32'hc03c4c72, 32'h3f987504} /* (8, 22, 23) {real, imag} */,
  {32'hc04c2576, 32'h3fee1a88} /* (8, 22, 22) {real, imag} */,
  {32'h3e8346aa, 32'h3f09cd94} /* (8, 22, 21) {real, imag} */,
  {32'h40735bc6, 32'hbff5c93b} /* (8, 22, 20) {real, imag} */,
  {32'h408ab9c3, 32'hc033b629} /* (8, 22, 19) {real, imag} */,
  {32'h400b3f54, 32'hbfa3323a} /* (8, 22, 18) {real, imag} */,
  {32'h3fbbaf50, 32'hbff13b0c} /* (8, 22, 17) {real, imag} */,
  {32'h3ee015f2, 32'hc08dd978} /* (8, 22, 16) {real, imag} */,
  {32'h3ffc70d4, 32'hc0557e76} /* (8, 22, 15) {real, imag} */,
  {32'h404425ea, 32'hbf824568} /* (8, 22, 14) {real, imag} */,
  {32'h4076f892, 32'hbfe935c3} /* (8, 22, 13) {real, imag} */,
  {32'h3f967a8f, 32'hc048a4b4} /* (8, 22, 12) {real, imag} */,
  {32'h3f289662, 32'hc016f8d5} /* (8, 22, 11) {real, imag} */,
  {32'hbfe6d5b4, 32'h3fbb6627} /* (8, 22, 10) {real, imag} */,
  {32'hc03e85a5, 32'h4046cd3f} /* (8, 22, 9) {real, imag} */,
  {32'hc06128f7, 32'h406afe66} /* (8, 22, 8) {real, imag} */,
  {32'hc029e028, 32'h3fd77921} /* (8, 22, 7) {real, imag} */,
  {32'hc075eaa8, 32'h401166b9} /* (8, 22, 6) {real, imag} */,
  {32'hc043bb24, 32'h400918dd} /* (8, 22, 5) {real, imag} */,
  {32'hc00cd918, 32'h400ab2fa} /* (8, 22, 4) {real, imag} */,
  {32'hbfad91b4, 32'h3ff313a9} /* (8, 22, 3) {real, imag} */,
  {32'hc025592c, 32'h3f3d3946} /* (8, 22, 2) {real, imag} */,
  {32'hc03d5b0e, 32'h3fb5f617} /* (8, 22, 1) {real, imag} */,
  {32'hbfe42941, 32'h3ff84c7c} /* (8, 22, 0) {real, imag} */,
  {32'h3f192a4c, 32'h4007fcf3} /* (8, 21, 31) {real, imag} */,
  {32'hbe2b1aca, 32'h40113857} /* (8, 21, 30) {real, imag} */,
  {32'hbf8a26aa, 32'h3edde5b2} /* (8, 21, 29) {real, imag} */,
  {32'hbfa1639f, 32'h402b6ec0} /* (8, 21, 28) {real, imag} */,
  {32'hbf41722e, 32'h4065f7c4} /* (8, 21, 27) {real, imag} */,
  {32'hbfabe012, 32'h40165123} /* (8, 21, 26) {real, imag} */,
  {32'hbfb4c298, 32'h3f7d4e00} /* (8, 21, 25) {real, imag} */,
  {32'hbf82e7a1, 32'hbf19c0e4} /* (8, 21, 24) {real, imag} */,
  {32'hbf7d4512, 32'h3ea2d26a} /* (8, 21, 23) {real, imag} */,
  {32'hbf4c1225, 32'hbf2c9017} /* (8, 21, 22) {real, imag} */,
  {32'h3fb57cd3, 32'hbf79792c} /* (8, 21, 21) {real, imag} */,
  {32'hbe851faa, 32'hc00d1962} /* (8, 21, 20) {real, imag} */,
  {32'hbb944ac0, 32'hbfb027f2} /* (8, 21, 19) {real, imag} */,
  {32'h3e666e80, 32'h3b956180} /* (8, 21, 18) {real, imag} */,
  {32'h3ece6b32, 32'h3f467e76} /* (8, 21, 17) {real, imag} */,
  {32'hbeaecdb4, 32'hbed084fa} /* (8, 21, 16) {real, imag} */,
  {32'h3fb56476, 32'hbf5c6d02} /* (8, 21, 15) {real, imag} */,
  {32'h401dcfb0, 32'hbef6e3fa} /* (8, 21, 14) {real, imag} */,
  {32'h3ff07350, 32'hbfb43bd2} /* (8, 21, 13) {real, imag} */,
  {32'h3dd6e1a0, 32'hc05e3c28} /* (8, 21, 12) {real, imag} */,
  {32'hbf662b40, 32'hc008295e} /* (8, 21, 11) {real, imag} */,
  {32'hbef9fe4b, 32'hbd055948} /* (8, 21, 10) {real, imag} */,
  {32'hc00bed34, 32'h3fbc2528} /* (8, 21, 9) {real, imag} */,
  {32'hbfc2d176, 32'h3ece589c} /* (8, 21, 8) {real, imag} */,
  {32'hbfeab9ea, 32'h3ee5dd75} /* (8, 21, 7) {real, imag} */,
  {32'hc0817128, 32'h3fc1eb11} /* (8, 21, 6) {real, imag} */,
  {32'hc023fa59, 32'hbefae98a} /* (8, 21, 5) {real, imag} */,
  {32'hc002c59e, 32'h3deedf50} /* (8, 21, 4) {real, imag} */,
  {32'hbfd37376, 32'h3eebfa28} /* (8, 21, 3) {real, imag} */,
  {32'hbf584d54, 32'hbf9208be} /* (8, 21, 2) {real, imag} */,
  {32'hbc198d80, 32'h3f811ece} /* (8, 21, 1) {real, imag} */,
  {32'hbf24dad4, 32'h3f65f520} /* (8, 21, 0) {real, imag} */,
  {32'h3fbb0387, 32'h3f8d1a84} /* (8, 20, 31) {real, imag} */,
  {32'h3f3334a0, 32'hbda9bc90} /* (8, 20, 30) {real, imag} */,
  {32'h3f915946, 32'hbf966ece} /* (8, 20, 29) {real, imag} */,
  {32'hbf071d58, 32'h3f86ff4e} /* (8, 20, 28) {real, imag} */,
  {32'hbc3cc700, 32'h3feb42da} /* (8, 20, 27) {real, imag} */,
  {32'h400e504a, 32'h4017cffd} /* (8, 20, 26) {real, imag} */,
  {32'h40159e86, 32'h3d782680} /* (8, 20, 25) {real, imag} */,
  {32'h40112b94, 32'hc00cfe19} /* (8, 20, 24) {real, imag} */,
  {32'h400acfb8, 32'hbffbdb7f} /* (8, 20, 23) {real, imag} */,
  {32'h3ff21ed4, 32'hc08140a8} /* (8, 20, 22) {real, imag} */,
  {32'h400e89bb, 32'hc0590254} /* (8, 20, 21) {real, imag} */,
  {32'hbfa4a2e4, 32'hc02c26ef} /* (8, 20, 20) {real, imag} */,
  {32'hbffb8f27, 32'hbf09f438} /* (8, 20, 19) {real, imag} */,
  {32'hbf14e90e, 32'h3ff9fbe2} /* (8, 20, 18) {real, imag} */,
  {32'hbf4849db, 32'h40309a47} /* (8, 20, 17) {real, imag} */,
  {32'hc01366f3, 32'h405a83bf} /* (8, 20, 16) {real, imag} */,
  {32'hbfca909d, 32'h405bcba4} /* (8, 20, 15) {real, imag} */,
  {32'hbee5dbcb, 32'h40142636} /* (8, 20, 14) {real, imag} */,
  {32'hbf3c9b93, 32'h3f8eb2ce} /* (8, 20, 13) {real, imag} */,
  {32'hbf7c7ce5, 32'hbf5671c6} /* (8, 20, 12) {real, imag} */,
  {32'hbf50e62a, 32'hbdf06c60} /* (8, 20, 11) {real, imag} */,
  {32'h3f9501ee, 32'hbf7da7d8} /* (8, 20, 10) {real, imag} */,
  {32'hbe6a3920, 32'hbfb27cb8} /* (8, 20, 9) {real, imag} */,
  {32'hbecfc20a, 32'hbf9a90d3} /* (8, 20, 8) {real, imag} */,
  {32'h3f52f954, 32'hbefc5e62} /* (8, 20, 7) {real, imag} */,
  {32'h3fa18f54, 32'hc00664ea} /* (8, 20, 6) {real, imag} */,
  {32'h3e009c90, 32'hc01e7f84} /* (8, 20, 5) {real, imag} */,
  {32'h3deedff8, 32'hbfe1532e} /* (8, 20, 4) {real, imag} */,
  {32'h3fa7260f, 32'hbf8a3751} /* (8, 20, 3) {real, imag} */,
  {32'h3f442d46, 32'hbfcb4702} /* (8, 20, 2) {real, imag} */,
  {32'h4001cf46, 32'hbfa62014} /* (8, 20, 1) {real, imag} */,
  {32'h3fcda652, 32'hbf389a89} /* (8, 20, 0) {real, imag} */,
  {32'h3f472eb4, 32'h3ede304c} /* (8, 19, 31) {real, imag} */,
  {32'h3ffe46ef, 32'hbf3ecd41} /* (8, 19, 30) {real, imag} */,
  {32'h402edf5c, 32'hbf59ffa8} /* (8, 19, 29) {real, imag} */,
  {32'h3e94702c, 32'hbce992c0} /* (8, 19, 28) {real, imag} */,
  {32'h3f458dc1, 32'hbf753bbe} /* (8, 19, 27) {real, imag} */,
  {32'h3febc7a1, 32'hc0002af8} /* (8, 19, 26) {real, imag} */,
  {32'h3fcceac6, 32'hbff911e0} /* (8, 19, 25) {real, imag} */,
  {32'h401f1bc0, 32'hbfc66b80} /* (8, 19, 24) {real, imag} */,
  {32'h4046ef40, 32'hc0364ca9} /* (8, 19, 23) {real, imag} */,
  {32'h40586cba, 32'hc024dae9} /* (8, 19, 22) {real, imag} */,
  {32'h402e6326, 32'hbfc1c319} /* (8, 19, 21) {real, imag} */,
  {32'h3f4c68c1, 32'hbfb5d1e1} /* (8, 19, 20) {real, imag} */,
  {32'hbfebef17, 32'hbf737aa9} /* (8, 19, 19) {real, imag} */,
  {32'hbfe89754, 32'h3faa8b1c} /* (8, 19, 18) {real, imag} */,
  {32'hc03f4516, 32'h404f3385} /* (8, 19, 17) {real, imag} */,
  {32'hc0646340, 32'h408a2f60} /* (8, 19, 16) {real, imag} */,
  {32'hc02be56e, 32'h40a842e2} /* (8, 19, 15) {real, imag} */,
  {32'hbfce11e6, 32'h40583aee} /* (8, 19, 14) {real, imag} */,
  {32'hbf877872, 32'h40483d30} /* (8, 19, 13) {real, imag} */,
  {32'hc00cb08e, 32'h3f90c8f3} /* (8, 19, 12) {real, imag} */,
  {32'hc0127bcc, 32'hbeb257e0} /* (8, 19, 11) {real, imag} */,
  {32'h3f7f3ba0, 32'hbfe58341} /* (8, 19, 10) {real, imag} */,
  {32'h3eac64a8, 32'hbfc9c229} /* (8, 19, 9) {real, imag} */,
  {32'hbf11e529, 32'hbe81c3e8} /* (8, 19, 8) {real, imag} */,
  {32'h3f3d65cf, 32'h3f5a5f84} /* (8, 19, 7) {real, imag} */,
  {32'h3fe12e96, 32'hbf8a50f0} /* (8, 19, 6) {real, imag} */,
  {32'h3fb302d3, 32'hbf7d4f39} /* (8, 19, 5) {real, imag} */,
  {32'h401efe2a, 32'hbfe95713} /* (8, 19, 4) {real, imag} */,
  {32'h3faa1d24, 32'hc0395ad5} /* (8, 19, 3) {real, imag} */,
  {32'hbf0a9a04, 32'hc001f870} /* (8, 19, 2) {real, imag} */,
  {32'h401ddc20, 32'hbf319c40} /* (8, 19, 1) {real, imag} */,
  {32'h3fec42f4, 32'h3de893d0} /* (8, 19, 0) {real, imag} */,
  {32'h3f0d929c, 32'hbf2527d4} /* (8, 18, 31) {real, imag} */,
  {32'h3ea94c1c, 32'hbfb1ee29} /* (8, 18, 30) {real, imag} */,
  {32'hbd10be00, 32'hbfc090ed} /* (8, 18, 29) {real, imag} */,
  {32'h3e3f85aa, 32'hbfc42553} /* (8, 18, 28) {real, imag} */,
  {32'h3f837958, 32'hc020cf72} /* (8, 18, 27) {real, imag} */,
  {32'h3e78bcd8, 32'hc014773e} /* (8, 18, 26) {real, imag} */,
  {32'h3ef8958c, 32'hbfdd6a52} /* (8, 18, 25) {real, imag} */,
  {32'h406d8dd2, 32'hbe936024} /* (8, 18, 24) {real, imag} */,
  {32'h3fce7c08, 32'hc0170e36} /* (8, 18, 23) {real, imag} */,
  {32'h3fa11014, 32'hbfec940e} /* (8, 18, 22) {real, imag} */,
  {32'h4030189e, 32'h3fac2285} /* (8, 18, 21) {real, imag} */,
  {32'h3edaa36e, 32'hbfb5a752} /* (8, 18, 20) {real, imag} */,
  {32'hbfc68f5a, 32'hbed1fe64} /* (8, 18, 19) {real, imag} */,
  {32'hbece286c, 32'h3fb94988} /* (8, 18, 18) {real, imag} */,
  {32'hc05b19ab, 32'h405047d1} /* (8, 18, 17) {real, imag} */,
  {32'hc02c2cb7, 32'h402c4176} /* (8, 18, 16) {real, imag} */,
  {32'hc012a841, 32'h4013cf91} /* (8, 18, 15) {real, imag} */,
  {32'hbf9d138e, 32'h3fa2ae92} /* (8, 18, 14) {real, imag} */,
  {32'hbf7e5dd8, 32'h40111b62} /* (8, 18, 13) {real, imag} */,
  {32'hbf4ba73f, 32'h3d37f3d0} /* (8, 18, 12) {real, imag} */,
  {32'hbfb99ff3, 32'hbf6d1c9d} /* (8, 18, 11) {real, imag} */,
  {32'h4015b803, 32'hbf109e1b} /* (8, 18, 10) {real, imag} */,
  {32'h3fdbc64d, 32'hbf178c22} /* (8, 18, 9) {real, imag} */,
  {32'h3f14f499, 32'hbfac21b8} /* (8, 18, 8) {real, imag} */,
  {32'h3f426eee, 32'hc04cc86f} /* (8, 18, 7) {real, imag} */,
  {32'h4012f465, 32'hc07d8850} /* (8, 18, 6) {real, imag} */,
  {32'h405e62d1, 32'hbfce0c86} /* (8, 18, 5) {real, imag} */,
  {32'h4070957c, 32'h3f1fbbc6} /* (8, 18, 4) {real, imag} */,
  {32'h3ffbfe46, 32'hbf887961} /* (8, 18, 3) {real, imag} */,
  {32'hbf4f577a, 32'hc01c9248} /* (8, 18, 2) {real, imag} */,
  {32'h40135098, 32'hbf0d1c2d} /* (8, 18, 1) {real, imag} */,
  {32'h401274ea, 32'h3f879d46} /* (8, 18, 0) {real, imag} */,
  {32'h3f550cda, 32'h3ed465ae} /* (8, 17, 31) {real, imag} */,
  {32'hbf03c1cc, 32'hbf102b78} /* (8, 17, 30) {real, imag} */,
  {32'hbfc15ea5, 32'hbed01c90} /* (8, 17, 29) {real, imag} */,
  {32'h3c8bf200, 32'hbec6089a} /* (8, 17, 28) {real, imag} */,
  {32'h40071424, 32'hbfc62591} /* (8, 17, 27) {real, imag} */,
  {32'h3fbc5da1, 32'hbf9da03b} /* (8, 17, 26) {real, imag} */,
  {32'h4028afe6, 32'hc0432088} /* (8, 17, 25) {real, imag} */,
  {32'h40495904, 32'hc0152b9e} /* (8, 17, 24) {real, imag} */,
  {32'hbf9044b9, 32'hc039e5ca} /* (8, 17, 23) {real, imag} */,
  {32'h3fdd40ae, 32'hbffc5d1e} /* (8, 17, 22) {real, imag} */,
  {32'h4055c3a4, 32'hbf6b4244} /* (8, 17, 21) {real, imag} */,
  {32'hbe81addc, 32'hbf95d64c} /* (8, 17, 20) {real, imag} */,
  {32'hbff9a458, 32'h3ffb96a3} /* (8, 17, 19) {real, imag} */,
  {32'hbf966340, 32'h4080510e} /* (8, 17, 18) {real, imag} */,
  {32'hc024b22c, 32'h4048c814} /* (8, 17, 17) {real, imag} */,
  {32'hc03c0316, 32'h3f057412} /* (8, 17, 16) {real, imag} */,
  {32'hc066fa88, 32'h3e36fe60} /* (8, 17, 15) {real, imag} */,
  {32'hc0467a48, 32'h3fb25e39} /* (8, 17, 14) {real, imag} */,
  {32'hbfe3a2a6, 32'h40294086} /* (8, 17, 13) {real, imag} */,
  {32'hbf878f43, 32'h3fc683b5} /* (8, 17, 12) {real, imag} */,
  {32'hbfc8e971, 32'hbeb18f5c} /* (8, 17, 11) {real, imag} */,
  {32'h4050e823, 32'hc05b8dd3} /* (8, 17, 10) {real, imag} */,
  {32'h403d4a6b, 32'hc00d8286} /* (8, 17, 9) {real, imag} */,
  {32'h3f23675c, 32'hbfd2c556} /* (8, 17, 8) {real, imag} */,
  {32'h3ecf2cf2, 32'hc0499ee7} /* (8, 17, 7) {real, imag} */,
  {32'h3fca6ec1, 32'hc08e491c} /* (8, 17, 6) {real, imag} */,
  {32'h4080e41c, 32'hc04800aa} /* (8, 17, 5) {real, imag} */,
  {32'h402fbc78, 32'hbf574382} /* (8, 17, 4) {real, imag} */,
  {32'h3f6aac10, 32'hc0229ee0} /* (8, 17, 3) {real, imag} */,
  {32'h3ffd9650, 32'hc05dc63a} /* (8, 17, 2) {real, imag} */,
  {32'h406fbdeb, 32'hc0140f37} /* (8, 17, 1) {real, imag} */,
  {32'h401b617e, 32'hbe85ee08} /* (8, 17, 0) {real, imag} */,
  {32'h3d2aba20, 32'hbe391dbc} /* (8, 16, 31) {real, imag} */,
  {32'hbdefd530, 32'hbf484c5b} /* (8, 16, 30) {real, imag} */,
  {32'h3fca8cf3, 32'hbfb2015d} /* (8, 16, 29) {real, imag} */,
  {32'h3f7e60ab, 32'hbfad0237} /* (8, 16, 28) {real, imag} */,
  {32'h403f1a06, 32'hbf0e60a7} /* (8, 16, 27) {real, imag} */,
  {32'h3f7e632a, 32'hc011c2a0} /* (8, 16, 26) {real, imag} */,
  {32'h3f8e5ad4, 32'hc045d01e} /* (8, 16, 25) {real, imag} */,
  {32'h3fb9feac, 32'hbfd3706e} /* (8, 16, 24) {real, imag} */,
  {32'hbe03d54c, 32'hc01650e8} /* (8, 16, 23) {real, imag} */,
  {32'h4006a772, 32'hc0096410} /* (8, 16, 22) {real, imag} */,
  {32'h3fb9f30a, 32'hbfc52de0} /* (8, 16, 21) {real, imag} */,
  {32'hbe5292f0, 32'hbf5c1c97} /* (8, 16, 20) {real, imag} */,
  {32'hc01d4e98, 32'h4025ef0e} /* (8, 16, 19) {real, imag} */,
  {32'hbf257b53, 32'h40164501} /* (8, 16, 18) {real, imag} */,
  {32'hbf868a00, 32'h3f280162} /* (8, 16, 17) {real, imag} */,
  {32'hc03e7f05, 32'hbf008212} /* (8, 16, 16) {real, imag} */,
  {32'hc04b4340, 32'hbee1d428} /* (8, 16, 15) {real, imag} */,
  {32'hc06c4866, 32'h3fe0a58a} /* (8, 16, 14) {real, imag} */,
  {32'hc03eca37, 32'h404c91d8} /* (8, 16, 13) {real, imag} */,
  {32'hc06d6552, 32'h40203290} /* (8, 16, 12) {real, imag} */,
  {32'hc00ddd5c, 32'h3f012fa0} /* (8, 16, 11) {real, imag} */,
  {32'h3ff6f2f8, 32'hc0525d22} /* (8, 16, 10) {real, imag} */,
  {32'h401663ea, 32'hc03d17e1} /* (8, 16, 9) {real, imag} */,
  {32'h3ffc8c41, 32'hc00a9d06} /* (8, 16, 8) {real, imag} */,
  {32'h3ff0ff14, 32'hc05d3610} /* (8, 16, 7) {real, imag} */,
  {32'h3f77c1ac, 32'hc0b7c6ce} /* (8, 16, 6) {real, imag} */,
  {32'h403d3d4c, 32'hc06a9e28} /* (8, 16, 5) {real, imag} */,
  {32'h40166dce, 32'hc00d5ae2} /* (8, 16, 4) {real, imag} */,
  {32'h4005e4ea, 32'hbfda93a6} /* (8, 16, 3) {real, imag} */,
  {32'h409fcbf8, 32'hbfe2e62c} /* (8, 16, 2) {real, imag} */,
  {32'h40424c5b, 32'hc03e4ce0} /* (8, 16, 1) {real, imag} */,
  {32'h3f9638dc, 32'hc00c7a43} /* (8, 16, 0) {real, imag} */,
  {32'h3ea1fee2, 32'hbf60a4fd} /* (8, 15, 31) {real, imag} */,
  {32'h40079e42, 32'hc0023428} /* (8, 15, 30) {real, imag} */,
  {32'h40792916, 32'hc05fd0b0} /* (8, 15, 29) {real, imag} */,
  {32'h40129747, 32'hc0302756} /* (8, 15, 28) {real, imag} */,
  {32'h40389a07, 32'hbfc2aadf} /* (8, 15, 27) {real, imag} */,
  {32'h3f8206d2, 32'hc0415238} /* (8, 15, 26) {real, imag} */,
  {32'h3f0a2028, 32'hc0314342} /* (8, 15, 25) {real, imag} */,
  {32'hbfb51689, 32'hbf1c9cbb} /* (8, 15, 24) {real, imag} */,
  {32'h3fc28ead, 32'hbf43b62a} /* (8, 15, 23) {real, imag} */,
  {32'h4020812c, 32'hbfac925a} /* (8, 15, 22) {real, imag} */,
  {32'h3f26f538, 32'hbef12188} /* (8, 15, 21) {real, imag} */,
  {32'hbf9e35cc, 32'hbec8c992} /* (8, 15, 20) {real, imag} */,
  {32'hc0296e24, 32'h3f853953} /* (8, 15, 19) {real, imag} */,
  {32'h3f01480b, 32'h3f98a9a1} /* (8, 15, 18) {real, imag} */,
  {32'h3fcdee00, 32'h3fa53c21} /* (8, 15, 17) {real, imag} */,
  {32'hc000dfae, 32'h3f8140bf} /* (8, 15, 16) {real, imag} */,
  {32'hc058c865, 32'h3fbb662b} /* (8, 15, 15) {real, imag} */,
  {32'hc049ab4e, 32'h3fb9b99b} /* (8, 15, 14) {real, imag} */,
  {32'hc02465c0, 32'h40321b74} /* (8, 15, 13) {real, imag} */,
  {32'hbfe5ed86, 32'h40033502} /* (8, 15, 12) {real, imag} */,
  {32'hbe16c150, 32'h3f9587f8} /* (8, 15, 11) {real, imag} */,
  {32'h3fffa1d5, 32'hbffc36a0} /* (8, 15, 10) {real, imag} */,
  {32'h402b1e80, 32'hc080e82e} /* (8, 15, 9) {real, imag} */,
  {32'h3f92b804, 32'hbf8ef401} /* (8, 15, 8) {real, imag} */,
  {32'h3ee8fa48, 32'hbeb6a368} /* (8, 15, 7) {real, imag} */,
  {32'h3fd26ddc, 32'hc01605f0} /* (8, 15, 6) {real, imag} */,
  {32'h4078a8c5, 32'hc0249826} /* (8, 15, 5) {real, imag} */,
  {32'h401fc872, 32'hc07630f8} /* (8, 15, 4) {real, imag} */,
  {32'h4071a139, 32'hbfee5b58} /* (8, 15, 3) {real, imag} */,
  {32'h40b8b2f0, 32'hbfd10475} /* (8, 15, 2) {real, imag} */,
  {32'h4018c947, 32'hc0655f61} /* (8, 15, 1) {real, imag} */,
  {32'hbc949be0, 32'hbf3716a2} /* (8, 15, 0) {real, imag} */,
  {32'h3f42d5d8, 32'hbf7c4e8a} /* (8, 14, 31) {real, imag} */,
  {32'h3ff2f50e, 32'hc07a4872} /* (8, 14, 30) {real, imag} */,
  {32'h4043ec25, 32'hc0b80fde} /* (8, 14, 29) {real, imag} */,
  {32'h404a5f03, 32'hc06a98b2} /* (8, 14, 28) {real, imag} */,
  {32'h401e01cf, 32'hc0631799} /* (8, 14, 27) {real, imag} */,
  {32'h3ee046ac, 32'hc07f5108} /* (8, 14, 26) {real, imag} */,
  {32'h3f8e1a83, 32'hc052e1ac} /* (8, 14, 25) {real, imag} */,
  {32'h3f4aaf18, 32'h3f2d0964} /* (8, 14, 24) {real, imag} */,
  {32'h3ff61fc7, 32'h3eb7b048} /* (8, 14, 23) {real, imag} */,
  {32'h3f4d856c, 32'hbfafc050} /* (8, 14, 22) {real, imag} */,
  {32'hbd09f490, 32'hbfc6e1c0} /* (8, 14, 21) {real, imag} */,
  {32'hc0296a11, 32'h3e3047a0} /* (8, 14, 20) {real, imag} */,
  {32'hc01a6d02, 32'h401b5df4} /* (8, 14, 19) {real, imag} */,
  {32'hbe4ee388, 32'h405fbf78} /* (8, 14, 18) {real, imag} */,
  {32'hbf0621f8, 32'h403a4cf8} /* (8, 14, 17) {real, imag} */,
  {32'hbfcd0e82, 32'h3f9a7f62} /* (8, 14, 16) {real, imag} */,
  {32'hbffe2876, 32'h40272b0a} /* (8, 14, 15) {real, imag} */,
  {32'hbf71b7fc, 32'h3ffe24ae} /* (8, 14, 14) {real, imag} */,
  {32'hbf85bbdc, 32'h40349d82} /* (8, 14, 13) {real, imag} */,
  {32'hbf1b9233, 32'h40448604} /* (8, 14, 12) {real, imag} */,
  {32'hbe3fe4f0, 32'h3fde4db1} /* (8, 14, 11) {real, imag} */,
  {32'h3fe1920b, 32'hbdf01b8c} /* (8, 14, 10) {real, imag} */,
  {32'h3fedfe54, 32'hbfd27c9e} /* (8, 14, 9) {real, imag} */,
  {32'h3ddbeb38, 32'hbfca51d6} /* (8, 14, 8) {real, imag} */,
  {32'hbd851318, 32'hbfecf4b2} /* (8, 14, 7) {real, imag} */,
  {32'h40199e7d, 32'hbf9eb2fb} /* (8, 14, 6) {real, imag} */,
  {32'h409f99e7, 32'hbf96a133} /* (8, 14, 5) {real, imag} */,
  {32'h405e64be, 32'hc02f8947} /* (8, 14, 4) {real, imag} */,
  {32'h400fdc76, 32'hbfb78f4c} /* (8, 14, 3) {real, imag} */,
  {32'h3f493394, 32'hc013b9e4} /* (8, 14, 2) {real, imag} */,
  {32'hbf2d41b2, 32'hc043ef4a} /* (8, 14, 1) {real, imag} */,
  {32'hbf8bc9a6, 32'h3ef40ae9} /* (8, 14, 0) {real, imag} */,
  {32'h3e125e98, 32'hbfa9c622} /* (8, 13, 31) {real, imag} */,
  {32'h3e66ba5c, 32'hc047e717} /* (8, 13, 30) {real, imag} */,
  {32'h3f55bfe4, 32'hc05fe2ba} /* (8, 13, 29) {real, imag} */,
  {32'h3fc77d9c, 32'hc01763d8} /* (8, 13, 28) {real, imag} */,
  {32'h40774740, 32'hc0836a73} /* (8, 13, 27) {real, imag} */,
  {32'h4005dcf9, 32'hc0879b2c} /* (8, 13, 26) {real, imag} */,
  {32'h3fd6f842, 32'hc03c1e33} /* (8, 13, 25) {real, imag} */,
  {32'h4062e27e, 32'hbee16bbc} /* (8, 13, 24) {real, imag} */,
  {32'h401f6c7e, 32'hbfed872e} /* (8, 13, 23) {real, imag} */,
  {32'h3ebf8baa, 32'hc088236a} /* (8, 13, 22) {real, imag} */,
  {32'h3f80551b, 32'hc015ed22} /* (8, 13, 21) {real, imag} */,
  {32'hc006070e, 32'hbeddc5c2} /* (8, 13, 20) {real, imag} */,
  {32'hc0241084, 32'h40038140} /* (8, 13, 19) {real, imag} */,
  {32'hbfd8f870, 32'h40710cb0} /* (8, 13, 18) {real, imag} */,
  {32'hbf8deec4, 32'h4040ece9} /* (8, 13, 17) {real, imag} */,
  {32'h3eaedff4, 32'h40805316} /* (8, 13, 16) {real, imag} */,
  {32'h3e32d778, 32'h40476776} /* (8, 13, 15) {real, imag} */,
  {32'h3f7967d3, 32'h3fed3de6} /* (8, 13, 14) {real, imag} */,
  {32'hbfe64bbe, 32'h3b8ed180} /* (8, 13, 13) {real, imag} */,
  {32'hbfedabd1, 32'h3f7efcbb} /* (8, 13, 12) {real, imag} */,
  {32'hbfc6e250, 32'h3fd3370e} /* (8, 13, 11) {real, imag} */,
  {32'hbe5236ec, 32'hbeafa781} /* (8, 13, 10) {real, imag} */,
  {32'h3f8a2938, 32'hc0043c91} /* (8, 13, 9) {real, imag} */,
  {32'h3ffe9ac7, 32'hc0319b00} /* (8, 13, 8) {real, imag} */,
  {32'h4066e5d6, 32'hbfde31f2} /* (8, 13, 7) {real, imag} */,
  {32'h405d3ac2, 32'hc014fd16} /* (8, 13, 6) {real, imag} */,
  {32'h40286ffc, 32'hbffe1d46} /* (8, 13, 5) {real, imag} */,
  {32'h40683378, 32'hc0251810} /* (8, 13, 4) {real, imag} */,
  {32'h4060a390, 32'hbfed1e3b} /* (8, 13, 3) {real, imag} */,
  {32'h3eeedf60, 32'hc03a70bc} /* (8, 13, 2) {real, imag} */,
  {32'h3d905840, 32'hbfc9c2b8} /* (8, 13, 1) {real, imag} */,
  {32'hbdf19b00, 32'hbf01e73f} /* (8, 13, 0) {real, imag} */,
  {32'h3f30e725, 32'hc0011c2c} /* (8, 12, 31) {real, imag} */,
  {32'h3faa9ce7, 32'hbff43e04} /* (8, 12, 30) {real, imag} */,
  {32'h3f405386, 32'hbf86c499} /* (8, 12, 29) {real, imag} */,
  {32'hbf67b75c, 32'hbf88145a} /* (8, 12, 28) {real, imag} */,
  {32'h3fcbdf9b, 32'hbfe4ac86} /* (8, 12, 27) {real, imag} */,
  {32'h4028326e, 32'hc0020680} /* (8, 12, 26) {real, imag} */,
  {32'h3ff93417, 32'hc076634a} /* (8, 12, 25) {real, imag} */,
  {32'h402a9670, 32'hc0626580} /* (8, 12, 24) {real, imag} */,
  {32'h3fd80655, 32'hc08a9b33} /* (8, 12, 23) {real, imag} */,
  {32'h401f903c, 32'hc0935b13} /* (8, 12, 22) {real, imag} */,
  {32'h4061fdfc, 32'hbfd09ff0} /* (8, 12, 21) {real, imag} */,
  {32'h3e945e2e, 32'h3bc22f00} /* (8, 12, 20) {real, imag} */,
  {32'hc00895ca, 32'h3ec2fd78} /* (8, 12, 19) {real, imag} */,
  {32'hc0083d6b, 32'h40147b36} /* (8, 12, 18) {real, imag} */,
  {32'hc00266a8, 32'h40341daa} /* (8, 12, 17) {real, imag} */,
  {32'hbf51ee04, 32'h40559df2} /* (8, 12, 16) {real, imag} */,
  {32'hbf67fecc, 32'h3ffa6384} /* (8, 12, 15) {real, imag} */,
  {32'hbed50a88, 32'h40002d01} /* (8, 12, 14) {real, imag} */,
  {32'hc022f4ee, 32'hbcbf48e0} /* (8, 12, 13) {real, imag} */,
  {32'hbff67c90, 32'h3e849d28} /* (8, 12, 12) {real, imag} */,
  {32'h3eb48870, 32'h3f5bc556} /* (8, 12, 11) {real, imag} */,
  {32'h3faed33a, 32'hc0145a06} /* (8, 12, 10) {real, imag} */,
  {32'h3fd921be, 32'hc00364ee} /* (8, 12, 9) {real, imag} */,
  {32'h40299991, 32'hbff6a152} /* (8, 12, 8) {real, imag} */,
  {32'h400a4f7b, 32'hbf8715d4} /* (8, 12, 7) {real, imag} */,
  {32'h3fc6fd31, 32'hc00d7ee4} /* (8, 12, 6) {real, imag} */,
  {32'h3f194286, 32'hc031bd0a} /* (8, 12, 5) {real, imag} */,
  {32'h4021f3f2, 32'hc03e90e4} /* (8, 12, 4) {real, imag} */,
  {32'h3fceeaa1, 32'hbf886f30} /* (8, 12, 3) {real, imag} */,
  {32'h3fdfb464, 32'hbf52b928} /* (8, 12, 2) {real, imag} */,
  {32'h3fec5a98, 32'hbf8192c9} /* (8, 12, 1) {real, imag} */,
  {32'h3f7e03c5, 32'hbf8fdc82} /* (8, 12, 0) {real, imag} */,
  {32'h3bab4200, 32'hbfd79722} /* (8, 11, 31) {real, imag} */,
  {32'h3f926dd8, 32'hbfc2f820} /* (8, 11, 30) {real, imag} */,
  {32'h40371931, 32'hbf86c480} /* (8, 11, 29) {real, imag} */,
  {32'h400b1bf2, 32'hbafd5800} /* (8, 11, 28) {real, imag} */,
  {32'h3ff9b382, 32'h3ef44294} /* (8, 11, 27) {real, imag} */,
  {32'h402b4dce, 32'hbe6c5640} /* (8, 11, 26) {real, imag} */,
  {32'h3ff69f20, 32'hc0563b15} /* (8, 11, 25) {real, imag} */,
  {32'h3efd28e2, 32'hc04663b6} /* (8, 11, 24) {real, imag} */,
  {32'h3f81c942, 32'hc08b8e35} /* (8, 11, 23) {real, imag} */,
  {32'h402a6b5a, 32'hc0871c47} /* (8, 11, 22) {real, imag} */,
  {32'h401f703a, 32'h3eaa71a4} /* (8, 11, 21) {real, imag} */,
  {32'hbed37b6c, 32'h3f93e50e} /* (8, 11, 20) {real, imag} */,
  {32'hbfe35caa, 32'hbe13a91c} /* (8, 11, 19) {real, imag} */,
  {32'hc04d9881, 32'h40138ea0} /* (8, 11, 18) {real, imag} */,
  {32'hc084c2af, 32'h402cd2ae} /* (8, 11, 17) {real, imag} */,
  {32'hc011ba02, 32'h4040440c} /* (8, 11, 16) {real, imag} */,
  {32'hbfe0672e, 32'h3feffb46} /* (8, 11, 15) {real, imag} */,
  {32'hbbeb9c80, 32'h3fa94e60} /* (8, 11, 14) {real, imag} */,
  {32'h3ee2dad4, 32'hbe4cf1f4} /* (8, 11, 13) {real, imag} */,
  {32'hbea2ce6d, 32'h3faf044e} /* (8, 11, 12) {real, imag} */,
  {32'h3f0250d5, 32'h4002400e} /* (8, 11, 11) {real, imag} */,
  {32'h3f22bae1, 32'hbf11e448} /* (8, 11, 10) {real, imag} */,
  {32'h3f8d79e6, 32'hbf122e74} /* (8, 11, 9) {real, imag} */,
  {32'h3eafb5b0, 32'hc0038ac4} /* (8, 11, 8) {real, imag} */,
  {32'hbf45d808, 32'hbfd757fc} /* (8, 11, 7) {real, imag} */,
  {32'h3f48b6ea, 32'hbfb7ba70} /* (8, 11, 6) {real, imag} */,
  {32'h3f1cd990, 32'hc076cfa7} /* (8, 11, 5) {real, imag} */,
  {32'h3e903ea8, 32'hc01142eb} /* (8, 11, 4) {real, imag} */,
  {32'h3f957454, 32'h3d7f47b0} /* (8, 11, 3) {real, imag} */,
  {32'h3f27e993, 32'h3e9c5fce} /* (8, 11, 2) {real, imag} */,
  {32'hbdc95e58, 32'hc016f962} /* (8, 11, 1) {real, imag} */,
  {32'hbe4af45c, 32'hbff5afc9} /* (8, 11, 0) {real, imag} */,
  {32'hbf5ade30, 32'hbf5dfa30} /* (8, 10, 31) {real, imag} */,
  {32'hbfce97f7, 32'hbf154d00} /* (8, 10, 30) {real, imag} */,
  {32'hbf98c817, 32'hbe8e0ba6} /* (8, 10, 29) {real, imag} */,
  {32'hbdde2d30, 32'hbecd1302} /* (8, 10, 28) {real, imag} */,
  {32'hbf9d8ffa, 32'h3efc3498} /* (8, 10, 27) {real, imag} */,
  {32'hbfb6d8e0, 32'h3fc00ab1} /* (8, 10, 26) {real, imag} */,
  {32'h3e202e80, 32'h3f88e666} /* (8, 10, 25) {real, imag} */,
  {32'hbe3fab04, 32'hbfc9f762} /* (8, 10, 24) {real, imag} */,
  {32'hbf7575b1, 32'hc0289f0e} /* (8, 10, 23) {real, imag} */,
  {32'hbf857610, 32'h3ea0adae} /* (8, 10, 22) {real, imag} */,
  {32'hbf67790c, 32'h40785870} /* (8, 10, 21) {real, imag} */,
  {32'hbdec76a0, 32'h3ea65db0} /* (8, 10, 20) {real, imag} */,
  {32'h3fc6a52f, 32'hc00afe52} /* (8, 10, 19) {real, imag} */,
  {32'hbefcc588, 32'h3fcbe24b} /* (8, 10, 18) {real, imag} */,
  {32'hbf681bc4, 32'h3e7a8e18} /* (8, 10, 17) {real, imag} */,
  {32'h3fba3a39, 32'hbecd2406} /* (8, 10, 16) {real, imag} */,
  {32'h3ffabc42, 32'hbfa2661f} /* (8, 10, 15) {real, imag} */,
  {32'h3fc931e4, 32'hbe8594e9} /* (8, 10, 14) {real, imag} */,
  {32'h3f1c0996, 32'hbfee0d6c} /* (8, 10, 13) {real, imag} */,
  {32'h3f28f448, 32'h3eac4ba6} /* (8, 10, 12) {real, imag} */,
  {32'hbf009212, 32'hbf2363c6} /* (8, 10, 11) {real, imag} */,
  {32'hbe6ab3cc, 32'h3f239800} /* (8, 10, 10) {real, imag} */,
  {32'hbf8eae55, 32'h405b2a05} /* (8, 10, 9) {real, imag} */,
  {32'hc0017c80, 32'h40272fb7} /* (8, 10, 8) {real, imag} */,
  {32'hc04029c9, 32'h40088d1c} /* (8, 10, 7) {real, imag} */,
  {32'hbffadb42, 32'h3fb1a245} /* (8, 10, 6) {real, imag} */,
  {32'hbf1e90ff, 32'hbe726d00} /* (8, 10, 5) {real, imag} */,
  {32'hbfb8b534, 32'hbf3a77de} /* (8, 10, 4) {real, imag} */,
  {32'hbfe30a22, 32'hbf99c7f8} /* (8, 10, 3) {real, imag} */,
  {32'hc00f46ea, 32'h3fa13f50} /* (8, 10, 2) {real, imag} */,
  {32'hbf8f116c, 32'h3fd18ea0} /* (8, 10, 1) {real, imag} */,
  {32'hbf533350, 32'h3ea7a952} /* (8, 10, 0) {real, imag} */,
  {32'h3d9c4128, 32'h3fa5c0c2} /* (8, 9, 31) {real, imag} */,
  {32'hc001dc16, 32'h3f10c832} /* (8, 9, 30) {real, imag} */,
  {32'hc0265af9, 32'hbcaabe80} /* (8, 9, 29) {real, imag} */,
  {32'hc01abbc7, 32'hbe7ff190} /* (8, 9, 28) {real, imag} */,
  {32'hc0848f46, 32'h3f4a28fb} /* (8, 9, 27) {real, imag} */,
  {32'hc0450942, 32'h40164118} /* (8, 9, 26) {real, imag} */,
  {32'hbdce2358, 32'h4012603a} /* (8, 9, 25) {real, imag} */,
  {32'hbeb1d9d8, 32'h3eb11464} /* (8, 9, 24) {real, imag} */,
  {32'hc014786e, 32'h3e041d00} /* (8, 9, 23) {real, imag} */,
  {32'hc03774fc, 32'h4065a411} /* (8, 9, 22) {real, imag} */,
  {32'hc0000426, 32'h4080bf08} /* (8, 9, 21) {real, imag} */,
  {32'h3fa7a90e, 32'hbf432c90} /* (8, 9, 20) {real, imag} */,
  {32'h40299260, 32'hc026f6da} /* (8, 9, 19) {real, imag} */,
  {32'h3fd75553, 32'h3ec7c3da} /* (8, 9, 18) {real, imag} */,
  {32'h3fde3f4f, 32'h3ec9642a} /* (8, 9, 17) {real, imag} */,
  {32'h4047865e, 32'hbfa58fdf} /* (8, 9, 16) {real, imag} */,
  {32'h4027a8e8, 32'hbff24afe} /* (8, 9, 15) {real, imag} */,
  {32'h4009283e, 32'h3edf1200} /* (8, 9, 14) {real, imag} */,
  {32'hbef4af40, 32'hbf6eb45c} /* (8, 9, 13) {real, imag} */,
  {32'h3fcb2eb6, 32'h3fdae580} /* (8, 9, 12) {real, imag} */,
  {32'h3fbda60e, 32'hbf34c9c3} /* (8, 9, 11) {real, imag} */,
  {32'h3e941183, 32'hbf51f754} /* (8, 9, 10) {real, imag} */,
  {32'hbf9b1c0e, 32'h402e374a} /* (8, 9, 9) {real, imag} */,
  {32'hc040784e, 32'h408a3750} /* (8, 9, 8) {real, imag} */,
  {32'hc06384bd, 32'h406283a4} /* (8, 9, 7) {real, imag} */,
  {32'hc003bc94, 32'h3ff30a9e} /* (8, 9, 6) {real, imag} */,
  {32'hbfa45eb7, 32'h3fb12a46} /* (8, 9, 5) {real, imag} */,
  {32'hbeb2e716, 32'h3f914973} /* (8, 9, 4) {real, imag} */,
  {32'hbfed8272, 32'h3e559048} /* (8, 9, 3) {real, imag} */,
  {32'hc04ac0ff, 32'h401a7df4} /* (8, 9, 2) {real, imag} */,
  {32'hbfea47c2, 32'h40539c46} /* (8, 9, 1) {real, imag} */,
  {32'hbeff1ce8, 32'h3ff6e7e4} /* (8, 9, 0) {real, imag} */,
  {32'h3f669044, 32'h3c9ad070} /* (8, 8, 31) {real, imag} */,
  {32'h3e4a7e9a, 32'h3f5fdb60} /* (8, 8, 30) {real, imag} */,
  {32'hbf20d376, 32'h3fbce18c} /* (8, 8, 29) {real, imag} */,
  {32'hbecb38de, 32'h3fd745a8} /* (8, 8, 28) {real, imag} */,
  {32'hbfd097e7, 32'h3f80b27d} /* (8, 8, 27) {real, imag} */,
  {32'hbfd174b4, 32'h401d2b2a} /* (8, 8, 26) {real, imag} */,
  {32'hbf35f0c0, 32'h4081e25a} /* (8, 8, 25) {real, imag} */,
  {32'h3f7a41bc, 32'h3f89e0b0} /* (8, 8, 24) {real, imag} */,
  {32'hbf845c45, 32'h3f83b85e} /* (8, 8, 23) {real, imag} */,
  {32'hc0429d8c, 32'h40827548} /* (8, 8, 22) {real, imag} */,
  {32'hbf1397ad, 32'h400ef4c6} /* (8, 8, 21) {real, imag} */,
  {32'h3fae22a6, 32'hbf5d3c46} /* (8, 8, 20) {real, imag} */,
  {32'h3fece4c2, 32'hbfbedc8c} /* (8, 8, 19) {real, imag} */,
  {32'h3ed8975c, 32'hc0108263} /* (8, 8, 18) {real, imag} */,
  {32'h3f86cc18, 32'hc01b2aec} /* (8, 8, 17) {real, imag} */,
  {32'h4068480f, 32'hc0508222} /* (8, 8, 16) {real, imag} */,
  {32'h4041954e, 32'hc01bcced} /* (8, 8, 15) {real, imag} */,
  {32'h4038cca2, 32'hbd36d380} /* (8, 8, 14) {real, imag} */,
  {32'h40456649, 32'h3e7fe214} /* (8, 8, 13) {real, imag} */,
  {32'h40840a10, 32'h3f2fe880} /* (8, 8, 12) {real, imag} */,
  {32'h40449c99, 32'hbf6bfaf7} /* (8, 8, 11) {real, imag} */,
  {32'h3fcdcba4, 32'hbf698e62} /* (8, 8, 10) {real, imag} */,
  {32'h3eb1078d, 32'h3f62e16a} /* (8, 8, 9) {real, imag} */,
  {32'hbfc8b6d0, 32'h3f984370} /* (8, 8, 8) {real, imag} */,
  {32'hc080497e, 32'h3f14cdbb} /* (8, 8, 7) {real, imag} */,
  {32'hc06455a1, 32'h3fabe074} /* (8, 8, 6) {real, imag} */,
  {32'hbffeae86, 32'h403f7df0} /* (8, 8, 5) {real, imag} */,
  {32'hbf8aa352, 32'h3fd1019a} /* (8, 8, 4) {real, imag} */,
  {32'hc0054324, 32'hbf2a9ec0} /* (8, 8, 3) {real, imag} */,
  {32'hc0625d86, 32'h3fc13b4a} /* (8, 8, 2) {real, imag} */,
  {32'hc084397b, 32'h40065452} /* (8, 8, 1) {real, imag} */,
  {32'hbfc2681a, 32'h3f8d05ed} /* (8, 8, 0) {real, imag} */,
  {32'hbfbed5c6, 32'h401a0f72} /* (8, 7, 31) {real, imag} */,
  {32'hbea369f8, 32'h40880462} /* (8, 7, 30) {real, imag} */,
  {32'h3ee75ca0, 32'h4052aaf1} /* (8, 7, 29) {real, imag} */,
  {32'hbd20fa20, 32'h3fd01215} /* (8, 7, 28) {real, imag} */,
  {32'hbf05f7b0, 32'h3fc12591} /* (8, 7, 27) {real, imag} */,
  {32'hbfb1e9cb, 32'h3fb5dc84} /* (8, 7, 26) {real, imag} */,
  {32'h3ea8acf0, 32'h407acdd4} /* (8, 7, 25) {real, imag} */,
  {32'hbe8f666c, 32'h400fb37e} /* (8, 7, 24) {real, imag} */,
  {32'hc00987c4, 32'h3f960c82} /* (8, 7, 23) {real, imag} */,
  {32'hc043b0c3, 32'h40071a17} /* (8, 7, 22) {real, imag} */,
  {32'h3f5f81b2, 32'h3f993822} /* (8, 7, 21) {real, imag} */,
  {32'h3f703f54, 32'hbfdf3762} /* (8, 7, 20) {real, imag} */,
  {32'hbe189554, 32'hbf71f348} /* (8, 7, 19) {real, imag} */,
  {32'hbe8e41a4, 32'hc026ac5c} /* (8, 7, 18) {real, imag} */,
  {32'h3fa52e26, 32'hbf87db17} /* (8, 7, 17) {real, imag} */,
  {32'h3fe13c2f, 32'hc0237a5a} /* (8, 7, 16) {real, imag} */,
  {32'h3e877432, 32'hc02387a4} /* (8, 7, 15) {real, imag} */,
  {32'h403a94e4, 32'hbf8c9748} /* (8, 7, 14) {real, imag} */,
  {32'h4053a9c6, 32'hbf915e89} /* (8, 7, 13) {real, imag} */,
  {32'h403d51b5, 32'hbfc24f26} /* (8, 7, 12) {real, imag} */,
  {32'h4028d191, 32'hbebcecee} /* (8, 7, 11) {real, imag} */,
  {32'h3df390a0, 32'h3f140fca} /* (8, 7, 10) {real, imag} */,
  {32'hbd92ef80, 32'h3fa5e870} /* (8, 7, 9) {real, imag} */,
  {32'hbe4f3008, 32'h400c3b5b} /* (8, 7, 8) {real, imag} */,
  {32'hc02b6e83, 32'h3ff6d92c} /* (8, 7, 7) {real, imag} */,
  {32'hc06f2e54, 32'h4027707a} /* (8, 7, 6) {real, imag} */,
  {32'hc0177d4c, 32'h4083e535} /* (8, 7, 5) {real, imag} */,
  {32'hc0177bda, 32'h405950e2} /* (8, 7, 4) {real, imag} */,
  {32'hc01a86f3, 32'h3f968aa2} /* (8, 7, 3) {real, imag} */,
  {32'hc03194a2, 32'h3f9a75f2} /* (8, 7, 2) {real, imag} */,
  {32'hc01c78e8, 32'h4003ea64} /* (8, 7, 1) {real, imag} */,
  {32'hbf9c8944, 32'h3f862350} /* (8, 7, 0) {real, imag} */,
  {32'hbfaff50b, 32'h40175aa8} /* (8, 6, 31) {real, imag} */,
  {32'hbe7eb44c, 32'h403772eb} /* (8, 6, 30) {real, imag} */,
  {32'hc00deff0, 32'h3fddfe4b} /* (8, 6, 29) {real, imag} */,
  {32'hbfe8c92a, 32'h4003e238} /* (8, 6, 28) {real, imag} */,
  {32'hbf6a349e, 32'h4010a3f5} /* (8, 6, 27) {real, imag} */,
  {32'hbeb0bbe4, 32'h40476c22} /* (8, 6, 26) {real, imag} */,
  {32'h3e50c120, 32'h405fd8e5} /* (8, 6, 25) {real, imag} */,
  {32'hc002d2b0, 32'h3fff40f4} /* (8, 6, 24) {real, imag} */,
  {32'hc010fd56, 32'hbe816524} /* (8, 6, 23) {real, imag} */,
  {32'hc00f0234, 32'h3f836ca3} /* (8, 6, 22) {real, imag} */,
  {32'hbf2e0bce, 32'h400aac50} /* (8, 6, 21) {real, imag} */,
  {32'h3f5cc01f, 32'hc023c868} /* (8, 6, 20) {real, imag} */,
  {32'h3e34d124, 32'hbfbb37ff} /* (8, 6, 19) {real, imag} */,
  {32'h3fa89d0e, 32'hc0189f94} /* (8, 6, 18) {real, imag} */,
  {32'h3fbfe70a, 32'hc01a5ef3} /* (8, 6, 17) {real, imag} */,
  {32'h3f138bac, 32'hbfd475d4} /* (8, 6, 16) {real, imag} */,
  {32'h3f51b5db, 32'hbfa1b158} /* (8, 6, 15) {real, imag} */,
  {32'h40060b86, 32'hc00b3148} /* (8, 6, 14) {real, imag} */,
  {32'h3f6a4e68, 32'hc037203e} /* (8, 6, 13) {real, imag} */,
  {32'h3f15ef3d, 32'hbfe6daba} /* (8, 6, 12) {real, imag} */,
  {32'h3f7bcea4, 32'hbe8d2ee0} /* (8, 6, 11) {real, imag} */,
  {32'hc018696c, 32'h3f937aa8} /* (8, 6, 10) {real, imag} */,
  {32'hc03d135a, 32'h405630f0} /* (8, 6, 9) {real, imag} */,
  {32'hbfe1bfc4, 32'h40828042} /* (8, 6, 8) {real, imag} */,
  {32'hc02f3d4e, 32'h3fec862c} /* (8, 6, 7) {real, imag} */,
  {32'hc051ed30, 32'h3fb187bd} /* (8, 6, 6) {real, imag} */,
  {32'hbff7f187, 32'h3fcbf671} /* (8, 6, 5) {real, imag} */,
  {32'hbff27b9f, 32'h406cdaee} /* (8, 6, 4) {real, imag} */,
  {32'hbf9f2d34, 32'h403f1dbc} /* (8, 6, 3) {real, imag} */,
  {32'hbf80f6b0, 32'h3ff6c60f} /* (8, 6, 2) {real, imag} */,
  {32'hc045d915, 32'h401e8f2b} /* (8, 6, 1) {real, imag} */,
  {32'hbfe7b605, 32'h3f5cfca7} /* (8, 6, 0) {real, imag} */,
  {32'h3d0a11a0, 32'h3f0abe2c} /* (8, 5, 31) {real, imag} */,
  {32'hbf4c7f56, 32'h3fa500d8} /* (8, 5, 30) {real, imag} */,
  {32'hc01db64a, 32'h3fccc286} /* (8, 5, 29) {real, imag} */,
  {32'hc030f21e, 32'h4068c3b8} /* (8, 5, 28) {real, imag} */,
  {32'hbff0a988, 32'h40248105} /* (8, 5, 27) {real, imag} */,
  {32'hbfe325d2, 32'h401f3b2c} /* (8, 5, 26) {real, imag} */,
  {32'hbd1c81f0, 32'h404dc922} /* (8, 5, 25) {real, imag} */,
  {32'hbf9acb02, 32'h3f97ef26} /* (8, 5, 24) {real, imag} */,
  {32'hbf94653e, 32'h3efe27ae} /* (8, 5, 23) {real, imag} */,
  {32'hbfa19bca, 32'h3ff32dd0} /* (8, 5, 22) {real, imag} */,
  {32'hc04cd078, 32'h400360b8} /* (8, 5, 21) {real, imag} */,
  {32'hbfb30e06, 32'h3e5b6e98} /* (8, 5, 20) {real, imag} */,
  {32'h3f565680, 32'h3fa79ac4} /* (8, 5, 19) {real, imag} */,
  {32'h400ef0d6, 32'h3e902e36} /* (8, 5, 18) {real, imag} */,
  {32'hbe4745e8, 32'hbfc081be} /* (8, 5, 17) {real, imag} */,
  {32'h3efb8796, 32'hbf8b5d12} /* (8, 5, 16) {real, imag} */,
  {32'h402b174f, 32'hbfb46558} /* (8, 5, 15) {real, imag} */,
  {32'h40633654, 32'hc02f75e3} /* (8, 5, 14) {real, imag} */,
  {32'h3fb2615c, 32'hc00271ce} /* (8, 5, 13) {real, imag} */,
  {32'h3fb5eb26, 32'hbf26809c} /* (8, 5, 12) {real, imag} */,
  {32'h3f897058, 32'hbe146fb0} /* (8, 5, 11) {real, imag} */,
  {32'hbf8c8aa4, 32'h3f953e88} /* (8, 5, 10) {real, imag} */,
  {32'h3e1e4916, 32'h3ff3695a} /* (8, 5, 9) {real, imag} */,
  {32'h3fcf4e8c, 32'h3ebdc0bf} /* (8, 5, 8) {real, imag} */,
  {32'h3fa0b0af, 32'hbfc97426} /* (8, 5, 7) {real, imag} */,
  {32'h3e3b2940, 32'hbd2170f4} /* (8, 5, 6) {real, imag} */,
  {32'hbd6c1a20, 32'hbdd5afa0} /* (8, 5, 5) {real, imag} */,
  {32'hbf684f31, 32'h4018d4e8} /* (8, 5, 4) {real, imag} */,
  {32'hbffa1032, 32'h40176292} /* (8, 5, 3) {real, imag} */,
  {32'hbfd46578, 32'h40208856} /* (8, 5, 2) {real, imag} */,
  {32'hc02bdd69, 32'h402006ce} /* (8, 5, 1) {real, imag} */,
  {32'hbefe3a12, 32'h3db2eae0} /* (8, 5, 0) {real, imag} */,
  {32'h3eae0f00, 32'hbf526000} /* (8, 4, 31) {real, imag} */,
  {32'h3f8f41e0, 32'h3e4a8528} /* (8, 4, 30) {real, imag} */,
  {32'hbf4fdcd0, 32'h3df93cb0} /* (8, 4, 29) {real, imag} */,
  {32'hc0632608, 32'h3fd59451} /* (8, 4, 28) {real, imag} */,
  {32'hbf5205ea, 32'h3f894189} /* (8, 4, 27) {real, imag} */,
  {32'hbfe5f033, 32'h3ee1a866} /* (8, 4, 26) {real, imag} */,
  {32'hbfcce55c, 32'h3fcf07d1} /* (8, 4, 25) {real, imag} */,
  {32'hc0222063, 32'h3fcfeef3} /* (8, 4, 24) {real, imag} */,
  {32'hbf7671f1, 32'h3fa020df} /* (8, 4, 23) {real, imag} */,
  {32'hbff65d0e, 32'h3f8d3cd9} /* (8, 4, 22) {real, imag} */,
  {32'hc03aa674, 32'h3fbffc78} /* (8, 4, 21) {real, imag} */,
  {32'hc0519392, 32'h3f9f4242} /* (8, 4, 20) {real, imag} */,
  {32'hbf9cf1c6, 32'h400a9791} /* (8, 4, 19) {real, imag} */,
  {32'hbee49210, 32'h401351e2} /* (8, 4, 18) {real, imag} */,
  {32'hbf8c7203, 32'h404dad4c} /* (8, 4, 17) {real, imag} */,
  {32'hbf488cdd, 32'h403a69b2} /* (8, 4, 16) {real, imag} */,
  {32'h400700e2, 32'h3d0d1d00} /* (8, 4, 15) {real, imag} */,
  {32'h40846746, 32'hbf800cd3} /* (8, 4, 14) {real, imag} */,
  {32'h4017bb2c, 32'hbebec31c} /* (8, 4, 13) {real, imag} */,
  {32'h3fa3e270, 32'h3fa001d4} /* (8, 4, 12) {real, imag} */,
  {32'h3f29a758, 32'hbf6477af} /* (8, 4, 11) {real, imag} */,
  {32'h3e587bb8, 32'h3e563e78} /* (8, 4, 10) {real, imag} */,
  {32'h4005e1c9, 32'hbee56be4} /* (8, 4, 9) {real, imag} */,
  {32'h4058895b, 32'hc01dd169} /* (8, 4, 8) {real, imag} */,
  {32'h40262b84, 32'hc0200932} /* (8, 4, 7) {real, imag} */,
  {32'h3fcca50e, 32'hbebfc7cc} /* (8, 4, 6) {real, imag} */,
  {32'hbf1c86cf, 32'h3f201f34} /* (8, 4, 5) {real, imag} */,
  {32'hc004ecb0, 32'h3fb50104} /* (8, 4, 4) {real, imag} */,
  {32'hc03b9b54, 32'h404157fd} /* (8, 4, 3) {real, imag} */,
  {32'hc0431a20, 32'h40271f8c} /* (8, 4, 2) {real, imag} */,
  {32'hc04d0d32, 32'h400228f2} /* (8, 4, 1) {real, imag} */,
  {32'hbfdcbcc7, 32'h3ebee4ee} /* (8, 4, 0) {real, imag} */,
  {32'hbf816eac, 32'h3f3485a4} /* (8, 3, 31) {real, imag} */,
  {32'hbe448f4c, 32'h401cd738} /* (8, 3, 30) {real, imag} */,
  {32'hbdcc3d00, 32'h40261ec0} /* (8, 3, 29) {real, imag} */,
  {32'hc021aa7e, 32'h40697d90} /* (8, 3, 28) {real, imag} */,
  {32'hbf65f7dc, 32'h403239aa} /* (8, 3, 27) {real, imag} */,
  {32'hbfa3f9ec, 32'h3f91c07a} /* (8, 3, 26) {real, imag} */,
  {32'hbfdceb5c, 32'h3f01309e} /* (8, 3, 25) {real, imag} */,
  {32'hc07620a0, 32'h3fdfb38b} /* (8, 3, 24) {real, imag} */,
  {32'hbf094c81, 32'h40170c94} /* (8, 3, 23) {real, imag} */,
  {32'hc02e3220, 32'h3fc24ea5} /* (8, 3, 22) {real, imag} */,
  {32'hc0691798, 32'h402333c3} /* (8, 3, 21) {real, imag} */,
  {32'hc0481fdb, 32'h3fa2d9d6} /* (8, 3, 20) {real, imag} */,
  {32'hc00a9982, 32'h402801c4} /* (8, 3, 19) {real, imag} */,
  {32'hc0768ca2, 32'h40452ed4} /* (8, 3, 18) {real, imag} */,
  {32'hc01f30fc, 32'h403c983b} /* (8, 3, 17) {real, imag} */,
  {32'hbf2ceed6, 32'h40036265} /* (8, 3, 16) {real, imag} */,
  {32'h3fc79254, 32'hc00d6c13} /* (8, 3, 15) {real, imag} */,
  {32'h40413332, 32'hbff758bf} /* (8, 3, 14) {real, imag} */,
  {32'h401d10d6, 32'hc03b13a5} /* (8, 3, 13) {real, imag} */,
  {32'h40061982, 32'hbed9eb50} /* (8, 3, 12) {real, imag} */,
  {32'h3fbe0145, 32'hbeb40542} /* (8, 3, 11) {real, imag} */,
  {32'h3faa4921, 32'hbf843f64} /* (8, 3, 10) {real, imag} */,
  {32'h3fd66e41, 32'hbf416bc4} /* (8, 3, 9) {real, imag} */,
  {32'h401ad6cc, 32'hbfe42d44} /* (8, 3, 8) {real, imag} */,
  {32'h3ff3ff1b, 32'hc027514c} /* (8, 3, 7) {real, imag} */,
  {32'h3f24c7fa, 32'hbf57197f} /* (8, 3, 6) {real, imag} */,
  {32'h3e5631fa, 32'h3fde5e86} /* (8, 3, 5) {real, imag} */,
  {32'hbf934e2a, 32'h40039cda} /* (8, 3, 4) {real, imag} */,
  {32'hbfcdd4da, 32'h4065754a} /* (8, 3, 3) {real, imag} */,
  {32'hbff31b5e, 32'h403d4d01} /* (8, 3, 2) {real, imag} */,
  {32'hbfd148d5, 32'h40039fc1} /* (8, 3, 1) {real, imag} */,
  {32'hbfe7b66d, 32'h3eba50e4} /* (8, 3, 0) {real, imag} */,
  {32'hbec07f68, 32'h3e72fbf4} /* (8, 2, 31) {real, imag} */,
  {32'hbf6858a5, 32'h3feda0ce} /* (8, 2, 30) {real, imag} */,
  {32'hbd9a4248, 32'h400b249a} /* (8, 2, 29) {real, imag} */,
  {32'hc01ac10a, 32'h4069fe3b} /* (8, 2, 28) {real, imag} */,
  {32'hc01ed8d0, 32'h401e17a0} /* (8, 2, 27) {real, imag} */,
  {32'hc009ae5c, 32'h3f53e40e} /* (8, 2, 26) {real, imag} */,
  {32'hbf3991b9, 32'hbe54f2a2} /* (8, 2, 25) {real, imag} */,
  {32'hbf35348c, 32'hbdc86650} /* (8, 2, 24) {real, imag} */,
  {32'h3f57f39c, 32'h3fab3a95} /* (8, 2, 23) {real, imag} */,
  {32'hc0131bcb, 32'h3e2585fc} /* (8, 2, 22) {real, imag} */,
  {32'hc0670370, 32'h40478fad} /* (8, 2, 21) {real, imag} */,
  {32'hbf79f4a4, 32'h401b4cb6} /* (8, 2, 20) {real, imag} */,
  {32'hbfa7ac31, 32'h400c6ec0} /* (8, 2, 19) {real, imag} */,
  {32'hc04770cb, 32'h403dd3b4} /* (8, 2, 18) {real, imag} */,
  {32'hc05abda5, 32'h3fd25ac7} /* (8, 2, 17) {real, imag} */,
  {32'hbc27d600, 32'hbe4ff738} /* (8, 2, 16) {real, imag} */,
  {32'h3ff05c26, 32'hc086faa7} /* (8, 2, 15) {real, imag} */,
  {32'h3f63e449, 32'hc03e453e} /* (8, 2, 14) {real, imag} */,
  {32'h3f7c3904, 32'hc08efd4f} /* (8, 2, 13) {real, imag} */,
  {32'h407591a6, 32'hc075c2a9} /* (8, 2, 12) {real, imag} */,
  {32'h40584641, 32'hc045e47a} /* (8, 2, 11) {real, imag} */,
  {32'h3fe60f87, 32'hbff1d5ef} /* (8, 2, 10) {real, imag} */,
  {32'hbf020194, 32'hbfc64d94} /* (8, 2, 9) {real, imag} */,
  {32'h3f2a70a1, 32'hc0028d2e} /* (8, 2, 8) {real, imag} */,
  {32'h4002b65b, 32'hbff3fc4c} /* (8, 2, 7) {real, imag} */,
  {32'h3ff408c8, 32'hbffefe3a} /* (8, 2, 6) {real, imag} */,
  {32'h404b7fcc, 32'h3e95d24f} /* (8, 2, 5) {real, imag} */,
  {32'h3f5b8353, 32'h406308ab} /* (8, 2, 4) {real, imag} */,
  {32'hc0011e86, 32'h40608bb9} /* (8, 2, 3) {real, imag} */,
  {32'hbf0b2d24, 32'h40435087} /* (8, 2, 2) {real, imag} */,
  {32'h3ff061c8, 32'h407a799e} /* (8, 2, 1) {real, imag} */,
  {32'hbdbd6834, 32'h4004aaca} /* (8, 2, 0) {real, imag} */,
  {32'h3fca2a1c, 32'h3f5db2e5} /* (8, 1, 31) {real, imag} */,
  {32'hbf12c9fc, 32'h40194de2} /* (8, 1, 30) {real, imag} */,
  {32'hc016bccb, 32'h3fb09c1f} /* (8, 1, 29) {real, imag} */,
  {32'hc095f85c, 32'h400dbaa2} /* (8, 1, 28) {real, imag} */,
  {32'hc082c7f6, 32'h4014fda8} /* (8, 1, 27) {real, imag} */,
  {32'hbfa68913, 32'h3fee4244} /* (8, 1, 26) {real, imag} */,
  {32'hbe9097d8, 32'h3fc52690} /* (8, 1, 25) {real, imag} */,
  {32'hbe5925a8, 32'h3f1d72de} /* (8, 1, 24) {real, imag} */,
  {32'h3f91ed2e, 32'h401d676a} /* (8, 1, 23) {real, imag} */,
  {32'hbf94e9a7, 32'h4029a8c4} /* (8, 1, 22) {real, imag} */,
  {32'hbfd0e044, 32'h40407348} /* (8, 1, 21) {real, imag} */,
  {32'h3e4587ec, 32'h40370448} /* (8, 1, 20) {real, imag} */,
  {32'hbf18246e, 32'h40477676} /* (8, 1, 19) {real, imag} */,
  {32'hbf88d695, 32'h4082e22e} /* (8, 1, 18) {real, imag} */,
  {32'hbfd14bc4, 32'h3fb97bb8} /* (8, 1, 17) {real, imag} */,
  {32'h3faf407e, 32'h3e6147c0} /* (8, 1, 16) {real, imag} */,
  {32'h40024234, 32'hc027f180} /* (8, 1, 15) {real, imag} */,
  {32'h3e0f1bd0, 32'hc0635072} /* (8, 1, 14) {real, imag} */,
  {32'h3f9c2e3e, 32'hbfa86206} /* (8, 1, 13) {real, imag} */,
  {32'h40084a76, 32'hbfdd2060} /* (8, 1, 12) {real, imag} */,
  {32'h40714cde, 32'hc02acbfd} /* (8, 1, 11) {real, imag} */,
  {32'h4045adfb, 32'hc0427c67} /* (8, 1, 10) {real, imag} */,
  {32'h3f08aab1, 32'hc009e869} /* (8, 1, 9) {real, imag} */,
  {32'h3f9ff604, 32'hc0107666} /* (8, 1, 8) {real, imag} */,
  {32'h40109026, 32'hbe953226} /* (8, 1, 7) {real, imag} */,
  {32'h4032f410, 32'h3e14cf18} /* (8, 1, 6) {real, imag} */,
  {32'hbe1668b6, 32'h3e9b3fec} /* (8, 1, 5) {real, imag} */,
  {32'hbfed39f6, 32'h40430626} /* (8, 1, 4) {real, imag} */,
  {32'hc00b5bf7, 32'h3ff2e35c} /* (8, 1, 3) {real, imag} */,
  {32'h3f26437c, 32'h3ffb601d} /* (8, 1, 2) {real, imag} */,
  {32'h401eaa64, 32'h3fd4be5c} /* (8, 1, 1) {real, imag} */,
  {32'h3fb71b68, 32'h3f880617} /* (8, 1, 0) {real, imag} */,
  {32'h3d8f6c84, 32'h3e98a277} /* (8, 0, 31) {real, imag} */,
  {32'hbf8b63d6, 32'h3e0c79a6} /* (8, 0, 30) {real, imag} */,
  {32'hc02514bf, 32'hbe209f2e} /* (8, 0, 29) {real, imag} */,
  {32'hc0690db2, 32'h3f4015c0} /* (8, 0, 28) {real, imag} */,
  {32'hc072fd0c, 32'h3ff106ae} /* (8, 0, 27) {real, imag} */,
  {32'hbf74348e, 32'h3fd4f560} /* (8, 0, 26) {real, imag} */,
  {32'hbf1bf4e5, 32'h3f224366} /* (8, 0, 25) {real, imag} */,
  {32'hbe7c37a0, 32'hbf5b9d5c} /* (8, 0, 24) {real, imag} */,
  {32'h3dbe8808, 32'h3ff7aa26} /* (8, 0, 23) {real, imag} */,
  {32'hbf29548a, 32'h403f9f0b} /* (8, 0, 22) {real, imag} */,
  {32'hbf1d04ed, 32'h3f648ce6} /* (8, 0, 21) {real, imag} */,
  {32'h3d7b6b20, 32'h3ee14873} /* (8, 0, 20) {real, imag} */,
  {32'hbda93d40, 32'h3fdb2e6a} /* (8, 0, 19) {real, imag} */,
  {32'hbead3ab0, 32'h3ff0c93e} /* (8, 0, 18) {real, imag} */,
  {32'hbed222d4, 32'h3f3d953e} /* (8, 0, 17) {real, imag} */,
  {32'h3f6539bc, 32'h3f349962} /* (8, 0, 16) {real, imag} */,
  {32'h3f4f84d8, 32'hbf359b88} /* (8, 0, 15) {real, imag} */,
  {32'h3f7225e6, 32'hc010dbe6} /* (8, 0, 14) {real, imag} */,
  {32'h400ce0a2, 32'hbf40171b} /* (8, 0, 13) {real, imag} */,
  {32'h3f2b14ee, 32'hbfab367a} /* (8, 0, 12) {real, imag} */,
  {32'h3fa75646, 32'hbff2a6ce} /* (8, 0, 11) {real, imag} */,
  {32'h3f64ec04, 32'hbfaa04c6} /* (8, 0, 10) {real, imag} */,
  {32'h3f39ad56, 32'h3f04b7aa} /* (8, 0, 9) {real, imag} */,
  {32'h3fcabc94, 32'h3dd4f8f8} /* (8, 0, 8) {real, imag} */,
  {32'h4011c5bb, 32'h3f39e498} /* (8, 0, 7) {real, imag} */,
  {32'h3f9c02ea, 32'h3fd5c74a} /* (8, 0, 6) {real, imag} */,
  {32'hbfb7f67e, 32'h3f0dc23c} /* (8, 0, 5) {real, imag} */,
  {32'hbffc3fba, 32'h3f85b6d5} /* (8, 0, 4) {real, imag} */,
  {32'hbf9ae831, 32'h3f31b52e} /* (8, 0, 3) {real, imag} */,
  {32'h3f5639ce, 32'h40013f58} /* (8, 0, 2) {real, imag} */,
  {32'h3fa4e7f8, 32'h3f464a7e} /* (8, 0, 1) {real, imag} */,
  {32'hbb4a6b00, 32'hbe8a287c} /* (8, 0, 0) {real, imag} */,
  {32'hbf8f6ba8, 32'h3e8e2108} /* (7, 31, 31) {real, imag} */,
  {32'hbf839c43, 32'h3f5197d2} /* (7, 31, 30) {real, imag} */,
  {32'hbfe2b12b, 32'h3d1e6080} /* (7, 31, 29) {real, imag} */,
  {32'hbf029e6e, 32'h3e7fa802} /* (7, 31, 28) {real, imag} */,
  {32'hbd206838, 32'h3f886002} /* (7, 31, 27) {real, imag} */,
  {32'hbfa4d401, 32'h3f5885d8} /* (7, 31, 26) {real, imag} */,
  {32'h3a179c00, 32'hbf0e26d0} /* (7, 31, 25) {real, imag} */,
  {32'h3f7b91f8, 32'hbfe109c0} /* (7, 31, 24) {real, imag} */,
  {32'h3fb5811e, 32'hbf8b1ce0} /* (7, 31, 23) {real, imag} */,
  {32'h3f991b21, 32'hbea66a03} /* (7, 31, 22) {real, imag} */,
  {32'h3f96b794, 32'hbf153dea} /* (7, 31, 21) {real, imag} */,
  {32'h3fa30cc1, 32'hbfae2479} /* (7, 31, 20) {real, imag} */,
  {32'hbd8be810, 32'hbf760419} /* (7, 31, 19) {real, imag} */,
  {32'h3dbb40a4, 32'hbf3e043e} /* (7, 31, 18) {real, imag} */,
  {32'h3ef74bc8, 32'h3f3fe5fa} /* (7, 31, 17) {real, imag} */,
  {32'h3f40902e, 32'h3e13c1be} /* (7, 31, 16) {real, imag} */,
  {32'h3e2f5f03, 32'h3f45cf06} /* (7, 31, 15) {real, imag} */,
  {32'hbfc07db2, 32'h3e32990f} /* (7, 31, 14) {real, imag} */,
  {32'hbfff7603, 32'h3fafb13a} /* (7, 31, 13) {real, imag} */,
  {32'h3ed0239c, 32'h40147afe} /* (7, 31, 12) {real, imag} */,
  {32'h3fefa61a, 32'h3fd65368} /* (7, 31, 11) {real, imag} */,
  {32'hbe0d0bc7, 32'h4001268e} /* (7, 31, 10) {real, imag} */,
  {32'h3e1d0d3c, 32'hbce0da90} /* (7, 31, 9) {real, imag} */,
  {32'h3f6398a5, 32'hbf62cd50} /* (7, 31, 8) {real, imag} */,
  {32'h400f4538, 32'hbe95e618} /* (7, 31, 7) {real, imag} */,
  {32'h3d897a70, 32'h3f00549a} /* (7, 31, 6) {real, imag} */,
  {32'hbe54c9c8, 32'h403022d1} /* (7, 31, 5) {real, imag} */,
  {32'hbecd2d9f, 32'h3fd424ee} /* (7, 31, 4) {real, imag} */,
  {32'hbfade374, 32'hbf0d0bd7} /* (7, 31, 3) {real, imag} */,
  {32'hbe79bc77, 32'hbeafa922} /* (7, 31, 2) {real, imag} */,
  {32'h3f464511, 32'hbf9a84c6} /* (7, 31, 1) {real, imag} */,
  {32'hbf84740a, 32'hbf32b4c0} /* (7, 31, 0) {real, imag} */,
  {32'hbfc86320, 32'hbf8914d7} /* (7, 30, 31) {real, imag} */,
  {32'hbfd0da86, 32'hbf9b3c08} /* (7, 30, 30) {real, imag} */,
  {32'hbfac0794, 32'hbf934f94} /* (7, 30, 29) {real, imag} */,
  {32'h3f81ff44, 32'hbeefa6ed} /* (7, 30, 28) {real, imag} */,
  {32'h3face322, 32'h3f9fc338} /* (7, 30, 27) {real, imag} */,
  {32'hbf3d221e, 32'hbe9ded64} /* (7, 30, 26) {real, imag} */,
  {32'h3eb89214, 32'hbf42b2e0} /* (7, 30, 25) {real, imag} */,
  {32'h3e748ed8, 32'hc029f24e} /* (7, 30, 24) {real, imag} */,
  {32'hbce451d0, 32'hbf4587d4} /* (7, 30, 23) {real, imag} */,
  {32'h3d8ebe02, 32'h3fba42cc} /* (7, 30, 22) {real, imag} */,
  {32'hbf0caa55, 32'h3d18d308} /* (7, 30, 21) {real, imag} */,
  {32'hbd295f30, 32'hbf421f60} /* (7, 30, 20) {real, imag} */,
  {32'hc018912a, 32'hbe7f5d94} /* (7, 30, 19) {real, imag} */,
  {32'hc0097128, 32'hbf32e9d9} /* (7, 30, 18) {real, imag} */,
  {32'h3fb186bd, 32'h3dd6dd32} /* (7, 30, 17) {real, imag} */,
  {32'h3f6349ba, 32'hbf9a5b7d} /* (7, 30, 16) {real, imag} */,
  {32'hbfd2080b, 32'hbe9a8c0c} /* (7, 30, 15) {real, imag} */,
  {32'hbff03075, 32'h3f6315c4} /* (7, 30, 14) {real, imag} */,
  {32'hbfcd0672, 32'h401d3506} /* (7, 30, 13) {real, imag} */,
  {32'hbe5606ac, 32'h40771ee5} /* (7, 30, 12) {real, imag} */,
  {32'h3facd87e, 32'h3f4a06fc} /* (7, 30, 11) {real, imag} */,
  {32'h3f14cf43, 32'h3e2a4b58} /* (7, 30, 10) {real, imag} */,
  {32'h3ef7e768, 32'hbfac9967} /* (7, 30, 9) {real, imag} */,
  {32'h3eda22ca, 32'hbfec78ea} /* (7, 30, 8) {real, imag} */,
  {32'h402a4eea, 32'hbe4acfc0} /* (7, 30, 7) {real, imag} */,
  {32'hbf90025d, 32'h3fb1f7d0} /* (7, 30, 6) {real, imag} */,
  {32'hc03cffe2, 32'h402e11b7} /* (7, 30, 5) {real, imag} */,
  {32'hbffa6b44, 32'h40122946} /* (7, 30, 4) {real, imag} */,
  {32'hbfa8c09c, 32'h3f274deb} /* (7, 30, 3) {real, imag} */,
  {32'h3d80ba10, 32'hbf393a7a} /* (7, 30, 2) {real, imag} */,
  {32'h3e03663c, 32'hc05c00c2} /* (7, 30, 1) {real, imag} */,
  {32'hbf86022d, 32'hc00a5e52} /* (7, 30, 0) {real, imag} */,
  {32'hbf3d74ad, 32'hbf66aaac} /* (7, 29, 31) {real, imag} */,
  {32'hbf38b68a, 32'hbf495aa8} /* (7, 29, 30) {real, imag} */,
  {32'hbf9282d3, 32'hbe5a53a8} /* (7, 29, 29) {real, imag} */,
  {32'h3fe03a80, 32'hc00cf7fe} /* (7, 29, 28) {real, imag} */,
  {32'h406c079e, 32'hbfbb034f} /* (7, 29, 27) {real, imag} */,
  {32'h3fa5bee0, 32'h3d9552a8} /* (7, 29, 26) {real, imag} */,
  {32'h3f22aec6, 32'hbe650fc8} /* (7, 29, 25) {real, imag} */,
  {32'h3b86d500, 32'hbfeb9a32} /* (7, 29, 24) {real, imag} */,
  {32'hbfb53e62, 32'hbee230b7} /* (7, 29, 23) {real, imag} */,
  {32'hbe288ea8, 32'h3f54355c} /* (7, 29, 22) {real, imag} */,
  {32'hbf8c519f, 32'hbfe5e506} /* (7, 29, 21) {real, imag} */,
  {32'hbff4fe24, 32'hbf8fe0ae} /* (7, 29, 20) {real, imag} */,
  {32'hc078936d, 32'h3fcba601} /* (7, 29, 19) {real, imag} */,
  {32'hc0550d76, 32'h3d3153d0} /* (7, 29, 18) {real, imag} */,
  {32'h3f0ff873, 32'h3f2853a7} /* (7, 29, 17) {real, imag} */,
  {32'h3f3de902, 32'h3dca16c0} /* (7, 29, 16) {real, imag} */,
  {32'hbfbe4430, 32'h3d717d10} /* (7, 29, 15) {real, imag} */,
  {32'hbd974360, 32'h3e00b920} /* (7, 29, 14) {real, imag} */,
  {32'h3f9f1336, 32'h3e28dd58} /* (7, 29, 13) {real, imag} */,
  {32'hbf1375ae, 32'h3ffe276e} /* (7, 29, 12) {real, imag} */,
  {32'hbf41c8ca, 32'hbefc2a7a} /* (7, 29, 11) {real, imag} */,
  {32'hbc40b880, 32'hc0033830} /* (7, 29, 10) {real, imag} */,
  {32'hbecdd678, 32'hbfa05eba} /* (7, 29, 9) {real, imag} */,
  {32'hbf4bff80, 32'hbffda430} /* (7, 29, 8) {real, imag} */,
  {32'hbeafd484, 32'hbf6ff917} /* (7, 29, 7) {real, imag} */,
  {32'hc032de7c, 32'h3f1addbc} /* (7, 29, 6) {real, imag} */,
  {32'hc0821e54, 32'h3f598410} /* (7, 29, 5) {real, imag} */,
  {32'hbf83e00c, 32'h3ede1872} /* (7, 29, 4) {real, imag} */,
  {32'h3f1f618c, 32'h401048ac} /* (7, 29, 3) {real, imag} */,
  {32'h3fa45796, 32'h40407793} /* (7, 29, 2) {real, imag} */,
  {32'h3ed8e06e, 32'hbf1a445d} /* (7, 29, 1) {real, imag} */,
  {32'hbfde07a0, 32'hbfde0056} /* (7, 29, 0) {real, imag} */,
  {32'h3e5a24e6, 32'h3f7c42f0} /* (7, 28, 31) {real, imag} */,
  {32'hbf9551e3, 32'h40069222} /* (7, 28, 30) {real, imag} */,
  {32'hc0629421, 32'h3f4ea468} /* (7, 28, 29) {real, imag} */,
  {32'h3ef0c24b, 32'hbfadb1b1} /* (7, 28, 28) {real, imag} */,
  {32'h4065801f, 32'hbfdf23e4} /* (7, 28, 27) {real, imag} */,
  {32'h3d945982, 32'h3fc45960} /* (7, 28, 26) {real, imag} */,
  {32'hbf2ae3da, 32'hbdf81130} /* (7, 28, 25) {real, imag} */,
  {32'h3f71bbb0, 32'hbf1712d5} /* (7, 28, 24) {real, imag} */,
  {32'h3f82d485, 32'hbf135252} /* (7, 28, 23) {real, imag} */,
  {32'h400b0378, 32'hc0482ab5} /* (7, 28, 22) {real, imag} */,
  {32'h3ff201d8, 32'hc006fd4a} /* (7, 28, 21) {real, imag} */,
  {32'h3f819a94, 32'hbfbefd65} /* (7, 28, 20) {real, imag} */,
  {32'hbfbbcf98, 32'h3ec17c40} /* (7, 28, 19) {real, imag} */,
  {32'hc0047c7e, 32'h3e359c28} /* (7, 28, 18) {real, imag} */,
  {32'hbf6cce08, 32'h3f931f60} /* (7, 28, 17) {real, imag} */,
  {32'hbf9003a9, 32'hbf7ae97c} /* (7, 28, 16) {real, imag} */,
  {32'hbf7135a0, 32'hbf719681} /* (7, 28, 15) {real, imag} */,
  {32'hbf0b083c, 32'hbd950da0} /* (7, 28, 14) {real, imag} */,
  {32'h3f9eb4fe, 32'hbf9020b9} /* (7, 28, 13) {real, imag} */,
  {32'hbf6d2f02, 32'h3df066e8} /* (7, 28, 12) {real, imag} */,
  {32'hbf779898, 32'hbf51b8c3} /* (7, 28, 11) {real, imag} */,
  {32'h4005f14a, 32'hc03df1eb} /* (7, 28, 10) {real, imag} */,
  {32'h40532fd2, 32'hc02a5d27} /* (7, 28, 9) {real, imag} */,
  {32'h3e850d13, 32'hbfab7aac} /* (7, 28, 8) {real, imag} */,
  {32'hbf777b89, 32'hbf97a525} /* (7, 28, 7) {real, imag} */,
  {32'hc0012220, 32'hbf3faf16} /* (7, 28, 6) {real, imag} */,
  {32'h3e975f24, 32'hbf53cfa6} /* (7, 28, 5) {real, imag} */,
  {32'h3fac2dd3, 32'hbfdf7c02} /* (7, 28, 4) {real, imag} */,
  {32'h3f605b49, 32'hbfcaa59b} /* (7, 28, 3) {real, imag} */,
  {32'h3f134f17, 32'h3f88d41e} /* (7, 28, 2) {real, imag} */,
  {32'h3f5aa6cc, 32'h3f9bb667} /* (7, 28, 1) {real, imag} */,
  {32'hbe977dc4, 32'h3f63fd4e} /* (7, 28, 0) {real, imag} */,
  {32'hbfeb98bc, 32'h3ef5f246} /* (7, 27, 31) {real, imag} */,
  {32'hbfdb3f62, 32'h3f8f481b} /* (7, 27, 30) {real, imag} */,
  {32'hbde312b8, 32'h3e98bc14} /* (7, 27, 29) {real, imag} */,
  {32'h3f9086b8, 32'h3fbb3382} /* (7, 27, 28) {real, imag} */,
  {32'h3fb0428b, 32'hbd463ea0} /* (7, 27, 27) {real, imag} */,
  {32'hbfa814a6, 32'h3e38c514} /* (7, 27, 26) {real, imag} */,
  {32'hbf8cebf0, 32'hbbfa33c0} /* (7, 27, 25) {real, imag} */,
  {32'h3f0d8315, 32'hbfa22daf} /* (7, 27, 24) {real, imag} */,
  {32'h3f149380, 32'hbf27e572} /* (7, 27, 23) {real, imag} */,
  {32'h4007fe44, 32'hc08876a9} /* (7, 27, 22) {real, imag} */,
  {32'h3ff7925b, 32'hbfe4385b} /* (7, 27, 21) {real, imag} */,
  {32'h3f42475a, 32'h3fb4e3b2} /* (7, 27, 20) {real, imag} */,
  {32'h3ebf1698, 32'h3fba7a60} /* (7, 27, 19) {real, imag} */,
  {32'h3f1652e0, 32'h3de47da8} /* (7, 27, 18) {real, imag} */,
  {32'h3e644b38, 32'hbde233d0} /* (7, 27, 17) {real, imag} */,
  {32'hbf453acc, 32'hbe851210} /* (7, 27, 16) {real, imag} */,
  {32'h3f2d5300, 32'hc0017102} /* (7, 27, 15) {real, imag} */,
  {32'h400a425a, 32'h3e0a6e70} /* (7, 27, 14) {real, imag} */,
  {32'h3fa55b4f, 32'h3fb8e2a6} /* (7, 27, 13) {real, imag} */,
  {32'hbf5c92ca, 32'hbc8fede0} /* (7, 27, 12) {real, imag} */,
  {32'hbfd939b2, 32'h3df808b0} /* (7, 27, 11) {real, imag} */,
  {32'h3ee5eed0, 32'hc000ffeb} /* (7, 27, 10) {real, imag} */,
  {32'h40225cb4, 32'hc01b1a3a} /* (7, 27, 9) {real, imag} */,
  {32'h3f55b975, 32'hbfe01d07} /* (7, 27, 8) {real, imag} */,
  {32'h3fa60c43, 32'hc0230300} /* (7, 27, 7) {real, imag} */,
  {32'h3f7c45d5, 32'hc02f001a} /* (7, 27, 6) {real, imag} */,
  {32'h3fbe5702, 32'hc03f9f3b} /* (7, 27, 5) {real, imag} */,
  {32'h3e03a588, 32'hbfe63392} /* (7, 27, 4) {real, imag} */,
  {32'h3eb1869a, 32'hbf088731} /* (7, 27, 3) {real, imag} */,
  {32'h4035152a, 32'hbe8d9931} /* (7, 27, 2) {real, imag} */,
  {32'h3f9706db, 32'hbf1c29b5} /* (7, 27, 1) {real, imag} */,
  {32'hbf87e43b, 32'h3ebd82b8} /* (7, 27, 0) {real, imag} */,
  {32'hbf8271a4, 32'h3f96b2bb} /* (7, 26, 31) {real, imag} */,
  {32'hbf5679a6, 32'h3f3730cd} /* (7, 26, 30) {real, imag} */,
  {32'hbe1d76f4, 32'hbe901a9e} /* (7, 26, 29) {real, imag} */,
  {32'h3f411830, 32'h3f53308c} /* (7, 26, 28) {real, imag} */,
  {32'hbd178af0, 32'hbee1e65c} /* (7, 26, 27) {real, imag} */,
  {32'hbfc45029, 32'h3e3020cc} /* (7, 26, 26) {real, imag} */,
  {32'hbee54b74, 32'h3f959280} /* (7, 26, 25) {real, imag} */,
  {32'h3f179d58, 32'hbfe104bc} /* (7, 26, 24) {real, imag} */,
  {32'hbf89b26c, 32'hbe966fbf} /* (7, 26, 23) {real, imag} */,
  {32'hbe8a5ef3, 32'hbf9d5690} /* (7, 26, 22) {real, imag} */,
  {32'hbea0b800, 32'hbf5b647e} /* (7, 26, 21) {real, imag} */,
  {32'hc00db592, 32'h3f9b5fda} /* (7, 26, 20) {real, imag} */,
  {32'hbf12a808, 32'h3f0f6d68} /* (7, 26, 19) {real, imag} */,
  {32'hbfa24e13, 32'hbebb5960} /* (7, 26, 18) {real, imag} */,
  {32'hbf87a9c6, 32'h3fb58c38} /* (7, 26, 17) {real, imag} */,
  {32'hbf5fbcf2, 32'h3fea6cfa} /* (7, 26, 16) {real, imag} */,
  {32'h3fccb344, 32'hc02abc9c} /* (7, 26, 15) {real, imag} */,
  {32'h404628e2, 32'hbfbaea29} /* (7, 26, 14) {real, imag} */,
  {32'h3eed8266, 32'h3fd0d444} /* (7, 26, 13) {real, imag} */,
  {32'hbf5e8892, 32'h3ed1edf2} /* (7, 26, 12) {real, imag} */,
  {32'hbf710c32, 32'hbeac8464} /* (7, 26, 11) {real, imag} */,
  {32'hbf3230d7, 32'hc02f9670} /* (7, 26, 10) {real, imag} */,
  {32'h3f64287c, 32'hbfff974e} /* (7, 26, 9) {real, imag} */,
  {32'h3faa3b2c, 32'hbf94966c} /* (7, 26, 8) {real, imag} */,
  {32'h4024933a, 32'hbfd45c72} /* (7, 26, 7) {real, imag} */,
  {32'h4048e5f0, 32'hc003df4e} /* (7, 26, 6) {real, imag} */,
  {32'h3f96a463, 32'hc0245661} /* (7, 26, 5) {real, imag} */,
  {32'hbfd135e7, 32'hbf9cc0a0} /* (7, 26, 4) {real, imag} */,
  {32'hbf94779e, 32'hbf0ef7d1} /* (7, 26, 3) {real, imag} */,
  {32'h3feac6ef, 32'hbf540d4c} /* (7, 26, 2) {real, imag} */,
  {32'h3f433e32, 32'hbfb17250} /* (7, 26, 1) {real, imag} */,
  {32'hbf8ea2ac, 32'hbdddff34} /* (7, 26, 0) {real, imag} */,
  {32'h3eae0817, 32'h3f673c9c} /* (7, 25, 31) {real, imag} */,
  {32'hbf6559c6, 32'h3fd3a1de} /* (7, 25, 30) {real, imag} */,
  {32'hbf6f8814, 32'h3fb9f079} /* (7, 25, 29) {real, imag} */,
  {32'h3ea5bf12, 32'hbf150aa0} /* (7, 25, 28) {real, imag} */,
  {32'hbf5c4538, 32'hbf24d1cb} /* (7, 25, 27) {real, imag} */,
  {32'hc02806ae, 32'hbf6be99a} /* (7, 25, 26) {real, imag} */,
  {32'hbfd4d6e4, 32'h3f90a8a2} /* (7, 25, 25) {real, imag} */,
  {32'h3f248f71, 32'hbf1d6cec} /* (7, 25, 24) {real, imag} */,
  {32'h3c22d040, 32'hbfda53ca} /* (7, 25, 23) {real, imag} */,
  {32'h3e2df1d8, 32'hbf965320} /* (7, 25, 22) {real, imag} */,
  {32'hc0083f15, 32'hbfb56e96} /* (7, 25, 21) {real, imag} */,
  {32'hbee5e020, 32'hbfb87af1} /* (7, 25, 20) {real, imag} */,
  {32'h401196df, 32'hbe5f4d4c} /* (7, 25, 19) {real, imag} */,
  {32'hbe132932, 32'hbe496fb8} /* (7, 25, 18) {real, imag} */,
  {32'h3fb1d3a8, 32'h3f7d2f3a} /* (7, 25, 17) {real, imag} */,
  {32'h3fadf4a0, 32'h4036ccab} /* (7, 25, 16) {real, imag} */,
  {32'h3ea31978, 32'hbdc0448c} /* (7, 25, 15) {real, imag} */,
  {32'h3dde6c78, 32'hc005c2b2} /* (7, 25, 14) {real, imag} */,
  {32'hbf3b9950, 32'hbf75dd89} /* (7, 25, 13) {real, imag} */,
  {32'hbf550070, 32'h3f76c0e6} /* (7, 25, 12) {real, imag} */,
  {32'hbf5d5dba, 32'hbf671d05} /* (7, 25, 11) {real, imag} */,
  {32'hbf580836, 32'hc031d176} /* (7, 25, 10) {real, imag} */,
  {32'hbe2b0f78, 32'hbefc55ca} /* (7, 25, 9) {real, imag} */,
  {32'hbfd2d146, 32'h3f40bac4} /* (7, 25, 8) {real, imag} */,
  {32'hbebee08a, 32'h3e85fef7} /* (7, 25, 7) {real, imag} */,
  {32'h4046216e, 32'hc0022b38} /* (7, 25, 6) {real, imag} */,
  {32'h400e8301, 32'hc02f77cb} /* (7, 25, 5) {real, imag} */,
  {32'hbf9bff70, 32'hbf24b117} /* (7, 25, 4) {real, imag} */,
  {32'hbf8c2c25, 32'hbe68993a} /* (7, 25, 3) {real, imag} */,
  {32'hbf3d3af6, 32'hbfc26885} /* (7, 25, 2) {real, imag} */,
  {32'h3f72d158, 32'hbfb97679} /* (7, 25, 1) {real, imag} */,
  {32'h3fb18062, 32'h3f3eecf1} /* (7, 25, 0) {real, imag} */,
  {32'h3e32f0f1, 32'h3ea2eb0c} /* (7, 24, 31) {real, imag} */,
  {32'hbe830478, 32'hbe92ae9b} /* (7, 24, 30) {real, imag} */,
  {32'hbfd5426b, 32'h3e2d43c0} /* (7, 24, 29) {real, imag} */,
  {32'hbfb1b37f, 32'hc014ead8} /* (7, 24, 28) {real, imag} */,
  {32'hbfa7de1c, 32'hbf984618} /* (7, 24, 27) {real, imag} */,
  {32'hbf747451, 32'h3ec0989a} /* (7, 24, 26) {real, imag} */,
  {32'hbf485845, 32'h3e5a0176} /* (7, 24, 25) {real, imag} */,
  {32'h3f95ef69, 32'h3f135375} /* (7, 24, 24) {real, imag} */,
  {32'h3fb96a6a, 32'hbf2d6d62} /* (7, 24, 23) {real, imag} */,
  {32'h3dea4e10, 32'hbf80e666} /* (7, 24, 22) {real, imag} */,
  {32'hbedff3c9, 32'hbefc782a} /* (7, 24, 21) {real, imag} */,
  {32'h40162fbe, 32'h3f5479ff} /* (7, 24, 20) {real, imag} */,
  {32'h3fef54e3, 32'h3ff741b1} /* (7, 24, 19) {real, imag} */,
  {32'h3fb64789, 32'h3f8486a0} /* (7, 24, 18) {real, imag} */,
  {32'h4065eb98, 32'h3f826482} /* (7, 24, 17) {real, imag} */,
  {32'h3fb5d904, 32'h3fb66eee} /* (7, 24, 16) {real, imag} */,
  {32'hbfadf8ec, 32'h3f0c40f0} /* (7, 24, 15) {real, imag} */,
  {32'hbf938944, 32'hbf5dad46} /* (7, 24, 14) {real, imag} */,
  {32'hbf3095f0, 32'hbfa3a8c3} /* (7, 24, 13) {real, imag} */,
  {32'hc0863dbc, 32'hbf4e183d} /* (7, 24, 12) {real, imag} */,
  {32'hc02edfea, 32'hbf19f6b7} /* (7, 24, 11) {real, imag} */,
  {32'h3f96d64a, 32'hbf396b44} /* (7, 24, 10) {real, imag} */,
  {32'h3f7f82db, 32'h3fbe6ba4} /* (7, 24, 9) {real, imag} */,
  {32'hbf3eea9d, 32'hbda885a0} /* (7, 24, 8) {real, imag} */,
  {32'hbf2d4110, 32'hbfd533e6} /* (7, 24, 7) {real, imag} */,
  {32'h3ff1d04a, 32'hc0284914} /* (7, 24, 6) {real, imag} */,
  {32'h3fdb9ac0, 32'hbfe70aa0} /* (7, 24, 5) {real, imag} */,
  {32'h3f1dd20e, 32'hbf19abce} /* (7, 24, 4) {real, imag} */,
  {32'hbdb45430, 32'hbf949132} /* (7, 24, 3) {real, imag} */,
  {32'hbf46711f, 32'hbfe215c4} /* (7, 24, 2) {real, imag} */,
  {32'h402decef, 32'hbf6c09c6} /* (7, 24, 1) {real, imag} */,
  {32'h3fd59f2e, 32'h3e943bde} /* (7, 24, 0) {real, imag} */,
  {32'hbf78a0db, 32'hbee09a7e} /* (7, 23, 31) {real, imag} */,
  {32'hbf173140, 32'hbeed7677} /* (7, 23, 30) {real, imag} */,
  {32'h3efb5014, 32'hbfb19657} /* (7, 23, 29) {real, imag} */,
  {32'hbe057e40, 32'hc00eae75} /* (7, 23, 28) {real, imag} */,
  {32'h3d6c3dc8, 32'hbf4afbb6} /* (7, 23, 27) {real, imag} */,
  {32'h3f9841e6, 32'hbf8d9c0a} /* (7, 23, 26) {real, imag} */,
  {32'h3f0f4760, 32'hbf95f9c8} /* (7, 23, 25) {real, imag} */,
  {32'h3f84e5bc, 32'h3f29e91c} /* (7, 23, 24) {real, imag} */,
  {32'h3fa4a017, 32'h40192aa2} /* (7, 23, 23) {real, imag} */,
  {32'h3ec5e244, 32'h3fd46b80} /* (7, 23, 22) {real, imag} */,
  {32'h3f945588, 32'h3f640990} /* (7, 23, 21) {real, imag} */,
  {32'h3d169620, 32'h3fa36fb9} /* (7, 23, 20) {real, imag} */,
  {32'h3f81877a, 32'h3e026a36} /* (7, 23, 19) {real, imag} */,
  {32'h3ffeb2c0, 32'h3efb522d} /* (7, 23, 18) {real, imag} */,
  {32'h401040af, 32'h3fe23fc2} /* (7, 23, 17) {real, imag} */,
  {32'h3f5b814f, 32'h3f4a09c2} /* (7, 23, 16) {real, imag} */,
  {32'hbfde2f6f, 32'hbec475a4} /* (7, 23, 15) {real, imag} */,
  {32'hbf888d71, 32'hc01d96d8} /* (7, 23, 14) {real, imag} */,
  {32'hbf87ba68, 32'hbfef7971} /* (7, 23, 13) {real, imag} */,
  {32'hbff404d2, 32'hbf959064} /* (7, 23, 12) {real, imag} */,
  {32'hbfa08bfe, 32'hbf7de26c} /* (7, 23, 11) {real, imag} */,
  {32'h3fd7f2cf, 32'h3ea2538c} /* (7, 23, 10) {real, imag} */,
  {32'h3ff268eb, 32'hbe2e519f} /* (7, 23, 9) {real, imag} */,
  {32'h3f18c320, 32'hbf6b0fee} /* (7, 23, 8) {real, imag} */,
  {32'hbf474aba, 32'hbf8577c1} /* (7, 23, 7) {real, imag} */,
  {32'h3f17520c, 32'hbfea58a1} /* (7, 23, 6) {real, imag} */,
  {32'h3fd41ece, 32'hbff09530} /* (7, 23, 5) {real, imag} */,
  {32'hbe81ff28, 32'hbf8d6552} /* (7, 23, 4) {real, imag} */,
  {32'hbed6a758, 32'hc00b9490} /* (7, 23, 3) {real, imag} */,
  {32'h3f16657d, 32'h3f233aea} /* (7, 23, 2) {real, imag} */,
  {32'h4034314c, 32'h3fde341d} /* (7, 23, 1) {real, imag} */,
  {32'h3f407d46, 32'h3f26c838} /* (7, 23, 0) {real, imag} */,
  {32'h3fb79b7d, 32'hbe9c2dcf} /* (7, 22, 31) {real, imag} */,
  {32'h40044032, 32'hbfb75af6} /* (7, 22, 30) {real, imag} */,
  {32'h400330c4, 32'hbe191e20} /* (7, 22, 29) {real, imag} */,
  {32'hbe8a2994, 32'hbf92143a} /* (7, 22, 28) {real, imag} */,
  {32'hbf064bb8, 32'hbf9d5864} /* (7, 22, 27) {real, imag} */,
  {32'h3f92a61a, 32'hbf3f10ce} /* (7, 22, 26) {real, imag} */,
  {32'h3e9dc692, 32'hbc6a3100} /* (7, 22, 25) {real, imag} */,
  {32'h3eca997b, 32'h3eabbb56} /* (7, 22, 24) {real, imag} */,
  {32'hbfac1ebc, 32'h3f2dea52} /* (7, 22, 23) {real, imag} */,
  {32'hbfd9f5f3, 32'h3ffa2848} /* (7, 22, 22) {real, imag} */,
  {32'h3efcaeec, 32'h3e868811} /* (7, 22, 21) {real, imag} */,
  {32'h3e648d48, 32'hbf05329f} /* (7, 22, 20) {real, imag} */,
  {32'h3f86d549, 32'hc053ab83} /* (7, 22, 19) {real, imag} */,
  {32'hbd845508, 32'hbf9eb66f} /* (7, 22, 18) {real, imag} */,
  {32'h3fd87ada, 32'h3f06411e} /* (7, 22, 17) {real, imag} */,
  {32'h40225285, 32'hbee6583a} /* (7, 22, 16) {real, imag} */,
  {32'hbee0885c, 32'h3f5918fe} /* (7, 22, 15) {real, imag} */,
  {32'hbfd67223, 32'hbf7a4cfa} /* (7, 22, 14) {real, imag} */,
  {32'hbffa01d7, 32'hbfddc95a} /* (7, 22, 13) {real, imag} */,
  {32'h3f56c312, 32'hbfb46c18} /* (7, 22, 12) {real, imag} */,
  {32'h3f8350d6, 32'hbdbaf130} /* (7, 22, 11) {real, imag} */,
  {32'h3df4843c, 32'h3fbb5dc6} /* (7, 22, 10) {real, imag} */,
  {32'h3c8c4140, 32'h4018dc78} /* (7, 22, 9) {real, imag} */,
  {32'h3f20379e, 32'h3f52fce8} /* (7, 22, 8) {real, imag} */,
  {32'h3e2f2668, 32'h3fc3deed} /* (7, 22, 7) {real, imag} */,
  {32'h3d8398f8, 32'hbf8aa682} /* (7, 22, 6) {real, imag} */,
  {32'h3ff2b544, 32'hbfef11d5} /* (7, 22, 5) {real, imag} */,
  {32'h3f9f4452, 32'hbe1f418c} /* (7, 22, 4) {real, imag} */,
  {32'h4012a1a6, 32'h3f4d81dc} /* (7, 22, 3) {real, imag} */,
  {32'h3fc62a98, 32'h3fbe6c8c} /* (7, 22, 2) {real, imag} */,
  {32'h3f40abb6, 32'h3e4027e8} /* (7, 22, 1) {real, imag} */,
  {32'h3e940b43, 32'h3f2844d5} /* (7, 22, 0) {real, imag} */,
  {32'h3f7704f1, 32'h3f7f7e55} /* (7, 21, 31) {real, imag} */,
  {32'hbc68e3e0, 32'hbf34cca6} /* (7, 21, 30) {real, imag} */,
  {32'hbfb5601e, 32'hbf2f10ba} /* (7, 21, 29) {real, imag} */,
  {32'hc045af35, 32'hbf766773} /* (7, 21, 28) {real, imag} */,
  {32'hbf8f2b34, 32'hc0248de5} /* (7, 21, 27) {real, imag} */,
  {32'hbe966e08, 32'hbfc04564} /* (7, 21, 26) {real, imag} */,
  {32'hbfb908d4, 32'h3f02fddd} /* (7, 21, 25) {real, imag} */,
  {32'h3e023c74, 32'h3db45410} /* (7, 21, 24) {real, imag} */,
  {32'h3ea31f15, 32'hbf8c3a7f} /* (7, 21, 23) {real, imag} */,
  {32'h3e28df90, 32'hbfa5d5ec} /* (7, 21, 22) {real, imag} */,
  {32'h3ec6d2d7, 32'hbfbe8fff} /* (7, 21, 21) {real, imag} */,
  {32'h3ffa4ab0, 32'h3f2c8c09} /* (7, 21, 20) {real, imag} */,
  {32'h3ffb3b9c, 32'hbf5f1250} /* (7, 21, 19) {real, imag} */,
  {32'h3fad7c34, 32'hbf58d5e6} /* (7, 21, 18) {real, imag} */,
  {32'h3f9e8ad8, 32'hbe93a452} /* (7, 21, 17) {real, imag} */,
  {32'h3eaea62a, 32'hbf52b81f} /* (7, 21, 16) {real, imag} */,
  {32'hbe46df90, 32'h3d129c88} /* (7, 21, 15) {real, imag} */,
  {32'h3f0d37a6, 32'hbf1d17ff} /* (7, 21, 14) {real, imag} */,
  {32'h3fbabc8e, 32'h3e231d98} /* (7, 21, 13) {real, imag} */,
  {32'h3f61b892, 32'hbe85c28c} /* (7, 21, 12) {real, imag} */,
  {32'hbda45be0, 32'h3cfd1240} /* (7, 21, 11) {real, imag} */,
  {32'h3e9a07e6, 32'h3fbedee2} /* (7, 21, 10) {real, imag} */,
  {32'h403ac5e1, 32'h403b4f77} /* (7, 21, 9) {real, imag} */,
  {32'h401f3784, 32'h3fd12052} /* (7, 21, 8) {real, imag} */,
  {32'hbed8b152, 32'h3fc66819} /* (7, 21, 7) {real, imag} */,
  {32'hbfaf6e34, 32'h3dba2e3c} /* (7, 21, 6) {real, imag} */,
  {32'h3f5958c5, 32'h3ef528f5} /* (7, 21, 5) {real, imag} */,
  {32'h3f329604, 32'h3f40f4bc} /* (7, 21, 4) {real, imag} */,
  {32'h4003a2fa, 32'h3f9956d4} /* (7, 21, 3) {real, imag} */,
  {32'h3f0b2238, 32'h3fb208b9} /* (7, 21, 2) {real, imag} */,
  {32'hbe8ae62b, 32'hbfab5e90} /* (7, 21, 1) {real, imag} */,
  {32'hbd5f0488, 32'hbf6df0fe} /* (7, 21, 0) {real, imag} */,
  {32'h3ec222f2, 32'h3e814846} /* (7, 20, 31) {real, imag} */,
  {32'h3f2d28d4, 32'hbf4b0ffe} /* (7, 20, 30) {real, imag} */,
  {32'hbfaf6f0a, 32'hbf3c8b9a} /* (7, 20, 29) {real, imag} */,
  {32'hc033b117, 32'hbeeb0f86} /* (7, 20, 28) {real, imag} */,
  {32'hbfc05aca, 32'hbfe53bd4} /* (7, 20, 27) {real, imag} */,
  {32'hbf81afae, 32'hbf91f7f2} /* (7, 20, 26) {real, imag} */,
  {32'hbfab99ff, 32'h400c4c82} /* (7, 20, 25) {real, imag} */,
  {32'h3fbc662b, 32'h3fedfc05} /* (7, 20, 24) {real, imag} */,
  {32'h401ac61a, 32'hbf966456} /* (7, 20, 23) {real, imag} */,
  {32'h3f852a74, 32'hc0505892} /* (7, 20, 22) {real, imag} */,
  {32'h3ed077a8, 32'hc07287af} /* (7, 20, 21) {real, imag} */,
  {32'h3ff5bde2, 32'hbfd7fe67} /* (7, 20, 20) {real, imag} */,
  {32'h3f9108dd, 32'h3eb84738} /* (7, 20, 19) {real, imag} */,
  {32'h3f3ef7b0, 32'h3f45c61e} /* (7, 20, 18) {real, imag} */,
  {32'hbeb3e832, 32'h3ed1ee4c} /* (7, 20, 17) {real, imag} */,
  {32'h3e924a30, 32'hbf97f314} /* (7, 20, 16) {real, imag} */,
  {32'h3f674a81, 32'hbeaa48fa} /* (7, 20, 15) {real, imag} */,
  {32'h3fe8b48e, 32'hbfa969f5} /* (7, 20, 14) {real, imag} */,
  {32'h3fb0d3c4, 32'hbebc009e} /* (7, 20, 13) {real, imag} */,
  {32'h3f4eda6e, 32'hbf0e40d8} /* (7, 20, 12) {real, imag} */,
  {32'h401a3857, 32'h3ee4d320} /* (7, 20, 11) {real, imag} */,
  {32'h403ed83b, 32'h3fb9b1f4} /* (7, 20, 10) {real, imag} */,
  {32'h4054ccb9, 32'h3e8cd5d4} /* (7, 20, 9) {real, imag} */,
  {32'h400af2fa, 32'h3e84ff60} /* (7, 20, 8) {real, imag} */,
  {32'h3ed64a30, 32'hbde49c50} /* (7, 20, 7) {real, imag} */,
  {32'hbe85441e, 32'hbf52c06c} /* (7, 20, 6) {real, imag} */,
  {32'h3f1bc1b7, 32'h3f891c49} /* (7, 20, 5) {real, imag} */,
  {32'h3f689508, 32'h3e89a6ea} /* (7, 20, 4) {real, imag} */,
  {32'h3f828be0, 32'hbe841184} /* (7, 20, 3) {real, imag} */,
  {32'hbf5b6649, 32'hbf0d8fa1} /* (7, 20, 2) {real, imag} */,
  {32'h3e3fac8c, 32'hbf8289b3} /* (7, 20, 1) {real, imag} */,
  {32'hbdc37548, 32'hbf93f738} /* (7, 20, 0) {real, imag} */,
  {32'hbe0327d6, 32'h3eaeb760} /* (7, 19, 31) {real, imag} */,
  {32'h3fc6bf03, 32'h3d899b40} /* (7, 19, 30) {real, imag} */,
  {32'hbe0926d8, 32'h3ed454da} /* (7, 19, 29) {real, imag} */,
  {32'hbf94f579, 32'hbe68239c} /* (7, 19, 28) {real, imag} */,
  {32'hc01ee5f7, 32'hbed7437e} /* (7, 19, 27) {real, imag} */,
  {32'hbfd76a66, 32'hbf040031} /* (7, 19, 26) {real, imag} */,
  {32'hbe1c66f6, 32'h3fe8c48c} /* (7, 19, 25) {real, imag} */,
  {32'hbebd5839, 32'h3f4b04b0} /* (7, 19, 24) {real, imag} */,
  {32'hbfab45f9, 32'hbfce82e7} /* (7, 19, 23) {real, imag} */,
  {32'hbf2aec00, 32'hbfa7a7da} /* (7, 19, 22) {real, imag} */,
  {32'h3e241f80, 32'hc04571ca} /* (7, 19, 21) {real, imag} */,
  {32'h3f499a6c, 32'hbf4831e5} /* (7, 19, 20) {real, imag} */,
  {32'h3f2de360, 32'h3fc010ed} /* (7, 19, 19) {real, imag} */,
  {32'h3f0f90a7, 32'h3fc76e4c} /* (7, 19, 18) {real, imag} */,
  {32'hbfa3449a, 32'hbf737270} /* (7, 19, 17) {real, imag} */,
  {32'h3e98b592, 32'hbebc3571} /* (7, 19, 16) {real, imag} */,
  {32'h3f944889, 32'h3e1e1e26} /* (7, 19, 15) {real, imag} */,
  {32'h3f96cd84, 32'hbf2649e8} /* (7, 19, 14) {real, imag} */,
  {32'h3f1ff8c3, 32'hbf7df400} /* (7, 19, 13) {real, imag} */,
  {32'h3f166947, 32'hbfdc71d4} /* (7, 19, 12) {real, imag} */,
  {32'h3f5db09f, 32'h3f0531fe} /* (7, 19, 11) {real, imag} */,
  {32'h3e8f6176, 32'hbf2ea5ad} /* (7, 19, 10) {real, imag} */,
  {32'h3fd78390, 32'hc04aedd5} /* (7, 19, 9) {real, imag} */,
  {32'h3fbdf997, 32'hbff47783} /* (7, 19, 8) {real, imag} */,
  {32'h3f93e592, 32'hbfb2fbb4} /* (7, 19, 7) {real, imag} */,
  {32'h3e7a9cd8, 32'hbf900f4e} /* (7, 19, 6) {real, imag} */,
  {32'h3f387c69, 32'h3f5034ec} /* (7, 19, 5) {real, imag} */,
  {32'h404ddeb4, 32'h3e5468f6} /* (7, 19, 4) {real, imag} */,
  {32'h3f138393, 32'hbff78acc} /* (7, 19, 3) {real, imag} */,
  {32'hbfad7c7e, 32'hbf93ae00} /* (7, 19, 2) {real, imag} */,
  {32'h3f316a51, 32'hbef0a88a} /* (7, 19, 1) {real, imag} */,
  {32'h3e0c5e08, 32'h3edcfe07} /* (7, 19, 0) {real, imag} */,
  {32'h3f591882, 32'hbd9eac40} /* (7, 18, 31) {real, imag} */,
  {32'h401f86bb, 32'h3daf22a4} /* (7, 18, 30) {real, imag} */,
  {32'h3f552fc8, 32'h3fa1b477} /* (7, 18, 29) {real, imag} */,
  {32'hbebf60f4, 32'h402c19f8} /* (7, 18, 28) {real, imag} */,
  {32'hc029a9bd, 32'h3f99d8b2} /* (7, 18, 27) {real, imag} */,
  {32'hc04b5265, 32'h3f13d1d1} /* (7, 18, 26) {real, imag} */,
  {32'hbff91306, 32'hbe7b1ca4} /* (7, 18, 25) {real, imag} */,
  {32'hc044cf5c, 32'hbfb87e2b} /* (7, 18, 24) {real, imag} */,
  {32'hc049fa00, 32'hbfa51650} /* (7, 18, 23) {real, imag} */,
  {32'hbf858d7b, 32'hbf0d1ee4} /* (7, 18, 22) {real, imag} */,
  {32'h3dd732f0, 32'hbfa4f357} /* (7, 18, 21) {real, imag} */,
  {32'h3e1d2358, 32'hbe64d230} /* (7, 18, 20) {real, imag} */,
  {32'hbf237c08, 32'hbcdd5a50} /* (7, 18, 19) {real, imag} */,
  {32'h3ed19d68, 32'hbf9b72d2} /* (7, 18, 18) {real, imag} */,
  {32'h3e2b97b0, 32'hbe4e926e} /* (7, 18, 17) {real, imag} */,
  {32'h40051237, 32'h3d7d7640} /* (7, 18, 16) {real, imag} */,
  {32'h3f9d29e2, 32'hbf70d016} /* (7, 18, 15) {real, imag} */,
  {32'hbf83620e, 32'h3e88fc74} /* (7, 18, 14) {real, imag} */,
  {32'h3e362948, 32'hbfd23ae8} /* (7, 18, 13) {real, imag} */,
  {32'hbf0d9780, 32'hc0059b16} /* (7, 18, 12) {real, imag} */,
  {32'hbf4d9680, 32'hbfacf886} /* (7, 18, 11) {real, imag} */,
  {32'h3f02a132, 32'hc010a3ef} /* (7, 18, 10) {real, imag} */,
  {32'h3fc627c8, 32'h3e694508} /* (7, 18, 9) {real, imag} */,
  {32'h3ecc4778, 32'h40092811} /* (7, 18, 8) {real, imag} */,
  {32'h3fb46214, 32'h3fca458e} /* (7, 18, 7) {real, imag} */,
  {32'hbea992e2, 32'h3f2c3ee2} /* (7, 18, 6) {real, imag} */,
  {32'hbf995c68, 32'h3e4b4350} /* (7, 18, 5) {real, imag} */,
  {32'h3f39d7a2, 32'h3da2c700} /* (7, 18, 4) {real, imag} */,
  {32'h3f4dbd54, 32'hbf797c72} /* (7, 18, 3) {real, imag} */,
  {32'hbf45d323, 32'h3ed38b6c} /* (7, 18, 2) {real, imag} */,
  {32'hbf003dde, 32'h3da9a9e0} /* (7, 18, 1) {real, imag} */,
  {32'hbeb20614, 32'hbedbd9f6} /* (7, 18, 0) {real, imag} */,
  {32'h3fac5102, 32'hbf78a39c} /* (7, 17, 31) {real, imag} */,
  {32'h3fc2ef7c, 32'hbf06695a} /* (7, 17, 30) {real, imag} */,
  {32'hbfa75b46, 32'h3d0b24b0} /* (7, 17, 29) {real, imag} */,
  {32'hbf6cb1a1, 32'h3f030276} /* (7, 17, 28) {real, imag} */,
  {32'hc01ab8f5, 32'h3f1087d8} /* (7, 17, 27) {real, imag} */,
  {32'hc068d566, 32'h40390f91} /* (7, 17, 26) {real, imag} */,
  {32'hc039c38e, 32'h3fb90d3c} /* (7, 17, 25) {real, imag} */,
  {32'hc064b788, 32'hbe2d3ad0} /* (7, 17, 24) {real, imag} */,
  {32'hc045d406, 32'hbf05241e} /* (7, 17, 23) {real, imag} */,
  {32'hbfe44125, 32'hbef39964} /* (7, 17, 22) {real, imag} */,
  {32'hbec8f662, 32'h3fc6a2ea} /* (7, 17, 21) {real, imag} */,
  {32'h3edda1be, 32'hbd995bdc} /* (7, 17, 20) {real, imag} */,
  {32'h3dc45f6a, 32'hc0214f6b} /* (7, 17, 19) {real, imag} */,
  {32'h3ee82634, 32'hc05ef112} /* (7, 17, 18) {real, imag} */,
  {32'h3fa54513, 32'hbfb54a43} /* (7, 17, 17) {real, imag} */,
  {32'h3fcafccd, 32'h3bf2d580} /* (7, 17, 16) {real, imag} */,
  {32'hbfb3edf2, 32'hbf17213a} /* (7, 17, 15) {real, imag} */,
  {32'hbf278b24, 32'hbfb2d56c} /* (7, 17, 14) {real, imag} */,
  {32'h3e1815b8, 32'hc02899c0} /* (7, 17, 13) {real, imag} */,
  {32'hc05729df, 32'hc01cbda8} /* (7, 17, 12) {real, imag} */,
  {32'hbfcee157, 32'hbe8fe206} /* (7, 17, 11) {real, imag} */,
  {32'h3f53d424, 32'h4012f904} /* (7, 17, 10) {real, imag} */,
  {32'h3e5030f0, 32'h4025f8f9} /* (7, 17, 9) {real, imag} */,
  {32'hbf628548, 32'h3fd98a48} /* (7, 17, 8) {real, imag} */,
  {32'hbf77b0ee, 32'h40438266} /* (7, 17, 7) {real, imag} */,
  {32'hbfa16202, 32'h3f985e95} /* (7, 17, 6) {real, imag} */,
  {32'hbfd32582, 32'h3f5f93ee} /* (7, 17, 5) {real, imag} */,
  {32'hbd14c9e8, 32'h3f141444} /* (7, 17, 4) {real, imag} */,
  {32'h3fc9f370, 32'h3d499990} /* (7, 17, 3) {real, imag} */,
  {32'h3e6704ca, 32'h3eff71ea} /* (7, 17, 2) {real, imag} */,
  {32'hbf09aebc, 32'hbefec35c} /* (7, 17, 1) {real, imag} */,
  {32'h3dd1f0a0, 32'hbf886876} /* (7, 17, 0) {real, imag} */,
  {32'hbee2895d, 32'hbfa77912} /* (7, 16, 31) {real, imag} */,
  {32'h3d92f3a0, 32'h3f2bbb46} /* (7, 16, 30) {real, imag} */,
  {32'h3e9716ac, 32'h3e90bc58} /* (7, 16, 29) {real, imag} */,
  {32'hbf944950, 32'hbd8ff4c0} /* (7, 16, 28) {real, imag} */,
  {32'h3f3788a0, 32'h3fc25461} /* (7, 16, 27) {real, imag} */,
  {32'h3e06f830, 32'h4022b70f} /* (7, 16, 26) {real, imag} */,
  {32'h3f48862a, 32'h3fa44fd3} /* (7, 16, 25) {real, imag} */,
  {32'h3f9e63df, 32'h3f357a39} /* (7, 16, 24) {real, imag} */,
  {32'hbf1f6200, 32'h3db122c0} /* (7, 16, 23) {real, imag} */,
  {32'hbef7a89c, 32'hbf8241c1} /* (7, 16, 22) {real, imag} */,
  {32'hbd247e40, 32'h3f80c6da} /* (7, 16, 21) {real, imag} */,
  {32'h3eeeed98, 32'h3e9f9f60} /* (7, 16, 20) {real, imag} */,
  {32'hbcdfd2c0, 32'hc01341d2} /* (7, 16, 19) {real, imag} */,
  {32'hbdf21af8, 32'hc04b908d} /* (7, 16, 18) {real, imag} */,
  {32'h3fcfb7c4, 32'hbfc6aac2} /* (7, 16, 17) {real, imag} */,
  {32'h3e2817fc, 32'hbf5af5f4} /* (7, 16, 16) {real, imag} */,
  {32'hbfab79df, 32'hbf9a4ce4} /* (7, 16, 15) {real, imag} */,
  {32'h3f37f543, 32'hbf9c3e24} /* (7, 16, 14) {real, imag} */,
  {32'h3e98a534, 32'hc00c6d12} /* (7, 16, 13) {real, imag} */,
  {32'hbf14a69a, 32'h3f0d827f} /* (7, 16, 12) {real, imag} */,
  {32'h3ff15dfa, 32'h3d7c5d20} /* (7, 16, 11) {real, imag} */,
  {32'h3fdc8e32, 32'h3f3ef707} /* (7, 16, 10) {real, imag} */,
  {32'h403543d5, 32'h3fd35924} /* (7, 16, 9) {real, imag} */,
  {32'h3f85b580, 32'h404fde76} /* (7, 16, 8) {real, imag} */,
  {32'hbe534aa6, 32'h403e0bf2} /* (7, 16, 7) {real, imag} */,
  {32'hbfa32644, 32'hbf1e2b96} /* (7, 16, 6) {real, imag} */,
  {32'hbfa87286, 32'hbe4ca8f8} /* (7, 16, 5) {real, imag} */,
  {32'hbf3d466a, 32'h3e612b72} /* (7, 16, 4) {real, imag} */,
  {32'hbf6ac45c, 32'h3f4b7490} /* (7, 16, 3) {real, imag} */,
  {32'hbf271e44, 32'h3fa46ef5} /* (7, 16, 2) {real, imag} */,
  {32'h3fa2e2df, 32'h3f3f08a4} /* (7, 16, 1) {real, imag} */,
  {32'hbea15e60, 32'hbf145322} /* (7, 16, 0) {real, imag} */,
  {32'hbfa9a0b4, 32'hc012969f} /* (7, 15, 31) {real, imag} */,
  {32'hbf56f7c4, 32'hbdd99160} /* (7, 15, 30) {real, imag} */,
  {32'h3f9002fb, 32'hbfc9dd81} /* (7, 15, 29) {real, imag} */,
  {32'h3ef68dd0, 32'hbfb0c0f0} /* (7, 15, 28) {real, imag} */,
  {32'h3ff538d2, 32'h3f85e233} /* (7, 15, 27) {real, imag} */,
  {32'h3fd05509, 32'h4003787b} /* (7, 15, 26) {real, imag} */,
  {32'h3fc78926, 32'h4027a9c8} /* (7, 15, 25) {real, imag} */,
  {32'h3fe980a4, 32'h3fcefad2} /* (7, 15, 24) {real, imag} */,
  {32'hbf8cfbe7, 32'h3faab764} /* (7, 15, 23) {real, imag} */,
  {32'hbff64801, 32'hbf0f9100} /* (7, 15, 22) {real, imag} */,
  {32'hbfc23ca1, 32'hbff7fc55} /* (7, 15, 21) {real, imag} */,
  {32'h3f31d427, 32'hc0007d3e} /* (7, 15, 20) {real, imag} */,
  {32'h3fb785ed, 32'hbf2b784c} /* (7, 15, 19) {real, imag} */,
  {32'hbd3c1930, 32'hc024a97e} /* (7, 15, 18) {real, imag} */,
  {32'h3fabb40b, 32'hbfd8d066} /* (7, 15, 17) {real, imag} */,
  {32'h3eef0810, 32'hbfefec56} /* (7, 15, 16) {real, imag} */,
  {32'hbfa943c2, 32'hbf6f4f3e} /* (7, 15, 15) {real, imag} */,
  {32'hbfc8f92c, 32'hbeb2916c} /* (7, 15, 14) {real, imag} */,
  {32'hc0475cf4, 32'hbeab1bc7} /* (7, 15, 13) {real, imag} */,
  {32'hbfdcb3f5, 32'hbf419356} /* (7, 15, 12) {real, imag} */,
  {32'h3fc7e146, 32'hbf89f907} /* (7, 15, 11) {real, imag} */,
  {32'h3f6b5fed, 32'h3fa37d5a} /* (7, 15, 10) {real, imag} */,
  {32'h4009a1fb, 32'h402844ba} /* (7, 15, 9) {real, imag} */,
  {32'h3fc4ebd4, 32'h401ad136} /* (7, 15, 8) {real, imag} */,
  {32'h3fa1ec3b, 32'h3f6b8f30} /* (7, 15, 7) {real, imag} */,
  {32'h3e85d850, 32'hbf73b258} /* (7, 15, 6) {real, imag} */,
  {32'hbef140ae, 32'hbe87b553} /* (7, 15, 5) {real, imag} */,
  {32'hbededae8, 32'h3ef62720} /* (7, 15, 4) {real, imag} */,
  {32'hbfa07f51, 32'h3fa7c76e} /* (7, 15, 3) {real, imag} */,
  {32'hbf555668, 32'h3fb2fc7a} /* (7, 15, 2) {real, imag} */,
  {32'h3ff8cd47, 32'h3f56d6aa} /* (7, 15, 1) {real, imag} */,
  {32'h3f61fb3a, 32'hbda27180} /* (7, 15, 0) {real, imag} */,
  {32'h3ed7daac, 32'hbf03f862} /* (7, 14, 31) {real, imag} */,
  {32'h3e8ad90e, 32'h3e4eed48} /* (7, 14, 30) {real, imag} */,
  {32'h3ed68232, 32'h40074a5d} /* (7, 14, 29) {real, imag} */,
  {32'h3f371491, 32'h3ec28e6f} /* (7, 14, 28) {real, imag} */,
  {32'hbf80558a, 32'hbf418346} /* (7, 14, 27) {real, imag} */,
  {32'h3e72f064, 32'h3f9a747e} /* (7, 14, 26) {real, imag} */,
  {32'h3fa3d306, 32'h4007e594} /* (7, 14, 25) {real, imag} */,
  {32'h3fe13bc6, 32'h3fac1123} /* (7, 14, 24) {real, imag} */,
  {32'h3f5d19f6, 32'h3f37fe08} /* (7, 14, 23) {real, imag} */,
  {32'h3f6607e2, 32'h3f3437bc} /* (7, 14, 22) {real, imag} */,
  {32'h3f277d26, 32'h3f167704} /* (7, 14, 21) {real, imag} */,
  {32'hbf291b7c, 32'hbee952bc} /* (7, 14, 20) {real, imag} */,
  {32'h3f708766, 32'hbf322ba5} /* (7, 14, 19) {real, imag} */,
  {32'hbe64743c, 32'hbffe0b3c} /* (7, 14, 18) {real, imag} */,
  {32'hbf30454f, 32'hbf195d74} /* (7, 14, 17) {real, imag} */,
  {32'h3f74a05b, 32'hbfa06f82} /* (7, 14, 16) {real, imag} */,
  {32'hbfbfe443, 32'hbf5a705f} /* (7, 14, 15) {real, imag} */,
  {32'hbfcaa908, 32'hbf7dcf16} /* (7, 14, 14) {real, imag} */,
  {32'h3eb767b6, 32'hbf9a7e3c} /* (7, 14, 13) {real, imag} */,
  {32'h3f109198, 32'hc00bb12c} /* (7, 14, 12) {real, imag} */,
  {32'h3f931382, 32'hbf9d8624} /* (7, 14, 11) {real, imag} */,
  {32'h3ee0e6b9, 32'h3fdff212} /* (7, 14, 10) {real, imag} */,
  {32'h3fbd4cc6, 32'h3fe50055} /* (7, 14, 9) {real, imag} */,
  {32'h3fc56750, 32'hbf52a536} /* (7, 14, 8) {real, imag} */,
  {32'h400b3749, 32'hbdf53f50} /* (7, 14, 7) {real, imag} */,
  {32'h3fc59064, 32'h3e32f4ce} /* (7, 14, 6) {real, imag} */,
  {32'h3f1714f6, 32'hbf432c5c} /* (7, 14, 5) {real, imag} */,
  {32'hbcbe86c8, 32'h3ebf2dd9} /* (7, 14, 4) {real, imag} */,
  {32'hbf40e5d6, 32'h3ff34a10} /* (7, 14, 3) {real, imag} */,
  {32'hbfe3a70e, 32'h3fea2489} /* (7, 14, 2) {real, imag} */,
  {32'hbf31ea8a, 32'h4013bf20} /* (7, 14, 1) {real, imag} */,
  {32'h3fddfd76, 32'h3fcd4a2a} /* (7, 14, 0) {real, imag} */,
  {32'h3ee55966, 32'h3edc98bc} /* (7, 13, 31) {real, imag} */,
  {32'hbf1ce290, 32'h3d089358} /* (7, 13, 30) {real, imag} */,
  {32'hbf2fd704, 32'h3f0dc15b} /* (7, 13, 29) {real, imag} */,
  {32'h3f3ff07c, 32'hbf2be2e6} /* (7, 13, 28) {real, imag} */,
  {32'hbe851e2a, 32'hbfcbec6c} /* (7, 13, 27) {real, imag} */,
  {32'hbea37e10, 32'h3eaba59e} /* (7, 13, 26) {real, imag} */,
  {32'h3f27a74b, 32'h40042f6a} /* (7, 13, 25) {real, imag} */,
  {32'h3f36e286, 32'h3f202168} /* (7, 13, 24) {real, imag} */,
  {32'h3fbe2006, 32'hbf6cf9da} /* (7, 13, 23) {real, imag} */,
  {32'h4038a7e8, 32'h3f3a45ba} /* (7, 13, 22) {real, imag} */,
  {32'h404f1cae, 32'h3f58825a} /* (7, 13, 21) {real, imag} */,
  {32'hbf7a976c, 32'h3f77c6b2} /* (7, 13, 20) {real, imag} */,
  {32'hc01b9520, 32'hbfe76fba} /* (7, 13, 19) {real, imag} */,
  {32'hbfff794f, 32'hbf9fe219} /* (7, 13, 18) {real, imag} */,
  {32'hc0236762, 32'h3d685b00} /* (7, 13, 17) {real, imag} */,
  {32'hbfc1dc93, 32'hbf1c8eb6} /* (7, 13, 16) {real, imag} */,
  {32'hbf5533c8, 32'h3e646be0} /* (7, 13, 15) {real, imag} */,
  {32'h3e96916d, 32'h3edd9dea} /* (7, 13, 14) {real, imag} */,
  {32'h3f8f5795, 32'hbe0ca5be} /* (7, 13, 13) {real, imag} */,
  {32'h3f78db26, 32'hbf2584b0} /* (7, 13, 12) {real, imag} */,
  {32'h3fd40add, 32'h3f7ec947} /* (7, 13, 11) {real, imag} */,
  {32'h3df88b98, 32'h4035b3e6} /* (7, 13, 10) {real, imag} */,
  {32'h3e16b5c0, 32'h3fc908ef} /* (7, 13, 9) {real, imag} */,
  {32'hbe9c5454, 32'hbe761ff8} /* (7, 13, 8) {real, imag} */,
  {32'hbf083280, 32'h3eca2e70} /* (7, 13, 7) {real, imag} */,
  {32'h3fcb547c, 32'h3e1f7d57} /* (7, 13, 6) {real, imag} */,
  {32'h3fcd3a80, 32'hc003538c} /* (7, 13, 5) {real, imag} */,
  {32'hbf16ee16, 32'hbe1fd95c} /* (7, 13, 4) {real, imag} */,
  {32'hbf87f790, 32'h4003ddfe} /* (7, 13, 3) {real, imag} */,
  {32'hbfab7ae7, 32'h3fbd97c0} /* (7, 13, 2) {real, imag} */,
  {32'hbf965c7c, 32'h40174bb0} /* (7, 13, 1) {real, imag} */,
  {32'h3ecc3b68, 32'h3fdbb972} /* (7, 13, 0) {real, imag} */,
  {32'hbf56da6a, 32'h3f828d10} /* (7, 12, 31) {real, imag} */,
  {32'hc04cc0c0, 32'h3f5e2992} /* (7, 12, 30) {real, imag} */,
  {32'hc0098099, 32'h3eac049e} /* (7, 12, 29) {real, imag} */,
  {32'h3ebd68ac, 32'hc0011d48} /* (7, 12, 28) {real, imag} */,
  {32'h3f2169aa, 32'hbfa32672} /* (7, 12, 27) {real, imag} */,
  {32'hbed5440c, 32'hbe98f15c} /* (7, 12, 26) {real, imag} */,
  {32'hbeaabbd8, 32'h3f2ceb6b} /* (7, 12, 25) {real, imag} */,
  {32'hbf96172d, 32'h40055066} /* (7, 12, 24) {real, imag} */,
  {32'h3d268d50, 32'h3f8f2bdd} /* (7, 12, 23) {real, imag} */,
  {32'h3f3d96cc, 32'h3fc91971} /* (7, 12, 22) {real, imag} */,
  {32'h4027585c, 32'h3f8bc75c} /* (7, 12, 21) {real, imag} */,
  {32'h3fa03c78, 32'hbde1a4b8} /* (7, 12, 20) {real, imag} */,
  {32'hbf484d8e, 32'hc012e7a6} /* (7, 12, 19) {real, imag} */,
  {32'hbeae0928, 32'hbf8f9a32} /* (7, 12, 18) {real, imag} */,
  {32'hc015c328, 32'h3f050404} /* (7, 12, 17) {real, imag} */,
  {32'hc00731eb, 32'hbf87ba5c} /* (7, 12, 16) {real, imag} */,
  {32'h3f4a85d2, 32'h3f925ec7} /* (7, 12, 15) {real, imag} */,
  {32'h3f4e329c, 32'h3e9c25cc} /* (7, 12, 14) {real, imag} */,
  {32'hbf9ea922, 32'hbf6907e6} /* (7, 12, 13) {real, imag} */,
  {32'hbf234118, 32'hbfdffef9} /* (7, 12, 12) {real, imag} */,
  {32'h3f1458e0, 32'h3f9a65ce} /* (7, 12, 11) {real, imag} */,
  {32'hbf3ceb42, 32'h3fa75602} /* (7, 12, 10) {real, imag} */,
  {32'hbf7c7308, 32'hbf7ae16f} /* (7, 12, 9) {real, imag} */,
  {32'h3ea4060c, 32'h3e1c76a0} /* (7, 12, 8) {real, imag} */,
  {32'hbe8e3a34, 32'h3efe8912} /* (7, 12, 7) {real, imag} */,
  {32'h3f907e9b, 32'hbfbd80e8} /* (7, 12, 6) {real, imag} */,
  {32'h4035651b, 32'hbfb44f30} /* (7, 12, 5) {real, imag} */,
  {32'h3ea901d8, 32'h3e871dcf} /* (7, 12, 4) {real, imag} */,
  {32'hbf0b35d1, 32'hbf370c25} /* (7, 12, 3) {real, imag} */,
  {32'hbf7aa316, 32'h3f0e5f57} /* (7, 12, 2) {real, imag} */,
  {32'hbf637af1, 32'h402023c7} /* (7, 12, 1) {real, imag} */,
  {32'hbeb40b53, 32'h3f994033} /* (7, 12, 0) {real, imag} */,
  {32'hbf71e8cf, 32'h3f040cae} /* (7, 11, 31) {real, imag} */,
  {32'hbfbc1ff2, 32'hbf456cc1} /* (7, 11, 30) {real, imag} */,
  {32'hbfa7ec9f, 32'h3eb8fb16} /* (7, 11, 29) {real, imag} */,
  {32'hbf09db34, 32'hbf8906d2} /* (7, 11, 28) {real, imag} */,
  {32'hbf2f3602, 32'h3d83bb88} /* (7, 11, 27) {real, imag} */,
  {32'h3d3773e0, 32'h3f638189} /* (7, 11, 26) {real, imag} */,
  {32'h3f952231, 32'hbde32b38} /* (7, 11, 25) {real, imag} */,
  {32'hbf3bf695, 32'hbf17e9de} /* (7, 11, 24) {real, imag} */,
  {32'hbe6fff60, 32'h3faeaa2e} /* (7, 11, 23) {real, imag} */,
  {32'h3fae3351, 32'h3edad5a8} /* (7, 11, 22) {real, imag} */,
  {32'h3f07973e, 32'h3feaf2f6} /* (7, 11, 21) {real, imag} */,
  {32'hbd968490, 32'h3f8cb838} /* (7, 11, 20) {real, imag} */,
  {32'hbf051f95, 32'hc02ac1b0} /* (7, 11, 19) {real, imag} */,
  {32'h3ea80958, 32'hc0128a41} /* (7, 11, 18) {real, imag} */,
  {32'hbf2966ff, 32'h3f80877b} /* (7, 11, 17) {real, imag} */,
  {32'hbf8a80fc, 32'hc0433ec0} /* (7, 11, 16) {real, imag} */,
  {32'h3deff4e4, 32'hbfe8403c} /* (7, 11, 15) {real, imag} */,
  {32'hbfda3e4f, 32'hbf2c367e} /* (7, 11, 14) {real, imag} */,
  {32'hc00f0bf5, 32'hbf5cb702} /* (7, 11, 13) {real, imag} */,
  {32'hbf1f032e, 32'h3e5a1fe8} /* (7, 11, 12) {real, imag} */,
  {32'h3bb40400, 32'h3e518c18} /* (7, 11, 11) {real, imag} */,
  {32'hbf71eaff, 32'h3fa31589} /* (7, 11, 10) {real, imag} */,
  {32'hbfd980a2, 32'hbc2e7100} /* (7, 11, 9) {real, imag} */,
  {32'hc01a3db8, 32'h3f9abfd2} /* (7, 11, 8) {real, imag} */,
  {32'hc0349e4f, 32'h3f8851e0} /* (7, 11, 7) {real, imag} */,
  {32'hc00e7c50, 32'hbfef984e} /* (7, 11, 6) {real, imag} */,
  {32'h3ebc39e4, 32'h3d1cc900} /* (7, 11, 5) {real, imag} */,
  {32'hbd1bdca8, 32'h40206ce0} /* (7, 11, 4) {real, imag} */,
  {32'h3f350007, 32'h3fad0cb4} /* (7, 11, 3) {real, imag} */,
  {32'h3e8ab62c, 32'h3fce46ce} /* (7, 11, 2) {real, imag} */,
  {32'h3e946711, 32'h4001e8a2} /* (7, 11, 1) {real, imag} */,
  {32'hbeaae442, 32'h3f15cfe3} /* (7, 11, 0) {real, imag} */,
  {32'h3dbcef4e, 32'h3f085bbd} /* (7, 10, 31) {real, imag} */,
  {32'hbf0276e9, 32'hbf878be8} /* (7, 10, 30) {real, imag} */,
  {32'h3fd07793, 32'hc086ff07} /* (7, 10, 29) {real, imag} */,
  {32'hbf4ddc0a, 32'hbfa03486} /* (7, 10, 28) {real, imag} */,
  {32'hbff1146b, 32'h3dbd4c98} /* (7, 10, 27) {real, imag} */,
  {32'h3fe505a6, 32'h3e8ca096} /* (7, 10, 26) {real, imag} */,
  {32'h3f175ea2, 32'hbf156912} /* (7, 10, 25) {real, imag} */,
  {32'hbf03d49a, 32'hbfac3210} /* (7, 10, 24) {real, imag} */,
  {32'hbfa63862, 32'h3e272b18} /* (7, 10, 23) {real, imag} */,
  {32'h3fb9cac4, 32'hc010e3b8} /* (7, 10, 22) {real, imag} */,
  {32'hbfb6fcd7, 32'hbfa32840} /* (7, 10, 21) {real, imag} */,
  {32'hbff7b1c0, 32'h3fecfe11} /* (7, 10, 20) {real, imag} */,
  {32'hbf6fcc3e, 32'hbf57bda4} /* (7, 10, 19) {real, imag} */,
  {32'hc01095ee, 32'hc0190108} /* (7, 10, 18) {real, imag} */,
  {32'hbed67a14, 32'h3f61d735} /* (7, 10, 17) {real, imag} */,
  {32'h3ec6d5ca, 32'hbfed0042} /* (7, 10, 16) {real, imag} */,
  {32'hbe772338, 32'hc0752d7e} /* (7, 10, 15) {real, imag} */,
  {32'hbfac447d, 32'hc017b5d8} /* (7, 10, 14) {real, imag} */,
  {32'hbe47fec0, 32'hbed9df44} /* (7, 10, 13) {real, imag} */,
  {32'h3e525988, 32'h4026fae4} /* (7, 10, 12) {real, imag} */,
  {32'hbf2cf9c4, 32'h3f9ef54e} /* (7, 10, 11) {real, imag} */,
  {32'hc029f9f6, 32'h3f532651} /* (7, 10, 10) {real, imag} */,
  {32'hc00d8558, 32'h3f74b200} /* (7, 10, 9) {real, imag} */,
  {32'hbf9abbea, 32'h3ffc684c} /* (7, 10, 8) {real, imag} */,
  {32'hc0832a93, 32'hbeb83d40} /* (7, 10, 7) {real, imag} */,
  {32'hc03cc236, 32'hbf79f9f5} /* (7, 10, 6) {real, imag} */,
  {32'hbf85884e, 32'hbf980344} /* (7, 10, 5) {real, imag} */,
  {32'hbf131bec, 32'hbe83d3a4} /* (7, 10, 4) {real, imag} */,
  {32'h3fb8b905, 32'h3f52c829} /* (7, 10, 3) {real, imag} */,
  {32'h3f701ce2, 32'h3f380373} /* (7, 10, 2) {real, imag} */,
  {32'h3f269a5c, 32'h3f72a5da} /* (7, 10, 1) {real, imag} */,
  {32'h3d072554, 32'hbe935976} /* (7, 10, 0) {real, imag} */,
  {32'h3ea6e190, 32'h3f4e4785} /* (7, 9, 31) {real, imag} */,
  {32'hbfd2d0b2, 32'hbfbc4530} /* (7, 9, 30) {real, imag} */,
  {32'hbf3d0200, 32'hc084d786} /* (7, 9, 29) {real, imag} */,
  {32'hbfdeba38, 32'hbfee691f} /* (7, 9, 28) {real, imag} */,
  {32'hbe38ea84, 32'hbf8c6eed} /* (7, 9, 27) {real, imag} */,
  {32'h3f4c96e8, 32'h3e8f261d} /* (7, 9, 26) {real, imag} */,
  {32'hbf4b359c, 32'h3ff165dd} /* (7, 9, 25) {real, imag} */,
  {32'hbf897122, 32'h401a19e8} /* (7, 9, 24) {real, imag} */,
  {32'hbf9939e4, 32'hbf85592c} /* (7, 9, 23) {real, imag} */,
  {32'h3f3178a6, 32'hc02f8dec} /* (7, 9, 22) {real, imag} */,
  {32'h3ec1f42e, 32'hbf53df04} /* (7, 9, 21) {real, imag} */,
  {32'hbfb237e4, 32'h3ff27060} /* (7, 9, 20) {real, imag} */,
  {32'hc03d5650, 32'hbe24f2a8} /* (7, 9, 19) {real, imag} */,
  {32'hbffc59c4, 32'hbecc4434} /* (7, 9, 18) {real, imag} */,
  {32'h3dbb4e50, 32'h3f2b6422} /* (7, 9, 17) {real, imag} */,
  {32'h3f4e2e9a, 32'hbf500bc0} /* (7, 9, 16) {real, imag} */,
  {32'h3f492c93, 32'hc0434cae} /* (7, 9, 15) {real, imag} */,
  {32'hbf9668f2, 32'hc06a2816} /* (7, 9, 14) {real, imag} */,
  {32'hbd6d20e0, 32'hc03e5f33} /* (7, 9, 13) {real, imag} */,
  {32'h3f6488ea, 32'h3e360ce8} /* (7, 9, 12) {real, imag} */,
  {32'h3ecb6bde, 32'h3fd5729e} /* (7, 9, 11) {real, imag} */,
  {32'hbeb4e35c, 32'h3fc0768d} /* (7, 9, 10) {real, imag} */,
  {32'hbe9c5d70, 32'h3f1ccfba} /* (7, 9, 9) {real, imag} */,
  {32'hbf8b6ef6, 32'h3f676122} /* (7, 9, 8) {real, imag} */,
  {32'hc03eb8bc, 32'hbf56aa80} /* (7, 9, 7) {real, imag} */,
  {32'hbebba2b0, 32'hbf69bde0} /* (7, 9, 6) {real, imag} */,
  {32'h3f8d6848, 32'hbebbbe99} /* (7, 9, 5) {real, imag} */,
  {32'h3f7fcff4, 32'hc03010ec} /* (7, 9, 4) {real, imag} */,
  {32'h3f96e160, 32'hc029f073} /* (7, 9, 3) {real, imag} */,
  {32'hbd78ae80, 32'hbca57780} /* (7, 9, 2) {real, imag} */,
  {32'hbf81b1e4, 32'h3ea8a7c3} /* (7, 9, 1) {real, imag} */,
  {32'hbea73632, 32'hbe3a3a98} /* (7, 9, 0) {real, imag} */,
  {32'h3f0b0e56, 32'h3f7abf84} /* (7, 8, 31) {real, imag} */,
  {32'hbfd0ec63, 32'hbff66896} /* (7, 8, 30) {real, imag} */,
  {32'hbd666b80, 32'hbfd19dc8} /* (7, 8, 29) {real, imag} */,
  {32'hc000122a, 32'hbe359a42} /* (7, 8, 28) {real, imag} */,
  {32'hc001737a, 32'hbf88a9a4} /* (7, 8, 27) {real, imag} */,
  {32'hbf82054e, 32'hbf812153} /* (7, 8, 26) {real, imag} */,
  {32'hbe3e172f, 32'h400458e8} /* (7, 8, 25) {real, imag} */,
  {32'hbf164ba8, 32'h4085dde6} /* (7, 8, 24) {real, imag} */,
  {32'hbed3a1d8, 32'h3e3c5af8} /* (7, 8, 23) {real, imag} */,
  {32'h3f942633, 32'h3e869308} /* (7, 8, 22) {real, imag} */,
  {32'h3feb7d23, 32'hbf670090} /* (7, 8, 21) {real, imag} */,
  {32'h3f9a50e8, 32'hc00cdb71} /* (7, 8, 20) {real, imag} */,
  {32'hbffe02ff, 32'hbf969f5b} /* (7, 8, 19) {real, imag} */,
  {32'hbe91847f, 32'h3f7e56f6} /* (7, 8, 18) {real, imag} */,
  {32'hbd88aa78, 32'hbf065b96} /* (7, 8, 17) {real, imag} */,
  {32'hbf611d04, 32'hbff14604} /* (7, 8, 16) {real, imag} */,
  {32'h3ebc1994, 32'hc05b1157} /* (7, 8, 15) {real, imag} */,
  {32'hbf925db5, 32'hc0121aa6} /* (7, 8, 14) {real, imag} */,
  {32'hbfa07e10, 32'hbfad31e0} /* (7, 8, 13) {real, imag} */,
  {32'h3fea8b6f, 32'hbec67b58} /* (7, 8, 12) {real, imag} */,
  {32'h3ef09620, 32'hbf7190e0} /* (7, 8, 11) {real, imag} */,
  {32'h3f34fb1c, 32'h3b975000} /* (7, 8, 10) {real, imag} */,
  {32'h3ff84add, 32'hbe04adb0} /* (7, 8, 9) {real, imag} */,
  {32'h3e874ec8, 32'hbf6421f0} /* (7, 8, 8) {real, imag} */,
  {32'h3f9ed4af, 32'h3ffd7bd0} /* (7, 8, 7) {real, imag} */,
  {32'h3fd9b75e, 32'h3f0f952f} /* (7, 8, 6) {real, imag} */,
  {32'h3fcd75fd, 32'hbfaf85f9} /* (7, 8, 5) {real, imag} */,
  {32'hbf0add29, 32'hbfe1e01d} /* (7, 8, 4) {real, imag} */,
  {32'hbf54cb78, 32'hc02f13a8} /* (7, 8, 3) {real, imag} */,
  {32'h3eb3e2ec, 32'hbfb5ce5f} /* (7, 8, 2) {real, imag} */,
  {32'h3f945147, 32'hbf3d0a6c} /* (7, 8, 1) {real, imag} */,
  {32'h3ed68cec, 32'hbd040660} /* (7, 8, 0) {real, imag} */,
  {32'hbf3f1ae3, 32'hbf4abea3} /* (7, 7, 31) {real, imag} */,
  {32'hbf17b6ab, 32'hbfe6977a} /* (7, 7, 30) {real, imag} */,
  {32'h403ae15b, 32'hbfa115a3} /* (7, 7, 29) {real, imag} */,
  {32'h3fffd40b, 32'h3e3eaaf4} /* (7, 7, 28) {real, imag} */,
  {32'hbeb5b9fe, 32'hbf0d0913} /* (7, 7, 27) {real, imag} */,
  {32'hbe7deaf4, 32'hc03bdbad} /* (7, 7, 26) {real, imag} */,
  {32'hbf0573ba, 32'hbd55dea0} /* (7, 7, 25) {real, imag} */,
  {32'hbe8f6e32, 32'h4037efd4} /* (7, 7, 24) {real, imag} */,
  {32'h3f92ccb5, 32'h3f77d34c} /* (7, 7, 23) {real, imag} */,
  {32'h3fd74811, 32'h3f9859a6} /* (7, 7, 22) {real, imag} */,
  {32'hbe010878, 32'hc0074730} /* (7, 7, 21) {real, imag} */,
  {32'hbf2d603c, 32'hc09d8d02} /* (7, 7, 20) {real, imag} */,
  {32'h3eed0e46, 32'hbfb67800} /* (7, 7, 19) {real, imag} */,
  {32'h3ffebe02, 32'h3faa457c} /* (7, 7, 18) {real, imag} */,
  {32'h3e909bea, 32'hbf1e42a6} /* (7, 7, 17) {real, imag} */,
  {32'h3fdccdd1, 32'hbfc06252} /* (7, 7, 16) {real, imag} */,
  {32'h3f8706ce, 32'hbffa4b62} /* (7, 7, 15) {real, imag} */,
  {32'hbf637307, 32'h3bdebd80} /* (7, 7, 14) {real, imag} */,
  {32'hbfd537df, 32'h3f2312b2} /* (7, 7, 13) {real, imag} */,
  {32'h3f804050, 32'hbd094a00} /* (7, 7, 12) {real, imag} */,
  {32'h3fa2927e, 32'hc002a6e7} /* (7, 7, 11) {real, imag} */,
  {32'hbf24cb62, 32'hbebaa43c} /* (7, 7, 10) {real, imag} */,
  {32'h3f9b8a3e, 32'h3fb6c00c} /* (7, 7, 9) {real, imag} */,
  {32'hbe4aee3a, 32'h3e3af180} /* (7, 7, 8) {real, imag} */,
  {32'h3ffe4621, 32'h4006ae57} /* (7, 7, 7) {real, imag} */,
  {32'hbf24d720, 32'hbe250b94} /* (7, 7, 6) {real, imag} */,
  {32'h3ef01e34, 32'hbfe8d295} /* (7, 7, 5) {real, imag} */,
  {32'h3f30ccdc, 32'hbeb60f5b} /* (7, 7, 4) {real, imag} */,
  {32'h3d904410, 32'hc00ce86b} /* (7, 7, 3) {real, imag} */,
  {32'h3fbd03fe, 32'hbf5f5880} /* (7, 7, 2) {real, imag} */,
  {32'h4035e1e6, 32'h3f963df0} /* (7, 7, 1) {real, imag} */,
  {32'h3f516d8c, 32'h3f6191fc} /* (7, 7, 0) {real, imag} */,
  {32'hbe057844, 32'hbf8882fc} /* (7, 6, 31) {real, imag} */,
  {32'hbf71ed84, 32'hc0196b2b} /* (7, 6, 30) {real, imag} */,
  {32'hbf3d8851, 32'hbed4151c} /* (7, 6, 29) {real, imag} */,
  {32'h400a4a16, 32'h3f728c62} /* (7, 6, 28) {real, imag} */,
  {32'h402031de, 32'hbfa4caf4} /* (7, 6, 27) {real, imag} */,
  {32'h3c5ff040, 32'hbfd5a010} /* (7, 6, 26) {real, imag} */,
  {32'h3da27bb0, 32'hbd904ba0} /* (7, 6, 25) {real, imag} */,
  {32'hbeb4d0a0, 32'h3ec6e5e5} /* (7, 6, 24) {real, imag} */,
  {32'h3f89a74c, 32'h3f121aa6} /* (7, 6, 23) {real, imag} */,
  {32'h3f5418bc, 32'h3fbba6a2} /* (7, 6, 22) {real, imag} */,
  {32'h3df46050, 32'hbde104b8} /* (7, 6, 21) {real, imag} */,
  {32'h3ea07079, 32'hc01eca8e} /* (7, 6, 20) {real, imag} */,
  {32'hbf364e3b, 32'hbf916f95} /* (7, 6, 19) {real, imag} */,
  {32'h3f0bc0ea, 32'h3f8cb9a3} /* (7, 6, 18) {real, imag} */,
  {32'h4011d40c, 32'h3ec97d29} /* (7, 6, 17) {real, imag} */,
  {32'h40045af8, 32'hbf4e08b4} /* (7, 6, 16) {real, imag} */,
  {32'hbe8223fe, 32'h3ea234a7} /* (7, 6, 15) {real, imag} */,
  {32'hbe8b005b, 32'hbf566a6d} /* (7, 6, 14) {real, imag} */,
  {32'hc02a5c51, 32'hbfdfeaf0} /* (7, 6, 13) {real, imag} */,
  {32'hbf068f07, 32'hbed32bb0} /* (7, 6, 12) {real, imag} */,
  {32'h3fef8c1b, 32'hbf3441c8} /* (7, 6, 11) {real, imag} */,
  {32'h3fbbb156, 32'hbf55f3d3} /* (7, 6, 10) {real, imag} */,
  {32'h3f5fceb5, 32'h3f00345e} /* (7, 6, 9) {real, imag} */,
  {32'hc02ee8a2, 32'h3fc4c265} /* (7, 6, 8) {real, imag} */,
  {32'hbf648dce, 32'h400e447e} /* (7, 6, 7) {real, imag} */,
  {32'hbe1d85f0, 32'hbf7f3ad3} /* (7, 6, 6) {real, imag} */,
  {32'h3faa76fd, 32'hc014e267} /* (7, 6, 5) {real, imag} */,
  {32'h3fe4ac41, 32'hc04bec94} /* (7, 6, 4) {real, imag} */,
  {32'h3fb0354f, 32'hc008fc75} /* (7, 6, 3) {real, imag} */,
  {32'hbe6c8290, 32'hbf399906} /* (7, 6, 2) {real, imag} */,
  {32'h3f347812, 32'hbc4eb700} /* (7, 6, 1) {real, imag} */,
  {32'h3b14bb80, 32'hbed861e8} /* (7, 6, 0) {real, imag} */,
  {32'h3ee7e750, 32'h3ef01a2e} /* (7, 5, 31) {real, imag} */,
  {32'h3f1d4b9a, 32'hbf58c622} /* (7, 5, 30) {real, imag} */,
  {32'hbfcfa360, 32'h3f429e50} /* (7, 5, 29) {real, imag} */,
  {32'hbf94e611, 32'h3f3dfa67} /* (7, 5, 28) {real, imag} */,
  {32'h3f31eb80, 32'hbffd91c7} /* (7, 5, 27) {real, imag} */,
  {32'h3fa6cd10, 32'hbfb8576f} /* (7, 5, 26) {real, imag} */,
  {32'h3e7edc70, 32'hc0067f35} /* (7, 5, 25) {real, imag} */,
  {32'hbf8465a4, 32'hbff98907} /* (7, 5, 24) {real, imag} */,
  {32'hc004d290, 32'hbe5fc024} /* (7, 5, 23) {real, imag} */,
  {32'hbebd6270, 32'h3f08ba56} /* (7, 5, 22) {real, imag} */,
  {32'h3fe25224, 32'hbee9cf88} /* (7, 5, 21) {real, imag} */,
  {32'h3f494f61, 32'hc016868a} /* (7, 5, 20) {real, imag} */,
  {32'hc0490780, 32'hbf7f80be} /* (7, 5, 19) {real, imag} */,
  {32'hc0270934, 32'h3fd580fe} /* (7, 5, 18) {real, imag} */,
  {32'hbecff6a2, 32'h4004dd40} /* (7, 5, 17) {real, imag} */,
  {32'hbe3ebf3e, 32'hbf972e88} /* (7, 5, 16) {real, imag} */,
  {32'hbeb8ab4a, 32'hbf1fad74} /* (7, 5, 15) {real, imag} */,
  {32'hbe124b14, 32'h3d985ea8} /* (7, 5, 14) {real, imag} */,
  {32'hc013d509, 32'hbee21b90} /* (7, 5, 13) {real, imag} */,
  {32'hbf40ed50, 32'hbdf91b18} /* (7, 5, 12) {real, imag} */,
  {32'h3f097bf1, 32'h3ff6eb0b} /* (7, 5, 11) {real, imag} */,
  {32'h3d918490, 32'h3f92c842} /* (7, 5, 10) {real, imag} */,
  {32'hbf8d64c6, 32'hbca84300} /* (7, 5, 9) {real, imag} */,
  {32'hc04ff316, 32'h3fbd3c02} /* (7, 5, 8) {real, imag} */,
  {32'hbffe6458, 32'h4025fb16} /* (7, 5, 7) {real, imag} */,
  {32'h3fa9868b, 32'hbf507be5} /* (7, 5, 6) {real, imag} */,
  {32'h4027e931, 32'hbf89c314} /* (7, 5, 5) {real, imag} */,
  {32'h3ef7df34, 32'hc03b87a6} /* (7, 5, 4) {real, imag} */,
  {32'h3fdc4aac, 32'hbfc9d738} /* (7, 5, 3) {real, imag} */,
  {32'h3e3c6488, 32'hbf3a2fe8} /* (7, 5, 2) {real, imag} */,
  {32'hbf525f28, 32'h3fc55e0e} /* (7, 5, 1) {real, imag} */,
  {32'h3f335052, 32'h3f44b006} /* (7, 5, 0) {real, imag} */,
  {32'h3f036484, 32'h3faae32c} /* (7, 4, 31) {real, imag} */,
  {32'h3e843d50, 32'h3f24abc2} /* (7, 4, 30) {real, imag} */,
  {32'hbc4c66c0, 32'hbf9af1f6} /* (7, 4, 29) {real, imag} */,
  {32'hbf26a128, 32'hbfc6ff81} /* (7, 4, 28) {real, imag} */,
  {32'h3fee5f78, 32'hbe912116} /* (7, 4, 27) {real, imag} */,
  {32'h3f7c6d9a, 32'h3ebe6300} /* (7, 4, 26) {real, imag} */,
  {32'hbf83e2e6, 32'hbec64d50} /* (7, 4, 25) {real, imag} */,
  {32'hbdb04938, 32'hbeda57a9} /* (7, 4, 24) {real, imag} */,
  {32'hbfc235ea, 32'hbd8d7100} /* (7, 4, 23) {real, imag} */,
  {32'hbfabfb46, 32'h3fcd28dc} /* (7, 4, 22) {real, imag} */,
  {32'hbf6c5239, 32'h3fc6a57e} /* (7, 4, 21) {real, imag} */,
  {32'h3ed30140, 32'hbec5fcf8} /* (7, 4, 20) {real, imag} */,
  {32'hc031fba9, 32'hbe275406} /* (7, 4, 19) {real, imag} */,
  {32'hc044e03c, 32'h3ee7f6e8} /* (7, 4, 18) {real, imag} */,
  {32'hbf7683ce, 32'h3e29df70} /* (7, 4, 17) {real, imag} */,
  {32'h3f4049c2, 32'h3f9bee90} /* (7, 4, 16) {real, imag} */,
  {32'h3f84b6cf, 32'h4033f9d6} /* (7, 4, 15) {real, imag} */,
  {32'h3ea2087c, 32'h400f49af} /* (7, 4, 14) {real, imag} */,
  {32'hbfdae6c0, 32'h4002a88a} /* (7, 4, 13) {real, imag} */,
  {32'hbf8b4e30, 32'hbde48422} /* (7, 4, 12) {real, imag} */,
  {32'hbee9186e, 32'h3fd36037} /* (7, 4, 11) {real, imag} */,
  {32'hbedb104a, 32'hbed1e7c4} /* (7, 4, 10) {real, imag} */,
  {32'hbf2a8b7e, 32'hbf83e0ce} /* (7, 4, 9) {real, imag} */,
  {32'hc0133e2d, 32'h4020a836} /* (7, 4, 8) {real, imag} */,
  {32'hc0082ed2, 32'h400ee874} /* (7, 4, 7) {real, imag} */,
  {32'hbf9a96d2, 32'h3eafb481} /* (7, 4, 6) {real, imag} */,
  {32'hbe2aa7f0, 32'h3fe0a974} /* (7, 4, 5) {real, imag} */,
  {32'hbf8c2b29, 32'hbf9ae7bc} /* (7, 4, 4) {real, imag} */,
  {32'hbf16e942, 32'hbf52471f} /* (7, 4, 3) {real, imag} */,
  {32'h3f6eefeb, 32'h3ea789b8} /* (7, 4, 2) {real, imag} */,
  {32'hbef3b1e2, 32'h3f0b7532} /* (7, 4, 1) {real, imag} */,
  {32'h3f9da22e, 32'hbdab31d8} /* (7, 4, 0) {real, imag} */,
  {32'h3ea6b3d8, 32'h3ecf45a7} /* (7, 3, 31) {real, imag} */,
  {32'h3f5e45ff, 32'hbee74000} /* (7, 3, 30) {real, imag} */,
  {32'h3f906779, 32'hbfea1179} /* (7, 3, 29) {real, imag} */,
  {32'h3ffe079f, 32'hc01e3428} /* (7, 3, 28) {real, imag} */,
  {32'h40867072, 32'hbf4d42fe} /* (7, 3, 27) {real, imag} */,
  {32'h3fa8916a, 32'h3f8c24b6} /* (7, 3, 26) {real, imag} */,
  {32'hbdba8fb0, 32'h3f5913b5} /* (7, 3, 25) {real, imag} */,
  {32'h3f99f02a, 32'h4014f98f} /* (7, 3, 24) {real, imag} */,
  {32'hbf67eada, 32'h3faa03fa} /* (7, 3, 23) {real, imag} */,
  {32'hbfebcade, 32'h3fa31f1c} /* (7, 3, 22) {real, imag} */,
  {32'h3f24186c, 32'h3f8f205a} /* (7, 3, 21) {real, imag} */,
  {32'h4024fec6, 32'h3f616a14} /* (7, 3, 20) {real, imag} */,
  {32'hbddc5998, 32'h4003e618} /* (7, 3, 19) {real, imag} */,
  {32'hc004f228, 32'hbfbc9ddf} /* (7, 3, 18) {real, imag} */,
  {32'h3ece5088, 32'hc001b6e8} /* (7, 3, 17) {real, imag} */,
  {32'h3fa6f2e6, 32'h3ea7a875} /* (7, 3, 16) {real, imag} */,
  {32'h3f39846e, 32'h40783dee} /* (7, 3, 15) {real, imag} */,
  {32'h3faf4291, 32'h4088a319} /* (7, 3, 14) {real, imag} */,
  {32'hbf4bd963, 32'h3f09d3ba} /* (7, 3, 13) {real, imag} */,
  {32'hbf237f4c, 32'hbfce2cec} /* (7, 3, 12) {real, imag} */,
  {32'hc000889a, 32'h3f165add} /* (7, 3, 11) {real, imag} */,
  {32'hbf38c3d5, 32'hbf17ef3e} /* (7, 3, 10) {real, imag} */,
  {32'hbf958a5d, 32'hbfb35d14} /* (7, 3, 9) {real, imag} */,
  {32'hbfadacba, 32'h3f86f743} /* (7, 3, 8) {real, imag} */,
  {32'hbf874efc, 32'hbeb0c2ec} /* (7, 3, 7) {real, imag} */,
  {32'h3e51e4e0, 32'h3f11fd61} /* (7, 3, 6) {real, imag} */,
  {32'h3f64dea1, 32'h4046ee91} /* (7, 3, 5) {real, imag} */,
  {32'hbf44cfec, 32'hbe267f10} /* (7, 3, 4) {real, imag} */,
  {32'hbf8f0385, 32'hbfba6d5d} /* (7, 3, 3) {real, imag} */,
  {32'hbf8c1708, 32'h3ea85cec} /* (7, 3, 2) {real, imag} */,
  {32'h3fd395c5, 32'h3efa3420} /* (7, 3, 1) {real, imag} */,
  {32'h3fc35abd, 32'hbed0eba0} /* (7, 3, 0) {real, imag} */,
  {32'hbf4e6a75, 32'hbe4702ee} /* (7, 2, 31) {real, imag} */,
  {32'h3e97e542, 32'hbf684344} /* (7, 2, 30) {real, imag} */,
  {32'h3e081caa, 32'hbf8101ca} /* (7, 2, 29) {real, imag} */,
  {32'h3f134ed9, 32'hbef3d4d6} /* (7, 2, 28) {real, imag} */,
  {32'h3fe451b3, 32'h3f4d1504} /* (7, 2, 27) {real, imag} */,
  {32'h3dafeeb0, 32'h3fe8a074} /* (7, 2, 26) {real, imag} */,
  {32'h3f0eeefc, 32'h3fc55d90} /* (7, 2, 25) {real, imag} */,
  {32'h4019c1e8, 32'h40423fa3} /* (7, 2, 24) {real, imag} */,
  {32'hbf9205bc, 32'h3fd2696e} /* (7, 2, 23) {real, imag} */,
  {32'hbfa8ca9e, 32'hbe8df8dc} /* (7, 2, 22) {real, imag} */,
  {32'h3fc037f5, 32'hbf844cfe} /* (7, 2, 21) {real, imag} */,
  {32'h3fbf1d47, 32'hbd97f7d4} /* (7, 2, 20) {real, imag} */,
  {32'h3ea83b3b, 32'h3fc8ebb8} /* (7, 2, 19) {real, imag} */,
  {32'hbfce007e, 32'hbf7d155e} /* (7, 2, 18) {real, imag} */,
  {32'hbeafd307, 32'hbf8dd544} /* (7, 2, 17) {real, imag} */,
  {32'hbf6e7ebe, 32'h3f1d5ce0} /* (7, 2, 16) {real, imag} */,
  {32'hc020584a, 32'h4037a6d0} /* (7, 2, 15) {real, imag} */,
  {32'hbf86f7e2, 32'h405bbe0f} /* (7, 2, 14) {real, imag} */,
  {32'hbf48b442, 32'hbf74a392} /* (7, 2, 13) {real, imag} */,
  {32'hbed6c818, 32'hc015c5d5} /* (7, 2, 12) {real, imag} */,
  {32'hbec529c8, 32'hbea46598} /* (7, 2, 11) {real, imag} */,
  {32'hc0145114, 32'hbdd12768} /* (7, 2, 10) {real, imag} */,
  {32'hc0659e2e, 32'hbfe4e40e} /* (7, 2, 9) {real, imag} */,
  {32'hbd2db750, 32'hbf31ed38} /* (7, 2, 8) {real, imag} */,
  {32'h3edc3ae0, 32'hbf804e1b} /* (7, 2, 7) {real, imag} */,
  {32'h3f919348, 32'hbfbbf67e} /* (7, 2, 6) {real, imag} */,
  {32'h3f8a8eba, 32'h4001366c} /* (7, 2, 5) {real, imag} */,
  {32'hbf046330, 32'h4034baab} /* (7, 2, 4) {real, imag} */,
  {32'h3d5d2da0, 32'h3fd7cf47} /* (7, 2, 3) {real, imag} */,
  {32'h3e8a51fe, 32'h3f76add2} /* (7, 2, 2) {real, imag} */,
  {32'h3f149fd7, 32'h3fd52142} /* (7, 2, 1) {real, imag} */,
  {32'hbefb606c, 32'h3f7646d3} /* (7, 2, 0) {real, imag} */,
  {32'hbee3eacf, 32'h3f219ae4} /* (7, 1, 31) {real, imag} */,
  {32'h3ee77ea4, 32'hbd91440c} /* (7, 1, 30) {real, imag} */,
  {32'h3ebae542, 32'hbffc3201} /* (7, 1, 29) {real, imag} */,
  {32'h3fdf95a4, 32'hbfa308b8} /* (7, 1, 28) {real, imag} */,
  {32'h3f1cf6d8, 32'h3f0a349d} /* (7, 1, 27) {real, imag} */,
  {32'hbf6d26dc, 32'h3f872f64} /* (7, 1, 26) {real, imag} */,
  {32'hbe60c8d8, 32'h3f2ae6fe} /* (7, 1, 25) {real, imag} */,
  {32'h3fe1cc28, 32'h3fa26b7c} /* (7, 1, 24) {real, imag} */,
  {32'hbc9601a0, 32'hbe2405b0} /* (7, 1, 23) {real, imag} */,
  {32'h3f8567fb, 32'hc00fda00} /* (7, 1, 22) {real, imag} */,
  {32'h3f8a39d2, 32'hc016e08e} /* (7, 1, 21) {real, imag} */,
  {32'hbe86f49e, 32'hbf7d2ebe} /* (7, 1, 20) {real, imag} */,
  {32'h3f1c1efd, 32'h3f16a2fd} /* (7, 1, 19) {real, imag} */,
  {32'hbfe67871, 32'hbe9652c8} /* (7, 1, 18) {real, imag} */,
  {32'hbfd239ca, 32'hbea07b2c} /* (7, 1, 17) {real, imag} */,
  {32'h3e318fc8, 32'hbeecf2eb} /* (7, 1, 16) {real, imag} */,
  {32'hbe85b3ae, 32'hbe91038a} /* (7, 1, 15) {real, imag} */,
  {32'hbe8dc553, 32'h3f5ff5f4} /* (7, 1, 14) {real, imag} */,
  {32'hbfee67f9, 32'h4015832d} /* (7, 1, 13) {real, imag} */,
  {32'hbfe979eb, 32'h3f2a629c} /* (7, 1, 12) {real, imag} */,
  {32'h3e53c854, 32'hbf1301a8} /* (7, 1, 11) {real, imag} */,
  {32'hc01dce47, 32'hbe873b8a} /* (7, 1, 10) {real, imag} */,
  {32'hc0284bac, 32'hc01277fc} /* (7, 1, 9) {real, imag} */,
  {32'h3f727250, 32'hbfeebd90} /* (7, 1, 8) {real, imag} */,
  {32'h3fbc31af, 32'hbf63d29a} /* (7, 1, 7) {real, imag} */,
  {32'h3eac26d0, 32'hbf8c49a8} /* (7, 1, 6) {real, imag} */,
  {32'h3f0b2831, 32'h3fb4671b} /* (7, 1, 5) {real, imag} */,
  {32'hbe3e9988, 32'h405a8bce} /* (7, 1, 4) {real, imag} */,
  {32'hbfd4ea4e, 32'h4021149c} /* (7, 1, 3) {real, imag} */,
  {32'h3f05931a, 32'h3ea3ff92} /* (7, 1, 2) {real, imag} */,
  {32'h3f2f0e72, 32'h3f8baef6} /* (7, 1, 1) {real, imag} */,
  {32'h3e788d04, 32'h40049185} /* (7, 1, 0) {real, imag} */,
  {32'hbf76eca2, 32'h3f1a9764} /* (7, 0, 31) {real, imag} */,
  {32'hbeff48d0, 32'h3d557c08} /* (7, 0, 30) {real, imag} */,
  {32'hbf702360, 32'hbfd2d172} /* (7, 0, 29) {real, imag} */,
  {32'h3f3ef1e6, 32'hbf973008} /* (7, 0, 28) {real, imag} */,
  {32'h3e1f62ec, 32'hbf1f0c04} /* (7, 0, 27) {real, imag} */,
  {32'hbf9adecb, 32'h3ebd8352} /* (7, 0, 26) {real, imag} */,
  {32'hbe8c0b94, 32'h3c952180} /* (7, 0, 25) {real, imag} */,
  {32'h3fab9e82, 32'h3e962dbe} /* (7, 0, 24) {real, imag} */,
  {32'h3f20ad12, 32'h3c776c20} /* (7, 0, 23) {real, imag} */,
  {32'h3f957e54, 32'hbf2163be} /* (7, 0, 22) {real, imag} */,
  {32'h3e97d5d0, 32'hbf7e2464} /* (7, 0, 21) {real, imag} */,
  {32'hbef1a132, 32'hbf4092e1} /* (7, 0, 20) {real, imag} */,
  {32'hbde8b260, 32'h3f915024} /* (7, 0, 19) {real, imag} */,
  {32'hbd9d435a, 32'h3f1ad1a9} /* (7, 0, 18) {real, imag} */,
  {32'hbf25d009, 32'hbe0d4878} /* (7, 0, 17) {real, imag} */,
  {32'h3e2ffbb0, 32'hbf9a9129} /* (7, 0, 16) {real, imag} */,
  {32'h3f30431c, 32'hbf454ee2} /* (7, 0, 15) {real, imag} */,
  {32'h3fdcfe79, 32'hbe904fe0} /* (7, 0, 14) {real, imag} */,
  {32'hbf3862c8, 32'h4027f8e0} /* (7, 0, 13) {real, imag} */,
  {32'hbfb1eaa0, 32'h3ff4ce91} /* (7, 0, 12) {real, imag} */,
  {32'hbf903dac, 32'h3f195238} /* (7, 0, 11) {real, imag} */,
  {32'hbfcea005, 32'hbfaf75b2} /* (7, 0, 10) {real, imag} */,
  {32'hbf6101e6, 32'hbf4f9054} /* (7, 0, 9) {real, imag} */,
  {32'h3f330295, 32'hbf424038} /* (7, 0, 8) {real, imag} */,
  {32'h3f05c102, 32'hbe8c1926} /* (7, 0, 7) {real, imag} */,
  {32'hbfa660ef, 32'h3ec5ac5b} /* (7, 0, 6) {real, imag} */,
  {32'hbe54d64e, 32'h3f7159b1} /* (7, 0, 5) {real, imag} */,
  {32'h3eeb5784, 32'h3f853738} /* (7, 0, 4) {real, imag} */,
  {32'hbf906bfa, 32'h3e5922e9} /* (7, 0, 3) {real, imag} */,
  {32'hbea86ada, 32'hbf86a56c} /* (7, 0, 2) {real, imag} */,
  {32'h3ddbf910, 32'h3caa3080} /* (7, 0, 1) {real, imag} */,
  {32'hbddc8db4, 32'h3fb21a1a} /* (7, 0, 0) {real, imag} */,
  {32'h3eb8ed12, 32'hbeafd44d} /* (6, 31, 31) {real, imag} */,
  {32'h3f1f0261, 32'h3e7a1fa0} /* (6, 31, 30) {real, imag} */,
  {32'hbf39ba04, 32'h3fc854b0} /* (6, 31, 29) {real, imag} */,
  {32'h3f3c28c2, 32'h3e8f6842} /* (6, 31, 28) {real, imag} */,
  {32'h40411b32, 32'hbf223875} /* (6, 31, 27) {real, imag} */,
  {32'h3fb1dd32, 32'hc0282e34} /* (6, 31, 26) {real, imag} */,
  {32'h3f17ad3a, 32'hbf4183bb} /* (6, 31, 25) {real, imag} */,
  {32'hbf2e28be, 32'h3f8a685a} /* (6, 31, 24) {real, imag} */,
  {32'h3da1db08, 32'h3cd7fd20} /* (6, 31, 23) {real, imag} */,
  {32'hbf2b29da, 32'h3fe38665} /* (6, 31, 22) {real, imag} */,
  {32'hbf0f29a9, 32'h4021feb9} /* (6, 31, 21) {real, imag} */,
  {32'hc01a9a83, 32'h3ec1c3f1} /* (6, 31, 20) {real, imag} */,
  {32'hc014360e, 32'h3fe36b9f} /* (6, 31, 19) {real, imag} */,
  {32'hbf640bfc, 32'h3feaf9c5} /* (6, 31, 18) {real, imag} */,
  {32'hbf8802a5, 32'hbd8ab4a0} /* (6, 31, 17) {real, imag} */,
  {32'hbf539d04, 32'hbf2703fe} /* (6, 31, 16) {real, imag} */,
  {32'hbf915c2e, 32'hbffc1407} /* (6, 31, 15) {real, imag} */,
  {32'hbfb94b35, 32'hbfcc79fb} /* (6, 31, 14) {real, imag} */,
  {32'hbfa26463, 32'hbe8c92f0} /* (6, 31, 13) {real, imag} */,
  {32'hbd8278c0, 32'hbd0242e0} /* (6, 31, 12) {real, imag} */,
  {32'hbec7de23, 32'hbf229546} /* (6, 31, 11) {real, imag} */,
  {32'h3f723f84, 32'hc01141ba} /* (6, 31, 10) {real, imag} */,
  {32'h3f7eace8, 32'hbeeacf04} /* (6, 31, 9) {real, imag} */,
  {32'h3fcd1d5f, 32'h3f8ca9b2} /* (6, 31, 8) {real, imag} */,
  {32'hbf40fb5e, 32'hbef54444} /* (6, 31, 7) {real, imag} */,
  {32'h3f36fdbd, 32'hbc12aa80} /* (6, 31, 6) {real, imag} */,
  {32'h3f9d1f9e, 32'hbe89a1b4} /* (6, 31, 5) {real, imag} */,
  {32'hbe06e804, 32'hbfe55ae2} /* (6, 31, 4) {real, imag} */,
  {32'h3f403b5f, 32'hbfbda512} /* (6, 31, 3) {real, imag} */,
  {32'h40422443, 32'hbf0790c1} /* (6, 31, 2) {real, imag} */,
  {32'h40368687, 32'hbd1ac280} /* (6, 31, 1) {real, imag} */,
  {32'h3ff823fb, 32'h3e524754} /* (6, 31, 0) {real, imag} */,
  {32'h3f53d6c4, 32'hbf02b434} /* (6, 30, 31) {real, imag} */,
  {32'h3ff07be2, 32'h3e19cc40} /* (6, 30, 30) {real, imag} */,
  {32'hbf1b04ce, 32'h400cb18c} /* (6, 30, 29) {real, imag} */,
  {32'h3eafd1dc, 32'h3f00e864} /* (6, 30, 28) {real, imag} */,
  {32'h40460ee6, 32'hbf36e17e} /* (6, 30, 27) {real, imag} */,
  {32'h401aedaa, 32'hc0165540} /* (6, 30, 26) {real, imag} */,
  {32'hbf36faec, 32'hbf67edac} /* (6, 30, 25) {real, imag} */,
  {32'hbf820cdc, 32'h3fbd55da} /* (6, 30, 24) {real, imag} */,
  {32'hbf2c724c, 32'hbfa9cc66} /* (6, 30, 23) {real, imag} */,
  {32'hbfcee29f, 32'h3e97bfb8} /* (6, 30, 22) {real, imag} */,
  {32'hbe7ee898, 32'h40793ec1} /* (6, 30, 21) {real, imag} */,
  {32'hbd0f5e00, 32'h4007de78} /* (6, 30, 20) {real, imag} */,
  {32'hbf3389d3, 32'h40363e8f} /* (6, 30, 19) {real, imag} */,
  {32'hbeeae7e6, 32'h404a6128} /* (6, 30, 18) {real, imag} */,
  {32'hbfa6dab1, 32'h3fcd4105} /* (6, 30, 17) {real, imag} */,
  {32'hbf6da475, 32'h3ec20cba} /* (6, 30, 16) {real, imag} */,
  {32'hbe3e7d1c, 32'h3bab4700} /* (6, 30, 15) {real, imag} */,
  {32'hbff6adf8, 32'h3f918d4d} /* (6, 30, 14) {real, imag} */,
  {32'hbf432c20, 32'hbf1f0616} /* (6, 30, 13) {real, imag} */,
  {32'hbf49baab, 32'hc009c74e} /* (6, 30, 12) {real, imag} */,
  {32'hbfc3c1d9, 32'hbf4b7660} /* (6, 30, 11) {real, imag} */,
  {32'h3e424ea4, 32'hbfa75274} /* (6, 30, 10) {real, imag} */,
  {32'hbed17bee, 32'hbf0ff126} /* (6, 30, 9) {real, imag} */,
  {32'h3f87b600, 32'h3f5085c2} /* (6, 30, 8) {real, imag} */,
  {32'h3fd56919, 32'hbfc79813} /* (6, 30, 7) {real, imag} */,
  {32'h3ec175c0, 32'hbfd352e5} /* (6, 30, 6) {real, imag} */,
  {32'hbeff6108, 32'hbea7c080} /* (6, 30, 5) {real, imag} */,
  {32'h3f0625ca, 32'hbff99898} /* (6, 30, 4) {real, imag} */,
  {32'h3fd1c968, 32'hc018cb4a} /* (6, 30, 3) {real, imag} */,
  {32'h3fe3d8a6, 32'hbf5f5530} /* (6, 30, 2) {real, imag} */,
  {32'hbf879fae, 32'h3eb40b58} /* (6, 30, 1) {real, imag} */,
  {32'hbf7479e0, 32'h3ffcc0ac} /* (6, 30, 0) {real, imag} */,
  {32'h3f258f1e, 32'h3e4db7dc} /* (6, 29, 31) {real, imag} */,
  {32'h3e91ac6c, 32'hbeb5ef50} /* (6, 29, 30) {real, imag} */,
  {32'hbf3a2dd6, 32'h3df6b610} /* (6, 29, 29) {real, imag} */,
  {32'h3fbf73a2, 32'h3e94f58c} /* (6, 29, 28) {real, imag} */,
  {32'h402ef59b, 32'h3e20baec} /* (6, 29, 27) {real, imag} */,
  {32'h3fd82dac, 32'hc010824a} /* (6, 29, 26) {real, imag} */,
  {32'hbd4a2210, 32'hbfeccc6a} /* (6, 29, 25) {real, imag} */,
  {32'h3fda64de, 32'h3fba0b9e} /* (6, 29, 24) {real, imag} */,
  {32'hbf81a156, 32'hbf4dda1c} /* (6, 29, 23) {real, imag} */,
  {32'hbeb35b82, 32'h3dc1a8c0} /* (6, 29, 22) {real, imag} */,
  {32'h3f8db77a, 32'h3fea45a8} /* (6, 29, 21) {real, imag} */,
  {32'h3fb995fc, 32'h406e444a} /* (6, 29, 20) {real, imag} */,
  {32'hbe2f5924, 32'h40296a64} /* (6, 29, 19) {real, imag} */,
  {32'hbf2c4174, 32'h3fac4ad1} /* (6, 29, 18) {real, imag} */,
  {32'h3fb0ce7e, 32'h3f5678ef} /* (6, 29, 17) {real, imag} */,
  {32'h3fba8f14, 32'hc00d16ec} /* (6, 29, 16) {real, imag} */,
  {32'h401e72fa, 32'hc0007709} /* (6, 29, 15) {real, imag} */,
  {32'h403f8adc, 32'h3fafd9f4} /* (6, 29, 14) {real, imag} */,
  {32'h4014fabc, 32'h3f0fba90} /* (6, 29, 13) {real, imag} */,
  {32'hbef34fae, 32'hbedcb68c} /* (6, 29, 12) {real, imag} */,
  {32'hbf3cc61c, 32'hbf25540e} /* (6, 29, 11) {real, imag} */,
  {32'h3e88cdd4, 32'hbf9de02a} /* (6, 29, 10) {real, imag} */,
  {32'hbf97f64b, 32'hbf46646a} /* (6, 29, 9) {real, imag} */,
  {32'h3f8aec04, 32'h3e5439a8} /* (6, 29, 8) {real, imag} */,
  {32'h40525093, 32'hc006f804} /* (6, 29, 7) {real, imag} */,
  {32'hbf3d7286, 32'hc00e1940} /* (6, 29, 6) {real, imag} */,
  {32'hc00e9236, 32'h3f5de2cf} /* (6, 29, 5) {real, imag} */,
  {32'h3dc4e7a0, 32'h3f6c5e0a} /* (6, 29, 4) {real, imag} */,
  {32'h3f83e598, 32'hbf4462fa} /* (6, 29, 3) {real, imag} */,
  {32'hbfe570d2, 32'hbed9ed38} /* (6, 29, 2) {real, imag} */,
  {32'hc04ba56d, 32'h3ef74d6a} /* (6, 29, 1) {real, imag} */,
  {32'hbf3b00a3, 32'h3fbafe72} /* (6, 29, 0) {real, imag} */,
  {32'h3ec67e6c, 32'h40203788} /* (6, 28, 31) {real, imag} */,
  {32'hbfa10bdc, 32'h3f20461a} /* (6, 28, 30) {real, imag} */,
  {32'hbf1bb9a8, 32'hbf9e18f8} /* (6, 28, 29) {real, imag} */,
  {32'h400e78d6, 32'hbfb10c9c} /* (6, 28, 28) {real, imag} */,
  {32'h40353528, 32'h3c226300} /* (6, 28, 27) {real, imag} */,
  {32'h3fb89bf8, 32'hbf8325d7} /* (6, 28, 26) {real, imag} */,
  {32'hbeffb00c, 32'hbd81d240} /* (6, 28, 25) {real, imag} */,
  {32'h402c20b6, 32'h3f48f1d0} /* (6, 28, 24) {real, imag} */,
  {32'h3fad650c, 32'hbc544f80} /* (6, 28, 23) {real, imag} */,
  {32'h3ff21cd8, 32'h3f95ed7f} /* (6, 28, 22) {real, imag} */,
  {32'h3fb512ba, 32'hbeec4af2} /* (6, 28, 21) {real, imag} */,
  {32'hc054925c, 32'h3f149c81} /* (6, 28, 20) {real, imag} */,
  {32'hc0271f66, 32'hbd296000} /* (6, 28, 19) {real, imag} */,
  {32'hbe0bbfcc, 32'h3f83d3b4} /* (6, 28, 18) {real, imag} */,
  {32'hbf2130cd, 32'h3f8bbff5} /* (6, 28, 17) {real, imag} */,
  {32'hc00da723, 32'hc019e9f2} /* (6, 28, 16) {real, imag} */,
  {32'h3d0c3340, 32'hc0353e62} /* (6, 28, 15) {real, imag} */,
  {32'h401fc758, 32'hbf1a58d2} /* (6, 28, 14) {real, imag} */,
  {32'h401f99cc, 32'h3f47259e} /* (6, 28, 13) {real, imag} */,
  {32'h3f494c2a, 32'h400142c0} /* (6, 28, 12) {real, imag} */,
  {32'h400e0966, 32'h3f4283d1} /* (6, 28, 11) {real, imag} */,
  {32'h4021f100, 32'h3f9ab006} /* (6, 28, 10) {real, imag} */,
  {32'hbee0487c, 32'hbfc29abe} /* (6, 28, 9) {real, imag} */,
  {32'hbf9c4bfa, 32'hbf4f6a7c} /* (6, 28, 8) {real, imag} */,
  {32'hbe424c50, 32'hbf23bbfa} /* (6, 28, 7) {real, imag} */,
  {32'hbf48184c, 32'hbf12922e} /* (6, 28, 6) {real, imag} */,
  {32'hbf5aa14f, 32'hbf44abe0} /* (6, 28, 5) {real, imag} */,
  {32'h3f4d9178, 32'hbf875932} /* (6, 28, 4) {real, imag} */,
  {32'h3f547080, 32'hbf55adc2} /* (6, 28, 3) {real, imag} */,
  {32'h3eec14a6, 32'hbf2366cc} /* (6, 28, 2) {real, imag} */,
  {32'h3f79ae2f, 32'h3e85034e} /* (6, 28, 1) {real, imag} */,
  {32'h3f07555a, 32'h3f3fd885} /* (6, 28, 0) {real, imag} */,
  {32'hbeb6c85e, 32'h3f301fb5} /* (6, 27, 31) {real, imag} */,
  {32'hbfaabd13, 32'h3f38880c} /* (6, 27, 30) {real, imag} */,
  {32'hbf4e94ad, 32'hbff33082} /* (6, 27, 29) {real, imag} */,
  {32'hbfb41334, 32'hc07a471c} /* (6, 27, 28) {real, imag} */,
  {32'h3e9fef52, 32'hbf475cea} /* (6, 27, 27) {real, imag} */,
  {32'h405f5621, 32'h3ffa907d} /* (6, 27, 26) {real, imag} */,
  {32'h3fe22904, 32'h401513ef} /* (6, 27, 25) {real, imag} */,
  {32'hbed6bff8, 32'hc004c36b} /* (6, 27, 24) {real, imag} */,
  {32'h3f7ad5b4, 32'hbf669c92} /* (6, 27, 23) {real, imag} */,
  {32'h3f55707d, 32'hbf1252bf} /* (6, 27, 22) {real, imag} */,
  {32'h3f7c7c10, 32'hbf11a9c5} /* (6, 27, 21) {real, imag} */,
  {32'hbfb3d9ba, 32'hbeafd170} /* (6, 27, 20) {real, imag} */,
  {32'hc02ead05, 32'h3f0cf096} /* (6, 27, 19) {real, imag} */,
  {32'hc0069107, 32'h3fd4735c} /* (6, 27, 18) {real, imag} */,
  {32'hc017aa0b, 32'hbf8b8f7d} /* (6, 27, 17) {real, imag} */,
  {32'hc001465e, 32'hbf641c35} /* (6, 27, 16) {real, imag} */,
  {32'h3dff66d0, 32'h3f7d95e2} /* (6, 27, 15) {real, imag} */,
  {32'h3f1a650e, 32'hbf54379a} /* (6, 27, 14) {real, imag} */,
  {32'h3f07fe3e, 32'hbfa06012} /* (6, 27, 13) {real, imag} */,
  {32'hbd8ec9c8, 32'h40034e2e} /* (6, 27, 12) {real, imag} */,
  {32'h3fffd3f0, 32'h3eb263aa} /* (6, 27, 11) {real, imag} */,
  {32'h3fd0ea1a, 32'h3f056220} /* (6, 27, 10) {real, imag} */,
  {32'hbfe3aed1, 32'hbfd2a02c} /* (6, 27, 9) {real, imag} */,
  {32'hc05cd75c, 32'hbf68dd14} /* (6, 27, 8) {real, imag} */,
  {32'hc03ab422, 32'h3eead05c} /* (6, 27, 7) {real, imag} */,
  {32'hbebc3016, 32'hbe404138} /* (6, 27, 6) {real, imag} */,
  {32'h3f7be7f8, 32'h3f0a1d35} /* (6, 27, 5) {real, imag} */,
  {32'h3f196656, 32'h3f494bec} /* (6, 27, 4) {real, imag} */,
  {32'h3f035b5b, 32'h3e1c2038} /* (6, 27, 3) {real, imag} */,
  {32'h3f4efadc, 32'h3fb15e8c} /* (6, 27, 2) {real, imag} */,
  {32'h3efd4e2c, 32'hbf2680a6} /* (6, 27, 1) {real, imag} */,
  {32'hbf97c180, 32'hbf8c0d30} /* (6, 27, 0) {real, imag} */,
  {32'hbeecd59e, 32'hbed393fa} /* (6, 26, 31) {real, imag} */,
  {32'hbfb8c3cb, 32'hbe11917c} /* (6, 26, 30) {real, imag} */,
  {32'hbf951d1a, 32'hbfccc106} /* (6, 26, 29) {real, imag} */,
  {32'hbfacd871, 32'hc01f294d} /* (6, 26, 28) {real, imag} */,
  {32'hbcbe0438, 32'hbfaaf29c} /* (6, 26, 27) {real, imag} */,
  {32'h3f959911, 32'h3e88808c} /* (6, 26, 26) {real, imag} */,
  {32'h3f19eafe, 32'h3efb783c} /* (6, 26, 25) {real, imag} */,
  {32'hbff87bb2, 32'hbfcc83d4} /* (6, 26, 24) {real, imag} */,
  {32'hbe942e72, 32'hbff5789d} /* (6, 26, 23) {real, imag} */,
  {32'h3c2db580, 32'hbfaaf530} /* (6, 26, 22) {real, imag} */,
  {32'hbede3b16, 32'hbf285add} /* (6, 26, 21) {real, imag} */,
  {32'hbeb7c714, 32'hbece062e} /* (6, 26, 20) {real, imag} */,
  {32'hbd5e17c0, 32'h3e0a2e58} /* (6, 26, 19) {real, imag} */,
  {32'hbfd35895, 32'h4019f8a4} /* (6, 26, 18) {real, imag} */,
  {32'hc03db6dc, 32'hbf503bf5} /* (6, 26, 17) {real, imag} */,
  {32'hbe9efa02, 32'hbea8f856} /* (6, 26, 16) {real, imag} */,
  {32'hbf3d5a35, 32'h404fc2d0} /* (6, 26, 15) {real, imag} */,
  {32'hbf3e2c50, 32'h3fca7dbf} /* (6, 26, 14) {real, imag} */,
  {32'hbe95a5f0, 32'h3e9e30e4} /* (6, 26, 13) {real, imag} */,
  {32'hbf2d6318, 32'h3eab90b6} /* (6, 26, 12) {real, imag} */,
  {32'h3f1e326e, 32'hbf47ee6d} /* (6, 26, 11) {real, imag} */,
  {32'hbf8ef085, 32'hbf443e3b} /* (6, 26, 10) {real, imag} */,
  {32'hbfe18672, 32'hbfcec66b} /* (6, 26, 9) {real, imag} */,
  {32'hbf9aee5c, 32'hc0130914} /* (6, 26, 8) {real, imag} */,
  {32'hbfde002b, 32'h3f96eddb} /* (6, 26, 7) {real, imag} */,
  {32'hbfd06acc, 32'h40353361} /* (6, 26, 6) {real, imag} */,
  {32'h3f4d0a98, 32'h3f9dee2a} /* (6, 26, 5) {real, imag} */,
  {32'hbfb488f8, 32'h4009c9ab} /* (6, 26, 4) {real, imag} */,
  {32'hc007bd18, 32'h40782adc} /* (6, 26, 3) {real, imag} */,
  {32'hbf34919a, 32'h408d2880} /* (6, 26, 2) {real, imag} */,
  {32'hbf94e038, 32'h3f6e6828} /* (6, 26, 1) {real, imag} */,
  {32'hbf95d82c, 32'hbf1e956e} /* (6, 26, 0) {real, imag} */,
  {32'hbfb9cd65, 32'hbf8dc7e8} /* (6, 25, 31) {real, imag} */,
  {32'hc009b8ce, 32'hbef28876} /* (6, 25, 30) {real, imag} */,
  {32'hbfc09ebe, 32'hbeec9cc6} /* (6, 25, 29) {real, imag} */,
  {32'hbf40a07c, 32'hbfa9519c} /* (6, 25, 28) {real, imag} */,
  {32'h3f4e0d22, 32'hc01ba548} /* (6, 25, 27) {real, imag} */,
  {32'h3ef6ba7e, 32'hbff6ce00} /* (6, 25, 26) {real, imag} */,
  {32'h3dc5b4e0, 32'hc00855cf} /* (6, 25, 25) {real, imag} */,
  {32'hbfc2662a, 32'hbf752d1c} /* (6, 25, 24) {real, imag} */,
  {32'hbf4407aa, 32'hbfc1059c} /* (6, 25, 23) {real, imag} */,
  {32'hbf8bad89, 32'hc01aace2} /* (6, 25, 22) {real, imag} */,
  {32'hbfe1cf11, 32'hbf8767b0} /* (6, 25, 21) {real, imag} */,
  {32'h3e90302c, 32'hbf311826} /* (6, 25, 20) {real, imag} */,
  {32'h400c355c, 32'hc003175f} /* (6, 25, 19) {real, imag} */,
  {32'hbe5830e0, 32'h3f3e8776} /* (6, 25, 18) {real, imag} */,
  {32'hc022e036, 32'hbf303456} /* (6, 25, 17) {real, imag} */,
  {32'h3ff8d0db, 32'hbf808a14} /* (6, 25, 16) {real, imag} */,
  {32'h3ffec784, 32'h3ed40a5a} /* (6, 25, 15) {real, imag} */,
  {32'h3fdd8fa8, 32'h3f50b738} /* (6, 25, 14) {real, imag} */,
  {32'h403b6078, 32'h3f5b8e02} /* (6, 25, 13) {real, imag} */,
  {32'h3e32b5a0, 32'h3dec4f70} /* (6, 25, 12) {real, imag} */,
  {32'h3f562d46, 32'h3de22590} /* (6, 25, 11) {real, imag} */,
  {32'hbf88a8da, 32'h3fca1418} /* (6, 25, 10) {real, imag} */,
  {32'hbff1ecc7, 32'h3d38ee20} /* (6, 25, 9) {real, imag} */,
  {32'h3f599ccc, 32'hc0263375} /* (6, 25, 8) {real, imag} */,
  {32'h3fc607e9, 32'h3f8587d1} /* (6, 25, 7) {real, imag} */,
  {32'h3e386414, 32'h4034b730} /* (6, 25, 6) {real, imag} */,
  {32'h3e05b464, 32'h40198208} /* (6, 25, 5) {real, imag} */,
  {32'hbfa5c849, 32'h40170fde} /* (6, 25, 4) {real, imag} */,
  {32'hc00b0613, 32'h405ba6cc} /* (6, 25, 3) {real, imag} */,
  {32'hbf396e18, 32'h3fac6e7b} /* (6, 25, 2) {real, imag} */,
  {32'hbf24bed2, 32'h4020a5d9} /* (6, 25, 1) {real, imag} */,
  {32'hbf27ac52, 32'h3f0d140c} /* (6, 25, 0) {real, imag} */,
  {32'hbfcf9ba5, 32'h3fb2cd24} /* (6, 24, 31) {real, imag} */,
  {32'hbe454338, 32'h3fdff0a9} /* (6, 24, 30) {real, imag} */,
  {32'h3f90c89d, 32'h3f8fdb06} /* (6, 24, 29) {real, imag} */,
  {32'h3f9f0c6e, 32'h3e1f3058} /* (6, 24, 28) {real, imag} */,
  {32'h3fc7b9c9, 32'hbfce0003} /* (6, 24, 27) {real, imag} */,
  {32'hbf1a2a10, 32'hc0007ffa} /* (6, 24, 26) {real, imag} */,
  {32'h3da91e28, 32'hc0985f9f} /* (6, 24, 25) {real, imag} */,
  {32'hbc47a840, 32'hc02f0b02} /* (6, 24, 24) {real, imag} */,
  {32'h3f8af200, 32'hbfdb4228} /* (6, 24, 23) {real, imag} */,
  {32'hbfdcb314, 32'hbf07884e} /* (6, 24, 22) {real, imag} */,
  {32'hbffd7104, 32'hbff4c4e4} /* (6, 24, 21) {real, imag} */,
  {32'hbe0d1118, 32'hbfd27bd8} /* (6, 24, 20) {real, imag} */,
  {32'h3ff86ad9, 32'hbf3e9734} /* (6, 24, 19) {real, imag} */,
  {32'h3f8306e7, 32'h3fc41db6} /* (6, 24, 18) {real, imag} */,
  {32'hbfaf3526, 32'hbf271a52} /* (6, 24, 17) {real, imag} */,
  {32'h40193f26, 32'h3efad2d4} /* (6, 24, 16) {real, imag} */,
  {32'h3ffa5fbc, 32'h402f2ad3} /* (6, 24, 15) {real, imag} */,
  {32'h3fc5b277, 32'h404121c9} /* (6, 24, 14) {real, imag} */,
  {32'h40d16606, 32'h3fade0ef} /* (6, 24, 13) {real, imag} */,
  {32'h40205827, 32'hbec283d4} /* (6, 24, 12) {real, imag} */,
  {32'h4002050f, 32'h3dd0c5e8} /* (6, 24, 11) {real, imag} */,
  {32'h3ffb290d, 32'h404cdd32} /* (6, 24, 10) {real, imag} */,
  {32'h3e55cb10, 32'hbea9052c} /* (6, 24, 9) {real, imag} */,
  {32'h3e6b4fa8, 32'hbfa9ebb8} /* (6, 24, 8) {real, imag} */,
  {32'h3f22dae7, 32'h40001fee} /* (6, 24, 7) {real, imag} */,
  {32'hbeb8b406, 32'h3eadf734} /* (6, 24, 6) {real, imag} */,
  {32'hbfbe590b, 32'h3f89d837} /* (6, 24, 5) {real, imag} */,
  {32'hbfa841a4, 32'h3f0716b7} /* (6, 24, 4) {real, imag} */,
  {32'hbf0af1a1, 32'h3fdb0f1b} /* (6, 24, 3) {real, imag} */,
  {32'hbf01fc54, 32'h3e8aaa18} /* (6, 24, 2) {real, imag} */,
  {32'h3f41c800, 32'h3e393eec} /* (6, 24, 1) {real, imag} */,
  {32'h3f16de4c, 32'hbe88d377} /* (6, 24, 0) {real, imag} */,
  {32'hbf1df689, 32'hbdac3240} /* (6, 23, 31) {real, imag} */,
  {32'hbdbdc5f0, 32'hbf314bb4} /* (6, 23, 30) {real, imag} */,
  {32'h3f37343a, 32'h3d8235f8} /* (6, 23, 29) {real, imag} */,
  {32'h3e574540, 32'hbe074c20} /* (6, 23, 28) {real, imag} */,
  {32'h3fedd428, 32'hc057e526} /* (6, 23, 27) {real, imag} */,
  {32'hbea8ab64, 32'hc05dd35a} /* (6, 23, 26) {real, imag} */,
  {32'h3f3d401e, 32'hc06076b1} /* (6, 23, 25) {real, imag} */,
  {32'h400754e7, 32'hc04fc388} /* (6, 23, 24) {real, imag} */,
  {32'h3dd3f3e0, 32'hc02292a9} /* (6, 23, 23) {real, imag} */,
  {32'h3ef9d2e4, 32'hbfeb2d86} /* (6, 23, 22) {real, imag} */,
  {32'h3eedaea3, 32'hc00bbbda} /* (6, 23, 21) {real, imag} */,
  {32'h3e81871c, 32'hbfa402f7} /* (6, 23, 20) {real, imag} */,
  {32'hbfc57397, 32'hbc3b9880} /* (6, 23, 19) {real, imag} */,
  {32'hbfc39a53, 32'h3f8fd005} /* (6, 23, 18) {real, imag} */,
  {32'hc0417b1e, 32'hbfcd107a} /* (6, 23, 17) {real, imag} */,
  {32'h3f43f8af, 32'hbd3ad480} /* (6, 23, 16) {real, imag} */,
  {32'h3fbc575e, 32'h4025ff94} /* (6, 23, 15) {real, imag} */,
  {32'hbec55bae, 32'h4046c4b2} /* (6, 23, 14) {real, imag} */,
  {32'h406f73be, 32'h3f6c20b6} /* (6, 23, 13) {real, imag} */,
  {32'h3fac416d, 32'hbf06cc0e} /* (6, 23, 12) {real, imag} */,
  {32'h3f1a5811, 32'hbf287798} /* (6, 23, 11) {real, imag} */,
  {32'h403c80e3, 32'h3f31b7fd} /* (6, 23, 10) {real, imag} */,
  {32'h40001812, 32'hbef6965c} /* (6, 23, 9) {real, imag} */,
  {32'hbdf488f8, 32'h3d458a70} /* (6, 23, 8) {real, imag} */,
  {32'hbe4ca6c4, 32'h3fa2f991} /* (6, 23, 7) {real, imag} */,
  {32'hbf2b9986, 32'hbfc8d5a3} /* (6, 23, 6) {real, imag} */,
  {32'hc0370b69, 32'hbf646f2b} /* (6, 23, 5) {real, imag} */,
  {32'hbfe1fcf0, 32'h3e4aacd8} /* (6, 23, 4) {real, imag} */,
  {32'hbf0928a8, 32'h3ef7eb2c} /* (6, 23, 3) {real, imag} */,
  {32'h3e8d02dc, 32'h3f8ca284} /* (6, 23, 2) {real, imag} */,
  {32'h3ff5578a, 32'hbe5b8d90} /* (6, 23, 1) {real, imag} */,
  {32'h3f84aabd, 32'hbdd380a8} /* (6, 23, 0) {real, imag} */,
  {32'h3dae3c20, 32'hbdcc81d8} /* (6, 22, 31) {real, imag} */,
  {32'h3f6a6249, 32'hbfd7dd47} /* (6, 22, 30) {real, imag} */,
  {32'h3f230010, 32'hbfa6f478} /* (6, 22, 29) {real, imag} */,
  {32'h3fc4a038, 32'hbf629200} /* (6, 22, 28) {real, imag} */,
  {32'h40443c77, 32'hc0430430} /* (6, 22, 27) {real, imag} */,
  {32'h4008bd74, 32'hc05a11a8} /* (6, 22, 26) {real, imag} */,
  {32'hbf11738e, 32'hbfeda1e2} /* (6, 22, 25) {real, imag} */,
  {32'hbf48f87a, 32'hc000ab6d} /* (6, 22, 24) {real, imag} */,
  {32'hbfa97b06, 32'hbfc4b56e} /* (6, 22, 23) {real, imag} */,
  {32'hbf8e7dba, 32'hbdccb568} /* (6, 22, 22) {real, imag} */,
  {32'hbf588a53, 32'h3fe47342} /* (6, 22, 21) {real, imag} */,
  {32'hbdef8408, 32'h3f200846} /* (6, 22, 20) {real, imag} */,
  {32'hc02b0ff6, 32'hbe840f00} /* (6, 22, 19) {real, imag} */,
  {32'hbfea38ca, 32'hbd60f7c0} /* (6, 22, 18) {real, imag} */,
  {32'hc03762ed, 32'hbfd620b2} /* (6, 22, 17) {real, imag} */,
  {32'hbfe7ad64, 32'hc0054b13} /* (6, 22, 16) {real, imag} */,
  {32'h3ec17f0a, 32'hbeb6a20e} /* (6, 22, 15) {real, imag} */,
  {32'hbfebda4a, 32'h3f49cd8a} /* (6, 22, 14) {real, imag} */,
  {32'hbf1385fc, 32'h3ff75a70} /* (6, 22, 13) {real, imag} */,
  {32'h3f71abcb, 32'h4024288b} /* (6, 22, 12) {real, imag} */,
  {32'h4007d7f7, 32'h3fd92914} /* (6, 22, 11) {real, imag} */,
  {32'h4011036f, 32'h3df4a598} /* (6, 22, 10) {real, imag} */,
  {32'h4023808f, 32'hc0106c78} /* (6, 22, 9) {real, imag} */,
  {32'h3fb9324e, 32'hbf85c4e7} /* (6, 22, 8) {real, imag} */,
  {32'h3ef3b7ca, 32'hc01a64be} /* (6, 22, 7) {real, imag} */,
  {32'h3cbcac00, 32'hbfca8354} /* (6, 22, 6) {real, imag} */,
  {32'hbfdb9ed0, 32'h3e837190} /* (6, 22, 5) {real, imag} */,
  {32'hc0038781, 32'h3f563c82} /* (6, 22, 4) {real, imag} */,
  {32'hbf8b32f9, 32'hbed01a70} /* (6, 22, 3) {real, imag} */,
  {32'hbecb4b40, 32'h3f9e7de6} /* (6, 22, 2) {real, imag} */,
  {32'h3fa8660a, 32'hbf7690e4} /* (6, 22, 1) {real, imag} */,
  {32'h4028fbf2, 32'h3e55db0c} /* (6, 22, 0) {real, imag} */,
  {32'hbed10dbe, 32'h3f9e27bf} /* (6, 21, 31) {real, imag} */,
  {32'h3f9158ad, 32'h3fdf7204} /* (6, 21, 30) {real, imag} */,
  {32'h3fb4f2fe, 32'hbf82e369} /* (6, 21, 29) {real, imag} */,
  {32'h4005528c, 32'hbfb3dc84} /* (6, 21, 28) {real, imag} */,
  {32'h40249ea5, 32'hbfe5d972} /* (6, 21, 27) {real, imag} */,
  {32'h3fe4b485, 32'hc018d902} /* (6, 21, 26) {real, imag} */,
  {32'hbf07080e, 32'hbf892300} /* (6, 21, 25) {real, imag} */,
  {32'hbf6af5fe, 32'hbf1a0f90} /* (6, 21, 24) {real, imag} */,
  {32'hbf44e6bc, 32'h3f19ff8c} /* (6, 21, 23) {real, imag} */,
  {32'hbf2d8fef, 32'h405f51fc} /* (6, 21, 22) {real, imag} */,
  {32'hbdc60c30, 32'h40a7cd40} /* (6, 21, 21) {real, imag} */,
  {32'h3ef10fa4, 32'h3f006d5e} /* (6, 21, 20) {real, imag} */,
  {32'h3fc3870f, 32'hbfe5964a} /* (6, 21, 19) {real, imag} */,
  {32'h3e1ddbc4, 32'hc0139316} /* (6, 21, 18) {real, imag} */,
  {32'hc00f1a82, 32'hbf9af7b1} /* (6, 21, 17) {real, imag} */,
  {32'hc031540e, 32'hbee4b87e} /* (6, 21, 16) {real, imag} */,
  {32'h3fbab2bc, 32'h3ed996a8} /* (6, 21, 15) {real, imag} */,
  {32'h3cb1fe00, 32'h3f257cad} /* (6, 21, 14) {real, imag} */,
  {32'hbff9ad44, 32'h3ede5cd2} /* (6, 21, 13) {real, imag} */,
  {32'hbed53cc0, 32'h3f539673} /* (6, 21, 12) {real, imag} */,
  {32'h3fba3935, 32'h3f41eba1} /* (6, 21, 11) {real, imag} */,
  {32'h3f3ea733, 32'hbfd39faa} /* (6, 21, 10) {real, imag} */,
  {32'h3f48cc38, 32'hc028ae4b} /* (6, 21, 9) {real, imag} */,
  {32'h3e120d50, 32'hbf974da3} /* (6, 21, 8) {real, imag} */,
  {32'hbf1b665a, 32'hbfc311f5} /* (6, 21, 7) {real, imag} */,
  {32'h3ffd53fe, 32'h3f6010d2} /* (6, 21, 6) {real, imag} */,
  {32'h3fadc4b6, 32'h4010cb4d} /* (6, 21, 5) {real, imag} */,
  {32'h3f88094f, 32'h3fff2021} /* (6, 21, 4) {real, imag} */,
  {32'h3f4ea6fd, 32'h3f04f016} /* (6, 21, 3) {real, imag} */,
  {32'h3ec7494c, 32'h40057e97} /* (6, 21, 2) {real, imag} */,
  {32'hbf1aecbc, 32'h3e5f7a4c} /* (6, 21, 1) {real, imag} */,
  {32'hbd47a920, 32'h3f2b3498} /* (6, 21, 0) {real, imag} */,
  {32'h3df9f644, 32'h3fd0a96e} /* (6, 20, 31) {real, imag} */,
  {32'h3ff202c7, 32'h400b1c16} /* (6, 20, 30) {real, imag} */,
  {32'h4015ae20, 32'h3f2624b8} /* (6, 20, 29) {real, imag} */,
  {32'h3f93e160, 32'h3f93d694} /* (6, 20, 28) {real, imag} */,
  {32'h3ed04264, 32'h3eb522d8} /* (6, 20, 27) {real, imag} */,
  {32'h3e0c82c4, 32'hbf506de6} /* (6, 20, 26) {real, imag} */,
  {32'hbf859dfd, 32'hbf1685d3} /* (6, 20, 25) {real, imag} */,
  {32'hbe1622a8, 32'hbfa616eb} /* (6, 20, 24) {real, imag} */,
  {32'hbfac9548, 32'h3fea805a} /* (6, 20, 23) {real, imag} */,
  {32'hbf6756c4, 32'h40755e80} /* (6, 20, 22) {real, imag} */,
  {32'h3ed9d2f2, 32'h40451008} /* (6, 20, 21) {real, imag} */,
  {32'h3fb90996, 32'h3f814171} /* (6, 20, 20) {real, imag} */,
  {32'h3fb9002c, 32'hbffd31c7} /* (6, 20, 19) {real, imag} */,
  {32'hbcd88128, 32'hc074a9b9} /* (6, 20, 18) {real, imag} */,
  {32'hc007ea2a, 32'hc02f2f82} /* (6, 20, 17) {real, imag} */,
  {32'h3c44ca20, 32'h3f6a60c0} /* (6, 20, 16) {real, imag} */,
  {32'h40286915, 32'hbdf96810} /* (6, 20, 15) {real, imag} */,
  {32'h3f88c29f, 32'hbe87e1ee} /* (6, 20, 14) {real, imag} */,
  {32'hbfa80fb0, 32'h3f438213} /* (6, 20, 13) {real, imag} */,
  {32'h3f12068a, 32'hbc2bd6c0} /* (6, 20, 12) {real, imag} */,
  {32'h3f01d76e, 32'h3f57eab2} /* (6, 20, 11) {real, imag} */,
  {32'hbf91a355, 32'h3f9092ff} /* (6, 20, 10) {real, imag} */,
  {32'h3f8f8344, 32'hbf28b93e} /* (6, 20, 9) {real, imag} */,
  {32'h3fb4f664, 32'hbf93cb3f} /* (6, 20, 8) {real, imag} */,
  {32'h3eaeec4c, 32'hbfcf5328} /* (6, 20, 7) {real, imag} */,
  {32'h4002c7fa, 32'h3e3cdfd0} /* (6, 20, 6) {real, imag} */,
  {32'h3f9b853e, 32'h3fd994f0} /* (6, 20, 5) {real, imag} */,
  {32'h402e3532, 32'h3e79cc90} /* (6, 20, 4) {real, imag} */,
  {32'h40381cae, 32'hbf4515e3} /* (6, 20, 3) {real, imag} */,
  {32'h3ff62b0a, 32'h3fe15cbc} /* (6, 20, 2) {real, imag} */,
  {32'hbf8d692d, 32'h3f5e750a} /* (6, 20, 1) {real, imag} */,
  {32'hbfc4a533, 32'hbe6713b3} /* (6, 20, 0) {real, imag} */,
  {32'hbdbda960, 32'hbdcbc080} /* (6, 19, 31) {real, imag} */,
  {32'hbdc01418, 32'h3f346124} /* (6, 19, 30) {real, imag} */,
  {32'h3f1a4bba, 32'h3f9cc31e} /* (6, 19, 29) {real, imag} */,
  {32'hbf3d13b9, 32'h3febf3a6} /* (6, 19, 28) {real, imag} */,
  {32'hbf3c507d, 32'hbe7ede70} /* (6, 19, 27) {real, imag} */,
  {32'hbf1cee66, 32'h3f18681b} /* (6, 19, 26) {real, imag} */,
  {32'hc057da16, 32'h3e9c9db4} /* (6, 19, 25) {real, imag} */,
  {32'hc083b8b2, 32'hbe0c0bd8} /* (6, 19, 24) {real, imag} */,
  {32'hbe08f4e8, 32'h3f08ed3a} /* (6, 19, 23) {real, imag} */,
  {32'h3ef8bd92, 32'h3f2faae2} /* (6, 19, 22) {real, imag} */,
  {32'h3e98648e, 32'h3f0a85d7} /* (6, 19, 21) {real, imag} */,
  {32'h3fc89290, 32'hbfaf6505} /* (6, 19, 20) {real, imag} */,
  {32'hbde60300, 32'hbfd81ac8} /* (6, 19, 19) {real, imag} */,
  {32'h3ee4d21c, 32'hc0256536} /* (6, 19, 18) {real, imag} */,
  {32'h3d587a70, 32'hc0886b42} /* (6, 19, 17) {real, imag} */,
  {32'hbd7b75e0, 32'hbf43cca7} /* (6, 19, 16) {real, imag} */,
  {32'h3f5997e4, 32'hbfb1cfe4} /* (6, 19, 15) {real, imag} */,
  {32'hc0042d35, 32'hbe2aaa00} /* (6, 19, 14) {real, imag} */,
  {32'hc010c0a1, 32'h3fe893be} /* (6, 19, 13) {real, imag} */,
  {32'hbe7eb91c, 32'h4008ad50} /* (6, 19, 12) {real, imag} */,
  {32'hbfa7b388, 32'h40508f39} /* (6, 19, 11) {real, imag} */,
  {32'hbf8de790, 32'h40644528} /* (6, 19, 10) {real, imag} */,
  {32'h40177949, 32'h3ee6f1e8} /* (6, 19, 9) {real, imag} */,
  {32'h401465a3, 32'hbff51f78} /* (6, 19, 8) {real, imag} */,
  {32'h3fdfe1f5, 32'hc06cbf86} /* (6, 19, 7) {real, imag} */,
  {32'h402bb444, 32'hc038e3e4} /* (6, 19, 6) {real, imag} */,
  {32'h3ea9017e, 32'h3dd51a80} /* (6, 19, 5) {real, imag} */,
  {32'h3e87f780, 32'hbffdb377} /* (6, 19, 4) {real, imag} */,
  {32'h4010cbd5, 32'hc046a437} /* (6, 19, 3) {real, imag} */,
  {32'h3f8d4f6f, 32'h3e11fc78} /* (6, 19, 2) {real, imag} */,
  {32'hbe326df8, 32'h3e7b6170} /* (6, 19, 1) {real, imag} */,
  {32'hbfb28940, 32'h3ed6681a} /* (6, 19, 0) {real, imag} */,
  {32'h3f723f73, 32'hbf65ea5e} /* (6, 18, 31) {real, imag} */,
  {32'hbf7214c4, 32'hbe517aa0} /* (6, 18, 30) {real, imag} */,
  {32'hbf0507ee, 32'h3fbba18a} /* (6, 18, 29) {real, imag} */,
  {32'hbf8d6f09, 32'h3f86fa5c} /* (6, 18, 28) {real, imag} */,
  {32'h3f4875e6, 32'h3f9cb64e} /* (6, 18, 27) {real, imag} */,
  {32'h3f8c30e5, 32'h4019d864} /* (6, 18, 26) {real, imag} */,
  {32'hc01e5736, 32'h3fbacb79} /* (6, 18, 25) {real, imag} */,
  {32'hbfc906d8, 32'h404168cb} /* (6, 18, 24) {real, imag} */,
  {32'h40261ec0, 32'h3fccd071} /* (6, 18, 23) {real, imag} */,
  {32'h3f04fe0a, 32'h3ff1e895} /* (6, 18, 22) {real, imag} */,
  {32'hbf4875cf, 32'h408095ce} /* (6, 18, 21) {real, imag} */,
  {32'h400dabd0, 32'h40033dd7} /* (6, 18, 20) {real, imag} */,
  {32'hbd575fb0, 32'h3fe7c308} /* (6, 18, 19) {real, imag} */,
  {32'h3e8081c3, 32'hbf6fa56f} /* (6, 18, 18) {real, imag} */,
  {32'h3f1e88fe, 32'hc060d21c} /* (6, 18, 17) {real, imag} */,
  {32'hc01ab4ea, 32'hc014bc3e} /* (6, 18, 16) {real, imag} */,
  {32'hbea2eff0, 32'hbffdc744} /* (6, 18, 15) {real, imag} */,
  {32'hbfa80ca8, 32'hbfb32e29} /* (6, 18, 14) {real, imag} */,
  {32'hbf71686a, 32'h3f541f1a} /* (6, 18, 13) {real, imag} */,
  {32'h3edc7be6, 32'h404d6b8e} /* (6, 18, 12) {real, imag} */,
  {32'h3e5adc18, 32'h40597d3c} /* (6, 18, 11) {real, imag} */,
  {32'h3ea8b47a, 32'h3e6293b8} /* (6, 18, 10) {real, imag} */,
  {32'h3f9fc2d0, 32'hbffd3e8a} /* (6, 18, 9) {real, imag} */,
  {32'h3f1bf54c, 32'hc0456718} /* (6, 18, 8) {real, imag} */,
  {32'hbf82d8d0, 32'hc0852c60} /* (6, 18, 7) {real, imag} */,
  {32'h3f7c5894, 32'hbed022c0} /* (6, 18, 6) {real, imag} */,
  {32'h3fa0479e, 32'h4037ed97} /* (6, 18, 5) {real, imag} */,
  {32'h3fe81c7a, 32'h3feaa674} /* (6, 18, 4) {real, imag} */,
  {32'h4026e9ac, 32'hbb82b200} /* (6, 18, 3) {real, imag} */,
  {32'h400fbf03, 32'h3ee00da6} /* (6, 18, 2) {real, imag} */,
  {32'h40688041, 32'hbe730350} /* (6, 18, 1) {real, imag} */,
  {32'h3f42e974, 32'h3d446fa0} /* (6, 18, 0) {real, imag} */,
  {32'h3fc2240c, 32'hc0102ae7} /* (6, 17, 31) {real, imag} */,
  {32'h400c5854, 32'hbeeca2e8} /* (6, 17, 30) {real, imag} */,
  {32'h3f3f7755, 32'h3fc085b0} /* (6, 17, 29) {real, imag} */,
  {32'h3f470846, 32'h3fe61771} /* (6, 17, 28) {real, imag} */,
  {32'h3f30f11e, 32'h40347fb7} /* (6, 17, 27) {real, imag} */,
  {32'h3faa0660, 32'h40873c6b} /* (6, 17, 26) {real, imag} */,
  {32'h3f520e4e, 32'h4028688c} /* (6, 17, 25) {real, imag} */,
  {32'h403922a3, 32'h4021927a} /* (6, 17, 24) {real, imag} */,
  {32'h402a8c96, 32'h3f34eb88} /* (6, 17, 23) {real, imag} */,
  {32'h3fc0e128, 32'hbe8f4d1e} /* (6, 17, 22) {real, imag} */,
  {32'hbe7845d4, 32'h400f4b70} /* (6, 17, 21) {real, imag} */,
  {32'h3ff62f60, 32'h404953f4} /* (6, 17, 20) {real, imag} */,
  {32'h3f55183a, 32'h4009da60} /* (6, 17, 19) {real, imag} */,
  {32'h3f2b530c, 32'h3fc0023a} /* (6, 17, 18) {real, imag} */,
  {32'h3f31b71a, 32'h3f75c74e} /* (6, 17, 17) {real, imag} */,
  {32'h3f3bbf84, 32'hbfc1ecec} /* (6, 17, 16) {real, imag} */,
  {32'h3f3e83ec, 32'hc037edf3} /* (6, 17, 15) {real, imag} */,
  {32'h3f55d8e6, 32'hbffe83e2} /* (6, 17, 14) {real, imag} */,
  {32'h3e97f5ee, 32'h3e049674} /* (6, 17, 13) {real, imag} */,
  {32'h3ed55ab0, 32'h3fea6098} /* (6, 17, 12) {real, imag} */,
  {32'h3f8aa296, 32'h3f84e4fc} /* (6, 17, 11) {real, imag} */,
  {32'h3fb20069, 32'hc0232005} /* (6, 17, 10) {real, imag} */,
  {32'h400078c0, 32'hc0a32772} /* (6, 17, 9) {real, imag} */,
  {32'h4056ec0b, 32'hc06cb6d9} /* (6, 17, 8) {real, imag} */,
  {32'hbde8ddd0, 32'hbe106e20} /* (6, 17, 7) {real, imag} */,
  {32'hbefbf430, 32'hbd34b8e0} /* (6, 17, 6) {real, imag} */,
  {32'h3fc4cb26, 32'h3fb2df84} /* (6, 17, 5) {real, imag} */,
  {32'h3fcfd877, 32'h4086b098} /* (6, 17, 4) {real, imag} */,
  {32'h3f2e46c4, 32'h40743790} /* (6, 17, 3) {real, imag} */,
  {32'h3ecce480, 32'h3f55265a} /* (6, 17, 2) {real, imag} */,
  {32'h4051a6d2, 32'hbf4119b6} /* (6, 17, 1) {real, imag} */,
  {32'h3de14d30, 32'hc00b9a04} /* (6, 17, 0) {real, imag} */,
  {32'hbef15470, 32'hbcd7cc60} /* (6, 16, 31) {real, imag} */,
  {32'h3e2120dc, 32'h3cb90a00} /* (6, 16, 30) {real, imag} */,
  {32'h3eb91d34, 32'h3e289054} /* (6, 16, 29) {real, imag} */,
  {32'h3fdc3677, 32'h40412236} /* (6, 16, 28) {real, imag} */,
  {32'h3f22233e, 32'h3f81f9c8} /* (6, 16, 27) {real, imag} */,
  {32'hbe95fa2c, 32'h3fc3fa93} /* (6, 16, 26) {real, imag} */,
  {32'hbe950a68, 32'h402e5dbf} /* (6, 16, 25) {real, imag} */,
  {32'h3fc42384, 32'h3f3f8d76} /* (6, 16, 24) {real, imag} */,
  {32'h401aeb7a, 32'hbf926868} /* (6, 16, 23) {real, imag} */,
  {32'h4013f1a2, 32'hc00638d2} /* (6, 16, 22) {real, imag} */,
  {32'h3efbe088, 32'h3edc513a} /* (6, 16, 21) {real, imag} */,
  {32'h3fea5019, 32'h3f9d4d94} /* (6, 16, 20) {real, imag} */,
  {32'h3f8fea62, 32'h3fec0b9f} /* (6, 16, 19) {real, imag} */,
  {32'hbe62d538, 32'h401ff778} /* (6, 16, 18) {real, imag} */,
  {32'hbfeb9283, 32'h3f26cc5c} /* (6, 16, 17) {real, imag} */,
  {32'hbe8b2cc8, 32'hbfa8badd} /* (6, 16, 16) {real, imag} */,
  {32'hbf49fa8a, 32'hbffa8579} /* (6, 16, 15) {real, imag} */,
  {32'h3e1c26f8, 32'hbf99db78} /* (6, 16, 14) {real, imag} */,
  {32'h3f5c0ef2, 32'hbeb13ae4} /* (6, 16, 13) {real, imag} */,
  {32'hbed3fe58, 32'h3f855f2b} /* (6, 16, 12) {real, imag} */,
  {32'hbe97423a, 32'hbf9fc6fc} /* (6, 16, 11) {real, imag} */,
  {32'hbf1297e5, 32'hc03454ac} /* (6, 16, 10) {real, imag} */,
  {32'h3e4752c0, 32'hc07d2a15} /* (6, 16, 9) {real, imag} */,
  {32'h3f205c10, 32'hbfd5f677} /* (6, 16, 8) {real, imag} */,
  {32'hbf6ce1a4, 32'h3fd176a6} /* (6, 16, 7) {real, imag} */,
  {32'h3f38048e, 32'h3ffd9283} /* (6, 16, 6) {real, imag} */,
  {32'h3fb8cdec, 32'h3fbe0411} /* (6, 16, 5) {real, imag} */,
  {32'h3e732fe0, 32'h4041aed2} /* (6, 16, 4) {real, imag} */,
  {32'hbfc4b3ca, 32'h402cd37a} /* (6, 16, 3) {real, imag} */,
  {32'hbfd8c784, 32'h3ea719ec} /* (6, 16, 2) {real, imag} */,
  {32'h3ebd0898, 32'h3f8ae200} /* (6, 16, 1) {real, imag} */,
  {32'hbf6b9bb0, 32'h3fdef3bc} /* (6, 16, 0) {real, imag} */,
  {32'hbebb5991, 32'h3f3536a1} /* (6, 15, 31) {real, imag} */,
  {32'h3e3ff114, 32'hbeb0c0b8} /* (6, 15, 30) {real, imag} */,
  {32'h3fdc7953, 32'hbf303ee1} /* (6, 15, 29) {real, imag} */,
  {32'h3f986494, 32'h404de3e4} /* (6, 15, 28) {real, imag} */,
  {32'hbf1e444e, 32'h3e206480} /* (6, 15, 27) {real, imag} */,
  {32'hbfe5ea31, 32'h3e481188} /* (6, 15, 26) {real, imag} */,
  {32'hbfa49401, 32'h4011074a} /* (6, 15, 25) {real, imag} */,
  {32'hbfe1d576, 32'h3fc1b99e} /* (6, 15, 24) {real, imag} */,
  {32'hbd4e5b60, 32'h3fb8b388} /* (6, 15, 23) {real, imag} */,
  {32'hbf0f2f06, 32'h3f100b50} /* (6, 15, 22) {real, imag} */,
  {32'hbecc3416, 32'h3f6d28fe} /* (6, 15, 21) {real, imag} */,
  {32'h3ec890db, 32'hbf15dffe} /* (6, 15, 20) {real, imag} */,
  {32'h3f874163, 32'hbe32c9fc} /* (6, 15, 19) {real, imag} */,
  {32'hbecde4c4, 32'h3feffc10} /* (6, 15, 18) {real, imag} */,
  {32'hbff0cad2, 32'hbd9654c0} /* (6, 15, 17) {real, imag} */,
  {32'hbf6e8787, 32'hbee91260} /* (6, 15, 16) {real, imag} */,
  {32'hbfdecd56, 32'hc02bdbfc} /* (6, 15, 15) {real, imag} */,
  {32'hbfa71072, 32'hbf88650b} /* (6, 15, 14) {real, imag} */,
  {32'hc00639da, 32'hbf7c2515} /* (6, 15, 13) {real, imag} */,
  {32'hc0571beb, 32'h3f3c2b38} /* (6, 15, 12) {real, imag} */,
  {32'hbfc9e875, 32'h3ee9a57c} /* (6, 15, 11) {real, imag} */,
  {32'hbfd84718, 32'hbfd7fedd} /* (6, 15, 10) {real, imag} */,
  {32'hbf104042, 32'hbfcf5ac0} /* (6, 15, 9) {real, imag} */,
  {32'hbfe6cda7, 32'hbfb11aae} /* (6, 15, 8) {real, imag} */,
  {32'hbf5f657c, 32'h3f2962a8} /* (6, 15, 7) {real, imag} */,
  {32'h3fddcf3a, 32'h3f573d76} /* (6, 15, 6) {real, imag} */,
  {32'h3f2a46ac, 32'hbef03bac} /* (6, 15, 5) {real, imag} */,
  {32'h3e5f638c, 32'hbf424f08} /* (6, 15, 4) {real, imag} */,
  {32'hbfaf0036, 32'hbcfbe5c0} /* (6, 15, 3) {real, imag} */,
  {32'hbf881f37, 32'hbf52df08} /* (6, 15, 2) {real, imag} */,
  {32'h3f02a8f0, 32'h3fde1d3d} /* (6, 15, 1) {real, imag} */,
  {32'hbf235db0, 32'h3ff37094} /* (6, 15, 0) {real, imag} */,
  {32'hbf4612dc, 32'hbd1a5400} /* (6, 14, 31) {real, imag} */,
  {32'hbee814a0, 32'hbff5dd15} /* (6, 14, 30) {real, imag} */,
  {32'h3f057b54, 32'hc0298865} /* (6, 14, 29) {real, imag} */,
  {32'hbfd2637a, 32'h3e77e5b8} /* (6, 14, 28) {real, imag} */,
  {32'h3d98d1f0, 32'hbed1b35c} /* (6, 14, 27) {real, imag} */,
  {32'hbfa98e4d, 32'hbf05a485} /* (6, 14, 26) {real, imag} */,
  {32'hbffc6df6, 32'hbf106053} /* (6, 14, 25) {real, imag} */,
  {32'hc04b3c62, 32'h3fae8ec2} /* (6, 14, 24) {real, imag} */,
  {32'hc024147a, 32'h3ff08563} /* (6, 14, 23) {real, imag} */,
  {32'hc0008dc8, 32'h3d1dcb20} /* (6, 14, 22) {real, imag} */,
  {32'hc05c79f0, 32'h3e73f9f4} /* (6, 14, 21) {real, imag} */,
  {32'hbfa892ce, 32'hbf18d173} /* (6, 14, 20) {real, imag} */,
  {32'h3fa57250, 32'h3f946862} /* (6, 14, 19) {real, imag} */,
  {32'h3fba5690, 32'h400b3169} /* (6, 14, 18) {real, imag} */,
  {32'hbd29d3d0, 32'h3d613e20} /* (6, 14, 17) {real, imag} */,
  {32'h3f25b88e, 32'hbffcc9ea} /* (6, 14, 16) {real, imag} */,
  {32'h3dd180e8, 32'hc03cec38} /* (6, 14, 15) {real, imag} */,
  {32'h3f3a9d08, 32'hbe116404} /* (6, 14, 14) {real, imag} */,
  {32'hbf9de086, 32'hbe83af60} /* (6, 14, 13) {real, imag} */,
  {32'hbfc0437d, 32'hbeddbc50} /* (6, 14, 12) {real, imag} */,
  {32'hbfc3542a, 32'h3ebcc6a8} /* (6, 14, 11) {real, imag} */,
  {32'hc005c333, 32'hbfbb53bb} /* (6, 14, 10) {real, imag} */,
  {32'hbf6f6d96, 32'hbf80abef} /* (6, 14, 9) {real, imag} */,
  {32'hbf64a192, 32'hbe8b4c2c} /* (6, 14, 8) {real, imag} */,
  {32'hbe57f1ec, 32'h401a9fb0} /* (6, 14, 7) {real, imag} */,
  {32'hbeede1a4, 32'h3f953806} /* (6, 14, 6) {real, imag} */,
  {32'h3e31ebc9, 32'hbf4ecc3a} /* (6, 14, 5) {real, imag} */,
  {32'h3f88cf29, 32'hbf692aac} /* (6, 14, 4) {real, imag} */,
  {32'h3eed582e, 32'hbfa6d66a} /* (6, 14, 3) {real, imag} */,
  {32'hbf40f5a4, 32'hbf7ee122} /* (6, 14, 2) {real, imag} */,
  {32'h3d098880, 32'h4020a262} /* (6, 14, 1) {real, imag} */,
  {32'h3e9a6f5e, 32'h3f04e4b8} /* (6, 14, 0) {real, imag} */,
  {32'hbf8c238e, 32'h3f41ba8f} /* (6, 13, 31) {real, imag} */,
  {32'hc0117cf7, 32'h3f1d62fc} /* (6, 13, 30) {real, imag} */,
  {32'hbf4e4235, 32'hbf78f3e6} /* (6, 13, 29) {real, imag} */,
  {32'hbfb18f64, 32'h3f78aae6} /* (6, 13, 28) {real, imag} */,
  {32'h40145366, 32'h3fe58ff4} /* (6, 13, 27) {real, imag} */,
  {32'h3f8f172e, 32'hbf77ffee} /* (6, 13, 26) {real, imag} */,
  {32'hbfd5a220, 32'hbf1a44f9} /* (6, 13, 25) {real, imag} */,
  {32'hc03b12b6, 32'h3ef1a8f0} /* (6, 13, 24) {real, imag} */,
  {32'hc06d2ba5, 32'hbed5317c} /* (6, 13, 23) {real, imag} */,
  {32'h3e50df10, 32'hbee6563c} /* (6, 13, 22) {real, imag} */,
  {32'hbff2f282, 32'h3eb25c32} /* (6, 13, 21) {real, imag} */,
  {32'hc0304186, 32'hbf4e3752} /* (6, 13, 20) {real, imag} */,
  {32'hc016563b, 32'h3f8846ec} /* (6, 13, 19) {real, imag} */,
  {32'hbf856847, 32'h3f1cf69f} /* (6, 13, 18) {real, imag} */,
  {32'h3f711f90, 32'hbea647e0} /* (6, 13, 17) {real, imag} */,
  {32'h3f0a39c3, 32'hbf129d94} /* (6, 13, 16) {real, imag} */,
  {32'h3de2fba8, 32'hc00f6adb} /* (6, 13, 15) {real, imag} */,
  {32'h3faa10bc, 32'hbfe9ba2e} /* (6, 13, 14) {real, imag} */,
  {32'h3fadecde, 32'hbf6f084e} /* (6, 13, 13) {real, imag} */,
  {32'hbf84ece2, 32'hbe683898} /* (6, 13, 12) {real, imag} */,
  {32'hc02eab8e, 32'hbe09a6a8} /* (6, 13, 11) {real, imag} */,
  {32'hc00871c7, 32'h3f13d2d2} /* (6, 13, 10) {real, imag} */,
  {32'h3e648530, 32'h3f5a982a} /* (6, 13, 9) {real, imag} */,
  {32'h3fd16e6a, 32'hc0290810} /* (6, 13, 8) {real, imag} */,
  {32'hbe4f2698, 32'hc026ccf6} /* (6, 13, 7) {real, imag} */,
  {32'hc00b554e, 32'hbfae5513} /* (6, 13, 6) {real, imag} */,
  {32'h3f30d40a, 32'hbf7e74ff} /* (6, 13, 5) {real, imag} */,
  {32'h4011847f, 32'h3e97f093} /* (6, 13, 4) {real, imag} */,
  {32'h3f8c689e, 32'hbf4dab68} /* (6, 13, 3) {real, imag} */,
  {32'h3fb7f518, 32'h3fe2fefe} /* (6, 13, 2) {real, imag} */,
  {32'h3f710ec0, 32'h3ff6715b} /* (6, 13, 1) {real, imag} */,
  {32'h3e16aa00, 32'hbf45236d} /* (6, 13, 0) {real, imag} */,
  {32'hbf98d850, 32'hbf1d2216} /* (6, 12, 31) {real, imag} */,
  {32'hc00bd6de, 32'h3f4e3eeb} /* (6, 12, 30) {real, imag} */,
  {32'h3f3af68c, 32'hbdf4af68} /* (6, 12, 29) {real, imag} */,
  {32'h40298b25, 32'h3ff672da} /* (6, 12, 28) {real, imag} */,
  {32'h404c19da, 32'h3fd28e1e} /* (6, 12, 27) {real, imag} */,
  {32'h3d794710, 32'hbf75857a} /* (6, 12, 26) {real, imag} */,
  {32'hbeca6734, 32'h3eb432a8} /* (6, 12, 25) {real, imag} */,
  {32'hbf1888b4, 32'h3e03a8d0} /* (6, 12, 24) {real, imag} */,
  {32'hbfd8b7d2, 32'hc013912e} /* (6, 12, 23) {real, imag} */,
  {32'h3f0bc792, 32'hc00be16c} /* (6, 12, 22) {real, imag} */,
  {32'h3f17abd2, 32'h3f5350c1} /* (6, 12, 21) {real, imag} */,
  {32'hc02014a8, 32'h3ebb172c} /* (6, 12, 20) {real, imag} */,
  {32'hc0a29628, 32'h3fc735c6} /* (6, 12, 19) {real, imag} */,
  {32'hbf3b67f3, 32'hbedfaa44} /* (6, 12, 18) {real, imag} */,
  {32'h404df554, 32'h3f8e3955} /* (6, 12, 17) {real, imag} */,
  {32'h3ffadaf7, 32'h402700dd} /* (6, 12, 16) {real, imag} */,
  {32'h3f9f7783, 32'hbefb23de} /* (6, 12, 15) {real, imag} */,
  {32'h3f9ec309, 32'hc02106f4} /* (6, 12, 14) {real, imag} */,
  {32'h401d6497, 32'hbfc6fe88} /* (6, 12, 13) {real, imag} */,
  {32'h3f3f1554, 32'h401aa1da} /* (6, 12, 12) {real, imag} */,
  {32'hbf74aaec, 32'h40145e37} /* (6, 12, 11) {real, imag} */,
  {32'hbf5052da, 32'h3fdc2cec} /* (6, 12, 10) {real, imag} */,
  {32'h3d387b90, 32'h3f6b74aa} /* (6, 12, 9) {real, imag} */,
  {32'hbf9d9f8b, 32'hc0208e13} /* (6, 12, 8) {real, imag} */,
  {32'hbf27590a, 32'hbffe63ec} /* (6, 12, 7) {real, imag} */,
  {32'hbfd58922, 32'h3e492c94} /* (6, 12, 6) {real, imag} */,
  {32'h3e3b67c8, 32'h3cf7d700} /* (6, 12, 5) {real, imag} */,
  {32'h3f920dac, 32'hbe2bf854} /* (6, 12, 4) {real, imag} */,
  {32'h3cd55a60, 32'hbfcc4157} /* (6, 12, 3) {real, imag} */,
  {32'h3fe61dfd, 32'h3fb1ac14} /* (6, 12, 2) {real, imag} */,
  {32'h3f2d5014, 32'h3f86bcfa} /* (6, 12, 1) {real, imag} */,
  {32'hbea7d01c, 32'hbfa40d82} /* (6, 12, 0) {real, imag} */,
  {32'hbf156432, 32'h3fa1f1ca} /* (6, 11, 31) {real, imag} */,
  {32'hbf730a94, 32'h400f755e} /* (6, 11, 30) {real, imag} */,
  {32'h3e5f4324, 32'hbf7cc184} /* (6, 11, 29) {real, imag} */,
  {32'h3fc7e691, 32'hbdb5a010} /* (6, 11, 28) {real, imag} */,
  {32'h3fea9341, 32'h3f9a0e4b} /* (6, 11, 27) {real, imag} */,
  {32'h3e08530e, 32'h3ec2453e} /* (6, 11, 26) {real, imag} */,
  {32'hbf2fad8f, 32'hbe5f7738} /* (6, 11, 25) {real, imag} */,
  {32'hbcf701e0, 32'h3e54a9a0} /* (6, 11, 24) {real, imag} */,
  {32'hbf1d916c, 32'hbf309454} /* (6, 11, 23) {real, imag} */,
  {32'h3e55ff88, 32'h3f032c19} /* (6, 11, 22) {real, imag} */,
  {32'h40145a68, 32'h3f22c028} /* (6, 11, 21) {real, imag} */,
  {32'h40097c14, 32'h4011bbf2} /* (6, 11, 20) {real, imag} */,
  {32'h3e9543f9, 32'h3fd2082b} /* (6, 11, 19) {real, imag} */,
  {32'h3ff886a8, 32'hbf800e07} /* (6, 11, 18) {real, imag} */,
  {32'h3fa2ec10, 32'h3fb88038} /* (6, 11, 17) {real, imag} */,
  {32'h3ed813c8, 32'h4099278b} /* (6, 11, 16) {real, imag} */,
  {32'h3fd84c51, 32'h402fd49f} /* (6, 11, 15) {real, imag} */,
  {32'h40213a92, 32'h3ecf921a} /* (6, 11, 14) {real, imag} */,
  {32'h3f93862a, 32'hbfbeee44} /* (6, 11, 13) {real, imag} */,
  {32'h3f198fd4, 32'h3ffddcad} /* (6, 11, 12) {real, imag} */,
  {32'hbed3199e, 32'h406dc2af} /* (6, 11, 11) {real, imag} */,
  {32'h3f1cabfd, 32'h4076594c} /* (6, 11, 10) {real, imag} */,
  {32'h3f033fdd, 32'h401a340d} /* (6, 11, 9) {real, imag} */,
  {32'hbd729520, 32'h3c2f5940} /* (6, 11, 8) {real, imag} */,
  {32'hbdaba424, 32'h400ab998} /* (6, 11, 7) {real, imag} */,
  {32'h3f2cbc96, 32'h40643945} /* (6, 11, 6) {real, imag} */,
  {32'h3fdf6a1e, 32'h3fb86f6a} /* (6, 11, 5) {real, imag} */,
  {32'hbeaea53a, 32'hbcc15460} /* (6, 11, 4) {real, imag} */,
  {32'hbfc45519, 32'h3d997538} /* (6, 11, 3) {real, imag} */,
  {32'hbf1387c9, 32'h3fd5f21e} /* (6, 11, 2) {real, imag} */,
  {32'h402ed45e, 32'h3ff51aa9} /* (6, 11, 1) {real, imag} */,
  {32'h4016cc51, 32'h3fa87d8b} /* (6, 11, 0) {real, imag} */,
  {32'hbebd7422, 32'h3fd3b4f3} /* (6, 10, 31) {real, imag} */,
  {32'h3f1d7750, 32'h4040f412} /* (6, 10, 30) {real, imag} */,
  {32'hbf619e12, 32'h3fd9ea17} /* (6, 10, 29) {real, imag} */,
  {32'hbf5d6b78, 32'hc018bc7d} /* (6, 10, 28) {real, imag} */,
  {32'hbff688f8, 32'hc00d097a} /* (6, 10, 27) {real, imag} */,
  {32'h3f8a6039, 32'h3f0fddf3} /* (6, 10, 26) {real, imag} */,
  {32'h3efbfc46, 32'hbfef834e} /* (6, 10, 25) {real, imag} */,
  {32'h3fae1ce2, 32'hc0542866} /* (6, 10, 24) {real, imag} */,
  {32'h4010eb29, 32'hbf9fb11a} /* (6, 10, 23) {real, imag} */,
  {32'h3fda16c6, 32'h3e9391fc} /* (6, 10, 22) {real, imag} */,
  {32'h3fa71975, 32'h3e79cae6} /* (6, 10, 21) {real, imag} */,
  {32'h405f24dc, 32'h4046ab84} /* (6, 10, 20) {real, imag} */,
  {32'h3f6ebc98, 32'h3fe45e6e} /* (6, 10, 19) {real, imag} */,
  {32'h3f06458c, 32'hbf18abd6} /* (6, 10, 18) {real, imag} */,
  {32'hbfd310dd, 32'h4029460c} /* (6, 10, 17) {real, imag} */,
  {32'hbf03d07e, 32'h40852fe9} /* (6, 10, 16) {real, imag} */,
  {32'hbe3b5fbc, 32'h3db16398} /* (6, 10, 15) {real, imag} */,
  {32'h3e3fd894, 32'hbfaa664c} /* (6, 10, 14) {real, imag} */,
  {32'h3e38d43c, 32'hc0715d70} /* (6, 10, 13) {real, imag} */,
  {32'hbe61e768, 32'h3d906828} /* (6, 10, 12) {real, imag} */,
  {32'hbfd9d8c7, 32'h406082df} /* (6, 10, 11) {real, imag} */,
  {32'hbf7e6357, 32'h40009dfa} /* (6, 10, 10) {real, imag} */,
  {32'h3f169b92, 32'h3d37d300} /* (6, 10, 9) {real, imag} */,
  {32'h40149d06, 32'hbe087335} /* (6, 10, 8) {real, imag} */,
  {32'h4005ce0c, 32'h401b56da} /* (6, 10, 7) {real, imag} */,
  {32'h4062d1a6, 32'h3fe816f9} /* (6, 10, 6) {real, imag} */,
  {32'h3fcebddd, 32'h3f69ce9d} /* (6, 10, 5) {real, imag} */,
  {32'h3f0f9237, 32'h3fbf86b2} /* (6, 10, 4) {real, imag} */,
  {32'h3c790d40, 32'h3fb817ce} /* (6, 10, 3) {real, imag} */,
  {32'hbfbcbbfe, 32'h3fef2718} /* (6, 10, 2) {real, imag} */,
  {32'h402f6d06, 32'h3fa37415} /* (6, 10, 1) {real, imag} */,
  {32'h401c590b, 32'h3edd3bae} /* (6, 10, 0) {real, imag} */,
  {32'h3f83aba3, 32'h3f1211b0} /* (6, 9, 31) {real, imag} */,
  {32'h3f6097b5, 32'h3fb01ada} /* (6, 9, 30) {real, imag} */,
  {32'hbf3135e8, 32'h3f0e36da} /* (6, 9, 29) {real, imag} */,
  {32'h3f88d3c6, 32'hbeefd6dc} /* (6, 9, 28) {real, imag} */,
  {32'h3ea702aa, 32'hbf4c9939} /* (6, 9, 27) {real, imag} */,
  {32'h40045dd4, 32'h3f5855a1} /* (6, 9, 26) {real, imag} */,
  {32'h3f37cf57, 32'hbf4fe79b} /* (6, 9, 25) {real, imag} */,
  {32'h3f045818, 32'hbfaa83bc} /* (6, 9, 24) {real, imag} */,
  {32'h400a0b5b, 32'hc0079cd3} /* (6, 9, 23) {real, imag} */,
  {32'h3fab7c5b, 32'hbefbe81c} /* (6, 9, 22) {real, imag} */,
  {32'hbe8be266, 32'h3e46e948} /* (6, 9, 21) {real, imag} */,
  {32'h3f896ad5, 32'h4047d9be} /* (6, 9, 20) {real, imag} */,
  {32'hbece811a, 32'h3f6621e2} /* (6, 9, 19) {real, imag} */,
  {32'h3f3fb592, 32'hbecbc87a} /* (6, 9, 18) {real, imag} */,
  {32'hbee08e12, 32'h40133b4c} /* (6, 9, 17) {real, imag} */,
  {32'h3f13c444, 32'h3ff87a87} /* (6, 9, 16) {real, imag} */,
  {32'hbf29f3f6, 32'hbffc2c4c} /* (6, 9, 15) {real, imag} */,
  {32'h3ed46814, 32'hbf87a1c6} /* (6, 9, 14) {real, imag} */,
  {32'h3f8d276a, 32'hbfe72e0e} /* (6, 9, 13) {real, imag} */,
  {32'hbd481510, 32'hbd736e40} /* (6, 9, 12) {real, imag} */,
  {32'h3e39b4d8, 32'h3f94df86} /* (6, 9, 11) {real, imag} */,
  {32'h3f675ef4, 32'h3e0203f8} /* (6, 9, 10) {real, imag} */,
  {32'h4022b74b, 32'hbf8f4f7a} /* (6, 9, 9) {real, imag} */,
  {32'h3fe6e470, 32'hc0015910} /* (6, 9, 8) {real, imag} */,
  {32'h3ef6b904, 32'h3ddbf420} /* (6, 9, 7) {real, imag} */,
  {32'h401d1794, 32'h3fa2ad8a} /* (6, 9, 6) {real, imag} */,
  {32'hc0030a2c, 32'h402b3e4c} /* (6, 9, 5) {real, imag} */,
  {32'hbf19b191, 32'h403312ba} /* (6, 9, 4) {real, imag} */,
  {32'h3fae010e, 32'h40192fa0} /* (6, 9, 3) {real, imag} */,
  {32'hbed27235, 32'h4003c0e5} /* (6, 9, 2) {real, imag} */,
  {32'h3f1698e3, 32'h3f1de93c} /* (6, 9, 1) {real, imag} */,
  {32'h3e1ed1b4, 32'hbe9e3398} /* (6, 9, 0) {real, imag} */,
  {32'hbf1b1690, 32'h3f5cd652} /* (6, 8, 31) {real, imag} */,
  {32'hbe03dfa8, 32'h3faea5e2} /* (6, 8, 30) {real, imag} */,
  {32'h3fad3ea0, 32'h3e029ae0} /* (6, 8, 29) {real, imag} */,
  {32'h402ade29, 32'h3f013056} /* (6, 8, 28) {real, imag} */,
  {32'h40775728, 32'h3fe1f80e} /* (6, 8, 27) {real, imag} */,
  {32'h3ff45410, 32'h3e3765b8} /* (6, 8, 26) {real, imag} */,
  {32'hbf3de9e1, 32'h3ef0f164} /* (6, 8, 25) {real, imag} */,
  {32'hbfc7fede, 32'h3fa009e6} /* (6, 8, 24) {real, imag} */,
  {32'hbf235f38, 32'h3de01fa0} /* (6, 8, 23) {real, imag} */,
  {32'hbe254424, 32'hbfc25a36} /* (6, 8, 22) {real, imag} */,
  {32'h3cb10fe0, 32'hbf6acea6} /* (6, 8, 21) {real, imag} */,
  {32'h3f1ca228, 32'h3f9681fa} /* (6, 8, 20) {real, imag} */,
  {32'h3fa084e0, 32'h4017cdfc} /* (6, 8, 19) {real, imag} */,
  {32'h3d99d4a0, 32'h3fd4bf9c} /* (6, 8, 18) {real, imag} */,
  {32'h3f5d4aa1, 32'h3f89f81c} /* (6, 8, 17) {real, imag} */,
  {32'h3e470408, 32'hbdafee50} /* (6, 8, 16) {real, imag} */,
  {32'hbe02ea40, 32'h3fc12ba6} /* (6, 8, 15) {real, imag} */,
  {32'h4051da5f, 32'h3dfba548} /* (6, 8, 14) {real, imag} */,
  {32'h3faf90ee, 32'hbff9c3ce} /* (6, 8, 13) {real, imag} */,
  {32'hbf938f3c, 32'hc060e6e2} /* (6, 8, 12) {real, imag} */,
  {32'hbd9836e8, 32'hbf62b63f} /* (6, 8, 11) {real, imag} */,
  {32'h3f9959f8, 32'h3eb1fb2c} /* (6, 8, 10) {real, imag} */,
  {32'h401332a2, 32'h3ff8292a} /* (6, 8, 9) {real, imag} */,
  {32'h40599234, 32'h3ea2ebce} /* (6, 8, 8) {real, imag} */,
  {32'h4050c55e, 32'h400cc6b5} /* (6, 8, 7) {real, imag} */,
  {32'h3ff3afe7, 32'h40456b71} /* (6, 8, 6) {real, imag} */,
  {32'hc0132a50, 32'h402f039b} /* (6, 8, 5) {real, imag} */,
  {32'hbf9d104b, 32'h400babbc} /* (6, 8, 4) {real, imag} */,
  {32'h3fdc1c36, 32'h3ffdcfa2} /* (6, 8, 3) {real, imag} */,
  {32'hbfa0441a, 32'h40013b4c} /* (6, 8, 2) {real, imag} */,
  {32'hbf532533, 32'hbf8884e0} /* (6, 8, 1) {real, imag} */,
  {32'h3edadfa6, 32'hbfe2120e} /* (6, 8, 0) {real, imag} */,
  {32'h3e837eec, 32'h3fc62576} /* (6, 7, 31) {real, imag} */,
  {32'hbfa580f0, 32'h3f174018} /* (6, 7, 30) {real, imag} */,
  {32'h3d2a73c0, 32'h3f5f960a} /* (6, 7, 29) {real, imag} */,
  {32'h3fc79dd7, 32'h3f5aafdf} /* (6, 7, 28) {real, imag} */,
  {32'h4047c7cc, 32'h3f2ebbbf} /* (6, 7, 27) {real, imag} */,
  {32'h4006dc46, 32'h3f836e04} /* (6, 7, 26) {real, imag} */,
  {32'hbdcd92c0, 32'h3f8f14aa} /* (6, 7, 25) {real, imag} */,
  {32'h3c8aba40, 32'hbed7eabc} /* (6, 7, 24) {real, imag} */,
  {32'h3d9928d0, 32'h402c4c39} /* (6, 7, 23) {real, imag} */,
  {32'hbe476a28, 32'h3efd85f4} /* (6, 7, 22) {real, imag} */,
  {32'h3ff948b8, 32'hbff895dd} /* (6, 7, 21) {real, imag} */,
  {32'h3fcd29c0, 32'hbe615e9c} /* (6, 7, 20) {real, imag} */,
  {32'h40368d35, 32'h408ebf56} /* (6, 7, 19) {real, imag} */,
  {32'h3f94300c, 32'h3fefa77a} /* (6, 7, 18) {real, imag} */,
  {32'h3e582b90, 32'h3f258b34} /* (6, 7, 17) {real, imag} */,
  {32'hbf16097a, 32'h3f874f29} /* (6, 7, 16) {real, imag} */,
  {32'hbf19b58c, 32'h40220a82} /* (6, 7, 15) {real, imag} */,
  {32'h3fdcfbd4, 32'h3f9e0cea} /* (6, 7, 14) {real, imag} */,
  {32'h3fe10bbc, 32'hbf56490e} /* (6, 7, 13) {real, imag} */,
  {32'h3ebbaa9a, 32'hbf9aaa9d} /* (6, 7, 12) {real, imag} */,
  {32'h3fac9a57, 32'hbeaa5ed2} /* (6, 7, 11) {real, imag} */,
  {32'hbd916cf0, 32'h40286dfb} /* (6, 7, 10) {real, imag} */,
  {32'h3ea13420, 32'h40852c73} /* (6, 7, 9) {real, imag} */,
  {32'h3fb2aeca, 32'h3f9a2e31} /* (6, 7, 8) {real, imag} */,
  {32'h4023e852, 32'h405a5a93} /* (6, 7, 7) {real, imag} */,
  {32'h3e83636a, 32'h4090ec44} /* (6, 7, 6) {real, imag} */,
  {32'hbf59e2fe, 32'h3ffae81a} /* (6, 7, 5) {real, imag} */,
  {32'hbf56d9cc, 32'hbf6db777} /* (6, 7, 4) {real, imag} */,
  {32'h3f1fbc23, 32'h3f0e6f58} /* (6, 7, 3) {real, imag} */,
  {32'hbf96143a, 32'h3fad052b} /* (6, 7, 2) {real, imag} */,
  {32'hbe6d926c, 32'h3fc3a9df} /* (6, 7, 1) {real, imag} */,
  {32'h3f8039e4, 32'h3f8bd933} /* (6, 7, 0) {real, imag} */,
  {32'h3e756870, 32'h3ed0aa88} /* (6, 6, 31) {real, imag} */,
  {32'h3ebda694, 32'hbd8e9f38} /* (6, 6, 30) {real, imag} */,
  {32'hbf27065e, 32'hbee55db4} /* (6, 6, 29) {real, imag} */,
  {32'hbf537536, 32'hbed077c6} /* (6, 6, 28) {real, imag} */,
  {32'h3f43e10c, 32'hbfcd576e} /* (6, 6, 27) {real, imag} */,
  {32'h3fe0cc50, 32'h3eb53034} /* (6, 6, 26) {real, imag} */,
  {32'h3f99a10d, 32'h3f660d92} /* (6, 6, 25) {real, imag} */,
  {32'h3f89204c, 32'h3fcea037} /* (6, 6, 24) {real, imag} */,
  {32'h3f438c03, 32'h4070bc50} /* (6, 6, 23) {real, imag} */,
  {32'hbdd0ad18, 32'h4020309c} /* (6, 6, 22) {real, imag} */,
  {32'h3f959ed5, 32'h3faaf5f8} /* (6, 6, 21) {real, imag} */,
  {32'h3ff3ca49, 32'hbf2c3120} /* (6, 6, 20) {real, imag} */,
  {32'h400c91ca, 32'h3fc54760} /* (6, 6, 19) {real, imag} */,
  {32'h3e4e5ec8, 32'h3fa4f2d0} /* (6, 6, 18) {real, imag} */,
  {32'hbedadf10, 32'hbf77d0cb} /* (6, 6, 17) {real, imag} */,
  {32'h3f7fb6d2, 32'h3f4e96e2} /* (6, 6, 16) {real, imag} */,
  {32'h40033092, 32'h3f3358c8} /* (6, 6, 15) {real, imag} */,
  {32'h3f7da980, 32'h3fbbe416} /* (6, 6, 14) {real, imag} */,
  {32'h3f781329, 32'h3f34910b} /* (6, 6, 13) {real, imag} */,
  {32'hbf2635cd, 32'hbd4f19d0} /* (6, 6, 12) {real, imag} */,
  {32'h3fb4df81, 32'hbf349ebd} /* (6, 6, 11) {real, imag} */,
  {32'h3fffbf39, 32'h3f877a67} /* (6, 6, 10) {real, imag} */,
  {32'hbedf9db4, 32'h404ea182} /* (6, 6, 9) {real, imag} */,
  {32'h3fd4215e, 32'h3ee3e7a6} /* (6, 6, 8) {real, imag} */,
  {32'h403c46e2, 32'h400e8fc0} /* (6, 6, 7) {real, imag} */,
  {32'h3f63a0ce, 32'h3fe7f4bc} /* (6, 6, 6) {real, imag} */,
  {32'h3f8ad952, 32'hbd4c4db0} /* (6, 6, 5) {real, imag} */,
  {32'h3ec6aab4, 32'hbfcc8c78} /* (6, 6, 4) {real, imag} */,
  {32'h3ec1d5e6, 32'h3e0e85c4} /* (6, 6, 3) {real, imag} */,
  {32'h3f25b8b2, 32'hbe189ff8} /* (6, 6, 2) {real, imag} */,
  {32'h3fcc1236, 32'h3d518700} /* (6, 6, 1) {real, imag} */,
  {32'h3f86c974, 32'h3f9f6fb9} /* (6, 6, 0) {real, imag} */,
  {32'h3e9c441c, 32'h3ef58270} /* (6, 5, 31) {real, imag} */,
  {32'hbe7ea4fc, 32'h3ee38b92} /* (6, 5, 30) {real, imag} */,
  {32'hbf5cf1c2, 32'hbe8d9da0} /* (6, 5, 29) {real, imag} */,
  {32'hbff14e4e, 32'h3f6d9aa6} /* (6, 5, 28) {real, imag} */,
  {32'hbefb5bac, 32'hc0010788} /* (6, 5, 27) {real, imag} */,
  {32'hbd086cc0, 32'hbeb63172} /* (6, 5, 26) {real, imag} */,
  {32'h3f8e64ec, 32'hbfb46f7d} /* (6, 5, 25) {real, imag} */,
  {32'h3f95ecd4, 32'hbf286a42} /* (6, 5, 24) {real, imag} */,
  {32'h3f5fe954, 32'h3f3d99cc} /* (6, 5, 23) {real, imag} */,
  {32'hbfd53a05, 32'h402b8a5e} /* (6, 5, 22) {real, imag} */,
  {32'hc06d6ddc, 32'h3fa778a0} /* (6, 5, 21) {real, imag} */,
  {32'hc01bd3b8, 32'h3f2eff9e} /* (6, 5, 20) {real, imag} */,
  {32'h3e5aac04, 32'h3ebb2a7e} /* (6, 5, 19) {real, imag} */,
  {32'h3fb570a9, 32'hbf9e491e} /* (6, 5, 18) {real, imag} */,
  {32'hbfc3daae, 32'hbfe84e5e} /* (6, 5, 17) {real, imag} */,
  {32'hbfbebf69, 32'h3ffc5285} /* (6, 5, 16) {real, imag} */,
  {32'h3f3241c2, 32'h3fefe0c9} /* (6, 5, 15) {real, imag} */,
  {32'h400c4ca2, 32'h401cf5e0} /* (6, 5, 14) {real, imag} */,
  {32'h3f453aef, 32'h3f503bf2} /* (6, 5, 13) {real, imag} */,
  {32'hbf9983c2, 32'h3e842848} /* (6, 5, 12) {real, imag} */,
  {32'hbf8bd8a4, 32'hbf8252b6} /* (6, 5, 11) {real, imag} */,
  {32'h3f989bbe, 32'hbf897732} /* (6, 5, 10) {real, imag} */,
  {32'h40290a04, 32'h3d205b18} /* (6, 5, 9) {real, imag} */,
  {32'h4037c756, 32'h3f8a5578} /* (6, 5, 8) {real, imag} */,
  {32'h402195e4, 32'h405cbeeb} /* (6, 5, 7) {real, imag} */,
  {32'h3b711c00, 32'h401c7e30} /* (6, 5, 6) {real, imag} */,
  {32'hbf39cd18, 32'h3d2a8440} /* (6, 5, 5) {real, imag} */,
  {32'hbf339d51, 32'hbdfb8430} /* (6, 5, 4) {real, imag} */,
  {32'hbf6facbf, 32'hbf08a71c} /* (6, 5, 3) {real, imag} */,
  {32'hbfc476ad, 32'hbeed3ff4} /* (6, 5, 2) {real, imag} */,
  {32'hbe7e6e88, 32'hbf90109a} /* (6, 5, 1) {real, imag} */,
  {32'hbf613a34, 32'h3f346ea6} /* (6, 5, 0) {real, imag} */,
  {32'h3f81cff4, 32'h3f55485f} /* (6, 4, 31) {real, imag} */,
  {32'h40016dfc, 32'h3fc1fde4} /* (6, 4, 30) {real, imag} */,
  {32'h3f3e57a3, 32'h3eb860c0} /* (6, 4, 29) {real, imag} */,
  {32'hbfa2dfbb, 32'h3e03f660} /* (6, 4, 28) {real, imag} */,
  {32'hc004f95c, 32'h3fa3c21d} /* (6, 4, 27) {real, imag} */,
  {32'hbf411f53, 32'h40785c09} /* (6, 4, 26) {real, imag} */,
  {32'hbd966314, 32'h400b54d6} /* (6, 4, 25) {real, imag} */,
  {32'hbf1bba5f, 32'hbf688270} /* (6, 4, 24) {real, imag} */,
  {32'h3f83063e, 32'hbfd8e372} /* (6, 4, 23) {real, imag} */,
  {32'h3f8f1904, 32'h3fd55830} /* (6, 4, 22) {real, imag} */,
  {32'hbfb5348c, 32'h3f1818c4} /* (6, 4, 21) {real, imag} */,
  {32'hc016539c, 32'h3f82dc7c} /* (6, 4, 20) {real, imag} */,
  {32'hbf6201e6, 32'hbfa9543b} /* (6, 4, 19) {real, imag} */,
  {32'h3f0371b9, 32'hc09b09bc} /* (6, 4, 18) {real, imag} */,
  {32'h3f1e8c2a, 32'hc01c1732} /* (6, 4, 17) {real, imag} */,
  {32'hbf8b30cd, 32'hbde7c220} /* (6, 4, 16) {real, imag} */,
  {32'hc0036b89, 32'h3fcfc9bc} /* (6, 4, 15) {real, imag} */,
  {32'h3fb115d2, 32'h405589e6} /* (6, 4, 14) {real, imag} */,
  {32'hbd0d0d70, 32'h40029086} /* (6, 4, 13) {real, imag} */,
  {32'hbf38639e, 32'h3e94bc0c} /* (6, 4, 12) {real, imag} */,
  {32'hbe8de412, 32'hbf9b86ce} /* (6, 4, 11) {real, imag} */,
  {32'h3f0b8d0a, 32'hbf8da1b1} /* (6, 4, 10) {real, imag} */,
  {32'h3fdb79e2, 32'hbfdf2635} /* (6, 4, 9) {real, imag} */,
  {32'hbf4b6cbe, 32'h3fada844} /* (6, 4, 8) {real, imag} */,
  {32'hbe8c35a8, 32'h3fedb118} /* (6, 4, 7) {real, imag} */,
  {32'hbe9eeb7a, 32'h401768e7} /* (6, 4, 6) {real, imag} */,
  {32'h3f4f66d0, 32'h40024ba0} /* (6, 4, 5) {real, imag} */,
  {32'h3e7ee268, 32'h3fb0b6f9} /* (6, 4, 4) {real, imag} */,
  {32'hc00ab8fa, 32'h3da90ee0} /* (6, 4, 3) {real, imag} */,
  {32'hc02556a2, 32'hbf0abfa0} /* (6, 4, 2) {real, imag} */,
  {32'h3ee48794, 32'hbd9d2800} /* (6, 4, 1) {real, imag} */,
  {32'hbf0a84d3, 32'h3f751d13} /* (6, 4, 0) {real, imag} */,
  {32'hbe9c5ab0, 32'h3f947c88} /* (6, 3, 31) {real, imag} */,
  {32'h3fa679a2, 32'h4010b770} /* (6, 3, 30) {real, imag} */,
  {32'h3fabb16f, 32'hbf67c4e2} /* (6, 3, 29) {real, imag} */,
  {32'h3fa66b21, 32'hbff21b34} /* (6, 3, 28) {real, imag} */,
  {32'hbfc50bda, 32'h3f7ae8f0} /* (6, 3, 27) {real, imag} */,
  {32'hc0072554, 32'h405a4ca2} /* (6, 3, 26) {real, imag} */,
  {32'hbf9a1c68, 32'h402073a5} /* (6, 3, 25) {real, imag} */,
  {32'hc003588d, 32'hbec5bfa6} /* (6, 3, 24) {real, imag} */,
  {32'hbe74ca08, 32'hbedfc52e} /* (6, 3, 23) {real, imag} */,
  {32'h3fc4e584, 32'h3f6d5018} /* (6, 3, 22) {real, imag} */,
  {32'hbe9f117e, 32'h3e97b70c} /* (6, 3, 21) {real, imag} */,
  {32'h3fae32ef, 32'hbf3eda2a} /* (6, 3, 20) {real, imag} */,
  {32'h40143319, 32'hbe99462c} /* (6, 3, 19) {real, imag} */,
  {32'hbfe33621, 32'h3e8a88ac} /* (6, 3, 18) {real, imag} */,
  {32'hbf13ca1e, 32'hbfb4efb4} /* (6, 3, 17) {real, imag} */,
  {32'h3f87f8c2, 32'hc00c5539} /* (6, 3, 16) {real, imag} */,
  {32'hbebe78f1, 32'hbfff26a2} /* (6, 3, 15) {real, imag} */,
  {32'h3ec280f6, 32'hbf244460} /* (6, 3, 14) {real, imag} */,
  {32'hc000af84, 32'h3d5537a0} /* (6, 3, 13) {real, imag} */,
  {32'hbef812c0, 32'hbfbbd5cb} /* (6, 3, 12) {real, imag} */,
  {32'h3fb02355, 32'hc05620ae} /* (6, 3, 11) {real, imag} */,
  {32'hbf2cd5a6, 32'hc0080708} /* (6, 3, 10) {real, imag} */,
  {32'hbf27f3d0, 32'hbd97d198} /* (6, 3, 9) {real, imag} */,
  {32'hbfe38bf1, 32'h3f6eefc2} /* (6, 3, 8) {real, imag} */,
  {32'h3e1a4ba0, 32'h40248e4b} /* (6, 3, 7) {real, imag} */,
  {32'hbf2f19bd, 32'h4078063e} /* (6, 3, 6) {real, imag} */,
  {32'hbdd56e14, 32'h407da054} /* (6, 3, 5) {real, imag} */,
  {32'h3f29a2f2, 32'h401d8390} /* (6, 3, 4) {real, imag} */,
  {32'hbf76e542, 32'h3f81669c} /* (6, 3, 3) {real, imag} */,
  {32'h3de505dc, 32'h3e8039c4} /* (6, 3, 2) {real, imag} */,
  {32'h4007806b, 32'hbe360d80} /* (6, 3, 1) {real, imag} */,
  {32'h3f41b860, 32'h3f8bce09} /* (6, 3, 0) {real, imag} */,
  {32'hbf1edfea, 32'h3f1c2741} /* (6, 2, 31) {real, imag} */,
  {32'h3f5f4a93, 32'h3f8fee7e} /* (6, 2, 30) {real, imag} */,
  {32'hbf59e182, 32'hbdf48630} /* (6, 2, 29) {real, imag} */,
  {32'hbea75850, 32'hbffc28c3} /* (6, 2, 28) {real, imag} */,
  {32'h3f0b298c, 32'hbfaaf4b5} /* (6, 2, 27) {real, imag} */,
  {32'hc0397f8c, 32'h3fa34728} /* (6, 2, 26) {real, imag} */,
  {32'hc00a91ad, 32'h3f2b82c8} /* (6, 2, 25) {real, imag} */,
  {32'hbfe12932, 32'hbf6f69db} /* (6, 2, 24) {real, imag} */,
  {32'h3c86dc40, 32'hc02bff32} /* (6, 2, 23) {real, imag} */,
  {32'h3f9238c8, 32'hbfbbf398} /* (6, 2, 22) {real, imag} */,
  {32'h3fa535a2, 32'hc009520b} /* (6, 2, 21) {real, imag} */,
  {32'h4085f3a6, 32'hc07300c0} /* (6, 2, 20) {real, imag} */,
  {32'h409a547c, 32'h3ec688d0} /* (6, 2, 19) {real, imag} */,
  {32'h3f9b80da, 32'h401e139d} /* (6, 2, 18) {real, imag} */,
  {32'h3f10778a, 32'h4041ed86} /* (6, 2, 17) {real, imag} */,
  {32'h3faa767a, 32'h3f56fc64} /* (6, 2, 16) {real, imag} */,
  {32'hbf1855bc, 32'hbf2a25ee} /* (6, 2, 15) {real, imag} */,
  {32'hbd78c3c0, 32'hbfbc94da} /* (6, 2, 14) {real, imag} */,
  {32'hbe9619e0, 32'hc019f3bf} /* (6, 2, 13) {real, imag} */,
  {32'hbf56adef, 32'hbf5fe2a2} /* (6, 2, 12) {real, imag} */,
  {32'hbec819dc, 32'hc0698906} /* (6, 2, 11) {real, imag} */,
  {32'hbf5fb3f4, 32'hbeed2824} /* (6, 2, 10) {real, imag} */,
  {32'h3f188d26, 32'h3f599c68} /* (6, 2, 9) {real, imag} */,
  {32'hbe00b360, 32'h3e9086a4} /* (6, 2, 8) {real, imag} */,
  {32'hbd375030, 32'h3fbc7c1a} /* (6, 2, 7) {real, imag} */,
  {32'hbf84d459, 32'h3fa8aae3} /* (6, 2, 6) {real, imag} */,
  {32'hc0109e0a, 32'h4032f131} /* (6, 2, 5) {real, imag} */,
  {32'hbfb47204, 32'h3f0447d0} /* (6, 2, 4) {real, imag} */,
  {32'h3f7cfc2b, 32'h3f099087} /* (6, 2, 3) {real, imag} */,
  {32'h3f8acfda, 32'h3f5ac0b0} /* (6, 2, 2) {real, imag} */,
  {32'h3f46ba52, 32'hbf0260a6} /* (6, 2, 1) {real, imag} */,
  {32'hbea6b6e4, 32'hbed0d324} /* (6, 2, 0) {real, imag} */,
  {32'h3f8b66c6, 32'h3ca28600} /* (6, 1, 31) {real, imag} */,
  {32'h40030aca, 32'h3e764c08} /* (6, 1, 30) {real, imag} */,
  {32'h3f66a61b, 32'hbec4a988} /* (6, 1, 29) {real, imag} */,
  {32'h3e62ce40, 32'hbfd89acf} /* (6, 1, 28) {real, imag} */,
  {32'h3fc0973a, 32'hbf7e988e} /* (6, 1, 27) {real, imag} */,
  {32'hbfdb18bc, 32'h3faa59bd} /* (6, 1, 26) {real, imag} */,
  {32'hc00aed21, 32'h3fe7db67} /* (6, 1, 25) {real, imag} */,
  {32'hbfa788e4, 32'h3e0ca958} /* (6, 1, 24) {real, imag} */,
  {32'hbe65ae48, 32'hc05ba102} /* (6, 1, 23) {real, imag} */,
  {32'hbf67ac4f, 32'hbf9836a6} /* (6, 1, 22) {real, imag} */,
  {32'hba2a4400, 32'hc099634d} /* (6, 1, 21) {real, imag} */,
  {32'h3eabce68, 32'hc02b739a} /* (6, 1, 20) {real, imag} */,
  {32'h3ffe7c8c, 32'h3f5df26c} /* (6, 1, 19) {real, imag} */,
  {32'h3f651da8, 32'h3d87d760} /* (6, 1, 18) {real, imag} */,
  {32'hbf0d38ae, 32'h3fb7a6ce} /* (6, 1, 17) {real, imag} */,
  {32'hbf53db6a, 32'hbd877c68} /* (6, 1, 16) {real, imag} */,
  {32'hbfc8480c, 32'hbf1b8473} /* (6, 1, 15) {real, imag} */,
  {32'h3fa2af52, 32'hc029cde9} /* (6, 1, 14) {real, imag} */,
  {32'h3f9174c0, 32'hc0644110} /* (6, 1, 13) {real, imag} */,
  {32'h3f5342d0, 32'hbf8d1db8} /* (6, 1, 12) {real, imag} */,
  {32'h3e005e50, 32'hbfdd6fc0} /* (6, 1, 11) {real, imag} */,
  {32'hbefafa6e, 32'h3ece91cc} /* (6, 1, 10) {real, imag} */,
  {32'h3f57b870, 32'h3f7463a0} /* (6, 1, 9) {real, imag} */,
  {32'h3f3bdfa8, 32'hbf5e98ba} /* (6, 1, 8) {real, imag} */,
  {32'hbf71c51e, 32'h3e145b68} /* (6, 1, 7) {real, imag} */,
  {32'hbfb223ca, 32'hbf305602} /* (6, 1, 6) {real, imag} */,
  {32'hc023b622, 32'h3f2d58bc} /* (6, 1, 5) {real, imag} */,
  {32'hbfcd5595, 32'h3e637068} /* (6, 1, 4) {real, imag} */,
  {32'hbf24ac61, 32'hbf4222aa} /* (6, 1, 3) {real, imag} */,
  {32'hbef80bf7, 32'h3f967d27} /* (6, 1, 2) {real, imag} */,
  {32'h3fefa6fa, 32'hbf8ce932} /* (6, 1, 1) {real, imag} */,
  {32'h3f0936d1, 32'hbfe27d22} /* (6, 1, 0) {real, imag} */,
  {32'h3fab7342, 32'h3f12af5f} /* (6, 0, 31) {real, imag} */,
  {32'h3fd0d210, 32'h3ede6772} /* (6, 0, 30) {real, imag} */,
  {32'h3fb08fcb, 32'hbed05c10} /* (6, 0, 29) {real, imag} */,
  {32'h3fe72478, 32'hbf3d70e8} /* (6, 0, 28) {real, imag} */,
  {32'h3f60b7fb, 32'hbe906b6a} /* (6, 0, 27) {real, imag} */,
  {32'hbfe268dc, 32'h3f23faeb} /* (6, 0, 26) {real, imag} */,
  {32'hbf37043c, 32'h3e6973ba} /* (6, 0, 25) {real, imag} */,
  {32'hbe44f1a0, 32'h3e4b97b4} /* (6, 0, 24) {real, imag} */,
  {32'h3cf343c0, 32'hbd7e8fa0} /* (6, 0, 23) {real, imag} */,
  {32'hbf8ac449, 32'h3f18bbd2} /* (6, 0, 22) {real, imag} */,
  {32'hbf2a2be6, 32'hbfe584a3} /* (6, 0, 21) {real, imag} */,
  {32'hbfdd4f1e, 32'hbf567398} /* (6, 0, 20) {real, imag} */,
  {32'hbe4815e0, 32'hbe8b972e} /* (6, 0, 19) {real, imag} */,
  {32'hbf2349be, 32'hbd1db850} /* (6, 0, 18) {real, imag} */,
  {32'hbfcf0b44, 32'hbf1e355b} /* (6, 0, 17) {real, imag} */,
  {32'hbfc9ab66, 32'hbebe88c2} /* (6, 0, 16) {real, imag} */,
  {32'hbf4b9ace, 32'hbe797ec8} /* (6, 0, 15) {real, imag} */,
  {32'h400413e3, 32'hbff0236e} /* (6, 0, 14) {real, imag} */,
  {32'h3fba0535, 32'hbfb8d942} /* (6, 0, 13) {real, imag} */,
  {32'h3ff7b938, 32'h3f84bb18} /* (6, 0, 12) {real, imag} */,
  {32'h400ed162, 32'hbe201a20} /* (6, 0, 11) {real, imag} */,
  {32'h3fc9e64f, 32'hbfbffd6e} /* (6, 0, 10) {real, imag} */,
  {32'h3edca77e, 32'hbe6c1190} /* (6, 0, 9) {real, imag} */,
  {32'hbf1c15dc, 32'hbfa7a0be} /* (6, 0, 8) {real, imag} */,
  {32'hbfff8945, 32'hbf8347b4} /* (6, 0, 7) {real, imag} */,
  {32'hc01f47ef, 32'hbf25f69e} /* (6, 0, 6) {real, imag} */,
  {32'hbf6f4e72, 32'hbf7e00a5} /* (6, 0, 5) {real, imag} */,
  {32'hbe79acf0, 32'hbf532ece} /* (6, 0, 4) {real, imag} */,
  {32'h3eb4b83a, 32'hbf903a80} /* (6, 0, 3) {real, imag} */,
  {32'h3f7e7832, 32'h3f307c09} /* (6, 0, 2) {real, imag} */,
  {32'h3ffcf58c, 32'hbedd6140} /* (6, 0, 1) {real, imag} */,
  {32'h3f44131e, 32'hbf8be2da} /* (6, 0, 0) {real, imag} */,
  {32'h3f86cc84, 32'hbec18892} /* (5, 31, 31) {real, imag} */,
  {32'h3fdf1535, 32'hbee77387} /* (5, 31, 30) {real, imag} */,
  {32'hbe061118, 32'hc01076e4} /* (5, 31, 29) {real, imag} */,
  {32'h3e4449ec, 32'hbfcf2648} /* (5, 31, 28) {real, imag} */,
  {32'h400272b3, 32'hc01c52d6} /* (5, 31, 27) {real, imag} */,
  {32'h402e0a5a, 32'hc05accf5} /* (5, 31, 26) {real, imag} */,
  {32'h40192240, 32'hc0025582} /* (5, 31, 25) {real, imag} */,
  {32'h400943aa, 32'hbfc65a0d} /* (5, 31, 24) {real, imag} */,
  {32'h3e80fc19, 32'hbf785c01} /* (5, 31, 23) {real, imag} */,
  {32'hbeafc95d, 32'hbfb0e738} /* (5, 31, 22) {real, imag} */,
  {32'hbfcb4d89, 32'h3f516cfb} /* (5, 31, 21) {real, imag} */,
  {32'hc00ff9dc, 32'h3f9f0c16} /* (5, 31, 20) {real, imag} */,
  {32'hbfc41404, 32'hbe40b88d} /* (5, 31, 19) {real, imag} */,
  {32'h3d16c210, 32'h3f4e7b24} /* (5, 31, 18) {real, imag} */,
  {32'hbf30c22c, 32'h40238b02} /* (5, 31, 17) {real, imag} */,
  {32'h3ecf103f, 32'hbdbd2790} /* (5, 31, 16) {real, imag} */,
  {32'h3f1ae8e8, 32'hbe76c586} /* (5, 31, 15) {real, imag} */,
  {32'hbf7f3012, 32'h3d795850} /* (5, 31, 14) {real, imag} */,
  {32'h3e117bcf, 32'h3fdb5c0c} /* (5, 31, 13) {real, imag} */,
  {32'h3f48669c, 32'h4015dac6} /* (5, 31, 12) {real, imag} */,
  {32'hbe0062b2, 32'h3f99349c} /* (5, 31, 11) {real, imag} */,
  {32'h3fb7ee3c, 32'hbf478444} /* (5, 31, 10) {real, imag} */,
  {32'h3f647396, 32'hbf04af19} /* (5, 31, 9) {real, imag} */,
  {32'hbe846a9c, 32'hbf3fee78} /* (5, 31, 8) {real, imag} */,
  {32'h3ec1a468, 32'hbe9cf84a} /* (5, 31, 7) {real, imag} */,
  {32'h3e92bae4, 32'hbfc9d1da} /* (5, 31, 6) {real, imag} */,
  {32'h3e46a7e2, 32'hc013c3cd} /* (5, 31, 5) {real, imag} */,
  {32'hbf10964a, 32'hbff121ec} /* (5, 31, 4) {real, imag} */,
  {32'h3d5d36c0, 32'hc01f142d} /* (5, 31, 3) {real, imag} */,
  {32'h3e58e068, 32'hbfb91aad} /* (5, 31, 2) {real, imag} */,
  {32'hbec240d6, 32'hbfc422f1} /* (5, 31, 1) {real, imag} */,
  {32'h3f186bc4, 32'h3d8533d6} /* (5, 31, 0) {real, imag} */,
  {32'h3f84cf59, 32'hbf0e53aa} /* (5, 30, 31) {real, imag} */,
  {32'h403ef993, 32'hbfdfa33c} /* (5, 30, 30) {real, imag} */,
  {32'h3fc3f0b0, 32'hc0603b9a} /* (5, 30, 29) {real, imag} */,
  {32'h3f76e93e, 32'hc008fe3c} /* (5, 30, 28) {real, imag} */,
  {32'h3fc7d8d8, 32'hc07db2b7} /* (5, 30, 27) {real, imag} */,
  {32'h3f4f42b5, 32'hc09bb444} /* (5, 30, 26) {real, imag} */,
  {32'h3fcb3439, 32'hc056957e} /* (5, 30, 25) {real, imag} */,
  {32'h3ff34eec, 32'hc02c00f8} /* (5, 30, 24) {real, imag} */,
  {32'h40185fcd, 32'hc021d02c} /* (5, 30, 23) {real, imag} */,
  {32'h4047c284, 32'hbfe1f5e0} /* (5, 30, 22) {real, imag} */,
  {32'hbf2d82d2, 32'h3f4b33ce} /* (5, 30, 21) {real, imag} */,
  {32'hc08e1466, 32'h40695309} /* (5, 30, 20) {real, imag} */,
  {32'hc0b3e85e, 32'h3fbe79b5} /* (5, 30, 19) {real, imag} */,
  {32'hbfaae44a, 32'h4036ecee} /* (5, 30, 18) {real, imag} */,
  {32'hbef71f6e, 32'h40953d31} /* (5, 30, 17) {real, imag} */,
  {32'h3f72d973, 32'h4056221a} /* (5, 30, 16) {real, imag} */,
  {32'hbf7ec28f, 32'h3ffafb1e} /* (5, 30, 15) {real, imag} */,
  {32'hbf9133e2, 32'h3f3bc508} /* (5, 30, 14) {real, imag} */,
  {32'hbd1c2910, 32'h3fe4e679} /* (5, 30, 13) {real, imag} */,
  {32'hbf51f00d, 32'h4081ff34} /* (5, 30, 12) {real, imag} */,
  {32'hbfda083e, 32'h406bdefe} /* (5, 30, 11) {real, imag} */,
  {32'h401726ff, 32'hbebe7211} /* (5, 30, 10) {real, imag} */,
  {32'h400a81f4, 32'hbffd28a0} /* (5, 30, 9) {real, imag} */,
  {32'hbec4d87c, 32'hc00afbf8} /* (5, 30, 8) {real, imag} */,
  {32'h3f1581db, 32'hbfec728a} /* (5, 30, 7) {real, imag} */,
  {32'h3fd99ea3, 32'hc04d6876} /* (5, 30, 6) {real, imag} */,
  {32'h3e6ac088, 32'hc08a3f40} /* (5, 30, 5) {real, imag} */,
  {32'h3ea2e182, 32'hc010faf4} /* (5, 30, 4) {real, imag} */,
  {32'hbea90298, 32'hbfee4112} /* (5, 30, 3) {real, imag} */,
  {32'h402b34f2, 32'hbee70914} /* (5, 30, 2) {real, imag} */,
  {32'h3d264f70, 32'hc0074ee2} /* (5, 30, 1) {real, imag} */,
  {32'hbf5523e6, 32'hbf897266} /* (5, 30, 0) {real, imag} */,
  {32'h3eac693a, 32'hbfb690a5} /* (5, 29, 31) {real, imag} */,
  {32'h403013f3, 32'hc0469abe} /* (5, 29, 30) {real, imag} */,
  {32'h40139ecc, 32'hc03b58cc} /* (5, 29, 29) {real, imag} */,
  {32'h3fb49807, 32'hc0269228} /* (5, 29, 28) {real, imag} */,
  {32'h3fe2c84f, 32'hc0686954} /* (5, 29, 27) {real, imag} */,
  {32'hbf78120f, 32'hc035d4ad} /* (5, 29, 26) {real, imag} */,
  {32'h3d8c4a38, 32'hc064729d} /* (5, 29, 25) {real, imag} */,
  {32'h3f483d04, 32'hc01497dc} /* (5, 29, 24) {real, imag} */,
  {32'h400b5a68, 32'hbf901336} /* (5, 29, 23) {real, imag} */,
  {32'h3f963edf, 32'h3eea6be8} /* (5, 29, 22) {real, imag} */,
  {32'hbe1cca98, 32'hbfd19d8c} /* (5, 29, 21) {real, imag} */,
  {32'hbff7ec54, 32'h3f256b10} /* (5, 29, 20) {real, imag} */,
  {32'hc0c807c5, 32'hbe4917c0} /* (5, 29, 19) {real, imag} */,
  {32'hc077175b, 32'h3f0bf190} /* (5, 29, 18) {real, imag} */,
  {32'hc07f163e, 32'h403e8162} /* (5, 29, 17) {real, imag} */,
  {32'hc05c6a56, 32'h40963db2} /* (5, 29, 16) {real, imag} */,
  {32'hbfe81e9c, 32'h408881bb} /* (5, 29, 15) {real, imag} */,
  {32'h3fcdfa14, 32'h4005201e} /* (5, 29, 14) {real, imag} */,
  {32'hbe68e174, 32'h3ee8178a} /* (5, 29, 13) {real, imag} */,
  {32'hc0592792, 32'h40012244} /* (5, 29, 12) {real, imag} */,
  {32'hc04ae31e, 32'h3ffaecaf} /* (5, 29, 11) {real, imag} */,
  {32'h3f5a3e72, 32'hbf9c822c} /* (5, 29, 10) {real, imag} */,
  {32'h408c797d, 32'hbfdc052d} /* (5, 29, 9) {real, imag} */,
  {32'h4017080c, 32'hc03076fc} /* (5, 29, 8) {real, imag} */,
  {32'h3f8944ba, 32'hc04fb234} /* (5, 29, 7) {real, imag} */,
  {32'h40402ec6, 32'hbff71c51} /* (5, 29, 6) {real, imag} */,
  {32'h404a4d4e, 32'hc070715c} /* (5, 29, 5) {real, imag} */,
  {32'h3ffa049e, 32'hc0007e30} /* (5, 29, 4) {real, imag} */,
  {32'hbe76a1d6, 32'hc00d697d} /* (5, 29, 3) {real, imag} */,
  {32'h4084f2d5, 32'hbfb76f5c} /* (5, 29, 2) {real, imag} */,
  {32'h40774c0b, 32'hc012e410} /* (5, 29, 1) {real, imag} */,
  {32'h3f3bfebc, 32'hc018f62d} /* (5, 29, 0) {real, imag} */,
  {32'h3f617fca, 32'hbfbb3e70} /* (5, 28, 31) {real, imag} */,
  {32'h3fcaca16, 32'hc0264b7d} /* (5, 28, 30) {real, imag} */,
  {32'h3f172494, 32'hbf2d0948} /* (5, 28, 29) {real, imag} */,
  {32'h3fed6410, 32'hbfbfcb25} /* (5, 28, 28) {real, imag} */,
  {32'h4052ee49, 32'hbfa9f988} /* (5, 28, 27) {real, imag} */,
  {32'hbfd264b4, 32'hbf5f834a} /* (5, 28, 26) {real, imag} */,
  {32'hbfce88dd, 32'hbff114db} /* (5, 28, 25) {real, imag} */,
  {32'hbe3c6f24, 32'hc06968d9} /* (5, 28, 24) {real, imag} */,
  {32'h3f44635e, 32'hbfc67ffd} /* (5, 28, 23) {real, imag} */,
  {32'hbfabd2dd, 32'h3e1fcad4} /* (5, 28, 22) {real, imag} */,
  {32'hbfb48f46, 32'hc0263ea8} /* (5, 28, 21) {real, imag} */,
  {32'hbfb2e1f1, 32'hc00bc9fa} /* (5, 28, 20) {real, imag} */,
  {32'hc00b04c0, 32'hbf848c65} /* (5, 28, 19) {real, imag} */,
  {32'hc02add5e, 32'h3f2466e0} /* (5, 28, 18) {real, imag} */,
  {32'hc02068b6, 32'h400a1dc2} /* (5, 28, 17) {real, imag} */,
  {32'hc062d24b, 32'h40525abb} /* (5, 28, 16) {real, imag} */,
  {32'hc05bf708, 32'h403643f4} /* (5, 28, 15) {real, imag} */,
  {32'hbf75b00e, 32'h3ffa04ba} /* (5, 28, 14) {real, imag} */,
  {32'hbfc31d9c, 32'h3fb88b75} /* (5, 28, 13) {real, imag} */,
  {32'hbfeae1b2, 32'h3fb7da6a} /* (5, 28, 12) {real, imag} */,
  {32'hbfc9528b, 32'h40898ff2} /* (5, 28, 11) {real, imag} */,
  {32'hbf48390c, 32'hbf39d560} /* (5, 28, 10) {real, imag} */,
  {32'h401bb740, 32'hc08636b8} /* (5, 28, 9) {real, imag} */,
  {32'h401b073e, 32'hc0524066} /* (5, 28, 8) {real, imag} */,
  {32'h3ff5b338, 32'hc00b2f2f} /* (5, 28, 7) {real, imag} */,
  {32'h403877ea, 32'hbfe976f3} /* (5, 28, 6) {real, imag} */,
  {32'h401057ce, 32'hc0559e44} /* (5, 28, 5) {real, imag} */,
  {32'h3f68ac31, 32'hbf9133e2} /* (5, 28, 4) {real, imag} */,
  {32'h3fe66992, 32'hc04547ac} /* (5, 28, 3) {real, imag} */,
  {32'h40853d8c, 32'hc044ef97} /* (5, 28, 2) {real, imag} */,
  {32'h3feaa412, 32'hbfe7bd43} /* (5, 28, 1) {real, imag} */,
  {32'hbe56d964, 32'hbfb0f1cc} /* (5, 28, 0) {real, imag} */,
  {32'h3f7b3a48, 32'hbf6c4fd9} /* (5, 27, 31) {real, imag} */,
  {32'h3f16a2c1, 32'hbfaefa26} /* (5, 27, 30) {real, imag} */,
  {32'hbfe71616, 32'h3f82894f} /* (5, 27, 29) {real, imag} */,
  {32'h40163643, 32'hbedb9452} /* (5, 27, 28) {real, imag} */,
  {32'h406a91b2, 32'h3d0596e0} /* (5, 27, 27) {real, imag} */,
  {32'hbf5a5545, 32'hc00f00c0} /* (5, 27, 26) {real, imag} */,
  {32'hc06ac3c8, 32'hc08fcddc} /* (5, 27, 25) {real, imag} */,
  {32'hbeb959ee, 32'hc08b3c8a} /* (5, 27, 24) {real, imag} */,
  {32'h3fe1e5a8, 32'hbf81f666} /* (5, 27, 23) {real, imag} */,
  {32'h4012a858, 32'hbf8c68d0} /* (5, 27, 22) {real, imag} */,
  {32'hbde9f658, 32'hc08b4374} /* (5, 27, 21) {real, imag} */,
  {32'hbf5e20b8, 32'hbf8cf9cc} /* (5, 27, 20) {real, imag} */,
  {32'hbf7034a0, 32'h3ec8a6a4} /* (5, 27, 19) {real, imag} */,
  {32'hc05ac066, 32'h404d423a} /* (5, 27, 18) {real, imag} */,
  {32'hbfe1e0fe, 32'h4080ad29} /* (5, 27, 17) {real, imag} */,
  {32'h3f25248e, 32'h406f8716} /* (5, 27, 16) {real, imag} */,
  {32'hc015c8a5, 32'h3fe63150} /* (5, 27, 15) {real, imag} */,
  {32'hbf6964c5, 32'hbbe30a80} /* (5, 27, 14) {real, imag} */,
  {32'hbfdcb2f4, 32'h3f90b8b6} /* (5, 27, 13) {real, imag} */,
  {32'hc05790d0, 32'h40449b74} /* (5, 27, 12) {real, imag} */,
  {32'hc01ed7d3, 32'h40a2e0d2} /* (5, 27, 11) {real, imag} */,
  {32'h3c7ee200, 32'hbfca3089} /* (5, 27, 10) {real, imag} */,
  {32'hbfabe7f8, 32'hc09d59cc} /* (5, 27, 9) {real, imag} */,
  {32'h3f7e882e, 32'hc01038d8} /* (5, 27, 8) {real, imag} */,
  {32'h3f9ed8a5, 32'hbfe2430b} /* (5, 27, 7) {real, imag} */,
  {32'h3fd24db8, 32'hbfa1bd2c} /* (5, 27, 6) {real, imag} */,
  {32'hbf42fa43, 32'hc08011a2} /* (5, 27, 5) {real, imag} */,
  {32'hbf68ab9a, 32'hc08a0eb0} /* (5, 27, 4) {real, imag} */,
  {32'h3fe5767e, 32'hc0531c10} /* (5, 27, 3) {real, imag} */,
  {32'h401cb186, 32'hbf7bdf4b} /* (5, 27, 2) {real, imag} */,
  {32'h3fe465d5, 32'hbf993498} /* (5, 27, 1) {real, imag} */,
  {32'h3f86490c, 32'hbf84c6a6} /* (5, 27, 0) {real, imag} */,
  {32'hbdd2ddba, 32'hbf13bff3} /* (5, 26, 31) {real, imag} */,
  {32'hbf05eca5, 32'h3f10cc74} /* (5, 26, 30) {real, imag} */,
  {32'hc01b01ae, 32'h3e35e1cc} /* (5, 26, 29) {real, imag} */,
  {32'hbc8b8d40, 32'hbfa20009} /* (5, 26, 28) {real, imag} */,
  {32'h403404e4, 32'h3ef7dccc} /* (5, 26, 27) {real, imag} */,
  {32'h403f66f5, 32'hc0897228} /* (5, 26, 26) {real, imag} */,
  {32'h3f7fdb84, 32'hc08bb020} /* (5, 26, 25) {real, imag} */,
  {32'h3ffd8e05, 32'hbf645638} /* (5, 26, 24) {real, imag} */,
  {32'h404cc058, 32'hbf350f48} /* (5, 26, 23) {real, imag} */,
  {32'h401c9db9, 32'hbf9d531c} /* (5, 26, 22) {real, imag} */,
  {32'hbfb22e0c, 32'hc03d8ae0} /* (5, 26, 21) {real, imag} */,
  {32'hbfadc356, 32'h3f48670e} /* (5, 26, 20) {real, imag} */,
  {32'hbded7c98, 32'h3ff3ec7e} /* (5, 26, 19) {real, imag} */,
  {32'hbf9d4ea8, 32'h408433c2} /* (5, 26, 18) {real, imag} */,
  {32'hbfd31cbb, 32'h40602168} /* (5, 26, 17) {real, imag} */,
  {32'h3f32119e, 32'h405948c0} /* (5, 26, 16) {real, imag} */,
  {32'hbfb57610, 32'h4017422f} /* (5, 26, 15) {real, imag} */,
  {32'hc00a2265, 32'h4004edc6} /* (5, 26, 14) {real, imag} */,
  {32'hbfcf7d2c, 32'h3fb2f8fa} /* (5, 26, 13) {real, imag} */,
  {32'hc01f66b2, 32'h3f36209d} /* (5, 26, 12) {real, imag} */,
  {32'hc023c0d3, 32'h3ead35ac} /* (5, 26, 11) {real, imag} */,
  {32'h3e04fb38, 32'hc02354b9} /* (5, 26, 10) {real, imag} */,
  {32'h3e706dd8, 32'hbf962cc4} /* (5, 26, 9) {real, imag} */,
  {32'hbe3ec0e2, 32'hbff0647c} /* (5, 26, 8) {real, imag} */,
  {32'h3e84f96a, 32'hc0069af8} /* (5, 26, 7) {real, imag} */,
  {32'h3f88b21e, 32'hbf45c97c} /* (5, 26, 6) {real, imag} */,
  {32'h3eff166c, 32'hc0791ec7} /* (5, 26, 5) {real, imag} */,
  {32'hbc2b3f00, 32'hc0863e82} /* (5, 26, 4) {real, imag} */,
  {32'hbf5a82a3, 32'hbfd7da05} /* (5, 26, 3) {real, imag} */,
  {32'h3f3515cc, 32'hbe57b9d0} /* (5, 26, 2) {real, imag} */,
  {32'h3cb14c80, 32'hbe60c904} /* (5, 26, 1) {real, imag} */,
  {32'hbfb05ca9, 32'hbf22527a} /* (5, 26, 0) {real, imag} */,
  {32'hbea50bbe, 32'hbfdad0b0} /* (5, 25, 31) {real, imag} */,
  {32'h3ed8299e, 32'hc01df9ae} /* (5, 25, 30) {real, imag} */,
  {32'h3e291f1c, 32'hc0405598} /* (5, 25, 29) {real, imag} */,
  {32'h3ebaf7a8, 32'hc0233f50} /* (5, 25, 28) {real, imag} */,
  {32'h3fe35c29, 32'hbfc49e83} /* (5, 25, 27) {real, imag} */,
  {32'h401661bc, 32'hc0179c18} /* (5, 25, 26) {real, imag} */,
  {32'h4033b69a, 32'hbfa5d505} /* (5, 25, 25) {real, imag} */,
  {32'h4099294c, 32'hbfe92160} /* (5, 25, 24) {real, imag} */,
  {32'h4065d8e1, 32'hc0708824} /* (5, 25, 23) {real, imag} */,
  {32'h403252f2, 32'hbfd297c3} /* (5, 25, 22) {real, imag} */,
  {32'h3ef8cc02, 32'hbfe430b1} /* (5, 25, 21) {real, imag} */,
  {32'h3ecf66f0, 32'h403dbfe2} /* (5, 25, 20) {real, imag} */,
  {32'hbede3cb6, 32'h408650cd} /* (5, 25, 19) {real, imag} */,
  {32'hbf73c6bc, 32'h3e67f078} /* (5, 25, 18) {real, imag} */,
  {32'hc06de39c, 32'hbf9f934b} /* (5, 25, 17) {real, imag} */,
  {32'hc03a45dd, 32'hbf102759} /* (5, 25, 16) {real, imag} */,
  {32'hc00ad25a, 32'h3fe32046} /* (5, 25, 15) {real, imag} */,
  {32'hbf20b0be, 32'h40447947} /* (5, 25, 14) {real, imag} */,
  {32'hbf187ffb, 32'h404ff002} /* (5, 25, 13) {real, imag} */,
  {32'hc0536004, 32'h3f1afee6} /* (5, 25, 12) {real, imag} */,
  {32'hc0804fb3, 32'hbf892b52} /* (5, 25, 11) {real, imag} */,
  {32'h3f1e9a15, 32'hc03a9ab2} /* (5, 25, 10) {real, imag} */,
  {32'h3e297358, 32'hbfa22f7e} /* (5, 25, 9) {real, imag} */,
  {32'hbff52631, 32'hc07e4d78} /* (5, 25, 8) {real, imag} */,
  {32'hbfc7c368, 32'hc00ad3f1} /* (5, 25, 7) {real, imag} */,
  {32'h3e0cc50a, 32'h3e9079ce} /* (5, 25, 6) {real, imag} */,
  {32'h3ffa22d5, 32'hbf61c766} /* (5, 25, 5) {real, imag} */,
  {32'h3c5fb040, 32'hc02ce42f} /* (5, 25, 4) {real, imag} */,
  {32'h3f2a00b6, 32'hc007b8f2} /* (5, 25, 3) {real, imag} */,
  {32'h40121e04, 32'hbf71582e} /* (5, 25, 2) {real, imag} */,
  {32'h3d5a7c00, 32'hc028b508} /* (5, 25, 1) {real, imag} */,
  {32'hbff4e120, 32'hbfc0696e} /* (5, 25, 0) {real, imag} */,
  {32'h3f9e26fc, 32'hbfaa045e} /* (5, 24, 31) {real, imag} */,
  {32'h40324540, 32'hbfda1b0c} /* (5, 24, 30) {real, imag} */,
  {32'h40894b38, 32'hc02d4d2c} /* (5, 24, 29) {real, imag} */,
  {32'h409c6304, 32'hc0a3fd18} /* (5, 24, 28) {real, imag} */,
  {32'h40853ceb, 32'hc09bfb37} /* (5, 24, 27) {real, imag} */,
  {32'h4025f578, 32'hc033106b} /* (5, 24, 26) {real, imag} */,
  {32'h401a6100, 32'hbfd5aa58} /* (5, 24, 25) {real, imag} */,
  {32'h4062e0c8, 32'hc03606c8} /* (5, 24, 24) {real, imag} */,
  {32'h4004a277, 32'hc0915d39} /* (5, 24, 23) {real, imag} */,
  {32'h408224ae, 32'hc05779ac} /* (5, 24, 22) {real, imag} */,
  {32'h401338b7, 32'hc0206b7e} /* (5, 24, 21) {real, imag} */,
  {32'h4037f372, 32'h3e7cd9ac} /* (5, 24, 20) {real, imag} */,
  {32'h3e778f74, 32'h4021a59a} /* (5, 24, 19) {real, imag} */,
  {32'hbfe8aec6, 32'hbf91f51a} /* (5, 24, 18) {real, imag} */,
  {32'hc0ceaeea, 32'hbff8ec70} /* (5, 24, 17) {real, imag} */,
  {32'hc0cdd1cc, 32'h3f1dfd22} /* (5, 24, 16) {real, imag} */,
  {32'hc001fdbf, 32'h40966f56} /* (5, 24, 15) {real, imag} */,
  {32'hbedb4bc8, 32'h409c51cc} /* (5, 24, 14) {real, imag} */,
  {32'hc06f6c90, 32'h408a9f2a} /* (5, 24, 13) {real, imag} */,
  {32'hc0cc2a86, 32'h3fecc373} /* (5, 24, 12) {real, imag} */,
  {32'hc054c62e, 32'h4001efea} /* (5, 24, 11) {real, imag} */,
  {32'hbec5ac72, 32'hbf9de423} /* (5, 24, 10) {real, imag} */,
  {32'h3de6bbf0, 32'hc0538ce9} /* (5, 24, 9) {real, imag} */,
  {32'hbfbdf01b, 32'hc0b205be} /* (5, 24, 8) {real, imag} */,
  {32'hbfe27e3d, 32'hc01d7590} /* (5, 24, 7) {real, imag} */,
  {32'hbfd5290a, 32'h3eb95e05} /* (5, 24, 6) {real, imag} */,
  {32'h3f1c528a, 32'h3fcd81ee} /* (5, 24, 5) {real, imag} */,
  {32'hbf58b49a, 32'hbf1d88a0} /* (5, 24, 4) {real, imag} */,
  {32'h3e6aec5e, 32'hbf94ad00} /* (5, 24, 3) {real, imag} */,
  {32'h3f8ae594, 32'hbf890978} /* (5, 24, 2) {real, imag} */,
  {32'h3f874a58, 32'hc059e61c} /* (5, 24, 1) {real, imag} */,
  {32'h3c8847f0, 32'hbfa93d4c} /* (5, 24, 0) {real, imag} */,
  {32'h40064b23, 32'hbf39e86e} /* (5, 23, 31) {real, imag} */,
  {32'h408c7ee6, 32'hbf66ddaa} /* (5, 23, 30) {real, imag} */,
  {32'h40475b7a, 32'hc0393d30} /* (5, 23, 29) {real, imag} */,
  {32'h40529a1d, 32'hc0c003db} /* (5, 23, 28) {real, imag} */,
  {32'h40ae55d3, 32'hc0b725ba} /* (5, 23, 27) {real, imag} */,
  {32'h404b6b4c, 32'hc04a17bc} /* (5, 23, 26) {real, imag} */,
  {32'h40084dca, 32'hbfb459fb} /* (5, 23, 25) {real, imag} */,
  {32'h3f881d44, 32'hc02e06a1} /* (5, 23, 24) {real, imag} */,
  {32'h401e604b, 32'hc08ce065} /* (5, 23, 23) {real, imag} */,
  {32'h40119e70, 32'hc08b3d0d} /* (5, 23, 22) {real, imag} */,
  {32'hbf26c9b8, 32'hbf3866fb} /* (5, 23, 21) {real, imag} */,
  {32'h3f19816c, 32'h3f1847c8} /* (5, 23, 20) {real, imag} */,
  {32'h40027994, 32'h3f9f5d29} /* (5, 23, 19) {real, imag} */,
  {32'h3f679f60, 32'h40134334} /* (5, 23, 18) {real, imag} */,
  {32'hc03fd97e, 32'h4051ad1a} /* (5, 23, 17) {real, imag} */,
  {32'hc028893e, 32'h40321930} /* (5, 23, 16) {real, imag} */,
  {32'hbf2e1a33, 32'h40a53cb6} /* (5, 23, 15) {real, imag} */,
  {32'hc04ca205, 32'h40abdc34} /* (5, 23, 14) {real, imag} */,
  {32'hc0a18c83, 32'h4081bd93} /* (5, 23, 13) {real, imag} */,
  {32'hc06f949a, 32'h40679e6a} /* (5, 23, 12) {real, imag} */,
  {32'hbf5340e3, 32'h3f44e1b2} /* (5, 23, 11) {real, imag} */,
  {32'hbf4a020c, 32'hc017c142} /* (5, 23, 10) {real, imag} */,
  {32'hbe8c3c52, 32'hc07d8856} /* (5, 23, 9) {real, imag} */,
  {32'h3fce7fe9, 32'hc0ad3b93} /* (5, 23, 8) {real, imag} */,
  {32'h3ebfcf5e, 32'hc0835c7e} /* (5, 23, 7) {real, imag} */,
  {32'hbfa346b3, 32'hc0461a3e} /* (5, 23, 6) {real, imag} */,
  {32'hbf5e54e9, 32'hc03e9627} /* (5, 23, 5) {real, imag} */,
  {32'hc00cefaf, 32'h3da93270} /* (5, 23, 4) {real, imag} */,
  {32'h3e0c81a2, 32'h3e207404} /* (5, 23, 3) {real, imag} */,
  {32'h3f4e81df, 32'hbfb9f427} /* (5, 23, 2) {real, imag} */,
  {32'h3e518e70, 32'h3e8c7bbe} /* (5, 23, 1) {real, imag} */,
  {32'h3f8577e5, 32'h3e1d6988} /* (5, 23, 0) {real, imag} */,
  {32'h3fbe1450, 32'hc032c3e6} /* (5, 22, 31) {real, imag} */,
  {32'h402357ba, 32'hc076e3da} /* (5, 22, 30) {real, imag} */,
  {32'h3fa8f815, 32'hc0bd2944} /* (5, 22, 29) {real, imag} */,
  {32'h3f7865aa, 32'hc0a09120} /* (5, 22, 28) {real, imag} */,
  {32'h40364efb, 32'hc07775be} /* (5, 22, 27) {real, imag} */,
  {32'h3fb9fe74, 32'hc0476152} /* (5, 22, 26) {real, imag} */,
  {32'h3fb75e98, 32'hbfa09e06} /* (5, 22, 25) {real, imag} */,
  {32'h3f6c822a, 32'hc0269e8c} /* (5, 22, 24) {real, imag} */,
  {32'h40481868, 32'hc04d140b} /* (5, 22, 23) {real, imag} */,
  {32'h403a02a2, 32'hc049f1e1} /* (5, 22, 22) {real, imag} */,
  {32'hbef73f8c, 32'hbe46df52} /* (5, 22, 21) {real, imag} */,
  {32'hc00119be, 32'h3f59672c} /* (5, 22, 20) {real, imag} */,
  {32'hbf3ebde0, 32'h4005428c} /* (5, 22, 19) {real, imag} */,
  {32'hbe356b48, 32'h40781bea} /* (5, 22, 18) {real, imag} */,
  {32'hc00b200b, 32'h406bd553} /* (5, 22, 17) {real, imag} */,
  {32'hbe975bc6, 32'h3f9589a0} /* (5, 22, 16) {real, imag} */,
  {32'h3ef852cd, 32'h3fafae8a} /* (5, 22, 15) {real, imag} */,
  {32'hbfabdfbb, 32'h3fcd873b} /* (5, 22, 14) {real, imag} */,
  {32'hbf5e04f2, 32'h3ec9e12a} /* (5, 22, 13) {real, imag} */,
  {32'hc009a80b, 32'hbf15f522} /* (5, 22, 12) {real, imag} */,
  {32'hbfad9bc8, 32'hbfb63c12} /* (5, 22, 11) {real, imag} */,
  {32'h3ec6d3a8, 32'hc02cdeaa} /* (5, 22, 10) {real, imag} */,
  {32'h4023f948, 32'hbfd04b04} /* (5, 22, 9) {real, imag} */,
  {32'h409ba3a3, 32'hc06b1e3e} /* (5, 22, 8) {real, imag} */,
  {32'h404138e8, 32'hc0631773} /* (5, 22, 7) {real, imag} */,
  {32'h3ffdd81f, 32'hc051df24} /* (5, 22, 6) {real, imag} */,
  {32'h3f590478, 32'hc06c9183} /* (5, 22, 5) {real, imag} */,
  {32'hbf82ba8e, 32'hbf33b62f} /* (5, 22, 4) {real, imag} */,
  {32'h3d1c3d30, 32'hbf41d6ed} /* (5, 22, 3) {real, imag} */,
  {32'hbf023496, 32'hbf25a06e} /* (5, 22, 2) {real, imag} */,
  {32'h3ee1f0a4, 32'h3f26daa6} /* (5, 22, 1) {real, imag} */,
  {32'h3f748112, 32'hbf423fb0} /* (5, 22, 0) {real, imag} */,
  {32'hbfa417f5, 32'hbf859949} /* (5, 21, 31) {real, imag} */,
  {32'hbf8ce5e8, 32'hc022b9f6} /* (5, 21, 30) {real, imag} */,
  {32'h3ef65c7a, 32'hc06357ec} /* (5, 21, 29) {real, imag} */,
  {32'h3fb8c68a, 32'h3ef9b606} /* (5, 21, 28) {real, imag} */,
  {32'h4012a3ec, 32'hc01831ee} /* (5, 21, 27) {real, imag} */,
  {32'h3f5b9422, 32'hbfebe71c} /* (5, 21, 26) {real, imag} */,
  {32'hbf8ba480, 32'hbeec1d1b} /* (5, 21, 25) {real, imag} */,
  {32'hbf995bd6, 32'hbf5b9ce8} /* (5, 21, 24) {real, imag} */,
  {32'h3e8dab0b, 32'hbf2284e4} /* (5, 21, 23) {real, imag} */,
  {32'h3fc7282c, 32'hbff0abd8} /* (5, 21, 22) {real, imag} */,
  {32'h3e07a1c8, 32'hc005a818} /* (5, 21, 21) {real, imag} */,
  {32'hbf6190a8, 32'h3e073d18} /* (5, 21, 20) {real, imag} */,
  {32'hbf9463c9, 32'h400558cb} /* (5, 21, 19) {real, imag} */,
  {32'h3efa5824, 32'h3f8ad3a3} /* (5, 21, 18) {real, imag} */,
  {32'hbf9b7078, 32'hba8b6a00} /* (5, 21, 17) {real, imag} */,
  {32'hbf09fa4d, 32'hbf5318ea} /* (5, 21, 16) {real, imag} */,
  {32'h3f19a8a0, 32'h3df89c78} /* (5, 21, 15) {real, imag} */,
  {32'h3f88b9ba, 32'h3f7d8e3a} /* (5, 21, 14) {real, imag} */,
  {32'h3f95a7f1, 32'hbf6939f8} /* (5, 21, 13) {real, imag} */,
  {32'h3f0142cc, 32'hbe8166f0} /* (5, 21, 12) {real, imag} */,
  {32'hbf190370, 32'hbec59360} /* (5, 21, 11) {real, imag} */,
  {32'hbfbfaf15, 32'hbf3c2926} /* (5, 21, 10) {real, imag} */,
  {32'hbe7333c6, 32'hc001624d} /* (5, 21, 9) {real, imag} */,
  {32'h409267e3, 32'hbfa20f76} /* (5, 21, 8) {real, imag} */,
  {32'h3ff9ee27, 32'hbfc6d0f0} /* (5, 21, 7) {real, imag} */,
  {32'h4031e47b, 32'hbf90c6a0} /* (5, 21, 6) {real, imag} */,
  {32'h3fea4cd6, 32'h3eb8a38c} /* (5, 21, 5) {real, imag} */,
  {32'h3f727290, 32'hbe8f52ee} /* (5, 21, 4) {real, imag} */,
  {32'h4046c22c, 32'hbfff36e3} /* (5, 21, 3) {real, imag} */,
  {32'h3faecdff, 32'h3fb707e5} /* (5, 21, 2) {real, imag} */,
  {32'h3f70d256, 32'h3fea2d10} /* (5, 21, 1) {real, imag} */,
  {32'h3f35a54c, 32'hbeaf68be} /* (5, 21, 0) {real, imag} */,
  {32'hc005738a, 32'h3fdd2c67} /* (5, 20, 31) {real, imag} */,
  {32'hc0509a6c, 32'h3f78c875} /* (5, 20, 30) {real, imag} */,
  {32'hbff0eeef, 32'hbf1f7a7e} /* (5, 20, 29) {real, imag} */,
  {32'hbda99b78, 32'h40340606} /* (5, 20, 28) {real, imag} */,
  {32'h3f49a0f2, 32'h40068338} /* (5, 20, 27) {real, imag} */,
  {32'hbf8ad6ce, 32'h40369dfb} /* (5, 20, 26) {real, imag} */,
  {32'hc05f89b7, 32'h3f73980e} /* (5, 20, 25) {real, imag} */,
  {32'hbff07ae6, 32'hbee0d208} /* (5, 20, 24) {real, imag} */,
  {32'hbff575db, 32'h403a52d2} /* (5, 20, 23) {real, imag} */,
  {32'hbe89f4d8, 32'h3fa16870} /* (5, 20, 22) {real, imag} */,
  {32'h3f2fe53e, 32'hbef003dc} /* (5, 20, 21) {real, imag} */,
  {32'h3f0d0244, 32'hc0033f3f} /* (5, 20, 20) {real, imag} */,
  {32'h3e28bee8, 32'hbe9123ba} /* (5, 20, 19) {real, imag} */,
  {32'h4056b254, 32'hbebd7fdc} /* (5, 20, 18) {real, imag} */,
  {32'h405cb2f8, 32'hbf0450c1} /* (5, 20, 17) {real, imag} */,
  {32'h3f867684, 32'hc0271159} /* (5, 20, 16) {real, imag} */,
  {32'hc0163712, 32'hbeaee06f} /* (5, 20, 15) {real, imag} */,
  {32'hbf929415, 32'hbf7051e3} /* (5, 20, 14) {real, imag} */,
  {32'hbed5fdb6, 32'hbfacb945} /* (5, 20, 13) {real, imag} */,
  {32'h3f652dc3, 32'hbf8742e9} /* (5, 20, 12) {real, imag} */,
  {32'hbff8a86a, 32'hbfbe3521} /* (5, 20, 11) {real, imag} */,
  {32'hc08ed6b8, 32'h40011ad9} /* (5, 20, 10) {real, imag} */,
  {32'hc059d288, 32'h3fba0c3c} /* (5, 20, 9) {real, imag} */,
  {32'h3f8577ba, 32'h404b2da6} /* (5, 20, 8) {real, imag} */,
  {32'hbf8c3b9d, 32'h4023c44c} /* (5, 20, 7) {real, imag} */,
  {32'hbf129df8, 32'h3fa4dfe0} /* (5, 20, 6) {real, imag} */,
  {32'hbfe04136, 32'h402e4475} /* (5, 20, 5) {real, imag} */,
  {32'hbff70ed4, 32'h3f998cbe} /* (5, 20, 4) {real, imag} */,
  {32'hbecc63b8, 32'hbecf7d98} /* (5, 20, 3) {real, imag} */,
  {32'h3dc33938, 32'h403ee305} /* (5, 20, 2) {real, imag} */,
  {32'h3f4ebf28, 32'h40897aef} /* (5, 20, 1) {real, imag} */,
  {32'hbe1886f6, 32'h400a84e2} /* (5, 20, 0) {real, imag} */,
  {32'h3fbb4fb1, 32'h3f769471} /* (5, 19, 31) {real, imag} */,
  {32'h3fbb565f, 32'h3f8ba292} /* (5, 19, 30) {real, imag} */,
  {32'h3f3b7331, 32'hbf010fa9} /* (5, 19, 29) {real, imag} */,
  {32'h3eced446, 32'h3f333b48} /* (5, 19, 28) {real, imag} */,
  {32'h3dec14b8, 32'h40312b0f} /* (5, 19, 27) {real, imag} */,
  {32'hbf8a2f38, 32'h401969dc} /* (5, 19, 26) {real, imag} */,
  {32'hc012c232, 32'hbdf75020} /* (5, 19, 25) {real, imag} */,
  {32'hbfe2b922, 32'hbe722c30} /* (5, 19, 24) {real, imag} */,
  {32'hc045706a, 32'h3ff525cd} /* (5, 19, 23) {real, imag} */,
  {32'hbfc06eea, 32'h4007cac6} /* (5, 19, 22) {real, imag} */,
  {32'hbd5d6be4, 32'hbe6d8418} /* (5, 19, 21) {real, imag} */,
  {32'h3f8b50ee, 32'hc05b5527} /* (5, 19, 20) {real, imag} */,
  {32'h4023c4d4, 32'hc066beb8} /* (5, 19, 19) {real, imag} */,
  {32'h40638130, 32'h3e27bbb8} /* (5, 19, 18) {real, imag} */,
  {32'h402f2ce1, 32'hbf100b96} /* (5, 19, 17) {real, imag} */,
  {32'h3ff05b23, 32'hc00f2f0a} /* (5, 19, 16) {real, imag} */,
  {32'h3fa251ed, 32'hbefc2062} /* (5, 19, 15) {real, imag} */,
  {32'h3f339bb8, 32'hc0001416} /* (5, 19, 14) {real, imag} */,
  {32'h3faa6bad, 32'hbfaeff5d} /* (5, 19, 13) {real, imag} */,
  {32'h3ff5ca72, 32'hbd5eb330} /* (5, 19, 12) {real, imag} */,
  {32'h3ef4a9f2, 32'hbfc93916} /* (5, 19, 11) {real, imag} */,
  {32'hc02d2ff4, 32'h3e1e77d0} /* (5, 19, 10) {real, imag} */,
  {32'hbf2904d7, 32'h4024ef1a} /* (5, 19, 9) {real, imag} */,
  {32'h3f7bc0e8, 32'h4080257c} /* (5, 19, 8) {real, imag} */,
  {32'h3ee6d872, 32'h405cf702} /* (5, 19, 7) {real, imag} */,
  {32'hbe387130, 32'h402ed1ce} /* (5, 19, 6) {real, imag} */,
  {32'hc019b1b2, 32'h405d4a46} /* (5, 19, 5) {real, imag} */,
  {32'hc00699f0, 32'h40327d44} /* (5, 19, 4) {real, imag} */,
  {32'hc00f8d08, 32'h3f344ca6} /* (5, 19, 3) {real, imag} */,
  {32'hbf4d258d, 32'h3fd2445f} /* (5, 19, 2) {real, imag} */,
  {32'h3e386d1c, 32'h3fdda522} /* (5, 19, 1) {real, imag} */,
  {32'h3f4de2d8, 32'h3f158f0c} /* (5, 19, 0) {real, imag} */,
  {32'h3fe88a7c, 32'h400b44a8} /* (5, 18, 31) {real, imag} */,
  {32'h3f796d52, 32'h406dd126} /* (5, 18, 30) {real, imag} */,
  {32'hbfaf6c12, 32'h3fdce0da} /* (5, 18, 29) {real, imag} */,
  {32'hbf464d60, 32'hbf4ba29a} /* (5, 18, 28) {real, imag} */,
  {32'h3e92acd8, 32'hbef036fa} /* (5, 18, 27) {real, imag} */,
  {32'hbe8635e4, 32'hbeac63e6} /* (5, 18, 26) {real, imag} */,
  {32'hbf41e133, 32'h3fe44e5d} /* (5, 18, 25) {real, imag} */,
  {32'hc0698f6d, 32'h40455029} /* (5, 18, 24) {real, imag} */,
  {32'hc059551a, 32'h4076ba20} /* (5, 18, 23) {real, imag} */,
  {32'hbf4bd4f2, 32'h40820970} /* (5, 18, 22) {real, imag} */,
  {32'hbeac6eeb, 32'h3fbeac36} /* (5, 18, 21) {real, imag} */,
  {32'h40032110, 32'hc00dd637} /* (5, 18, 20) {real, imag} */,
  {32'h404eb98c, 32'hc032ad68} /* (5, 18, 19) {real, imag} */,
  {32'h4019e04b, 32'h3f290432} /* (5, 18, 18) {real, imag} */,
  {32'h403dceba, 32'hbfcce1df} /* (5, 18, 17) {real, imag} */,
  {32'h3f707793, 32'hc03db9bb} /* (5, 18, 16) {real, imag} */,
  {32'h4016ed38, 32'hbfb51203} /* (5, 18, 15) {real, imag} */,
  {32'h403db41a, 32'hc05a29dc} /* (5, 18, 14) {real, imag} */,
  {32'h3fe9d642, 32'hc03a1522} /* (5, 18, 13) {real, imag} */,
  {32'h3cfabac0, 32'hbf3341f2} /* (5, 18, 12) {real, imag} */,
  {32'h405e3b33, 32'hbfe0db91} /* (5, 18, 11) {real, imag} */,
  {32'h3fce40ca, 32'hbe18a498} /* (5, 18, 10) {real, imag} */,
  {32'hbf796e74, 32'h400e9cad} /* (5, 18, 9) {real, imag} */,
  {32'hbfa0d485, 32'h40044d00} /* (5, 18, 8) {real, imag} */,
  {32'h3f94e65a, 32'h3eae6540} /* (5, 18, 7) {real, imag} */,
  {32'hbe2f1e68, 32'h40817894} /* (5, 18, 6) {real, imag} */,
  {32'hbf3cbfd6, 32'h40730970} /* (5, 18, 5) {real, imag} */,
  {32'hbfb02bd0, 32'h403bbba2} /* (5, 18, 4) {real, imag} */,
  {32'hbf488698, 32'h402f7dbe} /* (5, 18, 3) {real, imag} */,
  {32'hbe0eb2e8, 32'h3ecf281d} /* (5, 18, 2) {real, imag} */,
  {32'hbe7d41b0, 32'h40404ac0} /* (5, 18, 1) {real, imag} */,
  {32'h4012ac98, 32'h40057180} /* (5, 18, 0) {real, imag} */,
  {32'hbf446644, 32'h40465cb0} /* (5, 17, 31) {real, imag} */,
  {32'hbf03de94, 32'h40cb6b4c} /* (5, 17, 30) {real, imag} */,
  {32'hbf330a48, 32'h406061d5} /* (5, 17, 29) {real, imag} */,
  {32'h3f8f1b4a, 32'h3eb49618} /* (5, 17, 28) {real, imag} */,
  {32'h405e7b89, 32'h3fd8f43e} /* (5, 17, 27) {real, imag} */,
  {32'h40387b07, 32'h3f03272b} /* (5, 17, 26) {real, imag} */,
  {32'hbf10248c, 32'h406072ec} /* (5, 17, 25) {real, imag} */,
  {32'hc03fe108, 32'h40a8b77e} /* (5, 17, 24) {real, imag} */,
  {32'hbfd9bdf4, 32'h40b297fc} /* (5, 17, 23) {real, imag} */,
  {32'hbf923a3c, 32'h40311d7e} /* (5, 17, 22) {real, imag} */,
  {32'h3f004ebe, 32'h3f7bf433} /* (5, 17, 21) {real, imag} */,
  {32'h40452bb7, 32'hbf577e59} /* (5, 17, 20) {real, imag} */,
  {32'h4059a834, 32'hbf843a5f} /* (5, 17, 19) {real, imag} */,
  {32'h4032a0c8, 32'h3f9d1bf9} /* (5, 17, 18) {real, imag} */,
  {32'h402ea3dc, 32'hbf098c1c} /* (5, 17, 17) {real, imag} */,
  {32'h400e8728, 32'hbf834455} /* (5, 17, 16) {real, imag} */,
  {32'h4075f217, 32'hbf5334fc} /* (5, 17, 15) {real, imag} */,
  {32'h40592463, 32'hbef18da8} /* (5, 17, 14) {real, imag} */,
  {32'h402625c5, 32'hbe4018d4} /* (5, 17, 13) {real, imag} */,
  {32'h4018711e, 32'hbf882328} /* (5, 17, 12) {real, imag} */,
  {32'h401d0750, 32'hbee486da} /* (5, 17, 11) {real, imag} */,
  {32'h3f8dc9aa, 32'h4009aceb} /* (5, 17, 10) {real, imag} */,
  {32'hbfda1290, 32'h4023919c} /* (5, 17, 9) {real, imag} */,
  {32'hbe1c8ef0, 32'h40445b01} /* (5, 17, 8) {real, imag} */,
  {32'h3f9f7d73, 32'h3fc18fea} /* (5, 17, 7) {real, imag} */,
  {32'h3f97b6d1, 32'h4006126e} /* (5, 17, 6) {real, imag} */,
  {32'hc009e36e, 32'h402d1cc5} /* (5, 17, 5) {real, imag} */,
  {32'hc03c95e0, 32'h40186d14} /* (5, 17, 4) {real, imag} */,
  {32'hbf980918, 32'h40295c2b} /* (5, 17, 3) {real, imag} */,
  {32'h3f437e26, 32'h401fd304} /* (5, 17, 2) {real, imag} */,
  {32'hbf13ff0c, 32'h4007d9c0} /* (5, 17, 1) {real, imag} */,
  {32'hbec7ada7, 32'h40033e7e} /* (5, 17, 0) {real, imag} */,
  {32'hbf53f77d, 32'h3f905cdc} /* (5, 16, 31) {real, imag} */,
  {32'h3d86e010, 32'h408da47a} /* (5, 16, 30) {real, imag} */,
  {32'hbea62352, 32'h40690f5b} /* (5, 16, 29) {real, imag} */,
  {32'h4057071b, 32'h3ff755cd} /* (5, 16, 28) {real, imag} */,
  {32'h403b80fc, 32'h4072ad82} /* (5, 16, 27) {real, imag} */,
  {32'h3ef3df2a, 32'h401a3369} /* (5, 16, 26) {real, imag} */,
  {32'hbf54f634, 32'h407eafb1} /* (5, 16, 25) {real, imag} */,
  {32'hbf4db1d2, 32'h4072e79a} /* (5, 16, 24) {real, imag} */,
  {32'hc023e7ec, 32'h40ba1ad0} /* (5, 16, 23) {real, imag} */,
  {32'hc08ea251, 32'h408493a2} /* (5, 16, 22) {real, imag} */,
  {32'h3e4ab06c, 32'h3fc08314} /* (5, 16, 21) {real, imag} */,
  {32'h406720cb, 32'h3dc651d0} /* (5, 16, 20) {real, imag} */,
  {32'h406fca26, 32'hbf87d4c8} /* (5, 16, 19) {real, imag} */,
  {32'h40750b28, 32'hc00a58ec} /* (5, 16, 18) {real, imag} */,
  {32'h4027d8be, 32'hc0582f33} /* (5, 16, 17) {real, imag} */,
  {32'h4015ee10, 32'hc0603913} /* (5, 16, 16) {real, imag} */,
  {32'h403b4954, 32'hc029133e} /* (5, 16, 15) {real, imag} */,
  {32'h3fab35ab, 32'h3e8130cc} /* (5, 16, 14) {real, imag} */,
  {32'h40059482, 32'hbf715223} /* (5, 16, 13) {real, imag} */,
  {32'h408c51ca, 32'hc06dfdcc} /* (5, 16, 12) {real, imag} */,
  {32'h40223ac0, 32'hc03c5606} /* (5, 16, 11) {real, imag} */,
  {32'h400db6ac, 32'hbf6cbcb5} /* (5, 16, 10) {real, imag} */,
  {32'h3f9065c4, 32'h3e979d3c} /* (5, 16, 9) {real, imag} */,
  {32'h40255cae, 32'h40597a33} /* (5, 16, 8) {real, imag} */,
  {32'h3ff6890a, 32'h407819f9} /* (5, 16, 7) {real, imag} */,
  {32'h40559ac4, 32'h4021ab18} /* (5, 16, 6) {real, imag} */,
  {32'hbf116cc8, 32'h401d01b8} /* (5, 16, 5) {real, imag} */,
  {32'hbfd38f38, 32'h4020ae06} /* (5, 16, 4) {real, imag} */,
  {32'hbff0af78, 32'hbd407a40} /* (5, 16, 3) {real, imag} */,
  {32'hc001399a, 32'h3ff54de2} /* (5, 16, 2) {real, imag} */,
  {32'hc03cbf06, 32'h3fe9caf9} /* (5, 16, 1) {real, imag} */,
  {32'hc01599e5, 32'h3f038e1b} /* (5, 16, 0) {real, imag} */,
  {32'h3e90d4a0, 32'h3f6686b1} /* (5, 15, 31) {real, imag} */,
  {32'h3f18dafe, 32'h40050d3b} /* (5, 15, 30) {real, imag} */,
  {32'hc00cc3e6, 32'h402388d7} /* (5, 15, 29) {real, imag} */,
  {32'hc00c511b, 32'h3ff7402e} /* (5, 15, 28) {real, imag} */,
  {32'hc05b390e, 32'h409a9335} /* (5, 15, 27) {real, imag} */,
  {32'hbfcd4f2e, 32'h40a1e643} /* (5, 15, 26) {real, imag} */,
  {32'hbfb53348, 32'h402de67a} /* (5, 15, 25) {real, imag} */,
  {32'h3f2a482d, 32'h403b8f75} /* (5, 15, 24) {real, imag} */,
  {32'hc053374e, 32'h40d12b50} /* (5, 15, 23) {real, imag} */,
  {32'hc0a4c4e5, 32'h40d4f11e} /* (5, 15, 22) {real, imag} */,
  {32'hbf870453, 32'h40232ecc} /* (5, 15, 21) {real, imag} */,
  {32'h4023209e, 32'h3f56e7aa} /* (5, 15, 20) {real, imag} */,
  {32'h3f482a42, 32'hbf7b340d} /* (5, 15, 19) {real, imag} */,
  {32'hbea3b68e, 32'hc05473d9} /* (5, 15, 18) {real, imag} */,
  {32'h3ecfca9b, 32'hc08b1283} /* (5, 15, 17) {real, imag} */,
  {32'h3f053c2c, 32'hc088fa60} /* (5, 15, 16) {real, imag} */,
  {32'hbf10526a, 32'hc053386a} /* (5, 15, 15) {real, imag} */,
  {32'hbf90ca0e, 32'hc018f6b0} /* (5, 15, 14) {real, imag} */,
  {32'hbecef88e, 32'hc09267a6} /* (5, 15, 13) {real, imag} */,
  {32'h3e3dfa5c, 32'hc08be1ab} /* (5, 15, 12) {real, imag} */,
  {32'h3d4cafc0, 32'hc051aeb7} /* (5, 15, 11) {real, imag} */,
  {32'h3d409bc0, 32'h3ea94dc4} /* (5, 15, 10) {real, imag} */,
  {32'hbe7c6070, 32'h3fd515b1} /* (5, 15, 9) {real, imag} */,
  {32'h3f8a1fa8, 32'h3fffaf7e} /* (5, 15, 8) {real, imag} */,
  {32'h3f41da06, 32'h402bbbec} /* (5, 15, 7) {real, imag} */,
  {32'h3faccaaa, 32'h404917a7} /* (5, 15, 6) {real, imag} */,
  {32'h3fef859e, 32'h3f89d848} /* (5, 15, 5) {real, imag} */,
  {32'hbe6b2dc4, 32'hbf0b332c} /* (5, 15, 4) {real, imag} */,
  {32'hc02e6464, 32'hbedc6ea0} /* (5, 15, 3) {real, imag} */,
  {32'hc072b1c9, 32'h3f56cf68} /* (5, 15, 2) {real, imag} */,
  {32'hc088c7fe, 32'h3fe6b1cb} /* (5, 15, 1) {real, imag} */,
  {32'hc04bb62c, 32'h3fccaf35} /* (5, 15, 0) {real, imag} */,
  {32'hbf657fe2, 32'h3ee28506} /* (5, 14, 31) {real, imag} */,
  {32'hbf409042, 32'hbf8bff6c} /* (5, 14, 30) {real, imag} */,
  {32'hbffccc18, 32'h3f85fd66} /* (5, 14, 29) {real, imag} */,
  {32'hc014f7a0, 32'h40707842} /* (5, 14, 28) {real, imag} */,
  {32'hc0498304, 32'h4086dc13} /* (5, 14, 27) {real, imag} */,
  {32'hbfa4f4f1, 32'h3fea5e8d} /* (5, 14, 26) {real, imag} */,
  {32'hbe576e20, 32'h3fb0f818} /* (5, 14, 25) {real, imag} */,
  {32'h3ea315ae, 32'h3ff84344} /* (5, 14, 24) {real, imag} */,
  {32'hc07ed662, 32'h40998f6a} /* (5, 14, 23) {real, imag} */,
  {32'hc086026c, 32'h409d3e6c} /* (5, 14, 22) {real, imag} */,
  {32'hbed32604, 32'h3fc5e22e} /* (5, 14, 21) {real, imag} */,
  {32'h3fb24982, 32'hbec63c70} /* (5, 14, 20) {real, imag} */,
  {32'h3f810e03, 32'hc0312a82} /* (5, 14, 19) {real, imag} */,
  {32'hbf4358be, 32'hc05e69fb} /* (5, 14, 18) {real, imag} */,
  {32'hbff7c78e, 32'hc065c2ce} /* (5, 14, 17) {real, imag} */,
  {32'hbe90f1a6, 32'hc02c5b10} /* (5, 14, 16) {real, imag} */,
  {32'hbf06b22f, 32'hbfc59d6a} /* (5, 14, 15) {real, imag} */,
  {32'hc01a4480, 32'hbff7ac9a} /* (5, 14, 14) {real, imag} */,
  {32'hbfe4a077, 32'hc07d9c84} /* (5, 14, 13) {real, imag} */,
  {32'hbf5c8970, 32'hbf999af9} /* (5, 14, 12) {real, imag} */,
  {32'hbfa346f1, 32'hbf23be34} /* (5, 14, 11) {real, imag} */,
  {32'hc082f4df, 32'h3e4d236c} /* (5, 14, 10) {real, imag} */,
  {32'hc001dfa6, 32'h40225830} /* (5, 14, 9) {real, imag} */,
  {32'hbf8ac0cd, 32'h3fdb4ab2} /* (5, 14, 8) {real, imag} */,
  {32'hc0632cb0, 32'h4013cc22} /* (5, 14, 7) {real, imag} */,
  {32'hbfe9d608, 32'h3fa2217a} /* (5, 14, 6) {real, imag} */,
  {32'h3ea7d384, 32'hbf0213d0} /* (5, 14, 5) {real, imag} */,
  {32'hbfc3f4aa, 32'h3f25a1d7} /* (5, 14, 4) {real, imag} */,
  {32'hbfdc4cd5, 32'h3f2aeb74} /* (5, 14, 3) {real, imag} */,
  {32'hc031a250, 32'h3e2559dc} /* (5, 14, 2) {real, imag} */,
  {32'hc084228f, 32'h3fbcf976} /* (5, 14, 1) {real, imag} */,
  {32'hc05ea6ad, 32'h3f3c7d7d} /* (5, 14, 0) {real, imag} */,
  {32'hbf9a4d9b, 32'h3c7cbce0} /* (5, 13, 31) {real, imag} */,
  {32'hc01e0336, 32'hbf891e5a} /* (5, 13, 30) {real, imag} */,
  {32'hc05aabe4, 32'h3ee63f98} /* (5, 13, 29) {real, imag} */,
  {32'hbfb97817, 32'h40248ca0} /* (5, 13, 28) {real, imag} */,
  {32'hbf1902a8, 32'h3fc9db73} /* (5, 13, 27) {real, imag} */,
  {32'hbf23fb22, 32'hbeb3f918} /* (5, 13, 26) {real, imag} */,
  {32'hbee57b84, 32'hbe270410} /* (5, 13, 25) {real, imag} */,
  {32'hbfeb6cc6, 32'hbe88c408} /* (5, 13, 24) {real, imag} */,
  {32'hc0210c00, 32'h3ee2c3a0} /* (5, 13, 23) {real, imag} */,
  {32'hc0707a3e, 32'h3f698f56} /* (5, 13, 22) {real, imag} */,
  {32'hbfc23e05, 32'h3fd99f2a} /* (5, 13, 21) {real, imag} */,
  {32'h3efc557c, 32'hbfefe0be} /* (5, 13, 20) {real, imag} */,
  {32'h3fda560f, 32'hc0079492} /* (5, 13, 19) {real, imag} */,
  {32'h3f80d20b, 32'hc04a245c} /* (5, 13, 18) {real, imag} */,
  {32'h3d8822c0, 32'hc03ec888} /* (5, 13, 17) {real, imag} */,
  {32'hbfa1664a, 32'hbf6d09f0} /* (5, 13, 16) {real, imag} */,
  {32'hbf427134, 32'hbfa2e816} /* (5, 13, 15) {real, imag} */,
  {32'hbfa5526f, 32'hbfbea2b1} /* (5, 13, 14) {real, imag} */,
  {32'hbfc25eac, 32'hc009a635} /* (5, 13, 13) {real, imag} */,
  {32'hbf30a732, 32'hbf9cdb18} /* (5, 13, 12) {real, imag} */,
  {32'h3e9f50d2, 32'h3ef35bc0} /* (5, 13, 11) {real, imag} */,
  {32'hc0126ece, 32'h400e2688} /* (5, 13, 10) {real, imag} */,
  {32'hc02f00aa, 32'h4020652e} /* (5, 13, 9) {real, imag} */,
  {32'hbf53a7bc, 32'h3d194a10} /* (5, 13, 8) {real, imag} */,
  {32'hc05b3a57, 32'h40144e05} /* (5, 13, 7) {real, imag} */,
  {32'hc0176532, 32'h40083495} /* (5, 13, 6) {real, imag} */,
  {32'hbe04c35e, 32'h3ecc6840} /* (5, 13, 5) {real, imag} */,
  {32'hbf455ed5, 32'h3f6bed12} /* (5, 13, 4) {real, imag} */,
  {32'hbfd9f92c, 32'h40077a71} /* (5, 13, 3) {real, imag} */,
  {32'hc0352ffa, 32'h3fbd4e08} /* (5, 13, 2) {real, imag} */,
  {32'hc05a6a38, 32'h3ece06e4} /* (5, 13, 1) {real, imag} */,
  {32'hbf6dd414, 32'h3f0fab08} /* (5, 13, 0) {real, imag} */,
  {32'hbf5ca718, 32'hbcf85c60} /* (5, 12, 31) {real, imag} */,
  {32'hbfaecb5e, 32'h40011c2c} /* (5, 12, 30) {real, imag} */,
  {32'hc09b5b24, 32'h405c64d9} /* (5, 12, 29) {real, imag} */,
  {32'hc077e169, 32'h407fd708} /* (5, 12, 28) {real, imag} */,
  {32'hbf35fb86, 32'h4003e6a6} /* (5, 12, 27) {real, imag} */,
  {32'hbf77a4ce, 32'h404d256e} /* (5, 12, 26) {real, imag} */,
  {32'hc0325b6c, 32'h407cb926} /* (5, 12, 25) {real, imag} */,
  {32'hc07fa9f3, 32'hbe333b24} /* (5, 12, 24) {real, imag} */,
  {32'hc007bcc2, 32'hc023f987} /* (5, 12, 23) {real, imag} */,
  {32'hbfdd7493, 32'hbf315fca} /* (5, 12, 22) {real, imag} */,
  {32'h3f65c185, 32'hbf89f2d5} /* (5, 12, 21) {real, imag} */,
  {32'h3f85d2d0, 32'hc0494517} /* (5, 12, 20) {real, imag} */,
  {32'h3f07f3c2, 32'hc0657be0} /* (5, 12, 19) {real, imag} */,
  {32'h3fc20064, 32'hc02550e6} /* (5, 12, 18) {real, imag} */,
  {32'h3ecdf280, 32'hc031a804} /* (5, 12, 17) {real, imag} */,
  {32'hbe885e2f, 32'hbf5ffd18} /* (5, 12, 16) {real, imag} */,
  {32'h3fa9afd8, 32'hc00fc2a0} /* (5, 12, 15) {real, imag} */,
  {32'hbf62b597, 32'hbe845612} /* (5, 12, 14) {real, imag} */,
  {32'hbf56c4a9, 32'hbfa18e78} /* (5, 12, 13) {real, imag} */,
  {32'h4007f2cc, 32'hbfeabd96} /* (5, 12, 12) {real, imag} */,
  {32'h3fc8f960, 32'hc026b8d2} /* (5, 12, 11) {real, imag} */,
  {32'hbf3d9ea4, 32'h3fc4002c} /* (5, 12, 10) {real, imag} */,
  {32'hbfc424e5, 32'h401f0bb9} /* (5, 12, 9) {real, imag} */,
  {32'hbf86498d, 32'h3f8f24cc} /* (5, 12, 8) {real, imag} */,
  {32'hbfe93eb3, 32'h3fdafba3} /* (5, 12, 7) {real, imag} */,
  {32'hc07253ff, 32'h3fdb3cfd} /* (5, 12, 6) {real, imag} */,
  {32'hc00fadc6, 32'h3ebb955a} /* (5, 12, 5) {real, imag} */,
  {32'hbf6854d0, 32'hbcabce60} /* (5, 12, 4) {real, imag} */,
  {32'hbfea8ac6, 32'h401ef62c} /* (5, 12, 3) {real, imag} */,
  {32'hc01e4354, 32'h40351a5e} /* (5, 12, 2) {real, imag} */,
  {32'hc0183a94, 32'h400aceb9} /* (5, 12, 1) {real, imag} */,
  {32'hbe8c0139, 32'h3f62d5f7} /* (5, 12, 0) {real, imag} */,
  {32'h3e2a4df8, 32'hbfb14ce4} /* (5, 11, 31) {real, imag} */,
  {32'hbf8178f4, 32'h3e2c6b60} /* (5, 11, 30) {real, imag} */,
  {32'hc0620fc2, 32'h3fd4309f} /* (5, 11, 29) {real, imag} */,
  {32'hc02b2d63, 32'h405ec191} /* (5, 11, 28) {real, imag} */,
  {32'hbf7d8d83, 32'h3fd4325c} /* (5, 11, 27) {real, imag} */,
  {32'hbfe1123f, 32'h4071f1b5} /* (5, 11, 26) {real, imag} */,
  {32'hbf9d7efa, 32'h4073d0a4} /* (5, 11, 25) {real, imag} */,
  {32'hbf26f034, 32'h3f32e83a} /* (5, 11, 24) {real, imag} */,
  {32'hbca33c00, 32'h3f8bf648} /* (5, 11, 23) {real, imag} */,
  {32'h3ea488d1, 32'h3fab6a0c} /* (5, 11, 22) {real, imag} */,
  {32'h3f94d79c, 32'hbdbdf9e8} /* (5, 11, 21) {real, imag} */,
  {32'h400805e8, 32'hbf675a99} /* (5, 11, 20) {real, imag} */,
  {32'h3f943084, 32'hbfddaa43} /* (5, 11, 19) {real, imag} */,
  {32'hbe1795ca, 32'hc0008b3a} /* (5, 11, 18) {real, imag} */,
  {32'hbf159bea, 32'hc0070207} /* (5, 11, 17) {real, imag} */,
  {32'h3f7a05be, 32'h3f211bb9} /* (5, 11, 16) {real, imag} */,
  {32'h3faf0478, 32'hbf63ec98} /* (5, 11, 15) {real, imag} */,
  {32'hbf568694, 32'hbf09d171} /* (5, 11, 14) {real, imag} */,
  {32'hbeddf32c, 32'hc02451d5} /* (5, 11, 13) {real, imag} */,
  {32'h404a1a9c, 32'hbf186d7a} /* (5, 11, 12) {real, imag} */,
  {32'h4012ed98, 32'hbe1cfd38} /* (5, 11, 11) {real, imag} */,
  {32'hbfa0cced, 32'h3fa041ea} /* (5, 11, 10) {real, imag} */,
  {32'hc0915c95, 32'h3f2bee3d} /* (5, 11, 9) {real, imag} */,
  {32'hc06a6ed8, 32'h3f079964} /* (5, 11, 8) {real, imag} */,
  {32'hbf4aef1a, 32'h3fb5c122} /* (5, 11, 7) {real, imag} */,
  {32'hc0686e7b, 32'h3fc3e3c3} /* (5, 11, 6) {real, imag} */,
  {32'hc0a3df53, 32'h3f86813e} /* (5, 11, 5) {real, imag} */,
  {32'hc05f7946, 32'hbfdf17e4} /* (5, 11, 4) {real, imag} */,
  {32'hbfb4a5ad, 32'hbfdabaed} /* (5, 11, 3) {real, imag} */,
  {32'h3e362754, 32'h40168150} /* (5, 11, 2) {real, imag} */,
  {32'hbfa83912, 32'h409e8267} /* (5, 11, 1) {real, imag} */,
  {32'hbfa5cc70, 32'h3fb60756} /* (5, 11, 0) {real, imag} */,
  {32'h3fff1d42, 32'hbfc3c34a} /* (5, 10, 31) {real, imag} */,
  {32'h3fb352a7, 32'hc00685ce} /* (5, 10, 30) {real, imag} */,
  {32'hbf363150, 32'hc07bf4ba} /* (5, 10, 29) {real, imag} */,
  {32'h3eab7364, 32'hbfeaff6e} /* (5, 10, 28) {real, imag} */,
  {32'hbf5f86c0, 32'hbf74be41} /* (5, 10, 27) {real, imag} */,
  {32'hbf95f683, 32'h3ed323dd} /* (5, 10, 26) {real, imag} */,
  {32'hbfb7bd86, 32'h3eee0d30} /* (5, 10, 25) {real, imag} */,
  {32'h3eb05932, 32'hbfc3ecca} /* (5, 10, 24) {real, imag} */,
  {32'h3f4cc386, 32'hbf9fa0ea} /* (5, 10, 23) {real, imag} */,
  {32'hbf884e50, 32'hbffdf89a} /* (5, 10, 22) {real, imag} */,
  {32'h38390000, 32'hbfcf814c} /* (5, 10, 21) {real, imag} */,
  {32'h3f846a13, 32'h3e818338} /* (5, 10, 20) {real, imag} */,
  {32'h3f41ef02, 32'h3ff77068} /* (5, 10, 19) {real, imag} */,
  {32'hbf2ba190, 32'h3f9b5b86} /* (5, 10, 18) {real, imag} */,
  {32'hbf3f1bbf, 32'h400e30ba} /* (5, 10, 17) {real, imag} */,
  {32'hbf6a34da, 32'h4023a703} /* (5, 10, 16) {real, imag} */,
  {32'hbe81f0c2, 32'h40246ac6} /* (5, 10, 15) {real, imag} */,
  {32'h3dc98654, 32'h3fef8038} /* (5, 10, 14) {real, imag} */,
  {32'hbf7fd2e2, 32'h3f14f2da} /* (5, 10, 13) {real, imag} */,
  {32'hbe5e2ba5, 32'h404702d8} /* (5, 10, 12) {real, imag} */,
  {32'hc0169799, 32'h408b1fe6} /* (5, 10, 11) {real, imag} */,
  {32'hbf653144, 32'hbf0f24ac} /* (5, 10, 10) {real, imag} */,
  {32'hc0183e08, 32'hbf8db5d2} /* (5, 10, 9) {real, imag} */,
  {32'hbf2acced, 32'hbfb46482} /* (5, 10, 8) {real, imag} */,
  {32'h3f91c5b8, 32'hbedef88c} /* (5, 10, 7) {real, imag} */,
  {32'hbfdd1f58, 32'hbf76bc62} /* (5, 10, 6) {real, imag} */,
  {32'hc040bd78, 32'hbdff65c0} /* (5, 10, 5) {real, imag} */,
  {32'hbed8cda8, 32'hc0004d32} /* (5, 10, 4) {real, imag} */,
  {32'h3fb03af4, 32'hc0628870} /* (5, 10, 3) {real, imag} */,
  {32'h3f89f141, 32'hbfdfff96} /* (5, 10, 2) {real, imag} */,
  {32'h3f4ee5f0, 32'hbdec6528} /* (5, 10, 1) {real, imag} */,
  {32'h3eb82210, 32'hbfc0e50c} /* (5, 10, 0) {real, imag} */,
  {32'h3fd6917e, 32'hbfba1e0c} /* (5, 9, 31) {real, imag} */,
  {32'h40385302, 32'hc033cd8c} /* (5, 9, 30) {real, imag} */,
  {32'hbf1fdc26, 32'hc08ef262} /* (5, 9, 29) {real, imag} */,
  {32'hbfd3c30a, 32'hc0656c52} /* (5, 9, 28) {real, imag} */,
  {32'hbe36a130, 32'hc0307e18} /* (5, 9, 27) {real, imag} */,
  {32'h3ed064ea, 32'hbfbfc08e} /* (5, 9, 26) {real, imag} */,
  {32'h3e260864, 32'hc00f08f5} /* (5, 9, 25) {real, imag} */,
  {32'h3fd7d0af, 32'hc089fc4e} /* (5, 9, 24) {real, imag} */,
  {32'h3fcccbed, 32'hbf7ac47c} /* (5, 9, 23) {real, imag} */,
  {32'h3ff77d28, 32'hc0090ba4} /* (5, 9, 22) {real, imag} */,
  {32'h40263963, 32'hbff990dc} /* (5, 9, 21) {real, imag} */,
  {32'h3db09e60, 32'h3e9ceb20} /* (5, 9, 20) {real, imag} */,
  {32'hbf452f04, 32'h3ffdffca} /* (5, 9, 19) {real, imag} */,
  {32'hbfd2b4e7, 32'h40bc5480} /* (5, 9, 18) {real, imag} */,
  {32'hc01b3299, 32'h40ade52e} /* (5, 9, 17) {real, imag} */,
  {32'hc019138e, 32'h403b3ac6} /* (5, 9, 16) {real, imag} */,
  {32'h3eaac192, 32'h4083f90d} /* (5, 9, 15) {real, imag} */,
  {32'hbf08fc20, 32'h40720c08} /* (5, 9, 14) {real, imag} */,
  {32'hc0340618, 32'h409e98ea} /* (5, 9, 13) {real, imag} */,
  {32'hbf836a70, 32'h40402102} /* (5, 9, 12) {real, imag} */,
  {32'hbf31bf9a, 32'h3f5ce314} /* (5, 9, 11) {real, imag} */,
  {32'hbe2d0710, 32'hc00b3088} /* (5, 9, 10) {real, imag} */,
  {32'hbe1c5d64, 32'hc01032df} /* (5, 9, 9) {real, imag} */,
  {32'h407a7cec, 32'hc00105ca} /* (5, 9, 8) {real, imag} */,
  {32'h40477198, 32'hbd470ee0} /* (5, 9, 7) {real, imag} */,
  {32'h3e14dddc, 32'hbfd4e5e6} /* (5, 9, 6) {real, imag} */,
  {32'h3e9eadaa, 32'hc01ca331} /* (5, 9, 5) {real, imag} */,
  {32'h3ef0c3dc, 32'hbfd51801} /* (5, 9, 4) {real, imag} */,
  {32'h3f9593b3, 32'hbfba09d1} /* (5, 9, 3) {real, imag} */,
  {32'h402960e6, 32'hc034e680} /* (5, 9, 2) {real, imag} */,
  {32'h40063670, 32'hc05967c0} /* (5, 9, 1) {real, imag} */,
  {32'h3e4d3d20, 32'hc02a7c15} /* (5, 9, 0) {real, imag} */,
  {32'h3fbe5ebb, 32'hbfe15aef} /* (5, 8, 31) {real, imag} */,
  {32'h40125754, 32'hbfed7b18} /* (5, 8, 30) {real, imag} */,
  {32'hc0384e8f, 32'hc0795c30} /* (5, 8, 29) {real, imag} */,
  {32'hbf0f9fdd, 32'hc079746d} /* (5, 8, 28) {real, imag} */,
  {32'h3e229b78, 32'hc0167e07} /* (5, 8, 27) {real, imag} */,
  {32'h3f08f944, 32'hbfded139} /* (5, 8, 26) {real, imag} */,
  {32'h3e58dc97, 32'hc03288f7} /* (5, 8, 25) {real, imag} */,
  {32'h40371e84, 32'hc0122ecb} /* (5, 8, 24) {real, imag} */,
  {32'h3fef3067, 32'h3e39aaf0} /* (5, 8, 23) {real, imag} */,
  {32'hbaee0c00, 32'hc028240a} /* (5, 8, 22) {real, imag} */,
  {32'hbf50fc2a, 32'h3e7dd6e0} /* (5, 8, 21) {real, imag} */,
  {32'hbf60e8b5, 32'h3f826c56} /* (5, 8, 20) {real, imag} */,
  {32'hc004a49e, 32'h3f990010} /* (5, 8, 19) {real, imag} */,
  {32'hc002da67, 32'h40a25daa} /* (5, 8, 18) {real, imag} */,
  {32'hc01f4fb8, 32'h405ee326} /* (5, 8, 17) {real, imag} */,
  {32'hc0667012, 32'h4066fa2a} /* (5, 8, 16) {real, imag} */,
  {32'hbfdd6a8a, 32'h4061c06e} /* (5, 8, 15) {real, imag} */,
  {32'h3eacf902, 32'h3f11fda2} /* (5, 8, 14) {real, imag} */,
  {32'hbf6b9dba, 32'h40837c86} /* (5, 8, 13) {real, imag} */,
  {32'hbff05e1d, 32'h4073b0bf} /* (5, 8, 12) {real, imag} */,
  {32'h3f66b7dc, 32'h40352d39} /* (5, 8, 11) {real, imag} */,
  {32'h3fc2595a, 32'hbf699778} /* (5, 8, 10) {real, imag} */,
  {32'h4020e12c, 32'hbfeda017} /* (5, 8, 9) {real, imag} */,
  {32'h409720b0, 32'hc0328cf0} /* (5, 8, 8) {real, imag} */,
  {32'h4024cd42, 32'hc0473ee2} /* (5, 8, 7) {real, imag} */,
  {32'hbe3c0fa4, 32'hc0b84690} /* (5, 8, 6) {real, imag} */,
  {32'h400171ac, 32'hc0a5a14a} /* (5, 8, 5) {real, imag} */,
  {32'h40005d37, 32'hc0126cc4} /* (5, 8, 4) {real, imag} */,
  {32'h3fd1f30d, 32'hbf4db8f4} /* (5, 8, 3) {real, imag} */,
  {32'h3fa4c52c, 32'hbfeb5dfc} /* (5, 8, 2) {real, imag} */,
  {32'h3e7bc294, 32'hc022bc0c} /* (5, 8, 1) {real, imag} */,
  {32'hbee21331, 32'hc02ee007} /* (5, 8, 0) {real, imag} */,
  {32'h3f71460a, 32'hbf2d94d8} /* (5, 7, 31) {real, imag} */,
  {32'h3fa9b1a4, 32'hc00e12b6} /* (5, 7, 30) {real, imag} */,
  {32'hc048988b, 32'hc00c80be} /* (5, 7, 29) {real, imag} */,
  {32'hbf8d46ce, 32'hbff1a5f8} /* (5, 7, 28) {real, imag} */,
  {32'h3fcd3620, 32'hbfd8dba7} /* (5, 7, 27) {real, imag} */,
  {32'h400b8532, 32'hbf7219d6} /* (5, 7, 26) {real, imag} */,
  {32'hbed910c8, 32'hc03b3b0c} /* (5, 7, 25) {real, imag} */,
  {32'h3f1a9f26, 32'hc067830d} /* (5, 7, 24) {real, imag} */,
  {32'h401a2e0c, 32'hc03400bc} /* (5, 7, 23) {real, imag} */,
  {32'h3fc51d8b, 32'hc045f23a} /* (5, 7, 22) {real, imag} */,
  {32'hc00c30dc, 32'hbf571c4d} /* (5, 7, 21) {real, imag} */,
  {32'hc0090901, 32'h40109917} /* (5, 7, 20) {real, imag} */,
  {32'hbcb7f000, 32'h406684d0} /* (5, 7, 19) {real, imag} */,
  {32'hbf062611, 32'h40966009} /* (5, 7, 18) {real, imag} */,
  {32'hc04fe8c1, 32'h40a7e684} /* (5, 7, 17) {real, imag} */,
  {32'hc03d4d73, 32'h40264d18} /* (5, 7, 16) {real, imag} */,
  {32'hbf8710f8, 32'h3f988b5c} /* (5, 7, 15) {real, imag} */,
  {32'hbf98656f, 32'hbeefb5d4} /* (5, 7, 14) {real, imag} */,
  {32'hbfe8b1e6, 32'h40207fd0} /* (5, 7, 13) {real, imag} */,
  {32'hbfc125b7, 32'h4013189b} /* (5, 7, 12) {real, imag} */,
  {32'hc0457f56, 32'h40889118} /* (5, 7, 11) {real, imag} */,
  {32'h3f6910fc, 32'hbf1d8fa4} /* (5, 7, 10) {real, imag} */,
  {32'h400c9a66, 32'hc04c4748} /* (5, 7, 9) {real, imag} */,
  {32'h3fce6f04, 32'hc091f98a} /* (5, 7, 8) {real, imag} */,
  {32'h3eba6e73, 32'hbfa94294} /* (5, 7, 7) {real, imag} */,
  {32'h3f7c0ee5, 32'hc043d01d} /* (5, 7, 6) {real, imag} */,
  {32'h3e982430, 32'hc05140ca} /* (5, 7, 5) {real, imag} */,
  {32'h3fe8c095, 32'hbfbe9a43} /* (5, 7, 4) {real, imag} */,
  {32'h401f7eff, 32'h3facacc9} /* (5, 7, 3) {real, imag} */,
  {32'h3ec43580, 32'h3fde82aa} /* (5, 7, 2) {real, imag} */,
  {32'hbf92bef4, 32'hbfd8e47c} /* (5, 7, 1) {real, imag} */,
  {32'hbd057ae0, 32'hc01e2092} /* (5, 7, 0) {real, imag} */,
  {32'hbe4da3d6, 32'h3cb2fbb0} /* (5, 6, 31) {real, imag} */,
  {32'h3f0f9c30, 32'hc006c30f} /* (5, 6, 30) {real, imag} */,
  {32'h3f8b3142, 32'hc07a41a2} /* (5, 6, 29) {real, imag} */,
  {32'h3fa4c70a, 32'hbfa20c29} /* (5, 6, 28) {real, imag} */,
  {32'h407f0e84, 32'hbe8a958c} /* (5, 6, 27) {real, imag} */,
  {32'h40398812, 32'hc00f0a67} /* (5, 6, 26) {real, imag} */,
  {32'h3fb64a27, 32'hc05217c0} /* (5, 6, 25) {real, imag} */,
  {32'hbf1cf722, 32'hc04afc71} /* (5, 6, 24) {real, imag} */,
  {32'h3e14e8dc, 32'hc0748d60} /* (5, 6, 23) {real, imag} */,
  {32'h3fd7adfc, 32'hc08dd33b} /* (5, 6, 22) {real, imag} */,
  {32'hbef58e78, 32'hc04af78c} /* (5, 6, 21) {real, imag} */,
  {32'hc004aef2, 32'hbef34cda} /* (5, 6, 20) {real, imag} */,
  {32'hbf93629e, 32'h404ac6e8} /* (5, 6, 19) {real, imag} */,
  {32'hbf1cf8b6, 32'h4050dc91} /* (5, 6, 18) {real, imag} */,
  {32'hc02867b1, 32'h401c8c4b} /* (5, 6, 17) {real, imag} */,
  {32'hbf959bdc, 32'h3d9376c0} /* (5, 6, 16) {real, imag} */,
  {32'h3e829736, 32'h3f49112f} /* (5, 6, 15) {real, imag} */,
  {32'hbea56f96, 32'h400a7da4} /* (5, 6, 14) {real, imag} */,
  {32'hc0094f1b, 32'h404b3b10} /* (5, 6, 13) {real, imag} */,
  {32'hbdb42508, 32'h3f9fc3bd} /* (5, 6, 12) {real, imag} */,
  {32'hc02723d8, 32'h3f99942d} /* (5, 6, 11) {real, imag} */,
  {32'hbdc371f8, 32'hbf120737} /* (5, 6, 10) {real, imag} */,
  {32'h400cedca, 32'hbfbe9bb7} /* (5, 6, 9) {real, imag} */,
  {32'h40461ec9, 32'hbfa5b1e1} /* (5, 6, 8) {real, imag} */,
  {32'h3fb8499b, 32'h3e02d7b8} /* (5, 6, 7) {real, imag} */,
  {32'h4025067e, 32'hbfcbdc64} /* (5, 6, 6) {real, imag} */,
  {32'hbf85d34e, 32'hc04ddd92} /* (5, 6, 5) {real, imag} */,
  {32'hbe91231e, 32'hc085a002} /* (5, 6, 4) {real, imag} */,
  {32'h3f2d27ee, 32'hbfd3f724} /* (5, 6, 3) {real, imag} */,
  {32'h401c033a, 32'hbfa433e4} /* (5, 6, 2) {real, imag} */,
  {32'h400a72dd, 32'hc04dba13} /* (5, 6, 1) {real, imag} */,
  {32'h3f8da5f8, 32'hc000f5ca} /* (5, 6, 0) {real, imag} */,
  {32'h3ed1455e, 32'h3cc34ea0} /* (5, 5, 31) {real, imag} */,
  {32'hbda8a308, 32'hbf93038a} /* (5, 5, 30) {real, imag} */,
  {32'h3fd636d9, 32'hc06bdaa4} /* (5, 5, 29) {real, imag} */,
  {32'h3fef4fb3, 32'hc07f27d4} /* (5, 5, 28) {real, imag} */,
  {32'h403c7e11, 32'hbf965e66} /* (5, 5, 27) {real, imag} */,
  {32'h401b1563, 32'hbc290ec0} /* (5, 5, 26) {real, imag} */,
  {32'h400274f8, 32'hc0573922} /* (5, 5, 25) {real, imag} */,
  {32'h3eb169b4, 32'hc0650529} /* (5, 5, 24) {real, imag} */,
  {32'hbeb9eb18, 32'hc0060b54} /* (5, 5, 23) {real, imag} */,
  {32'hbea45154, 32'hc08b28fc} /* (5, 5, 22) {real, imag} */,
  {32'h3f408ea0, 32'hc093a6d2} /* (5, 5, 21) {real, imag} */,
  {32'hbf1418be, 32'hc09d5e26} /* (5, 5, 20) {real, imag} */,
  {32'hbf9142ae, 32'hc0044c1e} /* (5, 5, 19) {real, imag} */,
  {32'hbf7adb04, 32'hbce434e0} /* (5, 5, 18) {real, imag} */,
  {32'hbe993f11, 32'hbf416d15} /* (5, 5, 17) {real, imag} */,
  {32'h3fc1f95c, 32'h3f4455b8} /* (5, 5, 16) {real, imag} */,
  {32'hbfa53e68, 32'h3fed65ba} /* (5, 5, 15) {real, imag} */,
  {32'hc089f20c, 32'h40762eed} /* (5, 5, 14) {real, imag} */,
  {32'hc044637a, 32'h4006c9d0} /* (5, 5, 13) {real, imag} */,
  {32'h3e2262a0, 32'h3f1b2fec} /* (5, 5, 12) {real, imag} */,
  {32'h3f4488f5, 32'hbf42766c} /* (5, 5, 11) {real, imag} */,
  {32'hbf8bfe4a, 32'h3fb8ec45} /* (5, 5, 10) {real, imag} */,
  {32'hbf758334, 32'h3f3be7be} /* (5, 5, 9) {real, imag} */,
  {32'hbff93f81, 32'h3f7765e6} /* (5, 5, 8) {real, imag} */,
  {32'hc00a282a, 32'h3f224ce5} /* (5, 5, 7) {real, imag} */,
  {32'hbfe9cac6, 32'hbee7bb7e} /* (5, 5, 6) {real, imag} */,
  {32'hc00c9a2e, 32'hc0588c3f} /* (5, 5, 5) {real, imag} */,
  {32'hbeef24ca, 32'hc00c9977} /* (5, 5, 4) {real, imag} */,
  {32'h3f3a3f3e, 32'hbf283d62} /* (5, 5, 3) {real, imag} */,
  {32'h3f7f6148, 32'hbfe36d9e} /* (5, 5, 2) {real, imag} */,
  {32'h3d47df10, 32'hc054d7a4} /* (5, 5, 1) {real, imag} */,
  {32'h3f2033ad, 32'hc01d060c} /* (5, 5, 0) {real, imag} */,
  {32'h3f18c680, 32'hbf4a1d45} /* (5, 4, 31) {real, imag} */,
  {32'h4022e5f8, 32'hc0219400} /* (5, 4, 30) {real, imag} */,
  {32'h3fc52fcb, 32'hc066772f} /* (5, 4, 29) {real, imag} */,
  {32'h3f0a3f3e, 32'hc093ba69} /* (5, 4, 28) {real, imag} */,
  {32'h3f98b6e2, 32'hbfaa5788} /* (5, 4, 27) {real, imag} */,
  {32'h40298ee1, 32'h40434833} /* (5, 4, 26) {real, imag} */,
  {32'h4036a730, 32'h3ff96190} /* (5, 4, 25) {real, imag} */,
  {32'h3f43d3e7, 32'hc01c5be8} /* (5, 4, 24) {real, imag} */,
  {32'h3fac1bf6, 32'hc06865f1} /* (5, 4, 23) {real, imag} */,
  {32'h3fc202c0, 32'hc0a11ebb} /* (5, 4, 22) {real, imag} */,
  {32'h400bb3c2, 32'hc0affbfc} /* (5, 4, 21) {real, imag} */,
  {32'h3fdbd92d, 32'hc02d8bac} /* (5, 4, 20) {real, imag} */,
  {32'hbebd045d, 32'hbfdafaa4} /* (5, 4, 19) {real, imag} */,
  {32'h3ed4b624, 32'hc008c4f2} /* (5, 4, 18) {real, imag} */,
  {32'h3f132a63, 32'hc0107b40} /* (5, 4, 17) {real, imag} */,
  {32'h400b4958, 32'hbf01fe40} /* (5, 4, 16) {real, imag} */,
  {32'hbf4d1a18, 32'h3ec99c56} /* (5, 4, 15) {real, imag} */,
  {32'hc097baa9, 32'h3f604f30} /* (5, 4, 14) {real, imag} */,
  {32'hc055cd6c, 32'h3fc91f68} /* (5, 4, 13) {real, imag} */,
  {32'hbf9ce882, 32'h3fb77687} /* (5, 4, 12) {real, imag} */,
  {32'h3efdd552, 32'hbd21bcf0} /* (5, 4, 11) {real, imag} */,
  {32'hc01addae, 32'hbf0b14c8} /* (5, 4, 10) {real, imag} */,
  {32'hc0612674, 32'h3fb52539} /* (5, 4, 9) {real, imag} */,
  {32'hc04ac067, 32'h3fca405d} /* (5, 4, 8) {real, imag} */,
  {32'hbff152a2, 32'h3ed18e0e} /* (5, 4, 7) {real, imag} */,
  {32'hc0700ab3, 32'h3fa43262} /* (5, 4, 6) {real, imag} */,
  {32'hc0193114, 32'hc02a7e14} /* (5, 4, 5) {real, imag} */,
  {32'h3f679882, 32'hc098e85e} /* (5, 4, 4) {real, imag} */,
  {32'h3ff75ee3, 32'hc04a812b} /* (5, 4, 3) {real, imag} */,
  {32'h3f9d9032, 32'hbfb14c3c} /* (5, 4, 2) {real, imag} */,
  {32'h3fc9a178, 32'hbed27ff1} /* (5, 4, 1) {real, imag} */,
  {32'h3fa46c53, 32'hbe7a8e7e} /* (5, 4, 0) {real, imag} */,
  {32'h3ff9e249, 32'hbfa8f971} /* (5, 3, 31) {real, imag} */,
  {32'h40a7d4dc, 32'hbfc1657f} /* (5, 3, 30) {real, imag} */,
  {32'h4032a0cd, 32'hbf915aa4} /* (5, 3, 29) {real, imag} */,
  {32'h3fd33b48, 32'hc06c610e} /* (5, 3, 28) {real, imag} */,
  {32'h4004a288, 32'hc040b55f} /* (5, 3, 27) {real, imag} */,
  {32'h3ff872cb, 32'hbe6a4d90} /* (5, 3, 26) {real, imag} */,
  {32'h4042fc02, 32'h3fd76853} /* (5, 3, 25) {real, imag} */,
  {32'h3fd53ea8, 32'hbf8ff66b} /* (5, 3, 24) {real, imag} */,
  {32'h3f909b94, 32'hbfd8c1ff} /* (5, 3, 23) {real, imag} */,
  {32'h3fe946a3, 32'hc029a855} /* (5, 3, 22) {real, imag} */,
  {32'h3fac9610, 32'hc02c6056} /* (5, 3, 21) {real, imag} */,
  {32'hbf79c520, 32'hbfc13282} /* (5, 3, 20) {real, imag} */,
  {32'hbfba1c1b, 32'hc0201bc2} /* (5, 3, 19) {real, imag} */,
  {32'h4049d2de, 32'hc0a49ca2} /* (5, 3, 18) {real, imag} */,
  {32'h3fa26937, 32'hbfe7fadf} /* (5, 3, 17) {real, imag} */,
  {32'h3fb7a111, 32'hc0213197} /* (5, 3, 16) {real, imag} */,
  {32'hbf59bc4c, 32'h3eaabf7a} /* (5, 3, 15) {real, imag} */,
  {32'hc09353c7, 32'h3ed6673a} /* (5, 3, 14) {real, imag} */,
  {32'hc03ac4fd, 32'h4089c132} /* (5, 3, 13) {real, imag} */,
  {32'hbf83d2e0, 32'h405d44c0} /* (5, 3, 12) {real, imag} */,
  {32'hbfb6ccd8, 32'h3f22a140} /* (5, 3, 11) {real, imag} */,
  {32'hc03c3c2c, 32'hbf0c552d} /* (5, 3, 10) {real, imag} */,
  {32'hbff6a01b, 32'h401d23a1} /* (5, 3, 9) {real, imag} */,
  {32'hbec10c9e, 32'h3fa657e3} /* (5, 3, 8) {real, imag} */,
  {32'h3f9c2c41, 32'hbe3c2000} /* (5, 3, 7) {real, imag} */,
  {32'hc01a8732, 32'h3e41fabc} /* (5, 3, 6) {real, imag} */,
  {32'h3d88ec90, 32'hc01db864} /* (5, 3, 5) {real, imag} */,
  {32'h400d272b, 32'hc099d501} /* (5, 3, 4) {real, imag} */,
  {32'h4023502a, 32'hc097c59b} /* (5, 3, 3) {real, imag} */,
  {32'h4013ea19, 32'hc00853ca} /* (5, 3, 2) {real, imag} */,
  {32'h3f22139f, 32'hbf89e719} /* (5, 3, 1) {real, imag} */,
  {32'h3f3dbcff, 32'hbfd3b6b4} /* (5, 3, 0) {real, imag} */,
  {32'h3f5885b3, 32'hbf142448} /* (5, 2, 31) {real, imag} */,
  {32'h3fe38d45, 32'hbfa1ebce} /* (5, 2, 30) {real, imag} */,
  {32'h4053636e, 32'h3e623976} /* (5, 2, 29) {real, imag} */,
  {32'h3fe3ef70, 32'hbf4ed799} /* (5, 2, 28) {real, imag} */,
  {32'h40076cd9, 32'hc03ecb4e} /* (5, 2, 27) {real, imag} */,
  {32'h4088fd81, 32'hc0499588} /* (5, 2, 26) {real, imag} */,
  {32'h408420d2, 32'hbf1c8f70} /* (5, 2, 25) {real, imag} */,
  {32'h3fff1ae9, 32'hc0024e78} /* (5, 2, 24) {real, imag} */,
  {32'hbf53a4ec, 32'hc014a4ba} /* (5, 2, 23) {real, imag} */,
  {32'h3f8953ae, 32'hc0236e9c} /* (5, 2, 22) {real, imag} */,
  {32'h4086014b, 32'hc019d7c5} /* (5, 2, 21) {real, imag} */,
  {32'h402da5ea, 32'hbff05191} /* (5, 2, 20) {real, imag} */,
  {32'h3f96894a, 32'hc0ab63be} /* (5, 2, 19) {real, imag} */,
  {32'h4021a4f8, 32'hc0cc2772} /* (5, 2, 18) {real, imag} */,
  {32'h3fcf4cca, 32'hc0c07053} /* (5, 2, 17) {real, imag} */,
  {32'h4015f1e0, 32'hc0a55ad5} /* (5, 2, 16) {real, imag} */,
  {32'h3ef69545, 32'h3eee41d8} /* (5, 2, 15) {real, imag} */,
  {32'hc02e8321, 32'hbde6a60c} /* (5, 2, 14) {real, imag} */,
  {32'hbfc16c1e, 32'h4010beaa} /* (5, 2, 13) {real, imag} */,
  {32'hbf9f4cb5, 32'h405b875d} /* (5, 2, 12) {real, imag} */,
  {32'hbfa0da0e, 32'h401116ec} /* (5, 2, 11) {real, imag} */,
  {32'h3ed8fff4, 32'h40139bf7} /* (5, 2, 10) {real, imag} */,
  {32'h3f6a59db, 32'h4095b350} /* (5, 2, 9) {real, imag} */,
  {32'hbf998b22, 32'h402bb511} /* (5, 2, 8) {real, imag} */,
  {32'h3e51fc54, 32'h3f884678} /* (5, 2, 7) {real, imag} */,
  {32'hbe32c23c, 32'h3f1557c2} /* (5, 2, 6) {real, imag} */,
  {32'h3f7d31bb, 32'hc028ff6e} /* (5, 2, 5) {real, imag} */,
  {32'h3fba47a8, 32'hc0235d3a} /* (5, 2, 4) {real, imag} */,
  {32'h3fc85d95, 32'hc04db895} /* (5, 2, 3) {real, imag} */,
  {32'h4088bfb6, 32'hc051cb9a} /* (5, 2, 2) {real, imag} */,
  {32'h4017c5a1, 32'hbfbb0b08} /* (5, 2, 1) {real, imag} */,
  {32'h3f8d95fc, 32'hbfb1d088} /* (5, 2, 0) {real, imag} */,
  {32'hbe0b1848, 32'hbefb366f} /* (5, 1, 31) {real, imag} */,
  {32'h3ef76a22, 32'hbfd663e2} /* (5, 1, 30) {real, imag} */,
  {32'h3f7953a1, 32'hc0002ba2} /* (5, 1, 29) {real, imag} */,
  {32'hbf063a34, 32'hbf55dc5c} /* (5, 1, 28) {real, imag} */,
  {32'h3fcf9f20, 32'hc01ca0f3} /* (5, 1, 27) {real, imag} */,
  {32'h405317b4, 32'hc013bcfc} /* (5, 1, 26) {real, imag} */,
  {32'h40403348, 32'hc029b606} /* (5, 1, 25) {real, imag} */,
  {32'h3f9b0e19, 32'hbf83d3b6} /* (5, 1, 24) {real, imag} */,
  {32'hbea1b6ae, 32'hbfa3687c} /* (5, 1, 23) {real, imag} */,
  {32'h3e67ad98, 32'hc05cd8cf} /* (5, 1, 22) {real, imag} */,
  {32'h3fe201cd, 32'hc06e0f86} /* (5, 1, 21) {real, imag} */,
  {32'h4076d79d, 32'hc00313ea} /* (5, 1, 20) {real, imag} */,
  {32'h3f761ff8, 32'hc0b373c7} /* (5, 1, 19) {real, imag} */,
  {32'h3d416ce0, 32'hc0d4023c} /* (5, 1, 18) {real, imag} */,
  {32'hbecfa014, 32'hc0f4e042} /* (5, 1, 17) {real, imag} */,
  {32'h3fcb36ef, 32'hc0a4a253} /* (5, 1, 16) {real, imag} */,
  {32'h3f76139d, 32'hbeb044ec} /* (5, 1, 15) {real, imag} */,
  {32'hbf942c57, 32'h3fcd815c} /* (5, 1, 14) {real, imag} */,
  {32'hbf944889, 32'h3fbf6c09} /* (5, 1, 13) {real, imag} */,
  {32'hbf129211, 32'h3ffe6bbd} /* (5, 1, 12) {real, imag} */,
  {32'h3f992399, 32'h404999e7} /* (5, 1, 11) {real, imag} */,
  {32'hbee82508, 32'h4067dcb8} /* (5, 1, 10) {real, imag} */,
  {32'hbe883eb8, 32'h40af76db} /* (5, 1, 9) {real, imag} */,
  {32'hc00b9933, 32'h40a4b02b} /* (5, 1, 8) {real, imag} */,
  {32'hc008e69a, 32'h401383ff} /* (5, 1, 7) {real, imag} */,
  {32'hc0165d50, 32'hbf18734e} /* (5, 1, 6) {real, imag} */,
  {32'h3f8b2fd9, 32'hbf81a75c} /* (5, 1, 5) {real, imag} */,
  {32'h3f886ffd, 32'h3ee514b5} /* (5, 1, 4) {real, imag} */,
  {32'hbf133b1b, 32'hbff24b90} /* (5, 1, 3) {real, imag} */,
  {32'h3eafc7ea, 32'hc05af4e4} /* (5, 1, 2) {real, imag} */,
  {32'h3ff2cbe3, 32'hbfba1748} /* (5, 1, 1) {real, imag} */,
  {32'h3fca0c38, 32'hbe8825e8} /* (5, 1, 0) {real, imag} */,
  {32'h3c77c3f0, 32'hbdd56508} /* (5, 0, 31) {real, imag} */,
  {32'h3f498e21, 32'hbf0a4718} /* (5, 0, 30) {real, imag} */,
  {32'h3effb5af, 32'hc0011877} /* (5, 0, 29) {real, imag} */,
  {32'hbf223992, 32'hbe8ad38e} /* (5, 0, 28) {real, imag} */,
  {32'h3ff15a78, 32'hbef80e34} /* (5, 0, 27) {real, imag} */,
  {32'h4060b48a, 32'hbf9d709a} /* (5, 0, 26) {real, imag} */,
  {32'h3ffcf6cd, 32'hbf91b86a} /* (5, 0, 25) {real, imag} */,
  {32'h3f9668a8, 32'hbefc3847} /* (5, 0, 24) {real, imag} */,
  {32'h3f96d8f6, 32'h3f0b4476} /* (5, 0, 23) {real, imag} */,
  {32'h3f31989a, 32'hbf489870} /* (5, 0, 22) {real, imag} */,
  {32'h3f107932, 32'hbfc10338} /* (5, 0, 21) {real, imag} */,
  {32'h407fd350, 32'hbf8dea08} /* (5, 0, 20) {real, imag} */,
  {32'h40172c40, 32'hc010b356} /* (5, 0, 19) {real, imag} */,
  {32'h3fcf79c4, 32'hc0382734} /* (5, 0, 18) {real, imag} */,
  {32'h3ef7ff18, 32'hbfcd7986} /* (5, 0, 17) {real, imag} */,
  {32'hbf54d43a, 32'hbf6cc9e1} /* (5, 0, 16) {real, imag} */,
  {32'hbf1d52a0, 32'hbe00e47b} /* (5, 0, 15) {real, imag} */,
  {32'hbfbfa2d6, 32'h3fad490e} /* (5, 0, 14) {real, imag} */,
  {32'hbe791d0c, 32'h3fb93300} /* (5, 0, 13) {real, imag} */,
  {32'hbc2864e0, 32'h400c0678} /* (5, 0, 12) {real, imag} */,
  {32'h3e485812, 32'h3ffb04aa} /* (5, 0, 11) {real, imag} */,
  {32'hbfabd68d, 32'h3f97babd} /* (5, 0, 10) {real, imag} */,
  {32'hbf39993b, 32'h3fc89ba0} /* (5, 0, 9) {real, imag} */,
  {32'hbec6cb85, 32'h4046b0ca} /* (5, 0, 8) {real, imag} */,
  {32'hbf658b20, 32'h3fc939a3} /* (5, 0, 7) {real, imag} */,
  {32'hbff1a2b8, 32'hbeda0001} /* (5, 0, 6) {real, imag} */,
  {32'hbd58bcc0, 32'h3f3dd043} /* (5, 0, 5) {real, imag} */,
  {32'h3ed89e86, 32'h3ef07906} /* (5, 0, 4) {real, imag} */,
  {32'h3e2538a8, 32'hbfc6a460} /* (5, 0, 3) {real, imag} */,
  {32'hbfebcc72, 32'hbfce4cb0} /* (5, 0, 2) {real, imag} */,
  {32'hbf239bac, 32'h3cf018c0} /* (5, 0, 1) {real, imag} */,
  {32'h3fac9f5c, 32'h3f946464} /* (5, 0, 0) {real, imag} */,
  {32'hbb2a1380, 32'h3fe55793} /* (4, 31, 31) {real, imag} */,
  {32'hbf90e643, 32'h408b3cbe} /* (4, 31, 30) {real, imag} */,
  {32'hbff18948, 32'h409a93bb} /* (4, 31, 29) {real, imag} */,
  {32'hc0111137, 32'h40940d86} /* (4, 31, 28) {real, imag} */,
  {32'hbf8b6595, 32'h404f7456} /* (4, 31, 27) {real, imag} */,
  {32'hbee810ca, 32'h40492ab4} /* (4, 31, 26) {real, imag} */,
  {32'hbe184ac0, 32'h4070082b} /* (4, 31, 25) {real, imag} */,
  {32'hbeedb80c, 32'h401c1d48} /* (4, 31, 24) {real, imag} */,
  {32'hbfa55d48, 32'h401de1e0} /* (4, 31, 23) {real, imag} */,
  {32'hbfe326f3, 32'h3fdd8fb0} /* (4, 31, 22) {real, imag} */,
  {32'hbf24f4e7, 32'h4008b007} /* (4, 31, 21) {real, imag} */,
  {32'h3f460b86, 32'hbe333028} /* (4, 31, 20) {real, imag} */,
  {32'h3dcc10e6, 32'hc0138e36} /* (4, 31, 19) {real, imag} */,
  {32'hbc029b18, 32'hc0514078} /* (4, 31, 18) {real, imag} */,
  {32'hbce60810, 32'hc0674750} /* (4, 31, 17) {real, imag} */,
  {32'hbf46230e, 32'hbf51c62e} /* (4, 31, 16) {real, imag} */,
  {32'hbed6b442, 32'hbfef3ef9} /* (4, 31, 15) {real, imag} */,
  {32'h3f6feee3, 32'hc0703adc} /* (4, 31, 14) {real, imag} */,
  {32'h3e56eaca, 32'hbfd0d051} /* (4, 31, 13) {real, imag} */,
  {32'h3f1245c8, 32'hbfee9fb4} /* (4, 31, 12) {real, imag} */,
  {32'h3fc36aca, 32'hc0425026} /* (4, 31, 11) {real, imag} */,
  {32'h3dd57516, 32'h3e4ae007} /* (4, 31, 10) {real, imag} */,
  {32'hbfef6c3a, 32'h40274b40} /* (4, 31, 9) {real, imag} */,
  {32'hbf03cca6, 32'h3ff60e7e} /* (4, 31, 8) {real, imag} */,
  {32'h3f4574ff, 32'h40109768} /* (4, 31, 7) {real, imag} */,
  {32'h3ea04386, 32'h40126892} /* (4, 31, 6) {real, imag} */,
  {32'hbfedc90c, 32'h404fab11} /* (4, 31, 5) {real, imag} */,
  {32'hc0308aea, 32'h3fedadf2} /* (4, 31, 4) {real, imag} */,
  {32'hbf8a19d3, 32'h403aaa7f} /* (4, 31, 3) {real, imag} */,
  {32'hbfbb08b9, 32'h4063a80d} /* (4, 31, 2) {real, imag} */,
  {32'hbeb3282a, 32'h4083d19b} /* (4, 31, 1) {real, imag} */,
  {32'h3db72ce0, 32'h3f86f732} /* (4, 31, 0) {real, imag} */,
  {32'hbdc034c8, 32'h4013bd4e} /* (4, 30, 31) {real, imag} */,
  {32'hbf07a3f6, 32'h40b6c985} /* (4, 30, 30) {real, imag} */,
  {32'hc0156a5f, 32'h40d50de8} /* (4, 30, 29) {real, imag} */,
  {32'hc025f80f, 32'h40b662d6} /* (4, 30, 28) {real, imag} */,
  {32'hbf747d9c, 32'h40a59a7a} /* (4, 30, 27) {real, imag} */,
  {32'hbe4f82f4, 32'h40dd9762} /* (4, 30, 26) {real, imag} */,
  {32'hc00b6af0, 32'h40baa496} /* (4, 30, 25) {real, imag} */,
  {32'hc010b3b6, 32'h4096e4a4} /* (4, 30, 24) {real, imag} */,
  {32'hc019ad80, 32'h40983df3} /* (4, 30, 23) {real, imag} */,
  {32'hbf88fb76, 32'h40aaba8b} /* (4, 30, 22) {real, imag} */,
  {32'h3e254958, 32'h405e82f6} /* (4, 30, 21) {real, imag} */,
  {32'h4004878d, 32'hc094def8} /* (4, 30, 20) {real, imag} */,
  {32'h3e808c24, 32'hc0bf083a} /* (4, 30, 19) {real, imag} */,
  {32'h3e9d3cb0, 32'hc0d878d1} /* (4, 30, 18) {real, imag} */,
  {32'h3faa11d6, 32'hc0eb3d2c} /* (4, 30, 17) {real, imag} */,
  {32'h3ea3113b, 32'hc0a6342b} /* (4, 30, 16) {real, imag} */,
  {32'h3f19b7d0, 32'hc0d5dc40} /* (4, 30, 15) {real, imag} */,
  {32'h4010b6e4, 32'hc0f5aba5} /* (4, 30, 14) {real, imag} */,
  {32'h3e50516b, 32'hc0a43b5d} /* (4, 30, 13) {real, imag} */,
  {32'h3f0cdaa8, 32'hc07b3916} /* (4, 30, 12) {real, imag} */,
  {32'h3fd0ca79, 32'hc09960eb} /* (4, 30, 11) {real, imag} */,
  {32'hbf92456a, 32'hbf78f616} /* (4, 30, 10) {real, imag} */,
  {32'hc0a974a2, 32'h40992024} /* (4, 30, 9) {real, imag} */,
  {32'hc068fea2, 32'h4095a244} /* (4, 30, 8) {real, imag} */,
  {32'hc0048eaa, 32'h4096d4fe} /* (4, 30, 7) {real, imag} */,
  {32'hbfbbe76c, 32'h40b281d4} /* (4, 30, 6) {real, imag} */,
  {32'hbf8e0f6a, 32'h405749f6} /* (4, 30, 5) {real, imag} */,
  {32'hc0889d88, 32'h4085f3b7} /* (4, 30, 4) {real, imag} */,
  {32'hc0ae5a0d, 32'h40aed984} /* (4, 30, 3) {real, imag} */,
  {32'hc040e772, 32'h40c292fa} /* (4, 30, 2) {real, imag} */,
  {32'h40043288, 32'h40cc3f6e} /* (4, 30, 1) {real, imag} */,
  {32'h3f005c94, 32'h40509a90} /* (4, 30, 0) {real, imag} */,
  {32'hbf47c2ec, 32'h3feade69} /* (4, 29, 31) {real, imag} */,
  {32'hc02496a6, 32'h4086ec38} /* (4, 29, 30) {real, imag} */,
  {32'hc087ba82, 32'h40ab6893} /* (4, 29, 29) {real, imag} */,
  {32'hc046d46c, 32'h405a19ae} /* (4, 29, 28) {real, imag} */,
  {32'hbfdf22df, 32'h40634daf} /* (4, 29, 27) {real, imag} */,
  {32'hbfce3c82, 32'h40b0fad6} /* (4, 29, 26) {real, imag} */,
  {32'hc02e0596, 32'h408d2941} /* (4, 29, 25) {real, imag} */,
  {32'hc03cba01, 32'h40c41a2c} /* (4, 29, 24) {real, imag} */,
  {32'hc06161b6, 32'h40a8e8e4} /* (4, 29, 23) {real, imag} */,
  {32'hbf09144d, 32'h40c2fb5e} /* (4, 29, 22) {real, imag} */,
  {32'hbfbf2ab7, 32'h40011eac} /* (4, 29, 21) {real, imag} */,
  {32'h3f1c87fe, 32'hc1085f15} /* (4, 29, 20) {real, imag} */,
  {32'h3fd82dce, 32'hc0a3368a} /* (4, 29, 19) {real, imag} */,
  {32'h401c927a, 32'hc089cba2} /* (4, 29, 18) {real, imag} */,
  {32'h40396f4a, 32'hc0dc199a} /* (4, 29, 17) {real, imag} */,
  {32'h3fdeb468, 32'hc0cfdbfe} /* (4, 29, 16) {real, imag} */,
  {32'h3fc702f2, 32'hc08fdfaa} /* (4, 29, 15) {real, imag} */,
  {32'h408e720c, 32'hc0ce3d04} /* (4, 29, 14) {real, imag} */,
  {32'h40360b6c, 32'hc0aedb02} /* (4, 29, 13) {real, imag} */,
  {32'h3f9bbc5d, 32'hc03e5fe8} /* (4, 29, 12) {real, imag} */,
  {32'hbbdd3200, 32'hc04eed4a} /* (4, 29, 11) {real, imag} */,
  {32'hbf6a4468, 32'h3f80b78a} /* (4, 29, 10) {real, imag} */,
  {32'hc0601efb, 32'h40903ba1} /* (4, 29, 9) {real, imag} */,
  {32'hc09175f2, 32'h40aeb010} /* (4, 29, 8) {real, imag} */,
  {32'hc08eb3ea, 32'h40a18ea4} /* (4, 29, 7) {real, imag} */,
  {32'hc05a39ec, 32'h4084bd91} /* (4, 29, 6) {real, imag} */,
  {32'hbfbb9a0d, 32'h40a210f5} /* (4, 29, 5) {real, imag} */,
  {32'hbfb0814f, 32'h40ba5900} /* (4, 29, 4) {real, imag} */,
  {32'hc09cb02c, 32'h40c1b964} /* (4, 29, 3) {real, imag} */,
  {32'hc093d571, 32'h408d877d} /* (4, 29, 2) {real, imag} */,
  {32'hbf164c1d, 32'h408f6657} /* (4, 29, 1) {real, imag} */,
  {32'hbd86e7c4, 32'h4064c9fa} /* (4, 29, 0) {real, imag} */,
  {32'hc016c7e0, 32'h3f25b102} /* (4, 28, 31) {real, imag} */,
  {32'hc0ab7c2b, 32'h4085a30a} /* (4, 28, 30) {real, imag} */,
  {32'hc0a61fc4, 32'h40e85491} /* (4, 28, 29) {real, imag} */,
  {32'hbfa71630, 32'h40ca9aea} /* (4, 28, 28) {real, imag} */,
  {32'hc02e86b9, 32'h4065476b} /* (4, 28, 27) {real, imag} */,
  {32'hc078dbec, 32'h40b20909} /* (4, 28, 26) {real, imag} */,
  {32'hbfc18f70, 32'h40a0f07a} /* (4, 28, 25) {real, imag} */,
  {32'hbf4a4dd7, 32'h40988319} /* (4, 28, 24) {real, imag} */,
  {32'hc007a982, 32'h406897b5} /* (4, 28, 23) {real, imag} */,
  {32'hbf610d54, 32'h40987f84} /* (4, 28, 22) {real, imag} */,
  {32'hc08a8d4b, 32'h406010b9} /* (4, 28, 21) {real, imag} */,
  {32'hbea3f1e3, 32'hc09dde1f} /* (4, 28, 20) {real, imag} */,
  {32'h408a37d7, 32'hc05b1728} /* (4, 28, 19) {real, imag} */,
  {32'h40e01572, 32'hc0848f96} /* (4, 28, 18) {real, imag} */,
  {32'h40a69e65, 32'hc0ba0cd5} /* (4, 28, 17) {real, imag} */,
  {32'h403efab7, 32'hc0447d1b} /* (4, 28, 16) {real, imag} */,
  {32'h40274cd4, 32'h3f8e8b4d} /* (4, 28, 15) {real, imag} */,
  {32'h40488b07, 32'hc073afa8} /* (4, 28, 14) {real, imag} */,
  {32'h4050fc47, 32'hc05bd2ae} /* (4, 28, 13) {real, imag} */,
  {32'h40291dc4, 32'hc0031ab8} /* (4, 28, 12) {real, imag} */,
  {32'hbdc27239, 32'hc05088d4} /* (4, 28, 11) {real, imag} */,
  {32'hc0426f54, 32'h405bfde2} /* (4, 28, 10) {real, imag} */,
  {32'hc0743e51, 32'h4095fc97} /* (4, 28, 9) {real, imag} */,
  {32'hbfee131e, 32'h40967b94} /* (4, 28, 8) {real, imag} */,
  {32'hc054cec0, 32'h40a61689} /* (4, 28, 7) {real, imag} */,
  {32'hc07ca72c, 32'h40192f76} /* (4, 28, 6) {real, imag} */,
  {32'hc053d66a, 32'h40655256} /* (4, 28, 5) {real, imag} */,
  {32'hc01aa901, 32'h40782550} /* (4, 28, 4) {real, imag} */,
  {32'hc056480b, 32'h408f1f36} /* (4, 28, 3) {real, imag} */,
  {32'hc0a09c37, 32'h4026859a} /* (4, 28, 2) {real, imag} */,
  {32'hc055a9f9, 32'h3fcd5630} /* (4, 28, 1) {real, imag} */,
  {32'hbf9f8c05, 32'h3f9fa1f4} /* (4, 28, 0) {real, imag} */,
  {32'hbf169ff6, 32'h4008b328} /* (4, 27, 31) {real, imag} */,
  {32'hc09cbe4e, 32'h40a9d4a4} /* (4, 27, 30) {real, imag} */,
  {32'hc0caa516, 32'h409921f5} /* (4, 27, 29) {real, imag} */,
  {32'hc025eef4, 32'h401de5d0} /* (4, 27, 28) {real, imag} */,
  {32'hc0628fe0, 32'hbd132b08} /* (4, 27, 27) {real, imag} */,
  {32'hc06a927a, 32'h408ce195} /* (4, 27, 26) {real, imag} */,
  {32'hbea2df6d, 32'h40c4c861} /* (4, 27, 25) {real, imag} */,
  {32'h3feab81e, 32'h406061a2} /* (4, 27, 24) {real, imag} */,
  {32'h3e0caf6f, 32'h4032e1c7} /* (4, 27, 23) {real, imag} */,
  {32'hc028eed8, 32'h40aaccda} /* (4, 27, 22) {real, imag} */,
  {32'hc02c8fcc, 32'h40d207ff} /* (4, 27, 21) {real, imag} */,
  {32'hbdcd27b0, 32'hc00c4e4e} /* (4, 27, 20) {real, imag} */,
  {32'h40803974, 32'hc086525b} /* (4, 27, 19) {real, imag} */,
  {32'h40e95260, 32'hc07b7c08} /* (4, 27, 18) {real, imag} */,
  {32'h40574d74, 32'hc047c8e4} /* (4, 27, 17) {real, imag} */,
  {32'h400fbcc6, 32'hc03fb99c} /* (4, 27, 16) {real, imag} */,
  {32'h3f0c9959, 32'hbfbd191e} /* (4, 27, 15) {real, imag} */,
  {32'h3eb15fb4, 32'hc0946206} /* (4, 27, 14) {real, imag} */,
  {32'hbe92c52a, 32'hc0aa950a} /* (4, 27, 13) {real, imag} */,
  {32'h3fa519f4, 32'hc04ce1a0} /* (4, 27, 12) {real, imag} */,
  {32'h3feae9ca, 32'hc073678e} /* (4, 27, 11) {real, imag} */,
  {32'hbeb0378c, 32'h4088142a} /* (4, 27, 10) {real, imag} */,
  {32'hc081bfd1, 32'h40c23e38} /* (4, 27, 9) {real, imag} */,
  {32'hc03fe1e6, 32'h409307cc} /* (4, 27, 8) {real, imag} */,
  {32'hc040192a, 32'h409e8c84} /* (4, 27, 7) {real, imag} */,
  {32'hc03d3ca2, 32'h4099bb48} /* (4, 27, 6) {real, imag} */,
  {32'hc007f916, 32'h40913fd5} /* (4, 27, 5) {real, imag} */,
  {32'hc030c9cf, 32'h40356a6a} /* (4, 27, 4) {real, imag} */,
  {32'hc0800b18, 32'h406a34f1} /* (4, 27, 3) {real, imag} */,
  {32'hc03ce924, 32'h405c81e2} /* (4, 27, 2) {real, imag} */,
  {32'hbfac887f, 32'h40008524} /* (4, 27, 1) {real, imag} */,
  {32'hbe566e50, 32'hbf43e9b6} /* (4, 27, 0) {real, imag} */,
  {32'hbfd5c54c, 32'h3febb8d8} /* (4, 26, 31) {real, imag} */,
  {32'hc097cb72, 32'h40756506} /* (4, 26, 30) {real, imag} */,
  {32'hc06bd624, 32'h40902e08} /* (4, 26, 29) {real, imag} */,
  {32'hbeb9e438, 32'h40950e7a} /* (4, 26, 28) {real, imag} */,
  {32'hc04c131f, 32'h405af4a0} /* (4, 26, 27) {real, imag} */,
  {32'hc086f3be, 32'h40928714} /* (4, 26, 26) {real, imag} */,
  {32'hbfeaa5c6, 32'h40908790} /* (4, 26, 25) {real, imag} */,
  {32'h3fd56e5f, 32'h3f62958b} /* (4, 26, 24) {real, imag} */,
  {32'h3f46e86a, 32'h4012815d} /* (4, 26, 23) {real, imag} */,
  {32'hbfc93e91, 32'h406cf66e} /* (4, 26, 22) {real, imag} */,
  {32'hbdf04118, 32'h406c533c} /* (4, 26, 21) {real, imag} */,
  {32'h3f7fad97, 32'hc04fb3a2} /* (4, 26, 20) {real, imag} */,
  {32'h3fb08e5a, 32'hc05ab486} /* (4, 26, 19) {real, imag} */,
  {32'h4033323a, 32'hc0140fb6} /* (4, 26, 18) {real, imag} */,
  {32'h3fce4922, 32'hbfd2c397} /* (4, 26, 17) {real, imag} */,
  {32'h40437fd0, 32'hc095fbca} /* (4, 26, 16) {real, imag} */,
  {32'hbd59a328, 32'hc06e9d5a} /* (4, 26, 15) {real, imag} */,
  {32'hbfb23083, 32'hc0a7d15c} /* (4, 26, 14) {real, imag} */,
  {32'hbfdc182e, 32'hc0babf64} /* (4, 26, 13) {real, imag} */,
  {32'hbe23c0f3, 32'hc0970b3c} /* (4, 26, 12) {real, imag} */,
  {32'h3fe8af80, 32'hc0696bc0} /* (4, 26, 11) {real, imag} */,
  {32'h3f713c70, 32'h3fbcd5bd} /* (4, 26, 10) {real, imag} */,
  {32'hc0807cf0, 32'h404a415a} /* (4, 26, 9) {real, imag} */,
  {32'hc074fb93, 32'h40bad20f} /* (4, 26, 8) {real, imag} */,
  {32'hbf98a13c, 32'h40bf9a9e} /* (4, 26, 7) {real, imag} */,
  {32'hbfdd403a, 32'h40bab092} /* (4, 26, 6) {real, imag} */,
  {32'hbfbea09f, 32'h40b68e2c} /* (4, 26, 5) {real, imag} */,
  {32'hbfbd60a2, 32'h4041086a} /* (4, 26, 4) {real, imag} */,
  {32'hc0391268, 32'h408961f5} /* (4, 26, 3) {real, imag} */,
  {32'hbff74f58, 32'h409e7692} /* (4, 26, 2) {real, imag} */,
  {32'hbfe1cc50, 32'h40a33945} /* (4, 26, 1) {real, imag} */,
  {32'hbf817817, 32'h3fe02d97} /* (4, 26, 0) {real, imag} */,
  {32'hbfeea039, 32'h40715f54} /* (4, 25, 31) {real, imag} */,
  {32'hc0932852, 32'h40c9f1be} /* (4, 25, 30) {real, imag} */,
  {32'hc0959131, 32'h40664a66} /* (4, 25, 29) {real, imag} */,
  {32'h3ed68204, 32'h407cdc56} /* (4, 25, 28) {real, imag} */,
  {32'hbe245276, 32'h4101a504} /* (4, 25, 27) {real, imag} */,
  {32'hbf016e98, 32'h41125cb6} /* (4, 25, 26) {real, imag} */,
  {32'hc06117c8, 32'h40abaf5f} /* (4, 25, 25) {real, imag} */,
  {32'hc00c791c, 32'h4038bf4f} /* (4, 25, 24) {real, imag} */,
  {32'hbe860814, 32'h4082ef2e} /* (4, 25, 23) {real, imag} */,
  {32'h3ee53bd4, 32'h40a5300d} /* (4, 25, 22) {real, imag} */,
  {32'h401eb90b, 32'h3fe43bed} /* (4, 25, 21) {real, imag} */,
  {32'h4064b7f4, 32'hc100116a} /* (4, 25, 20) {real, imag} */,
  {32'h3f5cced5, 32'hc100324b} /* (4, 25, 19) {real, imag} */,
  {32'h3f0e2af6, 32'hc0593e39} /* (4, 25, 18) {real, imag} */,
  {32'h3fda8bce, 32'hbfc881fb} /* (4, 25, 17) {real, imag} */,
  {32'h407f1270, 32'hc084330a} /* (4, 25, 16) {real, imag} */,
  {32'h3f29b61f, 32'hc0902648} /* (4, 25, 15) {real, imag} */,
  {32'hbf3204ac, 32'hc0ca1779} /* (4, 25, 14) {real, imag} */,
  {32'h3ec98a7a, 32'hc1045d61} /* (4, 25, 13) {real, imag} */,
  {32'h3f1401e6, 32'hc0ebbc4f} /* (4, 25, 12) {real, imag} */,
  {32'h3e81a4ed, 32'hc068939b} /* (4, 25, 11) {real, imag} */,
  {32'hbf84696c, 32'h3fc04698} /* (4, 25, 10) {real, imag} */,
  {32'hc0a4b30a, 32'h40977de6} /* (4, 25, 9) {real, imag} */,
  {32'hc07508df, 32'h40b65d29} /* (4, 25, 8) {real, imag} */,
  {32'hbeab72f6, 32'h40a0578a} /* (4, 25, 7) {real, imag} */,
  {32'hbe0b4f58, 32'h4063840e} /* (4, 25, 6) {real, imag} */,
  {32'hbf25cbaa, 32'h408c64da} /* (4, 25, 5) {real, imag} */,
  {32'hc02883ba, 32'h402846ce} /* (4, 25, 4) {real, imag} */,
  {32'hc033c344, 32'h404c9c8d} /* (4, 25, 3) {real, imag} */,
  {32'hbead1c86, 32'h406e262e} /* (4, 25, 2) {real, imag} */,
  {32'hbfa1bd32, 32'h40f280d4} /* (4, 25, 1) {real, imag} */,
  {32'hbf8f893a, 32'h408a629e} /* (4, 25, 0) {real, imag} */,
  {32'hbf6fe70a, 32'h40b03064} /* (4, 24, 31) {real, imag} */,
  {32'hbf2921ef, 32'h40c7ec20} /* (4, 24, 30) {real, imag} */,
  {32'hbfab73b4, 32'h406c7136} /* (4, 24, 29) {real, imag} */,
  {32'h3edf5b6e, 32'h409685ca} /* (4, 24, 28) {real, imag} */,
  {32'hbfc7b1ba, 32'h4026c2f8} /* (4, 24, 27) {real, imag} */,
  {32'hc0377e28, 32'h40d686ab} /* (4, 24, 26) {real, imag} */,
  {32'hc091dd84, 32'h40ef1046} /* (4, 24, 25) {real, imag} */,
  {32'hc05f876d, 32'h40d0375b} /* (4, 24, 24) {real, imag} */,
  {32'hbf24dfac, 32'h40eaa6ec} /* (4, 24, 23) {real, imag} */,
  {32'hbf96c9e6, 32'h41011bd1} /* (4, 24, 22) {real, imag} */,
  {32'hbf9ea10f, 32'h4039f105} /* (4, 24, 21) {real, imag} */,
  {32'h3fce41ec, 32'hc0becf6b} /* (4, 24, 20) {real, imag} */,
  {32'h3eea9b16, 32'hc09a42f4} /* (4, 24, 19) {real, imag} */,
  {32'h3fbb76a7, 32'hc054aff6} /* (4, 24, 18) {real, imag} */,
  {32'h4080c10f, 32'hc0a3bda8} /* (4, 24, 17) {real, imag} */,
  {32'h401dacf0, 32'hc09a09d2} /* (4, 24, 16) {real, imag} */,
  {32'hbd28e638, 32'hc05a4ca3} /* (4, 24, 15) {real, imag} */,
  {32'h404c733e, 32'hc0e83cb6} /* (4, 24, 14) {real, imag} */,
  {32'h4037bbe3, 32'hc10625d3} /* (4, 24, 13) {real, imag} */,
  {32'h3f7c02a8, 32'hc060e198} /* (4, 24, 12) {real, imag} */,
  {32'h3e23f470, 32'hbff20748} /* (4, 24, 11) {real, imag} */,
  {32'hbfea4ac2, 32'h40418c38} /* (4, 24, 10) {real, imag} */,
  {32'hc082fd76, 32'h40c5936e} /* (4, 24, 9) {real, imag} */,
  {32'hc095ff48, 32'h409ee504} /* (4, 24, 8) {real, imag} */,
  {32'hc03aeeec, 32'h4057d958} /* (4, 24, 7) {real, imag} */,
  {32'hbd833ff0, 32'h40442b3a} /* (4, 24, 6) {real, imag} */,
  {32'hbf11c679, 32'h40c1b09f} /* (4, 24, 5) {real, imag} */,
  {32'hbfd37f0e, 32'h40a8905e} /* (4, 24, 4) {real, imag} */,
  {32'hc023cb79, 32'h40ae6df0} /* (4, 24, 3) {real, imag} */,
  {32'hbf13da50, 32'h409d0a9c} /* (4, 24, 2) {real, imag} */,
  {32'hbf824eb2, 32'h40ecc0f4} /* (4, 24, 1) {real, imag} */,
  {32'hbf49ef68, 32'h40936584} /* (4, 24, 0) {real, imag} */,
  {32'hbf856529, 32'h408d8594} /* (4, 23, 31) {real, imag} */,
  {32'hbf257b7e, 32'h40b29cd6} /* (4, 23, 30) {real, imag} */,
  {32'hbf134114, 32'h40b242e9} /* (4, 23, 29) {real, imag} */,
  {32'hbf2baf05, 32'h409ef4c8} /* (4, 23, 28) {real, imag} */,
  {32'hc04fd332, 32'h401e6eb1} /* (4, 23, 27) {real, imag} */,
  {32'hc0bcc9ca, 32'h40a4bf30} /* (4, 23, 26) {real, imag} */,
  {32'hc0466fb0, 32'h40c99a8e} /* (4, 23, 25) {real, imag} */,
  {32'hbe99fae7, 32'h40a0108e} /* (4, 23, 24) {real, imag} */,
  {32'hbfdaa9a2, 32'h40b685ae} /* (4, 23, 23) {real, imag} */,
  {32'hc01057ed, 32'h40d906ca} /* (4, 23, 22) {real, imag} */,
  {32'hbe46fd90, 32'h404700da} /* (4, 23, 21) {real, imag} */,
  {32'h40157965, 32'hc03f5b5a} /* (4, 23, 20) {real, imag} */,
  {32'h3f750364, 32'hc007953c} /* (4, 23, 19) {real, imag} */,
  {32'h402d4c63, 32'hc02fd7e0} /* (4, 23, 18) {real, imag} */,
  {32'h4027655c, 32'hc0a85842} /* (4, 23, 17) {real, imag} */,
  {32'h3f9e9bee, 32'hc0c1e3fb} /* (4, 23, 16) {real, imag} */,
  {32'h40026fb4, 32'hc0b81080} /* (4, 23, 15) {real, imag} */,
  {32'h402209a2, 32'hc0e4d275} /* (4, 23, 14) {real, imag} */,
  {32'h3f2be564, 32'hc0d8c63d} /* (4, 23, 13) {real, imag} */,
  {32'h3f31c713, 32'hc0533152} /* (4, 23, 12) {real, imag} */,
  {32'h3fb3247c, 32'hc01bfeb2} /* (4, 23, 11) {real, imag} */,
  {32'h3f877d8a, 32'h3f819d98} /* (4, 23, 10) {real, imag} */,
  {32'h3c866b70, 32'h408a86cd} /* (4, 23, 9) {real, imag} */,
  {32'hc023eb7f, 32'h408e00da} /* (4, 23, 8) {real, imag} */,
  {32'hbf9c9340, 32'h400bf10b} /* (4, 23, 7) {real, imag} */,
  {32'hbe76d970, 32'h40513e52} /* (4, 23, 6) {real, imag} */,
  {32'hbf4beec5, 32'h40ee7801} /* (4, 23, 5) {real, imag} */,
  {32'hbebd4834, 32'h409da75c} /* (4, 23, 4) {real, imag} */,
  {32'h3feaea31, 32'h406b0a30} /* (4, 23, 3) {real, imag} */,
  {32'hbe9a50d9, 32'h40b10610} /* (4, 23, 2) {real, imag} */,
  {32'hbff43eba, 32'h40b5def8} /* (4, 23, 1) {real, imag} */,
  {32'hbfad80cd, 32'h40519d5b} /* (4, 23, 0) {real, imag} */,
  {32'hc04f5c96, 32'h40630b19} /* (4, 22, 31) {real, imag} */,
  {32'hbfbf13a2, 32'h40788804} /* (4, 22, 30) {real, imag} */,
  {32'hbf35d336, 32'h409c72ea} /* (4, 22, 29) {real, imag} */,
  {32'hc007d5d8, 32'h40d48d26} /* (4, 22, 28) {real, imag} */,
  {32'hbfcc8be0, 32'h410085a0} /* (4, 22, 27) {real, imag} */,
  {32'hc0308f7a, 32'h40ad62e5} /* (4, 22, 26) {real, imag} */,
  {32'hbf8e92c8, 32'h40421cef} /* (4, 22, 25) {real, imag} */,
  {32'hbe85756e, 32'h40959b15} /* (4, 22, 24) {real, imag} */,
  {32'hbf837aa1, 32'h40e5b0ac} /* (4, 22, 23) {real, imag} */,
  {32'hc05b26a7, 32'h40dcda19} /* (4, 22, 22) {real, imag} */,
  {32'h3f2fe722, 32'h4053de04} /* (4, 22, 21) {real, imag} */,
  {32'h4071e552, 32'h3f15256a} /* (4, 22, 20) {real, imag} */,
  {32'h3f9c7d00, 32'h3f185e81} /* (4, 22, 19) {real, imag} */,
  {32'h3fd75238, 32'hbfdfcaa8} /* (4, 22, 18) {real, imag} */,
  {32'h3f9314ac, 32'hc0c519e7} /* (4, 22, 17) {real, imag} */,
  {32'h3fd433fd, 32'hc0d0f9ae} /* (4, 22, 16) {real, imag} */,
  {32'h3fc57ba9, 32'hc0c17e48} /* (4, 22, 15) {real, imag} */,
  {32'hbb4733c0, 32'hc0c3b0f6} /* (4, 22, 14) {real, imag} */,
  {32'h3ff40b98, 32'hc0ac474d} /* (4, 22, 13) {real, imag} */,
  {32'h404ce806, 32'hc0bf7bc2} /* (4, 22, 12) {real, imag} */,
  {32'h407bcae6, 32'hc0913555} /* (4, 22, 11) {real, imag} */,
  {32'h404d96d0, 32'h40010cec} /* (4, 22, 10) {real, imag} */,
  {32'hbecf8556, 32'h40ff9e2a} /* (4, 22, 9) {real, imag} */,
  {32'hbfc8b5ed, 32'h4113ccfc} /* (4, 22, 8) {real, imag} */,
  {32'hbfe97b96, 32'h40cab56b} /* (4, 22, 7) {real, imag} */,
  {32'hbf52bac6, 32'h4070eea1} /* (4, 22, 6) {real, imag} */,
  {32'hbef83099, 32'h40e3c8fc} /* (4, 22, 5) {real, imag} */,
  {32'hbeecec14, 32'h409cf7db} /* (4, 22, 4) {real, imag} */,
  {32'h3f56f27c, 32'h3fbc6ef2} /* (4, 22, 3) {real, imag} */,
  {32'hbe98295a, 32'h40977c84} /* (4, 22, 2) {real, imag} */,
  {32'hbf95ccb2, 32'h4072bfe8} /* (4, 22, 1) {real, imag} */,
  {32'hc00fae0a, 32'h3ffad31e} /* (4, 22, 0) {real, imag} */,
  {32'hbf86d980, 32'h4026f694} /* (4, 21, 31) {real, imag} */,
  {32'hbf2e52ff, 32'h40858314} /* (4, 21, 30) {real, imag} */,
  {32'hc0199b30, 32'h3fdb6894} /* (4, 21, 29) {real, imag} */,
  {32'hc05817fe, 32'h40578f66} /* (4, 21, 28) {real, imag} */,
  {32'hbf8ab0bc, 32'h40d58741} /* (4, 21, 27) {real, imag} */,
  {32'h3fcccf00, 32'h405159dc} /* (4, 21, 26) {real, imag} */,
  {32'hbe807315, 32'h3fb9d74c} /* (4, 21, 25) {real, imag} */,
  {32'hc051f121, 32'h4057cd55} /* (4, 21, 24) {real, imag} */,
  {32'h3f516faf, 32'h408b8716} /* (4, 21, 23) {real, imag} */,
  {32'hbe0c3ff1, 32'h40113750} /* (4, 21, 22) {real, imag} */,
  {32'hbf20065e, 32'hbf40e47c} /* (4, 21, 21) {real, imag} */,
  {32'hbe3c72af, 32'h3f781422} /* (4, 21, 20) {real, imag} */,
  {32'hbfb34cd4, 32'h3f4306ca} /* (4, 21, 19) {real, imag} */,
  {32'hbe9527c0, 32'hc00ca6b6} /* (4, 21, 18) {real, imag} */,
  {32'h3f07751a, 32'hc09c8d9c} /* (4, 21, 17) {real, imag} */,
  {32'h3fe89a26, 32'hc09f54f0} /* (4, 21, 16) {real, imag} */,
  {32'h3f3fe40e, 32'hc02bbe4a} /* (4, 21, 15) {real, imag} */,
  {32'hbf5c44a5, 32'hbfbb9d47} /* (4, 21, 14) {real, imag} */,
  {32'h3f8d7080, 32'hbfae431c} /* (4, 21, 13) {real, imag} */,
  {32'h3fda3c8c, 32'hbebd6096} /* (4, 21, 12) {real, imag} */,
  {32'h3dfeab74, 32'hbb862fc0} /* (4, 21, 11) {real, imag} */,
  {32'hbee60ea4, 32'h3fbd814d} /* (4, 21, 10) {real, imag} */,
  {32'hbfda77f2, 32'h4104b877} /* (4, 21, 9) {real, imag} */,
  {32'hc00a23b7, 32'h4102e422} /* (4, 21, 8) {real, imag} */,
  {32'hbfce30c7, 32'h4089764b} /* (4, 21, 7) {real, imag} */,
  {32'hbed94aa3, 32'hbf7c2a1f} /* (4, 21, 6) {real, imag} */,
  {32'hbfa85e3c, 32'hbf34f66d} /* (4, 21, 5) {real, imag} */,
  {32'hbfacddda, 32'h3feef9dc} /* (4, 21, 4) {real, imag} */,
  {32'hbf8b2bd6, 32'h3f44af87} /* (4, 21, 3) {real, imag} */,
  {32'hbe02090e, 32'h3ef73d12} /* (4, 21, 2) {real, imag} */,
  {32'hbd1d5630, 32'h3f88c5aa} /* (4, 21, 1) {real, imag} */,
  {32'hbf4242ea, 32'h3d221440} /* (4, 21, 0) {real, imag} */,
  {32'h3f195046, 32'hbf484645} /* (4, 20, 31) {real, imag} */,
  {32'h3e9346e2, 32'h3f85a9fd} /* (4, 20, 30) {real, imag} */,
  {32'hbf122617, 32'hc04a9985} /* (4, 20, 29) {real, imag} */,
  {32'hbf6f7e65, 32'hc0bb60f4} /* (4, 20, 28) {real, imag} */,
  {32'hc00543ad, 32'hc07549b2} /* (4, 20, 27) {real, imag} */,
  {32'h3fa01c37, 32'hc0299cac} /* (4, 20, 26) {real, imag} */,
  {32'h40169192, 32'hc03c928d} /* (4, 20, 25) {real, imag} */,
  {32'h3eef75a2, 32'hc070a94a} /* (4, 20, 24) {real, imag} */,
  {32'h3ff24446, 32'hc0bc48f0} /* (4, 20, 23) {real, imag} */,
  {32'h40815946, 32'hc0b2fbac} /* (4, 20, 22) {real, imag} */,
  {32'h3f18fdc5, 32'hc00d48df} /* (4, 20, 21) {real, imag} */,
  {32'hc005cdfd, 32'h402ae7c6} /* (4, 20, 20) {real, imag} */,
  {32'hc07ddc20, 32'h3fe6fb64} /* (4, 20, 19) {real, imag} */,
  {32'hc06ba4bf, 32'h3fe094ad} /* (4, 20, 18) {real, imag} */,
  {32'hbfec15ea, 32'hbe794bf4} /* (4, 20, 17) {real, imag} */,
  {32'hc008f951, 32'hbf3f44ff} /* (4, 20, 16) {real, imag} */,
  {32'hc0240404, 32'h40847555} /* (4, 20, 15) {real, imag} */,
  {32'hbf8c0851, 32'h40cc8308} /* (4, 20, 14) {real, imag} */,
  {32'h3f820389, 32'h409b94f6} /* (4, 20, 13) {real, imag} */,
  {32'h3f17410f, 32'h40d2bb36} /* (4, 20, 12) {real, imag} */,
  {32'hbfb6134f, 32'h40a8d832} /* (4, 20, 11) {real, imag} */,
  {32'hc008d79f, 32'hbe6eaab7} /* (4, 20, 10) {real, imag} */,
  {32'h3f940372, 32'h3e22c148} /* (4, 20, 9) {real, imag} */,
  {32'h3fb9f7cb, 32'hc0529b25} /* (4, 20, 8) {real, imag} */,
  {32'h3eb95997, 32'hc0a9431e} /* (4, 20, 7) {real, imag} */,
  {32'h3f001623, 32'hc0b1bc02} /* (4, 20, 6) {real, imag} */,
  {32'h3f0f8a65, 32'hc0491458} /* (4, 20, 5) {real, imag} */,
  {32'h3f8d12ca, 32'hc0510e5c} /* (4, 20, 4) {real, imag} */,
  {32'h3fb2834f, 32'hc085aeb2} /* (4, 20, 3) {real, imag} */,
  {32'h40358db0, 32'hc0a3ab8c} /* (4, 20, 2) {real, imag} */,
  {32'h3fe12170, 32'hc076e4b9} /* (4, 20, 1) {real, imag} */,
  {32'h3f4b62a3, 32'hc048607a} /* (4, 20, 0) {real, imag} */,
  {32'h3fd8f79d, 32'hbffca8ad} /* (4, 19, 31) {real, imag} */,
  {32'h402b927d, 32'hbfc47ab4} /* (4, 19, 30) {real, imag} */,
  {32'h3fd26972, 32'hc04d1f44} /* (4, 19, 29) {real, imag} */,
  {32'hc0114250, 32'hc0b9cd5c} /* (4, 19, 28) {real, imag} */,
  {32'hbe41540e, 32'hc0ccac62} /* (4, 19, 27) {real, imag} */,
  {32'h3f92ff1c, 32'hc0a86a4e} /* (4, 19, 26) {real, imag} */,
  {32'h3e9f85ae, 32'hc0edb42a} /* (4, 19, 25) {real, imag} */,
  {32'h3e922ae7, 32'hc0ef8a1e} /* (4, 19, 24) {real, imag} */,
  {32'h402a8cb7, 32'hc0e6680d} /* (4, 19, 23) {real, imag} */,
  {32'h409b5e3c, 32'hc0bcd85f} /* (4, 19, 22) {real, imag} */,
  {32'h405e5822, 32'hbfaa3b94} /* (4, 19, 21) {real, imag} */,
  {32'h3f225fb6, 32'h40ac6ca1} /* (4, 19, 20) {real, imag} */,
  {32'hbf8a1ed8, 32'h40d6bcdc} /* (4, 19, 19) {real, imag} */,
  {32'hbfa246ba, 32'h40fc0577} /* (4, 19, 18) {real, imag} */,
  {32'h3fb4f2d8, 32'h40a84ee5} /* (4, 19, 17) {real, imag} */,
  {32'h3ef61188, 32'h3efdfc43} /* (4, 19, 16) {real, imag} */,
  {32'hbe3e73d8, 32'h402fa427} /* (4, 19, 15) {real, imag} */,
  {32'h3f8d4f65, 32'h407eaf27} /* (4, 19, 14) {real, imag} */,
  {32'h400194ed, 32'h40952e8a} /* (4, 19, 13) {real, imag} */,
  {32'h3e43d0a8, 32'h40ecd1ee} /* (4, 19, 12) {real, imag} */,
  {32'hbfc1436e, 32'h40b9dc85} /* (4, 19, 11) {real, imag} */,
  {32'hbe2d29c4, 32'hc0060f48} /* (4, 19, 10) {real, imag} */,
  {32'h3f365377, 32'hc0a835ba} /* (4, 19, 9) {real, imag} */,
  {32'hbe4172ea, 32'hc104071c} /* (4, 19, 8) {real, imag} */,
  {32'h3fc3e328, 32'hc0f85663} /* (4, 19, 7) {real, imag} */,
  {32'h3fedbc78, 32'hc0093458} /* (4, 19, 6) {real, imag} */,
  {32'h408d83c8, 32'hbe55b1d0} /* (4, 19, 5) {real, imag} */,
  {32'h401cf4aa, 32'hc07f3e7a} /* (4, 19, 4) {real, imag} */,
  {32'h3e0340aa, 32'hc09bb1c1} /* (4, 19, 3) {real, imag} */,
  {32'h40476878, 32'hc09983d2} /* (4, 19, 2) {real, imag} */,
  {32'h4021157a, 32'hc0e62c16} /* (4, 19, 1) {real, imag} */,
  {32'h3fe43afd, 32'hc0a2221b} /* (4, 19, 0) {real, imag} */,
  {32'h3f8f60c8, 32'hc07ee72b} /* (4, 18, 31) {real, imag} */,
  {32'h401597a8, 32'hc08dc00e} /* (4, 18, 30) {real, imag} */,
  {32'h403e7efe, 32'hbfc16ac4} /* (4, 18, 29) {real, imag} */,
  {32'h3f959319, 32'hbfadb0a4} /* (4, 18, 28) {real, imag} */,
  {32'h40636dcc, 32'hc08d502c} /* (4, 18, 27) {real, imag} */,
  {32'h4045450d, 32'hc0aacbcb} /* (4, 18, 26) {real, imag} */,
  {32'h3f742d54, 32'hc09fb03b} /* (4, 18, 25) {real, imag} */,
  {32'h3fc8d634, 32'hc0ac40c8} /* (4, 18, 24) {real, imag} */,
  {32'h403c5948, 32'hc08d025e} /* (4, 18, 23) {real, imag} */,
  {32'h4099ee2e, 32'hc0742e95} /* (4, 18, 22) {real, imag} */,
  {32'h409d3f51, 32'hbdc9c858} /* (4, 18, 21) {real, imag} */,
  {32'h3fda04a6, 32'h40cb9846} /* (4, 18, 20) {real, imag} */,
  {32'hbfff6f9c, 32'h40dc69ac} /* (4, 18, 19) {real, imag} */,
  {32'hc059d9fa, 32'h40e4b872} /* (4, 18, 18) {real, imag} */,
  {32'h3f804285, 32'h40efed22} /* (4, 18, 17) {real, imag} */,
  {32'h4089780f, 32'h4014a00c} /* (4, 18, 16) {real, imag} */,
  {32'h4019b0ac, 32'h3faccb05} /* (4, 18, 15) {real, imag} */,
  {32'h3e5ba62a, 32'h4066c0bc} /* (4, 18, 14) {real, imag} */,
  {32'hbf867339, 32'h40aded96} /* (4, 18, 13) {real, imag} */,
  {32'h3f956954, 32'h40ba0d74} /* (4, 18, 12) {real, imag} */,
  {32'hbe8e8470, 32'h409f22f4} /* (4, 18, 11) {real, imag} */,
  {32'h3ff72bfc, 32'hc06a1f90} /* (4, 18, 10) {real, imag} */,
  {32'h40303042, 32'hc105f7fe} /* (4, 18, 9) {real, imag} */,
  {32'h3c0d4558, 32'hc0dc7d48} /* (4, 18, 8) {real, imag} */,
  {32'h3fa4e7a2, 32'hc092a322} /* (4, 18, 7) {real, imag} */,
  {32'h3ff88099, 32'hbf8f8be9} /* (4, 18, 6) {real, imag} */,
  {32'h3ffc2836, 32'hbea030f0} /* (4, 18, 5) {real, imag} */,
  {32'h3f74c3b0, 32'hc061ffee} /* (4, 18, 4) {real, imag} */,
  {32'h3e5d8734, 32'hc0775aae} /* (4, 18, 3) {real, imag} */,
  {32'h4031b714, 32'hc08972b1} /* (4, 18, 2) {real, imag} */,
  {32'h3f23ce58, 32'hc0971cb3} /* (4, 18, 1) {real, imag} */,
  {32'h3e6edea8, 32'hc094d72c} /* (4, 18, 0) {real, imag} */,
  {32'h3f06d937, 32'hc06c9fa4} /* (4, 17, 31) {real, imag} */,
  {32'h3f137066, 32'hc0cdc758} /* (4, 17, 30) {real, imag} */,
  {32'h403df83c, 32'hc0900445} /* (4, 17, 29) {real, imag} */,
  {32'h4098c18a, 32'hc0234d47} /* (4, 17, 28) {real, imag} */,
  {32'h4020c2f2, 32'hc0c8c232} /* (4, 17, 27) {real, imag} */,
  {32'h3fa81de1, 32'hc0c5c5c7} /* (4, 17, 26) {real, imag} */,
  {32'h402180fc, 32'hc05b752a} /* (4, 17, 25) {real, imag} */,
  {32'h4077620a, 32'hc02b90e1} /* (4, 17, 24) {real, imag} */,
  {32'h4098f478, 32'hc04605bd} /* (4, 17, 23) {real, imag} */,
  {32'h40946642, 32'hc0adb354} /* (4, 17, 22) {real, imag} */,
  {32'h40a1e6ac, 32'hbe38d06a} /* (4, 17, 21) {real, imag} */,
  {32'h3f8f7544, 32'h40b04e16} /* (4, 17, 20) {real, imag} */,
  {32'hbf7718fc, 32'h406cafb7} /* (4, 17, 19) {real, imag} */,
  {32'hc0189e97, 32'h3faabdbe} /* (4, 17, 18) {real, imag} */,
  {32'hc024bf76, 32'h40ad03fc} /* (4, 17, 17) {real, imag} */,
  {32'h3f127b28, 32'h40b3a1a8} /* (4, 17, 16) {real, imag} */,
  {32'hbf2694f3, 32'h408504ed} /* (4, 17, 15) {real, imag} */,
  {32'hc0866a12, 32'h404010ff} /* (4, 17, 14) {real, imag} */,
  {32'hc06a99e2, 32'h40556404} /* (4, 17, 13) {real, imag} */,
  {32'hc026733c, 32'h4086c80f} /* (4, 17, 12) {real, imag} */,
  {32'hbf5646bc, 32'h4000e5a0} /* (4, 17, 11) {real, imag} */,
  {32'h3f980bfa, 32'hc0bb046c} /* (4, 17, 10) {real, imag} */,
  {32'h40224060, 32'hc0dd5b91} /* (4, 17, 9) {real, imag} */,
  {32'h3fdcc6ad, 32'hc0951a4a} /* (4, 17, 8) {real, imag} */,
  {32'h405c5578, 32'hc0aca6ca} /* (4, 17, 7) {real, imag} */,
  {32'h4010473e, 32'hc0cfb23c} /* (4, 17, 6) {real, imag} */,
  {32'hc0337f36, 32'hc08358da} /* (4, 17, 5) {real, imag} */,
  {32'hbf984851, 32'hc0863d52} /* (4, 17, 4) {real, imag} */,
  {32'h3e854cb2, 32'hbfd15608} /* (4, 17, 3) {real, imag} */,
  {32'hbffc3f47, 32'h3f0935f7} /* (4, 17, 2) {real, imag} */,
  {32'hc00a2801, 32'hbfd5516c} /* (4, 17, 1) {real, imag} */,
  {32'h3f0a5755, 32'hc05d71fc} /* (4, 17, 0) {real, imag} */,
  {32'hbf101bea, 32'hc0022428} /* (4, 16, 31) {real, imag} */,
  {32'h3da94208, 32'hc0a01d1a} /* (4, 16, 30) {real, imag} */,
  {32'h40340356, 32'hc0bb55f2} /* (4, 16, 29) {real, imag} */,
  {32'h4067fe3b, 32'hc059a41a} /* (4, 16, 28) {real, imag} */,
  {32'h3fdcb534, 32'hc0a2431e} /* (4, 16, 27) {real, imag} */,
  {32'h3ede4ca4, 32'hc08d8f76} /* (4, 16, 26) {real, imag} */,
  {32'h3f8ac3bd, 32'hc075dc87} /* (4, 16, 25) {real, imag} */,
  {32'h403ab86f, 32'hc0bd5cd0} /* (4, 16, 24) {real, imag} */,
  {32'h4083f552, 32'hc082db37} /* (4, 16, 23) {real, imag} */,
  {32'h405ed41c, 32'hc0c52915} /* (4, 16, 22) {real, imag} */,
  {32'h4004d860, 32'hc035a2c9} /* (4, 16, 21) {real, imag} */,
  {32'hbf6e7eac, 32'h40ab0fd5} /* (4, 16, 20) {real, imag} */,
  {32'hbf659db8, 32'h40c37966} /* (4, 16, 19) {real, imag} */,
  {32'h3f7a54ea, 32'h405e4636} /* (4, 16, 18) {real, imag} */,
  {32'hbffd56bc, 32'h40c7da92} /* (4, 16, 17) {real, imag} */,
  {32'hc013760e, 32'h40c4291a} /* (4, 16, 16) {real, imag} */,
  {32'hbf3729b1, 32'h40d7f1fa} /* (4, 16, 15) {real, imag} */,
  {32'hc03ecbd2, 32'h409eacbe} /* (4, 16, 14) {real, imag} */,
  {32'hc0460af2, 32'h408cd396} /* (4, 16, 13) {real, imag} */,
  {32'hc0941c2a, 32'h4093b986} /* (4, 16, 12) {real, imag} */,
  {32'hbfb900a4, 32'h40212c86} /* (4, 16, 11) {real, imag} */,
  {32'h3f8947e2, 32'hc0743fd6} /* (4, 16, 10) {real, imag} */,
  {32'h4023c67c, 32'hc0a5627e} /* (4, 16, 9) {real, imag} */,
  {32'h3feae2b6, 32'hc0a923f6} /* (4, 16, 8) {real, imag} */,
  {32'h4056827e, 32'hc1099040} /* (4, 16, 7) {real, imag} */,
  {32'h4021b516, 32'hc1103d3a} /* (4, 16, 6) {real, imag} */,
  {32'h3d373cbc, 32'hc0a05c77} /* (4, 16, 5) {real, imag} */,
  {32'h3faea607, 32'hc03f10f3} /* (4, 16, 4) {real, imag} */,
  {32'h3f575fb4, 32'hc03c448d} /* (4, 16, 3) {real, imag} */,
  {32'hbf8a6e31, 32'hc06c0fa4} /* (4, 16, 2) {real, imag} */,
  {32'h3f99f5d8, 32'hc0b6aa04} /* (4, 16, 1) {real, imag} */,
  {32'h3fc841d0, 32'hc0706166} /* (4, 16, 0) {real, imag} */,
  {32'hbf9f3f0b, 32'hbff0f968} /* (4, 15, 31) {real, imag} */,
  {32'hbf84d7f7, 32'hc0382a5d} /* (4, 15, 30) {real, imag} */,
  {32'h3f8709b8, 32'hc08fd70c} /* (4, 15, 29) {real, imag} */,
  {32'h4016c760, 32'hc0ae988c} /* (4, 15, 28) {real, imag} */,
  {32'h3fe16804, 32'hc0a1dbe7} /* (4, 15, 27) {real, imag} */,
  {32'h3d88419c, 32'hc066415a} /* (4, 15, 26) {real, imag} */,
  {32'hbfd46514, 32'hc05d0c36} /* (4, 15, 25) {real, imag} */,
  {32'hbf2d20ba, 32'hc0972c15} /* (4, 15, 24) {real, imag} */,
  {32'h3f48a65f, 32'hc0aee574} /* (4, 15, 23) {real, imag} */,
  {32'h3f010900, 32'hc0d570e2} /* (4, 15, 22) {real, imag} */,
  {32'hbedd8aeb, 32'hc0a7c5ed} /* (4, 15, 21) {real, imag} */,
  {32'hbfa4a130, 32'h3fbcebce} /* (4, 15, 20) {real, imag} */,
  {32'hbf9eb5ab, 32'h40d12f7a} /* (4, 15, 19) {real, imag} */,
  {32'h3f32437a, 32'h40a5d2a0} /* (4, 15, 18) {real, imag} */,
  {32'hbefdac28, 32'h40bf4332} /* (4, 15, 17) {real, imag} */,
  {32'hbfe89059, 32'h40d92264} /* (4, 15, 16) {real, imag} */,
  {32'hbf3d4459, 32'h40ceb5dc} /* (4, 15, 15) {real, imag} */,
  {32'hbf739b16, 32'h40e84ad4} /* (4, 15, 14) {real, imag} */,
  {32'h3f2448c3, 32'h4094ce2a} /* (4, 15, 13) {real, imag} */,
  {32'hbfe48c60, 32'h403a167a} /* (4, 15, 12) {real, imag} */,
  {32'hbf0ae2b8, 32'h4017fafa} /* (4, 15, 11) {real, imag} */,
  {32'h3fdd1d46, 32'hc04f35dc} /* (4, 15, 10) {real, imag} */,
  {32'h40032ec6, 32'hc09b6288} /* (4, 15, 9) {real, imag} */,
  {32'h3fd9eacc, 32'hc09ba0e2} /* (4, 15, 8) {real, imag} */,
  {32'h4039b959, 32'hc0fbd5ef} /* (4, 15, 7) {real, imag} */,
  {32'h406e9acc, 32'hc0d4e2f2} /* (4, 15, 6) {real, imag} */,
  {32'h4004932e, 32'hc08bbaeb} /* (4, 15, 5) {real, imag} */,
  {32'h4013a4f3, 32'hc00b2602} /* (4, 15, 4) {real, imag} */,
  {32'h3fe3d24c, 32'hc058c6b5} /* (4, 15, 3) {real, imag} */,
  {32'h3f9dfc81, 32'hc0c99c92} /* (4, 15, 2) {real, imag} */,
  {32'h3fce52cf, 32'hc0d4468d} /* (4, 15, 1) {real, imag} */,
  {32'h3feac00c, 32'hc0551500} /* (4, 15, 0) {real, imag} */,
  {32'h3f18cd8b, 32'hbff14911} /* (4, 14, 31) {real, imag} */,
  {32'h3fd611f8, 32'hc01ac97c} /* (4, 14, 30) {real, imag} */,
  {32'h3fd4676e, 32'hc0b52a2e} /* (4, 14, 29) {real, imag} */,
  {32'hbf8c15f8, 32'hc0d185f8} /* (4, 14, 28) {real, imag} */,
  {32'hbe8d56f2, 32'hc091e0e5} /* (4, 14, 27) {real, imag} */,
  {32'hbe3cd9e4, 32'hc031ff92} /* (4, 14, 26) {real, imag} */,
  {32'hbfb0a2ae, 32'hc020f3b6} /* (4, 14, 25) {real, imag} */,
  {32'h4028858d, 32'hc0606eae} /* (4, 14, 24) {real, imag} */,
  {32'h408480bf, 32'hc08cbb6e} /* (4, 14, 23) {real, imag} */,
  {32'h3f1b1f58, 32'hc0c15e56} /* (4, 14, 22) {real, imag} */,
  {32'hbff27688, 32'hc06039b2} /* (4, 14, 21) {real, imag} */,
  {32'hbea45f68, 32'h403d8e24} /* (4, 14, 20) {real, imag} */,
  {32'hc08224f8, 32'h40b29e1c} /* (4, 14, 19) {real, imag} */,
  {32'hc04c5584, 32'h4094774e} /* (4, 14, 18) {real, imag} */,
  {32'hbf2bb8b0, 32'h4099c866} /* (4, 14, 17) {real, imag} */,
  {32'hbfa55495, 32'h40fd4fa7} /* (4, 14, 16) {real, imag} */,
  {32'hbf3795ec, 32'h40d72160} /* (4, 14, 15) {real, imag} */,
  {32'hc02e12c6, 32'h40ef9bad} /* (4, 14, 14) {real, imag} */,
  {32'hbfa73d30, 32'h40a334ae} /* (4, 14, 13) {real, imag} */,
  {32'hc01a8eac, 32'h3fdbb394} /* (4, 14, 12) {real, imag} */,
  {32'hbfa04b10, 32'h3f9acbc0} /* (4, 14, 11) {real, imag} */,
  {32'h3fc63c73, 32'hc0913361} /* (4, 14, 10) {real, imag} */,
  {32'h3ec4d3ea, 32'hc0b00efe} /* (4, 14, 9) {real, imag} */,
  {32'hbe0a9ac4, 32'hc081a47f} /* (4, 14, 8) {real, imag} */,
  {32'h3fc53bd4, 32'hc09a530e} /* (4, 14, 7) {real, imag} */,
  {32'h3fc3a150, 32'hc0acac57} /* (4, 14, 6) {real, imag} */,
  {32'h3fb86d70, 32'hc0944764} /* (4, 14, 5) {real, imag} */,
  {32'h4065beef, 32'hc06f9877} /* (4, 14, 4) {real, imag} */,
  {32'h409f44c4, 32'hc0d637c6} /* (4, 14, 3) {real, imag} */,
  {32'h403bffea, 32'hc0f42494} /* (4, 14, 2) {real, imag} */,
  {32'h3f944ca2, 32'hc06f3bfc} /* (4, 14, 1) {real, imag} */,
  {32'h3fd2909a, 32'hbf34bd1e} /* (4, 14, 0) {real, imag} */,
  {32'h4016d642, 32'hbfef3c45} /* (4, 13, 31) {real, imag} */,
  {32'h40719df4, 32'hc0b777d6} /* (4, 13, 30) {real, imag} */,
  {32'h405b031e, 32'hc0dba3dc} /* (4, 13, 29) {real, imag} */,
  {32'h3ff2a66a, 32'hc0e11c2b} /* (4, 13, 28) {real, imag} */,
  {32'h3ecf4a78, 32'hc0a8dcca} /* (4, 13, 27) {real, imag} */,
  {32'hbe50d8b8, 32'hc064030b} /* (4, 13, 26) {real, imag} */,
  {32'h404edbb2, 32'hc0ae1bde} /* (4, 13, 25) {real, imag} */,
  {32'h4083c9c6, 32'hc0f2e9a4} /* (4, 13, 24) {real, imag} */,
  {32'h4017007a, 32'hc09ee4ac} /* (4, 13, 23) {real, imag} */,
  {32'hbf9788c2, 32'hc073e05b} /* (4, 13, 22) {real, imag} */,
  {32'hbfd73af2, 32'hc023f1b9} /* (4, 13, 21) {real, imag} */,
  {32'h3f386c74, 32'h4047b682} /* (4, 13, 20) {real, imag} */,
  {32'hc039c226, 32'h407be793} /* (4, 13, 19) {real, imag} */,
  {32'hc09fde33, 32'h3f8d8c0b} /* (4, 13, 18) {real, imag} */,
  {32'hc01a81aa, 32'h409e8817} /* (4, 13, 17) {real, imag} */,
  {32'hbffaa4a5, 32'h41062e90} /* (4, 13, 16) {real, imag} */,
  {32'hbfafc154, 32'h4100dc1f} /* (4, 13, 15) {real, imag} */,
  {32'hbf2a9c16, 32'h40f8ce13} /* (4, 13, 14) {real, imag} */,
  {32'h3f603c69, 32'h40919955} /* (4, 13, 13) {real, imag} */,
  {32'hbfdd997c, 32'h402c5656} /* (4, 13, 12) {real, imag} */,
  {32'hc00aec5c, 32'h3f319418} /* (4, 13, 11) {real, imag} */,
  {32'h3fec85a8, 32'hc0886c58} /* (4, 13, 10) {real, imag} */,
  {32'h3fdcc792, 32'hc0aaafd8} /* (4, 13, 9) {real, imag} */,
  {32'h3ff65524, 32'hc0a27734} /* (4, 13, 8) {real, imag} */,
  {32'h40577191, 32'hc09ea676} /* (4, 13, 7) {real, imag} */,
  {32'h3f9aa62a, 32'hc0a0f17c} /* (4, 13, 6) {real, imag} */,
  {32'h3f5317ca, 32'hc0af46eb} /* (4, 13, 5) {real, imag} */,
  {32'h404f824e, 32'hc0b0957e} /* (4, 13, 4) {real, imag} */,
  {32'h40a6c779, 32'hc0ff7f2a} /* (4, 13, 3) {real, imag} */,
  {32'h4020d361, 32'hc0d1b175} /* (4, 13, 2) {real, imag} */,
  {32'hbd35bcd0, 32'hc051011c} /* (4, 13, 1) {real, imag} */,
  {32'hbe89e5fe, 32'hbfc78322} /* (4, 13, 0) {real, imag} */,
  {32'h40778010, 32'hbfdf719d} /* (4, 12, 31) {real, imag} */,
  {32'h408e5bb6, 32'hc0bc539a} /* (4, 12, 30) {real, imag} */,
  {32'h403bd002, 32'hc0e3bf1b} /* (4, 12, 29) {real, imag} */,
  {32'h4056f851, 32'hc0ccef86} /* (4, 12, 28) {real, imag} */,
  {32'h400893b8, 32'hc0baff12} /* (4, 12, 27) {real, imag} */,
  {32'h4021622d, 32'hc0a3d2f0} /* (4, 12, 26) {real, imag} */,
  {32'h406e88b3, 32'hc0e89c98} /* (4, 12, 25) {real, imag} */,
  {32'h4085a2f8, 32'hc0f8ad7f} /* (4, 12, 24) {real, imag} */,
  {32'h4010eb3f, 32'hc0a454b1} /* (4, 12, 23) {real, imag} */,
  {32'h3f0ed524, 32'hc080be71} /* (4, 12, 22) {real, imag} */,
  {32'h3fb563ed, 32'hc052c9c9} /* (4, 12, 21) {real, imag} */,
  {32'hbf010075, 32'h4054ba3c} /* (4, 12, 20) {real, imag} */,
  {32'hc0bf76db, 32'h40aeff4e} /* (4, 12, 19) {real, imag} */,
  {32'hc0f55e8d, 32'h40333e07} /* (4, 12, 18) {real, imag} */,
  {32'hc095bb62, 32'h40b1656c} /* (4, 12, 17) {real, imag} */,
  {32'hc0860537, 32'h40e55258} /* (4, 12, 16) {real, imag} */,
  {32'hc015f434, 32'h40d854c0} /* (4, 12, 15) {real, imag} */,
  {32'h3f5c4630, 32'h40abe1b4} /* (4, 12, 14) {real, imag} */,
  {32'h3fbd3641, 32'h40ad4589} /* (4, 12, 13) {real, imag} */,
  {32'hbfdefc0f, 32'h4104e4c2} /* (4, 12, 12) {real, imag} */,
  {32'hc06a044c, 32'h40c1be48} /* (4, 12, 11) {real, imag} */,
  {32'h3e839cf3, 32'hbe8fc052} /* (4, 12, 10) {real, imag} */,
  {32'h3fa470b2, 32'hc0881fda} /* (4, 12, 9) {real, imag} */,
  {32'h40050388, 32'hc0b6beb6} /* (4, 12, 8) {real, imag} */,
  {32'h404b334e, 32'hc0aa04d5} /* (4, 12, 7) {real, imag} */,
  {32'h408f687c, 32'hc0a2f794} /* (4, 12, 6) {real, imag} */,
  {32'h40912b0e, 32'hc067530e} /* (4, 12, 5) {real, imag} */,
  {32'h400bae76, 32'hc053c7a0} /* (4, 12, 4) {real, imag} */,
  {32'h407e6900, 32'hc0c8ce92} /* (4, 12, 3) {real, imag} */,
  {32'h40b5f4c0, 32'hc0be396a} /* (4, 12, 2) {real, imag} */,
  {32'h408c5f0c, 32'hc0c05424} /* (4, 12, 1) {real, imag} */,
  {32'h3feeb9ec, 32'hc08571ff} /* (4, 12, 0) {real, imag} */,
  {32'h401a521e, 32'hbf67dde6} /* (4, 11, 31) {real, imag} */,
  {32'h3ff04cfe, 32'hc0736f2e} /* (4, 11, 30) {real, imag} */,
  {32'h3f148a53, 32'hc0c74b76} /* (4, 11, 29) {real, imag} */,
  {32'h3f81bfb6, 32'hc0923f32} /* (4, 11, 28) {real, imag} */,
  {32'h3efbb496, 32'hc0567b8a} /* (4, 11, 27) {real, imag} */,
  {32'h3fec483d, 32'hc02430fe} /* (4, 11, 26) {real, imag} */,
  {32'h3fdcf1ff, 32'hc06934c8} /* (4, 11, 25) {real, imag} */,
  {32'h407612c1, 32'hc03bbe8e} /* (4, 11, 24) {real, imag} */,
  {32'h402a2504, 32'hc099a0c0} /* (4, 11, 23) {real, imag} */,
  {32'h3f83c14b, 32'hc0839d42} /* (4, 11, 22) {real, imag} */,
  {32'h401fdf5e, 32'hc0a073b9} /* (4, 11, 21) {real, imag} */,
  {32'h3eeb1def, 32'h3f353671} /* (4, 11, 20) {real, imag} */,
  {32'hc01c48b0, 32'h40820673} /* (4, 11, 19) {real, imag} */,
  {32'hc0637e7a, 32'h409b8a28} /* (4, 11, 18) {real, imag} */,
  {32'hc08853f8, 32'h40caf940} /* (4, 11, 17) {real, imag} */,
  {32'hc07274f0, 32'h409885b6} /* (4, 11, 16) {real, imag} */,
  {32'hc017aa97, 32'h4026fa15} /* (4, 11, 15) {real, imag} */,
  {32'hbecc037e, 32'h409cffcc} /* (4, 11, 14) {real, imag} */,
  {32'hbf133b60, 32'h4094955f} /* (4, 11, 13) {real, imag} */,
  {32'hbfa8c687, 32'h409c878e} /* (4, 11, 12) {real, imag} */,
  {32'hc007f51f, 32'h40a7f78a} /* (4, 11, 11) {real, imag} */,
  {32'hc03abdc8, 32'hbfc482d9} /* (4, 11, 10) {real, imag} */,
  {32'h3fc2fc36, 32'hc0ec2e51} /* (4, 11, 9) {real, imag} */,
  {32'h40662ca4, 32'hc0babfd8} /* (4, 11, 8) {real, imag} */,
  {32'h409a633d, 32'hc0b039ac} /* (4, 11, 7) {real, imag} */,
  {32'h40c36b7e, 32'hc0de74fe} /* (4, 11, 6) {real, imag} */,
  {32'h40808802, 32'hc0c13ad0} /* (4, 11, 5) {real, imag} */,
  {32'h402cf1a6, 32'hc0729936} /* (4, 11, 4) {real, imag} */,
  {32'h4045b3fa, 32'hc06a92d1} /* (4, 11, 3) {real, imag} */,
  {32'h404af6e1, 32'hc04cf7ae} /* (4, 11, 2) {real, imag} */,
  {32'h3f59df00, 32'hc081e1bb} /* (4, 11, 1) {real, imag} */,
  {32'h3fd0cca4, 32'hc04b0e41} /* (4, 11, 0) {real, imag} */,
  {32'hbfd253cc, 32'h406992a8} /* (4, 10, 31) {real, imag} */,
  {32'hc04026b5, 32'h4045ec32} /* (4, 10, 30) {real, imag} */,
  {32'hbfe14e06, 32'h3ff80f44} /* (4, 10, 29) {real, imag} */,
  {32'hbfb4734c, 32'h4074382c} /* (4, 10, 28) {real, imag} */,
  {32'hc02759be, 32'h407a4fd4} /* (4, 10, 27) {real, imag} */,
  {32'hbf9d2de9, 32'h40955d22} /* (4, 10, 26) {real, imag} */,
  {32'hbf7904e5, 32'h408691b8} /* (4, 10, 25) {real, imag} */,
  {32'hbe2c4758, 32'h40770484} /* (4, 10, 24) {real, imag} */,
  {32'h3d90c036, 32'h3ea3a29c} /* (4, 10, 23) {real, imag} */,
  {32'hbf19fdb9, 32'h3f1d72f6} /* (4, 10, 22) {real, imag} */,
  {32'h3ee3877b, 32'hc069a158} /* (4, 10, 21) {real, imag} */,
  {32'h403d49c2, 32'hc08a062a} /* (4, 10, 20) {real, imag} */,
  {32'h3fb0712a, 32'hbf0598b2} /* (4, 10, 19) {real, imag} */,
  {32'h400b8880, 32'hbe082ea0} /* (4, 10, 18) {real, imag} */,
  {32'h401893b4, 32'hbfab98a1} /* (4, 10, 17) {real, imag} */,
  {32'hbf988c53, 32'hc01d228d} /* (4, 10, 16) {real, imag} */,
  {32'hbff8a099, 32'hc0941a4e} /* (4, 10, 15) {real, imag} */,
  {32'hbe2e9128, 32'hbff0b422} /* (4, 10, 14) {real, imag} */,
  {32'h3f5cb248, 32'hc01483c2} /* (4, 10, 13) {real, imag} */,
  {32'h3fa8b28d, 32'hc020caeb} /* (4, 10, 12) {real, imag} */,
  {32'h3ef2911e, 32'hbfc0ba04} /* (4, 10, 11) {real, imag} */,
  {32'hbf5ab3e8, 32'hbf3662bb} /* (4, 10, 10) {real, imag} */,
  {32'h3fa55964, 32'hbe3d2630} /* (4, 10, 9) {real, imag} */,
  {32'h3f8725a7, 32'h4025d318} /* (4, 10, 8) {real, imag} */,
  {32'h3e439e80, 32'h3f0c95db} /* (4, 10, 7) {real, imag} */,
  {32'h3fcde138, 32'hc0009fea} /* (4, 10, 6) {real, imag} */,
  {32'h3ec1486e, 32'h3e5b1e45} /* (4, 10, 5) {real, imag} */,
  {32'hbda8b564, 32'h3f73a9bd} /* (4, 10, 4) {real, imag} */,
  {32'h3ea090f6, 32'h405a4f4d} /* (4, 10, 3) {real, imag} */,
  {32'h3e132a39, 32'h40ba6621} /* (4, 10, 2) {real, imag} */,
  {32'hc05b5ac2, 32'h40a87b95} /* (4, 10, 1) {real, imag} */,
  {32'hbf95c5ec, 32'h4065f720} /* (4, 10, 0) {real, imag} */,
  {32'hc01f841f, 32'h4080deb8} /* (4, 9, 31) {real, imag} */,
  {32'hc04ebc12, 32'h40c3880a} /* (4, 9, 30) {real, imag} */,
  {32'hc02a7d45, 32'h40098cb3} /* (4, 9, 29) {real, imag} */,
  {32'hc01f90c4, 32'h408f29c2} /* (4, 9, 28) {real, imag} */,
  {32'hc076f58c, 32'h40c5ebe3} /* (4, 9, 27) {real, imag} */,
  {32'hc02d0d02, 32'h40f6e8fe} /* (4, 9, 26) {real, imag} */,
  {32'hc014d262, 32'h40dbc6d2} /* (4, 9, 25) {real, imag} */,
  {32'hc03b90bc, 32'h40b5f12e} /* (4, 9, 24) {real, imag} */,
  {32'hbfae09ab, 32'h4083a901} /* (4, 9, 23) {real, imag} */,
  {32'hbff19077, 32'h40d84cc0} /* (4, 9, 22) {real, imag} */,
  {32'hbf28c779, 32'h40221f25} /* (4, 9, 21) {real, imag} */,
  {32'h3fb8f130, 32'hc095211b} /* (4, 9, 20) {real, imag} */,
  {32'h3ff5bcd3, 32'hc06a4895} /* (4, 9, 19) {real, imag} */,
  {32'h3f00cfe6, 32'hc0710180} /* (4, 9, 18) {real, imag} */,
  {32'h401ec09f, 32'hc0bd3bdd} /* (4, 9, 17) {real, imag} */,
  {32'h4029a758, 32'hc0939c66} /* (4, 9, 16) {real, imag} */,
  {32'h3e82f99e, 32'hc0c5868e} /* (4, 9, 15) {real, imag} */,
  {32'h401e9476, 32'hc0cfcd12} /* (4, 9, 14) {real, imag} */,
  {32'h3f828f39, 32'hc0378679} /* (4, 9, 13) {real, imag} */,
  {32'h3fd47c1e, 32'hc088db5c} /* (4, 9, 12) {real, imag} */,
  {32'h3f95e725, 32'hc080c478} /* (4, 9, 11) {real, imag} */,
  {32'hc023cf39, 32'h3f75e2aa} /* (4, 9, 10) {real, imag} */,
  {32'hbf954d6d, 32'h403cc59d} /* (4, 9, 9) {real, imag} */,
  {32'hbfa38906, 32'h4049caeb} /* (4, 9, 8) {real, imag} */,
  {32'hc0218fa6, 32'h405f1c5c} /* (4, 9, 7) {real, imag} */,
  {32'h3f524a0b, 32'h3ffad769} /* (4, 9, 6) {real, imag} */,
  {32'hbfc2095c, 32'h40ce8d55} /* (4, 9, 5) {real, imag} */,
  {32'hbee025fc, 32'h40d4fb5c} /* (4, 9, 4) {real, imag} */,
  {32'hbf936917, 32'h40d6a489} /* (4, 9, 3) {real, imag} */,
  {32'hbf846d03, 32'h41058f28} /* (4, 9, 2) {real, imag} */,
  {32'hc018e616, 32'h410219df} /* (4, 9, 1) {real, imag} */,
  {32'hbfce068f, 32'h40aa5884} /* (4, 9, 0) {real, imag} */,
  {32'hbfc050c5, 32'h4093f578} /* (4, 8, 31) {real, imag} */,
  {32'hbefac69c, 32'h40d503da} /* (4, 8, 30) {real, imag} */,
  {32'hbf2b1128, 32'h403cad75} /* (4, 8, 29) {real, imag} */,
  {32'hbeebb18e, 32'h4057cc29} /* (4, 8, 28) {real, imag} */,
  {32'hbf5f271f, 32'h40387652} /* (4, 8, 27) {real, imag} */,
  {32'hbf0897c2, 32'h409369aa} /* (4, 8, 26) {real, imag} */,
  {32'hbf5603fe, 32'h4062e252} /* (4, 8, 25) {real, imag} */,
  {32'hc02c75e6, 32'h40757320} /* (4, 8, 24) {real, imag} */,
  {32'hc0099894, 32'h4075a6d7} /* (4, 8, 23) {real, imag} */,
  {32'hbf9acfa2, 32'h409db6fa} /* (4, 8, 22) {real, imag} */,
  {32'hbf933457, 32'h4009fb9b} /* (4, 8, 21) {real, imag} */,
  {32'hbf9f3d6e, 32'hc08b1fc2} /* (4, 8, 20) {real, imag} */,
  {32'hbd0f901a, 32'hc0a84f4c} /* (4, 8, 19) {real, imag} */,
  {32'hbf6a76d7, 32'hc046af56} /* (4, 8, 18) {real, imag} */,
  {32'h3f890413, 32'hc03e98d8} /* (4, 8, 17) {real, imag} */,
  {32'h40931506, 32'hc0891a27} /* (4, 8, 16) {real, imag} */,
  {32'h3f99eb77, 32'hc0750af2} /* (4, 8, 15) {real, imag} */,
  {32'h4036d118, 32'hc0c9129a} /* (4, 8, 14) {real, imag} */,
  {32'h405a77e2, 32'hc092548b} /* (4, 8, 13) {real, imag} */,
  {32'h4025f046, 32'hc0949d3c} /* (4, 8, 12) {real, imag} */,
  {32'h3fb0d1a9, 32'hbfee243a} /* (4, 8, 11) {real, imag} */,
  {32'h3c366ac0, 32'h408b06d5} /* (4, 8, 10) {real, imag} */,
  {32'h3d8397f4, 32'h4084a422} /* (4, 8, 9) {real, imag} */,
  {32'hbf7a1625, 32'h3ffc3934} /* (4, 8, 8) {real, imag} */,
  {32'hc01beeeb, 32'h4033599e} /* (4, 8, 7) {real, imag} */,
  {32'h3f15e495, 32'h4056fb1e} /* (4, 8, 6) {real, imag} */,
  {32'hc016f64a, 32'h409a4960} /* (4, 8, 5) {real, imag} */,
  {32'hbeed48ca, 32'h409ac014} /* (4, 8, 4) {real, imag} */,
  {32'hbe73f4d4, 32'h40ea9d78} /* (4, 8, 3) {real, imag} */,
  {32'hc07f31c2, 32'h40f148be} /* (4, 8, 2) {real, imag} */,
  {32'hc08467eb, 32'h40d35e12} /* (4, 8, 1) {real, imag} */,
  {32'hbffb33aa, 32'h40aff3f1} /* (4, 8, 0) {real, imag} */,
  {32'hbf4ae59c, 32'h4094e537} /* (4, 7, 31) {real, imag} */,
  {32'hbf46e7d8, 32'h40c72c3f} /* (4, 7, 30) {real, imag} */,
  {32'h3ff9704c, 32'h409d198c} /* (4, 7, 29) {real, imag} */,
  {32'hbd191c60, 32'h40a002bb} /* (4, 7, 28) {real, imag} */,
  {32'hbfcb51f0, 32'h404040dd} /* (4, 7, 27) {real, imag} */,
  {32'hbfdb155d, 32'h4080a250} /* (4, 7, 26) {real, imag} */,
  {32'hc00384eb, 32'h406d93c4} /* (4, 7, 25) {real, imag} */,
  {32'hbfb374b9, 32'h40b98f68} /* (4, 7, 24) {real, imag} */,
  {32'hc06e0fc4, 32'h40965484} /* (4, 7, 23) {real, imag} */,
  {32'hbfe98c6c, 32'h40a130b3} /* (4, 7, 22) {real, imag} */,
  {32'hbf36e7c8, 32'h3fcfad43} /* (4, 7, 21) {real, imag} */,
  {32'h3f9287e6, 32'hc0d785f3} /* (4, 7, 20) {real, imag} */,
  {32'h3f6ffb62, 32'hc0ac7c92} /* (4, 7, 19) {real, imag} */,
  {32'hbe8ebc52, 32'hc082749b} /* (4, 7, 18) {real, imag} */,
  {32'h3e1ea2f6, 32'hc0815a46} /* (4, 7, 17) {real, imag} */,
  {32'h3db56784, 32'hc067816c} /* (4, 7, 16) {real, imag} */,
  {32'hbf73e91e, 32'hc0b4050b} /* (4, 7, 15) {real, imag} */,
  {32'h3fd0e542, 32'hc0e0a67c} /* (4, 7, 14) {real, imag} */,
  {32'h405c7f26, 32'hc09a5a86} /* (4, 7, 13) {real, imag} */,
  {32'h3fb56270, 32'hc0940c91} /* (4, 7, 12) {real, imag} */,
  {32'h3f081141, 32'hbff8ffa7} /* (4, 7, 11) {real, imag} */,
  {32'h3f0c664d, 32'h40b17481} /* (4, 7, 10) {real, imag} */,
  {32'hbfe2cd8e, 32'h40d3416b} /* (4, 7, 9) {real, imag} */,
  {32'hbfb3e6cc, 32'h40b3a5f5} /* (4, 7, 8) {real, imag} */,
  {32'hbf92179c, 32'h408df42a} /* (4, 7, 7) {real, imag} */,
  {32'hbfe9332b, 32'h407e273a} /* (4, 7, 6) {real, imag} */,
  {32'hc01fc5a6, 32'h409f9fd6} /* (4, 7, 5) {real, imag} */,
  {32'hc02ae63a, 32'h409bc6ec} /* (4, 7, 4) {real, imag} */,
  {32'hbfc4d5c6, 32'h40bc0c6a} /* (4, 7, 3) {real, imag} */,
  {32'hc0c2a92a, 32'h40e2916a} /* (4, 7, 2) {real, imag} */,
  {32'hc08f1fb6, 32'h40b807f0} /* (4, 7, 1) {real, imag} */,
  {32'h3d81c520, 32'h4041c7f0} /* (4, 7, 0) {real, imag} */,
  {32'hbf2f1181, 32'h403ece16} /* (4, 6, 31) {real, imag} */,
  {32'hbfb6f213, 32'h40e8d8c8} /* (4, 6, 30) {real, imag} */,
  {32'hbe5ceb64, 32'h40be8afd} /* (4, 6, 29) {real, imag} */,
  {32'hbfd3d302, 32'h404c4732} /* (4, 6, 28) {real, imag} */,
  {32'hc00bfd08, 32'h40218c98} /* (4, 6, 27) {real, imag} */,
  {32'hc06d842a, 32'h40634524} /* (4, 6, 26) {real, imag} */,
  {32'hc08b096c, 32'h40b890f4} /* (4, 6, 25) {real, imag} */,
  {32'hbfde7c87, 32'h40e434a0} /* (4, 6, 24) {real, imag} */,
  {32'hc0538da0, 32'h4085250b} /* (4, 6, 23) {real, imag} */,
  {32'hc0881583, 32'h40a0349a} /* (4, 6, 22) {real, imag} */,
  {32'hc088575f, 32'h401829b4} /* (4, 6, 21) {real, imag} */,
  {32'h400108b4, 32'hc0cd7fe8} /* (4, 6, 20) {real, imag} */,
  {32'h3fc036b5, 32'hc09cf15e} /* (4, 6, 19) {real, imag} */,
  {32'h3ffcea60, 32'hc046759a} /* (4, 6, 18) {real, imag} */,
  {32'h3f6db947, 32'hc0c2b57c} /* (4, 6, 17) {real, imag} */,
  {32'h3f802ece, 32'hc0845a54} /* (4, 6, 16) {real, imag} */,
  {32'h3d8317d4, 32'hc098047e} /* (4, 6, 15) {real, imag} */,
  {32'h3f238b2c, 32'hc09784eb} /* (4, 6, 14) {real, imag} */,
  {32'h4015b0b0, 32'hbfe5e003} /* (4, 6, 13) {real, imag} */,
  {32'h3ff6f9d6, 32'hc0a64b95} /* (4, 6, 12) {real, imag} */,
  {32'h3fe5194b, 32'hc077e18f} /* (4, 6, 11) {real, imag} */,
  {32'hbf304632, 32'h3fc073e8} /* (4, 6, 10) {real, imag} */,
  {32'hc0934811, 32'h40a9f355} /* (4, 6, 9) {real, imag} */,
  {32'hc03c965b, 32'h409b61de} /* (4, 6, 8) {real, imag} */,
  {32'hc0391d0d, 32'h405b098d} /* (4, 6, 7) {real, imag} */,
  {32'hbf472c43, 32'h40a718d2} /* (4, 6, 6) {real, imag} */,
  {32'hbf21b40f, 32'h40d09c47} /* (4, 6, 5) {real, imag} */,
  {32'hc059ba83, 32'h40db4b56} /* (4, 6, 4) {real, imag} */,
  {32'hbfe31331, 32'h40ab9bf2} /* (4, 6, 3) {real, imag} */,
  {32'hbfdd3520, 32'h40dec746} /* (4, 6, 2) {real, imag} */,
  {32'hc012af6c, 32'h40999654} /* (4, 6, 1) {real, imag} */,
  {32'hbf311dbc, 32'h3f1e1072} /* (4, 6, 0) {real, imag} */,
  {32'hbfee2cb9, 32'h40ac44b8} /* (4, 5, 31) {real, imag} */,
  {32'hc093431a, 32'h40c3729c} /* (4, 5, 30) {real, imag} */,
  {32'hc06f1dfc, 32'h40b988e0} /* (4, 5, 29) {real, imag} */,
  {32'hc02d6b6f, 32'h40a7d448} /* (4, 5, 28) {real, imag} */,
  {32'hbfe6404c, 32'h40155981} /* (4, 5, 27) {real, imag} */,
  {32'hbfcea652, 32'h3fb8affa} /* (4, 5, 26) {real, imag} */,
  {32'hc0093ded, 32'h4062bb9e} /* (4, 5, 25) {real, imag} */,
  {32'hbe4d4134, 32'h40c8a45e} /* (4, 5, 24) {real, imag} */,
  {32'hc0189aaf, 32'h40a11d3f} /* (4, 5, 23) {real, imag} */,
  {32'hc07e2ed7, 32'h40983ddc} /* (4, 5, 22) {real, imag} */,
  {32'hc0c693ec, 32'h40132f6f} /* (4, 5, 21) {real, imag} */,
  {32'hbfb5f994, 32'hbf8ccbc9} /* (4, 5, 20) {real, imag} */,
  {32'hbf511a96, 32'hbe8a4b47} /* (4, 5, 19) {real, imag} */,
  {32'hc0085c8c, 32'h3f953a78} /* (4, 5, 18) {real, imag} */,
  {32'hc017029c, 32'hbf93e58f} /* (4, 5, 17) {real, imag} */,
  {32'hbfa76626, 32'hbe4a7d5b} /* (4, 5, 16) {real, imag} */,
  {32'h3e88a274, 32'hc0340a48} /* (4, 5, 15) {real, imag} */,
  {32'h3ece4391, 32'hc0248f94} /* (4, 5, 14) {real, imag} */,
  {32'h3f4ba5ea, 32'hc040d5ea} /* (4, 5, 13) {real, imag} */,
  {32'hbf48846b, 32'hc0b86a6e} /* (4, 5, 12) {real, imag} */,
  {32'h3fcbd78d, 32'hc0a5689c} /* (4, 5, 11) {real, imag} */,
  {32'hbe8bceb8, 32'hc0973b0e} /* (4, 5, 10) {real, imag} */,
  {32'hbe8ee5c5, 32'hc0545a52} /* (4, 5, 9) {real, imag} */,
  {32'hbefbe734, 32'hc0457438} /* (4, 5, 8) {real, imag} */,
  {32'hbf98ba52, 32'hbfdfa18e} /* (4, 5, 7) {real, imag} */,
  {32'hbce5cd20, 32'h4011c794} /* (4, 5, 6) {real, imag} */,
  {32'hbf6870a7, 32'h4097d7fa} /* (4, 5, 5) {real, imag} */,
  {32'hbfcb260f, 32'h410affe6} /* (4, 5, 4) {real, imag} */,
  {32'hc055e617, 32'h40946546} /* (4, 5, 3) {real, imag} */,
  {32'hc0574e8c, 32'h40935e27} /* (4, 5, 2) {real, imag} */,
  {32'hbfe896b8, 32'h40786222} /* (4, 5, 1) {real, imag} */,
  {32'hbf75e182, 32'h3fb3a299} /* (4, 5, 0) {real, imag} */,
  {32'hbf8575bd, 32'h4090793c} /* (4, 4, 31) {real, imag} */,
  {32'hc08e548e, 32'h40ac5ad0} /* (4, 4, 30) {real, imag} */,
  {32'hc085cdd2, 32'h40afae46} /* (4, 4, 29) {real, imag} */,
  {32'hbf9d1158, 32'h40a47174} /* (4, 4, 28) {real, imag} */,
  {32'h3f1acf57, 32'h40906be8} /* (4, 4, 27) {real, imag} */,
  {32'h3f429b82, 32'h404724bc} /* (4, 4, 26) {real, imag} */,
  {32'hbf5fcdd4, 32'h400877f3} /* (4, 4, 25) {real, imag} */,
  {32'h3f98c703, 32'h4085f451} /* (4, 4, 24) {real, imag} */,
  {32'hbf6d1495, 32'h40be2ca0} /* (4, 4, 23) {real, imag} */,
  {32'hc02ff7e0, 32'h40ac022a} /* (4, 4, 22) {real, imag} */,
  {32'hc08f6ac5, 32'h40b1144c} /* (4, 4, 21) {real, imag} */,
  {32'hc0b89366, 32'h40a29934} /* (4, 4, 20) {real, imag} */,
  {32'hc033b29c, 32'h4085235f} /* (4, 4, 19) {real, imag} */,
  {32'hc05dec88, 32'h40a1fbca} /* (4, 4, 18) {real, imag} */,
  {32'hc0be9192, 32'h4099f629} /* (4, 4, 17) {real, imag} */,
  {32'hc0a83a98, 32'h400a9385} /* (4, 4, 16) {real, imag} */,
  {32'h3ec0b611, 32'hc09c2768} /* (4, 4, 15) {real, imag} */,
  {32'h3ff7004b, 32'hc0a07a92} /* (4, 4, 14) {real, imag} */,
  {32'h3e1d5a7e, 32'hc061803f} /* (4, 4, 13) {real, imag} */,
  {32'hbfccd680, 32'hc09db210} /* (4, 4, 12) {real, imag} */,
  {32'h3e9c54ce, 32'hc0db5718} /* (4, 4, 11) {real, imag} */,
  {32'h400450cc, 32'hc1004f7c} /* (4, 4, 10) {real, imag} */,
  {32'h403bfe3c, 32'hc0f0a5f1} /* (4, 4, 9) {real, imag} */,
  {32'h402bf483, 32'hc0e6fefa} /* (4, 4, 8) {real, imag} */,
  {32'h4000bc2e, 32'hc0b2ab3c} /* (4, 4, 7) {real, imag} */,
  {32'h3f57a28e, 32'hc03a296a} /* (4, 4, 6) {real, imag} */,
  {32'hbfe992d2, 32'hbe230d44} /* (4, 4, 5) {real, imag} */,
  {32'hc0679d2e, 32'h409bb19e} /* (4, 4, 4) {real, imag} */,
  {32'hbfbf6c12, 32'h4072e4c2} /* (4, 4, 3) {real, imag} */,
  {32'hc0371a3e, 32'h4016929a} /* (4, 4, 2) {real, imag} */,
  {32'hbeb3de0e, 32'h40924226} /* (4, 4, 1) {real, imag} */,
  {32'h3ea11006, 32'h4018b3ec} /* (4, 4, 0) {real, imag} */,
  {32'hbe69b537, 32'h404b7258} /* (4, 3, 31) {real, imag} */,
  {32'hc034eaa8, 32'h40717a28} /* (4, 3, 30) {real, imag} */,
  {32'hc0813f5f, 32'h4050fcd2} /* (4, 3, 29) {real, imag} */,
  {32'hc084aaee, 32'h3fe95426} /* (4, 3, 28) {real, imag} */,
  {32'hc06dc496, 32'h40ae48f1} /* (4, 3, 27) {real, imag} */,
  {32'hbee55cd8, 32'h40b61a6c} /* (4, 3, 26) {real, imag} */,
  {32'hbf542c2d, 32'h4081c89e} /* (4, 3, 25) {real, imag} */,
  {32'hbe25fee7, 32'h40addac8} /* (4, 3, 24) {real, imag} */,
  {32'hbee55a2b, 32'h409ca7df} /* (4, 3, 23) {real, imag} */,
  {32'hc0077fb6, 32'h40d6f37c} /* (4, 3, 22) {real, imag} */,
  {32'hbfecaef2, 32'h40a282f0} /* (4, 3, 21) {real, imag} */,
  {32'hc01ff259, 32'h4096ccd2} /* (4, 3, 20) {real, imag} */,
  {32'hbf5f8408, 32'h409c9f6a} /* (4, 3, 19) {real, imag} */,
  {32'hc07b46b7, 32'h40ba6a2e} /* (4, 3, 18) {real, imag} */,
  {32'hc081f5d4, 32'h40993e5a} /* (4, 3, 17) {real, imag} */,
  {32'hc0132f04, 32'h4007f1e8} /* (4, 3, 16) {real, imag} */,
  {32'h3fa4a7d6, 32'hc047cb5c} /* (4, 3, 15) {real, imag} */,
  {32'h4030309c, 32'hc0a976f3} /* (4, 3, 14) {real, imag} */,
  {32'h4023165f, 32'hc0aac019} /* (4, 3, 13) {real, imag} */,
  {32'h3f3fa6bc, 32'hc0e77eb3} /* (4, 3, 12) {real, imag} */,
  {32'h4042a3de, 32'hc0ff9648} /* (4, 3, 11) {real, imag} */,
  {32'h405a5c58, 32'hc0d2ba78} /* (4, 3, 10) {real, imag} */,
  {32'h3fdb0d44, 32'hc0cb6684} /* (4, 3, 9) {real, imag} */,
  {32'h3fdaa7b0, 32'hc0c0215e} /* (4, 3, 8) {real, imag} */,
  {32'hbfe32990, 32'hc0affb44} /* (4, 3, 7) {real, imag} */,
  {32'h3f10b5a2, 32'hc081226f} /* (4, 3, 6) {real, imag} */,
  {32'hbf8055ee, 32'h3f61e053} /* (4, 3, 5) {real, imag} */,
  {32'hc06f9419, 32'h40a36c6f} /* (4, 3, 4) {real, imag} */,
  {32'h4018015c, 32'h407777aa} /* (4, 3, 3) {real, imag} */,
  {32'hbe32d42a, 32'hbec3974c} /* (4, 3, 2) {real, imag} */,
  {32'h3fd01547, 32'h3ffbb3c0} /* (4, 3, 1) {real, imag} */,
  {32'hbec1d89d, 32'h3ff7c3d2} /* (4, 3, 0) {real, imag} */,
  {32'hbf816a42, 32'h403330d7} /* (4, 2, 31) {real, imag} */,
  {32'hbfb79e36, 32'h40c3a1f4} /* (4, 2, 30) {real, imag} */,
  {32'hc0146bf6, 32'h407a6ca6} /* (4, 2, 29) {real, imag} */,
  {32'hc066f9a6, 32'h40833f3a} /* (4, 2, 28) {real, imag} */,
  {32'hc062084c, 32'h40ab7326} /* (4, 2, 27) {real, imag} */,
  {32'hc022f3aa, 32'h40a73f12} /* (4, 2, 26) {real, imag} */,
  {32'hc014bbdf, 32'h406c047a} /* (4, 2, 25) {real, imag} */,
  {32'hc0211f55, 32'h4042ffc8} /* (4, 2, 24) {real, imag} */,
  {32'hbf1ffb40, 32'h4018a3ae} /* (4, 2, 23) {real, imag} */,
  {32'hbfe2c754, 32'h40b0f66e} /* (4, 2, 22) {real, imag} */,
  {32'hbff9eb4b, 32'h409ce697} /* (4, 2, 21) {real, imag} */,
  {32'hbf8d40a5, 32'h4093ada9} /* (4, 2, 20) {real, imag} */,
  {32'hbfb7b439, 32'h40a0b937} /* (4, 2, 19) {real, imag} */,
  {32'hc09627f8, 32'h40fd3d5e} /* (4, 2, 18) {real, imag} */,
  {32'hc04cac32, 32'h40aa0a7f} /* (4, 2, 17) {real, imag} */,
  {32'hbfa4a6f6, 32'h3fc38de4} /* (4, 2, 16) {real, imag} */,
  {32'h3f96d335, 32'hc04e902a} /* (4, 2, 15) {real, imag} */,
  {32'h4061350d, 32'hc04a0ca2} /* (4, 2, 14) {real, imag} */,
  {32'h40b728fc, 32'hc09edadb} /* (4, 2, 13) {real, imag} */,
  {32'h4046cfe2, 32'hc0ae9708} /* (4, 2, 12) {real, imag} */,
  {32'h4070458a, 32'hc0bc8e14} /* (4, 2, 11) {real, imag} */,
  {32'h4093a0fe, 32'hc0b00e82} /* (4, 2, 10) {real, imag} */,
  {32'h403b4ce8, 32'hc0bed87e} /* (4, 2, 9) {real, imag} */,
  {32'h400e5b6b, 32'hc06a7a67} /* (4, 2, 8) {real, imag} */,
  {32'hbf0f33a2, 32'hc0b18e08} /* (4, 2, 7) {real, imag} */,
  {32'h3faf2393, 32'hc08e5d1c} /* (4, 2, 6) {real, imag} */,
  {32'h3ed6ef1c, 32'h402822f5} /* (4, 2, 5) {real, imag} */,
  {32'hc02374a1, 32'h40d22542} /* (4, 2, 4) {real, imag} */,
  {32'h3f3f7885, 32'h40c7602b} /* (4, 2, 3) {real, imag} */,
  {32'hbe4ef712, 32'h4022d2d4} /* (4, 2, 2) {real, imag} */,
  {32'hbcb96ef8, 32'h404586b4} /* (4, 2, 1) {real, imag} */,
  {32'hbfab4f36, 32'h40091a4e} /* (4, 2, 0) {real, imag} */,
  {32'hc0057caf, 32'h3ffcc127} /* (4, 1, 31) {real, imag} */,
  {32'hc025cfda, 32'h4078d922} /* (4, 1, 30) {real, imag} */,
  {32'hbfc3ae48, 32'h40390198} /* (4, 1, 29) {real, imag} */,
  {32'hbfad28b8, 32'h407158ae} /* (4, 1, 28) {real, imag} */,
  {32'hbfbbca7b, 32'h3fff0e14} /* (4, 1, 27) {real, imag} */,
  {32'hbfc36b72, 32'h3fc7ea62} /* (4, 1, 26) {real, imag} */,
  {32'hbf0a45f0, 32'h40198c48} /* (4, 1, 25) {real, imag} */,
  {32'hbfd61b0a, 32'h3ff5951b} /* (4, 1, 24) {real, imag} */,
  {32'hc013c9c1, 32'h4002fccf} /* (4, 1, 23) {real, imag} */,
  {32'hc03a2e55, 32'h405f97b7} /* (4, 1, 22) {real, imag} */,
  {32'hc00b724c, 32'h409903d4} /* (4, 1, 21) {real, imag} */,
  {32'hbf9602dc, 32'h4059f9fa} /* (4, 1, 20) {real, imag} */,
  {32'hc0633efe, 32'h406f0a98} /* (4, 1, 19) {real, imag} */,
  {32'hc09b0667, 32'h40c0d0f9} /* (4, 1, 18) {real, imag} */,
  {32'hc0441ec2, 32'h408eba62} /* (4, 1, 17) {real, imag} */,
  {32'hc05d8ca6, 32'h3f9648b1} /* (4, 1, 16) {real, imag} */,
  {32'h3fa2c447, 32'hc00dfb39} /* (4, 1, 15) {real, imag} */,
  {32'h4087bf1a, 32'hbfd8aa9c} /* (4, 1, 14) {real, imag} */,
  {32'h40a31a76, 32'hc03801c6} /* (4, 1, 13) {real, imag} */,
  {32'h4094b97a, 32'hc07278a6} /* (4, 1, 12) {real, imag} */,
  {32'h40325418, 32'hc0d97ff9} /* (4, 1, 11) {real, imag} */,
  {32'h3f337f6a, 32'hc0c36918} /* (4, 1, 10) {real, imag} */,
  {32'h3ee010b7, 32'hc098c4a5} /* (4, 1, 9) {real, imag} */,
  {32'h406410ae, 32'hc0734d26} /* (4, 1, 8) {real, imag} */,
  {32'h400bcd64, 32'hc08fc52c} /* (4, 1, 7) {real, imag} */,
  {32'hbe37ae58, 32'hc0a334a4} /* (4, 1, 6) {real, imag} */,
  {32'hc002db93, 32'h3de5a610} /* (4, 1, 5) {real, imag} */,
  {32'hbfcac572, 32'h4091921d} /* (4, 1, 4) {real, imag} */,
  {32'h3e9d205f, 32'h40aa292d} /* (4, 1, 3) {real, imag} */,
  {32'hbf7d133e, 32'h4080ce41} /* (4, 1, 2) {real, imag} */,
  {32'hbfc0aaa5, 32'h4057c38c} /* (4, 1, 1) {real, imag} */,
  {32'hbfff3f60, 32'h3f9820c2} /* (4, 1, 0) {real, imag} */,
  {32'hbf2022f7, 32'h4016a72e} /* (4, 0, 31) {real, imag} */,
  {32'hc00aa408, 32'h3fd4c7f4} /* (4, 0, 30) {real, imag} */,
  {32'hc006bc70, 32'h3fbff62e} /* (4, 0, 29) {real, imag} */,
  {32'hbf9fda7d, 32'h400eb574} /* (4, 0, 28) {real, imag} */,
  {32'hbfdc0bbc, 32'h3f93220c} /* (4, 0, 27) {real, imag} */,
  {32'hbfa5d875, 32'h3ebf8ca9} /* (4, 0, 26) {real, imag} */,
  {32'h3e941138, 32'h3fbfddb2} /* (4, 0, 25) {real, imag} */,
  {32'hbfaa8dcc, 32'h3f95e9bf} /* (4, 0, 24) {real, imag} */,
  {32'hc04339e4, 32'h4018f072} /* (4, 0, 23) {real, imag} */,
  {32'hc0437bb4, 32'h402bdb96} /* (4, 0, 22) {real, imag} */,
  {32'hc00b4ae0, 32'h40752c79} /* (4, 0, 21) {real, imag} */,
  {32'hbfcfcb12, 32'h4003fce7} /* (4, 0, 20) {real, imag} */,
  {32'hc03729c4, 32'h3f94a770} /* (4, 0, 19) {real, imag} */,
  {32'hc01d8a8c, 32'h3fd0cade} /* (4, 0, 18) {real, imag} */,
  {32'hbf1ae02d, 32'h3fc718f6} /* (4, 0, 17) {real, imag} */,
  {32'hbf85f9a8, 32'h3ec6649a} /* (4, 0, 16) {real, imag} */,
  {32'h3f33aafe, 32'hbfd36aee} /* (4, 0, 15) {real, imag} */,
  {32'h3faab354, 32'hc02dc358} /* (4, 0, 14) {real, imag} */,
  {32'hbeeef802, 32'hc055550c} /* (4, 0, 13) {real, imag} */,
  {32'h3f458595, 32'hc03d2462} /* (4, 0, 12) {real, imag} */,
  {32'h3f5c8b1e, 32'hc0741187} /* (4, 0, 11) {real, imag} */,
  {32'hbf83d288, 32'hc064803e} /* (4, 0, 10) {real, imag} */,
  {32'hc025a006, 32'hc02951b5} /* (4, 0, 9) {real, imag} */,
  {32'h3f51d1f0, 32'hc01aa48c} /* (4, 0, 8) {real, imag} */,
  {32'h3fc180dc, 32'hc04eb7cd} /* (4, 0, 7) {real, imag} */,
  {32'h3f9a3c56, 32'hc077031a} /* (4, 0, 6) {real, imag} */,
  {32'hbf327cfe, 32'h3d379986} /* (4, 0, 5) {real, imag} */,
  {32'hbf46a603, 32'h3fed28e4} /* (4, 0, 4) {real, imag} */,
  {32'hbee01b5e, 32'h407553cf} /* (4, 0, 3) {real, imag} */,
  {32'hbfea9794, 32'h4070801a} /* (4, 0, 2) {real, imag} */,
  {32'hbeed8c88, 32'h400f4184} /* (4, 0, 1) {real, imag} */,
  {32'hbd127990, 32'h3f25bdbc} /* (4, 0, 0) {real, imag} */,
  {32'hbf23fc40, 32'hbe9e3f56} /* (3, 31, 31) {real, imag} */,
  {32'hbf986902, 32'hbd7bed00} /* (3, 31, 30) {real, imag} */,
  {32'hbf9489ba, 32'h4023d0f0} /* (3, 31, 29) {real, imag} */,
  {32'hc03c8b61, 32'h405b652e} /* (3, 31, 28) {real, imag} */,
  {32'hbfe7cba2, 32'h40703c0d} /* (3, 31, 27) {real, imag} */,
  {32'hbf74ef53, 32'h3ffd8d3b} /* (3, 31, 26) {real, imag} */,
  {32'hbf38be58, 32'h4083a241} /* (3, 31, 25) {real, imag} */,
  {32'h3ef0fc4a, 32'h408e397a} /* (3, 31, 24) {real, imag} */,
  {32'h3f094a32, 32'h405db876} /* (3, 31, 23) {real, imag} */,
  {32'h3f37bb82, 32'h40853850} /* (3, 31, 22) {real, imag} */,
  {32'h3f8dfa78, 32'h403fc80a} /* (3, 31, 21) {real, imag} */,
  {32'h4006992a, 32'hc03ad95e} /* (3, 31, 20) {real, imag} */,
  {32'h3e2c0e0f, 32'hc0321a18} /* (3, 31, 19) {real, imag} */,
  {32'hbd0d90c0, 32'hbe75d1ec} /* (3, 31, 18) {real, imag} */,
  {32'h3f0cf424, 32'hbd904708} /* (3, 31, 17) {real, imag} */,
  {32'h3fa80d52, 32'hc020ca93} /* (3, 31, 16) {real, imag} */,
  {32'h3f76770f, 32'hc010e2c0} /* (3, 31, 15) {real, imag} */,
  {32'h401901b9, 32'hc086ffb0} /* (3, 31, 14) {real, imag} */,
  {32'h3ec7c43c, 32'hc0b4ce6a} /* (3, 31, 13) {real, imag} */,
  {32'h3f0bdd0f, 32'hc096f3d4} /* (3, 31, 12) {real, imag} */,
  {32'h3f2b0a28, 32'hc000717a} /* (3, 31, 11) {real, imag} */,
  {32'h3e1eb758, 32'h408d694a} /* (3, 31, 10) {real, imag} */,
  {32'h3d319ca0, 32'h408e51f2} /* (3, 31, 9) {real, imag} */,
  {32'h3edf2d4d, 32'h40817d77} /* (3, 31, 8) {real, imag} */,
  {32'h3cfb3ac0, 32'h4073c158} /* (3, 31, 7) {real, imag} */,
  {32'hbe696f4e, 32'h40039ab4} /* (3, 31, 6) {real, imag} */,
  {32'hbf3abd8f, 32'h3f915aba} /* (3, 31, 5) {real, imag} */,
  {32'h3eafefbb, 32'h402309d5} /* (3, 31, 4) {real, imag} */,
  {32'h3f84013e, 32'h401e9cc4} /* (3, 31, 3) {real, imag} */,
  {32'hbf5f2439, 32'h402b9034} /* (3, 31, 2) {real, imag} */,
  {32'hc02cd63c, 32'h408b170b} /* (3, 31, 1) {real, imag} */,
  {32'hbf064877, 32'h3fa31383} /* (3, 31, 0) {real, imag} */,
  {32'hbfb544ce, 32'h3f0a03d8} /* (3, 30, 31) {real, imag} */,
  {32'hbee7308c, 32'h3fcae33a} /* (3, 30, 30) {real, imag} */,
  {32'hbf5d86be, 32'h405a15a9} /* (3, 30, 29) {real, imag} */,
  {32'hc0a2ad46, 32'h40d9177b} /* (3, 30, 28) {real, imag} */,
  {32'hc0571a76, 32'h40c5f076} /* (3, 30, 27) {real, imag} */,
  {32'hbf294ad3, 32'h40741462} /* (3, 30, 26) {real, imag} */,
  {32'hc01073da, 32'h40cc82a0} /* (3, 30, 25) {real, imag} */,
  {32'hbff8cc74, 32'h40c13f58} /* (3, 30, 24) {real, imag} */,
  {32'hc043d842, 32'h409bd6d8} /* (3, 30, 23) {real, imag} */,
  {32'hc01c5278, 32'h40b6761d} /* (3, 30, 22) {real, imag} */,
  {32'h3c8bd518, 32'h408bbe38} /* (3, 30, 21) {real, imag} */,
  {32'h407a3a1f, 32'hc0a2724b} /* (3, 30, 20) {real, imag} */,
  {32'h3fbe7a91, 32'hc08deadf} /* (3, 30, 19) {real, imag} */,
  {32'h3f798c5c, 32'hc02ec78a} /* (3, 30, 18) {real, imag} */,
  {32'h3fdac6e0, 32'hc0560ca5} /* (3, 30, 17) {real, imag} */,
  {32'h40551773, 32'hc0b59719} /* (3, 30, 16) {real, imag} */,
  {32'hbece87d9, 32'hc08b6ad6} /* (3, 30, 15) {real, imag} */,
  {32'h406b03d7, 32'hc09e8dc0} /* (3, 30, 14) {real, imag} */,
  {32'h3f9ddd02, 32'hc0db20af} /* (3, 30, 13) {real, imag} */,
  {32'h3f9161e8, 32'hc101e577} /* (3, 30, 12) {real, imag} */,
  {32'h401cc9c0, 32'hc0cadcf4} /* (3, 30, 11) {real, imag} */,
  {32'h3f948c3c, 32'h40696537} /* (3, 30, 10) {real, imag} */,
  {32'h3efb69e8, 32'h40bb95b0} /* (3, 30, 9) {real, imag} */,
  {32'h3f8754d2, 32'h40bd9eb8} /* (3, 30, 8) {real, imag} */,
  {32'h3f5b06be, 32'h40bfb12c} /* (3, 30, 7) {real, imag} */,
  {32'h3eb852ac, 32'h406f5754} /* (3, 30, 6) {real, imag} */,
  {32'hbf646352, 32'h4093d86f} /* (3, 30, 5) {real, imag} */,
  {32'h3f6cc4df, 32'h40cd1018} /* (3, 30, 4) {real, imag} */,
  {32'hbf05ecf7, 32'h40b8dbce} /* (3, 30, 3) {real, imag} */,
  {32'hc000c539, 32'h40bfc374} /* (3, 30, 2) {real, imag} */,
  {32'hc0612333, 32'h40b74cf3} /* (3, 30, 1) {real, imag} */,
  {32'hbfea4ead, 32'h3ff1631d} /* (3, 30, 0) {real, imag} */,
  {32'hc02def62, 32'h401d336b} /* (3, 29, 31) {real, imag} */,
  {32'h3eb79030, 32'h40a5f7f0} /* (3, 29, 30) {real, imag} */,
  {32'h3fc38429, 32'h40b7ea9c} /* (3, 29, 29) {real, imag} */,
  {32'hc09edc68, 32'h40af1d68} /* (3, 29, 28) {real, imag} */,
  {32'hc064871a, 32'h40ad6af9} /* (3, 29, 27) {real, imag} */,
  {32'h3eacc596, 32'h40c71a10} /* (3, 29, 26) {real, imag} */,
  {32'hbf82a415, 32'h40f94aee} /* (3, 29, 25) {real, imag} */,
  {32'hbfc57e52, 32'h40b9e780} /* (3, 29, 24) {real, imag} */,
  {32'hbf5d3aa8, 32'h40492a25} /* (3, 29, 23) {real, imag} */,
  {32'hbfc5a17d, 32'h40a7f4f8} /* (3, 29, 22) {real, imag} */,
  {32'hbff68f01, 32'h408262c3} /* (3, 29, 21) {real, imag} */,
  {32'h403551fc, 32'hc0cb400c} /* (3, 29, 20) {real, imag} */,
  {32'h4087edda, 32'hc0f6616e} /* (3, 29, 19) {real, imag} */,
  {32'h406cc163, 32'hc0b90aa1} /* (3, 29, 18) {real, imag} */,
  {32'h3fba669a, 32'hc09d776d} /* (3, 29, 17) {real, imag} */,
  {32'h3ffa4dbe, 32'hc097cfca} /* (3, 29, 16) {real, imag} */,
  {32'hbf8706ae, 32'hc0b3faae} /* (3, 29, 15) {real, imag} */,
  {32'h402c73e8, 32'hc0c3fef0} /* (3, 29, 14) {real, imag} */,
  {32'h3f68f91b, 32'hc093d4bd} /* (3, 29, 13) {real, imag} */,
  {32'h3f7541cc, 32'hc0f24cd8} /* (3, 29, 12) {real, imag} */,
  {32'h3ff78d4b, 32'hc0cd30e4} /* (3, 29, 11) {real, imag} */,
  {32'hbf6e20ec, 32'h403bb69e} /* (3, 29, 10) {real, imag} */,
  {32'hc033defa, 32'h40ae6c4e} /* (3, 29, 9) {real, imag} */,
  {32'hbfd8b5be, 32'h40b76ff5} /* (3, 29, 8) {real, imag} */,
  {32'hbefa651c, 32'h40ae6494} /* (3, 29, 7) {real, imag} */,
  {32'h3b387400, 32'h401edf16} /* (3, 29, 6) {real, imag} */,
  {32'hc06e3917, 32'h40431da6} /* (3, 29, 5) {real, imag} */,
  {32'hbfb8470e, 32'h40c8a480} /* (3, 29, 4) {real, imag} */,
  {32'h3f0bcb7a, 32'h40f55459} /* (3, 29, 3) {real, imag} */,
  {32'hbf0bd209, 32'h40de12c5} /* (3, 29, 2) {real, imag} */,
  {32'hbf6b584c, 32'h40222eec} /* (3, 29, 1) {real, imag} */,
  {32'hbfbc23d4, 32'hbeb79dd4} /* (3, 29, 0) {real, imag} */,
  {32'hbfde23e8, 32'h407d8172} /* (3, 28, 31) {real, imag} */,
  {32'h3f44b39e, 32'h40f2f644} /* (3, 28, 30) {real, imag} */,
  {32'h3f0f2800, 32'h40e6bd12} /* (3, 28, 29) {real, imag} */,
  {32'hc0901b98, 32'h40309942} /* (3, 28, 28) {real, imag} */,
  {32'hbfaf7cb6, 32'h40874a9a} /* (3, 28, 27) {real, imag} */,
  {32'h3faa1aec, 32'h40d8e472} /* (3, 28, 26) {real, imag} */,
  {32'h3f5724f2, 32'h409828fb} /* (3, 28, 25) {real, imag} */,
  {32'hbf628b81, 32'h40202446} /* (3, 28, 24) {real, imag} */,
  {32'hbf9efbf2, 32'h4039880a} /* (3, 28, 23) {real, imag} */,
  {32'hc08b3c32, 32'h40d54f00} /* (3, 28, 22) {real, imag} */,
  {32'hc0c08e16, 32'h40869d4b} /* (3, 28, 21) {real, imag} */,
  {32'h3fef62e9, 32'hc0a59976} /* (3, 28, 20) {real, imag} */,
  {32'h40b8348d, 32'hc108fce5} /* (3, 28, 19) {real, imag} */,
  {32'h40049d60, 32'hc0a4f019} /* (3, 28, 18) {real, imag} */,
  {32'h3f45f52a, 32'hc04df096} /* (3, 28, 17) {real, imag} */,
  {32'h3fd474ef, 32'hc04f392f} /* (3, 28, 16) {real, imag} */,
  {32'h3f851f82, 32'hc0a1456c} /* (3, 28, 15) {real, imag} */,
  {32'h3fb2704c, 32'hc0c64dac} /* (3, 28, 14) {real, imag} */,
  {32'h3e9965ba, 32'hc0ad9486} /* (3, 28, 13) {real, imag} */,
  {32'h3eff8202, 32'hc0c0500f} /* (3, 28, 12) {real, imag} */,
  {32'hbe8beb17, 32'hc0a1f3dd} /* (3, 28, 11) {real, imag} */,
  {32'hc0a4daf1, 32'h40834e07} /* (3, 28, 10) {real, imag} */,
  {32'hc0b94788, 32'h40f1d89a} /* (3, 28, 9) {real, imag} */,
  {32'hc0a4e688, 32'h410319ca} /* (3, 28, 8) {real, imag} */,
  {32'hc05485d9, 32'h40f251f5} /* (3, 28, 7) {real, imag} */,
  {32'hbf942c08, 32'h3ff2889a} /* (3, 28, 6) {real, imag} */,
  {32'hc07991f3, 32'h4041c93e} /* (3, 28, 5) {real, imag} */,
  {32'hbf70caa1, 32'h40ea0ae4} /* (3, 28, 4) {real, imag} */,
  {32'h3ede7f90, 32'h411ed1dc} /* (3, 28, 3) {real, imag} */,
  {32'h3e1ae764, 32'h40d1891d} /* (3, 28, 2) {real, imag} */,
  {32'h3fe790f2, 32'h400d925f} /* (3, 28, 1) {real, imag} */,
  {32'hbfc6f680, 32'h3f81d8f0} /* (3, 28, 0) {real, imag} */,
  {32'h3e7515c0, 32'h3ffeaeb5} /* (3, 27, 31) {real, imag} */,
  {32'h3f203383, 32'h40372341} /* (3, 27, 30) {real, imag} */,
  {32'hbeb1a052, 32'h4056a084} /* (3, 27, 29) {real, imag} */,
  {32'hc085e5da, 32'h40325fd3} /* (3, 27, 28) {real, imag} */,
  {32'hbf95c87f, 32'h40ddeae0} /* (3, 27, 27) {real, imag} */,
  {32'h3fd567a4, 32'h41219ab9} /* (3, 27, 26) {real, imag} */,
  {32'h40286f50, 32'h40cc28ac} /* (3, 27, 25) {real, imag} */,
  {32'h3f1e7969, 32'h40a17f90} /* (3, 27, 24) {real, imag} */,
  {32'hbf39f02c, 32'h40840a53} /* (3, 27, 23) {real, imag} */,
  {32'hc026ca4a, 32'h408fb5f6} /* (3, 27, 22) {real, imag} */,
  {32'hc0af1a89, 32'h4023bc00} /* (3, 27, 21) {real, imag} */,
  {32'hbeb568d8, 32'hc0ad9c68} /* (3, 27, 20) {real, imag} */,
  {32'h3faf7631, 32'hc105feac} /* (3, 27, 19) {real, imag} */,
  {32'h3f83720a, 32'hc0dfa610} /* (3, 27, 18) {real, imag} */,
  {32'h40184354, 32'hc08d83c0} /* (3, 27, 17) {real, imag} */,
  {32'h3f122cae, 32'hc0890d88} /* (3, 27, 16) {real, imag} */,
  {32'hbf8bce37, 32'hc0559b8f} /* (3, 27, 15) {real, imag} */,
  {32'hbed32a52, 32'hc04e5475} /* (3, 27, 14) {real, imag} */,
  {32'h3fe47c68, 32'hc0f53bf4} /* (3, 27, 13) {real, imag} */,
  {32'h3fe668ad, 32'hc0bde93c} /* (3, 27, 12) {real, imag} */,
  {32'hbf37daff, 32'hc09fe602} /* (3, 27, 11) {real, imag} */,
  {32'hc05d752e, 32'h4065fd16} /* (3, 27, 10) {real, imag} */,
  {32'hc01ec614, 32'h41000dfa} /* (3, 27, 9) {real, imag} */,
  {32'hc06e4d5e, 32'h40c0a397} /* (3, 27, 8) {real, imag} */,
  {32'hc01be1e9, 32'h40c1d964} /* (3, 27, 7) {real, imag} */,
  {32'hbfdd9e1a, 32'h4008d24a} /* (3, 27, 6) {real, imag} */,
  {32'hc07a72ed, 32'h4091dd0a} /* (3, 27, 5) {real, imag} */,
  {32'hbd046d78, 32'h41036f99} /* (3, 27, 4) {real, imag} */,
  {32'hbf768735, 32'h411ef222} /* (3, 27, 3) {real, imag} */,
  {32'hc01a895e, 32'h40d645ae} /* (3, 27, 2) {real, imag} */,
  {32'h3f22de14, 32'h4066f10e} /* (3, 27, 1) {real, imag} */,
  {32'h3e9bf91b, 32'h4018a690} /* (3, 27, 0) {real, imag} */,
  {32'hbceb5dd0, 32'h400457b9} /* (3, 26, 31) {real, imag} */,
  {32'h3dc4dc20, 32'h405ebd8d} /* (3, 26, 30) {real, imag} */,
  {32'h3cf4c940, 32'h40c8cb48} /* (3, 26, 29) {real, imag} */,
  {32'hc01d38c2, 32'h408f6f5c} /* (3, 26, 28) {real, imag} */,
  {32'hc00f8aa4, 32'h40ce955a} /* (3, 26, 27) {real, imag} */,
  {32'hbfccb0e0, 32'h40fc4f95} /* (3, 26, 26) {real, imag} */,
  {32'h3ffdc514, 32'h40b2aae2} /* (3, 26, 25) {real, imag} */,
  {32'h3f43085e, 32'h41021434} /* (3, 26, 24) {real, imag} */,
  {32'hc02c0808, 32'h40a9b795} /* (3, 26, 23) {real, imag} */,
  {32'hc0343645, 32'h40578528} /* (3, 26, 22) {real, imag} */,
  {32'hbfd25ef6, 32'h3fd1bad5} /* (3, 26, 21) {real, imag} */,
  {32'h3f908fe6, 32'hc0c8b6b0} /* (3, 26, 20) {real, imag} */,
  {32'h40199b31, 32'hc0e15986} /* (3, 26, 19) {real, imag} */,
  {32'h4081173d, 32'hc0d9e55a} /* (3, 26, 18) {real, imag} */,
  {32'h408616ed, 32'hc0bdf192} /* (3, 26, 17) {real, imag} */,
  {32'h3e0b9268, 32'hc090789e} /* (3, 26, 16) {real, imag} */,
  {32'hbfac4c58, 32'hc0a81742} /* (3, 26, 15) {real, imag} */,
  {32'h3f93c0f1, 32'hc09652df} /* (3, 26, 14) {real, imag} */,
  {32'h406a1186, 32'hc0845b7a} /* (3, 26, 13) {real, imag} */,
  {32'h40612a9b, 32'hc0672fe2} /* (3, 26, 12) {real, imag} */,
  {32'h4046d639, 32'hc03d0f46} /* (3, 26, 11) {real, imag} */,
  {32'hbf178a45, 32'h3faa64f0} /* (3, 26, 10) {real, imag} */,
  {32'hc0219b78, 32'h40ed009f} /* (3, 26, 9) {real, imag} */,
  {32'hbf6a3b5a, 32'h40597766} /* (3, 26, 8) {real, imag} */,
  {32'hbef6141c, 32'h3fe9268a} /* (3, 26, 7) {real, imag} */,
  {32'hbfde61f7, 32'h3ff90f3e} /* (3, 26, 6) {real, imag} */,
  {32'hbf620598, 32'h4049275a} /* (3, 26, 5) {real, imag} */,
  {32'hbf67a844, 32'h40956d2a} /* (3, 26, 4) {real, imag} */,
  {32'hbfdc7822, 32'h409c3c6f} /* (3, 26, 3) {real, imag} */,
  {32'hbf3d4e36, 32'h408bb40f} /* (3, 26, 2) {real, imag} */,
  {32'hbf2aa87c, 32'h404c6ad2} /* (3, 26, 1) {real, imag} */,
  {32'h3eeabc78, 32'h40182784} /* (3, 26, 0) {real, imag} */,
  {32'hbfaf1b18, 32'h407d9958} /* (3, 25, 31) {real, imag} */,
  {32'hbf3eda1c, 32'h40ea79e0} /* (3, 25, 30) {real, imag} */,
  {32'hbe50191c, 32'h40d56060} /* (3, 25, 29) {real, imag} */,
  {32'hbcd91310, 32'h409d67ce} /* (3, 25, 28) {real, imag} */,
  {32'hc007c7da, 32'h409bb400} /* (3, 25, 27) {real, imag} */,
  {32'hc003e261, 32'h40c410a1} /* (3, 25, 26) {real, imag} */,
  {32'h3ffc8561, 32'h40ca16a4} /* (3, 25, 25) {real, imag} */,
  {32'h3e3d7fa8, 32'h40d7a09d} /* (3, 25, 24) {real, imag} */,
  {32'hc0458c02, 32'h40a85d4b} /* (3, 25, 23) {real, imag} */,
  {32'hc0326a71, 32'h40563d19} /* (3, 25, 22) {real, imag} */,
  {32'hbfc55014, 32'hbfcbc695} /* (3, 25, 21) {real, imag} */,
  {32'hbf4df390, 32'hc0d2f698} /* (3, 25, 20) {real, imag} */,
  {32'h3fed69ac, 32'hc092dd1a} /* (3, 25, 19) {real, imag} */,
  {32'h4080ec14, 32'hc0be22f5} /* (3, 25, 18) {real, imag} */,
  {32'hbf2732c2, 32'hc0c11eda} /* (3, 25, 17) {real, imag} */,
  {32'hbf97bebe, 32'hc073f4ec} /* (3, 25, 16) {real, imag} */,
  {32'h40201f26, 32'hc0eb703e} /* (3, 25, 15) {real, imag} */,
  {32'h40a32925, 32'hc11ee4d0} /* (3, 25, 14) {real, imag} */,
  {32'h3feb7421, 32'hc01dc00c} /* (3, 25, 13) {real, imag} */,
  {32'h3f72cb7d, 32'hbfcbd431} /* (3, 25, 12) {real, imag} */,
  {32'h3dea0cf5, 32'hc0306052} /* (3, 25, 11) {real, imag} */,
  {32'hbfc5b5c0, 32'h4013c836} /* (3, 25, 10) {real, imag} */,
  {32'hc04b058a, 32'h40d3851c} /* (3, 25, 9) {real, imag} */,
  {32'hc04a840c, 32'h40b052f4} /* (3, 25, 8) {real, imag} */,
  {32'hbff3f80a, 32'h40929998} /* (3, 25, 7) {real, imag} */,
  {32'hbfdc859a, 32'h40a36bbe} /* (3, 25, 6) {real, imag} */,
  {32'h3e8d8eea, 32'h40f9ec00} /* (3, 25, 5) {real, imag} */,
  {32'h3e99b21c, 32'h40fe0274} /* (3, 25, 4) {real, imag} */,
  {32'h3edb95f5, 32'h40946513} /* (3, 25, 3) {real, imag} */,
  {32'h3f0c61bc, 32'h402cebf0} /* (3, 25, 2) {real, imag} */,
  {32'hbfb568c6, 32'h3f107271} /* (3, 25, 1) {real, imag} */,
  {32'hbf407f32, 32'h40259504} /* (3, 25, 0) {real, imag} */,
  {32'hbecfa7da, 32'h406b466e} /* (3, 24, 31) {real, imag} */,
  {32'hbf84d274, 32'h410d8ece} /* (3, 24, 30) {real, imag} */,
  {32'h3e08c794, 32'h40a8356b} /* (3, 24, 29) {real, imag} */,
  {32'h3ef19bc0, 32'h40a679d4} /* (3, 24, 28) {real, imag} */,
  {32'hc0148564, 32'h40bb1b7e} /* (3, 24, 27) {real, imag} */,
  {32'h3e163950, 32'h40fe03d0} /* (3, 24, 26) {real, imag} */,
  {32'h3fa38c62, 32'h41117cb7} /* (3, 24, 25) {real, imag} */,
  {32'hbffe1d74, 32'h406ce2ab} /* (3, 24, 24) {real, imag} */,
  {32'hc083eecb, 32'h407e125a} /* (3, 24, 23) {real, imag} */,
  {32'hc0318fee, 32'h40802488} /* (3, 24, 22) {real, imag} */,
  {32'hc059f07f, 32'h3ec92274} /* (3, 24, 21) {real, imag} */,
  {32'hc03d11fe, 32'hc09ed97c} /* (3, 24, 20) {real, imag} */,
  {32'h3f3c392d, 32'hc099d75a} /* (3, 24, 19) {real, imag} */,
  {32'h40293788, 32'hc0bea5ea} /* (3, 24, 18) {real, imag} */,
  {32'hbed1ddac, 32'hc08c15cc} /* (3, 24, 17) {real, imag} */,
  {32'h4041cd07, 32'hc0774f7c} /* (3, 24, 16) {real, imag} */,
  {32'h409e5f72, 32'hc0fc1686} /* (3, 24, 15) {real, imag} */,
  {32'h40c1a9c1, 32'hc11e1afe} /* (3, 24, 14) {real, imag} */,
  {32'h3f65d0cc, 32'hc0601c00} /* (3, 24, 13) {real, imag} */,
  {32'hbeaf6ac8, 32'hbfcf5082} /* (3, 24, 12) {real, imag} */,
  {32'h3ef0458a, 32'hbf98d3b2} /* (3, 24, 11) {real, imag} */,
  {32'h3f075db3, 32'h40a18718} /* (3, 24, 10) {real, imag} */,
  {32'hbf1c25bb, 32'h40bdd440} /* (3, 24, 9) {real, imag} */,
  {32'hc08c2a00, 32'h40ac2238} /* (3, 24, 8) {real, imag} */,
  {32'hbff4186e, 32'h40c750fa} /* (3, 24, 7) {real, imag} */,
  {32'hbfb07c76, 32'h40dbc094} /* (3, 24, 6) {real, imag} */,
  {32'h3c1ba2c0, 32'h40e97b70} /* (3, 24, 5) {real, imag} */,
  {32'h3f3874e0, 32'h409d7ad9} /* (3, 24, 4) {real, imag} */,
  {32'h3ef25373, 32'h40d4302c} /* (3, 24, 3) {real, imag} */,
  {32'h3ffc1394, 32'h40e82fdf} /* (3, 24, 2) {real, imag} */,
  {32'h3f02eb5a, 32'h4081d758} /* (3, 24, 1) {real, imag} */,
  {32'h3ebf2cda, 32'h403add63} /* (3, 24, 0) {real, imag} */,
  {32'hbf69442f, 32'h408132f6} /* (3, 23, 31) {real, imag} */,
  {32'hc030dce4, 32'h40c4ecd6} /* (3, 23, 30) {real, imag} */,
  {32'hbfcaaf24, 32'h40bd589c} /* (3, 23, 29) {real, imag} */,
  {32'hbf22389d, 32'h40a69e34} /* (3, 23, 28) {real, imag} */,
  {32'hc04413cf, 32'h41070e10} /* (3, 23, 27) {real, imag} */,
  {32'hbfaada2a, 32'h410c4b3c} /* (3, 23, 26) {real, imag} */,
  {32'hbd93c438, 32'h40db12a7} /* (3, 23, 25) {real, imag} */,
  {32'hbfd6898c, 32'h40085fd0} /* (3, 23, 24) {real, imag} */,
  {32'hc005dcba, 32'h4083cca2} /* (3, 23, 23) {real, imag} */,
  {32'hc006e09c, 32'h40a25fc1} /* (3, 23, 22) {real, imag} */,
  {32'hc063a0e8, 32'h3fd41efe} /* (3, 23, 21) {real, imag} */,
  {32'hc022e8de, 32'hc0750465} /* (3, 23, 20) {real, imag} */,
  {32'hbf01dd62, 32'hc0b54a40} /* (3, 23, 19) {real, imag} */,
  {32'hbf005f81, 32'hc0cccd82} /* (3, 23, 18) {real, imag} */,
  {32'hbe480b5c, 32'hc0aa0abe} /* (3, 23, 17) {real, imag} */,
  {32'h4032d2fc, 32'hc004819a} /* (3, 23, 16) {real, imag} */,
  {32'h3d8b6708, 32'hc08d148e} /* (3, 23, 15) {real, imag} */,
  {32'h3fb63798, 32'hc0fe4697} /* (3, 23, 14) {real, imag} */,
  {32'h3fb63d7a, 32'hc079dbd4} /* (3, 23, 13) {real, imag} */,
  {32'h401de69e, 32'hbfc44fba} /* (3, 23, 12) {real, imag} */,
  {32'h3f568fc0, 32'hc06e2ee9} /* (3, 23, 11) {real, imag} */,
  {32'hbe06b5ee, 32'h3fc7fd36} /* (3, 23, 10) {real, imag} */,
  {32'h3fe89e28, 32'h40b151ac} /* (3, 23, 9) {real, imag} */,
  {32'hbfefe5e8, 32'h40cdc9a5} /* (3, 23, 8) {real, imag} */,
  {32'hc0137507, 32'h40fcf237} /* (3, 23, 7) {real, imag} */,
  {32'h3f30e700, 32'h40bb2d28} /* (3, 23, 6) {real, imag} */,
  {32'hbed9377a, 32'h40a8e7a5} /* (3, 23, 5) {real, imag} */,
  {32'hbf6c3daa, 32'h40838c8a} /* (3, 23, 4) {real, imag} */,
  {32'h3ed46497, 32'h40c5bb74} /* (3, 23, 3) {real, imag} */,
  {32'h401e4263, 32'h40ce9a8c} /* (3, 23, 2) {real, imag} */,
  {32'h40082e3b, 32'h40c8ed6f} /* (3, 23, 1) {real, imag} */,
  {32'h3fc12d42, 32'h408f58a4} /* (3, 23, 0) {real, imag} */,
  {32'hbf60637c, 32'h4013a220} /* (3, 22, 31) {real, imag} */,
  {32'hbf2b9c69, 32'h4082ccc8} /* (3, 22, 30) {real, imag} */,
  {32'hbff8a947, 32'h40bef31b} /* (3, 22, 29) {real, imag} */,
  {32'hc05b74e0, 32'h40742bb2} /* (3, 22, 28) {real, imag} */,
  {32'hc0a66d03, 32'h40b3e254} /* (3, 22, 27) {real, imag} */,
  {32'hc006bc85, 32'h40c0e5b2} /* (3, 22, 26) {real, imag} */,
  {32'hbde416b8, 32'h40bd3c61} /* (3, 22, 25) {real, imag} */,
  {32'h3e6be200, 32'h40add610} /* (3, 22, 24) {real, imag} */,
  {32'h3ea35d9f, 32'h40b853b7} /* (3, 22, 23) {real, imag} */,
  {32'hbf201a46, 32'h4099e864} /* (3, 22, 22) {real, imag} */,
  {32'hbf19cc94, 32'h407dc18a} /* (3, 22, 21) {real, imag} */,
  {32'hbe249e96, 32'hc07c17ce} /* (3, 22, 20) {real, imag} */,
  {32'hbf93f0e0, 32'hc0e59640} /* (3, 22, 19) {real, imag} */,
  {32'hc0136e42, 32'hc0bc1b2e} /* (3, 22, 18) {real, imag} */,
  {32'hbfc94d88, 32'hc081d5f2} /* (3, 22, 17) {real, imag} */,
  {32'h3ffdad48, 32'hc03d4d4e} /* (3, 22, 16) {real, imag} */,
  {32'h3eda28df, 32'hc06d4526} /* (3, 22, 15) {real, imag} */,
  {32'hbf00d638, 32'hc0ee6f89} /* (3, 22, 14) {real, imag} */,
  {32'h40011dfe, 32'hc0c854c8} /* (3, 22, 13) {real, imag} */,
  {32'h404f3072, 32'hc03cdc2e} /* (3, 22, 12) {real, imag} */,
  {32'h3ea74c55, 32'hbfd8564e} /* (3, 22, 11) {real, imag} */,
  {32'hbfe446b9, 32'h403c29e0} /* (3, 22, 10) {real, imag} */,
  {32'h3eaf3140, 32'h408af502} /* (3, 22, 9) {real, imag} */,
  {32'hbff8f87a, 32'h407e2c2a} /* (3, 22, 8) {real, imag} */,
  {32'hc0215e9e, 32'h40b8bb97} /* (3, 22, 7) {real, imag} */,
  {32'hbf7b5874, 32'h40b7d416} /* (3, 22, 6) {real, imag} */,
  {32'hbf999740, 32'h40e511f6} /* (3, 22, 5) {real, imag} */,
  {32'hbf8d275e, 32'h40a8b746} /* (3, 22, 4) {real, imag} */,
  {32'hbecbcee4, 32'h40f68bfe} /* (3, 22, 3) {real, imag} */,
  {32'h3ffdb84e, 32'h40a9abae} /* (3, 22, 2) {real, imag} */,
  {32'h3eabb3f5, 32'h40195e2a} /* (3, 22, 1) {real, imag} */,
  {32'hbd8a282e, 32'h40196510} /* (3, 22, 0) {real, imag} */,
  {32'hbf638c8f, 32'h3e9c2771} /* (3, 21, 31) {real, imag} */,
  {32'hbec2c233, 32'h3f2102f0} /* (3, 21, 30) {real, imag} */,
  {32'hbe0623f0, 32'h3fac584d} /* (3, 21, 29) {real, imag} */,
  {32'hc0134002, 32'h400e4c96} /* (3, 21, 28) {real, imag} */,
  {32'hbf801725, 32'h40218ee3} /* (3, 21, 27) {real, imag} */,
  {32'h40236db2, 32'h3fd5f0b8} /* (3, 21, 26) {real, imag} */,
  {32'h3fa2c210, 32'h40045f50} /* (3, 21, 25) {real, imag} */,
  {32'hbe1f9e4c, 32'h3f7f50ae} /* (3, 21, 24) {real, imag} */,
  {32'hbd4350d4, 32'h3fa42e6c} /* (3, 21, 23) {real, imag} */,
  {32'hbf351d7b, 32'hbee3a63a} /* (3, 21, 22) {real, imag} */,
  {32'h3e7a7991, 32'h4007db9d} /* (3, 21, 21) {real, imag} */,
  {32'hbff667ef, 32'hc0288880} /* (3, 21, 20) {real, imag} */,
  {32'hc07c1d8a, 32'hc0599368} /* (3, 21, 19) {real, imag} */,
  {32'hc002a86d, 32'hc04aac98} /* (3, 21, 18) {real, imag} */,
  {32'hc0019fb6, 32'hc061f3c4} /* (3, 21, 17) {real, imag} */,
  {32'h3feb3220, 32'hc0493bda} /* (3, 21, 16) {real, imag} */,
  {32'h3f8a307c, 32'hc00c5a8c} /* (3, 21, 15) {real, imag} */,
  {32'hbf4d894e, 32'hc08d7af2} /* (3, 21, 14) {real, imag} */,
  {32'h3fd7f5cd, 32'hc0379ba7} /* (3, 21, 13) {real, imag} */,
  {32'h4079c864, 32'hbfbcdeae} /* (3, 21, 12) {real, imag} */,
  {32'h3f9468ab, 32'h3eb4e695} /* (3, 21, 11) {real, imag} */,
  {32'hc04a70d0, 32'h402c9dea} /* (3, 21, 10) {real, imag} */,
  {32'h3e7972c2, 32'h3ff3c444} /* (3, 21, 9) {real, imag} */,
  {32'h3e30d28c, 32'h3f5e4f79} /* (3, 21, 8) {real, imag} */,
  {32'hc021b1e4, 32'h3f4bcb25} /* (3, 21, 7) {real, imag} */,
  {32'hc018c56b, 32'h3fae4ed4} /* (3, 21, 6) {real, imag} */,
  {32'hbee90c91, 32'h4035d740} /* (3, 21, 5) {real, imag} */,
  {32'hbe9c9d84, 32'h40357de7} /* (3, 21, 4) {real, imag} */,
  {32'h3ee258f9, 32'h408b5126} /* (3, 21, 3) {real, imag} */,
  {32'h3f17bece, 32'h400ec0c6} /* (3, 21, 2) {real, imag} */,
  {32'hc0091ee3, 32'h3ddc529c} /* (3, 21, 1) {real, imag} */,
  {32'hc0057da2, 32'h3e367b26} /* (3, 21, 0) {real, imag} */,
  {32'hbf14b2bc, 32'hc02d7bdc} /* (3, 20, 31) {real, imag} */,
  {32'hbfcf166a, 32'hc0a373ea} /* (3, 20, 30) {real, imag} */,
  {32'h402447a6, 32'hc0c433ce} /* (3, 20, 29) {real, imag} */,
  {32'h40235fdc, 32'hc0646992} /* (3, 20, 28) {real, imag} */,
  {32'h40926ac2, 32'hc063a1f6} /* (3, 20, 27) {real, imag} */,
  {32'h409a51cd, 32'hc0aff5ec} /* (3, 20, 26) {real, imag} */,
  {32'h40a8f873, 32'hc0f91b59} /* (3, 20, 25) {real, imag} */,
  {32'h3f762dd8, 32'hc1158cc2} /* (3, 20, 24) {real, imag} */,
  {32'hbf824351, 32'hc0f9b904} /* (3, 20, 23) {real, imag} */,
  {32'h3e11132e, 32'hc0a5687a} /* (3, 20, 22) {real, imag} */,
  {32'hbd5b9b20, 32'hbfff5a47} /* (3, 20, 21) {real, imag} */,
  {32'hbfd41847, 32'h4043f9aa} /* (3, 20, 20) {real, imag} */,
  {32'hc0901cb9, 32'h408862ce} /* (3, 20, 19) {real, imag} */,
  {32'hc09c67d9, 32'h404efeb6} /* (3, 20, 18) {real, imag} */,
  {32'hc09a26d6, 32'h406cfeb0} /* (3, 20, 17) {real, imag} */,
  {32'hc0037637, 32'h404aa1a1} /* (3, 20, 16) {real, imag} */,
  {32'hbfe1d432, 32'h4064f980} /* (3, 20, 15) {real, imag} */,
  {32'hbfe89bc0, 32'h407007aa} /* (3, 20, 14) {real, imag} */,
  {32'hbea523e7, 32'h40ab1c44} /* (3, 20, 13) {real, imag} */,
  {32'h40212432, 32'h4035a3cd} /* (3, 20, 12) {real, imag} */,
  {32'hbe8c20ce, 32'h3f0fc6ee} /* (3, 20, 11) {real, imag} */,
  {32'hc00e02f1, 32'hbe0a5984} /* (3, 20, 10) {real, imag} */,
  {32'h3ec845bf, 32'hc052377f} /* (3, 20, 9) {real, imag} */,
  {32'hbde4a018, 32'hc09842e3} /* (3, 20, 8) {real, imag} */,
  {32'hbfcbb702, 32'hc0bb399e} /* (3, 20, 7) {real, imag} */,
  {32'h3c967a40, 32'hc0d0f33c} /* (3, 20, 6) {real, imag} */,
  {32'h3fa78757, 32'hc0a2da33} /* (3, 20, 5) {real, imag} */,
  {32'h4010469a, 32'hc0c3c12b} /* (3, 20, 4) {real, imag} */,
  {32'h40278782, 32'hc0979f28} /* (3, 20, 3) {real, imag} */,
  {32'h3fda2fe3, 32'hc04c49be} /* (3, 20, 2) {real, imag} */,
  {32'hbfcef41c, 32'hc08c92a8} /* (3, 20, 1) {real, imag} */,
  {32'hbfe6505b, 32'hbf8f4962} /* (3, 20, 0) {real, imag} */,
  {32'h3f2be11c, 32'hc0b182bc} /* (3, 19, 31) {real, imag} */,
  {32'hbfca5dfe, 32'hc0c0d088} /* (3, 19, 30) {real, imag} */,
  {32'h3fde29d7, 32'hc079b290} /* (3, 19, 29) {real, imag} */,
  {32'h3ffeb5a3, 32'hc087e267} /* (3, 19, 28) {real, imag} */,
  {32'h40956758, 32'hc086d96a} /* (3, 19, 27) {real, imag} */,
  {32'h40041548, 32'hc0bba6a6} /* (3, 19, 26) {real, imag} */,
  {32'h40541987, 32'hc0d1ddaa} /* (3, 19, 25) {real, imag} */,
  {32'h40372f08, 32'hc0c1e542} /* (3, 19, 24) {real, imag} */,
  {32'h3fe0b42c, 32'hc0d7632e} /* (3, 19, 23) {real, imag} */,
  {32'h3f694bb1, 32'hc0e38736} /* (3, 19, 22) {real, imag} */,
  {32'hbf83d3e1, 32'hc0183be2} /* (3, 19, 21) {real, imag} */,
  {32'hbf3ef815, 32'h408ca3ea} /* (3, 19, 20) {real, imag} */,
  {32'hbff7b877, 32'h406d5010} /* (3, 19, 19) {real, imag} */,
  {32'hc0806fa6, 32'h40a6b9fc} /* (3, 19, 18) {real, imag} */,
  {32'hc0715701, 32'h40e0334a} /* (3, 19, 17) {real, imag} */,
  {32'hc0385063, 32'h408e93c4} /* (3, 19, 16) {real, imag} */,
  {32'hbf9e94b0, 32'h405c283e} /* (3, 19, 15) {real, imag} */,
  {32'hc01936b4, 32'h40b7712d} /* (3, 19, 14) {real, imag} */,
  {32'hc087197e, 32'h40fd2aae} /* (3, 19, 13) {real, imag} */,
  {32'hc01434d1, 32'h40c38558} /* (3, 19, 12) {real, imag} */,
  {32'hbf4de5db, 32'h4039efd4} /* (3, 19, 11) {real, imag} */,
  {32'hc020fc66, 32'hc04c437c} /* (3, 19, 10) {real, imag} */,
  {32'hc040649e, 32'hc0c59909} /* (3, 19, 9) {real, imag} */,
  {32'hbf777267, 32'hc1011f99} /* (3, 19, 8) {real, imag} */,
  {32'hbf859eb4, 32'hc0d58af7} /* (3, 19, 7) {real, imag} */,
  {32'h3f3050bc, 32'hc0b8972e} /* (3, 19, 6) {real, imag} */,
  {32'h3fad9290, 32'hc0d64199} /* (3, 19, 5) {real, imag} */,
  {32'h400eafd9, 32'hc0d0dd1b} /* (3, 19, 4) {real, imag} */,
  {32'h4053f36a, 32'hc0cc6d56} /* (3, 19, 3) {real, imag} */,
  {32'h404d1b97, 32'hc0964aaf} /* (3, 19, 2) {real, imag} */,
  {32'hbead93a2, 32'hc096c350} /* (3, 19, 1) {real, imag} */,
  {32'h3e6db6f6, 32'hc0088f29} /* (3, 19, 0) {real, imag} */,
  {32'hbfa291cf, 32'hc0cdc03e} /* (3, 18, 31) {real, imag} */,
  {32'hbe3d9f90, 32'hc0e2ea12} /* (3, 18, 30) {real, imag} */,
  {32'h3f28ac68, 32'hc07408a4} /* (3, 18, 29) {real, imag} */,
  {32'hbf0f346c, 32'hc0984229} /* (3, 18, 28) {real, imag} */,
  {32'h40052839, 32'hc0b468fe} /* (3, 18, 27) {real, imag} */,
  {32'h3faf4a5e, 32'hc0bb6a34} /* (3, 18, 26) {real, imag} */,
  {32'h4042e15a, 32'hc08d321b} /* (3, 18, 25) {real, imag} */,
  {32'h403565d8, 32'hc09d934e} /* (3, 18, 24) {real, imag} */,
  {32'h403a854e, 32'hc08a5c54} /* (3, 18, 23) {real, imag} */,
  {32'h40039e74, 32'hc0a301e7} /* (3, 18, 22) {real, imag} */,
  {32'hbfc30d8f, 32'hc009ce51} /* (3, 18, 21) {real, imag} */,
  {32'h3ee1c54a, 32'h40d7f2e8} /* (3, 18, 20) {real, imag} */,
  {32'hbfa50815, 32'h40ab65fe} /* (3, 18, 19) {real, imag} */,
  {32'hc09ca92f, 32'h40aee8a7} /* (3, 18, 18) {real, imag} */,
  {32'hc089188e, 32'h40c80b48} /* (3, 18, 17) {real, imag} */,
  {32'hc07dabda, 32'h40564dd3} /* (3, 18, 16) {real, imag} */,
  {32'hc012a05b, 32'h40a353ba} /* (3, 18, 15) {real, imag} */,
  {32'hc042b0aa, 32'h4105da74} /* (3, 18, 14) {real, imag} */,
  {32'hc03b30aa, 32'h4106b9a8} /* (3, 18, 13) {real, imag} */,
  {32'hc0015ce6, 32'h40e3b5d5} /* (3, 18, 12) {real, imag} */,
  {32'hbf47dcf2, 32'h409258f6} /* (3, 18, 11) {real, imag} */,
  {32'hc026fcc2, 32'hc0278d26} /* (3, 18, 10) {real, imag} */,
  {32'hc0344b7f, 32'hc0bafd5c} /* (3, 18, 9) {real, imag} */,
  {32'h3f01c9e9, 32'hc0e2f7e0} /* (3, 18, 8) {real, imag} */,
  {32'h3f1e3130, 32'hc0de18ac} /* (3, 18, 7) {real, imag} */,
  {32'h3fa2f134, 32'hc0901cc7} /* (3, 18, 6) {real, imag} */,
  {32'h3fe321b8, 32'hc0669469} /* (3, 18, 5) {real, imag} */,
  {32'h3f28383c, 32'hc088e7d4} /* (3, 18, 4) {real, imag} */,
  {32'h3fd89e92, 32'hc0c03108} /* (3, 18, 3) {real, imag} */,
  {32'h3f790fa4, 32'hc0c406ae} /* (3, 18, 2) {real, imag} */,
  {32'h3e83e67c, 32'hc0a12cf4} /* (3, 18, 1) {real, imag} */,
  {32'h3fbc0a6c, 32'hc01c9cea} /* (3, 18, 0) {real, imag} */,
  {32'h3f23b8bc, 32'hc0dd3ca5} /* (3, 17, 31) {real, imag} */,
  {32'h4018d5e6, 32'hc11ccde4} /* (3, 17, 30) {real, imag} */,
  {32'h400efc42, 32'hc0c2cf16} /* (3, 17, 29) {real, imag} */,
  {32'h3f205307, 32'hc0bb637f} /* (3, 17, 28) {real, imag} */,
  {32'h3fa5de4f, 32'hc0a774ca} /* (3, 17, 27) {real, imag} */,
  {32'h3f6715d2, 32'hc09de2e4} /* (3, 17, 26) {real, imag} */,
  {32'h4087c0a6, 32'hc0b9c3a2} /* (3, 17, 25) {real, imag} */,
  {32'h4009c262, 32'hc0cf8898} /* (3, 17, 24) {real, imag} */,
  {32'h4018cc7c, 32'hc0b83e3c} /* (3, 17, 23) {real, imag} */,
  {32'h3fab1069, 32'hc070b69e} /* (3, 17, 22) {real, imag} */,
  {32'hbf53dc68, 32'hc01b20cb} /* (3, 17, 21) {real, imag} */,
  {32'h3fd670fe, 32'h40a16e69} /* (3, 17, 20) {real, imag} */,
  {32'hbfb10ae3, 32'h407d69be} /* (3, 17, 19) {real, imag} */,
  {32'hc090db56, 32'h4092231a} /* (3, 17, 18) {real, imag} */,
  {32'hc09dcecf, 32'h40eeddca} /* (3, 17, 17) {real, imag} */,
  {32'hc040d146, 32'h406d50ce} /* (3, 17, 16) {real, imag} */,
  {32'hbffbc713, 32'h40a52148} /* (3, 17, 15) {real, imag} */,
  {32'hbfa54d35, 32'h4105e5c0} /* (3, 17, 14) {real, imag} */,
  {32'hbecb3b8c, 32'h40dcba60} /* (3, 17, 13) {real, imag} */,
  {32'hbfab47ac, 32'h4094aec1} /* (3, 17, 12) {real, imag} */,
  {32'hbf973e32, 32'h409df11e} /* (3, 17, 11) {real, imag} */,
  {32'hc065c9da, 32'h3e482854} /* (3, 17, 10) {real, imag} */,
  {32'hbf9ad68e, 32'hc08ed0d2} /* (3, 17, 9) {real, imag} */,
  {32'hbfa47677, 32'hc098691e} /* (3, 17, 8) {real, imag} */,
  {32'h3e1e1b8e, 32'hc0aabaee} /* (3, 17, 7) {real, imag} */,
  {32'h403a25b4, 32'hc0bce1b4} /* (3, 17, 6) {real, imag} */,
  {32'h4035454b, 32'hc03ba606} /* (3, 17, 5) {real, imag} */,
  {32'h3ed19a60, 32'hc06b00d3} /* (3, 17, 4) {real, imag} */,
  {32'hc004a79a, 32'hc0ded42d} /* (3, 17, 3) {real, imag} */,
  {32'h3f034cf4, 32'hc0b4cff5} /* (3, 17, 2) {real, imag} */,
  {32'h4029dc37, 32'hc066eef5} /* (3, 17, 1) {real, imag} */,
  {32'h3f737831, 32'hc02d1a14} /* (3, 17, 0) {real, imag} */,
  {32'h3f867462, 32'hc08ab702} /* (3, 16, 31) {real, imag} */,
  {32'h403a6aaa, 32'hc115bd52} /* (3, 16, 30) {real, imag} */,
  {32'h40054f77, 32'hc0bd5767} /* (3, 16, 29) {real, imag} */,
  {32'hbea2741c, 32'hc0936682} /* (3, 16, 28) {real, imag} */,
  {32'h3fac9137, 32'hbfdf44e5} /* (3, 16, 27) {real, imag} */,
  {32'h3ff72225, 32'hbf899d8e} /* (3, 16, 26) {real, imag} */,
  {32'h409205e2, 32'hc09d0b40} /* (3, 16, 25) {real, imag} */,
  {32'h3f937ac8, 32'hc09148c0} /* (3, 16, 24) {real, imag} */,
  {32'h3f3524fd, 32'hc0a45d7a} /* (3, 16, 23) {real, imag} */,
  {32'h405848dc, 32'hc09180de} /* (3, 16, 22) {real, imag} */,
  {32'h3f22b54b, 32'hc00f2258} /* (3, 16, 21) {real, imag} */,
  {32'hbfe44120, 32'h4065ae04} /* (3, 16, 20) {real, imag} */,
  {32'hbfd5a360, 32'h408e5d4e} /* (3, 16, 19) {real, imag} */,
  {32'hc0262495, 32'h4073c0de} /* (3, 16, 18) {real, imag} */,
  {32'hbfd949e2, 32'h409d6b12} /* (3, 16, 17) {real, imag} */,
  {32'h3f9445f9, 32'h40cdf196} /* (3, 16, 16) {real, imag} */,
  {32'hbf3a1ce7, 32'h40d7c7d4} /* (3, 16, 15) {real, imag} */,
  {32'hbf1bc8ed, 32'h40971f26} /* (3, 16, 14) {real, imag} */,
  {32'h3eafc692, 32'h40867266} /* (3, 16, 13) {real, imag} */,
  {32'h3f1fb225, 32'h407466fc} /* (3, 16, 12) {real, imag} */,
  {32'hc010419e, 32'h4023c8fe} /* (3, 16, 11) {real, imag} */,
  {32'hc0851f68, 32'hbfe31309} /* (3, 16, 10) {real, imag} */,
  {32'h3f310be0, 32'hc07ad4d4} /* (3, 16, 9) {real, imag} */,
  {32'h3efd83c0, 32'hc08d90f8} /* (3, 16, 8) {real, imag} */,
  {32'h3fa0dcd4, 32'hc0b1420c} /* (3, 16, 7) {real, imag} */,
  {32'h40283e8a, 32'hc0fad32e} /* (3, 16, 6) {real, imag} */,
  {32'h40310a9e, 32'hc0a9f578} /* (3, 16, 5) {real, imag} */,
  {32'h3fe3ec54, 32'hc0c672f0} /* (3, 16, 4) {real, imag} */,
  {32'hbe65b428, 32'hc0f6739c} /* (3, 16, 3) {real, imag} */,
  {32'h3fc85017, 32'hc10c1f8e} /* (3, 16, 2) {real, imag} */,
  {32'h4054b614, 32'hc0f1116c} /* (3, 16, 1) {real, imag} */,
  {32'h3f0da093, 32'hc091a7f6} /* (3, 16, 0) {real, imag} */,
  {32'h3ffd5b98, 32'hc0512254} /* (3, 15, 31) {real, imag} */,
  {32'h4053879f, 32'hc0d9da49} /* (3, 15, 30) {real, imag} */,
  {32'h403429b9, 32'hc09a8462} /* (3, 15, 29) {real, imag} */,
  {32'h3f89f639, 32'hc087800c} /* (3, 15, 28) {real, imag} */,
  {32'h3fe34a12, 32'hc046ae4e} /* (3, 15, 27) {real, imag} */,
  {32'h40782f17, 32'hbfbc108f} /* (3, 15, 26) {real, imag} */,
  {32'h40d85be7, 32'hc05e2ae5} /* (3, 15, 25) {real, imag} */,
  {32'h3fe49ae6, 32'hc0831c69} /* (3, 15, 24) {real, imag} */,
  {32'h3f01eb9c, 32'hc05b6949} /* (3, 15, 23) {real, imag} */,
  {32'h40682d4d, 32'hc02d6a8c} /* (3, 15, 22) {real, imag} */,
  {32'h3f903327, 32'h3fc05654} /* (3, 15, 21) {real, imag} */,
  {32'hc07b5097, 32'h40c6ea7a} /* (3, 15, 20) {real, imag} */,
  {32'hc04ad2e3, 32'h403569af} /* (3, 15, 19) {real, imag} */,
  {32'hbf1ec740, 32'h40285b5a} /* (3, 15, 18) {real, imag} */,
  {32'hbd6c36c8, 32'h407f7248} /* (3, 15, 17) {real, imag} */,
  {32'hc01b681c, 32'h40be5368} /* (3, 15, 16) {real, imag} */,
  {32'hbf58e613, 32'h409eb10e} /* (3, 15, 15) {real, imag} */,
  {32'h3e1409bd, 32'h408ca6c8} /* (3, 15, 14) {real, imag} */,
  {32'hbf972830, 32'h40c6f1f6} /* (3, 15, 13) {real, imag} */,
  {32'hc031d010, 32'h40ae6c77} /* (3, 15, 12) {real, imag} */,
  {32'hc0a0834c, 32'h3e96af30} /* (3, 15, 11) {real, imag} */,
  {32'hc07b16ec, 32'hc045a54f} /* (3, 15, 10) {real, imag} */,
  {32'hbfb063fc, 32'hc088f22e} /* (3, 15, 9) {real, imag} */,
  {32'h3ed26e10, 32'hc0a3acb9} /* (3, 15, 8) {real, imag} */,
  {32'h40046604, 32'hc0b309f0} /* (3, 15, 7) {real, imag} */,
  {32'h402e2f1c, 32'hc04ae68d} /* (3, 15, 6) {real, imag} */,
  {32'h4086028c, 32'hc07f4f0c} /* (3, 15, 5) {real, imag} */,
  {32'h403d3ff0, 32'hc0a4d9c7} /* (3, 15, 4) {real, imag} */,
  {32'h4072c38b, 32'hc0ba0a7a} /* (3, 15, 3) {real, imag} */,
  {32'h4095257e, 32'hc0cdc506} /* (3, 15, 2) {real, imag} */,
  {32'h40355430, 32'hc09fb21c} /* (3, 15, 1) {real, imag} */,
  {32'hbef22ba7, 32'hbfd0d544} /* (3, 15, 0) {real, imag} */,
  {32'h3f9f7290, 32'hc090d176} /* (3, 14, 31) {real, imag} */,
  {32'h405509f2, 32'hc0c66895} /* (3, 14, 30) {real, imag} */,
  {32'h407dc35e, 32'hc04adb77} /* (3, 14, 29) {real, imag} */,
  {32'h40666b09, 32'hc03dd1c0} /* (3, 14, 28) {real, imag} */,
  {32'h400ce2e8, 32'hc08d2511} /* (3, 14, 27) {real, imag} */,
  {32'h408352d6, 32'hc0954fb2} /* (3, 14, 26) {real, imag} */,
  {32'h40f1dd86, 32'hc0a873a0} /* (3, 14, 25) {real, imag} */,
  {32'h40c94e50, 32'hc0bb5326} /* (3, 14, 24) {real, imag} */,
  {32'h40a6b5d2, 32'hc0d9b15c} /* (3, 14, 23) {real, imag} */,
  {32'h404de288, 32'hc0b40ca1} /* (3, 14, 22) {real, imag} */,
  {32'hbf837c8a, 32'hbf2d7c33} /* (3, 14, 21) {real, imag} */,
  {32'hbffd3d83, 32'h408772d3} /* (3, 14, 20) {real, imag} */,
  {32'hbef01cf8, 32'h4029f946} /* (3, 14, 19) {real, imag} */,
  {32'hbfc81883, 32'h40545dd8} /* (3, 14, 18) {real, imag} */,
  {32'hc0044bc1, 32'h40948ca6} /* (3, 14, 17) {real, imag} */,
  {32'hc03aad95, 32'h40b0ed78} /* (3, 14, 16) {real, imag} */,
  {32'hbff89288, 32'h403c1138} /* (3, 14, 15) {real, imag} */,
  {32'hbe5114d8, 32'h40215408} /* (3, 14, 14) {real, imag} */,
  {32'hbff51b5a, 32'h40c272ac} /* (3, 14, 13) {real, imag} */,
  {32'hc04d93ce, 32'h409e2144} /* (3, 14, 12) {real, imag} */,
  {32'hc03da8fc, 32'h4036ea74} /* (3, 14, 11) {real, imag} */,
  {32'h3f228186, 32'hc0448403} /* (3, 14, 10) {real, imag} */,
  {32'h3fbafa33, 32'hc1077e24} /* (3, 14, 9) {real, imag} */,
  {32'h3ff979b3, 32'hc115c190} /* (3, 14, 8) {real, imag} */,
  {32'h4045b407, 32'hc0c0f325} /* (3, 14, 7) {real, imag} */,
  {32'h3fe75410, 32'hc00b64b0} /* (3, 14, 6) {real, imag} */,
  {32'h40579a54, 32'hc0d08ba2} /* (3, 14, 5) {real, imag} */,
  {32'h402adbeb, 32'hc0a3cefa} /* (3, 14, 4) {real, imag} */,
  {32'h404834b8, 32'hc0bbbc88} /* (3, 14, 3) {real, imag} */,
  {32'h40a160dc, 32'hc0476944} /* (3, 14, 2) {real, imag} */,
  {32'h401ebbd1, 32'hc0037266} /* (3, 14, 1) {real, imag} */,
  {32'hbfa57640, 32'hbfe3618e} /* (3, 14, 0) {real, imag} */,
  {32'h3edbefe3, 32'hc0876fb1} /* (3, 13, 31) {real, imag} */,
  {32'h400420c8, 32'hc09099a0} /* (3, 13, 30) {real, imag} */,
  {32'h405acdb6, 32'hc0c1ac32} /* (3, 13, 29) {real, imag} */,
  {32'h3fc2a08e, 32'hc0dbb699} /* (3, 13, 28) {real, imag} */,
  {32'h40080788, 32'hc0be333f} /* (3, 13, 27) {real, imag} */,
  {32'h401cacaa, 32'hc0d83d82} /* (3, 13, 26) {real, imag} */,
  {32'h40287188, 32'hc0d7d249} /* (3, 13, 25) {real, imag} */,
  {32'h406bea3c, 32'hc1015b30} /* (3, 13, 24) {real, imag} */,
  {32'h40466922, 32'hc10dd926} /* (3, 13, 23) {real, imag} */,
  {32'h402c9498, 32'hc0fbd961} /* (3, 13, 22) {real, imag} */,
  {32'hbc2dc600, 32'hbfd4f1d0} /* (3, 13, 21) {real, imag} */,
  {32'hbf29f668, 32'h40af83a0} /* (3, 13, 20) {real, imag} */,
  {32'hbf922a1a, 32'h40c585f0} /* (3, 13, 19) {real, imag} */,
  {32'hc0157600, 32'h40b45812} /* (3, 13, 18) {real, imag} */,
  {32'hbfd7c7bf, 32'h40c697bd} /* (3, 13, 17) {real, imag} */,
  {32'hbfbe94be, 32'h40de6bec} /* (3, 13, 16) {real, imag} */,
  {32'h3f240703, 32'h4058f851} /* (3, 13, 15) {real, imag} */,
  {32'h3f11ba20, 32'h3f137f9d} /* (3, 13, 14) {real, imag} */,
  {32'hc01a585d, 32'h40683492} /* (3, 13, 13) {real, imag} */,
  {32'hc068471e, 32'h40bee69a} /* (3, 13, 12) {real, imag} */,
  {32'hc066d065, 32'h40af6c56} /* (3, 13, 11) {real, imag} */,
  {32'h3f45b14a, 32'hc082dc9e} /* (3, 13, 10) {real, imag} */,
  {32'h408c1990, 32'hc117753c} /* (3, 13, 9) {real, imag} */,
  {32'h403be916, 32'hc0edbbef} /* (3, 13, 8) {real, imag} */,
  {32'h4077300d, 32'hc0882d2a} /* (3, 13, 7) {real, imag} */,
  {32'h3fb579c3, 32'hc09dfbeb} /* (3, 13, 6) {real, imag} */,
  {32'h3fc5d83c, 32'hc1113100} /* (3, 13, 5) {real, imag} */,
  {32'h3f9b1a28, 32'hc0cf0daa} /* (3, 13, 4) {real, imag} */,
  {32'h3f8822e8, 32'hc0be0823} /* (3, 13, 3) {real, imag} */,
  {32'h3fdac35f, 32'hc067182c} /* (3, 13, 2) {real, imag} */,
  {32'h3fa6fc35, 32'hc09d2ca0} /* (3, 13, 1) {real, imag} */,
  {32'hbe8b88a5, 32'hc07c1950} /* (3, 13, 0) {real, imag} */,
  {32'hbf32d99e, 32'hbfe255f2} /* (3, 12, 31) {real, imag} */,
  {32'hbee9fcc4, 32'hc05ab1ec} /* (3, 12, 30) {real, imag} */,
  {32'hbf0c2ace, 32'hc092950a} /* (3, 12, 29) {real, imag} */,
  {32'h3fb1c7b8, 32'hc11152c4} /* (3, 12, 28) {real, imag} */,
  {32'h4023d1b8, 32'hc11df772} /* (3, 12, 27) {real, imag} */,
  {32'h40209c82, 32'hc0f2567e} /* (3, 12, 26) {real, imag} */,
  {32'h3fe97ef0, 32'hc104d0b4} /* (3, 12, 25) {real, imag} */,
  {32'h3fb27715, 32'hc11d57c4} /* (3, 12, 24) {real, imag} */,
  {32'h402310bf, 32'hc0d53659} /* (3, 12, 23) {real, imag} */,
  {32'h402978c8, 32'hc08e8612} /* (3, 12, 22) {real, imag} */,
  {32'hbf9b3170, 32'hbec10af2} /* (3, 12, 21) {real, imag} */,
  {32'hbfb8051a, 32'h40b65841} /* (3, 12, 20) {real, imag} */,
  {32'h3f58ec9d, 32'h40d3eba4} /* (3, 12, 19) {real, imag} */,
  {32'hc004d0b0, 32'h40cb7691} /* (3, 12, 18) {real, imag} */,
  {32'hc059442a, 32'h40b8fb3a} /* (3, 12, 17) {real, imag} */,
  {32'h3f9113ad, 32'h40bc1d0a} /* (3, 12, 16) {real, imag} */,
  {32'h404174d0, 32'h4087defc} /* (3, 12, 15) {real, imag} */,
  {32'hbc4aa870, 32'h4005bb47} /* (3, 12, 14) {real, imag} */,
  {32'hc089a2c7, 32'h3fe0bfd4} /* (3, 12, 13) {real, imag} */,
  {32'hc08b59fb, 32'h408b6f4d} /* (3, 12, 12) {real, imag} */,
  {32'hc0991358, 32'h408e0b2d} /* (3, 12, 11) {real, imag} */,
  {32'hbfd67e20, 32'hc0657e66} /* (3, 12, 10) {real, imag} */,
  {32'h3f81e89e, 32'hc0d4d477} /* (3, 12, 9) {real, imag} */,
  {32'h4034f774, 32'hc0a783b8} /* (3, 12, 8) {real, imag} */,
  {32'h40000254, 32'hc0923f3e} /* (3, 12, 7) {real, imag} */,
  {32'h3e99dbd6, 32'hc0f68f40} /* (3, 12, 6) {real, imag} */,
  {32'h3fa212c5, 32'hc0ecbb74} /* (3, 12, 5) {real, imag} */,
  {32'h3eea2ed6, 32'hc0b33296} /* (3, 12, 4) {real, imag} */,
  {32'h3ed54984, 32'hc09f2878} /* (3, 12, 3) {real, imag} */,
  {32'h3ee0f9ce, 32'hc0d61b4e} /* (3, 12, 2) {real, imag} */,
  {32'h3f644a5a, 32'hc1185e24} /* (3, 12, 1) {real, imag} */,
  {32'hbf73334f, 32'hc0bd00b7} /* (3, 12, 0) {real, imag} */,
  {32'hbf6a6f29, 32'hc0108b0c} /* (3, 11, 31) {real, imag} */,
  {32'hbfe96428, 32'hc068be15} /* (3, 11, 30) {real, imag} */,
  {32'h3febc604, 32'hc04435de} /* (3, 11, 29) {real, imag} */,
  {32'h400fe54e, 32'hc0b4d082} /* (3, 11, 28) {real, imag} */,
  {32'h40027764, 32'hc10884a3} /* (3, 11, 27) {real, imag} */,
  {32'h40673494, 32'hc0a9eae0} /* (3, 11, 26) {real, imag} */,
  {32'h401341cc, 32'hc0cb0d6e} /* (3, 11, 25) {real, imag} */,
  {32'h3f647fba, 32'hc0e21f3e} /* (3, 11, 24) {real, imag} */,
  {32'h3f9656d0, 32'hc028dc46} /* (3, 11, 23) {real, imag} */,
  {32'hbe167e58, 32'hc08bda4e} /* (3, 11, 22) {real, imag} */,
  {32'hc075dbbc, 32'hbfcf5fae} /* (3, 11, 21) {real, imag} */,
  {32'hc03a36e6, 32'h401add60} /* (3, 11, 20) {real, imag} */,
  {32'h4015a686, 32'h409e6aaa} /* (3, 11, 19) {real, imag} */,
  {32'h3d8e005c, 32'h409ff11f} /* (3, 11, 18) {real, imag} */,
  {32'hc024f3f2, 32'h403b8694} /* (3, 11, 17) {real, imag} */,
  {32'h3fcfe389, 32'h4070609c} /* (3, 11, 16) {real, imag} */,
  {32'h3f17e0c0, 32'h40a99bb1} /* (3, 11, 15) {real, imag} */,
  {32'hbf7b1dca, 32'h40834a47} /* (3, 11, 14) {real, imag} */,
  {32'hbf960516, 32'h408ad824} /* (3, 11, 13) {real, imag} */,
  {32'hbfe36012, 32'h408d834c} /* (3, 11, 12) {real, imag} */,
  {32'hbfe11412, 32'h4084e4fb} /* (3, 11, 11) {real, imag} */,
  {32'h3f302583, 32'hbf849ffe} /* (3, 11, 10) {real, imag} */,
  {32'h3eb94eaa, 32'hc0a1d45c} /* (3, 11, 9) {real, imag} */,
  {32'h3fa1c922, 32'hc0b0ad3c} /* (3, 11, 8) {real, imag} */,
  {32'h3fec4ec9, 32'hc0ce01c0} /* (3, 11, 7) {real, imag} */,
  {32'h3fee3e2e, 32'hc0b24c0e} /* (3, 11, 6) {real, imag} */,
  {32'h3f844d8c, 32'hc08c349f} /* (3, 11, 5) {real, imag} */,
  {32'hbb88c780, 32'hc02e830c} /* (3, 11, 4) {real, imag} */,
  {32'hbe21961a, 32'hc076c964} /* (3, 11, 3) {real, imag} */,
  {32'h3f24382e, 32'hc0b254fa} /* (3, 11, 2) {real, imag} */,
  {32'hbf5a3840, 32'hc0c288c8} /* (3, 11, 1) {real, imag} */,
  {32'hbf9e2e9a, 32'hc07169c9} /* (3, 11, 0) {real, imag} */,
  {32'hbc2bdfa0, 32'h3f3b55de} /* (3, 10, 31) {real, imag} */,
  {32'hbf99d21c, 32'h3f1f6742} /* (3, 10, 30) {real, imag} */,
  {32'h3f659762, 32'hbecdc93a} /* (3, 10, 29) {real, imag} */,
  {32'h3d9f3718, 32'hbd790510} /* (3, 10, 28) {real, imag} */,
  {32'hbfa3401a, 32'h3fa1f6b8} /* (3, 10, 27) {real, imag} */,
  {32'h3ea206a0, 32'h3f9f3838} /* (3, 10, 26) {real, imag} */,
  {32'h3fd91645, 32'h3ff8286a} /* (3, 10, 25) {real, imag} */,
  {32'h3d98a490, 32'h3f422630} /* (3, 10, 24) {real, imag} */,
  {32'hbfb7cd60, 32'h409da647} /* (3, 10, 23) {real, imag} */,
  {32'hc04c8029, 32'h4031bc1c} /* (3, 10, 22) {real, imag} */,
  {32'hbf34a51c, 32'h40493dc7} /* (3, 10, 21) {real, imag} */,
  {32'h3feb2830, 32'hbf665a07} /* (3, 10, 20) {real, imag} */,
  {32'h3ff4f516, 32'hc02ba6a8} /* (3, 10, 19) {real, imag} */,
  {32'h3f6b7a73, 32'hbfe84883} /* (3, 10, 18) {real, imag} */,
  {32'h40249b7e, 32'hc0b567d8} /* (3, 10, 17) {real, imag} */,
  {32'h3f6dbafe, 32'hc07e26ee} /* (3, 10, 16) {real, imag} */,
  {32'hc0332004, 32'hbf6fd99e} /* (3, 10, 15) {real, imag} */,
  {32'hbf17b9fe, 32'hbf8fc9f6} /* (3, 10, 14) {real, imag} */,
  {32'hbd47c7ba, 32'hbed1f63a} /* (3, 10, 13) {real, imag} */,
  {32'h3f281464, 32'hc00cf29c} /* (3, 10, 12) {real, imag} */,
  {32'h3faa88af, 32'hbfdb9ae4} /* (3, 10, 11) {real, imag} */,
  {32'h3f985f19, 32'h3ecb7a4a} /* (3, 10, 10) {real, imag} */,
  {32'hbefd1332, 32'hba4f3a00} /* (3, 10, 9) {real, imag} */,
  {32'hbe9487d7, 32'h3faf55b8} /* (3, 10, 8) {real, imag} */,
  {32'h3f8f5f50, 32'h3fce7413} /* (3, 10, 7) {real, imag} */,
  {32'h3f4fd752, 32'h4016b3d7} /* (3, 10, 6) {real, imag} */,
  {32'h3e77de34, 32'h3f3a61df} /* (3, 10, 5) {real, imag} */,
  {32'h3f0889c4, 32'h40728d2b} /* (3, 10, 4) {real, imag} */,
  {32'hc000fbe4, 32'h408a31dd} /* (3, 10, 3) {real, imag} */,
  {32'hc000e00a, 32'h3f68e017} /* (3, 10, 2) {real, imag} */,
  {32'hbfffa6d4, 32'h3fadb452} /* (3, 10, 1) {real, imag} */,
  {32'hbf89ed43, 32'h3ffde762} /* (3, 10, 0) {real, imag} */,
  {32'hbff440fc, 32'h40c3e124} /* (3, 9, 31) {real, imag} */,
  {32'hc02c520c, 32'h40fa84b4} /* (3, 9, 30) {real, imag} */,
  {32'hbff92a26, 32'h40d72a14} /* (3, 9, 29) {real, imag} */,
  {32'hbe9ee5bb, 32'h4062f9fc} /* (3, 9, 28) {real, imag} */,
  {32'hbdb78ff0, 32'h40948044} /* (3, 9, 27) {real, imag} */,
  {32'hbfcbc558, 32'h406c311e} /* (3, 9, 26) {real, imag} */,
  {32'hbf9fbe38, 32'h40a70491} /* (3, 9, 25) {real, imag} */,
  {32'hbfd97819, 32'h409a169e} /* (3, 9, 24) {real, imag} */,
  {32'hc052be3c, 32'h40e9939a} /* (3, 9, 23) {real, imag} */,
  {32'hc0982956, 32'h40e4591c} /* (3, 9, 22) {real, imag} */,
  {32'hc054bf7a, 32'h4073b006} /* (3, 9, 21) {real, imag} */,
  {32'h40263b42, 32'hbfb10eee} /* (3, 9, 20) {real, imag} */,
  {32'h4020c176, 32'hc0acbec9} /* (3, 9, 19) {real, imag} */,
  {32'h3f2bf702, 32'hc06eee5c} /* (3, 9, 18) {real, imag} */,
  {32'h3fb3d29b, 32'hc0ac6642} /* (3, 9, 17) {real, imag} */,
  {32'hbfdc5136, 32'hc0baeff1} /* (3, 9, 16) {real, imag} */,
  {32'hbf6916b7, 32'hc05c072c} /* (3, 9, 15) {real, imag} */,
  {32'h3dde2a98, 32'hc019cb29} /* (3, 9, 14) {real, imag} */,
  {32'h3fa968eb, 32'hc0b20b45} /* (3, 9, 13) {real, imag} */,
  {32'h3f8b22d8, 32'hc111f0a3} /* (3, 9, 12) {real, imag} */,
  {32'h3fca34d3, 32'hc0c1be30} /* (3, 9, 11) {real, imag} */,
  {32'hbc7d7120, 32'hbf3e4c40} /* (3, 9, 10) {real, imag} */,
  {32'hbf88d5cd, 32'h3fcf2878} /* (3, 9, 9) {real, imag} */,
  {32'hbed039b2, 32'h4098be91} /* (3, 9, 8) {real, imag} */,
  {32'hbfffab2e, 32'h40b014b3} /* (3, 9, 7) {real, imag} */,
  {32'hc045ba3e, 32'h405ee25b} /* (3, 9, 6) {real, imag} */,
  {32'h3d5379b0, 32'h403a723e} /* (3, 9, 5) {real, imag} */,
  {32'hc000ab3a, 32'h40982774} /* (3, 9, 4) {real, imag} */,
  {32'hc074b346, 32'h41140d3c} /* (3, 9, 3) {real, imag} */,
  {32'hc07476fc, 32'h40e1d47a} /* (3, 9, 2) {real, imag} */,
  {32'hc03d1121, 32'h408ad423} /* (3, 9, 1) {real, imag} */,
  {32'hbfc6a05a, 32'h4039aa2e} /* (3, 9, 0) {real, imag} */,
  {32'hc00cfa62, 32'h4070dd73} /* (3, 8, 31) {real, imag} */,
  {32'hc07d1817, 32'h40ae174c} /* (3, 8, 30) {real, imag} */,
  {32'hc013257e, 32'h40f660cd} /* (3, 8, 29) {real, imag} */,
  {32'h3fb26afc, 32'h4063ae25} /* (3, 8, 28) {real, imag} */,
  {32'h402d0d2f, 32'h408bf33d} /* (3, 8, 27) {real, imag} */,
  {32'h3f6bba6c, 32'h40b8fca5} /* (3, 8, 26) {real, imag} */,
  {32'h3edb7348, 32'h40aa2508} /* (3, 8, 25) {real, imag} */,
  {32'hbff4da6e, 32'h40ab0901} /* (3, 8, 24) {real, imag} */,
  {32'hc05f3722, 32'h40da8135} /* (3, 8, 23) {real, imag} */,
  {32'hc0d29a70, 32'h40d7c1f0} /* (3, 8, 22) {real, imag} */,
  {32'hc08f07f1, 32'h3f4bf242} /* (3, 8, 21) {real, imag} */,
  {32'h3f8796d0, 32'hc060a864} /* (3, 8, 20) {real, imag} */,
  {32'h401818dc, 32'hc0a73a4d} /* (3, 8, 19) {real, imag} */,
  {32'h3fc1f52f, 32'hc0d14b4a} /* (3, 8, 18) {real, imag} */,
  {32'h3f1d9ad5, 32'hc0dd9599} /* (3, 8, 17) {real, imag} */,
  {32'hbf5a2850, 32'hc0a3907f} /* (3, 8, 16) {real, imag} */,
  {32'h3fd2bfea, 32'hc05b163a} /* (3, 8, 15) {real, imag} */,
  {32'h40673d3c, 32'hc091902e} /* (3, 8, 14) {real, imag} */,
  {32'h406b34ea, 32'hc0ced7f1} /* (3, 8, 13) {real, imag} */,
  {32'h3f54558e, 32'hc1136d05} /* (3, 8, 12) {real, imag} */,
  {32'h400c33f2, 32'hc0a53e11} /* (3, 8, 11) {real, imag} */,
  {32'h3f5c07df, 32'h3f4e6fd5} /* (3, 8, 10) {real, imag} */,
  {32'hbee8655a, 32'h40695e66} /* (3, 8, 9) {real, imag} */,
  {32'hbf7a45da, 32'h40d68e46} /* (3, 8, 8) {real, imag} */,
  {32'hbfffd0b7, 32'h40cfddfb} /* (3, 8, 7) {real, imag} */,
  {32'hc0075820, 32'h40868211} /* (3, 8, 6) {real, imag} */,
  {32'h3f908306, 32'h40421943} /* (3, 8, 5) {real, imag} */,
  {32'hbf16025d, 32'h40bf037e} /* (3, 8, 4) {real, imag} */,
  {32'hc0631b0a, 32'h40eb0f26} /* (3, 8, 3) {real, imag} */,
  {32'hc073c2ac, 32'h40c3a29c} /* (3, 8, 2) {real, imag} */,
  {32'hbf8cc938, 32'h40b15390} /* (3, 8, 1) {real, imag} */,
  {32'h3fe1591e, 32'h401d5970} /* (3, 8, 0) {real, imag} */,
  {32'hbfaba2e2, 32'h3f69882e} /* (3, 7, 31) {real, imag} */,
  {32'hc04d5930, 32'h40542640} /* (3, 7, 30) {real, imag} */,
  {32'hbd5a4c30, 32'h40e37dee} /* (3, 7, 29) {real, imag} */,
  {32'h3fc1f19e, 32'h40edf586} /* (3, 7, 28) {real, imag} */,
  {32'h3f88de0a, 32'h40c5563a} /* (3, 7, 27) {real, imag} */,
  {32'hbfab0d0d, 32'h40baa85e} /* (3, 7, 26) {real, imag} */,
  {32'hbff2fc19, 32'h40a77a79} /* (3, 7, 25) {real, imag} */,
  {32'hc0202a42, 32'h40d3a3b4} /* (3, 7, 24) {real, imag} */,
  {32'hc06105cf, 32'h40c4c2d3} /* (3, 7, 23) {real, imag} */,
  {32'hc082652c, 32'h405dabe0} /* (3, 7, 22) {real, imag} */,
  {32'hbf835650, 32'hc0033ec8} /* (3, 7, 21) {real, imag} */,
  {32'h40133d5e, 32'hc0c6712a} /* (3, 7, 20) {real, imag} */,
  {32'h40569c8b, 32'hc085c39d} /* (3, 7, 19) {real, imag} */,
  {32'h3e3b9408, 32'hc06831b7} /* (3, 7, 18) {real, imag} */,
  {32'h3f8e0a0c, 32'hc0e3dacf} /* (3, 7, 17) {real, imag} */,
  {32'h4007f3c7, 32'hc0d002a6} /* (3, 7, 16) {real, imag} */,
  {32'h4073cc74, 32'hc09964ca} /* (3, 7, 15) {real, imag} */,
  {32'h40941af9, 32'hc0c38676} /* (3, 7, 14) {real, imag} */,
  {32'h40778623, 32'hc0b76cf3} /* (3, 7, 13) {real, imag} */,
  {32'hbf8466d0, 32'hc089e83e} /* (3, 7, 12) {real, imag} */,
  {32'hc06bec38, 32'hc023e113} /* (3, 7, 11) {real, imag} */,
  {32'hbea46b22, 32'h40187458} /* (3, 7, 10) {real, imag} */,
  {32'h3dfcb200, 32'h40c6ebc5} /* (3, 7, 9) {real, imag} */,
  {32'hbf882ca8, 32'h40d3f2bc} /* (3, 7, 8) {real, imag} */,
  {32'h3f94fad5, 32'h4057a684} /* (3, 7, 7) {real, imag} */,
  {32'h3f2a977a, 32'h4050ea5c} /* (3, 7, 6) {real, imag} */,
  {32'hc01f2868, 32'h40b8b79b} /* (3, 7, 5) {real, imag} */,
  {32'hbe46bb9c, 32'h40db7c7c} /* (3, 7, 4) {real, imag} */,
  {32'hbfca062b, 32'h41017026} /* (3, 7, 3) {real, imag} */,
  {32'hc0a02c1c, 32'h40ed7df0} /* (3, 7, 2) {real, imag} */,
  {32'hc002561e, 32'h40c000c6} /* (3, 7, 1) {real, imag} */,
  {32'hbd0e6618, 32'h4012529f} /* (3, 7, 0) {real, imag} */,
  {32'hbef0f380, 32'h400f07b8} /* (3, 6, 31) {real, imag} */,
  {32'hbf9b25d2, 32'h40774eed} /* (3, 6, 30) {real, imag} */,
  {32'h3fc5750e, 32'h40ea971d} /* (3, 6, 29) {real, imag} */,
  {32'h3eb3c5be, 32'h40fb6f46} /* (3, 6, 28) {real, imag} */,
  {32'hc07f6577, 32'h40bace02} /* (3, 6, 27) {real, imag} */,
  {32'hc08df2e4, 32'h40b4c673} /* (3, 6, 26) {real, imag} */,
  {32'hc04cefbe, 32'h408fc8b8} /* (3, 6, 25) {real, imag} */,
  {32'hbf557ffc, 32'h40c36dce} /* (3, 6, 24) {real, imag} */,
  {32'hbfd74202, 32'h40b2bf3e} /* (3, 6, 23) {real, imag} */,
  {32'hc08f804c, 32'h4056d0ac} /* (3, 6, 22) {real, imag} */,
  {32'hbf866d14, 32'h3f147aa4} /* (3, 6, 21) {real, imag} */,
  {32'h40869b38, 32'hc05cce8a} /* (3, 6, 20) {real, imag} */,
  {32'h4059c510, 32'hc00baec0} /* (3, 6, 19) {real, imag} */,
  {32'h3d82735c, 32'hc00255b0} /* (3, 6, 18) {real, imag} */,
  {32'hbe4cfbca, 32'hc090f409} /* (3, 6, 17) {real, imag} */,
  {32'h3e3440cc, 32'hc0baa8c4} /* (3, 6, 16) {real, imag} */,
  {32'h405aef0d, 32'hc0c06559} /* (3, 6, 15) {real, imag} */,
  {32'h3ff8891c, 32'hc0c83b19} /* (3, 6, 14) {real, imag} */,
  {32'h4032b8b0, 32'hc0c17014} /* (3, 6, 13) {real, imag} */,
  {32'h3fb5728b, 32'hc0c10400} /* (3, 6, 12) {real, imag} */,
  {32'hbfec3f0a, 32'hc0b479fd} /* (3, 6, 11) {real, imag} */,
  {32'hc05f5166, 32'h400b3b53} /* (3, 6, 10) {real, imag} */,
  {32'hc0906dd6, 32'h40980e14} /* (3, 6, 9) {real, imag} */,
  {32'hc06319a8, 32'h4047457e} /* (3, 6, 8) {real, imag} */,
  {32'h3fbdae13, 32'h40876fde} /* (3, 6, 7) {real, imag} */,
  {32'hbde35a54, 32'h40bc6bbe} /* (3, 6, 6) {real, imag} */,
  {32'hc08d0c1a, 32'h40f2c7eb} /* (3, 6, 5) {real, imag} */,
  {32'hc0156b48, 32'h4089875f} /* (3, 6, 4) {real, imag} */,
  {32'h3ed983fa, 32'h4075f7c9} /* (3, 6, 3) {real, imag} */,
  {32'h3c72d580, 32'h40b81c46} /* (3, 6, 2) {real, imag} */,
  {32'h3f74b34c, 32'h40b88e2e} /* (3, 6, 1) {real, imag} */,
  {32'hbe84322a, 32'h405abd48} /* (3, 6, 0) {real, imag} */,
  {32'hc0409ec8, 32'h4088cc55} /* (3, 5, 31) {real, imag} */,
  {32'hc05025d5, 32'h406b08ca} /* (3, 5, 30) {real, imag} */,
  {32'hbe390230, 32'h40a100d2} /* (3, 5, 29) {real, imag} */,
  {32'hbfa04f53, 32'h40f0e0fc} /* (3, 5, 28) {real, imag} */,
  {32'hc05492cc, 32'h40cc4bfe} /* (3, 5, 27) {real, imag} */,
  {32'hc00a4f3e, 32'h410c1f89} /* (3, 5, 26) {real, imag} */,
  {32'hbfb6a9d3, 32'h410a4273} /* (3, 5, 25) {real, imag} */,
  {32'hc044435a, 32'h40d44398} /* (3, 5, 24) {real, imag} */,
  {32'hbfa5e8eb, 32'h40c81f12} /* (3, 5, 23) {real, imag} */,
  {32'hc0248e56, 32'h40c9ab02} /* (3, 5, 22) {real, imag} */,
  {32'hbf9c1336, 32'h40bbf53a} /* (3, 5, 21) {real, imag} */,
  {32'h3fdb65bd, 32'h40a20cad} /* (3, 5, 20) {real, imag} */,
  {32'h4023c2e7, 32'h405953ba} /* (3, 5, 19) {real, imag} */,
  {32'h40104467, 32'h3fc2dfb0} /* (3, 5, 18) {real, imag} */,
  {32'h3f166a8a, 32'h40286461} /* (3, 5, 17) {real, imag} */,
  {32'hbfa8fc38, 32'h3fcacd0a} /* (3, 5, 16) {real, imag} */,
  {32'h3faa3188, 32'hc09180df} /* (3, 5, 15) {real, imag} */,
  {32'h401708c4, 32'hc091b1f6} /* (3, 5, 14) {real, imag} */,
  {32'h40474bba, 32'hc0c792f1} /* (3, 5, 13) {real, imag} */,
  {32'h3fa862fc, 32'hc0ff8a1e} /* (3, 5, 12) {real, imag} */,
  {32'h40387b80, 32'hc0e10c44} /* (3, 5, 11) {real, imag} */,
  {32'h3fd751f8, 32'hbfdd477a} /* (3, 5, 10) {real, imag} */,
  {32'hbf766ec2, 32'hbea5bbe8} /* (3, 5, 9) {real, imag} */,
  {32'h3fa36036, 32'hbf1c378e} /* (3, 5, 8) {real, imag} */,
  {32'h3ff4ef0d, 32'h3f8aa11a} /* (3, 5, 7) {real, imag} */,
  {32'h3f1d2e04, 32'h3f93f626} /* (3, 5, 6) {real, imag} */,
  {32'hc0169a8e, 32'h409a39f4} /* (3, 5, 5) {real, imag} */,
  {32'hc0423246, 32'h40881f33} /* (3, 5, 4) {real, imag} */,
  {32'hbf9fc77d, 32'h403e2292} /* (3, 5, 3) {real, imag} */,
  {32'h3fa826c7, 32'h40873b66} /* (3, 5, 2) {real, imag} */,
  {32'h3f82cf17, 32'h40e4408f} /* (3, 5, 1) {real, imag} */,
  {32'hbf7ba3b4, 32'h40b1b16f} /* (3, 5, 0) {real, imag} */,
  {32'hc020a680, 32'h4060e288} /* (3, 4, 31) {real, imag} */,
  {32'hc005d34a, 32'h4095073c} /* (3, 4, 30) {real, imag} */,
  {32'h3f51a2bc, 32'h40825e46} /* (3, 4, 29) {real, imag} */,
  {32'hbf94c211, 32'h40fc21db} /* (3, 4, 28) {real, imag} */,
  {32'hc01e2685, 32'h4113d960} /* (3, 4, 27) {real, imag} */,
  {32'hc0207459, 32'h40fe1e6e} /* (3, 4, 26) {real, imag} */,
  {32'hbf9f894d, 32'h40d16aa4} /* (3, 4, 25) {real, imag} */,
  {32'hc091ce93, 32'h40bb837c} /* (3, 4, 24) {real, imag} */,
  {32'hc001b111, 32'h4087a940} /* (3, 4, 23) {real, imag} */,
  {32'hbf264955, 32'h40129e66} /* (3, 4, 22) {real, imag} */,
  {32'h3eb4b4d2, 32'h3fe723b9} /* (3, 4, 21) {real, imag} */,
  {32'hbf676bdb, 32'h40c63d8c} /* (3, 4, 20) {real, imag} */,
  {32'hbe45bbfe, 32'h40bfd534} /* (3, 4, 19) {real, imag} */,
  {32'hba8e4100, 32'h4092e091} /* (3, 4, 18) {real, imag} */,
  {32'h3f4e0678, 32'h40acdccb} /* (3, 4, 17) {real, imag} */,
  {32'hbf5c34f9, 32'h404dff78} /* (3, 4, 16) {real, imag} */,
  {32'h3fcc3c1e, 32'hc0cae614} /* (3, 4, 15) {real, imag} */,
  {32'h4076be20, 32'hc04939f4} /* (3, 4, 14) {real, imag} */,
  {32'h4015fb5c, 32'hc08b02c0} /* (3, 4, 13) {real, imag} */,
  {32'hbe0ffdd8, 32'hc0dd6402} /* (3, 4, 12) {real, imag} */,
  {32'h3e77d3a0, 32'hc0cad47b} /* (3, 4, 11) {real, imag} */,
  {32'h4032df9c, 32'hc0a1968e} /* (3, 4, 10) {real, imag} */,
  {32'h403b5299, 32'hbf9acb90} /* (3, 4, 9) {real, imag} */,
  {32'h4003a506, 32'hc0095675} /* (3, 4, 8) {real, imag} */,
  {32'h404892da, 32'hc03750b1} /* (3, 4, 7) {real, imag} */,
  {32'h3fe7c51f, 32'hc09d037a} /* (3, 4, 6) {real, imag} */,
  {32'hc031df10, 32'hbee7f9c9} /* (3, 4, 5) {real, imag} */,
  {32'hbfa1f2e4, 32'h402db69e} /* (3, 4, 4) {real, imag} */,
  {32'hc04f9281, 32'h4095f957} /* (3, 4, 3) {real, imag} */,
  {32'hc029ec14, 32'h409d413e} /* (3, 4, 2) {real, imag} */,
  {32'hbfe825ee, 32'h40bb5e0c} /* (3, 4, 1) {real, imag} */,
  {32'hbfb34724, 32'h4086589d} /* (3, 4, 0) {real, imag} */,
  {32'hc0176bd6, 32'h400db347} /* (3, 3, 31) {real, imag} */,
  {32'hc036a821, 32'h40ccb838} /* (3, 3, 30) {real, imag} */,
  {32'h3fdef498, 32'h40f92023} /* (3, 3, 29) {real, imag} */,
  {32'hbfbec5e8, 32'h41089daa} /* (3, 3, 28) {real, imag} */,
  {32'hc08182a9, 32'h4102f916} /* (3, 3, 27) {real, imag} */,
  {32'hc043fd00, 32'h40d5fbd3} /* (3, 3, 26) {real, imag} */,
  {32'hc00f8b9b, 32'h40b8651f} /* (3, 3, 25) {real, imag} */,
  {32'hc004b038, 32'h40b277c4} /* (3, 3, 24) {real, imag} */,
  {32'hbfceb00c, 32'h401ac16f} /* (3, 3, 23) {real, imag} */,
  {32'hbfa0302e, 32'h3eaeb4d6} /* (3, 3, 22) {real, imag} */,
  {32'hbf73dc22, 32'h404a115d} /* (3, 3, 21) {real, imag} */,
  {32'hc011a93f, 32'h40aa748b} /* (3, 3, 20) {real, imag} */,
  {32'hc0267a0f, 32'h409a2a5c} /* (3, 3, 19) {real, imag} */,
  {32'hc02dc48d, 32'h4071e2c0} /* (3, 3, 18) {real, imag} */,
  {32'hc00ddcea, 32'h40aef9cb} /* (3, 3, 17) {real, imag} */,
  {32'hc009ae40, 32'h409a1f7d} /* (3, 3, 16) {real, imag} */,
  {32'hbf3cc29a, 32'hc01b6bea} /* (3, 3, 15) {real, imag} */,
  {32'h3fec06b4, 32'hc0963dee} /* (3, 3, 14) {real, imag} */,
  {32'h3ff764e4, 32'hc0c87840} /* (3, 3, 13) {real, imag} */,
  {32'h3ed86a66, 32'hc0dd206f} /* (3, 3, 12) {real, imag} */,
  {32'hbfe6cf48, 32'hc0c2919e} /* (3, 3, 11) {real, imag} */,
  {32'h3e926560, 32'hc0ccafd2} /* (3, 3, 10) {real, imag} */,
  {32'h3fb4f755, 32'hbfdf2b2a} /* (3, 3, 9) {real, imag} */,
  {32'hbfc1217a, 32'hc02bbf0c} /* (3, 3, 8) {real, imag} */,
  {32'h3f4ce0d2, 32'hc0e3d674} /* (3, 3, 7) {real, imag} */,
  {32'h3f7a8397, 32'hc101d836} /* (3, 3, 6) {real, imag} */,
  {32'hc0417429, 32'hc04b9a48} /* (3, 3, 5) {real, imag} */,
  {32'hbf939c9b, 32'h3ff6ba1c} /* (3, 3, 4) {real, imag} */,
  {32'hc0ab3be8, 32'h40dcf364} /* (3, 3, 3) {real, imag} */,
  {32'hc091924d, 32'h40f47d6e} /* (3, 3, 2) {real, imag} */,
  {32'hc0311a24, 32'h40d0f5ef} /* (3, 3, 1) {real, imag} */,
  {32'hc00c633e, 32'h4072fef0} /* (3, 3, 0) {real, imag} */,
  {32'hc0447305, 32'h4017e3ac} /* (3, 2, 31) {real, imag} */,
  {32'hc0b7f99b, 32'h409e9d2f} /* (3, 2, 30) {real, imag} */,
  {32'hbff1bd5f, 32'h40fb14ac} /* (3, 2, 29) {real, imag} */,
  {32'hbf8a097a, 32'h40fb2db2} /* (3, 2, 28) {real, imag} */,
  {32'hbffb72d4, 32'h40c835d1} /* (3, 2, 27) {real, imag} */,
  {32'hbf132d95, 32'h40cd8666} /* (3, 2, 26) {real, imag} */,
  {32'hbfd1f94f, 32'h40cd054a} /* (3, 2, 25) {real, imag} */,
  {32'hc0356a8b, 32'h40801a82} /* (3, 2, 24) {real, imag} */,
  {32'hc035e6e6, 32'h3f94e2a2} /* (3, 2, 23) {real, imag} */,
  {32'hc0b5b828, 32'h40841513} /* (3, 2, 22) {real, imag} */,
  {32'hc08b5da0, 32'h410b427e} /* (3, 2, 21) {real, imag} */,
  {32'hbfa4f828, 32'h4113543c} /* (3, 2, 20) {real, imag} */,
  {32'hbf327ba6, 32'h40e1b94a} /* (3, 2, 19) {real, imag} */,
  {32'h3f9b5b16, 32'h40835031} /* (3, 2, 18) {real, imag} */,
  {32'hc016e6d1, 32'h40cb0f92} /* (3, 2, 17) {real, imag} */,
  {32'hc0bf7418, 32'h4018a166} /* (3, 2, 16) {real, imag} */,
  {32'hc05e9d17, 32'hc071dff3} /* (3, 2, 15) {real, imag} */,
  {32'h3f33f07a, 32'hc09efd54} /* (3, 2, 14) {real, imag} */,
  {32'h3f5fb81d, 32'hc0927e8a} /* (3, 2, 13) {real, imag} */,
  {32'hbf957517, 32'hc0ca1687} /* (3, 2, 12) {real, imag} */,
  {32'h3ec94c34, 32'hc0f50460} /* (3, 2, 11) {real, imag} */,
  {32'h3fa22ed2, 32'hc106fcdc} /* (3, 2, 10) {real, imag} */,
  {32'h3fcc2107, 32'hc10e4d94} /* (3, 2, 9) {real, imag} */,
  {32'hbefe1e76, 32'hc098f0cf} /* (3, 2, 8) {real, imag} */,
  {32'hbff2ffea, 32'hc0e5c952} /* (3, 2, 7) {real, imag} */,
  {32'h3f85b46a, 32'hc1219c84} /* (3, 2, 6) {real, imag} */,
  {32'h3f3524c8, 32'hbf9db1e9} /* (3, 2, 5) {real, imag} */,
  {32'h3db4ddc8, 32'h408c22c3} /* (3, 2, 4) {real, imag} */,
  {32'hc079fa98, 32'h40ad9b03} /* (3, 2, 3) {real, imag} */,
  {32'hc09705bc, 32'h40732f24} /* (3, 2, 2) {real, imag} */,
  {32'hc067d582, 32'h40a745da} /* (3, 2, 1) {real, imag} */,
  {32'hc017bfce, 32'h408ced7a} /* (3, 2, 0) {real, imag} */,
  {32'hbf9df608, 32'h3ff9d01c} /* (3, 1, 31) {real, imag} */,
  {32'hc015264d, 32'h4048b739} /* (3, 1, 30) {real, imag} */,
  {32'hbfbdb12c, 32'h4076e5df} /* (3, 1, 29) {real, imag} */,
  {32'h3e5bafda, 32'h4092f1ee} /* (3, 1, 28) {real, imag} */,
  {32'hbf5affa0, 32'h40bb7be4} /* (3, 1, 27) {real, imag} */,
  {32'hbf140ebe, 32'h40c86882} /* (3, 1, 26) {real, imag} */,
  {32'hbfa2b647, 32'h40d4a30b} /* (3, 1, 25) {real, imag} */,
  {32'hbfbe9011, 32'h408fed5e} /* (3, 1, 24) {real, imag} */,
  {32'hc067c494, 32'h400c36a2} /* (3, 1, 23) {real, imag} */,
  {32'hc06d1cbc, 32'h4083213c} /* (3, 1, 22) {real, imag} */,
  {32'hbf939799, 32'h40e4bc8e} /* (3, 1, 21) {real, imag} */,
  {32'hbf3f83f2, 32'h4089e6c2} /* (3, 1, 20) {real, imag} */,
  {32'hbe0ec798, 32'h40a33d8e} /* (3, 1, 19) {real, imag} */,
  {32'h3fadf332, 32'h40b148bc} /* (3, 1, 18) {real, imag} */,
  {32'hc0143646, 32'h40bfec40} /* (3, 1, 17) {real, imag} */,
  {32'hc08f6d25, 32'h406827f2} /* (3, 1, 16) {real, imag} */,
  {32'hbfdbe7e5, 32'hbfdb2fac} /* (3, 1, 15) {real, imag} */,
  {32'hbf0661fb, 32'hc079355b} /* (3, 1, 14) {real, imag} */,
  {32'h3eed5d84, 32'hc09bc014} /* (3, 1, 13) {real, imag} */,
  {32'h3febdcc2, 32'hc0d112a8} /* (3, 1, 12) {real, imag} */,
  {32'h403b4306, 32'hc10cc7a0} /* (3, 1, 11) {real, imag} */,
  {32'h40126db3, 32'hc0db73a4} /* (3, 1, 10) {real, imag} */,
  {32'h409dd165, 32'hc10d4d0a} /* (3, 1, 9) {real, imag} */,
  {32'h405e45ee, 32'hc0d1ee00} /* (3, 1, 8) {real, imag} */,
  {32'h3f5c9f08, 32'hc0c5c8a8} /* (3, 1, 7) {real, imag} */,
  {32'h4079cc94, 32'hc0ca592f} /* (3, 1, 6) {real, imag} */,
  {32'h40313855, 32'h3f2d8496} /* (3, 1, 5) {real, imag} */,
  {32'hbfb0ce43, 32'h40b09469} /* (3, 1, 4) {real, imag} */,
  {32'hc081cf32, 32'h40ad8334} /* (3, 1, 3) {real, imag} */,
  {32'hc055396a, 32'h40299013} /* (3, 1, 2) {real, imag} */,
  {32'hbf95143e, 32'h404c8fea} /* (3, 1, 1) {real, imag} */,
  {32'hbe913799, 32'h40286d07} /* (3, 1, 0) {real, imag} */,
  {32'hbf25587e, 32'h3f755ab3} /* (3, 0, 31) {real, imag} */,
  {32'hbfd90625, 32'h40039709} /* (3, 0, 30) {real, imag} */,
  {32'hbf294938, 32'h40310656} /* (3, 0, 29) {real, imag} */,
  {32'h3ee2f69b, 32'h3f993268} /* (3, 0, 28) {real, imag} */,
  {32'hbfce76a9, 32'h401a830c} /* (3, 0, 27) {real, imag} */,
  {32'hbfdcdc88, 32'h404a3fd8} /* (3, 0, 26) {real, imag} */,
  {32'hbe9194d2, 32'h4056ce43} /* (3, 0, 25) {real, imag} */,
  {32'h3f8926a2, 32'h4040f377} /* (3, 0, 24) {real, imag} */,
  {32'hbf398d3f, 32'h401e98ef} /* (3, 0, 23) {real, imag} */,
  {32'h3c84dcc0, 32'h400e36b7} /* (3, 0, 22) {real, imag} */,
  {32'h3f47b63e, 32'h3fce6d69} /* (3, 0, 21) {real, imag} */,
  {32'hc00952cb, 32'h3d8a98dc} /* (3, 0, 20) {real, imag} */,
  {32'hbfbca118, 32'h4000e4ca} /* (3, 0, 19) {real, imag} */,
  {32'hbf14cd99, 32'h407354a8} /* (3, 0, 18) {real, imag} */,
  {32'hbfe994a8, 32'h4040bc88} /* (3, 0, 17) {real, imag} */,
  {32'hbf932fba, 32'h4007a172} /* (3, 0, 16) {real, imag} */,
  {32'h3f98dd81, 32'h3d9e1ec4} /* (3, 0, 15) {real, imag} */,
  {32'h3e29a290, 32'hc06092da} /* (3, 0, 14) {real, imag} */,
  {32'h3efda7f6, 32'hc0a99562} /* (3, 0, 13) {real, imag} */,
  {32'h40080915, 32'hc08ac17c} /* (3, 0, 12) {real, imag} */,
  {32'h3fc7be93, 32'hc01edb8a} /* (3, 0, 11) {real, imag} */,
  {32'h3f7f7c20, 32'hbf1830a2} /* (3, 0, 10) {real, imag} */,
  {32'h40119950, 32'hc04137b4} /* (3, 0, 9) {real, imag} */,
  {32'h3fc88348, 32'hc0453b65} /* (3, 0, 8) {real, imag} */,
  {32'h3fa82e97, 32'hc0543dcb} /* (3, 0, 7) {real, imag} */,
  {32'h3ff9e7d7, 32'hc031e8f8} /* (3, 0, 6) {real, imag} */,
  {32'h3f4b4e2a, 32'h3f9996fb} /* (3, 0, 5) {real, imag} */,
  {32'hbd8b9742, 32'h40537325} /* (3, 0, 4) {real, imag} */,
  {32'hbf69412a, 32'h407f6a44} /* (3, 0, 3) {real, imag} */,
  {32'hbf7d2994, 32'h4071d448} /* (3, 0, 2) {real, imag} */,
  {32'hbf1bf15a, 32'h400ee712} /* (3, 0, 1) {real, imag} */,
  {32'hbeb9f424, 32'h3ef83b38} /* (3, 0, 0) {real, imag} */,
  {32'h3d01967e, 32'h406484f2} /* (2, 31, 31) {real, imag} */,
  {32'h3f571cc3, 32'h40c5fae4} /* (2, 31, 30) {real, imag} */,
  {32'hbfcc8416, 32'h40d66968} /* (2, 31, 29) {real, imag} */,
  {32'hc06914d1, 32'h41002642} /* (2, 31, 28) {real, imag} */,
  {32'hc035e531, 32'h41232dcb} /* (2, 31, 27) {real, imag} */,
  {32'hbfab88b7, 32'h4130cc3c} /* (2, 31, 26) {real, imag} */,
  {32'hbff75967, 32'h4116bc59} /* (2, 31, 25) {real, imag} */,
  {32'hbfedaf13, 32'h4111b4b6} /* (2, 31, 24) {real, imag} */,
  {32'hc01bc83f, 32'h40f37ce0} /* (2, 31, 23) {real, imag} */,
  {32'hc01f56fc, 32'h40fee966} /* (2, 31, 22) {real, imag} */,
  {32'hc00dbc31, 32'h40668e8a} /* (2, 31, 21) {real, imag} */,
  {32'h3e40eda6, 32'hc04ebf0d} /* (2, 31, 20) {real, imag} */,
  {32'h3f0a4e8f, 32'hc096e0a9} /* (2, 31, 19) {real, imag} */,
  {32'hbf85b1b8, 32'hc092b51a} /* (2, 31, 18) {real, imag} */,
  {32'hbf30783a, 32'hc09218d5} /* (2, 31, 17) {real, imag} */,
  {32'h3fa5e0a8, 32'hc0bfe476} /* (2, 31, 16) {real, imag} */,
  {32'h3fb6a424, 32'hc10171d2} /* (2, 31, 15) {real, imag} */,
  {32'h40271418, 32'hc1156335} /* (2, 31, 14) {real, imag} */,
  {32'h3fa26cd6, 32'hc1380c3f} /* (2, 31, 13) {real, imag} */,
  {32'h3f96b9ce, 32'hc102e7fc} /* (2, 31, 12) {real, imag} */,
  {32'h3fdd53ae, 32'hc0c5f0bb} /* (2, 31, 11) {real, imag} */,
  {32'hc0244d94, 32'h3fe2cc68} /* (2, 31, 10) {real, imag} */,
  {32'hbf625198, 32'h40f997be} /* (2, 31, 9) {real, imag} */,
  {32'hbfdb148c, 32'h40e5fcc8} /* (2, 31, 8) {real, imag} */,
  {32'hc086896d, 32'h40bd8844} /* (2, 31, 7) {real, imag} */,
  {32'hbfc4a4ce, 32'h4104697e} /* (2, 31, 6) {real, imag} */,
  {32'hbfb5f2a3, 32'h41173129} /* (2, 31, 5) {real, imag} */,
  {32'hbfa11c2e, 32'h41024bf7} /* (2, 31, 4) {real, imag} */,
  {32'hc006f431, 32'h40ea75a3} /* (2, 31, 3) {real, imag} */,
  {32'hc0119f1d, 32'h41262d3e} /* (2, 31, 2) {real, imag} */,
  {32'hbfb78eb0, 32'h40f4f4b9} /* (2, 31, 1) {real, imag} */,
  {32'hbfb3e2eb, 32'h407c73d8} /* (2, 31, 0) {real, imag} */,
  {32'hbff97500, 32'h40f2f2b5} /* (2, 30, 31) {real, imag} */,
  {32'hc02cc1c3, 32'h412f9ede} /* (2, 30, 30) {real, imag} */,
  {32'hc0add34c, 32'h411cfb2c} /* (2, 30, 29) {real, imag} */,
  {32'hc0eb2d76, 32'h4159af2a} /* (2, 30, 28) {real, imag} */,
  {32'hc0b53924, 32'h417678fb} /* (2, 30, 27) {real, imag} */,
  {32'hbffcbee2, 32'h417dcb0b} /* (2, 30, 26) {real, imag} */,
  {32'h3f956ad0, 32'h418bf9c8} /* (2, 30, 25) {real, imag} */,
  {32'h3f091831, 32'h41836d46} /* (2, 30, 24) {real, imag} */,
  {32'hbf5dc9e5, 32'h4173635f} /* (2, 30, 23) {real, imag} */,
  {32'hc0383bd8, 32'h416fac52} /* (2, 30, 22) {real, imag} */,
  {32'hbfe496ab, 32'h40dcf8da} /* (2, 30, 21) {real, imag} */,
  {32'h4059d509, 32'hc0dd545a} /* (2, 30, 20) {real, imag} */,
  {32'h407a7f15, 32'hc130790e} /* (2, 30, 19) {real, imag} */,
  {32'hbf2031c4, 32'hc13f5978} /* (2, 30, 18) {real, imag} */,
  {32'h3e51746e, 32'hc1472484} /* (2, 30, 17) {real, imag} */,
  {32'h403704b5, 32'hc150356a} /* (2, 30, 16) {real, imag} */,
  {32'h40484edc, 32'hc161a592} /* (2, 30, 15) {real, imag} */,
  {32'h40670428, 32'hc1803eee} /* (2, 30, 14) {real, imag} */,
  {32'h3fa0da62, 32'hc18af233} /* (2, 30, 13) {real, imag} */,
  {32'h3efd8fea, 32'hc17dcbf4} /* (2, 30, 12) {real, imag} */,
  {32'h3f877cf4, 32'hc117c0e8} /* (2, 30, 11) {real, imag} */,
  {32'hc04ffd9d, 32'h40cad558} /* (2, 30, 10) {real, imag} */,
  {32'hbfca73b4, 32'h417fc247} /* (2, 30, 9) {real, imag} */,
  {32'hc03be682, 32'h4148d753} /* (2, 30, 8) {real, imag} */,
  {32'hc0d0378c, 32'h413df1b8} /* (2, 30, 7) {real, imag} */,
  {32'hc03a25f4, 32'h41784a83} /* (2, 30, 6) {real, imag} */,
  {32'hc02ebc94, 32'h4176ac4c} /* (2, 30, 5) {real, imag} */,
  {32'hc0c4c026, 32'h4185bdf2} /* (2, 30, 4) {real, imag} */,
  {32'hc08ae32b, 32'h415df9e8} /* (2, 30, 3) {real, imag} */,
  {32'hc0d8f1e8, 32'h414eeb80} /* (2, 30, 2) {real, imag} */,
  {32'hbf16643d, 32'h4120e0b6} /* (2, 30, 1) {real, imag} */,
  {32'h3f566ce9, 32'h40b0a7ec} /* (2, 30, 0) {real, imag} */,
  {32'hc08fa42d, 32'h412704b7} /* (2, 29, 31) {real, imag} */,
  {32'hc08a9e6d, 32'h41887bfa} /* (2, 29, 30) {real, imag} */,
  {32'hc07fb06b, 32'h4150b0bf} /* (2, 29, 29) {real, imag} */,
  {32'hc08f8282, 32'h414279fa} /* (2, 29, 28) {real, imag} */,
  {32'hc00b76cc, 32'h4144be26} /* (2, 29, 27) {real, imag} */,
  {32'hbf28eefd, 32'h415bbc2e} /* (2, 29, 26) {real, imag} */,
  {32'h3fb4a9aa, 32'h41912eef} /* (2, 29, 25) {real, imag} */,
  {32'hc0398dcb, 32'h4185e91c} /* (2, 29, 24) {real, imag} */,
  {32'hc03ee124, 32'h418944f8} /* (2, 29, 23) {real, imag} */,
  {32'hc010471b, 32'h4166f80e} /* (2, 29, 22) {real, imag} */,
  {32'hbf015566, 32'h40763bb8} /* (2, 29, 21) {real, imag} */,
  {32'h40906642, 32'hc147e176} /* (2, 29, 20) {real, imag} */,
  {32'h40759a4c, 32'hc182d0d4} /* (2, 29, 19) {real, imag} */,
  {32'h4017e9a0, 32'hc1743d3f} /* (2, 29, 18) {real, imag} */,
  {32'h4025c351, 32'hc182e302} /* (2, 29, 17) {real, imag} */,
  {32'h4058be03, 32'hc189af5e} /* (2, 29, 16) {real, imag} */,
  {32'h408b1f7e, 32'hc174035e} /* (2, 29, 15) {real, imag} */,
  {32'h4066c90a, 32'hc16d87ef} /* (2, 29, 14) {real, imag} */,
  {32'h40909910, 32'hc16cdc6a} /* (2, 29, 13) {real, imag} */,
  {32'h40756f2a, 32'hc17cfc76} /* (2, 29, 12) {real, imag} */,
  {32'h4050d7a4, 32'hc1128a2b} /* (2, 29, 11) {real, imag} */,
  {32'hc02eccb9, 32'h40beb67b} /* (2, 29, 10) {real, imag} */,
  {32'hc0918eb0, 32'h41662d39} /* (2, 29, 9) {real, imag} */,
  {32'hc099aa87, 32'h413e4b4a} /* (2, 29, 8) {real, imag} */,
  {32'hc083fbe0, 32'h4138436f} /* (2, 29, 7) {real, imag} */,
  {32'hc0745f33, 32'h4156363c} /* (2, 29, 6) {real, imag} */,
  {32'hc0860080, 32'h41687ecc} /* (2, 29, 5) {real, imag} */,
  {32'hc109ff19, 32'h418b6154} /* (2, 29, 4) {real, imag} */,
  {32'hc0e327d4, 32'h416af390} /* (2, 29, 3) {real, imag} */,
  {32'hc0a120cf, 32'h4130babc} /* (2, 29, 2) {real, imag} */,
  {32'hbf63b60d, 32'h4136758f} /* (2, 29, 1) {real, imag} */,
  {32'hbfb07cd1, 32'h40ed4158} /* (2, 29, 0) {real, imag} */,
  {32'hc062570a, 32'h40f60d90} /* (2, 28, 31) {real, imag} */,
  {32'hc02e7abc, 32'h4183801b} /* (2, 28, 30) {real, imag} */,
  {32'hbf7df1c6, 32'h4179a8d8} /* (2, 28, 29) {real, imag} */,
  {32'hc02fe32d, 32'h416d36ce} /* (2, 28, 28) {real, imag} */,
  {32'hbfa78496, 32'h417401ad} /* (2, 28, 27) {real, imag} */,
  {32'h3ea5f1a9, 32'h416f687a} /* (2, 28, 26) {real, imag} */,
  {32'hbf16715e, 32'h417687e8} /* (2, 28, 25) {real, imag} */,
  {32'hc0ba2ace, 32'h4184789d} /* (2, 28, 24) {real, imag} */,
  {32'hc0ae36c0, 32'h4186c194} /* (2, 28, 23) {real, imag} */,
  {32'hbfd4e9c1, 32'h416f07ce} /* (2, 28, 22) {real, imag} */,
  {32'h3fb40d97, 32'h40a6bc74} /* (2, 28, 21) {real, imag} */,
  {32'h40306d4d, 32'hc14c80a3} /* (2, 28, 20) {real, imag} */,
  {32'h4012cc22, 32'hc18bdbd6} /* (2, 28, 19) {real, imag} */,
  {32'h404bf77e, 32'hc16bc2b4} /* (2, 28, 18) {real, imag} */,
  {32'h4058f32e, 32'hc168ae62} /* (2, 28, 17) {real, imag} */,
  {32'h40599de7, 32'hc1882094} /* (2, 28, 16) {real, imag} */,
  {32'h409fec38, 32'hc1807ed9} /* (2, 28, 15) {real, imag} */,
  {32'h40a35f5e, 32'hc14a690b} /* (2, 28, 14) {real, imag} */,
  {32'h40baff0f, 32'hc1433171} /* (2, 28, 13) {real, imag} */,
  {32'h40862042, 32'hc16e5923} /* (2, 28, 12) {real, imag} */,
  {32'h4024afe2, 32'hc13254ac} /* (2, 28, 11) {real, imag} */,
  {32'hbff6cca6, 32'h406c8f43} /* (2, 28, 10) {real, imag} */,
  {32'hc06385d0, 32'h4178d51a} /* (2, 28, 9) {real, imag} */,
  {32'hbfa7377a, 32'h4180bc54} /* (2, 28, 8) {real, imag} */,
  {32'hc0478616, 32'h41604f44} /* (2, 28, 7) {real, imag} */,
  {32'hc03dff8c, 32'h416a1b2c} /* (2, 28, 6) {real, imag} */,
  {32'hc07323b7, 32'h416d1e73} /* (2, 28, 5) {real, imag} */,
  {32'hc0d6b6ea, 32'h416cac17} /* (2, 28, 4) {real, imag} */,
  {32'hc0b50d72, 32'h414389c3} /* (2, 28, 3) {real, imag} */,
  {32'hc08ac776, 32'h41479271} /* (2, 28, 2) {real, imag} */,
  {32'hc008a0bf, 32'h414dda9a} /* (2, 28, 1) {real, imag} */,
  {32'hbf986316, 32'h4112f82d} /* (2, 28, 0) {real, imag} */,
  {32'hc04c1ee4, 32'h40f6dd73} /* (2, 27, 31) {real, imag} */,
  {32'hc01f0f72, 32'h417f78c6} /* (2, 27, 30) {real, imag} */,
  {32'hc0492120, 32'h4183b549} /* (2, 27, 29) {real, imag} */,
  {32'hc030266c, 32'h4184bcdc} /* (2, 27, 28) {real, imag} */,
  {32'hbe3151c8, 32'h418ca6e4} /* (2, 27, 27) {real, imag} */,
  {32'h3f1c0601, 32'h417e9f0c} /* (2, 27, 26) {real, imag} */,
  {32'hbf81189f, 32'h417f9b12} /* (2, 27, 25) {real, imag} */,
  {32'hc0968457, 32'h4182acd8} /* (2, 27, 24) {real, imag} */,
  {32'hc1055670, 32'h417ac879} /* (2, 27, 23) {real, imag} */,
  {32'hc03b7457, 32'h416e2e40} /* (2, 27, 22) {real, imag} */,
  {32'h4038bf7c, 32'h40e7fc3e} /* (2, 27, 21) {real, imag} */,
  {32'h40adb724, 32'hc10cddc8} /* (2, 27, 20) {real, imag} */,
  {32'h4093ace4, 32'hc163c620} /* (2, 27, 19) {real, imag} */,
  {32'h4046d3a5, 32'hc16b9b61} /* (2, 27, 18) {real, imag} */,
  {32'h40a8e5b8, 32'hc166ee20} /* (2, 27, 17) {real, imag} */,
  {32'h4088d543, 32'hc16020e3} /* (2, 27, 16) {real, imag} */,
  {32'h4089a02b, 32'hc1879417} /* (2, 27, 15) {real, imag} */,
  {32'h40a83880, 32'hc15eb8a2} /* (2, 27, 14) {real, imag} */,
  {32'h408159af, 32'hc13ad5fe} /* (2, 27, 13) {real, imag} */,
  {32'h406caec0, 32'hc14d2f4f} /* (2, 27, 12) {real, imag} */,
  {32'h3fdb74d9, 32'hc13fb2f6} /* (2, 27, 11) {real, imag} */,
  {32'hbd1873a0, 32'h40b27098} /* (2, 27, 10) {real, imag} */,
  {32'h3f1552fe, 32'h41812fdc} /* (2, 27, 9) {real, imag} */,
  {32'hbfb5a81a, 32'h4183682e} /* (2, 27, 8) {real, imag} */,
  {32'hc0a1668d, 32'h4179d131} /* (2, 27, 7) {real, imag} */,
  {32'hc0266652, 32'h418c6e24} /* (2, 27, 6) {real, imag} */,
  {32'hc082f97c, 32'h418f7ef6} /* (2, 27, 5) {real, imag} */,
  {32'hc0acfd90, 32'h4171eed2} /* (2, 27, 4) {real, imag} */,
  {32'hbf84d202, 32'h415f33e4} /* (2, 27, 3) {real, imag} */,
  {32'hc0381f15, 32'h41696f32} /* (2, 27, 2) {real, imag} */,
  {32'hc09ef037, 32'h41557ef2} /* (2, 27, 1) {real, imag} */,
  {32'hc02f7741, 32'h4114bc07} /* (2, 27, 0) {real, imag} */,
  {32'hc0597787, 32'h40d22497} /* (2, 26, 31) {real, imag} */,
  {32'hc0577822, 32'h414d3ae4} /* (2, 26, 30) {real, imag} */,
  {32'hc042d31a, 32'h415f004d} /* (2, 26, 29) {real, imag} */,
  {32'hbfd72f06, 32'h414e9584} /* (2, 26, 28) {real, imag} */,
  {32'h3f413b22, 32'h4158091a} /* (2, 26, 27) {real, imag} */,
  {32'hbf2e56ce, 32'h41651f9c} /* (2, 26, 26) {real, imag} */,
  {32'hc02d2e70, 32'h418f994d} /* (2, 26, 25) {real, imag} */,
  {32'hc048e3ee, 32'h4193844f} /* (2, 26, 24) {real, imag} */,
  {32'hc08004a5, 32'h417cf510} /* (2, 26, 23) {real, imag} */,
  {32'hc0370346, 32'h415f445a} /* (2, 26, 22) {real, imag} */,
  {32'h3fc9d830, 32'h40a81412} /* (2, 26, 21) {real, imag} */,
  {32'h4096eb5e, 32'hc11c04ce} /* (2, 26, 20) {real, imag} */,
  {32'h40803979, 32'hc1482370} /* (2, 26, 19) {real, imag} */,
  {32'h3ec027ca, 32'hc15b9c7c} /* (2, 26, 18) {real, imag} */,
  {32'h4056eab4, 32'hc16815da} /* (2, 26, 17) {real, imag} */,
  {32'h4048e249, 32'hc16a0b57} /* (2, 26, 16) {real, imag} */,
  {32'h404d3e7f, 32'hc18c4606} /* (2, 26, 15) {real, imag} */,
  {32'h40a78b48, 32'hc17e13b6} /* (2, 26, 14) {real, imag} */,
  {32'h40788fea, 32'hc1595f06} /* (2, 26, 13) {real, imag} */,
  {32'h40104e11, 32'hc1725806} /* (2, 26, 12) {real, imag} */,
  {32'h4013fd9a, 32'hc1274984} /* (2, 26, 11) {real, imag} */,
  {32'h3ebe3786, 32'h4087eda8} /* (2, 26, 10) {real, imag} */,
  {32'hc086f1ab, 32'h416d2ff0} /* (2, 26, 9) {real, imag} */,
  {32'hc0a95b3a, 32'h41881d28} /* (2, 26, 8) {real, imag} */,
  {32'hc019d0e2, 32'h415a7c25} /* (2, 26, 7) {real, imag} */,
  {32'hbf8b5922, 32'h414ad9c2} /* (2, 26, 6) {real, imag} */,
  {32'hc087d0c0, 32'h41553276} /* (2, 26, 5) {real, imag} */,
  {32'hc095c716, 32'h41419e8d} /* (2, 26, 4) {real, imag} */,
  {32'hbf32cd1b, 32'h415c6620} /* (2, 26, 3) {real, imag} */,
  {32'hc06d9aea, 32'h417ef46f} /* (2, 26, 2) {real, imag} */,
  {32'hc0c4fc10, 32'h415818dd} /* (2, 26, 1) {real, imag} */,
  {32'hc059fd4f, 32'h410c9b3a} /* (2, 26, 0) {real, imag} */,
  {32'hc008c0ca, 32'h40f945dc} /* (2, 25, 31) {real, imag} */,
  {32'hc0103faf, 32'h414fcb81} /* (2, 25, 30) {real, imag} */,
  {32'hbffa9420, 32'h41673317} /* (2, 25, 29) {real, imag} */,
  {32'hc031f468, 32'h416a0e09} /* (2, 25, 28) {real, imag} */,
  {32'hbf431873, 32'h417bc2e8} /* (2, 25, 27) {real, imag} */,
  {32'hc00e9591, 32'h417bb100} /* (2, 25, 26) {real, imag} */,
  {32'hc0156ab6, 32'h419aab18} /* (2, 25, 25) {real, imag} */,
  {32'hbf99551f, 32'h4187b78e} /* (2, 25, 24) {real, imag} */,
  {32'hbfe2f5fd, 32'h4164064d} /* (2, 25, 23) {real, imag} */,
  {32'hbfe307b1, 32'h4186d0c8} /* (2, 25, 22) {real, imag} */,
  {32'h3d344cb8, 32'h40fb1c0f} /* (2, 25, 21) {real, imag} */,
  {32'h405db358, 32'hc14aab16} /* (2, 25, 20) {real, imag} */,
  {32'h40abc648, 32'hc16dda26} /* (2, 25, 19) {real, imag} */,
  {32'h3fbbfe65, 32'hc16a55ed} /* (2, 25, 18) {real, imag} */,
  {32'h3fc7af9b, 32'hc1787799} /* (2, 25, 17) {real, imag} */,
  {32'h3fe2cccf, 32'hc16c4e5a} /* (2, 25, 16) {real, imag} */,
  {32'h405bdc97, 32'hc1800671} /* (2, 25, 15) {real, imag} */,
  {32'h3f808440, 32'hc18179ee} /* (2, 25, 14) {real, imag} */,
  {32'hbf78214f, 32'hc169c6d2} /* (2, 25, 13) {real, imag} */,
  {32'h4011058e, 32'hc1745a83} /* (2, 25, 12) {real, imag} */,
  {32'h40b743fa, 32'hc13a6962} /* (2, 25, 11) {real, imag} */,
  {32'h3f8e91a0, 32'h409b8f27} /* (2, 25, 10) {real, imag} */,
  {32'hc0b62fa0, 32'h4185442c} /* (2, 25, 9) {real, imag} */,
  {32'hc08c087c, 32'h41a65d98} /* (2, 25, 8) {real, imag} */,
  {32'hc0598fbc, 32'h416e6062} /* (2, 25, 7) {real, imag} */,
  {32'hc01e9f24, 32'h414e868a} /* (2, 25, 6) {real, imag} */,
  {32'hc02d8a1a, 32'h41735ebc} /* (2, 25, 5) {real, imag} */,
  {32'hc050325f, 32'h41674787} /* (2, 25, 4) {real, imag} */,
  {32'hc01aed4e, 32'h414f58c6} /* (2, 25, 3) {real, imag} */,
  {32'hc0869e79, 32'h4181abc0} /* (2, 25, 2) {real, imag} */,
  {32'hc0c77a0a, 32'h414e992a} /* (2, 25, 1) {real, imag} */,
  {32'hc0330ce2, 32'h40fd2c58} /* (2, 25, 0) {real, imag} */,
  {32'hbff96bc3, 32'h40c5f43a} /* (2, 24, 31) {real, imag} */,
  {32'hc00e3698, 32'h413f4091} /* (2, 24, 30) {real, imag} */,
  {32'h3f621614, 32'h415866ec} /* (2, 24, 29) {real, imag} */,
  {32'hbffaf4dd, 32'h41601451} /* (2, 24, 28) {real, imag} */,
  {32'hc0a7fdb2, 32'h4176b026} /* (2, 24, 27) {real, imag} */,
  {32'hc0b81b27, 32'h416bd699} /* (2, 24, 26) {real, imag} */,
  {32'hc0504354, 32'h417e1b6c} /* (2, 24, 25) {real, imag} */,
  {32'hc0419962, 32'h41711b77} /* (2, 24, 24) {real, imag} */,
  {32'hc013c6ac, 32'h4160c720} /* (2, 24, 23) {real, imag} */,
  {32'hbf85dcbe, 32'h4174543f} /* (2, 24, 22) {real, imag} */,
  {32'h3f63c68b, 32'h40b0eb6e} /* (2, 24, 21) {real, imag} */,
  {32'h40d815fe, 32'hc16ce95a} /* (2, 24, 20) {real, imag} */,
  {32'h40cab6ba, 32'hc1828528} /* (2, 24, 19) {real, imag} */,
  {32'h400ffc6e, 32'hc17778f9} /* (2, 24, 18) {real, imag} */,
  {32'h3fb48675, 32'hc1734ff8} /* (2, 24, 17) {real, imag} */,
  {32'hbec8c092, 32'hc1811c12} /* (2, 24, 16) {real, imag} */,
  {32'h3fd6c809, 32'hc185474e} /* (2, 24, 15) {real, imag} */,
  {32'hbf4587ce, 32'hc183df40} /* (2, 24, 14) {real, imag} */,
  {32'h3f967bdb, 32'hc153994e} /* (2, 24, 13) {real, imag} */,
  {32'h40b7138c, 32'hc172fe7a} /* (2, 24, 12) {real, imag} */,
  {32'h4062733b, 32'hc155b8f2} /* (2, 24, 11) {real, imag} */,
  {32'hc0ae1b33, 32'h40ce1a20} /* (2, 24, 10) {real, imag} */,
  {32'hc0d84288, 32'h419c959a} /* (2, 24, 9) {real, imag} */,
  {32'hc040964a, 32'h41b513a0} /* (2, 24, 8) {real, imag} */,
  {32'hc03d13ec, 32'h419397ca} /* (2, 24, 7) {real, imag} */,
  {32'hc0339986, 32'h417699d1} /* (2, 24, 6) {real, imag} */,
  {32'hc00beac7, 32'h413e3e3c} /* (2, 24, 5) {real, imag} */,
  {32'hc016dbfa, 32'h41300aa9} /* (2, 24, 4) {real, imag} */,
  {32'hc02cbefe, 32'h4166473f} /* (2, 24, 3) {real, imag} */,
  {32'hc0ae24fe, 32'h41827d6e} /* (2, 24, 2) {real, imag} */,
  {32'hc0a8f2ac, 32'h414261c2} /* (2, 24, 1) {real, imag} */,
  {32'hc00a6af2, 32'h40d2d48e} /* (2, 24, 0) {real, imag} */,
  {32'hbf99b3c2, 32'h40c5b6e7} /* (2, 23, 31) {real, imag} */,
  {32'hbfcf2aff, 32'h414f4ecd} /* (2, 23, 30) {real, imag} */,
  {32'hbbdf1680, 32'h41649f21} /* (2, 23, 29) {real, imag} */,
  {32'hc01c65e3, 32'h416d10a7} /* (2, 23, 28) {real, imag} */,
  {32'hc0bd678e, 32'h4170a1e8} /* (2, 23, 27) {real, imag} */,
  {32'hc09a6115, 32'h4151c546} /* (2, 23, 26) {real, imag} */,
  {32'hbfdf426b, 32'h412b6ba2} /* (2, 23, 25) {real, imag} */,
  {32'hc024db88, 32'h414de7e0} /* (2, 23, 24) {real, imag} */,
  {32'hbfa98bc6, 32'h4181a5d2} /* (2, 23, 23) {real, imag} */,
  {32'hbe33991c, 32'h4176c391} /* (2, 23, 22) {real, imag} */,
  {32'hbf50d3e6, 32'h40d6eb04} /* (2, 23, 21) {real, imag} */,
  {32'h408d1869, 32'hc154bf02} /* (2, 23, 20) {real, imag} */,
  {32'h4082711f, 32'hc18bd736} /* (2, 23, 19) {real, imag} */,
  {32'h3fc8525d, 32'hc1929d8b} /* (2, 23, 18) {real, imag} */,
  {32'h3f894077, 32'hc172267c} /* (2, 23, 17) {real, imag} */,
  {32'hbdc07718, 32'hc16be15c} /* (2, 23, 16) {real, imag} */,
  {32'hbfa29050, 32'hc14b28ef} /* (2, 23, 15) {real, imag} */,
  {32'hbe8e5856, 32'hc16be773} /* (2, 23, 14) {real, imag} */,
  {32'h408447e8, 32'hc151091a} /* (2, 23, 13) {real, imag} */,
  {32'h409d1556, 32'hc15dd9c0} /* (2, 23, 12) {real, imag} */,
  {32'h406891da, 32'hc1415546} /* (2, 23, 11) {real, imag} */,
  {32'hc07228ea, 32'h40af59be} /* (2, 23, 10) {real, imag} */,
  {32'hc09db60f, 32'h4179ca1a} /* (2, 23, 9) {real, imag} */,
  {32'hc07dc1b6, 32'h418e0b05} /* (2, 23, 8) {real, imag} */,
  {32'hc031d48e, 32'h4189ffee} /* (2, 23, 7) {real, imag} */,
  {32'hbff50aad, 32'h415f198d} /* (2, 23, 6) {real, imag} */,
  {32'h3ebace82, 32'h415048a8} /* (2, 23, 5) {real, imag} */,
  {32'hbef7bfec, 32'h414d5724} /* (2, 23, 4) {real, imag} */,
  {32'hbff42819, 32'h4181a1ac} /* (2, 23, 3) {real, imag} */,
  {32'hc08c60d6, 32'h416feaee} /* (2, 23, 2) {real, imag} */,
  {32'hc0291170, 32'h415e3d20} /* (2, 23, 1) {real, imag} */,
  {32'h3f4c755c, 32'h40e4e965} /* (2, 23, 0) {real, imag} */,
  {32'hbe664b64, 32'h41011560} /* (2, 22, 31) {real, imag} */,
  {32'hbedfb97e, 32'h41881d72} /* (2, 22, 30) {real, imag} */,
  {32'hbf909aa7, 32'h418b5d39} /* (2, 22, 29) {real, imag} */,
  {32'hc05db881, 32'h417d350e} /* (2, 22, 28) {real, imag} */,
  {32'hc0c79db0, 32'h4145b610} /* (2, 22, 27) {real, imag} */,
  {32'hc0b5ed42, 32'h4130743c} /* (2, 22, 26) {real, imag} */,
  {32'hc07460d8, 32'h41086ebe} /* (2, 22, 25) {real, imag} */,
  {32'hbfdc6d6a, 32'h413f3eac} /* (2, 22, 24) {real, imag} */,
  {32'hbfb204a2, 32'h4180301b} /* (2, 22, 23) {real, imag} */,
  {32'hbf77aba6, 32'h4161b7d2} /* (2, 22, 22) {real, imag} */,
  {32'hc042607a, 32'h40b549b4} /* (2, 22, 21) {real, imag} */,
  {32'h3fd5d75c, 32'hc14ab91f} /* (2, 22, 20) {real, imag} */,
  {32'h3fc2f339, 32'hc181c484} /* (2, 22, 19) {real, imag} */,
  {32'hbf6ba41c, 32'hc16e80b2} /* (2, 22, 18) {real, imag} */,
  {32'h3f8664f8, 32'hc14e6e33} /* (2, 22, 17) {real, imag} */,
  {32'h3f3263be, 32'hc14b334e} /* (2, 22, 16) {real, imag} */,
  {32'h3e6388c8, 32'hc116b692} /* (2, 22, 15) {real, imag} */,
  {32'h4078ed4a, 32'hc14c8c9f} /* (2, 22, 14) {real, imag} */,
  {32'h4078ffa8, 32'hc16ca544} /* (2, 22, 13) {real, imag} */,
  {32'h3f975a96, 32'hc148b194} /* (2, 22, 12) {real, imag} */,
  {32'h3e6432f8, 32'hc11cd6e9} /* (2, 22, 11) {real, imag} */,
  {32'hc050a57a, 32'h40acaf4a} /* (2, 22, 10) {real, imag} */,
  {32'hc0543203, 32'h415a7c82} /* (2, 22, 9) {real, imag} */,
  {32'hc0593bc6, 32'h4168eb24} /* (2, 22, 8) {real, imag} */,
  {32'hc030b0f4, 32'h416ff3de} /* (2, 22, 7) {real, imag} */,
  {32'hc015d188, 32'h4145733c} /* (2, 22, 6) {real, imag} */,
  {32'hbd7b0130, 32'h414ae50d} /* (2, 22, 5) {real, imag} */,
  {32'h3faf658c, 32'h41687224} /* (2, 22, 4) {real, imag} */,
  {32'hbffceab1, 32'h4179b170} /* (2, 22, 3) {real, imag} */,
  {32'hc083dbe7, 32'h418bc943} /* (2, 22, 2) {real, imag} */,
  {32'hc00c3e33, 32'h4192fc22} /* (2, 22, 1) {real, imag} */,
  {32'hbeccc8f5, 32'h411f83fe} /* (2, 22, 0) {real, imag} */,
  {32'hbf908741, 32'h4084b31c} /* (2, 21, 31) {real, imag} */,
  {32'hbf9f9087, 32'h40ccf566} /* (2, 21, 30) {real, imag} */,
  {32'hbea55982, 32'h40d101ae} /* (2, 21, 29) {real, imag} */,
  {32'hc03cf67f, 32'h40a14d9d} /* (2, 21, 28) {real, imag} */,
  {32'hc0ac3783, 32'h4052459d} /* (2, 21, 27) {real, imag} */,
  {32'hc0952e2f, 32'h408b7560} /* (2, 21, 26) {real, imag} */,
  {32'hc008434e, 32'h3f15193c} /* (2, 21, 25) {real, imag} */,
  {32'hbf2dc041, 32'h405cae9e} /* (2, 21, 24) {real, imag} */,
  {32'hbed0d976, 32'h4089e9ec} /* (2, 21, 23) {real, imag} */,
  {32'hbf8fc93e, 32'h40a19827} /* (2, 21, 22) {real, imag} */,
  {32'hc04741b1, 32'h40900ad0} /* (2, 21, 21) {real, imag} */,
  {32'h40010dbc, 32'hbfe86169} /* (2, 21, 20) {real, imag} */,
  {32'h402e0886, 32'hc0f0c79a} /* (2, 21, 19) {real, imag} */,
  {32'hbf91531c, 32'hc097eeca} /* (2, 21, 18) {real, imag} */,
  {32'hbf62a262, 32'hc0729006} /* (2, 21, 17) {real, imag} */,
  {32'hbec3d879, 32'hc0833532} /* (2, 21, 16) {real, imag} */,
  {32'h3f8914b4, 32'hc091c06a} /* (2, 21, 15) {real, imag} */,
  {32'hbe1d126c, 32'hc0f3c040} /* (2, 21, 14) {real, imag} */,
  {32'hbff18174, 32'hc0c6c987} /* (2, 21, 13) {real, imag} */,
  {32'hc0338ab0, 32'hc07e1a66} /* (2, 21, 12) {real, imag} */,
  {32'h3f536a0a, 32'hc097ef96} /* (2, 21, 11) {real, imag} */,
  {32'hbf23f6b6, 32'h401444d2} /* (2, 21, 10) {real, imag} */,
  {32'hbf0f2ed6, 32'h40dcab18} /* (2, 21, 9) {real, imag} */,
  {32'hbe833504, 32'h408e9da6} /* (2, 21, 8) {real, imag} */,
  {32'h3f070205, 32'h409d6582} /* (2, 21, 7) {real, imag} */,
  {32'hbfb19111, 32'h40824589} /* (2, 21, 6) {real, imag} */,
  {32'hbeb90d37, 32'h403fecff} /* (2, 21, 5) {real, imag} */,
  {32'h40021654, 32'h40efd75e} /* (2, 21, 4) {real, imag} */,
  {32'hbfa04006, 32'h40e046ac} /* (2, 21, 3) {real, imag} */,
  {32'hc0827c18, 32'h40d70af2} /* (2, 21, 2) {real, imag} */,
  {32'hbfecc51a, 32'h4107c4fb} /* (2, 21, 1) {real, imag} */,
  {32'hbf815597, 32'h40a475cc} /* (2, 21, 0) {real, imag} */,
  {32'h3e36e7ea, 32'hc0ca08e6} /* (2, 20, 31) {real, imag} */,
  {32'h3f8d8ba4, 32'hc150bf8a} /* (2, 20, 30) {real, imag} */,
  {32'hbece3a24, 32'hc1436925} /* (2, 20, 29) {real, imag} */,
  {32'hbfa1c225, 32'hc16a96a6} /* (2, 20, 28) {real, imag} */,
  {32'hc047e75c, 32'hc14debcc} /* (2, 20, 27) {real, imag} */,
  {32'hc0365f14, 32'hc1024d8a} /* (2, 20, 26) {real, imag} */,
  {32'h40353848, 32'hc16a7aaf} /* (2, 20, 25) {real, imag} */,
  {32'h400a30fc, 32'hc17fce40} /* (2, 20, 24) {real, imag} */,
  {32'hbd97b7b0, 32'hc1372cd8} /* (2, 20, 23) {real, imag} */,
  {32'h3f3629be, 32'hc127246d} /* (2, 20, 22) {real, imag} */,
  {32'hbfc8a0c4, 32'hc032c8ec} /* (2, 20, 21) {real, imag} */,
  {32'hbf8fed04, 32'h410b3c12} /* (2, 20, 20) {real, imag} */,
  {32'h3da85340, 32'h41003e74} /* (2, 20, 19) {real, imag} */,
  {32'hbf9304aa, 32'h4119bbc2} /* (2, 20, 18) {real, imag} */,
  {32'hbe8722da, 32'h4144120c} /* (2, 20, 17) {real, imag} */,
  {32'hbf251f1e, 32'h413cbd86} /* (2, 20, 16) {real, imag} */,
  {32'hbfb3941f, 32'h411f38f2} /* (2, 20, 15) {real, imag} */,
  {32'hc0559ec0, 32'h411599f5} /* (2, 20, 14) {real, imag} */,
  {32'hc0400bc2, 32'h41432304} /* (2, 20, 13) {real, imag} */,
  {32'hc089fb10, 32'h4144dab2} /* (2, 20, 12) {real, imag} */,
  {32'hbf194392, 32'h41011956} /* (2, 20, 11) {real, imag} */,
  {32'h3f8f3142, 32'hc0a181d7} /* (2, 20, 10) {real, imag} */,
  {32'h3ffb5890, 32'hc1044714} /* (2, 20, 9) {real, imag} */,
  {32'h40454258, 32'hc1003b87} /* (2, 20, 8) {real, imag} */,
  {32'h402d7ef0, 32'hc1262899} /* (2, 20, 7) {real, imag} */,
  {32'h3d99fb08, 32'hc14cc296} /* (2, 20, 6) {real, imag} */,
  {32'h3fd3f01c, 32'hc179d006} /* (2, 20, 5) {real, imag} */,
  {32'h3fc2b674, 32'hc11f88ba} /* (2, 20, 4) {real, imag} */,
  {32'h400aa68d, 32'hc12224e4} /* (2, 20, 3) {real, imag} */,
  {32'h402bc168, 32'hc159d878} /* (2, 20, 2) {real, imag} */,
  {32'h3fd6a2c8, 32'hc1160dd2} /* (2, 20, 1) {real, imag} */,
  {32'hbf08c9fc, 32'hc069bdf6} /* (2, 20, 0) {real, imag} */,
  {32'h3f89c3c0, 32'hc101939e} /* (2, 19, 31) {real, imag} */,
  {32'h400e03d8, 32'hc1714ef3} /* (2, 19, 30) {real, imag} */,
  {32'h3ffe87fb, 32'hc16684e3} /* (2, 19, 29) {real, imag} */,
  {32'h3fa1354c, 32'hc18024fc} /* (2, 19, 28) {real, imag} */,
  {32'hbf347415, 32'hc170dcde} /* (2, 19, 27) {real, imag} */,
  {32'h3f492915, 32'hc13261fe} /* (2, 19, 26) {real, imag} */,
  {32'h4087cc45, 32'hc153ef83} /* (2, 19, 25) {real, imag} */,
  {32'h40c8bde2, 32'hc18965a8} /* (2, 19, 24) {real, imag} */,
  {32'h404f0c54, 32'hc16f58b9} /* (2, 19, 23) {real, imag} */,
  {32'h404dd98e, 32'hc15fb9ad} /* (2, 19, 22) {real, imag} */,
  {32'h3f5f82ad, 32'hc08a0d4e} /* (2, 19, 21) {real, imag} */,
  {32'hc05ddf86, 32'h414a3092} /* (2, 19, 20) {real, imag} */,
  {32'hc026097c, 32'h415a799a} /* (2, 19, 19) {real, imag} */,
  {32'hbef65a27, 32'h414d5e90} /* (2, 19, 18) {real, imag} */,
  {32'hc021fa2f, 32'h415191c7} /* (2, 19, 17) {real, imag} */,
  {32'hc077508a, 32'h4181d836} /* (2, 19, 16) {real, imag} */,
  {32'hc0a74bba, 32'h4197e2fc} /* (2, 19, 15) {real, imag} */,
  {32'hc08307e0, 32'h4170174e} /* (2, 19, 14) {real, imag} */,
  {32'hbf4f46ad, 32'h41736589} /* (2, 19, 13) {real, imag} */,
  {32'h3e568d6c, 32'h417c5194} /* (2, 19, 12) {real, imag} */,
  {32'hbfb0ce62, 32'h415aeb46} /* (2, 19, 11) {real, imag} */,
  {32'hbdcb70e8, 32'hc073c605} /* (2, 19, 10) {real, imag} */,
  {32'h3fe16f16, 32'hc14fba21} /* (2, 19, 9) {real, imag} */,
  {32'h4092e571, 32'hc13267da} /* (2, 19, 8) {real, imag} */,
  {32'h3fd9debe, 32'hc1693aad} /* (2, 19, 7) {real, imag} */,
  {32'hbfad3ff2, 32'hc13d0892} /* (2, 19, 6) {real, imag} */,
  {32'h40372dd4, 32'hc174a9ba} /* (2, 19, 5) {real, imag} */,
  {32'h407e83a6, 32'hc179e1c2} /* (2, 19, 4) {real, imag} */,
  {32'h40a2e9be, 32'hc14ace70} /* (2, 19, 3) {real, imag} */,
  {32'h40c20f1e, 32'hc1704afd} /* (2, 19, 2) {real, imag} */,
  {32'h40a1dfbe, 32'hc163832c} /* (2, 19, 1) {real, imag} */,
  {32'h400e5635, 32'hc102e9fd} /* (2, 19, 0) {real, imag} */,
  {32'h3fa5a41c, 32'hc10501aa} /* (2, 18, 31) {real, imag} */,
  {32'h40814c8c, 32'hc172b0be} /* (2, 18, 30) {real, imag} */,
  {32'h4024b6ae, 32'hc16cbab6} /* (2, 18, 29) {real, imag} */,
  {32'h40266029, 32'hc1722c34} /* (2, 18, 28) {real, imag} */,
  {32'h407dcd86, 32'hc15017c6} /* (2, 18, 27) {real, imag} */,
  {32'h40922adb, 32'hc1426b3e} /* (2, 18, 26) {real, imag} */,
  {32'h40a40cb2, 32'hc13ee2da} /* (2, 18, 25) {real, imag} */,
  {32'h41190b2c, 32'hc16356c6} /* (2, 18, 24) {real, imag} */,
  {32'h40c2fc05, 32'hc18047e0} /* (2, 18, 23) {real, imag} */,
  {32'h4005ec80, 32'hc16354fa} /* (2, 18, 22) {real, imag} */,
  {32'hbeb018db, 32'hc0fadd75} /* (2, 18, 21) {real, imag} */,
  {32'hc073d2ee, 32'h41013cf8} /* (2, 18, 20) {real, imag} */,
  {32'hbfbfeece, 32'h4152e299} /* (2, 18, 19) {real, imag} */,
  {32'hbdcbdbd8, 32'h416f3f34} /* (2, 18, 18) {real, imag} */,
  {32'hc09f2374, 32'h4145ce40} /* (2, 18, 17) {real, imag} */,
  {32'hc0b7a824, 32'h4166b24e} /* (2, 18, 16) {real, imag} */,
  {32'hc0aca078, 32'h417b1dc9} /* (2, 18, 15) {real, imag} */,
  {32'hc0852ae8, 32'h4159a55c} /* (2, 18, 14) {real, imag} */,
  {32'hc062f5e6, 32'h416cadb4} /* (2, 18, 13) {real, imag} */,
  {32'hbff2b08f, 32'h417693db} /* (2, 18, 12) {real, imag} */,
  {32'hbff0ab29, 32'h416dd0b0} /* (2, 18, 11) {real, imag} */,
  {32'h3fcb31ec, 32'hc0918978} /* (2, 18, 10) {real, imag} */,
  {32'h400dc286, 32'hc15a929f} /* (2, 18, 9) {real, imag} */,
  {32'h4056c8f2, 32'hc1663c58} /* (2, 18, 8) {real, imag} */,
  {32'h3ffd7706, 32'hc180cee0} /* (2, 18, 7) {real, imag} */,
  {32'h3e6e1524, 32'hc1705960} /* (2, 18, 6) {real, imag} */,
  {32'h3ff2937e, 32'hc184bb00} /* (2, 18, 5) {real, imag} */,
  {32'h40b3f756, 32'hc17a704e} /* (2, 18, 4) {real, imag} */,
  {32'h40c5b7b4, 32'hc1472763} /* (2, 18, 3) {real, imag} */,
  {32'h408704aa, 32'hc1449405} /* (2, 18, 2) {real, imag} */,
  {32'h4026e35c, 32'hc16e585a} /* (2, 18, 1) {real, imag} */,
  {32'h402c61de, 32'hc121d978} /* (2, 18, 0) {real, imag} */,
  {32'h40248ce2, 32'hc0d929f2} /* (2, 17, 31) {real, imag} */,
  {32'h40c7ac8c, 32'hc166da44} /* (2, 17, 30) {real, imag} */,
  {32'h408dcdb4, 32'hc177a93a} /* (2, 17, 29) {real, imag} */,
  {32'h408bb4cd, 32'hc182159c} /* (2, 17, 28) {real, imag} */,
  {32'h4083947e, 32'hc181bc46} /* (2, 17, 27) {real, imag} */,
  {32'h405bc536, 32'hc157e101} /* (2, 17, 26) {real, imag} */,
  {32'h40837c7a, 32'hc14fad3a} /* (2, 17, 25) {real, imag} */,
  {32'h40c38844, 32'hc160dae1} /* (2, 17, 24) {real, imag} */,
  {32'h4089882e, 32'hc1950560} /* (2, 17, 23) {real, imag} */,
  {32'h4022a194, 32'hc173139d} /* (2, 17, 22) {real, imag} */,
  {32'h3ea8ff22, 32'hc0e6dbd4} /* (2, 17, 21) {real, imag} */,
  {32'hbfb1765e, 32'h41039cd4} /* (2, 17, 20) {real, imag} */,
  {32'hbf36ef18, 32'h4167e81c} /* (2, 17, 19) {real, imag} */,
  {32'hbfa53181, 32'h418445c7} /* (2, 17, 18) {real, imag} */,
  {32'hc0947edc, 32'h4180a4d6} /* (2, 17, 17) {real, imag} */,
  {32'hc098db82, 32'h416d57a6} /* (2, 17, 16) {real, imag} */,
  {32'hc07982a1, 32'h4155e8ec} /* (2, 17, 15) {real, imag} */,
  {32'hc0507893, 32'h41458740} /* (2, 17, 14) {real, imag} */,
  {32'hc04647c0, 32'h412eeefa} /* (2, 17, 13) {real, imag} */,
  {32'hbff1a5c1, 32'h4152ddf5} /* (2, 17, 12) {real, imag} */,
  {32'h3e87ed8c, 32'h4139f290} /* (2, 17, 11) {real, imag} */,
  {32'h4097d742, 32'hc0c4ef6c} /* (2, 17, 10) {real, imag} */,
  {32'h40913a58, 32'hc141e8ca} /* (2, 17, 9) {real, imag} */,
  {32'h40730958, 32'hc162d3f4} /* (2, 17, 8) {real, imag} */,
  {32'h3fdc9c43, 32'hc14a3b46} /* (2, 17, 7) {real, imag} */,
  {32'h40305274, 32'hc17fedb2} /* (2, 17, 6) {real, imag} */,
  {32'h3fce0918, 32'hc18631ae} /* (2, 17, 5) {real, imag} */,
  {32'h405b41b4, 32'hc18aaa95} /* (2, 17, 4) {real, imag} */,
  {32'h40bc7e0a, 32'hc181bfe0} /* (2, 17, 3) {real, imag} */,
  {32'h407f6122, 32'hc17ca7c6} /* (2, 17, 2) {real, imag} */,
  {32'hbf21b2a8, 32'hc16a4c1e} /* (2, 17, 1) {real, imag} */,
  {32'h3e614880, 32'hc0ff8926} /* (2, 17, 0) {real, imag} */,
  {32'h3f7c2d8c, 32'hc0fcb814} /* (2, 16, 31) {real, imag} */,
  {32'h407702ad, 32'hc175ea4c} /* (2, 16, 30) {real, imag} */,
  {32'h40810b34, 32'hc160bd5a} /* (2, 16, 29) {real, imag} */,
  {32'h40c5ac54, 32'hc1502a26} /* (2, 16, 28) {real, imag} */,
  {32'h40c06b03, 32'hc179dd76} /* (2, 16, 27) {real, imag} */,
  {32'h4036de60, 32'hc16d4cfe} /* (2, 16, 26) {real, imag} */,
  {32'h400c4e65, 32'hc1817538} /* (2, 16, 25) {real, imag} */,
  {32'h3f919e17, 32'hc187970c} /* (2, 16, 24) {real, imag} */,
  {32'h3eb64abe, 32'hc190ac72} /* (2, 16, 23) {real, imag} */,
  {32'h401befb1, 32'hc1681114} /* (2, 16, 22) {real, imag} */,
  {32'h3fce5eec, 32'hc07747fd} /* (2, 16, 21) {real, imag} */,
  {32'hbf7b9aa6, 32'h41601302} /* (2, 16, 20) {real, imag} */,
  {32'hc00ed286, 32'h41861d00} /* (2, 16, 19) {real, imag} */,
  {32'hc0480112, 32'h4179eaa7} /* (2, 16, 18) {real, imag} */,
  {32'hc09eaddb, 32'h417b662e} /* (2, 16, 17) {real, imag} */,
  {32'hc09831da, 32'h4183e67a} /* (2, 16, 16) {real, imag} */,
  {32'hc0bdb1ce, 32'h416f0c4e} /* (2, 16, 15) {real, imag} */,
  {32'hc0927377, 32'h413e02de} /* (2, 16, 14) {real, imag} */,
  {32'hc0777918, 32'h4163cc96} /* (2, 16, 13) {real, imag} */,
  {32'hbfe48bed, 32'h41812aa5} /* (2, 16, 12) {real, imag} */,
  {32'h3eb407aa, 32'h4138dacd} /* (2, 16, 11) {real, imag} */,
  {32'h407e1018, 32'hc0c771c2} /* (2, 16, 10) {real, imag} */,
  {32'h40b8dc94, 32'hc163d402} /* (2, 16, 9) {real, imag} */,
  {32'h40c5c3b8, 32'hc1693a3c} /* (2, 16, 8) {real, imag} */,
  {32'h40129c5b, 32'hc14863e4} /* (2, 16, 7) {real, imag} */,
  {32'hbf4872ac, 32'hc13eb3ec} /* (2, 16, 6) {real, imag} */,
  {32'hbfcdfb54, 32'hc15bfd55} /* (2, 16, 5) {real, imag} */,
  {32'hbe611498, 32'hc164ffac} /* (2, 16, 4) {real, imag} */,
  {32'h40828ce3, 32'hc172c833} /* (2, 16, 3) {real, imag} */,
  {32'h4092307a, 32'hc15bab00} /* (2, 16, 2) {real, imag} */,
  {32'h401b47ec, 32'hc156d3b2} /* (2, 16, 1) {real, imag} */,
  {32'h3eb0b51b, 32'hc0f9a560} /* (2, 16, 0) {real, imag} */,
  {32'h3f6df2ed, 32'hc114d7a6} /* (2, 15, 31) {real, imag} */,
  {32'h4036884a, 32'hc18c1504} /* (2, 15, 30) {real, imag} */,
  {32'h4072cd34, 32'hc1858f04} /* (2, 15, 29) {real, imag} */,
  {32'h4069061e, 32'hc1603b09} /* (2, 15, 28) {real, imag} */,
  {32'h40973be0, 32'hc15f2bca} /* (2, 15, 27) {real, imag} */,
  {32'h4083aef2, 32'hc183b880} /* (2, 15, 26) {real, imag} */,
  {32'h40751733, 32'hc178aec2} /* (2, 15, 25) {real, imag} */,
  {32'h4034e0ac, 32'hc15f051a} /* (2, 15, 24) {real, imag} */,
  {32'hbdd3c05c, 32'hc1787658} /* (2, 15, 23) {real, imag} */,
  {32'h40880f95, 32'hc16fb11b} /* (2, 15, 22) {real, imag} */,
  {32'h401ba26c, 32'hc07aafe0} /* (2, 15, 21) {real, imag} */,
  {32'hc013894c, 32'h4138d42b} /* (2, 15, 20) {real, imag} */,
  {32'hbfbafdd9, 32'h4150d61c} /* (2, 15, 19) {real, imag} */,
  {32'hc0089aae, 32'h414c0378} /* (2, 15, 18) {real, imag} */,
  {32'hc06f5296, 32'h4144a71c} /* (2, 15, 17) {real, imag} */,
  {32'hc055b716, 32'h4154e291} /* (2, 15, 16) {real, imag} */,
  {32'hc05ab234, 32'h4172efd0} /* (2, 15, 15) {real, imag} */,
  {32'hc043a42e, 32'h41437a6f} /* (2, 15, 14) {real, imag} */,
  {32'hc079482c, 32'h417e6541} /* (2, 15, 13) {real, imag} */,
  {32'hc0718df9, 32'h4191cb4a} /* (2, 15, 12) {real, imag} */,
  {32'hbffb4c58, 32'h415f6e78} /* (2, 15, 11) {real, imag} */,
  {32'h403e79be, 32'hc0ad9adc} /* (2, 15, 10) {real, imag} */,
  {32'h40b7e82b, 32'hc16bea90} /* (2, 15, 9) {real, imag} */,
  {32'h40b60bbe, 32'hc181cdae} /* (2, 15, 8) {real, imag} */,
  {32'h40a7dea2, 32'hc18bf8f3} /* (2, 15, 7) {real, imag} */,
  {32'h3fcc2f29, 32'hc15ed9e4} /* (2, 15, 6) {real, imag} */,
  {32'hbe054b14, 32'hc166313f} /* (2, 15, 5) {real, imag} */,
  {32'h404f8163, 32'hc1698046} /* (2, 15, 4) {real, imag} */,
  {32'h40a36b83, 32'hc16b87a4} /* (2, 15, 3) {real, imag} */,
  {32'h40d59c49, 32'hc14cdf3d} /* (2, 15, 2) {real, imag} */,
  {32'h40b3d0a8, 32'hc16e9026} /* (2, 15, 1) {real, imag} */,
  {32'h3fe8591a, 32'hc115ed41} /* (2, 15, 0) {real, imag} */,
  {32'h3f2e44b8, 32'hc10ccc4a} /* (2, 14, 31) {real, imag} */,
  {32'h40045784, 32'hc184a7c2} /* (2, 14, 30) {real, imag} */,
  {32'h3fdba09b, 32'hc18e7b40} /* (2, 14, 29) {real, imag} */,
  {32'h40080326, 32'hc1834504} /* (2, 14, 28) {real, imag} */,
  {32'h406aa9b8, 32'hc15e4ce4} /* (2, 14, 27) {real, imag} */,
  {32'h408a549e, 32'hc1569b14} /* (2, 14, 26) {real, imag} */,
  {32'h40891db7, 32'hc147824e} /* (2, 14, 25) {real, imag} */,
  {32'h3f81df8e, 32'hc14c4068} /* (2, 14, 24) {real, imag} */,
  {32'h3f1a00a8, 32'hc16132a4} /* (2, 14, 23) {real, imag} */,
  {32'h40aa0708, 32'hc186f8d2} /* (2, 14, 22) {real, imag} */,
  {32'h4069b2c2, 32'hc0f22889} /* (2, 14, 21) {real, imag} */,
  {32'hbfeffc48, 32'h412ba3e5} /* (2, 14, 20) {real, imag} */,
  {32'hc067685c, 32'h4151e210} /* (2, 14, 19) {real, imag} */,
  {32'hc0413113, 32'h4146cb30} /* (2, 14, 18) {real, imag} */,
  {32'hbfadba1b, 32'h4157617f} /* (2, 14, 17) {real, imag} */,
  {32'hbe407ed2, 32'h415c0017} /* (2, 14, 16) {real, imag} */,
  {32'hbf825958, 32'h41759822} /* (2, 14, 15) {real, imag} */,
  {32'hc09baae3, 32'h4159ac36} /* (2, 14, 14) {real, imag} */,
  {32'hc0a0cb84, 32'h4159cd9f} /* (2, 14, 13) {real, imag} */,
  {32'hc04dac30, 32'h4168f73c} /* (2, 14, 12) {real, imag} */,
  {32'hbf03ff20, 32'h41438bdd} /* (2, 14, 11) {real, imag} */,
  {32'h4051db1e, 32'hc039987c} /* (2, 14, 10) {real, imag} */,
  {32'h40a3c585, 32'hc161c732} /* (2, 14, 9) {real, imag} */,
  {32'h4049b4ff, 32'hc1886413} /* (2, 14, 8) {real, imag} */,
  {32'h403b4157, 32'hc184963a} /* (2, 14, 7) {real, imag} */,
  {32'h3fb9d12a, 32'hc14d94cc} /* (2, 14, 6) {real, imag} */,
  {32'h3d7d6c00, 32'hc137ceb8} /* (2, 14, 5) {real, imag} */,
  {32'h3fbbdefb, 32'hc12f265c} /* (2, 14, 4) {real, imag} */,
  {32'h40832c30, 32'hc141c34d} /* (2, 14, 3) {real, imag} */,
  {32'h40d1915e, 32'hc1529554} /* (2, 14, 2) {real, imag} */,
  {32'h409c5a0e, 32'hc1885cfe} /* (2, 14, 1) {real, imag} */,
  {32'h3edf19b8, 32'hc1324645} /* (2, 14, 0) {real, imag} */,
  {32'h3f7230b0, 32'hc107254e} /* (2, 13, 31) {real, imag} */,
  {32'h404a2108, 32'hc17f7f5c} /* (2, 13, 30) {real, imag} */,
  {32'h408e5b3c, 32'hc18bd9a4} /* (2, 13, 29) {real, imag} */,
  {32'h4032ad42, 32'hc18fb20c} /* (2, 13, 28) {real, imag} */,
  {32'h3f1be061, 32'hc15ec1e2} /* (2, 13, 27) {real, imag} */,
  {32'h407be294, 32'hc13d5c26} /* (2, 13, 26) {real, imag} */,
  {32'h40a7fcdb, 32'hc13a4b45} /* (2, 13, 25) {real, imag} */,
  {32'h3f9519e2, 32'hc14d8f06} /* (2, 13, 24) {real, imag} */,
  {32'h3e0cb07c, 32'hc1450bb4} /* (2, 13, 23) {real, imag} */,
  {32'h4027dcce, 32'hc1891bf4} /* (2, 13, 22) {real, imag} */,
  {32'h3e22f6b0, 32'hc116bf44} /* (2, 13, 21) {real, imag} */,
  {32'hc04bcfd2, 32'h41297bc2} /* (2, 13, 20) {real, imag} */,
  {32'hc0054a34, 32'h418774f8} /* (2, 13, 19) {real, imag} */,
  {32'hc0100e5c, 32'h416cff8a} /* (2, 13, 18) {real, imag} */,
  {32'hc043ccb0, 32'h4172c18e} /* (2, 13, 17) {real, imag} */,
  {32'hc041f0ef, 32'h41485542} /* (2, 13, 16) {real, imag} */,
  {32'hbfd1108f, 32'h4132762e} /* (2, 13, 15) {real, imag} */,
  {32'hc03ec7bf, 32'h415bda37} /* (2, 13, 14) {real, imag} */,
  {32'hc03f66d0, 32'h415505fa} /* (2, 13, 13) {real, imag} */,
  {32'hbfdc1127, 32'h4145e167} /* (2, 13, 12) {real, imag} */,
  {32'hbf9b7a30, 32'h412b2d48} /* (2, 13, 11) {real, imag} */,
  {32'h3ffd092c, 32'hc0848cf6} /* (2, 13, 10) {real, imag} */,
  {32'h40a067e0, 32'hc1475582} /* (2, 13, 9) {real, imag} */,
  {32'h4014f1c8, 32'hc1862f5e} /* (2, 13, 8) {real, imag} */,
  {32'h4006b3fc, 32'hc183adfe} /* (2, 13, 7) {real, imag} */,
  {32'h3e8346f4, 32'hc143fc1b} /* (2, 13, 6) {real, imag} */,
  {32'hbe1ab5d4, 32'hc12ec3b0} /* (2, 13, 5) {real, imag} */,
  {32'hbed16703, 32'hc10d597c} /* (2, 13, 4) {real, imag} */,
  {32'h408f5434, 32'hc12d37e0} /* (2, 13, 3) {real, imag} */,
  {32'h40c2bf2d, 32'hc14d20a5} /* (2, 13, 2) {real, imag} */,
  {32'h408673f7, 32'hc184ef24} /* (2, 13, 1) {real, imag} */,
  {32'h3f5c4113, 32'hc130b131} /* (2, 13, 0) {real, imag} */,
  {32'hbe777d66, 32'hc0eee60e} /* (2, 12, 31) {real, imag} */,
  {32'h3faf8b52, 32'hc15e1a63} /* (2, 12, 30) {real, imag} */,
  {32'h4079a5bf, 32'hc163fce6} /* (2, 12, 29) {real, imag} */,
  {32'h40583f1b, 32'hc1809afb} /* (2, 12, 28) {real, imag} */,
  {32'h3fd6a3ee, 32'hc162ee44} /* (2, 12, 27) {real, imag} */,
  {32'h4050e364, 32'hc12883b4} /* (2, 12, 26) {real, imag} */,
  {32'h40c444ac, 32'hc1258680} /* (2, 12, 25) {real, imag} */,
  {32'h409ec35d, 32'hc14bc10e} /* (2, 12, 24) {real, imag} */,
  {32'h4041d396, 32'hc167d02c} /* (2, 12, 23) {real, imag} */,
  {32'h3fbd3f7e, 32'hc190366e} /* (2, 12, 22) {real, imag} */,
  {32'h4018452c, 32'hc1006618} /* (2, 12, 21) {real, imag} */,
  {32'hbf475efa, 32'h4123411c} /* (2, 12, 20) {real, imag} */,
  {32'h3faa49dc, 32'h419c9c8a} /* (2, 12, 19) {real, imag} */,
  {32'h403d405c, 32'h41861e3a} /* (2, 12, 18) {real, imag} */,
  {32'hbeb2c9e8, 32'h4187b7ec} /* (2, 12, 17) {real, imag} */,
  {32'hc06e02c8, 32'h416e0364} /* (2, 12, 16) {real, imag} */,
  {32'hc08dd4d7, 32'h4137356e} /* (2, 12, 15) {real, imag} */,
  {32'hc085a03e, 32'h41683f1c} /* (2, 12, 14) {real, imag} */,
  {32'hbf9e9ace, 32'h4156373a} /* (2, 12, 13) {real, imag} */,
  {32'h3e69f514, 32'h41303cd1} /* (2, 12, 12) {real, imag} */,
  {32'h3fcf2f5a, 32'h4111f349} /* (2, 12, 11) {real, imag} */,
  {32'hbde92edc, 32'hc0eb70a4} /* (2, 12, 10) {real, imag} */,
  {32'h402734b4, 32'hc14ec5fe} /* (2, 12, 9) {real, imag} */,
  {32'h3f3cf854, 32'hc162eaef} /* (2, 12, 8) {real, imag} */,
  {32'h4062e213, 32'hc18054e0} /* (2, 12, 7) {real, imag} */,
  {32'h408950fe, 32'hc1670ac4} /* (2, 12, 6) {real, imag} */,
  {32'h402bbbd0, 32'hc15416eb} /* (2, 12, 5) {real, imag} */,
  {32'h40106ac1, 32'hc142474e} /* (2, 12, 4) {real, imag} */,
  {32'h403e7cf2, 32'hc174083c} /* (2, 12, 3) {real, imag} */,
  {32'h400f836c, 32'hc170f980} /* (2, 12, 2) {real, imag} */,
  {32'h40110265, 32'hc18b031e} /* (2, 12, 1) {real, imag} */,
  {32'h3f9177ae, 32'hc1097857} /* (2, 12, 0) {real, imag} */,
  {32'h3e5eee54, 32'hc095946a} /* (2, 11, 31) {real, imag} */,
  {32'h3ee96381, 32'hc10c50a8} /* (2, 11, 30) {real, imag} */,
  {32'h3fde0ba0, 32'hc10c3f93} /* (2, 11, 29) {real, imag} */,
  {32'h3fd489d4, 32'hc14d8e01} /* (2, 11, 28) {real, imag} */,
  {32'h3fadbb6c, 32'hc12b531c} /* (2, 11, 27) {real, imag} */,
  {32'hbf518947, 32'hc10c4d49} /* (2, 11, 26) {real, imag} */,
  {32'h3fd0443a, 32'hc10b1500} /* (2, 11, 25) {real, imag} */,
  {32'h3fdddfee, 32'hc11fd9ec} /* (2, 11, 24) {real, imag} */,
  {32'hbfa47d48, 32'hc1365fce} /* (2, 11, 23) {real, imag} */,
  {32'hbfabfee8, 32'hc135757c} /* (2, 11, 22) {real, imag} */,
  {32'h406f449a, 32'hc0550988} /* (2, 11, 21) {real, imag} */,
  {32'h3e967070, 32'h40e9d56c} /* (2, 11, 20) {real, imag} */,
  {32'h3e311f45, 32'h414983bd} /* (2, 11, 19) {real, imag} */,
  {32'h3f76c4c3, 32'h41437e86} /* (2, 11, 18) {real, imag} */,
  {32'h3fa7230a, 32'h41702826} /* (2, 11, 17) {real, imag} */,
  {32'hc02b0c6a, 32'h4145d38d} /* (2, 11, 16) {real, imag} */,
  {32'hc09dc27e, 32'h41256b5c} /* (2, 11, 15) {real, imag} */,
  {32'hc083f2ce, 32'h4140f63a} /* (2, 11, 14) {real, imag} */,
  {32'hc01a5e88, 32'h4140413e} /* (2, 11, 13) {real, imag} */,
  {32'hbfe8c569, 32'h41202157} /* (2, 11, 12) {real, imag} */,
  {32'h3f0b5df5, 32'h40bac488} /* (2, 11, 11) {real, imag} */,
  {32'h3f2370b1, 32'hc1084442} /* (2, 11, 10) {real, imag} */,
  {32'h3f615a6f, 32'hc131839b} /* (2, 11, 9) {real, imag} */,
  {32'h3f9c303c, 32'hc11e3a32} /* (2, 11, 8) {real, imag} */,
  {32'hbe5b2dda, 32'hc14207d2} /* (2, 11, 7) {real, imag} */,
  {32'h408f0f0a, 32'hc1483840} /* (2, 11, 6) {real, imag} */,
  {32'h40aa971f, 32'hc106830f} /* (2, 11, 5) {real, imag} */,
  {32'h402e15e9, 32'hc102ec99} /* (2, 11, 4) {real, imag} */,
  {32'h3fe80430, 32'hc1378e16} /* (2, 11, 3) {real, imag} */,
  {32'h4039670c, 32'hc127817a} /* (2, 11, 2) {real, imag} */,
  {32'h4054e744, 32'hc1383d49} /* (2, 11, 1) {real, imag} */,
  {32'h3f65b1e5, 32'hc0c086d3} /* (2, 11, 0) {real, imag} */,
  {32'hbd6ce0f4, 32'h40bc47ec} /* (2, 10, 31) {real, imag} */,
  {32'h3dd04e50, 32'h40e4bcec} /* (2, 10, 30) {real, imag} */,
  {32'h3fd2bf4f, 32'h40ed4cae} /* (2, 10, 29) {real, imag} */,
  {32'hbf816082, 32'h40e14596} /* (2, 10, 28) {real, imag} */,
  {32'hc0629b4b, 32'h41084f32} /* (2, 10, 27) {real, imag} */,
  {32'hc076035f, 32'h40d9335a} /* (2, 10, 26) {real, imag} */,
  {32'hc016b34b, 32'h40b8da0a} /* (2, 10, 25) {real, imag} */,
  {32'hc058ee37, 32'h40f8ffc1} /* (2, 10, 24) {real, imag} */,
  {32'hc08bbbc8, 32'h40dbd30d} /* (2, 10, 23) {real, imag} */,
  {32'hc02591a7, 32'h41050b4d} /* (2, 10, 22) {real, imag} */,
  {32'hbf8602ef, 32'h4099445a} /* (2, 10, 21) {real, imag} */,
  {32'hbef103af, 32'hc0950036} /* (2, 10, 20) {real, imag} */,
  {32'h3f9756f0, 32'hc0e36416} /* (2, 10, 19) {real, imag} */,
  {32'h400d5dbe, 32'hc0a9a037} /* (2, 10, 18) {real, imag} */,
  {32'h3fe795b8, 32'hc04ccd0a} /* (2, 10, 17) {real, imag} */,
  {32'h3f8cd445, 32'hc0c1ba76} /* (2, 10, 16) {real, imag} */,
  {32'hbf91b779, 32'hc0d4e461} /* (2, 10, 15) {real, imag} */,
  {32'hbeb9e4f6, 32'hc07189a4} /* (2, 10, 14) {real, imag} */,
  {32'h3f76ad58, 32'hc067c845} /* (2, 10, 13) {real, imag} */,
  {32'h3fdc2cbe, 32'hc0e4dbb6} /* (2, 10, 12) {real, imag} */,
  {32'h401b9282, 32'hc0d78261} /* (2, 10, 11) {real, imag} */,
  {32'h3f334d67, 32'hbeca6a65} /* (2, 10, 10) {real, imag} */,
  {32'hc000f4cd, 32'h40b4495a} /* (2, 10, 9) {real, imag} */,
  {32'hbfa3cf0f, 32'h40ae12c2} /* (2, 10, 8) {real, imag} */,
  {32'hc0baa72c, 32'h40d6461b} /* (2, 10, 7) {real, imag} */,
  {32'hbf85b150, 32'h40fe01d1} /* (2, 10, 6) {real, imag} */,
  {32'hbf6c6867, 32'h4117857b} /* (2, 10, 5) {real, imag} */,
  {32'hbb09b800, 32'h4119ef8a} /* (2, 10, 4) {real, imag} */,
  {32'h40459a6a, 32'h40cf786c} /* (2, 10, 3) {real, imag} */,
  {32'h3fe8ac23, 32'h40e331e6} /* (2, 10, 2) {real, imag} */,
  {32'hbebbf837, 32'h40f0147a} /* (2, 10, 1) {real, imag} */,
  {32'hbfcdabb4, 32'h40c83a28} /* (2, 10, 0) {real, imag} */,
  {32'hc0254c98, 32'h410c36b4} /* (2, 9, 31) {real, imag} */,
  {32'hc055f853, 32'h4165e18a} /* (2, 9, 30) {real, imag} */,
  {32'hbf59642c, 32'h41806803} /* (2, 9, 29) {real, imag} */,
  {32'hc01a0926, 32'h418debe0} /* (2, 9, 28) {real, imag} */,
  {32'hc03473d5, 32'h416c75eb} /* (2, 9, 27) {real, imag} */,
  {32'hbfa881b4, 32'h415b6a70} /* (2, 9, 26) {real, imag} */,
  {32'hc0338633, 32'h4140c15a} /* (2, 9, 25) {real, imag} */,
  {32'hc00f0674, 32'h41739bd6} /* (2, 9, 24) {real, imag} */,
  {32'hc086cf16, 32'h414e38d4} /* (2, 9, 23) {real, imag} */,
  {32'hc0a67042, 32'h415c31f6} /* (2, 9, 22) {real, imag} */,
  {32'hc0307e90, 32'h410ec7ac} /* (2, 9, 21) {real, imag} */,
  {32'hbeb9ecb0, 32'hc0f17206} /* (2, 9, 20) {real, imag} */,
  {32'h404325bb, 32'hc1491124} /* (2, 9, 19) {real, imag} */,
  {32'h40283b6e, 32'hc15dbd00} /* (2, 9, 18) {real, imag} */,
  {32'h405086ea, 32'hc15f022e} /* (2, 9, 17) {real, imag} */,
  {32'h40918270, 32'hc1863786} /* (2, 9, 16) {real, imag} */,
  {32'h407b73f8, 32'hc197f9e5} /* (2, 9, 15) {real, imag} */,
  {32'h3fea1e35, 32'hc15d5ae2} /* (2, 9, 14) {real, imag} */,
  {32'h4058b657, 32'hc12ec9ba} /* (2, 9, 13) {real, imag} */,
  {32'h406460e6, 32'hc1783314} /* (2, 9, 12) {real, imag} */,
  {32'h40257886, 32'hc13f68c8} /* (2, 9, 11) {real, imag} */,
  {32'hbee81c51, 32'h40c0bcee} /* (2, 9, 10) {real, imag} */,
  {32'hc02617ac, 32'h417a4a8a} /* (2, 9, 9) {real, imag} */,
  {32'hc031d668, 32'h41541c9f} /* (2, 9, 8) {real, imag} */,
  {32'hc0991bec, 32'h41413ba8} /* (2, 9, 7) {real, imag} */,
  {32'hbfab6dd5, 32'h41596413} /* (2, 9, 6) {real, imag} */,
  {32'hc0260c18, 32'h416a5b05} /* (2, 9, 5) {real, imag} */,
  {32'hbfba99db, 32'h4181c03c} /* (2, 9, 4) {real, imag} */,
  {32'h3f7a21c5, 32'h41741581} /* (2, 9, 3) {real, imag} */,
  {32'hbf7047f4, 32'h414dcea1} /* (2, 9, 2) {real, imag} */,
  {32'hbfec943e, 32'h4150720d} /* (2, 9, 1) {real, imag} */,
  {32'hc010b2bb, 32'h410e086b} /* (2, 9, 0) {real, imag} */,
  {32'hc05be5bb, 32'h41000b0e} /* (2, 8, 31) {real, imag} */,
  {32'hc040bfb1, 32'h415a4770} /* (2, 8, 30) {real, imag} */,
  {32'hbff7fce6, 32'h41790fc2} /* (2, 8, 29) {real, imag} */,
  {32'hbfcabbe1, 32'h4178df1a} /* (2, 8, 28) {real, imag} */,
  {32'hc022a408, 32'h417958a8} /* (2, 8, 27) {real, imag} */,
  {32'hbff25a4f, 32'h418980db} /* (2, 8, 26) {real, imag} */,
  {32'hbd735550, 32'h415c9464} /* (2, 8, 25) {real, imag} */,
  {32'h3dc1ac48, 32'h4167d216} /* (2, 8, 24) {real, imag} */,
  {32'hc09956fc, 32'h4152896d} /* (2, 8, 23) {real, imag} */,
  {32'hc09388b6, 32'h4165d60d} /* (2, 8, 22) {real, imag} */,
  {32'h3edba324, 32'h4100fd68} /* (2, 8, 21) {real, imag} */,
  {32'hbeb9f780, 32'hc1064036} /* (2, 8, 20) {real, imag} */,
  {32'h40087b96, 32'hc155f265} /* (2, 8, 19) {real, imag} */,
  {32'h403cea72, 32'hc17052ae} /* (2, 8, 18) {real, imag} */,
  {32'h40893214, 32'hc158f286} /* (2, 8, 17) {real, imag} */,
  {32'h40c0f56e, 32'hc159bf23} /* (2, 8, 16) {real, imag} */,
  {32'h4079008b, 32'hc19a2c71} /* (2, 8, 15) {real, imag} */,
  {32'h4052b547, 32'hc17b2e80} /* (2, 8, 14) {real, imag} */,
  {32'h3fd9774a, 32'hc1150dc6} /* (2, 8, 13) {real, imag} */,
  {32'hbda93f24, 32'hc16312cc} /* (2, 8, 12) {real, imag} */,
  {32'hbe4ce4a8, 32'hc1541082} /* (2, 8, 11) {real, imag} */,
  {32'hc0837890, 32'h40bd6183} /* (2, 8, 10) {real, imag} */,
  {32'hc08c04a6, 32'h4171190b} /* (2, 8, 9) {real, imag} */,
  {32'hc022e856, 32'h414f2f86} /* (2, 8, 8) {real, imag} */,
  {32'hbf873892, 32'h413a8d5c} /* (2, 8, 7) {real, imag} */,
  {32'h3e4fd640, 32'h4165bc08} /* (2, 8, 6) {real, imag} */,
  {32'hc008059a, 32'h416217f5} /* (2, 8, 5) {real, imag} */,
  {32'hc093fea0, 32'h4165e434} /* (2, 8, 4) {real, imag} */,
  {32'hc012d35d, 32'h416119d0} /* (2, 8, 3) {real, imag} */,
  {32'hc01d5a19, 32'h4151828d} /* (2, 8, 2) {real, imag} */,
  {32'hc02a57cc, 32'h414d8cf0} /* (2, 8, 1) {real, imag} */,
  {32'hc05e6fa0, 32'h40cfb576} /* (2, 8, 0) {real, imag} */,
  {32'hc0353c1a, 32'h40f38f3d} /* (2, 7, 31) {real, imag} */,
  {32'hc0345b08, 32'h413fa5b9} /* (2, 7, 30) {real, imag} */,
  {32'hc0286922, 32'h415b2d8a} /* (2, 7, 29) {real, imag} */,
  {32'hbf71d983, 32'h41435194} /* (2, 7, 28) {real, imag} */,
  {32'hc04135ca, 32'h4161c90e} /* (2, 7, 27) {real, imag} */,
  {32'hc0795b88, 32'h418c8cca} /* (2, 7, 26) {real, imag} */,
  {32'hc003891c, 32'h418f69e6} /* (2, 7, 25) {real, imag} */,
  {32'hc05623f9, 32'h41898c53} /* (2, 7, 24) {real, imag} */,
  {32'hc0725166, 32'h414a8ca3} /* (2, 7, 23) {real, imag} */,
  {32'hc065d886, 32'h4159823a} /* (2, 7, 22) {real, imag} */,
  {32'hc072ad98, 32'h4109f6be} /* (2, 7, 21) {real, imag} */,
  {32'hc02754a4, 32'hc12e9ab1} /* (2, 7, 20) {real, imag} */,
  {32'h3fa35d6d, 32'hc1718477} /* (2, 7, 19) {real, imag} */,
  {32'h409a2e72, 32'hc175247f} /* (2, 7, 18) {real, imag} */,
  {32'h40b79a3a, 32'hc1844084} /* (2, 7, 17) {real, imag} */,
  {32'h40af33e0, 32'hc1698897} /* (2, 7, 16) {real, imag} */,
  {32'h40c4f368, 32'hc17bb7f9} /* (2, 7, 15) {real, imag} */,
  {32'h40c373fb, 32'hc1676f5f} /* (2, 7, 14) {real, imag} */,
  {32'h408f0756, 32'hc1196658} /* (2, 7, 13) {real, imag} */,
  {32'h406e733e, 32'hc15b6c08} /* (2, 7, 12) {real, imag} */,
  {32'h404b71b0, 32'hc13f5ea7} /* (2, 7, 11) {real, imag} */,
  {32'hc0171887, 32'h40b29a24} /* (2, 7, 10) {real, imag} */,
  {32'hc0a1a356, 32'h4138ed86} /* (2, 7, 9) {real, imag} */,
  {32'hc04f7fa0, 32'h413fe5b8} /* (2, 7, 8) {real, imag} */,
  {32'hbfc9fad6, 32'h41689ef8} /* (2, 7, 7) {real, imag} */,
  {32'hc00ef2a4, 32'h41806acc} /* (2, 7, 6) {real, imag} */,
  {32'hbff03aa7, 32'h418a161f} /* (2, 7, 5) {real, imag} */,
  {32'hc0ad888c, 32'h4192d084} /* (2, 7, 4) {real, imag} */,
  {32'hc0829f18, 32'h41821926} /* (2, 7, 3) {real, imag} */,
  {32'hc016433a, 32'h416de660} /* (2, 7, 2) {real, imag} */,
  {32'hc0377c56, 32'h41446287} /* (2, 7, 1) {real, imag} */,
  {32'hbffd5208, 32'h40b240bb} /* (2, 7, 0) {real, imag} */,
  {32'hbf9ba987, 32'h40d1c411} /* (2, 6, 31) {real, imag} */,
  {32'hc059d930, 32'h4102fe34} /* (2, 6, 30) {real, imag} */,
  {32'hc08646b6, 32'h415375fa} /* (2, 6, 29) {real, imag} */,
  {32'hc01601f9, 32'h413f12f1} /* (2, 6, 28) {real, imag} */,
  {32'hc0754b05, 32'h414c6112} /* (2, 6, 27) {real, imag} */,
  {32'hc0c96764, 32'h417943c6} /* (2, 6, 26) {real, imag} */,
  {32'hc0b31774, 32'h4186c383} /* (2, 6, 25) {real, imag} */,
  {32'hc0979de8, 32'h4159e994} /* (2, 6, 24) {real, imag} */,
  {32'hc019fd9c, 32'h4122edd1} /* (2, 6, 23) {real, imag} */,
  {32'hc053e515, 32'h413c0afa} /* (2, 6, 22) {real, imag} */,
  {32'hc076f21d, 32'h412d8eae} /* (2, 6, 21) {real, imag} */,
  {32'h401467aa, 32'hc0a362ec} /* (2, 6, 20) {real, imag} */,
  {32'h405d4dec, 32'hc1262b18} /* (2, 6, 19) {real, imag} */,
  {32'h400d403b, 32'hc1564b0a} /* (2, 6, 18) {real, imag} */,
  {32'h4011959d, 32'hc1545a84} /* (2, 6, 17) {real, imag} */,
  {32'h408f3d67, 32'hc163087a} /* (2, 6, 16) {real, imag} */,
  {32'h40a0c56e, 32'hc16789fa} /* (2, 6, 15) {real, imag} */,
  {32'h406db0ee, 32'hc18b3ade} /* (2, 6, 14) {real, imag} */,
  {32'h406fe94a, 32'hc1761d52} /* (2, 6, 13) {real, imag} */,
  {32'h4085f678, 32'hc169169a} /* (2, 6, 12) {real, imag} */,
  {32'h4070c070, 32'hc1314468} /* (2, 6, 11) {real, imag} */,
  {32'hbf3a5ea9, 32'h402395b9} /* (2, 6, 10) {real, imag} */,
  {32'hc087e63c, 32'h4126223f} /* (2, 6, 9) {real, imag} */,
  {32'hc0769526, 32'h413c3408} /* (2, 6, 8) {real, imag} */,
  {32'hbfaafb90, 32'h413d6f79} /* (2, 6, 7) {real, imag} */,
  {32'hc003a184, 32'h41540f97} /* (2, 6, 6) {real, imag} */,
  {32'hc0a04c7c, 32'h4142345d} /* (2, 6, 5) {real, imag} */,
  {32'hc085cdbc, 32'h416d8a42} /* (2, 6, 4) {real, imag} */,
  {32'hc04c9e71, 32'h4170da3e} /* (2, 6, 3) {real, imag} */,
  {32'hc0a0c842, 32'h4160d6b2} /* (2, 6, 2) {real, imag} */,
  {32'hc038d7be, 32'h41520940} /* (2, 6, 1) {real, imag} */,
  {32'hbf46790c, 32'h40e0a89c} /* (2, 6, 0) {real, imag} */,
  {32'hbfd88a78, 32'h40bcf6be} /* (2, 5, 31) {real, imag} */,
  {32'hbf53b20a, 32'h4140703d} /* (2, 5, 30) {real, imag} */,
  {32'hc0163ee6, 32'h418b33c4} /* (2, 5, 29) {real, imag} */,
  {32'hbfe799a3, 32'h41705050} /* (2, 5, 28) {real, imag} */,
  {32'hc093f1f5, 32'h4183193e} /* (2, 5, 27) {real, imag} */,
  {32'hc09cd44e, 32'h4184dc7a} /* (2, 5, 26) {real, imag} */,
  {32'hc07d52d4, 32'h417b9a4d} /* (2, 5, 25) {real, imag} */,
  {32'hbfdcd53b, 32'h41720bb1} /* (2, 5, 24) {real, imag} */,
  {32'hc09f6272, 32'h414f0a34} /* (2, 5, 23) {real, imag} */,
  {32'hc0ace72a, 32'h4149de0d} /* (2, 5, 22) {real, imag} */,
  {32'hc005b348, 32'h4164b32a} /* (2, 5, 21) {real, imag} */,
  {32'hbf17e261, 32'h411fea44} /* (2, 5, 20) {real, imag} */,
  {32'hbfa40210, 32'h40900374} /* (2, 5, 19) {real, imag} */,
  {32'hbfb2748f, 32'h3ffac7e8} /* (2, 5, 18) {real, imag} */,
  {32'hc035e0fa, 32'h40960959} /* (2, 5, 17) {real, imag} */,
  {32'hbd16cfe8, 32'hbefe768e} /* (2, 5, 16) {real, imag} */,
  {32'h3fb6c016, 32'hc10e0306} /* (2, 5, 15) {real, imag} */,
  {32'h4007e0be, 32'hc160fc60} /* (2, 5, 14) {real, imag} */,
  {32'h402e1f86, 32'hc1540993} /* (2, 5, 13) {real, imag} */,
  {32'h40898652, 32'hc163fab1} /* (2, 5, 12) {real, imag} */,
  {32'h40632818, 32'hc181d21b} /* (2, 5, 11) {real, imag} */,
  {32'hbfc269fa, 32'hc11cf982} /* (2, 5, 10) {real, imag} */,
  {32'hbf78d2c7, 32'hc032aab0} /* (2, 5, 9) {real, imag} */,
  {32'hbf4af91a, 32'hc063137f} /* (2, 5, 8) {real, imag} */,
  {32'hbfbc1048, 32'hc0b9a1a7} /* (2, 5, 7) {real, imag} */,
  {32'hbd33c4d8, 32'hc01bebfc} /* (2, 5, 6) {real, imag} */,
  {32'hbfc64b67, 32'h40cc2f81} /* (2, 5, 5) {real, imag} */,
  {32'hbffc1679, 32'h414570bb} /* (2, 5, 4) {real, imag} */,
  {32'hbfbd31f8, 32'h4176c134} /* (2, 5, 3) {real, imag} */,
  {32'hc0a5d6b2, 32'h415f64be} /* (2, 5, 2) {real, imag} */,
  {32'hc0b5f0d3, 32'h414dd6bc} /* (2, 5, 1) {real, imag} */,
  {32'hc019788d, 32'h40ee8942} /* (2, 5, 0) {real, imag} */,
  {32'hc0227103, 32'h40dfaf08} /* (2, 4, 31) {real, imag} */,
  {32'hc064d6c6, 32'h4166acfa} /* (2, 4, 30) {real, imag} */,
  {32'hc05bce11, 32'h41906d3e} /* (2, 4, 29) {real, imag} */,
  {32'hbfe561a5, 32'h4181f9ca} /* (2, 4, 28) {real, imag} */,
  {32'hc0482d6e, 32'h417e9be9} /* (2, 4, 27) {real, imag} */,
  {32'hc00be1bb, 32'h4156b2d8} /* (2, 4, 26) {real, imag} */,
  {32'hbf08e2c8, 32'h41439a2e} /* (2, 4, 25) {real, imag} */,
  {32'h3f4b6805, 32'h417985a6} /* (2, 4, 24) {real, imag} */,
  {32'hc040d33a, 32'h417699d4} /* (2, 4, 23) {real, imag} */,
  {32'hc081ee9b, 32'h416fe47b} /* (2, 4, 22) {real, imag} */,
  {32'hc04d5bbd, 32'h419479b8} /* (2, 4, 21) {real, imag} */,
  {32'hc0670d08, 32'h41906ed2} /* (2, 4, 20) {real, imag} */,
  {32'hc03eea3d, 32'h415e9d1a} /* (2, 4, 19) {real, imag} */,
  {32'hc023bc0e, 32'h41569dac} /* (2, 4, 18) {real, imag} */,
  {32'hc0997415, 32'h417152c4} /* (2, 4, 17) {real, imag} */,
  {32'hc00db662, 32'h4120451d} /* (2, 4, 16) {real, imag} */,
  {32'h40110925, 32'hc0b4c20a} /* (2, 4, 15) {real, imag} */,
  {32'h4045345a, 32'hc136a7db} /* (2, 4, 14) {real, imag} */,
  {32'h3fadc388, 32'hc13d57cc} /* (2, 4, 13) {real, imag} */,
  {32'h409568c3, 32'hc127c508} /* (2, 4, 12) {real, imag} */,
  {32'h40804d1c, 32'hc165b6ab} /* (2, 4, 11) {real, imag} */,
  {32'hbe716550, 32'hc180b914} /* (2, 4, 10) {real, imag} */,
  {32'h3fbf8557, 32'hc1683f2a} /* (2, 4, 9) {real, imag} */,
  {32'h40334b90, 32'hc1777614} /* (2, 4, 8) {real, imag} */,
  {32'h3fba6b75, 32'hc165fac8} /* (2, 4, 7) {real, imag} */,
  {32'h401f3834, 32'hc13b1850} /* (2, 4, 6) {real, imag} */,
  {32'hbeafa313, 32'h40bad6a4} /* (2, 4, 5) {real, imag} */,
  {32'hc0320b2e, 32'h415bb8f6} /* (2, 4, 4) {real, imag} */,
  {32'hc0342d5a, 32'h417e626e} /* (2, 4, 3) {real, imag} */,
  {32'hc0515c0b, 32'h41752ff9} /* (2, 4, 2) {real, imag} */,
  {32'hc0bbb685, 32'h412cf854} /* (2, 4, 1) {real, imag} */,
  {32'hc0353f81, 32'h40ba6936} /* (2, 4, 0) {real, imag} */,
  {32'h3ded73f0, 32'h40f6dcef} /* (2, 3, 31) {real, imag} */,
  {32'hc094dde2, 32'h4186d9c6} /* (2, 3, 30) {real, imag} */,
  {32'hc06bdae6, 32'h418f2a68} /* (2, 3, 29) {real, imag} */,
  {32'h3e953541, 32'h417ce517} /* (2, 3, 28) {real, imag} */,
  {32'h3ed1eb4c, 32'h41623a4d} /* (2, 3, 27) {real, imag} */,
  {32'hbfb3b025, 32'h4138bccd} /* (2, 3, 26) {real, imag} */,
  {32'hc0815b91, 32'h413629b8} /* (2, 3, 25) {real, imag} */,
  {32'hc089f202, 32'h417286f4} /* (2, 3, 24) {real, imag} */,
  {32'hc04023fc, 32'h417c9c14} /* (2, 3, 23) {real, imag} */,
  {32'hc02a4cc0, 32'h418176e1} /* (2, 3, 22) {real, imag} */,
  {32'hc04ce9a6, 32'h41752e62} /* (2, 3, 21) {real, imag} */,
  {32'hc02de4ae, 32'h41736ac6} /* (2, 3, 20) {real, imag} */,
  {32'hc0c4e470, 32'h416967be} /* (2, 3, 19) {real, imag} */,
  {32'hc0d1a4f9, 32'h417aca91} /* (2, 3, 18) {real, imag} */,
  {32'hc0696006, 32'h41803bf0} /* (2, 3, 17) {real, imag} */,
  {32'hbf030670, 32'h4125b570} /* (2, 3, 16) {real, imag} */,
  {32'h3fbcdd00, 32'hc10038dc} /* (2, 3, 15) {real, imag} */,
  {32'h3f94120a, 32'hc14c3c06} /* (2, 3, 14) {real, imag} */,
  {32'h3fbad72b, 32'hc15f1470} /* (2, 3, 13) {real, imag} */,
  {32'h404623d2, 32'hc154a672} /* (2, 3, 12) {real, imag} */,
  {32'h4062228e, 32'hc168e039} /* (2, 3, 11) {real, imag} */,
  {32'h3ffbe354, 32'hc1749ff0} /* (2, 3, 10) {real, imag} */,
  {32'h4070880c, 32'hc16193f7} /* (2, 3, 9) {real, imag} */,
  {32'h40a311bd, 32'hc15c5243} /* (2, 3, 8) {real, imag} */,
  {32'h4040ae40, 32'hc1578a6c} /* (2, 3, 7) {real, imag} */,
  {32'h40602a44, 32'hc15558db} /* (2, 3, 6) {real, imag} */,
  {32'hbf45ddb6, 32'h4089abd0} /* (2, 3, 5) {real, imag} */,
  {32'h3d904a30, 32'h415ef3c0} /* (2, 3, 4) {real, imag} */,
  {32'hbf9e2abc, 32'h417e4387} /* (2, 3, 3) {real, imag} */,
  {32'hbfb17a7b, 32'h41907018} /* (2, 3, 2) {real, imag} */,
  {32'hc055d48e, 32'h415b2b54} /* (2, 3, 1) {real, imag} */,
  {32'hbf289ee2, 32'h40b3dd52} /* (2, 3, 0) {real, imag} */,
  {32'hbf82607a, 32'h40ff89c0} /* (2, 2, 31) {real, imag} */,
  {32'hc01ab8a3, 32'h41852ef1} /* (2, 2, 30) {real, imag} */,
  {32'hbfeadd8a, 32'h4180b616} /* (2, 2, 29) {real, imag} */,
  {32'hbf52ed5c, 32'h4172671e} /* (2, 2, 28) {real, imag} */,
  {32'hbf80c270, 32'h415eb8cb} /* (2, 2, 27) {real, imag} */,
  {32'hc00e4d78, 32'h4153d746} /* (2, 2, 26) {real, imag} */,
  {32'hc0cd6eaa, 32'h41632b34} /* (2, 2, 25) {real, imag} */,
  {32'hc098f1cd, 32'h417d3946} /* (2, 2, 24) {real, imag} */,
  {32'hc034ce82, 32'h41800f8a} /* (2, 2, 23) {real, imag} */,
  {32'hc0480fa2, 32'h413c795e} /* (2, 2, 22) {real, imag} */,
  {32'hc01d2590, 32'h413b0f04} /* (2, 2, 21) {real, imag} */,
  {32'hc03c5d51, 32'h417038ad} /* (2, 2, 20) {real, imag} */,
  {32'hc0c8385f, 32'h41841b06} /* (2, 2, 19) {real, imag} */,
  {32'hc11c4fba, 32'h416b6cda} /* (2, 2, 18) {real, imag} */,
  {32'hc0fb8c0c, 32'h416b0750} /* (2, 2, 17) {real, imag} */,
  {32'hbfd8833b, 32'h4108a8f8} /* (2, 2, 16) {real, imag} */,
  {32'h3f9837ea, 32'hc1148f80} /* (2, 2, 15) {real, imag} */,
  {32'h3ff75afc, 32'hc14fc892} /* (2, 2, 14) {real, imag} */,
  {32'h407a43d0, 32'hc1653e5f} /* (2, 2, 13) {real, imag} */,
  {32'h3fe8f713, 32'hc166c89e} /* (2, 2, 12) {real, imag} */,
  {32'h4083e4b7, 32'hc1522277} /* (2, 2, 11) {real, imag} */,
  {32'h4099567e, 32'hc15fc42a} /* (2, 2, 10) {real, imag} */,
  {32'h40890d95, 32'hc17c8b68} /* (2, 2, 9) {real, imag} */,
  {32'h40b5170a, 32'hc1599fac} /* (2, 2, 8) {real, imag} */,
  {32'h4030c3a6, 32'hc151b358} /* (2, 2, 7) {real, imag} */,
  {32'h3fc74f40, 32'hc171c01e} /* (2, 2, 6) {real, imag} */,
  {32'hc02d9c68, 32'h3f99459a} /* (2, 2, 5) {real, imag} */,
  {32'hc040acc4, 32'h4167ed73} /* (2, 2, 4) {real, imag} */,
  {32'hc017a68e, 32'h417e892b} /* (2, 2, 3) {real, imag} */,
  {32'hc05b05a2, 32'h4188b10a} /* (2, 2, 2) {real, imag} */,
  {32'hc0b5af07, 32'h4170bdc6} /* (2, 2, 1) {real, imag} */,
  {32'hc044c696, 32'h40c38da2} /* (2, 2, 0) {real, imag} */,
  {32'hc017d2a5, 32'h40c994e8} /* (2, 1, 31) {real, imag} */,
  {32'hc048b23a, 32'h413dedc5} /* (2, 1, 30) {real, imag} */,
  {32'hc065dc5b, 32'h415ee71e} /* (2, 1, 29) {real, imag} */,
  {32'hc02463da, 32'h41554bf5} /* (2, 1, 28) {real, imag} */,
  {32'hbfc6107b, 32'h4171bd89} /* (2, 1, 27) {real, imag} */,
  {32'hbf6c20d5, 32'h415ad129} /* (2, 1, 26) {real, imag} */,
  {32'hc08a87fa, 32'h415adeaa} /* (2, 1, 25) {real, imag} */,
  {32'hc08b522c, 32'h4174b13c} /* (2, 1, 24) {real, imag} */,
  {32'hc008a0f8, 32'h4183c354} /* (2, 1, 23) {real, imag} */,
  {32'hbf684378, 32'h415020e8} /* (2, 1, 22) {real, imag} */,
  {32'hbf126e63, 32'h41395606} /* (2, 1, 21) {real, imag} */,
  {32'hc015de9e, 32'h415fe496} /* (2, 1, 20) {real, imag} */,
  {32'hc0706d43, 32'h41788ffb} /* (2, 1, 19) {real, imag} */,
  {32'hc10eb30e, 32'h418da710} /* (2, 1, 18) {real, imag} */,
  {32'hc0a42dfa, 32'h418a329f} /* (2, 1, 17) {real, imag} */,
  {32'hbfd5a4a8, 32'h40f3d5f1} /* (2, 1, 16) {real, imag} */,
  {32'h3f4c58e8, 32'hc1179a4c} /* (2, 1, 15) {real, imag} */,
  {32'h4017cc2b, 32'hc16b9cf8} /* (2, 1, 14) {real, imag} */,
  {32'h40c1755a, 32'hc17c8a3b} /* (2, 1, 13) {real, imag} */,
  {32'h40a256b4, 32'hc176052e} /* (2, 1, 12) {real, imag} */,
  {32'h4053fe52, 32'hc14fdfed} /* (2, 1, 11) {real, imag} */,
  {32'h40210d5a, 32'hc1794304} /* (2, 1, 10) {real, imag} */,
  {32'h40268b5c, 32'hc1847a92} /* (2, 1, 9) {real, imag} */,
  {32'h400fd340, 32'hc165bf40} /* (2, 1, 8) {real, imag} */,
  {32'h4041cb22, 32'hc17422a4} /* (2, 1, 7) {real, imag} */,
  {32'h401b28e8, 32'hc1884e3e} /* (2, 1, 6) {real, imag} */,
  {32'hbf886cee, 32'h3f921506} /* (2, 1, 5) {real, imag} */,
  {32'hc0b5b47e, 32'h41673e26} /* (2, 1, 4) {real, imag} */,
  {32'hc0889218, 32'h416fcc1f} /* (2, 1, 3) {real, imag} */,
  {32'hc01646e6, 32'h415c1128} /* (2, 1, 2) {real, imag} */,
  {32'hc0a594f1, 32'h414b82df} /* (2, 1, 1) {real, imag} */,
  {32'hc08665e8, 32'h40d59646} /* (2, 1, 0) {real, imag} */,
  {32'hc01ea9c2, 32'h405573a2} /* (2, 0, 31) {real, imag} */,
  {32'hc01017e8, 32'h40b2bdf4} /* (2, 0, 30) {real, imag} */,
  {32'hbfec5a25, 32'h40ed2504} /* (2, 0, 29) {real, imag} */,
  {32'hbf9c33eb, 32'h40f6f3e9} /* (2, 0, 28) {real, imag} */,
  {32'hbf8ce83c, 32'h4106f129} /* (2, 0, 27) {real, imag} */,
  {32'h3ef73516, 32'h410d1a9e} /* (2, 0, 26) {real, imag} */,
  {32'hbfd28671, 32'h40d6e410} /* (2, 0, 25) {real, imag} */,
  {32'hc03fc071, 32'h40e20e80} /* (2, 0, 24) {real, imag} */,
  {32'hbfdaa77d, 32'h411d2d1c} /* (2, 0, 23) {real, imag} */,
  {32'hbff02ee3, 32'h41013334} /* (2, 0, 22) {real, imag} */,
  {32'hbffb61cc, 32'h40c2936a} /* (2, 0, 21) {real, imag} */,
  {32'hbfb90842, 32'h40f8398e} /* (2, 0, 20) {real, imag} */,
  {32'hc00b4cc0, 32'h410067e1} /* (2, 0, 19) {real, imag} */,
  {32'hc08b0743, 32'h411d988a} /* (2, 0, 18) {real, imag} */,
  {32'hbf971482, 32'h4117f687} /* (2, 0, 17) {real, imag} */,
  {32'hbec1e074, 32'h400c2d24} /* (2, 0, 16) {real, imag} */,
  {32'hbd891488, 32'hc0c63af6} /* (2, 0, 15) {real, imag} */,
  {32'h3ee15476, 32'hc10fc311} /* (2, 0, 14) {real, imag} */,
  {32'h40024147, 32'hc1298237} /* (2, 0, 13) {real, imag} */,
  {32'h4061874e, 32'hc111df22} /* (2, 0, 12) {real, imag} */,
  {32'h4051bad4, 32'hc10111a5} /* (2, 0, 11) {real, imag} */,
  {32'h3fc0e5b0, 32'hc0f09574} /* (2, 0, 10) {real, imag} */,
  {32'h4008a9a3, 32'hc0bd340a} /* (2, 0, 9) {real, imag} */,
  {32'h3f304bbe, 32'hc0cda0eb} /* (2, 0, 8) {real, imag} */,
  {32'h403a82fe, 32'hc10c8e4e} /* (2, 0, 7) {real, imag} */,
  {32'h4046b414, 32'hc10e26f4} /* (2, 0, 6) {real, imag} */,
  {32'h3f0bd734, 32'h3fdb67e6} /* (2, 0, 5) {real, imag} */,
  {32'hbfd6a6b1, 32'h40ebe3c6} /* (2, 0, 4) {real, imag} */,
  {32'hc022fbb1, 32'h40fb4586} /* (2, 0, 3) {real, imag} */,
  {32'hbf5c161f, 32'h40d9dc42} /* (2, 0, 2) {real, imag} */,
  {32'hbfdb09f6, 32'h40ec5f82} /* (2, 0, 1) {real, imag} */,
  {32'hc01e342c, 32'h40bde6ae} /* (2, 0, 0) {real, imag} */,
  {32'h3f3e33ba, 32'hc0406ff4} /* (1, 31, 31) {real, imag} */,
  {32'h3df0f9d4, 32'hc0f3cc9e} /* (1, 31, 30) {real, imag} */,
  {32'hbe930cb6, 32'hc0c28aa6} /* (1, 31, 29) {real, imag} */,
  {32'hbf3aa0a1, 32'hc08a903e} /* (1, 31, 28) {real, imag} */,
  {32'h3da09cb4, 32'hc089860d} /* (1, 31, 27) {real, imag} */,
  {32'hbe03f53e, 32'hc0a25dba} /* (1, 31, 26) {real, imag} */,
  {32'h4018811e, 32'hc08b8e38} /* (1, 31, 25) {real, imag} */,
  {32'hbed25468, 32'hc0a37598} /* (1, 31, 24) {real, imag} */,
  {32'hbf8f21b5, 32'hc0a48d23} /* (1, 31, 23) {real, imag} */,
  {32'hbf5c8ddd, 32'hc0d2a772} /* (1, 31, 22) {real, imag} */,
  {32'h3f60a13c, 32'hc02eff23} /* (1, 31, 21) {real, imag} */,
  {32'h3fa1f960, 32'h405c68f2} /* (1, 31, 20) {real, imag} */,
  {32'h3fb7bf2e, 32'h40675295} /* (1, 31, 19) {real, imag} */,
  {32'hbe7cb3c4, 32'h40824455} /* (1, 31, 18) {real, imag} */,
  {32'h3e8919da, 32'h40474011} /* (1, 31, 17) {real, imag} */,
  {32'hbe508a40, 32'h40b2d2b2} /* (1, 31, 16) {real, imag} */,
  {32'h3f7df615, 32'h40beb4d2} /* (1, 31, 15) {real, imag} */,
  {32'h3f6a5189, 32'h408d614f} /* (1, 31, 14) {real, imag} */,
  {32'h3fb4254a, 32'h4086056e} /* (1, 31, 13) {real, imag} */,
  {32'hbef07825, 32'h40922bbe} /* (1, 31, 12) {real, imag} */,
  {32'h3ebb1666, 32'h403ae851} /* (1, 31, 11) {real, imag} */,
  {32'h3d6c1b4c, 32'hc08647cc} /* (1, 31, 10) {real, imag} */,
  {32'h3f3f4f88, 32'hc036def2} /* (1, 31, 9) {real, imag} */,
  {32'h401dae88, 32'hc06702fd} /* (1, 31, 8) {real, imag} */,
  {32'h3f65fc5a, 32'hc0826525} /* (1, 31, 7) {real, imag} */,
  {32'hbfdf4916, 32'hc08f9dfd} /* (1, 31, 6) {real, imag} */,
  {32'hbd618a90, 32'hc093e12f} /* (1, 31, 5) {real, imag} */,
  {32'h3edf7962, 32'hc05b6c55} /* (1, 31, 4) {real, imag} */,
  {32'h3f2036d2, 32'hc02acd4c} /* (1, 31, 3) {real, imag} */,
  {32'h3d01148c, 32'hbfd78983} /* (1, 31, 2) {real, imag} */,
  {32'h3f45a380, 32'hc07e3bdc} /* (1, 31, 1) {real, imag} */,
  {32'h3f338ca5, 32'hc020666a} /* (1, 31, 0) {real, imag} */,
  {32'h3f8d8e6a, 32'hc091158a} /* (1, 30, 31) {real, imag} */,
  {32'h403c8724, 32'hc1299a68} /* (1, 30, 30) {real, imag} */,
  {32'h4099d85c, 32'hc11dd9f7} /* (1, 30, 29) {real, imag} */,
  {32'h40064a5e, 32'hc0de3687} /* (1, 30, 28) {real, imag} */,
  {32'h4030b5c6, 32'hc09c984a} /* (1, 30, 27) {real, imag} */,
  {32'h3f3ff99e, 32'hc0a421e6} /* (1, 30, 26) {real, imag} */,
  {32'h3f6694fc, 32'hc0d209dd} /* (1, 30, 25) {real, imag} */,
  {32'h3e6152cd, 32'hc11fb032} /* (1, 30, 24) {real, imag} */,
  {32'h3f8c2a69, 32'hc0f24654} /* (1, 30, 23) {real, imag} */,
  {32'h3e9aa86e, 32'hc11f393e} /* (1, 30, 22) {real, imag} */,
  {32'h401fbec6, 32'hc05a5ef2} /* (1, 30, 21) {real, imag} */,
  {32'hbebe9b8e, 32'h41171088} /* (1, 30, 20) {real, imag} */,
  {32'hbf9033c6, 32'h410006e9} /* (1, 30, 19) {real, imag} */,
  {32'hbfa51a8a, 32'h411a2e18} /* (1, 30, 18) {real, imag} */,
  {32'hbf08c376, 32'h40d4fb80} /* (1, 30, 17) {real, imag} */,
  {32'hbf5e4760, 32'h41199259} /* (1, 30, 16) {real, imag} */,
  {32'hbfacd556, 32'h4114fa20} /* (1, 30, 15) {real, imag} */,
  {32'hc090f5c8, 32'h410ed162} /* (1, 30, 14) {real, imag} */,
  {32'hc07135ae, 32'h41049922} /* (1, 30, 13) {real, imag} */,
  {32'hbfb0b31e, 32'h40df1bd8} /* (1, 30, 12) {real, imag} */,
  {32'hbfaa849c, 32'h408745be} /* (1, 30, 11) {real, imag} */,
  {32'hc0627ba0, 32'hc096b352} /* (1, 30, 10) {real, imag} */,
  {32'h3e1d8cf2, 32'hc09ffdca} /* (1, 30, 9) {real, imag} */,
  {32'h404a156a, 32'hc1082ec6} /* (1, 30, 8) {real, imag} */,
  {32'h3fc58f4b, 32'hc0e1fb70} /* (1, 30, 7) {real, imag} */,
  {32'hc016c686, 32'hc0b3456b} /* (1, 30, 6) {real, imag} */,
  {32'hbfbe3c6e, 32'hc0f8dbff} /* (1, 30, 5) {real, imag} */,
  {32'h3fb080d4, 32'hc0cf08b4} /* (1, 30, 4) {real, imag} */,
  {32'h4029ab14, 32'hc0b9f85c} /* (1, 30, 3) {real, imag} */,
  {32'h3fca2fa0, 32'hc0d2f373} /* (1, 30, 2) {real, imag} */,
  {32'h3ff7440c, 32'hc10a2035} /* (1, 30, 1) {real, imag} */,
  {32'h3f80fb6e, 32'hc080f559} /* (1, 30, 0) {real, imag} */,
  {32'h3fe26e4e, 32'hc0a1a97a} /* (1, 29, 31) {real, imag} */,
  {32'h400e7512, 32'hc11d636e} /* (1, 29, 30) {real, imag} */,
  {32'h3ff23e4d, 32'hc0c08b68} /* (1, 29, 29) {real, imag} */,
  {32'h3fe52446, 32'hc0a0dd0a} /* (1, 29, 28) {real, imag} */,
  {32'h3ee5d564, 32'hc09fceba} /* (1, 29, 27) {real, imag} */,
  {32'hbfd9e8f8, 32'hc0c34258} /* (1, 29, 26) {real, imag} */,
  {32'h3ea06c74, 32'hc0d5e27c} /* (1, 29, 25) {real, imag} */,
  {32'h402e894c, 32'hc0cf07ba} /* (1, 29, 24) {real, imag} */,
  {32'h3fa7ba30, 32'hc0c518de} /* (1, 29, 23) {real, imag} */,
  {32'hbf80e7e5, 32'hc106ca24} /* (1, 29, 22) {real, imag} */,
  {32'hbff032b0, 32'hc0a9426b} /* (1, 29, 21) {real, imag} */,
  {32'hc0ac7af6, 32'h4102ace9} /* (1, 29, 20) {real, imag} */,
  {32'hbfb1637b, 32'h40f568ee} /* (1, 29, 19) {real, imag} */,
  {32'hc028bbca, 32'h41189014} /* (1, 29, 18) {real, imag} */,
  {32'hc05b5cc9, 32'h40c049cc} /* (1, 29, 17) {real, imag} */,
  {32'hbfb1a6ad, 32'h40b0a810} /* (1, 29, 16) {real, imag} */,
  {32'hbfe8500a, 32'h40fbf634} /* (1, 29, 15) {real, imag} */,
  {32'hc08de528, 32'h40e26604} /* (1, 29, 14) {real, imag} */,
  {32'hc0b22285, 32'h40e85e0f} /* (1, 29, 13) {real, imag} */,
  {32'hc00f2632, 32'h40cc3302} /* (1, 29, 12) {real, imag} */,
  {32'hc02bc2b6, 32'h40933b41} /* (1, 29, 11) {real, imag} */,
  {32'hc0a78254, 32'hbf9b741e} /* (1, 29, 10) {real, imag} */,
  {32'hbee0b086, 32'hc08b8a6c} /* (1, 29, 9) {real, imag} */,
  {32'h408b2f2e, 32'hc1218358} /* (1, 29, 8) {real, imag} */,
  {32'h3fc69bb2, 32'hc112e0c7} /* (1, 29, 7) {real, imag} */,
  {32'hbeda995b, 32'hc0a87132} /* (1, 29, 6) {real, imag} */,
  {32'hc0023d00, 32'hc0963c0a} /* (1, 29, 5) {real, imag} */,
  {32'hbef64539, 32'hc06159ae} /* (1, 29, 4) {real, imag} */,
  {32'h401b25c3, 32'hc0c4c8d8} /* (1, 29, 3) {real, imag} */,
  {32'h3ff46b51, 32'hc10f2413} /* (1, 29, 2) {real, imag} */,
  {32'h3ed9a390, 32'hc13f422c} /* (1, 29, 1) {real, imag} */,
  {32'h3fad3bb1, 32'hc092e6aa} /* (1, 29, 0) {real, imag} */,
  {32'h3fe6fd5a, 32'hc0ae522a} /* (1, 28, 31) {real, imag} */,
  {32'h3f804398, 32'hc1061616} /* (1, 28, 30) {real, imag} */,
  {32'hbe106590, 32'hc0cbd3fd} /* (1, 28, 29) {real, imag} */,
  {32'h3fa4163f, 32'hc0c2e2f5} /* (1, 28, 28) {real, imag} */,
  {32'hbf46b255, 32'hc0b7b5f2} /* (1, 28, 27) {real, imag} */,
  {32'hbf8078fe, 32'hc0ce4218} /* (1, 28, 26) {real, imag} */,
  {32'h4066aeeb, 32'hc1116fcc} /* (1, 28, 25) {real, imag} */,
  {32'h40baf834, 32'hc1253f2e} /* (1, 28, 24) {real, imag} */,
  {32'h3f60cd8a, 32'hc12bd523} /* (1, 28, 23) {real, imag} */,
  {32'hc005db3d, 32'hc12279cf} /* (1, 28, 22) {real, imag} */,
  {32'hbee260b2, 32'hc0c8926e} /* (1, 28, 21) {real, imag} */,
  {32'hbfbad340, 32'h407c24c3} /* (1, 28, 20) {real, imag} */,
  {32'hbe2b2f11, 32'h40c90ddf} /* (1, 28, 19) {real, imag} */,
  {32'hc0094472, 32'h4132ae34} /* (1, 28, 18) {real, imag} */,
  {32'hbf4d0dbf, 32'h410f0788} /* (1, 28, 17) {real, imag} */,
  {32'hbd1df618, 32'h4107abea} /* (1, 28, 16) {real, imag} */,
  {32'hc068b29c, 32'h4124d76f} /* (1, 28, 15) {real, imag} */,
  {32'hc09c91ab, 32'h41059ce8} /* (1, 28, 14) {real, imag} */,
  {32'hc080ba32, 32'h40ac4f79} /* (1, 28, 13) {real, imag} */,
  {32'hbfb9fa06, 32'h40ee52e0} /* (1, 28, 12) {real, imag} */,
  {32'hc00c5b4e, 32'h40f07383} /* (1, 28, 11) {real, imag} */,
  {32'hbec9143e, 32'hbfd2f5b0} /* (1, 28, 10) {real, imag} */,
  {32'h3fd79bee, 32'hc0c53143} /* (1, 28, 9) {real, imag} */,
  {32'h3fbe7681, 32'hc0ec81b8} /* (1, 28, 8) {real, imag} */,
  {32'h3faf62e8, 32'hc0ea3220} /* (1, 28, 7) {real, imag} */,
  {32'h4010d493, 32'hc0e1f2b9} /* (1, 28, 6) {real, imag} */,
  {32'hbec3bb45, 32'hc108eeec} /* (1, 28, 5) {real, imag} */,
  {32'h3dc39caa, 32'hc11e3d1e} /* (1, 28, 4) {real, imag} */,
  {32'h401456f4, 32'hc112ed8e} /* (1, 28, 3) {real, imag} */,
  {32'h404d5afa, 32'hc1003eab} /* (1, 28, 2) {real, imag} */,
  {32'h4001fa5b, 32'hc114890f} /* (1, 28, 1) {real, imag} */,
  {32'h3f936de9, 32'hc0895519} /* (1, 28, 0) {real, imag} */,
  {32'h40286a18, 32'hc0aa60b7} /* (1, 27, 31) {real, imag} */,
  {32'hbf2805a4, 32'hc10b2b08} /* (1, 27, 30) {real, imag} */,
  {32'hc01f7092, 32'hc1191bfe} /* (1, 27, 29) {real, imag} */,
  {32'hbf04da33, 32'hc0e968cb} /* (1, 27, 28) {real, imag} */,
  {32'h3f2bc5ca, 32'hc0f568d0} /* (1, 27, 27) {real, imag} */,
  {32'h3faa2744, 32'hc128ef7c} /* (1, 27, 26) {real, imag} */,
  {32'h3ed9972b, 32'hc12c8f1b} /* (1, 27, 25) {real, imag} */,
  {32'h400d96b7, 32'hc133cd78} /* (1, 27, 24) {real, imag} */,
  {32'hbead19a1, 32'hc1367e68} /* (1, 27, 23) {real, imag} */,
  {32'hbfff158a, 32'hc100a812} /* (1, 27, 22) {real, imag} */,
  {32'h3f8ca4ae, 32'hc04b712c} /* (1, 27, 21) {real, imag} */,
  {32'h4003c7bc, 32'h407a8483} /* (1, 27, 20) {real, imag} */,
  {32'h401b7c2c, 32'h40e34cdd} /* (1, 27, 19) {real, imag} */,
  {32'hbea8b4a0, 32'h4115ee26} /* (1, 27, 18) {real, imag} */,
  {32'hbedd594c, 32'h4118890b} /* (1, 27, 17) {real, imag} */,
  {32'hbed91f6a, 32'h412b0334} /* (1, 27, 16) {real, imag} */,
  {32'hbf826200, 32'h4114ed43} /* (1, 27, 15) {real, imag} */,
  {32'hc05ed63c, 32'h4106ade9} /* (1, 27, 14) {real, imag} */,
  {32'hc04a02ce, 32'h40d1fbfa} /* (1, 27, 13) {real, imag} */,
  {32'h3f3310b0, 32'h40e5ad19} /* (1, 27, 12) {real, imag} */,
  {32'h40157cdd, 32'h410a392f} /* (1, 27, 11) {real, imag} */,
  {32'h402ccc1c, 32'hbf83751d} /* (1, 27, 10) {real, imag} */,
  {32'h409102a7, 32'hc119d613} /* (1, 27, 9) {real, imag} */,
  {32'h40745090, 32'hc10d646b} /* (1, 27, 8) {real, imag} */,
  {32'h406fb87c, 32'hc1003f7c} /* (1, 27, 7) {real, imag} */,
  {32'h3fe5a972, 32'hc1096692} /* (1, 27, 6) {real, imag} */,
  {32'h401424a0, 32'hc13c9936} /* (1, 27, 5) {real, imag} */,
  {32'h40587ff3, 32'hc16180d3} /* (1, 27, 4) {real, imag} */,
  {32'h40064d51, 32'hc111e618} /* (1, 27, 3) {real, imag} */,
  {32'h3faf2f84, 32'hc0ca4951} /* (1, 27, 2) {real, imag} */,
  {32'h3fee6d36, 32'hc0f5f82e} /* (1, 27, 1) {real, imag} */,
  {32'h3ea1c760, 32'hc0b04fe7} /* (1, 27, 0) {real, imag} */,
  {32'h3fe30119, 32'hc073f22c} /* (1, 26, 31) {real, imag} */,
  {32'hbf8cd09c, 32'hc103f50d} /* (1, 26, 30) {real, imag} */,
  {32'hc059e721, 32'hc1499391} /* (1, 26, 29) {real, imag} */,
  {32'hbfc535eb, 32'hc1320b80} /* (1, 26, 28) {real, imag} */,
  {32'h400cf535, 32'hc11c55db} /* (1, 26, 27) {real, imag} */,
  {32'h4002fbf6, 32'hc140a36b} /* (1, 26, 26) {real, imag} */,
  {32'hbff7c4e7, 32'hc1491e84} /* (1, 26, 25) {real, imag} */,
  {32'h40090f22, 32'hc1072ed2} /* (1, 26, 24) {real, imag} */,
  {32'h3f0c9cac, 32'hc0dc41b8} /* (1, 26, 23) {real, imag} */,
  {32'hbef6efd7, 32'hc0efac28} /* (1, 26, 22) {real, imag} */,
  {32'h3f7b8df8, 32'hc08444e8} /* (1, 26, 21) {real, imag} */,
  {32'h3f410203, 32'h404f2f8c} /* (1, 26, 20) {real, imag} */,
  {32'h3f230e8c, 32'h410aa014} /* (1, 26, 19) {real, imag} */,
  {32'hbea7fdd7, 32'h40eabbbc} /* (1, 26, 18) {real, imag} */,
  {32'h3f2e3908, 32'h40f826b4} /* (1, 26, 17) {real, imag} */,
  {32'h3f87fffa, 32'h411b68e2} /* (1, 26, 16) {real, imag} */,
  {32'hbfd7368d, 32'h40b8fa7d} /* (1, 26, 15) {real, imag} */,
  {32'hc04041df, 32'h40f38238} /* (1, 26, 14) {real, imag} */,
  {32'hc077a4e1, 32'h410f47ec} /* (1, 26, 13) {real, imag} */,
  {32'hbf514abe, 32'h40c3c0d6} /* (1, 26, 12) {real, imag} */,
  {32'h3d205250, 32'h409062ce} /* (1, 26, 11) {real, imag} */,
  {32'h3fbf4df1, 32'hc0bfd2f3} /* (1, 26, 10) {real, imag} */,
  {32'h40070209, 32'hc14d53f1} /* (1, 26, 9) {real, imag} */,
  {32'h406ec56d, 32'hc129f7bd} /* (1, 26, 8) {real, imag} */,
  {32'h40176ae6, 32'hc12826e2} /* (1, 26, 7) {real, imag} */,
  {32'h3f77631c, 32'hc0f5ba39} /* (1, 26, 6) {real, imag} */,
  {32'h400c50c8, 32'hc0d9145d} /* (1, 26, 5) {real, imag} */,
  {32'h400fca36, 32'hc112443a} /* (1, 26, 4) {real, imag} */,
  {32'h3f4a9f86, 32'hc0edd56d} /* (1, 26, 3) {real, imag} */,
  {32'h3ef35f05, 32'hc0e9466f} /* (1, 26, 2) {real, imag} */,
  {32'h401453e3, 32'hc116a864} /* (1, 26, 1) {real, imag} */,
  {32'h3fa4d427, 32'hc0b85ea7} /* (1, 26, 0) {real, imag} */,
  {32'h3fb3afb5, 32'hc0a0f3b0} /* (1, 25, 31) {real, imag} */,
  {32'h3f29415f, 32'hc10eb610} /* (1, 25, 30) {real, imag} */,
  {32'hbfd3151e, 32'hc129e9fa} /* (1, 25, 29) {real, imag} */,
  {32'hc02b4110, 32'hc12f22a7} /* (1, 25, 28) {real, imag} */,
  {32'h400da622, 32'hc10d41f6} /* (1, 25, 27) {real, imag} */,
  {32'h404c428e, 32'hc10c05b6} /* (1, 25, 26) {real, imag} */,
  {32'hc028fca2, 32'hc12779e4} /* (1, 25, 25) {real, imag} */,
  {32'hbfa815c2, 32'hc0f313d6} /* (1, 25, 24) {real, imag} */,
  {32'h3f8ee2fa, 32'hc0a41b1f} /* (1, 25, 23) {real, imag} */,
  {32'h3f475121, 32'hc0ced002} /* (1, 25, 22) {real, imag} */,
  {32'h3ecc40bc, 32'hc0853b64} /* (1, 25, 21) {real, imag} */,
  {32'hbf17f57c, 32'h40a24d44} /* (1, 25, 20) {real, imag} */,
  {32'hbe1c7110, 32'h412130e0} /* (1, 25, 19) {real, imag} */,
  {32'h3fa4aff6, 32'h410dae24} /* (1, 25, 18) {real, imag} */,
  {32'h3fd9d589, 32'h412070b6} /* (1, 25, 17) {real, imag} */,
  {32'h40522e7c, 32'h411d6f3a} /* (1, 25, 16) {real, imag} */,
  {32'hbf7a0346, 32'h40985339} /* (1, 25, 15) {real, imag} */,
  {32'hc07e2e62, 32'h40f26b04} /* (1, 25, 14) {real, imag} */,
  {32'hc037e23e, 32'h413148dc} /* (1, 25, 13) {real, imag} */,
  {32'hc031c6b6, 32'h40ffa739} /* (1, 25, 12) {real, imag} */,
  {32'hbfc71602, 32'h4017da24} /* (1, 25, 11) {real, imag} */,
  {32'h3ff3892e, 32'hc1079c7c} /* (1, 25, 10) {real, imag} */,
  {32'hbf9ea37e, 32'hc14937d3} /* (1, 25, 9) {real, imag} */,
  {32'hbed686b4, 32'hc10d218a} /* (1, 25, 8) {real, imag} */,
  {32'h3f2933b6, 32'hc101504f} /* (1, 25, 7) {real, imag} */,
  {32'h3f2fe4bc, 32'hc0e8161a} /* (1, 25, 6) {real, imag} */,
  {32'h3e7779d4, 32'hc0d70052} /* (1, 25, 5) {real, imag} */,
  {32'hbf3ac76a, 32'hc102c86c} /* (1, 25, 4) {real, imag} */,
  {32'hbec234b6, 32'hc10c669d} /* (1, 25, 3) {real, imag} */,
  {32'h3efca8ef, 32'hc10a7408} /* (1, 25, 2) {real, imag} */,
  {32'hbf2f815f, 32'hc116a046} /* (1, 25, 1) {real, imag} */,
  {32'hbfb6842b, 32'hc08c47e6} /* (1, 25, 0) {real, imag} */,
  {32'h3dd67418, 32'hc0722b44} /* (1, 24, 31) {real, imag} */,
  {32'h3fe028ee, 32'hc0dc5ef8} /* (1, 24, 30) {real, imag} */,
  {32'hbf475944, 32'hc0b2648e} /* (1, 24, 29) {real, imag} */,
  {32'hc00f14e6, 32'hc10aa046} /* (1, 24, 28) {real, imag} */,
  {32'h3fe27fc2, 32'hc0ddbf10} /* (1, 24, 27) {real, imag} */,
  {32'h402c91ed, 32'hc0901bbe} /* (1, 24, 26) {real, imag} */,
  {32'hbd86acf4, 32'hc0e486e2} /* (1, 24, 25) {real, imag} */,
  {32'h3e0e781c, 32'hc0e11f44} /* (1, 24, 24) {real, imag} */,
  {32'h4063baab, 32'hc0c4401d} /* (1, 24, 23) {real, imag} */,
  {32'h40266d6c, 32'hc0f67ec0} /* (1, 24, 22) {real, imag} */,
  {32'h400a372d, 32'hc0836a4e} /* (1, 24, 21) {real, imag} */,
  {32'hbcd3afe0, 32'h40df4f65} /* (1, 24, 20) {real, imag} */,
  {32'hbfdceb0e, 32'h410bc4c6} /* (1, 24, 19) {real, imag} */,
  {32'h3f1244e4, 32'h40dd5787} /* (1, 24, 18) {real, imag} */,
  {32'h3e9e62a3, 32'h410fbd9a} /* (1, 24, 17) {real, imag} */,
  {32'hbde2d010, 32'h410cbcca} /* (1, 24, 16) {real, imag} */,
  {32'hbf668b19, 32'h40f14e5e} /* (1, 24, 15) {real, imag} */,
  {32'hc013e0bd, 32'h40e7a852} /* (1, 24, 14) {real, imag} */,
  {32'h3f11ad4d, 32'h41187580} /* (1, 24, 13) {real, imag} */,
  {32'hbf2fd0c3, 32'h41006caa} /* (1, 24, 12) {real, imag} */,
  {32'h3fad57e9, 32'h40286abd} /* (1, 24, 11) {real, imag} */,
  {32'h3fdd1c04, 32'hc0e86704} /* (1, 24, 10) {real, imag} */,
  {32'hbe55182c, 32'hc12569ee} /* (1, 24, 9) {real, imag} */,
  {32'h40244481, 32'hc105d348} /* (1, 24, 8) {real, imag} */,
  {32'h4028aaf6, 32'hc111a38d} /* (1, 24, 7) {real, imag} */,
  {32'h4048ef0c, 32'hc0fb8250} /* (1, 24, 6) {real, imag} */,
  {32'h3f4b4015, 32'hc0e12a4c} /* (1, 24, 5) {real, imag} */,
  {32'hbf2c3f15, 32'hc1130e00} /* (1, 24, 4) {real, imag} */,
  {32'h3ff37078, 32'hc1306de2} /* (1, 24, 3) {real, imag} */,
  {32'h404693f6, 32'hc10f8a3e} /* (1, 24, 2) {real, imag} */,
  {32'h3e4bb654, 32'hc0d71c0d} /* (1, 24, 1) {real, imag} */,
  {32'hbff3ae2c, 32'hc05576da} /* (1, 24, 0) {real, imag} */,
  {32'hbec471f2, 32'hc03bbac5} /* (1, 23, 31) {real, imag} */,
  {32'hbf147dcc, 32'hc0f6b335} /* (1, 23, 30) {real, imag} */,
  {32'hbfc8a022, 32'hc101e6f4} /* (1, 23, 29) {real, imag} */,
  {32'h3d493200, 32'hc1079497} /* (1, 23, 28) {real, imag} */,
  {32'h3facf260, 32'hc0c46d18} /* (1, 23, 27) {real, imag} */,
  {32'h3ff54f94, 32'hc0b26ead} /* (1, 23, 26) {real, imag} */,
  {32'h3f9df6cf, 32'hc0e431c6} /* (1, 23, 25) {real, imag} */,
  {32'h3fe33bf2, 32'hc0f3fadc} /* (1, 23, 24) {real, imag} */,
  {32'h40b8ab12, 32'hc126443e} /* (1, 23, 23) {real, imag} */,
  {32'h409d96bf, 32'hc10d42c5} /* (1, 23, 22) {real, imag} */,
  {32'h40811e26, 32'hc056f11d} /* (1, 23, 21) {real, imag} */,
  {32'h3fc62e26, 32'h41011642} /* (1, 23, 20) {real, imag} */,
  {32'hbfb8f2cc, 32'h410fedd0} /* (1, 23, 19) {real, imag} */,
  {32'hbf17f75e, 32'h40c6bf84} /* (1, 23, 18) {real, imag} */,
  {32'h3ff67d20, 32'h40ec893e} /* (1, 23, 17) {real, imag} */,
  {32'hbf949112, 32'h40f5b4c8} /* (1, 23, 16) {real, imag} */,
  {32'hbfbdd10a, 32'h40f2f51d} /* (1, 23, 15) {real, imag} */,
  {32'hbf83f461, 32'h40fc531c} /* (1, 23, 14) {real, imag} */,
  {32'h3f9d0328, 32'h41150166} /* (1, 23, 13) {real, imag} */,
  {32'h3f9eb3db, 32'h41111d97} /* (1, 23, 12) {real, imag} */,
  {32'h40886c1c, 32'h408d00ec} /* (1, 23, 11) {real, imag} */,
  {32'h404e5136, 32'hc060b16e} /* (1, 23, 10) {real, imag} */,
  {32'hbd831ce6, 32'hc0cfddd2} /* (1, 23, 9) {real, imag} */,
  {32'h3fc80c4e, 32'hc0c8808e} /* (1, 23, 8) {real, imag} */,
  {32'h3ff255ae, 32'hc10a3dbb} /* (1, 23, 7) {real, imag} */,
  {32'h401a8308, 32'hc11c2082} /* (1, 23, 6) {real, imag} */,
  {32'h3f019c4e, 32'hc133358a} /* (1, 23, 5) {real, imag} */,
  {32'h3f2a80b3, 32'hc130d0ce} /* (1, 23, 4) {real, imag} */,
  {32'h4019bbc0, 32'hc1017669} /* (1, 23, 3) {real, imag} */,
  {32'h406266e3, 32'hc0be9750} /* (1, 23, 2) {real, imag} */,
  {32'h3f1572c3, 32'hc0e390cc} /* (1, 23, 1) {real, imag} */,
  {32'h3d32fd78, 32'hc0736f1b} /* (1, 23, 0) {real, imag} */,
  {32'hbf6c5cb2, 32'hc06b597c} /* (1, 22, 31) {real, imag} */,
  {32'hbfbe93b6, 32'hc0ed9135} /* (1, 22, 30) {real, imag} */,
  {32'hbfee9fd0, 32'hc11700b4} /* (1, 22, 29) {real, imag} */,
  {32'hc009e994, 32'hc11c5ea0} /* (1, 22, 28) {real, imag} */,
  {32'hbfb6b14b, 32'hc0fc6490} /* (1, 22, 27) {real, imag} */,
  {32'hbe10791b, 32'hc0d61af4} /* (1, 22, 26) {real, imag} */,
  {32'hbe05d6c2, 32'hc0d0daa5} /* (1, 22, 25) {real, imag} */,
  {32'hbf18c4d6, 32'hc0eb0308} /* (1, 22, 24) {real, imag} */,
  {32'h403113a2, 32'hc13c0223} /* (1, 22, 23) {real, imag} */,
  {32'h408fe4cb, 32'hc1252c56} /* (1, 22, 22) {real, imag} */,
  {32'h40105a0e, 32'hc05362c4} /* (1, 22, 21) {real, imag} */,
  {32'h3f8d2c52, 32'h40d178aa} /* (1, 22, 20) {real, imag} */,
  {32'hbdc26ad4, 32'h411fec44} /* (1, 22, 19) {real, imag} */,
  {32'h3f124189, 32'h41237056} /* (1, 22, 18) {real, imag} */,
  {32'h3ec0b9a3, 32'h4102fe6e} /* (1, 22, 17) {real, imag} */,
  {32'hbfd32efe, 32'h41052ca9} /* (1, 22, 16) {real, imag} */,
  {32'hc02522f8, 32'h40ead6ac} /* (1, 22, 15) {real, imag} */,
  {32'hbf233b02, 32'h411222c0} /* (1, 22, 14) {real, imag} */,
  {32'h3f4da032, 32'h412f7e86} /* (1, 22, 13) {real, imag} */,
  {32'h3fe47fde, 32'h415383fd} /* (1, 22, 12) {real, imag} */,
  {32'h402b081f, 32'h4113c8f2} /* (1, 22, 11) {real, imag} */,
  {32'h40105e8e, 32'hc0131490} /* (1, 22, 10) {real, imag} */,
  {32'hbea4caa8, 32'hc103da72} /* (1, 22, 9) {real, imag} */,
  {32'hbe940136, 32'hc101c844} /* (1, 22, 8) {real, imag} */,
  {32'h400ce6f2, 32'hc10f25e5} /* (1, 22, 7) {real, imag} */,
  {32'h3fd8e1e6, 32'hc100ca11} /* (1, 22, 6) {real, imag} */,
  {32'hbee49a24, 32'hc10cced8} /* (1, 22, 5) {real, imag} */,
  {32'h4037cbc7, 32'hc0d49660} /* (1, 22, 4) {real, imag} */,
  {32'h406879cc, 32'hc0cfb8a4} /* (1, 22, 3) {real, imag} */,
  {32'h3fe71258, 32'hc0de7304} /* (1, 22, 2) {real, imag} */,
  {32'h403e8ae0, 32'hc0f68604} /* (1, 22, 1) {real, imag} */,
  {32'h3fc39e77, 32'hc078ced0} /* (1, 22, 0) {real, imag} */,
  {32'hbf7c4bd1, 32'hc0189a02} /* (1, 21, 31) {real, imag} */,
  {32'h3fe9cd3b, 32'hc0bb32a6} /* (1, 21, 30) {real, imag} */,
  {32'h4036796c, 32'hc0c98723} /* (1, 21, 29) {real, imag} */,
  {32'hbf0b57ee, 32'hc0de8062} /* (1, 21, 28) {real, imag} */,
  {32'h3def6460, 32'hc0a49d54} /* (1, 21, 27) {real, imag} */,
  {32'h3fd630ca, 32'hc01d3d96} /* (1, 21, 26) {real, imag} */,
  {32'h40048cc1, 32'hc0ac2ac2} /* (1, 21, 25) {real, imag} */,
  {32'hbf597418, 32'hc08885c4} /* (1, 21, 24) {real, imag} */,
  {32'hbe9c2c22, 32'hc08075ec} /* (1, 21, 23) {real, imag} */,
  {32'hbfe15c09, 32'hc0713c00} /* (1, 21, 22) {real, imag} */,
  {32'hbfde3f4e, 32'hc00377e6} /* (1, 21, 21) {real, imag} */,
  {32'h3ee7a064, 32'h40050ec0} /* (1, 21, 20) {real, imag} */,
  {32'h3e76fed1, 32'h408ab9e4} /* (1, 21, 19) {real, imag} */,
  {32'h3fdcf0a8, 32'h40aed4dc} /* (1, 21, 18) {real, imag} */,
  {32'h3d98c6dc, 32'h408644de} /* (1, 21, 17) {real, imag} */,
  {32'hbf95bc5a, 32'h4002f5d7} /* (1, 21, 16) {real, imag} */,
  {32'hc07f9749, 32'h4000c370} /* (1, 21, 15) {real, imag} */,
  {32'hbfcc9002, 32'h40ab3c8f} /* (1, 21, 14) {real, imag} */,
  {32'h3fad6ef6, 32'h40e4b98e} /* (1, 21, 13) {real, imag} */,
  {32'hbe7cbbf9, 32'h40deef85} /* (1, 21, 12) {real, imag} */,
  {32'h3fd8aa5a, 32'h4022c329} /* (1, 21, 11) {real, imag} */,
  {32'h405da10a, 32'hc08e0e8e} /* (1, 21, 10) {real, imag} */,
  {32'hbec3376d, 32'hc0998e0f} /* (1, 21, 9) {real, imag} */,
  {32'hbfe13e80, 32'hc0c1e174} /* (1, 21, 8) {real, imag} */,
  {32'h3f0b2724, 32'hc0aace6a} /* (1, 21, 7) {real, imag} */,
  {32'h3f9b0220, 32'hbf525b27} /* (1, 21, 6) {real, imag} */,
  {32'hbf8abd1f, 32'hc01d9d17} /* (1, 21, 5) {real, imag} */,
  {32'hbed2fa79, 32'hbffa6cd0} /* (1, 21, 4) {real, imag} */,
  {32'hbe6e9655, 32'hbfcce369} /* (1, 21, 3) {real, imag} */,
  {32'h3f904190, 32'hc05ce936} /* (1, 21, 2) {real, imag} */,
  {32'h3fc491aa, 32'hc06ef1c6} /* (1, 21, 1) {real, imag} */,
  {32'hbf3fd7a2, 32'hbf85104c} /* (1, 21, 0) {real, imag} */,
  {32'hbed8ea6c, 32'h4066c033} /* (1, 20, 31) {real, imag} */,
  {32'h3ff4c8bc, 32'h40d20571} /* (1, 20, 30) {real, imag} */,
  {32'h40886c0a, 32'h40bd4076} /* (1, 20, 29) {real, imag} */,
  {32'h407861e4, 32'h403e0628} /* (1, 20, 28) {real, imag} */,
  {32'h3fa76193, 32'h40a6a2ae} /* (1, 20, 27) {real, imag} */,
  {32'hbd5a4bd8, 32'h40e47666} /* (1, 20, 26) {real, imag} */,
  {32'h406a6eaa, 32'h404685e2} /* (1, 20, 25) {real, imag} */,
  {32'hbf84349e, 32'h408b0e90} /* (1, 20, 24) {real, imag} */,
  {32'hbe468b90, 32'h410f451c} /* (1, 20, 23) {real, imag} */,
  {32'h3ef9500e, 32'h4113cc44} /* (1, 20, 22) {real, imag} */,
  {32'hbdd276e0, 32'h407d41a0} /* (1, 20, 21) {real, imag} */,
  {32'hbd7dae18, 32'hc083bd05} /* (1, 20, 20) {real, imag} */,
  {32'hbf89045e, 32'hc0c56495} /* (1, 20, 19) {real, imag} */,
  {32'h3e11b292, 32'hc09ceb59} /* (1, 20, 18) {real, imag} */,
  {32'h3e253054, 32'hc0feede6} /* (1, 20, 17) {real, imag} */,
  {32'hbe2f243e, 32'hc0f199a2} /* (1, 20, 16) {real, imag} */,
  {32'hc0403cc8, 32'hc0c78932} /* (1, 20, 15) {real, imag} */,
  {32'hbfe32829, 32'hc0938362} /* (1, 20, 14) {real, imag} */,
  {32'h403f2aed, 32'hc09919b5} /* (1, 20, 13) {real, imag} */,
  {32'h3f53d00d, 32'hc0b78a2a} /* (1, 20, 12) {real, imag} */,
  {32'h3fbd33c8, 32'hc0e99769} /* (1, 20, 11) {real, imag} */,
  {32'h40383e6c, 32'h3e527498} /* (1, 20, 10) {real, imag} */,
  {32'hbfcb085c, 32'h40d769b6} /* (1, 20, 9) {real, imag} */,
  {32'hc085760d, 32'h40d0e030} /* (1, 20, 8) {real, imag} */,
  {32'hbf3afd98, 32'h40ba4b7a} /* (1, 20, 7) {real, imag} */,
  {32'hbf8a2605, 32'h40de58f8} /* (1, 20, 6) {real, imag} */,
  {32'hbefa2e36, 32'h4073e354} /* (1, 20, 5) {real, imag} */,
  {32'hc00f44b8, 32'h40c8a28c} /* (1, 20, 4) {real, imag} */,
  {32'hc06b81ee, 32'h40f2d848} /* (1, 20, 3) {real, imag} */,
  {32'hbefd424e, 32'h409afaac} /* (1, 20, 2) {real, imag} */,
  {32'h3f5cb598, 32'h40d70775} /* (1, 20, 1) {real, imag} */,
  {32'hbef3cbc8, 32'h4096a236} /* (1, 20, 0) {real, imag} */,
  {32'hbc9630d0, 32'h407bb8d5} /* (1, 19, 31) {real, imag} */,
  {32'h3fe37603, 32'h41056942} /* (1, 19, 30) {real, imag} */,
  {32'h3f4c7f9b, 32'h410c3afc} /* (1, 19, 29) {real, imag} */,
  {32'h3f205430, 32'h40dcca6c} /* (1, 19, 28) {real, imag} */,
  {32'h3f5e1696, 32'h41049d56} /* (1, 19, 27) {real, imag} */,
  {32'h3da60492, 32'h411b5dde} /* (1, 19, 26) {real, imag} */,
  {32'h3f378110, 32'h40eb990b} /* (1, 19, 25) {real, imag} */,
  {32'hc01e067a, 32'h410ccb1c} /* (1, 19, 24) {real, imag} */,
  {32'hc05eeb97, 32'h4136d108} /* (1, 19, 23) {real, imag} */,
  {32'hbf9966bc, 32'h413269a9} /* (1, 19, 22) {real, imag} */,
  {32'hbf47a643, 32'h40ae22b4} /* (1, 19, 21) {real, imag} */,
  {32'hbe4c2715, 32'hc0c0486b} /* (1, 19, 20) {real, imag} */,
  {32'h3f8349da, 32'hc0f856de} /* (1, 19, 19) {real, imag} */,
  {32'h3eeb1b06, 32'hc0ece5dc} /* (1, 19, 18) {real, imag} */,
  {32'h3e09bc06, 32'hc1103b0c} /* (1, 19, 17) {real, imag} */,
  {32'h3fa45ca1, 32'hc11986dc} /* (1, 19, 16) {real, imag} */,
  {32'h3f8b2704, 32'hc112a94b} /* (1, 19, 15) {real, imag} */,
  {32'h3fabc60f, 32'hc10e1498} /* (1, 19, 14) {real, imag} */,
  {32'h403a4484, 32'hc10e77a2} /* (1, 19, 13) {real, imag} */,
  {32'h3ed7a569, 32'hc10ef5bc} /* (1, 19, 12) {real, imag} */,
  {32'h3fdad3c3, 32'hc0b0b13e} /* (1, 19, 11) {real, imag} */,
  {32'h4054c45e, 32'h40704152} /* (1, 19, 10) {real, imag} */,
  {32'hc00c6e47, 32'h40fd2a72} /* (1, 19, 9) {real, imag} */,
  {32'hc0937f48, 32'h41022e58} /* (1, 19, 8) {real, imag} */,
  {32'h3fc572c2, 32'h40f0e1a0} /* (1, 19, 7) {real, imag} */,
  {32'hbeb39ba6, 32'h40de984f} /* (1, 19, 6) {real, imag} */,
  {32'hbea370c8, 32'h40a76244} /* (1, 19, 5) {real, imag} */,
  {32'hbf2b83ce, 32'h40dce896} /* (1, 19, 4) {real, imag} */,
  {32'hbfe6ecbe, 32'h40e06f20} /* (1, 19, 3) {real, imag} */,
  {32'hc08ec1f2, 32'h40fce337} /* (1, 19, 2) {real, imag} */,
  {32'hc07f57f8, 32'h4109dcd8} /* (1, 19, 1) {real, imag} */,
  {32'hc01b893c, 32'h4096076c} /* (1, 19, 0) {real, imag} */,
  {32'hc02e05aa, 32'h40d7d3ec} /* (1, 18, 31) {real, imag} */,
  {32'hbfc7771e, 32'h412e4310} /* (1, 18, 30) {real, imag} */,
  {32'hbfcfc400, 32'h410eab25} /* (1, 18, 29) {real, imag} */,
  {32'hbf2d763a, 32'h40ef3e53} /* (1, 18, 28) {real, imag} */,
  {32'hbfb23210, 32'h40f24569} /* (1, 18, 27) {real, imag} */,
  {32'h3ed55cc6, 32'h40bdb049} /* (1, 18, 26) {real, imag} */,
  {32'hbfff5f19, 32'h41045102} /* (1, 18, 25) {real, imag} */,
  {32'hc05da901, 32'h4142c301} /* (1, 18, 24) {real, imag} */,
  {32'hc0493b3a, 32'h411a03d0} /* (1, 18, 23) {real, imag} */,
  {32'hbf1c67e2, 32'h40bce0bb} /* (1, 18, 22) {real, imag} */,
  {32'hbfd8c593, 32'h40477bb8} /* (1, 18, 21) {real, imag} */,
  {32'hbf90236e, 32'hc0df4f71} /* (1, 18, 20) {real, imag} */,
  {32'h400e0674, 32'hc10d33e7} /* (1, 18, 19) {real, imag} */,
  {32'h404a4b4c, 32'hc0f7513e} /* (1, 18, 18) {real, imag} */,
  {32'h402b95f7, 32'hc10ca71d} /* (1, 18, 17) {real, imag} */,
  {32'h407daee9, 32'hc113aacb} /* (1, 18, 16) {real, imag} */,
  {32'h40588684, 32'hc1181e53} /* (1, 18, 15) {real, imag} */,
  {32'h3fda4666, 32'hc1098ac7} /* (1, 18, 14) {real, imag} */,
  {32'hbee001f8, 32'hc104bf3b} /* (1, 18, 13) {real, imag} */,
  {32'hbe7d4ccc, 32'hc10873a7} /* (1, 18, 12) {real, imag} */,
  {32'hbdbf4df8, 32'hc07874e0} /* (1, 18, 11) {real, imag} */,
  {32'hbf5dec64, 32'h409c5292} /* (1, 18, 10) {real, imag} */,
  {32'hc09c6032, 32'h40e14d00} /* (1, 18, 9) {real, imag} */,
  {32'hc04da3f3, 32'h410a0147} /* (1, 18, 8) {real, imag} */,
  {32'h3fc7be50, 32'h41073c52} /* (1, 18, 7) {real, imag} */,
  {32'h3fd52d02, 32'h40e56285} /* (1, 18, 6) {real, imag} */,
  {32'h3fb098c0, 32'h40b5fa17} /* (1, 18, 5) {real, imag} */,
  {32'hbffa2733, 32'h40bb3274} /* (1, 18, 4) {real, imag} */,
  {32'hbf10115c, 32'h40da00dc} /* (1, 18, 3) {real, imag} */,
  {32'hc0134c64, 32'h411133ea} /* (1, 18, 2) {real, imag} */,
  {32'hc09237c4, 32'h411ef9f2} /* (1, 18, 1) {real, imag} */,
  {32'hc0842470, 32'h40d73eb0} /* (1, 18, 0) {real, imag} */,
  {32'hc04165c6, 32'h40a0467a} /* (1, 17, 31) {real, imag} */,
  {32'hc060d77a, 32'h41088456} /* (1, 17, 30) {real, imag} */,
  {32'hc02bf998, 32'h41118fb8} /* (1, 17, 29) {real, imag} */,
  {32'hbffc724a, 32'h411a50f0} /* (1, 17, 28) {real, imag} */,
  {32'hbf42c016, 32'h4111402b} /* (1, 17, 27) {real, imag} */,
  {32'h3f76793a, 32'h40c13cfd} /* (1, 17, 26) {real, imag} */,
  {32'hbfca35c0, 32'h4106ebaa} /* (1, 17, 25) {real, imag} */,
  {32'hc07d9fd3, 32'h41560c62} /* (1, 17, 24) {real, imag} */,
  {32'hbf1127e1, 32'h41360f7a} /* (1, 17, 23) {real, imag} */,
  {32'h3fb59523, 32'h40f2f5d8} /* (1, 17, 22) {real, imag} */,
  {32'hc027c148, 32'h3f9223f4} /* (1, 17, 21) {real, imag} */,
  {32'hbd2937f8, 32'hc0e02cb0} /* (1, 17, 20) {real, imag} */,
  {32'h3fa59d10, 32'hc10ed796} /* (1, 17, 19) {real, imag} */,
  {32'h3fbb5b02, 32'hc108b9b1} /* (1, 17, 18) {real, imag} */,
  {32'h3ff522f3, 32'hc0d13328} /* (1, 17, 17) {real, imag} */,
  {32'h401c6164, 32'hc0e436f7} /* (1, 17, 16) {real, imag} */,
  {32'h401bd18a, 32'hc10fc79b} /* (1, 17, 15) {real, imag} */,
  {32'h4081b80a, 32'hc1070308} /* (1, 17, 14) {real, imag} */,
  {32'h3f3a66b2, 32'hc109a9d6} /* (1, 17, 13) {real, imag} */,
  {32'h3feedef1, 32'hc126204a} /* (1, 17, 12) {real, imag} */,
  {32'h4014a9d6, 32'hc09a7202} /* (1, 17, 11) {real, imag} */,
  {32'h3f5dc6c2, 32'h408a7cd3} /* (1, 17, 10) {real, imag} */,
  {32'hc0155ab7, 32'h410b81f2} /* (1, 17, 9) {real, imag} */,
  {32'hc04ebca3, 32'h410b3a62} /* (1, 17, 8) {real, imag} */,
  {32'h3eb761f2, 32'h41129218} /* (1, 17, 7) {real, imag} */,
  {32'h4097bc86, 32'h41274ca6} /* (1, 17, 6) {real, imag} */,
  {32'h401aaf5c, 32'h4107c71e} /* (1, 17, 5) {real, imag} */,
  {32'hbf907c2c, 32'h4106dc6e} /* (1, 17, 4) {real, imag} */,
  {32'hbf417ad5, 32'h4116b366} /* (1, 17, 3) {real, imag} */,
  {32'hc030958c, 32'h41127ed8} /* (1, 17, 2) {real, imag} */,
  {32'hc065a9b6, 32'h41143c0c} /* (1, 17, 1) {real, imag} */,
  {32'hbffe9d73, 32'h40c6f233} /* (1, 17, 0) {real, imag} */,
  {32'hbf7a5aaa, 32'h40921fdc} /* (1, 16, 31) {real, imag} */,
  {32'hbff52826, 32'h41270204} /* (1, 16, 30) {real, imag} */,
  {32'hc0409d46, 32'h4113d9e2} /* (1, 16, 29) {real, imag} */,
  {32'hc00f2c4c, 32'h411ad5be} /* (1, 16, 28) {real, imag} */,
  {32'hbfac1d2f, 32'h410fe8da} /* (1, 16, 27) {real, imag} */,
  {32'h3d6db3b0, 32'h40dd3190} /* (1, 16, 26) {real, imag} */,
  {32'hbf78c02e, 32'h40fe75fe} /* (1, 16, 25) {real, imag} */,
  {32'hc05802f7, 32'h41293d70} /* (1, 16, 24) {real, imag} */,
  {32'h3f58b67a, 32'h412b7ec6} /* (1, 16, 23) {real, imag} */,
  {32'h406aad8c, 32'h41129095} /* (1, 16, 22) {real, imag} */,
  {32'h3edd5f60, 32'hbe93ca03} /* (1, 16, 21) {real, imag} */,
  {32'h4023c096, 32'hc107dafa} /* (1, 16, 20) {real, imag} */,
  {32'h402bdaf6, 32'hc115cd5e} /* (1, 16, 19) {real, imag} */,
  {32'h3f60c905, 32'hc119b166} /* (1, 16, 18) {real, imag} */,
  {32'h3e056dda, 32'hc0fb6ccb} /* (1, 16, 17) {real, imag} */,
  {32'hbecef594, 32'hc0dfead1} /* (1, 16, 16) {real, imag} */,
  {32'h3fa2878e, 32'hc0dd9b53} /* (1, 16, 15) {real, imag} */,
  {32'h403eb18e, 32'hc121c4c8} /* (1, 16, 14) {real, imag} */,
  {32'h40172034, 32'hc12c2200} /* (1, 16, 13) {real, imag} */,
  {32'h400d3368, 32'hc1146def} /* (1, 16, 12) {real, imag} */,
  {32'h3f0889ac, 32'hc0b2d5ad} /* (1, 16, 11) {real, imag} */,
  {32'hbfb556fb, 32'h404e6c68} /* (1, 16, 10) {real, imag} */,
  {32'hbfadb7ad, 32'h410c525c} /* (1, 16, 9) {real, imag} */,
  {32'hbfc6b589, 32'h40d83e4b} /* (1, 16, 8) {real, imag} */,
  {32'h3f8dbefe, 32'h40f82cce} /* (1, 16, 7) {real, imag} */,
  {32'h3fefbc3b, 32'h410b4106} /* (1, 16, 6) {real, imag} */,
  {32'hbf1dce0d, 32'h40df07f2} /* (1, 16, 5) {real, imag} */,
  {32'hc012db1f, 32'h4104d541} /* (1, 16, 4) {real, imag} */,
  {32'hbfda21cf, 32'h412a455b} /* (1, 16, 3) {real, imag} */,
  {32'hbfe8ac0c, 32'h4128af99} /* (1, 16, 2) {real, imag} */,
  {32'hc031fef1, 32'h41165ca4} /* (1, 16, 1) {real, imag} */,
  {32'h3ee91d0c, 32'h4087d8d1} /* (1, 16, 0) {real, imag} */,
  {32'hbd19c1b0, 32'h40890dca} /* (1, 15, 31) {real, imag} */,
  {32'hbfa56b4a, 32'h411bfe10} /* (1, 15, 30) {real, imag} */,
  {32'hbf957958, 32'h4117d5aa} /* (1, 15, 29) {real, imag} */,
  {32'h3eb9fda3, 32'h41275287} /* (1, 15, 28) {real, imag} */,
  {32'hbb86f240, 32'h411bb30a} /* (1, 15, 27) {real, imag} */,
  {32'hbefed505, 32'h4117b846} /* (1, 15, 26) {real, imag} */,
  {32'hbfd9f66c, 32'h4105983e} /* (1, 15, 25) {real, imag} */,
  {32'hbf818f1a, 32'h4111d680} /* (1, 15, 24) {real, imag} */,
  {32'h401c40ad, 32'h411f98ec} /* (1, 15, 23) {real, imag} */,
  {32'h3eb8ec8f, 32'h408dd8d0} /* (1, 15, 22) {real, imag} */,
  {32'hbfcaa4a8, 32'hc01a12ef} /* (1, 15, 21) {real, imag} */,
  {32'h3fa8eb14, 32'hc117e0bf} /* (1, 15, 20) {real, imag} */,
  {32'h4037f2a8, 32'hc11848be} /* (1, 15, 19) {real, imag} */,
  {32'h3fa32266, 32'hc11be3b0} /* (1, 15, 18) {real, imag} */,
  {32'h3eb40f39, 32'hc12d92f6} /* (1, 15, 17) {real, imag} */,
  {32'h3fc652d4, 32'hc12757ec} /* (1, 15, 16) {real, imag} */,
  {32'h400ca3d6, 32'hc0d78a16} /* (1, 15, 15) {real, imag} */,
  {32'h3fccb0b6, 32'hc0f4397a} /* (1, 15, 14) {real, imag} */,
  {32'h3e645052, 32'hc0f79099} /* (1, 15, 13) {real, imag} */,
  {32'h3d7dc440, 32'hc109623e} /* (1, 15, 12) {real, imag} */,
  {32'h3f3be06f, 32'hc0e29e0a} /* (1, 15, 11) {real, imag} */,
  {32'hc0443a75, 32'h3f69b30c} /* (1, 15, 10) {real, imag} */,
  {32'hc047ca22, 32'h40be3c86} /* (1, 15, 9) {real, imag} */,
  {32'hc0350eda, 32'h40eed412} /* (1, 15, 8) {real, imag} */,
  {32'hc002bccc, 32'h4107e1f7} /* (1, 15, 7) {real, imag} */,
  {32'h3f24d2ab, 32'h40e165ce} /* (1, 15, 6) {real, imag} */,
  {32'hbfb43ff0, 32'h4093353b} /* (1, 15, 5) {real, imag} */,
  {32'hc041c6c8, 32'h411a84fc} /* (1, 15, 4) {real, imag} */,
  {32'hc0850986, 32'h413fa0b4} /* (1, 15, 3) {real, imag} */,
  {32'hbebca06a, 32'h413a2cc4} /* (1, 15, 2) {real, imag} */,
  {32'h3eecd992, 32'h412ab2d8} /* (1, 15, 1) {real, imag} */,
  {32'h4008da78, 32'h40bff4ea} /* (1, 15, 0) {real, imag} */,
  {32'h3f28feae, 32'h4061de68} /* (1, 14, 31) {real, imag} */,
  {32'hbf10f828, 32'h40eabbc5} /* (1, 14, 30) {real, imag} */,
  {32'hbeb062c6, 32'h40ee178b} /* (1, 14, 29) {real, imag} */,
  {32'h3fd641c0, 32'h41103554} /* (1, 14, 28) {real, imag} */,
  {32'h4022f844, 32'h411738cf} /* (1, 14, 27) {real, imag} */,
  {32'h3f37dd46, 32'h411aa0f4} /* (1, 14, 26) {real, imag} */,
  {32'hc01a65f6, 32'h4115cd2a} /* (1, 14, 25) {real, imag} */,
  {32'hc08410ba, 32'h410657b0} /* (1, 14, 24) {real, imag} */,
  {32'hbfdf4b53, 32'h41223cf4} /* (1, 14, 23) {real, imag} */,
  {32'hc05aed4f, 32'h40cd0939} /* (1, 14, 22) {real, imag} */,
  {32'hbf4e51a6, 32'h40108f1b} /* (1, 14, 21) {real, imag} */,
  {32'h3ff6c0dd, 32'hc0a9566a} /* (1, 14, 20) {real, imag} */,
  {32'h400e223b, 32'hc0b38851} /* (1, 14, 19) {real, imag} */,
  {32'hbef0f788, 32'hc0ae98c4} /* (1, 14, 18) {real, imag} */,
  {32'hc041aff3, 32'hc0d993bd} /* (1, 14, 17) {real, imag} */,
  {32'h3f299fc0, 32'hc0f547ee} /* (1, 14, 16) {real, imag} */,
  {32'h3fdfe74a, 32'hc0e74d17} /* (1, 14, 15) {real, imag} */,
  {32'h4003bb65, 32'hc0fc7bc9} /* (1, 14, 14) {real, imag} */,
  {32'hbed3bbda, 32'hc10c748a} /* (1, 14, 13) {real, imag} */,
  {32'h3f12d1e7, 32'hc10b8ef0} /* (1, 14, 12) {real, imag} */,
  {32'h3de40668, 32'hc0fcff2c} /* (1, 14, 11) {real, imag} */,
  {32'hbfc3feb3, 32'h3f971177} /* (1, 14, 10) {real, imag} */,
  {32'hc04a731e, 32'h40dc35cf} /* (1, 14, 9) {real, imag} */,
  {32'hc02d8f33, 32'h4108eb47} /* (1, 14, 8) {real, imag} */,
  {32'hbe15e6f0, 32'h41267d56} /* (1, 14, 7) {real, imag} */,
  {32'h4005c1e4, 32'h41042dc8} /* (1, 14, 6) {real, imag} */,
  {32'hbeb40918, 32'h40ce37f4} /* (1, 14, 5) {real, imag} */,
  {32'hbefc74d8, 32'h411d2347} /* (1, 14, 4) {real, imag} */,
  {32'hbfaa32b5, 32'h4105ef56} /* (1, 14, 3) {real, imag} */,
  {32'hbcad1260, 32'h40ff93b4} /* (1, 14, 2) {real, imag} */,
  {32'h40298d1e, 32'h413adda3} /* (1, 14, 1) {real, imag} */,
  {32'h405292ca, 32'h40fc16d0} /* (1, 14, 0) {real, imag} */,
  {32'hbf20e0f0, 32'h40821875} /* (1, 13, 31) {real, imag} */,
  {32'h3f07f2dc, 32'h4108984d} /* (1, 13, 30) {real, imag} */,
  {32'h3f952d84, 32'h40d588c8} /* (1, 13, 29) {real, imag} */,
  {32'h4000db60, 32'h4117d4b2} /* (1, 13, 28) {real, imag} */,
  {32'h3fca6a8a, 32'h411ddd7a} /* (1, 13, 27) {real, imag} */,
  {32'hbebb15f8, 32'h40cd96a6} /* (1, 13, 26) {real, imag} */,
  {32'hbfac1539, 32'h40bf48a5} /* (1, 13, 25) {real, imag} */,
  {32'hc0147e7e, 32'h410be176} /* (1, 13, 24) {real, imag} */,
  {32'hbed43dfd, 32'h4131faee} /* (1, 13, 23) {real, imag} */,
  {32'hbe542db4, 32'h4116dde6} /* (1, 13, 22) {real, imag} */,
  {32'hbf15e04a, 32'h405cfb9f} /* (1, 13, 21) {real, imag} */,
  {32'hbe8b2d31, 32'hc09273e5} /* (1, 13, 20) {real, imag} */,
  {32'hbe9e2841, 32'hc0df469a} /* (1, 13, 19) {real, imag} */,
  {32'hbfc3a9a0, 32'hc0b3318c} /* (1, 13, 18) {real, imag} */,
  {32'hbfd6f9e6, 32'hc0b331a8} /* (1, 13, 17) {real, imag} */,
  {32'hbf4d8127, 32'hc0d97f05} /* (1, 13, 16) {real, imag} */,
  {32'h3fe62839, 32'hc0ffab5b} /* (1, 13, 15) {real, imag} */,
  {32'h400d7a6d, 32'hc0d916be} /* (1, 13, 14) {real, imag} */,
  {32'h40154680, 32'hc105298b} /* (1, 13, 13) {real, imag} */,
  {32'h3f3f9810, 32'hc10b659c} /* (1, 13, 12) {real, imag} */,
  {32'hbf8b6178, 32'hc0fe9376} /* (1, 13, 11) {real, imag} */,
  {32'hc01aba80, 32'h407f618f} /* (1, 13, 10) {real, imag} */,
  {32'hc0b6b01a, 32'h412c065b} /* (1, 13, 9) {real, imag} */,
  {32'hc0cae482, 32'h410c086c} /* (1, 13, 8) {real, imag} */,
  {32'hbe814249, 32'h4116fb9c} /* (1, 13, 7) {real, imag} */,
  {32'h3f520e64, 32'h41206a44} /* (1, 13, 6) {real, imag} */,
  {32'hc004e79f, 32'h412dd538} /* (1, 13, 5) {real, imag} */,
  {32'hc02f15f2, 32'h4128e182} /* (1, 13, 4) {real, imag} */,
  {32'hc0539854, 32'h40fadf48} /* (1, 13, 3) {real, imag} */,
  {32'hbf08759e, 32'h4081938a} /* (1, 13, 2) {real, imag} */,
  {32'h3ff495f3, 32'h40eab581} /* (1, 13, 1) {real, imag} */,
  {32'h3fe6ed38, 32'h40ba5245} /* (1, 13, 0) {real, imag} */,
  {32'hbf3fe50a, 32'h409f9b2b} /* (1, 12, 31) {real, imag} */,
  {32'h3fa3f1e2, 32'h411259cf} /* (1, 12, 30) {real, imag} */,
  {32'h40621f46, 32'h40eca033} /* (1, 12, 29) {real, imag} */,
  {32'h3fe4b9b4, 32'h41193717} /* (1, 12, 28) {real, imag} */,
  {32'hc062fdda, 32'h410aef92} /* (1, 12, 27) {real, imag} */,
  {32'hc0a49f72, 32'h40edb72b} /* (1, 12, 26) {real, imag} */,
  {32'hc0021522, 32'h40c2e610} /* (1, 12, 25) {real, imag} */,
  {32'h3ffdee3a, 32'h411d279a} /* (1, 12, 24) {real, imag} */,
  {32'h3e87a363, 32'h412eb661} /* (1, 12, 23) {real, imag} */,
  {32'hc033a2ca, 32'h41008246} /* (1, 12, 22) {real, imag} */,
  {32'hc03d812c, 32'h406885c2} /* (1, 12, 21) {real, imag} */,
  {32'hbfdf26b8, 32'hc0c4e545} /* (1, 12, 20) {real, imag} */,
  {32'hbdc47dec, 32'hc1183002} /* (1, 12, 19) {real, imag} */,
  {32'h3e30a54a, 32'hc10630f4} /* (1, 12, 18) {real, imag} */,
  {32'hbdd92cfc, 32'hc11ba262} /* (1, 12, 17) {real, imag} */,
  {32'h3dd3a6b4, 32'hc11f7072} /* (1, 12, 16) {real, imag} */,
  {32'h403a7d75, 32'hc111a9e0} /* (1, 12, 15) {real, imag} */,
  {32'h408616af, 32'hc0d174df} /* (1, 12, 14) {real, imag} */,
  {32'h4072c05e, 32'hc0fd651b} /* (1, 12, 13) {real, imag} */,
  {32'h3ed5f730, 32'hc134dc68} /* (1, 12, 12) {real, imag} */,
  {32'hbf81c814, 32'hc0d4b932} /* (1, 12, 11) {real, imag} */,
  {32'hbf6ee4f4, 32'h40efd7de} /* (1, 12, 10) {real, imag} */,
  {32'hc05cf7bb, 32'h4135f8b8} /* (1, 12, 9) {real, imag} */,
  {32'hc094bdd4, 32'h410ed303} /* (1, 12, 8) {real, imag} */,
  {32'hbf7633db, 32'h410e799e} /* (1, 12, 7) {real, imag} */,
  {32'hbf1baeef, 32'h41240bac} /* (1, 12, 6) {real, imag} */,
  {32'hbfa79fc0, 32'h411b9be8} /* (1, 12, 5) {real, imag} */,
  {32'hbf8d1397, 32'h40ec5399} /* (1, 12, 4) {real, imag} */,
  {32'hc0069d0e, 32'h40a187d2} /* (1, 12, 3) {real, imag} */,
  {32'hbfc67b62, 32'h405f943c} /* (1, 12, 2) {real, imag} */,
  {32'hbf163cf4, 32'h40500ec0} /* (1, 12, 1) {real, imag} */,
  {32'hbee26648, 32'h40143ec8} /* (1, 12, 0) {real, imag} */,
  {32'hbf20baa1, 32'h4027db46} /* (1, 11, 31) {real, imag} */,
  {32'hbfc0e177, 32'h40bc74d6} /* (1, 11, 30) {real, imag} */,
  {32'h3db7341e, 32'h40951eff} /* (1, 11, 29) {real, imag} */,
  {32'hbebe8073, 32'h40c7fc07} /* (1, 11, 28) {real, imag} */,
  {32'hbfea5576, 32'h40d4d02c} /* (1, 11, 27) {real, imag} */,
  {32'hbfda9fde, 32'h40e19714} /* (1, 11, 26) {real, imag} */,
  {32'hc005d541, 32'h40cd2d56} /* (1, 11, 25) {real, imag} */,
  {32'h3fc10c3b, 32'h4126fbbc} /* (1, 11, 24) {real, imag} */,
  {32'h4002fcf8, 32'h410cee31} /* (1, 11, 23) {real, imag} */,
  {32'hc04c228b, 32'h40cb10c4} /* (1, 11, 22) {real, imag} */,
  {32'hc0169eaa, 32'h3fc384ee} /* (1, 11, 21) {real, imag} */,
  {32'hbe29b734, 32'hc0a13f68} /* (1, 11, 20) {real, imag} */,
  {32'h3e2fbe7c, 32'hc0a3d17c} /* (1, 11, 19) {real, imag} */,
  {32'hbdeb72f8, 32'hc06a36ab} /* (1, 11, 18) {real, imag} */,
  {32'hbe4e2150, 32'hc0a3f6dc} /* (1, 11, 17) {real, imag} */,
  {32'h3ec7fbac, 32'hc0c358cc} /* (1, 11, 16) {real, imag} */,
  {32'h3f2983e0, 32'hc0992c89} /* (1, 11, 15) {real, imag} */,
  {32'h3fb78725, 32'hc09e1e6d} /* (1, 11, 14) {real, imag} */,
  {32'hbe063a0c, 32'hc0af94b9} /* (1, 11, 13) {real, imag} */,
  {32'hc02e197a, 32'hc0fd8164} /* (1, 11, 12) {real, imag} */,
  {32'hc07edc3f, 32'hc0a62986} /* (1, 11, 11) {real, imag} */,
  {32'hbfaedca6, 32'h4076f4e9} /* (1, 11, 10) {real, imag} */,
  {32'hbfa75016, 32'h40d275df} /* (1, 11, 9) {real, imag} */,
  {32'hbf663456, 32'h410863da} /* (1, 11, 8) {real, imag} */,
  {32'h3fb5c943, 32'h4112fb07} /* (1, 11, 7) {real, imag} */,
  {32'hbf1a50ea, 32'h41111db4} /* (1, 11, 6) {real, imag} */,
  {32'hc03d2eba, 32'h40c3a51f} /* (1, 11, 5) {real, imag} */,
  {32'h3f9f0ea7, 32'h40960568} /* (1, 11, 4) {real, imag} */,
  {32'hc01065a4, 32'h400e7c6b} /* (1, 11, 3) {real, imag} */,
  {32'hc09bc2ca, 32'h40be0f4d} /* (1, 11, 2) {real, imag} */,
  {32'hc013b5bb, 32'h409fb3d5} /* (1, 11, 1) {real, imag} */,
  {32'hbf3118e4, 32'h3fdc0b74} /* (1, 11, 0) {real, imag} */,
  {32'h3f843d40, 32'hc0069f0e} /* (1, 10, 31) {real, imag} */,
  {32'hbe3d032f, 32'hc084fd73} /* (1, 10, 30) {real, imag} */,
  {32'hc01613f4, 32'hc0e67c36} /* (1, 10, 29) {real, imag} */,
  {32'hbfcf2840, 32'hc0be9a84} /* (1, 10, 28) {real, imag} */,
  {32'h3feef866, 32'hc0ad64e1} /* (1, 10, 27) {real, imag} */,
  {32'h3ef844be, 32'hbfeff1dc} /* (1, 10, 26) {real, imag} */,
  {32'h3fc2bbbb, 32'hbfa5d730} /* (1, 10, 25) {real, imag} */,
  {32'h4037e6eb, 32'hbe324d15} /* (1, 10, 24) {real, imag} */,
  {32'h408e39c4, 32'hc06f3758} /* (1, 10, 23) {real, imag} */,
  {32'h3e1187ac, 32'hc0959077} /* (1, 10, 22) {real, imag} */,
  {32'hbfcee815, 32'hc08a685e} /* (1, 10, 21) {real, imag} */,
  {32'hbf5804b3, 32'h3f4316f2} /* (1, 10, 20) {real, imag} */,
  {32'h3f3c6314, 32'h4094a474} /* (1, 10, 19) {real, imag} */,
  {32'h3ea907a6, 32'h40cb15e5} /* (1, 10, 18) {real, imag} */,
  {32'hc001d244, 32'h408e8a75} /* (1, 10, 17) {real, imag} */,
  {32'hbf6039f8, 32'h40f17913} /* (1, 10, 16) {real, imag} */,
  {32'hc06de258, 32'h40c12574} /* (1, 10, 15) {real, imag} */,
  {32'hc00f7250, 32'h4031eaa6} /* (1, 10, 14) {real, imag} */,
  {32'hbff1f4d7, 32'h4035bfcb} /* (1, 10, 13) {real, imag} */,
  {32'hc042b2ec, 32'h405699fa} /* (1, 10, 12) {real, imag} */,
  {32'hbe499ef2, 32'h402aa641} /* (1, 10, 11) {real, imag} */,
  {32'h3fa0e8fa, 32'h3f413653} /* (1, 10, 10) {real, imag} */,
  {32'h4002db33, 32'hc01cfb4c} /* (1, 10, 9) {real, imag} */,
  {32'h3f286e0d, 32'hbfaaeef5} /* (1, 10, 8) {real, imag} */,
  {32'h3fef621c, 32'hbfbf19fe} /* (1, 10, 7) {real, imag} */,
  {32'h3ffbeb9e, 32'hc0137c6c} /* (1, 10, 6) {real, imag} */,
  {32'hbeb14d5c, 32'hc09e82d6} /* (1, 10, 5) {real, imag} */,
  {32'h40217930, 32'hc09dc264} /* (1, 10, 4) {real, imag} */,
  {32'hbfb96968, 32'hc0c26433} /* (1, 10, 3) {real, imag} */,
  {32'hc03e3f00, 32'hbf400d3a} /* (1, 10, 2) {real, imag} */,
  {32'hc002995c, 32'hc0063c94} /* (1, 10, 1) {real, imag} */,
  {32'hbcbd1688, 32'hc01c0571} /* (1, 10, 0) {real, imag} */,
  {32'h3fdfc816, 32'hc03ce72d} /* (1, 9, 31) {real, imag} */,
  {32'h4050d0f0, 32'hc0b4caac} /* (1, 9, 30) {real, imag} */,
  {32'h3fbe5b68, 32'hc11293d5} /* (1, 9, 29) {real, imag} */,
  {32'hbf33d006, 32'hc129b5a3} /* (1, 9, 28) {real, imag} */,
  {32'h3fbd2496, 32'hc1408898} /* (1, 9, 27) {real, imag} */,
  {32'hbd9c17cc, 32'hc10d5694} /* (1, 9, 26) {real, imag} */,
  {32'h3fd3980a, 32'hc0f1bf3f} /* (1, 9, 25) {real, imag} */,
  {32'h3fa2cb2c, 32'hc101a3bb} /* (1, 9, 24) {real, imag} */,
  {32'h3fea7170, 32'hc10dd6c4} /* (1, 9, 23) {real, imag} */,
  {32'h3fdb4699, 32'hc0eeb038} /* (1, 9, 22) {real, imag} */,
  {32'hbf03999a, 32'hc0bfef7d} /* (1, 9, 21) {real, imag} */,
  {32'hc0077152, 32'h403c8507} /* (1, 9, 20) {real, imag} */,
  {32'hbe8f7a25, 32'h40bea81a} /* (1, 9, 19) {real, imag} */,
  {32'hbf5e1bba, 32'h411cb8fa} /* (1, 9, 18) {real, imag} */,
  {32'hc0972cc4, 32'h41120f44} /* (1, 9, 17) {real, imag} */,
  {32'hc08bd0bc, 32'h41227f9c} /* (1, 9, 16) {real, imag} */,
  {32'hc082e936, 32'h4112c55c} /* (1, 9, 15) {real, imag} */,
  {32'hc02e7350, 32'h4117892b} /* (1, 9, 14) {real, imag} */,
  {32'hbf98745d, 32'h4103e816} /* (1, 9, 13) {real, imag} */,
  {32'h3f43de2d, 32'h40b8a6c2} /* (1, 9, 12) {real, imag} */,
  {32'h402cf976, 32'h409a5275} /* (1, 9, 11) {real, imag} */,
  {32'h4001081c, 32'hbfad21f4} /* (1, 9, 10) {real, imag} */,
  {32'h408144f9, 32'hc0bab180} /* (1, 9, 9) {real, imag} */,
  {32'h3ff0a9a0, 32'hc10db0f2} /* (1, 9, 8) {real, imag} */,
  {32'h402770ad, 32'hc12d8f0a} /* (1, 9, 7) {real, imag} */,
  {32'h3ff77dde, 32'hc10e7b98} /* (1, 9, 6) {real, imag} */,
  {32'h3fd34f43, 32'hc1062826} /* (1, 9, 5) {real, imag} */,
  {32'h404acd6c, 32'hc0e69190} /* (1, 9, 4) {real, imag} */,
  {32'hbf1fa756, 32'hc1045453} /* (1, 9, 3) {real, imag} */,
  {32'hc008b703, 32'hc0be14c8} /* (1, 9, 2) {real, imag} */,
  {32'h3f73b32e, 32'hc0eec5d1} /* (1, 9, 1) {real, imag} */,
  {32'h3ffdbf93, 32'hc0a34e83} /* (1, 9, 0) {real, imag} */,
  {32'h4027cd70, 32'hc038bf84} /* (1, 8, 31) {real, imag} */,
  {32'h405c52f6, 32'hc0aefd8f} /* (1, 8, 30) {real, imag} */,
  {32'h405b55b9, 32'hc119d27e} /* (1, 8, 29) {real, imag} */,
  {32'hbe2daeda, 32'hc11887ac} /* (1, 8, 28) {real, imag} */,
  {32'h3f1b811b, 32'hc11718e2} /* (1, 8, 27) {real, imag} */,
  {32'h3f84a788, 32'hc11150d2} /* (1, 8, 26) {real, imag} */,
  {32'h3f35a4e5, 32'hc0f639eb} /* (1, 8, 25) {real, imag} */,
  {32'hc02531ea, 32'hc130ed38} /* (1, 8, 24) {real, imag} */,
  {32'h3d77d3d8, 32'hc130ba5b} /* (1, 8, 23) {real, imag} */,
  {32'h3fdb96bd, 32'hc10bc3a4} /* (1, 8, 22) {real, imag} */,
  {32'h3f982473, 32'hc095df1f} /* (1, 8, 21) {real, imag} */,
  {32'hbf1bc038, 32'h408d9e5c} /* (1, 8, 20) {real, imag} */,
  {32'hbf298b52, 32'h409617bb} /* (1, 8, 19) {real, imag} */,
  {32'hbfa12b4c, 32'h40be806e} /* (1, 8, 18) {real, imag} */,
  {32'hc0345bec, 32'h40e9dcf4} /* (1, 8, 17) {real, imag} */,
  {32'hc01f5393, 32'h41020708} /* (1, 8, 16) {real, imag} */,
  {32'hbf1a0160, 32'h412386b8} /* (1, 8, 15) {real, imag} */,
  {32'hc08dab9e, 32'h4113baf7} /* (1, 8, 14) {real, imag} */,
  {32'hc097d45d, 32'h40fce002} /* (1, 8, 13) {real, imag} */,
  {32'hbff9171a, 32'h40b57cf9} /* (1, 8, 12) {real, imag} */,
  {32'hbfc1dc15, 32'h40a58d4c} /* (1, 8, 11) {real, imag} */,
  {32'hbfba5338, 32'hbfa65716} /* (1, 8, 10) {real, imag} */,
  {32'h3f350172, 32'hc0826c68} /* (1, 8, 9) {real, imag} */,
  {32'hbec8a572, 32'hc1119ac8} /* (1, 8, 8) {real, imag} */,
  {32'hbeb152bb, 32'hc1335012} /* (1, 8, 7) {real, imag} */,
  {32'hbe78b661, 32'hc112e9d0} /* (1, 8, 6) {real, imag} */,
  {32'h3e98b813, 32'hc0ea2b75} /* (1, 8, 5) {real, imag} */,
  {32'h4005d022, 32'hc0b5fc8a} /* (1, 8, 4) {real, imag} */,
  {32'h3fc76e66, 32'hc0c265c5} /* (1, 8, 3) {real, imag} */,
  {32'h3f6f2e06, 32'hc1023619} /* (1, 8, 2) {real, imag} */,
  {32'h403c7b13, 32'hc101336f} /* (1, 8, 1) {real, imag} */,
  {32'h405afba6, 32'hc08339b8} /* (1, 8, 0) {real, imag} */,
  {32'h40708508, 32'hc0912fd6} /* (1, 7, 31) {real, imag} */,
  {32'h407bd172, 32'hc1014d50} /* (1, 7, 30) {real, imag} */,
  {32'h3f74b5d5, 32'hc130b132} /* (1, 7, 29) {real, imag} */,
  {32'hbfd22eed, 32'hc10dc78c} /* (1, 7, 28) {real, imag} */,
  {32'hbf3e3fa4, 32'hc0dbf53a} /* (1, 7, 27) {real, imag} */,
  {32'hbf2958d6, 32'hc0a948de} /* (1, 7, 26) {real, imag} */,
  {32'h404554f8, 32'hc0ae2e47} /* (1, 7, 25) {real, imag} */,
  {32'h3e835d62, 32'hc106c0da} /* (1, 7, 24) {real, imag} */,
  {32'h3fc40c41, 32'hc12183df} /* (1, 7, 23) {real, imag} */,
  {32'h3f8463e2, 32'hc140a466} /* (1, 7, 22) {real, imag} */,
  {32'h4052ed34, 32'hc0cdc551} /* (1, 7, 21) {real, imag} */,
  {32'h4046737f, 32'h40ac01a3} /* (1, 7, 20) {real, imag} */,
  {32'hbfe0080a, 32'h40f09e44} /* (1, 7, 19) {real, imag} */,
  {32'hbf9810cf, 32'h40e12830} /* (1, 7, 18) {real, imag} */,
  {32'hbefa420c, 32'h40bdd6d2} /* (1, 7, 17) {real, imag} */,
  {32'h3ef70f4d, 32'h40ff00b0} /* (1, 7, 16) {real, imag} */,
  {32'h3fb1deb0, 32'h411c1faa} /* (1, 7, 15) {real, imag} */,
  {32'hbee8e36c, 32'h410eaa6c} /* (1, 7, 14) {real, imag} */,
  {32'hc00caf5c, 32'h41089bd8} /* (1, 7, 13) {real, imag} */,
  {32'hbf902b00, 32'h4115dccc} /* (1, 7, 12) {real, imag} */,
  {32'hc086abbc, 32'h40c3ac6c} /* (1, 7, 11) {real, imag} */,
  {32'hbfec6974, 32'hc032def3} /* (1, 7, 10) {real, imag} */,
  {32'h3ff8d2ce, 32'hc0cfcc14} /* (1, 7, 9) {real, imag} */,
  {32'h3fc13a96, 32'hc146d839} /* (1, 7, 8) {real, imag} */,
  {32'hbff76513, 32'hc12308bd} /* (1, 7, 7) {real, imag} */,
  {32'hbe17a84a, 32'hc107c88a} /* (1, 7, 6) {real, imag} */,
  {32'h3f936704, 32'hc10082c6} /* (1, 7, 5) {real, imag} */,
  {32'hbdcd8728, 32'hc0f57e3c} /* (1, 7, 4) {real, imag} */,
  {32'h3f192e3e, 32'hc0ff0e87} /* (1, 7, 3) {real, imag} */,
  {32'h402b813f, 32'hc1225155} /* (1, 7, 2) {real, imag} */,
  {32'h3f8e8706, 32'hc10a5a69} /* (1, 7, 1) {real, imag} */,
  {32'h3fbe68c6, 32'hc056ae7a} /* (1, 7, 0) {real, imag} */,
  {32'h4022da9c, 32'hc071531d} /* (1, 6, 31) {real, imag} */,
  {32'h40858d79, 32'hc0b30a10} /* (1, 6, 30) {real, imag} */,
  {32'h403cda72, 32'hc0a85978} /* (1, 6, 29) {real, imag} */,
  {32'hbfaa41f7, 32'hc0fe21d4} /* (1, 6, 28) {real, imag} */,
  {32'hc02f5306, 32'hc0e3b088} /* (1, 6, 27) {real, imag} */,
  {32'hbfc92da8, 32'hc0ade30a} /* (1, 6, 26) {real, imag} */,
  {32'h4047cfee, 32'hc0b2d036} /* (1, 6, 25) {real, imag} */,
  {32'h3fe0ff50, 32'hc0fc36c4} /* (1, 6, 24) {real, imag} */,
  {32'h4001fcf9, 32'hc10dbc8b} /* (1, 6, 23) {real, imag} */,
  {32'h401cced0, 32'hc12156eb} /* (1, 6, 22) {real, imag} */,
  {32'h400c3eb0, 32'hc0c09188} /* (1, 6, 21) {real, imag} */,
  {32'h3f01108c, 32'h40a4cf48} /* (1, 6, 20) {real, imag} */,
  {32'hc0157938, 32'h40d9989a} /* (1, 6, 19) {real, imag} */,
  {32'hbfbaa637, 32'h410b42ac} /* (1, 6, 18) {real, imag} */,
  {32'hbf8d2f14, 32'h40ea42f3} /* (1, 6, 17) {real, imag} */,
  {32'hbf1bdf41, 32'h410b8f82} /* (1, 6, 16) {real, imag} */,
  {32'hc0321f02, 32'h412446ae} /* (1, 6, 15) {real, imag} */,
  {32'hbf8fd547, 32'h4118385c} /* (1, 6, 14) {real, imag} */,
  {32'hbff34b9f, 32'h410c337a} /* (1, 6, 13) {real, imag} */,
  {32'h3f40d9f9, 32'h412b8bee} /* (1, 6, 12) {real, imag} */,
  {32'hbfb59126, 32'h40b92f58} /* (1, 6, 11) {real, imag} */,
  {32'h3f7d7424, 32'hc007c224} /* (1, 6, 10) {real, imag} */,
  {32'h404ce793, 32'hc09f818e} /* (1, 6, 9) {real, imag} */,
  {32'hbe8dc1c5, 32'hc120a8f8} /* (1, 6, 8) {real, imag} */,
  {32'hbefb9ee4, 32'hc0d88214} /* (1, 6, 7) {real, imag} */,
  {32'h3f930089, 32'hc10c0fc8} /* (1, 6, 6) {real, imag} */,
  {32'h401346b8, 32'hc11b1547} /* (1, 6, 5) {real, imag} */,
  {32'h3fa43282, 32'hc100d77b} /* (1, 6, 4) {real, imag} */,
  {32'h3fe83424, 32'hc11389c0} /* (1, 6, 3) {real, imag} */,
  {32'h4040378a, 32'hc115583c} /* (1, 6, 2) {real, imag} */,
  {32'h40000662, 32'hc116bed8} /* (1, 6, 1) {real, imag} */,
  {32'h3f1ff264, 32'hc094184c} /* (1, 6, 0) {real, imag} */,
  {32'h3f8db188, 32'hc0b7c7e2} /* (1, 5, 31) {real, imag} */,
  {32'h40050c3c, 32'hc0f31b98} /* (1, 5, 30) {real, imag} */,
  {32'h40753cfe, 32'hc0e6b6a8} /* (1, 5, 29) {real, imag} */,
  {32'h3f0d2537, 32'hc10822e0} /* (1, 5, 28) {real, imag} */,
  {32'hc03f3724, 32'hc12583b5} /* (1, 5, 27) {real, imag} */,
  {32'hbf6404a3, 32'hc0eb24b6} /* (1, 5, 26) {real, imag} */,
  {32'h3f675e98, 32'hc0bd16c9} /* (1, 5, 25) {real, imag} */,
  {32'h3f86e3e8, 32'hc0b8f815} /* (1, 5, 24) {real, imag} */,
  {32'h3f787e7e, 32'hc1093498} /* (1, 5, 23) {real, imag} */,
  {32'h3fe87647, 32'hc1137a34} /* (1, 5, 22) {real, imag} */,
  {32'h40420d02, 32'hc0b71014} /* (1, 5, 21) {real, imag} */,
  {32'h3fe6604e, 32'hc014bc2a} /* (1, 5, 20) {real, imag} */,
  {32'h3f90193f, 32'hc024cf2e} /* (1, 5, 19) {real, imag} */,
  {32'hbdcc6988, 32'hc0136a7a} /* (1, 5, 18) {real, imag} */,
  {32'hc053aee9, 32'hc0384229} /* (1, 5, 17) {real, imag} */,
  {32'hc04c73f4, 32'h3f8c9c87} /* (1, 5, 16) {real, imag} */,
  {32'hc0250978, 32'h41170d00} /* (1, 5, 15) {real, imag} */,
  {32'hc004a2ba, 32'h411e14c1} /* (1, 5, 14) {real, imag} */,
  {32'hc01c9d95, 32'h40b01c80} /* (1, 5, 13) {real, imag} */,
  {32'h4013d11d, 32'h40eca9bc} /* (1, 5, 12) {real, imag} */,
  {32'hbf8f7a9c, 32'h41123310} /* (1, 5, 11) {real, imag} */,
  {32'hbf627a67, 32'h4090ffb9} /* (1, 5, 10) {real, imag} */,
  {32'h3f6a5728, 32'h404e84d5} /* (1, 5, 9) {real, imag} */,
  {32'hbfbd5a0c, 32'h4083561f} /* (1, 5, 8) {real, imag} */,
  {32'hbe100d90, 32'h4056fdc4} /* (1, 5, 7) {real, imag} */,
  {32'hbf9d5b8d, 32'h3ec1473c} /* (1, 5, 6) {real, imag} */,
  {32'h401672b5, 32'hc0e0e1f4} /* (1, 5, 5) {real, imag} */,
  {32'h406ad54c, 32'hc0ed65b0} /* (1, 5, 4) {real, imag} */,
  {32'h403c6bfe, 32'hc1290389} /* (1, 5, 3) {real, imag} */,
  {32'h40130c42, 32'hc1187565} /* (1, 5, 2) {real, imag} */,
  {32'h3faab43e, 32'hc1261c37} /* (1, 5, 1) {real, imag} */,
  {32'h3f686682, 32'hc0a4408e} /* (1, 5, 0) {real, imag} */,
  {32'hbf9885d4, 32'hc0a65d5c} /* (1, 4, 31) {real, imag} */,
  {32'hbfcd4fe0, 32'hc10eb819} /* (1, 4, 30) {real, imag} */,
  {32'hbf47b3ed, 32'hc0e45f0e} /* (1, 4, 29) {real, imag} */,
  {32'hbf9c797b, 32'hc0ca7cf2} /* (1, 4, 28) {real, imag} */,
  {32'hc02efdb1, 32'hc133e12f} /* (1, 4, 27) {real, imag} */,
  {32'hc0258eae, 32'hc10f112c} /* (1, 4, 26) {real, imag} */,
  {32'hc0499fa8, 32'hc101c264} /* (1, 4, 25) {real, imag} */,
  {32'hc0009dda, 32'hc1022be2} /* (1, 4, 24) {real, imag} */,
  {32'hbfab6683, 32'hc1138249} /* (1, 4, 23) {real, imag} */,
  {32'hc00f2a79, 32'hc127090a} /* (1, 4, 22) {real, imag} */,
  {32'h3f06f58a, 32'hc115de73} /* (1, 4, 21) {real, imag} */,
  {32'h40036d71, 32'hc12987a1} /* (1, 4, 20) {real, imag} */,
  {32'h3fd4096a, 32'hc11324ca} /* (1, 4, 19) {real, imag} */,
  {32'h3f8b623c, 32'hc10f64fe} /* (1, 4, 18) {real, imag} */,
  {32'hbe2f509c, 32'hc11c898a} /* (1, 4, 17) {real, imag} */,
  {32'hbfc75118, 32'hc08ee8fe} /* (1, 4, 16) {real, imag} */,
  {32'hbe822c00, 32'h4105f316} /* (1, 4, 15) {real, imag} */,
  {32'hc00dd65e, 32'h40e85edc} /* (1, 4, 14) {real, imag} */,
  {32'hbfa1a482, 32'h4096b1cf} /* (1, 4, 13) {real, imag} */,
  {32'h3e875943, 32'h40ff5804} /* (1, 4, 12) {real, imag} */,
  {32'hc0218d48, 32'h4113684d} /* (1, 4, 11) {real, imag} */,
  {32'hc02bd995, 32'h40c97328} /* (1, 4, 10) {real, imag} */,
  {32'hbf1ff08a, 32'h41049600} /* (1, 4, 9) {real, imag} */,
  {32'hbfd3cb65, 32'h413d2652} /* (1, 4, 8) {real, imag} */,
  {32'hbf24343d, 32'h41170ee6} /* (1, 4, 7) {real, imag} */,
  {32'hbf279aae, 32'h40efb04f} /* (1, 4, 6) {real, imag} */,
  {32'h4071972f, 32'hbf5135b2} /* (1, 4, 5) {real, imag} */,
  {32'h40a1b5ae, 32'hc0cd6fe8} /* (1, 4, 4) {real, imag} */,
  {32'h3fbf7a2e, 32'hc1071afb} /* (1, 4, 3) {real, imag} */,
  {32'hbe0464aa, 32'hc0e5cba6} /* (1, 4, 2) {real, imag} */,
  {32'hbf882409, 32'hc10ecf96} /* (1, 4, 1) {real, imag} */,
  {32'h3e8a3045, 32'hc0a70a44} /* (1, 4, 0) {real, imag} */,
  {32'hbfb7bf67, 32'hc08dbf94} /* (1, 3, 31) {real, imag} */,
  {32'h3fdab86c, 32'hc0f87aea} /* (1, 3, 30) {real, imag} */,
  {32'h3cfa8e10, 32'hc0fa002d} /* (1, 3, 29) {real, imag} */,
  {32'hc00af643, 32'hc0e940a2} /* (1, 3, 28) {real, imag} */,
  {32'hbead4cc9, 32'hc108d6f8} /* (1, 3, 27) {real, imag} */,
  {32'h3eaf6e02, 32'hc0da27de} /* (1, 3, 26) {real, imag} */,
  {32'hbf82af02, 32'hc11694d8} /* (1, 3, 25) {real, imag} */,
  {32'hc03c64ee, 32'hc146cc10} /* (1, 3, 24) {real, imag} */,
  {32'hbf90dd96, 32'hc1253761} /* (1, 3, 23) {real, imag} */,
  {32'h3e92a0dc, 32'hc11f129a} /* (1, 3, 22) {real, imag} */,
  {32'h3fb2bc49, 32'hc11c0a3a} /* (1, 3, 21) {real, imag} */,
  {32'h3fb1d09a, 32'hc10ff323} /* (1, 3, 20) {real, imag} */,
  {32'h3b3b3c00, 32'hc0ebb832} /* (1, 3, 19) {real, imag} */,
  {32'h3f709766, 32'hc0e7f70a} /* (1, 3, 18) {real, imag} */,
  {32'h3ffee701, 32'hc0fb44f4} /* (1, 3, 17) {real, imag} */,
  {32'hbfa030ab, 32'hc06ec0d4} /* (1, 3, 16) {real, imag} */,
  {32'hbf51425e, 32'h40e08a05} /* (1, 3, 15) {real, imag} */,
  {32'hbff78a00, 32'h41086eb8} /* (1, 3, 14) {real, imag} */,
  {32'hbf9c8e1d, 32'h41078a48} /* (1, 3, 13) {real, imag} */,
  {32'hc015e8b0, 32'h411fcdc0} /* (1, 3, 12) {real, imag} */,
  {32'hbf87dfe7, 32'h4128ab93} /* (1, 3, 11) {real, imag} */,
  {32'hbff15dfa, 32'h40d76f1d} /* (1, 3, 10) {real, imag} */,
  {32'hc0159a3f, 32'h410c2102} /* (1, 3, 9) {real, imag} */,
  {32'hc02a3af4, 32'h4142e808} /* (1, 3, 8) {real, imag} */,
  {32'hc02e094e, 32'h416ccb7a} /* (1, 3, 7) {real, imag} */,
  {32'hc01c3205, 32'h412fb5b8} /* (1, 3, 6) {real, imag} */,
  {32'hbff0c5e0, 32'hbff32004} /* (1, 3, 5) {real, imag} */,
  {32'hbf4e47b3, 32'hc1310fda} /* (1, 3, 4) {real, imag} */,
  {32'hbf6ffa00, 32'hc0fe504c} /* (1, 3, 3) {real, imag} */,
  {32'h402a3362, 32'hc0f366ce} /* (1, 3, 2) {real, imag} */,
  {32'h3ff67885, 32'hc11bacd5} /* (1, 3, 1) {real, imag} */,
  {32'hbd85e9c4, 32'hc0c5bf04} /* (1, 3, 0) {real, imag} */,
  {32'hbeb84a55, 32'hc0600214} /* (1, 2, 31) {real, imag} */,
  {32'h401842e7, 32'hc0ded0a8} /* (1, 2, 30) {real, imag} */,
  {32'h3e2833b8, 32'hc10bd75f} /* (1, 2, 29) {real, imag} */,
  {32'hc033876e, 32'hc10f4b8e} /* (1, 2, 28) {real, imag} */,
  {32'h3d1e25a8, 32'hc0f986ca} /* (1, 2, 27) {real, imag} */,
  {32'h3fda5011, 32'hc0cd1912} /* (1, 2, 26) {real, imag} */,
  {32'hbc6422a0, 32'hc115f4b4} /* (1, 2, 25) {real, imag} */,
  {32'h3e63c7f8, 32'hc139c046} /* (1, 2, 24) {real, imag} */,
  {32'h3fc2db00, 32'hc131d8a7} /* (1, 2, 23) {real, imag} */,
  {32'h407cbfe9, 32'hc10b46e6} /* (1, 2, 22) {real, imag} */,
  {32'h401bbd52, 32'hc0d572be} /* (1, 2, 21) {real, imag} */,
  {32'hbf28974a, 32'hc0e75a1f} /* (1, 2, 20) {real, imag} */,
  {32'hbeebe65a, 32'hc121b5a0} /* (1, 2, 19) {real, imag} */,
  {32'h400628c1, 32'hc12c440a} /* (1, 2, 18) {real, imag} */,
  {32'h401c2ceb, 32'hc10aa99a} /* (1, 2, 17) {real, imag} */,
  {32'hbf74836b, 32'hc0ca84da} /* (1, 2, 16) {real, imag} */,
  {32'hbee18916, 32'h3ffeda6b} /* (1, 2, 15) {real, imag} */,
  {32'h3e8e8ae2, 32'h40f60b56} /* (1, 2, 14) {real, imag} */,
  {32'h3f11caa8, 32'h410b4dd7} /* (1, 2, 13) {real, imag} */,
  {32'h3f142b2f, 32'h40f9967f} /* (1, 2, 12) {real, imag} */,
  {32'h3f4f152f, 32'h40e78a94} /* (1, 2, 11) {real, imag} */,
  {32'hbfa3d9ec, 32'h40d4dcca} /* (1, 2, 10) {real, imag} */,
  {32'hbfc9124c, 32'h40e5f85a} /* (1, 2, 9) {real, imag} */,
  {32'hc0012881, 32'h41151f37} /* (1, 2, 8) {real, imag} */,
  {32'hbfcdec8a, 32'h413f1d7c} /* (1, 2, 7) {real, imag} */,
  {32'hbf5d1549, 32'h41257ca0} /* (1, 2, 6) {real, imag} */,
  {32'hc086fb92, 32'hc0328fc8} /* (1, 2, 5) {real, imag} */,
  {32'hc0896375, 32'hc1210cd6} /* (1, 2, 4) {real, imag} */,
  {32'hbf3646a1, 32'hc1043156} /* (1, 2, 3) {real, imag} */,
  {32'h3fe08413, 32'hc131a6db} /* (1, 2, 2) {real, imag} */,
  {32'h3e8a2987, 32'hc1069f5a} /* (1, 2, 1) {real, imag} */,
  {32'hbf7646d3, 32'hc04d5ee4} /* (1, 2, 0) {real, imag} */,
  {32'h3e1f8b68, 32'hbfca4872} /* (1, 1, 31) {real, imag} */,
  {32'h3ed4f557, 32'hc09446f2} /* (1, 1, 30) {real, imag} */,
  {32'h3f4ece2a, 32'hc10f7e00} /* (1, 1, 29) {real, imag} */,
  {32'h3f0b788a, 32'hc1397801} /* (1, 1, 28) {real, imag} */,
  {32'h3ed30fc5, 32'hc131c037} /* (1, 1, 27) {real, imag} */,
  {32'h3f03dd47, 32'hc1046014} /* (1, 1, 26) {real, imag} */,
  {32'h3fb1ad2f, 32'hc0ea3142} /* (1, 1, 25) {real, imag} */,
  {32'h40411f24, 32'hc105c18d} /* (1, 1, 24) {real, imag} */,
  {32'h401bb2b6, 32'hc0ed940c} /* (1, 1, 23) {real, imag} */,
  {32'h405bbbf5, 32'hc0228dba} /* (1, 1, 22) {real, imag} */,
  {32'h3fdf5cb9, 32'hc09e115c} /* (1, 1, 21) {real, imag} */,
  {32'hbe79f0d7, 32'hc0de606b} /* (1, 1, 20) {real, imag} */,
  {32'h3f813268, 32'hc0ff4e5c} /* (1, 1, 19) {real, imag} */,
  {32'h4082c4b4, 32'hc1129040} /* (1, 1, 18) {real, imag} */,
  {32'h40b3154e, 32'hc10a6673} /* (1, 1, 17) {real, imag} */,
  {32'h3eeebcc1, 32'hc0bf84e2} /* (1, 1, 16) {real, imag} */,
  {32'hbf8f69d1, 32'h4009e19e} /* (1, 1, 15) {real, imag} */,
  {32'h3f63b0a4, 32'h40ca0202} /* (1, 1, 14) {real, imag} */,
  {32'h40202784, 32'h40ce2cc9} /* (1, 1, 13) {real, imag} */,
  {32'hbe6d0dac, 32'h40ed7988} /* (1, 1, 12) {real, imag} */,
  {32'hbf773530, 32'h40f08e75} /* (1, 1, 11) {real, imag} */,
  {32'h3f318ef8, 32'h40cbc8fa} /* (1, 1, 10) {real, imag} */,
  {32'h3e84aeb8, 32'h40d61749} /* (1, 1, 9) {real, imag} */,
  {32'h3e488e20, 32'h411b58fc} /* (1, 1, 8) {real, imag} */,
  {32'h4066fd9c, 32'h40fd4aa9} /* (1, 1, 7) {real, imag} */,
  {32'h4059bf28, 32'h40b7ee34} /* (1, 1, 6) {real, imag} */,
  {32'hc0067c51, 32'hbd68abd0} /* (1, 1, 5) {real, imag} */,
  {32'hbf745343, 32'hc086e9ea} /* (1, 1, 4) {real, imag} */,
  {32'h401e0858, 32'hc0e09d4f} /* (1, 1, 3) {real, imag} */,
  {32'h40125fe1, 32'hc0dbf98e} /* (1, 1, 2) {real, imag} */,
  {32'hbf2434da, 32'hc0babb36} /* (1, 1, 1) {real, imag} */,
  {32'hbeeb5f14, 32'hc0041de9} /* (1, 1, 0) {real, imag} */,
  {32'h3f2253fa, 32'hc009cb42} /* (1, 0, 31) {real, imag} */,
  {32'h3e8c7019, 32'hc0524b3d} /* (1, 0, 30) {real, imag} */,
  {32'hbef5413c, 32'hc052dc8f} /* (1, 0, 29) {real, imag} */,
  {32'hbf2f94a6, 32'hc0befcbc} /* (1, 0, 28) {real, imag} */,
  {32'hbecc3bff, 32'hc1241210} /* (1, 0, 27) {real, imag} */,
  {32'h3ead008f, 32'hc107f058} /* (1, 0, 26) {real, imag} */,
  {32'h4008d35f, 32'hc081d6cd} /* (1, 0, 25) {real, imag} */,
  {32'h3f9923f6, 32'hc0698ac6} /* (1, 0, 24) {real, imag} */,
  {32'hbfbd361e, 32'hc0134fc0} /* (1, 0, 23) {real, imag} */,
  {32'h3f9fa477, 32'hbf24c766} /* (1, 0, 22) {real, imag} */,
  {32'h40289836, 32'hc006b68b} /* (1, 0, 21) {real, imag} */,
  {32'h3ffef21d, 32'hc03b2764} /* (1, 0, 20) {real, imag} */,
  {32'h3f4b26fc, 32'hc0164ba4} /* (1, 0, 19) {real, imag} */,
  {32'h3f6712d3, 32'hc03624eb} /* (1, 0, 18) {real, imag} */,
  {32'h4031c478, 32'hc08b793c} /* (1, 0, 17) {real, imag} */,
  {32'hbe439c74, 32'hc00c26c5} /* (1, 0, 16) {real, imag} */,
  {32'hbfa5ff47, 32'h401d95f6} /* (1, 0, 15) {real, imag} */,
  {32'h3f8a8e13, 32'h408ea482} /* (1, 0, 14) {real, imag} */,
  {32'h3fa7cc36, 32'h40474116} /* (1, 0, 13) {real, imag} */,
  {32'hc00eb34c, 32'h408e16da} /* (1, 0, 12) {real, imag} */,
  {32'hc01b622c, 32'h40b30860} /* (1, 0, 11) {real, imag} */,
  {32'h3f1fb5f8, 32'h4080bf6c} /* (1, 0, 10) {real, imag} */,
  {32'h3e9d2039, 32'h40971bca} /* (1, 0, 9) {real, imag} */,
  {32'h3e8ee750, 32'h40c83518} /* (1, 0, 8) {real, imag} */,
  {32'h3fbb5e17, 32'h404e868e} /* (1, 0, 7) {real, imag} */,
  {32'h401e2ce4, 32'h3ec7268f} /* (1, 0, 6) {real, imag} */,
  {32'h3de617a0, 32'hbcd6fd38} /* (1, 0, 5) {real, imag} */,
  {32'hbd3bdd64, 32'hbf9b5364} /* (1, 0, 4) {real, imag} */,
  {32'hbf4821e7, 32'hc08ad53b} /* (1, 0, 3) {real, imag} */,
  {32'hbf1584c2, 32'hc0590231} /* (1, 0, 2) {real, imag} */,
  {32'h3e00f1b0, 32'hc089d1b8} /* (1, 0, 1) {real, imag} */,
  {32'h3e3903ca, 32'hc01235b4} /* (1, 0, 0) {real, imag} */,
  {32'hbfa0b8fc, 32'h00000000} /* (0, 31, 31) {real, imag} */,
  {32'hbfb1c9e2, 32'h00000000} /* (0, 31, 30) {real, imag} */,
  {32'h3eb9ad36, 32'h00000000} /* (0, 31, 29) {real, imag} */,
  {32'hbfa6993c, 32'h00000000} /* (0, 31, 28) {real, imag} */,
  {32'h3e9defe2, 32'h00000000} /* (0, 31, 27) {real, imag} */,
  {32'h3fccc140, 32'h00000000} /* (0, 31, 26) {real, imag} */,
  {32'h40450f1b, 32'h00000000} /* (0, 31, 25) {real, imag} */,
  {32'h3f99a583, 32'h00000000} /* (0, 31, 24) {real, imag} */,
  {32'h3e1c89ec, 32'h00000000} /* (0, 31, 23) {real, imag} */,
  {32'hbd327380, 32'h00000000} /* (0, 31, 22) {real, imag} */,
  {32'hbf862d64, 32'h00000000} /* (0, 31, 21) {real, imag} */,
  {32'hc001bb36, 32'h00000000} /* (0, 31, 20) {real, imag} */,
  {32'h3fdda560, 32'h00000000} /* (0, 31, 19) {real, imag} */,
  {32'h4009d148, 32'h00000000} /* (0, 31, 18) {real, imag} */,
  {32'hbf9fc478, 32'h00000000} /* (0, 31, 17) {real, imag} */,
  {32'hbfd4646a, 32'h00000000} /* (0, 31, 16) {real, imag} */,
  {32'hbf08bb72, 32'h00000000} /* (0, 31, 15) {real, imag} */,
  {32'hbffcfa8a, 32'h00000000} /* (0, 31, 14) {real, imag} */,
  {32'hc0503055, 32'h00000000} /* (0, 31, 13) {real, imag} */,
  {32'hc06e18d0, 32'h00000000} /* (0, 31, 12) {real, imag} */,
  {32'hbfaa6d50, 32'h00000000} /* (0, 31, 11) {real, imag} */,
  {32'h3fe7ee54, 32'h00000000} /* (0, 31, 10) {real, imag} */,
  {32'hbf50c844, 32'h00000000} /* (0, 31, 9) {real, imag} */,
  {32'hc052bc39, 32'h00000000} /* (0, 31, 8) {real, imag} */,
  {32'hbf999db3, 32'h00000000} /* (0, 31, 7) {real, imag} */,
  {32'h3f8c1996, 32'h00000000} /* (0, 31, 6) {real, imag} */,
  {32'hbf399ce9, 32'h00000000} /* (0, 31, 5) {real, imag} */,
  {32'h3f633605, 32'h00000000} /* (0, 31, 4) {real, imag} */,
  {32'hbd0ee930, 32'h00000000} /* (0, 31, 3) {real, imag} */,
  {32'h3fbd591c, 32'h00000000} /* (0, 31, 2) {real, imag} */,
  {32'h3f7cc984, 32'h00000000} /* (0, 31, 1) {real, imag} */,
  {32'h3fe6157f, 32'h00000000} /* (0, 31, 0) {real, imag} */,
  {32'h3f88fa6b, 32'h00000000} /* (0, 30, 31) {real, imag} */,
  {32'h3eebaa62, 32'h00000000} /* (0, 30, 30) {real, imag} */,
  {32'hc01524ce, 32'h00000000} /* (0, 30, 29) {real, imag} */,
  {32'hbffac39a, 32'h00000000} /* (0, 30, 28) {real, imag} */,
  {32'h3f9dc155, 32'h00000000} /* (0, 30, 27) {real, imag} */,
  {32'h3fa9bf44, 32'h00000000} /* (0, 30, 26) {real, imag} */,
  {32'h409ca36a, 32'h00000000} /* (0, 30, 25) {real, imag} */,
  {32'h40505b87, 32'h00000000} /* (0, 30, 24) {real, imag} */,
  {32'h407d19b6, 32'h00000000} /* (0, 30, 23) {real, imag} */,
  {32'h3f967040, 32'h00000000} /* (0, 30, 22) {real, imag} */,
  {32'h3e19f7e8, 32'h00000000} /* (0, 30, 21) {real, imag} */,
  {32'h4028081a, 32'h00000000} /* (0, 30, 20) {real, imag} */,
  {32'h3fe20b4c, 32'h00000000} /* (0, 30, 19) {real, imag} */,
  {32'hbfb09652, 32'h00000000} /* (0, 30, 18) {real, imag} */,
  {32'hbfe194df, 32'h00000000} /* (0, 30, 17) {real, imag} */,
  {32'h3f9108a4, 32'h00000000} /* (0, 30, 16) {real, imag} */,
  {32'h3eabda1a, 32'h00000000} /* (0, 30, 15) {real, imag} */,
  {32'hc058ac2f, 32'h00000000} /* (0, 30, 14) {real, imag} */,
  {32'hc0828308, 32'h00000000} /* (0, 30, 13) {real, imag} */,
  {32'hc06db30e, 32'h00000000} /* (0, 30, 12) {real, imag} */,
  {32'h3f6f52bd, 32'h00000000} /* (0, 30, 11) {real, imag} */,
  {32'h4053d51a, 32'h00000000} /* (0, 30, 10) {real, imag} */,
  {32'hbe1cc884, 32'h00000000} /* (0, 30, 9) {real, imag} */,
  {32'hc01447bc, 32'h00000000} /* (0, 30, 8) {real, imag} */,
  {32'hbfe910e3, 32'h00000000} /* (0, 30, 7) {real, imag} */,
  {32'hbf8d6f5b, 32'h00000000} /* (0, 30, 6) {real, imag} */,
  {32'h4007b1f6, 32'h00000000} /* (0, 30, 5) {real, imag} */,
  {32'h40439540, 32'h00000000} /* (0, 30, 4) {real, imag} */,
  {32'h3fa83954, 32'h00000000} /* (0, 30, 3) {real, imag} */,
  {32'h3f811e13, 32'h00000000} /* (0, 30, 2) {real, imag} */,
  {32'h40a0d8c9, 32'h00000000} /* (0, 30, 1) {real, imag} */,
  {32'h408a6636, 32'h00000000} /* (0, 30, 0) {real, imag} */,
  {32'h40292f9e, 32'h00000000} /* (0, 29, 31) {real, imag} */,
  {32'h3fbb1904, 32'h00000000} /* (0, 29, 30) {real, imag} */,
  {32'hc08b0838, 32'h00000000} /* (0, 29, 29) {real, imag} */,
  {32'hbf97750d, 32'h00000000} /* (0, 29, 28) {real, imag} */,
  {32'hbf76bc26, 32'h00000000} /* (0, 29, 27) {real, imag} */,
  {32'hc035956e, 32'h00000000} /* (0, 29, 26) {real, imag} */,
  {32'hc086bd14, 32'h00000000} /* (0, 29, 25) {real, imag} */,
  {32'hc03e5f89, 32'h00000000} /* (0, 29, 24) {real, imag} */,
  {32'hbd0f7350, 32'h00000000} /* (0, 29, 23) {real, imag} */,
  {32'hbeb4b226, 32'h00000000} /* (0, 29, 22) {real, imag} */,
  {32'h3f92c6e6, 32'h00000000} /* (0, 29, 21) {real, imag} */,
  {32'h3fd59868, 32'h00000000} /* (0, 29, 20) {real, imag} */,
  {32'h403568e0, 32'h00000000} /* (0, 29, 19) {real, imag} */,
  {32'h3f089509, 32'h00000000} /* (0, 29, 18) {real, imag} */,
  {32'h4084c12e, 32'h00000000} /* (0, 29, 17) {real, imag} */,
  {32'h40355c08, 32'h00000000} /* (0, 29, 16) {real, imag} */,
  {32'hbf8f997e, 32'h00000000} /* (0, 29, 15) {real, imag} */,
  {32'hc06551df, 32'h00000000} /* (0, 29, 14) {real, imag} */,
  {32'hbff905fa, 32'h00000000} /* (0, 29, 13) {real, imag} */,
  {32'h40312acd, 32'h00000000} /* (0, 29, 12) {real, imag} */,
  {32'h3fd0af7d, 32'h00000000} /* (0, 29, 11) {real, imag} */,
  {32'h3fb4c433, 32'h00000000} /* (0, 29, 10) {real, imag} */,
  {32'h3cd59c00, 32'h00000000} /* (0, 29, 9) {real, imag} */,
  {32'hbff79884, 32'h00000000} /* (0, 29, 8) {real, imag} */,
  {32'hc0608f43, 32'h00000000} /* (0, 29, 7) {real, imag} */,
  {32'h3e990ba8, 32'h00000000} /* (0, 29, 6) {real, imag} */,
  {32'h40b9426a, 32'h00000000} /* (0, 29, 5) {real, imag} */,
  {32'h408fa95f, 32'h00000000} /* (0, 29, 4) {real, imag} */,
  {32'h402e089c, 32'h00000000} /* (0, 29, 3) {real, imag} */,
  {32'hbf115ed8, 32'h00000000} /* (0, 29, 2) {real, imag} */,
  {32'h3f82878e, 32'h00000000} /* (0, 29, 1) {real, imag} */,
  {32'h3ef01c3c, 32'h00000000} /* (0, 29, 0) {real, imag} */,
  {32'h3f1773ca, 32'h00000000} /* (0, 28, 31) {real, imag} */,
  {32'h3f52ca18, 32'h00000000} /* (0, 28, 30) {real, imag} */,
  {32'hc0193aa6, 32'h00000000} /* (0, 28, 29) {real, imag} */,
  {32'hbff1cdb8, 32'h00000000} /* (0, 28, 28) {real, imag} */,
  {32'hbfcb90e9, 32'h00000000} /* (0, 28, 27) {real, imag} */,
  {32'hbfaf300f, 32'h00000000} /* (0, 28, 26) {real, imag} */,
  {32'hc0e90d1c, 32'h00000000} /* (0, 28, 25) {real, imag} */,
  {32'hc09f15fd, 32'h00000000} /* (0, 28, 24) {real, imag} */,
  {32'hc0198224, 32'h00000000} /* (0, 28, 23) {real, imag} */,
  {32'hbfdea987, 32'h00000000} /* (0, 28, 22) {real, imag} */,
  {32'h3fcf10cc, 32'h00000000} /* (0, 28, 21) {real, imag} */,
  {32'hbf910d6b, 32'h00000000} /* (0, 28, 20) {real, imag} */,
  {32'h3e4b58e8, 32'h00000000} /* (0, 28, 19) {real, imag} */,
  {32'h40321586, 32'h00000000} /* (0, 28, 18) {real, imag} */,
  {32'h40708754, 32'h00000000} /* (0, 28, 17) {real, imag} */,
  {32'h405197c2, 32'h00000000} /* (0, 28, 16) {real, imag} */,
  {32'h3e899ba1, 32'h00000000} /* (0, 28, 15) {real, imag} */,
  {32'hbff737fc, 32'h00000000} /* (0, 28, 14) {real, imag} */,
  {32'hbf9efa9c, 32'h00000000} /* (0, 28, 13) {real, imag} */,
  {32'h40c77482, 32'h00000000} /* (0, 28, 12) {real, imag} */,
  {32'h40a96afe, 32'h00000000} /* (0, 28, 11) {real, imag} */,
  {32'h4073f85d, 32'h00000000} /* (0, 28, 10) {real, imag} */,
  {32'h3ecbd9e8, 32'h00000000} /* (0, 28, 9) {real, imag} */,
  {32'hbf137be8, 32'h00000000} /* (0, 28, 8) {real, imag} */,
  {32'hc0259214, 32'h00000000} /* (0, 28, 7) {real, imag} */,
  {32'h3f809279, 32'h00000000} /* (0, 28, 6) {real, imag} */,
  {32'h4032778f, 32'h00000000} /* (0, 28, 5) {real, imag} */,
  {32'h3f202bf1, 32'h00000000} /* (0, 28, 4) {real, imag} */,
  {32'hc01b0812, 32'h00000000} /* (0, 28, 3) {real, imag} */,
  {32'hc01614d1, 32'h00000000} /* (0, 28, 2) {real, imag} */,
  {32'hc059a57e, 32'h00000000} /* (0, 28, 1) {real, imag} */,
  {32'hbfb5bbe2, 32'h00000000} /* (0, 28, 0) {real, imag} */,
  {32'h40117a0c, 32'h00000000} /* (0, 27, 31) {real, imag} */,
  {32'h3f94603b, 32'h00000000} /* (0, 27, 30) {real, imag} */,
  {32'h402096c2, 32'h00000000} /* (0, 27, 29) {real, imag} */,
  {32'h3f8f4273, 32'h00000000} /* (0, 27, 28) {real, imag} */,
  {32'h3f1bbbc1, 32'h00000000} /* (0, 27, 27) {real, imag} */,
  {32'h3fdfe6cd, 32'h00000000} /* (0, 27, 26) {real, imag} */,
  {32'hbfe92c8c, 32'h00000000} /* (0, 27, 25) {real, imag} */,
  {32'hc07f63d8, 32'h00000000} /* (0, 27, 24) {real, imag} */,
  {32'hbfb9f404, 32'h00000000} /* (0, 27, 23) {real, imag} */,
  {32'h405b0776, 32'h00000000} /* (0, 27, 22) {real, imag} */,
  {32'h40a7add8, 32'h00000000} /* (0, 27, 21) {real, imag} */,
  {32'h3c540280, 32'h00000000} /* (0, 27, 20) {real, imag} */,
  {32'hbeba8d3e, 32'h00000000} /* (0, 27, 19) {real, imag} */,
  {32'hbf2835a2, 32'h00000000} /* (0, 27, 18) {real, imag} */,
  {32'hbf1e8d69, 32'h00000000} /* (0, 27, 17) {real, imag} */,
  {32'hc0664e0d, 32'h00000000} /* (0, 27, 16) {real, imag} */,
  {32'hbff5af53, 32'h00000000} /* (0, 27, 15) {real, imag} */,
  {32'hbe8fb9d0, 32'h00000000} /* (0, 27, 14) {real, imag} */,
  {32'h40143ab2, 32'h00000000} /* (0, 27, 13) {real, imag} */,
  {32'h40902e72, 32'h00000000} /* (0, 27, 12) {real, imag} */,
  {32'h402f4200, 32'h00000000} /* (0, 27, 11) {real, imag} */,
  {32'h3f0c7488, 32'h00000000} /* (0, 27, 10) {real, imag} */,
  {32'hbf33ceba, 32'h00000000} /* (0, 27, 9) {real, imag} */,
  {32'h40060c1a, 32'h00000000} /* (0, 27, 8) {real, imag} */,
  {32'h40754716, 32'h00000000} /* (0, 27, 7) {real, imag} */,
  {32'h3fa1ae62, 32'h00000000} /* (0, 27, 6) {real, imag} */,
  {32'hbfa0b70b, 32'h00000000} /* (0, 27, 5) {real, imag} */,
  {32'hc020a6c4, 32'h00000000} /* (0, 27, 4) {real, imag} */,
  {32'hc0610c7e, 32'h00000000} /* (0, 27, 3) {real, imag} */,
  {32'hc0a0fbec, 32'h00000000} /* (0, 27, 2) {real, imag} */,
  {32'hc035f805, 32'h00000000} /* (0, 27, 1) {real, imag} */,
  {32'h3fab4ed0, 32'h00000000} /* (0, 27, 0) {real, imag} */,
  {32'h3fa9f44e, 32'h00000000} /* (0, 26, 31) {real, imag} */,
  {32'hbfdea655, 32'h00000000} /* (0, 26, 30) {real, imag} */,
  {32'h40007d76, 32'h00000000} /* (0, 26, 29) {real, imag} */,
  {32'h3f4b05e9, 32'h00000000} /* (0, 26, 28) {real, imag} */,
  {32'h3e25a348, 32'h00000000} /* (0, 26, 27) {real, imag} */,
  {32'h3f86b7e6, 32'h00000000} /* (0, 26, 26) {real, imag} */,
  {32'h3fecf0a8, 32'h00000000} /* (0, 26, 25) {real, imag} */,
  {32'hc03fe187, 32'h00000000} /* (0, 26, 24) {real, imag} */,
  {32'hc09971fa, 32'h00000000} /* (0, 26, 23) {real, imag} */,
  {32'h3df1a9b0, 32'h00000000} /* (0, 26, 22) {real, imag} */,
  {32'h3f2ca4c8, 32'h00000000} /* (0, 26, 21) {real, imag} */,
  {32'hbff6d1b0, 32'h00000000} /* (0, 26, 20) {real, imag} */,
  {32'hbfa5b27a, 32'h00000000} /* (0, 26, 19) {real, imag} */,
  {32'hc049ba02, 32'h00000000} /* (0, 26, 18) {real, imag} */,
  {32'hc046fa80, 32'h00000000} /* (0, 26, 17) {real, imag} */,
  {32'hc0e9d6c9, 32'h00000000} /* (0, 26, 16) {real, imag} */,
  {32'hc0515981, 32'h00000000} /* (0, 26, 15) {real, imag} */,
  {32'h3f6b86ca, 32'h00000000} /* (0, 26, 14) {real, imag} */,
  {32'h3d880438, 32'h00000000} /* (0, 26, 13) {real, imag} */,
  {32'h402b5d9e, 32'h00000000} /* (0, 26, 12) {real, imag} */,
  {32'h3e8586e4, 32'h00000000} /* (0, 26, 11) {real, imag} */,
  {32'hc0543d27, 32'h00000000} /* (0, 26, 10) {real, imag} */,
  {32'hbf4d7c92, 32'h00000000} /* (0, 26, 9) {real, imag} */,
  {32'h402dd483, 32'h00000000} /* (0, 26, 8) {real, imag} */,
  {32'h40756105, 32'h00000000} /* (0, 26, 7) {real, imag} */,
  {32'h3f0114b7, 32'h00000000} /* (0, 26, 6) {real, imag} */,
  {32'h3f8811e7, 32'h00000000} /* (0, 26, 5) {real, imag} */,
  {32'h3eed2b8c, 32'h00000000} /* (0, 26, 4) {real, imag} */,
  {32'h3f2714b2, 32'h00000000} /* (0, 26, 3) {real, imag} */,
  {32'hc0247a1a, 32'h00000000} /* (0, 26, 2) {real, imag} */,
  {32'hc027da26, 32'h00000000} /* (0, 26, 1) {real, imag} */,
  {32'h3ef65b4c, 32'h00000000} /* (0, 26, 0) {real, imag} */,
  {32'h3e1e5de6, 32'h00000000} /* (0, 25, 31) {real, imag} */,
  {32'hc075ca46, 32'h00000000} /* (0, 25, 30) {real, imag} */,
  {32'hc018c318, 32'h00000000} /* (0, 25, 29) {real, imag} */,
  {32'h3e32b3c0, 32'h00000000} /* (0, 25, 28) {real, imag} */,
  {32'hc025ef8a, 32'h00000000} /* (0, 25, 27) {real, imag} */,
  {32'hc03740aa, 32'h00000000} /* (0, 25, 26) {real, imag} */,
  {32'h402e0e70, 32'h00000000} /* (0, 25, 25) {real, imag} */,
  {32'h3ecdb186, 32'h00000000} /* (0, 25, 24) {real, imag} */,
  {32'hc06e44f4, 32'h00000000} /* (0, 25, 23) {real, imag} */,
  {32'hc018ddcb, 32'h00000000} /* (0, 25, 22) {real, imag} */,
  {32'h3ed33858, 32'h00000000} /* (0, 25, 21) {real, imag} */,
  {32'h40c758fa, 32'h00000000} /* (0, 25, 20) {real, imag} */,
  {32'h40af9d9e, 32'h00000000} /* (0, 25, 19) {real, imag} */,
  {32'hbeeaf702, 32'h00000000} /* (0, 25, 18) {real, imag} */,
  {32'hc0abbfc6, 32'h00000000} /* (0, 25, 17) {real, imag} */,
  {32'hc08d4686, 32'h00000000} /* (0, 25, 16) {real, imag} */,
  {32'hbef0b508, 32'h00000000} /* (0, 25, 15) {real, imag} */,
  {32'h3e454320, 32'h00000000} /* (0, 25, 14) {real, imag} */,
  {32'hbfb762a0, 32'h00000000} /* (0, 25, 13) {real, imag} */,
  {32'hbe67fc80, 32'h00000000} /* (0, 25, 12) {real, imag} */,
  {32'h3f1e3a66, 32'h00000000} /* (0, 25, 11) {real, imag} */,
  {32'hc03a8d74, 32'h00000000} /* (0, 25, 10) {real, imag} */,
  {32'hc01a395d, 32'h00000000} /* (0, 25, 9) {real, imag} */,
  {32'hbf893950, 32'h00000000} /* (0, 25, 8) {real, imag} */,
  {32'h3ee95b1e, 32'h00000000} /* (0, 25, 7) {real, imag} */,
  {32'h3f2097e8, 32'h00000000} /* (0, 25, 6) {real, imag} */,
  {32'h40c47f6c, 32'h00000000} /* (0, 25, 5) {real, imag} */,
  {32'h403a8d8c, 32'h00000000} /* (0, 25, 4) {real, imag} */,
  {32'hbfd88784, 32'h00000000} /* (0, 25, 3) {real, imag} */,
  {32'hc09f10cc, 32'h00000000} /* (0, 25, 2) {real, imag} */,
  {32'hc08b1622, 32'h00000000} /* (0, 25, 1) {real, imag} */,
  {32'hc009fec9, 32'h00000000} /* (0, 25, 0) {real, imag} */,
  {32'h3f5f57b6, 32'h00000000} /* (0, 24, 31) {real, imag} */,
  {32'h4023bfe4, 32'h00000000} /* (0, 24, 30) {real, imag} */,
  {32'h40177a89, 32'h00000000} /* (0, 24, 29) {real, imag} */,
  {32'h4011f9e7, 32'h00000000} /* (0, 24, 28) {real, imag} */,
  {32'h3f7c4aca, 32'h00000000} /* (0, 24, 27) {real, imag} */,
  {32'h3ea43166, 32'h00000000} /* (0, 24, 26) {real, imag} */,
  {32'h4018074f, 32'h00000000} /* (0, 24, 25) {real, imag} */,
  {32'h4014f738, 32'h00000000} /* (0, 24, 24) {real, imag} */,
  {32'hc02295dc, 32'h00000000} /* (0, 24, 23) {real, imag} */,
  {32'hc0208aa6, 32'h00000000} /* (0, 24, 22) {real, imag} */,
  {32'h3f9c335e, 32'h00000000} /* (0, 24, 21) {real, imag} */,
  {32'h40920725, 32'h00000000} /* (0, 24, 20) {real, imag} */,
  {32'h407234b6, 32'h00000000} /* (0, 24, 19) {real, imag} */,
  {32'h4051f3b6, 32'h00000000} /* (0, 24, 18) {real, imag} */,
  {32'hbf5f4cd4, 32'h00000000} /* (0, 24, 17) {real, imag} */,
  {32'hc0364cc0, 32'h00000000} /* (0, 24, 16) {real, imag} */,
  {32'hbfd22728, 32'h00000000} /* (0, 24, 15) {real, imag} */,
  {32'hbe80f498, 32'h00000000} /* (0, 24, 14) {real, imag} */,
  {32'hc046750a, 32'h00000000} /* (0, 24, 13) {real, imag} */,
  {32'hc09002f3, 32'h00000000} /* (0, 24, 12) {real, imag} */,
  {32'hc0817c5c, 32'h00000000} /* (0, 24, 11) {real, imag} */,
  {32'hc084adf2, 32'h00000000} /* (0, 24, 10) {real, imag} */,
  {32'h3fc1ca9e, 32'h00000000} /* (0, 24, 9) {real, imag} */,
  {32'h4007a6a0, 32'h00000000} /* (0, 24, 8) {real, imag} */,
  {32'h404f3804, 32'h00000000} /* (0, 24, 7) {real, imag} */,
  {32'h4013e28e, 32'h00000000} /* (0, 24, 6) {real, imag} */,
  {32'h4056dad0, 32'h00000000} /* (0, 24, 5) {real, imag} */,
  {32'h403fbe9e, 32'h00000000} /* (0, 24, 4) {real, imag} */,
  {32'hbd7de3a0, 32'h00000000} /* (0, 24, 3) {real, imag} */,
  {32'hc04ecabf, 32'h00000000} /* (0, 24, 2) {real, imag} */,
  {32'hc06cf546, 32'h00000000} /* (0, 24, 1) {real, imag} */,
  {32'hbfecb296, 32'h00000000} /* (0, 24, 0) {real, imag} */,
  {32'h3f371838, 32'h00000000} /* (0, 23, 31) {real, imag} */,
  {32'h40c125cc, 32'h00000000} /* (0, 23, 30) {real, imag} */,
  {32'h3ff0cb50, 32'h00000000} /* (0, 23, 29) {real, imag} */,
  {32'hbfe473fc, 32'h00000000} /* (0, 23, 28) {real, imag} */,
  {32'hbf547854, 32'h00000000} /* (0, 23, 27) {real, imag} */,
  {32'h3f7f24dc, 32'h00000000} /* (0, 23, 26) {real, imag} */,
  {32'hbff11e25, 32'h00000000} /* (0, 23, 25) {real, imag} */,
  {32'hbf9f1c02, 32'h00000000} /* (0, 23, 24) {real, imag} */,
  {32'hbfb378df, 32'h00000000} /* (0, 23, 23) {real, imag} */,
  {32'hc005fb6a, 32'h00000000} /* (0, 23, 22) {real, imag} */,
  {32'h40063068, 32'h00000000} /* (0, 23, 21) {real, imag} */,
  {32'h40816857, 32'h00000000} /* (0, 23, 20) {real, imag} */,
  {32'h3eebb024, 32'h00000000} /* (0, 23, 19) {real, imag} */,
  {32'h3df1c6f8, 32'h00000000} /* (0, 23, 18) {real, imag} */,
  {32'h3fd588e2, 32'h00000000} /* (0, 23, 17) {real, imag} */,
  {32'hbea3a72c, 32'h00000000} /* (0, 23, 16) {real, imag} */,
  {32'h40262a86, 32'h00000000} /* (0, 23, 15) {real, imag} */,
  {32'h3f595db6, 32'h00000000} /* (0, 23, 14) {real, imag} */,
  {32'hbf9f7356, 32'h00000000} /* (0, 23, 13) {real, imag} */,
  {32'hbfb55032, 32'h00000000} /* (0, 23, 12) {real, imag} */,
  {32'hc04992de, 32'h00000000} /* (0, 23, 11) {real, imag} */,
  {32'hc09ebd78, 32'h00000000} /* (0, 23, 10) {real, imag} */,
  {32'h40009959, 32'h00000000} /* (0, 23, 9) {real, imag} */,
  {32'h405daa56, 32'h00000000} /* (0, 23, 8) {real, imag} */,
  {32'h405eef36, 32'h00000000} /* (0, 23, 7) {real, imag} */,
  {32'h3fd2724e, 32'h00000000} /* (0, 23, 6) {real, imag} */,
  {32'hc014b1ba, 32'h00000000} /* (0, 23, 5) {real, imag} */,
  {32'hbf1d0cf8, 32'h00000000} /* (0, 23, 4) {real, imag} */,
  {32'hbdf85cf8, 32'h00000000} /* (0, 23, 3) {real, imag} */,
  {32'hc00dde50, 32'h00000000} /* (0, 23, 2) {real, imag} */,
  {32'hc0b4fcda, 32'h00000000} /* (0, 23, 1) {real, imag} */,
  {32'hbfec8983, 32'h00000000} /* (0, 23, 0) {real, imag} */,
  {32'hbf8d67c4, 32'h00000000} /* (0, 22, 31) {real, imag} */,
  {32'h4036ec74, 32'h00000000} /* (0, 22, 30) {real, imag} */,
  {32'h3fb218ac, 32'h00000000} /* (0, 22, 29) {real, imag} */,
  {32'hc0692e4e, 32'h00000000} /* (0, 22, 28) {real, imag} */,
  {32'hc0898323, 32'h00000000} /* (0, 22, 27) {real, imag} */,
  {32'h3e48a960, 32'h00000000} /* (0, 22, 26) {real, imag} */,
  {32'h3e0abef4, 32'h00000000} /* (0, 22, 25) {real, imag} */,
  {32'hbfe49958, 32'h00000000} /* (0, 22, 24) {real, imag} */,
  {32'h40551ae4, 32'h00000000} /* (0, 22, 23) {real, imag} */,
  {32'h404f5ad6, 32'h00000000} /* (0, 22, 22) {real, imag} */,
  {32'hbf521df1, 32'h00000000} /* (0, 22, 21) {real, imag} */,
  {32'h3f2fdce6, 32'h00000000} /* (0, 22, 20) {real, imag} */,
  {32'h403e74be, 32'h00000000} /* (0, 22, 19) {real, imag} */,
  {32'h40390abe, 32'h00000000} /* (0, 22, 18) {real, imag} */,
  {32'h3f41d585, 32'h00000000} /* (0, 22, 17) {real, imag} */,
  {32'hbe61a43c, 32'h00000000} /* (0, 22, 16) {real, imag} */,
  {32'h3fec45da, 32'h00000000} /* (0, 22, 15) {real, imag} */,
  {32'h400182aa, 32'h00000000} /* (0, 22, 14) {real, imag} */,
  {32'h4089a0c4, 32'h00000000} /* (0, 22, 13) {real, imag} */,
  {32'h3fa28d99, 32'h00000000} /* (0, 22, 12) {real, imag} */,
  {32'hbfc35e81, 32'h00000000} /* (0, 22, 11) {real, imag} */,
  {32'hc0023386, 32'h00000000} /* (0, 22, 10) {real, imag} */,
  {32'hbffeb9e8, 32'h00000000} /* (0, 22, 9) {real, imag} */,
  {32'h3ef82a0c, 32'h00000000} /* (0, 22, 8) {real, imag} */,
  {32'h3f81a701, 32'h00000000} /* (0, 22, 7) {real, imag} */,
  {32'h3eb2a5a8, 32'h00000000} /* (0, 22, 6) {real, imag} */,
  {32'h3ed8ae30, 32'h00000000} /* (0, 22, 5) {real, imag} */,
  {32'h3f0339fd, 32'h00000000} /* (0, 22, 4) {real, imag} */,
  {32'h3f9e3e71, 32'h00000000} /* (0, 22, 3) {real, imag} */,
  {32'h408d8253, 32'h00000000} /* (0, 22, 2) {real, imag} */,
  {32'hc015db06, 32'h00000000} /* (0, 22, 1) {real, imag} */,
  {32'hc02b67be, 32'h00000000} /* (0, 22, 0) {real, imag} */,
  {32'hbff056e2, 32'h00000000} /* (0, 21, 31) {real, imag} */,
  {32'hbeafb1f5, 32'h00000000} /* (0, 21, 30) {real, imag} */,
  {32'hbf8bfbe8, 32'h00000000} /* (0, 21, 29) {real, imag} */,
  {32'hc00e3b77, 32'h00000000} /* (0, 21, 28) {real, imag} */,
  {32'hc0239ff4, 32'h00000000} /* (0, 21, 27) {real, imag} */,
  {32'hc0595ea9, 32'h00000000} /* (0, 21, 26) {real, imag} */,
  {32'hbfc02318, 32'h00000000} /* (0, 21, 25) {real, imag} */,
  {32'h3e759e58, 32'h00000000} /* (0, 21, 24) {real, imag} */,
  {32'h3ede1c6a, 32'h00000000} /* (0, 21, 23) {real, imag} */,
  {32'h3f953cdd, 32'h00000000} /* (0, 21, 22) {real, imag} */,
  {32'hbf103ac8, 32'h00000000} /* (0, 21, 21) {real, imag} */,
  {32'hc086a880, 32'h00000000} /* (0, 21, 20) {real, imag} */,
  {32'h3f5e9b37, 32'h00000000} /* (0, 21, 19) {real, imag} */,
  {32'h407ccf11, 32'h00000000} /* (0, 21, 18) {real, imag} */,
  {32'hbf1b439d, 32'h00000000} /* (0, 21, 17) {real, imag} */,
  {32'hbf68d887, 32'h00000000} /* (0, 21, 16) {real, imag} */,
  {32'h3f584d30, 32'h00000000} /* (0, 21, 15) {real, imag} */,
  {32'h403a5671, 32'h00000000} /* (0, 21, 14) {real, imag} */,
  {32'h40b5c9e6, 32'h00000000} /* (0, 21, 13) {real, imag} */,
  {32'h408326ac, 32'h00000000} /* (0, 21, 12) {real, imag} */,
  {32'h3ff97b48, 32'h00000000} /* (0, 21, 11) {real, imag} */,
  {32'h3f1e0afe, 32'h00000000} /* (0, 21, 10) {real, imag} */,
  {32'h3ff41e20, 32'h00000000} /* (0, 21, 9) {real, imag} */,
  {32'hbef1bed6, 32'h00000000} /* (0, 21, 8) {real, imag} */,
  {32'hbfc95313, 32'h00000000} /* (0, 21, 7) {real, imag} */,
  {32'h3f2cdae4, 32'h00000000} /* (0, 21, 6) {real, imag} */,
  {32'h3f762be7, 32'h00000000} /* (0, 21, 5) {real, imag} */,
  {32'h3f6f5228, 32'h00000000} /* (0, 21, 4) {real, imag} */,
  {32'h3fe9e048, 32'h00000000} /* (0, 21, 3) {real, imag} */,
  {32'h407fb257, 32'h00000000} /* (0, 21, 2) {real, imag} */,
  {32'hbf66ffbe, 32'h00000000} /* (0, 21, 1) {real, imag} */,
  {32'hbfbd34c6, 32'h00000000} /* (0, 21, 0) {real, imag} */,
  {32'h406baa8a, 32'h00000000} /* (0, 20, 31) {real, imag} */,
  {32'h40a145f2, 32'h00000000} /* (0, 20, 30) {real, imag} */,
  {32'h3e45f6b4, 32'h00000000} /* (0, 20, 29) {real, imag} */,
  {32'h3fb38cee, 32'h00000000} /* (0, 20, 28) {real, imag} */,
  {32'h405dfbf5, 32'h00000000} /* (0, 20, 27) {real, imag} */,
  {32'h3ed9bb4a, 32'h00000000} /* (0, 20, 26) {real, imag} */,
  {32'h3f0d7408, 32'h00000000} /* (0, 20, 25) {real, imag} */,
  {32'h3ffda643, 32'h00000000} /* (0, 20, 24) {real, imag} */,
  {32'h4012bc3c, 32'h00000000} /* (0, 20, 23) {real, imag} */,
  {32'hbf161ce4, 32'h00000000} /* (0, 20, 22) {real, imag} */,
  {32'h3f948b8c, 32'h00000000} /* (0, 20, 21) {real, imag} */,
  {32'hc04a90ed, 32'h00000000} /* (0, 20, 20) {real, imag} */,
  {32'hbf8d4c65, 32'h00000000} /* (0, 20, 19) {real, imag} */,
  {32'h4051406a, 32'h00000000} /* (0, 20, 18) {real, imag} */,
  {32'hbfc536d2, 32'h00000000} /* (0, 20, 17) {real, imag} */,
  {32'hbe962f90, 32'h00000000} /* (0, 20, 16) {real, imag} */,
  {32'h40322324, 32'h00000000} /* (0, 20, 15) {real, imag} */,
  {32'h40519e15, 32'h00000000} /* (0, 20, 14) {real, imag} */,
  {32'h3ff1664c, 32'h00000000} /* (0, 20, 13) {real, imag} */,
  {32'h3faaec7e, 32'h00000000} /* (0, 20, 12) {real, imag} */,
  {32'hbf54d5a0, 32'h00000000} /* (0, 20, 11) {real, imag} */,
  {32'hc01815d4, 32'h00000000} /* (0, 20, 10) {real, imag} */,
  {32'h4019745d, 32'h00000000} /* (0, 20, 9) {real, imag} */,
  {32'hc04ea5ea, 32'h00000000} /* (0, 20, 8) {real, imag} */,
  {32'hc095639c, 32'h00000000} /* (0, 20, 7) {real, imag} */,
  {32'hbd6c63b0, 32'h00000000} /* (0, 20, 6) {real, imag} */,
  {32'hbeb76580, 32'h00000000} /* (0, 20, 5) {real, imag} */,
  {32'hbfdc5e4c, 32'h00000000} /* (0, 20, 4) {real, imag} */,
  {32'hc01a3596, 32'h00000000} /* (0, 20, 3) {real, imag} */,
  {32'hbfe0c9dd, 32'h00000000} /* (0, 20, 2) {real, imag} */,
  {32'hc08cfe9e, 32'h00000000} /* (0, 20, 1) {real, imag} */,
  {32'hc0024106, 32'h00000000} /* (0, 20, 0) {real, imag} */,
  {32'h401845e4, 32'h00000000} /* (0, 19, 31) {real, imag} */,
  {32'h40234e1a, 32'h00000000} /* (0, 19, 30) {real, imag} */,
  {32'hbeb83b04, 32'h00000000} /* (0, 19, 29) {real, imag} */,
  {32'h402bde40, 32'h00000000} /* (0, 19, 28) {real, imag} */,
  {32'h3fceb682, 32'h00000000} /* (0, 19, 27) {real, imag} */,
  {32'hbfd4c9c4, 32'h00000000} /* (0, 19, 26) {real, imag} */,
  {32'h3f5f2b7c, 32'h00000000} /* (0, 19, 25) {real, imag} */,
  {32'h4059e3a6, 32'h00000000} /* (0, 19, 24) {real, imag} */,
  {32'h401c65f7, 32'h00000000} /* (0, 19, 23) {real, imag} */,
  {32'h3ed73764, 32'h00000000} /* (0, 19, 22) {real, imag} */,
  {32'h3f83aeec, 32'h00000000} /* (0, 19, 21) {real, imag} */,
  {32'hbf7c57bc, 32'h00000000} /* (0, 19, 20) {real, imag} */,
  {32'h3f289661, 32'h00000000} /* (0, 19, 19) {real, imag} */,
  {32'hbf3801a4, 32'h00000000} /* (0, 19, 18) {real, imag} */,
  {32'hc00d74ac, 32'h00000000} /* (0, 19, 17) {real, imag} */,
  {32'h4037a9a6, 32'h00000000} /* (0, 19, 16) {real, imag} */,
  {32'h40b34aeb, 32'h00000000} /* (0, 19, 15) {real, imag} */,
  {32'h40a24d2c, 32'h00000000} /* (0, 19, 14) {real, imag} */,
  {32'h404a2cb4, 32'h00000000} /* (0, 19, 13) {real, imag} */,
  {32'hbf63bfaa, 32'h00000000} /* (0, 19, 12) {real, imag} */,
  {32'hc04121f4, 32'h00000000} /* (0, 19, 11) {real, imag} */,
  {32'hc0137c5e, 32'h00000000} /* (0, 19, 10) {real, imag} */,
  {32'h3f0818ca, 32'h00000000} /* (0, 19, 9) {real, imag} */,
  {32'hc06a495d, 32'h00000000} /* (0, 19, 8) {real, imag} */,
  {32'hc027abf8, 32'h00000000} /* (0, 19, 7) {real, imag} */,
  {32'h3f797ee8, 32'h00000000} /* (0, 19, 6) {real, imag} */,
  {32'h3d726290, 32'h00000000} /* (0, 19, 5) {real, imag} */,
  {32'hbf8405eb, 32'h00000000} /* (0, 19, 4) {real, imag} */,
  {32'hc02622b5, 32'h00000000} /* (0, 19, 3) {real, imag} */,
  {32'hbf9f2ffd, 32'h00000000} /* (0, 19, 2) {real, imag} */,
  {32'h3f79ca6a, 32'h00000000} /* (0, 19, 1) {real, imag} */,
  {32'hbf9c72e3, 32'h00000000} /* (0, 19, 0) {real, imag} */,
  {32'hbd863990, 32'h00000000} /* (0, 18, 31) {real, imag} */,
  {32'hbf7dee08, 32'h00000000} /* (0, 18, 30) {real, imag} */,
  {32'hbdade1f0, 32'h00000000} /* (0, 18, 29) {real, imag} */,
  {32'h3e3f1c0a, 32'h00000000} /* (0, 18, 28) {real, imag} */,
  {32'hc0141ebe, 32'h00000000} /* (0, 18, 27) {real, imag} */,
  {32'hbea2f10c, 32'h00000000} /* (0, 18, 26) {real, imag} */,
  {32'h40739c98, 32'h00000000} /* (0, 18, 25) {real, imag} */,
  {32'h3fdb7172, 32'h00000000} /* (0, 18, 24) {real, imag} */,
  {32'hc0656cc4, 32'h00000000} /* (0, 18, 23) {real, imag} */,
  {32'hc06d5dc1, 32'h00000000} /* (0, 18, 22) {real, imag} */,
  {32'hbeeabb64, 32'h00000000} /* (0, 18, 21) {real, imag} */,
  {32'h3f703a3b, 32'h00000000} /* (0, 18, 20) {real, imag} */,
  {32'h3ec5e06a, 32'h00000000} /* (0, 18, 19) {real, imag} */,
  {32'hc0501f86, 32'h00000000} /* (0, 18, 18) {real, imag} */,
  {32'hc03e69e0, 32'h00000000} /* (0, 18, 17) {real, imag} */,
  {32'h40035988, 32'h00000000} /* (0, 18, 16) {real, imag} */,
  {32'h3fc4a452, 32'h00000000} /* (0, 18, 15) {real, imag} */,
  {32'h40179352, 32'h00000000} /* (0, 18, 14) {real, imag} */,
  {32'h4060464d, 32'h00000000} /* (0, 18, 13) {real, imag} */,
  {32'h3f9b2f0a, 32'h00000000} /* (0, 18, 12) {real, imag} */,
  {32'hbef129d2, 32'h00000000} /* (0, 18, 11) {real, imag} */,
  {32'hbf03fddf, 32'h00000000} /* (0, 18, 10) {real, imag} */,
  {32'h3fd6ea06, 32'h00000000} /* (0, 18, 9) {real, imag} */,
  {32'h3eb4de2a, 32'h00000000} /* (0, 18, 8) {real, imag} */,
  {32'h3f873b09, 32'h00000000} /* (0, 18, 7) {real, imag} */,
  {32'hbfb4bc83, 32'h00000000} /* (0, 18, 6) {real, imag} */,
  {32'h3f5af476, 32'h00000000} /* (0, 18, 5) {real, imag} */,
  {32'h3eb2f1b8, 32'h00000000} /* (0, 18, 4) {real, imag} */,
  {32'hc0a570d4, 32'h00000000} /* (0, 18, 3) {real, imag} */,
  {32'h3f940be8, 32'h00000000} /* (0, 18, 2) {real, imag} */,
  {32'h40a5ab4c, 32'h00000000} /* (0, 18, 1) {real, imag} */,
  {32'h3f8be6aa, 32'h00000000} /* (0, 18, 0) {real, imag} */,
  {32'h400045be, 32'h00000000} /* (0, 17, 31) {real, imag} */,
  {32'hc08a2710, 32'h00000000} /* (0, 17, 30) {real, imag} */,
  {32'hc04ca0a6, 32'h00000000} /* (0, 17, 29) {real, imag} */,
  {32'hbfa3cc74, 32'h00000000} /* (0, 17, 28) {real, imag} */,
  {32'hc058773a, 32'h00000000} /* (0, 17, 27) {real, imag} */,
  {32'h3f6c2294, 32'h00000000} /* (0, 17, 26) {real, imag} */,
  {32'h40014f10, 32'h00000000} /* (0, 17, 25) {real, imag} */,
  {32'hbf3f235e, 32'h00000000} /* (0, 17, 24) {real, imag} */,
  {32'hbfdc1153, 32'h00000000} /* (0, 17, 23) {real, imag} */,
  {32'hbfe227da, 32'h00000000} /* (0, 17, 22) {real, imag} */,
  {32'hbffcb2b9, 32'h00000000} /* (0, 17, 21) {real, imag} */,
  {32'h3f5876e9, 32'h00000000} /* (0, 17, 20) {real, imag} */,
  {32'hbf390e43, 32'h00000000} /* (0, 17, 19) {real, imag} */,
  {32'hbf7e6f92, 32'h00000000} /* (0, 17, 18) {real, imag} */,
  {32'hbf8ec117, 32'h00000000} /* (0, 17, 17) {real, imag} */,
  {32'hc046c733, 32'h00000000} /* (0, 17, 16) {real, imag} */,
  {32'hbf2d6d26, 32'h00000000} /* (0, 17, 15) {real, imag} */,
  {32'h3fc28510, 32'h00000000} /* (0, 17, 14) {real, imag} */,
  {32'hbf4f6669, 32'h00000000} /* (0, 17, 13) {real, imag} */,
  {32'hbf022eec, 32'h00000000} /* (0, 17, 12) {real, imag} */,
  {32'hc060dc46, 32'h00000000} /* (0, 17, 11) {real, imag} */,
  {32'hbfa21f9c, 32'h00000000} /* (0, 17, 10) {real, imag} */,
  {32'h405ea072, 32'h00000000} /* (0, 17, 9) {real, imag} */,
  {32'h402a31d0, 32'h00000000} /* (0, 17, 8) {real, imag} */,
  {32'h3fc40516, 32'h00000000} /* (0, 17, 7) {real, imag} */,
  {32'hc086d5de, 32'h00000000} /* (0, 17, 6) {real, imag} */,
  {32'hbf6def1e, 32'h00000000} /* (0, 17, 5) {real, imag} */,
  {32'hbfdfd686, 32'h00000000} /* (0, 17, 4) {real, imag} */,
  {32'hc0decaba, 32'h00000000} /* (0, 17, 3) {real, imag} */,
  {32'hbfbe2d74, 32'h00000000} /* (0, 17, 2) {real, imag} */,
  {32'h406a4aae, 32'h00000000} /* (0, 17, 1) {real, imag} */,
  {32'h409d66f0, 32'h00000000} /* (0, 17, 0) {real, imag} */,
  {32'h4016b56a, 32'h00000000} /* (0, 16, 31) {real, imag} */,
  {32'hc0373a70, 32'h00000000} /* (0, 16, 30) {real, imag} */,
  {32'hbf0e1168, 32'h00000000} /* (0, 16, 29) {real, imag} */,
  {32'h3ed6e19e, 32'h00000000} /* (0, 16, 28) {real, imag} */,
  {32'hc03e6a24, 32'h00000000} /* (0, 16, 27) {real, imag} */,
  {32'h3ed76eec, 32'h00000000} /* (0, 16, 26) {real, imag} */,
  {32'hbea56086, 32'h00000000} /* (0, 16, 25) {real, imag} */,
  {32'hc01fca0e, 32'h00000000} /* (0, 16, 24) {real, imag} */,
  {32'h3f35083b, 32'h00000000} /* (0, 16, 23) {real, imag} */,
  {32'hbe27aab0, 32'h00000000} /* (0, 16, 22) {real, imag} */,
  {32'h4006ddb7, 32'h00000000} /* (0, 16, 21) {real, imag} */,
  {32'hbf8f8360, 32'h00000000} /* (0, 16, 20) {real, imag} */,
  {32'hc007529e, 32'h00000000} /* (0, 16, 19) {real, imag} */,
  {32'h40190ccc, 32'h00000000} /* (0, 16, 18) {real, imag} */,
  {32'h4000262a, 32'h00000000} /* (0, 16, 17) {real, imag} */,
  {32'h3d9f88b0, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'h3f27ba10, 32'h00000000} /* (0, 16, 15) {real, imag} */,
  {32'h3f8630a9, 32'h00000000} /* (0, 16, 14) {real, imag} */,
  {32'hbfd11f3a, 32'h00000000} /* (0, 16, 13) {real, imag} */,
  {32'hc07feeb2, 32'h00000000} /* (0, 16, 12) {real, imag} */,
  {32'hc0bccaba, 32'h00000000} /* (0, 16, 11) {real, imag} */,
  {32'hbe63abcc, 32'h00000000} /* (0, 16, 10) {real, imag} */,
  {32'h40dc5aea, 32'h00000000} /* (0, 16, 9) {real, imag} */,
  {32'h404ad3f2, 32'h00000000} /* (0, 16, 8) {real, imag} */,
  {32'h3f8a39a8, 32'h00000000} /* (0, 16, 7) {real, imag} */,
  {32'hbec64f50, 32'h00000000} /* (0, 16, 6) {real, imag} */,
  {32'h3ead22a0, 32'h00000000} /* (0, 16, 5) {real, imag} */,
  {32'hbf92f090, 32'h00000000} /* (0, 16, 4) {real, imag} */,
  {32'hc004d3da, 32'h00000000} /* (0, 16, 3) {real, imag} */,
  {32'hbfdc0e6c, 32'h00000000} /* (0, 16, 2) {real, imag} */,
  {32'hbf637c1a, 32'h00000000} /* (0, 16, 1) {real, imag} */,
  {32'h406c4afc, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h3f011650, 32'h00000000} /* (0, 15, 31) {real, imag} */,
  {32'hbfb4d63a, 32'h00000000} /* (0, 15, 30) {real, imag} */,
  {32'hbeba13e0, 32'h00000000} /* (0, 15, 29) {real, imag} */,
  {32'hbe1725ec, 32'h00000000} /* (0, 15, 28) {real, imag} */,
  {32'hbf348de2, 32'h00000000} /* (0, 15, 27) {real, imag} */,
  {32'hbf61fe78, 32'h00000000} /* (0, 15, 26) {real, imag} */,
  {32'hc0be02ca, 32'h00000000} /* (0, 15, 25) {real, imag} */,
  {32'hc00c356c, 32'h00000000} /* (0, 15, 24) {real, imag} */,
  {32'h3e9663d8, 32'h00000000} /* (0, 15, 23) {real, imag} */,
  {32'h3d0fadd0, 32'h00000000} /* (0, 15, 22) {real, imag} */,
  {32'h40db2c54, 32'h00000000} /* (0, 15, 21) {real, imag} */,
  {32'h3f9863d6, 32'h00000000} /* (0, 15, 20) {real, imag} */,
  {32'hc0201f6c, 32'h00000000} /* (0, 15, 19) {real, imag} */,
  {32'h4004dddc, 32'h00000000} /* (0, 15, 18) {real, imag} */,
  {32'h3e85f9b4, 32'h00000000} /* (0, 15, 17) {real, imag} */,
  {32'h409c7384, 32'h00000000} /* (0, 15, 16) {real, imag} */,
  {32'h402e50b2, 32'h00000000} /* (0, 15, 15) {real, imag} */,
  {32'hbef5ec0c, 32'h00000000} /* (0, 15, 14) {real, imag} */,
  {32'hc03deee8, 32'h00000000} /* (0, 15, 13) {real, imag} */,
  {32'hc0b24692, 32'h00000000} /* (0, 15, 12) {real, imag} */,
  {32'hc09524ba, 32'h00000000} /* (0, 15, 11) {real, imag} */,
  {32'hbfa2fcf2, 32'h00000000} /* (0, 15, 10) {real, imag} */,
  {32'h3ff0acf0, 32'h00000000} /* (0, 15, 9) {real, imag} */,
  {32'hc0172536, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'hc0ba352e, 32'h00000000} /* (0, 15, 7) {real, imag} */,
  {32'hc0a745de, 32'h00000000} /* (0, 15, 6) {real, imag} */,
  {32'hbf98d0b9, 32'h00000000} /* (0, 15, 5) {real, imag} */,
  {32'h4040c04c, 32'h00000000} /* (0, 15, 4) {real, imag} */,
  {32'h400dffde, 32'h00000000} /* (0, 15, 3) {real, imag} */,
  {32'hbffc1ccd, 32'h00000000} /* (0, 15, 2) {real, imag} */,
  {32'hc052765a, 32'h00000000} /* (0, 15, 1) {real, imag} */,
  {32'hc0011eac, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'hbe326638, 32'h00000000} /* (0, 14, 31) {real, imag} */,
  {32'hc03e23fb, 32'h00000000} /* (0, 14, 30) {real, imag} */,
  {32'hbf83251e, 32'h00000000} /* (0, 14, 29) {real, imag} */,
  {32'hbfdfbf1b, 32'h00000000} /* (0, 14, 28) {real, imag} */,
  {32'hbfc967e0, 32'h00000000} /* (0, 14, 27) {real, imag} */,
  {32'h3edde2a4, 32'h00000000} /* (0, 14, 26) {real, imag} */,
  {32'hc0dd59f5, 32'h00000000} /* (0, 14, 25) {real, imag} */,
  {32'hc070c146, 32'h00000000} /* (0, 14, 24) {real, imag} */,
  {32'hbf107afe, 32'h00000000} /* (0, 14, 23) {real, imag} */,
  {32'h4008fa61, 32'h00000000} /* (0, 14, 22) {real, imag} */,
  {32'h40196fee, 32'h00000000} /* (0, 14, 21) {real, imag} */,
  {32'hbf30f81e, 32'h00000000} /* (0, 14, 20) {real, imag} */,
  {32'hc0b6c294, 32'h00000000} /* (0, 14, 19) {real, imag} */,
  {32'hbf3fac58, 32'h00000000} /* (0, 14, 18) {real, imag} */,
  {32'hc02fd746, 32'h00000000} /* (0, 14, 17) {real, imag} */,
  {32'h3f61529c, 32'h00000000} /* (0, 14, 16) {real, imag} */,
  {32'h4018b1f2, 32'h00000000} /* (0, 14, 15) {real, imag} */,
  {32'hbdf05840, 32'h00000000} /* (0, 14, 14) {real, imag} */,
  {32'hbf99d460, 32'h00000000} /* (0, 14, 13) {real, imag} */,
  {32'hbf53fdf1, 32'h00000000} /* (0, 14, 12) {real, imag} */,
  {32'h3fc89f75, 32'h00000000} /* (0, 14, 11) {real, imag} */,
  {32'h3fa882f6, 32'h00000000} /* (0, 14, 10) {real, imag} */,
  {32'hbf2e7369, 32'h00000000} /* (0, 14, 9) {real, imag} */,
  {32'h3ff3e620, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'hc048fb78, 32'h00000000} /* (0, 14, 7) {real, imag} */,
  {32'hc0849969, 32'h00000000} /* (0, 14, 6) {real, imag} */,
  {32'hbeee3714, 32'h00000000} /* (0, 14, 5) {real, imag} */,
  {32'h4018eb3d, 32'h00000000} /* (0, 14, 4) {real, imag} */,
  {32'h3ebd2380, 32'h00000000} /* (0, 14, 3) {real, imag} */,
  {32'hbfd567b9, 32'h00000000} /* (0, 14, 2) {real, imag} */,
  {32'hbfca18a9, 32'h00000000} /* (0, 14, 1) {real, imag} */,
  {32'hbfc78232, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'hc01a9510, 32'h00000000} /* (0, 13, 31) {real, imag} */,
  {32'hc07afeb7, 32'h00000000} /* (0, 13, 30) {real, imag} */,
  {32'h403448d7, 32'h00000000} /* (0, 13, 29) {real, imag} */,
  {32'h40691f18, 32'h00000000} /* (0, 13, 28) {real, imag} */,
  {32'h405fc07a, 32'h00000000} /* (0, 13, 27) {real, imag} */,
  {32'h40b3e6cb, 32'h00000000} /* (0, 13, 26) {real, imag} */,
  {32'hc03ded18, 32'h00000000} /* (0, 13, 25) {real, imag} */,
  {32'hc0db6591, 32'h00000000} /* (0, 13, 24) {real, imag} */,
  {32'hbf19f535, 32'h00000000} /* (0, 13, 23) {real, imag} */,
  {32'h405a6d83, 32'h00000000} /* (0, 13, 22) {real, imag} */,
  {32'h3ef12d20, 32'h00000000} /* (0, 13, 21) {real, imag} */,
  {32'hc050fcc8, 32'h00000000} /* (0, 13, 20) {real, imag} */,
  {32'hc09d0b63, 32'h00000000} /* (0, 13, 19) {real, imag} */,
  {32'h3fe6f6a1, 32'h00000000} /* (0, 13, 18) {real, imag} */,
  {32'hc035c8c9, 32'h00000000} /* (0, 13, 17) {real, imag} */,
  {32'hc044f82e, 32'h00000000} /* (0, 13, 16) {real, imag} */,
  {32'h401b160f, 32'h00000000} /* (0, 13, 15) {real, imag} */,
  {32'hc01d1f90, 32'h00000000} /* (0, 13, 14) {real, imag} */,
  {32'hc043d782, 32'h00000000} /* (0, 13, 13) {real, imag} */,
  {32'h3fcfcb56, 32'h00000000} /* (0, 13, 12) {real, imag} */,
  {32'h3fd6505a, 32'h00000000} /* (0, 13, 11) {real, imag} */,
  {32'h3eec7671, 32'h00000000} /* (0, 13, 10) {real, imag} */,
  {32'hc0504f39, 32'h00000000} /* (0, 13, 9) {real, imag} */,
  {32'h40171f57, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'hbfac1a9e, 32'h00000000} /* (0, 13, 7) {real, imag} */,
  {32'hc0887325, 32'h00000000} /* (0, 13, 6) {real, imag} */,
  {32'h3f69a6d1, 32'h00000000} /* (0, 13, 5) {real, imag} */,
  {32'h3e26ba58, 32'h00000000} /* (0, 13, 4) {real, imag} */,
  {32'hc0563c70, 32'h00000000} /* (0, 13, 3) {real, imag} */,
  {32'hbe9bc0b0, 32'h00000000} /* (0, 13, 2) {real, imag} */,
  {32'h3fb83808, 32'h00000000} /* (0, 13, 1) {real, imag} */,
  {32'h3f552817, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'hbfbccf34, 32'h00000000} /* (0, 12, 31) {real, imag} */,
  {32'hc04a990e, 32'h00000000} /* (0, 12, 30) {real, imag} */,
  {32'hbfb2b186, 32'h00000000} /* (0, 12, 29) {real, imag} */,
  {32'h3ed3b366, 32'h00000000} /* (0, 12, 28) {real, imag} */,
  {32'h3d176e20, 32'h00000000} /* (0, 12, 27) {real, imag} */,
  {32'hbf196dbd, 32'h00000000} /* (0, 12, 26) {real, imag} */,
  {32'hc0126309, 32'h00000000} /* (0, 12, 25) {real, imag} */,
  {32'hc033d738, 32'h00000000} /* (0, 12, 24) {real, imag} */,
  {32'h4068aeae, 32'h00000000} /* (0, 12, 23) {real, imag} */,
  {32'h40d5c40b, 32'h00000000} /* (0, 12, 22) {real, imag} */,
  {32'h407c79d4, 32'h00000000} /* (0, 12, 21) {real, imag} */,
  {32'hbf994ab6, 32'h00000000} /* (0, 12, 20) {real, imag} */,
  {32'hc066154f, 32'h00000000} /* (0, 12, 19) {real, imag} */,
  {32'hbf108d4b, 32'h00000000} /* (0, 12, 18) {real, imag} */,
  {32'hbbeb5e00, 32'h00000000} /* (0, 12, 17) {real, imag} */,
  {32'hbe344fe0, 32'h00000000} /* (0, 12, 16) {real, imag} */,
  {32'hc00f505e, 32'h00000000} /* (0, 12, 15) {real, imag} */,
  {32'hc080d4d8, 32'h00000000} /* (0, 12, 14) {real, imag} */,
  {32'hbf37e591, 32'h00000000} /* (0, 12, 13) {real, imag} */,
  {32'h4052bafd, 32'h00000000} /* (0, 12, 12) {real, imag} */,
  {32'h3ff83185, 32'h00000000} /* (0, 12, 11) {real, imag} */,
  {32'h407c0d9d, 32'h00000000} /* (0, 12, 10) {real, imag} */,
  {32'hbf7a7ab1, 32'h00000000} /* (0, 12, 9) {real, imag} */,
  {32'h3f0c4488, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'h3fcd6178, 32'h00000000} /* (0, 12, 7) {real, imag} */,
  {32'hc036c1b8, 32'h00000000} /* (0, 12, 6) {real, imag} */,
  {32'hbf624bfc, 32'h00000000} /* (0, 12, 5) {real, imag} */,
  {32'h3ed9e3b4, 32'h00000000} /* (0, 12, 4) {real, imag} */,
  {32'hbf0e3047, 32'h00000000} /* (0, 12, 3) {real, imag} */,
  {32'h3fc1569e, 32'h00000000} /* (0, 12, 2) {real, imag} */,
  {32'h4024b154, 32'h00000000} /* (0, 12, 1) {real, imag} */,
  {32'h3f96e8f7, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h40762173, 32'h00000000} /* (0, 11, 31) {real, imag} */,
  {32'h40d3071d, 32'h00000000} /* (0, 11, 30) {real, imag} */,
  {32'h3f3bf165, 32'h00000000} /* (0, 11, 29) {real, imag} */,
  {32'hbe3fbedc, 32'h00000000} /* (0, 11, 28) {real, imag} */,
  {32'hbf95fc88, 32'h00000000} /* (0, 11, 27) {real, imag} */,
  {32'hc019f508, 32'h00000000} /* (0, 11, 26) {real, imag} */,
  {32'hbf3889dc, 32'h00000000} /* (0, 11, 25) {real, imag} */,
  {32'h3fa23b06, 32'h00000000} /* (0, 11, 24) {real, imag} */,
  {32'h4049ca48, 32'h00000000} /* (0, 11, 23) {real, imag} */,
  {32'h40ff39cc, 32'h00000000} /* (0, 11, 22) {real, imag} */,
  {32'h4067cd98, 32'h00000000} /* (0, 11, 21) {real, imag} */,
  {32'hbfa9764f, 32'h00000000} /* (0, 11, 20) {real, imag} */,
  {32'hc084c7c2, 32'h00000000} /* (0, 11, 19) {real, imag} */,
  {32'hbfd71d25, 32'h00000000} /* (0, 11, 18) {real, imag} */,
  {32'h400c8b4a, 32'h00000000} /* (0, 11, 17) {real, imag} */,
  {32'h40917e0f, 32'h00000000} /* (0, 11, 16) {real, imag} */,
  {32'hbf9c005c, 32'h00000000} /* (0, 11, 15) {real, imag} */,
  {32'h3f3dd080, 32'h00000000} /* (0, 11, 14) {real, imag} */,
  {32'h3ffa46b6, 32'h00000000} /* (0, 11, 13) {real, imag} */,
  {32'h3833e000, 32'h00000000} /* (0, 11, 12) {real, imag} */,
  {32'h3fa5fb44, 32'h00000000} /* (0, 11, 11) {real, imag} */,
  {32'h3fccff1a, 32'h00000000} /* (0, 11, 10) {real, imag} */,
  {32'h3f157817, 32'h00000000} /* (0, 11, 9) {real, imag} */,
  {32'h4068d354, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'h40d0fbbc, 32'h00000000} /* (0, 11, 7) {real, imag} */,
  {32'h3f813a74, 32'h00000000} /* (0, 11, 6) {real, imag} */,
  {32'h3fc16bd2, 32'h00000000} /* (0, 11, 5) {real, imag} */,
  {32'h402bf3ff, 32'h00000000} /* (0, 11, 4) {real, imag} */,
  {32'hbffa2a0c, 32'h00000000} /* (0, 11, 3) {real, imag} */,
  {32'hbfa5367b, 32'h00000000} /* (0, 11, 2) {real, imag} */,
  {32'h3fce1580, 32'h00000000} /* (0, 11, 1) {real, imag} */,
  {32'h400ae074, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h40845d1c, 32'h00000000} /* (0, 10, 31) {real, imag} */,
  {32'h40aaae3a, 32'h00000000} /* (0, 10, 30) {real, imag} */,
  {32'h408b54d6, 32'h00000000} /* (0, 10, 29) {real, imag} */,
  {32'h40696b90, 32'h00000000} /* (0, 10, 28) {real, imag} */,
  {32'hbe14cd80, 32'h00000000} /* (0, 10, 27) {real, imag} */,
  {32'hc0691426, 32'h00000000} /* (0, 10, 26) {real, imag} */,
  {32'h3f136705, 32'h00000000} /* (0, 10, 25) {real, imag} */,
  {32'h3f96052c, 32'h00000000} /* (0, 10, 24) {real, imag} */,
  {32'hbe04694c, 32'h00000000} /* (0, 10, 23) {real, imag} */,
  {32'h4025be35, 32'h00000000} /* (0, 10, 22) {real, imag} */,
  {32'hc0645348, 32'h00000000} /* (0, 10, 21) {real, imag} */,
  {32'h3e82b658, 32'h00000000} /* (0, 10, 20) {real, imag} */,
  {32'hbfb4dfb7, 32'h00000000} /* (0, 10, 19) {real, imag} */,
  {32'hc07b0e06, 32'h00000000} /* (0, 10, 18) {real, imag} */,
  {32'hbc70ee00, 32'h00000000} /* (0, 10, 17) {real, imag} */,
  {32'h407fc4e5, 32'h00000000} /* (0, 10, 16) {real, imag} */,
  {32'h401b2950, 32'h00000000} /* (0, 10, 15) {real, imag} */,
  {32'h3f8b2138, 32'h00000000} /* (0, 10, 14) {real, imag} */,
  {32'hbe8f2e9d, 32'h00000000} /* (0, 10, 13) {real, imag} */,
  {32'hbfb45762, 32'h00000000} /* (0, 10, 12) {real, imag} */,
  {32'hbeb3a3ca, 32'h00000000} /* (0, 10, 11) {real, imag} */,
  {32'hbfd8d76e, 32'h00000000} /* (0, 10, 10) {real, imag} */,
  {32'hc0569734, 32'h00000000} /* (0, 10, 9) {real, imag} */,
  {32'h3fafe321, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'h4103aa31, 32'h00000000} /* (0, 10, 7) {real, imag} */,
  {32'h4081ae96, 32'h00000000} /* (0, 10, 6) {real, imag} */,
  {32'h40a57dea, 32'h00000000} /* (0, 10, 5) {real, imag} */,
  {32'h40345f06, 32'h00000000} /* (0, 10, 4) {real, imag} */,
  {32'hc08da3a6, 32'h00000000} /* (0, 10, 3) {real, imag} */,
  {32'hc07d42de, 32'h00000000} /* (0, 10, 2) {real, imag} */,
  {32'h3f1db5e4, 32'h00000000} /* (0, 10, 1) {real, imag} */,
  {32'h3ff7ed3a, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'h3faac776, 32'h00000000} /* (0, 9, 31) {real, imag} */,
  {32'hbdf4d540, 32'h00000000} /* (0, 9, 30) {real, imag} */,
  {32'h405695c8, 32'h00000000} /* (0, 9, 29) {real, imag} */,
  {32'h407e7cf7, 32'h00000000} /* (0, 9, 28) {real, imag} */,
  {32'h3fa1e7dc, 32'h00000000} /* (0, 9, 27) {real, imag} */,
  {32'hbe4d9f48, 32'h00000000} /* (0, 9, 26) {real, imag} */,
  {32'h404af54e, 32'h00000000} /* (0, 9, 25) {real, imag} */,
  {32'h405531c6, 32'h00000000} /* (0, 9, 24) {real, imag} */,
  {32'h3f9030fc, 32'h00000000} /* (0, 9, 23) {real, imag} */,
  {32'h3f8d0e62, 32'h00000000} /* (0, 9, 22) {real, imag} */,
  {32'hbfb3524c, 32'h00000000} /* (0, 9, 21) {real, imag} */,
  {32'h3fcc8e4c, 32'h00000000} /* (0, 9, 20) {real, imag} */,
  {32'h3f3e0e25, 32'h00000000} /* (0, 9, 19) {real, imag} */,
  {32'hc015d8c6, 32'h00000000} /* (0, 9, 18) {real, imag} */,
  {32'hbff3d4aa, 32'h00000000} /* (0, 9, 17) {real, imag} */,
  {32'h3f88126c, 32'h00000000} /* (0, 9, 16) {real, imag} */,
  {32'h40895a1a, 32'h00000000} /* (0, 9, 15) {real, imag} */,
  {32'h3fc8f958, 32'h00000000} /* (0, 9, 14) {real, imag} */,
  {32'hc03ac079, 32'h00000000} /* (0, 9, 13) {real, imag} */,
  {32'h3fcbe4d2, 32'h00000000} /* (0, 9, 12) {real, imag} */,
  {32'h400d9e62, 32'h00000000} /* (0, 9, 11) {real, imag} */,
  {32'hbf9c46d8, 32'h00000000} /* (0, 9, 10) {real, imag} */,
  {32'hc058214e, 32'h00000000} /* (0, 9, 9) {real, imag} */,
  {32'hbf7abae8, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'h408360e8, 32'h00000000} /* (0, 9, 7) {real, imag} */,
  {32'hbf043fad, 32'h00000000} /* (0, 9, 6) {real, imag} */,
  {32'hbfdc06d5, 32'h00000000} /* (0, 9, 5) {real, imag} */,
  {32'hbf0499a5, 32'h00000000} /* (0, 9, 4) {real, imag} */,
  {32'hbed0b70c, 32'h00000000} /* (0, 9, 3) {real, imag} */,
  {32'hc02a9d6c, 32'h00000000} /* (0, 9, 2) {real, imag} */,
  {32'hbdbfc1b0, 32'h00000000} /* (0, 9, 1) {real, imag} */,
  {32'hbe137aa0, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'hbf1e9adc, 32'h00000000} /* (0, 8, 31) {real, imag} */,
  {32'hbf302852, 32'h00000000} /* (0, 8, 30) {real, imag} */,
  {32'hbfdaca7f, 32'h00000000} /* (0, 8, 29) {real, imag} */,
  {32'hc06bc200, 32'h00000000} /* (0, 8, 28) {real, imag} */,
  {32'h3f88d536, 32'h00000000} /* (0, 8, 27) {real, imag} */,
  {32'h3f1bcab9, 32'h00000000} /* (0, 8, 26) {real, imag} */,
  {32'hc05f554d, 32'h00000000} /* (0, 8, 25) {real, imag} */,
  {32'h3fe7cfee, 32'h00000000} /* (0, 8, 24) {real, imag} */,
  {32'h3fc010e7, 32'h00000000} /* (0, 8, 23) {real, imag} */,
  {32'h3fb63e9e, 32'h00000000} /* (0, 8, 22) {real, imag} */,
  {32'hbf6366cb, 32'h00000000} /* (0, 8, 21) {real, imag} */,
  {32'h3fa40222, 32'h00000000} /* (0, 8, 20) {real, imag} */,
  {32'h4040428f, 32'h00000000} /* (0, 8, 19) {real, imag} */,
  {32'hbf85eb60, 32'h00000000} /* (0, 8, 18) {real, imag} */,
  {32'hbee75f4e, 32'h00000000} /* (0, 8, 17) {real, imag} */,
  {32'h3fec45c9, 32'h00000000} /* (0, 8, 16) {real, imag} */,
  {32'h4011182c, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'hc0071d8c, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'hc04b90f2, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'h3f693770, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'hbfcf1aca, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'hc0270a50, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hc00ec354, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'hbf74d45c, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'h40200bc9, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hbdde66a0, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'hc081d0bc, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'hbf922e63, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'h3fcded0a, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'hbf28d64b, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'hbf588450, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'hbf8ee719, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h3e530ee4, 32'h00000000} /* (0, 7, 31) {real, imag} */,
  {32'hbfad5060, 32'h00000000} /* (0, 7, 30) {real, imag} */,
  {32'hc0a292c4, 32'h00000000} /* (0, 7, 29) {real, imag} */,
  {32'hc0e32b51, 32'h00000000} /* (0, 7, 28) {real, imag} */,
  {32'hc03a0d4e, 32'h00000000} /* (0, 7, 27) {real, imag} */,
  {32'hc09e9819, 32'h00000000} /* (0, 7, 26) {real, imag} */,
  {32'hc1205b46, 32'h00000000} /* (0, 7, 25) {real, imag} */,
  {32'hc0917553, 32'h00000000} /* (0, 7, 24) {real, imag} */,
  {32'h3f0ee442, 32'h00000000} /* (0, 7, 23) {real, imag} */,
  {32'h40670dfc, 32'h00000000} /* (0, 7, 22) {real, imag} */,
  {32'hbf8a382a, 32'h00000000} /* (0, 7, 21) {real, imag} */,
  {32'h3fa5141a, 32'h00000000} /* (0, 7, 20) {real, imag} */,
  {32'h3f276acb, 32'h00000000} /* (0, 7, 19) {real, imag} */,
  {32'hbf9236ec, 32'h00000000} /* (0, 7, 18) {real, imag} */,
  {32'h4006c8ac, 32'h00000000} /* (0, 7, 17) {real, imag} */,
  {32'h3ece57f4, 32'h00000000} /* (0, 7, 16) {real, imag} */,
  {32'hbea76da2, 32'h00000000} /* (0, 7, 15) {real, imag} */,
  {32'hbf6141b6, 32'h00000000} /* (0, 7, 14) {real, imag} */,
  {32'hc021b134, 32'h00000000} /* (0, 7, 13) {real, imag} */,
  {32'hbe9196ae, 32'h00000000} /* (0, 7, 12) {real, imag} */,
  {32'hc041f979, 32'h00000000} /* (0, 7, 11) {real, imag} */,
  {32'hc04a8ac1, 32'h00000000} /* (0, 7, 10) {real, imag} */,
  {32'hc013d7a1, 32'h00000000} /* (0, 7, 9) {real, imag} */,
  {32'h4089985c, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'h40d3b218, 32'h00000000} /* (0, 7, 7) {real, imag} */,
  {32'hc030ba35, 32'h00000000} /* (0, 7, 6) {real, imag} */,
  {32'hc0291e92, 32'h00000000} /* (0, 7, 5) {real, imag} */,
  {32'h3f7ad5f0, 32'h00000000} /* (0, 7, 4) {real, imag} */,
  {32'h402d4c60, 32'h00000000} /* (0, 7, 3) {real, imag} */,
  {32'hbf69edee, 32'h00000000} /* (0, 7, 2) {real, imag} */,
  {32'hc01fd64c, 32'h00000000} /* (0, 7, 1) {real, imag} */,
  {32'hbe442410, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'h3fc4c88b, 32'h00000000} /* (0, 6, 31) {real, imag} */,
  {32'hbf04938b, 32'h00000000} /* (0, 6, 30) {real, imag} */,
  {32'hc08d5251, 32'h00000000} /* (0, 6, 29) {real, imag} */,
  {32'hc06638c6, 32'h00000000} /* (0, 6, 28) {real, imag} */,
  {32'h401c161c, 32'h00000000} /* (0, 6, 27) {real, imag} */,
  {32'h3f225892, 32'h00000000} /* (0, 6, 26) {real, imag} */,
  {32'hc0783e91, 32'h00000000} /* (0, 6, 25) {real, imag} */,
  {32'hc00ce397, 32'h00000000} /* (0, 6, 24) {real, imag} */,
  {32'h404ceb04, 32'h00000000} /* (0, 6, 23) {real, imag} */,
  {32'h408b8741, 32'h00000000} /* (0, 6, 22) {real, imag} */,
  {32'h3fe45132, 32'h00000000} /* (0, 6, 21) {real, imag} */,
  {32'h3f4ef8ed, 32'h00000000} /* (0, 6, 20) {real, imag} */,
  {32'hbe7cf484, 32'h00000000} /* (0, 6, 19) {real, imag} */,
  {32'hc02dce8e, 32'h00000000} /* (0, 6, 18) {real, imag} */,
  {32'hbf600661, 32'h00000000} /* (0, 6, 17) {real, imag} */,
  {32'h3ebec7f2, 32'h00000000} /* (0, 6, 16) {real, imag} */,
  {32'h40333484, 32'h00000000} /* (0, 6, 15) {real, imag} */,
  {32'h4004356d, 32'h00000000} /* (0, 6, 14) {real, imag} */,
  {32'hbc5c8280, 32'h00000000} /* (0, 6, 13) {real, imag} */,
  {32'h3f032c0a, 32'h00000000} /* (0, 6, 12) {real, imag} */,
  {32'hc04a8fc9, 32'h00000000} /* (0, 6, 11) {real, imag} */,
  {32'hbed36008, 32'h00000000} /* (0, 6, 10) {real, imag} */,
  {32'hc01f13c6, 32'h00000000} /* (0, 6, 9) {real, imag} */,
  {32'h4024a20a, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'h408f849d, 32'h00000000} /* (0, 6, 7) {real, imag} */,
  {32'hc00679d5, 32'h00000000} /* (0, 6, 6) {real, imag} */,
  {32'h40a061c5, 32'h00000000} /* (0, 6, 5) {real, imag} */,
  {32'h40b896c1, 32'h00000000} /* (0, 6, 4) {real, imag} */,
  {32'hbef53b8e, 32'h00000000} /* (0, 6, 3) {real, imag} */,
  {32'hbec94cb2, 32'h00000000} /* (0, 6, 2) {real, imag} */,
  {32'h40244cf6, 32'h00000000} /* (0, 6, 1) {real, imag} */,
  {32'h3f9601d0, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hbf655d5e, 32'h00000000} /* (0, 5, 31) {real, imag} */,
  {32'hc067d8c4, 32'h00000000} /* (0, 5, 30) {real, imag} */,
  {32'hc05c273b, 32'h00000000} /* (0, 5, 29) {real, imag} */,
  {32'h3f991867, 32'h00000000} /* (0, 5, 28) {real, imag} */,
  {32'h406cbd1b, 32'h00000000} /* (0, 5, 27) {real, imag} */,
  {32'h3f9d755d, 32'h00000000} /* (0, 5, 26) {real, imag} */,
  {32'hc0431ff8, 32'h00000000} /* (0, 5, 25) {real, imag} */,
  {32'hc025240f, 32'h00000000} /* (0, 5, 24) {real, imag} */,
  {32'h402d0301, 32'h00000000} /* (0, 5, 23) {real, imag} */,
  {32'h409a2140, 32'h00000000} /* (0, 5, 22) {real, imag} */,
  {32'h40a20ca3, 32'h00000000} /* (0, 5, 21) {real, imag} */,
  {32'h40204ebc, 32'h00000000} /* (0, 5, 20) {real, imag} */,
  {32'h3f84461e, 32'h00000000} /* (0, 5, 19) {real, imag} */,
  {32'hbf221b7e, 32'h00000000} /* (0, 5, 18) {real, imag} */,
  {32'hbf46d66d, 32'h00000000} /* (0, 5, 17) {real, imag} */,
  {32'hbf851500, 32'h00000000} /* (0, 5, 16) {real, imag} */,
  {32'hc057b8d1, 32'h00000000} /* (0, 5, 15) {real, imag} */,
  {32'hc06b4f37, 32'h00000000} /* (0, 5, 14) {real, imag} */,
  {32'hbf3f594f, 32'h00000000} /* (0, 5, 13) {real, imag} */,
  {32'hbf88baa8, 32'h00000000} /* (0, 5, 12) {real, imag} */,
  {32'hc0c1dd20, 32'h00000000} /* (0, 5, 11) {real, imag} */,
  {32'h3fc35cfa, 32'h00000000} /* (0, 5, 10) {real, imag} */,
  {32'h3dd5f06c, 32'h00000000} /* (0, 5, 9) {real, imag} */,
  {32'h3fc79ca4, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'h3ff8a664, 32'h00000000} /* (0, 5, 7) {real, imag} */,
  {32'hbca53de0, 32'h00000000} /* (0, 5, 6) {real, imag} */,
  {32'h407877d4, 32'h00000000} /* (0, 5, 5) {real, imag} */,
  {32'h3ffce4fe, 32'h00000000} /* (0, 5, 4) {real, imag} */,
  {32'hc01256aa, 32'h00000000} /* (0, 5, 3) {real, imag} */,
  {32'h3f455000, 32'h00000000} /* (0, 5, 2) {real, imag} */,
  {32'h408344a4, 32'h00000000} /* (0, 5, 1) {real, imag} */,
  {32'h3f9983ac, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hc00e78fa, 32'h00000000} /* (0, 4, 31) {real, imag} */,
  {32'hc0b79553, 32'h00000000} /* (0, 4, 30) {real, imag} */,
  {32'hc0ea720a, 32'h00000000} /* (0, 4, 29) {real, imag} */,
  {32'hbfef3212, 32'h00000000} /* (0, 4, 28) {real, imag} */,
  {32'hbc2f8900, 32'h00000000} /* (0, 4, 27) {real, imag} */,
  {32'hc00322f0, 32'h00000000} /* (0, 4, 26) {real, imag} */,
  {32'hc0a6004e, 32'h00000000} /* (0, 4, 25) {real, imag} */,
  {32'hc0f940a2, 32'h00000000} /* (0, 4, 24) {real, imag} */,
  {32'hbf79cf47, 32'h00000000} /* (0, 4, 23) {real, imag} */,
  {32'h40ecc214, 32'h00000000} /* (0, 4, 22) {real, imag} */,
  {32'h40e4add7, 32'h00000000} /* (0, 4, 21) {real, imag} */,
  {32'h3fd0d3ad, 32'h00000000} /* (0, 4, 20) {real, imag} */,
  {32'hc049b9d6, 32'h00000000} /* (0, 4, 19) {real, imag} */,
  {32'h40432cff, 32'h00000000} /* (0, 4, 18) {real, imag} */,
  {32'h403f942a, 32'h00000000} /* (0, 4, 17) {real, imag} */,
  {32'hbfdecee4, 32'h00000000} /* (0, 4, 16) {real, imag} */,
  {32'hc0b54f9b, 32'h00000000} /* (0, 4, 15) {real, imag} */,
  {32'h3ef9f004, 32'h00000000} /* (0, 4, 14) {real, imag} */,
  {32'h3f90562b, 32'h00000000} /* (0, 4, 13) {real, imag} */,
  {32'hc018e2bb, 32'h00000000} /* (0, 4, 12) {real, imag} */,
  {32'hc07ca5d9, 32'h00000000} /* (0, 4, 11) {real, imag} */,
  {32'h3f9afc8e, 32'h00000000} /* (0, 4, 10) {real, imag} */,
  {32'h407204a2, 32'h00000000} /* (0, 4, 9) {real, imag} */,
  {32'h408ff843, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'h40b1f41b, 32'h00000000} /* (0, 4, 7) {real, imag} */,
  {32'h409ed874, 32'h00000000} /* (0, 4, 6) {real, imag} */,
  {32'h40675f62, 32'h00000000} /* (0, 4, 5) {real, imag} */,
  {32'h3ed95b5a, 32'h00000000} /* (0, 4, 4) {real, imag} */,
  {32'hbe5bf098, 32'h00000000} /* (0, 4, 3) {real, imag} */,
  {32'h400ebc68, 32'h00000000} /* (0, 4, 2) {real, imag} */,
  {32'h40320548, 32'h00000000} /* (0, 4, 1) {real, imag} */,
  {32'h3ffbe14d, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hbeb6baca, 32'h00000000} /* (0, 3, 31) {real, imag} */,
  {32'hc015e929, 32'h00000000} /* (0, 3, 30) {real, imag} */,
  {32'hc02b3892, 32'h00000000} /* (0, 3, 29) {real, imag} */,
  {32'h3ec07364, 32'h00000000} /* (0, 3, 28) {real, imag} */,
  {32'h3e805ad8, 32'h00000000} /* (0, 3, 27) {real, imag} */,
  {32'h3fb20c22, 32'h00000000} /* (0, 3, 26) {real, imag} */,
  {32'h3e293784, 32'h00000000} /* (0, 3, 25) {real, imag} */,
  {32'hbf8f8aaa, 32'h00000000} /* (0, 3, 24) {real, imag} */,
  {32'hc0938893, 32'h00000000} /* (0, 3, 23) {real, imag} */,
  {32'hbe408bd0, 32'h00000000} /* (0, 3, 22) {real, imag} */,
  {32'h403b25d7, 32'h00000000} /* (0, 3, 21) {real, imag} */,
  {32'h3eb14668, 32'h00000000} /* (0, 3, 20) {real, imag} */,
  {32'hc014bdf2, 32'h00000000} /* (0, 3, 19) {real, imag} */,
  {32'hbf8eaae7, 32'h00000000} /* (0, 3, 18) {real, imag} */,
  {32'hc00ab022, 32'h00000000} /* (0, 3, 17) {real, imag} */,
  {32'hc0771941, 32'h00000000} /* (0, 3, 16) {real, imag} */,
  {32'hc00aa00b, 32'h00000000} /* (0, 3, 15) {real, imag} */,
  {32'h40895609, 32'h00000000} /* (0, 3, 14) {real, imag} */,
  {32'h408acce4, 32'h00000000} /* (0, 3, 13) {real, imag} */,
  {32'h3c393f80, 32'h00000000} /* (0, 3, 12) {real, imag} */,
  {32'h3ea51a32, 32'h00000000} /* (0, 3, 11) {real, imag} */,
  {32'h3fc9cc9d, 32'h00000000} /* (0, 3, 10) {real, imag} */,
  {32'h3f5a13d2, 32'h00000000} /* (0, 3, 9) {real, imag} */,
  {32'h3fd8229e, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h405c9c49, 32'h00000000} /* (0, 3, 7) {real, imag} */,
  {32'hbe97778a, 32'h00000000} /* (0, 3, 6) {real, imag} */,
  {32'hbfb7062e, 32'h00000000} /* (0, 3, 5) {real, imag} */,
  {32'h3f15bf9b, 32'h00000000} /* (0, 3, 4) {real, imag} */,
  {32'hbf4da2d7, 32'h00000000} /* (0, 3, 3) {real, imag} */,
  {32'hbcc17080, 32'h00000000} /* (0, 3, 2) {real, imag} */,
  {32'hbf4b19b6, 32'h00000000} /* (0, 3, 1) {real, imag} */,
  {32'h4022c48e, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'h3fe98aa4, 32'h00000000} /* (0, 2, 31) {real, imag} */,
  {32'h403460f1, 32'h00000000} /* (0, 2, 30) {real, imag} */,
  {32'h3f8c5278, 32'h00000000} /* (0, 2, 29) {real, imag} */,
  {32'h3ec47898, 32'h00000000} /* (0, 2, 28) {real, imag} */,
  {32'hbf37037c, 32'h00000000} /* (0, 2, 27) {real, imag} */,
  {32'hbf0650f0, 32'h00000000} /* (0, 2, 26) {real, imag} */,
  {32'h3fee8234, 32'h00000000} /* (0, 2, 25) {real, imag} */,
  {32'h40fef2e5, 32'h00000000} /* (0, 2, 24) {real, imag} */,
  {32'h3e87e02c, 32'h00000000} /* (0, 2, 23) {real, imag} */,
  {32'hbdc6a258, 32'h00000000} /* (0, 2, 22) {real, imag} */,
  {32'h402721b2, 32'h00000000} /* (0, 2, 21) {real, imag} */,
  {32'h3fa97851, 32'h00000000} /* (0, 2, 20) {real, imag} */,
  {32'hbfdd3a66, 32'h00000000} /* (0, 2, 19) {real, imag} */,
  {32'hc0f567f0, 32'h00000000} /* (0, 2, 18) {real, imag} */,
  {32'hbfac4333, 32'h00000000} /* (0, 2, 17) {real, imag} */,
  {32'h40174af6, 32'h00000000} /* (0, 2, 16) {real, imag} */,
  {32'hbd4f8330, 32'h00000000} /* (0, 2, 15) {real, imag} */,
  {32'h400e9e2e, 32'h00000000} /* (0, 2, 14) {real, imag} */,
  {32'h40a2eb9e, 32'h00000000} /* (0, 2, 13) {real, imag} */,
  {32'h400ec1a8, 32'h00000000} /* (0, 2, 12) {real, imag} */,
  {32'h3f41ce94, 32'h00000000} /* (0, 2, 11) {real, imag} */,
  {32'hc03d3dda, 32'h00000000} /* (0, 2, 10) {real, imag} */,
  {32'hbfdf26ae, 32'h00000000} /* (0, 2, 9) {real, imag} */,
  {32'hbfeef75c, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'hc0035403, 32'h00000000} /* (0, 2, 7) {real, imag} */,
  {32'hc01326f9, 32'h00000000} /* (0, 2, 6) {real, imag} */,
  {32'hbfb42b49, 32'h00000000} /* (0, 2, 5) {real, imag} */,
  {32'hbf988fe2, 32'h00000000} /* (0, 2, 4) {real, imag} */,
  {32'hbf714992, 32'h00000000} /* (0, 2, 3) {real, imag} */,
  {32'hbeb2d838, 32'h00000000} /* (0, 2, 2) {real, imag} */,
  {32'hc02c9964, 32'h00000000} /* (0, 2, 1) {real, imag} */,
  {32'h3f85a64d, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'h400afd6e, 32'h00000000} /* (0, 1, 31) {real, imag} */,
  {32'h402df90a, 32'h00000000} /* (0, 1, 30) {real, imag} */,
  {32'h3ecd0d44, 32'h00000000} /* (0, 1, 29) {real, imag} */,
  {32'h3ea96314, 32'h00000000} /* (0, 1, 28) {real, imag} */,
  {32'h3fcf26b8, 32'h00000000} /* (0, 1, 27) {real, imag} */,
  {32'hc080bef1, 32'h00000000} /* (0, 1, 26) {real, imag} */,
  {32'h3f6f4bf0, 32'h00000000} /* (0, 1, 25) {real, imag} */,
  {32'h40d1e54f, 32'h00000000} /* (0, 1, 24) {real, imag} */,
  {32'h3ec7221a, 32'h00000000} /* (0, 1, 23) {real, imag} */,
  {32'hbf8cb756, 32'h00000000} /* (0, 1, 22) {real, imag} */,
  {32'h3f99c908, 32'h00000000} /* (0, 1, 21) {real, imag} */,
  {32'h401bc9c6, 32'h00000000} /* (0, 1, 20) {real, imag} */,
  {32'h3ecd5580, 32'h00000000} /* (0, 1, 19) {real, imag} */,
  {32'hc06fdce8, 32'h00000000} /* (0, 1, 18) {real, imag} */,
  {32'h3e98a070, 32'h00000000} /* (0, 1, 17) {real, imag} */,
  {32'h4040fb17, 32'h00000000} /* (0, 1, 16) {real, imag} */,
  {32'h3f77c8c1, 32'h00000000} /* (0, 1, 15) {real, imag} */,
  {32'h401677b4, 32'h00000000} /* (0, 1, 14) {real, imag} */,
  {32'h3fa310b6, 32'h00000000} /* (0, 1, 13) {real, imag} */,
  {32'h3eb2445e, 32'h00000000} /* (0, 1, 12) {real, imag} */,
  {32'h3fb3de98, 32'h00000000} /* (0, 1, 11) {real, imag} */,
  {32'hc03faada, 32'h00000000} /* (0, 1, 10) {real, imag} */,
  {32'hbfda96a2, 32'h00000000} /* (0, 1, 9) {real, imag} */,
  {32'h3f1b8cc6, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'hbf813d94, 32'h00000000} /* (0, 1, 7) {real, imag} */,
  {32'hbf7dc5d4, 32'h00000000} /* (0, 1, 6) {real, imag} */,
  {32'hc0236260, 32'h00000000} /* (0, 1, 5) {real, imag} */,
  {32'hc09fd2f3, 32'h00000000} /* (0, 1, 4) {real, imag} */,
  {32'hc000956b, 32'h00000000} /* (0, 1, 3) {real, imag} */,
  {32'hbe6ddbf8, 32'h00000000} /* (0, 1, 2) {real, imag} */,
  {32'hbf8aa668, 32'h00000000} /* (0, 1, 1) {real, imag} */,
  {32'h3ddbaba8, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hbed7d248, 32'h00000000} /* (0, 0, 31) {real, imag} */,
  {32'h3ed371b7, 32'h00000000} /* (0, 0, 30) {real, imag} */,
  {32'hbfc394f0, 32'h00000000} /* (0, 0, 29) {real, imag} */,
  {32'hbeca5ae4, 32'h00000000} /* (0, 0, 28) {real, imag} */,
  {32'h3fcea8c6, 32'h00000000} /* (0, 0, 27) {real, imag} */,
  {32'hc06a3604, 32'h00000000} /* (0, 0, 26) {real, imag} */,
  {32'h3f0fb004, 32'h00000000} /* (0, 0, 25) {real, imag} */,
  {32'h402600d4, 32'h00000000} /* (0, 0, 24) {real, imag} */,
  {32'hbf10bef8, 32'h00000000} /* (0, 0, 23) {real, imag} */,
  {32'hbf3e1240, 32'h00000000} /* (0, 0, 22) {real, imag} */,
  {32'h3fb770ad, 32'h00000000} /* (0, 0, 21) {real, imag} */,
  {32'h3ebe42fd, 32'h00000000} /* (0, 0, 20) {real, imag} */,
  {32'h4020665a, 32'h00000000} /* (0, 0, 19) {real, imag} */,
  {32'h404b9767, 32'h00000000} /* (0, 0, 18) {real, imag} */,
  {32'h3fb1700d, 32'h00000000} /* (0, 0, 17) {real, imag} */,
  {32'h3f1ad83a, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'h3e42572a, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'hbf36a84c, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'hbfdcf965, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'hbf5149db, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'h3fb871ac, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'h3cd74d30, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'hbd85879c, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'h3e254cf8, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'hc0065116, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'h3f0131bc, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'hbde24dfa, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'hbf83f2b4, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'h3fb18025, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'hbf4a8514, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'hc07cddc0, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'hc01becd0, 32'h00000000} /* (0, 0, 0) {real, imag} */};
