-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ugJesKeIdzf8NPG2XWIhQHgwbvMwubZbbQVzozO3Gyx8cbtgt5gEKvem0a3dSP6U
6k5X4EKVf/pMSaL3Rh0GcarTX6JRv0TnEAEvzIC7vVre+5SdqHwhMGwkCDawzow1
0oHIrMhcGsAO0xQGOUlvP6/9cYonPGi9S6PpLu4tksw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 47984)
`protect data_block
IhsiViMw77Q/qdpDF/SUT9l9idQCPrXken6/V1Zn2pDFEUGGpMedFB8IWlsRp0LG
uHuweIxt4uUhNIFR+nIlBP8GJL9RDA8LAkuqXnLJYgYngt+VYXZXuun5FT0K5WzM
JDMMQBsyss7X19mkNE5OFmch8lSm4RFn2yvZlAxzrTDWoMPPXutZQx51oK8Qil6m
VgXT2SP3n+JFdWvv/B3N4SCSQCo55ll1BnVmOEl+ReQk9nE1Mi8MNKsOueydVoJz
s/lv4sJnr4NSynTPEM1oYtDq/q0f0jJBQEj/KtXE74sA6rvSULOIcUs4wn8/hPA/
CXT4MvuqiCvnADfmMYzVwTIq96MnzXzmOpVaAHI7/MeEkyMkfT/FEt8p0o13tYGo
cuRiKgLu1mfKax7E0Fjrntu8jpM1n6TBrhrjghr2CIM/yRdtixuKbrG0Jeaz1c1W
meSyySvzPebxzIMninv+BeN0KDf+wJkFTXBDgp+J2q9OD11xlcH4UY0TVmA9LtrE
IoKdz4W56W3IygFR5FN90++qZ52SX1Ignlvz3/kSD4DogmqkayLyAMS8fV1UNznr
1IfSwRz5wZGH85DaUnFyFhQ5DUAXhep2+uBKndKiU3Rgtx3qqU3S3DCjO3ibw7u6
8K/ehvR83/FjGbVzCNs5/rD3Zi+QMVP6PRwLibJ43JmJPvZQcQWsSv13IHMXX0Ze
vUVopkpRA6I8Y2eBbXle4fvooiTqXzmlDVzxSV+mjCXyuYZK2TPcm0O2uCNhIJEo
xWSTtTNyGJKBYtk6WlzEipLysQroU6cc/sho9oe6xTB2KZqHUut9YSMpn9i3sKLG
4Q666Xiu/awMPiPJ6iX0FVus895NulB/RV03sp9SNPP+8OqErVZA7N9kG7SfUL8b
eXEKg7Og+ivwaY15x0AQ2jrc1Mb+V5kWylSPkak17kUyEIZLvS1CHrVVFLFWusBR
pV7kRpyAlT9M20/uf/1pYEZk9WL1qbecPXKEwq4LeD3WXHXidav9ji9YEok2Ldov
u/SUz9SuVfWj0CQetmVlnkb5IJQunYI6SEQ4ReKZvCmYoalVkZnsoDCCqdyZx5J0
gLEWu+hiTSmWmDv/cT4fUnp75mcIdFzWburVkPNJycsdWWTTAv9eUtjENM5SE/D4
Ex1+Oh5Pnx11a/zlQHCWN7lkdX/2jhBXmFcaZgXUpUwMBxPuCrXZdtJMPie1gHtG
HRkp2aiLNN4jGdDaZqy/cnP98P+euUozcX7vB8x/xPJouYIq39ex1hNtAuw3mlK7
biu7OLiCAcmmXRTzCRnytQsqzkeuGQg6IhUsaADWJu03fyoLjbtHZ91tfYng4kcn
Y02WQv9XADueYaidORB5+yabBl1uhPka44hTE1no20YcH2rIP6iAeU+PyTt743fN
u8pLsSmAfCXKUAsWOnVkRbuBp48xsrCNGOB9hPuARvfkN+VZlQ9xiyAO31vXJ60K
8cXyzj6hJ8M9tbl6qTuK5S/09e2ErhLu5nQ9AFHZRPFZLMMpVh57RQvSTv0tibm4
kvpFgm27yQtCVl3NjNlSQozQCOOORBYRAi2xaoA6u9tzfjUt9oIEa7wghsRaLmjV
yZ0hHOvdkfgvR8nQKyjueuPybaUigvoLjMffufumMEpeK3k3s7WbVUnA/hpVDMo3
Pn7Rn6MK6yvK6mX8KpiOjP3kkVZO+sa0q7Kb6ptAyMyKp06FPdN7qjUORQBpm8YE
7M/Q8zL3URBbzvACOkqasVNKHb7VxH9OAsGCVdpVFJZ8y6AVdQ24vPbgRbEdCgs1
1Ng1VQiueDqX++dWsNAJ7RLOIfdiK2exM/0wTwJkBH6nRRQoqmhJu5C60pVoBjJ/
pZlQIj45lhEua1Wsb6NQ6b7aiehQSXSgK4qwDC/BrwlqldHRfqJDuHIsCD5yW+mw
4y1U4ojNQRyjfJeKHxdkYwQqPqMB5p3Np+bNekYy11zwfxT9nW8lVS1AVOMUh2bV
SAcGDKYhE4XWr6yAiAEKznRfRu75i/cE4E4lqSSdhXyTs0HUpl3elbB08r2C4xOx
xsg9rOoVa2RTwKxMCnmMXI4GvFCmK9m0Iin0XgoD0ZZ3fgG+mLN89y151Q2bA4DO
CqXupKzB54wvfLhcnShEZYCWK0Qet0hD4AzluifY2O4FnXSG0kFTOvShho+XkWvv
ckZ/OmxdL651pnLsdCTzZRWncnVDmbR34oGkgX5mjIo0JygtfbgRcVYmuFQNCgiP
hpfZloLtWTOJFWB7sawzIw+MKjrfbqm6TBvJNzeZGjTthezL9Os5gO94G8T7LnwM
ePM7fXjiBk/WY3fZ6Xq5hQj0Y6hNdO/WVCv0wqUH7/47SjrZdPXzibqZdoJglQCM
7VO9X28asd6XWTGiaQCk8FXHPit6yoeIUdpn0Mpt602ZxYUx1CawaG7G88IJiOyF
AhChQUpv3gGJxOtaFpaLqPTb9titkt/LmrtiL2Y16oJi+deTUmyDMnMvnyY/H7M2
6tMgFAzne5e0YzStQtp0fr1A+vBGVZaWU5D6/ROpdbd4nIdPDQMTKNcym6kwErM6
jE+lYLmLN3asGMjMWIgMiCZNDQNdi9rbET8H3JxyhHk6YhIzz1NpVjTlcbgPKICC
iyzi5KTdN72ph/ZP6sEjv9ua5yc7dMwbkE5aLoE21yZeX3K2ae2dscVDksNgLqTm
ThY5EfUQIh+c7TQQUrpjDnH3QqFUgDglpGQm01HCfy9yoO9w/kbwC9pdaNr3tgiM
/41Fk5A9A8RJu15HLMgZOxW7OpRl8LqxF2SfL91rbBzxSXKFYWlTq91fiC/JzZmw
RUQLz77P6IgUrgdUJAEKVYTDPeDWX5BC7DLjijDQBi4TOa+D+VrSwNhGnEYSHhF5
4TftNgZczIcJOyeJADYHfnK3hgKVmkdR6+D6o1SzospWem69yGl5iJ3T0mEl3VXn
0vCZnyw3mSQOHl6V0wI4dq/Vu6mvF2jSBQoag5kOtTylfA99T/5pSeMxyFq9jR9n
H07/J81lqGsRgpd6o+fprX13JaoZksDhwgc/3l3pD1lfOpAb3sVNaYVU5GJebCzs
Nhq/Q7pxti+9lPpqJ5alhgmzHJKXccNs1P2Wj7hAG00jKmbuEHq2JiHXRQZc/JLp
bzcIeVZiQ1X8rnCvcaKfHF+OsqlVRmSTizl3eFdzg5h8UTVmxX51bomS4kF9jEam
5qgM7+Vfs067JnMHlEfDQ34HNV8y2u/seYWxxh4+GUW8bjhCGpYylpxohpxRCKEx
ApFmgx5X3A3FvEF1X2MweZBVoU9IlTQzQkZvR42SDjEhQvTjNMityLfzda8tzWcS
0ae8kHq5fB6dfvSEz5byjNdpGMpnRfdBBqBvXOYuTlFMMG1jI3oGUZVT1qCLrL4C
duC5wNf4KQjbpPhg3L0a3vImSQmoS8pu+q5XOPJ8hl6FwweH1RsDb/gI2G1nHy/E
etaeRGEFNsildwtyjbERaT26rtuyMCxW3+Jbdfs0NcEkrOihpYOQ1EJScIjfe0Ma
e4h0c3uxMfqtCY65TJrWkjfG4H4dU/rCV/d+4yj8xv9IYfcw95Bpb+yd2QKUkWFW
lOXMQASMELhlE6j/PjiaBnRvQbIDu2CAZJmxSE9nvn4wWsD3EIu+BFDg6aPATEgw
k0XPwXxGKG70g2oFNgw4WggMlymdRHIHmU+fuwRVaMS1BRcVaZLNYtA9YMXhOMfY
wWJA2VSB6oO7s/x6vfA7ajNgJFfIXBjz5JHkMGL0vBFiW+3IDlOosfhHgD6zlWli
zSKWdCk5peXPw+EN6ZTqvABN1hKn7cWGQ6sGyRApQBxQvbyxweS2EVGjRFzcbCgp
lRwfliifSNUARU0pUv2RI89gMbKlDdRpXnR1HI1SqkwxvmmRdt5emhyAVktSgFYL
RJPGyfYeGLXqTcdKv7FX5kcPgtW0fkyu771Ps1KhiCas4reyyHWGy70iNOTgYceD
Qi/HveWIoM70aMvcCvevpJRaGCLJ7/AzN8MtcoabvhE7hPMhI60fIT7QIGhGSm68
hxpHBos9Ev+q/ARVHmUFOdwK2XLMIWHmUKT/2P+CFtPNtMUKQbluAW0EjduUVb29
YHGYG7RcyANOVUEsIojBVvneah+rRq7HTcD7D/wolID6jijjj/LE/dj89arZHtLu
7hp0t3xNJpucExwmwwOz+FmiT2Y5Lcof5v3g5t+7Wx2paUyQZIFMW2Rf5LNyv5eJ
PUpbeBeogOcDUEgzGZ4kbN1XEt6A1g12tQgOTc9HkJUTLN+wA/CL0OQelzEqZljG
QUCvgyMoBcJ29sbDoAT2WJRxYvfLI96qzax5e2MylW2qiJJft34oNyaqeeAXGTqh
aQQlW2pZ12Mu8s36K2RBJB9j9QoEJyTL0S9q9/1Ol+4ShvelK5+k3z0qCKwWE24J
FhZwDqRVadjO4ymtcUI9vT+7ToDtGYw4omylrg6B9EndBaQhPmmkkejFW3OFzdyo
MGYHDOV0TUwGvW0JIgkfIeg8aZA5910oUmFd626Zw5C+HmL+1Mb5mj8lWGrMD89y
fUcqAPWZ1yaYyl2PEiigB4kgF1F4z+gsX37PalngJxJkDZMJicSjpW/AazW4Gg0x
+Nft7hv5G1GHGVf7c8MwTWf4p4GYIJSXZg9rWRfGL6udAzYGfJUYpR5rU4g8+v9I
KoB7l/ffQvdYL0Iu6BCcvp2KHLBarlMy+DsFHeLuX4c3qpnm8z55IARqepS7UYHB
59yO7vUP+EbERU0No40q9wPpq3y1Cr796Boq60lOzXZRlrzmBhrA0W8qa/65BJVG
s5YnHVfyXnfR5dzXu0yU6izy8Rpe2lMYir4QPziieuxCwpRKB0jessEBB3ojvAte
sHic7zQ8bgGmmCmvL19ph+zzq5eGKve0cXIOxNKk/F5t0j1DUpa8T+CWvI5ohjE9
/ojkc2LyGke3EYqQDwB30kxXsfoDZhzGgzEYzL0tJnQJL0UljwN/SguGmv+aRzJy
n+S+QTydmwJoDJ2wZl+6PJ/vnesteB3m+/+tBMgTGaMmjmMZcnCXJWAK2oUpxboS
LltR9XFIYs+nYH6xxSpyojYcjfRpwKKmMyAfyUBgT0gyezuovFD9Bqa+cZbAftMe
cmhexiYB3S9aieRZ0yPJbDuFoXiHket+6JkK4mgOAH8KOAmkrXcm6339T9aLC+Lz
2lFxxjNJ/BR/xT4p+Yt1+IPGsKPJ8E/psFVkWM1FLnjo0hL0dDWDPdI+X1PuwM+4
dYPT3rBZAlWRWd7jWCpaHfelQAu+kNUIoV+0H8Li7krXqpx1wNBVeX0mXJOHKbG3
rbpdt9vw9ZsNYynAXTXD2Aor/KkeBoaNZojlQKPqEZRqzqRuf1/YnDVeMhA3+PPK
JMMozk3bL9woekfMStNjpMx/cZ2ETksBvlYneDlgHcsHjavR6ReKD9/iSghMU42L
EZ7WVxi/cUO9qQApLYi2lFmPN8AKZNJwMdFD6F3oWFCDhe+xCledXU+w6Hza0DiB
u4aa6Woy/OqbPZYJ7S5514A2Saf2dzEPXmLPNk/czQtgqPngG/0viYttZwUozJrj
dFwoHXEXIXwWGVwPTgkcX54BLBV0fKDjsc3CTiQ0CpYW7N/Ynw7ZYgj3JdmzhnYd
dGBybR2QyVn0yCoNJaOx62vTvwJEaWq25oM32SFtudtBxpYHTwSiTy5qTnFNHHH9
fFjBIn5dt5YebZg0Uqi1+0jeOouYJRZmiS+4wv1Jyv2P1YRSNGl6sVnzyhzgYM3U
yGU4W/jQNAYChuW4iVv8gREPfq51PfjjXKMqsfcva6xgkvEmvDEzZUySKPjN2JwE
8lDFK6kGYBtnimpX6KH8CeRJNPEPWwQbJvkJ2GUgYmqSUJfwUWzb/6h7uiivfP0j
by+enjyzXmasuj/RayZm9pGNp7Zk6tOqWuUvLKF0rMRWi1xsTfCPp8nJVI8VYqMw
tT+f/hOKJGzneA/u4RRInkMj2cSTkx6woh8gNYaJQNkFrZx/080C8oYd/6wyN+TP
u5Setn1lE4lw0NXuVsQ2Uw3GnsoolVrSgl4rGhTwN2p/tWu4oj7zAPsbBXrwmwA/
stzSwoYPjBHXDtyj4M7c2jo5Nxd5cnTF6SaOkNJJDm0Miy3CpX1LGvcKVJ3NiOC+
vqYrSByyaTe8IlHqk81AgWB3HpcD1TCI38iRbsc18y7rN4mn5+t5D068h+t6BnWf
GHlHvGqd8M2SveZutlYH0f2lmHbvgdaG+BEsodc88WMCxZN70n2EkO/UqXV/wbxx
37c/e9w6GUlxCBiCzhl8LsoZ7rnm8YjJ5aaozf9TQaHdsTD+2zCBYOA/9J4fNBW2
kWv8i4k1iWAQaa3oTHpdidm/WDs04eJEoAss50/YG0cvpC0hUlMLdhzt38AEdEY/
xKj5rpUU5rBktF+ozFP0tK5Ts3xS9+xrMqugEf4aGZcDNZ2ZEYjK3K2o+Z/Vz4wu
86oHQEuYSwjHu4IerRIlYkLinowvnPJU1J2EqgYhZ9v9Dw5TYdlK57tfkzaU8EWu
RQruJdNbp/6a8+oL6/RJF9I6Lknn1KncCdvJgD1B0yHwuWVeEaL0qK0WYWLE1R5U
hOO5MaHQIbdwrq7r2/0d4REin0BmPBY9ffwCv5meSMzyHjlOMhKbcQd5nmaX3RcS
JdcUcGqB+7yVYaKTGU4CB+ZkN0nwJsB5q9TTfRK1iGyTHFUE21DgbuMPwFHUFBtQ
xSBfndLFuZUillAC+8ryN4VaeploVLxp5LxOWHWiIZZw48HY4m/uSebqep0uUgmc
J38bMB9s5qryrqjCNVAv4ExxpYCczCuloTVOrL7d5L9xkdcVYRt49RC4Btq1yuwZ
GJFHUcWh0VZpH4/bo6au0ScD+MRJN2J+81Z/nr5du34qDsTPNru7rSbfdSrxdssF
RJZdm7PcTjhk6iO9HnFte/f2zXLnrBmTUiLszWQNfgyXWL+Ks4fwdq4TrE0F2Gs5
skZoDE2kAtvL0btvpIWAY2aIuzsn4wZQ0WoH/7otU8NmbKuSieU/3q/G3n2ZkzjX
qVmgfQfM5H+4E4wGsCtfzQ+/A0TVlrMRaS//Mrb5EkqC/jxqjGsrqY2vTxbNtDTN
ygtoRYueNxxxrxqBYi5VROqiUnDKLZmHQUCIqEgnH4gdBBWgWpksUvO6bSoSDYi6
5xQgaOiAepZcXsCGX1eP7UgVlVYDpiAmDRNo23YuqxuYhtDYRnlsSRGNftH/ouG2
YZn2j74JRTRfr6EQZnu/lCPnh9P9l2zxpTaTcRyui3j2RQzc7Dp5OWM/XUOVxo+B
/sN8p+Q//z9Sap7LsMFZCn3ND/C5Yh8JsbJLRyjn4umYIRy0kIFQFSOd2d0lIkSK
OFWdRn9CNZxOLEkKF0qIG102q9Q+nmHvFFd5wXhT9c66pzK0vYel6QjX4g6Fppno
Wul1H4wuv0SPuBzhX5bMs8HCLcNOqr80eVYUfDRbwBKa+NOSuDUA0ajR6l3wA97T
sl9HbjCL6J2iVwcHvH5s2bGPO/lovjarQeO7ZZ5awHUjcnFeiNFqB9rUz5JRwo/5
yrzHv52GCLYh6CKoAjhonOxkSCSQUgbv48omIcz9CG9jVyQ4zGljOPkpcxAQOEt1
NGeC0g4xUp36lQE+enG3R3tNcgO9X8yq1SJJlCfz1Tnrs+WS31zkLHeRmm2arQSy
jav1trNCKNJ58U9dVSL8kJn6ZgyrX9V5Y6vbYYHsfMOcz7A2QTucNMfmEe6m91Q7
sOGkDiOYX7Cy0s7N+el0Jd3gFcU7cVBDxJQU5ehUaq/amdre/YzA+Ef5tWfvv+KL
Qf3eaZXikNxGutG5fPXxh1KN+t2v1vTcJSMKGNNHrE9wcizrpnTqa/2Igp3WnvmM
H7/PZ9SayKuS9y31QoGjCiJZzbIpbzelGSRR17PKuTceS4x1mJG9yNP1Lx+B0azX
tluRGCT+axJAgxEa6mu1rLA+04pe5H5YYsN4VKYnLgbBK607zhwm8MdXsk2SZr8n
QsCyvaeowIXKqqefE3Iaqw4bwcGWYt6/Ex7L3f0OheYTeIUqNfFeOoDwkOa+0FgS
lKuYCsD923wwt8b/5z/8XdN80pLp9mrJbf2ySaC+NJSsW19Js8MVKk9Px3uD3OV4
fCjYKkOLxC/qLHOUM6p+ROx6j51iqPPDDdjLUizL+83gietsvn+w59mVr4cK7GB8
afoErUY6k5XUK+yom0nWAVYaPNQhuS+xd/OOBxY2m4MF7VSbYO5TMAkhMKUdpdlG
5xC7iPjIj4xvo6GiGF1B8yDVGS2KSL5GTZL4mvpB4UQKfc4YVL5qHj4FP0O0tdmj
a0t7WgjkfkNWk8EmpasJ7rUu/2mnqE9BZK8J+5g/uN1j6Sw+Bzr02oOBskTiNMsK
yyHclhUwtaJeT9pPicOOVX2wVCuoIr9i893Iq14ArgMQfMhk2kg2FwHPolBYmO70
wL57HYdcdV72LwCnGUfwKNX0fhUdYtC6rUCUoeUxAbDY8kpx/FCa66H6mAYRlxs7
xKGGi2BI35XwsLDyNNclEaEQP+ivqc3JFCHby3RELUkTGAq2RUI6a4subObbWxlk
sk3AngP9CFLUDanO5WH/+eK8vW0GMF9lrw1o9VXacBTIghX4qan/jYgQpiTr1Khk
1vgXUW6r3pNp9CJ17uSx1VurasSZ0kjo1qREBJmvLb9vB0OqbCIFFd9ASBtPKwaz
xS1f9NhS8dE+WUFJaNEYeMYvZbMoRIo3WzYDmlCAFJlENv1yEcaevEoO+2NeAmPb
/h5uMAJLjGYfn3M4ZncCXDUSUnMm336Ag1cRiwAKO0Dmi9N6b+3SIedxvFG38GSs
u0OvlwTn5bszObHGSHinWI5wCZLquZbmP8h4gSUYcR0S1uU5fmWVYSFpzMpuMyAO
x+0H84WxDl2fNFytGJemZnR4I9XbD3kUyymxCwVHZlmrPo40WaM/qmDq8VV6Vari
naMUVwKtporEtDVub1I2P6fp1VxOs3mnQXwa7GsOYwXqyWgpupaLm/DX2dJYUU8D
M/hnYCbLbSk+Hbe6wktGxC73Nwvo93LZUfjHhGrdItZx1HBPv59aDYi1NL1wp2Ko
HbVnri5mGo86/PRW9mxIyteXomYQ9cAJ05867nbV4LX4hkAdnnnIqdbJbeHVOcDc
p3hq66AIBQeQ+D4juM9jHK2tmSpDIN4FopCkk3L9Kfc7VJhcx3I/N8mc5Jeya/QB
pnYDYQ35gmSno3vsZPWIZmI0McIqK6DSDJWBkSrc5i7L6El1H51MubQ90MK2ABwK
nf0UncmAp8+X6pX1xbVbuzF9/vN5sqnws5sEg/EoItGZwYja0B/RX1aWkQ67GKfQ
4NV86W8AlICOkQns5pV3mldaChScdBo0E2TTf57maPwLsxx+PfRkujD1Ev8ia3Kj
22p0Gv5W+YhpBU3rP145OSb1dmL2ubcX9Usk7kvhMTcxGaBbrXMRw2Ky2+uKrIW7
BfXk3SWbS+4ty07KVtc5P8C0nqDn5/R7CfN4OHkmNglSxyRUOwL6c2rDuj6YucJE
dY85AT3BlLobSJ7/NlInqKVD5n97QbaJ7VCuakQbTAjeT90vhAS/kwWPC+LOQMzl
1VIok5+mZ1jB37gCcLtok3slWi26joOh/GTxZJyf4+p+MDe/OVPZeLQgex880nTz
HQ1OIAPRxPRhi5im+W6jUv8ZYnpUA6fpC7Zi9OgLTFoznakAsttkVF5Rm8GxwCKb
Xztrfpi/WEfg+ABrYRhhj3yN5TpyjJHixFfhEtEWgq8djKg1JNR9ojXLgeisMR4a
bwNnZr01VkamjxjYpeKJbi5RfE/60TXqWegH39pnrFg+5nMJWl/2wFuuioHBxptk
YdFa1hSrLroHaMKKVSicTajnBQe79g+V+fJSGiYjoDaz5CIs42ryAqHLve6v52mb
ZzPQZqZ0PSStpn5AmgekB6ng+gSOmplJAls7Wzjvi2pWnmiLOZDr0Rc3exT98Jtu
RRM6g9LOmG+m/4d0lYYg/24WomSitz3z4HMTf4mXLEGS99Ye6G1VVHhYLogncNLn
F8esnYmcQNRsQ47+Ze4hqbKX7HRs7QNlbE+4sqOZKrbH7uoXZWGmGSZ4ePSujVuY
EiW30DkYbq72P03sZdqGzp+FfU68mfWHvxAdcDhirhK+Qt6l3DWmd2iCTOF40/DB
dN2hINpSUwWWGCpjnjaRHxggQfAunZHnp7MueCvBOlaCSuHfE/XJKrZQ36YYWUlM
EF7rYkk0VekE4YA7pqH0xseBKDDtRBGK0WuEQO8Eane8knCzKOVLO+9KWZhUVEpK
pHqVU9OJ6oHfkyU3QUKynzOgX891vFbLhxYGLTcq/DO+9p9Dc6PP6jF5esRU3puT
pGVlPTERa67guEVnP9Unp0V6CFNNCLH2psLO0YexHUOwkhOWuXhZyL7tSzfftsGA
Pmu8DNBKDFHrRlyA+lns6S2rpG4rh0nFjmzMzFRtuCHXdC1fSM8qq8N4oyBA2Sz/
d89i/rkCxsy0NZMlI0+tHvbiDuTlq8rL90hWNsmcnSvrVaB+K2AGzoXx/Z0w3nBr
2AkaCoQ5H8sK6Y07DpZ1VFvCmvwgLHyxER+eI8uMhPgGyoizgXQT0LrhNcHPSjHY
iWCzAPzFEos9cGABmYWsE7CyxFUwi6W5TEwKO46NtxBxjAY2UlvUCVlQCDpu3q3w
liuRczuOARY5e1SYeW/kUdQnVLBXOe2a7JjSfMRYQY0He+ZfOUsEFmyhnD2OYmvu
xvU6cVhUV/zRpUj0NYvBOsieInrXOdGvKRGDTLYqLOcAQpup2FCwAYYz4CLx7y1z
VvEO2UtvTsjctYtlrDn2Mm0r9Ekj0OEgQKIvw73x8HAoYiP6mlBTE7Wyn1rULYxI
VNAfGs5cvFBXlHSYfw9TVSfeJpc4qra5Y+jmVQvz5CTHKqBj5cXvbcT1no+x3k6P
2BCHWeBYfbaNGhm9Uea19ZHuytnmjT79jJCX0clghIa0Oz5JtubpisNJXHJm6Xvb
sD23hPPjLothHfe4usCa6xVbGM+TZd9oxuVxzY+G+hd9JRagkicFNaljjl6Z3OpZ
ilnLlMicwYHj8aXzRPbAljFDKP8zijPTOKj04rTU7DqIjpBqH/iF8ahMkFDxKei/
NQykirrlnMsvAi0t+Ax6mpl9OiRK9UvgDKiU5fWkJDEJlnr5s9yzN+1ElVwrOasK
7k/6x/WAIrJIn5BeodtCWkNQoSTVK3QiSIWkXp4JUdQWdWlnEszDeD6/A35LoCcw
RH3s47FgDmnMgUeB4GJwFwA6cHuaPgXkIkBtj8a0oe5ZCy59isCaBkbtC7F3VNxv
XZeqhpdsQfC33R+CFydbommY3h8Ojn66+TIVKGVqMIdiLr6zEFlJyGreAmer42Ze
dHRllQeQlhpTk3ngjoesxXjhSV+XQhbuv3yL9QyB0kHUgvw39/2lLw1/CvEmwHFV
fOjEFhEMub2JJApJNrU/45ZjMACR/cR9jwOA/PIqyzoGMsouHkIV2JepIF/Lzoar
KcRxdE34ma4DU5HMqTuEg47hICtGZFdaDX+oBYJLZ0o+yCRbUbPKu/dRb2Cjhbm4
Nvaw6xDoZmeWvb1zE1USQ15QUZDej7S+zX305FOgquBEm/z7zWeBAQAbv/StJqEw
5EX1cnTk68A/pxF1FQ2HVOv7M1ReFM+s2gBeGCam9+YiDsRGcI9tnyzCjCm3V8Jr
ZN/VpBS0OUrn8bYXvar8XW4a2vkNUQpouJFJj8m7HeOVt63ffbIMEPXcWmXuXUqe
TkKxvi43HjPq3dRFyxX0hsPRskQU3V0aQZWll0ANmeYdi03KyAYgt+ls7ykWUX5l
ZkcFVDIGSNg7qCQmfGJ6pKLa3rJoovEcmP5ykA/V3y0s1lu7HUqLrQjv9jYXxoG8
w2iY7Qqv7ZogRDCdeiyqA3R3+bSuu/UeWEtZVfipPoTgNFSFJeOGdhasp68WlH3p
FPcuEFauTs36Ltn6LxyAXZAG/6yprtV8O988oRZBdShoMpAYi5CAJzbeqpJshSKD
5pBmivtS1Wzrl+BilpIkp+SF4TCHUPa0RV0YJUFmHN/aefXnkdjJwua2sT020Anh
Ox2k4otpM55h3s/FsAXi+Tp75Xlc0T/ufb54Ezt66MVS1E8omxOrTO0fKkmtVCNk
9RcyG5JL+AR+NIySenTKJgev0KOOD8er2ySN8ZHkHAaRAHfYzbOKUIV+2WS/LN9b
6HeD8EPC4ZV5vspHcN6CUvN0nDU6LeiDXpD+5muFuqiBh5Y/4wC6QGI9hADa/nQH
vQ+xIbU1kV8KcPVWOAKxUqkMNt21mVqmMzKUIANYwOP/S8nj/1kasoVD12Cod///
SUc9W6BX4my+nysLf5q7pF68J7Wsc3nClSJZPV2Y6cbXCEPijoOnPrFnx3/GTZq7
81YQNsmDysbL1+KSYEqt+jmV1qfamJspNNaLC9WNvrwPnIPZcsF+Qlo6sAacKgMC
dCILt5sbblQc++1W6iOxxgouGnQmmrP3BWs0zCUUXhrtKIibfQHcyVOEH+SwFP6Y
ORMCYH+Uy+NrWNpDZfgGLb/x5f9XVqrQ9Pai/KFUxr0+7hqAndAdyxNaJ5N1M61y
ynlgPeyE1vjRIOc4ffcQSG8fYPIdD12KE56FMKKJ3YJ1D2rf8ubUhHeeDHo9K6qC
H+pX0x1fmwyCJmFoFncshcITGlUcDIlse4jAS899gDOBzu3AP6jvQV4RihBHT0Da
AoCo7mlRaDob7f/7xMSvxep1m6Hmd6aKEOhzazmBeoYcCRVO6AeSqZz7986uG7/H
x26TKZxHMhmlnTqJcIA1l6G2dlZ7qruCBrnIv1Ds4/igeRnWuWpVf635PfNZJOYA
VaiIiQLtMuiqjnfRnoPcqWjR5R5a/Ci+LOXkV9VFiQpFGaScufy/oh6Nfli1VVcc
9HjKMFJ02qNOzr/s4yusQeZHZmx+ATYjjIOpqeIAkBxTq+RWkUrcWa/UOMKOMocX
L15V3UpBKYdtDvqD/+/NvW4DCwrZIJHxSWjNv4u60v8c8wpEsp6sXqHQnDkxhyoo
u/64oeT+d6azcA37y0SkQTVRGZ9JLAB7ENgIpJYhWzWdf5My5AT6uwNAYMLrWFrl
6AOlVUQ4ZfvnbtfxFuhdHLomSC4+IF6dIqzzH/lQqj+u4IpwH3Qtb6u2DawPjl07
Vm+Ckyh6GBSfbGAVxjVeVY6CCTlmGpEi0o2A6AZQLmTMOAaGqzbfUEyKy9uemzON
aAx3sSKKAyTOC450ghQwduwyN2FnM7f5XHXjvdrzL+Q/3IuZHZJi/jC9yO2EV5iH
u4HEuX48SU0N/0xVhqbWUrcOJHN56RsbrSLZ6TbqbHrGIUbOkLoii2cphLE2WKqH
GQTW4I+B3A6iYi+IKVf6mU1k3wYK+gBENs2Bie7L3YMmV2pDO9sZflXrQJmad2+N
BPPXmUa6lX+vF0QYvVTLcSt8609bB+wo3MJqrSWhv1igJ/oqRZ7jQwBx0WpMaQK/
NiTFZGrrXf/aROJy0DQFS+2gBDhswLlwD1K9XpVRJoXbMjRnCozJx1wIwXgegHfQ
emczBkLmyCxcHfytlKf/wm7+3t7IN3Tobifuf7XmphDD6ooS1WeMj0kmhuGNPsx7
28Nj2uwRcXWnjIpTdGDi0XMyEq6Yx0Y+1Km/3Qnqa8AfHmu09h0tRvs/oW/QExa0
SKl1W16KFbN1E9j5+PPElcw9uejNAUP6Rr0W9+xsC/xee0QJEqamqo0D6mOpirlQ
ncApcQXoTxcfgPeQE1HKJ7HtKPRkYOLtRB/i8MsrVNPHa7QGCTJEfpkenh65M1lE
EHdJOwFtFipJYP6MmEkS/FVf7DltHpRYDsnoeBQ5AwshYmE23iXAFlpbBB1LPE2I
ootUE1Yd7SqRn71raDdwkv22KcbOISRZ69wVkWbi1MUN2cZTGtI5wRLOSuGBfqQu
APMhKPUH8CAy9jc9t+ZQPX73pT3VHUyEGP1Wk4N3N+nKq46WOl/+EtcAnX9LEhGX
pa24vJ3284mVkmLlNXDHruMY/ZKk80cS3wOR13BcvtX8z8/o34t3bMh3nrTIhnCY
RKjO3eYGbB7r+XOaPGFBmoz6KxMWl584lg7roJj5vSTTxAywnn2E1ASLl1aLcaq5
XQpmR1FAhiIa9FNpxWudCQJeBFkkh2O526Bm8cnGaA2srE9pjb079QHCBA1Vbknp
TW+jKmBDQn089jK3ElRuwMEfJgFzW9CcE2gjXARs4e71fJn1J70ACeZyP9NFxYWN
FUvkoExA6cAJvxcxSNixdMgVdWb2Upubb7PjoqAClYp/yfeq9A3fldkZE7gPbFiU
KW20d7jJgA0zFZTfZiMDe6b6SLTgnoHCeCWsdHAyog0xvqftx+vOqFdosGqA3Eqx
ZUG/wDwR2VOPSYeQtWjDt1QuU7ffqRzqVIhC477eqUJZfZr01dMKPIRRiDjJTqtP
YBzcDJKN6MuJoI0/vGmgcuWOP4ndzsGp3WZF8VslF2vdedCA5UySyMDejXwvfIWb
+O8GZtUaj5Z7exIkYzo9hxdP96viepHVmcgOgpdf0p5NQMUdwRi8JASaVDZfg/aa
bondfenAwVo3aCagiUj5DP/eul9umEkVPChtyhN24o9OSRaelaDzKzylKMtpLgqQ
wuIGJbs36i71akoFiUQ3UZBIt0j3GW1o2ybYSNGnHXfHUyAcbKyKrCGkzOJ2ZBTs
r8YSa8m8QJ7p2Fuo47aslSkomHz8U/LOvfCqKxoWefpTckhefe0d96FmqoXEwRXi
f+E+em6FU2d+pDB7M6+DETMvptIoYQ6+w7McUex9hEPYzytPvoFdBZMa/Q9JCmiJ
XdxVwyPbg8O6rimcfSLZ578Ba02JJEQzNdbNvOPzlrZ+YweP5lJ+otMrTyAbxcDy
p6NJOzR0Xz+qxDYAoKBGdyBCmW0vZ4ZeIGun4Lv6Bld7YWGlBtgVZURGRJYvwSNP
LUpjjFT6J7IcAqIINXXoHQeCAQCidOPYPgVl5Lj9NTbRkY1gmyZMwFCeVX3dlUqw
2U6+3kXkN8C2OgzPuDuLP3ngG0Rc8lZurSJDogsiFKhBv9Vdm7ihuQwfMHUaOm/v
mwJiKj5aNmt8r5WLmDlfheFuQmhCDgc3KvCPtFXLPTcIEYNr128wnnx3H0ckQEDv
KzdiyLavul3yGX+RlFouDYnp/4oRsvGQeNkjgg3zhLlIP3I40Jq8l9tsRYAY1HeU
a5ygGxc8cjx5M49yFNx5tJYnaCh4KienFs0amZXxtlVDeBAO2EjUehq9hnmoa3HK
cbtAMvyVdY7OtoCyaRkniKj0TucFrASUgErFCOQ3g9aKTGoV3GTYe9w7BEPRk1lL
piMfUUdzkbdB76xqTauJdu3kAvn50lV6TRboSHNEkuCf0T4QpkT8dl56UQnS9BIR
Aztn56yPkJ3/OfHZLxX29gTZAxzlRtb6A7nL1drKLCsTQRX08bS1QtKl2zui3OH9
xeYWWo5gNzKQkq9dll6LVt0ld46mztdZp0gWnsyNHzI7SSIIDoL6G2hM6f5ciJS2
RSdhEmXl/aAjqjG/Nk993FT/LkNIC4nysze/f2NX0jekhJ+1mFeo7zEqBlHfbSDj
Z6Po1iNCh1HCLNh0DgLwWpK0KHYFh9rDsCMLAoXjLhRhW2//7pZ2YWLWTbmxkDSm
Vv3eCS0+WgxsRWQwTAv5tU1MxxHumhXhjmh4/KlxD7oycLiGblcCSHUad2jsMHly
0qWU2QTARsnC1g1BJqOKSDKimDZfxwelaYaH5mvGERvISdpf0wggvKppcwUqtHiu
Rfdn8U5NZq6kGCrcn8LPzIwqNEeFkisXqXaIgZqtwJb9JDNhxTeFD/+IAYYrTGu9
wHTQd8KLh4K4OJEE26f395Png+zkhO0ST4oHH3snz+XrDb+fEVSmRH+MwQLAgL3K
wfjxnbAohGmj0jaZxRfcnSzNbNoLOTTI2LbVP5WOq9ZRFigyEcxj0PppCGhubwxE
Z/jdem/bTdX/Z1UIb0PQ0l1YZZRKo95ykv48Un56cNuJdrLHdg8AGe4gAd4lchyo
WkjBuYw1wX+muaZRD+rpT7Ijb9E/PsMutEEOgvObJzcCqKGTbWWyI4oSOJLc++4d
pYwC4iVRHtsoK4y8OfI2f7eFy0Fq8HdlcGlH/CGUGSMBcyRbniNx5GyKqrN14UN+
cwXeTyB5ySypMnT9iESVUrL23fBMz+GyUC7orD0c1kVtU77opE0WbnNfDErsIsNc
ePN18Y3ODtoSrHoSqs+hzdYxZGEvoS9YX+a6GmANuzFP+vyb7/2ABLfeqZrW0rhe
uVumWq+diSxcTnFIIDq+Z3FLNl+TeDLWWmEyYWUNXF8x4lfph8e6v+FUSwPZMeV+
zlXflvA3KbdkVM9vp2TQkjHcGhvmEGMsIZhD08dzIk8AJLn7WQ1td4ko0IrygT+H
/BvLv9ymMDWKWToVAJuFxRuj6Qg+SjnRvJJu8HRE8kCXYwiXGcobYlXMVok1Prea
VoglEzU2S7xnHl6laO9KTkGa0+MupiiyrjSUdPW+FNJtgqVUr1eZXRQC8YoNB2T9
77OJPl3VAghGEqTd+hS38/gjRRt6WQ8dciPS5SL50jrnxHsiT2XBoJK5Id5z8Hl5
aTyvIIMBDrGvWo7DzMw40Onhu6uj/iYSE/FYFMdUr8QS0ONhpnRatuD1tUlIhLlS
eNZjiFA0IfDb3SSpUi8ewI8FFQduyC5w4m8GMcM+/ecwO3hExDJPHI4QH6vN8LLT
cGepdFzihYSGpz4hTmzuy8f4BpF+VPyuT/LStpfNOFeW4G2RIZ7hh5UlOBZ9Ol9N
Oqp2oxpO0y9CCeeMlopPc693gYul/HEO6Ud1ecFa+XUQ2rxiGNmqNTZWAzuARWlk
oGi34orhKD9APAW8lbNVQss50Bu5IH92TBzG9BuU4ZkDK/2c0zGXwhxxBPnqSCh2
Ov+EdTe4LORLWOsEgkh/tNNuxLAzI8kNHZFkWjFut5mtvFJ+Jy57SReeyY9eaC4m
4OAYd7UB+sygUWZVRU010p4TxPn0fMAGo5o8SVpPkVzUI/MB6CVPpvEK7DVOT9hD
P2JJqv5LA6S/YBmVmQSgR3Mj2e8D2J8yQBi9nAgqe8w1QYBql9KnHsT4d5ianA/7
L/8xnmAgpBT9TtR1ZojgrTs0tK6UKrppIXzMlTDz4d9nPesTSjGtlyh6H598JTIR
tpp9QjywcIBk/3MBpte2fbXwTluj03YKt5hNFQ80daxolyAkMqEwpyQ8lTsnr7Hn
cYG/P7WI29AmQ7DNvw9XSRfHUMhzRrN5MQVk+7w4BKf2UB0n+cmcnkgxCjFZyhjN
IR+k0PlkXMwMCLY1AUzlrbRrigmlhRqUO6W4V6m6AAiYkhwzQrXhhM5daZJNSJbH
ASHzK5CRcNZg7+RzQDyxLc3M6nl5AH6yeTt0OPNPpOKoViWEZ7PlT9kzDwXNHJIa
sVQtVbMGOmOPiuj4nQmg2D6YIuwDkD48WYAUOBf4WlsObwa9sW1hnXrsVU9aRuPh
T7nSM4GmFZSsPSk8o8zi6FUSSLokYgQPhNWzK26H0YDdGmH2oiH1oeRPICK/ryyY
l/3oOEU0BofPZGWNSZcqWf2+wPuZ4/1c3+pjyYUAw0ElhLCRoUlqEQNyI8/zflu4
vrfK12n8NmItl9XEKdQl9Q4YC5NMx0Z7P+l7dc7/BVAczaubU8Qq2tMdaG3uWMUC
Yx9JGIZctGtHntXuykhNPyfJS9G+Ilyup9Bv5PdOwuFsKMspGhJgAPePJlZAS1Mb
cutIK5rPN8Pruk3EJ7G5eXq6AULXREMd0SZAf1ON8cW/H6Ts5quwLT5bIrGJZ1RY
Tv81+ZRW9zr0ICMLj+eratn6GzOQqJ1vHw9HsFu0q5m6NfPdC3YTgoghqTxrJZMs
L1+RKjrK0jn4DkeVx41miTzbPisI70iBgAoR0pFpKrMkANN6KXBnVcDgkQPjPYwo
8jM9PSUwKip1vKuYEsNrBYDGNoErCpWuG9WSylXi5itYXAaXiy3eiK7WP5my+wI9
5hVIq//Wp0ketiLEJ78en7F61gx9t+C31zS50+b04RgC6QVXyfRz2NIZ0Poux10f
0RhhfvDvYATsPwUG4AummDlfz4Nw/6rczCi0UpDh55zMxiif7jEFR+YWosjMG6g2
AT9NNLaPS41JvlVrgISqkAOK3SBgoKPicy4GtGZYRZYs1rmlQtWxoBWT8S8H5SIa
4i/ABYShb6isevf+KbEE3vVLOOnnrv17Qj1bBo9ZdSv0EqOc4jAtSlWEw28qQyKM
V30Ae44QFw6WvdYZT7RVgwprOejB49nBKPRx3X1Cf2RcNk0ZMwBIngPpfeUt0Pmg
LSLemwKhmCgnGVsSgPMlI+whPzwyzu3SsmqEZLvSenYb8xMc9gZAJbS+Xt/bKTxq
QNFVT8FZdAKXB/D+cBNKGPsQteax4gckFK7DhFKOxhj34ASPjNQMyqqks8vousnu
fbHVZ6TPqf6PifHe5YNFb93Mp6Qp7fZr9HR0Q6CMkAOiT2KlgWtQAwwgXERgXAVI
xa9bToFmv1CzYHnNc1MF785XREH6OPaM0Zgqv4vQzS1dSS0oDcGhF7xHzZmUVqUm
B0JEzP8G0V1RMRbFbAwGiJvATMjT2NR5ZqjwA2Lrr4dvzTKGzBGjrzhRBMeSvXga
pwkKFdp92+9sipdJ2ZxrOE+xDndu/M0o0P+2TaDcnpe/46g+Ho6pBPe7QUhTaPGy
GwQ2WJr08u9Uk913Vcsa/DyWLuGnGDklNeF1qzyEcMzj1BHW0wTMnzdmuMryfBAz
7tYRow9a1c2NoNzOVwvtDjelYe47xKmq7Q4PWWvX4KQMnO6a7/Fn2Pm3ivIRUM2u
CSCY/ivbcsoj4NtiBKJywcMuUdAxrqOLCZlzOxCmJWKViI6PDimYIqaSUEyyQJ4w
uGl2l/w5QPwHyZXEX/PhPVvd4iYGijRfyaCacxA2aQPZUVWYWCL154E/IohbNFtY
2ZVM7Pc9iIRghsZWxoCnNWwCM8MXFY5wD3KafmhZS3AdupSx58KOUEoZWtqBtUgM
CNw/WQ+YbblbC3/ohf38GmjJ9F2C1p6UUp/I/MRtXr7OgZbtwlBFw+C0XayhO73s
noJA+GeirTnhC9BXMFV67F7iTO3c9j+cXOHc7cTcCQJ+ll6ePu0Y3aNz4+k52+nm
Ee4ms0k9aoJ7Rn8CtYWkdkbEvIsCUh7NpvnKGxzteBjQe/ok+Vw7yWcaHw0FzF5j
VF/Bq6Sw1L4RWupHRn7BV4V63N2Td5i/7he7t+NORmc5XrHvX0JOxVCAssI7EB+5
rGk3xssSe2sXfDosuS7dlsC4limgcGKNY6z6Yvg7rcQJMhWxZ0K9Xq6j4kgWa/oT
uIwu7WhOCLS8w4LUUEVULaM8g6ZHn9krePebEJBwCfcw57fCmvGvxyt8sRHiiEPW
9zm11KvJl1/Z1sKTzHKXJjRbfGnZhxmili8DVUS14wLs8K0stwC+SWHMvzJaXwk6
lS19XlOem1KTmIfvOSJBToEpt6M2jrx7t0EpX4UQzV5HbWL+ZJFOKAVKq9N0N6AQ
kByCvGlQiGStiBhViMZiIHIY7/PTLHhC3j6ZascQZDPqwuNrpo5AgvEhkS9R3/FO
JDsJrEEUfwprX4uxTsCXYqUQV+XwWGhJzXswBcVlxks0oDiGYBsbCAQ+WB/Y3JYE
fTAGo85S8dRw4ZDEaSLk3wrhr5OCb/P5rTgXmnCdq9V3Nz5zR7Hm875+4tFsHPUA
PI5CBs2AoUpuTVli6pcccH3jjWAmByfWdOXG3uhVblKDsHCelCardkOCS1SBpkAU
QyNLvlDiSRlJ189u2mvEU6uFI6h5liW1AbDsvlxaJjzkq8DQ9f6rXbvK0t6jz9l0
KYNMa4+31yRS8cOEM3qheaEFDH+0M95UivwCYJwEoxjuErAo2z1/1LN7U1v8VGCt
WFB1H2Ot56cGc853ufAnSiY9c9ClQiITf3/5b3/RIIeE/EXKwL5zlukrXMON1Z7n
rHcVmUOqp1k1SUTJZ2z4u4AYf5HYRm0ZMk2iHi0IArSo9cW3RDzoJ4YlDR4baArZ
NDStZKgPR1R2NqzvBorMNUXDxJ6j5az5R2XVY0I6fN/G76MAszsC2qYH6/iatB4w
VpVJfDNi7P39SwTFAK4wr+OWqi5bZEPUTGRTIWrT4WAC25QTJVRiWtVV3bisRsg8
oZVD7KExdmN7CDXfmKHevQ7tT3+ujQ0rD/qQHidzLpHMujccD2q763ke8FwfCqYf
4ZJGO1xUdgAgsZPHk8X5fhkEbyLNPpq5FX2ISBYeptqDGxAYCqV1V06tKqq8dSfk
MqnLU9uBOvlpz9gZZ8Q4JBpUEWLGmO+Zl9nTfI9n/qAhu+rNGmxyz3u+lM64mXiN
4O/4AuWvO3pA23OTA1JEhxjbr4VvezvYIsNlDk9/LVgabWPV+as57Eh3QEX6cqBG
GE+2mv7DplMxRjd55iKYupfdJaVae1qE8HnNgPZG+rosMpn2dAdtcZ+SYSbmp6tG
LFJVjtGSlVVF9/UrAsQloIOtGduYkprz3qlhPlCtWk4/thg3V4K0yRRd65ZRBZIo
sc/Dvm3DPoR22IOcypJqwT2/oX7t0VbQRIuIS6lXkKbZKj6Knueoq2SxzxWDVoXD
q8EWu8HKSJmEKtO9mM4DA91ftBCats/q1y+ZEuQ2pWTsv8boI9ylL3XjjVz7adnt
a9X4Ozh9rdzJ7UgYsf+VgxcKXVE/WvIq/cbSpRI4Vtq97/DrYoBY2G3D1QRndJWL
lZeW4VMEGN+iN3xqwwb5Ek4vVED+6lXEvZd+QmD3XIMq9LX0pffKwBHH3GuCzNCp
MqefX8b1hUSGi+6g+9r8QpGGOqyQNxYAAKLrTu486iUxzPaAE/SnpPBmnWOr/KPK
w+UE1arFOX1PUW4qGfd6xJR37izWLYY+nYBTGTMsd+6snjcwMl+pmov1tXMzGMoJ
ZQGB65215LqykICZw3ft4MxVAKqY2TOppYt8lrYe8zUToYnXMDYyr09vxNriHMTK
Wyu+z77q2tI/qc9a6VMdP0PMRAivEyKZgU4mDWJsyN5PkytuzPXcaWVzWDqZd7PA
IV9zJjvLaLii7FkItVn9RkBfQ1Qoh2rcliG68iMJUQVzmDNCuWw4mO7PBm4j7Lec
jQG/GPw1IraMu3ANyStma/2aothQUufL0Lu8vI4LqY0PodbBOZD54OeyLIUBOyMx
sQlMXyR93lgpAzBTmEnj4l6u1Qv0o+H5joshW4VRyBhiOfmWbSZls52rYMWr5PFz
8VR2ZDR/Idq28tYEbeWpdigbtJ6SIBamv3VLFKHO/ghPS3vxhiYMZmjv3T228iIq
Ws3KiS99Z/SBQlJxsMcqV8p1+b18Ul5PGeXZYL1KobAtKmk8YIWo3LIG/ox++SAL
LfWjmRwOoRFXQWuG7b1QIXhMf3QFQEe4FSZHXU5TbBoQuXh9wuzl+XTBmHgJ6qnn
vwI5XDk1GVuluOBPXEKSBtiSne49kKpE/xO5nWv7Mk1cwGu161ywOv97nxauxEry
IchuYGeYzcj6X7oU2DKLdhDkyhNU6Po4skFCOCEoCr05QY0yGsfpMOGWv/VJgRi+
Q6Y5xrtoKNfNf7mWwAL537elSbViVKYFkNGvuaPmuLKfHnWNJIL49Ke0xAh7Kwdb
SgQg6tDbuuxSLMNDujptIMUozSeXlQfiKYq4YI3sNgJXv/AcJ8yadFARZd7x5goi
iWzB/NzHXhnGyiRbhCHm67Lb6zodO9EE+I/wwxZVK+e3RJvCKyaqbR1yBIVsOahF
7apRhEzfeklchyEkC0QXAbxF3y2okbMpDl1tWI1cj+i4Aq6AB78n6SO89hO3SPJm
o6kZttjA6w6wOuWNYgeOKlGzVKZtA4b0/Oqgn62qslu8VnpBX5MRxwnB90Pv/6Bj
A25mDJrRkGMZ1FObYLdwHXpj/KY6u3UozMbHikyOs37CzUh6FvYrufdfEsttrVlj
auoowhDoh0ysHsmyd7oi8SmMVCkOdki0XyM24fMUUNkZQmZdjgAPrk8klW6TM+0v
gbeOtGtYfv6oE+crKwrhR/uzw5VlqL71mn7r5btJyEpilbscm8/YMG+yzYTmt7IH
5J4d+oFCO/oIQov1foXtHMLR28waY8pCWlnsFLDzqIs2Xc5XCQygvq0uHrjq+Xvh
/Go5H+IFa69Gs9rMeHE7g2lkxTw2TOshke5+1BfNCOvvED7zvlmxnnfRyxn7Ck2C
YhlXXd9zztJauMw286YBFMXiZI2Zf1X6/mrItxTs0EMA3DH+twWkuqWgLnHQrhPA
nETdyxxsk67Qewm5m9SsKwWLA/Zan13tZogn7KLWcG5hRW21aClFe8igSzbr7QHd
eOIfzw9hFh+R99x5/W7aEC/tmpZv0grAQthSLX+mhQsV9k9PiJ5hBX4iSCnrdJAu
GXIx9UVXUzf383kXIyqINxwqUePrf/K0LgC3gjVqsEZ5iolceAnmKnJKosP6EZF6
Lge+TVcvBXQg1gjJF3J0theqZN2vDE1Gtj6PHkO14tu6MjptDcqiyeh/FQnak3tB
dEkYG6BvD7LJEPrqH8ZIuk7CPY0T0PgOj9i6a2FR4rwBhPAX4Ru7L1NMt8GdLZOH
X4xjXktBfKW7bDfneaQex5POJg1zshKzn+Bq8Vg5njL0tN0Jfiwa/PLHR++VBKPb
VULr+I+pHJ4/6CcYlMTEM8LW9TPoRiGMIGD46eYtd5FFokq8iNcMeKk6Ti3kdLdT
f5kiGUSuFyswPFfoWvtXBgCTqUx9N0mOfxNiVKbhl5p4F8RvHlFrB3Aj5w6iW0o1
5/547j6mI9Mux09C/bVq/71vLGyUrxQqvC5MzMa/ml83oF1zwtpC5ANJgY1v90Q7
Kf/fClfTjGlt/i3GeOdErSs2QurllSI8uTrNsb3TwBeU1772ZoATiLqlXNwcIsHH
dsx8TqmGbeCqSJ7ngRZgqo/hM8csxH7kR9BMSZQN+LN1D+mrutsFxOOD4rn4O1Og
rDE6JPlxsOKad27lb4j8tRBMoCSEs5Fmq06c+cS93+pUpYClFMgZvPIkjeun9VUu
WC9FNbjIjs+EvHwv7B4B5hFOTkk7C4LcFeW/Lc2uDJ6eHTn4z448Dut0H+eHwDX6
wOl6yR0Ff2jXjrfvgsNsXgq1aLraHjY7ur4tzOeLThTR0tq+frz6aRuo52v7shjz
Qb7/KEqyjMhYgrQ4j7qYgIdvO08EUTHYSPnMUoIvLO4jtYh0+ktm244Awos7xfhQ
2sXtHcRH51zt1OGiVNh50SjNx1unfzmnLAqpsegwqrtzPfLJ1QkIiWYd7P6jDV+K
B3ppbAzCKsmpRgg43ulDMwG+0Bxq83H8ByUFNVIL2tc61Jp17n9a9welxrkLtb9E
+QywkeibaZ4vx7GlUrylB1GfSimgq1UQKxtGb9imEAvl1727IFqx9rIWNR62mw9/
DWsxwkYwoDiSThtNRS6yQQT/zx7jSHY16Az24a6LXxYPF2agjPYelWGa56wN8ULD
v+QprzDMaphnP0J4rdwnak0ygkvyfmLWECTLbj6st13GWT1b3kgeTt+r2kd53B9U
2jDC+wjVBJ9dY/L9t490m0fhYHxWU26C3AdsoWITpyqGH6wegiT7fmx4Uvz2pPgi
BivQbkJQ8Ig86KV67rbQoZjjIh/ygWeigpyHMbKaZQKJTix+lPb8CexqOhdkLMqu
p7pa4I+b6lwhQxcjWt0Bi9MVedlmUM5HigS/1GZDjFbV/LxCd3A+lm0TR8Jn6Iwu
4dkW1Rz1JfD/7/XQeu3e0t8DS5jFcnmexBq5lzHLEfuf94Rmf7guWddOQAeXIlHW
nbVN75mjChcEbaT+WAfDy/4x2CPGFhdOtpTdBQXUCisldfZY4Qa/NO3Ie2RqV/pY
bb3uiLH93HycHVsDtaFd9oJwZao207r6xB2CQ/nM1HFIDfXWJrUz1NmjIh6mZhC8
jzUcPMc0ENGJOZD35JAsAEAIZs3CGKw/+zDvvRsaLZoaV9U9b2HRkLoedJFJXuP/
IkLvQz4iTUtmZYXrZDkzlgUhOZkZNXttC20x0MVclY5aYBLrScasZ00nvmQk9NG+
bbhuBxlccT5xJd8F5gKFUTBH+1gnoCzK+ZTmsx2bHL5cta28/BljKvEWlGRqBF4E
Vc0XedQhMsmds+0b1N2+esTQla2i9eGyf9gjmQLl+DDYyckKV9j21axjAqloknLY
SepuAQqIQNcOETLmfcSKTIecL1XrLN98K7AwZXD71ZyUeCy4fnvP5kaGTS/db9gk
ZJ6pn4C9ERio8fOMHNUcJRy+OSTAl/oiAhUdGCbLKDPl6cM7+1tj5WAV/R4emghi
U0ukMHZMuQqT7d2gb+hJ2JxTp8e7OzZVPt7kznzjiooQchLsusdGF0gyo6U4MBjA
Qj1Df55io6KjrBtRlSbw5z+P/6IxRpc3Abc6XU4DUKlITO5U+QVvc6mI3UwjtBVP
WqQjHZM6zBXMu1AViExAjpJUfiuFyG/m53/M/AWjhWRm5HnaaY+dQrTbvQznpv4R
LT+MjVX794/Cp5/PZZXBrUHxVBRnzO6fv7UOM9aH6DAsa0O0G56Hgam10aZThMV2
16fAgzo6LNlFFwLuRvZOr5tsINvvv1Jve+ESCv6ib1qNS5li4qNa1fmpwp2uiX28
l6K2jHZwv8BTxRokB4eBjSfLLJ5WBEy7Vmrh8jER6faVnK0OTyFJE/9U2hVgMnLP
z9Kh0oHp9//R1Li5/yGzhQ6l/rPxGXxPB/4VbSBKfu8s8b9XMw+zB2YKTZksOK0d
3/lxJEaYtdiNy/yUYlANES7GSla7JHevRKk0zqCLiRASY8/9pRWOOlp17SJkePQy
ejZcrWWvrAU5WufaBRRI0uqun2+w5rONjW8U9sX0349TbQ3tZTPvmIX1SvMI8evc
+tQ/qzqIwozD8nPTGVgVgaiYxkhR03BdiecwCndoT2+ONx6FzdAWXhxgN30lF6K4
hiL1rLAXxURHx/gs4foYjf+n3EOJN7VLZEF5qlywIDxABt9Ra+xqn1CNFN5DM4vg
fEuUFDxO9t0/wX1ZnK65YD8nVQM5j0PbVDRDkJd8aKvGW347QhFOMVZ7h1WAbBRo
Kz4/5JGr9wS0ChZy9ElqMItY+9POQzFIgI51e84WC3mKf3vTvXhyco842ebEcl9f
baw5rFTKyNgR/xupCQCAnlPl3P3CTsFEsifctSbQNAv4JAvZmVTnVmkY78a5g3w0
Idz8o4yGT6fge360ghpfOgjeTLfUTEqAhH1bUfbh1RvPqmo9ovAwy2+/Hz275UsN
j4DnE0zJjdNG7xXRn7EQ78E3iX6ptQ+5V5xLWZ7YzG6v6HzZufdkonyrHnOvuHTk
NFiXxLk+IZb0ItDWvUX8l4kVPMog0v2/n5VESwD2ItFm7RhAAivXvjWi2NEybDVE
uDEu4qIq/n25tpN5m2c19VMswg9KPbfdh7oUJMkGzu2jFNo9PLPoXQ0xNRUW4A/+
r344hCHK5DWR7RbmwwNgnS5IdnukETdF58FP67XbS6C4F0FvdLDTrVuyf8vwVbqR
4FKiaYD2Wecq3H/J70yj2ODKK6kC+Lsm6zBkFkTAV/VapnuOKuJ9cGINKw9M8rqo
rugNRa3mq+MdNiLkUOwM/73X7u/NcU8ma0x3uOzaMa1BsSLV3RicvXhdlpQ2SkkP
e8g9dF6ZZu4I87SnrUEMCYgYZ0YlIU5yLyQytgqd7tTp4pVcQydhVmwAtS/AltNK
CRSh4KpGBV5XKgvrwhDe38fqpjdQZeBHSRUL/ZBU/mxd/k9O2Imts+uU+xdIdq7y
4Q3OYo/yyVv5TSEFlQCezyLaQTIcAKjXpL/DbiPZxwkmtAPtXJa3cqecCKPvbu1H
3eWz9441bll5Iswys9OQlvWUc6YuxmzAEV+JMRe7rpweRmmHPuYXjgtZDo65V1AN
ahtgG76OsGBuhivHFvlIyutdRH+Of9t/wAE3jlg3Mo6tIgPEYsoqot4X2Ufub1/U
ZQHP74B6o8vr5PnvObMBwUx0xcpllRO1kIvVB9NNTeJsLOmPwP5nSi9mK6eLwz+U
XwZJkFWAcvkinrRKBbT3fy93rC49NWA4okL8A/lecs9VwVf3r00iYhEAgzC3Jx6w
vCGVQffNJcljEi27XuHV2lcsRmu+hc6cdm+MoTdBRJTAVnyV3N3eOrbhjZa0t9Ey
a0S4aOa+38PZGeU2Na7lcmKsjHCLwfURsWoApo9T1WlzVZO5ADew0+xLC/I1R7x6
SRsfOV4QoxZnHLc/byfp32AV6DR4kXd+C0UOzkQFXqG7AImUZKPveg4dh3NjHA3D
m5OVl2mxk/cJuY9xkOJbUNjK+h9azax2G8ZTZ/TKMUno8JOteOhw2LKL37fyOG6v
1xGxLWv0sTwXJ/Gg+uaQcvZpMXaztV43OZt74iOG3V4NQhsDOMI7sC78DyjZfdxr
FjoX4Ol3vChD2hzpZMp5fB2DgYReKMskPvWJ10o8Wt6GXuC4jyCkP8vgk8pPDbCs
CEUR3S0uW2EDHzLYSUi88XBGY7WVjf+c6Bp3NzkxaOkGjWjqx480Y3stD5YjB2Ag
Im04kFeA4vhbFsWOhDoZymZSoCbxgluRid6ekHkfWCX3jFmeZPgi2pN7yrG34UVQ
1tUTf+1nFAGfIBRBROU+o+03ML2ZUULmawtc+KCoBMzve5GS1nMIoPyV1ar4/ouI
4YfeXUeAAeQ2sbsLLwftVx6fb2UlmTmrVFlnlkQr8EA/tOBMN8HubgWtKmDvzcL5
f5xs9hSvW44BA/Lr32P2metwLu404wq5LFQKEAyHEQhW+mQRqvN/hzFXZgEog0dX
pVa3uGXRfzC7tgTOUIBCJ5gQoY7voZKLcAhJwTdA5/FmfSNab7ZmNWxOsYUr8oXs
EcUcIVgXf0lUrt7UwcLwhK5vUxvWNDyEofEeQfzOIN1Zrz3YuK+r6H0ZGZM9Yss0
wE0W+wF/C5aZ0o3axYGmngAr0694b03nGEaptYrxt7phO9nv6gC12fNIWhd1t5a4
tOrbKWx6BNZOYeB8+YBDlPei1+1qv/R/DFRB2ptS52dlPDIe23BEymYcyeUjJBPy
fZOuSCQJRJPF7QI5MvVw9LQ5mp78FlQwd10yWdlUEYBtEhDfGvr82tVK1HmP5QlZ
5ViRThoh2t4mruQMTYpDb7/GfIqvLZqF1TFQdC4pRD7jVbIJA7M4ADjMQNzwcPTC
hkSqtwgB8r+DJjNcGXfiIrJkupsj2JwYv7DdZILcBAuUMqJn4Z/Cs4zMjefr9A6P
CPisQjKDes+/aZWUkMbXrPvabE8EhXJrdxoH+c8uEWpLRM9VeBiKPGpsLdhA8d+z
mdMBQrQUSaCLuRLBei5yuNuD1n55HPlOobuyX3JYOdl95Q4bbjo8kV/+HvHufqqb
S4o9QXa2abETg9Y8CeR2sBktpbAHqmXQfG0dR+nlRMKZYfOpZoKbKWQ/bvik/6/J
NYQAE+1q/IdwDUFP43v7KOsRdHJWxtqnV4OJqeX8vnY8DAohNY7l6pvpHE9kHGFy
StUz5ACShBpcca79kArmM+ShDpC7NBoXaSxKmQ9vKKXTm7sZGDgO7wYbGI+T6nDi
iGvaX1fmA6E6Zny/5E3RmVRbbX2Gp6hSr+s6zQJaUHVZkJwV1EN7b3Og9wtMogu6
Hvikfxn9gqQOHsU8wXQUoTRD4CFphXZM8l+Rc35o8KiYx7l8LI0nhNzO7PSzsXUF
rUzv34Wl1oZM81HWcEkNKpfaVrcvSjIrrOEryVgjT6pxiEeaapCDJZby36Ga5K/f
vWV+3xE6vPSCBh+LBY755j9nern+kOOBF+3WTawiBPzrPS5WYr+zVPp9/tfzhXqW
+wECF4rmGMvu+Shdt+M2AmWa6fRozsPHlVimxayYEzR3fGDuy8WUipUuLgzgyr1d
nsFZy2A6P9G1gsZbli95AYJSjiyFjtOewT3JLUyJewpFF32c1MQ/NKnU+/xYl5CC
MEakBdTsnRmfyZ1wzTq6s87hUCocTBDa1K4co2l+5EjdUI4S0yqkIvb9xP3QYwOj
wxN/i5FyzkhBI/2LpyXFHu9it2D4erRXPWQaObQ3AtKdMKfcVl4SzOB+woVo+Ats
uRFoJH1f4u4Lv88FQw644dFd9uPaSgRe0y1Pd2D0/XvSI9isk/jHkCiCPouIKuud
XptmirDJKPy8zxTB4cqmUgiO6q66zx/7HMgpqYbbC7xdciZ3u3KKd7+l+Ev9W7X0
KtVp8GRcHUFI+tDxWfN7VV3XwSaNPS2Z05UnD9koHK1fjlCFXcA168BGBUIcz8Y4
fsbETQ/nWcuZUdhJe0zJpRVhbVTpBNUpZGsKBDj5+TNW/NSgeVMEPvIY0drl9gEI
DkN13LY/nsNk0X/UHRcD3orNG4lqlwHmQRLHXg+39mNw7/ifmsyLw6826U8mghYi
T1QfyIK/qlZn8zWrTdvxMx2jnpAizaH2goitYODqjJ7X+HudTztqLIDlKrgFKyNc
vYNMFeU4fwEwoQJn2yrjAN7PY1wvZN0smT7Z72gLpgooA8BCcN052b/pvdO7focg
wiVXy3Lo9pSFfAmIXeI4/hqdz9D8DXmWXy9n9X++SIfBOkB9khknItyI2jUDLMLw
f4Im06cNbmDAFLMxfWuUImTP0M+trJ1jDTgrpLfMK++OBSQlsJYthu9k/36zkPZe
WRMncfUusmzO+3mE1hanYlNFg75x3yceVSMIm3I47Uj9pqFkxLluCS0ZjSLgWaMJ
ROSKD2RSV0PGyrb7hxHowQ2C4MbtBkk9rutP5ltB2MYzMc2vzyN/txo7Ri9l/TQC
0l6GFMR07H05lFg3Zb+FyKgJsoqOpniv0LTc1lmyquMsMDNZQ2DiWr8HTUJZn1O3
jTnFCrGE841tH2oVj1BRTJbyBbX/mEV9B8mYIkDc8cdJEZQBfiufC8RvmUOyMgSJ
QTf+hwQWE+PKiQZf90qcu9prmEdKhtnUVserc2wGJPMFLOJe9yAKqTyhLpuOxoYP
HtjfoJPRi/Kdd21OwmW8r/x/bEqtrfGh1/SXZhr9acmeaaTr6ge+XcgbSBGrm1m3
cnhhvpg0kqAk35ynEjCKRsmW8izlAIPgeuzouXh3EWJgtV4yXj4nSQ1/3mrH1uh3
PZd0mqroTM67Tw9Ys/tuIFxceHn/zN1U+HlBgjqYISwCEfKsyejvoWzxNS5gvUA2
l6xV2s1zYKCqti7Az7hVNJb+CdVyFJGGm0Llk//houcLOqYQpjyYTn51JlhOVRdb
lVSekRRaA5DITCjV63Bp+wQxp9LNeVd9Muiimubq1TMuBpKD89KjCLy0HWoMt+wA
xW972mmU1M6p/3bBDDYqmYQXml/KkNRT81uqQRvI5sfVKr0/8BtJCFoRT0SUFsw8
zFFlOKdiYCRsKPyZCkX2W7aRcPxzr1oKyrzlDpD6IxJHdNuNRXpc2CVlJIujO01F
8poTEoL0jJFgtLS5hDQ9uv119mBC5fJbKjRijsFTFbfduUT2nSrc2dX9HGQ54LLh
YAZfbiOFycPWAk9xC+lADUDIKXqJlo9fDVrDQ7jOs4ktRqapFbI8e8ywOtQDvGrn
6MZj0B7FSeZcWjkQZ0l/gUvUw4vSgawJSnL8jzPM7LbowsQvigGH0sxvpqnCpl6R
4CQw7TOoUngLfGMehVs24inFZ55+VgRQQVa2casl4/TASNQW3Or+q229emlmR3hS
JSKEnp/utG0LUfFYtWIlW0G08IIU0lLzx45psVdAnZZNRG4gpKEAta42idp7olvn
nAWH2fv6QNg1vDUwRgKp8VVemfMnvtIvtmUC+Ek23XxBgKFwb7tKiV6CF94d8XP1
iayQQ9mCwxgoueuyJUvvRKvhNY9k5r64NmcUXeLS2oa9kewFawI3d+1Qz6Dk0+d6
S6HUfnlbmhlmVDX7dPn4wfkVbGnJWJ598lRCCTmoj3A2cGnOnDXypEtbqNdGIrBj
px3r/DDjZlp/vaLJ4jLL/c93NXfzjO2VS9R8svk0rDS6aj3VQZDrJJNU2XcS22oR
MLagF+1Ck/Dlr28sosc6QYrEKaNwAliD5z5zMrZTjaO881p10cqvW9044gH+NjjJ
dUCeBbjjI48st9OGzglTqES62i5XGvwGmourbEKZFnDGPVnpU0ENGOszR6m3OTnJ
fKalBkkxxepJSAamzazD2efJbN23u0QScuLXNSGlitaEExyO7LFjk0zOyICO2++z
08c+/gD4Hb3clzEmCcuBG3RUm2kdH1L4z/FJHEJKmwmqlklmuhjYWiZGFuZQ/CAW
OjiWbgich/c2gKn7an0ffaxvNqGsNndi6q6wRovc/lhsytRnWZ7wARh0u3nPpmeV
UFqYHjAG0xiA1e9sxwlJYCcXXnuCVh6++QC6hp0myVBkRL/LGK7ytVUsxA70f/Nk
QI0XKv+iFnEXk5tLQ0+nTf16MeKoB0WXGjCmlstzK/NEQF3Z6If4SUck3pOIJhTH
/5bx95ulGEGRDXaKX/n4wsLMYcLqpfrgmzbuZ5eKj834Yw3e9GmczALsCR8IfcuO
spDHrztpTRxeymlh032k9HDjuyF8h2khk1pELAHGIZyZfky/DhNpX+Xiz58qTGr/
ectrssjBmAuD1rNgEb1l1ODTh8R9yk48mBYXrPxu/iVFSNfIZQhY25GufIidHCcx
ALtl8BhB68+aMkZcW5AynokZiLwgd2Pmgvce3uEQh6Xtp5aggC8MyHYxW7e5bC19
3qxnw2owgNAiw0BxI2xXa0lBZRY9fDkUYUs1Ze9WFhCwVscpVTkkCIRmmrGIVfi+
eHs+ly13F3ZFBh4cIi0TFIdz00e+7+HqJC+5Vc+q0IjKX9cygmnQu9gf/I9n9NNj
BP3bZRl7oST9hGeh/065y7S97uzUUa9byN3xmYaU9OLLWD4f7ACeGTeYVE06Yf5h
nnd3FQKz8mvdGJf8izRorScrvb+0UeUhM5AHDIXQklgShH7rxsz64p3cYKSI8LjF
UBIIjrzCAKXandJG1h+TPjFcq5VNb/39upRYBJz9xQX3EN6MJkcnzwQWFN4X649j
dK0jl+LStfPVMOj8DzA4CIk+I7ewaNRjFp6KiLXX9zwtSzqlfElJmXzbBVIXgJYI
A46OMDkN4Y2qQOMctN2bBgV3KF3rAQxTh0HHJZ93OKu6P46toH0V3gYO+2K1lOwU
0UqxAjPRkxAl0eYk/gjnITadWtX/RbgiC1/lwCWJFWxhaJ29XZ0zS8ZXDS8vOBjC
o1jBs9WDFLMmk6W1WH/tlhxfGtkMdCnFT0SwdUJJwMltbz5mOxxbszV+IoLWt7zg
OfzdNPUkmRA7Ag9PygBEp8fQEDFYlAYryOM0ubxC5uEBhsMY8dwNS/eykDEg9uYd
IZMYHjyrnwIoiP394jJsBDIdkbhJZ7URmrTenBuyhMUDQRFL35x+heZyvKQ6oA8T
XBjH2/fkxKnhqj0MSAQpzkaK845JQz2y2IT9u6/AVrXyK1IRacBAdpj694uETH2z
nf7p4c1CIVVOG8uJwv51KV7TYshhxngvCFKv1XGHBz4NPmvMs2R8upTLa9NQZfzG
7GX0TqrgabFZgTED3UgtRlRS0B/HSd6Wp/XUL6FtDWVtvRfGBfmPyQu1mG5u9PUA
1Z1AJ2X7as4gO84t1o2uJtDyL0j96HhEJIyYPjMjvPzJI9adp+9ezLj8Q0iD35er
N+Cjr9+ugk1JnV7sh4h3VAmXsFlc9fwF3T9vNKfy3nUwmymH4tGyWZ1LR29ywjyj
DGhgPPz7escUB921/Esw/j6n2xoED/wOOsskyJmOCaEFpdd3zGlazCH7oMvMDoQy
UPK0gsr+Ghft5wPC7np6gUZygBQLuWI8P6EWQEeIscvCPhv3N5/hphxoyTjS1hYy
ffeOcTHSzeP9IzlW2OX7Ph+9OkZE/Lr2Xv4PYTBjO9wvu8cp5J+UouyaldtvT5Fp
JiNS5wipcO5h1B9xNgU6PXsO7s+ZDuxj5zYjRxpNJP61ipG0oBqqXxUvxoTW0Uu0
/8JPbVKpsamDQ7Ha3+0pEjXABK56L3pmNsFc5dOHtNWXzhabivK/425DUF1LkhFo
JMokDaGS6N41fPhxNKkr+emX+GkWDeHpRDjDGWE3tUyMdvShw0S3u1T1V5agLaMN
P+L76KFlj96NibC9o2/5HpwEtBu8nMopSTamrMwjbLqFOwFrWD1bt/+n4aO0vF7Q
Npt8d8r6vnQ1fUVNYLUIi84JgN497c1w1dVtN+NjwM4yZOcoNPtM+MhE7lumEGbn
d/hOvC9aO2lKlF/TTJq3Bai1tlZFCR2IPfrlGhDbaCx70T8ybM4ewYgeSSMEJGm3
F58gYRtQydjtXtRVmJKni7jShaGikYtWqtkzdqZagNSqwByvYhYaUbkvCS7vB9Q0
XnSw0M+ORzpsdR2LC3KLFNVvtrpyhcL5dOlJoCBynzJhCzLK5iwtzFlRFBhE7fok
xB7TvpKt6uDyZYntmgafXMM8M/E6HBZv1QWinLwhUXIaG1VIfqPBWrxzoJDRjwI4
YW2wC2RbXnZ3613Vw2OExGuV5Xis/l+JLPwpLNgR2RUP5QsfRwGsLPudKw00aGdX
of13nDSXOOavl6eYTgGOxQ3IF3rMzjRASpM9AqtTbosPt/XLxyk/yrd4npKlt877
TLBpeAso0kFT1VOlzKuMb+jHljubh+RmoEqdolJal8lNWpFPlklpvqNf9wz9Hx9O
heKJy/4UoFQxxRXC6kanqQ3YeztZ6AgbJKaoGnRbCy069bTxBCw8cOkuUxNRRJtA
hFO/te5II4dxXaFI9f/LqERTgwgPreruGe/2IkioCcz/akRqZVWUycJ8aixlO+Eg
E4XrThKQLppK6TZrZnqfSgUFVoqVEkVTNbT39gMa4YF5AG93HugYZfFzwr6WS566
xqx3v/OBOViPnqDqV0kV/wNCbQjCTpRY2wye0Gs6wTDVe+Ks2fIgEeedA7kl4KiB
wpghbpFJW4kCMhmO5VdLMGs3NfV5EwUrAnY9m1A8u+bBIf8tA6CM39jfHGLgPY8O
/FOypR8Wxhv45bFwIuIcus9A8Mux6Ue4RaULw9KJ0TOvI7uV1v2TbqdxqDVEenME
EYpS+QUktjXh5uHU50GT3UXqZduiD/CfyV33ZmygZ4EixiOGjqmEkbTtw8Qr/vIF
XWw7be8iMzPQ1Wjyug2m0GgQzdfBbgXHNQ6j8aZBlK60mxp+lYnuuu9XeFYHW2ca
VV/SGyWvck+7xRzeMtCLOpQFDspqIadSJFCRd32Txu3BlNrw9sCHLcRluoiNCeCc
c+LQVhbs7O0Kw/dqiJtvuEAqauDTx5gDjymLpHahga6cC1l2/ofMA7Zj/6hOlice
nI08TUUig4uJAFkZ+n8SHqiGfSGeCqiOD29kia73O8/jkz3FcrnFJlxNHNowR7k6
dwI/LIyAIfnyyxy3ku3baOtIzaNFWBdcIdifq1H/lHSwFu7gBrSAeUvv3oiWEGxB
3rhBbRnJrIN9wkeefCFO1sfDwR4uDxsiNOYGK2vbXGU7Fb9/cSnITXk1qjltwGZ9
5bP7HFPBwyo8P8DloxEJrEXI68SSvfSnbE7SstkbpuaGm50E/PXqSCZxh/K/ubJz
cswepbFczLi3jN65iQSds6k+YpWXlcX3MHtvCeRbTUG5JM+Nx1r72/a7M7GlxAHu
V6mDZg/Q8XDCaKm/4YM0UcKNXlq8Sss1K0FWKeYGoBDwlZvFCO+srEjq1b982b5g
1OKpg/Lue84Od0kmV7dcogFTtuE2Y4KboQChZ6Wte5t0O8p9qb/AeCHF8uj3qeYh
JqvPsJwrSxNldf7U4UpaUjDpCV9Hfis0T0ZWbllWokKjIASuRzj1LXkz5MQD79vL
TOEvn9AZ4Lgu65OtXxWGONVEcfo8bEyaWaymjezxZqyIp/8JboJL7/N8gHXAWqzj
11MQHnlEgXQKJf3Zo79/qwFf7g5Ks4hjocZGBA54W+ozSM+24I1akpPfhniuvLWp
CRqfBaHqULHSIfa4e8f3BA+nb2Q6w8Pcfn059VhmTkSULeZZ1zXHE1C7pn4Jwqn6
fGAEGkj3Qnbhvk/pEdCPbIpgeGUPskcBQa+aQWFFvcFgnQJwVHkamSWa5ZlQdA+2
4bgfv+NAdEfj52FTOC+y1a0CObNocKIMfrAkjzpUUHhUsJt7Rkzqe/uFgsJf3Aig
VJxi5eqHJRTa3HWMkDsAH+EaiQqCrjjonz5fEEuqBe8ENmPqRZm9BN8o/oed8vZ2
YGt7xXvbl+FyFMU3inEZT5LzT5iH7BmgFkQqJteHC1mBlgC9RciVilVO6NMmSnHm
wwkderMiJyHFpKVx7HPRQxZPjt15BW0YsBJFSK6RNyzNMIT9FdTCWiOkDvPkG9fI
S1JrbSnaCQqqZz3rbOtauELLRghfjkQQ47YpVD9VrC5x2PQ09cuRsT/pqbTRnBb3
s6AchthK3sou0/mFNs9ZhyTwtY/AKqi7FbgNB/sXqpdDkPMiqLFOQt8Jhz3mGsEz
ifGCX1Weh7ZBCAn5Kn+VYFVvrAadcVI9aef4jACg0y1PPeRsiA1avnE64HqObJ9Y
WpbvYFJoeKRJwHXhH7VMiTZ3mSpWxDxBOCrDF8gQYLedI7cOnZUFzSvQXozVqX41
0Nbr+ajuV+wltjzFiiJDCYKqavNgotyKZqftGvTEHpOivVFRq+VBpTUB4xX2+jaA
lR7Nwamotq/LWs2i6chnxYBfNG1tVImxzi/FRrjmlY8fEG/+vb1bXXEdUea0yRG4
m1gEqutxsDgip+lLuqnB/vSYtqpyK375QEiS4DTsit30yu585tDsPXoxQa5G0JIq
g7L5/uG8h6D53OBPWHobZDKrTjvYpdQM2Kqr+cT4biqQnmvKLsvaB2DBRMG5O07s
9eFtUKHEo4BXzUDY/GMN/Y6dG2Fl58FJPYciNqv5rJvLtaDZmL8gDx1ZODRaVyPD
cINTSSb+oVVH0UA1fWQUk8HA+DmlnO/eoEm8y45pYgtjyTCZVbw2e/nAYDQD9OYr
mCuVqtL1CyXbcSMiHr17cPe8YcyzA9LPWZtPmdXKXoXRRTkg1kBplTX32HLET+sJ
8PzMt3g++HtF2cp5JmNL7cf2z6Dhr44SIJLX5PnA8uQ/HG+1IOU2J2r/tLMxlwcz
psGklDvwYU18v8q/HnGkrd69zyqCsCxt1VtxLGQh3Ze5aO/2BT9G+zjA3e+U5gjP
bBiPypckkp2aiauiCyQQ0n98zagI2ubrwGv7p2+xSfAukIPJvfrqywRpVq5yKfkB
rcFRX2rKF9/Luw5rDPp5lX02DUm7hoTgpBCFqbXlPv8pnUS5LXFRpRBCEs1yTf+W
qqdIExJ5IKTR6GLvkt5Ka1RS4lyvJyVtFWEQpWSFWj0OH2x0MzpCFrPm8B5lcXHn
l9+1SSGiYqDK5EzBtINtR315hnzFGVsZFKl74lX05kYC4lit603TrpQe8pDUB9BE
810WXuspSWCsyWEhBNysw/fPcrEhvBsHQT1U8cFgC2Ax1xBHp/1vdkwjXX7jhuYX
4Mv+pT9l99KdJrPOg1AUniUsSKvoKwZ0YPBu2vluVQeQEhxdi8MMHOPiAHwbBMWC
eMYJ/JaeH1xQ4oe2mJnBXbAAyXDyol9K6wmvN+rcriSgGip0qHnkgFb5XLbBsBYt
YldMEqxFZ2TOuHkE+Je/hPdqEAhJ0CO5/MkvJhJjYrK2VBakWyiJcduczu4niyp4
3jlQ7nwuG2kojZ9nZ80cl9S2UXm2O2x6oHrLvYk913YjhYiiKVM8xx0hgU9Q1aj1
FuCl4MyqErI6GQRUg7cdsbWqX3kCEH1fIqa688uEzwdfWualJebfTwwJarx23I2d
TXsGFdIbp1FB+d73lQ5ARFqR4QpbRtmbMUN8RPC4V8f5ERVS4bUp9gdigV85ebQF
EKnWAF0sV3en7PPSpxVqM1sXyAGm+2jldJGC6iHEvVQ1xGoDVxjLBDzBM1yxoAv3
aLRYEMjW7QnEHZ+ST5ceLwsj2YgiC2CNhBa9unXSNVee3qxyY2bxGlg8WPr1+E3k
6yXdRjoYngDqlsfAekQBvtMi76E7UPpsZfNZtWJptTjlik+hRNkqjTNK2MgWO3+p
i6t1tFfpESMAd6fErIdNOfAObBMb7RvPpQjxanDHEQNsU/shL+UHuPrAwe/c30VX
6lI4x0OthhbehUR6jkmCa/KC0QLVqhw9v1plBe/crGBRpsksYHOGoiG79gtRB2X3
7SB2ivqsSbyr3KbYQR3IkZjLk4sFKvzdhj+K3WR4SQg6j3iuShC/bAsMC879/Pxp
A7Dxltsy0ISwsI+zanuoz6GIRtklhNdm+n75+BvLta0D4A0PicWq6U8DEsP8q1Q5
M5nWFMm+yOVvIl2zjhFTlrFu/KsH1UpT9qwN1J/FkEwifi+k226aafQnLCof897s
J/kGg/Mhx8Ub8gNFuUc7d+bqNeo4lwqDERq+uwB46ZwAIcumPI0LY2I2PT5xILVA
+yArF3JS7nVj/hMalr8PZj3g5s14MUS0T5x8/qXH2MlNsfLMOcQAxrHAgUfKrcaf
F9HNhWQM1bWWCbhZsZGC7z8VmJpJ87yvgtrT9mgmiatz4XNHxrTwhPNOheFsm/MA
/RzI+Om1uymufp/vp7Eod3FcKAVUFenMkStB50DMHx72GYcHfp8hUNaA23Poijeu
LmHnMJy8smWwnDU0KoNeiubK1aaq+JAatXyWAxUxcVBG/HAhYCLw26k0/hiDvoIh
qtt05XQUIzeUr2j5EOMzVlSNTXOutGYLbzRZp+gZX9742bTm2PdYqZMDsgrxpCBw
Lf+WgJ6ZWt1nU59vNs1o4ZjfsVvspdy62uh0DLl6vRcLlLY7/f+I0K5UDuN5IoiJ
GowNXepJTR+H2laVrzCqeZLywwLgltpKLkxeKfiDLpcenGBsXhjZaVWmcWpN5pr3
ZB7PdMG6ER7zkiH8X4RCPqMFKQ4awzaYBi5XRfvbaie3XzZozObupZT3XEFx+JID
nsNG1DsiuBwzrLY2vC/zdPzyTlr6QzBQKYZlaqXMn0gZXjkqvwlFDmBHjm6rngYE
eaiYQjyV1H4KcoM7Cyxe6zLA1p+BANINiArFPnjvf1tdpnOtXtvs4Xu9ehIZ7ILp
e5zqMyo35VEN+6uCGBUQar2YfASda+u7U69+1FQONvZt7sX82caa/PjMSjfgTGxn
WA1TLuwgzImKibHP0jf+DVsm3o6drIdI9RYpz0Oa4NfXNuekGpYOTNs1nPg+hOmo
PktPVWrTaOF222hN3fp3NN53QyoGJzAGNbYJbT2MSrhkcvL7xEMz7zJrjP8+qVY1
Gq77dOmhcK7ne/ZKG/VAKn2dzkB8Jg5gE74ke2Pzw1SRCV9qtToBuJtDiC08VhqU
W3RlxiFqckDZDzirVAyn3ajcUX4Rdogm7V47r1dKw9bz65VkFkEftr/84BoNdoZN
T+pE8v7gjP0Ekyu0WWrIg3lTFD0LcUyzhoSVNFruozTdPFg03OG4ypoQlRKD8Yh4
PdIRAAq1SGNaL8D9xPZJe/GX5jU3WEU6MHvM7svmcOMOmWfNNlcaRlqF9R1F8LPi
K0nguZo3NmKXeHJ7BVz9IasIhGhrEx69sXCWrfrvh7SkyjHPvAX5l9Q0n18laII7
sk6cXSrTp4L8Qr45EomdyBMk5ooHFd6UWlC4phTjfRvZdZWc7Wk4m63TvpMo92hL
Zhdwunj9dQ74+4CyIFgNlGC+N0zbJwNz9qdtKxTmcBlH6qg8lRmeN4ONg5spvZh0
ZjYhl6zyuKMpc4mNA7T5FkP1cy2SNUiaEeYqt+sO3IJfDjOA2/c88FFG3ocIYTMR
rncs+me3v/lIWwelxC9XufLKfkDIk+Jkr7HCz5mpPRAOjwVMEZz9p6mat0sYMNAk
B/NbAmDq4saHjpNYWWZD9Ta2pA5g7kLvcfCoQF9o9pr/YbaMNCImgsRiA9B/bHyz
zT50FIFNfoY4cPVb7E86ObcIJcFmeRRuu2I7A3zgcSUEvec38S2ttSB+imLsWO+x
q63Id1LD1AJB09R9yr+doU19LvbUZDzQbZn5qjF348yEejHdKWbccwUj6KGUCWur
uEBrrBj8Y1Kuuxoh2auqJOYVkmrV2S7ZLGg6XUTT14rq7pfx3ghDw6KkAUUSeaeU
z7xvlLARR0cS1UpSQzQaIE1kSVOqtn2ZZO8oA8imL5x8+FGWxq33v3vFnyZV2Yn0
RNkXNARt8bFRiWkovixvRVJ5I3zmAkeI9ORLQFoFueC2Jx5h3C+cumdWS2S/GeYn
6N9HpaS6rhm7gtAG4J1zXGmhfKUgAkxEPe1eDxqBR7510heZDYB2uFunO9FdpS4m
9HA2Ie6Bu0Cas61YBntdjlOC11H1ZRs1JK0BqRbvlgQ31iRr1yZQK63I3EQFSbmo
uGtERgBWd+kW+iaiyldIu7c+BaFH60flvL7A3bEksht6NYaDlKF4r1GYyEA1PguS
ETC6S0vgCsUm+s7ZX3QX2zr4SDIE0PfJYZ66uB8RYHs+HEXDysN1Yhzsd7Q+ji42
kNC6g0rWjfLVgrBbYVuo3hf018IpvtC+QJ1vb0LRrObRMT6+D4krdJC38fNwl4Qc
WYO2QVyxjttLN3vq7S2ljGqPTv3wj+w7SHrusLlw1pWgfxV3Z7+uwnC21D7yT3wh
tuACDA22BjBeAGo4VkC1V4/AlnGDEyy+wwbXtxAwasFS+rTbHmnCXxDdMcKLQThd
vGI89exOE8s6c2fDlfhC3rzG3mKGdr6R8bS/e9E0zld3UodaC78EHm5XSPnv/0x0
6Pxg6JF0D9u2Tm8QlvX5sXl5d+CanPa+BVUSX+RuX/J6lw/0yRE471nh5Qwvn0B6
kCRt40qNsPet9tXGoX+bYyMWVoXm96LQvbFUxMBnKmKDEobHxZM2yQMCdCBoMM2q
lf9bHhDT318BPUAUfeWyfDAQljGyhj++o5n1Zm0DZ4C4rbhfmJWkhQF8cKm/PG2E
Mr16GgjLgDolr2V0fCMXYp/adervnry0V92q0TKCZRkpKIXNp98i8ErdOmW2QQCb
TRfWKQAofaVy2zgoHq0lP/0Cgbl1KKPn06XJhPPipr8AKldXe5JPYPfe01fcNGVp
Ll9I1br88c4GOloFCzL+lgie8OtE7XaF+nDVG4igl17KGripGlwwhrxr+TLkK9eJ
cFds6lDm9N769lN6jW3bYqRR/rSUJjSmkDofbw8+DY0jKEwT2b91z7a4PrTTEgc6
oOL/emC9SYpYFJdqIDuJJAfN+0xQ3X/ESmsan4PovXs5ydSMVMqaeB9ns7X9j+uh
BecJE7Ss4yvNr5DA1kaCv865Ki367LS7FaKmgqciOgqAGO0bciG5tfn6KRYSI7ZV
XdhnYvpA5gkVv5PUiaMp/VGo2vBCUyBTGJ+Mtvof2/RQUqmhIELTZKD/wtqgA3qh
ZP494u8/nJqHSCl3KGaRpGNA8Xtw35dffmPmnghIbiGWoATc1/hHndGPbklfZasi
klU7fCPKMSzXIfhFIYrZTxYxyx9E2UylHz5C/3gGWOqYmkirE0dY9vuJ/Am3zJSI
7WdxJNU8CHftTdvDKshnD2Jh4//nG4gIyskRgm2ZlwCpdW430swLolrnwz9s0qu6
6flr8dm/ORreC7XMBEkndw9xLW8pu4APgGheA7K9Sv0Pt0DIpThXW/d6i+Ldat9Z
GtytI+UATLJr+MfxIqrjYE4n7UT/ELdLLxZbOoGmCg2A8Dn/YKbt2q03udMQ080o
rdgrv2psDdAg7+++/Z10Ivc7oK5fjpZJn4TIIY6dNcNbLwBmWFG2LD8zHLNcNn67
Ng3U2yNFnFmExFe6I0eDTGXAc6MV5lMb3nFH6Z4u3yeTqxIPG2P1MX1BGzQLz4R+
t829qunD6p3cFvtd8TlD905VUL4CFrEMbxSIAA3GXOTJM3dA63z9ZTosFLkPlqc9
zKFwUuR37CsYGdFc69JOSBfsWW5TuzsGwhz8gL9Y9zW2zVQn+Ck+Xfh8j+tObbs8
vQGptpx87GpzMx6vmq7giTISitO2F2PfnLZBaNIP7jV9qb9KLoDoQbiK+2Ad/b9O
X2nusJTing6UDk3LiILJI5VcrG0OXuy3BYlFvCAsbU2Tz4nRabB5mAHdrjEETBTX
Uv8w9jqd6Fg1VgArfN3jkqJ9Cr6/3L9yMi7kB5II/COANpAN1SObhrkXXltDmwXg
ClCR46ORQD8BjLZH+g6G9uGgBCAqYafW4NGPiE3K8l6WVLpYkF9kYk833EgJHKPp
0tvicM4f2pnoNepXzfgZ/3pG+dncQVXLhdMhtNiuuKfAUzkrGqRUFXPjakLl4CCe
dp7IWRxVHk7ofBPZ1O+cACi+TxrsUraWDQPDdyt8CBGsCannvMrURqk5ChCwtlN5
fJo9F9DWb5Y6Nq3Kfd8NHqVhM4+m12hr7p6g/4kn8o0J6Ub3d59vuhanpOZFVPer
/GShD2aRDwo/C7KMm2Urj6P7R7eMtRQ1An4y141IuJTlBFZQvx/KtvW2YPSquWYO
i4h8dCgIly0xEuxh8F4nE1IwS+b8/fMdmX+8Urff7GlBcqnIahMMzZcrHJ7jR6Ho
vVR2MTP3weMAQ2I/5H7CFCPP6+Qe2vsUy2RzZ9M5lW/H9X7OYHYQ34NkbjWNksg+
Maw6mi/OQv5uIcus2ijzvY60gT/BAkCv3j0PUl45W998UbBUtJ4Uv0hphTYpYYlp
pCbXWVqxYj1LE6Kvt3iiPpfRUt2x9is+VXunHLxu/vMJHjDIK7bRvNVDZC5PXzdw
AK4MmiNC/hIP+C5r1rMVKpG/NGMB4iFJZCTDv3l8IV+rPaiTVo/XzJxxpkB/sAhI
MbUHQ/PmyujaQSnMe2a8jypBa36Z7rPe1LQJWg+TQoYb8+E6lkqbTeh+iFAhVV5y
5uv7ofsu9HQc9L1PLRnfzrniiyRy5ajWbig26RgidxvvBnAzGJf5MDSeSc+jaQ+9
uMT385GAuPPcsJKswkSLiF9pRQOF/lRyazuf3zo0K/dYcqCGJ8odIfSddp3lGuJV
Yc+bqL5G7VWGViFlJRbhFHjMUqCSKJWD+Evp8+cZdzlHk3Sb8gBgHXQ3+Z17+opi
ly+7lMxOuo8sxj4o+P2Ac2NY4xXoInN/vanF9nupdDS64kBz1PQo9mxTu4g+nn1U
p81/cbI6ohsRJz75djU7IJ5NO8l/PkusSk+iB+d3pGAz4Hfr9ORccO/Zgdg1+OeN
bdnsX50ZGdTAdM0E3jqiJ51xWEQ96XPhrRk5BrC+koikAyu9dRuOWx7FZJFC3hHH
5ruxB7sdeqgZdOWBsb5U9PX/YxnrhQyd5p/VqsbCbB1xCd1/teYtPIw1d1ZKmrjz
ULTeyhy2yE9INK0L9sFpk30My3BZ1/ZV+wmSh8ZdM9nHzKiPGJfwN0Q5qW//DBzy
q5c4x1RjaMPuFrhhsNRWZR1NMm+dVSdpcRYJ1Qp2dHmkG5JmsQUUaequcsvwc4WG
zliCmGf0rmKNTA0Zh0l9NsExYEOkR8rox3e3sk/i5yvDxHFhzXDQH6F26SR34Kes
IF6Bh0+tMv2xG9uS5/wN3DZ6SCoiqgSyuqzAiI+vOaBmY+mp4qjDY+GkXsv8l8kV
k8olLJrPFb86F55V68QRHFO2u0GM15he/v8v5jD/Ddn3w4+z0eDhjkjvCgrne92v
bH8UmvP5Skq8rQVBpgUtfYY5Dwq3CEQLo8UYLjfe9WhGsCIrAuZqqwSlEiyC2Qzv
f5KRZMBn3P4DocNlrpAvr7R4k+V6rlwSUWJmgdh7le1x05dfJuXQwqpffgakvrzs
qJP1v1oCI+udi5wJ99bMtPxIIXbHsS6k8sLeIs1NMf9SCMqLNxJH5EBWq2GuUdZg
MQ4JSSdYNjzkbA4MNm22GJQo5TEkKu5DqdBxJYtaqAAX2IUnsOY+E+WO1cRLITXK
bRlCiHXvAEUhGGOP6mCes69RjBYqDhdtL0wZu6Odu4v1x9hnift0Bahus+El2Lf8
YFNAoKFzmQUA7dRsfkxmPb2RSNLwFIvaqVjfNRkMTRpaHzk4D87nsNN67qbjbNhc
H2Up/qdSDntXPKNx3ttNiYCRwVAIHp4XUViaFGVs2OYouDHDtLA2G5EFZTOLeTxW
q+cU44U2WcEd45Ug63K6nD+gDOIhhriBt+dKVxFwxYePpVqeGeoN98HKBPBstKFD
7qkrzsm2jZUoV2Lqi9JGqZ4GO5x1PXn8Ng0ciUEkQaCqQqhsIi6idzLZGmIIjOgh
fjptayQ5JkUVnaYUPWdDTDTaW6rbqGEIEq3854xUXClVl9CDKPTOZl2/U1uSWzg9
6N2yI/gIu9JO8HRu54rGgHDeoTeIu/Ba9xwn2dLpZUCSIuUUxyzkurjwE96PCdVR
i3NAPWlAabx97FxWVuCyuB+x8J6CaaiOAX9pHr9454Vg8708KJFpP4qu6DVMGSHc
FwY0vWx262aY2eIEIxcrpZ71dG06AaL0wfNyV1SeQJLqdItO4pZzGbP3DJqvLmTP
v8r3Z0R/X+1Idjd77/vuKcdJPoV+/j65LHKQehwDcbKaJsh7TrIlBeyPl5wfCQj3
SgKdoKs6T9zwQ/KdOiIt+mSQJlvStqE6vBCP5DHbWX1oHhbCDZfBkAjK4PjjIMBj
vKnbtDkwyR/NWRTGv1b8A5C74oKa01xXpbXZqRAnTbiUYBPHRNclGrgZ5hiSJ6VQ
YVYnHUEJzQfvwG89jHxEoWB6ZjC2a8tMbvK3P6/AWQXUFZf5IQZNKKkrvAyW6SvS
y8QBEdOytcAfF8P/ryHz1Q6QI8bPi7ZjAMthP4yL4wQhw+sPRaCXGCPrDyIaWAKG
Qi58mcXlZLJyZru1+qgl1AUcOnitwX51f+3zuBEjgaTgMEDaJQM75XlQP1izIM4j
GZin6MqYJDiGLrDuZeqxhtczEBooWzVr/MdZi0+r4s4wjhsJe8zk4+zCV+Gx9t3o
pXgoos0vpXXvM+M7S4BGvnWbnStwwtRIrswApPCjxPWG73DDXabo7FGFKRJwkGqm
lCU4dv9uC0bVZBRn9zpswr1NESCTIafxdiSpmMcC6+LD7TkX5QB+3/HT5ojqcpGM
RT6rSzwHU+8v9H2k9D/CWabjGZOzvk0cq50b4F3vY3h4lxGkTx0GFU0aMsCvlpDj
T97ljJ0MKRtiNCQo+ngMw3JjT6IWMH6kUS/py2HGQhUd7i4ciT1/IexlcGTUH2Pi
Ojuo2KUAtKuSsSRe5d7KDZL90bLHKd3mi0q9TXQIv+MrDSllQcNlQ1m63ai6Q5h7
VEglrz0uEjt1Ebs7zl06bzjY4Ny/TQMLfHVi5aXhngRI0KsTL7fx4TrngRAOzddO
njDX08VLaerm4/1lnoDxh2YnDILUuRoaju5TKec7yASd/brq3fQG0RpMfzRU6sG1
uZjWgWDYjXFtJDIpL4EmlkklF/z1WF/MbMNnGZHRqIfomNf3pTLzIJtcJ/tvOtUW
/Gr2SG0efNWIswHR2M177e4eaGwsWiOzmuhjQCYvFswdA1JFGHEiRbYJ47kD7mEm
yiPkw8rESfRHwooCJVoY1AO/MoScdmeABbSIyEbfj1iBmAbf5x0EShaFiDaeoKwS
D1rtkhj8k7ScCcpTg5u7eobfA4Ul4v9gsDfg41SLzNvxNoCaWD26Eq62YiI1MoQP
i79WcdU/SgE0J/Se3+0QOw1zoKNzkhmPum3DP0HrMlBeLphjTbCEAJ+f9zRl/I/T
oIV/jJOielePQUcleR28igfBIZ8e3Htj+n7GN4EU9d3Wc9rR84o7EcsPIolgvJfw
IhUx5iQIF2tKBR4ID6rfLNcKMpFxiGPpVaEPioDyhq16hfTbTxMdl5IXaLnokWWX
fxRZiQ8nTgrcqPX7rqXHXUlTcGWwCGicmlukD1l+p7ts4ipG9s7a5ZC0ke6dH8W4
Pw3/b3GR2Y+EezoyCuJLE6WZhFMBy5YLIdvRX/jOc59znrRtHfXufchzfGPbKbSs
qe87L54vg5KCWnFuKx4Ig/buEUSGWlult5Vjt6zIS4mCqicpIeXdrE0aelw/Os/i
Im9MQzRcX2M7ey6p+ZpPjGhrExyNMjw6p3htb7kyMr+TwRZmeWEJaJ7othatkXCH
fwPJcfw6DTb6C917yL4r/6aFcsu05jpQ6KuWZV6W6rbcO0CFnfxPP6I/mjdaX911
gd1D5LvaTIpoK/JsnWPQHW4VJ9KhjcFR9ilnTAlB5fjluYEWCweKxg+HY/SEKLUQ
MW2dGhTy+/CJbuEpYhzVe4sAsUyHEO/XTOX9QxFxJ0F9Ui8RAdwnZ2QC5ETYSnzF
wTqRvyzQDbmXVJiOKwGB0E1A79TK5vex9KqjSPEyy8f8Vi8yTIfIGAllS45SpHBr
HeKnps2osRWamn1hiAab/k4DQy9nNSyE6mh5l9U7LNa6AnBdjSS0hZErRJIRnp2k
lym/Fz4B+lzMV8pVj1uxfWUPHvyEfAhezh8HRSZGb/e2apZonyscb7Ix1wZHbuDr
62L/gnd2bNwbyRmYmpiIw3KmFefc5qS008aAIYLFGnk2HiKYP432+ADZOGZScPB9
NnoHr4PwNY9qZlbyzamXoqOiiSA7dgoUTleqB6tQVpGG+PtpXrQ24MFmzrHz7mVT
zbRdJvM6cJBSR2PMimp2m32oZ04vycgFih4PJ5MXglrJIFsPkIvNTBmqIkPhtB8r
dekghKlBhmG0I8tprY6IipTkaiVcrgXXmHkbPaFHTsHcaJjkAe5EXUVlk0nFeKLt
Z5rIpW2WK+M3S/V81Hblxkd3wJmKSzkEOt5K3+Fq2prgcY2RAPk1A+iI3+fggV7i
Lnnztva1ONSImspNPtxoT+KN4GdbtCBBRFKqTfWXSwnnqs5MmG30tKShGe8JfCc+
3PTKDSIWyPpl2ghEOZmRuhUyQZSirfNvih35i3zyglqSJM5gRT0/aeq0ZAzaFbiY
6a0IPETLzag6Io+njJUxsuYlYeSc7T4h1VWAGhMf/UQzziqmvQPj3kq0ufMjZh7o
/JXSWzH0Ttq8LK0pXrjplNlyCQX08Xnq737F+P832x89YUiaLgL7Rq8VcyNgohUw
mdm/plD+steWOOxNS4FPV3FETS2c2WRFRMTPMlTjG8KuImNqHFGynW6+0vC4WJ9V
nt1ilaZ5Hu1S7hX+GBXKgGOW66KUlvozYdmjzanr6Ezuw3mzxt6TkGIIrKzy9ayC
b1vpm9V9CP6K+Xj8UuMBKXJXO0fcrdDP3gbvSvIJFj/850RpmUF3wjC5uJIJ9+XY
5DCXlQLerAX57SRBvHKsKCPCK/PDc+YBTvseaxgWBQ5w+fBXDocLSjd1bnUihfvt
qHohvJXwRCyr4CM1YNmcl53LY5upEOr0nkolYkiScEKeDqP9FzoXyU0Kgo+xZ9xX
Gux0pFbqSsmvarPBIh/SRAq6FGN93xRBxhesUeZ8lZCgWlwFQHVF96Cf59wtg53e
2uquEeMzKqTSGXtvPphzfvw6jbPNXoW+JLFmymXsy1byVjLKIYTYRJ2nzC2JwNMZ
mEmai++yMmQXylsDHbYWZhJIHDI/tq4cC4vrCGaGryRR5AhhRF+KXPzk9eMnfekR
nW8STrqHwW2YrHU/pLHkypAufaQxcpMXhjKc3I1MSGO/gU2yYkfiVTBsNuzmC132
91eRdEl1yPkY5WUX7+YnQUdcQfBWiQfxWbx7ze2cUhtNt9L8EX+c+rROQEAAa4o4
j45KOU1ObLQaMTwTzuI0CovWL2LjGKm5wFGbNWy8o7YvzxAJC3Wd14DboxnbvgeU
a5Benq8eINag67K1vJZ941EyxW7XT766LQLYa9De+xxXRy/bvifSut9eosu0e2tV
4x2PqVwOj/15xJrQAJWap32HCqDyFQub8mojRIJTCRTcNb2ccms5t7NynRKABtp6
nBjafBPIAHsQj4ybH8bdeWkI7yJOt7mpAbKlW8lUHIYkrNRRE3e/JmWY1Dh1OtZH
Usq7CqmxdTs1ouXOAD6Cqm2QIg1nKCDrGu1QZeBXwdRuruQSFUL7cPtu/sGYwViS
914bhQ1HlDrRL6wMJr8aZzygPl5ViNgximO36uM2pSHi7sh4ovGj3AG8DI3QC07E
EzhtFt06FS/vuC8HD8rtNzstPIsIHZIDCgHpa4tqILVr59BB3L9u/cOwphDFBEnq
yh7Kcq1g0NRXfVU4BrTmuBb4LbTxj+iEwCxNzf9rsogii5eGntNXVO2mhRsBk231
HoHZuFc26BCa35AMXTdDVT9dPE0KG8sbyP3JfDj6pREKtA5RAHfKhRr2Y7ZvCDfb
ym0rM57R10NsWUpJeBnzww6oLUBVyn2d43+1SZL9Bg6UfFUWYNkqxJkLPbUwkN4/
l3dSQkWz07Xyse1iyDhVAooL3760guEnll02W0unThNfkdrUNLDm3TsHphAnnDCO
185A2wL2l9brtW/AI2lmoUKI4lahEYO5WEg9K2hsAD8SteZW2Ud6mkCq/uwmvgyt
6blU4j4lJbYEf+oiNCPWkSqoo0d19e9SUK+mCCuq7EPnTX5nJxmOXBJXUkn0j2LZ
rTgd4/B38cEhJ1Vbpeky7iuCgL6wshypACHK7H0cO7QW2cslQ4kmBI+tmjWB2jnJ
oWvTOx0A1HBPQUmUjh6ILBT398szuer5zvg72bXPz63vQjlXuTWCj/AMBVy/pan4
6otg5rSrGbONWTavL6W+bW6bbKaLIdTNw+6ywWybYP4oFXbDTUJose3aLAk+/Zvp
aggZnzTZKeyKqI3H05FqjzzENkYm/OAwuTAGoKaD9TF1zQFUextJ4jUWQ797RI1a
w86TYEz1ySnPVDBVfdz83B6PtaVvbOoKtayeidMIArn5PK3cNlgxMd93xXMMF01y
AWTw2GkSPMfuFQtBS/hdIGpyVRcgyzsXdF8JwEOVYzl4KDtzkiOCd6Aw0DpCxwro
k7PJhCJxGMUTo6yGxc+oAProNQwy0foteiLNaOELieBVbAi3MYBZh0EB0WbuHh5V
wOA2vWc96LZyh5jxIPIUJCfnikR4Lyg95VmeWhwABzqgE9p8CflZAt5F5vXONxzB
0Q++YXxNCcc6FwXnigVGr/SGzy+S6lS11+Lfv7NEGIt+HkCQvxkeuxLySbhAoC8i
nUuVvP9LuthvX6y9XZu5SbJi8klY/sDZcPnF2JZOlNV0F/47mIqplrjb9U3LWIqu
/gSZ3LLZJFZDyHNF0/Nr11Y2s2z7ELvJ4B7o8vCKFpQbgA/j7UH0PWVcpveWU9vg
2tODQ8BYeZ1klhshA1FNJttnWHZ2BvcytRwpYmhu8dV8ptBfciOabCM/fWKDvMja
A/qKyWUSLW7R6FXQM7Ap5rNFcNckxruMdJT0QOWznF6YVQc7CU8tKVJlKizWgOAL
9Yg3mJLAUmpB3qA3IB78vrmASeIYQBe9zkymI9q3S0F7dOsBvdWghLjbiPzpy8kM
CWz/af5Ssd1+Zn+rGSkWrewZz7h1ujBR4boh9i6Pg7gLyw8uKTooilyGHO5Tx+ow
3/ONAnXxgeepfCyp3SHIGpAzSkuUKHyB5EbSyd1rZM/iE7Cip3EYQRMdBTglvgx9
Oh4KPb9/NGj3LiFHd0YX0Joa8sWK5YnEu76soyO7FZap4agxw4ix1FBRHfPHFWqo
wotYkLPSQR0405U0gBsqPiTo8QvyD1nVPIr8hqUgoajQuuyDhiY30T0VMRXEGwMM
0FEUCmLL/djwZptYz/+UI6zBDgiahVHvI2g6/ecAHFA7jZkaEEpnTW+fGuwvJ7w0
KXabzBIUwJqNYGuh2GhIZnFmR/Vgyyd+bG0aYFF+S0Ea7V1E5A+utAt7T12o7U/Z
SQLQXUnvfr9hGwEIn1dursIgQExczsdkvAvgFeo7glNyDmFPlmBs0MOnaa/xxToQ
XWp0sOevEKfMlJw8uI5V6x6iPfOcCTJxUvykOAcIeK1WxqPVp9P8Pz/5a1iMhWF4
ndM3rsyT5Hwqu/BcWD2Jof6wpdWe7qTPGD7qj3LLRzVsGKpg0acgkOWr2bUwZq4J
1d+pn/s3jVLhFFmH2IBZ1kAeqGxv+n8Wvq2S4J5Xs2iQh3SoZ+oKcVyPlK+XM2zv
70ETtqBA22quzmrQFeaY5juLdin2KwpncpO1vEVTZhhuglHorxIInyR6QOF9j/Ld
a/c24GOHdMZWG8iExNkiq3y9XwMNn9LcD6BbzhT1k3AFAKKcHEiIkiKr+It2e9AO
/nYYS/62eyPOeNoImX4BJrF4b8exiXY+hOT6mCjkEVXnTCJCb5+nhNJMkzOJhTeC
ZWIxV4PrTFdL4t7WTF+M0QQ4WVMAb6NYy086gbxQDIplcVFg3QZ/M0uoxXU7/Q6i
wLS7TUMABq8fLMD7ZyP1pu0VuoNvRn6p7uO4sSby8KbTPq/POcjzumNLzuzJ0zHx
0t3iRfwQUf82+6vlMoAiV3Ny6j/Mh5fsi5lD700Z40gaM5f5n2mbKcTWFzD/FSQ9
34YTv448G/p7oZvLDweULueJcW08j3Og52YogDbD2uSu8MuKhPHByTslpOcIn1Jx
bVadHiMAdK556PdQwL8/aIW4TJ1cjSUzZdZQvA0xAqqlb0kGgZOKyx10fmubL3Ut
+wNIoS3PwkwGW40Cx4ZE91zyF/R2Zd2zba3weqdhKo5SrNaso+c6PfD63hH8wtdR
HtTCy2EYEB6lVmkA8X0hws2Ij3pm39GI46NtowN7GyBxoGTkyKck1Sj0+6bzy3Uq
o2ou6pswfoWMhhSHiscv/CUZ58p2AlSFP98OEXEj2MJYkTsUKdIN+BoibmlILptK
0karFgNvOrmhGebsudWM5Hpf/6aus4Lj1ZO9sCjGfK9yjo7HUMh2tLnxDKDU/a6P
XVl9lIA/+SnCQB2up9yWeFXnCDWuQO+EY/oALmprvteR9mymLozqi1S59tn7QwEH
xtupN51Z9eymY+b38D+DQkZkxVo50Ivl7htw2ZMsGSFfdLFR8u5xI678tXhoenN1
p2HoGsRVQX4TJUpXiQKRIZrhJccYlyHyqavINan0vC06q5E1iKu59duOsAdIjIaG
ctuhJJtSIJmF/pTJP2FEn9PaQE8tBSs6BCA4O9DbnfIGaigdjMFo5X0QK6nFvWUs
++WkcWAKNhZ6hjzdAHOG7jCGg5RfP3hqCYsSUN/0FvM/OiOL8M8WhT0ehVD6ve1+
PcHQywbr9S49I6yixGfaCCZ9JJGLWHIR5mY7vhluXxmyI3mo0zIk9C7SDzbVtdkG
PAMeXwFWDOiOjTtREBjGeT5wXnmEretStZOkCUyH1oc5N+FqSXch2b2YAX5rL2Q1
yH0D5rY/afwG7Wa3KGbLWswhxOdbRw/4QvYGJlElpKl5S6QuxGaevABqW+uPqtwb
jy0uJGKRETG5Ov3TVrNZcRv7hDSUq6p4/HwmlnDkKHQQ3utXr/S3AUeHkZFlVXIb
wliW/A+wAtUWXB9Ay88X72Hp87mgyXBWmynty33baJYsvQuGSQltQanDIfIIGsOd
CBn0G9piM3PzV1xrG4CAMmOf4cIt3y5dZjA6blubuCb/uMvX9PAzGdtkHN0UpDj9
YOqPoYmIqjeYYwjmXr2/del4kzxlWJBUHkGjHkNHUAcJ/r7SLFWxhv4iVqc+fbk9
7wK/sm1/+fLrY5mCSS89vF8cw+B0EQRbPNpa/O/T2C9/8fP/kCa7KjKquqQ6IxUD
vLah+FcaAMqbl2duGdu5/TjG/9VpG+izrmoqjbiOXuC1ZYuOv+rHs1tvvXD+sdpb
xSHTfHBfRZyswJMQxkl9LpkB+gDWvMJAEKrhPRRRq5bBLuBz6Rs03fsDg3BKHFyS
0uCK2eH4SbSd0NFMNiQygJiWo7MJGsPKBgLwWp20LrgprWZqcebk/NDZ5x4dhuba
pn4VIXl1IVIEa1S3yKARns5rqqMWj3rMlfxFzWnxzEdfk13bT2XvhE1AjFSpxxBi
ZGwZhS0209Gr8f7mKfzqxdghaWLdhsqtgvlH0Y4i65W8YzppjyiE8jvoFGehAC5j
SX4VM1AWUHgdKiKuem5iR5X803YXyprO1/p1/rd6Gn5eNVjwj17z8D9bGN/Jwsva
rz8UCJJW6rsqjsgiDRsdX37TEQw6iGAHkzFnnwS1j7FOBebzQGHyjcWb1k1DJ0Ur
zEvK0fDzriBVpl9ERgpOtlU6sICBCf/mgn909J+YPC8JepX74fKzGt49GmJ4Uigu
BKowFvx2pORm733QFPcxZcoRTmA0m0hUtEXxZlQCFO/atVVOgElD60Su5GVXlpTk
vzDmf/bfuJfwl4V9XKtDcRCFP1WrmFkvQrNqQUQs07LrFtNkp9VmC0CsCIF2q9Md
Spe25ZFWCU3yrd3mGFjRdsd+Ir9d5EPlzdGVbXOBTUFEn3VfQ1z1r6neg/U76q3+
VoX6YhQOpwcz0+yaDnTH6QcRyNPPM/gjG0JWX5fRgvepG5DzQ9PC4uYhUuv6nFRV
F+hdNz33a/Aki6VthSFhSWCvMh7475Jc8JZcFZ+UXsMsb6O7a4ef1AABm5+dWa+U
d5fLqvzZMJjM6mExv+mKzMkiTlgZWWxxodMTD7Zf3oSCwjK3K0GbieZCLcPpsLWL
cowxynx3b+tqen4NsV/jUnxeF88pdlKfVCV7nn/IMf8s0k3OaP067Bry0foTIWyp
ZInmtW5WM1bq4Wp/aqZvs+4uT4d3GwWOFsee6uUQCFi5u5bk4Wr+v88sN5FQHHzw
YdgNDz6jyKYvM2ZLmqK8tQFExvGKyuh56EeVEzr2nkvMwJG2QkwPa2Hq0TKKr3wC
0cZ+JmuRitxmo1e8EvtpOUZ45JJjIr8XE6Oc4pLoLowHVQc8yzK2mI2MZb/Rq4Ux
QCB1RE/b2ZpelOzGJA3VYJhXuRGB4g7/xGYfpA6GEbf2KcNcYRmtTtxNPPVJWSSP
x1qnJGams9612y4ZpPA3qedTP/7OrXef7gGo4FXwj/VOMZYXiQDi8XETSAGgzcYo
fmAqhxsvS0hkFNcGZZoExzVnV6Rofu7G1XDC/8Vt+JGLvABEGSHdsYh/L2pNCCvv
Q29PoRKf+5vq1Rd2gNPJZ84oMWrh6eXX7Ls4MM4JKvVwfOSCLrtMBpVokVk0KMiI
pc7v+3FOIzEGrEA727Vp14hKglC+7qJUdh/A0zmR2R/m2rNxKvnoDax8NjM/PIOo
vD8ecVpv1FaX8UMlVF4I4pCyLo63pMTp5uwqVDR6G+aNCAXHTBy7lrT2uqMoB4jd
P/o+sKf/rp1bm8cdyw2fYcTeyL+TLHUp6lSyT8UQRMo6crUApn0Av/ZStoJDx8fA
lLQcmjFB7rwmlO+0trmgw22QJOCrx6o/4Ybtn2mhBPF/zeweU1T9Uimk276TQM0N
WEpJBecRQY/R59hIID/UoCawd3S7J1xOyOLzgPFPt0VM5WczNi8BtyFkGeoEJkki
fgkPC6QIBsKW6nLa0CB1UOsKfZA/rtrT2FVjoMOnLBNxFGMM0MkBVIZf4ihpHABB
bVUQQwHR82HDzMs5snMUovyxqnOyxMDn1CdJv7djOw/qmk+e9fRsaJyZ8VimY0eT
+CUxQlMvUlJA8siG9i94zH4DBe/ngOzugAnJrJeX773E/00ftfgBABVfsGX3bdmk
y4+wHiM/aLM3OqGOM9zlPoJgUyb9BXeHDbYFoyUP/K3MelyhcLinaB3O9S52NFBy
QGkdoX+7K/fPkUSWzuvHEJE76TzPI3aoBitDV0tSXOk0s6Kx36RjErNkBUiNnDJv
hOCCJ9MGZd6guOkLfdDYwNEqxGmsGhnQGVN041gFJVUvoKl9H8EZnDunDZ6LSS4H
7IF+sMt905xSW+4yJN+gSxMB/PAXvx1dReQ3X/mDWj2gCjuBLn58e6AZdpQLhUuT
iSed/kSffWf87C45Xyoxou4dHw76+6IgxYoHEtEbBWprY7qBbZzGKwSstaC5+Mor
BxsFqg5aU96DrJnZ3a3XXRdNYjEMvbawyD5+ethEF0eGKbMpFqJemXgtKdZp+b51
7jqYLCDc5lQdgZz0Y7XTlC08UMhH3f9IWOYMi0q50FNigU1DNb1tpQC4fHIprTDa
j5+CX9cMAhML1Llvfw+qG58zh5reO2AoQ6eXn4qDt/U+ziE+KVKR0x22PlsLeHeZ
DLVq8UNhh9iUdeepLktxCsBu5PRCc68EgXh5+Kwb9ca7Ea4ITdvHQMgoQ0qmTC+t
b8kZvrZxA1I758DoPDsEHB25s9GZS2AiARpKNdZ3gVikU1aKXYtvi8hA1Z8hpJ0e
UqqzZ7KztO2TdvN5ODDQwMxeEP8UH7YhHnv5OXzUh5qBL+a3VPYUFbhSdvon1IBG
dgqhZwlTg6WDo07xm5Judo98ybZnb5/POg1Hrw8TAkfRI6VCXdWz4RiBKbkFDJSN
/i3NDB0U6HfWEouGtYepgVQ6ulk44lUaBst2z/ehC9XkZ65Vb1WzjtfozNpoDz8T
I985g8jJaSF87TTj2cahFOiiAbhiWx03u4o4+/v+dM8d5E/3LT3A8LIuD/T3z52L
NbbsFl9jxmgfZrsPexbYJc8o0VKkcdqz9BmLDyYgicTzHLz3NnbytDcXQ41KoVmz
JWb7WhWn2tN3uB4bA7rQzUzMgPAmWHxKmFxMA6cHrBvghiAqP3yqcfeoYn/8/29B
gaLW6nIGR9xzWqjy6KcHFFZv2x2kig6WkKyu3lNj7d7YVaimGZAjDbUaPIk8LpaV
7XurgcAOLrTNj7Vx7GVSD/AiQQ/CdySt7bvWq5ecFhCpf1B6C4uyJ5IyoimtBHKR
CiBp4QpSF+e8Ajxs8gkqYN8+7XpbSg5zQiZ0z7/1fG2Oo6WeDYcUDlrqL/iOtsZn
3e8yeqZFtEdiHreadCZS6OO6oXwVFQZ84rqI3qraq9ZVihWNGucCURB47qZooIkx
2/awPwWKqKVJUfkADmfXRwJR0tlq8vpirsRO/J1Vd/8j4ilKAMalcCEYci6y/dTG
BBcnpVmuc09+58tGwBsRkwVl6GUgzWoxvrOyX8VA0MgY7RPQwA+B9VAd4K0UOodP
YO81fjBtGOkDldLnPaox8IBPaAbWZDXW6jvI3TIfoOeRTfW68ZBHCNZrKWA/ey4G
FDyPafGVNJKVvSE5uDCgGzN5fKTpMJOlDIXn20ogWAQGB7D35vblWVy11WWPOXfA
hzqDcCjlea/4UmBSZ4XwRqGwivWLkL/PztXqUDExdQsgAd0rDdscMqOjAapLMnuW
n5R9EBwPtaPBpBt66NR236ATNW/lIynyO4Zi4WrZB9ACkn+IWnlD4/UNnxUFhAFj
q5C4x/26+ujCauwEmb6m48EybjLKS/33XKUxKR5zsxjZufQ0goKY/ymfbR+8eGMD
UQkW8cN2VCbSslI8Y283bma6SDLN39W537sOQDr7Ka5SMLkk9euCjvmLF+bOiRAI
D7+55ghwUimNiFo3hcX5y9Bg7weFcXwOH3BkHRpcoyDc7Xp9SijYhjoGv/sZG04x
cvkU/2I4udCcRt/DLxoVRp4Xy8yJKeAlx7Rhr9M2dUZ5Safn0pp5x6xaag/D4E+2
zU4V9UXfOG72vDtBEy0yjTyPPQFKAYOomPqFhfBJiR+0dNAYJWGR+v4GFz+AajHZ
Z6Lkq8dC6Ghk5cmypm25jVYtuJDH+tU6Z5XwKDMSJrUmQFE4kDTHPMnRK9M8PzWv
Nxjuib67eY5O4rgXG3u2w8XBaBCa2O8uGmYzKzQRfwwloCjNysuA6ZK3z3ivufBO
D5Rxv3UP3LjqhaLDORoPvcpFokN7Lfhv1va53sbCshhMCuf0I4h9Q5VA9ULZFBeZ
2++LOgEnyf5+ouq3qaJdHiot+K5lWQkaWgAqPWVNAY9DJpYTCmyu0/itSjuL4fJU
5JtgUtCJa1DSpdaYqCKYaFAqVgrNu4UZdnLCL35seEvisVb5dngpTrHLGfvDezj1
jOQMH2JtELAbCTSQ9POOOt8QTy+Q5fRchz2aaHUFHds7fEKUGGwlQS7ofL7wssim
JEXUH8bvs6sEle8N3zIAMrK5rTESu+XHtWxNWTDJ+DzZ7llhaZuZnKhrQ4oTvAE8
YP3ud4vlxQiaGxk0oCJRk9mokJwjDG03J5FmJNBluyzSpl2NDJ6isZtxgM24C5mN
vDykeala9/6QSeP33Xv+rSFZ/U/xoUa2myaAoMlyyTI1qaDqjHamCfkzm5dN0rLB
xUp5kjRTrOt8uzH2m4GhXFONj/5yew8LUtbyuufXWF4FDtD0ND28MMwOXTtUKSnR
9rwqS1bvJ/YxbOVdl3YMSB226/+LZYZ+anbBcPtNqKLSNy+woiUlt7bITilSWqaD
9vKTptG3JHvqLHMtZ/Kn9NwCap5uk++3e+otJ+Tob1ic5I/CicOSnEcU+uezg3ka
M11SMdUH2XARL/vGW8PYODMTQ8zjy7jkk74BvQ9WWgqRfI7yDuv9cdR6eYKf3SCs
/s03xsuSPAXm0DjZFyGTp4vvUsjU/MPnCMs4xFpJi7/hyjd13W4CcPD3tcaQZK8M
dvhLfdbqU2g/0vULQFqKodKpwPC95mR5HGQoLrkRi6wJR6aZESxrryCdD1e+A/H+
gk9I3ZrfIFhqw2CNVGZ3LxkyoPk0W+6Pv2vL41HNOj1KdXnQUuLL/J5SulQj/7+U
CphHiUPNJgf1ESk/5K4MIIY9IoItb0EjtuzuIZjeVyb3Rn2jTN1lQUtw8LpqH9oH
d3MfgNZH2qTbUqUQ681TiBJC/Hps8QUnvS1r7Gk874pREcm3uscVVvgzF68BpiWo
mk13I1pPiwVUT5UhDy7Q9WAu5XOhbgi14NG09byiV3QGi3R4rQi619zwr3yUkmfh
t1zePJFY9SErJDhYgshYnIqxlQJFUX6UgaYEIpsnJMKkk8mOoLpd8YRdcKX26A96
y0T1+gdUhoA1lCXjunm4b8o0THK9D5ui/nrAv/zWx2eNE3pgpF2mFzsnyD5MDMq/
COYQD3mTIre1ydi2SrnOqoJi+g+1MYg5qlKDUvEfuUUlXoazdGZPR4NiPnhGbvbv
/DRKYvTk3HGT5EvTML2rNjighfnZLDAEF0KWiLseQIdqjI3cegRILE+T7I9rr3IR
ZUsjyCMNM6oEC3Tcp+4QCDzbx3wVQm4qFi8kwd/rvasPWJXOEOa1Wh2mHFJBz7Rn
SNfpgx/rvSzWGnlF2uqIW0cazRbjSaTTehkqdJ7r8wzIuF+sugdFoLX8jo7F+AtE
ul6+bvw1EiGOx2ugDnzgiBnhnZpqY66NhKOlR8b67Ti3FEXYDOi6KrLsfTSPzMsB
p+WZyciVxIo05dcuVWAeSFDU875s4yo75vDg4ydGAUiH4IMxEHdT1buSHDl4vOnA
8LLf1fz8v7pkwaQNA3QBhDMhM1OzugbELvarg1bII7QfB14j50vi3cn0J15WI8T2
06NAUBUhtOjgnYDNCtsWJ15fmR3xRmxBoCUV2o4/M1SheFhUprLlZmjnMNmBVe3m
UA9uVNgXkvpxwnvDd+fqKDq8rPu2ytdemrczj0D0FxlEMoY1kgN/vRfSnCyUmSGp
PHOZMEWIfWuh7G8lt9+FfqAx2NvEJidQPsUzrprPwiR5WzkE9vZ5sdVtQfOIcDF+
wP7YSkDMuH9E7W1vAa/VjIZCfbmQewqzJkg3MfPiZenHfskL/EFnnQKiZ+7/Z8wp
5RPGKxeQpjCOAWWq3eTGfxoWqvvuYWERBVES65Q80GkLw2KcesFhkKtfMXWb73xN
PbpUf1x1y10U2UHbqwOHQn9uMNG5y/YD8mEc5CfR0ZMY/LLs6kDO1hskZCQdQ8D/
MuIcbUbDkbypt2cC2PsfUM0w0nstY93+E0pQUA13anwkjF1sE9Ij2rNDYnSyGyKR
gIsolnsObJHqswdYu9GEMGaZ2T9gt7I/D4wFr5OppIApSKsay7mIEN+5ZYjnA8AL
CLzx6oqVcYSe5sxbbC3wy6JvxjgnYp23U4osLzteELhsf+XboxRhyualpG+3PNLA
JqhoJ6R9lY173Zarm+8ktbkVyJ4m0lIY3gKU7ylwZchlgVpcSXNMSevqpNFUsllm
cBOzansJy5GLmsq79XH7mFEh16v3R8s73xA4Zh+QYO7U4tMrO5Nmo7cmUsXj1KO1
8UgSQdycWSIZRo0wgV/55fC6S4rPigdHshJEyX0ZCjfKdNW02GCuU4arLULf1FVx
clq8xDmfodmlR+DZs35nOht5QXlf9OtotEfV+KJ4DrQs2DhhCSGL9AjkPPMSgrHC
EYOPCaTIpDkPhBqy5lfK8RfdXOPh4/OKB2XN7nENhSbTt18anmpgl1UbEf+j3CWD
1U4fNDctHFamrd2ZYz77Z22Agd0H75+pbHs8IhvOzuVt9fN8ZQkV1jg1IXIUKdb1
fqtKDRn5ccPHa+8LMQhZP2E6Pr7igafSEWWCDnK+2goeW2M/4HR0kABM47P6It5S
mplB+jv3lo/9eU8yDGIL4hhHDx0+sFtMonsUpxckOR7pLT/y8Pu+0dX2iZBrUbel
6l3QbbiWslWjMweLa2T6gweHwqHTLOst4sGXsqmeuEv4cAxX72A8kTKpGDfYKMDM
uvb4jQj3AtplBBb16RBpYbWQu6qLWz9HSTMuNeNUYq/cEqZRK8qao/oP4sS1k0WM
52j5hsMO6ntD15MgmS4QxvBcCn2Yhyw69l9J4teT+IBvJUxF7eTwmpoIhD0cRCTy
Br/mMDv6drGJNwkAIWQCCNmVPKvPZjC3qzzr9GVIW+G76yweKVZAysiGOhQKno+6
o96LLKOMVLIggyu++TZahacVD+vkHENXT1TqFp45v6zJJG/LzVr9brfcXWiFfRSy
SIxs8mXh/03sjYVLMYzsCG8nic9yIYBj0IUG0Q0vEdoO8h1Y/W9BBkrw9XcbRh19
5e4CPYy2COGgsPuUOFMdTxRa/5RAxTTmL24INC0mQd8EkyftALHGmDvui/9vTOCf
8rjFbYrPeMhWXmy41W+hWDdsO0EKSSHiv8F2zagVeF4HylkLbTjRAfZpG6xtw398
K2qHQi935j6blL/kCxYdyT2khrNnkO3h4QkiFQGKcvqEti5SaP1BJir9WesQCULT
J3YrInd8vardkVfjC6ar3Lz8fsMkm1yqAyiUZVLbH6cpYh0lRLxgVpUfHRTxvdkN
F+hKEntGSKDNRSIaJ1wAwgf9khf1OYFFTBGkRgJzV36VWm2eKZ6fexA/4e2QKP5u
QfaLRG5OaqwnD6pcQ03yWWmJyC00PpMgpNiQ+9T41IYBpgAHvd5UgUtWVCNmnoM7
A1BryEXqsZjwVjQhxCUUcy3wYgpxAsf6bA4g2WwQJQlYXzGp8sWYRtdpyIolZ8ay
cCWeYOOzHLXb/JDCIBvKqWQ9QHpnFDeFlh8ER2KagteifkJGraC+QxbdS5qSEsM9
4f6u3R82nEsLL2W1uf55VOlePHhOqucu0hLQtebO9y28vkLuWVeXB/VXf0gu7SD3
6dJ/CepiC7XbySFf1/qALQeOSa9V3OGA6axECp0WVeKV1KQt4SCw6lPYw2KIFN7G
cLK36SoUpe5ux2bnFw8/61SaTdlS06DP41ZWZv6NGWQs48pZSaU6JcdAzW0Ak9Iy
UFDrflNaI6dQ6uL1iGGztr2zC3r3AKUPfNtjVk/i4qwPyrEjcMswraefeSDh5fyy
865F561fvZ9rqGBmfmzqpcIwo+cMXqcpiTM+jfghBOztt/bSSOu78MgenQAWPdDN
oNolXV9DhZcibvi9+DJ2usSuAxfcnKREQCgEm/IXcTaKJuamK2JWAoDDZn2pgYLr
+7+Fr95SWxjS+1x7+AEZ9q7nPZDMycrsMHjxVgriWS/2bINgX/RGg39gUIzDFuD9
NV2akQw/QoxkCvYaY3gr2F35SQH+1tvv/vdM/XgFOM32N745lidWyoykBUy2OLio
+m+0npVE6Kc1Q2pdN3xqK2dmDpwBqE09vRIq2URRqXXLYgK4WOOQtDV1iCqp5D1q
Tf/dWu7028UqHckLrLMEKhjuxcPCSw6XDDSxUL8so55evflPI5sb/xVJuJC0U25Z
WGWBJyzZpCdax1wGIP/tLlqjBcbGqqWKbt9/5yNBViRkqaT/fxlw6wStMWwzCMTx
93lR8sLZb8KxIWafx/X26LBuIQkk6E7ufBsaxTT0pCUTF6/Q20gyIpnZ6alL8G38
WEHviRiLTiDqJR+fm9q1GrB4JLIp78NlHNhClj1SGguIaJSRsfU01nCD4sjp8uKZ
JqydVBhJZC2mRQdfhHjV1Ztob7IYbaZ1ocwQdKTbU5FYr0hCyxxSvMtROb4y+Hts
gLVdlP62x6ZRb3GG7Bc3SpqPbvAHIZ7/t3cdDFfWjYPctpZUusrwAUW2NVuHdpRN
6C5woj8b6+QQsVHZXrQ5doVJUqGe4JXSnRi3eueseOQxlRcXc/f7vEBbRarDotIO
IuwZPSQ0YqtgzCuf+Hl3n3mwZrka40squPjCTl0TWdPWGwqzekbNsRp/KpyNX16O
taOnQSR+iElFht4dT6KXmDR3pyQtPOFJf1iKQT4CPaJdiVJAanrB76uA1W5GGvdI
iQu8hs0AJYCQHwjntuwLUhOlWvDJ1wZgr9XCgasOlHUUNXmiB39XoE4uMQttNKhr
vpzYj6JTPtXTrsl/3aCLNLcYOFn3WlCuA+0lTL63Pj5rxx+X/TmDqEwAAMWeyCFu
IJCjT+yAtiQCOOk/x3zUhEamMDgPdNYlI36V2OP73MTDRzi8Vo3QzJMYAHlFz1W0
s2RscVBnxKS9YTpmDthhplejPzQRA95HjluW9QrzUV6RJmf4tE6S++Lq670GzkMs
MASso/XSLhbCI2Ja0flBbcZ7kZ3nPVWLC9nL6rC6f2nJwF8X6Ln2g3xCRuKkBnl5
nddCzTkVCj/2yxzQH53sbmKVADeahIUr7ntSSnACXJa3Y3LavLV0N78Q9LXIqxig
3A/s7Afdpv4N+4D5EXI8xB5tO7XT/3yPnYORztF33wut1/iVWrtk0X65eKqg7mcj
gABe8zDc15Y0vYlgtB0G67M4ACm/I0M08O3b5b1axySKE4jXIp4JW/GpAOnSFEnu
zgmXRLN0PTJeQCUZsHzSpPdDDu2DGBR+wN5cMJz/XMZIt+cGfHJwpfu6eHj4z7xZ
sn28anagbQ8QyOyIBUiIYrxH8TF3+EWZWec9q2wxEobJ7dBk9j0KwEmY3Mag2p6m
J2FgVvvU9lQG3Me3NZS5RWz2eXLsmaxdMy4Y/8CmOaew624Uf0KUeTEAdpM+TvC+
Vnjop3ouefoCLTtcPQq3AlNMrNO6Q15erGgCYwra+A9nIXC9IKqAx395754A1QBi
8j9DT3BpcXgTfa/5lolUN65lIVo83h1jEMdheUpQOKdX3QnDzRuks37yrdImoTNK
wGpHiqk39W58jqlnpMCc2Fzk31lQFiCW6TwcU45Px/cR7gn9kAcNo0j+4zoiHKd6
VKTdBIgIeyM6IJ+mW+2ktwBePzg3ocvoAN/MeOywCbb66ESddY1NcGpoFArRCS66
8/tiy1yljsn5EtEaMQJJYwVKe/DJ5rx2g1I1CW7uKiSYdeotU4etEaz/aB/coC+j
U07hErB1ch2hvEm4m96FY4qq4x6SMnOdTsrKpZEhAVgnoqy29RSNT+XWT0ICsm53
oENRw2myTOasN493aB/5DZlhX3dtLefiYyQQByUze2zdAKBOb5FM7SrDjAFdegiw
iqdNlgMIvdMluRfWJ+rtP9LhPEodF/0pQe06Hbrb+JWmoKXpnIrIrMSunH042VSC
IFHUvRUM4n85mleBB5BJn17V0l89uzK+MlXMcW476AGPoP2YYQwVwaSfMAp/oSwU
1r+NujrorMHqx6+ZZU86MWU5tSMKAEWWMKCYIbUbJDIvTc68z/wUuXhyODriN165
WfqwVhW3biAdPjjkuFojYUnvRKusngSOqWTa9a9WmnWY8pMZ/xVRL/ZlDp3fAKb5
JxJHdOCoKwRtXlcRc/fa9EPkLTqFMObezcakCEUE3DcR2nRlQfNfGWHtV4gYKHSn
y2hcYnNH+cPrWA7iRBUOIXRleEhwEqz9q98TP1i09iCYxC6kn3Izr2ZNTTMW1roA
1WIxm1Hn+vtEU+TExJXHBWOUjZpmw+QgN+8/5VnSRmZDlJvMiSeYxgolxdgwwcz3
nK05p4gA8ONRQVBHc27Mbnd3F9AmiPvbnObIWoiCuzrmiQ+NkH6nl2xxGiOF9Xsd
Ux5m1DxYxPVu+HLcQwuIEQHv+rIE8xPo7EmImREAdH/kEfLtZgGFppzme+bAHDWy
ZPWX/ibGz2nb+kBfr9pPx/4G0vv9UlPy2a4ifXeJ8/1KbmMaZCYL6t1FzP5tGFgB
oaCReaAQWa+FLkD+AaAXRQZ7xm8P4acJaYAZLkV5/zgGJWQrLiNFCJjMQ3ztjGuE
MyJ085e/oa5rkQIqh+ppk94kqEHhFcmrKqHS7gcROJkYpXo06e6JAqkMwd7GiJkr
kTBWs7qdXMGMN6uxHouCTinEPTh0vRRhDFCGICn1TxHmL9ZjtMaA+dJMtIltbPzo
nsAfwBnZ+5AqxzZPIb/eNLasf2AEe80Z+K4LWFDnRcB38bNzuwdfDmSGB+0o2ldH
MUqZSgQyTWmpD263yrbRFwQnMLBXY2h7JSLoviKU4QhZ+WjBLGSJsa2JKXVpuHhb
A0XlyuTRFLeZFvKT6liHU9Te8UrCxUB9CnSTcgPozpj2gPwUKH47KWXedNDfL9vm
B0y4+tY2UO6kHjqqVs9FFvzb9pNM5dm0gcdGTUBGKdEXanoFLh9C3gFjZ1RuYhY5
kmmNJUnp9U3ae6MrcFUfiq8Ps8gPZ1FAxgIr52r+GbxrJHpZIJo8YRIvVMl7+p0X
10LQ5gtpDZtXhb8MVNLIASsVqAYkTZ6ydq71Ka6VFC10rAIWwp4PZ3QMssuWej+J
F09oAmAZcyJj1d54cA9eHFHXRDXBR/8hmnd/pN1vm8mmvHC3oVJjlteUC9sM0zeu
id+aDOV6DnZaclYpa7RH2Z6lcoYOtcb3ZCvd0lqHNRDDLG3x3gu7+9GJNjcCMSBw
JuWLh/lnKzvctqndDN5r4iucyq/QIhRn4FCEnGKClg0kCVDL2ecZbI3PL32TbHnE
dsM6DuEAWamdhYwLSTwXBF063qqS1VZk1fynl0nmgnyTDHn06pJpeMdOlaY/QZm3
5Mh5CPK0YHlYdbZ2Y/ObO93D3oVa/H2+DoPOiIZ+zYTLZEtn1zk8L0YJLFKnhvzO
Exsl/2LOcMhc1RhH0z/1/p8ef8PjLD1zN5ypeF96pFX9HkATej0bjugJPWRC4IEr
dk17Y+5+pkEtydv8xoWRDZzVDpkh0FwuYx9t1j2FUL4mPLyjrpi05NXRsL4dCg65
7og7AB0Sqr/wMdwyvX2SgFvaDhymaYj1x8aZTCILndGi+fJep0W/bX3KOwGfivRO
U0HUaWPtGCADijOLV8sXy14PGybf0Q63tin7NvF7MlcJoRFg1tNDiE5ZLQhHKuJa
cF492nXUtD8SJS4V2iftD+W5irFCwMx28Nky9KgPlGYGE/kaciavnA9DbQH6Ez9q
t2ekb8XP5P9j4o+Jl5iQ7JiYYAvoRZ1iAA56Hg4kKUq8Qa1Zuy+Nd1jJHKHinAP+
rh9fQ+rq01Py3RhJiQ6zH/Ttvqst2FeOd04vjvGEAG9oZ20hqh1xHuzinNyPZiTJ
MhBwcYSHaOqWtAF8CCLE+ZbMpZyhvv8lDl4GlSrm5OwvIMdbhys2y30vKhPg4la/
9IexZXG7sFG+4TU1NqtchttOe/nyjAK5/zFU/AWw4uSBb61ffZuZsdFC1mXjaFAO
jLDoCm9EIQjV1rueuhNz8RADyqtxoMk3HVvo5BZyQxtjDdUaqiAG49WyLs0z8GBD
406nMxCz6cMRZDmoayXFEaPMQH8U8wcNPQzBBXKxrvbzFTciCHqDMZSeaqp5KI1+
5duNbTqMk9ykV7YXwgwXfZ9VDG4BBG0HzZnFyGCKt0ENzmKETmhLxFMS4HgYEyjb
1labjGcV5ufpmF6sRpZX+LLbOjn0uLnJfqGHHLmXlBJIjRpQqM3pKpny4i2rzzRw
W3l6vfIU94GO5Xqr5OsOFYrcc64JAAJJqS1pZ6CIJOjRr9T6FD0Ap5zkaRyb4qyR
zUgQmk5IAXBLwCAvEt66ea9PPYN/T5q3wR3e8W1baM9kVjNZMFH750vwQFYTVXKt
IXRND395Mr+qbjg+4CJKmE/SeBRfslo5V3Y2FsmoKeNwo5SODnaOsF1gqMe1h96s
p4+CqA4UObuylQP/67++Viivb/jGu2FlrhdDPU20XKu5LxylLTLBtlFotwNZA3rV
wq/ikP8qutxz80pgsBPTo4rcN4iJy/Z4WX4EnAO+md5VyP/1S1ksV4lHwbB35T3+
73IEt739QEYyP8C+fFJsFVA5Jmk7Tz2oq4w9Q2LK7fj6WfKud2QRId4hNvZUkrCt
jfacNDkE6lmIqNv4E4BIgZx26YK1M8E5FkD2WQ+LmTMrQh3okQG8doGbzLgpL7DL
0+hh7Df0vnf7B1mFOvsxMaP4SezBG7OkHhfMt1fRJ8rlYaxVYQ+jueY8Vy6dlSRm
JuMGqHhTYB/USr3nMSVIqArQCXaNlSQK0+8KDQmSMKZ0vu/z6tK3X2mbWm+omlW8
sNtZKcn+JllRrE/W1MMMRH6pucUP1oQp8NqVW9b5UR/4BXx9xXoAPpuMC1gbgWe2
/2yMyM+INfJ034M1CkQpeLUSrTDj4JAh97ndcHZFxrii2R0yBWxBtKG4r4aUVwwv
8DMc9ZOADvBa861Upc32ZU01npT+U69pYgF5Q8qDB+s/CbN+GAlLoxIcjYPov60+
/pqilgmAxnkJ3eI6uWXUKI/rkt6eMubzwbH7cimegyk5qHtJ2+IZUoIpwQbH4tfk
EvLk75hkJyIwQk3VH12AryKGW/F3elVAcUNQJrLGKbNYGSed8QzOJkAklTa3rheY
J6yx6nabc+9sC50ZPS4QuS0ZXjQEM1F2xja9mSZOyvnPqqqlSpB9ATk0tUS59OVL
oCa1Vv3F3/ngH8kfKoCDyAfF4jJo3pCXG/J1M3veOanTvS7m5x+FgZYJlM1aWCP1
iN6nrVH3nVGFoQFarxQXKHiYbEQQLjUXac48l67rtlX0FYr0bcFn0zyxsldzEx8P
rOVasqlUItCtyIR+BUa5OtfLivytNUOiPuck2v9/yn4ZxT97g2HLOJbLN3vHII52
Wn/3pA1Tmx8n+7ql3pT+CfdUz7mWAJ9GwN+m6g66SjrNaylXudE9c1ReMjyvLH7i
IWFwVP4xyVEsKmE2bjJ+e7PCwqDo51s3jf37fTWfN+kKy8Ulv4uG+aae19B8dvP8
vNTRlXBqNeaEsJHsf7j3rhqs6AsHtPTZW5WVa0xWb76C3/fxZ90dPcnyIc8gTX11
3ODYueOp6gKtPgPQD+bjEVkJVxKklr8Bc61KLd/Kvf5DQ3CiqBBUG66x5n9ICc36
jIcVu5HjWpBUhc0b5pFeVE/0QgkHElQ0cOeOpIvOYV2M8VZsAbuFdRaXWrZ2s9eL
qrfrfiij5raMzF53HXV8SV2j917F5fr/wg5/7Fri/T0xLtjlKY9baLZM5566VvWK
kQvCOyopeASquxePOXQweRoDciNijaHX5oJ0Vp3HsDWZC8ExJHjpD06abXhsl4yL
4xQ3mxaoTr8zMPDJoxSc+xWjdLufL5C3LXb4FY8GyH982FOOfFmLO3Op3YgHuHOf
HyW+uOk1qWw9PzSLqMWlip57DXpkxQ1GbWg5gj5n66L8sQdzgKOi5whh32M4435B
kfWGmurRpRtQgLd0Mg3mbrxJGjx4l/njglR9BP1anaO9x3G+a+KNEJSb18LMav/J
BpSEPB4ccsz81VYJxQwVP5098/C9nhQcCJHMNtR4eY5VW7Sw7kWiY1JPApM9PhzE
X5M/fizS2Ch/LXiymviVCZx4tjvGcavVBLeeKcWofy0=
`protect end_protected
