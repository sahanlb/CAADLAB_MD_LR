-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ab/e6VY370lE0UERMzPzmCOnO0/T1BJzYvtDc82eWEiCNQirsVl++5ACQtQhanae89oMyoeauEQ6
audNwe3VBjbvGBTnEy9EzXJaGyqeE3/TEMG6LjAcI1GM13+ACNogjYKwvWJxhboFW1rCouFy2xE2
bm27q03vvJ1VG/7lgHHHujzorTGgVvfbLoVSzZrrogury8UqgoZJx1x1WKo7Cq4stQddxRbZz4iD
Qi5gst/rwf25kaXd7GKPOxPKVPEyM9oovG0DfAEKR7x1766y62OKpPkPWx3Zxs/kuitXE66vSjHp
e2iomEr0ZOi6les90MHH5QG+fVc0sga/TaQ8yg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5984)
`protect data_block
sS/LR6rXihjQEagBk2uBl+a9jnm8vI7IP0YK3dYyRkweTK+Y8rrCvcLUixtKYG7ftrRU5dqwxMMX
3ISKe1mklFW+SvZb4KcKJ0fYjmitLI9sDnv8GKz17zI0Y/BROcRPHzJI8tzLadZ5aP9enObTgLEZ
Dy/jQlY6qOBmhxXvfwbCAKytub3LDyzSbgUmU191dDxHoreL39aucsbd2oiIFfV8Mp0H/7QOcuiF
6S7XxKxgaBak+wzrj+2K6N9EtHbxXwnZpX/zRjWKJsE57wvhrRt9dYQ3p8s4MHVdtVMI3myb6uZ3
suIeejdzAPilHK+hO1sMpJt4vbVz/5iq5UWZ1XY4FolNBcYCyChquo5re/aIUTUccOJ4Ziwbi8Fn
M89lYZ319/+jlbjUE54Ayd9ukuVFjZ4xYkSaJskrlUayiiK8v1GZ5laE8pGfEYblM8JLiELjU+9R
XF2QhB4hSEfJCh02z+jlQCsTirV/mNiXJI8yVe3WEYz1WIYt7shkdZXWvFyHTqOzAn03efrYpZaY
/K1/Chm/lkuuY3+FCixurX/0e0rVL5Agz/6q1Kj5claqA6FVi6Z5CVHGQlW5zRniQUMFJH2kT6fx
p0Nku00VcF/qajns+zM7jMrRSWnSUjlRhYjfEH4CxZP7psgtN8dZK8PvVLibrxrhkX/Nr2dfOOd6
7Jy88cVspBjiKVgJHcnoK8Rrr76Y1namYWwqBKxg4t3A8pZb6bNXkcZhTc/M1bl+Gr/77wlCrtmM
cWfss68xssw6OFFcfa9akXv6dqf4eZ4IjEIIQFxcqO+YDBFeMWn7y4Cr/vdwMrsIsX8ecTI369Ei
VBDecVs958QWXDzneCBRCqkCTrfOObfSqzCYCtWokyLRI00fk1OI6lm2QDjZJ0QJyIzuuX4hd58x
ZQygUNbzszXTzAsubwvIy1x9Jp8GOvTRMdFW/OIJQQD8ti5Q7F0XlHKhys6WR4kGslzhXbFKbatw
raLLgYQGPybl1gtH3AJH34OwTaqtB+csFocyQ3W7BQmDQJyU0v0wWyG1Az/WZMmVFbvbIqS7gogA
/QtaxHzx3RG3mI2T5Bf1iz702kq2TgT7qIdB0utPfH74zHcLnaodgmB7aPb4RlFrRbCsQtQ/t+mD
LNDhAp+LAC4kO5r24Q5qR/w9FanjZdZF8EoGBL6plc4jOFDGEdho2eqRaZpjcc23BzU5MBhsVdQ6
PTziDrx8wna35ud14ByHyfP3GNBYs7o0QoFeqZGpbEkpJIXNxfq6EG9zFMphoVsjJWzJYyTWE2cU
y1cqLN0Hq4iP52Sl07ZCkm4zon/HureXXIlltauaFqK4Dc92pfxlLoKwt62zXN0OYPyuScVRCC78
anbxfsROL5LBsVHMeKT+TSZarGoSL3H0r5g7Vu8445zGbHYukfdY4OXKnvvBQnbnYUJrz1+7oydh
h9rJHGC/9dHuqlEPeNo2mlOuCzfXXT1YcANtLxpD4DzP9UxFdhMzAQfRSrX4U3rCM8CbIGPaF5uW
UUF/f+MMFJ+0htcRwU7AWCEgQTc8oDHdyll7ei/WhsgabwAuzOIx67qJEqcYqS8MKfazUg8IvJHj
OSuxMrdusIu3MkIF/huPHF3/NrXQUEilJAsNXHgRA2Ix+eTcKf61pc+4UkQ23djkW9Z0qjDU8Sdb
rH3ZPIovdiLoYH0yT2l13xg4ivzJI/eiw2CiNP6jRahKhyjcxNX/WVte2U96IJrkZIoKt+gJs96N
sY8xX3bDKqcWK8lNH4wPb3gDS7PxuPf0zkqgCKMJR5A4F//DJU9qKC7BynfDhmTvMBHEwou2NUFW
/jehx/f0LX7tfXUBIqeVnnDEuz9VSLfoxnJWJsxeRqeNwLHW2bM6UI/nOPGCBYh+zb/RUXFi+h4O
I+4hfrr2wB0HgOyx5+vqi4jG8I6ZtD2T1TP261uqiY8NfULXFUug/NqjDxtV3C8QZaEgPeOonD5j
/NzWU5ZFybni5V9tpJy1ap9Z3XnwxuWnKyqE6b7p99QPnbeNE6lhXnHchhkN6ddwHDsG+5AcLb9v
8Biqnbtbo73cjh2scaBB+qjeblRR/uKV3b9/SET9g+8knmSg4uMBZjZrSQMwSU/7NhRYlbZRISRt
/H3tk9ZyHx7XIADiQXlURvWo0EfXr8XlrYA83RFVH+2MH9W1X+UEPiuZCrKbvTPnsmvernsgOB2q
Gn+qwvQvABgmUVyBo/9W26Ker+w6AzOw8NHsQ+DlAiOdGYMFnUpmHviyvQTKgZf05fm1R5zQPzgu
FiQCmK6iT/QA839ki03QrTSMRCk7n7OAIV+x3/Bmir+OJUxiLnkMHzCNV1mfMdyoFIyyLBC+9HD5
dzR/TyAPrxnDiNjXmQoiPBjjsJ/dkTJgmx2u+jLUZengN1Yve1TXYd0480mf7OO6z7TIkl7HS77l
FESC9tS/njFGA8KY0v/XT+bTEkq08/6b07D0BA+Uoi5UYnWM5cIVi0mSg2gtlXbOXirOjdnAJHe0
yFBY7bm0ir3Mn4b2Ms9LSTWJ3O1FIAswHMkDevgJfmsYPzdO1uHvTmVzkpjsAM3exDDDGe/LmFla
NTToSexBk+MK0nn5cFotes07qVaMPptA/ERbqCH0wggz+bq/GesG0QHwCmQ6AdCjBg63ux3Yhlo/
FLw26Ly6jFJB8nCYPckdmQy0jv3mDi0czRry1QrghKQenZ4Dl2GoQYDgLsJjzK/a1UYF/jl2WGLQ
a1u7SV+j0HmCdZ92CkBe4xGaP8+GNzIHetZiuKoWV4Tp+Lx2sW7drowf90LuKk88NeZ52dARTStG
Q2yEfZ3XgHc04YSTQNIiRuSyM4gA93D/pLRclu1H3pX4CCLGVp8E8ot2A8mIx5VS6yHkG1JkAEyT
1Q5VgqG+es0oPRuSgsr9kFGQJkpN5GVRRRTpVQThi67X4nWNawAfqHkPuIS66+GVTfVMfPzJrDPH
63PaKgmEyLWR/9g36cU0qeLTHOfg7YCMrLrRTR6JZ/3tuhfswdx9uvQx/rZ6IE3IrMiShetWxoJs
erqs4X0cWPDi942xPPsiTAWC2WtbZ1AxzBYMao5o9fDpRL4eXSuH8wdLcoQZ3OmO421iF6B3oZmI
/tyXowDu6Vk9TCV47S1YUYpFpuUnIxGO5OIDFo9RBlvA4YX0/UnES69FMytQdfOGreCumeqqLMWX
Dl+ymE6Fc+5R+lTTvprUMtEhNFpC302z9zZjkvvrAhF4S2X+4OzUXBONyKKinhIJHxdF9qMtfQRs
ehP5bw1z6Z48o9nsa6BscUqymRWTly9n6cCUHcGYE7maaqSFcEWxNT22FBLK0wRQK7CJHgiThUUn
AAlmAlejfZ0BxgQDGZJ0dOMAB5BE+qncKAdrcoKiPqbMceZayLC5N8EsRlSmioslHseT0jlgizSE
k72Y9Kf3BwRzBXFIUUTCP/sm/lkLcimCAJfRreeG8TLElBVRu6JeIK9R1Ex42yrWks2j1QhIEScq
tvS8LAZ3giMBlh77+G6KTr25c6Y9KwHEszPiXDNDH9rzElBNyNjGW1C6rUJLvD+VTNV4bCj6MToV
Y3YPrn3utPX++kP2BJB/XB75aMflFWIGmj/9xTB+kSwwgoHQf5XRLWTwy3Xsingq3DAHZECbkW15
X/AMc/6SYrbcspB+dMKw50ZUTFfw12u2elkGyLYcM0oT4yqSvkHWKgWIbazxYdfpnEgMOt41W4mh
a6uTcq5QCivLwTdE0jWowbVDchx23QLWE1cyFmUDruCiiniVbF4C0IHLBgxI3xpT4XEhFPJ+8fbQ
Ml0yfUcJNqtrUtjt3TiTrSkpDTZCWWGT2xtDgFeEwy1rOVJRZiVKXTFe5GjPSP1Zns+F/HCjoheW
G8TCWsGlfBi4vcnMDmp469l1Yi5RSLUPbsxPiBefBdQm1qW7ONfZROKbiCzrAaOBuaAh3tQVzpx6
/MkZs2WtFVYL2uDq10/wlRie29+ICLZak4c4LRfc6Hzv9INJtQIcWS0DYwQtREcYrSpBiydiSRLi
GDUP+SZSkSqlmC6wp3MQ7p1FDWkGNylQoogX8VBX4H2u8k6z/IVrX6RJwvrbV4JTocF/NWG7xmy8
nFp/BDFEddh4Ydx40J433X16yASHjdhIVrozzUFNzMjPA/G7FSobMHeygFzZGldb7vrFBEQXi1El
HzfJsP3B9laP+tCEf40A0m1T7RGgQ/Kd3XF1VTgtqZKBN+qWPfAdHaILlGs9evjLyr/B4Z2A0j8x
+ps+cPLJabwyTZ/fm6frbEFHgHyz/bS26ZC3w1Psk0m0xEeOBVZ9Hi73mtj4JxzmvGAtf+vrdkSN
8FSZytCnqzv8N7DR5cGPAc/Janty/xgfIFYmaQgHbtoI8uaAKq9zVG2VBPxDrsbJXJmwfpy+rm0a
cu8/fIBKE1Bvy3/ImHmOqAaasP640mZTa1kR7Eb0/6YnWZ+jvrsYUaQQ+jy30kGldIzURfwxWm9+
fEeMXNr1RSp9ph0c8A5yjIscEbueU8YRCdHEzCDRF8EVqvA1hiGbfB00z/gi4M9aBPsov4JYMad8
usJeCWphkcIDecbLZVD7hskmYZpEtyb3LRgpPsoYhH0sGsSee/xYB3yn3+Cpx6MENh7aeoeuAREJ
1XhDP2UTaBRh6s2el2uFFCVFVu9UrkNUvlgXqZMVkpxzXsnd/pR5FltujmLbEU7LX+B2zEqAY0Cx
UeFTj73oBaOTnpalIeeAdJO/9AnIbpHQjYgBwfiYmZ/ywMo8F2bm/t3FnUR6TPRNL0+DhvGRncKW
OxKLdC1zxh17I4Yg8ZIz7a8uk9yhvx1KrBpLheTc7YrVdM7Won79Kl3S5Nuq/Jbjacb0J2QrCyIt
DnBU+3AwH9eGCK9wPYxdggt5OU1a7RgZIsRkXZvBJI7iZQhLlx/VSmTdl0j0adhVDXS+eTKphEk0
WM1agdJXKTtI8dVtpAc/7W08+ifZKyG3RJ0fuf3BsCdPgrzUW1zckNzxmCN6e0Xs9Ahzfr8h9Pu4
iAV+y6LlDNcgXNlNsAGC6Ok0x2i4v2AFAOfMKUIhcLHwLALLLiSClXanvIFiiDPgBwo8h3i9A7xK
AGoQttzD/GVOemomTTsu4tLjxKJTNym0BuE9gULg3U/cDCZ+h3FDrpTOJRzmRFj057sbq0pDCjjb
8WurfDBB8HjupKOJsDW5UZg0NJI1alZItau6tZp4Vz4DzwFzrmKyGWWyAX3eSRrFPXfy+7hpa2Oq
orh86MjNrU3bghsouLpDeRh2avvWPgxoddTvmhnoeEm1ysdTTP5AJX+dDiAWC7JMjeQx8IAB3JMp
ehUN54xRiUwrVFlcs9yD3gepDSXY8ZnA5QQxzIVLYiOj7B8Id24ioGoggOSN+hWilFQ61Za/KuRF
OtleDxWswzYtYGqTS11FpaVmbyrH7qvdteckqManY8GS/6rKLKSChBx4wJJlNM5SBTWvrw02u4Fa
5xXSlf5l+kWbPk8lLZI+eXS1L6NedSWPDgnJV6HAphZRqzUBnKqLfQG7/W2zS8yGL5Rebupa9WMg
enNBHbfTDTc6Y6QRAFI8B+5GDhOGB5HlrDWob63+EVtzbnxWV5QQbTCXc0xb5sgRh0KlsTwiRcTn
gaPaaMplwrDvIp/1QzxM4/VClSW9q/UzFRzF3gBvmeaMh9BWgMavKPeZ0GTlfa1eCR5XPUxRtY2b
jc94NXU0m+b4hTsS+6lFHRvibjkdGY6LSiuNrG/Rq9p8DE1Si3T+hKdiHKb15ZulTsFj/LTKjZl4
r3l6FRKIvRar4g2Uw0vyU7T+Mj+TJwxPpIWGIczNXPPJnvGmzv/o6/gCfGDvvjQK1Zn7M26dkqwP
I0p9hxxTISaaPHPEsIRTo/srnuJasK8AZXL7oLQY87jzf2hVWwvPyRwROA8dKZB5lfAIow6fqLe4
biMNzhvLzNhWQzmiBlDVRaASSJliGUAQ85dTJCrvwn4hm1QijmbC2W/qEl/5USNP/RukE/Kzjf9d
wQty6UuVC+s/WK3s30FISZCSjcXdQnGeRqeA/IGw+A4azzyAMlETx7ySU6h0NSnP3PZiwZYmhvQg
8mYS8HCgl3Nlu6I8GxHacuUks0bLcUDu+nl7/P/viVx5YSBHqA7tFk6aREjqJszdtcXc0sdWY+t+
1lJlJ/ruSQ92WiUCiJOs+AYT9hO8vnhhagQBmk4VxbSe8uCC8Ercj3akDjrlLFNYv/ezXUJ5e9vV
hdSTOBLO8PmpMIsHbvzlWlJ9pKpyqC6cREZ/kdTJWMQT1h9V8VhRCov77KckL6zEmBDK4WfUO17q
sm2OMyo6x1Kn1z86n+4yOm9vKYcoIhvd6+AFF2LCzckNBSFPoF05CoZK0G2JKFgulCUlEFuCTbOD
F6KfYG5D5lvHmlRLq5ITBxZF+ouhuJy0tTE8DcIw59R+p3+U6SuXrHy/ZFhJiAIDvqgB0NFGsGFz
i+h9rajDF3w08huVUdEJa8ocJUhCSJdJSrGnxxvGcH7Bm35BPkv76wmzljZWdmZEWjuOs24iwSyg
xckuXwHSWh1sdLPJN0euTrQvGTDGzVbqwNolLttZKbZeEdDk7toUsqHbJGDtXpT4xCOMH6evYdVC
x9Ugpv3kwVdtmR/AaX38dfrA+OXAJ8Fko+yl9s72/myqCVRJ+YTQOSDAIigbh720hL+VxrdF6TX7
fTRstr75NKelWJEKxTDmL3A+bOnMK5NjyaeUmVRviU36kzs4PhlygTuedK+sg20KuyA0m3cpwka9
cS3dtwg7R6N/7hyRTmTAYairwkIQDoa1c3IDSkTdz3Taj1AL18XnEyIC4CFC9I0CZ7IQxHXL2ibc
UaIu9tsSgkzN5gkSyiFUxG6PELeZKVpJoAaj+FKIg4prxms3MUe81MT1iO4KYKEQPoW4IxBEzKQY
bwQOUsiJ2F5zTGRKIaWk1paYHKBfAoySuizhmdQwjYnBQw2dAIG2cFE3yYvMHJbdYImlzMk9UhPP
WWEcvVnko2wcQQbSicxBLOFeKN0TIvi37/cTmkykquCH+pJu1bovWtgcpSwLaypy27Wz6Wnwzc8X
WO+2+nCDBlFBrYPBh1IC11lgd9bOHsg1ueQyYGAhlX4c0CYVi7p1Xbg0BgEcMmzQ7VQqdmddNnLR
ODWCVwlXzVShsmwqn0rw1UhCASoV7yxARM5koHe6FbeowwkTcrY9n+4I2lwj89/OwvXoCayiTOnS
+2x6Zyoi2EQYcm83GJUUL/J5VuARLLgbu2L71Y5hBij/FarHfHM82nlzMOUkweqCD8DJ+y7e/wmZ
Soh0nTyHZ1RfDWIHfYVS4qNGBg+Av40h6Z/yyE3KVM5Mf0Oa4qlj4cTuzBkRl9caAc93kSQ+YN49
XgmHbZImB4BjT+l/1raxy3wIetxOEqcqMbKuQWnrNOHq+DcJzYAWCtc2zAF17HyOTQSnRHiFcmxl
r0VWVRuq1lrZOOnIZrbyW3AZ8CMpHSswnzsLKZWgC9DuMFpTcps8NHBPJVIU/g0QM513yeDKBUAb
ZdUINmoLcEKvmIrVyKFKJZM0v/PyqZmYiSoE4F04epdORwLvqAPia5XlMMVwTxzIUYsmKv7xnzJp
t5iCs2H4siTx5vuQO/CKkZS5F42LrSsQiv306ZhrVdcswwWVzzszwTvp9wYy9D6V0uk/q99Kpco0
4SnQkkJhhEVMx0NzeK1JE/yECysba0lyzRmF5rNjp3Ndu3d6OOZVSR8y4XO+bXTfKtJkJqgb5y0E
cmheyMekOcgnmKYkOElKHrxEnaQLOniw8seJHpi18nFXY8kP39QEs4+kPzb2Qek3A9++fVf5u6KK
hXoHuvY77fO5LhSMt3j+qKGgrxKLk/Y6QHp8XDOPgZgcflk+Bwqyv9bdQ061NdXF/6Bl6CiQLYtm
6tR6WSZPP9ctNV6CsY7DTGYTNks8lK08kEkNFuWe7gBPZ1gzKb56Z/RuocS166BI6zWOIOebgYg=
`protect end_protected
