-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
JfTcKk6rcpp202RRTFFt3Mv/74xlDCT3BGjyhzojf3L0ETtACgtxRvfqFEVjTFv/
9Kc2F/k0H8KyZuiO1DnT5JCJreEN+H/UX0lKl+cLFLfj7lNR//fcP23g37Awg17S
rqQRrYt1PVoJQdUHq2FlEGLjevwWcsee5NmHAkrfMI0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5200)
`protect data_block
VIsWaAZYIXRjh+4METI0P2IckIn1UG0diaF1seQuogjZ3ondVlx/zlGoroSegeLR
ofA1qHRWH696XpejFTi7H3XyJRWbiYx/Q5O/uyylKuDfTMn8i6+IVcIk6LZjBUlU
ZKi0ObFHd+oWXpa4hq6Zwxd2ibNOow4r92PMCsCXUl0i6Nr6sUQFrGd2eFZl5gpJ
XPw92krW0JUSiTzLRD/fOeChJXSj6IJR94LgObOXDXa7bLjj5SSbXmpahhyonw80
Fy14nPct1ng90bZ+WQymb91y5ZQPMXs6U/oLwNO+Ar14ubeDYMojNnC0eXCPRjUh
CMZwgUaQPtJau6Hv7/ZsgR/NCzyfGDvVlQ1cwuTH2u5BYnNwfJdveJPhs4+9yqIy
LoSwtNHIV8jdC+TjFoVkDR3oAwdtXXkFf0hXJIWDiZvTHtFpdBizR/cSCrwctmsX
9/ZM4PoiEXc3GwsKQD3jnQRtNZTY2Tmag1hXyyWrF9IFod7/rGlafeLGzhwNeCoY
QxHA5XyHfse6VP7jafkh4Al+bydhf7jXTy4/i4Xq/I3HWHklsotR3izW2hXgWDwz
UEbgtSIZr5iP2poNMu7snVok1qj90KJ0nMyTtYzEiZ/At4LrTYatvY+VUY0XOrtb
nqoYhdcCMJL0DULM6OfmtjELVdlkcnslQ2ONg/7o9XwU+JgeYyO9Ce4XXZ252BG1
TZhYjWqILGnURP7YNHnETa5mJ3BUEkcOOx5bvRIK7juKRotK3BhHADYr6NI9xH0T
PIUvKWe3E2jJjDbCqiKkRliGgGcvF29Rk4Hz3hx6GNmGo0gwwfrfELH/9awpFQDP
ppf/AevQE6u5Y1vH4ckhNN3kH8J8YeZ93YNEaj0H31fUhLtMEv2KbrYW8D6JMmmW
36ndbTC0QyJOUq9GhNfR2C6oyJ64QojfS+bmebjCnyRHvs43FUeK/d8iNPLfVIVv
ihRvAVCD2KGe5m13wzpVB1zh7XX5jGbAhRqsyNYenzI/JLJK89GE1FJkC8G01SJE
RtoA7e3XkTx+kal6cbjLlXr96/Iptnr6Qcyb2gvk3JsAFaLYw5kJUZRsLVhFre2L
EMhJ51MH06xsM6luQe/ViuyrKwUW6ZO52eGxYtx7QhM6BSkiES2PXqt7PfqtZO9E
3uep5EzNK9nwj6pZmPDDysE64JPd7oYUuBUFwhjGx3sGUStwHLlgixjaqMcz5mON
dbq1lHqQHpjlonUgt4ekoMx59mzsSBza72+K0IwOVGGm/W18ua4kLcohwkin6OaT
WVu4z1OmP+2TxHQDrNNIIeVzAhXidGKa80hVKS4j5CVmUfOZqxAiaz5GkMtECKIf
ctpxmddPtPlD/Q2Tto/Plwz/5QDYiZjsuDLPPg/csDD7JyLOfxvnU6VGnITF8E9d
KZMtxaB7cNVlYSUoS767XAvUHrFd93XfYag3+cISKksCqYrIuWxVsdBUbkon6SOh
whQCRKnLwmeZ88S9JEvKReKS5j8lZ5oP3MDuqlVscW4F7CcIdk9GdHBOpnAIFzOL
oU7pbcSHhw9rbPg/E3z+YQ5tkrGBeEkmsOBlePeFPkhcGxu9Jlf305pOV7y3x1AJ
9iydzTZY8gjkbNtNxB1/aWA+a4v7N0Z8b8ZBoKjjzFjUs5S5B9f+1IThDLOrjZ9R
8eiws0+6AWM40Ucgs0VTjeC/9k9cqMLxzNz/lzpxC/b70858WHeORg/4jzp+WbmY
aL97mtRvhG0eBar+mUJmuRLrtscA9akrPZmIQtuoleKYbCbM9nbA71R6Y1OFepid
RxIR5xBRVCYb6quvqvMmRZRdhB+c7R7LSSYk4IfuyDF8WnG340uihFY5X1sXRYs3
iDbKIPWLTmCICcJZGdlbnRRmzav2RE8vThoE5l6Ify+pIMhz9XybbRc4He/uf8we
HrhTC/0i25fPQ6EN0/bCgXdIT95Tz0EZ/eZd0YsUMOStaRvtjWYiBc6PU0fWJuS7
etdDqM2KS/3w/fXwlDDpxoAx00zZsiB1NGKzXtnVfOmYgSfWuwiLDvj9ZSZD2+4W
+uZvzsye5rPlwFV5LoF3ps3gv5ZlX7ed0UyRWTbB3inOhL5hEtHv1xorm76z6rHV
jlWY5SVJyzsVwQ1v6Zhv5vMohtRutlO1T3nwiAN/a1RTzan3aVOrYL8YV+so8U6G
fdLljKvcHHL/g0WXKcUP+ahsYO4MSssnuBCNrSbOdAUyajqovMTO3mjr0pHJ6hcr
3c8WR6a0zEC5Al+JunCMUeR7hmJ+p9we7bIQUOlnWMaGlHQrw5BhqdyaTioKYlwe
6jpi16svw/bBr9QxoZYhlp3VRWmAlqAbNJrcCQzxmP6IFmBfEwD0qUCG/A+M3XHL
M7QSGyJgSO8jHq6SpSDKbfLh4HRNQPM546cOgnYzJTUvOUwrDiDcv3bih61iNGn9
sqKKwaSV9PG0YdMi7LcTd1XtDTjmkut5F0ucDfrYGCrwmOg7h/Za2FUwLK2hXzIx
CBxizhlPbRAUdASyevs/gQitMyvRXNGdjIz/IOjhO+sXJ6MfUL/5SCoPLOA895k4
8nCGAw3K4hbtXj6hsEittIgn9QjBGaK/Q1v3xqL7KRQy2dr8tOSbjwkKCk+ZqO7Y
fXITyHkhIAgKb8AhaZ+RB4iPUDfSQ8/KBTDX0UVdvoOyVvWx/Z1XQWiMr0qChreM
fHSsl9U5ObtQzF5XOQy8fDhw5bCeGZyIuD6XQctdxYe8eN0YJd01ePs7dqXl075d
zA58BCyrI0gZJeA31flzRsnH0PbTMpSm0oJeeFCvNP4IX+32XjJHFLMl73hsC6L7
JmUJSZzcKvXGVJWvmkeJOhR+KK/QYV3z07akb/parQ5rtIYq61EpAy0B14OPZp5K
c4nTj6pxhE23CRM9ezsN8xgBmBEOEzZkit9kTECuB3YVY0ULUnBMeK6u3hJ9TKXT
5BQCx3JnEE1bkosbKHoeiiSpH5ib6i+/TvfLZf7KFNDV8F8VM4gUSiNRFKOY/Lou
WEi0Bi27fcMQ5WcelLXFGJZrkhzdaMft7FuVjpOZ0BaPb6i5RlleVOQt7AYE1BFG
ybQggDvtvjKsK9NWIwrRmB0u0SOSVdod/dRWxYPl+QZDVCXE4AfGNaPPhLzwAszn
m9jy8OKyIU1PRahvchmwfYnkWxIyzEI5ZngkG9yhgEFfgOEFBVWZ4kIAGDcFsYC8
6aeNzf9eoAwmK/5r8ehyRDr8B3thApZzN0xWw86hG2ts7W+pberXFRufD4eU5+wa
Il9MLr6m5O9huUWoTrsbVoRmipYklCEIlctNYdpu1+sPqp3CRKKd+0Wvjt9ndjAB
nPqdtg9FJ/uNPPf15JQcDFeLMST9XF0cAy77VdafRTzrd7PkXQwikc3totU5yciG
dJI8xD+Ldw/O3EFzXhRjr+yHw6kp3/cH3w8m8Z7ApSFaU1g5ZYKMXs/JlWt9ywP9
N+kJFjKIGzlO8l1PupzNrwP6EkaMDfoT75C6BJncg9K4JwLXMu1teDBO2Zl0/0Ol
4KtcooU/HAMWZKSO0188MBWRJjeguzOdlm/E9jMhhh863+eN+iB1v4yoNh40r3Oh
Qax3tmpxAd8PP/j7c/+vpmYVVejOIbLzameRrSr5jqw5vVEqzDMHiIm1BZmHg0qH
97dX13szKTVwduejGmXghwpv2Zjog5ziz05ZQmYP20KFq/90hFJIaXu5OS2EdCF+
vKV103ODwZQ+g+1QqoEkC2xEg85lFCZw9OFUMRiyBtOYRuo6qG0zYsFZcw7z4irc
BtmIUPGORD/jwaNS2JTFsEvUGu6O4fTLp+04e6m1Bgwf0+qE95L0nsJLvb2BOa4n
nUXidaLGdMfXzPyk/KdcqmYB2AYO/1kiq3S8t8CIw/fJzUY+3anqWYmVqELs2vmS
wFkjFywWKXsrtBizdT6XhLJSBcwfZSc5WBRa2fPlMvXfK8lj/I1NhPoKksJDKVYP
lt2cyJik0+FYlj3Xopoy9NnidCO4BSQR0CIQq3lhLj27tQxxZe2Uz/cS57R8V+sL
a//9Dg3tTqV61Pfg9PfXFDGxJixMnIjPH2Z9cG8OyIH2KNMGNE9BbWMDGgAc1JTu
WpA8GgZw/9K59c9YigfrWpqKXmtsbIHw8vmKYTwvqLm2aKrDUmCu5OuOQGFgIfWZ
Hp8T+qEX+Jj8mnwgL6AY622VDXBe/izUX7pAE3jqQRGh0PlX3Hrdu2dIfKMEXTrp
DkkyfLQIRO51sCQRoBMag/h3Kvcnqwd9iPhGq8thZNcCp0qGtHSvv+kAd1xrDomD
fqG7UGnQqcX/DKU8lKY+jugt2Dy/7VVM7CfFX0HX9+Q8t5ew5t8jR37ZsTRyPW3Q
Hwsq405s/q0iHwoJfflVpwv2ltj4d8A+PbxmqdkeeOdf9SMgbqmp2s0i577ZfFtY
71TF49om/DjpH3ha18QsEq/urqvQz+hB+v5mgbwe02ToQyHSM2nZfLPKQeKDWZc3
akPYVxJZCN7qxx+WSVmJmNpTe2ihpRZJrv223BHMBFF6hapmiN2u79yCgZLuv97v
gAYbt/G6e0ecjmoM4Epn1i3aIkeRDYwbuPlUlsoXKGckj+H9oK61bgqvFbBi3NkC
nx8BM8PynR3c77fzmx3jcOKfQ5/gOvrfstejduRKFgSA48QkNdg7sTlJzw8w9rnU
E3kjVNM6qKw0oXF63IlERLx5WIxbURCisquKHOPd3C8NfDXk44Arb47KKH4xJM2a
XpAsDsiVD68Qd842aVU/V2FaU7M+MhGH1L0Jfg/b+ZMWG4JjBUfxfUms/9p4Gg1+
iMTO5krvMroWxq1Qm5AnMcC68ti2b3VMsp+xKKVFjt9HG6ZeFPyWZunJ6Xs+pihe
eJWfN+/8fxbeeTSnno9yulctf6c8i/Tog7bzhJjSdjYbkAvJ0PRRaYIuNOo0wrun
nG24bX2e3m1TaUEh7KHTCiAqQhhuf/oT2yarULouldTl43l1Tnn9y4EIUFU9hmt+
lwPBiA5777RRNtUy6OgS+KUgvJ7yxjyAzTqOTDfxAaqfAkoPDdPqh+vafpAaSO6E
NmFsrsqBwdbSk37AYxmHTt1cidNV5XJaKemJOPkIWc2cXvUCHODMdLPm/GQu/zTB
vwiKe+v+MrnGkohx9X1Wn3sMrBkanvadQ8S8USXZb7veGRNIuVVu4ZqNclbyGIU0
lA0180QmutQ/kOiNGD1HhXlGjbxnabLge689pAQUQkSTdZsTyRoK2UaBef64VstY
gNTGb6jq94A6MU1juM36Uj/A8LMGuRH5apB09yQlfw/lBe8890/onmUDWhRdnQL4
/91H28u/9vAMbrE1MDlAlTlTnFDNJ/BXKa49bPUrsk1wmNp9PBJQTzCVm9fPmiJc
3bMY47282lu60IoSPLFYLlhE4JEHI23Xw15y75njAjPBOBvrSlMrJPCF39LTJ/vv
z9ntirurwC+wc/DmFf+8Ju8NPf7rbHYDLzthGghjItV6WAP5SZueZ2kZndmdhN6Q
TyXQvJjrkC2TbKIvRFxjjuheLZ35TunAhWMlJZGUZgqzuV4mjS/AUlQ4Go3gED51
7S3wgozqnrg1SGy46fUPcGktTOYyJ51RpXqftJZHc2+lNB0Un34eoKvtYHQM19zu
2ycoT+OV7r62q/tT8DnrsMbwMWLGcvhDL13HWOs+YhRzvoDtO+t0PDc50o1JH2Ln
O6MBBC/0LezpV9xGA1XvZV2QveXbJ/K3cPuyXptY3g0FebN2QblLn/krOTmIQxiy
Jwbf7OfacPemlBjMeIcEFG2NGTnWwXdK26HF5lpZrLyGsSiIc2LHNcLqtUx0q7sJ
DbU0biQdQ1m1t1y/f6iKnvNjy+e5SgJUltc8D0+H0EDWE6fqW3Ee9kWgsNz8EoYw
MgD7g7VMiP+kN7zj0WucJhGQ7q7Vr3Y7VJ5+VhPCrW2GVgv/6YmQgJ0uAI7QGqFT
Xhe774Pmd1mC6eFpG4vowK7d5WmdsxyX5ITfj2u8nML+Xtd2leWN/HDeNDO6sidP
AmukMVSNMSRFGqyQa273ILAPtwAbA4lDHBHHXnwMYIKdmakUsH+QKsLUP/I9XRma
Pxp7n2I95ALzSW7I/cFEoO2qFXSHuxvpcj8RLU749U2l7W1o1P/UJ165Zcbjqn5v
G9ypc6r+vrIAhxaPszLFn1t1iLmIztkTkpjeXdjzHL1mU5S25da0BFbeqHOyqAJu
F7371IZ8vo73PUiBRg1SG/TPWVezZsi1BHAtjaLhpsW40lu8E9mZs/0NJWrnlyQQ
gIZmx4hmToL+kqW9n+3OdE9BrvV09Lafq4FpFXKMe0Xt2PZPQBPkDSih6nmhXxu9
yCkqIfoGrJKnutnDo0i0zNhp9BdZ1FQh+1Up7br4CIVcaZxH+l20VUTsoHEA8UMF
ZoslnbM2OFNnrF7GPbSwGj1Ak8J0i9LSc0o51MKK4+HLx41tqcC6r1Ea49wXAk3N
dWf4c7bRdvmi4H1se18nq3eaiQv8NHQmiLgSuDEQYOygsQSbcczgpywNZIcqLlN6
9FiQK6FaaZgn3VNnSr1Ckvnw2Fzf8WAWoGgXDSJfe0NXhF0wBADIUWANWdAWVpwf
ubIRVYoLe20N1sTAv0eTg6wC+8QX5VSKf9pXRU/AsTABCtVCvr5VTjC0xvrkpADG
skIhD8OX/QqFg0pdOaB/xDQgCTrVUfjqZ+LHYgGgLAnhFt6oMNandHj0hUkgvMmV
HGVOnQu6OArUlpaZNv9eTNs1NFfwhmAmEEag6wNuntfEA2u4aWZqO9ymnnKHVZ9C
IXzIleQZ3sVejZhYyT/b962Ls5vYmnHxLDwQ094db5RHapXyynaXcQzuDhNNtxJe
sVHmVANplXtsuXVUSPVfh8y6ZFUegnYRCj6GjbGOON4Atj2rbLPVSeynpn0a8kBR
3bayABhM9nJ5F8adf8I93A==
`protect end_protected
