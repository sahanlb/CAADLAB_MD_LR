-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
GegozqWDg1dY+S8B0r+OOrGYDAO7KGdzrMKNUw9udpMuRWqNbcjF9+YCn1ri3xkb
gWA4SUEQ3lxKmqyyoihJp/X7oAj7vWqete3iNAwTuTlnTtHHuTgp2PTJt33FDcaq
gfP+/2vIQ3X4iTftvD5UNNDwV8Wizlx1TOE0NC0qaqs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 17110)

`protect DATA_BLOCK
9aPFarPYftGpcJRDjsjJZTyqKG385oalqsmFUOWyVcvzEfG4s6xTyBF4P4M+Pb+7
xYCY1AAukDQygIVAxFBvDMqW+LqtC0TOCCYZ8HSZp8NasdqI+10u2JT7OV+QtNY9
NIw33EnX8rDSR3xn6lv4lZwaTQOin20kOqrmucFE6n4ai8s7Ak2axzzjmqvuRQdw
VmS2tbw1SB7URddyiny7s39QYZEF6MUKvLJRGktQOmO0DqT4b3a7FS5XBWFJ2i3a
9dkFufJXkvAY04sOJeYgchA8qC1mHt0t+S7D6UVNv6Yh9I1HZI+laxH2/Bt2M8gN
VYYRNJlw946R3FWmNzIQSsl4rrGNovxWKE9SgxZKyIxEI2mtQFC4N8zIHYQ0NWFm
7UFS4fs57e++idFaRPlpG8sE3eh9T+M5c0GSavKJuqh9pklgtnl5X/IKHXG5ZT6l
4v0SHtsaO8WP7MBRr0yqU1FNAlviGgDuIKkzEQdMsHRYVNuxZKx4qLLzzCddaqRK
k9nxoMdzFSmmvK5knXfTLQ8QT19p3Gy2apftDd+SoA4Hl1w+itStUE8stqMObZV9
b52lWPHegc0fy2+LbJ60iWnmN8kTGRBO+VLb8qxw9AStAziakunslilcdJAHvsmd
SRkVYa0ibDFgP2kuHvwVzSjtjncf4UuDQcbwfmZl0Seo6zm5PuCiCJazgtp6e8Ry
n6PTh0B8d9a8r4HP1laghdY3UQrqIIjqNSuumz6f5cq/RApCWzel8HKxARcohKka
Y5/Npl/1B0xjqFK9tzgRgTq6ycluZ1rOWgwUiQ4ywZSmISg/T54YBLDBWAuEwRB4
0sq7dqfoELAPmx1X43o4yQY5hrD5suDA8PZ2RE0UCf3G9Fu8Wbv4IyvceQvbDrO5
C/aRzqxiegMDKHOint/LeluNMMvSGB23ioleaUR95VWGB00tEwFBgkiUDZST/Gxr
k9cACr/7UjlpbpDbkytFUAdzgSbjbrYipXf3UZoHjWe4nIri7MT2Ekxuhpj4iXW1
y2WYWbiFC3rxDiz99FO05IXX8nDzJQDadmcacZy4fdW0TpNnpMYAe7Oy/J+Msj66
3QljH3euvVWPk4MBk8ZdRUpBcQ7NTfOQerWck/Dcr4q9cAr4AQkwBc0bek5wNBxF
DGxodU/a3QFxER9q4rO2EGtIaaSvRrtxvE+r+FaaTmC5K2xEtb2x/2V8pzFsO49l
t4KOml9oie5MfyP03iDj4TIlWPwXFDWusbWHlJ/jk74LHUDjcEQWW2WCrhqForxW
YGba7/rvQWJ9fnVmJB50e1wIDK1Qbu7v+/2Y1pUeYrO21QepRROCScrIqioXBu0h
lKVvGhfg1BmU5ZsyeLmNHcKrRDu2jFfCfAnnjJi1BYYlKxD0pE3t62WUhX0xWtdG
cUJD9nznV9ygX+ma7R6tIFkE0TJ03DfX2fS1h560/yqHtc4SrPUUYU2pxgCPcmnI
N6w2mOnWQcpRynm1yDwSgFTgRR5JgHQf5Jwva0aoKNdQk4DrRfgAWQebxFq4CCi9
neUcXRVeUnrD3/gI9YfSNvRszSiqF4oqpvl3MQrjOjW9x3yAJL1LtEoxN59M4mQs
1EY/YHDXxA1a1LOGZpQMflJgy2J3TSuvt9W92I9XWhLmxNUTYIQDQL9SRmPXrtIt
/qVVlEFLSRfvULm/NrmTdfB0tIS0Ff2pMIMt7xYPx14bu8T6Nm3EMnw4uFGiGlr8
JbgyLrdUNnn7gRlsPXWKJUFZV6Vx2YogYPSKztUNvKssO5St9RKDTNW9qA0GXH2M
xZFI+f/Dy5t3bJEmcOHBxavEk8dFEV23/lFuC0jh8kOqCsd/MRcrIvkVRQpQ2PxQ
AWPejri7bgYTbN03SBNo9OhevYBDBwXO+hGgTCZ9nfoedvvf7MXYpHkXIrFwE2iF
B8YfjrqwZqK0N0ckL8HTIXT0FiQQNYxl4JJNArnifK+T3X78GDqEaSw6sd17eUbV
ZfoFRTZlrssgLVnDFKrf+tNWomQr5eHq1PrxiGeEeHprFVIivcchytlSp5tlSv/0
BGgBkzdOqXUEs+JYt38+BerYNNxONPDQxwOnMKlz2SC+5D4cDk+brX1Dv+OaquX5
ljzraAnRKw15aoyknx3bVdSxIgx83cLadkdb4D6UcAjvBdUtm+tpTMoKVJeLufw6
Q2+XWyva9m1oEKhP1bB8J75wh1rTMtFsViHHi4yxgMW/b8SmFpx8qbY3Sw03e+Sl
2NXc4q8zO1JuYUXXUGuJ33bEbasjuBPBm8KHl1lhWj+D0rTGzDIHrwMtqLP7Qphf
V/vSLvo1n7YoqN5dks1aoM6XXm0dgqjUMtfL1TtvR/4QN8lGVMeSQuyQ5/g8NNSx
qcCDonF4eFuNG3une3aL/h3L0MQlymkZK2MUiBMdT6xui/JchBld/Htt3cBAy/Uj
1Va2TiN4HZsuhKvVfRr/uBzp+tCDQZpOr3HQNHqKVWhZ0+ebWD2LYBMGf8AQ7lKE
U1j5wnhZIG13wQBSSRqaf8gAdKwk50TpbuARhKTiQbWgPIUhPdlrpaCHGY7y5sOL
W66D6rPoruKETDSxDeFlYJ0Ei7uswCjJrhVuq8cntVSrnsWFGXmXAdbd2sruvKq8
USyrGZJ9JjHoN0ZHlFtWR5BX4eZQyAVeOGeKkKdj8RfWhG7Lg5UFom93+v4yWasb
sTqV5G2LH2pAVEypFAwscg2pWKALDuoWSK4V4hjxYLdZJ/gpL47sG0hDLGAtV7OU
sBtAZf8Oo77snqHAnOTME0mCFPxB0L14AVICYjBZj9WNBn09eMaJnttxLzaBjaUy
TnlnnbQiSYOxAhlfMAyLV6a3JLg1DVLxX4cqZGtQppK/4yB8f7M/u3xy9qbaHG8E
yfE7JK1WcW/oRvFgUNOe7ww4N/2IiUztNFzYyrr/7AlTjqxMDSOj8nisJTuop4Oe
YMwB+MJH/pyEg3GmyEEle5HDLJyScj9FJVa0J4vEUDydPUlW50rldKSZi82C3RZx
/SX3dtg923083IUIIGtzTWQPd5nxKt8aWEXCoMPAQX9r5rpUBQt50JtOAZGbvLUt
xPdqFyTT0Bq2lGHgxT9S9v+IfK4DPYZJsWrtF0TzPndaLEiJ42Db2CwgUKRH7O0l
DbpXLHcyjLTfJQPWkMvAvjiThggB0eLWnTmufsS/DZ/rUJZCQjhBQMMTJCdy0Wbi
9v/dNyYbBt08LEjCOzWFHoR0APX6Co+tJVJ47uJo/zPvmgW1auspJTgbbbRFqDJ4
JKFdDvnP+WJgXdd/j6QosTUC3jmTF8FL2+9PP3Td+opSeJ+VGLS1y6MFOsFmQmG/
84pNpejwEv5leX+r3UKgnIT8n4Xb9Od+IbFuXD4AB6WJc1Voj6wxi90fdFukiZVc
Ygue4wOLEMHES5Vv/u6TR5vbjXjf1dYVuWrTa6ltlX6AmZ1IIbM2pTVthI9wKQe/
kDRcdMoAxfHpB9o3x1cCQ1lvhHxqTj+s4TkhgI49ze9TdlTvUM6+TbV9DlZHkXTV
GnwpWUc0YR5ONj2/Lvs5ly8cJYA/SHaI1Xt2WhZPvaA3m/2vtdQyaOERblp4FDZJ
SVjCwctbzgGQcykUe0zZ9lfWDVdT9DULDHWLmicBXCz0sEzYXbZ5ekj9sdyERi05
ne2F/v+b/x3yZms40kQWwg8igy5vMZqlN8V+RnQXz2GPSToq6An1r2EuRTAyxVTG
rvvVbs5cmlDDUJRnz6WLrqURmd9zA/fyCIhNn3TzNTA0t2Wsp7TeQRAdx/K6Fcvk
Mr750Gfn7NIr3IPxqfsVB2b2hxNWn5LyhaiU3EBh708TrVeXdJu6Pm8Tqr/feU9b
g/+u5pEpV5gtAZkxJMrEd5RYRWV4pEaCK3+GGZb2/28uM3Pcyu0f8sOfwPpPIQbL
5S7TvQh6Gv05OXqSlou9G8NQw0piR7/UsQkc6k6+Mn/DTVD6VG4Bt9x0rP3uUfdT
IwuYTeUH5KCwEml/zZpN4+6+ILPubs8eZ6cAczfzu4wu6kwcA+slyBufoMNkebhJ
1pFf781Yy15aveVMgt10YABwu0PxTDslni1u0iFIDqaxp1v05Pu47x+TFLow7OQk
yLBMY6P09htrMFnIKppM/UiGJFPSO3HNYqSiJcCj1uYrEI+uIksRVv+eJav2Isvz
y1wEhSj5GzkwlN+c224Fq7dGPrXjinkMv17HVe+T7cRVYV7rq/UGlDvjhieimtMr
io4qwvwyoHRIrzvbskGOgDY0SKLHLbcGcno1X8HCxvck3syCYaxZwRSjbss3fkEE
K/Q3TTQaclIZehhRJyWech+L7RrTQ+lKi/AXcDywAF+KTWv/0+BGhHS/oLQ0+oMK
bDngmrpcH4FRyZ5zd+oGOJk0CTPDeLCWfhFfECa4AA6H8kAzogJiorFTWypVfk3D
TEZbBlg//sLSFpcyVGiuZao19XZ6atMbSJjBBn4vCe3jObRcI6ZBnSVwAXGInC6/
fNpnjqrhkOhdCy15oKQm6QeDJkdRhZqvKnUDmOMMkvCM58KBIpLoKwvhiTQG35IG
ZmFpiPqJ+MsKI1DAjA5uhpbzsh9Pz+qT8HgT4eyYndV/HEPF2cLhI5gotjpZy3fA
m2w6r4xR6j/dI/qbtkoCN5I8aOFvmbUmqvPRDcs9NsVmbWtluPLQGc3vvLW27RB0
jDArgVd9W6ko33M3UB9+xfB2XKK/0vlMtHhfZVs6g2rmcQMB0BORBgDx9J7gk4hl
RynR46rR8DW5rnWTHa1OV5LtwS5NlJXFZzuEbgI5QGkea7XuDQVYg00LBjB2osos
L27+2y6jd/ON5ynzJR+iC4UOjwGhit4Ax8hLqm7XSN2LZTuziC8riBNNYrwKEegL
g2xdtrbuv6wIu00y5RK96tGzdK6LaIS9el/RpkgUj/IRVSGuE39/yFZLRmEsXSP7
0DcQsXWrjxQm5P+COc2n14xyEJHSLTQzdYrNT9Dhfeuu8TZZ5VHi4sJ7O90WFgXt
btDGw1MQFugxFs79tvxayBQA1UP7+N6ZLM4MBFoESWpSr9qv64R/tGbgbYHvHdIw
ZL9BfVaAH8ZQCOPzmDG7X2w4Ju5naaCY0kwrJn7yPdoAk0lOq6pEuxHCVg4eZL5p
xnHv+zmDqVAHztn4Ux5QiEwAifd9v25AG9nnwEgIboh5XjAxNEidGYXznkkhSG43
o4ayh12iH7AsgxOlDhX2ysBhzsFZlEKsHgLplDDJVMu+wYX/7IQpQOWQCfmvfNDy
dm6yq1hW+s13YTDSG34Kzemz9InGkV6mVxsQcBg72vR66N1Eoe3lYA44DuzFTwNu
6/weaPx29b5eFUkvzlj5JRkQAQKDIb/w0/22E5HSWZlunGEPuaCcRNGZOz850Ofo
S+ugBPj7nGAouKByv7h9niOkj+tXCrAxtOW8yxNXGSSCMLavLC6XV9NRPwwi3DTV
N6MXXQkMo4hNPvGzvXqs22wkNR8DYrYF097nqo6KKiIdG35i1F5KZm3XmM2qgvob
ruZL/UzGmItaSjgNcWTUi0hZYs/gjr5goR+xmbKKe1z9Pkqr0HxL2YY6VWSgDjxM
nQBP3ZscW5Lg6D7jXKcPXET+LpudiKHf9k/iC7PYTl1E3ysxvqiYJBvFksPKhARL
fWXqNZF/CC2X/uAxaWZ2jKJ/HH5YSZV6z/fbvqKszpbCn9XJ9QF/K8FGwGZ3sDot
aagfS1gWUCmC2hpEe+aGcZYY5EAR/AkWbc2T+JJ4ruV/+qCOBONJKe8T2VwrM7F1
011xBBsqT9wRUr3V7Ig06y+YqLlbw/bIOgM/JfbU33YrJvYtFewgKb/liIh5Fr5A
bb7YMalhS4C+u4/66rgEQbgXo6YntjMFHfA9SGF/DmgCr4RHm7VpjBQnzl/GFkES
Tqi7s3mBP/glsP/IlYzsGVgxV8e3h1EQmKATYx/GIxrOtOlJ5hgFCflp7egX5ogk
eVdYw2PljyDYPtnqzdssvM3KTrhiO5/+BjEIvyZmTr0c3LJyVYQXmTR99UqgP+7G
OVcf5wXEk4+QfYIga/c4nfxREZ1CSqrTItIGsZh3xkdnAkUweriB2mGReZQ4b7Ra
omBZO1acs8oQJ66BTIK64bmo80N+rAASr8Db+0Afij72FC7tXwQ0q1DsUYaFirRH
WmZivasXT+aAxgKydaadbSGY8QvJu49QZvTeSf7Q/7FCZNjad27x18O/WhTlHhHW
fWshSs8X1V+a/4RYVo4GQ/l6DzO8OQ6Gs0aRvtODkjL+HV9gKIneSIEdXXlHpius
CVbrCHwJQWcAu7vSyjeVUcbji8QI2Ti6jHWZehXX7gQZer76NDSBhyl2E/vXsHUf
OERmJQm8/fdaaxvKvIvzz1HjqO7jKv39KMvJuO95k3Dskx2xYBcYJarvlGjv+w+F
s0RtEZ/VvPmWp68G1lt/uA62vhKKCuf6IdxiXS8zsKDEU9SqvMqcByDKlyNJDVvv
tHfbn0MpYF3isNfsLMN00fMi2+cv8/nIKzxuBvXbpHJW8Lqr15cSS5ZXbcxSdyGu
cvvPTEKltQXb3vQlkbZXwOSSK3spd/SX/kA8q+E1lhcu8UJpcOMUj2wecLuH19EZ
KbliUVXQWahcCBwOzrEAgaW3gDcaGVcOlQ+3s8WXld9ubftxp29gd/KRItGqRVPN
ZR1If5lA+Tn7RJM9V7IVOPGy3qPDeQd02X4A6Q98a79qcKQqOSc8Q52223Uv4Kni
Fj9rCrOx5Ej4XtmxdRKtLnaujJIvg18rMQGpMcE3YaDFI1DmwRgtdenecJk2qQUJ
vd6/4D15rQSBu2T0FHfSg6PvUhaQvkIVgkAqjwOqwcQObFVchq+ZBUguLgAjghlm
/t5CnRt3xVPNuvY56VF5KF+cI/08lNYG8lY1adFpWt4H7C5+UMzLTmA52tP+WZM0
y7nJL1kL4PrdI8qwM2hqFGONLnrolK1QTGMA1esKC50kO4PUX6+nsypvSizrHUC3
0vqy4gxu6w1qe5d9LyfUD10x5SlhajCUgtYcGun3QUi0v/OqNuikZwhgYd/PFc58
/vgO/jmUdvm+BcF5j0HOb657kCVXFIoJ3zsbOFxgTQ8KYZDKAUZ1EjnPp/3fmMV+
lHlGGDdUErS/lYT/B0ZYAZZPBq/T55IDPr5QtM4Czu/LCF2WW4P6M/4H6h6orlhE
aWlao7dsHM71HPxI/XkJvw1NueJbnySHGyyLoMn6Vdf/T680cOtQbEK6ECKmRUXM
JpHf/Jb+F1MO4aD3NGfNMuIqodHgzu/zNPst+qXRmwNH07TY3ZuvboMERW3BHAWs
GB5Q3+khM6JWP4MTMwPXZXnrxIFpSAcnBXXBUaTbv9HdvlnzbfoTpVmibISXc0+j
bLPi7prPquOYmGGtP3b9eg8LiGxwr09aTQBgtZPkgIq1pTDo3d8k8fHt3rAuaMLi
l9hJ5tAUO84/nxwIhZFyH4xBb2CuZJqx3nG8h3QAMWNSE5lmJiEl0mbkO452Wrhw
UYX4Y7sHshlPoWBWyy3OCiPHkXdakBGccruSiSNPtlrvTaGDj4DLFqrzZVST94B+
gJoApwkx3e3IY8Qg8CLNoRpnW1DntSNp8qk2ZAdZZkO2y29AWR36p6vsCUu1tuqm
pDrcwn9doSwLkvINcQywVZgQQ1dXwX+7qFOxJQ0ckeKLz8Ul0OOAvGzsyq2KIAbC
ru+7NhzV1//wWFbWrEZ5kEiJIVTzy8OLyGDlEtLxBbuO2nuLc5lu8u6G4Veaqmjp
mUV8jv39l3I3KX69xsIgYKGriuT9wymTnxZGOhGn4vwHImEiuTF47IvN8vZDahWs
zHX1AsrhsbNrWTG3BY1wWjTBwH2IQfGjAX5UXykV40YWbuM/xfNeWpmRXEHkcebY
35OQxOjDqSpbXKzK++CMn9XfBtFeRM4OHviK9SoKYk6w8Vsp3U6RsXjL+8LG8bDk
sWwfk4qmi2rrDfiyayetwon994t6J0foVwaXRcT6Y7DY8lxSNHYa28LqXTnkFW9m
r3Wsy49M1NXShAFcM4kZZIhokfjWIh2HQIJBNced2Zkhnv+Rkj2DiXs8o7hmrssO
bBJf4D1dYoYRCBw6Ny/yzyQZaSoUbx0B30XO+kXGS7vSHGhmzW6hJof+bxH/GScD
1BfB2g5UlCsmbxWYBosdJOWaomewOo179S9ZtBOxLvZtDVjC98KPoSnchxzojpIJ
J43l61YeRXhRry8NPyGrIu1qdDQvZgdRY5F1QtNy0Ue1M0t0VFKXF9rnU1oq3j5N
sTX9Wir7BJnvV5uaIQ5E23kqgkqvjeQEMhXGtLVHhzwJK/wl1k7HCZX4NbhBeo9m
RxrPu5kZnFy6Pu+5M1LQcaYmmjnHRdFGB7nsB0yR2nPM5SZUU0gcYiFTFZldV8g7
WVdzt04rTulDJQRFzJn94NhY8xY9p7TIKZuygM9cyD3WQOTzjQB0lo1CAQG47CzR
SrVHlGdxsyfrzwnua69rJhk91VF2RIdKb6Iog8N6QLX3CbcSiu32gLJx3TfbqrPU
AIOL44OtNM8ZpwRXkJtnMvYjNEtGuUBtuwC0DeMCrMarIwKjMWTG/Gk5FLW/hQP1
sldmBCOi5EZl+D8HXFWDGQeZmROgPhNZNoai4UcnEMvLOAuENYsgKUetmyzHu9iG
g0FCe05UH2y2y/U2mIMY5yldqxmYHK7Rkjd0cHASpBpiW8LGxDZI2LrwekLqEqng
8AQqVMqWO2DgUQaQFZByeB/bCT1Kkre+CAHp/A59mOeI1mFhCEzDTD46Ki9ESGBW
z2HPm34CMG0M4uydYckrmxqEd7DHcv4sJxst3B15Aq7nuiQ+MUMhrS2mKd5qazbg
s+NHBxfgAKNA9/+WZUl+r8JetViXihTqL7f5cZYyDe28taBUFbRHLLQEOnK2i/bB
4d2MO6LoTnq6w8yw9QZwe25zVznaxLC2oRUnDPlxXZJH2n4dDWPBJ5GnveJdxVYa
jLTgCplE4EIbNVv340xKLf9C3TVBzXSVBmi4RIhjRSPKa11sVsKJ5CVjAgiQM8Z1
oPhtdROj7w71f3gVlHVxjS+DREAgfmKG0C8kF4UncPLie3sUwpPR2VyZavOs9Swk
sSwdVTqOkQnRvUEo+F2ye5x/K5jWs4U/X/tVHCAydMEIlBmVyeBqsDTtE2eMpvls
syfT4iXn8wiqgIAiCYD5KXsxfzu395xeN0Rkm8bbQBOgAozNrie12reWqCrloFWP
wbpixftgD9tccTvPpC3FN0F6Az0oRhdpuSYs3uZaOA56OEmqibk3tzqxCpDqDehN
0YRfMBQcQzXau3Fs9Rp2AUS8IABdw1p2ULfC7scCp67zT/PjU/Ta8uzDb+6m0t70
yK4tSYPfQN/5ys0uaDMMGx20Udn7/8TC2HpwYqscp2nkuC7w9/3GBetHlcDiVL+y
lMp+FCO3x1mT6kM5zW9e/uV5JL+dm7nzFja3FKcHVLo6+pm1LFZgnFgjPY05MTRI
+AtpOhHEWWSJ4YkadZ6q/x3zKKghxGbJ8HNGdN1NBkyTQLIP30vMz6f6+5hNpV4S
uDru9zZTfMOd7WipbmkkJj1r3Ge5CirNQcz3j8rnPJHxVUV1kXJQ+Y5UuY7c6qXL
uOCyzgsrrbjvtAD0CmlI6m7apLHtkU4mP92p/KS27fBrbxnLOOVA1M7GZ2DpEEAq
QFch/6vgFv2RBD1SR3+TatKwc01/iNLAoIMJcePET2UmW66QgtLh+c9AVpLXQu7k
U21mFB7Z5Lctuc1uOKGob/FTjcikxIxiEmOHQpBwqRggMbHRNLjP0hpuKySYzmPL
93ygneQMnkOcsno/GQOfSm5oj5O1Zhu6HkegyV1n7HaPGhqGfIvP/NdbIi/hVXPp
fhHbKlb/LDxYOnt9Mxe6/V4rKmZq+yuQVio4jXlyPcXUgMpL43IABzexJqj9EQxV
HCLzk1m2q2WQQhDLTzADSi6WES48zXb9GGU7RKU1QarLk1FqfeiciVt+TWy5KxEc
4oB0EZ1a9nnMb4H30uAsMRAF4I8SlSKHUsUjKD1+XfpiJiETvwP/ld4PDQCm4D95
RB7G3L59oXJvvYf+TGV6bNhoXR1ntAwWCc1TcMZg0gp7eyOP2jGttAt08dHVvSaE
NS+Fy2IkS10q21minDe3hZwQ/m7wO41VYNzxqt/qFDPFit7Fww6SS2GmmhdazAZ+
cXtJCL3qZSsE1v9fzN8aZ/sD/5lgPx9nBx6NgxgHo2XK+6sQFHIajYdGazdmBABC
sLGz1pnJwy7q8kiTh50sbrjG5mm1hkwEE7QeYmavI880cq77gleMY/nRDjWZ9FPA
pcXw7CFDGZ3GlUEkXcs9zO2QlbSU8RXPw83Lcc1Fk5NwXW6RSZTQ5fxiJFnACpMe
3kjAYD3Rz8FRLiBLMYKaKFwhFND7/IWRz7v9cpzD0KEdvRcrKsHW/NyRn35WuO3F
u6D4XSTUkeTu+eyXdXNgjSH6b6NTx/Ft5Mye6qof0cA5TLRyWwOXWbvdBHzHy5rJ
Znl0e9f4Uq0ALPhYxDMQC4G2OysAE+2DVGd+VvzLjMt4sGxbSXswOL6tdQ3cI6GD
4LtGZxqP7aIdiMrhiX/cLDkQB1iFO3c4cqIMB4v+L1zBKo3ETnA27BEnZ8JaHfp3
DnXDvHnLegkGB911NpadkjM0aCUMSqBdSn2JOANtw8auFrksG7CQOXsl8ciceH5X
22cYBYFDb9cKzizRmiU2G+Xvg9mk903SoaEfp5/pi5JZcdewBRaZDeddxCJjW6eX
KIfNGF3H/MD1+weMgWMe9U7WuL3K3loc76kM971sId756ybZkpnokokUyQivU9Ga
Y6hLbKirLDxAFSDGc2MjIPnUOC0vnOarQQT1FYL5sRR8ZiQnoG45Ox7QwoWPQrCM
tDvFvwfGC5Y5bIe954u30YYe/Td6X7rat+oJlBGat2qmX5NrvZpVt5iKJadApTkU
LE5Ca8iVgpaCoFW1lbtwHVZBBLzpCXndOtwQp/X03oFKTXou2U/rzzFSxwPv5giC
d4WNscEQ0O5WxNoIbXZ5FLx30KewbyxhBIYquZpFgINnIM2viFNnzysvrumcp+hZ
ym7b7/yiEPPeiDHL93HxG4I7HaNS6cxdqtGxTtNkX/lV6HVceRGYFBGSJlGOVEkm
4MrYi5a93PyIe5shyZ3thU5ok5Q7SyGzI+dhLsSaMBIQROvS2DpnsDF6jhEWceZO
KqsAUhYse0bwKdvHXdG43Oanrv/25ZNSU71YBOzotHprPUjy/CdHrkM7ubidEY05
tlrsH3UHu22Co9Mu1d5Pqw6SZB5oiY6Jh/sxz8SHm8cOKIceNuNfMmgjlsJGLlAL
RvaFbqDTQUrniDHDuEUveW55tdcXOjnx+2LIiT8+Wh08CPaZjNUOrKcXhP7y3hUI
3sG6d7/z+trRQPb+fMtFheScBcxFRZcy3/aw6PQe9nJ4OpWn2hUgbfIoIMUjQt7D
4DXzxKbqkx9T9wFQg4bwrcbNP7U6FV2BjbEUGC/Y9BRRpHzf4ZDoa43yscTAhKpN
kWx7M2cAaD206llX76rbup618azUZNZpv+E7EvWeMQ61QnLcA2RzWZ+AfY6nkEUS
6RRw1n6skXQtm1IpAOnlKK9fmWCdB3jA0+PWWvxJkttYKEG30AoymxVlpgutA9MB
cPUuVzer1oQYI9hnecN7yXPUxnn59Ul96Tr7T4Mj4KJwySwOFcMR/LTKX/s9eMKL
9lS6o9+HBnUh8VmddAaPPsvSNagXmzEx6H5e5SFQOt6dmr5VoRhV/yKUaqGEeL31
r0Q0L5O+EuKhzlVkTnKd9ij8kNLpf4IyBCI26YWIEQEHockQITj69Fj32gYeYne4
AUFIzetoBtekb8q3HIUulI80WcO2sPeohMQ2gsXtPLgVvLwcvfYBxT4MIPspuhQK
MLgJqwDW6UlMXzH6rIJxLH/qkbmWef+DfldZJnxTFv0KVGu6qLfuoLPjWdAYpbUy
wnp6fv0w4G0MoEnSutzvAuYlBuLDiF+ga9HosT4jqcP5qCMV4pbbPPVqlMG7oJlf
JsSKd2XKCPmNwfhztCgYwTOEB2NN4XXQKKqiJclGCAD4MxUK/k4XafnGPPpWmcvP
JRxLbsI/Fg+YFuScal89yFvfYN6Y7le8Y2I4Rc5kSd/Q5K01RwIz4z1SLdTvTsS3
rTSXfJnPJpAljooC0iniDllEfILbzyithSnAO2Q1RvafEgvcPivaCZCsEq/5H98p
fjrPBdHNW3TUIaOl4ZxItqhullLV1ZIKqkdu69UTSzSIqGOhO6v1qqGennC7k6XJ
9a5XxqNhsF7Ia0jlQmWLg+zKVFINHAwOaEtpOVjp5vHJMVQ4MV9ihDiCvfgK+uxI
zoa6oLrlhkgzV6QmvKW9Q9NfoePe5NkThK0i8g9qQvvLtLYm1Xqz36bliRPVfXSN
W1aHDgcSx02RvOw3MAjCbliQqRer1hal2AD952gDrvNditF8/ikImctf9kn8XAEr
iXYVvU+KZ+UGBqmaFwGTn2ynSlPiGXJ0tL2YsP69ziXR5pMls51/LVT1PF3volGT
oGsBywn6digiL3ZsJyY+A6V/GkMdEKob7zHdG/4x0dVy8Wj110hBM971i1MsPb8w
n9c+52K2s8S7oYyhe+AQQK/h8aF4TN0CvGG+7EhBecBcyqbujCkndrqjIoKocrJX
4A9mAF89Z3zjpzvPvzN8Erbigovuini+DkQSZqJ2ryPjLSIK9pELVMKRHwuB6XzC
hxR1R2O/FRt8an2KvPaTs64xn/HpvRjX+nIDQMyMiCMP+2nPjfv4X6HYddSh/Vmh
R4CA4+mcgnqaDe0oN9u3sWdJ2IGsFuYSUlpSNN64wZW3CWUYnz1re1lk9SSpEpGg
mJcJvoSNFCZGUFQTjsy/Qp4Y7V6kz3ZL4wxlmBKIZ45H+cxE7Rez8C5NAo4SRbry
cWeThFEoWmtOErSBnVSZYEMzcRAI0Nb3z02068gx006UPBvwcT4awO/CLa+bFrSZ
9pOdGx/QHGYydUGGrZY4i1ccOMiDc7gIyaDhziAiAI7PdYChZhJOTDa6nefY5sNg
vbKza3QOJKTcIBd2ivNuoIKPQ/KlNPt+34+TgWRsh3W24B8BTmjx6dEoUqOVHr8Q
cK0G4NluTyvorXowgIVSUN3r+gOFaOP5I0uKuX13zwcdEOTpOj/7AOk7+Gsr5rnt
YF9zHh+cSlFqD1A6C8rEQfkX1tifyKug+jCW/lxkwEzRiY5vmVfB/i1Fwgmfzqke
3YN5FHtvxat04qDqX8xTv+OBaynHPRIEJVZ7xDzg8s2QLeiNkziv3DNHhKtXAmW2
/51sIp4guHZHOU7WAcNgefmNE//GGz6e863oq3qxn/gXBcK9Yj/BKsktblH33a/B
AcmL+Cc/EPaRK3YUq1RkmbhN7EuBFlvy963C1B3kXSyWyn6z+4Q6JfwiOtqj+H/+
p4WCt6s22fBFJ/MbJk+d6ZeCQ9NHV0pYwGBvz/29ULbOONqL9wuZ0jolV0OH+ZdG
Rjc7xlRwyPZOTPkSoqNbjUZg+NbxPLMF5fVvTuignP/fE9apGJN9LjN+OjaRhgOq
zj0Tl9ITD0cBdCoUTP3/61TGGdC19a9aFTojZ0ie1eNKn56sgEC5K4tdj0WHau1a
2YxiApJc2jms6zJeD+1lMAqge4nSy+kSwDjwfhOGiwuCUWMbmrc+6gR1lPJChsoZ
K2ALAHKEdlQiQ9Lb4hiCmrHQtPuYdxvprQgcpDorzUXW8+lgHaTKBsgnjAsOrPV5
j/3c1LUZgvAWTCYButxShUyOGPxyTYMUCyWBpxVbLq0PKd/yJmXrck8rjNowWpE6
GfdJq6kzvyqFvUHagRfXhIMMQrgGnxQH/Z+QGaU/BlOto7e4zH+ZigaaZvw+ubJV
Yu2IRxxlxkcVK2Brl8e6Ol/VlIBEGrVUIBHaIydv5V8yHJZK+ezMC/FMKqQANrzY
cOY/PBDIM1HB06wtLLGll6pu+7ZeZi8qR9b0RdslEOhRxcDUlbKqGVxd7p4eyjOJ
VoNOLrlfmqD4MsISsgenDVhv0PQG6EWZostQeOf6rQrqB2rzOVCkw52j4mm6srgq
lgsbkDvjZBRrW4VMfXWs8BRs+9UYqSgOxS+do3H2iid90xl06KMGVkS7o5OPkw8n
5y2S8y7CISlIWKYwYkyEI2Z8D2fnYrC1rxdHQevd501PtUgsuoKt7Yj/5K5mUlzP
mn4N2LhuMMR0POZoOLMt+C/CEx2V/wNuK00RVIPLVLHEjWAK3yAWjhJR8qxkpr4t
freLjJT/avwBm2zBT7heXU8jDAOBc7kiF8H2Xaihlc5cR89e9Ep0iQni6lchbPuO
+4VFXAbVcpfG+/qgcJ+dI9nMIbye1ZIzRrGku1BTYdQE1o7Gj6JGPp2vufssA8Ro
7Zq9QelomdrS8deJlBJum/LM+ZXZVYkCwWD1fs0MMgyd6JIyvLUjqazyJJ005tTV
K4/D+5NSg/ae/QyNl/aVOhuePN798wBQfvsxMkjc0sj2ouHW+eJVgjkHEgbKQx2H
dhFCEnRU8QbgKyrM3COi/Kt+ShEj4fYadgHPChu9WkspsCHylQ9/A0qJAsfOcjcB
oIwQNUIA4lukCWT0zZl5y/1kyQr26B0dBdHbf89WqwDsZgFkqTW/tORFx5BPVPyM
RKV44/tku0mwD1LYVqPyY3JaI9WK57NdQztPBKu0Y6+CU6sekMY4JrfSHEHkv65Q
7LfOUW0WYNLe58w+9AulJUYZVBLV8DKfbni2I9HLZBbW8WRAg++oRpOXhA/zNpPa
78F8y768FMTp2pzUIeINDR2cOFk9kxGrrRi1cvN0QH4bsDmlrzfIr6+DS5k+D1xI
OmxVytdN0bTYwW5ubJNzzb3u8pZKx9me/dYqfd6SUH+7fXbc12pqvKodza+nBSDh
Hy6Wuw3k04neMQ+HMf/Of/3fJjOivQHTnKMGj9XTlTeKnXKhogNqRC0GYE5OAZGm
F4hBqEeJ09HJxWRdW54zgMYrCznr0LdzCkelNf0K1fAIi3j18YhPxQcdFZ0fqfAw
edAA8p13sJaJqid48a7Vw1pJYAnnYmOxhRLnyLvwF0dhhLFcu5XvUgQ+nVXNh57u
v9H0jDoE9/gCCaFJo1CX2SGBLi9uujptBok4NtsLGWsCvTWtNse3jgZVFVmKPdkl
65ccFijuLKDX/EBkg3gqGXnsD8OXuLjgDR8cbkwq1cNUTDR6naldQ0xSuGUTg5Fo
4h7WnfP7xVa3uUriswM3d4eSwLm2IAlR/NU822VqxK7Bq9IzjMSI+4liuN/8Az2n
pdpto1dUiZ1lpCkUrSltmszlDzYk+xlpw2kb+k551JyYnyCPOcY7xvkqaHLFBxv4
SvHB5fhQe9flvOB8ZcDqG9OEi5s8jbi94aUJjIvVWc0P+QJfXs5LJVTz4+bmpynG
XoVZZNSN61aY8YhyoPvDhE+pCh4Lki+DSB5yW9l7gI14sqR4LKG1dcNaQOie5V80
sleEuvNMQ7lsZdBTbKMEMYnNDfS+8I2iVt9R/Vk+O7fWXZZqfSChsvUNM6UiTWj7
dMfUo+5eMRpTXYWk2Ptj00kPPnN4TquKMbHjSuYVp94oBV+mFYb+qdm/fywR44Wu
N42d8zquI7iuTdaI8yUSLI2eXsBw4wubBCg5s0MrEzVyAlhxJAyZrFs6+63G/fd5
Lq8v2HsK7CSPjhRApmIXzWpCxbFrvgIyxyb6a9vhFzikeImIzqSvtEMAEot+SVkN
BTDZ1t63objfzcIGpgDq3zUMV2VISNt8aAXwcCpZFEWeZjoZJPLMZLbVE+iMWJSU
FKQZN2jFYa3M4PCPatJorbx4JKfBPHPgxwamD1FUktObsQ5u5KJH1AMlP8xXQhPM
jxQGP0XIuxaKOK5RdN1snXOqvCBsHE8aVbpJhKIJoZIjmxOQTHIe5ne1xmKQbJVO
CLvBMQJ5dg0Nq1K+9ToIa8artO/Gvr+ezbV4n0HqnzyRftjFeTijj7nPD2ZePQux
t2TWME3EP4xLYhyjuA29wCPcxG2k2JetLgTNwlb0Rjmb8Dr4xMJkKG7t1IIrDVo1
76wvmP14m56oebHERC8mgce16nwA3fB2Mv1XvPCDNQDzcUHdPutmbTWy+8orINWW
2Z8z+AFPk1wRIJ44LE7Ep0d28z+2T1Z2/Rc4AzGWCfa7Z5brmdoSxioiCW6Dd+bM
CHrOkODD0Iyyhkcf2DUtEhq2FZGxpcOk7Vv5UTWmTWnimz+XWcH4vUTb0XiGihlI
dwirajoehEKGL+b1epfJ9rHh4RJZBhQYr1nWZRdfHZJZGexmtPY12T6wFKDhYIdD
pjsS4iIILH6ux4Zu3hgHQfBcsBhuwhYkp9JKrrO5mv64SVL5QuDb8f8p8eLLAbFN
DFsixPH3geCh+SdSxxQgp3WO8P7UXpnSE0gnlQxWG0+4CYWs+iKYfvFQ0fpMMCXK
Pqmf4apFMQg32WX6YOMy6SY1PCV16yEmM0u/IPU02fuTBr6sdWXZCVIKlkoad2r8
3c0LsUyHe2x1gD/twO4nG4uo9RNt229vy8pJzc9ALPy2/SG2I/LtvYPGo2NnP0fo
JjSguLy40QmVG19MPTtxUiC4KrftJE5R5ZjLhFUR8gIa+fMKjBy10gUWuFaCDQcT
0DLpby/Qy/joC3xGUWvvKS/aC+5pejBe7y5+jyeHXElnfv+6KXYtlk7iSsu2vESs
zSCQsS+owMbcuKYqY0e4LOcfqU4RsfNpzKFs7j8bxt4W7Q/wQA1ges5vMClE5uf0
AEKInJ6yxZSCFK+Y8GGgqS8TeaSMqcC1sVgpgncX1AFKblLx1pRAKf2OyY9Mf1ou
fzuthRSu/gnyrydCO7A+BVyBM9glIKq9pnw1dY75B47Rsursfvzpc6+yRvh5CNek
LdqZMMnbGyziGZaibMkXBVxVK0LY3zHDUt8mFmjAyKGfGPWDPtLkUpj29fpYbyq7
AQdudUAZI+Oj6bCWP+2Qaq7bG96wM+EkpEM4rhWBs8gNbBZP0vqkYF2DC16XRwKU
bBzIHbggdcclPR7+6PdH3TH1Cvkn0qyYIrb1M37e3WZcOMxwNyyD/ff7osLDJbCz
y5yo7DY3qcRjLGmKqbWg9aG/DH+gohydjzl36hu3CKK1/xsiDZ2O1Ywn/8C4bJfx
wc32h8RwrIAdFkpkVA2baTZFm/UBXJdsxZTL8hx6IJVnR71o0bEmmgeHTrhVbqW0
+WbYXTHRph8Ye7uUJkUPVobhLWpRr014kuzq6BqaTs2XojQuFxjhqM0OxIRmg4sy
uMwg2vDK2K3+0IhcVU8iHLX8PHwTb6OC1c5PZJ79pUlQ5PyYF9aQome6N9y7FC7f
E5qx5FYjrn2bW0QKfeQj1uWBWgkXCtg8nLT4vEPZpEBpddB5s2HAhaRz9zuah7xm
+hf+gGavvhqAAk/4xCmOR82xyZ+WA5ota3YKFV0fksHpicNJA70LEvfRFyOF1vpE
DlRetYckI9krypJc4hSEgdc6xX+Ew076l/WMp1nLzgsOCxh2SV8QCIcE4tnqzZZZ
nDQyG4kgznEQhX66AqV5N6IkRhp1EfTt1b/KY2/3c2LznLfI1ZE5dZBjIsB7a1P/
RLsEr5WDDzvbveEOTzdbzY3lDD8m5cXgdMAYd+oFIMdzlcUh85O2kqBq5UFQyJop
Q5kQz/O0R1GrkX9NZX56bG0vMYDOBkibPoEjOKDlkfnZfFucqaicd+3Ro5DZ18Y5
WdOxDvDtGBBlb50OcZrwP7BiffPenM75TSgA0QlXkGR/NK2nUqJQGfINoouall/A
fnxk78Us/y6T2aC2cVUhlNU9+E7sbNJf/eb8XHV8kTJxRgS4zoOMJdGHAogssrUG
u/77UBHbl50EmseACNRn1SjTcH/lWF0yaDC8Oud2Vz10hvnxz1FlR4WzcBT26hZx
w5u4nGC4qcRDMIyAK9qtr35nYJyQVOjn8PwqXETjpk6wqLdnNoOGDBbGkZz/GZLP
2+dONSxe4plPJuYeCWrBH93IPnSb/UCYX6TJLeCYLKlHDVGva1gW8UfGTmgSLxne
v9/MVQTsv0PW185nqPozV4NlixUCw8f6KyUzfYFZtjsz1rgW/tCuISIDfLMreJQN
Rv3R/ud1Avy89JXd4L/wiiG27nyNN9MiBmSOdH0gbwYZqgu4L5lqqrdqr/DpoT0G
Uk7CyCrfdQtuUI7pu0PUC9UaQciiT11jTv5TWkei9eB7XN0wTN0mscm3JGmJMZJ5
3clY9El8FtedkDmLdZkSk0zZZxw6h7gKpE61/64zee5HMaCfICJN8CnJvx6p6qc5
uet4FoeSdhe/mkcAmQM6Qw5fijOXjNIBmIe1QMjC1r9ab+rsLASnZqzn9JY2lFmt
30DHoPoaCVv4GKQbaZFkbW2jeaK9ETdd/jLQZvUYjsZYYpFwNo+0pt2oCdAqG0fH
q+qtPmscoNSOyUaGqoiVXfTJrfK3C8NNu6xjVpSTw9TO3vo+M4Q/+9jIyxjdSnwH
4CZRR9mh1cC1jua0+DJYGPwxMZrZRJZ/ebyFT5JnzNDoe+rSqb4d2mnyskKtGBGT
pFWQMveEog2LHEdFEonq6rQJqsbwyD5V5QUddfZ0gv/wH3+Kbv75wTgAu6u5iC0+
QgQMkIi5oAkKZefGadwKFtNm5hxNL7eN1CEycZiYU1by7dV43gVk47jZqyR8FvyG
hs6MI2YTF8Jt7VAVwXn2vX2pKWcmfR5nZuBa/TPylcCc4+fFrjTvoW8XOTpRzjzi
giL9plkWx8k5IhdPOL+Axi2ADypAk5+sWg+Y41Y1mNe5LHgZ0qDcI1EwIJe22hvH
Gtmnn4dt2R0JCnwY6Tdy85LCTRy6RhLJ91Qf2+JxE8bvtkS4Hcw2kifZkefzQgUP
l+0jaPUkEbqsHqUVi2c2i/ph3Uz6OHTdBWMTkasewCrTpChJqfOqYAbw0fZubk1W
4r5ufcN7+fPgIBFl6tMU0S2sl5UsXg24ULJHFMjtRF9roxLx5aTS87axD0OPIXf/
3ChzE9vyUiKkw/wgGeuFVC/0RsiQFG90bgyTK25YqKvbuIC5bVxRl9MPHBsqnrRL
6gIyjEYwu0P3G/wGvGskL26uuNAj4+VcQBMeRSxBu8XbSoBOFRPD5c98yCTu1CD4
HZV3Fb77iVb/oHtqmVFBX6O/Lc8ReLvl+5hWmfmDSCAhlsUsXK46hWTBgCFysPOa
bhwRGqLxRDk5Fj4GlKmsWX8V9LMglK3icwDpcE6stpijQCC3RkjxP9AiugpNoy6/
FCNsIjdRAZwEWrLOPN/4qywxAaeSCbtWIf3FBarq52Agau5qXngO9dySi2ZV0bN8
1LwbmDgWaOlloBsVMUG7v/jRs88nU8zIUrC1JYxDKDti1G97J6Rigg1/0kkkSbId
2YNeVEwxruWFRVSNCxG4Bj27iQLX1NOau4M9BJ01wgcx/dT0vNvqmcKV7/xbvSdi
z1k6gI49k7CuEFChpifx+QIVo3reEfM7FnomhgbOvKW+vVPWwLDwrXZl+qhAOJPs
0SKrh7Dhs5IeYxIluizWh14H0A0Z4uxnioo9rMoR5vqqZXqvpOmdchAYa02EvaN4
xAviuUmL14TUF/11BECY6r1bnHmX9SBuDe6AOuo2jEs6Zeh0FOOiNM9AqbwitOR6
6zenoFmL8fMVkOUb3eTh+JsJz0pZ0LKxyp3fy49KcBXIuZrWX4eCrxcVkaGnb6dq
P7a7PBLP08/ZJ+rs3ylX3v6LkS+CVkmiODqjBU82sC+95IpVf7AtnhlWcnOahzS/
6WME7WxV5gkTwiNPPDO1zoHYejWCOch7CXhodIAvubp1/n+UmJJEXW8++9A7JOEu
LOcsKrbr+0lm1uMm1NXm++Kcp6QBjupGwM6kdyVOkxzMbKSx0RKJCfa0y468jBO3
Uuvs59zVUwMJHabDtxlTDGhdc6llOV1kgK0+XUmnBSPqgbB1l0LrOUXD5RRSAPKU
NihfjOFkIWoXLuq/yxQ9aSyMz374YQsmo7uscpm71kgr+8p/ape1FyUUArSFYqDG
t3kFf63LdBXr3NA4IzxIzyBXiRQroYPirhPYIPtfTQNIxzeTxjtrQvjXi6IPiYX/
WuxD14vjXoOrZMP9OIjXpLP2xNQj21xKgUWvxFm+khfDFfHDMiSPxo/tI2bIyzfK
bcilRtXBhCeesHsZCuPT1JyPg7Sz9AbnSb2nNfAklCXvITTyyx5OfT/Vp6cZ8g4M
qdZyVSYATceQD+sht8t8ErMF+5ZDBdT7gDVGu4JUpZK9jqWIOV6OS54yXvsal2Hx
FQLCLs2YLyKPHhMO04S8fYxNWH4+DoEPegh2QZxylgQLF0wazJZ9NkgCjwWEtr5g
cudaea3X/7z2NGpoSM1cR5EA+OHwTG9F14QGNLhAnbiZc7qZq3h5+9vFFmA53AbD
F4w3dG5lb0sSZuO88fcRC8lErLOMoe/n4XZCkq0EkFearwimXNcIXOGYG0XDA8KN
Q1yguvKG36fjNzARglINrgQitZAz946craNHAIlQ+ZoGQafSXlLwQ4Zk1wgldOBZ
GjaZaYCXSbpnjKJNbBEZTjvyK8CBipMqyLpkGcfDI8hAo3+sbGadlqSiX2wjphtD
vtAm8UVhPYZQ80x1XNm7TvVJtAv4WkWmwpJihrgfkza2GyVx5bVmB+zHTQOiBHW9
FXozIK85MIOtP41e8RwHaM9EtFXDY63R7xFVITw1GzYBsE8qggrNmhWEp5hda/S2
C6iS+UwblVk7OtzMBIWrW2C0y58scKClXKYhyt+XsU/nSPflYFIidNk+oXTNoom9
8RFfbwl04QFuXNyPByO5E2yj9MCdP0LNJJ1EQCZSkhGPOsD7brqqSmXS0okQQwvE
k0cNA0qQE0N7UwZdzlFsNVvqsJ9yXVpQhqjsbUVtUvhUfT//WbaRinBunmthb5bI
Y92UelaBYZ4CVSBPzReHeEDvnNcV+R6FLaQAN1Ko2N1m0vn3tR8LVvf9Naih+mLA
yyXSJU5eYYZbMPlInfQGwpVfDuBKUHhlicONTAjtAzkPxfqD4WyXRoFQs0O0USpi
83C3xx3yO2NgdaR2IGbv0+M5SnOabc0JiZLr2BqAoQ5ojQ4r2s/AR3J7lwXqUsPP
kdWjqLeo6x16Is4Y1KRmQOr2Csx5uGg+fBE4iu7FcpLkDGpic/USauKHBKAhEbuW
yCsFTjvWhPzERu5GsJI/1JCUULNkXWe1GUhqgJNSbITJhTKz1Mrg0m6Gj2NetbM+
r6is08kRiAPT+Ry8cH+Zb5veTxtklI+eysgssX/Bj2yGkPO9oGYZdGrspSt4LlSY
KlewqdaZkdZS6wuhsXhS9Y5HvKnHZfnLR0kheoeYJVshFIUkQTIXtC0HtdmkIz+H
lPLNUXzIaCZbSsNPDP5BrP+7Dm5kBAFP3+D6nb0Uin693JuztvXAu1HUIgLUFnB8
TSR6yvyFUFJVGqVGr6M7pwUHIQaUQIrX8aFFb1ItLY0aSm6OExOt66214BJwjnhC
CXQ2z0PdLukVadc0+OhbX2GGFPDSi9zjAVNponUcrOsuH7kxQaY5ymkptSfMjnmw
K6rPyOxx00uHOAumw790ZZYNO3ntZTH0XSQHMV6xHi451cyyWKo4JN998s+ZJCOb
LJ9z/B3oiGckktgM5Qke8eZT17e6HrTyLkCX6upjgmTHlqupuSDc/gPooT3F1KPp
RmWScSpiY0ansvt7tMijc2/ZHJyjLXnUMqILoMdqgkbyU/ql0h65HrSs1n3tT82T
wpUixyU85CwgUrS2llnE12KnOzguAEgv6+KyIxN4BjLnUZN32etFCfPgtN22TVJp
6uIvVE1llkvwDDHHxgcYC2YraNbhzJE5eCkqOGWAleC1DNx0pXuc4L3SOZmhAPxr
/pA8TlYfmIOgkKKKUDw9l6QR3OLdcfDLXAzgEioQcCywCsJJ4utRd+UVw9UiqNBv
37LCP7IrmuwfmU27pZmeyyXjmwUJH6sDSp27zNID65FDaHNyqI895YheA0Rsz5Xv
iTUprIhcvGAZP5nYXtSz6XvZmp8UiUBviz/EB6OTpzpVkvB87apdab6L9CeJGPsL
ZxfRdhUH8TpjI/OUEUCXhlj6PhcUaydAieb0+qXVRFCTPQ1IN0FCpaYTq8mFgmUh
3LhqX/CS4tR5+qcpcKnSy9y+4WNhXmBd/90+IxGmFxZOp7tYyuJaHtYFkj5x9CqY
nCO1+KlcfMCQGjWwV6N2ddAV79hOW+ADm+vEQVBPXquVxgHpJF+5Wvz1EHUDP+rS
GZRHZKX/3FAUNYkAgGWiHCGvpZ+eqx4RzijVJNb5LPaidQmCsJveK4Zb3IYd3q0A
SNG+Ms/hFxterQijUElSQnO9ccM9ZixZcwI8QXnUtHfspJdD+R7Yugx2uTOd1hBA
tCtIMAejAakWCr7WbtUNNGydoPNYOkAOK2f1vKMLatJveU1ch+thjpJJZ6GmP76k
k2D4XtZcJKDPqXEYTfa7TWv8pSLf0lWxYHoQuWO2SFr3u7b7xMd4SF7gRBOU94/D
5uhZiKHli1lxHQEKYW8IbN+NwI9jA0PfzJdW7KKukhhvLiLAfr9oFfFvusm7hegc
G1+aKQY5y7uwNRnptU/F+9eFZ5MM/itNkajKd9kvFQ344Pl1cCCZ667FDuDcUasS
Z2RJncKe7k1KvrfS9XGd6JCMHZj3797k487FOcwEZ7iIEAbdlP8ibcPWxLaBJvLh
rnSuWCOc+rkKLNmXomO2tNtX5plLy6WztQgbgLaJkYwZs7RnJnRb6L+vrFJcX2rP
ND0l0kEUXyzoSaU8dKqPD4maCm+yJHNhPsGxuq25DFPIR+YEJq6KSfxk8wPWwr/B
`protect END_PROTECTED