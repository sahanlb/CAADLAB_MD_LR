-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
jBKbdtQhicEXjJVqM/8+w+mHcK5hTQSAQL8Pbj/QPyZNodlcQmrKwPbPIJy1ASZT
u1Qvdog10XqEUFY4f+w4ogxh0wW9apxj5fpBspXIhSljZyefmGkSuMPJJzh2y3cp
ul6NSbU+700GzDngSd2Ji+sMJ6dqf3A3KmXMB3mniqs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5629)

`protect DATA_BLOCK
JcihUmqin4UKgZ/ehs8CKTLGMNcsf6gt9oSrNAOcRHB+osSgjEx65bJyhFWmDZyh
J4m3OC3H72+Ko5XYjPpDytPsEdPxo9CluC3HPXVvQdPDXstj+/XHkIgJb/6KKbOx
uufGSx9oe2R3UPv6hu1CBVYKqtC5dj3zExY0/S5+bAOV0iUtGe+VVpgEFt+JMS74
JyPxphfK8Ou8tzsTjqefdHdR0ZXmHEOinDGIVBtPA3aDKmdfhivN7onBZ3jG8Lde
x8W5oYMZdqE9U1464vqknwz4IosxsF8p7Zb6sOXYNHwaR3uWTalnMOyL8E5rDuKL
RURpM0yd2RhkQi8Bl3Di57gSc/U/cPh3+QOZCZSK2DXip5PO0tOnqhIp75VNk0TP
nJtv7kt/wUaQG9vCNBfIAvKYrgFjYTVh6AgB7aNoYz0deC+edj1++ZMAdnYUJe5Z
kuE/BRNqUjEZHkp33QmWRmgKIMG7Eaf6LNYtBgLO2MyNRv9jPmDEAhIgmAmo8j5+
8EXlNUE/24ibpjJ3GLtLBW08KaJp74u2SZYrux37C6l+C2H/dP5Wg4FtmveDyl7J
zubW/fha0dCiPTqMNoBaCGziiSz9ffZiqTUPfOU6v8GbkXSXQ7rrfx+/qx51WLDq
jwjgn3ykTb2WM6C8caHvquarUtxXNHpl6xiF4XUXmqR/FKNFsTqaqnChldIZPkr5
jK7xfnb7uq2GSE/SnW4d/A/1617Ge82vpiWEaO6KHqJRFZU8HaRsLxzsSm+TyDgM
S8DT4JegqV1WieOB8+HFs+C2NrfAH3mDlV//2hUJLZWgv8dUNEU0Cm0Fg0+V1Zva
lpAtgizZL0bZgJop+lFlvKy8lTGrjEgv8/49m5TE/YSg44mVHHAoS66ho+zTt6Sg
2TmOuvUvlr2EAJI0VRpemD5ETdNtIBEmWxgmwCXcd9LNOirX0z4txYcYfvPspKhR
qyZBcGzzHzRAjqNYTgAvSCMZUeM+T/m65ytjuUXo87O9fbTX0LCq7RplF8Silgtf
w7cBnAny41DFfoNes08f/IyDL2y2/Mz0AU5sdGNufyqYUAgOTamTeLTMKWlAJY+H
LtSYIZsFK7/uCfYZ+WVQoPZpcW4Pqt10DulilJyAMu5hysiw8I92C9MusfFq+iKs
+mxJ9FKmbKo5b1gP96QDmpaY2Q+6WMz2ye8vsYY/Dij+kTB2PmvXrUhYa/0So41J
azZR+H8wEKopm/8qYmCuzLol2JeCFyxGllJHapyffuRhdQEbeb66q5g6LUrhQCPH
ntDZJGgiHM6Gmf8GIxxj8X0oEg0yRmLpQFs0OjNenJ+I32x9zcb2++5hk7v/Y+2m
tGLEi70xH/BmXo1m8gQiEy6w4GnaVo7OgPFE+4LEs4kOeiay1bjUz6ltsF3Hran0
jK8dxQ3IWCQwqQoBx/ZdQ8jF3V6Zi/BVug4r7I78inWFA91fsBaJa+2kfPXu4WDQ
+pt9b+cJ7TxluBTwmFlOSgjcpvCt66cszPzFA0amPxKrQSgaEku7HB6C5ap4kzlQ
tQoNfwF8HnHZyjWdZt8Ws2xFLnObB434dgaAQqV5b8VqZnKEq4keqd6FaaKey23O
acpr9kfpiQtHGtudEsAw2Dx/GCdtmBcuMj6eqmbqWetJfT+tTRQjTWxCIMlLHQ54
vU4o4P9MU0hLPJOb+jpWT/fLIugBnmtME2DvicbRisGgf2Iwz7sVLOsmhfPOep65
5N9Px0MTMRelM98IkbafAvhu0PUJKs0KaWAV1xtnpK+SE3SbqpH6cohzv7/g0yvc
HMxU/xFx3rTpTTllppgRx9Nu4i1d54cceSnOXI7HnCiRbObZJgBp2SFi0kWRy5b+
0DwbA3OFWtw2+P8Z1qL/qvbMdCRTQHkZaYeLELjCKE2epzBLVspaESL6/mTPB5tn
NJvVGRoc2Nuf9Xabsx7P4QMiQ5fPa0p4P/jqiRRCTgG6VxcVgw+QW3l4i6uNbA2L
Y0IN4vYexYR50E66jjQu+TzwbibSLcZJDA7WB8vhjwoqKe6GWCLrXiUnxUuCIvoO
xBUtl/fIB+u5LYkmlVDvs+q7RzfEF181UuWAPyAdkCzd3r1bz1k8GEmi4h/BJr8P
+9CXAZh3svby2xzkgnDOr9TLx5be1707WvHhdjU0BYQzBLxDQzyR7kpXq2es6oAt
dRGnQuICItMxTFrfsxEhr/SXhPnFiMgM/t0CZZf8zCuSzh8t22sn540hhnfmGfgF
i4oK2vxQwlQN87moSfodnfl02LXpI8z8EUT7rWdQk3BMUEjnjxFF/fiwrlnbgRA7
pmbird89DNzMfWLYBpQa9rS1Hwwsm6I1Jm+X4Xwk+4sTX01u7lN6qQ21m5wg4Yel
2Fh2OkbGW+bEgkJHLzyr9hM4V86WFIWg/FGYPyH3my3IxDSvwCwPFOueDYx3r00A
X4I1cyIvXnIAku/3P0bmISjM0vgiLmUVv5d8ManmVNTFIQwVZuoKudIjJat9bgsK
CAfDYFwpvS7TQGliQjaLVil7xa8GKXqjZrZNmtEv8NBw+DkwWFbXyfBDDa4V5lRr
SRoj7s4YldEmZD2vCYZJpcJEW9OkZ3zRB7eNLq7YXed/N8LX9HjK3yw9L9/nPUTG
ionbY9ziEV47Z1a5NUcg2/wLm1QjZwFJ+iGhIrIJX4+fi4fF9J1ElW2yRFd7AukU
J/uyPxfe7ouWFEA3+tMIbh3onJWg5bO+s24tUifyhn+iGmbfeWCpyfdOQi12bH0e
rlj5YftReVsg860Mx4M2VYGsLw1fdGXWovM9fb9YgTCUJVg0nMQThniu8bGfgqPT
nlBlsHc+7sMLt9K6KRDDZEAANlCpbmnFhZNvKhVwDH8s+ybg+1vraigORGjBdhQQ
Ng5zdRqoTehn9R9kQktSTujc8UQa9kY+NUUQZwuTspk3fFmBpuSY3mNXSZ6Yla5O
MFeKoEIEsvUzLGxPYn+qZ4GpjtWD6TZHDmadLnr0v06a1u+9MRf5OxBde0IdiUpN
JNo7sSci8ZkCXDaB6sd2NkWGBQ8EEa6n971kt6GQmGLWPt59nS3ZiYIRcHkbbrQ5
vNu8djbwswUOFlvWdr96lF/tisEmJERYTKnCWYyKzhKTyAj/fuASAEDJJ0z6B5Vj
JAAP206FiEjSUSxjPUdvV/7lhGK8nNOd3lC0AcI+eYkOPGh7Viu7P1IT0L+k9Sku
85GZsBA2LsdiLuG0kSMru3xnf0zKs5lK3tnwDnlSjsd7Om1wwtRcIPcRELosQ36N
hM2gOtKOVgSA+WTeZLDbS9HrFecyQUKqW/Pojl5ZtpWrkEKJ2dfQLwsCWxrwMJKI
OJ5LrOFGJhMcY9YU02oVFsS1iEdtRCNL29byw98RVisHMfnJR1w9xmlKsuV4u6In
ygLjmNe7ZeWQ+CINeKmK6FqCnDHsX9FkzhqRltl6BSfyxVoWT9/ep8OMxO7/spzO
j+zdQpAGMZGb2kXa0JAoaqvrW9j9dAOtFRx+ZK5uRqEpEstPCneLdCxjCWbw6sen
sX8CNVCwbFahc4k8FoZsXMbIEY2rBKBci9Vpv8Mey55Uj06xHP3zNFZveW/B3W7Q
xiCU3A2y5rqBRtqlx3h8oFghD4KOXf9GDL5QeDy6xuUu2Zu9Rdki/KSLE/3YCDzo
Xg9oQbIAY2QVTUS/R9yYH3mlcSjsLZB4uWrs9fW6qIC5NOMBqaQoQiGLSepKI1Pg
vozMJCF2pFwwTihlKHIZDGws8Aj5q0JyPe1J0eRdnwXWu86fedAOLe8lEGvi1BcD
UG1z03shxmH7qW3vwDkVYIr6P/z7E8vpw0Z03Vx0t7hdqtqVbUwEXv0CWTlvqyRf
wnvOUJcFWeKrVn1OAb8ub5xw88xO64APPyz1q1BsKWsfrwQzD72mLKaLQDRJbgv/
dTHG8YF+879YDbv5ygzVlCrp4zyI5rfL1Ap5DsZOtEaT37xpWAcOX2IFS58k6/3T
XuFW18j1DVWVqbijOYzX0Db/KYzhtfN+hxOgyVQX4xLSRgpVHeoGL0bxbhatdBrp
i/1Dj372LgsN1Tjrg7d0BLt2S4C/lPumx0JriwYY9cmzfw7feWhrNZIY7AhfO4Y7
ucxpoy0mQGkHtu2HLCl4yye9NLxYo4Axq/jkkYRojo+CHJTx8s2EwEveG1hNs3ac
CMZ4tfnC0E/RBh+fJ0r62eVu5oknaKhjI/8rMk6yHctKFaoMXm3pziS/QuB1WheS
H1piBL/WWNTVgn4QlHozuDYK5uhloBUGBkClxMpTtTxQbxXJwVx/sjMNOijuKA5I
gSQlTKIZ/PoWd9UsocMd4qAA1L+7exYcPfOqBb9L1Q82OdkzXKrv53G+PCMHDd+S
dInz0o5uKP0cWgA3kG0mUpZUPqM1M/IbVnj5tl02j6hztDmM1bdL7iUTQgtj9D+Y
V/fGezyCHmRUtE171ZP3OCYECOLKGbd3B+Eg4NC0NsYt5V+oaIBklt1ytochjrIf
7rXXS5ZaAv643Gky7+5D0R4fFPk3dDc2KyYvas7uTL26/s1thkrE3eXF6asU1JoU
EGU0Q029poQ6XQEHERKaGaerytqgWK1T7LwAeDlTqFGkDbxt2rAY0H2dIukIjCvl
1p0Xr6Bf63PTjc8A1lYJgEcPcHasc020NJbaXqNgrnvXXO/MiqIK4ktJjsiFTBI4
FSinF45wFuzPd+tmL0zBlEnxJSnarPAG24bvuy5UxWgQnd/JjZw3LuiQnmQm8JNL
pI4NrQLY2HdFppYVubmn43zTV5NrJ37yhNIKGE6mvA7XiaH41eiB6x7MTiAq1I5x
zMg/DCut3cAlI1InrBRBbF9s+jELJ0MBX7EZNbw2HvcsBn6kNAsIMxyxZqg3ail1
h6RoaGSj5YTJtVUzIIBVPmJWt/oAalmJqCL9hhrILfOheUUtiDw/DpX/wYH+qZEk
SLMxAqOqKe8A0ExuEv9TSwTsCAFA+P2Y/Hdlj8qP+AjK9rgPayJW/DYKVslj2aoB
AOr0NPo/R7GwzR4mx6v8Q9suiCrmSO+4MMmR9jSHKr/4a2EI1ek2323cjspAqdIB
YlpCoP9oVIKB5yS7pFZuj3HklB+ACPQKXmWaKtgyIKafd36dEDKLutHtxWFQ+x/l
n9teZHGO/ZGmHpOSjOhLYu1cyRsR2pwHTK9Kf3yFL0uc8zG3vbON/vw+ys23WmRF
EWmKo9M4bvqNuj5+JFBb8D46noYfbL8Qlqp0YQI31+mvtF79fdHgfjEwzMhf7U4v
fR0evJXNSqiJenucra3fPVwPvGo+7XMZrbo9trXE2SCsGzszh0kGdmNASxre60vJ
T3ZafwWjaFHtwXUjKdGWyb2HLix9eocnaAItwO4jItUo5B5irY6LlRtTy3eoBApR
Bjix34S8Hk3x85EUUHdufH2jDSrCClRn6qDZNRbG/+AI+QWQ4gKc0X9Rek6LLaS3
LSlqhAAc+fXS6sGmJBhUHRVUVwb4jQO3gXqrJAwdmeoZLaNBahHAdFB5+LjmfX/n
C5tVIyyanZXq3QVAXq+klvVsCi7c3n+kYSgBYMAJeesfUgKy85lW3opGCwYcpxQQ
fxbdoNibJ3YK5sz9lCEPP9ZCURlD5a/jYVaxGrphT4a7pzchrfj9dvgSmC0hKxCE
V08+rcmziFB6n6lJdp2dL06OVrHeosPDGTMANCSFMlo8Uj+OeJda7nK1pqI96pW7
SCA0UAFOA/juEQR5m8MzgpXuWcMmFFO3FtHxUy39qu7FRwEDuBiWRJAeyfLXcwpM
9XDVgFCUl8tC32JRXNoArsPshUZggZOUXypY5wcLgP8YfE26jHgwJli7R/mSTqed
weZE3fX981ts6gPtNmETd16zWKHAYXyNRcJJ8PMKhBcEspeQiz4rZ/ffQfJWuSDX
lqAGKGI0pH9c2+DN9B2WIW6u1Ia13FVXKITMNmY5dnkK+jNUgVo1qY5vueLt9YVD
C47N2f2EhZeiTCxZvxkV8CRVopNTlmcMvANVnlvUpO4PaA3vOxN4hrZkHJFKCzcx
ePOesJMtaUgD3dTPYLP2Tl0wOAiRC+U5/5cEWHhzczbmMGfnHOfXs0YDyVEQzjEE
vG/iNici7ppojlYtnwzkew00fFpEQdBXisZBQ2ALISmRU+GRcovpyKl3QOEIrZ0F
QpAk+hrd0cSYqK/pdpoZ2/20VYTGoj6k8srlAyQNKGa+dlueWZqbk/gDg7RgzD9Q
chjYGIqZYvNvm9e93QjL9YtW3rG/Xjo/LOLRDuTWnPCdHNhzw7s+hmGvqxqGzl+4
Z1fbstowO+LmwFuNilCTzBaxusRQ9B9RZxPTzPXKdi03keiyVH3BaIVNUFwVZJsW
Ido07a8M2ZBKZY3qNdf8TEd2cxx6LCiwlDPdLRF/AcMEiT91Tgr3pB/XJgkTtd1P
u+BvMtz5vqTNVu9hU8DAAaGWFsuQ2/+AR/w6txeJOjxBzJVSmEjsLxAuHTYNUYSE
eOsH6C05lWbAkXbS2KZy0E2cXGsblq6dBzugLf+rs3UHPFKFH6g0XzTHCw0MeUvF
NtSWax/+LYVGMCmHftvhs5beZMbRUkEiCnYDTYg1HDO8qDA5DQ3oZVt35rjUVgTz
cb4um0tUvThHgoGWMz9Jy9+BLyjYleqWdJtHYS6R+p88bfUTepizF1kMEH+IN2C3
Th76/2yn3BXZy8Kzv68tDGIGF3B1S6VirQzC+3mxEL6354jx2t3Fl71dW+8dzJaU
delEZzSHESRsmNVTndhvbHuDxrk5WMSzu9AFDu1CssiCfyn6pFXIewBsd2AG/4MY
SacV9w3JXkkFNCm54OWZG2mkiKCEGvbpRYOP3TQtxggcJX60GqtgyKKEM2xUkcds
mY+PAZNls9EmqzxMORRdbJHDQbTqhJmxaJZkDKMJASgVNXDOPJvgBDLgJYwstLEO
Uoebu7ZCxuYYtpllVv4EjbRjy+Le/qH7OkF7rBMW+Tn2KT7W8p3byqoSDG6oJN6D
9eYl+yPSV6FZJgOJeMu7hHhS2rmx1dZhxWavfAM9PmJxEl7sOxtSoi3txCod0ab/
/RXT3OzPTrHDyC7Y0iUlx1vJdrAOdiLyLzYcRLMPJjIgeCyxMIhOnajqThyABDrh
JnIeQwOvn0Cc9i6XwseA4Fi1r3NGyyo36AWQGkMveLrDyET06kj78JTMdUsm7m1q
esTtVdy1haEnEljtAnIsyLKAgTUi9VkKfemUSGrsD7wcgwPp80vsi/C2G31eVBox
VBq7JuA3wITbXyj2kgngjGUuhUt50417ZUtgMFDIHsiQYhYxpwa25Uaz2yPqdUC0
EZ78uVHrAxayIv8dZKMFCQ41p+tAyBduDQdNZQy6SlNFdvrCwtcRDdBSpAvLUV8m
Sj3rb5utSH7WHg2QXOcQDcIgTYBY7ViDDecJhl9TCJmnq75P23jwlrXQzX7IHzcy
B6GhLaV8ZpV4dEfKkRnG8eG9i3q7PTsGUZgggm4m33InoDg0t57GitrEgRCvHQgI
qGrHhvBFqIhZ4vZ7IJGGT84AmiEU5OC/fTlXZDm5v9Q=
`protect END_PROTECTED