-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
fa3a4lAFZ8eVZ846T6m8q9uhhBBD/s6hSEeo8ehYJ74RM0UGpEzwpYBSd2Mv11ME
Bnhiom1E43Tdnaqbqel7aeWqmXUnvGxW7ikTtZnayKHNcYVRKiYeJHoZFXDfVklo
RUCulOIwk0yxr/opbNqSjH5ByqWpPAsciA7WgzrHd1AgrWM04uKQZw==
--pragma protect end_key_block
--pragma protect digest_block
PDLSCMGt7h/oSAxlVqplewpIppI=
--pragma protect end_digest_block
--pragma protect data_block
m8H4aLVgu3wkUsoaK57jfMqY3eMfgOgdk8QUzu8x/leU8j8Wu3Z3I5Fhfq1Avw3Y
OjGrKlgrN5EN07nvLMflTrKoprw/wQvHEsHa8nX+yX+BUa+lKCfDL2RHDmG+DxPn
rRF+AVHpqCtRCKyLFREc3yn3kYqgAOxzucrvYWCiehwZFYVUT8k7Z2haDU5ZeZxF
e9TKbjrloNoqvCI7phrtVZyNaxLDjoXnAUN5kft3hd77S/wferJ0eQ5Im1WeeUZo
skIW94nVMHtVHEIdHmwjCJjGGuYMkx8zI7DBrneWiG4HhnOcrhd/GYl3Lb0WWXto
JAEaYY69v1SLW71s083+Wpej7URaMAOr+fbuQEYN9xwD0gvWOnqcDTmxSG9dU0+K
4YzK2poXqZQoypxq8otXiXR11Cxi80OzaA6STRXP79Jt1dWrKWCOLtNZOLeiQFeq
oestD3er+eIFWGehoFbiiksdF5yN9f0a2vT8w0FJkxO1SK17ZPLgE+TM2ymZN3uK
sGkq7NnlKpKJUIwUNrBxoZyZT1JVfcAc8Ke/+Ath/dY7wnPamdZxw7fJC3ZnkhoK
Gk90BHRm5j5uCut9wZ8AztVsVZR+dz4mkbjj1+gWNIMGtmQojLjyDONYiuJzBXX0
ftPPjoiEHxk+yoe7NtJa7Ijf9UciQWz4ChZMTSCbg8EVwyZ3LOPLlCzTRZoUH2Tu
ZsM46XedbLPM+KDon7wqAcMmz4jaGwPRov/iZ//emFly0xU9uMpDOAgPfbq2H3tn
JNniceY8pKmAmOHvQ6lJHb32QVH2isivAwx6HY/5qc2XtO7fVdTi3lFzRgz7F8sb
Qzc+wpTqSEIP0QwPh97u3rFLYpTlk+7xnSkigDmyvIkGuA1uOsa+6IsVJC/Kuv5w
5gWhGmGhkMXwqejYi1xz4vZf+ht9nNrD5ECOmHkBY/RYPn7fi+m1UjTJfjuuBits
P3AA0r+U+MpnMsE51bUuw5Tylg74J272VDMX1+HFfvgkOt0avZOK8y8TekqHEYQT
IUIfJumJCGoGQH7V/rjBj9fbsWyP5lGehpQ9ISrfJD1PvY53jRx+N2ybl2pOL4wq
8uJtE2E2Gn95+q5gJPgdQN/14L0tAOUgutQK0F1r87PHkRkl4YaUOoef+QGMeScC
XqAEId6A87OyEArBfS5XZkCzwjSQ9enT1fJyOVd8aVuAaAkgjb4vRYMueXc4hzBX
ovRBspnDUhmroOlAxQY12Fy8EI6RQwQm2ud4S7RQkMJ3r3y7G9qh1hLZ7A5/CiYw
ErOzxZTPyjItjzQPxKMiBDggO7xG8NZHuejJi0bcc6Y06zGJAmAPFbx1lyE0tif6
XPPFXAAiZYoWYfvWGZwapv2WHtKI6kTZsHkp2nmAi6mD4/8FKgehRwQzAyK/41cZ
rYTnzb4PIz10C6B8sxKS40bmF8XxLJgxLscbgwa+3hnln8Io4iDjWsZafl27tdTA
Cw3QyiqptlgjVjhtXc9pu01Dk73F32b2g6iZOvgouuTQE+hkyQiNk7hMrq6fGlDC
VpE5h6jZ82zVKjOaNQ0ifiLoLKHyW++Edpk2R++lfFlCc9V6DjjtjmnQj7w7UY/o
LFPwAGjmU+qlFKDksJateawPdo5w7zFuIaDTGcuDWirrOeNbpaWZEv03bHu960Jr
GM/qhD9sxl6H3+OiHm8uULAtTgnGUHQ/G2HSq0+Wi5i90Lfy8Bgy/Li5GwF7njB5
MiSlPmstUpaBZvGa+nDaCFCiit45MzU9siRzSyCxeD+WRPFHSFglV2oKtYBkyAEl
clkUSFz/boHO+xyZFKrG2815v4+yrTatqiEJHRa44aRQRK37jcE114Mg04KTizBG
RqaY1GgoAts5XjmCnqaJZy8UNQMZnFR7a2CKhk39tZtiZ06wGCVL0W6w2hGYiAps
g0wyA/Lz0Y2cMlExqK5EvBHbC5TNiAFvfh+GGzjUa+MtSh6z4wQn1ym5KfReuu4Z
ojSp6qAYWlEexYOswiDXm/Nz7njQ/Ifw+mcv8en0zsNdpRBvMuzFH1V2QUGv7uVX
g8CfK4bGQbhx+ZExH6+qc52Jl8v2qZ9WrbtDqu0GJO88+jPHq44L/ugVIh+Mnflc
FsbjnnVlDtsPaK/Xcp+lOyYwd3TqO2zDyr8mPvdGBX0AoTKcjizKceRzNpqG0FRP
Wtw/Mp37LXkGtl5jVKWiIRnsNM5r7FPCPaefBQss7ZciL/2+9xq/0nldxCxNUCcz
tTIHDQ2eSM5jlN6gjFB6eFuHTYzFqVTffvvk2pSh0ipsxvsxLdsAeezIJ7B5PQ8Y
o5QMnRUp8jakdHmoMXb2VdkEZQcaEuxtMFnt3dL03+D6Ze0J5tSR9atJOgoDXDKU
DEEnparq3loQc23E36mzv4E9NHnxzebcnNo11zEuXJ/oNRWAr34jUoYR4LQRvkwP
aLn+8ja42FhdGi0zEpFZeNFPYQ7NV+fsO1d2Jq9c6WhQVNVr55cy43PLfgH+A3sQ
xu+Mv5lYvxUDncDB1F4qUI1DwFmMEIHV0K3tp11SB7c0oGm1JcAUkq0lmxdunEYF
2foVAQsgfAFExdqQtSK+rEDbfyi6IOj3vD7KWqcDnY8wel7wTGhehU3Ik+ZSEunq
VD4vfAm6QklEyIXdrgD5PtNdrkkECUxtfacWLDTaIkCik8w0aaWbVDiBiadqTPfa
B2g4n/OEzI9MX81VKXUXlSWI+Rh75Iae6pwbmq4JDKqd38qNzy4vY1cuD+WigveB
nITxciO1FWPTkRNdFbm/2kNJ7Vlqte+pRsUT8NMVeIlD1YAE8gCTMvazpyOhdiGz
itwWjxrBayoZTdkBbAO7zq9ZJFiCJwX4rQibWiLh2RPIgbPd6kUSKJpVuXb8kjNW
a0GGReWMQuWC355W43DSSmwjQtbivaqXmoygSWxE/h4FMDkMvsJ4PjBUAXPjo3FW
YgLCA/sGR1CIAAubg4mZvHdSPIOSf7XDevslJrUQSg4NlvdhogvDgw8QqiX/8hsw
wPC+Shy70JCCYoqQMXLg8LzKRZsYUBAi+pN2jqNP2eHHkPt/UXwkjffmuIsZMeIR
X/Ec8sRepYlggTIhh50fFs41YdhRXT0lz6PFUiQRD7E9HTG89BPEfv2fp7okISwH
XysjZtl+n1GZt9nHBEIdRXRuI7Ds5Ii03vKQ+CvR7AXCFWpK1JSRlRSBK7ru0se7
BOu9IWImVH3cOI2Ol3dfyR3ImKaLIJ6ko5jJsh7VhnpHfQf0kXMKzQ/sRvkNuUIo
hHChSBMluvD2fomll33MKTnRCLMbKg0AGekcGfp/zSPX+Zxo1s6k7MpUGbHoRNT2
06QLkQrAaoiLGNwPxbYtv87Zs6J+OwLHN8/BHW+DgNaigP7dNDFbHx9dNrwvIWu4
mxmpWnISJ+ooCv8K3Hmude1QZ28iHMRxzRX36tYai+/Sn1Aca5fTn3NfZiaGvcni
z3UPYn+1FOvMb6eKoATOjYDEP5nRpFeyNUHfCiidfh6NRpq06iLCo9jSTCrFLR9E
ABdBmq1UqEXCi7XQo5B/I7A7Jj1TB+5QKn7Tqqa2J746wamdDhPVL20CyB6v9hYu
MWTmAvZ0ftMsLClDIhprt7dyVoaQw4DzsUa/Pzxgt6YMORUHCmUTe+o5CHcHvyVl
Ckeg3NmMN2xz5c4kdHXUso4tiNFKzHGu+Lw/e4KDNuT2ohyK9mykwWgnNx373ku5
jq/P49j+eH+UFnRv75scDnjEmyXJlHY04nCELJ1NnliAcpmlcoct5wJ+W0ILYL3s
g8XzpEB2KDA8TlgUbaNFYFp3cALcnDX2KGVENNeiXGTD9uu5ZrSfD+gZI81cLUTI
8hgyPgZ2i2Gd93JOWCoYMaCRtPixxobH808YPkdlrLfYO4PjH+7jYET4ChvttOmj
E0mgpfWJZd5dxjWNTYyRCz0A0MXdPSXZ5LxNSZtt+2XeZVKWIA9Udyzz7J1tNSmN
48fwaBe4k+wbcgPeXJTAiW7u+jiYdRBFT3MBzvWuhDKByfYAhiAct76B9shQOJ8v
w2XGuTxKVHEPrLmwTjKC7g6NOtxAdc38ihRVLv1SlbFPv0tQYPtp5xFi61d4CdVa
UnAeYkOobLTMwAhMNE9G0z+zTQOXVG4L6WuKdQuEybje39PsKLh2hbqnwpbA0Y4s
9jqmSlP88x6egSDz94IH3ltfdVDiWNoXW4haXBsWW6c4FS6T/fcnBcaxY+qgUiPc
qEKbeWT1TJBbX3oKpVQHjpKGrD2jqEHULVLRvk106gPvUNuicI16dtv78EFoUF+W
+QhWUjXTXbsaUzfO0TggZv6ONse54oM4R022BlOod4FE1bUhNGv/WoEzx94gc+cB
6Ay53spepYw0XOBgw2xBVk1bldOqBGkPiZ/vtgjOCKJSifAYVVvx5OuUmR63p3rt
JUnHDnQWEkgOUJDYkVcKMn7/ZXDkBp9H+lLKiics79t8XMDnSV05jFVV3hZv53UH
yFlOb9GP2lgym+/9O3e3rW0GD0YvK77Ev2+6lkae/oEdxrzjbA8k0LOQ6FwcgPag
79fdSwVr1PlxlT1MGRzJrNSbUokhX1SV6zmwNgHiB0COMUtIlt1LTvlsQnKWdo5U
PiZFmUJxGx76WUqBqrB8pAEpvaz0e4Y6snINka6RFfY1vS1n7YU0gwYqCa1vOg2L
/t6nFJ5B0MBywa4E73hbFIAm3sYihkdK7y94l5e9pInwWXcYPzQfLTxODGHFeTjr
w0msV5dYFD4fd1kUPF/WsxWV0OW08nVXT9Br+qcfSJ1qztdotxsM97OzhGfcPolX
pjAhd/sGtGFljL+mZUJ2Hy2zuWBpku3YpNlUqRHcxqXTazw4rY6rsrNrvCDlhsly
tk0TuCAku3wmlIBTtCebhgXjAPAhzqGlReE/8ri4KfQkQdHdp/8ej4bzDKxgKOHG
Pnw/TIkuEGrobz9Q/qjFCFMXrnrjH0Vxv+7A9in0+/nMPvxnxChc2e6zOv2roXB5
3wb0DAS96r5zWwOLqSKrvGy688TzKUfAVpM4mRUqOzrRfbRJJZ+C/uVEz8DX4HDg
yqelR4AFTwYRZnpySukVVx+z5fPe/ZodPwBD8Slts7+DsaehPwhvrgjTeCZWnZ9x
d4u2xutaiUiREp/nT8xdL46poVWeIB2h55YNYAOYlnBt7tDXk4xXh8bdAi7V8YgE
DMWjNXDloWqZ8gk2yw73DpZ4GKDyw0Etaeamz1ECBEL2WF5izqhK4jmEoiuvuWlM
g0dg0Hd3WK+Zo0M4yyZzyqUlEw2UO6A5Zzzuc2cgdTNMGdAz38+aa7qCqCMWJqQ6
1bLr0wBsfog5Q8HbZ8Ztbw2PSwrE60PF300+ifHcSVQy8d1RM41za1ZjNak6vDwS
qtg9T4jkMhAhF0RlBaCT0pB0tiZ7OoKdTWIrpwYZNcroErnI0eHxkqJeoxF7SX6Y
ceiRm9NYlt4tSa/H+IqIywqzFVWx68mganI1OlZQA00Ek43Yc5vHxflC+Czzm+1i
NI1zIEXpOJND5Jb6yF5YcQsGiaBjb24idD0NfIvoNaBM9XYaNr6bFbtfxWFBdVcI
8kHj2eNmMSSXpiiRYL2LkOTeaHTL0WelYLh/FEKSbF761Ah5zIQrIGI1Gl0gR5J6
qREuBksp9vuxxYjXUgE1VOrFSQfeJCX2WPUipU4TIlVpEsdtlIq/Yn9Ff4LF+x82
x2Gn2Y06Fxv7YvphwKEV0L71FJ/yvSIGeZz4F9BqUsPM4Xb+/iKxn7r+dnpgyDUG
HUvZIIQD7m0NthPhDT4thla4odQ5avetmlERBlC8ivFk2C1CBKXB87XBdrJE5B2X
rta4bchjKEucWJHsE4nUubx6VYwsWqKADfb1yYCStwNGxCSyVR/Fgzydk1A+fo3m
yenVYOD6dtwUosrNUdpJEFOak35Dcz1/GgDfUDK9MlP8lMmL3IDr700A5s/sDvv+
CS3KRw4r8V6xdJlTvokScr8+3zPDKvOHokNvxRcudoUgNsHKcY13JSyS55/4f/os
S9SbE0/Ws5u6fTpEMhA4i2l7Ai8ERlQBzIMJH9c//EMJocDNDWH2/939Ux3MrJ2G
WaQrHjXGHtJaR3txtjEqTbLmDEtarNAQkwqsxK7tVQpUfsKEA0rvstkKyAyazhCQ
jCGC5rrWROZXtMIvt6OGCOjKKUsLIjj3r6WSp5j7eVQ7zeMq60cdkeqf+MzfMlef
8HYpsd0WQw8EutsL5ZVKZOh+pFGtOVnw5OVsRioiBkyvEPQJ4oMIqW/gGuX+YIdn
YfTTfp+8AFZ62G305IjtggDvLh9W7dVRpZd2HYw7Ea1/m6Sd75ozKomCIlcXbULB
G664ekXEBa4iWCU99USeqHERKDO6NrwzNo8wfxXImZD9z0hc7EMvwuCbRKTuKV7C
KNq7LMrZjjICDrhX1nHnoyB7Vpo9xLzVi5c8uFAQAWp0RWuxgRf6RjILg9Wg5XBy
OiIzPAU3kxZpQqqqgra7S3efGxyWiOarf6JTvcZr/Tz1JTgWAcFJdvDKXnDgtz05
B3ETTJ3477+qtBkQeV3KJkboCK7X93vjsQOwXa+sDQAhlWbhuYw13zPhQIx5KC5w
qHkIb9i0y8pout5TK6UUE+Slq1QlR7npsxLOSoCeMJtSL2yxOSR4JVI11ySXBTP0
EZ8EhvMJR1wAhTUFfcfC+YXrWUNHeLUNBfvGG1BoWlZLxsGo6QW/MNjUW17hs7dA
+818HfCd/IKa5gsM6JVSjK+QhPQCUrNOFG36uFCb/Zr01aGfH6cObRkbNazYLXas
zVvt4t9S6+Lg2B88aq0UXdSRdTQAkkzJNiU19ucZX/QcyD64MniV2VcqZ8UfHzEw
Zk3thLMiKky96qMwom4f+nicvu0pYUYUPWXn01c9i22SMklb2CXM85gu1kp7Wci1
cYzHiqtapbYPVKFxnR+VOivfxj2ZNz9NOrIJUoDVlUAXn0YhDyPtVnMXTcZS/zq5
7uqo+rME8iI4ow1ib584zpR+QFdBTIfpMYnCKI6hs/OtwaD4boxYhdzLhwaeiV1T
13Qkjpo3wI6j0wytJ7UqFGLzhR4huDvTCHb43c0UQHsyDqgrVxYlfoa1FVWQ0pZc
gz0NTmgOk0I5jYseOmg8fsKCJAan4REqNRxiqhW+y8tJIJyqrq8IR6gPzebP6X0x
yz39tfaqX3pYmswxc3sv0CXzepEmojESrT+Z6kjHk25lAnpGrW8j0MwmsdU5bVh8
aD0mlQeFeBaquuELzMG3WSZkHPwkhvJmCpG7psIQbhNCIltLNBlOCb0xQOI/Acoy
LPfwZNfy8GVnedB4ENgAzXfwn8hBUNNcSC9bJBAmMUk0Ei1qGihWWStBG/alyXUy
R9Erw6vLEMAnYdykbrf6evJc/J7/8jaAr66aP+yAUQU0VixqUfXuBx6hKYRYU3bT
Pd88z49v8ix+TXMEOr9AAbLNQQ+DTnTMknTx+YorIc63IMA2Jt4SIzFBZmHePnus
IxeXy/ZXKkfWaRdEeJobC7YC5eCuIRSUgulBq7hEo+J3S9dlY8V8xE41rw0A/fmL
jGXq1khu4gM9dTchHqOLITD5x62nqylD3+5qLrBeQuHHBNuVwmEJCm4AaWrjmVgX
M/i385XbMWdYGGhc6XYeUbaaXOGD1JE3VrcvzbEcQxGmzgyBIoNykk/0X6okxwIs
kdIt2D9vJ6EGlXn2/++bJhyhsfFWyAixMX3cwY/xJUDj+ICYJeZcz7tUxIuEHRYH
BOJ/KRq1O6lMoLGfpia+pfjHTzYml/whNUtsRDSjwvkbj8SdiKO4tX5T3vunjOCe
mKl5mX+vpjn4WT3ICsQccsROjuopa3WbBBAnvdg10u8J2rJE/+2Xwc4bOlojlFRW
iawVj8fNjX4PImQJaOeQHGqReE1WM9k36xETmugcSEPsTQ5BzrYw8E0cqI1LmNC5
yh4XewLiN+SgXZRoQUM/2Kpmjf5dCrhyldXIF6f2n9wdSxWUGzNfv2xG6ff52uo9
RHE0ix3NfaKkKcHJv6/QlkUE5de/CuFn6WjUmlUGAxPieKpy3hbfclNiJ4NmWdWl
c06iUTysrZBo3gdRCaNOtRhn6qKVZVo+tzRKKnHtkkBojMhtSWOwQJTLj+t/lFUH
WHFRWL2T402uv6oV/C9k5VhvOLtDuVLp/s4FYIyl98knGQI9eESZ/NjjGAiPNCwN
yjP9UKas5rdrgroESdRyoCYLCIzEpPX1/COUetNy7a+N4cJATmarrH412GmD7G1a
Fs8E1qztYciDpYRKbkF1eDlbL9PODGA4VZDYM8YJhlEvE173VbEd325A8rxWtPv5
LjWQdoktBPh20IhhcE5yG452OxnikSev5g32f2pf+i7d+GVh/SWmEKkBMekwP/gc
F6pLnbbqEjU5XLtiWFa9KepcClcTDw2JoVBVEu2TXVjFDwIxtjc0B+CYVQX8+Qyg
FWbavbo1S5B0G7iUIGtp+BV0XwtqowgTVkxoZ4vHZeKnH2XfjuWkSOzpxF3KJJJi
AkVWggxYluw4eIgieMQ/rO/72w9lKFAx2sUQ12it2xaE5/uvrs3tRtQZy9mCM8GZ
Nx21IDZ8AujJ1GzqWAAqZFIdKL99b1uG7VlCsub/qwN/NM0j1RVVOZeZhxfwSrNI
bqjG/dpQf/kzEpc1uIN5ggJJ73Gj8MU8GTv2h+yfRcSma5prDo29KDpUEZp2IktL
HMvWWtIiWvZYtYbKnYLp2xQsyQJztFJRILLlkCTrVmS8ub6YzbX0CabYokq/RSSW
rkUtTq7KsOD4Y+7QoMJUIq+aXku0rPADPagRk5GH+JVKIuDaoKaDU5QOrddgS0f9
vN8XYqRaXwMZVfzNITGXLPG3C1gh+BdoQT6NCnbMxeTFDAi9bGVg9Sgj0YylIese
4DYLy7YO+pqQMYwfGK03qYh4SpnxTXPoYLhAdDHHl56Z6NLRRs2lfB8AgRhXI/0W
NhHzbQY2/K228hpxd3kf81L1AtRZ8xkZ5vYVx53mczA4Wclg1NZ/wX4sa+kNC6+m
0DC61ZEh8SQFtISG4e6R8B5wzXAgJ5sDbOWDICZ00h0G7LbAA1sjimPLythaDk8Q
XI2Cyq1pCQpQRNPsuHWub6TNrJFMbOu+EeygqrppeNlzG5xj5j3CIQmzWPWveRKk
F5DKzZR2lL6Mzd5DoHbuoL5I1CATwxX3tpE6fEsH2+IH3pZ9iZ2Be36UE5D77+XM
j7VAkb+9MrbX4+1/EhAORAZrATaF8j6NsqfWbILxi6zCpT8YX0tGl37OXQvW+HGL
ZOe3OltoA0xNhrHHxVKG6RppA5oiuJcICzv6Jw3G3HB8woDOPBfM5JEez9Q1jV4y
MArzJof0m3Kycm+gJS50gqEeoecQxZteBW7aj+qEx/cJhc+Uz30ZxEm5O1lZ/lEW
yiLZYDQ7dCNpMVEHEVIefytSk/E+txXj9bYpRbV7BpxmRC+5CFwvA0ti+i9VUrT8
djKpNmRJycnJsOCcYIrJiyEgb5ABslC7nyOW/bmk9pxCT3HhO6RKvIsEjkwd8nWU
htUTReDT9qLYPqI4UCU6C0roEKiX6POpBsahsxbINi9pbIV4poOFB8GkdySfSugq
JyyWgHW2KT+LjdLfEJtdLNM+K1HxoUomzLh1pITfUUNFc8Z4FjYpMJy7tFEdgBiN
Z9hD5ki47NOA2eiLsCtopJKUdamlQ7ZYvLBksMF5RZq38NIbdi1frq1ELT5U0tZA
obAFDcupzjTHrSChzrpkr54bvNZWEfNJbH3oHZWzpjpyKr5MlVTNkJdWjWID8WWO
6wxV+LUX1jWyHwiAljS43CUwmmDyLOPXuTcfl7CkQsXNLq21C+gO2i+MvpCvl+cC
5MEHB+ta9Hs67np1TCfBhRkzC8WtxAplzTKUjrAWo4JwaF9RMqE8Iaejd6FvpNPZ
tX06Pe0uzKii87QaG7EDWDj7suLPZ0GsrB4bfsoH5zS1+QHWdslM796UC6b4In8v
6aAbyHYImStrafpMMMPkaIheOZmar9vCktwAhKVzbvYJVjSJhI5Okvddybh75j9f
9AXD8/EtGkn8BtxE/QZqYcfiP+/RfUDLKK449SqOCbTGMrz/Lajf2iS9iGXuHc5d
Za440+OXkSwBzS1engw0xQ784y8/U+wAuIBJvirXGj+F0Wmm8Vu/mNJa/Y2WXxtZ
94oK/qjZ5Te4cpkAav8a5spMW9nGvC7cJL9/NzIvHGOSAzK76QS7nxNn3MsHaqCm
hCCG0PYPWItZl3yqO01kwGcK4N/PLdNwN4Pe1J7rFL9VlVgITVmzFvG+pvvuL/ax
OrFLgg/MP8/wd6kIWHKakVjjkODmNnd1XQBap3pb349H7zu1emHGxbxbK9G3I7Xh
aA9HX7ocqtpY1AIH2EjMh76HtjiUfqWiEmym/h1VYVV60fbUT0OVmCsfsSXPMuYE
8EJy0sFvOr1Ccs0ymvnRP1vcjUWyePkrGQ47Ga6gFfirt0rfe0Rf8vTzllzZXlEM
1HYBIY+PxBRnWmOh39TIMwlSCWsiAmhQwbJ1ctl8CUUc2Wlt/pUznwg9k0hlPYw8
HUpETo97eEvRdlqgWtVHkw4RCISAzCFeCo31ePFihuHW3eAaufLIOCSieeCoaD8E
Y3Gmu2BSy8BKYEXEIOdVBEQGL4jNakFwi5g6i8dZeacCvfd+2jB0xgoC/f095oIK
vqYwamk8yp/NNq/iayI8pNzmPQcVeWD8NJl35K+dptuPi1qVa9GSSaMgsaaOyFJo
FDpogLxZBoWUGNV7jeDoPfvp2fEH3s69QRt2QgtqvlgPiNhDYzJkUbaGq2g22lqL
EyerNHD/d+9cVI7T0IeXoAZaLfndG/K2OsUBQa30yeyqKXjnl/87+su1DIDvibpF
T55F9jgc/+QLbvLbqDGmVpqCR75sDhShTPZeFCPocrRvjmuCLx4yHifK5BszCJMg
chFyEoPHiSs2T87peefzrRP+PsCAROuuhRq5YYx7LZbV75t1O2zlllqiHPLxhq+p
siig0u4Dn1lIXytKm+RSfWlscjCy0Doml3RVvo+GHqkK0yF3PMq7sKD1qcVkaM46
cjby7My6/635qPyR/3VR9g6n/ticFpg8kY87YqV/FwWA6V+yqlTFrKuYAzPVILnN
CXiSOlOyePhBsNR9StTZWBm0Fes8zKGc+FswpxBILffPvdU1EBzNTb1DpBh+ob5/
nt6OMd5T1SUJKFrehaqoMSbqgz2IKKgdVUy8AwDM8tyjWTBrOvJ5hjIUY7vLmuvX
5zbRHs9GdoD9KMkAH/vP+vK7w4PMbzTXtyO0YWb2L0VwIRe6nmk6r4DJeGXzkT9X
xxEczrX9DDAju+xqE4hZ7/Bi6EpFSeuC+82nq2TrwvVnb/oSXzRPbwEZ9CDvPzLe
2reYoOZV4vaUBb9F3zFMrillkEilOIFIVpLFeLCf5ygIM6+QVOe7SDzUJFGf4vwE
uT/n/GOWd3WGe6eO6u4O5CRK2gdw6bQGFEWRSbBgc2d5doF54gC54rPVT1Zjtflw
Jpi3TvZ/wHXByAVqQTv3+Ml2IkzLV/V5K7mOZ6ypOtjecqeaYPoDAiVW0io+jfEV
X/t0JDblB25+00PGBISMoF39Jpvcx6ZiG0VUg+3xV5Ltzq4l/zuirdXcUicQZdve
vPv/Ny6747s4PqPMHaaGJVgq/Jobc3bnyFF9OJJyAPMALI+PSs6tU4u0shaKMDDK
jy/TBMCgdyAfwNPJkrwuCrHUnpyujwB2eAFkHFYDR3GvktP0LHTvwlwmRyKsP+P/
u9Lp0yfX8T9NYd8lVY9F+pmUyLWYtJ+m1OEgBjLjk6oD/f14lPDa7QCUzCJDqDM6
38CmdrHz+1NhNfD3DxzSkk7U8y7GKeN+MIer3j9ApJGBGntPW81GQB42AIFNWhFH
xQps5ktj+EXYg0eQYh08TrRF/y/iDc0l4yiZtc7VvjmCIjd74k+hWszZR1TI7+y8
Kcreob8NbCzPgDV+08c0Yxj+TQz6nCi361TfNM0/eY4VnaSd+IdKIVecb7lklQzP
B7PZLb5cfdVDTcHQ/SDWnuGfWbShcrs7c2w87z7Ppshb2oHJItuqMISUtyVVKumf
FMBo0Rm3EbSH/eCt8GRL0WsJNib3MVe01PNIfEDz99o68O8aQ4oyvv4fk/dCakFJ
cAzzxLlTn/pSMLLHuR3C7CYOTrSLQwXhIEJ1NTORYZt3k35lL7m6lE9EGhsWyCNC
Q0DW9GdEXUYj/FEJR3P3452nkoZPoEmGLaLBQ7bBnvZEg36Spop8xKG/wEsVaItT
V7oDtCffBpA7ytyfBTFAo58XiHQ6gPx9THRWZM3/YRXnSVO3kQx/9tC/IqsA31Yr
fuuj9NBfxSgpDOEy2YZKH4yLv1GIX+ns7o2clZZvtyaY81CFgli5QXYnHGDJc5+y
0ZzRtYoryZpgEVU9FkG3rZFywc8IsUC9hOQtYE4NVwuBEREN+ri3zGnmFNTgjN9G
1FfYZ2i+ajGBVy5lPe53MrP5jHWNodS5kddo5lZOCpYGMjqBIdf/p7IzSkvrk5Ah
QvtJSgHowSZfHhCeWouDG4pf2Yx+QZ3mZ1IqsXQcYqsOa3R0tr8UHx5TlnsZt/sP
hihOKBUR7dsgOPa/c+TK9OOZsxM0Luh/tGDkSzuZoOPSKk96X6qXmewV951h6Fx1
DObaO7stiMvgfbBaWre8JdXH9eAKFB1p/egzD/ADp9jgjlXHed63fYr9OnYRVfkW
kTu7ghfjFw9u9lM2dfycUcWgWPD/5M2nAe+gZM1QcirsMLmtaDEJGYczgTENy+VS
xT6PHkCorNtA+Cn4Ahvvn9nabNwLjqDFGgh7cDaGQykmIWTa3gZw73uAHT/6Juxk
JxbhFxtY6tsFJosttDo+V5x9KyeNRrMbKFFETBfV4fCS4IHxVdH/0SrBU2pp1wt9
POz9fD20luodA6Unl7sQlJ3/y7u2yuSdcmGFuVPHkNzEA3uHN4Bt8I9zA/Ur+1QD
tw6zV/wgufYzWmXOKb4QKBUsn+WbSf1EeN8sEYDEVOWa79D2Mo2zTSMcY3KOS/md
jQPy7hUQwPaN0EAm+zDan6kRz8g1lvi0J2oN4GuhyXUz/fiCcoV73k2e5FnVsJFh
OIQRJKrfWnzGIxfRyFAAzwVqVAHNmFcfMDDralwb4IcXVlLzov8zQUjYdc6cUfUB
C5ZNS+lDy0WCkAZKdNDQgvR3pl3t2JyfJ1f1jr/AkaTRpLutJ5FChHDQrs+wH7yz
5ixMoQezhl4kAdKiNRd5ryNHdP6LJt7HT35xyoMhpExxlbfUgQ7sRwUskORjKnb7
/6oRS2Cq1KplaXcetgcB2Fv2SPUkE/n5aZT/GBiZTTtzQsrMczZLdMBf0m3VWo5K
mVXBQlCH/TmBO3nXSpKYQgbdYjE1ctXbCuexdQw1ElFBqS0woFRtvG6J8PXbz+2p
hbXQ78MOMu6AY+MFVvDkU5iKbf56gpSgBhHIv70cJhZTeSYOZnp7HXa1DeE6kPrh
ZZOiWzVKlBfQrdGdrIteFF4lu6FtvOqKcw9Z78sS7SceFEjj+r4hZQDZaXHB0nXj
83pKBwxAcz54LjVFR0pD/eUcSy9vi28jEBWIUCKe0FsSp2mTOu6zdIMOhlxjKtBX
rbsZVzMefzfKkjJRArS3cDz39pSx/WR/jK8p/6KVc3Qqmf7/7Hgf8+GJkNUmcSoD
UpGTb+kEhNzXvagMAd8mXVYG92fZwP+migRDimZblCqcVk2UWHgMFTjgQlx7rcYz
UwICpbTte2gj2+jaLswgx7EhoiBaPmlGlJ0jtfFsGztahLSqEBSeD8SAyP1G93Zp
FJautPDYmfHzkoW5EQmz8s0muv9MZKHngdc7rvpaEkBTYExXkS8HCs/f/QTdtTmF
CId/ahoEjhHAtIqtd7y+SedbE8MWP9oMEEv2jH3qpD3Tzdm5p2plXn/cHHCT9Icf
Rzgr1tSqiTge52+bvLDqpR9WK1YXJiYPB7WtLIJYHE9/uVIuCK/wwUysnmqZH6oI
UeJUaH7UgF/wJ5L0hpyyGOw/kbS5KlF+Wl11JxJEb70oEXFi0j5liJxx5ZvgA6Yp
NmtCKu5imyj6bytbZ3WnxyX+69NHXGBcHEcm++ADg4inulV/jBDh2bRpaj0Y1s3f
MtCa8ImAhoUdQatVJ867qNWjSWZ3id5iup7VLglNYra/VNbaxbgjS6jd0CR0rkuE
XdIl3OuU9MzYG3MHRABRAdqxkLWsdOdng4yzh/Rgo4TOQloiBkfiowmLclmtGTlV
jS9jSuTYutngl/m12ys8IZL1LiwedD4ffUfl50HXG/y011OSbrveP7cXuP8LbW/A
AbPaLvwQReVM9y0pV34/7QAkC2kWwP/U4FcQI9ocZoXuDhUuHmZopqDyDIJ3YpJn
pXzrosliBcbp7kS/KUIEvnxqewz93CH4d0XoosK69wJW7oJZXlpFqdsHL/DjlddU
IknQNAX0+4HV1M6LpBpOrO8tr/aXhJ+i+HJW/Du+emjKN9U0iCZPmll14oj+6RLc
AE7fJwiva+8lFVkZ9/dedt0MILUKt79XHE2pSAdVDoTOJUduajFfp41ylHNZY4NJ
+z04Y5PNw4v4uBRCeZK0PWlNWUWjMEalW1XKs7Nd8Nzi9wwlqd4HKQ5pLU/ylNHU
Q49g0ZsKRahpRr83zjf9o67/34CeKUF6CLl/FBx9TsTvL/Z6xsGQj6P3J/EiosAs
U3koDGjzTSfCf79pjdxEIyxVfSlS7ca6p1/AMNGQWZSBP9oX/0j2idWMyslNF+W8
Jr1ZGPG+t/JGUCnwKU29AIxPVG9OPzCjfm8ZgxPc60zPaSFcHomOFGRTyV+lePWJ
LKnjEXW42K92jhsE94DknZEEEAGGoihNZzQKysWsy9PDAj/S5ROBV5OSvDFZoPHq
IvJZotkcwHMEK7Kh6S0E6Hazvn6IudogovLQqVw1AiELGhEcYjNaKU1fV5gFr65A
RXp3rdxapUZqNVQV7l62yS5IbChAJ6mYSEjmX6YvPTppFMjuvRsD/UBon8pkwJ/F
LO0t2PrGP5H86GrG4oSVN01UKOeSMWLWb2Pp3Hm7sGe0P9/olBo8TRjeDCvwCMFX
VbTJXpTg86d4uKSRC+FD2n6s5+NdQZSqF8tcaTUwr2MIAuzRz2mNGAEBM9Z4FDxy
QOdOyn8f3jEwUY7a90+mmGX3nZgaR9NKazt3aBJXw13KvhbqbGhcoFME11ZUQoYe
7GFxaF9m11lPcA4M/DB/Y6oVdd7NOMEu2TILCzmmRz7DBpReuE7ccRvG+w1w3h3q
ml4UGTL6cmDQBuw3Bt+85AHT6zm96uXSrSf26bQA8jvjGJyF3Juw9vS+x19m1kqh
Bzk+zF8jI3vy7hyNIiE7/uBaAzmL8qtTTsjMW5pizKyJBWnz25yPUi0a/9Eq5p5S
PIWHrGBLparWaWdQrzpu0R1vata8IOSWMd/EWpcZRP7ZHeUjRhAe0R+k1+/JTm21
kjXa2saOOFBGQw1Ag+yKxe0H1wXOq7vI+0XUHYp3jdpr74Mu/ZAGx1pUWkrXpRpH
w/TxxBjQBZjQKzVncgWz643lOtLS96HIutFduJG7NK6dERbc9S1A2R07Xr2Hqg73
k1ofG4lpF0IXTibXRD4jn6uDVWh8LUqEFbkFEWAm74kBiwBgA/R1zlZUvXao5ukO
e2zDelDDAWwS3OBIack72lXP72s1GL5u0aInqSuAofCFCwr45fXiqC3xxARoQOAN
gOPMDXkU1XJXBV8Nwd6SNTWqhI8K93ECJM8J0FSPpAvD0bDkVJVZDsvlwOd0KYXB
b+3+Q89I9/C/WdwbAj4F4Bmputgx6rF//3oFl4Xs1+oZx0HmrM9mBFJnD28jhsoG
Vq15QQCbNErjh9PGqZsnLi5lYKioTzlHOHkn1Z5oR3lo/PjIU557nCZStRYgM+pN
JiAhRMBqmkgSUvKR3dguxRZEQN04ybUa0DYN335eYpcjVbcko/XpEO8ZUDC/Xxg4
Yo0UaPtlQGJ3gl9vff5QKF9d6WlHG0aYamk8U6m7NkwaFGrPsj5CZxnQ/NX1KpBP
RU/Tg4omGRiqrtjox79s6AMtz8QBdxpv9/MR4zrUnqXAAEa7bps2AaRmDH2QH1Ku
Kf4DCNdn6tTgFDwf5rop7DQhQVQEXpMYfMklOsvVfpF8EQE9GGLYzYSIKUfzn4Bx
ho5TJ5EBj3Aff3UMp7A9A0yqb0yKD4ZELpgAMYP61kzftU/2LdreTEIr3eIunrSp
tokThrY1ZApKF9LwEoqjJtxPJ1HalvAGXS9zEv5RPwse1CFjM4Y82pmzDmJqzsKY
s0DIiYMQxpLA2EFGMr5H8foQcNlmJrep3HPX/81/5BQKiOuRDUsw2FhULn/OWWsq
2OMzBTsHN5ag7HLHIfLUJmst8v8FUO85NAtf8w+NFaIQQe6dvxK2mlVysu4SoU82
nDO5i8gVls7yOW5ECSQqC7eZ+P0H0qtSjTJCx/WRPaIzP6r49uY2CjIYyHbXaPtc
chGJbq+HuE7A2rQe8XjGjpQ5Iwzz+HMJY4HmJKMPdgRCBfTzDMutvveBHb5ZKWu/
T/XGIW06NW+DNNKtcDPHCTAQrbxI/XM87m9UY6m9uyw6HVXSTqW153jhchpC0Ruu
rwAzPUayonwGzSd0kV9Xt1wG/l2OqWUZad8lVX80aal6Hj6Vy92kb7oKIX5QU+Z5
aU9xOgsjzW2sjtpYONAcjr/5Ke0r3jWb5oAu7qiuDOD9qOpWQE7fjTtrQxcyYmQR
41TyzqGI7rvotglqT8NXoPS2mP6XoRrHQbg04ypRqK9haZ5JzbkLJehT/YwwEEQx
Ia9F5/0nxs46fV57vGOlFgWdHlXP74iLjxEO7acL12cFOAeZuOItWGqWT3DbkDwt
aXCi7NdncYQ/xZZV6FmZNvSaFS77RHZXylcRyeo1vZmZy9ALE0b+uHWMkidACU+5
LfQHbIZ+N4lmZdo184TcA9AC9BMYkBtqMlE1HdbD6Q8m9BDRXSaFrzfXeXoojDeF
wVuoA5HtKorHnRQ1wSh9q8WBVhVIegBo2ziSfOeQnP1s5D9bLxJ2LYFTX8FLNGbI
Vd3E9IiJYmsnTjHRYCPGUPUZ1Q4oslg0Z4JsKX0xhDb2eeI2JccrPs4AAZVl358e
ep9zyDnqZEuSMarNRyOlaKN5WsuL9V6SmOmc3ZpcCeMRHDr4QC7QSa9c1F31WT16
R9607rCfGYwJGm8APovtoBetqFc9deiAAOzWusNL9swTLTPx+lud7aR46eI5jm1s
MhS1acgmHBg/2GWwhKvil78kG8Qj0H7Qc01omadK6mntLb4T58/4CmNPyZE9fued
TxOXD+BThPnzjyiApuObkKW+gUM6R9VCvXJMyJAcyQxcFFHQ0tW0XUyH/RNaAMS0
YPgl9qrfSzxMMGEtGMSC+0PJDwd3aM7SMx+8+/eP7TlEXgWLsCYaOk3LoZNdCn6A
NNWp4evQa2IJPR+iBonfvZrVVF9C5mYQU8u1YiWyTn/kGFHwPnSw8w+d2rGExu1/
KFCW+bwd+8Lkn3QNAqFTc5qDbL84/9tGEGUZFygOTQ2TeWIFDJNIIBzA6RJdQ8la
Jy7pclQnD8geiZZY/tCHoS7q73neIe+vM3FZxfJBdaxIMHLYhFoXszG2WkvHvYiL
9+5KPMxoTr7UnyBhDiuRimY8EZ7mgmDxsHFgF6tJGFhbvd7AApK69N8bVP6FYeeH
6U4NmLZUSrLgQik9x94mb1XheUprK1qZLkYB4t3Kncii6Jgbwn5lr7FvC2rhqd7Z
+tYKvrxLO44OQMllh9nuSdI0qWvme9HztBhmQFzT/rSXPb3/UAx2R9218jISPCS8
tl3j0LHpTdmrS7/GIq97EtDtJovKXDcTsnvaCzMCKPOqTDLfEEUQ0pVPC3D0VLO9
W3H9A+eZxGBrzwa32oT5NL+6xkQYzi5q9JciBgSoscCdAkUSNzjNf2crp/3d2IUO
W1IziZife7BRu2MAEMHCpg4KLvdDiE1RVCGXC5FS5c90H56ZZkZGTy0lfk+ccANb
CK0pCJlT/vAYrUzeRC8HVzXSkcbFY3EAO0zxzqtYIU01+b6Oh+m6QxlHKiFE+a6x
hauXkLRDmjEbinUi5R819y3gRxSqSX3C9cecKRkcjJ1JfHg7Q8xmRmbU5YYJItjG
eCvZfupEtpiGmCgXLuzL/bOeoWl20W0ovqmmsJg3NrpEgP1UeBrnIhmhQjQ0qQxt
W6sjpAiKtffe+Ac2kNL7vRPAofgEmMGf5rdsLiSrFLbZcS9gaPGhMUvED7r+UDz1
8RU9ZXAsFcfqzynPH1LbRl4lYLrB+lqXJsCtm4/d7POHGd+AFOu+9XgbfQtI4qA3
ZeDh4peNCX+2Xkz4LjUjrRnhfb9aOOotqXZQiGr0Fcr3SZL7pvaYoNeS3kLdP2Ht
j6Ite22QpagLE8S0wq4j0Dw00sgMCent7dkapCJnlmPmLhyRL8xzqbgj2dk5yKqI
3frs7neNaE73qz9kMVxF3+Xxz3LBny1l4t3NynwKxRSo29D5uFdKYCpYprcZ6YDr
qKask8LPdgHhPgwAwMe1njdzCIq5SmierZnfIXehXYPHoVKkEL3jNHDqVq3Vek6U
6GKTEi3GwOOH+tNuVQ9wlz3hXslsrCrMp0809c1evGEW4QTYNrY0DBTyevWLrLpY
DLsJeS6jwTU8wNswY9V418B2ySipgtTXV1CocgLqM3RcJJ04xpWtrzD7qT+XIAcP
ZTZoY0Wq0J2DNQdHBdip7FKTrWZr8tab88SuFXaZImZBejTFv6ZPMEOo0uA2joz4
tTM3A7nqeQ9W0+Hlypt/HNFibeq0ANXiabut8aThHJq6oFsr6FeqRiPIDSL+H+u+
wRrmkfmH8u0tRoPw+Mx9LtLSKfzr2QUtHjGEdIMwbwCPbUOdLj/aALsyvHnllWRk
GsGKvNpcwt+Hu4zlp77HMyxkFzt5Ed5lpmTur7nhVhoByoIA2kIa6qU327WRirIZ
8YYsDKg32H20j7ZDTbZQl9xcZJza2axJLsyP7lUTRCsEQ3IKhOYTZDfGeihpvEVP
+NqpY45wIfR65V4yIpgXFIlpyyepyKN4YehyZFMgYKAmPA1vR2+1HrQB3XDNYomO
yA0wL0vVFcTDIBGjYMI8O8xkEuli5KeOW3Cyz1odKGdcDAu7Cqpa6H7Hw71/ky1J
fJyw/g6Q1eKmjtUJ0ApLY6KjPwyFkhxnEgsaCsF8W94L/eR5LcKhr+Qua/+3lblQ
14C/S6BbzXZLBnpI0Y1nfBKxwO0vCJGPZe0ydGpXCZvCDSiWi1TsaSzXIkbJ32VC
t/GFNH/bQTpXracVBMZniY4GPzCnlD3XAEZ1aEyuLfbCH/GXN+SioiWrw5qUimXk
tS/7uk71foqml5Gs3c7CGurH5lXHmF6BTqPUESfKJItXeNikm9pJ/IWhQfH7rlHl
CA3XDoC66zcfy4klZCLegH676Cac7iSfmMpIgfHS+/kbYNwmjSdSIbafa2mlvR/D
EU/dg27YMZt8w60x54UklbFfr6B0J7lKyIDjDAKmH1DbAJcA1v1+wGSxd/gRkcFb
d86eqZ2jd6T900gmGVZQCANB69DqBg4y20R6g5KSKS1zn+9+0m2x8KucgbqPSo4K
5CGYjALsbrD1ylejDcO0Qc90/RcFqx8ZA3NQqm4lgc0KFM2q0H74LXvnNdz5WumH
EtfHYt3X/T+UrH7QOAa0sv0s3G1meZgmfYWJFq1yvbUELoCdB1GFwB4LZSAJHDiA
6o3zVe40bf5i0panvRVeXf3pPWzo0tNI/eX3aIMtd2u4toVJasm6mVi98CSb8ILK
zEZI2N7jVhCvtPBnyw0O2E3ANa1TmYGiL2jGQ4f0STSDZenRzdpJPNP2sqz+tH99
gkRr6QowhmRIHVYM8Jq3EOUEDdV+Ge4l+zJDRE/6X5eEumR0k6cfnUd7w/82CLBe
NAdPAlDOuxzAdBOE9QjYEchZstrSzLS0MQyqJfrZwPbOYry2hLeBpgX5rCEVai03
pVDemkb5nYUBIQzbeHo2AYxWqQm1+kB77h8wmc6CyTySMSUqiNBiuendmRh9Dg1B
jkSyetlZzBVAtPVLwC59/bQ6etZQw/ONIrAPOnJKVGkxBu1YUrjakwfxMC706NdC
nytzE03yw51rcmLPZQ2UC7WDqV1kW1KJsm4k7/vZ5l2YX67ZSaYBND+0UHCGvHfv
JWziKYu2Jsp/CLvrf8OjMZZQZzLqonCYS/7qvRjHRjo7w5Hh3Si+IWnWY6vfT8oH
gOS2vwfvtHnfdebjnvH1m8qoDmO+c1+fQl+Z9bRP/bKL5CxVkgcog3lcfuCVC8Ep
GBWJUXv8KQ+L0jwsbAcHzQGNKluQPjgli/jeauRUwCKSKrXtX+j7HpKEI8Y0EDYr
PuNLu9vUVZ26W29NsMAOemF3dxYrq4qjoWgkYY/DEYxjk6R0ir3vEjrMG9rhear0
it0cOGAZZhs/DDfRX8bARF84LgCXZ8QW/10R7z/rEMMgFR0oEq2VkCg+l8BaoRiL
RlR/qKrt/fbKh7WckYU/Wxqxdp6rpD1VXCfxA2NZGOYd4vk7/wulKWWi9Bm1dLeT
2oDv3LTySnUaZ/I1Kl/PMn1ojekW3EUSOXNAjO3bvu20aptZ6qg6AqooD1cWFNtx
nJlDgOU0DQjU8wtvMpCjSG3IGg5x5Oe5gZp9XcG8qr2UdOkRXw2Dq8ugw6JLAdQd
AjRXIsStShXrbdqgb91zJ3EWhnXc7sJJ++eV43wq90iyMU+inL7kEMHQZAR1s8JH
mTfg/2E/THzPSWMcRZS5BM7Aa5qAaOlsyiJHOkZx4LXe1/RHT6xVVAywPLNGpCXf
+otD4dVEjYOwRJBS2DJMJH5I9JLR8iURlyUcBFGfRUCsEKqsuoDTHoCF2Fei6jx4
/rGjK/M9NDdLM4uiOPpkibvIryjSwqX52yKZK/xGKzai7wdf5UuBf2PnbzNoTM7Q
tKNHjnA2ZttexAVezrf6bStghX2i2mzHC0Wen5sgVP5kCFf88+Qvj2T3SUfFNCEs
+WLHbfVhRJVX9CWLlFm8JTCWeACJGW0Xmphd68KQxFjFFKtYCHmO8G2EuuD/tzU3
N1fh0VU5RxLxYpNEPoCuzIWF7jcKhzDl37t/YJnJb5rBzwOvEyZJpeO/wm35FmrF
Sy7i6TdRnKp9zc9L7DLyovXWPCNnnAMQmTDWtQ3rqcyI8Zs7D+Nykjp8pPLkGNlk
XH3sS/yHhRYx71ppOu8SPzU2VVfRzFrsO3cqdvKmr4f20D9xFpJoJ3/Su02knSfe
qtO+zPFfdt8ysqYIfbf0Oh6Et5vPtHJGtvdEN+ULUEa0VLBjcBQ8rwrKN0jO4tjv
rOt3kuKul5W301pHNvC3SMcl4c+rdbENANx0+sFXeOb0mJ/LbcI+HsEn+wWnyqjC
36m5gWHuARuMRBByj5/mAM/WVliYxbWdVN2ZKg4jfUDnKvuk9B6m39dUBBaBHiHf
xibtkmo2vlY0qlrfnBCRO8ihMk81HXEvZ2P4KF9QH1ioklhMKaqKoTPcqy/5gtga
vgFtR4fgkfdITp+AehxPPxYh+uOdwlPmYKhl1KBjoCC5Z3hV6p5BzI+cdrbi2rqT
r9g5uLtuzh7iLl5u9J73VDvwQH/z70Lfi2F4n0ddU72pPUN/qS3PpDTg2t/dtzfP
Mwnq25l9PeK2yBmvFnbJK12dBIV5IcvAOHw3wQVC6myl421CLKrEtnIQJsgy8e5l
9RFyqhop+JUBbDvAbHsa5DQF07/DJcVeovYJZ0Kh98iTXq7cs4l9p8AYLF0QNdea
440pTmrCvoIwuDNtXdNrpeNNqoX1DWPZzM80cBGMfBKXVFoQte1TWI0+3Am27AsB
kfcwkqCpwR/fqdFMIJqPm5hGNqbyBQyLz6aZB56RYsAQb/LDrgJChuHId1vSxF83
TZaTXaE2FIBHMxt7rmPcMr0+ojROYdyRZOrWCjo2eWclDcSwnCOOn84PYMQha6FC
zHfk6fa7vp0BlMh9K3pH6XAGyuiw9O1GAPm2LHvOd63HCRc6/GZWNgzKnPkeKGrU
WJmc5Ad5HMzhigpXFjaKMFzPA4tk5AIoJzB4e0m6/iFwddMZyYJF6HHVK+F4GxqS
1bLMKKkNuiwCv0pSDku94kve5106Nt5xFFJFaTGuHE4+vnw1YsXB4oJ2W9SBT3Ks
ESRgvFwbEeYjQHsoVC/qEghfyPuEgq6EqDj9aSFB9v/2i1gnF7lqEhaAwLY9T4u7
/D64wjuztisE0Pyt/x8OhiOCg1wU/VXgnqVLXwAVdxa3PAHhzLcPsviwjPIFMHMc
mdujDoJ66kIASHduotBhkOkK6jUOebvULVxDugqqCPqempTJqpl5bKIa9ZHuPbq5
ATEt+GJHTfwiDy/rEQX5DSojvvpnSyQ9wDOLK0r2rvP6OJ3GG1sQvRwo1S8eBU6w
trYt0H+rh0T8Eeiyy9hZN/QugJhJW/jdyDNq4eJmzibHS2bBkbfqfrN39ck6rwEu
1+A66z3E9ePfvJgYq+iM76zEdEB/5RGdyyD2pGyXMlKGbbsbFIP6ab0K2m6M9Emf
1QycR9q8cZhiarYMJPkF25KxwHz5+ZvpDDINhrBvlFEQbKZ436tQItxoPNI48TpF
Pw/1kX51/LJixWkZQjNZse4yfHkYC6eQzSKsuuQ5P9ODLzhbY/W9hu5DHMWvHudm
wim4tAap4Q4R4oKbGgWN154aNAuGNCLEzceapPx/pWVy4N2QRcb3vTZxdDNoj/qY
bZj8yXgCD+YBX9i8B9aE6uNjemxOKyaZ5KUOTfyHEYW8ieRwv3lIDXaFq2kL1CQE
NMOZTzDdMZJoW+JenGMCtqJ+y9nlbAIzGiBfrJA8pnTeN8NWCOm/HVfJfykM7Ggs
aeDXtn4WV12QTnkEOt8SlOH662h9gH8LhtWRcAwefWFc3ERLQemSZ+0KnrCtv3qy
Zh6UiZGbOU+aGvXW2bdDUkYTepFnMA7guzgirhPyOCoxn/PNURn9YLhMz3xxYzoY
51EUd0B3Df+YG8uB0Q5NvMCugfcD8ziAHyjvNqAPd9fMz9fh/sPh2PAEdhbBrTJ4
gW2q1o5WiTqab5kcft6pVtpRrO5u9Ei6memMfie4Itz+0T1NXKDvwN/EQx74go/e
jCXV5RwsviXm+ULP2iwHoc6zFW5lf/bqNlhdgFEFd3D/n/6+fph0thOkAeKXnFyG
qv+8S84wwF1xcb3EX0nUfSVTZWfbCeMoUUHgm7/4cOgWtETav+rF6hMOo9S1ud+k
Lo9gYKXtTDUvrrSMf6ndG1KhTf/6WfS0K68sPTD3wLoh8qjEz7r5bD5ZIfGt61Hf
/hpTAniAzdzAwl4z2x3TQLpLrc5PTW5BmbyabX0c7o0ylchb3RnHyN1wCpK9eIlO
hX4OzPDbYHXbQPMrElJ210HJOfc2wW9mygfPErjbEjOK5SapCtSSdYMGkiO3kHqa
HYJAcB0GJOgwKBAMm3yp7Et5EOkkmRuaCuB5oIQPCwyy5JOZPpa2HXbrx/H+M8vQ
2pGNggotf75Zf5vqqmz1EaxbLOup92QnHXRNGH+Inm80e11bxVyVZ8pg2YAmNZta
nzzqzBFECx2LyArIpeXa642MAByFulr6SIm2jXN8beVXajaMvKVHY8gBWRbaJHAh
uhdjehuFJrv64PIydxGhfl8eLLgJwzowHvIfiex1GHQRC5Mxxw8PwddcbiOKvJ3E
5aKXF3Z8kLMHpMHQbxVlzgyzUDc/w2ZyzafNHfLUj8pzFLsW7Zt8b9YfJkG964MD
Dgwkw1eUXohtOaib8ltlLFlTgIA9NMkC75EdGC688JCuwi2WKcUn9woXsTlf50o8
0pWSzxgGsaUICFM8yczC01MKp7m/VNiTFz2flC1ZFdFd13EgKte0E9M3pEsN7W52
+c5OWVrGsaSztih7vD49fElI0m8yhN72ES4dwG0Ve39DT5x4kKEt54iFpmnJfzpG
LQUmVjoxow/OHQS3sO3v+bJ51JPYbk+qf7G3U0E1UtH9ScbhXIsteCqGLuyuo/Z2
xRx51HqlBxuM9o9jvqcFwLsD/EXtltoPCXFu2r1WD40TcghUx7gcTBMBcdgKFAMF
jUEExGLKEEsJruWfUv+yO48Sms4EVLNlagCKkNft7BcUPZuyPZZ2Hx0trwGUjNWA
q6MerP4jYnLd6fxzZcItuNAoGuggGWNsMJwx4nYh5zFy1WgubmPzCLPOljmgdiTg
RlaEqdpzV/aBYPTiQnvake9dk/Ukey/nePRobHS8Sp22vJuUXvoVvAZDimiwBE1w
lPw/yhUgn9QleIzKX22mw6Os8zbO7fB4V/VP6+ETkg27qBrShjNAVcruOGMKU93X
PEjM3GueAIan8lVPQdCZBFgoO9zkrI8IvFziVrZ9WLGIWpVWvhSg+AJ1z8+FRBxz
aLx68YrCSYYL+RavJ3D0RKh+PDunrKQ+J54msFxNOoj8I36I/8yB1YGykRfotiq6
3MGNehwk3Sbx10oF4hbtc/3FAo+QuljIqosZTwm9t/1hL3oHYtOWxUu3qog8Br28
3Z1PafLK408Cp9BfEM8xC3WEW2c6uwaJ5Zva3gzCPVFR2z5yE1EU6YRIyKb78D0k
q5yWkxVPk5WyMwcdQ8LnW/Wltraqw8tEGpE+gt1P/KmCPRhkf+MzOY5IEZroDd9m
z4L09gbihucA0JGGRYfz6+eKFJ7rB040pFbDOcRXBdNSKrKn8HdVn/fqiyJ+taYe
CAod2p7+txcpZUL79b6sXFTVhdaPMWD/ZcKXAhF8ynXQc2xA7mBpXYxVxID+bSax
ksU8HHafm8fEzNrV5/QP34KnPZZ3IUuswc6S8bw5GoM9dJNG7Y7AbMcKyDeY3JJN
QRPx7cbL76Do0I0rf97iYRRhYW/PMKXtCAiI15MmbGAeUv60iZ+iOeMWBp+ClaL2
7K2MDzj77xUBfxT+Wp9Pk/GuRTgCfBJN7MLGbcExc2Hx2qPuzVZ5nPXJiJZD3Ecv
28tWPOHFiTuGUihnD0dsAGLmKZre6uxvfAw1ohFfUh7wfDZITk/1pUSye7/HOKsD
UxTlsW03/fmRYE33/iMOUaqezWQIvQV32BJlRqidIcH7aQbQ+3+X0gWV8OVy7rEo
iUrVMSqPJ1cbuDWnfvZCgZdRPm9KOVBL+5XPWy802vL2lc44R7lhRkqlkxXfthgC
EceeF5f69fG41Ado324HAFAv53ybRGEyvRDVOSH7/0Llg07Xa04m+YwXZN5vOv+a
sIc4Oln3+UjgHAdlvShoY+yrL0JXb8ZDZY9uYGpoh8DDG8jmr/Cwk0jHR3h3Isvn
q2wXHpXchhJTdFGZX4iIWibV/QYEsY7V2KdkfrRMRA/L6xjqm/xDEdAQmmgzP7kA
OrZ1HVtoicRD1GeFD0FhU25e2j6hvtJ2ONp8VK8bwQ5vegP99eIFBYJ80QXHom7Z
X1K/XpQw6pJ+4HSMwfNUj4QP3ZB2C1bf7qoB34EEu/Ta3fghqJxyo2LSi/2xsIqv
Jd2jaPPAGp4awEpiQCqureKQaJW9gkJ2Sln/+9SnvPGz2VeTeUIBb/1aBgXRStgj
0oVfVRxaIO2YomdXXB/PWqxYsO/cESEnyoHrMvheTrkGcEjd5aj3IqqKqVoRjXgD
oI+x6wpFtLLU9NePfjm2FkIuJU1jF5QmzNvbPM6f1fDE8/MtNhQV8puW7E+vp2rb
PmUrLPKWHxbc0k9brASIifBD25Ygf7s5+LDXvGKklvFPYJU+DW0ehHVNYRWIK/yU
+svaXpRrJ9BwYNorWEf1Bjt5AGj0/Zz7KSF5CFwnW38uPQ53CFop5Z+YUXrktFlf
Iup7GZP4pg04pFBTK6EWp8dRj9ZHBhL5zjzel6VVzlb/3dSJyhJERJPLYgcWfqmk
WY1Ys0zYso07uKXXzIyfFCVULQ2GcPG7lvMWKF5uPkoT3/aTfp8RUr82IDZYyXS7
MQgxs7pJOeJ7A0xEmj29a+LNU5vlN8vub064Z/AK430yGjQA6kAvMwEu9YOwwLy9
+yh4Ayi5NENF9UUV+HNZIWp6XvHoOK5WD1/Za+J5xQSUlDKsza5MIoQx8N9jEHlx
8rs1KKiekoqaP15oKY+RlJNFIoHUOxA+3OPqCYAwx4dA4h0GzLW4aU4FSGIhc1t0
SFGrddCDiLyvEQ67lutAKmvT+eGzy9/YwI0fXiOIrgX72uTWeB2Y4AFTQOtNUPqX
DEgV/CzsUlmiC/V3MyMcz4U6SlBGqxxCly+u+d4NfyYqx3ziivThis17iad1BHn7
ZYZBVbNN+1fWGZnBMFC9Sru9QMUOh3ZNQ7oobBOwELd/a2kL3dePVPjnF3R0YDic
E/8AqBhL2QQXgnynY7QzaXWUfvhPJ9CJe1Y/uzQjRsWrC3RrfSrxX7/IETMvfbKz
9/OH8lR/gef/T1n5M8E9X1ut72dUZhVmJg9al9E5ybOc4jeUCTAlliq1z1hnuqXf
b5l/uwpj07IClBI8HGWiRXgqJsgR1SrV1aT8+DqLdkCrlUPr02MEjlPfN7izIlZJ
H/Mf73ccgqREImX3Io/eSttBw97eze7pD+8HYstOkCW5BnuP6PrOAIHBal9xfCaG
a66ht2ciPY1l/l98O7pZLtxbKjLF30M3bCcAx2xGF7gRghmriDND3PwmS7+eZb/0
XjITUJs4JV20hlZN28KQbod3UJHAy3eTiubtt/UkMt/w7EE8FYy2WyEI24mGlgcI
anDet9CqhmY1NdMUDfsgauYY5kTFan6UaadfOryCOSAKxvrnZHEpAGpL9gaY+JOF
XaxvY36PmEw9k0dyReJ9iIelyUz6GT3BlVCHilN8MGnNnN0fJ/MLb2zk5GSWmPHY
6HdHjUyIhR4SvWRnkJcOaX+e3ueuR87zAZFlzBTBx8h3nrW6woWmErJFWBWaj5kP
DtqTXcFRr3LiNLgsf6nuuxdOspTZ/MohcVaX72g0Z4OlVc8GSwXCfQgCDXBMWgU3
9FWxJcyaAg1hFyo3XDAU1XD4nTSS0SqWvead8sk8GKRV/RF3lLVCJiXi9SeOXxCz
9pb9hU7WnV4Ly614ptOCP1KjUagYkbKF/KFVcaPZ9sA+7M5cqcbKeETrcz4Mcj5R
JEABViksUiQ2mquRpwwaf9QryFlB2IG0kRfPptG1T2GSv5uxHoAiXiV6gx4jhIdO
xKHaJssFQ2wW+jMpRbBa7demD9XC//J+GjOdHzYCzm7S8bYxj1hBr7CdK0sA9wS3
Qpr05R6UaMZmaFoszuY52WQePR6Bc8NifF8Sq3rbMc2wrMIp8sbbFbLejOr/fcmT
xfRICailM/4MJg43m9yQBOkieATymhyLMaTCbGd912pzNuGmFWcQ86wXH3veMxMx
GyuWZ9GUtqKx7Kburcm9VS6Lvcn7yB+kpKtRQJbyp/2gTcDHWJR5O3+VLwJUbYyN
JzPJ3M4ZjUYwZWWlGQQQEhB4yEZxayQPXdDmhLu6eJSBxE87KpQ5WuEzXZGSntnT
vjAWwl6bIly/rLVPzgT9pcnuho9HgEfBbQUEGz40NTNmzpQ+jocGkv8SWAZE5ZoX
c+LBKGPiavCMg686d4DI3uwhEAhZrxwVcBSeD9ltmTmzf2li5JceZjNl8OqncNwO
2EtQnhWdy+g6aXwEixv2FEkmuDenjdf1x8zitPYP/D7YxnJu+bWpm9xQY9X1dW2Y
G0YUCeDA8rbpN7XNqKUsnjpdFGjKorGf0mKZ+8wuXJdyXgzN24TNoSeCPKY2BBsW
PnNldZSnrgA8aPStDTYkfkByH8yR8oZzWRTAn3OrCgAbLwyfHOF0NfeZ+soln5Yj
IjIEETnp2kF4p/T0J2gcOBATiEJMREh3y4QCFOvli0RB3UbkiLw/VSSNpMc4SZd5
lbJTFXuW3iZiBLTX7Ny0upehpj5luZKkyBzD4BDUYZvQeseuE1RlrAbjJmARl2lP
sRFvLXFYUeDXiefRAQBvwo7Oda0LpwIS7kzgRka0WkYYcrkzCfjgk8ArjQrOO6Bs
0TIQLcOIRVW3fWA/M6m8PTWfP5CH8PsH2xoVnOXll1w0i5eB9GkBK7EjhovTf2kx
9emQmVIA/cYTouvpx18wMcBCbM7BHxAZoXyt0rWQMfUP4tm3KKU1SUgBSXR2jKXM
AB4sxcPsf5H8sgoCpDcCSCMfBhmrGWmtZKgcXhv7PIK1ARGTjKzogoT+ZLfYjoeS
FA/wSkwgf9OqH67dUp4QkwQS+RX3RXg0PPGOtI5iZ++hOb+qeyGMCf/SzlbtZ27Z
1IGjA+DXo5ml0Yioon3dIj+VCbxGN3jZakB0qSjm7DzgFMQBmb91pat4blORjQqZ
nVFyqFaGu8wGsKA7DGcnrAZoo8a5OvNB1thE5TAHllPYeoCGYeUWqY5r2zgjbCPp
RiGuD1tPaEGqQPN8qNqpZ0jXPDm3M1vByTesGTClyG1OR/jfE4HTwzmH+CF2Qrlv
l8BcJTo68oW24ZQUoce2cdkc1Il+SFSfA4FM/S3cEvUYO81aA0liMnmvnujw8zPe
Oe9LRsMSecaYzw4m3lb3NKSzhL5AYTi3mUQ6GUt0G0BQflBOAsGB0nJD1ln5Rpj9
I3I2sbne4795PVppxQxJoGsk2gp9uZU6VWN7rq6QddCPN8x85o1TFEum3QlE3j9b
GgtHx06M1CGG5929FQMUtGeQxByb1hShvH6Jv60+E6Op2tss9tHUp6TMCzXgqjpK
3nhxnnvAR9MjnTregtz2iqw1xbnMyQCF3C6HU4FWW7xpFi9lMbx3d046+fTGiqMP
pcNiDvNEbCy67RF/TRwG2mRXdG2H7ThB2AZ1mSARv52ddlfuRH9bb1Vz8D4hhWvN
iwSnSiBdZBn/XD2O4Ya6AuUOxbEwf6ruwBlPH5Zs/t1++NqY3vLgqgXF9JzG5WPv
o5C8cYx+tjDRD1QaNYS4Uk2nVg3CSJhKh8SYORwuqPZAcCY90JhyVE4vyW9v9k4Y
oK9Ck7/7bLx4VlSjoKkAFLdIGOWcsgmwqOFKPmprMSAo6HVwkeUkOXXDiHX0lXrm
Lz2YKb5TXhzk+3etWtdykm+/d8Hrp97NB6a3KWj2V0QVPMu51XXl/L52qIGWunTm
ia0PEpnMT3BPJZx8Zv8aUK0gbOT/Z4FzFfHxvn3KjLlNHHY4HbZVfMPh5rVp/l//
OCiiIv+G7qJpwh+ucmamWVPMGPgAWeU3w9S0LxTVCIpSPvbXiNyo/Ih4QbGxRU7E
Rm8oiOJg7eHyPPp9aM7TyALqoxDX+Ed5nRfu+UBmgYVJWkzjnDuZeD97J7ygoXkf
OOwGhLvWNamY42z9qlB8MTApHaeuJInuORFD0lRiaEgZmtE+5oW29Ep7q24OFlh4
ZVMTsWoT15dPcT/CNdPVRWge+w0kcmyLTny6eV14t2L7ztAil/REwYmCLB17ptcM
CqexwPBGBhhXfYBPq8jforcG9BjYfAMATddm7kSV+EmRPdkjj+XddMQPg3DK3MvP
XpyoyLAPwXJULLmOqKXq1Hfp9l9+jNLv0SbCDETVr6z4+5hnyoAJ4t4k0fpH5lCX
QDtn+3DsUzUYyMQ9va8NhQSP5lmZcoFa0DxVAkrQvsSz2RzoV/lJtdqADZNkqoVy
eHmTH4Fv/sPz0dAdabzcy6XSRCyy/KaGeAq0DwVoY2NVquKGTR3EX+h2wQlR5Mil
2tGHxOTQk56LtM8cT4eLE1eju53IjH9OaJ4fJHc6udt/98sHzyOIaGXZ7I3sQDV2
M6guB6ZHf15yY7ApG0jI/O2zkGzRokFeqwQGMRzVokf+Rgnz5k5padRLZIi/24g3
PiWQWP2SE8fGT8dvts2FksiS6CDklZU7LZTUdSpggyaDAXGMN9vsIFGSPYUykuPT
IEJxxdXaQ351tDVmkxlMuILUukj51nTktpoqt/nf/x5t/X9wRcVntsSeMjOqjJs7
SQwtvF7udUsoRTKVYRnJj6A0VjL6wR4krfA8jmzgJvQWkPT8fCpK2G7N0SEoIpjg
hMNGbhjAR6fed5xNpChIAZkot77r0WAlSNIEAuG6vklMZNMhNR1ndRRwrIcYS4aD
xMKwMS2NGAHgXOlirwGrc6nPOyuqFi90jGGHWvEVhc8C+1/MDeS4XTiWQ1EUdZHE
HJM/FVDuKee4qGC8m3EfPEnUllQwWFZdElZiNqYcF4k1lYUyyTymGjfF5mOYlUcb
lTehJ3t+7XGY8xhNBiPIdeXl1ymgENU3186+E5au9nBUMYvXGujvwBEmLehgO6CO
cGyKT8XlPAgrSqgT7rb0nr/hpCi0KQ8LIA18jn7zNdGV1PGXHvTMCuFXcyCKhi+3
2GWEYzX0FSoS6ARslNkrWzuXVeKu4eQl5ju7O1UBfIy3CnXc6IX4yn9Oa55xtGmL
hMv6rrOXGCAiRfOelHFjVXY2CCHCBa6rB1dOzXTtUHMIHMdJVRu4XSunP8VuyDxd
uuHudvzUBm+349voFqGbL2BUM7vP8Mg1R+8M0w77RfWz/B26DrUnmQLukQBUqDl3
/MOXKqOR3kGxomA7oZk3751XCh+FLnqzyBCm/eExsf1umxSEqQFyr19PXUjMb7OA
Ta0x/orLVNfv0cmPL17TwOB+zAym6BoLZU/s9WQm8qXeuoCLE8Dft9zKvQgIDnxd
/pnelzM1m3pQeK+JR4mSkp+2rZzE0iwNvw+GsZKXM4sfRe41qo/2kX4vlNP7XsvH
SCXqBl9EgaynvGrhG5mvuLNEEDC1I0z4RE3lS4xricMNN5p2hWqWNrNV4JvkSsjg
SDWThrcSJZ1EseIwX42izpAJo61VJ9OrMULupX0VtcC6xbZg+JkxCsbymNXWD/fR
iSDQHlfSqsTmo4oMDVUC9g1JCX5KCVOj3V5xVYgPY37ACKO6dfLB04lyfFqGHexz
QU6ylLRNkqsloQa3+kYfyZV086ffYcbrI5OjgTtpn4KpZaseRUUJwD5GLuUk8+Vz
avPkvJptde1ypzVV++PSDAf71iqBWb0bEvRWWwvXqQzWzDmHhzM/AvDOu2oTyIlz
XZS62SlCmY7d7DRimXQE3UkFhorpXMP65cdF7N3bePhc71ESMGcHd28NwBOaF6NZ
QL20VplNb/Ta6BWcp4r0xmjYN8rUEzRIFWtL+hojui1r0NGQ9RM8e68sDKHryrgE
7BwE64wGvALCS+VMz8IdnjMNO1yxLEh7xjc4x+yC+0ADzge8qRHV/Y9pQJfe1Z4V
Mapnv4ggOUbCUpvNLwE/lvj0FbYDWvgiuNjyoKq1rhGXNREDPuU5PqK5m3KXnKTA
mimR05aiuTNGe9q7P2tVh0KS+EIst+izfLVGEbjwMVd8vvQo7vDR8hhlflt1wTJw
wqK3rzWKXQ/Fo1ZZsyO/YKYypP0aRNMJBDdW2uiuKtGQF3ny6Qm4F4Xm1Xe+hE23
U3fI7Mf5+nOZCUxIqWdpVCrzHm2JS9OXaEHc7Iuz8GAIo8MdaQMH88PreYeEo4mR
eImI8k9mhGuiqZkGOJ7qNn8JwwKIO3R3zy2u26kbww952M/BVai4aPu/rlIi1BB7
4MhgH7KsvTH9vQoEem2k3l1vMgR/qfwK612SCtU2bCVUQf6FslkfbD9YfrZBjjgH
mvWU0HsEFDXLPUDYxzk/k6u+jxfLZN3+wYXVBOBder1ofwTHt1V8Etf1Bqn9vgGA
gcya2oQ5GGtYdpCdVdbTb34C6CS3FRpO+v9pCs6yls4w58+gINYhJmKzWWhtoH0A
+l8hrL2mxmL6pI67fvdV8xbexvNZZnZwNmJ7VXccgBGgKId/MsmUa3w5KvtixFYf
8fk0Ofbg16nsJrYrDbDHoYDkiobSz4tohra8e7E2CK4Suf/Zu433H5dDuGkfhzGf
WCvGogRAqWfPgEkEA8QOhS6aIb5XiChh4m87kZEAaAwrQbcW+509vfjIMEF2H6HU
flmSQUBm+qhzhZPjddIURqwUvr7IYTuypfJciS8mAyqERQ5CyoV4BRY2lBLYsOJ1
7uL0IpnFEpTUJH8Xb0MWNkYN74XAHd+x1hioHM39N0B/oqQKXLlBDKhIajQIZ/U0
So2zyNyHgXd+sqrOVQHiYXph5oJ521gmWOjPKKkcW2G7ZBYX5ZCvxCB0thZslK4B
/18GXRvPMy49zZGAuUFFGxPs+jquArIF6TRlPajUR8Hswr2bFygPdoQ4qHp9AYsn
la4SSI3ONm49ebnUyVfZUvSg/Ju+xytNhje/0UkpzozonxARlC4D1JCcqlGtdPgI
eJUjECeizt6/ET9U7Z4CBlviNcbAekChby8RS5Y/uPjADohgQg7BcDOwph6aIIBb
i0UUt2S9NtI056uj78tVfjb/dHvnn+DO9wlk7XyntMniznvINrsM1FouMsDwd5VG
VKYWACYOx/OhB8T8ngeQW9KqcZHc+DaciEMX3wzsDgpa9i9l8AGWAfVZFUGM+yz/
N2vyK7yslaPd9s0+hSbWOwJqrfVtZh6ku+zVgNLlOVm2B2lheekmLINcybfnxoHN
aP+yZhdZBjSRS0N6hZmxG6+sUUoFZWvO+t70CLAnd3WyEBDB7tlVoT3MFnWeaNC2
ThDOYbrI7R90K1TR8lJpYySPuZDDyUZQC27Wnoa00eYtZmWONLR11tbfOwyODxY+
W1k7bN63gjGzXxleo/aY2pjVR6T/RexPhPt1Nu0R7MHpfAj/fXp4vUv+oKxCGJU3
XseWp4SZXbOYn/orSGUWIr5ygsNXR/8gOwmPu4NyyoxdUlugAEyMJ97BHbu3WGN0
QHaUjzSVPMRZa+WqUQ07kqUIPsjvgasG5VKs1gslvula/ZCj9eT2LNnEe06yDwSV
eIWetGMaoy07czA2afJ9bdO/8ul1A0Uc/YsZW/SgOkMvrHY8FjpIbam0Rw5gQOzE
/qBhAK6JiFNwLqSn32fAt2Q/YOiNjRGhXRYB2+iok/Dew7yGeeL86MNfrN/p5wRw
NOnv52EnSRvl5U5e8MeYafMi6npjHuqCJFedODubCeVYY4hk0o01sjnsrdhh0ekg
sew9MRIPBo5FmZWnTiFiQW+XpasoCBW6ysm9EUw3dFI7TqowiokZYLt5NQNFHmd+
QlYntqX1ZFkcZpkXQTSV+oeFCG55am07ov3u4RPnRjzTkfGGBiiCWzOvL0F6W9aT
UvK6xppV5HIpnLF0popadaJsdZXsY7taYqDinoPFhcnO9BlOlC7P7m6QraEMN0CN
qwCh0Js+W7/2HN8/Ae+hQCjguivZe0sZobNpV+9AX9sDWOnG6vMRBV+VFR/n5z32
7nV6ustQpksyjMUJ0DdVQDxp3ZkwVLrxhhDTF7jmYICdqIiIwPSPNOVz70z8zbQw
OM7yp+bkyIXx2brDoIfAG/4btei1xceoNrRYBIk7xYf0whp+WNcMZq2n8iM9uXdd
U2knu2fsyVa2Edzu3nYTAdZVdvZDCd1koH7NgaDJywqqRuLd8vZGGzxG1hBSOoto
sv4jx8GoAwCkWtiCpg3cyYEP3wWvYD8jhqc6k0aBm8/4noQFCKpuchMFttngkmyi
NqgB8Yu8E+5/4thjrYXiTPJCDcsDJQszZaifYgvXQO2n5LmQBj8F378dh527olxK
GLnwwPZ76by1nRCJubvf8U1uuxeokqtnOsc2PC9369a6/ocrb7F2nTunFgifggRF
wcwM/qphb8mCM7Z4eMQKt9CwG7Vq8ibMB36UetB9+0g5ZBG6AJNaZMTrwG9NxzYC
E1+LpYDTd61rGxRId+tk8uO8lNTj1SKKRY8E3YV8blZsT7GB5TicE/ln+BmEarma
hGdgWBmXrsXxNofKpTo05IinojJ1m3O3qzeLPZWfxj3ZuEXAwXPrzqRB6fcgxow1
k7jiKAj5JS2vi5/P61D5wA1ZuEE+GDRzDCvPcCWFIHLcuttlFffeCydwLmzJhvrC
BUldg23+WTnbehw5d2APqxlBRfNHtNds2f19TTuofRDiVmpM6zVKGxSCIcriN+kD
FVzLTQszNGHk/mV863aD8z5Ak96Pje1rxKr7JowlxBIWvM6MSSIq9gPZq5FgU6gP
nW5I/FQOxCDZoeP7O2NbjHeHe8h/XWZXSUV6WxiQmqLnqFyfi6Z2k5KLbENpi3Tb
4XRSdzpZuZ2Bn6n1GO348o+AorAZ7yjwrsYoXVX/kG2D0A5gRrlUI6NubU0tdY/F
SR/89bHbsx0heq3RoL3KfjR7ubJ/rW3uyeY0YEkOggINqw8BTseEMF9P2XdHUs52
eAvMjGxSzfFZYA7g5xijnPz+bWYv/LJDnsk3SEq0BkkBJ+FjdAIB0m99rmFcrWGu
hZyy7hSxCQdT+AaP2ajReaJdYQijBMpMYfX6HYcO2yIshB+dY0CoPiFujF4AibTh
Y5rAMUSgdbHy+skT9YkVmjUSTi3LVQRLaqcT1vEGGrXTRHraxfOHrMgvNyu0mwtr
EDmJpD1vOOTE5ts/k1dCsbqUarfhU6sxl25Q067rCXKUEinpO2YZF+q8T8keiZ3o
Sjh+qDl3cBra9EXHuo1z1yoyqFcNzO14XaozuCcnJWY5hsOEaBRSI8yvnOlIFos0
UV9gHJ8JH4vn2T1sdFO0L+QuHNXTql3VRYCnpuElNnxoBEEaEtU4bK4creiH3SVy
tBYxJE/SW4HLnzS6c4eAJA2CJGEwXCbV32yG+H649O6FjFjdMootPMgzhu1VH7vn
Om5VTnhhcBaHmufNNW9p4mriVZUy/cqrnmVDjB77ueqvpVt2h2djAUKbF3qs0LJu
EIiNEDSz0PZpmL2A3L/n7+koHCPwUFnxNhw8YZNN1ASBtgXq5eN0n0kYaiJbv/B/
EzMf9mOrl5wqz5y67d8PjtyI7pkgA4ycAPxngnPe6xeray0sWIp9IOzCspV76ZFD
e4dhuPtsg7zYzvkHnZy0XuFhm8dsaN92OZlb1pM3Cx8tm+XBn2H1yik0TQ7O167T
6haWTInLnrtoZ+5/rn8y4hJQwY5CZ1wM82YSI2vnDvTLYGfghx0Q6s/WvxZpyQDK
jkL02SRIHBjkyLEA//qDr9YNstVa1wiQEQi2UhP/RXthOKQoAU2tYjOtRvFCMV20
xsPKgA2XpFO+aOfy0nGY2zYsAtQrO7Oncu8mA8WQt+Tx2KlyXMEMvz0y9YDR5Svx
DutAEkGkKQDxQYHcZwDYKeOZykBUVWwJfpvkK2cmvqHlFjF4qymu5LwYmygZ2eRJ
+GSVLSANx51XJmm185tuM6HMijGha8bUHaMPTqFpD3C98vmqZBtjYKCSeqhSHzbA
xVDJP6TRIUQg2611sPevmfElq6g1H4NzM9xgenBsZZirZQSvRJ/Iz6WQUqYy+d7d
jnoY1zARludA2hmkH9WCilT/p30kfAQaUIh5qpIK7B1gvP5Nzb0/fdmg445P5TCf
yWNtakR6L3Xjs8B/ACfThl+sMi2ztQwkVrFxYjYCQlph7stclJvWEqhAlNceGUK2
pLdIGRkWH8RjmDf+Wph1UWlTijvhK9DRU+B0ft5dA/wt+SOF/4I3Xtu6L3s51D4R
bcpOCzuPxMZ2TIB+Agbx5vUEe0RQnosSkIrg2u+Sr4CODMWhQIH1mEvmy++0Sryn
sKO9mgcXHEwy/TOiIwozKgCMZ2WWNtHjvW55CaorxhQ1We8nYuBdP223emDjgA1G
yZDsq9xdSUinYDLRBrLM5ScbtxeZNlF24dhksfKxFlL77uwRW6qeNFT3uxvGUKRp
TEN4YCpcSdErm98q0Sr1hVm7FXgCaRky9o2JpAQsWvpMXulACJA5nz2IxH/QI/QH
Hwfyvf2YyhNPGvsVZyR+r/Hbxoh959a2+j7aOmirsHGeOAI4X/TlnfQvWhdbqdtU
ObibYVmuInhbseFKb6FrzTSZjjzQtbysh3OkAIHVh98BaIkxiQbsOTwhJFW8Qdud
MbZ1hpg/xvziYdp9MGmpxCd/rQQnWcWpbfILjea92ZPIEiGn+IMjsybZvONbYEhJ
KN3y5wi8C/mqpUMxnQlzYLXnArqsHCV1vW5AElotpYWKSg8/vlTkUv20ODuQjhef
XJPg0VLsd0i5i9r9mba7l+5bhK88AqLRFr3mQY36I1mGXeu8L049SVxGbbz5OEkX
+ddOevyZtjM6aTknoh2d6odfnnTBznPROpRj45+TGjwfth4vpC94KJbSV3imuUHU
DuSFlJS4Wj/ds+Y2nwPN4m0TkKw3nT4wv127rI+4il8WSoJDOW5q78UbcKddMLvb
GzXvkFIjcbzWaX1RcT7hcl04aahcTX98BR4IDO1MNdK31zXCMns/6p5DSbAIJfSK
0zjZULw5ZTESvd586CXvC9UecxWWAOZ2n+RFTNFpO2P/sbzjU5IarCpuGO3lq5O+
AWirN7bs9Qog6lVdsmVi0HS2TOyB685/rSv4c30lWSAmL2u1MBrprzW4oLl+khki
qL2dlWZ61nxUazAAqQnCZKOwSkHDfljYqF1fc/4EwVqdyFUu5Cm3eNFyCpArZAPR
CL0qOQvGXXSuu++mSVrjf/y2+q2REdLvGTlYS1XYwyN00PoAflAoCQF1um4V05GM
JZnCEsaYioYGtJMGN7kT0OSEfGXl8s0NsSqhr/0jBMX3LqC8bBx7SKEKeN/NF/A9
l0jKb+Afx3OwLQSGfbODRYLZ3+VXYM9RsTdLUJspmRvJ5EvbdKpcLavuWHUtiIYh
3c4vtjXPt1c+E4RBTjECeXTt9kjcmehPC4rAyqGrBuUOxmCDkvlKsgL/aUWKLFkP
MmlVDvEhIFXof+0cAST++7fJqsVzXY/+TJMHPmooYYDvyZkcnseGFpgLYqnm4RA0
bO62elIsfj4e+DEMIVXGJlajmpAYauMiTWBFu9T/2rWz+9K57Q8V4Y1ElfjN2glX
2qpehkONe5nH68DUKUIve3XOrndDSt09b2ac2SSCCGEdwLctHa4Ri3vkqRG1siRV
DwrR8ggc/+FZaz82RH1caI8+o1mwGK5nJMaW6xPBCa+hVHafXVYKApjNVG2b9LRx
tPVJsfMRHf0hkh4GAoQTMQflxK6gXBjGxqy3bCATZ72+Z3RwV4BZ5bDaVAdN8CMk
8eefvpmMO5XyHe6P0WdHVahiB/9Tq6uXQFnoKuTOkByiH54nqDcDks09TRM/tRQ9
DRFQ6ILDLNInzMX/2AND9fVBNKva2bWgC+ipKpiE++IDGf1AtWXBiu7tRJcSRuEo
4DJu64w5g5+mPmQH5qtzqd1Gt7zue2KMhPP9FsmjbtzEjAwdPu9lfBfUXepdervm
FZYRr79Y2xl+K8HriEerzZtULYZSYmrl93s5ec2FOQcOknOekbOHOnPjZ7Cp2cG6
gt1SbRzfu75JH9OGE7sW86y6cPOgqsTd0ufTKdQA/AMrAj1ELAi9emrW4jn0as1B
UbqD0AyE0MFB2Y/MaIqhCSV0iLqqIgGHZY2Qji6nvgctawmQ9deDgPFjNMyGmFAW
xFNA+WjCbTqCZVsunNQbMHCrn692Tc4guy3dI2AZKpcH1Rf6nXT9d0U22cU1YAH3
y3JN5VYhIgU2HI2i92o3KmOUD+GQPg1gCTfhD/d2Z/6RG9cNeq+manpu9OzSFkgt
r53PCPFZIb531Sg0+2x1F0GM8PVCM0Oaulb9bWRbKzUa57ezg7krOUhc7ZMR/ew4
NAIC7N4ZiwEWLwHfx9ruZDHSynH5tIp4YqevCInUVZZ7SjjDSJrdwLhvoe+GNDE4
NHfCjeQj5B0IMRGFX2OBHaAi3Dz5FG6JLqSSZDuZ0JxjtYJDFGWi6CCBu/KFWkGp
xQ7UA/Ld5dN6GVJ343qHYciqK23H2KNdBYDwuEQAzHZo8cN51nrB9WVW+zrdyf7n
PrpTYmSCBnVtTYxtp2c2VYXJKPdtpOtCKiSTMEDFBZuElVsfT9fNzILdc4cV0UHD
kFCCG0bvr0qt9geMglB3Po9aAlfnxCw7bEzdYM6vFBl790tby3QCPT6ESN3BjzzF
2csFgvFi3KlNd52T0Wve0qM8B5pJzgTZH1JRfBNCH2szz6xTkak/oKh6iGYSr7Uh
MIywarBx3i8RMDkyhGezetOZWsiBujNU0gWbuoFvYNK4PyCKKJNncBB+l3PxAo/b
nF/rFzT94h9bdYmUSFB55vjG7YHWu5yemqdVnrF/bS9dr6Pj14d0EAJsHen4xFe0
FyvxTmmed0rVTl63HjWTPiS1OggFhwy447GOwP/JfpcbB5blK55EpOByUYrHK1oC
Wc+Vr33yfOE/APOdgJC7AWZaO10LfZdOFxfn5dFE97vqVaGGpUnbaERG7gkKCP8n
dJSRfz6atqrlOPVg3CpIdyd7kzL13fSLqmNqnttc3z/37HOpAxdKfnnsA1FfWByE
PzsJEkJH9QBbwDMhtMTW0sAYUkRRWXyTQQEcJxlWZNpqehrsoRQvaQ9juuzo6elM
yzmovM77lJeFCKsECracXpj+gtzyJW8ZYpnd4cKt9Dw+4ZlFQX7IAbyRGpvNN1gv
yaKbDM0ORtZwwP3uvj5oRu5xU/pvDgpkvSjRONXWcbugiXva9GxjcbKnT91oqVFT
K05CZQr3T5xFj6EXSDApWHz59A6DjmQ1MIATxOPUnKZ7fR8CQIqWY5k7CDeQiX8Z
WcXnL0jBHhBwK6EFW28gipL+jZuKcv6+KJj7MFdYPkV1XUhGm0ktCupwSzkheFLK
l3nmi1HvyyaLiHZcOJmhcyuJ/6mTj4IHDcmmD7xyVv37saKyc+MI+/WZRGSm6DB1
vNnE1CekzsJcEUD2rldWveToHc4Z06+vGedjoMxGxbYsBoL/FijdfXcLElky+u3T
z/Rs7x2avDYgmI6dqdTbNWK7xetoy8CiThXiSdD2qX8ZOhynnR1jPilhoIm/huK5
7T43FJkj6a9Gv/AsOJFP79tyGN49QS1c5vZh82ZvuE5CuS7sgsrLpIozn98bs3Mm
B9EUGH098iohMtPAfQEPW05BNv+2UhERRCE89FCuJpmcQmeKWOxnm+6VG+4ywB50
bEkRbETzfb3T6EdGUaR7jlGniXnjQ/u3UZGe6Ox2LGZyYi+65CuDcIjR1pdv2nUU
1uwMsE6sB8RNrlYqfXmBPH2YfJJ7JeO5DnqSMhoDIWL9KRmPLLvwgw/T5qV1ZnQk
sljq8TaBANyTi+toceSFMm/1kUTRnDTn7wous2sOS+QzLViLEAMNqZPMKvpJZ3xH
ZsEDUNIDqU4ocKAeKjdNGoDto249UznDjmh7sgpPZwUhYnPFuFU5+5ER0HHcRncE
jNdMyuGIHhaTYefobDAgE1hfeUwJBH1bbVJtT/NHIA+5y6pnyHT1eoxnPMu8jIeD
KX1jBzCI6CGjF7Q+rSFEZSez0LTxDgEsm0pkrPFyBkZSK4DjcZnM9WiHRs7DmBeT
UMJ5jYu+yj7omPJzYW4m+1j0pP6jTxl104k/I7QO3nRNbby+9mIX1M+HJj1yFAfe
sm57E88ti5evYFSIjVaMheq8fKG+UlxKZuA210bANG74nabcVD8rw03YevExxQB1
MbwUBlnGMTyBoaZKRm/AQA0FG6bwVktHuagsOTM43KzHmA9KTstGqbXZX7C66OLp
A53zoFwnNOF4kYnX4UAFfBKl2A7fsYBP69dYighzzgg+20vy4GoxWNHAZMffGQkQ
mxhl5RocaqetfYETmwQ+fXT/PF/RRvuKRG7lE8a5dpNmQYurFYGbwQsTqnV5facl
Osy3TdX1w4Bp0v4+PP5REPKGGbmkRYF1xRRw8r5/6oIiMZHcM1/PZI+7Svz5/yUL
wfgzXnjVnEz3PwG/GEvrBKRTAc2csFs9k8lBaUaSJFt6XgB6ZfV/NVNnNurU4xIJ
eeQUu+EV74Hnen3nXvEOcTrTBAfJTRbfC/PoyDm0+AaC1ukNwAAFCgcp4sfYv2V9
lGy2nOMat/28oXyWusLjfAIbolgLf6rw4iGH/YfN9lYclhGFeOnP1NOWM1StayX2
kcTj0ad8fuCGd/YmtGdbyNaqSiLolCRCtuu3A8byXKVVseOUx9/JQPn/hK7y3Hex
jyv2PnjZ7wjwJZE0HB1DTeedbDsWYQ7wlDflIbrJxF64Zb2qQ5eJAR5vp+8Uhxjd
ZKjiF4alw3oGpQwM7y/OTBmvL4Jte7P3iSpcBjbG2RXtDKS6VTjNzX8CVzSlLO9H
qe46noJjUj89rY+0BPJdbFiZVNKhoHoeYG2xhyssRvIv6HZJbZ5iMiLGN4kjq08o
U43WA6yDUEIlzfNzO0eczvkmn+mKAxlTUTmLrQSvNpahB5HVr4j38i+evRR7MYA/
b0D5SWh6XPUBNCZk3I2JR/7MxNUni7YNv2nbNw7R7Dk6ziV175CugJ3MZZk5JzoF
XpmgG6AbCITIVDR6TTrBRDTI88jiK0RxLav8ogDaOlooZhLUXC7mON9aMEKyR+z2
NvUz/de2LKElewelJy1riaxYe0uvWLAZ/BiQC28QsJsLBXRdGi7zWckrBjNFYk6Y
S/qmDNkcjpD7t82eYYwDS8DeNMr5Vb8RPo3z+ZViozq/ApnDI37l+yVxt2zjs1U0
YbAlXpu4EAVlMax+9rYnR0K2C8RSgfQ4MwZZjAOsLY8Ta8Hzav+vEVCNokpFQ12p
k4Nb92mln3TegzZKyIxSZOs0eV7Q0J0RUfwY+TFuNIUr5eQ76kM9CKTZSP/E59Ph
HWY/DrxQ1Jzgp4iZeo5kpRZ0gg9c5TN3yar7Ff7m005SEHArnT0a/lUlTCDxTBsc
MgwMdZhEkfABzHiw5O0E/ePp0MDQQHjuqxjGBGzc4kTDAS4gglL2tFsonbdB1X79
jBh9x40uT/aqnlyxtPIMgEmtUarn4klW4xTcu2Y3UUBwgUNhIZa8H3OCkwJtggJA
sHjE7tsSVmc/kt/wbTei7CIn+4j1P4H+mahl0q5Ha3gcctTROzV4htdIZfqGKW6r
B+YBolyzJ404U9mbB0MvO+nMPQUG7QWbSELzHgebyusnvAeVHY/CoLj63C36vlCl
mYNxi0NNm4wrAs+7yR502JQeSKYYAKl+TyiLGd00fEXmVOptGiroExBPrwgZaZhY
SxH4Cr8rq0DDWYqbEy5AZIxe0KwWhsAbd0gjrvByMzXeLdn0KonWK0ADzbkOB0l7
UHavsxEY5eMmvXgRc7Der5ZEdgiRKrBOaHswJgrdt1KHpd3pClA+TpZ/01emT/gm
OJ+ZktORMtQDpCnsjJG5l7X4+HjtFPYiFGLCzu+dtveZPqILcYU8kiJVKzDMffuc
k1tnliUET10GFbBHnqwg7twSKL6Lbl7kJFVhg8np1mWOgD4pmpoGlUiyNEYu9GpN
FpR5EeFJhhgAVZ0G6zyFKaxZLruN+IbvnXgqo6XOV/Jy2+OWGS4HT/aNg0L3Di14
DlBjGNJAacvz4+1NWX/YBNKa7J7pw1BQ9/jaYbL2vo9kYDXO6O0fJ8oKduvamtL2
djx5tGxQG5Z1Q1qWhNU4vqUB0j7ukKso6KS8WMI9BYLTlYSjP0XSBt96M3b3ueWX
03FpyTuyjcQTVrdWTc/T45tBbwG8T38gREMvx1xP74fCgnelObbeWoeQWgGCuZgR
ZEtPmtnZCsqBpQgC6bsozTZDt3F99xxJg8IebblUct3DxIH7MKMRBRGFBJZCnBzU
LEkCQ8X7EoeXhZfU4W7ohASSalItYlg7PhW9s0r5x7VtCbloo1lCnSsa00Mp2Ttt
X5/NDqB4TEYQuNR8Elq6Yt8grmC+h2HNgRAhwbme6pzCzNHL/Xg6NFl0MqFkMtku
bNl3eWLOnPAnDyantMWvBcP/WYEo/mCx1fFwJLP5xYaWkrcFRYpz8FXE+VhASvOV
fFuE5kcI4J+BvJrkA8/akZ4gugpt4wHkA9YbZ45aze0Fpgw1NsGHLutqvQT+soyQ
HCFd1787X44xNFXQD5tPW6IsGsbOUq4SsWqHMrTUgCNRa9n+QZhA66kfFLcUBFUr
M76/fI8LTA9QGAaEnREuctyBEn9JUl1Cs+FHNSc67gx0yIOo55RiC36yZXouqOms
6ALe/V/rcsGW1EjZrDEYr18xt/sU6GcMOCfj/g7ZbZJZ+BlfbVs3WLyMB5gd0JhJ
bO72NI0S+Sg6CZc5ZTKXRkvO97+fXlmFzO/G1ciEWn+g1zw60ref1CcDUlgwHvRO
z/o7HoG0glZ2qRKAfE4BXbt9zbZw4k+sINgS/h06+6DxFj8PjXSvsUxF3umym1ml
Yg6zQ3y5oURYb6WMqZeTmvVhPZdjhF76cLlr8SDLj63sV6o7pezMFw6hUjMUWNq8
AqMmxiTGJ1jWGolc5QNS5aI5ZwZSI2l7TlTgqSxmgqzfveTL/bltKeGGv1R0sGj8
uT4C2FaGCSGDZTfdi1VlgZFu4Go6/XuKRwrDY6j4y9cxtVd0sL/fHr3vp/lu22up
7ueTPgJX6elif0hqKlP0aFyGkzw67wGavI7yp+QMtR+YAMEl9jqucCRiVQM+3TnI
A5yNNdiDIUNeG3gMbGRIkv5/Fa2CH3H6Vtsj3WxCp9uQlHzpxqca9uwUx3daQx3T
9e4Xqc+5aWndhxLdIKi2trIAEeheC7NSX6z6i3cw2xbO8CduI5auh5VxmjcNU9d/
aDj9Pjlldi0oZAjkrj5AaZ3Isy0wYKErCPubNExd6n8/XBKmnceiwYMPaojL1iKI
px5ymtJB5Q1QPmrJVPU8ysSqNc+jibm7pCDLmu/s5FiICa8Bx+TIB+tkMcqaT48U
C8X39wF3acrUMOcR6a2w3yFHaXD5UooVUyxVctXVdAW/SBAj/MSwUD8XUDlkoS6C
8ufNh2kZtLkaZ49KN3ojupNBxLlBBGcT6aaFgZvUUB4oX/SgTrLtXYPaFDjt9G8u
vldF6fo1xFotZljF7e1yV5PnS1FYBO0LNI7Zto39EfoyeFvnFgmN6TCoTLGof+O6
zcGOrgDL68MjpcbOYyK1AGB6xxqWt3mQwGcvb2tBVX8sUEz55GDfVnNZAuAKknCq
8+AszW8MJMToKh8WwMvU0he69EobZFzpJitArJj0CelfQwV2epWrJBrw5Qsnv2c+
nxlwt8u/yB7uYW6ulvTJYyo89y1aqMJ5go4e0ouU2/CPo8+s2k8OOH36NvEv2Tyx
tTLwAUyK0ZSVCmL8HCbBa2WmmuwFDnQC4b+MuMC0XY9EWLhyMzgUGMQAgZicRat3
ZjHboG9CXh2ZQS+JsejG9kvNiuB5bqdynGp0CKu9fWjpdQRNvsCmbYE+QHN8ypVH
aNsuI2exAIxl641UnYUy6tildwVJiuRCKQzyOFgRh0xy2X4w/wtfECmZxytnUPo9
XxaXKmKBzQO6OUVafBCm+DtsScK/x0ijmiO6C6mTAYZvDWOf0kFkIN0336cU2cxP
prBdhWmqit1OdZNs4NGR8ajsnA7nE+zRBpmc2/u1L56w3yRnoAj1GNvC+fwA59GI
AmI1h/XZMNHgRIiVJrVSDjxt2tUWY6UIzsa7iZd0FRq3wtRY4prnlGttkE1qCEJe
nRzxbAN0KdgDKCCv1iFUZ96bbMkG/IFOME2PugnOzUdReZYkZfV/2R36P3GOR6X8
EKGGJb+w+2QwUOkpgZC620HWB3OJi+y6PhV6MnaatPqrV/zDtmi1xF3dsniqjpDW
c64E3kns0o5WblnHrMFgvD85cPQk7YqHYs76B5flCSlEic6ByzMjWLIR/lbpi4qD
nf2Ip4LQrmt1P07EqvKHBRmUAq6WjFPvvG7xAS9OSvpXIAd0pN80bEopfB7EoUca
qig88IzqcOOFthp1G9YUjsX9KJJTnpoW1m59doPUxoqMtTrDOQ6ZJuV9tN5Yn7eT
1irF3p7V6TSRBacBLAnH2I2CSPfZg6qFwMeRrdml/l7Bb6T1SfateldFgRuSeHhY
yty6KVTxeyVUOB0SHnM2rLbzoEpkkRMoOoMn0eWZYJJib0QCaFvLghlYJZAfjQKH
hJnbS4tyfEgMmyUNIZy0DNKyGGp2NKBI220nxlUPvRgoG8hcQHjDH3KMyGqkAOUf
E6ORCp82g+Mtt9Z1vcP7/4DEF5liQzyC7pkpb3jLdC3lE5JIVKIEknepe1rsXQ3S
TUItRBy7oYhe6NOVsKgUVfSC+qUh/PYivqs2zIQECAPARUtqnQP9pmBTnpPtEu/P
5UgHKt3ApQFKnouMBJzlnSALyy0Do8qvn+zrRSF62wLlI+YJ9ndXYPqWApY3DOt2
mN65L928mGLjUqReLe3dkkGxn5sWcp22FSCKw84YB+FzIdCu8tPxFmF/0tZpblbl
4M/8EGdUB17+3PVSbuGNRfTPBpSK7+GHOdProY8tI23ufmEZohU6gQUnfan7+FNb
clTcR/EWlQ1h2ykPRuO2FWyGF79/xC68lKbhoshx4A/DC6hSen5d8zTqr6Rvnfgd
/su1lCdi7nlldBsNy7sv8RmP3kxUMlPPNKWt0SGNdz7m725ymhj3tkC5v0eKAAl1
WaQvbOT6ZQH55TEm+lQ8nHmX72BOT8B7Exe6e0t5w71O9h9Pcj4H46Igg/bXi+aD
fj0N1j4uLtsxyJe9qBPsWrbJesTlpQGU+vkVA9PQa8GANvbDkTgBjkisCJ/f70t2
vBlCRkraS3PBxf6JBAN87Rg31L+1DLmzyqCUvoVgNfLvoFPTK0j7aXM6ihF/q6EG
0hau+QLn2lIBVW3AhiZFy/eErn2e6wMVxAnWBdG9HqoA2lkh8+RJmPnr1WEwl5LL
rsGZAFgqiV1D27ZdyMlJDhnjbzHcqJLTCoD+BIaQYroKe+GONolqU40HotdH5XLD
k3kFZ63FPaN3Bj7RN/O5veWV2tSvDFsP4Af+uW1Y1nu3bQuLWTHGZ9LaTKnRHIb5
C0fWzOfBkcdkratNZUREiAa6NuBcI9XTNkB0nVcBXWy3nffIj96JVrdkVehvltPa
+jOJL71H1733Hr9GUdkgGDp3LJhFxowu+KHPc6/VmIy8iitAmenKQ8xxQ0wIIphz
yDWXFIQDsYIBurLKjPnERwovtSaoTZzW+fnNVTC3Oo/CX273qI6CGp2FnQDVWEyy
JLLaA0a8/S5wblYCCkqvAFeeUHAzwTE7B9n1UoZUHLGdZxL8kIfaZiA7W5TyHOiy
3AceBfdeP2Q9SAu6x/+1TW0UKcMzp0ga6lcoblj93UrpGc6xXRyxRw4J96z9mUfF
WC+xtAZz/GqAz9IGRV+5wQp3G+NPNDMWHrZcy2W0kIVTPFJANexK0eMIeJ8Zeklt
h4hD/ZQ/oPXeg9hUp84ATSp0hmbm/YqrA2VtU17RrrCPDWZbqV9HWfttEIpPsOv3
Icl+1JqTtHQkSTR/I7saAEmvGPjyoZfCAEabP/JiNu37W8eLcDiftHKMSGRc+esy
RIloTGhM+GGOYzxaekms/emoKXbB4b6BQjLhycB+u8tafHFy5P/bsNQVZC2/isSK
w9L2ob/Rit90900ybuK6RxO7o8KSC99JH8duG5TKjoexFp4+rAT3makH0p+I+cQ0
2ugKnIzdJOEndjRNulrzhxkdp7NiD7M4kYTXtdXyqo4lmjBhMfJ0AwMUvOytUrWL
fVKibq5vHeA5qz2+Ybe/6T17akKpvF8f19Uyb7FKencgtN1w9iFbWRc/mu0/lLGx
tqfgnmtDLMds6knSWV4ca6JNAAogsr0hbMdcfvORSv2XRROieOsgjmrD8LxaRsMu
7dgVAI9Y4UAWeL+BW6kd5lu6zuVWYOcVlx9EeiTJeIZoRm+cDzOcmQ+xMt98Ygfl
SfH0q5yJZbtpJ1FSo/8rzMjVGQ9nb+IqJwSxYFQv1Nb7w6ciHrvrO/FdylhhEa6n
1VQSmgpolbznBx0EuPeWDsAgEFSo6aUnEYwD3RKSX3LVT6S9N3E5tFvshbh1fCr5
fVKqEqALa/vbS8JM90JptkI2ZLcU3V3AwoCwLgiIRFseVWFeIx04ZZtC7nuVKnYn
hrg8t0AlMM8h3OTcYeGZY+mggJlnmm643Z+/LXfU9vyrQndlvV5wWl+Uc2mudobJ
vbBiIe9+rQ9NzJi9RSXtu2Vf7UbofvSglucaok9GDT4f0FkWgrLHXTBenKeXjMge
T9cnU4utBTYsu/baJ1Z0kK+Glh/VCkRpAYWYLMA90K4rgHwzFU8sxnQtCDEHrz5E
tn91wOQ27rbAjKLZ7gTyRfTNJIorK9LlcREe1J0SRvSKd+ybr0jfd/xkevna5VuY
ySmZPlYa0KlGofJVPnmZl/YPS3bLw34lNWqlHbsvWrla8mLMDARvF/462bW+ZK4k
muM7dHcZEeyk+lJzOQpicIjYFAJSwE0HbwNekkLBx1ky3sHD8vLZdW9smzMSel+M
NA/8Qzgzy4uK/hIxRKdv6AjVFF5z3mWonlE1Ml6IlXcQoypJiolMxOuSsasrHLjg
1viNtMJAOOiQ4VGEYZwvYb/fZh7/mEtu0mCp0Y6ZOqNZ9opstGqTJ9SlFQZUW3Pt
VlB3QGu9TpELwIfAgCHSECmy6TKFIPi9H4hOkjHZiIvZGTl/SWsIXUbUzvIj5sFT
p4+oosF8vH1JBokAIULqtyaNl1kwxajBS6o9sIy9XGz4WHYLZmdER+D6nwjyASR/
2laRPQWBJmsyaxvM9WCLHJtJ0V+k6+LTgAZilpV5UgpSKVacpmqWbiCc1Ux36FPM
0mhHT/W6Ja76h3UX4eqs4ooKSP10FaTZMinioBcUov7elz5c/nLwOF6NcPl3csSA
0wsbN24LgoapewZcCGEG8tK81R8k42CaUlmN/iv+bqeoO6jTAowKc1ZvlKstfa+J
ehSTlCCutBHRw07UMRp4CWxX4EIUUg2C6TBkrr3S+HSv0zhEFlX811b74mB5xbDo
DcPVSPENf80ZpmKLcu8DTSTuGOsrB8Q2lwrGxhTBiMQanK087vyao2Nlcsz7R+zl
yS60WsAp7ytPbgfbPN4gezowYFoZ/62Ujel0ozB3NxMxQWD+NwwXQf9AS5ePW0uE
Ia4bVz6AAiglotZN9TkSx54Ir7Cp+e9wiBj1HO4APv18BicI9nAHVfYQs/8j2uLy
fI6mJLVJi+nP/7Ls++S0ClWOIajhSio84jRZrd+jKXom6g7tDPdQ5pFC9mdKI9Fq
lodk5Cj6n2jGwvESmdCJHmif9UZj/NwOnYNdJt1toMRUCyYs3TFjPpOZHLVJHkUm
0KdIBq2VoyEyJunLHW+nj8WpeGg0kiLhLkyIF+wdkTA4OCYUAbp7+ZYeu4+tWqPS
kHwF9nKEGXhMTfdd1kJFYHNuE2QgzcbC4ODVTLZApeGkWtQ+DPjZ6Qi+on8skssR
aTLLY7o6oQVkmX+0roX9bLpn/ZdEHy7SGMxRZWoVGzAkDpG5pfAvF6kEuxY5gt6C
Lh2JzaPj6xxpJ6iOa5080d2QDJVdRuevkVTkr3UkuJlMBNQ4wk+K/FoKIX650HEU
pHT6tOk8gM7WtlL9AechwTSv8ANmSbSm2uTLkG14OEUBaIWGZ68xsf1C4qYcG9ZX
NnTDG5svy6PeoTGiZQakU38OaP+3MIvm/QOnkcErS3662iSilAiQkanL6Yhu6Yn6
pWZQLjbpSPsSK3ase9WNEjnLC8I0CIT+6WOTVZWqKpINaHR3AqX/jGldzS769QLI
xE2YBSg6eYh/tZxzgPUeNTtUkt6KtVv51g3JcaXx31/GEYdXExh8WQWqpwbBL1ds
SmMlSHT1U99ntN4eObMOLjw5SMBS8fTRFSzwEWIMv2T2MP16XHXVYa8TSuljoiSZ
x0HGHSNP9ESjFnZdam6+1zp5CcdasDdYyS2h1o5wmzwtt/lIBZhlDqPtpMeuf9M4
ugEtsxNLA9aSWtinZnUzXM5w/lV8PmL6wH4N0oQnGH5usdG9qZIfuZ2SRDGrYhOY
H5NH8b8q6RBGJun2pKraIGLQ24qyoaHXoC9LVrKatbxKHiD6TSRVONzlfU98EYk+
cmjBiJ5d6+hWepdHkWBUNHE+0nDHdS5MX8lwWReG/8E356omZ/ocoMo7vkQvuTLi
jBW6E2VwxFMw4h/fS6xO6xgmQkb2GwlpQYrO1k88CbXTxsMOkNfY0g01F8Z4fV8K
Qq4MsnSvhrRt7cGaKsJ3+DdCfH1vs4ndDrDDY8teympmpNblvYlMPHcXS+3YzU/U
e56ozKS8L7HsOiTBWIwmOwnsKP9ds8csCyZCkuwliIb1O/SZgdocbaqZZdRUcUQd
0a5OUhal7LoR0+UyoOYuoRFwrLn1diyNz4x9BS971gnRtJ8Eir1jD4qwQcC6//NP
tOCnHMsoB8Th+Df/yU8pZ/GS1BkD6V4R5g2sOs2HlXEVNDDD6VkBtOvs610d+fiK
SjCLTKusG6X5T1PNdcXyDA7cxvRzubAJ3TvkfyP1bpaw/DU/tYIs+v3nRZXYFKEs
n3a7H7D4F/SM5y39gC6UyHtQ7wB4r5RfkX50I7/DecvkJrQ5E6xrs+2+GID0IisR
WbCrvv1oJ8wRUiDwzfaEIJ3q8gQ/ESu7mNV9Nn+klaYyqWF4fkzUU23TPrCDp2ab
dFdqIM2jtQWkLb5P66ZRufKgTvy6SmMILF3MfE8yL/n7F5yK4u7pOIlkDy4jPGBJ
f3o1Dxr7wmbyx+ZgmUeBJJxRsuX5BxTmjYLeBO7n3iMfcKkYO90rKZTyXd+mMc78
YkZ0R9epBJad0Y3pmmu+aITCHi6hmW6KN4jG5fifcwl8DzpXsUvB6MK2iLTQ03PG
H3uuaE0nJlhdeV2z3Q3Yr7QVPK9kyJrjoWITFKyykc5B40PSQ9L7fOdsraEZI5ZZ
ZP1j12fQeQKUGXhmvjd7vU28fIphW2nEjmfKKJZsFpr+PV4CvNp1wB2gt5d7Rrsf
dWa1O1Eg8i6yj2u4wRK1iGZtPw4uua7baNSdmiFguZ7g5QtIj3uy3r8y+gAROWr/
Qoyui8f0pxGIvPICy2iP+GsNUzEnzVnKxahekZG0bM4tcRvGwPD2dga0Xi5w6AyO
iE5PGGOorb5TCPAnDy7DLLyEq4Zq4Sd4eyCs9E5d1+BETI3AXZnBp8nvXnKdPNg7
Cyu+plOR+8C/4GeC6rHdDIe6+d0wWqyR12hCi8oYXO8tQdRcEhV2bltZeeTk3b60
+y76WS9avf03JhDZXW/TKM6UdRY8BhGS+m+GK5ijCrLeKOlQkdloXpnm2FJ6fDNR
7xEjCBEn18oE3X4Us9L1FFrRl3YFTj+Vn0+qqqawoZHN5JN7uDRjMflrvfIVJ/P4
HVFo9k8zp86Pso8P6n6qAHr5HTOrqtv+3j+zLBRepDfdbj9YMkK0qPDnkjnqvm62
+hoUCmDPwxGZ7cPwSYUg+OTRJWKRli6PtzmJMSWe93Uh2GIbpc8fJkmBujkBvrfV
cXq5xIam269LyWXPEPySPEi0de+9IbUwfT2ceuOSbretu9tirooyMGEqYJiZvVAS
pY0w2qc0Pomb4vLonoxWB0VB22XU8/y3KNMdtQfTiwrklf/+JC8HBcSBNZx56CKo
3/p4Gnn+g8cB/EXpg750drYtNklP6mOJcoKPQnxnDiqmi3TpXzT8xQqbkQ/VQpp+
nltPeKthaGbr+1/YMVkI33rLYe5u2xDFNrz61EiJN+lbMHQV/N5GkUG19bSL+0WQ
X58aKDY/lk4h6QWpOWKSSoRSl7Lqp3q1Ti6k2DFVqURV0522YAujE7sXYrfXfz8G
E8+msHPzH0f1do/p9IJjHAecTlWzqEBZNNncWrmH/Jmd0PtLCGqwefeF3kGtpCB8
ANOpfduwVtMGdvKGWHemG0RAt0fp1ewiidfWwTDO62zxDGAuyQOiKarSLWjn8cgj
TBlkhhNFcTIIlhyp4OCzbWfkimjCzGDKPsEHD9lzxH4BAT5fHwdoIgSqnHL4Jtx6
xh3Gd6tgBRROYi1QMj+F4murY6iWroNHbZ5XrQaJB2lCR4OLCOCUeycr0iEy8mHh
b27HT8rzGapIB75AqSrfs5IybC0Ojd+PKCOfuQEUQ190MccM6u9HwjunmO70FGof
R9v+HlxCpzOD2S0Ra5gaMMxu0iqpqRJqHdESMEAjROPH+0I5LRknBM73a92GzzTq
IfW9YyhAcrXduZ1o/FNqap8py8OWUR+O6+HCsm5+0KTVL5oMBCaxKsR/mbuwvCBK
DUaW7B0cPeBK1apwrlZlOh3Pw2zDoxdvsYoh+Z4qj9za207dt3qLfCC9qbQ+uC3z
hQhTHtqg3589/6yj2aeRK+vpANgYl0htmTREUQgHeQ5KqvwQ5MHQoVWTkp05YUhV
I4Tu8ktdnSmU6EQ/oA61ApCakpBPSeqiFpWQsEKWTTk0G0JRR8Nl1408vq7oXMtT
lj7zc37GvMhu2ylzbV/ZAKr/GN/qfKq43d+Z61uGou2fic0izXNlXf8T0PLfS5BV
JKaFwG0S+MKH6r9jKPTdG/Tzv5lJcBb1hg3Ok9by1VlAu2EuPaPpRBJxMWGrWwqi
g7ap4pX6ArAlR+f5y9e+u7sF+jSvCJROqBx9dzOneT2sWmuFmLbtiwu0tdMlpNpb
oir52LvICClB9CH04dqXJX5NSX1166Y01S3KdPWbm/IB9pQDAjE/A+0sqD37aDNQ
2c1IhwJmeqDLZ8j089aRAgf4T6eBSzVDu4rZ6ipveICZz9SvQ4jIQ0HwlfGpiUU0
MVqUwBeQYjjj9f77WRt7YRziIzaTLUVTlqIDRtXU6207a1+yFzezil7hSIZbnff1
9bF13KH/YphmAvq76FO1HYTUCkHcb+nJxC4o9aOEQ8Kqf+R247EHjbRPaRRt7mvL
B7GxiMWvfIzY2Mhx7lZxXXw6HtRcwPViH1Y6G382sht2xa05pvcawP8bMoVqq117
vQRnZshZKhKQCEdXu5aCoZ9lTr/VY8SNhph71o24BBYxnm9RKVJYWlmkWPtiS8YJ
+ecH4wlXCVBqPSNWrUs6JvVKGF7yM0A1V72bmRfQ3M1ps8TOzxM21woHKPE9/Pfz
x6uaHBb1hlSW0/GXxB1rU6WM2h/CFygChoFscSJ11hmWx3hkzELSkGjJM8nlGAbG
p0yrlkbP1IoS7+l+bnMYzmsUVNkI2ZW4URDG/um4id6Ma+d5q8T7yShQvMFquVkY
Z5x5RHeG+9lVKYrVEnkd7VkCJj+9W7KaHjFB6Iwl71iJJLyne8QGj52zYUa1Vuwh
VAJJ/sX8DFNtPqQn/jX/wCSaJf0vk0ugIv7hphvtW0G7OA2NkChk3I5smWHnJReM
fdA3EzPjF+BuKFKUzFnW8+bS7nU1Hdqf75Cfa21rJ9HyKawvOjlzDDVDuzsWE9PH
UiIyJTRgvUwwSnQcU28/Uj+1glWkiZUWUnFFbA8aGtnIV1W20TdrlP6FWJ6Ns/id
Bseqa5H0ABU52/Mho2BxRv6WqCCqV026b9fObGLJZNEIqXhtUqA3gsJmi//lffUt
judVtjXNToWX3yiZAF62exwYHQZiwDuooBFSyKAfkGq8AkkWAeAu7PoBiQdonzb/
XIDSGtaqtaLGWPI9xjgLNM+0dn+0G2Wc5yUgTSiLpWIsIgrcV4jvUMbH3hXjwe/H
gHk7vCsZ9awLJiIE/b3v8BsnsMtbnLCDUIP/Z81+/SD+xVnvUidhfs9Zjz5qdsU8
I5hVmZ4Xi1RWxBUUD5CJVs5Wb7yGwrILd2Cr0QAkOZvNXfPB2LJfPVK6WBSSQcZU
kjgg/Sp/uoLVJ7DsytVDe+TvfNSZrIENEAIT50h1tOZ/zkCvvyYdgS1FntOvzVRp
Y/vp0wuV1ziXNnVHEyY8HAXDG/h9QWcbXLI34MYoDN0Buwf17pxVf5XrP1BJtglV
kchwq0kOr9vFBROcPdSPFVuoaFWdgzkWVfPM0tcKHrI8BGaBa+ZrZ3NUrSLmtAes
T+MVuI/URPkm3aPXHO9cp3E0XX/CrXBe+w9rdSIumKB2gcxWN8PCe2S70S4G3OUu
AbACCHCpYiKYMZovTPCPcs8T2TtgT7NKC2HxUAp0yhp83PnM9b+BqgjGYujy9s1W
uP2LzcKOexQYiEAQ4Zn8iCBEcXnGtneWycu3eUn6fX//JNcBe4poAEPbaeDogm/4
0+Xl1WCATJiMOvDe9qMH1QKxM+pYeUxqC1LeDrWTSRGj5n/LOJUC6EQlydGdsz0U
f0/DIDwVpJj4CCCSEZfnHWaBOjEV4FxiFp9ROaUk9JshOqmPrziJvsuO5+djvc20
cnh6cux8b9nqwVqhW0IEbVBsEzdVdqgrpAjeV4BYfPJxBlDjxgWXnMWMdSTR7WZt
/aVAoLztpiLTjpmXuJTuda7M1Gm+ENyEjWLao2c6fh98arTnKEnw/HSSUAvAJ6lQ
8koUMl9Qv2lIz6QdwCbzoKSBBnoF1Itl/hDmZ7Rxxg2xLIDFen8s28SQzriC0ei9
HDZT1o+UwIjV3D/nahWi3Vh76XiZa4t8+pbZrbSD2eqjgreMgv5VdDscPRPOKQ5O
Kv05ogPUU+piJ4Ngx6Fk/Vpi9lONObLTzdl28ju6V63BZqD2oNLqjtZKhyYtCWFz
0h28Lgp3SQybGYsSvUrSyBHwVD47DC4dqIsTshSqpVqkL/73exUhyjumpOht2tN8
ttqgk+CjV4b4Md7uIa+aYVJziYXbUetaOr6Mm+vIqIXdWeQIWR636Z4rG6P7iPdM
mJWFydy5QxqqNT6xzZhjDsRehUWHg463TAMNKptP7DScmf0rZ6HUUIsAXo+7U/SC
LNT/uPBgQwVF39CVJlt6/soBp52I+HQsTFna8vAE72iPx2IsWAdTL35Lk7yyevnV
7zGuJytG5n0I5yN77mKpuv4T43VofMhHYCaSZEQVdP0Ay1SyFSe8T/+ZXI/0oJFo
wdTgPAKhkxYOe7yPjWjZjXcBwtxyw4B5ri4IjaotuiWlajitgtbDAjQuqX4hhetd
S/n27HT4sk5QUKoBhNsihA1qKVbqiCs6jY9Ib9vf9GGGu5mCcYSxHs5LdHpNMB5M
tIIuCYBkrWXW5K+WHuNvO53uPCgmSmZ8vLgwaFYltBa74Fq4ibQ9XvqVo1eyjw6x
KWvOLp2c1FxB9j0NaqXgjhm4/P2Ma9poW65eO58TmfPm2HIW81Pe9dd9X6mVLqbO
y0jPl72Xw8Xy5abIGZZ9vHR03OkfRtgPnTdlv9ise4iFoqs58j75EUuvY3Sm70ec
JC/BB73NxPsAFg1BYupYmKhJYlIh0sWEEVQRdlzfA4tI7fIfAsQoN0f5vB0Uxhny
a1TDYUI6268/0TvVkS3QtkcDRiolUEQ8YO3zvMXJ0MdzYxCj+lYF9Qw5Zq6AR8Qc
mYsf5uJw2LvyealOp2/1Q1Qyp9ktjMt5VvyytFhPCXrocbd36HMguAzz8Lrs3Cg/
oaS/AMX/981DbFCD9YpLwdiAaOVPjXItLo7K3mGSt4K8K+y/siQ5RIqOZhso7B5A
XlaHMn0wnpyY26rNGDAS6HF83ADEYyLOxlUlkorOyD9BUb3vW8O+oCpspD2lZoJ5
rVO6DDxtp4gYA2CIbYjaiGj1NghOFW5mQPIwiJi6NS8ooBbLMO63uxQf49Lc4m4j
YrP2iiPnSN2KJ7vpCM+dlXrxMEhMbd8KdjogmOJrZD+3akgdhtwX3MdZ4ZWizM3+
6MIm+AQRB4yq90CQYqAQsGsMkrHUVxWzDSk1MUSZkafphFjbzo/o21KnUPEKc0dL
X4JpLo5bFvzl9a6Mqx8M6q3/41xMJVO45QLpqEL8f2TPR27aFOI5oNtex9doLYHa
4Cybs6MFe1cdTEFLqFY8F1b2/YPkfdDECTgnozK2Z92rVcfdfQMxoCOZ+izjJQo7
HFVSV6qNEm8VUd/O7IAIowZlIYsk/G5pjSWDkvl7jiOnT3hngFLrDhgN0Vmeg0wt
IzRPMfjxoUGCOxeuqexEJTThPdqb9pediLq2jA+D/r4m9tr2E4IlrYr3372i4UgH
skyiOUdF/qGnWkMiC+BM+nqQBa4I4E2O7zKTqBwcZ9IRHKJ8ojEDzdooyPsM6ORB
M3grtrfjp2LRK5HgozaOGAUoEYh3qpcwK/hBYDn13GLssZTxJcSADn0phn3DlvSO
IAB1lxDGxsT/TK13GtFnsCYhV1OfYMNcf57dUB4JrNsvCHg0qjYrQBSvQDkdgP2o
daGo/1pAX9xkec8vlucNhewduyTU2qATFs/PrxAJAzLKtuPCyE7Rm9E1KzTVZoau
iQ9A+N4dFwZFYCERqJFDCjBIH95d9xTO2Q2N23Zj2Bnd4JLbsfKcm7GrnWXHTSxS
9XMxrQHzBBusFEPLz4lbrBdNC0OK7ZnuPji8QW1D4Ug4WYfGn/sK+G3Pk1AETvhB
NprPjRGShQYYe9Y7J2FjvbqVFsAtS8xwCJxkiAHegZf4GqPZ06h9fpqVWhQfR73H
ZLSpxO77y5d81cRsvzpxBLoly8y+SRu1ZoTzWnsnnTLDuOEJlOjC4rWjRQlOYDI3
41djEJAqHGWYEFmqr2PLiyI2KuNMVL464kSAd5joo3E4LHyEAGTXUGlKGhYCHF2E
KDt+Dn2hyYmUQVRW+/XUTRPqAmqaCJTFiYFdrxDVNvi5kopTnqbLQWD99rIPBQf2
be2s7AQGlBlF5oxwZD6pkat64ayDtQ2TO1onpoKU8UhsNDg5MYf8eRgcDyPdM04g
M/Sc+YaTHz2CU5ihS7u8TUsDQnWeK4WzpsAE64Vwr77YKJf5YYuUHOTWuGqOcrqu
RA6BeBXk9XQxUvIyuur6f8iBvh+clYFI9PwLUsUYxus6L7Wy0YoiKhfLpCxRWAeI
UKeh+GU2wIXSyR+1F6Wb8FA0qtGAYwMbhitclK2HY4N5mnNFbYouvE+z+9z7EJBa
uUPnsUst4nS3IyqqUc4qLbtXouZTHntaNYa3qMvr9ubDAIarC8xZJSyF1WXyB8SU
kNXhTTRJaVG/V980Z6DR1j7brDDVcWejY7m8L3yhpBBWRQvZauJ/IqNGD3qaMjtl
E8ij8HQ58zEdVQz5m+SEwpUpuEr8ozBoQc25h9leDRrXZzO0NcehnbFEZN8NUKD0
vvAAmyXLnbFDOJgOZ4IChZZoo2kHqLb5SEW7fkQC+49yS/LFTnohHPKKmxLIuxIJ
J2Bq3v/ltyOeHASFRcF9/dXPk7Y5mdoUPdRXLUj0orErONma8vBkWV/LixNItFwu
16AeC6Jk9sw8WN8bDGHM4+Phjunjg/QFluEe9fphFN8hfvaGAmbeh5kjwPluaf/q
PhlyM9qy13oN0a/Fw38+keisdRYN/DDh9+EFQfveCc7eKUWCCCbhklO0pxKH1FWG
pz8XeVHiDH9gm6x2wyj+zlNisPtO55ogLADB7/u6e2eSL5s/3PX3wqD9b78ep5kk
epBki00u/a1hOCN9CfSoBeJ3ZRQg5/NZYNOWqywi4uwL2lAo+mhA5AFAsDNUr3wa
djN+INSaSRQCvC1JW7zI6xs5jmI4QFk7qzKufgEOSuyclNr/wPCArNODmW0TBvjh
1ZMXys067YQ++nHG0cy3IKxkCwyKJB3UIAT4mN+rCbVIo99hPUx78OnfgdWmGIOG
jV24tA1j1Obov8tkS3tHGAGcVpEbhPDpRhqz2mLcEyFfxsXqYfnSLCgD0boVPHIk
e/CkFhG/R4EWKxNqMrrBWpiIlYkSG08ZKEX7jELZHsOAI1w3uc7lCmGAZdUAvij7
094WbntC2gyjOhU5oiCgWT03CxSV9rt6vvNB8DIIpVUnsBREx4zA+QHHCDmjw/kD
LzMAn7+O9cmKOi6IHEn4+uZNkdX52GTO/IemauYwPGC4xHEVBmC1wyONwj0TfsxY
UxXlfUOKD6Mr4EWwD6A403RhMGHKn3k7K6B3w2d9p7k6BfGw/Xx12lMJbNK+jL13
lTQDi456ZtxqSzwt22WfiSw1uvjabIU7o8WnxuBTJyMpyLL5QiVCb9WmTUtjlTTu
RXDLIS1NQbQloGpzhdxf/kwZr48DwibdHEZui037pTj0iSTnl5Dz482OtK9qg5Nv
exIVyf6cYbRJmLIbh9Dss6F1uAGkkwtRS8pupYLGNP90DNlts9Ehk6jpzqNBN85m
XnMYj8MCXv+UcjQqYpENwuTsGXpEjcdo/xBhgKAJEjvAYJZ/6rAMQVOWRgZP1l/7
iiqu8HT2Oslsm8jbKxhO/214ilx9lJ5YtyEKF3Y4dc3eafBbHa1+Ab2eJdBIb33X
lijikFEeX+xlNiS/iu5PvTLdHbtyeXU79kEiFps2ILELU0H/xfAeEIXWGeDc9a1q
epYtbJfyIN9TRnHebS0/JihlS5Mu8HjOnwrzkKoLh9rQuhPMVITpRcS4vQMMnfIj
B+ROByw9SFBKhbGDpc/Po3zhLjIHvGwZFstgXyoY7fdF3bQf8S+pz5QF8HKoS/bb
DnBa44YRL4t+0TM3rvflOl954vNPxXF0kmKwWXPGZjk=
--pragma protect end_data_block
--pragma protect digest_block
eTaA0zNfCnRLL3OY/o2H1lE9sNo=
--pragma protect end_digest_block
--pragma protect end_protected
