-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
6YsI/YmapRsxBHS3i0zAFfgYcCR/Zut+XXAfGaIEcqUi6Qxk9yTsJ19V6oNimBBG
aQ3Jjbb9nFmsO6D8SoX5Qx9hIIN8Yk2lAus8KZjYKpL4aiam3/i7gXqD/HQ8s7gE
vPj33kJTloqSGUN9uySPaNj0BaT1VRuP7n0HDHNgaTB9n8js4oQmsQ==
--pragma protect end_key_block
--pragma protect digest_block
EcBm6JCNGDtgVmlCYQZ9DBQ1quI=
--pragma protect end_digest_block
--pragma protect data_block
4lPDc+jtWP3Qu0Hn7NRI4VeQIAMcPNypgNSKX5S0LlZKdKoBa30JMVOaMkPXxGUP
bWZGldZlLikhE6S2QBKmXmwDcAfIVHV9lw/+X0XvoQRJAzr8ESlp7BT7COjs+pUp
yezgqGohboAsihY2x/VTe17sYbotn9OToP3pKzO6E+WgmWLpKC5nPSG/NdlrN0GH
NiDIlv8JzSKKuNoTAsN188JieC0KoauTbq02fkLFDURiOlwtv1C7UsaA60vAZRNR
SULp2S9azUnbqJiElcZG2v49ZPorHXpmvjod9rj7WjkQ5NEw7i3XSpu9DJ7EhN1Y
+khFmDqy0kxLPSObALy7fFTIRI5WprraJUv7oesoaJ68tCa8l1eCXbFfGE2xzbGS
2TPI/KY8O7kt2khrZSebW+Yt2Mbq3diI7qJm1WTFW6pAA428Z1r7ZvacLMaj+2pq
R76Ym6HzGk6FaLFHjnzj4tO9qjyTQ8AJdEgXz+BQKYcjWlgjsJgbWvCOwBcYYC6d
Rput5FMLujxv4Wakxw11K9LD7dPl8cLcGiGww5wpLArznBMUuNxtOZduIShuuBlx
wo8H5qMsdY6e1MQq/D8YktAif3qdW/iJFXpv7B5RCePx2iVHHEYw5+8bkuOPvTuY
lUqR+McLZNTNpvnZCNu1J49fWr6wAECZkiugyodn2WuAs1E/30iEGG6EwkHSEqRJ
V81J1sQp/hFhtV4iM3iSEqRS9tCc5bZjNfJ4W3tCuUnYCic80e6PBc487IDlsOhU
Tk9STeuHMYAVpdyH6/ol/l0fY6/MYImjAQXgNFfj+QUe6GuVQ7mG+U+Bon0EMjqU
yQa7ChFo3KmcKbXqXm2ZFtiNhX4RyGUQhuZw2AssUKHkCLQYOpYxHQtLyeiGuebX
ZpEeV/fyY6nqEz1RwE6OdkzbSZ3PdsWRVlwAWvdtkMvjdp+X4grF/Yf8cRY9lfPp
7kduxHZVuchwd6je3tbqw9awqPkKoT4aiqqpILHBsgPwvPKTL6DWyk9cErPHlJEa
OcK79c+HmWYFylu9GeY4OfkhEnf1x4ahRoIwX8b0TR/XVPYCCIUuPDebaw4vjRCh
Ga1CyZ5prool6QDDj3RH1Fs/H/qfblMpVMPSfAcfyfMWESQ53wBU+vOg63O53xAn
bRMKgUbVIyVgPzuK8sZuiWULl2PKFDOj6FbDf2Hes5xv1Y+RCPf/ylRqxktJCGGK
xthZavlmyDwcfu9EXnnA+eZBHtPlq73WmFbNaG1a6mxlAqAynGOtvXp+VvkbG3vP
5dHFJtuzffXwfozAczIrpJo6+b777GR58eJjPn+ON9CHqFbQLOjiALX54wv5HM5u
Zz0GnfonGzEa+oIWkYiobjr56uAEO5gGyR7hgjYJIFOxOtbIdgXeSmjFKsUGDAs6
HzB5jR5OWseIymrtlYZgz8vx5q/kd6u4XPCSUPzK6f1HEVmFjyEU9rbebBpO16Kx
MOYsVYl2Rhx+BAH1M3selmcWTGDfEuUE4Rl1/eyi93iie2QLmjBV6CJ5Ar64OVKP
6x4Cy7247CX6iy+Y024Lq3iyb6chdDhmHK6n3psIVIpTByr9Cv3eToB47/hNstbz
LSuQPEVz3mfsdqP6dj7evItCExtC2o2f/EozWDk5m4EPIhSoqhmVOC5FPNZOrX0B
TF8rWYpzXkzKTApF6HTTHW4l7fOF7mhB2jmQ8GdNM7BTK4/nS4mJ2HmNL/T4Bahq
Fi/x53v+HQyJAhK66hgB7W5zMOoJlCHV/NzzpgFnEMrpD9udMmPFk1J1JEkjQeeV
7E0beqDwzMDsR5/PnGoA/pwG5nZXBUg53ETfYIYigAuQEE82VQyMGoU0qHV+WYqI
sgpriZ13K4H27UoRotawYhl162JIiaG8n8W6VqfHygLywWbGhdQXth6kHQQK0ypn
dwggDvBhIpQkWEXy3USxi8Pp37QnQJ4RVWLYsBu/TKztz6CGMV8MLdCSIEMQ3z50
3l+XsqsmIFnqvJ6XZNahT7TeCq2LsoebJVFivItDTDg1lLoHWmgBR2KXvDodyltA
qrMw5em4FNtWLHOk+WmHZFvhwIpNU7M+4l+I++zHIGAg5Lj/qsuEmXudCowqbYW/
Y4f3ecy1J0Etu7w1ZrJehdLbqekqunCO3QMn4WBZJ+aoDOSr+2LGulv8Hd30Om0Y
EGxmmEvZ6+qvkHN2+DhTi8jEfTlhl7wZ2VUoB/3X2sYdkUHWHx7CguamkUHQnw9b
R52ypbXimi5YvQ/HrnclTz0ch37EuCjnzEZCdtd+IiCTL+yuVqWM6FTTAmcNGkrU
fwGy44CCYr4jakdiB1BfIjPmDbJorLAQfpLbh6p7/uxUlrukNEuSuRyfTrez/H+W
W5AknYZpUKOGpnRSBoU6R6HK0fNIZa8KwCbikV1Y9hwlp6N4XPrqGzckXoY5zn67
b3alZ1xFR+Dx9VxvLm0XzkmwnrVK7dV6hxIrJYnSGQ21dbJ5LRTbrzdDL7/o2YIM
H0n9K91tLaUoms9mdajW5yhBIVHBASoUi/BrPxWUTymSYElM1sC7y3bVg3i1WO5E
hqRAM29Qo3TL1zj4btE7qHLZpD8NoD5PZXVW6DfRLk9KVSRK66rLsHn+6/xOq8B8
M44esNXFi3D/pS57ZzQ/olE12wMTa9Ue2gku06IIDD8h4cXlo7ziCRUoDsKxK+Qr
G+00F+USsTwxxIk8QJzJagNMxnZHWTQsZD32kh+GWv69uXVhwoMeYFjaT9rN1nIK
q1DXGcmugdEgTj0k7++fSoJZN1IDWiTn2yV99BsPavf2cQDE8iOjAQWEVyyHV6uY
vr/UgJOZ/AEVbCI6lE1HyUv6CxSB4nNwUcmaybXkQYCxVkmICUj1V6lYU56X1mhz
CqdLC9Li4XH0s3FCpAJ8WeJgvnE9YcT1h+xvZxsFR9Ao2CZnK1IkIrEtjtOzIPCL
Bl33MA2TkHo5Pb2qo2jhNFIvj6Dv5kHsa2FUhuWmuaowHH4BQWpE3I6It2Ok8O29
o3gfSpr103V9grLE04fahEoaHrqdcNUdv737IQI0Lw5AAt55Pw9R1faYIG796nIq
0r6ts854UmZQDu1qsqwHDAHSsO6H44I/q8nVUermEewNT9aUCwWZ/T45ccPZp0Iy
iYCH88bloMtAm3Zovr9dAn4j6w1ffhFujwmO+BVtKGUVf6RPUF4UROc+xiACb4Oj
iEPguI7SZeDPEWYbg+QuW/M6SMyW7mdWshO9Om2I6Co7BL5LYrYIYRfve+7YMfCD
UjSJ1ATSg1ajeSKFZ9j4ESfyH/h7O+rUSvVFUvPqDuSLmPIk8/mRmIxpB8cvaoyN
Z4CfhxDiWgTnx6ipMR9LPrBi4sBk/ZmIjssgmEsECj9GKDcmNTJ+HECHuxtiaD5Z
J63bfXAFcUndkjrSij0Czk/r+qEg1FsOavlCHD/3oHD7l9/wPBu3WjzvMeRbfnTY
upJX7F6xlnlBwHkvmLkZIB/MYG8kmFMyFuDkTj7cH3bQRcos5eE3lHBAQViSA8Sz
izn+w6EtFjlXf/DeKsmbmRiZZdOy73eF434W3RjO+bPF0rG+TPtuWYHYqm6c2lPb
a6ox1Wazz/yKHCLz7CmG5QGvH0g/WNO+0hle9qXgyP4d9QMHXcOsBevkFVlXDOeA
X1uAnj6Ubz7fJaU4IPpOjexISGHqovr7ypMCk2/yAapElNBipqdl8yTvQ/n4lhdL
CbrK3T3uj8dxGLuXWrrvlALP9eV01wlQEtHsPJHgVCwPyg9KqVgMrNOkODBDBrW4
oLymXodP2fe5dqarZX+OhbPw9SUab4YLIEnctIjbOV8t5OmoWRiZM+kbAb/ZyGNP
lwYI3Eqe/UQpUqCsE5ltxyMhmDxc5CHDC4qAVZl25MZ92lp25PrqfVzn/NJMGgpb
/O+zBL7izKcvFVwGkmG0AicXC1XXyh597NyYLDFBlpaU0r9LGJR5ZCPQc4EzutMc
q7zSRP7MfBSUdHANa+OT8RzIhUpgcj+ltkfh5TMAxUB7GFz4nzn54S5maaRtaSA7
XmFy2VgfosHBqSsIvSU/ioRoYVwjzbC83okx3wW1owMawBLgN/zYFW8Ty7Y0M4i0
Wh/nKGRPo2dGK887bsZH88NE8MHb126gqPrz++apSvYnFtFSyBI57sNys0i2eXsb
2sOAuYCSCo6ZGnUCtw3DFfN/qKIDXMxA3ii8CRYE1OfUFXBI604vqZdxQKA0TbB8
2pKdccBQlSVUOl2JquQuqGO8kTjN4YdiosIZeL6oHhhtpxj4RH/RrBb8JsxLBZfC
3pjdLnVAfYBlEylmvAdV2V5DQ8FxPKAYSoApmHLhGah3Ah5LBC3oD59lvsMtajxV
eUhpwdzXxsyIbUDQdmLyUYqqkSK+mJIpJXcr91scuf5dzF6aLnXXppW0K4Y1iBQk
uppv1Zfvo+ob69n1342q3GpsTeHOzFxtkoZHNr1X7jerWEYOB0ChSrV68dVLamaW
U+nbyyd5+EJE3tDe5Efa1Ujb46yL2p4UWaZrbXPub02Q6HZ1s0ocZo22NkLtwxh5
AnnHKYniNfqhbvLFDPF2h8ISV3ciOwBbOBSzqcsct4ICp8T8OUTmEAY01waGHbmn
FQVbeGy9is+1F9kAy3cRWWFS9WPvfkETVJgxWuJ1DlHfZdEuFyadiM1OWIhNT3rX
low00nmoazOu1+b1pxJVj/GDa11hcZVabHWNeXeRQrRBOEp04mgX6HwBg9gihCoc
GgWzPhDQcQ1NABrP1yRthoVoJPHe5NokZLUXcAfo/XuzxSGPpsaLQJ0QLMMvKjN+
35kbVnOYCQqsF6n5fec6rnKP1OOdbt1/C6DQmyTcc9ZkIg6gpHaG10doZXw15kwu
x9tKFr+GRlLUFPedj9WdxHwBJSzjKrml5BQGeFJqawD7liZtXeRilvngQ7FlVoT2
HnrwJJ/AZf+DTpmgIgmxMq0S8ZBm67DzWgY9726z4fbw3uUqSMxm/GlJhkOcv6Dc
Z98eEjV/AqUBXyblxS0QrQs/+yKVfSMrzlYCGv+PvOoL5KrWABNvzMAFvdSToLMn
00YuwonmNJ7TzXsXaBdt4mNOwsx5z5DKSM1lQPwrMJqAzQo/OU5Jrs9YNj3FZsdA
rcRbGrOHwZvAiOmQnzU2nnWfubVZ8+fosIteQpACBCIka5S9G4ExB+4kyNXMEpyW
ephO2Ihmi/XN/CVIQwzeYoLNNel2iAVcPl0JEKTs8CUUbrHExUKrE2sxyPjk+DB0
nLu1lc/NVeaQDiKYJ8iUTRlWI6Tq+s1npsS+E5TLp9dhdrQ34TC30kmtL4+9zYJd
dSTYIgvAYRgJxdE2N3H3EJoXfGIqXSyA4bFlfEWaFeU1k9LR1qloI/MQ0wiNNX1U
s6CC2LEd05fwqMgignqhJaa22A5djaBFEl0ebpoFPv0VFYRdeE/aG9Uzy2S4pB3H
otHdxkv0zFsyvOvuj2IMOYP0Q7Qs8m1epx1tYk1N660lItKMxqjGTbAgHFbhvLKd
xcZqqQcrEEWkN4ao2mAO4QzfvV6cV7mA8b8KeW4Tw7ejTdANjtBbZnResmUSPj45
d88hb3OS8TZ1Ygw0szuBMOKVEsDnafpfus5Vv4rxo4c+TXToTo4M4ZlMXiwjQMF/
lZ0jRTh8sB3IseZS2v0sDZXOeCX9XHWWlU0jUPLfkqY1kfrq8kUz5Rybgvl/KJps
JhsQohIOM42QySc2fwvjKQdm9yJHghtHoMkL627nX3XjjlWRRkH792chMwwYcLwY
+A5KZNULpRmYUIkBm1wVxcDtxpFsqZPvoikd/dxDQcIUH+0nh+2l8bOyLIQN/icZ
oUt+kHlrshH96gDUjNCcGWbkjSboNnM8+2KXJgg3aiDrQf8z/NhTa2iNSwP9pQ/F
xVctY37mdb+pPH5ZqD1QoNHbFh/YMmmXr+YOUwqX+bGHYYcpLvK+yMExKZOFnwwF
RSxAjEL27fS3nSEB1skAE7vqxvUNKKo4BOKdL7RseSnJwCvbo8YjhfxsvSeN/RnK
b1HOBlscoAsBHzF5lm++plsvv7QUfSrP4zGkbkUa1gG4Zthpfgt3TFlH9JfbSvWE
vSyFU7c9/i3Cazw7qBG7PDguoLzdK5oEEXgirka2T8IPoaNmADKQsiHRs3zN4V8H
3AoniHtvDIr5hfU42TwFI/bLgoaagw/0UMggMxtCyY3p2aIkDbiuF5ZC2dVFsjUN
lVxubitjSLQHip9/yyHN1Lecd6aT1uxX1agxWLKeemLh33t1gOyqqmYLwAKywc/K
w7O1jIlcThMuPeJ/L5NvJOTmFTn4QeM8xRentrXRhZK6IN/0vGF99riQnzfCLTrB
+9NjTzOYRL/rK/oZVnE2aCkQzuNScSoLo2uHKEeBwapip0n4bqv9zqI88oX6Ww51
Y6SCtFlrrYrN8e1Po429LhN/KLW4cZIetCoVbAd0xguGtgneFJunmAdkAIPKEqGt
5OBET02adRfSKRla/u5902e7SzJGh6H7M7bJKlB9YXpVkHID3DCuGzvvBdvIsAwh
0rndw95ZMpluIWr2IjpP0zyJ7V8QHiLvZqFqoL2gYNQFkN0IiZ9HpOY7BHLseA0Z
TzZn9v5B/H1wRG6Cg5dPGlPdO95squmTO4XftqZmdB/pEeRCZPcw+PVm31E9t0j8
kNtFC9gFqTGvj+TWQtcv6nHOpLML7kgRbUp9AhTNp6uKGh2NoPGr+q6gmjX6KIIk
pezlxvNvu17Ce/UPYhFPrurHmyko0curRrw6iLLWz3okHfmXgSxgO/iQJhEqivKl
ppQqXzZBDAtCiRipC1lJmRxMADHDO+vvsFFm8GshwRy6H/D8l8oTs2WzcRYOVG7H
DY7mkWODgoYodisxyNkkku2jI6L0QIZqKChllJCwR3uUZSg7J3R6blnJo0KkP7Hz
tKnJlR7FJwOzSIk4JaylwYJ+lWA1P3CE2IeUBfwbNV5Z7L0BzdP8lMykBccAA0l9
eri4kSXNL00NBX57b2GEdY2f8CaguQ1CvqfQmS0/uYYz03vOUTlnOGNbLxe2EXu0
uGy7QZ/ZVpPpZGwz+pPtk51Lmevo1uv7dHINJYAsbXilf/IwG6xVtr8R4tu7tcld
NpUDNuiv8Nj3h+JoKR261rUyY3gJZLeajegJNm/fU52wDeKRPHYgimLwhpjiwDa5
6mpcUu5Cw1tCFFaiNkIMTxk8IcC9WmP0sF/WMvCtyymumdFB+roHHdaokIlLvlH3
HgCP+Ljqdn2wJ5IRM4cqXVjtpRADwUIkxpd3HGBGpVKuNNCXcsXs92pZTFdCQyfW
9Jw9D3rPYZPRwk+6K2SYUQstwU+BmSMCJ/GqGc0fzjFiFh6Gw4sNdtla3uzfsZMH
HavNeGp6UWT2Ig5oLIsugD3Q/A6Gq1pt5n8DyG/w639yiC13vuT6a4pw4VzKv1T0
FjF2YZpgBDW7lm82J/wp/H9CL6tvCDhUacNzEJkLa4v5mJmh3FHolno7ITlCUQwp
FUp44Nt+uFP2aDjINDF+C6oV31BS6DlYYD3pvPZ4GYwWfzI8gkxHv3wpIlNunAdZ
bw1hUdjojxus9GmYRb3bIs9rJEhRxFBC7PN8xOBSHaY=
--pragma protect end_data_block
--pragma protect digest_block
nfDaYGhvuKM4vL6ETUjKw4skuyg=
--pragma protect end_digest_block
--pragma protect end_protected
