-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
chg4UMkY+5J3JIXufALdcOznXvSqUXx9wPCf+gKt05oJL8WdPbOqn8pF4hKZRMXi
6xDOg2RIkXdyxzi83l6bz5k/I+yyyrwwv4hlYYL3nHnFEWv5S7P7fKhwSP38Myo9
as0KLxgYPK1eVreBHU9F8TTKnsdXochXDG5cQnVVrQesSVOOg6KK+g==
--pragma protect end_key_block
--pragma protect digest_block
xxbRw4iKy+tjlClEN/vOdDI7F1Q=
--pragma protect end_digest_block
--pragma protect data_block
VrC5bA57mXRA0PjEl08fJbjL8q56mOP2wRJt4oXuPQpPDgZkBb39dwLxVcHKL63K
xvrjCIFT/UXgtRUTaQdoob6+0R4II+W5b8Cl5xM2yNPET3eHuuCsuZUz5pdCUtYY
iyYN0igiQucpQyp9lufPPhqkZxDkXHIJhpATzlbxkCtbDsQuJvWUq0J2GTGbKKjR
kxtC61fTj6MpA/No3p/7jd36GJidiwYND36Q0qLEiVcLxaS9vOsStAUEbYu7tjSZ
siWpu0jpCH0zH4viTdQ70tyGI2AWSDD/AtZuJJb3IvKjgppKvF8QzYwIHCucL3FA
Uw4UVhMyXH9s0dzDzxZz+KNAYhl9AsfjBdvjTuoSEcm1RaJqO7jdqooZgbxwsX+T
5kPLM9LnDdS/S6ORxAduZ6PrJo03+oTkj6km045WxlyT8fON6f3SJW0BHjaSGSdB
2AZdqWEVgZCu6kBrklx48rBOx8zPl3x042fbgNLmXBi0z7CXsj0QbLE2+eGOHBN2
eYR5gPgsR4uHehgZPdtvy4x8uWpgdUPOWZvz1C8Jz/sl9x3bBaH1RHlSxwLAEMoj
qZq1HQWkmfvSnnwvUmw3XQQZFKIrX0jKivNWluwBG0XT3X81Pk31SEynf9pkn1GJ
iJ4K6Y9rs6pBPYFpQU7CZIrDR5J6t7JNaMEJpE1aKRbPZ9cojk482PZ9TON64mAh
fquJHv/g8HAXCiB17p2VxAIXZp/klzTcY1LG8drSj6nqE6KoOdagSyuT3jY0yE0Q
rS97efiLbU3w5nMtb/jkcA+yVnvtjEK/jwHGcTHQokSASeI8FvA6j+feom2YTe1S
vclPbyxjtxuWLEhWqxtSWQ7ZG/DszOeMCJTYHwZt0bpA9FMbKIwzOGnuWkPrYvBu
jTuoteQjcKI373UvBY22QS6z8oqcLbBFoL8Rs3pQGjFZZ3Au2capsBZwzNBib4hg
6CKObBuTFac3+QI5/x1RoxUyHFK90Xi4cue/0IYmVeDf+7VKO2Zk+4Ul7VgJXP6m
qofXG94c0kW/Fyy4l9i/APAFmB93hv1R8t+2QcUtAjDVrjMnVjZl7UMzF/fZOiL/
GLrhmRtZPqaPkU5JxmnbMVGsOCxmnPcsBn8vYOOHNmeF+nTuX5jLpHrLHV/uW7xk
L9fdCkD1JqKnPVP8yfY4knXnGxrI1QF10HFDHm3qrQCRqZ5iSRC2moEYXic1U+v/
L3SdbXYCNYi0beF3sMwrMGefIHqOSGWBawSzOwyTmt9QScl1J/BgZH54knVcjJl1
a1xFHpQ3FIn4q1csMuhUsqh1kGcgVhbU9fOy547kDml78th5Pzdio25PnZBh23bn
a6+6JaoW+bDdrj/8qA04bQ8IUrTo1iR1h3KHvqqQaUkKNuDzDHW6388tTvxZ64Am
mksppyqamHP4J4e67tTkk+zO/Sv2QOdN0YbnTAc5ib9eyCChs8TRosoSKCSoD75H
Oi2pbBikjq2UbQcqFkBNPTiTkPUT1hXemPDDid7H10qrmEAdDCrAPh1kKNJMA7hu
AD/8uMzTxVAZ7Wi7Xtpt1qu5j+V+abctbiVUd3VfUX3ywr0vm2cLBs6jrelg5e/N
UCR5nR1syxX8YxOOn1inrpu6T+eNQposxyGpRhWBaCazm9mRQ6BS7LLKweYfhn7m
Y6OoOLTIOLLFEPPtOuMvvhKLrdxaWokG5/AePYR5xV56Grr4Drwwgt+LLNi4szYB
hwOmd8oQXlFfkYimySCAFGeZ7fj1HrdyW1rxTTnEilaK6jeAJd92mc9KzRZrzN4f
YU//ARBeqV2jsZQYJ54wpKvdh60pTn/otwOj/hQPAWueRzfRAj1pphY0aD0UM+zB
dtcb3+oAxeTbbhtVYXOTh0oVcEgDLRTIwTT1871WowxaouZI/EhvWDSal+8KQOPt
sFU1iCI6jRukQR4Tfos+JHIrrpBKxDu4R63xhPmg4i94VnLzNipHu9VrPBckZMwX
37o1RLQR2aeBURtg1qWNnPrNjYuxbZeqXZc0zaeWw0FR81JWNJLxPm7Zd4A2nwOI
nmW/Eg9c4pJ8gazNU2rcGq21ta2f1wpBNdarZXdmViFMKkJkDnDeAXgrVf/+PFZK
RGclAhlNGKNPJn1iVtz35g9O8+wg3ZA6x/K7vMEAr1+3ZuDrLttPArqIZVNhF3us
0X687eppXAY3vhwSlCZL/pIhyfI9ox/v5i5BQMsvmV+zy96sIVI3ntuUsbrc3z8O
fU4ALes/sXHUyU6UYuQUZaeyJITRb8tNrEX5sQAaLtv6xx/5L0Y/yDAnHDN+TwSM
KEHZ8GsNqeVEYDcdM75Paz0NwOdQP5C7QpH47aJEew5Vg0Ok7qrCtp0cZbySjg1/
qYHqSDCoZf0iiYhmRTJgPASGVY1qZZk33nxnSkk+VzfZIjnKS2V6vY+LYgYuUQpJ
EBolJzR/TD+kHKrtwErrYYvQVD0uAACRi1KpNPFgrzP5uYMckYoDaNRBHzzBa4vX
vIt9H60EP8QXTEJ/SLXWeQ8eUFqSN/0WxWmGdW9sxzHwYUwvhmCBuLqJybQOYoxK
4D4vztAugyzCkkZPO4JgaMx6W3Wm99ckOpYKCYz2MStePmt0gRrV43N3vbpMTiBm
GEsdVNJccQb09Fqry5c21o4FOKPwVha+j4m/HDInPNxWCzgbmD9c46gHlnZ53Rpw
7eZMJc2OMBi6NJh9RJ0ZHLe5+84wZuGmLWRV39aMY/Q86YtrHg4eTaD1CY5l1zsG
lZYPiSG6WOyeuY1d6kFE22ydRk5CcTkJOfns0VC6JRMu9TNrMCky1pzhKXRC3YDJ
yy/uIcinsp4l0UOEIapBKFOO/98RVViGoH8NrjRkitdL0w7ZEN6ZPHAs6qCGEdEA
w172f3DuJC08pCB3eYMidJSKHmVm5/LaObzkj6Dh0MvGpRPMowsjON1a3yRPUtVQ
owPAJ4iCFvNlrlxe3jk64jOlSl4wrKvgknIRcDli2xddMH3M8CyHVuyruCTcYi7G
O9E3Pz3E3yY8b5emHPNNDyQMb+9IpmdjDrblm9gmmJcAnxlNAjLHZU093kpDQiUU
h3lDTYRfPD4K2NpNEfU0zeV4GRcA4hAY8mkMnXs459PZS+emvypqLnu5vKyfB2hX
VeiH104s2ZjGM88lInOtsKIYfzQ3KHsxq87oDjqQLe6mZ31R6YjXlx2C6VC4kCpP
TD49S/ex6CHaz/DSUyKV60h8gF3qhGTlSCeJZ9Qgl1SUWJ65HZmFMWJHfSdi5G0X
5UFWaagU9ABm/fz5MtIgAPkOhssESJR4rCMFFaBlOiKI18XRbCCyGw4N5lDqlPIQ
0D4v8yoZPH1JZ5Yjf9pUnCTyIrhJf2mijkIRfZDUNdmggkJdYc9ous/D5iymcYR0
FGTrdvVbBjuyJUzF4LZ3gVeHICgfojOsALt1zbxZQLdlQfE3AYrc79+87PzJ/hQt
spyAAMC4n7b/nBzETg4I/XJwwwQoPOzOmxFW3OR76GRRVqoL9j56GQY5CjywS+xM
OXosSbD0FqHPJdPDYDCL7h1i7NASK9TrliBB5mtY6OdlQMdH4VQPw1vwoSdr0nt8
2b1x2VhD+8tEznGgYoIn9J8vsUNXU4lyu9hqIzvF9zikugvXy/j4P8lF0ndibt8p
RV/PxB2u4EqEaOhpowPABvRgq5tRMjTHdBT8SRRdfcnR1/R0uvi8f2pV7guUKNy9
8Efukc4YS3JLKMgzEULJ1GCsUQ1N1N6ZEhdUCDHZJkPY312Rw/mJOGYaM05xB7A2
xyG5CpUc5cXnZOBGXJNL5g+fjqJgB6TLV3sXVF3XCOTo/BDa1o4xNPhwlUxebzrL
O/cllC0VnDCxcdl8/s0b7l9QJiq9aULakmdHe14guWe3XAsvK01Pad3GPutd7KtM
EnQjjxQbV/d3Idb4JfAX3+BsTVUAsZ+z70bcScPHmX9/Y7eIkKnQwMLr5QL+ZBCu
8jpwIpDktsHQIzK1sSL48Zw6JROJWb+sa5NXK2Cu3/AcfaeMzegHiCOXdoZplvit
W2ZWkYiqxVBpyDVzy2qqwPfD1DugpZOK4Kig6zCzkAWwdIIQGcQN4xsr4PS7e13E
1YjWeUDkywXbhIKYWLnpST6gbQnXO0MLkGf2Jdy5VsCZ6Wsg6HpYjp7cEVk61PGd
q9MfiX60aB+ZOKdaVinihUQqo+yojzUJFJr9CR5RKoPqpsgmz1X9FsQBHhdNQIss
AwedJlHVq6+3bDVoXodbzDPnuFaY85ze1rV3r8SECYu/rj8cyS6NfFa0ehR/LFMG
1dW4scTCmKSuz4oHjO4WsKUtZwe7bxUlwJDJT1S2PUDpKvMwvAXQshjX8wUdaww3
aFlzns3oMsu1WWA03Xi0nA1s4mC9829Z7jmcrWof4j3EpFDYSZ0hMsjKhdb5aF6/
vw08iHCeRZ2uZzyJKFxvH1poag4R7QKsHu+7qXXEU0dqNA5mCOkQhMjd//jahHpE
RD7GF2O5zL9hRjxxml+6P1gb3KkfdGxxtDJkBvv6ZOQX6eXygbClq312dQpfNBUc
hZMl9zKWHAEIJaUUK7mT109Mr/dcLiKBMiXq9d2MPAm8lrIdmd0ideVYS15DQPDD
53ZujRsc7M3nCwhYN3iC5I/44PpbrvQgg7WmdA+FesfacnzkfAXpqiRIa3+RkqrS
t20CqtzfnBzrMdXLWGAfEBu//eRwQ8TIAoyJagJSDNBGXKCNADHiY67/UY6uXrDB
WMLlhX0tAvopBASv5lEVMK2uFoWNqlFya+mLuGrvzZiZetXIeJXzmRGyrHrN3c6O
5PEqBMEahWktMOUbnmDGl7b5bqvCynKHjqSrTZzzGuxLHvV5D7XrmYMSZkvGJAtU
Bc+yx/E+2H56GTgnB+0UNd2jDYusTkl1KLpiTWa1BX6Ep4XYNQL6d/J+wRVKPxJm
uTtuOgf/2O3p0Ds1q6tCH5kvwGc7plP44cO0f+INKtQ2T/1Pk9wjROmc68GB5xns
ppX4Fm2JHNNXz7TKPt1SH7mIPig4GJ0EHMlaB+KBNEv/stRaMnVMgQWqIJkQ1dZC
7Qd7lij42fiNsGc38n68xy1slyo94gdUBEPUuziJercxiE4lBigbLuBHtPJw41dE
zHgEhvivqtchz6L+J1vqiUf1qf6Q+koDQ6WIqYa3xL7SfXrZA1dZnh7cuhQisBWb
0LlW1EASypmTNs51YBbUQt+6DCxCDtSRon38QdUn4S67EEwCvh7Stom6iXlHs2J0
Gonnt3l3lwSUdCAFlgNvSvrIiMhgK+jUicRBsmx8JwD2QAxvIClj5KMS/yHSHYes
Rclv7lEbyzhHHT2y7X98LrXJAhSHLpxfLk+XYbTa7sGPA3NSUA/G4mWIKPfWI7EI
EkBh+dBGf+hQcaSr6hvdcwFUYUacRlVmGzTFwLmpnixA0cNMD2h5gCE9RSJBYE8C
A81ssLSOROoNJ1KnwEnbv5ntVDCjXqOQnl5Vz6oRqyrlNS4ZHI0MG1R9LQVSdh3I
JghyfYQwqbdjaOUGb5kvF3rXTAd9u+aIA/Tc4iBtL38wI9s8PWXNwZxShINEu0cN
60VtnS19CLma8DGV8im7HqEXadRvPZSTOcAMYCX4hq4aeNTM5lUSLsCcpsb6Muyq
mF9eTYdBluy+7sMPxXFNh00qXQMFJ80LWnWFZAjwA19YBtV3ePeFIW2y1An2Q3Zq
69/DAY1+i8eQEbmMJPfClMinkfJqdW2JrGqpBjoKEA8MjfgQgFteL0SKNg48v9c8
NaHy6oLcSvbVTKx/yAUyO2ZoHtXpQUPPiWS+sNM81Pvp+Eu4VmeljEFqMu+DQDrL
AG5tjsrvcM/n/DnObMLL7gGXH6PoM+EMiXr3UUesODIKm+foI42meoPznu0lygLh
BiAboe8UBoKAxshdTg12tZnM8jqezSBx3eaYCvKl/7DUxyI5IFuJpM5xFYoECAD0
iJI6sZKiTnbsgtCNwAqWrcS93+e/upyDgpVv1nzmR35kkZspOkUDcwhB6PDAinq/
5kUt/ZxESqzJtUGNfmgUXFT2sdP2/9QOzzvglC8dBKuASZ+zgGazGryKWcvhVy4y
V26eFlDJKRjIpJbBlrwfmQLAPcwTERh7kVl9RVgC0xhHz5UH5icDeFMjx/gF0841
aMg8NB6u1ZwDGzjo8g3BBEwfTUugUMRq55XgYG81d/emxqqxWCY1JdzpX09gUVzk
FMdcIspjhaahptPmz/hc8ZBMefodJXzkaTk0tfb/zsK2arhrJJA03LEVlrJfI+z8
+YQAVzXe7a7FMFVA3fvpG9GVTcEK44/oc85m55tuk8/ldikmbiOI97PpDvxBjpiz
+mkwk23vwUxRlR73nTht00tciQH0QjCql+b3AZB0vSiATr/RsF7cEdtp6LoydJZJ
vFa+1ki9R8C+H1X3LKI1cKckIEdKUgde/g0CzKFVGI6fzycuI1KO9WGe9Ffb5I31
Zs6sPfH/EHfvXoXxV74pXT+ridYjTuHOc6NYZiNQmQ5DupMJ4/8MXq2oY82Ltohc
pZ60LXtmoPC8XU4I7t7ywkGPAfgJ2RTPeKL4QsUK1BGqt2+OYouFdxPMJMRFnO4h
I2PkQR8d5jBcPUeqqi7YN4nQmPc1QOCr1usbb9Bmw4wm1FcrDT6Ai7sz5AzZ+nsl
6y5HaunBCoylJ+6wRYIzBNvHWEQgMj+/t8EUpQ6ChfFf67LLxHam2x4sxyLg84+X
Pl0swRCnEh72mqdIt9CWXj8XLWPnqnDaXzw72T+bstWn2LR5OuvvHRoszXwha19Y
0U9QoCnK/ELwAJZmsn0T6sTsemc8aoSfqDTKNwnWSJnw2FJ7OMGW78EANrkpvYFy
Lu/kruT4njpz6XyXxDCEy0EWEOHmPOjtwTpLb2v0LQKdthiSc8olFz7xMRD5XRvx
cUFrvGYA6cmB9R4k82wwm/vVucjXu8W3Kyj2xadeZr67ppkToCrwK4K+y3ZfIm+T
c0FNa5trUgvL2YjFygMLD99PsZ4DoWFS4Vx3g/NPaD3X0EoHs89VENu20CYGH8RF
sKHC03/fZ52vOojzHKVXIWmkNbOBzs0EgWm5XwSq1zCyu/UYIbr+rFGiF4+DKc98
y4Zvy/q+O6KnkR0PUl6oON3qPjpDxhXURevywZ4LwhqU7h/8QDZxoNdJvhRg7piD
1pZF0WOXp0cG1a6cd64hOFUQxvuhsQJI2ByGhsL3KEFBW29PcmTyInClq3JlX3mi
2Zfuw3RW1+Qpjk/tNlYt8aGNaozDLZ5koV8j0byLGTRZ/INmp9UV5IbQWUOHzked
UwAh0nP9/FhlOD3mriZDbYgI33K1HMt90RGPtYYUSmkGtTWn4yFh7yUZt7tTCEuh
CfeFtRxCD3xyrEQYrfeecttteBa6kjikgUuB2bWPrdk8JlMSIzTFKb8iJWr3DgqA
LkhuL0YQD0Yrqf0Vgh8juJF02M2SGVeUzQ8e7YBmHeEgSv+unLyjlGMAeSWYZVWP
HFfXTnfbiin9SHyDhBBxM2HvfzOCb5kBbQJvqJFChSHuj4QAnSLQTc5y0duNnSAP
XBe+liaIdH+6ntNBA2OPfA/Nc81uB6lFQvEG0/9idgrLxp+Qeam8tbSzedStOzLS
Q8jyOwtGDZ4koZAmJga7kRqA8t+4+J5BNrKtjic34yime3mPAYnoZCkFZQ2vKnII
/CBbyg8QdmpgxAQzRRfRKM2L/ER34/zC9o2/tFqllKp+m1Y0JXdCkTK8Fvt1xIll
S3YSlclwT+mM2SKoZJeafNrfwfItjwIBP/r0qfzviTlUDtS2pOEc2qx37HLGaouh
4iPOJK6LDPAXUFdZST9+BKo46JKTAuTFVIfowkWFXlEnC5WWx11/Dr5d0E3nPM/O
RqXsghQ+uckLNVBBh0SrBO8XWQhj/M+0CmMk5KXoZvKdKBKsSmkB6FObkuje32AD
wJobX9D/cwKAPo6cP08M5mUBPqnsrWh2Fl/p+n2K64cWajAWXfgt/1rjpwfpF3UV
7yXP1y3iyfJGZyO6/Y1gJs9GC5YNN9PV9sUPiGfDtr6UEbs5jV/hIt9OXOnBoenU
6gHzBZhKbhz51rbrqU9WfVQ9XcQksxVbJviKVwUhPTxao/cmnFsHz/Pq9+MaxCy9
yrH5efiTZQym8Inr67Yrq9KAj40ZcnQx6YeFNAkQiW/Ebjk2OqYIE6GzV8f3eO4x
RE4HBUjGKme5UwYDfJGtToFkHroBZ4/ug4Q7AmQjTabIqw3avFVzOo59r6cSFuJj
F0RsFjJxxCX+vWnm0sqTDSkmt5seAEgdX7WyjMAHmdBq5jpeAoUpt4m9jPoJqsUS
kArozLjkI5IxEBAIDxgO7CHDZqt1yG192Od8BRpyXyaUZJ55kScuNUXuaIekIu/8
S2gi+XoA/bErKPFzqIoYQQo6TIFCgjVZ1TQpzLp48Iq3q3WwR/1nmC74Ib5XkhUa
p1BRS9Hj4Lkafly+4AI/oSrm4yzG2fOXl+qTSfgEO1rvur/Tr+NN5tKc1F0uQT01
xnZKt5MLmvvLUoh2oc/YS6rQBHbfQj5yFszhcm6M4qXcWOYY7rRVUaEJM4NzlwM6
5KywHCq9vvDAgEdixs4kCoasB3wXOBAbcX20hzQU4wfeIiHDUvhDG9DuIeVaAysI
b3jc0GyAtR+im4Euk8neO0cD7Hg1cu1HwKVOc7bB2XjX25rkh3gudNOjYZJLsaNW
tOST8ddOft4KkX6wCuWeUa/bhjZNfqrNDC0pOmTpI4X1Cuye8ItS1T9jKxw2qH2D
8zaLYNe75F6GVlxxfe8i6JOleN32zcXofZeqX3KDVN6Y7LS23wj2O79I7sJoqxQ2
IVpULiwiuPGkvQK6IXIY+iPdZlcgHNrf1vyU5aNt03vwkaP4VrkScvnGK0YyjCyB
H4zrj93DYbsfUrlm4DDQJ0aKqz2L9z0hi1551mqkpWVcCtM6RxEkRyMyqSvSNjmB
Olvc/w0yH1sZht4s03VqMugeOF3sXYl4O7FrAvAgyIZKr9hbjgig/2X8S2zdelnc
9G6AO8lN6rEQM8mzFwlbGFHNtvdU7xgQb6dDiE44MDpbaSIznxoJI0LRlErXnNuZ
ZNTXZhpK/dnuA81+ueXxVC3V1VNrTCPM44ER8UOT2a9wwNy91oVJuErbzspr+Qo6
66lm5LgRlp+B+OR/WnMFDMhzIXPrfZzCmerWxROJ1FeBcxLbUg1q5rF9C/ZeYk+k
sTMGmxctEyXaX9UG+o8VM70XflkJ1iQu/y6FRsoa0rqAhc4v4pDvbigG7E/606SF
YPiaR/ju1Se8ALQ+BUumtg9MuGapOU/QC9qkkzwO1e3b8MwozbPoUB3ubv7dzn2B
AyLu9AIs7fwMzTK/0FUu+qdlC1NmP4wqnD0lUTIyjmoGpK4O64Mr0sKX32fSKyam
f2QPGN6dNVuYjwjc0jxRH62fAK/9Qzfm8L1cJy93zQ2FNPnSkeZ5HK+RlfhDtgzb
CUx65Hzo5kwf3l0tYM7k8GenzMp9A2Cc35Gi52Pm31XYihO7AzpuHrIKmQHQ3fLs
gaWQY/PPQaZ8OgBEDklZuOzUNsHtrUGdBNFZf2u064bn+QDfQqQQED64d1avr2rb
GOMaZFYyn3mhyVjVwBrmidTNfuHklth8iTx2XnI7k14kiD4vsQ1zV/52YFxKzcAz
jnPj8YEDyYNRf34XKED9kMp2N/5pjVrTX4h7AvCmkla6jOCIOoGG2QJlSSzzEyuk
E+SjpjytuS7CA7hq20FzBABemtJgQ8xoefQnjIACGU+2W3xKWW+b+9o1hNhtryGt
GPN4m/0xxguLi28U53dXRwZGmprmWnSrAlzLoEWLtctXZYFEtGkstTPJE6Fqxb9f
aaa0oYOjwLAjnut/ZvwVeX1uvZEeiRSVOyZ5cx516PsNSoU0o97Ax0I0T5aLT7yV
VoZ7KQGQiznQ2lT23ate8z3E6xfu83/fCPZTouoQDr1usIjNdvSraYFPhPYZb73d
WyQogb1HeA4qzHSvcapUtkrT4PvchPRnx/rJacMETFSesPwW+PyUHsNX3W6mF+L0
h3PbQIbkeYRZs+/a5OQ0aEucgpet31Ou9gOnNO2Dgra1wFlSj/iB56zEwF1L8n8L
i6MU+rGQ/8xyA77jLRea50jJzN1XKzRJwR0RWWFLhpTUWAHinUDhBRC0Hb7rDywD
M9R8ZAhsr4NHLhKoYygfU8BORc8y9NYyii6BM8P3Tual8Thc5fnd0Jd3oqkpDYCT
y1eWBc2RL15r5Y9yUxSqt+qPxJMGZOYpDKxIo1CwNgbQPxQuJW6KwSfwFLD+GHuc
FGcXznB+lsWOuyRep9tm22flN2XTVOqQI9KCCvBgZLUok6pGwmHWjnHiwB8eUY3y
OBefmgk3W912gI/7raqVppWzQnp7LrlCB7atj8e9AqL/jTwe/BOxL6cLHeBB9FQY
ugQcTnLRA45+eUcZusIUW2Q8siMLF3ppvd8Z1Pft60lUiMYU7ElihYzH4muQm7ro
nVywUJEco2foBNcQbswxItnGnXVmX0UbrL2j5fwijMFcote97HlJhcVIAp5h1BuB
2V83NmGqXAswlrEZVvU1bPJvNCxj2R/EfcEEO/X0TEf/UXesyULJ1+HU4UGgVTuS
Nbv120mnix725al6SPoNrKqABeD+3Z/8ZkFN3bvORmQJ915Rribh7wMvVEJUNX/O
4aIMSgVHR3a/AWJgR39T0cqb0m7yeShGDUcaOF3Rl+L3/WKg+mSTwDHXf4LznZsz
xW6nrW+iaqT8LBGdEFHQwRWzQ1KVClXaeyyn1U35QVYOl3teI/cRtiMqlaFoUBVj
/9++Eu5VfpPb5shG7wMJegWY43CNI41sbQvtHyhce9iX9Gl/wlJic/W83tCQ+OXm
d0fGOlCngVf7tnQqlZgt/aAMju2KSOzwsA2x1NXjEBpitaKZXwCl9LE/0NGhOyu3
5SRkBLsvuWak3PgmUwhqccvRsA9r6LbjmS62ut0miwf2VU/FSpj8Sj+1JjzLdi6v
q8DClmTRN9r3Z3dy8ay1v/IenHp+kH0HZEsfcYGEj8nBxGOlN9BjNyk2KGXFVw7L
meb8FHhPzk2n9DL+h/zqSfX+e7DmLHlMJbqrc3C0Swbivm+yzX2ONpvo/9GYiiol
s9+n0g1Xk57QiGGc092ymZP3+5XV4VBmJBT6BXZ2f+2T0hPvHZybCZ5ZKaQ/A9fo
THzmlrpBzela20E3WjvzQVjSl6zwt20iOOHuE/pwhiv77M/kk0CUWY3nnAm78w4P
/rrAyMsGUJVR0P+memzDhToo6OHvxq61PZ3CwVYli6IS/VnZS+eGukjcmuIitUV+
dpOYDQKhIW7JuJx7Sc9veS6fSpJ0KJCjOi3LqMF79lnWVsB9Tr9atSudM0ep6MHF
eukjIi1ikFdGixEXUAy2wyT/AaC0wbgNJj4i/sfMa+o7RdRikJGK4syzHYXOaCGu
71s0aWF5AH4WY0QyAVUoEkiMlyo+oAr+AZdqvZw8ZrbJSfvzAmI9lGZRT5y3kYk5
8xk8rZwKbW9t+Y8pZlsKSXwdFDM+5O75IPD4zBoJa7k/dLX3QmLLdwa8WuSZS11U
1+jrPlO4h8eXccl1VvIYA262rmr84ITE6i88zyb7zKH05mymPezdwINQ1Sj0mQxw
zM1pabyb1duaFUI6l13NkQUhYRcffUDzZJ+RuutBu7ucW75aXYxZPqOlpG4Mpdj9
4itpiDJOS1xNaTL4GvttaavEIJ7H2Fz89DY+nUCNhjuvYJ801E1JhyuL/TOTwwSI
3rLoT6ZZLsA5MLF2wbS4B3AlMnqRZ0WdAUWi3aYGqAwORgwvLwaN2dM4FyFMqBYh
mThGwv50Hcc8e62+gv7Zqt1CxSeCi52D5dvxKat6w+Ly1hGteS8N4rISoV9VFkgp
qAQk+dPSs73Al/bR4tVTjQqj1XG6X5/8HQskpnJx5b570TRIZlzIFAcBQVQBIpYR
gSdBB+jfPng6xVMqwf1yhBnVH+FvzWOtZ34FME1IBidgOQDr0S2Sh0dKb5OXUWnq
Ix8UDDJ0tLA8aZIXQdVhy3yWY565VKfCpxBXaV6zIyzZ4dgOsbM7pMMPpOCOwWt6
ge6LjmOfeOM9tKIXMquXuZm/NvR6dylWwat+zKZH1ifi1DnRxEUfRHRT1lhXCwEA
8Ef+mHG0BrbWUQKL6phxyX4RKIWUeIgOv0Wew3FdzaukSR0iT9Gh7tJpU5UnSCde
dVGwiVQtccs8Q6Zv7GKbMQyZ3QbKLtbV5hSf6ySq4ixkyLeHBJcRX3XNgjqCA1jC
BHe9nhWyGJauYJasnnle0IpvTOr5tn4DEIs/05/YOi4HpXzkHnXJom6CFeGGAANU
tsVUKy+b8+DrvgYF/mbILMhen12y2EBcSw4J3jsClbF9S5GZuIYUPVidFagWj8kV
FASQ5h9yzsW20heh5Bk56xnH5msfAjppPJ15RBtm4nMbZCuQX2FiynAe4Daud8Vk
B2eYndmRlDbuRjI8rPBmI77HBX2RzXholDajc9zvPj/8FLPLf+bD5qXdKi+MplPZ
YBhKvuPPNRSi4thqzFhRC4i8rl1iaKuY+/7UQb+6NJQ+CBMWpTbRDIEKeiacIN9M
Bd5mPdauevYdh9WyXjbw9J98dd3062gTzYJv/mSDF42pOr/pRdmQ7g/A8wW8aeIX
vRR39n+tWxhL/SyynN7Xtc712haZPCG2v/92YhIsRr87dOkIVFWL/+LKBSh+lN+Y
z6QXkuJZC+Z1Yfws4XdVyffbEohq211TAGfM5bq7Xo1wLIgzrcJEOIYSEY4p/KY2
wNwSotMwjIQm8oJG9n6lbJ6odxLpT6kVA8Ile85AXD+AO8gyOYf0C6+odAERy1+4
U0jJcWQ6e/azdcmf5I7lYk8yv+BN95KC0E/FCiGZjI7Ry91wyr2vHL5NfBA5s0a6
G2S/hmLKhMwXnVEHnQNkKDabYu0+TzTqd9ggEbB11rnb1EUAStBEzQuPrpqt2AmK
/QV5wRkjh3Jsi1tRTsrOR2o6gKBGf+t5V0gJCggW2IxD7vyEws2idbmdRSJIaeGy
AFAD996emxs1XnNtQ+sNX6xUC3OCcYHTda0cDV1bPFJv+SxamhcO/qjMIlJQLoYz
XBzxXytP7LOIVNvz90pCfqDfzKVO+XzowJZ8MziWtHq06/MT1ZKkUnPLuhn+kGLK
D4tnkvUw0v9IOnFKFy69i5GY2u2jS+mTA29MSkO6FJqIjR2JzGQsPvtqZP2iReep
2iWxXqOi+M9NdNB22feP+oUsXFq03X35iwXMEVqgtTT/vXVFkNpgNicWYnDLT3G8
dFOwYpvX4N55hVrfkE6UBEI6Kzz4YQpO+9ZjArqwU8+7twk03D6AzUTxhS4yV/r4
V/d3ZZmgoAEBhsQ4kvSiUYW+ujeAcziAmpYb0spUZ46PMTvX+sEi1oREkHhc1M86
IznEN5G2l7eX94JUeAEOT8Nz5iT0FnJ+pSTiw9hR3OdntadbWHOjsB9Ka3Y+QIyD
HzSRD+Bg9iOUkUk0eAFhN9ruIXIQ5iO5ONMSsMSunEv869GZO9UfA2AqTNXKjjJl
BKd/dkxbnvbb5w0Bnb7VGMfqHijXithOdtulaCTxMvMGFCMNwCBQGtFoNrjDgOYe
n8BXMtdIUjpOAlahUzSV8kuSqbqmJUKP3ZBNGooaWGlC6xnLCY5JJSXYgVW+brx9
ygkuj+Uz0ICBabJDDt3c6s6HsQJ0A2Fr806jr6fEaJX20PIDN9fcfC00iqhUtPns
moFBioiEyf7Xj935niI/6GCmnSh4mQSH2uODPXG1vOawj3koMuYuFCw/faITK/jR
bilj7EabDvqPyFn/q4nqxB7LJR7jkxygqhtiA00iHEMhqE+F0Jqcw6iaC5HB95bK
FdRU/wbOH7/l0ImCsPo8rn84TLaMhFBB3Po2dMagYSmpv7bMx3PuPA5AcLbX8WFy
i0Kd8EtjVve1fx9R4PYUXW0IhBMpgIjMUZAJ78uotwncwyQC080oQPfkj3HPTgyb
mI2yCTQb7omMwnXYlABNd/7XgcZJWOWAdBMd96OYOBoexNtawV6kEfALt8nNMqjf
Ikd4Y6OihjRVqxAE+TpIrPvrcDsEU/trfosAvafd+hwVLZAMC8ybOdc03Ubvxrdz
T+Nbn33xQWUCsftIO657XEbpPSN2dBiwrdSXeBRXhNtdAb0u4M2Y2t5BfbDfP5Vk
2y308/hgM2dYXtY+mT41rxYef5pkbtfFuQYrSjDMeQ5CtgZvdFv+S7qMGR2wQwoa
YsL3WzqcnhJVAkz9lSez3ZvidhgLm3zwYIj6jPZHH4xVJopiLcgK6yuj2u2EFTGD
Cy+jJXNuqf6MlgkpPZ++JJqAHUuPNsJNTqDFGmH7raOoyWP1TECVYKDBE0+d7ijD
4Vm7yyGSd6ziHSmRdyIjin9GWUWHvhKQoZZDEFv4u5oPuT1f4VkD+SX8um25wzhT
yS+gVqwz+FfptqPacOEKvdFoPFOK35BE+41LN4K1HpzIvNGBYTBU6G6GJPvbluzd
MdtmU40B+LgUZbFe3iQZa7u+az2Ij86WtfgKHGuQlmeaY2jw15cTIMpo2EDkJ1da
jVIiCLbGDCdXK4Ylt/lJqYwl5LL3JHtxE7Ux0B8uiSvSr7KauyJ4wFYcDod7oAaL
jsD3ErmUCQb0P/ssMt1dm1HoW9x2+bDyz06WBHZXg/o/WpnXBAvSZfwp7oc1JQo4
sHnYHPCbuBAZk8ro5zV1U6b9OFBasUJJZPs2ZMRTsgmww7xVBxwftvvtG84L+Rg1
FrbCb35RcyaQ0OFanQB4IYbWtNuSY2zi9U1PpbKHjeBkaBpSSwk3cwmf3m/vePQ6
YXKhpgXTPmO0pZvyNg3vAQe4BJ8Cr2HRNQ6zO4tuAnwvtDjR30r0uE5cCnG8eIh8
ZhjCYG+1PxvptQE67mki0FmmrWCChOjC3+ojQfboPaFx9cF0UlN0hSPa1+DUlsRQ
ZAxzePQxWhUNqx6rXTg33VXYKPd8K+aRDI7UlNSUvqwqtQDH8xZI3DX7mF4H4Sw+
aNkzX7vZMxGkSXuw1FDrETuvBulUStoN4CTq8EBAIgMaGXwYp1VRNw3tK16eNNF2
FgNUigdooXJt1Xcs1enj7/snDjFx1pRENiWCVnYd+CekmEjxggIJCYsiZI7w9eau
2XB0U+gpfhl2Se4J/IYwswd8sF4JrxZgRGDaENRnLxIkNt6MvZmelmbrFAyv3pxr
yYWUJ0cOJPtLi+N8qXawefsiRJLmM+04QKWNn3qtIsamOTolz7eItCJ/6jk7zWHO
JyY5JYPpshjrFScQJAQszLRkPc7GZePKs4BQzcBee4mipVl/0jyLycpZXfQHQla4
m/HvP428jrkGQ0k85PcVsGlxNbsch5rAXPLURNq7iCFJbBfAgKuwHQdAxI7TSDsB
s+M1QFYTla1PBwZIdryqnzA6lSlo2EwTDaJLXKnYCiOwF6bIqQfkprTazL/wAgtk
faFTiAj5EpAQsZOrXKwaG69bklLV3dthp1aPt4hRsbMRUYozONj1rPV2RmprZuXe
AiRR8Rdfb5IevFk6YLwmPP4//uiNsDFaxFw29aooIF8iLq8De0UafXER+xGEYT/p
+Gaa1HbjVhGV8WtMoJdf6Zmk9Z71/ELC7we0hwTpGh6tn7t5zJUoxN7IGbmsBVuE
7ggLX9JkV6CDMsrQeLXdkEaIe7j0BePACJOS7cPOeEWzVDXeIIczcIHMCxfLQYAP
UuTgh7LykDf8GVsczgDWmI023rhQO6sl8fgSE9xX9WqRYiQ9EGUZytSiXZdi1kcu
zeEMJBlTpHXtxQ6xL0Ui3nQhj4ia46cec0127L3gBmc8n2y1zlozh2Y/eyku6bjK
zq1uqubAFQ9Tb68DWuOhgnP2KHNLvpxiXk/UWwzxzov47unm+ogIDKLPFCXH3ur8
YqGj4RoTPnXFZsqbyJu/ic7aNVNMyvBmnvrXoDm5KJJUJBuXTpIpQPFT53EAqWVc
BcM7w/4eDLkSPkadaT4Tgyx11PtynwWziUKovrS/EdamT1Y9DNdMos+HaRMbedxO
rrMXqxMXsEdGL8KbYxxzC2cJxM96EvIDXHALqxCBRdRg5kpZ4eVdXUSQfRCLoxFa
gu/ctdjlq5Vrvidd56XbyRa1ynrdSxTluHR+7aRos0uMC3XvTcWX2wbTfgOqn8Jt
RmP4M7qxEs8Ip2h3Yl/7ZnR6nIZnxTH/vLAL7LPByNgU+4viL31A/pTLKJoch3cB
yK1X/3nQKXAvKtW67/92NCilw4ym4uIxujZSjWBOkL/iYGFnEvdSSmW3hpLD04Q+
Mh6wx8dmj2MTuhfKeu+nrJ49gYgtHEOWt6CLi5hhx1F+Fu3xV1yjqLCI4ZTgZZ6l
jDgmJQ1+ZxTsBU/9dxX8QDlLROx9VXWABgG3AVE04SOG/H8s26EeiS4Qt0l8MEfx
lYNvRCNP0uFi4UdHJJ1mNl83LybtkkzoKlpblH8hUJKCS8RKu5wNlZtKPzKyomqr
UNA2YoWz9V2dcf2JyLzgXJGhyLYruPmDlJcEydnHgw/h5zu1Wg0AYn4SkSsEZS0H
QI/ZJ2rPqn7MIOmJp52svqOu5j3gkRMIX7NL468uBwHHWScYl/wM/aKuMQ0LkuBH
QDN64uaUZozkoZCNIAucJW8JYlZ8jqTtyGz+5/TWGN2wV1PJDLK3H1nwryWTNLA2
RijX/ttiWhgboSRAfGoWXp2xFZTQTNmSJQOIwH1VQ3hMJp2nW59lrqcr5+i4q76v
Lin99jeX+n8PMC7OAetA7mcaF4oGP0j228v/RR6gC6fcloihBzzscKvOGskcGw5p
K9tU1j74RULzF+0wMB7N3lwgHUwaHfUeqkKJQ+jLO5mFoxSmF5UEbfFSya+VhzcP
txF1nmZdA5D6gYH2pZs5eiPaRH9W7shMxkw0LP9gN/ggEZTpw915PSoQqMlwxLIj
KeGJx3pchf868bwRhNX7wlXGZzqBCI/eMWUjwTcsLMPlHzPDRGpW+TGXFAFuph8W
wqlogyd3J96QQSWU+FaOSIlIq7OJ/DXfPDe8oZry6yH3UOKma+69KbmzzBbML6Rf
YJggWSCidhJl3ImZvPLJsiMij+KnDPbS2YmxI7RJK7sKykzAuaGvaSpto3sX3zwn
PhHwONmd44CVAkTbiPm4kHDWRhmEt8mijHsu6b4yYpqc7kOeyGMfgGiSgKzMLALj
7iSxrt9q6Hc+TsuVDSXFy2yapUB5xSIKpXo/VIjClzRFLdW3jD65N16rFw82pT7t
v+xuh2dgqZdCgUg7+FDwk50+XmMLZeBnki1L8imex/3Gng4vbGwcUQpXXkG/d23H
WdRqjmCU6lvPmhJsFDV+eHSa2+inpMlnlBkMrBJom1g9hiA9mpO/nxCR028LyuRJ
pbHGqLejzFR6OTC9oDoiHbkNyrLWiQj1DuoWoV1C3lP7TgGOZyLNqLnEX7YK54qf
C4MUWTj7BzfNsN3au7VqgXzgTAqU0y807pd3AuzoR/SJ+TlmfXlwGG7FFylxJTP2
RwvlB63oHWFQrzNnlfnh+DXufvgd+pZDIzfFhpszv0QeSkzo4SZKquNknCivSeSH
lQnFdTaSnXn3ZvFemlsZWklW4qKuoF0vwrGtr9eI4vvHB26YJ6J5q1JICW0PMCf0
SGGDR+NjzhDr35zNoDSBCp5EbarGoImEMoqOjbwtliTkDERL8mMV5fOIm73qzFez
UZRX2pij0QrnK5XiONH1Rc24/9mAVcqTdkfgr5lJ1Fvuw60n7zW+2i3gELP6xgY1
gnK32PrNCiWqy1Zp8RHWlsqXTb5KYqa469mo/MyV6wH+zvR/dXRqBFxvwdfTDSfL
CMDl/BeQvMX6E+EY2oqnRAxa5/3v9ODBastgu08WugdUIx5fPq2rgu4yDhfhjjA0
juOGFzg2CGEb5pCXbO5Wk2uANUHfqIRfuddVdp8cVFYy+pH+7j/qPUBvlWSN/4Zu
cCMA6ngevsbz/KeW2AktS9x5fh8gz0XrgcVHUUw4X7QITHL+I+3/T2oMsvinpAMl
gYMbkjrOb97z8vz67mpB8JRPmwCSwnjtZHoOMgEHvGNc/xSWF6tTnVps0fN3wvPZ
DDaJkoajxdJekaCrlfOluvGR9UNcOOeM86Vy/0pbWsw+yJoxxAu7dbeJw0jUYvJ5
nJanMRqcK3fgi8LBnuLlJAUXxR4X818mx9AZczaQox3sMRqaEmmuT2teOGmF1Td4
UovEN0OnvLfdkAuEfLhLYbI5Khryr3tZ4zy8ytGS7E7NKWP3+3iDsmzrDjUUrPeU
oirPWeod1db5VUngtx4HqteuVeQMiVATbmwkwdkzvTUi0omnIgI3CH9KC0iLN7w2
iBQrKiYSmS/Ru+LZ7BNn11AgDtX22qxod4dAipIzoIoT85/O3GDPtsuYoGzSOrpb
9bY9S74Q6ls3yZ1YoBhYOPngKdOUBNEUt4ir8u4NIdgM/V78w2m4CEgZQoX2huIN
OVoB3K94gzxSyPhzFBiwCOm4K0v53vO9DFwsY4D//mOculFhE0B9zvj5u2bel2RJ
WGfN0LPcSAmQaibNBP/YcZitHbNVk/oglLjXxMMVnCUzSXUZ0knCIDBKGJ/fgYYo
cvI/V93aEHlndAM+0tgWTx6tTWpbmGY1meW+hXlIQTnCscKIw2TO7iU4teMQv76+
6pbP9Jw/JBdMYNUr2XHJ0c+A9E2c3P8KmMGCbg+ysKba83Zs8+gXwbzeEs0jAXpZ
ku8mRppwOcle6godiMw3vxy+nE8Bvvos9osohp6a/lRPEZ/DR2+tAlmH5x3TyNY9
Svs8EIZXZmeyQsAaDut/iQya1n9bCCDChOVD/r2VsUPeSBOlcZufz0nsXVUnmiWF
cAy0LfqISMTZzOXfNrR6VGOFDjrmdrYSzgIY3uitFvN30JO0/JMFlow76sUsOK26
5T2Wj0tzzBswsknMQi55Hxx8yKra36UmhRXjqwIydq+TFJwuEjGxX0EOm+WHnZog
L9388kYRCvlu5Ll3hozDuhSWuM7N8tLqLhPxCAdlQMUidG74cXgsehAKmo3+THud
Tlp3aRWSMm3ik9WCQICV4bwQKqNaNus2cwL6yVIL1aBodPn5WHWqMgF0MC2Ovqzh
BCRwn3cpQ6gV/WsIuRy59MrFCQOvVT69jl26ouAR/TVIPkXPEpIqFVciUOH2gsau
4oi7OwyEYWU66KYUzFwnBi9QDGMSb/u2fxIwFPHotGfKDQ0U2A8wPshefaVyjaHy
880K/YaJRNu6qhJKOJdtUzc4/NAW2r33SW8BV7ai4wo6xFU0r1lhomVqOlFM4r/G
7VAzTClS7e/CUvROe+ObdsGhOUhKFCh+8H7FPvWLsNnnOVi5vvHC3TmvIegYtG0f
37vXVe/uoldLRVmbJ3VD4czR8kudzviAOUGcZa6TpFX12wOjsqPer/0L3J+L8qsl
+71M3ejhIzujfihYDU+x4QGDDrx+lziwybQ6F482b5PjtL2mpH03cKjnxzpYrLJH
OOrP41OlEWoHutI5TdNdNwOvY0eJ1K3EeoRvgVDblxS2ixLyd/FdJ3xX11YQx84g
0i8kXFGTFxWVaKZtM28RQ0XeDJOs1SGr+yLE1VzRwgNril4NoGh2YeqcxsXtHZSb
9WFinYl0CI3zt7hCgPOeaJXXqfzRPs738ZQV6NUz1nVNrt2R+iYtSh6OmAVIZ04g
5tsV9lvhbLUMRkUb622cN0ypea4qnVHWyYnU2nyDrPZKRVr8U1DvIQxz4liE8eGJ
3T2MkpfgLkHCg/ywlzKVcrdP5hSOZ0lFlL2RUqHSkMft8Ls4sKNzEvFXawPSaJyH
WP3neTr1KC4wxgRa8FcCGUpWZv7tXi5cg1l+QTz0GJlXqzvHpg2Nz/oMoOurahqU
2uQGsxuK7ZL+ZT5+H9yKMIfLNvig3jJnzUc4V5edoncjv5b7YfYA80A1PvaUz1Ah
h+bFAMHwDJV8m04pDXA+uhUPcBX1iq/f8NSsYfs0j7ole48LUISzrO/ycXSZIkyI
dAomaIzwPHJFgCPmVBRDnzZt8yrMjpmCEicTPkMwiIbO4BwbXd+aD4uiEzRbWjIS
Gc/jIVz8HOm2KM1ZltiYVkO8ghLtKzdKKCmj8u4+fpcr+nrq3auoTuPl6Xg7sKZC
uYcJQRs3Ao4RsTD5Zxz9m/SIkTdY7PgGMFrCVXuGHRi5D385r3syEZgJXCPYTs1I
FZ60EQ+22UROXJpEIRSmEw6V0bIrny64u8SAULT9k9nbm/qZ/serEQeMbmQJ6Ca5
Wz9iXkdJwe34MUTwe9o4rMDpoe0AK+w+u6gB2movlqemjx2U+Z8+KcRZA5u2mBk5
Dxt+m0ELk/K/O2J2V7O+nCIIK0IbzFLtxhmrOLkxOgH8XpJUyXULKD9nJcBTSWDz
jivVHFh4J6sADz0qUdxxmI5bCCNvkrS25K/DZUyIvGxTZByedtVqcpP5Xafp+LV4
BhQM2gAkawEWq3cMGM7t5bFx0qzX10CjpLiz4syramv2v36wTYjwPx0PzqpvzBHd
5VPdfuRvP53eWLH3pKbNwc5sFY9KPngf9RKhxjvNHHhZdltnj8l4v7gC13hIIQs6
bBMHN+80jB+E5daUGWax0zo/Ro2eQfoSaOtscvf9xP9fOoeGClLs/Zt2L3yMWvVY
slQbiJMYxoBcGvkgWErYP2Pr/63KH8stUClVmUZ3CrF17eHfgfNcYzs7E8T/UhTt
/eetqG41I6UmWXbt4vPSjym8iwmn+Zgg6RAMuG37ZDRWiKIf9lHkuShkyTolgnHJ
UWn0bDUp/mhR9DjM6Pf0bLrStp6pdRssrTmYsWyAod/nEBdasxaIv3XKKABzYokx
SWmfhdt6hgXwTcrS/kgiWHIsZISZU0K7BXDh0R3f4J58u4lkdnnePCNoQZ1W59WO
cz81M/xJoMZZgmTqdgaUFmfXgRdT58yt04GWK9Moi1PIK/WfzZ8AQavP2RFNlsmf
wD/+gIqzK6B8z+aWrdPMFRGVDsxQng1a8t3tdCajp0fwPy0I14cnSDNna3C8pzox
wRJqY7HBb3w4ZqviLu4I8pUs1Jp1Z6YlRI4XA0+eU5DT5Yi84HPNOb9AGRqAV2Pm
TZC+Szr432jMftuqrrxUbo3COB44EC6bEFZ9A1UNBCUqBkrShRfisx5psMR+5rvr
kpm4kXzw1Un9PhR1lBVm6ldeJond329aG9zMDtxg5kkmm6F47aU6D0OmVm4gjT8+
gL+ZCbD6KJC2BGk/IRpoctEnVu+vg0XtrQSsAJP4LyUBQMNM8L8ohJGppFx8b3zb
JORDfuOujWxbk4BtAYPQaxPGCot8FL6YdBS8LQlRJIVEZkwCePvpd0/W1GCAo7uG
mfa1R/3eRRhiQw5KbUu5SaYqCLOsCMs1ZU1C9i9JdoED0cuUqa4zNaYHFWIjGSdc
LtLNm94cxpWROd6/+aliDi4SYe6HtJYQGbnHiDic+2PglEBcdwm7uG78yGn3IkVL
ad4kdFNnsTththt0W9NJhlvg+WbpI6NSumcCi74OdI15NGk3eyi0Ry8d4zvUi23b
LWlyCprLt1eFDtZ66gZa2J8Pyx6jYWkf3/uNFHlY/+dCdmu7jpHL/o/beT285cPu
JLZ4UuIsF83XPQVQN8EmrVCyjXbrqkMhu00q8zoaM3Qgtq4M0EI1zrwFq/6I9eFb
IzyycQMQQWBW2oe5YiFPtSbE5OFEKwaIdu1+BsEuYH798vaR3URwPlz4QzGyIFpX
688NnFCKKrlDzRxZcecwzkWAvBiF4J8VnL+gfGwv7Y/K/QBpJMcZ5jY4bsrrsCh1
I0WGQ0+2yyEFB+VuSpM5IZ5zn4p6O4WJXkb+Xyp6tFpHxGBJmpEVzHrJA+6pcj2p
RDzwBi2/auUEZ/58dZz3eatNzre1bvtpk5GLFmJFhPVJoVxc+5wOKX5LIZxc2veF
6Je/4l2AzHyKznCDbXdfmx9zTEcI4Jwj+CgFOfFrEpDUAWnj0V88eb82E+3Wnobf
D+tEd5fBEzwU/BGJGTX1Vwslv2HJslJe3l2tIB04Ab9xAnVwcBPw6iRKGPg/OcEk
eRwehm2XCn+ANo7xJ/3UqixBNjrMd0HD+B38/2uPLSghDfAzeoPzT+D3VDFSsJVq
xnpFNWGdBXm48QyUlI4+9pOSRnjFkLQ7ROdLE7fdWAlCWbvarP3AGr7yKLJeWow1
WzoG71PIszt6bnDDucJwZKM/8dYztypWhp8p0ksCZKnyX9GMxEpIiEr3DHYn2ZfV
YzNmjADM36rXccvadljVgdabrI5QFPGzqlqS7zJ9VIMkU8gT55O/MdCCf1vulr+v
Ui1eAJ0OKatTlzYD+amvVyzAXQzSuDKsgYwGKtdH7hCMMfyhysoNco6HVkJgly1N
SnUKgNuOHMeGDnywyUCKA/3x19Oi5xHMEWKiX3QTiu45Hr6RCEKYaj5Yefb4/4IG
AFD5K0F9mg5hp6lRJ1SDGxZMF44xWMCRf2cz/7wtUfRP4ZcLkr0Sv/YBD8VucePT
vUrqFxFs3XHlnDHZqHkPllFcdJUlY07RzchqcpR06HutJCfH22kcplupyO+Hbhy8
uWlEqQltHF3MlKRzJLg9BfjKYnYWq3uI4jFOPXd2oOKBRBTRcvF08E9RtuueKNwn
4ffmd42MdEh9FJgw4kop7QnHd6zAezJjouezDsIFCTX94hn3HYXFGn0+/soZ60fa
LUKtvOIwVbP3qPYY27DratqaR7BTAnc2IbQaYzyoOoTj/8YtS/lGl1zoc6a33jcF
HF6prkgznATf2zaGY0sYEXVxOPL+pBPTYfCPkyhufsqdIzHK8eFP8F3TYfUnJeLT
WTHYDiDQDh0F1/oPUEeY4sF1YRfun5WTQ/sXKVKmVgIsYV+iJWH4IK2LAKpL6/Xj
u4bix7HWXQpivfnJrzjguykHnWvK2ocbk3Iu3tIo9Mm6/KwdH7NX+cT7s9x8d5Cp
hJG5X0o2D15crY1HuiwbwOPohqy3fwbyE8kiO8qA3fbeQe2Oth2kMFQO1+nn6vDH
T+AaB/aaMSt6eQ2VjCMZgpJ6gCPfZFJwAK6WTDhOH4oHoxxSP5Mjtm3OMhT2rrQZ
R0FWo5wqJPVHwxZCrpl56buxis+2PihHr3KixdXn68s8/YQxkaMmr7ephV8W2mDa
93/bBUjQ0dte7I6IpSpcxkpy17hRETI7HFn1gb2J2VQMFib4DtgsvrY9hSthnRHw
VoiIvZqL15qYyboZlu9rYFa7sasBEzKbbnD38ggbbXcgeEWIH0UYjR8p1V0HmGXu
z7Ag0vS+2wy/oLRD1CG3RI/sa+sa4tXiJiwY5yzVtuxC/Saoe+aRIczX4upLNt0K
f0SGzeZJu0E3vHzoy7pTb4QOgo+FbcUbXg2RqX4aSs3QayWbs8UaulpQwZKeys/s
DXjHIrG3GJ7KQsYrjNGkHDFbbveataruOlVFjNXO/H6Rhuo12a99VC7+mcyT2QGO
8eSBpXkIViwNXqel70+yN3ocPxo463hhSwZMuJWjko7ltHaVP8spK+Q6BuCAAzsV
wkRA6llzm6bg7Vog6sTC0u6fvkVE7YsQLlr3UpQCecL0BBpX0X3D+EwDv1eLK392
XMCKmDRgCspBI1DGIsZ2SjnxSvrT124Jdlc7iOa6bYoOLSLOQlIySfpSEWBRB5OO
MvcJYDeS5AP3X585ZTCUB8p9A497lg760Y3K3/+H9r5nXohu4S2YaIpzlTVZB7ZE
UkyHOFeP/P2wasdPL3cY+Td8AuxY2nFAHfq8A281NT2eBRSqwHU36XPreYJJPMAD
OcmbdwO2zN8RKQlpnyZIYr9QWuDw5VUsOWtN5htIQAl8Jlt9cdRkBytFtJMOip/S
iCuocIvGYxvCbx17v2UYlWaq0g6nvT4GvXrkhJFehpX9AGIT1WpkOqVugI9MkuqQ
8AU0Gw8ofnVDJlmNtp2LsIgF0rkai3uGLCyx7lMiSokissWbSm7KRDex0kjSu1DE
B9ozZshQvHnZ7wp1QR2vH7lBLaHinzcEIyxsd/awHIjSSQeVA/p/Sr7oV5EaXXNH
SSbJ7wWRiCBoZveX375IshPxZwB+Wob7+hAvjJKnjb0SLn+6fYF9/lJ18k9+F2n9
ENZL4KmMsQYWaBDzaz4kgPMKf6zKOz+tQQyhOrlzqGrTSjnrtUYeVqa4NCIdGVta
DSQdTV9gfdRQbABIEqHHBgRA6l7JGPkv6Nw1r+0XDziFFIyv3q1rbFtfBVrwoxyg
MhL5UGuBhFfpJDf9c2RoMVqCySZLBA5LCBTqQI62OdGX0Gio6+EaGPkNTsMm0uPv
rXgCcVbacPJoGbozCUvOhpUmIv98ejaJ1/UJ6P7hGFYbTq21wWQCPBDcFaXxp54a
GmqmddDqUFuq80AGVyLl9Fjza3JcKjAxkrz0WFRVRBSso+u0iqJLI69SukljVy0C
skV5lEl2ZETn9tgw0ebi+9fEZ5QShVUcJJ/msiCZ4XfiHcRId8glo5leQGZY6R5+
saLv3y0gyTf16rNprbGTDfiYlprPN9JzamUuF4APOV3nsNVKSdNKacPZI5Iv7LHm
lLo1Kp2VjtB69HpCEpdqXXBv4VCWrvXhZvWJBcW8HU6sLRkalTFixo6jOvgKOQDw
xFKfDZhPjgcs1HH4C9eBpfvCa2FUoKKhDF1D8rmbGU3optteQ/x+VM6yaHuTd5JV
KP2WU+TwzQjYR6TxidQCLAMT0b9Ed8sCJi8OcjTrCLbqRwGBIi5537Pzz5Zq2cFX
elCFpNVmLvAf4KzY6VOGwDDk84+s5XH33V140cUPfyP0TFC6RJ1FlMKpK/RuQaeC
LbpptSX9QWbKNqxaG8TGWMCuxbnawGBjMhRt/UE5r+WMcjTcmIJ/3fafM4ZFcjCD
WaOxj77muiviV/7rwRzDjfq4r9hOKmsggHAllyIomiqtad1nONvlCxUkLgKKoa2x
hJ5tK/FDnMy+shuL2giwDf+L7gIyqRyOjkAlMPxvOsgSeCsw66iR1LWMFdlAJUWi
G523CC8o9wyhjUjyveIJ+h/rpie3PWI7Q89fXwg2XYLvE7tOYPrmSAGUB58RYcS0
/xmccRHGHGhL8CLqcbml19TtcvG8Vcf/nDoi9luKb3vgZma4276VcCU0DCld96e9
LScRNK0YOIpMqtDQaBJiIkqPdauTyTBWLn8eO6jWmU6Kd2HYtdomn5iFKbA/HfF9
zF6CGcfU3LODms+23Z6zzFQaCIMS3CQkpjcfDRA8hs0CcPLc4YLK5kuiiI8OR3vz
MjJrIoJIVY7MD3fHYJkeKRb87ejqUGzpb0xPEace7dxAEqv/PcB8UKOSKKQ/duvr
jHXi9dY5yuFgAxoPxqP6c7gqLmcw8iheHB6V9nqEgPz92FkPibRst5v/Zgwgx8bq
kwVwQnaQ+jA5XDJP2G2AwEbWiL22f/ErkYeWAGd25cqvoJfoL8KsIAulWq4TOaE6
xCj+Ks3/YVFeyUw0pAlhOfc7ps4tzmcRfJ0PftDi5J19oQ84KWWwlaTzLVDFLt2h
us6199iI96U8lqrA23RlC+MWckko1aDiW625O7Ft6XO3JSpmu+zlMmEWtkv6rrJO
soRxNkEj/IqEomC1AF5XPk0E9Qj1Ob3w0LjJqpjBiI24imWIcvBMBnvEbhfWSDtJ
MfcXlCxsgWjR5Fw7lEwClwNxwwO3IfxmIp4LCgkfQcrAzrAlU8940B9RMSD0p2lj
Xh/vbttn2vNcjxV0PH3Ha+ri/iP4rqc56CWc+HSLVcbJhooOUpDAPD+TY9WHkXyN
ocAt146Bqb9LnVS9m1gfy5eXuZysJv3uTCavzLCYcNAA8rKvblJXdQuxnLDE0+zf
3zX4EP7/K6GZdidoaHyIrzS8G6uwIAwzpAk6Imy0h3IDN3W1ap2Y6AyBB2buqJBA
TJ3Y89Pu8EcJQoRA5hV1VzVJBaHImM1iKtiZo3q6lkyDJxwM7uBDAaaoRzqK8IG1
hCn3Ajavk+PLR1TxBN+MpXwBPYTPiafnSJ0aXRn2ZWFbpQgoGPFdEYELDe2PynR7
ZcHbarcxd67UDU5TH7gobBQPN3Zv97LiNnObuFRnePHjfAtIzEsoE1F+u8vjSUET
TRMY1H2Dap4dklrywwtdAMtnW4137dra4sVlBezgLU4oyVG+xuL4hF6Arls4jLk+
qJZbR6sCxZp8bH/6WwYOVm8PvBsX+xpBpmqee3pr1ieIykU86QQmuojFT5SPYlIW
jSRF4Ems6RtyGBHvobrhqYF1Lzgs2OvZEob9kBITI3bm2iZ8iBUyJ3x0g0zUPhD2
ZWIGviOvtaOJPbZmU7Swgi6jtbFCIXODXKh74Amm9MCrpIA+yKtM5odc9J9kNVTY
xXrIVNAS8YTPv2a7Jo/BRWGpmi1cGb8bY2BjvgLxspz7ajf9At1yHiAy7rZO7YDJ
/S3ua51ypaBHBIDnW4fbxXAsXK3g1ulESmrX7Kn7xZd77afqRmkDylHLnNgKp4bh
QlUVCSZ52CetS6uChdZXPnt8wbA8MczgOQ2SUlueLPB6DHl06cuq9hpLO9MtGAVt
IbvqChne7uc+c8w6KyYNggS8ZtehDWW10qJ6InKeodnaeF3m/GI05MTSgWKX0veF
RDfO939zWTArH2ifb0W2UJuFss3xE8CFyEIBebxyV++OgI0j3ZTmCgJbt4Lbtn+7
CLBalmJHybiJxO574cJiL0KFOnRkMB4JCdNBUxQVCZ6v3clE/UvaILlDigA7Da4h
MTLLToGGKhvL5xMcB+x/TcgNlsO5lABjxbEjSrGNbZC8IoXujRTyDAV18L5c4nsp
H+yEJ0p0ArPiaIPxo87gm/f085kNy8pFoOfzSRL2OEWJ81vghYD2uMLq41MAuBXN
WssA1sH4g0JxOb4dbv9Tb6nkaPpopNrS0vnctKQh/lA2K24RChrDRoDXTGD1q9Yf
8do4+6bwnY/etB0kcr4Qtn83xHzyLtbbPlEopn30Ss+oeFW7o8CGsG4jRdEIZJ0M
wYj3OHaWbpnf9pEbY4/JsMn78k6hbtJLVuWUwSd48Zboz1gWNduvaAjIpEAaz9Lo
J+r5C/aZJRab9nCkkPRMeZZFn+do3IZsX+pjL3/wbyTxwRlVc4VlbigF7sUJlWE6
vSlF0qB98JD2JpL71dXClmrdLe83GNwunBJUzEzjSOAgazmqKIeGF5UtdqG02Foc
EAuhSwZkTZlEmbdqLuvmj3f7L3X84AJaV9KRFpS6BCc6jvPYixwKudtUnWJmEGPj
yQb29zYFjYzdB4dOfKM9Ezkgw0GSSOwahYPADO3o+BKKfIZ6x3Velit6qpb9hOVt
vkPlWRaZjg8whV7GLBGzpAj99YAQYE9XP1RbS45OX84KzrHUvW3qs2CSZuArXZQE
njtyiiqbvreV4VVxc9xeqdS/bLjVK+kYFPCMQ53Vv2Q84yduqtzDbmfb5Zpdqt3k
ezbO1V75NHYvuWc2b326s9QQDnI3BoFoJFtDrrIZZ73l7htKOtdyQlo3EJ81dqpS
EBrLPa64WMMZUg/V8cYwVBARWWdNXMyJOhLDWZAhW+C/kIt3hh7UXIzj9tVggK5u
rPKin7LpvLcTbG4n+DwaKTr28NlQSYCbDGDIi69yZMXXHmek5RKIQYlSfg3nO1C1
CIsBEiN7UCkO2V0SDCFy1IMSO05HaXeKxNI81U7OLDe8+sRqcfJqmU/PP7eFvfSs
0I9uHNc8jqw5KhVRRfhVp7Myy3T9CJWnVKENdlY7c1tevYCRxvYhV+Sa1qn1NE31
1WS6/9n29OQO6js5vPU6yqklmCRhcGaI3tgw+UAlJ2CuRfhkRFpgmiyjL3SM/N34
fZj75L9AVJquk4sJVFCt2jvqRJhbE75MABC9sF78aM895pMYkUMz8voJc5kVId5b
MAL8vyBj3Hf7IS47HUovBFPFVXIdo8mpiPu/NNVUx5UanxI4FtBbLCy8YC5wYdBA
1kB+zOEbNnAu+AowdoDUweF5Jp05CmQ2LylJgt7IgiWuqsWRD89yVmlU1QP7usvg
tkAQLzeX3jh2gbgj9Onn4Vsgc1uhM6yhtNYzpDYsBht5NHl/5WPysA5oyTtvsawu
L24inA3f/TqWQ/kR6dTtVeDKJkPcRJLe8HxNqufxe4XaUJgjEE4+noJIW6I0mkME
WrMcyjHfl1+7M31kfHb/4BivVF26Lzv7JfLz6YsRxHBY8XxJblyW7ix1JCM+8spS
l/rkBOaEhpi349Bs41flK/XoBEk61yEW+vTF23TozRSjsq6jU//xrWm3M+WI8VVZ
NNGy+3IcBZ9RsOMR84OfIZB8wEWY+JSebadzuYMDosoPExXLorlhsxukAnylnYUo
tpXaGoZLgzmOEdckwrtj5+ng3ZEnUoIIGRK6jidRu3+UYsOUU1mSB56S4h2YCOmB
KQ/dbiF4rCMNqKItFk+F9/gCngymrGzppfP+cAJiAQx7qunUOZYXdNOMogX7iGCx
FRg9kTdEOu+9paN08CyeRwFhqrmKYCP/IoXqY2cJ84n8yWUWS5wOUlKjteNlaAR5
LDCO/Ied8Rz2WBoE0k9J1V0Cu0/pPI0CCSrLgAwXYkLoH3k2zoMpHmZANM2WAlyc
P+U/CYcUBOy5n/5oGl5KFHJbPWI5NMxjSx/n1jaNJ5gZPE031nb0pCLbE4dCXKEf
GdvrWZl2BTriYij8CcBfJ85D05EW5MLrTDZGgD8bhf+2X1iBGt3fyBMa0QsTbLF5
c21YckZpQ80jD4l3jOs4mKsVwveoBWsksLlyn5gJcuESZ3XpUPuSju8/LgihpiCv
4Mn+1yC72vISbPnlDbvH3eond96gK+EcUbJP696+1GElUOQc4fZO01mgavCpI3EL
vhTt9BWsNUAa3FL6Q0Yvae//gwbPWKilLsquitSbtSiC/NFrj3LAOGXwehIF8E2T
XD0sFf+6OFMWhoj8q+tAH7WQa82pwf9+999XUibzWA67jatU1DMMFIx7t+Z2lnMk
YvGP19+BVRqOxzg+2oWdY7wz0a7n+sRsyo4J0HR1x4nH8QotFkGi4yGnqUnw1faq
UK50A1KuYZlEsb0SNSlGVX//NLS8Liz8GPmmStbZOM/zb2lKmpIlses0OVNtOZk0
QIrLdB6ypX420CiHsxVgviHDCdKYe4zDa8xglRBKuBNljQlG/KYdLk2h9F0Bp6R9
XvLGCMjoG1zmWzmxvT0mWh+Uv+WGm1QOH32S5EZY+/l1Jq347QCds6Tw3SaWfJnb
FZnYTPTFaF/Pz7Zaa8b09RDNGgDToC9MtYvNaJECZ7b1sdD4TMFRQpiRXcukqm+y
sRAfDs/j5Z16mWXS2tZd+lXGg3o37aI5kSO+lFx9NiAn74ZVNdhdFflFsInOytCJ
jbydHFYAwIMRhseR9utyIZwkPVbVMh6XcZUt+FmoH4Zcx1rwz8DB7zhgiJYsMZp7
9IkrnDwFhh73/qmDnpQReLUINpfGFycu4qD1rt2a9SWvyFyQYduPBHSbJsR7+Ntk
4u6fg9wgLQ5s3rOmWOmR0gw20QuU/M38LRgV37oOaq8zymk4npueoL+zt9aFisFg
tTIoS+16DqnDvzrdscEcB3b+0c/8FqryjwbEQhM73vtE1+La+ubZhO7vdbM+3S32
n8OsnPxRjOzfLnuBBGYEVTAm8QqHqCuINOPmgcjacmlXyvdU9amYosJ0dJH1vwgu
Bz6gRLcfBsxNTtzqcqn4V3vQE4OcwB+xSVIHYyi9wk9gIMj2cf082EW9XAmV2394
+sar+3btj2vs6dy8jakTW2Ql7f0qaJK9d8vQjVPhWVFnThBr+Rbjs7aFVCBNAsUw
ubbPsi8NZiIfHdanxU0tnyhzg56WpeYoe3XiMp2aHTHEg/renpH3KHXL389mLitl
RfhNvL8V5XbgyNU0PEv9xAjuF7axYCjD/Rxlv7rCKmxhvPud64vfrUA6vBBu8q30
r0ekAfn2R1uH344M5hVSbFtTu1PQeaiOVl8BcGo8xhH2sJmjZ2oUNLAYEKymgBOG
Tu7sMF25QKPuzRUQOfud7HbTqSRNcng6ep599HwXdyOtzssfaPCiyq7U34Ub51vU
wMnjR+f45nVBzGNzeIOpeFv0nb2xnTqfT4RWyvWUtH6FdywekOANX7dSjMU1rCQH
RJ0cZqjR4G5bErelb6lecRyDVStLJNnQeoj9PDES6JiDPadrvXkCvNlcsRp3dnGC
MsZBlJpCCfh+wpq9As7PJW+khm6ScIEDmfflRclUto59iVOF6m51ZsnqYcnL2i7u
oZdad37Ybh6fGPEs5e90OxmaV1mG0pNfTJfqCh/Pzf9ZRLRypgTFIajVYoUjK4mY
xsGcW8xAUqnMrEWVn+fZfi6/xM/K8WmTPHHtd8uXhQrrjZokeml4PrP51wS0v9yF
YLwWYOVm5Yku/wV/y6l8ANUBTMoNw8CDHqXkmvUcjzMJnYXiYxMgEFVo8BwsNl56
gL/CwiG+YAPmuD399H7GkPa1v7kLF9LJ2SN10HSdOWTu6EalIj/T6YcmA6uQ5UNa
3pJOV9yKbcAMFy3GVgS7++f3iXpKBKeo58c+ebgNbHNXKGHXyCGAssuQ+ymHT+eP
54LM6fJR4mxd/eIVYELEEmgswhtpobw/2SsC2T3+Hfyqj8rkE4A1+AHAyBN38xWD
Zj9d5Fr+QWkS6LDGa86tt0HcQZwkFzaCE6RyO8iExaxstbnbTaZWv+OdTga4pV/K
4MzApVNHa/7mwOeMwjafUIlb7nznz2pHDbv3EsB+ugI7i5hvKcJn/Twy4hZ03XpO
gCYBo94EmclxjwdS/a5QXBwR6Sp+LOSZTrgLuMRrHsAnt/RooymhFLEWkV/ZXJc+
SCD3xV9RicDS4Z+bgC9MhoQ4kTVE6CNKdGZMQSXxCYhQNmIotNv6cYIj0CPQQvcL
orc/ddPtqC0OUR/miDbJfymzjzxmAgXGpu9wPEwasSoZvD9eih23GXj/85qogNoj
CJ1AJ0UbYh6KmdzNAjfQXNwt3FcUSQq2kh5VKttobG4s/0M5ScLddFGfC52dmPoA
fF4bfJnmmEx1vThazWniWggnLvrJ0rhWvxKUk7bbaeik9N2jPByDM1iO1ZMjhG4Q
wI18Vtp8km+TgNyuTQyoNtABNV2FnOwRNU/KM0aEE9TIWPdq/kWOeuaiT3BDIT6m
ISo72OB/1jO0ZBMxjNheS/HwwX2HPCtt7VvQp1OqP5xMwPhi6khNGTbiTlguXcio
aSKN42bIJGPY3rEOSNoQz6tQg3zx4Xp6vI7YDcSsshgjVSptWR3wbhesOpXpPDzM
VbGaWCWAuHXeaQ9FdAtBJ25f3TrtDoUFVSNk2ZOSDJnLSRM5QkDqQs8potaKEKYe
wI6r05w7kgKgt7tXAS3zEvnieGPprfHOIH293ZDM1alcaKS6VXIlKFcdqtePrz8m
ezzx6D1hnxOuQ5YRL3uxCJkTCsS/hFquhGEvqFytSfebqydshJnmTcoa7MNSBWPQ
/MNlx4XHQ1f80H8/kOdS8iP7uN82sGZG+K4Di5tDfEuhmnG38N2KOSynzV9ygpXa
EeEujpctP29rjoY28I5OA3RdiP4B1IiT4nSrqekObt287IU/vR2Ts3EegKWD5rS1
Ovw2clbbal7JebRmYdi5H8iJ9xYtIS9GDnku3uWvCJiKL1cC8O054GN3bC5pKNiY
tDFVI8PgyRe0BEPvkmpDXGxaVarH9K0vEnt7eYXwyaalP7AfO/pJOhDKfw1fZEHV
ydcEuAQMdqxDa26ipSZbkpDRg4TcQ5QFXUQS09bpyJFyU25hmmFZpOAIXcj5dDjc
UsFtlh98ze96N0fptJLeUnSat6mb0xn/iiClZ8KoTKLv3okY48ALU5tRCz5YVo02
E2RqkOUriHXBx/ws/x+/VTfn9jJk5MkEzkI72NZBWtI8GwvRIUjvFqpyNOnEbxtS
r8l3rDgmtvhnp9LRCkvIfJ8GbTsxf1xwTHSVSeG/lvoOWwVaRlWcKElWOZPH+sU7
sNpZA39YIUNE7m1gJwvqgNk3jWkRiarNnDLSg2Owl/pIHTLLoZoJRABlwMSkg6xk
q6D9XcQqzf0r3c+fphOOEIwVOSeDZegWJjRBJ2UUEWgWbLJSHF3G9GYkdgOVOQO0
3hk9kQV8pT/E0FETqjYbKkvzd7PEKE4twIRUqkSKVlaXoDE9TAFoTPichu+U22KS
HBB5CJvyIFJD1hnCEVzBGImAUaxiZLwln+QHwNyNWLQ5BPmrn2TCDcUDC7z8Fh4+
z3dRK5rA8l+clIuTdkzGbBmErlbFVUnYIB0Liv1YQU0ijKXZPTNotddJOdEAxv+p
tao5IIpupDlT45Aj2pmqbfQrJVgpHSK7fh3iUh6jdGoDCb5t6NVM5BKb3ODt/Ta1
dRmDcO4dH5hM0ULFG1qT3EwWFvHIiQXvRatILzxDXnk8SiZdoGgrHk+kPRDUO2cQ
Qq9YPAePEHPBWs4fHxq6ZNwAMrksYvK/ex5XHINEFzDr8eLpjBi5QqkSMkvAyJoC
nI/wmml5PeI8v7Jg/vmX3BpnBVzAwi2h2RTFyaSKlqgVOOVe4wSW+VKobRZpOkgF
6Yy3PEgI/3GzjMyNgTD5lYsqcFAUnsomPFKlOMekBG2U2/teZ9ChZnr+aKMhTqR3
ncvUDR92OeRcHLYfiFOuzO1LfISYxr97CMzUuoBGNgxo4yi7YlXAJmocpG//AALM
OR5j4dvSD+iB/7BcGG5ykczDpcvc8Fdjjpzmvo10rFZSEK/Euj7ae1EJ93QXflaR
JYzcXc0uGOp2sXDaBEyCf9ltoMBO9cNmpKCjIRxEWHWQzMC+h8mRXWjwuiydVpTi
cIG6jIZupe14DBX1qG8cqLseZCj+ILxEgFrq3X5ecUeuWggozPnP4O03qNLwCtaY
M7TG5PN2zm7hGBzQUdJCRvGy9vPplUN3IEhQsHSaMZQYe728Nf0RZVEYKwY1jANV
EyBmSZV7HS3jTojvpaDEMZbBxgopOppiIIG4NDUpgNagRp+l+yxI5emSmxAm5HNo
hQllbbHN3eoOc/XUjR8QyCay0CsUw0nd08Ofj/coXmvNvAiYZK3NMa648FgXEr6V
rvoMqG0g0/n0beF4XI6atjEeFSz3QhFonSWUczUSQXUbKx0w0FUQnOSDfO6QJphj
ZKvlf6e25qQDe5uL7BlfbFpMOjtUz8b2IcvfAyPAs4livYxNh98QJ34XgkUQapMD
VqcKGHiLQizWB0ymYnGBhXK9vYp59P74tLHc04/YLnbe3aidDozzp7FpmpcUFOgm
2b70y3J/TqlI9Wn/NvvKZCLdyYMeoUjt5SWIms2IMJO8nxrdIXCj0JTco/xxngSO
nakNxkl1c78Lor1fCork4Zy8/FMcTB8laKgnmTdSwaXe08A3jqPMug/dgEvTahd0
gE2ADfo3xlkUWCw572mSRV2+EOtJ2l09IFNBGPl/ac7OCS4k5Cc+/WNGaw/nTWzl
O1gKZ+a5oekG1PZ6Qm3LzinvY6nnLCGV+8CW9r42EZ/RY08VLueVirgiwHS+ddah
dv9C866SXbJkYdfLbUqWv+pprdXZEzWJXXPGQj1kZOvG0f7Q3IQZXTLf+qK4OyGW
l+NWI6wystdBe7QntAWiLW1npf4iSawK0gFFcyg8YoOjOcOrpAJg5Bnskrno8vle
0XiTHYoFsx0mjG1ZSdXOvKKu/4dudyYvZcN7gXm9Wpyn2ZdTiRaYFO8qVCcXL4+a
4PdB+EvGU+EOvV9bkUEqVUl6edg8cjZHFsgxPHz0xrMR/Xh2SzxNCWGlPztjD2xa
FbRRSybzgXSpI7xM7sYQ7doSNgDuGcNtSkj/2Bo8x4PA0R0IoVyiUbRWtJuXW25X
rUCRSE4lSDIz/wqxCJ849mue2aoRAGOpBPsH2J7Mhzq0+sAVZTz2HiwugiYE6LsM
6FNV49F/0jEAMJgIXh9MyQaRQ7atxmB+M3QLaoVZN99Y4LRXqFZfX/qdomxdpig2
PnXNm7yFIxpWcseyeYWvNlomtnZQSJg/q3gJTTFu/B/k2w4vAPd3hkP0y1aupfmM
nN7jbRFMAe/+93vElYAj42Z/ldB1xT9XvgDAaciUwnNp3oXUCzZzReIrjaXl1gRl
N5J6o9ENInezcQ6Dyq0/nPIjOv1ol0vi3AQTsPgyUWL1KwjvlljFdsySD2zwESzj
I7XazihBJM0Fn+F71oFg9omQ15xQUsMS8FiV+E7I8JzLZtU/qHEG9D36qibw/jOq
bzbO5l7I7sblGjqrHPu1rp9jTqbhJPqEMi7IfrAZ3y5wS4+xIS8FBuDLI0qopT1H
dplVZ44SqGC5Ehe7WSJqMOQpKml/UCSDn+9Yjy8L7zfNcF4qFW3QQXkv2g9O2tnK
u5SHM6WqkVLieNI1cwKJa/sYMK+/Iy3Y09SfvxRvYvIi9YgYXIGnbkW9OqqhBNzE
eAWdVCOS+1By57/j37Gwg33TjXf2NX5+U0k3XTj/ZYlDuTkFtymSt+cwHtZGnFIt
a+2JlWuVNEzcb/AQNNs1kcf7HVpAAkDVnUZNmLIZVjkcLN1j8YKVIPHde8ldpxxL
qTwRV5v8VzWIu09xKxTJmiMBI8ho6+BliNM+EYVX7RXHq541IUw8r3yT/OuYcISd
TYXp9vgtFFn05n9Os7PXh4V9Ax9XTwWqww5pw0GHhXDRTDEt/NnqzZD9bup9FVjJ
eUV8hWAEJriKbOEzJbbM0TikhSC23F1ckRkHA80ixdDbYqd25xp4t7pufJwOH9WQ
CILqLu/eAD72BM7lPZCL/x0rpeX7IwEBYVymHLF/5kxPcesk09ru35Ot71oXCR4V
u2dYe/noNbwAoXQ3tJdged+fEPN2+4ESkjkIWaF0Avu06smsLEP4bLlnC/+UCp8j
+/w72Jlfgg8+KdwfIffRLypPcY+/6H1vNGU0AY7XEY2Hy0n1BJBBqcEcg9T0Av3G
7TH5TlncvcueG40bFVSP9LiyvpLQyTYT3kPqun76wtjhxQeTl9KudHbXMcu+0Tbs
VshB+yIjSelslwF4RmtgwfV+aZ1iXtL5/X11qLmup1S+Tt4fufJ+4kvEy1NRhrDi
ZF7PwztYqWldbBGlNw3XpTqmn4gF1dLCQwisyhawG9Di4KhMMqZq13Czw9/ue56h
ICQNOQFz2BpZzzTIS+A8JIApKwmUv9yOrgIMSZs1m0j/U+9Q4jcunqqM1XPRgTJH
0rvmj2EBe3Q36K2uXBjK/OwrF/4HccpcHr2PH6mBRjnpSYeyiun9vgFLCwUXTqDY
6v0c31oJwnhaAT8PvLLazShZ3xnWyw7hqttGfSMtRa8IGvKwP8T0bJQKXGI+0B8U
I3NGd8hHWBKzA/s4cyesU/PRrzREa5L/alXYA0cCL9OlZSuf6bj9e+Z/LVKC0bw4
k1TK2p5jVWCNa9pjp+G9QDc5RHEApUJ9qiI7dI2xOu2rJ58vK7me3NpVNx42XMNs
X1ADCZHWmuEYSG9vq0OUdCRaFT8df3crtmPhvgPgywuPJfQ9V7PM4DHavgEg+rzU
JVZMkkpbiSSSb0jBkjL+n3cgQhCZltfNdZObIJafirlw9Gnja2Umr8vjqjz7YWS5
sSHeWuoNW/SjfOqJWnhR3qux4FhIIVKE16CAPU/3gxgWCF2bhJ5CcGNHtyeStRlt
Kh7QsxpLhNvrd4WMmcreoOZtbHMW1/GI2Nh7yDxO1oPtOmjehknPZmIs44Iborx4
NZ15GE/jqETbv9zuneDWoADFKw/+g4pRHJximNVFlO8+A5JcTyE60MsmlyzqS8Jy
YnimSxFIGE1UybLR4FGtuxYzSkRplYJG4M8V2TrA9goLc9JYLDSc6nok/i9Orguw
HyImaWXe1t4QFKv4F6t5ZiNW/9MWFJKMFUaWBHdZHE/DsdSbxBEPMte1hABcXUwM
Io//oYvBNb3KbG411CdxCr8MXYHP45VXYo0rE/VboxSKsQdgvb8GHFjh+Py2297Y
IClWOIRWYzlLYxV51fI9dEgrExn0qMqa5PSSpOjhIiSgKaCNdvxqQqK3uHEeOHAQ
6ed/U778SWr7jM/phD+feWqBByiBI/2OjhFyqAcULWJ188rEw/Mz3QMT3rEU6ukG
/3C+xSAkLFFOJ2DAgrPbzqI+hAyiOYOw832Gzm3WmzZBxC1bLFKNPNe+3DhZpX2D
9dcjXQNWmC2t5uS4/KJzozFgpzdSo/hwsRuqb1XTYO5QzV7qIuWOUdaa/RbzOBXf
idzvKrrqHZjs4WulPA74QTSAmZsTLuvnDdgLs7l3ibpnExPHhnFxj6YmjCANnS3s
dGkWhBXKkhL5qJsS9U7ib1AJeEH3h/Okg1Waa6ByzqUZ9tbPgCR8GDQO/2DVLTq5
hIGvqoYpM+h+U8b9ffk9rJwWw6WCgb3S3cw0qecdguarrKRl/BJMF+TkY0+brflK
F/e/PxzjvDP3oMAE2gV+AQ4q/lb9bU/t7sAR1i9O/lDCn2HIfvnafYVDq0BfMfaL
5rLddwPt8rg1okOXKC0xjmJqP6fGK8oVKGlczLQ34HAjPJ8kVCfhKqoM0ZORWnsk
FIsdxiknO8Ah5NyqxUfZtWpU4pTzp+wNL9oyVTdFrT89J1/20yjIcJGZolLrj1iV
1WG/rBVSRwHA2RhtzhbDf8BM75oZURJ9FR6CAefnPEOco0tKfoZoJVPC46DMBdFt
ZbCjtM7QdWQIDaKLgi5EUFky2rEgbmynnFhQPE04qIStSkgWyM8o07Oc72Djxpiy
1mYoCfoU1pmCAiimM2ZPsWJdxg3YW6HR3NLBz/VPoeMjLpnn0yyK4SjNn6Bg1X9a
Xrfs+A7bk61wonFI91Oyj/yTaEF1/KlIzolWAowegraVDxZ8GPXxl0kDakNe3OWC
82L+b3mvZ6nLzqwrweIP12evQW6L4nqDAjn828Z4p7o9RmFqE9kpcjZ1sTXs4tY3
RSYdElfNYKK5YvrthuRHwrc8ShLzpE3574M9CrfFRNPyu1AESpNwEBA8veFXYSGp
ZaNZxMhJfrNDsXXopH7q5f3jwDja8mIokxkyECp033fwqowQgsSQ6UyoUU+clpRM
q61rGKvczZseH3hNRlMOSm1H6wGeVj/ZGuYl5hEWC0Meyg5o9MSCysIP+BA7Ypgd
ZoojVoEzckvQi0GuSohzADzE9DGksaH4zaJPRViWyiFZmuQWsiiBfM084rU49iu5
csTxufaPmJxtHcn35K/2Swz0Uszz6WERVuFTG5NEl4pxATcFDJiQF9J74l8CvYYq
1e6kOpCyU6Q4mo29XqiBqwvf+ZYgemaZCue93nyw6c1dBye4oZBDGaDDa/2DiuXV
QKQd2VK0cbvQ+rO3obD/grX3cvqzAol0Aa4GANkSnix/bWbm6FL/aSULgzEIYF8/
CwSRulKCgU5qP6sur0PTAqa0fTbOglFNDJgJiMl6J7Fqzo4EJ1tXE78/+LMH8qSe
GRHNNSoe5Ws4fFArWJHAgE5bzThndKE7Py/ADwWGzypG0SgpVhtFSMtw7U39sg2Z
+9WviWqYVHSpQfarZsUwf5z26fSYr9NAw5k57hzpCI2R3c4IN368SdymuIk1V1xD
mN3dhht+gj/eM3hscuoGloYxSPoCjZbhrNv106B5nHPDumeLHNT32m2XeRjXf880
wisonigJVbkLHaCh3EG3GrODNA1rNnj5wQqh22o7MoTsy2+MmyhJk2RQSGKii0hC
ptwHBBJtOU/R0GEIvtMZAucNLJazLTL9EhaG+AHyv8UTBt0YI3hHNWORF5MlW6Pw
qmkJKYjdkgqQhD2lCQsZjnHm2ttMSbIQ611jcguFEASxtcDHtkRyWod4nrPYtOAg
yX/A0v1uZbisQvXmOWJktQpd+n9Vixq2jmPyzWZl4W6059lOaKiBnPsUxjust5o1
QgA5fY9vFmm70BvzPg4c1+T1gDs+nx3FaFJiwc92Tm97WPrBpTUOSM4kUm49NSjC
Fb5opXFH8jXOEZYZPANlXA23Mboyt0FNe+jOTIWWE7+uGZyAUxsenuWrr2QvcyOS
7ZgDOTiB5efhEt72bXWHxb7a0NcJ+4w2hikg3khTPoAfat/ANLm+PijNLDhxiA5W
zy4Ikyl2nB/du7DJai04iLmDvI1B3PvA/nORJ/BIlKDVA3fVTtIunpnkEedF0EKU
x9KJNq/P82IEjBxJvd2PEJWfc56JjUGiJK4LUV2tDb/ot4LOQSRp9iTENePsL3qc
g/pkIuJhGTS82mXhgCuQiLgjqqCeXo3nGEJ9gHGdttG5HFhAKSp4rx5ge0U8GpT0
MxkMEvViIOuhNUL9p5zcsn4p2aIxf8p8Pw0SJyAn8DPzUCjzWZJO5kzI8dKhv7SK
imlRQuk19/sSObqSRqSqhmKLYNuG3M0gyrfl5yhb22QEtfbSu0WdQvIPE0KLq5eG
ryBTmA/HKX0FIpVXPb1uDfSZoju+44Rk0IOLWjTzqULRUF+x7t4gRGIWRgW9ubx2
AjVC437NPsHnIO/O2HQQz7xQb9F6RKiTeAekcjR2sh4d8QKBzII142RiKslaQBDi
Rvipz1z6FRheigiFXCXpmzNPJw9gnuQaFILFIfP+XVS4hJz754OOqqrQK4RkE64A
xg6XP4H2Zvy0GJ39WAI49H1UrS2M9bDjUwA37QOI/ETFCP2Mi3WJjfQR+rdb6ZTa
epqkxr0/V78/xnVvr++4Ux19qP0yh0mBj0rU7edlqhCnus8q2kbg50NyjzO2cGRw
TpOPMeg3n6QKpGw8h6Vk+kwBU+xfylSqe3wxHCgVY3Md6ceCiGIYc39vX2b1+LJg
L6BrIMdJV6DtDusOyFTLlMPLQc5TwbT6X3XvdHzkF3j6esVmpoeGprXNewX098d7
zsCDw+IOKXZaXwGujHS26sRH0LbvIozEmmqe351v1QBGW0ru3Uh0wIOjDLox0shj
h3GgbJssqIDpBtQyIgbDZ9jP4u9rBCH51dbnJlQEKn97l0rF4ia09QxFkr6z9U/q
9/2zBB1xH9k/2/tv6KXgrq5naoVMDWoJGulG9B9oKZE8s8jYyfZbXnDOusWVHZZf
/eQfEorZt3/QDwijkhK4LFiqZydubA47/MhrnHlz5GS2nmzlqmAk4K4W3rdX7ALe
//Mg7zcD468ynkxaDOnPSE1Fb0ZdUFzTiPwe+urIN+cl+izrHgVbrW3gWPig8KBH
fnMF6shioZcY1MmrelreT3YzKmFI8ddEDv9RYsLBuA9ITAof2mFI/Nz2bf+Fgb/s
3pyKgJcxTa2ywY3hIGHvSjCPvXIYfrdMLnMSl4G5Mi/umrDmBs4+LEyu6MDk9ao6
ENTI7oaW+9kdmX9+TkXWaZBXr6F8f358MIdv9IRRz9cZpMcU93s9ZHEMKfO868lS
cnS8gK0+ZFKL3zWiRDe64sP08y/R9OyHkbMESaqrfd4GimIesYzy4pYUvxcz0zwT
JlxOS5NXOww0M85ZjoNHqT3HF+5YLMCU17FHOamfVt096R2AWTUQqIeGVICcLNQD
e8Ir77Zoj7b4koPdCc2hkdI13b5ivuMO5uFCSk2dNRphvAFRr0FMnZCuHZOGZ+kV
NZ8hHWyLNC95Q4m/fpVmOdp3oyDendgzSjuuJz92TFuZCDQLeiM/ojf+6u5k5ugU
kkTDv/pirzRaw43JM6W7fHgeqtFMgvNjPCQzEnzaO6ivnBH2DDhwYYKii/FmCFtd
jG0YpPNTKpLzw2o5Nyvy7ASGr2HND4uSOgYRoJlGgKn9be8X58SSRS4iSGIbW1U9
BFOO2ZiNIYdPVOxdeclipyDpMI7hhVbWW+7OLX1rLYdnmFiuLMnEbPze4qySKm8x
RJDGkFA75T5icjLKaPKZt5hyxBDrwneuA563D+mEtxSFHf3lGNCjX4zQDglRZSQT
x9WpeltdxIKEMDNJFTOyjlZjKgYFCuySB6rMoruczqoF/14FQQmLFf1gehxxy7UC
eTbO6nC6UARCgR6QN92S1PxmZ7N9lhyn4NuGlLMiT1d7HAuYQCQi3AKxTCO0T2A3
WT12deqt3CreaMYislyfOmAfLAIdnAH7xtRKG6YnBO5Pw2ohW4PEDfhoMesqky9f
u0iIXl9I+/EJirHrLYLUjCZg5VYVwChxwuIiOF5tK4UOj2NaIUEXQ8apTlhba8jq
srNnwPMQOLJEOvRuqokY/wmeiT/YDySLWuk/1GfevjCVLk3xFFUYipg3kAzP+r7Z
g/73gE2LBa6lZDTmFxiUC4MITiqDSGei9/LDfnSCr9Bd6cnhl4UQwCW+WWo3Gw79
cJN3rbSSWeZCLMFl/NwU9yh+lx6X//6aBA8uNowh1ZehrsRnGSj1rVb0wKRwKJtZ
YTsZ1iGmsFJmLw4k1AIqIWZGMde1puPoBFGF5+2WJj6EKqJnkmCkSeQGAplQXxIX
yb/55sD++Q4MZ6Qs7LaKtbiMWn78xtg+jelzYksh6MgTzqyVRdxgAJwEYmQB43Zr
2PpcqgZqwUxiyFHx0N3lgR170IKd5d0hURz+78/A2ff6fL1OJCSemKvR4+UmGqwx
HtchXhMrddnmI925DrXy+6m/4n6KsHp1oys1z00aM3f+jTs5oeEG3YkCZj1LFOIX
8nRSTYTst48cHvdn5aMllIFoGo/dCijmqXnw15VPdGcwT2gGg8f4StnauEyt8SGW
OkeK2f9UGEDU7jKRhlZZVUB17dpuKz4U7PAtSJhDsnwdNAKwxs7mBVBCBGFx4QC8
0NQosMQfKg3hngbsMEi8LasIHAXCTQMDqOmRCAT47uciVOYLDDfaN0QM2ZlSWq8o
uXdyVwQphjd+j7AKR/SKrBblW2QTkxOlGyE8oT6FPsVxBRHmNW0uY6x4/LEmjE2Z
DLDn5DorPD+WK37MuBm9hTBgI3dWRXLTMJThEssrP0rFMccyuUWZFLILLKnxTUbj
woCOxPlp9JbwiBsQuOPulwFv8jODf0u+UiI8+1sqyBCM9g64NOsMe8HWLIGIbn+V
rzwVZiGyt4Ba2hyAuugCI8cfDQuB7kWkuF8kB/ZaaACkOL1QS1uJ/a4i2FlCPt/k
jyQBRBh8/fAjOt/eNtdDgZ4431UNnkRJQ/k45uHyhmfPg15Z741QdqWeASu2uDpm
6Y1GaznZnursVXRVbLrVgWjaBsFQ8R3E8yFwtJhYgUVKkP2lZ+4pRdtB+Vxzvxww
EdKCqrj/bVaxr5sikY80q7wIKafwaMES/u+Av7SFppVlA681egm4WqEFL4gxb4AH
RpzCkLVcmu9FIwthA3Wc3Lz465kzhIk2OWWkoq8+9u0kwSTzmkC5lfB2Hfs0AwY9
uspl0vxRxt8PB0vsWwz1FDQ/4Oliqjfyqk7G/KArik09XkHv8EmOJrHH/jcfHCx0
bp50IkK12u2ziaUOTi4CRwqlcoXyA4wfkaqaYO8bwKw4s4xdJbuScbtixsf4Pe3A
paW6K/dUIm+K+PQBKRdBrJhb4tlWhCQEXmhVg0VCEh/7tGvpUB1R2f5HBiwxAwE+
ED+a1wg28rEhpMaW0pVLLqKAvVIdVVa9SemDWI+D8C4DbVu/NEWHQPiBDNu8Rb7X
AIbt/PpDzG2wmIxcDM/kfr+sOQjVASNypjK6HIdtFvVqbZbqjtGyL7edS2VvP1WQ
zwDMPeusiKlBpzybuuhzrtvlEXBEAnDWXG0/EU0c63aVFb3wz7sywbjxsyij2JUu
ONnJVZV6I2LGuHEdYMS9WPSxeQfEKtWD28exaW64VLga8zgojZiHeGGPIHQy4HxA
qtlik9qHGOCyDcUgsg0hiCI8Dz3lJnZY1J9ryI6WmxVk6JwtX3dyU0YhUO2r2VC6
zqckX9wgY+EHeEKsqc2IF3xwDe/D6viGcTINJccnxqrXkFsWRXHeSu9tS8tOGf7L
f7Sjm/+CYuM4EauIt7urRplXzIE4Lo1WueOKiH/lETqQzm/MEdaS2JAnZNTS7rfW
LdQtsZI4LYjcSIEdjbP8wwogwM6bhDtcOho5jZFn2EHdQzX7fgt4tZjNI+a+CqE7
I7DTeqa0kMq1HRbmZAbbDWnXnejvyIGK1iqtL1nihC8XEA8y+Ea2hBqNCBpcSzRV
v+dMhiFFJpG/PXAl9Cay/XtycxqCGyiDHsOcpMg8VCAmi/lZDGm7fnqsQKuihSDF
n3eCMtB0/Baxzbu1Km0qQ9nPDEXVGAkjwWzrYjhS4h8CWv817C+CzYdoZsR/H3qn
GBcHWzVDsCm1fn3wIWaZilLqCpWHhBXj8S2ePcOKOVLUCna0DcshSwk7sD4nyiis
eOt1Y64Mbn6piCWJEob9Hgi3FuopMZzSJe3DtCjDgTVKqiz8iKH4n3j0Ke4Pp8Mn
GmP/3OzgNqG5wcQT3ZUb9S9FlOJDX4uWe0w2yJaSpOJ2XLd8I1VbWBb1U/YyOD1a
Ai4C/pmbMClMhdHemyQetfGjAkVGvIAcrHASkNzhrsO9UoRkMk0Zl2uiJQy+8Cpl
o9sn+PMr0oI3OIgNpi2gx6Wi7uGopIRy1pGWkMcG4NIjWOcBYsfMPBgt2JKpuItK
QyfgFVUdWNCduZkPl2fye95atEBAD4/2B0Tgc3mgeb2uFvedNjPpwjM+ayQ6zVYv
2uVCs56ZvGvlQ4D4CEY7/M+85T57IMkd1r6cxWSKzpVnMMdkGSbJHX6zSNNRgVXg
gVVUbfhnavxOTZhEJ8kRNxpSq6L32tRBw+sGe1y8jZRb6jQwYIlqwX0sSjnpUZwX
fVAmtLtSXhPsy/3wlEi/JTyQ/K4qZSMnrZU5QSE2U3/zgmapJir9opZQLWG7RL2y
1fzG8crOXiL4ZW/OLFlinS33m1TyQnXJtdk63wxSODIq8GZc01UBjFb25tV7/EwC
gbddRKDiDtFAmHq8t8uOJ7xsBIgo6SShtODA99tM6+42kQZn+lf6d+BGWVETiFLt
WgUtz8zgWw69CXtRz5QsrWPfi1BEZw+fTH4feS5Qu5iB3/gDlEkh89WrD+LMTLxY
5w+BeNAYhu3sEKBTohKzCZzfdi+ppKu9HNMH9oE8OEqx4BUF/QzXwaihZrGNd4Bm
gJ+/kot/Y6sDtODbNvdFfaQuNaPyMzd8DCx4h6I+ffreBvnEfLrhc7jLw6ETlP/8
iaAiWggFhtTfmaCEo3wvRhzG37U/VIIMZ8C4icrNRi4ACgsxxH1j7hheXoGXBtDM
fmYCeu9ow+oicxopBLw/t1V4ugCfWhukphHH4WYPjzCEKqUFezaGLpKBzPPLAMPz
+/6NqU63FzVJ1ozhPyJjFeyA6hWB1UqVz2Ul20+twN3NC/BImDJZUH6uU48JW8B4
QYilGoYI//QB4G1jxNHL5uVPKQX99VWi5RL3pINEBzlJGxKzb591ipQy223Ez285
YnXKZM1axOEixiTZIkMKAw/S3WhEpwXiAIKyiRfVytIC0nUTf0Of8UoGgZNh5/oc
YEZZt965HZNf+mKTbnAKnmJeIY44HXs4eOUttfElclQFFG+HlfkmA+HVED8PuChs
VwJYnw52LiKvQlma2lxmY11QDpx1ZolXEjojn5Hok79Kh6yhOSW7b7cfOga0Nach
wuwtz/AtTnH+BEFvw8z6+vPt6zOIk7E6G7otFa6Ei/zthjjF+OpBftlVU9CtqihC
8yr2EskxK9hktRBBcWSUHf4K1cK6EA6z0NnFuS7pDTPKrBNlfKptmR0lbYLjZnZI
BHKgGAKIJ46YR+CDB29PScIgnI2f2XtUEFB4a+JeOZBtH95euzINkYkljkXcKuY7
uQsUOw6/Jz7fJjg/smpmjWiChxHa0unUdOX9QUspMiZVNhe7Ma8oQdTQj+OCDgO8
HBbs1Z39T4G9lGCkIWP5lBoOWz+f9u6xDcXTERBdOu+iW+zpaov+D8YUOtWloZox
mwl7bcI7R837A4H8/9+mT4oB8J0gvOqEzMjWtQC46ssw/OOCP8EqGrdPfrKg6VI9
eZwEy+/sar2iYGPkmqAIEg4BAGNvw4ZOgZr5gUY1PMcr7EUEpczpmyOmJa3JFc0+
mysKexaiZUZAi1KD4I5RE1nINoxMmWrAzaoqzY8GoqHZG+QNt/vdm8Rl8VH/KWxU
5GeSTej/AXB2tyF1vTaebtCLdfqN/9UehKfdwjdaNutPQJfgcywfJN3IrKPzZ2i5
6O8BX9l8wYUH0zs5J33mxWIGutl50Vm++q7mxcFb/UfVWBg17gPthXh3aAh5OFKS
Ltf3/lJo9ztd/epPOrb7/HlOy7/yR0QS6qklIBO3n/gt+vYuc1IN2qHayvg1tXzD
3SSaoOF210rih/E/6xLjTmvWKVbyujZ/fZx5tv8iLvNZPX0LHIuXQfCrR6z+zSyy
ZOGUEtK/TVE28KI2i1xEQBlcoMCRl0vOSgCxdHcrhDETVgtRZtjW3XWZB29ejmVx
RU+nvS850Jn40P/kjpFQfs0aQ6Zm+ofaa9Ugvt4OJQnZh9gCl/KfWpZkY+CU45ZC
LgByxqukrFKIkxRpt33KXoBiJ5DAPAFbUz3Mtfq6XLkEfwe24MyVD/3L/pjsP4B+
iO9vpdy6K0kp/OlzWoN4u8NTCiDu80z3B3VMhfUIwRu8yf9HAGOBPh2zBxt2ocPp
q2ENYIjHWnRhpLVnBcmBh1J4TNBEBZS//gG9X1f+lJ7Ym+jIaAj7F8E2lVD9cCv9
ZIZz8puXFMcH5xDtgjerGnZN2+WhYo2EBKU8hoVtzmuPS5ROYT3Do7MogFo08Gi3
/jLgTdy1HLT6/Jeko8FZpKNh1BTfoJPZ68A9hVspvGGvGFExwXbeitntlyQMmY3Q
JS+m8BNGnFyX6cid42erDWwTYhQHyBMo3RBxf7i087DReytXWvlgg2X7Bu9QUELb
1SVpybT6CyjKsCfdjkquG9JzFMG9JU90SdVLw9u8WKRJAOk5CAQf1W26ElktRGHV
zhYvwwlBmiM+MIY5EU0ED+Y/K/XSkaG5pri0lzAlqFO12IhLHLyCkPDdSYHJjwh1
C5D86HqIwJhnZZ1CIAEVxhk27oS3Nt1530pC80sFzlYNjkWttHbfJ6/x9RQRoPi/
sqgfpOrSVwZMIsQWpuO4q2RYkjHhkA/KgvaYFfSsJ+i9wqeCBQpzrpuyziI8CQDX
3d1ahOxuuRKHKsGx9cZdcLi3Uu8pH8vA/ZuvU7prPm2KbrwfrxqMA6cMemrQhezn
VBtJkfpfQwYoqoecXEwi+scr9DZExHL30j+ahZHaH9NghKmJ/9cqYAunCWLzbFw6
oErpLZWtePgoxaUNV5qCETzoIL/gWa2zCR7GOpUhQS+r6+2qq9rZtDipu1tW2f6b
Mg8rfMdvHHLG3DyAaBlx/0V36E+jXqlCQFhipHnQ7lLiUTs4hHEA0YfZrs3OR2nI
cu74mdd3E9bU4/FOY0e5BVGHKYZpGSMPJAjNguxalsrJs57mtLsPogpsbAlvaLAI
g4qBi43VzHoTkewozoZXUEPzT+0ZzJDDmu8jy9iaFXp6xmhA08VzfIaKUNq6BPNF
CT+zjdFGBmi/9HPXEhV88WLfwG9ihQXpCPxXOGw0qt9nu3MH74J7BMv5KeBOUfXw
2muocrKGHrDaYmm7d4kWdXlUI2/z0RTVbuh593zEpNQAA1QF5PuT832kj5yaVetW
9Ig5SSsYXx1NGSPF55vRMcEkcG8ovh0a+jmkNZmKSXoKzCnyup3JBieAljQt7Jk5
l+CKgPjnfXg4dMS37mqszcU35gmUbh9sYWZTtkdCcXsDzv+ZoMvpTCLbscN/xsSu
EsjHiUq6motlT2bBZqFQrx4bmN2O/siNy9hCOClQWPriz5n07XkRF+cwd3qwRIXa
mKfYQ8FSkpDNPz5guKh6Lw/4dUz6X+ZakZNXe6+N0gVQykfCQi08toJcVz7yZWTL
onaqKq2Uqtd+nq11oX0YhIbN8ucBPtaiPzceSO1OUsd4Z0DnlnLZZhQAxJtF4BeR
laWGFVJcjGW0nWpje7zr7PtrrXA9tHDzRTUlemVU8sVIqHqKwFqqECOiD0AipDt/
2iBQm/imsvoG58isOPMh5aKMgBnH+MJlYbA6S4qFFn2evH80bGeJGmLq37GFHgYt
fAm6JGa99Uml8YjamrGDt4M/vS5zoNnEzOlxLqboijq2zoIy2nz5SsRnpfdIDR/V
5ZDYXyqquE0SyAVeI/1ZM4Whx2yWXT8nJyFtmir2xLrjFGde02hfM425ZB+StbFm
fK1ktyRth3KXOOv5HWo4MjokhnxMdM89SUQ8vSxmC6FDFw1kU6PwOVNemi4wzrKA
/3uABIV8l18DzlgvLY4Qdlaqf/m/yBGlDTVeuZpQmFFVyzuYIWgJ0LzpMx3N1znU
bsqI5hys11vJjRKub6WpNo2vgNAbMnuTdlnKOqNIsLXyEEBwN/J0+vmNe7JhSpkt
LEmyyqgCzMZbJlzhzK/aANAmIsglGko7x/KrKyoRW5i2GN/6Pogq3BW4kImMoQeT
mwZQOl0r/h6tYMTfFVDHKsN+KFJQ7LRsaK3eSkQ6G0kaNapngMMt0+buo48w5SEI
XOGtjJwK5FEpE/JFuCetBMwGOVumtZq+PwpxViKBp0cuYQv+u8+HJSfO3Uo94JZB
dbkM0Dg1jzrqcfsc+Sx77rrPV0OSRYnYi1xcwpv2oD/vkznlN3v/fKew9R07zhpX
rVNwJCfGypUVdGQp4sN6TE/9RNlORZZCwakOzEiuKW7ZSLiuOCfIYBvsOLihKodD
8XAQyrgqKZy6MZ1wXYgixnn/o6rBy3ZLPRprxH68hCcZK4ip5kHHijPq+FEDbP4R
VZ4xoh7C4QHC8QnqPNNdwd2o/JR/+yYiacfGcLuclNMaN/Qjj18n+6j4CsQ0yNFe
dL+UIFmop6MBAXx44Lu95FchkkJ9/LU9aTo7JA+AbO8zRmqrb/+wxBqN1LTHmM75
083FK0p9ebI8brqE2l4mGt7p/4swcL/kPNLauIW4bSwXawSnnXyh02QPYWbSfctX
UClRLwJg6o8j916xngOAM5PV6YxCkkOmpSumRkVz/mJQw3OvFRotWdPc5nEBN3tb
Y7uH83ZwtRTyAMWa+2SOzENLnxwk3ox0pQupAogXjMCQcIuZzuVUzySKCxOSZmu2
PsNpT1pDWe7UXEnrtkKCFdR28k7qnNzxZ+0Cw6Xlveg2NPE7xrv9wcLudinVnurz
o6JG8ctAr/XF2wXGhn+3zkOAMmIss4qe/sgqL2c1EIEehPsjnp/OX+VxcNeitqXB
NUIgMJ03uF5Gi6HUFJhrMa4rLOlBq4799O3WCDESVArDUDWnV/pziya3RQdExCDa
sSB53jKokcmBoFaUNgVSfJLZarextuAbdqjYrsKbtCnpjiZ/0EAXCXwOo5lUVbrZ
+nRnVUU1/rjCz76ytzbKzGRN6VcrpaWrtkk5Na9eBq/O9KE5Rskxtv6ZabPdzhpv
tF30KV1BkThTLg1XSIYj1y1DC8LeJgFv4diUoZCV333oJJf2/iun0iIa84tl2jGb
ivrYVCCTMjQSm/wKs6eB438WI4kBzkeYKiGKUDuCGvRxpEGMWc3UIs5tSnxf9t6o
yVopJUaIPoGHidLhEDQ6d4FEJCUaM5Ic95Ptt8rbc3MEKfdHkAOTgi2rpYgFcrMS
2J/U9iHfU1tpDSJ+7vfK0i4iHqiq7OcoupJfTU0CLmIJ9+ACZ8LQVOqgdJCYiFwz
KKOCHit+tRIhRpUYHmRqpmwC4eBI/ZJLxxLdCV84pUJX2pQsobQpQF1W0Yre5Y3s
Y1l//BiBFqU6iErzQro7a1uITQNJJtNX7zZq3VF+OhcS6upbHI4NjlFmZxhBauOl
z+x/zluSpcYkiw7nVZR3zNyE7FL/Dey+wm/SO7x6YbtDAlOg8O/Fv2JyKuyVXWik
r0pmAu+jb3tQCue9W9cSKJlOXLEiEKugbCVM7yxLvJsnsl3/OtkjIgv4YIiBghvx
sBgOAaw2hW/8KDcVZX5saVjdHglUuJ81tTtt9rzAcQvQzvw00i7Ohh/y6GNUuLnc
bKCLHeb4oAn7bqHs+hpQhauWBwQihA6zdQHfa6JUbwF1MNuoUyOGfBNvvHYhsxeq
ijBi/1lDXdDMcsGAA6lDfBBZMOyvvM9fezBi+BAu31lv8QfJm6Z2lIzFOf72iLON
p71vH7PUB4UxM4eyBdTQryCPQAbAFbkkJBojey5HlM0ckajyYrqpYDuV3KwvvIRy
ybWnK0zBszOfIi0zRd4+a+N5NHQhWm6KaBrmqldwz/8RoDMpNnP0LuoDORen4A3A
HpirIuldHHden6eo/9gz+66ISEeBjaZKbB9zE7EGfvC9ea+pHqnCCukt1FZhCN43
nwtAXm7L9ji5OUtUskoEmYO8qnixSHFVJjWuyukgoGOU6fUlOPEv/q5mhBCD+1OH
rwlBiyyqOuq0pkhZre+V7klWKi7diGQUXqSv53fIliALJHJRX6ssVsMObt17Ierd
ek2f+cLpfCjHl7Dq0YQv5Nd0l8UQqKX/xHRN7rIpxs/A2TLu3x9b6JMjbt+Jydpx
QLTZM/VChqSSaIqq+XDq3DSyjFQdx17FZLb/zQMCj/JHOMCeNLRoayix5Hx9u9u9
a8ujgFenz/sKafxzY/pQL/kDTjr623acWMYFgDzL2uVVZjGaviQx7aAIIwDeuGpo
VNMZLcX+smlCXZHQLaossrJqc/ehu2kO7zGIbPGdbwb2Fc3w9GTuoJLl8GhAF/dd
ldY5X+nPZjBiF79z1R82eKOjdS9PfrLfyqsVKGH2npmAWFWnw5izOLA1SykaSxIO
wiisEdb+zaQpHLIX/JQtJat5F2JAx1CUynBrYkxX8SM=
--pragma protect end_data_block
--pragma protect digest_block
kYm+3xoogugM725lqD00zrTszjM=
--pragma protect end_digest_block
--pragma protect end_protected
