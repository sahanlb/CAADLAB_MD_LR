-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
tN6uSX9cTQvTcwnIxaVAw6UN4xuKS1GINgpEcsJrj10j0Bu6UgBxZs726UZDVJ7T
X0gojstJ4jquE7G+SGIygnS6p/Al4PzstFjUV3ws4YBx7q4xeJmrpJe9VGVDiEPT
npF2igpEt2F3DUEEZh+FaGs2URZXrtCum1BVUHY4pSQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 42976)
`protect data_block
BvvabmBU9ImWMo+4XIDfeILhWwGmCwicAnrnnGGoSf0hp35UMtvq892oNLZebknz
g3v7DS6pYtC1s1GIovrxf9PQLcq7uXHFlc+i3+8Y7Mm8vUEHhVM4lcwFiYNzI/AX
2fXEtYk8cWHz4lqiGX92C0MaYIe2GUkvRW8T1+GkWHzieddGeC8oeZ0fbM27qW5v
iu8+aitQVXX5ZjzDElx3xLUFrZTvJjIw6TiNgloFvESLIhMoYYJ4xWV2+EIPZiNQ
FqHyu6d4eiIAE3hZtc6SA7K+M3P7cC/G/a18Glct8u0wHStmqJGdo1/jLo7bRM86
h4k+LBB5gy+/FQMOxTBANQU3F5yr9epHbuFJXAsm5F8hu9Vf0FL42T31g2Y+Y0vt
xe5nPwX7EnGunHBSpiWB5oZquD4fHMQUa07hx75j+uSImryTQHKG3azloIGuMXxE
qgaCMsFaEvmX0aQSv0tRzHwtyqCzz3AkAgbTfm2fRrt6Y6ogN8aydL7HAAfc5XQE
TXucMc3QNmjb8f/qpSMedrGa/fXXj4oxPG/VwRKQ0jp7+E6o/oSf962GmyQMGj03
iClgg8OVrpUO0H9UeD3HGdYSVsMTbReX0tJV2CPamd2gykYr6g/l6Ex8z9cvKfJc
uzewWYz8IyQ45y4xe1zPlfKenTogQVBY3iHUBXsfz12S2WMbfDe7iPyfeWyw85I3
FQCC8UO+/w865HssZuDfL5MdVxg6bGhztep11n1z5e7+vf5nbT/hpuJB2mWWNT/R
neFgwYLnU+DCNH7d+Awa1H4pHD4Va5uKFwpJKB5dbnDBsJq0jOX+GNTpmxF0M/Pc
DLfEJK4h7582FRD8/GFjW+oeoiwWkCQFrbtc33fdlahr8e9BjwvmYCoFw5qj6FXs
I3TF6R8l5JsWi12AcTf5puM6qtb9eExPPUcB2vHZbotQS7aWZX2aDxNxuO6SkeVQ
QcoFXUio9jWzqKBKGbqVFKt+ggHVH9I9R5R8Tudzm6RMVRG7SkZVRuOVtOtXWxOB
VfFJLtI+uDOzUZljUVbIsxjVOdlmk19AsTA2R/AFyIg2B3T7ivqbGvbrS8i3XAt9
UQZ+L0RjgG6QPVKsTWmp9iAEImQpPmkQ46ssZ8mesN4iASTBsjWGDM5wFVmBn+/L
LgZp8zkexlDIs0yxTw7WU5USKTSs965NOXdrVypW57tSpISxQxGrkKnlabH4R9DO
09FtxdMqfgwQpHpwC1jWeUrkauWNH3NBNFeLp9D0UuAghN0JRvAOaD4LADwTO9pE
YjlM7N1nsgX0wjiCNT+U9eiZwjwI/Q5WYhAotEDXzudMenkYu4cNZnNunFH5D4hx
oo8jI2yHIW/bCBrgLal4EquEktGtOIVH9oeppCkW/X3Gk6ozo0A8BsuJwNwFZ3ZK
6qKxt53b5XnF/3He9Vy8XNlNVg8copi3ESkt+bfXnTUJqgWfivV++8fMqaGYOybI
VQrBf7viVMd5ePNKBhku26p3lfoRi8cKmmUUAG0Fdugryzyl//1QAEcWSus9+Mee
W7U+CCTRS6V7MSPkPtc1LLPy2CffaVGvdPRaD2TfYV82RHgcJJe3YzAnZjR+O2YM
843mu/cqpc+wkKWTQ00gDOSwS+zPZF1ZKkotjwk9yCha4/oIlvUSvOgZI/+Pb3Z+
XEeGCqzwajKcfoX1xBgl56IJ1YAT19hho/HCRksLuUpUFKdzXVNabpLL937ibnFg
t5IjI4hLqBV3qxWBb+r5I2cKXJ2QvIXeClc9um07CsW1Fz3dOzSrdAIY2cSRuhNH
BeWMXxFQw6DTp4bPooVC+yTiSG/lcpukQX2Vwfmpjxab2+NF2nin/ZFSzIlalfqh
q7KoQrH7XB3lpPBtNdEV0sxogS20z+iRkubi8KNdUAqOlQ0J3d9gSuebfjlvxMen
G+LngIsSqnckdYIRhRhIRdsIT1IZ5EoEft6G7ertm8DyfMNdM61YE74L+eMPOc2f
Up2regDlHq5iPSq6wPR7pZ9Ao0uw/2hq1tz+VvS9p3tbkp4Hlu/PEJuELZqVezgd
PnVdFMcCTP6y4iEv7Ff6GfuJT5McU7grMQw4AMNDDxCKMB5rpmXuukIcpji0s7zs
3D4n7tl9nJpZagqNowRl3iaZunSJSDVcywY6kxqzdFKlp+Ss0B7jC3c5ePr1TmQQ
7pu4Fnx3li7vk6TYYIn1d6jq8lDEYDrH7GRw+WsBYVVQ+e71sC494c+hOvJomhr5
JpWMUI+GGvfqjyoJPy9RUYwPPpgXUuIHkPgZRbISC332zBAWnw8tIj1OR52u8kEW
2tYN9TURbJQLarGZEpJUJqvJ9Wcx9sfKWkMBv6/o1b9jbRi12IX1yqroMaz7Mhdq
gGF93eBHzoO7YHm7Dz7KTvGSSmLBxc/JcAf7awh+77e+V70HxANtPK//gUDxCp/E
nG3QkVH3CghNzmRoREDRbEhE9Ocef7B6EEpyuBUOQWOMf2L1TRGYeoEKCyR2hprF
VIYNr19VQf8Vzjf36rUaBhZO15gT51ZOqcoEzFF+xk4z13IXQkk2R92qdYlaqYdy
veugN0Zsvo8dMF32zk3HmL8UU5Qf6xHOwCfw8JHA0EuKmTStM7Pgz3fuuX+eb4R7
DjLxAlADVAgNO0tR2wg3q801eoNQa3J+HFdNNeezTDiV/P0qFthp5X1WXSMTT7YA
gwBUUhtOjuZrBHg5xp7yp6YYiZZojRr1EXOgyCwfBm3dMLtrWJE9003AJDsjyeSi
e+Wsi69m4QK1pgKyQeCH31bC7/2xEMuxp0shM6pdtQ6fU3lY8B2xg15Z9HANlCf3
2arSmUyApKcfhlcWAqOkbQBhIkba9OO67Refca0jY/f5egg4a4wFivR0L/gbPfOf
BXbl0OLVyRcJWL6kGfmStGmwE8JKPgFsIiueU8SfsphWRHHo2YDkbOfoB5rUfo22
pkdnfHflUIrXXI0keuehVdmXFcEzuC9jfUy/WIaBawCddDhysTkGLrwr8+J4oh02
h3EI89nssL2224T+hSppAR+bcCioKLbcf+iu2Krt67eKNW2sawc0p8iXs10Ftymu
VqYhmDaPVlFlb6Hf1JbUHicVYBsIGDvPzqwhF2r365TdfgVNfbz6BoqqlTYwSKNY
YZrgBg/0xigxkjOyW5Znp4CNHpQF4ZkzYixm2Qrt2uUh1/+rTdsUc7XrZ3ORh6Ce
ZqzySBzokPVa0H98GqmcWq+fFHl9/bngse4ul2XvhSMpSngk5uVjSRG7NBaIogEb
N1w/F7+SEdpdiBH1iNMkQz2xV4pwGaQwsrxH54v/QlkCemEgqCdS8sOu7ot057qP
1o2eMVTBw7tNMg/blr8DPNrFJ/++WQVfKdESctg7lpfbwfCIOzQNfmaCvRMb7f0y
/9k31MtffmnqIuJiRHWI2cNl/PefbI6/hVDoEvdj5f45q4Mgecw+1LksB3tSCln7
0uVmI6eDplWPPePXL8KJLM1U1nxRu1/qS9/ZvZEgUZz3pab5F40xezDbqh7MDDso
kHcruTlMF1jA3tSdkbl+6ke+XJnKP8bsBQwlS1DVvE7EB+5OrA+RnUYBnETOpL/R
lXdbzrT21I77pJ51fFXbxvjN34Hp/q+C8FbEON4ZHZT6SKvJh5siazt349oCwaQy
2DrzeidpTJFj0I+jN5sUPXBQPZgAdN08nabXN8bv6B9vRkgc1CwuQRvgQ/xc7XL3
bZjC1F5C7xmtLhMzIu57PDZ27SWuVDew32zhSt3kXCC8SOKof14bCb7zwV1mDXi5
FrS6YJ9cTxii2cQkZJ7334xIcnWPpRTNcWRbiR65J6OQLqywtp02YR7fZHTayrFI
q3ySFwk5IP3n+0D/ZgQx5S4/bIh1D6N1sTjPssyALYp3huS8MboLgG1jfMol+cJ8
6pqDoB80v97Pvd7AIZ6y5Zkhy3JW5mzjmzOYPjXYdPTy5lPqePTPD4pNSM6omBwu
HCyzLvCLM/rJ4WtjA0EN2bJ0c6yzOABd7gY171td4xAQMTiuJaScOXUVBHV5Scab
eATaWq62KNFKEKyHU8W9l2YadnY8SpSb6Z7aciJopFKifMvNgYy8cdGbQIwrsJPa
WzZLQJ+B3xl5+bHYB20xlX1QeD+jZl9QYdH2TkIXLbh7gUSi0IC7G8JKm01JFWY/
Sw3vPPMGL+NHRLnhVyqkFu7gSq+1LzWfAQvMZtPFBdhtrQFPfJH2DfD2UJGIZBWx
70H7QDjuMl5rQzk5ADtN2a4glsegfjaEIV3DRuic7UMBw+WS8p5gncGTJgE/mgGV
WmD7dHoJa5x/NNXtSceOSB0MUMNHolt/zadZzwUrRYZPN+X2bBDzP6bfOtMgb3Us
irijan0+wontUOcEXn5gO4hZsJcOZ2ykdXMXf07QlqFHRWA8U3PON4VS0wrTlhnX
DQf+R8pi2lO9j2MBPLysLgULRWLz9tgCYMKi50gOg9PsbJMzKTTol/q9YCzTgNQS
SOceeIv809SGQ7NyeswuN8njgbWkDGAFhbYlPLqo993oiXBQWY/8auyFoG03rmy7
WQ6oQrTQi+MaEJyRd3WIot66eES0OCv1l93eZi+xxgkO5vtoo8OHSHnjviK89rK6
brAqIE6WGG4jQk0GmTK+zEd8EJdr7Ep22kEockjScESBqO0gjZ27Wh8+AHPjqrBd
FjUD94ti0/FDK19pwzpCHZxOz11J7trQ3fNYdlEmpcy4itQit6gnoBGkCGfgjSUn
48kAJgRSUhs4a4aY055CODZ/AAVwnb6PGxupCzGTJcmJ98SSUlUkvNvw7Mp8p1PK
bDWMA+Is++qGBcxGB2i7ZilVL5NU38VE7dQFbeeXiAA8yE/FSp9029ZzDsdM5wiR
UdGYF7Kcbpmu5RNpurzSf7Rqw3ZK+LPCf4WW2IWRVvpzwsfh2lIxkmrz9P8hD3/P
+j2hPsW4EV8Hafeba4BlCXLKEidoVuarWkAT5GlngprjEBQ243pIOnCnvO5g7ru8
Egd7kCGYEAKTVqHCBcZD2bg7OW6Sk2CRWTiPXlnwsYAB9laUG+by4aZhIUt9fMif
hNqMAVQgDP1M3hkJwYTW2FhTRyPOL1OtIHJ+OPW4ClPftU+Xk6c1Q457LRfe5x9q
Bj5LvyLJmdtxDuRd2ylsg7Blgfwr57Mpu3V+Ob6mn1lGi6y1lmC79n62belerwHx
A1DNMZXxkVAK+qBX2CJLKzA5jow+odScGuj6sPr7Wz7L3rgCbXr+gsfya3l04qnd
iYWfyHGz1YeMuy9ubkM5rZdiyGBfAFFzqA3u9YErutgugk9UDRh0Kpk617C/AfdG
lRxOHCRx62NU76g/4mJzzZHJBsuCKI9nvePas4NSGyqiN7fy/GXAsSdcQ11RSnht
j2mUt/20S5oSrAsS+5bZe5i410ub+DuGz1sHDgz4f8fmNJXnhUKVwcdLMt4AxbWD
pdm4eWrbA/XM5GwIItv23QgmhWLyl84LG55hb5H8a/i1csnZVjS/W8lWMRWNgc3x
nCIOwnq7z6PKUUCEQt2FQcSSG5SgvmISRUgQJrBrMTdiFbP3H4UTlrWi8Q6X8QUd
kG7OUamkkZFEc8WNpbSSNjtM7LtAZtqSdNUXlIDVmp26G1if5aEm9bZJSdrsVKrh
NKNPu3JZb+x+iyzmogCUfSyVEe8SO4CPtGIUH/WX7Ik44fYjvoYJDAVQa+Eqes+m
nDw3i6f9Mk5/IkKBFOvMGUUVLjvIFyg0KAPEHRY618p8INaz3d7qR8f7DvPj0qJ5
jc/KHeGQsvqcre3elsjP6jWdcOYhRAlRR2NIFHnjyLlOs4bSyjaAiQjJxrX+FPwp
XqTkJ5hcyMApUDrtA1EdWB4irm/rFSXsBXvBv2O0eQ6i/uYoYZmq3jN4ZObPUpnS
Ha0bhvFkZchcotSvAPHm//cKI+6SpSBF/qRm53VEGmYPretPq0A8RLNQgp7BcOVO
v5vGN+0/OwItwpkBVxCRyfqGZtIsbldUWKKFULWXj6WVZgpQVdxVe0sROJJINB68
0DgZiSzB2VdY7wd72/yUBS+/GeWVM5OEgzOkCF+kAFzujCDZ6GXssnP31+MK3EJz
BQuRn1gabo0Mg1WZ824RmU/Aplk5ufZjYtJ3/cbjfpetscvMGnakoNZ/8A0gmnOk
K4BxgROx7+hbySCBeQcpSZZCKRPBLjei7R7TcZTvvz+YaSj6NPhtn7HtobmTXLh0
mdhT6KFXmOilAaOBo4NBkBPtL2Qgfg9BWEoUWd9hzz4IL2kio7tetUTMlnWqCTm5
RYf3O8PBsk3BsJwmAfptjDp2OXgEKDNSnnFSRWEfRgACdWhvDn4n+gJBzaTCENiD
JL3Va+EW4VThgDtHMBeq/39RYBB9+pzv5TMzTh62AtENV3xf+kCkLuEOn0nFE+W4
JBQmTMOaYYhM21VAAnQh0gcqvlcz6R3cHk1YzAyf3BxpaR/X9iyNFQq4cyQYoArt
ibOR0fLxaIlUuoq507QOPRlNrR3pvmNv5S9EXBYcuef/aVraN4ARQSAVWqnbtHdp
R9CFprjKB13jqSGoCrYiHUz/QdsE8iQAcm/MNu695vgv0npcTvomdS6WqIdZif9r
58tjbXU2rt0ysKPs30rVJqMNOtVaJBG/6LIlKAvz7x2JEEFIWjcaJ4ybjoFQO8nr
gw082in4zJjX8qFI1Cl6d6bNgfYaNWf7He8Zi8WWSbSMJtyNu9RklNNZwmwTWKaE
kR2xzPsjpmetKOtfG5jb6kzYD4Pi/PfkWdN6GLJqbiSHbFC25utIS7wUOPUN7bVr
t7fcmPuvxpxt7MXy9/we7l4S0Qa1xMHFM5QOuNYscfmRpVYWiG5EjVWOO+QldZkh
iOelKJckl6aud72v80K0KU0i+7faQ0EAI9HQMskC2D+v64BWjIYyxCkL+xXj8cTl
t3AOS5L22DjHExYgjYNBO1mmJMcn+2eZojX4u4mLB9vspRMx4xyjXpUHU1gAb6G6
Js05AktKYNNexc7D+CsFF/HrsY0zf6vzM0GBBnlu8ipU9GzOQNMTg4Cc89gDnKaT
tu7YyBPXp04MvCj3iACPN8WXB/sgZIyjurqJ/Nw0O3MCBVnb46fXkdPV+Q3fRNqf
zyt8LbwHIMsBrh2eKzECPfpmP9E5VOCUDmlMc88BRTPCc6Dwu7KeLn4PIGXlwrcT
eZcnWwBuTxkyohAG8kTRBJGKE3UL7OnnuPO2pDJWeziVLpeMx+NfRFsdK/CpSK9b
WTJg4g0YHvZQskBYEUZHlmbCZyqzvslbtix9jbh4G2iMIh3Jg+0pNlb1+L9yhT9D
PeW27v6GWLzI2F255gcaomneO31yWmaL69kyF1zj9i6WjIDnxIzwVG1q0ExOSSRa
nvyJJt3A3WSGoDOxHejQ0j3zscBsPKXSpgQc1Rr1Y3uOKjuFmR3MHr9SbJ/DpBjb
26fzLouP47DQEDP1wBSV7zGHd3hjDneI73b5AlcsVIOvMEDujbPojZo5KnnBlV4G
Kjs1tYwSj8FT9L3Xvt4SfoWIylRqACNLiu5kiqdDbB3eL9OvctUndEEe0D06WbNs
8qBnV+g4P7i9cdBH5ktkT5lxjRzGE1vkPZKUdP6Y0ol6Is0oERxkbNZnY6ZvgkNj
BEKkTf8VLiCYqGy/V0gUpVhWi0n91JzfRJC+RhyAdsw33FRBeqxDLivh1HKXs8yH
+fDVJrRaP0GSQViSC4e9p45EgFkcxPx3o4KbaHvYXEL8Us1Upq3pJbHo1cKRXzeB
rSqdsAYw879WDUzfKNEey0nY4qhFUZzcORcGy1ncZEe5WmpEWy5r8f/FFslSeJ2t
bkQrPfVXaIXYUCA1+eslQlc47o8tVXx8L6kKj6vjYMwbCtaasgnmpUhJaZhb7xzR
vmte804egO/drPEFJbkE2r4DxLa8wXTMp91wPasVK2RBKm6fvhk1IuCbHHl2Icz2
jS7UwHlRa9J06XO5xCwnYUTQRJgHlcv26iNpSbPQ0p6Pnvzu0oNxY+S1BbKiAMQu
XYJ6vb1lvdMTuOZg5uPMHpQPNy3VUIBJvxd3E6S9d6qsBS/6G9DmPkpwEslLuHz0
gMzlwQA03w6XdFye2oPnsD2BFTa4B+NzzqRVeK/+TVI8b8Fv4B8PS3kGhz6yUCuN
pKkJqTxsaxOhg2EfGGcOX6c++LYMIt8kCNV+/6COWl4xGxKvqHNTBT7F9Or2Tg1j
BQXEE/NWBMHw7QeFeRKWAF5MWiCpxkQErHp2b0dMyYlCdfHEQwhVrB5EYnFmCyk7
+E+/VWpufTT2oy0UHeyI29iNTo6rGkX0sjhLVnwefu87ljWwcmPxhc+h4zjbyMAo
a/7N2heKuD1mnPnh2/D/S9RHY8XkQPvRKoFp16iYdeq9pAxcUbaO5e14qcbnTnw2
BhLpXLc7HvicjKg5/3p9dwuWlVZcVPU4rKeWNyeCmBLKhELEsVFbiwjI1CjrOOmb
IBrFD/G3F3Bn2WB2QQzKwUxwxxBHqCMQDizSpTzyzh1Rc7keZ9eFCjq8z5kZ+EGw
kb5IYga8G1dFdwNFs3Oh1Gkt2wEcr2ECE25BTlTvWvlLrj+W8lTqUxPdp0RP88Vr
w4QoVgo8y2YEg/z5k/HrDEIrJXgFKSpGY07zuNTl5CpjRZfvuS7917eJfJd1a+CX
0LPptRFE75i+NhrdZT7+Mb8xDZeQ8WCPgN4VuhTmn6vyWUOuCZHARTM/JtnMD7oC
p0eX+832rSLDxW6hMvIFYI3mX89+viJ/sgTwSHB8bKmYIbgJplTtDHNnPb2D2h89
jrFiGCwKlBJIKudwJ80ilhi5r+VvaofX8td/Ke5JLoY0UVe3F+Gt3/b3ZahRVbmv
tF/19lMU10Qxn3yYMxDfbxVl+xtDN+FpME7xc33Wd80yjUqRxwUVIptTuAHOAAiG
HIgtVvkrqgYRfHRiU4O5t8P6MTt+KiToXFxi4pDF9iaFG16531MkiN4uT/wGzeN2
vRzm6vYwN227ueMi0JC/Cx2k5Zld4TrtgRSjYqZc/ZbkMwbdsg2lW9+9G8MZeGzR
7m5A3D+E5WXdZY9Nm3xDAWtBCQNYK8QSaP9nJ9aRrsxg9/UFFqyhrPfwq1sLQd11
yko7wZyquIARhUeJfgntfUbURNWzp0e5cyFg1a815EdJjDFXUcLWY0UfQ5VRGvfn
oSVT3bPR/12Em5/rSKop7zaMHzRr+t1meKapU/zse8SCwV4yagkL0FBVYvjg/3S6
gwy9UpcPusHENWRhZh5HRTqjuh+2qv82kJv1k306L1GwjcNCedMguf4rbaQQbUAl
HB1ds4HWQg3MBpRusG61ijX6MzoXrwEgVbO7unnTUPoaC9DTqrmGAUVgcYSyc3LO
8spgtLUTEWo65F7lI1mF3t6QPZvN2Z++sIda1n6Z6EznDtMbzrkYGeEZdMqhQQ3N
Fh+ik3V8uz+bGTt8rtM/IxJzjlUSH8/pHtmmxF/3rVlYuFROb3VLa+BltMA3lPO2
s0OjCQsAnELnF71aPJXWbLX1ZMidVSYpItkE4OqOGFbsZdq1k/hFSpRdu+pPsfFN
vOdeRTEfJkP8lE24c39aXmR6V/H9J9mEvAeEh034/isPmH7Yi0h2lMs402OINgM9
/4R9xBH49WREtq+Ceul46BNfBrsZVfLlQa9iVuwRrTq8G/sWlOpHguNcfYe3mNYO
zk/+AtwWgNMxmKn5YLlYlSu7ds/QrZBkupDQRP3mijntrL3CL/EdORXgQglVCdby
iIwA75fmRVjtHFozffp3uNj9GQ8LcbldpGQMPSb3begyP9i726t5ZAGTScuPIKWw
DowWRIvUtok/Dy5IWYFYxLS11bvte0pqKtSAOHsMEqAm86zArPReCDnSMN+iKJPH
c0eL7VnlinpAoVgRM4GMrvzLacwnMqKz5JNGcn1vyKsKfGVuk/gixaAHthWP3URG
kmcuJ9OQVG8Iiz5MqMLIvslr0UPWKea/r7eCz26ItSIfeMJTz7C5DEcZPtcHqjIx
qyUbdpvcdw2xv6hdKfvx2SnMy591u3hptsotNRai78+zfRLOw6m16SDG0Y2Yf5Wb
BR3AgnQDhsuPhC8ayHvMUg6ftYex11ltuSXmzL7xswLrpF7TtG0SJxILNUjdB3yq
dyausFhllE9DG+BEdgV2qc1VCHLlYi71uf9ydH9mig7NvKZnPnfAfsm66HAPJj7r
L6IN38mITFM5XuA0w913tbkQ4k6A/PjMtFFDjc4Uwupp1CbI78mtub852a+gCxMI
tpf6vR45OuwTQBDILXnx4jSFSV3PqowJ7a1lrTszVig+Oa1+q6kvRD+cskHAW7NH
CCh3z0RwbW4cAIkP4XO2YHdISvpCgNw3HjfRG0C3hIKXZs4zVzERtsmmgDOIvAPT
IeWRjQTVyq1jmX1irP4W9kWv3ya5H1s734KcZ/NdQdglZnMg73zF35AK332l2SCy
hFoH2mkL5IBTKiAxqG2KjT25m8cUXWeQVY1T3gw+J1FJnKGJvlukaEZmJQHfEQBF
cutkXyUAJ5X6XY/MVHqZ7yZ8zrazr04zLGfd4dDDImn2yioSvjOydRx+e2krRoFL
oqv8GIQyUr5U9CzXqMU6/G/EoIycEdf0pI/eivq4sT4Uty5IO0iH0sz1bM6rHum8
Qkdbi4i9k/31MrNa+FO4iNr82wOaq4iRuMJNzWQYlTrFeTanfXIj0QaS0HczE6+p
8St+Fb7dAUXKxKxGnujYgI2LmGsoL42K0uzJvUI6KJ+ADZs6L8cUm9qztWr8uiN5
z/KsAbbHBufDRwBSkixb8ztbSh8xRdvc+ax3NANMncb/z0xx9xbq/lIgpUMLk+rZ
IkGny+wu7i9baLQvHpYBoDiopFiSJBKOCbWPwLFnu2sUbnzlKZKqCaLmNx6PjAbI
4aJ2SKbfuatkudsQx/mXssdl2pWvo0J91yOIGvdS2Y+PKZRuQxeE+6n2P8ppBEw8
a0owwn8Dx/JAXYeCsLEBjiN1mezi2LYYn/kETASRJ6PV2z2UVJhDKWwDUQtdg1fC
Ecqh5Pg8elKyp+0HrTy8XVT+pfjHbuOmTO43VLP/MDIslURnVfSBDAV3t1yiAt21
sga3OOBCDPGlpY0zUBViESWrXoCVnSKHmR0TEunJ7RvhPaNeZMM8cG/g4gOw01cQ
UgdlshSKv8E84DXZwP0gGErs74TLIZxHJca865AGhGdM8OcSirVoB6h2H2EpBkjJ
r352xnD6VXxw/ERt4zRh8K8qgagnWyVbLIE/VyXyPzQS/pVn9INdm9EBY3yFrMDM
iyeGFe7i/5JTTfA+iAT591urFHRd+ptTstfzeQubE7gIH5JHX5ZCTD7eG1dSs+7x
uYNMR5toz3Gl+Xff0ilxGENKNcbDBwTifiaG7DVOvWQOahJ8vxJzg0pK53HohnEh
RB4ZZVUdOLYDzClpPNQWNXuE2A83FjjLfEtR31rTWwv5MxtaDq8JhKpqolXyZLPH
8O1GZkJaY/jML6W874o/MIec3YumkKR3zR0IL7G6Wb+Z6qCwla7P7+rOHRVa9fnc
D69/6T1ilvR77u3WTmI+5i0OTPASDakIpzgARv5zv54x4IIJ1lFrsHH/DciKHZXB
tNQ6oAfeS1LzLn9nLWuUi+DRVCqQ9mhk0KCD9D29JPN9ZBpluBF6Bg9mpbvzK52r
lUbxctRvxg+n5uAZ0WBKSrwROpirsJqv4ZE2FD7CFfHkr0zC9SkNTFZmqzOCea15
IpSFJQTJK466u0HDxUgOhY5rT/PlgTzZ7CtTExdkU73Yt9z9uzeVGEnAetXwYyVZ
yCeyYv0KJ2i0P6Ut2xp4odkVjiptakGBZGg/m9DbWOf/cIoxgvuxI833Cx4yWaCx
ADqgP4Q8W9rrj/slvDT0L5GWUxGJGMDHpZFbhwrdkpGgW+QS87dWnkWQjPRf1haC
IAMTGkOZBeAxg5uyhNbdCnXxZpdEYlgSjT2+M1ZbkfhSob5o1K6BZPbs3qK/yFnB
E7olwPSybkJgQX6+gH2SXd009wrULwbsBiiQz9glmzWNpUPpdhdgRSmhtAiHFrf+
KbgDrXfYXThTFs+Qj5tmk6hwtiJQIZawaaqTBXmUbRUPcz0CxibM1XIcyPSd15za
5nNrMAfXYP80FbAX9qkmfIYHtzAVvRy7xd3R6t2M7K8uFKI81iiYXOYDwzTpB3sS
62eBe6Bi28ZgWMe4GJQZRtPftzqFOZ+rQmEdJVMR5h2lhuTCIjF4dalG9fX9nJov
BmhqvtSE67pQGp1A/5sWafT0/l98IgKpmgG2buiE/Dt/l9Izt39Y5XJI+qOxQKoO
uF5S/uwcA3LQNgqnE6bMGhBK6kicu+141s+iV4UZYG+okZFdKFl0Rce5H/b3hHdm
//LMShcN9DoH2Pzx750J3xk1oZYmOlYG1BN9azN91OM+FIUJfqJ8JQ0kqhB42W++
RdyvDZTLBsZhsWCxyC1i9pa3oj/wLY8BMH/dppcz7KFSaMt52NvV1h83yENuaEDk
6savHoadznBwS17OJOSLpSXukxEJxwIxUCL66zAo+8i9isSlliU+jnCOm6+1Jlhq
crf8H5gbi6SjH9iMcyM7ycPCo/b9lDRfPPj778F9rBqHnALKPk1N4tguEO8l2kVH
ZWg4ksmA2EuVBemLeOiEy4KDAtrUYPdg5LHsnGGZ/KaHqSLRpD5yeQbqzXjfAGZu
LFKh/n8ikg6pViQikhDXhgzR3hFF8f4BhXunKN/H9CGKolCY8WC5OlA7fVXA6sPa
SKyqret1nnnK4q6G/bk4GpitfZshCHx23k2CLUwEsNzzw3VtL9db9Es/gpYKtmOx
HlIOer5zpPdtoZMyyfvC3z0Uk+8PXzx2bSFl8lWMfvraRTr6gCX7HmwWxcbzYKTk
70ezMNlbzV+jXMzH2Xjd/g6egjGAXf11XmIrtkFr6jmeXOkJ0MTZznbYwiXshQF1
KxTl6GOwIQ7MkiqVu0Ef7DlMXvIH+wNltW6ua5kFN8aVUesoQNq/72d/Fnzh3ulj
VLlrL41qd3L7kbAG6siqIg4eBRTMWJ7cxv+BKcOxWF9Onm/ndx95NEK5Zhro4LDq
4P2kj7gFd17PsXVTlKF6gH2H8onrpJ5YEgd+o4q13sxTisehOkthx+cdix2k6PM5
GcQZDlFgu3NtlVpO/sKG1vxAF97MQZTSKud6SWV9fxZhZaCYI8DLt8b+6ewzbhWV
HC06bR/n5sUDw2K3W47vHoULM3SpIRLgH29wiG3iHodsCPyeSUwHizX5q/eNgIPx
BcYPkLniKGmtArjkXVPYJToxLpr+/17rltAAThlpMn2U/3pStBzNb7LRqtwbpY8K
+OPQHowtWVh+JJ264+gehp5SPueG6uh87X4rdi+1Y2HD9e4HB2w++wq6VIIcnDom
4y8si8823HKvPtRMJBPVrdXIXqNJZMJNb2zsnrJmKBW62FXsSqYCY9yzKwPeWzcP
MkV0j21BVvoP14BY4oGt5IQrkCFkXqx3LkhL23LUXAz7x3VjIJDHuCo+5y67ZJuM
hXYM4pkMslSTRhjL7cZ/vaiuhRcML7I2TZQ2tpVpngOQydYiR1LDt/fGVWBAVknw
kiIWkbWkgHeM2QeDR9Ub+cvewBViuM+7jemwMx8PvPX2/MZ8bdTdR+Q1FCS0G5QQ
3Doj4/imwIiE9PGyU6BrIaXELY9JOr3JB67DJ3rP7nR6Jq7e1jISPih0xMypU4Vp
j8W0foJ0yTjPcNAe3UngNaR4Xuq6QPvhD99/zxA3+Bpta5QGYk2EoT/yhBaWn08y
3A6/jfRR76tRUngjdBQWZ4kfcnZ1NhaQw2iBd8l4Bvx6pQomGVr0caoRL9F5mUfv
6ZY4XD8VoZ+vF9Dum/tpWsub5U896JC/a6T+8iWkTQFQlvV7w8aDYfOMyB01q8h/
I64yrDsUkPjvoc7vU7E521yULOzno6ZVz2U0aWogyCxuny+NvbtgXbXxYZVTb7LM
kdN0cf8S4upErWcyNo9hvWwa8/VbDvDdOTuHrAsnGU1lepIPFKoe9nGuDWFP6TEo
S4F7cEpBBGYQ1u6ElGkXK+MtEAUxRAbRiYahEQr08cqEFxcIhhgFrUpQTdHRSeD4
WGQod/GdXuEpq6qNgn1JedfE+wDE/CFYzqylvKm5FndxSrDFC20ulkxKtsBgtxm/
SXdyMI/bvyr099s2OA2dGroqo7wLFKDV7DH0SB4piaUr1JN7bAIUFN2f+Ws1R+kq
AmsrUmBOcIqNPAQI/lbczfpxgH14Dkx7DTaJEe/4dw42fd2YpwFQtYGqFPhI+RZb
rJkyrdEs8m49qiHAWHP7ux6HTuEFAZllIvAiBzGAaQSBlmO/ZTD21sRvhrE0MMOl
AOLtzG0UgYTRN7XqGLKJtvYff04Do4saJwRpvF7yRQWPYp7gmj0ZgjowA8kfMV2E
s+tmYX1DtZsTxO1WTKgRV5DLwHA9v7uBwJwsCdJbRVSY8j9KVuV/pFZZbg5O5UM1
RW0VH1h1YoCcDJKnwfCfteL3YVoguYoCRTpAz+ASpl3klAhhvCAERKGzYa4hyivV
4LxWrMEQI7OGg92yREb0b0Y+OkOPZ7JzW6ZilSuYDg4XCZI1LZaAUrzDcrylKQ4H
r0BocX1BSEfGgUMDoE0AJeoS2JXKs2/GP46Esy8hnfKCMGkdPXwEBpiYCwMt4cfp
LRSFn5L5DjGIIBT3oAv3eMhZRffiR+27PTJzL1cNN8eCiaaeHqqxjIw78c4dKeiR
S0nrsENk32WsCcL+67JlwryctpoCPNfUBrjZti+udvXOUBU9WfTrjaIwJpNsM38z
wc7Qi9eBBwcb0Mirgi14pm9l6nIzosaRncptiq4wKt0wDKvzc1BMjF/EWkxKydim
q0bL2QsgWpOgxS95+1gHpgPYx4DaXgeeYUWBKk2bB29FQEKgXIrcN5gJqqGV9+xL
p6S/pSE81qcptWCJG0YTfy6U1O6DZrBF7C/EdsLGim4SR7eqDY45wIeAJZcNd9XE
EINg/mAmZuzv7/ynbGopfbyqJGyX8VBTydZe8f7Oi45/gxnotxJ+EXIecg4ncXti
RK/wdxzVY/ZaLki4R6bwfQeHPb7bva7apV8TVA04UBLW3Ku9Frh+7UM24Bp+ZF1Z
HHQbC3FUKRKpb2bgFqq0Rzeb7MIlbhXzCTADYnaVW7O4USBobj8Xfo/WWDN+ZNJp
7+dosfTcNT0veTB8J1iz4kbGdFFiBbT47Q4+Biw75KuVUeLqshMM3kUDeIb+/A+I
iiXsga/0xU41HRULsp1ZwBzwx4j6peYhJXPBNLk+2HwyBe56FFcshe1WIskVZcrf
lJAK1fkUBjo3lw5JxRBedGJzpu0DfSxmeRCg8w7JPxJFl8eDZEpt4xUJcw//cdtF
0XOi6pWlgmiATRrPzvKwJMyA5Y2KZTRodM2dxypaVBPPq3eOV8hYkvcyiZ0K97/f
xiWMIm4rDQcVO2Ku57l3NID7nMdOjbDKS+I2p/I5999kKg8FHniIRFinYixsxKZd
MXtLoTsu/nMhwPEbHCppS8SFSgruJ2qJjE19DqfkEwrK6yFxpt8eNNKnwYBhDn0p
WDIbm1/iFEuyYiaKcgy01Jg5SSaIPd/3fG5FzUYKeKB53QGzQFyF/0GE8xVlbYUL
q9uRe+kqfGFM3r5uypxIM+gl6hptCMMx0fDfaPbi9yr79CvAZ3UJMZwEL658VVk+
+OCVWUW0S0A/z2/YtpuPAYrcIRriy0oU1uL9sU3Xbk6bbHhshFPLHW1k0204abE6
kkubyWbZ/8ll5gogjhXsJBt0+fDx4SnNToeK8R/BYDDx+kLStzv4/hqHcC3+Rw4Y
JsGpDrpy6+n+6YCEYlJa0q8BCcNlrWLPhab2jYa+8Ajk/yv0tuPhr2tM3S2Gm4uU
qwAK2A+2SPYH9d9+OolYisETL/zcXKOBVfB+sBjQb89GLn+eE1vlcdq9zBNvPxIF
S4cBS+5LB1QjHcq/TTNWT8XYE5xiGmg2Zm45WqX3CdQc1vhZWysGm+4ywhhZkKc7
JKPDo3olH99EuRQ1gamChqTcNbw6tCqhengMJHpoNUlP/KvSWEFKFfIjiyzRA3lu
1vy6O6CQi676DmnmpAIctMb3tdRKbu5cF0zGEzz2cN4rwh9Ac9nB7dVLIptx6TE1
z6CbCzGwcRzaXpRhch6iNieO57POnJ+LutdOa6NXv8cE0Ha3ehgp9dzYdQjKawR6
KpTVSj/7LPblB91Bt7g7/tPDwBVSFI1sSCRr0oggtMns3+UQhi2w9rtV+G3ArYO1
A1y8rW7dkovr7IqjfS2GDbAArgiAulAJSUmZnl9RmwZaJr8rMcqiLsSpZ9inMXsY
o4fhIEVpOhlOnvacVeit73DpiccphL7vX9lW3angmWYBf04eznTmvXvTqwmgN4GY
yr3UTkn7Y2MK2fFgdeU/NYCVf1g3t7Qg7HiLRFdF88Zu/fH9tALY6zbYsxQGnnvM
o3pdfbLSHWuzKDNwRvvs6/lXhnJMdpm5BkSHSmPZ/EkR9UbxxaWhRXEwe9HwQp4t
5or9dcEuzQe8DoSO6Kcx6zkJXdOxfAcMY7VjrD1mLoFmfCN+o9YInzTyO7x/bJ9z
1J2KgZ13UZdfYTL+kmKFHhHoCIiODnMxpkHF1NC2tJ9m85BOgD+O05LUuquwkrVg
O+9EJf1IFo6JijPQ+KEa1zEA4Ikgtzy3jCxRrltJbjVXKlNam78ZO8afr4t1X405
yu/B8KS0hp/u9cS6dDZ9g+nBYKPBZzLuqgHYdH+avYvZdSEuVfRuP6u2+6sxOgID
poB+v1Jj0a+Ec8Sk8at9teJhiPk46ZZFKGrJuBnt6bWccghriuTuNo5qGZ+gZEWU
oW1+tZ7aTGmU566Voc/iB9dkxSecEscejEALCKo65T5gvXq80GZk0dnlKXuAqC/P
PjK0fS2NuP4Szj2OT/EXZMAf3eDXNKfky0cHDvDiOpxPmqKapoOTbTavTmV2KiOH
tYIaGpgsOMdLk+3gi8LNQT51FE2u5zD3QQuiXZuFz3b/sSXCGjGEmw9HQDCBJY6z
rfwFQx7Kygj9OXG9UZYKLVCzqYR849QjOz0j2x5mYPVd+pSAyH9ivyorAummKTmm
P2atCChJvgj6qOofLHrPVX9XmCtmm51ide7eWZtYlqaDNJzYGI+wosNCUlmehA/q
eW6u/Aw2UFUmsFfZOxoKHS9ZfCKsXJIU2DRoizypaxq3wIsJbMNZlX3+PbeTUXkI
jCewzP2NF82X/UaUK5iBHlz7vdAA5lyRiCPniZpqZRzLzrx0pThaNNFKzCFNUfMz
w3VfJAJIutWSCQPuUWSbJfbHM1UMZ/jGLZg+xiLUj7nkWduUmi3ZOHuFni3bOEb9
HWGqP/41j+/l6XjHNE4oXdJQZMcGIYP2F0bnP+35Q1GmbQYSGc61TWs+mWPVpsZF
HuXMzlPQfjSqSnEDZPooDM8wVdZ+hmAaG+f/EmmwzinjJNuPl0abaEkx1UYq2FKY
ar4ILY6SlvekjuuEipjtdrwDBVEiajK3OXRi2rkyeO4iZn4KuUy/n5Y/IsKvhTE5
VeOeCAogf95Y5P8VZlyG/IwC/LIV9a63RNbTIrT8akVJo+bO2gtm1pO95wGlW0I7
3/i2oosE5ALYdLBaxNO2aHrS+X9WbRzhIANW9Lj3u/W8vJM8TqrZ1Qu20ngm3H7u
imHoXaXfvLEFfxw/vhjLapHGrWCXs0Xxev42GmSZOXfwXxQ8AaIcCasmVg7Oss69
TIub1ObN6BNh32uiZ2+vRVx9VwKoYS+DRJ78t3V6scUzh0CTVhQn0fMMvIrcb3/5
vXKLtpZmrNtlTK6lR4BvSszPKFiKMT6ZoCHTsJEguv2o1zSSrJ0buFBdjqWpGsR9
pGfMZ1+HNfA8qVvHR2Gzn2Nh5i7M3hS3udQM8mb2E2DbrrMZdOrJpW+xm9/uqDss
PXVST6CjcFbgfXF+4CGM9Aj7Od5QfgI+5brHMAGird0vx6P2AVHolRT0LkHsLdEJ
W8tl6yYTUKSS7NPtkis4FHZVRbIJd2zFh0f+f1X3V+HGXyVw4y+zUTdlr9aBim0i
mjEgUxxEJxbC8b8n6xwikZ+244u0HSO3owXCeRiUuHXCw1oiv9qw2V0tzAwq76PC
RMeZSk+v4AsEITZSczdFLHmBnPA2H6nXH0WjJVjdy1mVI6dte0XCnumWG0XMSQ5y
ibFuCOAfRL2B7cSBVXFsN5YxFurcXSCYPjkag5P/6jP5vRy8YKjp3EPXwXR1uchC
3IlAw9F8ncRMHXSRTqfhdI84L3Ltunw8phr86d7v6a4IvQfWYYS2FqG0aqA1Q3xH
0BxWD8NK68N77GKILvxcM3hu09X2j3S1scgx4VynGJuA0Q+8R07+Y1/xfDB4+r3Z
GcsbNTYnBGMPfIEeJI6iMdGR1Ys2W357JJeH8054dxfMkO5gHCrJ4WqBl+CBA8iv
tVLII1VSv/1QO9pk0gEixYvM1z4kGx+9iZraYZqkyFIt2mVgLbvJbHPHXAy5LotT
nojktOMoyiWxo1Y1Xy4pkSM5cvCrDQW8xoOES5TVYikvyNsJhJaNaMcm0aeB7/LZ
pAB+4ex961J3y7Gxf7TEnUEUXtvF1CIrGVLTxNI1t8Z020E/pt1N7auV5LHbOcKd
+MzdaiDVtaCLEojtAZpPWZ+WCxIvsFOr7HigE7n0UKsJitOms/LFKj8H2r5G4Sn/
1W/G8wByEBV3KjoCerhCGCSLwngbgvHR1Vokeu1QKKzsXqvpDpuG+7XdYGeXir2i
jIkWhQEiRQb8/PRdK05feCmX/ap7O8wb2YrcWcdvzIZaQJE0+D8g0gmXuq7sxaXu
LOEm1ZVzL3ST1EaHWN5GjVEwyPyTNGr8qC805Iac12Mt7IpYM+KuPveLk0+8aey4
Evi5rHkoYKO9mCgENT0WHz/d8FWJRXCdMsQ4L8BghTAwOm4iBmXTsntw7Y66Sa4T
tIK8UrXs8WzdQzBAxUIETGk/RValwsF6UbB+cX89Dvt5WmoqxgkHiwKpu0tvt7VR
7FZEgV2Qt/HlmQZR9cBt0YCqPiwg+CuocuaYxTTpbVn1bogETxrPryp0YKsRNxBg
IkgIFc0wcPSsRPDlECbmFqLwuE4zOs6HzL3h/f5h5djDHRSaMn1ZtOr/7n/Ec5aD
1rG47mmQITnY5AsvYjUN+Gd2NdgLalfW4Fvy7cSItB62Z4d6jLEQnPyaFHN/43ry
2pbODWu6WV/j7fzwFQvcM4dsCpIvknc6N/fPi0ksVXdvoyMKqw0cp+jNerPV8/BE
7PQ/xXPY8nQY2Z9MdwaHQcaD4IDXQnstjDlGZuEmwmdhL2WTL26//4I0vrEcutdb
ssMQgle8ybrf4A082NqhGuGmx9LXKzR/dhrri3Bzz6YM/aAUTIrLc6lB6EzhTZjF
NcEzIdXBxULv2KPr7wBWEaIAoBJc6xcn5P7/3fIELKZ4qbFKmMga5RlZD5rJ+Wp0
jnFbW+0tUG8wGYuRzjWCH7nJpLaeoHF/ZoQZbXcUDC4P4GvbjYuMlI1jkE1hEHlW
ITcn57mbaiQXXomTeh+/9qQmlLv/q4iLjfTcNPUjCvK9lNtbU9RMNiIrq10PmEmD
QmW3AGqE5TFXhyZuUo6xZnMYl2vrZtggUXinzjDUejQKID6f0f5h7p1ZkX/v37pD
zcwrjTRovu8TObDl83aknQw4o6VihbwbdajN343DDo7Dk4bdnp5HWqtKAkXMnjka
BWa5cZ8Ik+B4LojbdQpiT2muUoepcN37gJ6/roVjuhtBohIf2zeul1aSzKdjHtUN
1hq44VdMLcJMaLYMm4sfysS8As6Ykerm77SWlNk9tswKZT3GXFhuD3ZEUuoeqywc
KvYdLg/TUySlmAKQjcRvXeezlUYyFvvk8D5pvUm/62m4wh5zFjjQQbrg/Jc/Eq+T
tz0xmDFi/eKT4k8jUwlvyGVXMTDjBoNTCxGNIB4qmJP8wKwQATkIQzK1UW9/7rbk
Kzwj1fGglWE7O8N+kXpltm4gy14uck6m+4abKYqMVrgpH3QLqijNUzKw7gqgZG0L
W6Hzmtdyq2RtLqyQUYmJqAAKeckaXD2ZleC9Z3heTA39Rh5UEA3CJLN/QtUW+g6I
YuYenvYLN0/q7GE3YKjkX4npge/vdgBwzRhgPem9Vv94ML/lSRv5YD780Bcb7fth
1lUrjEkSouwSk+VqqPfLFuCopGoo8ge+lljnfCFLyL4rnEwvFgl3bWIsXwXbO2G+
LYQDjMIWd90I8pEKH68MUfLIpU7YPY3t+l02/vbqqZueupUan3yapWxVVZrV1yp5
camffgafPaAvYgbTecanTlHNTN75qbfNX+egzVp7fNGPxqzAuFSoPeqZ9GtIJdtS
7pXXrBWTofP5EmOmRYP9EAg0PY8h649O2CtDpa6mynwdtBYJB5Oe/ZJFeRMwOJWe
damF4W4RDZWIWspRsznuFPUszJjqCQXrZDnfgrt+d7YXt4lnQERbM/YAHcT/tO2X
FH/Vm/ygwjzvVwAix3BwWvi5ITsynuZWggmBd+e5zI34HXcRxrSKs4hDm0JMvRPy
IltmsayTIfml1haHuAkITaPJJ032e8Jv4J8Syw0wX2dJjEPBiX/eiQTFOAR43knv
XcfEtP+OFzkN7HE04nICWbVgdwUVEGeEKm2k+36c8CPEJ3wRnShf+I6JZGVSkaoU
QqIEZwnkju9IMYKvAh6lnflJgfkeg4+t2jt5K00RSCfZnaKKMa9YpLaZt4eSGho9
kh2bash0GNtgTa8izO4OgK+86TiGjYhyngl/3D+Yrwywa4uIzi+7Lv1ZEFQ9dhSv
1pvU0DIvpBh4fBvUGkGLI6HQW6IZI83fczWNmZ0b2OwtQK6YtYRKCYEOHoIBEvE9
yNs4YE3uWdk5VXM0TYbr5ClLWB6HbXgOjiNaTTZD2p0cYlTJlk1d5okJkZZ1ES/O
btEwP1UcEn/l02tUgoamln3rbsM+xnVe+hvVRJ8E1jYtvDSAkj+YjUqmR+K52QNO
rPrtWJejcfmq+J1WfGlaHNVots64FEcmESczQc2vW24yooQh6qBfr/w1UR0sD3Nr
l46HnEtrQGrL62XbG2YVMWGuZAn7uzxLtBN4flIMgonvUZ0ZAFlCSWNyQRNbqh7+
WGn1eIsuIKPQhDX8HdluzZz/U156YAzVBiriEC3kB62smtkM8M4l475qODbyyFX3
GS5klZ2JbfHlj+ZJX6XC3wCjoQB/0zDUS36zDLvvWf3Sx6ktJsS8Pxkonc6AE4YF
q6rD8nUb45f+8Y7I+7uucnLoVPDLLlHLEx04WMUbTCqL3NGFw8pqEYTLjIDmn9ij
8tI5lU2fxH+B6JDmr2aa1LfBavafIM0NybXIsow8VBneuD1UQrDckkH7mkzlRsoM
KyxAsmLki0d+2+W2he5BkZTe+ZnYbzxrVfps/5UkQSxYmw0run4nbcha8R48FFL8
GM6t3ding6ocgPueF5IKY0YWPBys7uhOouMcR4lFPMmLdwHxbBiofSD9TbzC5ezu
Qf0CIfqfV5XTkWYqHb+RXh39meyaw+TfIG0FGioMltDSZa8bGhbXLAkDnAQldgs8
OuvgmkjiVp0qFNvCyWWJ+Nyzb7bXrhYBO6bR5zfGkCxAAaNGeyvUmObam01yCPiP
0Npa3bcrWkBGTNREiYH9dtuXlG/ZykwhGlKozs3eyYr3NZXo+X3cYZMfnjgJK2tr
KeethweFQXzhInCYe3QbLuZvGj+NxQap4aNr4lG4Lzxd2hRhogpEPijuAIGreoAf
+IMU0bXWqT6zkEFRpgmkpX8UBl6tBBkyAohhPWUB9fwxqIXvF4JXF0jed6b7MtlG
ZqNUfXQKkb/H0hJ6a3shx9XckZvFpiA8qbdWJoY3E9xJD3WwLmFP2KmHr5onj/ke
zm8SOghyOXVdWJSg7jaAtjT97qmeHfEgwD/H5d1xs13ER/b+5+mIXYJLTexVDDlC
4llpbyQM5b30udjNnb8JARzqdyZZrSjQKRqhU5BiBDLf0hubXsFfaJ0R6y6CyRKm
jYsMH7zn+cGifa3K2ThrYWu3e8hF8hRI//FgLSqFeGuHzZRb9fRLFdyG7jaWeHgj
l3L1PnRCTYb6DJms37u1lSwGyYz80Bs3OQ7DKAwXqQrZjfDsWcgXobFyN0XAVWS8
dMCw5xs2WPwaXZ1w2Q1TqvigCXYZo2HpI8GPdOe+7xP6NIURDoRqulkuEKqWLBvZ
nDNOJmIrnqbKmZPK1UDZANhhBoEhjbG3Ws3zyYxgCgw3bMCSktrj6L6ToKJwV06r
m/b9ka0j1kDuKEUpLSL8mFS0MrbT8fZ7h6F253hG35gy1vgKoYjS4UQEC4bGkCef
sqJfsug3YQmNpHTbzCB8VUyeTjzGMOA2wBVwdooY6Xc4hPhhO1iPdPv4ciWg8adj
qim4Nc7P6+6BJeMWGCoD1RMNPa7+8o8tZj5rU6DKwUBiJ+p0LBvhrfOWcbdsRdg3
ub0O/qMnb1hDu2jScQUhY8ze6THq4xND5J5GsCTQeMlrwl1GiSu0+3Mbsa1VnGZu
TX1+DUHjfFXKRsL3zknmM2AzOth6XTmNkPAXudN2WqRkZqK1pYYN+rx8VS63e9Xo
sqq9OTs4cjYZYFs4/jkcf76pg8UttBwgmyT6i4iFSCqeHIjc5z75gkZc1IXzRa7h
9w/w+ChgO1B5f/RvIKFdrLeeA6pv2bmk2h2L50XigpfrKa5BFq1FCTuK/o1xW0Ro
yxgnVb0msouDk9GXGlbC4T2hKPyfNjz37xxFW4dv/7S0z1GWiYkOcAzPLbyjGBZU
i7Xn82vZnnwnL77VxGJNgMUwAh53FkggC0ckgemsiMjWEc52zgUaTWeMKcXbczOY
LByC3RAi3xHi6aJUwcVD7h03IYUezW4pqYdCdK8mUPEWk4SetmwqEGSOQ7zMcq+J
F66IXgkv4ea6RGuTmYlEom8FEwtmQN0YT3jcbKNM8QwPrb6dhZ4UxEEkPHGarC++
9D2RS36utocswa5dP+g647Zpu9h0q4BkPQu20tTg0uUW1BMbq68j28uDDrxF0Q+O
I1Ml2PcaYiauTpNXhfH0yjs6rpy7Zi19mYCFGUmilhsWkTqOLizu+zHUIghx9Ogk
OFMSqbq4+s8VTD/NSFsJh+HygKr35/J0/GSJa2cnHFY88gdzrseLCrB8ideXsJ7+
FGCqtl85bzqde95FDksAZ0UgQ6l+XCUCcJVN/aKvQVHctFaO8VnVxGCwQluEWkFS
BT1t4dxdZD67guH0/NUXUICPrI1pZPtx/0i2dRLHrnzqLW8TQy45JjfGQfd+j1vU
xn+Hrp3h12CRA6dtLIqXGYLVQACVsUmUs4RhHTlju3kEm7UQT5fiW4qnHO++yUrV
OsQpmNdr8SEUQUqR/yRODZ7SOAsSQlPBk0wK62A1KdAzbuBtOqtQSRTM17yOwgfP
25eIrx4UA1y4bRKzmemFBkcBTiTVqW6NnzdNHTlVgjUm4WGj6XPzEqQVrbYgy5Nl
/u/1J23Ffcvq7y5DGffly0rjyHC4eNVuN1tCf0XxZY7btMzfFdxB+efO07gAP4qM
E5nX2l5qVj1zz4HtQ1dVex9xqV5tsR33dYYot38cZnxyE1PmVK+OstEVjFsRF/fb
sZphSBB4lZc6YIWyKFfvzYcAQWl97gfDWjL/mmWWTGdwFBsZLWBwAPTx1zesbkHq
WgWNF0hVT66qN+cddp6MyIMUvi+URCBvOncM9XzsUvD2bVxxbjKzxXXGNJ5iPv0F
ruGAxsDtl6sv/VRCOzc6t0i6auRw1Hrnk7q4mu93pTfMHlxl0N3unifKBz0MG1yv
V0nVfqzNp1XRyiuu1vyyDxFg0K1K7Z/76T8fQrD+B8JmeDl5Q5yVWLjWRKLSjz2n
O1M4GvyZgMxV5AfvsGipGtAGiX+VITrlqahqdMNGjfvs34PtP30y+wG08v5qVmb2
TgIoHV2qxIn0jSPFJimZ+ey/gl7I0iIeiDHmmK/BSNZLzfGPKF9Pu1UYsk74X9eh
SLpKNsKActf0FzxXo36ERJv+WItSQy96cYPIWlabsuLNb856DFbFGponZzw9luwg
Y8Wk+a6mG+f+ihbMKyMk7UMkqH4vPgKt6HbT9lFw5vUUWPeXKOxcdLgxGyQUASBb
/S4oqA6wx2SOcsri4+l0vnLeA7iexzHOvUAGN8RW0MkDbncONzSSo44XAAEZK+NE
qOlsrR7EloG2tcFkeL1h9JxvDI+7jzzlJ+qpa8zk2FAwhLsSxAVPAt4vvi2VQpuL
If+SfODwIAUtVKNI97mCff/n5JL9+6AdvKmhwef1aL2Ul1bFBQtkixmhq/tJOA35
RFt8IjY0XNhTElfwBD4Pg8nksqAmDRs3vysQsXFkENh64e1IjyfFolPmO5fsR86q
Oq7JNAK9I3iHoQlSQlZq2c3hpOmU8E8ubZ+h5mTlBn5Zrc7KlbLVes0N+xY+lByv
5c6v+q2ifsOs3qGWxidMO+cqXnLJpfkfWZAYCXx//3Zjw3iTCw9z5GC8dn9A9HKF
A3bDmAwHX1D7ARCmDiaIwCVZFWVQUvIy7dJRLlk6vZ0fmk+CxSD7IHbUDAnDZD38
qPiAEX3WfVly/3wLBMfjH7hvLreoSe1+W5mbpDH/e21KsnOTuknV60OVqg6ZWTZ+
ndUZbNAsWDPvExXe/0yqxf5MSLjhLlvv4P/QLxUVyLo5ETO2Mz7NgUVr6ztFnPyl
4O43dCxp5ab7fvApim79GjN4SK+mQb4ZkQ2ZI8aaeikR/2EPP0JMi7si3KbI248L
F7kWn2rpQETjYGh7Hw8cgz9j6ML7Yoh5mkWWFjccz3Y/QVW1Z+FWGuejyLSBRpph
1gDd9NmrSKOPjNU79+LQ8Hl+EFityqa78gwZTnTgMELZwZ/TVv/7TiV3uc298Q0c
GJJ5aEIwCyL34YU6LQCyLOUN+jW3Lr+43FgT/sWdhl0qFpPKVXfNmU5Rr0aAj2BB
QK2wOp03fOjIsNdH8ZzNaQpY4tlVRxFilegNyUt+i2GrvNPYAzbsvSIcx32Q6YPx
fJVOPO7oEPN5r+pIq14/8/M+6h+vpBWRJOlFnyduK/632C3fXybKjbxQTzqQD3Vl
mK6zhHzOHC/nQhJwY77x1J8cZ5m9oDPqNdRtKYov4E+1Eg2fkvLORbB7Y4StwD34
kRm8/qrW46NbxB3fkmIqwV8LK6yKKYf3fx5h0dmMh6udIrH58RUwhAagrHPxt0t3
hq7K6A4Q5/1qWbo2GSELi7rUMhclNGtCMFQtSsCn61rzGDK/NAQJ6Y2hHdTPGC2I
kodrnQK+iN6gSNfpMQTqH29hMRgqqUyDJskqnuikN4TW7CWhzajmlPea0zCynaU4
jO+BXTfWnQdOcdzoKjqrsVTA6oUuXENgy7NxD07c2ZySLtu9IVJecJBYKbrwMd1f
1ovVUZeV2jAlBcpU1gCRW54fUR6yMMjOoxtgIQK3T3Iz/t09fK3UuSut77dA41nF
SlHkSDxdFwT2ExSZNb1GCmL6oPx+5b/r7FXqrAjtWFk4eh6jEjjWimhn2Ta049ls
8rxjlvn1yNcuCGFHtY9HedqjxepiPkJ+zXrKdaoJlnhhrHC/dgvi60wpe9JCxc7s
+8WRUEqQxSUd4+CSMTKKoxQazzMcVDdppBSmNxF2N18kD/1IdR7K8Df5ePGr7RY4
capt1XTT9XbjvplArYLkqkCfUHLLSpJ3EQYKWJcoYk29OVWBr2xJqDjfjox5Q/nT
vktJuM759dQMfxFE+7pG8FDLCbyK1HRLDQjbNKBIgfwzb7r/CdmDEKJucRmg2DPT
bNEQ2kIbGquGLs0zHzdExELYRnH7B3CDmegBnr6p8Ova46hOKNR2Ojr9u2ZCQize
vM2btlOEtb2mZAPOAbY/fY1O1i1g1jnyi7ietiZhXLg025yqTBAJbZ+8qgnrisAS
Wdak7EL7HGuh0RZoKnBl6C6lCD+SbbdL2Kb638uJlXIvvC036ypS6FW4qFYRCbNe
/KQ2LrnziPOAisP6n31Q7ujZKsZjyO3MAre32z1AgG+iZ2UxDCaixGSV0HHZSKZU
1GKkx9RZkcJ7K4Xerpd8Y7oLDAB50DBcLJ6f0NmGdoJ7vMHmgBSkjgD4XcBvNqsl
EmP3vy5IbMr7egvuWnIzutiv/oHMOoYuII5fy3ScQteoMYjG8cW5dnOxTtvM7N0j
vfin6dqIq7rwKxwgt8up/pT2Sqcn310/PYmD/rEUl1dlGWUKECPpfDaqA16pGuNy
eReS1QMXBjbCnnIGd0nEmdplTlGKNMIh1vEhS7jMY5JWHa2OzaF4/izQKIQ3Mo7k
KZ1COEf6RJSwdr1x71aUFge95fgf5NBAH8q1I7bLxulBosbt41waCURny7NHyilm
9KXaqzSJ3hIZOkpvoKKfUUeH16ZhJJs6Vrc017R9bvqCgGqQK9D8Uq1+FjOuyaNv
zgwelDKFmzkqwkTr1yhiXAAobyvsbMaTJHKQ/RdyAXHidysOIZLG7i0E1PfAdOEJ
IWl3UnaTr1DJZw3Apm/qVuu8hxYqbQy3JkNLnPOxoHirgKMGLteP/lx0SFRiMhZm
7ytemr3vqKjr3kWtvlVerawflYdCuYxUOz5fAdFnCH3O/Rf3inDXpjfg0wNgbI47
MHBZ78gbKcoySVgpLUYSxIDEVfIBPSTXO7D7kervS4ZG/J0GieKA0rK71kL7pamL
Qq8lRENANksdZ6KGUGq/ILLDsEogqjy1r7mlzBC0Cubd8Om5InXgKW1xmLcWabCh
o1eQhrZqDy6o8i3EzzZ1VUuI46nJ40eh73fnkcOev9IJueZl3Ay7UbrMmJaJbKUB
BB/1PmAnkAxNKY6m9jKVzeIXHmJrPdUSOCCfH/QBcwexxQTEunFP4rBGCnEwP5X8
hHDtJYDDKquAldjpfz1pXVchVmQSIHXAKl9Dxnx0gtKnGnWra8iOr4MdDnHFETl8
AbmHlm3kK8A7wZCOd537rjTDeEOIO+veAm0Yl5aZMN5ipGZQ6WULQrxVPnNQoHME
2RD28tTzkHGmOW7LUySinLAnyF7BMuX8ZpqkBABArUxfKfhb/KbtVySzJ7Eev2OT
CyvM3d3T6eCfQPIWj4+rSWxrEy4ZzIWC2z8spgf01H/plIV+d8PUcT6y058uvdVH
XSgWWS+DHvixDUvrCG2aE+TtnmgNtDFN+1pgrj6g2oNDAddYmxNM/DjV2d5glu5I
rJszsGxMLWPE/UBf5w1D0DD4fV+MUWue0Q2M2CsBvooXEaXpo67+l+UVUOrXPAgR
FBNIt+WqOAnyxEkBhibZB0o05WNhXjQsIQybTTRqybm0FRr+N636moT7qdSsz/6v
A+1yeEei4p2WBWprdghZUjirS6444fJEMuJv82vw2FuM0CRjf0Iovr+PMR823ErK
+witQ/bdI3hH5aNdzkKYVw8/BjIaoqZ3aeS8wDIdvVCQUO8zxXD7lwJrfvJMUogU
kaZGFM7WeZIBTalvyarTgw06IpWobfb/w9wzQQ8LZpuwelCZHWiNugakFA0Le5jA
K+y1kv5/Xt6VutCBzh7KW7o8fcoOfMy/jYRkkU0ZY2Kzbtul6JBd+Q8J20ew4vVq
iTZeaSQkZGyuHzMuWlFd8JlnNC6TjZD8+2zNFLnvXXigdz08z/JmwrP7+ynDGmZr
VchCLBelZIRljnu0ccMqeNuX6jtsCc/OJ5fz4zqCSgtDGkcTNY7GiD/F0HNox/NE
cFX4/Ua9oEjOp6ULKXtLodS7o74A8cSSfEYiNE5GDgfb39jPv3SrHxyQw+Jmq8rf
S92NokAhZzCdRBT6okgg1N/cT/3mxYK3mJGA2WMiZX7A5L1hIyChgYvJ+Oep6DpZ
bsBekzNxgj5ATky/TMmouxIT4eNUuzbH/zN3Y/7nOXwANn4FTKpJnQ4Tmp9cQqOK
3FWVKTA6sWqczFlSy9mMpUsSptnj/1NHX6/X78WZsWW+zhtGj1UzZ5xLrjih5kyl
+jD1pSBjodjrm5hSjQ1ZsaXtBJZmMnuno2NmmUXEDBceS4AXFWnGttWh0IpDP9GH
/rc7LNZi1jkFeAeHLk0uZ/iwLmgsuwEyvE55WE0FzOFr0eA/xUfSfo8suDhEhwhr
5qx9zIEGGJRd57dDjN1zAjViZIZo3pqfATi94u0Wa+b+5QftxEiVDltJutC9UuXS
bPkuH0rA4nNKOXTYO7PRWkFYHQy7Vt6yw3uL48bJA86KYKuNtCmUvyw0RWEsq6ce
5jDVQItLq7v2hFD9ah4pElvXdAJROMdHE6p/dXntw3RqhMJxBacOuuRBRtzR4TPr
892tv8AJNeGJwdzdlNNHWloD+oFSLQp0bp62VKv/fSzSoJWTu3plzzeLuHCoEpuB
HI0O8qFHgmJyo+fYRkmSY8e9d3Pbeef9qShd6/bvaUBuYggDB6LM/M6OzF20TRQx
IGx9zFKHjq9Keq3r79jROZ+N5IqR91KlsHA0ArOHao0w0Mw4lXAkpuHlxQqIpdHd
3vgWLNK0aIi/RvqcTFksKGO2gBISzkp2tMHKL4alS64l/elva52KX51k5hX1mBdp
I07OTdSDimCl6PSr588SVjAFxBN1aldj3kvTErgBvmzgBl7pdGgj2p0k+KgAslr3
th3skW9AlVLB1zCl2cwzdBTsG4M7i5SBfPbr+ah2D1tALaWZE4UkRAlZ1kYt5ivv
v1Mvv3WwwYQniPW+TBgUyyzj1k0o3BB4pIka7Ei3VJCqLOHC4XxtF3JtArlJPFFV
ZB13OF+3N2XDG1KbMKyzIuQJ1liFc6FqQTeLW3y6cwIzqjiPzEjmuAwo7YxqzG+y
h0oJBW0UNXL9JTVd0+HdtO8aCb644wY3aD2bza3qjvTiRE5AZmDMXR3HamGPsV3s
0Xxzb04FaE/hMALlr01TGon6g7mC/8RURINH247pfhpANqmv/qdDB2372LskR1aJ
XUsCTxr8+/a9O3te6/jbEUfJYYG8PG+IJaukokjI7Al+m+RtV5/BdcN5T0i+5nkf
whk1erOdnHYx7aTE2BMEjidanF1HA89AhT9MXxwU3TPdl9SCY3jcamIaa+LSsAO0
jetP7IPrOSlykZsP1qLOBJEzFIaKWSbVOPT0Vwf6Cpnq0tL6++5RpnkssM9q/xRR
OUEnKZuKoSdSFnNkWWuy36X0bOn3ZrOctnZm5dN8b2I+ZOuzBGd9WZyFECoKq1Vh
OJGAqfL66hUtzTwz3LuSSq8ZYIQUCW7hHCrBcq6aP1gld6HOftlI5V7jhMyhld6V
olb3MV7556R7c6LEG72Y17LW2mkI73gpnISYA2WuAb2mNYKsg68jzaOC2e+0hbWJ
HDgShXDedd/P+dYsqGYhPmUdVDoHA59ViPOZMyBoQuQwz4IGypdFjzcFYJWabGol
QuLQWcjD4G6K8VpzD1lrdT2yZM6YhdiXIZ9kaelWN0Bz25awyWLxEQvwL6hpl9Eh
Tz4PfY89iEzwCvbmjmG0WrWTAbSOhzuMzq+D9QmyBEbRHMU6N3wRm1OdbzCh+AUJ
/a/5uAmaXGceL5ReN8Kcv7epm8SAmPEYMYYnE99kUn54aiZ4n+KgDsLZLY8cVDsu
7qg4IVo+jWm9XXbneORKUXYu8eO8wigg68cgN37ZQRh1dV9dLksECOhLzOkQtaAN
4CchGzajp2lfssbEQSxOxnnZlH247fdiBWOkLByIq0TlSLSacrhsQF8rCM5V0/iY
gtg7ZjICtkwGPm6VNlYiFF/BOoNA8E1DuhTvQp/OEcMeV9CvHKrXpi2KS93JaczI
zx8g9C5OJDNGWdAN5UjjBNo1DtsNM4e4MO5jRFgJ1dZgucKMK9tXy0vkEKY7n2Jk
pCDRPgfMu9osV1ZMbDJOE43KLCBSDt1r2FyckdSkPd9RHtf3bCm13e4SsKri8aET
IRVv5+MYoZ+/Gr61l2nX7rZG7NtwHGl7c++EH2mYuJAPJXlpd5vj1mt6cMaG1evp
R12OVZhgrqT05TalI+D/wuZM2sPy6FPv08yYK1GUcZNyvi+0N642RK93+ITjVeRT
NWQDuFq/qWOuWbjwtamBrbV6hhkMwoJcWTq84gPPkSbu+w2VPv5KAlr2b5VY4pAi
FlNZOdl3pHyfgZRQRqSGeIWK7E/Qe+dFuT7M1ILozRyJXh0FgwOjxjEG6zzF9d4n
T431SZNcWRmPpKVUUaUWYguUGNMUH/i1bnWOcbWvcc8q+X8oVIC9fDb/HpRAIJUO
nqRQ4ghEdMj5I3R9P12lxr0GamMVBy4IwEJeci04jigj14ZYlEMOuu1N/JXlQePd
VkN1Seo6ba6U4xK0P7aCYKh1IFQPfcRAa9jxS2QiUj5e5G2OWvJncCJiSBmCd2Hq
EcmHylNi3PqbfBYaRDG0nZlccLq4qYUIElQxX7kKJxfoGcSHoeWVmA71IBGgVAvz
Tqu8uUKLGisfeqwccNYGVu3MLlBz68C9sWutrkYvl4AEB1k9RAhIjmrSyuWEjqbJ
oSGB7toJy0pjAkrGwQuIJvggrWBIrwdmzeLpsxMUjNh9IAsq7lB89okq42/Up4C5
fJie3FyH7VwDQhSzu2gkGmbr0HhxwtirW5tEdtZyu73xq5TuOnCDKEnIUA0mh2h+
bodATg6M6tL/o+jvdniL74HX/f9+bzTCAv/ylsf/LlN/NFHKfMwucYEXE2Ad0+up
ZIgKTpWQRbgrSpleq1gStXN7gMaDdYTPS/Y5eVcn8ZhJ0bcenyv9MS2YPFBdvong
bOWpeHdbwaCxGkZkq45TDQWHecc/NW+9bAl8I+jm5UqB/+78o3x5tKNLwYDhwc5r
KKMhhe4QXEVWe3Wetm5/acgkoTyAu8WQ3JhgKCwEBGoksyA5iXL5Op/OQJpJFGfA
OuY0sPF946P6YduYpp9PxZZG6DmViI28YH/1aXeM92VDyitcWXfCbTLd+BuW1Tqj
ORIDNq6DONCq8VrV9OAIr4QM/GP9wEPKxzFnAMsY36/MlYAfpHRyZoRNshRfKX1Y
XoAWYDfMT/fnWyb0qJY16HuN0F9jZPibDUHp7QPuRRtdjrVyyBDEoKuHwY73uNvY
siMpkE2CIvcHGOAZYOBI2Cupnb1Motp6eyeSqg3rzFC4PAbRSlj9YDYumJL+zrlA
lEIlS94Lehxb2EAbKb5YZrDQvZFPtnF0C/bj2QnCO5+NdPI99BUSaTtYAhwXI6Hx
tvOgPe9Eaw79SQ7lT6VS/kCNQ5zpHK4yxA7xHsAR85B7IdXV5zefmj4dYhCfI4hO
K6Qgrnu1VbEOn+gFGU0cW9h/Q9V4HkGd5OyOPo34+X1Z1FzDdrMuw4fBDOFYo7eO
rmnwkjclFN0534/Mw8QC3eXQEYCCXAiD0Jq5/p2WO4zZRDM+DWatXXZtyucOpv6m
D+bHlvGwyus4mLwGaXsfoLRPbaAFroGIJG94TqgmDwNYdNUXE8l7lcgqyYEoHKwP
nHxRid1iK/8MYstftAs5x+2ZuCyyN+0ce9DMUBwGlFZkvF7HGn6XpmpkKkOta4z5
p5Z4HlxvudE3cXzsq0NAJ0TVK6fORtAXw6WS+juwNVPTUh6B5G+/KVd+RpwVQJqq
H96rJtAHIRBj1xxBL3vZqNIqCDKybiDFCScSuS5EfqsIv6N1F8nQz1ORG2g0VjN0
5LBnU1PsVHw1II9SiyIxlz6KqQeCkIqqR0HwEiITaljc6gGxX0K482jjHab4FoWZ
Na4+merhQM3yTsvqY/+PaqzA1zO0rsS0dQW+q3BeJgYBwQ+HxgM880DWfCESK2fY
2HlotitcXvuAw+z8ax8W/W3WaUDE5c2EYPQZr4iL/uIRDtiPBZoDFGA2HR47+Ym9
8nh8DVogMWsIpk3YB84t+J+I8kcprufj4wWe1tkJ03xT0DVXHFki3Em8z/aT6XjF
3dcEbEhNTDI1pn12alje3hP25hDMQ5oeWDqcJT8NxemKPiF91F8JloMYiYo6kCW0
qolw+SDxklWwtwNfkyEaBtbQgTUX8uflIpnyvz8ATltx4YvDThkPiKikvWUDK3R1
HuVv5wFY02aUtnmJpidTsRP5etfmZSppQqE1amGwnpkXXVePr+v9/QuDNCDv7aEn
5SpZhgJLzddJB5xVCUxJcrwWO7lYuO9LRwMQGfTep6qUYFgQycJIZjoZtGoVcOZc
VvdA+s3i9LquaV+QORwmMWaU7L1q6H3iyoXGCHqZ+f7wmaog5mapnL7s4ciKf2xa
lierfQLHK5NwOW1dYGSPQmRrooEperqjQn/1xMd9QuRPaNOYpIeLR/nlGI6An1hT
vmBCtFEfirh37dyH+ya+qXVTG38rv8GsuUzsYWwZcG9Tr7M/J9C1dwR7tjWpe534
m/mr37eVGmnkrKXCQ/1d8gSmfwuWshHU8Ko5N3e7qzi82hQ4xLSmuyee5OKzViFA
qnUx8s/a9iKrjdDCTw55audTFoTKX21z/KEqxOlixBSSybXaVTfyki6R6XdbXULn
zAKBFyiVgEwcRg52kVl1nrkCmjUZjlXRazTFQGuCLTmdE4hrHQB6CLDrH28g7TFL
xM3qcd10n/0iBP0UrHaO5Zsc9XHsuxXD/EiL7u0rFUwE5oJaOkSC7VaCow2ty9JQ
ZLXLog2qFcTEPoiBh3wl8Ns4QcbJdfJzTZ1l9TzwMMZoqR8WoZcVBgJn2PA7mMqq
sQzzjHXL32KliVGODQ7UZVKVcfep/Cf2qE/XUWLH6G/LbxNzo0k05EuQ2C3HbtYM
mFZo2OPVnmt9NLDM9JxNmgBoTrHPCDC2QfuKiRLTZ5mgR/Dx/S/Gi+d8dbhtP5iA
yC6LNvHXAqCAzFrUK+rs4gsYNrdDOHDAc/6MK0Tzk21frfuYYF4lIaqkuk+dE4eb
hbWfgQJpTLxiOfwJmmDO2DVePsHRYz0V1u7fRvq8vz5fcZ3Cogq8CNZSymH0UEtn
GwkdxGKZYEeDJR2Lpy1X6ql9dpZ885wkH/UZeJ6M5AmkBweOEMxoFfsoIiVVADb4
1CR9K5ZzhLxJwKEEd/vFZvyTms7w55AD8Tb/Zy0iMzvUXcNEAyMf1BgXYT2UETbw
Nt/ltD/f/RPgHXrj8eEKQxVuB/SheHVpAn6xpZR/8rIlxWNhvDpLgYdMg5whOIdY
fpbgviwF6/v1QAMNZFbYphlHsHsucWjiPQKxbyvwIXxG3wHmaVE8CHx4kFd9T9Ud
wFdRh7SZkkD3MNkmk2rTWswzPG/rF6zK5zAvkUOXgKKQWW+PNcVGMK9iesiDV4Vj
kg2uyWwcOo2Gn9+k7rhFmckwOM9GaLgikThAdSs2/26SSHA9uZfqCfazJxWgrr5U
6CNhp0IkSDE5XNaBpcNVYU1CqnbFgGGCe/E1m0ffi3PlTR5RkShxPRY/RSlEmrav
fitWlJLFKP2d1hPgt/0R5o0nzFJUpzpi+08EVNbbkTQI3bmRqwtVJpOJrd7w6kq3
whd3WLe6/ifvClYKPim1dYMak8wyEZfNd2KhVQbj+eZVQJpoL+tJsGQpQ+eHhflX
Ah10C4BffjfSVXvUhR00EpmfoEF+oQSoS9x36OZBtK0T5RJYxgbn6ouWknJz0snF
8HeB92UkO7eoyqsS+9Sfu/EkhXgsJ81XQX7v5d5THAX6IkgdVNBfvTCPjhgrPNEf
M2rLxqc5icNJWOazwb9cABK3wJpE5NP977svf5WMaf0ET1CAUBbzovRu0/Ph1gT8
9fXA8DQc59rBNiSyFr9+H7LuhDWsiEFnvyQLxxhSZowX7unC7yvswtEhCsTAvIT2
dib0UAhai0eHlLOeELlFSu86lCCM57iGNs68oYHLV+buTOqf7jJyzpGRI7u4bAX5
gEFZVEXokpG102QgHZ6UfhLO9KR49LhinQ3YMf5+TF+KOo47nZC9a6KBSsKjwI7s
33BtDvK6q+L4idJLNTQ1RdYF2ZEtgnaVgfpBiLROct3rkcjdC7FDEIvqZnWqlL6N
HEzeI/CeMQZvgWNtCcs3wjiVVnu8cWzwUSl5nqcJyyZPsZToQemH8t+Eex6j/6L4
hojbL4V5NPEXAzDXIep4yry0DhdH/fbIawhyiQgWSRhylBF8I0SETxLTJpXzHalt
YtTotvzxDU61HLwb3Sfw/q+trLDkpUmPT2hwC7USSPAFlrMuIcvAQ2KwJXW/Zmrc
lJgwsETn101LkIEzjW4VprkCrxABUbQG3AlU5ZuQT07apHDQH4UnVOiElyj0QrSS
k3Oyz6YsOYNJxFt/HhjAJJ3t4LaJ3qgNcnSNKrM5zc3ZKtQnFdlOifwIFsRPdyGS
e3mq4koQAz78mX1j3TVphf07e/oXhRD+X7PRy96caGvBKxk4JDpHi99oOn50aDSf
LQ5JbE1bXQug8smVRjJjwVeQr33WiYgbseQeIpT2kmJLGf9RRNVAeV0Qd8kA6SPX
2eZIHaLKJ3fq2C/8J0zaZe/Cx9isaX44u0X7dxKzBVVexIg7leX9MYNp7gHpVrCc
aXWVThOz6neCTsAMggVxP7PdS+Ucw8U2WPfK3KeUBjMmAFHRCE76+BlcOxkSTQ6s
NPQcEjmJ0f+NlH4ufijKCmvOFnx91QWMdPhrjtBwImVNOVYzHfgRbcE12axbRvOZ
CHVQ14iDT4jx5gvvPwHxI0lyvwuBlaAaMAtEkdCBM2RsRV+u+3Cr317H2i0G19Ed
0lMKj6o6s4NSjNAJj5TJ7Aq+yN0sNgMPdxpg+YQRu/XW0d6B5eaY6GfCI9VySVD/
wUoXD4ulLHiNjnSgk5AnKUSJiKTeo6o8CGGhmewXgYdUfxbKRwuRI4a70ES+VyIN
GVZ3xpzwJyJ77q4GuCoaJeWMilaIfX1vk7U0oFiKe16XW5OlI6V5vlLXPpZsIaQi
XrcMbJV/3T3CTIWFMX8rOQSSFGTDR3CbwAuMvWBywpibe3T7Vjes54T9OJQBQMpN
0EQiNeXH6sMn7hh906hXQaEe4b50WgFjL9utzTsg/3+YX7UUGovmjSZkPXB8Epg/
FQ6BQVOsrQ8UHFJWm9q+yKt9xmJtOZ31dW0xid7ZaTUC8gp2wvAxA6BKPlH88kk9
h07xs105kMi8ZtSig8Einh7iKz+EkwSsYaxFIoXvHyU9NOzq6ojXu1azIWSuzdqL
ihRhdaMS2S/94M5P4F4d+rUh1hXthMn77VzS3SWZ8U1lMNcHLwTVirvTk/lUYwgj
Y0lrdc+JkAq8VX+l4h6vAD8Oo6+A7x4I6G9zhU944CIG+Rdrd1xKhvRHMZqYX8PN
4lLXP/Stbm+xsG4IXYws5Th8HRlh7A+eOV5NlJubKobIf+8URmPqG419oIHQcWn2
WZVVCxmOUcfzJjOdsmLvJTqjeBCqUI0LlW3TE0cOroWp/gk98A6QweI0xvOyguW2
BtZG4R4Qn1oCHmjS+5jnzcFv8GP1WyrjXgGbPsMeiFIboeoOR6PX24gIGKWPgTWM
mXKR5HsSXu7+NIgVrWKaKD5oTTzMNxP96UfdH8b8dCl7yC3TXmp4hgwc7ixLgaRW
mP48T6HH5CmbhI5OyPiAxqmL2G5ukWMIln4C//IYaFyDCpyaGRVakBeWXeAuaOzH
Py9jtSItyeZZzV8/vXbpOwd1MdxXardEc7xKQ1NF2FWny1jC7EyjoLhqfy5DOBJ6
3URyK6byOPTVWDlbGgUVKK8M9g+MhRLmDTR3MTPg8fDXGYUCRU3lYg6sk5xByWWq
3nWJJ9eHSXybfPiW363UYSxPbCrtSTU7dpX5M1rfB9aaEZqVqbx9wMsCpDFCL/nK
vV41BQtWcEfRAg1M7skS2/Qz0dKMkvXwlKIk4x5dzNqtfYyC7NpqQlSUzVBtF13X
mRQDwTYG5EJjNRmnZ2Xw6RNxDWo0bQhu5Z3G8uusRa6AhAL0MXrN5oVhPiSw9FTG
wUs24BwY6ZbgiOvBOA9JGsfQPhnMc5+529NtaMTxrmizv7g1E/c8KC9X+kWrFOUO
2TM5+MH272z1pIsHRWkN41sWSyAFneUvXDuiLoS80bGSF99H0AmTEuIhRt5zWUlu
SJOFmqjjfB2IDv/v9dMsjaUiKQTRFs0CryrxNv3Wep26LG5sSnjiiYB0B8u5/zLE
ECw7Qir1y6FEwROEYuv+hujxta8seUcHEWtZ8x5bqZlBVe+MqonMCQ3I4J3PdxL1
bsqRfmMu5LU5fgQfmP85oVZTjf+rgrDuwsL4O4g+WFuJiffdOSVIrP01081ksEvb
H9jHMrK2BWkpXbRGKInhAsFw/GwmvnWnp+UtanN8ZT1tK83NhMwF7LD1Dmit/kWg
nX7C9CyTdizJrM/QQ97zrqSCW31p1RTb2idaC/TAPTIBv/Ol/ixDdKqc0tpH835M
FG4StIBjERtLaAKikCwZAKqF20kedZziNVWOFfuuifFbAGMcN86GBMlmMAedEa8N
DbroyFglGft6XRr6EWxIeeg6UIAzaG6XJC5p1Tm8Yzu2L7nQYi81rbsiG9o1GehW
2OjwjtCvlbr/FRGNdTnsck6FU1WV/u6Nwo7iVa+RPqFEM1o3tUwMaeAtsAzDs1x0
4TWn3eO0uZhSydUFCbaq8zO5SriLgtwQ7GJcdaLZ01jXfdFjn2uBn45G7AMQuu18
+zy9SCg1iI30MShM2ten9e1zhRrnf1WK2SccMQSzpACCN7jmfJ0EIYl3gIWFKgly
7GzzNkE3VYMdzuxeIWvjbL6D2BRJAk3nRu9hgAKyAVPQYfi4loqvPvUcmYLlAK1l
34z9DXHvlTo9ECnUg+jPyRib/s5utwHPrJJ6tk1BYfQeuNNbfDdueQEJEoVOKvoR
5vhH5dt9POOyDW32zjYqpih8TeBttlIp8o3UOSy/y3wqHs6M5omBkuDNyeP7rchE
q2f8pbmvUMo1Vg/B3EErkHQhab0wKjT+UIq8zCHh6Om2xbughmqcXBSTEUaea3UN
hGqICbfS9gwKBCLlha9X6vWGidz1N/Bu8syjpD8HrrTUy9KzxtQHQLe1R8y1gwyW
Qg9+Y9pVDJbBBjM5gW7hXq7kGNVY3fN9txyiJBKCoecarNPWilij+Ifp+ROAPSub
5K63ON0Iy/ad02vBdlk6CG0ixfwFrCQw0aC9x4tLjldyuzYCx3ewBRHqyKhYwzV2
/ZDIyoOf2392nbC5lx09CvakeD2jjKIbGs7WeA+fU0Dkc9XbesRsljDybU39AUsR
Wky+HHzncEtDtZWX1uxUpjg2kdzjuEfca4wJFPrEYauKL14qFx0lB2IOAco2xybu
r8qVv/h/fgBSSOO/KSn/ZVZZg5BrzYvVAnEIMjdqy7IrH2Nzp4ffU6rZXo/oe7+T
PRWoL14taGVO/M+bbNITND/TyLERWvnCnVVJYiy7XGpJ0p/ne6nmc1yHBzbK1h8h
JOir72PE4KHlJBuxiPXsdwO30aQCnxDwqu//zrtiDzFGIwsjd3r7v5z0VcEpN1Er
KNWTuQJYdpDntAwbayfnXYOd0OzeGvg6n4/HmkTvS5i0GQCQfqmq/hzILL2Hwvrc
nPwlW7a3z2xaGiCg7kE17zjgNbFXWNHTDBSXaAUqldQv5H3uPjBRhbdGvcgfW3WT
kyRy0Xb+Or8eh2Pwg8Mm1XjOsngPc/qBZAB5CvEHEGJ1VbHQK99NV9LaLyogVvdn
AiTrUrpDANs+DJT/YUQNL+Srwv14czVYiBsufkAEH4Gq5W+lgNQoOVwwiyNwbBet
nTZWIcxGUCB459CtF7tyApVsQKDXOoXLZsOocozhpI0O7NUVqygAN0OEEurFuuIb
IqFe8l3i66JxjAfVNTxH7lQnu0PotU9rX9qAYJaCa6PmDsNK5SffhhLqlThAYEUM
Ra6Y3mdhlR/HN8EVQqxoFlYOuCRJa+ztSufDZQGe6vj301S1S1hiXy4RZY4huqzw
hJQtf95hrrZxa/I1DQPiwR4htMXkJwGWftOgFrx0X4nmZ0A1cim24mfICGsr8WyW
IC+xUSsTYpEQn8esbnWoQxVjzRcm8DI3QPMOkS8p6ihYDZSCIq8iTay/+pTfY394
v/nqBeEqMN6N9h6n6dbPWQOmijfvd6QTZWebkfSpW7BYf+/oJdKkMbbqxe8v/Wv7
gZyljJv+Sr0iZPRs2G8tLX2d7H9+7uizOGOTqAp561MEnnLPZzh4JEF5h1j7Th1U
X91raRp3+gNB5pkAhAsn0EDSxR1584vpHnFhC8AsWFbJCOwNQef0wnaeYAgWRiHy
6/qkaf/oh7nb1TiWrK06ijH8g4bWRL/f1ixJotNZ05JmQ41yTRbzBrmlHKTBBXIW
M8eeMBm6i1AZIjQu60v0tqIZwo7A8ebRrGvR1Jdrf21AqQPT98n3ytpy8+RfqMdE
KvVcdsbhGfZDHvGM1Pa1s5OFV1LyzH+VfMEzt2jfkxl6c8B1nw6fN/IGPRtps1eF
zz+s7ajB/Z4QDePN7+FTs1+oH4v/QX4oMVK+J3Oma1VkFkSNTwgldu5yTlxVqUTd
W84tW+NfO93QvmhjbqFrviZcGlSj0ij7qwwPkrvKrYwXi+cRrecSE4g8wm5tBund
GupcqX5jr4wcYMX06GwuFT3bRQ7PvbZ5yjmrz3Me3BwyHbwCPOCVY7r4Rv+K6hW/
kPi/7YlLUrCd1W136eVwIfa5cvnpkQ3r8UEsP+TzrbW0oVZvGNOX6XjXTkveQZjm
kw22aB5ezdAmSEeMf2QaBkNZG1bWMgbxYZ3LWeKX9QHVKl8oW1b38XKb9VJNX1Eb
Y0QbD+YzHXrUPYFc/6x8NVG+aeXvmwlg70he9tObMBifWpsXj9Ohd7x6utndLkyY
C5ZsH2zCNnIv6RLIuS2Snxx9kVcOc7iVPUS6OlDFUVj70zFOfOvQpvDVSwnwZZvg
ihBNmYJmDu3KQobbD/ctX4JWHQ1MIArB0OaVveNNZytWLe+Z0DMuWs4wsXr9Lg6W
pRBjYd5TZdLNSdvYpdRzgspRiqF8vZ0EgntyDB4TYRivCjvr/HDqHtnoK0YW1Noq
//PvonKUsWOciP14uO8q/oCOLN6ATzRjW3GRLBJchjOS58tTv01io59MCb38Zi+5
ONCqFIDAGsm8VUsAQvcM3cvjAr18KgHhXA+EfGV4ZRK/hQNBqSawFjIRB/v1eNSG
+hCYGCbJ84JuVAifb7XiVcvujvE4e50Kah4Mq+BIVeHOYtAOJxnPM4gA6MbK3jFC
a9O0xskFlAgpIDa5yWueR8YU4if2/d7Bco0pFh3IptJmUhtu0hDMf0bHOGpscO6X
ARuAP2N+3mAe3jByZplNm41gY5KnPWg30yUeL6TxJi34c92PulzO2VXND4fW9aKE
2Cbh1fu0Q1oHnZy+owHsZ3h2ZpltytjSlOIEUUASE1Fv2HMEWpFsLoTfmwNdsOdP
T71BA/s9ZJrCjdhvHVN8+mgktrGb2J+sMDmjM73f3OKOcAbSzhspZqTjsM/eUu5u
Q0iN3pmG/tE86Sd58z94oknQ1f3aOpICWClABh2v0pHlUEqTWQSbxm+43gZW57s+
Rs0i+ABwUbLWo7TsGx7ZUpa8J4Oi+Pi4vJR6DpfjMxsQ6EUJg4EqXuIzo7MHJJh9
fWUXnuwV8cSuG2GcgLk12e+qybmynP2zi+oktLfFMx0jTTuqGlArqAloOmX1UioA
9UVsodE77XAW2YraelEbmqPYI9AyCPig/vH+srlLTJYeHAT/kEEtJKZ7fuy/RZ1s
nB2A51NFVzF6w0HPR0MGFjYsJ8mZgHleHoVhL7Vxlb9QKpLaHv0Ys7OxXdP2916h
vf6xJcR1xUMc3PyjiwIPCHz+JzTUqoN+y4x5XLV4gPMybXNz3MGKhQ8QkMi88JPp
P3SQzSHFBiZD7wNKqQ3LXJ6L83i2kk37w7FaTv/OI+3yfnVKcH6ciL68bbnGPOEr
f04pAyUa6UpZ5NaxojF/MFzmBLTPu0oT45QjZqJE5xZ/3KQ3y3q5ldLD+BQk0lJ7
MNKPlcXzzYCDEfbHJpx/IBCljI/zB4EC91fA/UeBlf7kqSRrbfQ/we0cfrwRXCuj
/iLZBgDenMTQlpu10qE8HeV4KTMdEfkglhepvYwnwsQ8K9zI8+oBrJalbooYBRMq
LDBmnQykd0ka6HjhjLC2o3aafB1ce56uJ7akUY3YdH88IjWU6XTYY8sj4xBzdbFd
fr79lSMvqh6p+64Aj/kMpL1gwXWxP9lQ2G8BMNwhVPG9WxKbLlPugnUz81LF1KJw
WpCo62EzRXNcD8Ramxq8YNro6uDK4FasA5ezayxipl2HHMmG0k5tDXp9g9OeFaf+
CtNf0eZQa0iXKm30TA2lWVaU2iBLPWDqt+7UOEHgqj+qr8u5yHOOeoBunAd+RqFt
xsgmz5p9G5MWNTiP6bYppNguBWQ2I/3x+jZdPyAbK2bcDsL4uLgacds19gX1S7+O
knLA6kz+Gsb3NpGyCqI7rDSRQrldVLZbFuvV2qxPcXw/wRFyew2Rj1/qDyEYmcAH
BpI+AkMIxKBYgu1pQp92pSuXYEnooUjnXZ7QnAFZz2XBKgLETldUFb0TsA/ddj4m
dIGNHN1JvKa9iAYst5p36KKEnHYvaNA59JTwNuAeqajzGGye/AmYailg1hIYuIMQ
/ORUy9TwYqNjKMjkXH68ncGJD4TtPORt8el3uh+S75dR+bkM6cdwuwbLKkffkXzE
VZcd7EdhS8e8LKjqCjMzoBTTWrksUS77t8RcsL2e3sgNpJU8nUMOWXE6T0X0lBDP
COFg9jHkOEgCF+5uzqCloEh77Mn62oft3AI0/BJ24eDfOMdNIdx73e9LNDzo7MV5
V5vRLD+q+vB/41ojYmHw1H4WkEirxKvFyjpeKHKKQIGFj2vMJAKx7lA1QdBWlnpD
v4B8ZSs33hr0+T2wUAPQ6ljSZUR1CMeQW9MBahHuqA8mYaEWFFJxXAwrje1H3C1C
JuaQAHOqn3T+5RVatcWKom5pThdzp++srNNyoJLZ2UW5ncveEiGxIcV95f1YS1GN
vYtOgTXdvySEmNjxTv/8ZgZ7LiVb890ytqeQdvSpHD0EG71mIaDRF8l+6XO4Xv7r
DO9GL/Y5OyGduF9Juj8TRLudOAb+ICska3LlDw14H6P3Vcrq6VnjVdeKOdEw+O90
OmgilTADUyIu+OBpOXBTV4AQmp9jMExrPLOX6+VRL92xipHBYDcXDFUJ1H1HMNyk
fbX4L9rBdgSKa4v4wIO2bhQF1guq84v8WuSlNn1EEqLL04eY/idnWWVsjNfVb1LC
LZkRc1kOB+EL8joG5b48R67LXCVnE/po3afFLopcka+2E3GBy+gG7aKCPcEohZRV
qJy/QN6Qbok1MzZIMto+PgYeiV/gZadK9c15IsEw31r7zXttbiUVtg5ODD2w89g7
2U01qIJyUeGyB4uGVBaEHOAKYSPbkqoTLAyEylJYyy+emZIGHScI59tnUZ+jiyjA
WV3fYYqTOjG2VWaAzECb7y0yJLKBOYwU7wlGn6mPTLZpmFbZJJubN8/zST1J5t77
r83kGOu6HbJLans2hysZiRmy0okgWPAjzqFuga00/Qm7PMioH+cQeSIJ+vD6BBMz
ehfFQvFDvLM/m9vhzUC23T0r8PLX1Qoj+w5QY+eimELhgKb7hXG9uKoVtpGk3OfU
jm3qyt0EDRRsfZeJAfBh6cBVei5fu4ZmUffCKqyzOdwLy1JzTvYrkgCpB/142pfp
ixw88YlBDXkIHveyAnlhTK7lwenVbLjPF7zOcUyoh5bX2U0RhqxBzgC+wPPfae45
q6YnUFU1VS912U4Z8StdLSYxGuSK9WtZ/DBKP88vRIGPVaWOxbZFHIEJgKrNjzHJ
q7LmdEqOzMnfb09PnGGQG77HoFt3nYpD0KH/Xz5AWeBA8luAcClUpuYZEvAWBqoK
ba6Ce1dRGfHAcoXTRhSVZuuWyqVvP/DqZtrpb2KHdbxELo/771hzb1E1gZ4BZQF9
nA73u4GVErNmDz2NeRxlvzllP56/0lxIYbTGBruhms7gaOBO2FeLiHMNo0kj3a7W
B4OxT0mIyBEMpXv6xQauMQav7v3gdm2r1rCHZJNku7uGPRX8xm6NXEqeqFa5yZAI
SOSrjXDLdOPb94aQHvl81Ak30FVRoJmVo0es0fa/0riLQTAsoGFmPXaCRawevWrw
ZnuZHpniP339PhI7km6KyPXqXZwG/abHgmdX+/gNFqYP/r9kNrRw4QlOVyZGdxi8
F4yvl8wCDNwG1jnPfzaebmjmSA3syY7C7cWVud4+IR1DRcHg6m1AdbzArTNlmVQm
cU5z/SKeSakA0ZrIF2rpPhFUnfWqK+uxdYHRRFlJPlk+1x6/O3INnlLyEEsXhPzO
FJhltlm3AcBBH5GBPIXZ/iw7bHxIJ0FUjpZAQwYeOnbffTvOZMXyiiZwKOlISbge
OBv1Uzxmno/LDTXmB74ZIaIDrAdeD/fqQEG6eByHJQGdbcowu5i3dac/xoN8po08
1dDM72rWAyxLaQmA9CFfejSybq8USSC/WmJwdAuJssxzejc2Q8ST8qPhICBgWw7D
jBe6Wu4Cn/qRIEodeeEh0aKAIKUXRXf1+vLbD9RLstHhnpEPdgWkYDSxtMq9fmWU
ofozJ4gfpqKOAHsZMqfG7z3REvDriNKXtafcbOXppEbGAELQFQxChSDxvOdjoFvz
eEfFMhdDVtXshGooa7ZtkaloLxMxFFgw81lxn8T3cV7j/YEUvFrp+jm7vIb5A7kK
+curYOG3LMAn1H5hQe70CZnkN8WKUasDx4pB+2bXQvhS0kw0ifV1SDjPHIxW84VE
+TN7d7yHGBYeHRTN8M7CIKSbCXdAbean86A+4V9f8nZLKZ3RTOXmPKgEiXrmHq84
MWzpyAdR+RdzJEtVaTh4FRxCeka3EW27Tv/VH3pFiEnUVpxM5WR9ecgIPmDOML4T
Ea3g2b6j7PSWG53jbz93vYRN7bZrqRL4a3LC7nr9PhxOvQOFjTqE49yYnMJhPDq/
5JHvfXu8FGc8pABWOmxQZ5tZhy3xVfdUTKygeSNizTCS7P3PSlhMg/FCtPg+7kw0
cTTK8t2SLugKbRdj5JplgMBH23urGLeQzxSv0B03FodMpCKqpdhe+TOIRPHAtL6l
OobwHFKaSYcG+lR1zpfvX2VovxYXtg0HNQS6skSovbBgD62RW87rOyR9l7ot9+rV
qbWDsmDsrjzjvyGnsAAIj1u9Pfd1AfnUTFrYse1hG8sqgHU7+h9bwSVAZCyS1Bl1
U2Vaugu8s3GP8adnkTd1//lFDGY/PUl795lhbgDbDEQR/2o7mpSinziKjEB4p9wX
oflZNPRbDUlZtgrKRq3ngdcUX6gTqeSZHGiQjAusIKW6SZDRuvmCyj59eP3BaFUM
5qqiDqFth0CJUQSkW47EHWGmuBhdMtMzsiUKuUJbRaf6SwxH7fVdxEimFwslZlCM
52shJ9J7dQETB2x+xBiAwoWZZ6foHRpy3jqgQwi6nwTsyGpUvjPDhiPPqk5OUqWF
9UfP3+JynFHmnsdP8WjB+q479M4cO71p1YWBcfGfVsrMJ4pIwbgYAKw6fli496M1
ENOryI/Mj+UeGeEl6WI44rbpNxYMd+cSqlMfkBlk+dyjtb5/inltDbq68fEL1ybP
LDVzhO7oUWioBS95PrnxByk617MhaMiSuzJ8aDwwwDb7e5XR8KgVDAKbQhX2hDWD
rkLgXL969PfgcIo0FAuOYIncmWwxNKTmf1YJqjfRlE2bkGqGsRD07Lh7j3hycnkV
nZ7lpD09Thb8AW9WfBuMoONTTMfo2sI5COLWSOI3lRRUyvhX14RiNOImABuXDtcv
X0vulXL8QIjqLCdM5FMY/Neikem9yP3eQ2WQBj0Yaid6cuNu+2hk3lnP2xf7TS4C
mAwjmgg8FE7sSiauq7FBieKpMW9Vh0HaP9VxMCh2/3bjSMyGP/Cp1BtHWOP8PT7g
5Mi8dcn6uNkye78tKGMCboQR210lghGQt4O530tZ2ZSLsJtHI0G8TzF4Gvstu/uL
rFb85duWwosOGBOoIUvw+aDmoCHBy29L7SJvGRyWplY6rhXdFoiyctXs8aalRooK
0tfh4pE8Nwudd1b9bzPC1LHAK5lsKfzagxnEU0tvbWeZBxeQlhbYf4GF4OowVoHN
OVT1tZCFy9H4CZcuzmQZmXynyOr8yaXZKqLyXbPBICbikQJ7HURIVaKNXtGo5mN9
GkqoDRqbjt5E4maQMNHjqvDvBM8hF/oLX+KhxYLM7SC36mHZ5MIEO58hY/S94Fr3
lkX0zb273PIrzTlmd047AODTG+rQY0hwziFy6yLGPO7v7vmd+9axO0LPK8K+AXxO
d3QJy5WL1I/SziwbT8mVKdoKNsIcZFnDsQPOmqPqDiogassP89GLd6fCJbALi4EW
Lvl2QW7QoXNyPkAkELS6YHvyoXHl4vkaZZezWKTx+wVt0/OWLRDU4gImDC1lO57H
vbB+qiLyozhALQHh1fp6azNNWJXSc2Ddm5RdP8uqoEBVoeLIc9AaFzjrVK22f5pt
u0qSp6aYFvshjdKZ0R0Mw0iktexkLsXC4tyfc33qV/iAYZ9UmxXNdcTo7mKyC85G
I2diABMOkldG1Rou6MoimVxbwfRRgQZwAHUlvlLCOfVwtkXy9joCsatDORmfpkYw
t+HaudK28WZ0OZxvXyjJ8vqz5v1/0nU1N/YOm20F8hVVCzgQ1gWxIMfdDZtAC+sU
iXbawWkusCFAOL9Tc1AQqHQaa4S5h9Yo6eflEkQzoixnDlk5iszS36Ks7b394vsy
54wtdEaPb737LK2Y/wTAhVmaUuKY4JrMLCBlx1Fu8FRMduknAeT7Qf6Z/17gQs5X
csP2nJZWGEiwTpd5WaaJhKvVUOc/rVKdMVQ9Ouf+C+XiG2/dJIuu73yej0FkypGP
85FAUb1O6FqSO8Pi0DNXvEb7O8dBA9efJzRkfMRf9DZVMtIFYnYVAVE7LTrhP+OC
+EB2zGadQhOb4Udt2NkgdnbbLMRDozUtOZddxTQrihmcUqs5QanD6zn1nRxU4Oez
6b5BOWSv1QaZ+06NTvI6AVyq90GrvsPLpAyPqg1nAs6V6Q0uPxqXCIxq6jsBW/t3
SXpzHN0N91qaFpj70j1/Z+TmEUmIywh/ZK2y23oEJvDxC8PKjr2eUGB4jgJFtQEI
k7QywuJ4x5dGORfapiRj0ZCWW27760IARN6BZ7r4wVvWqrONwH3Ocn1LBw5TGa2H
RmwTSwlR1/5JMqZmcVUFelaO1leLmHg4lPkbbviqaHTTZnVz4v5sYwkb99zlPTT3
Pv7F+sWLjkePWZ0sVlOUCQ2gsS+pA2aGdi82UV/mbi8A30qgQJtUWH8r2IG8+8De
7Mfg/FhPj+6dSKYJjBZhZ15O4hwpZz1QJkwQT9g/43fus2HYcNMK/ZbcwXL5+bVt
dvnhemZcovwL2PErmeXNK2IDjpnPRgPKJp8DaxLtjk00iued07DS9bY96nECiB7X
+0Kxbj9ezfW3g+pLfxBu0n8uQ+C8eXU5MtD91IUUiyRggB//UzdJDEkPvMSJPPwW
SoUOIgJpbOWKug5H+3w6XqVf9+FTX08Y30QEg+aKAv4jX/najVhCbjSnol6ftGot
k2NxMOlOxIrCRiHzZyIJ0RXJg6W08dmf27kqGNefS6462ysVpU2xS6JvcOisvNHD
Ae0owlYHR9bmsyzAEHObbFb6AtqCgeg459x+wnOqRRKUMKcOthUVdL6rxmfQDb8W
Hap/b3AJnw9f+waDfBDxoTslUAwYhClBe97encBjALDvYJJmDk7iQ9CqrX33613R
LRBvdnc3bTq+vjbVacz/9BUI4XdMlGCAGfvwBfhJ8YUo63SuXtESqjJdNeLRIEyF
YFOHQd9mS3KEfUQD/zxFR9yJ4Gj7C6pCYFG23XPfXqh4jlgFDi/QxGb/s0u5Ycpf
lBXKzSkdiTSNacJfCNGs+/4QVYp5ZZpY5e2Fe8s9vOV/46Sq7E70jLmzNdlVygI/
fEovxp/3bPWWZ6KkSzJoUY8HDk5U0d0Zu+4nYTFKCLPY00OJagq3LOCVxHUS7N4h
Sg8z6uMsl3lgu15c5AvDX48m31hm6Mj/Ro0oXVt3aBPpY5vaQtEwPEMW03bWj7T3
wE8GWKnTnOGzddx4Pzu4fZUSGkCLisucBSOKpN0UnpTQ8CjM+coDiWVoWp0HIDwB
vcPRgaHCdeGHay2iqDFFxQYrqHy3XuweLw3xsuYIFMFiKPjB3VOEKlRRx7pB0nnG
Nb3Ry5g/RFyeBFuYC5Hy8SOKfBDF+W7S5JRCoyUsBzs5mQuYVNYeBNYleKCHkMrP
IC72FFG5OQuvHPPXWw0fxT9TwtAhaw9EVg7/ufSW8Ooc469S3PwY5g2eB4dC0vxc
ac4o1+r7wKvMsFhGYKJIe4/2WIgpIUvSL8GOOvsrrD3cYURfFSGMLr/0UKT/IAUX
F5cIw4XPRpWNj2KF9lcHeA4+B+dKMSYIjm9ovtd5CmeBiI54Ag/UaKHEiihonsjO
bEmtq26IpSj3lny0dzcuwgSK8XAHtujfVydwa67b8CoevEUPOCTJidJpfVl7drVD
0/W62haN0Gft+M+A1KL6d0QSJBd8DVWQ+WQhgocmj+RHTL0upu7yH3IovpGJluKT
OaENe3FO0SKle8pQ6H8DOaxQaMX5zUinmHVzSUzgFtSAp2ccBc5I4DeV/qL40rJA
ijobcIKzjPR+ChY8aIL3B+9s/B8ZVtL+Gv+MSy6l6oRGF/wMEzKs+d827Gj/khxi
6Ak1RqxKYFbXSBanf4mF6GW5D7azeuJoViVE0a+UzP5p4++AI/XxOWHBILNYbO3L
p4TqnrOBSebvN7E5Jjq5CLFedXkTcRfjUZGAJWf2ffyT3xdNkkog3GrsbEw88Hcp
/YJACNPTvKwRXI4ccb0FEZ3EveAC6FoDQWZdNG71UPbQDVYvyrQ2LQKjUzc7mCKN
SRJnFN5Vwx1z5EWVjt8KNvFerZkzM7CuKokECZ5tUvzYzohGjX0vj+/2Gebm5H65
qMijK6XmOf/rxV3w+4Jobrr+YcXv9BiqcgJmKLjdfFMvgxP86KR3RR46Yi6INgO3
voKLHBxBNZuci+Lx0u9UOgjziAdfwKcbsdk3pRohe9XJFXaTOvBdK5+8xh6t1JYn
Ih8JIC7NdUt2+bPhRDugAWtX7Lfj5moc6vvqFqXvSFNsCpBjYnypacmQ+Wrmx2dZ
g0ir5SA+slRQ/5sI8sVLmhjqP0L9ojhdxSjQ4susTExg1R0gp5NQ3i05b8kqGhZ4
2RY1U4dwMZghWpf3zDQtNBB2wN/9nL/W2Ke5EMAJnZ6q2bF67CmK4wV5g4dYYRbX
Gpw48Wk9miFdIl4oCr2J6P4BDiLH5hRpeAm2GlS8huDju/TlcPfRBV3xoIn837kb
P0ZZYOqwxBPJUyARxjzB8NwGMNCXJcW7dWunIO+TXfw2+K9O41dNosTMjWwq88en
sQ70zSFkto1vTRF9Y66dqKN0Wz02fMnzj+JPpgkKfvfED1gRyV+zch6mnPVKx3Mu
6cHN3Dy0L9urC1cI7q7A/XMTLvigxQ6c/TbT7BZF8NIdwmMwRXdH/xnqvN3mEStx
CkKsGCF0CSQAQST4qhmU9m4HqY6iy3N61MtcQF9ERMtECWbGshjaf2a1B0a3Yegb
zhhDTj0TBvWLDF0vqyqpGKDC22FlbEnPxZl7xpjX0cNmsjNtnQGG6i/UET+BOJ1b
XQSMGS4JkEj4BeLKnpEmbLsRWjsEXtMUsCPfV9qaIKWgmQdr9I/np7cryDF5XAHm
2K4v9jspkMwqy7PamXezWvlfCVn7HkjHvFGNGXrvfuGOadiomS+nZ+lKkl6MDBcb
6M7sLhSO6kb5A4ZUs61kYindnr7llhbWGufnxfz1+Tc5bbc551AG7MOLwm3c+2XE
UzQ1kvMsRrNtUB8x89u/T3DeJcVw0zfluXNcFWrmcsw+45J/nPE8sq+UAt40YeIA
cyZBDtyt75o2lHQS1whNlQ8yWF/n1Jd+K9suFbrMvF3TcrBygAoIELP5JuAtmg/t
FM72GV9IO5CHbC1BU/wTK6iNplJm/lyRaoebSpSCzLh/eRMYIxODYsFTNEJBPP+O
YNWQVcOb8dCvq33ffWEJgZ5TUZ7e35wv2j1gi/DxrH7cDC5f3y86JahZKSud7LPa
oSxkoTZAScK+NZ0jW1a0scJqsTAqWhFgntlZAyy/A5FUbVZsyvUAbUlNam5iX/II
rdLletfA/3W03dDeG+VUD7gG+O1bI4+OhzidGRo+6lwT72MFJo1ST5PzZ/qAJ54n
m6TU7YF5uQsi/nFwGJ8n8LbiH4Y9VeTQjTzZnn5556WhU2nHlWpZPj1fIWwPsbBD
jimg0baPNWLwT5/LVQzlI1sJUeBEbW09mAMfPYc84h++/5th4EYYkDUMFagGZnzD
8mNmMS632JoC1edSx/WJC5NLYF2puzwo/K1IGJWBEu1CGB76BOgOZKBcX3huOP7U
/z7h9l3O6U6FFzDThPt7tqnDYFqRQ+2F9bgA9jluBdpOYGWxtSPdjSbjJr3t/1Fu
wHZkjQgHcfOqf5QlKtE7m3WGt9wFBlVYkE2UpfHDpjDwDP86emwm96U3GcxK+izM
Fp/9ab3oSEhTO5RQDxOqcxGvFomA0IpsH2nE4kIAYUzMLsbGYXW2neHW9zy817RL
OupTIYyYR/AdfbESXHvDpgF2rNm3ZqTeF6mob8aRXwCEIS8/+b+8roJKgwSYljqr
JKSAn0hkWDVRJOB1ZTxRilMNU9uVYaSJ3awOQy+2QCG3DyKIn4IyWN6MNl+zBK4C
3ghyfWPBfkqJbip4pI2trUIs7xTV2jDZ0FyMmXp3LzaFxWK471B93kJYwt7nAfl2
FQbywhnVB0w5NLVD8Mc0aa/eK9DWdcQw+5Um6xcbPCsRe2nsWxuIXtSo01nbOnkp
mlYQRbuzo5waiALg5XeMf8RUNsluoKepYxZcTCv+6Mbip9MimTpfenJESIQVKAiP
9DHnzazjf5T3fA4eYVONCYQwTsj2uL0KWIMjmcR/yHXyAEyWDVpAECn8J/f70hvc
AuBT/4dWr08IEydimOItXwROYaTlLIOb6ZwuWsNtGfenyhlZTVz9iE5fdW1UzhUp
XMUJEaf2cm54Xw09RmgOVJ0G0rHO9CWqfsNYC+zFrIPegwfry8AgbR/OR3PJCCMZ
uxnz3v372SgPUkeXTGfGC42JmMjuN7+lNX08WdiI7D63hRo4th+NMLwWdipNS8CH
d/IcD4bDwTRiJ9IQGZF47Aa0E+IaW6cJ93ghtMCbniSlGkzGoweVHKtffc5ahGK4
PkxwM35aTrfODiacW4m4TlMFU9hKzBdQefoIql4txhLqIhYT/FaxlUdjILq/jprb
vGlozP1DwqMvjFijCSJkoGVB8SL+5i7/5G6uZglesLshYKnQR5+W6M+P9LGaJcX6
usVNoTsbVYJUeaH4apw5RrFX+CdLhKpE69J49UKR5TCTf04kh+ULxeR5OztwIfwh
oJFH1VHZ3Za3lhAmhRiht4Lwqtu2pWnE5BFbWYLZPQFRYQaXk3THzDVOrJ8FhvgC
gDp4mewYKZxScyOyqA6/TMwJ5egihSNYH8AeK4zhUZWNE51DRV7G26fadYedZdWa
9lAbHzkf2BSFiAmYtAsZyU4iuCUaKaIkvOFbZBQASArk2Rl3wwmHzRN5cMtC4LuK
iEMK4D2v9JsKm660mdrn37o0X3laJzjFfiXLn9a8pOUUXVf6hY993e/pHinuooDs
3TjD/HVavlxrh+vqYu/W4FAkhjOAubR6L4icyAVOE2goyH+fRIa4RZ104GUTUb0q
mRDC5gsGX1V8l9WLCgrEYOhGO5VQcByMPSsPylBlvE1yovdXM8blSC/EiznxyJgC
A5tuyRsrffy7POPa9ZP15Vu0NbeDjWIbLL4I55jSQG4geGrLqPs9PNgKMnIz1uBa
JxPF1ELNEUrTBkagqWhhy7CrVpbeymbRrLlIuZS3jTJkBUU7Qh3HCg7cRSpBsmkS
Tp8FqnJTpZmEXk6dpwHaY6TcVQM/HegydjIHa+O4I1TlTStCMpY0cl5gQKgJBgcN
U01CFwShr5d2ue3/Ct5TKj/pdqR8zsA4PpRlWmQ645Bez5WoR/561tRc+/VUP+y8
9TAjxjsDrCyMvrTqRyVER56CkVX8+Bzf16xa1YL6r177ciSjRvNrKM8OXvFHpwJK
LtTvs1B3H6zWr7g8lMy20EULK2jjm3PMaouUjUvhaSzpCduq3lHAhOCfRrqJoint
+U0VERVO8kg4OPeKl++1m6DLcjbo4RigpVlKuYGf0wVLtyicj10e1efo6IReqwd0
ssDiH9pcNnHCPFQWwzeFy5ocuXDAE6olFoE40Tg550jYITtejeRsTGUqcLH8N/iq
F1E/FO1GUaIpeDpRWtMpaGdwS3gSbpCxzRUx8LcNP4uMlJMcG8I0PjHyD79SQiUQ
yrhy9ymZsarkJgMpo0bGdeig0WaJoINpWd+ePSzO3l7tJNpwoOvmj/ON8XFqWuPH
O4Ygs4k8QtTy3mckz+5ZMwjF/T8qJYwX1dkoc48gn8WlaNoS1tnIfNv7o5sgBixN
7wGLEy6bfwqkwAa427w9YpnRcJSkuE9N4tVnN78sO42jXmSeECztQ5JB1sRFdEot
BxrEnOLG0Hh2AXp+E1wnwUQ9Wsvc9XStP4B2ArCT4F/5IfDb0sTDob7NJGKmbt6z
XNXHhVBr3pzlRGkX2TFso+HNym1MI62JUCfqIP9wbJMEnTrNv7imYvFqHFafznpN
0/2h9L/EE0dizMbgq6b7M0wVeGyAoNshIbchDEeKGxrT2VuZTzHs9IgHSSL78O6T
6ofaY2v+gNrj9Tx1m9nkn89DabTonXOkZYvFNnTceJtX+wU+tfQjCg6JfMMRWbRk
b7B5RJ0w6lQ+XObfRb8U/NjqouhS3MsYarAfBFZm95M8dU2h0PhChjy/V5Ta7FR/
wDLswGs1SMoUg/8AYd580bPB4NpyqJ9TtBARb9FOXq6BbgDhSfMjkCFeSppffjCw
hglN/vfqfQpUMsKc9bBhVtW0xVUV28HyeD5vWxbz/TXwLJjdgLWjbp8uAIfWWQWe
ltxSzgDYv2rUHGiG7ENyiqC/pgwL0mBDnF370YkSlt7h+q0AKJf7iNz71Wm04+6h
ZO+ZxYX5YXBYWlVutbFo1oIHSjPlkN764Z49eiksnuO5ZXkh46IGDqG1dVzmU9L8
78SNSwfagWnhhL2ccju7rEPjwmn0VAelgW5/twmXd3fo+dSVPe+INpdy8MYrxgz8
gyx1+U1wV5Y2LQxUqXOobKzjky9EYh6uXjJcED2tHIBwrXwBsYgd+UqmfRuf8US0
sgDv9VlD89VkH/c0aX8lqt+cHFjgJmy6I/xuBFo0sRwOqtmwsiFe2kuFh4ioz9XU
SuBGhkjmdhFLVKPwh6lgb4Iu4XkuK2lyj7/TA910XFaEtzMychAOS2RB1n9rXncD
ZdzbogQBazO4+LrVG7PvYz7KYo63TtL8pQpc/uGwLO5eijcfDv7LpxIbbEfHtQ2p
+zVP+arl4Z2QS5xTA3ZHvZ5dIQAxjTJpv4FRHIkRAffE8YjpRPU16T8mQD2CQAxG
qqPcmALA6tUJe0JG2G1L5gLO5j9ncpDuLuCTO4dvhgchuue+ArQv1tFbjF0nSWAC
kOFRWg9tW2r4zaNWYtOS4rtudf83656VoIp41bwFHPcHoshHFwwhA4OMPJ3iRmCM
DunDbEnZzFtfrs9xJddLxTwazqFtLHyNXLZ3/4JSrs/NiCvJa6x3jZn1E9fNi5dJ
chjHNlnuynXUZu1MNP95rWrP1jmmIxKH4s6PlzBpQohEsEtCeKr0xnFi0juEKkwM
zR7+klyzof4nl/jhFDpjGCEA3owSgoXCJbJk3x/qCk3cRblaTQL71k3Py77rFy6/
ATD2CSUACQlhiK7wExBpj5oeXGyssIb0d9nxJwHiCKxVTLO0RZfUYiJbwdIZ6Boe
9hdJ+Ba0fN+6rS4LfwOyUH5Lc99+HsrP9o0aan2LR1m0zUy1w5aJSrVmTslo048C
4Xq2J5q6O4gO9RGrN7YiqacO9Ho0i2WeBT2wME7sbzW5e98qJ3Hl7PWrJFNWMcW7
W/gZUHjSeairM5hBfKgotRC44kEe4MifoZcpGBNBSUW4NPlIVltt3qbHT2aIbGQp
+EXN6e9AeHS4c2EjY5ZPRQm51TgtCZip2Qt2q4aSThGiHcg8lJAXUUYhD6O9CE2W
JF4OwDUvZOoIResZUR1dLc13dk/0He0k81lapHSb1fh7S6TUlncMXK4zXuk+VKVs
VeonjoIM6jFw9GK2ncc9rv5U7EgoO5sM9tTTT6eyVDH04U503PtScezdBoDy8WuA
kJgVWQ+YOtCiqToV+Ukj42bS+vDHaR7CWHP5DGNCpqlw9ynXB39/YZVpHXioAtnn
lD37J2KjrlUaPj4XM2pOx4wXYHZwqfAjfEPdu/rDj4Y7LxzVofCp/rgxLmNDacBF
LQgjsz1D2C9yGtfLdL/k3wQXCSs4Nreq666dv5W2Fo/bEWFXMhEojoF8uqV9MNCV
Doom9+C0kUqMfsElclPqzHYyRdzXDm3nOZZM5aiSjnzgmXYBuZz9XR1zkeetUDuA
xuIDAX27RYG0+vmo0/aJ+V0PNCwq3g5aJRPyaBl6DoW7Aw2WJ9QtjCuOFcO+cSCe
iXbdIzOr3VTDwIfHdFFD2U/DS++bWjLFS5SyBCvF/qbE89O4ISByfDsfU6n23w9A
5EyLKYyAksDqwzXgNQ9zDM4mExr7zsOxjUNt9ukP9fVvulDz0UnwgVTqb4o1yR59
tiplGjnixRFFGXVhFINwiDW46iv2YgbLKSx34lUf5/LI+oSqU7kN+R2MOV9b/YNr
8zpWIydlVh/+VmR5Uqb7du2gNYQj/IAl0Pmq6RxAsDz0iqoCh91AxR8LkIKRiQZ5
ejRlTKKzXRMhJELUXhEmcgOk8ncciq6dm3Z11xPD4K6BqLue1DNEjHaRLlKyQ+JS
AyDCowG3p8ayn6opL+0eJZoHBUUYw0FAEsRKzlruhRFt+J3KheOMXYe3WUPSzPI+
rBeYeiG+SoaVGY6b5izEpcfCZJCNbxoNRwyttYagH9WiG+2WUpyaTXNgnFmN0Yy2
8ThBubPH5+/JFF7CRD3aTl78+VMrZgMd8XnSJ39wS6B4XwOBhKRDpR59dpG6LrXD
wFNteaaF74mlIii6gIaxaODVG0Uqs8eXqbpRAsIbNgQc+Rq468cXaHUv/CI6pbpo
CjvicSDOC3pnZiWL4ZELpmCJjBu+qUra2WgIoNIrllUpkHZFgQ22PAPA304A6Ikk
/hGkV+ALSObtlzab4F1eO1fHQq0NTtcCxFk6YhqcT5+/X8VCFPhVxKBNzaaEEWir
zCbPO++jhoG++9bdh7by45J1GJe1E0LFZ0xK+fKCJXU87/TWQohGV7fcjcew9pen
Hh5CZ+L3vNtYTz8aW52h1PFJcatwWsQzOnBsKNDBW+m2dhojrUhCk6DLDMwfh2Xj
v2yU81Pc8nlNcm+cTwOWuEf2Nyopm8jP9ce1vjCUJuqU04a9uFpqgMW64kq12VKL
5jX2XjTCcuTU/HBxSFYFRNTHWoKbymCYNUaAA12YQWnc+FsurlIyVfL3L10RKpwY
DmfbUm5KBTMTGTvYzcXlVVzyIWHP/+NS5kYcZX5mUYwrSL4FqGH/l2ZkTsIuCYLV
tEjGkiwTsH1Eai9xhndUctvf+lVVfnqyEXh9jvii+LfLtalma+mOdKpmYbervI4/
gs95f2kg6qCHViERico7Rmj6kjAePMdU9cmsHYG+fupzhBUd8x6n4D7ONr9dF/Fd
ej11B2KXegRBY5zvHyzbhR0jaVlbu8tokyhthnA9vGQ/i+RG5ddyONGpAiW3PTVY
gG7tOx5DiTiNfg2gGY+FDYIQZYE9Zavzr8cqmOOKmyoLhgiR7X2QHkYc6NQiSnSH
K3ARemUZfrP+F/doikkTknFBogHtSnKNOnfDWJlpEL+uP+jaQHTay7mZ/pKsauq4
wsQSCzIdIJeqEHAfVXp/79KKHuko4jkXh4VCdQD9LBaMTL5kNpCDI7dVNbAHXvmT
36JAdnxn+jgYVVdl7SGwkymTgw3BO+r4mIYDplFDPZgexKvCqLuf0/cePuf9W2PC
8sP3TScqgJEnjkQwzcb32PHD2KWU62Ahu1Odjy87qbp6+Gl6pMPgK6GOdGkbwKA7
zrU5PUWkYreNYWbT4YccFsN9v5ALYj5sHOETWuXh8zlZeHM9Ak0CV7LJFgpb8hKd
6IcXt9mUOX3xOvrXQJAtO7pWXhsYvJzcZoMaSe6dCivL7QwupId9VMcBl+h9Qiu6
DuBQuvKDXXkeo//qrCHmsniQq976stEYkMehfw/UaudCKPE8MuYeTFIaTZPl208L
2wCfDvD0aZkP3gU5Q0+nWL7yEU1caUhNL6c8ofFCAudfGJa1X+qw6zv5DdzFfGjM
M4MvHkCGkkVacR5ZmWNMdzLdD5BOdLJvsIJ5pCdjuGJo81FgxMTNnQJzIqFkJl2O
Cy400l4IAMJr6zeQcJNZGg2bV6nBqTPqLqg/iOAMtbR6WBrgWg4c3L+FdCDZDREY
4SKiSMn5J0COUJG+kgPZbxHHVShNBcgz8hUbE3k3qbFMjvou8KvtHiyGsQgxWtFO
ZeA1+EtE4kc7+bxKeWJzy3kRPNfDVYVaHmpN8gG+6arwehZHUda3bRDF2uHjfoyv
k7Hzp1j0HaG4ftcGwLUP3IfqvXCgjDmSbHFB4sRiXMNe1G0cu6LNRqchqnWc8P15
5Flkc5w+LMDyvVuJ8imEghSvFIPVTq5OVM8GL73VCEaI59yzH9rNq4sJKJpdHwO2
aR5kuIDS10wCKFkFenqr3Sa5MT0oRlAQxruw+DHEEiooCVhu//MYlBAA/hH1244P
8lYmTCcihc2s/gR3jQXzNuFFj9on0cNbRoxbqTmxyqQFcDblZxgox4Lz68fWh8N/
DzHWHg5v3cjpsLHbIif08sBCbF+e1RdrcrkVifz/q7kY6NwR/zzjA0zKvlh6eEVg
HX/5UIGEBU6qY6Gg+gkCLDaeQchFkbkJe1biXa+23fzoLdu9Em+NUNUVfja6QkDf
ulLoYnShX+4+jLJy9FJ8t8/APfY1C3IpThKf4lU/yAYVZhD+u+cdoJLbuWHOc8r4
8+oVKyzNf/Df3uUkRjCcvCPk1p/oBqaxlUBJqAztoeeQpuZPyJO71afgMy6uRELf
ov27IdPgWtTg1g89DJfKLyZrItHhiHDO7+g5HQrmM5BgiligDf1+0AIxhF1IZYPV
RqgbCWqhGcVV0Q3FLwQyyYvZeIb9RXuV9CU4s0EZLC531CQThiw6+3WRXdk1flJC
Q9GRUvl+hGx2bcjz43aZmuozlWxqdRqRzltWQi9uQldgOnI5kJy4BWENXlTkE8XH
iR5b1cqNA/uMi8C4bqtxI8ftarSGXrw1Evnkvrxjrs5FKB18N6rtPAU1f9GaySRT
rpRmjiTe+NrULf4BCIrs8GLttgZhyhkp3iiRlb9uOKowN9ca57BcvWq3nhYaGNoJ
uXNHpkTuL1bWESdOVuipg7StfiZ0jWD2NwsfshJhxbMFsfGyTiAyDM/LyahoKcOk
K1+UvoSDUxMPZb5rN+hNdRqXov8w/jrX4bbfjKcHBjTZ8+PzGvjIYWNkrTwkqhuS
6czLUaQjJwccdNyTI3MB7KRlAFh5BzcIKdw8H7wk3O9IKM6qxShupbtKKmV7rEO1
bhKcGHcdBXgkxgxUtSg4FpyDFZAiRyza77QQ8CM7R+zuN+7KfUqQ4ST4pDjs9zwK
ehkCMMbYZCHG3AnhcgOeHpGu20X02LqCfjncYcXCqIKTJGnpIGKFBOwghGkCRpnt
BlJ2cl+9trVH8wnENz6ag6tsytWz9/wWLqQoX2g5ebPm3dHin5BKy8kWPFVB/8Cc
QJuRRH9k9qCtjsQRW43nOwkRe1nF+iB601Z4891xJbhPLZUVKKwPbg4NrNLy6L9O
dycUntBRA1k86McJTAOOcMY6Rg5AMzf+4BZSFOuY2WPYwXN/qBiQCAiyz5GWMGAf
KDT59GBZybRmaOEFG7OXNUju0goFFGazmiODd7jiDxYfz5M+PCnqe+j0T8OaD/lE
wJ0YyChhjdbevXOAitFN4Dfiij3f3dxf+9Sn762tLQIB85jHZZk0VYyUU5jW5mNv
K7GMjV7ZmndDkmuQCIu8ES1kl9rWFJWb142nnRhANGf+0IVNW1vvjFy30uhpTQzF
OKEknmbR+zaAmM6LgnJi0OJt9dvCzWSA56sZhQFc2Kki3jkn6s8cXvZb4BUNpkC3
ypSQVSMmgvNjWZijLY3LCc+IOqYb6yEtV2zLxds4B6dp3es5znqQ/DXUlhfKRcS3
Rk9tYvqOc6bgjXxMcrrb/sO/Ygi0fp7ynmaaoJxeoFnQHrbNeyg8WHB91pGsbDxs
VpSbnO4kRF0sfsj69ZV4UEqNggPWQqBo3KT88iXgY4TO/V6H37fHYp34ltNfckxE
ppmGlFtz1swyxttfFOgNhztwbmWH9tRn6S7puMehJsCz3QIKK/riCpervAu4FtA5
xKMSNWuARllI4tJrLe5jgOl9+C73yzBJ4lszhuXAm7C0f9h/uHjzzIAwdgir+GM7
8kIsfwvHSRxg9GoyAAcat+qpdU6auuiqhoGvldLja2Rwilm8xSBgce6qgkY7ShS/
7m/ISISQklfI/km0pcszZ8fxzVoZzJqWNMEHIqCSQoO103tYXjsAeK1zADv6z0fj
APWFLmDxDphsOeSoLfKciHErdC98THXDqcaVl05wDrO7gZzjt7hOToI98nl1xMgu
aNLwnAb+m8qBz1HESuKyB3mW++9Mjwj5/0M02lhOwoP/h/E3udNhmgmUfEenuf+Z
wft2rhLjAqP7rjCHhD+Iv14PiJd/eAx81w+zMfQGsr0CCj75HtWfHPZidbp0SwkN
M3yzMe/AtB0wU3xoSq8cth5VkXMSWP9RhX+d8zjEUjvTLWzYjXY/LeJ6ZrxKpZtX
IcKpgmDolBEIQMo8iw6NQlEgZkkSwuu8pgYaW/WDyapiQ5PNMvVdQVHwyrulOiX/
VhJE/y7rJZd+MI6gmmJv0EqgbHpRX48juIQDX3MtJg/XfvK/Z+HuSjeUEb6JCy7Z
ePYQ84bEU19bVZo6esCNz8Aezxwk2rzanC8Xz0lAJrUPcJZReUiRZEZB9AjIJAzF
VEpQrXe7DivskVOtmalEHV1I8cmMRy96WLywZDeRZRsNava6N1LqH81ATk4R+C/X
o0HNrVbwCALjgTANQoCicQuxCibuUBokVCh94dGD0t7Fj80SOgO5CPaGv8Km8zOU
0uCBvOyvpwBHMpLIFXAX3w==
`protect end_protected
