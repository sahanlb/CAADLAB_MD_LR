-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Yo3HU1OOgehfjGR9RjbHLk9vjD9VcmeAq3uIaBjTgtxVectkjU4NDTqtHO+R9u6x
60TJBLKsBkntJ/MTCyiGaRiY7lHIs4jgdWl0D2qI9SC5iDJnoIDdhiDXTAcvz4Sj
ZplTXnWaZ+4VHZrbyWfOIoIniO2YDouMEtHh7do42S4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5980)

`protect DATA_BLOCK
fr6yuGiGaySO6OHGJxEUP55f0Un9KP5kppdJGCAUeDMb01N/RPuKkYhrXkYccBpT
uuKhrY7z+/XYTCNYTm5FtyaAWWnwXzrWtG6qdoEMynL8DH8jiapQd05TiT8g/Ayt
PPQDE5Dp4jIbJDwSKQrAnKLt4RuBjQ+H4k4hfNAVJHEq8jR86dkv81k2+YQrtlGZ
2xQHRpoi3RiUhA6XfwrqPa3PJBYfkqrGVZt1vTT8ZXaIwAd86ciM9eJFwcY/pmP6
B5ia9KQmMAx5ih7qGxUP5CJ/47dc736uD5qf09Qxs/dONT3GLS3gIdrTh96J6Cy3
HXOMElwu0Y1cJQzGjks6X2pU+sbHUOw3fye7XrWLV5umIyhRM9tsdjwYOPZwW4NO
0PqJI9DK6vZ7Ok+vF57E36YoY26Yn16bME5rh3kq3uIfrGZv6W71wBk0bzgk+J++
9hC2aNq/ibuaCIaemhLUPo0ZGs7Sa03D8IpJqLjJMCfEx2f4NDexcPvf/MjKPh2W
uVBAzcudHs750Bch8F23O7LylCdputCBDkkT4SSYLyDSrB2n6W/zZQ74Q1gQPcBx
bbw4OCdSAxat+WxlvUOfC7uKWRJUn1Vw7CGMo2SVmz5IWk2Tay1dVb/cSUBRcpfu
qcFL9o01Hek5LVoa1SmlhQRIMEahYNN4JKnD90IY4SQS2xBHFdfalU1ahz9nkUKo
aHs4/dtw0SdVk5pG9Nw0UUZmuQ09l9joHYOQREmh8iwtz51BPh6dwnqUIx35NrTF
0G1WyA6mmDUswOaY4AbaT+/w+2+WdBCVhFqw0OBT/i5LnLZNW9rpm1bBfJ3Bs/on
O4Gm1k/bBv1sxhdoNtqL1xHymSVzOtA9IrLmmava6FZbjklqc671DHjPNJ7kAv6o
19arJi9cPaJT/UP/XI3515nEExcY3+SP77qtSYXC9UohvZUPWUJVSu2l4XOneDxh
YjORCij6VioK0W8CA1tABWNv5LWiQam01GIS7/I4QPRsmAoh3e5pc9/kWJhA8XBJ
1MjJWfzBPv9B/zm90+vvY6DwMaLTSioLC38EB3G2/Q0fbTak+HSlSULQbkWcD4FO
PL/Gi4eAxY+qGCuf/BJCtpkeVZ7xQhZbCYF6wO5O8ZiEl4BqXp6q6fNRSDod1nnE
zrqagI/HJnU5M+lhnGDDfRrhojQk4LdQwuIdgZHSRRJGlREyOHLDRets496TyIf2
iT378b1HDU4ZWzXZA5oDsK44P+EoGN2BiJ2PJ7dTdMTorrDnDAfHw99+RGCLb1uk
c66cKUcgr3ZFdtJWCsPHTW1m0Cc2+UPoRVmL68RlvVQiS4DKJHNR1GE99hkdnBcr
DTev38ZH7rX1RQ5wqy8/rwbslr1TrjYLYTxcaOEtcBDdlLSm5b4UP4JFct+XKTcT
oFT/cQ+cZGOsLEfHtNpn10I+eQrGTE8lKJd+ZWEhbIbsblFeM+gO04rj2nUcSQ6u
+VYl7go5OB1e/YK51YzAaU9D19Gz0MYZe9uDLuoJ7jiyPcVKqzol5B1Qo1jNrZEy
w6Tyr3+r1wumqS02XzO30UOePCCbigWirXMmkRDK2VpatMSSMEQm9pNxx45Ng6i5
vqH91AWpJbMWGJRUAVpiVWTKOXaCp3npxa8R9wrhYN4tZnuz7gbUoV7RMXPK59MX
JaT6MGAVxYDkqhJYceg+luP7YCJMrWQA2bLcORcLeWuR7I416nSxUESPFXKfL/r7
THvshAMEwqRXMgzrAoAk7TDztAKqvkpbyWLKLjIjD5ksyj6C4k+zy45I5JUZudZt
VFpQGhKA9nAoJJVPO7TWF5WDkDu86Z5zaOfisSGxdg4G/gFjWlkgWqZRVJJtSaNi
4PGMjTkmKEdIUmAwJe6rva3ZvlIgvCop9GWgXCkHA+K5ICd5kfIVX/f+IbcPS95M
wrcx4BBRn3pc1sdwcxMLsiJ5dpJZojhtL7eLbEqJMxRGq8uiDS4FA+MEfyqmEjNM
s6lH/Zg0S3ZSkV0SrZOkniaL5nyrSf5Qvcb9W3VGUpN4+OUuVJhNjUwBvDowd0H4
e/ZGB2K1huwAilVX/ntGn91l67VjIVVcq7BQlc6RqRy+HYzPO8W1MESzEE090jOz
y4dVBGrmZSSmxYuOsg/0RTK598dAmwkPVUf6MvaG2JNKPK2hyuIW1i4EFZzNfOJQ
+sKk/6MNRWM4j0kcvOPUtlfaUvBniFxRB9mXY0pX3KSvxy/1Ci5ahev0lK96Dfit
5QSPh67KG0HCkgUx+tmYGiKvnEUazVFaVsv5OlQrtR45otcXSI/IHSvoALCobvKi
6R5U6eA1LGB/+8EXTut6Pl4ceE5+5wa8hrXCOkCalpTlWB9YnEbdeGZSTydO5xTP
5glTazsrevPId9Klv8vuGOmdhBGpVpg7Y1cLcm/LhfeK5IhNMDT2+bseB2znQsBG
lCTWO59yOEX7N382CX7ktS/BwbR6A6+Pgzz8gvnZELWwcv59LzYMSeZ5LxHxbfWY
XevpGeroCpFWOidjEV2kXq0fyU9td37NNHR9mkguT6/bPIRT82pUqO/wvDhOjk+I
4ZYeCW/PZ8fcXXN2AvVopxhvXFqTX5nDeSKEcB2HSMrYi3hJEX+CdHKy+NH6aIqr
HGDRTUmrJDxnk2F6w7mY/KAbg+EiTHPP11JiT7ZxRhFyOXO2ZjUe4cvaYDcKKBFG
ockp2lc/VXVsyC1PQvL069puvKktK4j41iGpF3FOZo8Yz3OXdtZxCBP0DA5IltPd
LvYcxBCIXhvou+7P4V6hCYz6CEgWiJTaqqgqxF1N38F6fdr/oAqTTort5s00LGeI
PXbmcdMPazV071wJS7Zaxdtf02nL2SZSzrUVXp0sE9SbXXaDW0QFm37Ut40T3TcN
ddIxAV4gleDxw6q+wnojzAnxyhANbB8hNFgksEc0qQkUcfJkRKuoGuK6mUrDL4je
2AWbcii3NxMx22/1FiMxJvXqPVBAkrCFhJfoQv5lJM4ffCcMSK/nKZExJF8km+8o
+U8mq1wRAHqeDvGiUkLNqnUsSIBprJnS2Z1E9ydDQuCgT3fH7pDTNxu1vfmhuouH
MbQyA10AkJWIyey/DfDvgEJDX1vLPHDaqoDEADy/1bMlVqyY8P0BnJr1hTpxcCIQ
yuMN6IV/SUzWrC+6FuMAA+okZ2iYxlz5v/hVLshFO+lJowqdLea5hkpDpkrN/N93
39lJH0ocmkTD4XbWMtCQTATZRf2Ih/AeJ0KKFcHa+RHbBUEqZiEweGvarjC8PSg/
WaBo7izPhlhvlJrKHNz/8PoKwQA8m3/O4R903ezbZIMqngo9TCCs2fZaiKVsUgBc
7Ap8v+TXUzdMjbsDLZ1RPEyhn5J5cGH30lgkYee47s33R0RRaA0MawQJJmVKJTtR
4vnBBhdIuf89fVM/lj45YVmbzs0mQK8i69NjDhw1JtRuZ7KDv5Ze17OqVDOd5Dv5
DiYH+Sl6tq6TbO05rrwmOKitL+mXj9PMRKlpXNxxGIvo2rv6R4ZOTZPlKomzFF6B
tfD/500VYO96eXUxzww9SXiMnothy+5IwncZdrt8Yk5fawyLH+9V9J6pFAnwdHr6
xRfkJTRwSPsDiCfHVV380WduJJ25+9vVMEJVgcE6AxBYSbcYzFQxzXE/K5JO0LMf
qqnH3yfnpfr4Lec2toiik2eU/6neFmeE4mG4GlNlI1gbU/OdLBSP4SjxumSACekY
vJtk3EGm/fSBihk16e0oCkFEnoDnN1Ik3TDryIAjM1UeQfrA0ZjrTCANstBpSwe6
mB+U8n7SNFNFXLjHDAxT3H6KDqvzleOJTdkasieAgcmXuvmwOw+mRQosD0XSYapY
qB7tN5/KsQaHIW1tXIWO5JZOwv1dxmfts2EJFXw3OzwHYiQL8SmQx4Y2uWBaihni
1L1biClWD6aTMPoRbR/H6JZW4ARyOUHzA5ti4Wo0KXejTDc7pDs05XiNiH/jSiKD
QXRFJ3/8uQAu6gUWe0n4ia93djotqV/uFGZYZmHIEoAq32/AaBJ7fVmZjKSg+FQ2
FD/BveRN/lZw0jeAfRIq9xOJguMty+rPtvd1tXQCRPt2U1KAClaLLhBofgFbssEK
ULOiXsyslTHQ15tzujcMeV6m2l9zAoIAU6dMqhLb/hXEw6hFu3vIb0v7Qr3wERi1
QausLXBe+zeEdfpBv8+fpr58I/jC/mVhT0rUxB0GftTZ9OY0qZN/071n4xz4nVyh
j2B7f7tsqUeswur/pxGtW1yNOtUdEAl1ihEknlfSf+ERbGcqmH4Hh5hfhfx16UuO
40wmaBVWmJvqo9EtMxraM6NjvH+dFlp1EympbMTgQ0RoFRYnupZwuOdLazAj/zrp
W8PRY1Ivoy28vrfpZ6BaEkfm23CtBvC2krHF+i96PC195ueRZF47QCnz05ooSFYP
GNY0XvNgK9E2OW9826AaRJ4KUg/RTRC5kFbl7hk3KgOKoX8aVFrZNhSSrJdzd3zz
2KV31Dhotrtz5Kuwh1XDynu7ipbysJo2ERA83iVFtgeZTQWtIOyLOQVr5UdkimcO
xBhPGJzuCd5r4xwnPwoJEXcKaGma/B+xTVr4dGSCnkUYcWweoz+dVWpLcNc3BcEL
ks5VUa8WvJiX9+HIvWBVgLwrOnGgA9SffOSyfkow6hnQYlSvEA4IyUUI0n61X++c
BJr1gwATQXc4EsVjZ9oq647cOuSEOW6kxiAJ/UmXe2S/VOgYDdrp07iPrNPPBSS2
YgZLU8OJciFicoiFlL/0dSb3RWbznn7I5xEhChTruQCpfUlUCT040i48Wsiyf209
ielb4NxV3zpSDbZj1WlTQZ2kxmKI+ul794n3qesE8jmpSzXYNghvGc9/ieSgqA29
tfgs1rxwwKaVxcNmUxVfWRB3JMK9/Gk2uq0M/Zuh34eyh2Y41CAI+BJrg9wYj3CD
sNhy2oXu07PtHWVDAnaMpW09jJaKpr5BRSoXLSl1cASUSXZbBTCA8dXTiZwkJrmD
BUOM5UO1SC/7BcvAssquwca2dPaN+ih7voyCGPsuewGaBoUGu1h5KgxeQbCCT+cH
iiCq5DbbOvmUheD+576eLtot5UuHuPBEacko/+3CX868R8b8vFGokx26gsnsx8kg
6FmIy/g1cnFEoV1jS2hRVl21+UjrTOo3Qjt48AWc5ZERG8w5QWQQjTnBBMFyJu58
BEwi1S+QnmdKOYFVvGakg7zAFuc97bvc8P+O8LLmWGOCsHgSkiEOhXFZfnJd27Tx
fN0pYgxU1bsq051aNpmzsu+PHjCkmIrCUoqlPm9oc3V0baVKsNakFDhoYVqOpPFR
S4IIeUisq8jdfk0bo45l+Pxn/jfDIH4QEP9U/tt7IO9XyJeKWdHqtFIf6S2G9qXk
1UD5F6Z648smkMAf3qpdBBwty40qioyvEQ7ukSUQ+Q3gab9RnKpjCCGnO4dql7+T
TxMC6puiK6xSz12eSBI5ZofJUp0Dcubg6MP7rbgWOdN1enf7EQZBYY4/v2LFyc8i
X/WUZhqqHF6t9QBv6BcHQjI8telRFfDkF2JGKYi5vlEGkfRp6vFzmZ51rXWk8UCx
skZwozjQ0qof9tRt4TqD/PrZC7/yDaXOTLndok+reSVF0oE+SzS1ZTnUSmvyIQBO
bpLKE4TqTRDriCOCZZsBAzBob9ryEM+r/rORse4aFqcjUtutECZFrGKgGYjhktTh
T8VAWm1MZeFYFVI/mVVjLb0NKv18TkbJI+4Y5ytm48qCBvvJ+U/cHmWIMXPhihmI
wleAwJqLH2cTkd1Qds3AaNXxRXcHlA43P+yAopvtYd+0njF7XaDY3/MzSGcxzPrS
dopfQwZCN/6yNkIk9wCPHqiUdF88kKI0PmPeIgCSHd8HVLPqW1+x285YZthTNnvn
1YfY00Ojw7seFIPmcu7DUQWNy0ubPbyBp9f3TxkvGSX7VJ+M7DEYtMkmZHnDFSA0
olHKsDqyE4vAGTaTcpxy/1ZIhhw4/qCqsj/g+Nv2U0fJF5/wfGEwsy2VVZ6anSgG
Xx2n6Mp1N6wB+/z4aiT2mIVhsA8ABW7NVUIXtkuNt8Pu+IxVUhV0HTviLAinkaAn
U/cGwBUhiUuZe3Mw766GJ5glhqu3d5OkrxIlRBkC8VMJ3RdU80eoQGxk974mL+gU
7nnggGZKsnkDC0CEmMWQZO9HZBJiIsR+WavqpkFSNh/0oPy3sT+8CCQkdt6O2ntd
0qekHZDiipn6IxKcBwfdt5xDsSC7b7vuUKmD3LB10uBOL89TSeC3ZqJ6aMjXSnTa
8ThVvG/7BM7SKizuRpKeDvBfbVGuxDkvH2vnygUhaKy1LAZrn99kvikm2G6mtj3w
rOp/7Wp1b9sAGM2CtO4kkTzYJPgNTV8dJ2jHYR/dM6gz1JQ0q7GFbhwuj+E1NmPB
+VXSAjO9JQaTjHj1jEUIjQAByXcPT7xkW1Fets8oa74nxC3IJ/95OFDJ+38Tal+h
NOknyUndyX8dEA6/3vqkaiO9VPrGzDzyhGpuAIXofIXz/ARjVCzX6EHHYmS7z4XP
IGvthtT8eS428mZRweKbHGUKUaJrp3CSYvX7+dp9rOqgeObGhDm4vPZng0+k4ZRD
iySFPs1vnph9B39HKfuFAFmgWIE5+XgMLPNGGc6j/0VwpA9P+2+Z6KuqPPN77zHs
CSd0siryZ1/HIOtxHE2j7tXUxN8xzDNpiVrg4KszHIa5x4RpBL9y9lzWNx3BHKZH
YkpXSc/TNt6GhpFk/um6USMtfo80mU82LrtIJizQgpV0Qr8Xl0J8d1qFIxh738Yu
o72k7rs84g43YbTun7JGL25XLD/eyrKpal2C1gFQT38xMDJ2hUmY2NqlPsW9xdCc
Ba1E0ltJo1G0k47n1G1iFSltE4rG2MAqru6WZnCh2uY7wTCKko0tYX7P05WI75p+
Ki0Dba/7w7LzGQpqzcY5gEDT92g1m6PIwwrHlhQ1w6oHe39t2fKm/9Z4cVj2w66w
q92pullmZIj/YvOu4Veujd5E5tVcsCVtei4w8KrQ9VWHAgsqO84D/hlFGq+VnqzY
C9Nv2tS4kmw/K7MI/Sv635BHsnK6w4vPFgs2CZ/tPLJSup8TD1nST/Pf2aWnjLdh
PlZMRaAUYuJsRUdeyKZR+bF4EEDOg+sqyhD+9zyzEdoboArJ68If6OJthOoZnMLR
DeQydnJMLdx7mCHNrlD6Z1R2AxGMTHUbYeQ3D2NIJEarC3j/gMDa35VJ1jQOjXlG
E5CEeQAY6zHbEwtdLeXg5UZR+kVKJlnjhdwKq5z3b/ORMn2i91VtiwF1rrAzKIxg
N/CYDC8w7DHTX02T+Dgzh5lENrjA5e1JK45HLkKtBn+IJxSTZPS3jTGs4NfI4A1/
2bWfTRqUsmezhnWidP8Iv2Rmvbu5OaU2mNYg90lWtdhMusTLgxIFbdgS8L3gwneO
+5EqwT5/UCXAQQCaB17y0b6XoMonce67YsMvlxiSsL5+JXiHErUTZdcIwIygoxvu
jqpAJMITjhJbLhXCkyPVPZk6t4/wHTtUX0g+WzodMBw4A3kkG0PoH9WzkvoQdZs9
WUwyO1rtilsV9QzoEm9/ljCxWSsR0JBVB6epq6rM5wJwJruk+L+1HoRUBBDH/n28
uzr99x+B5DrfRQysfBBT3zuH7rxOLC3K0P7zRfFEEtTWoAc8dBe3D9hUhu7vXYp9
FphhjB/JbCw8q8XhjHn0ODhAQOLrm7KXR8ZotgCq/v7b8B8JY6FavqhOkZRwzMn5
3hg4UKCj4ATwjVdV9PCT8t0tPT11Cq42XIQhT3tLO5U4rsO3I7yO7c4f3qgoX3gz
yuvGYv/Wb+mYDCXG8Xfcu1MFEO1UICiD1wjlNSyeUN1PLF4HyVKb1BlpKVcmfHo1
9Dj2vnxtrIvtx2GyQy4pniV4L8pF2DhTcnkVntQpnuxx3PYd4rIhvdnYfTFzX0dN
wxe4OE5TvrHxUpLuDLUQ+NmueKiuz+otW993NYlKQ12n1iojOp64gwvsHpr33JNq
`protect END_PROTECTED