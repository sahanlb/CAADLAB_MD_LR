-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Yvy2yvogGcSvS/QgOOgvnp1MA9GtIfSh+aY1jEt4HOdccXAAJqmfnYEFWYKkh3hw
E8mmng3ROztwENDgGS6SJFgG64FVlmqOxEd3Fkyy7lOzha/egeW0NW6ibynTbAlG
GSFyQfWP5q1xWScPyQX+WcET2duDKLh1IEGcstN/84U=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 29978)

`protect DATA_BLOCK
WKJqYPWtnIXpaxYYpXlqpRh8xsbEPvzazWMtDBiJ/9Nva2FmjBCTnfVAwyxbw8aE
OcdWl7oZJ/Pe7Nt0XhTbhAmPxi9LqyTP38SvI4dnYlU1wufZJZ5xM5CivvTKUytZ
5Yy2I64SqazZQ3bDymitGZktrVELrLd09wJfIS8ihhj3B6CPKZynFpIjkjh1Y+Gm
MrtOYtwAqjF0hN1Xqt/lt0O4U5D87uEO7T7lTVRLb6wjLX/TLjZc1dkWoB5FtgG4
g5/KwT6TAkGeXjTnL+eWhEyH10gCPNtVUIv7ZB7MAvuIa73/27oNIMYtzGd+Da6j
qvyAZQwFKOtfaFnC/+sMMidun+BIQIr6EdTQYhDAa8OBI2xHEz10rUrqIDsP9D7X
ItPs4NOS4AnUIO5D5U2KMJJW0K5o1ujYzaLvRUCN/zLnh+eBBF5tpNdpjVF5tz1c
nVutcz0pp5lg5I26Dv4GwW495ve/ZofVkq+BBJdzLQhR8aBSLpQgL9lpR4QULtau
MORktH3XEBQBAV6kYv1qsopgUIz3kSBeXrwGpgvHN2lHO+m2wiOcX5N5O3e6ILj/
8Oaf+EDfaMLn8elCsvrvi5CA6jv4d4eDJOQWTNZRkjToSdDw5Dp/Rf4zH0QAsDTz
h8Q02duJ2w1sBeLbFqZPCFqoRAzqt9CNDzCa9ytCbFPaUVXFoXNhaLZTE6yZgFN2
vUFAcryWPmJX7KcstA1zLwH9YNj12SlZXIrnjyPKHj6qxwmFuiZxVNim0CWPqiF3
JCtNOHl9ODea5k97Bv9cQ8xJ/5278b4IfkiO1WjSCOMWbjmflaD1ggWzfFTt86VR
XM/eSsbHgiGtAJf8SY71tToOXkBgYq/AUYT8jqIsCcdQny711nG1KFHNDR7qU35J
IYDvpZIxsWx7iu54FYYUzlXctlP01ScOpTDxP5PIkdeJ1OEGnQ9RMW57mGPG3Uq/
5w0E9PfbMpaDBOJFncnL+2EtClBvJheXH7Qmgx64q09qX88BloeUxWujAIoKXuQP
nOP+gFOXnZKVF5N6wAHoXgn86M5eEZ8B4fewoHaPHippkM+GCz9GkOhDbMX/xUtv
QjKU4Wtha4diUIYnYztxmzo4squRuvkw+p2A+LGn4LWfVP3WX7JAEY3Th87yLKz+
NyREzx+kjRW/liUMK017XD/Bjr93Gbwx1G8H/CAgQWRfyhJhMODdB/N8ex9tqmYM
EikO0PmwTpGup7uKt8U3V90z9Qbi5YoWZeYjc7tpgsZ3OOzMAaM54n8PIBQjkuCg
Han5vJpe9Ka0oTnjP35fSuql+qfMEJZOD3RAs3k6nTF+k8/IoUxqD0H4tpkfglVs
njYriinIw5dqB4RmNSKWHxl8UEronrZUKuncasZ+jI6B37r5N/c3kxbisdXnipX6
J1e+NByXB437JHnYqpyhd7uexdjxarnBOYeTfPyFilxvrJk8sjM/u/lsyZvbhTK7
O/G2Z36OElvHtp+YnUyQGNBxzjgOfdmLZKD26F8AjEFZrsGS6Y6eirXDwdPDjJ0F
WpEMB5Q0vKah6Vyd7Y8HSEVK8Y/FjXZutRz4f6MgDoPiIuhvDSlqpS3J1wUIIwuw
dwyBoTO3gg1Op0cQ3KtVEHGoomQbRV9ixDeUi68CKaazEDSeuAsFvhR1WC34oWHf
FRy97++DF767gT2sRESFDgy/B7e4dPsi/k9CyWmdywnD/yDPYoVOs+RZIxFa3Y2T
f5X1qGwd/3niXpvT+hvIf9pTQ1ICJUiQc9Ttmx735givAkKwMcvcMb+/656QPUz6
Hd4RbVcGaWvXthdsLRTTOCp1meYERg054dvUP8WRFncQ1qWmEuRswFtCWgDDf6//
wqzxkPlda0fdxKSpQKntH/k+SqdPvFkunw+5QC8GN3PrYyhWciLZltV2ogJvulSt
zSX8WWNHwqf01Hn7Q3/4Q12P1gSDPqnfufd1HQkokypf5aOrKqjgGI1rKqQ1pEV4
Q45DIrY69Wh4SyMczGvGZ2njnhjWKbHVI0Lsn4woqFzM/d0BYbVtWE77oi9f237s
REOeGDZtDe+zQe+G99eQI8nt9rSCcsXYVKhuwxdsCZXCqAr5ik5gcOXhYENy3GGY
oJpkm0FsA43IJmZADRVsRcVqRxNzlLV9hReEg+Gl99q/3xLFuLVg8mirCuBz+AJp
vvkLIrty0oaCE9gzUy5roOwBu6wNZzHvqKAkM0S69PtmCl40Mp8gSiwrQiHoYFj5
aox5IrJWy2Ka1P59ngIUMewP5vg6m48XNmYh13V1gA9gACuHfYhXMb39uNRlhmCo
fH5QEvU5tSP3SnZ9/2yTaQMqAcls8Xk5FrnvON9PGfFPVJHsCvDEIefD/L68Dpbs
rsv6IWaoYJW80z0YnnNbKNNSl8s88j7dkZDTwW/dRVsiiQm4w2V6/fNGNgdLxD0X
16mdNyyyPYPN/52AP5Xn9RJHsKEpy/+sVXLyXWHc7sLSuv7hXH2CQsxiXEC+EJ6o
dxLbdi9Gv2lrDk7gmkGQ1H8fvXlYWQGCj4LK+vtIMPmDpjUzt4H4w/blA969OglQ
/YSaljeOW35ULrXT8wBYj9jQ6Hzaxd3xla5orJbF1QYbVTiFi4BP/ZDH4SYyJ5m5
ZfMTqJycY0WEAtK9g6ZM0yex1JXXNqg5T5Vgbn0RZQG/66a0r0RxUJAa8Me1Ihuk
JNwS55WhinG1Gvkt/WfK+qY4TaNj0XpLFomovmzLzXJdRw/Wz2vUcw/mbY+tVKJp
FA9SZ6LFs7xSwnACUR0cTrP4fl2q6by2l4ZoA/nJtJ47wCEcoTFDd6krS9dI43Xi
/7PsFh39xzql+IAUB31y5LU9caj1biZKdGKXG/qUG21r9Cdj7xM7EhLA/wKEouFr
2iQS5ycTofE54BMOD8XIHTIH0i5tVgNqy3euxY+0QNP0nrP4HQKs5TgQyafCJfWI
C57Ofr7BJRDFMtm2zL1lMnG+clNnG8lekoG5bm5NvMFU4m8KJjkvVJCPM+iNJJtV
iRXT7Pbv0ZQBHOHmx8bO0C94kbaKv6KDqCmVstEDgLLW/bXY1ySj/iqP7dEbUV0c
ZA+5J9Nw29+/WkhXHQLlnn72+WR7M9IIS1FJTMxw0sZUgqYMZizZQJ+HWAxS0g6A
jI91K37Kk3VVlXrWd1Ce2L+0M+MXkFyjcUM9hM2Zk76XrBPNO4r3JLRuGCs2toUu
Zszz6unpLNC5Eofb01Q/fS/gRjYUsJnmDiKQKqNFCYe7hoQcFGy3Xa/+EZyuyxij
KPbUpapQ735L1ZLtHXwbpdWkvP9A94oB0P3ERMYCSRqHhgbUtzso1iVS7gOQu7UZ
tUYzi6ZtARHTtGhcKbPjuyD2/2Ct4jKcGcw+j3S77V66bddiDUpgx4Xp4Lk6DEtU
ZW7C/NCe28PUIlHTef7noHpYLouUseSRbPvP0na8aL3/Vr8zSBYGvxnYMJQy4d17
6/4OlEMlhgSWffmF4vFiXB03aTTxTP2OpwwLw+VeqiqjAd93t4Cp8McluVDfoeEe
VQ6pGtl3dtKy0C/5ne6SW2X/+V+MMmI092G1PVtd8Kq1KFmkfgAPy9o+bBGzxj7+
aMN/AMnjwnbYUqQScT+qEJT5h6kILBV5Uqoc5s/vnYFIbjEil1tcb/dSuEWTlqd6
MSdxBLM/JPi2bkgS3v8ciL4PS5yfl6u9dXkCaqAklsHMGm5gWaRXZmdPC8NDuDdz
h3ddzjHD65eQBVUzum6vN1StXTfsNVyu2al3cuuNrtBZzb9wQIFI8l0PQb9mqj4o
PDiQyJKRm8/rz662dBqzbU+PQQM2k/EjWUtJeQbapct4Y318B2nNTvKlzruE+ffv
zbWNsaNp3ioa6BQ9oyxwenf/Xq+l2QrvJZ1MjjKJWOULsIQwcWSoX10NexukXyPM
gaLheEZpqC3dlCh1YUgHB/zqMZ+Hl+B1b0/xxGrL8AkX9q6dWZUCedF9JqWGVvtr
FaUDZ6P/3hacJakoLg2x1Y6u7R6Rq0oXdVmVW331GZ9k70PbkXLg1bdcr+4oDdKs
8JdJVBLFeVZ1m2Clg0KerWG04TyWno3lckYlzk4sX/lwyi25OtJucHxskM710xf8
eiGjedpkm/LFYukq8f28GcmaHEhLUrOPk8sdEvQPq3BmqD1/OJ+vrFyl5cBmAXij
yvasTLOIsVKz4m8m4rPn9uPKlXT3JrswzDX12/MPsLlP/qIqFZof/NO/yHhWIGq/
OWcnBOLEWb1PY9H/NL9wLD73pa8rvfm1j08ZznITyrwc8Qtp+3MbvUbd4Zhvk0Gv
cR4cnyeUCI+Pe+2d+qmn3RkOMlFC4tWzwAq1I/pQGl1dYv9vwN6upIYZDWQ26UyH
r74gsAuUIXG+yES+zm76bPZA+lXlmh/eK6D+bybZivx47p31CorR6znTJjlzbaVJ
3X4wL4LgWLMnjbGWN3U4lTBTVNlDMgqLr6bXeV7NKLcaXKp76Qj/nBlaTA2/QHVR
/60JvDoIT2iU2OlZ1hwxgJY+ekzt10/QmtTxYKNPWHX7YO35V6GSdyMYmNCNpDOk
z6PwvKZSzMlrpa8vWIVugZwftVsVq5D0fyF2+q/fhmUu1Ix0I92l3i/VlJD7nX+u
nLU1hymjRd4JVOQ3OWwcQ0Y/BzKD85WDyiaBIIrBkwykXXmCEJP0dNiW8ezwK0Xp
+z7lFc8IlfbygbB7G2rDFsL/JeIGfJ2VODYqJkUvCCutRyj9T1Mgrt0x/62d3qyW
JjfRtDYechrB24WEqwGFVGwPly6Ub+Wyesdsno09t3z5WjP712KHyUvTf3SR1K5N
XMqUiIrjgXHyzUGldpZdegbk+K9C9wpCUq4T9wmyCjhe/x/8C5R5wcMAThE+5fV5
1mU3Cu/KIx4LELQAxrJkAB0lGSNfuKZymhW6jzect13CBvat8f7l9N1PQe2N9FCe
35lnHB832GG0LSQSSl4aHVGYrduL/24X2yYOMbCVun1vqFLjijxgfJbX71/9hMHv
9tWfQutEkGimlA0MB+pi6YgyXpnrheiTSt7sbD4a3lOEvLkox8erO6haMzfjV4Bu
Fm8MnGZPPKzOZi0+taKM8sVc6AHvlPUjvn9vBfK9ucv74aC6v6lqmA6qEd7YLqT1
tPoNlvKBHaVuJ7jk5tQl1uDl7DuPqBf4Sz4nanA7NVt5+2tG6/rO1TVeDwAxd6A/
gexEaKfvz7IhfOUhpIvQG2dbECdxh5z0HweM3SIvSeoxxqRhNLH29BP1WYVij6+w
xYSYU8abOz3+8ZnTeK5G8aVJ8bN7mhD3AHeq6zdXTR4ih7kNbgwhGAHXtgCGp9I+
T4APnl85GzDgqmle/c+7aaC3DtD7m8NZo20DaGOfCYJcqHYLB+z3Wdik4NEKcKw6
zUy/3PwLwWwU4V8h5ndf2oVwmspIKszy4OA893FnJplKkuJtIZ0vFlPtSjBnI1gi
w8TA4rgOooERglK7BAySFlWs90DmyVSH28+LB3/UMFsyszpc4FNs5g0uqlZKUd84
8ksW3pMpT52h3ME0XFiJ3MT+N3j72eLuZ3/aTMITNFfDNgx1kEvP9xb51syI9vLg
HZ3+jI+4Lpo4gjbMML+X0vj/4sC9VWSbHiuWxQgAz4BtdacabcFh3eEvzZEe+DJX
cTJOFf9hO2nBWvEZ7qrxYktkGBuV4SeHD1th+w++YV2z2X2RW0PC12uWUt+zwFQQ
5O+OkpA//f3JWYZJOGpytYQcAj1zir2WXZvn0iZ6vBwxT3tv0bQVzjlHze++8zku
FuBq8alPMaMsl53pyUL8yUzmUOL348NfRsczOQhjFmoZlth5CeKRGMYDg7psdlyu
cFrIHVq3wAdU9uVFNexhvm2Zb/RUquIsjYgaQOhMCrWHMOKwXnZbFivAiV3rBlyB
K2iRuGLqmIA9dxszqy5A2eGTjf2ugIgMcgMZ/xECURQqD9GpjHDRnOfCBAnq9mKy
GXsCCJrszFSK6yCWWVgJMFR5iUMHh4wnNgz2pnkpyz/lFTcMxg/OgtVhNxlRz59P
/HEJD4LhbohA2kTd5Cn44YKqATOw/CpEQD8WUOv4p21/cbu/Kas0/PgsOKDsEdtt
LS2nfuIp9SSgExyPcAvfL4LbFNkAgSlJ646BBtfHoUNB3/A9YT31k1xwJsXPEnlZ
a3TnkCUAWTPGHm42jqT75ZuxQcVs4uhCYPKXmjX4D62pvLxrGzo2Lt3yTHa6Yvbw
DKjg/Nzq3R6KP4dEO6bcuuTifY8/kM4DN8M+CgGucUb/Xkuc2i05wuHnIVkm9W3z
tFuc1ux6HcgBsCDn7I+3R8537AXpmPya0TKYTJHwhYnbRf6L5i+ppyItVvXyNPq4
v1BraBi7aWDCBCpRLGFl5CKPH/morGgYDXyFCLtZDQlvLzenIN+YrM4Ko1XaMZSQ
e4p4ix791UL2IUAiykV+utfWuZtU7+cHdzACUeZAxPAjUtIN34/xxj/9jrLJJB84
59cM2JeSxCz5el5Lko1G1VaY8mkMDKPV+WQjFPgUuvWpQtC6rAOHI2QXe1pFg+VE
Q3HC6pnRAr3bSo010xT2BB8/HTpCixE+sHYwy+jpQfvDLLAhrTt575QOSws1aolM
PiyQxT9zMQ1mEU8kfYCiWzip8BINJYTjipptuJrnBrM/zqhxazFzDdJ78s2dto2Q
i2qsedtindu3HBlrqJUXs4HNHrZA/UOC16GGm/dtJJGdTqoyXezi9M4kV3w2mI1H
xQZKjM8UvCyZmHRg4/SA1lkixWiWKoZRWautXB2UyFDRad6mW/p9l0wkhBG+feLq
Z/maVqis285x8PgbIP4Rhc1/dX8bMU8MTz8gBE+spVwYLeJj8Cn6DtVWwuVuWSLC
ILzfNaeL8HIFOE+O+CVgcMSTlLkyw/6GwAZoRybs6aLra+K33QkO/lYiCmdoiAJ+
8FO67EWQCeUwx/yVSgIms7hk/u+xxd13MfqpvY5pOj1kG9MhmdF/+0LQ8+4F8OYK
gbu4QeFYe024rLISFPcYAG+ybVD6Su5Cz3U0QNhbsiUwNAs4yJWIMXzfNkr3/k5b
mLim4psO5koyXF4xsX3c2DCAhqaq4a1lHHpSjJLvEiv/eRsPw8d5MMX1WvDmd4D3
5r3ONZvYZ+zUtxs4XowsBxn1Elb3JnUjrxjxX/fVN4JGRZmikBYXTLnC9zx1d+XA
Ri1k7ZRQNT1OkZ0+Pk5PTO+VE8Ru1YMTX92eeLM9wSp+NESs62KArrNH5CIwjFjd
TYVUd5uukjTLzNpV5i/SKTTP9+RFTHj2m6J14GzLeE1LUQlcfx/GfH2geewucmb/
TNiNos12Fi77WpEtOshk6rXeOq+S5ScjZJgXObHOg9IsyDn/QJSIkXE2kxjP5wwW
inoB+squV7l32nJtI3IJQQouBDnfUfUB8ba8KWQkWYncb1Q46/xJKOOy4Lk1ML4q
qr+jMNwz6A1mcfhg1MBUgz4XJFK8H2iQlSuryWEcbLJVeAMODaMpPsCNSOPgzxUh
EbPJnLhTIBqaDYKwGZOV6IMg8R7wJwx4C1kyRn6JkUpG7H/L2u7g9XDF8bNr0po3
SKOMTtIya2o4+gZRRC8O5yDtiUNqM5IVAnOu6kk53shB/6clpHBbayWdxzjYL45c
06VCvy7DVWKwe+d5EcPAkE5GaJ0fpHMhLcoVCwy1k4oZOHAWTAvIe97L/XyNr25N
CmPbMcCZlwnLE+QilrmsL/JDne+8PBPlJAB283ZWInT35QIzGlb4Ha8/TW97e25X
xMhV6kUuV//AWzXRPJARQDaJMCuiA2EHXd65dK28Zg9PwEJ8ZmFd4GGbMlyovtE7
eBGxW8HWGMdLVjsQ8U4Lch9p9KJ+W1DL+CtcYjmdxjwiMZ/oi8Sfbw9x9SS9LkqE
U/BI6SPpg2UfcQnKiHLYQjO5bHR5JlNRobpDrRZn4AGB5t99mlWohrEYnLzU2Tir
/dAcsyz6bEGMUgBuD/vEKN/9NErvjjgzF0yNkS3OLYF+BS2mwnl0frTk465U/0LO
gydJ5AGmsPeMMVD9d2BlMn8LwcgvmtWF9vRdQGO9xk7hSwIv1HLdXqgzPDNVf8hR
yV4C+4jzFY4CdqKh11dDgJ5y9T/vfn5TeoBvh/jnFRXtZ2BJ4L5xGxQN2Rc+hFPi
eSweurVPzHijBPiJtTsnks+O2Umt1nD/2TT46qx+YMeyKKy+U/I7qW61+arR7pwU
gR/+8GHSr+aFWHghut9ot3xIJcfy8ehqPQ/A+5M0V1lmICzgb0fUAWtq+aSwupc/
z3OoWTKy5hg8fzxd+ti7M2z1gWvvHmn/EkCSj3CGfUix7eGIsRmMv8sa+duvSeAe
xFUEpcebLNzcr0OGHd+PbJnbkc6aTRmxUUKGc8hqWqDVWtFLNwX2vAUdJQXJD2Pp
VGhLt8II6uOfEJmWZKieQzjndFjysyMRzhPTp/V7cPCvewGElAjszPNDMAu8GkHI
EsJNEymVq6Yz5BMgrY6dY3BA+CsslK6LZfm/sTsGAjgtNh4PhSK8/c+r1/vQrAMS
ieWvXvGeJNFC3emZM/pazYnqwzh63xBra2UW3hUOIQB7mzXb7z3p9IaUck91j04u
5uqDbXb1vnlTRNKWFVg4eD1ZmQPJIQaXvjtV4s9flTrTChIijBCV/xR9DkbSD0Pb
uwZ/WYeqRuw4uNADIPgR8uiBSUzOOu5dic8btMH/f6E5O5qc/fREBXUEf7wirnPq
lAP9OD0nQcFivwPyMf+kgIs1azwisEJbJ8LXj+7N5zjLWa8OR/4JJhNhqPYjp7aU
Q0FFUMRzke4hNMemxCA4rvWFv3m8+eaY3NNMr/FNk6f90dURDcauS6EJGo9WcEiS
Ravolmdb95D9vKwVbjXhIuF5UokBXR4QFEiyxD0od9ri4emBog0afykw+0rmyMFN
YsqxQCKGlVITslN3hvoV+JyeyRP7JpSx8q009bQiAuxXAU28R2+Yad0gG1M6As5N
XWGHL5AqrVfc42JtsSdcfngMjsHNJQsV7wRdzqIAK3SzZQj1l8UjVKpHly/lCZNV
FlyE9VmI2LVYs78SRKm/nK068UJVnHUyfwYoMpO4dTwuw0jiGvMkf3jw8eX0pIU2
G2CgW6MI7O4gKE6+/l8Wxej6jpq5EeLewTf4UVnnEb1T0AuXgKQdoPmb22fEc+Zy
X8D8+MK9Ci5OQB0a49DBqxBG65KK30kPLiOlsHWgO62XALcE/3J/Icxi0AaSwwk/
Dk3VILm390WX/6srd8l3tlplynQgFJW26opul+3ExUEDdVN5Z2uInnSyoCAv6gc8
zKdBS9zdIh0YXeQGHYpVzNwyLtrT+NBLv2wLa7iBWRr39jVCwBWSKdSq3rWyIkA7
9gNoMZffdq1gn9B2OclPzsXPCpnZF9ORTTvxUY6q+oKmrbm9pUm9YrRGqhaZSZcy
wKkPLCw37XD22L11dO1yrbSwglNoZfnChCDsX6++zVRiD88bZqoY3M3qWlPSpKY/
Cv9rI2gBdJlWQ4KooQ6tPxIymH2NG8EQCLFMNaJKDA3wp4rTm7FyDN4BG44fIq92
QNmmKnITtC4VRrsXDq1hrN9dk9O4HUfrbynhKPToYOcVlhO2QwFq5NofnOyxr0Rk
0AYWAcq275st3kyHDc5+7J50S3PefvSsaaEmAQSRkcEAfr76/9/fA+v9Unm5KnJ6
oQr97h0dLPFpcdADF0e5RPnw2iHUGBysxiwj/UoznGlO24fZVe1WlopTfbUB6Umu
32FShsgFlsEr+b+iGMJs1anUtWroQ2E/VddN/2Vzw30a4rxJw4wMdu7iNFHD0acP
LO1JFikdkA35dj4TouDDO/bW79o1v1PBPt46zKBtdEMc9k024EOoMmbzWE29FAmj
JucZl0NpVPqlUcCmELO+cFKoZvoZWuck/v6iGa+q2HA96/L17Jne5jFm+FAgIwEE
whAMOQSGNb66u+GPu9MyrBdLZaVATf9SrEf9R66rhPo6HM4nNcVEmsymwHcxt8WI
KhV7WgOsqU5A7lPaQHD43SySniQXKPKkwKWlWY/VDcoZ4FYcPwNcDFWJCc75s/yw
IMSKWqGFGPGKGc4lYKhMlK1+sHKvdupGV12ccGCK8IwmCCDCflyOqoreHw9KQhWH
Qjov5gZLTzPAnEhFXU/WTMzsUTsluiWVfjvhLJmXs3YgbrL9wOBVjfz74EcZkUHa
uHJ2gumxtISm5gkfpwBWeyx0+fRQLHo5PnM1J1DnoO2epcs+T+d3RrQx5rr4TPxj
dpnJfWFkBlt3nD8FbZs1P9Pd6QlD/ajY4di8aui+rukoeSeywYdQHfJzzqFRXYf/
oys13rGDDuZHb5jHsV1ppDAcaRJkm8g4ndpcC27vUBbEwHYun4OJjbI37+HLnlCF
9/k+pg1aWyduk5oWOi6IfbW3qDNE/uqXKHASVTxHMysOztDtVOibyQVTWqe+NjjK
rkOyS5byuRItAY/VRE/I5/2kbvif0OVAUL+g+02rGw0n2dGe5PIaG1j41kn0cPLa
XqXkw7UZkSh1L2N6Q4HtxxrBC9kv1trrhPgnbjsMvygg7NgXeFzXOmgO0zJibaKT
0Aqdl2P7fVtOgtbZ4mikR6515rsYezC6RUJJfBwJUgbacs/geIGN03yBCsIsEl5r
rBUiT8RW7xBvSSbeCk8XaTL3LuOkrFxA7mySmOInd5EQZ+lG4tyzKFlULo4PZRLb
oxONIqhlpJ1gGqdIYDS2QP0QqXo/1roMt5clE7ALTlvfNEduqAniXW9kSHX3Mb3j
ji2Nhsun1L+eF44/p86brtYLf9nSiAAk8I6b28B1lQP0oBEN5PdWt1X3v2gGL/2U
A4FmhPJwWKjQaxZ/3BOsVxmFnAQCmfbAaZUo/7WOA3Ia2qTB+M7p8784h8zKhkD5
4eJCeNEY0wp0JFfsHsH5in4nkI4y/1hownovkhKXse1X0CQk8cg5mFr6XLOmns6H
64ZTBb86pHr6M/qU5/9n9aPkbCuSPahXRAdLS1wGpQXeIdFXok3kSNq29oK4jpJx
a3TiA/zy1Y3dEQrfKeWkENtmLckItsZuEDmxfqVIslFsNRMO+cm8tro7tvq1M/8f
CQOoco7UbcnYYpRlRDSNBzX2UDM4DY1lgce7qfaFXteKR+kbCYeyDDfsB1FuydO5
967Q93XQm6J/xHyKY4ucm+V525f/0cQiZejTsXm/4U8n1qj8+YjiVFAYkaJ6I3Gz
SVileETH3QIE4IsOLHB8S77TACDLfTAYri+qOpaqRbairZjDGy67LICR6qGDymjV
XL1fEB2tphm55tEdHN7Y2tUhnO7Vv9GrPZdTjMWNn1VInVBNS7Z4xhRI/aLau0lm
8fgTK7pq94c/rcgjMyaAS19zFs5NUGFmR0IdaaXHjqssiUYsmrSsXFYmxMg4TfCd
XdgqMhR9LZZ9E9U8Nxvgn5NAWlBUREJMi5jsox+pgcwgD22Sawr0qGv0cVHorIcG
GapXfX9BWsxFCRftBi1f8IYOIOdMzLucRwzZCHH9TkoFLPXzsKQv3Bl0ewsThFE2
n6DiLpTSMLIyLHfXQUZCLuJsKAkmmQcis+0oP8kqMj1xvpRegd5e6QnhRRXciIxq
Lx9xHxT9oUtAzX72Q4Izqkmu624mAQnOaVrzHBZPWbt2PkvhqIBypawYcCo3vLLL
OYP/gYNefiHvntG/7ucJtnIIF7M5spBKNUDtWGjWBGAho8QnM9GJ/feMfTMlhSj5
4sNZuIxKuHJ6S4TAX5OCU11qle5KDqwddbvXU4szcfn/3QgMyllHzJvbhG4MhvQu
PG1mBuyWW6BDStBxqTBjeEVoC3zvkyLTRz0C7YwK6+IccBBvju9UqhP89RBf5COs
R2HKfVM83XK7cuK5qkHTmpbB8gp9WKwR3UCstc9j7g+p82H2CJspyeco2cNlJiQz
Rz/K/vmVUUAgTrBHpijbtMvAvYStiGpZiwtztfhi9/TY6+UYRKNsFCxW3r0Tclkn
FixZtqi2gt6/S+/7J4RQnggp1X1JlshzLI6q2fA95xUXo68RI1Ooy6C+hisJ2XDq
tkW+X1ZnD/OyKkZJMitSFK0YcYsxESnITdn23GSMazFcwcU3wlJlcAKSDXF6xCw+
1U+TcD0uHru7KS3GDdPK8f+PJaMwdgkzvecwpIbhMRYyyaQHjGAfyzGHndkvm7K9
zS5gLGKtgzZXXw5ZApUdqqOsTDOldYEa04DFwWtHfKf4istskhxvuh4TB6xqtc6e
RvHNEj2LLZnL9WA1ayX/cMC6FYtazGJOsHtoWcFYtTuLZ+gonbAEhyK9DvwwKPHf
yb+bfeQnaKjVNn0Wo3tpxJQaSO2bA6+sZlPTHD4u/ZaOKgohWXY5xoWCpVvHahvY
4P05sg0JPLbfxdocMmHth3HcRUQgNfsAwEC6RcIIjUZVc+zzNYA2GFmOIg5ukHAj
MJLVbYVafipfrrjswgi7ZqAqxpwfmYRroa7xfTecXiODZGdTMtK1XnLmL/njak5x
bsqvIJj3O5hzLpVZWITboaWlFyfXsLs4yvC6e0XCihw7yV8d7I9+UHg9LolSW/hQ
5It4ggJwdadQcbNXZoky3jrd37X72I/z/n7r0tVfSvR0nI5jcCInpt4HthqpzUnx
/3nk/809BXfjK1wmT49tl6MQsJLlk86U+OEM3MPzpqGCT46H7mrDErnL/bAfwQyj
US5z3cysOyxrs/cKANZ5AaUWin3NWri+9zRut5ppnX92VzmlDDW0PpEY3NOOWVP5
I9DiasGJHosO9OZGldAjXlGJb1ztEnIi2Pd5HkcqcwpP3mgCplN3gg9fZvvo69s6
LY01+DDnlxRRaDweXp1qnR3nahvi0vqxYy32atn7xSYaEBkbDSFHDQsMN0rbY+kw
6d2/fRQwek/W2Lj4nbxpLE6ynyDNmf8UxcNfWL6aRC1p5s/R3isyi4fyHU1RaTPX
AevvZ/g39XZDIWMfMn9MGFSQNvNp5nEfwxMgqYgtYsaFQ0ZqFdcmlkbPAxvkdPNT
nnswQa1pWLy55f6r5j/yqzZDkFiD/lcFoEhrfscJnO1lN+WtRfPhPoWSbaMdeAID
2ZI9XoRuWqULUano5vtELH4kUbJAKes1WK3xcjtLNVmg6bfAI+ZNr7i+ChVTt83Y
pwRDJ6KZX+RGBv1VLEMesuF3jJIKLwiTUk83kFrHxvHIW/aGuiEdrMiGuZx10Nep
AJEFktEx99vIkAoZfPkm5/TuqQKBnkx/y21aCP+SKN4k/RH8WyaGKH60uUdfiCiJ
wDxznMPsggg9JXsak1o2DMGtLsG9xIxsDXBJhqFl7AjCz3WLEw8wXqeA8+YIkrkz
06EWQyE+1l0MdfqIgKz+hIxph65TQb/z+zBVAEVLnZoPT/wezpe6VFAQyJNI5LIP
dY3aJdcW9eaWBCSmxkI65tJzv/6XVlj4TaqTlmfNgaLHYxYQCeBkLcmqbjUsIdZH
ubBB12eHjOZqjF4lOtiIlgRQ8JqIHLFfkqcHGcoBxwoioGI3B4UTPLMoAZf/wO/v
TGU2/b0T/poi4WMuTJ92XegEmzjeqPDlPrz4vJZh9NxLV3zSK09V8Ev8NkzH2jFU
BHqIPNbOiZMTBoZaET/cSz4LkzO11fp7eDrrA1ujiyPjewgSw4IUwHv8jqSjQlgj
mVOT4cUn+BMKUk9+3PwqBJwt7J9M7sSbGsAMSbBgUMpbgpeYXPk7RPh3d0M0YgSc
HiFGGMBtdx+ITFyVTD/+zelScBut6tcbSXqXo1tuEiHSV2SqwPA302B4CWqsYsZk
0ZS3VSoZb7Y+DOaWV1CBgPY5NZbyIWsgymbwBsyYW7/w/dVtgDic5msEgiKsRMl8
AwjURtkvNiegFeRtzdvPqfBOl9kwN9q+2001LXyssY8S1aSb8vIELwa6DCieGhjr
8LpBMYYCj560UDWx36+8HuTgoL5ruMdHSnwPoxnGyAo2fCuJy+hII0x8Xa8xfhnu
t3cgLOmZwJy+Z0C4Y+2fIoVpprNfqpTuajZI7mbIw72nQ8Dd3d1KDvLq/4RrSUvL
T0dYjDyKWItiLG3wdiYD8PoCUB8w5lNO289CMIviqAWNYdiq/qtEVb6wFMd9LPLR
o/PbRkkGl4S+B7KOGcA7BTxMfto1ijFP6ZrF/GuvdMlFqyr2on/Ccz0wot1k+txx
Nbsli6w7Edx17LXyn03QiPEOecGZNnZwZP/TjMlrHTzoNefysxZPy3BTG08ngBGV
AuZzMNZvaoML45a3Rn3BxHOHkujxJZK0N8tiYUOOk9tJ9kAfF0+awI+OiYujZbVU
FPMDJYizqcOw9+FzXq87CoaquKBzymd4fA9OOKFc+gdhPJLrNPyQ3qxBWQqJqAQZ
1IZgDqmEj5RT5+348CdYAiA6SpCYapxE4wcnJTZsUcKCWihKqeg/HSjBN7ljGhUu
XHyoZifAJhIc6JVffi5a6TpjdXx9Fdbp0oPmNtDpPzuIgDImzMZ2mhd69UHDGdok
+bTkLarGbsIMX8p2vK+fD21x/aRXRqZ8nfENOIjy0xTCreSVD1RvVUIQ/rffWZC/
YbJsdT7Yl1ndx377tRenyJBgTW1Wcu6YZ2xS7med1Y3u6i3gr5fmgTiGyQlRFWIA
AvwdWAk7t105L4tVH2AFYj4pxCLc0lkI65LT7qGByU2CwZhSjBuGlHfdEMNMg0W/
tPpFbE0lDCQPHB1R6dCsTn89VWAAgnuT1tGKAtCXcndcmLRyQwpxrtSurWwfhKQ/
NZgVReTMU7W6yBMQVdZHq/yKuo5EQrqB0VDb8p6Vfy7tFS2EXT8/R8no+z/6YeH/
2W+kHbeDr8Udbo8rrrxuk8PE2sKLkeRp7gi02lTKwYax1SRhc4CVqa/KfiWq4xLi
/teqOMHkhFAxhphkk0CAOpsHsfxCNVd7AuzuFQBb/NZnjlE7zPgM0cctoYI/w1p+
kJr0hKpTgBlG8RJzTpzKNN7Hc0ow2SqqG2iPon+pi1tVODu3VXhGcjWqWl0D4l0D
tASf+xfaa9mtxqQ0uAu4AfE9mf9XfwudAXHx6mJhxUyMAC4aOduwf/zxI1gsjQMT
0zMP2o6cohcgUubN3/pJHVqZIuC/wCQMUGitHOcjnQt5ys1JurQws9mOw6An8635
ZjNC59JkoTK7xZWDpHu3D459c8DNflK6MD/BaMNeCSkhknPcx+Lw2g7OjLJCqLSF
162VDvY4L6oKYTdKOW5jNczibJ9hrg1233Zsh2xi8zK+XFqgYoH/KCrjJfY2tWKs
foXSeXy/WAuqzASl0opPMCkeAwecaG8V7ymFtOI8HoLKJzrggZlEhEE+vSpyWImP
4CUvpV53sct++OcC/BMh9enzOw1q4plkm2fBDlpwafb5XUntjSERv1RMIUBpAvdG
zXjRiTLTaD543QSDsWhl8KQMWCc9iJUhi39am4Xniv4pzVvFXiKsjKwkkSpCnDQG
IPi2k7ifgpHzCI4WR8XQjmE9lF/SN0pG7L98qtyfqeOLLnfvEaLciYGEnGePjsJY
FPf6rW4xN85R9XqNOSlV/Iajwjrx0SXG1/ei05xYQLIjNBTxY6fUcTBkS6jCtQOK
1z/wNLnR7LuzH8kRYGlObUHGH3KvWmrS6Xfh1DxkXGoUpZolkdn/fmDQ05u6/vFo
AUrdBo1ALUkMAVcL0pA3vlMUtPIfrnN2iPe3topQF2i00rMjqL2b/OKFviGWrwlb
9IsK6Y9ET6j7gp0hYT/jM12NhPULYss/8hTey3c93yIuHMomSy0PZJAmW3e37adS
aQlL/DvyANn8iNzJgIOWVxPMcLCBSgXVeO/kudnF4yenBgRL0VwKuoRPVQ8zlGIP
Muah5Zkw85WawH4RTfLAVNLaMCSzv55/KXTGpfQMNDPFA/63yUSaz1INnXTNHT6H
H5oAddUp6wrjIw+9Ftc6sS8ewZBcQ1EC6wZZHlBP5RkW9kvqZq/vN26bmdMvwLIS
uAqjgeDFPEh3bXeKJgo3uNrvTokBaxOUbsDk8mP0NZGkw12d4QgHymRnzpQM/Jv6
j8ydTR3fHIyB91c6GSFn9j30kLsT0FZb+BwuLEYdUljbXrbEUj/OlTOm+fSYX+jw
UvsXfPj+xiOELaIfisJgo00MMZkyHFrDp4pYvq4HxSBXoKu30vfmjNQwhmsf7QDQ
U8cfVrKF715a69uqIaK9WCUn/F4111W0zfxKfbqfkS5chBoDWw400vuPpw2UlRY8
522++bWZM8vNF/k6v21M9XQzxGygyZYycAw5uz8vf1dcCvTUQIeHINV+yA1maJfq
mL9yfnaHwsQweBnQRlscVFwF2IbcHhi6zKR0Gdu/5aEesIfTAwCvjYw0l/I9Df0j
HW6iXs1gF2IxR85Z/ZtG8rU9tFxqBREUOlcDMPLJ5w3CtmK2CRk5VYH/guq+4OCU
uKWbWSWMUng9I61bLwUAZkeK+zjqk5txW/obe+mohyE4bS6qcdV2Djzms0bZKuat
bRb/0yqLfaFK3dyhFiG4NF2ohd02W9ebmGyiEjQRMslcsF6hKow9rPcuAPs6PrHH
79/UczlSIEBcBiJz4IfVAvSuik4RO1mQDKNP2dnPDcMnd92U4XYk+InS5s+oJchv
inTeFRm8C5cgZfXZrAuHul/c3EDnwTOQznnTumUr5qVM/hkiWrlX7ImYaLpNLgiR
XO4DL4yG1nRItACeu0NOYcLMBtMHEQmVgOVwjXxGYmoJ6lG69Oy3Q7OxM6oNeD0B
DNJ5ohQ/EPD/ppRnARIgrcopRrnJsypZhtoQ8CoLRz7vau65bwybleFADNRYkLai
UHTZLHiqLvh398llZqPnxqGlF5479yRXt7KGE3KE8O6Jw5KYHmCWTUlKdhrpTg+l
s9J/a7DS1xNBo+4UKdnYxkapJLx0eVe3m11z7qD6QpgZWVP+clnCaZ0qxPSpjoCP
mWNPZhYqe48OgdP3uhBV38dWd1RPyfNDKZQiXpiXsIBvcJ9SO7Fnh1bAJGejV/br
xf1TkTllWizhuz2kSAoxywKWL72c1zIbplSTWnyhAxorvvr+xFttgliKxqfT7aAs
vZyJ51jn64ptrk5AjszhN4GbvA/hI0BrhoNZsSx7/G2rphlKqgaOoCf6vdG3msKi
uhmqaLrsQjJF8Rl58E3Xh2I9uib8fzWF9RbpehTussxTrgyMforJ6PLDZkyweRO3
ySeohguFyVlYIBoN5Q648rNHOlNFOsOPONUge5l+kgqMv0VULEPqJAOPhTeh2N85
gVo2UD6wRDqvkUzxC3r47RQhp3HjfxMcHVVwsyS4nabT51AxYOIUJD6aogvqrDq4
JB/TFPOwMhaKbkgVzdD7CS6Kq/UPum7Z5rWwTLGXsVulcciZT4u41thUXSAVTMeB
UJgKE3hRW3lZXqth6lf728Ohj5yHTSCe2JZJQknN0vE0KdsSa2aYP0nUa/Ln5W2Z
ZkKaxWBmaRMOZNklMLkuDsrwXCzJpyd9iHPfYpmN/MDabw9W4x20gnCHR93fcqPE
v/UECnVK5T/PY7hAAT9xtIyrJIx989kvpgRJjSoxuQyRkE70BRCfUXhfsmDvtt3O
pExx8LBaoeSmFD2nXQUphpTd9lFXxCiGsm9iMZW+/7y7n/j/l+Q9UfACAZ7/FCa4
oT5ceSH+tjboK8IIs9SMyUAjGAxjyj69hQNd2NKpntUKVD1S1/nlXlywuk/V9ET6
Vh84Mmq1ejdLOGiWM/e8ynEz2rIhbTkfhGhCWpUiSIecE23aN/trniO3lIs8cE2r
NaRPKWndGK0LM7FkLAfcFPNt6mv6FrfA3ghZpyQOGWvR12ShtaePZIjHL8qKFPAb
9XrXrx8h+JTytyMqIDwKjw+BA7sO7EYkw4HyrZjsVDHynca99nz3Wm7ycwmZJ79e
HygN7ym2GgTLuIYK9xT9azDvSEWLx24OHRFWm1bJQtxlYoyTQDnclkwas1hODxDE
JGUAC97VYyGF4oH7im2cBpKjP4pPzF0m4sqnE/bRsA0Zhq0oOGHFdplNUAyiZ2oE
meuxhAxLf+JvgtK2Z/0Ktb8qqPCJ6/mVbZihCifEhX+X4+bnt7kkm+Bc/ACZs8TM
rNEtfzYC4F7HXtmFFk61OtbqRO/wZ89KjKewTDeS3z6Hu37SUyhODIB2rjJShGz5
g7RKqo1Z7eC2ruSAUseG7HVedilI/BiKJfgz36FlEmZFCWW+LqpjqiTJNZs9uC8A
VK+1qDLYQJg73YNfkcaEi3eiokiwo7C4Su402I7axOxxtebKVaGOPhIRu7ETzKye
g89a0gQmu6bhCSpl52IU38KQ18LWophgWyyxA40fzXIpMcmODNcAjavOZBhhxcJi
OFEXzBdiGiYfmYeom1Ph/IRKykhbajtBl13+YJ88H0vlPJs3Fu9wr0d8lrOSZkdP
gN2IQgXF66FflQTMl4JwBwCegFBnuk3R92SwqZih7fiX3W1LxrZzORQSj9ma55+v
5RFfnIkJNhAQ7FyHoOUNL7QzFceHuz0sEdFUK/9ZpbIfnItH1GCQh3mUjrTVmWjW
m7+qR5XSo4cW17UgRu/qgUA80Zu++TLTQMKUgVz6kiLlxgjufpgOWJjyP3sRKAbW
2DUAQ6XU/qEmcdaR1vy5AIHL5C3RJCUqTImhqDDJgEB+Wqf7TU9SA/pKP0nk53as
qqfQrO1pZ4/i6nZiBVbODDgraIZC4jsi/bvhZbNCmoWtnlx2F5Lz2wKUAFPA5o5U
RGSIkYeRe/2IMkyONIZWCy0SzkZxSndDapTPoKkhWd52fVSFp6owmDWqIiR+yO5z
Wg51EDGLh3WFcU93s8GOO+6FSxg1rLs1Wdqdb5yuNl/Ywc2yuG5R5J4Ann5agaKA
lLYLQXc8y4BT/I8GXslguLm4AfzSeILYEfOvC5qNpDhFOHPHPROVvErCc3XlYuBv
oCB2VmxnHU2+t7ZD9Hz0qERIEEoq6OBdtYqd93J/7wbc9DWR6F7sqMqq0E9xVB/M
T++IohdwpPoWXkZD7O9SW6BsTg3Lrew4P4cHkV+7bKkP4b53g/m8go/vTerN1/QU
R00xiLeNjOM5/w0G2/M3tLZLisTCBpntj6TwhDZSHife5cqkdtJ2asuylR6dKcOS
1KffvdDUYPOTE3VymSWledeLT24UQ/bb7DiGAqvp4CStkOwPLb8nWrofuaOS9Eg9
BDjePXwV8wNAM7Nu++oc4gXgUJcEw8xgzYF7iYfR6JSG5K5iadggvlQALnUBhIwE
x8OtxI0s1AxAB1rco7+ise8oK+06tJCiwQlhwUSVO0iMfOmsB++qM3zB8ZKZPJeS
HBInYPyjjZN5pocTgTiJ+Wc12zuJIXHG88QlM1Mdbg8aQ1TAD2tOhlT3booU6h4V
5ODjFZVO3kyJExg+zKYbdLJat8HlnLNtNdrDaW0NLSgM/HPQCgJ1gYvmTaKarQ2d
L6IyRaC+m3emHVYA9KOXQ47nWvNSgXCU9UjlKbm0aWiBWFBy6SH5ttdF8Lkxd6I3
Y85nsDL8TLWf+svBZpueJUGl4oEmCmoRKFIuYdLLES4Isdn4ybThJJV1CtYckTV8
MM1z58WMm5ek5u/i7cnw9RZrCQdEJcKb4CMKfeD5AtirzzB7kHDf0gPdYqG8NVC3
9niQfmwo/yj5HxashvWOVxzsq1uh5NlHPOyTuy9Z7MK731S55E9do5IXtxjzZcbK
gdTQNaoitpiP8F9pfbau5qvFgMYW20ATvl6qRoxJ7zXTqNMf0NNBy+9ML01/aI2i
eGaW0jTcfo06w8deSdUWnDAQCu+uz3JArw8sBhYExZdplvKsq7wAnusEROwFF3oK
mzBL2PoJ10wMrsW/WDUhnphPEWZymHgXt3W6gdCe8r765kxbCO7P8eKjWRMXXmUe
ZDCMnFcrkQKoEm+gS/Nv1lpFt0l2utUHQ5s2dWRlcf5SfjwijCI3SM7AzenZmkoE
XLeu4SmhCbPv8Yvr5Nl4n/n+qOI6ZoaHUKfjNGIrwN5/Ulm/RcqL5SJgIHrLzHVS
ok9/T39u73Y8aKRO5gi0sOMTWn/G+08C4RoJEbeHA8jf2RtA/6zNdvbJzyi41m4+
MhDcu/YnMWbFMPXsOsLiFQJVtG4DhOo4qnOjesWb1KqbaRYs3RJ3WzqxzKPMuIS7
YKHLpB26uBW/bNA0n8/5dEu0U790hXC0hGaJ7NHTGt9e3PXyluD3rfbVG1iKupjv
tuRhqE1OdnhjZcTTqyVAKkMYe5A2Oqs3kt2r5c8OJOMqrZyCxLUChH9E60I7ek4g
vh3+BibShatv7E1SjfeQFp+JjnRPhOkjGk1N/5eh760ozGlIOmljocO15dABRQyZ
i9vxDN/BHCPJG0Ul57LvKPu89rr7TYeVrC7DO5QejtO7oI9nM7t/8RR6tVL/IH+I
gU3zauvxPMmEtalb1rgIyFXBstTmraVLPPK3SWqLOfpC2OqKw4mlGZJDmnaKPARd
siLAqNcDjU7aGJgjFf6xdw9Yb/guAdZt8FZ9rUXSrWeo6J4/HridFb2i2vrmSihW
M9ZLa+zKosBj4eMIaFkrr8/zLzZxmvubCfUEIupWcxB5DKoRKrU0aLlEmEWYvc6d
/P1LNwd9QHt9moGx7WJU57+STcdmmHSlaaoTVwHhjNOAOBd9O0NrysHwjc5AaRpi
fVCqKejI1nn+ez8ihs9fHIezTPlV2duxWVZ6mwYk4Y/qDOiTPUbfBL+nnQcSBjRr
hvUQHSvN1iwQ0V20QpoVa687c3tbl/2v05uwwSuQKn90lPuK+r1EcwKea85ktZBz
GJa1gwfWLbyYH3ii32P8B6+7SSljlxfSzTBsGTBBqsJRuALTX8E0bEwhaHSiIIrK
FLxFPl5iCACoLruhmtkZz2b+RsuMueKTZ/x7zEMHG2v7sq1iCiQr1pTumS8tKjDJ
QH+2Qh+kvGdpXfXEbqDU5B1Ipnanz+p5ytvlsq2KhYG7m39d5o52/yJaaB9HdnoM
5kPWpUiZ+iGLSKoxAEAuKHkOeuNdX5RMqjJMo4/FsxBEQ/GS1I/lgmfGnAymOhjE
CpA2iVNJrjsAOyS0foywEWNW8cz8A/E4SUPcXhP2pHlJ3LRnhToSIRetBAyEQl0L
KSJvl8bmZG1LftqLs1y670C+/8ZYXfbylFOVLoWkwA8hspacPqwGGQseEKRlBmTa
pwnzmOAFPujDIfxgxtlr34CKpUK220q4b96UK/E5HIaD60UufsaNotoffCWIrdHh
H49/qQm9q54hqZdE7rMLVdQfkF3iq2YvYwRHRq0mY8W+2UOjuD8hFZYNwAY76zzW
ITOnubRL9gzsNrtYVinKetdYby7r0vueUILendqzC9eILgwc0y5XZ8qB/4eTzymi
yVFBR5bqK6Il3EEOl6zwTNWskkuP5+5wXaBiqAlGTlzqbXOpXKOwVt00MnkgftCn
IBX5yjBPTYxfDKWQDqFwuKDtRQpRBl7ZyxPjregvTFcczbZSATE0E0gCYC3bFalr
tRti5jJAkPPZmJLyLGfVVlOTmGXxQnEhJHOlP2s+h9l0HIvOgZffIPhzx2b21JCu
gF1MzPeQyB4jaSDR8rLPJZiY/Grvi0Aif034HX3ShHrKOnGn2jskpueKl2CG2E9Q
vzcojADrmQTCJ2GUXaqY4GybBQm7gD0Wcy2XSV3FOsTrup1Iv8WVuwRfPudbSX+a
eEHky+nSWGwT6RDHKsMs0y/E0aPDs2dkL1vxTXce1mTvwWZIUMsvRvgchhFmgxLr
9K7hYt0IaQUmCTmDvcNo+LvuPUiNRLoGKCcEnWUly6pmUuOwn797au9CUI8yhFwb
H11RObLsT1G9UvLbhhabG3/KqOaqVvVGSODQVrJLj1g1AaeOQ728/DfhXdYroYfo
prgq+abJaYbHC9Zu8qFLP6AgmFt4whg6Zq55XlUT09Xs+lKtagqXTR7Sc1PCgSKc
fexr+doIdedj3bkhVdUpksoV7Jte2XyssUjss+tLunv9cFRNna3yn8PewSNdahwQ
Xv6YWM6WUgZeozT7XTRj2m2KZrvG81dpdTUHp/xAqTblc0XxvSt+uMTsdNF5ByTg
nnueG4AYoSFeMB0IODGqCjAMg2w+jlCO62ROkPufvRqQzzjSi9Cy609IvzNzQLVo
I47YfGTq6EFvq31lQtQzNubIcwlsPNrldcXWp2tFN5rl8ElpWgBosHBGmUwL7jBE
9axfKLVetvU9d/KCckk1wCiEFYzIxueF8ll87FyQwrvYWxKTD5CoN2tPBPBUfBkA
5TFdKuJ12Qn7eKlbq902PjtcxkrDhdjbOLt5a88pFj+ZT9e98ASuT0C10is0wD2v
0HsUtXdRDCg5wB9rTjDWCU3S9n0lFtLV4H54T7uuU1dui2/7GhjZdsFA/IL6X0ra
yn0A4GaG0M/L7kuS+iUIO2jIlzFwHUsYrPPiRayRMCjaChAaNpp+1T1JaNASRWQf
gTQeGLPBXvuOXiB3GPVUVhXDNePpLdGqhW5UhbDvpP4b+rkckJmWtNJJNze0DjA3
MP7dMIxLqbhCj9h0SVOmCMHS187cORmJx4fZPW3iw6E5tn5CmE5D7uSV9RGRnK9l
eoeE3sAtzWER7wlMTSvwEv7h6bEKkGWK8O6zGysPzX34hnIbsJC9vYsHLasf7bvu
uYPL9oSjQboJzb2+FMNwrxZ62/OzYbrtZ2gfX3fcpMl6MjgL0JE8Od5EDxnAuaAl
ER6GoF627vPreCSAlyMiSc0rpWBSb6cfHHSAZBnkwureptkPjJr4rls0vaU5HRav
us6NVvw8jv9h4l7XJTmE+VqGH4Fj9uPB+Apv+QblguGk4WSf25XaZsyB+Fp2LR2U
WEf14kn3VoU5TPqaeDTScc04/au8JamTPbES9lNBKZIonfJhut6Pr96A6/XHOkkr
bwVmyxD2onQ3Ocx8EIblkVQA415lAY8k6kb2KqWrFxj/AB9ekOV3zVahyJesVOMK
jVKmvjxAbQsugu5YS9R9pR7Z1I6nBnDUXmc2l1HbrnIRZDF348Q7YJS/tzB9O3h6
Qa3yyHMX/X1314/U8l35oYVkN/qCEWCfBBwVdfmafb1MrI+SfmLRh1W2aDE0GxZE
uXmgHq74ius9559FEHpAc1lIeU1SLo0oMA6GlrXHL25pox+5TT7sw2Sj7LgkWbLt
2DEkdMHaGDpChlx24MxxCm9zZjzWtRxXmjFwWyouhMAPgbDMvgi5j4PdLn9DvAgP
4016zTTH7+2RazGyoeZ6etN9aJ+4bGyNtKnB/GDGPOc1asIO/IeYnzF8qfCXcCEs
QqmuOJJi5kzx4P/ye8kPavLay1/CyEaAglFsYsZ4rIjy5ttJbNhuDSM4zcnVecnD
9FE1odE7vxqdUVRTs6wxgUcoNtqVtJYcEyHwzP3TBnLEPf68SQu8AdUGZ/IzV+tK
3gBdMfVn6gmvq1r+tyZGftyHCY4/knID3ef59d8lhW+6eNcNTP4MkooYhX9Dw0Cy
Z0hl0oSQi2ONYcqxHgedVRn1Qb6n9VJITSpcOqNzADTft+0yD5gG2x86RhnbN+fy
IVOm690BcnEaI87AF2aNjM2wn/kwnGHYrw1lisRDKelIbWTewYN+kHe3ETJ4RNjA
RwV1RcS7C4QktV93t8bKtH2dlXKw23hOVpWA+cb7B4m0wf5+4hAgSdsNUrVyqCce
p84wl/px5bmFaijlEL3JLgaNhN+3scVaQgJCAD5KN84vB/73rfKK84qJa3JZFHxa
kgCeqIevspJJ59LHwUn87mLFIb5Ne92ud4zc+TWYr4+vvpMR1/HJYKxCOgALkyIO
YJ6ezjc+fP1d+9MuvlTaFvLbxuysnmOLY4xh57Y4UnTRUN3TYi2giv3AKqcT+7sJ
6EySS7eb8Ttvm0Fl0vm+ke0LNqeBgZDk5wxAivk8Z9vyjcg+eRS95/rPle4a6OKj
P32rf1q9hbLjVBy+/tGuelu9DMWw0T/j1bEb+AVI3ilmuTFrGGi2XVWm/CSDrTbp
vEE4mZ1SfrpjonbGHj/mtvl6RQMVkViC2Xy+uxcOrOA0ZJVip9Wys9PQHczYTrZ8
Dm8Nb7sl2zb8t7yNbTnIQAnGIZ6IsFGJOznyXJdP0oy+h7RTyVIfVMqOFFaa7sNR
tHJif8xB8H4H2GjyA//S8giApPIU060elGRvw6q62oNJiNI9GYexl0vO4cxtJkSc
47EunUxjF/fmJWa5LHNzSfyk9F4pnVqXoaSA29tOEYa7LOLgARCFDREyUQ+COO/Y
OgPZD+4q7h/tdxpR7ARH0Rq3VSLYx4Wq2DdDFezyfK34EvX1ksNNfq5ndMiWyqy1
vhulXwl7JY9o5efNkMcw+W+tpWCunxG73TqC3tyHRxWciOwmKFCt7ub9JnKaIIm9
EEI5qSQuCOoeLEon3LnSGa972xYJqCgPv20HcHY86Qi3QfNbiliD2Y9loGcEkHQG
wMRFY5vR7ESwx19AJVoOFhgq8sHwBMPgBo2jg0IxeDOvUwUmlRpxHGyL9pkAvmYH
5DLzrloZa01U/olCWEX3sqxr3ntrFLjHJEnujftSsD8ycNvx6cy/MwNrhNlD7QH0
XaXkcT17qEY42+i676DCAFyKgzR6Tvs5i928hMiVRKUKqPH74wwUMQXIfFxVRLgL
taKyDJMUSghvi5ZkSRp4nJK9QAWNcwKTy4Hst6T4F9ruqX1EWZTKPkvLmJY3yleB
B4A5YQZ2YyJXE9p4b1LTWw/9vhdVwNsi8oVXrMqSYBsEfMjASH8ad71frUB0LhT8
5BdlBDO9lPg57XaevI6XGAndIjPwI9AOZlAyKiaDApmk62zz7ViMzRhaN7y8oPfY
csFMmGWVUGftmFmIr5lcO9nS1stc33RtCpo8TLtWdkDXQuoXZR44DNsOCvW2tvdE
NusJWNhhAITZCCRo9++KmSjjYXISqEiMBmX5XmoBGHM28xWm9hbOjpxP7Jw8tN+i
OAmpQtl5lNMPBj+sVKE5O+ZLPST/V5Pgc04i4YUU8x9oBJavmd17gMoPr0teik1G
ShJ195WifqCv0qt1opFdye/AOuBAnrQgAJfcxvTrP9RJ0/aRc4xsPqD985xTb08d
ETf5kF42NvFFYaEXyw8/NV9fn6G8qS2KJMQ4WRTIu+gszA8IUPNv8dydmnYIY0Bo
/d8zmtl1K+yEfWeKOTmR7SXmQFAE9BeYJBcW3j27jPBJ5SkpfaFWJPt+jJPYtGLO
toS28ncrLpM+5yC6QE+4eAx4T64i79CVRZ/YL2XnAoS0ZxmPG/0v0CWXfIxtjzDf
a23n5Oo/QUuwUt9sP/k3gh7ScRzUGTw79wj/2M+afNtFcrPQAX0eyswzO2Hl6Rhr
cKAkc8nbH6o4cS2ayz1oWPwucDUOHlpLUguGCVx1xFmw8bC8pIn5WTxqqGkSrtAW
iQlYu2H8DGxfyqDGVifZnT4qK+LkTHWfqwIqi/p7Rc2fjOthio7VaUiKIss5VoDs
1Ck2pMw++2t1WsXubX+Cfq6NoV8cGbgVoRN+QB+pTlSK8thBEM1ICwWvZ8AOw7Rn
+fLQU3lJ6VzWd1fmzvqAN3yFu9APBZpuC6u32cZaqzMziA7L3jYQHIjh7+p5HGY1
hy1tyl61cl/kxmG5bRxM3PqtqDYCRPPXmdJwwGeHMs2iC6+eBUBKYTr83AYz29YI
lcMEKLsNnDBEU4/Sa3B6n0j651sAuv+YVt/Oil51i1WBCyJAqMTK50wXLwnbLw8s
PzaUqsKut5Hl7k3UcmxdgfOicnu7Ry4OYLeL4eaLVN9EDwUiPnousXPRyjrB3zyk
oi0guuvmTwzQEraq0SI1MELilJ1LCSYEi7Pw6VM6afdsSJiShDdNYZ3EcWAf0cwZ
S361NhYg4UaucB5QCbx7cFt6uhfutJfuqlDCsX9BGe5JN/IqNoq3SqfCs5g3azI5
Px7wXyaBmeJHefq8By7KNVC3oI9NlSMVcCENtIiE0KbWEqkywiqfTefNKnwitGpY
QjOPa4Bht7iTepJ+n3+5pyz1pGTacMUt7GI3VW7+lN0jo87sq6zFACcY9FCP1l8M
66vRRTxd1D32MngN6Q1b28ehuPebhnz4XC6S97IxcKyLuiO2/lqE9HN0XyzpTFW5
NGZnPblMuI3AktvhwfvSzQUkr3SYKqTAoMoBC7WmGGobsRDIA4FwDalcLld7Fb+1
H/+w0hQ9pG6CB3AzgaHZD9nXpCiOFWQCM1wtw6m/MH9k7jBOqxChnTW+UF46EwOz
QFb6wbZ4dkKW5FdNQuKa+VowaMZs581smAeLKobpxjQrlkMD3g3laCjuiTCy66SD
wcZXnvEzcBqTrbQCyGK1b1Avwz1l9RubL5m/hH4737Ec8SdKnfGjwby7hGQsa1uk
HHEGztDiIotJf0Pm0OgCo8KbAUjfvXE9fEL/Jv8Xng6TA1vtdgrgDf2RUWYo30yj
3H9SnrnBuQs1ZSWExRNg1ubZiuEyZceMkOX2USkQ/Ry0ElRlNNz3OjHqbjB6cYhN
3DAJJlpoWJPGZNh6ZgPIzi33fADKMkn1tHshglneXBDQVbunuYHOgmiQooOiZyCt
MymeZqzWKaJwISWqhndrO6o19ZqB5WzQjUG/9A5pkoIzgllzIrMjhqnEid0mwmYt
+3o6RijzElvAkReoDJ4iXanGc4Eo/umlW8jQuxh7u809PX+atuO62Tt1HseuZbjH
tWDjMGj7D2f2mzBks2Iq0Tx9oKkY6NzUL/m5E1m9jvSfEMsLczCBq07O1lG4ViJ6
Y0mturv+lBc/r3y6f4iTGhORYdYk4kdPAvewu4XwGjx1Vx4BgDa2YAu118glUPXG
eCTqVO6fjbvRuvsYDDxQxU1m0w3hmFjVMh6tVKjb0loCOrGrOJ2kFhf228Rceydi
Q0HTx84N8ESuuBk9lBHKF5XUc/VvoSnG4XsZQLH6xshcLGLeycDUey5u9gQodShr
+nTef/0kZHhJfMIGbD1z+HM8S3ay+NsjK386VnHsiNV3JY24D67cxWyrPbzsZ9hl
OLH3npn1MGhPWqQkxIXXj3lPFz6F/49DgDvjQEzpNqEtkFIf7QX/oa0rNiSbNSqw
XG/J7UVd7krG4B4A7GP+x37S5MeP+mN9b5pmP8TQt/ePKWs1OWHLe56f0Q8dcNJz
7XhRRh7+eY6x0EJCytNi0uMjX8qkHfqQKpzVFEt0RVr001k3NTZxRLuRmHsoQPlP
T1253Y0nvxTvFC92AqdsbVC6B2e6zpgu3zIKgI2seup1KCKL7KIh58+Uc4aDInoq
vy6Rd+mpQzCpjTyoXM5LTkKecXMWWjdHjejpIV9kSu2ZhQiXTbK/mcbZo3e5JVSr
8caxQo/ElCCeWMPg1uFZZUAdO6voMPRTIH6ePk61HgYOPdo5MEwmmBSA1oSVSrPN
u7/E51o+SiET47xKeZzNLkKlQaiSICIbO4ER6jRvF26BiaX/1TtJr/aaeSLb51bo
8LceVr/1EJWqSamBteoVjYfNmxQDF4IL1NNz9c8km5MXmB44OsqUOtdcqBOtajv6
5yJT+zhTIiT3G6Mve1fgpV5IlmVoTJJwCzcX+NIykBsq6y+zQM/+usjmDfYnH+Ya
NImBYVDIs6TXk3i82jce1qKaDAopd0Hrz08/E15zLh+m7ok/P4ul4fTL+ZjL/jgv
IQeAm/jOpVzbJCiNm0BhWWVvjq0mJoSJ87pOvbhPfrDlzQPz+Z+8h68drAoL9pd8
Q6WFlnLVLxdQFLJsG3cZ9cER4reQOoefpBDqYmg1dr+HfFnSWSnoQl4VlEYRNpMY
+jaSEQUV0wlDpKCa+jQxdnPT3LIVoUsWwW0Ly0QDqkOVU1RzTqoEwFZUImp3G85i
aBPCZDEHJsOIyoe9Qr8M1Q594PgdQv8AswikIa7iS/bTuR47v/IkfSNxdegrXk9W
6iyxl5S/Vh3ifH1eKcyfv/Nk9FcTMU6apNGmhN//fh5hLH8ePATDyMI4UT4lgW6P
egvAqNSXisjbqoJg3qeLVCaxuH2L1FlmBND1krqxttc+NXOq6LD+tu6pDhb4dntH
NwEK+uzPqMf8AX1w+FTVrQZiLuOks7oigG1pDCkWEskzR/Xm0FmVAoMVqEsdotOX
+Ckm/n+UJvwZTJAnAmSIB6IlECHwaVOos4os1i23HyO+fbeLkJh/GnSXYrcMpDNf
7o2bVTCGoc0AGDOs2loKTlXKhPu0HoaLDMnswa44jrxQg+ovtngOsYR/wJnmTx4b
LUSw0Wow5AgssImTMfRtQIHkI5gN0J8FWVuNXCdaQMTkB+8ctYawTtPWCSGsaK2p
8RolBkQqASv8dfe26Q58b0baJat6AlJI582IVCgH8SLr4c90xnZAI04spnxNSgK5
RlsFCVbQsqCxQrELeLG/6wjObVLsQexrnEiYtfDnTV97HZf+fJ68Rio+Cv21s3P1
qHNBs0j5tZjOZXzgiW8hu/C2gNAgzIfaID4cM13bbRKUk1J3ZhYGnXutgDDxVdrj
MPENkTV+lGFbz2d2mQXls5grYMB7nBsW7fq59pV3Jfr5P93yzabXF9g11fI3n6S2
ATrc0JN5tusQldCu+XUVx4JSfPVi880P+1WyZDP4hvV1l0WtAIgSiM8HElbRWWBq
xo3BJ8AnT/q0xnxPTRAeKuAZ/5+jTydl1sXvQKACOM1aQC0IP5VQ7u8QnI9nLHH1
g0zWJEpwEaeIa/fTQM/qLCA/3i552/h7Z/kum6FFekqgY9iUFrThZkf0Cfz9f9zK
XIbVGPqpDsGBWZ1KpB1Z8/1vFKl0MsxTerkQ/qJUjfnmX3Atq4bvIJm0TSK2OKSJ
+WS2DG/nN5E3WgEaUIx7iCZd2xRBXyc0bftyDDKwrYKinVU71yyfLG+4i7MEw+5A
N07TBDlSJJy+6Ib9f0AixllyVgTWlADWzVsC23O+FooVnCk1TqpqgtbHzjuaI0eY
JPFdNGmTmrUnJji6/uZlxLIPxoDwJAWmH3joXU8mxufJp92yX1eN0oVphu6Q6otR
fFc8Dol6ofZafAed58r1AQXgYL1+4SkDkQb72xgJuxLfZN80N9E/Q9ycamkjymm1
09L3kaWzhvWtJ2w4qCQKGWaDwxIegAp7E6Qj6nBGeVIgknxduX5QmC+kO3uYMe70
rjHEwm9iVOUsjobnC3KHfMV3CrMq8u0RbkZ1gjd1FSOgdjk76x7lYs4wkyXt4Hzg
mYZ2U8B+VyY2oFusgVTuac42CpHjO6diTDREnlHe0RA6qE0+da9BiAUvZNa9yy3E
bSt0hqinRy/I9c6/uOzUrGIX60R73BPtkZhkcn51xaleoRmUWRPr92t7scDPr9mu
KONGcsNCeXWpUMJ8stRmyDDXL6pdmcgDnXg7RDtcLH3poqqF4/4ceQ/iqv1oew1e
5ST5xuw2kf53Mrs7xA6zIAGdsQf2qDKjG+nJl2cXZ0DttCeS5VxuxaPXF+zL6Jvw
wx7HCVvLqEAjgmnzd/ckr6SPzWAkOivzqbBYOWIxva/QH7vIupBF2zI3Gwg5VyvS
rbgNhIuy9l6OR1Sr3y2Ny2zwJtVBa019cxCwXDe/rWu/yifhAQ2gZDPzxv/JfAcY
yNB6GGg+3yorKFK/WjtOamFulx+/F8evNYDiZNGIS/UI2grvT5mjxjiWUJzaiwkO
46Vb+9o/ScFkDx/597gpYBQCABqdWi1koGptWbaV2s0XALwhVFrGZN4roQlUAmek
UUV8biGyFu5yjJHfz+yfisLH3Njz9hKLbOlmS4v7I3L5D8vQhmXWCzMm/wFVeEFy
afygvUudvHXXyr6/JUHiuGzXu7v0oz1X+lgxF3E/+iqaceSOBcbx3hEd2q8/O9iZ
t1D3vU3j6JH2yjo/Vx5EvPKIszyiZAiwci9FC+jZoXkEABrxyi8WV0c1N3P7FFGM
/TdL2xblPsBRkCcnduOl15IRbLKQIw4cQxHEKkXBwMxmem0eEQ+9J1Zyh5Jp5K0d
grmUPUu6WCEQgPxSKkblbNDfeJFMXvx88woJHhwtxcXQMnHHTBltxxG8IXGNwteu
4+a3xWCe1ZmwdjuCv9AvUOV2aVivWqhRi6ikvVvpJ9RnNEtZmHvXVWEhu5Kc76G9
DknxU1kXEWrTzQxm3Z5LF7IbusKfvz2wY8xI2qUiRl3dI9sjPZ1GMRJYEZP5r9yQ
s2lTlE2AB3aaa3xsi8QJb7pK/4FU52+85v0uJ8qPtESjuWVLuMofFsomLCDhZkbX
RIu3NHvRfoqlvqtGhpk5SyA777CeJbYz3hfBQTlkzq7nZcHUzsIzvC2+RdXrhP/S
czzUV6dmGugWE1oZRMOiIqVhLP9eUvFc/adp8MjfDXZAQF063hiEJnHpQrqZtqDI
5Y8+AoWW3EzHFBq8xPW/7NfBWZ0bJRFXFDmmlcYNAOZAjBlOGZTg/0E+Ff73F/PE
JRkwmApyiXw8UfGNpx8CL9Ypr4FlK1PvHivTVPsPb/JZCxFM2UqMU31kl+BlmFAs
jaa9dJlgDd8uePfHsv7Sv4xL5t53IxP+mWYyIcjc4OUJkZRDDGg9nFuZlGEmp6Ya
J7gs4lblLJD131JKrnQSPgBfPofZiPkUkmVbL+WivkntauhbOARCSUyUmDSbFsDG
1e4J1/m7DKAhvokwKZe2B/dvQ7GduyhhcrJDiqlraKCLRFF9Ay320Ptc19EfrCYZ
H7lxqGYBUgfHRpLcP6ewjkao5UPrG9O0RJze9IMrojEwI+rUxR3XBCAnCQPc1dDo
0cR4gXL0Oryufb0HIee0fWEWAOfpjDOuvknh4UrkSSWxjGhGT6VQLcqxN8bhQPIX
N+UUDWy+4U0/ziqMMaTlMTgHxvtRaiLGdRkZ7Y/CYNBa2aNxN4bRHP9SbRcF3NtQ
mC1E1w6jgCwm/arP9YCnsNdDCqTQTzrwLy4710rCkIValzwQUgzcY0U7ZCVjCVcW
BY6GrnjLs5l6We5KOMLDylXnp0/j6HA+PnURkSw9EpZSsVWyRD+0hBqoXXgQ2vPK
8gEhMla0JNHdj6g33zRf2UtQZQRssXJ1X7IPi7r68dv2IA/ymdviAvy0CXvqhkhl
zWbtJ33IsjdWRXkNvbBFmREFYPcGujX9WQJrVvZdvnoSqBUHpWLe5kBWpMNP57VV
Qa7IK78AZPAtNMITSRuVOq8pywulJxEXU+cEvxLrPD+kp5AoR26mz8Gl6Qj4+Aml
qx0PGD53/Bw6xzSaUW6HS2bscNDLaQ7xYgLqQOKELyL09xrH9vupCn2nChW0QA3y
P5GLu58bLKcPgG+hoYLMFeo2pEx6xSUeB29ZZVoTBmJjC/1oD2XQpel2PNXNHZFu
UcWtms0SAhDomDepqa3Enrzqo9B9V+cidOfDcq5KWJkba2oGnhhrmYvp8V7sRkfj
9fAppk6k64eKJstlRs5MryezOjxQwLHWt8GFX+29EFWF4z73K1c82K/LQsjXvmoY
ClGDk/YL9PXarSugYHCemjOP7uITT9VA8MJP2jAi9H2k43MLCtt5ILtpCnAcUxwy
guGzXb5hJNX3f9ebCy+Bcl1MzRWSm1rCET6NaSVlwzbqda5Par1ESMXQulKpwqq6
dxTrGutdlEqtKi6vorxVT+R47RSqaKiVihPT0etWXvsYBOZk/MCF4t8RQXeMVMUh
6az8CjitHBEzm6VuqxsZ5m+X2wzLtiZvzd1epjbM2udVZIcdLt8Q80pwa8I+Uylb
NKF1D4XPPkeeuj9PUMN+qlRYDguIlX3Qv5By+3zLG3QE2sYB6to9O7rbz9IsxPWK
BixNmm2pVVWs1EAxH8c7s/Xzlh43Uo1xMv90+d0pS1q5U2MZuu5AZO6pMsVaZn8u
38GB9T2GsOyOaJ8IunwFOGC/C80aKQpPgYL1OM0eP5c2AWohG80ocy3sGw9gkwN3
xAR8cFaTNZnRmx5QYahuN64wZcPYpWVO7d/Tgzqx118MMRNZeyHvMgo3JPBkM6Wb
nLccyzR0npOud8NFIF6cWNDnb3r/QJUg+BV2jAdO8DCwROgkfN2GznjUw3uQWRca
Kll91VdxhapldvOXNxob3EEz6UcYaVUNNkecNrOurwDjNNrW5m0sJS/VhtpqxTMN
0vE8nRZsGBifgzjdy7XKHihljlviyFoiG3WUWjToU6UF80AHmUQ0Hbc+QYYi0qd2
ioX94R9JkrTut40VQ7M5oIbwAOwbV/4bofFrNESthk8Pny6qENgPpDZSHK1zt3Cs
UAIES0KMJ4EneqVMbnPe61yuoUiEEU7/6leOtjtn5LzqAapGkkKzUkxUI1CdOkkI
Iqwv887ixXQZ1xfm1kUl2PYHlQ7EtmnZCuN1vTkuKWxSmenVHEZgA46O7PaJ5FOy
SBB4Mhgts3kIjufacOLeu3wSVt6Du4EGGi6tYS7QCwovB2PmJqNUNXqCLjiSVsSI
KK2QYt+4b1VrfB/Rr5cR1H87KihsIksIrd8+uJfkW2ZZn3OJlFjly6le96/S1mrL
2NWdZDXnLArr5jNho3Mmt0kiFpUgcYrWUgtp2khz2rwz1YvLUpiGsJawbcXrzA7C
zWktX50e9ttWyliHTri0xuKX9QsuUIj5FWRpR7sn8y7KFy91Ex43+81rnTypgzWu
KH8g26QpbI0wxnxlapkhpu31wdMkEVmuNCgIn43NLjT010QUUmJXLs+YoSUagiX/
OupUJ10iw0nQKUQZslOz37EevcoVjdo4Iqk2Ugd2eCwvkAySYSTgZcr4DpAXDDpJ
lQLzU1us0hmPKusDy5BQS7aH8ksmxsmmwbj2HMpOQgHjt24mPNwE1QyksnPV+wzY
tp6IZrlk5OKU/5WtldpwUr5jZGgCsLpsVyBFQwd6LYS6zMI8Jh0HIaaRMcKjTpWo
Xh5VTh5+zkWn37vHn5wmK877m+JKb+Cuo0qo3yougYJjJjs9xdY+a9hlUj2CcuB3
ugnHrVY+S/V5dF4foPemCG3nVEpOOqqHWZ3W1ZJqK7n+jNYeiVJSO61ayQL428lm
zXMsIMqZ8SpyIsOaZC+BOKSy7eFh9ZXVtnJBsm4u+cUhHo7rN5I8TyFj6op/rlbV
F7VcWBuFYqIpyIsbjp0L0MDIq2YZZxB7a9ee5JOK6EDx5Oh4sGLn1/ekloGKVhW/
jr9mVQ/vPFy0CAn+lXI/HpZ0OURDEEvypNJ+SnJhWfJ6pXtlrTiadkDlm0XemPwO
S/UAjYS35v7MMXqrc+eYRQhK2BHm3HjUpLa9Z8ofrEEMjzRpe2KCs2K0L2BT7YUw
EyaN6Pfz+ypwliLQJ3KMmCYPETf8bsVKl/6i8lcoJB1u7jt/znqoB/XqjTQClAx9
lJYhL57mrcZwe9dguGRefK6SMMGbSO/rLtkgP0P6G2PwgBovsV6IB5/KJtwwW7Ed
0OlPhIdve+ckDXm/ODP5mlmUvT28oKYd8EavmfoGdi7yeOHQEeuRnqzPhKLZbqB5
k7RNdhsVZrHMoPtDhecywF8dYCwVOFD4LRzFbmTuyVsnJVRvviWwfeZ5Zwh2LtDn
iE44EMNmwbLtnoNngMFswCPZhE+xudW7ME4IKHcVhMB8rHTUtBo61rdnT0XS/Vr0
CtXoVNcTgmWMZdpYzQYnAku7dN9EUoIovv1znjUB7eK0kq8n8p6k+KlSR/SkNkMK
e5VwIkBUZhIBtRarv+fXji5XW+A7L4fYvUMtqMpuFIlnnG95DBICn/2BNdQBdZFD
bbuHw3qFmrXLmtaT0N26FcbR8zj+WsMS5rjCvbRj5Z5UqIDF9LUZN/yhGk2+Lx7+
F7SWZ5JozLc/GgvuKuh29PwdRC3BSe/0ajAX9vx74zanqJQkkOEwhuVKX8eStyTQ
n5loikTeBMzmrGkZHTcFGHT+sKLLkdcukIiIWPcunwdFHsEQ1hURAj+jusHkvARK
zavDJ5sAIZZB/aBjZPU3OQ2RLJJf4wH8Bn5q/d9exevsdEFJmdz780mgPYl2JAFX
PPmmHiQOInfPFlCjdBv3lR2XryW0/qC6sghWeM0St5dOIO7LJ1deGBQQaHFcqGSS
H6U65BnQIluIQuWXlWJSUithcBiLMfcmFxXoq8utlbGVbCBrh+3+aHS372Oo3M38
ccNLLozBlb5SI3om/JCEWgib7mMqNHnypUZznTkwsF7pVgnzGmZLkpVJ8wz53l6g
sp2jYFDecI/41LnOcDmWJzyNm/X/4nH8r4n0Gb/poV0mRBuPhM86WvpQtc6oOyGj
7uv2O/xUipCkvjiKfMkyln/FdHCu2uktiSCtxBpNG7IIvAd+suHPrm4YewNo4NpK
R81RLBnD7McVtJ35aJQgyE77eadV15XUtH2iZY3HafHrKSP//gQTo0zpTQAOzbam
ELhge020J0IwmvK9VGhcWx6A6vPzbGJPw+GaAmN+kztKe+vN+fxHZqCFHHjzGn0P
xAlNE8gPrF32GqhDSJSrjgF3rcCrWAQ0JPcpNBkqxIlGAcZRicm9DUuiUZB38VfB
nsZ3oWZbXsw0HPn2LJ99AxMd+L2m8GTfCRMuAZchcktSUqhNhTpFg0HACfDD+cYp
tZf2Z1QtsiDSfPw7+c1Fs3PwH6rmv2xjYY8XObqPZMEXFkcHHRxORvdPFYOe1qsW
0fex//F2Znh4L+r5TFhsKMZ4dse0ld5tRjg9UIw17iUBaKSB01tJmM6bXc3kaApM
AF/OC1ZTDSyt/BSFzB4kny98gyoQ1tI4nhz5B6cxIAFnglgwgpfYviHByMkNgy1c
PIe9+fm9JAaCw7RFWCyZZWakMym3OwVYZTpj5i96kQo64XuKGReFB3KqpNUJE3Zx
Tc0T0eC+vbXiZiJeSSjgUMopLniOwHAFuN6bw7RsRUz9uQR7AXYZ0NQp5Y2XuzJM
VjwzTOcvc+f0psCpTPRsN4PeQWfBnEXH9n0BYD7bxEOFTguUQoYbpeGQJOCAUDQd
GRCTsGZGMRyOvOsQK5IVa68Eh61sYbZ7o2TSMd749uLf5Xigc0DIxJL14AXXW2l1
ye9A7z5NlBzi6Gsk+nO2ZvYE0vLIE1gx4QHcjthRguJKwzMk8Rx1qm3Nf7E+b+i5
upkiV5UicQKbyfrnitTp2FeO9fVRVkqWJskL2F46VXpr3TRmMfkXjVF1nubJa6FE
8rD+FoBgwG35xf7LNwA2VMQyb+aF0/gub9GwG+2m6vvSL8UlqHUh3M0NjSz88+rZ
+XzuhSCWD+zjDeIwXFva0HZ+o6f8Sd2pGg/uvvK6t1iXWtDsMzox2kZpVot8D9A3
7WFlrpPUoeCNwcCbbnlipUWmgfqsXNkcc6lbQxrFiEUxCxR2LJ/0GPcnmTfIqe7j
E8822sjzy8pWuD9h+KhNA6hKvhVjamKHqTBBiCQVBYpO67TnddSh4GhVmaUf8IeS
PButkzBbQsJWjSbrSnBHNZ9LRdz7oPly0+hEr9g8JaEVD0pbWh5hTa8AH7ZpAzzX
z/UPbgL+fFve6iLBsJni01B6oDxF3mKja4JyyyiIZ7ZDdRo9LRy/T+7VLQfyqP13
zurVfSPLnKEwe0lWYkNQaAujz2HqIvNKWJosClj4mltkF1zfqh3rpW2gxnZmVZz+
mh64DZSS+wX7pjY343k6F/qI1ipk+mcGcXMt6ckZ54RP9oenus/kYfpGvLVkRKqF
9/y32SvyrKdkJN6lL+M6uIlsr+YQ0hm31i92RcoaxA+4nCohq9+g0Dc0ON2N3Bil
2HeTaLu5ifLs0RdH9d2H0nxGYraBfNxtGg4LFpNJqdy2KYKKuCIwmGE3c1gyQVQP
UxbyeOEpAYntA4XeBftYZXk/TFYl7LZxEthDEnE2LvgToQl7Hth9asAgvYvZWDHP
7QHVolmauTu/B2Lh8YLTvs8HIhiJZ8No7JIPDgwMbEvuvjiuazcL7NWLCe1DYvxu
Bhz4keOK5zo7aTpw2OmaRCZ23776+dO3GEOvkbaqqQx6RQFgiPWqENVssDdqFmT9
yjZeWMqzyun2z7LQOIps8DPNS/OX+6kqEKk0mh4s/RwYJ7iQFmGxIvR9tFa/zkE2
e0QrJhqib8m+sUftBsYQy3Qg6M1bw7TcOkjpZTufUipPMOTp3/HtLQuLOU58ZKI6
q3kzXsld7pXqv/RaKwVB3Zr8skQlrxcxh/jJGwREP7DXejXsLVBX4d+9Uy9XaP6Y
NBAvQYOb9c33vHC/K4jBMayk64/sbhzSXK3bw6+DEWfdaWHwwXIZnHzfMYnQS5IA
HUO1bNWz7T+6kQKJD4UoJjkG6nOFwjOdxeCr9TRxHQtRzTwqpFDXDJpRIJtxSgf9
F1fnk5F1HCVJp7ZfYoH0osBNamKZ0On3B+zsIvEISkrER7Pij+xncZgSlwf/95tw
HMJgxm7zW65xGM4jppAA4patYxot4S29Vb2QdFWbRubGz+p1PE2EAcYpdsmB6/I9
TBWdbYtEuAq6Mpl8VPk6IM3HY9gJtzITRKTsxBR7pleXAMAhy4/xaF7AyqCQtaUH
rYMhTlPUklt4pzLRsW9/dLXr9NurENdTCXrUUj8DxWf0o0OrbRMJK0mfM8NfKCMV
nsZwx/ROOOQ2RQ0sSlHSS2u6NutJFJ/E8Ap6mGyiOeheT8WzZX3Jx9ynJcJ5xXkD
unSF6lTDHX555ceIODVzX1HiYZCKDrme2E3LgBcAz5O1gwUPVeQHt1YcRXKuIrUZ
ZDgcYHtjGoSs8T13gcPPr2Ju4yTI1a6wrCjpdCNGkI8zY69eHINGkTM5gZVX4sgb
2GNQNW6yrJkJIz1MvbEegZPztRD0WMCfzmG3jfVAwwHJCGszOYg8yiI3VgsqwNdC
crs8mEBi+1z2Oi+gKN7OzFhIOSnD0TNcSuqq3l9aQWwhcH6fgGHsD/Pp6Qo0KiVT
aVc71C2Jkdn4w93LyrI1NGl09CT6eXe4qY1fjmbXuZe0erfq2wFsOsUBP4HFvVxb
DV5UlDj3O9QzP6LOLJnSXS2MRuP2BzMoYD/WMidIlwlBE6NrcBoHkH9C3r8c1cxQ
hG6avGqJnw1z+jtUR/O/HRxUBALJjLpq0+A0w7Rs4MJ5XBgRsK9rdS0MKU5F7PmH
y8lWeVHMyg8DhSsj1Tuuhchpp244ucyTZhvgnyXtEIDZ04bac3DbHv9TMVzAGN7w
QaFSS8Pr7hKqIV8PxDUImHbryAwOInNSiWcKGLKtYPPRAvBD4ocbOsqVrXqRkTjU
SgBN+432gb7zCxfWFLXFkJXALy0O7wUvwVCKo+m4B55HEPNwvNTpP7PN+Y8NfrDu
A5NAcSTu7QqJwwJD77TUTNFNXVS5oLZqfU69sb7faSGli78pOqbHxY8TbwNIdfbJ
xsDmTgR3rQ9sM2kjPw4qO86MjY764A0AG8/2cbjI1/7o5Kyzq0p9TTdkG0Y981ZD
IDzg68h7ghlxyPkpTdrfoGgamQ8LyujcQNjzhM52kOP9WY9ZOKwT3ctWn488Y5DD
wXupzljBneRwJ1L6xcFBwn5baaS4IzvvoL+c18uHZpPO9M6LwYNSryF9kODs10nf
LrAo278kU8BVT+M9IgDBO9OtsOW+dCDYZiJk2q1OPfSHCE84z0sgUULEf9GdmWpj
T56sch9O9pDhKFOsip4SoNgbrufTcw7wGKH8mnMG+KfDrVzFuu8TCIP41ntHjG4Q
wSOF+IXl5SSGB43ugXP5M3vLouFv5AfjsOalWjPip3S4m8HtkqeYE9BEs8RVgIAU
hZQYxJJH5XfIhNQkPcHuuwwTa/TRGFl2QSGEr9nKg8GtVzPBw/xaIQgZHE5X8OsG
MBXlxIYTE/KT0/Ciep0DqUNFgfG62nk0OYyf8398nzg+SoogotwG/F90Q2yh4hbd
t5pW2JUWgx4gzg89tR5FygaAKO3c/IY5Qq6b6ZfCIdW9VHcsnp5uowGszs9BrXpm
aJJVwZ1Fkunh6q2YYYqF2+gYNjJ0SaH2OuMuz3ZyLP4AkD0cJ/oB41GH/DUwf+nL
f8CJsbJeIWH6wlAfgGnv1j5Omk4OvpBU/ASg+Em/x9PyIGqZmw4jqSkEtIbh4Htd
9yb8GkaTxIcD7mJLchVBTfWnBg5f5RcS6Zo5Mf+vNZ5UZoOvoqOiVMinNDiahUm2
swTOjEbv1Q42IrhEZ+I0z9V18Eq39ka1xOaa3tAQPeIjjJ0OZ5vKU96lcX4qfZ69
z41i5rVGVvXEoZKZhouWHlIfJjK3v2RN5JQb35Fs8BRGvOQzbIKQkksf9nj2oM62
zB5cIFhZrNvvOLbT9qOs+IPtCtUPf1JOkXxCywGhmUOhHhwU8+ctd2n90KcXC/c6
7IAQdqNm6uHhWmhmTb0xWPI78RmqjciH+wfMDU1Ddf/CfJREYGHZMpAWyWAiU2Bd
TF3H50WA/1b+M5SL7k9ebdRdSsvFTlqnSLQIwIkU4ajHBOBxTHIPVeBmI74w0g1o
EN0IRaPnxgvLKa5ffOf8635kcgT0mfNnyitHtbginguIER29TZDLBEQyyjJ1DxsS
+vtq0LC8RyAUHlQFn0mxiQfj3EWfoDvQWgVTJI5K8K1957PuVUKOxK/mJrwIMF+H
h4MRTRFoWkZsIeYu3e3XIHhJ+9MIV+nsttBAnQ54ei2Q0a69j5FFnIqUObsu+Bhv
CG6hORLZBNhbk62hEhuGFi1MmkGzms5C+yMesYc8bUheoIZMKno34cwYuMhDf3nU
ASOoMsxiau7m7sTnbI5Ae7U3PLyCExDnYLrHV/cbKFnQNnChqmleNfTo5UNXF1B5
pGv6ykaXpwJngzOxXk0J46DJJeugSX9jLwd2LWjngxnyTGAcUxlPGQ8hSmPsApeN
cAoM9v/fvhEdGc7ifAXANVOdU1icpilQUED6sszu9GbDln6BmZG/sW3d4PZ0CSG2
qL0R/mPyo4y5zr2Jmaj1TCIqb7aIWBBcPBxE79QmMFVoUm3hLWG5+Wni6B8c00H1
RVKIBDvnqnkKa4j31k0VfmzvArgMwpRITfb+AVFVMtUUXWtDImtjSAXvxxvxuIoH
8SRZEpzvWVYXf/or1LHs4SVtgkshqbfwX7rTDYbxoNMqXV4xNCDwVLMKAVujxbeK
8IQeE6ehH7mgV8En7M97QCHg7eA92bhwwUhhTPwigSK/lg0WbQ0zkwCzyrWHonth
figrFNgu6/zGuvU3xuf6MUOMfLR0NkItp1/iXnK6jGEVRpjYV/NEXh6nhhW/EXuB
cLNQ/afFhRH7Geowp3zVgR+8KQwm2t2kx2ylXifreD3lfxLrL2fVyPddUUshN17K
DWqhf2ULwQzfKFU6wCyy4Mqxe9jdI2jF9SUDZ3UBnD2QbCTjx0NF3yQxPpwyCl+G
s9PjbtY7LEPlv3Jfi/I8VOhF/3ipdthzi/QXUUiYC/oacd7sX3/qSqfl5A6KWuSm
JYiDdW3r+t6AmfEbZmgOV+vCiYgDOw/Y0JrPh1F0pn9bRrjwpSH/FCoPjjS+iMUC
NFe/kHeGQSsYtj9x2Uf5WCtVMDbphzqwyG2XzKMgWNy5+oxTLuyUbYKIcq76ikWl
ECnLh5j5AJuqTxRDsMsIX6Hn1OaYKTv2syLgaD2XNPZkWrpvHTonu8lHcSaheh4M
RUltMoRp+ZO/NudzgShqZ53E7/SysnfqBsqwa5jrHC1r4QaTcMoTe3MQrXrl4rYp
o2xoJidU6p66Hem2fgbS7xjN2CURbznjiOvtmg10pR0ZagHS22/7womR4Bfz2OzU
GIS5kKbL9WcbNjgf9OadK2XL+f9Wcb0vra/4A9mLVgzERXWKI20L5UaVs1ZkdSal
DScjByh7IfTPMEYc8Y0NPMq9DqnHv5vt91Qszc71kdGkH80QgbOQFPQ5VXiTmFoH
A4INIe00/x4dsOVJOpDBNX3jcsOP+HzjQTA1WKgS0XW5ssso2140agPLss/WJIc6
yYXnq16xFreYsLhkDX+aG9lDED6VhINnTarzUTns7fDGk649fE1g6Mf5yFozxtET
an25jYcF2TmEIcHq9Egp3deuS4aJHyZNzLpzbRIxQ7Q6Xi/KOMMgdUOYYWEDMgLH
7e0vPAKXG4AhtEokEOzweihUTFQ6tyd7QETqkI/BszUUz5nd3779jQMqa0JHVPTw
c2WyDnvNvOn/o68T5jmWES7friGzBFih9FD8Er1oS/zI+qhn664F/fpYr11kFZBc
`protect END_PROTECTED