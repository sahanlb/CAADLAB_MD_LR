-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SxkXxb3rQJi7/x4UCQ6sQ+ZCsLiSUErFAYQ3Fllx6IpHgmT6awN6cw8HabOs9qhGNW9INBGxFQd/
yOFhSYoLTDsSpQqrGzDrY0jXCuhFSO/MGLdfRNJDSTFYzGCsseSkptGk46r/EB406KRnjX19wGKb
qrolN4vjovtVUujptuQjbSRG9vSQI3orGtqSGfk69T0FDwlaY9DOzLqu1sbVjlexI97/qUtTwsHy
A23G+EU0FOWYrXKdbCAh5XtQ4tPp74t4RomBwsu3ROvXl5EYWgnEhcZzm/rvPRD+y0VQc68156Eh
RYDOPd91yU2dsPn6QrWDpV3awbTO+2EmrIBSQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7952)
`protect data_block
P+8mOOGmA/P3lCljbNzHnPGTEMJ69fh3nloz/HOSTaHe4nXNWpYRvPpKPEmnxm5EKYiLIRKGLXOy
Fu15xux2zM1GTy/ATt+ywEgRqdQ7HJroLpUK+s+s1N7eUY2vLgcMBdMJZ5BR/2ZcV7X5H13rMhKU
/9y56+UeJkbJC3cm+ccglkxTM12S4Un7ACoyyciqJz+5Cys4WzrN9KJsmgqD0w3UrA9vgLPSlpkr
77OsPbI2IdejoV5+VmqnL46TbdLF8c+D7YcPKkWj+S85FYUvJQXoODuUbN3Vd22JdIeQfueyXgXj
1YIzF08qFDcubhSH/SLH43cEcvu54I1FVrAXOTTyeIpcICfTiOb0UI/HFYekCCmDWjxMNTepaQek
uysh3iYk+p7B+vl/ByughgRPABxoguUw4kv1G/KuZjUTObW9D/Cn/o48DWFQKikzCTN6/O1bnoeU
GB/jexlqaMn0Q3QYtUw74xpizdkDOo7IwhZGBLZGH9UFf0V++oV3e0isDBZ7frP1sO0cGb6bHDq7
y/Bkh3CJp7tJwA2fR7GHfUSEJOiMnwlU68zcGcYMAmb+LnqWhOBNzpTPspplsEoF6+sz7j9zKuWo
/OnaHwwX4CUriyvnR6O8XfJsTI8Xn9uEuYjItkrcIJ5aUZwCLtXxb0RWd8HNhbCZl0ZMglaPzyZe
87/mCzthfJlt/CCdoufhV1Gz6aVBB7G33gZZfOoyW/HOzVVLcxVFvlO34byLIqfr6PQIIowID/tX
ReHtBL0A1yQeMKsOB6c4DZ8I1JBXWwW0k5TTpFGBw4vcHBsgM1jylbRSKEY/hJLNlRpVJ6HwKtSU
6yzo7CE1iiMFQK3PruVC0SGiXk1YYqjAyfLJa4+aVx5jl7mNFL++WeofFKBazq9tnQ7a6ls1tOa9
BoTShXsx97Bo04ZNyQTzvlh+qRCt1p+Jwl4FckZTkNAgwmfpuH02UApf3SjiPyYPFYt/zlyihpmk
j/yQzBiI67hOAzUUS8TJjypZ7zVrbt6a+JHQbAyCwVDxqoA+66+hG4llY6weNEbpJAHrch+FZqkR
IyDEUdF/pP6K9nEGS1CsCfFpbdLq/kO/Ku+oZnL0BrHpW8Kg5afSMyPRK1X0WT33Yw7wxthOmTA/
Ok5dDEFnpslEcO7r16yGjuQ7Txw4tI05tD9UMKIkOSlRlme3f0gW3xY237fgj/v+sDuOaW8FbJyc
jquYmxA4dkriY6XX+snKqjB571gdtwwADRmVuFbbxtoH/dzTYnmEYmO5A+tFwO8a4qxie8dNSIhc
pgxoKYfhx4g/bafIBN8y9VX7fuB8o1pHII/IM8NnU7usVqhCMPsst8aLCFmg7DGlnEiDp3CtcyMd
pLa/rT6KUYVUqANb53kNfMaYvRc7cLfW5PUsaBWSoHSiqnaENTMNK+hJn0CFzRIb9glYvC6aIO7B
jeQl0KprthfM6jPcbx2q74rQP9tc3YmMHMpcZ+VKUgb9QP9SCOfrIm2RD9Rex9aCYJ5yq4grQ9pk
vWuKDf7Rz0davCd0iJMKABYwSjWqNokXIq3fRkDMezVrwKXzHx9S3rQd0nyI0gmDgJFhnSDfPtpx
o6Z/Wuhbs/3O7T3ZWfsFL6smG4zRgF5zI0gtMPqzQE97zW+1Qi4VyaiBr+DElKlPJwrHNT//KiAj
ueZj9D4T2axUywVU7wohRxCPgWcGcTSgqRGA/lKyNh3i7uZJFXZZYLQ6LbgJGTtzee5H2WX01k8V
ZQTUi605zk7TMuBNx2xlr6Tc4o+VF622GEXX3cFQRXCquK71Cu1BEEJIqaCfoZ/IPcbXM3hmfYmU
4XVWnE1WX3zXh6a8b6uA/MQ7sCmY0pF3C0rVvFGbcxZxqM0YSjxqIVFN9PGTjiLClwbPuRr2qBKb
KklN2OcUW7pnV8dsY2oyqE7uBENw9tAVRzpis+zcHj2sNjCTMlBZ/0ec0XHH3MPbZ7Bsw4jxmbLS
QIrjpckJdT1flJyvfh4uE2OFreVIJCRf2m6wxvmwIQjsCmbfSXycKNvBMxQdTGTfnvYNL/p+myLt
LwixazQLhSZYsYVxzd18WEkc9zgfGVPUFADv9IYhvmJyYx2PQdre0vL6pmJekI8CKVrUnvqMw+0z
Z63nq1E9HLKQDl3dGLlWyUy5xBwI0a4a/42PznobQqNs7Qqq+VHh9Gj2SGfjffthjP7rVcFi3QiS
JsUOXR/Nocj5JO+bxsUeh/IV8Xk7WnNPUWg26hNmd/zSY1NLtch9p0yxjQTZxmHeFQposws8fl27
tpjbBgbmEu7Qcm9TOTmnShIeB9tCPqzqP3sb8CbnkZl3h1tmPzmjJH/T/QPEdgkE/50jhAIzcwZc
73p1UL40lMVQJq7A6h216iKmqZMUiGssHACRbamYWLA8UAuqeevRohuVJkNj9uSZE8sUT6YPntsv
uB+kc9ubY9engQGUs1VCYZkjSzOkpNAq3PRrWAmLshztHUBvw+geIUAY8g87Xht16l3nfzgduv0h
DyE8/3snAwDYmSW945Niv8gPqqGnuKmrRQjSrMqX1dAsM75gDHpUYs1fPFIQRHzcKbtHxZEZwjFk
ZGCh6TI+h6Dl7WBc7CuRT2U9duwPhhaWQbanrG3gYwwuJsrVnz7jCU9riTjLrl4GbtcucRhoLnVL
XAV3BOJFxYPw3/CNnaDdCWZI4EtEKD+/YB4Xj2arNYf6JIbLV8MQ/eW5wJyVO1ikbWYCRffxiPXv
33TiuVgnbDX5IQ6ygiNiNGW39zC+LmCHQqu/rA1i5AS7Ygb2Tf+J6QVXtMLCAR9yWaiEAEx8/agc
M3COoXycN4usmHaGR6/50AdKsWFyEtqhGaNzJuzLHozWtXXiSLoCwC6UxAaPO1CQAl8u/SJxJN9A
s3T7vaygsV4voEYAZk/LdLmvSGouz6dl+hMmEh0OJftLAZN6ijVLpfFj35nYIZoCzLOkvg8QvscI
DBjzYVmn/fAkxaNglobN9/R1BWdjFXTjpgHMNKcvlxGZU7Ce6azFPaEgtekl+gZ/uz+zPSxOaGU7
7+6dixf1HLeyH+ND0uRzUgxRYHGnff74eJmppuzlbkKjQIil60Co+Rh/RuR8NcVP366hK0MzPuBo
mxItSY8SgS/Rd2RZEuhEfPysctk+1pU+njGiVYKyE8c4TVScZS5xWcFnzmEYJIc4StSUI2O3wCG1
ehKPbJ5sMoQpU3dbbHksoXvyudag0luH8TrY8oPOPQn8CFNZ8iKY1RIDqTH2AXghiz027hwt/QKF
MVNJIgV+YdpA7PX/1yw71JtKAuASdbqDu1fJfdg7qWsGSm0VNIKUmiR4uIph4NqadffPDcDI0QxL
acwLaomO9UZSExMiU8VfIDD+keMPiFhDjFgHvxXGEH+UrvIUsrRp9jxofOVuu5SCr1KnHXGfuAk9
Ziplh2gJscr2Kxn6kZHstOosBp+BKHiG5xmG3LZncsHPbIq4GmK9dbAjXjOy1fwZ9S3IpwX1OnD9
n2uK1IuGiv9Ucgv1Ijlg5NEHNchdP2zi0brSjUCYJOOk9RNsa8y5FxPwoc5p44d3GPuH91jg4PHn
iISBcFjo7TgRfyhvWvSCMDKdaMAdCFAcMW+iCJTigmL378gpjMb8r/AJhPG8Bt52DtHF1l7fDZ3U
gTPJ9xUItZMZdcIg6bGATjfNQhrWG+o8Vyh3VWQ5Gvf/arSE2H3T1XaRIfjB1Imd/OaAhLOJHB0X
+wzq3uUxXaXnxrXjgLaPbD07EcSYyCr5TBICEqH/intvu0TC7BRc+z4HSdhjKlz+jYQl6l7rCV17
DRNOjVx4V78Mancb6d802xuNkiGcCuqFO6oXjaqgebz/o7Jp2clEX9PGbzEhHPsBIhEXGfUWtMAb
mWtONkcuwUTtwkiEL6xZgkvrxjU3L7JdZeb84wlu4/I0ItnVdpiEq7fphEjNq3jRTHX7B5WhEmfo
rGDqqlzFKTaSlcua6g97WhgDPlM/FlTLAHQrfxxUTkoAW8al1S21s+YxWtsxdP5B9K6ChJnD3OuC
zTNcqtnef0Vpc1uT9GHpFREnQKWDylouidUowS6wy+VyIgCuk9s2VBEuWDz1jbGblW6ic/7U+Av7
ouui1TArYU7+7J3/bMUpKX//tBjYSWBxkIOKmMM+pdLtUIYn2qNeCkcc2peGr7hGB4/35N4bth/4
UW8zLEbuSsbIk7AZoI7iqk2c8SV1HBhmo3JXz+SWm1KpJj0m6ds3iyTTtZB3byhgsvqQ+h+Yjpof
1UMZ9yJ1sNTo3+b7hhHpOWhT80xlOD2DWfvop60ebjDqmIHW0kfBLAPm6+eMEWUOU2kXa3MAlj6U
5qmKV9hN7gKLFIYEIIe02cDS/u5mtN7ZxPGwpR6mS+B5ZoBjy0GFqW2YriXEQQmRozFNpSjqaOhP
rxN3O3LOKiMVeYJp6htmuSWVOkbWQHanM1gFR6638WDzNDFEwIWBTy3+HoISwyjiLzIxck8xaWaY
v0bJ6aZYLn0zR4DOJpuSdIt5YUGsQa5ci3764/pKMXF4cp8sYxoO36XhvKop2QxqBqW3bqIFasGj
mQdbPSs0gUBZq5mTY39Yb8HS+xFiQSCHXfM7jUBnABdT7IgQVkTLuUv1eEtuvz3W7hxSVtiRS8AD
rodJ7alDBKk8saAlx/9gv/CU8FqX3tEVGiTbaXQtC9kwuwQBvLHJZJjevxJRATq9jOwxM8m9HS10
YAMqTQLrDF2e5z0rUmME1sOr/9AohkzB1KSs1dmAiotqrBq9h5HgRJcTBu4z2Zcg7lz4iZe0elXl
jVtU86h6q/aSzaAAvZ0/bB4jXZvSZxA8ngBNmVs9p5mZ5U158J+dqXcIHemaDllpOfE75DIlB110
fq43Fw3mAj+cryogi0unou2nLS5Cnq/Mr+LWb/9aUtNVACnPH7w3PRH+VFNn9B4rdz2T9dFtYoIv
3EDfuCCNxGxk7wyBNj165MQiEKpWqZOyxQhSIxjd5GqwLC7WRni7WxtuhQBFh8/oWQkbfWAsJId+
dser4CnDuN15okLm6amyilYqbYmVdqIehgcmSl9oQ9u368WRTsfrRsiy0iASzqkn/4l+ROgac4SK
naf2sqXOviskNRyh1xB4TI/Hlkr879Zpw8mNTK9BQhHCFUHXyVZ1unsZd/UW5HEQLz5cO4sENbXX
8YQAMIsU+kRBFEIebWia6kR4YvkgQ6tkJWVboollRNgHuYPMssDxFRoUx2esBY6YElKMzIuqy52i
lQPYawMiXt+C8dTxVPNYi7dTku1r03SlBBEtxcQQYwfgK3g2HTR7VRjL6SBJzvIB0uM92Mh+oRPq
7Uj81OC0ZD8bTc7NMTLd0dME2e669dS+cSiWo4eWygTFgcxecGD1GkoIKJ7Nh6sDtwI7TTcv/5li
D+/ZDoUA2/LCK5XVb7cVqTEsgjFQUhaGGFb9WU5NpymkjqU/3kZ6Bw23UaMGFBuaWe+O8TS30lur
0DnFMZ3kn51fH9hp38UDkziwx2J6GTEJyGSFJX4zgEtIQcadAts79wJZS5Gu9knFKiqLAob7vxvz
tt2SP/MfJm0ADUux/S5wFNxiexhP1ZmZgJxdxZ5U4CRFbD5a85hLYEnvrqnmWgee2TMflhW6BpSK
koyYJK8BfMIb9aG6Oo1xbvCQ7IZM+ob64tVZOh6mWIRPcNuSSMPpNGPFFYI+1EyMssWs1w3EYnY7
aBsNM+EVDlH7SvQjoB4RoRTOceeqFAe7BhZ1NHbTMec2U0WmmvL+pOQkDA85xeEdd7u7NTR7ciA/
xpaPvT5nzQUhEKb6o+E827xJpEWTRIsUx1r1uXH1cMXBg7NJ2+vG8zBNGhKbOmauBAIDEpCbblj9
lI+I+a+BUIG1givXk1Qvj1RDEW7O8qD83826OdI2wxSn8rVrDOt1tpxo1SteEOQmMlk03K0zw0B9
6gbBhPgqmvtby85aQZHKAf3Cw9r19Y50Ff1UFsxTm8onoVeIYMy7cOsMHfbSJZBu14BE9srXpbUB
DIvAwQz27PuX6CCDKFIbJS27Xcc44F3nExRa4CMe/oBgS2Hs7oRY4MHiRB2IRahoUXARsGQ49ldm
YZS3b+zHevMBH7+C8iqEpFGfifp0jus3ApsfMi5cnwZDXQDIG3ymrZnrQaAZiu9biKgGZau9zsGu
IeXsssnw+OQt1TWTmYCRxQBPZwk9AGIWW4FsufAarTlCnra90FMGtmlJwg0zz8FfbTSiyjUskU8i
CMlkki3C6BPhsTdcW4O6fJogPKqLfb8IH/IxYyvsc0C+NY4A2tYnLTiP5sfjd2+uSg2irvrCbEza
2CD2g0CVFVFc2+LZxudTTRP4IrsUfGO0tQfz7DhaXFkltjaU/EkUlm0Tl8xjXfRJ2oVhgB7nekj1
CFrj8WjYHlzf+9MVKfo/wSHGl9a/1lMEXwCp9WZ+J7ZMIakx0wMfbDBt8wFqAXLQyrFy/0gemH84
3EHZh572ZBNX/E5Ce7cChF+Xn6q8MNJ9lhBBI0C10xAFktdmvhhrK79oFhRLC+UmX35DoiI82enb
WkJxtRrZB5nWpKC3Avo9uXOJrZOh0pagEysfkqpsAZ/dzlQRWaDU34bgs/hUB/em6NhLN51ertYk
9FQ1X1RkCCNED1/gIT/sN6SqojkLh3/n31y65OoIeN2ZowrBBXoI1ZrYvAsP1Z5PL66DgHDr1sAx
j2VQ33kyiQUok99AJKHmqJ0ufs/w+mxuiX/WyriGPsSNVMRKhsr8q/ol0+lDVwulgtBWg/80UHCv
pcKp6Ub42wwDQwo27GNeDUT6SNSQsTXgceg5pwm6HZKcDA5OM9W8JwkK+0qqyUNdIyKrH2BMq4h6
Bcg/Mms4h6tehWB6Z0i4T+JL3k7hJ11G3Fs60B2TSZxvDeUUGZzQYYpzCvMllo1IhgWimrob1uCE
SJRrCLPQnWasiNpFQsYt5wsPADxJkz+uFpol5/c9S8G/pCZhlbbIzHW3QB65h8W9Ta856nmrPXuF
qQK5fgQpEgYBaypNDPYyiGMxX28tH0EoTzS9rPfDxOMZrGQN96/XZAo+WJP6InTq3d/VoumlMfvc
/9PoIGZqM6nJFJHuIcThGsaQfRU2LhUQYE/ARMmbdt5oKhxqSuPHZD24OIch4r6rIjUNkFIYbx/S
80EQ+ZuIxS3CSDgaNjn5+h/O1nWMlxD506u6k783ZnkRLpnLzyq5PpWdsEQxdmPPvBr6JCCqd0m3
UJDBVuUK7pz4flUPhr7eheIo6FnlyR1eerVC9HjZ0DWGuRi7sgArVuwy2ZKpPRIS188K/KUvbjke
30IT3PgI5M6oXe7bx+jYQ0c4SyN9oAsVJlinGTE08ZoAMBib9dn98TDhm+xKSSl/gowHjQGIS3Yt
1p6F/6vXnTmtWYR4tp3436semKM4iFCIqGbFcTiJ99A8OM3q4GhrJMMSSiF1ckp6h4Le0GyZCqn3
/h3TxabVBsBYkpGfG1LuNzUE6u8iH76341eFRqtcG4fFhUVxpqUUwqrXr8v/YaRCLs7IxKNIL1RN
lpczItYEfW8jKT85Yk/MpfEMO1FIJq8AQkBvWr4fCuppmJc7Mt4Cw1VqlFQyT6nqJ0qNfLpCM1aN
ER8RburLRkOmSi6FNkap2T5ZpIACyWZD2mI+eMyivbtXhC04JtU7T6nbxKwiZgQ1Jr201PS3Qaun
HO2rlzD9OuDDlco/WQ4H9vDQC3cyCsLEusQ+C1FVBzTyVSc3Mbgk2gVnkCYBQ2KMIM9wxBBhrggP
DuUK9aXRUAmSd93dV4KG8tPIfjNwoYud8moaZBTfw+2HKk1oWO5Zxa9wmn6Yvlx6PEnEzZvWpRA7
U99X/lEzxfEcoJ/OXusMiipT8TFyiyEqrduzeyNCij7keEcCjybKvLOmYD/Z9zr/fU1JHIP7/ReB
xEwWmePstBYg86sLK7eQvP3FD/2Mwxsb6jYsdow+zcZP28btH8ErErTvwh2fBw0BNXnRsOL8oL1t
fRhRUtYmtRs9DT5VR8QvqqHrnyJZOMTTWewRdiLVc17OvmkhgrWkZUII7tgiJQPhjhmq4LETcVqD
VH1NqeGQDx9YjDLDUm/x7pmiM2sVlzdvPF7cU21SAcZqpjGZlg+YJEZL5N1mwm7sDH1HTDyFLqJB
SioVD+fIVIu42tbaGdEsz2Y7AJUwFfoIE5AsvcbDo/z8ZFTSODC0Z9BtT+7rlrlafE6eXD3VqxjN
zocL11JgGtZC9eygBD3F9J3mGJrcIylW+9d22fyrZAhmRHtksYEu84t4XMm5j/gba3n7Y+bwoyTl
Yi/JhqsRtkcsECejhNwuD5KW2Um1QCLq8jyrXpiqT0HwGQTBCjNxQZhRFeKHj5QGQLP+ZIKmeC0r
cNhMiUeuXH8KyM+XOSyifFKUXi5TOq6cTRceF0u20SeVZr76Aldbw98Kkvbi0V4iK7X7XIA8iiJG
7p0ekdgeLu8E5jAXJBMtAcbYW7yKHfYxtzrARCTQS3OYKYeWro4N5XWECw6E0IWK5BRZVuRZVdFl
kIBhh1pBdHgQKmQ2vedR6qCKSwRvDoQemozk9ei3Zzhq4hoDaOF+XUf7Tqh5/jeiG8vS7oLq8jP1
26mG7Yrtz+kfUGu/rn+/XRn+TbRehPPqonMZRKZw6CD0nRmSCaacSU6m74BLFYqdNCj8ZEmKaxMp
J4ZZLKfyRn2yb+xmG6hELnvQPI7Lb+2YxSBYUrv0G+8cCHfj56m41UgdEdO9D1yOa56o6ycKJfY0
6f8z/Xet0mIoarpw+blQP4YegMUoFJzoVAdYBBayMbP0Ip1R1+VfsvSWVX3cxPc0RSHdnioMe67S
f4pFZ3T0t1+Qt4lT6/8aRqZvzFxGvTVYyP8rFJ7encOS9602sSIIliUC8Qpi4dahjmJButR0/EV5
T7iC7wheQ50uAtgoGanxiAuSc4xZl7otmmf9c4Mago+uJs8W1Ait3+1zfCpOYuCz0TTZSMj/l3U1
kv2GngGiyNvg+6ibdCvEiksbJlcAP7sqWbfT21gl2sPsXlQRgdiatjjRd26D8Q9NhIaOdPYpI6K8
Jyo5G0s24RBfbQMg3xQSrwI8Wn/fXImJgz2oeubZSyJK73LEz70RPbrnexk+1/2PZxtfpZkH4IQq
jv12D7N1ayoVYs6C+hJbp1b3smxxW3L051WfnEK36RS2GUdUfUwVFRtOEE4GHy+SWBD2jEqtP83L
LGCZSj53rK0uB+AcZqvqAiDCi0kJ9y0yUs0BwRDIx7D7qGdebEy/6alkwXVclt/n0ufYb605h/dI
dWrw9k+o3p/sVLdPlHrbID4ptpbgabk/O2xryLB8rPTLMo4QZFoB8VYeDR9tr8PFHwEiowcBlSmc
ARcfFUoNsPIEBejT/TJs+R3ZvGfivdYWnBoAooVsKA0Lo/BLAWbdRgask5S47JPtX55FR8hqi6fq
ktu8Y4ZkhRypScJyLJet26fPPXS4sNtT1mTAwwk2PIsicA7ftlubNYBIqFop8Lwfjms+xqoQk6pr
tk3JE8duYcb0FNXQaQmNcyvws5qQ/RfO7ddzxbjh1kPGOty+HYE3bAzV5rJIRs0H+5a4EEZ9H27s
W68eTPvG1NxTZWhOzj4ARwj1vVouYMilyCn7hMl374/bsT/kWacEeTdynfw9AERvgyUMw4d4SLpG
ih/u7QYSZiiG4CHuBRYUeCg9iFJWohESPHoz337V6t6FaUwOom5B0P/hgAUm+TtOPMvZv8wllnW+
JVejIdrzJ0JX9u7S1ho14YD8gFU3wEcd7AWc1/S8LXUp/2+u2Zf+qlHtgAmOEpazK4sS3c9Ledlq
NDDxzd2DKM8J/GriuWMjPSHx+6yOeKytsyQYkXabKfxaHje0Z9YxK8U0TAQGP7o40PEGylazrT46
sBOYaxVgyGjVl9kmXlwooiOy0AqKhuA093N9X7HuwA9gjiApzO4dcXsC7/7fZ2tsdlIrSwP9jsee
rMQOtdbN8HIXZWk+kJwCJTxRP4aknJYyk/P0hUMDreKdRVYlQkyMHvwnofDJ8Czy+pmwNy0KXT+2
RsnbLdqnRC4VBFVYVsTfZirrsXc5cOgEfwpyUFSRAjetzHsJdd9at+wZpVsB6snHr0Gn6EURZQ+x
aTTW7S0XtbammvBsCrZM0pnXH54vsfGZN3Jy1EzOtiRqoMO48THrGegNEq2ifYyWQA8mGUDmB/jL
ezgFMp/OrqDYL8VHQ39uinIr/uYYTMAHAE4DAIgeZ0qnUX1eNQmSa4BqWchVfS7KCONjRKd7F0CY
BYQSFhZb+y3FDt66bp4kLq6de/Od/6b3+M2DXMMGpmmgMqRvgpXEmAqpJJmZMSRuEmb+cfkAnS4a
Yj5LJye+gO1jCcrPLut5YM5JM12PImaX87craAb7dv9dX5VxxEOAvln+2wnrinSRFD8+aHwU1LMr
qAzuWes2uBmyprePCMO4UFrHJtdkQK3ipqYXGU2O84nk7LulteczP/pUryeM14i61N2Cytn4Tz0B
EVdIQdGvs8R+xeLkZcPaYeoHBNb/YMhkxEaifvK3KW+1LkrEFFit6mnu37xT8Pc1lHLtvbEIN9AS
eccnlLUMrUpdcGhh48y//1Ug2jUns3acP1uOlIM=
`protect end_protected
