-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
k7qeO0H3l8LES56uP13ugSda83fb3kTWyuz+OIRvvJjVQojTSsw8q7XLptN3ghEP
SNuy68sHSrmBN+s/b6dFLrT4DfXRlW3wczX+R0jK7GHsMM/R9k6izPGK50jFzshn
pT//8EWmIUlKcmVJpWG/4lNzfzgHVVjp9ciivumxBpY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 3280)
`protect data_block
Xbv5ua9hoPlE3UfKhm8MzwH0JQf5MJhpdkrpsDqDXiIoNudzCGJA4o15znSyuwfA
P3FYU6Kr8eWNwVRy6FmlTRuYHvupzuDZuZfkgXJRnQ3Hp7MxXtZmUU94T9ooZ2/H
P6SBPrxq8mDeebMZQNy6n+8aZnHFPupk/vTlrzUydSU3yLun6rNCzxXj8dnvjUsg
0dS/hq9HkiQsoLPNsn851hGGt04dzqj5kLc4cL9OYApxeDKX8L/Xwvkzts81iBKX
U80nLwyQCkgtyn36m8GklV11f5r1tr4um1NDKYbgViZ1Vs9vwJoqzsIaCSNaSfTp
5ydRWJ35D+qy3Nnbw5nhzaL9djOA4f1hOOZJPIXExJDopinqWyOR07+DJs8rHYO0
/5gVA5oAMaCe9yiDxMVA1epDwMrpa4rW+aH9mRw8iJo+HVbxCod9l5KwszCmh/il
WWKTbb2YdvdZo9W55wlyVOXYCKcVwfdpp8lQRhlVBN7KvVfBh/wWVQhyLm+HtQ8j
IlLrMZTL0MZxr/5qoMJq4WJtoTDACxJo9rChiVn4klF53HeDi6j4V0W7vEN6LFHe
grxqUTA7F3q8+m5gkcIBxeLCbfKMJSVkDwQ3tuXnaSmU+63Gw3E7kUOvsno6+SaH
xHIqG0YlEWuD7OeFhCrwtjsz8JOWNx9NtrkrEQzX/3roxYNRSyjGpD574Ws+fbsD
Kw/xTak/ZdpSX27mhd/vsaIu8K4ldWde2IMlX4BZRPaE8azTJH+Zi6q0s9YVUN0u
UkCayYCyh2daYAfzfaTTNBRUDLz+Y02Tkhh6RQj3PmFu8j5GakoGHYLxqyZhw1jN
8pRDmCRIm1HfUdGWnJm2P0Tatwnt8GCEnkTwQcFLIOjb14PrwotyXRqQleagVBqP
/pX9EniNszo3aIvYS+VfVIDOjWSOGIQ616xPXfDC0yYQkrt85t+gRu6an9znaqkY
gSQFQpkEBrQYP+Li0pbPXVi4HgMiQ0Ol2CvlQGgJsqhAFKSVdpgmoC0YoFkbxb9R
Y550vljyP8rqGuvh2JLH1IF2AtapKExcQvIUgFKGtGH/hZLLxFJaLeLycE8/BVxu
VVMupKAMkzzfb977kh5xVVoeNESUTEg8nvthK/7dc+AeRIuXTUs/WPyxxhsoXKCS
bhhwmA7vm2p3Nl3F0tn5dDc1ZHLlxTj+krv7ELpx6jZqQoGpOHyMABY09cnv2IlG
dFmv9dqrsQPVC0CmXb26naaWOHJD0krebV86GaVBOsSeV4XQudobbfdEo6eD9YnO
EBegrqmWkafy/b9kPk/zTRVEfinHDcH/LdM9LgsKePVbQnXpEEMal8p/xzyEZpTo
uePWmaoRi25jR7c/pnv51ffu1WvSN24nGd2pun8cWDXPIT2YdKBNLUGA1RxL/Pw2
/BLHdFdoKlnUGuRCRAG5N8qMPm/qHOF4ZOqZkz+XlIC3mIoIWuMqQPpen+cRLcR0
aGx8czQmn5glY0b0X7zARWWpFLJDceCtUYfkH/qdSsWXfthHSOnEYa0ACXwAaC9f
knSyfaV69DIpenk2qFEVSvvBvbgA9ON4ZRdu0X0/3s+VKU7fz7VJeGH3jyXQhDPw
ddghDrCt3rEnBdqtJcY5WXrp9pwx0fNXAOIAdofiBX3XwvcDo/XgwUFq938D9eGe
pMxwDzufrsN1/kNzEtfsFtcYlpajbF3ftL3qDhXll3J1MNP3tqEmJhtdm+l4E/m9
QCipK84O+Jq3SDa3m7aaPUif7WRhmFY0TK3V8FqRLUwE8j1XNnYJTcVDIusohfvh
laitFOFkSVgQ0fZ8q+GQHR/cypqcKSLuVURTTNAFuUEnnAWIwDTMPJKlrMfAK0n6
jXS9CKo7bQZsJtX8ojxCRiNPGj52FLRAsdlhrNt0PyBQTxLloAnfckmSKurLgeMf
qKVtd6aU6l5QJZuV0Bb7NsTV/Ez2Httj+PX5QJ5MJfx0B1gycPSUrJEVoo3D382s
IC7QLCP9iv3o8ij/U7L+6HIrEpH+1QIHVQDJGj2SU7Ia0Ov2CYYT70Dvw9lKCO7A
wxCHnuQTHj+5AGghyeLLdbrzFmCP9fZYcQ6k8nabvDWqqGHP+8lio3fGNNkOlo4j
UrOspTunKYzZ9ay8sn8qgEHNzaGoiEhk8yrNqUsgIyHWXe2orY9Ls4l6Y/kPcrs1
zxxjFtNe25iUHPx3yXRKjtbInMwsNnGJ1IFQvu1vjr5w1uiXcaJQhyVyNn9RBswL
ggkPAVNIw72SVCrMnOrDf0FaA7CSd8KbdTYE8e0cYmuCbf7hQYvfLJZlUUSTKmaT
4Fvq6lv9Jkq+Z14cW1VoGIfgyJwZ2RTNwFhe/bRXdrhL5COoYE5MWZ4NRFRm+G/+
1bSqrWPbpIt0v52Qnv/6TL3lc3w0BkjBsn0YXxL7g2x4BQ8AWrgq0IKmoSu7HFic
aT7tKkGblQRCJzXPqnyZohHSqlx7mhDFCaDQJ7h9YYhIgycPuevIc8eT0jQ/G6fC
6ceq68KSazt/kCqCnjPuYRhP2DSDbbV6vu7hNu5ts/cbRvd7PRnxdeSYQk9cGf4I
HBBlIsXaYpH262gnDE4O0yYzjaFlrjK8b4L8D56jJvBs4xREpd7jmepPi5qPxnS5
gZ1zJbpeOwju1pU+1Sg7d4lPeK6BwLYrAnT1GhE1aslmMz5uSbe6p3VJ/knSbA+Z
oCwpPt0LKKv5/y16SLD43rE8B+q3GJ7u6cc6QfAj7EYtoyoySxWIrYdug8Wc5vul
mDxLGjQcF61eRG43DY2XBROiUDCiAMGpksKmqATaaEgvURH2zR+LJItg44/yW3IC
iTdX3DlVmWTbXSOF53PbPxDEx2REbegFMHf73z++H8Pe7fzkuXTsrhoeFdVKyiox
38hY8mA/i3J9GeiOnHzdmHs2Ai5KCYCao6tru3GJDofG5umEbZKroxvexVvUhoG3
sqrgsvEGRPa2gdh2pkv++Tay19Zf0wB7R465N0KM6SBaLVthbMb6FWQ5nZrnz/1C
g+3MzZ5AsdoU05QEEaWD6fRloq5ZSHxKtntP7Dd54Mx+9jVScW+GALS+NYh1N8z0
b2hPuZ+BQ8+Ofndkxlsk6clrFMEmuoGed+9ZlBtZZWF8Op8vS5KRni9RvX8TOSaa
tQ/3NSe5gmX2mP//tgu0lDKx3NqEesoTsSzPUSwdvKfdzpvlSWiSR48XzDJW7dQ+
Ee3BDWQgZNsAQ5VRZrzz+k8XtcXZAze3Td5yOkOfc/Is+DbpxuMhlGCTHc7KzbFq
W9O7sKNM7U4B9LojmY2pgsdFAOGizcL+nufHmNuQJVgT41VQDp5+xLMcu0Zx3knE
X/VqPBd4iG5hZPxis3IqL1M8vRG3fy1W6FEGhRNx8kWMGSfrWFrhQyZYjw7oxepn
lxn/mE+qeK6sp0apGfgtdDQpCanHmul+XtdpGPg6F3hY5Q2htRitBL/8xSHIKJn1
Cmx+F6VbqdH4XQIkaM7kQrmJFq5t6bosobU7241GiNnLYWuKgbzKIpVqpoo3oBAW
HatnRzg7YaTHq+NsxM5er108qHU8iZdf3LdK3Zww2bRrTkPpsXmQU1lrrHLsiX9n
XS6rIZ0MYnc8ZL7pjM2t4jcCJQNRjyZ70HRNk9pFTFx//Q+YiH2ai0I6rou9qU4u
1JFvFIFhzeKpvttTuGKbihDHBKMFklsk+gOWVbtPzLGd/RaIOyj6u0SjfDl0l23k
vPjKkO7qlFapOFAGAhMA2D5aOHel3N9QmF2tah1KtpeLPHezFFZtHa1xLL+WuXtW
Nu3AyM7QE4alITu+SDr4QZuK1H/LD+ay28nRSJgMT37zGVoFIKXnYQP5/MUZ9j8u
dvWcThPqOOW2NzvmBlpjBROMRHSUD5kmidSeaq4w2P1Ma4aQmNQ/MU9iK46tuWHO
9pm4GhzEo/D10WNRfLxW5MPMY8q5LUuIDMe8JiZ0W2myxByKME8w7Wluh6IJdH+e
rK9Zm6goD2F7IzB7JSv/l/A/ZmpYA5QfZZdtl1Enn7LcMJyNBOvs0kmQ0GqK4+e/
BVNxImj9hoPiTGS0vIR0FGPTnQClDreHcEel8VkOd9O+MqtBcZiG/OxCHUwFK/u1
S+4r6DcmjLpPtLAo4oDMmMXsvOddFOFaETJoF9mPBZ8ZcGoF8YIxhc+3yYcXDgkl
PnEYcJCeDuUh5cLcmRjBdmTevd1btSF+ntnErvhkgGpn6aOJq5p/cfyv8vN2dhwQ
CNbfuSuCmMiP8f0xLF08aXSR6Ps0NM9oO/FvTHlwAf42NgN8o8iueG9aoAVc9l8T
jkWmbAgM8V2yQhQuPUw8R/BIcj2O1zfyb/OkiLpYPIEnyIs8mZLjG17Y6gNkWvGd
IT00eYEjsA2FfS0G5R698Q==
`protect end_protected
