-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
BY9AXwznp5sDDXkITu9vYzWI8sQOg2g7ZEIYvG9bXtvb9OitIkFscX6jjetKP5s7
urzstjHkicLsYFQtb1dQ+gzEPPLWEo9i8D9cyBeHvhjU9Mywf37EqKNp6LwUnvsL
zGcI6gXXktxc98q1AQztajVd66ui+Bqh0bc3vokq4x0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 11519)

`protect DATA_BLOCK
w+r9iVq5l9nk0fWjisvDDpw71UNKgSS+r11TDHxd6iKi5BgP17IgbVwDj6uqsJ2l
kRvCnXsng71vNKKi6PeM/Quop5WYpCZaqKtX+wnipsvmPlzRKqDu+cRqZ90ibgph
/NSF7MbCta6gSXo6O57bAPhKTMRmgO/93/O0wI/RKD9IaSdMTF7TyRhajE0cN/o1
F41cRmvV8+JjzP/8RLblsj3uv7LUd+HC90wU/40YcS00vKARy+kzJSrSXp4q1tcO
O4J13BX+wJ33E/rxZ3yTUaB4oLR99dC2NZdsT8S6gi+A2GJsFad4R6ByisC6X2zy
2tyT8QX60qLDjvj60WeLoSmrjV4pGNQ5Oe6tbZu0XzdS0PLLcIA0I3OJ7lvTkTqY
ZGn8Q1NXjYUrGTx8IAgCMNPa6scVBlPIY82TFyx4lT1vjxElaq38tTV0Ti8p5xJW
k7JN2xuDa1kqMICatKdqaLRerbTxoy+0qKr1UFv1nVnIVXIsbpjQS7aUvPw78gC3
eD3aLZJ2kBAoF5bawlhXWaYHgUm/RGG7FNKAWmySbXpWHbvK3QSx1L0HJXSWNmLp
30kXaN3Yv4fBWdwn7Q9hVz5AztJhGoZbQEAXoHGurzjUbJNSm2/rhXXnWInPyc4V
P6qZJL/C1xADgOIJRyaUTAuQY4TM1+HmtEGhl58dRLVZCEEkU8PmNpRo14dNkgL2
UL4WQSxJkmr4Lmrv3snZ8h7enIVaBOfwH7LgVfM2m02xM1meugGkfXeh+VBsApmP
Z6d00uBjpfanuYQPY1J368JiV/L94XGiYlVWC86PqE+aeRQtwYpRgm0aSHcRVkAk
XUYjdfwypCoJQwz/shUr62OVU++ZZVLvYCETST3dEApDRJTJmyfXEKd/aW4qUiJ3
uQZoM5f8NWLenqShmhZyVSbDKb3ShLKbZYTaDrzoDibQ2PjWaw4e+a37/z0oIL46
8e2gVyGXHGJwA8IZUUQG5y9D+x6Z09sy7KCkLq4peZdZjSeSozF834eKrAxfIV/E
cEC43/KYNWI3upGwAjbas1V5Sky9Gyu3q8KtlfTTrTQghvWH6OVjAiVyeda1iqyU
CjkQ5PS3iU+5FjBvmTZFhPxJKdwhjkRxjgBoD6CAa1o37YyfGIXG30ubh0jw7EOW
ZfBbgAXNN+8z+f3fuHh+dc+cQOx7WVOvyCrnCg81Iu2i5yxNYSO8F3jb/fruJuHA
ikp8OXfLFCqsn2Qi/lFae94Gy6RHVgqCAyF0rTyopjIyaa9mqhuhoR7jXX/36sLc
rSztiH1uwqXI6NaQxx0bOJsg78k7UmNOyb70cvDKziOcQpNOqQ85Kuhl5GC1CQMt
TCs9NxqsA1k9eLqKzt/hHnvyr8ZzzsINidZ47AUydspQ9LPloewZxkObD/Ce23as
eDxBGg20s2L4FGbCK8bFxLL20z+arwtCv9gbsXsS/GO6xyxTT8eynQqKzYJ9Wf2y
2ikBMYChTGhNVpM1kJ8wQa2Sylei3zTnzG2Q/OLjtwMcv0vbpx5xIKERwJFA5a+V
mJxVcSo/C9FY3iXAavoMLCBxmF0c4VV/V7RPxIkdtiMqGkJkMmj9G7ZGt2ABeqgD
wH3lsGuMeXEFiDCcYmrVH6GEabw4PqwtV8GTL6DQD84+5cby70lM/kEM5d/s612t
aWbVnt2GA7jwWNNXSEPXUBer5c21zHRnf15she4RP6dgPebZbLETsu53dESTlR86
Mb0KaxLihTMNGroe9LORUl2I0IPfCInC7l9r5ugdTCJmwpoMXtB5kcQZJ1d/jqEY
llkGWe2GcYz9Cejchi161fnsjj4a3e9llqYwIlLsYN5k41K5I87ahZzV6TJHOdtk
lO21MDjWnGrvQMg4Ps218eoh9wZYiFiUQzz9+JCOz3HlztA9T552zmtOgecPhUg+
9Q57VRWiovpuUjD3tzonXDIpZw62V9dcPQlSRPm2dqfexiv/o7Dy8YBwRZgpuyvm
PEy5gjGQVL8ytb3vBzm6oLL6xH/PXqOrKRKmP9021SNZcjVtoPT1/PnSp7HsSYnV
bqBIaZbJZZpSDPEwg5R8UXU5YCgIczSI32MWEIAGRQ5FXPwzkaDSatJdAUgf35ww
5xRNPfvNomHBaAgmhMNB4zhVAuQJbpDpXdoz+/QNHY1ay0nubFB5V2CLUhpA2kQb
Gg4jg3qHQiGM/K2OcSqwWParSTCulpxMarZFteCClCcCNAAKkzJZqiLWk6wvi8KK
XF4pVS27zSDGj3v+vUVqdZWa7xB+HdxM7zIM1Noo6fKkAC+sdB66ZeFCoTQc5pdm
w1ata+GQFmGYF4dAljuWPzKdoVgwlOfataj/pUWBeOE6hehaAGKbKqPJ+nBTpLwG
Jjtr1k+DCc/GDR0AgLRSg35JMAjpUXpDKnt0zBWa/a4nUZIO290UUtST3ExiMtql
sIwc+lqPmnS6hVKPbzipXd8CFWpc/dBnanLmPcg5Nh8/9QSNRi/qIZbNzWtK76rV
kFkD5U3P/yfcRca2dgsGHze7wEE3/cNHt/9bNbWYZ8FK6vFEwdy7AJRoqAn0mW3f
JXmIz7Ck+DlSud5XfR2onxGZVoLO79aOms/CH+rnp7Zcr68wLUR9NdTdxq/L7urX
dslSyuntYYqfnhRPrCHUoEsDO60PtJDQzpmU8omVFCCUzbD2CplR6WPYqh9Hf6W/
DLJTifMxlk0poLOf2RC3DHQDiywDUhAXA22t/FGAmTapVKAcXiTx4LM8VIyaRPPn
rY1FGw8/oCS0fOZktEUV2H4/exbwDgJM38OU6M8L8n1NP9bBrtCBoGJ+zMlqTvQO
Hwg3aKK9X1h3veJJ/Z9z+O4nbFmaXzg6XI8PXPiNbMlbFxiGB0fzFhrdjZFes4rs
a6TSS1dSd/Ba0hjMzmuUbju76eZ2g2W7xJ+p9GU7OqJaPpl5/KW7bJ/EXiaQr9Rs
STSWI/SNuTDVKmflr5x9mb2qRnZiCKZPIINLOlu1B5KBn4qgu3dp7+PNw9lBiAyX
+k+kvSad70+/PCQBvunNGoKmxTTWb+Fl1Ht8TJfaSqVdDYlU/RgKGoX2ot1U2aqc
ocJakX7NzfZHXh2WcathPWcAToI4xemV3qNrm7vhgfoIK/WwnqKDqSdeTI3x9pDa
IUDQDyJA/KPesn9F+sd8vd0z2fmEpatFeYaQWMqpA+M145rRCEOPI8xztUFMQ0/9
wFrwexUbrt3upwFSSI7/bJDW/QoOrKvUtcfMF6Emtapg8c+e53jWAn9pc7fhi+3v
oUrG/SZltPOP0nA+YOGv+WYMNvlwcNYe945Y+Gy7awlEUqZx4QsR37m39whqsmBm
WgmX1nLeoGNtvOnnU88yasUqQfvanGxNk2z6qYXHPttzzmpp8NA9iA6EpF+e11nq
1ivEIFy1oO74y3fJKYlgiLjYbt8mDHGdZtoyf5b1t76Lo3OZ4vorUMmGQnsDW1CH
oHQwj34FUuEIUh2HK+QCrpftabQ90p9giv5xrHPzcb6XI07LFIu2p2w6U0Eqpuig
v9oLe2dwtQijDgVWfzaq7FNd9Q4jCzkLcap8NCJnMPUuZob5I+y2SwzwLPKjBGYA
cYQ+nppyAJauPdfMFmVszjwFA+58furDsv+SMwEyb4eOU6i+CFiOrF9Jd2qZp9t0
8w8UHuVWb1a6BXIFAyZo+SKYxgTj3NHug3wXjOOwyYs6lGXqIoaKcHmT9djc9y+t
jnh7cxlRsPIxf41jrjrhb/C7yBt28ME2rdTxnzB0oTmwLeyhPpFc3/UPdOkOfrDk
rrIzCKIFSEvJQaP46n8mDb6OYmI6UevM3PeFstYOpe36axUOqYlouaOwnWBZow97
niWO9UZLE/jBQ3H1m3yvnqHMUFzUZI/DG7q6q8eVRMLiG62Y3ls7V1ErmmFTPiXi
16dx+t5MYuHxwpdluTDaNDHM4FHtUMxKRvXxHSTjTo3owbR/tSeC1qvH7CVbtIGB
77nnyCdVQQKdIhcn3iQBD1Dwk+SgMaTjptW0e7m5YCKMOgR44NKAXmx4MVbnTo/+
Au5OM20etwKBow/rC1MBMBVC0ijaFxGI/Q66dF5r9qjSnh4gt1D1KHNxypDJ82Wm
Tnl61zVwap17NUIP0a0pfd3yGRxaSvrGBVRc4ID9Y3uuRxygrltdyHQ42JT83ia2
OZLmfQsvSJcidxvyHroh1J80afvwOqb0TAw3xfMf+6/QM4YeExzX3reGYhSImKGj
jcydWzz8MpUTcLffhsmlyeDshkba6gLUqsyQIF2rXl5KPBqC1lzeAnEdAtgmlZ0V
08uvGkCz7js5Su9N27nbs29o83NmHHkszNtg5IKuU7teoDncEV26Nz/MIQ32JVNU
Bjr4dXL/226+XnBoBFKh+brfcq92bkBP3JFUfeK2m2wMrHYAhZG54xPQZUXAEJHm
ZmRhMs8NzHszrFEED2q8IBGAa687YKXV2hzfPfbm1uHmlKgTIsn2pCJi/r3IWV6J
YbTzAR4+hydQNOT1K3x0z4/voRAU/+BAApbXkK6qqdqYVlFJOft26FSZUT0wAM2A
VwDQ2N9E/zngQlk8CItM0m1u1V9NsRlrSZ3d/StObHDuxQhMWKHhiTKtbcEBhOiP
8dQ8RQi46qeIxIDOFrSrYp3P77GtIV5tnkC8hGzoKQlhLz0k1qdJG/oBOHYrzCxL
OlSaOkfXBXp66BOaLnMMbz6q5pmmJruANctG/2DQPRMRDWqGl5uJkg1LK6Qe3hRl
Doxu0oVkzC+p0DQSQkKryOFxsCbU4jI/0eOH5ypnkyyKV7V3mrxalWkJOv2+lapt
bD050KLFnMQXdeXUgJHiDzZyjdMk3kAhdeYkcIFUpUGBg4x6coCl/12DofJZixKP
tYho/QtovDZHsAwI1RxQDO2qvOw7E6BlnzFeyuT6SEYRyjjvyn+5PQFtoHb/p9SC
KFYYueURUgFBkTj8HFtJkwSPJIOAUqUkAIs9fPg5Duc49Gb0EbPnMdZam2VD/HbX
sJ44RMuavBIJfp6pUJaMryn8rx30CTnnyx36dWD2LxOoKdG3+gb5hALSigOFsQGk
Ns/umfalcSCQajUNQtjgbA0eThgu0OFnbH4ebNvFo2wAI/nCSB4QC1Ul+51qs7se
bxGC8XLkaqycynlx4UrSQ1lw3KbXUtUEbUXmRj0r3BO9zTB4/vMkW+Uy/kSBPcUb
6WfNI78Q+2I2+p46+bSyrPtGHO9dBXrlgxXFsJh69mOnDNt7j4HmHVAMKYx3eb94
U+TuHMtkbDE0E/tK5trNPpsEOF8u8u87i+YZ/sDsZL2VNlLYRISIucq971Y8GJCd
OAApw7SjuaMricWrxjFArcQCr7g2ca5WNirRdIUNiQiK0SvShIHtzkjaiw9bLuv5
4XxJ8b/8mgIWq+02ID4uIPUwdAz6pp2CUanoumvR3gyW71cwqeXh6vtfanqgJnkW
d/gk4l34OSwG2CzUFmPsSJici5shU9iU0MakpnoeDcbFrRoIbvtieOvE+l7TDpNt
Nnx8fw8f98OQsPWnG/4HTGzvsNKZDcdwtPCmyJMhRusYp9PZoSp9qzTnK6iA9u6j
dzI9uMjn/AWwby/+NSJr8OV/TY4K/3yceUzURx8rk2ambgtsu9Zw1JEB4wW/iTGn
DcJSsG6ESpiVCh/ZXHmKCbwtaZ/zu/TdVqJDm62u3yYz1NMK+ERC6HCwfWdYyK6f
K3exj+4yVGhr6JFz2k+4qPke91PCfWX/5QoYkcOKXjvw+uFmV2bb5w8jZa6wIHFF
j4CdaCYKWZDJ/aoRc7WIME2rQ5X0Mxo5Y/ppFx2jSiDQZjsGqAwkLsecXNioZksv
3MSD0WEsrciI1mjw1RtsA7j/pEVGAVwNSJPobPgt1fONK+pP/vzg3CXctjJ0K+6d
dz1fKVzGMsRuE1MocfIWUIIJW8/u1McBCDm6jYF7BBZ90gxoVK59QvxjYyVV94h2
68g+wlb/qDJ8ttQVC9aq9RkVJr1SlijR8z/J5UdjRLuV7C4Trjts3HGjFhR03nHE
2ZPK7+fGe/ymPq/tO5W3chuU4GPumhPjrB3l1YmtXYSxuq0gY4zzz04gU2ktj5LK
QJz1LKP7khkLWym592Upe2+Q6qeitAXDs8tqm5j8NNG8HEgBH7xAuJZGILQZuBKg
9C4EmTD3EybbCjVGu1SO0T+V4st8cLIEydh1kPEf6ueePVBSDMXztbH9SGMbuzqQ
tYkQaAPx91/3FbZtUnsG+W6uwbrYPRPoLZOJqHDxc1cxvcJ+2ptpTHlnLd1mcgK6
oHKZoL4beGmec9TCJ5LTEfVUIGt+YnrC83843kEgWfl+fHbDy9zP7bhqSFpgJ3r6
Mc9J3MthERzElwJW/Uukamn56JRvIO+waqOUx/ymaS+UfGb+2L3MSLXvgo7AneIZ
Krm+ZQsxaUJ0FkRyh4XDaxi9WyqwjX5DVDM6Ob2snzOIroDfBvOFfzTgPbKMK6DH
vLyL1K4HqMq7T4NiQQarXuBw3Rlg5m4FxcPBc1dMAebrLuChQl6ijHExGewKyvSb
bjVYrks4vpw9KRc0jH6K1xYjAC9jjIYUjsu5r5oAGW8TaapVG6onzyqG/qp0sN2x
JZ3aLDiNwZmCGscF3aPGRvCQrSRIWC/exEKr82myofJjsU21z9C0ROOCSUtelUOg
OofPIPY22J8doAqvgMqunBNZ2NHHr1tfn2YEjdtUy57LNkdXdw9V86cNzADTCuLV
STwC3tWSIJZD0WMAyJ/cCynFsZdNa5eBQvAZ8ybCzwiGrI/Y362Oaod2khf7jk34
691kXQvg6RFw853D+c1TPcjqxP9im7LjR7hrs/w8R8jqUsyBlranrerQcag8AG6U
50Mnwhz9a9ZClcxnu0JI7ZuA6uR2HFL64oK8eOkSlyMJw3Y6TtJ7DWgo23NvxrDG
6xvcLirDi8gWhBCGSIG50Hs8N3XdTZK095ES4LPKXSQqKiFIkdu2MWkM3rj7NL6G
pXOI2urgoKI45a8KhcGn+wf55T+NUoWcYv9AWXK9wmfj2ZeThvsTmJaSH6HoMij3
uKnrFduzF7+wIVXB95qRXkr5cS/IQRBw7W/0uP16dTyKTqRwFkSpxkacIIIza6DZ
KXsgI+/20C+plqpDJKqyZ5daXQ1cHnDSbwjDxhID0yTJcUTee/36IvBYoOUJiyAo
/AfqA8tj8Bs7ooKJmMcQcNjeQIFYS0n8EcedskRqENqLvs6Aa9YpBjGov+qrxxAR
pDVlVVjSlDJKJaPFb89NtPSXvglQnqljC959HbmQ5qcgpH7kmgLWgqvjvuG8/q5W
YPs/AZ+QXjCP6OyUZmud6/8yRtrxOkrvTZYJFfhPjaTwUZvyKUvmYSe3nAJ0AwjE
sVLljq/N+LKvLPo8zehlG+7cBy2nWL2L6SEHxAl5ssjna5lZH6A4Q1IyJOpQnQMq
y1rkugGd+8wQDxRN6x3Hv1d1bOk0dxdrx+5clI6Yap5fT8jG36azvVFOgkHtbDmt
G3g2R1k7J3qDTN1Xhg6O6W1EIrO0qhwK0dKyEJ0XQUBpFMBm6aDYIfMlgNaD0ACi
bNOFiEbxaziIAUb7of9USfV1VXJrEHDHxfo307cnzUQIo9GmOCoLIABmPCCiK0y+
pJNcqxvEzYeob9dxkq+2NeZazHgw6crJh0fZXe4biPBPaxVZB7i2kF7AUJWHsMgn
Fb5JyciS2NoSHD+++85RzmNXbLx9VLraebyCRVwjf7Ha3ENNE0J0CwJsQnZsdD8O
Ksebr3mfa6oNJypkUSkU9Zeeq6mCdJCDOLiUvNrsG6mCm3GFqUUMfvZqvPDTkDuI
zgALXdAcUNzF/aWw62CMfFNScysqQuvNgpJsu4FTU7sdBJZk5Am9qTG9vVMw198I
JZtUFZICPdrdSmeDdPkomLePFC2IvvIYaVs8Qmot0SpwjTzGwKAToL4nmqKEBD1o
FBH7oRXLJKSRlw1nAq5icwBMenclY1QTd6+8n7xf562YINQ4F1FhZjbIENeWeef2
LJ4DuoYLsZKLcYrXxx2QM3oLt7uDf+XjwlroGldNx4oDmpHIAnPxU2zutfcAYAes
37wMOhnOS9E69nJId4cXXwrxyjGPaVWS+B32tKzsoo/sf80Fs3psJXyIgghxmFSe
KDNwdojzHCof4I46RCsKdO/Xl0eDLi+gkGLgjJO37wMcauq1kAtqwyJbitgJPh1p
abLSJU1XA0EWZ3NBBSD5l+qkfm7mh2buV+LxFqy3WMzoeU03NfV828b0Zxp5XWYi
2YWPl7ZWKgbuX7Uw4/ThEZ1CIjh3cvkknk5voHwOEyqsVSDqStW8dKVoPsYVqTcJ
6UcPggIBJaZN2kyzx80/dVrdoz1p677gI0riQCtQ7hRGBB8NjdxmoAMEF032Y35P
50jDhBHi8/B6GTfee9N6TSG32AY6V51S8P+C7WTQz3nJLqNC3hUt18RDbWLmQG/R
O8JkK951vhfXErdwVbKklvE3wI8Nj/QDCoGh1Tw7tkfTuo8ZfMp7+M4MZld5wrK8
vd68L395nsOBrhojIEE9XZaS545c6hKCeNcw6sjbxtkGpQcUaVFROXU9NJxb38+N
iHo+/RV+/Oxr44imUT2AnpUJLISnNoDg/DSZsh3bBbS1Lv272bwQSzSaP6gTdMxe
M1Xr06FF/VEXtkq8M9lWgu9riFvkAZGuk6JaNAah50oWJt9qsw3grKRuPYTj69Ua
ka9/pxf1Rv3SNopw53jrHzxynsGudc2YeznM0D0d1CDnlK575/R076krquKmU3MA
c4Pg6LfNC5INEkAWoKfkOLMv+o91OPnyaT0SvSGRR/fcp3oP5DKlfYEe+ickn12c
fc9M/CJp5Z47O4lIpZCQrfpSNR6MQfyeMRkS2AC0uZwQazMRrN7WesEc7hGRvdoV
NwkKsMSrA70oDG0fM+IJQTytKe+snJWcGODQn050MLiZBTreb+sTPjbX0Z9GWBgL
CUXhyn9q1ba9ektjPeoSNfgkBK4El/16MpY2EEj5HVGLRL4LEZDiKta0HNf7Lth6
plXD0hzvi6Or+gxi3HcO572cbvgiops6Ia2bdsWN9oI7iHP/UWm+0cDltjejQg/r
hTg+zG0OzZscO3ZfFubuHaU9UBRPVrXFKIwuh8TH+5448QRT4tPBJwqjSaWyQ/Q1
4SRYXSOoQrwpyXSKoea93+CyXhsgpnToFIhDebxTSb1lN3BimzRiNoI34A1mO93y
ugZs3SD8iWcrr176C41Jk+u5jW/LhfFv+5lgnA3+44rMLXPhIg4z4RA6ie7hH2fY
3JUXqOxTRRbZh7qt9yAPCHCTSgWujrUdHfTd/qm0GVDBXJAoA9/ArfImZUV/fZRo
8zpHVftmFwNVWp9Et7SSJ4Gty0l220SCtRJwRGkQvP1CUpLTrBWob/Ancp2PDp0p
/636GZhtpO8oReTarDAEparNuuhjniCNdH0bbYm8r4ForQjkdKf60Jm4dX7WhIM7
mL378GyuX8FAaKc+EJ8QUcNATBBAQnRUYjMYQjDmGOCFuqvpmQ4yW/6upEtqVLhY
3Xmt7XXNdhsd3/ZUco6ZvrwQ5QtvLMp2tqpP09Owi5KNmk2lkkHbHa3u5b7pDGyu
e3ku5LXlskdLZPKrA4ZnwR1BSJ7UnqbDjPfjnaQX0dbmoRRNnv6Xje7CTcs3vP8u
CO7igKEn/mlBCPNxTrGZ8gQvp/8rzttOLvcw9Bzw1WE0jtIa/t0OQMNmsWIFQ0IT
Q/fswSEg8WpAnhrO6yazHaM8SbKHU9+YDNMFOxW50sWBFUdDRBp2f25vhwwbruXL
w9jWIOyaROWcaMI6JRUsnef41+8MSV622hWibddPhk7c0Ejkhbn4cREyYBFYAPV4
Wq1peR4fAwSysQT/cVHD1xwuxAK02zZWk2LMjiMRd2U+Je77nxHoFBGk2RWFOq7M
F/h56jpo+Ep8nVfhHCwtm3+Qn7g8FzBLoFmX12PgPrCQmXdtZa1lOG1gunIpOAiN
9pMIy60oTvdukZG7cb8LLv/pQ/BogCLezmA0Xf/XzxwP7DTdq+88E47CoEY+rjeP
LLRm31N+ACfmpSi02K29gWXvkbbmM32APt01uq02kA9rD+1jfMAZuZZThaDo4qOT
dxV9qEZMpAOEnfXh+Pr07YYrR5djq3vnkGL93szt16tmreaeGXDntF6U83uMhiqB
7VbS8b80VEPhaaN4JipCymu5dROtyg4QOE1Ou1V6te5tpe0L5P/mdg4idT1n/m8K
Z4wYGIwx6W1j7IQ5AnpidEcBSAo/3HZbNdaxeQjR3zNW27L0a7yhSe14iNxg8Gnz
BQk1F4OnHEL/+VFqubQhxDPQuQ5qaQTpH4VXWY53hAc3jWl70Y7UKZATMv1EJ3DF
YFF5JJdRw/+R6jzVX2l8mH4l/LpvRW/1LxshhiQU8FS0QQFur1mbLM5I+LBgAAbZ
ZgSLOJX04EyWSo17nJ4QQNS5FPKiu/7X2TJum4BiuH7v+EQgJZJBK9yKJX4swIqV
MFRHb7mnqLzd5Mrl6bAu6MJb0Z0GQsNAPtraY+9NUudHIdUdci5c+QMDYy8kiuBj
YJSp/9Q41k/ie1Zi6viktnfIPHLWqLmSnbg1eH34qoag8ew4hIg9XG2xIhVTAB7M
Y4SeHrnSRuBaAIrUFPEO25wuM/1IUa24dNqWcoACe6vyUmBfzH3sgjwLiy38aWlC
GZH0QY/yKLosvvQPTIEkCrbqfQ37kddjuQ44gCjJPhcgnImIc2NdZJWmWBZAwb2D
Rmy5b4LH82p2mG+837lQjaU4IXZsr6OdkffZf79280ZqArBspxZGk9+qSFAJbEOH
2NP7PxalDxGbFATHED4id+b2PVbbR6ttPSIwwd0xhEDqdNt9xh3dysN/0heofyPA
N8nP81VKJIyR35mOpcKH4dxOPSNI5YcmbtLzqkdFkFOsy2g/h4c21oLKojFv0R+j
iNX7zEKqVD1mPC/qYYCY/56xxuuZtcmvYMh+KJ5BIkZ9sGIvHBOxlwSgD3UEXaiN
ltccTPEpoRgfeddojxg9RL3+Pv/TBbBQ2xcvP7a1bztpv+UXnuzCxMA5fW/ZKDJD
By3PqWqtzJwKY4JFUSHXrWnfta2KRxseFJZc7PGIBkr5itDvoPfalzKORceFYyZP
a6v6xzz8dLkYIfsv0bmLwhImJm12LEGT18BM+2TjyqSoLEYr7vlOZO96o735M4UQ
yDGGMHL9W64ROcJlI4E6JTRqwhPT7+QJpdkt+k3u+21N0r44tHzQUvY4dUnt6+kD
NFuuq1uD9aRTsGheeWIv11jR4UOf9L4vNW8VQV56H+lk3/UsT/kqpnImis315Zxc
NkwVP2+gsNUknFnyAWQa0QD6BCT8ssn88DOoMOWGJs6lXeXGUEsNiZnrdQt2WQP/
J5sjt3USLIbV0BCHODvFP6vTO5Rc5bZeYYSOWxnO0AMRIS60byX6PQX6Gkuoi+Ef
3GhCqRtuFc0D6wx54Ty7/K6X/lnBAUa/hDwdzvgIFaFoDoIXLu/Dk+kQV+bn2xYV
CLGPMPfclTJqRsJGU48nGxdAMHzSffxfwMbv1hTzXTH0700mKaSzkVCrDwrkG/4E
9XT2FmpCo7QMBO0XDn/O25Hza29BbfN2gMSHQRyLktkjPNrVy3CSXtk+7oGgsZ08
EfcnUgvbkEKm80dGxFFH0U/8fjzme01e6evk/trUuVk/VE+pjjcs3GBKSbyWkcO9
SgJFnchTjA1OhfWNOlgFcPdtWB+a4FtWllre5gIRqb+/BtIE2L3DTpVmw5xV9ruQ
WgwRJJdgE+C8vAzHoek3LmRwMglgTPIW0WEa5hOcOunXEveb5t4I2RLzYGFVvUkK
XbbH4Xu80g6aiCwJ403lejel2rg/qTPOOLxa4e5HAlC7eJ42jjUe5OSX+x1GZiMN
vH/PB9UA5sGmCOqWOOEOuZqQHVJI36l2W1Q7u9bydy5VOtWz8tb8N/r75Hy+ibSg
w4W1Cehmf0SNhVJhtMug1K+W7Aad5yRGhm0B1cT6IHOECI4F9+K6IZms1TZw58S9
X0gNpzvIFPF8EyDZvB1MNHMWVcGgaoKzc9LyJeh5M0SAiW5qUN7PnToi9q37dUDK
BbDIMccxxxLNtn7jeVA+t6sLH8tedrc3xf7XFb9WxzzWXp1uix9wiNH5LeRNgpwX
86++Bejszn5S3Dbh+vHH1ZYQGuaZep17fyC/Y9SHaJdLdKzohPi36QaTJmW0kP2u
Px7NLJG4D9f/x1BnG5kmTnlCuCdXpn1+7nEScHTNpyI7YvJh2amCOEEfKbT174H1
rEOg2AK2dGDLaHZGJR90bjRKGi55k3xpkfE6abh1UDNjd7t2HuToVeQ5x9let9MG
sjjL96HU+0K80Q9a32bCvY51FOkteVEk8GdbGnPHs7fHlYdS25fWlSYQ1BknlbQV
nVWHNIOiSQGmM7FKmfMR1E4bys/5FD/s27aDlGSQv+126/VhPntbJjIiLoAq2qkD
/3OML0iTt9LFKxvpOzr7B4h43h+Mc3bjguIVoDL6hCtzmJ3A3xyc55hRLZJ2/Fu3
99ah1RfmKAPKPERGBMKSXfi06qpHlq4IoJ0QCKWO3zGN5q5fEYlS+D+OhEpvwHpm
ertU+hm4/lDaU1KwS8vyiPQbuP53kkzjrHGBcFLfevNH42hHq6fdHo+1e6lfq6Xa
5xCcJoG+woG9cR5ULdcr6Vy0k/Qf0cL7m/LWm6UPIF50M2HHn42+KJrvbjRRXk0t
P9jvK5pSpFDhQRX0FHA+SnkFK3C+hN6sReRn1cU7gK2F9eFdaXUFJi/XisClkItP
NPv4/IGX4TfOoWZ/QgnC52f1IhVI5Fl4XBzLZGAn7g5VWkdc7wDFhtirliQtBa1j
xQaGPgh3d3W3DH0SNSWqjr5fd21E3MRkAKm1stKHC2bYxTCW0xkHbmA7qvcAfmQi
qNxscxOmPypwrJRmTuMelDUxfDJXX4OyHpjnvac68xpAE6Ee8TgpARIuGjnwElHq
m4wFl1sTRLKyxOpT6BLwjFl8j9cp25Vc57wM0osdYuj/3U0dsSFmlbJYJqogi4qP
+/XuEipVvv41z23peeIOOtQKfsOTnTbb4l86+x5DPKdkN7wQPECwbltdzwxmjdXr
98fu8+JMl3jTRT6J5+tcorrBX7sh2Gn3BOerqGuaRVMKmHw9uCvGnNqDK2p4FSnH
tdatEPKWzE01BGeiewMwbTG/czcFlKFaXmcD0rfCgr5vaTwqbhEuxmVmhHckFCwD
BNdb1hRxjdAr6tUVAtUQHvxzW1oMv3ORwkQrApYFWQ1q3PUozL7JWK4ZoEWWsDBA
Zgmfif1Kx0cBrkDBv5nyW5mUhMKazbf+d1uZb37XZw7Xz8KVBYvzdOHHXvDzhwfS
g3Rn2KT0prc6RTgIjAA2vLTCrw+r2nDetDTMMzjOX55Dqpzv2hy6wd4L88TTva/v
/Xsnmms+psGep2k0QlAaIcr0B8BFrCW3+S1HndwKaLFo8WYMlfKlvm/XUdwi65mE
JAytiImvTMkDGvmH9JyC1xCpZOsq7bPHfhftzG/MllKvKnbM1LsQv7PjWrmrUPTV
onlsrqliQgsRBZicDaVukZ7NqHviSJovLebGgQEcjoXg5XNQutj5b3IkQDigAV0m
CF4mta9/S+tJdwAYEW0M3dWqiGm0wogJbcbE66DgDkVdAdANm16OMxE0635JruDV
Rptph8KI+lOH79PtKni5aqPVeO/nahbVkZxuTo3BD634BU6MzIpJt3UWmOFO/AiN
k3QjZ5fkRUAGzM3AScfwVnwIP+GPjP2RJ/6eVtRhcrv0F0xJCrxyvkU0E5tC51Xn
c8AkyL/7dBKWtQyo+aq3pb9YGsq1tTwDLZvwSTicGjCWsvtqTMx7Qjy6R/4xGfCz
WSIEMD0s4aW9HDPoakmOk2xIc14UIqX6+Yp4uLfM5tUZY60i8KlRqc9QqUJLW1G5
DLiDf5Qk2j0c2t10chJhcqjpMwvH6+ARThT1rLPKxsOQ4/34omcCFKWkULYJQ2bJ
6pcFF43HNQYGQ75+CBR/iCHaPFJFVtug7zCmO71uL9Zzp1NTay1L6ymXuRM1QPb3
ozNEjJFfRjt14oGqLemdQqxpaAPGhishkJLFFrkoY1q5AMqS4MJPCTjZMM7XvXPC
BzdA64Ac4wyk9pPtMlsuK+KRRf1f7uHya4V582QAgvCRgAg+m/MF5vVt/8WR06F4
8KbXt0RuzWikg2z5eRiHs81dO2XYG/pa28OYPNuVomGXmCNFvHklQoyrwYLEyLbG
n/2N0oUXdgmvPo7iwaW+2pzqgWjB1z0j5Q2o8X6weO2bSOEngfj39cFkICUM2/GA
ZUxcXP430eLpOHgh4loCyeFM2JgnzlFcDJHWSBg8jOPYs73ph72Ciu80goRA2JKl
soBTg/QKRZOA5T62IpbQ6BTGa0ljH3TlC/GKPeila1mKtlQOwjGGRVjzoh8gEpYX
K0GxH4YMHnlnbfnAj1bP+B0+XDHwtoGyBgZPjxu7Hp5UogEqm/fCln5WeAlLx7TE
wS+q2tFpeyQVI2KhkWylFtWwM6fMhOFH2F11GOEuEfk9MMVIR2Ir1qzdMvkUPHtE
DRI7OmdOZSiyAJulyhOD47OvnuvFdes4r4FMqpDTXqZzBLuEuO29hMP3jXdrrEAr
NTuyWNtn+asydo4G6PW0WWLa1C+fd6hOck/4mTVjpYwbM52Btce2dDK4pi6VQHFL
s67hIvUO+W+COVLcDIBuSzqmz2rqJF3i7MBFD2cx1yIB/01CINbdmNYfgUKwxtTX
+jH9Vr4US3q4mQUAslqxLVg8wtTQbBbuOU/sSbsQO96UgfnrZtArog07+8r2LiMe
jL0Gg7Jgbiy73BP3wC/bA11jhwkJz4sYPDgBLH06dPN7duc/dCALgt68K2kl7YNi
aJyuV8R9fvxhUIduJjGb5zX12xcOUNCo5r8DfTSo2JKT0ys9TL8exzJTcVXk8cqZ
Zwk9gZqSQlg+Wgm/uUji+K3WiLX8Rm2aJVyDisw7HVuVWmT3iR6TIuJ7gNLNNmJr
dmgz0zhxZN4ojg8l692cp3JwndW17CrSHn6/E7d5GSIm0P8amvkBzpjTre54QCvk
uafM503Ks/NH8Tg0dXyJ924GK5xoD0QchdZl0D0vza+HZn1MTme/ECPybofYeAb2
7ZfajeI/OhxelO3ODkuG3uo5JLwA91drHGFUR8H/yqW0iLy92jxf5maGicvl5pGI
2scnmvAH3CwTZ2ROhmhLmA4MKVXN9cEuaxKgXMUjGgKba7wC0h7hrADbIk+5Wzmr
i5CYqBD6NXas52MGUwTVq+jOOPCEDQ2LE9feAkuqKoOrSg/zW5Hnmhkuso3Mk3ji
qBD9XGJVnwlKBjRPCBoD+g==
`protect END_PROTECTED