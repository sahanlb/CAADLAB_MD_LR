-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
hAx7c7Nqx+5t8Cffeqcb5ftRgmxbQkRX18NWFhSOh854k5p0i/wJxlJMii5yNJ6i
1mi33/jltQ/HvaESP7f2mJWNq92mUr3Oq1bczd9RXh9BV2ezEvFylgjaxa3btytZ
HUeXQk4rvFCN3X7XoMl5Jv/umI1AAH+o5XQbtPnQse4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 4304)
`protect data_block
KifA06dyjx8higL9wCRfMlTxfyVLalVczANfCSZNBWRLXYxvu7YQ0EbJEBhglZKr
IwKe5i+walnI5v4R5Xt1vJKzoT5dM3wb+Xpde4EFO522EdydkgEzG4IrJeqDGKK5
5OHvO9x2IKyJplnWRDj6kFGgGgqfZEjT0AcVw9E4jGnkJb9rkg6erIcYFn8ppnsD
eldCxY+UpMlTGu7qvoz5g6ZeiafXF2jZS+6bI99nJOnLzB6E75vxW3zMW7Wk94H/
51sM2iA7tjNKFPzBAVtb4Zt431NiHVDWDClQ4zgCbOBdXSl+QzHsJs+NH4WVfj+d
3kc63ETp+1wA1JuvDyTlljgEDCKwDAuR8Bia6GGL4ubpHlHMj/38N2m2dSpG1aoK
IwEmkfJukv1dzs016OEaN0g0qD4APB+9bc1XLmov54dOp8eahUXvoFa8PCxokot6
TrqotnKBcaPKS5EKgDPU1P/la4T9nSY0efPz0q2iCleZwJ0UCx5XfhB/VibOR14K
dbmnbonToeCWyQcUr83S5Dqp6utgWle8TbpqQmWFre76wKP4w8e57/QKO6TBdr49
qVSLBuBi0ZjWN8rrOtxuN01GUTIKt0Qb6pLuZZispXjtrYs7uYHyL8ZlwJECF0lU
rpf+H5Wyz98WiJ3D0wthujDd5iU/bfYPeJ6fbPOcKdRYd+j+C+bR7RzzQm5JKE1g
swb4aX/sIPHVyaKDK62k6wAHvwAj3zTBMn9UJ3mXEfCeLhTSAez6LxSnqoTnA+dC
kYIhN5uPYsKf2CK9W6g5XXcKa3UaTnhceYw5PiGgs43GwtbbX4s2HTB9DK0S+2R0
7Uqv1rSvAmYXitV2E/9fvyyracU3dq15T7yc+OIinbb6YEWHIeEqwLGSOTA1DGNL
ByvA4mxPmiCDmUST8mQfe6Jegcl1rsMQA93Rg2N8oD/C0Chz2HdPFB4wJI0UVKOy
0V46+NTXhwe5P0mrfwooOomt83Z8d8u8T+rVVjK1T1wHRnw8gXgoGcWWxs6konZf
lwCNpoTtcE0IQT59Tq4Rk2DP+U0W4GLf6l8WC7rgloOfQqQ+NPYgHwmoQEyVYdkn
62b7v4aT4h9yaRYz+WoMeXBfcPWkozOOQxyuPd7GHDtX9069W2FXQ41a5kLp915d
s6Gu0s6ImlUupSWSJUiWjPXmTDjYauBRDLchEUWjuGXvB5Lz3q7EcpUQ51RGogvn
76RTS7fqhZ03PVbdktQjTdLvugEviEgFYN7sdyfnoIhHEYECRSAbPNS+gAPXN4NE
AGLiwfrlUroh23Yuzc2wYOz1I/Q76FV3yysbDawUKpx53wWkPBQmAi14b9012RIU
sZOMm8vW8YTTPjqUjjd7JZRNCJJei1x9AQGD0tRAMoQ//Hk+ie+FzVHEY34On/SS
6hiXr5irYepDc+PDjUiTq83a8BQECEg5wLbz2a2W1pRF3BEEeAJJE7wTRks3JcHW
NmNHB+k4dFMZeWSEQmq3gl+LrtHKQAhIRhFnEgIPgmFNPERtkWMJe8+GPXNWs+V+
lYmVSDdRXTGzdjj1sZxMA8Uv+9zFrEGIcYL1FknLBI/rppgOQPCc89KR2oxDjppT
44TGdT19JkET0Tzuv6WuLgt+MzmcdxEcMEETSsvAsusZ4r8QKlo7g1Z3HzkOc1cH
d//KXlfVhwhWR9JbumVY/z99G3AGcoc1y24cncWkp3Di4mnOhNoKBIa26XImjHQT
GLce23eAeg19WgPAYYc7tzAg1RxsXumcluTAAmw51FJSmR1UaI3xzy82BnHaUYZy
o5RPOL+izmipLbCu2gSt8ngiZJ21iVCbxSVvgc/L0dZR0YystUJi43zpG2gPBBK8
fWDThmwgkvcx0u4k9g/eU75GAPSSHzJukH1Kcgq8jHcIhdYJ1axI+J6xIbW90bA6
xIFdi3j12M5VDQi9Y5yHciTdfry0VKt3uSNfhl+hYzXX+KrZVpayx6QnNNndO5Hw
5YDcfcRpx7t6TdfCPzQPY95nnHUHQh5SoklsPPRvgfZGY1Np9rQV2dOzKVYZAMZi
c6G3UMQUj0SfWG4YCj6j/mt2RPeCCFBTOTZDOE3zNfKA/KHJp4oJ7RFTFGz03Evj
q39kh9jzs2uBu5ew4wKLTDU6LaDC6oNRRwbxa46awNtAU+XOKYuenAX2X0oChh8U
khMB43fUDbc0E4bgS6oRJ9jbt2HdyH8dinPEGNs4nmr7s6ZVlJ9r3p1BVlJSaZkH
qkHAxxjZUsN6MQWsN5TSt/+KVWzgM3X2ZHM6TNwV6U70GadP63xlXgPWh0o1Tleg
+AG8SRbzimtN68Wsg8CxDLAE0mWywd4/FV/yJ8TS0KU6BR0P3wfchuG/K2BwK4F9
kDRQAYnHq00QWxrdKstHRIziT0A3zV1CdR68wb4KUPhvGToWH3D2uMphas8y4ETl
LacTFnBG0PKUCXr5wVQVSY14hClK43q+qrivZA+QkgUMdGGsNMRQBE8KyXKfSLYI
Htj/J5tJj5Z/VMBIF7rargKw1qLTSIal6ypCn6Td9Xsa1sdXW9Y+vuE3ujgWb0bz
UhdFmY3KD6+AHUUfmY0D6T+CotSPHxeQ9I1927GdhgR4i/WDGuZfL3bgZx0eMEtx
A8J4tKjK5u0f7V8461wc+MryKcvu9thiwodDZsQsPrH4jbxJeCX8v2xITQah9lhh
q5iZqa2E0GoY1shfiIGxspD9aTq6qWwSx6wUAvc5Ldoe3KQWEvcAf+PuZjeO+KYt
QbtQ3X7lGha1u5UsQS1ASjDGUb1op6sVCpwLl60lZ7t9JZb3ONkIvM/lWP4SWde6
1pSRMl+tYe4tS20OXhOq4tesjB0sVDvbTa6PYyU1iopguvM01RFqZuQbBA6r0hIK
/1DazG8tD9FJBoVi1uXKY26pKgAjTcj996DzWe+6pJnxMOvbdSnnxaVpfcTS9RZb
r3NQfjSIU57Ax4Gugw2Bc8GTLl/O2BvHfTsQnHUJPlGMZSzV1E8L8dvqkpqkwI+h
vRMlN1Ghj3GVjiIBhSGgOhHwHM+w2LSaHP+iA5x5plkw9p3x66BNgzZ8colCkSLq
pV1hU8snJlYwSkkckq+Dv02RwgFEpqIe+buifDTBJVDT8fC4yVgHuN2pC9dJg1SD
aN97M1a7y9kIELcv4TCIHe76BZCgqWe0I1wHQ77Yiq/I7NreELisc05qctD7eTKk
pz+oIeOTAqnBGfKbqc1bWd+PojxhCwi72vD+kaE0Dlyv3eI9H24zwEfnr6dQ4n5B
4Ywc+yOo417sOFYrNUOElynUWIHypc4LAYKbPyYm8qTeVOuXNQCXAuYw/Y9YfkN6
axRgXZSmM9KserVj2WeOoV5Ijia4tQRrnybE0+oMQezJ8cpiVNCFUxsvAuXKLTPw
NGhZgsXyFDvWU1h9utODBfRIimKc2Lrw2EmggAVx9+rfDwCwLTFNUxM3Bx0prHOc
vmMuB7pNRqjIU3G4C4XR6W7kI51Y9dnGAI3qQOH23O0V9KUSJQWVwS6+BsR0BTwL
82jIroEtJNUYYsXeRjYuS8748Z/9mgjCdexPEUFEQcir/lo0flJ3Ec8005fRg52P
DnVYhzLOGssHq4juJ7jHlLeJsCQm04oEvC75yX6X+A2oPPQDhl/TZVVxFK4jatzU
dobGV31eMl+SNods0oRi97d3NDXs1S/9x3JVJJAhnFimFHjJv382KSuKyo7fcRAD
sZ7vSF7UyWo5pawAbfqa0v5VWxAdZyTmJrduAFhy2zDu1VlqbL55HXk3nI8Y+ljo
c2fX2QDRoqJQfxoCbL5yiXDF73KIZQSPOXaV8L7VgGf7zXdD51Pz1WwNjIQKinrQ
HGXU9tRZTJn9K41nYL/DJ3rRVtjVcs2DM8Jc7JNSkdCeKs83QxRSHMBjHqZOmX8k
s7qsogIq589YXhF5wW0nmSHG2DrNJk5E+girHBFCbE4mQAofiAmGM6uAJFuJRYAf
mMhdGP1nDX4NHO6AFnB2PuCXoqJw7Bm7+hFHRHc3Ldoo2bg69fJQM1wuA+ecooGl
SwGUnXsmVnuqZoc/nqeX5oMuUJyMbweQA/4VOvg3/6G+OwCE5jbcUVGef+ZuzZUb
3ZNngAeuC/UPrXJwMmGKvEMPtYBl6x8mn/8tRja90BsOLga7U1svU2G7QZ7zWfeh
IkC1j1WYqnZ39bY2skHZextiuBSIiAQlxDDpmS6na4cCrYuy4C+QpBQi8h4G/IqT
ydJf7yB9wXUw0NRr+R1QSTVn7/LpU76pD8xnux5zxoCYJIPtTVmr0wR27BNWXm/d
vBxm07TO3XbItdA1uqXPr9KKGqELzg69LI3HSrhXSVImedqeciynZSVnNO7PRai1
JHDgilotB4A3SCGfkA6EEIHvV44gDERc1WltrOkGYdadAHjlDAEnPXsS3zpkSAJD
jbuUGqwU3SCucPcy86oNHI+vj9Eontee5NvuH3aOCPDvwxIVXzxf/iwTCIb7VlNQ
MgP1lLACe5VWQZfMv/NPaXQehr2gsByfm7fVjy2NaVLyNpY7KJiEgAP9L3KjioWl
LYAv/APY3rsq3Kg7tx5eGrtJ9xPTs3Ga5Ra3YB0uS9AwRxe4ySbg58Gktkg7A0U4
pklIDQVJdTeA7ke3dEWHLwRyLPz0bjIJ62OEQYI76+gCX9h9Dw99Cy/OHtmC/667
UQy58wQ97SX5s8krU94sNB7pmK9ZuaW9DmfFpcXQj/JwrLgVSyMjPmR1sXX59tZI
wyTcU8wTj/nv85CmZrDxnbHI5z1vVGreXYvXa/zGPQaqDZoen5gI0rFIgC+KSGlr
Vz9SrtCgwyb1gPPv2rx1lvgLZ7jd6G/e7aVCdC5+9rPm6/cMrsT8flYN4WWaHkLf
vUWAxY05Htik5ZgoPP0R2JiKbZ9XXgALOAGKEKAAEfs7aeVVk5Y1+S5G+Ai8RlpA
UlapIvooQX2KeT1qKXgMY9Jckj67FfIBer4bhabz01NNHPgiM6r/X4Yy4RO2A0iw
wCYT7TRzRe9V3NyPv9Ff7iw4o/mP4uhQO+27ZAUlA8tG3U6z7CdXlxEKdr+REtPg
uerdS0nMITMXK4wVAbEbm1be5skHlz5V+nETESEE1cJ683CFBWUM4CazHAqPc0wG
1ENWg0UdK01JswrA1akVg97i9X+za0LrvZEsT8R1xZo6Znkr9xF4f0S7yLzP1gvt
iY+RgbQSqCXSYU+idLIMORSqpzycODSoD/5ORynDkCvetIB1wJKfGyeBFOsCy6t7
APXS79MvbHhx/x5hZ6d87gASYIgb/VGQedSxcZyNEfuhVnvmReuuB7LMK2AJ/Xhd
+eLV+lXySAbqhLvS9OgXhz5VxNJ3cCDCKK2ahW0NXTyXlACAjhQzglHeexcWo+3M
J2NJJuuORojeozvoOQ6rltZLV5Jq8qvnyk9rcjDM/gbcRRXKCOhHxIDffj/rto5m
D7jEDDdB+HcJLUgrZuGbE6B2r0/FpSbCbuq+b1ON3l2qxH4zu0xUw3UIaGHnnnrA
7s8Oz2f1N7qxE9ORx51Es/MuTh7Sp8tDgnSxwy8l7OgXWC3YQ8C9eoK0g+g/7WR6
OFuQ/RoDasYWwdMoMbGPzGtXpbuWhOuhDPnbRibaZPOWxXZwAsC5hZklxz+D9bc8
N024GovJGiSps7N5NeWZd/8fSBMEhGJAgIXAPw1Kl6o8zQ3usFyG9YGcirsbEoh+
yogz4RI44hXtcybIFyHEffbRPQQXDV9kglimLVKH/dQ=
`protect end_protected
