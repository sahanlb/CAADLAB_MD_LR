-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
QyWFYmXDq52dtdRBYlHaIYVBVTb/dxCXZpqLlW357rhwmvE37ziIsU/RDS5mMRqM
mWa3qk3a+02WbFuQop/PRA8a35KuR2WoxYzvTIV5npuwUqhAa2y9D5A1GrFcll7/
XNk419qVhZxSfKbHYVCK1FN9JEoH6dq3RkKZDg8Acf0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 36304)

`protect DATA_BLOCK
id8OCXJ0Zsm3A18fCPDEPxkex8AcsKB5gtBBobM5Zu8nkVbOTxgGEgw/Cx3TLXDi
0wPnuuNU6xtHfcOk6OfNlAybO/3U/rvD6I+Gfk0cziSoSPPKhpZJ3sctjJy1QBMz
Fm8QYvan9SMa5KrjESVCtxaHVdIR2bRjcxZWGkagEpsvdkVfljFUbNoXNWJAk1NI
Dmwy+sy10t9JCN/iUKT5Ccj3o36yjsnewgBpP3Juxx1OTQOfoxIQegN4fH/dwxPM
hLwhbr0B/OcbxmyjJyhNB6u1srUJQkSuM7wpbB9esbCqu0Z7m/Pn4jWEjjO23SBN
U4S+4SjtNT6vX+9igYt3LWLeuCXA2SJzn8i4pcg3LJSl9vNmvHNlfJuScIbNLF5D
VnhbN8iWD54O9/978hO+m7s/ohzIfGvQWjAbTs00EL+bBqC0Rfcfk7zlVc3OPeAp
jflw56CtT21xDh9owJcRLq9+yUarJNdnuqRoFe4tY/UIif4kmpKoJnLgK7gY0J8H
vz1WjjSL1tmg6eWVjtaj9OiE1h6MpwZTcpFY/jR2S2zwOgJbc0/tLVBIa+8q9juS
vr83RJ6UZskmxvVYcpL9D7fbNji/EwqXyJhesuETRGug2c6MMF2BkqsEib0Etgzw
LsTPcFDBxhkGFBecPoMJrFLI5Sb1GiciyYn3KRNF+IFVoeTCYwdSdMtO6pusX8DC
f+RYThKeFs1n5e+K0FNPNlUiRkjVGi2IUh+i4CLfo8RsEaYEqSF8j1cbJj6aEHW8
hIFBPiPfrOhLfsdkGgkNn8tTxp+nZyBxd9kP8sf0dEoYY98fkpO4ioi4mHKfUc9/
j2uKRE2mQv0lKHjTFWkLNwBFBy88JAfKMWmtkAB3gSqsdbDHQlIgETkV8+Cmudrz
z0Q9MjjMn0esttq0rUqqZAzbgb0rWFCsbCi6GShRwgZlgcudnqBKSrwmynfWaKYv
gftsanNs0n/arxhwYnkj5PiPF1rhCwvNKUECZKzQ17I7ZuatshIZyAVjS6cd/JyC
zx2vsB9JR8KfAyOSrZdKm609p9mGSBqBULMDnkr9LJZE2kgRBLdqHoHiJRa7d61B
C0ao5e2S6PnusA1mqp1c8GH/7j78dZYpL5HRDtgjrdrdjsoz51JuYoQLSoH5MFxB
A6AmBxw72NJ4fJT8G74UUn4Ly20n6fOtiarMzDI2Iq0UZ5guOwnGetD7n9uWgM9E
lNmFgl/kqqre38mKPw4zEZxVt4dqRClp3di8H4aV0bFYfcorJTdDNbs5M+njN2gV
2n09pxTPiaeM9t7oi67vULXhioahMywTQcmeyZVRu0tIBYMTUdgas/3YSuRKclly
3ir62agHNwDQY38UdAvKY4gWWJxwon3dfanJvfLVVT2+KU5iLubxlxy2GzqzCumU
7+12BWCYg7z1Wj7k5TqnPBHBKlNdg4R+TqRlp7djGPq6c+ZzfUPcfHiUouBLZ5SA
xXaKdZdAfZ3zYTYzAHtSUn20119i48veltVwtbDkzHlu8CK9GKWvoBqYgFBn7SN2
xWWHKpgJCyFEBYo0f3axfmb0uINE34PdWtIdEGEYEPRVRZ0gXAwGHzaBXzGpLFPq
/tcRssAOi81aZre5BjemKZKILMP1uqo1n1kqTw3Kl7xL/F98dixV5oCwdP1p18VG
UFzWoC6HtTIM3MGQK1dqQcXIAyyTb/2LoVFVEnLL3MtVfln7Y+xnYdHm6rF6kcXS
MbaC7jVIL3zcMe37lKMgkTEeRFQyyG5+mMX71U42QT9ZuPh1pvXAbNZbk0EW7fSY
x1r4y4z6JGBijAQGms5x14Ky73/T5nA7DJPQtvY4QNhwpgRmCA09Gvd+a1HbG0Cy
cMdYXSQ3RPoFYJexwemmYmzJ2xVbu6Pr3W5Y/GloFOC9dddg+8XYzFA5WT6lPWiq
cRXIfoGYcy/e2thDblvg0qbHul+BCXTAGvbfOcuzRF4Unb3D2/0iUwWwK1XOq/dM
evLyVb8iNcnIaR7Eb+Q6RXKwlblRTUvedHLNEGdeYe1ksVfvq1YRCMKOT6Oyq2ND
f8ddyGC+2HL6IARzU24Y/FqlOkmovpORHrAwxrANi1aQpFNkiq7WPkP7lcrW3wxA
RF2LhjR8u+SWV7OFG+CDjzmStFEp5RXxYJfpihV+XEYRRSfH/Padb5zTn1jYto3z
l/rIo5YS4pH0AEbSYpfZOOsoT2CtxZzGjRF0O/Lg2EHhJ/Ffe0xuW/p1dFGIzkkL
3P9f+xEfiQbUat7mvXfxyCInJvjGblXLD0OjznZQzVwtgpsiUbdkZyCYP2/raCaO
EZyR7IBMAZ7J1/qgtr0YKBSjt1U4CPSmJQ+9q+71mw4Kf3yOF70EWXuZcUFLcHNX
CVELiaiio97OR/ywDll68OJq9TYP3HA5J4c+ZUQ+IkLsByeWvteitfI2M5U3uH5U
l1zb5tAi+AaxnFE1kP7J96Nh42BA9NN/kPbuSUItUA2jpcYG9/FkT7g4UgARtkJN
hf5tDjjxJrS5S6VDXVf6Emm8pGBzfp2CipcrACwKZiiyFG+05f6TXLoDs3wByRCA
LG/FHihwfNXcVgCFN/jS91N+PXM8zrsEt2FIOPwmvhM2g6iuaZ873FDs7uinVTMi
S/llMbtAWCl7vt6bkgRkTXYet+06j6pPjicUFjl+Ahdlnxf33GqZrOK51BxGoZ9L
FcV0jqCKwrGQRhowQuDhLpChnpM5bMOqOTYi0WysirMOEzGzLmkERLcOok8baGyc
d+6miQs3BjH0vj8lq+IbvNtchmQ8t2TmyM082EV8imDz4nIjtDw6lZ8EQHfge7Hl
k+cmxFpYPK/ygfVAD21/jwjmXcGHk1ZOsNoSWijoKFhwZappZAkbEy4qDF480yAn
ErOp0CzjK3I52gpNZ2YPP9NPuGEVDpO0cDpNV6xufbEkT6/vJQ/QK9E6a6v+EJRz
QiAHy49XpjKkjeCQw7baZ6eX7O2MihqGgYA4hJXzQjxxlTfdmA7a0kcQJn+94Rsy
m/CDgZRtTuWukm1PeTUCDQyP95ID8VEfbtMJSs6WKgq0FT2RKtlSoRVWDhMV4et8
XgJY9KlvJ2pWOf7QwamsnlE6WqNlsnBghvh8Yw3IIsc3121CqDkwficwBE9yDC5s
JWnsNmtZ/1699yO0ptpcO2S4F3AHT8AZdA7nE1XhIckt2MFlG5wsZYgR9PckgIhe
Y3ZmnrfMTlxXhxUIx7mMQTZ3O5W3my+3rUWReTZvYt0VrS0YJcqMlQ7H6Jf9qR67
whlIOhQEFM/0CS8FI7u++2Pqk7PFsJCyeEgy7SaJbVXpHpp94HBtlMGV1Af7KIKK
wknm+TX6PSDyoH+An1n14cxRcHKmALhnIqFfRAymXi6LG+VW0EmhF4OA8SPZCX8o
1L/3pAkNpOipmRD9jKiIR6aUIeGnRj0cH/l0O3puCxc2roJwevCjFOIo/xJV+yfJ
89rnMrBHQnmDzoqSj3kpiEvjxQRwHpixZZI801OnlxeMDKK6Xjdt0//eHjExWNzX
bENJfDJcYvIuA1t0W7X3FxgzLuM+MLySPrIqZRS8LfVevXgGQPRXhheOwDlh6J7n
PTAmD+E71QaUXZs6thuTdFyc9FszwlNK0sYpJp9P5pigYcDQMdEwGHoCbtcG2xD3
19dOwatzqjrnIEYbIZnS9fzeHsYLFvESVZdlzTgNx0hF0JKP35HT5jZaQUVOHdSU
SrMjkBBJ4CMPk2q+xeVDeW/nLHuCP0SG7lpmWUiJwMn25BkuPLf5E7PagawMr89j
INgah/T82JkOsY6Bvi59Ykc6XCnEmsRn5IVCndT8FIFhMmzGxGRb9lKiMX+ERWbM
YpTUy033q9FY8WI8WY4pJ5u7JSGYVi1LT7VUcGVEtVPhJYuJ0aEqhxs04tptKPMw
3FFv0cqOWXYzvJj6xdCGfqRSk28LO/q5AT32BfkPPdQaF0mYmEeVjBDpotiBOLby
RPI509vYlT/e7MHfp7h10KixZ2ac4PY4m+Z6FwJjGpbO+RoAVfOU62+NZ/iGlAAc
emwZlowHS8f2F+VKE2EDrai2vNUvgGFjBeJdb6eUiWIPyXKRDsb4rfhO/cz5lt+c
iz0VRvaAhxX7xOCmkWog6AhpUFrkcjKTVjxkyQGL9VR4dwczz6eayE8cnZBW42Ru
32FK0uENMoWY0C1SS+qveGnLMQHwGrk8M4ShjSr5846mlNFHnTJWLBf1664J0j4+
0sE4odC5WbEwbPXSjksGEKIFWgh+w4dCKD/f1k9twnfHCPv+wB7+IUzZ53LjRRw/
YSypS5LrrZKC9x9IwyMA5FZxeqUwV6JumGu2lRAFXsxNxYqziBf/0ku9/wSuEWWv
iEFbPBLgseQJdWhYksl+YvaPd/O+l2UOXZvuUDq0LnhtiaNlD5jB9jaxXvxPwn4x
QVMymaZpqL4pe78jm0Pobhz4wRN1fB2QnsUBU4otMerB/x6CF2mgk/Aov6xVV9uA
Ywscr8lIXDfO8diaS2kJWcuoIzm0SJNDaNmQc8RN7V9I7ojpyTSER/gpi3ImOQcr
4uwJiGzHCScCcbawHJopOiUD6EMR9HDArrDkxUs1yXYIqDfTp1P68DYYXWAQ2YyC
cfFio/TGx0tTNwcXuD1XKKzqpMoH+PpWmvYrXVdPrVVuIgtCHBnwq9CxrOupGF4z
O8OgDWqNmKhTC1Cwknw5MkOInr6bedqfyvwDTQYYCEXjZSLgMh9X+lLmnX45O7CM
4jZ/pwRj7nY3ymZOnKidccTOY1iH+nH3vdoqi+bLSqVvwsRnWpef5lro2IEelyQe
PBgUYxRxhWEIUS3Nnzs5apeGZjn8Z0MoSRhNymL9seIVHWnYIzINRTSf8/yVOteW
XAR6128FvObIlzVA2vGpWzHF+ZBcPMm1KVT8olZ2aQO/1kcptE+S77EcGG0XmUI3
teml80noZbUyL55CR4AsmcFWOTh9y+ZXQF9fpgvofmAz2Wz1ML0oNI9cm2kLZt3/
bbyMUazj+kkhbMaV6Ovxx1VmZT9KLsVFOFOVRzcuDlL42NQkHc3heQlwrkKQA+lV
HRMmfpKi/1Q6/q1FaTEoAtfT6UNkEL3cyA6XEhQq1CqGH0YQe447u7qThmTAw/7B
6idOSQyVd6ANbr7GXQWsraQ/CnXjGkKyC2n02nA/aeZbN7FrRziUS3eawD5BZmr+
htE/2lI/y/a09g+7W7FUPeqOBGsNOS1cT0qZVAuaxPepSs3fpc9Wn8uRFM4vBmPi
HBzmXAiNGN2HOy9jlph7XQ84iCP6s/+gz5RQ9GneKuUUdbvbzMV6tRZBNA1+IwRN
EBjw9yG/eX0xK+xSfUqmSCnRawjuEjXCYQw66vehhJCpy+nk6PpE+y2wtFu8Dkyr
/kE29Esy7SOPitfSylctCSgiu0yEEDMWB/a1HD+8FUpIh/qWZPxg6y9UELrp4zY9
vczZzh7QRcRWPgGAsAgFezFyqddfYClJW/8C6Nk8jGbmAo8tPjFfSqfKW/KkTkJZ
E1CHDZ/7o240gog1WNOnuOQsxw1Ytx/h61vG4fUVG/8lK8Xhhm9dDoSo2yRyvbWO
KKizBJWi1bffAqRJnUud5VuIbHbcQxyRp92ECnNtOEdesXIsd0QEukiphSQJvxDG
LrmtDzPW3I8jNXSeZxHy/E/U+xsoSesidUZPYsgJaFn3SiVYICE6B2fki/7tYJKA
m5BpFU0urqvgW70tzAHBW4Tc78im9CcZ3Phyqyn9aP/zMsgxZTe9qdYAe8OsSgp4
gUTeFe6wTTETOr2MlzgHwBYThpu0lBmie6spWhx2ZdafNfFiBm0tTbFkyuhJcld7
98Ixa9wFYxhlGbf8tuIayRhyBZN/rVNW7fkqwOQeGbr3/OfP6JoWqzKIvi1Zg0am
sHxe6QYhjA1vhicvcHoEMA1vkEiZgOykew9cDkBxYYsZdsD/SrGpFv/qoknp6T7U
nEA1/cAqBWzeTtGTrABmCjW1MRfVZg9cxxNR8Q2inwsfvvoHAuRgBuU7EhdPcmYI
MrRN3NINrDklvsQeFvCbJiQEVfQHtng/4XWsS0qs/kbo/CrXrSXzvjpbqVb8LrKE
73OarrdA5IauFcoYkhBYHs20rrAlyw8v984aGkRTAsIbGwFPx83yJEHqDr1P5RG4
MQvToYhdqnS51+N73Rt0wALWTiFFzgHKjotwCHK6NYoBrBXWbyBK5qzexaiHvejX
8nwyXvBYK+TMQZF7eJ2ygEpCJe9r3nLO+1WPn3TzBaMS17wQs4wfMOsuNIib1p93
f6yAWDc+0M5VIgorjikUL9kJPAxoxhChpa1vFR1wz7Lcn9lzwo2HKx192aQUKa8K
QbQDTtziOfR0gaJ/eippOcU4CpDb3PAZLKP8hB4spueiurID3oq4ds0EcaJxIv91
Cs9jbkT7GWfFXUeXGu3fvaM4j8mbf/elErTVnIfIjFtqoYCkzs2yVtwLBtMJIl72
GJRyyWVEfIGu/ISclDJDOpSBWWmpy3u7+j01/UMEBtVlRy3oSzNF6iyeCBwCXQ2p
mPx9WnMEQKKSYrAxR/8T7AUEqOhY5h806mtwclI+gblTrrpgiv9TAtIv83fu7s6f
QWXkcB6aORiQ3F4aoEeqWfGQOr+4VDkAtsqTk655JUOflS0Jq8gzRORA+Nvb7RtV
L4qOzB4TO18W13avAkcSSDg6k7SBplJGXkKPIzmcQAlISrtFydv2uTzLSIMfLHsP
SSpxhRTXUjr64shjXH29TKnNWoz6kesHo1k46UgpgSoeP7PCvZlWu7gnETg8QFUV
pKSGhvd/gbg9RE/AjvWixQnvbIr6goHyDbk76isfLmu4kLZ4pTy3uWLk5b9xN4vk
zB3BqqDhfDIYPQF14DP5IbWRXWhR+fcK5ySy5simox8FZ0f/Lfq1QWhd3+wDJYam
IHNt7i0x6w2xA/nUIToyXUu/DZpTyJPz+u/D6uRGbqic22+iVCENmv2aVzMQK1x7
rMb5FHACbqAGzCE9LfdPr8BGzP2aVKFy9PKs8XvzCnDi6RkZYWeEROYK77duSawM
sDatcm6wJlRMsWcopwbuNMR1cXIwxIGMTdMbUJ33BBaVJQ6J3AEFcoC3iBHaIErs
eobKIbIJZeFRxncTf/4jAfnvo3r3mtoipm3vONfcj90tVJB2ypQbsY4jBQpjKvEf
uJ6DJrHBtu+Elo1NHQkd8AlUIsDqez4fqDXmfUpwrIvicKtofACkMQABSWUUsPWl
kM7b6wTt4pTA1bHYM765fVqqI+yBGG0nzXoFwprjfqTdtD/ZVArsbv4vd6PnxghP
3OinVl5kZgFy99YPBBQMIO6m+G2WokBMMXCWmUg/gxcqnsbsj9zimkMA7LG0pFHv
zF0uR2e1Pgq8mI5Ho1NBTMbRSB5bJq7yvvY5k25Hq2Ivd6Shr1rwoa0r71lPrQH5
kkdX0omCcpinXUDd/WW3gudoXLkcoi+F7HFk9qDWRQOmHUkxuFvB2cpxPqZ6ERpx
C2W9056CEZF+LbD8BHKjrd/ZLv7fCcNsod1FbjCBj2Q3rBjkTC1dvakc9mgKiYko
YE+dXyHfXqZRbWxAIiGjVN916S/l+N+lHsy6GDA1lA4gliUglFj4N0+TpawILqoI
Q0Oe+TwrOg64bw2ugITtlup5EDKWWXol06v202xLmy5/nfrB85rUtFn70bNVL2jp
TFD8HTL89kN7i9JBAkpPxoeihM8TSEHsKqeliyOPfUHxIZ0ewvE+w6QNLFRdlevo
rSMDuViYXgpQK5ZQOIYvfsEqpyhz3aA/ve/yyt6smKsNrIk3QqoKSmACJ8ylV68b
mzBayXjQ+/fxNkvLhc/SYgiMGOxXR+kTFom+v4RDGb0md7f7e0VTYSo1Xb68oxbN
BSVPCG9pEhSO2nBkAEhXSLIG6zXzmRB+xkBC2qciJTtWEXmWiOmgoDo1sdUREMBu
QL1NqjXZm2LMnB7VpMoeIz4xGEzvel0Sobhv8wqSfoDy3YhqTqjYaqvsWzGflJ+X
RzIbADqVvuWdzzxyBMGtWSoa08s8U41nYXfPx99rMItPfq9B5dXARqkdlhC88KGi
HXIlzIvwtpcjCmgQl9evm0sfI3S8WUPlc2Cs3Btitv13BhJe+RMaeS0JI0ydhjNs
ZxsY+8aisgwGWcpuxO3gtbJ3mJQ8vQw0DJ15psjRfBQVRKZJ2yc0l1R3jRyDogVo
O+hKP2ciVGdAD5j6FL45UtxTJ++lVA6B7aPNJbVkEQoljShO7adURa/p98ubguXR
tv14I3vhY3/VrlMP/hk1KsSwryMPOtokFpfu0wZePSezRJFwMhJ3Z8ajDKnGNA8W
moCuAJmofKKaxAHiLlHDlMfDzNjBX3dZdHEpPr+miPT/Mf+xwXHv5RAR8SkPSQpL
HyKOl1y3UfuC4GPgCZ+nD3Vc6H+T3XZXICaVImFe13CGTfbCN4lazLsBDiczTYax
J6zQXdVdyxR7zPfm1DvxXsQwJt3aLJDoQSTHmLt0ShiM4cIRDh2PluBmB7mi25a9
HPwvvuk7xFuj5bqV2evlFkQRSFNmM3aQ2L1hV/+1CCKAsHCB5Bmkh2/INQslPTrF
fDDp/uz6dbsWCr8DVnmNsSDzht9laPVoVlqVZkK9SKCYSSTWusKJxAl83SNiYMfj
Jpv5bUcF2HQO/5+5r5mjfhkDFXakUomPuOFcUtW21KTiFmtNpn3f+6xI3a/iISb0
H5VWDBVg/GKz1dOYSsqMykTfxAlhiMiwqF6mg5CwB4ZuN2kpgDKkwIKiH1u0H1ZU
MiP/8331S9cQtAMjZ0aeUre7Gtj3aCZ31XhwU4Yu+dn5iUMdLFIsq6mC0nbl/Qpn
sJzBcWQZyi1TjdLx8/s6BAnWrjZ89w3Av36eYtAsaGCxMW3C4xV3xiTRHJ/QFwLX
UWcUlYKa6lgmEKQBjWGUabR6RA7pRiYBiniN9IEJAOkkbQPFOZKzB1EHqUm3Tc5N
tpyer5lFP2fhiI2x7nnJqjt4dCcR7EhK/f6KaW4G8f/cbNmdX/QXNrT9XKsAvrkt
0LQ1ppdjaSRwT99MZmXNBO/Fy8dr2oBFo776quMBSVAVRxIIuyKaQtBbYxhveiiM
2qXHa/0Vl33Y4lMxN4QW9avcL6Pt1VW4Y68Nzk7qaq4paYRGQyif4lukPBL9kXFa
lgSBJ1OTloL+tOWwO1T+PGIGEsYz+wIdjbPmaY03ZIRV1MHVpg3nacr7KelkqEX9
URuTpaZ5+hBGtgOvrHU3DOcdU+m7lAOT6QDy50QIMP+pCIFErW+ixYSD14etkOnp
ZhapLjDdE1/2G+uTRZadUhnVPrc+dfbGYpTd0+JUi97SEn+uEpRo9czzukDp6mLj
3xFqVGjKtTkVc7o04hN8Sxj+rUOaY+RAHlCRL3LG90ZBeaPg52P0cAwkphx9OMlk
pfxI083gd9e2LGAPBN8EfMooW1MjFC5DzMibKvBU91lXXm6CtknIxampqRqgotjk
ZGA6siOOnhB+QhtXPXoqqfcFOR1g7qH1qBYt+HXmdyKegnafXqbjULY2ek1DG7eO
AQ6nHaEwICAgJqonRbAmdjDG1dhhGEIOUU0jHIfsK1y97aYhjy3QGZUmGhS0knnZ
cAUI8478D9sYqLXCfkV1UTYyqRJ6PYbO+4ur+fYhqrPnuO8N53ClM1aiXw/klol8
E9ijqYMmbTLsmXXrktYccUBdpXRSqFwHaREqxsEnUrcTCxOpYjuLVSkGu2wzmAWP
ojXdtkyDZZ/kFyvAXQFXZVvhhZqepxYVO6QJX6/5vt4ZacSJBtnFY2LOAWDv2XQV
4aY9kxsqQv5T8HqZN/DgeUFiO8QBGlDR57eAeU0fuh8PHWQYQ7EQv8pCllP5U8ob
c693H2rT0d/9+DEDBN7wCtAcYSlB1UQmcB7/H2imQjg51XuxVX9TF03EMk50H3SQ
alvhWCjib6Mp8ifYVQgBXWwcpfbFH0h8qboFDxeFml4Dh9x8wbG7NTAzx1MmHU8u
QJIQ0k/F7essLU3eti84WUse1cXr1lik+6w51GwsfSy3YlUqAe/mMJHftOmQm+1t
iuK5dASYwvZsFkDmsFtpZNJHasHwwBfXw3k4q/Vx7QuouabusTiWHx+12zU6FRHd
jGAXJOWzZLgQOB0VTOrGuSucvNsHhZtYM8Sjv0/nZF0In08pscm7XrIgt6dIBJuF
yMKEhhWNzv4JpCmnNGtbRD26LKmMYKA8Y8UBJbw475bxU1yqQ58Q/SogGPQ1sp7x
k7yvUhb4DlV1KP1ir7U+SrIUSkWaqAJ7qlMbfrWsYTyOqevK8zF86A5Dek30x1VP
YafvvIAX+x8md4iN6in/zrNppAD1OmxFBKPwVtoGMAw1/NR0uWRvuH4ujrr00cm2
EutE3BztxEbUBMlD9mNiBaNOTF/D87F1Fhts1sPW+ZGQqzS5R4DJwMPD4fXgGzqS
KbrhLkYSAerFueEF2LKhfFNcnMPVJjBjJjMl9JnRHuFrtMMeM0FXrxohKA5z31VN
Sl1NAxeP2HLiWDVCrQRuk3JaqmQIH8yg7KqEYmAepJQ1jUQ2C50tJpbXKPqnrThd
Kbhf3GbaSWV7h80eD0MylgNdUCrXZgDMe2TYITYtkbXatu6a0p/9VpLkq4DP2HIk
E2wJbmQCz/scMiZF+1edtb2tzva1E5kIu7rTUghnR0q/HlE4LBc0ea6rhxJ5F+wj
RLZIj/UrNxBQFTLu1Pmj22ni5tgU+d5mYZjkoNKZKtfS6wH9w39SrOO4VYP4XAwp
c0yYRGcytakX5n2UxbsINvtFa2hhXNsyG3oSTBy56QYPxMfUMqqt9qJ5J5AgJoGU
zsGK2FltFFp+ZKWC5v37m2VLvevcJMAh/Ksn75oY+K4d55OpQiW/3u0KWaUqUvjG
bazBYYzpVdZHQubUbLbevHvHw1bEf5LWI3XSw8M1eWPlEwAFoh7JtL1sF8Jxnuun
lpGiL5LGJ7zm9AC+BGLyBLmOHb1ixgeoz5BbiCIFwQ4Yv9X2E/LMQM46MdSNxBAN
S0IPWlCE4pxxJVs7LqpO0303rOni0J4LkHkbWWJhVw9UB5eYTZliOXPspGtrHUoh
X0zholc0UjNJZF4TxPZqQTvGJ30zG7Q9K9qBjw/kltVV4qOkAIwkQFUApwpnUTVY
HmYDs2kYMTiNmz9X8c48I2gcrXFLCbaTcgJeoTp6qezychVlyS3TMwov1+O0qs+X
2DIF0Bh3pL0h5VHxYbouEXXmzEOawgoIbaagFt5WGPjhWdfLSocZs+IFY8+tRM1t
2Gf2ZaEAG+Z+MY7/8VSrW4VU9KcKLrSIY0hqgBgd+jEYCONGq2rzD9z6oKUo3Gyv
K5thvbY6iyMewUYz+sZ3pU++7Q9fNIr5EZ7ET4IHPY72TTjaKq33zMeFMHcss1JV
FBJHmvgvSFpKsXLoV5p13MrmXaAQiJcly9EJ0yIRohT+JvnNml95D5R2WGRYWiAn
Od8sPeGDeeyhsttarC8AKtqxcsgTDolP0sysGc0gRI6y0QpMT16X1aIGS1xYjelv
IXOpIy6AJqktzMqofUGrQ1jjdEntv1xKQiB392iDLijX2/7UoX/XX+8qqYTYDkCm
RNYaAW7zO+Hig8U8wQPJjIuLe7NPFqUK+Qh6FYR4OxVO1/z8ILFjg4nHLOnXyexB
qYSYjyjfJ2ygRGrZ/XDQwXNyfFCFpq5douF9S71LcooMLYdxpJnK9SeBwllyCQkx
iVI17xHLywEHHJGLUuvY0qjUY9isZtcua9cG23dvyJMcRGP8IkW/Sw1ZIJ5gkJie
/QY0bRjjmvBx2S+aQjRtw65W13mD0uUD1P/7HFbdqHfbHC9tJ7ic4mMMwF/T43WR
yXSLhZkBc0ZZAaxSElMPe9gOc8aPECgEBFs8xGHGAbpydI4+fyNFROU9aFUR+mib
p6E4JEtnrQce20s1SN/fECaje6uF/ZWjdj3dKaGbT9HLbnIand0zOqNyOgd+7y2Z
3FpdmT5ddz+6DGPquxm1LED9dByQ+Ktu3Z5xRYOiw9rs+wLum2Z1xxJXE1+QzvKi
Tn7gLpaMpz6VvkNiolKb3yZ0BgTj1cnPmw9fLBpOcAKL9XwJ2fm7+9PBu38U6A4X
98uHTuQ0DhU9PGdRTSfI4Y/Q8RCaXqdnPyYcAsFCXlaouU3brg70E1Fu9Hh/E1vO
/G2UcdofsBpbT9Z54yjraiik/IGF6e726c2hTeGlo0tw3hG2mzY0NIBkLEWZXc2A
5Yr3CXg8YsMNJlqtCerfXze8bjIg63wDb3/gY1sSWxG2Xf1s+BeHomjVta/EA8/I
+ivBax/s31PmIBqdBNiFg0HcSFG5ZfrYAwwllF6qz5ZOmtEJsajh1nBdAoImr+yM
IYIB6Bi+8uUH+Wdo5YC4QUicFfi18VuHwlDjl3t4TRICB6HPc84XJYZbBo+alvbj
rkrUa87L8wN9EmBSrrVdbGPsKpMryLtCMekx2K6AqDZVQ8RALB4Oz/iQdNGIrAmi
KkhfVMxBPidEkWK3ypXaT7Nok8HEhn1zyyhIBRp+LSYDAZu899zq0iUlTvnpLHdm
b2lD3H6d+EeUJm1UlYZd/DmX5gA48lwPFDDFstD4952PcVlctf+1Ejk6JemYo53z
Ik6LmWZUauXXP0f6gdttUUv/St1uq5qWjUvT1+AgTgiYuyvemn/f2Qj6LVJd7gdj
jlCiNPN1swCFNToSlcTQF4iAtLG7Phx9m7v6WO34ftUEKkgFdGODRJT9EaJo7wVg
niCLKdmK0o+FwxAirMQLyV3P2WiNNFVDvXe90R01bamU29ha3BbhwPSXOBszvQQU
RoJ5MFGOSI6BXnM2T/HUGD0YglfZpBtvMr/7/fJY6cDS5VKH2i18DMrAhy8ckEZA
sSrkQisThYcWj9M4XFftlZ0DcPBHLC/6Ldg2pR9/Kh07pelQ9Mmus+iK7Fi0xZEB
eTLCVC2IIa6cTZjoBTn/cN7BC4osqL2ZfsZ2zcydrH54RgIT9YS3ny3MYVeMxfrr
D+0X4eCxxf+F0dujroSNT+KYKqdXzrTgf0oVaUczurPFcNOk/7Gmsg62TBjHwToa
/pNgo2rB9WO/6G9DywYLncu10axEbuKYqT9Ka6s2I4rCEwlG2kMplOtLTiKId3Q/
c8ZsNWeCE3lyLrs6mmuSe11VGoOuag9u4igzKlTf4O5ys8pukArAnsNplBEVmG7z
55TUox0IrsHspLCbvXl8JZnk9vFKpReDReEl0kv3gXp1dzqzUwle7UtPMMErOgWm
TwbMAibQlTnEIb2NWTgEWyux2yeQu/gzHMmsuLyX1mtPIUCK1OtS8ozukZUDkBOv
s+V589MbDTJpAEEVLJOXXe5k7AnKGyEdJ6wHHGS9iFMV5+2bjQPucXIE6VGgYZcx
pJRnLFmnJgVtj1bsB8cIfN9+pGr9CfN5747bapQMW4PIrxYkW/9LqVRv03Ha2e40
9RB3fiaMdZGhbmADoWpaVZmU6ujxom1clzzOaa7RQgDiBSUUNGsf+MU4R+ttq+KM
u7gn1/eedPdbV/2goXABxsE+XdJMZ1pJ/rlRfVKGMdu5eAVbrbukeLFEPKInBA+A
k0t/za2eSx3nhT3vM+w1aXkz76ka757wgIHiKkKo4b0JUbPHr+WXLgF9XfL4DxVq
WGCd+gavQo7d/PEox9BKjrL00Po5xPVghIu+PO7QH+/GqD2ehJf1T8MGnHhqXqXQ
dmvLQT5SCIK1DsGgwMcCTCwK0aYRMtMUr9rzcoO6cCsNfNwq/MUrZI2UFpsMHzKY
nkH21rnqsCqDpRrES8IwsNxjNvhumRFM+wtPHXqEvjDh1zpXZ0uNbeL684tPRMWG
/giya+dwazcJMoGgaQTUsO7/O1FQdtRW1TKLmtoWIu7SSJhiQLrHQBwwDa8xp7sI
K8v4wOgto1fQzPu4qkkzFiNsbFW0L77oLimJtMMPYr8gNEztynadIL1U6uqAqpcJ
uQdT5gQgSXDTyBE6hH9L0wrf/sz7M7VH3VHxt/iQuKCE0yCOF4UeCynUi3Ftfk7z
a7cs6vhQa+Zek8psRtzXmbg4yDV1BfQhuxCjzUTuu1U1dhGD2dNnOKlvr07SMMuf
rwq5M0RZedcE9Av/PU4UO4KycIGqooMAp/wav3cXuFyAUPLNja7H4ewc4+ijCcEY
OKQTA0I4fmf8yn3BIOVeW9FDFvXMIQjPXzgjlTjxXQhDpyXRlWagtKHucIpW6os9
pYsAghSHWPoxH4VOBsyEMhdQZk+BNXB5WTZLgrSgHSY67MvCyN7O8VcbolTfwQBo
gmDPYvnf+7ndYoXtXqLHdWmGXbvwD8iyb15oni2XG1fAGfVlU5Tl9Nd1MiumY6ot
iw93sD5yCEEuw4PGuEhpfBf/4o2+CHEO9RQ7/W2JGUxtbySeGzL4hskCpcVZElpL
Z6/AC+qx50ZUoK8g2Z4MEncAQIHzZxSkDnmvk8Xp1ycKcbFuL6koHlphtCRw9gKX
IiJwmoszdu4XJ/PjszHfmL0fq8FiBF6sJEHaqKgUYGyhtjsviOM+5ZImBr01thCn
h4siPI1k3ALAGHcKGNZiX8iWwCMyeb4wfuG8YkPkwPd0l2XlP6JFigISnwNfw/Im
mIC+H7Y5HYlf6c/ug34VcIxkd/kDVOTPu9k3WoNoI+QQRM6AkftUgwpgkh7x8bbd
DIPg0hx1wLf7exmQfo7MWyTNHyen9DYKnbpVKJjw+yNxVd4epXFHnALPOocgCP6g
CrMFUNEXdVEP96OoVNLfyPwcakUG0IM4zymFIJtMPSHxnpvx/OzxlHsKZA1CX+J6
iF7ImZCPfUcbAhhvyfS9xUvXy9R1RShvjbdLdTFuPr11Y5bE6CWBqnNdLcUOZJHM
ub/5v7SEKh2/ziax0ogGm9gQlzUrWfUFiMrg7kctZgmN+k7M+a2OwUiKZ3LTWjyp
NYz9WR+4xmm6D76iApjQR4BS/3sr/10C2qsJcqK58sIPh/EYW4JL7IURoqC2gNnj
u71LqvpxnaF7OkSUE5NpIJq8Khm1Ed56Un5hP5+Y2fv4ZCYQB3Zxe9t40ucxHNnX
rFVA17bScgeleF9OGLZ+CpXqzpa0NaF9MbGOaSGfOdufYsPVcuAbjwQlfnx958eC
JbkRbmiUYDyt8qD7UMyGjAhYDtVZwTa/d3Lgv6fYofu5ZII7sqmbt8yjO0YbGrcn
nQaOo/rtMcDwndW6n8L3JFjJ2f07OOKik0V60vdFmqbXOpfacO6lGTXaw7aHelfm
lLy1P6tBseOM2d5iNd2Pv3G3CrKmdhXZPf0U4AMQHCqwIvF3gWm8B0hbYznx26UN
cdtXtCjadGbp+kqzt7QfF58kkn1HwFh7TQRcuxuI/9SXbtDbcOmSXJmXhXqw9ggX
SLuE4UawQ+mZs6H0Y8No0XdePwpoW3gLC4IljKC1wRcL3rcAzDELDmt67qRmAazw
1dw/okaumdWi4g3D8cO1ZFjeJbfoNPelzoA7EIQo+23+Vh/oc3Ug/DyHTt1o+w76
mLvMZz4hdW8idmyiJc4Z1L0FtlaPKOqWNsJ2+K9EXu4FhxF/ZZgekHViejnLNeBZ
iFCBY9wCOinMI+70u6NpM62kVJ/QDGR/RkrP4/34U+PPBXnbe/wNhIYia5VhB6mq
dU8gvDk8OV/LmCEoNJNTjWUZ5UeG8wFjK8LhbOyBnNOBXiSESqtnrbL37vkrkPg8
17wAWvkCDvkq9TGJXHgCgDYyhT61+Gx9c2PwKFCK4FAIpNRTb4godBVeJFdZ/Xrh
XZIQX+A4mVrfPbaUEvzzPNC5Z2SMOBry6NuGsCA8bUxBxCWrnf+o6tgoMjZIWFGZ
xfTI483M0GQIzRIgMNcqtY5/NFMZ8qMDp67GmwRLr/P0wbTyhs/0A12xj5SJCZpe
xgYED7qi/bMOT6TI9KgXB8wILpD9qbbeWELXbYcyWqFRCUi7HRlGa9ba5buxi2dE
3+2yORprkskTlXjGTlN8MMXtf2fiqJ4NeWsxBb+wSmDbAPf4Z5uw56/ZfSuXBtQ1
Le0JHCtxNx0Q9S1HXdOX7zhXIOFxmH8mxKH+/kDkkapr5gJ+Z4//1MJA/T7TiDWU
U+jWNdtDkIm1C93xgzHMUEMONsfvMoZQEibQinVOsnP2aNkCeY8YhkfkeyH8zr2S
belDHmbf5p1vsXC6pfkUuEwZcNASxQr3d0N6z3ahZWpk7Ukk6uRJz+rVaUGAIPYM
rRZxAgOLADRcg9Df23/8Odb8MLuMHvM5glj+J42uwRME8jNFYVKeA3ddpR6JAkDH
3RPlZOHYbp0EPu0YhqlJ8ygyoIRHcfHdyOsKHRMquiE84RmGV053xPC/PPTONoT2
t8NjYMO/qK2PVaXr8ceM9cvViKksWMSwxya8teH/cgEqOV88vUC9+PdXMLt+t4vp
gqjgMG4UMjrbBb1nCik1pOiOhYnqHyDn6CgoRD2GiTBLbw5CAxfIL9LvWKaUTsqC
9MutSyICZohycp/Xt0F2kJ4+o/TjnnjoUmM7Ir0cP5UxjdmUnJRbHzVzbPZbMLnC
/BKHSkSPca0boEvHnmNaUv1l3nMqzA9A9SyWMELQbdCeA60qXUYSM4ssDlWMnoXC
xUNK0Wa9DU38PcBKOrE3gjluCyE1SpPYeYzpWVKNtAFSXhzaXXzArP3pzOJkBRJQ
y++ma8EeoMRaN1UnOTnwOL2CbE4ovNR8d7m7fMRDrPSOChSjSncIv31RIvK9d+Rq
C4HXFcdqdDTc1+1onpSYaFdoecNAk61gaUqllZ4oT2bbuoblX2iG+zGu5arC7Stc
sU0H7zvPd7l9ltyZMmRyngwD+mpFx8boMKHIWDCyVitAgza3oN/ng1+Q785g7n6f
en/aU7Kn/SpbF1ebh+5Lu79Yr65APNyowy6nf6bsQqrQTquLEQksTdYtNg2S6Dkp
Kg9T2+qIZxZg5wdJODyka/DaHqBOBLdavjapAp9lb8gHQYxbdb6B56DfB/+WbJ1q
2R2NcOAIIJSpCk8Ll5+ZPPXGv3QkrvQ/9ijPenLH9L8XC/Y69LxFu2dMs1fv+06T
j5hJdA1sAvuszaHObcvB2A+2sl6weSR/G95EbvQb2iXkZdHtIlvQvMbb26J6PWO2
+VmUh87YRUmwY7ycpew7VE2pRmorJ4F+qhi6/LmRz5W0QuJ3anKwLctioytlCIgC
Yq1tLMMkzn4Sbmah6mQmiiaLbA4cz9LWKqhQXFI01aFjKjkAWu/Qv+i9/q0ef2D4
IoKJ55t+8q8MmDz27J6hfNgFw3ZmZbCkgUqDl7rwq4PicLSu9hHxzby6KoXzY4ii
OXdDSyh+mKFKXc/JrAZMI1bWNdgDLCeSUGbIkkTrYgGAgfsyvZ2SClddY86JHE6I
QDO6CyTShGKShkvApgs5lI3mkbnnPK7KWbwumNEAK15LPUONYh79PwcfLlpWZLEI
5xA6+vDb75QT6dTOyb54DDb1ReypLrVqS3EuCySqSmz62buOmMIlBD+Elh+VHTCw
jsFLyJqwLezpepv4ad2ZbkkBET12cMEUdA0HfGp4yH3fAxRtAbY9L2qhn67py2m+
neduOrD8XNNwfZ9s9lp4UmKPVdPX11AwK1Sshi2q4iiUj/xmmzuUmI/0QNujeVcS
Ql79A1l5/ULrw0mgK2mWJ80GuEeCtohde7AuOpXecLFrmVzUgUzmubbuRbLjDJgp
yZ+Z9fy3zR4lzfM8+yPoImjcMJzqieCcCuAvjTYboFKATyi5EqBmZ6w6gwHxz7Br
8w2XBcgQSpwC62Q0bT5wOn/iwxai+VW3LSNNAGUWftl1mKHrmKnABo03OyrSxAl9
EuxbtNy7o74blDzkqtro6V3xFP5Vhh/II/1my71Op53XLfklp4juVTca4QI87hbu
w3gpLVqMBJ5FOKbLPXVtbSwiSINivtQjYOKIQuT4GwCc72aMVR/5VJuSpboDyETJ
xTvHURPYeoj3da2g0K9jfnVNp17ad+Xx3v1Tcdp/XmuFs/HDQuLIwSr2n3wCCF/Z
9MUAHy0/Jjh9UdGVM+EEr/SXe3Bi5gLTH4njKDCR7+5NfFps5W12ZEOQ04wazu/y
CBG2it8VWNH8C78iklsji4912CCr4xKYeDGcxXdMMUTVp+0/pfwVPVy24O2J9RD4
/fkVZ1LyrWqnVqwgJuaLEuMh5hzjB28aJfZI5DZRJSBL+S9bsAmF3/YF5OuA5QBa
QPhgYpvhctVDstN62IsGXHr18MOPNTHyi25EMjRHNcYy0wfsnqtG51k6OL/GKSZ5
NjTdyQK2zZo4JWBh6Ynlobs9T/5SmqtAz3K0ZXR366sBhRq0M1h7nAyFWmYbR2Wo
/+TqKghe1PpRexjfHNsEEqqL1pNINDaHoy7+8KqGPvLVC9SfvCRBKeetKL4W/6nV
2SyD4hPnZwBWiOhILF0R1GLCdGAy12mrBoddf/y4gU8d1NSDJudCRE2X4siomXS4
JbaZ2CADwjPNAQ9N5cnWmKv7x6tKuhyy3ubaUy09+ZLQ1J14AW3FG+pbrZqd0WMH
NCC1Mz7mHEYyyTG0r8nErqiIZQEtu1B0lF24/9beC3YceUqTgmoxkkWleG2LHiWt
2m55gp6nphf/tEroskoB9+K7EAytp0hgxS0HXlShqLlRVqv27+KCMWOoY5/InRlu
lTQjr0lsV3GqRF6R4PVN4uuB0dHxJgOMx8vk40bgz5g+BqA2TN8BUHbQLTu0cDti
xxF2uLd3jBih73QIxtvrISLv3mv1NPcI/UJjGDknuefWQ7keWaCOplf1OZckJfkm
fTeuuLhAK6QHuCDTz/u+UjoqhTRDXIxZxCA3BWSxCkfpdibqRSv+lCogm1qqJ90G
8ROU3xl78HgWqEvgoAbkIqCWpV3FEGPadAAK9nlh3RI2VHEj9BL1/TfkvE8RFDev
9ADj/9RPHLElvIvMaFPyPRngojnnzOp2RtawRqkZcV8rQ/igpxNlZpANazifY4Wq
hqqA8W3QS7zhUu+QYB5KlGgVNSK7rDNHRBGv8Rby9/+t4TZTedQfnB3tJ1pnGS3l
DHdKgqYBct1FXbEZ79ijHrIkHg7/68qAqPoRrGL8Q7epPXiKeWXptzVYreJmE5hr
GRprBhlmgxgnWa7dyOWSaSZoNOVh9qNKRc4uQB6o2wDthJJqS5HiIeay7MDj+BBO
3wnJPvFB2XavxupOESTTxsIxA8wWUzqL2x7kyKcf0sSehcrbIXNqwxKRNKOKIkOv
lQF0fuwUpQ3ryaaiG2NfHpwAivWU7m0EWDuH+XqNsI2Bwn7MejnNqNRVLTBtxypV
0ziR3ss5O0sUsSwYaI60OLi+V+L2YTTYOGSq/5nvF9L+3nVgvynPm73ruBgl186V
rSuVsnrPrguYEN4gLFOkoWWgCZTmN5sG0hZLr0SACJCU+4Fj68G3hlkuVL4erNAs
FVQCh0zPBJU26CjPwZ9DUJGIby36Mk/vyIjem3AqAsuyx4qz+MXqJ7svHMKq/bI8
5cWC08B96Cm4aech3R/qU+k8BIR8IN392ny+/Usw+oSleUFmAieWwF25I3yLCurC
2W1dPGbPjCm/yfVggrqhdDOrHX6tsJidXtpvBa0YZffHeatnqhKiOgeOVDdTxc27
gF4KBWBJbtoD8vKPYOMCIo7UyoGOGZsXIUd8Z4327qTu2w0ryxgpmQSIiDf3mBhB
U7mt0ZM5G3eeq9BzycQJ5DBs0dYH7rt7KXRLIkbza2ffyVO2a23i9P4xMhFdGZSt
rjBagvSCzTnSZmEzrpkn3sNLZV8waqnDKproYedgMiPOFSUGrZ/vbS5pN5nCGwkZ
HYuDE3wbQYw3scQHY07YAGrpsF63OUvihrcA4hQwmGqfsMCjJ2/fonHsr6Lp0hL7
lhmHaByW3K7Dh8vBcy9s5Ce283kObk8umt+5XEQxVSwBVWQOliHTdsZzPxnNQkYY
O1UppS3rNOT7SDlsQTbuaAIqXKQUimqARrG5vLUXkQS/0FAld086PurKwYZWef1A
QrbJ1wRJbfr7+Br2u0nMJgVyjTy2sHAr0VWCoPOsvaTgMSxJ3JBU90+8l3FWXgL1
Ws8pEQaESqS9Ha4zx5Q7K7GFFYR3hLa6viUNm7qsvVL+INNXT4dRxXACvSbFmc2W
zG9mRu09V+gkBcEvTkB5ZK/M5HVYWJsWIFLfCHbtvdrKgYbqBlSztz6ZCNt7jWGe
xwL5hBmkTsB/AacNNHlv0IoWR0gUP1Pdkmpk9ABjSdxLAp5T7g0EMlBPdXipjsEr
dP2DH2If1Qzr+jLHwpc/SEXbLc6/pWhQaBX9b5m3RWS7Zy2WA6QNEXg9QNl4DE46
od8THm4yFucr8k2YVOjBDWC/l7kzh7y+hgf6c76a0MGuKr8i035T6Hf0iv6nKBKP
zafasHtExmsHYAgLSA69cwo1I6ZhDF0sdZ1TphYcqIPktLavnOVL0Lk9cp03rubi
/uV5RGn1KMc1B2ITy0FG2YizIxgtY45sNqFzUrNPxkKuGCa8jsMVY1YB3CZlTM83
p0sXbPZHAImJjryzwraxz4sWzY1YwcXVnrC8HJBLU69M46UrRvWbVmh3+e+dsHXy
E3iYNgogsuCs9JEuBV+ThhnCx38E2N1hcT1hJ4SB2sO6+PaJ6rn+H8v3Ly1BnS1E
tZ2bISElbH7h2vdveaPb+2D6zrQLAOSnoBhPXXN1jFmLmu8oEXej4J3MMCNubksV
DSU+oACDZXHAlr9kMm3M4Noc6/XeYv53xCeCf15wFpcPHD1g/r1rYijcOc/6BjpI
vHS89vDn+N65RpuhvYQeSPf4d4QOUf6A4IY9FjNTD/7TDB04lzW12CrcMJ8BJhCk
g4mXI9JQkqZs94SooHRcFEOHpAUGaG0xV4jc9SVN+03lLURMKnhYGpZzcP6Hgx5u
WhwHhEivrFBfds+xUI71ZYtFBv1VrEl7ztdK5rjPELXBYSQd74EdDJ6RMrPxxjm2
DQgMq8nhzbNQmvG35iSUC+fJ2395yndnnNW+o3BUJAqn9Q2O4XhYUlcY41aq4udY
yHwxujS4gWhDSmo8TT7yXcY9sM8AQUBF7ntC08/2TepnhQRkRH9PN2Qggn0Y9dCW
49I4F+idk5Tz5q6sWqHOL9kulxS0s26/ziJlKZdze+/XBcz9e+Dok/Ydlh9+fuOz
td5q+AD8pbLytjJskgJ2oJG8MS2ye5xB/OTgMXZpzJBJwB2opu/+Utz83HpLSqTW
kv0JvmaQyT3W+psE46yx3zzCCj07ZyKMCPI38AB4Svss0usqS15VXz49ec19u/S9
cEBAzO6DJ1HF1Bwh9GLKau1o6ap3b4QuA6QnIIWcxD3Dzx5Thcv7Mlkg5RmKPBZW
q1B693KheI3vH0zJgky8YxqABgA5dxy56Yd/IqcxZ1d8FMPp/feXY0cBySvmUFiN
fKY1vOqPHRTSpq10cFkaHkfyobBpTsNNdoecLe+sTftXd20k0jYyYqw0hDxz5dnx
73IQoC1Xzm6GDy2Tc2vjMGC9CYPl/fBC5Pio9LnAPhkvqB2+7dydWxrNwcB9a5Hv
6Cz0k82GfpupH3NwyexvJimbstLHfxAZCKbMb8WF9JdPQnLMbLjEaUcy4w7o59iU
m1hGFTNdVRlw+eCt4pGzCL+2JAApk/3tEaV3HlJvHucA6XgaxYpea/7iJ9ocFf+i
4Lf/lcxkBQOfIyyxM+cqiEQTaJBnDFGqd8j/M6Tb3TNZH1l2AVt0S1v6U/5RZA1r
JU3mwG2SRgip+nWdwUPW6p35TjDrbWN3mZOL89yGB37wjPu0BnHZuZJEcivPbrib
Mo3fSOF8SXj1oa22Mm2ZMQpqquba5Qgc+iTay+efljvCyT1tSvFlxNLFUiE36qss
Y8A5zpHWpISygrFI3a5P551JNN8SLmPlZvVWgVid1VvNxSXMJkzMPLyvhgDHA/av
GURCmmp+Jqxq3OmhxVuk4R8sB/41WOA6CL8fgtJm2WZmtADH6DkMlE4YxVXMCpBi
QH/YCutaic83V9yM8uT3EK3KO44G7vEw3VOojgoWEFdx37tJ1gainjEDId18SZlr
kiu6SU7Bbge0AgJHmBjJqQgwQcAaCYpQSrktMFOEMdIg/mOKFze3OQcSgi4GLiZ1
4G0FYNCPM9qWhyAuV5jvOmTngF49t4tXDL1EhqPsBipWQI+fM++dj5MUvsqC8Rhd
RysRw/1g9XL3Vo9tyyZPF1sQ+nrHxZDh0DHHDw6K6JJO3cOWJNxnML2MRgSfnrYF
zuO54dO9FMoiGcJIYzsmRdZ2o0YuNJbo1GibAyt2Pff8IhW2whlbYcFSZh2+J/6F
3Zpo9PjURaSJ4a+4RdjH2YGxRxHVBPOEznRP4gcZXShCSlxjlQWavxNbcz0Ebc8c
+qT0+H9cO0qA44mBIK7Ka3YYrIj5flDEm4gf1TdHRJSFoCvQcsDPmIJL5o0Wx8m+
Gy07rwlnxTccKCFOb9fCQsoPnboY5tWl2ZIGspYMslBoTh07/ddCUK6Tq420Q7NQ
hgbzN2lvXP/DcIXuBdPjAgAb6Va/aO8ciUWo2NZhvc1/xuiZMFZuqiGhWrZsWfps
V6prOCidNnR5S2197SBBCYPYQX2JJzaEBwGBJo/ZJ+T1MYE5wIP7GkERhu2+haX9
q1f+Z9xbsB5Vq/4XS6XGi7T3x/QQ85LI9rMix+7hTuvP5pg9kjiGgeVLKfj8UQzK
bgH+OdrisvHgDT+MvoLyZ2CwW2TiWPSiZLKu15zGdWWe0HDyniN/68DXUuhKm6Vy
eKTC+/dWUe4PkwaiZFn/Fqugcmxk6u71mTgKUrHQSBnv6sHI9RUXSHdeu5R+ieKC
79wmu5ZFRgv9yEbduAIKchwVm2BDSVlGDyC/Db8tl+hRnKUZu17Iqh3nfRaBvWWN
Gq8kniCyFgzlYx1dwYHhCvsCidBPihz8b6X50yssI2rj6TQ+hGjzRDBXVSPmMrnX
RYb4geJ+jpsNEhg+DMCZASPlidbpSkBKHBeaAUCFIWhlaAEK1OLLeNPBcTHzr/0t
R0+nJjszrGqBrMaaOdiDqvZdvx5ybXOMLcFV2n1Z/Hcyb/3Xgvd4n8iiydkveL5n
sqsquFOjqQOST6Ujj17kn++Kkq/ma8fAzrXJMmKYH6+gunAqVv2J0r5Q5a76yQyk
AhFkWjFgLk06leyA69o2KOWQWa+bCJFS8aCWYhtf2CyMzdaKwAqxImmM3WL3Ntzi
Yn5jLeunTSgloMdZghNFRCRHuLvD3zWXOls0wpl8PUoIrRNnfFd3vXtdSEwVlqn4
A6muyohQho+V6pu/FKUWiKuYOw8ALWMp5tqcrk+z1ouvmfyCD0RedKNbylNOvL54
gPORmGMyNVLQVd+3D8HpOP296j2qQ90/ygbGVZuLJRGSLXg5x4AZFK1x8Q8t/Sfe
ILuOlIdJdythRMa9FulWEng4+Nvj8Bog8ZQ2b59UbBH4gU86BM0qlzkPBp9slsNa
ynSjHWTeychnub8XaigOBVD2hvuqAa69+MeSvzGpoBC8tRX6o8VooVZ7D2IKpyeh
mZpCJr5GQjEnigggyiDvqPNuxjR1WzYMwwuwC8/PrnNFNfTlavKx+v0x/TCupSU7
oNIlN7ksXvriNewpTVHPuE9oTz7mukwGTy/Uz0hb4YFUsRE7GLeGxZek2Vk1YsJX
A+LQEgSbsjrtiL9dnRAlYyTy+XiCEzBn2LeZbYrIs1XJiQ1rxbqzxwOTs+wuQzxL
QmU+jlCfGTXHbWrjF4OTtBJfjLVflOUHIAtYAfm0hhj/C6T+2iP4M11zDBYEEFxx
3GSXNw8eqcDHRct3+VGrMgQpej8tzvrxLh0qHS4nY4D5yrRAcgdKThotWRFNdJJ+
2VQ1EIKlPqFPQ9LspbvUqWZHHRpkbqDEVFKdWfyiM9TAXCW7091tFp3DuxRPyU//
4br/zbkfkPR1S4InjUUgJfiYuXQOs5gqiy/Hzo5kXcISDAzX7wm6Xnq5bslTILeK
P70KYn/2qxdoc41aqSPEGgi91dNjfGLgtiAHf2akKcfrB9AZ86Mz8IAwg9BWTFwU
DW+3Nf8Br3OOVcCSLGIjc5CzM4qlYaS0uvfzQvhyE7t7ew9oLOIWdgct5omPo18+
O3AMDTUsi8RMglwNnVaSZPwDzh20MvAk9Bn62LtdQh73AKZCbtX5qT8Zrv5jukwS
CIG4ME9t6V4gphIHNfaa9lAvGSmCQVANSGHLXBdtfMICUrHaL+yZ4w7nPSkSfn30
V7mT0N9IxW8iZyF7Z8IF+zT/7i6aCzhQ1l2r1as/XhVHMbDq3zeXIXtzcFOH10S1
RG38wc7+kZKe/PnCk2xdPPP8IgpJ8Ph9VLGwClLnbKKN2ki7xwmV4sP2rKdeaa45
2BvpmTr/u0Bb3rgd+dDdeHuEwfOAgO2zA3cYKPPB6Vw4VIm/u+t7DjzaHwLwFKY/
ufIzwksVg/vgQ3X0eo5FhSH63ICHamUzOJL+lbVjgyirRbyYUjLNVAhlfxa7uRjm
ej72FeU+E51n0/V5s8TL4lDvS5/I9uT7QpPBWv82Rku0/BdTKajuOXCdtqDimeUL
j5udMre3mv9VPkF0G4N9A3dtzM0t+yJoJETvbHgpUaoER/exXBMcZ5fZdsFoqqPy
8H4L6IhL8/es5Wkw207mUiNClxocBea0Ope23xqZK+x8xORsvSqyCiQGB7Vrd7CJ
Hd7BNxUlHFbz2UX6P3xIBUS0N7tsVwrrSaEosiR5J6dROcKcX/D2UjX0n+RBHElp
FkU+1jrXgPRrCsEyf9W0KfXlx5KW0a+HtHoTgXFGKuby13WKfoTi1tc+TqcB09jr
vre/6Y32vuvMmNnYQtzvmnH1+jEGTuzs3NnZVCIXxTgcQPL4f6pt1WQmD/I5aOOd
dz1lbyQ2KxNd8Ll7D7mQMWy+wueBnZfFtIRRnAmZ2OO/TKdVgAOayYcKzlmJAtDI
03oDX15bjYKK1hUFLhSTSZ7Ab4Luua9Pj62V5K0x56pxlrSajjtih/jjBwz4zvaH
uxk8q+N1UL1Ks/lZLTicOFvr2QUlzs54FC348U2+YNDL6iH4GeH3jEdp53ppztny
4nht/3lknAzsp4yzBIMMADo8BNw/bOS0ZwyM9bCMOtbOyMgl9Ym2592D22cN0uGW
/hF2yQLe7TzI4qd8oh3apwnzGGCQ1D93cZEbzXTEocAQp4vIoe2gkB+MMy2eR8XD
oF6xdJ6HfwS9qUE0+hbarLLR72gg84FygSQfXywMY92AjGkGzdmsOfs6XHHZp4oh
Wx4SKFnq6wmJ3TtEQZ0zv+e8OLPu2yIOGugHM8HGhe3hnD1ty5g+WlDlpHRqALDf
UNuIwuh2F8w/Dm5Y++AedVJol6fYZa4/b8u5KZVO+k5M6/7VcXijqj2Wu/rznGkX
1non4c5Yp0Bi0mg4vf1joskPMeQcxAHUJ2ugcUXuyBZDOvPiC9K93MSL2R4BE9o/
6OiuHXUOqq0m7db+qno2CLnVtzpWMGkzB0Eopv0OliGCJ8/3kaq8qW+p4b/thXVi
t/W4UI0CJSuksycLQ06ooDUovoVbhtUnfBC8lFhPVqscrTEo4qxd4+ehjJy9GMdY
E9Nb6OqsC/kohp8gwwUUBcbY1DAk4YlCVV5+omKsqxJOYaHhdD3YggAbd55LSAia
uInzs6CR5pO59EdLSKWE4bpb/4pmOAIM+JRoG5uyEF31Q39y0Lj4Pc3gFSlxisdJ
+BCOo900SsVx7Z9bHRDe4yqglVlS3j0sRFpa+FfGsUgV4jeu4sv5lrM/i2dqe8D1
Usr+JsbL+xI2hyl36yULTbdn0PbEDO8L7+Mkb+z0zYDHlNm1Ef51PPbTW2WonxtV
odJ2vPs6N/T/z1dcY4Ew+PmDSdRpY+r+NxYPcGCB+guGmEScOL+ClqH/gHalD+Sy
BW8eCAnhdPVzIYzRKqkL8Hq2bvkThUtaSCz4/6Db3GUqj/FtlvtYZmNXd/QsuX4H
i6b9ElCO/4/LAD5MFu62420CNWw7KJB/MlF3qmlu7sXsIPgv3mpTqTp+u2sCL0+j
4hLbad7H/Lb3D8xys+KuwnQGIg3gKgwMlwg1R4qD7PHe96oVSm738G2Y6JJ1tvvq
krtsNXnxGBZY8cfkTKryVGQu5Fo6axaG0l0iBwtOz+RmLB7mjatNXLmJDAbtHRTf
+Yz24frKhVGQMVkw5iIvOb8jd3fujJsZ1xuJsa1+WvX4uab6Qn/vVHv4MhnRBPwH
sk9qduGOuWuRPKNr8iJE6wDLqxX21JsD/N5cavCEXwC9y+3rufGT4ZcEbCKbWi0S
LG8Mg9AfPlW4zCM+T3RfuPxOo9ZD0gc6HLs4fCoptJMgFdDJETNFJQAo5QpF4GuS
rPuoOKjudQm1/VrTGn0cWc4ysTbEH2d4EXijPO3/pR/uWJAxEl2nJEXVOqyf86BZ
ZoY7uPSrknDKHwfZFo/p+E1HRhW4bMHQEHZJErJI2sFi6n0aTpqbEEL1Vx8LXqxE
BduosSZvI50xdSL4XkxLe1zZQ4N0kmJ9R2SMAnSYgmG59W2WWjwpPc0x52BZzdc8
kAu/oL5fz11ONfH9ZtkwKzOAUpMU42ZtfkbDITV/Ynp1l6wh9DqKBv6zysYJowM1
Z41MN/IE9yJ2doiMwwjlHBjQMFSeD4BuuzsT9mwDQ/UKRxHR7DKORx13DymEhZ+s
pbSVmRBCgRd4x3FF4c8pAhBHDRolVb0mDxoq3v4pU7vF4SX5Hk1ao9u+Z+IniVIM
d8BmcpAucAeMZIvMgtvfcI3zyasfz9a1nje0ryYuH7G6kiqXN8CAMV+7XJNN5xyq
/VqSaGrlE8UwoZhy+3v25CyJt2JzbcWq03ifIKtXvCgZvaiUVVw+0l/btEpdlihN
VO/UzTCGqb013fvkLMvlkwYwCotr8OnFs05QcGsObYf1/wsetc7XogvM/svBusR3
0cn24h38TjRziIiX4HUx/j2Z/I/m1grHHdEFGfMU6j2dxGN2dB+yvDUmW6S+oEmU
pTqDl6a3TfeggOGayoCen9JxJBzWSp7gXQBPrOmibd4MdpAAfpDaBOcZVaP/WerP
oJlaJp7++wRtIl+u0MAwN/8kXjho5tpvI4R08X1ebUqRsPBj2d2exYZ0IX5z/vGM
B9newGLUZkGX5ZzFkkHZlx9pRNFSYJmE1Kun3mmoOBTy0HMENEn76wH0kIFHxpI/
kGpNcZzs45RZ7qPo56nlc9NIKtg12uaiO/kODfVhGxXT/1Rt3p7S+pa0RQ2hpw3L
2AS/YzcXq4/W6qcWU1N3zQZyYT+CA6rHayJrf5oHBd/CRBmBILiViOKTPC67yiZa
gfVMfZFdcGtCmJ+nQhLq9QOQyfazefxlNVWMxGtiLXWmkb63TUGuK+ycPn+r+ZnT
Vtt2Ck1zvjl3MDFH6r1CR9TKwK0SI6N4Gn0KNr/ENPspbdBuzblS2wAI+Wt5nKSt
asyjEUcxn+x6gHMhoX9nZKTpEeAQ+uE9WzR/vRCyXtUPjPoYVoKDvZAi0ra0V8j/
mBkMP/98+GVS0B7SAudtophqMlWKVhaewiG4fdeBHaqF1SCalTZJq/hg7t7O39nd
76b42DuKqOaLNVSDzrU9NumUnHHgkaELGv7GmnMjoOep6cVXcFnMxDs52B7XYPzM
cSGav3L1hxeWyElGpEu3pdrm6jwmd+9eK2wUCFquheHPxn7aWSBLmCajjtE95PsP
j6soeXpfioNHC2Z8jBSmS0AY2Q6K3yxDnjAsEnn44/eXppkd7P127fecBBKONbz7
XaMSbV8mc8FHaKvkNTDvUa2SkD0ePr6zoSTR9N+L8wbytxQW0fCoJbEkriRUPalF
Pu4YzhichF+xbjDjUwJwhJtGmkL4u46E6Q0mXZ6kcuzSXMVy1NtrxD+DihfhYrvy
OZ/Vc6XxRQRa5M9GJRC1mlWk7GadoyKESpvVCyFXyuITIPZRoXkTBvilO4gaBNJj
63FUF7p71UZhvj06Oa/AU7/DCRWkbD/q/fweqLSvp1wDXns3K2kbwbOJo8AED+lq
2BcPpR+N06oeyJrGINmnUU1M3bpnczjxCYUL5K1cIwQhIwgqty/OQ/3PCVTKP9jW
Tkku7LpW2PqRq98koDun+T/xQ8Qt0ntHZjP2bOWRkaDMKXS+gY3TZHqKrsLosZ1A
anEH7kzXljZKcLmt7RkDehujBtdtI7WcecPKUEoja1aTGvFbivlnWu6BAtZkeceU
GzaP6xc38Fta8ZDM7EY/fuXSepabOucllFg/bYti/GSoTMPFKE/WzFl5i2rUVxNP
Qwas6eZCf/ProwAWsTHJ+OL/aQjPAaNsuHakPDW4YEc8m+S8WhlgBLI8M34KkauZ
MxXyHQLudMisk0sFb1Zm2IMz7Cvg9V+2S2vH+evJYbZtY85lstmYidU2us4tKcxA
J8G0NOwjCDBIhhNEZyi0oOnf5oLA0eRR932cmZk8sqYf6HzcTakBkUfGQP+hB76s
VlUlSQ0YLXxH1vtfwpVOur6+8Fjc0bCWakrbCxFDNzB7/aqaV2v4BFGkLsVPGRX/
t+KoTNi1n9PlkuvnZSH89uVi2Jy5oXqnVhDvMWk93b1RGMwgqOnQLgGd61HXGbdi
yVWRsgyC5s+JrSmZYShxgBTPfchSkKDorRZPa3cqwD67Qudw4QwLgG8FJfENjwhh
Fag/fozvAuEFeeF8bxMFGG0+MoTaemHm7vnf6hjUv1CIRea57RPtugAj5m4ZUfz+
FEa/ijAYHvuXDF8A11onMIuTtmgBy3eYORoAYOd5x/RT5hODOGg+QAwDyV+779RZ
u/zEWJ4Syep5X2b8O0IeD+h4h7Q1ggVB9w4UvibN/NHp9aHnHcRP7mEa5+yc5omB
9Bbuv1wOvW4j5SEsFr5PTEjKPxabdf9q9w59GVWCt/TLMaKgfvU0QuJeoAzQBq9q
e8a9quE9JPoZcpMdF+VzLZxiTM+2NuDr3uCwZIGJH+yEyojISCuEVv88LStvUJgW
MLjhK8adFLEQ3JKS/44PBp8v1Jsj+eDUXFd6fxpTYSgPqVaxM0MTgu12nExcGc8s
FMz9yle0Nk0dMmX0Qdpx17jJ+QV3WA6k9IIHhnGnkgtqhdvglq3jVrybiHVWwaZ6
z8XRMrPgUSHe6Qyj6OXUIo+4+PBsOEEYQUWhYd6XSrfn/GWqQZsREfUpq8VxxvDz
X9KhwcfeVpeqaUPrlhJQdIkFrfXFMBKYawyd9ouML5UHQzvZQkWqU1v60g9PQrGp
N292FjAx3zGTT+Fx7BlOtYVKWThYwxESS92Bp1F7a4YLBim3FrFVk/9aZgqOfWAj
ae5m6nHsWIbZqKbd1QyLqqPulvg+JuVyKSxcJJeOXQUPfdAn3FYHMHmFSKSGjk2F
bh/G2kifGWW1z2ZqK46lrbeJeR2WmRX5I7dfTRFcBqzgC5Y6rXK4EGY1ngutjcnT
5VVyerfT0xoYoUw0SFIOWJ9fbu/rdO/VYoWdSb5ltR6TWcr4Tg9nxBpwTxLnDr4M
0y2jLcWgGLslsXZfMUQ+darPVeJW9bmVYaOB+ENsfGrPs/qPjj4Gk4N6iTWwTwD9
ba98iqOTMBSgiloNaFgW/rsJ12pdI5Qe/o5pH6fBePJwkpw8Je3ZFvay8O71bY4w
S/5DhB1dHUmqFuh1VUlR6O286Cksn0nscqW6/A7YyC88p97KcnnK7nSSM0wJ3RdB
k4cP8QHlRX2ly6gg8O6U9nYj9tJ60I30B0kAwuGm35Uo2CJsqLzIcCTyHIghmUvC
cz48PBInROd89UPYfltF8Q0yP8jq6GK/z4XqT/zMhJlgRh5I7irNqKMHz2y+/Inu
fCNDHo/aPmhvSetgH8QbWlIXi4PByuzZ2/aHTtUa9+VaM/rzb4HtRnT55AYfT+YN
kJ/kPsDI/O3a0jSDRMge5B7nRVhARFJyzVx5UWKgXxMF8DUoWh6hX96gGKz2/wFr
CSWHR61sHGcZ8oxSca5cGSgKenfEZzA6Y+at96l5JGW6a2EbYXu6TCYIH7+0Bzcc
BRIaGmDAjZS6Gy2THkWf5cjcDyPRdrflxqLVZ+GnZAfBe0xM7eN/ZdWk5DCzVU3G
uSOTk9krYYFLzWT1ui2kQHGprPXzApn4z2wCAEpEutZcjb5S+MxREWUQCWmdfnbt
RNKy6i5jmSrmb8hVIqA8v+pK1DB+gJHXcgxYLXOcg4bq8ebquuDyM/KpvR9iWRiM
90iQw2vvFA31ftZNl9jgIDlAjOLHQPxQPU0jyOfZBvkKHxptBonlIjVAuIx3wpKV
s2HrpBP4RGg/9uvEGnrNUGPPd+DMOGFVSKAhZu8sc6qUodZTncmH872bbEtoE1qD
5HU/LVmvgPXdc73gxijB7h9O3sBormL+8E1D0ZZbQXdcbslTPn57FgdgQ6xAdOL7
zB24aVtFWvpMHzKHec6mGEzP/o15VIRfh+vqhp+c3DHJNnyFXRYG+a24airyfZV7
dtppwdecwyLRpl1hTakjoVrSYtgD9ajJLkskarO5QAxoWYiDJ4J2WeQrhw5dY1K5
+IGebO/EU+hk686kXe7QSAF4THHDHmvGMNUaz9r93/2L8gyDNHEYpO+7V49zhNty
+AWPUaSRP19YygcOAsvNNlcCuX2hVvhZ7fPjfayE+eT8ZhR9L91+0oQNkdxTYhYR
hWYFt5blaHc5FKW3Ufx8mo8Ngmobd4CpjD4UA0c7wcHHx+gUxFfjgE1EO3+YCElE
FezGSFGX68xdwLIsoduPO0KaJjhy0kU0mTIchV1AzXdbdcNt9YzHQSvThExAZkNs
pRre1ucAyROoBRSzertexnLY1DV8AS/6IZsB6Rup3DRNtT2e4ivxdVL0C7VBUHPY
tk0OEYM/3AebprEav6Exj4KUFm7IvCsRGCPSliuXqcTqQO+K46sXs4nwusTtIOg0
t6UkdMPNUGpX4NYh8KYBMciRpVAuZcG0MiMqGcE2UZyBj7K5+7kWpw5DRw4nf5JZ
AOYr8UXpkJfQm/IPJ8oN2nTcpHAnQIq9G9/i4298NFWTQnMZczbyGjRKwA8iFwjC
/vsGSowfmoJZPlWEI7jSyhZG9GGFmj1ymnCmZK2RxpLiyKwIUGuhoJF35rbzZPYm
SMIChJt6NYWZ7W1DpxusVGSkYJY//slZiCkA5j2eFknUoBarLwydpuEPwDCkPUct
HfqffH82Zhbjgjyw8Rw6stdmVY84l/BbGxoGrD5k5t4P1NYfa9cPcyMLkcx7t76q
39KE/ax16QodiaxUveUG00r3o+9KyVbNKS9Sq/0j+esXqGqXslWTUgK9V4pm+PyI
9t9kPIoz7d0DUGrWKfGD/YdsnHKnqoiXRqbyxjn73u6/14Bwc0jCxdFs6VNDxFdd
dFVgLItz5p5AQp/SgfFLERlqC1HE0Pd0KZ+N9EygB7GJmO9XW208O23i6jcKszYZ
2smp3HiMKV3XQ9LsFz/Wkpa5/1siZQS4p5w5h+7XDVTQGD9rBcFqY5wrNneLVz/4
7v14Rhc57zNPqrnFpFCQAlbkVqUzDgKElfk3+C3u/mBcfziJ2jWwS0uAEtWg3krP
lbwaD3iAhB1rfJDz62ZWtW59h98ko3TKF7ahsvat8JlyMnencRgQ5kLD4ZGnKTGm
4KiuN/FPBMwqveJ9KnhVyflnsyyelsfD/WKuzW3t0jmHWOK+Q7PlFHsGjw5cZirE
1vx9NcIzDP2bhSdA6bR4JfwEp3icjLue3W0y6Ym4zEXO0uD4xYIXLm/zeYWS5S5r
8hEeIcSgrDzG6myjToFMuozU8Hwmpejh76kBnbmvpexMMOTkVl3QFmdupkxmA7Ot
2RTl5bP+sNpAwNFS7YCoD1Dnhlkp3KPjYf1YLXZ9Lbm6km7ybTpdFGh1Nerv3zNL
2OW7NgAIcbAQE8yZ/eTFF0GjBgUA2P3nj2zb32pIbF7tA2KpGVdOLbRRR+TQdiM3
EfuC/54z3EUkLxR49SfEgZPsXLbU9X1XTTZFTsWFAOglYxF2YMo2SfSFju9gLM5Q
lQaGFFXIIk5cB8YR1ItGB5h7CtfEchKL0yR8NW5Aamy7uI6oGLnL8idADFVum6uT
JQtx8C8ldhYiVDQ3G+s1rNVxOhGlXuSuE3cjAREXU5iJ7/5Zzw71yFlFkCdr5vDM
U7iJN0tm3YF6PXVzN02ctUIsT4OhFGXIfm8Wpy5QSd/kKBZIV0RyU5MEWwHfkUHC
fdO+h1D0Fwu/yeRyeMth8j+Rapw5Gl0RYl4s4fd5XNkfxrmElxohTOAQ6odYEY7I
ShSDzUd9yMrgaFoc25xxht+TmWITODnSIfw8g/qfNNj+NorRXfoi+2S/h2kYne1q
2Bu95bPGhi1geid7Wo6FsgUwK850kpy4V/+oFwtJ6PjzkWsN+Es/3tgheU11EYuh
yGsWPc17hN2sOFOAp1BHBni6eAUEeKCzY62HmcKwcIGWd6/CEB+JVqLLSdYUxeFE
d++a9cs2AjS5Au08owrQuTNfdpbQq4P82Nh+c22Vs1EqWKcJDMidKtA+FpOdr2ZG
JpJoGUMavkmt3xgGnrHNAd8LIm74veu1v+7yMP37qCvb9zI/d6n3iEQGr7X7rIwt
115HdurF8yy6I0NczJM6BSZR2sfyCK8TyeG6zd/1kqgfurpcr4UQGZbKHfHos7kY
Od7Qsa+yxd+9nhZ3W7hXxhHHMmZqZ9xkk2Am1rQv0i6cBdc4iuVX6AZ/lGwUPTRu
FMEdTYhCjKfitbNYeowGifmp7pb9i0rS1IegvtB2XMLSWGU33ONEKrwj2pMDqIPj
JhjUNm7HSCsueUHZ7S0KdenFvC9KtiRsLPlX1QDFg3BtrTkCwrTg4kopj7vExsJw
zGXrmrSBENKLchtMBje2KanjKaB5PnyaiDEb+0tfDAVHGaXQ1M1/20ygX8cia6cP
a6pmlSkHvV94F3oEiiVDpQ7/ZsaX7lvg3ZfPfd8fNbEM37sKpWr6ifjc39AVkwqb
micbewbdY7YtoUH1DYIc01qQcYTrBbdwipIeh9exImMeBEahvCO/UiNgUoWNS1NB
/OxT5rz8gpms6dpFTqQMD/eHTcT2bZ5bZUAOy8A+LX3mvMPUyVlgsGd9VvdJkwde
Gn69DwTy6Yy7uh9RK/DlWcxCqe4Qiqygu/f9urSb1X1gdV8oo/Sn78L+HlTXUNi5
nHUIzMdnOaHtkIivc3sZBNaNlkcP5rCP+ZvBkbXLL7BiTHGElqWphDXiIhB7YB5S
YE4USnoqvG3VjFcQYEhR34WAVVt70dqMq0QC5Zetmus7zIrsPQyjvBM74isD6HKM
8VOw7bctDPprt2kriAMJXuNbkKpUqxXtF5eYR7SCwxvbnfEQQTY/ZfgjfeLzPf0D
Nt28zFOxQjHAi2tfISVKqcjbW+RErGcZHSaoOUe43YAhRaSKO5yWqfQd1vzFs8dF
otMszNjgEmn/PY1IQ3Oc7Tl0E1ZR8lHeJERCG3jlhnOK7l6AD49sYbo/6TPr8Phi
tm6J4m4ZtB5rhP9Y1thrLEal6EMSh3L6ZrkNTKgOHeSzEcLz6UqXGCTJ0sewsldw
tHf5bOqvRf63r44cvvAoFLVnJaf0qX5zClDqp8o3pospfI6TLy0UwLk0iIvhruCQ
Czz/DAYeT7DZMrQ6TJlUhsHB136WjYIzy1jY7MRmSM+ctjH0BW3Dfcxq621+V3AX
lIfVlEAguYoRJ1egy+xGLS1Ag1iDbyUxQhh6n1PyQjgWA2yxg0XtOu2Cs19NlA/D
wkJqfyl3bxNHF/0sW9MqqtyVJg+5WDF5naeqR2fr3roNZ8NbIrWDHZvOhvIOljnY
l/zo39p5kGm+rC+2Hn2GCH/QBd4YOWD8PYj+I07KfuY4Wx7FycJU8ddl6XE8yMDN
DC3YT/A6sim4ddAx5RBbg7iDK//BgmbcQqKVL7B3VgIZVeZ2poHqjoVAV8u/b370
O5dRJmlhhQ/G65vSxtpP1Kncslsor6ZNhTGpKiHhdFlFaHYF3BJit+ZgNW5YE1GB
FTdtyNkiVvoaSVEpVNaB3od44koLstKJoFIddSIYfJGCcUChcNfYYbuLBsj7iuBd
GG4aN9lmmnNVabqLdbiUGqPqwq8phx706UeKCj6gfI8SpilY1gM8O6DXSELz4rHR
ikbn7l+sYfdybbXLZPjPJJY/zLG+lgkh9TfsUo/b9pIBseBQYpMe+kfW47p4cyDP
ppq+9P1HsdkQajHLGHVfSS6IGimgTDfMAPfXmKXrpFVd5D9qVDZJ+G5VioWdApSX
dDx4a8ylv5aVgvCeX8RD+yBaOBa8w7ZakwC1aJSROHAWZR9SDU/sQpCOKa2roFBm
M6EU9DmNlFvy0UEhy2+6Cvt+Uvn5TYEB6fmwj3MMob0/njViep8THQPXuyee89fM
BkZo1B2F7H2oVDna484ZO2UB9VsY38jVbas1APHCY6nHCsARuVEq8VM7Dm+yF+ck
xhvCWD/g5CJjjy5BbBJfs9l5XsSaXTBIKrpBczMGmjrakEya07UWLoprYcY/o3rU
KlEJKa8EV2maFmPXijO8ya2BK2HkBuUQnFyRWjrz34lIjhe8pzh/KTO0uSBGsXbz
KLofD9yeODvu/MhkKIPcVPQ8D7ZFtPnxJaOBsU+S+13qiJmBCAMIgSwpAajgxo1r
jLweM8NUGM8/BHao0V91futLJxiS+83sQjog4Nq2O1J+bLyJts0zLzr/9IeP3bpm
wm6WVoCGRjdE210C5TdMOMPzm5ocRP6OiA4v4Tn66hMRHNksUuAqDLVoucsxjonF
FO+yym0J3E/nIuu8GC95FDiysvZkHUlLPTE5SbgQD0neMxhZXU8ViB6jSj0apFiw
r4KZQx7+YjLqtIYpE4hFhJ1l4Nnw//6RBZSKWZ1HAoMMmSfHYFr2F2PCm2kuHgug
2hLD4GnMC8tUvJEIDDWtBRQ4c34yF0QDFr5jxwMFIKrittMluHW95jb3Hz9v3T/O
ECi46wIGyttEZ4OLzLOkVQcCWjZrgv3g/FuXuKfmQ3QlhJH98v//+sfxPUivDeAr
ww82qr7OmccH4bQJq8N8lQIbaIh8HSV6LaAPik5140km3s+/qIDa5zsucrLZ9l7O
CdAjbtM2OPpJ3t16kaQB8A+a/iESQ5fmBfbjRVuL1uG+d8QNjiPZg+6nmXe/TvGD
5rk2l3ul7L4FxN6MMFycM2WMNuOcVuixDqDQVR/R4UhsqnzwAQnFgxFOUVop4gwp
4NqJ4fYABhZ0Ms+Uk0CpwJ6iFtXhbESmUObtl4vW2ZZ6Nv4MOKv9J2gVT4PTCz/w
RM6cXmFQrRT97Qc7ENwLMNY2bJWtGemvjpDkhwcyFvbWQWp+lQEuY7bA20cgJsN8
Yhf1aP7dBqcNkUFxoXBaGEPo5yBkm3TgQkpBfcgBse97p45lBf78yXVi6VfKGODF
EKzgr8OYJjRvdDgObP3QqkV/hUl8ZMq1OBp5GBoj1cIC3ttcIDIjSGyc42sIIxD4
oArK62lQoBrAOPxPIgIEnAChi0mVghLyLs5Lp6XmE15YPrXSK2VSUIoeGEjdfcYq
DKpiMPu+BRTU00zE4hN6eD31vbJc2eFe6XMnoewbXw4rN8hFeMonphNoYWdN3PQ5
UVEai5BusPvxHdHLU8FO/yu6KLYQ4cSy+f/fJdw1Fkd4EdbyYIOIkbi+koFSSMJS
wK6KFwEUqjgeyxRFgCkTNirF2zafzI7LWzaPEVSY3tVA7TTNueFn9w09aGfyTQqb
hcaYReXYTJxeDzrJSdx1rlOdHlBrTHukQMPUQzDjWXOkFUi/mxnBSLblSuCyPYvv
4q354AFEM2CO17oMkAWGwD3HOz62hrMYmTLbKY2fr0r20kRlIH6eFDSKVqWNzGVl
HVLyUd5Nbhyl6fCjmGQyFvSPxwqFrdNi2Tk8Rc4SIZyDobjZDAvhjHDhU7CqsE0c
d7FrNMdLtrYD7gaCy5u2jtBcWoE0/LCBXKwSrJDa6SqosoC5eYFH9V+6QMK+EEJW
HFA7m9VQ/2QU5+nsiKDlJpWx6d+qPsKb6Ip4+8DR945apBXKqmPaPzQtKDXz5973
lflO+YRfDK8i2s1dV0QJiIm4tR2qxyLsRPRWdkvT6+q7nfigFnylhLFo597gCfwY
eZYWubFcEXqec1WAenYwwaTMZiWhQYI5gRcM7vje6KXCVwIYn0q30neJcc8EFbVC
eFl7vmmVmuFbGlUmtQ6u78F/1KXEuYRfUnhg3LpBNBnlFpUNNYcOUNKVsVXyJWGo
7l1NgbtvwIuAnvCjnq5idNxZM2F5m6fm/222dpzd1Hfc/TSBTpcpYzXgeEUIPW+t
DRl6Qdfgf9xv4Nd9Gv1j/mUI3kv2NgikHH6oImFH+IBY5M20ARnREti2Zl9U5wSu
f56b6K8kOh8CZdLxNGLS7+B/NJwQe6wxUlT/MdNnL49aB/K4R9dd07On3YzTI0k1
VB5Jmj58GuB/zkvjqTM5yk70UwubGm2EmRUrClAYzGoYVgkc3J1PilOLpyiCApsd
6s7ejQGqfi6aY9fwCek/x0N6Wa4+EoJiGZMqZHFEpUBQj3/H+h6dg42DOUAt3g9k
PHuSsO5GfJPAHMlEUwH4J2hkRJXYFnZJr3SHiWnY787VkMyVnGbWF4HFCVJbNivi
jN01FP2Fup6LYU3ycOwR2eRTctEEyN9IA69ylbEpe+b/2y5PEEWtEnw3wAKWJV5Z
qUM+zFjnlmIiPLMdf2eumSBjq0dtRFQaUoUXAdbtiMLFXdNVutB9Zz6mCuXyMM4/
pLm+HAd4v716s82gFQh4LbEsS5wPz9lSCKu6RMe3KPoaFWPZLncNRkFoB4RzRcSp
L4VbMaODgcExKL1Cv7A9maG/I/Hm7PivyIRggDkBTq7Yfa1svGxhrUtDwGUuEwQs
CXPrVyH+6mkuWCjhS3K8TTh+ujsWr6FTQvSI7tmw1i1zuLaJGxfjzBIdQ8xUjVen
NAgaDgXgghvtwRgMjRNwB16kS4TDaWmOY12iP8KCYWHzh1rVBDXiTpIpektzYVxk
/b82LRQK9HrvTAazo2NdwOACX+ZfpaeEDcb/KLHY6uvM2OpL3KjMygXcnKg+5E0H
M0b48c7Kq1aLnVEaSaBv6TzVQdH0N+WV+uVKPu+6k8dVck283/XdhbXgBuniIp3x
i8pTpm2dLC5bi0fOmUn3DG9PKCV5R4vUQuhKK2cXV4dkmHW0KpHTaUJ1Kwk1mmOu
ukJ9URfuTrLSg6mYfbO/ueuABLwg1vNBjq/+e2e68obV/vgFfVTJEuVx5iYLgf+9
+z9wvTQZz0jvMxE+cjnQxG4pvv163c6pTIt+S0JXqBYNF4Kt6CRo1iLx8oCxPnrB
1cNUIGXnMUGArajD0wKdkRkwx5cRcloBsDA4H2F4bvhtAHZ+7YHOSqzCVJFMxz1g
ZC67gNqvxD5lRIeS01feaG9EJhwusV4LJHjibQMuqtEZHIIKe7QmaXNSwO1SqPJr
39e82wz8/tLGxnNS3k9PULCjciOE15tyx0AwWU5gUP8lk69TqYSpNcbT6DBED51y
laRV2o8s6nUPM846bzV+FcdADsQExjwCsp/LxvO49xm5MzlQso0wwQkdGEEYzvsS
FfyATT2HQXZxdAttdNnDVb0TG6/mdpASGsky/um015qC8pA02YMT6QUGW8iVOLTt
eDY+phiy6RAUWLW7CjCfo5RWfh6wYO/7yRe64yNVktzUU0UG6cHBCc2giyTV6SM9
H4T/oD+OwyR784ME5GpNDQywZWl5Rb5FAVE4obOwt6K/28cxOQSDxAZBkhFe1afI
pbxHS6xFF/d2i49uPvSRceansNS8d7XtbRiKVuBdWLOrgx0S9aweksYB8EK4DAY0
h4Ut7NKGCe9T6iTKRsdmcEYtG2jasy9KiXIjFZCtFeeZM7OvHIZeML0J/onJ0OVP
ygtZ6cbECv2GYfPOQENj6IgLCHRtAIbhF4vnUeP7ROrhaA+4+NEazxB4fVzAx6fQ
G0TKAjHlxMixw61eJwDCY2rYa52mXwV0CqGkxcCqkNoBlm51HTzbq60aY5ZMHcab
Ai+uPcR0701phWOXUWgz7tfC8Bb56OzezXUktzBqdkYsIRAzhKJ8YdRZxLl8ly+z
U4AdiCDFzYr84hlVLdQld7QSKTqO67Uct3wYwrg5zk68MmxwuG4aCKRaUR9ZjjQK
0nZLNdzJW/xmhcVYT+DnpLe2tV9Aojm1tvt6x7yLo4UH8p27bVeBg13KkjOpM0Yn
NU5Un2++6ogflRnXbacJyjqhBqC8gy0tSYkhCk9nE2HZE+qOz1n+2uVF3Co4appQ
GLxvjzi46bel/mkvRWATgyrPp07CVa1MJow+JgOmxM+3qs6VN++/sZRICiKv1Sc3
wxIk9U1JaCxwR9pV/DtVvyY6K7+muyxAXF/Z7wVDIiP6D9NTLUTTWu9SWIt7EHpW
3l+s9WHLxyyt6HphDa/oezsE0IIc3JuW4pFbqNDxa8UXExuq4Ho0DLJvhsyLCV/h
FkhHlmV9sxzUl2LYNp00UkXQRhiwbuIgohXz+cU+AwJ+p+V0iph6qGwB3ddUKbyt
vxu7XTAkRlHm6/dZsarbjdvpsO8jmBiwdaZG/codpbo+NPWB4p0imJxujI8xO+bz
dTcg5DrsIrC8je5okxTQWdpTj8ypc++sBgKoovCfz36gE8BuGGwTRvPod3YsCF6Z
aELSuuiUWLgrLVDBt9jfKdK/uwjqMuD+eVn3Gu9mPCReQfasEi9TdIA2gWD+jLt6
iKHYHBLRZjC58N6NYl/q0fjEPFkLW6p0uVLeRtV1ZrRHAUSLly4CWoK8XWmL6r5C
JwUot/nNS2lhFcS38w43ibnQyQHwcJhATmHjXMYj/fkGih7B3VeKuI1Vlo3uG9Ba
mXjLDJy094UsfoAAfBzoYLSAJ4gqAOHlwaMqS8SJqHkGVZYTv9IAKRk672QGz97Y
tj/ghFXDl1AfqQD09Ws/tGTt5A9p7S/OAWrtL12sZjjVXFqH0K/SA+qpOVNx/qYp
nATPBcoMgJKNsuYSelIFYwaAb0ZJgtmGL/0v54qQNL23U8orpH+D+LnWnU+pNOKn
kKavvvnYr6x6D50mTwLG7i8nXsjEjJpDiFes37MHAx+YdNhngZhDMeqbKfxXH3V0
RtmCfZb+ngWx7BoyTuEQCHJkYvc7L0cfAL/i3RPAT3RkXqf9tH33iNXwopTTzmIm
Fh1Yf+GoGWrpKZ/bwr1r7LZx8Twc04fFidC5G/9sNObqpJN4NHxUjwkHCsDBBWZv
vhyCiO3O+dWlUOe/CSd57lYA9Ib2wt9GT71Yd7PHS7udLS2SsCnhjsIz5r1TPXrq
ecTUW4JRPe0w7V5TCWKnzphftloop4ntO30ri49iEnMjsGRSDKiqZWZzvL25vNV+
llPA9yWnAffnLk66L3WNLRQoQaXdMRj+RJNd5qHLYlOKDALaT+zFbf789GyvqEtC
Ep2i+zhBtBRpOCvhqyXEVtNLTj/2LBNGOUHjCca3PUCDesmrn+YZ/56Xv+2uJZ76
f3ndHEDhml+Apeb8EgsMYvMv/7Z8X9goMrFFnDuzPt5xlLP62/HZ9XJW5q7xRUAH
zCE986LyUWvy9nsj+ByoZlrPEVBgqyaPI9lR6hQx4XZcsPy0Y8cO4riRyNIFNpJU
pFvyQN7I5EQWcUL7cJDrHjPfzChrfqCUx3VMicNDwezT3Fw5T8wwYihNVMygFAux
wYdNMA9EWYqNmMssr4X/q/cXbyEAmrQwMVgPSPbPV5HOGkeVXH/LTMCRZJBD6nKc
ROG/S2iWgD/BO+FeIctfUMx5csPl1VzvWnA2vk8Gtqyz1G2yClwPHmTsHUGv8xP0
TdOgrQyP/v4WzpPBvpiFdV4QXYiRfqiiLVKfd+wRaoUyMc1XyOTzn+iDE+7gpoGq
Jx6x9d5lWmvNUnHRF7HZ3SCzE2XJw7BWVmBaqzMODEwn9plY91/k+NY41tJ92CXa
Da5B943TcOMOOOXQVTNaYWKUUUnCW8kcpwNX4lFRqCypcgaESJ58XiSt26ezcWNu
lGCAYNIzruQ6qRxZyWrYvAfGngV3BZ0G2MCsNEwjSoxIDNALaViBVpTzmDKwuLUO
B4PLVoXpjiZWfKTJTIqoCblPqh1q86oD3RS4Mi70Rmrp5mNUn/qPSa0kd8ggqDN1
j6MkWjs8YYrCPXxGHVsEUlXGeEO2sc8TfQb5RTjCVHjTK4B6WEUrsKhI8A0gTNsW
BrL/G7QnRu4IdxH429Ck7hW9I7GtQkZTOYkFLh4zshOZ68gz+hcitSXSJRJZqQkD
rOCpkPInsLl/aVW4teza4oqvk5QNBlsI+hJc6ViJmcLrwE1qma0N83uMhRmkvbMe
cJ7NFgfiVZRC2SzSO/rGXlLokqObGZUjOYacqqOJjPUDP3jJ4uTb9Zv1X6eyUR6a
UOc+Cg8xoVoPH6xBiWka3VYlY05xrdMtixuJj1KIByy90MAIfMlppibJSCrFEs3V
qhtX6iUPNIWmhbaFAB4YbiuPAOHBIbV1PAtUGuMkn5/sskoYJa4l19BlSm17a4V1
yTRmcmairY21i/0H+iiSW/2DvdcJRPLumGS6NaUbTRV7hlCxBjOrKfZepyogDl97
ibi4WeUaeR6uvYfTZ/bb0QoNDMb0JnfplUCaWFo1RAVvtnLl0Fa5huiAH1f00uB/
qtATFXPeCcz8SzjRnVDXhW3GpaYz4PEI7wyHk8haFhsYr8uJPhlaiQvUSYDHZLbJ
RAXJGtnj/Fotfrnms3G8+z2U3GWqce9VbgloraqXsBxnMpiKHJ7MH4BH6CgRvm+4
5KsYu6SEC9SkXnqsmM5NjIZd3RqTp2vVWPnyr2Z/t4tIo5tRQsUyRAji9aI8P/ql
RyCibKj+t3dztk8VtwOOj2QfapQz9pDyVLDEAr88XLpCOFUs+NUq3n6ygBNiUnKa
54g+xxDGT7TtCEe9TatN1uKd3T3At6Kin84LYIHJDxkNBSJfI50Exm0orwBl4YwW
DMA+VHb/7ul96ylnwO4Uck+vUpV4WHP0zpBNEByqANnoKAa7vXkEXHx4ePPyGUH8
Uio49hZ15r8Q3Rfs/oNlImcG+TSsLlkvrvauZMfmZkRUmOvAdI7IR+14SEqNnhaK
ji6isLL+8uT28jcK48qcMuy/0cHFEFCppRvrjAoqc4ZFM9Wh47sr620tJE5TwrQ+
SSxwzkS3hAyKoeAAW7gzM2fkJULZEM8Dyf0ApJpDOl3XJjpdmdGYJ27rQxnom//j
pVm2uW0hEAoFIQyS8BwrXeD977b+XgEry93ZWIQHHuQKd5obsiCqDIhDzyBYRAfK
oRuec1nEWEKbUDH6Ep2SI6vpXPex3kqv2gPbSteXPjSUke8rnTnaCMTzjcASaIYE
M/bfewoFjJNlgd9jQVSn8FCzDCmBBbOkt5lToHa+x64VuVlrLphdc7hjXhYIhit4
3b+qQdHUbKhvHBhZljsxRjaDNs4qCJTh3ZfDnjF4uP4IB9ERvWzg8hp0bQink8L0
jAgfBG4faI0uYENmNESMmQFsew3aTISYVeQQv7xLOfShhw+eE4Pw0xS8Q93vUNUV
MCBedtreIl+2GQSdr+YA0O7bcYu21uvD99q6m4S+2h/CUuuUZjOFWTAda3COQ9nd
lg6RmM12C6od3u9Ztr65cE5t2F1Ibc7h3Ru6bHqvkM/HTt94RatNorwQaXHYca4y
Rbq5w2uPAsWXc/WG8ulq/uOnO1xCKPkUKHhrT2KsDsQkFikrAv3VAhMWzNxQArd9
BGpuNdqnBc5Y78avHAGYkhewZ5wJljSbN/xwGAmPLlq5YyzsQxairzElH+6Kum0d
hId3ReB2+NNZtThOL6QDvVwSMCczQhINTRMQ2dZa0duxC9JpDjm9pgMH5xf8AeK0
aZihUBrabOoksqUUoEcjnE5yWjsgNQmDE9oDwrcufDK1kNFU2lDBcKgDToTb6kZg
zSNqgcLQdf3gF/Kn3vniATowKDRQt4psuiXAIjrbIJ4CtUyAdA6Xb84PcfASDATC
h1CN62LpawcV4BunQZStjKVOo47Q1a0+cgwkyc62VJcVUOS7cmsZ0VRnUtQxpgwM
cRz7XnqL6OjYgpMe6G/YAMftQGG1Kgbvla+bWiepW8g4qrzHP4mF10TnU196GUa2
9v8+gFoDKHuYDwSfsDtbmGSwIlUgh/n/Ol12nwEqire1ZZSZ+jRn6z0DKNlRHeK8
FkNLyuGeUJyh4JZErZF2uTEKiKjCijBhC/Iiib5+JCRODGALHUDGIxmNxm8pCRxw
wQD6jfgvV1Y6YYNleVHlsWOVDd7Ij46hkmM8sa0Lyq+UyDd8hBc/RdfGSIfIye9J
vXF1pEdMKxbfiXcpkzYg2Eiysa8/AhYZVFX8pU8PpZEsRw5uzseDkm0tKiZhHcQn
dPsM5gORj/c/l9CBMClZt8YzqyieMU/fQPzZxAAmNQGBcdEpZqPk29JNQw7MdSnj
jCVR3UR7NyoO+03P66FaVjuF09XkK1CTJQ5ZxkT+Lu6g4OOKazRhnr4lbzPbNbgk
d36QTccdkPi3KaQpsdMDP5q1o9Hsa2UxTm/QMUB0+OBUgNlgqKQIfpjS6mvUe/jq
ZOAxnzeZbaYUNyPZ/tSHWVGtKYASIBpbZyRA9zST51rAe8P6HUeo3ZE0UXBWExQx
EviXlleqWvlQJizOprT628EGX9hyUTjNvgzrDYDJfvOwjVuVfQ3/uNMG4dGHpXKW
ooNvHAFGSkKYrmQclwHaZKZEB6/MbZ/dBtt7GUImYMupMjUN889YLSMfgIXWv+Mj
oxgzaGmQwBpFYTw7j+6SConZ/jLCjDV6b+l1MmlK8xHkiCpsolTW1kZ0oYDj0c22
SinRqNTkgNx/IVxpM8u10fcoZazA4G6nYexOFbWI9w0flz36Dz0C8TghGTGL8aU+
KMtS6jakCCMSxw7wxpJ/KhE2ZbhtoU6PuJoieV1WPwhvomaEV1cRDbU4dw589aa4
oj3uAMCuEeJv+B7YQ2NPmXdM/7vTDV7tD8MVxevF5r5l4P3skYTMIVv0BeKlkx7T
tW9Ot5vMRsIqD12L3dBR/FnEKuf8IRgFpow1XrILAzvKSi/CsliJHlB5+79BdrPj
/Xu9Hy+tqYNHjNQf8fzvctH4Zrz3twcjp/Jx2K7zfb1yfb89EEAmPhEp5/XVpinv
iT9W3YL/ZFX20jT6y9Jcuzv8Oeg1ipQu+TLfBDaEZbp2i23asSj5FqZzwp2ttZrD
fE/FiCF25pClEKJvxQ4fo0amy5sUR2zjbzBi2CCBFQXDvEGw4LOPP/Y5pzBB4Mog
Vq1a4oQeahuxCyXL+dKgW7GiVgm3BN857NoqT5i0/KlnYU2xqc7VfvGxqe/kcGcx
ASbCAN858fUhwklH+lEuDl0RzpkHFlSqmsG3aovtK02PvPEwFFbl/634Ry2ETmR9
jONFoFOxjgnp0Mh9zwYmdvIqd1tNQ8Gm/lS3Eze4iKS9cOxIDCNFxw1UcLw7ySFM
dax/pdUh/3YzU2vy3BGypwQg5EGdUOXMuR7//7Pm7QRUdGe/Z4FeFbYlEQVGg7ob
FJTrID+nDTSU5fjFt07egXN8ZBlAl8rKTzw3akxyQxn3XLrdNWY3HK9byVPXaKBq
25qzICy1L0iEukOzqb7dfdt2tTS+4RQQu0FyQf1emzAuAQGkRayn93VFjf9xmAhR
G392nYrwhNI70Mh+AhKVNoU8FCwlTHYGH5R5LjSqn8sclvhyWV5iQN4SNDl5zIJl
9U//2HmW3HOYZZ9SlXurZkagSzEDub4kL9uE6K/xS6P3bzlsvV9ds66BKsWmqgZ6
lPVCHMK53OztVs5eL0Ue6k0GeVwAb7EPcavAA2sD72FgBcYMVkyLTgs45FnCI65W
SqCDAKu0KJ1aOKABh4X3LR7c/1p52ATfWCTGpX/KTjjPugDRAkMG7sIiDEu+sJy4
9v3JGbC0bf6rzdKZMw1IzNPkQZ9+yqnuH+IX/b991O4Fcz5412CjB8YtsSyIlUeA
R9PW7qwxrXo+iY+njTMW5v1UXJMLpwi5a+iNhoxIGS/VcguDtmBV1hPIXwsE6gLO
WKZAz3Nbc3mWDPrQFWNspssk7O1eDIQJTjm8HhqP9+gbc6oOwfz4gzQb09WuSDlC
ex+I+YjacRxb3KeiJ95RkHM1NvTmX0EVK2URTYghdaomdsXpqC6AvPoFbsbaJUzo
hPfdX5gpEqu+YtAr7+g0+w9tNsxOoL86gDrP18wK6qTymD5IX+ptGSB3Yl2I984C
JRGU2AN2Toc+C/SBqkQ7AMtWAvWj/wTOgSb6bop9s3IG5S1vKBPWhAF8xZi2d3BZ
TjLz3SYRAg2s3pmrfvAw7SlbFDdYiDEHgTUiN3s8bMwNSPCcN3K1HtBdCBgzxB2w
sSTQw9choMicxY0B/N4J8mw/XFa35kps2I1SCjcl+RZ7ls9x+DCAkE1VTk4YrblE
AnYvW6u/T2AslSdI7BzQdnPpCq8TCe2Y02hNDq/Fy7hIAmbvkDc7O3HHFoK5AlKd
Pul3YSXCOgeFQhy+FN0Na2M/nRNDIValZiZRaN/Ntlp54cPlyrWqXgC8K3ISTTPf
yRZjA4K5NChNV3nWKwchQpU3Suku6l/XJbfSpgmAy5EV+eg1eWyQrSZ+bM8x6Q56
p4jitMYXScKi0ampxRHBQLHwgDk8ojniZ0oYaUFN7yGXoI+/3byhL8G9NXSeeOxq
vEIfwVCt+BKGb8ZwXWterlDcHBLvtsfiN7ps2Ek1fTupxBAIZwCrWe6XKhddH3Ym
6XHn7eY2YfiKFPqmrwtnQSuI85YutHcxUxx+9VbahvkYd9gd1frzDaWx+tDFJobF
iU2z7Z4CQqMGf+nVqWrobudyWarRe5dKpy4NUrGEqlc5ynMSvg+W/2K93CP409Al
zYF1gMaT0hgyxGCyT0YfdV7wIrzZbODLXpir510EU3CYNvP5Z9BTk+27jvyXZGTF
cOzD11fTLrSmxxp+gqR6EHMz0zxeuU40ZFGT+rC0hersJGkoRCa5nSdFTFKx8pI2
JDvMITxy2fUNMigm3SHiU8klw8m9wuXdEhX3qHdZeQn/cUbAYFgVKSJaKnia396Q
9qYAoj0z4wXlQgxBKIffp+CMkWCIeuvR5HT6babsk1ZEJb6C8lOsF3zWAA8JbyHA
Ei+dwwPlgwQ3UDQyx6Dlc3S0aQV1sQPUwJU0XkyUaTyUJP3G68d2XBIHrETo1Jfu
8wp5CcvV/xhtOIMjS04o8y+8OlOyU2lQlLf6IPELMh8PEgP29MtuJUcBTey8hAcX
ca9SaT6b3OL3t50n6UHhN7tfMC0MtiiTuI/l6aTAoZtNo0jpSekXsCsosZqkHm5H
s8zS0xF9m/pdCztubb3n+MNsLtoui3CQX4LKo+eUUUV4oDsEGbrubG2MKVHfdR+q
ufUh1Dwrg6u9+gCkaQLz3NWFoXOPY23vyOz2vKm4HMggirk80JEMGpRUk0xZpiMy
KHPJAfj9vHfkuxRM2pTCZw2gpewutW/SlksNFMQBBRbrkBGReRygnvwOa9ApZEb0
XNA6s3tWsDTj5a7T8uiHo5uQKWOYW3QADpq4FiDg7uPjD1+YyRwTbndL+0vE0Wd6
VJX7a52j8ASPjgOKyMAdh2RcraIAXwPIZrsa5UU91+B0RakVkmHg7vLyhU+pfyv0
aI/Tv1ZUaIQuBRiU6UsFEzIBY8H5+SF4OxaT6mDTtOR4U56Usd7OukfDajf1DTEX
2CI7B/S6Plpw52ljJu2gNbREllSFQyn/CuXAIVj4A5M+H70FlKz0Hi05NS3aq3kU
ayJjqOW8kOmeYofb694mbgd/6GMuNKTv/UhMvqn18JZ/Q6yU/iMVT0CxninIZrgB
yL4o26hvFuparsVOGcEYvVGs7g8+LQqAQ5DXW3qLmPwrEyFHBdHU3HU+Y3IHw9nj
fhWHpodk76x1x3UPsI4QM9x1b6oweABrLxD5Y3zcstZTtwW7zIHqk5jAZiRu6G+L
cvG7XAAAScHKrsmKaEmmGW7rVFoitYJidqxTqStyEyxAXjaZ02xDd8idUIhLLF6Z
aqm4nw7NDxG+3gEI6uIFIHXf623fQ8mdcj7Rj04p0mxKRQtUa8DAvbnV+oxTm150
AlBxGbEGQUSbyMAWTDzzjKxv+Sv+MO29NhVvrXYkWpNQGaSqRYb6tFWClcmUkInt
3ld5PzsMBXMBt/e/lcgycPG1c5vq+IxzRKYWmGqwNCVRPbNX5r/kwTcccd+ef+jq
23DztRnrpaf2+H47SQ01LekMNJo8/ptahvebba5ZaPrQ3Pl06goN3rgba9KzoFH9
g56niNncD4TFZorhqrzIoHrZ2TqmRKdOOXoXSh4/S3BFmGbJd4hLNoo8UZfDs5x5
r91vWGYN4UOKp2KJqs9n+HnnkY6D7EX5eEk4q2+SLnFXe36+wpyDSBMiBShmtFkw
YakpEw2pi4NQvXwNr59n+iikbJ505JC+VDoQ8NiJ25nTEX6GfJtm857W5LmMAtsW
V6e9/4bv1y/KFh0GriCIhlMrNbSua5naAB2yu2Ft77bCot1HcVfJMlMyXt9IcSPu
L08mAZanBGczEzhsTZg6T1KJvoN2cUXrDpNYrHKdzn5kvicyv0BoixECyrKRBX7q
DtAklKKHCVYp82MabmnmHSgS0A88PwjqywPRYnpkXmxsbmRbyO8E/z3I9I/4Wbij
ll8bHw265EjD9JVZq6MiehwfJ1Rl0Q/8z+HA1SG4KoLY4HuRU4YoMuygASx00uOM
h+Uan0+uP3SHeyPZZ6n9eyApXtIYOIw7EsQrDAp5909J0548/P7pvmXVCT0wga9j
zouw6S4S4aySqHprWnM+f9mjU7P089EKjhEw+4DCqw8pZFdegLVvfwMDpg/DzjrX
SGTYCu4ewZtKluohTKaRyfykKaHLYfhxFgl0syHC7I9z2gz+xgNJoldmJayjo6Ck
pXpw/3ugRCaFcwy02q1NMHD5l66rCn5/b5NYow3p3nPkeLvNaYHeS/ZN3lmnGmzd
tNfP8eDlelRQ9hcLx/EA23wwh8ypWH3myeJ1OCSZ4IP7lQDPNtfERabTAaxohRjC
gGx7g+kMB6DxtHWdtZalv6qvRePy+P9T61CmdzZdXLLVXFj/U5Yx/xEI14EQDgyY
RC0DX1bZfkt7TCrQ/i228yt2mLp477GJLhtTE3AnYy9yaqbHriGHxywH4xReYmdn
Jt6JUh/bQkLXwUrJopfpQm31yfh3DHekJMl9iLHrJ/JXfnOxOQE+7fSWnzyCHDoq
EnglGRzxtl4KAl2nlLgCIHTgIZ4fYDcorKYqJJX0Zmx8/NHZBDJIwncghk5C4nxW
miWHoeC9CJwLKVM5h2u4cT6twcmrFKIyA6Tll0Zwt5pdsS8wORH5SqNUueusiidn
+EEcidudbZliVNWTIW24jcU9hM6HmqmwMExvYQMrqwNNlb68k192i4I7igvATYTm
BJQaoNsmDtwh+ppAJxbbGPHASS0bSuP36DgmoQQgpreDKIH4wz2aOttON47/7Gw8
dzjRT3TfE2wRXZd8Bog3jJCgv2UvtiHf0J/wb1bKy+IFEFzUeWpmJlRMns5UlTpg
94tW8nJEyILmm9CjnbHaDcH/oiBG3EDcUJMQoSZ0Z0EZDYKd7waVXNIZkJQvZW0y
ZvqlFKbQGeaaTVT/nKMQ288rVx2hgb2lc1FlLFvlS93NbgrSnd+1unhDSWOxkDj4
HcSl+IoSuckGqZFM5vQGBt41ZUEqBPFTYTKKhfx5W6afBnZ671kxy3iqizpAOuJb
1hJ/wQGYwhXso97qxrs1SpwDgAolVGIA9T4lrfIvwj+BgrUBJeDJB1IYY1oD9s2w
oUM0S6DtfAv8XNoJGnZhDOts8vodExDUX+y7lHQBHbUs1FLRba8XxPIthwqfizKl
X2iRdiZUI8JG3K/jgt1QJ2OwXpGy6MAld03xtTAtg32mxGrDPzftxDUhAnOt5XYD
yin12e+PHPPAMZ9Kw/GjS65c61B7e1o4uwvmEfi9TyekiRQHznXNj2yFjgA6nJmZ
BGmqM4lakLNMyw9rq174jlawlaiyGysQ1RQbEFu0yvjAm1mXy7DKKN3MBuU8V/Km
TkXgROgyMpRuv1LOCKhHYkzfolgQy/pyMpTNtLXjxjAx4lb9rG+Xdyxw6hy8cvfM
dZ4nawDkWClfiMyQOQiKqBRyY5/ZXzJoDPVHZQegE/VbT5SJvlLrB3j7MxaVigwu
lrt/lX73iSxoRR1dYldjRnXE/NK27fx6F3PK6Esle+SczaaubGhne90hFWddeo62
BlFq+vsHvEzMnFWRAWY5E21+lsYv/RWz9WzkqMzHqJ332bhrRkjSoG+5/0q5d5kc
36Y5FlEBmDkvYOEXnJNPbXF58pX3Vc/1fMJa86jtzgH+GgbmfYSxZP8kzHDP3Koh
BNQUcBxfC0rS4+iUg87CchxfDw/FeMwKmX3h5+8O0zGXtIP1bPMMv6Qg4EbqaMHy
Sigp5gv6D4HVe1y8fqzlJBpljBkUAMT1HfhYbaZwZzGn3Opn3Nvwpe5JpM7xV6hm
`protect END_PROTECTED