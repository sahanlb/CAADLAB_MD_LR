-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
jKB3vcR/Kv9FTUfLilnK9Gu+L4exwI66leULSsnQx0O313gnuHKupntr2bYwEWAj
5bUuwtzCS9M7vVcjbT8MnwfoKWwhaXgeozwYbBh4shPknz7mAL7OutMhoKO/fNKB
TnvnJhxXtzcAzQ/FYrP89blAqJa6Ldezu/RkoF/6Xn5c1VpUsjVBKg==
--pragma protect end_key_block
--pragma protect digest_block
UaWfylBky0wa/QN+WL+MfSOlk9A=
--pragma protect end_digest_block
--pragma protect data_block
FpTFQw8LOvK/0zs00p6DON36OzaW5ecQP4VXfI3HZBlBDdtOaJXBDEirmbCGHNiZ
OPbNT/KnfCy5pQaP6bs76AHcMKzUGpNkPHXsmb8RBwIu1Z4xJWAwxyuIToOXGlGt
SMACYiORMZEdVDYiSIly0KaThYpF4ENHFJLXNqsWxFNgaCDC5MBTyFRTAvVKWG1I
MbJEfy7d8XQq8dn3f1JPo0P/u/hNMWp60vGkwv+K2IwXOpP1yzWHNUnt9kCNu2o+
yPdhGwtdSa79oedezxHq3eZsPRnPSOafxffrSAd/GzQciE8o7f1ElE5EoGrJE/A/
A66fXRMpP0cP6b9Edr+eUCG3DXTbbXu7CCfnVNBarcNqY6YoiPSRN5FTo6C/MdzX
WP3zwkengsQBnpWS1ZxPz/9J/VrY1DFcNqceS35YMRS5XkbE4kAGHHlkzJtjdXjy
Ox957VG5wmkka8j2JvwnVSPOGpS7hIj7A4yMAMjgqxqLFOfGPLsOKUlia4AYJxTL
REG8+ZD/eaaCF98lNaC4rkVqxPlWDdBNFd60jrGR+/9WRc6M/3A0fAToiKOme8kb
Qrilm7D6zN5ZzOudV+9O4Ztw5E/N6dak1DxFcqnYuYl1vlnLhVPfIHAo7JQAAf5y
aDGGgWtd+pYW0gmMoDtL0X/NKp3VrvaWb2wyMP/OjlYa1EOJXiZ1BghBAK9ZX+7s
Xtm0kf3eU9BEOvUy4cRVHDWzUns1aS+TDyl8jQztSbD3xcqITeAuRBBs1blRvOAY
NBmv1fyJ04yc+DjAElTELMnX1YcHV3KEju+22YWPO+6OgSBJ5z6kTqooNxAkXk6D
5kdLP+vcnwWlebzNSw4quAQHLWO3lhVgN/ZVAPztjqRAkizVWq5m2sv1gY0hbMTN
slvQ/rT42SG9qXd0W4KJ4Pfv6oSRnxSN/zmkAJoorJasT4X1frrky+TMhZ3fTaak
YW2Het9qAlN+QBlsW2wVpdlFSkBgLTuQlmXVOp7hi97/ay+is68nvc6HrcnsuXN3
Y3HNk1QiXslxRhFRJJCjM+T7gvhVs06YKkNfD03l+HRbc2XEYhLUP07uZ8FGtDyW
5baxPSR49ZxoPxM3CgH+enQ6AQHsQeT9f8nV7g6lmQ1e2pTp7g12CpI3pCHYPzbg
61yEgJKFWx2FzFh9pPtMYJ13q4HEKrAHkDganSsDvBoq/26KQwVkhBWQiv33s9l8
LOyEEvL2PaUj/1le7tHhvznCSfB+UxBgRyTFG/lIhxgP0VBWhMhazqx+zlukz6U0
1gEyHd3kmfsGQsqijri9gKTsctHl4AHWk2ykCoQ10FxK7tK3pxZex0Q8O5ieOM81
tuJogXeWJG9AlUSZG0TIe6kBRja0PO26QFdQy6Kmi4/x4diMjTYmS2ESkfkmS1qf
QWiPgk4F1/iSOuC+BZObEdZ1umQt9lMVyx8OS8vFEmEa7pahnlsDhFC/93s37mdV
KL8yhIdqq3WIj4F3oi9t2IUseqUUeIASxR/kkryNt2uzqhSamrrl0JtnLbhuf5yl
ZcoXygTConvXFJHXmvoKWqI1D91J/nqoQ4pz91oc9dHpnVDoxAG8DR/3fGj++zsu
V1krucm0JVe0qnNrmRuB222yXUBOS95KFh4bJ8GBVSwCYCyYlsR8/BqpCEPHjMpI
aNfB6HCAJwv6NARZlnTdM8lmk6perS3mShPbImQ9aSMkKoSa1HOXE1tBDvGwrCki
NG8MeeWSNKyzE19HQwLZ/QQ+0VzbgavyBpKEjnJku7wdIshcyo/YT9Z485ZUW/E2
M3dxLnn76jfoMO0l4qnDfbO5MrWAG6RRYDyuF6yW1jbW+UVazYwWARBX6lAk4Trh
kY4mfMBozwoDP21j6kckV9kpfJ1aneBPasSwdVxKw2s7FJmy4h01sIojaQbrQraS
xOnoloFAAuEfukkAjhFzWktPVqs+p0GUrJtNewNPZH/AtKgFsRFEGWhTILfDyX2A
wwvgd+yUoDEqGeUXzS1WeZVSQ8r8losZaL7wwCff47QPJC6/njx8nLDBSy4lLa7f
w8KSfqruW7s2MaKFvLGAMecumFzpACEZi7bBUy2W39GN37xvQEr1vaW8iinKA29L
cVTfzd7ShDj6LnTfiJjg2ajVvoy7pqtuGIs8RILBmyj6Kjp8oOsGCn9fWxclFwed
jVLnK301ZeKV9FocNhNQ8jcj/EIv79T7tgCdLFPPpT9GhLTD+3gLVqnLRKiiUngR
2KPRtlV9UsrSwS7/b3Ax7juB2gzTi6fTez4F8JaFGqHTdfd4Sr/jCfi1aLYz66rH
O3TU/39JuuJfmVI34VEDHjVtDZXWK5sw1NYskFqiv7PnKiKI24vCoSmDsVqw+V2g
ekKww4Fx8xu3CkNoFTROa04skISf7wZQm1e7rV93td5SFFzq3kPXMhyPCT24qN4b
S+ujUijRXCXlvDUy6Y+BYSFDJPLgzq+OWqE47MfF7Tj8EkKkp3eZKb2N8LauIEKp
23VO5UDGOrH2PCEt4KKiNnIdkJE9C8emxfyGaf1J0xqwADgxItf0GiNtRrCsSafD
Up2Y+nY6xX8vI9t3fbna9jxzjOB1tgRHDLKlW5yx9o6mHOMnxcC6daPHCCCA8qOI
OCE4ucEzGUi0zUTi3gh+1O44IzlqAo9TWtYSRwJfT5zQN2V8lLX2wnl95AJvkfWj
6DZAUHe3SFe2Mg8dsgyZj4z7TLbAWUU+EAL8Thiye1U6Ft/GI5sjqvbq0ZyflBuV
3/yvchZqvl8qrjL8uKpUdZaTaf2H7gvnka45tp8rK8vzKwhDLOIPJuYSF0L5CZ9a
3sLwuuh4vD9PQKcxU6PV528iNCvzeLuiK/tmXRhKXqNe+xzH6hyv4qh6sEXibKRH
Z9pl66VAjQmcQTFBLwjt6WlUM/cTWFuOyFwEd75d2dvXOwyaUZ/IOUHS2QoYDGGK
zP6n0bYgpmvBVXj2eAaZOlQluzB/ucpLVAgB7oFOlwyiHa0YVK24jD57qr/5WCt2
rEbn0pOMHc7b5PSHTCSHt272NcfesJ/gKibfOM3D18BUxhK2Q/WBu9hB4mpZ3NCi
lgZ79+1DSFNGR3lJsSazhygoUA9kGQ/ltAQRhVSH0JE9T0GD/WaT4Midf+cpiWmU
IQcwkBE/lm57yN/RR7CKyulynhgyugm3GHWXWBdzWm4Pp8mLZcNreve8tk/hhTw6
3JV6ov+bn8h5j3aHYYR8FLrs+NNrIAhoTgZwZ1QGBanQfVfxFiBaBIJiBMo7iMLU
FdkWcsGd74it9Wio7oWfYfR4dhMXc50K/fcxgs8LjlJt3LZ6Q4+4/MOZOB6e/6Bx
N8BJ1uTCy3lGkKKQldfG0QU8uRnl92Xp8a5knnw3eyU+EM95A2VRB+YuUqXfkUpG
gX0oWK9vMrwWsQBHoRm/pyKv0HW9jQcGsSbVVjTyvKFEm0FAKHIiyQVljCLhN5Zi
L2YjSslS7gmKG56vccL6pxunmmKsn9bB4DSzKCzEKMe1EEE4+hALtvOlZ8dtQfY1
5ayeALEp463a7WI5w2NiqdFrhVAAxQ2vXbjssFaPoHojVjy6mg+nqeMMZ2Fgcpo2
oYLjPe17J0hWqKEI+y3tYxrziDbCzgpffTLGor0nHrtO1u8He6FLawnz2PJz0UNe
9+1wKWxfq3GQDgPPDarXV7RZNeOnrbncOWOkjokNRlEKSnLAsFBC+VG3zXVNTfu5
s9IFT+Ak1Jfwx8vel7lomVa0x9ub3/RcVXp3+dG4B5zLSyf8cw0c6OUgg2XuJMLT
o8XE/xL7LNLPEMvmJASJ8xZA4fJCcqp8imwlhUlfdM5uyXFdhuqrVc4xE4RNfC/i
Irx/+zh4GcIJMemqI52wNdeaWebe+iSgC3dn9z1AKdRolVZ1ybERVw07EPX70x8a
Np/F0r6mQa9IN+GTV4AopvlL5/pioCn4t8VLY+yU95w2nz4dRZVc883vofzaBas0
JgJInLoWTIBZBE5OQXP/hjk/lapMktRIxP2ZOl7TaxosicX/kF8Lu1XbD9TkmnQv
VaozXJoSAnwF8aGSWuYVGo/xPf0iKOtlbZkcA8dh0CBORxk8f2z+JHU6sYRJQT+g
6lQ3v+JuGAB+BIfn8ex1E4cyA9o42ua6ZWAGiR0CV3WjLSQGTRIMlJ3Q7w9nM/ox
JoJEOI2KQTKJsJ2IqE2QAb9wnnXQIjWKlsi26SXBLLOVLTFd1uJ5phQZ/+NlunPg
gqQY2rVwVNMUE3hoiCyZhMpoxNsaVGTZ0PRBYGMGETvxfqpFqNMG+LvLW5fmHvxd
KNtHn2YQzG5PlHSzEODX7Z8uwvygkObGpJKsC8i6FlMkSJugVZ7Y1mwg0on+h1Dm
emrU3fT1ztTQ9gGkw7NXEKnEXDlU4dyjZWbh/QYVNzVVxYl7HwbyjolfYPGOihTd
c8+ysKnxGzGFgBFw2D73yczI9ql8HXWQiH2gfJdj+V+i0VKTqVM0NBGM8WWYtRAR
3UFc24n/Ouz6JR2aqG3er5VlWhk83ZMD5+7HaFiMMoSFhA0vZr0Pb69vmTiN60TS
M1cjIY9UmhUVwy+QRUI1ge8LApAeqouyPI/okTf39IaTFfLAMHYc2l5u7sy9eZby
adn7iE+Xb9VglYR8IOkXV3t+93f+Zgcl3jWdvfg2HnmhKU96Ej3VVd7P+XTKhb2r
jeJtpethXxJjMkfGbxxqyAWQp1kLTA1CDomx0M87I4IfaPP9zg3AzPxsK7EYnP3i
x6fwRTrn9n6rJnzgIJYuCrGWOJOpq1VNPz8NHBMYwlSSlcYcw7dUaJoachaYxIc6
NrqkzKxsSD05+I4h+tL+/ied+AkN/1Cbt6la1FQ8BAcMHVKNuWX4h+Fbv4N/pYS1
ShTUwup/E/YT2PiqMPxXzFnjQmExO/UwcDnuJFvr0p2gLHqynADGGOkUQQCKXOdG
UfoExz0RAXiQ+aikyLVJEvsr/+yl0XK9deca81r/wbNqNLXGj1EYLDzQGWKsOrLZ
juZ87lVZI44y9X5iq/ov4XdHrrJK4i672cQgLSJlCi6VnT9i9wezne2mtHO5VPgM
UMMifXyNA/NwgtPMu4UtUc0djnN/mCLrxDmCQu1A54srcPspCWBWVqsz79s4w4Cq
2hGBTLp6CZS3HsUz+UvHBjr3lP9FV0w8qAxKTNM3r8UIV8nzaIQpcnV8k+21duOP
VpNgqn87VFRaSdmsA2o5CWXA3lWc9GZA5wlnFMkU5ST3biKuOMbjVFwXn2RZpys0
dPdj1kffZoiiT3Z5tG6sjGriHkFfXJnIYH/LUO2VzGAdbBA+t+EvJHx3RXBgafLt
mYEbDQ1061Akh00R/hrFTNax3qSA4J0Wc99hsC4jn5am0/nzuG/jIvz2VjYq2DX6
V9nyuxCQoqRZx2tkm4fPwqwiumAVI9yzLZUUKsNuOH0iesO0n/rU82NwTcgmz5E/
vQzkqJqk1TMcp8MQeV3DK2pEpEumiWRy+Sd1VjwtsCrAiPmJ45R1vvqAWT0vx6Y+
fWfN+FLdueHxe42lTnFgrEwRxBiTE7oxyPh2xfqVRuvn8SG4wCnlflCOEg8sL7u2
1bfYt5bdEbbffoJf0upVqHBvbp680QAuhDWpfWBciKsqC3seI5BLFuFbZa/nFXhz
rtmLONzULZyzv3WabpAQ4wWJU2bhvdah4r7pqpMLzSs5XIrxpGNx2z9btlhRadak
z+rfJLtHhYz6ZYAa7Wk2NzyU7W8Wz6t12njTbRIaFQiDLRItyuousWTQMqoVXJ70
nIkGHCJ70afviVn+X3z9fA==
--pragma protect end_data_block
--pragma protect digest_block
P7vlnctW1UqvISoJexDh5bqO4Z0=
--pragma protect end_digest_block
--pragma protect end_protected
