-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
7CNwmYqWVqovz9wz+qMxy8GvlX1eNVI/GmEOTTC3p+//mCFW6Jbo8Q9v7LbJNmbn
Ks4UYD4SpWEaOIbKNufjDBvngBzoa5o9TIrTRf3XAsXcS9Z026Xgc1yBR/UqQE6O
mFS7HHuseYf1ng2s++Z/qOlJh0YPon5r0S1D+E1ku2uoDslUROJ1AQ==
--pragma protect end_key_block
--pragma protect digest_block
rUvcWMgn/dIYaPcxHRv6dJnDTDM=
--pragma protect end_digest_block
--pragma protect data_block
jnqSd0fBL+102T0II15A5Bdi0hqvv6LMRMdISfGTqn/nDuD3dxHr/rZC/FwtipH1
+aJU5A+/HT3K9wXUmUE8nZuMmqlzZBCbJpEb1fsWmYVwKzcJLVKyKPmO4tlfA120
VOaqqa7oQQPebEOiKoUXFkajG9oGK4oyRrf6TzDVXFqVrzXShhM/8LKJc9K0FhZZ
E+CROtWmvHOLE6kXmTW+6DcgWQlQ9TFaEp17iL0y8wl0z1Dc7beqKtMWnqq5unve
YyQG67aGuKiTnolObS4JGemcKUBALr1nGODkRziPVqyd4bbYIj3jFFCtkzRt3/Vo
yMZocrIGSZpS/Sixp5kI3CvlD2hR4gl0st5kWB8mjuWBeOZh6wt+zUMfGG5/KeJr
epy0y832dVqqXwAiWJ0E1cd4cwodbJ01Ifhl1Nsfud8H3c+oBZAqbZnb4qtncvWd
eTE07cENrA/vkMrWNpQWoXIPmBJVYAwej7t26Cz6AdXEKVjFOj2doM3wtx5yl8BO
42q0DmOYj/3oae9eEssqsW3vm6qOmRFXxRg60BRXkm5Rx+b6I+m8NUmdNsYs7Gge
Eb37zG304XjJJ4bScaWBTomjv/EEm8Cgo4cs5IojA9gRsSUQcpZ/uJcw5fIJXgP+
u0/FdersgWrIyKnV9z/adqT/+zIJu7wO9wAIeOqhh7oeWKwcfz7erVHhzXAPsTed
uwuBew3siR/XKC94eYGWZILuIMAEAkLbN0UdL72kiPBu+MYNNoTyisWu+0Qr4ypn
d3z9y2H3L4i/hMQP0D9Y0RFLOWzt/srOnfJzodQd4LuTf59wH5lbbls12q+9P+CQ
dp2xssZwJU8VAg6fyq2llqF4J09OrFTEwQavqKMS33vvdxtGumA1Bm6myzWErySX
B4W+PF7qF9hzugvir1+WB4efGowda0ptIrBUPWyy8qupFL6H/cuh6Xj5jcG3JgxM
h8bIaMYjLzZtN1Ad/ah2/cYH2tbR17zsigwdmWkQR5OmkRL099B6yPDcma5ee3F8
qQE3cbC7RTk6Qu12pzS3ipBR2iu+PSNBiTUdOPrRlzM7+YKyoq7w2KPaEfSbxd/i
abLOH//l4SSqOaf7MYW4rp5je+h/5g1wNH91nWoJUxNR+jFKFeie2XlQBygYmpgg
wJMCNxQ0zQrwJNFhJGqtuSXp7UCSOBSJ6lrnt5IArw6UlXva9GZrqHssU4gm688c
uFXpzo6Kxf4hMPIRRz6DfdRcpooLZkGH9ilF3uoeKVjdu9Za/uMuDv0/l6qUPdQb
TnUH+ANZ70nuYWQVrMJn0q+KL/vwx6g7dCCIinR/0evBklLs9lkebhLAfC3wfrfd
QQNleGNbEKxx3Z4l2HfIc3njiHYZuIYCtbIBloqEIeszqXttC72r8DbPErZ39ETo
gaOOXRsuUrR/ToRfDk6uDlt7SHiBdk8ENarFzuOzq7Jer3K+jmvK7DMZiZMQu6hp
MCNCzR7TC351nRMKB6jcLqPdvbDmahsFTrcekB1N5KMEmoL5fAgBzKTEXlFIAtmw
+jEvQKkMIq3kaYof9EkVoJTUZad5cm1IXCel2Psq5Ea397ZJBht6a04UX922HR+f
sENlVlCCzVg08adSY9PPe0N4s/w7E/WJtYp/e/cWqnvcurrgeUJ+Ep14tfJnJRi2
uXunPQ1YAGB4HrpGiz7unUl2CfdicQw5eaWgX8PntR+APFQd1Jq07yNU8Raeaf7F
iPcbRyfYOAR/I+V+2fN4hpWHyk12cZQtc4Yo+VjsmxTbdq1+7MuuEi1Fk12JfHOj
cfwiHj6cQVN6LjiLzLukvr8kvsWUjNiEdQfQm1PticGD/SkqG05mVyNd7QobNwHm
IAZlYO28wbf9msyHJ4jqCqwMX5S31EZEKwVN8I5xiqHSxoU1rdO9l4rv5eUymv+R
SnlofClmaeRHdeDRIINVHsATtUj3D/SJGGLckz2FpN39hqWCxW+zaBtGcnBqjSC5
ZhEK3smJEIp6rPFVIjcjox2KW1I5iONteQEhTXffKDLW0bK5GsHsHz5L0V2J0aOX
FQJ2MgngOu8Ih7FSQVNrmO6eGEoqDTLxJCCY/CY+/hiC9sguRpk3HPush0evrFSG
w/mywUADnF2H93QvNIAX+vgaGzRzu6csU8t+ebKH+f6UtmUeVBry7jOaWlHGOMc7
Kxv9yvwi/9GLLehuDlUwoL48fLxIkaqGrYiw9KUDkfwab8eI4QFxAc/HmOVt5gpA
jed7DHTV0hGbAWictnaTubvxRGCjImogYacaQXNLlISZ0KJy0+U29g8z2+m8PR4V
XDlk6TEP/jD12z139i/3DvE4kbuOc6zOtSKsWkUfnjjWm1ZzLT0WFVTVEC9fWfKA
x/CU+/NzKGvAWsx3Yl+QbwxfBJSxpNK+x+9hB2Sx8J345XyNaDvihP2Yg/pfFe1L
UxrKPNh870cbpD+pGRITdrl+C3tuK0q2ATU6vhivX5ZNEftvpH3LkI5aZlDI/K6L
M8Dkv0ggaQRzTMl/+BnfYSXYj6UQb+1PuRajHDqojVgvzhaJb5NH4kirOlAX6grr
s9SEuPA0fUcQcg51MgBP10adcCfmGx5fuAiMpPVwnN6kjuRRw+x+xys6cRZVrB78
ihuXxKeoNElZ+ym7FVS+x4CG26wTZac0xr19ySLosajYT3jgvBqLV2b/y/EfxiRS
PgUERM7EoYHRPkX/ZNaxCxlrK73090Qd4YD+uyhBwuOfu95tZY86xRRVMAW2Xb83
VaIGtSoglf3j4ltp/QUQAv5CaOjrGh+X8T/x95YXUegQrPP/NvHgSc37+X9DCUp2
8HwWL719pqybar1e3E+/mT++bQqN5zTEL+dQp7wQu0K+N5aVTEydJUNNaVuvL73h
Nz22IX3qxA0A9DzrBRebj+GkoERpzW5x4QnDuYX8xLAHbgsIgAQW2vVYYttzIBVP
JCT4s8kJHVrfaY0XxpjtYeaZy7I6r3xMygp2oNpVHx6IanxOjipYzBBHE8eB1Kmu
deLQh+0h4LjZ3OPSgDWDG7fPQ7PVd765sHoj1pEUKsm7yVn9H1DBTHaoih7bVVAE
Y5DcZJ4PBv1gy8YaJINWSJuaftjRl+T1VT8m4AXR7VDHrQdvCifod+VjkXNDenR7
P5iValp2oY3Y57IoBk6sODrXuhktNcvIV7CWLEEUlTBhGZ4kyY4DJY+gucd6oBwC
9E6QesJcMnA8St8z9vwajYaxKZ9Dv1HADHJM5i87yroQSSW/8atFNLclfD1OKGV8
VsG3U9AGX1q9p1bzZV4Caw3RhcDp93PAmXfq/XjX/7VlzpgE8J1+z7m8j/rNX8H8
UrUfI+hFk/cfeSC1jrK69NzGcomNNVNR/V5e0aU9THgiqDicsjLMDW86OyEJ/yWI
/wOCezjqK0fcAXTFJGGSrtV8JzUoAlegriV0awfz1lnlaQLv734wVb7UsSUconZu
GyFrGtPH9Srw6toqE9U3AHVfXL9bB3XPv8Ioyg4IDFjgGO0wBBotU/3pclgzjlZO
LNj2gIkJzzzUKDCUIIcMako1bi2FdoF8WtY3Wi0XhmJKI1rD2ibGohvmHV6397+Y
nvjaFmxgV3+ac+QQB+EcfoQ9Zpivs8hgbSB5avKFhuhHY0Iip/EZHtsyQOu04sRn
8Atgd7fFcjNAWrslAaCEY9ALU8i1zOMddKwsWwOOcuvMqVNZVO1JbXaFg7ok7xhG
AYqrCO8G9GO2/lmTxz9YyKaZHWHtG8ul6xdi5vElcLOMx7K796R0RqD6nVGwJgn0
l6pFGtRVGGYiM2CltuxSLRMjaUv61PM1YW19cP1bUUCDDD3JLWVe1Y8z8hEZjJoV
MF/qQlo/7Rz9KgSkA1T00nd+4dQZVl27gtAseQF9yVX0DN2g3YsZSvKT2wtQQpMZ
kx3q7paJRopSuVqOGlCBmyA+6WkjamVjVKcjkiYgHjWOHHYJ7bVhF3l/85mtnXeE
T1TiHbBnzHcrsYR1gsszmxTxXMtPF3U81PSVx6fvMuF7pXeOunqeIJK/LkMcZgVn
MDTPbqlcoYEsciyAvgbzJgVYNJGaGLlOzeEF6elaBkF/+D6DWnXhfwXdFR5BAyrB
94B0uZ0SDxiA6vO+F85eZ/MLJu0B5+LcowefAedLRDSQjqDNvKwSWB+7dG4Z81rk
/V1z0ofcHlfiBKqM12Z1TcKOUI54++W/0fFOKWw5ow/EMwdsg9hV/SiDAqVK8TNT
XAjXRP+sGiyT07jJOJGWXKosGgDU1JHw22c7Ot+vvZYSxB67yo8y5ACbFNtsZx+D
QXNMR/gtvsDNwDs9dbUdfgmXxJFT/X8t8GW3SpeGVWhfzWcnjODpm0Kbzt2qfadE
HpnZ8eafiopQZf7wSpEtAbGuOW3tk4ZydiGaqPJzde5UsjaryO5V3sBbJlC3W5mn
5CUtB3AuB/NKqx7LGkVhK7mn9mYiTIMxeO9YWk8VlX6pjDbo4RJgBWr3upGylkut
lYTWH23VDAbDx1y5BTWMS0Q2PYsFegGJ5kbEbCikaLIbm1w0roRgiAVNceYEyKcE
L6N7f+ef+toGM6knE/dzkgnxhwNELwBTpMij4LyrjfQw8/wMs+1XdHwHHJnB49no
LiDmekDtsmwwusi2ooWoYhQWzfXB+0Qx5u5IF2z6e9h18BlDIDIIJruSvfb0kwRo
n3ENEejF9WCq0cClInU9ceYcIaffav4rKbnQrjfeFW11I9JODlQLx1Qb8jO9TzqZ
77re6Pp4T6f+FyN5LenuAM8ErmldEp4CmlqRYAvzb6A1hD9nGEn7qsGgJCzISeBO
W5g5sJWZ22GSGiPxKggFZzwlCtzJn/ovSIuwEG5ck4COVHnNfD4+Q2gljHhNfOne
3gzyc3ho69YWX9VWxjDD8CVz6MBE95gZR8M64yIRZNV+Zqc/VybrvgVm5BTjzfoA
/36qr0832N2+Es4NJ9t4FHFh9MGGfviV+mBOd7D+L4kMUafUYR/FrG7Gj5Ya8KSx
plYkLI2MGjj+PfQ5P17i0tAxpw5BRtzjLl1whhi9GGnzzRPBi4AsXwNefCEfkizA
9Ic5aDPddsz47fJnDWgFGQsOZlYDtOcsCLsWjG4B/0TtrV8xtolfKfjkpd7x2na8
ytwXl7NSlLk5ZCNN0qWejyQrDHwkrq1SjuAyXR+cC/nvvXS8F5ojCrcCdoAbswmb
wdXGjFjweoSKj5w7qul53dmzBYgAI1ZLhkRYTBaZsOS+RfPRFCp4xSmTuCORDGwY
xtgz9FtSUvbCGbKoXwmna+28zPPHEB2E0jABpOQoq/fyFW9+vr8WwvCXgURCayHS
B8j/ZRzOvlFonl/ebZep8asm1GOIjId0x+FrSL1IxIE1S7JU+MEJvW/saQ68UgzK
HGoX0C2qHZNi+kynp2SUFBhSaY5JjRc8W7AdGcTol3crhzKvRjZdo6mBzIsZeqaI
8QGDWUYcsSjsbaf9YL3R6MphlIZH/KWmfQD4wbhze5gkA4D065+eBIqSo+cXDXlB
krv7kukNXika6/VVnU3h6KeDcLP+1M+7Gn5RW4Km7Jq0qku1Yw00ymG7lNLVA4yw
JTotvGZg6/q2iPZiVMMWkPCXvsN1mLJw7IM3iiwcfQMfywHD6Aq/+8no9cR20R3g
bzcNe+bVGTq/aBC+xLlp/QIgVSfyOKqvF08nDCfhO6KKWKVL4ftw1Zoh9JSfnKwO
6XacE6XHQGcEanm25GpyrndAuAZKblwxaUC9ojyltkGaME7nothZtzAvK6VQQwSd
aLU6xScj/S6jjkxX+8XKkQ1Bsl+Cl4yKNwnOciTCqlwP71nifz9KeLo3jhL9xcF9
F3nuvfdRiuYe0WQsj3hi9J46OLtPrfe00UPI0dob2wQCA4xD/TlK5kNZPUz8n16Q
yo5iHHa2yWi6K3zvC9xpGJfnDKUuToZopt+PUnKnY6n7H6Evo9xHXjUpf5curcA+
lciFGyUUxkT/BX2eZ0JJpei/LbMcDRKXkC2NiuH5WKGMi3oEE3wG3tbL1lf79JIg
xECgINUMndF/Hj578HbJ3kLyIDuZnJ2w97fdWJymJ4n27hpKJQxsPgTKlFW2loV+
VFI/fPtdq1fEKiQew9nOMvc09E1HtXoqR0D9loA6cLKEwx4Qlaz10mtfwGiPEHnD
39RJ5jyzSj2qq7ErlVENAYaqH6znc9jN7FIAZ/4MkKfsXN0MjW0d/QnkaS1wn5vt
QaRDuRWgvv0tW89Bn0KaB/AOSYv7jkZSuerd9FpgrUluPSx2qcHP5MV8Hr71BV14
I/DMTll3XQWyZKmUp/gR50rcVDQKUghLjScCQff+0o2p4BFmpfjtM9DG0/kSJiSQ
wo8il6ROmdcVrfY4eEWGVVYCjbB97tEpo7iGlsl/dxw0jGePY6Qr1EuRZKZf4lt3
GYGQrSbG05ZzAHYcE0QFaLBRjAnU2aqh8AMSdr3xd8RFA9cPKO9kNAeSXgic4bxM
EJzvMPlrIomip5TOnlZE39lnNZU+ndZxw49B0pf8KiKU71ZW+QhVNnnUfri2bDQ+
91CE8fWnXqebXpdmNEnlVuxIg3f3Kc5dCPaNJZiOXzk323EWV0eH81wFQxVJ7169
Vm2AneWF/pGip6Ca4JnD1XgFrUtyoB8qkF3Oe8CcwwO/6bdgpxl8e4XKXsKNq1P0
Co2IlwwJWmeSYKc4hwk+eONdqeNugCqFOxwRS9YO6wQGgJgxCnKSp3yQjR/PI1Us
kmRcpQLNsMD2vAZ/7HdKn268dw25elALY2FqWPP6Oo9MFV4Irw+lqtFluOqTO4Uj
0c+GW87NLc3ibK78HE4k+rDgbYcJbJR5R/8kbFgFkmR4hgqPONQCDOd2hXgTDT3U
yIwBJCLI669rDnqoaF6dcV15+hPA/0610s/JZOyF6pYWHLD0uwXHcStuHDYy8mcH
RYhfaGl7Cg+ERIWxHWvpw+BVR2An4ukhYGyrK/smUWUUAU6mX6+AG2pm0VC5XXzi
CXkBOmubrqsOYPvFsHyzeX7Cc35hZ8gC2xFHwBhcYoRvBlEYMLFlEAbzAvTWHMH7
RB+RRQn97mwqZ2SRMgbakMHEjlSYiEM2GximCHoT/ZyogypEY6NMyuiGyslf7ey7
xfR8EUBl+vb1FaQXskBp659ALwildEO0zqUQoxoplqq3QaE3klsrWYp/TfV3Twvq
jxJLRf0xwPPxsmHA60FkKvQqUuKKtrgDXzY39ARtxOhZFcJO3CPS9YIA8iKDAXfr
wXlzsiC3S40AGiyA8+Fa7fAuRyCwJf9mXQfxWPwtC1HY/rpRm6qfka+oLE1acu/3
cjhlQzCgCrO2+/p3CrdyMooz10rXRRfuJY8xoLfly3Sj/lVfzYQwcZcGHd6OiXL6
AjvIGtgO2kNDalkJnWQtncZFvE0L2WfOBiZ7STsk43bbs7bVFfQplicK1uuKfLcF
KCXkkBFWYnOfDbMZGLGQjMHjzCX2qiruwOKDfOBYZ4kk8OsFEWeDi7hQSA5prnM2
p5PGNbu4UnSFOPQ+A4bJKuxGBd3UwbRMkTXUp1qOPqyVpwfIL2qqysgrOXFb66OX
fRAMid5nTgD//lD5woxAuLtnoKIzkxXsNwIgzkxo6UxXUwVWuzO2IOUQAlFV/7UB
V9kNRaGQ9bB9sAyFgYLUQR3araIAzqvXi/l0dbaiBwgwcJ2HafeR2595Wvf3anCW
tQisibaoUisK58RqcJ9vLfCfNV1lfygucu8whY/FFwId4MWJ+qxthgx8owpT3xKb
BFdFztaE7+mrt+zu5j7V1KIuq1cdQD5hKk8Z6KsLOQuudMN5W3NEJs4HZLgythPe
Cc0WvpOydJmdFyJlx6/0y+oibymcd6IC/oXbYDqHMP3EQ7jEkCGOuC8Sjj/cgwsd
XZbAN6v4b7eCiQuS3oeasPO1xS6oM7Ip4ydOTtJePczqLKVuOepuQpfQQfjL5Wd3
z3sUu2yve3XX4RvtW9S1XdrO3OJbricHiDb2GY2hFzCS4K4ATdXgseQZL3WnEgyk
QpxviCSuBmVgV6qkWexBP5GubTklFCLgpPUJRo3kXsGeZm+Qik3D9ZV6EyO9pTVi
MjteHVoQiBbE/d9HW/uIVzINtX89FSJHgkRRzNj1ws+kD7SIFwYIdNjAtVNC92Ib
vpbEYpJ73NyV8tD8aIqaGBLnZxoZnu13wQHk9k+mAXH+S5/kxHuwjJfHQvGCbKs2
khhCEkCUzLvUUv7dLAX1FJUthOe4n/yWi+7bWuyvFBYfn6UD/8XtWh6RF5fRZxiW
PjTchrRcN/fepl0HtjD3nB6D6eDioC1pkvZfBF2VYWE/0ryTno30OHHhj2T762Gh
1jVxLM9kH8xmK3Clup8c4oxPntM/M7apKz3Yem6DlwNYJetzcxn7K0f2rUlMsWS9
wIsxxNGU+rYf24Jh9f51XNTef549M5q+1DAXt5dRoXSN0DD6asYI3QYn9QprVwgJ
eLOeHR6xC1AkK4VRsmXwxsZrW/JQTioGPRbOMJgdOxS/SV4nO1I0Q4dMgn4S1Wjz
VkaEg4luEiaQs/BycyLJspaoE9omidi6nfd+3eH6AYQJGMvzVYdO46hI2D9zpkQu
hPkyCs62UXey20/4WlvEV6RpVehuMw0iR8qB6QybVv7fkd3DvbPJEcDstF0y7rZl
RIB13a03KwA2J/yB6yQzI/lZw7HXhh8A6SBoOIaaYnoMudUy2JVuF10xIt5mgoO3
KsH4yH83dPX2wkhIABK7CX+ucxaXvdCPBW1GzJm8E6ems3hgmIIgdSloH91hF46e
GqUQULOkK4n1VmKTlAtV/PawToK62/IBXgZyURGzoCokNnMreNivtKP08KnZeVqb
sOVCYyO5w54tWpuMi6JsqzgYXMcx0arHPxVI8tzKagNLgsJ0/VqpeSRWH4BGcQDo
wiCM/vzgs7OBGtVts/mwUyheWp9D557DoW67wR7KHBGEnUQP8oXcixuUw84mXjuk
FimsiFqFo0n69QSprRQRXj6ojRUgQvt+ozTSKFCpDOon2FBt8Tp636g2bpM/fmsi
zHAwWfDZa00vWIjjkUQupmf7uPBT/HaZ3yvoxWgqsUb7HMoox15TDSg4k/K1RxGO
C5NKCf5yjtijxKKRLyHy8dok7/NzAdAPlOEH6JKwHzIhIX912/wdQtDXXpru+5YP
VCMnKBJ2VhoQr+VVlSDTI0Ccv2HrCPwIToIrNu2yTeCrjcHHa8n8kfmGYJvueXov
nkPqH0RQgcVwOdaThpHEojwfuabM9l+2jynfaESGJxndDygNJcdd4E1xQGAmPKWt
U2qTYObuSQ1zvEcNSv27dyCAwZvnkx15MOxvYQwCL26OL6FpuDt4ptumTm9wN6nF
hi0FxP1Mg0XLzXNJPdk05+5I6b2fYgrSdsynybtbeE4fOq92cG9faFsySKpgCAdk
YS0u7oCWCIFnfm3Jw/OO+PjcNe2j94hsCd6RuEN9vFdLp6kiT4hiVtA8nPA0ED3f
CnyjX+nKVguo/aylfY0MctV30iRaShW3xc5XHJI9hV8Ws7NRwEc7FLCvUWwZOT5J
XSiQv5vPcYJwnBW7gBDAAf9BtK59ZDBfC5jiOX01Jy8YMfcgRFBK+qB6qOswkzb0
arMgUZy8Y3hDNSgCVbEphtc1+qJrDS35Q3o+uKviNpfCmngIginppJfvQ+Smh72A
IflhnRy93iwD38OHaf42jthUZcOOZyg8k11ObjQoBXvjMSpyiO+mYHQDsSxff9j5
Raa7fMr72wAWhjRjTScL0IX4wKp/1RQzpHrOkXwylm/yI73lDX8Rl/RWBXFT7DVc
0TSltUCux8g6w54Polozh7kViLsxE0DsN9BD1krzDD5nAp29+XXH8yq7FPiLgWbz
FuzW2FNhqofe7iZf1/ZGiifVUYB4UahEyvCIXPjlDRCHYBD7jgaLXPhWyP7+C9YI
W5APPkuxoFOdVCuZfFF5c6E0zDzJYMVQ21RQQr2jmVlyav0fpzWgUJYZ/Niiu3V2
NovG45qFuT00/g6IfwUk58Xu3ivTYDNtyk7capMU+SDMcwE+wf0WByGTuvmPf+tJ
pnCB6GT4O6z156Y6lWwR4TXa4voJEs7A2QN1umzFtMHYj9DceVUk/bvr2XC0hyzt
KTBcnqFOBEu8LFHNzRytwS66R5s8Y7w3lB6L+nuqOtdd5rQt4BGthyjGbBzAAcfO
WKsm6hq+X8jSRUyL+iwXjA+lfGI3GgWX4jdhzl+xg4+K/BuCBVFps/rEAuPUNxXs
HI80HK2omk0XsoIHvdDTSJxQ/5XGonqw9OE04VmgFd9oxBhk9PxuNNu4AQV7FDvA
UY+vM57kQUKW5v5BCUwkRlO1QqROOr8ZS5z41xeFWv7VVEZm+q0ddTRHbyxC1C9U
/GJACOxXg7t+WGixhs/qHrzKlrotkGdklZ0JXkyfKxMJ8d81qVpEIEJwSefWmpDD
C35sWeFsF+Ws4kdytW/9RtlRY+i9n7bG2tHiANwAJIyoCo5QyeCkqvp21rggUa9A
oyXfJKdWZye3eY5xaRMCRI5JqsjIHuncwoZys+o2EbawjhPzFTE4gd7aruFvodAR
Icyww7twqbOkaqM8rD2nm06Lhdxoui34gspbNnbNIWVNZb/RJFEctrGUGkRfPVui
RpNb0vrsYRQML2AvGodrVE0ZNK6imvs4pBUQ/+mgCv7/t/bQpVHXr15qNpXeFEQa
0bdPdcYocGyEGYRcuDwc+ygEoT3T/IJ2VqnbPVBI/553j8zpvnj5gDss4EvhBWjQ
RXyJGUS9qnExnBCZHhqIVtSG0uqgZvkqt08ZBvZ5oG/MJ+2Mb8OCE9zABL/0io+p
hIsegEMygK9rde51mdskrBL5IB5D5rms2LiOXEfc3+XLH9DlRluVS2ZYBhd8cj8C
eoscvq1V0mbMSmI655CRTiWBaJ2w4Kd7BrgoX0wU8NLzWbBsad4yBTQP4L40yOj3
KldcLGqICqvg8H9zVuhb0MLFMEu71D+8egsXsLU8Udi1vUzdQubnSrYnEAstqSZH
VwFyYnEsv0M1+HR2IrkyrVzFa5iqXlwB0rW9pOqHtPFwi7yGsIsKEQe9QGoyDFKt
D0y3J2Cm8oQyBIVBqa/2/XmhGahAx4TG6DD68fbdfA6OAgdgt6sKz9MrHwRlDlZf
gAuJgso4bI6V5zDh0SlmjuaJjkjVIAe9MoIp5JDJjLlXIjA/44ZN/aPAreXexBlw
lQn2IUG1XFLnMABipjr86J0oARsW04TLQNQC4Cb8ZcPgiRilrOuG5+jLE0Mi/pR0
hD1EEVOwKbhwmKXNrXQDITekpHlXEVkuUhvVUpfGgGc1x9Q1N3CVJNldJJXbnRQI
lQsPYVaoiH0e9WodmDVYVpgx6MAJT5UeVMW1DSL9l2+du+uqnDzGi5JTOjQyV7cH
tzbMjWXq+8jh73+2YIYn+8KKJkfjspp0Ub2VWOlnWvkwKw21HDP04ghFfYShte/p
/v4qQGkyCjvyvJCAfIcVnmOrbrtabQm4RoJC3Fmmxq3115UWTnaeNeR33ymZ09Se
cKmzZd0ILvdLlav+UswLzahcQw7haV2KbnGDckDA1Et4LIcfn/QSv8ukKguxZL0e
xHPh5Xd2p3//7DxTkCy2hlwctuKi6qdeuVuX2IRoA5EZCXFmNoRn4CTrvxeePwuE
HuaE5w4vyvJnlZi2zxZVcYZV51LVkSnQiMNQdibEtNz05y3NWVjroaKZto3KSR5a
tTqBx+M9foJZA+1QecmfNyJw4/PTb4euufnA7KB3i6JizAD/Za/9GRFTL0/OfhoN
3+fbs6a/F5Ru/lr5f9jxDs8tX1VtCD7sUNRmhSWVPOI23VfJhe3izwgKh1NpPpKh
20APWz2JLAg5rsvYMu3EH5MJA7fDCQ4rnok7UASyGaEve6ZSi9lS6VwiS79diGiN
vD7WLwBIvba+vaO4fgvg2sA3xDvqDQHLncuwwPEf3M53EYIpI3EJQXhYaW7IuDEv
QsDxeHhtdybIrR1cqWk27JoZe/twAxB5ztoF18ZRYHc4DCc3sCpY1fdrqlhuRsTq
GZYL/ieS+k10+hWP9Vjp89PSox966XubOLjigfNS7W0iwmO2OYgzHnr7smunjPF3
v/iU8qIuP4S1ehz2h5sl7vmQLN5A2oaS1WgX/6SOEkarnh2koal++hnYguOYDp0C
K970ITWk8BklIvhHinkTIqMJrcLRbI+1wR5sKHXbxO2UFaL8hDeXwy8FEZ5KKiyB
sDBhO6jqGeTqB2xhShImEvDXGBOl2f81/54lGPhGkt7YOKdzTZRGf0XKo8S8Q7Nu
CTy6R7bOZu39bViZz4PqNyk0iMERldl4e9APUDEi+PLO4dV8pFwGvrzW0xzmJUST
32gtfIiQ2YAbeQHZKW/c9GDXosLUj1ixJu43ZrA4SBO6/qBIUcIvfYcvcx2fszNk
qGptIyQtNX40iGiQ0pJLZPasHDWP85d50M0uMs+t/g2gQK4xrrMv5qo56VLm/btc
FfURgMCb+w5OaKDC5RaqX6B755YgTKCBA5tpk/RIGw08Ttya6Q+gTdvEKmAGeXKK
GSUJhPOGY3bB9bM/IdwPWLt0s3H7or66eTchOLCZBdUSCl2RPHpZ9tQkUgAHGuXy
GHhKtTGCDco3FIgQPsKyVsgCRPPHTAI5aJQ/qRdpW9ADXCq6b80/CBaQDJCj+q4Y
oPQAryFxQw+qVvLyL3dU7M+M2FFsnF/M0YeX44LTcWhXTa0PPvK9hKVgvMkEL9rn
nYPUGBmx8ttpRAtFxzXcDYf8RUDzr1c4lwgrifdOnMpCystRbt4Eh5aqevpeoTMV
2aPhZCMxxsF1qoxvQuTo3rRQURMKpCAdhfNNv1u3lvsqbDiojvRO965tcdzbvpMo
tmf0fOXkQSk8IaaH0CiMl7/G+mctC1Tx8PllTpyn5PiNm/XGO5csABGlGJhs+im5
5EEmcp/mfoR62Hmr6KSJYuhnL9k67eJKCzEPIf1LvE8NJ51A0c1fKBkq/rE2qeDK
KiQuvniEFPpc47q22SmzEKBuayQnTbIu/dpd0dYrNUyS6LlIiJtnLVeQXHa1CLjW
J5/J3i1X2FQgiMC9mBSfuf5ZfNYFQM5XMltMgkg7WM+XR5JQHAtZ6+FcFYLsn+xz
7t7nF4brRGUYuPTXaoxVql4XraqRD7+4R9Hg3uTZRIlHvox6V02Gz3Z3nOJbddC/
cIpxGA8cldCHxx1gsJKPNht8tmq7wifmHs+VZ+y3HxuuCHAPMT0AojMQsAL690GQ
O4kgc9WcgLJKC9nyCIK1YtFfxKgwQ84zf1r3w9TvO7O2qPY59kCHiVxMCCuso45q
wNGtx19o8YbLB6Gc/tHYm7nRk0rAF9kymH6zYl+uq7qwGtO2/OMTqsZvVJd16oP1
LB+N73djr+WvNj9wblDayeYV1aaKeFgcqe5lmA3TCfmVuq61SuwWw/XbaDGGL+xR
JQ09XBxAVq+fCvoc1aNF+R/Y2SyWrXPJpnqGzbmmq9mx6/tySVKad5Hlh6uMVB3I
7NbpoilrvU4loq/UaQw37fcIL7gwRBP332s8o2n4Y4drJBI6BBGnBF+R3VLl4gAq
zg3fLXfsqpJ2FSL2fXgjwtKojjZWYM+nIYH88EWKKHdDaK9gsK3U/XHLJr8e+E0H
awzSIE3bo0h7dfOerWbpm1cU1nDAmwYYzw3FhKzWXq8Fr3hVRJ+zIxDvccDJYgqL
YyKDkToYV0VHb6CcYlwty/rOfIn0NuShhQ8EJM7zbooI7F1c7OazxHervk0Hgu0S
uMuvIjQQsfrVDEHJVfCJnytMdmUrUeN1zOvFyUafDPUPyRdrT7N3npRV67Ke9Sip
C78Utzx/vkhkqKEv9ag2JtdEtZeqofTZtpO3s+Wfq+CWOqB9XZvemPPPxkFxRfp7
xrcA/6ulOV4oEZe1zIlau2n8jfXnIiLvUnxOU2aBLcWBwe0Mfic61ZSv+R0ER/U6
90FW8a/A7faRfMxiN8Y0aH5+nJZzSdechYvqhzpshmn1NEJQ3ZxxPyHVOG+zjQ3Y
8g6B1cCFtyNFF8otg9/7YvLPnOIUfVYtMVxOhFlbJV9duSfl6lPIAGOXGVwbi8dy
WhVg9Py8sGo7SL6r5olH0a5skyqCPzdPC9b1ku1+8FaF0qyrwSilSMFliHnggoRD
9uGyaI3zjzdgHveFCrh4H9LgYnT1COQVptpXICuLSpzfTDiRDrk142QoU+77SFUr
fsFO1dH0V1bKHiBfQ8ZvP9/xqOpkMKB321s05vHXmE1/t1VCr8dzB2OFDq/vlV3b
Bj04VcN6eO+3B/Z8s9cihnXq8tWhnUf+ncPPmFvVZKhSt7TD1CPXqb4yMJmBnCo6
0U/SVcYqbHyWMNmMr2ei2LdeuFvn+oHlXtTUwXSm63Y9Ca6aLX8Lzg+2jsg/R/ZK
mbrLVdrN0hXPShjJVgqFpi0TROF4aeMGe12OQVHZYPz425Koo/c5j4SlyUQpopry
a1VtAVUVtsCysTfn0Wf4HHKyAPDsHd7rFSm37FH8Uk7gk8p78gXk/NZEUrXH8tof
W8RkLUk5s+vYJvrxYtl2Rh36Dy629c4wwPwEcEFjKAs+je/xnjUgk7vHLu3BklrA
6e7XBPwWb4vZgDsLAelwc8sPX/riOY5zSg+9LlYNdKGAoujVsZzXmIv4mzp39ZXN
Ws8a3nGT/eqM4fCOocCU4k8dJ/vtk95lAYaYEf23RrI/MPs0E3Mme6EG93JXEAa5
twIJpr/DH0wAU5XlGJJ3d9iHJZ3cqRZb/NFZ3IMG00GGLa6gco6t//wUQ0ZrZkHe
rPZE7nRaSlzjX3KPmnAoRNTiniR6rqPe7BVKnHFWBQoKEGbvKqyzxZVHE7j2LtxK
T7XltwP5YDbkkSjgcH+6IdvxynUFFxxlt7ITNDoWjbmL/g1V9U2//K/j6uPNNYT4
1ACzJM7+RGCCzHIypO5RWYo4YA894kC5BF/oLPlPYo1e9jfcAjcEud1Dr4DLSIsd
3vS2ktukIEWqf88xulqw+cq8uuprAWTsVFxSdP/3hckk2oap+aZv/oERQsCLQMWQ
aMKkkM5pp8eBnRbyeW0KTd60nEq5gCMfHADc+VzapRA32lhY4ZIby1FD0JqhSa0Y
k+ry+0jprE998oqnt/actIKGkYbaJHeWBcN0ICA7yqiGNKSU1iHM+Zd7OvQOVG3O
Y1lmfEsm7c4ldzYenSp2QmCWTvvhZ+NygTvbfqgGkckfAPqvkOnIFmk6jpZvTHro
m6nCiy8VBr7aTom57egjmbPmI0P205+/kWR/u7mje+wEV0cLjY8bdO3s6AppTIL6
lS6M0uLrMg8a06RLcqaHvw/JapilmbK3N8DNI+zq7UcTwlYZ8m42fgSVn5qZ6+LT
7CQ8V6g8K0UiwuwVY2R4jfW8Q6MfEpFzuHTd3BIa2q6re5yyUnCdSwqPtsOyZ/bE
Dg3W4OxPYEIQGwrYtqkqF2PXaE82wvdG07tV50rMi1fYkCBpQFuA82jCJ+fTt8Uq
M9mQXOo8CoynKtJItEbR77wSRoJU2xc2nnVLBzHH2z5FOdbMYtO55HB3Q011z2d9
4nHMvfC15i7fM+kNVb4hRuo6BEvEssP0EBMsItJu4Ot23iGr7idaAxwqwEuW+QJo
VWdhTNlPPtzkLooNd6NGk1IMcg3CCZxnB2pCvvqVjkbhyqFMo1SosTdVeP08zEd+
MDElxu0KuKGWDVqzQgKnhkKg1h66YUe4NKRp/6jjzinmOtg8jS3GcVAhS/nTGy4y
H+0dTZryXgUPlmkktDyxxsS7ulScTB4yBZ31An866vjEN3cqPDEcJNQOLR6lIB6n
lSYEyrkZUiEVhPwEod/JAeXiG3Evlr9ju2qorPyLF4/639Vy8kuikcCeFLsIdWRc
/uE7XxFHo/uOw/X8MQM83z2ofK6++ysrsAyGsRikUICFVDW0bwBaVGI4qW5cDJz5
hbLkJ+XF/Ub9ACFUwd2iuyygc/KauY+QfvPrDDdvw2ndPIWYT0YTBPbWY5r94uEZ
cLxYzAKaJbnSqsUoQrCUhcqhQ/Xl5557q436fjKnPn78zuAaHEn3xZHxO40XCpqL
FAe1NAcnoEodVd+n2q/wnOQicKxQ83RgBWdGSXDAc55PH/Sqzx4yRmv5MTOVStoJ
n51q0UMpy2l1GOoqWpxzU+Qr7od7oEO7s9vC/ZLMj1DGbBpbrfxB8CKcgcsAFV8x
7QnYH02ncq0BRxN5ZnlnQWbIYcw8M7iTEqbQb3CSRv1XSqkEsBUePiTg5G5mU8cm
sd2SLlbSfCTHDXgX9Conz/p/uDslEWDhYb5dSbVzAWDtmBcwza1i2SNuunGEhM8x
5LmnEvBmSOSQDgy7PB7B+hPcSL/+6zMiRcDcnlh10m0a2Y7DCa02oUS0ono4Dwg4
qAeGm5yyd3iFiEwf5hHGXzXrV9wTnY9Ca5B1k8tOmPfS6aa3tsIOzrDpWxMDDv/9
Q56ChFSC5caT1iw+pD3kLgjpVAoHFQTAu9E9zyCvUnSRgsWY6fbC+Ud6TUd6utbw
3xDJxYzmseJ4cI0i8gTSWlC+JoAa73ebGglJLwqUSdyMOr1meedJWLXeB4HnRrJ+
0wEDp/hAu7RJzW0eC3M6WN+BhY73T5Ivym1Pyr2Mw+oR3tUNixnqSUuLaOh7T4IW
OtxquYsEM3dKTTMial0P8PNcyHHhJUGLiwAlBWMgQuhZ42DMFdZA+yg0KLj7NjOU
OzR6sGAUkzlvj2vw9p4+V9GasOiSLYw88BiL+WLnfHfBIfVkXWfVQXAS41z8o1yz
eI+QPSt7NHHspim00YVagEv/w/qmRnb3ZygXNGX65x3LIkbQBXRP925gs2iUffac
izq23DOpj2zBFNBhDvisdcis+0tKNFk9ZQrO26/k9Eg3+Sk9obmjjy2lhdY5y874
TpEo9zy2QQbFRgNRHs0KU+ptF78Td7kTLx6PVpYjfhdaQ3OZaxTOTZ1srjJ/aKhu
F67SQeaPiOTmNgMiXyGJ10C/Qnu8nZz3AZlpttoiHPGciSZYqcoinZkKMK/IKrC7
2zw4GMzS9eO1I/uroPlBs5pAteUtMknWTost8kzO/rDNdV1kQgT4PR4iQS74pQOV
QZBEPp76RvCNTQ4J11lcCBR9JME7dAq6Mnmqn03QJsP5mRwk3cylYISwGJqXZ603
V+BB2/N2WJjMmXqd1LV5wUE9BXiWziy21kcNdnc7rsgP2DR1JeW2R8uxN0gQVwx0
vmWp/A6OMU4dIjjIreOf7aOtq6vY3XmQjZoKJemsmQvN5i9Iao6z8U5IdduXsUnB
GqS4QgCHKacv0jl2ySpI8UKFwM/O0ALbgVnA2TwfTsuN3D882aksXLTFrWUyMvtH
8NxtX5I5Auchc598qBbchpRvUYfeesA1/+YY9hSqZQ3KlQhaHbN9m+PeBmg9tBRc
E2DmbD28OEuMMzSdMzL/DIimQb/ZvKVCQ8kWFji0SKSbl6TfJLECE1plCGZ3ZaLl
UyUaM/csIZ8jjofnkDJsynBf2XHb9XfLgsc1VRHXQXIdDOVbICpMLszoHahj5JlF
OTmpBGA52JxmB5MHRn1riWxB0RVZGZFFCV/IbDoF/qZSeo1RWPZcoyYeyaW6BVHy
hXANKROPI+VV6eyaOobPiZdB0T4uAnhkg2S6Th7LE5GLIbMiza5S+y/OUq2KGZ5Y
ESqSy94OBu8rdsFqPyW6uWyjTsbiLndllU3vj0xJEWwW4IasQdUP9r03dyhh3OfW
G1K/BkO7vqm3gsm/1OJ20gF5Q3SQ76VKhT7ZOOo8EF8vWQpm8d80D1oQZES9wOOp
qeX1HJzcyVi09bY7siNQ8yGUzIFFiXamAjlgf8nWph0ceK61cuW4iSaMnTfHnMBX
61BQGFKTnNEriLLp/HAW4KBfVfpxz6xunGCxGpnYTniVvRc58mbbU8Oop0g1dCh4
PodkzALOMmkLpvcxlDAOvjzEOvnb7HfnD/qTKmNLJb+7VVfoh2P2p+XGCqK1Vjbg
3NKmhbPLlbwi3lxTITtXauTj4ZsPzZE4tGX+g098zOgXFLiqCKY3pey07AdhYQVF
LKGEjqbB97P1EXuALnRbqTlCaXvssTFWI2v42jdMaePTFMxMREPSsYpijcnUMKG6
YtRTs79tUmULz9VFH2TPJm+0cDxjss894KIas6ocO6JH7MOnjTHREUJUwS5fgmE6
n/ObMnOAO1j7ckl0eqAfNo/83xQTW8IbdWEKVmCzZqWUsl0V0y9DI0TKFN4kxUqo
f96TlIw22ev7ZtO5MRvG7FZOIXyEMsI8OQju85rQdNYNde42tBOBAGK2q3XMAdGW
y6eh39vgmGjdFZQr9STLCcTOZGamnKc6gGHuzF44atqvYyreuUwNsWkvDFeOUII6
aqNMjk2bKcaZAd/l6DEVNA56lA1BrPPIb16cp2+brgc=
--pragma protect end_data_block
--pragma protect digest_block
iKg21QERN57ZgSqXhvcnH488oEQ=
--pragma protect end_digest_block
--pragma protect end_protected
