-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
edkc2sZgCLNPtF/AcJt+zUl8gaduv8JgT9gC7kTRat5liXK2hWVJMfBQnjKuMJ+T
V+v8IT4ZPrgigAjQ0pbAc0DJL9bGm4Xos+drZVm7de5DOGjXha3UdfYHEfm/bJsS
nfOrzrtxg8xyBNBtEwSC4drQM7b/zxGXGG3WeIhRLCo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 15457)

`protect DATA_BLOCK
aSlMa05uJn3nmJJKreS0Ifw2tWBmgtW1Q/qfb6bZ/MjmKPR+wjrk2mgWamfDh6Tc
VFyKXX+C++WkfcIoJkdhO23IERSLY7uhLw8362titxpyVHQxvG32IPLPtrLxXGKm
CdI6cHa9FgvLBcCjd3tz3aTMUBdCLzppIxE74VHrY7pT85i5NauVsTXY9AP/gxsB
RWJ7qivgZAFxMr1aBAvtJLOwjHDGzP3Bb+1T8j85iEav46XH1iP7Y4gBvk92GCUw
auMkEjbGISc2y15pZGA5wuLwOh+RejTXNwzNhroSJmHG8dt9JAu1rAJAZ+sKI8YY
kTXyevOEt6WUx2yjgL5MTfC6I/QqnIIdaZ0YQ+FBfXJGR8HwZ1bPV/vgOyLRTedP
0iuvuzYFDc35mx1qxu30IwiKqT+CBGPLeKssDnRpzojkwGigoYwouGKGdpEQvOV9
FtJSfNxdYlnW9JRBkJ+a9NQEdE/GxuuP+o5YgRZLLiL2pUp4EKDNWxgYB59GWbug
vF5kmPGMKNuIXn+eEj1jMlMJ6IPAp80nEseY3v50m8MN2aA5NzlStH3iUW+5hdah
Cw4M3xSHTPaPkpfPoZiv4xawPT5QiB+4TtzAsLhqXerT+BvItcjKC3hmffmiCkzE
4268Zl/mrID5gC1zrUc6i4oYxwXAQ6rLY5a/d+c/itHypRKEkS7cWQf+ZB89R6cH
6MgxuvvakowadlPRydTodShAhS7N+iRZ5rqP1KUl4OewOsGXZx8TibM8yfiQ0Xc8
1EJW3u6R+Eg+w47pltZ4MixYqZdDogFzCY+TSBbUuJPxYOr/TfcnbY4s/JbtE1MM
sh1kZxCDZoogTlktoqu+7bCmjGOqMQgxSUzCVPh8gvyp/MV/eUSc/kdRLBIO6XWB
JIGhPW0TpBsuHJONYQSwiRnt7fMfqtDS+6kvczvu5/A5wCxDWbHAb7l8lFwo3Pdd
hmGWMiwtuhHbGgzugDeXzsgy+XeNggDBfHdX5F/QzitlB/LJu8lj8fCaTaHa1Oqf
iZ1Qbtqc7Zv6RKkAAsJ4wVgfkoeW5b0InZd1Re3RealTlGb+nRWiGUTNEXVCMyYV
gL0xmFtCe/F5wuV9j9wAvZ/LTedxbKAlirHUSKuVegUnKdUn1scuw2nGSK0xgiA9
3nbWcZ5MSlIWEfttRCizFt4G0CPVuLb+lo1hey7lPvKv3rwZ1VL4bLma2hdZw+QQ
EVv/wElsLNtf7Jn82ZxC5EbyEoogeCfJT0K0A/PN+FOKbVRAQqRGjOqfm3p8o0h2
OWSIWPupKOVWmJMO/jdCp44sAtbu1N74YNUpROZ/0M1kVwTaUJqIXd5Qf0TTto+w
KEehbqBGFv2F8e8/nkBS0URWgpf/VOpZ+zEOX7EwoW9SHYwM+WipTl6yQh+MVpbs
ZeTC/kgnQVgChklK0JF48AqkoBVApgOQQLVghlrkPH+VQL9v6jAaEdO+ewwwttRu
GJNhTXJf+uDCFKPvcpkOdxwBc04HuYhzDftd8kJ+sXjyechBipBTV4IqOoP0VDPP
iywl89+9fA6j4Oxx7JTW1IeD6V1sj4XA3cHvHhM8fxnS2ECC+g9imtoXwEg86IjN
XObQM2HrH4eJMhmwnSIqu2x8p1mlYNzWqQMPSwy+0uX1Oz31fouzhuJS/bVU+EIQ
SECJz6YwTk269wUasri7yHkpNp6GEn98rfgbx9wjZkDaKMlW9rGXw7bKXRDOgBha
OByxjRMBJJlNayWrorYsMAY9sOlljyg+P+UTg/zPZy8XTNAjYkvR63Sxd0075IIx
qR8juSvNadz5hx2rFmEXh2sT8DBkVgIwp8L+eqAeoENHml35EgAqcTuz05978PPx
vPlZdvgFO8XDvF+9aLPUDoUBeVJTA6PZ+APJjTEopjHQkAKO8hWch3hhaDT8+xJf
mTxa7Pk+RB0FjzqYZ1J/EsmiQohBrwKlybV9VnFPoWpcROLDm/Q5mV14QiTS8/DI
0OOmjHD7fNGxVtXJLfeZICsO4e+h31ET4aQobugFR9lZzLNx8OqEkObrPPzDPK3w
BO0uTVbTMXur+68vibUAXNMhN1pyMAAHOeKszTM3pHXazIlHz2foGe7oo4iU1Hy9
15MyXPG+EUWSuvW17cJkneVMdOV6aPfEbkmilV/FwxHvETZSDX9gtGd0Y93J0Fcg
x+jVCX0hcPN+ifRQOwSRK3uzZrukQuUckL+JhnFW9V1Gd1ebsXz2cnrfBZFNKnCD
Yb+cifOWZQXdDVIR0oL+LIFbZsmfotZDkJwYvrp6wJ4mYn5RgFTxIo7JMRwJiBTb
al7vEKl14gvSQr4Q4TzNXPVCuNNv6V8n0lUOANuPr4Rg9NDbS+1WzrDqsG8HTMqS
Cfo37riJYrZ5GAUlZKIHUrXoScVEajbzHLGHBWz93pCdYylkSLdnW/2WyYY2a8f5
wSO0FkhWBICHh6uirJEyXn2eY1cQBRcLh2r1F4mcQN3gR0lvLxd1JvZimwLjI+Oa
jS4dJv6j/rqBvjbXrgkXpMyiCzaTfUu1MtlN8JskfKWGQvRHzQIlTGjX7EuTwuBC
Yu/gBBQ9bjKYjRhTG0ZfqZo4dyKqo5K1Yip69Mlcwzc1idV5TPG9kKcsF3MYHjWc
ZyrmcePFX/IJVUABQfyuL2wj4EH4TllY0r4pRvswoaR2EPziGebYhEjT/rr72971
o1Blx5zmTvWHv2Oe0eQLpPGdUCWcj6lwClE0Qaq7VnN/V8e9MpSMSSgbOXX6CWe+
BLAw+2Iq8S756+32fAKigEvaRpqB7I9HGkvYsfwxFppvjGO/Q7rQ8HUZK48shDPc
vX6/unBtrRrA0KYSXEA+h/x8fyD40qWydyaxT64nToYNgX8f4joOpv5DGElcoEjp
ewjBZVJLRz1SoYAobhoG5QsJ6xBnjzmFWqAyZkGq9nDUZkjGk9RKKipay7ipQDSM
UO7F26v66ZBdGCvEUwDxkPlP2WRzBWNs5ODj3ycJVvDHIr56ldF5+InAo2fGpgvv
pyv3mAcglJF+FGkwxlZaP6x9sNI7WLygix6snaJivEj6rE6X0J/E3BzZ9L8N0urv
fICnevB7fVhG1/GoBFiYLHdknk5wCt0o7FKat2P8sf3IbGGiJnrZqk/bJnmGA6fX
CCrdsL0fgiHPpPkZ+oS7PNv15qxyqNOhRrd5GdpJyEHZHan24ObNWHADnt0HNIJp
kx1fXr17xpsGOlhqcqWMLoepK66ooXrYau6VGwiGLKXb5tdYGvA/MU3nKVbP1zdb
q99Bc1w7y+4NSPxHYxndSaTeVqyQWOCf5l/OHdCNQVAlDOu6MACgbj2EjnCl3j2E
nueIUNc0FAGf0wSnHQwJRREmhyyxY+L11nFVeO+nk2fkwrCK8Bqsw1NLw+MzAqVz
kRfYPLiE5prsXke0u6iBNk3akvFRRc6vFF6FSh31Qww+uUnnkVfoxdJdzsoks01b
nmx2AnISs/NRvSLhekF7G1I39BULjcH4dle4VM+WMD8lhV32HSW8aWrUltkGUzlc
Zr65/Z/li3INXJJDn97dW+x0/mUQ8S4oiLkuQmGjEdleNbb6Dd51HWmSBCiWok4o
RSA64zvfljkiilw8RQ0ErK0KHbLa8FDq2fUAsjXopkfCvfOE3uIRqlzoNWjrMnvo
Oh62dtkwQAocOHuK92YYWT9VW276zES86BhvU7lo8yjVRJGWk5xOcY+DQXYw7v6O
lbNqLFl3MXtwd/DvWIX7H2CHJ7+blbze7PvRHIfRHVuC9PGDaC1vJy3+1VzfFgGw
G0xBgtIhPleIfh/Gk4og3Zk5R2Z7+HW0Nw5IYpl/bGgV0pAHf5P+TdL85rdmLyyj
aX5kkHPNCpsuEuyoVPzTIcwMH8NIyHXA5gkZqpve//f2VXC1fRBKCZaYP0MoHMcl
zvWTPYeeZ2fWXN6MkCoz/1hM0yMHRUXLJ7FYlbkXo1ZAZo6h2MsoPzy4wI+nY1l+
CyLXX8vXc/4CQOONuUjxMzmK5OEhztsnwlTUCT8aVcDiggn/KujVBvwdXOmCDagz
64nwaHcULsteR/l4Ru8jSXGTV4WUH+d9KhAYgchQw4PSgyyLb6JG17WTWy8l6S/A
srBEBcs8OhCgqDnNDUBnih3VXn9I8nvBWrg+z3ULhLzltGSBcXK6aGU/Yxg36TGk
XI2HCF8/+2H5XL9XO4Yuf+KYcJ87z9aKhnlaLJdeiB9M1HZzyCyp5mwepPcxvvX5
B/ZrfZVCmlTl4iCKG3AWdp3XiXuQGUsGLLMycHD4C8diIMN7I0NrqfHVUjnATbF1
7uDqucHA8B/y+QGrnmxdOgYUXtjUsr95PPQh3/ijgd668AQO3YN2xoEjrdRaK4ex
Eum+x9bw5Sp9gmfS8uCRCAIzCm/yxga2f2xmBvcevuL/u+zaztnueeWkYec8jhDN
wdFi+ZL6OltdmnTSdCWPSRa5IQ3wxxfUoleqsSDF/DPG93+WAMYex5ThASs59FC4
qbQAVGkGq6J/5d5agpGQR9nvo61uli1Z/xpDfcn7RulWnxqMXH4/9qD3tzLVHF3r
BQv/TTRdvqBxAF6909s4iB6LfVOA8nHLM3V0PRhJVyKsZTdbz2uZp1m3ziiv2dEs
KFy3/C8Md4NbcxZw9r8JKEjH3v6G4s7Tvgs+dPJ+i7gNaE64JXaqTBqWXQaMuXkj
cC2ISa1WRpV5+ZrIt66j3Fq3u27UyioQRPklbptls2pv3DHllEDOtmDP3HYyIrx8
ihd7/uueZl5UuHqZ+b3nBY5wmvTPDoUsiN66hQoaHhDiv9gHUPnCIcFdjmbcTQzQ
iIN83FCYcMpX9+XLeS0uPgtX5+XrW1xtq8Us5fpUiOdLz9jdSGkLIGlvPzdaw9u8
F8VSt8eybbnYaeNfiBBQzp5SBCgIgqbPC2Zxi1b1g0tzTkvoSmcgbiyeFZvZQCvT
WFyIKFiJoDrTqXjrf80q4VnCtM5rgGAa/15Ihoc/I6k3RHL1veTNhGWDgGzEUTdx
t0pwQqshEoHDutiVmtVF72UYGXT5mrMO1qvMWVVuZs8VaMFDc3Enfl/NoIX4fpFZ
2JnBoRgLXy9mmNL8QzmNlQwmW2lDXqJp3tui5s3u85Qzess2iBstYxFy+3AnOqnq
KkTNnBUuzFuUG0XCus0MbvTdMFcIbqFQvwQ3UUAQspqj9DQPDk7JutzV6/+KhJu7
jHfHdMgjYsMDvsXDWCT0RUZmyXnB1ViR8PMmLyeVIgj9d3ZXMxeoq6cVSE4dFnn+
70vD7I4ktMpDSvAuE4Yl7/iXNvMx5yPCv+puvYD4CZoedahoPg9kB2coStqTO+2f
QXPLov3fxxjmSd7tQicvl+jKqSH3qOsmsciyyhjl6p5t3UIO1bR+8/eORL7bBLsq
67btUolCBXZ86BfOS8/EHL8jFQfqgINceK5Gthrr84dE7lPRKm/VfsBaDG/8+OYq
Kj3o13q/iANWYpHunwu0PBDOxb4RmPtIu2E+9tA7ARju8hk7Y0DXKZqlo3/gJ2A9
7CZiSw9w9hVtMn8N7KBSogFqGtmOUfHEcqobMFvxmRmJespBOjOmZW3qFbWrB9J/
MXUPoYZivGspLIcB9F0S2LaGAFK2GRit64rf+o6QJGzMILL8/dycCqi4SCXMHFhz
6IbjXWdCTxBcSEucACPpz2om+Qs9XwTNjaIKUvwQ2j0QMW7MWfC5ENIy/hYskbpV
pDb5GhadEiLoemlwP60hTRDHycA2+m/V7cXfEATpjmS5s5PF6x7wxXJlyx6Lzaa9
ciL6n6Q0Z3lKONhYKdvrkbZfsgr/TnJJA/5VLLaGQEmaL/AmotW+RzdL+Sm1dxhF
Z7hsk5HPsHkKWsXH14smy0WOE7pw27YLGoIdtyoHqmRlMefqd7zLt+Lyrp62aPWZ
uowJrKLgSPDjjL/cmIbPfOlug1VsA/q0yVStjHHfPFzMVnxRCQSgkhAYt+geePfP
4dxlJk1Wbi1ZMpjPMSFL6jstjCqjAeVOG89ppHOTbZC94b7zmGdf8Zwp7VqbE50X
Wq9gSiA43N0fzlFTB5/Z2Vo4dUuD/bth898UaXaU+7I/lR5zamrg79KVgglfvaSd
wBDnSU4mK/ngAJYfY6LbNU0Oha5/oKqI1c5WaTqn2N308cYRQ09mhx8swCpRCjFH
qCBkfpa47N+Cme9UM1dwYFZF0f0noEGagoxpqHQ5OMJpKrnH02gyK5QIl62IJdpO
CptG7o7vTB7u7nHubsXCZsmtgQJGvMXoqyFP7cOsKxHnchuQyPcuYODil/tsCFWh
seVDruWGwWROwAM2yNle+BuyFmS5N+PsrO8xdjwX1j2/GFRw/nnMAtEBZRnlmbCR
dk1tb98BxkZow5DEkmQnm4CGB8aSocekyE6olVsED4/RsCHenAk/AUHnQ1xJwedc
RAYlI3/FWqW4s/wf6vQhrkPo5ddcLpARa8ozDW4Q5gwG4YAq/NGpHc0dEAIQjOsz
odqhtUbw9IbeiyAqGdA1cEwGpwJxHlUEIQKxHHCcKSaMH2GCJUPT7Jl4p2NH+x2b
+NdUmwB2AkCU7KAjN2keqTn9jfoM0omQY0tviZhQuXh+AAzdyJu7ppGAtX+5NMU+
+URnFI/Zrqdac/H4CxgRh19fWVaf4fo6G1BqO78P1kz9B4ZPmUPwVPG3DzbA99yL
wXQv34Puqj2OfNgHAuMwdU0K2jpl6BDuS7KxAI/4YkYb9cugBuGk8E7M7AK8DzdI
65PRngDb7PKiwYaO+7OuXVDzjgeUSuAWu1OONh7hBRx6p3tD2ALqQ/CeS8TmaAw0
hJKYLniHOD73XNyGTT8XigUvA4AhPrQxXP6aogNWIYbLV7d/GAED0bWTd11CaQ1s
uOlrjka7I4ekngG4ryOLro6F5HqdMj4M984yViHdm/kqMVLoVeG8Rei2JlWawHlo
U7iexBkeBx466VEDawlexjf5wW5rNtS1YNsFigPRbdP/lJlqAD92qT7Kawp1u0JP
Jz0rDvTC9gxSEHj5tQVEjdglwyK/64hdjzN1CeJi7KeuvjXhIWW1dYxwavABGJXB
2Pm4w1M2kc1P4TQV4Krr7KtmunHjtykVp6SK7szQWgvKYtDMOGGsOjaGRtyG+lPd
Xq5m1XA1dRY+x2OESiyKkKYGbWbeFifexvoQJpu6ZmnlwBLZe1qxDsIli9GVOHpv
WmXFTRQhDB4UZwMsU8NnGojgaTmzFpAFPcXBdEhA2xkSq7BDSWpv56+hhbR5rt5f
FzBcoCxOXjon/0+e2Y504co22ztoMAzDf8XEnVjmzVAGuEVdg1URvpf8aTWdbEDY
jb4z1CMWRd1SWcFs2XrcTudTyJ7NB8bNvvApe8RmwtPDfaPvo9lZmAemkbJtZh7G
MqSdCa71zb01fedAPK8ZWdE5Jws15gjap3GfVBo9qeI8Ot+JoxU11EyI3T/6q6s3
fzUq6ZUfg5VHmQ/8yZLQ2VpBAYfnxGzCf8Xw046Nl7XY82y1As1OwjRVerCt8scv
zfL18ckpJISuuhhMJjvAkjAWWWP2vtLxdxBiSdPYbJrxeR0Cjv9GLY1NLIGYJ5BR
KppcgXndf0F4doX1mB2u0Yi7+1o5Q0QCTMYRJ1+7mHv4Rdz9uZpryhxlZqYKbC9u
GuuMq+P0M2VVrsmpGu+K/9L9TA5Taddnl7Ifq8mZFCPDZ540f1lOUatvzi334AoZ
pyKQgVsM6bUxeaZj+3BT7/B6LJkBCkj7VYxwNwJyBjPsMeC/PZQFai8i94peXEsL
sPOBUNltOAKOojEo/aAZAlOMYZ5u8Hoo4GrBnbwu2poXcCMVDSDwoutoi/HShc/b
aapkaA4O1DTQMLi5FiB2No0RyRmEXx/EnQOOCKThethHQP4O6NZebs9ZUFhbW6fi
IX9wRtJaUWFNWjnR9mfkj2PKRnNbOIak/9qzjy1o2pOYkMlHxQnw7htb5GWIkB6h
nVWVjmyObiz3BpTL7SoLrE/0905J79ycFdl5UMhuRcwYbxdW9+z+GPJziaD74jAJ
sW2koxvlkROvh54tDMyJMPljl6y6K3RtscRpvulOhnupX8Oubl/a9fBBllIxD1DI
KP3Hei35X6oKxGnfbJUbGUtBcGpV3io0oaRicvtE51NSEVLMW9NJol5iB2r69uQL
7j5Vy6drUAxuiZNc1A8RD126851oIWvoVW1hxZb8dO8n4tQcalgz549i6gOqjr4t
fDDinyEEh5v2DBX30CgALKXTIN72AmVLLUd3QiZjifqym4eEltp0QnEQQgsMPzly
6SX7VM+V4qkYV5mIe0Fd9kgmxJIbGJahODTAAWqs0GRympt7ggrqRNw9phAm1/pZ
hHhd4Y/RAXOw8jQG0x/iK+i1FFXq43hpKnM93ny6MKfMsrdCAW5LRduCpAQB6IKB
fknjgBZoZOpn6+OAWBnN0r6Xmx+7GZwCHSqoJEPChxGVMjH6+ck8gKfCPk8g6y1z
4RoaTJD6oUveLiIyr42onCleIV+oiMNkG/MmeQr6nO4cvtkAyucP27kmysEgUtnr
cyrFWxteNkqkf8ODXNf11eFAJhd6k3nBSd5pCGpU6exs3pFd17EH6Ev73y12u0U+
LTxm6lHeFHXBCLAzfZAAThaDcIzakexWzZ4jx+zzlrbeT33AlywhyEKe6ndxxcIw
tiEp+jZ4IAlu9CpOS3OkYoPkBt1U2X2TZhBNjOhCcL8cmb+hAG6NuKlTpSNRlsWP
MKekETbCn0FIeq88LDhUn8IHuesJChlnCCFr0ajvKyUVtfViRUrxc3SHlTa0SIee
j6/X++h35GHKzUk9LN95mdPUARg1uxQHb0LXGIo/JowcyrTUcF4kMYDM2vp0Iyv7
rZgtgKZm0rthc1ZSb/BEm/qZXeAcC+gNmhQBTVujXgfgdFyPqgwIQ+mDDdlvpxIc
5hERqDo8aUhdTsNmkAnajfi2qGQ/kz55+0Sny+f2GAkVls6CDjdRvtt6q9iVONF6
k2eeesPtRYV6WqYW16hJJa2PxRd6pguPUy3QlWADaRMBWec9xhRTDZTKWkx2wa8m
H4RehsofTxVRAOfCn+Qf0rBnlqZ2Z54tzYupgcUAMYFa6gZW9FcGO9DcG3qbbgMj
/krteg0QJlA/VnveJVoFgSM76NqyRbApl2wsYFFVJut1KUI5JidvPS9mg57nPCVU
eU8+wN5fKXCq+4NWlM54y2PhwFAU053Hp9gGo+d2/ItL/zn9SpvvfWqRBkkOfn1A
x/zWVuWpCM85eaIdK8JcztTYmw924/J91ke5hdZIsHtuDKgskqNyUxhmaRm3yKy8
YnjwGc4uAeLJVw9byeSN9neb2ZsftJJmhw8Dm9G/gezpwa5UerL3PQIbOo+7Ohy7
1Tm3D4ulDgMc+9Y7YC7vEvmNZFWj/4atEqpUBbIbpUAvOCz4uHo3GaYhXxRCAjvz
9HjcUTHC0z5H5WAyR1NdslPlp6RHnbONsjbxZB6BL1CY6m2PzzfaDrvUbstBMnmb
hJPQvUT3DhXiEfVpyulCm+f5B7A0kg4xzAE8SBZN58lbjLI7D53Gc/SuzSthfDk7
eblb0sLgIDJcYNxJ6b1DtqEgOg4lLQDThWYp4q5poPR7W+p7rgCOZk7xBqLDoTZb
6xZVaHb5zLqhCflHwCUAISV1e+VOKhj8vrz+hLzSX3b/4L6+hon1AbJKIqPDWs+v
eI2HjDIsMGbg3E3QKvpQKA68Swr7SllLS3DaWn2bFOgu+JzuBMcRUjofJgMTdbuB
sI2p4fX6wFAHjNERtMhBOy5rT4Qu0vXCmiljLcAFIDgESNrASufOpLDTt93gDoFf
REvz8I0i030IzIY3LUF/HDCKF2z0TkH40ubjTBLsVoy/vK56rGNnRweXJnQ/XlSd
nyQR62zAbGCjRB4uliEWcXSCs0kARXTYRNvCxcDwN9ZO59PRMqVZGegAe0JrXAN0
a6xMUMNLo1xopts+a0P+GGL9ue+qJgE2G3xDjfzFhY9ENwZahlgKQ2wNKjmuN2dH
sTw9oJ9icKjwJqUi2P1t7QqZwmgTEPI11KxaKxNArNusa8gYydCmhyph8pS/TEVW
MK2OEUgDpZNXB/QypHKTaEY+BcSAuccazcbdj7bWwOZuJ5f8l6RJET5aOHJSojfh
rvnr8WsNEoz16uw0KU8nm4SC6v5edz3lyCv+vrRNVNjW779RexukUbzGalpSy60J
BGZdqSXEjLE0Id2Dl149f5grXWD7Mp8Xq8eZorWERlfeBlEH/xUt2CI5fEmH7WbZ
NwkYScyt1WJpokgJP6zjiNJfH+p6x3VtGShvGGDkE/Io7z13dJaLkl3IWdORpIXq
o8euJw9SXn7E3fwSvl66IGFAaCCL2tVfADYUPh8CPhtUpdoHMRzRoBRKS0tg4TTj
+VEb7Q4kB1Tsh1oyeEU1UycZptCrjRZYLcS5e7+iYv95NLNgxmTK9oS1fyYPS/CM
RRyhYHdmcWf/rUEDoVu4t0qDVLU4QaOaQCSFlpVfoa0nxOYV3v/qXMlEKUF5mIAk
cgpXh+nJZXwRmbpJu2qolf53fO1na04E7pKkQQ7QNpoKXl4WEiaTmHczl+OWC6HI
VGUrSnWR1iFw9fSM2arvfZlAfIarsElM6mGBejo94h9mIsp01EA+qEoFhPJwbeXs
ZO0I3WKWGFZpQTwtBbG6wyc9Es8Hw5SVInA5UNh+r6RrgESbiZxnnvpNZLifeGm1
JKwM7nJc59E7xYK51WeaghU0PeV6kcDDRwinOzFkKu586tAoHKTAIRYd6leLJhhX
ZqWCv2y4HRtSwY7GZUZmIZLBX0q/MS4qg3Q98AzCjEQ3yPTCdp4U1B1q9uryZTvp
MKlc68jJig7rMUH00HrSgzWsfjiLvOtS3FCKOkhfm3eBPYXRVG0CC6gNdCvSIyay
YIWfrbAC8L8+QOypE2OGIwI72TI399bf9jZVE4MCNAHig/kxij+h4gaNxse0OW3d
4Fet0DmxcncqZat46Ws7FqKgl65BgfnRkpdLfJoOx/v/6NMwwIx3YAl676+lxFhp
BW9hcYUOZpbkI4di85v2MTELMFZZqhn2BWb3watFOF/vCyfbRQsr3sdNEy6Fudzl
QWkDQ3RSf9FljfV0TuDTX5XJw6s9JZRh5uc38qZd6wceOTM8z5nqqUlEzRZdQkZO
YQNzf+jYvzTugTmZNghT/TbCyG+RFQko3fKE2iuCwH/rzyZvxk1HYJQdn697d0Zv
05Ssv+/R8YA1iHuWL5C6wwTDbbfwh28hCCYCB//7Ucx3MLi3eQvqd+Ax0tvlzqaY
hMdr8sMy2YwKsS8I7APhIWtX2rUs3X1nkOJ2oX6/LAguzyQEmqtLHHVW6EKQ2Ipr
A3g1L8ruIvDY/uEBu5x07tprCzGuoQwsnhtJQbExt5YEzmyzGp1bzwtHU6ushNtt
u4JDEL//0cB6A+JDaV9K+hBLgx12CpGoB+Pa6vNmaX07+RhlVotGDy/gOFDklZts
1JhNJFrHE6V0w89FDEyiR2XghcGOrZAauKT0mIe/jROg9eUVh/yZiZ3RkSk2iIhv
L3KIaG29TcITzvC22aqP44PBZ0A3ewwDzd0vSmPkHWg9YeZUHIBpc9WcId3h4suP
bVrIglAaytGU87MceN8oC4+rN89ZKCXDHnm1ic7PwI/BrhgD3q5mjbkrUkE36VRb
1J6gAlHNS8LYbga/LJLy+5hhdAOn+AZpDJ7B0LpBKxn84sf15EKlfBOuVvpgAFwt
W5pAx0rLjvGSKie2qTuQ+8wVN5eoEje+kywRdNfB4dCsPTkV1yNBSOChd39xWyy/
gYhjoDBh53cdluNDWSd1n8XZLZCDHvEucxYq2cQPQTQIkviJbymk9QZJ6UERJbsp
73FFpSpdsctEXCpaRs1qVow/QDsAZUX3/tooLpjxIArFYl3Q5hZ5Dgfb007GHpdh
FQbjiNYR3bfcrS2soms5qty1kO4N2wy7MrTRJlOaCuCdDqi1o1F7SG3vow2kTP7u
ihTVukFLuV5EYJV4vVr2Xil2Jzk+0F+YfjLAuMN54zV5OcQEkkn88AkqMHT1OsMG
sf11vLy7TR5+31e0cKk3JESdiWuDDl7XmALgPiRMVFSivlW387+zlicUeQOOvfcM
JvXW5B2/bSdyxHdC1vThuVN4WbfcIDKtpcPF1qzC3lepaW1xStvfErwRG3ypWa36
hr/hCMrfIH+1hvruvaZ3hSGqQhY6tFn8zHMSRz2521bBHVLeFsffAg4Fc2SlRl1T
6eLWXmwHZ2stoEZkplErlordgWmFKSNQr5q8qIqIM7oKjffXV2763raSlagD7r9X
vwhE0arLPvswragIyvFWd5jT+fwDDWXkqHXtfRKf+qDyaVgCXS/DQYUE+vq6ofHv
hUGV9SRiG7vwv/B9oYVAE0MFlMN9TVoSWbBLA9eX6MnnLC4DTPkFgMhNR0/V6VM+
TG5baW5cqWmUojtJBRbpQ2Ejq45jGpEeNf2AgIG8tWWnEuqU4WPYl4PmUnb9Q7U7
oWNygIxXm4bQHKdPVgP4yyNTIIIF7N1cQq/d06wESZsI9zoAoA0BBWIVlk8b38cq
rP0LrWKz3qlWKditfwPPxL0/QVreONQuOHL/TMlpSDzwoJhPxe/HlIArL5NLFleu
Qo6KM5dh+VA/nBHlcZp0i8FWlfqLOB1CqHnE74vf3Qp2qtYc4zNi8kxBvPS6ds4Y
UaY+EOfF/IJDBtrEoypkHw9fQu+9ApQ29fz2TfXBkiWyHtNzTYxnJGUJoHLBlxwp
fHXqipdW4KRKV9k2Hg1IQdG88ICtRphsKsdAO+WrUjV1pBMC776eHOH15Fgh90vI
fC5MXpMHDJHM06oNNcgFqogcD/soBBhVnAkQBPG8Ki26ZmaNtemjoDgxHn3WkFg8
jcIIXice8PwfpHAtZySkDCQ3W+LkCpcUWki2EkvcUAIYEov0ELtFyXGl4nHGR50a
3HNjJ1hKflVrKa6F/dzqJS19mH1WgcEgyBmJMahTMEGra98e2yP6Ph7ClRNixZ6b
mq88KPghDrRQ+UkUooS79Eoi/k5H+UIrnAbNdBuSJJCVwggus98pz/DeTQ6TWM5b
mi9a/erYD3lkbd8/5cq7tR05/c1CpX8tXQ+0uG8pYwliCant/TdQbph/kKXIGO/L
zB9SUdPz8MZes8AnLuXM8BNEOFV3Sfp+Rw9NylM5dGBGcjJcMEsxkDksPC9OGj4S
IqvDFwwsmr6eNfZeGNg1RbQQofVxxqMOIDPJsk6M31jiXzBbWLrTCOdguCN0i6bC
uY/Tse2PQMJ1aWLwrv9Lrz8dvLXYJ+SYwB3ByHUHInql42Ug6Xr7uPv8eLuMTNc3
ohqtC6ShnLsUkaeJGws9q+GAc1Bfvn7DZr0DnxMAWaild3KHGuml8u0Md88DCNhm
CY/6iSCnCAfpytSrp3l6yyJ87qvEWShhKhN+2/qeOAbHmmvYqLLvhqGV0S+fqkXu
Eb29tlQtaDKnnQeOWR4Ac6hQcj8dWV6mRsfU0vxcJrFiQSC5mFntFsr7CpKE4+8T
UUtUGgLLZ4K3A9fzlAioxT8oewWv+yVvVxGAx+jyJb4avSYwWtRjHWAQbN72j1pp
Y/t0thQ8wFQFSDKYPSX+5+kXPbUR2rRqmUmilqljPbPAGhWR9eL8SCvF1hE/hAOM
3bX55U3MeAeKIAGx/f99cmjH/UBE406LrYZww7tsY6QrywIfk0dZUo13FzrR9gmb
SRAHwKaFcTCSVbIyTG4orcc4JrppTbimutWEbs1YYhHrsSuUZY/T/zBTC1jvWkjb
N3+fpwC2q1RvTRf3H5AKNIKI36P138abmtht+2VA6gzj+0fcfroWGCVJKJjbXET5
lBJBjcfCTqjLdzNgJNVyKSZh+ZoP0YXT+xtGclqI5ntXMu3xOlqrwppPlSDKe1sX
8bYg/1Bs0aYycntFMsD1w8hL5NJEgEoawaRpHRw+hp3VATpHZCxHR0zahkDKbi9v
W99Ktd43nNnC8JesRVGiglMjmbczoImIVXFPMGDSvX6cGieqcvy5PMmoQmOJ4VUt
CFwE3eQ5RysoW+gJNxkFbRb44bUBhtaFBitavH0H7PsDN7945KBww/V3icRR9QAn
aKhIRM+CAKbvNj4tiiJm/ydicc5slSu1wzFumC1HWDh4USD4DXlqfn+w+nSfnQen
wiAP5SfilZtC2HxsTHVCvuxh8rbus/kGYwu+XTsRwO+iK3XWsFDH5KVcJSIp31FA
qXkzor/MoKOL1Zd1XSUAArxllApHder0eqUIOclU0No2hT1wi2yLHVUORG+usA8W
gE5yM+hTxhBJCuT+PXqf1Fykz9J4oWY4K/Z3FRX1gFUVPXZfEL2x1HSoqJ/MQn4i
8PhdFCPRp9/MugSgnyuBiFooozgSOklmqrYoBjt9WQleB1NXuxZjaxNNVr9qZPuw
zg+yc7NHdgu7Kv6nHhyglkYQSB/tuk6PjX0lExJCjXVfH6GsBGoTLcqA4vSay0Gy
rBCAh33wSMLg7mOhsAjHis11imSjiZOdWkuIqSWfUYICeq0T/vPnTz29df+/ww9d
b7NpKh3NSP86+csnzNkZvCVVjb1Uc/0wvl6Qih4sTDg4U7jCHdMGleQaRQls2Fkv
RKjS1YSATPiqTLQfaeRIG1C8Se67/ME3I8Ov2cRXJN7K7mGjt4DDYLexSYEiZ7kL
a7zFx39RjlGn4MmcEuEpdmzCOdnY2peaoGm7AhhwIPSFTkpg26Zqf0fUWU4Ea5R8
AmuuHD5L/Vv/EgjuA87btvaOzfgpNNYUALiSnELh3UeHsfdpvTUlPhD3OMtJUTHG
fVUjtHAIYfqYFJ81PC5LOBQYFtJ/ofoHSJUd8uEkZQoanxIWIe9b1N/D8ImGO3N4
EaAOF46vG9vAImIOxEglKsKtLSbcJftz++luPY8QcZ5EEvlpFzrfgam2ohCxUx1v
22kKg1Pni5QP+5UxqP6XcfmYsD7sRPBE+QUDA0ZM2QFFtU1LjuqkH+gjeSmyZhoo
Yh7l5DFhHCAYjh0JsiIXXTZLyiPLehEB9DwSLwDbRWA25wdQkARqozctNyIX0EFB
mOEL7IAw24XIF+s5yArngq48KOEHZvb9AnitYbGuj3Ry56PvuU83cal/yLYOrkEL
Nl/aIiV/HjDayGyUpQwTQyvyc3IcGs1OzYm3fzleFuNyc1wI0joQ6SqNKy0M6fU0
IIfIxwOepvgoHkKnL2OIo//REVMdr/ef/d8fTyq2qLsIxUFR3OU/pvLZHq3czDUU
0t062R7Y/voJYCms6WC/JZqeweh8K32UU0makL7QyWJG+eyW8QHB8X+GfQ/i3hvT
pTvTNF4sqcfjuEXw1HT3IulAGTtK8gfuY2reMCqhk2JLq8PfJAwvKbdW5digAXwE
dc5aCSw3D5yqdNPayAXQ+PGE4kTxCUWeScNHdbOiiDTUXn86Ioj1AzWDoiWPjNNJ
EzHWeLMnlr0b1hsletZXP553oVj7/F4mDq8dGnuAGnN92MKVH7vHfGw3aDGMeqmf
jjub6gnpr0vjgY/0mArSppvNoKR8P9QXiChVYZUV7ae1KEfWWvbkk6T+jlWNfnH0
gLlhtfMBfb66JN98D64AKF8LsWezdF2WDyDDpJ/4x8JMIOxgJ57PON8u/tF4yOKs
wqAw61sYwq/mvPt/udXAwsnwmqbp0/8phRHUBmp9QiBqSVASVidTXwPsEnLu+nHq
JIm7dH20lzR32mkIAqHMCpZi5R2Gz4fRMzjB3oHME0luvxHfZOxrF1bpe+mfRAof
X4b0HE8Z7vgJNLB17VPxbncS+8R4YehLeefSvewxSJ/xnGQMBIP9JUG0QmuWKTvd
whRO/tatYocm9BxMRxcH7/RnOHqQkjJY6FhKu6XV9xWvj8WGjpZuM2QjU5uFWGh6
a+CG9/trt5itHeturq8eeiVq4qeWr5HP5ccSXpq5DrloDfYCaXxvk57pGIQtzm/w
qEVQy0GpefTPHkod/gP2K/eD1Le99ROw9KjQLMWTU8U1euvB9go3D0rfle8J3vCq
rV3Hkq4dUPb34eQOhC+HgTQ1yrQuCE7MJgpsQK0iLms02ojfcm4UU0PnqwIw2VBz
u22qbcy4limPyjspgtYwLdnzB7I7vDTCJYSu2je3XmSCnfJoVB1GQ+CVhyozcXdn
VhlWxhGk5/xRE8Eu+rtSOfSPaah9l5Kn3LfhPHGPin/+7lBNznq+jz2OnUPCifim
ftyr5ZwHjQl7iY/CThj1PNUh6E9M61a2myjCOyVddH57LXQP8qbo1KDae1IvZaPZ
7BiUfv4vvhrIwMJXAUpvjZ/6KzLr7+4oCLkFnalUIkKDdUgxEDtG/PzQLFpdalhg
fauG2iN/AKcLW/ME4JZOJbVlPzW/eRCnzjBIHkTU4EZD6JodZPEJi/6T82nbmOEh
jRcW9eFXaQClvFOr8FIDQwy/aV65IahSqdDT0MyMED8BrEg3iZLazu4w/Z7Q4fQe
07O2OslAVtKdXxBSCHn4PtKyt0obJYqDo6P19L+wbm5/xKAMaIoGQgVcXrRe64LO
fCbHAqlk1XZo/33LWKegeWTDh2wUsfDuP9hi83Zrybmvj1z7Yqx5bJC/NiWj/+b9
qB5JkV9JjKQ6pL1e5QSWX7YUAzP6e0QaaBOm1vLsDOMDtl9jEOY9zQbIivypYkMg
/nI3xMwN8+A+ZY/+e4ZNmKZWqyW87IEs1eJwpMpjFhGGpoxfsLY/v7KuGJETDBCN
BFjMcOkL/5t6n/f0kXZAlaLh30rvaOepf16W72NOHapOXUK5Qz+YYQ60Ww8qC767
oc7HNTu7IuspgX1ZIe93yA1iVMA9z/vuvxmELgqLCQjyEsU9bpbhV6PA3/iyU2PK
KawKe1CnOFqeWdgBI8A5OavL9uFhB3PkNcZlRGLoWalv9jPdfxnS8Ij2bsMfxnyJ
013eHd9OUO7tShy1rEI9ScZeXEV23rBJS7Wki2Ner5Q3DcqhXbEQu1ZfoVJO3EJ/
Zd3N0cT5XoPHxBNlBZzzZX/D43rm1/EESdfF/nYpKcSr0wco5j789W2lHzuL0TjN
SmUVcwTSMq1em1SBo1hFi3dJK9vfv6vpu5jic0QMDskSN7gUdbiiYZhS7bUf8i7J
cXusPc82VjSErmUDWBtdXzWYDkq6l0TYLAAU3yb7E8GElJrFnhOYgldw4DMLbMuP
+O2eMgvbcUze0xCUEhzRdubqwLkhxGlm3rg0lEHDCDaD/8QpD2HmrPYIXBeOQUWQ
NcF2qZkPnkRqIVY4Mt4TtRnyEZzTNSNPhI4tZcU9sIG4tR0xcE8mL1UmffsKtVlq
RM8G4y0UEcqnO3UmB0OgHvajNO7DNXB7FCWB4sb3HWxNSH7TMDb9JmgePIRu94+6
5Lxb1NNgAHu7tAosAo1ot19uQLijhux17rFE8CdG/DdoRbsj3xAnUd2eofDbEOx2
a8AuCUTQ5Ft4205grZKHaJ8Rtdl9mYB211hjljGL+3BRj0LMbrCft8BgVX+dX/Xd
wW8qE3satjzxoPxjUW9wLQ4KhQ3XzdBZFJ8FIYDRAHq8z4TB9P2sVDCJYpzMiO/Y
jWdp58Djs5XyQRfA4T1v7Ljof2ADRyY0zwrG+ey3E/LdhyXeYmnt0z3P5OerM8Wi
45rEgRmsQjDPZYDzGS+Fmb7SCacWFZTrLUrRiop4WCVNPz5g5WrCICRYxjBWZ3Z+
pFjKPqTaes06J7XbSscQ69zoSpGGGeK4q23SPZbp77d6Dk4vXqYKwNBaOKgJ1SHJ
D2O9N9afxvQ7PqT9SQ/fmqKzyTxx1aH1ahWS4fo3VASSfDLZn5o9YsQAI87mLu3l
OhdN80jAZ4hpUinnE2zNVBuKS9uwBlBvYgKN5d7FysGRgVuQGF7NimVSrr70rZ42
VYxt5z1jNfuTjOkqNaYYayjnc7MCL1YsIFHkjxPVpYOODrm47dtGRhGwrTLLnVBn
z5JBWb2rGeW0DCRTyRQJd+cNWVcacUqSihoNHkqvDr+db4ODmjHVhnaPUy7H5mrU
owXoONnxeuvDxgJVflwsvVOcSlj5YeblGwvAAFLyEyz/JdlxBahbJQ25nbMJsBUA
2mWRLsGAmC3s2VcVzvdGUHpqeSJR3aNy8jmFl92KBVKi8L0n3+zeyvhq7HMerH2V
sJW/LK9cEujWIPoKbs+opfr+LDxmgcgLJoRSFq/NNkEzl+0Dfb7f6zBxB04roLGm
cIsD4J5qKLdjhCCpxlDqutEGvlkbn8VQ1WfhIjDD74zpQetw1t+d/8sRvGEq5c0u
IgKhEZmf1b8WHn9HBshBUmz+BfhAqrDY1UHrVbfF6ky8TzR7VuvcJjNnzLfZ0o6/
YQ3VHcVCqVKaYhpAY7v2Su0/SAnHzUKxdBBQ0VixhgIkqQnVmlGASv/B0cwClDEe
Xx1gS7rzkkq1efdcVqcznm+4ODEOdH3aFdYEiZOhqdy2ARX+hZO5OgWMqLoTaqwD
JlBrsS1HtBjSgKvDyVs1nKTHQsam7PRFvIS6VqV2x4HuX+LcgdOe/dy8KLiU4Iy7
0RpICafC4qrnp9IIogFDSpGpxX/ysWGCzdxIqa+ypW+tERMQxNdoLLkdbLRvElJS
Rb5LCWWXzOe5RInTS7NCI27EFvI2lUyS5fFC2HJH6QAEy+LKsCX7ByisarhNj5uQ
oFGyJLvA4Wb6HTsFYIV92n4euZbO6P7/b8FhaxyL4rMXaGeNkmJ6TxjPbJ69NX3m
iRECyHarZ4J6gVdjgwJmWuLyoqL1WAeNf+h4eyVUWb9aIfB78ZXYNiE/E3W7s+vN
rKWNLu2uzCPje7AfjR8IYhTFRFN0ogrGB6oQAW7gGd4OTdece5SCnMsn2lroiiew
/6hLSepMUA65pLI9fQ7cbn07MpL8erWAlnrL45QDGS4K/vaLueyELfvAIsfaYrID
1QbMonT59J4PCi4jKZKrLgKI6fMJymcXmO0oesMBXdN0Ozh8j44N4BjLrH6IpQKk
0ptBk1YXD3LfWjqDKXe4GNzGdxfqkWX41NDPoBnQmhdERxyvlVpO20faUKKCvO9P
kaSxf3sUPR/xJTmkmWatRF+9s7AbVo3XbDnC71NLV7tP91SPti1Va7ini7j+RRMz
aeY6WdYRR9k0Sjxb6OtRu2gO0gssUJw3LvLwGS4skPh3uBTR/un8jMjyc5H2ETn7
UXvtfotJNN9BgMH37AQ1inBVvN73Cd/pLFktq0eVwqUd+NbVnlaOSYm9w8ExM7ru
MFw4j9sF9tmHHvhjR5Z2q43XIoXinAVzUYV5nZxd8YKkO0bQBQZ2mOGhV9pyvjW5
jptHLXlygtMgqIqsEQYUqn/rYUqRIkci19b9amOeU04khOkuu3M4OGT6jUOZirrQ
GfJz29fq2LIVyi4nyzcqSwkbdeaW2prJOmHwLgcUOhZEjUoSqFSmCY7vfxH8yCOd
eMWO9DMo4pHK4b3LGbNPBWuxKQaNtqjWzRYf0TwDyiDsoU1Tk8piCJA48i2NBtgU
0v8Ak2kulvtMKqOmzd9Ey6FaType/Wb+e63T1+M7i80VU6f+LaSR6tKJIto7thZO
z+se0bDLaNn8z8sAP2A9Gvl86MSDOTdg2Mk3s1cr5R6icXyx0jNXyYykeJ7exmuy
WeIVnoQnbDwhFXx8kn26YEW1AxeO/AfWBy8Mwk4nksi7wrTzXgQxevgL3eit7oEy
rtO/qQe+lCuFljDm7rQVU3oktmY5emh5iB4U6bbG600EbmP5MWYAlb9c8WTqUK8T
PXY1jomEpm2IGrfuCm9oUlB0H7MmH5CyCr7ocRqPz7eKobsgNmpLkRh3biqzDrXG
4q1DtphOaoTfpkGzEJZOL5Qg0ZophBx+35EVnEoF8tujS3e7+1vI/2jPD6UBe939
EVdLl6zLcfnF6kxOyrl468rniAvqNaOFuJco/AOHF1IIWMxG7J0s99FIycIHIe9l
wpFu7YFZdQpnvc+a6MOE4aOdmPpWeFPX8zW+cwgGshi4RHIjhhn7IH3+rlpXfF1S
Hf2UxXhbJR6f/8pN/DqDW2klLrGD6xruyEffe+JbG7TDcBsccG1LYXQczbahkwAW
wIjVwJZicz9KqkWTUFJ+OrYYGG+iMOnTMRf0rDQqs/EX27QpJwNzMkoO/7NsR5Rg
85ZQWJ6NWq/HFTwuQ00Jx9D6Zp2tyvU/kANog8P2aWZ/wIDM3YL0m/cjGWkIMENG
PAocM1EqZIeG+B+FqRTeptJgakMalNJrSiclrFunl3GwQ3QFD7ZPOormQiRPpC0G
DMQFkuZYuaMf4lEje1tIewRR54KBcU/4xJZEbm0QyQQy4CdY8S8hznoXao4MsWCM
72IXB06tb2V8LP8PGcPt+H8sH2tjiDuGeQj4nZ+nNAWBwMg6TDTLsRmI2PhTgRS7
Mizevg9I3tG8SV0MtEEH7tekGUCYkB1zZKBpRHWHZiHaar7t8PFbKTtOIb9czicS
2FpS63hrKqtnEM3RGT2+otfYyFfrt746NKW7o9DUWapync2j10mWSd6dIxONj5Y5
8cgfvO5fA/jYDka1FbaPW2tWzZmLf+aZ/XTDy6SeNJOsGDItEAMzH9EkQH/wUOX9
i9pv2Jda8NVtFvUs3fl1RUUTQlP9+zPBnGN7hT+nps2vQloNKP/VclTSDYk8Qz4T
jCViq0Vcd4njGoDYWo7CTRkaDisEIwyOnQGQUdGUROg=
`protect END_PROTECTED