-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
dK8KodkaoOOIxXZ8I6uBf8R/tUiWjgSiMUJbdp797CW5gqkeeHPBBUBg+PfR0YyL
MATXbg3IYHBdFmyemeIA/i3Dd1nuGU35g+3sxVYhK0jUKLiXnSwXBJiHPNhyKJ3k
EOJA6X7rgPvhcH/xunobijmjJcz/qJBcLvLWS/t7kvU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 49772)

`protect DATA_BLOCK
5GAAT8ohlccvbcpgki9xP4fBWGTwtnf9yuRyk/058MGncBDNhNMjC5yW4XhHhYUs
Z3RelVJSZvDmD6UwAJXR5kaNJ1ypWPd5B8t5zw4wwmzlMaS6aZgqQSVFsylCc9yG
6sm0Wk4nXgttB5AF99NYYT9xmfMI3pquaWI9T7LOG4fVScQ/Ky6R2QSCLErJmsot
IVSGRQ27uokaY/zPdbExgzw6w19iAZfKE+5OR2A68xUiAvWVbsUQOutbquQ60rxk
jwZwVZyicdQ2OwCAwK2fNDxPU6MPGwbvJJxRPF3V7/BfOZna2HEUTxtlwAdrH8Tt
DlUt7vZbJ9KaCKWacP4WFxNyZFTfItppg9y9h2XWfE1ub1OBx1ZY+PdmpALb935K
PLtjNfI+6O/GEetruqCzqCMWjOGr6Vj2jrVuoev321adN8wzUZKWFxc3zap1EYs7
Vj0T2LHVipt8E5Bcbzujdabb4J5E+J215KkdbowXkITy0mzmG1CkJO/zP8O64CTG
ze3U+TUs6jadhsnU1sYtNakde9fJqbjdH3kJCS1pW/tCUS8foc7flT1wt97OAPjT
rBxSNv2FZK41PR5tLsdbiCxOLC7n2u92lyh7jIrXoMYwvsw+gioVgvNOJjMllfZa
FCkefwMiUSYCIbj/A8Zj5eAwdJ7lOZqA6GCGFeSFrMcCd7sDZgq8+yzmkfwtqnyI
TxyGEgfiEhizGHS4k+zSPT1Wqm6SUr9koXWyO/t8mc1MemDLg5bnPp6b3SnjJ0Xv
MuSI+tZmyZDzKu+bVqFIAkFCPXhfqWMOcddANzS+Lk72Rsh6IGG5vTXa7s4OYxBh
jOS8za330BRDhKk72p318X3AA7aV0+j5R8uNclhIm7v6J7kuAvQ9tWmFa0vbFCgz
rHsThlrp91dMy5S+zSMRMkWXefICl362hjwsXsA+CfYbgOUdxfJ1uE4DFipe9SlO
8AvkhIqrGvbQqz3EPmPCo2LYiC45BikvEqjt0RcKav3YbUeQbsWq2h2dmyPr68Z4
OBMtbEkuga4zR/jgus58FnbYMpc5jHovXuufNtf/F6DHsfpKeKvuMb9TToesb2J3
pY4smqpaqG6k7jUNp1RejG+bPiY/H3CY9pHYEmHp953Vbgq2Y/9qLw8M83f7Rr/D
tl9KXBhPWD5ETwhZTT3DzDHsiBsQnzybXkHJ7cCoHJ38rRuHpgSEK9llDBkLO+v1
vmsJnqST85YVR0zuu+X3rtwv2VIl9Tl+SRtqPgYhrZ9zkxiIaRkKtNJf5irzjiJk
piOrQxisQldMENPAgUAIA7XggVPdZ3iSzGv+RLOJVeC6o+Z6PUVblVRYKjIU8axb
x+q6HtPYkK+p25RjBKHEEwKDMzgYiZV0o31zMNUyylrNSLNQJMARKSgjgKOJ3HWp
RxzusNpsT4nbYB5/uiO/4xAbGPCoqwRUji0hD+m2MZE5WjPCHhIS/Nizz9/wuWfG
ejQTEaFzphB7tL0q7i+5pmVE4LIYyLsN4LhgpCS4xp2z0xaVOfATVM/LMT5lYXL2
M+yAYWwfGcKPAxzCmFVuPUv8WnOK8oC0gl2NcquHCDWR5dcZWojr1jq9CaKtUN4e
jbBnj5YAru9ScuA8zdSCiqGfQiCG0c2Tr4nSTbHJGqcRqXFODveeZj+dD6eFj5jt
HpAThNAKmvdAgznOjQ7ovbmQhsKil/Mno+YbO8WzjXMzaKqTyOEo3Wbk7KqmK+Vx
F5Qn6TAY++X+IYS7tAYGaN5wNVTVKQm8lI/phFmvfQ4FdIDlyMRl+D6U1KNQQgOb
Tqp+tkfMxHlu0MP3bh2+6exifj9XrMqepHYThkEBcMyigRVEJyk/OD5GWpCs7nMo
eqQ3sQnXz5Kb9hAO6KsuVFF6ox57cwpgJf0kKLCZU3vRu9CC+zVzvkq3ivAuP+mW
Av1JAOKrAADWazA9s/IK1cR3+MEV0DYPXc5z3KjLzdZuxzStvPDnp+L3XldGhTXP
B6ImpMvHMwnFfFjNBtzYWDCB9W3zj1RctYWs4Fitr7/OiMcpoBijV24x6DyD/2q5
pGBbxAfAtxO1YGx9DxalmUIGiCwezYbwhb2OuTiit25HKrwey3HBEq8B+w8FN910
mg9w1a+2X5nSZs/PWseoPyGTC7K4wcz8uwaaF1NZNj+xdQaFN5q6U9fKFjPX+cMr
/s9V7flGl9S9EMMswFIeEW9WMe0RK3O/4KUADY14JOIML+POXgbwEktq7G+VM2Xf
hmNp0v4g412evSnS+ozcyBrPMPfGY4zfzGpZaEJsBiuuTirW2mABh/js80MOqPgn
LoOXml+tG1w6Nbu4uB/CtGuatDjubCsZA7NIEdH0olHXU0mNR2uhgs7HBiSCb/x0
M6jYvRIO6znzC4R5KXUVRIZdVyD+J8COi32RCvqfaP4AjrUGGb2eLzcFGZyxZFKU
QzXggfyvn03DRAzacg5VjE1FeMFDdnza+x7jhdBQM1sfsCSHI8KrurDctBgViwFn
QQoMIDeCinQ4BPC87Ko/oxLd/42yOAL2w5GcO5LInbjDxWzQ+iMIZpYyrn22e9Ym
xRtiqLCOqTZiGo2Ni9CaW+GZI/XkAK0lHAewWroIiJEE5TCBk9PpAjuAVyZjuqxZ
5z/aAVQsWbxspai3z5bBrcyz0zYIczCP6Xm/ou6fbxIbtnys8tQw32/W2I4zQ/Ks
2HAj+4Ps5YCo+wZRc248DPmtIKWyWLbpMJDEeqwkT//WdjslfJ+h9rcauy7lHmuN
3x5SNphltq1AJTW4yWT6DScsdleZluN1XqE5fptU7F+eyNClBijaFVV6i4GgbcIb
HclTXld2zHfN8V5uYQcqQjqwijIDQrFtw2INBXE//bOdpi57pbrVAK2SXKpBdz+0
nMWcWagH88ccKbRqqR/TWuq/AtYwT23MSYqDfxumGZlhTw/Dkqkd0SaBAnCHkEc0
uPt7uvZhrjdfbZF39Jr+dKh76ZgRzw1MTGXqBGLGpLAgYa5hejWtLMclU6TsKcq9
cpp2kH7yoJ1nY2xpWkMVEGrUBLyNgIQc3sVuSZAVyfRgr6su1fDpmOKnV+Ap1rg2
dH6rWeXPwJtV9MIlp9do/cDUr5HLo3CHju04iIWyNezCP3gU8t8MDDCfMY6POY9N
p7DIxZFotYJ8YuFrBS4AEv3Q3rVkou4q8Rh7Gd9hgwKcnFkpyz5MQJ2t63JDAaNa
bxQd5bGk4Eceh9JhGPg19qZRGur9HBF+FDAI0Habw7oey/TmirB1qpnJG4FmSRoQ
0Qa2Y/DB6/nVtQb9onYaXejWKVIz+J7QpPvuY11pb7HTP6mf7braOVeDB47eDO4d
xRrABo/UU/+jNhNCPpy2fd/Xylih6sf5U05UjG+HCykGu0EK7WBLNMU3jXx+GlFv
woln3cENB6za1Aa01A+Q1VyEsml2/Htnv11gxHkNaaoltkmpuzPtP/1Qlxlely+0
AgkdwjE7o/uRV4WvpYmpPpP+5W6KaN1rhioTXYwZzk7Bw81Ml/ljXsva/4g8V9Sa
PD/56e2ARnRAU5kOifcsv2M/TlNbd6OGrWgS18/Ft3L+cFkgyYvKapM5iST6HA3H
6mm0dM/xQ74L2px4MpHAqCd8plAShwsznVHWATRg3QDguW60G4+O0KIv2mA6rAXr
baMrMM7wem9uT2PWOukbRecMs3xN82xWCArQAGqu7tiG/VRiMEnK1NVLwBURrwZU
uCqDuQ0EdEuVm3XExCFUkJ+96CzZsC3Zq3eFY9kNkxyJnZ+qPVx4WVxh/wr+l3cW
F/uKGMC/7wmQCNYj9+uzq8xKNzR7NWT7rfs4zDTyj1l5YIwbXgiObaGd5qII/Bp9
K8r8q9HBUmMG9rFHNVdBd3GDAdbhAnBtXtSUEN9pctgakiCfKOsEzmm2sS5pDcM4
i8lOyIujNVzat9SAd89rDEFANSA6mVMclMCwGqra1ng16+wm9sy5jki8Muj2H4w/
WVM/TplNOz52PKpYj8dI/886DnAOgTCw8O0xshsMNDeA/k6XCoWbKA/pNhEAtz4m
bbWgj7VxcQeMNajJQLV6p0OS8VwlMV5IbCdMGpSk62bCjBES774cVamPxEw9+Z4u
NkeZfLg1isei0BK2fvh0MnVQmql7U1zXhF6tS1L7BRtBtuCG13YXQAtHARVzDjmD
XF27VCgv/Sn/+1brV0YvgTfitNagkq+7y12lMEtv9EX0BJBq/XUN9NElTQUTeWhZ
CZdf4VOw6Hd4DAmku//bC9jB+jR/6kuxdcK9XrLNCsVGS7zTouSy3qdyyyjcRXgH
JimzYIEjQJTYM7H3tAFqfLxo5yOA9TVWqMSoZU9Ipk4lF42YE6jNo5B5+9kS0BqE
94s8U8mVUBorQcTnZEPlG2Ll55Re6Je6i8u2BXYoqqTOLvRNfBJ3bDMS85nrpd0s
Gz7oQrrE9kA6deC/uoEpr7b4S70cj9X97h/GvXxYx5ou9CIUhTMcC06kMcTS+y/G
GIMhQBZmSqbY0Vp2pcfcUycq5OFT0fq5K1YqT0vOzSE5Wsjso+h1QyOCl9hve5V9
v8QGIEpqO5SP+kF9lTCowCA9aoNfxCpAbEfxfLrkjge0oM1DvXknOLhEIX0lwVCu
yC3qh1juxyfZMzqvk3HLifXHFmPuyAmQbqkmK4CyFA7Z+fK/l3+xoEDCLSrvApv9
1+hdDYtTYmruZWRKoDGRCmkj9CkrxjTUDgh77MWXFvx3WuEB6JcSBtBve42BpQmd
3fuoNFQEW2nDep2tLwmeAzRixmMiX+kn3wL9HWGVlm3c4u3W6iot+Cwpf1azu9zT
HG0KyLxSjgN9AD7OqxRLU7F4KAIf+iE8WQBc3soOf6aZYgWqlNFaXVKSTwximlsU
A08DJ8owY/kdHPtZQkx0Lg+QG4omUhH/ttlsMPXnVTXdjrf1WP4+fmDWBnF+mm16
pBNbDQyxfqqKQRArJld3cjxmMJYxQHnVtPzku5lppLzf02rHLrbwjO7mGeyiMv/F
SBorURTYlZY1SpQhQHu/Eh4dHeW2kzvej0ZLm3dbtY/D6xaRKJc28oHFR7shwiNA
hGiyoab/4BZD2Jke+tWt1xrPYx4ZO3Q+xkNJHYsjy93PbbMAJ91cb0XxYrRgWV1J
JlSwytIXWn4uCON3dn5PwdzTrbwroO2q5vq+Wk9aLf/TdxnrYGbvf/LZmyiQg1gi
iufxm0Tqe1Rs27SUFZ/GGsK4VYQVJ7zjj6QHtCgLXz9pe9x+u5Hr9Q2xVm9khL2X
bxV0SV/XAAEh4uQBLj19bi/kh5unudIGwhcsuVYDTuebsLlfl21eonYLUM1P90UK
lr5/kr8jHjoB8FREzidShekum0kvm5V9UsuIvrTo+9yaXlNN5vOtEX9RaVMzOZei
YLaZ3/DiQKGDLNwVxe6XBzrS9/4SyQ3KLC3oFOBzlBEKNBeaMnBMHVN5xDehmAmW
YOGNeq8HQWtyZxyDJKbRVXYejdMDKGIQqQ4WlV1H6dnBJP5UKnE2/p4IEHzDRFGC
DnhW3hcCQuT114wFTu1ilwVL5qCXAm5/jpm9Nq2GJTtKxi5dDy+C4eZvY3+3LH/o
9nE/4iIqD2HHo8O2BXidzUCTe5wB4QoY7US1q3nFmHw5MY5lpGXC3MciYTsIKHCq
bVliuCrXiJbkyuiL3BSTallgQ3Slm+bnmV5+Ib7S41fMNYe1gM1TOTU8PCwTANNf
8zek6X7iz/HXQH+d2kl6wPvFmFdp7CpLg5lGvZ2neGPr9wacmMwC0kRpnk1uHLwh
tceFnIMsxOZg8uUzzHRLNsajCKcl2651pXL1cJznsBtjmkmwEclK3uqPLrwR6t/A
T0WtZgr7C3hB13xEzOfjm5PmBELkDT5SHFaL3BlMod4lQpYEzsM3U0GF9s8n99by
S1DTMfvtFK2NDbJUqMNW+XogttePEHZOM1Lh45GlHloktFvDtJ/CzZcJUrjghKR/
qH6JH3Cm3+81elKvbVSisZn9Yiyjx+6bCeVq/cCqKpJprhwG8y42sVzb0N9kbFwI
BPEHkUFS5ftPPNPVVpEImxxwCzLvYK1TsbQmb7MDpKhudKZZzvVQDsY6IyG1+bC8
cvmZvxkVti/xpg3zmZeErkl/0a2jv6zw9LpYxd/4qiV3J6uWDkm5wjnz8wGJp8M1
s9gW0kt2ruxshjUJbXQ3d5Kfp1NW9VebXoqtYDh0YA3oCa3bsf/oMoJ7qMv2Y4wc
+cXYPqlEteyMPnEHAT2LMhOS4jJSTWa41tvsleIT81DMLO4yRK0+Te/1y3VyfNbL
AdU2Hn9LrILZVqy50ZTpiVqcAzXBU+K4NpLLeOlS9B5WxaFxo6fteL1qFe62rtrj
j5aDfyr4A5mVeMG0WpSHG0BKepMOCSrg1tMocncucgZV2pTYN8AQDJXQnd3QlhWU
avP0jaXb/jJIoMoermhKJEAJQq6e2XBDNFvzBaky7y7LfjzCBVG/gwGSrFae/3Ta
ZTckfy+J0nQnhjZrBCTnZJlMh9KMIUgMBq/8A9sglL+oA87QcZGQQAk/uxsnmBW1
nmHf0JKoAEB42OQAejUsqNbBHEu9IXQOuyB3AA5G4Bfftx/4upSu6+tc5Udkju9R
Ubi2WOzuRxTc4SOm+MkOyzmiaIXCr6V3yQlj9TZzxFTEMpmVF/m7dH0ncctlXL26
f2qn4nJJwwWxPQlXVovWjrU3r7zULrA5amj1Gkr/pv/cYGErMDhFbcz035YZ78Vs
rVpRG+hiexfLxYGOYaJoRUJkymQq46Vjb4VMjumxpuZz1At89e01ADkg7GY6VodZ
8SUEwKYHNQxSxGRrDcSWMVEdVMmLsjEtxCecjv1IoGvUqG7BxhNmdZuWLDdvxmun
CPnMpdXzetLKup+o9tXVNtRzvwkSxw/Nb7TWEZaZx+E650WIKZa6iNFB1D0iMEJO
q3tP5ThvO6h7vT3ftm69kCpEXOFlkFIA2ZrJGBgXSLQb2Bs1wFgscS6yCptDMhZ2
+zubwtZQwz3yaLirvgvwedYiFKx2D0K88dP/Ildh789/de86O2fiXFIku08IRMa4
DJ81IKNL74qjWar4IOf/rPX5UxSGFpHTBWqzj+fj1rBWvnomHdDovpdwBfubBbgr
NorR4Ai3ATewz/gziZEbEhCD1vmmJgP/qCVcaa8kKawun1V9/MI1X86zqQZwInRf
AwTzwhgY4ig0w/SREEkAVcTBE2E7iel4wcjxf0CraKKopDq/XibdRNqqdB8g7QV+
30eBXun5NdXfvZwOokT2WvCOyVspHb6AqhRIg7N+DaWL7NNd+5zORW3mM1UXRfkv
ckXX7D4aJy7PgNE+Mi1thDS7ZBNsDP6Dizf67z+Qqy6EAR2SNn4FXE/ve1x+hUk6
IFrmhbTRJRqEmLbM2RGpxkynKDHcmMIQ66Pov+S2fJGU6P90/WSXlEhDflvc/pSK
IfzjEzR18hiDjobamvYHk5muRW7VvFktXKA7FvfJroNWeyzFRWfIWhDe5nFv6MQB
0RXQwhw0QNofH9aq+cpDx0lvdiG/4Eq2i+f27zF2s0scon5R9sRpMZ/VDoe7CimD
DYd7edXG2wTmbuOKs+WmOUBN0axn5TyxZsqaJTriY2gCmxdSOIcAYYK2LbGd0beI
SaNqDC1yryzNe9FvPba2zA8uFt4bSwl0UhSSAwGVBc7r8U58QC04hLAZVTyZgQ0/
k0RKSVCQDBawMMizhXo/IaHIgczaPPNUNQ1rf9BiPnLVBm2Y5pJAMV2ujMmzrqE2
NCQtAorhabv/KzjsA+Xbxh/l9il7OxoDgybBnenzwlaePbnHCapyTeKRr9o3lnbD
/VvD5nABH5Gd5r/8UiP3vwJ0/ChW972xDFIg2hHnfKoDjl/Y9bZ2RGA+MS1rWrq/
Xi9VfGvJejRkq44543Sp1rCx5u7MeGVsy3nf9+Xdm2CnKWq5QkFcawBcWfbQEhZC
E1DwfBxxUJaYCCOLFyYHZ6irb8HkNkZQFfnv2Do3uaLAJYpNaeffPKfGEjWGzs20
PW/POy4FvmSI7p7q0E39ANKnJqjazcU1Eb7ZMjlVXUsB3gbfiRhgWo4ZpRoOpBAy
m7ZgIi384TpT2LcmjzJXNDrtahnFP8XeXxfnYZ9Vtw+WHdfcTqq1bPZMybspcCwO
NLWdgoteEjhrB21T0j1odInxdA52F7Aa4AsQmCbhLSTfD+C59C3qLz3tUgLI3Cnb
D881esX0Vcx3OMTaRlG9VPGf01cfoPD1nz47cAAUUzX3XJu1t1kFgW8H4clbnAWv
9Kz6wtEJzRLcc60TjqlT2YmfrDPUMm37Dr/ZgOU8SRchmcEsW3SxerDdhPx13AjP
yDk3qpnlUHKd9RTGwsoKp/1pmCHk8/U/09RFpuyzSYz0R4KY5wNnokqRD7NWK3bi
Z/tL7NuYNRAjT5xtJehNVzAB/mbgl6W+e5a9ucjbrJh8hWDQtAwF4odmTEjaA/Dw
sRYo+Fow0EzEPmvWPF3OhBuciGAnyBPShV3KL7Dth65wzt/+YOhd8WudXAGxsf3b
qjz7weyy8jxAWx9YLWxuGUTKq35DlF8xMQNAjOEAxTFqbJ8s0Z0vypPE6IQCDUye
bLdzKmxpvVjslP5zQpjSyBOlYG3k8pcAZUehsKwlZ43tEkR2PXlII/JdJUthlJDd
T4vBJt1uEcQ1J6AEO7j12rs41VzCx3oOvwIN1zMlQ4zjBsnGzWVaZxMlmFs0P+KF
AFozitam4yRQAs1T//rDcOi/oWJ5Ecx8Y5PJwnSbkkNJgNtsnXzp5wQSGo2jSXxe
m+QBhjYM6IvTN9gpzmj8bGPLJi4FzHun4nSFXyXzSVAqBum8nyI5L1uBal20mVF7
SqYqGZvHBJ26jP42Pla5+JsFDhVLS1LDZQenF9k284kCyve0hwAo9TdtFxLpbajf
ZzP51tKeLEyzn5KsOwkZxOOLnx659YOq0tfhaVm23eo7+POd3Tvbuw9e3fM1Gy85
XtN7a7L98vNqGtlmyO8eYpWgqeE0fbdxt5VoI8ASox2qL0FiKR1XgJ2zOroy0x5b
tDy3zccJGS1pZqLZ/m5NI16UURyXUBu933EtrG2oosEO/UzETfczphH/SuMOkr6r
RujiSUbRt0nfnEvLdcsSJUEy3VFWnsZzHQDqO9dYr80GY9zceGOZufBtz7u0aqQC
B/x888T+P0bZddhrg9tDI9W6ynHgEvDkPWkLju7hyW0X6xEB4Ekaz+mUr6oYgspZ
GwqXaj0UJmWPZNpkVF35vUbkcLCcXIo5bbWglXkTk4avODXxatVCs8fb6gqblZxS
oX8x/yl7Uctn/CyxNxEZ65dq3shLXj6WlMFT6CBBt1Bxz+e3JxGsIYKuguWBTLIX
7BKxKVAu/ckkIrGh+VkomhOSJ9PZKLv8m7RcJyk5fwH5IoBEWcWEA81ilWq4jfI4
wA+uo6SP8UR0L/YcUGmu8sC7ImTQm8HNKg3ST7crT651sP/K7MASDQ2ZTTuDDju8
o+wL+exZKO/JlJF85RV4NN76ypFEgZvukWLzRpMV29g9JBIv3HAAPhMIDqJYIC9p
789Fi/T5zmRpNln6HTaIEkhK3lPqEkaRZQDzAvZsq16EhSYg7nXwSUXWiCAgbCC3
g0KA1+zUqgOLYK/0keqXgs8ajQgUkMF1bfrwkxIotFNFcDGEMFxpTP40b3S0l2Vs
c/xbSvS2J5PtlzvD19lLoL070I+1vnGmn1UhhaOjDC8YLh1Jthfz5TT+PJ9IcBa0
mJDXL/fmfbSYHc67ZRUIrYPhcjFY3wYQMZFVmHF5XGOx2yk1ZjtBGrGH8SN6rqVK
ziMSW7TRwd/7jcMLny8CQPTSg1dT5L7XMxsx//FvAhWRsEnHv5Z7wPwKMvouzGlY
HlJ9P7r18HCRWN//A3ztu5/xsV8VdSDFtXcjk3VHLOYyw58Z3dWQVfps8q/jc79t
wLnvc1N07rZomyl77lGQIG3iwJrveY908Pmx/uqHn2brzdQxsLmRMSlEL0jEW/WC
GDGu8E8LL4gXdarQD8ysxQ8UXHMVXUyDBKgI/T1H02ApBFS8cjDh9oiGOqeLu+aN
KaW42h3eg9Y0MRLIXY57GWnsrSVeTl5ViSvBjvt2h+R0uzhst9R+BlklGa7RH6YW
hnJZnpdgY+DFjLclwvAwoh7S6GT2kYUGc9uS952bxHHeq7uLOtMAM3stBsH9SfW+
/CNHZ76Fbg1Mu5mR4NKcgpbXQuhhC6TVaQRGpxz2yWjVzlHUZqvk9hQqSm9+wBi6
c2VJN0eGIZ5Ggm1gEaUnKWNS2C6mXZ8fHfJ2exjTQMZdi0aQhgGtLQvE5OfgFolr
jR3esyh43DWq0FXOLCihg3wU211LshonV7f42gIRM9WJAW1SdhvQ2j96jfKw3ZBz
B1DMJfGa96f3c5/SsZOrMXN9SknHsMIEtDezOYhQAnLEvQyb9uhSQ1Ud+c8MIK6k
C7Pc51zpo10QfnZDKwmfTOjXh+zLVD1uPV0WdVb9JjJ/d0t74/Z/0E/yWusQbqia
J7qxeuXb3d9RnaY1xHB8sk60B2zDCazEALT2qMlBcbcaISBnGhQcPlHeeZb0l+hc
gofFzwLQ2N7RSLwYgDS04q+DLiGCzR6PMOy3Ty3aIuBJtiNPv4XSGruGlsMn9Xxf
P01FWp0rN2Mp6pMWNHb2VeSTW62sQHtx3rahwPCZLTVPjL3jhPvSVhW/6EaH06D4
pn4sdJ4DybvdFjY7+eGuU4Py4JyciWwercikU3qGy2XiNWSN7ft3c1UzWV/7ChrQ
WG+W7xkMeklKjYSXFWQ/g7YP5Ufjj8+32C+Icv/15yFSXQPZf5P0XXBram+LXEc5
EwaoJN4fST5b4suB/1ST3Vd2Kcn4TcRJooK4fBUbnrym/H7yxkvo8hzOmCg9Lvom
AIWGpONQ6yu4J24za/V2ssjKrRV13lXTpHTAG/i9k7bsG++Su3cCognbjNH/tXgf
fvbMoHGHfhW/MfgDUvXhoeTRG+nIrrh4rNCXMLpXLIvvwTxJIp3jROsOAtoYbU+L
JQR/l2qeF2Gkr9+tzz7phoosHlMImZZnzbZEGTt5Z9KYThZDG9FJxy8fxeg7PjFy
1RpyhuImVQt6ia78FrzR9uvNSNzmBFvIHpUCB2OsCHu5+qbVpJISk2qO0u0CXwll
OKDvb8YRhGcb9wUXjI+RqZKMTVTAbXGPD8WoelhMoetkoUhmsN1ik6AkT63hB/R8
1x5YxVK0Ld1AYhvpjLAA8JKixFAEWor1vsSb7yNx/nkKn7qmSF8LK1HfwP3Yuam5
kLRWB/Zhxsd86Jz5TbNBCK9ZRkqJQbBtL0dDtpQm767ILWCAYwkup1wRy+gSaLpd
nINRJVMrK0mumiMsjA18xhXR6bekKiLrIQBoyS4YIsFZmM8JVhYgmmw/WoRhyz8n
K+lLc7Iq4f/Jq19lDmV3ad+mDx+umopZ3j1tCq/3439EdRXBoAcJuTOs7NSsQFac
FUizWniaj4NmaK/BAWCygILSx2dLDn6SuTHXPF7UG9uVYgRKC+OhZ4ydQIATXFg3
fiKzitvBgaq9jgbrI7r0fLsQbcUem3O3wHp0XKdu0iSZ/apODergLXHsGPEvidPg
RviB5zhltL/gXznGKbSbOaegequktf1koKAf504dL98QnkcIRk1VjnAUmiB44gS7
XKX0fOpSBuv8Syo4PNIS+zjbWQvGRGNVvbanx+BvhWwS1Q7zscUk3a8CBB6WpM24
fum1z6BVJ+ql32VMUs+NnMwcJGVUTRE9Nw0wiHRGnVEWqFjt0ef6pTxuguof2Tv9
OqctysWFa7a9xWqxSFRbaQgOQZ1Fo6vwgrrNGZs25MkD5oR9/Pn/u8xvU+43Xw2q
vpCR77r8ubL+SAkLPD7NHpU41e7wqTxOOxYYQaG4loOYJTRrX1XPzDZk8znzl+cm
Jo6TLv2NsUPOZ4HwRGv8oEKG5hxnyd/ni6Zk2sxrGoq5kxPQ523YBMs5Xn3d9rru
cz0NpLF8K8RnUDVP3ebxoxZyaVyD3SVUYF2x0cPNWEiYOynU0OqKkETUUgbFb8HD
V68vURs4yPtXGlJGfPhszGNNEytvufeR/h2iHEi9+k3VELFzNSCuHwjF3FVIz4mJ
J2XCKU1YgnmzUjNQn/6bzT/ix3e2yXmZqO8MI+xHFED8UqJZyCNjL3GhSQlptnmC
v+z57rRwbv0Nx07JaXEZOiPQ4RxS137A7jSCtwtV0QjeHDkGOr9OGTtxsIr7NZyy
5TGNNXSFbq4FYS2hLP+dd7QkmSIIfaSEtsA7u8eF2lzWRV7gj5O/NwKcFTSvZKA3
NzJ4WidXu/OkYicrYSmUqyTZ+wkSSUOW9/6WXLfstHM0zKpmgBOZjTvGquIRO3nb
ETbgfrC9hdaeNS3zoYLZmwY3mpseHigKfJlbClmXgHLWthBhvyvlaxShiiE6Sya7
OgavcJi0JImbApxZGio1oyj+eR4wLsO6SIVK7YP8GBQVhIrtfRtX8iWFO0I5aIto
ApzrjQTt3ltB0edbdA5z7V/QPjsbpMRwml7wcNk1Ja6BNkt8vIjOn2IQTmTyQI1z
7n+4PWNnTKmWUT87U1t2AN4SLKGtiSnm9gWPc3xuQWwAlc7JCgTly5/jos/vIGCV
Xw4L620mgUHHIcqX6MljCAslAFRgUepVfq/jQrP/a4W3pR/age4wZcyIxsr2bxbi
mXuvOm5nLlQVfxLi22JiY+CLe6fHeoKEgsHnBPFcwPEmnoJ3DAjpFelZ17t+i2nn
+292MKhjuMjxaIYS4udGFLZztkBpGVWIqDkY5GOY152cVqCATtVL5aOqLDdXSMA9
TX2OOTdqeqMUXR2gryDaZ8g5NfU2PniGDvhLsKJdtlUAONcSA2ljd/AXLVw6swOE
SlOUsExEJPtQGHd2OPGgwE5xne9YRxx8nZr92xJzQjnGTalCgFWtIAgp4clhKaf2
dZxwrMAgpYS6uSy/xmWr/z5INTXvs2lfKSXg1QpJlqI3lD7fXxyi9Ux2NR2MHO6p
eZj2TYKEBg/6Tvz/t840pPDXYOZNj38B73Ub7JV0C96UgNH/lIjNyDOVW6IW8+XL
jAbSUxVB4u//nEMYzaeOHgeaRHg8Ycb1IEddd/7Grre6ym6at91zOVxcHb3JCgOY
I27AT00vPzil7GmZ9uXoW6wrcM8Tz2/k3F9d9xoeDapR8K9smXF1XxPr67Xjn3Hx
FE2vqRzoOtiVV6evo46VVgtnltS+GtUOUUaOS6kmQ54X7SiOKXy+w/lovq98aBXg
SLKHq6kY6RIu0cNvBxoXIN1JJeaLqV59Ib5Yq4gOibI0S9g2XKO+WzIMtOXgCgSb
vpCILtUBkOKaDiNEAelMKDxPDjUpV5xty4MRO5C21lbHD6yBfy8DRvbSntSpC35u
AXleB8mM4IiOrUACqPkl93BmSGnWqaq/9LGev6G3oDGTeQ4CCtraTyIjQlKfa5Mt
KHvARayZeX6viABbet6yYu0aHh8kGyEZpEhUd5YQ/9w7NkfjALdNicbj7lHZ3ok/
tlBnEeowip4gjltHUiAM1jqxol+rv/5yVlqoA4/+cvqlA2jLWU1NgQAxTemgMxVm
kEfgV0hdpsYOOBQ/rAe8x/4DGGAlrQT3fcBIOCCyikXSSNEEWoeE4k7LQDyEJgoo
Zcqr5Q62CfWkYYakf7WFYcZLP6BG2uy2uiO/W+Ofu4/nJVAbCspQGLmu8VQwZ4Rc
L7MVFcAxUYl8pb2xqn0dhmAk9SngMCoEAkl1Wgw9Gc1oUERb4gdnzThFTHiH1tG/
t1+5nIb7sq60EJDiyhNn9n2gVB0nXZV4BGdE6knO9dLD47qv79qNJNIpKt4I4L4l
HGSawI/YDIyfTR6o80IOg+hsN22vJRAHvqgLbx+qMFGyVsfDVuv/6g4Ut6Jax4mk
pXUXjYew7LJJuJ4fPPFsWf0ckALettk/gMpjP1nKRvdqnPVt8SkwTJdeXazHKKou
86vOMvVEcUiHs92AnhzCbiMqcVrComRd4J3hFXpNsfK7hYLHBOQ6m2T4NrJnQT1w
hi61MNqSfH6aCfGaIQK1gOsBrzW9H585Bts0fE9qSrg6LWvFaCC6oK1W53UZgvFh
SbBVfLKwjtZUbC3gHPMi5ht1YymeYw/kwcr9Sb92Buyp0G6MtycWNoaqnvavommR
cuGxyboCCheRpVG0xKKRKU0N7vjKyAplVVzF7nmAByYSpOM1azi6bysDG3ZXEylL
kIuiZl5hTL45B2BnQVVSmhg00pa5dcpDwOZPb/j4Lr+B2+T0Nme4CbpV/EhWj6Fd
og9MPfAGgLmC/FqAp69Z9n9hA3eKU4uU48eQmbpfeAQD/w6FZmWv33rndXoa0B/5
2ttZT2pFYac+r+ijqleL7ImvPwSmz04U1C7rMrJ3YXhjt/xXWb012VdNxVOTMsDr
ZSORpOJkp8fMULp3HH2J/TzmQ26EvqTXhfqr168XF7PD5Tj2lWTjsSyJjTnVq1JD
/kq7VyY3QWbZ3irUMMxeo/KrRfCdp8YAaj8CqatIWCNlahgTDMbDtKJv53dsW6BB
UHjPMAOH9nWD9g0VyNwgb76TiN+ZN+b/zXy9rhyBn05ME+8Sdkrn28eXGIhX67ok
wSwOUsAB2DVDdXyCvGl0rOGnrGmACd3ES6WGTgMYmplAi+pVq/k2zWTQ0MTWbh3K
LCgHhxdzcuvxBf+n2l5Wo05A9A3nQC/BItF78az6Z202ncasCn2cAspQTtxDSbdh
mt1kh3ZIAmp697xrxBqsOzaxceEjKvpgDWwsB6RhqQb9ctSPLpdDFPl5711ZQXG9
rrkQeppExvGN5QTd9gixsppCNgL1flSiDguwOpD7BatfJYPvohgj89cPTNpZ4Kgm
tlbtcEF/vMR4RJcKHrr2e1BG+bMJLVx4ZSmPs+2laM+3nSNI2m9Kc24p2Pgmwc5H
ZsH+CCp85HtE4MANtCQ2YVWdUFXoKOVB1NIAgr3vjyRz/kWjy3nedUb15zbybJwM
LnBjhwS1Qez1LEML0I3k9eLXlLPzzr8LZ4IuWC7aJ5OhTQcEix7GvWp1dF4xzv2g
sWMwMFteURAzOj67NWuQy4IuXLVY9Y+QPXVRL2zBnSAqIBW94domdynu8RLDU8Ws
MQMV89W5cgE9VV1k28y0EZW4QT7QNzUKf/RHSqvWL7GdgeeBzPZq5fQcZguol5S4
Ucv+J1MjC6r8VBRYMvgHvqQn5YhfcCYXnEer1FDlBIno4Ihey0WAO3lJVlE1rlKt
TFU+2kDmN15DccHCQLGJTO1HkHuS7bVNw3vq7h8GNjATpixM0DXIfbHKSJa9FQq8
+iS7AuVCkLvHE+5qFpqcCD4rG2i+n3Q2r3KhFsz8RBqcqYBcf5DbSezLSh1K9eFu
uvtW7g+GmxhVhT8qM1IU0ChzZwvWFuXvE/kezE4IRT2YweS4KCuopP+Z12Imvg+C
5o8j+T76W37M7AYP0L+hX5/HeqtqgDMwbnVQFmT6hOvhBOh3olE/JJcS10TFoPOU
MFVcf3HXlo7Tct6ytZ921lOAvEU5WstuEqLQu8oryny73j6o6CBjmh/hiPQ6PwXY
Ox8SYojHTSqgdkNfCFw6ZVjoDmr89vJ9d1weJ2lKf8k3ZRuP0zRGmYC3WtN87voR
iMpXoN7StEtQpy308PKNELdlqbDbGPJ9if0DVym+kBHJHJ6yGeGEsiqGh1mczi5P
QgGt5d+Ff5nnZ6LtYGqN4SGjJBaudXlHvT3lMWUqCDWz5okYSh0RpUBIW6CYUyL8
uAmXZFHVG80+Nus+lS4TpWDJcjqV8F7oTnLwKcFnw1nQKKAqH6tztSgQMyPgMLsy
duFGEK2tR938AqRFnRYYHMxEDe3olCfsbuAOEx6g6cJIJcl+A2MG8yktxXX+MYxI
ToGyRMJpGX6ft4xi3jCchy6GwnQFR7bNSruRiBXp6i2ygtayEmV+HfJorLNm5fu7
Z4C8tYsia0PIePVKKEPfn/0BuhBds3uwFJpjUNpHdVHOdgGZTJo1u63yzqwuk3gU
4TlhMqvjeuGk0B6lW4O/5B+M2IhDM5kJwG5n4CUMuZaZP90bTtd2Lbc1KpsUGbpp
B9QOxUy5fu2Xf/hy434DRu4yEcW9bMAxv5di/qpRYnU5Cc/DqAz/JwIsmx0wQdJs
5A+kWd65/c2EKdpHdRQhrLrN6LvHkDgU3Woqob36EZ5eYoEfvgBANXFLZ7fAu50D
aWuzSyXxhOf/J/rfGi7To5VnORYMD7F6PO7K6BuoY59Ckp9YLN1sE/CFCum0FZYa
Tg1uO9Xmt29wC5MdsXCSHaXk/N5GLjsOOKwqS+29HZ7fdV6ygt0VtCHQMCZjmdRi
+3WT5HO7W2OswNjehnlkdTraM+7AiQFu4Z6eDpDGBZmPEsrsfu32qu8nZ87mPiNa
RM/4n8tu5DbFkDLSZgu6wQW7DD/LVu4pzAiqTxc0j9xKX6no7kc9Ku2EGamETtyp
WtZQawcsaIoNbmVjIqbUZhbP3qMl4l4GZFEaj4o+jXey1TNOhof153dHyfG8VmwS
B4nWi+yu2oL8VRGo60qe5cNtlSqR9m66VH18WGAn9kHZzdghJbVb9E/rLDCeeCin
vxRLgEYec+iex5+EeFnfvjcT1u6uSppVL+4cMmhrMAzAnn66+2cu9+cBuaPI/7p6
VuzRqSZ3xP4mJ5BYciBy4bGYHaFF4jj/OfSidpmus2uDBe7nHUbdmCDTPD0HzEhU
ep+LGe0qaAs5fY+wfO+0P6OSt9MCbwU6yYLw61i383QH5FiMqX9bF53uGQqeLsfo
qUD5ZAabSl0JbEj0h58xEq3COiA5HOBtsPcLm3avVKceM4XC2Au8Xj8JpHJq/glr
Nk7MCguypITTVzawLvbHTDD9wr1YlTY9BOh0FEodWTrStzkpcfwl32LCHwymeAlD
OxXDsU5W06LOeyBJh0EmYey7fnN4+pCoJzr1xGk6cel4f5FNPCNxM04M4DdgIw1P
yMvARN6DgnFFvf81l//JRYS9WADflHdizIHzQcemAq/4RPlWbBo8u+dvb/+NCp73
dJkUm7jlyDzDJ0R5qzRpXU/nwB9iPPB3iGH2GMBfjPOyTgdOrKdhOJtT5eHiYly4
OV+GgSQZRmM8JFqtdukzhvSYYXYp0EvuxypNZeS8LwrS91V7OBiTj2vHDRMhaaRm
pqFrjdoSFFYj7Jz9woCIPLKKl+NfU1Z1GGHThBsIp+v+UBvMhjmQ2aArILCg7ABh
5Bnflet7LBKwwhjyavi3pIJ6aUQM2Mf5zTrg3OLlA3c747hO0yK1VbBRgvT2lVFO
ft+XwDMr2LfP+VNNXGpjwv18uWV7Qi73bE3Xmq3AXhxN8E8opj6RltCbczReUgp4
b2Ls2xNURWuPYuti0W/gD9oDBeCZl4p92E5c3kfp3p5AfobsQBGPisqjXmQnJICZ
koUA8xMkSvtNJG+au9HaxaJ7rsWkHUXLd2HEWRFnvkJiWbNklxZqzuNa/o7uF6Ts
OTQmtPICh7CkWPei+24QA58QeFAvA4ugIm5Y2Q4q4z8Kgll9VFZeXja5TyjimbB7
CHe9HUXVdVVZSwRNQ088o7+i6IPh1WYI9TAyeusNsm+iZBCYHkR4ysa36Q3J6XsN
psxq9AEkMIA9lhlgRFW2eKC3j5sHtIUnNB2NlMobC/ywRZzL9xp5WDgRyP6V3qjf
15fxOWhrcc4smyJWgTk9Ffa6BIiit+dwsfOt/tWCk+0VfJJMRwPR+gUNCbotDKWv
Rsw53IzhOLmES6wRiLvN2E4GKhgVTHGj4VC1jpxynwI5ONPpHz4tPiQptTQG778F
bLtJQlNzAY9OofOoYU+xPyU8397xJ/2kd8CuJggzhiwBB2CAVU/o4BzN8Wgkww5Y
n0A4Y7p3afJMwvRylQbi79eKxI/3PU3RSgQks6fjgEwPUSSx4VvGlk3C/i4xc9Oz
84VgWENY6kvvY3UZl0Ph2eSfNWodOXOCMGsHxTP0SPznH6fBKewNUkPBw2iTI72K
yNOsz6d/CSSz/2KVdVgT27d8GlACuydSjCiAbZSameNjAOf9B3rELvVNUKfm06Ei
FNqLPpB+KFIifZTYHPP8+IRTXLiBtCI++H3aEK7LNgp5YFkh1I8b6XVqi6NNtSV+
WYquc4M9ClMWWcLDr7yUMaU3HF2zSyO3LLrnvYh8y2uccSYsUwu7bVuOJBpYPgFu
S09dWwDrVyPzLc6Yvhr77doStCyUmYWvBa3VQWTur1FxxqXcAPvrLBv5O2DShQ2Z
oqdcyepOJ4lf8l+jnoKMJhmuIGJXWQg3+fD+ZhZTBXy7Rpqor1ZFBXfuJMXbK5Dl
PmCpnVZ9FdaAvuiVCWuctM+J508vUsx35tCpH5oGGJxKiuezippWHLHbBb4dKhEf
JMVLaOU8hfs0Zb/XLq0AmgpHeApQLPC0XevTYI4r5sgcwp368K24DQLW7pgTPjiw
xLjBlah4+AWZbaqCYuXIKy060ocUQOHjpYbYyB0zMdjGjf7pBQNMeYyXkmFkNqd7
mpG2HJGghksEdtp8ulurAUkir03qGVTwM4ohsJjhdz7I8q8Ix7oK9DFJCRH3u/qg
80O1vlPxNctIVBiWndm0ZUAX8C26n7Swid5SkvkhaO7h0g0qiwPnI5hpd+ge4/58
ePsCpRmZKzAMm7owAtwgWgbGP4oQEmKPceFJqkmhNjqK/FQyTqFBk9o1Jui85ltQ
x3SKofjP2Tzf1O/wj6V6kLqUSw1v7p5S2FE/S8OeLw1bSd2DI3CSUJrU4T7ndRoB
ESgdb0Yqmkx8wsSV6QZPcu9LdyiQCcx1n+dRPzMsh6oLU2hDRY/ZcQWe+rzTSCu3
Th4smqenP0r41CmZLElsxexQQYhjgnUFtum9vJmsiRoIdSYWhKlzF4yQFAJRYdk9
O4VvNJOdu+55T2bvjxSP08GaYfbznrSSVlHPy70DxPNQjye763YsoYRSdqkujS41
EQiGANEmYQmS4h/XfZKTm+SsUggmML6dxl20BF8uJ5TWzuSgkGlE7RKUPvAJyf7n
lYX8vB2Zwz0PFHvYAgGo3tnRUg1E2mIx0xC/cuYhXUFq8ZmdyUBGKjYYNQ1FV45s
aUVK37EfO9W3U0DKsTedUBfXMsEMpQuk6h6PRjfINk/uI+S3eKlqd3EKIahNdNVV
uo9ivuZQJrECW2EEBr6y/1wMzFX8z7JViQ9d/sCi6fMV+8S321axvxmr7rm6IAYX
HEHPoaiM8jub2Mkn7voXacyJ0wfclcznylKw8aTHvMX6NELj/dsrBCSASc2KrtxO
ffLXcxEi+3hgdfk/yevqhfkM54SRdNTQV7LwdscXrxaz5wztRRpwqMU7AEKPmXXI
Y7XuEphzamIzJ8c/Opjz0YpbRW2lwwNskwOKBsILN6EYFUiCMQ3KApoJJ9sxNBX4
s3mZ90EgdcfqF1lWRsyNPGX7JCsAVzGnvCP/cpk0r8bBFFDS/VtLD8LFZN0A2zR/
1jyetcpeJu0CVSmua7VyOBejWGHNGkr7wYvs0ieJeowFWk4TLa7QrTrMmxVMewXC
ILX7X1145/DWEwaATlaCoQqWM5yWfnUJUbMojhqzoP9qXUVnBVbdd4D0xvAmKfLO
8ILKtf4BQwm9JbDKVlgfxKZAehUcK1f5pu7aW/XJBAEXhnUNjeDuiYB9LRtpSehX
WzMU/nFY0ibM6eoGNSs66HYm0Vsa9uSY7BNwGtcouKaO1KoOkyqJP8HwhcNr0Tl7
8/XRWQtIU/gaJE5c/miW3jH0OgMARamn0nwpva2HvX54RNzSjN0FuuLKKRdwKj9K
zCW492FOy9Vk0YUPT4xm34r7MlUUHul/amzR1mM9/42gNOIXxTCb5RiO8LJFcmq1
nXXVe2ow5VJGJpplPWoy7p253Pojuzpr/e62E1Etpa2/2wcnru2HYNsrencrcXkH
Z49/PzWtReRw92NnxD6ch+1WwtMbU8P02nYzHRhMngdjukN15xpAoElKUrYxAT9F
ZEN7vovr1O7Fa0kEF+iEKGhSWQIvG5xDyCAJypmM3T6S40krcC79U3sjICsfOKTL
v1jA1svFlxEvo+19im0W9kFG93NbxRNi4oVWMFhziEo61Q45VEk5cAfBjNYhzE+s
tgNi7w8b6YYakpxsdGGc5YERvsVDLe5NU37weSEOjBqJ7zwSSBnAg2oSbtuxXlJw
0rnirx01waVPdC8DBYsLl2+i3nBWKUV4DptdLcIJkzyy6ZLc4t5HKtfOyy+ZS9+8
gQVEu8Si+NRWSKfsHQTRs76HaE9XyBoKs+1WJ0O9dUyxqAVv3cFcuJwfkwjCVxd1
2N8Pp8L3jobff/ltqzwwWrGSPhrb4BfNiVagOfuOZVHKdNnH2Qb9LVZcyCmdkfBr
Xah0E5U/2vmEGj/9C+ijfvqc97TSIrb4/rqFhItxtw1UF2NCTx/5qSrApNbyY0HL
KErdPBgX71a5vWoT66bXUFEQWQwXtX2aRAOK84E+f8zy8tmvcUEyf1xqj9sopZ83
sVwZ6nVT9GPQpL7TFqdi4FI0AijE3YAMR/tgzZm3+4x7dwF6PUngqy89LVDHFAcF
1hrGGYqcITd/3wUYvN2+3fJlk48vBj0uSpFukpgo3+Co9ltEiQvMBPdjVsXEfpKN
zyUPCbAjFxvwWuEHhNiZBIMHqXgXFfYjcD4POfKYaWya7f5VULC1Uv/W9JD3P2AF
986sXuaDtP9tCz6ivzZd+paMJap2tY4iUmMxssnqnIcXvToy3qT1Hea+QyqjbnSa
/bB07kcZHqvgmYvK+IELaqH+ozHKvk2n0HyG0OLHbpYsUUZsb0kguyEIJDCSY9Fy
4Vq52xqVtVDjUGMNdNxhZq4XHdjMXyswvIbxrDyUQg1xk66oandhKzBrYrV1oF7Q
62xjtndGPbQy3qPlJQuStVUroxhIdqiTznIHfcCxXiwrsX9WQrZ5qUtrB2Q7MtQy
AMRNs14taG9a4RspVfonoazII0tB/l5bAo9xWGHdUIZYltspKiPy4rxPe+x8Hfrk
ZB+6ID9EOhRr+5JRjJVzLm2yZsuIP2o55ONyQzfQ6BRPwSi6toNHLyG33n+nO87+
weYBGZBuz7eLnm6JTSQ3o+7v9oHSvRO4UtLAKsQArAx937b3rHvvOr6MGCK0VpSP
TQ8LXjcyNdcl53RJRRWeQEfEeLLVQL/gELV8cUUVcZh1EffFkVtkydiMKM/nMM8G
226XiXa72w4y4qLekcw47XjnrJIBZRTgeW6u8PJuTQngWqiKkSnqeziKHbow6OdL
unmQEVJhAiqjPPWdcUCmnUfh1fvojozfppVm4DYerZU0JQVhT2Belsp3ORFp8rIu
oz5guZK7pP4+2ossLt3Vb5Ezc0woOIHHDoxifSIa/KaNv2sT/uDDkp4t5ewFFMLD
MP+kk0Uq1czAQe91ydU7jTWEVNBHVzt5cTB/xhoHgbZuQCt0o73LLfmkWkHbqrws
nxxGpEKSB7to54HhupoftF07/Wy2APYCVUfzX3h3CoZoUaOxzyno+fn0Vfebdcxb
4L7aPDYtxjIcN+peuHlObaDy+EdPtByjiWYPgDEG4Ou0+y90gE74hI29k4EJpVbO
iz0eHrB1IbHSyq5KKMf5naixfhCsBTvd5embPhqIKQPKHbUCxSrXsBuYQ8y6l24K
pFvF1yo7zrIZBZIPSgXwsjrIngBiRZpIcAdArM2ABjUm7VpIfhuj/2BjiTlrpPwp
bizw7oQE8iRlVfbrT/67lqL0QrPP81ojfME0x73M9ETU4vt1mr2l5EetzlwQhtA0
t6Y+G/5GjEEAfz2V0zRSgJzoSNXZmYsSl2kxCK/RM99IBounvBKATZdV72hHlc/0
rvAXqPkA9zYIbht21kCfnh0f9UMTlYx2UmFvbGwzip6z51DPaAHNV+OxNUoibkAi
q1ZDml6IBO5qDOHgOReszeArQMySr0RAmxkp4Mpem5lNlLLDczgYgxf+uJs6CJ4b
TtFIvGY5aZt+wcieouMA4qVc1MWNlFVkPrV/MawwkVAjTDm4mOt4kASeU2czbD8n
o+whQEAwGX1kD/Ys+0Eqzmwz+TaJlwieMa/2xWfD+dDua42KBDU9b5CN4QuhDa6T
9/wUluE9MMUph3EdrfBahQdabIGyQ+efJtT+NYglIT+x8NUXuGy3TyZyIl9S+C8x
rUtBmJUvyJm01v2nD70GD1g+16uL7VxsGqiPNnnr4/ASxySGs5hyCuw79p/3p4XL
62VXAbsuYzFNkYswQN2mtZ+ZdKqwJy49CghWm5znKVMnv/+EbU1P0fENl9MwnnKX
YYzwei/5T2zPFIv0UlC7Wr+/oSDtUPlZ5SPOav/p8yLYtbektxpdBnE4R1lkROOo
Kx+zMIOdr9904UKUVzjnNjTGQd3jxW/M8Q3Hfpay8aK1VxnOz4By1KLDYdz2Wt5q
jeQb1ara68Y/hqR/NxxOUMKdnq0Z2S1X1CgHMgBu8amn2j3K1XIvn7R3L3qexDMb
SBK1lf7987rZTRBlHGfNn95M6/MX3x95zlOS7GibKc10adh7twmrakf1bN8fdHDR
3LH3IDWX3LnALr8j9qHx9gsSMjdMF6lK4nqk49e12/D5+pTSFY1U/JbHEXMz0GDB
c3p1GiUUYXm/vVAoP4DD4m7z/GdHxMECK6Rx66tWFIhEymsLFcBafHy4RTHZnFV/
bDzPKBXQeUOhcbaA2vLezzJyvSMc7sIdhaDUS6Yakknj6fyL1dMHSH4e/tXt0FTj
QDUnVxoZgVzupYY6bT4KnEZAaEt5QNjRb5GFcjtz7Zqq2rkvCkDWrefkXwJHVhgk
SU3t4wGNWIorL0n4Th8o8gfpBn2plIetG7U1fPhcoeFG+rzrdXjVUhum9D8tketW
fc9vmOd8ety1JJPXrtbMpo7Q7ENx20Y4DYrpNputZP7rzJ5WgWpGBhfSKKl/2qj+
ETq23U80Akh7JBpvYcgEwOEGRhHPMSYEHIs7WoOFaVoC3+xy85hadO3BG0p2E+ad
XqxGTVX3OtHX/r1yQnIYjuvpDOXh9U2oy02tnJjrHxeuNqZ5ZiX8GUC4GkUdbY/q
GzFyl+uiFLiTrolxy6aKVGacNTgzvXMRZO6fSIqR5qGAzKrxmi65eA+c5wiFhkUy
dd+Zap5cU7jB71t5ye8X7TuGExeFXBalWjBp+8/sM14h4ynMKwc6oT/EH51BLCLF
S3o/nY7aWttFd/G3sUH5DPMjDdry2ZaJ6VUHwn4oAoaOiFM0rRTFiwsM4keqQBit
ZLDk9S3IWUhGyEDXY4FVLNTc+7Y02ooBRyg8w/stxYZBuvK0Cf3oxn8NL38yZVgL
uCQTZ8Sj/9Fh8UcwZSfPWSIzlXgLVItoPgVWkleBR1RNP4qhTY89hiFsnhG8utnD
pIjh18spLRilJhWI2jqzP/t59gYZ/jPVNPPjrhucIOaweDCm1YLVWZGowqiWXui/
4LUgt+WE6X4hpLGZXN1oGrUBI2+TnEpONOuiGvbBrNELD3glzwkpkdMx7dmf7Isw
/xnLbaZ42m7PgTaHYuXZY8rgH1E8G9Y9IWPwUYPp1ZKvOo6qsSN3AW+2sh/oJlWl
iXebA6ycUhNtUr4nwD5zKJ98z/nfhF3knYFcrQcwPu4BK8QKgzKzILAzeyUzAHkz
6x4KsqTo+N2gt56KioafNqZKbbsm1mxQx06otxU17+xG90KfX8sEOCyFScfGybtM
GlgDC+91XMCiolRYNwKwmzcWDggzAz/DUbiQFsyyVQxf5s9Tn4RuHxKa52KGBhQr
LM3MqpU70OA7BKsgDYrNgXhUSxZ8AeUAIzEdrZo8+VRzk3tl+R3eSampIkcEnSBG
FahhX79Gs2Szh2L6Eymofvfj4N7AHa0RTerCT7Aeh5NqtkinrD2Qh1bIcU4ItOjU
2h2rNn1pwLsnLvp/VJGiHXYUPSs0Jq0DJGiktrLP/bz30lVsjvcWVzl8ADI7IRCa
DT4kPoCO4QJQ5RnfPnG75kUHXeY8xU/9BIaXuch1P7x1TTgavss5xPczlpKoDfXn
n/pkjPxOoXS9TIuvoKDIxvUMXPAJCiH4vhZ1Hm0oHqapdKlnmMDWPLU09WhF5E4M
D66IaX5RmH97fbf2wFMEwsAIOdK8taUWFN+Kg6rQ9shQ9BNh3BgjYQKV2VeZqbSz
9QBmgfmcE1aDCLkbrLwdRYM3SiVtniaKiM/7TDopUCXCyJp8duwaTPyxBna9eGOT
0Ok+rBZGrjbc0pxxIZxd7yX/NT4itmA8/nQ/HctFnv8RBWHC9RzkzhF3INGE37uO
MO76gF3gM4ZHi9QL8JSJQLeXcH+pqI8YHNfRo5XV0i0IV9CwGMlIFCuz6tkh2EG5
8Rhf+ZfiIL3cDYZiZkqPe8vvP6oG/927L/VI/RgLu+2DQs1cSf9Xfjv2610fqy53
XUvTP85G+3ayRG8+uDWfaNEv438ISoipSngbeURnk80iqMU0SwuCDn0V3i7M/j9L
uCXz7ckw0liKtQzhnShWj+IMCllcDD2sYsJBbab6k8DJGH3bv+Bvh4bIFIQ+JYpt
4ekULfQwC5XCf7Id0sQiXmOsZw4nxbwxe/tubtxWs+BeYIh0seD4g2I5bOV6psl1
NL9EF9a0WOMh+/RPPwEnbuBzBu2cM48Iiuh0yNqrIhjmAonwa3G2N0gSi4cY7B83
cdo5nTpewGCBaF9eo9abI38lbpikQt8bp0Xk7Djx+D4nGnfFEa7kF0HRzfk2DbEM
zej2hFfSoRLmtbcaQmiYSNYFgdC7SNs1/zziHFa9PJonYJojSMgqWIkKsV3ruB/v
bAJrUdjxuqntHeV5cD8X2PNKEkUItDGob9hziooOG+pnN8XjXY4DJVCOXMG1WAsU
jqQ83i4uQ1laahZ0D3D0KJNY18irJeZifs38/IKZ2pS4gM34Z8cOPNvR8c8fo+Tj
UpFzz59+p/Gxk6KRb6EMgo/G6LblIvfHpArP50cGLpwP9JAopxBZZTnDaMwMrxlz
/dklGeE8O6NTYv9xIeGp74t9Hn/W09QU7VQ98pAx6zy/ob0lB6dtxxuZbMUutWiq
h0QcN3DR146y8ya10EyF8DsMPVSdED5gFMxYZq2MJHyOZeeY4B6tFS0ZhGpUVX6h
g4m/JJxoFhx21yhkEQsQGnhT8Rt+jmwXKLGoQKSe2xy+9DuG93ltWf39NdlE5FVS
xlce+TvuidTi/2cAAwRhkAnb31Wbq5wCNVifMMPDnxFKJHL6jQLUK+utFQ1eDyJK
WkJeaSAQFnER54qgLmlS4DWEbO7ZHL7ALsx8gc8AC5l4KAVYya0GgC05U/VcCl8f
YywNLr25mN2l0Q1CQto9V05QXJDVFFFjOWOwiYnHg04SkxxBqxaWyg00GT2RBlat
uPLtwRGG7u3b/uUW5ajOmWIOTlHjCryLzzEmWc0NgV45AhR4kiSPrtUSQzLA/vVH
JYmmOkQhFxkUQvT7wJaI6pk5knRvqozdO5FXn9cKfzOEl27qRF0ZDtKRpSr4UOEK
NhLC5hFyCbwmmQOzmfUKgGD2J0ZwqK4XVTt42At+2bqRp5iRUVerrbHrjhf9GkT7
JpxnjQoSptAPid8n81Y4bpfo2biiooka3KebN1z2Zf3c6fiLKqtVkLUpnUuiz+3X
H3ohpe4VvuFfrCmNHk4/L4mRb0CZ5PdTD+Hr7ur1HPTmNNKpaDfMn+kPQ0iKaX/A
KzAK1y5UijOlyAbkv8KBq+4L491wYusTKf0EV8W4rvO4Z0mVf1KdEsnw6gzXUneo
MqNIk9wNHvLcrftE4P90v6Ce3GxUO+OcLOvjQZdlBJO+SESfm1N/Xm6hUbAvAJhC
BevsFDdsbsxGUSTHwSJzoIprfurx84BvjTYaguvdl1FaTXNKYqvp4uJ+6sZDlWKO
lTjS4EAIJl7VfIwauCCmsTOkjmHLafr/kBIUip0yTZAEMuxr3p/yO2XkckCpLs3W
D3smjBNb8FmPX9XvIFBavPbmet+DQARsl01qFO825SrlLYinBZSjJUNLRebQQN7Y
MCnUiyWS+Y33hcO2LXLsCuvyi3ddmbEdD7Smu9+mk5tGPkT8fsNikH+TyWilrpj2
v5gFYeLKlklTQjolEERpNgJqBZ/wn4mjk9brxVrpE1z0n/TnwNnzCISH4l8Ksnkx
6iDZu/jeO96zbMubEeGtqUP/AqhtlIC4m1JUkAozlQbMyG2kd5y/AnDnX8KiDLLt
iRGWj0GwbvdNqwud0wC9gHlJLJQrt2GVZiREkLTiuCxU9NGctspO0AX9tyR4nYn6
C382PBjPDvzRAUUzu2njvpG+zkt9tuDZPleVQu1Wtk28bdrtXNAJa4ngBFblwds2
PISg7i4eE+SzNTK31sXYhBprQWOgr+05f2+IECI8tz0jxoWFHjkayDmLZ9ubfdYv
nFn/ka6Z1XDmQ7gA/7kjLZ2lxjx7PehbGqry0AMpM10tYr5imRJUfaxT8mqxKBgS
iQgyqKcKXIzGliZMkuZjYczCmxlRU8OP1Te1QQysweEAsbvc95BtdKjdpYtA3Fld
k7kal2ppGUb66e6SQocxtaId7eh/jjj4US+T6szn7V+Dg084RO/xO3v86yHUIJn4
XCmfuor5/nI22Fs69kFvXCgSO52r2XtHben3V2ldJfF1h/FLRnWGd8D5tQehDKiC
63mhqaCqwPnbD9OPZHXHEb17ImrpzTHdwF1+EtG8ePNBAYyHnR7V4ZTm4QvKvXD6
T8NJGR6D16gVRWDl1Mqw3/l4R6nij643yhQp9Y+aTpt7Yabyvl987rlcBM5eSSgQ
AxPVIcU8P4Z3CMWrsGzLUHDg280HP1blxydn3w6v7vGd3TgC4psQDAr/FfePgk+B
D6cZRPnD0qclQ+VEQ2WsG0/oq7Ub9rT7ZJjdZvUlNmW7qGx7TFrrHpMevzCeYvy4
GhGttTySPJGT6kxedNMFLsMs1/X64yVmBh92Pf+5hMvN5DBQg4yrYjcPQS0z9un9
wJXEqb1cbYx/n0P0wKfjKisjZ/LjNXHqi0Wx38BJM1pbW2YQHKWSRVjSwIGZsS8s
ShC5ILgyS6D2uVuLoSrmWHRAT0cNHZ3T4Dyf2lItYj9L9sKp5eRA5AxYNOZmOlJg
mat8AitZX8FAgqUnP2OpHovBm1HhfeYs/6Kkilzkw1gNN3DKogNOc06k2mDLt/tu
KezYcb7e6jrLd+9vgn2JIKjGTuvDX4sILohXgUwp2noc6Ku7ZP7gZ+0S1Byt7sci
HBuJTsaakROG8JfI/aP3nRKPB8xlbNpO/CJdkf4ghdHZ2eLj+UjAPMhjxQB1Yg/r
Ev1C8aMWiLhyRADF8vXJ/SlPfL278luiud8Q5YrOKuHPzgfNxOh2vrOYC5QQHh/+
h5mex1E/bCZzp0jcSfThmiq4s8rEAabVO4uGFLCoWmPK3J4bqlsQ+VxPpxudh25m
bux2mu3INMcnx6xb9kyqDRKs0LgGjoL2vVw4Vsif03EQr9vtallCHhtVWkTl9/8S
Ia6VHtDehspuSPs9KYTxcdFzRA+RVn5izqr+1ojdZk46lSqY5upK4sF3BmK697Y/
pJtArioyv/zd7Oy2lmxKCSt69NT2U9jbeXx2SDOJ/gYFDlooxu09ECKDriEUasSR
cXmw1v6bRTLlqnt3rbIlDAjPDAt4hHUKBaj1mqM+FnQWRzsqi1NOplpduIyfkS3A
+WZ4ocdf065kcXrqqNMJ9XCbMnmcPgjM+ts8W7vvPsXDqpNoyEm5SSuD77F0t4eY
mxvUl6s6eSb4PjqPU+QI0gyDe5pOXaJcVj80wBtK6XP+CB+mAlVkbRwSbZebdob1
DlnfwDNOd7vYc5ZLoejb7GbiNummU54ZAcwSBXuS9laKQFrGnEG8LSNVPf6mCqxe
HsSd5EDp339Ws2bSFNIuKfIRQ9okyE3XVFVtQsB3oGFqmkroe7nUo6+KsBOVI5RO
NNc53OlpYgcwVte6G/5McHuPmR1ckSrvFJqm0Dw6Mj5YZC40ckd6OtXijGHlxm5+
O0EKbfJ3ZhE9ccCpIU9H+jZSWNhHqOAIGBhLOzsbIHi76SfJclufm7Ep8kJJlzWJ
9tYIUs19gQF1N/UK9sYhzzK4lGeWkkBGVDa4QVb+W+l09vWp8/0EultszNr96ax9
PnfYz31Tfx+Z6j/tCjol+KVLD7j4nBsuV9S0eJPHeTzJKXiIf85zaJj1ZE+Zgz+D
TmlqUBcGcHtY327wCToRLoPOlC7yQ44u5RzAVD8pXCXcT3Yai+cOjiheohgwjFWW
ghtQRqBVZn7O14yYr5jztgthKQzuEEky6e9/05+0mRR8LlBhk+paGcflTBvBQGoF
EdwOCggMhMg/coj+RnbNxXa+DZGeL41rg9OmmTpjy58pvOknEKcRTpT0FYsVBL/O
Z2CCvGc2V6SzAsYeRil3P3MkITCtomIkVxW6YgPaGc/Nc4lYhH+nMaZXvLiz+3iw
ReBygv7Vk2h+ffXUtbg8u8TnYK7I0GCKGUX/QOBC2Pq11cm3ma/ZZ9PrgdF2CzBM
ZmPkx3VGwOhxa7PSsbx3Ipl9Uk3ICOFecBFWrbRI8SJ1ZSogqdZdCn3zXTQRk8Fa
mRVVy8GjSxo02RgUpSu16Cwq3I1/lgIgp+K6p/OPm2P+BjcfLPM0wDDrhS4ZjkC+
1c58VIsXCuTpDXwRzL0vzicWswtpX5035slO+GK5keGUs5l23NPso3g0hoQ1ksUV
gyGhhdUDLXGksxvUNAdYk/JgUdRYM0FDYmVbnHlX1uaAANA9QGW9kFWtfhSdXGbk
Xdjre/GCwgdTkjjVaaZ5+U2YzotnTTCp+Wro3J2KH56/Bicho70fTBr5r2W4U6Md
70Cbb8mSFheruARUzQRnTmK7rxhvPUNBNrFKRicT6N7O+wazPcLVpKV16Hswavj/
V8sGssbk+dyPH/S9EZNf/3VXKKQEwGq8BnHSD3IAUhwHt6U0nvgcAgEO8QKj8Qna
6r2ooLoEIja3PA8Hk3PFDeWuHkqzPbWnZrXoGp12vP0xD3WsKOlG0Yt1rZRfbeN1
XuVffwTRb4a3ClPPecBBQWMmw3hWcxW1AS+5rJRpu83m4Y50DDnchHeI0pd3Hxb2
u93xmlNIquaKEYktm6k7xNtClw+Evon+6yDAPMrDhgjpnUZHaJIfiCIKsttKoWTB
Y2On39xowzCxd62KmEnifJstb4wT3q9TsIwF+wZjCAxOQeUC7ZKfTYv5ZAwHqssj
HSsLrcZ8fmYxb4DL4pgRIPmZncD5hkQMqJcQtA3/zLjot9ivhFBCoJvRecHAyBPO
MmAseFzrORivMQggjLW+dB8aWPh3k581y7BO/Bu6HQHQCF5C2u5y9shDIMUCqwiM
8RsPGv17IcWYEW56WYgsFdGtqKBd3FrYj35egixySn711Lm+268BM+NFpF7NqUDO
kiEgBQElZ8nPgPH432BbVvL4E57/nktrPGAXLimtBkEZxyZE3TxZgECK6m5uteC0
7xD98UH/SEnCPrFUkc0IR0tZ4ozoD4VhGKZEloMPLtx+ezLcLC7Uuw8VmEgGfgyn
vnY0zde4ZUqGGnEmAVWWoHz7oaQcsaRv94BAgzA4zi2Xwx5EA7bC9GLut8S2HnxE
t8H4/GtIlyy49YqY7OFllLqHMojSiZSELdB11HfcvnXBneE4LaIGetV2uF6Q12Yp
gVbNY+sh/tHsrWT+SafZPTxyMBd+LL9sR/YzQ9M5FmqhspAswGeaFSjJPzpfXMAc
ThEmSSqXuci9y0o4QRRdd3XIsRg0SJlDR5mRylOF9Ksb2OpnNLsHwxzBkNIDj1tc
AKnQZ4elPPAAHJShHal8yYKE0mid9IE+HaQ0E39XxI2VtExKcy4emJnry5b37/r8
/Oa7IRnIayZJpoauBFOvBORn7CmTwAvJTc0+KhPC99uZ4SdxHIfcjBlUkmOOfeJ/
ZAoCwG1et9C1/C4fiKrAiOzaX2ftLpUjL3+jTuPddBv9pgyN5wupysQC9hmHT42t
MGrlNlZUKM6Ayp6bE8GguklbPpo5LxdX6WWkeQ6JNt5df+BIRscQB4C+vrewjCGW
jvJ+pCXtKQC6Pqgi6dxHOsyCaJtXdVTboAq2PebCr0tgw6GbyEVf/q4EOIBBIV8q
2HNfwOhH3UllEivZMeiHirtCns9VbiNhSpg3/SukLr/tHbjbomRKj1tq4TC43Vuy
yQa0XuHlTH9thslWSppsqAac4tIT3bF60K3HLWKhUVYDv0MdTPB5RjDYrFKgfUY6
edO2RtA95jh0dlv++njXfjLoqUW40GJOkMfx+vqgBtgBoc7PycRC3Gv59hsUwqPq
ihQSHGxbrMFssDoSCQX+gmaH3vGF4DxDh1zs873AWDyMKrmaC8CDd8AFDDrfiytI
lEyZylPtEYHwK+HuMngE+L7QxBX/9QkovIuYjDuLE9lKFXYm6n9UrGhD1yecLZ6i
tVfnXcbwjqzl/rHABRN5ZS1gDaJutMd3bvz0/ZfRwr42LmYRuxFUr8AjMjMgYuIN
x6wQmHADsc9gMV3mbTSVqz6pT17eDrcd71QdhvpZsrqoLv6e3q9UYZm3BD0K76/q
/MsjElFSXHP0VTf590FxrIfXwk+mPIcbC3LzjHoMiOkS/zxXE6xqgBSnXX0iSN9O
mvQzFO8OWn9zUU1FBl0HjYY5T6AlVWdD+Jrti0r5xdroOk7vAYMGdl/r0a0m04bq
/RArOXaYKPU9SGos20CWBM8jbeSt3eSf2GoMOUabGD1xtk48QjCoVx7AeiECeBmX
zelfc3Q2GLbsb2LsGPcoh68NMFHulTI5N8IXN+giJHEz0QJey2bnt67Kob034DI1
Y3+bKaBudCvMS+Af2C90d8O1VUs1npA3jMA0F86jQ+GdXRn09QSoOOkUp9MTIhd9
boJKC/iGRXO6CF0GUSoK5034MT4MAnmj7Inmkrw7eDBf+B5ZidbaxEuKtE50TbGM
tibGlszY/ebz5K5ghgdDHn1ybGHOYYmoE089cBxetGT81zsCReMRDZ4mfjqJ/OQ1
QAPGYNF2ZJ20/CoPQsF8LY6cVoZujAWtMgAc9ScmtmTAUTIo1dyhsYHe1qMHN+WV
hiLUoGwrgNgIgdABKiu0El4bQDOxljaXNS/rSwD+OWSQSz5tAjgcfTV5h68oPTEv
3VhdoBLcLmOZ0jVKVwqd9VOTXAy73DvzYoFPD2dhxGSX7dyZwx/JPPLE2Uyrn972
xXnX7k6uqpgokuaE1fgqQHbxhKOfcGnlkVU3u2QLSeKOw4wdGI/CuSohz8b+DVmz
cmbik2AbQ0LdyHtdo7r5Ec4IQAAVTmL65xwcjm3OUTiPindoad2MAfRDsBfzk8CG
wqkFBw2sfaBaq5wXzEiUnQp5VXKGDY6yuYq56WwlaCpgXFxlH7gOt/bIDiilTbkf
gLeCacISzcfFQfCWgPP0ucNJKKa7FYCySp8cHrlXkW/jISqniC3XWT+kII844BIS
JRknzSX0nMkHdx1qo7H84i35KTfrfVrJKNMHs4uQSpF2hRK/ng1O1aHiR6EbzbQo
w0YHI8B2xDxfuUNNocCvIbJeKG19edrby+Csf8hI1J7fCUio9gsDs642wiy1q6dN
jC5oGkxcTKNH2nDK2RqPGLTI7HIWPdTxBDqAcZ0iMk+yh8qE7/RmXlN89ce8RV/e
JFM2e3SwFGPLsuJzYicF8HiYXnRqswLbMYiUny45yFRUgZzUCZj6ZX1O+BfCiHJq
utCCJiClC/eAqMCJcQoLv+sMAqZLIqSeScBvQlw1aSt4eBVW3vTDHI8bHypBryc/
p6tHmhSsJr0qLklFFanUCfaxGMnQwag73GPw3xjUfX66W2OqCd4Otu74yRR19KWc
ddiKonA15fnRj/RyC3WAfIPSJc8w6vHhHYMoTFX3N6v2c5QwfZMClFqqmmEdASk+
YE1S1bclZaevg6ZuMFTsSDoygHwa4ZMTvnPmQHd+Bj0bPfrQlbl1GvGrPW8D4f+k
BLR/TUI2988hWlOH9pHGtUZ/Z3VNf0rsQ6O36eYWFXzCLDFYUnE/p2wfJ+tRfui4
pyCyUcpv5DHMBRkcIUeEfmTTSeceoRjquQANy9IDA1Jky/u5QFtFlRBal0/NEhVg
djHELGPocFAtijOTgilTbp6gy5ZJefB402ORVOcmWANAmJ0C76v5QopcC17xlGYF
quAX0XjMB/VKpivM2op/LY0gPcIG3Nw9WN+9UaxaBURo3BSZKirSYFe0vhK2Ek8H
givhfv02KJWAcesWfUPqeSQwcVhQpVMl+UA2FP1DIGqLF+dcXfPDlJKgUl5iHDS2
s/cFjn/fP6NPF5Bixg1lkuGOgimT/x0WYjB/9OFsSQ1zGFBoVRfIiCwj0GOOqNyr
UxIEd5e5mYOT0KN5aUFekukr7qMPRK6012UHcu0cw3Er7CknLIv+3lrRLviMz3bY
hEbGDJAnYMbETZJzlkLAZHjqfGac2Jdh8hLCle0OIgdTLDPAN5GDux1kYhVODMfV
dlGtaIoMUYgipknpC9zehBvjbKrL8swauFFgjzZCLWbNuv2PkvkOVdus6tThZ1kv
VJnoWqcBfkxebHtW9tmXgJBXOzc/RIzKzUwI+8lDAR9VCEdQiYpomE+hgF9Qomk4
gcpOJqWPngmFXcVNUF6By5L1oPQNdgkyDdR6TBFBGYcs+ZB9XxdekgqnX4SyIBFS
vvt8eGPccqMgIJmSfbx+p1CeGcvNVWdWmC5eb8ldSFs/vYE3Jz8WUISOYmUz3kHR
7NlFci4IEsiYSrzENI9TbdSW3foLpNGInMYd4k9W++tiKNP3UmpSOWMxftebA0XH
v6RCZhZarcNTvk8T244znp5E60+chQoqWPXSBq8zPyELBISIxlRahPSBy5oUOgik
Op1XTqULi/vPmjApRpBrkY93vTTPh1iBoksiBYGdir9wMcImHqa28L9VFWyGuzac
i6AITp7H77p7+HlNEfY3k22vKNd0tonJR228iKbzl/FXTl2InfZatvKTYiORfZHZ
LVykAPSvKSuaEBah90rhWgEQI689beAg2GA/n1dP6NHUwcId6GRo9vcocJSRjxu9
HU1Ck6k9cARO3n1uAnVEyAUayKQHGD7l/wdHfc6WUoqNlV7XuP369w5m0iOhigU2
kHq/jMRWLVP5xYDPQkgCjuoDnROq3gpcYFyKGwM8XCawPNyFadNpFIhuoPZClCke
WwfKKT9a4+SBFqUrpakhyRQO1adEAauVPCcLjzjAQCa2Ed/Snk8H+GxqLoemxRYg
LPs9mVamSEVMW09/kNPlYub7pthtxUqX2pw0rPWeNPCthS+0Cp5pQk6EV4yeB9Yg
iPmaMA89gJP0E/clvSlgsHWRt8MCUP3TBGd+vlFr6fP/IxnaN6bpRY9WE0rvd22n
40DDvGtTNnUj7B36c3U6wk0HNLoBvLve+0m1bgwl9Jle+cqmZw8y6iLJY9hnkwt0
iGFpCVpGzBpSsNdgz787pr0hpdkQQ95Ftjfg8hMV6YqCtBOWZXwKl2CWNt59CeRL
lLxUw3Q7ESHzdYbVBUoGThh/O1e7GgtvIsLJiSfLVvApBaIs+gt54u2oYjv7oHoB
Pu7ENve+w4JMyI+8dl72CLh/1YaQ7pqvLX/WhJdYa/PP2V/R0L+wwzuOpllsScb2
EHn6kcEVB3+Fu1EHWVGvU4pCwI3kbGnVEMP1xir52nvrqkC73yxTdqN6pUxU76x+
K5JsK8edTrMI+FOpSOlV2AxvQUh+ckOIiPtbGfPaDPxAkrpDWeJFgYmnQJR5+d6S
ACy5YpzRz4AcaTPtHzrmvAIr9/tTuk9nnIxFcxxm6tAwWeWeBNw3DazoTFLzVlN8
BkNMRMI2mJaAT760WtOXewDXElpBrpCzlQqAupJHYK77WdhZvQMQmGUlVQq531dC
9V8rOmAKVF1YtWAA9PtGzBGhjJK7pIAKNpM2f9boPK1C+E9443vTtCFTarzOtrqT
PEEAKG/IDfyVB25n6aLz4hpCc3EAv2Tp9BVLCTsosDceu9kf0TItxSho1zGVUJYA
iZbdMp5FZlL/cTULuhtyt3oBVtJwlBY64oovIT6hyJ4Q+t67Pf6XDAXuxciMQ0WM
bGia1PIYQcD3oWGYMxPxxlVvj3C8c9yfxEDusw/EGUKOAVtUughPQYmnGHILQ2bA
ytE3uguZPLXdESz3UmZdfY19k2PiWY3ZbhA4EQxN3iSEQnjdYimQm96mOT16ZAYS
oFG7vCj0MQHm558HnsKzwopQW7c3FARGSJACMWQb7DH+qqAJHq8f2vhcqXXcW6oS
ba6aVk6Y37S9I0F9HAKu1mJJb472nx4trk6agSaSDSIyHoVfCFAov1MmZy+7a3zw
un6OwHXFdaWWxk30E9yhF7e0vXedwpwC20knB3/Rfn6/XTdl5v3NpXwaxKsI/OnU
6sCVnFts6E5/FGqQBtRv7wSKNy067sMCg4L8a7D8B/J64ld/vSlIO+UT1Vn+o8Zw
E7lSh8gi+yqu1+v2iJW/QplB0KWAGk1kAnX2cpHc3/PgMhBTroihTPfWrKVWkI9R
lCl+fladqA4i8C9smSISzQe8PyaUEeomQDizsEKqSMD/M22xbA96vd0oK3gMykrZ
uH0Fd8KD0tScQinQKmpeiwF3qfIaGNBHbrCjbBvpiJsEvSCl7/lfr9d3+/ufjFRy
CW9JBO56g3sn8xay4yQN7/SJIZbRCtKzMHYLsWLHtfM0smbjDlWm8avEnsoi/Cfs
hhfaGWt1tQYHNt6DFGXpTwBogWc5U8u+HWTduwF3kKv7o6jv2RQ34UTqaX/f9pQc
Dkcdhb0/rOwCxliOIjFaxQ7YWiJ2zsf1NC9nJYfiHfgEv1xNUM4hh3ZEvVp7Tdmw
IQoiWVDmXy3JD/6u1LEEaMig6+r7HKtJOrm9hbZJ/vDHSf/Xt1riTGEl6zXhUOyW
VoVEfJXmTaofwLMhUXma++DOgXcy37utOmVQk+d61T0rpg3M8AShmZCXvQzKfzUE
WqbjVbBbBbVuJQyw7qAuITWTndTTzffs1rqpFK5I6EdNoIX4unM27tVj8lzhdPKA
OE9A4bcnKaD76r1niFtRIxjyD9+5+I1CR3k8AuMlAc0Jq4OGzyqjvFqgJOWFnVYh
LMzqtOk0kUnEihj9B68g7JXBuYOv9QrftlYP+HkUqH9ActYsF9yZK/vqNAsSoHmV
P7XaRW9iZJ2I6Rtm+LM4zBUFGN8Bue1DNPscDgV7asrz0X7F3vTg1kcCJ8Me1TFd
KYqT1Gy2Glu7WiZvNODs0uxggdui8ChaNzUiX7FTwJY6P1t82xscpN7F54bnvyqu
dIfIEKBPkQsukv8g+OViN7kn9Y2POgfmJBkmlQtfJba49R7b5RuqQYa9BSGwum8i
rN2R7BmKbF/kSW43pIjjfpygUZGF21bDAsJrgVKtS/+HVS74v9k1iKNtf2BQYo6e
CsS0grc44maf9J9lUlElUtJUc0afqHYZE3uyst5rMu3Gtll96/HHFzbQf0IM2txO
XvaRdpqBqtB+tdaPYS9nvSyLcf6alOJxDrpv95Lrqos0BL1XD4q8vhNc1rtOCmEG
3cystF3/9cqHgsRmVhVV0EyZMOkahqiqS7YqD1L58Q6Qhf5V3QuA68VpazKzl/6Q
ummI8Pr0r8ksLHUIoEj4hE4MtZEzIK7AvRM0pZjevVU/zklXPzuFRKaimWZgqdBR
s/rcKh3aShNMZC1EVmGnc+bMh82b/6PwkvqxfyoBjYpIdATtDZAT/RJRS1Zm2JoP
/NoJZu3rfLC/riEAifw/HjaQORJ09+5S2ZOVJH3dWB4m9cCHWWNEBGgM8MczzaGM
sHF2S4flaN+GmzY9XtMWITAysH9RPCSS6efrz5zfs2BTG+0hTBr49xhSh0zUsvxQ
qFBP469VEDyVnlv8PP3PUel1pWw/rtDIXDXj4GEIwykG8dqdt0dW2KGvMVFAzAs+
x7djLCL0rlDvSag5Jc+zgXiMFDQAVezeTNlZl1OYbf/Tf6y0RmuvrITf+U/02ouC
qZXL2Emq9QxCNAJm63slAVbO3hi8AGQK8+f/gOV4mywkgXDnqjRr4U7fQLL24szI
eDBVKguufm5hmTLTz743p9JEJBjJEezAutilQ85n+EwhmTxF+8ETgYA54vCJeky7
S8yYMKxcB+w2dwtlxzszG3DXvT7go4gzNezmavBUw1zl4rc6Ks5Flh2tSmGG1h9R
iyH3/6s33rmaKm6X2em+kyUxc/fYFikTJFyqjYwL6nSzXFsrbX6Fs68aqKlUUAmU
9hCeX3sxcNqAIN42k7jlvgXwvF198oCJZJuZUyjThmRyXXjwyqYcfyMuJXJJu4tX
73uClUBmJhsTe78WO1Nosk8lmsK1cOX+3IgTA7xd9nKrcJC+vsCFxmqKPJqZhx95
YspZKRElaZi3KVnR3x2mPFFouZ9A58uDWMS62QjHDOcdx26TrKddVeDd6sLoxqkK
UedUwmwQBeuwXrVB0h+ab8zxqI0HSPwYi07V11uxHM13y8hg7mU58nh6AMYBYoQU
DhUztwmiEhe+fOHIoxc5dIs19gT298PAx5Hqn0CUTY8xIlTddvXDbn6jQyILM4FC
WGAtWaMgvje/QOZfDvMdeT1NDP88gMBWGNbPhYscY6Gnao6SMOW5YSfjVERdPvnM
r5EzuZI7kPOjKIcnnBsDlkJbrUBDaNINQMdCCqLFxrMbrWh41xytuWLnPuCCvprA
q0QnS7jVtcRQWRQfSJllTZSvGO1LAgOxIdFF1BqONj3Z20L8rRjIHaJgxdWemOtw
y2Lp5vqBHIVJK2qtH1gLrIOYPs0YDopbKZRIKuDZfesOBYqjrdUVbHk70f2s3/35
Ljv67bMs0qpN0VhHgu8kbqTOZvvDnMq5Kf2WNYmyfDfq/Y9iOXUo70DmecCl4O48
sC7gxKx3wv/XkXnpgxn3eLUsJAAiN+PDOzTZMqP3q8JbQAA4pfKoAVhp9hgQqgrs
0Qd4OoXf3u1oy3oPZWryGJASlJ/CWbaGdNWUrHSbcpiO7GAEcMlYF5OOSVzBV8U8
/2M8VaJpX7qnlCGu78Q9wkT5XiUiv3vK+pjgOyyi3K3hxgRJnAn5kChbQp//X4Br
nfZG42k/gMq5b/ZoS+fmam6+bof4pCSpsSIWVxxrNIlKoDlw9LQaCbIuA+VYQb0E
L4h8LOoEu3ERZcO2COCZIHsqMw5Arz6Kw+GDY4jF1Izz3cAnS4zt7cNrSwkrsF/l
/t9AUA3Dd6x5VvJzTcgvjwN4hFosudE5mZa9xRfgvjCK6paoPnqtGcZAoSenkh9O
27g86XX2SFxYcYOQuaPhAtDdAQMJzJ3m0D/iSEYZjQ/XIrBI8jClgytjpYaiGPtc
OAoWT5ODmBYXUgStEMANZWM6hIBljETeRrOcs9jb+C8ObCPTdIPdu62Gkge6LB8f
fNuG5p+CikgS/6TdHFc4O4Ku/G3A5rAtZbcH6bRbZTM89SeLEmALgqFWED5EKpmp
78DiGUvYnaexkgd830qVpo5Om8kqoPmRzpk5BlEpovu6ytxn6moDp4vgSNnUibae
OEyeYhp4UNIry/PIPnR7xhLQs48StIFA+A2KqfkwbVdtFVGsHE6EPhjJsjK6RTjD
RPmaFtbQwZBz6rTmjMWcr1qE1t4awi/lWA6dWJMu5OG4oHW5laHLLrgRoSxd4KVq
Meo1aKJ4f45GBXcshfuR9YbQvtQm1rOiGrBi6KFS0oDqLNOb+a1KcAOHhYbXcITM
VXiH5XdkCnGB2r3RxJ1ZqAgZGxv/TCK9gnp4bqxnTFovchUXwEYXZ6LmGXIJLzEQ
wZzqwdTcswEg2mM99vr0dRGV3RZnNRiWN2ZQFr0CyS4/5P4fGH35U5lhhqGLlgNC
WJDo1vLhW7wsO/QhazDCaRflyycZgZKA+Q+Fdp+WNAOle1t/0k2mjUzpxBfWsaGK
RyLhNEyA5k1iT7Ni6pwbY7c6laZThOyvLJdWgJl/NJSD2NpK6LWUiSjj1fsvmgq3
vIts0uq4dvkFi97NJUhvDLCRe09NDghTaah+1CZMebCe5xC2tf97rB+xGtHzs90E
P8wUVfB/+4vK4pa9BkwY8MKJxMdyQAul5lt7qLKvWDJ7OzoLr5s69ICusKixnW0N
fAGjL39NPOMfLmyUZxIMTO+eSD2hFLBCyer8hQkZpyjIdvk3WThXE9yAhpUj1zw4
yl6dMMVscHc/RGTtgX560B9xkWVPF0O9Aeue5j6xo/59p7UQ9f6Z6IY1eB3SGi9I
ImGe5w7r+HfR85D7PDLH365433CM4+jiAAkMc10eLCHgqMxlwKjxKs3xZ7SRG8hb
p2qvPXMhntF8IL+2+ef+rK13nc6rQ5ZDHDtdUMu2ESSurnCHpD9rA8ilNXtbncOM
xb5lebDXbLkekYBi3+0sjb1gARtgKQsYAZEqtAxXwAQu8JdQOte2jwCPDTgJ+rUe
KVerSQWnEEM0CaoQCDWPEfTS4gXOv0bzT4DZsNTZFhQqy4NRh2vgxSQvqu3Y+/PE
jAhZATvt4Pi2BMsMLpeMNm+8710ufSLtVcgdet6zbmXuwRaqfnfSzXSncUBxjYJV
d9VDpW+/MtDmOesQQXAx2bV2olvDo+CSejVxRVSRlmHJGgK+6upsI0kzdn675eif
0Lv0bEYZaYEuF9ozllad5qtmK+uApuu18dK25ih7ZRNCDbUNG8NgGtlq2iqrMmCJ
QH0FPXz4hXoUhIhwoKmfWkTmVXf6/5K2W/KdVk0Ugvnu2uXcSO3CDTcq2vkgCQRs
QJCvSsXTFf5Am6pH1DhsQ0ykUyeo/qFKKLVemikIYuqmua/3QG9nb7Qlx+ryKjyN
EjEPXqR5+ZppY9wc4lGElkIsl0nuNjykaxTMRv6bgpNoXYckC4uTHi1Sh5mgR8ao
jd36ci/6DeWohRjQFGOX/CP3nIKkpKv9dhuVrNMTEnItlVyc5nOGMUoMUGLvpmCi
/JFAgqUj91L5/uxg6Gz5sMkt4NUnjRYLxlldpHLZG5Ugp5tiE4z0x3CYZfsZQg0k
i/0S3sAnDwzsAnhiwAl5OUJpuBm60UfBu85YaE1ctS9mO6NQIFh0v0FpOJgLXhTO
v/PnQB7sqYbdnLJh492sI6evTGRPRdt+9WRq+J8PlxkpimHW3mhJSfcPoHBIf3Pb
wivWxj87o6m8u8eSvP4x1J1IB9IeWhqgTMFJ7VAA6OHs+B67PdDI0YYVkylOUxAs
uEkk/sjLaW8h/7n+T0Y8sz++3lHE+xPZAzAz+Q+psiECcMwNKTNCSldGXiNMEP+/
ME+04hORGqs9q2PnEYzNmrr42ShxQMraIkYP1QtMC37o9lx72aeeEOg0e6RzE7nU
Pz6JSdAOn0jkGPmfmSJlszHJleMNE0uPCMm5Wg6GKxU3PExPrOddihqmVgbnPxnQ
d34b9rynXRdvOeZPF6u2bIZV5Ms8BPbMMB9aRcYiDfU43TSn8svOj4FPG/ihwcdg
pCz2CApKmfEj9vpOD5qhEdfUdOUgtWEePViou4l26zd0T9q9PB264yKoxhrEg+2p
zbcw7gUpAggGYGwt9+u7fCD218bCAFV9NaDRjjb0SabmLUfeYKmfqCdf0QMgFXCH
/zgAZTTzODkdpQ/VPuxuKA6D+Enq80QGqmjyFMsItclkfJN2KTZAo37njdm//JAb
3v38r1sv6KDmbRHqJzHGTnS8pQi8EG3pHpL+SWW/LfGHrSYz0dkQLoYb6Zq6HVsj
jZJYGPlzYHLRLCLq8CKjfKkk/QDr6eLJ1zOXPY2pi94/jbrnCEO9IaNcigKEyC2n
BrEzHxtnUJn1WOIm/ALs+1n1nAKzJeMTjk/g28SKFrrd+08FUp1J/vJwlKurEFDb
izrr3b9y4yEDdHfmtX23RKQfU9OX+BeEwXr/CZoXyFcOX/z6ozbM0CzKF0zqP65x
+UMV/0GuNgV5I/Rycycpmt2F2Rs3DqgugGclFEapS/usgIEW3bvnzCjLWD9YYUdZ
hK0ESP0OjgbD04qsZitqryQECsJMfFtvCB8aWnPC7K8TWSHKFvs8gmUaZyYkfGsv
rnSRMtAV9NhX4UWYNCTPetsbdX52V/CxgaQrlUs33k64NgJZqHLMFf5JK01Lo4yZ
sDBDD6KO/fpoUdjbbdsakQ/JWHeLLc5wiQd/A3nRFAE6RleAjBMGBd+SnUOZd9Yp
YEj+0ThESuBPDgbwWMsGh+XKDxOiJMGc6VJ1IYDnErd0dfVIFhJUL5nmyY0t7Zex
Ili8NM0+buz5HxEBzdxSrmWsST/n8oH9zFfDdNZPHJs1wXZVZKAlTQDKss1O6h4j
mUHxdXiHVGvP/ys/tNti+/9x4zuKuLt58N03z3RinpkDdCmMoiOnpYxOan8YTS8/
eiUrL75T/glcqWzOCDcjq/RZGTqxQ9Ff8cKdt/5FpatkBD+qE0Nd10PKK5tcxBRv
8cY6+tUcGKjP999C6amA+lopzmYQH6ohv7LtC75UsjDEnSSb9Yjq3Ad5mktbxsC1
OcwkotEOsfJ92sz6zvw/vTO8ET9ytwJRW/UnDi3Kr2mE0gBVnDwU6D7eDBqDvhQ3
IgXpoVafr4B5VAlsjejvv/i/eM6gqAxhXfrK5LFCHxbm6anHgdrkHcpbvdEeIw5+
UK/jW7Mh+h3Ttbo51W5VTmkZGqzW7rjmkabDTqOdNYiOGk5NEXa7gSGz+mZkNrBx
JqQuloDcDqrTzWTYQre6o7UH2aIwI0xPv+RNk9dHeejICBJsVM4TJpPNUZsNADJP
G6lqGuP6gZm+/MkuoAR79LVfHTr0pCM5Bd3sLWRrwRnZ6BW/cSP/Eqpf1NQM2aK4
rmvQ5Y3bHMInALc7Al6FJfe0YoRw3IXZ3HkMfGSymhvKxXOqBNTBDsf72i7Fp7+v
6fQJfmhW0G6vSB+RbiiZMZo5eXtePXIlm+V8V/bP1t6/dIu4NuUDYaskYAkqC6Zx
vDfKCAnFDPa2GSxztFHRX4unl6i7nAEsv8nj7KauT6Eom2fC2BOV9IEdNY79s5pQ
ph+DnnZ/sY+LXtKcRntReR7LaFCe6kieMO7WBMWv1XSRYSJxxbjoMC/u0vZ8xnYw
rnzr+m32jFtfZCrhQ4NNpfZ7u72GGX0tKd5XypvfLf68S2/Tkd/tl30TPJWh0hF2
Eeqlz3oUVI2NC55O+NoMg/zZzlrjsm9kZzbgBxdonuW7wt9bIxlKA2NVHGVZ3j1V
c615Un+SEHNiakIrsCha/ju/FCXRNpfM8acSmwniMfZV3nxUmnYI2DCoK/UikAy1
IZjyaAlFjjnCFR/OIke1zP7ZrgtMrWXU5vASywZgNAiGakW5pTvKklFVQS6SE+Bl
3FR2N0wx9C1K2bbHnrliA5vln2Xuia4klpuK30mRnRWD+0LuqHu0Fdwh01/Fg/to
ttplFQ33iKhyJ1tZTzhJC56VSnWIhOj1OaxsSIHTSfFvEInODKRtfVsjrHrirAgp
fV7plwqaPLAqXkhrcRm6M0USiqbfHzF7F46KMGWRd76LlNru8gfIOc0yTB71dcAd
6pFK05Tmb6mnFkSOtf52bnEzf0zS4xUkRuUbSH5SLs+TnVeMS2P7lejD4ev9Pw8/
gi8J/XCDABEXGoxMqEj4zfbjVFLk1/HHCgXUpu+UvDT0UWjzrLPOralghg+sVArs
NznE7Zs23vNMEAuoywtptutK8lbnl23i2Rtyyrv6DBIDBrqB/ieaOX4JtJ9Uqcz5
j59LKw/nSoEHeO5jQSNowF4ZdVwHEnK4Q2dpoGdnFiWwQYKWDglZRuQ3ycc6Au9I
YscwFKDwtwIjRFOlk0PU12V/JTUKEu9qDBXzKms56pvuCmB1q3zFd7fwEqi/alfY
SxGR0jWg01TXsQt0yH2Xcg8WblazySX0YVcDVtfvqybD5MPozOLrgGcUY8Nkv4Ma
xN5PapndL8KbdkD060H0qaU6/zVlQFk3HyzyUJhPWihYFtrSpd+xEWCQ7kGkPm1G
FFkqqyTAdSFbCFcEptYjnWEJW8b3VFhjXyMq/5iEA5W8BJiRAA53MIM4vraHp8FB
Khu9KRN9Zy6F2Rt5Zf7vk5eGU2vJ1SFgFwRjQq1nvE3diTpDq4djwHWa8rLf0Yfg
kpJXGuuqKg4J1xo2SnesAM/XmypUQOqurqMkD0rbk+A6YXUz58ODbyn67VJJpRKW
LnBd8y1TswE3phshLvKpWbQa/bHVc8kFv6+AN2kxGjRJ3KceJQQH11ui69iWAF0u
iaXNMJiSMUMTN4/Pr2LwNDyIYsZ+pHnQRAPjjvebuWhALbqJuu4eXZL8FVCbVJWF
TFOCUCAP8Dn4m5y1W7PkVCLplwmiHHlskT8gw600gh01GcZUXmJE9OoedJx4XCpP
9NgTVoaj0bkBvPrgDwRVpHYTAUESfdz0/in7xPWQ4HpDDlygISIp8vZVu97wj5sM
gzqYSmOAhjKgos+NGJLH4CuTtQB8Z2fyIBkOF2uTCvApBEQKoRmAemWvWRZ2R2qf
LxM3aWnm5DI58QvogStTBC+mU/IbTecHuhI8MiLWUz+mwQygfdDtbIbAXdVl4NfL
MV234YueQncTnjIQ+nc5PsFeukZ6ND84sKxgb1Cc/2Aa7RKreqyqRYMpTKxO34jg
JipheCzom9h8o4pNTy3HZ5z8TCcLWj4huTOr/O2tY8CXKGySb1ggt1oT9VH/bl0f
LodZqh+cAhP180K3fOBZds6N0YmbmiFVHAXLrC1qrVG5ae0g8R/zftq4BiSjk9Jv
q6iAAGQWQrf10XjllojidGWPAL7c9+iJcemSGIyadZ7cPFf8KxG1JHc2ndA5UnDV
mGefBVlUDE9IRA9eEB+gt1LQ229bkbT7wBC5CrwqJtfK0xuLhImHaivkNuic2Gl5
MkUXnsDp62+fKfnHxjoiHGscsAQfDCuCMgYcBityGc0fgVt+gMWQriGp0dPiMfUD
ofF4RLy5uFUSm3Wz/y3U8A4jhGr2PF4TQWBIrcKltMToZRtliGsQZ4SEfyBf+f+P
Ra2I9k7P+LgWWuVnvdi9+zabaYR92elG1XFvV4MsCoanH36NOAVmFYCRSyhA1Law
XUIeO7esAN2GGdYtGRrGyU8IaVUNqPjbM5POzqLOMBr5fN7DXawGwTQ67PeP1p8U
wSjKxSGkjScabK3Mzvg+VAWZ+lmz3ju3FK8h1JYdSVj0KMeMcCY/QL25rQqWXoW5
1c+V2SIraSN/Y2cQ2QIp+JdFtis0NBDuufcvs2Fkzj5TSxWYr1jjFz6z6IqKj/jC
9Uc5UimIEw5qgXpIKl4YTu5If+y1dI1mQ2pwzp7i/8KAzgcv9Gg/Cf//FzjMJI+z
ysY0Z39Y2oryaXlIMkuOwqTxspKEH8yu0FIyEgK3sSGnmJvX9VfXYFYYe4yn6ZSq
P2Iq+CWuyRx69iAlPPpplJdhyzyMTYXFBtX5xyf+FlgS0d6m86vLGvYJi0XmksQj
IIWhmDsou+dufzMc7DToViHg4GgzS5X1xlRYTN3FtD2BhdRp7zTDL4jv+RybRB4p
qFh5vX8uB76c1gBTJM9RTnKPxEUHEuyth3vM7cAUCpF/kweyXt6jBX9bR0GtVUEm
GLUTFdxOSC2NODIZli3nh7jp8fXb5mdF3jjmLa17RHIx0fKz9KaRJvtwrudUGPtX
zhh4XmbhIf30aCrDfTtRWxzZaOd9OJGslTlxEbUVgM8+WszbVopneADl66qBrNE2
Fb+NPipCeTVcEs/tJ+vg2yzFa2sJF1LRr5Zoho+YyDTbjH9puiMyklXU4LGZrdGF
kp1V7tZVEjQ9DO+cyGN6ns/CmrHtvDZ+FEcd3eeT6C36CkvCRk7lMGbN+AxTByU+
bq3yDSaILD0IMf1QQk4nTgnYbNUnuTv6MKuzLr6Hns9UnAZGeyi/FiBmaXXPN7FR
mRZVwlrT55hVIzvILcxG4/EDzpQ41YO+QBJ1srGJnZZZrnmYSMzKTkvu560SSwx6
KgbtOQ8iwxx/vfKESv2QEiRPuMMhgcD6fGIOBjfgxwYGToOL2wmNlaJYesAYrUVF
dFKt5Patgup6MMZ/KM5Hx+U06JC8O3gUymXQKlN9hf7nX30IvKTsNv5y75Cw4Sk7
2LVishhUcXJlssbHev/gNjOf/dSbI2V3fb4g+uMQ4niSkoIR9OVMI8SjWMSYuwU8
1daXvNknAPlwkGYJhmRhkvbYx3TQFEXIJOXV4uRQ5nc21JQ0qgbkxJXc5lwT93F4
JWj+DmNQ9GRnXR9gDSPsXJ+1+qwrI0EHuTTXN4zYzqbcLlNE3HMNmOyIyqIdwhCq
MODhwPs2vSCrcWZIb2ZRxxnf0eZiV7Aw4Rbhg8l/yPQu8zyBn/tI5OwwqwMVf5J7
xZgNML3EAzTOiEPGkrPTAWguZUWtzbb2cO5VSVQ++uDA9zIOU1joPymyBbZDex0f
VmdePxWRHdtq/m0NwoJigq+Otu/ml+1lmi4gKu6NPR8cznM14/0FEL8DQ/ZvV/Bg
je5u9HWC/50YQUpyxFwx0ENDPsLKtkyQQZXHkqFotA+geiMT6LuVTI3Jq5vF+pSa
j5mgJ6q45F80vJWHQpXXzbwBA7yJi+lqnZCNAfOP4HJOef3dc4wOJaqlOsFzh5BC
CGgwatX/DdQIBMu/KZtn37NWI6H6QsX1b+wFwzTap04fm6Q8hJhK6WjF3APteTnz
ybfQsuhn2l2YI2SA2MEltq24NqPxrtyJQWfdrYll9q0clXwIor+rggrZHL0hRKjx
bQhs5ivLI1v7cgBO/dGaHsnnLva5qNjPsVJ6YMTkc+uzLRd3XJfpUCVhjHVGzIuF
unDc+lz094XnleyCoD4RVAOOxrPnanEfnl3wbzwiQuwW3moYjC15rJ9pwH5e/JQH
URylL3zCpUvMIiWK/oVFPvjtxs4Qqfv2DqOdMeZ8/4Egs1FKDCkeE9HmPbTfscqv
RB4SdN3FyeZvIKvP4AzPrZ5YGAkgRxPaQzgWQm7yC4JZ3k3zC7D+XvZJ170XnoH4
MLGM6qYHzUGD0WSdq2ubgAamUczpugFDM1XJkyWzrots9JLA7ZSi9n1Z4RaUvrxV
OuE718BrjukxXuSUiLZqCq0qDz8K/OKwW6FzanaF/OsDQawtL+JdWPCXd61siho/
27c3TR8C8iR6LmKhK4NQIitksyJaoFcK1xMX3ZxJVTOUu+7FGViHo3ORS2Nk/1ZC
fCtsvbQkP0N0aQp8K/mLADUX2aCimjynBB18GM00WR/J/1ZyhFxtIlnH+92Ln17f
VPVA4QAgahTeCUmwzjq2s09M7WqT3PjHgHuWBHfO9ZiabPrwC/DlAaIlP/02ip4E
BNZfhLaXlGj655InvUZx4jGJbxFOp9XrnoKJmfj/Uto3HHhzKtl7oZplDAFy6Tnh
XGWtpfpTgFscgIse7WW33PKkg0icWyLV2/CJ1t3AIvhcw9+sZPzQKaEk4pAr1CAY
jPn8SPTFBNPejz4VccbwuCiOYRvuGkGKHpBLa3CjxBzsP3wuUfU/9ZSSIaLq4Zcc
stuPmEzkX1DGPbkZlU0ZL6bp+UBC6l+oovqake4LEatjjJZxvz4LOlYW9pcyyaNA
diFO+gf5XrNGty4rxZLiK7mMt3g0ebUIQN30cZLI2rAQbgdeFD25fVvSSAiGfhF7
kJfH8qXFDV//FnB/pooHfBi1lxX0SrvkBOzWV5vKVtpdMOKlNd1xL8PmtHIcSe0A
hfH4NF5hhDZMiXPVV904ElSEMFNLr/TzWbSpGijR1ViilLhSLF9UKl3EmkSX0FRL
oZgGFxikumED80JmtRrmqVNQi0lLhF/t2x9C04ARZG3L01QIpv1//im5LrUOjLI2
0ZArnJ0idHk1OthPM06jEcZ8E0wlr4pkuCtZgtx+4lwyoFbLNIknTUb8EM4RLSL+
zJ+y4NetJcdz3yvgfvjhwz42Fj5XX3GZFN8WbXhH81HpfcZf2wOV2cdxioZ1WdGx
bDWnpgtqP7ACl8FsTxI8rHJ8dlmxXQJWyx7zUwbTIumoUiflYBIQj0vEi4FVfwtt
oq9EGZY7n+rC2/9Dd09rESqXKAN2/dAZuAqRFVU3j0L2vuK4Pk9XqxiD7ctx5r77
BBcg2y35/VIS9cqkon+PZps6gNsbukxPlFzelm7j2+KIpenPkkusgUv7vmMzokOO
MZDCxMivo35zbW8pFyXbWZLxQj0TyXdOPN9mnOqYw67HvoD6EZllq3GgufR6oNNJ
s/wdJzrIV40KqAPB1GUOH+PTnJcVvsRwUd/0mq6ceWXdM2bRJgWDzE+K409oZK0X
b2DEGBBNVSoM3QHJMzvcbILk+W8yVuIJIkEDqQ/iulNgNdyoEkRP75qLp3vHc1ND
kNY+A/Bmcyk7eV1efs78wPSqZaMK3mmEjynvqNlehV+SLE+DKSY7jIZTcUApQfoa
qfOoz4UTamJ5ed7vVaQ14fIVMBn9/Mu1hQeQdyheSoBKyJgz0yLQb5ohq23mTOjS
Wl2loIE+ZfyY9Go2paSMG+XcVlD1mQSfHDWeEVq7v9RJ1GYLlG8pWiLke9BVMq7g
bN86ZfUnyEgNJWiGFO3xRCrRtQ4KLEkpdXFhQ1XbhsREMN44pfVQR8zvU7fNUoEd
Eg3kfZERcIvCT0UHulT98UN/k0sgerpEauSy6+jd/esdznC7G+eMbU/gEllBsCdc
op2hzcbH15He2AlRdRKe+r2AaqEiaJeqSuXu9w/08g0U3qKdusG2UM1aCiOOjhzL
TCBYie+ATWEjT6mfSmm87Uk1PXGXu1M1hIs0Ow9umS535YuDx98YUZEIOoolB7aj
QcWxA6yo0UOav1jEDcdZv1NOOcazVtierAFwFlGgX27CsiluaMqTcjXA77qjoBKi
FsEJ4LT1FyrN7skmiNA7uAktdDNwpLMoGXXUVM4rQtHCvLwaKiLme91b5HV41yJJ
DMIleqNL7Z3PqiZaOpkISGQYFbQIZo76e7nLmIOmgW0YDhxT3edAfz5pZgFdIw0U
ZvvcYWs0aZwiG2AoT5hemdGNGIShRlCwilwqqXc7Jx7uzEXqTeF1rWCkySWMCj/i
EQaOO3qwUcdUiXc9sljGKn2kc0SAcZv3ayeJoyL34QgefuG9BdLgOuS9d4QDmBWR
5FmP9Hr1CbXc8VLmie7iYjlek1AMyz2u3ovUPvEbkI6z1AF1zWfhCLIc5wCBF1ZI
RP4xD9A3jyOustbCfOyOoY+wF0ftid/XbzNunJGsb2t3Y0VzFjGjzuiS6tp4Ou9o
MIKYYEMkVdqgV2Jwbxn2jGkGes3O+zFhobnGxijS24qmdVV8j7rO6fp1gnc+D6Bh
FAKzVGNM7k53eXVKEby+CHLiMIvvUPK5mtrHXyAMyEaOZClD2k628q7OEaBg03FK
96pvCDLyI8FO0itFRFgwdqWi/klMwB8GcW40Xoir7V01gWvEJCcz26M6CUBFzmou
ChUJsKntkcSdz7g5t2WW8Q/KFHrAYDp+g60dPI7f8IOV8xJlp9qtI650xeAb+wCp
heuMzayRP8hkSDMK9xoggH0FKgmiIBlpLOk9nE166cf0b59nALW/BjtBSSyryYBM
G17oO73S7ejddkaUfG/ZpVQ7eS5XXmCQhRQPf/HW3nbiCtQU2kc6nBwfKhYpX4D3
mbzOQMvzXA6bXodQ2Oe1fbB4VuCsIt/MbC59OZIDzt9bxT/vLGYC0FYhalHbnpMS
DZL7oaAVycPF5/2/NFjYvX+IxCfUD4o9efIaEpUitpac1IUqPMzwG4PSu6i32+em
XUSiMQU3l7tLgF83yqjq9WDZW5yvqcHAT0gep7qaW2OfV8pN+yBS6Pc9kkzZetqp
sHGudJnE7UbXWzvkNqMpZJ31rrIViejKEx0Z2Q9Vsuw1eX5WnndM4B+ipJEVXOme
JJuiyHoJioRVDb2M4/j/PBOw+yYFWFo30SbojYgdIeGZm3ycm5Q6GHIRbmYca0nE
vKFh1S6h1VX9jsuaLlLGqR6KDVl7pU7e3hWOEOYB29Oh0E4D+pv2dDG9tIHWrhUi
gbPkK3FV36EXfnZKxlrdlIWsP1S+S8u3/VDCL9X58/TDXaAFZcbBK3Wuc4AmAVaj
d0BwguEZI+pLGKBQUv4UyMB4ETrrAwpXY6kBn8VtXHQSuaCvMVPTkSTeVgOK+JkW
BWQ+03lRB55DIhcr4cz6Va4ONb5kiYsU0AS3ROq9mNkshDH8cPr8J9Jitk2Yk8e4
2nWrrzIQUfQlTSuvBvu9YLXvwkiDC+BI9hYV3HL1UC5mAG/DmG7wCeqK/QeP3PFs
l8N+HJH0B9MJsApGxALhIXq2BLsd/HTsPtIfgUqoKNyTIcmItpoHyd+/EIuJJFIj
KL1zJH3SS3Mqn3GcEp5yu4A9jmeJZ55GW236KfzBxPz5SVasv3RoSU6rBPe2fScG
l2T1RUHCEEA3SQYh1jt/JeyogMqNZCLhF1ej7vjv6ON7AWAumUg3TDX0x5CTMPAu
VKDOJmWFkuaSwr9zj9/jfuld0N1A9ckTbr6EyuFmN0lm+mr5msgb3rYLjz8YyufQ
MypEr7/ScKYLWnAvr1e1kXU9a8uwcCCXs3T92zIUe/1xBwAFxWq3ZRIz3BdT2kY9
dLCBuXw5vTptzOm2l6JoX7woCbsf1/8GlIARQ+/xe+cBMTlJV4MmFzqflDNvMZrM
hGEtyVFijqmhUK81dbzJ0j7PlQThNz9M1wanoPfEWQ6k3yOkMbaxvnRelkmIoJiY
lHGEpj0nM9RZZYN+FoLnd2ztkY4aKcvOk4MtVXE9Qz1Q72Kkxfi+/WMc5Jt4IO68
3eiLEp21f1pBTramM80gUVLRL6KfettGcNbFtKqf8EsMsw4bR/oS+mEQPX4WR/R7
W7ZjGQ0kV5NdiOuHPXbopsDD77dXV7fL2lf0QfGHRXvEQCt0b7Fj0CeFj/7Uot84
h7mc61+ZShUrJOOmRBAMJF71Dd2x6Jcl2i/lPWqJ3xLLwC6grtHN86X0H7meezyV
02MawOJj4DLwVRsKrhrtXU1y9nuI/zRdMIPMCAdZyMvAT9JAbzGsfEHJIAqEmCes
qDIqL2rp2USAjksAdjZCvSY7i2kpRNLJccLO48dVbHoNgKGGY1Uj2NK6UBChCwyH
TWOwMdNCZjWokWss+VVIkXedwWsoDqC9pYzINaAKj4B2+c8hPiNi1Ur/e1sOx2b9
TLKY2aJjhfU2ft4zQJZW1OVVcJbs/KOZyzfMRZ4XiXcrmnQ8xqJLXqqKQgV7mJtR
+AVk/Mobp0EW7c3TFKgy7Cyxi5XMRiUeT0WyffXon7PTc+Enu5X/riB1oPdkLdlJ
dJ0DrSEWYExA+Lhxhlmp8AfjaPX5/+0bdTk1q0Q8P3IZeSbvl2hTnWg6rkf8AyuL
VbNLlzDBNIgtIdrw1h9rVT1AAIdFj82Hl9ICDzxILcf2PFxlqDZ02T5hDBYj9rPN
30vLo4zcPGS0r8H6Gdwm8EhDbdJAFo6rE05XPBCHVQZQC+QfnKFM5lnU135Y1NgY
B92wtaI/2U2inzi7fPOOhHW5Odlevuz1U3OQcYuJh3Pk65tzS4rhdG0Z51KK7Ibd
mUgUwq/Gy51YLvpsRgzzIuH5c1tW+3OWlo4u/e6pzewHc0R3grS3zr5Odx39IiaV
prS/0WdvgHTLRnyiS/3WZT6rT9T/36AtYfM7ZMz+56L/OPfJEUk+CbSMTk/S7bhm
JrtxEvSBBQ8hUHCtsFBvzEVT+R27wfR9rg1m9a67X6w9chNf1JdPNioHQ0kyE5No
sB9r+aPUNCwnvJMU6GDOqWXnMFw6bx45/sc3+6GftDwCLoSHqSesZ+GZ4dyKNime
780DSRA6M5+wG62Lxin1ZuJSEkNGoXIigXbZmbIb7iGuNcaQ9WpjgjJG6/MLxBEq
BUHnlemyuhv9TemiOOgO9Rn7qLJt4EUEZdT4sfrrCJUTSL7UYjY3JWY+HOGNmEOA
iHhnwDhex2XDZQQWJiNxT3TIvw2H4IfEGVzTH0USlkLU+bwiyDuF0sdIVLYr5CNg
/sybVxV5k+qi/Rdw010zardwRG/dsIs2p538378ugKjejEy+1hbLl+e26jbVcX5q
pm1UnswKpkGApBGdGS1ESZcXCpG4CzMeY+7ZiAgDG7NUYKFzs/o3/KU5tPe8wcMc
cmZFfqiqUPCy9BS+aGbR0txhaoLEdtLNTwDf4Ti1niSdD8inq7tSKyaf+FtnQP6N
zqjYX/+snx/Ir5tyyI4kKy2zhsC8Sd/TBep4mXIMJHymJPd8UarYgOszkKU/12nn
E0rxRth0PXmGkiJwdtDXBH9MtyMwXo8O+TxGrWyEwmaW/EnkIbS+ogzkB7Xg3tpA
PjHt6jZFhGRLlTcoSeby9c/0vZDvajuWjbZFstJ991glvQRsm99jks4SokblBoKS
oP9IN39FTTYsOB11UOp2/C2gMuFbPhaeCeMYePTdAAbBAoOpfnHwIvfgIvoI+sAq
BBYELk95Sz68or54kaoBLyXRpNPzJaAf+KJ04hDKrhWoMbXD1auVjlFlpOeKfzmT
ojdV33i8AJJjicFGeIX6wPtf3YcFJsWngr/X3V5WCA4B/UM1EF36zcZJkwFaXKWd
3VWxua5h0yJT9Cfgyqh39JWWDe8NQy+m/9kGwumtUBIp6UvcPHsI/oyBonSZDXEC
BKxagQQq5fTPG/FsgNUDSm4m+GXVPFfoLdlkUn12c876csJYDWu29orJ/DrPQjXU
2yRIu1/5DxkRZnrUgvm5tVsPD3Qj4BTs9t153aFlVv5u7XjalWfDG2AHx52Y843/
RrsEHtPjQj9Udw8GfWGm3T/EMSzHj//MK+I6kgLALsdgDmHDTxNXP99IUkezO90u
4Vk92w4DNeoLC9NrPZpY4L9FqQ/rEUTKVICSl63Rvb1hLzQb6A5OEVSs5DrYcPzp
RLv5yJ2JII8OvM9BQ3BVBJsp/O12rEzE0klnWpUa2K+irflQ0T3vPmNtYJlzBoKt
cZuUI0DcVKh4zx64YfR38BdD2bxCEjuhdWZmvmLDFhZcDJHeKxovHkHiewzYj/O9
hhLEpdXJBoiYauJKHwq5V2ZkKVWVSgYNV4rRwWNVd9cujOsweavHMaU3eQI7RVc0
3uvTPwx/rvVrdRxUv+nLdtE8iR4Oox8lSmytK5un8Fvd3rH8w/qrk8okoA5ehb6G
MN0VZ2EfrA9YHZ7I5P5T7iY1nU7hrqmW21Gpze0xY8TruDXASV5JtLWSjfaEc3JB
UcCcTbGH3HBLgfzZIXPoeC5hUUWyvD39w2/56L592BfvPmvC7NNOVYMgBc1sud+r
Hz5PC62uLBV8KlMC+mCkjIFVyl6A0xOr4S7ulCktdRZzSW8F3U35qYK4ExK136P7
GlpXmYAvz9lZxNyTrTELIfhKx3UHXFXAnNcScI2fBOjuyRg7zBEx44gDnOl4X7M0
PsHQLTzkxDf1GoU4Peb/O7C/tK4g5nF7VVtxY5WRdmJO42RiYwdwnMfVT5rDvX8a
I1dgPS898p2pVWlZkFW5g1/Swh0V4C/tHBUJjGjkn7QD1l2e6X958Ja5sZy/2YIZ
SnVLTSlhiNfhl+t+H+z+Pl8Jg6fkQUeB65CJXMPtC2BTzxz6WoKS24XzfNnrBX9s
P1zCzZKY1g2VTel51ieVBGk0AxMhcsxe+YeEx+9joUV6eAalGwCBlULB0X5DIwR1
xxCX1aQjuJsgFqMdJXJGeqrXdBfNVsYtw4rmVP9qNXPWyAQB9c2zx31EYG64gxmA
oq/ucZabr1UGlaEKNmG+FlE7Lcf1XQ7IIH/59PzeCFtNU+5IEU2rbaavSLQYP4vK
CDeJbGVIkfj5StkP75ihfaTrcugpAYoTcNgLiJDT1BXf+7c+NClR75q6VC7tbhHT
WHMb/2A5TLJp0xxARNfgjX/6Q7nQ/6mXtgSoW9v9wS4I7yDH/bUoDY0Rla9vsiKF
+GBYGzWMzlybV3iP4Nz2n4hw2Vsh9ZeOPQvsMGTce7LeFt30oG495RgS7emup+6Q
j/LSHpjGT9ZEyWTtyd8H3xJzueNadJyAlyhkkHpXN/9jNIvQn2xsG0NFzWX/8sab
MtS2NlBoNNxVqfPcH5RnXQK5A1oHVi1pFDn0Ofswt0su73iuxGnz/AHz3bRGQSqo
ebnQgSneP2V4a5BXJ8T9FWyDFJI2GsxUe+Td2HqgsHU6an/EKgQrnDt+Yd1LdWjD
pNGaRSQMgptNIioAaoTCLBw5v5nKnCpCU0/E9Ecduvrlm88+yyEMX86Vf/WS41wq
+YESzJOCq3ZKT+naeI6Ued2xZSqHEYXB4uUijTiYHr5faaMQUXvtDkMYg2sODzC9
CXgknd27rXFnOVaneX8Nzr119ikb3NUkyX9Hoaoxg20+N0Y6jzVuyHm13rdluQIB
1Y6TTk7FqwOiMHGVP8+ZZEejNN6rHCr5pkFcclvu5XJgIlba9Knd9aCC2cbx56W5
rXRj70L4A/1vvr+vsnkpXBtZoPJlViyflMeO/lZnX/gj2QgNaLZQuwx2XVUSq8my
VMXYDxWhcWwxO/9rGlCIJmibvbhyVDbfPfzrxAkYZtne0MWb3eRpK27hivIRzeW5
1eFOfXk3o6Dh086gD8hu1MNmj0YhZOQgEQ4Jm3ITaVgA9p1g92ZixEY1uwwD+gZB
8UMQPb1OqGnR2iP6DSX+brdTFPqdu4mC6784MXQntUxnXeEoscfHTmsjmyU3crGe
zxydSPBPNFjhy5Z/u6Dl4vvfpBMrbZ7LzBUC6CPNTWp3LmcOcrb7+ypbHtP2FQpl
7q0/tBq0QHk6j2pH+7lWqRrEyiI30A/UczCDNdzLLRE4bHPmxnhqGfY8nXDxomNh
81Oo3B4o/EnX7FZM+6OESx/yN63FTRWdrYwaUp3VGsZg7U7Vx9/qkdY9EXXW0LnO
BXyQKa/oiLuqCXqR/LrdSujOD2K8sPxbFGCymhXerxW5+KrS4UzSJ70cF3EfiWpZ
ehv1tLmC74I6cxKUtkooZY0Vb43sV8lhYpGZsAiNhRnjQ8EVSm8BL/FyQsEBZ89O
xDaTHD/3voB4RRP1gJzLRudc492z4b2QkP9/572y6qm0rte+NddojVAl60Nkp8NV
L2vSyGnZwgxTetkgfr5xEwWezjayqO8mCkAxmgmJ5Uy/YlfqOfcaR/Lat5aWM18+
ih3DXii3Gd7DIOJPRQ9titH3+m+x1Pc8Q6HyttZMPSPXpa8rddiTSaHP+UjTfEb8
vnIGb1ASFc9K+AlRlu0NqL89VuTCUQ1Vvu+ZAhaO/4Xk3bshdeyG5lxc3eKm3e9T
p+r3LU6EDf855oAQ8nmftHW1TnGVVint6dOqt1bka3f2zh3gwZrDfk5sSLP/hoNA
/gn0QMqSpcBcNd8gHoyK4jyaRCCv/TLf1cKmG6+uchGlUg+x8oxN3A0J0L/xaTIO
YcNEIUPQgDg25vEyVDXpKG9LJXWDEY3Rhk/9hFuT8WjwZerfpaXrYwU9cXqnnZIE
nIUStNIMt1j3f2GNd5r+XdLD4qwZlDwieNrrsc5ibk+jiiw5HWgUF3JrVuoMXps+
rN8aMZEWndVBjmQjwoRQo3UCKfhP9+e++sdh0OxteUqzI4HiHD7Lx/CdgBoGRBkH
UItakOj2LGy59jooMO2wyfr0yiX9zD4FKxVe/pEGt43YgMAjth/TN19tN7yQui+9
LBiWEmSKWnU8/Kq+NcJLWBRmaFOC7FywqdOw+85aV3ytbn/5omssYRxVfdM9wjT9
YrILcTflMjGN9Ggu7VvwqsESGpek0yflyat/zsp2ySaff+RArYpy+QCjl5pP0u/4
bW2UYzTHf+rE47ThQsVmtTb7dip7xuT+t0t4pmtQgnGuTPi/g9NdFjb+Xn4E8bhR
58UYOOn2yLfzieG0w4h7z1Y7FsP5hGG+Idwm6NiU9l5lgXYTl87K56QyQAEPQBpH
ocDxworO4rMRqB7xXNiz/SOR0b5Ia63/NAnr2b/g0ZKWosE4fjaM97Q8hNaE4GNG
6n8yo59bbNY0xsmyi3hYqRiqn/W6Ipz4N9HLPbKkA39j/XcnOdDYQ1CThZWBUgQL
loXCSNLGFk9w5zmJAGbVVXbrSZsfOs3OU4R4Tk92xqXaXvix5JjlEWFB6U89RxVn
0VBM3IA8Jl58fNuKigfsP58vNed5RmNv6WjIHgC58VUEqww/gXdeb19O/m/+HJpo
P6udthqZRlwDYGDaLKeFS7mUmD/MXTbNwKLY4e7klhGbn/XfbYCxfllm64KcKVE3
FZYv7JNtmtMMUKOEAJlkzOYcFiFtEg4FS7Drd3KJbI/jgvPVhl/nQbhd3D99oBJj
VsZ5+wlRRwwgX7A69XlpMzhroQN3y73SP7hbp2cEwikNUXH3RH7/JAlig311RhmJ
UZjl/e4SRlsnGGC86jnmRGqHRn8nOwZrU3MCHUm5GzVV4WpVVtiK1Ilo0JdnQLRq
AEchcROdCSHbDAa6IYwi8TzYyMfKrE8kciC7+Lo29SUy4RkwQ0aSJj21tiZewfP1
VQvR4im79olPkhTzhSeL5CbmJECEpuN8xmNTymnyNLjSL9bXt3hCss8Bw6UMAwu1
axmNGhPzk4KgUK9dRnBhvaKq2xXM1pNpVC7nCprpFekC0NXs6uMIWpkv44leb9Lf
XlXOZIQ4zAZKg7cDr7h7WNLFvrqIG/hBqpLQwG1rw4i/uG6QDJECWEgy4pN6G2t4
STc9tKgDjdlVJb6MxySnLWsIFx/W4KPlUzqr3HjbEGzP3S0GztHvXAhEUaBPuOBU
XTy+0JOYN7PfHH6Pq8SEBSr3Jjje+0dS3sbIC+51ONIaw6Xaop7Fvm6W6xaQftDk
08TNOxgj1m5AFY8cVPqr0V93ouOFsL5zBKSH1P/mhPe5E/BVCwO79KB46KKhEKfG
JOOQnjr7ZeGuk8ZCCBFWjvl0xMSWIcV27MLlowt7te+vul/uq6Ogb97UPc+S5XzO
JWv4aH939ZZmDzA3ILfhbrYy26jTAAPTv7ftIfJ9OM8ZMwfVS8xNuqlkaWCmGate
74tpTXEiNpMEGN/SVXKKus5ddgNg45i5Ptp3xRRszNGuqVXhHNi2CCw3KdXZlyN4
KdqukkfK4ZpVbtwNEZ3JNQsOJCEndNocoQxeiO5TGBZIWMy+wjv7i7E6uc2OpCaa
zBhcziL6i+cUKBPww5HfWkVyAytwR6lOYw1I/noK9ju5X3VRgGkKkJ58+BCxNBBS
2iUS6jdsk5ZqQr3pPMJsE1shwgXldPH6tIJup8awbdnvI5xIhQAknrvTec7yyOER
4HijaVewx0sV6oHb8NaLGDMXZtL13tDKy+qluif8bIDGG9E6yvHZGlAYrHNJa729
+0skdTf5kC1wG8KCgIZL2VCRorDbfDTrbX8LiyAifMs0xSRkDIR0k9tZlPtBetYr
cEYvKHdnZ+wn6pIEZyrK7+Qga7J7JcuujMaDh13tGUxheyZOP9c/XfQ4/m/bl5Ag
Bxw/79PYS5B3F1ZSbvFmFsSih9q4ITO1syzxWhY6xcJg833H2hVwlA56T4Dn+rDX
k2J1aeLeduEtKsCsn/7eTH+vEyQMEpMFMD7e1OCvpb9HSd/NhvEIQ8U28APMp74U
o9qhJ8+zBqImzi1zS++Ms8dNa039hoV67CSLvsxksqK99/Cm3KKf9WUAy7f9PN4+
H68Ap5d9MesL5730KzO9JAuRkpdns5U3dn8x7oL5H+KNcI70wV8lWtE3p8G+5/J0
SYLnzTIbn30lupzrXFGEKwMAmgIYxtsl7kv0kMehFM4tXyJt/ij4h35fr28QBMb8
KIrpyXktbQUywwfRSrqr6i16S3IVWqSI9x2FaE1PKEHj870AG5PAN99/1szQYgvK
9JYr2TmvwJunY/8K0RXZUZAcnVNugULA5RwXZ9tthEElPaKNXu15bb8yH64F1EBR
F2Zopd/MDYB9O2UH6az4OLTMA+cWzf3XQTgE4dNGxD+PvHOO8/uqhC35mfR62yAn
XfBBRl/rKEYJ2VkGom+aGU5HDDXdgT2NfEH+0j7wMkNOONz2A8eviqtlJdUm9cpd
zAbUustjKYr5wk0bd8pkhHl5U+Tmh1x3lcPlnzjB6HQRgmCt5Vobf60UC/fvHNBr
KE1A+0t03jWpsOyraWGYFc2HzJiCXJKDmsJKruBxDSkfUMGmy0FBqNuBgsKzAyWz
yTkNBnADfTlfFZSLNP+sJE4jngXxz+bR+zmWIPGhFL91+cjpTyBSNt9zj2Pc82ze
dMxcla8Z+hRdWN4IiTAECvapqvv0hsdOLzdgsRkiSmsMEUoKKuycX89WW8XMcURf
4iM5p9i/EzWZFtmlgxxKdfmho3HB2+0Oka/W5I1HvnUuSaUxeVykIeLYGtFFy59E
s62ocETFu2bhGPDhAJpk7XCKmCAsyzrBFyfO79uJFoty4cKVonf31iUQ7Tqusdmd
aJCw6+cQNIJXzBjv2S84A0a19a7T+kPBZCPSJ5yyQIH557zgqcjNMQqXrP83k+5O
jHwEH0Nb5WIxBPVujLnKe6vKWzezAZtlu/hDFhhB2Y+tPcY0WmkX2VTYij4/TpO/
O+xBm42XsWKDvTra1LhHWgk0qdhBteHZy6fUINtTFsCX73jn9TBoiJPl9mcXo8/W
tHb4PzqlyINr94W6qspgxpsm6cYWtzpzjQ8Wa9XeCAbofUWD5Ee9WDJZkEshPOri
8HPXhJgYIgDUxoL2lax6LQthmApdO4x2vx2lW+6Q/IIc/8skl9eXAM2PCxsnTG4S
+3OzGS8VSLjx7Uf8Ny0s19pORYQMDs4cUzf4WOizSuQtMFaiyG74zY//E/AkGV/a
H4pbsWC/nFz/hW8jD1ZrsTl0X9UlBx5LC+zdxpkkr+ZZVI5RoZfgsLCK+E1g8dfC
gGZkcalHnaZ3xzhmaAwF+7lT8+pp07ghbZj+rl8P6pjjkkNTtbglygk31yZsVRgU
gfALcqKQ69rDD/n9pUv2p6MBGtcfQoHa15Se2UZfjGWZjjR9oDSZPwZS1u2LUSs0
d+I1i5J8XyLQvvTGKM+eo5zyBRFIx7p6XC1u/d0I/WtOGpWTfL2GjiYe/rvr7LT+
hKPDDTnCJ5QR3nxp1JzhUKtEUQgLAWLcWU5+jS9Cx8zq0JPTRhjs2XkvT7u+wqA/
A3D0ZgcKm07a3Ec8p1i/10PJyoMEpAlnbJqvJe6zIVX6r6wSRV0kWr7zkl1r93ui
YhS8L0B4Wb31IEAbcxgQRvIbv4mCymjpGpUgbJnZf8eYQOyFFB9TtMojvRpNB0kc
iax/MQfoPce5Clu2l/e8ULVIxjHjRNXqxXFEjoU+9FUGiidlPzBDEWycegqsvGqP
3vy0pXHyJCa6HACoT1smiQ0yx6SKIBywdTIc2+5FDj3k8x6aZb00/+TCJWCL6XmA
43ZVwsEgMGoDSoT/zvxWnsj2Ge5Uqks1PilxHZuq3DGLeK8uNjUqj3lToOlNFJah
LTZvr1VCDt5ILjvUiyPd5yRHXLFxO3zsw1xbhJqOerRHSERR5BCM/FE1YkaNf7uD
ORtSgIPoqx0CtV8Ly+TaZytQ8puG63FX7Ci8/rh/8j+RG/yEkcmDh4lTdWaXvmAQ
Ecwv8n/iOY5umEB7XKoYrLHy3kRl0GW7N2lJCB+Y/nSF5kgQ6vqktuZCP3yv9sD+
jOosM0Pepkq1o0sy6B1OF8iIMxQPfSN5OBZg4sbSQKjjp+5BE8c8LfraI1Dh3RGq
yV8GzjQrmFvlIkhfbHDkijV/M/VATPU5OTDnG5lh+n6GP3sA8pVyvBfoY2VLV1UQ
P3Npg980zX/gNjzvQYpO17v2VhkG/mz+LQ3N7zSMzjUHOEnrsrp708/4WbIV9JZm
ZYg6lYypRomjKGNfzq2tL5HWWI4qxdwGDR1CdPD6cdaOndbYL5Xg8mOgTibbM+AV
xs+v+8LhVNHtYgo0bj7qJRslZLTvicAuB3dQu5ajwwS+Qa0ZxdsZeVL8NU36q/uN
CJpzkfgeBcHqeaXyChqFa9/dHF+dMCF6f85/hMOgsmN/a66lqOQxOwS4WGVpiHWK
p/rmQfQ16+54QS9c26rchkABDn7JqtPMwYOxu24WjEXi4Ul0n02GIkWcDLs9wApV
fBl3tZj4yfdZ8WFR4UuR8O23J/tg+dv+1pwHcCbvsNTe8xh2Zn8Dn7QBnVFiac/W
KeerzBCCg0kgklLPU3vg5hcvm9yJ+DE9rbbkhq22be+lx2HeyZbOc0oBAjViN4xA
aGkTSLShPtlisxvGORKS3LPvRHpEoaaTrm504V9tDQLShEEtln2Oon58EZoGFLvo
z/IxA+QHhvaUQSMybSVmwEhkz2HcoktoCR8TsVt5M4E2L96kEjYM/q0viFhyKP4+
+t+QPd5SyMZv6U1tlOPAtkcReVz5wqpYB18VMtNwiRkbdRj8VLHoJQYrttqfWeUa
tvCtODaW9Inb1dwbevbfcLnGxDJvaqbqdRJSY8BFx0wB3Tqqy7VOtK4CVAp0N4nU
jJBoW19eqi1S28HyWHuIG2T+cGYNR8R6k0UEINwHCu7jOuD0+YfowEQA/yqgkJX/
GbO2gmZiPzo4tPDxwfJBufpYxjSYGTvME3+DSq8Eu+Zhz0LVUSVL70JmbKHvJTsn
Pz6vR9ae5JgA89E6mQVsih4/EdKmCnCR0bux687tNbPQfpCrIISp5nbd78ip2xxo
D+LhM8yelnZifjvoOio95ey9xLKSWsKvT6lh08VtgbeCoBKdBTzznfYAcCbgnwRq
ogYYH9cPKpxBTdmWtfiAqFg9tf9lfAKoNWN17RlVjMM/bcdtAoILTX9t3XPlhyiV
V/1uJ4AbVFaJhPG+xOM1Cv/SE3EBa6FSo6PZTvFWQiCJ5Iab7GpGTnRhZBP81gng
4JA3yMmKRLR+EjiXgOxjd7AFL+wQo539/bVx7fk6f9/+KgGCBdY/zQYrDPbArItJ
YR75ebIsXdxiGFdOnD/ZFZBOcUflPTbzNw9EvXK2NFcUQXZG+hB5+wgdUpenCIMe
Xdos9UAX9IsGr+f9demWfTXFAMd2tzfs2Vzkq5tmo+DnUHg9nMrl5vElq/GwCwbd
86sf7sMoOlFXJtno0BDVdUjgyZJJnhbSVOR8fHCuj+BVPieW+4Jvz9v7eoF2qqjf
RBVedFz5wdn0E4wWZY1DAOXzxFyKffFAUhTdh456nIjdDLOAAha0L1GaEbsrWBl/
e1Bsm62lxnT0tY8VFzapWJOn2fU3ewm4AQOg32yDJNGfZn0e1Y91Ot1i/cIpMyBE
8a7ONH7E8RNbD1Mh4n4DCMCv6jpP7tJpYuo0G98hJ4pOG9LaKojcXBxCxM7w22CG
OKvBpVRnCw24mY8Nw4fXg+l7dS8ZLd9Vd677XJ2CAZ5BSRwYoeG+sVi2QrT2sByy
zbTDL0+IWWrYVEquFh3fnUpqMRG+VNpD+IaDBMt6lDRnOyzEegzc60g/FpyzXAHU
E9PDtl+xCAJs3WQQjgLMLrbVpWGLLa7YhqrO6AzkeSKL1/BNj0E85/rbvd7jIaek
hFdTqjuc9ZPrMMuNJ920hWTdUVKt/tO0nB2JsLVWXfxAlQA8wd3SNYAmUOLTtrF9
UtHNnOBGBRXS6+GAB/a7ft9q5R3nn5gksbseeP/wijlJ6n+nHkaDURlQrBWBdar5
6MuRCBtcsxCXvwcRl0PWg2xa7/9MVZayPBDa0n/WKkdiLsiUhAUGVgFhQpjq6WJE
cj0Hu11mEBAyj8VlWMNvZyYzv8AMEXFnWU0j3ZCAhZhvRRlwidpY1c1u3JYtBeLg
c6v4BXpgbrpmh7Gb2lb+AYG0QOrm+1gpVBgDGuNcI2l6xLqFtfp0tzIC6Vw10sdk
5E24S9ZXJxhmF6YM68in4VxcT50ywsDRC0wcLWSwjnckqv+Iftcm/BurSM3d/F5r
Hpu+AMKD3IriUvG0qT64t4aPEW0fv9xJIvd9G7vJhtPPlULRrcFYBVPR7JzJgmbn
fzsRiWMDKVyPCtwTwEDikMfQIAwf0DhMrKMVdd/bsYIZ9lZ7y6Z8fFwDdJwvSLYe
Ypu1fpD7M7PQzaqyl/PNuNIQoWPtxYck0FP3Qq7ZV79FwOABRdosJt8f0UUvPGkd
FOUJFkU0w78Z2uRYPac6LJ5xQG3yive+CDvkLRrYdGmENSHEZRk0UBsdfL5EUgdx
sBX6u43IY+RoqlkT6jn7lPuZIY+aFRZf4VB7D5jGRCfZS5KZQAyCGJsGni6N7x/8
iBL6yk+60aOhbBb9UIQKacnPysIv/SpRx/n2MvMVKS/mH1P6gSiLAhcYZ4fe0EQ0
5WsEonG49z1OegDDQ9eJQ+RGKrAax+tna31Gejq6dYZoz+hd6cOlUu16ghKVeTaz
Rlung4DJBCYrRoe6lX3bZGr5shc2f7hLThg/N2URx8anNajP1RaxJ9MPaUHkT4tL
b03jDtI6oX9wSe/kMGlqMRBJTNskorSHMrB3Tkjn6tlWIRmkbGle6kS+IjfC8JUo
VQNuipBqvPTK45cNL7XwBvdXR6+nSMxSEhFJ9Qm5f9Ji3m7hSkztDhtWdwHuhy36
O707To2dC+lYsMjnk5heXNQhlvQkAXPx+blKWSKlV5VoZ5bhUlUi66pxUfDiwEcV
dm1C7BC0t3aVe4AW5/eEaY8ZBlEzcgwkuehqIj199/8sC/eYDZkMFq33ykGwi65N
cljzc28F2sE9/+TKqX5NaI9+kcJE/rAiHH9PZeAy+zDtvfNwq6f1wYsC2zcpVaJg
BdJm3GSTnGXP8UX6mnAoqWdfza322FfV9pyOHm8gxHnRXdYAVqNbMjfxNEHVM1ob
Rmg/91jwsgoLz9vB+/D1eB5/39dGlumW65GHga0cms6lj5kPUAz8RpaoNWUDJERZ
jEY7SELY4tHuuPNG0KLtFvmT/SbYa/W6E12bjQ5+gWMhWuZ1lrUDKWlAMl05yfUw
yk3ukmFZGSL7ctzTSIPzNiFKQ2uKphxIhb4zT5e4OotFfQM8VPJYBGEN2iZDbq1a
CDRHvcsIlxyr1X7D3oTkUvKsx4Ex3nGGDMbFHDToeOdpj9n8qZI6xisGlnjvJ4Nt
diBJXnS4hbqQNHT1OrlBxbUultASRasL+9SoYCuk+iI9qtG5gFRD0hBfsRSKKWJX
YIdGC/+kUvVEU+M0j7sutdIM6ZHRYXQ+DHcddUET0rMvLlB7P5D1jwPrKYtRBBxT
t1k3G8ybXnf4CCK1ypIHgSV5EYKpQd5APMJD1sd0kn4hrgOMyKbS9hQEOc/laKX0
VM0zoY5h90nwPREKbx/Ip9JiSVN7EwosHiInaNNUC1DVXCirjTAH1GY13tr7y7qs
4UUVhTdqJHC9Wsu6ayeVSE/uYVXuu36miKIdy3cZiG8OU7WF0u8u5/MbXpLpFAKv
48aA1ywLrqf+yKVsS4WuhCsu4qqVUcTxAJaZ3/UJ5S3edExQbbHU+NVpJpEzci13
5HQGPiV16tv2TyISac0l05lPOuHCRAvrbSDAjngpw/gAH5caz1W6H2TpzgDoszqS
gU2OHbIOWXQcm7QxpmkXK8EtKHPJaN2ok4KNFg1HtTIIGB52ntdpGizKJ/QM825S
eIMI8T2u1YbJAvB57MIe4ssUFAzL7O7mWVJQkcXNhFOIYqsgWQNwF7U00FDtkKe9
u+6Ei73+qHA5WRrxpi4I9Vjb/9/QKob3OJOdiU72teKNBrwFgVMjm3gTrY5XI3gc
GPomdDethRcUEApIoS2gZFRboa+zoEwuuCZwUssUrw88fgrUPl89eoEFXRIzGFU3
0XAWh+G4WvQq8XU7CEkv1Fro5MvpfSY49vBh7KOXPWn57P2fP7q/rPsJetEiPRdF
dwiouFbFeMx76/Jrz/iQ8OMPzhj6aaBxPzRgB5S+5lt1YdNq4EEJFxLLGuHGdY8z
29K0agLzQ136Tp+Kar7w1dfEPEfYhhZ1CLl5fkxnZHbKOpqO9GDDpjvyV2KcAaxP
+k+JPm+zx/cqCErvhjtdlYXeUiurZsBuwcd7xjtcbQr1DuxJtmG3XYZWp3jOKHJF
H0rLGFEbTS1VgoEJS8c0G8UmlnLB4SpaAqKy6Q85Y3xKIKxYTQdg4tt+9BMHKcDE
zA2/QOh8jl8AyLSNym/MxRMJRvoyc9HLGNfR/pMLTpAr4bXLn91B0Bocfe2drtBS
KcHirYzRzBI/Sjfu71XJXDGcGRqt9PtlG3cBxuVPLjtyS1VKfx5fn2mAw3ew7JZZ
6R1cmcb8mbs5oNlUFs6vkcVar75/vdPpyz+YqlP6ajxTAHS0SxzOQ9YBzMoJr5oX
KGDNWM9fH9iPZuLv3FCaZ2sjH3TjZ+ZIrj5tFH8ZqhHsFzzvZsn9Lla8wLarZ7rK
xr1BpxXFzIlEpmaS2lLFxqwsWAXqu7HReIDgdQQARgsO2ellsT7ILYp/3aAHRLCh
D9wfUeb1mvmvV7IStjD+CrPjKYMhBqfrGy9icwF2gmRF8+coX0d703XsE8yaFa5M
rX6ld/6COxaFoJo98rXnWpCTzUp22naSjRyrIthK0ZQyR8B9U6VIIYYBJ7e6N/hN
N0IIDoZjUECllo2AcQ2MyxFdjOHz+e/PhxNcdVruQODGHwoGJ4aKgL5aeE9zuwrr
c7LuREF4QuPDSsI3ethXXWB04OyHbOjQXfmVKrXu4OGln5e/THd7a9IeNDG1jbo2
KuDBFqGBMkYj4XvujCn9T/dvQUrDIBPe4yAdPvpCVVc/Y9T7THEH72C+lSr9PLnc
mtrIC4pLOuFWT/Cc5YLic1nEFL0yZXWgSDBAYyKnezlyQH5UxONC7sUpceEjQVvf
TGgU1RO0cSEbSCBXMwmFzT5psTo8/LvBpAixYexUqAvsZdSkYyCGuI4ZMcncq15b
t2cjQenPRuzYvrFRu3C/8ZHAvu72g22jRQ/EIxL67JA/43McjeUmNI6Nb8edFW8P
5jxYicy9Mj4/a2JFqI/zMX1Jf4yLWBPJUSXEc/PhZ64EGZ+QcaNK8dJ3UHrcOoLp
5P8hsMT2XSbNilAAz0Hnu8kmAYFAeum0u4sd8ZqVrQkY8WxsQj8d2gaILmMsVZPE
ZmChsw0RebwbP0QnzlLIDM8QbvUc+eRFwLYB3vkds11wjCSmW/XmxbbuXWE+L8px
n25MPOgH0IGJxKQoysaE06pbrAQlUjKUKp7SE9JpOXo9QYR1CK+uuMqleqtl1N7a
7FGdQBQPDzRgeQtFFV0qopR14K3sjDGN07Sbe7VhiDQlHeFSybAyEoHyrWkJFSQh
L3RYShnGS+pCLq6x3z+tOPAvzZdPMisRNMc36eTGQdaQQgi2QWbloVgYDm69H7cB
wrQSXwS8Zoe//8UF/sLTCYvfxvx+BWKX2pZcRUmjEZ9i6SiIUKPlOrFLWpMuzX/Y
UTjqrJMyQqIabwMi7jas0DjxmiorJPFVIWBlIv601L3dVYYI/iNBA4oVtsgFes9f
u0hPwG+lpM5sD6DdwCabqAiO+hMVMBNwsZgXxFRowiV+YKTxTcUgZ6f11r40bMTN
+FkbERPYxap7EH5ZpiTb0a+cYtv1MxdUqodfjqFZrpBqu8H7/Od4wMmMsmDoyEQ4
sa28OiuHV1OMi4Lko1Dnr6QJRdp1T0zNPPvrZkjKcBxWz52RaD1UByt0fQqRQrPQ
s3HGbJMf9cdki9FzLmGCx2RatHBqgEzZPC7Suz3ySXcbF/FVRGZfGJvGhlKtbDQ7
DVQDWI/TJqI9CHhstIVkBFU6jqdemeIb4RhLu4SIrx4x2dfgNOAICFuTytAEBTvI
ytYk0kTUmsw8piBgWr+S2nZWJVvHsfZAVlnWHHDverzyyb83lX861H2EWiq+myZm
D4VgENt3u66/3gnqyjSJD0KutfcR8GL+G3Fp42Udl5ZNejkMtu2yVIZbJDbbPiM4
IyzyzIZ09+aqgs6tBAjOgeAF8zvyCVOt2qy68aESg6Mh6HvypKQUxb5oQX6rmJF9
y7AgtLJ2lm/5E+H8Al4wKq3QFuv0zmYXIaqXR2X2aP3QorALEnEnWbYL8Se0fw1N
DJ0Tzi+H3GNcSi1//d+NbL9hYut6AT4MQMkqHxW40aZHWZ2zkj21oi0mzXOJl+fH
dXt4zSzIv/4gX/DF2Voh0tyXQ7yvsnqCG2Y417RBa1NKhNIpAm3TlyQDrvgssXiK
JPHutuHhjLic6s1oaGJgX3L1oqbxn8oxjRJi1GX/VohaBn/3mvJ/T4ZEh8yfgM8f
eiZ8wVu8kz+SViDFAcz/yqkloDQL9hen717kEE5yQBhCbodkmSfSkMZ0eNU69Lcs
iwkkNVhfWPHwb/TMNG28OoHNTsAzvaHR9y/QqbAnROiy6dnN1K97cTU9a+mLNq75
t4NGWM3SL2aHD4gEREaK5qhJDlMRBnpm3Jkgu+fQRdrQgGvR+h61pkCOlsC1xYTe
aNlLD69cEB9dyOJwyj2O1SxBy97NITvaWpD4Y6unppYmhXCShkn85YS7WFfrsLhS
kwpB321IJv4khYvXYfSt0Jf8xrmTZOyIwYZgOrhHDQ8hiMu9YTkkfBnsB1BcALdP
GtfqtRh7vcrUy8CMyzhEFuLAotoAhPE+BJr7JdlM15OwXhV/X+0t83gP9tkD2nrH
ORUNfZ38pfo2w6E3IIzb4p4rYZEKvwiT7RZN45+OUQHv8Ka02ywR7hLmWciaUAJ2
HhBw5KbpvYW3LX/kwi9YvVn9O/VcBjITyJ7Hkrt0SYfpcOf49wpEP4p086oOtEaA
v0lSnWMRqvSxKY2OvS5LWcUusVL8iYywx2hcxITqTxOo4SzNu60NBn3uMztr0dtN
6GQC5eYaY7yEPkanGqD4lyFvLUTe+UkYKx/oSJDik+DejL9nac5a4D3wLSQKZij8
dTJ3p5GbhL0S9YbzHAxtVh/25EBS0Uikr4ykOwlJD+q8mMmbYRnpZ4fPuFBtqL4t
iS1DPRBzbEcS+vH9Bd2f+O5uY/ETfkj+CZKOGxbhpBqRVCXuuUGgggnb56g9jL84
kmNDjAMsO//LD0mOSVd8woyzT/qFrK+cFnER/aFKxZcBbQoo7skh3S+mzZ/bxtVH
JB7KlJA3Jg03o4wq+msN03hOqIeUbeuR42f1GW+DwpAlAH8yJ6LXqAUaVZsq5/9l
dWLU8xeQSsyuHYp31SKCLqoRMs//HFqIV24xBDBb7UvqPQGy3zXJtPi29QZ5AATw
yEBQ8KbCIOahlgMvU/i9F2FR/Q5VRy+f9Q4uerh7176YuxUtada6ZkrVVL2LSi9U
fDcKQtwA8/eWsTfRExQU16RNg0C5tOj/7Y58x1IGI3uLuIawWeSj6apTgynOd6ug
zujLeZDe0GBJ+ZXk6QKIidqavBKwpWyp8345XdGSzfU8oYl+7hWaXwOFo3zUzYfK
f2lzGa6dwG+FrBrvPjIr8HWAfr5FCxkMoleJF7GlVQhXo5FX2WCYjJC7yEA0t9DM
ZUli9pdw+Yu9putTcVQ1O1gxn0thUi6nEiw6HdVWhhGVt79GgsIjVCZIKxWiZnhZ
F8nuFWGNgFUPTARvtc/3mkwawlso/btfMUGmzvzXNnD3zZoKURDnhSIliWJex2MV
E6C/I8Qz1PJxdjkw0SHRVgylz+i4I4/O6NfcKrV5NJ3HDTqELaJEAyUbv51LJRxW
RPgmTZVXRV2/w6Ok0lBRSyTw8P32dD0pLSxLsHSWcYKvBnqWnrdbpNztvZUB1j89
ICZNEbzBW692AC9McBlJNezCWZ0KQEtTg9LWVYAZa5aTurBXoyGY+Z4zfkEy2YfK
7B/OkYDmc7SOfqdWz7rlA72xGW9BUnzmmuIyqmxxuJRZmwzOIj+JyvUBP3i/KiT8
AOFhYhrBVy9uAwRXvhawdDUQDR2FFF+q8s3Bo2RYIDKd4WxCFw1EeiKOiMXbFYCi
cFJAYW8GvtTH30gkVR5IVUpVvyn7NisVFlXtFUw72jKPvKf4jUWmf6sd4/jesTPc
QvITYoG3C1HnpMALFLT5ThPLdw3E815+KIBCBrO3ePYdiibUiEioNC3xDUEksWND
fuNMEcIi+uLwRZJFqZlNooWbjGiSNbSzHWnvlpyKsJYBvovCPK5Jq+WH0jcSJ8EX
6Yi3LRnhOvTNGY4PyOqqj8MM0GhEJPI0qmsxRCOC+phdQPXojr0f+XRaEDpoA6CI
qRwmynUkwHuk1VyUgSKU+d6HsQb9nyEBRltOQO5Z64/5vJYks2N2l5NwbjI8C2Cz
r/WYh+Oezo917OQ6ZNgBbE8F0NwJXNn7YRkOAGDLiucce7ewIRYaZdJ39Wm5AMo9
al936RabLQzrKLBvN5TBu+CXQQaoD3ynTFiztIcLJD49op/RcUML3NDUI5c0oOQH
jxcJBkovqJFV4KVYxUDrE2P1goRZXlql3Qsr6+oTTqNzjxHzm1Zl+iPRlJzAuj7d
yok7ujGRyv/8U7rajPvYEsbrLE68OLoSkK/7oz2ipk/d3kR0U340Ys5DP5BGDPQp
CBD/kFWKzlLAFWcvQdYemJ7kHKEu9KCc/ouvrOX2WbVEIeYDwN13Y+R4Af8z/5wQ
2eoI40pkISRi1Ay3iam1Eg==
`protect END_PROTECTED