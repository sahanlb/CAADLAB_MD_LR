-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qF2n1DA4DF5MfNx2qU+9uNT+Usx8znSkJKdzGkX3yFlALb7MlQS4zUH+7th6oREu8/m/ijb0vNcP
BrYWeIGW4BOio3Ae/1d0T2mu3CD/amz68UPHW3M+gRPD4qXfWcQyHxz9EMhH363IrhAAdd7mGBmq
Rvxablk5Kz8V2sUtPZ5pKc9sqEQ3jietJKslKX3c/O4qGtmLAso3HpnlCOQft6TNDMm9DvB2Lx2m
yhWhsn68U9GtryFj/p6TSwcK4T8Q/fjmQxZxE5cbUEO92PzUqdwtjeSHttXIaqsuwqNK2/A50MTt
3Jkek+n1CMQT+VC3tTMpvNnuUYcz6ej8H9Ou3A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5648)
`protect data_block
nqDgRkG2uWeAVBk5W+KgAHDWA/RUSxV+PBTgd3qbau50rhfCUqjxyUN1+JKfah7DXWbtJvRLG0r/
0SRNtLwVcsmiy8EVPRlpO/EfcXO4N/0nbmQiSpvjB07AkHdEbJBGdklpOz9gJ0qCtS/G/fB//454
1fegTYGvTluB0GQnhwgpTvexLB8Ek7SgtnW2IyzKdeqpDTPmA4v2HMnyo68jH97V5uvhHr0NqEk+
zvYaYCmJEoZRwjdDTqxO2VBzAR/EHRUi0RYxsChpavKDKw+SYFAXQUnQvZ7qtUu7XE9VkiMB5DUw
Jb9lZ+oqmor72VcgahzxmKdKtOgWClqEgdoptw9qodJsAeFQ7vKRErCZz0wmCcxatkZuQ59GmaNr
S8IYwBqyeyRTkFRFSjYlKPGZ5wIJnkS9fjfYjry/xcft8DEUJya2Njz2OjgvaAvD33K7QL3jWXWp
64+UOIRCghaJ814pA6pjDV77ToG1se9OcjWhYLBjd+rq3UT/qqTdtLxqaZJiBXIzG/GU/Ofa63D2
cTPp1yWRGLcsjFmw8Fan75kMs8uR5l4pY4H9fR6eRlSa/3qtIOo0PhxUGR09OpnDZQt12Zmj+qqS
kcUU/p6Sdih8wOyRjPU0ubppwMZrPSQV2dZVGbPrZK2gyQhIBaPUXN1Ydas3o9ttJDNPXirXobk/
fzzOgs3BKFI0ZsrXwOPsFHTg7sw6EzGndNZuZlU/aULdNKJJ2viKxXMTfSuPdP8lPK4oFhp4Lm4T
0PT6wKmeFHj9MTSINVokF12NuuXOzWVPR8irRECirY6PAk4BUkPtJ5WgfKAfLkVpgSTKUl3ifxbN
6S5q3jrF6k04WBH4QHar56cNo2zHQRDiFbCnyL8tS2/cmNbcBMS2MHRbUo7V59xhPtxjkOAdKgnf
DAhQsGzUzNScmANaZwKygdY/EKIjnWXaHPb+0uSsxydRCmXATuwW5uw++P1ID16gE+Fx4NY2kJwx
KoZwN7M5gxLn5e/qoZtGSY8KnlEE7MVUkGVNuKGpCVRp4rfPCmdnEpUtbZiFU6MCzfp5YJwmsdb/
ISha2qAArxXOk+dvLgbrbUFG5rnfF7wGY3Pm8Kal39rDXwB8Ysa8LZ3I8nain5EBcgYT+ytrHrYw
TlK9PQdhVIvrKLPAaKP7zTsLOdSlJaMAAq2ddIFN6yLC+YCSTZ4RQqYJyAApnz0P9BIrDe6C6TDz
z2I/h6zMHNeUaO3UaOuBWJQnJ1O7BBoxs2nKAnKfgRVj8rD3N6wIgklH7S8S7i7u4p5xD4x0Vvir
ywsnKvvfPuy7K62UUdZkgPHDzPTJxYmXZaPBc5mKvCeO84Y0RDErGNI6ma6yFUeeAkBN687A7bRl
zpECrPMbOmlvp1PxHbr150a2EuljWRO9XB6HzowvUdR7G8Q+gMVNz63v2I7uxRpgLIBjwjXcNNxb
uS5Iih4las6efaQ8CNKabh5bLXtQaxMZKRSBFa6YwTMvE7uaJKrh149yYp23qOSvebcdp3xU209K
BCDKPEJIuklusQkhrRPzeLDO7KJ9zlKHXcqZBp9snq79ScZt/YpLiNRk4/d52uGqFWFFjtGZAbSh
stu4hkqNaLF+tmJwuLuLEI0bEIKFZBrlYqFXqzgoSMj3mBO6n/LyR9Gj2JH3ndVQS6LbAVb0DJRu
+LbgCmZ1/RmzxrAtwBBelv71OcL7lbi+mZIEcOQjciLCpsGwmRMHFtc0kDjZiPE/Puz4x04pATOU
8mQlQuZ+mpNfdJNUnFyb/3iVNp4VOgckUz3G8DFuNqV+VIlEtna4JNh4gycwx4ZwwXSzLE1II8NR
buboWS+s45eBJPq0LrQCZQgz/gaO/zlamssWVWrvYAmdv+q1VWBkqN2DeBAUgWWdlhI7D2zZCvzm
tHcCOG3v8VEg/ivgJnRapPSS85goDSUiHgg0j+5aLSZzL87qADOyU616d0Hm0tyuwacmoMMNAsNl
POhdtVdZbnaZRcgXWHWTEtbPoR6u+ALa+S0x37QgRHWk9BL+6wli3FmTKB/rUrgr1QpdXGVP2bSB
gTbP1mCKpPSf2tv95hd5FIZlOyG/er+jkLkYyjDZxU8E1aAmdPqwHLFk609mxks9667yEC+eQKgD
0IfsFCAGYzNPKacFKf/2sMLoNI5Oi798OetC9IdKqg0E6SQz/SYFgRaSHd6FkA2v+8380/86y2zs
1nPk/kCHuI3WvATouh2/vepmW3+gZPAwc7k5qd8y4K466bxT+NTJWVh+4a3MQRhYqD2m2+3kYU3s
naCJUICPIUeAoHwfPCQdANxeK/H0EiMcKdtpiX//SI76RcUocGlwug2XojF0UbZf0RI2UCYlzSHK
cKxACJwyvdGIeT3u0cCsrQlpbUVtg3TkawnrR+y/Ho/Rg36dJd5PPXAKPqu64TMFyQlkUWSi86HL
pg2IvOReUc82RfOS3Vrrr1s7S6Qwe5DqSxOyhIXG8HrSKbKh7dAOqJe+xDzrWaFG7kb2Akq2DfZe
HclJI3oDfWDMdXe7lAG2rgRK0AKhGiyx0ZNhM3L2F0c9Xw4WmlfjW8KITk4/grJdMif+qeC8PZvY
3s2rGV451vv7AQC+xif+fRM86jDW5JdmeA4RQLfWuW6QwGyv54FyCLh58rFvsmlKKiy+AvbAuKaf
PrCb88nJdvAk8eRZzvzGKqaj/C4Bk58IGDop6aOgreuIfmcprHAIvPyxRG8xARyaXMbsJhGbmQ1h
U9xSw2DO39tb/VeVMcBsjYKV0TTHzItoOaW0qoBjymucXCZfCGQ+D3OdkwssoeEGxGx+co5BDIDK
vOzQiJwzZayHbaCaUe/DpCV3UmJU0Lfr71J1K/jJLVdR3dIQOQ+Ea5KcyfjcJzObraR8JKsrEohn
Z6KZWNFBHNDOkDTbHqCJpwXDVEyGjXZjzgnd5OvQ7pdag30/7szwhUbn9xFqj6KtQKChlqAdxKIj
XPw6BMsUdcmEqjbE8MvCtg1iFhx6Qg6eb2HOYKkLc7Qy1I+HLOER7d7MTGSYv245xB1KZSLJPNNH
Fb9wQEOtfqhUSGTcfyS/+psSYCtJI1MIGoHNPzzoCCQDd93uhikX+FCesANRvfEZjLu6qf3Lv6jL
qRKq8BmhjOEdtfso4GW05iQgu/AlHn42Tppq5Kk8CNYtwGLeS8dYUgqBkyJybCb8czMUYgCH9kMB
DZH/fQ52Z/oOgWlDe3GIpsRardEGA0rhm7XIbHFc17aYNN9dB3jlcFZyltLIdJNILzMDlEmy6ukV
2ESsQbdLBT/DFWKeftsAaYWSr5w+ysknIQQ26F+gH59Shg7CbfZNcZMoZeBuQoQiXB1oYQCl1q1e
2ZlNm1k40PFgFs3ggxVGXMVGHsagFvDrmMys2DasL+7fECqvb2ovlpEwCrH7Hrl+yYRyaq+LFZY8
aOmFNjMSzzkOk13NCXyfE7U1+BEwkTk69OG/YKbPwz4pmDOLqrQK0qTt9qN5rjPYr0U8Ra9st7pz
JPj1ReFRSTe4c6BwyAwHJeax1Kl5ow3zIxapSjKwQTnHx4A+wW02nLAIGjd9HWgr+FatPbCyn6S9
xu5gsWkLPPw7rzDQrvlpREuSypGwzf4WMDu9Sa1hBZgnEeZ2G7md6aBseQdszP2DTos22NjWfqfq
0q9183I354gQuqozdWwfqMdJc5Mt5mIV1OFgThmGVlLKKAtqcm4qnNn0Olp0QLgKlnTXEfA5X6dp
Ml+VfbyybohCD59kaPx00XNPCInh4M9ATZWTlSbNu9TzfYh9utM0sX5rRFSOxq8y2Xystrw1RUO5
MMm8VDyPZYDscwqJet4alQx3XOClEuQD2TMEXIYuwP5qjxA9hUZ8smzfJPTeo6+GLMlHOpORJtLM
r/08UJ2Y06WuQgOgYW9L/2jmZ6fkJk6yNWmWapKApHL7VQJuHB4xOd1c+dnETthBt0CcAG8SRWkt
7TLL9bTtv/5UhNQtdLQZ/YKColfd0cXj6/Ta3cjDcJ5HPJ4xMMjNIpaIDne7r6Kzslcv1eYTHLyf
JZ9v9uR+kX1rLicSvw5QgSpzwM+kniEbMx/fZnHn40uNR7wP0ARNJ+7Xw02kQB3zybqVkv0OiaWG
8xtZ2n6fhf6aWysiSyU0b8aUywXbwZ+OVMyeaV7GSTp5nJlneh9p3sSUPPk1ABsm9NJq21WI4eUa
fuaOyX9N0O/dd57/BqBYNB0lgYVPq4hdZ8pGFIxucclHOrB0aFWIM16gsKA9a9l1D+UkFo6tOA/P
2ZsgV+f9x+EnxlxiSJU2wd8m3uCJOL3LKBtdFgIIadPH3tK5htpWAQwWaqYENe8a7UTsTx2yAwbC
YWyfBQuDAXmoMNTjFGCOA/7LZX0zW434qOcmkhR6lapYXVyoV8VGWBdrogdRO0BMbwqsIDoMBiiF
i8BEOPFWvTfJVvp2D0l/nKrZQXZALfRtGAwVhQxkaQqpCMUz5zbsVGb9CUhA7Of4eSCAZ+t0Upe+
JW3aa0C2oks/k78Hh3HwQZrYnT893/OAbR7fTAAOLmXZnrVVg3O3XEaUI24cc524z1Cb+w1BTHod
M982YJbetJxaQvDXPof5+hLi9Swlsf18BvqAXxbYj41xdM4s8VrxZV4dhgA3/BFLVK2PG56fkYCg
YtCnOkBlLdSR/DhV8UQ4WDTCTm5EK2xWoR0KOAvC0mq+QECSjOPi8BqGt1JUJXji+2zh0Sf2yCHg
P7lpZXnDK9lJm7fz0QsAkHkMGd4A3gad0Pfm66DJMuKUWJ/djxGKkDjaTdvntCAjIFFNUMoxd+ae
G0gzb4p4VLBM7LB08ywZKCOh0QtAbHx5MkQElMLWGVJ/DA3MQgMPADzHrv0C/FQtF8O0DPTEQo0K
lBgXOYuDQNnNR4uvWg5FTMHw6klxg9HLJyPUUNnNiN3V6BKTyK9R5kYFZDzkVoAQra5tBDXMCPFR
3b8o4sXoewMJhfUtyOx1Vo7Qj1gOFYoxZA1tB6YPY5gXcY0gxL8qv8SeAZbJPQ/7Ke5csAuScUNa
rxcGFV+GU8Q5BKJ0cNnB5uSFcSetF0lsoxTYp4HUNmjFNV7p2qRL7wQ5PQFUBhVPE9bAhLXgXWlV
5es/gfFnvTe1PBNuGWCI2Dv47kQUeuHsF8KSJwR/SmdWup7I3NO+DHbxpfo0/OUqtik2V0FIiwCD
wTMwn86oWums+Wq+kg/Tq/VIcjXnTvgl0/EzGblvdE9+CbBOsQlUk/QYd9Z/2Y10E8FV0dQkRk57
EbCwnLReVNtUEYsjzdglgAQAZCBXKpBj9E5rvRyNSZJjLOVMKbhVmrQiLw0FzU+ceyRYyYNC/M1v
uH7kri8gDTjz4Fs4vAHcdBEE3nRDbxkoOobtdSCp2Fvd7EWlt4FB7fZt0ZOVEzJ8kaZe49dolQzh
udQzCttmgcFEs+toSwQG/VsJZ0xg5IFWZvcJffMY5dApG3ewYb11DOwNEHqaPESo0MngAwTaZWc8
dtgIfGLTNYZQK1AYSdNA+OdNSUo1V2uRZIMgf9WxWkqVMNivA1RpjuVM4ONZwKtihqoXUj0iaqIj
Q9re7x5uSLXIGp2+82CVnPYfJkq0ZpA7ukjO+TBW2KYdlrRqMGNbw9I6WpNTZr0l39ZWy1PFkHim
i48YrymmeHvo8C/2JLa63hQlHp4sShkuEV3WvdX2T2SK5EPpZE7AZV/57UeJx7zBQ7xkGEJOq9LM
SNMq9W0kcpi+KRHPEf2byYRlu9OaIUz6nBUMO+eumIMCK+KgJyUOGkZHxS2Rkv2THxhp+NLZ36qW
/8AnqDVYyubHnxsbLOoy9KfjrB1Wr/wxzh5mSslsPlyWdKJRMpzeXVBANgP56Pvwmo/DD4ovP5nK
w80vcxPjrvozr/3SPlg3W1R2sDAaOmI0xhm+UdTeL9MpedUtRQ+KboZurQOsKXOcrW5Rk24NrY3k
utAwKRCPSPP1F7EeznDXo9nqfMs0jKnLRkBdFljna8LJmeQU8H83tU1jbD25sC6n/LQMrSR2iiEl
QkUZpI1nk6NnkJDzTMf8ovhdChe70RXsWy8DIGyYTlh5AkPWXRRHV0TrFQufnS3EyolGWijfI3B5
+PDPaAJHZXwaF0xGD9hkqjqDWP7M3PHe5i6hq40PFTrA67haDCgb6zRMvdUlHvMmkWmq9CrcsEGs
BO3d0Ny0ERLz6Z07WMCCYp363WrY5FJ8XLMtNxTK9tza6gsFC+D5aRmVmG/zy9wVAAyQ5PmJUcoZ
M9HObVJsHtc2xydQSVTWPN0Nn6/ja+VP1tN7Jz3Gr91ZizirMwgiLexa3aaAkNssfjQf1/jnoUca
2TghHFGiMe9foMFIHO3XvNhVDMhlDqWN/F28ZjDU2nCEl4YRn/LkPosuaWL7o7a3mYmXY+KTX8aC
Rg4UUHC7JTQwVxb3sntu7z/j4UeCImR7cAr96cXlV3WHTiUOoBlV7z4G1S7zRpIkseRRPszMKwZM
tbgTAnRzFQKIHmbq5ot/PLxjkGuD3gPtXcEYGCaG/hr0ovLkM0L1cQ4BqGoP5TE197ko3Eawq1Q0
9PLLtFWBTRv31aiLWWCqMp2pTfNE89v9OovCir5bD7JG3OIKMPqeeBaW9wGwZTlLBfuDVqRU8bxh
J/lsMBTDlGe3d5TqN1lxyo1YdHLbRvINxOKPkT/TjUVW5BoH7cgxUgNG777pmjuNULqFKMyLEU3Y
enny3aj+lzfSt1k+EK3AED3pIkkj/2E0ihqWhKHkALEnf4dNA80h4zji0LTdP17NYhlUD2YO4uDK
iRhPFV0TyT1fQS295GtjjcNrln95R4ry5NW9FXcGia8NoABMj8o/PJL+e/jILpRgvcJGeUgz8u8r
uSJexvroAeKvJ44R0zhn1q/toYbIcIHURzAiNc9t3fTVU/BfHD6idG5IdkxMe3lS8wWyBSZCXDp3
VErJJKQU7umNQ3st336rHFF0YJSq2ngJch+S6wR1uhd7PgaBcbI/fPpka0yl+Jpjjug6asuJFyxX
m5Yv+yOVEsq/QS+pHLpOzp++t/j63SuYckoX+WDi92s1YazF8X85AtiIlIFvpNT3CZ6yuM/kSKBA
6jOS0kK/2amAcKzOlZOu3d+AQsgfU3RFH4oflg0e9tGsmpgOYe4N12hEjbzBvignK3f8A6pST4QE
dB4Vkd4ztXVmbPVNqDNJ/S3KQzVPaTdXeDRdyjYzARRuBko2ktvrZcIIzf7PCahMRUvmCtJ5Ohu4
JUpiZfDM3LLjy5tCeZ27B1wG25gP39E9F1Lumifa2nHHdHzDRJzdU3IgkIviNqAqpuacV9wV6srD
pJeuQmUVlRV/8EmacPz9U3SCtPuBJFSzimJgC727e8q/Sy+eK1YvuXSqDliXEL7CYK3if/SGbmbU
h67Ji9l0OhWcKLh6FPG+ok2l+yZMopGWJbK/t9RBTYEF6/XDGkTQCP0aEVlS9d2igjEe4bdqmIK1
V07nG8frJWHff8IJubjr2sM/xnzlPqsc6ekcJrWrXai5YVEiJeMIJpyxpqYjj6lG4Kp2zSqVH+vZ
rkWdByM=
`protect end_protected
