localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_IFFTY_CHK = {
  {32'hc1aa0dc0, 32'hc38220b5} /* (15, 15, 15) {real, imag} */,
  {32'h41a2a940, 32'hc0413a20} /* (15, 15, 14) {real, imag} */,
  {32'h42085f6f, 32'h40a89e96} /* (15, 15, 13) {real, imag} */,
  {32'hc11a6e6e, 32'hc0bd3cb4} /* (15, 15, 12) {real, imag} */,
  {32'h42a7e32b, 32'h422933b1} /* (15, 15, 11) {real, imag} */,
  {32'hc19b955c, 32'h40b86a98} /* (15, 15, 10) {real, imag} */,
  {32'hc0c61be8, 32'h40b0ede8} /* (15, 15, 9) {real, imag} */,
  {32'hc15bb12d, 32'h00000000} /* (15, 15, 8) {real, imag} */,
  {32'hc0c61be8, 32'hc0b0ede8} /* (15, 15, 7) {real, imag} */,
  {32'hc19b955c, 32'hc0b86a98} /* (15, 15, 6) {real, imag} */,
  {32'h42a7e32b, 32'hc22933b1} /* (15, 15, 5) {real, imag} */,
  {32'hc11a6e6e, 32'h40bd3cb4} /* (15, 15, 4) {real, imag} */,
  {32'h42085f6f, 32'hc0a89e96} /* (15, 15, 3) {real, imag} */,
  {32'h41a2a940, 32'h40413a20} /* (15, 15, 2) {real, imag} */,
  {32'hc1aa0dc0, 32'h438220b5} /* (15, 15, 1) {real, imag} */,
  {32'hc39c4dd8, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hc231d957, 32'hc30e3982} /* (15, 14, 15) {real, imag} */,
  {32'h423d0862, 32'h42678d0a} /* (15, 14, 14) {real, imag} */,
  {32'hc20f187a, 32'h420cb541} /* (15, 14, 13) {real, imag} */,
  {32'h421d89ba, 32'hc1acea98} /* (15, 14, 12) {real, imag} */,
  {32'h423913f8, 32'hc1b00685} /* (15, 14, 11) {real, imag} */,
  {32'hc2b6346f, 32'hc0bb0a3c} /* (15, 14, 10) {real, imag} */,
  {32'hc1c718bf, 32'hc2668f7a} /* (15, 14, 9) {real, imag} */,
  {32'h42040500, 32'h00000000} /* (15, 14, 8) {real, imag} */,
  {32'hc1c718bf, 32'h42668f7a} /* (15, 14, 7) {real, imag} */,
  {32'hc2b6346f, 32'h40bb0a3c} /* (15, 14, 6) {real, imag} */,
  {32'h423913f8, 32'h41b00685} /* (15, 14, 5) {real, imag} */,
  {32'h421d89ba, 32'h41acea98} /* (15, 14, 4) {real, imag} */,
  {32'hc20f187a, 32'hc20cb541} /* (15, 14, 3) {real, imag} */,
  {32'h423d0862, 32'hc2678d0a} /* (15, 14, 2) {real, imag} */,
  {32'hc231d957, 32'h430e3982} /* (15, 14, 1) {real, imag} */,
  {32'hc38441d7, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'h42e6e320, 32'h41c4ea54} /* (15, 13, 15) {real, imag} */,
  {32'h430341a9, 32'hc2b331cf} /* (15, 13, 14) {real, imag} */,
  {32'h42cfc984, 32'h4284bbc6} /* (15, 13, 13) {real, imag} */,
  {32'h4071d5d4, 32'hc1694bad} /* (15, 13, 12) {real, imag} */,
  {32'hc2108ca6, 32'h42851603} /* (15, 13, 11) {real, imag} */,
  {32'h42ad334f, 32'h4208b34a} /* (15, 13, 10) {real, imag} */,
  {32'hc29d8e95, 32'h41430050} /* (15, 13, 9) {real, imag} */,
  {32'h42217a62, 32'h00000000} /* (15, 13, 8) {real, imag} */,
  {32'hc29d8e95, 32'hc1430050} /* (15, 13, 7) {real, imag} */,
  {32'h42ad334f, 32'hc208b34a} /* (15, 13, 6) {real, imag} */,
  {32'hc2108ca6, 32'hc2851603} /* (15, 13, 5) {real, imag} */,
  {32'h4071d5d4, 32'h41694bad} /* (15, 13, 4) {real, imag} */,
  {32'h42cfc984, 32'hc284bbc6} /* (15, 13, 3) {real, imag} */,
  {32'h430341a9, 32'h42b331cf} /* (15, 13, 2) {real, imag} */,
  {32'h42e6e320, 32'hc1c4ea54} /* (15, 13, 1) {real, imag} */,
  {32'hc2825618, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'h42b90f00, 32'hc1fc4d48} /* (15, 12, 15) {real, imag} */,
  {32'h42b99074, 32'hc30656df} /* (15, 12, 14) {real, imag} */,
  {32'h41da4549, 32'hc22df25c} /* (15, 12, 13) {real, imag} */,
  {32'hc1fa1a78, 32'h4276138c} /* (15, 12, 12) {real, imag} */,
  {32'hc29db22f, 32'h3fbaeb60} /* (15, 12, 11) {real, imag} */,
  {32'hc1a91a94, 32'h4156c8c6} /* (15, 12, 10) {real, imag} */,
  {32'h4093c69e, 32'h41306f8f} /* (15, 12, 9) {real, imag} */,
  {32'h41d17b84, 32'h00000000} /* (15, 12, 8) {real, imag} */,
  {32'h4093c69e, 32'hc1306f8f} /* (15, 12, 7) {real, imag} */,
  {32'hc1a91a94, 32'hc156c8c6} /* (15, 12, 6) {real, imag} */,
  {32'hc29db22f, 32'hbfbaeb60} /* (15, 12, 5) {real, imag} */,
  {32'hc1fa1a78, 32'hc276138c} /* (15, 12, 4) {real, imag} */,
  {32'h41da4549, 32'h422df25c} /* (15, 12, 3) {real, imag} */,
  {32'h42b99074, 32'h430656df} /* (15, 12, 2) {real, imag} */,
  {32'h42b90f00, 32'h41fc4d48} /* (15, 12, 1) {real, imag} */,
  {32'hc00a96e0, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'h43146c86, 32'hc2ac4e63} /* (15, 11, 15) {real, imag} */,
  {32'h421bc3d4, 32'hc2eef395} /* (15, 11, 14) {real, imag} */,
  {32'hc20e8c3e, 32'h41aaf38c} /* (15, 11, 13) {real, imag} */,
  {32'hc25d8dbf, 32'h40860e32} /* (15, 11, 12) {real, imag} */,
  {32'hc19eef80, 32'hc2e59753} /* (15, 11, 11) {real, imag} */,
  {32'hc27ddb16, 32'hc1387630} /* (15, 11, 10) {real, imag} */,
  {32'hc1b5fb15, 32'h41980897} /* (15, 11, 9) {real, imag} */,
  {32'h422bcc0c, 32'h00000000} /* (15, 11, 8) {real, imag} */,
  {32'hc1b5fb15, 32'hc1980897} /* (15, 11, 7) {real, imag} */,
  {32'hc27ddb16, 32'h41387630} /* (15, 11, 6) {real, imag} */,
  {32'hc19eef80, 32'h42e59753} /* (15, 11, 5) {real, imag} */,
  {32'hc25d8dbf, 32'hc0860e32} /* (15, 11, 4) {real, imag} */,
  {32'hc20e8c3e, 32'hc1aaf38c} /* (15, 11, 3) {real, imag} */,
  {32'h421bc3d4, 32'h42eef395} /* (15, 11, 2) {real, imag} */,
  {32'h43146c86, 32'h42ac4e63} /* (15, 11, 1) {real, imag} */,
  {32'h425e8847, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h43214860, 32'hc2b36422} /* (15, 10, 15) {real, imag} */,
  {32'hc1c10c52, 32'hc100e374} /* (15, 10, 14) {real, imag} */,
  {32'h42e0d66e, 32'h419bae44} /* (15, 10, 13) {real, imag} */,
  {32'hc2f17fae, 32'hc2ade46f} /* (15, 10, 12) {real, imag} */,
  {32'hc237b5d4, 32'h42832d45} /* (15, 10, 11) {real, imag} */,
  {32'hc1806c67, 32'hc0869c5a} /* (15, 10, 10) {real, imag} */,
  {32'h4116df61, 32'hc0d36938} /* (15, 10, 9) {real, imag} */,
  {32'h4234515e, 32'h00000000} /* (15, 10, 8) {real, imag} */,
  {32'h4116df61, 32'h40d36938} /* (15, 10, 7) {real, imag} */,
  {32'hc1806c67, 32'h40869c5a} /* (15, 10, 6) {real, imag} */,
  {32'hc237b5d4, 32'hc2832d45} /* (15, 10, 5) {real, imag} */,
  {32'hc2f17fae, 32'h42ade46f} /* (15, 10, 4) {real, imag} */,
  {32'h42e0d66e, 32'hc19bae44} /* (15, 10, 3) {real, imag} */,
  {32'hc1c10c52, 32'h4100e374} /* (15, 10, 2) {real, imag} */,
  {32'h43214860, 32'h42b36422} /* (15, 10, 1) {real, imag} */,
  {32'h42da8954, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'h42faaa83, 32'hc25a4bb7} /* (15, 9, 15) {real, imag} */,
  {32'hc2192512, 32'h42e165b7} /* (15, 9, 14) {real, imag} */,
  {32'h41fe1a7a, 32'h42b274e1} /* (15, 9, 13) {real, imag} */,
  {32'h40c73d2c, 32'hc2900cff} /* (15, 9, 12) {real, imag} */,
  {32'h42ab3a9c, 32'h42861e5c} /* (15, 9, 11) {real, imag} */,
  {32'h41863864, 32'hc2dd6090} /* (15, 9, 10) {real, imag} */,
  {32'hc2435a47, 32'hc21a5ba4} /* (15, 9, 9) {real, imag} */,
  {32'hc200ab2b, 32'h00000000} /* (15, 9, 8) {real, imag} */,
  {32'hc2435a47, 32'h421a5ba4} /* (15, 9, 7) {real, imag} */,
  {32'h41863864, 32'h42dd6090} /* (15, 9, 6) {real, imag} */,
  {32'h42ab3a9c, 32'hc2861e5c} /* (15, 9, 5) {real, imag} */,
  {32'h40c73d2c, 32'h42900cff} /* (15, 9, 4) {real, imag} */,
  {32'h41fe1a7a, 32'hc2b274e1} /* (15, 9, 3) {real, imag} */,
  {32'hc2192512, 32'hc2e165b7} /* (15, 9, 2) {real, imag} */,
  {32'h42faaa83, 32'h425a4bb7} /* (15, 9, 1) {real, imag} */,
  {32'hc2af5be8, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'h42b847fb, 32'hc0ae1620} /* (15, 8, 15) {real, imag} */,
  {32'hc25f7026, 32'h43218d48} /* (15, 8, 14) {real, imag} */,
  {32'h429edb14, 32'hc1584a02} /* (15, 8, 13) {real, imag} */,
  {32'hc1bc6012, 32'hbd153300} /* (15, 8, 12) {real, imag} */,
  {32'h42b92ba5, 32'hc20a3be2} /* (15, 8, 11) {real, imag} */,
  {32'hc26b4072, 32'h40239d70} /* (15, 8, 10) {real, imag} */,
  {32'hc1a07be3, 32'hc2131344} /* (15, 8, 9) {real, imag} */,
  {32'hc2b63502, 32'h00000000} /* (15, 8, 8) {real, imag} */,
  {32'hc1a07be3, 32'h42131344} /* (15, 8, 7) {real, imag} */,
  {32'hc26b4072, 32'hc0239d70} /* (15, 8, 6) {real, imag} */,
  {32'h42b92ba5, 32'h420a3be2} /* (15, 8, 5) {real, imag} */,
  {32'hc1bc6012, 32'h3d153300} /* (15, 8, 4) {real, imag} */,
  {32'h429edb14, 32'h41584a02} /* (15, 8, 3) {real, imag} */,
  {32'hc25f7026, 32'hc3218d48} /* (15, 8, 2) {real, imag} */,
  {32'h42b847fb, 32'h40ae1620} /* (15, 8, 1) {real, imag} */,
  {32'hc2b5ea3b, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h41b14dc4, 32'h41dcd42e} /* (15, 7, 15) {real, imag} */,
  {32'h41ed4540, 32'hc27cfd42} /* (15, 7, 14) {real, imag} */,
  {32'h41806a9a, 32'hc293a7b3} /* (15, 7, 13) {real, imag} */,
  {32'hc1f4dbe5, 32'hc102c45a} /* (15, 7, 12) {real, imag} */,
  {32'h42804aa2, 32'h4125d83c} /* (15, 7, 11) {real, imag} */,
  {32'hc22cb666, 32'hbff32aa0} /* (15, 7, 10) {real, imag} */,
  {32'h41285ee4, 32'hbfa60640} /* (15, 7, 9) {real, imag} */,
  {32'h42252d2f, 32'h00000000} /* (15, 7, 8) {real, imag} */,
  {32'h41285ee4, 32'h3fa60640} /* (15, 7, 7) {real, imag} */,
  {32'hc22cb666, 32'h3ff32aa0} /* (15, 7, 6) {real, imag} */,
  {32'h42804aa2, 32'hc125d83c} /* (15, 7, 5) {real, imag} */,
  {32'hc1f4dbe5, 32'h4102c45a} /* (15, 7, 4) {real, imag} */,
  {32'h41806a9a, 32'h4293a7b3} /* (15, 7, 3) {real, imag} */,
  {32'h41ed4540, 32'h427cfd42} /* (15, 7, 2) {real, imag} */,
  {32'h41b14dc4, 32'hc1dcd42e} /* (15, 7, 1) {real, imag} */,
  {32'hc2a8073a, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'hc31ae212, 32'hc215ddf0} /* (15, 6, 15) {real, imag} */,
  {32'h425c71eb, 32'h3ff81100} /* (15, 6, 14) {real, imag} */,
  {32'h4208d579, 32'hc24e265e} /* (15, 6, 13) {real, imag} */,
  {32'h415e2724, 32'hc258738a} /* (15, 6, 12) {real, imag} */,
  {32'h4243a3d8, 32'hc100dcf8} /* (15, 6, 11) {real, imag} */,
  {32'hc185c73b, 32'h41d1ce62} /* (15, 6, 10) {real, imag} */,
  {32'h418f5172, 32'h422b5a2f} /* (15, 6, 9) {real, imag} */,
  {32'h42a66c87, 32'h00000000} /* (15, 6, 8) {real, imag} */,
  {32'h418f5172, 32'hc22b5a2f} /* (15, 6, 7) {real, imag} */,
  {32'hc185c73b, 32'hc1d1ce62} /* (15, 6, 6) {real, imag} */,
  {32'h4243a3d8, 32'h4100dcf8} /* (15, 6, 5) {real, imag} */,
  {32'h415e2724, 32'h4258738a} /* (15, 6, 4) {real, imag} */,
  {32'h4208d579, 32'h424e265e} /* (15, 6, 3) {real, imag} */,
  {32'h425c71eb, 32'hbff81100} /* (15, 6, 2) {real, imag} */,
  {32'hc31ae212, 32'h4215ddf0} /* (15, 6, 1) {real, imag} */,
  {32'hc1ff5720, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h4281198c, 32'hc3104a68} /* (15, 5, 15) {real, imag} */,
  {32'h428cb857, 32'h4277c2b6} /* (15, 5, 14) {real, imag} */,
  {32'hc1ed33cd, 32'h4270ae92} /* (15, 5, 13) {real, imag} */,
  {32'hc1b6eaba, 32'h41681e01} /* (15, 5, 12) {real, imag} */,
  {32'hc24766a0, 32'hc22270d2} /* (15, 5, 11) {real, imag} */,
  {32'hc2436a22, 32'hc15edea0} /* (15, 5, 10) {real, imag} */,
  {32'h41fd7661, 32'h4170988e} /* (15, 5, 9) {real, imag} */,
  {32'hc086ef2c, 32'h00000000} /* (15, 5, 8) {real, imag} */,
  {32'h41fd7661, 32'hc170988e} /* (15, 5, 7) {real, imag} */,
  {32'hc2436a22, 32'h415edea0} /* (15, 5, 6) {real, imag} */,
  {32'hc24766a0, 32'h422270d2} /* (15, 5, 5) {real, imag} */,
  {32'hc1b6eaba, 32'hc1681e01} /* (15, 5, 4) {real, imag} */,
  {32'hc1ed33cd, 32'hc270ae92} /* (15, 5, 3) {real, imag} */,
  {32'h428cb857, 32'hc277c2b6} /* (15, 5, 2) {real, imag} */,
  {32'h4281198c, 32'h43104a68} /* (15, 5, 1) {real, imag} */,
  {32'h4119c134, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'h4123cb90, 32'hc2b64da6} /* (15, 4, 15) {real, imag} */,
  {32'h406581c0, 32'h428ddadc} /* (15, 4, 14) {real, imag} */,
  {32'hc2460198, 32'hc0dd8290} /* (15, 4, 13) {real, imag} */,
  {32'hc1f1c48c, 32'hc2a022f8} /* (15, 4, 12) {real, imag} */,
  {32'hc0db2a30, 32'hc1bc7ab8} /* (15, 4, 11) {real, imag} */,
  {32'hc287e09a, 32'hc208235c} /* (15, 4, 10) {real, imag} */,
  {32'hc1e27de8, 32'hc1326273} /* (15, 4, 9) {real, imag} */,
  {32'h42d30913, 32'h00000000} /* (15, 4, 8) {real, imag} */,
  {32'hc1e27de8, 32'h41326273} /* (15, 4, 7) {real, imag} */,
  {32'hc287e09a, 32'h4208235c} /* (15, 4, 6) {real, imag} */,
  {32'hc0db2a30, 32'h41bc7ab8} /* (15, 4, 5) {real, imag} */,
  {32'hc1f1c48c, 32'h42a022f8} /* (15, 4, 4) {real, imag} */,
  {32'hc2460198, 32'h40dd8290} /* (15, 4, 3) {real, imag} */,
  {32'h406581c0, 32'hc28ddadc} /* (15, 4, 2) {real, imag} */,
  {32'h4123cb90, 32'h42b64da6} /* (15, 4, 1) {real, imag} */,
  {32'hc2bdf75b, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'hc1ceddee, 32'hc36c15f8} /* (15, 3, 15) {real, imag} */,
  {32'h41931f36, 32'h427d731a} /* (15, 3, 14) {real, imag} */,
  {32'h42272694, 32'hc1d4ad08} /* (15, 3, 13) {real, imag} */,
  {32'hc136e215, 32'hc07bb4f4} /* (15, 3, 12) {real, imag} */,
  {32'h42fbd187, 32'h41bfec37} /* (15, 3, 11) {real, imag} */,
  {32'h420a9e6e, 32'h425f0a1a} /* (15, 3, 10) {real, imag} */,
  {32'hc26e743e, 32'h42183547} /* (15, 3, 9) {real, imag} */,
  {32'h4313c3e2, 32'h00000000} /* (15, 3, 8) {real, imag} */,
  {32'hc26e743e, 32'hc2183547} /* (15, 3, 7) {real, imag} */,
  {32'h420a9e6e, 32'hc25f0a1a} /* (15, 3, 6) {real, imag} */,
  {32'h42fbd187, 32'hc1bfec37} /* (15, 3, 5) {real, imag} */,
  {32'hc136e215, 32'h407bb4f4} /* (15, 3, 4) {real, imag} */,
  {32'h42272694, 32'h41d4ad08} /* (15, 3, 3) {real, imag} */,
  {32'h41931f36, 32'hc27d731a} /* (15, 3, 2) {real, imag} */,
  {32'hc1ceddee, 32'h436c15f8} /* (15, 3, 1) {real, imag} */,
  {32'hc1e930da, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'hc0eb59b8, 32'hc3c19e55} /* (15, 2, 15) {real, imag} */,
  {32'h421c4264, 32'hc133cf06} /* (15, 2, 14) {real, imag} */,
  {32'hc2846543, 32'hc1a8cf5c} /* (15, 2, 13) {real, imag} */,
  {32'h42ed3cfb, 32'h424ae4ea} /* (15, 2, 12) {real, imag} */,
  {32'h426c46b8, 32'hc23c7e46} /* (15, 2, 11) {real, imag} */,
  {32'h42a9668d, 32'hc218122a} /* (15, 2, 10) {real, imag} */,
  {32'h41afac65, 32'h41e5dd10} /* (15, 2, 9) {real, imag} */,
  {32'hc1fb83c5, 32'h00000000} /* (15, 2, 8) {real, imag} */,
  {32'h41afac65, 32'hc1e5dd10} /* (15, 2, 7) {real, imag} */,
  {32'h42a9668d, 32'h4218122a} /* (15, 2, 6) {real, imag} */,
  {32'h426c46b8, 32'h423c7e46} /* (15, 2, 5) {real, imag} */,
  {32'h42ed3cfb, 32'hc24ae4ea} /* (15, 2, 4) {real, imag} */,
  {32'hc2846543, 32'h41a8cf5c} /* (15, 2, 3) {real, imag} */,
  {32'h421c4264, 32'h4133cf06} /* (15, 2, 2) {real, imag} */,
  {32'hc0eb59b8, 32'h43c19e55} /* (15, 2, 1) {real, imag} */,
  {32'hc339c00d, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'hc1f38a84, 32'hc3b7e28f} /* (15, 1, 15) {real, imag} */,
  {32'h42594286, 32'h431caa6a} /* (15, 1, 14) {real, imag} */,
  {32'hc29b0580, 32'hc1dcfafe} /* (15, 1, 13) {real, imag} */,
  {32'h421afdc0, 32'hc256b69a} /* (15, 1, 12) {real, imag} */,
  {32'hc1cddad7, 32'hc151d633} /* (15, 1, 11) {real, imag} */,
  {32'hc22810c6, 32'hc1fbe9c6} /* (15, 1, 10) {real, imag} */,
  {32'hc1a28faa, 32'hc232f6c5} /* (15, 1, 9) {real, imag} */,
  {32'h41ace45a, 32'h00000000} /* (15, 1, 8) {real, imag} */,
  {32'hc1a28faa, 32'h4232f6c5} /* (15, 1, 7) {real, imag} */,
  {32'hc22810c6, 32'h41fbe9c6} /* (15, 1, 6) {real, imag} */,
  {32'hc1cddad7, 32'h4151d633} /* (15, 1, 5) {real, imag} */,
  {32'h421afdc0, 32'h4256b69a} /* (15, 1, 4) {real, imag} */,
  {32'hc29b0580, 32'h41dcfafe} /* (15, 1, 3) {real, imag} */,
  {32'h42594286, 32'hc31caa6a} /* (15, 1, 2) {real, imag} */,
  {32'hc1f38a84, 32'h43b7e28f} /* (15, 1, 1) {real, imag} */,
  {32'hc3a76af4, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'h413991f8, 32'hc32c5705} /* (15, 0, 15) {real, imag} */,
  {32'h41af1d0c, 32'hbf4b5580} /* (15, 0, 14) {real, imag} */,
  {32'h414eb7e0, 32'hc172907e} /* (15, 0, 13) {real, imag} */,
  {32'hc17f1654, 32'hc1d43aa8} /* (15, 0, 12) {real, imag} */,
  {32'hc12e84d8, 32'hc1a57b52} /* (15, 0, 11) {real, imag} */,
  {32'hc1c34de1, 32'h4265da99} /* (15, 0, 10) {real, imag} */,
  {32'h41312058, 32'hc0939bfc} /* (15, 0, 9) {real, imag} */,
  {32'h401ef9d0, 32'h00000000} /* (15, 0, 8) {real, imag} */,
  {32'h41312058, 32'h40939bfc} /* (15, 0, 7) {real, imag} */,
  {32'hc1c34de1, 32'hc265da99} /* (15, 0, 6) {real, imag} */,
  {32'hc12e84d8, 32'h41a57b52} /* (15, 0, 5) {real, imag} */,
  {32'hc17f1654, 32'h41d43aa8} /* (15, 0, 4) {real, imag} */,
  {32'h414eb7e0, 32'h4172907e} /* (15, 0, 3) {real, imag} */,
  {32'h41af1d0c, 32'h3f4b5580} /* (15, 0, 2) {real, imag} */,
  {32'h413991f8, 32'h432c5705} /* (15, 0, 1) {real, imag} */,
  {32'hc380e323, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h420af4b0, 32'hc2a8ac20} /* (14, 15, 15) {real, imag} */,
  {32'hc2b63534, 32'hc3109a97} /* (14, 15, 14) {real, imag} */,
  {32'h429f7608, 32'h41571928} /* (14, 15, 13) {real, imag} */,
  {32'h404705b0, 32'hc26d6940} /* (14, 15, 12) {real, imag} */,
  {32'hc1ea4b6a, 32'hc2e5ea5f} /* (14, 15, 11) {real, imag} */,
  {32'h42039306, 32'hc2c92436} /* (14, 15, 10) {real, imag} */,
  {32'hc0625db0, 32'hc1f98e10} /* (14, 15, 9) {real, imag} */,
  {32'hc18029ca, 32'h00000000} /* (14, 15, 8) {real, imag} */,
  {32'hc0625db0, 32'h41f98e10} /* (14, 15, 7) {real, imag} */,
  {32'h42039306, 32'h42c92436} /* (14, 15, 6) {real, imag} */,
  {32'hc1ea4b6a, 32'h42e5ea5f} /* (14, 15, 5) {real, imag} */,
  {32'h404705b0, 32'h426d6940} /* (14, 15, 4) {real, imag} */,
  {32'h429f7608, 32'hc1571928} /* (14, 15, 3) {real, imag} */,
  {32'hc2b63534, 32'h43109a97} /* (14, 15, 2) {real, imag} */,
  {32'h420af4b0, 32'h42a8ac20} /* (14, 15, 1) {real, imag} */,
  {32'hc3a0aada, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'hc2092740, 32'hc2dbbf2a} /* (14, 14, 15) {real, imag} */,
  {32'hc1739f72, 32'hc20634ba} /* (14, 14, 14) {real, imag} */,
  {32'h42c2b1c2, 32'hc0343b30} /* (14, 14, 13) {real, imag} */,
  {32'h40958380, 32'hc2f847c1} /* (14, 14, 12) {real, imag} */,
  {32'h42824968, 32'h42467685} /* (14, 14, 11) {real, imag} */,
  {32'h41c4911b, 32'hc2bcebb9} /* (14, 14, 10) {real, imag} */,
  {32'hc1312724, 32'hc243bc18} /* (14, 14, 9) {real, imag} */,
  {32'hc220f9b0, 32'h00000000} /* (14, 14, 8) {real, imag} */,
  {32'hc1312724, 32'h4243bc18} /* (14, 14, 7) {real, imag} */,
  {32'h41c4911b, 32'h42bcebb9} /* (14, 14, 6) {real, imag} */,
  {32'h42824968, 32'hc2467685} /* (14, 14, 5) {real, imag} */,
  {32'h40958380, 32'h42f847c1} /* (14, 14, 4) {real, imag} */,
  {32'h42c2b1c2, 32'h40343b30} /* (14, 14, 3) {real, imag} */,
  {32'hc1739f72, 32'h420634ba} /* (14, 14, 2) {real, imag} */,
  {32'hc2092740, 32'h42dbbf2a} /* (14, 14, 1) {real, imag} */,
  {32'hc38f5c8c, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'h428828d4, 32'h41143cf0} /* (14, 13, 15) {real, imag} */,
  {32'h431f7468, 32'hc2b4a02a} /* (14, 13, 14) {real, imag} */,
  {32'h42a5cfd2, 32'hc321c8ed} /* (14, 13, 13) {real, imag} */,
  {32'hc1e87748, 32'h422e1ad4} /* (14, 13, 12) {real, imag} */,
  {32'h4248c145, 32'h42233a3c} /* (14, 13, 11) {real, imag} */,
  {32'h4132eb90, 32'h42d0049c} /* (14, 13, 10) {real, imag} */,
  {32'hc20058b2, 32'hc286748b} /* (14, 13, 9) {real, imag} */,
  {32'h423d9e78, 32'h00000000} /* (14, 13, 8) {real, imag} */,
  {32'hc20058b2, 32'h4286748b} /* (14, 13, 7) {real, imag} */,
  {32'h4132eb90, 32'hc2d0049c} /* (14, 13, 6) {real, imag} */,
  {32'h4248c145, 32'hc2233a3c} /* (14, 13, 5) {real, imag} */,
  {32'hc1e87748, 32'hc22e1ad4} /* (14, 13, 4) {real, imag} */,
  {32'h42a5cfd2, 32'h4321c8ed} /* (14, 13, 3) {real, imag} */,
  {32'h431f7468, 32'h42b4a02a} /* (14, 13, 2) {real, imag} */,
  {32'h428828d4, 32'hc1143cf0} /* (14, 13, 1) {real, imag} */,
  {32'hc2daac51, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'h435e8ecd, 32'hc2526614} /* (14, 12, 15) {real, imag} */,
  {32'h42f7ed02, 32'hc25a22cc} /* (14, 12, 14) {real, imag} */,
  {32'h4188bf5d, 32'hc1682ee4} /* (14, 12, 13) {real, imag} */,
  {32'hc1af1d20, 32'h42d5eaef} /* (14, 12, 12) {real, imag} */,
  {32'h42a730d6, 32'h4176b0d8} /* (14, 12, 11) {real, imag} */,
  {32'hc22e9c2b, 32'hc25e8514} /* (14, 12, 10) {real, imag} */,
  {32'hc2ad6542, 32'h430c40a6} /* (14, 12, 9) {real, imag} */,
  {32'h4170b478, 32'h00000000} /* (14, 12, 8) {real, imag} */,
  {32'hc2ad6542, 32'hc30c40a6} /* (14, 12, 7) {real, imag} */,
  {32'hc22e9c2b, 32'h425e8514} /* (14, 12, 6) {real, imag} */,
  {32'h42a730d6, 32'hc176b0d8} /* (14, 12, 5) {real, imag} */,
  {32'hc1af1d20, 32'hc2d5eaef} /* (14, 12, 4) {real, imag} */,
  {32'h4188bf5d, 32'h41682ee4} /* (14, 12, 3) {real, imag} */,
  {32'h42f7ed02, 32'h425a22cc} /* (14, 12, 2) {real, imag} */,
  {32'h435e8ecd, 32'h42526614} /* (14, 12, 1) {real, imag} */,
  {32'hc386aa56, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'h42ef56e0, 32'hc285c2de} /* (14, 11, 15) {real, imag} */,
  {32'hc28e7e09, 32'hc24e66c7} /* (14, 11, 14) {real, imag} */,
  {32'hc2d9d5d0, 32'hc257a427} /* (14, 11, 13) {real, imag} */,
  {32'h430dbd18, 32'hc194a175} /* (14, 11, 12) {real, imag} */,
  {32'hc2d73ca4, 32'h4269d710} /* (14, 11, 11) {real, imag} */,
  {32'hc1d2a4b6, 32'h42cfce12} /* (14, 11, 10) {real, imag} */,
  {32'hc18047bb, 32'hc28d5909} /* (14, 11, 9) {real, imag} */,
  {32'hc1ddbcfe, 32'h00000000} /* (14, 11, 8) {real, imag} */,
  {32'hc18047bb, 32'h428d5909} /* (14, 11, 7) {real, imag} */,
  {32'hc1d2a4b6, 32'hc2cfce12} /* (14, 11, 6) {real, imag} */,
  {32'hc2d73ca4, 32'hc269d710} /* (14, 11, 5) {real, imag} */,
  {32'h430dbd18, 32'h4194a175} /* (14, 11, 4) {real, imag} */,
  {32'hc2d9d5d0, 32'h4257a427} /* (14, 11, 3) {real, imag} */,
  {32'hc28e7e09, 32'h424e66c7} /* (14, 11, 2) {real, imag} */,
  {32'h42ef56e0, 32'h4285c2de} /* (14, 11, 1) {real, imag} */,
  {32'h42e7691a, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h42d15310, 32'hc1754d50} /* (14, 10, 15) {real, imag} */,
  {32'h4214658a, 32'hc2b6c534} /* (14, 10, 14) {real, imag} */,
  {32'hc1bdfc88, 32'hc25d1a66} /* (14, 10, 13) {real, imag} */,
  {32'h4265d96c, 32'hc2596efc} /* (14, 10, 12) {real, imag} */,
  {32'hc191e21a, 32'h4332248c} /* (14, 10, 11) {real, imag} */,
  {32'h41355f2c, 32'h42cecb2b} /* (14, 10, 10) {real, imag} */,
  {32'h422063f4, 32'h41df3fd9} /* (14, 10, 9) {real, imag} */,
  {32'h40c16a38, 32'h00000000} /* (14, 10, 8) {real, imag} */,
  {32'h422063f4, 32'hc1df3fd9} /* (14, 10, 7) {real, imag} */,
  {32'h41355f2c, 32'hc2cecb2b} /* (14, 10, 6) {real, imag} */,
  {32'hc191e21a, 32'hc332248c} /* (14, 10, 5) {real, imag} */,
  {32'h4265d96c, 32'h42596efc} /* (14, 10, 4) {real, imag} */,
  {32'hc1bdfc88, 32'h425d1a66} /* (14, 10, 3) {real, imag} */,
  {32'h4214658a, 32'h42b6c534} /* (14, 10, 2) {real, imag} */,
  {32'h42d15310, 32'h41754d50} /* (14, 10, 1) {real, imag} */,
  {32'h42e507d0, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'h42d4fd23, 32'hc3360fc1} /* (14, 9, 15) {real, imag} */,
  {32'hc2f96df0, 32'h42957969} /* (14, 9, 14) {real, imag} */,
  {32'h4349e346, 32'h42b97e1e} /* (14, 9, 13) {real, imag} */,
  {32'h430ab738, 32'hc3390d7a} /* (14, 9, 12) {real, imag} */,
  {32'hc1d6c114, 32'h41c3370b} /* (14, 9, 11) {real, imag} */,
  {32'h432edd5f, 32'hc2a59c28} /* (14, 9, 10) {real, imag} */,
  {32'h41d15e74, 32'h431fc997} /* (14, 9, 9) {real, imag} */,
  {32'h42d40a6c, 32'h00000000} /* (14, 9, 8) {real, imag} */,
  {32'h41d15e74, 32'hc31fc997} /* (14, 9, 7) {real, imag} */,
  {32'h432edd5f, 32'h42a59c28} /* (14, 9, 6) {real, imag} */,
  {32'hc1d6c114, 32'hc1c3370b} /* (14, 9, 5) {real, imag} */,
  {32'h430ab738, 32'h43390d7a} /* (14, 9, 4) {real, imag} */,
  {32'h4349e346, 32'hc2b97e1e} /* (14, 9, 3) {real, imag} */,
  {32'hc2f96df0, 32'hc2957969} /* (14, 9, 2) {real, imag} */,
  {32'h42d4fd23, 32'h43360fc1} /* (14, 9, 1) {real, imag} */,
  {32'hc19d39e4, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'hc22f3154, 32'hc08b8460} /* (14, 8, 15) {real, imag} */,
  {32'hc2680f8f, 32'h43627d84} /* (14, 8, 14) {real, imag} */,
  {32'h42554a8a, 32'hc2bdf9fa} /* (14, 8, 13) {real, imag} */,
  {32'h4293ccda, 32'hc1823ecf} /* (14, 8, 12) {real, imag} */,
  {32'hc1570ac0, 32'h4307e8b4} /* (14, 8, 11) {real, imag} */,
  {32'h4285e96e, 32'hc2d5e48c} /* (14, 8, 10) {real, imag} */,
  {32'hc2a4a06e, 32'hc274d0f7} /* (14, 8, 9) {real, imag} */,
  {32'hc0cf7e50, 32'h00000000} /* (14, 8, 8) {real, imag} */,
  {32'hc2a4a06e, 32'h4274d0f7} /* (14, 8, 7) {real, imag} */,
  {32'h4285e96e, 32'h42d5e48c} /* (14, 8, 6) {real, imag} */,
  {32'hc1570ac0, 32'hc307e8b4} /* (14, 8, 5) {real, imag} */,
  {32'h4293ccda, 32'h41823ecf} /* (14, 8, 4) {real, imag} */,
  {32'h42554a8a, 32'h42bdf9fa} /* (14, 8, 3) {real, imag} */,
  {32'hc2680f8f, 32'hc3627d84} /* (14, 8, 2) {real, imag} */,
  {32'hc22f3154, 32'h408b8460} /* (14, 8, 1) {real, imag} */,
  {32'h4116b648, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'hc34db59e, 32'h41ba4578} /* (14, 7, 15) {real, imag} */,
  {32'h4318e4b8, 32'h43033aec} /* (14, 7, 14) {real, imag} */,
  {32'h4322f946, 32'hc30dabd1} /* (14, 7, 13) {real, imag} */,
  {32'hc2cc0011, 32'h422ed788} /* (14, 7, 12) {real, imag} */,
  {32'hc23f3c86, 32'h3fe8c450} /* (14, 7, 11) {real, imag} */,
  {32'h421d07e0, 32'hc19da28a} /* (14, 7, 10) {real, imag} */,
  {32'hc1b0097c, 32'hc28f97be} /* (14, 7, 9) {real, imag} */,
  {32'hc28793ce, 32'h00000000} /* (14, 7, 8) {real, imag} */,
  {32'hc1b0097c, 32'h428f97be} /* (14, 7, 7) {real, imag} */,
  {32'h421d07e0, 32'h419da28a} /* (14, 7, 6) {real, imag} */,
  {32'hc23f3c86, 32'hbfe8c450} /* (14, 7, 5) {real, imag} */,
  {32'hc2cc0011, 32'hc22ed788} /* (14, 7, 4) {real, imag} */,
  {32'h4322f946, 32'h430dabd1} /* (14, 7, 3) {real, imag} */,
  {32'h4318e4b8, 32'hc3033aec} /* (14, 7, 2) {real, imag} */,
  {32'hc34db59e, 32'hc1ba4578} /* (14, 7, 1) {real, imag} */,
  {32'hc2c0939b, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'hc324e724, 32'hc32a9237} /* (14, 6, 15) {real, imag} */,
  {32'h4285517b, 32'h430f182c} /* (14, 6, 14) {real, imag} */,
  {32'h421ab283, 32'hc2052a3c} /* (14, 6, 13) {real, imag} */,
  {32'h4287aff6, 32'hc2e0c176} /* (14, 6, 12) {real, imag} */,
  {32'h4276bbe5, 32'hc1adf634} /* (14, 6, 11) {real, imag} */,
  {32'hc0e182f8, 32'h434c9406} /* (14, 6, 10) {real, imag} */,
  {32'h42a18d01, 32'hc100e09e} /* (14, 6, 9) {real, imag} */,
  {32'hc2c5dba2, 32'h00000000} /* (14, 6, 8) {real, imag} */,
  {32'h42a18d01, 32'h4100e09e} /* (14, 6, 7) {real, imag} */,
  {32'hc0e182f8, 32'hc34c9406} /* (14, 6, 6) {real, imag} */,
  {32'h4276bbe5, 32'h41adf634} /* (14, 6, 5) {real, imag} */,
  {32'h4287aff6, 32'h42e0c176} /* (14, 6, 4) {real, imag} */,
  {32'h421ab283, 32'h42052a3c} /* (14, 6, 3) {real, imag} */,
  {32'h4285517b, 32'hc30f182c} /* (14, 6, 2) {real, imag} */,
  {32'hc324e724, 32'h432a9237} /* (14, 6, 1) {real, imag} */,
  {32'h434b96e4, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h42876b40, 32'hc29674d6} /* (14, 5, 15) {real, imag} */,
  {32'h43120fc0, 32'h4324109c} /* (14, 5, 14) {real, imag} */,
  {32'hc221cb90, 32'hc28ed8b6} /* (14, 5, 13) {real, imag} */,
  {32'hc2ee09df, 32'hc23b7704} /* (14, 5, 12) {real, imag} */,
  {32'hc1f7cb80, 32'h4300ef74} /* (14, 5, 11) {real, imag} */,
  {32'hc22b522d, 32'h4323e735} /* (14, 5, 10) {real, imag} */,
  {32'h412ddbb6, 32'h422a1ebe} /* (14, 5, 9) {real, imag} */,
  {32'hc237ae6f, 32'h00000000} /* (14, 5, 8) {real, imag} */,
  {32'h412ddbb6, 32'hc22a1ebe} /* (14, 5, 7) {real, imag} */,
  {32'hc22b522d, 32'hc323e735} /* (14, 5, 6) {real, imag} */,
  {32'hc1f7cb80, 32'hc300ef74} /* (14, 5, 5) {real, imag} */,
  {32'hc2ee09df, 32'h423b7704} /* (14, 5, 4) {real, imag} */,
  {32'hc221cb90, 32'h428ed8b6} /* (14, 5, 3) {real, imag} */,
  {32'h43120fc0, 32'hc324109c} /* (14, 5, 2) {real, imag} */,
  {32'h42876b40, 32'h429674d6} /* (14, 5, 1) {real, imag} */,
  {32'h42cf5238, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'hc1cfcb28, 32'hc3333beb} /* (14, 4, 15) {real, imag} */,
  {32'h431609b9, 32'h42e8f6ea} /* (14, 4, 14) {real, imag} */,
  {32'hc1afc60b, 32'h41b7273a} /* (14, 4, 13) {real, imag} */,
  {32'h42cbc9cc, 32'hc2bf14a9} /* (14, 4, 12) {real, imag} */,
  {32'hc17c739c, 32'h42bcb9d2} /* (14, 4, 11) {real, imag} */,
  {32'hc2afcb00, 32'h42ab661e} /* (14, 4, 10) {real, imag} */,
  {32'hc2727a54, 32'h4010c860} /* (14, 4, 9) {real, imag} */,
  {32'h42e1dd11, 32'h00000000} /* (14, 4, 8) {real, imag} */,
  {32'hc2727a54, 32'hc010c860} /* (14, 4, 7) {real, imag} */,
  {32'hc2afcb00, 32'hc2ab661e} /* (14, 4, 6) {real, imag} */,
  {32'hc17c739c, 32'hc2bcb9d2} /* (14, 4, 5) {real, imag} */,
  {32'h42cbc9cc, 32'h42bf14a9} /* (14, 4, 4) {real, imag} */,
  {32'hc1afc60b, 32'hc1b7273a} /* (14, 4, 3) {real, imag} */,
  {32'h431609b9, 32'hc2e8f6ea} /* (14, 4, 2) {real, imag} */,
  {32'hc1cfcb28, 32'h43333beb} /* (14, 4, 1) {real, imag} */,
  {32'hc1cce0c0, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'h4348c7a6, 32'hc3c6aaea} /* (14, 3, 15) {real, imag} */,
  {32'h40d796b0, 32'h42c6c9fa} /* (14, 3, 14) {real, imag} */,
  {32'h40a22880, 32'h4300bca7} /* (14, 3, 13) {real, imag} */,
  {32'h419d37f0, 32'hc1109cba} /* (14, 3, 12) {real, imag} */,
  {32'h4293a82e, 32'hc3067ba9} /* (14, 3, 11) {real, imag} */,
  {32'h43397fb7, 32'h42eca908} /* (14, 3, 10) {real, imag} */,
  {32'h42e999a3, 32'h42833317} /* (14, 3, 9) {real, imag} */,
  {32'h406814a0, 32'h00000000} /* (14, 3, 8) {real, imag} */,
  {32'h42e999a3, 32'hc2833317} /* (14, 3, 7) {real, imag} */,
  {32'h43397fb7, 32'hc2eca908} /* (14, 3, 6) {real, imag} */,
  {32'h4293a82e, 32'h43067ba9} /* (14, 3, 5) {real, imag} */,
  {32'h419d37f0, 32'h41109cba} /* (14, 3, 4) {real, imag} */,
  {32'h40a22880, 32'hc300bca7} /* (14, 3, 3) {real, imag} */,
  {32'h40d796b0, 32'hc2c6c9fa} /* (14, 3, 2) {real, imag} */,
  {32'h4348c7a6, 32'h43c6aaea} /* (14, 3, 1) {real, imag} */,
  {32'h42a5712f, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h4339e0e8, 32'hc413b7e7} /* (14, 2, 15) {real, imag} */,
  {32'h420b5228, 32'h4187f34b} /* (14, 2, 14) {real, imag} */,
  {32'hc2a70432, 32'hc243be83} /* (14, 2, 13) {real, imag} */,
  {32'hc291eff6, 32'hc27fc526} /* (14, 2, 12) {real, imag} */,
  {32'h4318e31c, 32'hbe481b00} /* (14, 2, 11) {real, imag} */,
  {32'hc29d957a, 32'hc2cba631} /* (14, 2, 10) {real, imag} */,
  {32'hc2dc5c72, 32'h42acf80e} /* (14, 2, 9) {real, imag} */,
  {32'h436133c0, 32'h00000000} /* (14, 2, 8) {real, imag} */,
  {32'hc2dc5c72, 32'hc2acf80e} /* (14, 2, 7) {real, imag} */,
  {32'hc29d957a, 32'h42cba631} /* (14, 2, 6) {real, imag} */,
  {32'h4318e31c, 32'h3e481b00} /* (14, 2, 5) {real, imag} */,
  {32'hc291eff6, 32'h427fc526} /* (14, 2, 4) {real, imag} */,
  {32'hc2a70432, 32'h4243be83} /* (14, 2, 3) {real, imag} */,
  {32'h420b5228, 32'hc187f34b} /* (14, 2, 2) {real, imag} */,
  {32'h4339e0e8, 32'h4413b7e7} /* (14, 2, 1) {real, imag} */,
  {32'hc316421c, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h423bf260, 32'hc4071f0c} /* (14, 1, 15) {real, imag} */,
  {32'h42b4c2da, 32'h42e82cfa} /* (14, 1, 14) {real, imag} */,
  {32'hc36d447c, 32'hc3074f32} /* (14, 1, 13) {real, imag} */,
  {32'h4206a83d, 32'h423e9548} /* (14, 1, 12) {real, imag} */,
  {32'h42125b27, 32'hc332c228} /* (14, 1, 11) {real, imag} */,
  {32'hc25c0b3a, 32'hc1335414} /* (14, 1, 10) {real, imag} */,
  {32'h42655e53, 32'h40e1d690} /* (14, 1, 9) {real, imag} */,
  {32'h425e9cb7, 32'h00000000} /* (14, 1, 8) {real, imag} */,
  {32'h42655e53, 32'hc0e1d690} /* (14, 1, 7) {real, imag} */,
  {32'hc25c0b3a, 32'h41335414} /* (14, 1, 6) {real, imag} */,
  {32'h42125b27, 32'h4332c228} /* (14, 1, 5) {real, imag} */,
  {32'h4206a83d, 32'hc23e9548} /* (14, 1, 4) {real, imag} */,
  {32'hc36d447c, 32'h43074f32} /* (14, 1, 3) {real, imag} */,
  {32'h42b4c2da, 32'hc2e82cfa} /* (14, 1, 2) {real, imag} */,
  {32'h423bf260, 32'h44071f0c} /* (14, 1, 1) {real, imag} */,
  {32'hc3c4214e, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h431fd261, 32'hc373c671} /* (14, 0, 15) {real, imag} */,
  {32'hc22648f3, 32'h41e117f0} /* (14, 0, 14) {real, imag} */,
  {32'hc2f2da5f, 32'hbfc4e100} /* (14, 0, 13) {real, imag} */,
  {32'h4307bd79, 32'h42251bc8} /* (14, 0, 12) {real, imag} */,
  {32'hc2de317f, 32'hc259153b} /* (14, 0, 11) {real, imag} */,
  {32'h42827574, 32'h42789460} /* (14, 0, 10) {real, imag} */,
  {32'hc133e2d0, 32'hc1b7234a} /* (14, 0, 9) {real, imag} */,
  {32'h423e4556, 32'h00000000} /* (14, 0, 8) {real, imag} */,
  {32'hc133e2d0, 32'h41b7234a} /* (14, 0, 7) {real, imag} */,
  {32'h42827574, 32'hc2789460} /* (14, 0, 6) {real, imag} */,
  {32'hc2de317f, 32'h4259153b} /* (14, 0, 5) {real, imag} */,
  {32'h4307bd79, 32'hc2251bc8} /* (14, 0, 4) {real, imag} */,
  {32'hc2f2da5f, 32'h3fc4e100} /* (14, 0, 3) {real, imag} */,
  {32'hc22648f3, 32'hc1e117f0} /* (14, 0, 2) {real, imag} */,
  {32'h431fd261, 32'h4373c671} /* (14, 0, 1) {real, imag} */,
  {32'hc338f782, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h4385c56a, 32'h42793c44} /* (13, 15, 15) {real, imag} */,
  {32'h4238d3cc, 32'hc1e8883e} /* (13, 15, 14) {real, imag} */,
  {32'h421951da, 32'h42bb32e2} /* (13, 15, 13) {real, imag} */,
  {32'h42baf190, 32'hc290a1cf} /* (13, 15, 12) {real, imag} */,
  {32'hc1d568ac, 32'h4281b99e} /* (13, 15, 11) {real, imag} */,
  {32'h4202836f, 32'h41debe57} /* (13, 15, 10) {real, imag} */,
  {32'h42e74d68, 32'hc103ec7c} /* (13, 15, 9) {real, imag} */,
  {32'hc2055c7e, 32'h00000000} /* (13, 15, 8) {real, imag} */,
  {32'h42e74d68, 32'h4103ec7c} /* (13, 15, 7) {real, imag} */,
  {32'h4202836f, 32'hc1debe57} /* (13, 15, 6) {real, imag} */,
  {32'hc1d568ac, 32'hc281b99e} /* (13, 15, 5) {real, imag} */,
  {32'h42baf190, 32'h4290a1cf} /* (13, 15, 4) {real, imag} */,
  {32'h421951da, 32'hc2bb32e2} /* (13, 15, 3) {real, imag} */,
  {32'h4238d3cc, 32'h41e8883e} /* (13, 15, 2) {real, imag} */,
  {32'h4385c56a, 32'hc2793c44} /* (13, 15, 1) {real, imag} */,
  {32'hc28f782a, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'h43096bca, 32'h420b5cba} /* (13, 14, 15) {real, imag} */,
  {32'h427e8923, 32'hc3560d66} /* (13, 14, 14) {real, imag} */,
  {32'h42e419be, 32'h425784a8} /* (13, 14, 13) {real, imag} */,
  {32'h43135744, 32'hc3185ab7} /* (13, 14, 12) {real, imag} */,
  {32'h42148f32, 32'h4187c952} /* (13, 14, 11) {real, imag} */,
  {32'h41d1993a, 32'h425f3931} /* (13, 14, 10) {real, imag} */,
  {32'h4287ed1b, 32'h41540170} /* (13, 14, 9) {real, imag} */,
  {32'hc20f99be, 32'h00000000} /* (13, 14, 8) {real, imag} */,
  {32'h4287ed1b, 32'hc1540170} /* (13, 14, 7) {real, imag} */,
  {32'h41d1993a, 32'hc25f3931} /* (13, 14, 6) {real, imag} */,
  {32'h42148f32, 32'hc187c952} /* (13, 14, 5) {real, imag} */,
  {32'h43135744, 32'h43185ab7} /* (13, 14, 4) {real, imag} */,
  {32'h42e419be, 32'hc25784a8} /* (13, 14, 3) {real, imag} */,
  {32'h427e8923, 32'h43560d66} /* (13, 14, 2) {real, imag} */,
  {32'h43096bca, 32'hc20b5cba} /* (13, 14, 1) {real, imag} */,
  {32'hc3a9d3f2, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'h41258b10, 32'h40990ae0} /* (13, 13, 15) {real, imag} */,
  {32'h42073ff6, 32'hc1ba8bb9} /* (13, 13, 14) {real, imag} */,
  {32'h42863481, 32'hc204cdbe} /* (13, 13, 13) {real, imag} */,
  {32'hc2937082, 32'hc245825a} /* (13, 13, 12) {real, imag} */,
  {32'h42146d3d, 32'hc318e67e} /* (13, 13, 11) {real, imag} */,
  {32'hc1b41f80, 32'h41ffd494} /* (13, 13, 10) {real, imag} */,
  {32'hbf929504, 32'hc30b130e} /* (13, 13, 9) {real, imag} */,
  {32'h42513885, 32'h00000000} /* (13, 13, 8) {real, imag} */,
  {32'hbf929504, 32'h430b130e} /* (13, 13, 7) {real, imag} */,
  {32'hc1b41f80, 32'hc1ffd494} /* (13, 13, 6) {real, imag} */,
  {32'h42146d3d, 32'h4318e67e} /* (13, 13, 5) {real, imag} */,
  {32'hc2937082, 32'h4245825a} /* (13, 13, 4) {real, imag} */,
  {32'h42863481, 32'h4204cdbe} /* (13, 13, 3) {real, imag} */,
  {32'h42073ff6, 32'h41ba8bb9} /* (13, 13, 2) {real, imag} */,
  {32'h41258b10, 32'hc0990ae0} /* (13, 13, 1) {real, imag} */,
  {32'hc37e4b7d, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'hc24317ae, 32'hc3276da8} /* (13, 12, 15) {real, imag} */,
  {32'hbf252480, 32'h41b0cfba} /* (13, 12, 14) {real, imag} */,
  {32'h4111b408, 32'hc322a3c0} /* (13, 12, 13) {real, imag} */,
  {32'h42d18a36, 32'h430b70e8} /* (13, 12, 12) {real, imag} */,
  {32'hc0411900, 32'hc2ac0109} /* (13, 12, 11) {real, imag} */,
  {32'hc2a7befb, 32'h42685c0c} /* (13, 12, 10) {real, imag} */,
  {32'hc298049e, 32'h4125256c} /* (13, 12, 9) {real, imag} */,
  {32'hc309a56c, 32'h00000000} /* (13, 12, 8) {real, imag} */,
  {32'hc298049e, 32'hc125256c} /* (13, 12, 7) {real, imag} */,
  {32'hc2a7befb, 32'hc2685c0c} /* (13, 12, 6) {real, imag} */,
  {32'hc0411900, 32'h42ac0109} /* (13, 12, 5) {real, imag} */,
  {32'h42d18a36, 32'hc30b70e8} /* (13, 12, 4) {real, imag} */,
  {32'h4111b408, 32'h4322a3c0} /* (13, 12, 3) {real, imag} */,
  {32'hbf252480, 32'hc1b0cfba} /* (13, 12, 2) {real, imag} */,
  {32'hc24317ae, 32'h43276da8} /* (13, 12, 1) {real, imag} */,
  {32'hc1a33fb8, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'hc21dbd64, 32'hc361814b} /* (13, 11, 15) {real, imag} */,
  {32'h425e97b6, 32'h427c2bd4} /* (13, 11, 14) {real, imag} */,
  {32'hc26fcf48, 32'hc2c2f264} /* (13, 11, 13) {real, imag} */,
  {32'h4345510e, 32'hbfe08bc0} /* (13, 11, 12) {real, imag} */,
  {32'hc2ab3b1e, 32'h42e09700} /* (13, 11, 11) {real, imag} */,
  {32'h422d11bc, 32'h41e5f72d} /* (13, 11, 10) {real, imag} */,
  {32'hc1de28e4, 32'hc1cdf20a} /* (13, 11, 9) {real, imag} */,
  {32'hc2bb01f8, 32'h00000000} /* (13, 11, 8) {real, imag} */,
  {32'hc1de28e4, 32'h41cdf20a} /* (13, 11, 7) {real, imag} */,
  {32'h422d11bc, 32'hc1e5f72d} /* (13, 11, 6) {real, imag} */,
  {32'hc2ab3b1e, 32'hc2e09700} /* (13, 11, 5) {real, imag} */,
  {32'h4345510e, 32'h3fe08bc0} /* (13, 11, 4) {real, imag} */,
  {32'hc26fcf48, 32'h42c2f264} /* (13, 11, 3) {real, imag} */,
  {32'h425e97b6, 32'hc27c2bd4} /* (13, 11, 2) {real, imag} */,
  {32'hc21dbd64, 32'h4361814b} /* (13, 11, 1) {real, imag} */,
  {32'hc28202a8, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'h42087f9e, 32'hc30b67fc} /* (13, 10, 15) {real, imag} */,
  {32'hc2718e51, 32'h41ba790a} /* (13, 10, 14) {real, imag} */,
  {32'h420d94c5, 32'h431686f9} /* (13, 10, 13) {real, imag} */,
  {32'h42f1452f, 32'hc290eb14} /* (13, 10, 12) {real, imag} */,
  {32'h432b6d16, 32'hc2c8dac3} /* (13, 10, 11) {real, imag} */,
  {32'h419815be, 32'h43085da1} /* (13, 10, 10) {real, imag} */,
  {32'h4218e090, 32'hc116d8e8} /* (13, 10, 9) {real, imag} */,
  {32'hc2d42db6, 32'h00000000} /* (13, 10, 8) {real, imag} */,
  {32'h4218e090, 32'h4116d8e8} /* (13, 10, 7) {real, imag} */,
  {32'h419815be, 32'hc3085da1} /* (13, 10, 6) {real, imag} */,
  {32'h432b6d16, 32'h42c8dac3} /* (13, 10, 5) {real, imag} */,
  {32'h42f1452f, 32'h4290eb14} /* (13, 10, 4) {real, imag} */,
  {32'h420d94c5, 32'hc31686f9} /* (13, 10, 3) {real, imag} */,
  {32'hc2718e51, 32'hc1ba790a} /* (13, 10, 2) {real, imag} */,
  {32'h42087f9e, 32'h430b67fc} /* (13, 10, 1) {real, imag} */,
  {32'h43189e31, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h432e9522, 32'hc33f455d} /* (13, 9, 15) {real, imag} */,
  {32'hc2899548, 32'hc2a64151} /* (13, 9, 14) {real, imag} */,
  {32'h41dd64e9, 32'hc2dce9aa} /* (13, 9, 13) {real, imag} */,
  {32'hc2e1ef8a, 32'hc2743e9e} /* (13, 9, 12) {real, imag} */,
  {32'hc2ca42ee, 32'hc2375dcc} /* (13, 9, 11) {real, imag} */,
  {32'hc1c3e9e3, 32'hc2490fa6} /* (13, 9, 10) {real, imag} */,
  {32'h41d89642, 32'h42f55fb8} /* (13, 9, 9) {real, imag} */,
  {32'h42c747fe, 32'h00000000} /* (13, 9, 8) {real, imag} */,
  {32'h41d89642, 32'hc2f55fb8} /* (13, 9, 7) {real, imag} */,
  {32'hc1c3e9e3, 32'h42490fa6} /* (13, 9, 6) {real, imag} */,
  {32'hc2ca42ee, 32'h42375dcc} /* (13, 9, 5) {real, imag} */,
  {32'hc2e1ef8a, 32'h42743e9e} /* (13, 9, 4) {real, imag} */,
  {32'h41dd64e9, 32'h42dce9aa} /* (13, 9, 3) {real, imag} */,
  {32'hc2899548, 32'h42a64151} /* (13, 9, 2) {real, imag} */,
  {32'h432e9522, 32'h433f455d} /* (13, 9, 1) {real, imag} */,
  {32'h435f5414, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'hc2921027, 32'hc344f4ba} /* (13, 8, 15) {real, imag} */,
  {32'hc21f1033, 32'h42c93cf2} /* (13, 8, 14) {real, imag} */,
  {32'hc27f95ce, 32'h41f408c0} /* (13, 8, 13) {real, imag} */,
  {32'hc0395ad0, 32'h417069e4} /* (13, 8, 12) {real, imag} */,
  {32'hc3081566, 32'h411b378a} /* (13, 8, 11) {real, imag} */,
  {32'hc2298593, 32'hc29d55f4} /* (13, 8, 10) {real, imag} */,
  {32'h425535f3, 32'hc2789b1e} /* (13, 8, 9) {real, imag} */,
  {32'h4047dde0, 32'h00000000} /* (13, 8, 8) {real, imag} */,
  {32'h425535f3, 32'h42789b1e} /* (13, 8, 7) {real, imag} */,
  {32'hc2298593, 32'h429d55f4} /* (13, 8, 6) {real, imag} */,
  {32'hc3081566, 32'hc11b378a} /* (13, 8, 5) {real, imag} */,
  {32'hc0395ad0, 32'hc17069e4} /* (13, 8, 4) {real, imag} */,
  {32'hc27f95ce, 32'hc1f408c0} /* (13, 8, 3) {real, imag} */,
  {32'hc21f1033, 32'hc2c93cf2} /* (13, 8, 2) {real, imag} */,
  {32'hc2921027, 32'h4344f4ba} /* (13, 8, 1) {real, imag} */,
  {32'hc2574643, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'hc34b6e58, 32'h414d93b0} /* (13, 7, 15) {real, imag} */,
  {32'hc2e00004, 32'h4373d95e} /* (13, 7, 14) {real, imag} */,
  {32'hc221c65a, 32'h431fd51d} /* (13, 7, 13) {real, imag} */,
  {32'h4183bca6, 32'hc2758e56} /* (13, 7, 12) {real, imag} */,
  {32'hc28770da, 32'hc2e8111c} /* (13, 7, 11) {real, imag} */,
  {32'hc29f5704, 32'h430f6712} /* (13, 7, 10) {real, imag} */,
  {32'hc2f92e46, 32'h40b592c0} /* (13, 7, 9) {real, imag} */,
  {32'h4104df04, 32'h00000000} /* (13, 7, 8) {real, imag} */,
  {32'hc2f92e46, 32'hc0b592c0} /* (13, 7, 7) {real, imag} */,
  {32'hc29f5704, 32'hc30f6712} /* (13, 7, 6) {real, imag} */,
  {32'hc28770da, 32'h42e8111c} /* (13, 7, 5) {real, imag} */,
  {32'h4183bca6, 32'h42758e56} /* (13, 7, 4) {real, imag} */,
  {32'hc221c65a, 32'hc31fd51d} /* (13, 7, 3) {real, imag} */,
  {32'hc2e00004, 32'hc373d95e} /* (13, 7, 2) {real, imag} */,
  {32'hc34b6e58, 32'hc14d93b0} /* (13, 7, 1) {real, imag} */,
  {32'h435a8f48, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'hc37e3a34, 32'hc2056e4d} /* (13, 6, 15) {real, imag} */,
  {32'h4313e651, 32'h42ad7464} /* (13, 6, 14) {real, imag} */,
  {32'h41e4c1ca, 32'h4220e1bc} /* (13, 6, 13) {real, imag} */,
  {32'hc31ac620, 32'hc0c36060} /* (13, 6, 12) {real, imag} */,
  {32'h4330f992, 32'hc21ca732} /* (13, 6, 11) {real, imag} */,
  {32'hc2b4edc0, 32'hc31f45f7} /* (13, 6, 10) {real, imag} */,
  {32'h432a9fc4, 32'h4322fb86} /* (13, 6, 9) {real, imag} */,
  {32'hc213a52c, 32'h00000000} /* (13, 6, 8) {real, imag} */,
  {32'h432a9fc4, 32'hc322fb86} /* (13, 6, 7) {real, imag} */,
  {32'hc2b4edc0, 32'h431f45f7} /* (13, 6, 6) {real, imag} */,
  {32'h4330f992, 32'h421ca732} /* (13, 6, 5) {real, imag} */,
  {32'hc31ac620, 32'h40c36060} /* (13, 6, 4) {real, imag} */,
  {32'h41e4c1ca, 32'hc220e1bc} /* (13, 6, 3) {real, imag} */,
  {32'h4313e651, 32'hc2ad7464} /* (13, 6, 2) {real, imag} */,
  {32'hc37e3a34, 32'h42056e4d} /* (13, 6, 1) {real, imag} */,
  {32'h4387a9c2, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'hc288e685, 32'h4312e4b1} /* (13, 5, 15) {real, imag} */,
  {32'hc2768066, 32'h41e050e8} /* (13, 5, 14) {real, imag} */,
  {32'hc1ebb998, 32'hc28a7d16} /* (13, 5, 13) {real, imag} */,
  {32'hc2061588, 32'hc2399cfe} /* (13, 5, 12) {real, imag} */,
  {32'h42457b34, 32'h3f3bfbc0} /* (13, 5, 11) {real, imag} */,
  {32'hc1ee442c, 32'h40c36594} /* (13, 5, 10) {real, imag} */,
  {32'hc0e72b7a, 32'hc2bdc406} /* (13, 5, 9) {real, imag} */,
  {32'h41d21cc6, 32'h00000000} /* (13, 5, 8) {real, imag} */,
  {32'hc0e72b7a, 32'h42bdc406} /* (13, 5, 7) {real, imag} */,
  {32'hc1ee442c, 32'hc0c36594} /* (13, 5, 6) {real, imag} */,
  {32'h42457b34, 32'hbf3bfbc0} /* (13, 5, 5) {real, imag} */,
  {32'hc2061588, 32'h42399cfe} /* (13, 5, 4) {real, imag} */,
  {32'hc1ebb998, 32'h428a7d16} /* (13, 5, 3) {real, imag} */,
  {32'hc2768066, 32'hc1e050e8} /* (13, 5, 2) {real, imag} */,
  {32'hc288e685, 32'hc312e4b1} /* (13, 5, 1) {real, imag} */,
  {32'h43a47771, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h424af122, 32'hc2ffda90} /* (13, 4, 15) {real, imag} */,
  {32'h430af508, 32'hc1022195} /* (13, 4, 14) {real, imag} */,
  {32'hc31fcef8, 32'h4290013e} /* (13, 4, 13) {real, imag} */,
  {32'h420506db, 32'hc25ec848} /* (13, 4, 12) {real, imag} */,
  {32'h42b7d90e, 32'hc2842535} /* (13, 4, 11) {real, imag} */,
  {32'hc1605f18, 32'h42dd5eb4} /* (13, 4, 10) {real, imag} */,
  {32'hc2eb7c8e, 32'h42f4260a} /* (13, 4, 9) {real, imag} */,
  {32'h4227ffab, 32'h00000000} /* (13, 4, 8) {real, imag} */,
  {32'hc2eb7c8e, 32'hc2f4260a} /* (13, 4, 7) {real, imag} */,
  {32'hc1605f18, 32'hc2dd5eb4} /* (13, 4, 6) {real, imag} */,
  {32'h42b7d90e, 32'h42842535} /* (13, 4, 5) {real, imag} */,
  {32'h420506db, 32'h425ec848} /* (13, 4, 4) {real, imag} */,
  {32'hc31fcef8, 32'hc290013e} /* (13, 4, 3) {real, imag} */,
  {32'h430af508, 32'h41022195} /* (13, 4, 2) {real, imag} */,
  {32'h424af122, 32'h42ffda90} /* (13, 4, 1) {real, imag} */,
  {32'h4371eb6f, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'hc1b6e08c, 32'hc3a0b02a} /* (13, 3, 15) {real, imag} */,
  {32'hc25bebc2, 32'h42a03fc6} /* (13, 3, 14) {real, imag} */,
  {32'hc3829f92, 32'h43771ee2} /* (13, 3, 13) {real, imag} */,
  {32'h439f3972, 32'hc27dbefe} /* (13, 3, 12) {real, imag} */,
  {32'h4296d59e, 32'hc29225a8} /* (13, 3, 11) {real, imag} */,
  {32'h43221548, 32'hc31c29ee} /* (13, 3, 10) {real, imag} */,
  {32'h411e5b1a, 32'h418c1c4e} /* (13, 3, 9) {real, imag} */,
  {32'hc2c0f3cc, 32'h00000000} /* (13, 3, 8) {real, imag} */,
  {32'h411e5b1a, 32'hc18c1c4e} /* (13, 3, 7) {real, imag} */,
  {32'h43221548, 32'h431c29ee} /* (13, 3, 6) {real, imag} */,
  {32'h4296d59e, 32'h429225a8} /* (13, 3, 5) {real, imag} */,
  {32'h439f3972, 32'h427dbefe} /* (13, 3, 4) {real, imag} */,
  {32'hc3829f92, 32'hc3771ee2} /* (13, 3, 3) {real, imag} */,
  {32'hc25bebc2, 32'hc2a03fc6} /* (13, 3, 2) {real, imag} */,
  {32'hc1b6e08c, 32'h43a0b02a} /* (13, 3, 1) {real, imag} */,
  {32'h43965df4, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h4360486a, 32'hc3897d76} /* (13, 2, 15) {real, imag} */,
  {32'hc2542bc9, 32'hc2bcc43b} /* (13, 2, 14) {real, imag} */,
  {32'hc335400b, 32'h4302e34c} /* (13, 2, 13) {real, imag} */,
  {32'h42706aa6, 32'hc2c60471} /* (13, 2, 12) {real, imag} */,
  {32'h415c6868, 32'hc0caf056} /* (13, 2, 11) {real, imag} */,
  {32'hc2c75db2, 32'h4257f605} /* (13, 2, 10) {real, imag} */,
  {32'h42a57ccd, 32'hc14c5c40} /* (13, 2, 9) {real, imag} */,
  {32'hc2b09c15, 32'h00000000} /* (13, 2, 8) {real, imag} */,
  {32'h42a57ccd, 32'h414c5c40} /* (13, 2, 7) {real, imag} */,
  {32'hc2c75db2, 32'hc257f605} /* (13, 2, 6) {real, imag} */,
  {32'h415c6868, 32'h40caf056} /* (13, 2, 5) {real, imag} */,
  {32'h42706aa6, 32'h42c60471} /* (13, 2, 4) {real, imag} */,
  {32'hc335400b, 32'hc302e34c} /* (13, 2, 3) {real, imag} */,
  {32'hc2542bc9, 32'h42bcc43b} /* (13, 2, 2) {real, imag} */,
  {32'h4360486a, 32'h43897d76} /* (13, 2, 1) {real, imag} */,
  {32'h42cb0c1e, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h4325e3bb, 32'hc3ab5304} /* (13, 1, 15) {real, imag} */,
  {32'h4224ba5c, 32'hc2f0a316} /* (13, 1, 14) {real, imag} */,
  {32'hc2dc9b1b, 32'hc102358c} /* (13, 1, 13) {real, imag} */,
  {32'h41814b92, 32'h4389630d} /* (13, 1, 12) {real, imag} */,
  {32'hc1a200f0, 32'hc329ba4a} /* (13, 1, 11) {real, imag} */,
  {32'hc209dab1, 32'hc27c904c} /* (13, 1, 10) {real, imag} */,
  {32'hc1809b66, 32'h41893ee2} /* (13, 1, 9) {real, imag} */,
  {32'hc21ff850, 32'h00000000} /* (13, 1, 8) {real, imag} */,
  {32'hc1809b66, 32'hc1893ee2} /* (13, 1, 7) {real, imag} */,
  {32'hc209dab1, 32'h427c904c} /* (13, 1, 6) {real, imag} */,
  {32'hc1a200f0, 32'h4329ba4a} /* (13, 1, 5) {real, imag} */,
  {32'h41814b92, 32'hc389630d} /* (13, 1, 4) {real, imag} */,
  {32'hc2dc9b1b, 32'h4102358c} /* (13, 1, 3) {real, imag} */,
  {32'h4224ba5c, 32'h42f0a316} /* (13, 1, 2) {real, imag} */,
  {32'h4325e3bb, 32'h43ab5304} /* (13, 1, 1) {real, imag} */,
  {32'hc255096c, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h427b0232, 32'hc2f2da94} /* (13, 0, 15) {real, imag} */,
  {32'hc23879df, 32'hc242ca70} /* (13, 0, 14) {real, imag} */,
  {32'hc2edcad9, 32'hc14f61f4} /* (13, 0, 13) {real, imag} */,
  {32'h42f8c77a, 32'h42ee3158} /* (13, 0, 12) {real, imag} */,
  {32'h42220436, 32'hc2647646} /* (13, 0, 11) {real, imag} */,
  {32'h42491171, 32'hc223edf2} /* (13, 0, 10) {real, imag} */,
  {32'hc26ae427, 32'h41804358} /* (13, 0, 9) {real, imag} */,
  {32'hc1ae3ef0, 32'h00000000} /* (13, 0, 8) {real, imag} */,
  {32'hc26ae427, 32'hc1804358} /* (13, 0, 7) {real, imag} */,
  {32'h42491171, 32'h4223edf2} /* (13, 0, 6) {real, imag} */,
  {32'h42220436, 32'h42647646} /* (13, 0, 5) {real, imag} */,
  {32'h42f8c77a, 32'hc2ee3158} /* (13, 0, 4) {real, imag} */,
  {32'hc2edcad9, 32'h414f61f4} /* (13, 0, 3) {real, imag} */,
  {32'hc23879df, 32'h4242ca70} /* (13, 0, 2) {real, imag} */,
  {32'h427b0232, 32'h42f2da94} /* (13, 0, 1) {real, imag} */,
  {32'h42c265e2, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h4335610c, 32'h42d56467} /* (12, 15, 15) {real, imag} */,
  {32'hc2fe9607, 32'hc1be4384} /* (12, 15, 14) {real, imag} */,
  {32'hc1aa601d, 32'hc1b8b3b4} /* (12, 15, 13) {real, imag} */,
  {32'h41e38164, 32'hc30f90e2} /* (12, 15, 12) {real, imag} */,
  {32'hc10aff26, 32'hc298366b} /* (12, 15, 11) {real, imag} */,
  {32'hc1cdfdb4, 32'h428a8b4f} /* (12, 15, 10) {real, imag} */,
  {32'h4204acb6, 32'hbe6dd500} /* (12, 15, 9) {real, imag} */,
  {32'hc0373a48, 32'h00000000} /* (12, 15, 8) {real, imag} */,
  {32'h4204acb6, 32'h3e6dd500} /* (12, 15, 7) {real, imag} */,
  {32'hc1cdfdb4, 32'hc28a8b4f} /* (12, 15, 6) {real, imag} */,
  {32'hc10aff26, 32'h4298366b} /* (12, 15, 5) {real, imag} */,
  {32'h41e38164, 32'h430f90e2} /* (12, 15, 4) {real, imag} */,
  {32'hc1aa601d, 32'h41b8b3b4} /* (12, 15, 3) {real, imag} */,
  {32'hc2fe9607, 32'h41be4384} /* (12, 15, 2) {real, imag} */,
  {32'h4335610c, 32'hc2d56467} /* (12, 15, 1) {real, imag} */,
  {32'h415275d8, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'h430a4d74, 32'h43913342} /* (12, 14, 15) {real, imag} */,
  {32'h413e0c14, 32'hc310da8f} /* (12, 14, 14) {real, imag} */,
  {32'hc209f4b3, 32'h42728e5d} /* (12, 14, 13) {real, imag} */,
  {32'h41375790, 32'hc319553f} /* (12, 14, 12) {real, imag} */,
  {32'hc282da4e, 32'hc2899a2b} /* (12, 14, 11) {real, imag} */,
  {32'hc2dd53aa, 32'h431ea756} /* (12, 14, 10) {real, imag} */,
  {32'h41dc235a, 32'hc30a5fa6} /* (12, 14, 9) {real, imag} */,
  {32'hc30ded90, 32'h00000000} /* (12, 14, 8) {real, imag} */,
  {32'h41dc235a, 32'h430a5fa6} /* (12, 14, 7) {real, imag} */,
  {32'hc2dd53aa, 32'hc31ea756} /* (12, 14, 6) {real, imag} */,
  {32'hc282da4e, 32'h42899a2b} /* (12, 14, 5) {real, imag} */,
  {32'h41375790, 32'h4319553f} /* (12, 14, 4) {real, imag} */,
  {32'hc209f4b3, 32'hc2728e5d} /* (12, 14, 3) {real, imag} */,
  {32'h413e0c14, 32'h4310da8f} /* (12, 14, 2) {real, imag} */,
  {32'h430a4d74, 32'hc3913342} /* (12, 14, 1) {real, imag} */,
  {32'hc288c17e, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'h41fc3ab0, 32'h42748e25} /* (12, 13, 15) {real, imag} */,
  {32'hc110bfa6, 32'hc2ab64c9} /* (12, 13, 14) {real, imag} */,
  {32'h42aa41c4, 32'hc311a31c} /* (12, 13, 13) {real, imag} */,
  {32'hc1cf2f28, 32'h421394c8} /* (12, 13, 12) {real, imag} */,
  {32'h40fb5e18, 32'h425241ec} /* (12, 13, 11) {real, imag} */,
  {32'h41bd4aae, 32'hc24770b4} /* (12, 13, 10) {real, imag} */,
  {32'hc2842f8f, 32'hc2aa79f3} /* (12, 13, 9) {real, imag} */,
  {32'hc1fcdc12, 32'h00000000} /* (12, 13, 8) {real, imag} */,
  {32'hc2842f8f, 32'h42aa79f3} /* (12, 13, 7) {real, imag} */,
  {32'h41bd4aae, 32'h424770b4} /* (12, 13, 6) {real, imag} */,
  {32'h40fb5e18, 32'hc25241ec} /* (12, 13, 5) {real, imag} */,
  {32'hc1cf2f28, 32'hc21394c8} /* (12, 13, 4) {real, imag} */,
  {32'h42aa41c4, 32'h4311a31c} /* (12, 13, 3) {real, imag} */,
  {32'hc110bfa6, 32'h42ab64c9} /* (12, 13, 2) {real, imag} */,
  {32'h41fc3ab0, 32'hc2748e25} /* (12, 13, 1) {real, imag} */,
  {32'h42f8b6de, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'h41e4a45c, 32'hc304a6dc} /* (12, 12, 15) {real, imag} */,
  {32'h3f451c40, 32'hc29d2966} /* (12, 12, 14) {real, imag} */,
  {32'h42d6ded6, 32'hc36aaaff} /* (12, 12, 13) {real, imag} */,
  {32'h421bf5f6, 32'h41d21c13} /* (12, 12, 12) {real, imag} */,
  {32'hc2298e4c, 32'hc1e0fdb8} /* (12, 12, 11) {real, imag} */,
  {32'hc19cfed7, 32'h42c1d06c} /* (12, 12, 10) {real, imag} */,
  {32'h423c5832, 32'h431a94ca} /* (12, 12, 9) {real, imag} */,
  {32'h41d75822, 32'h00000000} /* (12, 12, 8) {real, imag} */,
  {32'h423c5832, 32'hc31a94ca} /* (12, 12, 7) {real, imag} */,
  {32'hc19cfed7, 32'hc2c1d06c} /* (12, 12, 6) {real, imag} */,
  {32'hc2298e4c, 32'h41e0fdb8} /* (12, 12, 5) {real, imag} */,
  {32'h421bf5f6, 32'hc1d21c13} /* (12, 12, 4) {real, imag} */,
  {32'h42d6ded6, 32'h436aaaff} /* (12, 12, 3) {real, imag} */,
  {32'h3f451c40, 32'h429d2966} /* (12, 12, 2) {real, imag} */,
  {32'h41e4a45c, 32'h4304a6dc} /* (12, 12, 1) {real, imag} */,
  {32'h431e86e9, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'hc2d97cfe, 32'hc3015a0d} /* (12, 11, 15) {real, imag} */,
  {32'h42d42342, 32'h428e3af5} /* (12, 11, 14) {real, imag} */,
  {32'hc1c5bc7e, 32'h4314b877} /* (12, 11, 13) {real, imag} */,
  {32'h4287cf3f, 32'hc24b7978} /* (12, 11, 12) {real, imag} */,
  {32'hc25543c6, 32'hc2aa1231} /* (12, 11, 11) {real, imag} */,
  {32'hc1119398, 32'hc2628e04} /* (12, 11, 10) {real, imag} */,
  {32'h42ad9cfc, 32'h40d9ab5c} /* (12, 11, 9) {real, imag} */,
  {32'hc28a4970, 32'h00000000} /* (12, 11, 8) {real, imag} */,
  {32'h42ad9cfc, 32'hc0d9ab5c} /* (12, 11, 7) {real, imag} */,
  {32'hc1119398, 32'h42628e04} /* (12, 11, 6) {real, imag} */,
  {32'hc25543c6, 32'h42aa1231} /* (12, 11, 5) {real, imag} */,
  {32'h4287cf3f, 32'h424b7978} /* (12, 11, 4) {real, imag} */,
  {32'hc1c5bc7e, 32'hc314b877} /* (12, 11, 3) {real, imag} */,
  {32'h42d42342, 32'hc28e3af5} /* (12, 11, 2) {real, imag} */,
  {32'hc2d97cfe, 32'h43015a0d} /* (12, 11, 1) {real, imag} */,
  {32'h43cd7f4a, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'hc2382a38, 32'hc35a008c} /* (12, 10, 15) {real, imag} */,
  {32'h42b40633, 32'h4302c86c} /* (12, 10, 14) {real, imag} */,
  {32'h42360cb8, 32'h42cb6164} /* (12, 10, 13) {real, imag} */,
  {32'h3f400b00, 32'hc2d62354} /* (12, 10, 12) {real, imag} */,
  {32'h4260478c, 32'hc1c659f2} /* (12, 10, 11) {real, imag} */,
  {32'hc2338c30, 32'h410cb640} /* (12, 10, 10) {real, imag} */,
  {32'hc2ebeee0, 32'hc2ada4ae} /* (12, 10, 9) {real, imag} */,
  {32'h42989616, 32'h00000000} /* (12, 10, 8) {real, imag} */,
  {32'hc2ebeee0, 32'h42ada4ae} /* (12, 10, 7) {real, imag} */,
  {32'hc2338c30, 32'hc10cb640} /* (12, 10, 6) {real, imag} */,
  {32'h4260478c, 32'h41c659f2} /* (12, 10, 5) {real, imag} */,
  {32'h3f400b00, 32'h42d62354} /* (12, 10, 4) {real, imag} */,
  {32'h42360cb8, 32'hc2cb6164} /* (12, 10, 3) {real, imag} */,
  {32'h42b40633, 32'hc302c86c} /* (12, 10, 2) {real, imag} */,
  {32'hc2382a38, 32'h435a008c} /* (12, 10, 1) {real, imag} */,
  {32'h43a35fd2, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h42ffa350, 32'hc38848fa} /* (12, 9, 15) {real, imag} */,
  {32'h42195522, 32'h43280ceb} /* (12, 9, 14) {real, imag} */,
  {32'h42f8788f, 32'h43239b8a} /* (12, 9, 13) {real, imag} */,
  {32'hc28d3c55, 32'hc1e16621} /* (12, 9, 12) {real, imag} */,
  {32'h422388f5, 32'h41ba1d4f} /* (12, 9, 11) {real, imag} */,
  {32'hc3090546, 32'h41de29e0} /* (12, 9, 10) {real, imag} */,
  {32'h4299aec6, 32'hc28bab0e} /* (12, 9, 9) {real, imag} */,
  {32'hc2d2de02, 32'h00000000} /* (12, 9, 8) {real, imag} */,
  {32'h4299aec6, 32'h428bab0e} /* (12, 9, 7) {real, imag} */,
  {32'hc3090546, 32'hc1de29e0} /* (12, 9, 6) {real, imag} */,
  {32'h422388f5, 32'hc1ba1d4f} /* (12, 9, 5) {real, imag} */,
  {32'hc28d3c55, 32'h41e16621} /* (12, 9, 4) {real, imag} */,
  {32'h42f8788f, 32'hc3239b8a} /* (12, 9, 3) {real, imag} */,
  {32'h42195522, 32'hc3280ceb} /* (12, 9, 2) {real, imag} */,
  {32'h42ffa350, 32'h438848fa} /* (12, 9, 1) {real, imag} */,
  {32'h42f9dce3, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'h419fa19e, 32'hc365c881} /* (12, 8, 15) {real, imag} */,
  {32'h4357e49a, 32'h420adf5b} /* (12, 8, 14) {real, imag} */,
  {32'hc23cdaa9, 32'h4238aab4} /* (12, 8, 13) {real, imag} */,
  {32'hc210cf1e, 32'h40a19df4} /* (12, 8, 12) {real, imag} */,
  {32'h414c6683, 32'h42672142} /* (12, 8, 11) {real, imag} */,
  {32'hc095cfbc, 32'h42e8dff2} /* (12, 8, 10) {real, imag} */,
  {32'hc23ebd67, 32'hc25a361a} /* (12, 8, 9) {real, imag} */,
  {32'h422640d0, 32'h00000000} /* (12, 8, 8) {real, imag} */,
  {32'hc23ebd67, 32'h425a361a} /* (12, 8, 7) {real, imag} */,
  {32'hc095cfbc, 32'hc2e8dff2} /* (12, 8, 6) {real, imag} */,
  {32'h414c6683, 32'hc2672142} /* (12, 8, 5) {real, imag} */,
  {32'hc210cf1e, 32'hc0a19df4} /* (12, 8, 4) {real, imag} */,
  {32'hc23cdaa9, 32'hc238aab4} /* (12, 8, 3) {real, imag} */,
  {32'h4357e49a, 32'hc20adf5b} /* (12, 8, 2) {real, imag} */,
  {32'h419fa19e, 32'h4365c881} /* (12, 8, 1) {real, imag} */,
  {32'hc25b2abc, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'hc387b79e, 32'hc1febbd8} /* (12, 7, 15) {real, imag} */,
  {32'h424160f6, 32'h43201dc1} /* (12, 7, 14) {real, imag} */,
  {32'h404eb9e0, 32'h42fced1b} /* (12, 7, 13) {real, imag} */,
  {32'h40ed6b70, 32'hc0c1309c} /* (12, 7, 12) {real, imag} */,
  {32'h4203a93f, 32'hc15527de} /* (12, 7, 11) {real, imag} */,
  {32'h42fb56f8, 32'h41d28b18} /* (12, 7, 10) {real, imag} */,
  {32'hc101edbc, 32'hc23b9657} /* (12, 7, 9) {real, imag} */,
  {32'h41f6be12, 32'h00000000} /* (12, 7, 8) {real, imag} */,
  {32'hc101edbc, 32'h423b9657} /* (12, 7, 7) {real, imag} */,
  {32'h42fb56f8, 32'hc1d28b18} /* (12, 7, 6) {real, imag} */,
  {32'h4203a93f, 32'h415527de} /* (12, 7, 5) {real, imag} */,
  {32'h40ed6b70, 32'h40c1309c} /* (12, 7, 4) {real, imag} */,
  {32'h404eb9e0, 32'hc2fced1b} /* (12, 7, 3) {real, imag} */,
  {32'h424160f6, 32'hc3201dc1} /* (12, 7, 2) {real, imag} */,
  {32'hc387b79e, 32'h41febbd8} /* (12, 7, 1) {real, imag} */,
  {32'hc19497f4, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'hc3caf2a9, 32'h434f42f2} /* (12, 6, 15) {real, imag} */,
  {32'hc31085a2, 32'hc2b9605c} /* (12, 6, 14) {real, imag} */,
  {32'h4283653d, 32'hc2b81270} /* (12, 6, 13) {real, imag} */,
  {32'h42da178c, 32'h408b3600} /* (12, 6, 12) {real, imag} */,
  {32'h40df6e40, 32'h425eaab3} /* (12, 6, 11) {real, imag} */,
  {32'h4306d0e4, 32'hc22e383a} /* (12, 6, 10) {real, imag} */,
  {32'h434876ac, 32'hc2563bd8} /* (12, 6, 9) {real, imag} */,
  {32'hc1fe7000, 32'h00000000} /* (12, 6, 8) {real, imag} */,
  {32'h434876ac, 32'h42563bd8} /* (12, 6, 7) {real, imag} */,
  {32'h4306d0e4, 32'h422e383a} /* (12, 6, 6) {real, imag} */,
  {32'h40df6e40, 32'hc25eaab3} /* (12, 6, 5) {real, imag} */,
  {32'h42da178c, 32'hc08b3600} /* (12, 6, 4) {real, imag} */,
  {32'h4283653d, 32'h42b81270} /* (12, 6, 3) {real, imag} */,
  {32'hc31085a2, 32'h42b9605c} /* (12, 6, 2) {real, imag} */,
  {32'hc3caf2a9, 32'hc34f42f2} /* (12, 6, 1) {real, imag} */,
  {32'h4359830c, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'hc23aae14, 32'h43399b0f} /* (12, 5, 15) {real, imag} */,
  {32'hc1a7e718, 32'hc2ff2247} /* (12, 5, 14) {real, imag} */,
  {32'hc26808a9, 32'hc0df7fa0} /* (12, 5, 13) {real, imag} */,
  {32'hc2f7e081, 32'hc1d4b450} /* (12, 5, 12) {real, imag} */,
  {32'h432637b0, 32'hc25dda46} /* (12, 5, 11) {real, imag} */,
  {32'hc325aac0, 32'h428fe1dc} /* (12, 5, 10) {real, imag} */,
  {32'h42eb6d38, 32'hc01bc478} /* (12, 5, 9) {real, imag} */,
  {32'hc1bbad8a, 32'h00000000} /* (12, 5, 8) {real, imag} */,
  {32'h42eb6d38, 32'h401bc478} /* (12, 5, 7) {real, imag} */,
  {32'hc325aac0, 32'hc28fe1dc} /* (12, 5, 6) {real, imag} */,
  {32'h432637b0, 32'h425dda46} /* (12, 5, 5) {real, imag} */,
  {32'hc2f7e081, 32'h41d4b450} /* (12, 5, 4) {real, imag} */,
  {32'hc26808a9, 32'h40df7fa0} /* (12, 5, 3) {real, imag} */,
  {32'hc1a7e718, 32'h42ff2247} /* (12, 5, 2) {real, imag} */,
  {32'hc23aae14, 32'hc3399b0f} /* (12, 5, 1) {real, imag} */,
  {32'h438ada3a, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'hc02d8ac0, 32'h42e52533} /* (12, 4, 15) {real, imag} */,
  {32'hc2ec86c2, 32'hc2bdd63a} /* (12, 4, 14) {real, imag} */,
  {32'hc26301bb, 32'h42d7b812} /* (12, 4, 13) {real, imag} */,
  {32'h42d652a5, 32'hc114d61a} /* (12, 4, 12) {real, imag} */,
  {32'hc2560b9e, 32'hc282ec4a} /* (12, 4, 11) {real, imag} */,
  {32'hc281af90, 32'hc2af3bc4} /* (12, 4, 10) {real, imag} */,
  {32'h41637416, 32'h42d246ac} /* (12, 4, 9) {real, imag} */,
  {32'h40931cbc, 32'h00000000} /* (12, 4, 8) {real, imag} */,
  {32'h41637416, 32'hc2d246ac} /* (12, 4, 7) {real, imag} */,
  {32'hc281af90, 32'h42af3bc4} /* (12, 4, 6) {real, imag} */,
  {32'hc2560b9e, 32'h4282ec4a} /* (12, 4, 5) {real, imag} */,
  {32'h42d652a5, 32'h4114d61a} /* (12, 4, 4) {real, imag} */,
  {32'hc26301bb, 32'hc2d7b812} /* (12, 4, 3) {real, imag} */,
  {32'hc2ec86c2, 32'h42bdd63a} /* (12, 4, 2) {real, imag} */,
  {32'hc02d8ac0, 32'hc2e52533} /* (12, 4, 1) {real, imag} */,
  {32'h43cc4348, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'hc29f2c98, 32'hc2bf0ef2} /* (12, 3, 15) {real, imag} */,
  {32'hc260561a, 32'hc3043f6a} /* (12, 3, 14) {real, imag} */,
  {32'h41cd4b16, 32'h427fdb99} /* (12, 3, 13) {real, imag} */,
  {32'h41bd4c5c, 32'hc233da54} /* (12, 3, 12) {real, imag} */,
  {32'h42bb4238, 32'h4248d57c} /* (12, 3, 11) {real, imag} */,
  {32'hc30c11e3, 32'h42bfef64} /* (12, 3, 10) {real, imag} */,
  {32'hc2f9566d, 32'h4203fa02} /* (12, 3, 9) {real, imag} */,
  {32'h4268f2b7, 32'h00000000} /* (12, 3, 8) {real, imag} */,
  {32'hc2f9566d, 32'hc203fa02} /* (12, 3, 7) {real, imag} */,
  {32'hc30c11e3, 32'hc2bfef64} /* (12, 3, 6) {real, imag} */,
  {32'h42bb4238, 32'hc248d57c} /* (12, 3, 5) {real, imag} */,
  {32'h41bd4c5c, 32'h4233da54} /* (12, 3, 4) {real, imag} */,
  {32'h41cd4b16, 32'hc27fdb99} /* (12, 3, 3) {real, imag} */,
  {32'hc260561a, 32'h43043f6a} /* (12, 3, 2) {real, imag} */,
  {32'hc29f2c98, 32'h42bf0ef2} /* (12, 3, 1) {real, imag} */,
  {32'h43a0ca36, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'h427f89c2, 32'hc306f4ee} /* (12, 2, 15) {real, imag} */,
  {32'h420adf83, 32'h426aa2db} /* (12, 2, 14) {real, imag} */,
  {32'hc20414e3, 32'h42d58eda} /* (12, 2, 13) {real, imag} */,
  {32'hc186fa02, 32'hc24f209c} /* (12, 2, 12) {real, imag} */,
  {32'h42f144ae, 32'h42576c46} /* (12, 2, 11) {real, imag} */,
  {32'hc2a03bba, 32'h417c0e20} /* (12, 2, 10) {real, imag} */,
  {32'hc2859ee2, 32'h4195ba3c} /* (12, 2, 9) {real, imag} */,
  {32'hc2cf26bd, 32'h00000000} /* (12, 2, 8) {real, imag} */,
  {32'hc2859ee2, 32'hc195ba3c} /* (12, 2, 7) {real, imag} */,
  {32'hc2a03bba, 32'hc17c0e20} /* (12, 2, 6) {real, imag} */,
  {32'h42f144ae, 32'hc2576c46} /* (12, 2, 5) {real, imag} */,
  {32'hc186fa02, 32'h424f209c} /* (12, 2, 4) {real, imag} */,
  {32'hc20414e3, 32'hc2d58eda} /* (12, 2, 3) {real, imag} */,
  {32'h420adf83, 32'hc26aa2db} /* (12, 2, 2) {real, imag} */,
  {32'h427f89c2, 32'h4306f4ee} /* (12, 2, 1) {real, imag} */,
  {32'h4211e624, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'hc2895861, 32'hc3273e0e} /* (12, 1, 15) {real, imag} */,
  {32'hc2048c8a, 32'h42905467} /* (12, 1, 14) {real, imag} */,
  {32'hc01c6618, 32'h426c5a26} /* (12, 1, 13) {real, imag} */,
  {32'h42a4d3ef, 32'hc25c0814} /* (12, 1, 12) {real, imag} */,
  {32'h3faec490, 32'h42a8c0ef} /* (12, 1, 11) {real, imag} */,
  {32'h42c56482, 32'hc2989ed9} /* (12, 1, 10) {real, imag} */,
  {32'h415bf9aa, 32'hc2f43608} /* (12, 1, 9) {real, imag} */,
  {32'hc1a36b7b, 32'h00000000} /* (12, 1, 8) {real, imag} */,
  {32'h415bf9aa, 32'h42f43608} /* (12, 1, 7) {real, imag} */,
  {32'h42c56482, 32'h42989ed9} /* (12, 1, 6) {real, imag} */,
  {32'h3faec490, 32'hc2a8c0ef} /* (12, 1, 5) {real, imag} */,
  {32'h42a4d3ef, 32'h425c0814} /* (12, 1, 4) {real, imag} */,
  {32'hc01c6618, 32'hc26c5a26} /* (12, 1, 3) {real, imag} */,
  {32'hc2048c8a, 32'hc2905467} /* (12, 1, 2) {real, imag} */,
  {32'hc2895861, 32'h43273e0e} /* (12, 1, 1) {real, imag} */,
  {32'h42b844b7, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'h42a333ae, 32'hc190cc78} /* (12, 0, 15) {real, imag} */,
  {32'h417bdee0, 32'h42702a47} /* (12, 0, 14) {real, imag} */,
  {32'hc226a949, 32'hc2112474} /* (12, 0, 13) {real, imag} */,
  {32'h4251ebcc, 32'h40cbfd74} /* (12, 0, 12) {real, imag} */,
  {32'hc103fa13, 32'h408c4010} /* (12, 0, 11) {real, imag} */,
  {32'h410f5ea2, 32'h3f405800} /* (12, 0, 10) {real, imag} */,
  {32'hbf51d940, 32'hc0eb2e0c} /* (12, 0, 9) {real, imag} */,
  {32'h42097b6e, 32'h00000000} /* (12, 0, 8) {real, imag} */,
  {32'hbf51d940, 32'h40eb2e0c} /* (12, 0, 7) {real, imag} */,
  {32'h410f5ea2, 32'hbf405800} /* (12, 0, 6) {real, imag} */,
  {32'hc103fa13, 32'hc08c4010} /* (12, 0, 5) {real, imag} */,
  {32'h4251ebcc, 32'hc0cbfd74} /* (12, 0, 4) {real, imag} */,
  {32'hc226a949, 32'h42112474} /* (12, 0, 3) {real, imag} */,
  {32'h417bdee0, 32'hc2702a47} /* (12, 0, 2) {real, imag} */,
  {32'h42a333ae, 32'h4190cc78} /* (12, 0, 1) {real, imag} */,
  {32'h4316b3dd, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h4315caff, 32'h420ee14e} /* (11, 15, 15) {real, imag} */,
  {32'hc33f3e80, 32'hc2c4ae8b} /* (11, 15, 14) {real, imag} */,
  {32'h4308dd44, 32'hc278314e} /* (11, 15, 13) {real, imag} */,
  {32'h41a26a30, 32'hc2553c4e} /* (11, 15, 12) {real, imag} */,
  {32'h4292ca1d, 32'h421fd062} /* (11, 15, 11) {real, imag} */,
  {32'hc300f1d8, 32'h43099add} /* (11, 15, 10) {real, imag} */,
  {32'hc2543fe5, 32'h41da9640} /* (11, 15, 9) {real, imag} */,
  {32'hc25fcb04, 32'h00000000} /* (11, 15, 8) {real, imag} */,
  {32'hc2543fe5, 32'hc1da9640} /* (11, 15, 7) {real, imag} */,
  {32'hc300f1d8, 32'hc3099add} /* (11, 15, 6) {real, imag} */,
  {32'h4292ca1d, 32'hc21fd062} /* (11, 15, 5) {real, imag} */,
  {32'h41a26a30, 32'h42553c4e} /* (11, 15, 4) {real, imag} */,
  {32'h4308dd44, 32'h4278314e} /* (11, 15, 3) {real, imag} */,
  {32'hc33f3e80, 32'h42c4ae8b} /* (11, 15, 2) {real, imag} */,
  {32'h4315caff, 32'hc20ee14e} /* (11, 15, 1) {real, imag} */,
  {32'h433bd86e, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'h4141d594, 32'h42bed0f2} /* (11, 14, 15) {real, imag} */,
  {32'hc30c9383, 32'hc31645dd} /* (11, 14, 14) {real, imag} */,
  {32'h42b99196, 32'hc2dd277a} /* (11, 14, 13) {real, imag} */,
  {32'hc2d5c2ca, 32'hc2cbcc56} /* (11, 14, 12) {real, imag} */,
  {32'h42b8b108, 32'hc1c22cf0} /* (11, 14, 11) {real, imag} */,
  {32'h41c58620, 32'hc180ac0e} /* (11, 14, 10) {real, imag} */,
  {32'h4242c7fa, 32'hc25d8c41} /* (11, 14, 9) {real, imag} */,
  {32'hc349f24a, 32'h00000000} /* (11, 14, 8) {real, imag} */,
  {32'h4242c7fa, 32'h425d8c41} /* (11, 14, 7) {real, imag} */,
  {32'h41c58620, 32'h4180ac0e} /* (11, 14, 6) {real, imag} */,
  {32'h42b8b108, 32'h41c22cf0} /* (11, 14, 5) {real, imag} */,
  {32'hc2d5c2ca, 32'h42cbcc56} /* (11, 14, 4) {real, imag} */,
  {32'h42b99196, 32'h42dd277a} /* (11, 14, 3) {real, imag} */,
  {32'hc30c9383, 32'h431645dd} /* (11, 14, 2) {real, imag} */,
  {32'h4141d594, 32'hc2bed0f2} /* (11, 14, 1) {real, imag} */,
  {32'h43de8af0, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'hc2d17b5a, 32'h42df6a92} /* (11, 13, 15) {real, imag} */,
  {32'h42f030d4, 32'hc3382e04} /* (11, 13, 14) {real, imag} */,
  {32'hc2ba6c4e, 32'hc2991cac} /* (11, 13, 13) {real, imag} */,
  {32'hc12c2cb2, 32'h41857db4} /* (11, 13, 12) {real, imag} */,
  {32'h3f9b3650, 32'h43974380} /* (11, 13, 11) {real, imag} */,
  {32'hc301c7b1, 32'h4272b790} /* (11, 13, 10) {real, imag} */,
  {32'h4325770a, 32'h412b9c0c} /* (11, 13, 9) {real, imag} */,
  {32'hc22d8c68, 32'h00000000} /* (11, 13, 8) {real, imag} */,
  {32'h4325770a, 32'hc12b9c0c} /* (11, 13, 7) {real, imag} */,
  {32'hc301c7b1, 32'hc272b790} /* (11, 13, 6) {real, imag} */,
  {32'h3f9b3650, 32'hc3974380} /* (11, 13, 5) {real, imag} */,
  {32'hc12c2cb2, 32'hc1857db4} /* (11, 13, 4) {real, imag} */,
  {32'hc2ba6c4e, 32'h42991cac} /* (11, 13, 3) {real, imag} */,
  {32'h42f030d4, 32'h43382e04} /* (11, 13, 2) {real, imag} */,
  {32'hc2d17b5a, 32'hc2df6a92} /* (11, 13, 1) {real, imag} */,
  {32'h440a20f4, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'h411b03c4, 32'h428ca0a3} /* (11, 12, 15) {real, imag} */,
  {32'hc20c7f56, 32'h43064659} /* (11, 12, 14) {real, imag} */,
  {32'h432c8bbe, 32'h42b1b1df} /* (11, 12, 13) {real, imag} */,
  {32'h43436cb5, 32'hc30ccb6b} /* (11, 12, 12) {real, imag} */,
  {32'h428a88dd, 32'h42ddee02} /* (11, 12, 11) {real, imag} */,
  {32'hc2cdc6b1, 32'hc011d510} /* (11, 12, 10) {real, imag} */,
  {32'hc201d62e, 32'h41a0401e} /* (11, 12, 9) {real, imag} */,
  {32'h424388ce, 32'h00000000} /* (11, 12, 8) {real, imag} */,
  {32'hc201d62e, 32'hc1a0401e} /* (11, 12, 7) {real, imag} */,
  {32'hc2cdc6b1, 32'h4011d510} /* (11, 12, 6) {real, imag} */,
  {32'h428a88dd, 32'hc2ddee02} /* (11, 12, 5) {real, imag} */,
  {32'h43436cb5, 32'h430ccb6b} /* (11, 12, 4) {real, imag} */,
  {32'h432c8bbe, 32'hc2b1b1df} /* (11, 12, 3) {real, imag} */,
  {32'hc20c7f56, 32'hc3064659} /* (11, 12, 2) {real, imag} */,
  {32'h411b03c4, 32'hc28ca0a3} /* (11, 12, 1) {real, imag} */,
  {32'h4407cf0f, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'h4224988a, 32'h4302dc20} /* (11, 11, 15) {real, imag} */,
  {32'h41b3e906, 32'h40a85290} /* (11, 11, 14) {real, imag} */,
  {32'h431ff28b, 32'h431617c0} /* (11, 11, 13) {real, imag} */,
  {32'hc15722c6, 32'h41f81742} /* (11, 11, 12) {real, imag} */,
  {32'h4132cf8e, 32'h41553b7c} /* (11, 11, 11) {real, imag} */,
  {32'h4211d546, 32'h4154b431} /* (11, 11, 10) {real, imag} */,
  {32'h40858668, 32'hc288d7b7} /* (11, 11, 9) {real, imag} */,
  {32'hc2a43efe, 32'h00000000} /* (11, 11, 8) {real, imag} */,
  {32'h40858668, 32'h4288d7b7} /* (11, 11, 7) {real, imag} */,
  {32'h4211d546, 32'hc154b431} /* (11, 11, 6) {real, imag} */,
  {32'h4132cf8e, 32'hc1553b7c} /* (11, 11, 5) {real, imag} */,
  {32'hc15722c6, 32'hc1f81742} /* (11, 11, 4) {real, imag} */,
  {32'h431ff28b, 32'hc31617c0} /* (11, 11, 3) {real, imag} */,
  {32'h41b3e906, 32'hc0a85290} /* (11, 11, 2) {real, imag} */,
  {32'h4224988a, 32'hc302dc20} /* (11, 11, 1) {real, imag} */,
  {32'h441e70b3, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'hc19d66b0, 32'h4342a3f1} /* (11, 10, 15) {real, imag} */,
  {32'h428a4cbf, 32'hc20923f9} /* (11, 10, 14) {real, imag} */,
  {32'hc04dc3c0, 32'h429dc72e} /* (11, 10, 13) {real, imag} */,
  {32'h41a0df0c, 32'h40fe5730} /* (11, 10, 12) {real, imag} */,
  {32'hc29d03e0, 32'h431c4da8} /* (11, 10, 11) {real, imag} */,
  {32'hc3086f35, 32'hc27aa5e9} /* (11, 10, 10) {real, imag} */,
  {32'h43015f52, 32'h42e1ea8e} /* (11, 10, 9) {real, imag} */,
  {32'hc24f69de, 32'h00000000} /* (11, 10, 8) {real, imag} */,
  {32'h43015f52, 32'hc2e1ea8e} /* (11, 10, 7) {real, imag} */,
  {32'hc3086f35, 32'h427aa5e9} /* (11, 10, 6) {real, imag} */,
  {32'hc29d03e0, 32'hc31c4da8} /* (11, 10, 5) {real, imag} */,
  {32'h41a0df0c, 32'hc0fe5730} /* (11, 10, 4) {real, imag} */,
  {32'hc04dc3c0, 32'hc29dc72e} /* (11, 10, 3) {real, imag} */,
  {32'h428a4cbf, 32'h420923f9} /* (11, 10, 2) {real, imag} */,
  {32'hc19d66b0, 32'hc342a3f1} /* (11, 10, 1) {real, imag} */,
  {32'h44457b80, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h41682786, 32'hc2d2d0da} /* (11, 9, 15) {real, imag} */,
  {32'h430362e6, 32'h432610ef} /* (11, 9, 14) {real, imag} */,
  {32'h41db3671, 32'h42d450b6} /* (11, 9, 13) {real, imag} */,
  {32'h42883f9a, 32'hc30d3e74} /* (11, 9, 12) {real, imag} */,
  {32'hc231b5ea, 32'h4315340c} /* (11, 9, 11) {real, imag} */,
  {32'hc2ee642f, 32'h41cd8618} /* (11, 9, 10) {real, imag} */,
  {32'hc25e186f, 32'h42251761} /* (11, 9, 9) {real, imag} */,
  {32'hc291508c, 32'h00000000} /* (11, 9, 8) {real, imag} */,
  {32'hc25e186f, 32'hc2251761} /* (11, 9, 7) {real, imag} */,
  {32'hc2ee642f, 32'hc1cd8618} /* (11, 9, 6) {real, imag} */,
  {32'hc231b5ea, 32'hc315340c} /* (11, 9, 5) {real, imag} */,
  {32'h42883f9a, 32'h430d3e74} /* (11, 9, 4) {real, imag} */,
  {32'h41db3671, 32'hc2d450b6} /* (11, 9, 3) {real, imag} */,
  {32'h430362e6, 32'hc32610ef} /* (11, 9, 2) {real, imag} */,
  {32'h41682786, 32'h42d2d0da} /* (11, 9, 1) {real, imag} */,
  {32'h43dd28ac, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h42cbbad9, 32'hc33127e4} /* (11, 8, 15) {real, imag} */,
  {32'h43126d6c, 32'hc218383e} /* (11, 8, 14) {real, imag} */,
  {32'h429eb42e, 32'hc31b6299} /* (11, 8, 13) {real, imag} */,
  {32'hc285dd3e, 32'h426d0b24} /* (11, 8, 12) {real, imag} */,
  {32'hc2af06aa, 32'h42ce37ec} /* (11, 8, 11) {real, imag} */,
  {32'hc1954f3a, 32'h41d2f756} /* (11, 8, 10) {real, imag} */,
  {32'h4206e3de, 32'hc2c138d5} /* (11, 8, 9) {real, imag} */,
  {32'hc31c57d1, 32'h00000000} /* (11, 8, 8) {real, imag} */,
  {32'h4206e3de, 32'h42c138d5} /* (11, 8, 7) {real, imag} */,
  {32'hc1954f3a, 32'hc1d2f756} /* (11, 8, 6) {real, imag} */,
  {32'hc2af06aa, 32'hc2ce37ec} /* (11, 8, 5) {real, imag} */,
  {32'hc285dd3e, 32'hc26d0b24} /* (11, 8, 4) {real, imag} */,
  {32'h429eb42e, 32'h431b6299} /* (11, 8, 3) {real, imag} */,
  {32'h43126d6c, 32'h4218383e} /* (11, 8, 2) {real, imag} */,
  {32'h42cbbad9, 32'h433127e4} /* (11, 8, 1) {real, imag} */,
  {32'h42cc74ee, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h3fb172f0, 32'hbf9a0300} /* (11, 7, 15) {real, imag} */,
  {32'h42aff3e8, 32'h42b20e78} /* (11, 7, 14) {real, imag} */,
  {32'h426d10fe, 32'hc25fcbe8} /* (11, 7, 13) {real, imag} */,
  {32'hc26d5eb8, 32'hc37bbbec} /* (11, 7, 12) {real, imag} */,
  {32'hc2e81be5, 32'hc172a7a8} /* (11, 7, 11) {real, imag} */,
  {32'hc24cfbda, 32'h4311418d} /* (11, 7, 10) {real, imag} */,
  {32'h4295f098, 32'h429f5758} /* (11, 7, 9) {real, imag} */,
  {32'h42a2f7c8, 32'h00000000} /* (11, 7, 8) {real, imag} */,
  {32'h4295f098, 32'hc29f5758} /* (11, 7, 7) {real, imag} */,
  {32'hc24cfbda, 32'hc311418d} /* (11, 7, 6) {real, imag} */,
  {32'hc2e81be5, 32'h4172a7a8} /* (11, 7, 5) {real, imag} */,
  {32'hc26d5eb8, 32'h437bbbec} /* (11, 7, 4) {real, imag} */,
  {32'h426d10fe, 32'h425fcbe8} /* (11, 7, 3) {real, imag} */,
  {32'h42aff3e8, 32'hc2b20e78} /* (11, 7, 2) {real, imag} */,
  {32'h3fb172f0, 32'h3f9a0300} /* (11, 7, 1) {real, imag} */,
  {32'h42fdadea, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'hc37911e2, 32'hc21f4fac} /* (11, 6, 15) {real, imag} */,
  {32'h42d6b465, 32'hc2f375ae} /* (11, 6, 14) {real, imag} */,
  {32'hc3398bf8, 32'h42be171e} /* (11, 6, 13) {real, imag} */,
  {32'hc019b0c0, 32'hc30db610} /* (11, 6, 12) {real, imag} */,
  {32'h4317c50c, 32'hc2fd1959} /* (11, 6, 11) {real, imag} */,
  {32'h42ab34c8, 32'h42b43768} /* (11, 6, 10) {real, imag} */,
  {32'h430f2982, 32'hc202181d} /* (11, 6, 9) {real, imag} */,
  {32'hc336bd40, 32'h00000000} /* (11, 6, 8) {real, imag} */,
  {32'h430f2982, 32'h4202181d} /* (11, 6, 7) {real, imag} */,
  {32'h42ab34c8, 32'hc2b43768} /* (11, 6, 6) {real, imag} */,
  {32'h4317c50c, 32'h42fd1959} /* (11, 6, 5) {real, imag} */,
  {32'hc019b0c0, 32'h430db610} /* (11, 6, 4) {real, imag} */,
  {32'hc3398bf8, 32'hc2be171e} /* (11, 6, 3) {real, imag} */,
  {32'h42d6b465, 32'h42f375ae} /* (11, 6, 2) {real, imag} */,
  {32'hc37911e2, 32'h421f4fac} /* (11, 6, 1) {real, imag} */,
  {32'h43ad9bd4, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'hc2d9a355, 32'h43808d98} /* (11, 5, 15) {real, imag} */,
  {32'h4313b7f2, 32'hc26433e6} /* (11, 5, 14) {real, imag} */,
  {32'hc33f8953, 32'hc2069278} /* (11, 5, 13) {real, imag} */,
  {32'h428c1e69, 32'hc1f083a6} /* (11, 5, 12) {real, imag} */,
  {32'h4239665e, 32'h41a400de} /* (11, 5, 11) {real, imag} */,
  {32'hc30c5308, 32'h41c7210c} /* (11, 5, 10) {real, imag} */,
  {32'h42d096a0, 32'hc2aaaa4f} /* (11, 5, 9) {real, imag} */,
  {32'hc19b7f70, 32'h00000000} /* (11, 5, 8) {real, imag} */,
  {32'h42d096a0, 32'h42aaaa4f} /* (11, 5, 7) {real, imag} */,
  {32'hc30c5308, 32'hc1c7210c} /* (11, 5, 6) {real, imag} */,
  {32'h4239665e, 32'hc1a400de} /* (11, 5, 5) {real, imag} */,
  {32'h428c1e69, 32'h41f083a6} /* (11, 5, 4) {real, imag} */,
  {32'hc33f8953, 32'h42069278} /* (11, 5, 3) {real, imag} */,
  {32'h4313b7f2, 32'h426433e6} /* (11, 5, 2) {real, imag} */,
  {32'hc2d9a355, 32'hc3808d98} /* (11, 5, 1) {real, imag} */,
  {32'h43eb17d7, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h4297bd20, 32'h438d7cdb} /* (11, 4, 15) {real, imag} */,
  {32'h42fea8dd, 32'hc23bc81b} /* (11, 4, 14) {real, imag} */,
  {32'hc2df901c, 32'hc294af1d} /* (11, 4, 13) {real, imag} */,
  {32'hc0553c80, 32'hc2e2941c} /* (11, 4, 12) {real, imag} */,
  {32'h408abfd0, 32'h4290b186} /* (11, 4, 11) {real, imag} */,
  {32'hc286419f, 32'h42dd1fec} /* (11, 4, 10) {real, imag} */,
  {32'h400acbd8, 32'h41c5640e} /* (11, 4, 9) {real, imag} */,
  {32'hbfb3b780, 32'h00000000} /* (11, 4, 8) {real, imag} */,
  {32'h400acbd8, 32'hc1c5640e} /* (11, 4, 7) {real, imag} */,
  {32'hc286419f, 32'hc2dd1fec} /* (11, 4, 6) {real, imag} */,
  {32'h408abfd0, 32'hc290b186} /* (11, 4, 5) {real, imag} */,
  {32'hc0553c80, 32'h42e2941c} /* (11, 4, 4) {real, imag} */,
  {32'hc2df901c, 32'h4294af1d} /* (11, 4, 3) {real, imag} */,
  {32'h42fea8dd, 32'h423bc81b} /* (11, 4, 2) {real, imag} */,
  {32'h4297bd20, 32'hc38d7cdb} /* (11, 4, 1) {real, imag} */,
  {32'h43a09bf9, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h42af3be4, 32'h4342fddb} /* (11, 3, 15) {real, imag} */,
  {32'h3e871180, 32'h425accce} /* (11, 3, 14) {real, imag} */,
  {32'hc289ab32, 32'h42303351} /* (11, 3, 13) {real, imag} */,
  {32'hc24f3e0c, 32'hc3525aec} /* (11, 3, 12) {real, imag} */,
  {32'h3e8d9840, 32'hc2a2ab04} /* (11, 3, 11) {real, imag} */,
  {32'h430e6967, 32'hc08ca310} /* (11, 3, 10) {real, imag} */,
  {32'h40bc4d60, 32'h425f8f3d} /* (11, 3, 9) {real, imag} */,
  {32'hc2b26a3a, 32'h00000000} /* (11, 3, 8) {real, imag} */,
  {32'h40bc4d60, 32'hc25f8f3d} /* (11, 3, 7) {real, imag} */,
  {32'h430e6967, 32'h408ca310} /* (11, 3, 6) {real, imag} */,
  {32'h3e8d9840, 32'h42a2ab04} /* (11, 3, 5) {real, imag} */,
  {32'hc24f3e0c, 32'h43525aec} /* (11, 3, 4) {real, imag} */,
  {32'hc289ab32, 32'hc2303351} /* (11, 3, 3) {real, imag} */,
  {32'h3e871180, 32'hc25accce} /* (11, 3, 2) {real, imag} */,
  {32'h42af3be4, 32'hc342fddb} /* (11, 3, 1) {real, imag} */,
  {32'hc10f34e0, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'hc2f6510e, 32'hc2aab01e} /* (11, 2, 15) {real, imag} */,
  {32'h409815e0, 32'h426f525c} /* (11, 2, 14) {real, imag} */,
  {32'h4300f850, 32'h42a8cd22} /* (11, 2, 13) {real, imag} */,
  {32'h424e5b83, 32'hc3233db5} /* (11, 2, 12) {real, imag} */,
  {32'h42987150, 32'h41e5a4d4} /* (11, 2, 11) {real, imag} */,
  {32'h4249ff20, 32'h42745179} /* (11, 2, 10) {real, imag} */,
  {32'hc2ca17f5, 32'hc2c0c27c} /* (11, 2, 9) {real, imag} */,
  {32'hc2573e2a, 32'h00000000} /* (11, 2, 8) {real, imag} */,
  {32'hc2ca17f5, 32'h42c0c27c} /* (11, 2, 7) {real, imag} */,
  {32'h4249ff20, 32'hc2745179} /* (11, 2, 6) {real, imag} */,
  {32'h42987150, 32'hc1e5a4d4} /* (11, 2, 5) {real, imag} */,
  {32'h424e5b83, 32'h43233db5} /* (11, 2, 4) {real, imag} */,
  {32'h4300f850, 32'hc2a8cd22} /* (11, 2, 3) {real, imag} */,
  {32'h409815e0, 32'hc26f525c} /* (11, 2, 2) {real, imag} */,
  {32'hc2f6510e, 32'h42aab01e} /* (11, 2, 1) {real, imag} */,
  {32'hc30dada9, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'hc294857e, 32'h41219eb8} /* (11, 1, 15) {real, imag} */,
  {32'h40f36380, 32'hc283846b} /* (11, 1, 14) {real, imag} */,
  {32'h41806490, 32'hc2b8961f} /* (11, 1, 13) {real, imag} */,
  {32'h41551330, 32'hc16f8146} /* (11, 1, 12) {real, imag} */,
  {32'h42a1dc6d, 32'h430c0384} /* (11, 1, 11) {real, imag} */,
  {32'hc287164b, 32'hc2843c32} /* (11, 1, 10) {real, imag} */,
  {32'hc11d5ca4, 32'hc035e02c} /* (11, 1, 9) {real, imag} */,
  {32'h40fd3470, 32'h00000000} /* (11, 1, 8) {real, imag} */,
  {32'hc11d5ca4, 32'h4035e02c} /* (11, 1, 7) {real, imag} */,
  {32'hc287164b, 32'h42843c32} /* (11, 1, 6) {real, imag} */,
  {32'h42a1dc6d, 32'hc30c0384} /* (11, 1, 5) {real, imag} */,
  {32'h41551330, 32'h416f8146} /* (11, 1, 4) {real, imag} */,
  {32'h41806490, 32'h42b8961f} /* (11, 1, 3) {real, imag} */,
  {32'h40f36380, 32'h4283846b} /* (11, 1, 2) {real, imag} */,
  {32'hc294857e, 32'hc1219eb8} /* (11, 1, 1) {real, imag} */,
  {32'h438ec7bf, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h42a95ca3, 32'h42cadcf9} /* (11, 0, 15) {real, imag} */,
  {32'h425d9892, 32'h42347ac8} /* (11, 0, 14) {real, imag} */,
  {32'hc246763c, 32'hc196ab40} /* (11, 0, 13) {real, imag} */,
  {32'h4079ee90, 32'hc1eeb420} /* (11, 0, 12) {real, imag} */,
  {32'h422c6d9c, 32'h42a1f954} /* (11, 0, 11) {real, imag} */,
  {32'hc236874d, 32'hc2ba48fc} /* (11, 0, 10) {real, imag} */,
  {32'h42a0f345, 32'hc25691b6} /* (11, 0, 9) {real, imag} */,
  {32'h42afe592, 32'h00000000} /* (11, 0, 8) {real, imag} */,
  {32'h42a0f345, 32'h425691b6} /* (11, 0, 7) {real, imag} */,
  {32'hc236874d, 32'h42ba48fc} /* (11, 0, 6) {real, imag} */,
  {32'h422c6d9c, 32'hc2a1f954} /* (11, 0, 5) {real, imag} */,
  {32'h4079ee90, 32'h41eeb420} /* (11, 0, 4) {real, imag} */,
  {32'hc246763c, 32'h4196ab40} /* (11, 0, 3) {real, imag} */,
  {32'h425d9892, 32'hc2347ac8} /* (11, 0, 2) {real, imag} */,
  {32'h42a95ca3, 32'hc2cadcf9} /* (11, 0, 1) {real, imag} */,
  {32'h431f0acb, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h41cfe2c8, 32'hc1821ef0} /* (10, 15, 15) {real, imag} */,
  {32'hc225d269, 32'hc2ed1ac6} /* (10, 15, 14) {real, imag} */,
  {32'h43048968, 32'h42addd42} /* (10, 15, 13) {real, imag} */,
  {32'hc2a9f629, 32'h42088974} /* (10, 15, 12) {real, imag} */,
  {32'hc1c02c36, 32'h41d0d7fc} /* (10, 15, 11) {real, imag} */,
  {32'hc27c8797, 32'hc2ac341f} /* (10, 15, 10) {real, imag} */,
  {32'h42254be7, 32'hc21f88c6} /* (10, 15, 9) {real, imag} */,
  {32'h40abf804, 32'h00000000} /* (10, 15, 8) {real, imag} */,
  {32'h42254be7, 32'h421f88c6} /* (10, 15, 7) {real, imag} */,
  {32'hc27c8797, 32'h42ac341f} /* (10, 15, 6) {real, imag} */,
  {32'hc1c02c36, 32'hc1d0d7fc} /* (10, 15, 5) {real, imag} */,
  {32'hc2a9f629, 32'hc2088974} /* (10, 15, 4) {real, imag} */,
  {32'h43048968, 32'hc2addd42} /* (10, 15, 3) {real, imag} */,
  {32'hc225d269, 32'h42ed1ac6} /* (10, 15, 2) {real, imag} */,
  {32'h41cfe2c8, 32'h41821ef0} /* (10, 15, 1) {real, imag} */,
  {32'h436d125c, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'h429597a6, 32'hc2fbdd64} /* (10, 14, 15) {real, imag} */,
  {32'hc30a62ba, 32'hc3c8ef5a} /* (10, 14, 14) {real, imag} */,
  {32'h4304480c, 32'h42226d9f} /* (10, 14, 13) {real, imag} */,
  {32'hc13a1ab0, 32'h422978e3} /* (10, 14, 12) {real, imag} */,
  {32'hc209b3f3, 32'h430cb4b6} /* (10, 14, 11) {real, imag} */,
  {32'hc21a90bc, 32'hc20cb1ca} /* (10, 14, 10) {real, imag} */,
  {32'hc1ea1ae0, 32'h41ea7002} /* (10, 14, 9) {real, imag} */,
  {32'hc1a2f20a, 32'h00000000} /* (10, 14, 8) {real, imag} */,
  {32'hc1ea1ae0, 32'hc1ea7002} /* (10, 14, 7) {real, imag} */,
  {32'hc21a90bc, 32'h420cb1ca} /* (10, 14, 6) {real, imag} */,
  {32'hc209b3f3, 32'hc30cb4b6} /* (10, 14, 5) {real, imag} */,
  {32'hc13a1ab0, 32'hc22978e3} /* (10, 14, 4) {real, imag} */,
  {32'h4304480c, 32'hc2226d9f} /* (10, 14, 3) {real, imag} */,
  {32'hc30a62ba, 32'h43c8ef5a} /* (10, 14, 2) {real, imag} */,
  {32'h429597a6, 32'h42fbdd64} /* (10, 14, 1) {real, imag} */,
  {32'h43c6aabf, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'h417bcc28, 32'hc20a4ec4} /* (10, 13, 15) {real, imag} */,
  {32'hc20d939a, 32'hc32274b0} /* (10, 13, 14) {real, imag} */,
  {32'h42ad5b31, 32'h42d393f6} /* (10, 13, 13) {real, imag} */,
  {32'hc2d49830, 32'hc2c4fc12} /* (10, 13, 12) {real, imag} */,
  {32'h413d23f4, 32'h42904d3c} /* (10, 13, 11) {real, imag} */,
  {32'h419e0ff6, 32'h43363316} /* (10, 13, 10) {real, imag} */,
  {32'hc2592e15, 32'h42a90868} /* (10, 13, 9) {real, imag} */,
  {32'hc20461c7, 32'h00000000} /* (10, 13, 8) {real, imag} */,
  {32'hc2592e15, 32'hc2a90868} /* (10, 13, 7) {real, imag} */,
  {32'h419e0ff6, 32'hc3363316} /* (10, 13, 6) {real, imag} */,
  {32'h413d23f4, 32'hc2904d3c} /* (10, 13, 5) {real, imag} */,
  {32'hc2d49830, 32'h42c4fc12} /* (10, 13, 4) {real, imag} */,
  {32'h42ad5b31, 32'hc2d393f6} /* (10, 13, 3) {real, imag} */,
  {32'hc20d939a, 32'h432274b0} /* (10, 13, 2) {real, imag} */,
  {32'h417bcc28, 32'h420a4ec4} /* (10, 13, 1) {real, imag} */,
  {32'h44253840, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'hc335089c, 32'h43937f72} /* (10, 12, 15) {real, imag} */,
  {32'h437cc0ee, 32'hc2bb638e} /* (10, 12, 14) {real, imag} */,
  {32'h42675d9d, 32'h4281a04c} /* (10, 12, 13) {real, imag} */,
  {32'h3e0e7f00, 32'h4232d2a4} /* (10, 12, 12) {real, imag} */,
  {32'hbf7aa580, 32'hc21ada88} /* (10, 12, 11) {real, imag} */,
  {32'hc2400440, 32'h42dc14b6} /* (10, 12, 10) {real, imag} */,
  {32'h3f971500, 32'hc2cc6da2} /* (10, 12, 9) {real, imag} */,
  {32'hc23d82d1, 32'h00000000} /* (10, 12, 8) {real, imag} */,
  {32'h3f971500, 32'h42cc6da2} /* (10, 12, 7) {real, imag} */,
  {32'hc2400440, 32'hc2dc14b6} /* (10, 12, 6) {real, imag} */,
  {32'hbf7aa580, 32'h421ada88} /* (10, 12, 5) {real, imag} */,
  {32'h3e0e7f00, 32'hc232d2a4} /* (10, 12, 4) {real, imag} */,
  {32'h42675d9d, 32'hc281a04c} /* (10, 12, 3) {real, imag} */,
  {32'h437cc0ee, 32'h42bb638e} /* (10, 12, 2) {real, imag} */,
  {32'hc335089c, 32'hc3937f72} /* (10, 12, 1) {real, imag} */,
  {32'h44070dac, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hc39b2350, 32'h4374d370} /* (10, 11, 15) {real, imag} */,
  {32'h4219f7b8, 32'h40b0b1a0} /* (10, 11, 14) {real, imag} */,
  {32'hc2076430, 32'hc300a952} /* (10, 11, 13) {real, imag} */,
  {32'h42a8c034, 32'h42f6d2ae} /* (10, 11, 12) {real, imag} */,
  {32'h422e24c7, 32'hc240cb6c} /* (10, 11, 11) {real, imag} */,
  {32'hc1d24e5e, 32'h42ccf8dd} /* (10, 11, 10) {real, imag} */,
  {32'h431272c6, 32'hc1cf96a9} /* (10, 11, 9) {real, imag} */,
  {32'h4184d5ea, 32'h00000000} /* (10, 11, 8) {real, imag} */,
  {32'h431272c6, 32'h41cf96a9} /* (10, 11, 7) {real, imag} */,
  {32'hc1d24e5e, 32'hc2ccf8dd} /* (10, 11, 6) {real, imag} */,
  {32'h422e24c7, 32'h4240cb6c} /* (10, 11, 5) {real, imag} */,
  {32'h42a8c034, 32'hc2f6d2ae} /* (10, 11, 4) {real, imag} */,
  {32'hc2076430, 32'h4300a952} /* (10, 11, 3) {real, imag} */,
  {32'h4219f7b8, 32'hc0b0b1a0} /* (10, 11, 2) {real, imag} */,
  {32'hc39b2350, 32'hc374d370} /* (10, 11, 1) {real, imag} */,
  {32'h44394c9f, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h41b5b482, 32'h438b24cc} /* (10, 10, 15) {real, imag} */,
  {32'h42c8ac66, 32'hc2811566} /* (10, 10, 14) {real, imag} */,
  {32'hc2c7cbc2, 32'h41eb0ec2} /* (10, 10, 13) {real, imag} */,
  {32'h41a39438, 32'h41cbebf0} /* (10, 10, 12) {real, imag} */,
  {32'hc2fcd62a, 32'hbec0aa00} /* (10, 10, 11) {real, imag} */,
  {32'hc2f8f90a, 32'hc1a10aac} /* (10, 10, 10) {real, imag} */,
  {32'h42268040, 32'h424910a8} /* (10, 10, 9) {real, imag} */,
  {32'h42b9cecc, 32'h00000000} /* (10, 10, 8) {real, imag} */,
  {32'h42268040, 32'hc24910a8} /* (10, 10, 7) {real, imag} */,
  {32'hc2f8f90a, 32'h41a10aac} /* (10, 10, 6) {real, imag} */,
  {32'hc2fcd62a, 32'h3ec0aa00} /* (10, 10, 5) {real, imag} */,
  {32'h41a39438, 32'hc1cbebf0} /* (10, 10, 4) {real, imag} */,
  {32'hc2c7cbc2, 32'hc1eb0ec2} /* (10, 10, 3) {real, imag} */,
  {32'h42c8ac66, 32'h42811566} /* (10, 10, 2) {real, imag} */,
  {32'h41b5b482, 32'hc38b24cc} /* (10, 10, 1) {real, imag} */,
  {32'h444fea53, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h434ad12d, 32'hc245b980} /* (10, 9, 15) {real, imag} */,
  {32'h4387ecb1, 32'h42e41e2b} /* (10, 9, 14) {real, imag} */,
  {32'hc3123c30, 32'h41c6077a} /* (10, 9, 13) {real, imag} */,
  {32'hc201f691, 32'hc20fe2e0} /* (10, 9, 12) {real, imag} */,
  {32'h4213c5fb, 32'h42a3a37c} /* (10, 9, 11) {real, imag} */,
  {32'h4084a798, 32'hc1b4382c} /* (10, 9, 10) {real, imag} */,
  {32'h42c8a86c, 32'h421edbc4} /* (10, 9, 9) {real, imag} */,
  {32'h40e30714, 32'h00000000} /* (10, 9, 8) {real, imag} */,
  {32'h42c8a86c, 32'hc21edbc4} /* (10, 9, 7) {real, imag} */,
  {32'h4084a798, 32'h41b4382c} /* (10, 9, 6) {real, imag} */,
  {32'h4213c5fb, 32'hc2a3a37c} /* (10, 9, 5) {real, imag} */,
  {32'hc201f691, 32'h420fe2e0} /* (10, 9, 4) {real, imag} */,
  {32'hc3123c30, 32'hc1c6077a} /* (10, 9, 3) {real, imag} */,
  {32'h4387ecb1, 32'hc2e41e2b} /* (10, 9, 2) {real, imag} */,
  {32'h434ad12d, 32'h4245b980} /* (10, 9, 1) {real, imag} */,
  {32'h440837fb, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'hc1296870, 32'hc37605da} /* (10, 8, 15) {real, imag} */,
  {32'h4317ecde, 32'hc213648f} /* (10, 8, 14) {real, imag} */,
  {32'hc3432b4c, 32'hc2a6bd02} /* (10, 8, 13) {real, imag} */,
  {32'h41cd0db3, 32'hc18c92dc} /* (10, 8, 12) {real, imag} */,
  {32'hc2c5a232, 32'h42b727ac} /* (10, 8, 11) {real, imag} */,
  {32'hc2a591bd, 32'hc22a6eca} /* (10, 8, 10) {real, imag} */,
  {32'hc11c7751, 32'hc2b18f55} /* (10, 8, 9) {real, imag} */,
  {32'hc31b826b, 32'h00000000} /* (10, 8, 8) {real, imag} */,
  {32'hc11c7751, 32'h42b18f55} /* (10, 8, 7) {real, imag} */,
  {32'hc2a591bd, 32'h422a6eca} /* (10, 8, 6) {real, imag} */,
  {32'hc2c5a232, 32'hc2b727ac} /* (10, 8, 5) {real, imag} */,
  {32'h41cd0db3, 32'h418c92dc} /* (10, 8, 4) {real, imag} */,
  {32'hc3432b4c, 32'h42a6bd02} /* (10, 8, 3) {real, imag} */,
  {32'h4317ecde, 32'h4213648f} /* (10, 8, 2) {real, imag} */,
  {32'hc1296870, 32'h437605da} /* (10, 8, 1) {real, imag} */,
  {32'h43bda29b, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h43230091, 32'hc23e7748} /* (10, 7, 15) {real, imag} */,
  {32'hc2693ea8, 32'hc33443c2} /* (10, 7, 14) {real, imag} */,
  {32'hc35c0892, 32'hc307560b} /* (10, 7, 13) {real, imag} */,
  {32'hc28a58d4, 32'hc336c66d} /* (10, 7, 12) {real, imag} */,
  {32'hc27b112b, 32'h42f3f796} /* (10, 7, 11) {real, imag} */,
  {32'h4120ac40, 32'hc2d2cacf} /* (10, 7, 10) {real, imag} */,
  {32'h42d249d2, 32'hc1942591} /* (10, 7, 9) {real, imag} */,
  {32'hc213ea6a, 32'h00000000} /* (10, 7, 8) {real, imag} */,
  {32'h42d249d2, 32'h41942591} /* (10, 7, 7) {real, imag} */,
  {32'h4120ac40, 32'h42d2cacf} /* (10, 7, 6) {real, imag} */,
  {32'hc27b112b, 32'hc2f3f796} /* (10, 7, 5) {real, imag} */,
  {32'hc28a58d4, 32'h4336c66d} /* (10, 7, 4) {real, imag} */,
  {32'hc35c0892, 32'h4307560b} /* (10, 7, 3) {real, imag} */,
  {32'hc2693ea8, 32'h433443c2} /* (10, 7, 2) {real, imag} */,
  {32'h43230091, 32'h423e7748} /* (10, 7, 1) {real, imag} */,
  {32'h43af449b, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h401bd350, 32'h41865728} /* (10, 6, 15) {real, imag} */,
  {32'hc3010777, 32'hc32e0989} /* (10, 6, 14) {real, imag} */,
  {32'h41acfa34, 32'hc30693f3} /* (10, 6, 13) {real, imag} */,
  {32'h42fe885a, 32'h4176dca8} /* (10, 6, 12) {real, imag} */,
  {32'h42d9cf8a, 32'hc2f7fb80} /* (10, 6, 11) {real, imag} */,
  {32'hc27c89d3, 32'h41ab59ac} /* (10, 6, 10) {real, imag} */,
  {32'hc08a06d0, 32'h419d0c67} /* (10, 6, 9) {real, imag} */,
  {32'h4313b319, 32'h00000000} /* (10, 6, 8) {real, imag} */,
  {32'hc08a06d0, 32'hc19d0c67} /* (10, 6, 7) {real, imag} */,
  {32'hc27c89d3, 32'hc1ab59ac} /* (10, 6, 6) {real, imag} */,
  {32'h42d9cf8a, 32'h42f7fb80} /* (10, 6, 5) {real, imag} */,
  {32'h42fe885a, 32'hc176dca8} /* (10, 6, 4) {real, imag} */,
  {32'h41acfa34, 32'h430693f3} /* (10, 6, 3) {real, imag} */,
  {32'hc3010777, 32'h432e0989} /* (10, 6, 2) {real, imag} */,
  {32'h401bd350, 32'hc1865728} /* (10, 6, 1) {real, imag} */,
  {32'h4393e71e, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'hc2ac8a9a, 32'h4337b72e} /* (10, 5, 15) {real, imag} */,
  {32'hc27fedd4, 32'hc3977f30} /* (10, 5, 14) {real, imag} */,
  {32'h42b84b46, 32'hc2bbdb18} /* (10, 5, 13) {real, imag} */,
  {32'h42bca8dc, 32'h421a3148} /* (10, 5, 12) {real, imag} */,
  {32'hc2f64142, 32'hc0ee3324} /* (10, 5, 11) {real, imag} */,
  {32'h4133ca5c, 32'h41f15794} /* (10, 5, 10) {real, imag} */,
  {32'h42bb05cf, 32'hc1b59fbb} /* (10, 5, 9) {real, imag} */,
  {32'hc2c3e318, 32'h00000000} /* (10, 5, 8) {real, imag} */,
  {32'h42bb05cf, 32'h41b59fbb} /* (10, 5, 7) {real, imag} */,
  {32'h4133ca5c, 32'hc1f15794} /* (10, 5, 6) {real, imag} */,
  {32'hc2f64142, 32'h40ee3324} /* (10, 5, 5) {real, imag} */,
  {32'h42bca8dc, 32'hc21a3148} /* (10, 5, 4) {real, imag} */,
  {32'h42b84b46, 32'h42bbdb18} /* (10, 5, 3) {real, imag} */,
  {32'hc27fedd4, 32'h43977f30} /* (10, 5, 2) {real, imag} */,
  {32'hc2ac8a9a, 32'hc337b72e} /* (10, 5, 1) {real, imag} */,
  {32'h42c43f40, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h43058f58, 32'h439a1054} /* (10, 4, 15) {real, imag} */,
  {32'h41dd3d10, 32'hc22d2e74} /* (10, 4, 14) {real, imag} */,
  {32'h4145616c, 32'hbea09780} /* (10, 4, 13) {real, imag} */,
  {32'hc264f577, 32'hbeac4d40} /* (10, 4, 12) {real, imag} */,
  {32'hc20053e7, 32'hc19e4540} /* (10, 4, 11) {real, imag} */,
  {32'h4326020c, 32'h4278be4c} /* (10, 4, 10) {real, imag} */,
  {32'h413a77e0, 32'hc29964a2} /* (10, 4, 9) {real, imag} */,
  {32'hbfba7260, 32'h00000000} /* (10, 4, 8) {real, imag} */,
  {32'h413a77e0, 32'h429964a2} /* (10, 4, 7) {real, imag} */,
  {32'h4326020c, 32'hc278be4c} /* (10, 4, 6) {real, imag} */,
  {32'hc20053e7, 32'h419e4540} /* (10, 4, 5) {real, imag} */,
  {32'hc264f577, 32'h3eac4d40} /* (10, 4, 4) {real, imag} */,
  {32'h4145616c, 32'h3ea09780} /* (10, 4, 3) {real, imag} */,
  {32'h41dd3d10, 32'h422d2e74} /* (10, 4, 2) {real, imag} */,
  {32'h43058f58, 32'hc39a1054} /* (10, 4, 1) {real, imag} */,
  {32'h4314a8c0, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'hc2b7f41f, 32'h43963a3e} /* (10, 3, 15) {real, imag} */,
  {32'h424fa962, 32'h425ba20a} /* (10, 3, 14) {real, imag} */,
  {32'hc1374b58, 32'h408e0dd0} /* (10, 3, 13) {real, imag} */,
  {32'h41598d98, 32'h42406c98} /* (10, 3, 12) {real, imag} */,
  {32'h42bed080, 32'h4290b992} /* (10, 3, 11) {real, imag} */,
  {32'h430ab863, 32'hbf57c700} /* (10, 3, 10) {real, imag} */,
  {32'hc2e3a5fc, 32'hc205dd43} /* (10, 3, 9) {real, imag} */,
  {32'h42b36038, 32'h00000000} /* (10, 3, 8) {real, imag} */,
  {32'hc2e3a5fc, 32'h4205dd43} /* (10, 3, 7) {real, imag} */,
  {32'h430ab863, 32'h3f57c700} /* (10, 3, 6) {real, imag} */,
  {32'h42bed080, 32'hc290b992} /* (10, 3, 5) {real, imag} */,
  {32'h41598d98, 32'hc2406c98} /* (10, 3, 4) {real, imag} */,
  {32'hc1374b58, 32'hc08e0dd0} /* (10, 3, 3) {real, imag} */,
  {32'h424fa962, 32'hc25ba20a} /* (10, 3, 2) {real, imag} */,
  {32'hc2b7f41f, 32'hc3963a3e} /* (10, 3, 1) {real, imag} */,
  {32'h42a1fd38, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'hc383e760, 32'h432f8684} /* (10, 2, 15) {real, imag} */,
  {32'h40dc5a00, 32'hc1ecb268} /* (10, 2, 14) {real, imag} */,
  {32'h41eb1dde, 32'h4285af14} /* (10, 2, 13) {real, imag} */,
  {32'h42d06e12, 32'hc2d9154a} /* (10, 2, 12) {real, imag} */,
  {32'h420baa35, 32'h42709e9e} /* (10, 2, 11) {real, imag} */,
  {32'h42a4ee35, 32'hc316e1dc} /* (10, 2, 10) {real, imag} */,
  {32'h429ae71d, 32'hc1d1abb4} /* (10, 2, 9) {real, imag} */,
  {32'hbe930380, 32'h00000000} /* (10, 2, 8) {real, imag} */,
  {32'h429ae71d, 32'h41d1abb4} /* (10, 2, 7) {real, imag} */,
  {32'h42a4ee35, 32'h4316e1dc} /* (10, 2, 6) {real, imag} */,
  {32'h420baa35, 32'hc2709e9e} /* (10, 2, 5) {real, imag} */,
  {32'h42d06e12, 32'h42d9154a} /* (10, 2, 4) {real, imag} */,
  {32'h41eb1dde, 32'hc285af14} /* (10, 2, 3) {real, imag} */,
  {32'h40dc5a00, 32'h41ecb268} /* (10, 2, 2) {real, imag} */,
  {32'hc383e760, 32'hc32f8684} /* (10, 2, 1) {real, imag} */,
  {32'h41d9f190, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'hc1d6ebf8, 32'h42d6ab34} /* (10, 1, 15) {real, imag} */,
  {32'hbd669400, 32'h42620b58} /* (10, 1, 14) {real, imag} */,
  {32'h431b8876, 32'hc1b35a0a} /* (10, 1, 13) {real, imag} */,
  {32'h42af0d3b, 32'hc2a7c010} /* (10, 1, 12) {real, imag} */,
  {32'h42be9e68, 32'h431d04d8} /* (10, 1, 11) {real, imag} */,
  {32'hc158d884, 32'h42c752cd} /* (10, 1, 10) {real, imag} */,
  {32'hc26604cb, 32'hc281e60f} /* (10, 1, 9) {real, imag} */,
  {32'h422d7130, 32'h00000000} /* (10, 1, 8) {real, imag} */,
  {32'hc26604cb, 32'h4281e60f} /* (10, 1, 7) {real, imag} */,
  {32'hc158d884, 32'hc2c752cd} /* (10, 1, 6) {real, imag} */,
  {32'h42be9e68, 32'hc31d04d8} /* (10, 1, 5) {real, imag} */,
  {32'h42af0d3b, 32'h42a7c010} /* (10, 1, 4) {real, imag} */,
  {32'h431b8876, 32'h41b35a0a} /* (10, 1, 3) {real, imag} */,
  {32'hbd669400, 32'hc2620b58} /* (10, 1, 2) {real, imag} */,
  {32'hc1d6ebf8, 32'hc2d6ab34} /* (10, 1, 1) {real, imag} */,
  {32'h4399d5ae, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h42a1b5c4, 32'hc2b6b463} /* (10, 0, 15) {real, imag} */,
  {32'hc2a14bc1, 32'h41191404} /* (10, 0, 14) {real, imag} */,
  {32'h42d2376f, 32'hc1c99788} /* (10, 0, 13) {real, imag} */,
  {32'h424e5a76, 32'hc2c5b8c0} /* (10, 0, 12) {real, imag} */,
  {32'h42b8f4e2, 32'h42ea37d0} /* (10, 0, 11) {real, imag} */,
  {32'hc0e4ff70, 32'h420a0d68} /* (10, 0, 10) {real, imag} */,
  {32'hc13e429f, 32'h41b974ec} /* (10, 0, 9) {real, imag} */,
  {32'hc26cf317, 32'h00000000} /* (10, 0, 8) {real, imag} */,
  {32'hc13e429f, 32'hc1b974ec} /* (10, 0, 7) {real, imag} */,
  {32'hc0e4ff70, 32'hc20a0d68} /* (10, 0, 6) {real, imag} */,
  {32'h42b8f4e2, 32'hc2ea37d0} /* (10, 0, 5) {real, imag} */,
  {32'h424e5a76, 32'h42c5b8c0} /* (10, 0, 4) {real, imag} */,
  {32'h42d2376f, 32'h41c99788} /* (10, 0, 3) {real, imag} */,
  {32'hc2a14bc1, 32'hc1191404} /* (10, 0, 2) {real, imag} */,
  {32'h42a1b5c4, 32'h42b6b463} /* (10, 0, 1) {real, imag} */,
  {32'h4394ca79, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h4283dce2, 32'h3f389c80} /* (9, 15, 15) {real, imag} */,
  {32'hc2cb275f, 32'hc23244df} /* (9, 15, 14) {real, imag} */,
  {32'h41ad8398, 32'h42bf6550} /* (9, 15, 13) {real, imag} */,
  {32'hc21e2552, 32'hc27a58d8} /* (9, 15, 12) {real, imag} */,
  {32'hc21c3f67, 32'hc1e70d44} /* (9, 15, 11) {real, imag} */,
  {32'hc181d7ca, 32'hc1b41014} /* (9, 15, 10) {real, imag} */,
  {32'h42289a80, 32'h41d61ee8} /* (9, 15, 9) {real, imag} */,
  {32'h4276d67b, 32'h00000000} /* (9, 15, 8) {real, imag} */,
  {32'h42289a80, 32'hc1d61ee8} /* (9, 15, 7) {real, imag} */,
  {32'hc181d7ca, 32'h41b41014} /* (9, 15, 6) {real, imag} */,
  {32'hc21c3f67, 32'h41e70d44} /* (9, 15, 5) {real, imag} */,
  {32'hc21e2552, 32'h427a58d8} /* (9, 15, 4) {real, imag} */,
  {32'h41ad8398, 32'hc2bf6550} /* (9, 15, 3) {real, imag} */,
  {32'hc2cb275f, 32'h423244df} /* (9, 15, 2) {real, imag} */,
  {32'h4283dce2, 32'hbf389c80} /* (9, 15, 1) {real, imag} */,
  {32'h435d3b4e, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'hc2ad325b, 32'hc317e586} /* (9, 14, 15) {real, imag} */,
  {32'hc322514b, 32'hc39dd6e6} /* (9, 14, 14) {real, imag} */,
  {32'h43094dd4, 32'h420c842d} /* (9, 14, 13) {real, imag} */,
  {32'hc112c8a4, 32'h4386a62e} /* (9, 14, 12) {real, imag} */,
  {32'hc1db15ae, 32'hc2e56fe1} /* (9, 14, 11) {real, imag} */,
  {32'hc2393488, 32'hc18a1616} /* (9, 14, 10) {real, imag} */,
  {32'h42bd226f, 32'h42f7c652} /* (9, 14, 9) {real, imag} */,
  {32'hc2b5ea28, 32'h00000000} /* (9, 14, 8) {real, imag} */,
  {32'h42bd226f, 32'hc2f7c652} /* (9, 14, 7) {real, imag} */,
  {32'hc2393488, 32'h418a1616} /* (9, 14, 6) {real, imag} */,
  {32'hc1db15ae, 32'h42e56fe1} /* (9, 14, 5) {real, imag} */,
  {32'hc112c8a4, 32'hc386a62e} /* (9, 14, 4) {real, imag} */,
  {32'h43094dd4, 32'hc20c842d} /* (9, 14, 3) {real, imag} */,
  {32'hc322514b, 32'h439dd6e6} /* (9, 14, 2) {real, imag} */,
  {32'hc2ad325b, 32'h4317e586} /* (9, 14, 1) {real, imag} */,
  {32'h43d84624, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hc2b5c6c4, 32'h41bd9b28} /* (9, 13, 15) {real, imag} */,
  {32'h41bf81f8, 32'hc336c84b} /* (9, 13, 14) {real, imag} */,
  {32'h420885f6, 32'h42923316} /* (9, 13, 13) {real, imag} */,
  {32'h40672760, 32'h4387e0db} /* (9, 13, 12) {real, imag} */,
  {32'hc04754d0, 32'h4248eff4} /* (9, 13, 11) {real, imag} */,
  {32'h4246bffe, 32'hc196ff24} /* (9, 13, 10) {real, imag} */,
  {32'h429ec90f, 32'hc1dd36fe} /* (9, 13, 9) {real, imag} */,
  {32'h428649bd, 32'h00000000} /* (9, 13, 8) {real, imag} */,
  {32'h429ec90f, 32'h41dd36fe} /* (9, 13, 7) {real, imag} */,
  {32'h4246bffe, 32'h4196ff24} /* (9, 13, 6) {real, imag} */,
  {32'hc04754d0, 32'hc248eff4} /* (9, 13, 5) {real, imag} */,
  {32'h40672760, 32'hc387e0db} /* (9, 13, 4) {real, imag} */,
  {32'h420885f6, 32'hc2923316} /* (9, 13, 3) {real, imag} */,
  {32'h41bf81f8, 32'h4336c84b} /* (9, 13, 2) {real, imag} */,
  {32'hc2b5c6c4, 32'hc1bd9b28} /* (9, 13, 1) {real, imag} */,
  {32'h438c3aa2, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'hc34ded3c, 32'h429c0385} /* (9, 12, 15) {real, imag} */,
  {32'h42fc26f8, 32'h41dbe000} /* (9, 12, 14) {real, imag} */,
  {32'h42bb8fe6, 32'hc2e56724} /* (9, 12, 13) {real, imag} */,
  {32'h431ce32a, 32'hc140b8ac} /* (9, 12, 12) {real, imag} */,
  {32'hc298b897, 32'h42a793c3} /* (9, 12, 11) {real, imag} */,
  {32'hc208af22, 32'h429b88e9} /* (9, 12, 10) {real, imag} */,
  {32'h411bdef8, 32'h42167a97} /* (9, 12, 9) {real, imag} */,
  {32'h404d8390, 32'h00000000} /* (9, 12, 8) {real, imag} */,
  {32'h411bdef8, 32'hc2167a97} /* (9, 12, 7) {real, imag} */,
  {32'hc208af22, 32'hc29b88e9} /* (9, 12, 6) {real, imag} */,
  {32'hc298b897, 32'hc2a793c3} /* (9, 12, 5) {real, imag} */,
  {32'h431ce32a, 32'h4140b8ac} /* (9, 12, 4) {real, imag} */,
  {32'h42bb8fe6, 32'h42e56724} /* (9, 12, 3) {real, imag} */,
  {32'h42fc26f8, 32'hc1dbe000} /* (9, 12, 2) {real, imag} */,
  {32'hc34ded3c, 32'hc29c0385} /* (9, 12, 1) {real, imag} */,
  {32'h43da6420, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'h424d64a2, 32'h439a4088} /* (9, 11, 15) {real, imag} */,
  {32'h429b258c, 32'h41a1bd40} /* (9, 11, 14) {real, imag} */,
  {32'h4294b4f6, 32'hc33730fb} /* (9, 11, 13) {real, imag} */,
  {32'hc3174887, 32'h4339728e} /* (9, 11, 12) {real, imag} */,
  {32'hc130fad8, 32'h42361ec8} /* (9, 11, 11) {real, imag} */,
  {32'hc2709518, 32'hc1f6e704} /* (9, 11, 10) {real, imag} */,
  {32'hc282ec97, 32'hc205d7f2} /* (9, 11, 9) {real, imag} */,
  {32'hc2159560, 32'h00000000} /* (9, 11, 8) {real, imag} */,
  {32'hc282ec97, 32'h4205d7f2} /* (9, 11, 7) {real, imag} */,
  {32'hc2709518, 32'h41f6e704} /* (9, 11, 6) {real, imag} */,
  {32'hc130fad8, 32'hc2361ec8} /* (9, 11, 5) {real, imag} */,
  {32'hc3174887, 32'hc339728e} /* (9, 11, 4) {real, imag} */,
  {32'h4294b4f6, 32'h433730fb} /* (9, 11, 3) {real, imag} */,
  {32'h429b258c, 32'hc1a1bd40} /* (9, 11, 2) {real, imag} */,
  {32'h424d64a2, 32'hc39a4088} /* (9, 11, 1) {real, imag} */,
  {32'h44251f21, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h41f070a0, 32'h43598de2} /* (9, 10, 15) {real, imag} */,
  {32'h43509ec4, 32'h4269a956} /* (9, 10, 14) {real, imag} */,
  {32'hc3583d60, 32'hc2253122} /* (9, 10, 13) {real, imag} */,
  {32'hc1a127f5, 32'h41d55aa4} /* (9, 10, 12) {real, imag} */,
  {32'hc1e6a467, 32'hc1079ed8} /* (9, 10, 11) {real, imag} */,
  {32'hc30bd69e, 32'h432a636a} /* (9, 10, 10) {real, imag} */,
  {32'h42d0da6d, 32'hc2f1f581} /* (9, 10, 9) {real, imag} */,
  {32'hc12af200, 32'h00000000} /* (9, 10, 8) {real, imag} */,
  {32'h42d0da6d, 32'h42f1f581} /* (9, 10, 7) {real, imag} */,
  {32'hc30bd69e, 32'hc32a636a} /* (9, 10, 6) {real, imag} */,
  {32'hc1e6a467, 32'h41079ed8} /* (9, 10, 5) {real, imag} */,
  {32'hc1a127f5, 32'hc1d55aa4} /* (9, 10, 4) {real, imag} */,
  {32'hc3583d60, 32'h42253122} /* (9, 10, 3) {real, imag} */,
  {32'h43509ec4, 32'hc269a956} /* (9, 10, 2) {real, imag} */,
  {32'h41f070a0, 32'hc3598de2} /* (9, 10, 1) {real, imag} */,
  {32'h43f9e038, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'h42d5e806, 32'h4399c5ea} /* (9, 9, 15) {real, imag} */,
  {32'h4336e98e, 32'hc1be1048} /* (9, 9, 14) {real, imag} */,
  {32'hc2a08efe, 32'h4225229c} /* (9, 9, 13) {real, imag} */,
  {32'h425e17e3, 32'hc257ba06} /* (9, 9, 12) {real, imag} */,
  {32'hc2a5162f, 32'h42f34817} /* (9, 9, 11) {real, imag} */,
  {32'h430fb1fd, 32'h431c520c} /* (9, 9, 10) {real, imag} */,
  {32'h428aa203, 32'hc284f9a6} /* (9, 9, 9) {real, imag} */,
  {32'hc2b9cbac, 32'h00000000} /* (9, 9, 8) {real, imag} */,
  {32'h428aa203, 32'h4284f9a6} /* (9, 9, 7) {real, imag} */,
  {32'h430fb1fd, 32'hc31c520c} /* (9, 9, 6) {real, imag} */,
  {32'hc2a5162f, 32'hc2f34817} /* (9, 9, 5) {real, imag} */,
  {32'h425e17e3, 32'h4257ba06} /* (9, 9, 4) {real, imag} */,
  {32'hc2a08efe, 32'hc225229c} /* (9, 9, 3) {real, imag} */,
  {32'h4336e98e, 32'h41be1048} /* (9, 9, 2) {real, imag} */,
  {32'h42d5e806, 32'hc399c5ea} /* (9, 9, 1) {real, imag} */,
  {32'h43e64afc, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h42c4b983, 32'h4279f683} /* (9, 8, 15) {real, imag} */,
  {32'h42ad8052, 32'hc318ce46} /* (9, 8, 14) {real, imag} */,
  {32'h4235624a, 32'h42f8d508} /* (9, 8, 13) {real, imag} */,
  {32'hc2c489ca, 32'hc14ad2c8} /* (9, 8, 12) {real, imag} */,
  {32'hc11980fa, 32'h40c5e6e8} /* (9, 8, 11) {real, imag} */,
  {32'h41185e00, 32'h4206e0f9} /* (9, 8, 10) {real, imag} */,
  {32'h4271d517, 32'h42bb85a7} /* (9, 8, 9) {real, imag} */,
  {32'hc27502f4, 32'h00000000} /* (9, 8, 8) {real, imag} */,
  {32'h4271d517, 32'hc2bb85a7} /* (9, 8, 7) {real, imag} */,
  {32'h41185e00, 32'hc206e0f9} /* (9, 8, 6) {real, imag} */,
  {32'hc11980fa, 32'hc0c5e6e8} /* (9, 8, 5) {real, imag} */,
  {32'hc2c489ca, 32'h414ad2c8} /* (9, 8, 4) {real, imag} */,
  {32'h4235624a, 32'hc2f8d508} /* (9, 8, 3) {real, imag} */,
  {32'h42ad8052, 32'h4318ce46} /* (9, 8, 2) {real, imag} */,
  {32'h42c4b983, 32'hc279f683} /* (9, 8, 1) {real, imag} */,
  {32'h438c1801, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h429a99fe, 32'hc23b559c} /* (9, 7, 15) {real, imag} */,
  {32'hc2c9dbd4, 32'hc386b1f0} /* (9, 7, 14) {real, imag} */,
  {32'hc302f6e1, 32'h43092711} /* (9, 7, 13) {real, imag} */,
  {32'h428a1e80, 32'h42158c1e} /* (9, 7, 12) {real, imag} */,
  {32'hbf5d3a80, 32'hc3372201} /* (9, 7, 11) {real, imag} */,
  {32'hc1630ff0, 32'h420493be} /* (9, 7, 10) {real, imag} */,
  {32'h4249041a, 32'h42166cb4} /* (9, 7, 9) {real, imag} */,
  {32'h41da851a, 32'h00000000} /* (9, 7, 8) {real, imag} */,
  {32'h4249041a, 32'hc2166cb4} /* (9, 7, 7) {real, imag} */,
  {32'hc1630ff0, 32'hc20493be} /* (9, 7, 6) {real, imag} */,
  {32'hbf5d3a80, 32'h43372201} /* (9, 7, 5) {real, imag} */,
  {32'h428a1e80, 32'hc2158c1e} /* (9, 7, 4) {real, imag} */,
  {32'hc302f6e1, 32'hc3092711} /* (9, 7, 3) {real, imag} */,
  {32'hc2c9dbd4, 32'h4386b1f0} /* (9, 7, 2) {real, imag} */,
  {32'h429a99fe, 32'h423b559c} /* (9, 7, 1) {real, imag} */,
  {32'h43574a67, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h42991394, 32'hc21cc2c8} /* (9, 6, 15) {real, imag} */,
  {32'hc2d59ca5, 32'hc38b4aa3} /* (9, 6, 14) {real, imag} */,
  {32'h42e91430, 32'hc1920fc0} /* (9, 6, 13) {real, imag} */,
  {32'h41a4bc97, 32'h4335dd70} /* (9, 6, 12) {real, imag} */,
  {32'h42800d4f, 32'hc27faa0e} /* (9, 6, 11) {real, imag} */,
  {32'hc31c37e8, 32'h42fc6ab4} /* (9, 6, 10) {real, imag} */,
  {32'hc042a9e0, 32'hc26dff46} /* (9, 6, 9) {real, imag} */,
  {32'hc31bb6a6, 32'h00000000} /* (9, 6, 8) {real, imag} */,
  {32'hc042a9e0, 32'h426dff46} /* (9, 6, 7) {real, imag} */,
  {32'hc31c37e8, 32'hc2fc6ab4} /* (9, 6, 6) {real, imag} */,
  {32'h42800d4f, 32'h427faa0e} /* (9, 6, 5) {real, imag} */,
  {32'h41a4bc97, 32'hc335dd70} /* (9, 6, 4) {real, imag} */,
  {32'h42e91430, 32'h41920fc0} /* (9, 6, 3) {real, imag} */,
  {32'hc2d59ca5, 32'h438b4aa3} /* (9, 6, 2) {real, imag} */,
  {32'h42991394, 32'h421cc2c8} /* (9, 6, 1) {real, imag} */,
  {32'h432a26e1, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'hc2af0237, 32'h42ed3572} /* (9, 5, 15) {real, imag} */,
  {32'hc2f6a010, 32'hc38c6e4b} /* (9, 5, 14) {real, imag} */,
  {32'h432e135a, 32'hc26b9a23} /* (9, 5, 13) {real, imag} */,
  {32'hc2e0aa7a, 32'h422a7b98} /* (9, 5, 12) {real, imag} */,
  {32'hc13b23b0, 32'hc31edc72} /* (9, 5, 11) {real, imag} */,
  {32'hc25a14b8, 32'hc03d0b20} /* (9, 5, 10) {real, imag} */,
  {32'h41f7173c, 32'h422310da} /* (9, 5, 9) {real, imag} */,
  {32'h42a3235c, 32'h00000000} /* (9, 5, 8) {real, imag} */,
  {32'h41f7173c, 32'hc22310da} /* (9, 5, 7) {real, imag} */,
  {32'hc25a14b8, 32'h403d0b20} /* (9, 5, 6) {real, imag} */,
  {32'hc13b23b0, 32'h431edc72} /* (9, 5, 5) {real, imag} */,
  {32'hc2e0aa7a, 32'hc22a7b98} /* (9, 5, 4) {real, imag} */,
  {32'h432e135a, 32'h426b9a23} /* (9, 5, 3) {real, imag} */,
  {32'hc2f6a010, 32'h438c6e4b} /* (9, 5, 2) {real, imag} */,
  {32'hc2af0237, 32'hc2ed3572} /* (9, 5, 1) {real, imag} */,
  {32'h4385e52e, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'h42835584, 32'h4370186a} /* (9, 4, 15) {real, imag} */,
  {32'hc39808ac, 32'hc3946bd2} /* (9, 4, 14) {real, imag} */,
  {32'h41973018, 32'h42688705} /* (9, 4, 13) {real, imag} */,
  {32'h425b7472, 32'hc25b6419} /* (9, 4, 12) {real, imag} */,
  {32'h429fea7b, 32'hc2acac41} /* (9, 4, 11) {real, imag} */,
  {32'h41f4d1f5, 32'h4287ebdb} /* (9, 4, 10) {real, imag} */,
  {32'hc1153420, 32'hc2f4a100} /* (9, 4, 9) {real, imag} */,
  {32'h428cfa74, 32'h00000000} /* (9, 4, 8) {real, imag} */,
  {32'hc1153420, 32'h42f4a100} /* (9, 4, 7) {real, imag} */,
  {32'h41f4d1f5, 32'hc287ebdb} /* (9, 4, 6) {real, imag} */,
  {32'h429fea7b, 32'h42acac41} /* (9, 4, 5) {real, imag} */,
  {32'h425b7472, 32'h425b6419} /* (9, 4, 4) {real, imag} */,
  {32'h41973018, 32'hc2688705} /* (9, 4, 3) {real, imag} */,
  {32'hc39808ac, 32'h43946bd2} /* (9, 4, 2) {real, imag} */,
  {32'h42835584, 32'hc370186a} /* (9, 4, 1) {real, imag} */,
  {32'hc13d8a10, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'hbf8d3a80, 32'h433f7049} /* (9, 3, 15) {real, imag} */,
  {32'h42e95c1e, 32'hc147ec50} /* (9, 3, 14) {real, imag} */,
  {32'h4152bff6, 32'h4229ab9d} /* (9, 3, 13) {real, imag} */,
  {32'h42c29d72, 32'h42ae242c} /* (9, 3, 12) {real, imag} */,
  {32'hc3005213, 32'hc1d93d9d} /* (9, 3, 11) {real, imag} */,
  {32'hc2b0b5c1, 32'h433a05b6} /* (9, 3, 10) {real, imag} */,
  {32'h431ad870, 32'hc2030da2} /* (9, 3, 9) {real, imag} */,
  {32'hc3309408, 32'h00000000} /* (9, 3, 8) {real, imag} */,
  {32'h431ad870, 32'h42030da2} /* (9, 3, 7) {real, imag} */,
  {32'hc2b0b5c1, 32'hc33a05b6} /* (9, 3, 6) {real, imag} */,
  {32'hc3005213, 32'h41d93d9d} /* (9, 3, 5) {real, imag} */,
  {32'h42c29d72, 32'hc2ae242c} /* (9, 3, 4) {real, imag} */,
  {32'h4152bff6, 32'hc229ab9d} /* (9, 3, 3) {real, imag} */,
  {32'h42e95c1e, 32'h4147ec50} /* (9, 3, 2) {real, imag} */,
  {32'hbf8d3a80, 32'hc33f7049} /* (9, 3, 1) {real, imag} */,
  {32'hc3344a7b, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'h40389fa0, 32'h437d78fe} /* (9, 2, 15) {real, imag} */,
  {32'h4304b96b, 32'h421b1180} /* (9, 2, 14) {real, imag} */,
  {32'h42feb9b1, 32'h421f7b35} /* (9, 2, 13) {real, imag} */,
  {32'hc27458e7, 32'hc2443792} /* (9, 2, 12) {real, imag} */,
  {32'hc2817d8c, 32'h432ffb45} /* (9, 2, 11) {real, imag} */,
  {32'hc1d2dbc4, 32'hc122f4d4} /* (9, 2, 10) {real, imag} */,
  {32'hc2ffed91, 32'h42c46712} /* (9, 2, 9) {real, imag} */,
  {32'h42bcc6dc, 32'h00000000} /* (9, 2, 8) {real, imag} */,
  {32'hc2ffed91, 32'hc2c46712} /* (9, 2, 7) {real, imag} */,
  {32'hc1d2dbc4, 32'h4122f4d4} /* (9, 2, 6) {real, imag} */,
  {32'hc2817d8c, 32'hc32ffb45} /* (9, 2, 5) {real, imag} */,
  {32'hc27458e7, 32'h42443792} /* (9, 2, 4) {real, imag} */,
  {32'h42feb9b1, 32'hc21f7b35} /* (9, 2, 3) {real, imag} */,
  {32'h4304b96b, 32'hc21b1180} /* (9, 2, 2) {real, imag} */,
  {32'h40389fa0, 32'hc37d78fe} /* (9, 2, 1) {real, imag} */,
  {32'hc286806e, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'hc32451df, 32'h42bf2be5} /* (9, 1, 15) {real, imag} */,
  {32'hc2a03fc9, 32'hc11baa64} /* (9, 1, 14) {real, imag} */,
  {32'hc19dd46c, 32'hc2510847} /* (9, 1, 13) {real, imag} */,
  {32'h434c2d38, 32'hc325b831} /* (9, 1, 12) {real, imag} */,
  {32'h427b4061, 32'h4353c60e} /* (9, 1, 11) {real, imag} */,
  {32'h409fe958, 32'h4345faea} /* (9, 1, 10) {real, imag} */,
  {32'hc237f400, 32'hc2c537fe} /* (9, 1, 9) {real, imag} */,
  {32'h4020e310, 32'h00000000} /* (9, 1, 8) {real, imag} */,
  {32'hc237f400, 32'h42c537fe} /* (9, 1, 7) {real, imag} */,
  {32'h409fe958, 32'hc345faea} /* (9, 1, 6) {real, imag} */,
  {32'h427b4061, 32'hc353c60e} /* (9, 1, 5) {real, imag} */,
  {32'h434c2d38, 32'h4325b831} /* (9, 1, 4) {real, imag} */,
  {32'hc19dd46c, 32'h42510847} /* (9, 1, 3) {real, imag} */,
  {32'hc2a03fc9, 32'h411baa64} /* (9, 1, 2) {real, imag} */,
  {32'hc32451df, 32'hc2bf2be5} /* (9, 1, 1) {real, imag} */,
  {32'h431a996a, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'hc2870703, 32'h41260b84} /* (9, 0, 15) {real, imag} */,
  {32'hc1700c70, 32'hc1c3c8f0} /* (9, 0, 14) {real, imag} */,
  {32'h424ea332, 32'h406cd100} /* (9, 0, 13) {real, imag} */,
  {32'hc12f4414, 32'hc2a16fc7} /* (9, 0, 12) {real, imag} */,
  {32'hc0b134b4, 32'hc1c2038e} /* (9, 0, 11) {real, imag} */,
  {32'hc298b5be, 32'hc25e72f7} /* (9, 0, 10) {real, imag} */,
  {32'hc2054331, 32'hbfef4f00} /* (9, 0, 9) {real, imag} */,
  {32'hbf0a4300, 32'h00000000} /* (9, 0, 8) {real, imag} */,
  {32'hc2054331, 32'h3fef4f00} /* (9, 0, 7) {real, imag} */,
  {32'hc298b5be, 32'h425e72f7} /* (9, 0, 6) {real, imag} */,
  {32'hc0b134b4, 32'h41c2038e} /* (9, 0, 5) {real, imag} */,
  {32'hc12f4414, 32'h42a16fc7} /* (9, 0, 4) {real, imag} */,
  {32'h424ea332, 32'hc06cd100} /* (9, 0, 3) {real, imag} */,
  {32'hc1700c70, 32'h41c3c8f0} /* (9, 0, 2) {real, imag} */,
  {32'hc2870703, 32'hc1260b84} /* (9, 0, 1) {real, imag} */,
  {32'h42a62f0f, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'hc0db6160, 32'hc2d91a02} /* (8, 15, 15) {real, imag} */,
  {32'hc214be58, 32'h41557878} /* (8, 15, 14) {real, imag} */,
  {32'h431b7c15, 32'hc22e022f} /* (8, 15, 13) {real, imag} */,
  {32'hc192d63c, 32'h4255f490} /* (8, 15, 12) {real, imag} */,
  {32'h418396c6, 32'h41ea8660} /* (8, 15, 11) {real, imag} */,
  {32'hc1d5b534, 32'h422a782e} /* (8, 15, 10) {real, imag} */,
  {32'hc1eebd86, 32'hc25426a2} /* (8, 15, 9) {real, imag} */,
  {32'hc289240b, 32'h00000000} /* (8, 15, 8) {real, imag} */,
  {32'hc1eebd86, 32'h425426a2} /* (8, 15, 7) {real, imag} */,
  {32'hc1d5b534, 32'hc22a782e} /* (8, 15, 6) {real, imag} */,
  {32'h418396c6, 32'hc1ea8660} /* (8, 15, 5) {real, imag} */,
  {32'hc192d63c, 32'hc255f490} /* (8, 15, 4) {real, imag} */,
  {32'h431b7c15, 32'h422e022f} /* (8, 15, 3) {real, imag} */,
  {32'hc214be58, 32'hc1557878} /* (8, 15, 2) {real, imag} */,
  {32'hc0db6160, 32'h42d91a02} /* (8, 15, 1) {real, imag} */,
  {32'h4084ace8, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'h4148d550, 32'hc2c2cece} /* (8, 14, 15) {real, imag} */,
  {32'hc2034388, 32'hc2df7c54} /* (8, 14, 14) {real, imag} */,
  {32'h4239cfed, 32'h41c3f49e} /* (8, 14, 13) {real, imag} */,
  {32'hc29e71b5, 32'hc2b488ff} /* (8, 14, 12) {real, imag} */,
  {32'hc2b7befc, 32'hc30a2e76} /* (8, 14, 11) {real, imag} */,
  {32'h4301db19, 32'h429aeb32} /* (8, 14, 10) {real, imag} */,
  {32'h41a6fec2, 32'h420dd77e} /* (8, 14, 9) {real, imag} */,
  {32'hc1c146f8, 32'h00000000} /* (8, 14, 8) {real, imag} */,
  {32'h41a6fec2, 32'hc20dd77e} /* (8, 14, 7) {real, imag} */,
  {32'h4301db19, 32'hc29aeb32} /* (8, 14, 6) {real, imag} */,
  {32'hc2b7befc, 32'h430a2e76} /* (8, 14, 5) {real, imag} */,
  {32'hc29e71b5, 32'h42b488ff} /* (8, 14, 4) {real, imag} */,
  {32'h4239cfed, 32'hc1c3f49e} /* (8, 14, 3) {real, imag} */,
  {32'hc2034388, 32'h42df7c54} /* (8, 14, 2) {real, imag} */,
  {32'h4148d550, 32'h42c2cece} /* (8, 14, 1) {real, imag} */,
  {32'h409b1160, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'hc30f98f0, 32'h42b050ac} /* (8, 13, 15) {real, imag} */,
  {32'h4191eced, 32'hc257285a} /* (8, 13, 14) {real, imag} */,
  {32'h433c924d, 32'hc187f428} /* (8, 13, 13) {real, imag} */,
  {32'h42e1bfe1, 32'h432b2eea} /* (8, 13, 12) {real, imag} */,
  {32'hc257a2fa, 32'hc332612d} /* (8, 13, 11) {real, imag} */,
  {32'hc2994e45, 32'hc0edb030} /* (8, 13, 10) {real, imag} */,
  {32'h42200a5e, 32'hc29ca54f} /* (8, 13, 9) {real, imag} */,
  {32'h428b1601, 32'h00000000} /* (8, 13, 8) {real, imag} */,
  {32'h42200a5e, 32'h429ca54f} /* (8, 13, 7) {real, imag} */,
  {32'hc2994e45, 32'h40edb030} /* (8, 13, 6) {real, imag} */,
  {32'hc257a2fa, 32'h4332612d} /* (8, 13, 5) {real, imag} */,
  {32'h42e1bfe1, 32'hc32b2eea} /* (8, 13, 4) {real, imag} */,
  {32'h433c924d, 32'h4187f428} /* (8, 13, 3) {real, imag} */,
  {32'h4191eced, 32'h4257285a} /* (8, 13, 2) {real, imag} */,
  {32'hc30f98f0, 32'hc2b050ac} /* (8, 13, 1) {real, imag} */,
  {32'h430803ac, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'hc09ece30, 32'h421fb865} /* (8, 12, 15) {real, imag} */,
  {32'h424a4119, 32'h42ccf41e} /* (8, 12, 14) {real, imag} */,
  {32'hc2b33b26, 32'hc2136342} /* (8, 12, 13) {real, imag} */,
  {32'hc22d0f57, 32'h41e5ef58} /* (8, 12, 12) {real, imag} */,
  {32'h42ee6ab0, 32'hc013fef0} /* (8, 12, 11) {real, imag} */,
  {32'hc23a8118, 32'hc1782ee0} /* (8, 12, 10) {real, imag} */,
  {32'h3ed1af80, 32'hc080abf0} /* (8, 12, 9) {real, imag} */,
  {32'h419a9138, 32'h00000000} /* (8, 12, 8) {real, imag} */,
  {32'h3ed1af80, 32'h4080abf0} /* (8, 12, 7) {real, imag} */,
  {32'hc23a8118, 32'h41782ee0} /* (8, 12, 6) {real, imag} */,
  {32'h42ee6ab0, 32'h4013fef0} /* (8, 12, 5) {real, imag} */,
  {32'hc22d0f57, 32'hc1e5ef58} /* (8, 12, 4) {real, imag} */,
  {32'hc2b33b26, 32'h42136342} /* (8, 12, 3) {real, imag} */,
  {32'h424a4119, 32'hc2ccf41e} /* (8, 12, 2) {real, imag} */,
  {32'hc09ece30, 32'hc21fb865} /* (8, 12, 1) {real, imag} */,
  {32'h435273c7, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'h4197d204, 32'h4309e85c} /* (8, 11, 15) {real, imag} */,
  {32'h4330e0e3, 32'h4283a41e} /* (8, 11, 14) {real, imag} */,
  {32'hc301363b, 32'hc35ccf59} /* (8, 11, 13) {real, imag} */,
  {32'hc2882c91, 32'hc0ca4a78} /* (8, 11, 12) {real, imag} */,
  {32'h42b30dbf, 32'h426d3b1d} /* (8, 11, 11) {real, imag} */,
  {32'hc2136b32, 32'h41d360ce} /* (8, 11, 10) {real, imag} */,
  {32'h41dec33c, 32'hc1c7132d} /* (8, 11, 9) {real, imag} */,
  {32'hc30bab18, 32'h00000000} /* (8, 11, 8) {real, imag} */,
  {32'h41dec33c, 32'h41c7132d} /* (8, 11, 7) {real, imag} */,
  {32'hc2136b32, 32'hc1d360ce} /* (8, 11, 6) {real, imag} */,
  {32'h42b30dbf, 32'hc26d3b1d} /* (8, 11, 5) {real, imag} */,
  {32'hc2882c91, 32'h40ca4a78} /* (8, 11, 4) {real, imag} */,
  {32'hc301363b, 32'h435ccf59} /* (8, 11, 3) {real, imag} */,
  {32'h4330e0e3, 32'hc283a41e} /* (8, 11, 2) {real, imag} */,
  {32'h4197d204, 32'hc309e85c} /* (8, 11, 1) {real, imag} */,
  {32'h4324a9d7, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h40aa0210, 32'h43948808} /* (8, 10, 15) {real, imag} */,
  {32'h42f8ff66, 32'h42967424} /* (8, 10, 14) {real, imag} */,
  {32'hc28f62e6, 32'h40993580} /* (8, 10, 13) {real, imag} */,
  {32'hc21aaa85, 32'h42f993db} /* (8, 10, 12) {real, imag} */,
  {32'hbfe78dc0, 32'hc3020dde} /* (8, 10, 11) {real, imag} */,
  {32'h42d17bd0, 32'h422a5733} /* (8, 10, 10) {real, imag} */,
  {32'hc3028a21, 32'hc2c283a6} /* (8, 10, 9) {real, imag} */,
  {32'h3f1577c0, 32'h00000000} /* (8, 10, 8) {real, imag} */,
  {32'hc3028a21, 32'h42c283a6} /* (8, 10, 7) {real, imag} */,
  {32'h42d17bd0, 32'hc22a5733} /* (8, 10, 6) {real, imag} */,
  {32'hbfe78dc0, 32'h43020dde} /* (8, 10, 5) {real, imag} */,
  {32'hc21aaa85, 32'hc2f993db} /* (8, 10, 4) {real, imag} */,
  {32'hc28f62e6, 32'hc0993580} /* (8, 10, 3) {real, imag} */,
  {32'h42f8ff66, 32'hc2967424} /* (8, 10, 2) {real, imag} */,
  {32'h40aa0210, 32'hc3948808} /* (8, 10, 1) {real, imag} */,
  {32'h43cca602, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'hc12d3e64, 32'h4355f84c} /* (8, 9, 15) {real, imag} */,
  {32'hc25aeeeb, 32'hc1926b68} /* (8, 9, 14) {real, imag} */,
  {32'h423607ee, 32'hbecac180} /* (8, 9, 13) {real, imag} */,
  {32'hc184ff64, 32'h422da93a} /* (8, 9, 12) {real, imag} */,
  {32'h41da0e44, 32'h42a47d80} /* (8, 9, 11) {real, imag} */,
  {32'hc23be39e, 32'h42124490} /* (8, 9, 10) {real, imag} */,
  {32'hc29298e8, 32'hc1c062cb} /* (8, 9, 9) {real, imag} */,
  {32'h41629028, 32'h00000000} /* (8, 9, 8) {real, imag} */,
  {32'hc29298e8, 32'h41c062cb} /* (8, 9, 7) {real, imag} */,
  {32'hc23be39e, 32'hc2124490} /* (8, 9, 6) {real, imag} */,
  {32'h41da0e44, 32'hc2a47d80} /* (8, 9, 5) {real, imag} */,
  {32'hc184ff64, 32'hc22da93a} /* (8, 9, 4) {real, imag} */,
  {32'h423607ee, 32'h3ecac180} /* (8, 9, 3) {real, imag} */,
  {32'hc25aeeeb, 32'h41926b68} /* (8, 9, 2) {real, imag} */,
  {32'hc12d3e64, 32'hc355f84c} /* (8, 9, 1) {real, imag} */,
  {32'h43af2f5a, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'h42b8861c, 32'hc2331945} /* (8, 8, 15) {real, imag} */,
  {32'hc1943612, 32'hc34cbf76} /* (8, 8, 14) {real, imag} */,
  {32'h42c81478, 32'h43753841} /* (8, 8, 13) {real, imag} */,
  {32'h427530cf, 32'h42c10c09} /* (8, 8, 12) {real, imag} */,
  {32'hc26ff4b1, 32'h42bd7352} /* (8, 8, 11) {real, imag} */,
  {32'h4299f146, 32'hc2b83472} /* (8, 8, 10) {real, imag} */,
  {32'hc28de1e6, 32'h41bcd85d} /* (8, 8, 9) {real, imag} */,
  {32'hc20a68c5, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'hc28de1e6, 32'hc1bcd85d} /* (8, 8, 7) {real, imag} */,
  {32'h4299f146, 32'h42b83472} /* (8, 8, 6) {real, imag} */,
  {32'hc26ff4b1, 32'hc2bd7352} /* (8, 8, 5) {real, imag} */,
  {32'h427530cf, 32'hc2c10c09} /* (8, 8, 4) {real, imag} */,
  {32'h42c81478, 32'hc3753841} /* (8, 8, 3) {real, imag} */,
  {32'hc1943612, 32'h434cbf76} /* (8, 8, 2) {real, imag} */,
  {32'h42b8861c, 32'h42331945} /* (8, 8, 1) {real, imag} */,
  {32'h42564728, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'hc2ce726a, 32'hc33b2920} /* (8, 7, 15) {real, imag} */,
  {32'hc19c4c4a, 32'hc32b9074} /* (8, 7, 14) {real, imag} */,
  {32'h420a0100, 32'h42eb2074} /* (8, 7, 13) {real, imag} */,
  {32'h423ce2d0, 32'hc2a68bdb} /* (8, 7, 12) {real, imag} */,
  {32'h42761472, 32'hc260f960} /* (8, 7, 11) {real, imag} */,
  {32'hc2a214f7, 32'h4221e9ca} /* (8, 7, 10) {real, imag} */,
  {32'h40ea7258, 32'h429d2b03} /* (8, 7, 9) {real, imag} */,
  {32'h43177014, 32'h00000000} /* (8, 7, 8) {real, imag} */,
  {32'h40ea7258, 32'hc29d2b03} /* (8, 7, 7) {real, imag} */,
  {32'hc2a214f7, 32'hc221e9ca} /* (8, 7, 6) {real, imag} */,
  {32'h42761472, 32'h4260f960} /* (8, 7, 5) {real, imag} */,
  {32'h423ce2d0, 32'h42a68bdb} /* (8, 7, 4) {real, imag} */,
  {32'h420a0100, 32'hc2eb2074} /* (8, 7, 3) {real, imag} */,
  {32'hc19c4c4a, 32'h432b9074} /* (8, 7, 2) {real, imag} */,
  {32'hc2ce726a, 32'h433b2920} /* (8, 7, 1) {real, imag} */,
  {32'h434e2444, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'hc2105262, 32'h4284b546} /* (8, 6, 15) {real, imag} */,
  {32'hc2fe0cb6, 32'hc34207d4} /* (8, 6, 14) {real, imag} */,
  {32'h43162ac3, 32'h4162df08} /* (8, 6, 13) {real, imag} */,
  {32'h41e7b78a, 32'h4293e711} /* (8, 6, 12) {real, imag} */,
  {32'hc37374aa, 32'hc1d5efcc} /* (8, 6, 11) {real, imag} */,
  {32'h42267ae4, 32'h429d8a18} /* (8, 6, 10) {real, imag} */,
  {32'hc245b553, 32'hc279ee25} /* (8, 6, 9) {real, imag} */,
  {32'hc1d7bba8, 32'h00000000} /* (8, 6, 8) {real, imag} */,
  {32'hc245b553, 32'h4279ee25} /* (8, 6, 7) {real, imag} */,
  {32'h42267ae4, 32'hc29d8a18} /* (8, 6, 6) {real, imag} */,
  {32'hc37374aa, 32'h41d5efcc} /* (8, 6, 5) {real, imag} */,
  {32'h41e7b78a, 32'hc293e711} /* (8, 6, 4) {real, imag} */,
  {32'h43162ac3, 32'hc162df08} /* (8, 6, 3) {real, imag} */,
  {32'hc2fe0cb6, 32'h434207d4} /* (8, 6, 2) {real, imag} */,
  {32'hc2105262, 32'hc284b546} /* (8, 6, 1) {real, imag} */,
  {32'h41acaa38, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'hc1155ad9, 32'h43015134} /* (8, 5, 15) {real, imag} */,
  {32'hc3521845, 32'hc371f569} /* (8, 5, 14) {real, imag} */,
  {32'h42a73316, 32'hc137a3d0} /* (8, 5, 13) {real, imag} */,
  {32'hc1779340, 32'h425b944b} /* (8, 5, 12) {real, imag} */,
  {32'h41076bc8, 32'hc1acb4b2} /* (8, 5, 11) {real, imag} */,
  {32'hc230b164, 32'h4213ac6c} /* (8, 5, 10) {real, imag} */,
  {32'h4245b9de, 32'h4187425b} /* (8, 5, 9) {real, imag} */,
  {32'h42566666, 32'h00000000} /* (8, 5, 8) {real, imag} */,
  {32'h4245b9de, 32'hc187425b} /* (8, 5, 7) {real, imag} */,
  {32'hc230b164, 32'hc213ac6c} /* (8, 5, 6) {real, imag} */,
  {32'h41076bc8, 32'h41acb4b2} /* (8, 5, 5) {real, imag} */,
  {32'hc1779340, 32'hc25b944b} /* (8, 5, 4) {real, imag} */,
  {32'h42a73316, 32'h4137a3d0} /* (8, 5, 3) {real, imag} */,
  {32'hc3521845, 32'h4371f569} /* (8, 5, 2) {real, imag} */,
  {32'hc1155ad9, 32'hc3015134} /* (8, 5, 1) {real, imag} */,
  {32'h42d1fb86, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'hc2c09288, 32'h42f015f0} /* (8, 4, 15) {real, imag} */,
  {32'hc2f5dfcc, 32'hc384cff2} /* (8, 4, 14) {real, imag} */,
  {32'hc3252861, 32'hc284d471} /* (8, 4, 13) {real, imag} */,
  {32'hc1e88086, 32'h42154110} /* (8, 4, 12) {real, imag} */,
  {32'h432f1b32, 32'h43021cd5} /* (8, 4, 11) {real, imag} */,
  {32'hc1ac0fe5, 32'h42e126de} /* (8, 4, 10) {real, imag} */,
  {32'h429ef340, 32'h41ce0654} /* (8, 4, 9) {real, imag} */,
  {32'h41380fa0, 32'h00000000} /* (8, 4, 8) {real, imag} */,
  {32'h429ef340, 32'hc1ce0654} /* (8, 4, 7) {real, imag} */,
  {32'hc1ac0fe5, 32'hc2e126de} /* (8, 4, 6) {real, imag} */,
  {32'h432f1b32, 32'hc3021cd5} /* (8, 4, 5) {real, imag} */,
  {32'hc1e88086, 32'hc2154110} /* (8, 4, 4) {real, imag} */,
  {32'hc3252861, 32'h4284d471} /* (8, 4, 3) {real, imag} */,
  {32'hc2f5dfcc, 32'h4384cff2} /* (8, 4, 2) {real, imag} */,
  {32'hc2c09288, 32'hc2f015f0} /* (8, 4, 1) {real, imag} */,
  {32'h430e11b9, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'hc315c040, 32'h436bf436} /* (8, 3, 15) {real, imag} */,
  {32'hc2357e16, 32'hc32ef804} /* (8, 3, 14) {real, imag} */,
  {32'h4287fbde, 32'h4315317f} /* (8, 3, 13) {real, imag} */,
  {32'h4154a4a0, 32'hc2b6bf89} /* (8, 3, 12) {real, imag} */,
  {32'hc2ad1123, 32'hc2e955f7} /* (8, 3, 11) {real, imag} */,
  {32'hc283c661, 32'h421ce0c1} /* (8, 3, 10) {real, imag} */,
  {32'h41c41e4c, 32'h4287120f} /* (8, 3, 9) {real, imag} */,
  {32'h42647bc6, 32'h00000000} /* (8, 3, 8) {real, imag} */,
  {32'h41c41e4c, 32'hc287120f} /* (8, 3, 7) {real, imag} */,
  {32'hc283c661, 32'hc21ce0c1} /* (8, 3, 6) {real, imag} */,
  {32'hc2ad1123, 32'h42e955f7} /* (8, 3, 5) {real, imag} */,
  {32'h4154a4a0, 32'h42b6bf89} /* (8, 3, 4) {real, imag} */,
  {32'h4287fbde, 32'hc315317f} /* (8, 3, 3) {real, imag} */,
  {32'hc2357e16, 32'h432ef804} /* (8, 3, 2) {real, imag} */,
  {32'hc315c040, 32'hc36bf436} /* (8, 3, 1) {real, imag} */,
  {32'h400dfd00, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'hc32c77e6, 32'h43b5d34e} /* (8, 2, 15) {real, imag} */,
  {32'hc28b511f, 32'hc287f958} /* (8, 2, 14) {real, imag} */,
  {32'h432b68a1, 32'hc2e66140} /* (8, 2, 13) {real, imag} */,
  {32'hc29bf565, 32'hc29457b1} /* (8, 2, 12) {real, imag} */,
  {32'hc237b093, 32'hc2c11c6c} /* (8, 2, 11) {real, imag} */,
  {32'hc155e29c, 32'h42cd45c8} /* (8, 2, 10) {real, imag} */,
  {32'hc16daab4, 32'hc28e18d6} /* (8, 2, 9) {real, imag} */,
  {32'h42c06c52, 32'h00000000} /* (8, 2, 8) {real, imag} */,
  {32'hc16daab4, 32'h428e18d6} /* (8, 2, 7) {real, imag} */,
  {32'hc155e29c, 32'hc2cd45c8} /* (8, 2, 6) {real, imag} */,
  {32'hc237b093, 32'h42c11c6c} /* (8, 2, 5) {real, imag} */,
  {32'hc29bf565, 32'h429457b1} /* (8, 2, 4) {real, imag} */,
  {32'h432b68a1, 32'h42e66140} /* (8, 2, 3) {real, imag} */,
  {32'hc28b511f, 32'h4287f958} /* (8, 2, 2) {real, imag} */,
  {32'hc32c77e6, 32'hc3b5d34e} /* (8, 2, 1) {real, imag} */,
  {32'hc323c8af, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'hc3844d74, 32'h4324da3b} /* (8, 1, 15) {real, imag} */,
  {32'hc141f9ba, 32'hc2af24a5} /* (8, 1, 14) {real, imag} */,
  {32'h41980378, 32'hc0166650} /* (8, 1, 13) {real, imag} */,
  {32'h41e65090, 32'h42f8063a} /* (8, 1, 12) {real, imag} */,
  {32'h414de5ef, 32'hc3793d0c} /* (8, 1, 11) {real, imag} */,
  {32'hc32a6ede, 32'h423f86e8} /* (8, 1, 10) {real, imag} */,
  {32'h428db042, 32'h41a686b5} /* (8, 1, 9) {real, imag} */,
  {32'hc18f8987, 32'h00000000} /* (8, 1, 8) {real, imag} */,
  {32'h428db042, 32'hc1a686b5} /* (8, 1, 7) {real, imag} */,
  {32'hc32a6ede, 32'hc23f86e8} /* (8, 1, 6) {real, imag} */,
  {32'h414de5ef, 32'h43793d0c} /* (8, 1, 5) {real, imag} */,
  {32'h41e65090, 32'hc2f8063a} /* (8, 1, 4) {real, imag} */,
  {32'h41980378, 32'h40166650} /* (8, 1, 3) {real, imag} */,
  {32'hc141f9ba, 32'h42af24a5} /* (8, 1, 2) {real, imag} */,
  {32'hc3844d74, 32'hc324da3b} /* (8, 1, 1) {real, imag} */,
  {32'hc2ae503c, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'hc35994b4, 32'h42a2016c} /* (8, 0, 15) {real, imag} */,
  {32'hc235ca21, 32'hc303218c} /* (8, 0, 14) {real, imag} */,
  {32'hc2a63950, 32'h424ad76c} /* (8, 0, 13) {real, imag} */,
  {32'h41dfce3e, 32'h425a00d6} /* (8, 0, 12) {real, imag} */,
  {32'h41401a2c, 32'hc22e6979} /* (8, 0, 11) {real, imag} */,
  {32'h4216d4c9, 32'hc26c5aa8} /* (8, 0, 10) {real, imag} */,
  {32'h41e4c006, 32'h40c74d2c} /* (8, 0, 9) {real, imag} */,
  {32'h41a2924e, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'h41e4c006, 32'hc0c74d2c} /* (8, 0, 7) {real, imag} */,
  {32'h4216d4c9, 32'h426c5aa8} /* (8, 0, 6) {real, imag} */,
  {32'h41401a2c, 32'h422e6979} /* (8, 0, 5) {real, imag} */,
  {32'h41dfce3e, 32'hc25a00d6} /* (8, 0, 4) {real, imag} */,
  {32'hc2a63950, 32'hc24ad76c} /* (8, 0, 3) {real, imag} */,
  {32'hc235ca21, 32'h4303218c} /* (8, 0, 2) {real, imag} */,
  {32'hc35994b4, 32'hc2a2016c} /* (8, 0, 1) {real, imag} */,
  {32'h42960e62, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'hc2b2c51b, 32'h41c658a0} /* (7, 15, 15) {real, imag} */,
  {32'h42a500f6, 32'hc33c7792} /* (7, 15, 14) {real, imag} */,
  {32'h42cdf092, 32'h42ad40fc} /* (7, 15, 13) {real, imag} */,
  {32'hc304e06c, 32'hc13bc0f8} /* (7, 15, 12) {real, imag} */,
  {32'hc1269540, 32'h407e8630} /* (7, 15, 11) {real, imag} */,
  {32'h40f83d30, 32'h41cf7a0e} /* (7, 15, 10) {real, imag} */,
  {32'hc115a374, 32'hc00e8ac8} /* (7, 15, 9) {real, imag} */,
  {32'hc2cb9e1a, 32'h00000000} /* (7, 15, 8) {real, imag} */,
  {32'hc115a374, 32'h400e8ac8} /* (7, 15, 7) {real, imag} */,
  {32'h40f83d30, 32'hc1cf7a0e} /* (7, 15, 6) {real, imag} */,
  {32'hc1269540, 32'hc07e8630} /* (7, 15, 5) {real, imag} */,
  {32'hc304e06c, 32'h413bc0f8} /* (7, 15, 4) {real, imag} */,
  {32'h42cdf092, 32'hc2ad40fc} /* (7, 15, 3) {real, imag} */,
  {32'h42a500f6, 32'h433c7792} /* (7, 15, 2) {real, imag} */,
  {32'hc2b2c51b, 32'hc1c658a0} /* (7, 15, 1) {real, imag} */,
  {32'hc3332b80, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'h41fbd7a8, 32'h4322868a} /* (7, 14, 15) {real, imag} */,
  {32'h4311955d, 32'hc32ce404} /* (7, 14, 14) {real, imag} */,
  {32'h42c83962, 32'h4274a0ce} /* (7, 14, 13) {real, imag} */,
  {32'hc28dc3fc, 32'hc260d254} /* (7, 14, 12) {real, imag} */,
  {32'hc31cc144, 32'hc21bd5b9} /* (7, 14, 11) {real, imag} */,
  {32'h4303d33e, 32'h41822154} /* (7, 14, 10) {real, imag} */,
  {32'h40ea1ceb, 32'h42151f94} /* (7, 14, 9) {real, imag} */,
  {32'hc2c2bd38, 32'h00000000} /* (7, 14, 8) {real, imag} */,
  {32'h40ea1ceb, 32'hc2151f94} /* (7, 14, 7) {real, imag} */,
  {32'h4303d33e, 32'hc1822154} /* (7, 14, 6) {real, imag} */,
  {32'hc31cc144, 32'h421bd5b9} /* (7, 14, 5) {real, imag} */,
  {32'hc28dc3fc, 32'h4260d254} /* (7, 14, 4) {real, imag} */,
  {32'h42c83962, 32'hc274a0ce} /* (7, 14, 3) {real, imag} */,
  {32'h4311955d, 32'h432ce404} /* (7, 14, 2) {real, imag} */,
  {32'h41fbd7a8, 32'hc322868a} /* (7, 14, 1) {real, imag} */,
  {32'hc35004ca, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hc31fcf14, 32'h42ff9664} /* (7, 13, 15) {real, imag} */,
  {32'h42168e04, 32'hc1f2d780} /* (7, 13, 14) {real, imag} */,
  {32'h42350a16, 32'h42995854} /* (7, 13, 13) {real, imag} */,
  {32'hc0f4e040, 32'h42de77a4} /* (7, 13, 12) {real, imag} */,
  {32'hc19cac3a, 32'hc340c88a} /* (7, 13, 11) {real, imag} */,
  {32'hc1f81810, 32'h437b8b97} /* (7, 13, 10) {real, imag} */,
  {32'hc2a98aef, 32'hc27380a8} /* (7, 13, 9) {real, imag} */,
  {32'h4305c111, 32'h00000000} /* (7, 13, 8) {real, imag} */,
  {32'hc2a98aef, 32'h427380a8} /* (7, 13, 7) {real, imag} */,
  {32'hc1f81810, 32'hc37b8b97} /* (7, 13, 6) {real, imag} */,
  {32'hc19cac3a, 32'h4340c88a} /* (7, 13, 5) {real, imag} */,
  {32'hc0f4e040, 32'hc2de77a4} /* (7, 13, 4) {real, imag} */,
  {32'h42350a16, 32'hc2995854} /* (7, 13, 3) {real, imag} */,
  {32'h42168e04, 32'h41f2d780} /* (7, 13, 2) {real, imag} */,
  {32'hc31fcf14, 32'hc2ff9664} /* (7, 13, 1) {real, imag} */,
  {32'h43554f2b, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'h423b20b6, 32'h42ddf84e} /* (7, 12, 15) {real, imag} */,
  {32'h42a80d46, 32'hc110de50} /* (7, 12, 14) {real, imag} */,
  {32'hc2e74841, 32'hc28dfe07} /* (7, 12, 13) {real, imag} */,
  {32'h41778f4c, 32'h42ad6e0c} /* (7, 12, 12) {real, imag} */,
  {32'h429e26d8, 32'hc2c437c8} /* (7, 12, 11) {real, imag} */,
  {32'hc18bd4cc, 32'hc1106390} /* (7, 12, 10) {real, imag} */,
  {32'h430328de, 32'hc249f85a} /* (7, 12, 9) {real, imag} */,
  {32'hc248b1ef, 32'h00000000} /* (7, 12, 8) {real, imag} */,
  {32'h430328de, 32'h4249f85a} /* (7, 12, 7) {real, imag} */,
  {32'hc18bd4cc, 32'h41106390} /* (7, 12, 6) {real, imag} */,
  {32'h429e26d8, 32'h42c437c8} /* (7, 12, 5) {real, imag} */,
  {32'h41778f4c, 32'hc2ad6e0c} /* (7, 12, 4) {real, imag} */,
  {32'hc2e74841, 32'h428dfe07} /* (7, 12, 3) {real, imag} */,
  {32'h42a80d46, 32'h4110de50} /* (7, 12, 2) {real, imag} */,
  {32'h423b20b6, 32'hc2ddf84e} /* (7, 12, 1) {real, imag} */,
  {32'h4166e1f8, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'h4212ae86, 32'h4370328d} /* (7, 11, 15) {real, imag} */,
  {32'hc185d0b4, 32'hc26a7250} /* (7, 11, 14) {real, imag} */,
  {32'hc2b33096, 32'hc304d44d} /* (7, 11, 13) {real, imag} */,
  {32'h41462440, 32'hc1c93263} /* (7, 11, 12) {real, imag} */,
  {32'h413954b0, 32'h428d3874} /* (7, 11, 11) {real, imag} */,
  {32'h41f175d4, 32'hc228b099} /* (7, 11, 10) {real, imag} */,
  {32'h424f1b69, 32'h422c2040} /* (7, 11, 9) {real, imag} */,
  {32'hc12888d4, 32'h00000000} /* (7, 11, 8) {real, imag} */,
  {32'h424f1b69, 32'hc22c2040} /* (7, 11, 7) {real, imag} */,
  {32'h41f175d4, 32'h4228b099} /* (7, 11, 6) {real, imag} */,
  {32'h413954b0, 32'hc28d3874} /* (7, 11, 5) {real, imag} */,
  {32'h41462440, 32'h41c93263} /* (7, 11, 4) {real, imag} */,
  {32'hc2b33096, 32'h4304d44d} /* (7, 11, 3) {real, imag} */,
  {32'hc185d0b4, 32'h426a7250} /* (7, 11, 2) {real, imag} */,
  {32'h4212ae86, 32'hc370328d} /* (7, 11, 1) {real, imag} */,
  {32'h4305d582, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'hc2bcd07f, 32'h438f5609} /* (7, 10, 15) {real, imag} */,
  {32'hc2ea68bf, 32'h4288484c} /* (7, 10, 14) {real, imag} */,
  {32'hc2f2c672, 32'hc31222fc} /* (7, 10, 13) {real, imag} */,
  {32'hc1cdffce, 32'h427cfd72} /* (7, 10, 12) {real, imag} */,
  {32'h42a2cb40, 32'h424f6e31} /* (7, 10, 11) {real, imag} */,
  {32'hc1072980, 32'hc32978d6} /* (7, 10, 10) {real, imag} */,
  {32'h422749e4, 32'hc1d35afc} /* (7, 10, 9) {real, imag} */,
  {32'hc1295a2c, 32'h00000000} /* (7, 10, 8) {real, imag} */,
  {32'h422749e4, 32'h41d35afc} /* (7, 10, 7) {real, imag} */,
  {32'hc1072980, 32'h432978d6} /* (7, 10, 6) {real, imag} */,
  {32'h42a2cb40, 32'hc24f6e31} /* (7, 10, 5) {real, imag} */,
  {32'hc1cdffce, 32'hc27cfd72} /* (7, 10, 4) {real, imag} */,
  {32'hc2f2c672, 32'h431222fc} /* (7, 10, 3) {real, imag} */,
  {32'hc2ea68bf, 32'hc288484c} /* (7, 10, 2) {real, imag} */,
  {32'hc2bcd07f, 32'hc38f5609} /* (7, 10, 1) {real, imag} */,
  {32'h43fa3e3c, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'h42214c8e, 32'h432dfca4} /* (7, 9, 15) {real, imag} */,
  {32'hc28c275b, 32'h4286b69b} /* (7, 9, 14) {real, imag} */,
  {32'h43039df0, 32'hbfa51fc0} /* (7, 9, 13) {real, imag} */,
  {32'h41d8b0c4, 32'h42fba728} /* (7, 9, 12) {real, imag} */,
  {32'hc3122f4f, 32'hc27005d8} /* (7, 9, 11) {real, imag} */,
  {32'h424d6e45, 32'h42a53c4c} /* (7, 9, 10) {real, imag} */,
  {32'hc219b97f, 32'h413d65ac} /* (7, 9, 9) {real, imag} */,
  {32'hc2bab0c2, 32'h00000000} /* (7, 9, 8) {real, imag} */,
  {32'hc219b97f, 32'hc13d65ac} /* (7, 9, 7) {real, imag} */,
  {32'h424d6e45, 32'hc2a53c4c} /* (7, 9, 6) {real, imag} */,
  {32'hc3122f4f, 32'h427005d8} /* (7, 9, 5) {real, imag} */,
  {32'h41d8b0c4, 32'hc2fba728} /* (7, 9, 4) {real, imag} */,
  {32'h43039df0, 32'h3fa51fc0} /* (7, 9, 3) {real, imag} */,
  {32'hc28c275b, 32'hc286b69b} /* (7, 9, 2) {real, imag} */,
  {32'h42214c8e, 32'hc32dfca4} /* (7, 9, 1) {real, imag} */,
  {32'h43733410, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'hc277f4e4, 32'h431be3d0} /* (7, 8, 15) {real, imag} */,
  {32'h41ab54f1, 32'hbfdcc000} /* (7, 8, 14) {real, imag} */,
  {32'hc0eb91e0, 32'h41e2347c} /* (7, 8, 13) {real, imag} */,
  {32'h41b95f10, 32'h41e9cae6} /* (7, 8, 12) {real, imag} */,
  {32'h42540e1e, 32'hc1b69092} /* (7, 8, 11) {real, imag} */,
  {32'h415071ac, 32'h4276c773} /* (7, 8, 10) {real, imag} */,
  {32'hc191c7b4, 32'h429acd16} /* (7, 8, 9) {real, imag} */,
  {32'hc2a05dfa, 32'h00000000} /* (7, 8, 8) {real, imag} */,
  {32'hc191c7b4, 32'hc29acd16} /* (7, 8, 7) {real, imag} */,
  {32'h415071ac, 32'hc276c773} /* (7, 8, 6) {real, imag} */,
  {32'h42540e1e, 32'h41b69092} /* (7, 8, 5) {real, imag} */,
  {32'h41b95f10, 32'hc1e9cae6} /* (7, 8, 4) {real, imag} */,
  {32'hc0eb91e0, 32'hc1e2347c} /* (7, 8, 3) {real, imag} */,
  {32'h41ab54f1, 32'h3fdcc000} /* (7, 8, 2) {real, imag} */,
  {32'hc277f4e4, 32'hc31be3d0} /* (7, 8, 1) {real, imag} */,
  {32'h43786abe, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'hc329fff4, 32'h41483140} /* (7, 7, 15) {real, imag} */,
  {32'hc2ace409, 32'h415884d8} /* (7, 7, 14) {real, imag} */,
  {32'h425300da, 32'hc0e87d50} /* (7, 7, 13) {real, imag} */,
  {32'hc2f6d867, 32'hc2e62282} /* (7, 7, 12) {real, imag} */,
  {32'h427d25e8, 32'hc2f5e8e0} /* (7, 7, 11) {real, imag} */,
  {32'h41f9f8fe, 32'hc3159647} /* (7, 7, 10) {real, imag} */,
  {32'h412d1ccd, 32'hc2817d74} /* (7, 7, 9) {real, imag} */,
  {32'hc18b4936, 32'h00000000} /* (7, 7, 8) {real, imag} */,
  {32'h412d1ccd, 32'h42817d74} /* (7, 7, 7) {real, imag} */,
  {32'h41f9f8fe, 32'h43159647} /* (7, 7, 6) {real, imag} */,
  {32'h427d25e8, 32'h42f5e8e0} /* (7, 7, 5) {real, imag} */,
  {32'hc2f6d867, 32'h42e62282} /* (7, 7, 4) {real, imag} */,
  {32'h425300da, 32'h40e87d50} /* (7, 7, 3) {real, imag} */,
  {32'hc2ace409, 32'hc15884d8} /* (7, 7, 2) {real, imag} */,
  {32'hc329fff4, 32'hc1483140} /* (7, 7, 1) {real, imag} */,
  {32'hc31c9efc, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'hc351c238, 32'h42c2c40d} /* (7, 6, 15) {real, imag} */,
  {32'h42e19ceb, 32'h41adb002} /* (7, 6, 14) {real, imag} */,
  {32'h42d11706, 32'hc247700a} /* (7, 6, 13) {real, imag} */,
  {32'h42f62d32, 32'h43059568} /* (7, 6, 12) {real, imag} */,
  {32'hc1a12386, 32'h42484d4b} /* (7, 6, 11) {real, imag} */,
  {32'h425b6875, 32'h430b1948} /* (7, 6, 10) {real, imag} */,
  {32'hc264af40, 32'hc2a009bf} /* (7, 6, 9) {real, imag} */,
  {32'h422fc8df, 32'h00000000} /* (7, 6, 8) {real, imag} */,
  {32'hc264af40, 32'h42a009bf} /* (7, 6, 7) {real, imag} */,
  {32'h425b6875, 32'hc30b1948} /* (7, 6, 6) {real, imag} */,
  {32'hc1a12386, 32'hc2484d4b} /* (7, 6, 5) {real, imag} */,
  {32'h42f62d32, 32'hc3059568} /* (7, 6, 4) {real, imag} */,
  {32'h42d11706, 32'h4247700a} /* (7, 6, 3) {real, imag} */,
  {32'h42e19ceb, 32'hc1adb002} /* (7, 6, 2) {real, imag} */,
  {32'hc351c238, 32'hc2c2c40d} /* (7, 6, 1) {real, imag} */,
  {32'hc36180df, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'hc37196e8, 32'h434f267d} /* (7, 5, 15) {real, imag} */,
  {32'hc10f6e48, 32'hc321cbc0} /* (7, 5, 14) {real, imag} */,
  {32'h42a7cdb2, 32'hc296f310} /* (7, 5, 13) {real, imag} */,
  {32'h4295acb2, 32'h42af54be} /* (7, 5, 12) {real, imag} */,
  {32'hc1c2a888, 32'h421fda03} /* (7, 5, 11) {real, imag} */,
  {32'hc2acedd4, 32'h42279197} /* (7, 5, 10) {real, imag} */,
  {32'h4243d497, 32'hc2cf0570} /* (7, 5, 9) {real, imag} */,
  {32'hc2ab0532, 32'h00000000} /* (7, 5, 8) {real, imag} */,
  {32'h4243d497, 32'h42cf0570} /* (7, 5, 7) {real, imag} */,
  {32'hc2acedd4, 32'hc2279197} /* (7, 5, 6) {real, imag} */,
  {32'hc1c2a888, 32'hc21fda03} /* (7, 5, 5) {real, imag} */,
  {32'h4295acb2, 32'hc2af54be} /* (7, 5, 4) {real, imag} */,
  {32'h42a7cdb2, 32'h4296f310} /* (7, 5, 3) {real, imag} */,
  {32'hc10f6e48, 32'h4321cbc0} /* (7, 5, 2) {real, imag} */,
  {32'hc37196e8, 32'hc34f267d} /* (7, 5, 1) {real, imag} */,
  {32'hc29d3504, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'hc3948899, 32'h429ed08c} /* (7, 4, 15) {real, imag} */,
  {32'hc32f6923, 32'hc347cd5d} /* (7, 4, 14) {real, imag} */,
  {32'h42d96729, 32'hc2cc2a2d} /* (7, 4, 13) {real, imag} */,
  {32'h43001173, 32'h43237439} /* (7, 4, 12) {real, imag} */,
  {32'h42106649, 32'hc29ba7be} /* (7, 4, 11) {real, imag} */,
  {32'hc09b89f0, 32'h43817908} /* (7, 4, 10) {real, imag} */,
  {32'h429fc312, 32'hc2dcfddb} /* (7, 4, 9) {real, imag} */,
  {32'hc2c5d3a8, 32'h00000000} /* (7, 4, 8) {real, imag} */,
  {32'h429fc312, 32'h42dcfddb} /* (7, 4, 7) {real, imag} */,
  {32'hc09b89f0, 32'hc3817908} /* (7, 4, 6) {real, imag} */,
  {32'h42106649, 32'h429ba7be} /* (7, 4, 5) {real, imag} */,
  {32'h43001173, 32'hc3237439} /* (7, 4, 4) {real, imag} */,
  {32'h42d96729, 32'h42cc2a2d} /* (7, 4, 3) {real, imag} */,
  {32'hc32f6923, 32'h4347cd5d} /* (7, 4, 2) {real, imag} */,
  {32'hc3948899, 32'hc29ed08c} /* (7, 4, 1) {real, imag} */,
  {32'h427af9d6, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'hc353fca8, 32'hc1ea9840} /* (7, 3, 15) {real, imag} */,
  {32'hc34b2bcd, 32'hc3959254} /* (7, 3, 14) {real, imag} */,
  {32'h414575b8, 32'hc1270070} /* (7, 3, 13) {real, imag} */,
  {32'hc2c6545a, 32'h428495c8} /* (7, 3, 12) {real, imag} */,
  {32'hc21bb873, 32'h42e62914} /* (7, 3, 11) {real, imag} */,
  {32'h4352b452, 32'hc10fb850} /* (7, 3, 10) {real, imag} */,
  {32'h429771f5, 32'hc0e81680} /* (7, 3, 9) {real, imag} */,
  {32'hc1e0fbba, 32'h00000000} /* (7, 3, 8) {real, imag} */,
  {32'h429771f5, 32'h40e81680} /* (7, 3, 7) {real, imag} */,
  {32'h4352b452, 32'h410fb850} /* (7, 3, 6) {real, imag} */,
  {32'hc21bb873, 32'hc2e62914} /* (7, 3, 5) {real, imag} */,
  {32'hc2c6545a, 32'hc28495c8} /* (7, 3, 4) {real, imag} */,
  {32'h414575b8, 32'h41270070} /* (7, 3, 3) {real, imag} */,
  {32'hc34b2bcd, 32'h43959254} /* (7, 3, 2) {real, imag} */,
  {32'hc353fca8, 32'h41ea9840} /* (7, 3, 1) {real, imag} */,
  {32'h41e1c398, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'hc329f1ec, 32'h424cba54} /* (7, 2, 15) {real, imag} */,
  {32'hc374cb13, 32'hc39a95f3} /* (7, 2, 14) {real, imag} */,
  {32'h42022d6b, 32'hc142c108} /* (7, 2, 13) {real, imag} */,
  {32'h422fffbd, 32'h41505600} /* (7, 2, 12) {real, imag} */,
  {32'h41aa5a54, 32'hc3204abf} /* (7, 2, 11) {real, imag} */,
  {32'hc21f2f0c, 32'hc2a09b08} /* (7, 2, 10) {real, imag} */,
  {32'hc18246a7, 32'h41e82b68} /* (7, 2, 9) {real, imag} */,
  {32'hbf54e8c0, 32'h00000000} /* (7, 2, 8) {real, imag} */,
  {32'hc18246a7, 32'hc1e82b68} /* (7, 2, 7) {real, imag} */,
  {32'hc21f2f0c, 32'h42a09b08} /* (7, 2, 6) {real, imag} */,
  {32'h41aa5a54, 32'h43204abf} /* (7, 2, 5) {real, imag} */,
  {32'h422fffbd, 32'hc1505600} /* (7, 2, 4) {real, imag} */,
  {32'h42022d6b, 32'h4142c108} /* (7, 2, 3) {real, imag} */,
  {32'hc374cb13, 32'h439a95f3} /* (7, 2, 2) {real, imag} */,
  {32'hc329f1ec, 32'hc24cba54} /* (7, 2, 1) {real, imag} */,
  {32'hc38c4dbc, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'hc311ac36, 32'h4340a772} /* (7, 1, 15) {real, imag} */,
  {32'hc326d274, 32'hc361272a} /* (7, 1, 14) {real, imag} */,
  {32'h428b4442, 32'hc2aec21a} /* (7, 1, 13) {real, imag} */,
  {32'h422f35be, 32'hc31d87b6} /* (7, 1, 12) {real, imag} */,
  {32'h431830ad, 32'hc23b8d79} /* (7, 1, 11) {real, imag} */,
  {32'hc312af96, 32'hc2294d85} /* (7, 1, 10) {real, imag} */,
  {32'h423f1ec1, 32'h425ecd68} /* (7, 1, 9) {real, imag} */,
  {32'h4246fe3d, 32'h00000000} /* (7, 1, 8) {real, imag} */,
  {32'h423f1ec1, 32'hc25ecd68} /* (7, 1, 7) {real, imag} */,
  {32'hc312af96, 32'h42294d85} /* (7, 1, 6) {real, imag} */,
  {32'h431830ad, 32'h423b8d79} /* (7, 1, 5) {real, imag} */,
  {32'h422f35be, 32'h431d87b6} /* (7, 1, 4) {real, imag} */,
  {32'h428b4442, 32'h42aec21a} /* (7, 1, 3) {real, imag} */,
  {32'hc326d274, 32'h4361272a} /* (7, 1, 2) {real, imag} */,
  {32'hc311ac36, 32'hc340a772} /* (7, 1, 1) {real, imag} */,
  {32'hc3351690, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'hc3128e5a, 32'h42fc0e98} /* (7, 0, 15) {real, imag} */,
  {32'hc0019118, 32'h411297e8} /* (7, 0, 14) {real, imag} */,
  {32'h429a890d, 32'hc1b3f57c} /* (7, 0, 13) {real, imag} */,
  {32'h428de68e, 32'h42880fac} /* (7, 0, 12) {real, imag} */,
  {32'h3f85af30, 32'hc22ba923} /* (7, 0, 11) {real, imag} */,
  {32'h422a9f21, 32'h428108ee} /* (7, 0, 10) {real, imag} */,
  {32'h423a735e, 32'hc1d60251} /* (7, 0, 9) {real, imag} */,
  {32'h423f81a4, 32'h00000000} /* (7, 0, 8) {real, imag} */,
  {32'h423a735e, 32'h41d60251} /* (7, 0, 7) {real, imag} */,
  {32'h422a9f21, 32'hc28108ee} /* (7, 0, 6) {real, imag} */,
  {32'h3f85af30, 32'h422ba923} /* (7, 0, 5) {real, imag} */,
  {32'h428de68e, 32'hc2880fac} /* (7, 0, 4) {real, imag} */,
  {32'h429a890d, 32'h41b3f57c} /* (7, 0, 3) {real, imag} */,
  {32'hc0019118, 32'hc11297e8} /* (7, 0, 2) {real, imag} */,
  {32'hc3128e5a, 32'hc2fc0e98} /* (7, 0, 1) {real, imag} */,
  {32'hc18f9e14, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'hc2b28212, 32'h421e05fc} /* (6, 15, 15) {real, imag} */,
  {32'h430c9306, 32'hc23397b3} /* (6, 15, 14) {real, imag} */,
  {32'hc10c5f90, 32'h414e7bd0} /* (6, 15, 13) {real, imag} */,
  {32'hc149f820, 32'hc23dc9f8} /* (6, 15, 12) {real, imag} */,
  {32'hc0fad260, 32'hc1ae3ed1} /* (6, 15, 11) {real, imag} */,
  {32'h42a14b42, 32'h4280a9a8} /* (6, 15, 10) {real, imag} */,
  {32'hc13f08ec, 32'h4266bd62} /* (6, 15, 9) {real, imag} */,
  {32'h41857e52, 32'h00000000} /* (6, 15, 8) {real, imag} */,
  {32'hc13f08ec, 32'hc266bd62} /* (6, 15, 7) {real, imag} */,
  {32'h42a14b42, 32'hc280a9a8} /* (6, 15, 6) {real, imag} */,
  {32'hc0fad260, 32'h41ae3ed1} /* (6, 15, 5) {real, imag} */,
  {32'hc149f820, 32'h423dc9f8} /* (6, 15, 4) {real, imag} */,
  {32'hc10c5f90, 32'hc14e7bd0} /* (6, 15, 3) {real, imag} */,
  {32'h430c9306, 32'h423397b3} /* (6, 15, 2) {real, imag} */,
  {32'hc2b28212, 32'hc21e05fc} /* (6, 15, 1) {real, imag} */,
  {32'hc392e42c, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'hc29fdb75, 32'h42c01356} /* (6, 14, 15) {real, imag} */,
  {32'h42dd6c7c, 32'hc0d2b800} /* (6, 14, 14) {real, imag} */,
  {32'h4284e5c5, 32'h41d63912} /* (6, 14, 13) {real, imag} */,
  {32'h42b1411c, 32'hc1d2e884} /* (6, 14, 12) {real, imag} */,
  {32'h41b07b88, 32'hc25d4c30} /* (6, 14, 11) {real, imag} */,
  {32'h4091c070, 32'h427345f2} /* (6, 14, 10) {real, imag} */,
  {32'hc26f4360, 32'hc20f9664} /* (6, 14, 9) {real, imag} */,
  {32'h41859404, 32'h00000000} /* (6, 14, 8) {real, imag} */,
  {32'hc26f4360, 32'h420f9664} /* (6, 14, 7) {real, imag} */,
  {32'h4091c070, 32'hc27345f2} /* (6, 14, 6) {real, imag} */,
  {32'h41b07b88, 32'h425d4c30} /* (6, 14, 5) {real, imag} */,
  {32'h42b1411c, 32'h41d2e884} /* (6, 14, 4) {real, imag} */,
  {32'h4284e5c5, 32'hc1d63912} /* (6, 14, 3) {real, imag} */,
  {32'h42dd6c7c, 32'h40d2b800} /* (6, 14, 2) {real, imag} */,
  {32'hc29fdb75, 32'hc2c01356} /* (6, 14, 1) {real, imag} */,
  {32'hc38ae7a8, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hc2b25226, 32'h42a6c730} /* (6, 13, 15) {real, imag} */,
  {32'h42b33b26, 32'h41ad1046} /* (6, 13, 14) {real, imag} */,
  {32'h428c4390, 32'h418e38d1} /* (6, 13, 13) {real, imag} */,
  {32'hc3388d81, 32'h3fdab240} /* (6, 13, 12) {real, imag} */,
  {32'h42400c23, 32'h4273e292} /* (6, 13, 11) {real, imag} */,
  {32'hc26c231e, 32'hc29f7cc0} /* (6, 13, 10) {real, imag} */,
  {32'h41ecac65, 32'h42349de8} /* (6, 13, 9) {real, imag} */,
  {32'hc12dffae, 32'h00000000} /* (6, 13, 8) {real, imag} */,
  {32'h41ecac65, 32'hc2349de8} /* (6, 13, 7) {real, imag} */,
  {32'hc26c231e, 32'h429f7cc0} /* (6, 13, 6) {real, imag} */,
  {32'h42400c23, 32'hc273e292} /* (6, 13, 5) {real, imag} */,
  {32'hc3388d81, 32'hbfdab240} /* (6, 13, 4) {real, imag} */,
  {32'h428c4390, 32'hc18e38d1} /* (6, 13, 3) {real, imag} */,
  {32'h42b33b26, 32'hc1ad1046} /* (6, 13, 2) {real, imag} */,
  {32'hc2b25226, 32'hc2a6c730} /* (6, 13, 1) {real, imag} */,
  {32'hc39dd480, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'hc2709ef4, 32'h434058b7} /* (6, 12, 15) {real, imag} */,
  {32'hc177f603, 32'hc136bc10} /* (6, 12, 14) {real, imag} */,
  {32'hc1723828, 32'hc20a7148} /* (6, 12, 13) {real, imag} */,
  {32'h421f0ea8, 32'hc2a2ffa4} /* (6, 12, 12) {real, imag} */,
  {32'h41883508, 32'h40db5060} /* (6, 12, 11) {real, imag} */,
  {32'h430e362f, 32'h4206ded8} /* (6, 12, 10) {real, imag} */,
  {32'hc2e99f39, 32'hc2f4be92} /* (6, 12, 9) {real, imag} */,
  {32'h40b71460, 32'h00000000} /* (6, 12, 8) {real, imag} */,
  {32'hc2e99f39, 32'h42f4be92} /* (6, 12, 7) {real, imag} */,
  {32'h430e362f, 32'hc206ded8} /* (6, 12, 6) {real, imag} */,
  {32'h41883508, 32'hc0db5060} /* (6, 12, 5) {real, imag} */,
  {32'h421f0ea8, 32'h42a2ffa4} /* (6, 12, 4) {real, imag} */,
  {32'hc1723828, 32'h420a7148} /* (6, 12, 3) {real, imag} */,
  {32'hc177f603, 32'h4136bc10} /* (6, 12, 2) {real, imag} */,
  {32'hc2709ef4, 32'hc34058b7} /* (6, 12, 1) {real, imag} */,
  {32'hc2bdeecc, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'h436b155e, 32'h438c8116} /* (6, 11, 15) {real, imag} */,
  {32'hc14be60c, 32'hc326aaa8} /* (6, 11, 14) {real, imag} */,
  {32'hc285fae5, 32'hc30265ea} /* (6, 11, 13) {real, imag} */,
  {32'h407cddb8, 32'hc204ff0b} /* (6, 11, 12) {real, imag} */,
  {32'hc2c58ce2, 32'hc225d163} /* (6, 11, 11) {real, imag} */,
  {32'hc258ff7c, 32'h42fe11c6} /* (6, 11, 10) {real, imag} */,
  {32'hc2c87819, 32'h430f0e4e} /* (6, 11, 9) {real, imag} */,
  {32'h4177ff6a, 32'h00000000} /* (6, 11, 8) {real, imag} */,
  {32'hc2c87819, 32'hc30f0e4e} /* (6, 11, 7) {real, imag} */,
  {32'hc258ff7c, 32'hc2fe11c6} /* (6, 11, 6) {real, imag} */,
  {32'hc2c58ce2, 32'h4225d163} /* (6, 11, 5) {real, imag} */,
  {32'h407cddb8, 32'h4204ff0b} /* (6, 11, 4) {real, imag} */,
  {32'hc285fae5, 32'h430265ea} /* (6, 11, 3) {real, imag} */,
  {32'hc14be60c, 32'h4326aaa8} /* (6, 11, 2) {real, imag} */,
  {32'h436b155e, 32'hc38c8116} /* (6, 11, 1) {real, imag} */,
  {32'h42df5a3e, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h4319fbf8, 32'h43dfc8d4} /* (6, 10, 15) {real, imag} */,
  {32'hc2197920, 32'h42c9636c} /* (6, 10, 14) {real, imag} */,
  {32'hc208a0b4, 32'hc32587c7} /* (6, 10, 13) {real, imag} */,
  {32'h428792d8, 32'hc2ddd199} /* (6, 10, 12) {real, imag} */,
  {32'h418cfb4e, 32'hc1f39abf} /* (6, 10, 11) {real, imag} */,
  {32'hc280bf9d, 32'h430a87b9} /* (6, 10, 10) {real, imag} */,
  {32'hc1e46d2a, 32'h428cd722} /* (6, 10, 9) {real, imag} */,
  {32'hc24ceda0, 32'h00000000} /* (6, 10, 8) {real, imag} */,
  {32'hc1e46d2a, 32'hc28cd722} /* (6, 10, 7) {real, imag} */,
  {32'hc280bf9d, 32'hc30a87b9} /* (6, 10, 6) {real, imag} */,
  {32'h418cfb4e, 32'h41f39abf} /* (6, 10, 5) {real, imag} */,
  {32'h428792d8, 32'h42ddd199} /* (6, 10, 4) {real, imag} */,
  {32'hc208a0b4, 32'h432587c7} /* (6, 10, 3) {real, imag} */,
  {32'hc2197920, 32'hc2c9636c} /* (6, 10, 2) {real, imag} */,
  {32'h4319fbf8, 32'hc3dfc8d4} /* (6, 10, 1) {real, imag} */,
  {32'h4391185e, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'hc31e1490, 32'h438d1785} /* (6, 9, 15) {real, imag} */,
  {32'h4306ebac, 32'h42c64a92} /* (6, 9, 14) {real, imag} */,
  {32'h4262fafc, 32'hc2782a90} /* (6, 9, 13) {real, imag} */,
  {32'h42770cf4, 32'hc2d91518} /* (6, 9, 12) {real, imag} */,
  {32'hc3531fdf, 32'hc2948304} /* (6, 9, 11) {real, imag} */,
  {32'hc2fd045b, 32'h41968e22} /* (6, 9, 10) {real, imag} */,
  {32'hc282f445, 32'hc2a5d3ca} /* (6, 9, 9) {real, imag} */,
  {32'hc28b62f2, 32'h00000000} /* (6, 9, 8) {real, imag} */,
  {32'hc282f445, 32'h42a5d3ca} /* (6, 9, 7) {real, imag} */,
  {32'hc2fd045b, 32'hc1968e22} /* (6, 9, 6) {real, imag} */,
  {32'hc3531fdf, 32'h42948304} /* (6, 9, 5) {real, imag} */,
  {32'h42770cf4, 32'h42d91518} /* (6, 9, 4) {real, imag} */,
  {32'h4262fafc, 32'h42782a90} /* (6, 9, 3) {real, imag} */,
  {32'h4306ebac, 32'hc2c64a92} /* (6, 9, 2) {real, imag} */,
  {32'hc31e1490, 32'hc38d1785} /* (6, 9, 1) {real, imag} */,
  {32'h43d24c9e, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'hc2e77078, 32'h434b5f2a} /* (6, 8, 15) {real, imag} */,
  {32'h42e62783, 32'hc2a1914e} /* (6, 8, 14) {real, imag} */,
  {32'h4287da96, 32'hc2c15cf4} /* (6, 8, 13) {real, imag} */,
  {32'hc253985c, 32'hc301a08c} /* (6, 8, 12) {real, imag} */,
  {32'hc21eceb1, 32'hc3130365} /* (6, 8, 11) {real, imag} */,
  {32'hc274d5de, 32'hc22c96da} /* (6, 8, 10) {real, imag} */,
  {32'h41f61b82, 32'h42a1fd04} /* (6, 8, 9) {real, imag} */,
  {32'hc28a0268, 32'h00000000} /* (6, 8, 8) {real, imag} */,
  {32'h41f61b82, 32'hc2a1fd04} /* (6, 8, 7) {real, imag} */,
  {32'hc274d5de, 32'h422c96da} /* (6, 8, 6) {real, imag} */,
  {32'hc21eceb1, 32'h43130365} /* (6, 8, 5) {real, imag} */,
  {32'hc253985c, 32'h4301a08c} /* (6, 8, 4) {real, imag} */,
  {32'h4287da96, 32'h42c15cf4} /* (6, 8, 3) {real, imag} */,
  {32'h42e62783, 32'h42a1914e} /* (6, 8, 2) {real, imag} */,
  {32'hc2e77078, 32'hc34b5f2a} /* (6, 8, 1) {real, imag} */,
  {32'h419fc464, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h42aec618, 32'h43a05d87} /* (6, 7, 15) {real, imag} */,
  {32'h4339a8a0, 32'h42b4bdb0} /* (6, 7, 14) {real, imag} */,
  {32'h42641cd6, 32'h412432c8} /* (6, 7, 13) {real, imag} */,
  {32'hc2c75358, 32'hc29b8f8c} /* (6, 7, 12) {real, imag} */,
  {32'h431a427d, 32'h41bbcaa0} /* (6, 7, 11) {real, imag} */,
  {32'h4199e884, 32'h4294a1c2} /* (6, 7, 10) {real, imag} */,
  {32'hc0cc8eac, 32'h4090f0a8} /* (6, 7, 9) {real, imag} */,
  {32'hc2539117, 32'h00000000} /* (6, 7, 8) {real, imag} */,
  {32'hc0cc8eac, 32'hc090f0a8} /* (6, 7, 7) {real, imag} */,
  {32'h4199e884, 32'hc294a1c2} /* (6, 7, 6) {real, imag} */,
  {32'h431a427d, 32'hc1bbcaa0} /* (6, 7, 5) {real, imag} */,
  {32'hc2c75358, 32'h429b8f8c} /* (6, 7, 4) {real, imag} */,
  {32'h42641cd6, 32'hc12432c8} /* (6, 7, 3) {real, imag} */,
  {32'h4339a8a0, 32'hc2b4bdb0} /* (6, 7, 2) {real, imag} */,
  {32'h42aec618, 32'hc3a05d87} /* (6, 7, 1) {real, imag} */,
  {32'hc39d2ffc, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'hc28d044f, 32'h43137c88} /* (6, 6, 15) {real, imag} */,
  {32'h42f01156, 32'h42047281} /* (6, 6, 14) {real, imag} */,
  {32'h43091d53, 32'h41a75108} /* (6, 6, 13) {real, imag} */,
  {32'hc320abd0, 32'hc2b08f8b} /* (6, 6, 12) {real, imag} */,
  {32'hc06264f0, 32'h4257151e} /* (6, 6, 11) {real, imag} */,
  {32'h42986be7, 32'hc12ab080} /* (6, 6, 10) {real, imag} */,
  {32'hc1ebf312, 32'hc2a15c16} /* (6, 6, 9) {real, imag} */,
  {32'h41eafb30, 32'h00000000} /* (6, 6, 8) {real, imag} */,
  {32'hc1ebf312, 32'h42a15c16} /* (6, 6, 7) {real, imag} */,
  {32'h42986be7, 32'h412ab080} /* (6, 6, 6) {real, imag} */,
  {32'hc06264f0, 32'hc257151e} /* (6, 6, 5) {real, imag} */,
  {32'hc320abd0, 32'h42b08f8b} /* (6, 6, 4) {real, imag} */,
  {32'h43091d53, 32'hc1a75108} /* (6, 6, 3) {real, imag} */,
  {32'h42f01156, 32'hc2047281} /* (6, 6, 2) {real, imag} */,
  {32'hc28d044f, 32'hc3137c88} /* (6, 6, 1) {real, imag} */,
  {32'hc3893920, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'hc3964ef7, 32'h42ce6cce} /* (6, 5, 15) {real, imag} */,
  {32'h429b6b56, 32'hc351b3c4} /* (6, 5, 14) {real, imag} */,
  {32'h4253bee8, 32'hbf44e080} /* (6, 5, 13) {real, imag} */,
  {32'h41ba0e21, 32'h420f2e79} /* (6, 5, 12) {real, imag} */,
  {32'h428a5c50, 32'h41bd217a} /* (6, 5, 11) {real, imag} */,
  {32'h42438002, 32'hc1334480} /* (6, 5, 10) {real, imag} */,
  {32'h4267bdb6, 32'hc2de2083} /* (6, 5, 9) {real, imag} */,
  {32'hc1420472, 32'h00000000} /* (6, 5, 8) {real, imag} */,
  {32'h4267bdb6, 32'h42de2083} /* (6, 5, 7) {real, imag} */,
  {32'h42438002, 32'h41334480} /* (6, 5, 6) {real, imag} */,
  {32'h428a5c50, 32'hc1bd217a} /* (6, 5, 5) {real, imag} */,
  {32'h41ba0e21, 32'hc20f2e79} /* (6, 5, 4) {real, imag} */,
  {32'h4253bee8, 32'h3f44e080} /* (6, 5, 3) {real, imag} */,
  {32'h429b6b56, 32'h4351b3c4} /* (6, 5, 2) {real, imag} */,
  {32'hc3964ef7, 32'hc2ce6cce} /* (6, 5, 1) {real, imag} */,
  {32'hc3d3c9f0, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'hc350c289, 32'hc292d272} /* (6, 4, 15) {real, imag} */,
  {32'hc1308b0b, 32'hc35d3dcb} /* (6, 4, 14) {real, imag} */,
  {32'h42a0f8d7, 32'hc27eea54} /* (6, 4, 13) {real, imag} */,
  {32'h41916808, 32'h434ffed2} /* (6, 4, 12) {real, imag} */,
  {32'hc2557bb4, 32'h40eca450} /* (6, 4, 11) {real, imag} */,
  {32'hc2f4b48a, 32'h41f10477} /* (6, 4, 10) {real, imag} */,
  {32'h41c170d4, 32'hc0a92558} /* (6, 4, 9) {real, imag} */,
  {32'h42fe342e, 32'h00000000} /* (6, 4, 8) {real, imag} */,
  {32'h41c170d4, 32'h40a92558} /* (6, 4, 7) {real, imag} */,
  {32'hc2f4b48a, 32'hc1f10477} /* (6, 4, 6) {real, imag} */,
  {32'hc2557bb4, 32'hc0eca450} /* (6, 4, 5) {real, imag} */,
  {32'h41916808, 32'hc34ffed2} /* (6, 4, 4) {real, imag} */,
  {32'h42a0f8d7, 32'h427eea54} /* (6, 4, 3) {real, imag} */,
  {32'hc1308b0b, 32'h435d3dcb} /* (6, 4, 2) {real, imag} */,
  {32'hc350c289, 32'h4292d272} /* (6, 4, 1) {real, imag} */,
  {32'hc376a1a2, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'hc2af89fe, 32'hc32054ce} /* (6, 3, 15) {real, imag} */,
  {32'hc2dbea1a, 32'hc2b0a54e} /* (6, 3, 14) {real, imag} */,
  {32'h422cd7ea, 32'h422b3e70} /* (6, 3, 13) {real, imag} */,
  {32'hc2c4ccde, 32'h4315d0f2} /* (6, 3, 12) {real, imag} */,
  {32'hc31ffb3a, 32'h42611cdc} /* (6, 3, 11) {real, imag} */,
  {32'h433cc7d0, 32'hc28844ca} /* (6, 3, 10) {real, imag} */,
  {32'h41d3f615, 32'hc2f03260} /* (6, 3, 9) {real, imag} */,
  {32'hc28cd3f1, 32'h00000000} /* (6, 3, 8) {real, imag} */,
  {32'h41d3f615, 32'h42f03260} /* (6, 3, 7) {real, imag} */,
  {32'h433cc7d0, 32'h428844ca} /* (6, 3, 6) {real, imag} */,
  {32'hc31ffb3a, 32'hc2611cdc} /* (6, 3, 5) {real, imag} */,
  {32'hc2c4ccde, 32'hc315d0f2} /* (6, 3, 4) {real, imag} */,
  {32'h422cd7ea, 32'hc22b3e70} /* (6, 3, 3) {real, imag} */,
  {32'hc2dbea1a, 32'h42b0a54e} /* (6, 3, 2) {real, imag} */,
  {32'hc2af89fe, 32'h432054ce} /* (6, 3, 1) {real, imag} */,
  {32'hc38aa168, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'hc3139082, 32'h429c3318} /* (6, 2, 15) {real, imag} */,
  {32'hc308c8d7, 32'hc30a0cd2} /* (6, 2, 14) {real, imag} */,
  {32'hc2900243, 32'h42c99b04} /* (6, 2, 13) {real, imag} */,
  {32'hc27ae127, 32'hc2decef3} /* (6, 2, 12) {real, imag} */,
  {32'h433d160b, 32'h41598356} /* (6, 2, 11) {real, imag} */,
  {32'h3fc90c00, 32'h42c63bb5} /* (6, 2, 10) {real, imag} */,
  {32'h424efb1a, 32'hc2f23cf2} /* (6, 2, 9) {real, imag} */,
  {32'hc23486c6, 32'h00000000} /* (6, 2, 8) {real, imag} */,
  {32'h424efb1a, 32'h42f23cf2} /* (6, 2, 7) {real, imag} */,
  {32'h3fc90c00, 32'hc2c63bb5} /* (6, 2, 6) {real, imag} */,
  {32'h433d160b, 32'hc1598356} /* (6, 2, 5) {real, imag} */,
  {32'hc27ae127, 32'h42decef3} /* (6, 2, 4) {real, imag} */,
  {32'hc2900243, 32'hc2c99b04} /* (6, 2, 3) {real, imag} */,
  {32'hc308c8d7, 32'h430a0cd2} /* (6, 2, 2) {real, imag} */,
  {32'hc3139082, 32'hc29c3318} /* (6, 2, 1) {real, imag} */,
  {32'hc3ead9c8, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'hc2df723a, 32'h43697f9d} /* (6, 1, 15) {real, imag} */,
  {32'hc36f9366, 32'hc30c8c1a} /* (6, 1, 14) {real, imag} */,
  {32'hc3553f95, 32'hc383cdf4} /* (6, 1, 13) {real, imag} */,
  {32'h430747cd, 32'h43241234} /* (6, 1, 12) {real, imag} */,
  {32'h422bebf4, 32'hc099e9bc} /* (6, 1, 11) {real, imag} */,
  {32'hc2313496, 32'h423da30f} /* (6, 1, 10) {real, imag} */,
  {32'h3fa92a40, 32'hc20612a2} /* (6, 1, 9) {real, imag} */,
  {32'h42a5f75c, 32'h00000000} /* (6, 1, 8) {real, imag} */,
  {32'h3fa92a40, 32'h420612a2} /* (6, 1, 7) {real, imag} */,
  {32'hc2313496, 32'hc23da30f} /* (6, 1, 6) {real, imag} */,
  {32'h422bebf4, 32'h4099e9bc} /* (6, 1, 5) {real, imag} */,
  {32'h430747cd, 32'hc3241234} /* (6, 1, 4) {real, imag} */,
  {32'hc3553f95, 32'h4383cdf4} /* (6, 1, 3) {real, imag} */,
  {32'hc36f9366, 32'h430c8c1a} /* (6, 1, 2) {real, imag} */,
  {32'hc2df723a, 32'hc3697f9d} /* (6, 1, 1) {real, imag} */,
  {32'hc39d3d32, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'hc2b7098c, 32'h42ca4c40} /* (6, 0, 15) {real, imag} */,
  {32'hc296f261, 32'hc2aa606a} /* (6, 0, 14) {real, imag} */,
  {32'h4231c4a4, 32'hc2b22d82} /* (6, 0, 13) {real, imag} */,
  {32'h425126b8, 32'h42fc7382} /* (6, 0, 12) {real, imag} */,
  {32'hc27f52cf, 32'h410573b0} /* (6, 0, 11) {real, imag} */,
  {32'h3f6da4e0, 32'hc2a31115} /* (6, 0, 10) {real, imag} */,
  {32'h423408e7, 32'h42110b58} /* (6, 0, 9) {real, imag} */,
  {32'hc20932ac, 32'h00000000} /* (6, 0, 8) {real, imag} */,
  {32'h423408e7, 32'hc2110b58} /* (6, 0, 7) {real, imag} */,
  {32'h3f6da4e0, 32'h42a31115} /* (6, 0, 6) {real, imag} */,
  {32'hc27f52cf, 32'hc10573b0} /* (6, 0, 5) {real, imag} */,
  {32'h425126b8, 32'hc2fc7382} /* (6, 0, 4) {real, imag} */,
  {32'h4231c4a4, 32'h42b22d82} /* (6, 0, 3) {real, imag} */,
  {32'hc296f261, 32'h42aa606a} /* (6, 0, 2) {real, imag} */,
  {32'hc2b7098c, 32'hc2ca4c40} /* (6, 0, 1) {real, imag} */,
  {32'hc3526efe, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'hc2dd92fc, 32'h432d0b16} /* (5, 15, 15) {real, imag} */,
  {32'hc2b81d0a, 32'hc188a3fb} /* (5, 15, 14) {real, imag} */,
  {32'h41e4aec0, 32'hc1ae177e} /* (5, 15, 13) {real, imag} */,
  {32'h4323bd7a, 32'h43011215} /* (5, 15, 12) {real, imag} */,
  {32'h42e5998e, 32'h429f5e43} /* (5, 15, 11) {real, imag} */,
  {32'hc1bf3d51, 32'h41a6b53e} /* (5, 15, 10) {real, imag} */,
  {32'h423061b0, 32'hc0da594c} /* (5, 15, 9) {real, imag} */,
  {32'h42b9f850, 32'h00000000} /* (5, 15, 8) {real, imag} */,
  {32'h423061b0, 32'h40da594c} /* (5, 15, 7) {real, imag} */,
  {32'hc1bf3d51, 32'hc1a6b53e} /* (5, 15, 6) {real, imag} */,
  {32'h42e5998e, 32'hc29f5e43} /* (5, 15, 5) {real, imag} */,
  {32'h4323bd7a, 32'hc3011215} /* (5, 15, 4) {real, imag} */,
  {32'h41e4aec0, 32'h41ae177e} /* (5, 15, 3) {real, imag} */,
  {32'hc2b81d0a, 32'h4188a3fb} /* (5, 15, 2) {real, imag} */,
  {32'hc2dd92fc, 32'hc32d0b16} /* (5, 15, 1) {real, imag} */,
  {32'hc3c70fc2, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'hc2866fa4, 32'h42e43d53} /* (5, 14, 15) {real, imag} */,
  {32'h430919bc, 32'hc2a8e99f} /* (5, 14, 14) {real, imag} */,
  {32'h433c2786, 32'hc110ced4} /* (5, 14, 13) {real, imag} */,
  {32'h42c28715, 32'h42789de1} /* (5, 14, 12) {real, imag} */,
  {32'h42ca9f6e, 32'h42f47544} /* (5, 14, 11) {real, imag} */,
  {32'h418b3f3c, 32'h432d77a4} /* (5, 14, 10) {real, imag} */,
  {32'h42f7dfb0, 32'h422ae515} /* (5, 14, 9) {real, imag} */,
  {32'h3f85b500, 32'h00000000} /* (5, 14, 8) {real, imag} */,
  {32'h42f7dfb0, 32'hc22ae515} /* (5, 14, 7) {real, imag} */,
  {32'h418b3f3c, 32'hc32d77a4} /* (5, 14, 6) {real, imag} */,
  {32'h42ca9f6e, 32'hc2f47544} /* (5, 14, 5) {real, imag} */,
  {32'h42c28715, 32'hc2789de1} /* (5, 14, 4) {real, imag} */,
  {32'h433c2786, 32'h4110ced4} /* (5, 14, 3) {real, imag} */,
  {32'h430919bc, 32'h42a8e99f} /* (5, 14, 2) {real, imag} */,
  {32'hc2866fa4, 32'hc2e43d53} /* (5, 14, 1) {real, imag} */,
  {32'hc3d3590c, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hc242b8ec, 32'h42d4bbac} /* (5, 13, 15) {real, imag} */,
  {32'h42c6f24e, 32'hc25c958c} /* (5, 13, 14) {real, imag} */,
  {32'hc1a4c3c0, 32'h41224b0c} /* (5, 13, 13) {real, imag} */,
  {32'hc31568a6, 32'hc305434a} /* (5, 13, 12) {real, imag} */,
  {32'h42589034, 32'hc10578a4} /* (5, 13, 11) {real, imag} */,
  {32'h42e82b14, 32'hc23f9681} /* (5, 13, 10) {real, imag} */,
  {32'hc208c64e, 32'h4155b1e8} /* (5, 13, 9) {real, imag} */,
  {32'hc22a827b, 32'h00000000} /* (5, 13, 8) {real, imag} */,
  {32'hc208c64e, 32'hc155b1e8} /* (5, 13, 7) {real, imag} */,
  {32'h42e82b14, 32'h423f9681} /* (5, 13, 6) {real, imag} */,
  {32'h42589034, 32'h410578a4} /* (5, 13, 5) {real, imag} */,
  {32'hc31568a6, 32'h4305434a} /* (5, 13, 4) {real, imag} */,
  {32'hc1a4c3c0, 32'hc1224b0c} /* (5, 13, 3) {real, imag} */,
  {32'h42c6f24e, 32'h425c958c} /* (5, 13, 2) {real, imag} */,
  {32'hc242b8ec, 32'hc2d4bbac} /* (5, 13, 1) {real, imag} */,
  {32'hc40ea07d, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'h42ecf0da, 32'h431fff60} /* (5, 12, 15) {real, imag} */,
  {32'hc223f0ae, 32'hc3458adf} /* (5, 12, 14) {real, imag} */,
  {32'hc32be070, 32'h4103fd40} /* (5, 12, 13) {real, imag} */,
  {32'hc2b39588, 32'hc22770a4} /* (5, 12, 12) {real, imag} */,
  {32'hc0bb1160, 32'h4336bedc} /* (5, 12, 11) {real, imag} */,
  {32'h4285652d, 32'hc2c94ab4} /* (5, 12, 10) {real, imag} */,
  {32'h42a6e931, 32'hc23a3a2d} /* (5, 12, 9) {real, imag} */,
  {32'hc182836d, 32'h00000000} /* (5, 12, 8) {real, imag} */,
  {32'h42a6e931, 32'h423a3a2d} /* (5, 12, 7) {real, imag} */,
  {32'h4285652d, 32'h42c94ab4} /* (5, 12, 6) {real, imag} */,
  {32'hc0bb1160, 32'hc336bedc} /* (5, 12, 5) {real, imag} */,
  {32'hc2b39588, 32'h422770a4} /* (5, 12, 4) {real, imag} */,
  {32'hc32be070, 32'hc103fd40} /* (5, 12, 3) {real, imag} */,
  {32'hc223f0ae, 32'h43458adf} /* (5, 12, 2) {real, imag} */,
  {32'h42ecf0da, 32'hc31fff60} /* (5, 12, 1) {real, imag} */,
  {32'hc3dea7dd, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h42a1e55d, 32'h43980962} /* (5, 11, 15) {real, imag} */,
  {32'hc28807c2, 32'hc29ed611} /* (5, 11, 14) {real, imag} */,
  {32'h4327f53a, 32'h423cf6cd} /* (5, 11, 13) {real, imag} */,
  {32'hc14b5fba, 32'hc36586c7} /* (5, 11, 12) {real, imag} */,
  {32'hc2a21126, 32'hc302ebd2} /* (5, 11, 11) {real, imag} */,
  {32'hc27bc0fc, 32'h42e252ec} /* (5, 11, 10) {real, imag} */,
  {32'hc18e2ed2, 32'h418d84d4} /* (5, 11, 9) {real, imag} */,
  {32'hc25ae07a, 32'h00000000} /* (5, 11, 8) {real, imag} */,
  {32'hc18e2ed2, 32'hc18d84d4} /* (5, 11, 7) {real, imag} */,
  {32'hc27bc0fc, 32'hc2e252ec} /* (5, 11, 6) {real, imag} */,
  {32'hc2a21126, 32'h4302ebd2} /* (5, 11, 5) {real, imag} */,
  {32'hc14b5fba, 32'h436586c7} /* (5, 11, 4) {real, imag} */,
  {32'h4327f53a, 32'hc23cf6cd} /* (5, 11, 3) {real, imag} */,
  {32'hc28807c2, 32'h429ed611} /* (5, 11, 2) {real, imag} */,
  {32'h42a1e55d, 32'hc3980962} /* (5, 11, 1) {real, imag} */,
  {32'hc3a0ba24, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'h41b838b0, 32'h43bd839c} /* (5, 10, 15) {real, imag} */,
  {32'hc056f440, 32'h422ab6de} /* (5, 10, 14) {real, imag} */,
  {32'h43134a89, 32'hc104a2d8} /* (5, 10, 13) {real, imag} */,
  {32'hc1592dec, 32'h4218ee4b} /* (5, 10, 12) {real, imag} */,
  {32'hc240494a, 32'hc2352a9e} /* (5, 10, 11) {real, imag} */,
  {32'hc187b90f, 32'h41f496d6} /* (5, 10, 10) {real, imag} */,
  {32'hc1d3a0fe, 32'hc28c4d18} /* (5, 10, 9) {real, imag} */,
  {32'h42136a93, 32'h00000000} /* (5, 10, 8) {real, imag} */,
  {32'hc1d3a0fe, 32'h428c4d18} /* (5, 10, 7) {real, imag} */,
  {32'hc187b90f, 32'hc1f496d6} /* (5, 10, 6) {real, imag} */,
  {32'hc240494a, 32'h42352a9e} /* (5, 10, 5) {real, imag} */,
  {32'hc1592dec, 32'hc218ee4b} /* (5, 10, 4) {real, imag} */,
  {32'h43134a89, 32'h4104a2d8} /* (5, 10, 3) {real, imag} */,
  {32'hc056f440, 32'hc22ab6de} /* (5, 10, 2) {real, imag} */,
  {32'h41b838b0, 32'hc3bd839c} /* (5, 10, 1) {real, imag} */,
  {32'hc2862014, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'hbfcbb580, 32'h4290de78} /* (5, 9, 15) {real, imag} */,
  {32'h42a8069c, 32'hc04c8600} /* (5, 9, 14) {real, imag} */,
  {32'hc1e52215, 32'hc3045e98} /* (5, 9, 13) {real, imag} */,
  {32'hc2ce4adc, 32'h42a9ea2e} /* (5, 9, 12) {real, imag} */,
  {32'h42446304, 32'h4322f018} /* (5, 9, 11) {real, imag} */,
  {32'h41e4f0c6, 32'hc30b54a1} /* (5, 9, 10) {real, imag} */,
  {32'h41b79794, 32'hc24e7426} /* (5, 9, 9) {real, imag} */,
  {32'hc30dfdeb, 32'h00000000} /* (5, 9, 8) {real, imag} */,
  {32'h41b79794, 32'h424e7426} /* (5, 9, 7) {real, imag} */,
  {32'h41e4f0c6, 32'h430b54a1} /* (5, 9, 6) {real, imag} */,
  {32'h42446304, 32'hc322f018} /* (5, 9, 5) {real, imag} */,
  {32'hc2ce4adc, 32'hc2a9ea2e} /* (5, 9, 4) {real, imag} */,
  {32'hc1e52215, 32'h43045e98} /* (5, 9, 3) {real, imag} */,
  {32'h42a8069c, 32'h404c8600} /* (5, 9, 2) {real, imag} */,
  {32'hbfcbb580, 32'hc290de78} /* (5, 9, 1) {real, imag} */,
  {32'h41231da0, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'hc1cd72ca, 32'h43648ff6} /* (5, 8, 15) {real, imag} */,
  {32'h437f81c3, 32'hc192a434} /* (5, 8, 14) {real, imag} */,
  {32'h42b12a61, 32'hc32531ee} /* (5, 8, 13) {real, imag} */,
  {32'hc1d18be8, 32'hc2a820fe} /* (5, 8, 12) {real, imag} */,
  {32'hc216b42f, 32'h43125342} /* (5, 8, 11) {real, imag} */,
  {32'hc26c3754, 32'hc2a9233f} /* (5, 8, 10) {real, imag} */,
  {32'h42903d40, 32'hc1e624c4} /* (5, 8, 9) {real, imag} */,
  {32'h41a31be1, 32'h00000000} /* (5, 8, 8) {real, imag} */,
  {32'h42903d40, 32'h41e624c4} /* (5, 8, 7) {real, imag} */,
  {32'hc26c3754, 32'h42a9233f} /* (5, 8, 6) {real, imag} */,
  {32'hc216b42f, 32'hc3125342} /* (5, 8, 5) {real, imag} */,
  {32'hc1d18be8, 32'h42a820fe} /* (5, 8, 4) {real, imag} */,
  {32'h42b12a61, 32'h432531ee} /* (5, 8, 3) {real, imag} */,
  {32'h437f81c3, 32'h4192a434} /* (5, 8, 2) {real, imag} */,
  {32'hc1cd72ca, 32'hc3648ff6} /* (5, 8, 1) {real, imag} */,
  {32'h41339e20, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'hc28ae46c, 32'h43964fd1} /* (5, 7, 15) {real, imag} */,
  {32'h4380c3a4, 32'hc31b31f3} /* (5, 7, 14) {real, imag} */,
  {32'h41e22233, 32'hc31f11e8} /* (5, 7, 13) {real, imag} */,
  {32'hc2e70c68, 32'h431010cb} /* (5, 7, 12) {real, imag} */,
  {32'hc1b50eb8, 32'h41e33730} /* (5, 7, 11) {real, imag} */,
  {32'hc23dc0dd, 32'hc168d91c} /* (5, 7, 10) {real, imag} */,
  {32'hc329e1be, 32'h42d97b71} /* (5, 7, 9) {real, imag} */,
  {32'h417292d0, 32'h00000000} /* (5, 7, 8) {real, imag} */,
  {32'hc329e1be, 32'hc2d97b71} /* (5, 7, 7) {real, imag} */,
  {32'hc23dc0dd, 32'h4168d91c} /* (5, 7, 6) {real, imag} */,
  {32'hc1b50eb8, 32'hc1e33730} /* (5, 7, 5) {real, imag} */,
  {32'hc2e70c68, 32'hc31010cb} /* (5, 7, 4) {real, imag} */,
  {32'h41e22233, 32'h431f11e8} /* (5, 7, 3) {real, imag} */,
  {32'h4380c3a4, 32'h431b31f3} /* (5, 7, 2) {real, imag} */,
  {32'hc28ae46c, 32'hc3964fd1} /* (5, 7, 1) {real, imag} */,
  {32'hc340ff2a, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'hc336810c, 32'h41cd3f08} /* (5, 6, 15) {real, imag} */,
  {32'h42f26c60, 32'hc35dd5d0} /* (5, 6, 14) {real, imag} */,
  {32'h430602bf, 32'hc3372b64} /* (5, 6, 13) {real, imag} */,
  {32'h417e660c, 32'h414d7091} /* (5, 6, 12) {real, imag} */,
  {32'hc145cf2a, 32'h42ce092d} /* (5, 6, 11) {real, imag} */,
  {32'h4235ab48, 32'hc1c96156} /* (5, 6, 10) {real, imag} */,
  {32'hbf433730, 32'h431af66c} /* (5, 6, 9) {real, imag} */,
  {32'hc0084150, 32'h00000000} /* (5, 6, 8) {real, imag} */,
  {32'hbf433730, 32'hc31af66c} /* (5, 6, 7) {real, imag} */,
  {32'h4235ab48, 32'h41c96156} /* (5, 6, 6) {real, imag} */,
  {32'hc145cf2a, 32'hc2ce092d} /* (5, 6, 5) {real, imag} */,
  {32'h417e660c, 32'hc14d7091} /* (5, 6, 4) {real, imag} */,
  {32'h430602bf, 32'h43372b64} /* (5, 6, 3) {real, imag} */,
  {32'h42f26c60, 32'h435dd5d0} /* (5, 6, 2) {real, imag} */,
  {32'hc336810c, 32'hc1cd3f08} /* (5, 6, 1) {real, imag} */,
  {32'hc3f8c0a9, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'hc36d79ca, 32'hc267e3d0} /* (5, 5, 15) {real, imag} */,
  {32'h41992571, 32'hc337dffc} /* (5, 5, 14) {real, imag} */,
  {32'h403c7400, 32'hc2771f7b} /* (5, 5, 13) {real, imag} */,
  {32'hc0e7200c, 32'hc2af417e} /* (5, 5, 12) {real, imag} */,
  {32'h41ebc7d9, 32'hc18729d0} /* (5, 5, 11) {real, imag} */,
  {32'h430704ed, 32'h4196b492} /* (5, 5, 10) {real, imag} */,
  {32'h43034f96, 32'hc11977a8} /* (5, 5, 9) {real, imag} */,
  {32'h430954b0, 32'h00000000} /* (5, 5, 8) {real, imag} */,
  {32'h43034f96, 32'h411977a8} /* (5, 5, 7) {real, imag} */,
  {32'h430704ed, 32'hc196b492} /* (5, 5, 6) {real, imag} */,
  {32'h41ebc7d9, 32'h418729d0} /* (5, 5, 5) {real, imag} */,
  {32'hc0e7200c, 32'h42af417e} /* (5, 5, 4) {real, imag} */,
  {32'h403c7400, 32'h42771f7b} /* (5, 5, 3) {real, imag} */,
  {32'h41992571, 32'h4337dffc} /* (5, 5, 2) {real, imag} */,
  {32'hc36d79ca, 32'h4267e3d0} /* (5, 5, 1) {real, imag} */,
  {32'hc40776d0, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'hc3696cfb, 32'hc29521d0} /* (5, 4, 15) {real, imag} */,
  {32'h4256d72a, 32'hc334d4fd} /* (5, 4, 14) {real, imag} */,
  {32'h4313f81c, 32'hc33c6bf9} /* (5, 4, 13) {real, imag} */,
  {32'hc314503e, 32'h42d587f0} /* (5, 4, 12) {real, imag} */,
  {32'hc31a8559, 32'hc1ef2354} /* (5, 4, 11) {real, imag} */,
  {32'hc2f3f4e5, 32'hc28bb6dc} /* (5, 4, 10) {real, imag} */,
  {32'h41528790, 32'h41866510} /* (5, 4, 9) {real, imag} */,
  {32'hc207aa1a, 32'h00000000} /* (5, 4, 8) {real, imag} */,
  {32'h41528790, 32'hc1866510} /* (5, 4, 7) {real, imag} */,
  {32'hc2f3f4e5, 32'h428bb6dc} /* (5, 4, 6) {real, imag} */,
  {32'hc31a8559, 32'h41ef2354} /* (5, 4, 5) {real, imag} */,
  {32'hc314503e, 32'hc2d587f0} /* (5, 4, 4) {real, imag} */,
  {32'h4313f81c, 32'h433c6bf9} /* (5, 4, 3) {real, imag} */,
  {32'h4256d72a, 32'h4334d4fd} /* (5, 4, 2) {real, imag} */,
  {32'hc3696cfb, 32'h429521d0} /* (5, 4, 1) {real, imag} */,
  {32'hc3a5a321, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'hc2cda748, 32'hc3a90453} /* (5, 3, 15) {real, imag} */,
  {32'h41c61218, 32'hc23cccdc} /* (5, 3, 14) {real, imag} */,
  {32'h4318151e, 32'h42af374e} /* (5, 3, 13) {real, imag} */,
  {32'hc335612e, 32'h420af34f} /* (5, 3, 12) {real, imag} */,
  {32'hc0ffe61c, 32'h42b050a8} /* (5, 3, 11) {real, imag} */,
  {32'h4326bd6e, 32'h41cc153a} /* (5, 3, 10) {real, imag} */,
  {32'h3ffe1880, 32'h42f6908f} /* (5, 3, 9) {real, imag} */,
  {32'hc31c3ccc, 32'h00000000} /* (5, 3, 8) {real, imag} */,
  {32'h3ffe1880, 32'hc2f6908f} /* (5, 3, 7) {real, imag} */,
  {32'h4326bd6e, 32'hc1cc153a} /* (5, 3, 6) {real, imag} */,
  {32'hc0ffe61c, 32'hc2b050a8} /* (5, 3, 5) {real, imag} */,
  {32'hc335612e, 32'hc20af34f} /* (5, 3, 4) {real, imag} */,
  {32'h4318151e, 32'hc2af374e} /* (5, 3, 3) {real, imag} */,
  {32'h41c61218, 32'h423cccdc} /* (5, 3, 2) {real, imag} */,
  {32'hc2cda748, 32'h43a90453} /* (5, 3, 1) {real, imag} */,
  {32'hc3d8d002, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'hc376306c, 32'h42e52089} /* (5, 2, 15) {real, imag} */,
  {32'hc33299f4, 32'hc30bbbc2} /* (5, 2, 14) {real, imag} */,
  {32'hc2c8df94, 32'h41aeeb2a} /* (5, 2, 13) {real, imag} */,
  {32'h4342a7cc, 32'h42446d9b} /* (5, 2, 12) {real, imag} */,
  {32'hc29567d0, 32'hbf3a40c0} /* (5, 2, 11) {real, imag} */,
  {32'h42c872b5, 32'h41e635c0} /* (5, 2, 10) {real, imag} */,
  {32'h42a7a1b2, 32'hc3095cb7} /* (5, 2, 9) {real, imag} */,
  {32'hc3430554, 32'h00000000} /* (5, 2, 8) {real, imag} */,
  {32'h42a7a1b2, 32'h43095cb7} /* (5, 2, 7) {real, imag} */,
  {32'h42c872b5, 32'hc1e635c0} /* (5, 2, 6) {real, imag} */,
  {32'hc29567d0, 32'h3f3a40c0} /* (5, 2, 5) {real, imag} */,
  {32'h4342a7cc, 32'hc2446d9b} /* (5, 2, 4) {real, imag} */,
  {32'hc2c8df94, 32'hc1aeeb2a} /* (5, 2, 3) {real, imag} */,
  {32'hc33299f4, 32'h430bbbc2} /* (5, 2, 2) {real, imag} */,
  {32'hc376306c, 32'hc2e52089} /* (5, 2, 1) {real, imag} */,
  {32'hc3cdd872, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'hc37629b6, 32'hc2f89f48} /* (5, 1, 15) {real, imag} */,
  {32'hc305ec61, 32'hc277bffe} /* (5, 1, 14) {real, imag} */,
  {32'h4203faa1, 32'hc2949a54} /* (5, 1, 13) {real, imag} */,
  {32'hc1f586b0, 32'h437d073d} /* (5, 1, 12) {real, imag} */,
  {32'h4120a4d0, 32'h4133cb50} /* (5, 1, 11) {real, imag} */,
  {32'hc28dc6c3, 32'h404efc90} /* (5, 1, 10) {real, imag} */,
  {32'hc1b657e8, 32'h419c9f2d} /* (5, 1, 9) {real, imag} */,
  {32'h42ae7d0c, 32'h00000000} /* (5, 1, 8) {real, imag} */,
  {32'hc1b657e8, 32'hc19c9f2d} /* (5, 1, 7) {real, imag} */,
  {32'hc28dc6c3, 32'hc04efc90} /* (5, 1, 6) {real, imag} */,
  {32'h4120a4d0, 32'hc133cb50} /* (5, 1, 5) {real, imag} */,
  {32'hc1f586b0, 32'hc37d073d} /* (5, 1, 4) {real, imag} */,
  {32'h4203faa1, 32'h42949a54} /* (5, 1, 3) {real, imag} */,
  {32'hc305ec61, 32'h4277bffe} /* (5, 1, 2) {real, imag} */,
  {32'hc37629b6, 32'h42f89f48} /* (5, 1, 1) {real, imag} */,
  {32'hc3b82760, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'hc2f87baa, 32'h42bbf833} /* (5, 0, 15) {real, imag} */,
  {32'h40170a40, 32'hc2a7dd55} /* (5, 0, 14) {real, imag} */,
  {32'hc2a8e6e1, 32'hc0eaaeb0} /* (5, 0, 13) {real, imag} */,
  {32'hc0373740, 32'hc23bf52f} /* (5, 0, 12) {real, imag} */,
  {32'hc27a1b6b, 32'hc12c0680} /* (5, 0, 11) {real, imag} */,
  {32'h431670df, 32'hc001b520} /* (5, 0, 10) {real, imag} */,
  {32'hc1edfc7a, 32'h3f8761f8} /* (5, 0, 9) {real, imag} */,
  {32'hc1e5070b, 32'h00000000} /* (5, 0, 8) {real, imag} */,
  {32'hc1edfc7a, 32'hbf8761f8} /* (5, 0, 7) {real, imag} */,
  {32'h431670df, 32'h4001b520} /* (5, 0, 6) {real, imag} */,
  {32'hc27a1b6b, 32'h412c0680} /* (5, 0, 5) {real, imag} */,
  {32'hc0373740, 32'h423bf52f} /* (5, 0, 4) {real, imag} */,
  {32'hc2a8e6e1, 32'h40eaaeb0} /* (5, 0, 3) {real, imag} */,
  {32'h40170a40, 32'h42a7dd55} /* (5, 0, 2) {real, imag} */,
  {32'hc2f87baa, 32'hc2bbf833} /* (5, 0, 1) {real, imag} */,
  {32'hc39ec29f, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hc29b5c41, 32'h41d7fe26} /* (4, 15, 15) {real, imag} */,
  {32'hc3201906, 32'hc247c2ba} /* (4, 15, 14) {real, imag} */,
  {32'h425dc218, 32'h41e71dd6} /* (4, 15, 13) {real, imag} */,
  {32'h41f9873e, 32'h4263bb3e} /* (4, 15, 12) {real, imag} */,
  {32'h41b3d450, 32'hc2124093} /* (4, 15, 11) {real, imag} */,
  {32'h41407fa0, 32'hc1bf2744} /* (4, 15, 10) {real, imag} */,
  {32'hc1a7d21e, 32'h4106921e} /* (4, 15, 9) {real, imag} */,
  {32'hc1a9e807, 32'h00000000} /* (4, 15, 8) {real, imag} */,
  {32'hc1a7d21e, 32'hc106921e} /* (4, 15, 7) {real, imag} */,
  {32'h41407fa0, 32'h41bf2744} /* (4, 15, 6) {real, imag} */,
  {32'h41b3d450, 32'h42124093} /* (4, 15, 5) {real, imag} */,
  {32'h41f9873e, 32'hc263bb3e} /* (4, 15, 4) {real, imag} */,
  {32'h425dc218, 32'hc1e71dd6} /* (4, 15, 3) {real, imag} */,
  {32'hc3201906, 32'h4247c2ba} /* (4, 15, 2) {real, imag} */,
  {32'hc29b5c41, 32'hc1d7fe26} /* (4, 15, 1) {real, imag} */,
  {32'hc31f0152, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'h4284cf70, 32'h4370aabe} /* (4, 14, 15) {real, imag} */,
  {32'hc2041d43, 32'hc1ed26ca} /* (4, 14, 14) {real, imag} */,
  {32'h431cc29a, 32'h4343f250} /* (4, 14, 13) {real, imag} */,
  {32'h42c5857c, 32'hc1cd42f8} /* (4, 14, 12) {real, imag} */,
  {32'h42759192, 32'h426955fa} /* (4, 14, 11) {real, imag} */,
  {32'h42674bfa, 32'h4239ee96} /* (4, 14, 10) {real, imag} */,
  {32'hc23d89ee, 32'hc2913920} /* (4, 14, 9) {real, imag} */,
  {32'hc26a12d1, 32'h00000000} /* (4, 14, 8) {real, imag} */,
  {32'hc23d89ee, 32'h42913920} /* (4, 14, 7) {real, imag} */,
  {32'h42674bfa, 32'hc239ee96} /* (4, 14, 6) {real, imag} */,
  {32'h42759192, 32'hc26955fa} /* (4, 14, 5) {real, imag} */,
  {32'h42c5857c, 32'h41cd42f8} /* (4, 14, 4) {real, imag} */,
  {32'h431cc29a, 32'hc343f250} /* (4, 14, 3) {real, imag} */,
  {32'hc2041d43, 32'h41ed26ca} /* (4, 14, 2) {real, imag} */,
  {32'h4284cf70, 32'hc370aabe} /* (4, 14, 1) {real, imag} */,
  {32'hc3cb0e22, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'hc25d0c80, 32'h4391155a} /* (4, 13, 15) {real, imag} */,
  {32'hc21f5b9a, 32'hc2fa72af} /* (4, 13, 14) {real, imag} */,
  {32'hc170ebb4, 32'h43286d36} /* (4, 13, 13) {real, imag} */,
  {32'h431eacd4, 32'hc32a051b} /* (4, 13, 12) {real, imag} */,
  {32'h42ad9f99, 32'hc269652a} /* (4, 13, 11) {real, imag} */,
  {32'hc28349c5, 32'hc22c3bb0} /* (4, 13, 10) {real, imag} */,
  {32'hc21d7642, 32'h42f83281} /* (4, 13, 9) {real, imag} */,
  {32'h42cbfe35, 32'h00000000} /* (4, 13, 8) {real, imag} */,
  {32'hc21d7642, 32'hc2f83281} /* (4, 13, 7) {real, imag} */,
  {32'hc28349c5, 32'h422c3bb0} /* (4, 13, 6) {real, imag} */,
  {32'h42ad9f99, 32'h4269652a} /* (4, 13, 5) {real, imag} */,
  {32'h431eacd4, 32'h432a051b} /* (4, 13, 4) {real, imag} */,
  {32'hc170ebb4, 32'hc3286d36} /* (4, 13, 3) {real, imag} */,
  {32'hc21f5b9a, 32'h42fa72af} /* (4, 13, 2) {real, imag} */,
  {32'hc25d0c80, 32'hc391155a} /* (4, 13, 1) {real, imag} */,
  {32'hc367ce66, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'hc187c188, 32'h431d3ec4} /* (4, 12, 15) {real, imag} */,
  {32'hc2ea009a, 32'hc30a1fe4} /* (4, 12, 14) {real, imag} */,
  {32'h4247efea, 32'h42a7d84d} /* (4, 12, 13) {real, imag} */,
  {32'h42535e3a, 32'h43896238} /* (4, 12, 12) {real, imag} */,
  {32'hc13e26f4, 32'hc26e9c2d} /* (4, 12, 11) {real, imag} */,
  {32'h42dd5a67, 32'hc1440cbc} /* (4, 12, 10) {real, imag} */,
  {32'hc297e42e, 32'h42c739de} /* (4, 12, 9) {real, imag} */,
  {32'hc2f4553e, 32'h00000000} /* (4, 12, 8) {real, imag} */,
  {32'hc297e42e, 32'hc2c739de} /* (4, 12, 7) {real, imag} */,
  {32'h42dd5a67, 32'h41440cbc} /* (4, 12, 6) {real, imag} */,
  {32'hc13e26f4, 32'h426e9c2d} /* (4, 12, 5) {real, imag} */,
  {32'h42535e3a, 32'hc3896238} /* (4, 12, 4) {real, imag} */,
  {32'h4247efea, 32'hc2a7d84d} /* (4, 12, 3) {real, imag} */,
  {32'hc2ea009a, 32'h430a1fe4} /* (4, 12, 2) {real, imag} */,
  {32'hc187c188, 32'hc31d3ec4} /* (4, 12, 1) {real, imag} */,
  {32'hc304e54c, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'hc0441600, 32'h43b241b3} /* (4, 11, 15) {real, imag} */,
  {32'hc2a4f168, 32'hc37f568e} /* (4, 11, 14) {real, imag} */,
  {32'h42e23ee4, 32'h42c3901a} /* (4, 11, 13) {real, imag} */,
  {32'hc23f415b, 32'h4310357e} /* (4, 11, 12) {real, imag} */,
  {32'h42e43439, 32'hc19f2a8b} /* (4, 11, 11) {real, imag} */,
  {32'hc24ff359, 32'hc2c0ebee} /* (4, 11, 10) {real, imag} */,
  {32'h42e58710, 32'h41bcc492} /* (4, 11, 9) {real, imag} */,
  {32'hc253576b, 32'h00000000} /* (4, 11, 8) {real, imag} */,
  {32'h42e58710, 32'hc1bcc492} /* (4, 11, 7) {real, imag} */,
  {32'hc24ff359, 32'h42c0ebee} /* (4, 11, 6) {real, imag} */,
  {32'h42e43439, 32'h419f2a8b} /* (4, 11, 5) {real, imag} */,
  {32'hc23f415b, 32'hc310357e} /* (4, 11, 4) {real, imag} */,
  {32'h42e23ee4, 32'hc2c3901a} /* (4, 11, 3) {real, imag} */,
  {32'hc2a4f168, 32'h437f568e} /* (4, 11, 2) {real, imag} */,
  {32'hc0441600, 32'hc3b241b3} /* (4, 11, 1) {real, imag} */,
  {32'hc10fdba8, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'hc04e8240, 32'h42c33efc} /* (4, 10, 15) {real, imag} */,
  {32'hc2b3f9b7, 32'hc30a5678} /* (4, 10, 14) {real, imag} */,
  {32'h4277e1ab, 32'hc1acc4f0} /* (4, 10, 13) {real, imag} */,
  {32'h42d567ce, 32'h419c3954} /* (4, 10, 12) {real, imag} */,
  {32'h41d67af4, 32'h423fbf5e} /* (4, 10, 11) {real, imag} */,
  {32'h428bd754, 32'hc29684c1} /* (4, 10, 10) {real, imag} */,
  {32'hc2601d0f, 32'h423e8578} /* (4, 10, 9) {real, imag} */,
  {32'h42a69c46, 32'h00000000} /* (4, 10, 8) {real, imag} */,
  {32'hc2601d0f, 32'hc23e8578} /* (4, 10, 7) {real, imag} */,
  {32'h428bd754, 32'h429684c1} /* (4, 10, 6) {real, imag} */,
  {32'h41d67af4, 32'hc23fbf5e} /* (4, 10, 5) {real, imag} */,
  {32'h42d567ce, 32'hc19c3954} /* (4, 10, 4) {real, imag} */,
  {32'h4277e1ab, 32'h41acc4f0} /* (4, 10, 3) {real, imag} */,
  {32'hc2b3f9b7, 32'h430a5678} /* (4, 10, 2) {real, imag} */,
  {32'hc04e8240, 32'hc2c33efc} /* (4, 10, 1) {real, imag} */,
  {32'hbed2b800, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'h41831d10, 32'h4284495e} /* (4, 9, 15) {real, imag} */,
  {32'h432e0638, 32'hc22c68a4} /* (4, 9, 14) {real, imag} */,
  {32'hc20a5c6e, 32'h4236e794} /* (4, 9, 13) {real, imag} */,
  {32'h4278db25, 32'h41c568a0} /* (4, 9, 12) {real, imag} */,
  {32'h4289d776, 32'h42e2f8d5} /* (4, 9, 11) {real, imag} */,
  {32'h42f0da62, 32'hc2ffe37d} /* (4, 9, 10) {real, imag} */,
  {32'h41ac4a90, 32'h42908c8a} /* (4, 9, 9) {real, imag} */,
  {32'hc258663e, 32'h00000000} /* (4, 9, 8) {real, imag} */,
  {32'h41ac4a90, 32'hc2908c8a} /* (4, 9, 7) {real, imag} */,
  {32'h42f0da62, 32'h42ffe37d} /* (4, 9, 6) {real, imag} */,
  {32'h4289d776, 32'hc2e2f8d5} /* (4, 9, 5) {real, imag} */,
  {32'h4278db25, 32'hc1c568a0} /* (4, 9, 4) {real, imag} */,
  {32'hc20a5c6e, 32'hc236e794} /* (4, 9, 3) {real, imag} */,
  {32'h432e0638, 32'h422c68a4} /* (4, 9, 2) {real, imag} */,
  {32'h41831d10, 32'hc284495e} /* (4, 9, 1) {real, imag} */,
  {32'hc354f67d, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'h42bc10ed, 32'h4298ade1} /* (4, 8, 15) {real, imag} */,
  {32'h43338e0a, 32'hc3599bd8} /* (4, 8, 14) {real, imag} */,
  {32'h4376310f, 32'hc291eded} /* (4, 8, 13) {real, imag} */,
  {32'hc2eb928c, 32'h42a080a2} /* (4, 8, 12) {real, imag} */,
  {32'h4203ee9c, 32'hc1bbc790} /* (4, 8, 11) {real, imag} */,
  {32'hc2e6fbe3, 32'hc21e4dcf} /* (4, 8, 10) {real, imag} */,
  {32'hc18532ec, 32'h40db92b8} /* (4, 8, 9) {real, imag} */,
  {32'hc2a5b4f1, 32'h00000000} /* (4, 8, 8) {real, imag} */,
  {32'hc18532ec, 32'hc0db92b8} /* (4, 8, 7) {real, imag} */,
  {32'hc2e6fbe3, 32'h421e4dcf} /* (4, 8, 6) {real, imag} */,
  {32'h4203ee9c, 32'h41bbc790} /* (4, 8, 5) {real, imag} */,
  {32'hc2eb928c, 32'hc2a080a2} /* (4, 8, 4) {real, imag} */,
  {32'h4376310f, 32'h4291eded} /* (4, 8, 3) {real, imag} */,
  {32'h43338e0a, 32'h43599bd8} /* (4, 8, 2) {real, imag} */,
  {32'h42bc10ed, 32'hc298ade1} /* (4, 8, 1) {real, imag} */,
  {32'hc313a7f2, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'hc2aae5e0, 32'hc0df0b88} /* (4, 7, 15) {real, imag} */,
  {32'h432b03f0, 32'hc2e9b7da} /* (4, 7, 14) {real, imag} */,
  {32'hc2538a9a, 32'hc2ff8ce2} /* (4, 7, 13) {real, imag} */,
  {32'hc212bfa3, 32'h428486de} /* (4, 7, 12) {real, imag} */,
  {32'hc0aefa94, 32'hc301674c} /* (4, 7, 11) {real, imag} */,
  {32'hc1e34d28, 32'h407390a0} /* (4, 7, 10) {real, imag} */,
  {32'h433aea88, 32'h42202010} /* (4, 7, 9) {real, imag} */,
  {32'hc2264a1a, 32'h00000000} /* (4, 7, 8) {real, imag} */,
  {32'h433aea88, 32'hc2202010} /* (4, 7, 7) {real, imag} */,
  {32'hc1e34d28, 32'hc07390a0} /* (4, 7, 6) {real, imag} */,
  {32'hc0aefa94, 32'h4301674c} /* (4, 7, 5) {real, imag} */,
  {32'hc212bfa3, 32'hc28486de} /* (4, 7, 4) {real, imag} */,
  {32'hc2538a9a, 32'h42ff8ce2} /* (4, 7, 3) {real, imag} */,
  {32'h432b03f0, 32'h42e9b7da} /* (4, 7, 2) {real, imag} */,
  {32'hc2aae5e0, 32'h40df0b88} /* (4, 7, 1) {real, imag} */,
  {32'hc3860da0, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'hc37edc95, 32'h42f09708} /* (4, 6, 15) {real, imag} */,
  {32'h4362e434, 32'hc311ad88} /* (4, 6, 14) {real, imag} */,
  {32'hc0fd22d8, 32'hc316bdb2} /* (4, 6, 13) {real, imag} */,
  {32'hc1a48296, 32'hc2187d89} /* (4, 6, 12) {real, imag} */,
  {32'h428551e9, 32'hc25ff056} /* (4, 6, 11) {real, imag} */,
  {32'hc211adca, 32'h42c215d9} /* (4, 6, 10) {real, imag} */,
  {32'hbf2792c0, 32'hc308616a} /* (4, 6, 9) {real, imag} */,
  {32'h4068a6b0, 32'h00000000} /* (4, 6, 8) {real, imag} */,
  {32'hbf2792c0, 32'h4308616a} /* (4, 6, 7) {real, imag} */,
  {32'hc211adca, 32'hc2c215d9} /* (4, 6, 6) {real, imag} */,
  {32'h428551e9, 32'h425ff056} /* (4, 6, 5) {real, imag} */,
  {32'hc1a48296, 32'h42187d89} /* (4, 6, 4) {real, imag} */,
  {32'hc0fd22d8, 32'h4316bdb2} /* (4, 6, 3) {real, imag} */,
  {32'h4362e434, 32'h4311ad88} /* (4, 6, 2) {real, imag} */,
  {32'hc37edc95, 32'hc2f09708} /* (4, 6, 1) {real, imag} */,
  {32'hc41a2b8f, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'hc399dba6, 32'h42c9fb29} /* (4, 5, 15) {real, imag} */,
  {32'h42548b15, 32'hc2a35d93} /* (4, 5, 14) {real, imag} */,
  {32'h42b06238, 32'h42511418} /* (4, 5, 13) {real, imag} */,
  {32'hc1821f4a, 32'hc2386d80} /* (4, 5, 12) {real, imag} */,
  {32'hbf6b2f80, 32'hc2378016} /* (4, 5, 11) {real, imag} */,
  {32'hc1f5959e, 32'h42f972dc} /* (4, 5, 10) {real, imag} */,
  {32'hc2fa3838, 32'h41d336ae} /* (4, 5, 9) {real, imag} */,
  {32'h4181a8aa, 32'h00000000} /* (4, 5, 8) {real, imag} */,
  {32'hc2fa3838, 32'hc1d336ae} /* (4, 5, 7) {real, imag} */,
  {32'hc1f5959e, 32'hc2f972dc} /* (4, 5, 6) {real, imag} */,
  {32'hbf6b2f80, 32'h42378016} /* (4, 5, 5) {real, imag} */,
  {32'hc1821f4a, 32'h42386d80} /* (4, 5, 4) {real, imag} */,
  {32'h42b06238, 32'hc2511418} /* (4, 5, 3) {real, imag} */,
  {32'h42548b15, 32'h42a35d93} /* (4, 5, 2) {real, imag} */,
  {32'hc399dba6, 32'hc2c9fb29} /* (4, 5, 1) {real, imag} */,
  {32'hc37fa3e6, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'hc3431ee8, 32'hc344651c} /* (4, 4, 15) {real, imag} */,
  {32'hc2717fd8, 32'h42d68c9d} /* (4, 4, 14) {real, imag} */,
  {32'h435670f4, 32'hc205f65c} /* (4, 4, 13) {real, imag} */,
  {32'h4125f1ea, 32'h42bd6392} /* (4, 4, 12) {real, imag} */,
  {32'hc0c3bda4, 32'hc2c35b4e} /* (4, 4, 11) {real, imag} */,
  {32'h42334b86, 32'h424de7b1} /* (4, 4, 10) {real, imag} */,
  {32'h4232b387, 32'hc0225450} /* (4, 4, 9) {real, imag} */,
  {32'h417f1434, 32'h00000000} /* (4, 4, 8) {real, imag} */,
  {32'h4232b387, 32'h40225450} /* (4, 4, 7) {real, imag} */,
  {32'h42334b86, 32'hc24de7b1} /* (4, 4, 6) {real, imag} */,
  {32'hc0c3bda4, 32'h42c35b4e} /* (4, 4, 5) {real, imag} */,
  {32'h4125f1ea, 32'hc2bd6392} /* (4, 4, 4) {real, imag} */,
  {32'h435670f4, 32'h4205f65c} /* (4, 4, 3) {real, imag} */,
  {32'hc2717fd8, 32'hc2d68c9d} /* (4, 4, 2) {real, imag} */,
  {32'hc3431ee8, 32'h4344651c} /* (4, 4, 1) {real, imag} */,
  {32'hc3df725c, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'hc38bbb12, 32'hc395be88} /* (4, 3, 15) {real, imag} */,
  {32'h42058d9e, 32'hc03c6ba0} /* (4, 3, 14) {real, imag} */,
  {32'h42c4b462, 32'h420a14bc} /* (4, 3, 13) {real, imag} */,
  {32'h42a46db0, 32'hc294e4d2} /* (4, 3, 12) {real, imag} */,
  {32'h4291dadd, 32'hc302c696} /* (4, 3, 11) {real, imag} */,
  {32'hc03e4ae0, 32'h428aad8e} /* (4, 3, 10) {real, imag} */,
  {32'h4344f5b0, 32'hc1eb2dcc} /* (4, 3, 9) {real, imag} */,
  {32'h42602efe, 32'h00000000} /* (4, 3, 8) {real, imag} */,
  {32'h4344f5b0, 32'h41eb2dcc} /* (4, 3, 7) {real, imag} */,
  {32'hc03e4ae0, 32'hc28aad8e} /* (4, 3, 6) {real, imag} */,
  {32'h4291dadd, 32'h4302c696} /* (4, 3, 5) {real, imag} */,
  {32'h42a46db0, 32'h4294e4d2} /* (4, 3, 4) {real, imag} */,
  {32'h42c4b462, 32'hc20a14bc} /* (4, 3, 3) {real, imag} */,
  {32'h42058d9e, 32'h403c6ba0} /* (4, 3, 2) {real, imag} */,
  {32'hc38bbb12, 32'h4395be88} /* (4, 3, 1) {real, imag} */,
  {32'hc417ef34, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'hc32f6aca, 32'hc38910b9} /* (4, 2, 15) {real, imag} */,
  {32'hc24d01e7, 32'hc213f1dd} /* (4, 2, 14) {real, imag} */,
  {32'h423fea71, 32'h43575f80} /* (4, 2, 13) {real, imag} */,
  {32'h42f2f780, 32'h4230708a} /* (4, 2, 12) {real, imag} */,
  {32'hc0687448, 32'hc1d94073} /* (4, 2, 11) {real, imag} */,
  {32'hc1e8e47f, 32'hc16a3413} /* (4, 2, 10) {real, imag} */,
  {32'h4110dde0, 32'h428d0b64} /* (4, 2, 9) {real, imag} */,
  {32'h4198cc32, 32'h00000000} /* (4, 2, 8) {real, imag} */,
  {32'h4110dde0, 32'hc28d0b64} /* (4, 2, 7) {real, imag} */,
  {32'hc1e8e47f, 32'h416a3413} /* (4, 2, 6) {real, imag} */,
  {32'hc0687448, 32'h41d94073} /* (4, 2, 5) {real, imag} */,
  {32'h42f2f780, 32'hc230708a} /* (4, 2, 4) {real, imag} */,
  {32'h423fea71, 32'hc3575f80} /* (4, 2, 3) {real, imag} */,
  {32'hc24d01e7, 32'h4213f1dd} /* (4, 2, 2) {real, imag} */,
  {32'hc32f6aca, 32'h438910b9} /* (4, 2, 1) {real, imag} */,
  {32'hc40f2b57, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'hc337d8f2, 32'hc30d2424} /* (4, 1, 15) {real, imag} */,
  {32'hc2be0f55, 32'hc2f0636b} /* (4, 1, 14) {real, imag} */,
  {32'hc18e6839, 32'hc22f93a1} /* (4, 1, 13) {real, imag} */,
  {32'h3fdf6de0, 32'h42be34b7} /* (4, 1, 12) {real, imag} */,
  {32'h422ee3cc, 32'hc0ba48b8} /* (4, 1, 11) {real, imag} */,
  {32'h42bc1e04, 32'hc2b303cf} /* (4, 1, 10) {real, imag} */,
  {32'hc0089f30, 32'h4254e1c8} /* (4, 1, 9) {real, imag} */,
  {32'hc21a51da, 32'h00000000} /* (4, 1, 8) {real, imag} */,
  {32'hc0089f30, 32'hc254e1c8} /* (4, 1, 7) {real, imag} */,
  {32'h42bc1e04, 32'h42b303cf} /* (4, 1, 6) {real, imag} */,
  {32'h422ee3cc, 32'h40ba48b8} /* (4, 1, 5) {real, imag} */,
  {32'h3fdf6de0, 32'hc2be34b7} /* (4, 1, 4) {real, imag} */,
  {32'hc18e6839, 32'h422f93a1} /* (4, 1, 3) {real, imag} */,
  {32'hc2be0f55, 32'h42f0636b} /* (4, 1, 2) {real, imag} */,
  {32'hc337d8f2, 32'h430d2424} /* (4, 1, 1) {real, imag} */,
  {32'hc3ac4f1d, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'hc33d0f06, 32'h42c51d1b} /* (4, 0, 15) {real, imag} */,
  {32'h41d15af8, 32'hc311ab22} /* (4, 0, 14) {real, imag} */,
  {32'hc222e33c, 32'hc2d08dd3} /* (4, 0, 13) {real, imag} */,
  {32'h4000fdd0, 32'h428c4584} /* (4, 0, 12) {real, imag} */,
  {32'h420abf68, 32'h41b99550} /* (4, 0, 11) {real, imag} */,
  {32'h42879511, 32'hc0e59738} /* (4, 0, 10) {real, imag} */,
  {32'hc205d0c6, 32'h41be3e1a} /* (4, 0, 9) {real, imag} */,
  {32'h420516d0, 32'h00000000} /* (4, 0, 8) {real, imag} */,
  {32'hc205d0c6, 32'hc1be3e1a} /* (4, 0, 7) {real, imag} */,
  {32'h42879511, 32'h40e59738} /* (4, 0, 6) {real, imag} */,
  {32'h420abf68, 32'hc1b99550} /* (4, 0, 5) {real, imag} */,
  {32'h4000fdd0, 32'hc28c4584} /* (4, 0, 4) {real, imag} */,
  {32'hc222e33c, 32'h42d08dd3} /* (4, 0, 3) {real, imag} */,
  {32'h41d15af8, 32'h4311ab22} /* (4, 0, 2) {real, imag} */,
  {32'hc33d0f06, 32'hc2c51d1b} /* (4, 0, 1) {real, imag} */,
  {32'hc3b22139, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hc351df59, 32'hc2079864} /* (3, 15, 15) {real, imag} */,
  {32'h4112a0d8, 32'h419ff050} /* (3, 15, 14) {real, imag} */,
  {32'h4192524a, 32'h42c4b8fc} /* (3, 15, 13) {real, imag} */,
  {32'hc2625086, 32'hc258a847} /* (3, 15, 12) {real, imag} */,
  {32'hc20672c2, 32'hc2bdfe16} /* (3, 15, 11) {real, imag} */,
  {32'h4292578d, 32'hc27e769f} /* (3, 15, 10) {real, imag} */,
  {32'h408508ba, 32'h420d9326} /* (3, 15, 9) {real, imag} */,
  {32'hc2e6f2b6, 32'h00000000} /* (3, 15, 8) {real, imag} */,
  {32'h408508ba, 32'hc20d9326} /* (3, 15, 7) {real, imag} */,
  {32'h4292578d, 32'h427e769f} /* (3, 15, 6) {real, imag} */,
  {32'hc20672c2, 32'h42bdfe16} /* (3, 15, 5) {real, imag} */,
  {32'hc2625086, 32'h4258a847} /* (3, 15, 4) {real, imag} */,
  {32'h4192524a, 32'hc2c4b8fc} /* (3, 15, 3) {real, imag} */,
  {32'h4112a0d8, 32'hc19ff050} /* (3, 15, 2) {real, imag} */,
  {32'hc351df59, 32'h42079864} /* (3, 15, 1) {real, imag} */,
  {32'hc361a5c5, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'hc2feabf5, 32'h4191feb8} /* (3, 14, 15) {real, imag} */,
  {32'hc261c09e, 32'h40877108} /* (3, 14, 14) {real, imag} */,
  {32'h42bb0770, 32'h40e3a608} /* (3, 14, 13) {real, imag} */,
  {32'h435fdeb8, 32'hc30f1ba2} /* (3, 14, 12) {real, imag} */,
  {32'hc34bafd4, 32'hc1b7ed64} /* (3, 14, 11) {real, imag} */,
  {32'h42dc9d9f, 32'hc261b791} /* (3, 14, 10) {real, imag} */,
  {32'h419496a7, 32'hc2191c95} /* (3, 14, 9) {real, imag} */,
  {32'h42a65fa2, 32'h00000000} /* (3, 14, 8) {real, imag} */,
  {32'h419496a7, 32'h42191c95} /* (3, 14, 7) {real, imag} */,
  {32'h42dc9d9f, 32'h4261b791} /* (3, 14, 6) {real, imag} */,
  {32'hc34bafd4, 32'h41b7ed64} /* (3, 14, 5) {real, imag} */,
  {32'h435fdeb8, 32'h430f1ba2} /* (3, 14, 4) {real, imag} */,
  {32'h42bb0770, 32'hc0e3a608} /* (3, 14, 3) {real, imag} */,
  {32'hc261c09e, 32'hc0877108} /* (3, 14, 2) {real, imag} */,
  {32'hc2feabf5, 32'hc191feb8} /* (3, 14, 1) {real, imag} */,
  {32'hc32764f4, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'h409f7550, 32'h430942ae} /* (3, 13, 15) {real, imag} */,
  {32'hc2b5b701, 32'h416dac28} /* (3, 13, 14) {real, imag} */,
  {32'h4262c0a4, 32'h42e87990} /* (3, 13, 13) {real, imag} */,
  {32'h431da954, 32'hc15371c2} /* (3, 13, 12) {real, imag} */,
  {32'h4080d420, 32'hc2d5373c} /* (3, 13, 11) {real, imag} */,
  {32'h42320be9, 32'h422c8787} /* (3, 13, 10) {real, imag} */,
  {32'hc2a35057, 32'h427a782a} /* (3, 13, 9) {real, imag} */,
  {32'hc1ac2f10, 32'h00000000} /* (3, 13, 8) {real, imag} */,
  {32'hc2a35057, 32'hc27a782a} /* (3, 13, 7) {real, imag} */,
  {32'h42320be9, 32'hc22c8787} /* (3, 13, 6) {real, imag} */,
  {32'h4080d420, 32'h42d5373c} /* (3, 13, 5) {real, imag} */,
  {32'h431da954, 32'h415371c2} /* (3, 13, 4) {real, imag} */,
  {32'h4262c0a4, 32'hc2e87990} /* (3, 13, 3) {real, imag} */,
  {32'hc2b5b701, 32'hc16dac28} /* (3, 13, 2) {real, imag} */,
  {32'h409f7550, 32'hc30942ae} /* (3, 13, 1) {real, imag} */,
  {32'h400e3700, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'h409adc70, 32'h42400e1a} /* (3, 12, 15) {real, imag} */,
  {32'hc301abc0, 32'hc363f352} /* (3, 12, 14) {real, imag} */,
  {32'h4250499f, 32'h43274e3e} /* (3, 12, 13) {real, imag} */,
  {32'hc0ead808, 32'h42c95410} /* (3, 12, 12) {real, imag} */,
  {32'h427049ba, 32'hc2f66464} /* (3, 12, 11) {real, imag} */,
  {32'hc0bc77d0, 32'hc2a7bf56} /* (3, 12, 10) {real, imag} */,
  {32'hc1cc0e02, 32'h4236e564} /* (3, 12, 9) {real, imag} */,
  {32'h404916b0, 32'h00000000} /* (3, 12, 8) {real, imag} */,
  {32'hc1cc0e02, 32'hc236e564} /* (3, 12, 7) {real, imag} */,
  {32'hc0bc77d0, 32'h42a7bf56} /* (3, 12, 6) {real, imag} */,
  {32'h427049ba, 32'h42f66464} /* (3, 12, 5) {real, imag} */,
  {32'hc0ead808, 32'hc2c95410} /* (3, 12, 4) {real, imag} */,
  {32'h4250499f, 32'hc3274e3e} /* (3, 12, 3) {real, imag} */,
  {32'hc301abc0, 32'h4363f352} /* (3, 12, 2) {real, imag} */,
  {32'h409adc70, 32'hc2400e1a} /* (3, 12, 1) {real, imag} */,
  {32'h415a0ea0, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'hc14f5578, 32'h4288089f} /* (3, 11, 15) {real, imag} */,
  {32'hc32892ae, 32'hc0e3fe74} /* (3, 11, 14) {real, imag} */,
  {32'h4208e560, 32'hc2e7071e} /* (3, 11, 13) {real, imag} */,
  {32'h431f1c20, 32'h420eac60} /* (3, 11, 12) {real, imag} */,
  {32'hc225f2f8, 32'hc1261b7c} /* (3, 11, 11) {real, imag} */,
  {32'h432eb906, 32'h416e346c} /* (3, 11, 10) {real, imag} */,
  {32'hc0f65c0c, 32'hc2d98d46} /* (3, 11, 9) {real, imag} */,
  {32'hc0804940, 32'h00000000} /* (3, 11, 8) {real, imag} */,
  {32'hc0f65c0c, 32'h42d98d46} /* (3, 11, 7) {real, imag} */,
  {32'h432eb906, 32'hc16e346c} /* (3, 11, 6) {real, imag} */,
  {32'hc225f2f8, 32'h41261b7c} /* (3, 11, 5) {real, imag} */,
  {32'h431f1c20, 32'hc20eac60} /* (3, 11, 4) {real, imag} */,
  {32'h4208e560, 32'h42e7071e} /* (3, 11, 3) {real, imag} */,
  {32'hc32892ae, 32'h40e3fe74} /* (3, 11, 2) {real, imag} */,
  {32'hc14f5578, 32'hc288089f} /* (3, 11, 1) {real, imag} */,
  {32'h42ec555e, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'h41c4031e, 32'h41606388} /* (3, 10, 15) {real, imag} */,
  {32'hc2803bed, 32'h431893c1} /* (3, 10, 14) {real, imag} */,
  {32'h4313df2e, 32'hc27a8b15} /* (3, 10, 13) {real, imag} */,
  {32'h43180d3c, 32'hc25ba2c5} /* (3, 10, 12) {real, imag} */,
  {32'h426b15e1, 32'hc1296b60} /* (3, 10, 11) {real, imag} */,
  {32'hc322f380, 32'hc29cc121} /* (3, 10, 10) {real, imag} */,
  {32'h40a6c5a8, 32'hc0a2e010} /* (3, 10, 9) {real, imag} */,
  {32'hc25f2df2, 32'h00000000} /* (3, 10, 8) {real, imag} */,
  {32'h40a6c5a8, 32'h40a2e010} /* (3, 10, 7) {real, imag} */,
  {32'hc322f380, 32'h429cc121} /* (3, 10, 6) {real, imag} */,
  {32'h426b15e1, 32'h41296b60} /* (3, 10, 5) {real, imag} */,
  {32'h43180d3c, 32'h425ba2c5} /* (3, 10, 4) {real, imag} */,
  {32'h4313df2e, 32'h427a8b15} /* (3, 10, 3) {real, imag} */,
  {32'hc2803bed, 32'hc31893c1} /* (3, 10, 2) {real, imag} */,
  {32'h41c4031e, 32'hc1606388} /* (3, 10, 1) {real, imag} */,
  {32'hc1271420, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'h429937fc, 32'h421db0e4} /* (3, 9, 15) {real, imag} */,
  {32'h42a651cd, 32'hc3046afd} /* (3, 9, 14) {real, imag} */,
  {32'h428ce6a2, 32'hc2839c4e} /* (3, 9, 13) {real, imag} */,
  {32'h42272adf, 32'hc1862aba} /* (3, 9, 12) {real, imag} */,
  {32'h423a92c0, 32'h4290087b} /* (3, 9, 11) {real, imag} */,
  {32'hc2f3ba39, 32'h426dd67c} /* (3, 9, 10) {real, imag} */,
  {32'hc180c090, 32'h41345ae2} /* (3, 9, 9) {real, imag} */,
  {32'h40fa440c, 32'h00000000} /* (3, 9, 8) {real, imag} */,
  {32'hc180c090, 32'hc1345ae2} /* (3, 9, 7) {real, imag} */,
  {32'hc2f3ba39, 32'hc26dd67c} /* (3, 9, 6) {real, imag} */,
  {32'h423a92c0, 32'hc290087b} /* (3, 9, 5) {real, imag} */,
  {32'h42272adf, 32'h41862aba} /* (3, 9, 4) {real, imag} */,
  {32'h428ce6a2, 32'h42839c4e} /* (3, 9, 3) {real, imag} */,
  {32'h42a651cd, 32'h43046afd} /* (3, 9, 2) {real, imag} */,
  {32'h429937fc, 32'hc21db0e4} /* (3, 9, 1) {real, imag} */,
  {32'h41324f50, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'hc30ac46b, 32'hc229dfd4} /* (3, 8, 15) {real, imag} */,
  {32'h42a1ff6c, 32'hc3956756} /* (3, 8, 14) {real, imag} */,
  {32'h42da236a, 32'hc3064102} /* (3, 8, 13) {real, imag} */,
  {32'h410804a4, 32'h42487ed6} /* (3, 8, 12) {real, imag} */,
  {32'h412fa3c2, 32'hc20edb5c} /* (3, 8, 11) {real, imag} */,
  {32'h42a02451, 32'h4347c5cd} /* (3, 8, 10) {real, imag} */,
  {32'hc2ae986e, 32'hc18119e0} /* (3, 8, 9) {real, imag} */,
  {32'h423bc6fe, 32'h00000000} /* (3, 8, 8) {real, imag} */,
  {32'hc2ae986e, 32'h418119e0} /* (3, 8, 7) {real, imag} */,
  {32'h42a02451, 32'hc347c5cd} /* (3, 8, 6) {real, imag} */,
  {32'h412fa3c2, 32'h420edb5c} /* (3, 8, 5) {real, imag} */,
  {32'h410804a4, 32'hc2487ed6} /* (3, 8, 4) {real, imag} */,
  {32'h42da236a, 32'h43064102} /* (3, 8, 3) {real, imag} */,
  {32'h42a1ff6c, 32'h43956756} /* (3, 8, 2) {real, imag} */,
  {32'hc30ac46b, 32'h4229dfd4} /* (3, 8, 1) {real, imag} */,
  {32'h4198c1e0, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'hc310b0b6, 32'hc332afc9} /* (3, 7, 15) {real, imag} */,
  {32'h4306b152, 32'hc248f7f7} /* (3, 7, 14) {real, imag} */,
  {32'hc2807d36, 32'hc33e0259} /* (3, 7, 13) {real, imag} */,
  {32'hc27fb9f5, 32'h4292fb24} /* (3, 7, 12) {real, imag} */,
  {32'h429ec169, 32'hc2819ec5} /* (3, 7, 11) {real, imag} */,
  {32'hc07a60a0, 32'hc0826850} /* (3, 7, 10) {real, imag} */,
  {32'hc1f1f024, 32'hc1d5ba8f} /* (3, 7, 9) {real, imag} */,
  {32'hc20380b6, 32'h00000000} /* (3, 7, 8) {real, imag} */,
  {32'hc1f1f024, 32'h41d5ba8f} /* (3, 7, 7) {real, imag} */,
  {32'hc07a60a0, 32'h40826850} /* (3, 7, 6) {real, imag} */,
  {32'h429ec169, 32'h42819ec5} /* (3, 7, 5) {real, imag} */,
  {32'hc27fb9f5, 32'hc292fb24} /* (3, 7, 4) {real, imag} */,
  {32'hc2807d36, 32'h433e0259} /* (3, 7, 3) {real, imag} */,
  {32'h4306b152, 32'h4248f7f7} /* (3, 7, 2) {real, imag} */,
  {32'hc310b0b6, 32'h4332afc9} /* (3, 7, 1) {real, imag} */,
  {32'hc3a605f8, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'hc3055c79, 32'hc291dbc0} /* (3, 6, 15) {real, imag} */,
  {32'h42a7bdeb, 32'h41116d30} /* (3, 6, 14) {real, imag} */,
  {32'h43035a02, 32'h41ea2a92} /* (3, 6, 13) {real, imag} */,
  {32'h41869a64, 32'hc290d71a} /* (3, 6, 12) {real, imag} */,
  {32'h42b65b10, 32'hc2c7b0ff} /* (3, 6, 11) {real, imag} */,
  {32'hc1d73ba4, 32'hbf387280} /* (3, 6, 10) {real, imag} */,
  {32'hc30175a0, 32'h42c6848e} /* (3, 6, 9) {real, imag} */,
  {32'hc2f832bb, 32'h00000000} /* (3, 6, 8) {real, imag} */,
  {32'hc30175a0, 32'hc2c6848e} /* (3, 6, 7) {real, imag} */,
  {32'hc1d73ba4, 32'h3f387280} /* (3, 6, 6) {real, imag} */,
  {32'h42b65b10, 32'h42c7b0ff} /* (3, 6, 5) {real, imag} */,
  {32'h41869a64, 32'h4290d71a} /* (3, 6, 4) {real, imag} */,
  {32'h43035a02, 32'hc1ea2a92} /* (3, 6, 3) {real, imag} */,
  {32'h42a7bdeb, 32'hc1116d30} /* (3, 6, 2) {real, imag} */,
  {32'hc3055c79, 32'h4291dbc0} /* (3, 6, 1) {real, imag} */,
  {32'hc404f434, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hc33d7322, 32'hc27cd2e1} /* (3, 5, 15) {real, imag} */,
  {32'h4356502a, 32'hc0ed446c} /* (3, 5, 14) {real, imag} */,
  {32'h42476260, 32'h4255087b} /* (3, 5, 13) {real, imag} */,
  {32'h4183f9d8, 32'h428d7507} /* (3, 5, 12) {real, imag} */,
  {32'h43358c36, 32'h4223e01f} /* (3, 5, 11) {real, imag} */,
  {32'hc2fc9d0d, 32'h42c72eac} /* (3, 5, 10) {real, imag} */,
  {32'hc0a8d764, 32'hc14d4350} /* (3, 5, 9) {real, imag} */,
  {32'hc1bccf88, 32'h00000000} /* (3, 5, 8) {real, imag} */,
  {32'hc0a8d764, 32'h414d4350} /* (3, 5, 7) {real, imag} */,
  {32'hc2fc9d0d, 32'hc2c72eac} /* (3, 5, 6) {real, imag} */,
  {32'h43358c36, 32'hc223e01f} /* (3, 5, 5) {real, imag} */,
  {32'h4183f9d8, 32'hc28d7507} /* (3, 5, 4) {real, imag} */,
  {32'h42476260, 32'hc255087b} /* (3, 5, 3) {real, imag} */,
  {32'h4356502a, 32'h40ed446c} /* (3, 5, 2) {real, imag} */,
  {32'hc33d7322, 32'h427cd2e1} /* (3, 5, 1) {real, imag} */,
  {32'hc3cd80a4, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hc35201ac, 32'hc35eee58} /* (3, 4, 15) {real, imag} */,
  {32'hc2112a6e, 32'h42ba0bcc} /* (3, 4, 14) {real, imag} */,
  {32'h421078af, 32'hc0c901d0} /* (3, 4, 13) {real, imag} */,
  {32'h42b25dee, 32'hc28d2302} /* (3, 4, 12) {real, imag} */,
  {32'hc225dbf2, 32'h42c62258} /* (3, 4, 11) {real, imag} */,
  {32'h43207022, 32'hc300e27d} /* (3, 4, 10) {real, imag} */,
  {32'hc228f99f, 32'h42b07780} /* (3, 4, 9) {real, imag} */,
  {32'h42b998bc, 32'h00000000} /* (3, 4, 8) {real, imag} */,
  {32'hc228f99f, 32'hc2b07780} /* (3, 4, 7) {real, imag} */,
  {32'h43207022, 32'h4300e27d} /* (3, 4, 6) {real, imag} */,
  {32'hc225dbf2, 32'hc2c62258} /* (3, 4, 5) {real, imag} */,
  {32'h42b25dee, 32'h428d2302} /* (3, 4, 4) {real, imag} */,
  {32'h421078af, 32'h40c901d0} /* (3, 4, 3) {real, imag} */,
  {32'hc2112a6e, 32'hc2ba0bcc} /* (3, 4, 2) {real, imag} */,
  {32'hc35201ac, 32'h435eee58} /* (3, 4, 1) {real, imag} */,
  {32'hc41700de, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hc3024d88, 32'hc2c66718} /* (3, 3, 15) {real, imag} */,
  {32'h41d476a4, 32'h43003c96} /* (3, 3, 14) {real, imag} */,
  {32'h428a9126, 32'h42a27758} /* (3, 3, 13) {real, imag} */,
  {32'h42c3f989, 32'hc20be44e} /* (3, 3, 12) {real, imag} */,
  {32'hc343a1ab, 32'hc0b278f8} /* (3, 3, 11) {real, imag} */,
  {32'hc224006b, 32'hc081c618} /* (3, 3, 10) {real, imag} */,
  {32'h4155cf48, 32'h41287508} /* (3, 3, 9) {real, imag} */,
  {32'hc30c8ba9, 32'h00000000} /* (3, 3, 8) {real, imag} */,
  {32'h4155cf48, 32'hc1287508} /* (3, 3, 7) {real, imag} */,
  {32'hc224006b, 32'h4081c618} /* (3, 3, 6) {real, imag} */,
  {32'hc343a1ab, 32'h40b278f8} /* (3, 3, 5) {real, imag} */,
  {32'h42c3f989, 32'h420be44e} /* (3, 3, 4) {real, imag} */,
  {32'h428a9126, 32'hc2a27758} /* (3, 3, 3) {real, imag} */,
  {32'h41d476a4, 32'hc3003c96} /* (3, 3, 2) {real, imag} */,
  {32'hc3024d88, 32'h42c66718} /* (3, 3, 1) {real, imag} */,
  {32'hc40c0c6b, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hc356b89c, 32'hc38f4782} /* (3, 2, 15) {real, imag} */,
  {32'h42194e58, 32'hc0044670} /* (3, 2, 14) {real, imag} */,
  {32'h4290a980, 32'h42e8f148} /* (3, 2, 13) {real, imag} */,
  {32'hc216a2c2, 32'h4253949b} /* (3, 2, 12) {real, imag} */,
  {32'h4299cde8, 32'hc22839c0} /* (3, 2, 11) {real, imag} */,
  {32'h421809b6, 32'h41488a7c} /* (3, 2, 10) {real, imag} */,
  {32'h42013cfa, 32'hc2187671} /* (3, 2, 9) {real, imag} */,
  {32'h42635d75, 32'h00000000} /* (3, 2, 8) {real, imag} */,
  {32'h42013cfa, 32'h42187671} /* (3, 2, 7) {real, imag} */,
  {32'h421809b6, 32'hc1488a7c} /* (3, 2, 6) {real, imag} */,
  {32'h4299cde8, 32'h422839c0} /* (3, 2, 5) {real, imag} */,
  {32'hc216a2c2, 32'hc253949b} /* (3, 2, 4) {real, imag} */,
  {32'h4290a980, 32'hc2e8f148} /* (3, 2, 3) {real, imag} */,
  {32'h42194e58, 32'h40044670} /* (3, 2, 2) {real, imag} */,
  {32'hc356b89c, 32'h438f4782} /* (3, 2, 1) {real, imag} */,
  {32'hc40f99c2, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hc2675cf4, 32'hc3257d43} /* (3, 1, 15) {real, imag} */,
  {32'hc3233c72, 32'h411fe3d0} /* (3, 1, 14) {real, imag} */,
  {32'hc26c2101, 32'h435e94e2} /* (3, 1, 13) {real, imag} */,
  {32'hc228e994, 32'hc25beac9} /* (3, 1, 12) {real, imag} */,
  {32'h4184abf8, 32'hc33f202d} /* (3, 1, 11) {real, imag} */,
  {32'h432a08fa, 32'hc2a562e1} /* (3, 1, 10) {real, imag} */,
  {32'hbfedf058, 32'hc1eccf78} /* (3, 1, 9) {real, imag} */,
  {32'h428c7b22, 32'h00000000} /* (3, 1, 8) {real, imag} */,
  {32'hbfedf058, 32'h41eccf78} /* (3, 1, 7) {real, imag} */,
  {32'h432a08fa, 32'h42a562e1} /* (3, 1, 6) {real, imag} */,
  {32'h4184abf8, 32'h433f202d} /* (3, 1, 5) {real, imag} */,
  {32'hc228e994, 32'h425beac9} /* (3, 1, 4) {real, imag} */,
  {32'hc26c2101, 32'hc35e94e2} /* (3, 1, 3) {real, imag} */,
  {32'hc3233c72, 32'hc11fe3d0} /* (3, 1, 2) {real, imag} */,
  {32'hc2675cf4, 32'h43257d43} /* (3, 1, 1) {real, imag} */,
  {32'hc39eb116, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'h4216a7ad, 32'hc2c74b2c} /* (3, 0, 15) {real, imag} */,
  {32'hc35017b2, 32'hc18bb638} /* (3, 0, 14) {real, imag} */,
  {32'hc2037df1, 32'h424105af} /* (3, 0, 13) {real, imag} */,
  {32'h4292d19c, 32'h4380a953} /* (3, 0, 12) {real, imag} */,
  {32'hc19ff3ff, 32'h42ffda94} /* (3, 0, 11) {real, imag} */,
  {32'h4187ef04, 32'hc208a8ac} /* (3, 0, 10) {real, imag} */,
  {32'hc23e5be0, 32'hc29fced1} /* (3, 0, 9) {real, imag} */,
  {32'h42cc9ab5, 32'h00000000} /* (3, 0, 8) {real, imag} */,
  {32'hc23e5be0, 32'h429fced1} /* (3, 0, 7) {real, imag} */,
  {32'h4187ef04, 32'h4208a8ac} /* (3, 0, 6) {real, imag} */,
  {32'hc19ff3ff, 32'hc2ffda94} /* (3, 0, 5) {real, imag} */,
  {32'h4292d19c, 32'hc380a953} /* (3, 0, 4) {real, imag} */,
  {32'hc2037df1, 32'hc24105af} /* (3, 0, 3) {real, imag} */,
  {32'hc35017b2, 32'h418bb638} /* (3, 0, 2) {real, imag} */,
  {32'h4216a7ad, 32'h42c74b2c} /* (3, 0, 1) {real, imag} */,
  {32'hc2e38ad4, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hc37c473c, 32'hc3273bc6} /* (2, 15, 15) {real, imag} */,
  {32'h4270bb36, 32'hc25b4462} /* (2, 15, 14) {real, imag} */,
  {32'hbf2ef180, 32'h4258433a} /* (2, 15, 13) {real, imag} */,
  {32'hc15f2940, 32'h40791cd0} /* (2, 15, 12) {real, imag} */,
  {32'hc18d6ff4, 32'h4304013c} /* (2, 15, 11) {real, imag} */,
  {32'hc2a72bd3, 32'hc1c84e96} /* (2, 15, 10) {real, imag} */,
  {32'h4151e1a8, 32'hc2359a7e} /* (2, 15, 9) {real, imag} */,
  {32'hc22b2674, 32'h00000000} /* (2, 15, 8) {real, imag} */,
  {32'h4151e1a8, 32'h42359a7e} /* (2, 15, 7) {real, imag} */,
  {32'hc2a72bd3, 32'h41c84e96} /* (2, 15, 6) {real, imag} */,
  {32'hc18d6ff4, 32'hc304013c} /* (2, 15, 5) {real, imag} */,
  {32'hc15f2940, 32'hc0791cd0} /* (2, 15, 4) {real, imag} */,
  {32'hbf2ef180, 32'hc258433a} /* (2, 15, 3) {real, imag} */,
  {32'h4270bb36, 32'h425b4462} /* (2, 15, 2) {real, imag} */,
  {32'hc37c473c, 32'h43273bc6} /* (2, 15, 1) {real, imag} */,
  {32'hc3637edd, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'hc28c0576, 32'hc25a928e} /* (2, 14, 15) {real, imag} */,
  {32'h42d4735a, 32'hc2ed3686} /* (2, 14, 14) {real, imag} */,
  {32'h40fb9bd8, 32'hc1dace70} /* (2, 14, 13) {real, imag} */,
  {32'h3f89ec30, 32'hc2b3821c} /* (2, 14, 12) {real, imag} */,
  {32'hc2188465, 32'hbdb66400} /* (2, 14, 11) {real, imag} */,
  {32'h4264bbde, 32'hc13e206c} /* (2, 14, 10) {real, imag} */,
  {32'hc0cc290c, 32'h42c33a2c} /* (2, 14, 9) {real, imag} */,
  {32'h422c13a8, 32'h00000000} /* (2, 14, 8) {real, imag} */,
  {32'hc0cc290c, 32'hc2c33a2c} /* (2, 14, 7) {real, imag} */,
  {32'h4264bbde, 32'h413e206c} /* (2, 14, 6) {real, imag} */,
  {32'hc2188465, 32'h3db66400} /* (2, 14, 5) {real, imag} */,
  {32'h3f89ec30, 32'h42b3821c} /* (2, 14, 4) {real, imag} */,
  {32'h40fb9bd8, 32'h41dace70} /* (2, 14, 3) {real, imag} */,
  {32'h42d4735a, 32'h42ed3686} /* (2, 14, 2) {real, imag} */,
  {32'hc28c0576, 32'h425a928e} /* (2, 14, 1) {real, imag} */,
  {32'hc33ded0e, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h421a6161, 32'h4249a864} /* (2, 13, 15) {real, imag} */,
  {32'h427b8b1c, 32'hc328b33b} /* (2, 13, 14) {real, imag} */,
  {32'h432e02c1, 32'h429d0a85} /* (2, 13, 13) {real, imag} */,
  {32'h434f1113, 32'hc30bfa15} /* (2, 13, 12) {real, imag} */,
  {32'h40be1500, 32'h421d33b8} /* (2, 13, 11) {real, imag} */,
  {32'h422e3fb0, 32'hc28ad844} /* (2, 13, 10) {real, imag} */,
  {32'hc28e6516, 32'h41c2ee84} /* (2, 13, 9) {real, imag} */,
  {32'hc14a8e70, 32'h00000000} /* (2, 13, 8) {real, imag} */,
  {32'hc28e6516, 32'hc1c2ee84} /* (2, 13, 7) {real, imag} */,
  {32'h422e3fb0, 32'h428ad844} /* (2, 13, 6) {real, imag} */,
  {32'h40be1500, 32'hc21d33b8} /* (2, 13, 5) {real, imag} */,
  {32'h434f1113, 32'h430bfa15} /* (2, 13, 4) {real, imag} */,
  {32'h432e02c1, 32'hc29d0a85} /* (2, 13, 3) {real, imag} */,
  {32'h427b8b1c, 32'h4328b33b} /* (2, 13, 2) {real, imag} */,
  {32'h421a6161, 32'hc249a864} /* (2, 13, 1) {real, imag} */,
  {32'hc3428089, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'hc29fcc00, 32'h428c74e0} /* (2, 12, 15) {real, imag} */,
  {32'hc0e62090, 32'hc34c39c3} /* (2, 12, 14) {real, imag} */,
  {32'h42b43432, 32'h41733b90} /* (2, 12, 13) {real, imag} */,
  {32'h42be0940, 32'h4307a51f} /* (2, 12, 12) {real, imag} */,
  {32'hc0e90738, 32'h411765c8} /* (2, 12, 11) {real, imag} */,
  {32'hc29c4ebf, 32'hc26fa915} /* (2, 12, 10) {real, imag} */,
  {32'hc1c5eeba, 32'h42181821} /* (2, 12, 9) {real, imag} */,
  {32'hc2852c3a, 32'h00000000} /* (2, 12, 8) {real, imag} */,
  {32'hc1c5eeba, 32'hc2181821} /* (2, 12, 7) {real, imag} */,
  {32'hc29c4ebf, 32'h426fa915} /* (2, 12, 6) {real, imag} */,
  {32'hc0e90738, 32'hc11765c8} /* (2, 12, 5) {real, imag} */,
  {32'h42be0940, 32'hc307a51f} /* (2, 12, 4) {real, imag} */,
  {32'h42b43432, 32'hc1733b90} /* (2, 12, 3) {real, imag} */,
  {32'hc0e62090, 32'h434c39c3} /* (2, 12, 2) {real, imag} */,
  {32'hc29fcc00, 32'hc28c74e0} /* (2, 12, 1) {real, imag} */,
  {32'h42b3058d, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h431ef980, 32'hc327aff6} /* (2, 11, 15) {real, imag} */,
  {32'hc2ca4858, 32'hc2ad832a} /* (2, 11, 14) {real, imag} */,
  {32'hc2e7d614, 32'hc16f67bc} /* (2, 11, 13) {real, imag} */,
  {32'h430ee49c, 32'h42c6d6e8} /* (2, 11, 12) {real, imag} */,
  {32'hc2942473, 32'h405f07e0} /* (2, 11, 11) {real, imag} */,
  {32'h430c95c7, 32'hc25904d0} /* (2, 11, 10) {real, imag} */,
  {32'h41ca385a, 32'hc2139efc} /* (2, 11, 9) {real, imag} */,
  {32'hc25f00d0, 32'h00000000} /* (2, 11, 8) {real, imag} */,
  {32'h41ca385a, 32'h42139efc} /* (2, 11, 7) {real, imag} */,
  {32'h430c95c7, 32'h425904d0} /* (2, 11, 6) {real, imag} */,
  {32'hc2942473, 32'hc05f07e0} /* (2, 11, 5) {real, imag} */,
  {32'h430ee49c, 32'hc2c6d6e8} /* (2, 11, 4) {real, imag} */,
  {32'hc2e7d614, 32'h416f67bc} /* (2, 11, 3) {real, imag} */,
  {32'hc2ca4858, 32'h42ad832a} /* (2, 11, 2) {real, imag} */,
  {32'h431ef980, 32'h4327aff6} /* (2, 11, 1) {real, imag} */,
  {32'h42fcf298, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'h433b122c, 32'hc2fed047} /* (2, 10, 15) {real, imag} */,
  {32'hc22e7b5d, 32'hc2e32dc4} /* (2, 10, 14) {real, imag} */,
  {32'h438c8ea4, 32'hbf9ec4c0} /* (2, 10, 13) {real, imag} */,
  {32'hc2e03b97, 32'hc1d073f3} /* (2, 10, 12) {real, imag} */,
  {32'hc282bb42, 32'hc1d8e4ae} /* (2, 10, 11) {real, imag} */,
  {32'hc24a0417, 32'h4239d1e8} /* (2, 10, 10) {real, imag} */,
  {32'hc0f3ce60, 32'hc2a4e2ad} /* (2, 10, 9) {real, imag} */,
  {32'h432922fa, 32'h00000000} /* (2, 10, 8) {real, imag} */,
  {32'hc0f3ce60, 32'h42a4e2ad} /* (2, 10, 7) {real, imag} */,
  {32'hc24a0417, 32'hc239d1e8} /* (2, 10, 6) {real, imag} */,
  {32'hc282bb42, 32'h41d8e4ae} /* (2, 10, 5) {real, imag} */,
  {32'hc2e03b97, 32'h41d073f3} /* (2, 10, 4) {real, imag} */,
  {32'h438c8ea4, 32'h3f9ec4c0} /* (2, 10, 3) {real, imag} */,
  {32'hc22e7b5d, 32'h42e32dc4} /* (2, 10, 2) {real, imag} */,
  {32'h433b122c, 32'h42fed047} /* (2, 10, 1) {real, imag} */,
  {32'h420d5244, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'h42520e9c, 32'hc21388b8} /* (2, 9, 15) {real, imag} */,
  {32'hc29dc343, 32'hc28e76f4} /* (2, 9, 14) {real, imag} */,
  {32'hc0a972f8, 32'hc2b9e516} /* (2, 9, 13) {real, imag} */,
  {32'hc2159258, 32'h41e80684} /* (2, 9, 12) {real, imag} */,
  {32'h425cd8c2, 32'h42cb2883} /* (2, 9, 11) {real, imag} */,
  {32'h410b96a8, 32'hc08d2b9c} /* (2, 9, 10) {real, imag} */,
  {32'h3f47c580, 32'h42c3aeb9} /* (2, 9, 9) {real, imag} */,
  {32'hc32e9ebd, 32'h00000000} /* (2, 9, 8) {real, imag} */,
  {32'h3f47c580, 32'hc2c3aeb9} /* (2, 9, 7) {real, imag} */,
  {32'h410b96a8, 32'h408d2b9c} /* (2, 9, 6) {real, imag} */,
  {32'h425cd8c2, 32'hc2cb2883} /* (2, 9, 5) {real, imag} */,
  {32'hc2159258, 32'hc1e80684} /* (2, 9, 4) {real, imag} */,
  {32'hc0a972f8, 32'h42b9e516} /* (2, 9, 3) {real, imag} */,
  {32'hc29dc343, 32'h428e76f4} /* (2, 9, 2) {real, imag} */,
  {32'h42520e9c, 32'h421388b8} /* (2, 9, 1) {real, imag} */,
  {32'h440693aa, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'h420a9cee, 32'hc333e8d0} /* (2, 8, 15) {real, imag} */,
  {32'h3fbf5e00, 32'hc347984b} /* (2, 8, 14) {real, imag} */,
  {32'hc3039fa6, 32'hc353067f} /* (2, 8, 13) {real, imag} */,
  {32'hc29accb8, 32'hc31ab8c8} /* (2, 8, 12) {real, imag} */,
  {32'h419b3284, 32'h42ca1c5a} /* (2, 8, 11) {real, imag} */,
  {32'hc21d943c, 32'h4299ae0a} /* (2, 8, 10) {real, imag} */,
  {32'h42fcccda, 32'h40d8a94c} /* (2, 8, 9) {real, imag} */,
  {32'hc1ea43d8, 32'h00000000} /* (2, 8, 8) {real, imag} */,
  {32'h42fcccda, 32'hc0d8a94c} /* (2, 8, 7) {real, imag} */,
  {32'hc21d943c, 32'hc299ae0a} /* (2, 8, 6) {real, imag} */,
  {32'h419b3284, 32'hc2ca1c5a} /* (2, 8, 5) {real, imag} */,
  {32'hc29accb8, 32'h431ab8c8} /* (2, 8, 4) {real, imag} */,
  {32'hc3039fa6, 32'h4353067f} /* (2, 8, 3) {real, imag} */,
  {32'h3fbf5e00, 32'h4347984b} /* (2, 8, 2) {real, imag} */,
  {32'h420a9cee, 32'h4333e8d0} /* (2, 8, 1) {real, imag} */,
  {32'h43c90b5a, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'h42b3d0b6, 32'hc38cb790} /* (2, 7, 15) {real, imag} */,
  {32'h429fcf63, 32'hc2e9dec4} /* (2, 7, 14) {real, imag} */,
  {32'hc29551c2, 32'hc11d7980} /* (2, 7, 13) {real, imag} */,
  {32'h434d4890, 32'hc2a05e84} /* (2, 7, 12) {real, imag} */,
  {32'h412bd936, 32'h42e32175} /* (2, 7, 11) {real, imag} */,
  {32'h432788ba, 32'h42110aee} /* (2, 7, 10) {real, imag} */,
  {32'h42151ce6, 32'hc31344d2} /* (2, 7, 9) {real, imag} */,
  {32'hc294ccac, 32'h00000000} /* (2, 7, 8) {real, imag} */,
  {32'h42151ce6, 32'h431344d2} /* (2, 7, 7) {real, imag} */,
  {32'h432788ba, 32'hc2110aee} /* (2, 7, 6) {real, imag} */,
  {32'h412bd936, 32'hc2e32175} /* (2, 7, 5) {real, imag} */,
  {32'h434d4890, 32'h42a05e84} /* (2, 7, 4) {real, imag} */,
  {32'hc29551c2, 32'h411d7980} /* (2, 7, 3) {real, imag} */,
  {32'h429fcf63, 32'h42e9dec4} /* (2, 7, 2) {real, imag} */,
  {32'h42b3d0b6, 32'h438cb790} /* (2, 7, 1) {real, imag} */,
  {32'h41a25b10, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'h42219b30, 32'hc3701f60} /* (2, 6, 15) {real, imag} */,
  {32'h419148de, 32'hc29ab260} /* (2, 6, 14) {real, imag} */,
  {32'h42403fdc, 32'h42b62d4d} /* (2, 6, 13) {real, imag} */,
  {32'h43321474, 32'h414cb7ee} /* (2, 6, 12) {real, imag} */,
  {32'h42aa0e42, 32'hc308b954} /* (2, 6, 11) {real, imag} */,
  {32'hc2cbe764, 32'h41e556e0} /* (2, 6, 10) {real, imag} */,
  {32'hc28bd40c, 32'h42821dcb} /* (2, 6, 9) {real, imag} */,
  {32'h40ff9bd0, 32'h00000000} /* (2, 6, 8) {real, imag} */,
  {32'hc28bd40c, 32'hc2821dcb} /* (2, 6, 7) {real, imag} */,
  {32'hc2cbe764, 32'hc1e556e0} /* (2, 6, 6) {real, imag} */,
  {32'h42aa0e42, 32'h4308b954} /* (2, 6, 5) {real, imag} */,
  {32'h43321474, 32'hc14cb7ee} /* (2, 6, 4) {real, imag} */,
  {32'h42403fdc, 32'hc2b62d4d} /* (2, 6, 3) {real, imag} */,
  {32'h419148de, 32'h429ab260} /* (2, 6, 2) {real, imag} */,
  {32'h42219b30, 32'h43701f60} /* (2, 6, 1) {real, imag} */,
  {32'hc3450796, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hc13663c8, 32'hc35ca142} /* (2, 5, 15) {real, imag} */,
  {32'h431cc83e, 32'h43229c2b} /* (2, 5, 14) {real, imag} */,
  {32'h41ef1938, 32'h42e52730} /* (2, 5, 13) {real, imag} */,
  {32'h4308612c, 32'h42b3c1c8} /* (2, 5, 12) {real, imag} */,
  {32'hc18a1a33, 32'h43114b82} /* (2, 5, 11) {real, imag} */,
  {32'hc2fc61ee, 32'hc19a1c79} /* (2, 5, 10) {real, imag} */,
  {32'hc29145b6, 32'hc1965774} /* (2, 5, 9) {real, imag} */,
  {32'h4106c560, 32'h00000000} /* (2, 5, 8) {real, imag} */,
  {32'hc29145b6, 32'h41965774} /* (2, 5, 7) {real, imag} */,
  {32'hc2fc61ee, 32'h419a1c79} /* (2, 5, 6) {real, imag} */,
  {32'hc18a1a33, 32'hc3114b82} /* (2, 5, 5) {real, imag} */,
  {32'h4308612c, 32'hc2b3c1c8} /* (2, 5, 4) {real, imag} */,
  {32'h41ef1938, 32'hc2e52730} /* (2, 5, 3) {real, imag} */,
  {32'h431cc83e, 32'hc3229c2b} /* (2, 5, 2) {real, imag} */,
  {32'hc13663c8, 32'h435ca142} /* (2, 5, 1) {real, imag} */,
  {32'hc3c8d206, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hc2c6c65e, 32'hc3627d60} /* (2, 4, 15) {real, imag} */,
  {32'h430bcc56, 32'h43305289} /* (2, 4, 14) {real, imag} */,
  {32'hc110d4d4, 32'h4261eb58} /* (2, 4, 13) {real, imag} */,
  {32'hbfb3ad00, 32'h4203759c} /* (2, 4, 12) {real, imag} */,
  {32'h3d1dd400, 32'h42831618} /* (2, 4, 11) {real, imag} */,
  {32'h42b8f0d1, 32'h41cefafe} /* (2, 4, 10) {real, imag} */,
  {32'hc2f67ede, 32'h422cc337} /* (2, 4, 9) {real, imag} */,
  {32'hc30bd4b3, 32'h00000000} /* (2, 4, 8) {real, imag} */,
  {32'hc2f67ede, 32'hc22cc337} /* (2, 4, 7) {real, imag} */,
  {32'h42b8f0d1, 32'hc1cefafe} /* (2, 4, 6) {real, imag} */,
  {32'h3d1dd400, 32'hc2831618} /* (2, 4, 5) {real, imag} */,
  {32'hbfb3ad00, 32'hc203759c} /* (2, 4, 4) {real, imag} */,
  {32'hc110d4d4, 32'hc261eb58} /* (2, 4, 3) {real, imag} */,
  {32'h430bcc56, 32'hc3305289} /* (2, 4, 2) {real, imag} */,
  {32'hc2c6c65e, 32'h43627d60} /* (2, 4, 1) {real, imag} */,
  {32'hc3a1089c, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hc2108d93, 32'hc34bf0cc} /* (2, 3, 15) {real, imag} */,
  {32'hc296dac2, 32'h4373e67d} /* (2, 3, 14) {real, imag} */,
  {32'hbe952000, 32'h427c9532} /* (2, 3, 13) {real, imag} */,
  {32'h41ed7ec8, 32'h42b57600} /* (2, 3, 12) {real, imag} */,
  {32'h42c7c484, 32'h426245b8} /* (2, 3, 11) {real, imag} */,
  {32'h42d7c414, 32'hc2e3d976} /* (2, 3, 10) {real, imag} */,
  {32'hc253d4e1, 32'hc26f6e2c} /* (2, 3, 9) {real, imag} */,
  {32'h4299d36c, 32'h00000000} /* (2, 3, 8) {real, imag} */,
  {32'hc253d4e1, 32'h426f6e2c} /* (2, 3, 7) {real, imag} */,
  {32'h42d7c414, 32'h42e3d976} /* (2, 3, 6) {real, imag} */,
  {32'h42c7c484, 32'hc26245b8} /* (2, 3, 5) {real, imag} */,
  {32'h41ed7ec8, 32'hc2b57600} /* (2, 3, 4) {real, imag} */,
  {32'hbe952000, 32'hc27c9532} /* (2, 3, 3) {real, imag} */,
  {32'hc296dac2, 32'hc373e67d} /* (2, 3, 2) {real, imag} */,
  {32'hc2108d93, 32'h434bf0cc} /* (2, 3, 1) {real, imag} */,
  {32'hc388b840, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hc2c676fe, 32'hc37abf70} /* (2, 2, 15) {real, imag} */,
  {32'hc1dcf0aa, 32'hc291d556} /* (2, 2, 14) {real, imag} */,
  {32'h41ba89ca, 32'h43052045} /* (2, 2, 13) {real, imag} */,
  {32'h424ca200, 32'hc303ab5a} /* (2, 2, 12) {real, imag} */,
  {32'h407ce110, 32'h42423a08} /* (2, 2, 11) {real, imag} */,
  {32'h41e2cfbc, 32'h42b4ac5a} /* (2, 2, 10) {real, imag} */,
  {32'hc18bd6ce, 32'h42be6524} /* (2, 2, 9) {real, imag} */,
  {32'hc01e89f8, 32'h00000000} /* (2, 2, 8) {real, imag} */,
  {32'hc18bd6ce, 32'hc2be6524} /* (2, 2, 7) {real, imag} */,
  {32'h41e2cfbc, 32'hc2b4ac5a} /* (2, 2, 6) {real, imag} */,
  {32'h407ce110, 32'hc2423a08} /* (2, 2, 5) {real, imag} */,
  {32'h424ca200, 32'h4303ab5a} /* (2, 2, 4) {real, imag} */,
  {32'h41ba89ca, 32'hc3052045} /* (2, 2, 3) {real, imag} */,
  {32'hc1dcf0aa, 32'h4291d556} /* (2, 2, 2) {real, imag} */,
  {32'hc2c676fe, 32'h437abf70} /* (2, 2, 1) {real, imag} */,
  {32'hc38469d3, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hc34f201a, 32'hc3429f78} /* (2, 1, 15) {real, imag} */,
  {32'hc2935edb, 32'hc0a9d62c} /* (2, 1, 14) {real, imag} */,
  {32'h432b2732, 32'h42f6aea1} /* (2, 1, 13) {real, imag} */,
  {32'hc296bb55, 32'hc17b0344} /* (2, 1, 12) {real, imag} */,
  {32'h431a37ca, 32'h4189c11c} /* (2, 1, 11) {real, imag} */,
  {32'hc296ba3d, 32'h42a531fa} /* (2, 1, 10) {real, imag} */,
  {32'h42d28247, 32'hc2c777a3} /* (2, 1, 9) {real, imag} */,
  {32'hc2b953a8, 32'h00000000} /* (2, 1, 8) {real, imag} */,
  {32'h42d28247, 32'h42c777a3} /* (2, 1, 7) {real, imag} */,
  {32'hc296ba3d, 32'hc2a531fa} /* (2, 1, 6) {real, imag} */,
  {32'h431a37ca, 32'hc189c11c} /* (2, 1, 5) {real, imag} */,
  {32'hc296bb55, 32'h417b0344} /* (2, 1, 4) {real, imag} */,
  {32'h432b2732, 32'hc2f6aea1} /* (2, 1, 3) {real, imag} */,
  {32'hc2935edb, 32'h40a9d62c} /* (2, 1, 2) {real, imag} */,
  {32'hc34f201a, 32'h43429f78} /* (2, 1, 1) {real, imag} */,
  {32'hc39cd248, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hc2e51699, 32'hc2d11d00} /* (2, 0, 15) {real, imag} */,
  {32'hc2bd6d80, 32'h42cdb8aa} /* (2, 0, 14) {real, imag} */,
  {32'h419db756, 32'h432c1823} /* (2, 0, 13) {real, imag} */,
  {32'h4086e140, 32'hc232ca06} /* (2, 0, 12) {real, imag} */,
  {32'h427c781c, 32'hc3099adc} /* (2, 0, 11) {real, imag} */,
  {32'hc29cd9c6, 32'h41841ada} /* (2, 0, 10) {real, imag} */,
  {32'h41a43cba, 32'hc0bd59a4} /* (2, 0, 9) {real, imag} */,
  {32'h4010f9e0, 32'h00000000} /* (2, 0, 8) {real, imag} */,
  {32'h41a43cba, 32'h40bd59a4} /* (2, 0, 7) {real, imag} */,
  {32'hc29cd9c6, 32'hc1841ada} /* (2, 0, 6) {real, imag} */,
  {32'h427c781c, 32'h43099adc} /* (2, 0, 5) {real, imag} */,
  {32'h4086e140, 32'h4232ca06} /* (2, 0, 4) {real, imag} */,
  {32'h419db756, 32'hc32c1823} /* (2, 0, 3) {real, imag} */,
  {32'hc2bd6d80, 32'hc2cdb8aa} /* (2, 0, 2) {real, imag} */,
  {32'hc2e51699, 32'h42d11d00} /* (2, 0, 1) {real, imag} */,
  {32'hc2a4c9c8, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hc3045048, 32'hc3432e8e} /* (1, 15, 15) {real, imag} */,
  {32'h424b7efc, 32'hc0f1858c} /* (1, 15, 14) {real, imag} */,
  {32'h421b554a, 32'h4216015c} /* (1, 15, 13) {real, imag} */,
  {32'hc215b266, 32'hc2957761} /* (1, 15, 12) {real, imag} */,
  {32'h416c91e6, 32'h4245a8c3} /* (1, 15, 11) {real, imag} */,
  {32'h41e1036c, 32'hc243b8e6} /* (1, 15, 10) {real, imag} */,
  {32'hc276dd70, 32'hc13569e8} /* (1, 15, 9) {real, imag} */,
  {32'h41da94a4, 32'h00000000} /* (1, 15, 8) {real, imag} */,
  {32'hc276dd70, 32'h413569e8} /* (1, 15, 7) {real, imag} */,
  {32'h41e1036c, 32'h4243b8e6} /* (1, 15, 6) {real, imag} */,
  {32'h416c91e6, 32'hc245a8c3} /* (1, 15, 5) {real, imag} */,
  {32'hc215b266, 32'h42957761} /* (1, 15, 4) {real, imag} */,
  {32'h421b554a, 32'hc216015c} /* (1, 15, 3) {real, imag} */,
  {32'h424b7efc, 32'h40f1858c} /* (1, 15, 2) {real, imag} */,
  {32'hc3045048, 32'h43432e8e} /* (1, 15, 1) {real, imag} */,
  {32'hc351178e, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'hc3273cd4, 32'hc300c558} /* (1, 14, 15) {real, imag} */,
  {32'h4213bb7e, 32'hc2d6f665} /* (1, 14, 14) {real, imag} */,
  {32'h4317252f, 32'h424826bf} /* (1, 14, 13) {real, imag} */,
  {32'hc183c6de, 32'h4173f0c0} /* (1, 14, 12) {real, imag} */,
  {32'h41f2b02a, 32'h42bc4581} /* (1, 14, 11) {real, imag} */,
  {32'hc2b00e8d, 32'h42ddafeb} /* (1, 14, 10) {real, imag} */,
  {32'hc2a0a221, 32'hc2dda806} /* (1, 14, 9) {real, imag} */,
  {32'hc083b2f8, 32'h00000000} /* (1, 14, 8) {real, imag} */,
  {32'hc2a0a221, 32'h42dda806} /* (1, 14, 7) {real, imag} */,
  {32'hc2b00e8d, 32'hc2ddafeb} /* (1, 14, 6) {real, imag} */,
  {32'h41f2b02a, 32'hc2bc4581} /* (1, 14, 5) {real, imag} */,
  {32'hc183c6de, 32'hc173f0c0} /* (1, 14, 4) {real, imag} */,
  {32'h4317252f, 32'hc24826bf} /* (1, 14, 3) {real, imag} */,
  {32'h4213bb7e, 32'h42d6f665} /* (1, 14, 2) {real, imag} */,
  {32'hc3273cd4, 32'h4300c558} /* (1, 14, 1) {real, imag} */,
  {32'hc278e0f0, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'hc10e495e, 32'hc22718f4} /* (1, 13, 15) {real, imag} */,
  {32'h4216d866, 32'hc2069bfc} /* (1, 13, 14) {real, imag} */,
  {32'h430acc0e, 32'h417a7338} /* (1, 13, 13) {real, imag} */,
  {32'h42c16128, 32'hc29625b5} /* (1, 13, 12) {real, imag} */,
  {32'hc16804f8, 32'hc22f015a} /* (1, 13, 11) {real, imag} */,
  {32'h42b576fb, 32'h42aa7097} /* (1, 13, 10) {real, imag} */,
  {32'h42090ebc, 32'h4278a806} /* (1, 13, 9) {real, imag} */,
  {32'h4284f8fe, 32'h00000000} /* (1, 13, 8) {real, imag} */,
  {32'h42090ebc, 32'hc278a806} /* (1, 13, 7) {real, imag} */,
  {32'h42b576fb, 32'hc2aa7097} /* (1, 13, 6) {real, imag} */,
  {32'hc16804f8, 32'h422f015a} /* (1, 13, 5) {real, imag} */,
  {32'h42c16128, 32'h429625b5} /* (1, 13, 4) {real, imag} */,
  {32'h430acc0e, 32'hc17a7338} /* (1, 13, 3) {real, imag} */,
  {32'h4216d866, 32'h42069bfc} /* (1, 13, 2) {real, imag} */,
  {32'hc10e495e, 32'h422718f4} /* (1, 13, 1) {real, imag} */,
  {32'h4205b7de, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'h439bc0ae, 32'hc28e47d2} /* (1, 12, 15) {real, imag} */,
  {32'hc2e53f80, 32'h4335c03a} /* (1, 12, 14) {real, imag} */,
  {32'hc242bd30, 32'h425bbc04} /* (1, 12, 13) {real, imag} */,
  {32'h42821639, 32'h426748aa} /* (1, 12, 12) {real, imag} */,
  {32'h42798cdc, 32'hc2738644} /* (1, 12, 11) {real, imag} */,
  {32'h42161acc, 32'hc21b8dcb} /* (1, 12, 10) {real, imag} */,
  {32'hc208f8a2, 32'h42063866} /* (1, 12, 9) {real, imag} */,
  {32'hc1c3aec4, 32'h00000000} /* (1, 12, 8) {real, imag} */,
  {32'hc208f8a2, 32'hc2063866} /* (1, 12, 7) {real, imag} */,
  {32'h42161acc, 32'h421b8dcb} /* (1, 12, 6) {real, imag} */,
  {32'h42798cdc, 32'h42738644} /* (1, 12, 5) {real, imag} */,
  {32'h42821639, 32'hc26748aa} /* (1, 12, 4) {real, imag} */,
  {32'hc242bd30, 32'hc25bbc04} /* (1, 12, 3) {real, imag} */,
  {32'hc2e53f80, 32'hc335c03a} /* (1, 12, 2) {real, imag} */,
  {32'h439bc0ae, 32'h428e47d2} /* (1, 12, 1) {real, imag} */,
  {32'hc2bad7ec, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'h4284d5a4, 32'hc38d1680} /* (1, 11, 15) {real, imag} */,
  {32'hc305e3df, 32'hc30f9be3} /* (1, 11, 14) {real, imag} */,
  {32'h418f43b4, 32'h418ac974} /* (1, 11, 13) {real, imag} */,
  {32'h42db148e, 32'h43714222} /* (1, 11, 12) {real, imag} */,
  {32'h42b06a38, 32'h421bb061} /* (1, 11, 11) {real, imag} */,
  {32'hc23f75a4, 32'h4071ebf0} /* (1, 11, 10) {real, imag} */,
  {32'hc2a66132, 32'h418de29c} /* (1, 11, 9) {real, imag} */,
  {32'h3edaa980, 32'h00000000} /* (1, 11, 8) {real, imag} */,
  {32'hc2a66132, 32'hc18de29c} /* (1, 11, 7) {real, imag} */,
  {32'hc23f75a4, 32'hc071ebf0} /* (1, 11, 6) {real, imag} */,
  {32'h42b06a38, 32'hc21bb061} /* (1, 11, 5) {real, imag} */,
  {32'h42db148e, 32'hc3714222} /* (1, 11, 4) {real, imag} */,
  {32'h418f43b4, 32'hc18ac974} /* (1, 11, 3) {real, imag} */,
  {32'hc305e3df, 32'h430f9be3} /* (1, 11, 2) {real, imag} */,
  {32'h4284d5a4, 32'h438d1680} /* (1, 11, 1) {real, imag} */,
  {32'h43a36075, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'hc2473daa, 32'hc3afdd14} /* (1, 10, 15) {real, imag} */,
  {32'h4211837c, 32'hc264b076} /* (1, 10, 14) {real, imag} */,
  {32'hc2ff63c6, 32'hc2a449b4} /* (1, 10, 13) {real, imag} */,
  {32'hc21aff44, 32'hc21d4f13} /* (1, 10, 12) {real, imag} */,
  {32'hc291698e, 32'hc2e2703e} /* (1, 10, 11) {real, imag} */,
  {32'h41ca3e5a, 32'h42fb91a8} /* (1, 10, 10) {real, imag} */,
  {32'hc27131f1, 32'h426e9dca} /* (1, 10, 9) {real, imag} */,
  {32'h424adb78, 32'h00000000} /* (1, 10, 8) {real, imag} */,
  {32'hc27131f1, 32'hc26e9dca} /* (1, 10, 7) {real, imag} */,
  {32'h41ca3e5a, 32'hc2fb91a8} /* (1, 10, 6) {real, imag} */,
  {32'hc291698e, 32'h42e2703e} /* (1, 10, 5) {real, imag} */,
  {32'hc21aff44, 32'h421d4f13} /* (1, 10, 4) {real, imag} */,
  {32'hc2ff63c6, 32'h42a449b4} /* (1, 10, 3) {real, imag} */,
  {32'h4211837c, 32'h4264b076} /* (1, 10, 2) {real, imag} */,
  {32'hc2473daa, 32'h43afdd14} /* (1, 10, 1) {real, imag} */,
  {32'h43c5f761, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'h429e598c, 32'hc2c17648} /* (1, 9, 15) {real, imag} */,
  {32'h41e90dfe, 32'h41ea1294} /* (1, 9, 14) {real, imag} */,
  {32'h430a7408, 32'hc22a5ce5} /* (1, 9, 13) {real, imag} */,
  {32'h420a2c0a, 32'hc21727ea} /* (1, 9, 12) {real, imag} */,
  {32'h4285d9a4, 32'h41b5982c} /* (1, 9, 11) {real, imag} */,
  {32'hc2c89d20, 32'hc28ddc88} /* (1, 9, 10) {real, imag} */,
  {32'h418c8b10, 32'h42b849ab} /* (1, 9, 9) {real, imag} */,
  {32'hc1e018de, 32'h00000000} /* (1, 9, 8) {real, imag} */,
  {32'h418c8b10, 32'hc2b849ab} /* (1, 9, 7) {real, imag} */,
  {32'hc2c89d20, 32'h428ddc88} /* (1, 9, 6) {real, imag} */,
  {32'h4285d9a4, 32'hc1b5982c} /* (1, 9, 5) {real, imag} */,
  {32'h420a2c0a, 32'h421727ea} /* (1, 9, 4) {real, imag} */,
  {32'h430a7408, 32'h422a5ce5} /* (1, 9, 3) {real, imag} */,
  {32'h41e90dfe, 32'hc1ea1294} /* (1, 9, 2) {real, imag} */,
  {32'h429e598c, 32'h42c17648} /* (1, 9, 1) {real, imag} */,
  {32'h43fc488c, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'h4321b04c, 32'hc1dac8e0} /* (1, 8, 15) {real, imag} */,
  {32'hc2497768, 32'h427a5828} /* (1, 8, 14) {real, imag} */,
  {32'h41606f9c, 32'hc3071736} /* (1, 8, 13) {real, imag} */,
  {32'h421671a0, 32'hc20524be} /* (1, 8, 12) {real, imag} */,
  {32'h4217de87, 32'h41edbbcb} /* (1, 8, 11) {real, imag} */,
  {32'hc2b77be0, 32'hc2d9046e} /* (1, 8, 10) {real, imag} */,
  {32'h42a57df2, 32'h428ea4a6} /* (1, 8, 9) {real, imag} */,
  {32'h415649f5, 32'h00000000} /* (1, 8, 8) {real, imag} */,
  {32'h42a57df2, 32'hc28ea4a6} /* (1, 8, 7) {real, imag} */,
  {32'hc2b77be0, 32'h42d9046e} /* (1, 8, 6) {real, imag} */,
  {32'h4217de87, 32'hc1edbbcb} /* (1, 8, 5) {real, imag} */,
  {32'h421671a0, 32'h420524be} /* (1, 8, 4) {real, imag} */,
  {32'h41606f9c, 32'h43071736} /* (1, 8, 3) {real, imag} */,
  {32'hc2497768, 32'hc27a5828} /* (1, 8, 2) {real, imag} */,
  {32'h4321b04c, 32'h41dac8e0} /* (1, 8, 1) {real, imag} */,
  {32'h43a481c0, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'h4395d8db, 32'hc2caa7e4} /* (1, 7, 15) {real, imag} */,
  {32'h42e4055a, 32'h42d53eef} /* (1, 7, 14) {real, imag} */,
  {32'hc0f652f0, 32'h42cf5d46} /* (1, 7, 13) {real, imag} */,
  {32'h433a31bc, 32'hc1fae2cc} /* (1, 7, 12) {real, imag} */,
  {32'h42656519, 32'h43198e52} /* (1, 7, 11) {real, imag} */,
  {32'h42660587, 32'hc2df79fa} /* (1, 7, 10) {real, imag} */,
  {32'h43062855, 32'h42e68a1d} /* (1, 7, 9) {real, imag} */,
  {32'h425213bd, 32'h00000000} /* (1, 7, 8) {real, imag} */,
  {32'h43062855, 32'hc2e68a1d} /* (1, 7, 7) {real, imag} */,
  {32'h42660587, 32'h42df79fa} /* (1, 7, 6) {real, imag} */,
  {32'h42656519, 32'hc3198e52} /* (1, 7, 5) {real, imag} */,
  {32'h433a31bc, 32'h41fae2cc} /* (1, 7, 4) {real, imag} */,
  {32'hc0f652f0, 32'hc2cf5d46} /* (1, 7, 3) {real, imag} */,
  {32'h42e4055a, 32'hc2d53eef} /* (1, 7, 2) {real, imag} */,
  {32'h4395d8db, 32'h42caa7e4} /* (1, 7, 1) {real, imag} */,
  {32'h419dce80, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'h42796c66, 32'hc3941638} /* (1, 6, 15) {real, imag} */,
  {32'h430eb85e, 32'h41cbda80} /* (1, 6, 14) {real, imag} */,
  {32'h42e5ded6, 32'h41f8ee32} /* (1, 6, 13) {real, imag} */,
  {32'h436dcb17, 32'hc1d64eae} /* (1, 6, 12) {real, imag} */,
  {32'h4335d0e5, 32'h435ff7f5} /* (1, 6, 11) {real, imag} */,
  {32'hc25ba96d, 32'h42621a9c} /* (1, 6, 10) {real, imag} */,
  {32'h42840b49, 32'hc1266f3e} /* (1, 6, 9) {real, imag} */,
  {32'h41d9573f, 32'h00000000} /* (1, 6, 8) {real, imag} */,
  {32'h42840b49, 32'h41266f3e} /* (1, 6, 7) {real, imag} */,
  {32'hc25ba96d, 32'hc2621a9c} /* (1, 6, 6) {real, imag} */,
  {32'h4335d0e5, 32'hc35ff7f5} /* (1, 6, 5) {real, imag} */,
  {32'h436dcb17, 32'h41d64eae} /* (1, 6, 4) {real, imag} */,
  {32'h42e5ded6, 32'hc1f8ee32} /* (1, 6, 3) {real, imag} */,
  {32'h430eb85e, 32'hc1cbda80} /* (1, 6, 2) {real, imag} */,
  {32'h42796c66, 32'h43941638} /* (1, 6, 1) {real, imag} */,
  {32'hc2a75730, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'h42de185c, 32'hc301b99d} /* (1, 5, 15) {real, imag} */,
  {32'h4224627c, 32'h432470a3} /* (1, 5, 14) {real, imag} */,
  {32'h42736cb0, 32'h43583b3c} /* (1, 5, 13) {real, imag} */,
  {32'h43048a0f, 32'hc2a0829c} /* (1, 5, 12) {real, imag} */,
  {32'h4193834c, 32'h42392a2f} /* (1, 5, 11) {real, imag} */,
  {32'h42afd0ca, 32'h41dc019a} /* (1, 5, 10) {real, imag} */,
  {32'hc286050c, 32'hc1935a04} /* (1, 5, 9) {real, imag} */,
  {32'h4271a53d, 32'h00000000} /* (1, 5, 8) {real, imag} */,
  {32'hc286050c, 32'h41935a04} /* (1, 5, 7) {real, imag} */,
  {32'h42afd0ca, 32'hc1dc019a} /* (1, 5, 6) {real, imag} */,
  {32'h4193834c, 32'hc2392a2f} /* (1, 5, 5) {real, imag} */,
  {32'h43048a0f, 32'h42a0829c} /* (1, 5, 4) {real, imag} */,
  {32'h42736cb0, 32'hc3583b3c} /* (1, 5, 3) {real, imag} */,
  {32'h4224627c, 32'hc32470a3} /* (1, 5, 2) {real, imag} */,
  {32'h42de185c, 32'h4301b99d} /* (1, 5, 1) {real, imag} */,
  {32'h40ab04c0, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'h4220c950, 32'hc2eae284} /* (1, 4, 15) {real, imag} */,
  {32'hbf76c640, 32'h435b2cec} /* (1, 4, 14) {real, imag} */,
  {32'hc1d6c838, 32'h437af957} /* (1, 4, 13) {real, imag} */,
  {32'h409da1cc, 32'h41fe864c} /* (1, 4, 12) {real, imag} */,
  {32'h431acb77, 32'h434cacc3} /* (1, 4, 11) {real, imag} */,
  {32'h42497288, 32'hc3227791} /* (1, 4, 10) {real, imag} */,
  {32'h4256e452, 32'hc1918e97} /* (1, 4, 9) {real, imag} */,
  {32'h42067b12, 32'h00000000} /* (1, 4, 8) {real, imag} */,
  {32'h4256e452, 32'h41918e97} /* (1, 4, 7) {real, imag} */,
  {32'h42497288, 32'h43227791} /* (1, 4, 6) {real, imag} */,
  {32'h431acb77, 32'hc34cacc3} /* (1, 4, 5) {real, imag} */,
  {32'h409da1cc, 32'hc1fe864c} /* (1, 4, 4) {real, imag} */,
  {32'hc1d6c838, 32'hc37af957} /* (1, 4, 3) {real, imag} */,
  {32'hbf76c640, 32'hc35b2cec} /* (1, 4, 2) {real, imag} */,
  {32'h4220c950, 32'h42eae284} /* (1, 4, 1) {real, imag} */,
  {32'hc3329d90, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hc20ddb7a, 32'hc401093d} /* (1, 3, 15) {real, imag} */,
  {32'h42dea385, 32'h43222b4b} /* (1, 3, 14) {real, imag} */,
  {32'hc31e1cc6, 32'h41c6024c} /* (1, 3, 13) {real, imag} */,
  {32'hc1d4a3ea, 32'hc2c5a5e7} /* (1, 3, 12) {real, imag} */,
  {32'h42723388, 32'h4293fe7c} /* (1, 3, 11) {real, imag} */,
  {32'hc2163fb2, 32'h42e5e0f3} /* (1, 3, 10) {real, imag} */,
  {32'h42ffb6a4, 32'hc2da339d} /* (1, 3, 9) {real, imag} */,
  {32'h4203eb5d, 32'h00000000} /* (1, 3, 8) {real, imag} */,
  {32'h42ffb6a4, 32'h42da339d} /* (1, 3, 7) {real, imag} */,
  {32'hc2163fb2, 32'hc2e5e0f3} /* (1, 3, 6) {real, imag} */,
  {32'h42723388, 32'hc293fe7c} /* (1, 3, 5) {real, imag} */,
  {32'hc1d4a3ea, 32'h42c5a5e7} /* (1, 3, 4) {real, imag} */,
  {32'hc31e1cc6, 32'hc1c6024c} /* (1, 3, 3) {real, imag} */,
  {32'h42dea385, 32'hc3222b4b} /* (1, 3, 2) {real, imag} */,
  {32'hc20ddb7a, 32'h4401093d} /* (1, 3, 1) {real, imag} */,
  {32'hc3820ba0, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hc38adf2a, 32'hc3844848} /* (1, 2, 15) {real, imag} */,
  {32'hc2310b56, 32'h40a93e80} /* (1, 2, 14) {real, imag} */,
  {32'h423daaa5, 32'h41ffdde2} /* (1, 2, 13) {real, imag} */,
  {32'h42868496, 32'hc316c332} /* (1, 2, 12) {real, imag} */,
  {32'h429bfa3c, 32'h42692e06} /* (1, 2, 11) {real, imag} */,
  {32'h42b09f17, 32'h40c1acf0} /* (1, 2, 10) {real, imag} */,
  {32'h43159b12, 32'hc1d74c5a} /* (1, 2, 9) {real, imag} */,
  {32'h4210db12, 32'h00000000} /* (1, 2, 8) {real, imag} */,
  {32'h43159b12, 32'h41d74c5a} /* (1, 2, 7) {real, imag} */,
  {32'h42b09f17, 32'hc0c1acf0} /* (1, 2, 6) {real, imag} */,
  {32'h429bfa3c, 32'hc2692e06} /* (1, 2, 5) {real, imag} */,
  {32'h42868496, 32'h4316c332} /* (1, 2, 4) {real, imag} */,
  {32'h423daaa5, 32'hc1ffdde2} /* (1, 2, 3) {real, imag} */,
  {32'hc2310b56, 32'hc0a93e80} /* (1, 2, 2) {real, imag} */,
  {32'hc38adf2a, 32'h43844848} /* (1, 2, 1) {real, imag} */,
  {32'hc34e6fae, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hc36288f0, 32'hc2a90fc1} /* (1, 1, 15) {real, imag} */,
  {32'hc28d924b, 32'hc14847a2} /* (1, 1, 14) {real, imag} */,
  {32'h431622aa, 32'h4351e797} /* (1, 1, 13) {real, imag} */,
  {32'h4342b770, 32'h42baf9f7} /* (1, 1, 12) {real, imag} */,
  {32'hc24bff5a, 32'hc18c3bd6} /* (1, 1, 11) {real, imag} */,
  {32'h425b6eac, 32'hc281843b} /* (1, 1, 10) {real, imag} */,
  {32'hc2f83c42, 32'h42dfe1c5} /* (1, 1, 9) {real, imag} */,
  {32'hc2abd4a1, 32'h00000000} /* (1, 1, 8) {real, imag} */,
  {32'hc2f83c42, 32'hc2dfe1c5} /* (1, 1, 7) {real, imag} */,
  {32'h425b6eac, 32'h4281843b} /* (1, 1, 6) {real, imag} */,
  {32'hc24bff5a, 32'h418c3bd6} /* (1, 1, 5) {real, imag} */,
  {32'h4342b770, 32'hc2baf9f7} /* (1, 1, 4) {real, imag} */,
  {32'h431622aa, 32'hc351e797} /* (1, 1, 3) {real, imag} */,
  {32'hc28d924b, 32'h414847a2} /* (1, 1, 2) {real, imag} */,
  {32'hc36288f0, 32'h42a90fc1} /* (1, 1, 1) {real, imag} */,
  {32'hc302f72e, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hc29d67cf, 32'hc3262e6d} /* (1, 0, 15) {real, imag} */,
  {32'hc21be232, 32'hc2d98190} /* (1, 0, 14) {real, imag} */,
  {32'h4262c17d, 32'h42d9426d} /* (1, 0, 13) {real, imag} */,
  {32'hc17b4860, 32'hc02aff50} /* (1, 0, 12) {real, imag} */,
  {32'hc280aba2, 32'hc14bc58e} /* (1, 0, 11) {real, imag} */,
  {32'hc2611d95, 32'h42659459} /* (1, 0, 10) {real, imag} */,
  {32'h40d6a800, 32'hc1575922} /* (1, 0, 9) {real, imag} */,
  {32'h413d7cb9, 32'h00000000} /* (1, 0, 8) {real, imag} */,
  {32'h40d6a800, 32'h41575922} /* (1, 0, 7) {real, imag} */,
  {32'hc2611d95, 32'hc2659459} /* (1, 0, 6) {real, imag} */,
  {32'hc280aba2, 32'h414bc58e} /* (1, 0, 5) {real, imag} */,
  {32'hc17b4860, 32'h402aff50} /* (1, 0, 4) {real, imag} */,
  {32'h4262c17d, 32'hc2d9426d} /* (1, 0, 3) {real, imag} */,
  {32'hc21be232, 32'h42d98190} /* (1, 0, 2) {real, imag} */,
  {32'hc29d67cf, 32'h43262e6d} /* (1, 0, 1) {real, imag} */,
  {32'hc37b28e3, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'h417a01d8, 32'hc2c2644a} /* (0, 15, 15) {real, imag} */,
  {32'hc0004b88, 32'hc2a9b496} /* (0, 15, 14) {real, imag} */,
  {32'h41755ef4, 32'h42983751} /* (0, 15, 13) {real, imag} */,
  {32'h41622f6c, 32'hc296138f} /* (0, 15, 12) {real, imag} */,
  {32'hc2a8a0e4, 32'hc15c1d04} /* (0, 15, 11) {real, imag} */,
  {32'hc1cbe260, 32'h412c2ae4} /* (0, 15, 10) {real, imag} */,
  {32'hc1dbf75d, 32'h417ea768} /* (0, 15, 9) {real, imag} */,
  {32'hc179ee00, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'hc1dbf75d, 32'hc17ea768} /* (0, 15, 7) {real, imag} */,
  {32'hc1cbe260, 32'hc12c2ae4} /* (0, 15, 6) {real, imag} */,
  {32'hc2a8a0e4, 32'h415c1d04} /* (0, 15, 5) {real, imag} */,
  {32'h41622f6c, 32'h4296138f} /* (0, 15, 4) {real, imag} */,
  {32'h41755ef4, 32'hc2983751} /* (0, 15, 3) {real, imag} */,
  {32'hc0004b88, 32'h42a9b496} /* (0, 15, 2) {real, imag} */,
  {32'h417a01d8, 32'h42c2644a} /* (0, 15, 1) {real, imag} */,
  {32'hc353a139, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h42a8c490, 32'hc2d22260} /* (0, 14, 15) {real, imag} */,
  {32'h41f6795a, 32'hc1f97d67} /* (0, 14, 14) {real, imag} */,
  {32'h4343f314, 32'h425ce1f2} /* (0, 14, 13) {real, imag} */,
  {32'hc0eb0130, 32'hc2d6f154} /* (0, 14, 12) {real, imag} */,
  {32'hc306b169, 32'h412ca858} /* (0, 14, 11) {real, imag} */,
  {32'h429cf75a, 32'h429c2792} /* (0, 14, 10) {real, imag} */,
  {32'hc25654ac, 32'hc200fd5e} /* (0, 14, 9) {real, imag} */,
  {32'hc22d3eb0, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'hc25654ac, 32'h4200fd5e} /* (0, 14, 7) {real, imag} */,
  {32'h429cf75a, 32'hc29c2792} /* (0, 14, 6) {real, imag} */,
  {32'hc306b169, 32'hc12ca858} /* (0, 14, 5) {real, imag} */,
  {32'hc0eb0130, 32'h42d6f154} /* (0, 14, 4) {real, imag} */,
  {32'h4343f314, 32'hc25ce1f2} /* (0, 14, 3) {real, imag} */,
  {32'h41f6795a, 32'h41f97d67} /* (0, 14, 2) {real, imag} */,
  {32'h42a8c490, 32'h42d22260} /* (0, 14, 1) {real, imag} */,
  {32'hc1ea6cb6, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h42d4c0b0, 32'hc30e799e} /* (0, 13, 15) {real, imag} */,
  {32'hc0d8da14, 32'h425f898b} /* (0, 13, 14) {real, imag} */,
  {32'h412e21e0, 32'h424eff2d} /* (0, 13, 13) {real, imag} */,
  {32'h40add2f9, 32'h424bc0fa} /* (0, 13, 12) {real, imag} */,
  {32'hc2813847, 32'hc0bc0ea8} /* (0, 13, 11) {real, imag} */,
  {32'hc21053dd, 32'h418d9c35} /* (0, 13, 10) {real, imag} */,
  {32'h42311295, 32'h41c96d04} /* (0, 13, 9) {real, imag} */,
  {32'h417e242c, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'h42311295, 32'hc1c96d04} /* (0, 13, 7) {real, imag} */,
  {32'hc21053dd, 32'hc18d9c35} /* (0, 13, 6) {real, imag} */,
  {32'hc2813847, 32'h40bc0ea8} /* (0, 13, 5) {real, imag} */,
  {32'h40add2f9, 32'hc24bc0fa} /* (0, 13, 4) {real, imag} */,
  {32'h412e21e0, 32'hc24eff2d} /* (0, 13, 3) {real, imag} */,
  {32'hc0d8da14, 32'hc25f898b} /* (0, 13, 2) {real, imag} */,
  {32'h42d4c0b0, 32'h430e799e} /* (0, 13, 1) {real, imag} */,
  {32'h4250d7a6, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'h43b61c53, 32'hc282cc06} /* (0, 12, 15) {real, imag} */,
  {32'hc2e4d0b4, 32'h4272563b} /* (0, 12, 14) {real, imag} */,
  {32'h41a358ab, 32'h430d40bc} /* (0, 12, 13) {real, imag} */,
  {32'hc250b8b3, 32'hc09e6e9c} /* (0, 12, 12) {real, imag} */,
  {32'h428ec84d, 32'hc0607938} /* (0, 12, 11) {real, imag} */,
  {32'h423c5873, 32'h4229fcc5} /* (0, 12, 10) {real, imag} */,
  {32'h42905182, 32'h410c4350} /* (0, 12, 9) {real, imag} */,
  {32'hc2b5ac31, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'h42905182, 32'hc10c4350} /* (0, 12, 7) {real, imag} */,
  {32'h423c5873, 32'hc229fcc5} /* (0, 12, 6) {real, imag} */,
  {32'h428ec84d, 32'h40607938} /* (0, 12, 5) {real, imag} */,
  {32'hc250b8b3, 32'h409e6e9c} /* (0, 12, 4) {real, imag} */,
  {32'h41a358ab, 32'hc30d40bc} /* (0, 12, 3) {real, imag} */,
  {32'hc2e4d0b4, 32'hc272563b} /* (0, 12, 2) {real, imag} */,
  {32'h43b61c53, 32'h4282cc06} /* (0, 12, 1) {real, imag} */,
  {32'h421187de, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h429489d9, 32'hc2ca2da3} /* (0, 11, 15) {real, imag} */,
  {32'h425ae24b, 32'h402cd1d0} /* (0, 11, 14) {real, imag} */,
  {32'h4230d70f, 32'hc1acf33d} /* (0, 11, 13) {real, imag} */,
  {32'h40faae41, 32'h41cc7e06} /* (0, 11, 12) {real, imag} */,
  {32'hc13f35c0, 32'h42c785c4} /* (0, 11, 11) {real, imag} */,
  {32'hc02ea31c, 32'h41848a45} /* (0, 11, 10) {real, imag} */,
  {32'hbfcd8e20, 32'hc0f0e500} /* (0, 11, 9) {real, imag} */,
  {32'hc1a02f07, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'hbfcd8e20, 32'h40f0e500} /* (0, 11, 7) {real, imag} */,
  {32'hc02ea31c, 32'hc1848a45} /* (0, 11, 6) {real, imag} */,
  {32'hc13f35c0, 32'hc2c785c4} /* (0, 11, 5) {real, imag} */,
  {32'h40faae41, 32'hc1cc7e06} /* (0, 11, 4) {real, imag} */,
  {32'h4230d70f, 32'h41acf33d} /* (0, 11, 3) {real, imag} */,
  {32'h425ae24b, 32'hc02cd1d0} /* (0, 11, 2) {real, imag} */,
  {32'h429489d9, 32'h42ca2da3} /* (0, 11, 1) {real, imag} */,
  {32'h42d680af, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h41848bec, 32'hc33e27cb} /* (0, 10, 15) {real, imag} */,
  {32'hbe512b00, 32'h42242efa} /* (0, 10, 14) {real, imag} */,
  {32'hc22d12fe, 32'hc2433786} /* (0, 10, 13) {real, imag} */,
  {32'h423fd0b4, 32'hc1d16f8e} /* (0, 10, 12) {real, imag} */,
  {32'h428a10ec, 32'h413e9d84} /* (0, 10, 11) {real, imag} */,
  {32'hc18ce1d8, 32'h429ed5dd} /* (0, 10, 10) {real, imag} */,
  {32'h41fb4aec, 32'hc24c3a36} /* (0, 10, 9) {real, imag} */,
  {32'hc1a4ea96, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'h41fb4aec, 32'h424c3a36} /* (0, 10, 7) {real, imag} */,
  {32'hc18ce1d8, 32'hc29ed5dd} /* (0, 10, 6) {real, imag} */,
  {32'h428a10ec, 32'hc13e9d84} /* (0, 10, 5) {real, imag} */,
  {32'h423fd0b4, 32'h41d16f8e} /* (0, 10, 4) {real, imag} */,
  {32'hc22d12fe, 32'h42433786} /* (0, 10, 3) {real, imag} */,
  {32'hbe512b00, 32'hc2242efa} /* (0, 10, 2) {real, imag} */,
  {32'h41848bec, 32'h433e27cb} /* (0, 10, 1) {real, imag} */,
  {32'h43202c18, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'h42a29d71, 32'hc0b46fd8} /* (0, 9, 15) {real, imag} */,
  {32'hc1f6005d, 32'h42a930a8} /* (0, 9, 14) {real, imag} */,
  {32'h43496c9a, 32'h4173dc44} /* (0, 9, 13) {real, imag} */,
  {32'hc2b5e96a, 32'hc15d7610} /* (0, 9, 12) {real, imag} */,
  {32'h42acad6b, 32'hc26fc3b3} /* (0, 9, 11) {real, imag} */,
  {32'hc25a63bf, 32'h42cbf10c} /* (0, 9, 10) {real, imag} */,
  {32'hc2211ee0, 32'hc214a941} /* (0, 9, 9) {real, imag} */,
  {32'h429473ce, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'hc2211ee0, 32'h4214a941} /* (0, 9, 7) {real, imag} */,
  {32'hc25a63bf, 32'hc2cbf10c} /* (0, 9, 6) {real, imag} */,
  {32'h42acad6b, 32'h426fc3b3} /* (0, 9, 5) {real, imag} */,
  {32'hc2b5e96a, 32'h415d7610} /* (0, 9, 4) {real, imag} */,
  {32'h43496c9a, 32'hc173dc44} /* (0, 9, 3) {real, imag} */,
  {32'hc1f6005d, 32'hc2a930a8} /* (0, 9, 2) {real, imag} */,
  {32'h42a29d71, 32'h40b46fd8} /* (0, 9, 1) {real, imag} */,
  {32'h439ee1d0, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'h434e68ba, 32'hc1bd7762} /* (0, 8, 15) {real, imag} */,
  {32'h407e4620, 32'h42f01e37} /* (0, 8, 14) {real, imag} */,
  {32'h426869ad, 32'h40a40490} /* (0, 8, 13) {real, imag} */,
  {32'hc22809f1, 32'hc2147861} /* (0, 8, 12) {real, imag} */,
  {32'hc24ac2d6, 32'hc1463abc} /* (0, 8, 11) {real, imag} */,
  {32'h401d72e0, 32'hc239c1a4} /* (0, 8, 10) {real, imag} */,
  {32'h42803111, 32'h42afbb3a} /* (0, 8, 9) {real, imag} */,
  {32'h428fbaba, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'h42803111, 32'hc2afbb3a} /* (0, 8, 7) {real, imag} */,
  {32'h401d72e0, 32'h4239c1a4} /* (0, 8, 6) {real, imag} */,
  {32'hc24ac2d6, 32'h41463abc} /* (0, 8, 5) {real, imag} */,
  {32'hc22809f1, 32'h42147861} /* (0, 8, 4) {real, imag} */,
  {32'h426869ad, 32'hc0a40490} /* (0, 8, 3) {real, imag} */,
  {32'h407e4620, 32'hc2f01e37} /* (0, 8, 2) {real, imag} */,
  {32'h434e68ba, 32'h41bd7762} /* (0, 8, 1) {real, imag} */,
  {32'h42b82f9a, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h42d46765, 32'hc2aab120} /* (0, 7, 15) {real, imag} */,
  {32'h42891b90, 32'h43320430} /* (0, 7, 14) {real, imag} */,
  {32'hc04eafa0, 32'hc26a3f89} /* (0, 7, 13) {real, imag} */,
  {32'h40369330, 32'hc144d490} /* (0, 7, 12) {real, imag} */,
  {32'h4240a6ce, 32'h40710670} /* (0, 7, 11) {real, imag} */,
  {32'hc1891776, 32'h419f6696} /* (0, 7, 10) {real, imag} */,
  {32'hc06025a8, 32'hbfcc0e20} /* (0, 7, 9) {real, imag} */,
  {32'h41ce55f1, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'hc06025a8, 32'h3fcc0e20} /* (0, 7, 7) {real, imag} */,
  {32'hc1891776, 32'hc19f6696} /* (0, 7, 6) {real, imag} */,
  {32'h4240a6ce, 32'hc0710670} /* (0, 7, 5) {real, imag} */,
  {32'h40369330, 32'h4144d490} /* (0, 7, 4) {real, imag} */,
  {32'hc04eafa0, 32'h426a3f89} /* (0, 7, 3) {real, imag} */,
  {32'h42891b90, 32'hc3320430} /* (0, 7, 2) {real, imag} */,
  {32'h42d46765, 32'h42aab120} /* (0, 7, 1) {real, imag} */,
  {32'h42a13dea, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'h4229457a, 32'hc33d7b8b} /* (0, 6, 15) {real, imag} */,
  {32'h42faa7d0, 32'h425dfd96} /* (0, 6, 14) {real, imag} */,
  {32'h43122308, 32'h40227b08} /* (0, 6, 13) {real, imag} */,
  {32'h4292903f, 32'h423d5e6d} /* (0, 6, 12) {real, imag} */,
  {32'h42782308, 32'h41c07f56} /* (0, 6, 11) {real, imag} */,
  {32'hc2897bb0, 32'h4178e1b8} /* (0, 6, 10) {real, imag} */,
  {32'hc1e52976, 32'h42179a20} /* (0, 6, 9) {real, imag} */,
  {32'hc2191690, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'hc1e52976, 32'hc2179a20} /* (0, 6, 7) {real, imag} */,
  {32'hc2897bb0, 32'hc178e1b8} /* (0, 6, 6) {real, imag} */,
  {32'h42782308, 32'hc1c07f56} /* (0, 6, 5) {real, imag} */,
  {32'h4292903f, 32'hc23d5e6d} /* (0, 6, 4) {real, imag} */,
  {32'h43122308, 32'hc0227b08} /* (0, 6, 3) {real, imag} */,
  {32'h42faa7d0, 32'hc25dfd96} /* (0, 6, 2) {real, imag} */,
  {32'h4229457a, 32'h433d7b8b} /* (0, 6, 1) {real, imag} */,
  {32'hc30522ac, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hc26c038a, 32'hc2d3199b} /* (0, 5, 15) {real, imag} */,
  {32'h425ca011, 32'h42c6b0be} /* (0, 5, 14) {real, imag} */,
  {32'h428107cc, 32'h4299f753} /* (0, 5, 13) {real, imag} */,
  {32'hc102af14, 32'hc1b94c14} /* (0, 5, 12) {real, imag} */,
  {32'hc11237f0, 32'hc04d02d0} /* (0, 5, 11) {real, imag} */,
  {32'h41ad1cd4, 32'h3fba2990} /* (0, 5, 10) {real, imag} */,
  {32'hc2917ad4, 32'hc295f0be} /* (0, 5, 9) {real, imag} */,
  {32'h42844e7d, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'hc2917ad4, 32'h4295f0be} /* (0, 5, 7) {real, imag} */,
  {32'h41ad1cd4, 32'hbfba2990} /* (0, 5, 6) {real, imag} */,
  {32'hc11237f0, 32'h404d02d0} /* (0, 5, 5) {real, imag} */,
  {32'hc102af14, 32'h41b94c14} /* (0, 5, 4) {real, imag} */,
  {32'h428107cc, 32'hc299f753} /* (0, 5, 3) {real, imag} */,
  {32'h425ca011, 32'hc2c6b0be} /* (0, 5, 2) {real, imag} */,
  {32'hc26c038a, 32'h42d3199b} /* (0, 5, 1) {real, imag} */,
  {32'h426a341e, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'h40c635c0, 32'hc370295d} /* (0, 4, 15) {real, imag} */,
  {32'h429bb9de, 32'h4278dee1} /* (0, 4, 14) {real, imag} */,
  {32'hc285a38f, 32'h418c4000} /* (0, 4, 13) {real, imag} */,
  {32'hc2366031, 32'h41b12c83} /* (0, 4, 12) {real, imag} */,
  {32'hc16c26a6, 32'hc220abf2} /* (0, 4, 11) {real, imag} */,
  {32'hc17c89e5, 32'hc1efe702} /* (0, 4, 10) {real, imag} */,
  {32'hc1f457d1, 32'h429beda8} /* (0, 4, 9) {real, imag} */,
  {32'hc082d370, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'hc1f457d1, 32'hc29beda8} /* (0, 4, 7) {real, imag} */,
  {32'hc17c89e5, 32'h41efe702} /* (0, 4, 6) {real, imag} */,
  {32'hc16c26a6, 32'h4220abf2} /* (0, 4, 5) {real, imag} */,
  {32'hc2366031, 32'hc1b12c83} /* (0, 4, 4) {real, imag} */,
  {32'hc285a38f, 32'hc18c4000} /* (0, 4, 3) {real, imag} */,
  {32'h429bb9de, 32'hc278dee1} /* (0, 4, 2) {real, imag} */,
  {32'h40c635c0, 32'h4370295d} /* (0, 4, 1) {real, imag} */,
  {32'hc250d680, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hc306d315, 32'hc3979851} /* (0, 3, 15) {real, imag} */,
  {32'hbfd28a90, 32'hc280394e} /* (0, 3, 14) {real, imag} */,
  {32'hc32ab064, 32'h4124f680} /* (0, 3, 13) {real, imag} */,
  {32'h418b1b88, 32'hc2ac0345} /* (0, 3, 12) {real, imag} */,
  {32'h407c8a60, 32'h42735c23} /* (0, 3, 11) {real, imag} */,
  {32'hc1a2f2c6, 32'hc1dd3ab7} /* (0, 3, 10) {real, imag} */,
  {32'h4273b7dd, 32'hc2b74e13} /* (0, 3, 9) {real, imag} */,
  {32'hc2c52a60, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h4273b7dd, 32'h42b74e13} /* (0, 3, 7) {real, imag} */,
  {32'hc1a2f2c6, 32'h41dd3ab7} /* (0, 3, 6) {real, imag} */,
  {32'h407c8a60, 32'hc2735c23} /* (0, 3, 5) {real, imag} */,
  {32'h418b1b88, 32'h42ac0345} /* (0, 3, 4) {real, imag} */,
  {32'hc32ab064, 32'hc124f680} /* (0, 3, 3) {real, imag} */,
  {32'hbfd28a90, 32'h4280394e} /* (0, 3, 2) {real, imag} */,
  {32'hc306d315, 32'h43979851} /* (0, 3, 1) {real, imag} */,
  {32'hc2ea4ffd, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hc3573240, 32'hc3720566} /* (0, 2, 15) {real, imag} */,
  {32'hc286d854, 32'h425241e0} /* (0, 2, 14) {real, imag} */,
  {32'hc1dca944, 32'hc2ef77ef} /* (0, 2, 13) {real, imag} */,
  {32'h42c667de, 32'hc0f9a948} /* (0, 2, 12) {real, imag} */,
  {32'hc1fed108, 32'h4333dc78} /* (0, 2, 11) {real, imag} */,
  {32'h41675720, 32'hc2e26d72} /* (0, 2, 10) {real, imag} */,
  {32'h429e30a2, 32'hc271b442} /* (0, 2, 9) {real, imag} */,
  {32'hc2bac722, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'h429e30a2, 32'h4271b442} /* (0, 2, 7) {real, imag} */,
  {32'h41675720, 32'h42e26d72} /* (0, 2, 6) {real, imag} */,
  {32'hc1fed108, 32'hc333dc78} /* (0, 2, 5) {real, imag} */,
  {32'h42c667de, 32'h40f9a948} /* (0, 2, 4) {real, imag} */,
  {32'hc1dca944, 32'h42ef77ef} /* (0, 2, 3) {real, imag} */,
  {32'hc286d854, 32'hc25241e0} /* (0, 2, 2) {real, imag} */,
  {32'hc3573240, 32'h43720566} /* (0, 2, 1) {real, imag} */,
  {32'hc204622b, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hc30e2ac6, 32'hc314ac39} /* (0, 1, 15) {real, imag} */,
  {32'hc21add0a, 32'hc21c02d1} /* (0, 1, 14) {real, imag} */,
  {32'h4247babf, 32'h42602f0d} /* (0, 1, 13) {real, imag} */,
  {32'h42f149d6, 32'h42f9e655} /* (0, 1, 12) {real, imag} */,
  {32'h427fa27c, 32'hc27ca9d3} /* (0, 1, 11) {real, imag} */,
  {32'hc1dc4f34, 32'h42ada766} /* (0, 1, 10) {real, imag} */,
  {32'h42237893, 32'h4187779c} /* (0, 1, 9) {real, imag} */,
  {32'hc23bfcb9, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'h42237893, 32'hc187779c} /* (0, 1, 7) {real, imag} */,
  {32'hc1dc4f34, 32'hc2ada766} /* (0, 1, 6) {real, imag} */,
  {32'h427fa27c, 32'h427ca9d3} /* (0, 1, 5) {real, imag} */,
  {32'h42f149d6, 32'hc2f9e655} /* (0, 1, 4) {real, imag} */,
  {32'h4247babf, 32'hc2602f0d} /* (0, 1, 3) {real, imag} */,
  {32'hc21add0a, 32'h421c02d1} /* (0, 1, 2) {real, imag} */,
  {32'hc30e2ac6, 32'h4314ac39} /* (0, 1, 1) {real, imag} */,
  {32'hc31982b9, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hc1d74bcc, 32'hc3140479} /* (0, 0, 15) {real, imag} */,
  {32'hc2b9b9e0, 32'h41174568} /* (0, 0, 14) {real, imag} */,
  {32'hc0a2dea0, 32'h430122c2} /* (0, 0, 13) {real, imag} */,
  {32'h424f8caf, 32'hc1d3a003} /* (0, 0, 12) {real, imag} */,
  {32'h40c30ebc, 32'h41939b98} /* (0, 0, 11) {real, imag} */,
  {32'h423a8cfc, 32'hc20c9238} /* (0, 0, 10) {real, imag} */,
  {32'h4187615c, 32'h42143420} /* (0, 0, 9) {real, imag} */,
  {32'h428e78dc, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h4187615c, 32'hc2143420} /* (0, 0, 7) {real, imag} */,
  {32'h423a8cfc, 32'h420c9238} /* (0, 0, 6) {real, imag} */,
  {32'h40c30ebc, 32'hc1939b98} /* (0, 0, 5) {real, imag} */,
  {32'h424f8caf, 32'h41d3a003} /* (0, 0, 4) {real, imag} */,
  {32'hc0a2dea0, 32'hc30122c2} /* (0, 0, 3) {real, imag} */,
  {32'hc2b9b9e0, 32'hc1174568} /* (0, 0, 2) {real, imag} */,
  {32'hc1d74bcc, 32'h43140479} /* (0, 0, 1) {real, imag} */,
  {32'hc3676cd7, 32'h00000000} /* (0, 0, 0) {real, imag} */};
