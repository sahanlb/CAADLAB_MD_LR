-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
KXqfdT4fFLgZcMT3YRzT30A7M27CDzzoGnyKpkVPGScr2P0RDMO838JVgwecHuCC
rBw6Pm7rLouVlw+/uGnj/UI20RFXwX5iOyRc5PZVIgtpYEAOArU+Da/s1vKqyzNx
BcGdLMkPMy2/J47gP1fEvXxwbTFth1R5crY0y8f4pXw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8848)
`protect data_block
3lW0B8hBodMYHjwmp/RrGGUerAvyIBbBRMq0oOA5mG/ZMEMJRlBH04sIzddL+8j+
85ZxGwuKclvu8nX8gNar2IEd5A+1A/Ebpuqi2Ekfo7wpbspZlqdWSVjnFQwStYjs
uOGNfOGcyd+0WVkUFOw++qYVZztRPez0k1BL0FJap/4MYXAbQsfq30A53lvuPzos
M1qK/EMmVPUQpzjt7ksWDQr1USBnpALWLAgnh55fb+uibG6PKR5xQSIofAKKeJ7Z
KcRavtMgGUyjGH1vajRcjJdVglEHaaYlJMfPU7NmETxkAvgLL3g08sWCXezgKXpQ
OlVRhKXYJJh2zx4zjlSgj/TKz4pvLnYGXRbJJbQF1J+a5zO+vBWuxMwU2O7lJF8s
hfoVJrMyAy0GhbunSpo1tAlu2+ukHgGChqztG1Jh/96KZ84Fq2U0sGgjov4OnB6y
kfTjAb8fDJD5mEA1FsVamIcXcr+/wM/Wg11cAO03nsxtsv5CryTC+Iv9PzBCZRTp
vUNNhxuZpcQru9XXZZrf8U3nstGITXefK2jmkQ06Zyl0i8/MXGekPTZu49uIMfMA
6BBI4md9rtIyQEZmMc+Y5H+M371MRlR9vBRd0QZL4aCKHvBTw/e+vrqZhr4/ehiE
B02Z0t4A1QVSFPJtCCm1WHAGKvD/c95mAjyx23/XaBnygL+K7opNt/1X4HF4Zat3
0YmowYdY1LB4smr01TyPBPrbAyJZKN995MYI6AKBq+pghlh1fi7nB9bJbhfE5cNV
xmUjs8TROKtZCuvQjY3d0z0paxSR0qskwj6D9E0Zch3B8OAzTxshm9JA043bENyr
scLS3EQCyOpKA5Ae0cFPht4lncEe9uryQS9tVMGH9Fo5izJFN1RAzUCvl1blzqgN
+yv+Wgq/dGrFQc/OoTBvdhlZ5PGqTu/bafahvhaKrEofcjFnuv3HeuQdtNxB2vXR
Yy7hp7KRkThJW2TSbB+hfRW3JPhzhOyzMJlKjgQ9dzGjdT0y+RJNQHDvmHx1Ie9t
sLEeafXjGuHKyBSvhqDgMkfYCZKJvcflAmAYh5tgNDls3hj1CQbdF9GC7SC+LyyP
CsOS6FnHpl0e7SMvO2fnMdr2PhIW28Q/HC2Bh/+o1OiXvAq6apOofx1U1EUTo8ph
0rkdsCBQi8WSPCTntZ4j8GNCRAGE9wQOfEKrjdCjMIKOr4grFt5YS088XlAxAyko
8vSD/sVPJi4Ey2c/iz3zqbSI8f6ip7adWdai9k5aKoiK3I+O87LM5SO7O53N6AUS
U+mP1AaWIwf0iVCtWcP4Y9A2rDXzTaLJMVK+rGyzd9bSvEDY8C5sg4Q3Se4msd4D
Q9rfjOCHvTTU1Ox21vnzPejTu3LGg0tzKfBeKoaanuSspDNDdhN5Ko2SkPcpzUpB
eYneXmwcmDNp6PVYcrq8vsQE/APFGR4dqpLwWQB87UGD/mTCoDUBEytQnDudtGt8
7J8Zuq0YECdqYHZ+Y72a7PkxKfmS1SCNxAubWYJzQcSU4Uj4pZSk57TCUY61jKsr
RhET8RyxnH/lYEbZCW5uttUUpmJXG/bymv3dfPTWmWt0zprBuCNRjSXHR3SkKgGC
u/khCV7AJ194PNnO+PIyqLA5SJmot7UIwcSvTrwD/I771ZHhPIc8X0rML8OhRvV0
L6n3kjvnX7d3WqAd9v4NW6NReJsxy/VYa05h6I86MCKShi+Se+QWAYBjPU2p6Wuf
l+KwW8nKZpWb1Bj9MRcv1OXYyenG3n3dzMwzPDJedbxXZr3O7lhM2+pj7mhPhbkC
nwZjzajfcwuzyfCfJSuEnk0cho4dSMaSjEUvSm68gMYf297vRF6AQie+2qno9JwP
Un+4W58YvwV+4IHN1HvYYmCMGz5xPm/IPP80P0GfcfsJIPnIuuV74HhxBdZUCIwh
JvgjL4qIrB2RkHAMWrgKamgMmRYVx3Lul7EX2vPMIcNQevzBIj1qpxSr0fE4i9uf
yZNR9Dv9lCk4pM1VNaOj7IcPmH83iIzKodU2jmDkmCduM+DRivpNQIVXX1ac1J9o
rPlleeiD++/B9ib9xP2KieoezRRdCro9diDXPPiiKuZV8C/Yu9Bz1dXMHtNUgjwB
sQS9CruqZa258Pkz+KTJv+itzWR216ii2nNGQMPPyLr1l3bl0EDRzmjqtdzIPOGi
MYP4Yz3SdOKKDoulqjvU8JG9JSBiXSCDWbouh14QYh+CtCp95hKVZeYNWI+9HsCo
BRpFqI1ebj5QAcOUPD3Q6BZCx7dmLT6yNBoWdRBUoATuMThWNeM8EqGV+hOmSqu3
q9JOYW0oInkBNXQ27pwZtf28/JISd0d2wxyC2AwW7ig2UUmQ3csEPO1WyfQteIeP
psVjlgjH8Z1Rg1GKk1nu3T7rGwMTuvm68PYjuhErQzdWJnq/J0e5EcOjv6ke5qwp
vyxwOu0SUjkjoEbTRGmraQMWBdrVuYqMGY3quPR017Yd9SQUGJWylgdqt/5b0Oox
TEOtYUfXZWXQwnNW4pcx4UHSfOy7KsPqXWmIOJQEW1nMXuNNXFk5+cktB7DrEJaL
q55crKqDUDGxLgHZR8kUh1+fpkuB0BEEcBXW82vu9eertm5DtfsgyACkrglmXOzC
pQ6aJFYs5FRgL1vKN6s6RTU186dDFRBdNCzvoXPwLL6FXjrLo53td/3SmH0BALqc
JABoSkkvwgwDIA3rt3Fd/HkNxaCe8VjqHnydMV7zmFfIDiMvcWN1iDWJpVsQ26GV
tlWV8/wY7A50Py9mzsADckLrXUZ8v1ZLVMbMnAM9YdxwBfHIDBds8cBrrSvLg9GN
xwrCKI6j/yD2suiJjQSftHyPBSM0KyB33scBCOOmhvcr+Om+107eMK/AnXacKowx
yGieTtFY3dY6J6TAuLLF7zvzjqVaCDJlJpzJAK4zqzvZnRzMeEZP5rYmwTrE0TvA
PQaSuJaWloV4P9D0onWLTFMuaswxjCvY2y61RNEsY3LUchwWZa8QRWZFepacGFnl
hHTP4e9UEuYsymyWA/Jir5Hor5+2aFHHU+V8IjHBM9LD+etYNdw1SRPpmh8lnH9d
qjPzCcZr5rtTu4q74E4JlRNWoj8PyMIl6VlvAKIozkQNWRAShWhpbns/e/RE04pF
UWxXoBkiGEdznL8A9QG4jn+KNHlXq6yd93IXXk+DlHWMnUJC1DLBImcgw5CDpBs0
tgtVLXLuogA5/B667VEYeMjynuZLDBw5RQN8xbgVFmzUmr91ttW8BpqGiBzchfsW
I875kS6n5P9AJPkbyQpwiIkD/N/fUjXFm8At8AArvQkv8o4DAG/0h8xI012pj044
h99Y1asVrfZvsYpNuqc1RvXjaxjSoOJejRXkrGYISXgBDVtXba8KI6nvf/CB1+d/
SW1noChKxcTmODv1zC3fQ8CP/FbkaYcsBipwTyN79KUg1mLJ5tkgRCM265hZxesx
04u0m834FgnlLo5fjVOW9lEIKl7RkRufxY4Xv9/kvbTBpYz63+I1KOHy2k9O92eg
bXbVF7gihdggrIT/yTJEmQOxEDRPLzZ6py5MOsVQvf/QMk+ZAuCJi7MAmHitwaRC
fl+t4yGttBi9yaXShwooZdWo8b71AD01HtT2DAauu5/ZYA1V+XRsJLq8LeN3splz
hUizljW+whVna3bTEdscNlYEsJt+1v4RbQq1N6m5wfVCjPsIfYEn5UIUHJqCdPem
MUnteGb79PLC5+QFZplkmyUB/ewW+vGYD/ljRvw1L30FSeLsKqllom/jaCn3uWXH
gZ+8qIZRdcl53mUpt+Oymri0j5ksl6Wuc4tnQ5BVyyrIWxYmKkk8yzsBHboLoEYC
zHVbnLCNP8rBOqsNsmV+nDtZ2UF+RxLT2l54rs9NmDDQfpxoRPYm2NiR8KoFFuHw
ZgtHt70pV8zBGaWW1S6tf1P2Ggd4e6ClSCp8U9cVm1izUKbLVQ+X9EXLP82XXbTM
QMwjNO7NFyRBSHfxXbYW5HKB/xsudvTQSu0yeohWLg2JeIxEFsQV7WlSMHa3Wxzd
kOjxxZoO2EXbSy4wQ9wGISIoqkbhsas757QKkhQMN4Mzjo7K95TQ1kZsp0OVPo60
fd1s2zAqAnXT+BgweSElLkn5R/9IswQ7YZ0ISnx1HTTjTrmaDsajMPy3Tik8Dgbd
DAbjccAwIQudAYzyL5nNp2IR8YgS/RXVZTh6TR5mJYj1ZnYfr6gRHn55uFutqiVc
AsZHnxMeUreOGyiVZ3D240pLgwAtbJvWhz0o9k0xjCpzSZAfdXxNIlJ8jrAX+b3N
4Xrpo+KiclrMKrZ91BISm+VDwIhhBJ1Z0Ntongcff15R2NV9KpY539PcuAZO0V8h
JvS7TKKOIwMyp3TzY6QGNbET93VQ9XmqUhgHSZOLkz+WunMWvwspLKWPx0PWRxzp
HubgcY+UzVedvIy78LfSaGEi77myMMrkcC+uK99rtGOwFpN3IDjPB13WRQ3br0ed
4sGAI6cAkfLm8Ihf5OOqJKcdHE4CQ33TAPVCnm+HCCsGjFV22ixwT0sLaxm5aET6
hH41eolV5ap1TRceipgCcgvfFNT8pC+DPE9qT2Yl05I1UUseOo5Oz9L08krslIZU
lFAWabk7hXrsaWRxCsH7IvLOFnVr3qSgFcZhXZmYUwmDH1Y89vL7Jhn2DP9kR1yH
qOHEmCpau+CQFnk1V6JHUJPikVLHMsV/PT6q/7dB2u71gsfFkdMMwR++/d3yOGxf
JRTqzwWh0GiyV8h3QaDWzlqmNTNbKvV3Eb5C5RidmTYfgSVAVjXEyYDp2GiXTxaM
lIKrU6kBVmJK1iOHXn2kYNCGVOI1Y0O6N/PKeiqVLu9bUaYxwIkm235dESxVPag+
vraIZGjt9A27QhCtaof6ELrOuzqoxQYMcLOT6jfb+6BT/kHE/CzJ3MtxEij4W18I
HT8NzSv/6PFya/0xA7emRZg9f0TsAWyPHrA2U8Txamjm0Oaf6VFKiLO41ayD/WJG
or7QZbGMDeLXI6VaxkaLPOQEv+8KqfsfL3+M3mIv7ANVSY6+pVNxgjIq8kHjh+A+
zoSqHW9CprgZww0WwECEqoGPJrV7f8hp382zHkX1x9sRgDZ+FHLmmGOnYpiZi+Z4
rISHWHdMNCQzUDeFBfCmkBFNE+DPl+3fD4+RtVsxWJ6AKH6qTQntn9S97vbwiVAp
Zj2V4r9xKULJmMNdFY+S41lcGIc7oDC7tJrbTkgDG0cDorINfTSxTMit0h34OTkA
Sl9qs2TUCC8oIMElSHm7fMd6++WfwjUKhNAu6BH3o01mdiCrXRPjKJgosxW9PJgL
R1L5yHRJydJjKgg5nToDqJmjLxp3PLelA9/kWs0FScuX+0Vee06mmuMtq5i/hqCK
fhaeEJGj87oKHAZVrTWhrPck1sn1iAMksr6ykqfNHWUtlZ+uL4tLJnQZ70wKHsyM
ITErhMoTx4t529t8saRpI+QSlwmR5Q4vHH+cwkILmlsFycDqiY+tgARzo8UAClAW
Ag9D33KHy/Dglv/8iTEDxEexDhgshIGolQcljLaTWm/i6w/EzgvK/RxztBHJEmZN
+k5CWNQJbv5Q1HvM/WV1kWXMX86pkv/oWkuFiQNqut08uNxIXiy6TZ+qenwQcwxY
Y5yE0Mvn4IiVscUl+B8iGrVgdw/mSa84HWOXg2W2gcxfO42LCaONqmWdD65cicQB
iNZyB5SZR0SxYg12nGSkbqb4Qgha3gDd2LLG1qTUHkke7lIspJCZxVWyvzvHLWSV
56+BbZEge3jcSefuTy1KMn4Pw5kp7hfquUAE+jFv8QltJgM7xL4jrjtiaJUvlvzA
MrODVyKua9WOCnIfzGpSN6ar3Oa5Ij/06vEmXNTNg1x7hycH8SN1DiuWPXyVSrjw
bCxZY0CS7eZeYe2jBwm8lZPUj27WXcDzlmaUVqrjISJIxs2JqW7pDxN3fP4U1A8E
K+8fYwWYEovvVeXqHLGloeN7f1DaiDMuvsaxBpUhd81epkJzeXw6DYFX/GbXNgtt
9Wl8JDI1lIXUp9rANGj1a/apF8uHkDkIwlIMJTqalATb7/TEebzqVfsl8ABnG1C0
kG04gs8xsFkBAMcQt/Zjk5EjSPi5vqmK8Y1q9xFzi4VZeaHrlgPeRnH5dWTqEln7
Uep9t21k/Z5A7qvl3X8k4f+EulODnn+OBQbAQu7fYlvDaOfCt7LpwE5QhV5o3E/3
iR08OIDjGbIBtp/ccd3r3Ox94cAWph0vyV0tjWuPkzoFvczrRVCH6awKN7PXZ7nd
n2fD4kysvv6NPesUeRH1RiGGNZFZdEGFgW3/7pVYz9Gf8+UU/ZVwiNvCXCdeS03h
Zvq0NEmAWCekd0U8rUaBXQ2AzSP25VYuZiD06rSXEiGNCg2EIMNEKiB1xbyVXY7T
G39kOlfsEl9NsP0E6crBk7nqVTR3rKhGSB3OAjBn+BAW+gMR1XAW8g/Ti+wBG3ib
iDBUrhUatz/a/x/gJP61TU0kUic9QJ7ZW+rJglwWKJ4sW5Y8SDOkKzb9iFSArg67
m5kyFA3pz6dTyPXPlDcPe0qZKElj/Mq2OLZmrV3hJDcUeBB8vozgOdcModOE2Yff
zfN2iD2ljUziETLRS4DICJANrCn+un1UBMYVpK1sWtj3s7BAmSaSPUTaEL8K4Aoq
Z94MTjX9u4O2L5TQXQESSrIhcqLsyWs2HDiXk/BxkruXEM0F9yqP1j3eIgVnGDJ3
X/oHtswVAzMosjPIRIndCrqaM8mV5mrpkRHQfeKv2h826vBv7xpeUe+GMK/D3Fht
FpkglbBJNmiyLR4wtVeywFQsS4fFxjaQ/V/Let3lFSsWveWgoffiDjHoI5tAA7Re
YZRC4jvYLmhoVIrCPgJRtEdbcbsr3hwjFV2AL8uMbW3J4qo+WzIe64u6qqob/LuW
pNrX/cLKqRW6WWtb16LJ8QPqoNYsKmE02Pm0fvVp/fz9uM1MCLrqdsM3DMbpy99I
gYFR7zpr4aAbOiCXMocUY4Umr9A4XHyjQJaQuTRDT9pFjCDFc8sv6LEuqyXvRFEM
PKkHkDPBjSmXxN4IeLeSVgwjoQHC9rNtqfP/Z5i9d/Vo8inA+/FUMa6XS3p922hr
GTmsuSSLioYeYFjydYB4uTysms71IMEbPJTB+JvVRTK8uFNTQYNFU01jTv7erqzZ
MArGva2UvX4BuOMQ+Loo/6lipLfAOthPUw7veh5/a2/uDimt/rp7cy6i29gabpdw
kFKyqf9g9xglaBPJ2wOsENaqZFJWNr/6mIDEEpN4XHL/Ow1oA7ki4BOngwEI4zRQ
TOhnf6vcjqDAOxqv3V86NYUqC/ljZdfVmQQH2+RMOlA0mpGOiwfyEgFTuVSFnZJu
vN55WyM3PnvvvYeHLVsZGEAL/8FdjuXuUk7RPP6yTQBe2W3WoSl7Siqbo8lc1oPD
TZyRmg2ea1c74Z2JztlIeMlQxCEJnnIHR35PQLBCoM/ZZMky7+ZG1V6IUCPyLU0j
788ACgoHJZ2HfaKHf6+av0k0mW16Xvgxggd21jWlJN/xytv4NI8YfwT+EiX1tMHI
YvuRhmzbiVf2FU5L/D9QSk09H5d2GrJ98A4bBHbysDoH5t0fq4lMMa3FrVumX8kN
AjXcTpOaKIFGfMChHqfMxLfXBvEjwXcjJecQdavECJkPLG5ASSY8mUc1CM8eSkeO
BX2A95b/dRuBDAFedkKPSKIgLC8Hp3bQKKAM+l7x/0USBZPd/2fFycqbGJv7fZWH
hHSLrOwH/XcuS9uxr7uXc2QN2pDixLxJV2U3BB15jPeqgCpJs83GVEB4XUJHjHKm
OzGZR8oXPC7fMgDolpW6Ky0EhKBe+/SnhqbdfbPObL4PR4ZCo3JVOprvaVtkjsT7
xJMAxTcwUD5lyhzwk6UulPtfrL4yIVg5ABHn2Nw7HmaP0UNbjPXmkWo1/DUP/6b/
c6gZq/OBGBf3wfSLabt9o89yinr9ex5kvLmjxnc1G6EY90vmDFlsECbyg96naRk4
aLBv0hhlNE5bA4Vhxly8IWrqWwwkbFgys6dCioEvXuUG+ujeTR1ZSkfOzDHVUoGR
GLSvmvBTt0VJPZLSWwS+ewF9Y6wa+2uG8eMvKgyEw34JpQpwHa4flDX+VXUc0k8P
KFkexz2fVUMvS10SJDS81Su14ws0yolOvcTAEw0kJUqH4phoM5jjIfu3fklWPlhj
OvEyEjQ1IWLCaBggkgLBXe1GUCwst00zUGuAt3mKO0IumoKa2pNMXCRVQpaX3sW1
j72craAzZUrgBkE8ECkaI0+LlyKTNSaPGL3z3IlJcLkgHLC8SExuOBv41B0PQa1i
3aeJ5Rfabb3zHrbCSivicL+PHBCw3L8kn7gApHT12hNuHdhhGad0GBiz+2be38rP
9iWEu7o6oDDUsux6UXOWeqWcDh6nLrxWjK6DgZMkpusRVenkwQ7COEo1gHQuLsPO
IjWjuOpj06aYhbuD38vtAifjx86sMlFnHrtG+3Za1hfr6sLEZjpZF53Uvm0DlP9R
P2teMxY//cxy/aIPKRe3hiZBEv9M3p7R77MWNedAbNFJ9yPoGmw93ge6fKV8EVei
FM74IMoAb+6bsXJQZhY+GaF89pG8FZXO3DFXa/ef9OedyTKdH/QM4Y2tWk2YhkCx
/8InOU28oRJtvQ0SJ/6f1Sf42Rcni0iHPdMOU7pU8Fv0jz3qbkYyduEiAWRWDw8+
cVMnj1ItYBROrVW+LcUFZYJzm2U4GbJYF2L0NgdrtNec5lc+V5H7Qu9QvqKMlfxN
SKin7oU59JCXea9rFgPfpMMM+dOpbWsah0p4F5i7ayXhF6M/0MLIZlIHmuRqF5M9
V23t+SCtQgP9MBp+syUCWu+2py7ZgtNsHvYrvGPH2p0Zp+hjZ5/XzUWYqfWsiGtu
27FWT9OShAIQuvOEBvcRUNBNj7TktnPmG0GZLSaSC+J5/esTUS33iyR5B/fjUoJu
X/ZCKGB7KWR2DWv76/6kIUAKqXYHRiQKIt3XeJWJnRBRvWrvROhKahlqd1/yr9mJ
ClRMZ5UcSCcJapEsynWF+10kYWRrR63VrJ+CkWNK1/S3YMGnqDRQ3jEeUrhqggSc
ajwSFxDs+mz6RkEFvVroDit/4NiU0g4sNp0dNVs1+nKH/03HHwjIyDbn0GlYlqvy
awAbTtZew2HO8RqhD/QtuoFg1qfkk50+08rNQcbO0J4n1ONQoJ32MwD42lAeB/BX
JvDWtDcgk/rpeEXsH4qiAfZv1kzoy16rpBB0L0YbMe4YMTTfRr6WNgq8gzUY6ZiJ
D3jodGb9/9POW9qnqLqdn1K9xxGb5putWzkv0qqniJ7vsXayFolZ4PGs2qLf/PVx
UKm9ujfBufMxkWv9ChEcbOnl5Tb3l/okcXUCfv2WgMgX44cYjX1SJ0CmBuqr2xRg
G5KAZGGHySUDcJtqQ5TKfb3pTDmKk6rUI9bc3JCN8qhEwdUQ9DRXkqKi0krQlJWY
piKxHHJCVZls7soe19xE0HyBXObyyel29K2dOehOruESwqAgLXgMZS5qjhwFwB76
wc5DiiWvVkYEOsy+x1hA8JO4XMRPVLf+D/aiyZu7+Q2U2DilYSgXYOldqKP0hBdb
6NSmZqOtErz9/vd2jZMbztKnqQ700CQO0MTx7a+yxYXGT170J3IABHR79e18qYWT
ekSgm54fKOFBUZxjl8HNytXaPP9s6kkhSlBaIrt6hT9zhE67h98pYcHZzPb92+uU
zTPjZc8xIcaY7C7yL6LK7xqakR7i7/w/bdz/CCzx96qRsTovn2BmpUqJfunrp3Sj
bkWIeud46L+9vYfpIYfeP40a8pbhiacNMZd8gl1VDm8/9qCy+EujH8HnSEgww5le
v0F1MqFHNVTYQGW54+zLTStCEIWgmo7u2T4IG1wOmPP59DBMInGHdcdkAyZfC+3S
oG2TrrKQnXEp5n5VUwuByDYoMQw6i77hgNATBiMaJUTB4JwRNb8D0O866/9+0SYm
bvQ0+MGmORgxXfI9+36X6jfNxvAixXKUbDPmbqSdj6oJa2bPlksTMQjqcRNxyigp
BUqAkfVBIByVTNBB8ryShDvALoZT1WYP6fm7hI1nGg0XeYMC84k6jF2X86P8DI0x
8dN1itg3g2G8u7eCIai2K6ltw010BbxVYVhpmwbZyLyPDDD2Q63UNjKS3WSEE3II
wZW64DfhCrAIgvUrYPo0t9XwRoDscqK62YJMjqlRMfKcK5KaYW9qWE3nq52XOVdJ
G8Onf8CHJ1CXPG1PH71ohrxblGxpcl7SWdNIFzEYOsTxHeNlkUKEl+HI6SQ+aDxV
cGZSCELfvNIsZbfpQZCyToZVamN1ShfnkUqn7eE6AYBSenmcy9Q+DNCM8eUfTPMB
T9kO4HrcCUZg9EROu8jaUwGSniR6usVddgas7QbitfpRFhj/9gsvHRSUy8qh8lXv
uQfviiBGW3iDnUMreOjiyUD2oVXIkAhHJLSrR3Fq0UANXNF//MaFVzPmrh/QL1qV
mY3t9cb23s1UTZHg0rqm2Tq8d+CSKw6TLmTtWNJCqdCaE43xw+JQdiIu+EXK4nqF
DCkJbzzXx9uKUtVJTipOeA7vYGKxIPmmiBckSvfo5uSgPIXXN/4+Focsx8dWpcRS
bLlcumOFMXV2VPPiN/OeOrJp6M9Y2NBFbeOb3Pr8/RtLp9kJ6cGRkPkMAvN2ie7o
4Woi1jD4C+DlR/aOZk1Q4gwK5gi58TDrxZzdb0rtoNEPjMF0/dTRrL9OnAisDPFT
q/ANFdzSGKEbbI7mq9L954Z4Qt0Ou8dfKhCYgjMS7lu74jQdq/SHG9a56jjxhqjL
a8ANgFjY7/cpD3QWBdWCGVxxFRvA6HWaafO2vU3fs9FNbDWxYZSdrB5Bu2zXbEOS
nLQXqKfvevOc5d9Qpreo1+1XLC5j6YZ2HNaI4Ak8wkeOXp3MUYxHRAP8tO+IQ79W
wwsvisBQWqYmG+8vK1NcAjGFLAtoKaur0lpwyyu3bDmMCsg2okiDgR+nB5LilEzi
WbrMhTClzwVzOoRy4Jgd3p1AwNU3U/kehbDUtYwwStMyK0oaZEYJWdYM39m4wpfR
dUOAaMEt7ETi2D6JIe3c8fswVohQa8t86cc9lnauiJVbSFQebskwmAlsKuHu8IjF
lGcqRhbcGy7MMvT8xF41c7L8IgjUmiV2FcJyf9JMkwg+hDWhFMfp2hhsMX38oSlL
TUm3lmipi+A9zAUvvgxOky/FXZ4eU6de/pwnsskwH2sVcUeegKRykAFUJUgGZNcH
odtg+0Ud6KOPDFXjnF4sh7KzbGvsbAkWrZHoa5rnFej2pPE8lqrtJQHowLP73ukt
2Tqu1ZU7MUhjDfRS7KS+tsqJcVhNAFfLavzg8WwOLbTkQEybD1ud83Q/rp5OcWpW
Z0IZ9fdCbpgKrgnOUH/6tfqR5olqTv4shCwcoyR7o/NZAR3aqdAH1wqws4Tv9nQB
ctd/hQikX+/CQbw4VVB1D0qo95nbZkDY6Vb7mdejn4h4cbkojD+2IKEu+0xpntnZ
tpGTVcZ0lGvVIaaNTJKfjzOt0PjYiHfXFAtxR5DAzr/ipgpWwUCMZG7iTj2ADPzg
Ten3fto2G5DFtj/8m6RpXYV99MqevKfo4ELDd3RAoUn9DaAEwDvBcLiwIAky0PoM
BJLi3uAHqYjTti/J7dmEigyigtNsHce9Rk9dguZM9jHqcVJE9ZIaiDA1pluwjd6M
ZGK+drBhWS8Ds7C+7SC8TLhCQRKl0GNLQGba0XmVYjf7nVLP2I3ZWepw5esNFde1
a+Hk0TrwB56gSY14t2F0fw==
`protect end_protected
