localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_CMAP_CHK = {
  {32'h3de324fb, 32'h00000000} /* (31, 31, 31) {real, imag} */,
  {32'h3e64c377, 32'h00000000} /* (31, 31, 30) {real, imag} */,
  {32'h3e25f3c1, 32'h00000000} /* (31, 31, 29) {real, imag} */,
  {32'h3e4c2c35, 32'h00000000} /* (31, 31, 28) {real, imag} */,
  {32'h3ed2d001, 32'h00000000} /* (31, 31, 27) {real, imag} */,
  {32'h3e80ed6b, 32'h00000000} /* (31, 31, 26) {real, imag} */,
  {32'h3f169433, 32'h00000000} /* (31, 31, 25) {real, imag} */,
  {32'h3ec6190f, 32'h00000000} /* (31, 31, 24) {real, imag} */,
  {32'h3e71d711, 32'h00000000} /* (31, 31, 23) {real, imag} */,
  {32'h3e6494a8, 32'h00000000} /* (31, 31, 22) {real, imag} */,
  {32'h3eac3175, 32'h00000000} /* (31, 31, 21) {real, imag} */,
  {32'hbde1143d, 32'h00000000} /* (31, 31, 20) {real, imag} */,
  {32'hbe7419f8, 32'h00000000} /* (31, 31, 19) {real, imag} */,
  {32'hbe78ef4e, 32'h00000000} /* (31, 31, 18) {real, imag} */,
  {32'hbe48071e, 32'h00000000} /* (31, 31, 17) {real, imag} */,
  {32'hbdd5b7b6, 32'h00000000} /* (31, 31, 16) {real, imag} */,
  {32'hbebd8207, 32'h00000000} /* (31, 31, 15) {real, imag} */,
  {32'hbf0badcd, 32'h00000000} /* (31, 31, 14) {real, imag} */,
  {32'hbeafca96, 32'h00000000} /* (31, 31, 13) {real, imag} */,
  {32'hbe45f263, 32'h00000000} /* (31, 31, 12) {real, imag} */,
  {32'hbdee4358, 32'h00000000} /* (31, 31, 11) {real, imag} */,
  {32'h3ce18155, 32'h00000000} /* (31, 31, 10) {real, imag} */,
  {32'h3ec8e997, 32'h00000000} /* (31, 31, 9) {real, imag} */,
  {32'h3ef798a5, 32'h00000000} /* (31, 31, 8) {real, imag} */,
  {32'h3e80796e, 32'h00000000} /* (31, 31, 7) {real, imag} */,
  {32'h3e1aec3a, 32'h00000000} /* (31, 31, 6) {real, imag} */,
  {32'h3eb8588a, 32'h00000000} /* (31, 31, 5) {real, imag} */,
  {32'h3e91f046, 32'h00000000} /* (31, 31, 4) {real, imag} */,
  {32'h3e1343a2, 32'h00000000} /* (31, 31, 3) {real, imag} */,
  {32'h3ea5413d, 32'h00000000} /* (31, 31, 2) {real, imag} */,
  {32'h3e0c1112, 32'h00000000} /* (31, 31, 1) {real, imag} */,
  {32'h3dc38a7c, 32'h00000000} /* (31, 31, 0) {real, imag} */,
  {32'h3e0d09ef, 32'h00000000} /* (31, 30, 31) {real, imag} */,
  {32'h3e4c4680, 32'h00000000} /* (31, 30, 30) {real, imag} */,
  {32'h3e14946e, 32'h00000000} /* (31, 30, 29) {real, imag} */,
  {32'h3e81e14d, 32'h00000000} /* (31, 30, 28) {real, imag} */,
  {32'h3f0c1ea8, 32'h00000000} /* (31, 30, 27) {real, imag} */,
  {32'h3ecf6c9e, 32'h00000000} /* (31, 30, 26) {real, imag} */,
  {32'h3f48e22e, 32'h00000000} /* (31, 30, 25) {real, imag} */,
  {32'h3f260ecf, 32'h00000000} /* (31, 30, 24) {real, imag} */,
  {32'h3f1425b0, 32'h00000000} /* (31, 30, 23) {real, imag} */,
  {32'h3f22a0a5, 32'h00000000} /* (31, 30, 22) {real, imag} */,
  {32'h3f35d295, 32'h00000000} /* (31, 30, 21) {real, imag} */,
  {32'h3d9949a0, 32'h00000000} /* (31, 30, 20) {real, imag} */,
  {32'hbf07fe24, 32'h00000000} /* (31, 30, 19) {real, imag} */,
  {32'hbf3004c2, 32'h00000000} /* (31, 30, 18) {real, imag} */,
  {32'hbf023029, 32'h00000000} /* (31, 30, 17) {real, imag} */,
  {32'hbed275cc, 32'h00000000} /* (31, 30, 16) {real, imag} */,
  {32'hbf719e8c, 32'h00000000} /* (31, 30, 15) {real, imag} */,
  {32'hbf70e038, 32'h00000000} /* (31, 30, 14) {real, imag} */,
  {32'hbf60171b, 32'h00000000} /* (31, 30, 13) {real, imag} */,
  {32'hbf1da4b7, 32'h00000000} /* (31, 30, 12) {real, imag} */,
  {32'hbed5022f, 32'h00000000} /* (31, 30, 11) {real, imag} */,
  {32'hbe58a8a2, 32'h00000000} /* (31, 30, 10) {real, imag} */,
  {32'h3ea4311b, 32'h00000000} /* (31, 30, 9) {real, imag} */,
  {32'h3f0468fd, 32'h00000000} /* (31, 30, 8) {real, imag} */,
  {32'h3ee79ebc, 32'h00000000} /* (31, 30, 7) {real, imag} */,
  {32'h3e906dec, 32'h00000000} /* (31, 30, 6) {real, imag} */,
  {32'h3f063631, 32'h00000000} /* (31, 30, 5) {real, imag} */,
  {32'h3f1d149b, 32'h00000000} /* (31, 30, 4) {real, imag} */,
  {32'h3eab2ae9, 32'h00000000} /* (31, 30, 3) {real, imag} */,
  {32'h3e9af77f, 32'h00000000} /* (31, 30, 2) {real, imag} */,
  {32'h3e8827be, 32'h00000000} /* (31, 30, 1) {real, imag} */,
  {32'h3e612552, 32'h00000000} /* (31, 30, 0) {real, imag} */,
  {32'h3d163b2c, 32'h00000000} /* (31, 29, 31) {real, imag} */,
  {32'h3e6aa9b2, 32'h00000000} /* (31, 29, 30) {real, imag} */,
  {32'h3eb290f7, 32'h00000000} /* (31, 29, 29) {real, imag} */,
  {32'h3d549614, 32'h00000000} /* (31, 29, 28) {real, imag} */,
  {32'h3d928bf7, 32'h00000000} /* (31, 29, 27) {real, imag} */,
  {32'h3e9ab9ef, 32'h00000000} /* (31, 29, 26) {real, imag} */,
  {32'h3f05740b, 32'h00000000} /* (31, 29, 25) {real, imag} */,
  {32'h3eeb50d8, 32'h00000000} /* (31, 29, 24) {real, imag} */,
  {32'h3ee2c90c, 32'h00000000} /* (31, 29, 23) {real, imag} */,
  {32'h3f3d953c, 32'h00000000} /* (31, 29, 22) {real, imag} */,
  {32'hbe0e976f, 32'h00000000} /* (31, 29, 21) {real, imag} */,
  {32'hbf345b0e, 32'h00000000} /* (31, 29, 20) {real, imag} */,
  {32'hbee9de45, 32'h00000000} /* (31, 29, 19) {real, imag} */,
  {32'hbf1b3a5a, 32'h00000000} /* (31, 29, 18) {real, imag} */,
  {32'hbf1a8a4c, 32'h00000000} /* (31, 29, 17) {real, imag} */,
  {32'hbf182f19, 32'h00000000} /* (31, 29, 16) {real, imag} */,
  {32'hbf3751dd, 32'h00000000} /* (31, 29, 15) {real, imag} */,
  {32'hbef3b512, 32'h00000000} /* (31, 29, 14) {real, imag} */,
  {32'hbf19bf1a, 32'h00000000} /* (31, 29, 13) {real, imag} */,
  {32'hbef7437a, 32'h00000000} /* (31, 29, 12) {real, imag} */,
  {32'hbf2075b3, 32'h00000000} /* (31, 29, 11) {real, imag} */,
  {32'hbec8ee7d, 32'h00000000} /* (31, 29, 10) {real, imag} */,
  {32'h3e444e71, 32'h00000000} /* (31, 29, 9) {real, imag} */,
  {32'h3ebe001b, 32'h00000000} /* (31, 29, 8) {real, imag} */,
  {32'h3e28b98b, 32'h00000000} /* (31, 29, 7) {real, imag} */,
  {32'h3e6342ee, 32'h00000000} /* (31, 29, 6) {real, imag} */,
  {32'h3eed5343, 32'h00000000} /* (31, 29, 5) {real, imag} */,
  {32'h3f4a3eb0, 32'h00000000} /* (31, 29, 4) {real, imag} */,
  {32'h3f1c921b, 32'h00000000} /* (31, 29, 3) {real, imag} */,
  {32'h3f1d3dc9, 32'h00000000} /* (31, 29, 2) {real, imag} */,
  {32'h3ed4184b, 32'h00000000} /* (31, 29, 1) {real, imag} */,
  {32'h3e0cd7da, 32'h00000000} /* (31, 29, 0) {real, imag} */,
  {32'h3e52330f, 32'h00000000} /* (31, 28, 31) {real, imag} */,
  {32'h3f0b399a, 32'h00000000} /* (31, 28, 30) {real, imag} */,
  {32'h3f10176e, 32'h00000000} /* (31, 28, 29) {real, imag} */,
  {32'h3e913973, 32'h00000000} /* (31, 28, 28) {real, imag} */,
  {32'h3e3641bd, 32'h00000000} /* (31, 28, 27) {real, imag} */,
  {32'h3f2162bc, 32'h00000000} /* (31, 28, 26) {real, imag} */,
  {32'h3f10bb95, 32'h00000000} /* (31, 28, 25) {real, imag} */,
  {32'h3e8bfb34, 32'h00000000} /* (31, 28, 24) {real, imag} */,
  {32'h3e4fdcde, 32'h00000000} /* (31, 28, 23) {real, imag} */,
  {32'h3e98e8d8, 32'h00000000} /* (31, 28, 22) {real, imag} */,
  {32'hbe8c20d8, 32'h00000000} /* (31, 28, 21) {real, imag} */,
  {32'hbf8dfb51, 32'h00000000} /* (31, 28, 20) {real, imag} */,
  {32'hbf17088e, 32'h00000000} /* (31, 28, 19) {real, imag} */,
  {32'hbe01761e, 32'h00000000} /* (31, 28, 18) {real, imag} */,
  {32'h3d52b4d3, 32'h00000000} /* (31, 28, 17) {real, imag} */,
  {32'hbe8e6c37, 32'h00000000} /* (31, 28, 16) {real, imag} */,
  {32'hbec9ae03, 32'h00000000} /* (31, 28, 15) {real, imag} */,
  {32'hbebb6c18, 32'h00000000} /* (31, 28, 14) {real, imag} */,
  {32'hbe88d6bf, 32'h00000000} /* (31, 28, 13) {real, imag} */,
  {32'hbe4fbd30, 32'h00000000} /* (31, 28, 12) {real, imag} */,
  {32'hbeb5270d, 32'h00000000} /* (31, 28, 11) {real, imag} */,
  {32'hbd180fe7, 32'h00000000} /* (31, 28, 10) {real, imag} */,
  {32'h3d0ea1e7, 32'h00000000} /* (31, 28, 9) {real, imag} */,
  {32'h3ea2322a, 32'h00000000} /* (31, 28, 8) {real, imag} */,
  {32'h3d7728ff, 32'h00000000} /* (31, 28, 7) {real, imag} */,
  {32'h3e31c840, 32'h00000000} /* (31, 28, 6) {real, imag} */,
  {32'h3ddb7fef, 32'h00000000} /* (31, 28, 5) {real, imag} */,
  {32'h3e44e48b, 32'h00000000} /* (31, 28, 4) {real, imag} */,
  {32'h3ea03074, 32'h00000000} /* (31, 28, 3) {real, imag} */,
  {32'h3f021cb9, 32'h00000000} /* (31, 28, 2) {real, imag} */,
  {32'h3f076606, 32'h00000000} /* (31, 28, 1) {real, imag} */,
  {32'h3e84bc9a, 32'h00000000} /* (31, 28, 0) {real, imag} */,
  {32'h3ea4a259, 32'h00000000} /* (31, 27, 31) {real, imag} */,
  {32'h3ee97714, 32'h00000000} /* (31, 27, 30) {real, imag} */,
  {32'h3e074bdc, 32'h00000000} /* (31, 27, 29) {real, imag} */,
  {32'h3e52f36a, 32'h00000000} /* (31, 27, 28) {real, imag} */,
  {32'h3f05b876, 32'h00000000} /* (31, 27, 27) {real, imag} */,
  {32'h3f7f939c, 32'h00000000} /* (31, 27, 26) {real, imag} */,
  {32'h3f2928f2, 32'h00000000} /* (31, 27, 25) {real, imag} */,
  {32'h3de0390d, 32'h00000000} /* (31, 27, 24) {real, imag} */,
  {32'h3e06674f, 32'h00000000} /* (31, 27, 23) {real, imag} */,
  {32'h3ec14da6, 32'h00000000} /* (31, 27, 22) {real, imag} */,
  {32'h3ed39770, 32'h00000000} /* (31, 27, 21) {real, imag} */,
  {32'hbe8b2afc, 32'h00000000} /* (31, 27, 20) {real, imag} */,
  {32'hbd28b1bd, 32'h00000000} /* (31, 27, 19) {real, imag} */,
  {32'hbe5060a5, 32'h00000000} /* (31, 27, 18) {real, imag} */,
  {32'hbe1d391f, 32'h00000000} /* (31, 27, 17) {real, imag} */,
  {32'hbeb4b88e, 32'h00000000} /* (31, 27, 16) {real, imag} */,
  {32'hbf1319df, 32'h00000000} /* (31, 27, 15) {real, imag} */,
  {32'hbeeb1ec7, 32'h00000000} /* (31, 27, 14) {real, imag} */,
  {32'hbe937551, 32'h00000000} /* (31, 27, 13) {real, imag} */,
  {32'h3d7a5e30, 32'h00000000} /* (31, 27, 12) {real, imag} */,
  {32'hbe1d5918, 32'h00000000} /* (31, 27, 11) {real, imag} */,
  {32'h3e51b897, 32'h00000000} /* (31, 27, 10) {real, imag} */,
  {32'h3e1f9ebc, 32'h00000000} /* (31, 27, 9) {real, imag} */,
  {32'h3e99f9dd, 32'h00000000} /* (31, 27, 8) {real, imag} */,
  {32'h3e334b2d, 32'h00000000} /* (31, 27, 7) {real, imag} */,
  {32'h3e63ad79, 32'h00000000} /* (31, 27, 6) {real, imag} */,
  {32'h3da80c3d, 32'h00000000} /* (31, 27, 5) {real, imag} */,
  {32'h3dc1e700, 32'h00000000} /* (31, 27, 4) {real, imag} */,
  {32'h3eba0df3, 32'h00000000} /* (31, 27, 3) {real, imag} */,
  {32'h3ebd240c, 32'h00000000} /* (31, 27, 2) {real, imag} */,
  {32'h3e70271a, 32'h00000000} /* (31, 27, 1) {real, imag} */,
  {32'h3dd8b7d0, 32'h00000000} /* (31, 27, 0) {real, imag} */,
  {32'h3e30f507, 32'h00000000} /* (31, 26, 31) {real, imag} */,
  {32'h3e333a70, 32'h00000000} /* (31, 26, 30) {real, imag} */,
  {32'h3cd98952, 32'h00000000} /* (31, 26, 29) {real, imag} */,
  {32'h3c64cea6, 32'h00000000} /* (31, 26, 28) {real, imag} */,
  {32'h3f118490, 32'h00000000} /* (31, 26, 27) {real, imag} */,
  {32'h3f2412e5, 32'h00000000} /* (31, 26, 26) {real, imag} */,
  {32'h3ef59179, 32'h00000000} /* (31, 26, 25) {real, imag} */,
  {32'h3f28ef3a, 32'h00000000} /* (31, 26, 24) {real, imag} */,
  {32'h3ec278f0, 32'h00000000} /* (31, 26, 23) {real, imag} */,
  {32'h3ee792a4, 32'h00000000} /* (31, 26, 22) {real, imag} */,
  {32'h3ef7a2fc, 32'h00000000} /* (31, 26, 21) {real, imag} */,
  {32'hbde200b6, 32'h00000000} /* (31, 26, 20) {real, imag} */,
  {32'hbe386d30, 32'h00000000} /* (31, 26, 19) {real, imag} */,
  {32'hbf07067e, 32'h00000000} /* (31, 26, 18) {real, imag} */,
  {32'hbea199e4, 32'h00000000} /* (31, 26, 17) {real, imag} */,
  {32'hbf12d7dd, 32'h00000000} /* (31, 26, 16) {real, imag} */,
  {32'hbf81f8d9, 32'h00000000} /* (31, 26, 15) {real, imag} */,
  {32'hbf07180d, 32'h00000000} /* (31, 26, 14) {real, imag} */,
  {32'hbea297f5, 32'h00000000} /* (31, 26, 13) {real, imag} */,
  {32'hbe8eafe1, 32'h00000000} /* (31, 26, 12) {real, imag} */,
  {32'hbedc1ea9, 32'h00000000} /* (31, 26, 11) {real, imag} */,
  {32'hbe40a0cc, 32'h00000000} /* (31, 26, 10) {real, imag} */,
  {32'h3e1f0893, 32'h00000000} /* (31, 26, 9) {real, imag} */,
  {32'h3ec656c1, 32'h00000000} /* (31, 26, 8) {real, imag} */,
  {32'h3ed6bc00, 32'h00000000} /* (31, 26, 7) {real, imag} */,
  {32'h3ecadd72, 32'h00000000} /* (31, 26, 6) {real, imag} */,
  {32'h3e8e8494, 32'h00000000} /* (31, 26, 5) {real, imag} */,
  {32'h3d9a3028, 32'h00000000} /* (31, 26, 4) {real, imag} */,
  {32'h3ed42d41, 32'h00000000} /* (31, 26, 3) {real, imag} */,
  {32'h3f13e53d, 32'h00000000} /* (31, 26, 2) {real, imag} */,
  {32'h3e9b192e, 32'h00000000} /* (31, 26, 1) {real, imag} */,
  {32'h3e0874c1, 32'h00000000} /* (31, 26, 0) {real, imag} */,
  {32'h3e1521f8, 32'h00000000} /* (31, 25, 31) {real, imag} */,
  {32'h3e9b2de8, 32'h00000000} /* (31, 25, 30) {real, imag} */,
  {32'h3d183ccf, 32'h00000000} /* (31, 25, 29) {real, imag} */,
  {32'hbd9d0731, 32'h00000000} /* (31, 25, 28) {real, imag} */,
  {32'h3ef3c31e, 32'h00000000} /* (31, 25, 27) {real, imag} */,
  {32'h3f1afd01, 32'h00000000} /* (31, 25, 26) {real, imag} */,
  {32'h3ef60661, 32'h00000000} /* (31, 25, 25) {real, imag} */,
  {32'h3f0dcf09, 32'h00000000} /* (31, 25, 24) {real, imag} */,
  {32'h3e90bbd2, 32'h00000000} /* (31, 25, 23) {real, imag} */,
  {32'h3f1bc763, 32'h00000000} /* (31, 25, 22) {real, imag} */,
  {32'h3d50d43f, 32'h00000000} /* (31, 25, 21) {real, imag} */,
  {32'hbf0221d0, 32'h00000000} /* (31, 25, 20) {real, imag} */,
  {32'hbe94e5ed, 32'h00000000} /* (31, 25, 19) {real, imag} */,
  {32'hbf052846, 32'h00000000} /* (31, 25, 18) {real, imag} */,
  {32'hbf79c0ca, 32'h00000000} /* (31, 25, 17) {real, imag} */,
  {32'hbf25c929, 32'h00000000} /* (31, 25, 16) {real, imag} */,
  {32'hbf23ecf9, 32'h00000000} /* (31, 25, 15) {real, imag} */,
  {32'hbf1e42a7, 32'h00000000} /* (31, 25, 14) {real, imag} */,
  {32'hbf082796, 32'h00000000} /* (31, 25, 13) {real, imag} */,
  {32'hbf600f13, 32'h00000000} /* (31, 25, 12) {real, imag} */,
  {32'hbf170ec7, 32'h00000000} /* (31, 25, 11) {real, imag} */,
  {32'h3d41a9ec, 32'h00000000} /* (31, 25, 10) {real, imag} */,
  {32'h3e0e59d9, 32'h00000000} /* (31, 25, 9) {real, imag} */,
  {32'h3ec12bc0, 32'h00000000} /* (31, 25, 8) {real, imag} */,
  {32'h3f0c98a6, 32'h00000000} /* (31, 25, 7) {real, imag} */,
  {32'h3f049f5e, 32'h00000000} /* (31, 25, 6) {real, imag} */,
  {32'h3f87cba3, 32'h00000000} /* (31, 25, 5) {real, imag} */,
  {32'h3ec7899b, 32'h00000000} /* (31, 25, 4) {real, imag} */,
  {32'h3ea82aa6, 32'h00000000} /* (31, 25, 3) {real, imag} */,
  {32'h3eb97e2f, 32'h00000000} /* (31, 25, 2) {real, imag} */,
  {32'h3d9af37c, 32'h00000000} /* (31, 25, 1) {real, imag} */,
  {32'h3dc89e5e, 32'h00000000} /* (31, 25, 0) {real, imag} */,
  {32'h3e94adda, 32'h00000000} /* (31, 24, 31) {real, imag} */,
  {32'h3f85fcfc, 32'h00000000} /* (31, 24, 30) {real, imag} */,
  {32'h3f6eadae, 32'h00000000} /* (31, 24, 29) {real, imag} */,
  {32'h3ec3f75f, 32'h00000000} /* (31, 24, 28) {real, imag} */,
  {32'h3e80e149, 32'h00000000} /* (31, 24, 27) {real, imag} */,
  {32'h3f1916e2, 32'h00000000} /* (31, 24, 26) {real, imag} */,
  {32'h3ecf4e21, 32'h00000000} /* (31, 24, 25) {real, imag} */,
  {32'h3eb892c4, 32'h00000000} /* (31, 24, 24) {real, imag} */,
  {32'h3ef250b1, 32'h00000000} /* (31, 24, 23) {real, imag} */,
  {32'h3f3b929b, 32'h00000000} /* (31, 24, 22) {real, imag} */,
  {32'h3ceba7dc, 32'h00000000} /* (31, 24, 21) {real, imag} */,
  {32'hbe908b01, 32'h00000000} /* (31, 24, 20) {real, imag} */,
  {32'hbd96af74, 32'h00000000} /* (31, 24, 19) {real, imag} */,
  {32'hbe61ff10, 32'h00000000} /* (31, 24, 18) {real, imag} */,
  {32'hbf68e6f2, 32'h00000000} /* (31, 24, 17) {real, imag} */,
  {32'hbf41f425, 32'h00000000} /* (31, 24, 16) {real, imag} */,
  {32'hbea4a1ad, 32'h00000000} /* (31, 24, 15) {real, imag} */,
  {32'hbefc9693, 32'h00000000} /* (31, 24, 14) {real, imag} */,
  {32'hbee1f939, 32'h00000000} /* (31, 24, 13) {real, imag} */,
  {32'hbf34f0ce, 32'h00000000} /* (31, 24, 12) {real, imag} */,
  {32'hbea26360, 32'h00000000} /* (31, 24, 11) {real, imag} */,
  {32'h3e8d2116, 32'h00000000} /* (31, 24, 10) {real, imag} */,
  {32'h3f0033a0, 32'h00000000} /* (31, 24, 9) {real, imag} */,
  {32'h3ed1a1a8, 32'h00000000} /* (31, 24, 8) {real, imag} */,
  {32'h3ef40806, 32'h00000000} /* (31, 24, 7) {real, imag} */,
  {32'h3f26709e, 32'h00000000} /* (31, 24, 6) {real, imag} */,
  {32'h3f81b1cd, 32'h00000000} /* (31, 24, 5) {real, imag} */,
  {32'h3ebda384, 32'h00000000} /* (31, 24, 4) {real, imag} */,
  {32'h3ed008b3, 32'h00000000} /* (31, 24, 3) {real, imag} */,
  {32'h3ef8e925, 32'h00000000} /* (31, 24, 2) {real, imag} */,
  {32'h3e400c80, 32'h00000000} /* (31, 24, 1) {real, imag} */,
  {32'h3dca1f93, 32'h00000000} /* (31, 24, 0) {real, imag} */,
  {32'h3e704ac0, 32'h00000000} /* (31, 23, 31) {real, imag} */,
  {32'h3f74ff38, 32'h00000000} /* (31, 23, 30) {real, imag} */,
  {32'h3f5b134f, 32'h00000000} /* (31, 23, 29) {real, imag} */,
  {32'h3ee9fc18, 32'h00000000} /* (31, 23, 28) {real, imag} */,
  {32'h3e8e3170, 32'h00000000} /* (31, 23, 27) {real, imag} */,
  {32'h3ee298ab, 32'h00000000} /* (31, 23, 26) {real, imag} */,
  {32'h3eb3f5fe, 32'h00000000} /* (31, 23, 25) {real, imag} */,
  {32'h3e7f714d, 32'h00000000} /* (31, 23, 24) {real, imag} */,
  {32'h3f59cfcb, 32'h00000000} /* (31, 23, 23) {real, imag} */,
  {32'h3f4ea371, 32'h00000000} /* (31, 23, 22) {real, imag} */,
  {32'h3ea007cc, 32'h00000000} /* (31, 23, 21) {real, imag} */,
  {32'hbda9143e, 32'h00000000} /* (31, 23, 20) {real, imag} */,
  {32'hbecf7e59, 32'h00000000} /* (31, 23, 19) {real, imag} */,
  {32'hbead5664, 32'h00000000} /* (31, 23, 18) {real, imag} */,
  {32'hbeca1e11, 32'h00000000} /* (31, 23, 17) {real, imag} */,
  {32'hbf22e29a, 32'h00000000} /* (31, 23, 16) {real, imag} */,
  {32'hbf0d2c21, 32'h00000000} /* (31, 23, 15) {real, imag} */,
  {32'hbf34536c, 32'h00000000} /* (31, 23, 14) {real, imag} */,
  {32'hbe850cb1, 32'h00000000} /* (31, 23, 13) {real, imag} */,
  {32'hbdf09aaa, 32'h00000000} /* (31, 23, 12) {real, imag} */,
  {32'hbe217f9a, 32'h00000000} /* (31, 23, 11) {real, imag} */,
  {32'h3e4921d2, 32'h00000000} /* (31, 23, 10) {real, imag} */,
  {32'h3f3806d4, 32'h00000000} /* (31, 23, 9) {real, imag} */,
  {32'h3ee5da88, 32'h00000000} /* (31, 23, 8) {real, imag} */,
  {32'h3ee85a50, 32'h00000000} /* (31, 23, 7) {real, imag} */,
  {32'h3ed84a6a, 32'h00000000} /* (31, 23, 6) {real, imag} */,
  {32'h3e8f2ae7, 32'h00000000} /* (31, 23, 5) {real, imag} */,
  {32'h3ec690ed, 32'h00000000} /* (31, 23, 4) {real, imag} */,
  {32'h3f4db94a, 32'h00000000} /* (31, 23, 3) {real, imag} */,
  {32'h3f6ae4c5, 32'h00000000} /* (31, 23, 2) {real, imag} */,
  {32'h3f2d77ce, 32'h00000000} /* (31, 23, 1) {real, imag} */,
  {32'h3f101788, 32'h00000000} /* (31, 23, 0) {real, imag} */,
  {32'h3cfd84bb, 32'h00000000} /* (31, 22, 31) {real, imag} */,
  {32'h3eddce5d, 32'h00000000} /* (31, 22, 30) {real, imag} */,
  {32'h3e831193, 32'h00000000} /* (31, 22, 29) {real, imag} */,
  {32'h3d0c0d82, 32'h00000000} /* (31, 22, 28) {real, imag} */,
  {32'hbd74f0ca, 32'h00000000} /* (31, 22, 27) {real, imag} */,
  {32'hba12a26e, 32'h00000000} /* (31, 22, 26) {real, imag} */,
  {32'h3e507a88, 32'h00000000} /* (31, 22, 25) {real, imag} */,
  {32'h3eb9cd72, 32'h00000000} /* (31, 22, 24) {real, imag} */,
  {32'h3f90c7fb, 32'h00000000} /* (31, 22, 23) {real, imag} */,
  {32'h3f8a96c7, 32'h00000000} /* (31, 22, 22) {real, imag} */,
  {32'h3edecf73, 32'h00000000} /* (31, 22, 21) {real, imag} */,
  {32'hbe083ef0, 32'h00000000} /* (31, 22, 20) {real, imag} */,
  {32'hbf2ec05e, 32'h00000000} /* (31, 22, 19) {real, imag} */,
  {32'hbef4caab, 32'h00000000} /* (31, 22, 18) {real, imag} */,
  {32'hbf25c53d, 32'h00000000} /* (31, 22, 17) {real, imag} */,
  {32'hbf6a0c15, 32'h00000000} /* (31, 22, 16) {real, imag} */,
  {32'hbf198ecc, 32'h00000000} /* (31, 22, 15) {real, imag} */,
  {32'hbf10e5a9, 32'h00000000} /* (31, 22, 14) {real, imag} */,
  {32'hbe451a3b, 32'h00000000} /* (31, 22, 13) {real, imag} */,
  {32'hbe3ef435, 32'h00000000} /* (31, 22, 12) {real, imag} */,
  {32'hbe63011e, 32'h00000000} /* (31, 22, 11) {real, imag} */,
  {32'h3eab2721, 32'h00000000} /* (31, 22, 10) {real, imag} */,
  {32'h3f6ffa98, 32'h00000000} /* (31, 22, 9) {real, imag} */,
  {32'h3f2b260d, 32'h00000000} /* (31, 22, 8) {real, imag} */,
  {32'h3ec8e206, 32'h00000000} /* (31, 22, 7) {real, imag} */,
  {32'h3e96c2ee, 32'h00000000} /* (31, 22, 6) {real, imag} */,
  {32'h3ec768dd, 32'h00000000} /* (31, 22, 5) {real, imag} */,
  {32'h3f76a992, 32'h00000000} /* (31, 22, 4) {real, imag} */,
  {32'h3f6a0567, 32'h00000000} /* (31, 22, 3) {real, imag} */,
  {32'h3f8b9cbe, 32'h00000000} /* (31, 22, 2) {real, imag} */,
  {32'h3f37fa7d, 32'h00000000} /* (31, 22, 1) {real, imag} */,
  {32'h3ee8b058, 32'h00000000} /* (31, 22, 0) {real, imag} */,
  {32'hbc502b2e, 32'h00000000} /* (31, 21, 31) {real, imag} */,
  {32'h3ea5286f, 32'h00000000} /* (31, 21, 30) {real, imag} */,
  {32'h3e20946d, 32'h00000000} /* (31, 21, 29) {real, imag} */,
  {32'h3e36743d, 32'h00000000} /* (31, 21, 28) {real, imag} */,
  {32'hbd218469, 32'h00000000} /* (31, 21, 27) {real, imag} */,
  {32'h3dd5b512, 32'h00000000} /* (31, 21, 26) {real, imag} */,
  {32'h3d99ebf4, 32'h00000000} /* (31, 21, 25) {real, imag} */,
  {32'hbd020e4c, 32'h00000000} /* (31, 21, 24) {real, imag} */,
  {32'h3eec61b9, 32'h00000000} /* (31, 21, 23) {real, imag} */,
  {32'h3e24fb05, 32'h00000000} /* (31, 21, 22) {real, imag} */,
  {32'hbc2c0cb9, 32'h00000000} /* (31, 21, 21) {real, imag} */,
  {32'h3c41cfa6, 32'h00000000} /* (31, 21, 20) {real, imag} */,
  {32'hbe7b559e, 32'h00000000} /* (31, 21, 19) {real, imag} */,
  {32'hbec2bc7f, 32'h00000000} /* (31, 21, 18) {real, imag} */,
  {32'hbf3bcb0f, 32'h00000000} /* (31, 21, 17) {real, imag} */,
  {32'hbedba952, 32'h00000000} /* (31, 21, 16) {real, imag} */,
  {32'hbe21cbc1, 32'h00000000} /* (31, 21, 15) {real, imag} */,
  {32'hbeb4edfb, 32'h00000000} /* (31, 21, 14) {real, imag} */,
  {32'h3ca9c948, 32'h00000000} /* (31, 21, 13) {real, imag} */,
  {32'h3db91413, 32'h00000000} /* (31, 21, 12) {real, imag} */,
  {32'h3d80d951, 32'h00000000} /* (31, 21, 11) {real, imag} */,
  {32'h3dd24f46, 32'h00000000} /* (31, 21, 10) {real, imag} */,
  {32'h3f148fff, 32'h00000000} /* (31, 21, 9) {real, imag} */,
  {32'h3ebac2e2, 32'h00000000} /* (31, 21, 8) {real, imag} */,
  {32'hbb7ee332, 32'h00000000} /* (31, 21, 7) {real, imag} */,
  {32'h3e24e202, 32'h00000000} /* (31, 21, 6) {real, imag} */,
  {32'h3e5e6d1e, 32'h00000000} /* (31, 21, 5) {real, imag} */,
  {32'h3f135b11, 32'h00000000} /* (31, 21, 4) {real, imag} */,
  {32'h3ebb17c4, 32'h00000000} /* (31, 21, 3) {real, imag} */,
  {32'h3ecd8785, 32'h00000000} /* (31, 21, 2) {real, imag} */,
  {32'h3e140c11, 32'h00000000} /* (31, 21, 1) {real, imag} */,
  {32'hbe41c9d6, 32'h00000000} /* (31, 21, 0) {real, imag} */,
  {32'hbdeea136, 32'h00000000} /* (31, 20, 31) {real, imag} */,
  {32'hbe5a5e8a, 32'h00000000} /* (31, 20, 30) {real, imag} */,
  {32'hbec0ce3e, 32'h00000000} /* (31, 20, 29) {real, imag} */,
  {32'hbd746893, 32'h00000000} /* (31, 20, 28) {real, imag} */,
  {32'hbe7fe2dc, 32'h00000000} /* (31, 20, 27) {real, imag} */,
  {32'hbe4b0b28, 32'h00000000} /* (31, 20, 26) {real, imag} */,
  {32'hbe0e5673, 32'h00000000} /* (31, 20, 25) {real, imag} */,
  {32'hbf7127ae, 32'h00000000} /* (31, 20, 24) {real, imag} */,
  {32'hbf3f0610, 32'h00000000} /* (31, 20, 23) {real, imag} */,
  {32'hbec18bb8, 32'h00000000} /* (31, 20, 22) {real, imag} */,
  {32'hbeb2cb2b, 32'h00000000} /* (31, 20, 21) {real, imag} */,
  {32'h3d472104, 32'h00000000} /* (31, 20, 20) {real, imag} */,
  {32'h3cabcca5, 32'h00000000} /* (31, 20, 19) {real, imag} */,
  {32'h3d985fc0, 32'h00000000} /* (31, 20, 18) {real, imag} */,
  {32'hbe3db503, 32'h00000000} /* (31, 20, 17) {real, imag} */,
  {32'h3d99cf22, 32'h00000000} /* (31, 20, 16) {real, imag} */,
  {32'h3eb860ab, 32'h00000000} /* (31, 20, 15) {real, imag} */,
  {32'h3e8bfaa5, 32'h00000000} /* (31, 20, 14) {real, imag} */,
  {32'h3f56f51d, 32'h00000000} /* (31, 20, 13) {real, imag} */,
  {32'h3f2372e3, 32'h00000000} /* (31, 20, 12) {real, imag} */,
  {32'h3e844226, 32'h00000000} /* (31, 20, 11) {real, imag} */,
  {32'hbda3ea49, 32'h00000000} /* (31, 20, 10) {real, imag} */,
  {32'hbddaa003, 32'h00000000} /* (31, 20, 9) {real, imag} */,
  {32'hbf0f05cc, 32'h00000000} /* (31, 20, 8) {real, imag} */,
  {32'hbf6798c0, 32'h00000000} /* (31, 20, 7) {real, imag} */,
  {32'hbf5990c7, 32'h00000000} /* (31, 20, 6) {real, imag} */,
  {32'hbeb60453, 32'h00000000} /* (31, 20, 5) {real, imag} */,
  {32'hbeec7d8b, 32'h00000000} /* (31, 20, 4) {real, imag} */,
  {32'hbf250813, 32'h00000000} /* (31, 20, 3) {real, imag} */,
  {32'hbea8afbb, 32'h00000000} /* (31, 20, 2) {real, imag} */,
  {32'hbed051a0, 32'h00000000} /* (31, 20, 1) {real, imag} */,
  {32'hbf0a03de, 32'h00000000} /* (31, 20, 0) {real, imag} */,
  {32'hbe805659, 32'h00000000} /* (31, 19, 31) {real, imag} */,
  {32'hbeade18c, 32'h00000000} /* (31, 19, 30) {real, imag} */,
  {32'hbe3531df, 32'h00000000} /* (31, 19, 29) {real, imag} */,
  {32'hbebe6ed4, 32'h00000000} /* (31, 19, 28) {real, imag} */,
  {32'hbedec4e3, 32'h00000000} /* (31, 19, 27) {real, imag} */,
  {32'hbf267b99, 32'h00000000} /* (31, 19, 26) {real, imag} */,
  {32'hbf34b518, 32'h00000000} /* (31, 19, 25) {real, imag} */,
  {32'hbf487a6c, 32'h00000000} /* (31, 19, 24) {real, imag} */,
  {32'hbf7cf2be, 32'h00000000} /* (31, 19, 23) {real, imag} */,
  {32'hbed04d88, 32'h00000000} /* (31, 19, 22) {real, imag} */,
  {32'hbe93aa5b, 32'h00000000} /* (31, 19, 21) {real, imag} */,
  {32'h3d98024d, 32'h00000000} /* (31, 19, 20) {real, imag} */,
  {32'h3ef77df4, 32'h00000000} /* (31, 19, 19) {real, imag} */,
  {32'h3f494efc, 32'h00000000} /* (31, 19, 18) {real, imag} */,
  {32'h3e756756, 32'h00000000} /* (31, 19, 17) {real, imag} */,
  {32'h3edcbfca, 32'h00000000} /* (31, 19, 16) {real, imag} */,
  {32'h3f5044bf, 32'h00000000} /* (31, 19, 15) {real, imag} */,
  {32'h3f2998e7, 32'h00000000} /* (31, 19, 14) {real, imag} */,
  {32'h3f8df596, 32'h00000000} /* (31, 19, 13) {real, imag} */,
  {32'h3f6fcb1b, 32'h00000000} /* (31, 19, 12) {real, imag} */,
  {32'h3f1078dc, 32'h00000000} /* (31, 19, 11) {real, imag} */,
  {32'hbe879ff9, 32'h00000000} /* (31, 19, 10) {real, imag} */,
  {32'hbf5d24d2, 32'h00000000} /* (31, 19, 9) {real, imag} */,
  {32'hbf8563b7, 32'h00000000} /* (31, 19, 8) {real, imag} */,
  {32'hbf45d8a5, 32'h00000000} /* (31, 19, 7) {real, imag} */,
  {32'hbf0ecd98, 32'h00000000} /* (31, 19, 6) {real, imag} */,
  {32'hbe46770e, 32'h00000000} /* (31, 19, 5) {real, imag} */,
  {32'hbf0d58f0, 32'h00000000} /* (31, 19, 4) {real, imag} */,
  {32'hbf7ecfa6, 32'h00000000} /* (31, 19, 3) {real, imag} */,
  {32'hbeff31b3, 32'h00000000} /* (31, 19, 2) {real, imag} */,
  {32'hbf3388fc, 32'h00000000} /* (31, 19, 1) {real, imag} */,
  {32'hbf186c3c, 32'h00000000} /* (31, 19, 0) {real, imag} */,
  {32'hbf1e4f65, 32'h00000000} /* (31, 18, 31) {real, imag} */,
  {32'hbee541ac, 32'h00000000} /* (31, 18, 30) {real, imag} */,
  {32'hbdf76f72, 32'h00000000} /* (31, 18, 29) {real, imag} */,
  {32'hbe607e40, 32'h00000000} /* (31, 18, 28) {real, imag} */,
  {32'hbe13fabe, 32'h00000000} /* (31, 18, 27) {real, imag} */,
  {32'hbe6e947d, 32'h00000000} /* (31, 18, 26) {real, imag} */,
  {32'hbe9dedb6, 32'h00000000} /* (31, 18, 25) {real, imag} */,
  {32'hbe9a012c, 32'h00000000} /* (31, 18, 24) {real, imag} */,
  {32'hbf117b4a, 32'h00000000} /* (31, 18, 23) {real, imag} */,
  {32'hbe60f4be, 32'h00000000} /* (31, 18, 22) {real, imag} */,
  {32'hbc5c0cb4, 32'h00000000} /* (31, 18, 21) {real, imag} */,
  {32'h3f1d2ddf, 32'h00000000} /* (31, 18, 20) {real, imag} */,
  {32'h3f4c8218, 32'h00000000} /* (31, 18, 19) {real, imag} */,
  {32'h3f28afa2, 32'h00000000} /* (31, 18, 18) {real, imag} */,
  {32'h3ea65c40, 32'h00000000} /* (31, 18, 17) {real, imag} */,
  {32'h3eaa3142, 32'h00000000} /* (31, 18, 16) {real, imag} */,
  {32'h3f0a1b4f, 32'h00000000} /* (31, 18, 15) {real, imag} */,
  {32'h3f0d8d7e, 32'h00000000} /* (31, 18, 14) {real, imag} */,
  {32'h3f5b7bf8, 32'h00000000} /* (31, 18, 13) {real, imag} */,
  {32'h3f6e2e28, 32'h00000000} /* (31, 18, 12) {real, imag} */,
  {32'h3f108f7d, 32'h00000000} /* (31, 18, 11) {real, imag} */,
  {32'hbeb5b1ea, 32'h00000000} /* (31, 18, 10) {real, imag} */,
  {32'hbf6564b1, 32'h00000000} /* (31, 18, 9) {real, imag} */,
  {32'hbf580500, 32'h00000000} /* (31, 18, 8) {real, imag} */,
  {32'hbf384494, 32'h00000000} /* (31, 18, 7) {real, imag} */,
  {32'hbec78edb, 32'h00000000} /* (31, 18, 6) {real, imag} */,
  {32'h3cd4183d, 32'h00000000} /* (31, 18, 5) {real, imag} */,
  {32'hbde5a99b, 32'h00000000} /* (31, 18, 4) {real, imag} */,
  {32'hbea3a33e, 32'h00000000} /* (31, 18, 3) {real, imag} */,
  {32'hbece6acf, 32'h00000000} /* (31, 18, 2) {real, imag} */,
  {32'hbf13ac7d, 32'h00000000} /* (31, 18, 1) {real, imag} */,
  {32'hbea01d3c, 32'h00000000} /* (31, 18, 0) {real, imag} */,
  {32'hbebcde44, 32'h00000000} /* (31, 17, 31) {real, imag} */,
  {32'hbeb3a125, 32'h00000000} /* (31, 17, 30) {real, imag} */,
  {32'hbe6ec996, 32'h00000000} /* (31, 17, 29) {real, imag} */,
  {32'hbd8a55d2, 32'h00000000} /* (31, 17, 28) {real, imag} */,
  {32'hbe00cfbc, 32'h00000000} /* (31, 17, 27) {real, imag} */,
  {32'hbd48965f, 32'h00000000} /* (31, 17, 26) {real, imag} */,
  {32'hbc07e1f7, 32'h00000000} /* (31, 17, 25) {real, imag} */,
  {32'hbd3ccc15, 32'h00000000} /* (31, 17, 24) {real, imag} */,
  {32'hbe08ca6b, 32'h00000000} /* (31, 17, 23) {real, imag} */,
  {32'hbe8ef961, 32'h00000000} /* (31, 17, 22) {real, imag} */,
  {32'h3d27f8a6, 32'h00000000} /* (31, 17, 21) {real, imag} */,
  {32'h3f8d8479, 32'h00000000} /* (31, 17, 20) {real, imag} */,
  {32'h3f30fc94, 32'h00000000} /* (31, 17, 19) {real, imag} */,
  {32'h3f0201fc, 32'h00000000} /* (31, 17, 18) {real, imag} */,
  {32'h3ee052b0, 32'h00000000} /* (31, 17, 17) {real, imag} */,
  {32'h3eb337cd, 32'h00000000} /* (31, 17, 16) {real, imag} */,
  {32'h3edafe5f, 32'h00000000} /* (31, 17, 15) {real, imag} */,
  {32'h3f0c3011, 32'h00000000} /* (31, 17, 14) {real, imag} */,
  {32'h3ee24bd2, 32'h00000000} /* (31, 17, 13) {real, imag} */,
  {32'h3f195f1c, 32'h00000000} /* (31, 17, 12) {real, imag} */,
  {32'h3efd3c19, 32'h00000000} /* (31, 17, 11) {real, imag} */,
  {32'hbe914f2b, 32'h00000000} /* (31, 17, 10) {real, imag} */,
  {32'hbf320a9d, 32'h00000000} /* (31, 17, 9) {real, imag} */,
  {32'hbf23d955, 32'h00000000} /* (31, 17, 8) {real, imag} */,
  {32'hbe8e657e, 32'h00000000} /* (31, 17, 7) {real, imag} */,
  {32'hbea647a7, 32'h00000000} /* (31, 17, 6) {real, imag} */,
  {32'hbeb7b1a8, 32'h00000000} /* (31, 17, 5) {real, imag} */,
  {32'hbe8e0430, 32'h00000000} /* (31, 17, 4) {real, imag} */,
  {32'hbea6968b, 32'h00000000} /* (31, 17, 3) {real, imag} */,
  {32'hbed2a181, 32'h00000000} /* (31, 17, 2) {real, imag} */,
  {32'hbf447441, 32'h00000000} /* (31, 17, 1) {real, imag} */,
  {32'hbecffd6d, 32'h00000000} /* (31, 17, 0) {real, imag} */,
  {32'hbe7b0f2f, 32'h00000000} /* (31, 16, 31) {real, imag} */,
  {32'hbeb4df01, 32'h00000000} /* (31, 16, 30) {real, imag} */,
  {32'hbed992ec, 32'h00000000} /* (31, 16, 29) {real, imag} */,
  {32'h3dabd3eb, 32'h00000000} /* (31, 16, 28) {real, imag} */,
  {32'h3da69a1a, 32'h00000000} /* (31, 16, 27) {real, imag} */,
  {32'hbdda7104, 32'h00000000} /* (31, 16, 26) {real, imag} */,
  {32'hbdfec29a, 32'h00000000} /* (31, 16, 25) {real, imag} */,
  {32'hbea2fd7d, 32'h00000000} /* (31, 16, 24) {real, imag} */,
  {32'hbe955d1a, 32'h00000000} /* (31, 16, 23) {real, imag} */,
  {32'hbe8213eb, 32'h00000000} /* (31, 16, 22) {real, imag} */,
  {32'h3d21b62f, 32'h00000000} /* (31, 16, 21) {real, imag} */,
  {32'h3f35f92e, 32'h00000000} /* (31, 16, 20) {real, imag} */,
  {32'h3f0a3ac7, 32'h00000000} /* (31, 16, 19) {real, imag} */,
  {32'h3ece05bc, 32'h00000000} /* (31, 16, 18) {real, imag} */,
  {32'h3e989c12, 32'h00000000} /* (31, 16, 17) {real, imag} */,
  {32'h3ebd4ea7, 32'h00000000} /* (31, 16, 16) {real, imag} */,
  {32'h3eb4d9cb, 32'h00000000} /* (31, 16, 15) {real, imag} */,
  {32'h3eeca9b4, 32'h00000000} /* (31, 16, 14) {real, imag} */,
  {32'h3f1e207f, 32'h00000000} /* (31, 16, 13) {real, imag} */,
  {32'h3f4f0fa2, 32'h00000000} /* (31, 16, 12) {real, imag} */,
  {32'h3def9582, 32'h00000000} /* (31, 16, 11) {real, imag} */,
  {32'hbf25a71a, 32'h00000000} /* (31, 16, 10) {real, imag} */,
  {32'hbf155dfa, 32'h00000000} /* (31, 16, 9) {real, imag} */,
  {32'hbe930ad4, 32'h00000000} /* (31, 16, 8) {real, imag} */,
  {32'hbe7ecde6, 32'h00000000} /* (31, 16, 7) {real, imag} */,
  {32'hbf37167a, 32'h00000000} /* (31, 16, 6) {real, imag} */,
  {32'hbf1f4806, 32'h00000000} /* (31, 16, 5) {real, imag} */,
  {32'hbee806af, 32'h00000000} /* (31, 16, 4) {real, imag} */,
  {32'hbea2aba4, 32'h00000000} /* (31, 16, 3) {real, imag} */,
  {32'hbed47a75, 32'h00000000} /* (31, 16, 2) {real, imag} */,
  {32'hbf4107e9, 32'h00000000} /* (31, 16, 1) {real, imag} */,
  {32'hbed5e609, 32'h00000000} /* (31, 16, 0) {real, imag} */,
  {32'hbebe68aa, 32'h00000000} /* (31, 15, 31) {real, imag} */,
  {32'hbf0a07b6, 32'h00000000} /* (31, 15, 30) {real, imag} */,
  {32'hbf1f16c3, 32'h00000000} /* (31, 15, 29) {real, imag} */,
  {32'hbe6d33de, 32'h00000000} /* (31, 15, 28) {real, imag} */,
  {32'hbdbd7e58, 32'h00000000} /* (31, 15, 27) {real, imag} */,
  {32'hbcb8c7bc, 32'h00000000} /* (31, 15, 26) {real, imag} */,
  {32'hbd9ed984, 32'h00000000} /* (31, 15, 25) {real, imag} */,
  {32'hbe2a9eb1, 32'h00000000} /* (31, 15, 24) {real, imag} */,
  {32'hbe8fe485, 32'h00000000} /* (31, 15, 23) {real, imag} */,
  {32'hbe494f87, 32'h00000000} /* (31, 15, 22) {real, imag} */,
  {32'hbd10d37d, 32'h00000000} /* (31, 15, 21) {real, imag} */,
  {32'h3e39c5f9, 32'h00000000} /* (31, 15, 20) {real, imag} */,
  {32'h3ea8255d, 32'h00000000} /* (31, 15, 19) {real, imag} */,
  {32'h3e970d83, 32'h00000000} /* (31, 15, 18) {real, imag} */,
  {32'h3dd6d3a0, 32'h00000000} /* (31, 15, 17) {real, imag} */,
  {32'h3e84738a, 32'h00000000} /* (31, 15, 16) {real, imag} */,
  {32'h3ee46865, 32'h00000000} /* (31, 15, 15) {real, imag} */,
  {32'h3ede91a3, 32'h00000000} /* (31, 15, 14) {real, imag} */,
  {32'h3edcc797, 32'h00000000} /* (31, 15, 13) {real, imag} */,
  {32'h3e758238, 32'h00000000} /* (31, 15, 12) {real, imag} */,
  {32'hbd6e87d8, 32'h00000000} /* (31, 15, 11) {real, imag} */,
  {32'hbf161d30, 32'h00000000} /* (31, 15, 10) {real, imag} */,
  {32'hbf085e22, 32'h00000000} /* (31, 15, 9) {real, imag} */,
  {32'hbec3d85c, 32'h00000000} /* (31, 15, 8) {real, imag} */,
  {32'hbef253f8, 32'h00000000} /* (31, 15, 7) {real, imag} */,
  {32'hbef9f290, 32'h00000000} /* (31, 15, 6) {real, imag} */,
  {32'hbf025b6c, 32'h00000000} /* (31, 15, 5) {real, imag} */,
  {32'hbf03ce2c, 32'h00000000} /* (31, 15, 4) {real, imag} */,
  {32'hbe9f4981, 32'h00000000} /* (31, 15, 3) {real, imag} */,
  {32'hbe9a4e9b, 32'h00000000} /* (31, 15, 2) {real, imag} */,
  {32'hbf0c0a96, 32'h00000000} /* (31, 15, 1) {real, imag} */,
  {32'hbe3dd784, 32'h00000000} /* (31, 15, 0) {real, imag} */,
  {32'hbe9e9540, 32'h00000000} /* (31, 14, 31) {real, imag} */,
  {32'hbf344da6, 32'h00000000} /* (31, 14, 30) {real, imag} */,
  {32'hbf2728fd, 32'h00000000} /* (31, 14, 29) {real, imag} */,
  {32'hbee0b50c, 32'h00000000} /* (31, 14, 28) {real, imag} */,
  {32'hbebe224f, 32'h00000000} /* (31, 14, 27) {real, imag} */,
  {32'hbe510695, 32'h00000000} /* (31, 14, 26) {real, imag} */,
  {32'hbe98a3b7, 32'h00000000} /* (31, 14, 25) {real, imag} */,
  {32'hbe30d6df, 32'h00000000} /* (31, 14, 24) {real, imag} */,
  {32'hbdb36294, 32'h00000000} /* (31, 14, 23) {real, imag} */,
  {32'hbec39880, 32'h00000000} /* (31, 14, 22) {real, imag} */,
  {32'hbe14bae6, 32'h00000000} /* (31, 14, 21) {real, imag} */,
  {32'h3edf988e, 32'h00000000} /* (31, 14, 20) {real, imag} */,
  {32'h3e7571c0, 32'h00000000} /* (31, 14, 19) {real, imag} */,
  {32'h3e2dc120, 32'h00000000} /* (31, 14, 18) {real, imag} */,
  {32'h3e08473f, 32'h00000000} /* (31, 14, 17) {real, imag} */,
  {32'h3eb027d2, 32'h00000000} /* (31, 14, 16) {real, imag} */,
  {32'h3f015881, 32'h00000000} /* (31, 14, 15) {real, imag} */,
  {32'h3def910f, 32'h00000000} /* (31, 14, 14) {real, imag} */,
  {32'hbd57a482, 32'h00000000} /* (31, 14, 13) {real, imag} */,
  {32'h3d16b26c, 32'h00000000} /* (31, 14, 12) {real, imag} */,
  {32'h3d6fa70e, 32'h00000000} /* (31, 14, 11) {real, imag} */,
  {32'hbe81cdca, 32'h00000000} /* (31, 14, 10) {real, imag} */,
  {32'hbef882c9, 32'h00000000} /* (31, 14, 9) {real, imag} */,
  {32'hbf269822, 32'h00000000} /* (31, 14, 8) {real, imag} */,
  {32'hbeab0fec, 32'h00000000} /* (31, 14, 7) {real, imag} */,
  {32'hbe919979, 32'h00000000} /* (31, 14, 6) {real, imag} */,
  {32'hbf1387ac, 32'h00000000} /* (31, 14, 5) {real, imag} */,
  {32'hbe95a531, 32'h00000000} /* (31, 14, 4) {real, imag} */,
  {32'hbe6e0d7a, 32'h00000000} /* (31, 14, 3) {real, imag} */,
  {32'hbe50be93, 32'h00000000} /* (31, 14, 2) {real, imag} */,
  {32'hbd102602, 32'h00000000} /* (31, 14, 1) {real, imag} */,
  {32'hbd27d926, 32'h00000000} /* (31, 14, 0) {real, imag} */,
  {32'hbea46dbd, 32'h00000000} /* (31, 13, 31) {real, imag} */,
  {32'hbf16a95f, 32'h00000000} /* (31, 13, 30) {real, imag} */,
  {32'hbeb98c70, 32'h00000000} /* (31, 13, 29) {real, imag} */,
  {32'hbe3bcba7, 32'h00000000} /* (31, 13, 28) {real, imag} */,
  {32'hbe9c612f, 32'h00000000} /* (31, 13, 27) {real, imag} */,
  {32'hbef534af, 32'h00000000} /* (31, 13, 26) {real, imag} */,
  {32'hbed4018f, 32'h00000000} /* (31, 13, 25) {real, imag} */,
  {32'hbf2efc09, 32'h00000000} /* (31, 13, 24) {real, imag} */,
  {32'hbf0eac7c, 32'h00000000} /* (31, 13, 23) {real, imag} */,
  {32'hbf16dacd, 32'h00000000} /* (31, 13, 22) {real, imag} */,
  {32'hbe9de47d, 32'h00000000} /* (31, 13, 21) {real, imag} */,
  {32'h3e8c7652, 32'h00000000} /* (31, 13, 20) {real, imag} */,
  {32'h3e92745c, 32'h00000000} /* (31, 13, 19) {real, imag} */,
  {32'h3def591a, 32'h00000000} /* (31, 13, 18) {real, imag} */,
  {32'h3e9b1905, 32'h00000000} /* (31, 13, 17) {real, imag} */,
  {32'h3ed1dcf5, 32'h00000000} /* (31, 13, 16) {real, imag} */,
  {32'h3f2897fa, 32'h00000000} /* (31, 13, 15) {real, imag} */,
  {32'h3ecf138b, 32'h00000000} /* (31, 13, 14) {real, imag} */,
  {32'h3e851e4b, 32'h00000000} /* (31, 13, 13) {real, imag} */,
  {32'h3e695ff9, 32'h00000000} /* (31, 13, 12) {real, imag} */,
  {32'h3d114db0, 32'h00000000} /* (31, 13, 11) {real, imag} */,
  {32'hbe04bd64, 32'h00000000} /* (31, 13, 10) {real, imag} */,
  {32'hbf2c3eb0, 32'h00000000} /* (31, 13, 9) {real, imag} */,
  {32'hbf9dde84, 32'h00000000} /* (31, 13, 8) {real, imag} */,
  {32'hbf205f8f, 32'h00000000} /* (31, 13, 7) {real, imag} */,
  {32'hbf299516, 32'h00000000} /* (31, 13, 6) {real, imag} */,
  {32'hbf3aee51, 32'h00000000} /* (31, 13, 5) {real, imag} */,
  {32'hbec99dab, 32'h00000000} /* (31, 13, 4) {real, imag} */,
  {32'hbec5c6f5, 32'h00000000} /* (31, 13, 3) {real, imag} */,
  {32'hbea5304a, 32'h00000000} /* (31, 13, 2) {real, imag} */,
  {32'hbe88ae3e, 32'h00000000} /* (31, 13, 1) {real, imag} */,
  {32'hbe87deb7, 32'h00000000} /* (31, 13, 0) {real, imag} */,
  {32'hbee67ee3, 32'h00000000} /* (31, 12, 31) {real, imag} */,
  {32'hbf21eebd, 32'h00000000} /* (31, 12, 30) {real, imag} */,
  {32'hbea33211, 32'h00000000} /* (31, 12, 29) {real, imag} */,
  {32'hbe7a9398, 32'h00000000} /* (31, 12, 28) {real, imag} */,
  {32'hbf351e75, 32'h00000000} /* (31, 12, 27) {real, imag} */,
  {32'hbf614abc, 32'h00000000} /* (31, 12, 26) {real, imag} */,
  {32'hbea1d2ba, 32'h00000000} /* (31, 12, 25) {real, imag} */,
  {32'hbef0c640, 32'h00000000} /* (31, 12, 24) {real, imag} */,
  {32'hbf41f11e, 32'h00000000} /* (31, 12, 23) {real, imag} */,
  {32'hbf60d557, 32'h00000000} /* (31, 12, 22) {real, imag} */,
  {32'hbe7ea972, 32'h00000000} /* (31, 12, 21) {real, imag} */,
  {32'h3e065e2e, 32'h00000000} /* (31, 12, 20) {real, imag} */,
  {32'h3e8a9b8f, 32'h00000000} /* (31, 12, 19) {real, imag} */,
  {32'h3e8d57c8, 32'h00000000} /* (31, 12, 18) {real, imag} */,
  {32'h3f2155ae, 32'h00000000} /* (31, 12, 17) {real, imag} */,
  {32'h3f4775aa, 32'h00000000} /* (31, 12, 16) {real, imag} */,
  {32'h3f04e484, 32'h00000000} /* (31, 12, 15) {real, imag} */,
  {32'h3f0179bc, 32'h00000000} /* (31, 12, 14) {real, imag} */,
  {32'h3ed2bb35, 32'h00000000} /* (31, 12, 13) {real, imag} */,
  {32'h3f2ff0ef, 32'h00000000} /* (31, 12, 12) {real, imag} */,
  {32'h3ed0b7d3, 32'h00000000} /* (31, 12, 11) {real, imag} */,
  {32'hbe818163, 32'h00000000} /* (31, 12, 10) {real, imag} */,
  {32'hbf41d99b, 32'h00000000} /* (31, 12, 9) {real, imag} */,
  {32'hbf9196cb, 32'h00000000} /* (31, 12, 8) {real, imag} */,
  {32'hbf10304e, 32'h00000000} /* (31, 12, 7) {real, imag} */,
  {32'hbf3d3e90, 32'h00000000} /* (31, 12, 6) {real, imag} */,
  {32'hbf170868, 32'h00000000} /* (31, 12, 5) {real, imag} */,
  {32'hbec2c5b6, 32'h00000000} /* (31, 12, 4) {real, imag} */,
  {32'hbef19a6f, 32'h00000000} /* (31, 12, 3) {real, imag} */,
  {32'hbea10da0, 32'h00000000} /* (31, 12, 2) {real, imag} */,
  {32'hbf0a8de9, 32'h00000000} /* (31, 12, 1) {real, imag} */,
  {32'hbf0f899c, 32'h00000000} /* (31, 12, 0) {real, imag} */,
  {32'hbdf74d91, 32'h00000000} /* (31, 11, 31) {real, imag} */,
  {32'hbefd9798, 32'h00000000} /* (31, 11, 30) {real, imag} */,
  {32'hbed9cd2d, 32'h00000000} /* (31, 11, 29) {real, imag} */,
  {32'hbec9e7a9, 32'h00000000} /* (31, 11, 28) {real, imag} */,
  {32'hbf195773, 32'h00000000} /* (31, 11, 27) {real, imag} */,
  {32'hbe9c5c77, 32'h00000000} /* (31, 11, 26) {real, imag} */,
  {32'hbe661029, 32'h00000000} /* (31, 11, 25) {real, imag} */,
  {32'hbe816005, 32'h00000000} /* (31, 11, 24) {real, imag} */,
  {32'hbeb91dc8, 32'h00000000} /* (31, 11, 23) {real, imag} */,
  {32'hbf315fce, 32'h00000000} /* (31, 11, 22) {real, imag} */,
  {32'hbd9b9911, 32'h00000000} /* (31, 11, 21) {real, imag} */,
  {32'h3eb32197, 32'h00000000} /* (31, 11, 20) {real, imag} */,
  {32'h3e90f33d, 32'h00000000} /* (31, 11, 19) {real, imag} */,
  {32'h3ee39619, 32'h00000000} /* (31, 11, 18) {real, imag} */,
  {32'h3f76f78c, 32'h00000000} /* (31, 11, 17) {real, imag} */,
  {32'h3f43d7be, 32'h00000000} /* (31, 11, 16) {real, imag} */,
  {32'h3e0289b8, 32'h00000000} /* (31, 11, 15) {real, imag} */,
  {32'h3ef7fef5, 32'h00000000} /* (31, 11, 14) {real, imag} */,
  {32'h3e3c84c3, 32'h00000000} /* (31, 11, 13) {real, imag} */,
  {32'h3f091768, 32'h00000000} /* (31, 11, 12) {real, imag} */,
  {32'h3ee6cf24, 32'h00000000} /* (31, 11, 11) {real, imag} */,
  {32'hbe3f93ae, 32'h00000000} /* (31, 11, 10) {real, imag} */,
  {32'hbee93af1, 32'h00000000} /* (31, 11, 9) {real, imag} */,
  {32'hbeb69d8b, 32'h00000000} /* (31, 11, 8) {real, imag} */,
  {32'hbc8396fb, 32'h00000000} /* (31, 11, 7) {real, imag} */,
  {32'hbe69863c, 32'h00000000} /* (31, 11, 6) {real, imag} */,
  {32'hbf107b8c, 32'h00000000} /* (31, 11, 5) {real, imag} */,
  {32'hbe550b50, 32'h00000000} /* (31, 11, 4) {real, imag} */,
  {32'hbee1d6b9, 32'h00000000} /* (31, 11, 3) {real, imag} */,
  {32'hbe425c6f, 32'h00000000} /* (31, 11, 2) {real, imag} */,
  {32'hbdc5b7a0, 32'h00000000} /* (31, 11, 1) {real, imag} */,
  {32'hbdff6c78, 32'h00000000} /* (31, 11, 0) {real, imag} */,
  {32'h3f1fb758, 32'h00000000} /* (31, 10, 31) {real, imag} */,
  {32'h3ec26713, 32'h00000000} /* (31, 10, 30) {real, imag} */,
  {32'hbe2e8360, 32'h00000000} /* (31, 10, 29) {real, imag} */,
  {32'hbe1e13fb, 32'h00000000} /* (31, 10, 28) {real, imag} */,
  {32'hbe3d2645, 32'h00000000} /* (31, 10, 27) {real, imag} */,
  {32'h3e06243a, 32'h00000000} /* (31, 10, 26) {real, imag} */,
  {32'h3ed3495b, 32'h00000000} /* (31, 10, 25) {real, imag} */,
  {32'h3e4a1044, 32'h00000000} /* (31, 10, 24) {real, imag} */,
  {32'h3ebd9380, 32'h00000000} /* (31, 10, 23) {real, imag} */,
  {32'h3d36b512, 32'h00000000} /* (31, 10, 22) {real, imag} */,
  {32'hbcacfce0, 32'h00000000} /* (31, 10, 21) {real, imag} */,
  {32'h3dc5200e, 32'h00000000} /* (31, 10, 20) {real, imag} */,
  {32'hbe1c7204, 32'h00000000} /* (31, 10, 19) {real, imag} */,
  {32'hbcec3034, 32'h00000000} /* (31, 10, 18) {real, imag} */,
  {32'h3ea13b72, 32'h00000000} /* (31, 10, 17) {real, imag} */,
  {32'hbd4ea600, 32'h00000000} /* (31, 10, 16) {real, imag} */,
  {32'hbf9a048d, 32'h00000000} /* (31, 10, 15) {real, imag} */,
  {32'hbf004f4a, 32'h00000000} /* (31, 10, 14) {real, imag} */,
  {32'hbeddf503, 32'h00000000} /* (31, 10, 13) {real, imag} */,
  {32'h3d32177d, 32'h00000000} /* (31, 10, 12) {real, imag} */,
  {32'h3e83f90d, 32'h00000000} /* (31, 10, 11) {real, imag} */,
  {32'h3e886837, 32'h00000000} /* (31, 10, 10) {real, imag} */,
  {32'h3f03cd59, 32'h00000000} /* (31, 10, 9) {real, imag} */,
  {32'h3f378205, 32'h00000000} /* (31, 10, 8) {real, imag} */,
  {32'h3f28ded4, 32'h00000000} /* (31, 10, 7) {real, imag} */,
  {32'h3ebf8266, 32'h00000000} /* (31, 10, 6) {real, imag} */,
  {32'h3e2eae35, 32'h00000000} /* (31, 10, 5) {real, imag} */,
  {32'h3ede0712, 32'h00000000} /* (31, 10, 4) {real, imag} */,
  {32'h3d219a78, 32'h00000000} /* (31, 10, 3) {real, imag} */,
  {32'h3e310c9b, 32'h00000000} /* (31, 10, 2) {real, imag} */,
  {32'h3e21a31c, 32'h00000000} /* (31, 10, 1) {real, imag} */,
  {32'h3dc6ec69, 32'h00000000} /* (31, 10, 0) {real, imag} */,
  {32'h3f270b78, 32'h00000000} /* (31, 9, 31) {real, imag} */,
  {32'h3f1a8c10, 32'h00000000} /* (31, 9, 30) {real, imag} */,
  {32'h3c9145e2, 32'h00000000} /* (31, 9, 29) {real, imag} */,
  {32'h3d7a1d0c, 32'h00000000} /* (31, 9, 28) {real, imag} */,
  {32'h3e995984, 32'h00000000} /* (31, 9, 27) {real, imag} */,
  {32'h3f20dcf4, 32'h00000000} /* (31, 9, 26) {real, imag} */,
  {32'h3f3b6cc7, 32'h00000000} /* (31, 9, 25) {real, imag} */,
  {32'h3f2b3105, 32'h00000000} /* (31, 9, 24) {real, imag} */,
  {32'h3efd8f95, 32'h00000000} /* (31, 9, 23) {real, imag} */,
  {32'h3f342ebc, 32'h00000000} /* (31, 9, 22) {real, imag} */,
  {32'h3e8b1981, 32'h00000000} /* (31, 9, 21) {real, imag} */,
  {32'hbdc36056, 32'h00000000} /* (31, 9, 20) {real, imag} */,
  {32'hbeab1a24, 32'h00000000} /* (31, 9, 19) {real, imag} */,
  {32'hbedb0fa5, 32'h00000000} /* (31, 9, 18) {real, imag} */,
  {32'hbee67567, 32'h00000000} /* (31, 9, 17) {real, imag} */,
  {32'hbefe74c6, 32'h00000000} /* (31, 9, 16) {real, imag} */,
  {32'hbf4c088e, 32'h00000000} /* (31, 9, 15) {real, imag} */,
  {32'hbef52eb9, 32'h00000000} /* (31, 9, 14) {real, imag} */,
  {32'hbeb8a924, 32'h00000000} /* (31, 9, 13) {real, imag} */,
  {32'hbe4498e7, 32'h00000000} /* (31, 9, 12) {real, imag} */,
  {32'hbd904fe9, 32'h00000000} /* (31, 9, 11) {real, imag} */,
  {32'h3e38ea44, 32'h00000000} /* (31, 9, 10) {real, imag} */,
  {32'h3f5111ce, 32'h00000000} /* (31, 9, 9) {real, imag} */,
  {32'h3f5e2cb1, 32'h00000000} /* (31, 9, 8) {real, imag} */,
  {32'h3f3c9dca, 32'h00000000} /* (31, 9, 7) {real, imag} */,
  {32'h3ea706ce, 32'h00000000} /* (31, 9, 6) {real, imag} */,
  {32'h3ee40692, 32'h00000000} /* (31, 9, 5) {real, imag} */,
  {32'h3f49c795, 32'h00000000} /* (31, 9, 4) {real, imag} */,
  {32'h3efc7520, 32'h00000000} /* (31, 9, 3) {real, imag} */,
  {32'h3ec95cb8, 32'h00000000} /* (31, 9, 2) {real, imag} */,
  {32'h3edab4ba, 32'h00000000} /* (31, 9, 1) {real, imag} */,
  {32'h3e3f136c, 32'h00000000} /* (31, 9, 0) {real, imag} */,
  {32'h3e99884d, 32'h00000000} /* (31, 8, 31) {real, imag} */,
  {32'h3ece32da, 32'h00000000} /* (31, 8, 30) {real, imag} */,
  {32'h3e51f415, 32'h00000000} /* (31, 8, 29) {real, imag} */,
  {32'h3e95f49e, 32'h00000000} /* (31, 8, 28) {real, imag} */,
  {32'h3f350ece, 32'h00000000} /* (31, 8, 27) {real, imag} */,
  {32'h3f627ebb, 32'h00000000} /* (31, 8, 26) {real, imag} */,
  {32'h3f54372b, 32'h00000000} /* (31, 8, 25) {real, imag} */,
  {32'h3f4dc212, 32'h00000000} /* (31, 8, 24) {real, imag} */,
  {32'h3eaaeb88, 32'h00000000} /* (31, 8, 23) {real, imag} */,
  {32'h3e92155c, 32'h00000000} /* (31, 8, 22) {real, imag} */,
  {32'hbc206216, 32'h00000000} /* (31, 8, 21) {real, imag} */,
  {32'hbf29ce16, 32'h00000000} /* (31, 8, 20) {real, imag} */,
  {32'hbec6ec65, 32'h00000000} /* (31, 8, 19) {real, imag} */,
  {32'hbec51700, 32'h00000000} /* (31, 8, 18) {real, imag} */,
  {32'hbf03357a, 32'h00000000} /* (31, 8, 17) {real, imag} */,
  {32'hbe80e434, 32'h00000000} /* (31, 8, 16) {real, imag} */,
  {32'hbe7e4218, 32'h00000000} /* (31, 8, 15) {real, imag} */,
  {32'hbebeefbb, 32'h00000000} /* (31, 8, 14) {real, imag} */,
  {32'hbecf8093, 32'h00000000} /* (31, 8, 13) {real, imag} */,
  {32'hbf45fb52, 32'h00000000} /* (31, 8, 12) {real, imag} */,
  {32'hbf00a5db, 32'h00000000} /* (31, 8, 11) {real, imag} */,
  {32'h3d63400e, 32'h00000000} /* (31, 8, 10) {real, imag} */,
  {32'h3f2b1338, 32'h00000000} /* (31, 8, 9) {real, imag} */,
  {32'h3edf7601, 32'h00000000} /* (31, 8, 8) {real, imag} */,
  {32'h3f374ba2, 32'h00000000} /* (31, 8, 7) {real, imag} */,
  {32'h3ed6c413, 32'h00000000} /* (31, 8, 6) {real, imag} */,
  {32'h3e1e51d4, 32'h00000000} /* (31, 8, 5) {real, imag} */,
  {32'h3ed6fa39, 32'h00000000} /* (31, 8, 4) {real, imag} */,
  {32'h3ee533c5, 32'h00000000} /* (31, 8, 3) {real, imag} */,
  {32'h3e9b094b, 32'h00000000} /* (31, 8, 2) {real, imag} */,
  {32'h3ec59ed5, 32'h00000000} /* (31, 8, 1) {real, imag} */,
  {32'h3e82e64c, 32'h00000000} /* (31, 8, 0) {real, imag} */,
  {32'h3f197efb, 32'h00000000} /* (31, 7, 31) {real, imag} */,
  {32'h3ef49de3, 32'h00000000} /* (31, 7, 30) {real, imag} */,
  {32'h3eb9c0dc, 32'h00000000} /* (31, 7, 29) {real, imag} */,
  {32'h3ed7a9df, 32'h00000000} /* (31, 7, 28) {real, imag} */,
  {32'h3ed8d4e2, 32'h00000000} /* (31, 7, 27) {real, imag} */,
  {32'h3e85b280, 32'h00000000} /* (31, 7, 26) {real, imag} */,
  {32'h3eb943fa, 32'h00000000} /* (31, 7, 25) {real, imag} */,
  {32'h3ebf5e38, 32'h00000000} /* (31, 7, 24) {real, imag} */,
  {32'h3eab738c, 32'h00000000} /* (31, 7, 23) {real, imag} */,
  {32'h3e858dd4, 32'h00000000} /* (31, 7, 22) {real, imag} */,
  {32'hbed7ab5c, 32'h00000000} /* (31, 7, 21) {real, imag} */,
  {32'hbf822f5e, 32'h00000000} /* (31, 7, 20) {real, imag} */,
  {32'hbe0929ad, 32'h00000000} /* (31, 7, 19) {real, imag} */,
  {32'hbd61dde3, 32'h00000000} /* (31, 7, 18) {real, imag} */,
  {32'hbe50dd8c, 32'h00000000} /* (31, 7, 17) {real, imag} */,
  {32'hbe1dda26, 32'h00000000} /* (31, 7, 16) {real, imag} */,
  {32'hbea37d45, 32'h00000000} /* (31, 7, 15) {real, imag} */,
  {32'hbeb4d546, 32'h00000000} /* (31, 7, 14) {real, imag} */,
  {32'hbe6c7ea0, 32'h00000000} /* (31, 7, 13) {real, imag} */,
  {32'hbf030bec, 32'h00000000} /* (31, 7, 12) {real, imag} */,
  {32'hbf3e8fb3, 32'h00000000} /* (31, 7, 11) {real, imag} */,
  {32'h3e8b6093, 32'h00000000} /* (31, 7, 10) {real, imag} */,
  {32'h3f216ce8, 32'h00000000} /* (31, 7, 9) {real, imag} */,
  {32'h3f0fe1a6, 32'h00000000} /* (31, 7, 8) {real, imag} */,
  {32'h3f958a28, 32'h00000000} /* (31, 7, 7) {real, imag} */,
  {32'h3f21a198, 32'h00000000} /* (31, 7, 6) {real, imag} */,
  {32'h3ec68eea, 32'h00000000} /* (31, 7, 5) {real, imag} */,
  {32'h3ec73959, 32'h00000000} /* (31, 7, 4) {real, imag} */,
  {32'h3f06a38a, 32'h00000000} /* (31, 7, 3) {real, imag} */,
  {32'h3ed058db, 32'h00000000} /* (31, 7, 2) {real, imag} */,
  {32'h3e8329cc, 32'h00000000} /* (31, 7, 1) {real, imag} */,
  {32'h3e8ea1f6, 32'h00000000} /* (31, 7, 0) {real, imag} */,
  {32'h3f1d753b, 32'h00000000} /* (31, 6, 31) {real, imag} */,
  {32'h3eb12314, 32'h00000000} /* (31, 6, 30) {real, imag} */,
  {32'h3eeaaec7, 32'h00000000} /* (31, 6, 29) {real, imag} */,
  {32'h3eeec0ca, 32'h00000000} /* (31, 6, 28) {real, imag} */,
  {32'h3d9783cc, 32'h00000000} /* (31, 6, 27) {real, imag} */,
  {32'h3cbeb6bb, 32'h00000000} /* (31, 6, 26) {real, imag} */,
  {32'h3e7c9463, 32'h00000000} /* (31, 6, 25) {real, imag} */,
  {32'h3ecda8a4, 32'h00000000} /* (31, 6, 24) {real, imag} */,
  {32'h3ed3d2a3, 32'h00000000} /* (31, 6, 23) {real, imag} */,
  {32'h3ee8bdf7, 32'h00000000} /* (31, 6, 22) {real, imag} */,
  {32'h3d3be160, 32'h00000000} /* (31, 6, 21) {real, imag} */,
  {32'hbf11af75, 32'h00000000} /* (31, 6, 20) {real, imag} */,
  {32'hbe3643be, 32'h00000000} /* (31, 6, 19) {real, imag} */,
  {32'hbec5ea3a, 32'h00000000} /* (31, 6, 18) {real, imag} */,
  {32'hbf5bcbb9, 32'h00000000} /* (31, 6, 17) {real, imag} */,
  {32'hbe9e51d8, 32'h00000000} /* (31, 6, 16) {real, imag} */,
  {32'hbe106ba8, 32'h00000000} /* (31, 6, 15) {real, imag} */,
  {32'hbee0ff67, 32'h00000000} /* (31, 6, 14) {real, imag} */,
  {32'hbee3193c, 32'h00000000} /* (31, 6, 13) {real, imag} */,
  {32'hbe49987a, 32'h00000000} /* (31, 6, 12) {real, imag} */,
  {32'hbf0304e4, 32'h00000000} /* (31, 6, 11) {real, imag} */,
  {32'h3d93215d, 32'h00000000} /* (31, 6, 10) {real, imag} */,
  {32'h3e98316e, 32'h00000000} /* (31, 6, 9) {real, imag} */,
  {32'h3ebec01b, 32'h00000000} /* (31, 6, 8) {real, imag} */,
  {32'h3f99d66b, 32'h00000000} /* (31, 6, 7) {real, imag} */,
  {32'h3f83254d, 32'h00000000} /* (31, 6, 6) {real, imag} */,
  {32'h3ef8cf06, 32'h00000000} /* (31, 6, 5) {real, imag} */,
  {32'h3ec69b88, 32'h00000000} /* (31, 6, 4) {real, imag} */,
  {32'h3efc881e, 32'h00000000} /* (31, 6, 3) {real, imag} */,
  {32'h3ed7466c, 32'h00000000} /* (31, 6, 2) {real, imag} */,
  {32'h3f1a0518, 32'h00000000} /* (31, 6, 1) {real, imag} */,
  {32'h3e800284, 32'h00000000} /* (31, 6, 0) {real, imag} */,
  {32'h3ed4450e, 32'h00000000} /* (31, 5, 31) {real, imag} */,
  {32'h3e4e3492, 32'h00000000} /* (31, 5, 30) {real, imag} */,
  {32'h3f29c67b, 32'h00000000} /* (31, 5, 29) {real, imag} */,
  {32'h3f7d6148, 32'h00000000} /* (31, 5, 28) {real, imag} */,
  {32'h3e3ec09e, 32'h00000000} /* (31, 5, 27) {real, imag} */,
  {32'h3eef4ffe, 32'h00000000} /* (31, 5, 26) {real, imag} */,
  {32'h3e666b72, 32'h00000000} /* (31, 5, 25) {real, imag} */,
  {32'h3ebf3cd9, 32'h00000000} /* (31, 5, 24) {real, imag} */,
  {32'h3f001758, 32'h00000000} /* (31, 5, 23) {real, imag} */,
  {32'h3eee95ee, 32'h00000000} /* (31, 5, 22) {real, imag} */,
  {32'h3ecc56fc, 32'h00000000} /* (31, 5, 21) {real, imag} */,
  {32'h3c85bcc8, 32'h00000000} /* (31, 5, 20) {real, imag} */,
  {32'h3e142752, 32'h00000000} /* (31, 5, 19) {real, imag} */,
  {32'h3cb53614, 32'h00000000} /* (31, 5, 18) {real, imag} */,
  {32'hbee7f25d, 32'h00000000} /* (31, 5, 17) {real, imag} */,
  {32'hbe13a7da, 32'h00000000} /* (31, 5, 16) {real, imag} */,
  {32'hbe1f31d7, 32'h00000000} /* (31, 5, 15) {real, imag} */,
  {32'hbeb210ba, 32'h00000000} /* (31, 5, 14) {real, imag} */,
  {32'hbef5ab44, 32'h00000000} /* (31, 5, 13) {real, imag} */,
  {32'hbe523c6a, 32'h00000000} /* (31, 5, 12) {real, imag} */,
  {32'hbef5306b, 32'h00000000} /* (31, 5, 11) {real, imag} */,
  {32'hbedd7f0f, 32'h00000000} /* (31, 5, 10) {real, imag} */,
  {32'hbe82c11a, 32'h00000000} /* (31, 5, 9) {real, imag} */,
  {32'hbe20c51c, 32'h00000000} /* (31, 5, 8) {real, imag} */,
  {32'h3e729eda, 32'h00000000} /* (31, 5, 7) {real, imag} */,
  {32'h3e9c3ec0, 32'h00000000} /* (31, 5, 6) {real, imag} */,
  {32'h3e69dee1, 32'h00000000} /* (31, 5, 5) {real, imag} */,
  {32'h3f0ff326, 32'h00000000} /* (31, 5, 4) {real, imag} */,
  {32'h3ec74dc2, 32'h00000000} /* (31, 5, 3) {real, imag} */,
  {32'h3e74c365, 32'h00000000} /* (31, 5, 2) {real, imag} */,
  {32'h3ed08766, 32'h00000000} /* (31, 5, 1) {real, imag} */,
  {32'h3dd9f363, 32'h00000000} /* (31, 5, 0) {real, imag} */,
  {32'h3e1b46fd, 32'h00000000} /* (31, 4, 31) {real, imag} */,
  {32'hbd9a998a, 32'h00000000} /* (31, 4, 30) {real, imag} */,
  {32'h3c87967f, 32'h00000000} /* (31, 4, 29) {real, imag} */,
  {32'h3f12b317, 32'h00000000} /* (31, 4, 28) {real, imag} */,
  {32'h3f037ea7, 32'h00000000} /* (31, 4, 27) {real, imag} */,
  {32'h3f21d355, 32'h00000000} /* (31, 4, 26) {real, imag} */,
  {32'h3e9828c0, 32'h00000000} /* (31, 4, 25) {real, imag} */,
  {32'h3e1dbef8, 32'h00000000} /* (31, 4, 24) {real, imag} */,
  {32'h3e573e5d, 32'h00000000} /* (31, 4, 23) {real, imag} */,
  {32'h3e906eab, 32'h00000000} /* (31, 4, 22) {real, imag} */,
  {32'h3e870c65, 32'h00000000} /* (31, 4, 21) {real, imag} */,
  {32'h3e5d1d6d, 32'h00000000} /* (31, 4, 20) {real, imag} */,
  {32'h3e98c000, 32'h00000000} /* (31, 4, 19) {real, imag} */,
  {32'h3e9a5cd9, 32'h00000000} /* (31, 4, 18) {real, imag} */,
  {32'h3ea8a82b, 32'h00000000} /* (31, 4, 17) {real, imag} */,
  {32'h3de8fa2a, 32'h00000000} /* (31, 4, 16) {real, imag} */,
  {32'hbe6d2a26, 32'h00000000} /* (31, 4, 15) {real, imag} */,
  {32'hbe269970, 32'h00000000} /* (31, 4, 14) {real, imag} */,
  {32'hbe92cbe1, 32'h00000000} /* (31, 4, 13) {real, imag} */,
  {32'hbe9751eb, 32'h00000000} /* (31, 4, 12) {real, imag} */,
  {32'hbf58a29c, 32'h00000000} /* (31, 4, 11) {real, imag} */,
  {32'hbf7c4dfe, 32'h00000000} /* (31, 4, 10) {real, imag} */,
  {32'hbeb4671f, 32'h00000000} /* (31, 4, 9) {real, imag} */,
  {32'hbe2b12f5, 32'h00000000} /* (31, 4, 8) {real, imag} */,
  {32'hbe0a540e, 32'h00000000} /* (31, 4, 7) {real, imag} */,
  {32'hbe3d4436, 32'h00000000} /* (31, 4, 6) {real, imag} */,
  {32'h3e1f2a10, 32'h00000000} /* (31, 4, 5) {real, imag} */,
  {32'h3eb4b36a, 32'h00000000} /* (31, 4, 4) {real, imag} */,
  {32'h3e7f1212, 32'h00000000} /* (31, 4, 3) {real, imag} */,
  {32'h3ea255a2, 32'h00000000} /* (31, 4, 2) {real, imag} */,
  {32'h3f00cd08, 32'h00000000} /* (31, 4, 1) {real, imag} */,
  {32'h3eb9163b, 32'h00000000} /* (31, 4, 0) {real, imag} */,
  {32'h3e9de6dd, 32'h00000000} /* (31, 3, 31) {real, imag} */,
  {32'h3ef96ab7, 32'h00000000} /* (31, 3, 30) {real, imag} */,
  {32'h3ec6cca0, 32'h00000000} /* (31, 3, 29) {real, imag} */,
  {32'h3ed8b827, 32'h00000000} /* (31, 3, 28) {real, imag} */,
  {32'h3f1575b5, 32'h00000000} /* (31, 3, 27) {real, imag} */,
  {32'h3f420d03, 32'h00000000} /* (31, 3, 26) {real, imag} */,
  {32'h3f0939b4, 32'h00000000} /* (31, 3, 25) {real, imag} */,
  {32'h3ef280a9, 32'h00000000} /* (31, 3, 24) {real, imag} */,
  {32'h3ee7bb27, 32'h00000000} /* (31, 3, 23) {real, imag} */,
  {32'h3edd8266, 32'h00000000} /* (31, 3, 22) {real, imag} */,
  {32'h3ea23e5f, 32'h00000000} /* (31, 3, 21) {real, imag} */,
  {32'h3ea0f425, 32'h00000000} /* (31, 3, 20) {real, imag} */,
  {32'h3eaf01c0, 32'h00000000} /* (31, 3, 19) {real, imag} */,
  {32'h3dd63c18, 32'h00000000} /* (31, 3, 18) {real, imag} */,
  {32'h3e942c20, 32'h00000000} /* (31, 3, 17) {real, imag} */,
  {32'h3d616e9d, 32'h00000000} /* (31, 3, 16) {real, imag} */,
  {32'hbed1d4d4, 32'h00000000} /* (31, 3, 15) {real, imag} */,
  {32'hbf11f6f2, 32'h00000000} /* (31, 3, 14) {real, imag} */,
  {32'hbf1c3622, 32'h00000000} /* (31, 3, 13) {real, imag} */,
  {32'hbf31bb9f, 32'h00000000} /* (31, 3, 12) {real, imag} */,
  {32'hbf51451a, 32'h00000000} /* (31, 3, 11) {real, imag} */,
  {32'hbf92c26c, 32'h00000000} /* (31, 3, 10) {real, imag} */,
  {32'hbedd9f62, 32'h00000000} /* (31, 3, 9) {real, imag} */,
  {32'hbe857c61, 32'h00000000} /* (31, 3, 8) {real, imag} */,
  {32'hbeeb2001, 32'h00000000} /* (31, 3, 7) {real, imag} */,
  {32'hbf03c26d, 32'h00000000} /* (31, 3, 6) {real, imag} */,
  {32'hbea40ce6, 32'h00000000} /* (31, 3, 5) {real, imag} */,
  {32'h3e4eacc4, 32'h00000000} /* (31, 3, 4) {real, imag} */,
  {32'h3ec93cfc, 32'h00000000} /* (31, 3, 3) {real, imag} */,
  {32'h3f2b6fe9, 32'h00000000} /* (31, 3, 2) {real, imag} */,
  {32'h3f376bb0, 32'h00000000} /* (31, 3, 1) {real, imag} */,
  {32'h3eac816c, 32'h00000000} /* (31, 3, 0) {real, imag} */,
  {32'h3e6cf57b, 32'h00000000} /* (31, 2, 31) {real, imag} */,
  {32'h3f1c2430, 32'h00000000} /* (31, 2, 30) {real, imag} */,
  {32'h3f0a7c7c, 32'h00000000} /* (31, 2, 29) {real, imag} */,
  {32'h3eb07287, 32'h00000000} /* (31, 2, 28) {real, imag} */,
  {32'h3f1ac5c6, 32'h00000000} /* (31, 2, 27) {real, imag} */,
  {32'h3f29f990, 32'h00000000} /* (31, 2, 26) {real, imag} */,
  {32'h3e8ea6b7, 32'h00000000} /* (31, 2, 25) {real, imag} */,
  {32'h3ec98ca1, 32'h00000000} /* (31, 2, 24) {real, imag} */,
  {32'h3e415498, 32'h00000000} /* (31, 2, 23) {real, imag} */,
  {32'h3e14012e, 32'h00000000} /* (31, 2, 22) {real, imag} */,
  {32'h3ea40aed, 32'h00000000} /* (31, 2, 21) {real, imag} */,
  {32'h3ee4e947, 32'h00000000} /* (31, 2, 20) {real, imag} */,
  {32'h3ea03925, 32'h00000000} /* (31, 2, 19) {real, imag} */,
  {32'hbda4d6b8, 32'h00000000} /* (31, 2, 18) {real, imag} */,
  {32'h3a9cb040, 32'h00000000} /* (31, 2, 17) {real, imag} */,
  {32'hbe17a6ba, 32'h00000000} /* (31, 2, 16) {real, imag} */,
  {32'hbf333a7e, 32'h00000000} /* (31, 2, 15) {real, imag} */,
  {32'hbeecefd6, 32'h00000000} /* (31, 2, 14) {real, imag} */,
  {32'hbedd2ace, 32'h00000000} /* (31, 2, 13) {real, imag} */,
  {32'hbf35f414, 32'h00000000} /* (31, 2, 12) {real, imag} */,
  {32'hbf101046, 32'h00000000} /* (31, 2, 11) {real, imag} */,
  {32'hbf22765d, 32'h00000000} /* (31, 2, 10) {real, imag} */,
  {32'hbf0b9957, 32'h00000000} /* (31, 2, 9) {real, imag} */,
  {32'hbeca9f48, 32'h00000000} /* (31, 2, 8) {real, imag} */,
  {32'hbf55ba4f, 32'h00000000} /* (31, 2, 7) {real, imag} */,
  {32'hbf6d3320, 32'h00000000} /* (31, 2, 6) {real, imag} */,
  {32'hbebad608, 32'h00000000} /* (31, 2, 5) {real, imag} */,
  {32'h3e40f7b4, 32'h00000000} /* (31, 2, 4) {real, imag} */,
  {32'h3f1f86c3, 32'h00000000} /* (31, 2, 3) {real, imag} */,
  {32'h3ef78870, 32'h00000000} /* (31, 2, 2) {real, imag} */,
  {32'h3e9a2ff3, 32'h00000000} /* (31, 2, 1) {real, imag} */,
  {32'h3e1b4bd7, 32'h00000000} /* (31, 2, 0) {real, imag} */,
  {32'h3e2b8708, 32'h00000000} /* (31, 1, 31) {real, imag} */,
  {32'h3ead05ea, 32'h00000000} /* (31, 1, 30) {real, imag} */,
  {32'h3ddfb74e, 32'h00000000} /* (31, 1, 29) {real, imag} */,
  {32'h3e87aaca, 32'h00000000} /* (31, 1, 28) {real, imag} */,
  {32'h3f1138c4, 32'h00000000} /* (31, 1, 27) {real, imag} */,
  {32'h3ec3d478, 32'h00000000} /* (31, 1, 26) {real, imag} */,
  {32'h3eca1bdb, 32'h00000000} /* (31, 1, 25) {real, imag} */,
  {32'h3f2c22c9, 32'h00000000} /* (31, 1, 24) {real, imag} */,
  {32'h3e6a3184, 32'h00000000} /* (31, 1, 23) {real, imag} */,
  {32'h3e42d15b, 32'h00000000} /* (31, 1, 22) {real, imag} */,
  {32'h3e46df2f, 32'h00000000} /* (31, 1, 21) {real, imag} */,
  {32'h3e86a8fc, 32'h00000000} /* (31, 1, 20) {real, imag} */,
  {32'h3e7b8723, 32'h00000000} /* (31, 1, 19) {real, imag} */,
  {32'h3d03bd6e, 32'h00000000} /* (31, 1, 18) {real, imag} */,
  {32'h3e131ca1, 32'h00000000} /* (31, 1, 17) {real, imag} */,
  {32'hbe0e342f, 32'h00000000} /* (31, 1, 16) {real, imag} */,
  {32'hbef3de5e, 32'h00000000} /* (31, 1, 15) {real, imag} */,
  {32'hbe912210, 32'h00000000} /* (31, 1, 14) {real, imag} */,
  {32'h3d9cbe97, 32'h00000000} /* (31, 1, 13) {real, imag} */,
  {32'hbdee08b2, 32'h00000000} /* (31, 1, 12) {real, imag} */,
  {32'hbed8a34c, 32'h00000000} /* (31, 1, 11) {real, imag} */,
  {32'hbf473643, 32'h00000000} /* (31, 1, 10) {real, imag} */,
  {32'hbf0c4433, 32'h00000000} /* (31, 1, 9) {real, imag} */,
  {32'hbebb3da0, 32'h00000000} /* (31, 1, 8) {real, imag} */,
  {32'hbedbb374, 32'h00000000} /* (31, 1, 7) {real, imag} */,
  {32'hbf1d5442, 32'h00000000} /* (31, 1, 6) {real, imag} */,
  {32'hbd3506dd, 32'h00000000} /* (31, 1, 5) {real, imag} */,
  {32'h3e92e930, 32'h00000000} /* (31, 1, 4) {real, imag} */,
  {32'h3ec486b1, 32'h00000000} /* (31, 1, 3) {real, imag} */,
  {32'h3ea05fd0, 32'h00000000} /* (31, 1, 2) {real, imag} */,
  {32'h3d4b839b, 32'h00000000} /* (31, 1, 1) {real, imag} */,
  {32'h3becadae, 32'h00000000} /* (31, 1, 0) {real, imag} */,
  {32'h3de1a70a, 32'h00000000} /* (31, 0, 31) {real, imag} */,
  {32'h3d485e44, 32'h00000000} /* (31, 0, 30) {real, imag} */,
  {32'hbdb38b8e, 32'h00000000} /* (31, 0, 29) {real, imag} */,
  {32'h3da267a8, 32'h00000000} /* (31, 0, 28) {real, imag} */,
  {32'h3e144c58, 32'h00000000} /* (31, 0, 27) {real, imag} */,
  {32'h3e1e0fd9, 32'h00000000} /* (31, 0, 26) {real, imag} */,
  {32'h3eb590f2, 32'h00000000} /* (31, 0, 25) {real, imag} */,
  {32'h3e968d11, 32'h00000000} /* (31, 0, 24) {real, imag} */,
  {32'h3e8eaf1c, 32'h00000000} /* (31, 0, 23) {real, imag} */,
  {32'h3ea6be84, 32'h00000000} /* (31, 0, 22) {real, imag} */,
  {32'h3e4a7b24, 32'h00000000} /* (31, 0, 21) {real, imag} */,
  {32'h3d931f4c, 32'h00000000} /* (31, 0, 20) {real, imag} */,
  {32'h3e19e6df, 32'h00000000} /* (31, 0, 19) {real, imag} */,
  {32'h3d4c1983, 32'h00000000} /* (31, 0, 18) {real, imag} */,
  {32'h3e023725, 32'h00000000} /* (31, 0, 17) {real, imag} */,
  {32'hbd825fe5, 32'h00000000} /* (31, 0, 16) {real, imag} */,
  {32'hbeb44129, 32'h00000000} /* (31, 0, 15) {real, imag} */,
  {32'hbefe9d21, 32'h00000000} /* (31, 0, 14) {real, imag} */,
  {32'hbe8561a2, 32'h00000000} /* (31, 0, 13) {real, imag} */,
  {32'hbcf0f43f, 32'h00000000} /* (31, 0, 12) {real, imag} */,
  {32'hbde8a584, 32'h00000000} /* (31, 0, 11) {real, imag} */,
  {32'hbee9ca15, 32'h00000000} /* (31, 0, 10) {real, imag} */,
  {32'hbe297364, 32'h00000000} /* (31, 0, 9) {real, imag} */,
  {32'hbe22d470, 32'h00000000} /* (31, 0, 8) {real, imag} */,
  {32'hbe360ac3, 32'h00000000} /* (31, 0, 7) {real, imag} */,
  {32'hbd880fa0, 32'h00000000} /* (31, 0, 6) {real, imag} */,
  {32'h3e2bb326, 32'h00000000} /* (31, 0, 5) {real, imag} */,
  {32'h3e84d996, 32'h00000000} /* (31, 0, 4) {real, imag} */,
  {32'h3d9d9d39, 32'h00000000} /* (31, 0, 3) {real, imag} */,
  {32'h3d98a688, 32'h00000000} /* (31, 0, 2) {real, imag} */,
  {32'h3c6d20c3, 32'h00000000} /* (31, 0, 1) {real, imag} */,
  {32'h3c899e25, 32'h00000000} /* (31, 0, 0) {real, imag} */,
  {32'h3e8d3a31, 32'h00000000} /* (30, 31, 31) {real, imag} */,
  {32'h3ed1ae24, 32'h00000000} /* (30, 31, 30) {real, imag} */,
  {32'h3f367a7d, 32'h00000000} /* (30, 31, 29) {real, imag} */,
  {32'h3eeca277, 32'h00000000} /* (30, 31, 28) {real, imag} */,
  {32'h3ea5a87f, 32'h00000000} /* (30, 31, 27) {real, imag} */,
  {32'h3e9e940c, 32'h00000000} /* (30, 31, 26) {real, imag} */,
  {32'h3f870f74, 32'h00000000} /* (30, 31, 25) {real, imag} */,
  {32'h3f2cdfdd, 32'h00000000} /* (30, 31, 24) {real, imag} */,
  {32'h3e830eb5, 32'h00000000} /* (30, 31, 23) {real, imag} */,
  {32'h3eb5a654, 32'h00000000} /* (30, 31, 22) {real, imag} */,
  {32'h3f0d9a8e, 32'h00000000} /* (30, 31, 21) {real, imag} */,
  {32'hbd9b18dd, 32'h00000000} /* (30, 31, 20) {real, imag} */,
  {32'hbe3883e3, 32'h00000000} /* (30, 31, 19) {real, imag} */,
  {32'hbe0be425, 32'h00000000} /* (30, 31, 18) {real, imag} */,
  {32'hbe26144e, 32'h00000000} /* (30, 31, 17) {real, imag} */,
  {32'hbedda31f, 32'h00000000} /* (30, 31, 16) {real, imag} */,
  {32'hbeafb9b5, 32'h00000000} /* (30, 31, 15) {real, imag} */,
  {32'hbf2909fa, 32'h00000000} /* (30, 31, 14) {real, imag} */,
  {32'hbf6cc036, 32'h00000000} /* (30, 31, 13) {real, imag} */,
  {32'hbf40d1be, 32'h00000000} /* (30, 31, 12) {real, imag} */,
  {32'hbf0cc790, 32'h00000000} /* (30, 31, 11) {real, imag} */,
  {32'hbce00a8b, 32'h00000000} /* (30, 31, 10) {real, imag} */,
  {32'h3ed2efeb, 32'h00000000} /* (30, 31, 9) {real, imag} */,
  {32'h3ec5928e, 32'h00000000} /* (30, 31, 8) {real, imag} */,
  {32'h3da5a992, 32'h00000000} /* (30, 31, 7) {real, imag} */,
  {32'h3e83e598, 32'h00000000} /* (30, 31, 6) {real, imag} */,
  {32'h3ed7a347, 32'h00000000} /* (30, 31, 5) {real, imag} */,
  {32'h3ef6e6c3, 32'h00000000} /* (30, 31, 4) {real, imag} */,
  {32'h3ec9913a, 32'h00000000} /* (30, 31, 3) {real, imag} */,
  {32'h3f06af8a, 32'h00000000} /* (30, 31, 2) {real, imag} */,
  {32'h3f1d030c, 32'h00000000} /* (30, 31, 1) {real, imag} */,
  {32'h3edd4095, 32'h00000000} /* (30, 31, 0) {real, imag} */,
  {32'h3f13b97e, 32'h00000000} /* (30, 30, 31) {real, imag} */,
  {32'h3f6d7400, 32'h00000000} /* (30, 30, 30) {real, imag} */,
  {32'h3f85b29e, 32'h00000000} /* (30, 30, 29) {real, imag} */,
  {32'h3f371dd4, 32'h00000000} /* (30, 30, 28) {real, imag} */,
  {32'h3f363493, 32'h00000000} /* (30, 30, 27) {real, imag} */,
  {32'h3f6393bb, 32'h00000000} /* (30, 30, 26) {real, imag} */,
  {32'h3fd452bc, 32'h00000000} /* (30, 30, 25) {real, imag} */,
  {32'h3fbaecf5, 32'h00000000} /* (30, 30, 24) {real, imag} */,
  {32'h3f9243c6, 32'h00000000} /* (30, 30, 23) {real, imag} */,
  {32'h3f721c4b, 32'h00000000} /* (30, 30, 22) {real, imag} */,
  {32'h3f967a8a, 32'h00000000} /* (30, 30, 21) {real, imag} */,
  {32'h3e0c56aa, 32'h00000000} /* (30, 30, 20) {real, imag} */,
  {32'hbea1a202, 32'h00000000} /* (30, 30, 19) {real, imag} */,
  {32'hbf1638fe, 32'h00000000} /* (30, 30, 18) {real, imag} */,
  {32'hbf2b3afe, 32'h00000000} /* (30, 30, 17) {real, imag} */,
  {32'hbf2f29c1, 32'h00000000} /* (30, 30, 16) {real, imag} */,
  {32'hbf4f5622, 32'h00000000} /* (30, 30, 15) {real, imag} */,
  {32'hbfb07f3e, 32'h00000000} /* (30, 30, 14) {real, imag} */,
  {32'hbffca469, 32'h00000000} /* (30, 30, 13) {real, imag} */,
  {32'hbfc965cb, 32'h00000000} /* (30, 30, 12) {real, imag} */,
  {32'hbf51beea, 32'h00000000} /* (30, 30, 11) {real, imag} */,
  {32'h3c24ab96, 32'h00000000} /* (30, 30, 10) {real, imag} */,
  {32'h3f5e96fd, 32'h00000000} /* (30, 30, 9) {real, imag} */,
  {32'h3f4e2184, 32'h00000000} /* (30, 30, 8) {real, imag} */,
  {32'h3ead4137, 32'h00000000} /* (30, 30, 7) {real, imag} */,
  {32'h3f1c5893, 32'h00000000} /* (30, 30, 6) {real, imag} */,
  {32'h3f7236c4, 32'h00000000} /* (30, 30, 5) {real, imag} */,
  {32'h3f9c49ee, 32'h00000000} /* (30, 30, 4) {real, imag} */,
  {32'h3f89bf33, 32'h00000000} /* (30, 30, 3) {real, imag} */,
  {32'h3f4d344a, 32'h00000000} /* (30, 30, 2) {real, imag} */,
  {32'h3faae7f8, 32'h00000000} /* (30, 30, 1) {real, imag} */,
  {32'h3f89491d, 32'h00000000} /* (30, 30, 0) {real, imag} */,
  {32'h3f0343ae, 32'h00000000} /* (30, 29, 31) {real, imag} */,
  {32'h3f9a475e, 32'h00000000} /* (30, 29, 30) {real, imag} */,
  {32'h3f9b3ff5, 32'h00000000} /* (30, 29, 29) {real, imag} */,
  {32'h3f0a3219, 32'h00000000} /* (30, 29, 28) {real, imag} */,
  {32'h3eca259f, 32'h00000000} /* (30, 29, 27) {real, imag} */,
  {32'h3f11ff52, 32'h00000000} /* (30, 29, 26) {real, imag} */,
  {32'h3f88c82f, 32'h00000000} /* (30, 29, 25) {real, imag} */,
  {32'h3fa9f218, 32'h00000000} /* (30, 29, 24) {real, imag} */,
  {32'h3f914992, 32'h00000000} /* (30, 29, 23) {real, imag} */,
  {32'h3f7558ef, 32'h00000000} /* (30, 29, 22) {real, imag} */,
  {32'h3ea6e832, 32'h00000000} /* (30, 29, 21) {real, imag} */,
  {32'hbf6224d9, 32'h00000000} /* (30, 29, 20) {real, imag} */,
  {32'hbf0aa84e, 32'h00000000} /* (30, 29, 19) {real, imag} */,
  {32'hbf1de3a5, 32'h00000000} /* (30, 29, 18) {real, imag} */,
  {32'hbf797c29, 32'h00000000} /* (30, 29, 17) {real, imag} */,
  {32'hbf95ee2c, 32'h00000000} /* (30, 29, 16) {real, imag} */,
  {32'hbf7a07d0, 32'h00000000} /* (30, 29, 15) {real, imag} */,
  {32'hbfb427db, 32'h00000000} /* (30, 29, 14) {real, imag} */,
  {32'hbfbf182c, 32'h00000000} /* (30, 29, 13) {real, imag} */,
  {32'hbf8aa186, 32'h00000000} /* (30, 29, 12) {real, imag} */,
  {32'hbf673e1c, 32'h00000000} /* (30, 29, 11) {real, imag} */,
  {32'hbe5f6775, 32'h00000000} /* (30, 29, 10) {real, imag} */,
  {32'h3f48cf1c, 32'h00000000} /* (30, 29, 9) {real, imag} */,
  {32'h3f421187, 32'h00000000} /* (30, 29, 8) {real, imag} */,
  {32'h3e8a9470, 32'h00000000} /* (30, 29, 7) {real, imag} */,
  {32'h3f11c10d, 32'h00000000} /* (30, 29, 6) {real, imag} */,
  {32'h3f7e25fc, 32'h00000000} /* (30, 29, 5) {real, imag} */,
  {32'h3f8a398f, 32'h00000000} /* (30, 29, 4) {real, imag} */,
  {32'h3fa44a31, 32'h00000000} /* (30, 29, 3) {real, imag} */,
  {32'h3f36c3f2, 32'h00000000} /* (30, 29, 2) {real, imag} */,
  {32'h3f2af15a, 32'h00000000} /* (30, 29, 1) {real, imag} */,
  {32'h3f12e894, 32'h00000000} /* (30, 29, 0) {real, imag} */,
  {32'h3ef4cd97, 32'h00000000} /* (30, 28, 31) {real, imag} */,
  {32'h3fcc9654, 32'h00000000} /* (30, 28, 30) {real, imag} */,
  {32'h3fee22f7, 32'h00000000} /* (30, 28, 29) {real, imag} */,
  {32'h3f2de866, 32'h00000000} /* (30, 28, 28) {real, imag} */,
  {32'h3f226e01, 32'h00000000} /* (30, 28, 27) {real, imag} */,
  {32'h3fa6c440, 32'h00000000} /* (30, 28, 26) {real, imag} */,
  {32'h3f8a9878, 32'h00000000} /* (30, 28, 25) {real, imag} */,
  {32'h3f39e3df, 32'h00000000} /* (30, 28, 24) {real, imag} */,
  {32'h3ed956a2, 32'h00000000} /* (30, 28, 23) {real, imag} */,
  {32'h3ed3ea4b, 32'h00000000} /* (30, 28, 22) {real, imag} */,
  {32'h3c8ad7ae, 32'h00000000} /* (30, 28, 21) {real, imag} */,
  {32'hbf91d55b, 32'h00000000} /* (30, 28, 20) {real, imag} */,
  {32'hbf85a093, 32'h00000000} /* (30, 28, 19) {real, imag} */,
  {32'hbf375a2c, 32'h00000000} /* (30, 28, 18) {real, imag} */,
  {32'hbf0fe9fa, 32'h00000000} /* (30, 28, 17) {real, imag} */,
  {32'hbf042f82, 32'h00000000} /* (30, 28, 16) {real, imag} */,
  {32'hbf11439b, 32'h00000000} /* (30, 28, 15) {real, imag} */,
  {32'hbf899a69, 32'h00000000} /* (30, 28, 14) {real, imag} */,
  {32'hbf856653, 32'h00000000} /* (30, 28, 13) {real, imag} */,
  {32'hbee13404, 32'h00000000} /* (30, 28, 12) {real, imag} */,
  {32'hbf23b455, 32'h00000000} /* (30, 28, 11) {real, imag} */,
  {32'h3e20c16c, 32'h00000000} /* (30, 28, 10) {real, imag} */,
  {32'h3f27b001, 32'h00000000} /* (30, 28, 9) {real, imag} */,
  {32'h3f7683b7, 32'h00000000} /* (30, 28, 8) {real, imag} */,
  {32'h3f2a3b22, 32'h00000000} /* (30, 28, 7) {real, imag} */,
  {32'h3f4bb325, 32'h00000000} /* (30, 28, 6) {real, imag} */,
  {32'h3f17f876, 32'h00000000} /* (30, 28, 5) {real, imag} */,
  {32'h3f1ec893, 32'h00000000} /* (30, 28, 4) {real, imag} */,
  {32'h3f4eebae, 32'h00000000} /* (30, 28, 3) {real, imag} */,
  {32'h3f1a6b78, 32'h00000000} /* (30, 28, 2) {real, imag} */,
  {32'h3f0334b8, 32'h00000000} /* (30, 28, 1) {real, imag} */,
  {32'h3ee6137e, 32'h00000000} /* (30, 28, 0) {real, imag} */,
  {32'h3f59482c, 32'h00000000} /* (30, 27, 31) {real, imag} */,
  {32'h3f9d8f39, 32'h00000000} /* (30, 27, 30) {real, imag} */,
  {32'h3f8a8bf1, 32'h00000000} /* (30, 27, 29) {real, imag} */,
  {32'h3f008c34, 32'h00000000} /* (30, 27, 28) {real, imag} */,
  {32'h3f84eacd, 32'h00000000} /* (30, 27, 27) {real, imag} */,
  {32'h3fe909df, 32'h00000000} /* (30, 27, 26) {real, imag} */,
  {32'h3f9e6d35, 32'h00000000} /* (30, 27, 25) {real, imag} */,
  {32'h3f0d7343, 32'h00000000} /* (30, 27, 24) {real, imag} */,
  {32'h3ea135b1, 32'h00000000} /* (30, 27, 23) {real, imag} */,
  {32'h3f0c2d6f, 32'h00000000} /* (30, 27, 22) {real, imag} */,
  {32'h3f249dad, 32'h00000000} /* (30, 27, 21) {real, imag} */,
  {32'hbea74ffb, 32'h00000000} /* (30, 27, 20) {real, imag} */,
  {32'hbf271068, 32'h00000000} /* (30, 27, 19) {real, imag} */,
  {32'hbf41b8e9, 32'h00000000} /* (30, 27, 18) {real, imag} */,
  {32'hbef6761a, 32'h00000000} /* (30, 27, 17) {real, imag} */,
  {32'hbeeb2cbb, 32'h00000000} /* (30, 27, 16) {real, imag} */,
  {32'hbf522ddc, 32'h00000000} /* (30, 27, 15) {real, imag} */,
  {32'hbf9c06ff, 32'h00000000} /* (30, 27, 14) {real, imag} */,
  {32'hbfa5bc91, 32'h00000000} /* (30, 27, 13) {real, imag} */,
  {32'hbe7f6c0f, 32'h00000000} /* (30, 27, 12) {real, imag} */,
  {32'hbedfabef, 32'h00000000} /* (30, 27, 11) {real, imag} */,
  {32'h3f2dd33a, 32'h00000000} /* (30, 27, 10) {real, imag} */,
  {32'h3faff51d, 32'h00000000} /* (30, 27, 9) {real, imag} */,
  {32'h3f9d2501, 32'h00000000} /* (30, 27, 8) {real, imag} */,
  {32'h3f8a7550, 32'h00000000} /* (30, 27, 7) {real, imag} */,
  {32'h3f605176, 32'h00000000} /* (30, 27, 6) {real, imag} */,
  {32'h3f1296d7, 32'h00000000} /* (30, 27, 5) {real, imag} */,
  {32'h3f424b9e, 32'h00000000} /* (30, 27, 4) {real, imag} */,
  {32'h3f7954b6, 32'h00000000} /* (30, 27, 3) {real, imag} */,
  {32'h3f4226b0, 32'h00000000} /* (30, 27, 2) {real, imag} */,
  {32'h3f1335c6, 32'h00000000} /* (30, 27, 1) {real, imag} */,
  {32'h3eed4900, 32'h00000000} /* (30, 27, 0) {real, imag} */,
  {32'h3f227dab, 32'h00000000} /* (30, 26, 31) {real, imag} */,
  {32'h3f83ad0d, 32'h00000000} /* (30, 26, 30) {real, imag} */,
  {32'h3f7f5c9c, 32'h00000000} /* (30, 26, 29) {real, imag} */,
  {32'h3f131feb, 32'h00000000} /* (30, 26, 28) {real, imag} */,
  {32'h3f8db17e, 32'h00000000} /* (30, 26, 27) {real, imag} */,
  {32'h3f8965d9, 32'h00000000} /* (30, 26, 26) {real, imag} */,
  {32'h3f74efee, 32'h00000000} /* (30, 26, 25) {real, imag} */,
  {32'h3f7a42e2, 32'h00000000} /* (30, 26, 24) {real, imag} */,
  {32'h3ee9585c, 32'h00000000} /* (30, 26, 23) {real, imag} */,
  {32'h3ee87cc3, 32'h00000000} /* (30, 26, 22) {real, imag} */,
  {32'h3ee534e6, 32'h00000000} /* (30, 26, 21) {real, imag} */,
  {32'hbf11b9a2, 32'h00000000} /* (30, 26, 20) {real, imag} */,
  {32'hbf3524bf, 32'h00000000} /* (30, 26, 19) {real, imag} */,
  {32'hbf069f5c, 32'h00000000} /* (30, 26, 18) {real, imag} */,
  {32'hbec2a441, 32'h00000000} /* (30, 26, 17) {real, imag} */,
  {32'hbf298287, 32'h00000000} /* (30, 26, 16) {real, imag} */,
  {32'hbfa1052c, 32'h00000000} /* (30, 26, 15) {real, imag} */,
  {32'hbf9a6c67, 32'h00000000} /* (30, 26, 14) {real, imag} */,
  {32'hbf8d3e20, 32'h00000000} /* (30, 26, 13) {real, imag} */,
  {32'hbf6d1717, 32'h00000000} /* (30, 26, 12) {real, imag} */,
  {32'hbf3ea7fb, 32'h00000000} /* (30, 26, 11) {real, imag} */,
  {32'h3e053e67, 32'h00000000} /* (30, 26, 10) {real, imag} */,
  {32'h3f52ffba, 32'h00000000} /* (30, 26, 9) {real, imag} */,
  {32'h3f7ac3d7, 32'h00000000} /* (30, 26, 8) {real, imag} */,
  {32'h3f8d1f13, 32'h00000000} /* (30, 26, 7) {real, imag} */,
  {32'h3f8a00f7, 32'h00000000} /* (30, 26, 6) {real, imag} */,
  {32'h3f49ffd7, 32'h00000000} /* (30, 26, 5) {real, imag} */,
  {32'h3f4405c6, 32'h00000000} /* (30, 26, 4) {real, imag} */,
  {32'h3fba4626, 32'h00000000} /* (30, 26, 3) {real, imag} */,
  {32'h3fa4a76c, 32'h00000000} /* (30, 26, 2) {real, imag} */,
  {32'h3f4f4d73, 32'h00000000} /* (30, 26, 1) {real, imag} */,
  {32'h3f15e3d4, 32'h00000000} /* (30, 26, 0) {real, imag} */,
  {32'h3f2bbca3, 32'h00000000} /* (30, 25, 31) {real, imag} */,
  {32'h3fb06289, 32'h00000000} /* (30, 25, 30) {real, imag} */,
  {32'h3f89f8cc, 32'h00000000} /* (30, 25, 29) {real, imag} */,
  {32'h3f2aa409, 32'h00000000} /* (30, 25, 28) {real, imag} */,
  {32'h3f9d477d, 32'h00000000} /* (30, 25, 27) {real, imag} */,
  {32'h3fa98889, 32'h00000000} /* (30, 25, 26) {real, imag} */,
  {32'h3f90ba2a, 32'h00000000} /* (30, 25, 25) {real, imag} */,
  {32'h3f49d140, 32'h00000000} /* (30, 25, 24) {real, imag} */,
  {32'h3ed4209c, 32'h00000000} /* (30, 25, 23) {real, imag} */,
  {32'h3f1cc331, 32'h00000000} /* (30, 25, 22) {real, imag} */,
  {32'h3ea6dda4, 32'h00000000} /* (30, 25, 21) {real, imag} */,
  {32'hbf8c0bcd, 32'h00000000} /* (30, 25, 20) {real, imag} */,
  {32'hbf81f25a, 32'h00000000} /* (30, 25, 19) {real, imag} */,
  {32'hbf439f72, 32'h00000000} /* (30, 25, 18) {real, imag} */,
  {32'hbf8eecef, 32'h00000000} /* (30, 25, 17) {real, imag} */,
  {32'hbf902b1a, 32'h00000000} /* (30, 25, 16) {real, imag} */,
  {32'hbfa46143, 32'h00000000} /* (30, 25, 15) {real, imag} */,
  {32'hbfeb454f, 32'h00000000} /* (30, 25, 14) {real, imag} */,
  {32'hbfb9c3eb, 32'h00000000} /* (30, 25, 13) {real, imag} */,
  {32'hbf946b1d, 32'h00000000} /* (30, 25, 12) {real, imag} */,
  {32'hbf1ded1f, 32'h00000000} /* (30, 25, 11) {real, imag} */,
  {32'h3eb698b4, 32'h00000000} /* (30, 25, 10) {real, imag} */,
  {32'h3f3da50d, 32'h00000000} /* (30, 25, 9) {real, imag} */,
  {32'h3f82a84e, 32'h00000000} /* (30, 25, 8) {real, imag} */,
  {32'h3f841986, 32'h00000000} /* (30, 25, 7) {real, imag} */,
  {32'h3f6f26be, 32'h00000000} /* (30, 25, 6) {real, imag} */,
  {32'h3fbbdb18, 32'h00000000} /* (30, 25, 5) {real, imag} */,
  {32'h3fa4fc74, 32'h00000000} /* (30, 25, 4) {real, imag} */,
  {32'h3f92563b, 32'h00000000} /* (30, 25, 3) {real, imag} */,
  {32'h3f66f496, 32'h00000000} /* (30, 25, 2) {real, imag} */,
  {32'h3eb39252, 32'h00000000} /* (30, 25, 1) {real, imag} */,
  {32'h3e9b9121, 32'h00000000} /* (30, 25, 0) {real, imag} */,
  {32'h3f62f80a, 32'h00000000} /* (30, 24, 31) {real, imag} */,
  {32'h3fcbb07e, 32'h00000000} /* (30, 24, 30) {real, imag} */,
  {32'h3fafbd19, 32'h00000000} /* (30, 24, 29) {real, imag} */,
  {32'h3f344c55, 32'h00000000} /* (30, 24, 28) {real, imag} */,
  {32'h3e96bc35, 32'h00000000} /* (30, 24, 27) {real, imag} */,
  {32'h3f806cba, 32'h00000000} /* (30, 24, 26) {real, imag} */,
  {32'h3f61a3e2, 32'h00000000} /* (30, 24, 25) {real, imag} */,
  {32'h3ee809c4, 32'h00000000} /* (30, 24, 24) {real, imag} */,
  {32'h3f1e3f8f, 32'h00000000} /* (30, 24, 23) {real, imag} */,
  {32'h3f81a15d, 32'h00000000} /* (30, 24, 22) {real, imag} */,
  {32'h3ec39133, 32'h00000000} /* (30, 24, 21) {real, imag} */,
  {32'hbf9ef985, 32'h00000000} /* (30, 24, 20) {real, imag} */,
  {32'hbf6f39b4, 32'h00000000} /* (30, 24, 19) {real, imag} */,
  {32'hbf3f603d, 32'h00000000} /* (30, 24, 18) {real, imag} */,
  {32'hbf8ae1cc, 32'h00000000} /* (30, 24, 17) {real, imag} */,
  {32'hbf92d0fd, 32'h00000000} /* (30, 24, 16) {real, imag} */,
  {32'hbf49aa13, 32'h00000000} /* (30, 24, 15) {real, imag} */,
  {32'hbfb3d3e9, 32'h00000000} /* (30, 24, 14) {real, imag} */,
  {32'hbf8fd5d2, 32'h00000000} /* (30, 24, 13) {real, imag} */,
  {32'hbf0eb6bc, 32'h00000000} /* (30, 24, 12) {real, imag} */,
  {32'hbefd3aba, 32'h00000000} /* (30, 24, 11) {real, imag} */,
  {32'h3e462a28, 32'h00000000} /* (30, 24, 10) {real, imag} */,
  {32'h3f5d2d9b, 32'h00000000} /* (30, 24, 9) {real, imag} */,
  {32'h3f9eef25, 32'h00000000} /* (30, 24, 8) {real, imag} */,
  {32'h3f95e865, 32'h00000000} /* (30, 24, 7) {real, imag} */,
  {32'h3f8592a5, 32'h00000000} /* (30, 24, 6) {real, imag} */,
  {32'h3fb2b4dd, 32'h00000000} /* (30, 24, 5) {real, imag} */,
  {32'h3f85d654, 32'h00000000} /* (30, 24, 4) {real, imag} */,
  {32'h3fbb5f3f, 32'h00000000} /* (30, 24, 3) {real, imag} */,
  {32'h3fb87c66, 32'h00000000} /* (30, 24, 2) {real, imag} */,
  {32'h3f16885c, 32'h00000000} /* (30, 24, 1) {real, imag} */,
  {32'h3ed80a9f, 32'h00000000} /* (30, 24, 0) {real, imag} */,
  {32'h3f445fa1, 32'h00000000} /* (30, 23, 31) {real, imag} */,
  {32'h3f973b35, 32'h00000000} /* (30, 23, 30) {real, imag} */,
  {32'h3f6d900d, 32'h00000000} /* (30, 23, 29) {real, imag} */,
  {32'h3f1cb2ec, 32'h00000000} /* (30, 23, 28) {real, imag} */,
  {32'h3e0e81a7, 32'h00000000} /* (30, 23, 27) {real, imag} */,
  {32'h3edfb2a7, 32'h00000000} /* (30, 23, 26) {real, imag} */,
  {32'h3efddbcc, 32'h00000000} /* (30, 23, 25) {real, imag} */,
  {32'h3ea9773a, 32'h00000000} /* (30, 23, 24) {real, imag} */,
  {32'h3f83bd9c, 32'h00000000} /* (30, 23, 23) {real, imag} */,
  {32'h3fa5b847, 32'h00000000} /* (30, 23, 22) {real, imag} */,
  {32'h3f09c244, 32'h00000000} /* (30, 23, 21) {real, imag} */,
  {32'hbf309bd7, 32'h00000000} /* (30, 23, 20) {real, imag} */,
  {32'hbf63b896, 32'h00000000} /* (30, 23, 19) {real, imag} */,
  {32'hbf68ee9e, 32'h00000000} /* (30, 23, 18) {real, imag} */,
  {32'hbf2da0a2, 32'h00000000} /* (30, 23, 17) {real, imag} */,
  {32'hbf612fb0, 32'h00000000} /* (30, 23, 16) {real, imag} */,
  {32'hbf34b1eb, 32'h00000000} /* (30, 23, 15) {real, imag} */,
  {32'hbf8a6bb1, 32'h00000000} /* (30, 23, 14) {real, imag} */,
  {32'hbf3a4c83, 32'h00000000} /* (30, 23, 13) {real, imag} */,
  {32'hbe177f18, 32'h00000000} /* (30, 23, 12) {real, imag} */,
  {32'hbef7fba1, 32'h00000000} /* (30, 23, 11) {real, imag} */,
  {32'h3b831965, 32'h00000000} /* (30, 23, 10) {real, imag} */,
  {32'h3f2bb58b, 32'h00000000} /* (30, 23, 9) {real, imag} */,
  {32'h3f80c63d, 32'h00000000} /* (30, 23, 8) {real, imag} */,
  {32'h3f84f15b, 32'h00000000} /* (30, 23, 7) {real, imag} */,
  {32'h3f42db45, 32'h00000000} /* (30, 23, 6) {real, imag} */,
  {32'h3f8111ab, 32'h00000000} /* (30, 23, 5) {real, imag} */,
  {32'h3f941e7d, 32'h00000000} /* (30, 23, 4) {real, imag} */,
  {32'h3fb0091c, 32'h00000000} /* (30, 23, 3) {real, imag} */,
  {32'h3fb513c1, 32'h00000000} /* (30, 23, 2) {real, imag} */,
  {32'h3f84297a, 32'h00000000} /* (30, 23, 1) {real, imag} */,
  {32'h3f76f85f, 32'h00000000} /* (30, 23, 0) {real, imag} */,
  {32'h3e831fc8, 32'h00000000} /* (30, 22, 31) {real, imag} */,
  {32'h3f3bf552, 32'h00000000} /* (30, 22, 30) {real, imag} */,
  {32'h3f29a568, 32'h00000000} /* (30, 22, 29) {real, imag} */,
  {32'h3e8eedd5, 32'h00000000} /* (30, 22, 28) {real, imag} */,
  {32'h3c8d53c3, 32'h00000000} /* (30, 22, 27) {real, imag} */,
  {32'h3e317ca5, 32'h00000000} /* (30, 22, 26) {real, imag} */,
  {32'h3ee58449, 32'h00000000} /* (30, 22, 25) {real, imag} */,
  {32'h3f178535, 32'h00000000} /* (30, 22, 24) {real, imag} */,
  {32'h3fb2510b, 32'h00000000} /* (30, 22, 23) {real, imag} */,
  {32'h3fc29973, 32'h00000000} /* (30, 22, 22) {real, imag} */,
  {32'h3f112c14, 32'h00000000} /* (30, 22, 21) {real, imag} */,
  {32'hbed67548, 32'h00000000} /* (30, 22, 20) {real, imag} */,
  {32'hbf34d27d, 32'h00000000} /* (30, 22, 19) {real, imag} */,
  {32'hbf361b27, 32'h00000000} /* (30, 22, 18) {real, imag} */,
  {32'hbf6e1303, 32'h00000000} /* (30, 22, 17) {real, imag} */,
  {32'hbf913a22, 32'h00000000} /* (30, 22, 16) {real, imag} */,
  {32'hbf887508, 32'h00000000} /* (30, 22, 15) {real, imag} */,
  {32'hbf5af3cf, 32'h00000000} /* (30, 22, 14) {real, imag} */,
  {32'hbf404110, 32'h00000000} /* (30, 22, 13) {real, imag} */,
  {32'hbf1f328e, 32'h00000000} /* (30, 22, 12) {real, imag} */,
  {32'hbf1d937d, 32'h00000000} /* (30, 22, 11) {real, imag} */,
  {32'h3e9dad14, 32'h00000000} /* (30, 22, 10) {real, imag} */,
  {32'h3f43f6d0, 32'h00000000} /* (30, 22, 9) {real, imag} */,
  {32'h3f1ce008, 32'h00000000} /* (30, 22, 8) {real, imag} */,
  {32'h3f7bdcaf, 32'h00000000} /* (30, 22, 7) {real, imag} */,
  {32'h3f4ccac5, 32'h00000000} /* (30, 22, 6) {real, imag} */,
  {32'h3f9950ee, 32'h00000000} /* (30, 22, 5) {real, imag} */,
  {32'h3fd78abf, 32'h00000000} /* (30, 22, 4) {real, imag} */,
  {32'h3fa6df7e, 32'h00000000} /* (30, 22, 3) {real, imag} */,
  {32'h3fb01856, 32'h00000000} /* (30, 22, 2) {real, imag} */,
  {32'h3f76dabb, 32'h00000000} /* (30, 22, 1) {real, imag} */,
  {32'h3f060382, 32'h00000000} /* (30, 22, 0) {real, imag} */,
  {32'h3d836439, 32'h00000000} /* (30, 21, 31) {real, imag} */,
  {32'h3eb89f0c, 32'h00000000} /* (30, 21, 30) {real, imag} */,
  {32'h3d70c022, 32'h00000000} /* (30, 21, 29) {real, imag} */,
  {32'hbcc6ddb4, 32'h00000000} /* (30, 21, 28) {real, imag} */,
  {32'hbd11d660, 32'h00000000} /* (30, 21, 27) {real, imag} */,
  {32'h3e40eecd, 32'h00000000} /* (30, 21, 26) {real, imag} */,
  {32'h3e6469b1, 32'h00000000} /* (30, 21, 25) {real, imag} */,
  {32'h3d50db6b, 32'h00000000} /* (30, 21, 24) {real, imag} */,
  {32'h3eb93128, 32'h00000000} /* (30, 21, 23) {real, imag} */,
  {32'hbd8b1ae9, 32'h00000000} /* (30, 21, 22) {real, imag} */,
  {32'hbe8cc3c5, 32'h00000000} /* (30, 21, 21) {real, imag} */,
  {32'hbea6455d, 32'h00000000} /* (30, 21, 20) {real, imag} */,
  {32'hbedb6bf0, 32'h00000000} /* (30, 21, 19) {real, imag} */,
  {32'hbed1cf93, 32'h00000000} /* (30, 21, 18) {real, imag} */,
  {32'hbf4f3d21, 32'h00000000} /* (30, 21, 17) {real, imag} */,
  {32'hbf5bcfdc, 32'h00000000} /* (30, 21, 16) {real, imag} */,
  {32'hbf3bfa90, 32'h00000000} /* (30, 21, 15) {real, imag} */,
  {32'hbf0dfb0d, 32'h00000000} /* (30, 21, 14) {real, imag} */,
  {32'hbeca56f3, 32'h00000000} /* (30, 21, 13) {real, imag} */,
  {32'hbeb25c32, 32'h00000000} /* (30, 21, 12) {real, imag} */,
  {32'h3d7e1e65, 32'h00000000} /* (30, 21, 11) {real, imag} */,
  {32'h3ed314d4, 32'h00000000} /* (30, 21, 10) {real, imag} */,
  {32'h3f544151, 32'h00000000} /* (30, 21, 9) {real, imag} */,
  {32'h3e0d0347, 32'h00000000} /* (30, 21, 8) {real, imag} */,
  {32'h3e8c20e8, 32'h00000000} /* (30, 21, 7) {real, imag} */,
  {32'h3eb282f5, 32'h00000000} /* (30, 21, 6) {real, imag} */,
  {32'h3ecbc252, 32'h00000000} /* (30, 21, 5) {real, imag} */,
  {32'h3f5c928f, 32'h00000000} /* (30, 21, 4) {real, imag} */,
  {32'h3f0f8e15, 32'h00000000} /* (30, 21, 3) {real, imag} */,
  {32'h3f35f608, 32'h00000000} /* (30, 21, 2) {real, imag} */,
  {32'h3ede1824, 32'h00000000} /* (30, 21, 1) {real, imag} */,
  {32'hbbbf14fa, 32'h00000000} /* (30, 21, 0) {real, imag} */,
  {32'hbdf26348, 32'h00000000} /* (30, 20, 31) {real, imag} */,
  {32'hbe672e3f, 32'h00000000} /* (30, 20, 30) {real, imag} */,
  {32'hbf3ee92c, 32'h00000000} /* (30, 20, 29) {real, imag} */,
  {32'hbf1de26f, 32'h00000000} /* (30, 20, 28) {real, imag} */,
  {32'hbf26c282, 32'h00000000} /* (30, 20, 27) {real, imag} */,
  {32'hbf21e138, 32'h00000000} /* (30, 20, 26) {real, imag} */,
  {32'hbf17f85c, 32'h00000000} /* (30, 20, 25) {real, imag} */,
  {32'hbfda1b5b, 32'h00000000} /* (30, 20, 24) {real, imag} */,
  {32'hbf86cd09, 32'h00000000} /* (30, 20, 23) {real, imag} */,
  {32'hbf6023db, 32'h00000000} /* (30, 20, 22) {real, imag} */,
  {32'hbf238eb1, 32'h00000000} /* (30, 20, 21) {real, imag} */,
  {32'h3d57f7ea, 32'h00000000} /* (30, 20, 20) {real, imag} */,
  {32'h3c941f2a, 32'h00000000} /* (30, 20, 19) {real, imag} */,
  {32'h3e55e819, 32'h00000000} /* (30, 20, 18) {real, imag} */,
  {32'h3ebf2ed2, 32'h00000000} /* (30, 20, 17) {real, imag} */,
  {32'h3e570425, 32'h00000000} /* (30, 20, 16) {real, imag} */,
  {32'h3effed17, 32'h00000000} /* (30, 20, 15) {real, imag} */,
  {32'h3f1cbf83, 32'h00000000} /* (30, 20, 14) {real, imag} */,
  {32'h3f8dfbe5, 32'h00000000} /* (30, 20, 13) {real, imag} */,
  {32'h3f502565, 32'h00000000} /* (30, 20, 12) {real, imag} */,
  {32'h3ee43666, 32'h00000000} /* (30, 20, 11) {real, imag} */,
  {32'h3d2ec2bd, 32'h00000000} /* (30, 20, 10) {real, imag} */,
  {32'hbe951740, 32'h00000000} /* (30, 20, 9) {real, imag} */,
  {32'hbf8ca58d, 32'h00000000} /* (30, 20, 8) {real, imag} */,
  {32'hbfa72f29, 32'h00000000} /* (30, 20, 7) {real, imag} */,
  {32'hbfa416e8, 32'h00000000} /* (30, 20, 6) {real, imag} */,
  {32'hbf40a115, 32'h00000000} /* (30, 20, 5) {real, imag} */,
  {32'hbf8c7d7b, 32'h00000000} /* (30, 20, 4) {real, imag} */,
  {32'hbf8df75e, 32'h00000000} /* (30, 20, 3) {real, imag} */,
  {32'hbed41052, 32'h00000000} /* (30, 20, 2) {real, imag} */,
  {32'hbeff16b5, 32'h00000000} /* (30, 20, 1) {real, imag} */,
  {32'hbee6f10a, 32'h00000000} /* (30, 20, 0) {real, imag} */,
  {32'hbecf2fbf, 32'h00000000} /* (30, 19, 31) {real, imag} */,
  {32'hbf3550e3, 32'h00000000} /* (30, 19, 30) {real, imag} */,
  {32'hbf42b402, 32'h00000000} /* (30, 19, 29) {real, imag} */,
  {32'hbf3a47c9, 32'h00000000} /* (30, 19, 28) {real, imag} */,
  {32'hbf428cac, 32'h00000000} /* (30, 19, 27) {real, imag} */,
  {32'hbf49f17b, 32'h00000000} /* (30, 19, 26) {real, imag} */,
  {32'hbf489a1e, 32'h00000000} /* (30, 19, 25) {real, imag} */,
  {32'hbf93a81e, 32'h00000000} /* (30, 19, 24) {real, imag} */,
  {32'hbf7728a6, 32'h00000000} /* (30, 19, 23) {real, imag} */,
  {32'hbf58420f, 32'h00000000} /* (30, 19, 22) {real, imag} */,
  {32'hbf17f81b, 32'h00000000} /* (30, 19, 21) {real, imag} */,
  {32'h3e862e3f, 32'h00000000} /* (30, 19, 20) {real, imag} */,
  {32'h3f0919b3, 32'h00000000} /* (30, 19, 19) {real, imag} */,
  {32'h3f5bb220, 32'h00000000} /* (30, 19, 18) {real, imag} */,
  {32'h3f3cc9a0, 32'h00000000} /* (30, 19, 17) {real, imag} */,
  {32'h3efa0f4c, 32'h00000000} /* (30, 19, 16) {real, imag} */,
  {32'h3f64659a, 32'h00000000} /* (30, 19, 15) {real, imag} */,
  {32'h3f7f37cc, 32'h00000000} /* (30, 19, 14) {real, imag} */,
  {32'h3fb510ba, 32'h00000000} /* (30, 19, 13) {real, imag} */,
  {32'h3fba8474, 32'h00000000} /* (30, 19, 12) {real, imag} */,
  {32'h3fa208f0, 32'h00000000} /* (30, 19, 11) {real, imag} */,
  {32'hbde53ca8, 32'h00000000} /* (30, 19, 10) {real, imag} */,
  {32'hbfb432cb, 32'h00000000} /* (30, 19, 9) {real, imag} */,
  {32'hbfdddfea, 32'h00000000} /* (30, 19, 8) {real, imag} */,
  {32'hbfdf97ad, 32'h00000000} /* (30, 19, 7) {real, imag} */,
  {32'hbfa36cd2, 32'h00000000} /* (30, 19, 6) {real, imag} */,
  {32'hbf1cb28d, 32'h00000000} /* (30, 19, 5) {real, imag} */,
  {32'hbf9f73d8, 32'h00000000} /* (30, 19, 4) {real, imag} */,
  {32'hbf9b8f93, 32'h00000000} /* (30, 19, 3) {real, imag} */,
  {32'hbf35be66, 32'h00000000} /* (30, 19, 2) {real, imag} */,
  {32'hbf7ec92f, 32'h00000000} /* (30, 19, 1) {real, imag} */,
  {32'hbf10ff65, 32'h00000000} /* (30, 19, 0) {real, imag} */,
  {32'hbf844a91, 32'h00000000} /* (30, 18, 31) {real, imag} */,
  {32'hbf852264, 32'h00000000} /* (30, 18, 30) {real, imag} */,
  {32'hbf0ae1b6, 32'h00000000} /* (30, 18, 29) {real, imag} */,
  {32'hbf23d5e6, 32'h00000000} /* (30, 18, 28) {real, imag} */,
  {32'hbf5d60d7, 32'h00000000} /* (30, 18, 27) {real, imag} */,
  {32'hbf117c32, 32'h00000000} /* (30, 18, 26) {real, imag} */,
  {32'hbe10be69, 32'h00000000} /* (30, 18, 25) {real, imag} */,
  {32'hbe1e345a, 32'h00000000} /* (30, 18, 24) {real, imag} */,
  {32'hbeac7de1, 32'h00000000} /* (30, 18, 23) {real, imag} */,
  {32'hbef88c0a, 32'h00000000} /* (30, 18, 22) {real, imag} */,
  {32'hbeb0af68, 32'h00000000} /* (30, 18, 21) {real, imag} */,
  {32'h3f0d22fa, 32'h00000000} /* (30, 18, 20) {real, imag} */,
  {32'h3f7b9c58, 32'h00000000} /* (30, 18, 19) {real, imag} */,
  {32'h3f83bdb5, 32'h00000000} /* (30, 18, 18) {real, imag} */,
  {32'h3f47200e, 32'h00000000} /* (30, 18, 17) {real, imag} */,
  {32'h3ec05e01, 32'h00000000} /* (30, 18, 16) {real, imag} */,
  {32'h3ef9db92, 32'h00000000} /* (30, 18, 15) {real, imag} */,
  {32'h3f54a30f, 32'h00000000} /* (30, 18, 14) {real, imag} */,
  {32'h3f8967a8, 32'h00000000} /* (30, 18, 13) {real, imag} */,
  {32'h3fc2303d, 32'h00000000} /* (30, 18, 12) {real, imag} */,
  {32'h3fbe0f15, 32'h00000000} /* (30, 18, 11) {real, imag} */,
  {32'hbf32fe4f, 32'h00000000} /* (30, 18, 10) {real, imag} */,
  {32'hbfe3a09b, 32'h00000000} /* (30, 18, 9) {real, imag} */,
  {32'hbfc1c674, 32'h00000000} /* (30, 18, 8) {real, imag} */,
  {32'hbfc11cf4, 32'h00000000} /* (30, 18, 7) {real, imag} */,
  {32'hbf518288, 32'h00000000} /* (30, 18, 6) {real, imag} */,
  {32'hbedeb083, 32'h00000000} /* (30, 18, 5) {real, imag} */,
  {32'hbf61ede1, 32'h00000000} /* (30, 18, 4) {real, imag} */,
  {32'hbf6fcfbd, 32'h00000000} /* (30, 18, 3) {real, imag} */,
  {32'hbf30afe7, 32'h00000000} /* (30, 18, 2) {real, imag} */,
  {32'hbf490799, 32'h00000000} /* (30, 18, 1) {real, imag} */,
  {32'hbf0a230b, 32'h00000000} /* (30, 18, 0) {real, imag} */,
  {32'hbf7af7ac, 32'h00000000} /* (30, 17, 31) {real, imag} */,
  {32'hbfad0dfd, 32'h00000000} /* (30, 17, 30) {real, imag} */,
  {32'hbf603084, 32'h00000000} /* (30, 17, 29) {real, imag} */,
  {32'hbf631ab2, 32'h00000000} /* (30, 17, 28) {real, imag} */,
  {32'hbf7649d4, 32'h00000000} /* (30, 17, 27) {real, imag} */,
  {32'hbec0e7ce, 32'h00000000} /* (30, 17, 26) {real, imag} */,
  {32'hbe4acc33, 32'h00000000} /* (30, 17, 25) {real, imag} */,
  {32'hbee1707d, 32'h00000000} /* (30, 17, 24) {real, imag} */,
  {32'hbe8c47c2, 32'h00000000} /* (30, 17, 23) {real, imag} */,
  {32'hbf0fc809, 32'h00000000} /* (30, 17, 22) {real, imag} */,
  {32'hbee1363d, 32'h00000000} /* (30, 17, 21) {real, imag} */,
  {32'h3f71b77b, 32'h00000000} /* (30, 17, 20) {real, imag} */,
  {32'h3f67785d, 32'h00000000} /* (30, 17, 19) {real, imag} */,
  {32'h3f47f509, 32'h00000000} /* (30, 17, 18) {real, imag} */,
  {32'h3f8b27fa, 32'h00000000} /* (30, 17, 17) {real, imag} */,
  {32'h3f111ab0, 32'h00000000} /* (30, 17, 16) {real, imag} */,
  {32'h3f16abb0, 32'h00000000} /* (30, 17, 15) {real, imag} */,
  {32'h3f7b44c0, 32'h00000000} /* (30, 17, 14) {real, imag} */,
  {32'h3f574d0d, 32'h00000000} /* (30, 17, 13) {real, imag} */,
  {32'h3f957b34, 32'h00000000} /* (30, 17, 12) {real, imag} */,
  {32'h3fa3d8d0, 32'h00000000} /* (30, 17, 11) {real, imag} */,
  {32'hbf208035, 32'h00000000} /* (30, 17, 10) {real, imag} */,
  {32'hbf92090a, 32'h00000000} /* (30, 17, 9) {real, imag} */,
  {32'hbf78bdde, 32'h00000000} /* (30, 17, 8) {real, imag} */,
  {32'hbf428ffe, 32'h00000000} /* (30, 17, 7) {real, imag} */,
  {32'hbf525ddc, 32'h00000000} /* (30, 17, 6) {real, imag} */,
  {32'hbf351998, 32'h00000000} /* (30, 17, 5) {real, imag} */,
  {32'hbf6d919a, 32'h00000000} /* (30, 17, 4) {real, imag} */,
  {32'hbf67505d, 32'h00000000} /* (30, 17, 3) {real, imag} */,
  {32'hbf3d1fd7, 32'h00000000} /* (30, 17, 2) {real, imag} */,
  {32'hbf45e3d4, 32'h00000000} /* (30, 17, 1) {real, imag} */,
  {32'hbefc70c6, 32'h00000000} /* (30, 17, 0) {real, imag} */,
  {32'hbf0d30b1, 32'h00000000} /* (30, 16, 31) {real, imag} */,
  {32'hbf9a9d35, 32'h00000000} /* (30, 16, 30) {real, imag} */,
  {32'hbf9aa629, 32'h00000000} /* (30, 16, 29) {real, imag} */,
  {32'hbf164de9, 32'h00000000} /* (30, 16, 28) {real, imag} */,
  {32'hbf1af9e4, 32'h00000000} /* (30, 16, 27) {real, imag} */,
  {32'hbed1ce1e, 32'h00000000} /* (30, 16, 26) {real, imag} */,
  {32'hbf37c7c0, 32'h00000000} /* (30, 16, 25) {real, imag} */,
  {32'hbfcb0866, 32'h00000000} /* (30, 16, 24) {real, imag} */,
  {32'hbf437c68, 32'h00000000} /* (30, 16, 23) {real, imag} */,
  {32'hbef5b016, 32'h00000000} /* (30, 16, 22) {real, imag} */,
  {32'h3d5dbb6e, 32'h00000000} /* (30, 16, 21) {real, imag} */,
  {32'h3f974599, 32'h00000000} /* (30, 16, 20) {real, imag} */,
  {32'h3fb8e06e, 32'h00000000} /* (30, 16, 19) {real, imag} */,
  {32'h3f67916b, 32'h00000000} /* (30, 16, 18) {real, imag} */,
  {32'h3f5a0e37, 32'h00000000} /* (30, 16, 17) {real, imag} */,
  {32'h3f545c12, 32'h00000000} /* (30, 16, 16) {real, imag} */,
  {32'h3f77ae00, 32'h00000000} /* (30, 16, 15) {real, imag} */,
  {32'h3f53e64d, 32'h00000000} /* (30, 16, 14) {real, imag} */,
  {32'h3f552434, 32'h00000000} /* (30, 16, 13) {real, imag} */,
  {32'h3f8514dc, 32'h00000000} /* (30, 16, 12) {real, imag} */,
  {32'h3ea757cc, 32'h00000000} /* (30, 16, 11) {real, imag} */,
  {32'hbf8ef420, 32'h00000000} /* (30, 16, 10) {real, imag} */,
  {32'hbf7b4e8f, 32'h00000000} /* (30, 16, 9) {real, imag} */,
  {32'hbf09ef12, 32'h00000000} /* (30, 16, 8) {real, imag} */,
  {32'hbf1b34e0, 32'h00000000} /* (30, 16, 7) {real, imag} */,
  {32'hbf963704, 32'h00000000} /* (30, 16, 6) {real, imag} */,
  {32'hbf9bc476, 32'h00000000} /* (30, 16, 5) {real, imag} */,
  {32'hbf8dc960, 32'h00000000} /* (30, 16, 4) {real, imag} */,
  {32'hbf8aa7d8, 32'h00000000} /* (30, 16, 3) {real, imag} */,
  {32'hbf8411e5, 32'h00000000} /* (30, 16, 2) {real, imag} */,
  {32'hbf80ef73, 32'h00000000} /* (30, 16, 1) {real, imag} */,
  {32'hbec14395, 32'h00000000} /* (30, 16, 0) {real, imag} */,
  {32'hbee17996, 32'h00000000} /* (30, 15, 31) {real, imag} */,
  {32'hbf89c6ad, 32'h00000000} /* (30, 15, 30) {real, imag} */,
  {32'hbf9c75c9, 32'h00000000} /* (30, 15, 29) {real, imag} */,
  {32'hbf5caae0, 32'h00000000} /* (30, 15, 28) {real, imag} */,
  {32'hbf020667, 32'h00000000} /* (30, 15, 27) {real, imag} */,
  {32'hbe82e210, 32'h00000000} /* (30, 15, 26) {real, imag} */,
  {32'hbf2c6ce0, 32'h00000000} /* (30, 15, 25) {real, imag} */,
  {32'hbf35ddab, 32'h00000000} /* (30, 15, 24) {real, imag} */,
  {32'hbea4c7bc, 32'h00000000} /* (30, 15, 23) {real, imag} */,
  {32'hbed2935a, 32'h00000000} /* (30, 15, 22) {real, imag} */,
  {32'hbcbfef6f, 32'h00000000} /* (30, 15, 21) {real, imag} */,
  {32'h3f0783ac, 32'h00000000} /* (30, 15, 20) {real, imag} */,
  {32'h3f828c1b, 32'h00000000} /* (30, 15, 19) {real, imag} */,
  {32'h3f7000cf, 32'h00000000} /* (30, 15, 18) {real, imag} */,
  {32'h3f00913a, 32'h00000000} /* (30, 15, 17) {real, imag} */,
  {32'h3f656150, 32'h00000000} /* (30, 15, 16) {real, imag} */,
  {32'h3f996f9b, 32'h00000000} /* (30, 15, 15) {real, imag} */,
  {32'h3f886c78, 32'h00000000} /* (30, 15, 14) {real, imag} */,
  {32'h3f52a6bf, 32'h00000000} /* (30, 15, 13) {real, imag} */,
  {32'h3f1d4331, 32'h00000000} /* (30, 15, 12) {real, imag} */,
  {32'h3da5f6cb, 32'h00000000} /* (30, 15, 11) {real, imag} */,
  {32'hbf7ce0ab, 32'h00000000} /* (30, 15, 10) {real, imag} */,
  {32'hbf96f4cf, 32'h00000000} /* (30, 15, 9) {real, imag} */,
  {32'hbf869a6d, 32'h00000000} /* (30, 15, 8) {real, imag} */,
  {32'hbf878f72, 32'h00000000} /* (30, 15, 7) {real, imag} */,
  {32'hbf812156, 32'h00000000} /* (30, 15, 6) {real, imag} */,
  {32'hbfc07db1, 32'h00000000} /* (30, 15, 5) {real, imag} */,
  {32'hbf87ef8d, 32'h00000000} /* (30, 15, 4) {real, imag} */,
  {32'hbf691a66, 32'h00000000} /* (30, 15, 3) {real, imag} */,
  {32'hbf45ddc5, 32'h00000000} /* (30, 15, 2) {real, imag} */,
  {32'hbf3728ef, 32'h00000000} /* (30, 15, 1) {real, imag} */,
  {32'hbe4f1d70, 32'h00000000} /* (30, 15, 0) {real, imag} */,
  {32'hbf16b58d, 32'h00000000} /* (30, 14, 31) {real, imag} */,
  {32'hbfa4a884, 32'h00000000} /* (30, 14, 30) {real, imag} */,
  {32'hbf92da8b, 32'h00000000} /* (30, 14, 29) {real, imag} */,
  {32'hbf4fc397, 32'h00000000} /* (30, 14, 28) {real, imag} */,
  {32'hbef44389, 32'h00000000} /* (30, 14, 27) {real, imag} */,
  {32'hbea4de6d, 32'h00000000} /* (30, 14, 26) {real, imag} */,
  {32'hbf4961e7, 32'h00000000} /* (30, 14, 25) {real, imag} */,
  {32'hbf5edaef, 32'h00000000} /* (30, 14, 24) {real, imag} */,
  {32'hbf1a6c21, 32'h00000000} /* (30, 14, 23) {real, imag} */,
  {32'hbf3d1c1b, 32'h00000000} /* (30, 14, 22) {real, imag} */,
  {32'hbe6dd925, 32'h00000000} /* (30, 14, 21) {real, imag} */,
  {32'h3f47507f, 32'h00000000} /* (30, 14, 20) {real, imag} */,
  {32'h3f0d0bcb, 32'h00000000} /* (30, 14, 19) {real, imag} */,
  {32'h3f1855b7, 32'h00000000} /* (30, 14, 18) {real, imag} */,
  {32'h3edc85e8, 32'h00000000} /* (30, 14, 17) {real, imag} */,
  {32'h3f819eb7, 32'h00000000} /* (30, 14, 16) {real, imag} */,
  {32'h3f99f2c3, 32'h00000000} /* (30, 14, 15) {real, imag} */,
  {32'h3f5c4038, 32'h00000000} /* (30, 14, 14) {real, imag} */,
  {32'h3efad3c2, 32'h00000000} /* (30, 14, 13) {real, imag} */,
  {32'h3edff944, 32'h00000000} /* (30, 14, 12) {real, imag} */,
  {32'h3f0f2fdd, 32'h00000000} /* (30, 14, 11) {real, imag} */,
  {32'hbec76dd0, 32'h00000000} /* (30, 14, 10) {real, imag} */,
  {32'hbf9ba0fd, 32'h00000000} /* (30, 14, 9) {real, imag} */,
  {32'hbfa19829, 32'h00000000} /* (30, 14, 8) {real, imag} */,
  {32'hbf5ef9de, 32'h00000000} /* (30, 14, 7) {real, imag} */,
  {32'hbf3fae35, 32'h00000000} /* (30, 14, 6) {real, imag} */,
  {32'hbfbd7940, 32'h00000000} /* (30, 14, 5) {real, imag} */,
  {32'hbf6b833b, 32'h00000000} /* (30, 14, 4) {real, imag} */,
  {32'hbf610530, 32'h00000000} /* (30, 14, 3) {real, imag} */,
  {32'hbede49bc, 32'h00000000} /* (30, 14, 2) {real, imag} */,
  {32'hbcd93b0c, 32'h00000000} /* (30, 14, 1) {real, imag} */,
  {32'hbe2bc164, 32'h00000000} /* (30, 14, 0) {real, imag} */,
  {32'hbf2a857c, 32'h00000000} /* (30, 13, 31) {real, imag} */,
  {32'hbf7b21fb, 32'h00000000} /* (30, 13, 30) {real, imag} */,
  {32'hbf44243e, 32'h00000000} /* (30, 13, 29) {real, imag} */,
  {32'hbf545360, 32'h00000000} /* (30, 13, 28) {real, imag} */,
  {32'hbf762a63, 32'h00000000} /* (30, 13, 27) {real, imag} */,
  {32'hbf32237a, 32'h00000000} /* (30, 13, 26) {real, imag} */,
  {32'hbf7ec23a, 32'h00000000} /* (30, 13, 25) {real, imag} */,
  {32'hbfd19264, 32'h00000000} /* (30, 13, 24) {real, imag} */,
  {32'hbfa4e93f, 32'h00000000} /* (30, 13, 23) {real, imag} */,
  {32'hbf81dde4, 32'h00000000} /* (30, 13, 22) {real, imag} */,
  {32'hbf1e1298, 32'h00000000} /* (30, 13, 21) {real, imag} */,
  {32'h3f282c26, 32'h00000000} /* (30, 13, 20) {real, imag} */,
  {32'h3f5300a4, 32'h00000000} /* (30, 13, 19) {real, imag} */,
  {32'h3f019833, 32'h00000000} /* (30, 13, 18) {real, imag} */,
  {32'h3f36918b, 32'h00000000} /* (30, 13, 17) {real, imag} */,
  {32'h3f830c79, 32'h00000000} /* (30, 13, 16) {real, imag} */,
  {32'h3f90f02b, 32'h00000000} /* (30, 13, 15) {real, imag} */,
  {32'h3f2c4cbf, 32'h00000000} /* (30, 13, 14) {real, imag} */,
  {32'h3ebe6384, 32'h00000000} /* (30, 13, 13) {real, imag} */,
  {32'h3f0c44a3, 32'h00000000} /* (30, 13, 12) {real, imag} */,
  {32'h3f172e61, 32'h00000000} /* (30, 13, 11) {real, imag} */,
  {32'hbe648dfa, 32'h00000000} /* (30, 13, 10) {real, imag} */,
  {32'hbf7745ac, 32'h00000000} /* (30, 13, 9) {real, imag} */,
  {32'hbfbbaa66, 32'h00000000} /* (30, 13, 8) {real, imag} */,
  {32'hbf929f1a, 32'h00000000} /* (30, 13, 7) {real, imag} */,
  {32'hbf9aac5e, 32'h00000000} /* (30, 13, 6) {real, imag} */,
  {32'hbfdd54df, 32'h00000000} /* (30, 13, 5) {real, imag} */,
  {32'hbfc06b60, 32'h00000000} /* (30, 13, 4) {real, imag} */,
  {32'hbfa4a050, 32'h00000000} /* (30, 13, 3) {real, imag} */,
  {32'hbeb6ed1e, 32'h00000000} /* (30, 13, 2) {real, imag} */,
  {32'hbeab1eff, 32'h00000000} /* (30, 13, 1) {real, imag} */,
  {32'hbef278f7, 32'h00000000} /* (30, 13, 0) {real, imag} */,
  {32'hbf0721e2, 32'h00000000} /* (30, 12, 31) {real, imag} */,
  {32'hbf077cf0, 32'h00000000} /* (30, 12, 30) {real, imag} */,
  {32'hbede2b82, 32'h00000000} /* (30, 12, 29) {real, imag} */,
  {32'hbf34eaba, 32'h00000000} /* (30, 12, 28) {real, imag} */,
  {32'hbfa82326, 32'h00000000} /* (30, 12, 27) {real, imag} */,
  {32'hbf726f38, 32'h00000000} /* (30, 12, 26) {real, imag} */,
  {32'hbf81bacc, 32'h00000000} /* (30, 12, 25) {real, imag} */,
  {32'hbf8599d4, 32'h00000000} /* (30, 12, 24) {real, imag} */,
  {32'hbf73bd33, 32'h00000000} /* (30, 12, 23) {real, imag} */,
  {32'hbfa80daa, 32'h00000000} /* (30, 12, 22) {real, imag} */,
  {32'hbf55c2d9, 32'h00000000} /* (30, 12, 21) {real, imag} */,
  {32'h3eb50ab8, 32'h00000000} /* (30, 12, 20) {real, imag} */,
  {32'h3f98baf6, 32'h00000000} /* (30, 12, 19) {real, imag} */,
  {32'h3f648b73, 32'h00000000} /* (30, 12, 18) {real, imag} */,
  {32'h3f778700, 32'h00000000} /* (30, 12, 17) {real, imag} */,
  {32'h3f92fe77, 32'h00000000} /* (30, 12, 16) {real, imag} */,
  {32'h3f5426d2, 32'h00000000} /* (30, 12, 15) {real, imag} */,
  {32'h3f4634a3, 32'h00000000} /* (30, 12, 14) {real, imag} */,
  {32'h3f3e1265, 32'h00000000} /* (30, 12, 13) {real, imag} */,
  {32'h3f3cf1a5, 32'h00000000} /* (30, 12, 12) {real, imag} */,
  {32'h3f16446d, 32'h00000000} /* (30, 12, 11) {real, imag} */,
  {32'hbe418f74, 32'h00000000} /* (30, 12, 10) {real, imag} */,
  {32'hbf4f2ee2, 32'h00000000} /* (30, 12, 9) {real, imag} */,
  {32'hbf8a6e08, 32'h00000000} /* (30, 12, 8) {real, imag} */,
  {32'hbf70bb9a, 32'h00000000} /* (30, 12, 7) {real, imag} */,
  {32'hbf904d6e, 32'h00000000} /* (30, 12, 6) {real, imag} */,
  {32'hbfa027e6, 32'h00000000} /* (30, 12, 5) {real, imag} */,
  {32'hbfa66662, 32'h00000000} /* (30, 12, 4) {real, imag} */,
  {32'hbfb0582c, 32'h00000000} /* (30, 12, 3) {real, imag} */,
  {32'hbf546ce0, 32'h00000000} /* (30, 12, 2) {real, imag} */,
  {32'hbf5f3adf, 32'h00000000} /* (30, 12, 1) {real, imag} */,
  {32'hbf4d9294, 32'h00000000} /* (30, 12, 0) {real, imag} */,
  {32'hbe4036ba, 32'h00000000} /* (30, 11, 31) {real, imag} */,
  {32'hbea27d88, 32'h00000000} /* (30, 11, 30) {real, imag} */,
  {32'hbf30d2a7, 32'h00000000} /* (30, 11, 29) {real, imag} */,
  {32'hbf514c58, 32'h00000000} /* (30, 11, 28) {real, imag} */,
  {32'hbf2cfdb6, 32'h00000000} /* (30, 11, 27) {real, imag} */,
  {32'hbedaceff, 32'h00000000} /* (30, 11, 26) {real, imag} */,
  {32'hbf7d3332, 32'h00000000} /* (30, 11, 25) {real, imag} */,
  {32'hbf091224, 32'h00000000} /* (30, 11, 24) {real, imag} */,
  {32'hbec86c38, 32'h00000000} /* (30, 11, 23) {real, imag} */,
  {32'hbf8a54ef, 32'h00000000} /* (30, 11, 22) {real, imag} */,
  {32'hbf11aee9, 32'h00000000} /* (30, 11, 21) {real, imag} */,
  {32'h3ed54825, 32'h00000000} /* (30, 11, 20) {real, imag} */,
  {32'h3f6e9a9d, 32'h00000000} /* (30, 11, 19) {real, imag} */,
  {32'h3f412bfa, 32'h00000000} /* (30, 11, 18) {real, imag} */,
  {32'h3fa3dd15, 32'h00000000} /* (30, 11, 17) {real, imag} */,
  {32'h3fb829da, 32'h00000000} /* (30, 11, 16) {real, imag} */,
  {32'h3f4e7d6d, 32'h00000000} /* (30, 11, 15) {real, imag} */,
  {32'h3f8406e2, 32'h00000000} /* (30, 11, 14) {real, imag} */,
  {32'h3f280e4a, 32'h00000000} /* (30, 11, 13) {real, imag} */,
  {32'h3e9e6318, 32'h00000000} /* (30, 11, 12) {real, imag} */,
  {32'h3f0c0865, 32'h00000000} /* (30, 11, 11) {real, imag} */,
  {32'hbe35880d, 32'h00000000} /* (30, 11, 10) {real, imag} */,
  {32'hbf89cc0e, 32'h00000000} /* (30, 11, 9) {real, imag} */,
  {32'hbf11fa2b, 32'h00000000} /* (30, 11, 8) {real, imag} */,
  {32'hbe250aba, 32'h00000000} /* (30, 11, 7) {real, imag} */,
  {32'hbec878ee, 32'h00000000} /* (30, 11, 6) {real, imag} */,
  {32'hbf181e1f, 32'h00000000} /* (30, 11, 5) {real, imag} */,
  {32'hbecdc9c2, 32'h00000000} /* (30, 11, 4) {real, imag} */,
  {32'hbf974d89, 32'h00000000} /* (30, 11, 3) {real, imag} */,
  {32'hbf229ce1, 32'h00000000} /* (30, 11, 2) {real, imag} */,
  {32'hbee8244c, 32'h00000000} /* (30, 11, 1) {real, imag} */,
  {32'hbeed9354, 32'h00000000} /* (30, 11, 0) {real, imag} */,
  {32'h3f21d28a, 32'h00000000} /* (30, 10, 31) {real, imag} */,
  {32'h3f243fae, 32'h00000000} /* (30, 10, 30) {real, imag} */,
  {32'h3ac494aa, 32'h00000000} /* (30, 10, 29) {real, imag} */,
  {32'h3d509d78, 32'h00000000} /* (30, 10, 28) {real, imag} */,
  {32'h3f113d66, 32'h00000000} /* (30, 10, 27) {real, imag} */,
  {32'h3f0945e9, 32'h00000000} /* (30, 10, 26) {real, imag} */,
  {32'h3f0650bf, 32'h00000000} /* (30, 10, 25) {real, imag} */,
  {32'h3ea68543, 32'h00000000} /* (30, 10, 24) {real, imag} */,
  {32'h3efdba54, 32'h00000000} /* (30, 10, 23) {real, imag} */,
  {32'h3e3c68c5, 32'h00000000} /* (30, 10, 22) {real, imag} */,
  {32'hbe3f4363, 32'h00000000} /* (30, 10, 21) {real, imag} */,
  {32'hbe38a50a, 32'h00000000} /* (30, 10, 20) {real, imag} */,
  {32'hbd8133b9, 32'h00000000} /* (30, 10, 19) {real, imag} */,
  {32'hbc911e01, 32'h00000000} /* (30, 10, 18) {real, imag} */,
  {32'h3d15aa48, 32'h00000000} /* (30, 10, 17) {real, imag} */,
  {32'hbd8c73ce, 32'h00000000} /* (30, 10, 16) {real, imag} */,
  {32'hbf033519, 32'h00000000} /* (30, 10, 15) {real, imag} */,
  {32'hbeba16ad, 32'h00000000} /* (30, 10, 14) {real, imag} */,
  {32'hbf14b476, 32'h00000000} /* (30, 10, 13) {real, imag} */,
  {32'hbefae4e0, 32'h00000000} /* (30, 10, 12) {real, imag} */,
  {32'h3e8a3f8b, 32'h00000000} /* (30, 10, 11) {real, imag} */,
  {32'h3e961ef7, 32'h00000000} /* (30, 10, 10) {real, imag} */,
  {32'h3e09f28a, 32'h00000000} /* (30, 10, 9) {real, imag} */,
  {32'h3f1ee731, 32'h00000000} /* (30, 10, 8) {real, imag} */,
  {32'h3f8f5691, 32'h00000000} /* (30, 10, 7) {real, imag} */,
  {32'h3f7e7327, 32'h00000000} /* (30, 10, 6) {real, imag} */,
  {32'h3f2ccddf, 32'h00000000} /* (30, 10, 5) {real, imag} */,
  {32'h3f6e35e0, 32'h00000000} /* (30, 10, 4) {real, imag} */,
  {32'h3ead82ef, 32'h00000000} /* (30, 10, 3) {real, imag} */,
  {32'h3ef96777, 32'h00000000} /* (30, 10, 2) {real, imag} */,
  {32'h3f05e981, 32'h00000000} /* (30, 10, 1) {real, imag} */,
  {32'h3ebfcf2e, 32'h00000000} /* (30, 10, 0) {real, imag} */,
  {32'h3f1e1ba6, 32'h00000000} /* (30, 9, 31) {real, imag} */,
  {32'h3f931a47, 32'h00000000} /* (30, 9, 30) {real, imag} */,
  {32'h3f5aab68, 32'h00000000} /* (30, 9, 29) {real, imag} */,
  {32'h3f533ce4, 32'h00000000} /* (30, 9, 28) {real, imag} */,
  {32'h3f793779, 32'h00000000} /* (30, 9, 27) {real, imag} */,
  {32'h3f7f66b4, 32'h00000000} /* (30, 9, 26) {real, imag} */,
  {32'h3f83f272, 32'h00000000} /* (30, 9, 25) {real, imag} */,
  {32'h3f45beec, 32'h00000000} /* (30, 9, 24) {real, imag} */,
  {32'h3f192cea, 32'h00000000} /* (30, 9, 23) {real, imag} */,
  {32'h3f2e2533, 32'h00000000} /* (30, 9, 22) {real, imag} */,
  {32'h3eae322c, 32'h00000000} /* (30, 9, 21) {real, imag} */,
  {32'hbec0675f, 32'h00000000} /* (30, 9, 20) {real, imag} */,
  {32'hbf00bf89, 32'h00000000} /* (30, 9, 19) {real, imag} */,
  {32'hbeeb9733, 32'h00000000} /* (30, 9, 18) {real, imag} */,
  {32'hbf630acd, 32'h00000000} /* (30, 9, 17) {real, imag} */,
  {32'hbfa7f852, 32'h00000000} /* (30, 9, 16) {real, imag} */,
  {32'hbf8ece9c, 32'h00000000} /* (30, 9, 15) {real, imag} */,
  {32'hbf88a882, 32'h00000000} /* (30, 9, 14) {real, imag} */,
  {32'hbf390e56, 32'h00000000} /* (30, 9, 13) {real, imag} */,
  {32'hbf7ac9c3, 32'h00000000} /* (30, 9, 12) {real, imag} */,
  {32'hbf0b0dc0, 32'h00000000} /* (30, 9, 11) {real, imag} */,
  {32'h3e318b38, 32'h00000000} /* (30, 9, 10) {real, imag} */,
  {32'h3f1a1dc0, 32'h00000000} /* (30, 9, 9) {real, imag} */,
  {32'h3f228725, 32'h00000000} /* (30, 9, 8) {real, imag} */,
  {32'h3f855fce, 32'h00000000} /* (30, 9, 7) {real, imag} */,
  {32'h3f48544d, 32'h00000000} /* (30, 9, 6) {real, imag} */,
  {32'h3f97b282, 32'h00000000} /* (30, 9, 5) {real, imag} */,
  {32'h3f902c00, 32'h00000000} /* (30, 9, 4) {real, imag} */,
  {32'h3f95d252, 32'h00000000} /* (30, 9, 3) {real, imag} */,
  {32'h3f805f4d, 32'h00000000} /* (30, 9, 2) {real, imag} */,
  {32'h3f8e8d8b, 32'h00000000} /* (30, 9, 1) {real, imag} */,
  {32'h3f2aedee, 32'h00000000} /* (30, 9, 0) {real, imag} */,
  {32'h3f01c23d, 32'h00000000} /* (30, 8, 31) {real, imag} */,
  {32'h3f75638b, 32'h00000000} /* (30, 8, 30) {real, imag} */,
  {32'h3f71e597, 32'h00000000} /* (30, 8, 29) {real, imag} */,
  {32'h3f37db44, 32'h00000000} /* (30, 8, 28) {real, imag} */,
  {32'h3f7821e9, 32'h00000000} /* (30, 8, 27) {real, imag} */,
  {32'h3f9da32c, 32'h00000000} /* (30, 8, 26) {real, imag} */,
  {32'h3f727a01, 32'h00000000} /* (30, 8, 25) {real, imag} */,
  {32'h3f3c0baf, 32'h00000000} /* (30, 8, 24) {real, imag} */,
  {32'h3f1e315f, 32'h00000000} /* (30, 8, 23) {real, imag} */,
  {32'h3f2b106f, 32'h00000000} /* (30, 8, 22) {real, imag} */,
  {32'h3e9b6d23, 32'h00000000} /* (30, 8, 21) {real, imag} */,
  {32'hbf50df75, 32'h00000000} /* (30, 8, 20) {real, imag} */,
  {32'hbf4adb23, 32'h00000000} /* (30, 8, 19) {real, imag} */,
  {32'hbf43023f, 32'h00000000} /* (30, 8, 18) {real, imag} */,
  {32'hbf729d79, 32'h00000000} /* (30, 8, 17) {real, imag} */,
  {32'hbf7deb4c, 32'h00000000} /* (30, 8, 16) {real, imag} */,
  {32'hbf7adf50, 32'h00000000} /* (30, 8, 15) {real, imag} */,
  {32'hbfe1c71a, 32'h00000000} /* (30, 8, 14) {real, imag} */,
  {32'hbfa38d5a, 32'h00000000} /* (30, 8, 13) {real, imag} */,
  {32'hbff0b6e4, 32'h00000000} /* (30, 8, 12) {real, imag} */,
  {32'hbf98b6c9, 32'h00000000} /* (30, 8, 11) {real, imag} */,
  {32'hbc9b0921, 32'h00000000} /* (30, 8, 10) {real, imag} */,
  {32'h3f0669ac, 32'h00000000} /* (30, 8, 9) {real, imag} */,
  {32'h3e82e396, 32'h00000000} /* (30, 8, 8) {real, imag} */,
  {32'h3f215054, 32'h00000000} /* (30, 8, 7) {real, imag} */,
  {32'h3f39b760, 32'h00000000} /* (30, 8, 6) {real, imag} */,
  {32'h3f2f6196, 32'h00000000} /* (30, 8, 5) {real, imag} */,
  {32'h3f658225, 32'h00000000} /* (30, 8, 4) {real, imag} */,
  {32'h3fb01f63, 32'h00000000} /* (30, 8, 3) {real, imag} */,
  {32'h3f8c9a9e, 32'h00000000} /* (30, 8, 2) {real, imag} */,
  {32'h3f859f28, 32'h00000000} /* (30, 8, 1) {real, imag} */,
  {32'h3f182a16, 32'h00000000} /* (30, 8, 0) {real, imag} */,
  {32'h3f31b075, 32'h00000000} /* (30, 7, 31) {real, imag} */,
  {32'h3f1e80a5, 32'h00000000} /* (30, 7, 30) {real, imag} */,
  {32'h3f2b92bf, 32'h00000000} /* (30, 7, 29) {real, imag} */,
  {32'h3f5714f2, 32'h00000000} /* (30, 7, 28) {real, imag} */,
  {32'h3f2b7855, 32'h00000000} /* (30, 7, 27) {real, imag} */,
  {32'h3f35f4a5, 32'h00000000} /* (30, 7, 26) {real, imag} */,
  {32'h3f6eed43, 32'h00000000} /* (30, 7, 25) {real, imag} */,
  {32'h3f54fcf2, 32'h00000000} /* (30, 7, 24) {real, imag} */,
  {32'h3f4ea3b1, 32'h00000000} /* (30, 7, 23) {real, imag} */,
  {32'h3f2f5acb, 32'h00000000} /* (30, 7, 22) {real, imag} */,
  {32'hbd95cae9, 32'h00000000} /* (30, 7, 21) {real, imag} */,
  {32'hbf7cc766, 32'h00000000} /* (30, 7, 20) {real, imag} */,
  {32'hbf3ef646, 32'h00000000} /* (30, 7, 19) {real, imag} */,
  {32'hbf272d23, 32'h00000000} /* (30, 7, 18) {real, imag} */,
  {32'hbf37d94f, 32'h00000000} /* (30, 7, 17) {real, imag} */,
  {32'hbf315548, 32'h00000000} /* (30, 7, 16) {real, imag} */,
  {32'hbf0e99db, 32'h00000000} /* (30, 7, 15) {real, imag} */,
  {32'hbf898a57, 32'h00000000} /* (30, 7, 14) {real, imag} */,
  {32'hbf44cdc3, 32'h00000000} /* (30, 7, 13) {real, imag} */,
  {32'hbf993747, 32'h00000000} /* (30, 7, 12) {real, imag} */,
  {32'hbf97065f, 32'h00000000} /* (30, 7, 11) {real, imag} */,
  {32'h3ebbfa5a, 32'h00000000} /* (30, 7, 10) {real, imag} */,
  {32'h3f6cf977, 32'h00000000} /* (30, 7, 9) {real, imag} */,
  {32'h3f41a2f7, 32'h00000000} /* (30, 7, 8) {real, imag} */,
  {32'h3f86cbb3, 32'h00000000} /* (30, 7, 7) {real, imag} */,
  {32'h3f89ad9c, 32'h00000000} /* (30, 7, 6) {real, imag} */,
  {32'h3f99d07b, 32'h00000000} /* (30, 7, 5) {real, imag} */,
  {32'h3f85e14c, 32'h00000000} /* (30, 7, 4) {real, imag} */,
  {32'h3fb87e3f, 32'h00000000} /* (30, 7, 3) {real, imag} */,
  {32'h3fc8cbd1, 32'h00000000} /* (30, 7, 2) {real, imag} */,
  {32'h3f80485e, 32'h00000000} /* (30, 7, 1) {real, imag} */,
  {32'h3f0437f3, 32'h00000000} /* (30, 7, 0) {real, imag} */,
  {32'h3f16fc69, 32'h00000000} /* (30, 6, 31) {real, imag} */,
  {32'h3f3c35c9, 32'h00000000} /* (30, 6, 30) {real, imag} */,
  {32'h3f83ec33, 32'h00000000} /* (30, 6, 29) {real, imag} */,
  {32'h3f2fb6e1, 32'h00000000} /* (30, 6, 28) {real, imag} */,
  {32'h3e4414ba, 32'h00000000} /* (30, 6, 27) {real, imag} */,
  {32'h3e5fe125, 32'h00000000} /* (30, 6, 26) {real, imag} */,
  {32'h3f5ff59f, 32'h00000000} /* (30, 6, 25) {real, imag} */,
  {32'h3f9da45c, 32'h00000000} /* (30, 6, 24) {real, imag} */,
  {32'h3f77ab0c, 32'h00000000} /* (30, 6, 23) {real, imag} */,
  {32'h3f3ef3e4, 32'h00000000} /* (30, 6, 22) {real, imag} */,
  {32'h3eb85828, 32'h00000000} /* (30, 6, 21) {real, imag} */,
  {32'hbf150e6b, 32'h00000000} /* (30, 6, 20) {real, imag} */,
  {32'hbeee95b5, 32'h00000000} /* (30, 6, 19) {real, imag} */,
  {32'hbf119b75, 32'h00000000} /* (30, 6, 18) {real, imag} */,
  {32'hbf87c4a6, 32'h00000000} /* (30, 6, 17) {real, imag} */,
  {32'hbf54e6ec, 32'h00000000} /* (30, 6, 16) {real, imag} */,
  {32'hbf480c6f, 32'h00000000} /* (30, 6, 15) {real, imag} */,
  {32'hbf8aab9c, 32'h00000000} /* (30, 6, 14) {real, imag} */,
  {32'hbedf25ca, 32'h00000000} /* (30, 6, 13) {real, imag} */,
  {32'hbf26dfe7, 32'h00000000} /* (30, 6, 12) {real, imag} */,
  {32'hbf95bb82, 32'h00000000} /* (30, 6, 11) {real, imag} */,
  {32'h3e4ed2b3, 32'h00000000} /* (30, 6, 10) {real, imag} */,
  {32'h3f8f949c, 32'h00000000} /* (30, 6, 9) {real, imag} */,
  {32'h3f2e3407, 32'h00000000} /* (30, 6, 8) {real, imag} */,
  {32'h3f8ee108, 32'h00000000} /* (30, 6, 7) {real, imag} */,
  {32'h3f85dad4, 32'h00000000} /* (30, 6, 6) {real, imag} */,
  {32'h3f63c4c9, 32'h00000000} /* (30, 6, 5) {real, imag} */,
  {32'h3f0ccd99, 32'h00000000} /* (30, 6, 4) {real, imag} */,
  {32'h3f494326, 32'h00000000} /* (30, 6, 3) {real, imag} */,
  {32'h3fa08439, 32'h00000000} /* (30, 6, 2) {real, imag} */,
  {32'h3f7bcb21, 32'h00000000} /* (30, 6, 1) {real, imag} */,
  {32'h3ede7f90, 32'h00000000} /* (30, 6, 0) {real, imag} */,
  {32'h3ef5c8b0, 32'h00000000} /* (30, 5, 31) {real, imag} */,
  {32'h3f4475a2, 32'h00000000} /* (30, 5, 30) {real, imag} */,
  {32'h3f9c7cf9, 32'h00000000} /* (30, 5, 29) {real, imag} */,
  {32'h3fa45fe7, 32'h00000000} /* (30, 5, 28) {real, imag} */,
  {32'h3ecba68b, 32'h00000000} /* (30, 5, 27) {real, imag} */,
  {32'h3f2aaa0a, 32'h00000000} /* (30, 5, 26) {real, imag} */,
  {32'h3f363619, 32'h00000000} /* (30, 5, 25) {real, imag} */,
  {32'h3f8bf38b, 32'h00000000} /* (30, 5, 24) {real, imag} */,
  {32'h3f6af738, 32'h00000000} /* (30, 5, 23) {real, imag} */,
  {32'h3f530d3c, 32'h00000000} /* (30, 5, 22) {real, imag} */,
  {32'h3f787b77, 32'h00000000} /* (30, 5, 21) {real, imag} */,
  {32'h3f354093, 32'h00000000} /* (30, 5, 20) {real, imag} */,
  {32'h3edee3eb, 32'h00000000} /* (30, 5, 19) {real, imag} */,
  {32'h3dec382a, 32'h00000000} /* (30, 5, 18) {real, imag} */,
  {32'hbe077c76, 32'h00000000} /* (30, 5, 17) {real, imag} */,
  {32'hbca5c8f3, 32'h00000000} /* (30, 5, 16) {real, imag} */,
  {32'hbf44ff22, 32'h00000000} /* (30, 5, 15) {real, imag} */,
  {32'hbf54006d, 32'h00000000} /* (30, 5, 14) {real, imag} */,
  {32'hbf2f546e, 32'h00000000} /* (30, 5, 13) {real, imag} */,
  {32'hbf551fb6, 32'h00000000} /* (30, 5, 12) {real, imag} */,
  {32'hbf9a6fe7, 32'h00000000} /* (30, 5, 11) {real, imag} */,
  {32'hbf160484, 32'h00000000} /* (30, 5, 10) {real, imag} */,
  {32'hbdae44c7, 32'h00000000} /* (30, 5, 9) {real, imag} */,
  {32'hbe68456c, 32'h00000000} /* (30, 5, 8) {real, imag} */,
  {32'hbda2e95f, 32'h00000000} /* (30, 5, 7) {real, imag} */,
  {32'h3dea2946, 32'h00000000} /* (30, 5, 6) {real, imag} */,
  {32'h3f2f2faa, 32'h00000000} /* (30, 5, 5) {real, imag} */,
  {32'h3f7ab68b, 32'h00000000} /* (30, 5, 4) {real, imag} */,
  {32'h3f51ba22, 32'h00000000} /* (30, 5, 3) {real, imag} */,
  {32'h3f7a01bc, 32'h00000000} /* (30, 5, 2) {real, imag} */,
  {32'h3f6b6264, 32'h00000000} /* (30, 5, 1) {real, imag} */,
  {32'h3eff32de, 32'h00000000} /* (30, 5, 0) {real, imag} */,
  {32'h3e406cf4, 32'h00000000} /* (30, 4, 31) {real, imag} */,
  {32'h3e931399, 32'h00000000} /* (30, 4, 30) {real, imag} */,
  {32'h3f16d284, 32'h00000000} /* (30, 4, 29) {real, imag} */,
  {32'h3f948bed, 32'h00000000} /* (30, 4, 28) {real, imag} */,
  {32'h3f7313f5, 32'h00000000} /* (30, 4, 27) {real, imag} */,
  {32'h3f8054b6, 32'h00000000} /* (30, 4, 26) {real, imag} */,
  {32'h3f37d734, 32'h00000000} /* (30, 4, 25) {real, imag} */,
  {32'h3f21f5bc, 32'h00000000} /* (30, 4, 24) {real, imag} */,
  {32'h3f1e755d, 32'h00000000} /* (30, 4, 23) {real, imag} */,
  {32'h3f4af0a4, 32'h00000000} /* (30, 4, 22) {real, imag} */,
  {32'h3f8a5596, 32'h00000000} /* (30, 4, 21) {real, imag} */,
  {32'h3f9b16ca, 32'h00000000} /* (30, 4, 20) {real, imag} */,
  {32'h3f6291b5, 32'h00000000} /* (30, 4, 19) {real, imag} */,
  {32'h3f2d36ea, 32'h00000000} /* (30, 4, 18) {real, imag} */,
  {32'h3f26eefb, 32'h00000000} /* (30, 4, 17) {real, imag} */,
  {32'h3ed6f0e4, 32'h00000000} /* (30, 4, 16) {real, imag} */,
  {32'hbf34807b, 32'h00000000} /* (30, 4, 15) {real, imag} */,
  {32'hbf195bb3, 32'h00000000} /* (30, 4, 14) {real, imag} */,
  {32'hbf15c0bc, 32'h00000000} /* (30, 4, 13) {real, imag} */,
  {32'hbf667543, 32'h00000000} /* (30, 4, 12) {real, imag} */,
  {32'hbfb19283, 32'h00000000} /* (30, 4, 11) {real, imag} */,
  {32'hbfc3162d, 32'h00000000} /* (30, 4, 10) {real, imag} */,
  {32'hbf6c3572, 32'h00000000} /* (30, 4, 9) {real, imag} */,
  {32'hbf1b3259, 32'h00000000} /* (30, 4, 8) {real, imag} */,
  {32'hbedc84dc, 32'h00000000} /* (30, 4, 7) {real, imag} */,
  {32'hbddf3c9d, 32'h00000000} /* (30, 4, 6) {real, imag} */,
  {32'h3f37e8bb, 32'h00000000} /* (30, 4, 5) {real, imag} */,
  {32'h3f766c51, 32'h00000000} /* (30, 4, 4) {real, imag} */,
  {32'h3f6e0d68, 32'h00000000} /* (30, 4, 3) {real, imag} */,
  {32'h3f3d941d, 32'h00000000} /* (30, 4, 2) {real, imag} */,
  {32'h3f14b8cc, 32'h00000000} /* (30, 4, 1) {real, imag} */,
  {32'h3ecfbd3c, 32'h00000000} /* (30, 4, 0) {real, imag} */,
  {32'h3eba9b19, 32'h00000000} /* (30, 3, 31) {real, imag} */,
  {32'h3f4c6370, 32'h00000000} /* (30, 3, 30) {real, imag} */,
  {32'h3f60fb86, 32'h00000000} /* (30, 3, 29) {real, imag} */,
  {32'h3f1aa26a, 32'h00000000} /* (30, 3, 28) {real, imag} */,
  {32'h3f7cb813, 32'h00000000} /* (30, 3, 27) {real, imag} */,
  {32'h3fba07ee, 32'h00000000} /* (30, 3, 26) {real, imag} */,
  {32'h3f86df9c, 32'h00000000} /* (30, 3, 25) {real, imag} */,
  {32'h3f45cc0c, 32'h00000000} /* (30, 3, 24) {real, imag} */,
  {32'h3f034012, 32'h00000000} /* (30, 3, 23) {real, imag} */,
  {32'h3f87f98c, 32'h00000000} /* (30, 3, 22) {real, imag} */,
  {32'h3fa2bebb, 32'h00000000} /* (30, 3, 21) {real, imag} */,
  {32'h3f6e2cfb, 32'h00000000} /* (30, 3, 20) {real, imag} */,
  {32'h3ed55c6f, 32'h00000000} /* (30, 3, 19) {real, imag} */,
  {32'h3ed05736, 32'h00000000} /* (30, 3, 18) {real, imag} */,
  {32'h3f3364bc, 32'h00000000} /* (30, 3, 17) {real, imag} */,
  {32'h3df6c982, 32'h00000000} /* (30, 3, 16) {real, imag} */,
  {32'hbf41d596, 32'h00000000} /* (30, 3, 15) {real, imag} */,
  {32'hbf3d1a25, 32'h00000000} /* (30, 3, 14) {real, imag} */,
  {32'hbf0dab24, 32'h00000000} /* (30, 3, 13) {real, imag} */,
  {32'hbfc934c9, 32'h00000000} /* (30, 3, 12) {real, imag} */,
  {32'hbfc3b56d, 32'h00000000} /* (30, 3, 11) {real, imag} */,
  {32'hbfa6fc0e, 32'h00000000} /* (30, 3, 10) {real, imag} */,
  {32'hbf285b57, 32'h00000000} /* (30, 3, 9) {real, imag} */,
  {32'hbf328918, 32'h00000000} /* (30, 3, 8) {real, imag} */,
  {32'hbf8a232d, 32'h00000000} /* (30, 3, 7) {real, imag} */,
  {32'hbf51644f, 32'h00000000} /* (30, 3, 6) {real, imag} */,
  {32'hbd276950, 32'h00000000} /* (30, 3, 5) {real, imag} */,
  {32'h3f37dc4e, 32'h00000000} /* (30, 3, 4) {real, imag} */,
  {32'h3f48daba, 32'h00000000} /* (30, 3, 3) {real, imag} */,
  {32'h3f9547fc, 32'h00000000} /* (30, 3, 2) {real, imag} */,
  {32'h3f368b8e, 32'h00000000} /* (30, 3, 1) {real, imag} */,
  {32'h3ea6b3f9, 32'h00000000} /* (30, 3, 0) {real, imag} */,
  {32'h3ed68635, 32'h00000000} /* (30, 2, 31) {real, imag} */,
  {32'h3f8f66e8, 32'h00000000} /* (30, 2, 30) {real, imag} */,
  {32'h3f91e698, 32'h00000000} /* (30, 2, 29) {real, imag} */,
  {32'h3f5d929f, 32'h00000000} /* (30, 2, 28) {real, imag} */,
  {32'h3f476e05, 32'h00000000} /* (30, 2, 27) {real, imag} */,
  {32'h3faa655f, 32'h00000000} /* (30, 2, 26) {real, imag} */,
  {32'h3f5d3367, 32'h00000000} /* (30, 2, 25) {real, imag} */,
  {32'h3f3c414f, 32'h00000000} /* (30, 2, 24) {real, imag} */,
  {32'h3e9b1567, 32'h00000000} /* (30, 2, 23) {real, imag} */,
  {32'h3f297ba4, 32'h00000000} /* (30, 2, 22) {real, imag} */,
  {32'h3f8127a3, 32'h00000000} /* (30, 2, 21) {real, imag} */,
  {32'h3f30c769, 32'h00000000} /* (30, 2, 20) {real, imag} */,
  {32'h3ec81368, 32'h00000000} /* (30, 2, 19) {real, imag} */,
  {32'h3e570283, 32'h00000000} /* (30, 2, 18) {real, imag} */,
  {32'h3f11223e, 32'h00000000} /* (30, 2, 17) {real, imag} */,
  {32'hbe0d66f6, 32'h00000000} /* (30, 2, 16) {real, imag} */,
  {32'hbf6d5da7, 32'h00000000} /* (30, 2, 15) {real, imag} */,
  {32'hbf0e85b8, 32'h00000000} /* (30, 2, 14) {real, imag} */,
  {32'hbebeb2cb, 32'h00000000} /* (30, 2, 13) {real, imag} */,
  {32'hbf92bceb, 32'h00000000} /* (30, 2, 12) {real, imag} */,
  {32'hbfa56011, 32'h00000000} /* (30, 2, 11) {real, imag} */,
  {32'hbf8c40b1, 32'h00000000} /* (30, 2, 10) {real, imag} */,
  {32'hbf71a7c3, 32'h00000000} /* (30, 2, 9) {real, imag} */,
  {32'hbf4b3cbe, 32'h00000000} /* (30, 2, 8) {real, imag} */,
  {32'hbfb3bd42, 32'h00000000} /* (30, 2, 7) {real, imag} */,
  {32'hbfbbc5e3, 32'h00000000} /* (30, 2, 6) {real, imag} */,
  {32'hbea63da7, 32'h00000000} /* (30, 2, 5) {real, imag} */,
  {32'h3f2205f6, 32'h00000000} /* (30, 2, 4) {real, imag} */,
  {32'h3f4997d1, 32'h00000000} /* (30, 2, 3) {real, imag} */,
  {32'h3f18aff0, 32'h00000000} /* (30, 2, 2) {real, imag} */,
  {32'h3eaa5b7a, 32'h00000000} /* (30, 2, 1) {real, imag} */,
  {32'h3e3c23ca, 32'h00000000} /* (30, 2, 0) {real, imag} */,
  {32'h3ea2ae65, 32'h00000000} /* (30, 1, 31) {real, imag} */,
  {32'h3f2b189a, 32'h00000000} /* (30, 1, 30) {real, imag} */,
  {32'h3f1b20f5, 32'h00000000} /* (30, 1, 29) {real, imag} */,
  {32'h3f275dd2, 32'h00000000} /* (30, 1, 28) {real, imag} */,
  {32'h3f314ba4, 32'h00000000} /* (30, 1, 27) {real, imag} */,
  {32'h3f4fbc40, 32'h00000000} /* (30, 1, 26) {real, imag} */,
  {32'h3f791d2f, 32'h00000000} /* (30, 1, 25) {real, imag} */,
  {32'h3f54290a, 32'h00000000} /* (30, 1, 24) {real, imag} */,
  {32'h3e8f6c42, 32'h00000000} /* (30, 1, 23) {real, imag} */,
  {32'h3f407817, 32'h00000000} /* (30, 1, 22) {real, imag} */,
  {32'h3f4ead91, 32'h00000000} /* (30, 1, 21) {real, imag} */,
  {32'h3ee9d850, 32'h00000000} /* (30, 1, 20) {real, imag} */,
  {32'h3f2141fc, 32'h00000000} /* (30, 1, 19) {real, imag} */,
  {32'h3f35af87, 32'h00000000} /* (30, 1, 18) {real, imag} */,
  {32'h3f9404cf, 32'h00000000} /* (30, 1, 17) {real, imag} */,
  {32'h3d7d7599, 32'h00000000} /* (30, 1, 16) {real, imag} */,
  {32'hbf65eeda, 32'h00000000} /* (30, 1, 15) {real, imag} */,
  {32'hbf1bc624, 32'h00000000} /* (30, 1, 14) {real, imag} */,
  {32'hbead61f3, 32'h00000000} /* (30, 1, 13) {real, imag} */,
  {32'hbf222dfa, 32'h00000000} /* (30, 1, 12) {real, imag} */,
  {32'hbfa53c9f, 32'h00000000} /* (30, 1, 11) {real, imag} */,
  {32'hbf8178e2, 32'h00000000} /* (30, 1, 10) {real, imag} */,
  {32'hbf599f2a, 32'h00000000} /* (30, 1, 9) {real, imag} */,
  {32'hbf5c7402, 32'h00000000} /* (30, 1, 8) {real, imag} */,
  {32'hbf69024c, 32'h00000000} /* (30, 1, 7) {real, imag} */,
  {32'hbf9bd61c, 32'h00000000} /* (30, 1, 6) {real, imag} */,
  {32'hbde1efd2, 32'h00000000} /* (30, 1, 5) {real, imag} */,
  {32'h3f503937, 32'h00000000} /* (30, 1, 4) {real, imag} */,
  {32'h3f80d578, 32'h00000000} /* (30, 1, 3) {real, imag} */,
  {32'h3f29cabf, 32'h00000000} /* (30, 1, 2) {real, imag} */,
  {32'h3e1f2c26, 32'h00000000} /* (30, 1, 1) {real, imag} */,
  {32'h3d70ea7e, 32'h00000000} /* (30, 1, 0) {real, imag} */,
  {32'h3e90c9e5, 32'h00000000} /* (30, 0, 31) {real, imag} */,
  {32'h3e901815, 32'h00000000} /* (30, 0, 30) {real, imag} */,
  {32'h3e84a190, 32'h00000000} /* (30, 0, 29) {real, imag} */,
  {32'h3eb472a4, 32'h00000000} /* (30, 0, 28) {real, imag} */,
  {32'h3eb83cee, 32'h00000000} /* (30, 0, 27) {real, imag} */,
  {32'h3ee86cdb, 32'h00000000} /* (30, 0, 26) {real, imag} */,
  {32'h3f3148aa, 32'h00000000} /* (30, 0, 25) {real, imag} */,
  {32'h3ed38b92, 32'h00000000} /* (30, 0, 24) {real, imag} */,
  {32'h3e8c65a4, 32'h00000000} /* (30, 0, 23) {real, imag} */,
  {32'h3f26d490, 32'h00000000} /* (30, 0, 22) {real, imag} */,
  {32'h3f255e5d, 32'h00000000} /* (30, 0, 21) {real, imag} */,
  {32'h3e678644, 32'h00000000} /* (30, 0, 20) {real, imag} */,
  {32'h3ea0a3f3, 32'h00000000} /* (30, 0, 19) {real, imag} */,
  {32'h3f0e515a, 32'h00000000} /* (30, 0, 18) {real, imag} */,
  {32'h3f56d3d6, 32'h00000000} /* (30, 0, 17) {real, imag} */,
  {32'h3dc178a2, 32'h00000000} /* (30, 0, 16) {real, imag} */,
  {32'hbef728e1, 32'h00000000} /* (30, 0, 15) {real, imag} */,
  {32'hbf5dcceb, 32'h00000000} /* (30, 0, 14) {real, imag} */,
  {32'hbf59d5aa, 32'h00000000} /* (30, 0, 13) {real, imag} */,
  {32'hbecb9d14, 32'h00000000} /* (30, 0, 12) {real, imag} */,
  {32'hbef282d2, 32'h00000000} /* (30, 0, 11) {real, imag} */,
  {32'hbeafc88a, 32'h00000000} /* (30, 0, 10) {real, imag} */,
  {32'hbe73d79f, 32'h00000000} /* (30, 0, 9) {real, imag} */,
  {32'hbef39358, 32'h00000000} /* (30, 0, 8) {real, imag} */,
  {32'hbf2e82ae, 32'h00000000} /* (30, 0, 7) {real, imag} */,
  {32'hbee017a5, 32'h00000000} /* (30, 0, 6) {real, imag} */,
  {32'h3e47581c, 32'h00000000} /* (30, 0, 5) {real, imag} */,
  {32'h3f0e1061, 32'h00000000} /* (30, 0, 4) {real, imag} */,
  {32'h3f0b6b55, 32'h00000000} /* (30, 0, 3) {real, imag} */,
  {32'h3ed58f63, 32'h00000000} /* (30, 0, 2) {real, imag} */,
  {32'h3dfa65e6, 32'h00000000} /* (30, 0, 1) {real, imag} */,
  {32'h3d7900e4, 32'h00000000} /* (30, 0, 0) {real, imag} */,
  {32'h3b6ee1f5, 32'h00000000} /* (29, 31, 31) {real, imag} */,
  {32'h3e450260, 32'h00000000} /* (29, 31, 30) {real, imag} */,
  {32'h3f2c0bf2, 32'h00000000} /* (29, 31, 29) {real, imag} */,
  {32'h3ed5da36, 32'h00000000} /* (29, 31, 28) {real, imag} */,
  {32'h3eae199f, 32'h00000000} /* (29, 31, 27) {real, imag} */,
  {32'h3eba73d7, 32'h00000000} /* (29, 31, 26) {real, imag} */,
  {32'h3eeee131, 32'h00000000} /* (29, 31, 25) {real, imag} */,
  {32'h3f037742, 32'h00000000} /* (29, 31, 24) {real, imag} */,
  {32'h3ec822fb, 32'h00000000} /* (29, 31, 23) {real, imag} */,
  {32'h3eca2cac, 32'h00000000} /* (29, 31, 22) {real, imag} */,
  {32'h3e826b5a, 32'h00000000} /* (29, 31, 21) {real, imag} */,
  {32'h3aff3f40, 32'h00000000} /* (29, 31, 20) {real, imag} */,
  {32'h3cf72032, 32'h00000000} /* (29, 31, 19) {real, imag} */,
  {32'hbe21beb7, 32'h00000000} /* (29, 31, 18) {real, imag} */,
  {32'hbe4f2fc7, 32'h00000000} /* (29, 31, 17) {real, imag} */,
  {32'hbe93f9a2, 32'h00000000} /* (29, 31, 16) {real, imag} */,
  {32'hbe4d9817, 32'h00000000} /* (29, 31, 15) {real, imag} */,
  {32'hbed8a96a, 32'h00000000} /* (29, 31, 14) {real, imag} */,
  {32'hbf139d5e, 32'h00000000} /* (29, 31, 13) {real, imag} */,
  {32'hbf3f61d1, 32'h00000000} /* (29, 31, 12) {real, imag} */,
  {32'hbf050d20, 32'h00000000} /* (29, 31, 11) {real, imag} */,
  {32'h3dcf412b, 32'h00000000} /* (29, 31, 10) {real, imag} */,
  {32'h3f33786d, 32'h00000000} /* (29, 31, 9) {real, imag} */,
  {32'h3ed51f5f, 32'h00000000} /* (29, 31, 8) {real, imag} */,
  {32'h3ea136fd, 32'h00000000} /* (29, 31, 7) {real, imag} */,
  {32'h3ec36218, 32'h00000000} /* (29, 31, 6) {real, imag} */,
  {32'h3e8b6479, 32'h00000000} /* (29, 31, 5) {real, imag} */,
  {32'h3ef22b24, 32'h00000000} /* (29, 31, 4) {real, imag} */,
  {32'h3f154ad0, 32'h00000000} /* (29, 31, 3) {real, imag} */,
  {32'h3f2103d9, 32'h00000000} /* (29, 31, 2) {real, imag} */,
  {32'h3f2a293e, 32'h00000000} /* (29, 31, 1) {real, imag} */,
  {32'h3e8ae892, 32'h00000000} /* (29, 31, 0) {real, imag} */,
  {32'h3e96b47c, 32'h00000000} /* (29, 30, 31) {real, imag} */,
  {32'h3f122bba, 32'h00000000} /* (29, 30, 30) {real, imag} */,
  {32'h3f485c16, 32'h00000000} /* (29, 30, 29) {real, imag} */,
  {32'h3f70c78e, 32'h00000000} /* (29, 30, 28) {real, imag} */,
  {32'h3f80f1d8, 32'h00000000} /* (29, 30, 27) {real, imag} */,
  {32'h3f82a2ec, 32'h00000000} /* (29, 30, 26) {real, imag} */,
  {32'h3fb1e2d9, 32'h00000000} /* (29, 30, 25) {real, imag} */,
  {32'h3f8ed572, 32'h00000000} /* (29, 30, 24) {real, imag} */,
  {32'h3f8d1ddb, 32'h00000000} /* (29, 30, 23) {real, imag} */,
  {32'h3f3f010d, 32'h00000000} /* (29, 30, 22) {real, imag} */,
  {32'h3f1d9565, 32'h00000000} /* (29, 30, 21) {real, imag} */,
  {32'hbe8d97f4, 32'h00000000} /* (29, 30, 20) {real, imag} */,
  {32'hbe443624, 32'h00000000} /* (29, 30, 19) {real, imag} */,
  {32'hbf1c8f17, 32'h00000000} /* (29, 30, 18) {real, imag} */,
  {32'hbf7b14bf, 32'h00000000} /* (29, 30, 17) {real, imag} */,
  {32'hbf2ccb63, 32'h00000000} /* (29, 30, 16) {real, imag} */,
  {32'hbf12c07c, 32'h00000000} /* (29, 30, 15) {real, imag} */,
  {32'hbf9110a9, 32'h00000000} /* (29, 30, 14) {real, imag} */,
  {32'hbf999782, 32'h00000000} /* (29, 30, 13) {real, imag} */,
  {32'hbf9550ac, 32'h00000000} /* (29, 30, 12) {real, imag} */,
  {32'hbf5aaf3b, 32'h00000000} /* (29, 30, 11) {real, imag} */,
  {32'h3d9985df, 32'h00000000} /* (29, 30, 10) {real, imag} */,
  {32'h3fb83c1b, 32'h00000000} /* (29, 30, 9) {real, imag} */,
  {32'h3f831ecc, 32'h00000000} /* (29, 30, 8) {real, imag} */,
  {32'h3f0a95a8, 32'h00000000} /* (29, 30, 7) {real, imag} */,
  {32'h3f6053c9, 32'h00000000} /* (29, 30, 6) {real, imag} */,
  {32'h3f239383, 32'h00000000} /* (29, 30, 5) {real, imag} */,
  {32'h3f838800, 32'h00000000} /* (29, 30, 4) {real, imag} */,
  {32'h3fb0bf74, 32'h00000000} /* (29, 30, 3) {real, imag} */,
  {32'h3f6e83ef, 32'h00000000} /* (29, 30, 2) {real, imag} */,
  {32'h3fa11daa, 32'h00000000} /* (29, 30, 1) {real, imag} */,
  {32'h3f48df83, 32'h00000000} /* (29, 30, 0) {real, imag} */,
  {32'h3f7864bf, 32'h00000000} /* (29, 29, 31) {real, imag} */,
  {32'h3f9a358e, 32'h00000000} /* (29, 29, 30) {real, imag} */,
  {32'h3f24f4da, 32'h00000000} /* (29, 29, 29) {real, imag} */,
  {32'h3f217587, 32'h00000000} /* (29, 29, 28) {real, imag} */,
  {32'h3f2e53b5, 32'h00000000} /* (29, 29, 27) {real, imag} */,
  {32'h3f76eff7, 32'h00000000} /* (29, 29, 26) {real, imag} */,
  {32'h3fa33e3f, 32'h00000000} /* (29, 29, 25) {real, imag} */,
  {32'h3f9b8509, 32'h00000000} /* (29, 29, 24) {real, imag} */,
  {32'h3fa31145, 32'h00000000} /* (29, 29, 23) {real, imag} */,
  {32'h3f306570, 32'h00000000} /* (29, 29, 22) {real, imag} */,
  {32'h3ea5c947, 32'h00000000} /* (29, 29, 21) {real, imag} */,
  {32'hbf9dda9b, 32'h00000000} /* (29, 29, 20) {real, imag} */,
  {32'hbf2b7c9b, 32'h00000000} /* (29, 29, 19) {real, imag} */,
  {32'hbf532c5a, 32'h00000000} /* (29, 29, 18) {real, imag} */,
  {32'hbfa60593, 32'h00000000} /* (29, 29, 17) {real, imag} */,
  {32'hbf53f26a, 32'h00000000} /* (29, 29, 16) {real, imag} */,
  {32'hbf76bf31, 32'h00000000} /* (29, 29, 15) {real, imag} */,
  {32'hc0032d62, 32'h00000000} /* (29, 29, 14) {real, imag} */,
  {32'hbfd82bb3, 32'h00000000} /* (29, 29, 13) {real, imag} */,
  {32'hbf638c1f, 32'h00000000} /* (29, 29, 12) {real, imag} */,
  {32'hbeca630d, 32'h00000000} /* (29, 29, 11) {real, imag} */,
  {32'h3ea8d035, 32'h00000000} /* (29, 29, 10) {real, imag} */,
  {32'h3f846a65, 32'h00000000} /* (29, 29, 9) {real, imag} */,
  {32'h3f738a46, 32'h00000000} /* (29, 29, 8) {real, imag} */,
  {32'h3f21aeb5, 32'h00000000} /* (29, 29, 7) {real, imag} */,
  {32'h3f4fb7bd, 32'h00000000} /* (29, 29, 6) {real, imag} */,
  {32'h3f45d898, 32'h00000000} /* (29, 29, 5) {real, imag} */,
  {32'h3f66c882, 32'h00000000} /* (29, 29, 4) {real, imag} */,
  {32'h3f8de665, 32'h00000000} /* (29, 29, 3) {real, imag} */,
  {32'h3ef79364, 32'h00000000} /* (29, 29, 2) {real, imag} */,
  {32'h3ee7a17e, 32'h00000000} /* (29, 29, 1) {real, imag} */,
  {32'h3f057ad0, 32'h00000000} /* (29, 29, 0) {real, imag} */,
  {32'h3f1588af, 32'h00000000} /* (29, 28, 31) {real, imag} */,
  {32'h3f9c608e, 32'h00000000} /* (29, 28, 30) {real, imag} */,
  {32'h3f8f8aaf, 32'h00000000} /* (29, 28, 29) {real, imag} */,
  {32'h3f25d11a, 32'h00000000} /* (29, 28, 28) {real, imag} */,
  {32'h3f1ee1fc, 32'h00000000} /* (29, 28, 27) {real, imag} */,
  {32'h3f868a3c, 32'h00000000} /* (29, 28, 26) {real, imag} */,
  {32'h3f6ebda3, 32'h00000000} /* (29, 28, 25) {real, imag} */,
  {32'h3f1fb3a2, 32'h00000000} /* (29, 28, 24) {real, imag} */,
  {32'h3f0f2aba, 32'h00000000} /* (29, 28, 23) {real, imag} */,
  {32'h3f6afd16, 32'h00000000} /* (29, 28, 22) {real, imag} */,
  {32'h3f7133f6, 32'h00000000} /* (29, 28, 21) {real, imag} */,
  {32'hbf07b1a9, 32'h00000000} /* (29, 28, 20) {real, imag} */,
  {32'hbf619c09, 32'h00000000} /* (29, 28, 19) {real, imag} */,
  {32'hbf497c5c, 32'h00000000} /* (29, 28, 18) {real, imag} */,
  {32'hbf3a4c8b, 32'h00000000} /* (29, 28, 17) {real, imag} */,
  {32'hbe8d5406, 32'h00000000} /* (29, 28, 16) {real, imag} */,
  {32'hbf3223b3, 32'h00000000} /* (29, 28, 15) {real, imag} */,
  {32'hbfae6a11, 32'h00000000} /* (29, 28, 14) {real, imag} */,
  {32'hbfb3eab9, 32'h00000000} /* (29, 28, 13) {real, imag} */,
  {32'hbf45bf38, 32'h00000000} /* (29, 28, 12) {real, imag} */,
  {32'hbed495f8, 32'h00000000} /* (29, 28, 11) {real, imag} */,
  {32'h3f379b02, 32'h00000000} /* (29, 28, 10) {real, imag} */,
  {32'h3fa9d410, 32'h00000000} /* (29, 28, 9) {real, imag} */,
  {32'h3fc151c7, 32'h00000000} /* (29, 28, 8) {real, imag} */,
  {32'h3fbda899, 32'h00000000} /* (29, 28, 7) {real, imag} */,
  {32'h3f6e214a, 32'h00000000} /* (29, 28, 6) {real, imag} */,
  {32'h3f1bf569, 32'h00000000} /* (29, 28, 5) {real, imag} */,
  {32'h3f2e3737, 32'h00000000} /* (29, 28, 4) {real, imag} */,
  {32'h3f4242b8, 32'h00000000} /* (29, 28, 3) {real, imag} */,
  {32'h3ed8c43a, 32'h00000000} /* (29, 28, 2) {real, imag} */,
  {32'h3e8654b7, 32'h00000000} /* (29, 28, 1) {real, imag} */,
  {32'h3f096072, 32'h00000000} /* (29, 28, 0) {real, imag} */,
  {32'h3f01622e, 32'h00000000} /* (29, 27, 31) {real, imag} */,
  {32'h3f55e95f, 32'h00000000} /* (29, 27, 30) {real, imag} */,
  {32'h3f671def, 32'h00000000} /* (29, 27, 29) {real, imag} */,
  {32'h3f35cd11, 32'h00000000} /* (29, 27, 28) {real, imag} */,
  {32'h3f913930, 32'h00000000} /* (29, 27, 27) {real, imag} */,
  {32'h3fa76950, 32'h00000000} /* (29, 27, 26) {real, imag} */,
  {32'h3f961c0e, 32'h00000000} /* (29, 27, 25) {real, imag} */,
  {32'h3f5c6484, 32'h00000000} /* (29, 27, 24) {real, imag} */,
  {32'h3eb7884b, 32'h00000000} /* (29, 27, 23) {real, imag} */,
  {32'h3f664a7e, 32'h00000000} /* (29, 27, 22) {real, imag} */,
  {32'h3f77bccc, 32'h00000000} /* (29, 27, 21) {real, imag} */,
  {32'hbeda8650, 32'h00000000} /* (29, 27, 20) {real, imag} */,
  {32'hbf90c495, 32'h00000000} /* (29, 27, 19) {real, imag} */,
  {32'hbf7440cb, 32'h00000000} /* (29, 27, 18) {real, imag} */,
  {32'hbee1fd05, 32'h00000000} /* (29, 27, 17) {real, imag} */,
  {32'hbf01dbee, 32'h00000000} /* (29, 27, 16) {real, imag} */,
  {32'hbf130171, 32'h00000000} /* (29, 27, 15) {real, imag} */,
  {32'hbf6e3b19, 32'h00000000} /* (29, 27, 14) {real, imag} */,
  {32'hbf90a911, 32'h00000000} /* (29, 27, 13) {real, imag} */,
  {32'hbeef6ace, 32'h00000000} /* (29, 27, 12) {real, imag} */,
  {32'hbe4e63b9, 32'h00000000} /* (29, 27, 11) {real, imag} */,
  {32'h3f613cf1, 32'h00000000} /* (29, 27, 10) {real, imag} */,
  {32'h3fe33ba0, 32'h00000000} /* (29, 27, 9) {real, imag} */,
  {32'h3fde9cb3, 32'h00000000} /* (29, 27, 8) {real, imag} */,
  {32'h3fe0ab29, 32'h00000000} /* (29, 27, 7) {real, imag} */,
  {32'h3fa88fae, 32'h00000000} /* (29, 27, 6) {real, imag} */,
  {32'h3f800dfd, 32'h00000000} /* (29, 27, 5) {real, imag} */,
  {32'h3f58ce3e, 32'h00000000} /* (29, 27, 4) {real, imag} */,
  {32'h3f9f58ca, 32'h00000000} /* (29, 27, 3) {real, imag} */,
  {32'h3f1e6a18, 32'h00000000} /* (29, 27, 2) {real, imag} */,
  {32'h3eb8ec4c, 32'h00000000} /* (29, 27, 1) {real, imag} */,
  {32'h3ece85ff, 32'h00000000} /* (29, 27, 0) {real, imag} */,
  {32'h3ecb251e, 32'h00000000} /* (29, 26, 31) {real, imag} */,
  {32'h3f1b3da6, 32'h00000000} /* (29, 26, 30) {real, imag} */,
  {32'h3f87c5e5, 32'h00000000} /* (29, 26, 29) {real, imag} */,
  {32'h3f62894e, 32'h00000000} /* (29, 26, 28) {real, imag} */,
  {32'h3f96437b, 32'h00000000} /* (29, 26, 27) {real, imag} */,
  {32'h3f89822d, 32'h00000000} /* (29, 26, 26) {real, imag} */,
  {32'h3f54efbd, 32'h00000000} /* (29, 26, 25) {real, imag} */,
  {32'h3f991643, 32'h00000000} /* (29, 26, 24) {real, imag} */,
  {32'h3f36428f, 32'h00000000} /* (29, 26, 23) {real, imag} */,
  {32'h3efbe507, 32'h00000000} /* (29, 26, 22) {real, imag} */,
  {32'h3e8db1f8, 32'h00000000} /* (29, 26, 21) {real, imag} */,
  {32'hbf6c53a0, 32'h00000000} /* (29, 26, 20) {real, imag} */,
  {32'hbf72865b, 32'h00000000} /* (29, 26, 19) {real, imag} */,
  {32'hbf6f3334, 32'h00000000} /* (29, 26, 18) {real, imag} */,
  {32'hbf1bf219, 32'h00000000} /* (29, 26, 17) {real, imag} */,
  {32'hbf78cf67, 32'h00000000} /* (29, 26, 16) {real, imag} */,
  {32'hbf85cacf, 32'h00000000} /* (29, 26, 15) {real, imag} */,
  {32'hbf6bb50c, 32'h00000000} /* (29, 26, 14) {real, imag} */,
  {32'hbf694710, 32'h00000000} /* (29, 26, 13) {real, imag} */,
  {32'hbf2f3c9d, 32'h00000000} /* (29, 26, 12) {real, imag} */,
  {32'hbe90e74f, 32'h00000000} /* (29, 26, 11) {real, imag} */,
  {32'h3e878e6e, 32'h00000000} /* (29, 26, 10) {real, imag} */,
  {32'h3f7dd6cd, 32'h00000000} /* (29, 26, 9) {real, imag} */,
  {32'h3f95a856, 32'h00000000} /* (29, 26, 8) {real, imag} */,
  {32'h3f6ef4ab, 32'h00000000} /* (29, 26, 7) {real, imag} */,
  {32'h3f563dcf, 32'h00000000} /* (29, 26, 6) {real, imag} */,
  {32'h3f642a47, 32'h00000000} /* (29, 26, 5) {real, imag} */,
  {32'h3f6bd795, 32'h00000000} /* (29, 26, 4) {real, imag} */,
  {32'h3fa05549, 32'h00000000} /* (29, 26, 3) {real, imag} */,
  {32'h3f2374b9, 32'h00000000} /* (29, 26, 2) {real, imag} */,
  {32'h3f058e9b, 32'h00000000} /* (29, 26, 1) {real, imag} */,
  {32'h3f0eadf0, 32'h00000000} /* (29, 26, 0) {real, imag} */,
  {32'h3f2aee9e, 32'h00000000} /* (29, 25, 31) {real, imag} */,
  {32'h3f654b4b, 32'h00000000} /* (29, 25, 30) {real, imag} */,
  {32'h3f73ca91, 32'h00000000} /* (29, 25, 29) {real, imag} */,
  {32'h3f539f47, 32'h00000000} /* (29, 25, 28) {real, imag} */,
  {32'h3f93ca49, 32'h00000000} /* (29, 25, 27) {real, imag} */,
  {32'h3facdc2e, 32'h00000000} /* (29, 25, 26) {real, imag} */,
  {32'h3fa5be12, 32'h00000000} /* (29, 25, 25) {real, imag} */,
  {32'h3f7be92d, 32'h00000000} /* (29, 25, 24) {real, imag} */,
  {32'h3f52ec3b, 32'h00000000} /* (29, 25, 23) {real, imag} */,
  {32'h3f3d3684, 32'h00000000} /* (29, 25, 22) {real, imag} */,
  {32'h3e81432c, 32'h00000000} /* (29, 25, 21) {real, imag} */,
  {32'hbf627f19, 32'h00000000} /* (29, 25, 20) {real, imag} */,
  {32'hbf2dfcd2, 32'h00000000} /* (29, 25, 19) {real, imag} */,
  {32'hbf664851, 32'h00000000} /* (29, 25, 18) {real, imag} */,
  {32'hbf14e577, 32'h00000000} /* (29, 25, 17) {real, imag} */,
  {32'hbf3d9c67, 32'h00000000} /* (29, 25, 16) {real, imag} */,
  {32'hbfacc31a, 32'h00000000} /* (29, 25, 15) {real, imag} */,
  {32'hbfe68ca4, 32'h00000000} /* (29, 25, 14) {real, imag} */,
  {32'hbfa52f97, 32'h00000000} /* (29, 25, 13) {real, imag} */,
  {32'hbf33b669, 32'h00000000} /* (29, 25, 12) {real, imag} */,
  {32'hbf0dcc74, 32'h00000000} /* (29, 25, 11) {real, imag} */,
  {32'h3e4ad0c2, 32'h00000000} /* (29, 25, 10) {real, imag} */,
  {32'h3f87a593, 32'h00000000} /* (29, 25, 9) {real, imag} */,
  {32'h3f9f072e, 32'h00000000} /* (29, 25, 8) {real, imag} */,
  {32'h3f68c5d2, 32'h00000000} /* (29, 25, 7) {real, imag} */,
  {32'h3f652443, 32'h00000000} /* (29, 25, 6) {real, imag} */,
  {32'h3f847b9d, 32'h00000000} /* (29, 25, 5) {real, imag} */,
  {32'h3f99d765, 32'h00000000} /* (29, 25, 4) {real, imag} */,
  {32'h3f2eafba, 32'h00000000} /* (29, 25, 3) {real, imag} */,
  {32'h3ed365e4, 32'h00000000} /* (29, 25, 2) {real, imag} */,
  {32'h3e86ff5a, 32'h00000000} /* (29, 25, 1) {real, imag} */,
  {32'h3ed08c7b, 32'h00000000} /* (29, 25, 0) {real, imag} */,
  {32'h3f128a91, 32'h00000000} /* (29, 24, 31) {real, imag} */,
  {32'h3f50c603, 32'h00000000} /* (29, 24, 30) {real, imag} */,
  {32'h3ebe5977, 32'h00000000} /* (29, 24, 29) {real, imag} */,
  {32'h3ece9d6c, 32'h00000000} /* (29, 24, 28) {real, imag} */,
  {32'h3f484621, 32'h00000000} /* (29, 24, 27) {real, imag} */,
  {32'h3fbfe526, 32'h00000000} /* (29, 24, 26) {real, imag} */,
  {32'h40013106, 32'h00000000} /* (29, 24, 25) {real, imag} */,
  {32'h3f9981d2, 32'h00000000} /* (29, 24, 24) {real, imag} */,
  {32'h3f5e3a61, 32'h00000000} /* (29, 24, 23) {real, imag} */,
  {32'h3f6198d0, 32'h00000000} /* (29, 24, 22) {real, imag} */,
  {32'h3f071691, 32'h00000000} /* (29, 24, 21) {real, imag} */,
  {32'hbf6f15c9, 32'h00000000} /* (29, 24, 20) {real, imag} */,
  {32'hbf8c6459, 32'h00000000} /* (29, 24, 19) {real, imag} */,
  {32'hbfa84e51, 32'h00000000} /* (29, 24, 18) {real, imag} */,
  {32'hbf6fccb6, 32'h00000000} /* (29, 24, 17) {real, imag} */,
  {32'hbf82252d, 32'h00000000} /* (29, 24, 16) {real, imag} */,
  {32'hbf92c089, 32'h00000000} /* (29, 24, 15) {real, imag} */,
  {32'hbfe0b376, 32'h00000000} /* (29, 24, 14) {real, imag} */,
  {32'hbf8953bb, 32'h00000000} /* (29, 24, 13) {real, imag} */,
  {32'hbed277a5, 32'h00000000} /* (29, 24, 12) {real, imag} */,
  {32'hbf0d55e5, 32'h00000000} /* (29, 24, 11) {real, imag} */,
  {32'h3e8653d1, 32'h00000000} /* (29, 24, 10) {real, imag} */,
  {32'h3f9e0e8d, 32'h00000000} /* (29, 24, 9) {real, imag} */,
  {32'h3fea8965, 32'h00000000} /* (29, 24, 8) {real, imag} */,
  {32'h3fdf8d46, 32'h00000000} /* (29, 24, 7) {real, imag} */,
  {32'h3fd2b476, 32'h00000000} /* (29, 24, 6) {real, imag} */,
  {32'h3f87b0db, 32'h00000000} /* (29, 24, 5) {real, imag} */,
  {32'h3f5355f9, 32'h00000000} /* (29, 24, 4) {real, imag} */,
  {32'h3f951940, 32'h00000000} /* (29, 24, 3) {real, imag} */,
  {32'h3f936d16, 32'h00000000} /* (29, 24, 2) {real, imag} */,
  {32'h3efe4f4b, 32'h00000000} /* (29, 24, 1) {real, imag} */,
  {32'h3e61d35e, 32'h00000000} /* (29, 24, 0) {real, imag} */,
  {32'h3f14f2cd, 32'h00000000} /* (29, 23, 31) {real, imag} */,
  {32'h3f06015f, 32'h00000000} /* (29, 23, 30) {real, imag} */,
  {32'h3ec94c17, 32'h00000000} /* (29, 23, 29) {real, imag} */,
  {32'h3ebe5c61, 32'h00000000} /* (29, 23, 28) {real, imag} */,
  {32'h3f174612, 32'h00000000} /* (29, 23, 27) {real, imag} */,
  {32'h3fb4295c, 32'h00000000} /* (29, 23, 26) {real, imag} */,
  {32'h3f949c07, 32'h00000000} /* (29, 23, 25) {real, imag} */,
  {32'h3f10d8f2, 32'h00000000} /* (29, 23, 24) {real, imag} */,
  {32'h3f48f700, 32'h00000000} /* (29, 23, 23) {real, imag} */,
  {32'h3f7642c6, 32'h00000000} /* (29, 23, 22) {real, imag} */,
  {32'h3f294779, 32'h00000000} /* (29, 23, 21) {real, imag} */,
  {32'hbf21aa95, 32'h00000000} /* (29, 23, 20) {real, imag} */,
  {32'hbf9bea74, 32'h00000000} /* (29, 23, 19) {real, imag} */,
  {32'hbfea0912, 32'h00000000} /* (29, 23, 18) {real, imag} */,
  {32'hbf69c618, 32'h00000000} /* (29, 23, 17) {real, imag} */,
  {32'hbf4ec180, 32'h00000000} /* (29, 23, 16) {real, imag} */,
  {32'hbf1cf08e, 32'h00000000} /* (29, 23, 15) {real, imag} */,
  {32'hbf66abf8, 32'h00000000} /* (29, 23, 14) {real, imag} */,
  {32'hbf19d3da, 32'h00000000} /* (29, 23, 13) {real, imag} */,
  {32'hbec8d664, 32'h00000000} /* (29, 23, 12) {real, imag} */,
  {32'hbf0478dd, 32'h00000000} /* (29, 23, 11) {real, imag} */,
  {32'hbd84d601, 32'h00000000} /* (29, 23, 10) {real, imag} */,
  {32'h3f25cd1c, 32'h00000000} /* (29, 23, 9) {real, imag} */,
  {32'h3fb1a95b, 32'h00000000} /* (29, 23, 8) {real, imag} */,
  {32'h3fbccfba, 32'h00000000} /* (29, 23, 7) {real, imag} */,
  {32'h3faa0f4a, 32'h00000000} /* (29, 23, 6) {real, imag} */,
  {32'h3f90cc64, 32'h00000000} /* (29, 23, 5) {real, imag} */,
  {32'h3f6ecb57, 32'h00000000} /* (29, 23, 4) {real, imag} */,
  {32'h3f969905, 32'h00000000} /* (29, 23, 3) {real, imag} */,
  {32'h3f82ab3a, 32'h00000000} /* (29, 23, 2) {real, imag} */,
  {32'h3f214311, 32'h00000000} /* (29, 23, 1) {real, imag} */,
  {32'h3e8e3710, 32'h00000000} /* (29, 23, 0) {real, imag} */,
  {32'h3f01a716, 32'h00000000} /* (29, 22, 31) {real, imag} */,
  {32'h3f0897c0, 32'h00000000} /* (29, 22, 30) {real, imag} */,
  {32'h3f31339f, 32'h00000000} /* (29, 22, 29) {real, imag} */,
  {32'h3eedbb45, 32'h00000000} /* (29, 22, 28) {real, imag} */,
  {32'h3eac281f, 32'h00000000} /* (29, 22, 27) {real, imag} */,
  {32'h3f53d55d, 32'h00000000} /* (29, 22, 26) {real, imag} */,
  {32'h3f2fe892, 32'h00000000} /* (29, 22, 25) {real, imag} */,
  {32'h3f50cd4a, 32'h00000000} /* (29, 22, 24) {real, imag} */,
  {32'h3f9188bc, 32'h00000000} /* (29, 22, 23) {real, imag} */,
  {32'h3f8edb14, 32'h00000000} /* (29, 22, 22) {real, imag} */,
  {32'h3f0c940f, 32'h00000000} /* (29, 22, 21) {real, imag} */,
  {32'hbf38004d, 32'h00000000} /* (29, 22, 20) {real, imag} */,
  {32'hbf019326, 32'h00000000} /* (29, 22, 19) {real, imag} */,
  {32'hbf157701, 32'h00000000} /* (29, 22, 18) {real, imag} */,
  {32'hbeee6e7e, 32'h00000000} /* (29, 22, 17) {real, imag} */,
  {32'hbf0bfcc7, 32'h00000000} /* (29, 22, 16) {real, imag} */,
  {32'hbf189b28, 32'h00000000} /* (29, 22, 15) {real, imag} */,
  {32'hbf2a4b5f, 32'h00000000} /* (29, 22, 14) {real, imag} */,
  {32'hbf43ebab, 32'h00000000} /* (29, 22, 13) {real, imag} */,
  {32'hbf166955, 32'h00000000} /* (29, 22, 12) {real, imag} */,
  {32'hbf1ab52b, 32'h00000000} /* (29, 22, 11) {real, imag} */,
  {32'h3ad4ed8d, 32'h00000000} /* (29, 22, 10) {real, imag} */,
  {32'h3e8045ce, 32'h00000000} /* (29, 22, 9) {real, imag} */,
  {32'h3f28b070, 32'h00000000} /* (29, 22, 8) {real, imag} */,
  {32'h3f92d9a6, 32'h00000000} /* (29, 22, 7) {real, imag} */,
  {32'h3f743d98, 32'h00000000} /* (29, 22, 6) {real, imag} */,
  {32'h3f9643a2, 32'h00000000} /* (29, 22, 5) {real, imag} */,
  {32'h3f997459, 32'h00000000} /* (29, 22, 4) {real, imag} */,
  {32'h3f9945f3, 32'h00000000} /* (29, 22, 3) {real, imag} */,
  {32'h3fbf8731, 32'h00000000} /* (29, 22, 2) {real, imag} */,
  {32'h3f95be6e, 32'h00000000} /* (29, 22, 1) {real, imag} */,
  {32'h3ed859db, 32'h00000000} /* (29, 22, 0) {real, imag} */,
  {32'h3e549272, 32'h00000000} /* (29, 21, 31) {real, imag} */,
  {32'h3ebb9b18, 32'h00000000} /* (29, 21, 30) {real, imag} */,
  {32'h3ec5862e, 32'h00000000} /* (29, 21, 29) {real, imag} */,
  {32'hbc85eb46, 32'h00000000} /* (29, 21, 28) {real, imag} */,
  {32'hbe1d05a9, 32'h00000000} /* (29, 21, 27) {real, imag} */,
  {32'hbe286fef, 32'h00000000} /* (29, 21, 26) {real, imag} */,
  {32'h3d8a9a6c, 32'h00000000} /* (29, 21, 25) {real, imag} */,
  {32'h3f0ecbad, 32'h00000000} /* (29, 21, 24) {real, imag} */,
  {32'h3e72ee71, 32'h00000000} /* (29, 21, 23) {real, imag} */,
  {32'h3e2e33e8, 32'h00000000} /* (29, 21, 22) {real, imag} */,
  {32'h3e3823c9, 32'h00000000} /* (29, 21, 21) {real, imag} */,
  {32'hbe8d57a0, 32'h00000000} /* (29, 21, 20) {real, imag} */,
  {32'hbe8641b4, 32'h00000000} /* (29, 21, 19) {real, imag} */,
  {32'hbd4984cd, 32'h00000000} /* (29, 21, 18) {real, imag} */,
  {32'hbe90cf59, 32'h00000000} /* (29, 21, 17) {real, imag} */,
  {32'hbf0080ec, 32'h00000000} /* (29, 21, 16) {real, imag} */,
  {32'hbf54c390, 32'h00000000} /* (29, 21, 15) {real, imag} */,
  {32'hbf30f543, 32'h00000000} /* (29, 21, 14) {real, imag} */,
  {32'hbe584494, 32'h00000000} /* (29, 21, 13) {real, imag} */,
  {32'h3df1bc67, 32'h00000000} /* (29, 21, 12) {real, imag} */,
  {32'h3e1c43b4, 32'h00000000} /* (29, 21, 11) {real, imag} */,
  {32'h3ee4c16a, 32'h00000000} /* (29, 21, 10) {real, imag} */,
  {32'h3ec235bd, 32'h00000000} /* (29, 21, 9) {real, imag} */,
  {32'h3dd38985, 32'h00000000} /* (29, 21, 8) {real, imag} */,
  {32'h3eef3b6a, 32'h00000000} /* (29, 21, 7) {real, imag} */,
  {32'hbda19917, 32'h00000000} /* (29, 21, 6) {real, imag} */,
  {32'hbe00af3d, 32'h00000000} /* (29, 21, 5) {real, imag} */,
  {32'h3eae207d, 32'h00000000} /* (29, 21, 4) {real, imag} */,
  {32'h3e6bdaa5, 32'h00000000} /* (29, 21, 3) {real, imag} */,
  {32'h3ed040dd, 32'h00000000} /* (29, 21, 2) {real, imag} */,
  {32'h3eed26ce, 32'h00000000} /* (29, 21, 1) {real, imag} */,
  {32'h3e696689, 32'h00000000} /* (29, 21, 0) {real, imag} */,
  {32'hbe7f8e32, 32'h00000000} /* (29, 20, 31) {real, imag} */,
  {32'hbe8f2103, 32'h00000000} /* (29, 20, 30) {real, imag} */,
  {32'hbf40c993, 32'h00000000} /* (29, 20, 29) {real, imag} */,
  {32'hbf8a3612, 32'h00000000} /* (29, 20, 28) {real, imag} */,
  {32'hbf51a093, 32'h00000000} /* (29, 20, 27) {real, imag} */,
  {32'hbf3fc6ce, 32'h00000000} /* (29, 20, 26) {real, imag} */,
  {32'hbf552b52, 32'h00000000} /* (29, 20, 25) {real, imag} */,
  {32'hbf7abd89, 32'h00000000} /* (29, 20, 24) {real, imag} */,
  {32'hbf2c99b0, 32'h00000000} /* (29, 20, 23) {real, imag} */,
  {32'hbf21fcb4, 32'h00000000} /* (29, 20, 22) {real, imag} */,
  {32'h3d14c81f, 32'h00000000} /* (29, 20, 21) {real, imag} */,
  {32'h3f1e82a1, 32'h00000000} /* (29, 20, 20) {real, imag} */,
  {32'h3f1adf39, 32'h00000000} /* (29, 20, 19) {real, imag} */,
  {32'h3f40927f, 32'h00000000} /* (29, 20, 18) {real, imag} */,
  {32'h3f27c84d, 32'h00000000} /* (29, 20, 17) {real, imag} */,
  {32'h3ef21566, 32'h00000000} /* (29, 20, 16) {real, imag} */,
  {32'h3ef2d9cf, 32'h00000000} /* (29, 20, 15) {real, imag} */,
  {32'h3f382a76, 32'h00000000} /* (29, 20, 14) {real, imag} */,
  {32'h3f8606a7, 32'h00000000} /* (29, 20, 13) {real, imag} */,
  {32'h3f3dcd24, 32'h00000000} /* (29, 20, 12) {real, imag} */,
  {32'h3efa4b8a, 32'h00000000} /* (29, 20, 11) {real, imag} */,
  {32'hbc749e96, 32'h00000000} /* (29, 20, 10) {real, imag} */,
  {32'hbedf46bf, 32'h00000000} /* (29, 20, 9) {real, imag} */,
  {32'hbf39af61, 32'h00000000} /* (29, 20, 8) {real, imag} */,
  {32'hbf2b66b8, 32'h00000000} /* (29, 20, 7) {real, imag} */,
  {32'hbf9689f4, 32'h00000000} /* (29, 20, 6) {real, imag} */,
  {32'hbfa4cd96, 32'h00000000} /* (29, 20, 5) {real, imag} */,
  {32'hbf83c730, 32'h00000000} /* (29, 20, 4) {real, imag} */,
  {32'hbfad5f7e, 32'h00000000} /* (29, 20, 3) {real, imag} */,
  {32'hbfaae262, 32'h00000000} /* (29, 20, 2) {real, imag} */,
  {32'hbf379f69, 32'h00000000} /* (29, 20, 1) {real, imag} */,
  {32'hbd09d924, 32'h00000000} /* (29, 20, 0) {real, imag} */,
  {32'hbf5a3816, 32'h00000000} /* (29, 19, 31) {real, imag} */,
  {32'hbf53f9b2, 32'h00000000} /* (29, 19, 30) {real, imag} */,
  {32'hbf9a4507, 32'h00000000} /* (29, 19, 29) {real, imag} */,
  {32'hbf853d21, 32'h00000000} /* (29, 19, 28) {real, imag} */,
  {32'hbf414330, 32'h00000000} /* (29, 19, 27) {real, imag} */,
  {32'hbef7b231, 32'h00000000} /* (29, 19, 26) {real, imag} */,
  {32'hbf09ad00, 32'h00000000} /* (29, 19, 25) {real, imag} */,
  {32'hbf0086c9, 32'h00000000} /* (29, 19, 24) {real, imag} */,
  {32'hbf4088ba, 32'h00000000} /* (29, 19, 23) {real, imag} */,
  {32'hbf92e28e, 32'h00000000} /* (29, 19, 22) {real, imag} */,
  {32'h3c23afbc, 32'h00000000} /* (29, 19, 21) {real, imag} */,
  {32'h3f7aefbc, 32'h00000000} /* (29, 19, 20) {real, imag} */,
  {32'h3f69b3ce, 32'h00000000} /* (29, 19, 19) {real, imag} */,
  {32'h3f603ead, 32'h00000000} /* (29, 19, 18) {real, imag} */,
  {32'h3f6a5a34, 32'h00000000} /* (29, 19, 17) {real, imag} */,
  {32'h3f4419e0, 32'h00000000} /* (29, 19, 16) {real, imag} */,
  {32'h3f446e03, 32'h00000000} /* (29, 19, 15) {real, imag} */,
  {32'h3f847488, 32'h00000000} /* (29, 19, 14) {real, imag} */,
  {32'h3f9ffe0e, 32'h00000000} /* (29, 19, 13) {real, imag} */,
  {32'h3f8f1421, 32'h00000000} /* (29, 19, 12) {real, imag} */,
  {32'h3f63e4fc, 32'h00000000} /* (29, 19, 11) {real, imag} */,
  {32'hbe0ba171, 32'h00000000} /* (29, 19, 10) {real, imag} */,
  {32'hbf846012, 32'h00000000} /* (29, 19, 9) {real, imag} */,
  {32'hbfa99d9d, 32'h00000000} /* (29, 19, 8) {real, imag} */,
  {32'hbf952a7f, 32'h00000000} /* (29, 19, 7) {real, imag} */,
  {32'hbf401075, 32'h00000000} /* (29, 19, 6) {real, imag} */,
  {32'hbf7c9edb, 32'h00000000} /* (29, 19, 5) {real, imag} */,
  {32'hbf823aa1, 32'h00000000} /* (29, 19, 4) {real, imag} */,
  {32'hbf4dfe90, 32'h00000000} /* (29, 19, 3) {real, imag} */,
  {32'hbfa21c94, 32'h00000000} /* (29, 19, 2) {real, imag} */,
  {32'hbf99f553, 32'h00000000} /* (29, 19, 1) {real, imag} */,
  {32'hbf3dbde3, 32'h00000000} /* (29, 19, 0) {real, imag} */,
  {32'hbf848eae, 32'h00000000} /* (29, 18, 31) {real, imag} */,
  {32'hbf84552d, 32'h00000000} /* (29, 18, 30) {real, imag} */,
  {32'hbf7603f4, 32'h00000000} /* (29, 18, 29) {real, imag} */,
  {32'hbf8dc54a, 32'h00000000} /* (29, 18, 28) {real, imag} */,
  {32'hbfa4b44d, 32'h00000000} /* (29, 18, 27) {real, imag} */,
  {32'hbf807cdd, 32'h00000000} /* (29, 18, 26) {real, imag} */,
  {32'hbedb4ab3, 32'h00000000} /* (29, 18, 25) {real, imag} */,
  {32'hbec08786, 32'h00000000} /* (29, 18, 24) {real, imag} */,
  {32'hbf9318f0, 32'h00000000} /* (29, 18, 23) {real, imag} */,
  {32'hbfb12fb9, 32'h00000000} /* (29, 18, 22) {real, imag} */,
  {32'hbf39ab6b, 32'h00000000} /* (29, 18, 21) {real, imag} */,
  {32'h3ef13232, 32'h00000000} /* (29, 18, 20) {real, imag} */,
  {32'h3f87ce47, 32'h00000000} /* (29, 18, 19) {real, imag} */,
  {32'h3fb746ab, 32'h00000000} /* (29, 18, 18) {real, imag} */,
  {32'h3f5dc512, 32'h00000000} /* (29, 18, 17) {real, imag} */,
  {32'h3f513582, 32'h00000000} /* (29, 18, 16) {real, imag} */,
  {32'h3f51609e, 32'h00000000} /* (29, 18, 15) {real, imag} */,
  {32'h3f7765cc, 32'h00000000} /* (29, 18, 14) {real, imag} */,
  {32'h3f5a397c, 32'h00000000} /* (29, 18, 13) {real, imag} */,
  {32'h3f66522f, 32'h00000000} /* (29, 18, 12) {real, imag} */,
  {32'h3f39d8c9, 32'h00000000} /* (29, 18, 11) {real, imag} */,
  {32'hbf1d2c5d, 32'h00000000} /* (29, 18, 10) {real, imag} */,
  {32'hbfbd53bc, 32'h00000000} /* (29, 18, 9) {real, imag} */,
  {32'hbf84c617, 32'h00000000} /* (29, 18, 8) {real, imag} */,
  {32'hbf2c7e3a, 32'h00000000} /* (29, 18, 7) {real, imag} */,
  {32'hbf033477, 32'h00000000} /* (29, 18, 6) {real, imag} */,
  {32'hbf282fca, 32'h00000000} /* (29, 18, 5) {real, imag} */,
  {32'hbf8f6a19, 32'h00000000} /* (29, 18, 4) {real, imag} */,
  {32'hbf91da42, 32'h00000000} /* (29, 18, 3) {real, imag} */,
  {32'hbf9223e5, 32'h00000000} /* (29, 18, 2) {real, imag} */,
  {32'hbfa2fba7, 32'h00000000} /* (29, 18, 1) {real, imag} */,
  {32'hbf964df2, 32'h00000000} /* (29, 18, 0) {real, imag} */,
  {32'hbf4986ab, 32'h00000000} /* (29, 17, 31) {real, imag} */,
  {32'hbfcabc89, 32'h00000000} /* (29, 17, 30) {real, imag} */,
  {32'hbf9ba528, 32'h00000000} /* (29, 17, 29) {real, imag} */,
  {32'hbfc736f6, 32'h00000000} /* (29, 17, 28) {real, imag} */,
  {32'hbfd7ad1f, 32'h00000000} /* (29, 17, 27) {real, imag} */,
  {32'hbfaad9b0, 32'h00000000} /* (29, 17, 26) {real, imag} */,
  {32'hbf446bdc, 32'h00000000} /* (29, 17, 25) {real, imag} */,
  {32'hbf533609, 32'h00000000} /* (29, 17, 24) {real, imag} */,
  {32'hbf9a0f82, 32'h00000000} /* (29, 17, 23) {real, imag} */,
  {32'hbf9268b2, 32'h00000000} /* (29, 17, 22) {real, imag} */,
  {32'hbfa5c074, 32'h00000000} /* (29, 17, 21) {real, imag} */,
  {32'hbd3642b2, 32'h00000000} /* (29, 17, 20) {real, imag} */,
  {32'h3f1294cf, 32'h00000000} /* (29, 17, 19) {real, imag} */,
  {32'h3f5d1543, 32'h00000000} /* (29, 17, 18) {real, imag} */,
  {32'h3faeb362, 32'h00000000} /* (29, 17, 17) {real, imag} */,
  {32'h3f6ef79b, 32'h00000000} /* (29, 17, 16) {real, imag} */,
  {32'h3f81a9a4, 32'h00000000} /* (29, 17, 15) {real, imag} */,
  {32'h3fa3df25, 32'h00000000} /* (29, 17, 14) {real, imag} */,
  {32'h3f0b4ed3, 32'h00000000} /* (29, 17, 13) {real, imag} */,
  {32'h3f147e16, 32'h00000000} /* (29, 17, 12) {real, imag} */,
  {32'h3ed87903, 32'h00000000} /* (29, 17, 11) {real, imag} */,
  {32'hbea0e4af, 32'h00000000} /* (29, 17, 10) {real, imag} */,
  {32'hbf2ed039, 32'h00000000} /* (29, 17, 9) {real, imag} */,
  {32'hbf8418bf, 32'h00000000} /* (29, 17, 8) {real, imag} */,
  {32'hbf5812ab, 32'h00000000} /* (29, 17, 7) {real, imag} */,
  {32'hbf3dc207, 32'h00000000} /* (29, 17, 6) {real, imag} */,
  {32'hbed5c8c8, 32'h00000000} /* (29, 17, 5) {real, imag} */,
  {32'hbf723113, 32'h00000000} /* (29, 17, 4) {real, imag} */,
  {32'hbf9ce642, 32'h00000000} /* (29, 17, 3) {real, imag} */,
  {32'hbf6fc7ba, 32'h00000000} /* (29, 17, 2) {real, imag} */,
  {32'hbf5e4046, 32'h00000000} /* (29, 17, 1) {real, imag} */,
  {32'hbef15de1, 32'h00000000} /* (29, 17, 0) {real, imag} */,
  {32'hbed831d3, 32'h00000000} /* (29, 16, 31) {real, imag} */,
  {32'hbfa45aaa, 32'h00000000} /* (29, 16, 30) {real, imag} */,
  {32'hbf727e3e, 32'h00000000} /* (29, 16, 29) {real, imag} */,
  {32'hbf91028b, 32'h00000000} /* (29, 16, 28) {real, imag} */,
  {32'hbfb4bd75, 32'h00000000} /* (29, 16, 27) {real, imag} */,
  {32'hbf361ea3, 32'h00000000} /* (29, 16, 26) {real, imag} */,
  {32'hbf621a41, 32'h00000000} /* (29, 16, 25) {real, imag} */,
  {32'hbfa9f35c, 32'h00000000} /* (29, 16, 24) {real, imag} */,
  {32'hbf640dc2, 32'h00000000} /* (29, 16, 23) {real, imag} */,
  {32'hbf2914bb, 32'h00000000} /* (29, 16, 22) {real, imag} */,
  {32'hbf400de2, 32'h00000000} /* (29, 16, 21) {real, imag} */,
  {32'h3f03a6db, 32'h00000000} /* (29, 16, 20) {real, imag} */,
  {32'h3f3f2847, 32'h00000000} /* (29, 16, 19) {real, imag} */,
  {32'h3f112123, 32'h00000000} /* (29, 16, 18) {real, imag} */,
  {32'h3f7ab9b0, 32'h00000000} /* (29, 16, 17) {real, imag} */,
  {32'h3f9bca9d, 32'h00000000} /* (29, 16, 16) {real, imag} */,
  {32'h3fb40601, 32'h00000000} /* (29, 16, 15) {real, imag} */,
  {32'h3f88c9c6, 32'h00000000} /* (29, 16, 14) {real, imag} */,
  {32'h3f1fd3b7, 32'h00000000} /* (29, 16, 13) {real, imag} */,
  {32'h3ef1da80, 32'h00000000} /* (29, 16, 12) {real, imag} */,
  {32'h3e3924b7, 32'h00000000} /* (29, 16, 11) {real, imag} */,
  {32'hbeccecb4, 32'h00000000} /* (29, 16, 10) {real, imag} */,
  {32'hbf166b28, 32'h00000000} /* (29, 16, 9) {real, imag} */,
  {32'hbf9e26ae, 32'h00000000} /* (29, 16, 8) {real, imag} */,
  {32'hbf92813f, 32'h00000000} /* (29, 16, 7) {real, imag} */,
  {32'hbf82f997, 32'h00000000} /* (29, 16, 6) {real, imag} */,
  {32'hbf50048b, 32'h00000000} /* (29, 16, 5) {real, imag} */,
  {32'hbf759316, 32'h00000000} /* (29, 16, 4) {real, imag} */,
  {32'hbf8a9086, 32'h00000000} /* (29, 16, 3) {real, imag} */,
  {32'hbf79784e, 32'h00000000} /* (29, 16, 2) {real, imag} */,
  {32'hbf9ad317, 32'h00000000} /* (29, 16, 1) {real, imag} */,
  {32'hbecc29d1, 32'h00000000} /* (29, 16, 0) {real, imag} */,
  {32'hbee19186, 32'h00000000} /* (29, 15, 31) {real, imag} */,
  {32'hbf8b8a17, 32'h00000000} /* (29, 15, 30) {real, imag} */,
  {32'hbf4136da, 32'h00000000} /* (29, 15, 29) {real, imag} */,
  {32'hbf0b62fc, 32'h00000000} /* (29, 15, 28) {real, imag} */,
  {32'hbf097935, 32'h00000000} /* (29, 15, 27) {real, imag} */,
  {32'hbf042f18, 32'h00000000} /* (29, 15, 26) {real, imag} */,
  {32'hbf75403e, 32'h00000000} /* (29, 15, 25) {real, imag} */,
  {32'hbf520352, 32'h00000000} /* (29, 15, 24) {real, imag} */,
  {32'hbeb06719, 32'h00000000} /* (29, 15, 23) {real, imag} */,
  {32'hbed9a199, 32'h00000000} /* (29, 15, 22) {real, imag} */,
  {32'hbb99c8c9, 32'h00000000} /* (29, 15, 21) {real, imag} */,
  {32'h3f55583e, 32'h00000000} /* (29, 15, 20) {real, imag} */,
  {32'h3f1552f6, 32'h00000000} /* (29, 15, 19) {real, imag} */,
  {32'h3f1320e8, 32'h00000000} /* (29, 15, 18) {real, imag} */,
  {32'h3f0ecfc0, 32'h00000000} /* (29, 15, 17) {real, imag} */,
  {32'h3faa535e, 32'h00000000} /* (29, 15, 16) {real, imag} */,
  {32'h3fcb368b, 32'h00000000} /* (29, 15, 15) {real, imag} */,
  {32'h3faf251e, 32'h00000000} /* (29, 15, 14) {real, imag} */,
  {32'h3f8838ce, 32'h00000000} /* (29, 15, 13) {real, imag} */,
  {32'h3f887e26, 32'h00000000} /* (29, 15, 12) {real, imag} */,
  {32'h3ed0da11, 32'h00000000} /* (29, 15, 11) {real, imag} */,
  {32'hbf3843d2, 32'h00000000} /* (29, 15, 10) {real, imag} */,
  {32'hbf7bb905, 32'h00000000} /* (29, 15, 9) {real, imag} */,
  {32'hbfaf921b, 32'h00000000} /* (29, 15, 8) {real, imag} */,
  {32'hbff9bed9, 32'h00000000} /* (29, 15, 7) {real, imag} */,
  {32'hbf9bd59d, 32'h00000000} /* (29, 15, 6) {real, imag} */,
  {32'hbf9129de, 32'h00000000} /* (29, 15, 5) {real, imag} */,
  {32'hbf2188e6, 32'h00000000} /* (29, 15, 4) {real, imag} */,
  {32'hbf3dc119, 32'h00000000} /* (29, 15, 3) {real, imag} */,
  {32'hbf35be92, 32'h00000000} /* (29, 15, 2) {real, imag} */,
  {32'hbf363142, 32'h00000000} /* (29, 15, 1) {real, imag} */,
  {32'hbea12354, 32'h00000000} /* (29, 15, 0) {real, imag} */,
  {32'hbf2b3563, 32'h00000000} /* (29, 14, 31) {real, imag} */,
  {32'hbf9cb148, 32'h00000000} /* (29, 14, 30) {real, imag} */,
  {32'hbf94d909, 32'h00000000} /* (29, 14, 29) {real, imag} */,
  {32'hbf12e133, 32'h00000000} /* (29, 14, 28) {real, imag} */,
  {32'hbe7c780f, 32'h00000000} /* (29, 14, 27) {real, imag} */,
  {32'hbea5fdaa, 32'h00000000} /* (29, 14, 26) {real, imag} */,
  {32'hbf5ca9b0, 32'h00000000} /* (29, 14, 25) {real, imag} */,
  {32'hbfb6f58f, 32'h00000000} /* (29, 14, 24) {real, imag} */,
  {32'hbf87250c, 32'h00000000} /* (29, 14, 23) {real, imag} */,
  {32'hbf90ff15, 32'h00000000} /* (29, 14, 22) {real, imag} */,
  {32'hbe782f21, 32'h00000000} /* (29, 14, 21) {real, imag} */,
  {32'h3f4f5da8, 32'h00000000} /* (29, 14, 20) {real, imag} */,
  {32'h3f23c13a, 32'h00000000} /* (29, 14, 19) {real, imag} */,
  {32'h3f1a2cb5, 32'h00000000} /* (29, 14, 18) {real, imag} */,
  {32'h3f3ab6cd, 32'h00000000} /* (29, 14, 17) {real, imag} */,
  {32'h3fa98af8, 32'h00000000} /* (29, 14, 16) {real, imag} */,
  {32'h3fa1006c, 32'h00000000} /* (29, 14, 15) {real, imag} */,
  {32'h3fabf06f, 32'h00000000} /* (29, 14, 14) {real, imag} */,
  {32'h3f74e150, 32'h00000000} /* (29, 14, 13) {real, imag} */,
  {32'h3f8da4c8, 32'h00000000} /* (29, 14, 12) {real, imag} */,
  {32'h3f7ad7fc, 32'h00000000} /* (29, 14, 11) {real, imag} */,
  {32'hbe8d578a, 32'h00000000} /* (29, 14, 10) {real, imag} */,
  {32'hbfa980d2, 32'h00000000} /* (29, 14, 9) {real, imag} */,
  {32'hbf9e841a, 32'h00000000} /* (29, 14, 8) {real, imag} */,
  {32'hbf9051af, 32'h00000000} /* (29, 14, 7) {real, imag} */,
  {32'hbf51641b, 32'h00000000} /* (29, 14, 6) {real, imag} */,
  {32'hbf92674c, 32'h00000000} /* (29, 14, 5) {real, imag} */,
  {32'hbf164145, 32'h00000000} /* (29, 14, 4) {real, imag} */,
  {32'hbf999ec4, 32'h00000000} /* (29, 14, 3) {real, imag} */,
  {32'hbf5f4e87, 32'h00000000} /* (29, 14, 2) {real, imag} */,
  {32'hbeba78e8, 32'h00000000} /* (29, 14, 1) {real, imag} */,
  {32'hbed5e14d, 32'h00000000} /* (29, 14, 0) {real, imag} */,
  {32'hbf4cd62c, 32'h00000000} /* (29, 13, 31) {real, imag} */,
  {32'hbf81a301, 32'h00000000} /* (29, 13, 30) {real, imag} */,
  {32'hbf8e513c, 32'h00000000} /* (29, 13, 29) {real, imag} */,
  {32'hbf9b8617, 32'h00000000} /* (29, 13, 28) {real, imag} */,
  {32'hbf3f67aa, 32'h00000000} /* (29, 13, 27) {real, imag} */,
  {32'hbf0a1a26, 32'h00000000} /* (29, 13, 26) {real, imag} */,
  {32'hbf9e375e, 32'h00000000} /* (29, 13, 25) {real, imag} */,
  {32'hbfd99392, 32'h00000000} /* (29, 13, 24) {real, imag} */,
  {32'hbf5f58ad, 32'h00000000} /* (29, 13, 23) {real, imag} */,
  {32'hbf890f54, 32'h00000000} /* (29, 13, 22) {real, imag} */,
  {32'hbf294ab5, 32'h00000000} /* (29, 13, 21) {real, imag} */,
  {32'h3f185857, 32'h00000000} /* (29, 13, 20) {real, imag} */,
  {32'h3fb40a4a, 32'h00000000} /* (29, 13, 19) {real, imag} */,
  {32'h3fa32248, 32'h00000000} /* (29, 13, 18) {real, imag} */,
  {32'h3f731d45, 32'h00000000} /* (29, 13, 17) {real, imag} */,
  {32'h3f8bc3fa, 32'h00000000} /* (29, 13, 16) {real, imag} */,
  {32'h3f575985, 32'h00000000} /* (29, 13, 15) {real, imag} */,
  {32'h3f3bb322, 32'h00000000} /* (29, 13, 14) {real, imag} */,
  {32'h3f5c966f, 32'h00000000} /* (29, 13, 13) {real, imag} */,
  {32'h3fa8b883, 32'h00000000} /* (29, 13, 12) {real, imag} */,
  {32'h3f7f77ac, 32'h00000000} /* (29, 13, 11) {real, imag} */,
  {32'hbeff1e13, 32'h00000000} /* (29, 13, 10) {real, imag} */,
  {32'hbfa3aa81, 32'h00000000} /* (29, 13, 9) {real, imag} */,
  {32'hbfca061c, 32'h00000000} /* (29, 13, 8) {real, imag} */,
  {32'hbf4b2ea6, 32'h00000000} /* (29, 13, 7) {real, imag} */,
  {32'hbf1a37fe, 32'h00000000} /* (29, 13, 6) {real, imag} */,
  {32'hbf87e31e, 32'h00000000} /* (29, 13, 5) {real, imag} */,
  {32'hbf6fd86d, 32'h00000000} /* (29, 13, 4) {real, imag} */,
  {32'hbfb056ea, 32'h00000000} /* (29, 13, 3) {real, imag} */,
  {32'hbf881e6d, 32'h00000000} /* (29, 13, 2) {real, imag} */,
  {32'hbf4ec3ce, 32'h00000000} /* (29, 13, 1) {real, imag} */,
  {32'hbf0cbb51, 32'h00000000} /* (29, 13, 0) {real, imag} */,
  {32'hbedaeaae, 32'h00000000} /* (29, 12, 31) {real, imag} */,
  {32'hbf171967, 32'h00000000} /* (29, 12, 30) {real, imag} */,
  {32'hbf0fa517, 32'h00000000} /* (29, 12, 29) {real, imag} */,
  {32'hbfafe54e, 32'h00000000} /* (29, 12, 28) {real, imag} */,
  {32'hbfefea7a, 32'h00000000} /* (29, 12, 27) {real, imag} */,
  {32'hbf7ad46e, 32'h00000000} /* (29, 12, 26) {real, imag} */,
  {32'hbf7c30fb, 32'h00000000} /* (29, 12, 25) {real, imag} */,
  {32'hbf89101d, 32'h00000000} /* (29, 12, 24) {real, imag} */,
  {32'hbef4e055, 32'h00000000} /* (29, 12, 23) {real, imag} */,
  {32'hbf3664bf, 32'h00000000} /* (29, 12, 22) {real, imag} */,
  {32'hbf35a696, 32'h00000000} /* (29, 12, 21) {real, imag} */,
  {32'h3f3b55de, 32'h00000000} /* (29, 12, 20) {real, imag} */,
  {32'h400c352f, 32'h00000000} /* (29, 12, 19) {real, imag} */,
  {32'h3fe1813d, 32'h00000000} /* (29, 12, 18) {real, imag} */,
  {32'h3f900d1d, 32'h00000000} /* (29, 12, 17) {real, imag} */,
  {32'h3f87f16a, 32'h00000000} /* (29, 12, 16) {real, imag} */,
  {32'h3f14993a, 32'h00000000} /* (29, 12, 15) {real, imag} */,
  {32'h3f3af028, 32'h00000000} /* (29, 12, 14) {real, imag} */,
  {32'h3f794988, 32'h00000000} /* (29, 12, 13) {real, imag} */,
  {32'h3f8d35ba, 32'h00000000} /* (29, 12, 12) {real, imag} */,
  {32'h3f8bf072, 32'h00000000} /* (29, 12, 11) {real, imag} */,
  {32'hbc91b532, 32'h00000000} /* (29, 12, 10) {real, imag} */,
  {32'hbf5e825a, 32'h00000000} /* (29, 12, 9) {real, imag} */,
  {32'hbfa4ac3f, 32'h00000000} /* (29, 12, 8) {real, imag} */,
  {32'hbf695953, 32'h00000000} /* (29, 12, 7) {real, imag} */,
  {32'hbf50cb2c, 32'h00000000} /* (29, 12, 6) {real, imag} */,
  {32'hbf6d74e1, 32'h00000000} /* (29, 12, 5) {real, imag} */,
  {32'hbf240bc4, 32'h00000000} /* (29, 12, 4) {real, imag} */,
  {32'hbf8a6229, 32'h00000000} /* (29, 12, 3) {real, imag} */,
  {32'hbfe6f679, 32'h00000000} /* (29, 12, 2) {real, imag} */,
  {32'hc0069713, 32'h00000000} /* (29, 12, 1) {real, imag} */,
  {32'hbf7002a3, 32'h00000000} /* (29, 12, 0) {real, imag} */,
  {32'hbe9307d8, 32'h00000000} /* (29, 11, 31) {real, imag} */,
  {32'hbeb7d7bc, 32'h00000000} /* (29, 11, 30) {real, imag} */,
  {32'hbebde6a8, 32'h00000000} /* (29, 11, 29) {real, imag} */,
  {32'hbf6ebce9, 32'h00000000} /* (29, 11, 28) {real, imag} */,
  {32'hbfb422b2, 32'h00000000} /* (29, 11, 27) {real, imag} */,
  {32'hbf71da0d, 32'h00000000} /* (29, 11, 26) {real, imag} */,
  {32'hbf190551, 32'h00000000} /* (29, 11, 25) {real, imag} */,
  {32'hbedfcc85, 32'h00000000} /* (29, 11, 24) {real, imag} */,
  {32'hbed0e052, 32'h00000000} /* (29, 11, 23) {real, imag} */,
  {32'hbf0d6aa3, 32'h00000000} /* (29, 11, 22) {real, imag} */,
  {32'hbf5ddb68, 32'h00000000} /* (29, 11, 21) {real, imag} */,
  {32'hbe1f9200, 32'h00000000} /* (29, 11, 20) {real, imag} */,
  {32'h3f8a8a7e, 32'h00000000} /* (29, 11, 19) {real, imag} */,
  {32'h3fabe8b8, 32'h00000000} /* (29, 11, 18) {real, imag} */,
  {32'h3f9346ef, 32'h00000000} /* (29, 11, 17) {real, imag} */,
  {32'h3f78b567, 32'h00000000} /* (29, 11, 16) {real, imag} */,
  {32'h3f04a5d9, 32'h00000000} /* (29, 11, 15) {real, imag} */,
  {32'h3f2bbd92, 32'h00000000} /* (29, 11, 14) {real, imag} */,
  {32'h3f8083d2, 32'h00000000} /* (29, 11, 13) {real, imag} */,
  {32'h3eb01af6, 32'h00000000} /* (29, 11, 12) {real, imag} */,
  {32'h3eb42106, 32'h00000000} /* (29, 11, 11) {real, imag} */,
  {32'hbe833685, 32'h00000000} /* (29, 11, 10) {real, imag} */,
  {32'hbf607b11, 32'h00000000} /* (29, 11, 9) {real, imag} */,
  {32'hbf1f9005, 32'h00000000} /* (29, 11, 8) {real, imag} */,
  {32'hbf7d97c3, 32'h00000000} /* (29, 11, 7) {real, imag} */,
  {32'hbf66fb9a, 32'h00000000} /* (29, 11, 6) {real, imag} */,
  {32'hbebd2626, 32'h00000000} /* (29, 11, 5) {real, imag} */,
  {32'hbe1b2614, 32'h00000000} /* (29, 11, 4) {real, imag} */,
  {32'hbf9f1bb1, 32'h00000000} /* (29, 11, 3) {real, imag} */,
  {32'hbfc8c2ee, 32'h00000000} /* (29, 11, 2) {real, imag} */,
  {32'hbfb30b15, 32'h00000000} /* (29, 11, 1) {real, imag} */,
  {32'hbf429efa, 32'h00000000} /* (29, 11, 0) {real, imag} */,
  {32'h3f072c60, 32'h00000000} /* (29, 10, 31) {real, imag} */,
  {32'h3f2206b4, 32'h00000000} /* (29, 10, 30) {real, imag} */,
  {32'h3f45a1e0, 32'h00000000} /* (29, 10, 29) {real, imag} */,
  {32'h3f5d801e, 32'h00000000} /* (29, 10, 28) {real, imag} */,
  {32'h3f9619da, 32'h00000000} /* (29, 10, 27) {real, imag} */,
  {32'h3eb93020, 32'h00000000} /* (29, 10, 26) {real, imag} */,
  {32'h3f2a688d, 32'h00000000} /* (29, 10, 25) {real, imag} */,
  {32'h3f389833, 32'h00000000} /* (29, 10, 24) {real, imag} */,
  {32'h3ec085d8, 32'h00000000} /* (29, 10, 23) {real, imag} */,
  {32'h3e9f4a27, 32'h00000000} /* (29, 10, 22) {real, imag} */,
  {32'hbf0d4d14, 32'h00000000} /* (29, 10, 21) {real, imag} */,
  {32'hbf952b42, 32'h00000000} /* (29, 10, 20) {real, imag} */,
  {32'hbec9ab65, 32'h00000000} /* (29, 10, 19) {real, imag} */,
  {32'hbe42044b, 32'h00000000} /* (29, 10, 18) {real, imag} */,
  {32'hbf2c300f, 32'h00000000} /* (29, 10, 17) {real, imag} */,
  {32'hbdfdf496, 32'h00000000} /* (29, 10, 16) {real, imag} */,
  {32'hbe4a414f, 32'h00000000} /* (29, 10, 15) {real, imag} */,
  {32'hbe3c9668, 32'h00000000} /* (29, 10, 14) {real, imag} */,
  {32'hbdccf49c, 32'h00000000} /* (29, 10, 13) {real, imag} */,
  {32'hbf6f836b, 32'h00000000} /* (29, 10, 12) {real, imag} */,
  {32'hbe777adf, 32'h00000000} /* (29, 10, 11) {real, imag} */,
  {32'h3ccd1a54, 32'h00000000} /* (29, 10, 10) {real, imag} */,
  {32'hbe4de039, 32'h00000000} /* (29, 10, 9) {real, imag} */,
  {32'hbde548fa, 32'h00000000} /* (29, 10, 8) {real, imag} */,
  {32'h3df35e99, 32'h00000000} /* (29, 10, 7) {real, imag} */,
  {32'h3eb0017a, 32'h00000000} /* (29, 10, 6) {real, imag} */,
  {32'h3f364cd9, 32'h00000000} /* (29, 10, 5) {real, imag} */,
  {32'h3f81029b, 32'h00000000} /* (29, 10, 4) {real, imag} */,
  {32'h3ebe24fd, 32'h00000000} /* (29, 10, 3) {real, imag} */,
  {32'h3ed7bd7d, 32'h00000000} /* (29, 10, 2) {real, imag} */,
  {32'h3f0fae8f, 32'h00000000} /* (29, 10, 1) {real, imag} */,
  {32'h3f29055e, 32'h00000000} /* (29, 10, 0) {real, imag} */,
  {32'h3f5946e2, 32'h00000000} /* (29, 9, 31) {real, imag} */,
  {32'h3fc72c28, 32'h00000000} /* (29, 9, 30) {real, imag} */,
  {32'h40012148, 32'h00000000} /* (29, 9, 29) {real, imag} */,
  {32'h3fd085fe, 32'h00000000} /* (29, 9, 28) {real, imag} */,
  {32'h3fa2929a, 32'h00000000} /* (29, 9, 27) {real, imag} */,
  {32'h3f46f88c, 32'h00000000} /* (29, 9, 26) {real, imag} */,
  {32'h3f5767d7, 32'h00000000} /* (29, 9, 25) {real, imag} */,
  {32'h3f78c595, 32'h00000000} /* (29, 9, 24) {real, imag} */,
  {32'h3f77594c, 32'h00000000} /* (29, 9, 23) {real, imag} */,
  {32'h3f657fc3, 32'h00000000} /* (29, 9, 22) {real, imag} */,
  {32'hbdccf4de, 32'h00000000} /* (29, 9, 21) {real, imag} */,
  {32'hbf8228c6, 32'h00000000} /* (29, 9, 20) {real, imag} */,
  {32'hbf3110da, 32'h00000000} /* (29, 9, 19) {real, imag} */,
  {32'hbf16489e, 32'h00000000} /* (29, 9, 18) {real, imag} */,
  {32'hbf808774, 32'h00000000} /* (29, 9, 17) {real, imag} */,
  {32'hbf7dad07, 32'h00000000} /* (29, 9, 16) {real, imag} */,
  {32'hbf8cea42, 32'h00000000} /* (29, 9, 15) {real, imag} */,
  {32'hbf4efd4c, 32'h00000000} /* (29, 9, 14) {real, imag} */,
  {32'hbf2364ac, 32'h00000000} /* (29, 9, 13) {real, imag} */,
  {32'hbfc60114, 32'h00000000} /* (29, 9, 12) {real, imag} */,
  {32'hbf729828, 32'h00000000} /* (29, 9, 11) {real, imag} */,
  {32'h3e15b317, 32'h00000000} /* (29, 9, 10) {real, imag} */,
  {32'h3ea6fac0, 32'h00000000} /* (29, 9, 9) {real, imag} */,
  {32'h3e43667f, 32'h00000000} /* (29, 9, 8) {real, imag} */,
  {32'h3f3a739f, 32'h00000000} /* (29, 9, 7) {real, imag} */,
  {32'h3f24601e, 32'h00000000} /* (29, 9, 6) {real, imag} */,
  {32'h3f72da71, 32'h00000000} /* (29, 9, 5) {real, imag} */,
  {32'h3fc6ab1f, 32'h00000000} /* (29, 9, 4) {real, imag} */,
  {32'h3fc92e13, 32'h00000000} /* (29, 9, 3) {real, imag} */,
  {32'h3f6c37ff, 32'h00000000} /* (29, 9, 2) {real, imag} */,
  {32'h3f6d93a6, 32'h00000000} /* (29, 9, 1) {real, imag} */,
  {32'h3f5616ab, 32'h00000000} /* (29, 9, 0) {real, imag} */,
  {32'h3f51a0cb, 32'h00000000} /* (29, 8, 31) {real, imag} */,
  {32'h3fc8144d, 32'h00000000} /* (29, 8, 30) {real, imag} */,
  {32'h3fbde631, 32'h00000000} /* (29, 8, 29) {real, imag} */,
  {32'h3f05797b, 32'h00000000} /* (29, 8, 28) {real, imag} */,
  {32'h3f1515f8, 32'h00000000} /* (29, 8, 27) {real, imag} */,
  {32'h3f50e691, 32'h00000000} /* (29, 8, 26) {real, imag} */,
  {32'h3ec83d88, 32'h00000000} /* (29, 8, 25) {real, imag} */,
  {32'h3ec4ba46, 32'h00000000} /* (29, 8, 24) {real, imag} */,
  {32'h3f768135, 32'h00000000} /* (29, 8, 23) {real, imag} */,
  {32'h3f8d29bb, 32'h00000000} /* (29, 8, 22) {real, imag} */,
  {32'h3f0bf74c, 32'h00000000} /* (29, 8, 21) {real, imag} */,
  {32'hbefe9491, 32'h00000000} /* (29, 8, 20) {real, imag} */,
  {32'hbf5fc888, 32'h00000000} /* (29, 8, 19) {real, imag} */,
  {32'hbf42ed87, 32'h00000000} /* (29, 8, 18) {real, imag} */,
  {32'hbf12ce87, 32'h00000000} /* (29, 8, 17) {real, imag} */,
  {32'hbece61db, 32'h00000000} /* (29, 8, 16) {real, imag} */,
  {32'hbf1dc47c, 32'h00000000} /* (29, 8, 15) {real, imag} */,
  {32'hbfc88ea1, 32'h00000000} /* (29, 8, 14) {real, imag} */,
  {32'hbf95d9d3, 32'h00000000} /* (29, 8, 13) {real, imag} */,
  {32'hbf93d3f3, 32'h00000000} /* (29, 8, 12) {real, imag} */,
  {32'hbf850f3f, 32'h00000000} /* (29, 8, 11) {real, imag} */,
  {32'hbcffb3dc, 32'h00000000} /* (29, 8, 10) {real, imag} */,
  {32'h3ec4c307, 32'h00000000} /* (29, 8, 9) {real, imag} */,
  {32'h3ebea08d, 32'h00000000} /* (29, 8, 8) {real, imag} */,
  {32'h3e8f916b, 32'h00000000} /* (29, 8, 7) {real, imag} */,
  {32'h3f178a8d, 32'h00000000} /* (29, 8, 6) {real, imag} */,
  {32'h3f4093ca, 32'h00000000} /* (29, 8, 5) {real, imag} */,
  {32'h3fb11972, 32'h00000000} /* (29, 8, 4) {real, imag} */,
  {32'h3fc6bdbf, 32'h00000000} /* (29, 8, 3) {real, imag} */,
  {32'h3fa29b37, 32'h00000000} /* (29, 8, 2) {real, imag} */,
  {32'h3fa10ab4, 32'h00000000} /* (29, 8, 1) {real, imag} */,
  {32'h3f1b8528, 32'h00000000} /* (29, 8, 0) {real, imag} */,
  {32'h3efa7306, 32'h00000000} /* (29, 7, 31) {real, imag} */,
  {32'h3f94a8df, 32'h00000000} /* (29, 7, 30) {real, imag} */,
  {32'h3f58dfdc, 32'h00000000} /* (29, 7, 29) {real, imag} */,
  {32'h3e93fab2, 32'h00000000} /* (29, 7, 28) {real, imag} */,
  {32'h3ef2bf54, 32'h00000000} /* (29, 7, 27) {real, imag} */,
  {32'h3f5e2117, 32'h00000000} /* (29, 7, 26) {real, imag} */,
  {32'h3f4d5b7d, 32'h00000000} /* (29, 7, 25) {real, imag} */,
  {32'h3f391d6b, 32'h00000000} /* (29, 7, 24) {real, imag} */,
  {32'h3f4b6261, 32'h00000000} /* (29, 7, 23) {real, imag} */,
  {32'h3f2168e1, 32'h00000000} /* (29, 7, 22) {real, imag} */,
  {32'h3f0ae25a, 32'h00000000} /* (29, 7, 21) {real, imag} */,
  {32'hbec5756e, 32'h00000000} /* (29, 7, 20) {real, imag} */,
  {32'hbfadbeec, 32'h00000000} /* (29, 7, 19) {real, imag} */,
  {32'hbf8aaad9, 32'h00000000} /* (29, 7, 18) {real, imag} */,
  {32'hbf4570d4, 32'h00000000} /* (29, 7, 17) {real, imag} */,
  {32'hbf25c6ab, 32'h00000000} /* (29, 7, 16) {real, imag} */,
  {32'hbeeba686, 32'h00000000} /* (29, 7, 15) {real, imag} */,
  {32'hbf89f922, 32'h00000000} /* (29, 7, 14) {real, imag} */,
  {32'hbf6a099b, 32'h00000000} /* (29, 7, 13) {real, imag} */,
  {32'hbf090484, 32'h00000000} /* (29, 7, 12) {real, imag} */,
  {32'hbee424c6, 32'h00000000} /* (29, 7, 11) {real, imag} */,
  {32'h3ea0288e, 32'h00000000} /* (29, 7, 10) {real, imag} */,
  {32'h3f308ad4, 32'h00000000} /* (29, 7, 9) {real, imag} */,
  {32'h3f490230, 32'h00000000} /* (29, 7, 8) {real, imag} */,
  {32'h3e53f39d, 32'h00000000} /* (29, 7, 7) {real, imag} */,
  {32'h3ef6ce40, 32'h00000000} /* (29, 7, 6) {real, imag} */,
  {32'h3f8eba49, 32'h00000000} /* (29, 7, 5) {real, imag} */,
  {32'h3fa1da39, 32'h00000000} /* (29, 7, 4) {real, imag} */,
  {32'h3fb2bf3e, 32'h00000000} /* (29, 7, 3) {real, imag} */,
  {32'h3fc1cc04, 32'h00000000} /* (29, 7, 2) {real, imag} */,
  {32'h3f63670a, 32'h00000000} /* (29, 7, 1) {real, imag} */,
  {32'h3e3e5c44, 32'h00000000} /* (29, 7, 0) {real, imag} */,
  {32'h3f28fdf1, 32'h00000000} /* (29, 6, 31) {real, imag} */,
  {32'h3f954873, 32'h00000000} /* (29, 6, 30) {real, imag} */,
  {32'h3f96b07f, 32'h00000000} /* (29, 6, 29) {real, imag} */,
  {32'h3ef4eff4, 32'h00000000} /* (29, 6, 28) {real, imag} */,
  {32'h3f046a3b, 32'h00000000} /* (29, 6, 27) {real, imag} */,
  {32'h3f4e975e, 32'h00000000} /* (29, 6, 26) {real, imag} */,
  {32'h3f6019b2, 32'h00000000} /* (29, 6, 25) {real, imag} */,
  {32'h3f4dcff1, 32'h00000000} /* (29, 6, 24) {real, imag} */,
  {32'h3f50bd5e, 32'h00000000} /* (29, 6, 23) {real, imag} */,
  {32'h3f1dc438, 32'h00000000} /* (29, 6, 22) {real, imag} */,
  {32'h3f1e3d44, 32'h00000000} /* (29, 6, 21) {real, imag} */,
  {32'hbe562375, 32'h00000000} /* (29, 6, 20) {real, imag} */,
  {32'hbf223f23, 32'h00000000} /* (29, 6, 19) {real, imag} */,
  {32'hbf4ac7d2, 32'h00000000} /* (29, 6, 18) {real, imag} */,
  {32'hbf427b77, 32'h00000000} /* (29, 6, 17) {real, imag} */,
  {32'hbf98fa72, 32'h00000000} /* (29, 6, 16) {real, imag} */,
  {32'hbf9d3495, 32'h00000000} /* (29, 6, 15) {real, imag} */,
  {32'hbf6e8f7c, 32'h00000000} /* (29, 6, 14) {real, imag} */,
  {32'hbf46b1e6, 32'h00000000} /* (29, 6, 13) {real, imag} */,
  {32'hbf5eb2e5, 32'h00000000} /* (29, 6, 12) {real, imag} */,
  {32'hbf817cf8, 32'h00000000} /* (29, 6, 11) {real, imag} */,
  {32'h3e4f3f69, 32'h00000000} /* (29, 6, 10) {real, imag} */,
  {32'h3f2f6174, 32'h00000000} /* (29, 6, 9) {real, imag} */,
  {32'h3ea95b36, 32'h00000000} /* (29, 6, 8) {real, imag} */,
  {32'h3eb6781d, 32'h00000000} /* (29, 6, 7) {real, imag} */,
  {32'h3ee874ba, 32'h00000000} /* (29, 6, 6) {real, imag} */,
  {32'h3f978ea3, 32'h00000000} /* (29, 6, 5) {real, imag} */,
  {32'h3fa42f81, 32'h00000000} /* (29, 6, 4) {real, imag} */,
  {32'h3f483b45, 32'h00000000} /* (29, 6, 3) {real, imag} */,
  {32'h3f77686f, 32'h00000000} /* (29, 6, 2) {real, imag} */,
  {32'h3f64003f, 32'h00000000} /* (29, 6, 1) {real, imag} */,
  {32'h3eca017d, 32'h00000000} /* (29, 6, 0) {real, imag} */,
  {32'h3f227e5d, 32'h00000000} /* (29, 5, 31) {real, imag} */,
  {32'h3f94b8a4, 32'h00000000} /* (29, 5, 30) {real, imag} */,
  {32'h3fb2f473, 32'h00000000} /* (29, 5, 29) {real, imag} */,
  {32'h3f71f354, 32'h00000000} /* (29, 5, 28) {real, imag} */,
  {32'h3f3f1fab, 32'h00000000} /* (29, 5, 27) {real, imag} */,
  {32'h3f7ae55e, 32'h00000000} /* (29, 5, 26) {real, imag} */,
  {32'h3f7da940, 32'h00000000} /* (29, 5, 25) {real, imag} */,
  {32'h3f82e4ee, 32'h00000000} /* (29, 5, 24) {real, imag} */,
  {32'h3f7f653e, 32'h00000000} /* (29, 5, 23) {real, imag} */,
  {32'h3f9d1a5b, 32'h00000000} /* (29, 5, 22) {real, imag} */,
  {32'h3fe93387, 32'h00000000} /* (29, 5, 21) {real, imag} */,
  {32'h3fa30b32, 32'h00000000} /* (29, 5, 20) {real, imag} */,
  {32'h3f180f2b, 32'h00000000} /* (29, 5, 19) {real, imag} */,
  {32'h3e2744d0, 32'h00000000} /* (29, 5, 18) {real, imag} */,
  {32'h3e9526a2, 32'h00000000} /* (29, 5, 17) {real, imag} */,
  {32'hbdf97e28, 32'h00000000} /* (29, 5, 16) {real, imag} */,
  {32'hbf796d06, 32'h00000000} /* (29, 5, 15) {real, imag} */,
  {32'hbf52d0b7, 32'h00000000} /* (29, 5, 14) {real, imag} */,
  {32'hbf800da1, 32'h00000000} /* (29, 5, 13) {real, imag} */,
  {32'hbf9889a1, 32'h00000000} /* (29, 5, 12) {real, imag} */,
  {32'hbfeb82ae, 32'h00000000} /* (29, 5, 11) {real, imag} */,
  {32'hbf4a3dec, 32'h00000000} /* (29, 5, 10) {real, imag} */,
  {32'hbea3ca77, 32'h00000000} /* (29, 5, 9) {real, imag} */,
  {32'hbe423cbe, 32'h00000000} /* (29, 5, 8) {real, imag} */,
  {32'hbe2fd720, 32'h00000000} /* (29, 5, 7) {real, imag} */,
  {32'hbe1eca26, 32'h00000000} /* (29, 5, 6) {real, imag} */,
  {32'h3f576cc3, 32'h00000000} /* (29, 5, 5) {real, imag} */,
  {32'h3fc61a6a, 32'h00000000} /* (29, 5, 4) {real, imag} */,
  {32'h3f75a47e, 32'h00000000} /* (29, 5, 3) {real, imag} */,
  {32'h3f7d0772, 32'h00000000} /* (29, 5, 2) {real, imag} */,
  {32'h3f8f3f52, 32'h00000000} /* (29, 5, 1) {real, imag} */,
  {32'h3f4706be, 32'h00000000} /* (29, 5, 0) {real, imag} */,
  {32'h3ea6daaf, 32'h00000000} /* (29, 4, 31) {real, imag} */,
  {32'h3eff4b6d, 32'h00000000} /* (29, 4, 30) {real, imag} */,
  {32'h3f60ca70, 32'h00000000} /* (29, 4, 29) {real, imag} */,
  {32'h3f82645b, 32'h00000000} /* (29, 4, 28) {real, imag} */,
  {32'h3f5cd696, 32'h00000000} /* (29, 4, 27) {real, imag} */,
  {32'h3f36382f, 32'h00000000} /* (29, 4, 26) {real, imag} */,
  {32'h3f07158f, 32'h00000000} /* (29, 4, 25) {real, imag} */,
  {32'h3f1d37d8, 32'h00000000} /* (29, 4, 24) {real, imag} */,
  {32'h3f26ec5b, 32'h00000000} /* (29, 4, 23) {real, imag} */,
  {32'h3f2ac148, 32'h00000000} /* (29, 4, 22) {real, imag} */,
  {32'h3fc5e2a2, 32'h00000000} /* (29, 4, 21) {real, imag} */,
  {32'h3ffa21fc, 32'h00000000} /* (29, 4, 20) {real, imag} */,
  {32'h3fa02b09, 32'h00000000} /* (29, 4, 19) {real, imag} */,
  {32'h3fa8d103, 32'h00000000} /* (29, 4, 18) {real, imag} */,
  {32'h3f90e5f2, 32'h00000000} /* (29, 4, 17) {real, imag} */,
  {32'h3ebb3eef, 32'h00000000} /* (29, 4, 16) {real, imag} */,
  {32'hbf6f09c7, 32'h00000000} /* (29, 4, 15) {real, imag} */,
  {32'hbf796cae, 32'h00000000} /* (29, 4, 14) {real, imag} */,
  {32'hbf4708de, 32'h00000000} /* (29, 4, 13) {real, imag} */,
  {32'hbf2a5903, 32'h00000000} /* (29, 4, 12) {real, imag} */,
  {32'hbfad6b81, 32'h00000000} /* (29, 4, 11) {real, imag} */,
  {32'hbfaf8311, 32'h00000000} /* (29, 4, 10) {real, imag} */,
  {32'hbf268b9b, 32'h00000000} /* (29, 4, 9) {real, imag} */,
  {32'hbf02455d, 32'h00000000} /* (29, 4, 8) {real, imag} */,
  {32'hbf295198, 32'h00000000} /* (29, 4, 7) {real, imag} */,
  {32'hbefcffdc, 32'h00000000} /* (29, 4, 6) {real, imag} */,
  {32'h3f0f1f4c, 32'h00000000} /* (29, 4, 5) {real, imag} */,
  {32'h3fa91b3a, 32'h00000000} /* (29, 4, 4) {real, imag} */,
  {32'h3f7e7166, 32'h00000000} /* (29, 4, 3) {real, imag} */,
  {32'h3f87e878, 32'h00000000} /* (29, 4, 2) {real, imag} */,
  {32'h3f157c48, 32'h00000000} /* (29, 4, 1) {real, imag} */,
  {32'h3ee7050f, 32'h00000000} /* (29, 4, 0) {real, imag} */,
  {32'h3e7e1579, 32'h00000000} /* (29, 3, 31) {real, imag} */,
  {32'h3f32f477, 32'h00000000} /* (29, 3, 30) {real, imag} */,
  {32'h3f6a8b7a, 32'h00000000} /* (29, 3, 29) {real, imag} */,
  {32'h3f3eba8e, 32'h00000000} /* (29, 3, 28) {real, imag} */,
  {32'h3f5d7dca, 32'h00000000} /* (29, 3, 27) {real, imag} */,
  {32'h3f4483b6, 32'h00000000} /* (29, 3, 26) {real, imag} */,
  {32'h3ed6a62b, 32'h00000000} /* (29, 3, 25) {real, imag} */,
  {32'h3eb5a2ee, 32'h00000000} /* (29, 3, 24) {real, imag} */,
  {32'h3e5ce5df, 32'h00000000} /* (29, 3, 23) {real, imag} */,
  {32'h3ee1aba8, 32'h00000000} /* (29, 3, 22) {real, imag} */,
  {32'h3f508398, 32'h00000000} /* (29, 3, 21) {real, imag} */,
  {32'h3f90d34c, 32'h00000000} /* (29, 3, 20) {real, imag} */,
  {32'h3f43ddde, 32'h00000000} /* (29, 3, 19) {real, imag} */,
  {32'h3fa60a8f, 32'h00000000} /* (29, 3, 18) {real, imag} */,
  {32'h3fac797b, 32'h00000000} /* (29, 3, 17) {real, imag} */,
  {32'h3eee7a44, 32'h00000000} /* (29, 3, 16) {real, imag} */,
  {32'hbee3c3de, 32'h00000000} /* (29, 3, 15) {real, imag} */,
  {32'hbf66a73b, 32'h00000000} /* (29, 3, 14) {real, imag} */,
  {32'hbf1991a1, 32'h00000000} /* (29, 3, 13) {real, imag} */,
  {32'hbf1a8037, 32'h00000000} /* (29, 3, 12) {real, imag} */,
  {32'hbf7147b3, 32'h00000000} /* (29, 3, 11) {real, imag} */,
  {32'hbf83ebdc, 32'h00000000} /* (29, 3, 10) {real, imag} */,
  {32'hbf19358a, 32'h00000000} /* (29, 3, 9) {real, imag} */,
  {32'hbf0f25bd, 32'h00000000} /* (29, 3, 8) {real, imag} */,
  {32'hbf2de01b, 32'h00000000} /* (29, 3, 7) {real, imag} */,
  {32'hbf6eb901, 32'h00000000} /* (29, 3, 6) {real, imag} */,
  {32'hbe90e33e, 32'h00000000} /* (29, 3, 5) {real, imag} */,
  {32'h3f1ec474, 32'h00000000} /* (29, 3, 4) {real, imag} */,
  {32'h3f27b960, 32'h00000000} /* (29, 3, 3) {real, imag} */,
  {32'h3f3271db, 32'h00000000} /* (29, 3, 2) {real, imag} */,
  {32'h3e5d2fac, 32'h00000000} /* (29, 3, 1) {real, imag} */,
  {32'h3e7d0e45, 32'h00000000} /* (29, 3, 0) {real, imag} */,
  {32'h3f52f0fb, 32'h00000000} /* (29, 2, 31) {real, imag} */,
  {32'h3fbcc6f4, 32'h00000000} /* (29, 2, 30) {real, imag} */,
  {32'h3f9b8505, 32'h00000000} /* (29, 2, 29) {real, imag} */,
  {32'h3f795d71, 32'h00000000} /* (29, 2, 28) {real, imag} */,
  {32'h3f356011, 32'h00000000} /* (29, 2, 27) {real, imag} */,
  {32'h3f516b76, 32'h00000000} /* (29, 2, 26) {real, imag} */,
  {32'h3f4a1987, 32'h00000000} /* (29, 2, 25) {real, imag} */,
  {32'h3f469e7f, 32'h00000000} /* (29, 2, 24) {real, imag} */,
  {32'h3f267e16, 32'h00000000} /* (29, 2, 23) {real, imag} */,
  {32'h3f8d6c76, 32'h00000000} /* (29, 2, 22) {real, imag} */,
  {32'h3f90384c, 32'h00000000} /* (29, 2, 21) {real, imag} */,
  {32'h3f60edff, 32'h00000000} /* (29, 2, 20) {real, imag} */,
  {32'h3f02f117, 32'h00000000} /* (29, 2, 19) {real, imag} */,
  {32'h3f551a40, 32'h00000000} /* (29, 2, 18) {real, imag} */,
  {32'h3fa2bbf1, 32'h00000000} /* (29, 2, 17) {real, imag} */,
  {32'h3eb7554e, 32'h00000000} /* (29, 2, 16) {real, imag} */,
  {32'hbea5525d, 32'h00000000} /* (29, 2, 15) {real, imag} */,
  {32'hbf14ef37, 32'h00000000} /* (29, 2, 14) {real, imag} */,
  {32'hbef63029, 32'h00000000} /* (29, 2, 13) {real, imag} */,
  {32'hbf0dd796, 32'h00000000} /* (29, 2, 12) {real, imag} */,
  {32'hbf55949a, 32'h00000000} /* (29, 2, 11) {real, imag} */,
  {32'hbf955bd9, 32'h00000000} /* (29, 2, 10) {real, imag} */,
  {32'hbf92fb54, 32'h00000000} /* (29, 2, 9) {real, imag} */,
  {32'hbf234bfa, 32'h00000000} /* (29, 2, 8) {real, imag} */,
  {32'hbf4227a1, 32'h00000000} /* (29, 2, 7) {real, imag} */,
  {32'hbf9b9517, 32'h00000000} /* (29, 2, 6) {real, imag} */,
  {32'hbeffe50f, 32'h00000000} /* (29, 2, 5) {real, imag} */,
  {32'h3f15ab3f, 32'h00000000} /* (29, 2, 4) {real, imag} */,
  {32'h3f0a61ad, 32'h00000000} /* (29, 2, 3) {real, imag} */,
  {32'h3dc59719, 32'h00000000} /* (29, 2, 2) {real, imag} */,
  {32'h3e6065c4, 32'h00000000} /* (29, 2, 1) {real, imag} */,
  {32'h3ed59590, 32'h00000000} /* (29, 2, 0) {real, imag} */,
  {32'h3f11f7fc, 32'h00000000} /* (29, 1, 31) {real, imag} */,
  {32'h3f496976, 32'h00000000} /* (29, 1, 30) {real, imag} */,
  {32'h3f45d81e, 32'h00000000} /* (29, 1, 29) {real, imag} */,
  {32'h3f7474d5, 32'h00000000} /* (29, 1, 28) {real, imag} */,
  {32'h3f4afff9, 32'h00000000} /* (29, 1, 27) {real, imag} */,
  {32'h3f4314cc, 32'h00000000} /* (29, 1, 26) {real, imag} */,
  {32'h3f693636, 32'h00000000} /* (29, 1, 25) {real, imag} */,
  {32'h3f98e635, 32'h00000000} /* (29, 1, 24) {real, imag} */,
  {32'h3f9486e5, 32'h00000000} /* (29, 1, 23) {real, imag} */,
  {32'h3fa1bd5c, 32'h00000000} /* (29, 1, 22) {real, imag} */,
  {32'h3fa61d63, 32'h00000000} /* (29, 1, 21) {real, imag} */,
  {32'h3f7c4565, 32'h00000000} /* (29, 1, 20) {real, imag} */,
  {32'h3f4ff66e, 32'h00000000} /* (29, 1, 19) {real, imag} */,
  {32'h3f9b43ea, 32'h00000000} /* (29, 1, 18) {real, imag} */,
  {32'h3fc7f818, 32'h00000000} /* (29, 1, 17) {real, imag} */,
  {32'h3f16b8fd, 32'h00000000} /* (29, 1, 16) {real, imag} */,
  {32'hbee291fa, 32'h00000000} /* (29, 1, 15) {real, imag} */,
  {32'hbf4800b3, 32'h00000000} /* (29, 1, 14) {real, imag} */,
  {32'hbf77222c, 32'h00000000} /* (29, 1, 13) {real, imag} */,
  {32'hbfa979b8, 32'h00000000} /* (29, 1, 12) {real, imag} */,
  {32'hbfaf860c, 32'h00000000} /* (29, 1, 11) {real, imag} */,
  {32'hbf5bcd05, 32'h00000000} /* (29, 1, 10) {real, imag} */,
  {32'hbf7338b6, 32'h00000000} /* (29, 1, 9) {real, imag} */,
  {32'hbf1c4973, 32'h00000000} /* (29, 1, 8) {real, imag} */,
  {32'hbf270cac, 32'h00000000} /* (29, 1, 7) {real, imag} */,
  {32'hbf675836, 32'h00000000} /* (29, 1, 6) {real, imag} */,
  {32'hbda456d8, 32'h00000000} /* (29, 1, 5) {real, imag} */,
  {32'h3f58d8c1, 32'h00000000} /* (29, 1, 4) {real, imag} */,
  {32'h3f9a2672, 32'h00000000} /* (29, 1, 3) {real, imag} */,
  {32'h3f602d88, 32'h00000000} /* (29, 1, 2) {real, imag} */,
  {32'h3edbbfd3, 32'h00000000} /* (29, 1, 1) {real, imag} */,
  {32'h3e95e812, 32'h00000000} /* (29, 1, 0) {real, imag} */,
  {32'h3de70365, 32'h00000000} /* (29, 0, 31) {real, imag} */,
  {32'h3ecce20e, 32'h00000000} /* (29, 0, 30) {real, imag} */,
  {32'h3f13fe3b, 32'h00000000} /* (29, 0, 29) {real, imag} */,
  {32'h3ea909c6, 32'h00000000} /* (29, 0, 28) {real, imag} */,
  {32'h3e42e2b3, 32'h00000000} /* (29, 0, 27) {real, imag} */,
  {32'h3e2aca23, 32'h00000000} /* (29, 0, 26) {real, imag} */,
  {32'h3eb6d6a8, 32'h00000000} /* (29, 0, 25) {real, imag} */,
  {32'h3f0f536f, 32'h00000000} /* (29, 0, 24) {real, imag} */,
  {32'h3f22e1f0, 32'h00000000} /* (29, 0, 23) {real, imag} */,
  {32'h3f11d7b7, 32'h00000000} /* (29, 0, 22) {real, imag} */,
  {32'h3f306423, 32'h00000000} /* (29, 0, 21) {real, imag} */,
  {32'h3f251b87, 32'h00000000} /* (29, 0, 20) {real, imag} */,
  {32'h3f0420af, 32'h00000000} /* (29, 0, 19) {real, imag} */,
  {32'h3f4c6a8e, 32'h00000000} /* (29, 0, 18) {real, imag} */,
  {32'h3f742c89, 32'h00000000} /* (29, 0, 17) {real, imag} */,
  {32'h3ec5f5d2, 32'h00000000} /* (29, 0, 16) {real, imag} */,
  {32'hbe360ce4, 32'h00000000} /* (29, 0, 15) {real, imag} */,
  {32'hbf0b6eb2, 32'h00000000} /* (29, 0, 14) {real, imag} */,
  {32'hbf839821, 32'h00000000} /* (29, 0, 13) {real, imag} */,
  {32'hbf86f31f, 32'h00000000} /* (29, 0, 12) {real, imag} */,
  {32'hbf2e5a03, 32'h00000000} /* (29, 0, 11) {real, imag} */,
  {32'hbe2e2a0b, 32'h00000000} /* (29, 0, 10) {real, imag} */,
  {32'hbe929d03, 32'h00000000} /* (29, 0, 9) {real, imag} */,
  {32'hbe7ce47d, 32'h00000000} /* (29, 0, 8) {real, imag} */,
  {32'hbef00ee9, 32'h00000000} /* (29, 0, 7) {real, imag} */,
  {32'hbef30791, 32'h00000000} /* (29, 0, 6) {real, imag} */,
  {32'h3eb7ef80, 32'h00000000} /* (29, 0, 5) {real, imag} */,
  {32'h3f172648, 32'h00000000} /* (29, 0, 4) {real, imag} */,
  {32'h3f493a3d, 32'h00000000} /* (29, 0, 3) {real, imag} */,
  {32'h3f58c872, 32'h00000000} /* (29, 0, 2) {real, imag} */,
  {32'h3ebc864c, 32'h00000000} /* (29, 0, 1) {real, imag} */,
  {32'h3de31071, 32'h00000000} /* (29, 0, 0) {real, imag} */,
  {32'h3c8c2211, 32'h00000000} /* (28, 31, 31) {real, imag} */,
  {32'hbe0f62ba, 32'h00000000} /* (28, 31, 30) {real, imag} */,
  {32'h3e1fc1b8, 32'h00000000} /* (28, 31, 29) {real, imag} */,
  {32'h3f11b8a7, 32'h00000000} /* (28, 31, 28) {real, imag} */,
  {32'h3f575f00, 32'h00000000} /* (28, 31, 27) {real, imag} */,
  {32'h3f78297b, 32'h00000000} /* (28, 31, 26) {real, imag} */,
  {32'h3f3a2d87, 32'h00000000} /* (28, 31, 25) {real, imag} */,
  {32'h3ec78d3b, 32'h00000000} /* (28, 31, 24) {real, imag} */,
  {32'h3eef839f, 32'h00000000} /* (28, 31, 23) {real, imag} */,
  {32'h3ef196f8, 32'h00000000} /* (28, 31, 22) {real, imag} */,
  {32'h3e8c173f, 32'h00000000} /* (28, 31, 21) {real, imag} */,
  {32'hbdec5549, 32'h00000000} /* (28, 31, 20) {real, imag} */,
  {32'hbcea5a48, 32'h00000000} /* (28, 31, 19) {real, imag} */,
  {32'hbe40d50d, 32'h00000000} /* (28, 31, 18) {real, imag} */,
  {32'hbee1ff90, 32'h00000000} /* (28, 31, 17) {real, imag} */,
  {32'hbe8ec181, 32'h00000000} /* (28, 31, 16) {real, imag} */,
  {32'hbec47716, 32'h00000000} /* (28, 31, 15) {real, imag} */,
  {32'hbf129c68, 32'h00000000} /* (28, 31, 14) {real, imag} */,
  {32'hbf3e6de0, 32'h00000000} /* (28, 31, 13) {real, imag} */,
  {32'hbf543018, 32'h00000000} /* (28, 31, 12) {real, imag} */,
  {32'hbeb80967, 32'h00000000} /* (28, 31, 11) {real, imag} */,
  {32'h3e84fc9a, 32'h00000000} /* (28, 31, 10) {real, imag} */,
  {32'h3f436a26, 32'h00000000} /* (28, 31, 9) {real, imag} */,
  {32'h3f19b814, 32'h00000000} /* (28, 31, 8) {real, imag} */,
  {32'h3f07cb23, 32'h00000000} /* (28, 31, 7) {real, imag} */,
  {32'h3e8e19fb, 32'h00000000} /* (28, 31, 6) {real, imag} */,
  {32'h3ee54b26, 32'h00000000} /* (28, 31, 5) {real, imag} */,
  {32'h3f63abc9, 32'h00000000} /* (28, 31, 4) {real, imag} */,
  {32'h3f233215, 32'h00000000} /* (28, 31, 3) {real, imag} */,
  {32'h3f6435d4, 32'h00000000} /* (28, 31, 2) {real, imag} */,
  {32'h3f216a3d, 32'h00000000} /* (28, 31, 1) {real, imag} */,
  {32'h3cd03ebc, 32'h00000000} /* (28, 31, 0) {real, imag} */,
  {32'h3eb65bfa, 32'h00000000} /* (28, 30, 31) {real, imag} */,
  {32'h3dc63e79, 32'h00000000} /* (28, 30, 30) {real, imag} */,
  {32'h3e8682be, 32'h00000000} /* (28, 30, 29) {real, imag} */,
  {32'h3f9095fc, 32'h00000000} /* (28, 30, 28) {real, imag} */,
  {32'h3fbd5482, 32'h00000000} /* (28, 30, 27) {real, imag} */,
  {32'h3fb52e40, 32'h00000000} /* (28, 30, 26) {real, imag} */,
  {32'h3fbe21c3, 32'h00000000} /* (28, 30, 25) {real, imag} */,
  {32'h3f844b5f, 32'h00000000} /* (28, 30, 24) {real, imag} */,
  {32'h3f95db48, 32'h00000000} /* (28, 30, 23) {real, imag} */,
  {32'h3f4eff38, 32'h00000000} /* (28, 30, 22) {real, imag} */,
  {32'h3eb1df53, 32'h00000000} /* (28, 30, 21) {real, imag} */,
  {32'hbee12145, 32'h00000000} /* (28, 30, 20) {real, imag} */,
  {32'hbf13896d, 32'h00000000} /* (28, 30, 19) {real, imag} */,
  {32'hbf6ddfdc, 32'h00000000} /* (28, 30, 18) {real, imag} */,
  {32'hbfa30048, 32'h00000000} /* (28, 30, 17) {real, imag} */,
  {32'hbf7f62d1, 32'h00000000} /* (28, 30, 16) {real, imag} */,
  {32'hbf4b71de, 32'h00000000} /* (28, 30, 15) {real, imag} */,
  {32'hbfa3a15d, 32'h00000000} /* (28, 30, 14) {real, imag} */,
  {32'hbf8b5aa5, 32'h00000000} /* (28, 30, 13) {real, imag} */,
  {32'hbf9dec14, 32'h00000000} /* (28, 30, 12) {real, imag} */,
  {32'hbf4fd566, 32'h00000000} /* (28, 30, 11) {real, imag} */,
  {32'h3e9bfcf3, 32'h00000000} /* (28, 30, 10) {real, imag} */,
  {32'h3fb96a2d, 32'h00000000} /* (28, 30, 9) {real, imag} */,
  {32'h3f85cc2b, 32'h00000000} /* (28, 30, 8) {real, imag} */,
  {32'h3f932be7, 32'h00000000} /* (28, 30, 7) {real, imag} */,
  {32'h3f3bf55e, 32'h00000000} /* (28, 30, 6) {real, imag} */,
  {32'h3f49211d, 32'h00000000} /* (28, 30, 5) {real, imag} */,
  {32'h3fc04c97, 32'h00000000} /* (28, 30, 4) {real, imag} */,
  {32'h3fb56923, 32'h00000000} /* (28, 30, 3) {real, imag} */,
  {32'h3f75842c, 32'h00000000} /* (28, 30, 2) {real, imag} */,
  {32'h3f0dfe2b, 32'h00000000} /* (28, 30, 1) {real, imag} */,
  {32'h3e24839d, 32'h00000000} /* (28, 30, 0) {real, imag} */,
  {32'h3f24832a, 32'h00000000} /* (28, 29, 31) {real, imag} */,
  {32'h3f3c223a, 32'h00000000} /* (28, 29, 30) {real, imag} */,
  {32'h3f4375b0, 32'h00000000} /* (28, 29, 29) {real, imag} */,
  {32'h3fb421f8, 32'h00000000} /* (28, 29, 28) {real, imag} */,
  {32'h3f876300, 32'h00000000} /* (28, 29, 27) {real, imag} */,
  {32'h3f8c9a01, 32'h00000000} /* (28, 29, 26) {real, imag} */,
  {32'h3fcc2cda, 32'h00000000} /* (28, 29, 25) {real, imag} */,
  {32'h3f89bdce, 32'h00000000} /* (28, 29, 24) {real, imag} */,
  {32'h3f7398cf, 32'h00000000} /* (28, 29, 23) {real, imag} */,
  {32'h3f3c3f93, 32'h00000000} /* (28, 29, 22) {real, imag} */,
  {32'h3e27283c, 32'h00000000} /* (28, 29, 21) {real, imag} */,
  {32'hbfa7b79f, 32'h00000000} /* (28, 29, 20) {real, imag} */,
  {32'hbfcf07c1, 32'h00000000} /* (28, 29, 19) {real, imag} */,
  {32'hbf9c4c83, 32'h00000000} /* (28, 29, 18) {real, imag} */,
  {32'hbf9a0b43, 32'h00000000} /* (28, 29, 17) {real, imag} */,
  {32'hbf8f97b4, 32'h00000000} /* (28, 29, 16) {real, imag} */,
  {32'hbf6a3231, 32'h00000000} /* (28, 29, 15) {real, imag} */,
  {32'hbfc68fc8, 32'h00000000} /* (28, 29, 14) {real, imag} */,
  {32'hbf82adcb, 32'h00000000} /* (28, 29, 13) {real, imag} */,
  {32'hbf7b84ba, 32'h00000000} /* (28, 29, 12) {real, imag} */,
  {32'hbf10509b, 32'h00000000} /* (28, 29, 11) {real, imag} */,
  {32'h3eedabbb, 32'h00000000} /* (28, 29, 10) {real, imag} */,
  {32'h3f68d89a, 32'h00000000} /* (28, 29, 9) {real, imag} */,
  {32'h3f4984cd, 32'h00000000} /* (28, 29, 8) {real, imag} */,
  {32'h3f840915, 32'h00000000} /* (28, 29, 7) {real, imag} */,
  {32'h3f59ef9c, 32'h00000000} /* (28, 29, 6) {real, imag} */,
  {32'h3f5ff1d4, 32'h00000000} /* (28, 29, 5) {real, imag} */,
  {32'h3fb37e4c, 32'h00000000} /* (28, 29, 4) {real, imag} */,
  {32'h3fb52b65, 32'h00000000} /* (28, 29, 3) {real, imag} */,
  {32'h3f57f17e, 32'h00000000} /* (28, 29, 2) {real, imag} */,
  {32'h3e51d3e9, 32'h00000000} /* (28, 29, 1) {real, imag} */,
  {32'h3e0ef66c, 32'h00000000} /* (28, 29, 0) {real, imag} */,
  {32'h3ea8cbf9, 32'h00000000} /* (28, 28, 31) {real, imag} */,
  {32'h3f4de20f, 32'h00000000} /* (28, 28, 30) {real, imag} */,
  {32'h3f82457a, 32'h00000000} /* (28, 28, 29) {real, imag} */,
  {32'h3fa292d1, 32'h00000000} /* (28, 28, 28) {real, imag} */,
  {32'h3f5037ca, 32'h00000000} /* (28, 28, 27) {real, imag} */,
  {32'h3f821416, 32'h00000000} /* (28, 28, 26) {real, imag} */,
  {32'h3f6de2fa, 32'h00000000} /* (28, 28, 25) {real, imag} */,
  {32'h3f69a29c, 32'h00000000} /* (28, 28, 24) {real, imag} */,
  {32'h3f5c6f17, 32'h00000000} /* (28, 28, 23) {real, imag} */,
  {32'h3f9dafd6, 32'h00000000} /* (28, 28, 22) {real, imag} */,
  {32'h3f8445c9, 32'h00000000} /* (28, 28, 21) {real, imag} */,
  {32'hbf7249d0, 32'h00000000} /* (28, 28, 20) {real, imag} */,
  {32'hbfed02ec, 32'h00000000} /* (28, 28, 19) {real, imag} */,
  {32'hbf8cca36, 32'h00000000} /* (28, 28, 18) {real, imag} */,
  {32'hbf8452c1, 32'h00000000} /* (28, 28, 17) {real, imag} */,
  {32'hbf6149bf, 32'h00000000} /* (28, 28, 16) {real, imag} */,
  {32'hbf492bff, 32'h00000000} /* (28, 28, 15) {real, imag} */,
  {32'hbf96ee28, 32'h00000000} /* (28, 28, 14) {real, imag} */,
  {32'hbf6dab1e, 32'h00000000} /* (28, 28, 13) {real, imag} */,
  {32'hbf817183, 32'h00000000} /* (28, 28, 12) {real, imag} */,
  {32'hbf0fbaf1, 32'h00000000} /* (28, 28, 11) {real, imag} */,
  {32'h3f854135, 32'h00000000} /* (28, 28, 10) {real, imag} */,
  {32'h3fe23374, 32'h00000000} /* (28, 28, 9) {real, imag} */,
  {32'h3fae7b3b, 32'h00000000} /* (28, 28, 8) {real, imag} */,
  {32'h3f9c606b, 32'h00000000} /* (28, 28, 7) {real, imag} */,
  {32'h3f665329, 32'h00000000} /* (28, 28, 6) {real, imag} */,
  {32'h3f89db6a, 32'h00000000} /* (28, 28, 5) {real, imag} */,
  {32'h3fa94154, 32'h00000000} /* (28, 28, 4) {real, imag} */,
  {32'h3fa20c77, 32'h00000000} /* (28, 28, 3) {real, imag} */,
  {32'h3f8fc112, 32'h00000000} /* (28, 28, 2) {real, imag} */,
  {32'h3e9d092f, 32'h00000000} /* (28, 28, 1) {real, imag} */,
  {32'h3e432df7, 32'h00000000} /* (28, 28, 0) {real, imag} */,
  {32'h3e7c44a4, 32'h00000000} /* (28, 27, 31) {real, imag} */,
  {32'h3f548dba, 32'h00000000} /* (28, 27, 30) {real, imag} */,
  {32'h3faa19f2, 32'h00000000} /* (28, 27, 29) {real, imag} */,
  {32'h3fa9247f, 32'h00000000} /* (28, 27, 28) {real, imag} */,
  {32'h3f5cfba1, 32'h00000000} /* (28, 27, 27) {real, imag} */,
  {32'h3f34809d, 32'h00000000} /* (28, 27, 26) {real, imag} */,
  {32'h3f068b74, 32'h00000000} /* (28, 27, 25) {real, imag} */,
  {32'h3f3a0019, 32'h00000000} /* (28, 27, 24) {real, imag} */,
  {32'h3eddd63b, 32'h00000000} /* (28, 27, 23) {real, imag} */,
  {32'h3f9d00c4, 32'h00000000} /* (28, 27, 22) {real, imag} */,
  {32'h3fad93b5, 32'h00000000} /* (28, 27, 21) {real, imag} */,
  {32'hbed435c8, 32'h00000000} /* (28, 27, 20) {real, imag} */,
  {32'hbf81ece5, 32'h00000000} /* (28, 27, 19) {real, imag} */,
  {32'hbf8c1c61, 32'h00000000} /* (28, 27, 18) {real, imag} */,
  {32'hbf55edc4, 32'h00000000} /* (28, 27, 17) {real, imag} */,
  {32'hbf909392, 32'h00000000} /* (28, 27, 16) {real, imag} */,
  {32'hbf25a287, 32'h00000000} /* (28, 27, 15) {real, imag} */,
  {32'hbf0a12c0, 32'h00000000} /* (28, 27, 14) {real, imag} */,
  {32'hbf22245e, 32'h00000000} /* (28, 27, 13) {real, imag} */,
  {32'hbf51cd18, 32'h00000000} /* (28, 27, 12) {real, imag} */,
  {32'hbf15a6a6, 32'h00000000} /* (28, 27, 11) {real, imag} */,
  {32'h3f59344b, 32'h00000000} /* (28, 27, 10) {real, imag} */,
  {32'h3ff257d7, 32'h00000000} /* (28, 27, 9) {real, imag} */,
  {32'h3fcdd8ca, 32'h00000000} /* (28, 27, 8) {real, imag} */,
  {32'h3fd08cc0, 32'h00000000} /* (28, 27, 7) {real, imag} */,
  {32'h3f8b74ca, 32'h00000000} /* (28, 27, 6) {real, imag} */,
  {32'h3fbf7ace, 32'h00000000} /* (28, 27, 5) {real, imag} */,
  {32'h3f969762, 32'h00000000} /* (28, 27, 4) {real, imag} */,
  {32'h3f86a5e7, 32'h00000000} /* (28, 27, 3) {real, imag} */,
  {32'h3f8a553d, 32'h00000000} /* (28, 27, 2) {real, imag} */,
  {32'h3f1cb9e1, 32'h00000000} /* (28, 27, 1) {real, imag} */,
  {32'h3e8d12ad, 32'h00000000} /* (28, 27, 0) {real, imag} */,
  {32'h3f018650, 32'h00000000} /* (28, 26, 31) {real, imag} */,
  {32'h3f0b033c, 32'h00000000} /* (28, 26, 30) {real, imag} */,
  {32'h3f140ebe, 32'h00000000} /* (28, 26, 29) {real, imag} */,
  {32'h3f1765bf, 32'h00000000} /* (28, 26, 28) {real, imag} */,
  {32'h3f44de6e, 32'h00000000} /* (28, 26, 27) {real, imag} */,
  {32'h3f61ec3a, 32'h00000000} /* (28, 26, 26) {real, imag} */,
  {32'h3f0deee0, 32'h00000000} /* (28, 26, 25) {real, imag} */,
  {32'h3f63833e, 32'h00000000} /* (28, 26, 24) {real, imag} */,
  {32'h3f453ed2, 32'h00000000} /* (28, 26, 23) {real, imag} */,
  {32'h3f8bf544, 32'h00000000} /* (28, 26, 22) {real, imag} */,
  {32'h3f4160c5, 32'h00000000} /* (28, 26, 21) {real, imag} */,
  {32'hbf47fd58, 32'h00000000} /* (28, 26, 20) {real, imag} */,
  {32'hbf503c70, 32'h00000000} /* (28, 26, 19) {real, imag} */,
  {32'hbfb95430, 32'h00000000} /* (28, 26, 18) {real, imag} */,
  {32'hbf95012a, 32'h00000000} /* (28, 26, 17) {real, imag} */,
  {32'hbfb256ff, 32'h00000000} /* (28, 26, 16) {real, imag} */,
  {32'hbf7411cf, 32'h00000000} /* (28, 26, 15) {real, imag} */,
  {32'hbef875b9, 32'h00000000} /* (28, 26, 14) {real, imag} */,
  {32'hbf2a4a61, 32'h00000000} /* (28, 26, 13) {real, imag} */,
  {32'hbf26284b, 32'h00000000} /* (28, 26, 12) {real, imag} */,
  {32'hbf183473, 32'h00000000} /* (28, 26, 11) {real, imag} */,
  {32'h3e1e448f, 32'h00000000} /* (28, 26, 10) {real, imag} */,
  {32'h3fa6d558, 32'h00000000} /* (28, 26, 9) {real, imag} */,
  {32'h3fda0dce, 32'h00000000} /* (28, 26, 8) {real, imag} */,
  {32'h3f477d00, 32'h00000000} /* (28, 26, 7) {real, imag} */,
  {32'h3f066e94, 32'h00000000} /* (28, 26, 6) {real, imag} */,
  {32'h3f84f97f, 32'h00000000} /* (28, 26, 5) {real, imag} */,
  {32'h3f393db6, 32'h00000000} /* (28, 26, 4) {real, imag} */,
  {32'h3f1db44c, 32'h00000000} /* (28, 26, 3) {real, imag} */,
  {32'h3f186ecf, 32'h00000000} /* (28, 26, 2) {real, imag} */,
  {32'h3f4e0d18, 32'h00000000} /* (28, 26, 1) {real, imag} */,
  {32'h3f27c515, 32'h00000000} /* (28, 26, 0) {real, imag} */,
  {32'h3f5e24f3, 32'h00000000} /* (28, 25, 31) {real, imag} */,
  {32'h3f4e208d, 32'h00000000} /* (28, 25, 30) {real, imag} */,
  {32'h3f05ada7, 32'h00000000} /* (28, 25, 29) {real, imag} */,
  {32'h3ee96ba1, 32'h00000000} /* (28, 25, 28) {real, imag} */,
  {32'h3f51baab, 32'h00000000} /* (28, 25, 27) {real, imag} */,
  {32'h3f5c60d3, 32'h00000000} /* (28, 25, 26) {real, imag} */,
  {32'h3f6ec878, 32'h00000000} /* (28, 25, 25) {real, imag} */,
  {32'h3f70d2b5, 32'h00000000} /* (28, 25, 24) {real, imag} */,
  {32'h3fa02333, 32'h00000000} /* (28, 25, 23) {real, imag} */,
  {32'h3fb1ba12, 32'h00000000} /* (28, 25, 22) {real, imag} */,
  {32'h3ed3c588, 32'h00000000} /* (28, 25, 21) {real, imag} */,
  {32'hbf4343bf, 32'h00000000} /* (28, 25, 20) {real, imag} */,
  {32'hbee8b210, 32'h00000000} /* (28, 25, 19) {real, imag} */,
  {32'hbf479e54, 32'h00000000} /* (28, 25, 18) {real, imag} */,
  {32'hbf0847f7, 32'h00000000} /* (28, 25, 17) {real, imag} */,
  {32'hbf1326a6, 32'h00000000} /* (28, 25, 16) {real, imag} */,
  {32'hbf6b2843, 32'h00000000} /* (28, 25, 15) {real, imag} */,
  {32'hbf70876d, 32'h00000000} /* (28, 25, 14) {real, imag} */,
  {32'hbf1f38be, 32'h00000000} /* (28, 25, 13) {real, imag} */,
  {32'hbf1f53a4, 32'h00000000} /* (28, 25, 12) {real, imag} */,
  {32'hbee155a1, 32'h00000000} /* (28, 25, 11) {real, imag} */,
  {32'h3e54e7f2, 32'h00000000} /* (28, 25, 10) {real, imag} */,
  {32'h3f6788a9, 32'h00000000} /* (28, 25, 9) {real, imag} */,
  {32'h3fc8fa98, 32'h00000000} /* (28, 25, 8) {real, imag} */,
  {32'h3f3291f3, 32'h00000000} /* (28, 25, 7) {real, imag} */,
  {32'h3f1aec25, 32'h00000000} /* (28, 25, 6) {real, imag} */,
  {32'h3f9c4f6f, 32'h00000000} /* (28, 25, 5) {real, imag} */,
  {32'h3f5f004d, 32'h00000000} /* (28, 25, 4) {real, imag} */,
  {32'h3e94864c, 32'h00000000} /* (28, 25, 3) {real, imag} */,
  {32'h3e94c262, 32'h00000000} /* (28, 25, 2) {real, imag} */,
  {32'h3ee1ade9, 32'h00000000} /* (28, 25, 1) {real, imag} */,
  {32'h3f257a8f, 32'h00000000} /* (28, 25, 0) {real, imag} */,
  {32'h3e9bd17c, 32'h00000000} /* (28, 24, 31) {real, imag} */,
  {32'h3f5081f8, 32'h00000000} /* (28, 24, 30) {real, imag} */,
  {32'h3f049912, 32'h00000000} /* (28, 24, 29) {real, imag} */,
  {32'h3f07097c, 32'h00000000} /* (28, 24, 28) {real, imag} */,
  {32'h3fb0b939, 32'h00000000} /* (28, 24, 27) {real, imag} */,
  {32'h3fa9ef5f, 32'h00000000} /* (28, 24, 26) {real, imag} */,
  {32'h3fc1d4e2, 32'h00000000} /* (28, 24, 25) {real, imag} */,
  {32'h3f9b2789, 32'h00000000} /* (28, 24, 24) {real, imag} */,
  {32'h3fa6951e, 32'h00000000} /* (28, 24, 23) {real, imag} */,
  {32'h3f84547e, 32'h00000000} /* (28, 24, 22) {real, imag} */,
  {32'h3f2ade02, 32'h00000000} /* (28, 24, 21) {real, imag} */,
  {32'hbe97a0c6, 32'h00000000} /* (28, 24, 20) {real, imag} */,
  {32'hbf1fbbe4, 32'h00000000} /* (28, 24, 19) {real, imag} */,
  {32'hbf230ade, 32'h00000000} /* (28, 24, 18) {real, imag} */,
  {32'hbe9e5463, 32'h00000000} /* (28, 24, 17) {real, imag} */,
  {32'hbf572e72, 32'h00000000} /* (28, 24, 16) {real, imag} */,
  {32'hbfdd3409, 32'h00000000} /* (28, 24, 15) {real, imag} */,
  {32'hc005e123, 32'h00000000} /* (28, 24, 14) {real, imag} */,
  {32'hbf614f18, 32'h00000000} /* (28, 24, 13) {real, imag} */,
  {32'hbf092409, 32'h00000000} /* (28, 24, 12) {real, imag} */,
  {32'hbf2d9ab9, 32'h00000000} /* (28, 24, 11) {real, imag} */,
  {32'h3e7047dd, 32'h00000000} /* (28, 24, 10) {real, imag} */,
  {32'h3f9d61dc, 32'h00000000} /* (28, 24, 9) {real, imag} */,
  {32'h40038c74, 32'h00000000} /* (28, 24, 8) {real, imag} */,
  {32'h3fc006c9, 32'h00000000} /* (28, 24, 7) {real, imag} */,
  {32'h3f97d361, 32'h00000000} /* (28, 24, 6) {real, imag} */,
  {32'h3f79a625, 32'h00000000} /* (28, 24, 5) {real, imag} */,
  {32'h3f38cdf1, 32'h00000000} /* (28, 24, 4) {real, imag} */,
  {32'h3f29b995, 32'h00000000} /* (28, 24, 3) {real, imag} */,
  {32'h3f1f1b65, 32'h00000000} /* (28, 24, 2) {real, imag} */,
  {32'h3f1926fc, 32'h00000000} /* (28, 24, 1) {real, imag} */,
  {32'h3e98e70c, 32'h00000000} /* (28, 24, 0) {real, imag} */,
  {32'h3ec60078, 32'h00000000} /* (28, 23, 31) {real, imag} */,
  {32'h3f84775d, 32'h00000000} /* (28, 23, 30) {real, imag} */,
  {32'h3f748a13, 32'h00000000} /* (28, 23, 29) {real, imag} */,
  {32'h3f76a8c9, 32'h00000000} /* (28, 23, 28) {real, imag} */,
  {32'h3fdfa571, 32'h00000000} /* (28, 23, 27) {real, imag} */,
  {32'h3ff0f607, 32'h00000000} /* (28, 23, 26) {real, imag} */,
  {32'h3f8653c8, 32'h00000000} /* (28, 23, 25) {real, imag} */,
  {32'h3f689425, 32'h00000000} /* (28, 23, 24) {real, imag} */,
  {32'h3f91ca45, 32'h00000000} /* (28, 23, 23) {real, imag} */,
  {32'h3f86917e, 32'h00000000} /* (28, 23, 22) {real, imag} */,
  {32'h3f9274ad, 32'h00000000} /* (28, 23, 21) {real, imag} */,
  {32'hbd959cec, 32'h00000000} /* (28, 23, 20) {real, imag} */,
  {32'hbf69b459, 32'h00000000} /* (28, 23, 19) {real, imag} */,
  {32'hbf90f034, 32'h00000000} /* (28, 23, 18) {real, imag} */,
  {32'hbeff3521, 32'h00000000} /* (28, 23, 17) {real, imag} */,
  {32'hbf7061c9, 32'h00000000} /* (28, 23, 16) {real, imag} */,
  {32'hbfa75be3, 32'h00000000} /* (28, 23, 15) {real, imag} */,
  {32'hbfa7808c, 32'h00000000} /* (28, 23, 14) {real, imag} */,
  {32'hbec2e315, 32'h00000000} /* (28, 23, 13) {real, imag} */,
  {32'hbeddd95d, 32'h00000000} /* (28, 23, 12) {real, imag} */,
  {32'hbf36df81, 32'h00000000} /* (28, 23, 11) {real, imag} */,
  {32'h3c991b8c, 32'h00000000} /* (28, 23, 10) {real, imag} */,
  {32'h3f8d1a13, 32'h00000000} /* (28, 23, 9) {real, imag} */,
  {32'h3fc23bf0, 32'h00000000} /* (28, 23, 8) {real, imag} */,
  {32'h3faf2086, 32'h00000000} /* (28, 23, 7) {real, imag} */,
  {32'h3f740c17, 32'h00000000} /* (28, 23, 6) {real, imag} */,
  {32'h3f377e66, 32'h00000000} /* (28, 23, 5) {real, imag} */,
  {32'h3f032b79, 32'h00000000} /* (28, 23, 4) {real, imag} */,
  {32'h3f43d914, 32'h00000000} /* (28, 23, 3) {real, imag} */,
  {32'h3f237a72, 32'h00000000} /* (28, 23, 2) {real, imag} */,
  {32'h3eebec5b, 32'h00000000} /* (28, 23, 1) {real, imag} */,
  {32'h3e412dd3, 32'h00000000} /* (28, 23, 0) {real, imag} */,
  {32'h3f27555a, 32'h00000000} /* (28, 22, 31) {real, imag} */,
  {32'h3fc77cd7, 32'h00000000} /* (28, 22, 30) {real, imag} */,
  {32'h3fc21379, 32'h00000000} /* (28, 22, 29) {real, imag} */,
  {32'h3f86c1bb, 32'h00000000} /* (28, 22, 28) {real, imag} */,
  {32'h3f8ecc7a, 32'h00000000} /* (28, 22, 27) {real, imag} */,
  {32'h3f93c56d, 32'h00000000} /* (28, 22, 26) {real, imag} */,
  {32'h3efddbe7, 32'h00000000} /* (28, 22, 25) {real, imag} */,
  {32'h3f26a731, 32'h00000000} /* (28, 22, 24) {real, imag} */,
  {32'h3f5c11f5, 32'h00000000} /* (28, 22, 23) {real, imag} */,
  {32'h3f6a55fa, 32'h00000000} /* (28, 22, 22) {real, imag} */,
  {32'h3f09256e, 32'h00000000} /* (28, 22, 21) {real, imag} */,
  {32'hbebf6df5, 32'h00000000} /* (28, 22, 20) {real, imag} */,
  {32'hbef7a184, 32'h00000000} /* (28, 22, 19) {real, imag} */,
  {32'hbf005d19, 32'h00000000} /* (28, 22, 18) {real, imag} */,
  {32'hbe666fad, 32'h00000000} /* (28, 22, 17) {real, imag} */,
  {32'hbf29ff5a, 32'h00000000} /* (28, 22, 16) {real, imag} */,
  {32'hbf290884, 32'h00000000} /* (28, 22, 15) {real, imag} */,
  {32'hbf0f1de0, 32'h00000000} /* (28, 22, 14) {real, imag} */,
  {32'hbeb363c6, 32'h00000000} /* (28, 22, 13) {real, imag} */,
  {32'hbe3fbea7, 32'h00000000} /* (28, 22, 12) {real, imag} */,
  {32'hbec05afc, 32'h00000000} /* (28, 22, 11) {real, imag} */,
  {32'h3d8c86a6, 32'h00000000} /* (28, 22, 10) {real, imag} */,
  {32'h3f016624, 32'h00000000} /* (28, 22, 9) {real, imag} */,
  {32'h3f475ed1, 32'h00000000} /* (28, 22, 8) {real, imag} */,
  {32'h3f5f4058, 32'h00000000} /* (28, 22, 7) {real, imag} */,
  {32'h3f181dfe, 32'h00000000} /* (28, 22, 6) {real, imag} */,
  {32'h3f1822f4, 32'h00000000} /* (28, 22, 5) {real, imag} */,
  {32'h3f778d75, 32'h00000000} /* (28, 22, 4) {real, imag} */,
  {32'h3f82a66f, 32'h00000000} /* (28, 22, 3) {real, imag} */,
  {32'h3f32eea6, 32'h00000000} /* (28, 22, 2) {real, imag} */,
  {32'h3f3fdd71, 32'h00000000} /* (28, 22, 1) {real, imag} */,
  {32'h3ee15c5b, 32'h00000000} /* (28, 22, 0) {real, imag} */,
  {32'h3db95193, 32'h00000000} /* (28, 21, 31) {real, imag} */,
  {32'h3e97841e, 32'h00000000} /* (28, 21, 30) {real, imag} */,
  {32'h3f53915d, 32'h00000000} /* (28, 21, 29) {real, imag} */,
  {32'h3eef15bc, 32'h00000000} /* (28, 21, 28) {real, imag} */,
  {32'h3e76dab0, 32'h00000000} /* (28, 21, 27) {real, imag} */,
  {32'h3d5532b3, 32'h00000000} /* (28, 21, 26) {real, imag} */,
  {32'hbd6fd1df, 32'h00000000} /* (28, 21, 25) {real, imag} */,
  {32'h3effde0a, 32'h00000000} /* (28, 21, 24) {real, imag} */,
  {32'h3e77077e, 32'h00000000} /* (28, 21, 23) {real, imag} */,
  {32'h3d6e8a41, 32'h00000000} /* (28, 21, 22) {real, imag} */,
  {32'h3e7e5091, 32'h00000000} /* (28, 21, 21) {real, imag} */,
  {32'h3debf84f, 32'h00000000} /* (28, 21, 20) {real, imag} */,
  {32'h3de13f67, 32'h00000000} /* (28, 21, 19) {real, imag} */,
  {32'h3e29e15c, 32'h00000000} /* (28, 21, 18) {real, imag} */,
  {32'h3da896e4, 32'h00000000} /* (28, 21, 17) {real, imag} */,
  {32'hbea46843, 32'h00000000} /* (28, 21, 16) {real, imag} */,
  {32'hbec149e0, 32'h00000000} /* (28, 21, 15) {real, imag} */,
  {32'hbea21ee9, 32'h00000000} /* (28, 21, 14) {real, imag} */,
  {32'h3e4a928d, 32'h00000000} /* (28, 21, 13) {real, imag} */,
  {32'hbc1c3c2c, 32'h00000000} /* (28, 21, 12) {real, imag} */,
  {32'hbe5aa734, 32'h00000000} /* (28, 21, 11) {real, imag} */,
  {32'h3ea01ccf, 32'h00000000} /* (28, 21, 10) {real, imag} */,
  {32'h3e6579a2, 32'h00000000} /* (28, 21, 9) {real, imag} */,
  {32'hbe6c568b, 32'h00000000} /* (28, 21, 8) {real, imag} */,
  {32'hbcee7f03, 32'h00000000} /* (28, 21, 7) {real, imag} */,
  {32'h3d136e9a, 32'h00000000} /* (28, 21, 6) {real, imag} */,
  {32'hbe0340d5, 32'h00000000} /* (28, 21, 5) {real, imag} */,
  {32'h3f027e8a, 32'h00000000} /* (28, 21, 4) {real, imag} */,
  {32'h3ed31e42, 32'h00000000} /* (28, 21, 3) {real, imag} */,
  {32'hbd74eb74, 32'h00000000} /* (28, 21, 2) {real, imag} */,
  {32'h3eba7f6f, 32'h00000000} /* (28, 21, 1) {real, imag} */,
  {32'h3e8ef798, 32'h00000000} /* (28, 21, 0) {real, imag} */,
  {32'hbec2ecf8, 32'h00000000} /* (28, 20, 31) {real, imag} */,
  {32'hbf1e74ef, 32'h00000000} /* (28, 20, 30) {real, imag} */,
  {32'hbeace76b, 32'h00000000} /* (28, 20, 29) {real, imag} */,
  {32'hbf489524, 32'h00000000} /* (28, 20, 28) {real, imag} */,
  {32'hbf38636a, 32'h00000000} /* (28, 20, 27) {real, imag} */,
  {32'hbf31dab8, 32'h00000000} /* (28, 20, 26) {real, imag} */,
  {32'hbfa6ad70, 32'h00000000} /* (28, 20, 25) {real, imag} */,
  {32'hbf86c4bf, 32'h00000000} /* (28, 20, 24) {real, imag} */,
  {32'hbf16784f, 32'h00000000} /* (28, 20, 23) {real, imag} */,
  {32'hbf303916, 32'h00000000} /* (28, 20, 22) {real, imag} */,
  {32'h3d33cbb8, 32'h00000000} /* (28, 20, 21) {real, imag} */,
  {32'h3f58d368, 32'h00000000} /* (28, 20, 20) {real, imag} */,
  {32'h3f84777b, 32'h00000000} /* (28, 20, 19) {real, imag} */,
  {32'h3f7934ed, 32'h00000000} /* (28, 20, 18) {real, imag} */,
  {32'h3f152c70, 32'h00000000} /* (28, 20, 17) {real, imag} */,
  {32'h3f2eebd8, 32'h00000000} /* (28, 20, 16) {real, imag} */,
  {32'h3f5a32a2, 32'h00000000} /* (28, 20, 15) {real, imag} */,
  {32'h3f5deecd, 32'h00000000} /* (28, 20, 14) {real, imag} */,
  {32'h3f88744e, 32'h00000000} /* (28, 20, 13) {real, imag} */,
  {32'h3f301939, 32'h00000000} /* (28, 20, 12) {real, imag} */,
  {32'h3f243a6a, 32'h00000000} /* (28, 20, 11) {real, imag} */,
  {32'h3e8cdc30, 32'h00000000} /* (28, 20, 10) {real, imag} */,
  {32'hbe865ef9, 32'h00000000} /* (28, 20, 9) {real, imag} */,
  {32'hbf89441e, 32'h00000000} /* (28, 20, 8) {real, imag} */,
  {32'hbf2e969b, 32'h00000000} /* (28, 20, 7) {real, imag} */,
  {32'hbf2fa1f5, 32'h00000000} /* (28, 20, 6) {real, imag} */,
  {32'hbfaa048a, 32'h00000000} /* (28, 20, 5) {real, imag} */,
  {32'hbf3c1594, 32'h00000000} /* (28, 20, 4) {real, imag} */,
  {32'hbf00b29c, 32'h00000000} /* (28, 20, 3) {real, imag} */,
  {32'hbfb03de9, 32'h00000000} /* (28, 20, 2) {real, imag} */,
  {32'hbf4cfb00, 32'h00000000} /* (28, 20, 1) {real, imag} */,
  {32'hbd384d64, 32'h00000000} /* (28, 20, 0) {real, imag} */,
  {32'hbf3df415, 32'h00000000} /* (28, 19, 31) {real, imag} */,
  {32'hbf700e21, 32'h00000000} /* (28, 19, 30) {real, imag} */,
  {32'hbf1a3b74, 32'h00000000} /* (28, 19, 29) {real, imag} */,
  {32'hbf3cdad9, 32'h00000000} /* (28, 19, 28) {real, imag} */,
  {32'hbf795b58, 32'h00000000} /* (28, 19, 27) {real, imag} */,
  {32'hbf615c86, 32'h00000000} /* (28, 19, 26) {real, imag} */,
  {32'hbf75c56b, 32'h00000000} /* (28, 19, 25) {real, imag} */,
  {32'hbf863c71, 32'h00000000} /* (28, 19, 24) {real, imag} */,
  {32'hbf743a30, 32'h00000000} /* (28, 19, 23) {real, imag} */,
  {32'hbf74b0cb, 32'h00000000} /* (28, 19, 22) {real, imag} */,
  {32'hbe74a944, 32'h00000000} /* (28, 19, 21) {real, imag} */,
  {32'h3f501b73, 32'h00000000} /* (28, 19, 20) {real, imag} */,
  {32'h3f8b064a, 32'h00000000} /* (28, 19, 19) {real, imag} */,
  {32'h3f4e67e5, 32'h00000000} /* (28, 19, 18) {real, imag} */,
  {32'h3f01e5ab, 32'h00000000} /* (28, 19, 17) {real, imag} */,
  {32'h3f66ac85, 32'h00000000} /* (28, 19, 16) {real, imag} */,
  {32'h3f93b42e, 32'h00000000} /* (28, 19, 15) {real, imag} */,
  {32'h3f840b9b, 32'h00000000} /* (28, 19, 14) {real, imag} */,
  {32'h3f80136d, 32'h00000000} /* (28, 19, 13) {real, imag} */,
  {32'h3f0177f5, 32'h00000000} /* (28, 19, 12) {real, imag} */,
  {32'h3f054476, 32'h00000000} /* (28, 19, 11) {real, imag} */,
  {32'h3def98b2, 32'h00000000} /* (28, 19, 10) {real, imag} */,
  {32'hbef4e430, 32'h00000000} /* (28, 19, 9) {real, imag} */,
  {32'hbf5523a7, 32'h00000000} /* (28, 19, 8) {real, imag} */,
  {32'hbf07f596, 32'h00000000} /* (28, 19, 7) {real, imag} */,
  {32'hbf1277dc, 32'h00000000} /* (28, 19, 6) {real, imag} */,
  {32'hbfc2c31c, 32'h00000000} /* (28, 19, 5) {real, imag} */,
  {32'hbf791562, 32'h00000000} /* (28, 19, 4) {real, imag} */,
  {32'hbf0bd921, 32'h00000000} /* (28, 19, 3) {real, imag} */,
  {32'hbfb14ee4, 32'h00000000} /* (28, 19, 2) {real, imag} */,
  {32'hbf92d4b5, 32'h00000000} /* (28, 19, 1) {real, imag} */,
  {32'hbf76e085, 32'h00000000} /* (28, 19, 0) {real, imag} */,
  {32'hbf19f645, 32'h00000000} /* (28, 18, 31) {real, imag} */,
  {32'hbf9335d0, 32'h00000000} /* (28, 18, 30) {real, imag} */,
  {32'hbf869d7f, 32'h00000000} /* (28, 18, 29) {real, imag} */,
  {32'hbf5bc2e9, 32'h00000000} /* (28, 18, 28) {real, imag} */,
  {32'hbf9cf703, 32'h00000000} /* (28, 18, 27) {real, imag} */,
  {32'hbfa447ed, 32'h00000000} /* (28, 18, 26) {real, imag} */,
  {32'hbf7708bb, 32'h00000000} /* (28, 18, 25) {real, imag} */,
  {32'hbf531344, 32'h00000000} /* (28, 18, 24) {real, imag} */,
  {32'hbfb5f91e, 32'h00000000} /* (28, 18, 23) {real, imag} */,
  {32'hbfe1497f, 32'h00000000} /* (28, 18, 22) {real, imag} */,
  {32'hbf9a9e1c, 32'h00000000} /* (28, 18, 21) {real, imag} */,
  {32'h3e69c55c, 32'h00000000} /* (28, 18, 20) {real, imag} */,
  {32'h3f58675b, 32'h00000000} /* (28, 18, 19) {real, imag} */,
  {32'h3f96b71e, 32'h00000000} /* (28, 18, 18) {real, imag} */,
  {32'h3f057664, 32'h00000000} /* (28, 18, 17) {real, imag} */,
  {32'h3f665d6b, 32'h00000000} /* (28, 18, 16) {real, imag} */,
  {32'h3f708fa7, 32'h00000000} /* (28, 18, 15) {real, imag} */,
  {32'h3f93b373, 32'h00000000} /* (28, 18, 14) {real, imag} */,
  {32'h3fa5f135, 32'h00000000} /* (28, 18, 13) {real, imag} */,
  {32'h3f2a82a2, 32'h00000000} /* (28, 18, 12) {real, imag} */,
  {32'h3ef7ce32, 32'h00000000} /* (28, 18, 11) {real, imag} */,
  {32'hbd6dfa77, 32'h00000000} /* (28, 18, 10) {real, imag} */,
  {32'hbf2bf1ff, 32'h00000000} /* (28, 18, 9) {real, imag} */,
  {32'hbf57a67c, 32'h00000000} /* (28, 18, 8) {real, imag} */,
  {32'hbf2fbb7d, 32'h00000000} /* (28, 18, 7) {real, imag} */,
  {32'hbf7364fa, 32'h00000000} /* (28, 18, 6) {real, imag} */,
  {32'hbfaa9b24, 32'h00000000} /* (28, 18, 5) {real, imag} */,
  {32'hbf8c0928, 32'h00000000} /* (28, 18, 4) {real, imag} */,
  {32'hbf55a590, 32'h00000000} /* (28, 18, 3) {real, imag} */,
  {32'hbf846ae5, 32'h00000000} /* (28, 18, 2) {real, imag} */,
  {32'hbf81580f, 32'h00000000} /* (28, 18, 1) {real, imag} */,
  {32'hbf6ff53c, 32'h00000000} /* (28, 18, 0) {real, imag} */,
  {32'hbedfb6bc, 32'h00000000} /* (28, 17, 31) {real, imag} */,
  {32'hbfbc8458, 32'h00000000} /* (28, 17, 30) {real, imag} */,
  {32'hbfccfc38, 32'h00000000} /* (28, 17, 29) {real, imag} */,
  {32'hbfa84666, 32'h00000000} /* (28, 17, 28) {real, imag} */,
  {32'hbfc0a8fc, 32'h00000000} /* (28, 17, 27) {real, imag} */,
  {32'hbfd4d8cd, 32'h00000000} /* (28, 17, 26) {real, imag} */,
  {32'hbfc837a9, 32'h00000000} /* (28, 17, 25) {real, imag} */,
  {32'hbf97083f, 32'h00000000} /* (28, 17, 24) {real, imag} */,
  {32'hbfdcdb74, 32'h00000000} /* (28, 17, 23) {real, imag} */,
  {32'hbf94e731, 32'h00000000} /* (28, 17, 22) {real, imag} */,
  {32'hbf7ea64b, 32'h00000000} /* (28, 17, 21) {real, imag} */,
  {32'h3e43ea23, 32'h00000000} /* (28, 17, 20) {real, imag} */,
  {32'h3f213de2, 32'h00000000} /* (28, 17, 19) {real, imag} */,
  {32'h3f7c85ce, 32'h00000000} /* (28, 17, 18) {real, imag} */,
  {32'h3f58355d, 32'h00000000} /* (28, 17, 17) {real, imag} */,
  {32'h3f254702, 32'h00000000} /* (28, 17, 16) {real, imag} */,
  {32'h3f27cf70, 32'h00000000} /* (28, 17, 15) {real, imag} */,
  {32'h3f97ecea, 32'h00000000} /* (28, 17, 14) {real, imag} */,
  {32'h3f427ca1, 32'h00000000} /* (28, 17, 13) {real, imag} */,
  {32'h3f2723b2, 32'h00000000} /* (28, 17, 12) {real, imag} */,
  {32'h3f0b3c75, 32'h00000000} /* (28, 17, 11) {real, imag} */,
  {32'h3d97630c, 32'h00000000} /* (28, 17, 10) {real, imag} */,
  {32'hbe94746f, 32'h00000000} /* (28, 17, 9) {real, imag} */,
  {32'hbf3e89bb, 32'h00000000} /* (28, 17, 8) {real, imag} */,
  {32'hbf7df908, 32'h00000000} /* (28, 17, 7) {real, imag} */,
  {32'hbf8a26ee, 32'h00000000} /* (28, 17, 6) {real, imag} */,
  {32'hbf2bcfe9, 32'h00000000} /* (28, 17, 5) {real, imag} */,
  {32'hbf85ab08, 32'h00000000} /* (28, 17, 4) {real, imag} */,
  {32'hbf9543a6, 32'h00000000} /* (28, 17, 3) {real, imag} */,
  {32'hbf5bd4a3, 32'h00000000} /* (28, 17, 2) {real, imag} */,
  {32'hbf2a1e0e, 32'h00000000} /* (28, 17, 1) {real, imag} */,
  {32'hbe719e30, 32'h00000000} /* (28, 17, 0) {real, imag} */,
  {32'hbebba993, 32'h00000000} /* (28, 16, 31) {real, imag} */,
  {32'hbfadfaf1, 32'h00000000} /* (28, 16, 30) {real, imag} */,
  {32'hbf8fa882, 32'h00000000} /* (28, 16, 29) {real, imag} */,
  {32'hbf9b570c, 32'h00000000} /* (28, 16, 28) {real, imag} */,
  {32'hbf91aa54, 32'h00000000} /* (28, 16, 27) {real, imag} */,
  {32'hbf92ff02, 32'h00000000} /* (28, 16, 26) {real, imag} */,
  {32'hbfc2dc00, 32'h00000000} /* (28, 16, 25) {real, imag} */,
  {32'hbf9b9a13, 32'h00000000} /* (28, 16, 24) {real, imag} */,
  {32'hbf9d3cb2, 32'h00000000} /* (28, 16, 23) {real, imag} */,
  {32'hbf1b789b, 32'h00000000} /* (28, 16, 22) {real, imag} */,
  {32'hbefdfbac, 32'h00000000} /* (28, 16, 21) {real, imag} */,
  {32'h3f0e1685, 32'h00000000} /* (28, 16, 20) {real, imag} */,
  {32'h3f04953b, 32'h00000000} /* (28, 16, 19) {real, imag} */,
  {32'h3f2c7a98, 32'h00000000} /* (28, 16, 18) {real, imag} */,
  {32'h3f9b3068, 32'h00000000} /* (28, 16, 17) {real, imag} */,
  {32'h3f983b88, 32'h00000000} /* (28, 16, 16) {real, imag} */,
  {32'h3f69a1a4, 32'h00000000} /* (28, 16, 15) {real, imag} */,
  {32'h3f24be62, 32'h00000000} /* (28, 16, 14) {real, imag} */,
  {32'h3f31b9c1, 32'h00000000} /* (28, 16, 13) {real, imag} */,
  {32'h3f3cc5e2, 32'h00000000} /* (28, 16, 12) {real, imag} */,
  {32'h3f56d480, 32'h00000000} /* (28, 16, 11) {real, imag} */,
  {32'h3e5412bf, 32'h00000000} /* (28, 16, 10) {real, imag} */,
  {32'hbec56052, 32'h00000000} /* (28, 16, 9) {real, imag} */,
  {32'hbf94f276, 32'h00000000} /* (28, 16, 8) {real, imag} */,
  {32'hbf9e728a, 32'h00000000} /* (28, 16, 7) {real, imag} */,
  {32'hbf914cb0, 32'h00000000} /* (28, 16, 6) {real, imag} */,
  {32'hbf79f383, 32'h00000000} /* (28, 16, 5) {real, imag} */,
  {32'hbf96179e, 32'h00000000} /* (28, 16, 4) {real, imag} */,
  {32'hbf35a9ef, 32'h00000000} /* (28, 16, 3) {real, imag} */,
  {32'hbf121d5b, 32'h00000000} /* (28, 16, 2) {real, imag} */,
  {32'hbf74c3d0, 32'h00000000} /* (28, 16, 1) {real, imag} */,
  {32'hbecaba24, 32'h00000000} /* (28, 16, 0) {real, imag} */,
  {32'hbefc70d7, 32'h00000000} /* (28, 15, 31) {real, imag} */,
  {32'hbf94255a, 32'h00000000} /* (28, 15, 30) {real, imag} */,
  {32'hbf301b27, 32'h00000000} /* (28, 15, 29) {real, imag} */,
  {32'hbf2415ae, 32'h00000000} /* (28, 15, 28) {real, imag} */,
  {32'hbf1a0761, 32'h00000000} /* (28, 15, 27) {real, imag} */,
  {32'hbf87646e, 32'h00000000} /* (28, 15, 26) {real, imag} */,
  {32'hbfb43644, 32'h00000000} /* (28, 15, 25) {real, imag} */,
  {32'hbf983605, 32'h00000000} /* (28, 15, 24) {real, imag} */,
  {32'hbf8a2cba, 32'h00000000} /* (28, 15, 23) {real, imag} */,
  {32'hbf7637d3, 32'h00000000} /* (28, 15, 22) {real, imag} */,
  {32'hbdb2f01b, 32'h00000000} /* (28, 15, 21) {real, imag} */,
  {32'h3f6b538a, 32'h00000000} /* (28, 15, 20) {real, imag} */,
  {32'h3f3c8317, 32'h00000000} /* (28, 15, 19) {real, imag} */,
  {32'h3f44fe00, 32'h00000000} /* (28, 15, 18) {real, imag} */,
  {32'h3f7ffbb9, 32'h00000000} /* (28, 15, 17) {real, imag} */,
  {32'h3fa86248, 32'h00000000} /* (28, 15, 16) {real, imag} */,
  {32'h3f99fcc8, 32'h00000000} /* (28, 15, 15) {real, imag} */,
  {32'h3f09239b, 32'h00000000} /* (28, 15, 14) {real, imag} */,
  {32'h3f84ee1b, 32'h00000000} /* (28, 15, 13) {real, imag} */,
  {32'h3fa5cbd6, 32'h00000000} /* (28, 15, 12) {real, imag} */,
  {32'h3f88bad3, 32'h00000000} /* (28, 15, 11) {real, imag} */,
  {32'hbe03fb60, 32'h00000000} /* (28, 15, 10) {real, imag} */,
  {32'hbf3acc4e, 32'h00000000} /* (28, 15, 9) {real, imag} */,
  {32'hbfa7ba2a, 32'h00000000} /* (28, 15, 8) {real, imag} */,
  {32'hbfc9a0c6, 32'h00000000} /* (28, 15, 7) {real, imag} */,
  {32'hbfa76baf, 32'h00000000} /* (28, 15, 6) {real, imag} */,
  {32'hbf94051e, 32'h00000000} /* (28, 15, 5) {real, imag} */,
  {32'hbf536420, 32'h00000000} /* (28, 15, 4) {real, imag} */,
  {32'hbf3f3701, 32'h00000000} /* (28, 15, 3) {real, imag} */,
  {32'hbf0f37a9, 32'h00000000} /* (28, 15, 2) {real, imag} */,
  {32'hbf6bf26f, 32'h00000000} /* (28, 15, 1) {real, imag} */,
  {32'hbee1aae5, 32'h00000000} /* (28, 15, 0) {real, imag} */,
  {32'hbecba417, 32'h00000000} /* (28, 14, 31) {real, imag} */,
  {32'hbf41bbdc, 32'h00000000} /* (28, 14, 30) {real, imag} */,
  {32'hbf47a140, 32'h00000000} /* (28, 14, 29) {real, imag} */,
  {32'hbf0513c5, 32'h00000000} /* (28, 14, 28) {real, imag} */,
  {32'hbebb99ae, 32'h00000000} /* (28, 14, 27) {real, imag} */,
  {32'hbf3b376c, 32'h00000000} /* (28, 14, 26) {real, imag} */,
  {32'hbf90399f, 32'h00000000} /* (28, 14, 25) {real, imag} */,
  {32'hbfcd5580, 32'h00000000} /* (28, 14, 24) {real, imag} */,
  {32'hbfab1294, 32'h00000000} /* (28, 14, 23) {real, imag} */,
  {32'hbf7b666e, 32'h00000000} /* (28, 14, 22) {real, imag} */,
  {32'h3c870339, 32'h00000000} /* (28, 14, 21) {real, imag} */,
  {32'h3f567bea, 32'h00000000} /* (28, 14, 20) {real, imag} */,
  {32'h3f70ddb8, 32'h00000000} /* (28, 14, 19) {real, imag} */,
  {32'h3f87da59, 32'h00000000} /* (28, 14, 18) {real, imag} */,
  {32'h3f73ae83, 32'h00000000} /* (28, 14, 17) {real, imag} */,
  {32'h3f9ed04f, 32'h00000000} /* (28, 14, 16) {real, imag} */,
  {32'h3f95a335, 32'h00000000} /* (28, 14, 15) {real, imag} */,
  {32'h3f6b34ad, 32'h00000000} /* (28, 14, 14) {real, imag} */,
  {32'h3fa88976, 32'h00000000} /* (28, 14, 13) {real, imag} */,
  {32'h3fa1758e, 32'h00000000} /* (28, 14, 12) {real, imag} */,
  {32'h3f4dfd54, 32'h00000000} /* (28, 14, 11) {real, imag} */,
  {32'hbc5be9c2, 32'h00000000} /* (28, 14, 10) {real, imag} */,
  {32'hbf6d262c, 32'h00000000} /* (28, 14, 9) {real, imag} */,
  {32'hbf8cd0a5, 32'h00000000} /* (28, 14, 8) {real, imag} */,
  {32'hbf7a1f56, 32'h00000000} /* (28, 14, 7) {real, imag} */,
  {32'hbf03c43e, 32'h00000000} /* (28, 14, 6) {real, imag} */,
  {32'hbee985d6, 32'h00000000} /* (28, 14, 5) {real, imag} */,
  {32'hbed5e0b8, 32'h00000000} /* (28, 14, 4) {real, imag} */,
  {32'hbf81c61e, 32'h00000000} /* (28, 14, 3) {real, imag} */,
  {32'hbf81b3c2, 32'h00000000} /* (28, 14, 2) {real, imag} */,
  {32'hbf83a88d, 32'h00000000} /* (28, 14, 1) {real, imag} */,
  {32'hbeaa7e6e, 32'h00000000} /* (28, 14, 0) {real, imag} */,
  {32'hbf18622a, 32'h00000000} /* (28, 13, 31) {real, imag} */,
  {32'hbf58f1ee, 32'h00000000} /* (28, 13, 30) {real, imag} */,
  {32'hbf7775b9, 32'h00000000} /* (28, 13, 29) {real, imag} */,
  {32'hbf293cc3, 32'h00000000} /* (28, 13, 28) {real, imag} */,
  {32'hbeb2145a, 32'h00000000} /* (28, 13, 27) {real, imag} */,
  {32'hbf175bf5, 32'h00000000} /* (28, 13, 26) {real, imag} */,
  {32'hbf8284db, 32'h00000000} /* (28, 13, 25) {real, imag} */,
  {32'hbf84b160, 32'h00000000} /* (28, 13, 24) {real, imag} */,
  {32'hbeafe550, 32'h00000000} /* (28, 13, 23) {real, imag} */,
  {32'hbe94fa2e, 32'h00000000} /* (28, 13, 22) {real, imag} */,
  {32'h3dc2d76e, 32'h00000000} /* (28, 13, 21) {real, imag} */,
  {32'h3f5db949, 32'h00000000} /* (28, 13, 20) {real, imag} */,
  {32'h3f77d9f7, 32'h00000000} /* (28, 13, 19) {real, imag} */,
  {32'h3fa6acdf, 32'h00000000} /* (28, 13, 18) {real, imag} */,
  {32'h3f83bebb, 32'h00000000} /* (28, 13, 17) {real, imag} */,
  {32'h3f46c2d9, 32'h00000000} /* (28, 13, 16) {real, imag} */,
  {32'h3f818d4d, 32'h00000000} /* (28, 13, 15) {real, imag} */,
  {32'h3f813211, 32'h00000000} /* (28, 13, 14) {real, imag} */,
  {32'h3f805a7b, 32'h00000000} /* (28, 13, 13) {real, imag} */,
  {32'h3f822bef, 32'h00000000} /* (28, 13, 12) {real, imag} */,
  {32'h3f09f66b, 32'h00000000} /* (28, 13, 11) {real, imag} */,
  {32'hbf2daab1, 32'h00000000} /* (28, 13, 10) {real, imag} */,
  {32'hbfc1d6c8, 32'h00000000} /* (28, 13, 9) {real, imag} */,
  {32'hbf8ac7b9, 32'h00000000} /* (28, 13, 8) {real, imag} */,
  {32'hbf10ed1b, 32'h00000000} /* (28, 13, 7) {real, imag} */,
  {32'hbe556b86, 32'h00000000} /* (28, 13, 6) {real, imag} */,
  {32'hbe492826, 32'h00000000} /* (28, 13, 5) {real, imag} */,
  {32'hbeb265b3, 32'h00000000} /* (28, 13, 4) {real, imag} */,
  {32'hbf7da22e, 32'h00000000} /* (28, 13, 3) {real, imag} */,
  {32'hbf9b47c8, 32'h00000000} /* (28, 13, 2) {real, imag} */,
  {32'hbf8856e3, 32'h00000000} /* (28, 13, 1) {real, imag} */,
  {32'hbf02ffc8, 32'h00000000} /* (28, 13, 0) {real, imag} */,
  {32'hbeeef5d3, 32'h00000000} /* (28, 12, 31) {real, imag} */,
  {32'hbf96f727, 32'h00000000} /* (28, 12, 30) {real, imag} */,
  {32'hbf69ca49, 32'h00000000} /* (28, 12, 29) {real, imag} */,
  {32'hbf8513f0, 32'h00000000} /* (28, 12, 28) {real, imag} */,
  {32'hbf981ae5, 32'h00000000} /* (28, 12, 27) {real, imag} */,
  {32'hbface6df, 32'h00000000} /* (28, 12, 26) {real, imag} */,
  {32'hbf8ef817, 32'h00000000} /* (28, 12, 25) {real, imag} */,
  {32'hbf52c16b, 32'h00000000} /* (28, 12, 24) {real, imag} */,
  {32'hbef002c6, 32'h00000000} /* (28, 12, 23) {real, imag} */,
  {32'hbf166de3, 32'h00000000} /* (28, 12, 22) {real, imag} */,
  {32'hbd9784d4, 32'h00000000} /* (28, 12, 21) {real, imag} */,
  {32'h3f70dc91, 32'h00000000} /* (28, 12, 20) {real, imag} */,
  {32'h3fa47572, 32'h00000000} /* (28, 12, 19) {real, imag} */,
  {32'h3fb278fe, 32'h00000000} /* (28, 12, 18) {real, imag} */,
  {32'h3f8a8d2a, 32'h00000000} /* (28, 12, 17) {real, imag} */,
  {32'h3f321fde, 32'h00000000} /* (28, 12, 16) {real, imag} */,
  {32'h3f1208fe, 32'h00000000} /* (28, 12, 15) {real, imag} */,
  {32'h3f6686d1, 32'h00000000} /* (28, 12, 14) {real, imag} */,
  {32'h3f68fc55, 32'h00000000} /* (28, 12, 13) {real, imag} */,
  {32'h3f2a1710, 32'h00000000} /* (28, 12, 12) {real, imag} */,
  {32'h3f29d6af, 32'h00000000} /* (28, 12, 11) {real, imag} */,
  {32'hbeaf0844, 32'h00000000} /* (28, 12, 10) {real, imag} */,
  {32'hbf650a3c, 32'h00000000} /* (28, 12, 9) {real, imag} */,
  {32'hbf614f9d, 32'h00000000} /* (28, 12, 8) {real, imag} */,
  {32'hbf37647b, 32'h00000000} /* (28, 12, 7) {real, imag} */,
  {32'hbf3e4730, 32'h00000000} /* (28, 12, 6) {real, imag} */,
  {32'hbf4cc42b, 32'h00000000} /* (28, 12, 5) {real, imag} */,
  {32'hbf45d3cd, 32'h00000000} /* (28, 12, 4) {real, imag} */,
  {32'hbfa798bf, 32'h00000000} /* (28, 12, 3) {real, imag} */,
  {32'hbfcd479f, 32'h00000000} /* (28, 12, 2) {real, imag} */,
  {32'hbfe2761f, 32'h00000000} /* (28, 12, 1) {real, imag} */,
  {32'hbf3ea405, 32'h00000000} /* (28, 12, 0) {real, imag} */,
  {32'hbec333bd, 32'h00000000} /* (28, 11, 31) {real, imag} */,
  {32'hbf03f511, 32'h00000000} /* (28, 11, 30) {real, imag} */,
  {32'hbec5618e, 32'h00000000} /* (28, 11, 29) {real, imag} */,
  {32'hbf4e314c, 32'h00000000} /* (28, 11, 28) {real, imag} */,
  {32'hbf8e1b7e, 32'h00000000} /* (28, 11, 27) {real, imag} */,
  {32'hbf887e2b, 32'h00000000} /* (28, 11, 26) {real, imag} */,
  {32'hbf397c27, 32'h00000000} /* (28, 11, 25) {real, imag} */,
  {32'hbf2c0394, 32'h00000000} /* (28, 11, 24) {real, imag} */,
  {32'hbf1a1496, 32'h00000000} /* (28, 11, 23) {real, imag} */,
  {32'hbef0b4bc, 32'h00000000} /* (28, 11, 22) {real, imag} */,
  {32'hbe1b1df5, 32'h00000000} /* (28, 11, 21) {real, imag} */,
  {32'h3ddc055a, 32'h00000000} /* (28, 11, 20) {real, imag} */,
  {32'h3f193ef3, 32'h00000000} /* (28, 11, 19) {real, imag} */,
  {32'h3f4c4d95, 32'h00000000} /* (28, 11, 18) {real, imag} */,
  {32'h3f5dedac, 32'h00000000} /* (28, 11, 17) {real, imag} */,
  {32'h3f145e7f, 32'h00000000} /* (28, 11, 16) {real, imag} */,
  {32'h3f061f52, 32'h00000000} /* (28, 11, 15) {real, imag} */,
  {32'h3f49a17b, 32'h00000000} /* (28, 11, 14) {real, imag} */,
  {32'h3f88c202, 32'h00000000} /* (28, 11, 13) {real, imag} */,
  {32'h3eb9e098, 32'h00000000} /* (28, 11, 12) {real, imag} */,
  {32'h3d87265f, 32'h00000000} /* (28, 11, 11) {real, imag} */,
  {32'hbf187b7d, 32'h00000000} /* (28, 11, 10) {real, imag} */,
  {32'hbf033a45, 32'h00000000} /* (28, 11, 9) {real, imag} */,
  {32'hbf0f22ae, 32'h00000000} /* (28, 11, 8) {real, imag} */,
  {32'hbf861cb3, 32'h00000000} /* (28, 11, 7) {real, imag} */,
  {32'hbfa77027, 32'h00000000} /* (28, 11, 6) {real, imag} */,
  {32'hbf7675d0, 32'h00000000} /* (28, 11, 5) {real, imag} */,
  {32'hbeefcb2f, 32'h00000000} /* (28, 11, 4) {real, imag} */,
  {32'hbf5fb4b5, 32'h00000000} /* (28, 11, 3) {real, imag} */,
  {32'hbfa5d2f6, 32'h00000000} /* (28, 11, 2) {real, imag} */,
  {32'hbf87647c, 32'h00000000} /* (28, 11, 1) {real, imag} */,
  {32'hbf0c99fb, 32'h00000000} /* (28, 11, 0) {real, imag} */,
  {32'h3ee56abb, 32'h00000000} /* (28, 10, 31) {real, imag} */,
  {32'h3ecc7c1c, 32'h00000000} /* (28, 10, 30) {real, imag} */,
  {32'h3e93a624, 32'h00000000} /* (28, 10, 29) {real, imag} */,
  {32'h3ea2136d, 32'h00000000} /* (28, 10, 28) {real, imag} */,
  {32'h3eda0fdc, 32'h00000000} /* (28, 10, 27) {real, imag} */,
  {32'h3e1367ed, 32'h00000000} /* (28, 10, 26) {real, imag} */,
  {32'h3f3bf6d9, 32'h00000000} /* (28, 10, 25) {real, imag} */,
  {32'h3f9e2cea, 32'h00000000} /* (28, 10, 24) {real, imag} */,
  {32'h3f726390, 32'h00000000} /* (28, 10, 23) {real, imag} */,
  {32'h3f8f678c, 32'h00000000} /* (28, 10, 22) {real, imag} */,
  {32'h3e82a49b, 32'h00000000} /* (28, 10, 21) {real, imag} */,
  {32'hbf81dba6, 32'h00000000} /* (28, 10, 20) {real, imag} */,
  {32'hbf2c2dca, 32'h00000000} /* (28, 10, 19) {real, imag} */,
  {32'hbefd54b7, 32'h00000000} /* (28, 10, 18) {real, imag} */,
  {32'hbf7c704b, 32'h00000000} /* (28, 10, 17) {real, imag} */,
  {32'hbe90234f, 32'h00000000} /* (28, 10, 16) {real, imag} */,
  {32'hbd1421f3, 32'h00000000} /* (28, 10, 15) {real, imag} */,
  {32'hbe7549a5, 32'h00000000} /* (28, 10, 14) {real, imag} */,
  {32'h3d272679, 32'h00000000} /* (28, 10, 13) {real, imag} */,
  {32'hbf4768d6, 32'h00000000} /* (28, 10, 12) {real, imag} */,
  {32'hbf413be9, 32'h00000000} /* (28, 10, 11) {real, imag} */,
  {32'h3c640224, 32'h00000000} /* (28, 10, 10) {real, imag} */,
  {32'h3ee29236, 32'h00000000} /* (28, 10, 9) {real, imag} */,
  {32'h3ea5ff83, 32'h00000000} /* (28, 10, 8) {real, imag} */,
  {32'h3e1d6290, 32'h00000000} /* (28, 10, 7) {real, imag} */,
  {32'h3e027b31, 32'h00000000} /* (28, 10, 6) {real, imag} */,
  {32'h3eb63f80, 32'h00000000} /* (28, 10, 5) {real, imag} */,
  {32'h3edba31f, 32'h00000000} /* (28, 10, 4) {real, imag} */,
  {32'h3dd578da, 32'h00000000} /* (28, 10, 3) {real, imag} */,
  {32'h3db8be7d, 32'h00000000} /* (28, 10, 2) {real, imag} */,
  {32'h3e93cf66, 32'h00000000} /* (28, 10, 1) {real, imag} */,
  {32'h3ead2b16, 32'h00000000} /* (28, 10, 0) {real, imag} */,
  {32'h3f8dbded, 32'h00000000} /* (28, 9, 31) {real, imag} */,
  {32'h3f99789c, 32'h00000000} /* (28, 9, 30) {real, imag} */,
  {32'h3f9500a3, 32'h00000000} /* (28, 9, 29) {real, imag} */,
  {32'h3f685649, 32'h00000000} /* (28, 9, 28) {real, imag} */,
  {32'h3f5c89f1, 32'h00000000} /* (28, 9, 27) {real, imag} */,
  {32'h3f3451ec, 32'h00000000} /* (28, 9, 26) {real, imag} */,
  {32'h3fa29eab, 32'h00000000} /* (28, 9, 25) {real, imag} */,
  {32'h3fcc3d71, 32'h00000000} /* (28, 9, 24) {real, imag} */,
  {32'h3fa2e392, 32'h00000000} /* (28, 9, 23) {real, imag} */,
  {32'h3fc648f8, 32'h00000000} /* (28, 9, 22) {real, imag} */,
  {32'h3f399c0d, 32'h00000000} /* (28, 9, 21) {real, imag} */,
  {32'hbf56ef73, 32'h00000000} /* (28, 9, 20) {real, imag} */,
  {32'hbf7c8566, 32'h00000000} /* (28, 9, 19) {real, imag} */,
  {32'hbf7d4a39, 32'h00000000} /* (28, 9, 18) {real, imag} */,
  {32'hbfd4ae75, 32'h00000000} /* (28, 9, 17) {real, imag} */,
  {32'hbf8433f9, 32'h00000000} /* (28, 9, 16) {real, imag} */,
  {32'hbf1992fc, 32'h00000000} /* (28, 9, 15) {real, imag} */,
  {32'hbefefdf4, 32'h00000000} /* (28, 9, 14) {real, imag} */,
  {32'hbee9027f, 32'h00000000} /* (28, 9, 13) {real, imag} */,
  {32'hbf6fc3e2, 32'h00000000} /* (28, 9, 12) {real, imag} */,
  {32'hbf31f1ce, 32'h00000000} /* (28, 9, 11) {real, imag} */,
  {32'h3f4d2372, 32'h00000000} /* (28, 9, 10) {real, imag} */,
  {32'h3fb1885b, 32'h00000000} /* (28, 9, 9) {real, imag} */,
  {32'h3f3456be, 32'h00000000} /* (28, 9, 8) {real, imag} */,
  {32'h3f13a470, 32'h00000000} /* (28, 9, 7) {real, imag} */,
  {32'h3ed974c4, 32'h00000000} /* (28, 9, 6) {real, imag} */,
  {32'h3f006db9, 32'h00000000} /* (28, 9, 5) {real, imag} */,
  {32'h3f835602, 32'h00000000} /* (28, 9, 4) {real, imag} */,
  {32'h3f88823b, 32'h00000000} /* (28, 9, 3) {real, imag} */,
  {32'h3f3399c3, 32'h00000000} /* (28, 9, 2) {real, imag} */,
  {32'h3f2bedd2, 32'h00000000} /* (28, 9, 1) {real, imag} */,
  {32'h3f1e8753, 32'h00000000} /* (28, 9, 0) {real, imag} */,
  {32'h3f6664ff, 32'h00000000} /* (28, 8, 31) {real, imag} */,
  {32'h3f7571c1, 32'h00000000} /* (28, 8, 30) {real, imag} */,
  {32'h3f8fb92b, 32'h00000000} /* (28, 8, 29) {real, imag} */,
  {32'h3ed1bed7, 32'h00000000} /* (28, 8, 28) {real, imag} */,
  {32'h3f1ccead, 32'h00000000} /* (28, 8, 27) {real, imag} */,
  {32'h3f8a1e20, 32'h00000000} /* (28, 8, 26) {real, imag} */,
  {32'h3f4c92ba, 32'h00000000} /* (28, 8, 25) {real, imag} */,
  {32'h3f537e3a, 32'h00000000} /* (28, 8, 24) {real, imag} */,
  {32'h3f532694, 32'h00000000} /* (28, 8, 23) {real, imag} */,
  {32'h3fa6e488, 32'h00000000} /* (28, 8, 22) {real, imag} */,
  {32'h3f410cfd, 32'h00000000} /* (28, 8, 21) {real, imag} */,
  {32'hbe872a02, 32'h00000000} /* (28, 8, 20) {real, imag} */,
  {32'hbf4bc613, 32'h00000000} /* (28, 8, 19) {real, imag} */,
  {32'hbfb08293, 32'h00000000} /* (28, 8, 18) {real, imag} */,
  {32'hbfa93065, 32'h00000000} /* (28, 8, 17) {real, imag} */,
  {32'hbf35fcc7, 32'h00000000} /* (28, 8, 16) {real, imag} */,
  {32'hbf1e6103, 32'h00000000} /* (28, 8, 15) {real, imag} */,
  {32'hbf7475df, 32'h00000000} /* (28, 8, 14) {real, imag} */,
  {32'hbf6dcea5, 32'h00000000} /* (28, 8, 13) {real, imag} */,
  {32'hbf43f42c, 32'h00000000} /* (28, 8, 12) {real, imag} */,
  {32'hbf67e3c5, 32'h00000000} /* (28, 8, 11) {real, imag} */,
  {32'h3edeeded, 32'h00000000} /* (28, 8, 10) {real, imag} */,
  {32'h3f7326fb, 32'h00000000} /* (28, 8, 9) {real, imag} */,
  {32'h3f11aae3, 32'h00000000} /* (28, 8, 8) {real, imag} */,
  {32'h3f03b283, 32'h00000000} /* (28, 8, 7) {real, imag} */,
  {32'h3eddbbf0, 32'h00000000} /* (28, 8, 6) {real, imag} */,
  {32'h3ec74cfc, 32'h00000000} /* (28, 8, 5) {real, imag} */,
  {32'h3f242adb, 32'h00000000} /* (28, 8, 4) {real, imag} */,
  {32'h3f6d8992, 32'h00000000} /* (28, 8, 3) {real, imag} */,
  {32'h3f8b47b0, 32'h00000000} /* (28, 8, 2) {real, imag} */,
  {32'h3f98de68, 32'h00000000} /* (28, 8, 1) {real, imag} */,
  {32'h3f33eeee, 32'h00000000} /* (28, 8, 0) {real, imag} */,
  {32'h3f032f03, 32'h00000000} /* (28, 7, 31) {real, imag} */,
  {32'h3f4d0b5b, 32'h00000000} /* (28, 7, 30) {real, imag} */,
  {32'h3f1a8a6a, 32'h00000000} /* (28, 7, 29) {real, imag} */,
  {32'h3e99692d, 32'h00000000} /* (28, 7, 28) {real, imag} */,
  {32'h3f298d4c, 32'h00000000} /* (28, 7, 27) {real, imag} */,
  {32'h3f90c4be, 32'h00000000} /* (28, 7, 26) {real, imag} */,
  {32'h3faa150a, 32'h00000000} /* (28, 7, 25) {real, imag} */,
  {32'h3fad0860, 32'h00000000} /* (28, 7, 24) {real, imag} */,
  {32'h3f517fc4, 32'h00000000} /* (28, 7, 23) {real, imag} */,
  {32'h3f442e35, 32'h00000000} /* (28, 7, 22) {real, imag} */,
  {32'h3f1b3251, 32'h00000000} /* (28, 7, 21) {real, imag} */,
  {32'hbf3888c6, 32'h00000000} /* (28, 7, 20) {real, imag} */,
  {32'hbfb47735, 32'h00000000} /* (28, 7, 19) {real, imag} */,
  {32'hbf829e61, 32'h00000000} /* (28, 7, 18) {real, imag} */,
  {32'hbf90a66a, 32'h00000000} /* (28, 7, 17) {real, imag} */,
  {32'hbf31e145, 32'h00000000} /* (28, 7, 16) {real, imag} */,
  {32'hbf789439, 32'h00000000} /* (28, 7, 15) {real, imag} */,
  {32'hbf758fbc, 32'h00000000} /* (28, 7, 14) {real, imag} */,
  {32'hbf64ff1f, 32'h00000000} /* (28, 7, 13) {real, imag} */,
  {32'hbf16e2de, 32'h00000000} /* (28, 7, 12) {real, imag} */,
  {32'hbf0453f5, 32'h00000000} /* (28, 7, 11) {real, imag} */,
  {32'hbd7e42f5, 32'h00000000} /* (28, 7, 10) {real, imag} */,
  {32'h3ef77cd3, 32'h00000000} /* (28, 7, 9) {real, imag} */,
  {32'h3f4c2673, 32'h00000000} /* (28, 7, 8) {real, imag} */,
  {32'h3f01538c, 32'h00000000} /* (28, 7, 7) {real, imag} */,
  {32'h3e9f9957, 32'h00000000} /* (28, 7, 6) {real, imag} */,
  {32'h3f74f57c, 32'h00000000} /* (28, 7, 5) {real, imag} */,
  {32'h3f9947c6, 32'h00000000} /* (28, 7, 4) {real, imag} */,
  {32'h3f8a61cb, 32'h00000000} /* (28, 7, 3) {real, imag} */,
  {32'h3f9f2d25, 32'h00000000} /* (28, 7, 2) {real, imag} */,
  {32'h3f5bda84, 32'h00000000} /* (28, 7, 1) {real, imag} */,
  {32'h3ea45758, 32'h00000000} /* (28, 7, 0) {real, imag} */,
  {32'h3f0cb859, 32'h00000000} /* (28, 6, 31) {real, imag} */,
  {32'h3f2f88ce, 32'h00000000} /* (28, 6, 30) {real, imag} */,
  {32'h3f48c656, 32'h00000000} /* (28, 6, 29) {real, imag} */,
  {32'h3f257311, 32'h00000000} /* (28, 6, 28) {real, imag} */,
  {32'h3f908001, 32'h00000000} /* (28, 6, 27) {real, imag} */,
  {32'h3fc59ed5, 32'h00000000} /* (28, 6, 26) {real, imag} */,
  {32'h3fbcae18, 32'h00000000} /* (28, 6, 25) {real, imag} */,
  {32'h3f638fe6, 32'h00000000} /* (28, 6, 24) {real, imag} */,
  {32'h3f5fc42c, 32'h00000000} /* (28, 6, 23) {real, imag} */,
  {32'h3f917196, 32'h00000000} /* (28, 6, 22) {real, imag} */,
  {32'h3f6a68e4, 32'h00000000} /* (28, 6, 21) {real, imag} */,
  {32'hbec7d09a, 32'h00000000} /* (28, 6, 20) {real, imag} */,
  {32'hbf87c839, 32'h00000000} /* (28, 6, 19) {real, imag} */,
  {32'hbf6d942a, 32'h00000000} /* (28, 6, 18) {real, imag} */,
  {32'hbf24b9be, 32'h00000000} /* (28, 6, 17) {real, imag} */,
  {32'hbf251a07, 32'h00000000} /* (28, 6, 16) {real, imag} */,
  {32'hbf6ac134, 32'h00000000} /* (28, 6, 15) {real, imag} */,
  {32'hbf87e07e, 32'h00000000} /* (28, 6, 14) {real, imag} */,
  {32'hbf9fc57f, 32'h00000000} /* (28, 6, 13) {real, imag} */,
  {32'hbf6544c4, 32'h00000000} /* (28, 6, 12) {real, imag} */,
  {32'hbf18db68, 32'h00000000} /* (28, 6, 11) {real, imag} */,
  {32'h3e365c84, 32'h00000000} /* (28, 6, 10) {real, imag} */,
  {32'h3f26df8c, 32'h00000000} /* (28, 6, 9) {real, imag} */,
  {32'h3f0aa6ab, 32'h00000000} /* (28, 6, 8) {real, imag} */,
  {32'h3eed1000, 32'h00000000} /* (28, 6, 7) {real, imag} */,
  {32'h3ee41f16, 32'h00000000} /* (28, 6, 6) {real, imag} */,
  {32'h3fa5f783, 32'h00000000} /* (28, 6, 5) {real, imag} */,
  {32'h3ff9ee16, 32'h00000000} /* (28, 6, 4) {real, imag} */,
  {32'h3f95db02, 32'h00000000} /* (28, 6, 3) {real, imag} */,
  {32'h3f24cfee, 32'h00000000} /* (28, 6, 2) {real, imag} */,
  {32'h3f0601a2, 32'h00000000} /* (28, 6, 1) {real, imag} */,
  {32'h3ea291a3, 32'h00000000} /* (28, 6, 0) {real, imag} */,
  {32'h3f09b299, 32'h00000000} /* (28, 5, 31) {real, imag} */,
  {32'h3f64779e, 32'h00000000} /* (28, 5, 30) {real, imag} */,
  {32'h3f8a6227, 32'h00000000} /* (28, 5, 29) {real, imag} */,
  {32'h3f853383, 32'h00000000} /* (28, 5, 28) {real, imag} */,
  {32'h3fa827ae, 32'h00000000} /* (28, 5, 27) {real, imag} */,
  {32'h3fac8fce, 32'h00000000} /* (28, 5, 26) {real, imag} */,
  {32'h3fb10f89, 32'h00000000} /* (28, 5, 25) {real, imag} */,
  {32'h3fac23ee, 32'h00000000} /* (28, 5, 24) {real, imag} */,
  {32'h3f98b195, 32'h00000000} /* (28, 5, 23) {real, imag} */,
  {32'h3f9b1072, 32'h00000000} /* (28, 5, 22) {real, imag} */,
  {32'h3fc7d08e, 32'h00000000} /* (28, 5, 21) {real, imag} */,
  {32'h3f7a1302, 32'h00000000} /* (28, 5, 20) {real, imag} */,
  {32'h3ebb264c, 32'h00000000} /* (28, 5, 19) {real, imag} */,
  {32'h3e6d35d9, 32'h00000000} /* (28, 5, 18) {real, imag} */,
  {32'h3e644234, 32'h00000000} /* (28, 5, 17) {real, imag} */,
  {32'hbd3fa79a, 32'h00000000} /* (28, 5, 16) {real, imag} */,
  {32'hbeb42fc2, 32'h00000000} /* (28, 5, 15) {real, imag} */,
  {32'hbf4ab14d, 32'h00000000} /* (28, 5, 14) {real, imag} */,
  {32'hbf918488, 32'h00000000} /* (28, 5, 13) {real, imag} */,
  {32'hbf40403a, 32'h00000000} /* (28, 5, 12) {real, imag} */,
  {32'hbfa62eb9, 32'h00000000} /* (28, 5, 11) {real, imag} */,
  {32'hbf4bbba2, 32'h00000000} /* (28, 5, 10) {real, imag} */,
  {32'hbe0ec7b9, 32'h00000000} /* (28, 5, 9) {real, imag} */,
  {32'hbe6d4111, 32'h00000000} /* (28, 5, 8) {real, imag} */,
  {32'hbec9c9cd, 32'h00000000} /* (28, 5, 7) {real, imag} */,
  {32'hbe1d9671, 32'h00000000} /* (28, 5, 6) {real, imag} */,
  {32'h3f83c2de, 32'h00000000} /* (28, 5, 5) {real, imag} */,
  {32'h3fa9775c, 32'h00000000} /* (28, 5, 4) {real, imag} */,
  {32'h3f88cd40, 32'h00000000} /* (28, 5, 3) {real, imag} */,
  {32'h3f4360c7, 32'h00000000} /* (28, 5, 2) {real, imag} */,
  {32'h3f1d6778, 32'h00000000} /* (28, 5, 1) {real, imag} */,
  {32'h3f04dc50, 32'h00000000} /* (28, 5, 0) {real, imag} */,
  {32'h3eeb121d, 32'h00000000} /* (28, 4, 31) {real, imag} */,
  {32'h3f59ff89, 32'h00000000} /* (28, 4, 30) {real, imag} */,
  {32'h3f882f31, 32'h00000000} /* (28, 4, 29) {real, imag} */,
  {32'h3f950eef, 32'h00000000} /* (28, 4, 28) {real, imag} */,
  {32'h3f433eb5, 32'h00000000} /* (28, 4, 27) {real, imag} */,
  {32'h3cbac340, 32'h00000000} /* (28, 4, 26) {real, imag} */,
  {32'hbdbcd8cb, 32'h00000000} /* (28, 4, 25) {real, imag} */,
  {32'h3f3edb9a, 32'h00000000} /* (28, 4, 24) {real, imag} */,
  {32'h3f698baf, 32'h00000000} /* (28, 4, 23) {real, imag} */,
  {32'h3f20eb88, 32'h00000000} /* (28, 4, 22) {real, imag} */,
  {32'h3f7458f1, 32'h00000000} /* (28, 4, 21) {real, imag} */,
  {32'h3f665c15, 32'h00000000} /* (28, 4, 20) {real, imag} */,
  {32'h3f4366c3, 32'h00000000} /* (28, 4, 19) {real, imag} */,
  {32'h3f9b4cde, 32'h00000000} /* (28, 4, 18) {real, imag} */,
  {32'h3fa30404, 32'h00000000} /* (28, 4, 17) {real, imag} */,
  {32'h3f2ff068, 32'h00000000} /* (28, 4, 16) {real, imag} */,
  {32'hbefac3bb, 32'h00000000} /* (28, 4, 15) {real, imag} */,
  {32'hbf2f14da, 32'h00000000} /* (28, 4, 14) {real, imag} */,
  {32'hbf5b8c46, 32'h00000000} /* (28, 4, 13) {real, imag} */,
  {32'hbed71cd2, 32'h00000000} /* (28, 4, 12) {real, imag} */,
  {32'hbf5f6cba, 32'h00000000} /* (28, 4, 11) {real, imag} */,
  {32'hbf85d8d8, 32'h00000000} /* (28, 4, 10) {real, imag} */,
  {32'hbf03b0fb, 32'h00000000} /* (28, 4, 9) {real, imag} */,
  {32'hbf43f7f8, 32'h00000000} /* (28, 4, 8) {real, imag} */,
  {32'hbf578623, 32'h00000000} /* (28, 4, 7) {real, imag} */,
  {32'hbf465eb7, 32'h00000000} /* (28, 4, 6) {real, imag} */,
  {32'h3f0b5401, 32'h00000000} /* (28, 4, 5) {real, imag} */,
  {32'h3f6d5365, 32'h00000000} /* (28, 4, 4) {real, imag} */,
  {32'h3f833a7c, 32'h00000000} /* (28, 4, 3) {real, imag} */,
  {32'h3f9c08b3, 32'h00000000} /* (28, 4, 2) {real, imag} */,
  {32'h3ede31ef, 32'h00000000} /* (28, 4, 1) {real, imag} */,
  {32'h3e7f8bc4, 32'h00000000} /* (28, 4, 0) {real, imag} */,
  {32'h3ec572be, 32'h00000000} /* (28, 3, 31) {real, imag} */,
  {32'h3f80722a, 32'h00000000} /* (28, 3, 30) {real, imag} */,
  {32'h3fa43c23, 32'h00000000} /* (28, 3, 29) {real, imag} */,
  {32'h3fdbeb03, 32'h00000000} /* (28, 3, 28) {real, imag} */,
  {32'h3fba8722, 32'h00000000} /* (28, 3, 27) {real, imag} */,
  {32'h3f121b73, 32'h00000000} /* (28, 3, 26) {real, imag} */,
  {32'h3d7aac15, 32'h00000000} /* (28, 3, 25) {real, imag} */,
  {32'h3ea06809, 32'h00000000} /* (28, 3, 24) {real, imag} */,
  {32'h3efc2b24, 32'h00000000} /* (28, 3, 23) {real, imag} */,
  {32'h3ed5700b, 32'h00000000} /* (28, 3, 22) {real, imag} */,
  {32'h3f098cc4, 32'h00000000} /* (28, 3, 21) {real, imag} */,
  {32'h3f71158c, 32'h00000000} /* (28, 3, 20) {real, imag} */,
  {32'h3f4045a0, 32'h00000000} /* (28, 3, 19) {real, imag} */,
  {32'h3f7e1598, 32'h00000000} /* (28, 3, 18) {real, imag} */,
  {32'h3fa52912, 32'h00000000} /* (28, 3, 17) {real, imag} */,
  {32'h3f7e79c8, 32'h00000000} /* (28, 3, 16) {real, imag} */,
  {32'hbee6c919, 32'h00000000} /* (28, 3, 15) {real, imag} */,
  {32'hbf3376f8, 32'h00000000} /* (28, 3, 14) {real, imag} */,
  {32'hbf73fa39, 32'h00000000} /* (28, 3, 13) {real, imag} */,
  {32'hbf2b526e, 32'h00000000} /* (28, 3, 12) {real, imag} */,
  {32'hbecccd52, 32'h00000000} /* (28, 3, 11) {real, imag} */,
  {32'hbf50c125, 32'h00000000} /* (28, 3, 10) {real, imag} */,
  {32'hbf555b7d, 32'h00000000} /* (28, 3, 9) {real, imag} */,
  {32'hbf145d53, 32'h00000000} /* (28, 3, 8) {real, imag} */,
  {32'hbee30761, 32'h00000000} /* (28, 3, 7) {real, imag} */,
  {32'hbf8c9a64, 32'h00000000} /* (28, 3, 6) {real, imag} */,
  {32'hbeddc4b9, 32'h00000000} /* (28, 3, 5) {real, imag} */,
  {32'h3eafe956, 32'h00000000} /* (28, 3, 4) {real, imag} */,
  {32'h3f8812a1, 32'h00000000} /* (28, 3, 3) {real, imag} */,
  {32'h3fc731f8, 32'h00000000} /* (28, 3, 2) {real, imag} */,
  {32'h3f69630c, 32'h00000000} /* (28, 3, 1) {real, imag} */,
  {32'h3edd1a39, 32'h00000000} /* (28, 3, 0) {real, imag} */,
  {32'h3f068e7c, 32'h00000000} /* (28, 2, 31) {real, imag} */,
  {32'h3f932671, 32'h00000000} /* (28, 2, 30) {real, imag} */,
  {32'h3f74ef51, 32'h00000000} /* (28, 2, 29) {real, imag} */,
  {32'h3f7d6599, 32'h00000000} /* (28, 2, 28) {real, imag} */,
  {32'h3f97cdd8, 32'h00000000} /* (28, 2, 27) {real, imag} */,
  {32'h3f49136b, 32'h00000000} /* (28, 2, 26) {real, imag} */,
  {32'h3f37abf5, 32'h00000000} /* (28, 2, 25) {real, imag} */,
  {32'h3fa41c24, 32'h00000000} /* (28, 2, 24) {real, imag} */,
  {32'h3f9409d9, 32'h00000000} /* (28, 2, 23) {real, imag} */,
  {32'h3f82a727, 32'h00000000} /* (28, 2, 22) {real, imag} */,
  {32'h3f7d9fe4, 32'h00000000} /* (28, 2, 21) {real, imag} */,
  {32'h3fa0fe96, 32'h00000000} /* (28, 2, 20) {real, imag} */,
  {32'h3f59cfff, 32'h00000000} /* (28, 2, 19) {real, imag} */,
  {32'h3eb2b996, 32'h00000000} /* (28, 2, 18) {real, imag} */,
  {32'h3f41da8a, 32'h00000000} /* (28, 2, 17) {real, imag} */,
  {32'h3f303ff4, 32'h00000000} /* (28, 2, 16) {real, imag} */,
  {32'hbf689290, 32'h00000000} /* (28, 2, 15) {real, imag} */,
  {32'hbf7a9681, 32'h00000000} /* (28, 2, 14) {real, imag} */,
  {32'hbf794703, 32'h00000000} /* (28, 2, 13) {real, imag} */,
  {32'hbf10f9ba, 32'h00000000} /* (28, 2, 12) {real, imag} */,
  {32'hbec0b335, 32'h00000000} /* (28, 2, 11) {real, imag} */,
  {32'hbfd0d4f6, 32'h00000000} /* (28, 2, 10) {real, imag} */,
  {32'hc0061a52, 32'h00000000} /* (28, 2, 9) {real, imag} */,
  {32'hbf64d623, 32'h00000000} /* (28, 2, 8) {real, imag} */,
  {32'hbf014bb9, 32'h00000000} /* (28, 2, 7) {real, imag} */,
  {32'hbf7a9051, 32'h00000000} /* (28, 2, 6) {real, imag} */,
  {32'hbf037865, 32'h00000000} /* (28, 2, 5) {real, imag} */,
  {32'h3eae9db7, 32'h00000000} /* (28, 2, 4) {real, imag} */,
  {32'h3f7afcc9, 32'h00000000} /* (28, 2, 3) {real, imag} */,
  {32'h3f7ba50e, 32'h00000000} /* (28, 2, 2) {real, imag} */,
  {32'h3f679064, 32'h00000000} /* (28, 2, 1) {real, imag} */,
  {32'h3f17e2e0, 32'h00000000} /* (28, 2, 0) {real, imag} */,
  {32'h3f08d4de, 32'h00000000} /* (28, 1, 31) {real, imag} */,
  {32'h3f410fed, 32'h00000000} /* (28, 1, 30) {real, imag} */,
  {32'h3f40c615, 32'h00000000} /* (28, 1, 29) {real, imag} */,
  {32'h3eff542d, 32'h00000000} /* (28, 1, 28) {real, imag} */,
  {32'h3f26bc04, 32'h00000000} /* (28, 1, 27) {real, imag} */,
  {32'h3ea7e9ad, 32'h00000000} /* (28, 1, 26) {real, imag} */,
  {32'h3f137962, 32'h00000000} /* (28, 1, 25) {real, imag} */,
  {32'h3fa6976f, 32'h00000000} /* (28, 1, 24) {real, imag} */,
  {32'h3fda4dc3, 32'h00000000} /* (28, 1, 23) {real, imag} */,
  {32'h3fca3a90, 32'h00000000} /* (28, 1, 22) {real, imag} */,
  {32'h3fa9d1ec, 32'h00000000} /* (28, 1, 21) {real, imag} */,
  {32'h3f4fc69d, 32'h00000000} /* (28, 1, 20) {real, imag} */,
  {32'h3f87c70b, 32'h00000000} /* (28, 1, 19) {real, imag} */,
  {32'h3fa4bd17, 32'h00000000} /* (28, 1, 18) {real, imag} */,
  {32'h3fb743c0, 32'h00000000} /* (28, 1, 17) {real, imag} */,
  {32'h3f89b00a, 32'h00000000} /* (28, 1, 16) {real, imag} */,
  {32'hbf03ba98, 32'h00000000} /* (28, 1, 15) {real, imag} */,
  {32'hbf4a3747, 32'h00000000} /* (28, 1, 14) {real, imag} */,
  {32'hbf936af6, 32'h00000000} /* (28, 1, 13) {real, imag} */,
  {32'hbf98d229, 32'h00000000} /* (28, 1, 12) {real, imag} */,
  {32'hbf4690db, 32'h00000000} /* (28, 1, 11) {real, imag} */,
  {32'hbfbca6b7, 32'h00000000} /* (28, 1, 10) {real, imag} */,
  {32'hbfee817c, 32'h00000000} /* (28, 1, 9) {real, imag} */,
  {32'hbf548862, 32'h00000000} /* (28, 1, 8) {real, imag} */,
  {32'hbf26f751, 32'h00000000} /* (28, 1, 7) {real, imag} */,
  {32'hbf237ac5, 32'h00000000} /* (28, 1, 6) {real, imag} */,
  {32'hbe168531, 32'h00000000} /* (28, 1, 5) {real, imag} */,
  {32'h3f067de8, 32'h00000000} /* (28, 1, 4) {real, imag} */,
  {32'h3f5d9fcf, 32'h00000000} /* (28, 1, 3) {real, imag} */,
  {32'h3f5aca79, 32'h00000000} /* (28, 1, 2) {real, imag} */,
  {32'h3f2cdd7a, 32'h00000000} /* (28, 1, 1) {real, imag} */,
  {32'h3ee2e1c5, 32'h00000000} /* (28, 1, 0) {real, imag} */,
  {32'h3dda59d0, 32'h00000000} /* (28, 0, 31) {real, imag} */,
  {32'h3e88fb6d, 32'h00000000} /* (28, 0, 30) {real, imag} */,
  {32'h3ed5d380, 32'h00000000} /* (28, 0, 29) {real, imag} */,
  {32'h3e57b212, 32'h00000000} /* (28, 0, 28) {real, imag} */,
  {32'h3e165640, 32'h00000000} /* (28, 0, 27) {real, imag} */,
  {32'h3d45bed2, 32'h00000000} /* (28, 0, 26) {real, imag} */,
  {32'h3eaaa152, 32'h00000000} /* (28, 0, 25) {real, imag} */,
  {32'h3f0ea6c1, 32'h00000000} /* (28, 0, 24) {real, imag} */,
  {32'h3f3e56ec, 32'h00000000} /* (28, 0, 23) {real, imag} */,
  {32'h3f3c9e25, 32'h00000000} /* (28, 0, 22) {real, imag} */,
  {32'h3f40f55a, 32'h00000000} /* (28, 0, 21) {real, imag} */,
  {32'h3f0ae261, 32'h00000000} /* (28, 0, 20) {real, imag} */,
  {32'h3f480f97, 32'h00000000} /* (28, 0, 19) {real, imag} */,
  {32'h3f4da27b, 32'h00000000} /* (28, 0, 18) {real, imag} */,
  {32'h3f28524c, 32'h00000000} /* (28, 0, 17) {real, imag} */,
  {32'h3eda3081, 32'h00000000} /* (28, 0, 16) {real, imag} */,
  {32'hbece6bba, 32'h00000000} /* (28, 0, 15) {real, imag} */,
  {32'hbea01ed6, 32'h00000000} /* (28, 0, 14) {real, imag} */,
  {32'hbf230831, 32'h00000000} /* (28, 0, 13) {real, imag} */,
  {32'hbf8e2b03, 32'h00000000} /* (28, 0, 12) {real, imag} */,
  {32'hbf2149c4, 32'h00000000} /* (28, 0, 11) {real, imag} */,
  {32'hbe0493ff, 32'h00000000} /* (28, 0, 10) {real, imag} */,
  {32'hbe355a0a, 32'h00000000} /* (28, 0, 9) {real, imag} */,
  {32'hbe1d4250, 32'h00000000} /* (28, 0, 8) {real, imag} */,
  {32'hbee02a79, 32'h00000000} /* (28, 0, 7) {real, imag} */,
  {32'hbef30e41, 32'h00000000} /* (28, 0, 6) {real, imag} */,
  {32'h3d876da6, 32'h00000000} /* (28, 0, 5) {real, imag} */,
  {32'h3ed0ba36, 32'h00000000} /* (28, 0, 4) {real, imag} */,
  {32'h3ec757c5, 32'h00000000} /* (28, 0, 3) {real, imag} */,
  {32'h3f00a56e, 32'h00000000} /* (28, 0, 2) {real, imag} */,
  {32'h3e89cdbe, 32'h00000000} /* (28, 0, 1) {real, imag} */,
  {32'h3db87bd2, 32'h00000000} /* (28, 0, 0) {real, imag} */,
  {32'h3d7df105, 32'h00000000} /* (27, 31, 31) {real, imag} */,
  {32'hbd80fb1e, 32'h00000000} /* (27, 31, 30) {real, imag} */,
  {32'h3db314b7, 32'h00000000} /* (27, 31, 29) {real, imag} */,
  {32'h3f2a1637, 32'h00000000} /* (27, 31, 28) {real, imag} */,
  {32'h3f541fd8, 32'h00000000} /* (27, 31, 27) {real, imag} */,
  {32'h3f3404f5, 32'h00000000} /* (27, 31, 26) {real, imag} */,
  {32'h3f84b5a0, 32'h00000000} /* (27, 31, 25) {real, imag} */,
  {32'h3ef6e4be, 32'h00000000} /* (27, 31, 24) {real, imag} */,
  {32'h3ed78598, 32'h00000000} /* (27, 31, 23) {real, imag} */,
  {32'h3e99ca0e, 32'h00000000} /* (27, 31, 22) {real, imag} */,
  {32'hbcd3e2a8, 32'h00000000} /* (27, 31, 21) {real, imag} */,
  {32'hbed82eee, 32'h00000000} /* (27, 31, 20) {real, imag} */,
  {32'hbe83be0c, 32'h00000000} /* (27, 31, 19) {real, imag} */,
  {32'hbc0aa3c8, 32'h00000000} /* (27, 31, 18) {real, imag} */,
  {32'hbd8f4466, 32'h00000000} /* (27, 31, 17) {real, imag} */,
  {32'hbe09b1ad, 32'h00000000} /* (27, 31, 16) {real, imag} */,
  {32'hbe384390, 32'h00000000} /* (27, 31, 15) {real, imag} */,
  {32'hbf4ea421, 32'h00000000} /* (27, 31, 14) {real, imag} */,
  {32'hbf9dbf49, 32'h00000000} /* (27, 31, 13) {real, imag} */,
  {32'hbf499947, 32'h00000000} /* (27, 31, 12) {real, imag} */,
  {32'hbee8c01c, 32'h00000000} /* (27, 31, 11) {real, imag} */,
  {32'h3e25f2ab, 32'h00000000} /* (27, 31, 10) {real, imag} */,
  {32'h3f113b19, 32'h00000000} /* (27, 31, 9) {real, imag} */,
  {32'h3ee837b8, 32'h00000000} /* (27, 31, 8) {real, imag} */,
  {32'h3e6a6db9, 32'h00000000} /* (27, 31, 7) {real, imag} */,
  {32'h3eb8fac4, 32'h00000000} /* (27, 31, 6) {real, imag} */,
  {32'h3f3469d2, 32'h00000000} /* (27, 31, 5) {real, imag} */,
  {32'h3f398a58, 32'h00000000} /* (27, 31, 4) {real, imag} */,
  {32'h3ede4d7b, 32'h00000000} /* (27, 31, 3) {real, imag} */,
  {32'h3f899bde, 32'h00000000} /* (27, 31, 2) {real, imag} */,
  {32'h3f4fdfba, 32'h00000000} /* (27, 31, 1) {real, imag} */,
  {32'h3e611b31, 32'h00000000} /* (27, 31, 0) {real, imag} */,
  {32'h3ebc4d28, 32'h00000000} /* (27, 30, 31) {real, imag} */,
  {32'h3e4f0f5e, 32'h00000000} /* (27, 30, 30) {real, imag} */,
  {32'h3eba9acc, 32'h00000000} /* (27, 30, 29) {real, imag} */,
  {32'h3fae6efb, 32'h00000000} /* (27, 30, 28) {real, imag} */,
  {32'h3fc0673f, 32'h00000000} /* (27, 30, 27) {real, imag} */,
  {32'h3f7fdbf5, 32'h00000000} /* (27, 30, 26) {real, imag} */,
  {32'h3fc0b359, 32'h00000000} /* (27, 30, 25) {real, imag} */,
  {32'h3f6b8132, 32'h00000000} /* (27, 30, 24) {real, imag} */,
  {32'h3faad91e, 32'h00000000} /* (27, 30, 23) {real, imag} */,
  {32'h3f56b39c, 32'h00000000} /* (27, 30, 22) {real, imag} */,
  {32'h3e0efe0e, 32'h00000000} /* (27, 30, 21) {real, imag} */,
  {32'hbf162373, 32'h00000000} /* (27, 30, 20) {real, imag} */,
  {32'hbf62381e, 32'h00000000} /* (27, 30, 19) {real, imag} */,
  {32'hbf1bc4b9, 32'h00000000} /* (27, 30, 18) {real, imag} */,
  {32'hbeed9c13, 32'h00000000} /* (27, 30, 17) {real, imag} */,
  {32'hbf3d2c0e, 32'h00000000} /* (27, 30, 16) {real, imag} */,
  {32'hbf40ef74, 32'h00000000} /* (27, 30, 15) {real, imag} */,
  {32'hbfce7aba, 32'h00000000} /* (27, 30, 14) {real, imag} */,
  {32'hbfd35023, 32'h00000000} /* (27, 30, 13) {real, imag} */,
  {32'hbfab7b12, 32'h00000000} /* (27, 30, 12) {real, imag} */,
  {32'hbf4bafe2, 32'h00000000} /* (27, 30, 11) {real, imag} */,
  {32'h3ecc59bf, 32'h00000000} /* (27, 30, 10) {real, imag} */,
  {32'h3f8810f9, 32'h00000000} /* (27, 30, 9) {real, imag} */,
  {32'h3f3828ea, 32'h00000000} /* (27, 30, 8) {real, imag} */,
  {32'h3f496d35, 32'h00000000} /* (27, 30, 7) {real, imag} */,
  {32'h3f1215e8, 32'h00000000} /* (27, 30, 6) {real, imag} */,
  {32'h3f7a186c, 32'h00000000} /* (27, 30, 5) {real, imag} */,
  {32'h3fb13374, 32'h00000000} /* (27, 30, 4) {real, imag} */,
  {32'h3f99e0d9, 32'h00000000} /* (27, 30, 3) {real, imag} */,
  {32'h3f92e685, 32'h00000000} /* (27, 30, 2) {real, imag} */,
  {32'h3f0da454, 32'h00000000} /* (27, 30, 1) {real, imag} */,
  {32'h3e4da374, 32'h00000000} /* (27, 30, 0) {real, imag} */,
  {32'h3f250518, 32'h00000000} /* (27, 29, 31) {real, imag} */,
  {32'h3f6c7e48, 32'h00000000} /* (27, 29, 30) {real, imag} */,
  {32'h3f6703c9, 32'h00000000} /* (27, 29, 29) {real, imag} */,
  {32'h3fbba98e, 32'h00000000} /* (27, 29, 28) {real, imag} */,
  {32'h3fb0b6d0, 32'h00000000} /* (27, 29, 27) {real, imag} */,
  {32'h3f288819, 32'h00000000} /* (27, 29, 26) {real, imag} */,
  {32'h3f950d7e, 32'h00000000} /* (27, 29, 25) {real, imag} */,
  {32'h3f9a2dd6, 32'h00000000} /* (27, 29, 24) {real, imag} */,
  {32'h3f8aaf35, 32'h00000000} /* (27, 29, 23) {real, imag} */,
  {32'h3f12ef24, 32'h00000000} /* (27, 29, 22) {real, imag} */,
  {32'h3eb95555, 32'h00000000} /* (27, 29, 21) {real, imag} */,
  {32'hbf2f998e, 32'h00000000} /* (27, 29, 20) {real, imag} */,
  {32'hbfa566ef, 32'h00000000} /* (27, 29, 19) {real, imag} */,
  {32'hbf9f0e58, 32'h00000000} /* (27, 29, 18) {real, imag} */,
  {32'hbf426657, 32'h00000000} /* (27, 29, 17) {real, imag} */,
  {32'hbf81334c, 32'h00000000} /* (27, 29, 16) {real, imag} */,
  {32'hbf68e4bd, 32'h00000000} /* (27, 29, 15) {real, imag} */,
  {32'hbf9a9a08, 32'h00000000} /* (27, 29, 14) {real, imag} */,
  {32'hbf5edf98, 32'h00000000} /* (27, 29, 13) {real, imag} */,
  {32'hbf7fe279, 32'h00000000} /* (27, 29, 12) {real, imag} */,
  {32'hbf3a7e17, 32'h00000000} /* (27, 29, 11) {real, imag} */,
  {32'h3ef0d5fe, 32'h00000000} /* (27, 29, 10) {real, imag} */,
  {32'h3fa5fe6e, 32'h00000000} /* (27, 29, 9) {real, imag} */,
  {32'h3f83a044, 32'h00000000} /* (27, 29, 8) {real, imag} */,
  {32'h3f4a2851, 32'h00000000} /* (27, 29, 7) {real, imag} */,
  {32'h3f1e268c, 32'h00000000} /* (27, 29, 6) {real, imag} */,
  {32'h3f94690a, 32'h00000000} /* (27, 29, 5) {real, imag} */,
  {32'h3fd451ef, 32'h00000000} /* (27, 29, 4) {real, imag} */,
  {32'h3fcf5109, 32'h00000000} /* (27, 29, 3) {real, imag} */,
  {32'h3f718a54, 32'h00000000} /* (27, 29, 2) {real, imag} */,
  {32'h3e814ec8, 32'h00000000} /* (27, 29, 1) {real, imag} */,
  {32'h3e70ff74, 32'h00000000} /* (27, 29, 0) {real, imag} */,
  {32'h3f299319, 32'h00000000} /* (27, 28, 31) {real, imag} */,
  {32'h3fa197da, 32'h00000000} /* (27, 28, 30) {real, imag} */,
  {32'h3f5e74aa, 32'h00000000} /* (27, 28, 29) {real, imag} */,
  {32'h3f82cba5, 32'h00000000} /* (27, 28, 28) {real, imag} */,
  {32'h3fa0f286, 32'h00000000} /* (27, 28, 27) {real, imag} */,
  {32'h3f6cde77, 32'h00000000} /* (27, 28, 26) {real, imag} */,
  {32'h3f086869, 32'h00000000} /* (27, 28, 25) {real, imag} */,
  {32'h3f90897b, 32'h00000000} /* (27, 28, 24) {real, imag} */,
  {32'h3f6aa2cb, 32'h00000000} /* (27, 28, 23) {real, imag} */,
  {32'h3ed62a3a, 32'h00000000} /* (27, 28, 22) {real, imag} */,
  {32'h3f487051, 32'h00000000} /* (27, 28, 21) {real, imag} */,
  {32'hbf61e9e6, 32'h00000000} /* (27, 28, 20) {real, imag} */,
  {32'hbfd7b7d4, 32'h00000000} /* (27, 28, 19) {real, imag} */,
  {32'hbf96ce38, 32'h00000000} /* (27, 28, 18) {real, imag} */,
  {32'hbf4c33c7, 32'h00000000} /* (27, 28, 17) {real, imag} */,
  {32'hbf837725, 32'h00000000} /* (27, 28, 16) {real, imag} */,
  {32'hbf7b3cf5, 32'h00000000} /* (27, 28, 15) {real, imag} */,
  {32'hbf450873, 32'h00000000} /* (27, 28, 14) {real, imag} */,
  {32'hbf49f70a, 32'h00000000} /* (27, 28, 13) {real, imag} */,
  {32'hbf499cd3, 32'h00000000} /* (27, 28, 12) {real, imag} */,
  {32'hbee7e8a8, 32'h00000000} /* (27, 28, 11) {real, imag} */,
  {32'h3f5f280e, 32'h00000000} /* (27, 28, 10) {real, imag} */,
  {32'h3ff2242c, 32'h00000000} /* (27, 28, 9) {real, imag} */,
  {32'h3f9a4991, 32'h00000000} /* (27, 28, 8) {real, imag} */,
  {32'h3f267bec, 32'h00000000} /* (27, 28, 7) {real, imag} */,
  {32'h3f6a58f4, 32'h00000000} /* (27, 28, 6) {real, imag} */,
  {32'h3fc4a1aa, 32'h00000000} /* (27, 28, 5) {real, imag} */,
  {32'h3f8097fb, 32'h00000000} /* (27, 28, 4) {real, imag} */,
  {32'h3f632e8d, 32'h00000000} /* (27, 28, 3) {real, imag} */,
  {32'h3f9c9c29, 32'h00000000} /* (27, 28, 2) {real, imag} */,
  {32'h3f3a79ec, 32'h00000000} /* (27, 28, 1) {real, imag} */,
  {32'h3f1da7dc, 32'h00000000} /* (27, 28, 0) {real, imag} */,
  {32'h3ede11c4, 32'h00000000} /* (27, 27, 31) {real, imag} */,
  {32'h3f5f6559, 32'h00000000} /* (27, 27, 30) {real, imag} */,
  {32'h3f7840ae, 32'h00000000} /* (27, 27, 29) {real, imag} */,
  {32'h3fb163c6, 32'h00000000} /* (27, 27, 28) {real, imag} */,
  {32'h3fb766b0, 32'h00000000} /* (27, 27, 27) {real, imag} */,
  {32'h3f8d1ed8, 32'h00000000} /* (27, 27, 26) {real, imag} */,
  {32'h3eff30d8, 32'h00000000} /* (27, 27, 25) {real, imag} */,
  {32'h3f13af39, 32'h00000000} /* (27, 27, 24) {real, imag} */,
  {32'h3f2dc011, 32'h00000000} /* (27, 27, 23) {real, imag} */,
  {32'h3f5a901b, 32'h00000000} /* (27, 27, 22) {real, imag} */,
  {32'h3f8d9ab5, 32'h00000000} /* (27, 27, 21) {real, imag} */,
  {32'hbeb9e86f, 32'h00000000} /* (27, 27, 20) {real, imag} */,
  {32'hbf7bc6ae, 32'h00000000} /* (27, 27, 19) {real, imag} */,
  {32'hbfba62ee, 32'h00000000} /* (27, 27, 18) {real, imag} */,
  {32'hbfb8925c, 32'h00000000} /* (27, 27, 17) {real, imag} */,
  {32'hbf8e5a0f, 32'h00000000} /* (27, 27, 16) {real, imag} */,
  {32'hbf6fa410, 32'h00000000} /* (27, 27, 15) {real, imag} */,
  {32'hbeabfda3, 32'h00000000} /* (27, 27, 14) {real, imag} */,
  {32'hbec227ba, 32'h00000000} /* (27, 27, 13) {real, imag} */,
  {32'hbf544fbd, 32'h00000000} /* (27, 27, 12) {real, imag} */,
  {32'hbf31984f, 32'h00000000} /* (27, 27, 11) {real, imag} */,
  {32'h3f10a85e, 32'h00000000} /* (27, 27, 10) {real, imag} */,
  {32'h3facee77, 32'h00000000} /* (27, 27, 9) {real, imag} */,
  {32'h3f859a28, 32'h00000000} /* (27, 27, 8) {real, imag} */,
  {32'h3f54ead6, 32'h00000000} /* (27, 27, 7) {real, imag} */,
  {32'h3f6c595c, 32'h00000000} /* (27, 27, 6) {real, imag} */,
  {32'h3fa4e7fe, 32'h00000000} /* (27, 27, 5) {real, imag} */,
  {32'h3f5bd677, 32'h00000000} /* (27, 27, 4) {real, imag} */,
  {32'h3f62c3ae, 32'h00000000} /* (27, 27, 3) {real, imag} */,
  {32'h3f855cf4, 32'h00000000} /* (27, 27, 2) {real, imag} */,
  {32'h3f569f59, 32'h00000000} /* (27, 27, 1) {real, imag} */,
  {32'h3f104047, 32'h00000000} /* (27, 27, 0) {real, imag} */,
  {32'h3f13e25f, 32'h00000000} /* (27, 26, 31) {real, imag} */,
  {32'h3f284b02, 32'h00000000} /* (27, 26, 30) {real, imag} */,
  {32'h3f02bf86, 32'h00000000} /* (27, 26, 29) {real, imag} */,
  {32'h3f06445a, 32'h00000000} /* (27, 26, 28) {real, imag} */,
  {32'h3f463b53, 32'h00000000} /* (27, 26, 27) {real, imag} */,
  {32'h3f81cb30, 32'h00000000} /* (27, 26, 26) {real, imag} */,
  {32'h3f515208, 32'h00000000} /* (27, 26, 25) {real, imag} */,
  {32'h3f47f9dd, 32'h00000000} /* (27, 26, 24) {real, imag} */,
  {32'h3f374c23, 32'h00000000} /* (27, 26, 23) {real, imag} */,
  {32'h3f5e5061, 32'h00000000} /* (27, 26, 22) {real, imag} */,
  {32'h3eddee16, 32'h00000000} /* (27, 26, 21) {real, imag} */,
  {32'hbf34fb3e, 32'h00000000} /* (27, 26, 20) {real, imag} */,
  {32'hbf42de3b, 32'h00000000} /* (27, 26, 19) {real, imag} */,
  {32'hbfc9f8b4, 32'h00000000} /* (27, 26, 18) {real, imag} */,
  {32'hbfc4b5fb, 32'h00000000} /* (27, 26, 17) {real, imag} */,
  {32'hbf7f1944, 32'h00000000} /* (27, 26, 16) {real, imag} */,
  {32'hbfb29bb5, 32'h00000000} /* (27, 26, 15) {real, imag} */,
  {32'hbf6830b4, 32'h00000000} /* (27, 26, 14) {real, imag} */,
  {32'hbf413e46, 32'h00000000} /* (27, 26, 13) {real, imag} */,
  {32'hbf83da50, 32'h00000000} /* (27, 26, 12) {real, imag} */,
  {32'hbf820760, 32'h00000000} /* (27, 26, 11) {real, imag} */,
  {32'hbe11a44e, 32'h00000000} /* (27, 26, 10) {real, imag} */,
  {32'h3f812a30, 32'h00000000} /* (27, 26, 9) {real, imag} */,
  {32'h3f900fe8, 32'h00000000} /* (27, 26, 8) {real, imag} */,
  {32'h3f10d52e, 32'h00000000} /* (27, 26, 7) {real, imag} */,
  {32'h3f024903, 32'h00000000} /* (27, 26, 6) {real, imag} */,
  {32'h3f4edbea, 32'h00000000} /* (27, 26, 5) {real, imag} */,
  {32'h3f0e67da, 32'h00000000} /* (27, 26, 4) {real, imag} */,
  {32'h3f1b5ad2, 32'h00000000} /* (27, 26, 3) {real, imag} */,
  {32'h3f522757, 32'h00000000} /* (27, 26, 2) {real, imag} */,
  {32'h3f2f8e72, 32'h00000000} /* (27, 26, 1) {real, imag} */,
  {32'h3eb9a76d, 32'h00000000} /* (27, 26, 0) {real, imag} */,
  {32'h3f0b8c6a, 32'h00000000} /* (27, 25, 31) {real, imag} */,
  {32'h3f3eaeaf, 32'h00000000} /* (27, 25, 30) {real, imag} */,
  {32'h3f2127a2, 32'h00000000} /* (27, 25, 29) {real, imag} */,
  {32'h3e8ef9ae, 32'h00000000} /* (27, 25, 28) {real, imag} */,
  {32'h3f2db75a, 32'h00000000} /* (27, 25, 27) {real, imag} */,
  {32'h3f372407, 32'h00000000} /* (27, 25, 26) {real, imag} */,
  {32'h3f241000, 32'h00000000} /* (27, 25, 25) {real, imag} */,
  {32'h3f7f47fa, 32'h00000000} /* (27, 25, 24) {real, imag} */,
  {32'h3f72af60, 32'h00000000} /* (27, 25, 23) {real, imag} */,
  {32'h3f4735f0, 32'h00000000} /* (27, 25, 22) {real, imag} */,
  {32'h3d4b112a, 32'h00000000} /* (27, 25, 21) {real, imag} */,
  {32'hbf41ef00, 32'h00000000} /* (27, 25, 20) {real, imag} */,
  {32'hbedff006, 32'h00000000} /* (27, 25, 19) {real, imag} */,
  {32'hbf392a13, 32'h00000000} /* (27, 25, 18) {real, imag} */,
  {32'hbf1f37d4, 32'h00000000} /* (27, 25, 17) {real, imag} */,
  {32'hbeae8c18, 32'h00000000} /* (27, 25, 16) {real, imag} */,
  {32'hbf9d61ec, 32'h00000000} /* (27, 25, 15) {real, imag} */,
  {32'hbfa4b510, 32'h00000000} /* (27, 25, 14) {real, imag} */,
  {32'hbed27af8, 32'h00000000} /* (27, 25, 13) {real, imag} */,
  {32'hbf591313, 32'h00000000} /* (27, 25, 12) {real, imag} */,
  {32'hbf61dc13, 32'h00000000} /* (27, 25, 11) {real, imag} */,
  {32'hbdcb469c, 32'h00000000} /* (27, 25, 10) {real, imag} */,
  {32'h3f542147, 32'h00000000} /* (27, 25, 9) {real, imag} */,
  {32'h3fd9b51a, 32'h00000000} /* (27, 25, 8) {real, imag} */,
  {32'h3f79830d, 32'h00000000} /* (27, 25, 7) {real, imag} */,
  {32'h3f20a4d4, 32'h00000000} /* (27, 25, 6) {real, imag} */,
  {32'h3f36eab2, 32'h00000000} /* (27, 25, 5) {real, imag} */,
  {32'h3f1065ad, 32'h00000000} /* (27, 25, 4) {real, imag} */,
  {32'h3eadc7f5, 32'h00000000} /* (27, 25, 3) {real, imag} */,
  {32'h3f10619d, 32'h00000000} /* (27, 25, 2) {real, imag} */,
  {32'h3ea32425, 32'h00000000} /* (27, 25, 1) {real, imag} */,
  {32'h3e15613b, 32'h00000000} /* (27, 25, 0) {real, imag} */,
  {32'h3e4d9df9, 32'h00000000} /* (27, 24, 31) {real, imag} */,
  {32'h3f63f03a, 32'h00000000} /* (27, 24, 30) {real, imag} */,
  {32'h3f892c89, 32'h00000000} /* (27, 24, 29) {real, imag} */,
  {32'h3f4beec7, 32'h00000000} /* (27, 24, 28) {real, imag} */,
  {32'h3fc39146, 32'h00000000} /* (27, 24, 27) {real, imag} */,
  {32'h3f9abaa6, 32'h00000000} /* (27, 24, 26) {real, imag} */,
  {32'h3f2c1587, 32'h00000000} /* (27, 24, 25) {real, imag} */,
  {32'h3f81b926, 32'h00000000} /* (27, 24, 24) {real, imag} */,
  {32'h3fb02593, 32'h00000000} /* (27, 24, 23) {real, imag} */,
  {32'h3f6c96fa, 32'h00000000} /* (27, 24, 22) {real, imag} */,
  {32'h3efba1e5, 32'h00000000} /* (27, 24, 21) {real, imag} */,
  {32'hbf004b28, 32'h00000000} /* (27, 24, 20) {real, imag} */,
  {32'hbf5dabc8, 32'h00000000} /* (27, 24, 19) {real, imag} */,
  {32'hbf2d4a57, 32'h00000000} /* (27, 24, 18) {real, imag} */,
  {32'hbe807218, 32'h00000000} /* (27, 24, 17) {real, imag} */,
  {32'hbf25d5b1, 32'h00000000} /* (27, 24, 16) {real, imag} */,
  {32'hbfc3bcc4, 32'h00000000} /* (27, 24, 15) {real, imag} */,
  {32'hbfbbe2ba, 32'h00000000} /* (27, 24, 14) {real, imag} */,
  {32'hbe8ff9ba, 32'h00000000} /* (27, 24, 13) {real, imag} */,
  {32'hbf830446, 32'h00000000} /* (27, 24, 12) {real, imag} */,
  {32'hbf9282be, 32'h00000000} /* (27, 24, 11) {real, imag} */,
  {32'h3e451e97, 32'h00000000} /* (27, 24, 10) {real, imag} */,
  {32'h3fa9c1b0, 32'h00000000} /* (27, 24, 9) {real, imag} */,
  {32'h4003e3db, 32'h00000000} /* (27, 24, 8) {real, imag} */,
  {32'h3f93932a, 32'h00000000} /* (27, 24, 7) {real, imag} */,
  {32'h3f691998, 32'h00000000} /* (27, 24, 6) {real, imag} */,
  {32'h3e9e202b, 32'h00000000} /* (27, 24, 5) {real, imag} */,
  {32'h3e6b4f6f, 32'h00000000} /* (27, 24, 4) {real, imag} */,
  {32'h3ea918cf, 32'h00000000} /* (27, 24, 3) {real, imag} */,
  {32'h3efa95c6, 32'h00000000} /* (27, 24, 2) {real, imag} */,
  {32'h3f23c738, 32'h00000000} /* (27, 24, 1) {real, imag} */,
  {32'h3e94edf2, 32'h00000000} /* (27, 24, 0) {real, imag} */,
  {32'h3e9e85ea, 32'h00000000} /* (27, 23, 31) {real, imag} */,
  {32'h3f856585, 32'h00000000} /* (27, 23, 30) {real, imag} */,
  {32'h3f8f30b2, 32'h00000000} /* (27, 23, 29) {real, imag} */,
  {32'h3f9772cf, 32'h00000000} /* (27, 23, 28) {real, imag} */,
  {32'h3ffa484e, 32'h00000000} /* (27, 23, 27) {real, imag} */,
  {32'h3fa8569d, 32'h00000000} /* (27, 23, 26) {real, imag} */,
  {32'h3f0755f5, 32'h00000000} /* (27, 23, 25) {real, imag} */,
  {32'h3f701711, 32'h00000000} /* (27, 23, 24) {real, imag} */,
  {32'h3fc8f8e4, 32'h00000000} /* (27, 23, 23) {real, imag} */,
  {32'h3faf9efa, 32'h00000000} /* (27, 23, 22) {real, imag} */,
  {32'h3f2d269f, 32'h00000000} /* (27, 23, 21) {real, imag} */,
  {32'hbed7f5df, 32'h00000000} /* (27, 23, 20) {real, imag} */,
  {32'hbf77a112, 32'h00000000} /* (27, 23, 19) {real, imag} */,
  {32'hbf87bbef, 32'h00000000} /* (27, 23, 18) {real, imag} */,
  {32'hbf3216d4, 32'h00000000} /* (27, 23, 17) {real, imag} */,
  {32'hbf385a6f, 32'h00000000} /* (27, 23, 16) {real, imag} */,
  {32'hbf71b621, 32'h00000000} /* (27, 23, 15) {real, imag} */,
  {32'hbfa4749f, 32'h00000000} /* (27, 23, 14) {real, imag} */,
  {32'hbf163295, 32'h00000000} /* (27, 23, 13) {real, imag} */,
  {32'hbf55e8fd, 32'h00000000} /* (27, 23, 12) {real, imag} */,
  {32'hbf2fc185, 32'h00000000} /* (27, 23, 11) {real, imag} */,
  {32'h3f456876, 32'h00000000} /* (27, 23, 10) {real, imag} */,
  {32'h3fa2de1e, 32'h00000000} /* (27, 23, 9) {real, imag} */,
  {32'h3fd38841, 32'h00000000} /* (27, 23, 8) {real, imag} */,
  {32'h3fa5e6ac, 32'h00000000} /* (27, 23, 7) {real, imag} */,
  {32'h3f551bf9, 32'h00000000} /* (27, 23, 6) {real, imag} */,
  {32'h3e8f69c9, 32'h00000000} /* (27, 23, 5) {real, imag} */,
  {32'h3ea04f79, 32'h00000000} /* (27, 23, 4) {real, imag} */,
  {32'h3f09fc4b, 32'h00000000} /* (27, 23, 3) {real, imag} */,
  {32'h3f3667b4, 32'h00000000} /* (27, 23, 2) {real, imag} */,
  {32'h3f0eb961, 32'h00000000} /* (27, 23, 1) {real, imag} */,
  {32'h3ee5aed6, 32'h00000000} /* (27, 23, 0) {real, imag} */,
  {32'h3f157848, 32'h00000000} /* (27, 22, 31) {real, imag} */,
  {32'h3f92b718, 32'h00000000} /* (27, 22, 30) {real, imag} */,
  {32'h3f9392e8, 32'h00000000} /* (27, 22, 29) {real, imag} */,
  {32'h3f86ab45, 32'h00000000} /* (27, 22, 28) {real, imag} */,
  {32'h3f90cbf0, 32'h00000000} /* (27, 22, 27) {real, imag} */,
  {32'h3f8856c6, 32'h00000000} /* (27, 22, 26) {real, imag} */,
  {32'h3ee26b5b, 32'h00000000} /* (27, 22, 25) {real, imag} */,
  {32'h3ec82c8b, 32'h00000000} /* (27, 22, 24) {real, imag} */,
  {32'h3f23387b, 32'h00000000} /* (27, 22, 23) {real, imag} */,
  {32'h3f41119a, 32'h00000000} /* (27, 22, 22) {real, imag} */,
  {32'h3d82d23e, 32'h00000000} /* (27, 22, 21) {real, imag} */,
  {32'hbf5b3f59, 32'h00000000} /* (27, 22, 20) {real, imag} */,
  {32'hbf548c46, 32'h00000000} /* (27, 22, 19) {real, imag} */,
  {32'hbf42bb05, 32'h00000000} /* (27, 22, 18) {real, imag} */,
  {32'hbf34bbbf, 32'h00000000} /* (27, 22, 17) {real, imag} */,
  {32'hbf32a690, 32'h00000000} /* (27, 22, 16) {real, imag} */,
  {32'hbee1a13e, 32'h00000000} /* (27, 22, 15) {real, imag} */,
  {32'hbf127db7, 32'h00000000} /* (27, 22, 14) {real, imag} */,
  {32'hbf50e70c, 32'h00000000} /* (27, 22, 13) {real, imag} */,
  {32'hbedbf2a3, 32'h00000000} /* (27, 22, 12) {real, imag} */,
  {32'hbc5ec156, 32'h00000000} /* (27, 22, 11) {real, imag} */,
  {32'h3f461734, 32'h00000000} /* (27, 22, 10) {real, imag} */,
  {32'h3f47f1ad, 32'h00000000} /* (27, 22, 9) {real, imag} */,
  {32'h3f628b5e, 32'h00000000} /* (27, 22, 8) {real, imag} */,
  {32'h3f93b6a2, 32'h00000000} /* (27, 22, 7) {real, imag} */,
  {32'h3f6ddfd0, 32'h00000000} /* (27, 22, 6) {real, imag} */,
  {32'h3f21870a, 32'h00000000} /* (27, 22, 5) {real, imag} */,
  {32'h3f365bc2, 32'h00000000} /* (27, 22, 4) {real, imag} */,
  {32'h3f976392, 32'h00000000} /* (27, 22, 3) {real, imag} */,
  {32'h3f6e12f5, 32'h00000000} /* (27, 22, 2) {real, imag} */,
  {32'h3f55ae32, 32'h00000000} /* (27, 22, 1) {real, imag} */,
  {32'h3f5d15e4, 32'h00000000} /* (27, 22, 0) {real, imag} */,
  {32'h3e72a915, 32'h00000000} /* (27, 21, 31) {real, imag} */,
  {32'h3e8d752a, 32'h00000000} /* (27, 21, 30) {real, imag} */,
  {32'h3e8594a2, 32'h00000000} /* (27, 21, 29) {real, imag} */,
  {32'h3e3552e9, 32'h00000000} /* (27, 21, 28) {real, imag} */,
  {32'h3f0ddc70, 32'h00000000} /* (27, 21, 27) {real, imag} */,
  {32'h3f05ed94, 32'h00000000} /* (27, 21, 26) {real, imag} */,
  {32'hbe7c5ca6, 32'h00000000} /* (27, 21, 25) {real, imag} */,
  {32'hbe4f4c6a, 32'h00000000} /* (27, 21, 24) {real, imag} */,
  {32'hbe4f1e89, 32'h00000000} /* (27, 21, 23) {real, imag} */,
  {32'hbdeae889, 32'h00000000} /* (27, 21, 22) {real, imag} */,
  {32'h3cd54f70, 32'h00000000} /* (27, 21, 21) {real, imag} */,
  {32'hbe1e8d61, 32'h00000000} /* (27, 21, 20) {real, imag} */,
  {32'h3dd51f85, 32'h00000000} /* (27, 21, 19) {real, imag} */,
  {32'h3efa40ed, 32'h00000000} /* (27, 21, 18) {real, imag} */,
  {32'h3e52c0a2, 32'h00000000} /* (27, 21, 17) {real, imag} */,
  {32'hbeec11ed, 32'h00000000} /* (27, 21, 16) {real, imag} */,
  {32'hbeb8336d, 32'h00000000} /* (27, 21, 15) {real, imag} */,
  {32'h3b909fdf, 32'h00000000} /* (27, 21, 14) {real, imag} */,
  {32'hbcc32e68, 32'h00000000} /* (27, 21, 13) {real, imag} */,
  {32'hbec1780a, 32'h00000000} /* (27, 21, 12) {real, imag} */,
  {32'hbe112c3e, 32'h00000000} /* (27, 21, 11) {real, imag} */,
  {32'h3f1facff, 32'h00000000} /* (27, 21, 10) {real, imag} */,
  {32'h3f78529b, 32'h00000000} /* (27, 21, 9) {real, imag} */,
  {32'h3e3ba6e5, 32'h00000000} /* (27, 21, 8) {real, imag} */,
  {32'h3e73c9e5, 32'h00000000} /* (27, 21, 7) {real, imag} */,
  {32'h3f43b751, 32'h00000000} /* (27, 21, 6) {real, imag} */,
  {32'h3eb8ffdc, 32'h00000000} /* (27, 21, 5) {real, imag} */,
  {32'h3ea47756, 32'h00000000} /* (27, 21, 4) {real, imag} */,
  {32'h3f60bba1, 32'h00000000} /* (27, 21, 3) {real, imag} */,
  {32'h3efc9963, 32'h00000000} /* (27, 21, 2) {real, imag} */,
  {32'h3ea669b0, 32'h00000000} /* (27, 21, 1) {real, imag} */,
  {32'h3eb582a2, 32'h00000000} /* (27, 21, 0) {real, imag} */,
  {32'hbe40d3f1, 32'h00000000} /* (27, 20, 31) {real, imag} */,
  {32'hbe85f6ec, 32'h00000000} /* (27, 20, 30) {real, imag} */,
  {32'hbf0b08ef, 32'h00000000} /* (27, 20, 29) {real, imag} */,
  {32'hbf764df1, 32'h00000000} /* (27, 20, 28) {real, imag} */,
  {32'hbecfe741, 32'h00000000} /* (27, 20, 27) {real, imag} */,
  {32'hbe8f1cf8, 32'h00000000} /* (27, 20, 26) {real, imag} */,
  {32'hbf999360, 32'h00000000} /* (27, 20, 25) {real, imag} */,
  {32'hbf752cc1, 32'h00000000} /* (27, 20, 24) {real, imag} */,
  {32'hbeebd504, 32'h00000000} /* (27, 20, 23) {real, imag} */,
  {32'hbf2bda5e, 32'h00000000} /* (27, 20, 22) {real, imag} */,
  {32'hbe497b1a, 32'h00000000} /* (27, 20, 21) {real, imag} */,
  {32'h3ea80fda, 32'h00000000} /* (27, 20, 20) {real, imag} */,
  {32'h3f269d84, 32'h00000000} /* (27, 20, 19) {real, imag} */,
  {32'h3fb78304, 32'h00000000} /* (27, 20, 18) {real, imag} */,
  {32'h3f8e9b7e, 32'h00000000} /* (27, 20, 17) {real, imag} */,
  {32'h3f6fc998, 32'h00000000} /* (27, 20, 16) {real, imag} */,
  {32'h3f373293, 32'h00000000} /* (27, 20, 15) {real, imag} */,
  {32'h3f360fa5, 32'h00000000} /* (27, 20, 14) {real, imag} */,
  {32'h3f28b725, 32'h00000000} /* (27, 20, 13) {real, imag} */,
  {32'h3e86eda7, 32'h00000000} /* (27, 20, 12) {real, imag} */,
  {32'h3d796220, 32'h00000000} /* (27, 20, 11) {real, imag} */,
  {32'hbe368d50, 32'h00000000} /* (27, 20, 10) {real, imag} */,
  {32'hbd5491eb, 32'h00000000} /* (27, 20, 9) {real, imag} */,
  {32'hbef378ca, 32'h00000000} /* (27, 20, 8) {real, imag} */,
  {32'hbf1bbbd6, 32'h00000000} /* (27, 20, 7) {real, imag} */,
  {32'hbed6c16f, 32'h00000000} /* (27, 20, 6) {real, imag} */,
  {32'hbf4d5baf, 32'h00000000} /* (27, 20, 5) {real, imag} */,
  {32'hbf1aea31, 32'h00000000} /* (27, 20, 4) {real, imag} */,
  {32'hbf10e4b4, 32'h00000000} /* (27, 20, 3) {real, imag} */,
  {32'hbf73cbd8, 32'h00000000} /* (27, 20, 2) {real, imag} */,
  {32'hbf1aa080, 32'h00000000} /* (27, 20, 1) {real, imag} */,
  {32'hbe6a0bec, 32'h00000000} /* (27, 20, 0) {real, imag} */,
  {32'hbee20c43, 32'h00000000} /* (27, 19, 31) {real, imag} */,
  {32'hbee8de22, 32'h00000000} /* (27, 19, 30) {real, imag} */,
  {32'hbf01b3d3, 32'h00000000} /* (27, 19, 29) {real, imag} */,
  {32'hbf239a5c, 32'h00000000} /* (27, 19, 28) {real, imag} */,
  {32'hbf607e6e, 32'h00000000} /* (27, 19, 27) {real, imag} */,
  {32'hbf27cf18, 32'h00000000} /* (27, 19, 26) {real, imag} */,
  {32'hbf374ae7, 32'h00000000} /* (27, 19, 25) {real, imag} */,
  {32'hbf93f442, 32'h00000000} /* (27, 19, 24) {real, imag} */,
  {32'hbf76c5d4, 32'h00000000} /* (27, 19, 23) {real, imag} */,
  {32'hbf38d783, 32'h00000000} /* (27, 19, 22) {real, imag} */,
  {32'hbdd8adfb, 32'h00000000} /* (27, 19, 21) {real, imag} */,
  {32'h3f1f9c99, 32'h00000000} /* (27, 19, 20) {real, imag} */,
  {32'h3f23c6e3, 32'h00000000} /* (27, 19, 19) {real, imag} */,
  {32'h3f52ac06, 32'h00000000} /* (27, 19, 18) {real, imag} */,
  {32'h3f4df76f, 32'h00000000} /* (27, 19, 17) {real, imag} */,
  {32'h3f98eada, 32'h00000000} /* (27, 19, 16) {real, imag} */,
  {32'h3fbbb5ec, 32'h00000000} /* (27, 19, 15) {real, imag} */,
  {32'h3f890e0b, 32'h00000000} /* (27, 19, 14) {real, imag} */,
  {32'h3f7fefcd, 32'h00000000} /* (27, 19, 13) {real, imag} */,
  {32'h3f0ea4ce, 32'h00000000} /* (27, 19, 12) {real, imag} */,
  {32'h3ee9eb46, 32'h00000000} /* (27, 19, 11) {real, imag} */,
  {32'hbc485ae8, 32'h00000000} /* (27, 19, 10) {real, imag} */,
  {32'hbe911dbf, 32'h00000000} /* (27, 19, 9) {real, imag} */,
  {32'hbf0b200a, 32'h00000000} /* (27, 19, 8) {real, imag} */,
  {32'hbf00b770, 32'h00000000} /* (27, 19, 7) {real, imag} */,
  {32'hbef6b3c0, 32'h00000000} /* (27, 19, 6) {real, imag} */,
  {32'hbf96d720, 32'h00000000} /* (27, 19, 5) {real, imag} */,
  {32'hbf684fe1, 32'h00000000} /* (27, 19, 4) {real, imag} */,
  {32'hbf76841f, 32'h00000000} /* (27, 19, 3) {real, imag} */,
  {32'hbfab684d, 32'h00000000} /* (27, 19, 2) {real, imag} */,
  {32'hbedbe79a, 32'h00000000} /* (27, 19, 1) {real, imag} */,
  {32'hbe6e06af, 32'h00000000} /* (27, 19, 0) {real, imag} */,
  {32'hbeb97a18, 32'h00000000} /* (27, 18, 31) {real, imag} */,
  {32'hbf533cbe, 32'h00000000} /* (27, 18, 30) {real, imag} */,
  {32'hbf61a91b, 32'h00000000} /* (27, 18, 29) {real, imag} */,
  {32'hbf2197ad, 32'h00000000} /* (27, 18, 28) {real, imag} */,
  {32'hbf61a5b6, 32'h00000000} /* (27, 18, 27) {real, imag} */,
  {32'hbf4ca37b, 32'h00000000} /* (27, 18, 26) {real, imag} */,
  {32'hbf6d5600, 32'h00000000} /* (27, 18, 25) {real, imag} */,
  {32'hbfb57bbe, 32'h00000000} /* (27, 18, 24) {real, imag} */,
  {32'hbfb0971f, 32'h00000000} /* (27, 18, 23) {real, imag} */,
  {32'hbf8c0eb0, 32'h00000000} /* (27, 18, 22) {real, imag} */,
  {32'hbec390f3, 32'h00000000} /* (27, 18, 21) {real, imag} */,
  {32'h3dbe8582, 32'h00000000} /* (27, 18, 20) {real, imag} */,
  {32'h3ebbb8de, 32'h00000000} /* (27, 18, 19) {real, imag} */,
  {32'h3f57d353, 32'h00000000} /* (27, 18, 18) {real, imag} */,
  {32'h3f70834b, 32'h00000000} /* (27, 18, 17) {real, imag} */,
  {32'h3f88bf5a, 32'h00000000} /* (27, 18, 16) {real, imag} */,
  {32'h3f8646ac, 32'h00000000} /* (27, 18, 15) {real, imag} */,
  {32'h3f8306b8, 32'h00000000} /* (27, 18, 14) {real, imag} */,
  {32'h3fada42f, 32'h00000000} /* (27, 18, 13) {real, imag} */,
  {32'h3f4de3fd, 32'h00000000} /* (27, 18, 12) {real, imag} */,
  {32'h3f4ce35d, 32'h00000000} /* (27, 18, 11) {real, imag} */,
  {32'h3de91588, 32'h00000000} /* (27, 18, 10) {real, imag} */,
  {32'hbe88d3e0, 32'h00000000} /* (27, 18, 9) {real, imag} */,
  {32'hbf0c1a18, 32'h00000000} /* (27, 18, 8) {real, imag} */,
  {32'hbf3f45d5, 32'h00000000} /* (27, 18, 7) {real, imag} */,
  {32'hbfbc5e1b, 32'h00000000} /* (27, 18, 6) {real, imag} */,
  {32'hbfbbb5f0, 32'h00000000} /* (27, 18, 5) {real, imag} */,
  {32'hbf6258ca, 32'h00000000} /* (27, 18, 4) {real, imag} */,
  {32'hbf4f3f49, 32'h00000000} /* (27, 18, 3) {real, imag} */,
  {32'hbedddb2b, 32'h00000000} /* (27, 18, 2) {real, imag} */,
  {32'hbdd74b01, 32'h00000000} /* (27, 18, 1) {real, imag} */,
  {32'hbdc408fa, 32'h00000000} /* (27, 18, 0) {real, imag} */,
  {32'hbe9123ad, 32'h00000000} /* (27, 17, 31) {real, imag} */,
  {32'hbf951007, 32'h00000000} /* (27, 17, 30) {real, imag} */,
  {32'hbfb524f0, 32'h00000000} /* (27, 17, 29) {real, imag} */,
  {32'hbf7ffe48, 32'h00000000} /* (27, 17, 28) {real, imag} */,
  {32'hbf561f6f, 32'h00000000} /* (27, 17, 27) {real, imag} */,
  {32'hbec0b84f, 32'h00000000} /* (27, 17, 26) {real, imag} */,
  {32'hbf91504f, 32'h00000000} /* (27, 17, 25) {real, imag} */,
  {32'hbfb9760e, 32'h00000000} /* (27, 17, 24) {real, imag} */,
  {32'hbfbcde51, 32'h00000000} /* (27, 17, 23) {real, imag} */,
  {32'hbf5785e4, 32'h00000000} /* (27, 17, 22) {real, imag} */,
  {32'hbf3191b4, 32'h00000000} /* (27, 17, 21) {real, imag} */,
  {32'h3dd87b64, 32'h00000000} /* (27, 17, 20) {real, imag} */,
  {32'h3f325164, 32'h00000000} /* (27, 17, 19) {real, imag} */,
  {32'h3f970e57, 32'h00000000} /* (27, 17, 18) {real, imag} */,
  {32'h3fc90e70, 32'h00000000} /* (27, 17, 17) {real, imag} */,
  {32'h3f6d667f, 32'h00000000} /* (27, 17, 16) {real, imag} */,
  {32'h3f10210b, 32'h00000000} /* (27, 17, 15) {real, imag} */,
  {32'h3f63eeb6, 32'h00000000} /* (27, 17, 14) {real, imag} */,
  {32'h3f502bf7, 32'h00000000} /* (27, 17, 13) {real, imag} */,
  {32'h3f16b7f4, 32'h00000000} /* (27, 17, 12) {real, imag} */,
  {32'h3f362457, 32'h00000000} /* (27, 17, 11) {real, imag} */,
  {32'hbcefb788, 32'h00000000} /* (27, 17, 10) {real, imag} */,
  {32'hbebe0b03, 32'h00000000} /* (27, 17, 9) {real, imag} */,
  {32'hbf01db93, 32'h00000000} /* (27, 17, 8) {real, imag} */,
  {32'hbf332a00, 32'h00000000} /* (27, 17, 7) {real, imag} */,
  {32'hbfab4a3d, 32'h00000000} /* (27, 17, 6) {real, imag} */,
  {32'hbf7c1fff, 32'h00000000} /* (27, 17, 5) {real, imag} */,
  {32'hbf62ca81, 32'h00000000} /* (27, 17, 4) {real, imag} */,
  {32'hbf7e4fb1, 32'h00000000} /* (27, 17, 3) {real, imag} */,
  {32'hbf833455, 32'h00000000} /* (27, 17, 2) {real, imag} */,
  {32'hbe926d83, 32'h00000000} /* (27, 17, 1) {real, imag} */,
  {32'h3dcb040e, 32'h00000000} /* (27, 17, 0) {real, imag} */,
  {32'hbeb8cc74, 32'h00000000} /* (27, 16, 31) {real, imag} */,
  {32'hbf861c78, 32'h00000000} /* (27, 16, 30) {real, imag} */,
  {32'hbfa083be, 32'h00000000} /* (27, 16, 29) {real, imag} */,
  {32'hbf62dacd, 32'h00000000} /* (27, 16, 28) {real, imag} */,
  {32'hbf5371fc, 32'h00000000} /* (27, 16, 27) {real, imag} */,
  {32'hbf47db73, 32'h00000000} /* (27, 16, 26) {real, imag} */,
  {32'hbfb3a791, 32'h00000000} /* (27, 16, 25) {real, imag} */,
  {32'hbf8912c7, 32'h00000000} /* (27, 16, 24) {real, imag} */,
  {32'hbf8cd0b7, 32'h00000000} /* (27, 16, 23) {real, imag} */,
  {32'hbf4475be, 32'h00000000} /* (27, 16, 22) {real, imag} */,
  {32'hbe12abbc, 32'h00000000} /* (27, 16, 21) {real, imag} */,
  {32'h3f45a671, 32'h00000000} /* (27, 16, 20) {real, imag} */,
  {32'h3f78f8b6, 32'h00000000} /* (27, 16, 19) {real, imag} */,
  {32'h3f6ca032, 32'h00000000} /* (27, 16, 18) {real, imag} */,
  {32'h3f83ebd2, 32'h00000000} /* (27, 16, 17) {real, imag} */,
  {32'h3f35ef6d, 32'h00000000} /* (27, 16, 16) {real, imag} */,
  {32'h3f2fff9b, 32'h00000000} /* (27, 16, 15) {real, imag} */,
  {32'h3f07beca, 32'h00000000} /* (27, 16, 14) {real, imag} */,
  {32'h3f378048, 32'h00000000} /* (27, 16, 13) {real, imag} */,
  {32'h3f5225cb, 32'h00000000} /* (27, 16, 12) {real, imag} */,
  {32'h3f33e609, 32'h00000000} /* (27, 16, 11) {real, imag} */,
  {32'hbe8d2ed8, 32'h00000000} /* (27, 16, 10) {real, imag} */,
  {32'hbeee986c, 32'h00000000} /* (27, 16, 9) {real, imag} */,
  {32'hbf143ffa, 32'h00000000} /* (27, 16, 8) {real, imag} */,
  {32'hbf4b193a, 32'h00000000} /* (27, 16, 7) {real, imag} */,
  {32'hbf83f259, 32'h00000000} /* (27, 16, 6) {real, imag} */,
  {32'hbf66d86f, 32'h00000000} /* (27, 16, 5) {real, imag} */,
  {32'hbf8f50f4, 32'h00000000} /* (27, 16, 4) {real, imag} */,
  {32'hbf6d1557, 32'h00000000} /* (27, 16, 3) {real, imag} */,
  {32'hbf473029, 32'h00000000} /* (27, 16, 2) {real, imag} */,
  {32'hbf41fad3, 32'h00000000} /* (27, 16, 1) {real, imag} */,
  {32'hbecf731b, 32'h00000000} /* (27, 16, 0) {real, imag} */,
  {32'hbf1d6bc8, 32'h00000000} /* (27, 15, 31) {real, imag} */,
  {32'hbf6bc8f5, 32'h00000000} /* (27, 15, 30) {real, imag} */,
  {32'hbf83fef9, 32'h00000000} /* (27, 15, 29) {real, imag} */,
  {32'hbf828c48, 32'h00000000} /* (27, 15, 28) {real, imag} */,
  {32'hbf8103ad, 32'h00000000} /* (27, 15, 27) {real, imag} */,
  {32'hbfa785f3, 32'h00000000} /* (27, 15, 26) {real, imag} */,
  {32'hbfb4712a, 32'h00000000} /* (27, 15, 25) {real, imag} */,
  {32'hbf53b9bb, 32'h00000000} /* (27, 15, 24) {real, imag} */,
  {32'hbf5647a9, 32'h00000000} /* (27, 15, 23) {real, imag} */,
  {32'hbfcebd6b, 32'h00000000} /* (27, 15, 22) {real, imag} */,
  {32'hbf05771d, 32'h00000000} /* (27, 15, 21) {real, imag} */,
  {32'h3f2eb0d8, 32'h00000000} /* (27, 15, 20) {real, imag} */,
  {32'h3f564b98, 32'h00000000} /* (27, 15, 19) {real, imag} */,
  {32'h3f1df77e, 32'h00000000} /* (27, 15, 18) {real, imag} */,
  {32'h3f0742e0, 32'h00000000} /* (27, 15, 17) {real, imag} */,
  {32'h3f30a748, 32'h00000000} /* (27, 15, 16) {real, imag} */,
  {32'h3f526fac, 32'h00000000} /* (27, 15, 15) {real, imag} */,
  {32'h3e94e02d, 32'h00000000} /* (27, 15, 14) {real, imag} */,
  {32'h3ef60424, 32'h00000000} /* (27, 15, 13) {real, imag} */,
  {32'h3f08f437, 32'h00000000} /* (27, 15, 12) {real, imag} */,
  {32'h3f50fe85, 32'h00000000} /* (27, 15, 11) {real, imag} */,
  {32'hbee07239, 32'h00000000} /* (27, 15, 10) {real, imag} */,
  {32'hbf5f9894, 32'h00000000} /* (27, 15, 9) {real, imag} */,
  {32'hbf5e41f4, 32'h00000000} /* (27, 15, 8) {real, imag} */,
  {32'hbf8b82b4, 32'h00000000} /* (27, 15, 7) {real, imag} */,
  {32'hbf8bdf82, 32'h00000000} /* (27, 15, 6) {real, imag} */,
  {32'hbf9121b2, 32'h00000000} /* (27, 15, 5) {real, imag} */,
  {32'hbf6a6568, 32'h00000000} /* (27, 15, 4) {real, imag} */,
  {32'hbf4a7810, 32'h00000000} /* (27, 15, 3) {real, imag} */,
  {32'hbf12fe4a, 32'h00000000} /* (27, 15, 2) {real, imag} */,
  {32'hbf530752, 32'h00000000} /* (27, 15, 1) {real, imag} */,
  {32'hbedfe02a, 32'h00000000} /* (27, 15, 0) {real, imag} */,
  {32'hbf1edd34, 32'h00000000} /* (27, 14, 31) {real, imag} */,
  {32'hbf9f0b8a, 32'h00000000} /* (27, 14, 30) {real, imag} */,
  {32'hbf7fade0, 32'h00000000} /* (27, 14, 29) {real, imag} */,
  {32'hbf9670c9, 32'h00000000} /* (27, 14, 28) {real, imag} */,
  {32'hbf900527, 32'h00000000} /* (27, 14, 27) {real, imag} */,
  {32'hbf6ce332, 32'h00000000} /* (27, 14, 26) {real, imag} */,
  {32'hbf9ab58b, 32'h00000000} /* (27, 14, 25) {real, imag} */,
  {32'hbf99981d, 32'h00000000} /* (27, 14, 24) {real, imag} */,
  {32'hbfa5db24, 32'h00000000} /* (27, 14, 23) {real, imag} */,
  {32'hbfb71c3a, 32'h00000000} /* (27, 14, 22) {real, imag} */,
  {32'hbedab973, 32'h00000000} /* (27, 14, 21) {real, imag} */,
  {32'h3ed3d4e5, 32'h00000000} /* (27, 14, 20) {real, imag} */,
  {32'h3f45faba, 32'h00000000} /* (27, 14, 19) {real, imag} */,
  {32'h3f7ed1c5, 32'h00000000} /* (27, 14, 18) {real, imag} */,
  {32'h3f1475a3, 32'h00000000} /* (27, 14, 17) {real, imag} */,
  {32'h3f36933b, 32'h00000000} /* (27, 14, 16) {real, imag} */,
  {32'h3f4f6e07, 32'h00000000} /* (27, 14, 15) {real, imag} */,
  {32'h3ef467be, 32'h00000000} /* (27, 14, 14) {real, imag} */,
  {32'h3f10ce08, 32'h00000000} /* (27, 14, 13) {real, imag} */,
  {32'h3f4b895d, 32'h00000000} /* (27, 14, 12) {real, imag} */,
  {32'h3f29a807, 32'h00000000} /* (27, 14, 11) {real, imag} */,
  {32'hbea7c66b, 32'h00000000} /* (27, 14, 10) {real, imag} */,
  {32'hbf7a1ec1, 32'h00000000} /* (27, 14, 9) {real, imag} */,
  {32'hbf76b215, 32'h00000000} /* (27, 14, 8) {real, imag} */,
  {32'hbf967fd1, 32'h00000000} /* (27, 14, 7) {real, imag} */,
  {32'hbf09f751, 32'h00000000} /* (27, 14, 6) {real, imag} */,
  {32'hbef87496, 32'h00000000} /* (27, 14, 5) {real, imag} */,
  {32'hbf0dd8a7, 32'h00000000} /* (27, 14, 4) {real, imag} */,
  {32'hbf1bf04e, 32'h00000000} /* (27, 14, 3) {real, imag} */,
  {32'hbf32aefb, 32'h00000000} /* (27, 14, 2) {real, imag} */,
  {32'hbf4639cb, 32'h00000000} /* (27, 14, 1) {real, imag} */,
  {32'hbd010200, 32'h00000000} /* (27, 14, 0) {real, imag} */,
  {32'hbf47ab2c, 32'h00000000} /* (27, 13, 31) {real, imag} */,
  {32'hbfa14da1, 32'h00000000} /* (27, 13, 30) {real, imag} */,
  {32'hbf84455c, 32'h00000000} /* (27, 13, 29) {real, imag} */,
  {32'hbf56915c, 32'h00000000} /* (27, 13, 28) {real, imag} */,
  {32'hbf1d9db9, 32'h00000000} /* (27, 13, 27) {real, imag} */,
  {32'hbed8d507, 32'h00000000} /* (27, 13, 26) {real, imag} */,
  {32'hbf6533a8, 32'h00000000} /* (27, 13, 25) {real, imag} */,
  {32'hbf73c19b, 32'h00000000} /* (27, 13, 24) {real, imag} */,
  {32'hbf4fe519, 32'h00000000} /* (27, 13, 23) {real, imag} */,
  {32'hbf3dff46, 32'h00000000} /* (27, 13, 22) {real, imag} */,
  {32'hbf027be7, 32'h00000000} /* (27, 13, 21) {real, imag} */,
  {32'h3d2b70fc, 32'h00000000} /* (27, 13, 20) {real, imag} */,
  {32'h3ea3c0ad, 32'h00000000} /* (27, 13, 19) {real, imag} */,
  {32'h3f834f0f, 32'h00000000} /* (27, 13, 18) {real, imag} */,
  {32'h3f7647ea, 32'h00000000} /* (27, 13, 17) {real, imag} */,
  {32'h3f1ea4e2, 32'h00000000} /* (27, 13, 16) {real, imag} */,
  {32'h3ebf2574, 32'h00000000} /* (27, 13, 15) {real, imag} */,
  {32'h3ef13ffe, 32'h00000000} /* (27, 13, 14) {real, imag} */,
  {32'h3f09afba, 32'h00000000} /* (27, 13, 13) {real, imag} */,
  {32'h3f2f3fe4, 32'h00000000} /* (27, 13, 12) {real, imag} */,
  {32'h3f2ccb46, 32'h00000000} /* (27, 13, 11) {real, imag} */,
  {32'hbed68e54, 32'h00000000} /* (27, 13, 10) {real, imag} */,
  {32'hbf956195, 32'h00000000} /* (27, 13, 9) {real, imag} */,
  {32'hbf665edc, 32'h00000000} /* (27, 13, 8) {real, imag} */,
  {32'hbfb399a4, 32'h00000000} /* (27, 13, 7) {real, imag} */,
  {32'hbf3c5fe7, 32'h00000000} /* (27, 13, 6) {real, imag} */,
  {32'hbe4d979f, 32'h00000000} /* (27, 13, 5) {real, imag} */,
  {32'hbec492be, 32'h00000000} /* (27, 13, 4) {real, imag} */,
  {32'hbf52d40b, 32'h00000000} /* (27, 13, 3) {real, imag} */,
  {32'hbf3d05e7, 32'h00000000} /* (27, 13, 2) {real, imag} */,
  {32'hbee74774, 32'h00000000} /* (27, 13, 1) {real, imag} */,
  {32'hbe042d06, 32'h00000000} /* (27, 13, 0) {real, imag} */,
  {32'hbf27ced6, 32'h00000000} /* (27, 12, 31) {real, imag} */,
  {32'hbf7265e5, 32'h00000000} /* (27, 12, 30) {real, imag} */,
  {32'hbf2dbb44, 32'h00000000} /* (27, 12, 29) {real, imag} */,
  {32'hbf6f0e3a, 32'h00000000} /* (27, 12, 28) {real, imag} */,
  {32'hbf4d3af1, 32'h00000000} /* (27, 12, 27) {real, imag} */,
  {32'hbf664a5e, 32'h00000000} /* (27, 12, 26) {real, imag} */,
  {32'hbf99ed0b, 32'h00000000} /* (27, 12, 25) {real, imag} */,
  {32'hbf2a487e, 32'h00000000} /* (27, 12, 24) {real, imag} */,
  {32'hbf11b5ab, 32'h00000000} /* (27, 12, 23) {real, imag} */,
  {32'hbf82fdb0, 32'h00000000} /* (27, 12, 22) {real, imag} */,
  {32'hbe3e16ac, 32'h00000000} /* (27, 12, 21) {real, imag} */,
  {32'h3dc81ba3, 32'h00000000} /* (27, 12, 20) {real, imag} */,
  {32'h3e0f6313, 32'h00000000} /* (27, 12, 19) {real, imag} */,
  {32'h3f70c85f, 32'h00000000} /* (27, 12, 18) {real, imag} */,
  {32'h3f99824d, 32'h00000000} /* (27, 12, 17) {real, imag} */,
  {32'h3ef0e2a8, 32'h00000000} /* (27, 12, 16) {real, imag} */,
  {32'h3ea631ec, 32'h00000000} /* (27, 12, 15) {real, imag} */,
  {32'h3f49c9b9, 32'h00000000} /* (27, 12, 14) {real, imag} */,
  {32'h3f32581d, 32'h00000000} /* (27, 12, 13) {real, imag} */,
  {32'h3e328f03, 32'h00000000} /* (27, 12, 12) {real, imag} */,
  {32'h3f19ebc5, 32'h00000000} /* (27, 12, 11) {real, imag} */,
  {32'hbe66d780, 32'h00000000} /* (27, 12, 10) {real, imag} */,
  {32'hbf4e8eb0, 32'h00000000} /* (27, 12, 9) {real, imag} */,
  {32'hbf178f3c, 32'h00000000} /* (27, 12, 8) {real, imag} */,
  {32'hbf6c9ba6, 32'h00000000} /* (27, 12, 7) {real, imag} */,
  {32'hbf91d87d, 32'h00000000} /* (27, 12, 6) {real, imag} */,
  {32'hbf35fc00, 32'h00000000} /* (27, 12, 5) {real, imag} */,
  {32'hbef7e69c, 32'h00000000} /* (27, 12, 4) {real, imag} */,
  {32'hbf5512e5, 32'h00000000} /* (27, 12, 3) {real, imag} */,
  {32'hbf3fedb6, 32'h00000000} /* (27, 12, 2) {real, imag} */,
  {32'hbf29b4d8, 32'h00000000} /* (27, 12, 1) {real, imag} */,
  {32'hbe9ac979, 32'h00000000} /* (27, 12, 0) {real, imag} */,
  {32'hbe44afe7, 32'h00000000} /* (27, 11, 31) {real, imag} */,
  {32'hbe3e9798, 32'h00000000} /* (27, 11, 30) {real, imag} */,
  {32'hbee88f0e, 32'h00000000} /* (27, 11, 29) {real, imag} */,
  {32'hbf67946c, 32'h00000000} /* (27, 11, 28) {real, imag} */,
  {32'hbf04add6, 32'h00000000} /* (27, 11, 27) {real, imag} */,
  {32'hbf28234d, 32'h00000000} /* (27, 11, 26) {real, imag} */,
  {32'hbf8041dd, 32'h00000000} /* (27, 11, 25) {real, imag} */,
  {32'hbf03509a, 32'h00000000} /* (27, 11, 24) {real, imag} */,
  {32'hbe83cc01, 32'h00000000} /* (27, 11, 23) {real, imag} */,
  {32'hbf06ee70, 32'h00000000} /* (27, 11, 22) {real, imag} */,
  {32'h3e9e65bc, 32'h00000000} /* (27, 11, 21) {real, imag} */,
  {32'h3efe22bc, 32'h00000000} /* (27, 11, 20) {real, imag} */,
  {32'h3d40534c, 32'h00000000} /* (27, 11, 19) {real, imag} */,
  {32'h3f56d3e4, 32'h00000000} /* (27, 11, 18) {real, imag} */,
  {32'h3fa1dbe5, 32'h00000000} /* (27, 11, 17) {real, imag} */,
  {32'h3eb7edfc, 32'h00000000} /* (27, 11, 16) {real, imag} */,
  {32'h3f2a101b, 32'h00000000} /* (27, 11, 15) {real, imag} */,
  {32'h3f896ccb, 32'h00000000} /* (27, 11, 14) {real, imag} */,
  {32'h3f496a30, 32'h00000000} /* (27, 11, 13) {real, imag} */,
  {32'h3e6e591d, 32'h00000000} /* (27, 11, 12) {real, imag} */,
  {32'hbd018581, 32'h00000000} /* (27, 11, 11) {real, imag} */,
  {32'hbef58f23, 32'h00000000} /* (27, 11, 10) {real, imag} */,
  {32'hbf19d391, 32'h00000000} /* (27, 11, 9) {real, imag} */,
  {32'hbeee0acc, 32'h00000000} /* (27, 11, 8) {real, imag} */,
  {32'hbeadecd1, 32'h00000000} /* (27, 11, 7) {real, imag} */,
  {32'hbf2c2dd0, 32'h00000000} /* (27, 11, 6) {real, imag} */,
  {32'hbecb36ab, 32'h00000000} /* (27, 11, 5) {real, imag} */,
  {32'hbdeafbda, 32'h00000000} /* (27, 11, 4) {real, imag} */,
  {32'hbf230fcd, 32'h00000000} /* (27, 11, 3) {real, imag} */,
  {32'hbf24f811, 32'h00000000} /* (27, 11, 2) {real, imag} */,
  {32'hbef95d15, 32'h00000000} /* (27, 11, 1) {real, imag} */,
  {32'hbe3dbb25, 32'h00000000} /* (27, 11, 0) {real, imag} */,
  {32'h3eb5537d, 32'h00000000} /* (27, 10, 31) {real, imag} */,
  {32'h3edeb8c5, 32'h00000000} /* (27, 10, 30) {real, imag} */,
  {32'h3de06dac, 32'h00000000} /* (27, 10, 29) {real, imag} */,
  {32'h3de55e34, 32'h00000000} /* (27, 10, 28) {real, imag} */,
  {32'h3e9d2744, 32'h00000000} /* (27, 10, 27) {real, imag} */,
  {32'h3ebd751b, 32'h00000000} /* (27, 10, 26) {real, imag} */,
  {32'h3e1eec2d, 32'h00000000} /* (27, 10, 25) {real, imag} */,
  {32'h3ed49e16, 32'h00000000} /* (27, 10, 24) {real, imag} */,
  {32'h3f361498, 32'h00000000} /* (27, 10, 23) {real, imag} */,
  {32'h3f67e41f, 32'h00000000} /* (27, 10, 22) {real, imag} */,
  {32'h3ef617d4, 32'h00000000} /* (27, 10, 21) {real, imag} */,
  {32'hbe75f92a, 32'h00000000} /* (27, 10, 20) {real, imag} */,
  {32'hbf5fc926, 32'h00000000} /* (27, 10, 19) {real, imag} */,
  {32'hbec9f385, 32'h00000000} /* (27, 10, 18) {real, imag} */,
  {32'hbed66255, 32'h00000000} /* (27, 10, 17) {real, imag} */,
  {32'hbe8b4d2f, 32'h00000000} /* (27, 10, 16) {real, imag} */,
  {32'h3e29ad32, 32'h00000000} /* (27, 10, 15) {real, imag} */,
  {32'h3e450411, 32'h00000000} /* (27, 10, 14) {real, imag} */,
  {32'hbcc03f8d, 32'h00000000} /* (27, 10, 13) {real, imag} */,
  {32'hbf03d933, 32'h00000000} /* (27, 10, 12) {real, imag} */,
  {32'hbf89fdb6, 32'h00000000} /* (27, 10, 11) {real, imag} */,
  {32'hbe979687, 32'h00000000} /* (27, 10, 10) {real, imag} */,
  {32'h3ea0ab33, 32'h00000000} /* (27, 10, 9) {real, imag} */,
  {32'h3f307828, 32'h00000000} /* (27, 10, 8) {real, imag} */,
  {32'h3f8c2760, 32'h00000000} /* (27, 10, 7) {real, imag} */,
  {32'h3f898f0b, 32'h00000000} /* (27, 10, 6) {real, imag} */,
  {32'h3f1df223, 32'h00000000} /* (27, 10, 5) {real, imag} */,
  {32'h3f11ac0e, 32'h00000000} /* (27, 10, 4) {real, imag} */,
  {32'hbd3cd53f, 32'h00000000} /* (27, 10, 3) {real, imag} */,
  {32'h3c072573, 32'h00000000} /* (27, 10, 2) {real, imag} */,
  {32'h3f0f2cb9, 32'h00000000} /* (27, 10, 1) {real, imag} */,
  {32'h3ef38eb1, 32'h00000000} /* (27, 10, 0) {real, imag} */,
  {32'h3f4a6453, 32'h00000000} /* (27, 9, 31) {real, imag} */,
  {32'h3f6dca0f, 32'h00000000} /* (27, 9, 30) {real, imag} */,
  {32'h3f7ee6fc, 32'h00000000} /* (27, 9, 29) {real, imag} */,
  {32'h3f5be04d, 32'h00000000} /* (27, 9, 28) {real, imag} */,
  {32'h3f075b8e, 32'h00000000} /* (27, 9, 27) {real, imag} */,
  {32'h3f0bda92, 32'h00000000} /* (27, 9, 26) {real, imag} */,
  {32'h3f32a3a1, 32'h00000000} /* (27, 9, 25) {real, imag} */,
  {32'h3f5ebc32, 32'h00000000} /* (27, 9, 24) {real, imag} */,
  {32'h3f5366e1, 32'h00000000} /* (27, 9, 23) {real, imag} */,
  {32'h3fa9029d, 32'h00000000} /* (27, 9, 22) {real, imag} */,
  {32'h3f47d717, 32'h00000000} /* (27, 9, 21) {real, imag} */,
  {32'hbf0af1d7, 32'h00000000} /* (27, 9, 20) {real, imag} */,
  {32'hbfa6229b, 32'h00000000} /* (27, 9, 19) {real, imag} */,
  {32'hbf5b2236, 32'h00000000} /* (27, 9, 18) {real, imag} */,
  {32'hbf747523, 32'h00000000} /* (27, 9, 17) {real, imag} */,
  {32'hbf6b8dc9, 32'h00000000} /* (27, 9, 16) {real, imag} */,
  {32'hbf571450, 32'h00000000} /* (27, 9, 15) {real, imag} */,
  {32'hbf0fb4ab, 32'h00000000} /* (27, 9, 14) {real, imag} */,
  {32'hbf692285, 32'h00000000} /* (27, 9, 13) {real, imag} */,
  {32'hbf3a9ded, 32'h00000000} /* (27, 9, 12) {real, imag} */,
  {32'hbf03bba9, 32'h00000000} /* (27, 9, 11) {real, imag} */,
  {32'h3f084a0d, 32'h00000000} /* (27, 9, 10) {real, imag} */,
  {32'h3f9dee22, 32'h00000000} /* (27, 9, 9) {real, imag} */,
  {32'h3f8151b8, 32'h00000000} /* (27, 9, 8) {real, imag} */,
  {32'h3f52f3a3, 32'h00000000} /* (27, 9, 7) {real, imag} */,
  {32'h3f657678, 32'h00000000} /* (27, 9, 6) {real, imag} */,
  {32'h3f06c1f1, 32'h00000000} /* (27, 9, 5) {real, imag} */,
  {32'h3f12b42e, 32'h00000000} /* (27, 9, 4) {real, imag} */,
  {32'h3ef5d724, 32'h00000000} /* (27, 9, 3) {real, imag} */,
  {32'h3ec35a71, 32'h00000000} /* (27, 9, 2) {real, imag} */,
  {32'h3f50dea9, 32'h00000000} /* (27, 9, 1) {real, imag} */,
  {32'h3f2a07b2, 32'h00000000} /* (27, 9, 0) {real, imag} */,
  {32'h3ef2ea6d, 32'h00000000} /* (27, 8, 31) {real, imag} */,
  {32'h3f26be35, 32'h00000000} /* (27, 8, 30) {real, imag} */,
  {32'h3f9bf7df, 32'h00000000} /* (27, 8, 29) {real, imag} */,
  {32'h3f3d14d3, 32'h00000000} /* (27, 8, 28) {real, imag} */,
  {32'h3f2f6a76, 32'h00000000} /* (27, 8, 27) {real, imag} */,
  {32'h3f3eb827, 32'h00000000} /* (27, 8, 26) {real, imag} */,
  {32'h3f38d65f, 32'h00000000} /* (27, 8, 25) {real, imag} */,
  {32'h3f183e93, 32'h00000000} /* (27, 8, 24) {real, imag} */,
  {32'h3f16d365, 32'h00000000} /* (27, 8, 23) {real, imag} */,
  {32'h3fced8f0, 32'h00000000} /* (27, 8, 22) {real, imag} */,
  {32'h3f36dddb, 32'h00000000} /* (27, 8, 21) {real, imag} */,
  {32'hbeaf2ffc, 32'h00000000} /* (27, 8, 20) {real, imag} */,
  {32'hbf724e75, 32'h00000000} /* (27, 8, 19) {real, imag} */,
  {32'hbf9e3b54, 32'h00000000} /* (27, 8, 18) {real, imag} */,
  {32'hbf7f85ed, 32'h00000000} /* (27, 8, 17) {real, imag} */,
  {32'hbf9b2334, 32'h00000000} /* (27, 8, 16) {real, imag} */,
  {32'hbfaf0f9c, 32'h00000000} /* (27, 8, 15) {real, imag} */,
  {32'hbf6ef27f, 32'h00000000} /* (27, 8, 14) {real, imag} */,
  {32'hbf69fb27, 32'h00000000} /* (27, 8, 13) {real, imag} */,
  {32'hbf58bedf, 32'h00000000} /* (27, 8, 12) {real, imag} */,
  {32'hbf8f3bb9, 32'h00000000} /* (27, 8, 11) {real, imag} */,
  {32'h3bfba3c2, 32'h00000000} /* (27, 8, 10) {real, imag} */,
  {32'h3f7ce0f2, 32'h00000000} /* (27, 8, 9) {real, imag} */,
  {32'h3f5bf1c6, 32'h00000000} /* (27, 8, 8) {real, imag} */,
  {32'h3f68f057, 32'h00000000} /* (27, 8, 7) {real, imag} */,
  {32'h3f7946cf, 32'h00000000} /* (27, 8, 6) {real, imag} */,
  {32'h3f36eecf, 32'h00000000} /* (27, 8, 5) {real, imag} */,
  {32'h3f257825, 32'h00000000} /* (27, 8, 4) {real, imag} */,
  {32'h3f1e2582, 32'h00000000} /* (27, 8, 3) {real, imag} */,
  {32'h3ed88ee8, 32'h00000000} /* (27, 8, 2) {real, imag} */,
  {32'h3f1a4d5f, 32'h00000000} /* (27, 8, 1) {real, imag} */,
  {32'h3ee38204, 32'h00000000} /* (27, 8, 0) {real, imag} */,
  {32'h3ec1edf2, 32'h00000000} /* (27, 7, 31) {real, imag} */,
  {32'h3f005f7f, 32'h00000000} /* (27, 7, 30) {real, imag} */,
  {32'h3ed2b630, 32'h00000000} /* (27, 7, 29) {real, imag} */,
  {32'h3f01737b, 32'h00000000} /* (27, 7, 28) {real, imag} */,
  {32'h3f639c43, 32'h00000000} /* (27, 7, 27) {real, imag} */,
  {32'h3f549283, 32'h00000000} /* (27, 7, 26) {real, imag} */,
  {32'h3f901495, 32'h00000000} /* (27, 7, 25) {real, imag} */,
  {32'h3f59731d, 32'h00000000} /* (27, 7, 24) {real, imag} */,
  {32'h3f559330, 32'h00000000} /* (27, 7, 23) {real, imag} */,
  {32'h3f868a96, 32'h00000000} /* (27, 7, 22) {real, imag} */,
  {32'h3f13cae0, 32'h00000000} /* (27, 7, 21) {real, imag} */,
  {32'hbec21479, 32'h00000000} /* (27, 7, 20) {real, imag} */,
  {32'hbf5cca02, 32'h00000000} /* (27, 7, 19) {real, imag} */,
  {32'hbf6c4707, 32'h00000000} /* (27, 7, 18) {real, imag} */,
  {32'hbf99ddf8, 32'h00000000} /* (27, 7, 17) {real, imag} */,
  {32'hbf630748, 32'h00000000} /* (27, 7, 16) {real, imag} */,
  {32'hbf5ce114, 32'h00000000} /* (27, 7, 15) {real, imag} */,
  {32'hbf655ab8, 32'h00000000} /* (27, 7, 14) {real, imag} */,
  {32'hbf5ae064, 32'h00000000} /* (27, 7, 13) {real, imag} */,
  {32'hbec3f3c7, 32'h00000000} /* (27, 7, 12) {real, imag} */,
  {32'hbf3e0631, 32'h00000000} /* (27, 7, 11) {real, imag} */,
  {32'hbe91492e, 32'h00000000} /* (27, 7, 10) {real, imag} */,
  {32'h3f1a0256, 32'h00000000} /* (27, 7, 9) {real, imag} */,
  {32'h3f36f980, 32'h00000000} /* (27, 7, 8) {real, imag} */,
  {32'h3f611a6c, 32'h00000000} /* (27, 7, 7) {real, imag} */,
  {32'h3f352da9, 32'h00000000} /* (27, 7, 6) {real, imag} */,
  {32'h3fa0d0a4, 32'h00000000} /* (27, 7, 5) {real, imag} */,
  {32'h3f877f5d, 32'h00000000} /* (27, 7, 4) {real, imag} */,
  {32'h3f15c750, 32'h00000000} /* (27, 7, 3) {real, imag} */,
  {32'h3f493e0e, 32'h00000000} /* (27, 7, 2) {real, imag} */,
  {32'h3f4dc056, 32'h00000000} /* (27, 7, 1) {real, imag} */,
  {32'h3ee928ee, 32'h00000000} /* (27, 7, 0) {real, imag} */,
  {32'h3eb59586, 32'h00000000} /* (27, 6, 31) {real, imag} */,
  {32'h3ee8988f, 32'h00000000} /* (27, 6, 30) {real, imag} */,
  {32'h3f0cb8b0, 32'h00000000} /* (27, 6, 29) {real, imag} */,
  {32'h3f11c0ab, 32'h00000000} /* (27, 6, 28) {real, imag} */,
  {32'h3f898b38, 32'h00000000} /* (27, 6, 27) {real, imag} */,
  {32'h3fa7f56d, 32'h00000000} /* (27, 6, 26) {real, imag} */,
  {32'h3fc16004, 32'h00000000} /* (27, 6, 25) {real, imag} */,
  {32'h3f2a94b2, 32'h00000000} /* (27, 6, 24) {real, imag} */,
  {32'h3f0b8806, 32'h00000000} /* (27, 6, 23) {real, imag} */,
  {32'h3f881ebe, 32'h00000000} /* (27, 6, 22) {real, imag} */,
  {32'h3f875ca3, 32'h00000000} /* (27, 6, 21) {real, imag} */,
  {32'hbe18c3c0, 32'h00000000} /* (27, 6, 20) {real, imag} */,
  {32'hbf4a629f, 32'h00000000} /* (27, 6, 19) {real, imag} */,
  {32'hbf5fec32, 32'h00000000} /* (27, 6, 18) {real, imag} */,
  {32'hbf01009f, 32'h00000000} /* (27, 6, 17) {real, imag} */,
  {32'hbe5cb905, 32'h00000000} /* (27, 6, 16) {real, imag} */,
  {32'hbee9c9b8, 32'h00000000} /* (27, 6, 15) {real, imag} */,
  {32'hbf83294f, 32'h00000000} /* (27, 6, 14) {real, imag} */,
  {32'hbfb45c6a, 32'h00000000} /* (27, 6, 13) {real, imag} */,
  {32'hbf00988b, 32'h00000000} /* (27, 6, 12) {real, imag} */,
  {32'hbeb010bf, 32'h00000000} /* (27, 6, 11) {real, imag} */,
  {32'h3f1d5655, 32'h00000000} /* (27, 6, 10) {real, imag} */,
  {32'h3f9b4c95, 32'h00000000} /* (27, 6, 9) {real, imag} */,
  {32'h3f3462ed, 32'h00000000} /* (27, 6, 8) {real, imag} */,
  {32'h3f58035b, 32'h00000000} /* (27, 6, 7) {real, imag} */,
  {32'h3f42f2c5, 32'h00000000} /* (27, 6, 6) {real, imag} */,
  {32'h3fa21a66, 32'h00000000} /* (27, 6, 5) {real, imag} */,
  {32'h3f9366c3, 32'h00000000} /* (27, 6, 4) {real, imag} */,
  {32'h3f061a8f, 32'h00000000} /* (27, 6, 3) {real, imag} */,
  {32'h3f44988d, 32'h00000000} /* (27, 6, 2) {real, imag} */,
  {32'h3f934fae, 32'h00000000} /* (27, 6, 1) {real, imag} */,
  {32'h3f12d809, 32'h00000000} /* (27, 6, 0) {real, imag} */,
  {32'h3e95986b, 32'h00000000} /* (27, 5, 31) {real, imag} */,
  {32'h3f326453, 32'h00000000} /* (27, 5, 30) {real, imag} */,
  {32'h3f7475b1, 32'h00000000} /* (27, 5, 29) {real, imag} */,
  {32'h3f757a7e, 32'h00000000} /* (27, 5, 28) {real, imag} */,
  {32'h3f75d85f, 32'h00000000} /* (27, 5, 27) {real, imag} */,
  {32'h3f906057, 32'h00000000} /* (27, 5, 26) {real, imag} */,
  {32'h3fb7b24f, 32'h00000000} /* (27, 5, 25) {real, imag} */,
  {32'h3f69f12f, 32'h00000000} /* (27, 5, 24) {real, imag} */,
  {32'h3f0c8e21, 32'h00000000} /* (27, 5, 23) {real, imag} */,
  {32'h3f837dc4, 32'h00000000} /* (27, 5, 22) {real, imag} */,
  {32'h3f98d62f, 32'h00000000} /* (27, 5, 21) {real, imag} */,
  {32'h3f4c6fe5, 32'h00000000} /* (27, 5, 20) {real, imag} */,
  {32'h3dd292ed, 32'h00000000} /* (27, 5, 19) {real, imag} */,
  {32'hbdde8f0a, 32'h00000000} /* (27, 5, 18) {real, imag} */,
  {32'h3e4563e2, 32'h00000000} /* (27, 5, 17) {real, imag} */,
  {32'hbc548394, 32'h00000000} /* (27, 5, 16) {real, imag} */,
  {32'hbec2544c, 32'h00000000} /* (27, 5, 15) {real, imag} */,
  {32'hbf8b2193, 32'h00000000} /* (27, 5, 14) {real, imag} */,
  {32'hbf8cc2d7, 32'h00000000} /* (27, 5, 13) {real, imag} */,
  {32'hbeec9836, 32'h00000000} /* (27, 5, 12) {real, imag} */,
  {32'hbf17c24f, 32'h00000000} /* (27, 5, 11) {real, imag} */,
  {32'h3e001b68, 32'h00000000} /* (27, 5, 10) {real, imag} */,
  {32'h3f06f545, 32'h00000000} /* (27, 5, 9) {real, imag} */,
  {32'hbdf6f375, 32'h00000000} /* (27, 5, 8) {real, imag} */,
  {32'hbdba554d, 32'h00000000} /* (27, 5, 7) {real, imag} */,
  {32'h3d0ec17c, 32'h00000000} /* (27, 5, 6) {real, imag} */,
  {32'h3f36e34a, 32'h00000000} /* (27, 5, 5) {real, imag} */,
  {32'h3f1915b1, 32'h00000000} /* (27, 5, 4) {real, imag} */,
  {32'h3f27a064, 32'h00000000} /* (27, 5, 3) {real, imag} */,
  {32'h3f507c7d, 32'h00000000} /* (27, 5, 2) {real, imag} */,
  {32'h3f665eb0, 32'h00000000} /* (27, 5, 1) {real, imag} */,
  {32'h3f0fbc47, 32'h00000000} /* (27, 5, 0) {real, imag} */,
  {32'h3e6434d4, 32'h00000000} /* (27, 4, 31) {real, imag} */,
  {32'h3f23a797, 32'h00000000} /* (27, 4, 30) {real, imag} */,
  {32'h3f3f55ab, 32'h00000000} /* (27, 4, 29) {real, imag} */,
  {32'h3f80f377, 32'h00000000} /* (27, 4, 28) {real, imag} */,
  {32'h3f0fafc9, 32'h00000000} /* (27, 4, 27) {real, imag} */,
  {32'h3bd70be8, 32'h00000000} /* (27, 4, 26) {real, imag} */,
  {32'h3d7c82e3, 32'h00000000} /* (27, 4, 25) {real, imag} */,
  {32'h3f140050, 32'h00000000} /* (27, 4, 24) {real, imag} */,
  {32'h3f59f0ca, 32'h00000000} /* (27, 4, 23) {real, imag} */,
  {32'h3f78645c, 32'h00000000} /* (27, 4, 22) {real, imag} */,
  {32'h3f7f43d6, 32'h00000000} /* (27, 4, 21) {real, imag} */,
  {32'h3f802953, 32'h00000000} /* (27, 4, 20) {real, imag} */,
  {32'h3eead2be, 32'h00000000} /* (27, 4, 19) {real, imag} */,
  {32'h3f27bec9, 32'h00000000} /* (27, 4, 18) {real, imag} */,
  {32'h3f871440, 32'h00000000} /* (27, 4, 17) {real, imag} */,
  {32'h3f5aaeb6, 32'h00000000} /* (27, 4, 16) {real, imag} */,
  {32'hbdcd0d5e, 32'h00000000} /* (27, 4, 15) {real, imag} */,
  {32'hbf2320ad, 32'h00000000} /* (27, 4, 14) {real, imag} */,
  {32'hbf5f09b2, 32'h00000000} /* (27, 4, 13) {real, imag} */,
  {32'hbef4ae3d, 32'h00000000} /* (27, 4, 12) {real, imag} */,
  {32'hbf299705, 32'h00000000} /* (27, 4, 11) {real, imag} */,
  {32'hbf2366ff, 32'h00000000} /* (27, 4, 10) {real, imag} */,
  {32'hbecf5e7f, 32'h00000000} /* (27, 4, 9) {real, imag} */,
  {32'hbf34b45a, 32'h00000000} /* (27, 4, 8) {real, imag} */,
  {32'hbf099ce9, 32'h00000000} /* (27, 4, 7) {real, imag} */,
  {32'hbeaf3ba5, 32'h00000000} /* (27, 4, 6) {real, imag} */,
  {32'h3fa06cf5, 32'h00000000} /* (27, 4, 5) {real, imag} */,
  {32'h3f99c9c4, 32'h00000000} /* (27, 4, 4) {real, imag} */,
  {32'h3f883791, 32'h00000000} /* (27, 4, 3) {real, imag} */,
  {32'h3f7fe022, 32'h00000000} /* (27, 4, 2) {real, imag} */,
  {32'h3eff4ede, 32'h00000000} /* (27, 4, 1) {real, imag} */,
  {32'h3e97ff31, 32'h00000000} /* (27, 4, 0) {real, imag} */,
  {32'h3e883daf, 32'h00000000} /* (27, 3, 31) {real, imag} */,
  {32'h3f9aeeea, 32'h00000000} /* (27, 3, 30) {real, imag} */,
  {32'h3f915b37, 32'h00000000} /* (27, 3, 29) {real, imag} */,
  {32'h3fb99ca5, 32'h00000000} /* (27, 3, 28) {real, imag} */,
  {32'h3f967bc5, 32'h00000000} /* (27, 3, 27) {real, imag} */,
  {32'h3ef7e772, 32'h00000000} /* (27, 3, 26) {real, imag} */,
  {32'h3eaf1fa4, 32'h00000000} /* (27, 3, 25) {real, imag} */,
  {32'h3f175e50, 32'h00000000} /* (27, 3, 24) {real, imag} */,
  {32'h3f336144, 32'h00000000} /* (27, 3, 23) {real, imag} */,
  {32'h3f4396f9, 32'h00000000} /* (27, 3, 22) {real, imag} */,
  {32'h3f8b77e6, 32'h00000000} /* (27, 3, 21) {real, imag} */,
  {32'h3f9aef97, 32'h00000000} /* (27, 3, 20) {real, imag} */,
  {32'h3f946e88, 32'h00000000} /* (27, 3, 19) {real, imag} */,
  {32'h3f731a84, 32'h00000000} /* (27, 3, 18) {real, imag} */,
  {32'h3f87160d, 32'h00000000} /* (27, 3, 17) {real, imag} */,
  {32'h3f5c870f, 32'h00000000} /* (27, 3, 16) {real, imag} */,
  {32'hbde7e546, 32'h00000000} /* (27, 3, 15) {real, imag} */,
  {32'hbdcdc9f5, 32'h00000000} /* (27, 3, 14) {real, imag} */,
  {32'hbf6faa3b, 32'h00000000} /* (27, 3, 13) {real, imag} */,
  {32'hbf44cfb9, 32'h00000000} /* (27, 3, 12) {real, imag} */,
  {32'hbf16474d, 32'h00000000} /* (27, 3, 11) {real, imag} */,
  {32'hbf46f803, 32'h00000000} /* (27, 3, 10) {real, imag} */,
  {32'hbf23ee25, 32'h00000000} /* (27, 3, 9) {real, imag} */,
  {32'hbedd3713, 32'h00000000} /* (27, 3, 8) {real, imag} */,
  {32'hbe99ddb4, 32'h00000000} /* (27, 3, 7) {real, imag} */,
  {32'hbf0502a6, 32'h00000000} /* (27, 3, 6) {real, imag} */,
  {32'h3f1c2c15, 32'h00000000} /* (27, 3, 5) {real, imag} */,
  {32'h3f3ac9c4, 32'h00000000} /* (27, 3, 4) {real, imag} */,
  {32'h3f708f17, 32'h00000000} /* (27, 3, 3) {real, imag} */,
  {32'h3fb2fee8, 32'h00000000} /* (27, 3, 2) {real, imag} */,
  {32'h3f7f9567, 32'h00000000} /* (27, 3, 1) {real, imag} */,
  {32'h3f04b02f, 32'h00000000} /* (27, 3, 0) {real, imag} */,
  {32'h3ed48979, 32'h00000000} /* (27, 2, 31) {real, imag} */,
  {32'h3fa4c6dc, 32'h00000000} /* (27, 2, 30) {real, imag} */,
  {32'h3f6ce9ad, 32'h00000000} /* (27, 2, 29) {real, imag} */,
  {32'h3f73ffa2, 32'h00000000} /* (27, 2, 28) {real, imag} */,
  {32'h3f91a3e9, 32'h00000000} /* (27, 2, 27) {real, imag} */,
  {32'h3f3ecc9c, 32'h00000000} /* (27, 2, 26) {real, imag} */,
  {32'h3f34c9ca, 32'h00000000} /* (27, 2, 25) {real, imag} */,
  {32'h3f919d8c, 32'h00000000} /* (27, 2, 24) {real, imag} */,
  {32'h3f5d84f9, 32'h00000000} /* (27, 2, 23) {real, imag} */,
  {32'h3f78dbb4, 32'h00000000} /* (27, 2, 22) {real, imag} */,
  {32'h3fc6669c, 32'h00000000} /* (27, 2, 21) {real, imag} */,
  {32'h3fb2c099, 32'h00000000} /* (27, 2, 20) {real, imag} */,
  {32'h3fb7d1b2, 32'h00000000} /* (27, 2, 19) {real, imag} */,
  {32'h3f206820, 32'h00000000} /* (27, 2, 18) {real, imag} */,
  {32'h3f976318, 32'h00000000} /* (27, 2, 17) {real, imag} */,
  {32'h3f855f4f, 32'h00000000} /* (27, 2, 16) {real, imag} */,
  {32'hbf145ee8, 32'h00000000} /* (27, 2, 15) {real, imag} */,
  {32'hbee9599a, 32'h00000000} /* (27, 2, 14) {real, imag} */,
  {32'hbf24aded, 32'h00000000} /* (27, 2, 13) {real, imag} */,
  {32'hbf6b8425, 32'h00000000} /* (27, 2, 12) {real, imag} */,
  {32'hbf807fa5, 32'h00000000} /* (27, 2, 11) {real, imag} */,
  {32'hbfa13e22, 32'h00000000} /* (27, 2, 10) {real, imag} */,
  {32'hbfa7ba07, 32'h00000000} /* (27, 2, 9) {real, imag} */,
  {32'hbf7b54da, 32'h00000000} /* (27, 2, 8) {real, imag} */,
  {32'hbed02ac4, 32'h00000000} /* (27, 2, 7) {real, imag} */,
  {32'hbf46c30c, 32'h00000000} /* (27, 2, 6) {real, imag} */,
  {32'hbe136f91, 32'h00000000} /* (27, 2, 5) {real, imag} */,
  {32'h3ec41bdf, 32'h00000000} /* (27, 2, 4) {real, imag} */,
  {32'h3f660f30, 32'h00000000} /* (27, 2, 3) {real, imag} */,
  {32'h3fb795c4, 32'h00000000} /* (27, 2, 2) {real, imag} */,
  {32'h3fac909a, 32'h00000000} /* (27, 2, 1) {real, imag} */,
  {32'h3f39a421, 32'h00000000} /* (27, 2, 0) {real, imag} */,
  {32'h3f62e751, 32'h00000000} /* (27, 1, 31) {real, imag} */,
  {32'h3fb9480e, 32'h00000000} /* (27, 1, 30) {real, imag} */,
  {32'h3f78b562, 32'h00000000} /* (27, 1, 29) {real, imag} */,
  {32'h3f0d6da4, 32'h00000000} /* (27, 1, 28) {real, imag} */,
  {32'h3f7f2971, 32'h00000000} /* (27, 1, 27) {real, imag} */,
  {32'h3f0428ea, 32'h00000000} /* (27, 1, 26) {real, imag} */,
  {32'h3f6ef418, 32'h00000000} /* (27, 1, 25) {real, imag} */,
  {32'h3f842aae, 32'h00000000} /* (27, 1, 24) {real, imag} */,
  {32'h3f900b24, 32'h00000000} /* (27, 1, 23) {real, imag} */,
  {32'h3fc1094e, 32'h00000000} /* (27, 1, 22) {real, imag} */,
  {32'h3fa2685e, 32'h00000000} /* (27, 1, 21) {real, imag} */,
  {32'h3f6688a5, 32'h00000000} /* (27, 1, 20) {real, imag} */,
  {32'h3fbe9af0, 32'h00000000} /* (27, 1, 19) {real, imag} */,
  {32'h3fb3bd02, 32'h00000000} /* (27, 1, 18) {real, imag} */,
  {32'h3fc1f590, 32'h00000000} /* (27, 1, 17) {real, imag} */,
  {32'h3f94a2ed, 32'h00000000} /* (27, 1, 16) {real, imag} */,
  {32'hbee087a7, 32'h00000000} /* (27, 1, 15) {real, imag} */,
  {32'hbf2e1c72, 32'h00000000} /* (27, 1, 14) {real, imag} */,
  {32'hbf354c68, 32'h00000000} /* (27, 1, 13) {real, imag} */,
  {32'hbf91255a, 32'h00000000} /* (27, 1, 12) {real, imag} */,
  {32'hbf82d6d7, 32'h00000000} /* (27, 1, 11) {real, imag} */,
  {32'hbf9575e1, 32'h00000000} /* (27, 1, 10) {real, imag} */,
  {32'hbfccb261, 32'h00000000} /* (27, 1, 9) {real, imag} */,
  {32'hbfbec805, 32'h00000000} /* (27, 1, 8) {real, imag} */,
  {32'hbf5a1c65, 32'h00000000} /* (27, 1, 7) {real, imag} */,
  {32'hbf502f6a, 32'h00000000} /* (27, 1, 6) {real, imag} */,
  {32'hbde80a57, 32'h00000000} /* (27, 1, 5) {real, imag} */,
  {32'h3f124ae8, 32'h00000000} /* (27, 1, 4) {real, imag} */,
  {32'h3f51eb18, 32'h00000000} /* (27, 1, 3) {real, imag} */,
  {32'h3f95d0a6, 32'h00000000} /* (27, 1, 2) {real, imag} */,
  {32'h3fa36e76, 32'h00000000} /* (27, 1, 1) {real, imag} */,
  {32'h3f77917a, 32'h00000000} /* (27, 1, 0) {real, imag} */,
  {32'h3e94ff3c, 32'h00000000} /* (27, 0, 31) {real, imag} */,
  {32'h3f1b752c, 32'h00000000} /* (27, 0, 30) {real, imag} */,
  {32'h3f010e09, 32'h00000000} /* (27, 0, 29) {real, imag} */,
  {32'h3e869959, 32'h00000000} /* (27, 0, 28) {real, imag} */,
  {32'h3ebb1a99, 32'h00000000} /* (27, 0, 27) {real, imag} */,
  {32'h3e64abdc, 32'h00000000} /* (27, 0, 26) {real, imag} */,
  {32'h3f00b2dd, 32'h00000000} /* (27, 0, 25) {real, imag} */,
  {32'h3eea8008, 32'h00000000} /* (27, 0, 24) {real, imag} */,
  {32'h3f1cde71, 32'h00000000} /* (27, 0, 23) {real, imag} */,
  {32'h3f6860dd, 32'h00000000} /* (27, 0, 22) {real, imag} */,
  {32'h3f0957e1, 32'h00000000} /* (27, 0, 21) {real, imag} */,
  {32'h3ec7a7db, 32'h00000000} /* (27, 0, 20) {real, imag} */,
  {32'h3f6bcc9a, 32'h00000000} /* (27, 0, 19) {real, imag} */,
  {32'h3f97d35e, 32'h00000000} /* (27, 0, 18) {real, imag} */,
  {32'h3f30685d, 32'h00000000} /* (27, 0, 17) {real, imag} */,
  {32'h3e36722c, 32'h00000000} /* (27, 0, 16) {real, imag} */,
  {32'hbe929c78, 32'h00000000} /* (27, 0, 15) {real, imag} */,
  {32'hbe8a5850, 32'h00000000} /* (27, 0, 14) {real, imag} */,
  {32'hbee8bda7, 32'h00000000} /* (27, 0, 13) {real, imag} */,
  {32'hbf276421, 32'h00000000} /* (27, 0, 12) {real, imag} */,
  {32'hbed496b4, 32'h00000000} /* (27, 0, 11) {real, imag} */,
  {32'hbe4d0ad5, 32'h00000000} /* (27, 0, 10) {real, imag} */,
  {32'hbe1aa299, 32'h00000000} /* (27, 0, 9) {real, imag} */,
  {32'hbef3a662, 32'h00000000} /* (27, 0, 8) {real, imag} */,
  {32'hbf2e71ca, 32'h00000000} /* (27, 0, 7) {real, imag} */,
  {32'hbf18a373, 32'h00000000} /* (27, 0, 6) {real, imag} */,
  {32'hbc6c7ec9, 32'h00000000} /* (27, 0, 5) {real, imag} */,
  {32'h3ecbf7f8, 32'h00000000} /* (27, 0, 4) {real, imag} */,
  {32'h3ee05a99, 32'h00000000} /* (27, 0, 3) {real, imag} */,
  {32'h3eee3fc7, 32'h00000000} /* (27, 0, 2) {real, imag} */,
  {32'h3ec92af5, 32'h00000000} /* (27, 0, 1) {real, imag} */,
  {32'h3e99bcf0, 32'h00000000} /* (27, 0, 0) {real, imag} */,
  {32'h3cd49734, 32'h00000000} /* (26, 31, 31) {real, imag} */,
  {32'hbe50e0f0, 32'h00000000} /* (26, 31, 30) {real, imag} */,
  {32'h3bd5ef94, 32'h00000000} /* (26, 31, 29) {real, imag} */,
  {32'h3e557f4d, 32'h00000000} /* (26, 31, 28) {real, imag} */,
  {32'h3f1d4f73, 32'h00000000} /* (26, 31, 27) {real, imag} */,
  {32'h3e9c3eac, 32'h00000000} /* (26, 31, 26) {real, imag} */,
  {32'h3e482204, 32'h00000000} /* (26, 31, 25) {real, imag} */,
  {32'h3df67802, 32'h00000000} /* (26, 31, 24) {real, imag} */,
  {32'hbe4304cc, 32'h00000000} /* (26, 31, 23) {real, imag} */,
  {32'hbe827d84, 32'h00000000} /* (26, 31, 22) {real, imag} */,
  {32'hbec3b2d9, 32'h00000000} /* (26, 31, 21) {real, imag} */,
  {32'hbf1d73ae, 32'h00000000} /* (26, 31, 20) {real, imag} */,
  {32'hbd1a28be, 32'h00000000} /* (26, 31, 19) {real, imag} */,
  {32'h3e92f71c, 32'h00000000} /* (26, 31, 18) {real, imag} */,
  {32'h3d4fbb7c, 32'h00000000} /* (26, 31, 17) {real, imag} */,
  {32'hbe0478f7, 32'h00000000} /* (26, 31, 16) {real, imag} */,
  {32'h3c8fe442, 32'h00000000} /* (26, 31, 15) {real, imag} */,
  {32'hbea9adf2, 32'h00000000} /* (26, 31, 14) {real, imag} */,
  {32'hbe5a347c, 32'h00000000} /* (26, 31, 13) {real, imag} */,
  {32'h3e0bb270, 32'h00000000} /* (26, 31, 12) {real, imag} */,
  {32'hbca280c3, 32'h00000000} /* (26, 31, 11) {real, imag} */,
  {32'hbca71768, 32'h00000000} /* (26, 31, 10) {real, imag} */,
  {32'hbe479f21, 32'h00000000} /* (26, 31, 9) {real, imag} */,
  {32'hbe5864a7, 32'h00000000} /* (26, 31, 8) {real, imag} */,
  {32'hbda94d57, 32'h00000000} /* (26, 31, 7) {real, imag} */,
  {32'h3e82b4c7, 32'h00000000} /* (26, 31, 6) {real, imag} */,
  {32'h3ed79694, 32'h00000000} /* (26, 31, 5) {real, imag} */,
  {32'h3cffb758, 32'h00000000} /* (26, 31, 4) {real, imag} */,
  {32'h3dc1c881, 32'h00000000} /* (26, 31, 3) {real, imag} */,
  {32'h3eeac695, 32'h00000000} /* (26, 31, 2) {real, imag} */,
  {32'h3ea9ce79, 32'h00000000} /* (26, 31, 1) {real, imag} */,
  {32'h3f0c31ff, 32'h00000000} /* (26, 31, 0) {real, imag} */,
  {32'h3ec4923d, 32'h00000000} /* (26, 30, 31) {real, imag} */,
  {32'h3e99021d, 32'h00000000} /* (26, 30, 30) {real, imag} */,
  {32'h3e0be9a2, 32'h00000000} /* (26, 30, 29) {real, imag} */,
  {32'h3eeb004f, 32'h00000000} /* (26, 30, 28) {real, imag} */,
  {32'h3f789f7f, 32'h00000000} /* (26, 30, 27) {real, imag} */,
  {32'h3e7731df, 32'h00000000} /* (26, 30, 26) {real, imag} */,
  {32'h3def15ea, 32'h00000000} /* (26, 30, 25) {real, imag} */,
  {32'h3de2f13a, 32'h00000000} /* (26, 30, 24) {real, imag} */,
  {32'h3ea762f1, 32'h00000000} /* (26, 30, 23) {real, imag} */,
  {32'h3d91ca6a, 32'h00000000} /* (26, 30, 22) {real, imag} */,
  {32'hbd441d35, 32'h00000000} /* (26, 30, 21) {real, imag} */,
  {32'hbdaf57c2, 32'h00000000} /* (26, 30, 20) {real, imag} */,
  {32'hbcab3c9a, 32'h00000000} /* (26, 30, 19) {real, imag} */,
  {32'h3ec34873, 32'h00000000} /* (26, 30, 18) {real, imag} */,
  {32'hbe1ec9c1, 32'h00000000} /* (26, 30, 17) {real, imag} */,
  {32'hbd6745a9, 32'h00000000} /* (26, 30, 16) {real, imag} */,
  {32'h3e3fcfd8, 32'h00000000} /* (26, 30, 15) {real, imag} */,
  {32'hbe9f3b2b, 32'h00000000} /* (26, 30, 14) {real, imag} */,
  {32'hbe4f9b33, 32'h00000000} /* (26, 30, 13) {real, imag} */,
  {32'hbe15a726, 32'h00000000} /* (26, 30, 12) {real, imag} */,
  {32'hbe6f5022, 32'h00000000} /* (26, 30, 11) {real, imag} */,
  {32'h3e6526a9, 32'h00000000} /* (26, 30, 10) {real, imag} */,
  {32'hbe398a67, 32'h00000000} /* (26, 30, 9) {real, imag} */,
  {32'hbf01fa99, 32'h00000000} /* (26, 30, 8) {real, imag} */,
  {32'h3d2297ef, 32'h00000000} /* (26, 30, 7) {real, imag} */,
  {32'h3f28cbd9, 32'h00000000} /* (26, 30, 6) {real, imag} */,
  {32'h3f322871, 32'h00000000} /* (26, 30, 5) {real, imag} */,
  {32'h3ef466d7, 32'h00000000} /* (26, 30, 4) {real, imag} */,
  {32'h3e744120, 32'h00000000} /* (26, 30, 3) {real, imag} */,
  {32'h3ecc655b, 32'h00000000} /* (26, 30, 2) {real, imag} */,
  {32'hbd5cac53, 32'h00000000} /* (26, 30, 1) {real, imag} */,
  {32'h3e5f6378, 32'h00000000} /* (26, 30, 0) {real, imag} */,
  {32'h3f7aa5b6, 32'h00000000} /* (26, 29, 31) {real, imag} */,
  {32'h3f44d244, 32'h00000000} /* (26, 29, 30) {real, imag} */,
  {32'hbd9c0cba, 32'h00000000} /* (26, 29, 29) {real, imag} */,
  {32'h3ef37152, 32'h00000000} /* (26, 29, 28) {real, imag} */,
  {32'h3f23b07e, 32'h00000000} /* (26, 29, 27) {real, imag} */,
  {32'hbe803a96, 32'h00000000} /* (26, 29, 26) {real, imag} */,
  {32'hbea371fc, 32'h00000000} /* (26, 29, 25) {real, imag} */,
  {32'h3e5b2860, 32'h00000000} /* (26, 29, 24) {real, imag} */,
  {32'h3eb2ee61, 32'h00000000} /* (26, 29, 23) {real, imag} */,
  {32'hbe416d9e, 32'h00000000} /* (26, 29, 22) {real, imag} */,
  {32'hbe14bc22, 32'h00000000} /* (26, 29, 21) {real, imag} */,
  {32'h3e6fa9f9, 32'h00000000} /* (26, 29, 20) {real, imag} */,
  {32'h3c9cd0e9, 32'h00000000} /* (26, 29, 19) {real, imag} */,
  {32'hbe6f5342, 32'h00000000} /* (26, 29, 18) {real, imag} */,
  {32'hbeb5c360, 32'h00000000} /* (26, 29, 17) {real, imag} */,
  {32'hbf118b7f, 32'h00000000} /* (26, 29, 16) {real, imag} */,
  {32'hbe9f1141, 32'h00000000} /* (26, 29, 15) {real, imag} */,
  {32'hbde3d331, 32'h00000000} /* (26, 29, 14) {real, imag} */,
  {32'hbebdbd9e, 32'h00000000} /* (26, 29, 13) {real, imag} */,
  {32'hbf236bb6, 32'h00000000} /* (26, 29, 12) {real, imag} */,
  {32'hbf2b1518, 32'h00000000} /* (26, 29, 11) {real, imag} */,
  {32'h3e4cd4e6, 32'h00000000} /* (26, 29, 10) {real, imag} */,
  {32'h3f1daf11, 32'h00000000} /* (26, 29, 9) {real, imag} */,
  {32'h3d444caa, 32'h00000000} /* (26, 29, 8) {real, imag} */,
  {32'hbd5b0f0e, 32'h00000000} /* (26, 29, 7) {real, imag} */,
  {32'h3f193bb8, 32'h00000000} /* (26, 29, 6) {real, imag} */,
  {32'h3f83582c, 32'h00000000} /* (26, 29, 5) {real, imag} */,
  {32'h3f3eea6e, 32'h00000000} /* (26, 29, 4) {real, imag} */,
  {32'h3e4e5cbb, 32'h00000000} /* (26, 29, 3) {real, imag} */,
  {32'h3db4d90b, 32'h00000000} /* (26, 29, 2) {real, imag} */,
  {32'hbe683de8, 32'h00000000} /* (26, 29, 1) {real, imag} */,
  {32'h3ea53840, 32'h00000000} /* (26, 29, 0) {real, imag} */,
  {32'h3f339bd0, 32'h00000000} /* (26, 28, 31) {real, imag} */,
  {32'h3ec06a4a, 32'h00000000} /* (26, 28, 30) {real, imag} */,
  {32'hbecf9d8a, 32'h00000000} /* (26, 28, 29) {real, imag} */,
  {32'h3ee39a43, 32'h00000000} /* (26, 28, 28) {real, imag} */,
  {32'h3f2b0cc7, 32'h00000000} /* (26, 28, 27) {real, imag} */,
  {32'hbeab259f, 32'h00000000} /* (26, 28, 26) {real, imag} */,
  {32'hbf28e5de, 32'h00000000} /* (26, 28, 25) {real, imag} */,
  {32'h3e938a58, 32'h00000000} /* (26, 28, 24) {real, imag} */,
  {32'h3eba869f, 32'h00000000} /* (26, 28, 23) {real, imag} */,
  {32'hbe0c39e7, 32'h00000000} /* (26, 28, 22) {real, imag} */,
  {32'hbd40913b, 32'h00000000} /* (26, 28, 21) {real, imag} */,
  {32'hbeb8896b, 32'h00000000} /* (26, 28, 20) {real, imag} */,
  {32'hbee55244, 32'h00000000} /* (26, 28, 19) {real, imag} */,
  {32'hbdb81d48, 32'h00000000} /* (26, 28, 18) {real, imag} */,
  {32'h3d80145b, 32'h00000000} /* (26, 28, 17) {real, imag} */,
  {32'hbf4badb3, 32'h00000000} /* (26, 28, 16) {real, imag} */,
  {32'hbfa4fa44, 32'h00000000} /* (26, 28, 15) {real, imag} */,
  {32'hbeaf0541, 32'h00000000} /* (26, 28, 14) {real, imag} */,
  {32'hbf173e09, 32'h00000000} /* (26, 28, 13) {real, imag} */,
  {32'hbe471bf2, 32'h00000000} /* (26, 28, 12) {real, imag} */,
  {32'hbc54abef, 32'h00000000} /* (26, 28, 11) {real, imag} */,
  {32'h3e39eb4a, 32'h00000000} /* (26, 28, 10) {real, imag} */,
  {32'h3ec433f5, 32'h00000000} /* (26, 28, 9) {real, imag} */,
  {32'h3ec9753e, 32'h00000000} /* (26, 28, 8) {real, imag} */,
  {32'h3e9b7248, 32'h00000000} /* (26, 28, 7) {real, imag} */,
  {32'h3f4e0598, 32'h00000000} /* (26, 28, 6) {real, imag} */,
  {32'h3ef880b1, 32'h00000000} /* (26, 28, 5) {real, imag} */,
  {32'hbd5ce0e4, 32'h00000000} /* (26, 28, 4) {real, imag} */,
  {32'hbe8af3ef, 32'h00000000} /* (26, 28, 3) {real, imag} */,
  {32'h3e7d255f, 32'h00000000} /* (26, 28, 2) {real, imag} */,
  {32'h3ec86279, 32'h00000000} /* (26, 28, 1) {real, imag} */,
  {32'h3f44af3c, 32'h00000000} /* (26, 28, 0) {real, imag} */,
  {32'h3ea8bfa3, 32'h00000000} /* (26, 27, 31) {real, imag} */,
  {32'hbe551b31, 32'h00000000} /* (26, 27, 30) {real, imag} */,
  {32'hbf0cb8b9, 32'h00000000} /* (26, 27, 29) {real, imag} */,
  {32'h3f0641a9, 32'h00000000} /* (26, 27, 28) {real, imag} */,
  {32'h3f540ee8, 32'h00000000} /* (26, 27, 27) {real, imag} */,
  {32'h3c8ac2b6, 32'h00000000} /* (26, 27, 26) {real, imag} */,
  {32'hbec7f4d4, 32'h00000000} /* (26, 27, 25) {real, imag} */,
  {32'h3d16c353, 32'h00000000} /* (26, 27, 24) {real, imag} */,
  {32'h3f233a9b, 32'h00000000} /* (26, 27, 23) {real, imag} */,
  {32'h3eabebf0, 32'h00000000} /* (26, 27, 22) {real, imag} */,
  {32'h3e682089, 32'h00000000} /* (26, 27, 21) {real, imag} */,
  {32'hbe0ccfc1, 32'h00000000} /* (26, 27, 20) {real, imag} */,
  {32'hbe8a05a7, 32'h00000000} /* (26, 27, 19) {real, imag} */,
  {32'hbf0f569d, 32'h00000000} /* (26, 27, 18) {real, imag} */,
  {32'hbf34a5f7, 32'h00000000} /* (26, 27, 17) {real, imag} */,
  {32'hbe4b8fb7, 32'h00000000} /* (26, 27, 16) {real, imag} */,
  {32'hbf5095c6, 32'h00000000} /* (26, 27, 15) {real, imag} */,
  {32'hbeaa6b55, 32'h00000000} /* (26, 27, 14) {real, imag} */,
  {32'hbe226e1d, 32'h00000000} /* (26, 27, 13) {real, imag} */,
  {32'hbdb04770, 32'h00000000} /* (26, 27, 12) {real, imag} */,
  {32'h3ec5e848, 32'h00000000} /* (26, 27, 11) {real, imag} */,
  {32'h3e8ab0df, 32'h00000000} /* (26, 27, 10) {real, imag} */,
  {32'hbf08fe46, 32'h00000000} /* (26, 27, 9) {real, imag} */,
  {32'h3e31a490, 32'h00000000} /* (26, 27, 8) {real, imag} */,
  {32'h3ec21215, 32'h00000000} /* (26, 27, 7) {real, imag} */,
  {32'h3ee54158, 32'h00000000} /* (26, 27, 6) {real, imag} */,
  {32'h3dcba157, 32'h00000000} /* (26, 27, 5) {real, imag} */,
  {32'hbe45f68a, 32'h00000000} /* (26, 27, 4) {real, imag} */,
  {32'h3dd69fc4, 32'h00000000} /* (26, 27, 3) {real, imag} */,
  {32'h3eb82292, 32'h00000000} /* (26, 27, 2) {real, imag} */,
  {32'h3ec3c4c4, 32'h00000000} /* (26, 27, 1) {real, imag} */,
  {32'h3f0c701d, 32'h00000000} /* (26, 27, 0) {real, imag} */,
  {32'h3db49546, 32'h00000000} /* (26, 26, 31) {real, imag} */,
  {32'hbe9688c8, 32'h00000000} /* (26, 26, 30) {real, imag} */,
  {32'hbf23f071, 32'h00000000} /* (26, 26, 29) {real, imag} */,
  {32'hbeb694b1, 32'h00000000} /* (26, 26, 28) {real, imag} */,
  {32'h3b9a6f76, 32'h00000000} /* (26, 26, 27) {real, imag} */,
  {32'h3db7a1fe, 32'h00000000} /* (26, 26, 26) {real, imag} */,
  {32'h3dc4b3a1, 32'h00000000} /* (26, 26, 25) {real, imag} */,
  {32'h3e6ec150, 32'h00000000} /* (26, 26, 24) {real, imag} */,
  {32'h3efa2e25, 32'h00000000} /* (26, 26, 23) {real, imag} */,
  {32'h3e0e0760, 32'h00000000} /* (26, 26, 22) {real, imag} */,
  {32'hbecc5887, 32'h00000000} /* (26, 26, 21) {real, imag} */,
  {32'hbee03d7b, 32'h00000000} /* (26, 26, 20) {real, imag} */,
  {32'hbe9a8f86, 32'h00000000} /* (26, 26, 19) {real, imag} */,
  {32'hbf12c425, 32'h00000000} /* (26, 26, 18) {real, imag} */,
  {32'hbf5289cc, 32'h00000000} /* (26, 26, 17) {real, imag} */,
  {32'hbd2aa927, 32'h00000000} /* (26, 26, 16) {real, imag} */,
  {32'hbf22faf4, 32'h00000000} /* (26, 26, 15) {real, imag} */,
  {32'hbf3dda24, 32'h00000000} /* (26, 26, 14) {real, imag} */,
  {32'hbe8c79b9, 32'h00000000} /* (26, 26, 13) {real, imag} */,
  {32'hbecb4330, 32'h00000000} /* (26, 26, 12) {real, imag} */,
  {32'hbe93de9b, 32'h00000000} /* (26, 26, 11) {real, imag} */,
  {32'hbec35d4d, 32'h00000000} /* (26, 26, 10) {real, imag} */,
  {32'hbe93dfc1, 32'h00000000} /* (26, 26, 9) {real, imag} */,
  {32'hbd9b5c55, 32'h00000000} /* (26, 26, 8) {real, imag} */,
  {32'hbda605e8, 32'h00000000} /* (26, 26, 7) {real, imag} */,
  {32'h3d07d59a, 32'h00000000} /* (26, 26, 6) {real, imag} */,
  {32'h3ed8f85a, 32'h00000000} /* (26, 26, 5) {real, imag} */,
  {32'h3e9e5b17, 32'h00000000} /* (26, 26, 4) {real, imag} */,
  {32'h3e71fd7b, 32'h00000000} /* (26, 26, 3) {real, imag} */,
  {32'h3e394fc7, 32'h00000000} /* (26, 26, 2) {real, imag} */,
  {32'hbebd5e8c, 32'h00000000} /* (26, 26, 1) {real, imag} */,
  {32'hbdebfb89, 32'h00000000} /* (26, 26, 0) {real, imag} */,
  {32'hbe2501b0, 32'h00000000} /* (26, 25, 31) {real, imag} */,
  {32'hbee6cf0d, 32'h00000000} /* (26, 25, 30) {real, imag} */,
  {32'h3d8767ea, 32'h00000000} /* (26, 25, 29) {real, imag} */,
  {32'hbdc462af, 32'h00000000} /* (26, 25, 28) {real, imag} */,
  {32'hbe016c9d, 32'h00000000} /* (26, 25, 27) {real, imag} */,
  {32'hbe4a7b1a, 32'h00000000} /* (26, 25, 26) {real, imag} */,
  {32'h3d97c766, 32'h00000000} /* (26, 25, 25) {real, imag} */,
  {32'h3e481ad3, 32'h00000000} /* (26, 25, 24) {real, imag} */,
  {32'h3e0cb251, 32'h00000000} /* (26, 25, 23) {real, imag} */,
  {32'h3d3e25dc, 32'h00000000} /* (26, 25, 22) {real, imag} */,
  {32'hbcf4d5a8, 32'h00000000} /* (26, 25, 21) {real, imag} */,
  {32'h3e950b1e, 32'h00000000} /* (26, 25, 20) {real, imag} */,
  {32'h3e2dbc85, 32'h00000000} /* (26, 25, 19) {real, imag} */,
  {32'hbec9a071, 32'h00000000} /* (26, 25, 18) {real, imag} */,
  {32'hbf221cb1, 32'h00000000} /* (26, 25, 17) {real, imag} */,
  {32'h3c8adc05, 32'h00000000} /* (26, 25, 16) {real, imag} */,
  {32'hbf1cdb23, 32'h00000000} /* (26, 25, 15) {real, imag} */,
  {32'hbf090966, 32'h00000000} /* (26, 25, 14) {real, imag} */,
  {32'h3e0431e8, 32'h00000000} /* (26, 25, 13) {real, imag} */,
  {32'hbe1a51e3, 32'h00000000} /* (26, 25, 12) {real, imag} */,
  {32'hbf10fbf8, 32'h00000000} /* (26, 25, 11) {real, imag} */,
  {32'hbe848872, 32'h00000000} /* (26, 25, 10) {real, imag} */,
  {32'h3e097a1a, 32'h00000000} /* (26, 25, 9) {real, imag} */,
  {32'h3ecf0803, 32'h00000000} /* (26, 25, 8) {real, imag} */,
  {32'h3e9ad89a, 32'h00000000} /* (26, 25, 7) {real, imag} */,
  {32'h3e330857, 32'h00000000} /* (26, 25, 6) {real, imag} */,
  {32'h3eeb871f, 32'h00000000} /* (26, 25, 5) {real, imag} */,
  {32'h3ed85257, 32'h00000000} /* (26, 25, 4) {real, imag} */,
  {32'h3e15f6c7, 32'h00000000} /* (26, 25, 3) {real, imag} */,
  {32'h3da0b138, 32'h00000000} /* (26, 25, 2) {real, imag} */,
  {32'hbe2f0f5e, 32'h00000000} /* (26, 25, 1) {real, imag} */,
  {32'hbdbae053, 32'h00000000} /* (26, 25, 0) {real, imag} */,
  {32'hbd5d8402, 32'h00000000} /* (26, 24, 31) {real, imag} */,
  {32'h3d648694, 32'h00000000} /* (26, 24, 30) {real, imag} */,
  {32'h3f03b0c6, 32'h00000000} /* (26, 24, 29) {real, imag} */,
  {32'h3e0a5f8e, 32'h00000000} /* (26, 24, 28) {real, imag} */,
  {32'h3f24ce03, 32'h00000000} /* (26, 24, 27) {real, imag} */,
  {32'h3e61b5c2, 32'h00000000} /* (26, 24, 26) {real, imag} */,
  {32'hbd886bb2, 32'h00000000} /* (26, 24, 25) {real, imag} */,
  {32'h3eff52dc, 32'h00000000} /* (26, 24, 24) {real, imag} */,
  {32'h3d402aa8, 32'h00000000} /* (26, 24, 23) {real, imag} */,
  {32'hbd9f60c4, 32'h00000000} /* (26, 24, 22) {real, imag} */,
  {32'hbcfd04f0, 32'h00000000} /* (26, 24, 21) {real, imag} */,
  {32'h3e851177, 32'h00000000} /* (26, 24, 20) {real, imag} */,
  {32'h3d8f84d7, 32'h00000000} /* (26, 24, 19) {real, imag} */,
  {32'hbe0f4fd4, 32'h00000000} /* (26, 24, 18) {real, imag} */,
  {32'hbef9b057, 32'h00000000} /* (26, 24, 17) {real, imag} */,
  {32'hbee640ae, 32'h00000000} /* (26, 24, 16) {real, imag} */,
  {32'hbe545ae0, 32'h00000000} /* (26, 24, 15) {real, imag} */,
  {32'h3d7bb854, 32'h00000000} /* (26, 24, 14) {real, imag} */,
  {32'h3e1f416f, 32'h00000000} /* (26, 24, 13) {real, imag} */,
  {32'hbf711bc6, 32'h00000000} /* (26, 24, 12) {real, imag} */,
  {32'hbf45800e, 32'h00000000} /* (26, 24, 11) {real, imag} */,
  {32'h3d931e63, 32'h00000000} /* (26, 24, 10) {real, imag} */,
  {32'h3f147984, 32'h00000000} /* (26, 24, 9) {real, imag} */,
  {32'h3f3399f0, 32'h00000000} /* (26, 24, 8) {real, imag} */,
  {32'h3eb0719e, 32'h00000000} /* (26, 24, 7) {real, imag} */,
  {32'hbd5add76, 32'h00000000} /* (26, 24, 6) {real, imag} */,
  {32'hbee4bf20, 32'h00000000} /* (26, 24, 5) {real, imag} */,
  {32'hbf0cc7fa, 32'h00000000} /* (26, 24, 4) {real, imag} */,
  {32'hbdca1989, 32'h00000000} /* (26, 24, 3) {real, imag} */,
  {32'h3e053942, 32'h00000000} /* (26, 24, 2) {real, imag} */,
  {32'h3c4649bd, 32'h00000000} /* (26, 24, 1) {real, imag} */,
  {32'hbe073690, 32'h00000000} /* (26, 24, 0) {real, imag} */,
  {32'hbda7bc72, 32'h00000000} /* (26, 23, 31) {real, imag} */,
  {32'h3df55ea6, 32'h00000000} /* (26, 23, 30) {real, imag} */,
  {32'hbdc6fe1d, 32'h00000000} /* (26, 23, 29) {real, imag} */,
  {32'hbdc90f71, 32'h00000000} /* (26, 23, 28) {real, imag} */,
  {32'h3f1c6b75, 32'h00000000} /* (26, 23, 27) {real, imag} */,
  {32'h3dea40bc, 32'h00000000} /* (26, 23, 26) {real, imag} */,
  {32'hbedb797f, 32'h00000000} /* (26, 23, 25) {real, imag} */,
  {32'h3d34edaa, 32'h00000000} /* (26, 23, 24) {real, imag} */,
  {32'h3d97617a, 32'h00000000} /* (26, 23, 23) {real, imag} */,
  {32'h3e2f2f07, 32'h00000000} /* (26, 23, 22) {real, imag} */,
  {32'h3d6a946a, 32'h00000000} /* (26, 23, 21) {real, imag} */,
  {32'h3d16a4e3, 32'h00000000} /* (26, 23, 20) {real, imag} */,
  {32'hbe4c4f3d, 32'h00000000} /* (26, 23, 19) {real, imag} */,
  {32'hbebb6da1, 32'h00000000} /* (26, 23, 18) {real, imag} */,
  {32'hbea4778b, 32'h00000000} /* (26, 23, 17) {real, imag} */,
  {32'hbe632d0c, 32'h00000000} /* (26, 23, 16) {real, imag} */,
  {32'h3f3c88b3, 32'h00000000} /* (26, 23, 15) {real, imag} */,
  {32'h3e232f03, 32'h00000000} /* (26, 23, 14) {real, imag} */,
  {32'hbe84266a, 32'h00000000} /* (26, 23, 13) {real, imag} */,
  {32'hbf47219f, 32'h00000000} /* (26, 23, 12) {real, imag} */,
  {32'hbebe7065, 32'h00000000} /* (26, 23, 11) {real, imag} */,
  {32'h3eb2c4e7, 32'h00000000} /* (26, 23, 10) {real, imag} */,
  {32'h3e60d153, 32'h00000000} /* (26, 23, 9) {real, imag} */,
  {32'h3f24f112, 32'h00000000} /* (26, 23, 8) {real, imag} */,
  {32'h3ef6a73d, 32'h00000000} /* (26, 23, 7) {real, imag} */,
  {32'hbeac8a04, 32'h00000000} /* (26, 23, 6) {real, imag} */,
  {32'hbf7fa421, 32'h00000000} /* (26, 23, 5) {real, imag} */,
  {32'hbf4275b1, 32'h00000000} /* (26, 23, 4) {real, imag} */,
  {32'hbd6df5b0, 32'h00000000} /* (26, 23, 3) {real, imag} */,
  {32'h3eb25d83, 32'h00000000} /* (26, 23, 2) {real, imag} */,
  {32'hbcc932e5, 32'h00000000} /* (26, 23, 1) {real, imag} */,
  {32'hbe862461, 32'h00000000} /* (26, 23, 0) {real, imag} */,
  {32'h3e31cca6, 32'h00000000} /* (26, 22, 31) {real, imag} */,
  {32'h3e78ac45, 32'h00000000} /* (26, 22, 30) {real, imag} */,
  {32'h3d92ff37, 32'h00000000} /* (26, 22, 29) {real, imag} */,
  {32'hbda77e60, 32'h00000000} /* (26, 22, 28) {real, imag} */,
  {32'hbdaf193e, 32'h00000000} /* (26, 22, 27) {real, imag} */,
  {32'h3dd711f7, 32'h00000000} /* (26, 22, 26) {real, imag} */,
  {32'h3d1a7bc6, 32'h00000000} /* (26, 22, 25) {real, imag} */,
  {32'hbe45fb39, 32'h00000000} /* (26, 22, 24) {real, imag} */,
  {32'h3da6aaba, 32'h00000000} /* (26, 22, 23) {real, imag} */,
  {32'h3eb1862b, 32'h00000000} /* (26, 22, 22) {real, imag} */,
  {32'hbdb73e9d, 32'h00000000} /* (26, 22, 21) {real, imag} */,
  {32'hbf302c73, 32'h00000000} /* (26, 22, 20) {real, imag} */,
  {32'hbf2ae7e0, 32'h00000000} /* (26, 22, 19) {real, imag} */,
  {32'h3e137750, 32'h00000000} /* (26, 22, 18) {real, imag} */,
  {32'h3bdd6b48, 32'h00000000} /* (26, 22, 17) {real, imag} */,
  {32'h3d0a8789, 32'h00000000} /* (26, 22, 16) {real, imag} */,
  {32'h3f083fb3, 32'h00000000} /* (26, 22, 15) {real, imag} */,
  {32'h3e17fd94, 32'h00000000} /* (26, 22, 14) {real, imag} */,
  {32'h3c6c0adb, 32'h00000000} /* (26, 22, 13) {real, imag} */,
  {32'h3eb70379, 32'h00000000} /* (26, 22, 12) {real, imag} */,
  {32'h3efc6941, 32'h00000000} /* (26, 22, 11) {real, imag} */,
  {32'h3f14adfe, 32'h00000000} /* (26, 22, 10) {real, imag} */,
  {32'h3ca209d1, 32'h00000000} /* (26, 22, 9) {real, imag} */,
  {32'h3ef18a14, 32'h00000000} /* (26, 22, 8) {real, imag} */,
  {32'h3f1ea4b3, 32'h00000000} /* (26, 22, 7) {real, imag} */,
  {32'h3eb62a14, 32'h00000000} /* (26, 22, 6) {real, imag} */,
  {32'hbe6d7c95, 32'h00000000} /* (26, 22, 5) {real, imag} */,
  {32'hbd200fa5, 32'h00000000} /* (26, 22, 4) {real, imag} */,
  {32'h3eea53a7, 32'h00000000} /* (26, 22, 3) {real, imag} */,
  {32'h3f25ee1d, 32'h00000000} /* (26, 22, 2) {real, imag} */,
  {32'h3ee480da, 32'h00000000} /* (26, 22, 1) {real, imag} */,
  {32'h3e9ecfe7, 32'h00000000} /* (26, 22, 0) {real, imag} */,
  {32'h3d82de0d, 32'h00000000} /* (26, 21, 31) {real, imag} */,
  {32'h3daa7ab0, 32'h00000000} /* (26, 21, 30) {real, imag} */,
  {32'hbd8826e3, 32'h00000000} /* (26, 21, 29) {real, imag} */,
  {32'hbeab8f75, 32'h00000000} /* (26, 21, 28) {real, imag} */,
  {32'hbf0d8880, 32'h00000000} /* (26, 21, 27) {real, imag} */,
  {32'hbea1703f, 32'h00000000} /* (26, 21, 26) {real, imag} */,
  {32'hbee6f380, 32'h00000000} /* (26, 21, 25) {real, imag} */,
  {32'hbebd1552, 32'h00000000} /* (26, 21, 24) {real, imag} */,
  {32'hbeb44091, 32'h00000000} /* (26, 21, 23) {real, imag} */,
  {32'h3e15b937, 32'h00000000} /* (26, 21, 22) {real, imag} */,
  {32'h3e5b022d, 32'h00000000} /* (26, 21, 21) {real, imag} */,
  {32'hbe95e2b6, 32'h00000000} /* (26, 21, 20) {real, imag} */,
  {32'hbe9a64de, 32'h00000000} /* (26, 21, 19) {real, imag} */,
  {32'h3f1a9b0c, 32'h00000000} /* (26, 21, 18) {real, imag} */,
  {32'h3e793260, 32'h00000000} /* (26, 21, 17) {real, imag} */,
  {32'h3cf26576, 32'h00000000} /* (26, 21, 16) {real, imag} */,
  {32'hbc6b2b26, 32'h00000000} /* (26, 21, 15) {real, imag} */,
  {32'h3e25a5f9, 32'h00000000} /* (26, 21, 14) {real, imag} */,
  {32'h3eafd1c8, 32'h00000000} /* (26, 21, 13) {real, imag} */,
  {32'h3e755fe8, 32'h00000000} /* (26, 21, 12) {real, imag} */,
  {32'hbd045ff3, 32'h00000000} /* (26, 21, 11) {real, imag} */,
  {32'h3d5134da, 32'h00000000} /* (26, 21, 10) {real, imag} */,
  {32'hbe68746a, 32'h00000000} /* (26, 21, 9) {real, imag} */,
  {32'hbea795b6, 32'h00000000} /* (26, 21, 8) {real, imag} */,
  {32'h3e40a516, 32'h00000000} /* (26, 21, 7) {real, imag} */,
  {32'h3f8bfd05, 32'h00000000} /* (26, 21, 6) {real, imag} */,
  {32'h3ef74702, 32'h00000000} /* (26, 21, 5) {real, imag} */,
  {32'h3eabe233, 32'h00000000} /* (26, 21, 4) {real, imag} */,
  {32'h3f14d528, 32'h00000000} /* (26, 21, 3) {real, imag} */,
  {32'h3f3b97ff, 32'h00000000} /* (26, 21, 2) {real, imag} */,
  {32'h3eaa4bc2, 32'h00000000} /* (26, 21, 1) {real, imag} */,
  {32'h3eae3879, 32'h00000000} /* (26, 21, 0) {real, imag} */,
  {32'h3e30634e, 32'h00000000} /* (26, 20, 31) {real, imag} */,
  {32'h3e5f6c62, 32'h00000000} /* (26, 20, 30) {real, imag} */,
  {32'h3dc9b1ab, 32'h00000000} /* (26, 20, 29) {real, imag} */,
  {32'h3e2f07a9, 32'h00000000} /* (26, 20, 28) {real, imag} */,
  {32'hbe43d673, 32'h00000000} /* (26, 20, 27) {real, imag} */,
  {32'hbe7c8c57, 32'h00000000} /* (26, 20, 26) {real, imag} */,
  {32'hbf175bd0, 32'h00000000} /* (26, 20, 25) {real, imag} */,
  {32'hbe10788d, 32'h00000000} /* (26, 20, 24) {real, imag} */,
  {32'h3ecbf110, 32'h00000000} /* (26, 20, 23) {real, imag} */,
  {32'h3e7b9ed6, 32'h00000000} /* (26, 20, 22) {real, imag} */,
  {32'h3e6a1850, 32'h00000000} /* (26, 20, 21) {real, imag} */,
  {32'hbd226664, 32'h00000000} /* (26, 20, 20) {real, imag} */,
  {32'hbde43ef1, 32'h00000000} /* (26, 20, 19) {real, imag} */,
  {32'h3ebd3c5c, 32'h00000000} /* (26, 20, 18) {real, imag} */,
  {32'h3e278fa4, 32'h00000000} /* (26, 20, 17) {real, imag} */,
  {32'h3ec75c31, 32'h00000000} /* (26, 20, 16) {real, imag} */,
  {32'h3c1add5f, 32'h00000000} /* (26, 20, 15) {real, imag} */,
  {32'hbda6483c, 32'h00000000} /* (26, 20, 14) {real, imag} */,
  {32'hbafc0d38, 32'h00000000} /* (26, 20, 13) {real, imag} */,
  {32'hbe442b8b, 32'h00000000} /* (26, 20, 12) {real, imag} */,
  {32'hbed6e8b3, 32'h00000000} /* (26, 20, 11) {real, imag} */,
  {32'hbf193589, 32'h00000000} /* (26, 20, 10) {real, imag} */,
  {32'hbe773722, 32'h00000000} /* (26, 20, 9) {real, imag} */,
  {32'h3e2ace82, 32'h00000000} /* (26, 20, 8) {real, imag} */,
  {32'hbd0088ce, 32'h00000000} /* (26, 20, 7) {real, imag} */,
  {32'h3d0bf11b, 32'h00000000} /* (26, 20, 6) {real, imag} */,
  {32'hbf17f19a, 32'h00000000} /* (26, 20, 5) {real, imag} */,
  {32'hbe6df1c8, 32'h00000000} /* (26, 20, 4) {real, imag} */,
  {32'hbd895643, 32'h00000000} /* (26, 20, 3) {real, imag} */,
  {32'hbd6bc8b0, 32'h00000000} /* (26, 20, 2) {real, imag} */,
  {32'h3b97e9bc, 32'h00000000} /* (26, 20, 1) {real, imag} */,
  {32'h3da31a4d, 32'h00000000} /* (26, 20, 0) {real, imag} */,
  {32'h3e991ee2, 32'h00000000} /* (26, 19, 31) {real, imag} */,
  {32'h3e9c7dbf, 32'h00000000} /* (26, 19, 30) {real, imag} */,
  {32'hbe128479, 32'h00000000} /* (26, 19, 29) {real, imag} */,
  {32'h3ddaa539, 32'h00000000} /* (26, 19, 28) {real, imag} */,
  {32'hbdeb123c, 32'h00000000} /* (26, 19, 27) {real, imag} */,
  {32'h3dac27d3, 32'h00000000} /* (26, 19, 26) {real, imag} */,
  {32'hbd14a2e4, 32'h00000000} /* (26, 19, 25) {real, imag} */,
  {32'hbe128631, 32'h00000000} /* (26, 19, 24) {real, imag} */,
  {32'h3e0d206c, 32'h00000000} /* (26, 19, 23) {real, imag} */,
  {32'h3bdd5570, 32'h00000000} /* (26, 19, 22) {real, imag} */,
  {32'h3c404a8b, 32'h00000000} /* (26, 19, 21) {real, imag} */,
  {32'h3b88ca43, 32'h00000000} /* (26, 19, 20) {real, imag} */,
  {32'h3e065719, 32'h00000000} /* (26, 19, 19) {real, imag} */,
  {32'hbe4c24ac, 32'h00000000} /* (26, 19, 18) {real, imag} */,
  {32'hbe481442, 32'h00000000} /* (26, 19, 17) {real, imag} */,
  {32'h3f669ee3, 32'h00000000} /* (26, 19, 16) {real, imag} */,
  {32'h3f4f4318, 32'h00000000} /* (26, 19, 15) {real, imag} */,
  {32'h3e7944fa, 32'h00000000} /* (26, 19, 14) {real, imag} */,
  {32'h3d9cfeff, 32'h00000000} /* (26, 19, 13) {real, imag} */,
  {32'hbdc8733f, 32'h00000000} /* (26, 19, 12) {real, imag} */,
  {32'h3e8abf8c, 32'h00000000} /* (26, 19, 11) {real, imag} */,
  {32'h3da7b70d, 32'h00000000} /* (26, 19, 10) {real, imag} */,
  {32'h3d4855cc, 32'h00000000} /* (26, 19, 9) {real, imag} */,
  {32'h3e50f324, 32'h00000000} /* (26, 19, 8) {real, imag} */,
  {32'hbc8a7324, 32'h00000000} /* (26, 19, 7) {real, imag} */,
  {32'hbe0e3f96, 32'h00000000} /* (26, 19, 6) {real, imag} */,
  {32'hbf2b5d92, 32'h00000000} /* (26, 19, 5) {real, imag} */,
  {32'hbf514746, 32'h00000000} /* (26, 19, 4) {real, imag} */,
  {32'hbf17479f, 32'h00000000} /* (26, 19, 3) {real, imag} */,
  {32'hbeacf5b9, 32'h00000000} /* (26, 19, 2) {real, imag} */,
  {32'h3d31ddd6, 32'h00000000} /* (26, 19, 1) {real, imag} */,
  {32'h3cfa1ab0, 32'h00000000} /* (26, 19, 0) {real, imag} */,
  {32'h3f001cb4, 32'h00000000} /* (26, 18, 31) {real, imag} */,
  {32'h3e4931fb, 32'h00000000} /* (26, 18, 30) {real, imag} */,
  {32'hbdc2707c, 32'h00000000} /* (26, 18, 29) {real, imag} */,
  {32'hbde8fffd, 32'h00000000} /* (26, 18, 28) {real, imag} */,
  {32'hbe4e3104, 32'h00000000} /* (26, 18, 27) {real, imag} */,
  {32'h3e2901ce, 32'h00000000} /* (26, 18, 26) {real, imag} */,
  {32'hbda19976, 32'h00000000} /* (26, 18, 25) {real, imag} */,
  {32'hbeeb211b, 32'h00000000} /* (26, 18, 24) {real, imag} */,
  {32'hbf37b3c2, 32'h00000000} /* (26, 18, 23) {real, imag} */,
  {32'hbefc4818, 32'h00000000} /* (26, 18, 22) {real, imag} */,
  {32'hbe39af6f, 32'h00000000} /* (26, 18, 21) {real, imag} */,
  {32'hbe252df0, 32'h00000000} /* (26, 18, 20) {real, imag} */,
  {32'h3d98f1a0, 32'h00000000} /* (26, 18, 19) {real, imag} */,
  {32'hbe0bd762, 32'h00000000} /* (26, 18, 18) {real, imag} */,
  {32'h3e2a1b4a, 32'h00000000} /* (26, 18, 17) {real, imag} */,
  {32'h3f1a9c47, 32'h00000000} /* (26, 18, 16) {real, imag} */,
  {32'h3f295879, 32'h00000000} /* (26, 18, 15) {real, imag} */,
  {32'h3e9b28cc, 32'h00000000} /* (26, 18, 14) {real, imag} */,
  {32'hbe760397, 32'h00000000} /* (26, 18, 13) {real, imag} */,
  {32'hbe645b9e, 32'h00000000} /* (26, 18, 12) {real, imag} */,
  {32'h3f1b86c2, 32'h00000000} /* (26, 18, 11) {real, imag} */,
  {32'h3ec59e1e, 32'h00000000} /* (26, 18, 10) {real, imag} */,
  {32'h3dc928b5, 32'h00000000} /* (26, 18, 9) {real, imag} */,
  {32'h3c235e7f, 32'h00000000} /* (26, 18, 8) {real, imag} */,
  {32'h3d73687a, 32'h00000000} /* (26, 18, 7) {real, imag} */,
  {32'hbda264a7, 32'h00000000} /* (26, 18, 6) {real, imag} */,
  {32'hbe789a99, 32'h00000000} /* (26, 18, 5) {real, imag} */,
  {32'hbef884cb, 32'h00000000} /* (26, 18, 4) {real, imag} */,
  {32'hbf145cfd, 32'h00000000} /* (26, 18, 3) {real, imag} */,
  {32'h3e206efa, 32'h00000000} /* (26, 18, 2) {real, imag} */,
  {32'h3e7b057c, 32'h00000000} /* (26, 18, 1) {real, imag} */,
  {32'h3ace6fc0, 32'h00000000} /* (26, 18, 0) {real, imag} */,
  {32'h3b61bf82, 32'h00000000} /* (26, 17, 31) {real, imag} */,
  {32'hbe5fa8f9, 32'h00000000} /* (26, 17, 30) {real, imag} */,
  {32'h3c0ac38a, 32'h00000000} /* (26, 17, 29) {real, imag} */,
  {32'hbdfc5b74, 32'h00000000} /* (26, 17, 28) {real, imag} */,
  {32'hbda5b3af, 32'h00000000} /* (26, 17, 27) {real, imag} */,
  {32'h3f13ad68, 32'h00000000} /* (26, 17, 26) {real, imag} */,
  {32'hbe1ac4c7, 32'h00000000} /* (26, 17, 25) {real, imag} */,
  {32'hbe9c908b, 32'h00000000} /* (26, 17, 24) {real, imag} */,
  {32'hbed23bdf, 32'h00000000} /* (26, 17, 23) {real, imag} */,
  {32'hbe8fdc5a, 32'h00000000} /* (26, 17, 22) {real, imag} */,
  {32'hbed0e83d, 32'h00000000} /* (26, 17, 21) {real, imag} */,
  {32'hbeae0523, 32'h00000000} /* (26, 17, 20) {real, imag} */,
  {32'h3da5f46a, 32'h00000000} /* (26, 17, 19) {real, imag} */,
  {32'h3ecb9092, 32'h00000000} /* (26, 17, 18) {real, imag} */,
  {32'h3f2af01c, 32'h00000000} /* (26, 17, 17) {real, imag} */,
  {32'h3eec07d2, 32'h00000000} /* (26, 17, 16) {real, imag} */,
  {32'h3ef0da3e, 32'h00000000} /* (26, 17, 15) {real, imag} */,
  {32'h3ebf481e, 32'h00000000} /* (26, 17, 14) {real, imag} */,
  {32'hbea6482e, 32'h00000000} /* (26, 17, 13) {real, imag} */,
  {32'hbdf2038e, 32'h00000000} /* (26, 17, 12) {real, imag} */,
  {32'h3e785eb1, 32'h00000000} /* (26, 17, 11) {real, imag} */,
  {32'h3ebb3b89, 32'h00000000} /* (26, 17, 10) {real, imag} */,
  {32'h3e9cb866, 32'h00000000} /* (26, 17, 9) {real, imag} */,
  {32'h3e28c8f3, 32'h00000000} /* (26, 17, 8) {real, imag} */,
  {32'h3f28fe51, 32'h00000000} /* (26, 17, 7) {real, imag} */,
  {32'h3ee8cb74, 32'h00000000} /* (26, 17, 6) {real, imag} */,
  {32'hbe217746, 32'h00000000} /* (26, 17, 5) {real, imag} */,
  {32'hbe34a53b, 32'h00000000} /* (26, 17, 4) {real, imag} */,
  {32'hbee102f7, 32'h00000000} /* (26, 17, 3) {real, imag} */,
  {32'hbf1b8683, 32'h00000000} /* (26, 17, 2) {real, imag} */,
  {32'hbe5b2b71, 32'h00000000} /* (26, 17, 1) {real, imag} */,
  {32'hbda7e2a2, 32'h00000000} /* (26, 17, 0) {real, imag} */,
  {32'hbe4b4b46, 32'h00000000} /* (26, 16, 31) {real, imag} */,
  {32'hbe00915f, 32'h00000000} /* (26, 16, 30) {real, imag} */,
  {32'h3d28d722, 32'h00000000} /* (26, 16, 29) {real, imag} */,
  {32'h3eb6c09e, 32'h00000000} /* (26, 16, 28) {real, imag} */,
  {32'hbe8ea81a, 32'h00000000} /* (26, 16, 27) {real, imag} */,
  {32'hbd039a9d, 32'h00000000} /* (26, 16, 26) {real, imag} */,
  {32'hbea060aa, 32'h00000000} /* (26, 16, 25) {real, imag} */,
  {32'h3d330a79, 32'h00000000} /* (26, 16, 24) {real, imag} */,
  {32'h3d99dfd4, 32'h00000000} /* (26, 16, 23) {real, imag} */,
  {32'hbed28c36, 32'h00000000} /* (26, 16, 22) {real, imag} */,
  {32'hbe1b1932, 32'h00000000} /* (26, 16, 21) {real, imag} */,
  {32'h3d957fb8, 32'h00000000} /* (26, 16, 20) {real, imag} */,
  {32'h3e5ffa53, 32'h00000000} /* (26, 16, 19) {real, imag} */,
  {32'h3ec93929, 32'h00000000} /* (26, 16, 18) {real, imag} */,
  {32'h3da9ae21, 32'h00000000} /* (26, 16, 17) {real, imag} */,
  {32'h3e571946, 32'h00000000} /* (26, 16, 16) {real, imag} */,
  {32'h3eb9cfed, 32'h00000000} /* (26, 16, 15) {real, imag} */,
  {32'h3e144742, 32'h00000000} /* (26, 16, 14) {real, imag} */,
  {32'h3d1d031c, 32'h00000000} /* (26, 16, 13) {real, imag} */,
  {32'h3f0b8a4b, 32'h00000000} /* (26, 16, 12) {real, imag} */,
  {32'h3e04af5c, 32'h00000000} /* (26, 16, 11) {real, imag} */,
  {32'h3e9e4259, 32'h00000000} /* (26, 16, 10) {real, imag} */,
  {32'h3e83cd3b, 32'h00000000} /* (26, 16, 9) {real, imag} */,
  {32'h3c59f8bb, 32'h00000000} /* (26, 16, 8) {real, imag} */,
  {32'h3f149336, 32'h00000000} /* (26, 16, 7) {real, imag} */,
  {32'h3f612c13, 32'h00000000} /* (26, 16, 6) {real, imag} */,
  {32'h3ca4315a, 32'h00000000} /* (26, 16, 5) {real, imag} */,
  {32'hbe32860d, 32'h00000000} /* (26, 16, 4) {real, imag} */,
  {32'hbeb7a9a8, 32'h00000000} /* (26, 16, 3) {real, imag} */,
  {32'hbf1008bd, 32'h00000000} /* (26, 16, 2) {real, imag} */,
  {32'hbe69300f, 32'h00000000} /* (26, 16, 1) {real, imag} */,
  {32'h3dabd660, 32'h00000000} /* (26, 16, 0) {real, imag} */,
  {32'hbeb3de3d, 32'h00000000} /* (26, 15, 31) {real, imag} */,
  {32'hbf281ab5, 32'h00000000} /* (26, 15, 30) {real, imag} */,
  {32'hbf489d95, 32'h00000000} /* (26, 15, 29) {real, imag} */,
  {32'h3e11a7c4, 32'h00000000} /* (26, 15, 28) {real, imag} */,
  {32'hbea6d978, 32'h00000000} /* (26, 15, 27) {real, imag} */,
  {32'hbee444fe, 32'h00000000} /* (26, 15, 26) {real, imag} */,
  {32'hbf3ac11b, 32'h00000000} /* (26, 15, 25) {real, imag} */,
  {32'h3ea0ba17, 32'h00000000} /* (26, 15, 24) {real, imag} */,
  {32'h3e97069a, 32'h00000000} /* (26, 15, 23) {real, imag} */,
  {32'hbf6b9578, 32'h00000000} /* (26, 15, 22) {real, imag} */,
  {32'hbeb21639, 32'h00000000} /* (26, 15, 21) {real, imag} */,
  {32'hbd2926ce, 32'h00000000} /* (26, 15, 20) {real, imag} */,
  {32'hbe95ce5e, 32'h00000000} /* (26, 15, 19) {real, imag} */,
  {32'hbef00fd9, 32'h00000000} /* (26, 15, 18) {real, imag} */,
  {32'hbf48f386, 32'h00000000} /* (26, 15, 17) {real, imag} */,
  {32'h3d8c1f5f, 32'h00000000} /* (26, 15, 16) {real, imag} */,
  {32'h3e54e9d9, 32'h00000000} /* (26, 15, 15) {real, imag} */,
  {32'hbd9ef4cb, 32'h00000000} /* (26, 15, 14) {real, imag} */,
  {32'h3e1e5ab4, 32'h00000000} /* (26, 15, 13) {real, imag} */,
  {32'h3ed04a5e, 32'h00000000} /* (26, 15, 12) {real, imag} */,
  {32'h3e73674a, 32'h00000000} /* (26, 15, 11) {real, imag} */,
  {32'hbe3a7f00, 32'h00000000} /* (26, 15, 10) {real, imag} */,
  {32'hbe846585, 32'h00000000} /* (26, 15, 9) {real, imag} */,
  {32'hbede909c, 32'h00000000} /* (26, 15, 8) {real, imag} */,
  {32'hbeb62699, 32'h00000000} /* (26, 15, 7) {real, imag} */,
  {32'hbd5465bf, 32'h00000000} /* (26, 15, 6) {real, imag} */,
  {32'hbefddba3, 32'h00000000} /* (26, 15, 5) {real, imag} */,
  {32'hbecd4a05, 32'h00000000} /* (26, 15, 4) {real, imag} */,
  {32'hbf273df6, 32'h00000000} /* (26, 15, 3) {real, imag} */,
  {32'hbf378d2a, 32'h00000000} /* (26, 15, 2) {real, imag} */,
  {32'hbe8f11bb, 32'h00000000} /* (26, 15, 1) {real, imag} */,
  {32'hbdfd4f70, 32'h00000000} /* (26, 15, 0) {real, imag} */,
  {32'hbe94196c, 32'h00000000} /* (26, 14, 31) {real, imag} */,
  {32'hbf520874, 32'h00000000} /* (26, 14, 30) {real, imag} */,
  {32'hbf5d2fb1, 32'h00000000} /* (26, 14, 29) {real, imag} */,
  {32'hbf075fdb, 32'h00000000} /* (26, 14, 28) {real, imag} */,
  {32'hbee0ee0e, 32'h00000000} /* (26, 14, 27) {real, imag} */,
  {32'hbec4b780, 32'h00000000} /* (26, 14, 26) {real, imag} */,
  {32'hbf71d1a5, 32'h00000000} /* (26, 14, 25) {real, imag} */,
  {32'hbebf160d, 32'h00000000} /* (26, 14, 24) {real, imag} */,
  {32'hbecac004, 32'h00000000} /* (26, 14, 23) {real, imag} */,
  {32'hbf761ae5, 32'h00000000} /* (26, 14, 22) {real, imag} */,
  {32'hbee540ea, 32'h00000000} /* (26, 14, 21) {real, imag} */,
  {32'h3daba51e, 32'h00000000} /* (26, 14, 20) {real, imag} */,
  {32'h3e208d9b, 32'h00000000} /* (26, 14, 19) {real, imag} */,
  {32'h3da12bfd, 32'h00000000} /* (26, 14, 18) {real, imag} */,
  {32'hbe7c4cd1, 32'h00000000} /* (26, 14, 17) {real, imag} */,
  {32'hbd82e0d4, 32'h00000000} /* (26, 14, 16) {real, imag} */,
  {32'h3e03eacc, 32'h00000000} /* (26, 14, 15) {real, imag} */,
  {32'hbcd31d78, 32'h00000000} /* (26, 14, 14) {real, imag} */,
  {32'hbe0d28b1, 32'h00000000} /* (26, 14, 13) {real, imag} */,
  {32'h3d9e59ae, 32'h00000000} /* (26, 14, 12) {real, imag} */,
  {32'h3d8be18b, 32'h00000000} /* (26, 14, 11) {real, imag} */,
  {32'hbe90301f, 32'h00000000} /* (26, 14, 10) {real, imag} */,
  {32'hbec371b4, 32'h00000000} /* (26, 14, 9) {real, imag} */,
  {32'hbe85ce25, 32'h00000000} /* (26, 14, 8) {real, imag} */,
  {32'hbe9dd6ea, 32'h00000000} /* (26, 14, 7) {real, imag} */,
  {32'hbe9cc83f, 32'h00000000} /* (26, 14, 6) {real, imag} */,
  {32'hbeef5914, 32'h00000000} /* (26, 14, 5) {real, imag} */,
  {32'hbc0f06e7, 32'h00000000} /* (26, 14, 4) {real, imag} */,
  {32'hbd122873, 32'h00000000} /* (26, 14, 3) {real, imag} */,
  {32'hbf1df9b9, 32'h00000000} /* (26, 14, 2) {real, imag} */,
  {32'hbe833729, 32'h00000000} /* (26, 14, 1) {real, imag} */,
  {32'hbd6650fb, 32'h00000000} /* (26, 14, 0) {real, imag} */,
  {32'hbe40111c, 32'h00000000} /* (26, 13, 31) {real, imag} */,
  {32'hbef127d3, 32'h00000000} /* (26, 13, 30) {real, imag} */,
  {32'hbf14af19, 32'h00000000} /* (26, 13, 29) {real, imag} */,
  {32'hbe2a5980, 32'h00000000} /* (26, 13, 28) {real, imag} */,
  {32'h3e815b19, 32'h00000000} /* (26, 13, 27) {real, imag} */,
  {32'hbd9d52f0, 32'h00000000} /* (26, 13, 26) {real, imag} */,
  {32'hbf09d6b4, 32'h00000000} /* (26, 13, 25) {real, imag} */,
  {32'hbf06767c, 32'h00000000} /* (26, 13, 24) {real, imag} */,
  {32'hbe8aace9, 32'h00000000} /* (26, 13, 23) {real, imag} */,
  {32'hbf0d8a44, 32'h00000000} /* (26, 13, 22) {real, imag} */,
  {32'hbefadaca, 32'h00000000} /* (26, 13, 21) {real, imag} */,
  {32'h3ce3db18, 32'h00000000} /* (26, 13, 20) {real, imag} */,
  {32'h3e762dfb, 32'h00000000} /* (26, 13, 19) {real, imag} */,
  {32'h3f2f822b, 32'h00000000} /* (26, 13, 18) {real, imag} */,
  {32'h3e311f3c, 32'h00000000} /* (26, 13, 17) {real, imag} */,
  {32'hbec6cd11, 32'h00000000} /* (26, 13, 16) {real, imag} */,
  {32'hbee72846, 32'h00000000} /* (26, 13, 15) {real, imag} */,
  {32'hbebed051, 32'h00000000} /* (26, 13, 14) {real, imag} */,
  {32'hbdcff264, 32'h00000000} /* (26, 13, 13) {real, imag} */,
  {32'h3daee134, 32'h00000000} /* (26, 13, 12) {real, imag} */,
  {32'h3e614045, 32'h00000000} /* (26, 13, 11) {real, imag} */,
  {32'h3e0fd305, 32'h00000000} /* (26, 13, 10) {real, imag} */,
  {32'hbd8405be, 32'h00000000} /* (26, 13, 9) {real, imag} */,
  {32'hbeacdabc, 32'h00000000} /* (26, 13, 8) {real, imag} */,
  {32'hbf3fdcc6, 32'h00000000} /* (26, 13, 7) {real, imag} */,
  {32'hbef18db3, 32'h00000000} /* (26, 13, 6) {real, imag} */,
  {32'hbcf7ee48, 32'h00000000} /* (26, 13, 5) {real, imag} */,
  {32'h3ea5fd2f, 32'h00000000} /* (26, 13, 4) {real, imag} */,
  {32'hbd7c6938, 32'h00000000} /* (26, 13, 3) {real, imag} */,
  {32'hbef9f318, 32'h00000000} /* (26, 13, 2) {real, imag} */,
  {32'hbecfc216, 32'h00000000} /* (26, 13, 1) {real, imag} */,
  {32'hbb133f2e, 32'h00000000} /* (26, 13, 0) {real, imag} */,
  {32'h3c047690, 32'h00000000} /* (26, 12, 31) {real, imag} */,
  {32'h3debaefa, 32'h00000000} /* (26, 12, 30) {real, imag} */,
  {32'hbc0ca6c2, 32'h00000000} /* (26, 12, 29) {real, imag} */,
  {32'h3dd40ac3, 32'h00000000} /* (26, 12, 28) {real, imag} */,
  {32'h3dfe80d5, 32'h00000000} /* (26, 12, 27) {real, imag} */,
  {32'hbdd996ea, 32'h00000000} /* (26, 12, 26) {real, imag} */,
  {32'hbec77c45, 32'h00000000} /* (26, 12, 25) {real, imag} */,
  {32'hbd2b752f, 32'h00000000} /* (26, 12, 24) {real, imag} */,
  {32'h3dd0b45b, 32'h00000000} /* (26, 12, 23) {real, imag} */,
  {32'hbdd2e03c, 32'h00000000} /* (26, 12, 22) {real, imag} */,
  {32'h3e119684, 32'h00000000} /* (26, 12, 21) {real, imag} */,
  {32'hbd32858f, 32'h00000000} /* (26, 12, 20) {real, imag} */,
  {32'hbe4d97d7, 32'h00000000} /* (26, 12, 19) {real, imag} */,
  {32'h3ea67392, 32'h00000000} /* (26, 12, 18) {real, imag} */,
  {32'h3ec4aeeb, 32'h00000000} /* (26, 12, 17) {real, imag} */,
  {32'hbd8d6785, 32'h00000000} /* (26, 12, 16) {real, imag} */,
  {32'hbe0072d0, 32'h00000000} /* (26, 12, 15) {real, imag} */,
  {32'hbe0e1fcc, 32'h00000000} /* (26, 12, 14) {real, imag} */,
  {32'h3d9933fd, 32'h00000000} /* (26, 12, 13) {real, imag} */,
  {32'hbe0b736c, 32'h00000000} /* (26, 12, 12) {real, imag} */,
  {32'h3df89b98, 32'h00000000} /* (26, 12, 11) {real, imag} */,
  {32'h3ea140be, 32'h00000000} /* (26, 12, 10) {real, imag} */,
  {32'hbc6a73f4, 32'h00000000} /* (26, 12, 9) {real, imag} */,
  {32'hbf010616, 32'h00000000} /* (26, 12, 8) {real, imag} */,
  {32'hbf0f0056, 32'h00000000} /* (26, 12, 7) {real, imag} */,
  {32'hbf0ed358, 32'h00000000} /* (26, 12, 6) {real, imag} */,
  {32'hbed9c680, 32'h00000000} /* (26, 12, 5) {real, imag} */,
  {32'hbe288451, 32'h00000000} /* (26, 12, 4) {real, imag} */,
  {32'hbf1931f1, 32'h00000000} /* (26, 12, 3) {real, imag} */,
  {32'hbee2bf4d, 32'h00000000} /* (26, 12, 2) {real, imag} */,
  {32'hbf0bf341, 32'h00000000} /* (26, 12, 1) {real, imag} */,
  {32'h3d6254c2, 32'h00000000} /* (26, 12, 0) {real, imag} */,
  {32'h3eb34882, 32'h00000000} /* (26, 11, 31) {real, imag} */,
  {32'h3f0d8935, 32'h00000000} /* (26, 11, 30) {real, imag} */,
  {32'hbdc83789, 32'h00000000} /* (26, 11, 29) {real, imag} */,
  {32'hbe507551, 32'h00000000} /* (26, 11, 28) {real, imag} */,
  {32'h3e3f47e4, 32'h00000000} /* (26, 11, 27) {real, imag} */,
  {32'hbdd3350a, 32'h00000000} /* (26, 11, 26) {real, imag} */,
  {32'hbe1f2a89, 32'h00000000} /* (26, 11, 25) {real, imag} */,
  {32'h3ee8ebb7, 32'h00000000} /* (26, 11, 24) {real, imag} */,
  {32'h3f02b36c, 32'h00000000} /* (26, 11, 23) {real, imag} */,
  {32'h3f02b28e, 32'h00000000} /* (26, 11, 22) {real, imag} */,
  {32'h3f2ea516, 32'h00000000} /* (26, 11, 21) {real, imag} */,
  {32'h3f227381, 32'h00000000} /* (26, 11, 20) {real, imag} */,
  {32'hbdb9106e, 32'h00000000} /* (26, 11, 19) {real, imag} */,
  {32'h3dfddd93, 32'h00000000} /* (26, 11, 18) {real, imag} */,
  {32'h3f05c573, 32'h00000000} /* (26, 11, 17) {real, imag} */,
  {32'h3eb13cc0, 32'h00000000} /* (26, 11, 16) {real, imag} */,
  {32'h3eade9c4, 32'h00000000} /* (26, 11, 15) {real, imag} */,
  {32'hbddf7822, 32'h00000000} /* (26, 11, 14) {real, imag} */,
  {32'hbe64915f, 32'h00000000} /* (26, 11, 13) {real, imag} */,
  {32'hbd836ff8, 32'h00000000} /* (26, 11, 12) {real, imag} */,
  {32'hbda9d9e5, 32'h00000000} /* (26, 11, 11) {real, imag} */,
  {32'h3e34f983, 32'h00000000} /* (26, 11, 10) {real, imag} */,
  {32'h3e5b9841, 32'h00000000} /* (26, 11, 9) {real, imag} */,
  {32'h3e9abe18, 32'h00000000} /* (26, 11, 8) {real, imag} */,
  {32'h3f00595d, 32'h00000000} /* (26, 11, 7) {real, imag} */,
  {32'hbe254c50, 32'h00000000} /* (26, 11, 6) {real, imag} */,
  {32'hbe8aa1bf, 32'h00000000} /* (26, 11, 5) {real, imag} */,
  {32'h3e1da12c, 32'h00000000} /* (26, 11, 4) {real, imag} */,
  {32'hbf06229c, 32'h00000000} /* (26, 11, 3) {real, imag} */,
  {32'hbe99b413, 32'h00000000} /* (26, 11, 2) {real, imag} */,
  {32'hbdc69abd, 32'h00000000} /* (26, 11, 1) {real, imag} */,
  {32'h3e4ca213, 32'h00000000} /* (26, 11, 0) {real, imag} */,
  {32'h3eb10347, 32'h00000000} /* (26, 10, 31) {real, imag} */,
  {32'h3f1f31e1, 32'h00000000} /* (26, 10, 30) {real, imag} */,
  {32'hbe259bbe, 32'h00000000} /* (26, 10, 29) {real, imag} */,
  {32'hbdeb5440, 32'h00000000} /* (26, 10, 28) {real, imag} */,
  {32'h3e9a3b35, 32'h00000000} /* (26, 10, 27) {real, imag} */,
  {32'h3e795e28, 32'h00000000} /* (26, 10, 26) {real, imag} */,
  {32'hbcb55bf5, 32'h00000000} /* (26, 10, 25) {real, imag} */,
  {32'h3ebe0043, 32'h00000000} /* (26, 10, 24) {real, imag} */,
  {32'h3ed6d483, 32'h00000000} /* (26, 10, 23) {real, imag} */,
  {32'h3e13aadf, 32'h00000000} /* (26, 10, 22) {real, imag} */,
  {32'h3a6539c0, 32'h00000000} /* (26, 10, 21) {real, imag} */,
  {32'h3f2858b6, 32'h00000000} /* (26, 10, 20) {real, imag} */,
  {32'hbc7822b6, 32'h00000000} /* (26, 10, 19) {real, imag} */,
  {32'hbe89dbae, 32'h00000000} /* (26, 10, 18) {real, imag} */,
  {32'hbdc0035a, 32'h00000000} /* (26, 10, 17) {real, imag} */,
  {32'h3ec38c20, 32'h00000000} /* (26, 10, 16) {real, imag} */,
  {32'h3df187e0, 32'h00000000} /* (26, 10, 15) {real, imag} */,
  {32'hbef039fc, 32'h00000000} /* (26, 10, 14) {real, imag} */,
  {32'hbecaca3a, 32'h00000000} /* (26, 10, 13) {real, imag} */,
  {32'hbe7d2c9d, 32'h00000000} /* (26, 10, 12) {real, imag} */,
  {32'hbe9588f7, 32'h00000000} /* (26, 10, 11) {real, imag} */,
  {32'h3bffc650, 32'h00000000} /* (26, 10, 10) {real, imag} */,
  {32'h3e34cd54, 32'h00000000} /* (26, 10, 9) {real, imag} */,
  {32'h3ea31879, 32'h00000000} /* (26, 10, 8) {real, imag} */,
  {32'h3f488bf0, 32'h00000000} /* (26, 10, 7) {real, imag} */,
  {32'h3f107bdb, 32'h00000000} /* (26, 10, 6) {real, imag} */,
  {32'h3e39b963, 32'h00000000} /* (26, 10, 5) {real, imag} */,
  {32'h3ee27812, 32'h00000000} /* (26, 10, 4) {real, imag} */,
  {32'hbe68a206, 32'h00000000} /* (26, 10, 3) {real, imag} */,
  {32'hbcaabdc6, 32'h00000000} /* (26, 10, 2) {real, imag} */,
  {32'h3f1816ae, 32'h00000000} /* (26, 10, 1) {real, imag} */,
  {32'h3f164605, 32'h00000000} /* (26, 10, 0) {real, imag} */,
  {32'h3ed918f6, 32'h00000000} /* (26, 9, 31) {real, imag} */,
  {32'h3f2dc055, 32'h00000000} /* (26, 9, 30) {real, imag} */,
  {32'h3ea94f5e, 32'h00000000} /* (26, 9, 29) {real, imag} */,
  {32'h3e553ea5, 32'h00000000} /* (26, 9, 28) {real, imag} */,
  {32'h3d3ffd84, 32'h00000000} /* (26, 9, 27) {real, imag} */,
  {32'h3e8cd20a, 32'h00000000} /* (26, 9, 26) {real, imag} */,
  {32'h3e0b21fa, 32'h00000000} /* (26, 9, 25) {real, imag} */,
  {32'h3efbd016, 32'h00000000} /* (26, 9, 24) {real, imag} */,
  {32'h3dfe6718, 32'h00000000} /* (26, 9, 23) {real, imag} */,
  {32'h3b91432a, 32'h00000000} /* (26, 9, 22) {real, imag} */,
  {32'h3e0b051c, 32'h00000000} /* (26, 9, 21) {real, imag} */,
  {32'h3eb5c12c, 32'h00000000} /* (26, 9, 20) {real, imag} */,
  {32'hbe354d7b, 32'h00000000} /* (26, 9, 19) {real, imag} */,
  {32'hbeb0ba95, 32'h00000000} /* (26, 9, 18) {real, imag} */,
  {32'hbe9384fc, 32'h00000000} /* (26, 9, 17) {real, imag} */,
  {32'hbe533ea2, 32'h00000000} /* (26, 9, 16) {real, imag} */,
  {32'hbf0ad02b, 32'h00000000} /* (26, 9, 15) {real, imag} */,
  {32'hbee1c713, 32'h00000000} /* (26, 9, 14) {real, imag} */,
  {32'hbf4146d7, 32'h00000000} /* (26, 9, 13) {real, imag} */,
  {32'hbef6a689, 32'h00000000} /* (26, 9, 12) {real, imag} */,
  {32'hbd43e2ba, 32'h00000000} /* (26, 9, 11) {real, imag} */,
  {32'h3dec992a, 32'h00000000} /* (26, 9, 10) {real, imag} */,
  {32'h3e9bf0e2, 32'h00000000} /* (26, 9, 9) {real, imag} */,
  {32'h3ebde7d6, 32'h00000000} /* (26, 9, 8) {real, imag} */,
  {32'h3ee4205c, 32'h00000000} /* (26, 9, 7) {real, imag} */,
  {32'h3f14241e, 32'h00000000} /* (26, 9, 6) {real, imag} */,
  {32'h3d92b2f8, 32'h00000000} /* (26, 9, 5) {real, imag} */,
  {32'h3ea0febb, 32'h00000000} /* (26, 9, 4) {real, imag} */,
  {32'h3d4dae22, 32'h00000000} /* (26, 9, 3) {real, imag} */,
  {32'h3e8b52fd, 32'h00000000} /* (26, 9, 2) {real, imag} */,
  {32'h3f0f0a4b, 32'h00000000} /* (26, 9, 1) {real, imag} */,
  {32'h3e596094, 32'h00000000} /* (26, 9, 0) {real, imag} */,
  {32'h3eb7c1b7, 32'h00000000} /* (26, 8, 31) {real, imag} */,
  {32'h3ef05411, 32'h00000000} /* (26, 8, 30) {real, imag} */,
  {32'hbd198c44, 32'h00000000} /* (26, 8, 29) {real, imag} */,
  {32'hbbcf40ce, 32'h00000000} /* (26, 8, 28) {real, imag} */,
  {32'h3e3eaa9f, 32'h00000000} /* (26, 8, 27) {real, imag} */,
  {32'h3d1d3c8b, 32'h00000000} /* (26, 8, 26) {real, imag} */,
  {32'hbe3f52ad, 32'h00000000} /* (26, 8, 25) {real, imag} */,
  {32'h3d688807, 32'h00000000} /* (26, 8, 24) {real, imag} */,
  {32'h3e14dfcf, 32'h00000000} /* (26, 8, 23) {real, imag} */,
  {32'h3e747fc0, 32'h00000000} /* (26, 8, 22) {real, imag} */,
  {32'hbd74e1b4, 32'h00000000} /* (26, 8, 21) {real, imag} */,
  {32'h3aee57b8, 32'h00000000} /* (26, 8, 20) {real, imag} */,
  {32'hbe26855e, 32'h00000000} /* (26, 8, 19) {real, imag} */,
  {32'hbeff573e, 32'h00000000} /* (26, 8, 18) {real, imag} */,
  {32'hbee187bf, 32'h00000000} /* (26, 8, 17) {real, imag} */,
  {32'hbf13a864, 32'h00000000} /* (26, 8, 16) {real, imag} */,
  {32'hbf3b9c3d, 32'h00000000} /* (26, 8, 15) {real, imag} */,
  {32'hbf18095d, 32'h00000000} /* (26, 8, 14) {real, imag} */,
  {32'hbf22ae1a, 32'h00000000} /* (26, 8, 13) {real, imag} */,
  {32'hbf25f4b5, 32'h00000000} /* (26, 8, 12) {real, imag} */,
  {32'hbf15220e, 32'h00000000} /* (26, 8, 11) {real, imag} */,
  {32'h3a3f37c0, 32'h00000000} /* (26, 8, 10) {real, imag} */,
  {32'h3f1b593a, 32'h00000000} /* (26, 8, 9) {real, imag} */,
  {32'h3efb3c76, 32'h00000000} /* (26, 8, 8) {real, imag} */,
  {32'h3f091828, 32'h00000000} /* (26, 8, 7) {real, imag} */,
  {32'h3f1c11fc, 32'h00000000} /* (26, 8, 6) {real, imag} */,
  {32'h3e2368c0, 32'h00000000} /* (26, 8, 5) {real, imag} */,
  {32'h3f0b3a8b, 32'h00000000} /* (26, 8, 4) {real, imag} */,
  {32'h3eafabcb, 32'h00000000} /* (26, 8, 3) {real, imag} */,
  {32'h3e7dd7bc, 32'h00000000} /* (26, 8, 2) {real, imag} */,
  {32'h3e4e4aa9, 32'h00000000} /* (26, 8, 1) {real, imag} */,
  {32'hbe39bf67, 32'h00000000} /* (26, 8, 0) {real, imag} */,
  {32'h3e5e3b5a, 32'h00000000} /* (26, 7, 31) {real, imag} */,
  {32'h3e2c8650, 32'h00000000} /* (26, 7, 30) {real, imag} */,
  {32'hbf26cc67, 32'h00000000} /* (26, 7, 29) {real, imag} */,
  {32'hbf4dd480, 32'h00000000} /* (26, 7, 28) {real, imag} */,
  {32'h3cfc65fe, 32'h00000000} /* (26, 7, 27) {real, imag} */,
  {32'h3ea3be0a, 32'h00000000} /* (26, 7, 26) {real, imag} */,
  {32'h3db0a85b, 32'h00000000} /* (26, 7, 25) {real, imag} */,
  {32'h3e2cb3f4, 32'h00000000} /* (26, 7, 24) {real, imag} */,
  {32'h3f214f43, 32'h00000000} /* (26, 7, 23) {real, imag} */,
  {32'h3ee5236b, 32'h00000000} /* (26, 7, 22) {real, imag} */,
  {32'hbc19c88f, 32'h00000000} /* (26, 7, 21) {real, imag} */,
  {32'h3d8f0351, 32'h00000000} /* (26, 7, 20) {real, imag} */,
  {32'h3d8c77cc, 32'h00000000} /* (26, 7, 19) {real, imag} */,
  {32'hbea7c03a, 32'h00000000} /* (26, 7, 18) {real, imag} */,
  {32'hbf34b071, 32'h00000000} /* (26, 7, 17) {real, imag} */,
  {32'hbf31fe3b, 32'h00000000} /* (26, 7, 16) {real, imag} */,
  {32'hbe9318a3, 32'h00000000} /* (26, 7, 15) {real, imag} */,
  {32'hbe206231, 32'h00000000} /* (26, 7, 14) {real, imag} */,
  {32'hbeadcd41, 32'h00000000} /* (26, 7, 13) {real, imag} */,
  {32'hbe8d4394, 32'h00000000} /* (26, 7, 12) {real, imag} */,
  {32'hbf341f5d, 32'h00000000} /* (26, 7, 11) {real, imag} */,
  {32'hbd21d9b1, 32'h00000000} /* (26, 7, 10) {real, imag} */,
  {32'h3ecc5648, 32'h00000000} /* (26, 7, 9) {real, imag} */,
  {32'h3df233db, 32'h00000000} /* (26, 7, 8) {real, imag} */,
  {32'h3e979f1a, 32'h00000000} /* (26, 7, 7) {real, imag} */,
  {32'h3ec25c26, 32'h00000000} /* (26, 7, 6) {real, imag} */,
  {32'h3e82b5f4, 32'h00000000} /* (26, 7, 5) {real, imag} */,
  {32'h3f17332b, 32'h00000000} /* (26, 7, 4) {real, imag} */,
  {32'h3eae4c40, 32'h00000000} /* (26, 7, 3) {real, imag} */,
  {32'h3624be28, 32'h00000000} /* (26, 7, 2) {real, imag} */,
  {32'h3da38c4e, 32'h00000000} /* (26, 7, 1) {real, imag} */,
  {32'h3e65bf27, 32'h00000000} /* (26, 7, 0) {real, imag} */,
  {32'h3d873d14, 32'h00000000} /* (26, 6, 31) {real, imag} */,
  {32'hbdb0bd18, 32'h00000000} /* (26, 6, 30) {real, imag} */,
  {32'h3dca0d4e, 32'h00000000} /* (26, 6, 29) {real, imag} */,
  {32'hbe6cfa20, 32'h00000000} /* (26, 6, 28) {real, imag} */,
  {32'h3eae4e49, 32'h00000000} /* (26, 6, 27) {real, imag} */,
  {32'h3f488c67, 32'h00000000} /* (26, 6, 26) {real, imag} */,
  {32'h3f33af89, 32'h00000000} /* (26, 6, 25) {real, imag} */,
  {32'h3e340541, 32'h00000000} /* (26, 6, 24) {real, imag} */,
  {32'h3f097d1d, 32'h00000000} /* (26, 6, 23) {real, imag} */,
  {32'h3f273fc6, 32'h00000000} /* (26, 6, 22) {real, imag} */,
  {32'h3f136dba, 32'h00000000} /* (26, 6, 21) {real, imag} */,
  {32'h3d0e0fdf, 32'h00000000} /* (26, 6, 20) {real, imag} */,
  {32'hbd4fc53f, 32'h00000000} /* (26, 6, 19) {real, imag} */,
  {32'hbdf8bf24, 32'h00000000} /* (26, 6, 18) {real, imag} */,
  {32'hbe97f9a3, 32'h00000000} /* (26, 6, 17) {real, imag} */,
  {32'hbe8faa7c, 32'h00000000} /* (26, 6, 16) {real, imag} */,
  {32'hbd6f75db, 32'h00000000} /* (26, 6, 15) {real, imag} */,
  {32'hbd94bb46, 32'h00000000} /* (26, 6, 14) {real, imag} */,
  {32'hbf0e1482, 32'h00000000} /* (26, 6, 13) {real, imag} */,
  {32'hbc61b9a1, 32'h00000000} /* (26, 6, 12) {real, imag} */,
  {32'hbec0338c, 32'h00000000} /* (26, 6, 11) {real, imag} */,
  {32'h3e9f1446, 32'h00000000} /* (26, 6, 10) {real, imag} */,
  {32'h3f219aa1, 32'h00000000} /* (26, 6, 9) {real, imag} */,
  {32'h3f11f680, 32'h00000000} /* (26, 6, 8) {real, imag} */,
  {32'h3e76d4c4, 32'h00000000} /* (26, 6, 7) {real, imag} */,
  {32'hbe5f6d62, 32'h00000000} /* (26, 6, 6) {real, imag} */,
  {32'h3bda1960, 32'h00000000} /* (26, 6, 5) {real, imag} */,
  {32'h3e487810, 32'h00000000} /* (26, 6, 4) {real, imag} */,
  {32'hbd94f120, 32'h00000000} /* (26, 6, 3) {real, imag} */,
  {32'h3d72a48b, 32'h00000000} /* (26, 6, 2) {real, imag} */,
  {32'h3e316559, 32'h00000000} /* (26, 6, 1) {real, imag} */,
  {32'h3e85d151, 32'h00000000} /* (26, 6, 0) {real, imag} */,
  {32'hbe687268, 32'h00000000} /* (26, 5, 31) {real, imag} */,
  {32'hbe2fb4b9, 32'h00000000} /* (26, 5, 30) {real, imag} */,
  {32'h3ede2330, 32'h00000000} /* (26, 5, 29) {real, imag} */,
  {32'h3e99be87, 32'h00000000} /* (26, 5, 28) {real, imag} */,
  {32'h3ea5007a, 32'h00000000} /* (26, 5, 27) {real, imag} */,
  {32'h3ec5d1af, 32'h00000000} /* (26, 5, 26) {real, imag} */,
  {32'h3dd0dd62, 32'h00000000} /* (26, 5, 25) {real, imag} */,
  {32'h3d35a47b, 32'h00000000} /* (26, 5, 24) {real, imag} */,
  {32'h3e4a98ab, 32'h00000000} /* (26, 5, 23) {real, imag} */,
  {32'h3ec0fac2, 32'h00000000} /* (26, 5, 22) {real, imag} */,
  {32'h3f66fd3f, 32'h00000000} /* (26, 5, 21) {real, imag} */,
  {32'h3ed0c703, 32'h00000000} /* (26, 5, 20) {real, imag} */,
  {32'h3d88efdc, 32'h00000000} /* (26, 5, 19) {real, imag} */,
  {32'hbe7ab5f3, 32'h00000000} /* (26, 5, 18) {real, imag} */,
  {32'h3d7f4012, 32'h00000000} /* (26, 5, 17) {real, imag} */,
  {32'hbe737b92, 32'h00000000} /* (26, 5, 16) {real, imag} */,
  {32'hbed84282, 32'h00000000} /* (26, 5, 15) {real, imag} */,
  {32'hbf12754e, 32'h00000000} /* (26, 5, 14) {real, imag} */,
  {32'hbf35d732, 32'h00000000} /* (26, 5, 13) {real, imag} */,
  {32'hbe583c73, 32'h00000000} /* (26, 5, 12) {real, imag} */,
  {32'hbee7dee8, 32'h00000000} /* (26, 5, 11) {real, imag} */,
  {32'h3df4a0eb, 32'h00000000} /* (26, 5, 10) {real, imag} */,
  {32'h3f08865c, 32'h00000000} /* (26, 5, 9) {real, imag} */,
  {32'h3ee28e53, 32'h00000000} /* (26, 5, 8) {real, imag} */,
  {32'h3c851a29, 32'h00000000} /* (26, 5, 7) {real, imag} */,
  {32'hbf47b326, 32'h00000000} /* (26, 5, 6) {real, imag} */,
  {32'hbec9cfd0, 32'h00000000} /* (26, 5, 5) {real, imag} */,
  {32'hbe694181, 32'h00000000} /* (26, 5, 4) {real, imag} */,
  {32'hbe51ac2c, 32'h00000000} /* (26, 5, 3) {real, imag} */,
  {32'hbcb3469a, 32'h00000000} /* (26, 5, 2) {real, imag} */,
  {32'h3ecfce6a, 32'h00000000} /* (26, 5, 1) {real, imag} */,
  {32'h3e94f351, 32'h00000000} /* (26, 5, 0) {real, imag} */,
  {32'hbdb19b44, 32'h00000000} /* (26, 4, 31) {real, imag} */,
  {32'h3d37d8fe, 32'h00000000} /* (26, 4, 30) {real, imag} */,
  {32'hbd1a8588, 32'h00000000} /* (26, 4, 29) {real, imag} */,
  {32'h3b193992, 32'h00000000} /* (26, 4, 28) {real, imag} */,
  {32'hbd6dc83d, 32'h00000000} /* (26, 4, 27) {real, imag} */,
  {32'h3ea0f6fd, 32'h00000000} /* (26, 4, 26) {real, imag} */,
  {32'hbca6a5cf, 32'h00000000} /* (26, 4, 25) {real, imag} */,
  {32'hbe609822, 32'h00000000} /* (26, 4, 24) {real, imag} */,
  {32'hbb2b4149, 32'h00000000} /* (26, 4, 23) {real, imag} */,
  {32'h3f3a7a30, 32'h00000000} /* (26, 4, 22) {real, imag} */,
  {32'h3f966d61, 32'h00000000} /* (26, 4, 21) {real, imag} */,
  {32'h3f04ed77, 32'h00000000} /* (26, 4, 20) {real, imag} */,
  {32'hbdc15419, 32'h00000000} /* (26, 4, 19) {real, imag} */,
  {32'hbceb59a6, 32'h00000000} /* (26, 4, 18) {real, imag} */,
  {32'h3b0d4d78, 32'h00000000} /* (26, 4, 17) {real, imag} */,
  {32'h3e44c0e3, 32'h00000000} /* (26, 4, 16) {real, imag} */,
  {32'h3e03945d, 32'h00000000} /* (26, 4, 15) {real, imag} */,
  {32'hbee2a2a2, 32'h00000000} /* (26, 4, 14) {real, imag} */,
  {32'hbe585d26, 32'h00000000} /* (26, 4, 13) {real, imag} */,
  {32'h3d18d5f4, 32'h00000000} /* (26, 4, 12) {real, imag} */,
  {32'h3ddb4b89, 32'h00000000} /* (26, 4, 11) {real, imag} */,
  {32'hbe103ad4, 32'h00000000} /* (26, 4, 10) {real, imag} */,
  {32'hbe86c71a, 32'h00000000} /* (26, 4, 9) {real, imag} */,
  {32'h3e31e5b5, 32'h00000000} /* (26, 4, 8) {real, imag} */,
  {32'h3da6c45c, 32'h00000000} /* (26, 4, 7) {real, imag} */,
  {32'hbe99f416, 32'h00000000} /* (26, 4, 6) {real, imag} */,
  {32'h3f639757, 32'h00000000} /* (26, 4, 5) {real, imag} */,
  {32'h3f276996, 32'h00000000} /* (26, 4, 4) {real, imag} */,
  {32'h3e9c6f19, 32'h00000000} /* (26, 4, 3) {real, imag} */,
  {32'h3f042864, 32'h00000000} /* (26, 4, 2) {real, imag} */,
  {32'h3ebfa3c0, 32'h00000000} /* (26, 4, 1) {real, imag} */,
  {32'h3e310a32, 32'h00000000} /* (26, 4, 0) {real, imag} */,
  {32'h3e1b4315, 32'h00000000} /* (26, 3, 31) {real, imag} */,
  {32'h3f4c7484, 32'h00000000} /* (26, 3, 30) {real, imag} */,
  {32'hbd8c471b, 32'h00000000} /* (26, 3, 29) {real, imag} */,
  {32'h3d13379e, 32'h00000000} /* (26, 3, 28) {real, imag} */,
  {32'h3949e02e, 32'h00000000} /* (26, 3, 27) {real, imag} */,
  {32'h3e9782a5, 32'h00000000} /* (26, 3, 26) {real, imag} */,
  {32'h3e59a6d3, 32'h00000000} /* (26, 3, 25) {real, imag} */,
  {32'hbddde9ac, 32'h00000000} /* (26, 3, 24) {real, imag} */,
  {32'hbe113f71, 32'h00000000} /* (26, 3, 23) {real, imag} */,
  {32'h3f0879b8, 32'h00000000} /* (26, 3, 22) {real, imag} */,
  {32'h3f0ad9dd, 32'h00000000} /* (26, 3, 21) {real, imag} */,
  {32'h3e81b2c0, 32'h00000000} /* (26, 3, 20) {real, imag} */,
  {32'h3ee5356b, 32'h00000000} /* (26, 3, 19) {real, imag} */,
  {32'h3f3fe603, 32'h00000000} /* (26, 3, 18) {real, imag} */,
  {32'h3e11d949, 32'h00000000} /* (26, 3, 17) {real, imag} */,
  {32'h3e7f73b2, 32'h00000000} /* (26, 3, 16) {real, imag} */,
  {32'h3e9bb06e, 32'h00000000} /* (26, 3, 15) {real, imag} */,
  {32'hbd08acfd, 32'h00000000} /* (26, 3, 14) {real, imag} */,
  {32'hbe89d4ae, 32'h00000000} /* (26, 3, 13) {real, imag} */,
  {32'h3c9f8eb5, 32'h00000000} /* (26, 3, 12) {real, imag} */,
  {32'h3ee80fa2, 32'h00000000} /* (26, 3, 11) {real, imag} */,
  {32'hbe73a8b2, 32'h00000000} /* (26, 3, 10) {real, imag} */,
  {32'hbee8ef35, 32'h00000000} /* (26, 3, 9) {real, imag} */,
  {32'h3df991e9, 32'h00000000} /* (26, 3, 8) {real, imag} */,
  {32'h3f2997ea, 32'h00000000} /* (26, 3, 7) {real, imag} */,
  {32'h3d488e97, 32'h00000000} /* (26, 3, 6) {real, imag} */,
  {32'h3f4d5982, 32'h00000000} /* (26, 3, 5) {real, imag} */,
  {32'h3ed6cfaa, 32'h00000000} /* (26, 3, 4) {real, imag} */,
  {32'h3f0199e0, 32'h00000000} /* (26, 3, 3) {real, imag} */,
  {32'h3f7805b2, 32'h00000000} /* (26, 3, 2) {real, imag} */,
  {32'h3ea2baf1, 32'h00000000} /* (26, 3, 1) {real, imag} */,
  {32'h3d58e4da, 32'h00000000} /* (26, 3, 0) {real, imag} */,
  {32'h3ec86869, 32'h00000000} /* (26, 2, 31) {real, imag} */,
  {32'h3f6b4eee, 32'h00000000} /* (26, 2, 30) {real, imag} */,
  {32'h3e17da0f, 32'h00000000} /* (26, 2, 29) {real, imag} */,
  {32'hbe27370d, 32'h00000000} /* (26, 2, 28) {real, imag} */,
  {32'h3dabe515, 32'h00000000} /* (26, 2, 27) {real, imag} */,
  {32'h3ea85fb2, 32'h00000000} /* (26, 2, 26) {real, imag} */,
  {32'h3efa6a7e, 32'h00000000} /* (26, 2, 25) {real, imag} */,
  {32'h3f28aab6, 32'h00000000} /* (26, 2, 24) {real, imag} */,
  {32'h3e39b067, 32'h00000000} /* (26, 2, 23) {real, imag} */,
  {32'h3e95d08c, 32'h00000000} /* (26, 2, 22) {real, imag} */,
  {32'h3efe47a9, 32'h00000000} /* (26, 2, 21) {real, imag} */,
  {32'h3e8132b1, 32'h00000000} /* (26, 2, 20) {real, imag} */,
  {32'h3ec818c1, 32'h00000000} /* (26, 2, 19) {real, imag} */,
  {32'h3ea2c415, 32'h00000000} /* (26, 2, 18) {real, imag} */,
  {32'h3f58ed93, 32'h00000000} /* (26, 2, 17) {real, imag} */,
  {32'h3f4331f1, 32'h00000000} /* (26, 2, 16) {real, imag} */,
  {32'h3eaa41a2, 32'h00000000} /* (26, 2, 15) {real, imag} */,
  {32'h3da0bc5b, 32'h00000000} /* (26, 2, 14) {real, imag} */,
  {32'hbe25ef9d, 32'h00000000} /* (26, 2, 13) {real, imag} */,
  {32'hbe71023d, 32'h00000000} /* (26, 2, 12) {real, imag} */,
  {32'hbea2c799, 32'h00000000} /* (26, 2, 11) {real, imag} */,
  {32'hbe83f7e6, 32'h00000000} /* (26, 2, 10) {real, imag} */,
  {32'hbdd655b4, 32'h00000000} /* (26, 2, 9) {real, imag} */,
  {32'hbea41bbd, 32'h00000000} /* (26, 2, 8) {real, imag} */,
  {32'h3e84cf09, 32'h00000000} /* (26, 2, 7) {real, imag} */,
  {32'hbe81bd9b, 32'h00000000} /* (26, 2, 6) {real, imag} */,
  {32'hbe7416c8, 32'h00000000} /* (26, 2, 5) {real, imag} */,
  {32'h3d21d2b1, 32'h00000000} /* (26, 2, 4) {real, imag} */,
  {32'h3efa66ca, 32'h00000000} /* (26, 2, 3) {real, imag} */,
  {32'h3f3cd25d, 32'h00000000} /* (26, 2, 2) {real, imag} */,
  {32'h3e8a4900, 32'h00000000} /* (26, 2, 1) {real, imag} */,
  {32'h3e18449d, 32'h00000000} /* (26, 2, 0) {real, imag} */,
  {32'h3e56c831, 32'h00000000} /* (26, 1, 31) {real, imag} */,
  {32'h3efd8b6b, 32'h00000000} /* (26, 1, 30) {real, imag} */,
  {32'h3e217db9, 32'h00000000} /* (26, 1, 29) {real, imag} */,
  {32'hbe543fdd, 32'h00000000} /* (26, 1, 28) {real, imag} */,
  {32'h3ed66f51, 32'h00000000} /* (26, 1, 27) {real, imag} */,
  {32'h3eca4f59, 32'h00000000} /* (26, 1, 26) {real, imag} */,
  {32'h3f194682, 32'h00000000} /* (26, 1, 25) {real, imag} */,
  {32'h3f4c9af2, 32'h00000000} /* (26, 1, 24) {real, imag} */,
  {32'h3e9a7811, 32'h00000000} /* (26, 1, 23) {real, imag} */,
  {32'h3e0e7c55, 32'h00000000} /* (26, 1, 22) {real, imag} */,
  {32'hbde69f10, 32'h00000000} /* (26, 1, 21) {real, imag} */,
  {32'h3f036a11, 32'h00000000} /* (26, 1, 20) {real, imag} */,
  {32'h3ee0c448, 32'h00000000} /* (26, 1, 19) {real, imag} */,
  {32'h3e87eeb7, 32'h00000000} /* (26, 1, 18) {real, imag} */,
  {32'h3f61b5bb, 32'h00000000} /* (26, 1, 17) {real, imag} */,
  {32'h3ed32b08, 32'h00000000} /* (26, 1, 16) {real, imag} */,
  {32'hbea9e6d6, 32'h00000000} /* (26, 1, 15) {real, imag} */,
  {32'hbec0e993, 32'h00000000} /* (26, 1, 14) {real, imag} */,
  {32'hbe7db8c9, 32'h00000000} /* (26, 1, 13) {real, imag} */,
  {32'hbe30931d, 32'h00000000} /* (26, 1, 12) {real, imag} */,
  {32'hbd40cc88, 32'h00000000} /* (26, 1, 11) {real, imag} */,
  {32'hbed07487, 32'h00000000} /* (26, 1, 10) {real, imag} */,
  {32'hbec91b47, 32'h00000000} /* (26, 1, 9) {real, imag} */,
  {32'hbe38f0b2, 32'h00000000} /* (26, 1, 8) {real, imag} */,
  {32'hbeba9a46, 32'h00000000} /* (26, 1, 7) {real, imag} */,
  {32'hbf69f179, 32'h00000000} /* (26, 1, 6) {real, imag} */,
  {32'hbe3f85e2, 32'h00000000} /* (26, 1, 5) {real, imag} */,
  {32'h3f385ca5, 32'h00000000} /* (26, 1, 4) {real, imag} */,
  {32'h3f25b273, 32'h00000000} /* (26, 1, 3) {real, imag} */,
  {32'h3ec8ee5a, 32'h00000000} /* (26, 1, 2) {real, imag} */,
  {32'h3da59c86, 32'h00000000} /* (26, 1, 1) {real, imag} */,
  {32'h3dd86539, 32'h00000000} /* (26, 1, 0) {real, imag} */,
  {32'h3d8661e8, 32'h00000000} /* (26, 0, 31) {real, imag} */,
  {32'h3ea3ec8b, 32'h00000000} /* (26, 0, 30) {real, imag} */,
  {32'h3e5600fc, 32'h00000000} /* (26, 0, 29) {real, imag} */,
  {32'hbd015b80, 32'h00000000} /* (26, 0, 28) {real, imag} */,
  {32'h3e2d70b0, 32'h00000000} /* (26, 0, 27) {real, imag} */,
  {32'h3e0bd544, 32'h00000000} /* (26, 0, 26) {real, imag} */,
  {32'h3e20f03e, 32'h00000000} /* (26, 0, 25) {real, imag} */,
  {32'h3e5d5c96, 32'h00000000} /* (26, 0, 24) {real, imag} */,
  {32'h3e332f35, 32'h00000000} /* (26, 0, 23) {real, imag} */,
  {32'h3dbd517c, 32'h00000000} /* (26, 0, 22) {real, imag} */,
  {32'hbb7a8440, 32'h00000000} /* (26, 0, 21) {real, imag} */,
  {32'h3f2a175e, 32'h00000000} /* (26, 0, 20) {real, imag} */,
  {32'h3f30e63c, 32'h00000000} /* (26, 0, 19) {real, imag} */,
  {32'h3f19914e, 32'h00000000} /* (26, 0, 18) {real, imag} */,
  {32'h3efa27ff, 32'h00000000} /* (26, 0, 17) {real, imag} */,
  {32'hbe39d8ed, 32'h00000000} /* (26, 0, 16) {real, imag} */,
  {32'hbe9e6738, 32'h00000000} /* (26, 0, 15) {real, imag} */,
  {32'hbe28e054, 32'h00000000} /* (26, 0, 14) {real, imag} */,
  {32'hbe00f7ba, 32'h00000000} /* (26, 0, 13) {real, imag} */,
  {32'hbcc70e81, 32'h00000000} /* (26, 0, 12) {real, imag} */,
  {32'h3d8a2947, 32'h00000000} /* (26, 0, 11) {real, imag} */,
  {32'hbe9e6c56, 32'h00000000} /* (26, 0, 10) {real, imag} */,
  {32'hbe50b1ac, 32'h00000000} /* (26, 0, 9) {real, imag} */,
  {32'hbd48b5ef, 32'h00000000} /* (26, 0, 8) {real, imag} */,
  {32'hbf2748a2, 32'h00000000} /* (26, 0, 7) {real, imag} */,
  {32'hbf28b9b2, 32'h00000000} /* (26, 0, 6) {real, imag} */,
  {32'h3d2a9ad3, 32'h00000000} /* (26, 0, 5) {real, imag} */,
  {32'h3ebe5d73, 32'h00000000} /* (26, 0, 4) {real, imag} */,
  {32'h3e37da84, 32'h00000000} /* (26, 0, 3) {real, imag} */,
  {32'hbdf70fe1, 32'h00000000} /* (26, 0, 2) {real, imag} */,
  {32'hbdfe6f72, 32'h00000000} /* (26, 0, 1) {real, imag} */,
  {32'h3e5ccfd8, 32'h00000000} /* (26, 0, 0) {real, imag} */,
  {32'hbe1be529, 32'h00000000} /* (25, 31, 31) {real, imag} */,
  {32'hbee5d484, 32'h00000000} /* (25, 31, 30) {real, imag} */,
  {32'hbecb55dc, 32'h00000000} /* (25, 31, 29) {real, imag} */,
  {32'hbed8bc51, 32'h00000000} /* (25, 31, 28) {real, imag} */,
  {32'hbe6ac0f9, 32'h00000000} /* (25, 31, 27) {real, imag} */,
  {32'hbe5f04e0, 32'h00000000} /* (25, 31, 26) {real, imag} */,
  {32'hbeaf2e4f, 32'h00000000} /* (25, 31, 25) {real, imag} */,
  {32'hbed209b9, 32'h00000000} /* (25, 31, 24) {real, imag} */,
  {32'hbf1364b8, 32'h00000000} /* (25, 31, 23) {real, imag} */,
  {32'hbed44b19, 32'h00000000} /* (25, 31, 22) {real, imag} */,
  {32'hbe35662a, 32'h00000000} /* (25, 31, 21) {real, imag} */,
  {32'h3ebfa7b9, 32'h00000000} /* (25, 31, 20) {real, imag} */,
  {32'h3f270725, 32'h00000000} /* (25, 31, 19) {real, imag} */,
  {32'h3f30bac5, 32'h00000000} /* (25, 31, 18) {real, imag} */,
  {32'h3e854c39, 32'h00000000} /* (25, 31, 17) {real, imag} */,
  {32'h3e157e2d, 32'h00000000} /* (25, 31, 16) {real, imag} */,
  {32'h3e960e32, 32'h00000000} /* (25, 31, 15) {real, imag} */,
  {32'h3ebbfe30, 32'h00000000} /* (25, 31, 14) {real, imag} */,
  {32'h3f3d1470, 32'h00000000} /* (25, 31, 13) {real, imag} */,
  {32'h3ee46e18, 32'h00000000} /* (25, 31, 12) {real, imag} */,
  {32'h3e365247, 32'h00000000} /* (25, 31, 11) {real, imag} */,
  {32'hbe32d497, 32'h00000000} /* (25, 31, 10) {real, imag} */,
  {32'hbeb523ef, 32'h00000000} /* (25, 31, 9) {real, imag} */,
  {32'hbec0b96e, 32'h00000000} /* (25, 31, 8) {real, imag} */,
  {32'hbecbe041, 32'h00000000} /* (25, 31, 7) {real, imag} */,
  {32'hbe9d486e, 32'h00000000} /* (25, 31, 6) {real, imag} */,
  {32'hbf0b7b70, 32'h00000000} /* (25, 31, 5) {real, imag} */,
  {32'hbf0e9b87, 32'h00000000} /* (25, 31, 4) {real, imag} */,
  {32'hbee17aed, 32'h00000000} /* (25, 31, 3) {real, imag} */,
  {32'hbecca6c1, 32'h00000000} /* (25, 31, 2) {real, imag} */,
  {32'hbf64011f, 32'h00000000} /* (25, 31, 1) {real, imag} */,
  {32'hbe393486, 32'h00000000} /* (25, 31, 0) {real, imag} */,
  {32'hbdc03ea4, 32'h00000000} /* (25, 30, 31) {real, imag} */,
  {32'hbee6eacf, 32'h00000000} /* (25, 30, 30) {real, imag} */,
  {32'hbf153306, 32'h00000000} /* (25, 30, 29) {real, imag} */,
  {32'hbf060450, 32'h00000000} /* (25, 30, 28) {real, imag} */,
  {32'hbe8ab4e0, 32'h00000000} /* (25, 30, 27) {real, imag} */,
  {32'hbf1d16db, 32'h00000000} /* (25, 30, 26) {real, imag} */,
  {32'hbf53d48b, 32'h00000000} /* (25, 30, 25) {real, imag} */,
  {32'hbf815ed0, 32'h00000000} /* (25, 30, 24) {real, imag} */,
  {32'hbf4a2de2, 32'h00000000} /* (25, 30, 23) {real, imag} */,
  {32'hbedc6c0e, 32'h00000000} /* (25, 30, 22) {real, imag} */,
  {32'hbb2f6280, 32'h00000000} /* (25, 30, 21) {real, imag} */,
  {32'h3f83d721, 32'h00000000} /* (25, 30, 20) {real, imag} */,
  {32'h3f52b8df, 32'h00000000} /* (25, 30, 19) {real, imag} */,
  {32'h3f92ce2a, 32'h00000000} /* (25, 30, 18) {real, imag} */,
  {32'h3f4bb7ac, 32'h00000000} /* (25, 30, 17) {real, imag} */,
  {32'h3f7493d8, 32'h00000000} /* (25, 30, 16) {real, imag} */,
  {32'h3f8c0fcf, 32'h00000000} /* (25, 30, 15) {real, imag} */,
  {32'h3f6cf05e, 32'h00000000} /* (25, 30, 14) {real, imag} */,
  {32'h3f8cff1c, 32'h00000000} /* (25, 30, 13) {real, imag} */,
  {32'h3f33f5e3, 32'h00000000} /* (25, 30, 12) {real, imag} */,
  {32'h3ef0a918, 32'h00000000} /* (25, 30, 11) {real, imag} */,
  {32'hbe64eda7, 32'h00000000} /* (25, 30, 10) {real, imag} */,
  {32'hbf1199ff, 32'h00000000} /* (25, 30, 9) {real, imag} */,
  {32'hbf554eab, 32'h00000000} /* (25, 30, 8) {real, imag} */,
  {32'hbf734736, 32'h00000000} /* (25, 30, 7) {real, imag} */,
  {32'hbf456026, 32'h00000000} /* (25, 30, 6) {real, imag} */,
  {32'hbf372ddc, 32'h00000000} /* (25, 30, 5) {real, imag} */,
  {32'hbf24caa1, 32'h00000000} /* (25, 30, 4) {real, imag} */,
  {32'hbf3ec897, 32'h00000000} /* (25, 30, 3) {real, imag} */,
  {32'hbf065183, 32'h00000000} /* (25, 30, 2) {real, imag} */,
  {32'hbf61ad90, 32'h00000000} /* (25, 30, 1) {real, imag} */,
  {32'hbea133cd, 32'h00000000} /* (25, 30, 0) {real, imag} */,
  {32'h3d48fb43, 32'h00000000} /* (25, 29, 31) {real, imag} */,
  {32'hbf24de98, 32'h00000000} /* (25, 29, 30) {real, imag} */,
  {32'hbf443bf4, 32'h00000000} /* (25, 29, 29) {real, imag} */,
  {32'hbf075803, 32'h00000000} /* (25, 29, 28) {real, imag} */,
  {32'hbf8304bd, 32'h00000000} /* (25, 29, 27) {real, imag} */,
  {32'hbfbb5761, 32'h00000000} /* (25, 29, 26) {real, imag} */,
  {32'hbfa8c158, 32'h00000000} /* (25, 29, 25) {real, imag} */,
  {32'hbf5374b3, 32'h00000000} /* (25, 29, 24) {real, imag} */,
  {32'hbeef06cf, 32'h00000000} /* (25, 29, 23) {real, imag} */,
  {32'hbf3bc400, 32'h00000000} /* (25, 29, 22) {real, imag} */,
  {32'hbf4ac09c, 32'h00000000} /* (25, 29, 21) {real, imag} */,
  {32'h3f56bf68, 32'h00000000} /* (25, 29, 20) {real, imag} */,
  {32'h3f2ae977, 32'h00000000} /* (25, 29, 19) {real, imag} */,
  {32'h3f65e8a1, 32'h00000000} /* (25, 29, 18) {real, imag} */,
  {32'h3f177068, 32'h00000000} /* (25, 29, 17) {real, imag} */,
  {32'h3ea8a8ab, 32'h00000000} /* (25, 29, 16) {real, imag} */,
  {32'h3f2719ae, 32'h00000000} /* (25, 29, 15) {real, imag} */,
  {32'h3f49c2e4, 32'h00000000} /* (25, 29, 14) {real, imag} */,
  {32'h3ee073e0, 32'h00000000} /* (25, 29, 13) {real, imag} */,
  {32'h3f139303, 32'h00000000} /* (25, 29, 12) {real, imag} */,
  {32'h3ed9f12b, 32'h00000000} /* (25, 29, 11) {real, imag} */,
  {32'hbeb027aa, 32'h00000000} /* (25, 29, 10) {real, imag} */,
  {32'hbebdd2f7, 32'h00000000} /* (25, 29, 9) {real, imag} */,
  {32'hbf6e55e1, 32'h00000000} /* (25, 29, 8) {real, imag} */,
  {32'hbf9b345c, 32'h00000000} /* (25, 29, 7) {real, imag} */,
  {32'hbec26aa8, 32'h00000000} /* (25, 29, 6) {real, imag} */,
  {32'h3d5da58a, 32'h00000000} /* (25, 29, 5) {real, imag} */,
  {32'h3d564efe, 32'h00000000} /* (25, 29, 4) {real, imag} */,
  {32'hbf4dd4c6, 32'h00000000} /* (25, 29, 3) {real, imag} */,
  {32'hbf721257, 32'h00000000} /* (25, 29, 2) {real, imag} */,
  {32'hbf343c8d, 32'h00000000} /* (25, 29, 1) {real, imag} */,
  {32'h3c80e4e6, 32'h00000000} /* (25, 29, 0) {real, imag} */,
  {32'hbe06e687, 32'h00000000} /* (25, 28, 31) {real, imag} */,
  {32'hbf7cf5e0, 32'h00000000} /* (25, 28, 30) {real, imag} */,
  {32'hbf83c46a, 32'h00000000} /* (25, 28, 29) {real, imag} */,
  {32'hbf28f146, 32'h00000000} /* (25, 28, 28) {real, imag} */,
  {32'hbf957df6, 32'h00000000} /* (25, 28, 27) {real, imag} */,
  {32'hbfbc7516, 32'h00000000} /* (25, 28, 26) {real, imag} */,
  {32'hbfa6d464, 32'h00000000} /* (25, 28, 25) {real, imag} */,
  {32'hbf4db9ff, 32'h00000000} /* (25, 28, 24) {real, imag} */,
  {32'hbf464fc5, 32'h00000000} /* (25, 28, 23) {real, imag} */,
  {32'hbf894c13, 32'h00000000} /* (25, 28, 22) {real, imag} */,
  {32'hbfab57b2, 32'h00000000} /* (25, 28, 21) {real, imag} */,
  {32'h3e475fe4, 32'h00000000} /* (25, 28, 20) {real, imag} */,
  {32'h3f3c07ca, 32'h00000000} /* (25, 28, 19) {real, imag} */,
  {32'h3fc6630c, 32'h00000000} /* (25, 28, 18) {real, imag} */,
  {32'h3f837f09, 32'h00000000} /* (25, 28, 17) {real, imag} */,
  {32'h3ed376b5, 32'h00000000} /* (25, 28, 16) {real, imag} */,
  {32'h3e8e6758, 32'h00000000} /* (25, 28, 15) {real, imag} */,
  {32'h3ef81bfc, 32'h00000000} /* (25, 28, 14) {real, imag} */,
  {32'h3e6035d2, 32'h00000000} /* (25, 28, 13) {real, imag} */,
  {32'h3f5e086f, 32'h00000000} /* (25, 28, 12) {real, imag} */,
  {32'h3f56df69, 32'h00000000} /* (25, 28, 11) {real, imag} */,
  {32'hbeb87683, 32'h00000000} /* (25, 28, 10) {real, imag} */,
  {32'hbf56465c, 32'h00000000} /* (25, 28, 9) {real, imag} */,
  {32'hbf48258e, 32'h00000000} /* (25, 28, 8) {real, imag} */,
  {32'hbf44e63e, 32'h00000000} /* (25, 28, 7) {real, imag} */,
  {32'hbedc6b68, 32'h00000000} /* (25, 28, 6) {real, imag} */,
  {32'hbf535f09, 32'h00000000} /* (25, 28, 5) {real, imag} */,
  {32'hbf572b26, 32'h00000000} /* (25, 28, 4) {real, imag} */,
  {32'hbf8b5379, 32'h00000000} /* (25, 28, 3) {real, imag} */,
  {32'hbf63b54a, 32'h00000000} /* (25, 28, 2) {real, imag} */,
  {32'hbf83e7dd, 32'h00000000} /* (25, 28, 1) {real, imag} */,
  {32'hbecf4a2b, 32'h00000000} /* (25, 28, 0) {real, imag} */,
  {32'h3da18179, 32'h00000000} /* (25, 27, 31) {real, imag} */,
  {32'hbeee3a25, 32'h00000000} /* (25, 27, 30) {real, imag} */,
  {32'hbf48fe56, 32'h00000000} /* (25, 27, 29) {real, imag} */,
  {32'hbf363b3c, 32'h00000000} /* (25, 27, 28) {real, imag} */,
  {32'hbf8cc8bf, 32'h00000000} /* (25, 27, 27) {real, imag} */,
  {32'hbfbe764f, 32'h00000000} /* (25, 27, 26) {real, imag} */,
  {32'hbfb98bbf, 32'h00000000} /* (25, 27, 25) {real, imag} */,
  {32'hbf839cfa, 32'h00000000} /* (25, 27, 24) {real, imag} */,
  {32'hbf09922f, 32'h00000000} /* (25, 27, 23) {real, imag} */,
  {32'hbf4bd447, 32'h00000000} /* (25, 27, 22) {real, imag} */,
  {32'hbf7dc601, 32'h00000000} /* (25, 27, 21) {real, imag} */,
  {32'h3e662808, 32'h00000000} /* (25, 27, 20) {real, imag} */,
  {32'h3f7d1055, 32'h00000000} /* (25, 27, 19) {real, imag} */,
  {32'h3fbdd4de, 32'h00000000} /* (25, 27, 18) {real, imag} */,
  {32'h3f5d3920, 32'h00000000} /* (25, 27, 17) {real, imag} */,
  {32'h3f5e4ccc, 32'h00000000} /* (25, 27, 16) {real, imag} */,
  {32'h3f0842a7, 32'h00000000} /* (25, 27, 15) {real, imag} */,
  {32'h3e435d61, 32'h00000000} /* (25, 27, 14) {real, imag} */,
  {32'h3e997351, 32'h00000000} /* (25, 27, 13) {real, imag} */,
  {32'h3f1680a2, 32'h00000000} /* (25, 27, 12) {real, imag} */,
  {32'h3f711c0a, 32'h00000000} /* (25, 27, 11) {real, imag} */,
  {32'hbea260e0, 32'h00000000} /* (25, 27, 10) {real, imag} */,
  {32'hbfe2c7fa, 32'h00000000} /* (25, 27, 9) {real, imag} */,
  {32'hbf61689e, 32'h00000000} /* (25, 27, 8) {real, imag} */,
  {32'hbee134ce, 32'h00000000} /* (25, 27, 7) {real, imag} */,
  {32'hbf1eca92, 32'h00000000} /* (25, 27, 6) {real, imag} */,
  {32'hbf8d5241, 32'h00000000} /* (25, 27, 5) {real, imag} */,
  {32'hbfb88f9f, 32'h00000000} /* (25, 27, 4) {real, imag} */,
  {32'hbfbc8a9c, 32'h00000000} /* (25, 27, 3) {real, imag} */,
  {32'hbf4c7b17, 32'h00000000} /* (25, 27, 2) {real, imag} */,
  {32'hbf348198, 32'h00000000} /* (25, 27, 1) {real, imag} */,
  {32'hbe94b9e9, 32'h00000000} /* (25, 27, 0) {real, imag} */,
  {32'hbde39db6, 32'h00000000} /* (25, 26, 31) {real, imag} */,
  {32'hbf3f338e, 32'h00000000} /* (25, 26, 30) {real, imag} */,
  {32'hbfb0d86a, 32'h00000000} /* (25, 26, 29) {real, imag} */,
  {32'hbf8b80d6, 32'h00000000} /* (25, 26, 28) {real, imag} */,
  {32'hbf72add3, 32'h00000000} /* (25, 26, 27) {real, imag} */,
  {32'hbf78c786, 32'h00000000} /* (25, 26, 26) {real, imag} */,
  {32'hbf86059e, 32'h00000000} /* (25, 26, 25) {real, imag} */,
  {32'hbf1e3311, 32'h00000000} /* (25, 26, 24) {real, imag} */,
  {32'hbe810470, 32'h00000000} /* (25, 26, 23) {real, imag} */,
  {32'hbeda187c, 32'h00000000} /* (25, 26, 22) {real, imag} */,
  {32'hbf3af1d5, 32'h00000000} /* (25, 26, 21) {real, imag} */,
  {32'h3e93192b, 32'h00000000} /* (25, 26, 20) {real, imag} */,
  {32'h3f502244, 32'h00000000} /* (25, 26, 19) {real, imag} */,
  {32'h3f8e2892, 32'h00000000} /* (25, 26, 18) {real, imag} */,
  {32'h3f0ceef2, 32'h00000000} /* (25, 26, 17) {real, imag} */,
  {32'h3f62d9e8, 32'h00000000} /* (25, 26, 16) {real, imag} */,
  {32'h3f104c1a, 32'h00000000} /* (25, 26, 15) {real, imag} */,
  {32'h3ec4fd5d, 32'h00000000} /* (25, 26, 14) {real, imag} */,
  {32'h3eb86235, 32'h00000000} /* (25, 26, 13) {real, imag} */,
  {32'h3eac2788, 32'h00000000} /* (25, 26, 12) {real, imag} */,
  {32'h3ebff461, 32'h00000000} /* (25, 26, 11) {real, imag} */,
  {32'hbefeece6, 32'h00000000} /* (25, 26, 10) {real, imag} */,
  {32'hbfb7ca30, 32'h00000000} /* (25, 26, 9) {real, imag} */,
  {32'hbf7ef434, 32'h00000000} /* (25, 26, 8) {real, imag} */,
  {32'hbf31955d, 32'h00000000} /* (25, 26, 7) {real, imag} */,
  {32'hbf100e69, 32'h00000000} /* (25, 26, 6) {real, imag} */,
  {32'hbf1ee635, 32'h00000000} /* (25, 26, 5) {real, imag} */,
  {32'hbee4f367, 32'h00000000} /* (25, 26, 4) {real, imag} */,
  {32'hbf12f6be, 32'h00000000} /* (25, 26, 3) {real, imag} */,
  {32'hbf0487e9, 32'h00000000} /* (25, 26, 2) {real, imag} */,
  {32'hbf11015b, 32'h00000000} /* (25, 26, 1) {real, imag} */,
  {32'hbe9a965e, 32'h00000000} /* (25, 26, 0) {real, imag} */,
  {32'hbf24b36f, 32'h00000000} /* (25, 25, 31) {real, imag} */,
  {32'hbf9f1f8e, 32'h00000000} /* (25, 25, 30) {real, imag} */,
  {32'hbfa2b36f, 32'h00000000} /* (25, 25, 29) {real, imag} */,
  {32'hbf4f49b4, 32'h00000000} /* (25, 25, 28) {real, imag} */,
  {32'hbf81f4f4, 32'h00000000} /* (25, 25, 27) {real, imag} */,
  {32'hbf4aa05a, 32'h00000000} /* (25, 25, 26) {real, imag} */,
  {32'hbf33e5da, 32'h00000000} /* (25, 25, 25) {real, imag} */,
  {32'hbf3fa94c, 32'h00000000} /* (25, 25, 24) {real, imag} */,
  {32'hbf05a0c2, 32'h00000000} /* (25, 25, 23) {real, imag} */,
  {32'hbee85980, 32'h00000000} /* (25, 25, 22) {real, imag} */,
  {32'h3e7f24ab, 32'h00000000} /* (25, 25, 21) {real, imag} */,
  {32'h3fa4be12, 32'h00000000} /* (25, 25, 20) {real, imag} */,
  {32'h3f28e23d, 32'h00000000} /* (25, 25, 19) {real, imag} */,
  {32'h3f3467fc, 32'h00000000} /* (25, 25, 18) {real, imag} */,
  {32'h3ea7e3fa, 32'h00000000} /* (25, 25, 17) {real, imag} */,
  {32'h3f1c761f, 32'h00000000} /* (25, 25, 16) {real, imag} */,
  {32'h3ef6236f, 32'h00000000} /* (25, 25, 15) {real, imag} */,
  {32'h3f818161, 32'h00000000} /* (25, 25, 14) {real, imag} */,
  {32'h3f8edb71, 32'h00000000} /* (25, 25, 13) {real, imag} */,
  {32'h3f17993d, 32'h00000000} /* (25, 25, 12) {real, imag} */,
  {32'hbdd2bd9a, 32'h00000000} /* (25, 25, 11) {real, imag} */,
  {32'hbf4d8fbd, 32'h00000000} /* (25, 25, 10) {real, imag} */,
  {32'hbfa4350f, 32'h00000000} /* (25, 25, 9) {real, imag} */,
  {32'hbfa30b85, 32'h00000000} /* (25, 25, 8) {real, imag} */,
  {32'hbf312a0d, 32'h00000000} /* (25, 25, 7) {real, imag} */,
  {32'hbefdee24, 32'h00000000} /* (25, 25, 6) {real, imag} */,
  {32'hbeb4cb0f, 32'h00000000} /* (25, 25, 5) {real, imag} */,
  {32'hbee08ba6, 32'h00000000} /* (25, 25, 4) {real, imag} */,
  {32'hbf06232b, 32'h00000000} /* (25, 25, 3) {real, imag} */,
  {32'hbebc6724, 32'h00000000} /* (25, 25, 2) {real, imag} */,
  {32'hbf228593, 32'h00000000} /* (25, 25, 1) {real, imag} */,
  {32'hbf24c368, 32'h00000000} /* (25, 25, 0) {real, imag} */,
  {32'hbeedc929, 32'h00000000} /* (25, 24, 31) {real, imag} */,
  {32'hbf457e88, 32'h00000000} /* (25, 24, 30) {real, imag} */,
  {32'hbf3072e3, 32'h00000000} /* (25, 24, 29) {real, imag} */,
  {32'hbf0d5288, 32'h00000000} /* (25, 24, 28) {real, imag} */,
  {32'hbec34ed3, 32'h00000000} /* (25, 24, 27) {real, imag} */,
  {32'hbf1ec434, 32'h00000000} /* (25, 24, 26) {real, imag} */,
  {32'hbf9189b3, 32'h00000000} /* (25, 24, 25) {real, imag} */,
  {32'hbf3b7fc0, 32'h00000000} /* (25, 24, 24) {real, imag} */,
  {32'hbf3de346, 32'h00000000} /* (25, 24, 23) {real, imag} */,
  {32'hbf5cbd97, 32'h00000000} /* (25, 24, 22) {real, imag} */,
  {32'hbdd7096c, 32'h00000000} /* (25, 24, 21) {real, imag} */,
  {32'h3f571774, 32'h00000000} /* (25, 24, 20) {real, imag} */,
  {32'h3f0cc551, 32'h00000000} /* (25, 24, 19) {real, imag} */,
  {32'h3f1855e1, 32'h00000000} /* (25, 24, 18) {real, imag} */,
  {32'h3e7e6afb, 32'h00000000} /* (25, 24, 17) {real, imag} */,
  {32'h3e592e04, 32'h00000000} /* (25, 24, 16) {real, imag} */,
  {32'h3f3fe766, 32'h00000000} /* (25, 24, 15) {real, imag} */,
  {32'h3fa63c44, 32'h00000000} /* (25, 24, 14) {real, imag} */,
  {32'h3f638c25, 32'h00000000} /* (25, 24, 13) {real, imag} */,
  {32'h3e417464, 32'h00000000} /* (25, 24, 12) {real, imag} */,
  {32'hbe7e9bd5, 32'h00000000} /* (25, 24, 11) {real, imag} */,
  {32'hbf697652, 32'h00000000} /* (25, 24, 10) {real, imag} */,
  {32'hbf907754, 32'h00000000} /* (25, 24, 9) {real, imag} */,
  {32'hbf4d73f9, 32'h00000000} /* (25, 24, 8) {real, imag} */,
  {32'hbeebd61f, 32'h00000000} /* (25, 24, 7) {real, imag} */,
  {32'hbf17e92b, 32'h00000000} /* (25, 24, 6) {real, imag} */,
  {32'hbefcb78e, 32'h00000000} /* (25, 24, 5) {real, imag} */,
  {32'hbf348a6f, 32'h00000000} /* (25, 24, 4) {real, imag} */,
  {32'hbf5070c7, 32'h00000000} /* (25, 24, 3) {real, imag} */,
  {32'hbf2ea801, 32'h00000000} /* (25, 24, 2) {real, imag} */,
  {32'hbf882549, 32'h00000000} /* (25, 24, 1) {real, imag} */,
  {32'hbf37d392, 32'h00000000} /* (25, 24, 0) {real, imag} */,
  {32'hbe91ba9b, 32'h00000000} /* (25, 23, 31) {real, imag} */,
  {32'hbefca8cb, 32'h00000000} /* (25, 23, 30) {real, imag} */,
  {32'hbf90cdd7, 32'h00000000} /* (25, 23, 29) {real, imag} */,
  {32'hbf82015b, 32'h00000000} /* (25, 23, 28) {real, imag} */,
  {32'hbf3857ac, 32'h00000000} /* (25, 23, 27) {real, imag} */,
  {32'hbf7a01b1, 32'h00000000} /* (25, 23, 26) {real, imag} */,
  {32'hbfabb94d, 32'h00000000} /* (25, 23, 25) {real, imag} */,
  {32'hbf3f26cd, 32'h00000000} /* (25, 23, 24) {real, imag} */,
  {32'hbf98833b, 32'h00000000} /* (25, 23, 23) {real, imag} */,
  {32'hbfac845f, 32'h00000000} /* (25, 23, 22) {real, imag} */,
  {32'hbd60c11b, 32'h00000000} /* (25, 23, 21) {real, imag} */,
  {32'h3f7db543, 32'h00000000} /* (25, 23, 20) {real, imag} */,
  {32'h3f2a79f2, 32'h00000000} /* (25, 23, 19) {real, imag} */,
  {32'h3f356cfd, 32'h00000000} /* (25, 23, 18) {real, imag} */,
  {32'h3f556ae1, 32'h00000000} /* (25, 23, 17) {real, imag} */,
  {32'h3f118bf7, 32'h00000000} /* (25, 23, 16) {real, imag} */,
  {32'h3fb52958, 32'h00000000} /* (25, 23, 15) {real, imag} */,
  {32'h3faa437a, 32'h00000000} /* (25, 23, 14) {real, imag} */,
  {32'h3f059f7a, 32'h00000000} /* (25, 23, 13) {real, imag} */,
  {32'h3e7d49ac, 32'h00000000} /* (25, 23, 12) {real, imag} */,
  {32'h3d8cfd7a, 32'h00000000} /* (25, 23, 11) {real, imag} */,
  {32'hbf216fd1, 32'h00000000} /* (25, 23, 10) {real, imag} */,
  {32'hbf510372, 32'h00000000} /* (25, 23, 9) {real, imag} */,
  {32'hbeca7c82, 32'h00000000} /* (25, 23, 8) {real, imag} */,
  {32'hbecdc591, 32'h00000000} /* (25, 23, 7) {real, imag} */,
  {32'hbf8aafc8, 32'h00000000} /* (25, 23, 6) {real, imag} */,
  {32'hbfc203a6, 32'h00000000} /* (25, 23, 5) {real, imag} */,
  {32'hbf8e2986, 32'h00000000} /* (25, 23, 4) {real, imag} */,
  {32'hbf128d9b, 32'h00000000} /* (25, 23, 3) {real, imag} */,
  {32'hbf410e40, 32'h00000000} /* (25, 23, 2) {real, imag} */,
  {32'hbfaba5db, 32'h00000000} /* (25, 23, 1) {real, imag} */,
  {32'hbf5848ec, 32'h00000000} /* (25, 23, 0) {real, imag} */,
  {32'hbf505d55, 32'h00000000} /* (25, 22, 31) {real, imag} */,
  {32'hbf6d2233, 32'h00000000} /* (25, 22, 30) {real, imag} */,
  {32'hbf839511, 32'h00000000} /* (25, 22, 29) {real, imag} */,
  {32'hbf8adc2d, 32'h00000000} /* (25, 22, 28) {real, imag} */,
  {32'hbf5ad867, 32'h00000000} /* (25, 22, 27) {real, imag} */,
  {32'hbf56bc19, 32'h00000000} /* (25, 22, 26) {real, imag} */,
  {32'hbf3b37a6, 32'h00000000} /* (25, 22, 25) {real, imag} */,
  {32'hbf67248e, 32'h00000000} /* (25, 22, 24) {real, imag} */,
  {32'hbf7f862d, 32'h00000000} /* (25, 22, 23) {real, imag} */,
  {32'hbf5a0e13, 32'h00000000} /* (25, 22, 22) {real, imag} */,
  {32'hbdb29405, 32'h00000000} /* (25, 22, 21) {real, imag} */,
  {32'h3f2ffb62, 32'h00000000} /* (25, 22, 20) {real, imag} */,
  {32'h3f60a2a7, 32'h00000000} /* (25, 22, 19) {real, imag} */,
  {32'h3fab978f, 32'h00000000} /* (25, 22, 18) {real, imag} */,
  {32'h3f76e3a9, 32'h00000000} /* (25, 22, 17) {real, imag} */,
  {32'h3f245479, 32'h00000000} /* (25, 22, 16) {real, imag} */,
  {32'h3f809571, 32'h00000000} /* (25, 22, 15) {real, imag} */,
  {32'h3f72ff6f, 32'h00000000} /* (25, 22, 14) {real, imag} */,
  {32'h3f9e5144, 32'h00000000} /* (25, 22, 13) {real, imag} */,
  {32'h3f9430d8, 32'h00000000} /* (25, 22, 12) {real, imag} */,
  {32'h3f43a2ff, 32'h00000000} /* (25, 22, 11) {real, imag} */,
  {32'hbeb08618, 32'h00000000} /* (25, 22, 10) {real, imag} */,
  {32'hbf992636, 32'h00000000} /* (25, 22, 9) {real, imag} */,
  {32'hbf67ea46, 32'h00000000} /* (25, 22, 8) {real, imag} */,
  {32'hbf8e9249, 32'h00000000} /* (25, 22, 7) {real, imag} */,
  {32'hbf88795c, 32'h00000000} /* (25, 22, 6) {real, imag} */,
  {32'hbfbf130e, 32'h00000000} /* (25, 22, 5) {real, imag} */,
  {32'hbf71f68a, 32'h00000000} /* (25, 22, 4) {real, imag} */,
  {32'hbf4f4f9e, 32'h00000000} /* (25, 22, 3) {real, imag} */,
  {32'hbf126588, 32'h00000000} /* (25, 22, 2) {real, imag} */,
  {32'hbf09f976, 32'h00000000} /* (25, 22, 1) {real, imag} */,
  {32'hbf107d9c, 32'h00000000} /* (25, 22, 0) {real, imag} */,
  {32'hbf290d16, 32'h00000000} /* (25, 21, 31) {real, imag} */,
  {32'hbf5ac481, 32'h00000000} /* (25, 21, 30) {real, imag} */,
  {32'hbeda1133, 32'h00000000} /* (25, 21, 29) {real, imag} */,
  {32'hbece513d, 32'h00000000} /* (25, 21, 28) {real, imag} */,
  {32'hbf3a3dc9, 32'h00000000} /* (25, 21, 27) {real, imag} */,
  {32'hbf0812c1, 32'h00000000} /* (25, 21, 26) {real, imag} */,
  {32'hbf0aa3a7, 32'h00000000} /* (25, 21, 25) {real, imag} */,
  {32'hbeee5bc4, 32'h00000000} /* (25, 21, 24) {real, imag} */,
  {32'hbea4f092, 32'h00000000} /* (25, 21, 23) {real, imag} */,
  {32'h3e651010, 32'h00000000} /* (25, 21, 22) {real, imag} */,
  {32'h3ec361e0, 32'h00000000} /* (25, 21, 21) {real, imag} */,
  {32'h3e759115, 32'h00000000} /* (25, 21, 20) {real, imag} */,
  {32'h3c8ee564, 32'h00000000} /* (25, 21, 19) {real, imag} */,
  {32'h3ef0ab88, 32'h00000000} /* (25, 21, 18) {real, imag} */,
  {32'h3f30d8ec, 32'h00000000} /* (25, 21, 17) {real, imag} */,
  {32'h3eae532d, 32'h00000000} /* (25, 21, 16) {real, imag} */,
  {32'h3e8b9732, 32'h00000000} /* (25, 21, 15) {real, imag} */,
  {32'h3f170b8b, 32'h00000000} /* (25, 21, 14) {real, imag} */,
  {32'h3f78b955, 32'h00000000} /* (25, 21, 13) {real, imag} */,
  {32'h3f8e1c1a, 32'h00000000} /* (25, 21, 12) {real, imag} */,
  {32'h3e91434a, 32'h00000000} /* (25, 21, 11) {real, imag} */,
  {32'hbf3e0a82, 32'h00000000} /* (25, 21, 10) {real, imag} */,
  {32'hbfebad34, 32'h00000000} /* (25, 21, 9) {real, imag} */,
  {32'hbfa40282, 32'h00000000} /* (25, 21, 8) {real, imag} */,
  {32'hbf706e4c, 32'h00000000} /* (25, 21, 7) {real, imag} */,
  {32'h3db064d5, 32'h00000000} /* (25, 21, 6) {real, imag} */,
  {32'hbe834744, 32'h00000000} /* (25, 21, 5) {real, imag} */,
  {32'hbe3b07b9, 32'h00000000} /* (25, 21, 4) {real, imag} */,
  {32'hbe6318ee, 32'h00000000} /* (25, 21, 3) {real, imag} */,
  {32'h3df3eb5c, 32'h00000000} /* (25, 21, 2) {real, imag} */,
  {32'h3cc31992, 32'h00000000} /* (25, 21, 1) {real, imag} */,
  {32'h3dc04e3f, 32'h00000000} /* (25, 21, 0) {real, imag} */,
  {32'h3e84e228, 32'h00000000} /* (25, 20, 31) {real, imag} */,
  {32'h3e580be1, 32'h00000000} /* (25, 20, 30) {real, imag} */,
  {32'h3f30ec6c, 32'h00000000} /* (25, 20, 29) {real, imag} */,
  {32'h3f50bd86, 32'h00000000} /* (25, 20, 28) {real, imag} */,
  {32'h3f4ec636, 32'h00000000} /* (25, 20, 27) {real, imag} */,
  {32'h3f255e68, 32'h00000000} /* (25, 20, 26) {real, imag} */,
  {32'h3ddc3e59, 32'h00000000} /* (25, 20, 25) {real, imag} */,
  {32'h3ec2b7cd, 32'h00000000} /* (25, 20, 24) {real, imag} */,
  {32'h3fa38b0f, 32'h00000000} /* (25, 20, 23) {real, imag} */,
  {32'h3fb6b772, 32'h00000000} /* (25, 20, 22) {real, imag} */,
  {32'h3f7feef3, 32'h00000000} /* (25, 20, 21) {real, imag} */,
  {32'hbe23484a, 32'h00000000} /* (25, 20, 20) {real, imag} */,
  {32'hbf21a53d, 32'h00000000} /* (25, 20, 19) {real, imag} */,
  {32'hbedb9359, 32'h00000000} /* (25, 20, 18) {real, imag} */,
  {32'hbe96a221, 32'h00000000} /* (25, 20, 17) {real, imag} */,
  {32'hbf16684f, 32'h00000000} /* (25, 20, 16) {real, imag} */,
  {32'hbf7fdeb1, 32'h00000000} /* (25, 20, 15) {real, imag} */,
  {32'hbf28c127, 32'h00000000} /* (25, 20, 14) {real, imag} */,
  {32'hbe67dc6e, 32'h00000000} /* (25, 20, 13) {real, imag} */,
  {32'hbe260eae, 32'h00000000} /* (25, 20, 12) {real, imag} */,
  {32'hbf1cb590, 32'h00000000} /* (25, 20, 11) {real, imag} */,
  {32'hbe91c269, 32'h00000000} /* (25, 20, 10) {real, imag} */,
  {32'hbe800d0e, 32'h00000000} /* (25, 20, 9) {real, imag} */,
  {32'h3e5a5f34, 32'h00000000} /* (25, 20, 8) {real, imag} */,
  {32'h3eff0606, 32'h00000000} /* (25, 20, 7) {real, imag} */,
  {32'h3f8a82ba, 32'h00000000} /* (25, 20, 6) {real, imag} */,
  {32'h3ec0d5e8, 32'h00000000} /* (25, 20, 5) {real, imag} */,
  {32'h3f10a529, 32'h00000000} /* (25, 20, 4) {real, imag} */,
  {32'h3ed34e25, 32'h00000000} /* (25, 20, 3) {real, imag} */,
  {32'h3ec980e4, 32'h00000000} /* (25, 20, 2) {real, imag} */,
  {32'h3f536084, 32'h00000000} /* (25, 20, 1) {real, imag} */,
  {32'h3f401e3b, 32'h00000000} /* (25, 20, 0) {real, imag} */,
  {32'h3f1d13e0, 32'h00000000} /* (25, 19, 31) {real, imag} */,
  {32'h3f37ba16, 32'h00000000} /* (25, 19, 30) {real, imag} */,
  {32'h3f2a10cf, 32'h00000000} /* (25, 19, 29) {real, imag} */,
  {32'h3f51c9e3, 32'h00000000} /* (25, 19, 28) {real, imag} */,
  {32'h3fa57785, 32'h00000000} /* (25, 19, 27) {real, imag} */,
  {32'h3f923b3f, 32'h00000000} /* (25, 19, 26) {real, imag} */,
  {32'h3f113e5c, 32'h00000000} /* (25, 19, 25) {real, imag} */,
  {32'h3f04f7ab, 32'h00000000} /* (25, 19, 24) {real, imag} */,
  {32'h3f8be81e, 32'h00000000} /* (25, 19, 23) {real, imag} */,
  {32'h3f9e180d, 32'h00000000} /* (25, 19, 22) {real, imag} */,
  {32'h3f287078, 32'h00000000} /* (25, 19, 21) {real, imag} */,
  {32'hbedc9ee7, 32'h00000000} /* (25, 19, 20) {real, imag} */,
  {32'hbeb89b74, 32'h00000000} /* (25, 19, 19) {real, imag} */,
  {32'hbf1d3de5, 32'h00000000} /* (25, 19, 18) {real, imag} */,
  {32'hbf30aca0, 32'h00000000} /* (25, 19, 17) {real, imag} */,
  {32'hbec1764c, 32'h00000000} /* (25, 19, 16) {real, imag} */,
  {32'hbebd6876, 32'h00000000} /* (25, 19, 15) {real, imag} */,
  {32'hbec97e2b, 32'h00000000} /* (25, 19, 14) {real, imag} */,
  {32'hbed65a99, 32'h00000000} /* (25, 19, 13) {real, imag} */,
  {32'hbf571d10, 32'h00000000} /* (25, 19, 12) {real, imag} */,
  {32'hbeec02ac, 32'h00000000} /* (25, 19, 11) {real, imag} */,
  {32'h3f2de2f3, 32'h00000000} /* (25, 19, 10) {real, imag} */,
  {32'h3f5cc9cb, 32'h00000000} /* (25, 19, 9) {real, imag} */,
  {32'h3f39de69, 32'h00000000} /* (25, 19, 8) {real, imag} */,
  {32'h3f7250da, 32'h00000000} /* (25, 19, 7) {real, imag} */,
  {32'h3f4b8428, 32'h00000000} /* (25, 19, 6) {real, imag} */,
  {32'h3ea70ec1, 32'h00000000} /* (25, 19, 5) {real, imag} */,
  {32'h3eb6d601, 32'h00000000} /* (25, 19, 4) {real, imag} */,
  {32'h3e454663, 32'h00000000} /* (25, 19, 3) {real, imag} */,
  {32'h3ea6a140, 32'h00000000} /* (25, 19, 2) {real, imag} */,
  {32'h3f071d10, 32'h00000000} /* (25, 19, 1) {real, imag} */,
  {32'h3ec73fae, 32'h00000000} /* (25, 19, 0) {real, imag} */,
  {32'h3f52b558, 32'h00000000} /* (25, 18, 31) {real, imag} */,
  {32'h3f41ea60, 32'h00000000} /* (25, 18, 30) {real, imag} */,
  {32'h3ea192e0, 32'h00000000} /* (25, 18, 29) {real, imag} */,
  {32'h3edc9775, 32'h00000000} /* (25, 18, 28) {real, imag} */,
  {32'h3f87c883, 32'h00000000} /* (25, 18, 27) {real, imag} */,
  {32'h3f7a3df4, 32'h00000000} /* (25, 18, 26) {real, imag} */,
  {32'h3f59c868, 32'h00000000} /* (25, 18, 25) {real, imag} */,
  {32'h3f6d6d11, 32'h00000000} /* (25, 18, 24) {real, imag} */,
  {32'h3f1e381a, 32'h00000000} /* (25, 18, 23) {real, imag} */,
  {32'h3f1efcdf, 32'h00000000} /* (25, 18, 22) {real, imag} */,
  {32'h3e98b1e7, 32'h00000000} /* (25, 18, 21) {real, imag} */,
  {32'hbece15f8, 32'h00000000} /* (25, 18, 20) {real, imag} */,
  {32'hbeacc694, 32'h00000000} /* (25, 18, 19) {real, imag} */,
  {32'hbf3289c8, 32'h00000000} /* (25, 18, 18) {real, imag} */,
  {32'hbf5c3e72, 32'h00000000} /* (25, 18, 17) {real, imag} */,
  {32'hbe97f2ad, 32'h00000000} /* (25, 18, 16) {real, imag} */,
  {32'hbeb8e2d4, 32'h00000000} /* (25, 18, 15) {real, imag} */,
  {32'hbeedecb1, 32'h00000000} /* (25, 18, 14) {real, imag} */,
  {32'hbf1dbcb9, 32'h00000000} /* (25, 18, 13) {real, imag} */,
  {32'hbf0c5774, 32'h00000000} /* (25, 18, 12) {real, imag} */,
  {32'hbe1d31b8, 32'h00000000} /* (25, 18, 11) {real, imag} */,
  {32'h3eb0813f, 32'h00000000} /* (25, 18, 10) {real, imag} */,
  {32'h3f4c5ea1, 32'h00000000} /* (25, 18, 9) {real, imag} */,
  {32'h3f45ceb6, 32'h00000000} /* (25, 18, 8) {real, imag} */,
  {32'h3f800231, 32'h00000000} /* (25, 18, 7) {real, imag} */,
  {32'h3f65feba, 32'h00000000} /* (25, 18, 6) {real, imag} */,
  {32'h3f00c2a2, 32'h00000000} /* (25, 18, 5) {real, imag} */,
  {32'h3e20a77d, 32'h00000000} /* (25, 18, 4) {real, imag} */,
  {32'h3e2a8736, 32'h00000000} /* (25, 18, 3) {real, imag} */,
  {32'h3f6cb1a6, 32'h00000000} /* (25, 18, 2) {real, imag} */,
  {32'h3f0e8874, 32'h00000000} /* (25, 18, 1) {real, imag} */,
  {32'h3e6b83f2, 32'h00000000} /* (25, 18, 0) {real, imag} */,
  {32'h3ea8387b, 32'h00000000} /* (25, 17, 31) {real, imag} */,
  {32'h3eddbde3, 32'h00000000} /* (25, 17, 30) {real, imag} */,
  {32'h3f2a0876, 32'h00000000} /* (25, 17, 29) {real, imag} */,
  {32'h3f6bb327, 32'h00000000} /* (25, 17, 28) {real, imag} */,
  {32'h3fa23ebe, 32'h00000000} /* (25, 17, 27) {real, imag} */,
  {32'h3f93a346, 32'h00000000} /* (25, 17, 26) {real, imag} */,
  {32'h3f999d02, 32'h00000000} /* (25, 17, 25) {real, imag} */,
  {32'h3fb9ad0a, 32'h00000000} /* (25, 17, 24) {real, imag} */,
  {32'h3f9a5a1b, 32'h00000000} /* (25, 17, 23) {real, imag} */,
  {32'h3f526af0, 32'h00000000} /* (25, 17, 22) {real, imag} */,
  {32'h3ec40044, 32'h00000000} /* (25, 17, 21) {real, imag} */,
  {32'hbe9bcb38, 32'h00000000} /* (25, 17, 20) {real, imag} */,
  {32'hbea7f924, 32'h00000000} /* (25, 17, 19) {real, imag} */,
  {32'hbebeb911, 32'h00000000} /* (25, 17, 18) {real, imag} */,
  {32'hbf23f4da, 32'h00000000} /* (25, 17, 17) {real, imag} */,
  {32'hbf07a826, 32'h00000000} /* (25, 17, 16) {real, imag} */,
  {32'hbef4a616, 32'h00000000} /* (25, 17, 15) {real, imag} */,
  {32'hbf406b03, 32'h00000000} /* (25, 17, 14) {real, imag} */,
  {32'hbf62dedd, 32'h00000000} /* (25, 17, 13) {real, imag} */,
  {32'hbf172e90, 32'h00000000} /* (25, 17, 12) {real, imag} */,
  {32'hbed7da54, 32'h00000000} /* (25, 17, 11) {real, imag} */,
  {32'h3e6fc891, 32'h00000000} /* (25, 17, 10) {real, imag} */,
  {32'h3f24d174, 32'h00000000} /* (25, 17, 9) {real, imag} */,
  {32'h3f71cd5d, 32'h00000000} /* (25, 17, 8) {real, imag} */,
  {32'h3fcdcfa3, 32'h00000000} /* (25, 17, 7) {real, imag} */,
  {32'h3fa8e6a3, 32'h00000000} /* (25, 17, 6) {real, imag} */,
  {32'h3ef6ecef, 32'h00000000} /* (25, 17, 5) {real, imag} */,
  {32'h3ea1feeb, 32'h00000000} /* (25, 17, 4) {real, imag} */,
  {32'h3f088012, 32'h00000000} /* (25, 17, 3) {real, imag} */,
  {32'h3f1506d8, 32'h00000000} /* (25, 17, 2) {real, imag} */,
  {32'h3e7dd377, 32'h00000000} /* (25, 17, 1) {real, imag} */,
  {32'h3e9abf0a, 32'h00000000} /* (25, 17, 0) {real, imag} */,
  {32'h3f00796e, 32'h00000000} /* (25, 16, 31) {real, imag} */,
  {32'h3f54fa67, 32'h00000000} /* (25, 16, 30) {real, imag} */,
  {32'h3f6e6b78, 32'h00000000} /* (25, 16, 29) {real, imag} */,
  {32'h3fa04518, 32'h00000000} /* (25, 16, 28) {real, imag} */,
  {32'h3f02e431, 32'h00000000} /* (25, 16, 27) {real, imag} */,
  {32'h3f102870, 32'h00000000} /* (25, 16, 26) {real, imag} */,
  {32'h3f702972, 32'h00000000} /* (25, 16, 25) {real, imag} */,
  {32'h3f68069e, 32'h00000000} /* (25, 16, 24) {real, imag} */,
  {32'h3f8df369, 32'h00000000} /* (25, 16, 23) {real, imag} */,
  {32'h3f3e8bc6, 32'h00000000} /* (25, 16, 22) {real, imag} */,
  {32'h3e9a1fdc, 32'h00000000} /* (25, 16, 21) {real, imag} */,
  {32'hbe90e090, 32'h00000000} /* (25, 16, 20) {real, imag} */,
  {32'hbeefb9c2, 32'h00000000} /* (25, 16, 19) {real, imag} */,
  {32'hbe3bef15, 32'h00000000} /* (25, 16, 18) {real, imag} */,
  {32'hbef68ce1, 32'h00000000} /* (25, 16, 17) {real, imag} */,
  {32'hbf38353f, 32'h00000000} /* (25, 16, 16) {real, imag} */,
  {32'hbedfef46, 32'h00000000} /* (25, 16, 15) {real, imag} */,
  {32'hbf4b24d2, 32'h00000000} /* (25, 16, 14) {real, imag} */,
  {32'hbf6d1d4f, 32'h00000000} /* (25, 16, 13) {real, imag} */,
  {32'hbf813606, 32'h00000000} /* (25, 16, 12) {real, imag} */,
  {32'hbf5cf348, 32'h00000000} /* (25, 16, 11) {real, imag} */,
  {32'h3e5c4e5f, 32'h00000000} /* (25, 16, 10) {real, imag} */,
  {32'h3edc9ba9, 32'h00000000} /* (25, 16, 9) {real, imag} */,
  {32'h3f328075, 32'h00000000} /* (25, 16, 8) {real, imag} */,
  {32'h3fde4553, 32'h00000000} /* (25, 16, 7) {real, imag} */,
  {32'h4017c84b, 32'h00000000} /* (25, 16, 6) {real, imag} */,
  {32'h3f8cf6c3, 32'h00000000} /* (25, 16, 5) {real, imag} */,
  {32'h3f8b5f00, 32'h00000000} /* (25, 16, 4) {real, imag} */,
  {32'h3f9323f0, 32'h00000000} /* (25, 16, 3) {real, imag} */,
  {32'h3f5586ba, 32'h00000000} /* (25, 16, 2) {real, imag} */,
  {32'h3f1bb842, 32'h00000000} /* (25, 16, 1) {real, imag} */,
  {32'h3f417810, 32'h00000000} /* (25, 16, 0) {real, imag} */,
  {32'h3f0a9720, 32'h00000000} /* (25, 15, 31) {real, imag} */,
  {32'h3f453dfa, 32'h00000000} /* (25, 15, 30) {real, imag} */,
  {32'h3f3cc16f, 32'h00000000} /* (25, 15, 29) {real, imag} */,
  {32'h3f9713a9, 32'h00000000} /* (25, 15, 28) {real, imag} */,
  {32'h3f014dd0, 32'h00000000} /* (25, 15, 27) {real, imag} */,
  {32'h3e81ee36, 32'h00000000} /* (25, 15, 26) {real, imag} */,
  {32'h3db6bec0, 32'h00000000} /* (25, 15, 25) {real, imag} */,
  {32'h3efe9f5d, 32'h00000000} /* (25, 15, 24) {real, imag} */,
  {32'h3f897d54, 32'h00000000} /* (25, 15, 23) {real, imag} */,
  {32'h3f08e4d3, 32'h00000000} /* (25, 15, 22) {real, imag} */,
  {32'h3ea82f0a, 32'h00000000} /* (25, 15, 21) {real, imag} */,
  {32'hbe4fe518, 32'h00000000} /* (25, 15, 20) {real, imag} */,
  {32'hbf3fe815, 32'h00000000} /* (25, 15, 19) {real, imag} */,
  {32'hbf0814dc, 32'h00000000} /* (25, 15, 18) {real, imag} */,
  {32'hbf6f3426, 32'h00000000} /* (25, 15, 17) {real, imag} */,
  {32'hbf749551, 32'h00000000} /* (25, 15, 16) {real, imag} */,
  {32'hbf3ffce2, 32'h00000000} /* (25, 15, 15) {real, imag} */,
  {32'hbf6001ab, 32'h00000000} /* (25, 15, 14) {real, imag} */,
  {32'hbf110994, 32'h00000000} /* (25, 15, 13) {real, imag} */,
  {32'hbf0154ab, 32'h00000000} /* (25, 15, 12) {real, imag} */,
  {32'hbec9b1cd, 32'h00000000} /* (25, 15, 11) {real, imag} */,
  {32'h3e7707e4, 32'h00000000} /* (25, 15, 10) {real, imag} */,
  {32'h3ef993f9, 32'h00000000} /* (25, 15, 9) {real, imag} */,
  {32'h3ee491d2, 32'h00000000} /* (25, 15, 8) {real, imag} */,
  {32'h3f25a226, 32'h00000000} /* (25, 15, 7) {real, imag} */,
  {32'h3f5fccc5, 32'h00000000} /* (25, 15, 6) {real, imag} */,
  {32'h3f2e8936, 32'h00000000} /* (25, 15, 5) {real, imag} */,
  {32'h3f796855, 32'h00000000} /* (25, 15, 4) {real, imag} */,
  {32'h3f494b65, 32'h00000000} /* (25, 15, 3) {real, imag} */,
  {32'h3ef84cd6, 32'h00000000} /* (25, 15, 2) {real, imag} */,
  {32'h3edc6d2e, 32'h00000000} /* (25, 15, 1) {real, imag} */,
  {32'h3edc819f, 32'h00000000} /* (25, 15, 0) {real, imag} */,
  {32'h3edadfc6, 32'h00000000} /* (25, 14, 31) {real, imag} */,
  {32'h3f1659f8, 32'h00000000} /* (25, 14, 30) {real, imag} */,
  {32'h3f1a5cf0, 32'h00000000} /* (25, 14, 29) {real, imag} */,
  {32'h3f3d4cf5, 32'h00000000} /* (25, 14, 28) {real, imag} */,
  {32'h3f5a260b, 32'h00000000} /* (25, 14, 27) {real, imag} */,
  {32'h3f1a5c3c, 32'h00000000} /* (25, 14, 26) {real, imag} */,
  {32'h3e5375ec, 32'h00000000} /* (25, 14, 25) {real, imag} */,
  {32'h3ee7d50c, 32'h00000000} /* (25, 14, 24) {real, imag} */,
  {32'h3f5b3afa, 32'h00000000} /* (25, 14, 23) {real, imag} */,
  {32'h3ee41c05, 32'h00000000} /* (25, 14, 22) {real, imag} */,
  {32'h3e9815fc, 32'h00000000} /* (25, 14, 21) {real, imag} */,
  {32'hbdd9adf0, 32'h00000000} /* (25, 14, 20) {real, imag} */,
  {32'hbf263c38, 32'h00000000} /* (25, 14, 19) {real, imag} */,
  {32'hbf25723c, 32'h00000000} /* (25, 14, 18) {real, imag} */,
  {32'hbf705ec4, 32'h00000000} /* (25, 14, 17) {real, imag} */,
  {32'hbfa9932b, 32'h00000000} /* (25, 14, 16) {real, imag} */,
  {32'hbf5dd43a, 32'h00000000} /* (25, 14, 15) {real, imag} */,
  {32'hbf3d7e05, 32'h00000000} /* (25, 14, 14) {real, imag} */,
  {32'hbf68348e, 32'h00000000} /* (25, 14, 13) {real, imag} */,
  {32'hbf22f19f, 32'h00000000} /* (25, 14, 12) {real, imag} */,
  {32'hbefc4367, 32'h00000000} /* (25, 14, 11) {real, imag} */,
  {32'h3dee3eab, 32'h00000000} /* (25, 14, 10) {real, imag} */,
  {32'h3ef18ff5, 32'h00000000} /* (25, 14, 9) {real, imag} */,
  {32'h3f28dd1f, 32'h00000000} /* (25, 14, 8) {real, imag} */,
  {32'h3f363af1, 32'h00000000} /* (25, 14, 7) {real, imag} */,
  {32'h3f048dd7, 32'h00000000} /* (25, 14, 6) {real, imag} */,
  {32'h3f402a7a, 32'h00000000} /* (25, 14, 5) {real, imag} */,
  {32'h3f78baf3, 32'h00000000} /* (25, 14, 4) {real, imag} */,
  {32'h3f25185b, 32'h00000000} /* (25, 14, 3) {real, imag} */,
  {32'h3e9f07a2, 32'h00000000} /* (25, 14, 2) {real, imag} */,
  {32'h3f05cd1e, 32'h00000000} /* (25, 14, 1) {real, imag} */,
  {32'h3e813234, 32'h00000000} /* (25, 14, 0) {real, imag} */,
  {32'h3f00e13c, 32'h00000000} /* (25, 13, 31) {real, imag} */,
  {32'h3f70abfd, 32'h00000000} /* (25, 13, 30) {real, imag} */,
  {32'h3f3f839e, 32'h00000000} /* (25, 13, 29) {real, imag} */,
  {32'h3f9d88b6, 32'h00000000} /* (25, 13, 28) {real, imag} */,
  {32'h3fa6a7a7, 32'h00000000} /* (25, 13, 27) {real, imag} */,
  {32'h3f23876a, 32'h00000000} /* (25, 13, 26) {real, imag} */,
  {32'h3f36e7d7, 32'h00000000} /* (25, 13, 25) {real, imag} */,
  {32'h3f6b494f, 32'h00000000} /* (25, 13, 24) {real, imag} */,
  {32'h3f946d3c, 32'h00000000} /* (25, 13, 23) {real, imag} */,
  {32'h3f469b27, 32'h00000000} /* (25, 13, 22) {real, imag} */,
  {32'h3ea12dd4, 32'h00000000} /* (25, 13, 21) {real, imag} */,
  {32'hbe9adc5f, 32'h00000000} /* (25, 13, 20) {real, imag} */,
  {32'hbed7c3f7, 32'h00000000} /* (25, 13, 19) {real, imag} */,
  {32'hbea3815e, 32'h00000000} /* (25, 13, 18) {real, imag} */,
  {32'hbf525dcd, 32'h00000000} /* (25, 13, 17) {real, imag} */,
  {32'hbfbf3bef, 32'h00000000} /* (25, 13, 16) {real, imag} */,
  {32'hbf8c523b, 32'h00000000} /* (25, 13, 15) {real, imag} */,
  {32'hbf2f217e, 32'h00000000} /* (25, 13, 14) {real, imag} */,
  {32'hbf0b473b, 32'h00000000} /* (25, 13, 13) {real, imag} */,
  {32'hbf275722, 32'h00000000} /* (25, 13, 12) {real, imag} */,
  {32'hbf118701, 32'h00000000} /* (25, 13, 11) {real, imag} */,
  {32'h3f2e73b2, 32'h00000000} /* (25, 13, 10) {real, imag} */,
  {32'h3f34e2b8, 32'h00000000} /* (25, 13, 9) {real, imag} */,
  {32'h3f1cb3d1, 32'h00000000} /* (25, 13, 8) {real, imag} */,
  {32'h3f558719, 32'h00000000} /* (25, 13, 7) {real, imag} */,
  {32'h3f7c85a6, 32'h00000000} /* (25, 13, 6) {real, imag} */,
  {32'h3fad97dd, 32'h00000000} /* (25, 13, 5) {real, imag} */,
  {32'h3fbb96b6, 32'h00000000} /* (25, 13, 4) {real, imag} */,
  {32'h3f58f095, 32'h00000000} /* (25, 13, 3) {real, imag} */,
  {32'h3ef00984, 32'h00000000} /* (25, 13, 2) {real, imag} */,
  {32'h3ee77a14, 32'h00000000} /* (25, 13, 1) {real, imag} */,
  {32'h3eaec47b, 32'h00000000} /* (25, 13, 0) {real, imag} */,
  {32'h3f3b9676, 32'h00000000} /* (25, 12, 31) {real, imag} */,
  {32'h3fa8bb05, 32'h00000000} /* (25, 12, 30) {real, imag} */,
  {32'h3f390c23, 32'h00000000} /* (25, 12, 29) {real, imag} */,
  {32'h3f8d4c2d, 32'h00000000} /* (25, 12, 28) {real, imag} */,
  {32'h3f755e83, 32'h00000000} /* (25, 12, 27) {real, imag} */,
  {32'h3f1387af, 32'h00000000} /* (25, 12, 26) {real, imag} */,
  {32'h3f78e65c, 32'h00000000} /* (25, 12, 25) {real, imag} */,
  {32'h3f94c12e, 32'h00000000} /* (25, 12, 24) {real, imag} */,
  {32'h3f69b583, 32'h00000000} /* (25, 12, 23) {real, imag} */,
  {32'h3f283a22, 32'h00000000} /* (25, 12, 22) {real, imag} */,
  {32'h3ea6f820, 32'h00000000} /* (25, 12, 21) {real, imag} */,
  {32'hbf37dee7, 32'h00000000} /* (25, 12, 20) {real, imag} */,
  {32'hbf923551, 32'h00000000} /* (25, 12, 19) {real, imag} */,
  {32'hbfa0c8b2, 32'h00000000} /* (25, 12, 18) {real, imag} */,
  {32'hbf8aba3f, 32'h00000000} /* (25, 12, 17) {real, imag} */,
  {32'hbf86168f, 32'h00000000} /* (25, 12, 16) {real, imag} */,
  {32'hbf84c0fe, 32'h00000000} /* (25, 12, 15) {real, imag} */,
  {32'hbf1609ef, 32'h00000000} /* (25, 12, 14) {real, imag} */,
  {32'hbe83d424, 32'h00000000} /* (25, 12, 13) {real, imag} */,
  {32'hbf369fcd, 32'h00000000} /* (25, 12, 12) {real, imag} */,
  {32'hbf4c209d, 32'h00000000} /* (25, 12, 11) {real, imag} */,
  {32'h3f8fd847, 32'h00000000} /* (25, 12, 10) {real, imag} */,
  {32'h3f84e43e, 32'h00000000} /* (25, 12, 9) {real, imag} */,
  {32'h3f2c2d87, 32'h00000000} /* (25, 12, 8) {real, imag} */,
  {32'h3f6c7540, 32'h00000000} /* (25, 12, 7) {real, imag} */,
  {32'h3f93f5f6, 32'h00000000} /* (25, 12, 6) {real, imag} */,
  {32'h3f8084f6, 32'h00000000} /* (25, 12, 5) {real, imag} */,
  {32'h3f41b8b3, 32'h00000000} /* (25, 12, 4) {real, imag} */,
  {32'h3efdc5b8, 32'h00000000} /* (25, 12, 3) {real, imag} */,
  {32'h3f556471, 32'h00000000} /* (25, 12, 2) {real, imag} */,
  {32'h3f54f1aa, 32'h00000000} /* (25, 12, 1) {real, imag} */,
  {32'h3efc65cf, 32'h00000000} /* (25, 12, 0) {real, imag} */,
  {32'h3f1ec64e, 32'h00000000} /* (25, 11, 31) {real, imag} */,
  {32'h3f7ca2bb, 32'h00000000} /* (25, 11, 30) {real, imag} */,
  {32'h3eba7607, 32'h00000000} /* (25, 11, 29) {real, imag} */,
  {32'h3f0bad04, 32'h00000000} /* (25, 11, 28) {real, imag} */,
  {32'h3eefbcd3, 32'h00000000} /* (25, 11, 27) {real, imag} */,
  {32'h3ec50175, 32'h00000000} /* (25, 11, 26) {real, imag} */,
  {32'h3f30e21e, 32'h00000000} /* (25, 11, 25) {real, imag} */,
  {32'h3f95bc0e, 32'h00000000} /* (25, 11, 24) {real, imag} */,
  {32'h3f837228, 32'h00000000} /* (25, 11, 23) {real, imag} */,
  {32'h3f8cb912, 32'h00000000} /* (25, 11, 22) {real, imag} */,
  {32'h3eb7f671, 32'h00000000} /* (25, 11, 21) {real, imag} */,
  {32'hbeadb6a9, 32'h00000000} /* (25, 11, 20) {real, imag} */,
  {32'hbf276742, 32'h00000000} /* (25, 11, 19) {real, imag} */,
  {32'hbf9c352b, 32'h00000000} /* (25, 11, 18) {real, imag} */,
  {32'hbf76b08a, 32'h00000000} /* (25, 11, 17) {real, imag} */,
  {32'hbe4d6766, 32'h00000000} /* (25, 11, 16) {real, imag} */,
  {32'hbe604104, 32'h00000000} /* (25, 11, 15) {real, imag} */,
  {32'hbe87d1ff, 32'h00000000} /* (25, 11, 14) {real, imag} */,
  {32'hbeba234a, 32'h00000000} /* (25, 11, 13) {real, imag} */,
  {32'hbf0b0624, 32'h00000000} /* (25, 11, 12) {real, imag} */,
  {32'hbf1f59f4, 32'h00000000} /* (25, 11, 11) {real, imag} */,
  {32'h3e8c29bf, 32'h00000000} /* (25, 11, 10) {real, imag} */,
  {32'h3f538f04, 32'h00000000} /* (25, 11, 9) {real, imag} */,
  {32'h3f9b225e, 32'h00000000} /* (25, 11, 8) {real, imag} */,
  {32'h3fea5268, 32'h00000000} /* (25, 11, 7) {real, imag} */,
  {32'h3f919e6b, 32'h00000000} /* (25, 11, 6) {real, imag} */,
  {32'h3f17afdc, 32'h00000000} /* (25, 11, 5) {real, imag} */,
  {32'h3ecfaffc, 32'h00000000} /* (25, 11, 4) {real, imag} */,
  {32'h3e6db6cc, 32'h00000000} /* (25, 11, 3) {real, imag} */,
  {32'h3f2adf1d, 32'h00000000} /* (25, 11, 2) {real, imag} */,
  {32'h3f49acbf, 32'h00000000} /* (25, 11, 1) {real, imag} */,
  {32'h3f15a757, 32'h00000000} /* (25, 11, 0) {real, imag} */,
  {32'hbcda21bc, 32'h00000000} /* (25, 10, 31) {real, imag} */,
  {32'hbe31292c, 32'h00000000} /* (25, 10, 30) {real, imag} */,
  {32'hbf45421b, 32'h00000000} /* (25, 10, 29) {real, imag} */,
  {32'hbf0428d2, 32'h00000000} /* (25, 10, 28) {real, imag} */,
  {32'hbf1147c0, 32'h00000000} /* (25, 10, 27) {real, imag} */,
  {32'hbf399784, 32'h00000000} /* (25, 10, 26) {real, imag} */,
  {32'hbf32a9e9, 32'h00000000} /* (25, 10, 25) {real, imag} */,
  {32'hbd49366a, 32'h00000000} /* (25, 10, 24) {real, imag} */,
  {32'hbd5913f7, 32'h00000000} /* (25, 10, 23) {real, imag} */,
  {32'hbe1b9b4f, 32'h00000000} /* (25, 10, 22) {real, imag} */,
  {32'hbebaa2e7, 32'h00000000} /* (25, 10, 21) {real, imag} */,
  {32'h3ec14335, 32'h00000000} /* (25, 10, 20) {real, imag} */,
  {32'h3f281dc9, 32'h00000000} /* (25, 10, 19) {real, imag} */,
  {32'h3eb69c3b, 32'h00000000} /* (25, 10, 18) {real, imag} */,
  {32'h3f4f84af, 32'h00000000} /* (25, 10, 17) {real, imag} */,
  {32'h3f68d43e, 32'h00000000} /* (25, 10, 16) {real, imag} */,
  {32'h3f353ff2, 32'h00000000} /* (25, 10, 15) {real, imag} */,
  {32'h3ec21522, 32'h00000000} /* (25, 10, 14) {real, imag} */,
  {32'hbc1854d0, 32'h00000000} /* (25, 10, 13) {real, imag} */,
  {32'h3e23d423, 32'h00000000} /* (25, 10, 12) {real, imag} */,
  {32'h3f0e67b8, 32'h00000000} /* (25, 10, 11) {real, imag} */,
  {32'h3e6c1b30, 32'h00000000} /* (25, 10, 10) {real, imag} */,
  {32'hbe10feb4, 32'h00000000} /* (25, 10, 9) {real, imag} */,
  {32'hbe446dbb, 32'h00000000} /* (25, 10, 8) {real, imag} */,
  {32'h3f565ee7, 32'h00000000} /* (25, 10, 7) {real, imag} */,
  {32'h3d940a3f, 32'h00000000} /* (25, 10, 6) {real, imag} */,
  {32'hbe494fb6, 32'h00000000} /* (25, 10, 5) {real, imag} */,
  {32'hbeb50f82, 32'h00000000} /* (25, 10, 4) {real, imag} */,
  {32'hbf2faabc, 32'h00000000} /* (25, 10, 3) {real, imag} */,
  {32'hbe9665ba, 32'h00000000} /* (25, 10, 2) {real, imag} */,
  {32'hbf35fa31, 32'h00000000} /* (25, 10, 1) {real, imag} */,
  {32'hbee941fc, 32'h00000000} /* (25, 10, 0) {real, imag} */,
  {32'hbed62d06, 32'h00000000} /* (25, 9, 31) {real, imag} */,
  {32'hbf02ee54, 32'h00000000} /* (25, 9, 30) {real, imag} */,
  {32'hbf4a2ce1, 32'h00000000} /* (25, 9, 29) {real, imag} */,
  {32'hbf471576, 32'h00000000} /* (25, 9, 28) {real, imag} */,
  {32'hbf9d62e9, 32'h00000000} /* (25, 9, 27) {real, imag} */,
  {32'hbf951d0c, 32'h00000000} /* (25, 9, 26) {real, imag} */,
  {32'hbf60689e, 32'h00000000} /* (25, 9, 25) {real, imag} */,
  {32'hbf2a1709, 32'h00000000} /* (25, 9, 24) {real, imag} */,
  {32'hbeecf3d9, 32'h00000000} /* (25, 9, 23) {real, imag} */,
  {32'hbf10f023, 32'h00000000} /* (25, 9, 22) {real, imag} */,
  {32'hbee9684a, 32'h00000000} /* (25, 9, 21) {real, imag} */,
  {32'h3f1af58a, 32'h00000000} /* (25, 9, 20) {real, imag} */,
  {32'h3f672c18, 32'h00000000} /* (25, 9, 19) {real, imag} */,
  {32'h3f655ddb, 32'h00000000} /* (25, 9, 18) {real, imag} */,
  {32'h3f6a5694, 32'h00000000} /* (25, 9, 17) {real, imag} */,
  {32'h3f5202d6, 32'h00000000} /* (25, 9, 16) {real, imag} */,
  {32'h3f38aa6d, 32'h00000000} /* (25, 9, 15) {real, imag} */,
  {32'h3f8848e1, 32'h00000000} /* (25, 9, 14) {real, imag} */,
  {32'h3f1723f1, 32'h00000000} /* (25, 9, 13) {real, imag} */,
  {32'h3f248e9f, 32'h00000000} /* (25, 9, 12) {real, imag} */,
  {32'h3f43ad3a, 32'h00000000} /* (25, 9, 11) {real, imag} */,
  {32'h3d394f84, 32'h00000000} /* (25, 9, 10) {real, imag} */,
  {32'hbf000d92, 32'h00000000} /* (25, 9, 9) {real, imag} */,
  {32'hbf4ea5a4, 32'h00000000} /* (25, 9, 8) {real, imag} */,
  {32'hbec42ab1, 32'h00000000} /* (25, 9, 7) {real, imag} */,
  {32'hbf0f40e3, 32'h00000000} /* (25, 9, 6) {real, imag} */,
  {32'hbf629f1f, 32'h00000000} /* (25, 9, 5) {real, imag} */,
  {32'hbf38714d, 32'h00000000} /* (25, 9, 4) {real, imag} */,
  {32'hbf63374a, 32'h00000000} /* (25, 9, 3) {real, imag} */,
  {32'hbf4acb57, 32'h00000000} /* (25, 9, 2) {real, imag} */,
  {32'hbf967671, 32'h00000000} /* (25, 9, 1) {real, imag} */,
  {32'hbf59e0c1, 32'h00000000} /* (25, 9, 0) {real, imag} */,
  {32'hbe0587cc, 32'h00000000} /* (25, 8, 31) {real, imag} */,
  {32'hbe453565, 32'h00000000} /* (25, 8, 30) {real, imag} */,
  {32'hbf95beab, 32'h00000000} /* (25, 8, 29) {real, imag} */,
  {32'hbf815ad5, 32'h00000000} /* (25, 8, 28) {real, imag} */,
  {32'hbf154c36, 32'h00000000} /* (25, 8, 27) {real, imag} */,
  {32'hbf35bfa1, 32'h00000000} /* (25, 8, 26) {real, imag} */,
  {32'hbf859a5a, 32'h00000000} /* (25, 8, 25) {real, imag} */,
  {32'hbf525115, 32'h00000000} /* (25, 8, 24) {real, imag} */,
  {32'hbf0fa731, 32'h00000000} /* (25, 8, 23) {real, imag} */,
  {32'hbf417863, 32'h00000000} /* (25, 8, 22) {real, imag} */,
  {32'hbedfff5a, 32'h00000000} /* (25, 8, 21) {real, imag} */,
  {32'h3f237361, 32'h00000000} /* (25, 8, 20) {real, imag} */,
  {32'h3f57332d, 32'h00000000} /* (25, 8, 19) {real, imag} */,
  {32'h3f52d0ed, 32'h00000000} /* (25, 8, 18) {real, imag} */,
  {32'h3f450b35, 32'h00000000} /* (25, 8, 17) {real, imag} */,
  {32'h3f5c1674, 32'h00000000} /* (25, 8, 16) {real, imag} */,
  {32'h3f6606df, 32'h00000000} /* (25, 8, 15) {real, imag} */,
  {32'h3f616700, 32'h00000000} /* (25, 8, 14) {real, imag} */,
  {32'h3f5173b2, 32'h00000000} /* (25, 8, 13) {real, imag} */,
  {32'h3f2710c4, 32'h00000000} /* (25, 8, 12) {real, imag} */,
  {32'h3f150537, 32'h00000000} /* (25, 8, 11) {real, imag} */,
  {32'hbd4cbd44, 32'h00000000} /* (25, 8, 10) {real, imag} */,
  {32'hbe97f0da, 32'h00000000} /* (25, 8, 9) {real, imag} */,
  {32'hbf28c8b3, 32'h00000000} /* (25, 8, 8) {real, imag} */,
  {32'hbf67dc20, 32'h00000000} /* (25, 8, 7) {real, imag} */,
  {32'hbf7367da, 32'h00000000} /* (25, 8, 6) {real, imag} */,
  {32'hbf8613b1, 32'h00000000} /* (25, 8, 5) {real, imag} */,
  {32'hbede6b41, 32'h00000000} /* (25, 8, 4) {real, imag} */,
  {32'hbe8bd134, 32'h00000000} /* (25, 8, 3) {real, imag} */,
  {32'hbf46858e, 32'h00000000} /* (25, 8, 2) {real, imag} */,
  {32'hbfa57f74, 32'h00000000} /* (25, 8, 1) {real, imag} */,
  {32'hbf675c09, 32'h00000000} /* (25, 8, 0) {real, imag} */,
  {32'h39bba480, 32'h00000000} /* (25, 7, 31) {real, imag} */,
  {32'hbf119367, 32'h00000000} /* (25, 7, 30) {real, imag} */,
  {32'hbfc9843c, 32'h00000000} /* (25, 7, 29) {real, imag} */,
  {32'hbfd9bd42, 32'h00000000} /* (25, 7, 28) {real, imag} */,
  {32'hbf3726bc, 32'h00000000} /* (25, 7, 27) {real, imag} */,
  {32'hbe92094f, 32'h00000000} /* (25, 7, 26) {real, imag} */,
  {32'hbf5f7158, 32'h00000000} /* (25, 7, 25) {real, imag} */,
  {32'hbf5c8181, 32'h00000000} /* (25, 7, 24) {real, imag} */,
  {32'hbf56189d, 32'h00000000} /* (25, 7, 23) {real, imag} */,
  {32'hbf5bf632, 32'h00000000} /* (25, 7, 22) {real, imag} */,
  {32'hbeb0ec07, 32'h00000000} /* (25, 7, 21) {real, imag} */,
  {32'h3f7e6a73, 32'h00000000} /* (25, 7, 20) {real, imag} */,
  {32'h3f51d240, 32'h00000000} /* (25, 7, 19) {real, imag} */,
  {32'h3f148e7b, 32'h00000000} /* (25, 7, 18) {real, imag} */,
  {32'h3f1409c2, 32'h00000000} /* (25, 7, 17) {real, imag} */,
  {32'h3edb3dd7, 32'h00000000} /* (25, 7, 16) {real, imag} */,
  {32'h3f126a70, 32'h00000000} /* (25, 7, 15) {real, imag} */,
  {32'h3f249106, 32'h00000000} /* (25, 7, 14) {real, imag} */,
  {32'h3f25684b, 32'h00000000} /* (25, 7, 13) {real, imag} */,
  {32'h3f0374a0, 32'h00000000} /* (25, 7, 12) {real, imag} */,
  {32'h3e6b2a8b, 32'h00000000} /* (25, 7, 11) {real, imag} */,
  {32'hbe753763, 32'h00000000} /* (25, 7, 10) {real, imag} */,
  {32'hbf2bd394, 32'h00000000} /* (25, 7, 9) {real, imag} */,
  {32'hbf7a4560, 32'h00000000} /* (25, 7, 8) {real, imag} */,
  {32'hbf3a6801, 32'h00000000} /* (25, 7, 7) {real, imag} */,
  {32'hbf16fcf0, 32'h00000000} /* (25, 7, 6) {real, imag} */,
  {32'hbf919d6d, 32'h00000000} /* (25, 7, 5) {real, imag} */,
  {32'hbf6a8a0b, 32'h00000000} /* (25, 7, 4) {real, imag} */,
  {32'hbeafd26d, 32'h00000000} /* (25, 7, 3) {real, imag} */,
  {32'hbf8930f8, 32'h00000000} /* (25, 7, 2) {real, imag} */,
  {32'hbfb52e90, 32'h00000000} /* (25, 7, 1) {real, imag} */,
  {32'hbedae288, 32'h00000000} /* (25, 7, 0) {real, imag} */,
  {32'hbea3ddf9, 32'h00000000} /* (25, 6, 31) {real, imag} */,
  {32'hbf36b693, 32'h00000000} /* (25, 6, 30) {real, imag} */,
  {32'hbf522071, 32'h00000000} /* (25, 6, 29) {real, imag} */,
  {32'hbf98d29d, 32'h00000000} /* (25, 6, 28) {real, imag} */,
  {32'hbec80454, 32'h00000000} /* (25, 6, 27) {real, imag} */,
  {32'hbde6d5bb, 32'h00000000} /* (25, 6, 26) {real, imag} */,
  {32'hbf3bbcc6, 32'h00000000} /* (25, 6, 25) {real, imag} */,
  {32'hbf5720f5, 32'h00000000} /* (25, 6, 24) {real, imag} */,
  {32'hbf1c4be2, 32'h00000000} /* (25, 6, 23) {real, imag} */,
  {32'hbeff8fa7, 32'h00000000} /* (25, 6, 22) {real, imag} */,
  {32'hbed59272, 32'h00000000} /* (25, 6, 21) {real, imag} */,
  {32'h3ed2bbac, 32'h00000000} /* (25, 6, 20) {real, imag} */,
  {32'h3eaadd7b, 32'h00000000} /* (25, 6, 19) {real, imag} */,
  {32'h3f1b2de5, 32'h00000000} /* (25, 6, 18) {real, imag} */,
  {32'h3f18c698, 32'h00000000} /* (25, 6, 17) {real, imag} */,
  {32'h3ef3f307, 32'h00000000} /* (25, 6, 16) {real, imag} */,
  {32'h3f2a242a, 32'h00000000} /* (25, 6, 15) {real, imag} */,
  {32'h3f5e3821, 32'h00000000} /* (25, 6, 14) {real, imag} */,
  {32'h3f458e64, 32'h00000000} /* (25, 6, 13) {real, imag} */,
  {32'h3f764291, 32'h00000000} /* (25, 6, 12) {real, imag} */,
  {32'h3ea129d5, 32'h00000000} /* (25, 6, 11) {real, imag} */,
  {32'hbeac69d3, 32'h00000000} /* (25, 6, 10) {real, imag} */,
  {32'hbeeecd8c, 32'h00000000} /* (25, 6, 9) {real, imag} */,
  {32'hbe56d555, 32'h00000000} /* (25, 6, 8) {real, imag} */,
  {32'hbe604d3c, 32'h00000000} /* (25, 6, 7) {real, imag} */,
  {32'hbf26b72f, 32'h00000000} /* (25, 6, 6) {real, imag} */,
  {32'hbf7ef36c, 32'h00000000} /* (25, 6, 5) {real, imag} */,
  {32'hbf8383b5, 32'h00000000} /* (25, 6, 4) {real, imag} */,
  {32'hbf4c8174, 32'h00000000} /* (25, 6, 3) {real, imag} */,
  {32'hbf396043, 32'h00000000} /* (25, 6, 2) {real, imag} */,
  {32'hbf73d86c, 32'h00000000} /* (25, 6, 1) {real, imag} */,
  {32'hbe7818cb, 32'h00000000} /* (25, 6, 0) {real, imag} */,
  {32'hbf256a68, 32'h00000000} /* (25, 5, 31) {real, imag} */,
  {32'hbf89a12a, 32'h00000000} /* (25, 5, 30) {real, imag} */,
  {32'hbf5835e4, 32'h00000000} /* (25, 5, 29) {real, imag} */,
  {32'hbf83010a, 32'h00000000} /* (25, 5, 28) {real, imag} */,
  {32'hbeee1b68, 32'h00000000} /* (25, 5, 27) {real, imag} */,
  {32'hbe8e2452, 32'h00000000} /* (25, 5, 26) {real, imag} */,
  {32'hbf6a6c4b, 32'h00000000} /* (25, 5, 25) {real, imag} */,
  {32'hbf44cc9d, 32'h00000000} /* (25, 5, 24) {real, imag} */,
  {32'hbed51946, 32'h00000000} /* (25, 5, 23) {real, imag} */,
  {32'hbf078e78, 32'h00000000} /* (25, 5, 22) {real, imag} */,
  {32'hbf22c0ee, 32'h00000000} /* (25, 5, 21) {real, imag} */,
  {32'hbeaacf77, 32'h00000000} /* (25, 5, 20) {real, imag} */,
  {32'hbe974f46, 32'h00000000} /* (25, 5, 19) {real, imag} */,
  {32'hbea34762, 32'h00000000} /* (25, 5, 18) {real, imag} */,
  {32'hbe6060e3, 32'h00000000} /* (25, 5, 17) {real, imag} */,
  {32'h3e508260, 32'h00000000} /* (25, 5, 16) {real, imag} */,
  {32'h3f4133bf, 32'h00000000} /* (25, 5, 15) {real, imag} */,
  {32'h3f06aa6b, 32'h00000000} /* (25, 5, 14) {real, imag} */,
  {32'h3ef629d8, 32'h00000000} /* (25, 5, 13) {real, imag} */,
  {32'h3f3ce0a6, 32'h00000000} /* (25, 5, 12) {real, imag} */,
  {32'h3ecce2c5, 32'h00000000} /* (25, 5, 11) {real, imag} */,
  {32'h3e1bc7db, 32'h00000000} /* (25, 5, 10) {real, imag} */,
  {32'h3e22c08d, 32'h00000000} /* (25, 5, 9) {real, imag} */,
  {32'h3f215285, 32'h00000000} /* (25, 5, 8) {real, imag} */,
  {32'h3f34d8f1, 32'h00000000} /* (25, 5, 7) {real, imag} */,
  {32'hbd6d97be, 32'h00000000} /* (25, 5, 6) {real, imag} */,
  {32'hbf835ace, 32'h00000000} /* (25, 5, 5) {real, imag} */,
  {32'hbf4c2be5, 32'h00000000} /* (25, 5, 4) {real, imag} */,
  {32'hbf7018bf, 32'h00000000} /* (25, 5, 3) {real, imag} */,
  {32'hbf5db7bb, 32'h00000000} /* (25, 5, 2) {real, imag} */,
  {32'hbf91b6f2, 32'h00000000} /* (25, 5, 1) {real, imag} */,
  {32'hbee0ad7a, 32'h00000000} /* (25, 5, 0) {real, imag} */,
  {32'hbecc5bf0, 32'h00000000} /* (25, 4, 31) {real, imag} */,
  {32'hbf4d06df, 32'h00000000} /* (25, 4, 30) {real, imag} */,
  {32'hbf60851b, 32'h00000000} /* (25, 4, 29) {real, imag} */,
  {32'hbf7dadd4, 32'h00000000} /* (25, 4, 28) {real, imag} */,
  {32'hbf8fbbba, 32'h00000000} /* (25, 4, 27) {real, imag} */,
  {32'hbebac086, 32'h00000000} /* (25, 4, 26) {real, imag} */,
  {32'hbf154336, 32'h00000000} /* (25, 4, 25) {real, imag} */,
  {32'hbf72ea75, 32'h00000000} /* (25, 4, 24) {real, imag} */,
  {32'hbf53f1be, 32'h00000000} /* (25, 4, 23) {real, imag} */,
  {32'hbeeb3319, 32'h00000000} /* (25, 4, 22) {real, imag} */,
  {32'hbeebb074, 32'h00000000} /* (25, 4, 21) {real, imag} */,
  {32'hbf498649, 32'h00000000} /* (25, 4, 20) {real, imag} */,
  {32'hbf68d6b5, 32'h00000000} /* (25, 4, 19) {real, imag} */,
  {32'hbf5529f0, 32'h00000000} /* (25, 4, 18) {real, imag} */,
  {32'hbf7d5d24, 32'h00000000} /* (25, 4, 17) {real, imag} */,
  {32'hbf3a71be, 32'h00000000} /* (25, 4, 16) {real, imag} */,
  {32'h3f0cce84, 32'h00000000} /* (25, 4, 15) {real, imag} */,
  {32'h3ec919ac, 32'h00000000} /* (25, 4, 14) {real, imag} */,
  {32'h3ece9707, 32'h00000000} /* (25, 4, 13) {real, imag} */,
  {32'h3f08aadb, 32'h00000000} /* (25, 4, 12) {real, imag} */,
  {32'h3f423a17, 32'h00000000} /* (25, 4, 11) {real, imag} */,
  {32'h3f10c457, 32'h00000000} /* (25, 4, 10) {real, imag} */,
  {32'h3f04d9af, 32'h00000000} /* (25, 4, 9) {real, imag} */,
  {32'h3f9f7f98, 32'h00000000} /* (25, 4, 8) {real, imag} */,
  {32'h3f9b9449, 32'h00000000} /* (25, 4, 7) {real, imag} */,
  {32'h3f5dc725, 32'h00000000} /* (25, 4, 6) {real, imag} */,
  {32'hbe07753f, 32'h00000000} /* (25, 4, 5) {real, imag} */,
  {32'hbf315fa7, 32'h00000000} /* (25, 4, 4) {real, imag} */,
  {32'hbed4faa8, 32'h00000000} /* (25, 4, 3) {real, imag} */,
  {32'hbed31812, 32'h00000000} /* (25, 4, 2) {real, imag} */,
  {32'hbeeed9f5, 32'h00000000} /* (25, 4, 1) {real, imag} */,
  {32'hbe745f5b, 32'h00000000} /* (25, 4, 0) {real, imag} */,
  {32'hbe8a97fb, 32'h00000000} /* (25, 3, 31) {real, imag} */,
  {32'hbecca6a0, 32'h00000000} /* (25, 3, 30) {real, imag} */,
  {32'hbf71e6d0, 32'h00000000} /* (25, 3, 29) {real, imag} */,
  {32'hbfb59e1c, 32'h00000000} /* (25, 3, 28) {real, imag} */,
  {32'hbfcac34c, 32'h00000000} /* (25, 3, 27) {real, imag} */,
  {32'hbf199056, 32'h00000000} /* (25, 3, 26) {real, imag} */,
  {32'hbecdddcd, 32'h00000000} /* (25, 3, 25) {real, imag} */,
  {32'hbf74a983, 32'h00000000} /* (25, 3, 24) {real, imag} */,
  {32'hbf643eb1, 32'h00000000} /* (25, 3, 23) {real, imag} */,
  {32'hbf1fb5e9, 32'h00000000} /* (25, 3, 22) {real, imag} */,
  {32'hbf3cca51, 32'h00000000} /* (25, 3, 21) {real, imag} */,
  {32'hbf902253, 32'h00000000} /* (25, 3, 20) {real, imag} */,
  {32'hbf38b572, 32'h00000000} /* (25, 3, 19) {real, imag} */,
  {32'hbe49a0c6, 32'h00000000} /* (25, 3, 18) {real, imag} */,
  {32'hbf4c6b55, 32'h00000000} /* (25, 3, 17) {real, imag} */,
  {32'hbf84cd0b, 32'h00000000} /* (25, 3, 16) {real, imag} */,
  {32'h3dacee35, 32'h00000000} /* (25, 3, 15) {real, imag} */,
  {32'h3eff5453, 32'h00000000} /* (25, 3, 14) {real, imag} */,
  {32'h3f932671, 32'h00000000} /* (25, 3, 13) {real, imag} */,
  {32'h3f68a1c9, 32'h00000000} /* (25, 3, 12) {real, imag} */,
  {32'h3f95ba01, 32'h00000000} /* (25, 3, 11) {real, imag} */,
  {32'h3f556651, 32'h00000000} /* (25, 3, 10) {real, imag} */,
  {32'h3f23adb5, 32'h00000000} /* (25, 3, 9) {real, imag} */,
  {32'h3f994084, 32'h00000000} /* (25, 3, 8) {real, imag} */,
  {32'h3fdf0454, 32'h00000000} /* (25, 3, 7) {real, imag} */,
  {32'h3f8f9b1a, 32'h00000000} /* (25, 3, 6) {real, imag} */,
  {32'hbdf5e398, 32'h00000000} /* (25, 3, 5) {real, imag} */,
  {32'hbfa09e93, 32'h00000000} /* (25, 3, 4) {real, imag} */,
  {32'hbf25bc1c, 32'h00000000} /* (25, 3, 3) {real, imag} */,
  {32'hbed793e7, 32'h00000000} /* (25, 3, 2) {real, imag} */,
  {32'hbf482a3e, 32'h00000000} /* (25, 3, 1) {real, imag} */,
  {32'hbf0b5a9c, 32'h00000000} /* (25, 3, 0) {real, imag} */,
  {32'hbde4c5d6, 32'h00000000} /* (25, 2, 31) {real, imag} */,
  {32'hbf0b824f, 32'h00000000} /* (25, 2, 30) {real, imag} */,
  {32'hbf4aa0b5, 32'h00000000} /* (25, 2, 29) {real, imag} */,
  {32'hbfb2d6f8, 32'h00000000} /* (25, 2, 28) {real, imag} */,
  {32'hbfa2114e, 32'h00000000} /* (25, 2, 27) {real, imag} */,
  {32'hbef41adf, 32'h00000000} /* (25, 2, 26) {real, imag} */,
  {32'hbe356c6a, 32'h00000000} /* (25, 2, 25) {real, imag} */,
  {32'hbef2b234, 32'h00000000} /* (25, 2, 24) {real, imag} */,
  {32'hbf2e469a, 32'h00000000} /* (25, 2, 23) {real, imag} */,
  {32'hbf022f14, 32'h00000000} /* (25, 2, 22) {real, imag} */,
  {32'hbf635020, 32'h00000000} /* (25, 2, 21) {real, imag} */,
  {32'hbf986767, 32'h00000000} /* (25, 2, 20) {real, imag} */,
  {32'hbf60d264, 32'h00000000} /* (25, 2, 19) {real, imag} */,
  {32'hbf47089e, 32'h00000000} /* (25, 2, 18) {real, imag} */,
  {32'hbf0b1250, 32'h00000000} /* (25, 2, 17) {real, imag} */,
  {32'hbe272eda, 32'h00000000} /* (25, 2, 16) {real, imag} */,
  {32'h3f2c495f, 32'h00000000} /* (25, 2, 15) {real, imag} */,
  {32'h3f2f68c3, 32'h00000000} /* (25, 2, 14) {real, imag} */,
  {32'h3f69c6fe, 32'h00000000} /* (25, 2, 13) {real, imag} */,
  {32'h3f99ff76, 32'h00000000} /* (25, 2, 12) {real, imag} */,
  {32'h3f77ddaf, 32'h00000000} /* (25, 2, 11) {real, imag} */,
  {32'h3f6aa47a, 32'h00000000} /* (25, 2, 10) {real, imag} */,
  {32'h3f99625d, 32'h00000000} /* (25, 2, 9) {real, imag} */,
  {32'h3f49cf97, 32'h00000000} /* (25, 2, 8) {real, imag} */,
  {32'h3fb4f508, 32'h00000000} /* (25, 2, 7) {real, imag} */,
  {32'h3fb5660b, 32'h00000000} /* (25, 2, 6) {real, imag} */,
  {32'hbe3f33f0, 32'h00000000} /* (25, 2, 5) {real, imag} */,
  {32'hbfa45a72, 32'h00000000} /* (25, 2, 4) {real, imag} */,
  {32'hbf568c29, 32'h00000000} /* (25, 2, 3) {real, imag} */,
  {32'hbf010e8d, 32'h00000000} /* (25, 2, 2) {real, imag} */,
  {32'hbf0bae74, 32'h00000000} /* (25, 2, 1) {real, imag} */,
  {32'hbe941dcc, 32'h00000000} /* (25, 2, 0) {real, imag} */,
  {32'hbe254c47, 32'h00000000} /* (25, 1, 31) {real, imag} */,
  {32'hbf19fa54, 32'h00000000} /* (25, 1, 30) {real, imag} */,
  {32'hbf09130a, 32'h00000000} /* (25, 1, 29) {real, imag} */,
  {32'hbf9865c1, 32'h00000000} /* (25, 1, 28) {real, imag} */,
  {32'hbf709d3e, 32'h00000000} /* (25, 1, 27) {real, imag} */,
  {32'hbf299726, 32'h00000000} /* (25, 1, 26) {real, imag} */,
  {32'hbe95035d, 32'h00000000} /* (25, 1, 25) {real, imag} */,
  {32'hbe55ff7d, 32'h00000000} /* (25, 1, 24) {real, imag} */,
  {32'hbee40493, 32'h00000000} /* (25, 1, 23) {real, imag} */,
  {32'hbef23e5e, 32'h00000000} /* (25, 1, 22) {real, imag} */,
  {32'hbfa162da, 32'h00000000} /* (25, 1, 21) {real, imag} */,
  {32'hbf29f3b9, 32'h00000000} /* (25, 1, 20) {real, imag} */,
  {32'hbf49e9f3, 32'h00000000} /* (25, 1, 19) {real, imag} */,
  {32'hbf514f27, 32'h00000000} /* (25, 1, 18) {real, imag} */,
  {32'hbf603908, 32'h00000000} /* (25, 1, 17) {real, imag} */,
  {32'hbf2aaeb4, 32'h00000000} /* (25, 1, 16) {real, imag} */,
  {32'h3ed6e6ba, 32'h00000000} /* (25, 1, 15) {real, imag} */,
  {32'h3f229e29, 32'h00000000} /* (25, 1, 14) {real, imag} */,
  {32'h3d993144, 32'h00000000} /* (25, 1, 13) {real, imag} */,
  {32'h3ee6c77e, 32'h00000000} /* (25, 1, 12) {real, imag} */,
  {32'h3f761e0e, 32'h00000000} /* (25, 1, 11) {real, imag} */,
  {32'h3f5fe02f, 32'h00000000} /* (25, 1, 10) {real, imag} */,
  {32'h3f697b55, 32'h00000000} /* (25, 1, 9) {real, imag} */,
  {32'h3f79a8ef, 32'h00000000} /* (25, 1, 8) {real, imag} */,
  {32'h3f36f924, 32'h00000000} /* (25, 1, 7) {real, imag} */,
  {32'h3eb70e66, 32'h00000000} /* (25, 1, 6) {real, imag} */,
  {32'hbe267a6b, 32'h00000000} /* (25, 1, 5) {real, imag} */,
  {32'hbf0915ca, 32'h00000000} /* (25, 1, 4) {real, imag} */,
  {32'hbf0d41cc, 32'h00000000} /* (25, 1, 3) {real, imag} */,
  {32'hbf017174, 32'h00000000} /* (25, 1, 2) {real, imag} */,
  {32'hbeb1587a, 32'h00000000} /* (25, 1, 1) {real, imag} */,
  {32'hbded086f, 32'h00000000} /* (25, 1, 0) {real, imag} */,
  {32'hbd2cc680, 32'h00000000} /* (25, 0, 31) {real, imag} */,
  {32'hbdf68405, 32'h00000000} /* (25, 0, 30) {real, imag} */,
  {32'hbe4c0556, 32'h00000000} /* (25, 0, 29) {real, imag} */,
  {32'hbf07951b, 32'h00000000} /* (25, 0, 28) {real, imag} */,
  {32'hbf08f3f6, 32'h00000000} /* (25, 0, 27) {real, imag} */,
  {32'hbf0b7aab, 32'h00000000} /* (25, 0, 26) {real, imag} */,
  {32'hbe22dc9a, 32'h00000000} /* (25, 0, 25) {real, imag} */,
  {32'hbda318f5, 32'h00000000} /* (25, 0, 24) {real, imag} */,
  {32'hbe55529e, 32'h00000000} /* (25, 0, 23) {real, imag} */,
  {32'hbe9e23d3, 32'h00000000} /* (25, 0, 22) {real, imag} */,
  {32'hbeedd7ed, 32'h00000000} /* (25, 0, 21) {real, imag} */,
  {32'h3d499042, 32'h00000000} /* (25, 0, 20) {real, imag} */,
  {32'hbce9da51, 32'h00000000} /* (25, 0, 19) {real, imag} */,
  {32'hbdc0e3ec, 32'h00000000} /* (25, 0, 18) {real, imag} */,
  {32'hbecb4dd3, 32'h00000000} /* (25, 0, 17) {real, imag} */,
  {32'hbec6a2a3, 32'h00000000} /* (25, 0, 16) {real, imag} */,
  {32'h3c16af66, 32'h00000000} /* (25, 0, 15) {real, imag} */,
  {32'h3e78322f, 32'h00000000} /* (25, 0, 14) {real, imag} */,
  {32'h3e38f3a6, 32'h00000000} /* (25, 0, 13) {real, imag} */,
  {32'h3e95e0da, 32'h00000000} /* (25, 0, 12) {real, imag} */,
  {32'h3ed071db, 32'h00000000} /* (25, 0, 11) {real, imag} */,
  {32'h3e85c216, 32'h00000000} /* (25, 0, 10) {real, imag} */,
  {32'h3e3969c7, 32'h00000000} /* (25, 0, 9) {real, imag} */,
  {32'h3ef89094, 32'h00000000} /* (25, 0, 8) {real, imag} */,
  {32'h3e7f9d75, 32'h00000000} /* (25, 0, 7) {real, imag} */,
  {32'h3db54e69, 32'h00000000} /* (25, 0, 6) {real, imag} */,
  {32'hbdfe45fd, 32'h00000000} /* (25, 0, 5) {real, imag} */,
  {32'hbe9d84bf, 32'h00000000} /* (25, 0, 4) {real, imag} */,
  {32'hbef4e7e9, 32'h00000000} /* (25, 0, 3) {real, imag} */,
  {32'hbf4d62b4, 32'h00000000} /* (25, 0, 2) {real, imag} */,
  {32'hbf1f05e7, 32'h00000000} /* (25, 0, 1) {real, imag} */,
  {32'h3daa196e, 32'h00000000} /* (25, 0, 0) {real, imag} */,
  {32'hbe84c358, 32'h00000000} /* (24, 31, 31) {real, imag} */,
  {32'hbf520208, 32'h00000000} /* (24, 31, 30) {real, imag} */,
  {32'hbf4f7068, 32'h00000000} /* (24, 31, 29) {real, imag} */,
  {32'hbf420428, 32'h00000000} /* (24, 31, 28) {real, imag} */,
  {32'hbf85b58c, 32'h00000000} /* (24, 31, 27) {real, imag} */,
  {32'hbf12967f, 32'h00000000} /* (24, 31, 26) {real, imag} */,
  {32'hbec1bee9, 32'h00000000} /* (24, 31, 25) {real, imag} */,
  {32'hbedfc90a, 32'h00000000} /* (24, 31, 24) {real, imag} */,
  {32'hbeceae46, 32'h00000000} /* (24, 31, 23) {real, imag} */,
  {32'hbf3d8b9a, 32'h00000000} /* (24, 31, 22) {real, imag} */,
  {32'hbe73ee3b, 32'h00000000} /* (24, 31, 21) {real, imag} */,
  {32'h3f1ea6e7, 32'h00000000} /* (24, 31, 20) {real, imag} */,
  {32'h3f301344, 32'h00000000} /* (24, 31, 19) {real, imag} */,
  {32'h3efa197e, 32'h00000000} /* (24, 31, 18) {real, imag} */,
  {32'h3e9c18ae, 32'h00000000} /* (24, 31, 17) {real, imag} */,
  {32'h3eb67f8d, 32'h00000000} /* (24, 31, 16) {real, imag} */,
  {32'h3e8bae1f, 32'h00000000} /* (24, 31, 15) {real, imag} */,
  {32'h3ee44733, 32'h00000000} /* (24, 31, 14) {real, imag} */,
  {32'h3edefa3c, 32'h00000000} /* (24, 31, 13) {real, imag} */,
  {32'h3eadaa36, 32'h00000000} /* (24, 31, 12) {real, imag} */,
  {32'h3e72fd0b, 32'h00000000} /* (24, 31, 11) {real, imag} */,
  {32'hbf2e0daa, 32'h00000000} /* (24, 31, 10) {real, imag} */,
  {32'hbf0b3e85, 32'h00000000} /* (24, 31, 9) {real, imag} */,
  {32'hbf0e43ab, 32'h00000000} /* (24, 31, 8) {real, imag} */,
  {32'hbe3a8738, 32'h00000000} /* (24, 31, 7) {real, imag} */,
  {32'hbf1736d0, 32'h00000000} /* (24, 31, 6) {real, imag} */,
  {32'hbf6271da, 32'h00000000} /* (24, 31, 5) {real, imag} */,
  {32'hbf0f99c9, 32'h00000000} /* (24, 31, 4) {real, imag} */,
  {32'hbece2874, 32'h00000000} /* (24, 31, 3) {real, imag} */,
  {32'hbec960e8, 32'h00000000} /* (24, 31, 2) {real, imag} */,
  {32'hbf0737bc, 32'h00000000} /* (24, 31, 1) {real, imag} */,
  {32'hbe558dbf, 32'h00000000} /* (24, 31, 0) {real, imag} */,
  {32'hbe8b4c1e, 32'h00000000} /* (24, 30, 31) {real, imag} */,
  {32'hbf7724fd, 32'h00000000} /* (24, 30, 30) {real, imag} */,
  {32'hbf6f25a0, 32'h00000000} /* (24, 30, 29) {real, imag} */,
  {32'hbf55e98d, 32'h00000000} /* (24, 30, 28) {real, imag} */,
  {32'hbf830faa, 32'h00000000} /* (24, 30, 27) {real, imag} */,
  {32'hbf235ff7, 32'h00000000} /* (24, 30, 26) {real, imag} */,
  {32'hbf541d6a, 32'h00000000} /* (24, 30, 25) {real, imag} */,
  {32'hbf36ac8d, 32'h00000000} /* (24, 30, 24) {real, imag} */,
  {32'hbf10b861, 32'h00000000} /* (24, 30, 23) {real, imag} */,
  {32'hbf8616fe, 32'h00000000} /* (24, 30, 22) {real, imag} */,
  {32'hbe8d936b, 32'h00000000} /* (24, 30, 21) {real, imag} */,
  {32'h3f9467f9, 32'h00000000} /* (24, 30, 20) {real, imag} */,
  {32'h3f4745aa, 32'h00000000} /* (24, 30, 19) {real, imag} */,
  {32'h3f82a3e8, 32'h00000000} /* (24, 30, 18) {real, imag} */,
  {32'h3f8138c4, 32'h00000000} /* (24, 30, 17) {real, imag} */,
  {32'h3f8463c8, 32'h00000000} /* (24, 30, 16) {real, imag} */,
  {32'h3f3444f4, 32'h00000000} /* (24, 30, 15) {real, imag} */,
  {32'h3f5651f7, 32'h00000000} /* (24, 30, 14) {real, imag} */,
  {32'h3f2ff502, 32'h00000000} /* (24, 30, 13) {real, imag} */,
  {32'h3f64b651, 32'h00000000} /* (24, 30, 12) {real, imag} */,
  {32'h3f857401, 32'h00000000} /* (24, 30, 11) {real, imag} */,
  {32'hbebc1d4a, 32'h00000000} /* (24, 30, 10) {real, imag} */,
  {32'hbf3fd0a1, 32'h00000000} /* (24, 30, 9) {real, imag} */,
  {32'hbf894514, 32'h00000000} /* (24, 30, 8) {real, imag} */,
  {32'hbf604ae1, 32'h00000000} /* (24, 30, 7) {real, imag} */,
  {32'hbf8d64f1, 32'h00000000} /* (24, 30, 6) {real, imag} */,
  {32'hbf90c39e, 32'h00000000} /* (24, 30, 5) {real, imag} */,
  {32'hbf4000ef, 32'h00000000} /* (24, 30, 4) {real, imag} */,
  {32'hbf850eca, 32'h00000000} /* (24, 30, 3) {real, imag} */,
  {32'hbf2bb8c2, 32'h00000000} /* (24, 30, 2) {real, imag} */,
  {32'hbee27252, 32'h00000000} /* (24, 30, 1) {real, imag} */,
  {32'hbe521371, 32'h00000000} /* (24, 30, 0) {real, imag} */,
  {32'hbefbf66b, 32'h00000000} /* (24, 29, 31) {real, imag} */,
  {32'hbfab882d, 32'h00000000} /* (24, 29, 30) {real, imag} */,
  {32'hbf9814c4, 32'h00000000} /* (24, 29, 29) {real, imag} */,
  {32'hbf351e7c, 32'h00000000} /* (24, 29, 28) {real, imag} */,
  {32'hbf575140, 32'h00000000} /* (24, 29, 27) {real, imag} */,
  {32'hbf7c52ca, 32'h00000000} /* (24, 29, 26) {real, imag} */,
  {32'hbf9c5f9f, 32'h00000000} /* (24, 29, 25) {real, imag} */,
  {32'hbf37d257, 32'h00000000} /* (24, 29, 24) {real, imag} */,
  {32'hbed71056, 32'h00000000} /* (24, 29, 23) {real, imag} */,
  {32'hbf275c96, 32'h00000000} /* (24, 29, 22) {real, imag} */,
  {32'hbeb2493d, 32'h00000000} /* (24, 29, 21) {real, imag} */,
  {32'h3f576223, 32'h00000000} /* (24, 29, 20) {real, imag} */,
  {32'h3f23e305, 32'h00000000} /* (24, 29, 19) {real, imag} */,
  {32'h3f68dbe1, 32'h00000000} /* (24, 29, 18) {real, imag} */,
  {32'h3f61a2e4, 32'h00000000} /* (24, 29, 17) {real, imag} */,
  {32'h3f53ee90, 32'h00000000} /* (24, 29, 16) {real, imag} */,
  {32'h3f3e01f8, 32'h00000000} /* (24, 29, 15) {real, imag} */,
  {32'h3f445035, 32'h00000000} /* (24, 29, 14) {real, imag} */,
  {32'h3f15fc8f, 32'h00000000} /* (24, 29, 13) {real, imag} */,
  {32'h3f8269aa, 32'h00000000} /* (24, 29, 12) {real, imag} */,
  {32'h3f5981f8, 32'h00000000} /* (24, 29, 11) {real, imag} */,
  {32'hbd16b8b6, 32'h00000000} /* (24, 29, 10) {real, imag} */,
  {32'hbef6db90, 32'h00000000} /* (24, 29, 9) {real, imag} */,
  {32'hbf92de3a, 32'h00000000} /* (24, 29, 8) {real, imag} */,
  {32'hbfbcf260, 32'h00000000} /* (24, 29, 7) {real, imag} */,
  {32'hbf21fc7c, 32'h00000000} /* (24, 29, 6) {real, imag} */,
  {32'hbe7b88cd, 32'h00000000} /* (24, 29, 5) {real, imag} */,
  {32'hbc0da526, 32'h00000000} /* (24, 29, 4) {real, imag} */,
  {32'hbf82afef, 32'h00000000} /* (24, 29, 3) {real, imag} */,
  {32'hbf849226, 32'h00000000} /* (24, 29, 2) {real, imag} */,
  {32'hbf3d9d6b, 32'h00000000} /* (24, 29, 1) {real, imag} */,
  {32'hbecdad73, 32'h00000000} /* (24, 29, 0) {real, imag} */,
  {32'hbf54cd90, 32'h00000000} /* (24, 28, 31) {real, imag} */,
  {32'hbfbfa52d, 32'h00000000} /* (24, 28, 30) {real, imag} */,
  {32'hbfa8cbc0, 32'h00000000} /* (24, 28, 29) {real, imag} */,
  {32'hbf165c1b, 32'h00000000} /* (24, 28, 28) {real, imag} */,
  {32'hbf48e21b, 32'h00000000} /* (24, 28, 27) {real, imag} */,
  {32'hbfaaa4c9, 32'h00000000} /* (24, 28, 26) {real, imag} */,
  {32'hbf5b4322, 32'h00000000} /* (24, 28, 25) {real, imag} */,
  {32'hbf42a559, 32'h00000000} /* (24, 28, 24) {real, imag} */,
  {32'hbf6ae916, 32'h00000000} /* (24, 28, 23) {real, imag} */,
  {32'hbf88430f, 32'h00000000} /* (24, 28, 22) {real, imag} */,
  {32'hbf84942d, 32'h00000000} /* (24, 28, 21) {real, imag} */,
  {32'h3ec701c4, 32'h00000000} /* (24, 28, 20) {real, imag} */,
  {32'h3f6e8736, 32'h00000000} /* (24, 28, 19) {real, imag} */,
  {32'h3f93747c, 32'h00000000} /* (24, 28, 18) {real, imag} */,
  {32'h3f8402c5, 32'h00000000} /* (24, 28, 17) {real, imag} */,
  {32'h3fa7cdfa, 32'h00000000} /* (24, 28, 16) {real, imag} */,
  {32'h3f980312, 32'h00000000} /* (24, 28, 15) {real, imag} */,
  {32'h3f265d9c, 32'h00000000} /* (24, 28, 14) {real, imag} */,
  {32'h3f12a0de, 32'h00000000} /* (24, 28, 13) {real, imag} */,
  {32'h3f890563, 32'h00000000} /* (24, 28, 12) {real, imag} */,
  {32'h3f96ab98, 32'h00000000} /* (24, 28, 11) {real, imag} */,
  {32'hbeb4e789, 32'h00000000} /* (24, 28, 10) {real, imag} */,
  {32'hbf826fbf, 32'h00000000} /* (24, 28, 9) {real, imag} */,
  {32'hbf864433, 32'h00000000} /* (24, 28, 8) {real, imag} */,
  {32'hbf8c3a0e, 32'h00000000} /* (24, 28, 7) {real, imag} */,
  {32'hbf10b2ee, 32'h00000000} /* (24, 28, 6) {real, imag} */,
  {32'hbee5bf25, 32'h00000000} /* (24, 28, 5) {real, imag} */,
  {32'hbf48b821, 32'h00000000} /* (24, 28, 4) {real, imag} */,
  {32'hbfa9fb52, 32'h00000000} /* (24, 28, 3) {real, imag} */,
  {32'hbf947a2d, 32'h00000000} /* (24, 28, 2) {real, imag} */,
  {32'hbfa55b42, 32'h00000000} /* (24, 28, 1) {real, imag} */,
  {32'hbf6850e7, 32'h00000000} /* (24, 28, 0) {real, imag} */,
  {32'hbedfaaa8, 32'h00000000} /* (24, 27, 31) {real, imag} */,
  {32'hbf580cb8, 32'h00000000} /* (24, 27, 30) {real, imag} */,
  {32'hbf3723ed, 32'h00000000} /* (24, 27, 29) {real, imag} */,
  {32'hbe8a3b41, 32'h00000000} /* (24, 27, 28) {real, imag} */,
  {32'hbf593254, 32'h00000000} /* (24, 27, 27) {real, imag} */,
  {32'hc0061308, 32'h00000000} /* (24, 27, 26) {real, imag} */,
  {32'hbfbae4f4, 32'h00000000} /* (24, 27, 25) {real, imag} */,
  {32'hbf818c29, 32'h00000000} /* (24, 27, 24) {real, imag} */,
  {32'hbf66de9d, 32'h00000000} /* (24, 27, 23) {real, imag} */,
  {32'hbf322af4, 32'h00000000} /* (24, 27, 22) {real, imag} */,
  {32'hbf59d008, 32'h00000000} /* (24, 27, 21) {real, imag} */,
  {32'h3d32c091, 32'h00000000} /* (24, 27, 20) {real, imag} */,
  {32'h3f75ad76, 32'h00000000} /* (24, 27, 19) {real, imag} */,
  {32'h3fc38003, 32'h00000000} /* (24, 27, 18) {real, imag} */,
  {32'h3f875adf, 32'h00000000} /* (24, 27, 17) {real, imag} */,
  {32'h3f730c62, 32'h00000000} /* (24, 27, 16) {real, imag} */,
  {32'h3f3419e5, 32'h00000000} /* (24, 27, 15) {real, imag} */,
  {32'h3eb81b17, 32'h00000000} /* (24, 27, 14) {real, imag} */,
  {32'h3f4dda4a, 32'h00000000} /* (24, 27, 13) {real, imag} */,
  {32'h3f9c30ba, 32'h00000000} /* (24, 27, 12) {real, imag} */,
  {32'h3fa76019, 32'h00000000} /* (24, 27, 11) {real, imag} */,
  {32'hbed3caec, 32'h00000000} /* (24, 27, 10) {real, imag} */,
  {32'hbf9c86c3, 32'h00000000} /* (24, 27, 9) {real, imag} */,
  {32'hbf193762, 32'h00000000} /* (24, 27, 8) {real, imag} */,
  {32'hbe75466e, 32'h00000000} /* (24, 27, 7) {real, imag} */,
  {32'hbf0336d2, 32'h00000000} /* (24, 27, 6) {real, imag} */,
  {32'hbf5e54de, 32'h00000000} /* (24, 27, 5) {real, imag} */,
  {32'hbfb11430, 32'h00000000} /* (24, 27, 4) {real, imag} */,
  {32'hbfce44f2, 32'h00000000} /* (24, 27, 3) {real, imag} */,
  {32'hbf89d2bd, 32'h00000000} /* (24, 27, 2) {real, imag} */,
  {32'hbf4bbd53, 32'h00000000} /* (24, 27, 1) {real, imag} */,
  {32'hbeeec334, 32'h00000000} /* (24, 27, 0) {real, imag} */,
  {32'hbe6c20c6, 32'h00000000} /* (24, 26, 31) {real, imag} */,
  {32'hbf45d060, 32'h00000000} /* (24, 26, 30) {real, imag} */,
  {32'hbf6e5136, 32'h00000000} /* (24, 26, 29) {real, imag} */,
  {32'hbf11f350, 32'h00000000} /* (24, 26, 28) {real, imag} */,
  {32'hbf90561f, 32'h00000000} /* (24, 26, 27) {real, imag} */,
  {32'hbffaaa97, 32'h00000000} /* (24, 26, 26) {real, imag} */,
  {32'hbfc1153d, 32'h00000000} /* (24, 26, 25) {real, imag} */,
  {32'hbf4edfcc, 32'h00000000} /* (24, 26, 24) {real, imag} */,
  {32'hbf282b45, 32'h00000000} /* (24, 26, 23) {real, imag} */,
  {32'hbeedeae0, 32'h00000000} /* (24, 26, 22) {real, imag} */,
  {32'hbf13d023, 32'h00000000} /* (24, 26, 21) {real, imag} */,
  {32'h3eadfc61, 32'h00000000} /* (24, 26, 20) {real, imag} */,
  {32'h3f7cb623, 32'h00000000} /* (24, 26, 19) {real, imag} */,
  {32'h3fa7d035, 32'h00000000} /* (24, 26, 18) {real, imag} */,
  {32'h3f84aa8d, 32'h00000000} /* (24, 26, 17) {real, imag} */,
  {32'h3f510435, 32'h00000000} /* (24, 26, 16) {real, imag} */,
  {32'h3f3a3207, 32'h00000000} /* (24, 26, 15) {real, imag} */,
  {32'h3f415719, 32'h00000000} /* (24, 26, 14) {real, imag} */,
  {32'h3f175c7e, 32'h00000000} /* (24, 26, 13) {real, imag} */,
  {32'h3f4df44f, 32'h00000000} /* (24, 26, 12) {real, imag} */,
  {32'h3ea298bc, 32'h00000000} /* (24, 26, 11) {real, imag} */,
  {32'hbf2c2162, 32'h00000000} /* (24, 26, 10) {real, imag} */,
  {32'hbf6b6dde, 32'h00000000} /* (24, 26, 9) {real, imag} */,
  {32'hbec4f747, 32'h00000000} /* (24, 26, 8) {real, imag} */,
  {32'hbee42f0f, 32'h00000000} /* (24, 26, 7) {real, imag} */,
  {32'hbf0052d9, 32'h00000000} /* (24, 26, 6) {real, imag} */,
  {32'hbf24cf9f, 32'h00000000} /* (24, 26, 5) {real, imag} */,
  {32'hbf5d305a, 32'h00000000} /* (24, 26, 4) {real, imag} */,
  {32'hbf7b0050, 32'h00000000} /* (24, 26, 3) {real, imag} */,
  {32'hbf112754, 32'h00000000} /* (24, 26, 2) {real, imag} */,
  {32'hbe9ab349, 32'h00000000} /* (24, 26, 1) {real, imag} */,
  {32'hbe959ffe, 32'h00000000} /* (24, 26, 0) {real, imag} */,
  {32'hbee15aca, 32'h00000000} /* (24, 25, 31) {real, imag} */,
  {32'hbfa55b47, 32'h00000000} /* (24, 25, 30) {real, imag} */,
  {32'hbfd8d769, 32'h00000000} /* (24, 25, 29) {real, imag} */,
  {32'hbf7378a7, 32'h00000000} /* (24, 25, 28) {real, imag} */,
  {32'hbf805d50, 32'h00000000} /* (24, 25, 27) {real, imag} */,
  {32'hbf89a114, 32'h00000000} /* (24, 25, 26) {real, imag} */,
  {32'hbfa7ed79, 32'h00000000} /* (24, 25, 25) {real, imag} */,
  {32'hbf4b9532, 32'h00000000} /* (24, 25, 24) {real, imag} */,
  {32'hbef78eb6, 32'h00000000} /* (24, 25, 23) {real, imag} */,
  {32'hbe81f857, 32'h00000000} /* (24, 25, 22) {real, imag} */,
  {32'h3db95b77, 32'h00000000} /* (24, 25, 21) {real, imag} */,
  {32'h3f8e973d, 32'h00000000} /* (24, 25, 20) {real, imag} */,
  {32'h3f872645, 32'h00000000} /* (24, 25, 19) {real, imag} */,
  {32'h3f825904, 32'h00000000} /* (24, 25, 18) {real, imag} */,
  {32'h3f971638, 32'h00000000} /* (24, 25, 17) {real, imag} */,
  {32'h3f1bbe88, 32'h00000000} /* (24, 25, 16) {real, imag} */,
  {32'h3f156b47, 32'h00000000} /* (24, 25, 15) {real, imag} */,
  {32'h3f9fae0b, 32'h00000000} /* (24, 25, 14) {real, imag} */,
  {32'h3f60caef, 32'h00000000} /* (24, 25, 13) {real, imag} */,
  {32'h3eb7cd99, 32'h00000000} /* (24, 25, 12) {real, imag} */,
  {32'hbe24505e, 32'h00000000} /* (24, 25, 11) {real, imag} */,
  {32'hbf5222ff, 32'h00000000} /* (24, 25, 10) {real, imag} */,
  {32'hbf9086f6, 32'h00000000} /* (24, 25, 9) {real, imag} */,
  {32'hbf977c15, 32'h00000000} /* (24, 25, 8) {real, imag} */,
  {32'hbf5822d2, 32'h00000000} /* (24, 25, 7) {real, imag} */,
  {32'hbed77c42, 32'h00000000} /* (24, 25, 6) {real, imag} */,
  {32'hbf3519cf, 32'h00000000} /* (24, 25, 5) {real, imag} */,
  {32'hbfa5b510, 32'h00000000} /* (24, 25, 4) {real, imag} */,
  {32'hbf90eca7, 32'h00000000} /* (24, 25, 3) {real, imag} */,
  {32'hbefc2364, 32'h00000000} /* (24, 25, 2) {real, imag} */,
  {32'hbee07b11, 32'h00000000} /* (24, 25, 1) {real, imag} */,
  {32'hbf21a962, 32'h00000000} /* (24, 25, 0) {real, imag} */,
  {32'hbe7d611a, 32'h00000000} /* (24, 24, 31) {real, imag} */,
  {32'hbf2e568c, 32'h00000000} /* (24, 24, 30) {real, imag} */,
  {32'hbf691bf5, 32'h00000000} /* (24, 24, 29) {real, imag} */,
  {32'hbf4a4d6c, 32'h00000000} /* (24, 24, 28) {real, imag} */,
  {32'hbf06ebf6, 32'h00000000} /* (24, 24, 27) {real, imag} */,
  {32'hbf298305, 32'h00000000} /* (24, 24, 26) {real, imag} */,
  {32'hbf8a27bf, 32'h00000000} /* (24, 24, 25) {real, imag} */,
  {32'hbf63df73, 32'h00000000} /* (24, 24, 24) {real, imag} */,
  {32'hbf41f97e, 32'h00000000} /* (24, 24, 23) {real, imag} */,
  {32'hbf169365, 32'h00000000} /* (24, 24, 22) {real, imag} */,
  {32'hbed2bd5b, 32'h00000000} /* (24, 24, 21) {real, imag} */,
  {32'h3f02c368, 32'h00000000} /* (24, 24, 20) {real, imag} */,
  {32'h3eebad8a, 32'h00000000} /* (24, 24, 19) {real, imag} */,
  {32'h3f174b67, 32'h00000000} /* (24, 24, 18) {real, imag} */,
  {32'h3f770134, 32'h00000000} /* (24, 24, 17) {real, imag} */,
  {32'h3f495c7e, 32'h00000000} /* (24, 24, 16) {real, imag} */,
  {32'h3f4971a5, 32'h00000000} /* (24, 24, 15) {real, imag} */,
  {32'h3fabc5aa, 32'h00000000} /* (24, 24, 14) {real, imag} */,
  {32'h3f2e1aae, 32'h00000000} /* (24, 24, 13) {real, imag} */,
  {32'h3e01dcb4, 32'h00000000} /* (24, 24, 12) {real, imag} */,
  {32'h3da3dc0b, 32'h00000000} /* (24, 24, 11) {real, imag} */,
  {32'hbf2a7107, 32'h00000000} /* (24, 24, 10) {real, imag} */,
  {32'hbf8647a1, 32'h00000000} /* (24, 24, 9) {real, imag} */,
  {32'hbfa01c47, 32'h00000000} /* (24, 24, 8) {real, imag} */,
  {32'hbf54d9b1, 32'h00000000} /* (24, 24, 7) {real, imag} */,
  {32'hbe95025e, 32'h00000000} /* (24, 24, 6) {real, imag} */,
  {32'hbeba8434, 32'h00000000} /* (24, 24, 5) {real, imag} */,
  {32'hbf25ce5f, 32'h00000000} /* (24, 24, 4) {real, imag} */,
  {32'hbfa4a67a, 32'h00000000} /* (24, 24, 3) {real, imag} */,
  {32'hbf6be22a, 32'h00000000} /* (24, 24, 2) {real, imag} */,
  {32'hbf478367, 32'h00000000} /* (24, 24, 1) {real, imag} */,
  {32'hbf114d60, 32'h00000000} /* (24, 24, 0) {real, imag} */,
  {32'hbe761025, 32'h00000000} /* (24, 23, 31) {real, imag} */,
  {32'hbedad290, 32'h00000000} /* (24, 23, 30) {real, imag} */,
  {32'hbf488170, 32'h00000000} /* (24, 23, 29) {real, imag} */,
  {32'hbf3b67f4, 32'h00000000} /* (24, 23, 28) {real, imag} */,
  {32'hbf6b946f, 32'h00000000} /* (24, 23, 27) {real, imag} */,
  {32'hbf6f2063, 32'h00000000} /* (24, 23, 26) {real, imag} */,
  {32'hbf43c958, 32'h00000000} /* (24, 23, 25) {real, imag} */,
  {32'hbf398550, 32'h00000000} /* (24, 23, 24) {real, imag} */,
  {32'hbf9a421b, 32'h00000000} /* (24, 23, 23) {real, imag} */,
  {32'hbfb04bb3, 32'h00000000} /* (24, 23, 22) {real, imag} */,
  {32'hbeb57ff0, 32'h00000000} /* (24, 23, 21) {real, imag} */,
  {32'h3f321217, 32'h00000000} /* (24, 23, 20) {real, imag} */,
  {32'h3f45be02, 32'h00000000} /* (24, 23, 19) {real, imag} */,
  {32'h3f76f5e1, 32'h00000000} /* (24, 23, 18) {real, imag} */,
  {32'h3f86e334, 32'h00000000} /* (24, 23, 17) {real, imag} */,
  {32'h3f22e481, 32'h00000000} /* (24, 23, 16) {real, imag} */,
  {32'h3f824e57, 32'h00000000} /* (24, 23, 15) {real, imag} */,
  {32'h3fca30c3, 32'h00000000} /* (24, 23, 14) {real, imag} */,
  {32'h3f568ee3, 32'h00000000} /* (24, 23, 13) {real, imag} */,
  {32'h3f251da4, 32'h00000000} /* (24, 23, 12) {real, imag} */,
  {32'h3edfefd5, 32'h00000000} /* (24, 23, 11) {real, imag} */,
  {32'hbedc1fc0, 32'h00000000} /* (24, 23, 10) {real, imag} */,
  {32'hbf2f6360, 32'h00000000} /* (24, 23, 9) {real, imag} */,
  {32'hbf772eab, 32'h00000000} /* (24, 23, 8) {real, imag} */,
  {32'hbf80f78d, 32'h00000000} /* (24, 23, 7) {real, imag} */,
  {32'hbf34c503, 32'h00000000} /* (24, 23, 6) {real, imag} */,
  {32'hbf827505, 32'h00000000} /* (24, 23, 5) {real, imag} */,
  {32'hbf00704f, 32'h00000000} /* (24, 23, 4) {real, imag} */,
  {32'hbeb54531, 32'h00000000} /* (24, 23, 3) {real, imag} */,
  {32'hbf68c031, 32'h00000000} /* (24, 23, 2) {real, imag} */,
  {32'hbfb78acb, 32'h00000000} /* (24, 23, 1) {real, imag} */,
  {32'hbf49f16f, 32'h00000000} /* (24, 23, 0) {real, imag} */,
  {32'hbf3c97fc, 32'h00000000} /* (24, 22, 31) {real, imag} */,
  {32'hbf42b070, 32'h00000000} /* (24, 22, 30) {real, imag} */,
  {32'hbfa74f7c, 32'h00000000} /* (24, 22, 29) {real, imag} */,
  {32'hbf903389, 32'h00000000} /* (24, 22, 28) {real, imag} */,
  {32'hbf8060c2, 32'h00000000} /* (24, 22, 27) {real, imag} */,
  {32'hbf70e60d, 32'h00000000} /* (24, 22, 26) {real, imag} */,
  {32'hbf167d27, 32'h00000000} /* (24, 22, 25) {real, imag} */,
  {32'hbf670f26, 32'h00000000} /* (24, 22, 24) {real, imag} */,
  {32'hbf9e92d0, 32'h00000000} /* (24, 22, 23) {real, imag} */,
  {32'hbfb21a1e, 32'h00000000} /* (24, 22, 22) {real, imag} */,
  {32'hbe1d67fc, 32'h00000000} /* (24, 22, 21) {real, imag} */,
  {32'h3f871797, 32'h00000000} /* (24, 22, 20) {real, imag} */,
  {32'h3fef1eaf, 32'h00000000} /* (24, 22, 19) {real, imag} */,
  {32'h3fcad467, 32'h00000000} /* (24, 22, 18) {real, imag} */,
  {32'h3f808f6a, 32'h00000000} /* (24, 22, 17) {real, imag} */,
  {32'h3f4fb5ea, 32'h00000000} /* (24, 22, 16) {real, imag} */,
  {32'h3f4ec279, 32'h00000000} /* (24, 22, 15) {real, imag} */,
  {32'h3fa33603, 32'h00000000} /* (24, 22, 14) {real, imag} */,
  {32'h3fc07f5f, 32'h00000000} /* (24, 22, 13) {real, imag} */,
  {32'h3fa0ae70, 32'h00000000} /* (24, 22, 12) {real, imag} */,
  {32'h3f24edef, 32'h00000000} /* (24, 22, 11) {real, imag} */,
  {32'hbea47e28, 32'h00000000} /* (24, 22, 10) {real, imag} */,
  {32'hbf6a14c8, 32'h00000000} /* (24, 22, 9) {real, imag} */,
  {32'hbf7f0542, 32'h00000000} /* (24, 22, 8) {real, imag} */,
  {32'hbf9d8d54, 32'h00000000} /* (24, 22, 7) {real, imag} */,
  {32'hbf70a614, 32'h00000000} /* (24, 22, 6) {real, imag} */,
  {32'hbf7f9964, 32'h00000000} /* (24, 22, 5) {real, imag} */,
  {32'hbf340ec8, 32'h00000000} /* (24, 22, 4) {real, imag} */,
  {32'hbf27c63d, 32'h00000000} /* (24, 22, 3) {real, imag} */,
  {32'hbf21d0b7, 32'h00000000} /* (24, 22, 2) {real, imag} */,
  {32'hbf711907, 32'h00000000} /* (24, 22, 1) {real, imag} */,
  {32'hbf65b3db, 32'h00000000} /* (24, 22, 0) {real, imag} */,
  {32'hbe0d6bc9, 32'h00000000} /* (24, 21, 31) {real, imag} */,
  {32'hbec82169, 32'h00000000} /* (24, 21, 30) {real, imag} */,
  {32'hbf70085a, 32'h00000000} /* (24, 21, 29) {real, imag} */,
  {32'hbf17eef9, 32'h00000000} /* (24, 21, 28) {real, imag} */,
  {32'hbe66b3cb, 32'h00000000} /* (24, 21, 27) {real, imag} */,
  {32'hbd919edd, 32'h00000000} /* (24, 21, 26) {real, imag} */,
  {32'hbee310c6, 32'h00000000} /* (24, 21, 25) {real, imag} */,
  {32'hbf0f1379, 32'h00000000} /* (24, 21, 24) {real, imag} */,
  {32'hbe3ed088, 32'h00000000} /* (24, 21, 23) {real, imag} */,
  {32'hbd127411, 32'h00000000} /* (24, 21, 22) {real, imag} */,
  {32'hbd7d70f7, 32'h00000000} /* (24, 21, 21) {real, imag} */,
  {32'hbdb50ff2, 32'h00000000} /* (24, 21, 20) {real, imag} */,
  {32'h3f02dd4a, 32'h00000000} /* (24, 21, 19) {real, imag} */,
  {32'h3f3a9c68, 32'h00000000} /* (24, 21, 18) {real, imag} */,
  {32'h3f0987b9, 32'h00000000} /* (24, 21, 17) {real, imag} */,
  {32'h3f358fe7, 32'h00000000} /* (24, 21, 16) {real, imag} */,
  {32'h3e7a2cc5, 32'h00000000} /* (24, 21, 15) {real, imag} */,
  {32'h3f4039f1, 32'h00000000} /* (24, 21, 14) {real, imag} */,
  {32'h3f93716c, 32'h00000000} /* (24, 21, 13) {real, imag} */,
  {32'h3f73fd4f, 32'h00000000} /* (24, 21, 12) {real, imag} */,
  {32'hbdf5ffb5, 32'h00000000} /* (24, 21, 11) {real, imag} */,
  {32'hbee930ce, 32'h00000000} /* (24, 21, 10) {real, imag} */,
  {32'hbe92b1d8, 32'h00000000} /* (24, 21, 9) {real, imag} */,
  {32'hbeb322d7, 32'h00000000} /* (24, 21, 8) {real, imag} */,
  {32'hbf08760f, 32'h00000000} /* (24, 21, 7) {real, imag} */,
  {32'hbeb01d54, 32'h00000000} /* (24, 21, 6) {real, imag} */,
  {32'hbed72183, 32'h00000000} /* (24, 21, 5) {real, imag} */,
  {32'hbf3d1a8b, 32'h00000000} /* (24, 21, 4) {real, imag} */,
  {32'hbf2d6105, 32'h00000000} /* (24, 21, 3) {real, imag} */,
  {32'h3de53fbd, 32'h00000000} /* (24, 21, 2) {real, imag} */,
  {32'h3e5f6150, 32'h00000000} /* (24, 21, 1) {real, imag} */,
  {32'hbc95e2d4, 32'h00000000} /* (24, 21, 0) {real, imag} */,
  {32'h3f23aadd, 32'h00000000} /* (24, 20, 31) {real, imag} */,
  {32'h3f45cbb4, 32'h00000000} /* (24, 20, 30) {real, imag} */,
  {32'h3f0903df, 32'h00000000} /* (24, 20, 29) {real, imag} */,
  {32'h3eb8a95e, 32'h00000000} /* (24, 20, 28) {real, imag} */,
  {32'h3f6445df, 32'h00000000} /* (24, 20, 27) {real, imag} */,
  {32'h3fbcbc35, 32'h00000000} /* (24, 20, 26) {real, imag} */,
  {32'h3f201402, 32'h00000000} /* (24, 20, 25) {real, imag} */,
  {32'h3f19633c, 32'h00000000} /* (24, 20, 24) {real, imag} */,
  {32'h3fcedba3, 32'h00000000} /* (24, 20, 23) {real, imag} */,
  {32'h3fcbc20f, 32'h00000000} /* (24, 20, 22) {real, imag} */,
  {32'h3f49b00f, 32'h00000000} /* (24, 20, 21) {real, imag} */,
  {32'hbf6399c0, 32'h00000000} /* (24, 20, 20) {real, imag} */,
  {32'hbf84a352, 32'h00000000} /* (24, 20, 19) {real, imag} */,
  {32'hbf23cab6, 32'h00000000} /* (24, 20, 18) {real, imag} */,
  {32'hbf7c0595, 32'h00000000} /* (24, 20, 17) {real, imag} */,
  {32'hbf484afb, 32'h00000000} /* (24, 20, 16) {real, imag} */,
  {32'hbf4ecc3c, 32'h00000000} /* (24, 20, 15) {real, imag} */,
  {32'hbf010894, 32'h00000000} /* (24, 20, 14) {real, imag} */,
  {32'hbee68146, 32'h00000000} /* (24, 20, 13) {real, imag} */,
  {32'hbe9479c0, 32'h00000000} /* (24, 20, 12) {real, imag} */,
  {32'hbf5e5281, 32'h00000000} /* (24, 20, 11) {real, imag} */,
  {32'hbdf4360d, 32'h00000000} /* (24, 20, 10) {real, imag} */,
  {32'h3f73cc97, 32'h00000000} /* (24, 20, 9) {real, imag} */,
  {32'h3f1955ac, 32'h00000000} /* (24, 20, 8) {real, imag} */,
  {32'h3f0254c8, 32'h00000000} /* (24, 20, 7) {real, imag} */,
  {32'h3f50f1a5, 32'h00000000} /* (24, 20, 6) {real, imag} */,
  {32'h3f1d3a30, 32'h00000000} /* (24, 20, 5) {real, imag} */,
  {32'h3f233fbb, 32'h00000000} /* (24, 20, 4) {real, imag} */,
  {32'h3ecedfa2, 32'h00000000} /* (24, 20, 3) {real, imag} */,
  {32'h3f2bb965, 32'h00000000} /* (24, 20, 2) {real, imag} */,
  {32'h3f8626dc, 32'h00000000} /* (24, 20, 1) {real, imag} */,
  {32'h3f3013ff, 32'h00000000} /* (24, 20, 0) {real, imag} */,
  {32'h3f0ad7a0, 32'h00000000} /* (24, 19, 31) {real, imag} */,
  {32'h3f7c3b14, 32'h00000000} /* (24, 19, 30) {real, imag} */,
  {32'h3f4c279b, 32'h00000000} /* (24, 19, 29) {real, imag} */,
  {32'h3ef265a8, 32'h00000000} /* (24, 19, 28) {real, imag} */,
  {32'h3f6084e3, 32'h00000000} /* (24, 19, 27) {real, imag} */,
  {32'h3f9f21ec, 32'h00000000} /* (24, 19, 26) {real, imag} */,
  {32'h3f442bb7, 32'h00000000} /* (24, 19, 25) {real, imag} */,
  {32'h3f4b0d83, 32'h00000000} /* (24, 19, 24) {real, imag} */,
  {32'h3fac386e, 32'h00000000} /* (24, 19, 23) {real, imag} */,
  {32'h3fbdbbab, 32'h00000000} /* (24, 19, 22) {real, imag} */,
  {32'h3f8000b2, 32'h00000000} /* (24, 19, 21) {real, imag} */,
  {32'hbf3fa187, 32'h00000000} /* (24, 19, 20) {real, imag} */,
  {32'hbf83d6c4, 32'h00000000} /* (24, 19, 19) {real, imag} */,
  {32'hbf8c4142, 32'h00000000} /* (24, 19, 18) {real, imag} */,
  {32'hbf8b61aa, 32'h00000000} /* (24, 19, 17) {real, imag} */,
  {32'hbf4cf3b2, 32'h00000000} /* (24, 19, 16) {real, imag} */,
  {32'hbf11762d, 32'h00000000} /* (24, 19, 15) {real, imag} */,
  {32'hbef2bcc8, 32'h00000000} /* (24, 19, 14) {real, imag} */,
  {32'hbf33dba2, 32'h00000000} /* (24, 19, 13) {real, imag} */,
  {32'hbf6d4ed3, 32'h00000000} /* (24, 19, 12) {real, imag} */,
  {32'hbf373b99, 32'h00000000} /* (24, 19, 11) {real, imag} */,
  {32'h3f3f61e8, 32'h00000000} /* (24, 19, 10) {real, imag} */,
  {32'h3f9be328, 32'h00000000} /* (24, 19, 9) {real, imag} */,
  {32'h3f3c62ed, 32'h00000000} /* (24, 19, 8) {real, imag} */,
  {32'h3f5398cc, 32'h00000000} /* (24, 19, 7) {real, imag} */,
  {32'h3f9338f6, 32'h00000000} /* (24, 19, 6) {real, imag} */,
  {32'h3f7bb6c2, 32'h00000000} /* (24, 19, 5) {real, imag} */,
  {32'h3f45e3a4, 32'h00000000} /* (24, 19, 4) {real, imag} */,
  {32'h3ebc3f08, 32'h00000000} /* (24, 19, 3) {real, imag} */,
  {32'h3f24bc92, 32'h00000000} /* (24, 19, 2) {real, imag} */,
  {32'h3f64fc41, 32'h00000000} /* (24, 19, 1) {real, imag} */,
  {32'h3eb9c925, 32'h00000000} /* (24, 19, 0) {real, imag} */,
  {32'h3f5d6ce2, 32'h00000000} /* (24, 18, 31) {real, imag} */,
  {32'h3f9b9f9b, 32'h00000000} /* (24, 18, 30) {real, imag} */,
  {32'h3f8110a9, 32'h00000000} /* (24, 18, 29) {real, imag} */,
  {32'h3f1fe94f, 32'h00000000} /* (24, 18, 28) {real, imag} */,
  {32'h3efba2e2, 32'h00000000} /* (24, 18, 27) {real, imag} */,
  {32'h3ee5434d, 32'h00000000} /* (24, 18, 26) {real, imag} */,
  {32'h3f71980b, 32'h00000000} /* (24, 18, 25) {real, imag} */,
  {32'h3f6d5411, 32'h00000000} /* (24, 18, 24) {real, imag} */,
  {32'h3f209661, 32'h00000000} /* (24, 18, 23) {real, imag} */,
  {32'h3f8ee229, 32'h00000000} /* (24, 18, 22) {real, imag} */,
  {32'h3f9bef52, 32'h00000000} /* (24, 18, 21) {real, imag} */,
  {32'hbf36156e, 32'h00000000} /* (24, 18, 20) {real, imag} */,
  {32'hbf92bf71, 32'h00000000} /* (24, 18, 19) {real, imag} */,
  {32'hbf877791, 32'h00000000} /* (24, 18, 18) {real, imag} */,
  {32'hbf87aa34, 32'h00000000} /* (24, 18, 17) {real, imag} */,
  {32'hbe0c2605, 32'h00000000} /* (24, 18, 16) {real, imag} */,
  {32'hbed0de7e, 32'h00000000} /* (24, 18, 15) {real, imag} */,
  {32'hbf3f16a5, 32'h00000000} /* (24, 18, 14) {real, imag} */,
  {32'hbef97738, 32'h00000000} /* (24, 18, 13) {real, imag} */,
  {32'hbef95a9c, 32'h00000000} /* (24, 18, 12) {real, imag} */,
  {32'hbebb371b, 32'h00000000} /* (24, 18, 11) {real, imag} */,
  {32'h3f723c0e, 32'h00000000} /* (24, 18, 10) {real, imag} */,
  {32'h3f880453, 32'h00000000} /* (24, 18, 9) {real, imag} */,
  {32'h3f070911, 32'h00000000} /* (24, 18, 8) {real, imag} */,
  {32'h3f17ded2, 32'h00000000} /* (24, 18, 7) {real, imag} */,
  {32'h3f36ca1b, 32'h00000000} /* (24, 18, 6) {real, imag} */,
  {32'h3f26b208, 32'h00000000} /* (24, 18, 5) {real, imag} */,
  {32'h3eaafff8, 32'h00000000} /* (24, 18, 4) {real, imag} */,
  {32'h3eb23438, 32'h00000000} /* (24, 18, 3) {real, imag} */,
  {32'h3f2187f7, 32'h00000000} /* (24, 18, 2) {real, imag} */,
  {32'h3f86a728, 32'h00000000} /* (24, 18, 1) {real, imag} */,
  {32'h3f3ea42f, 32'h00000000} /* (24, 18, 0) {real, imag} */,
  {32'h3f6059dc, 32'h00000000} /* (24, 17, 31) {real, imag} */,
  {32'h3f6a19ea, 32'h00000000} /* (24, 17, 30) {real, imag} */,
  {32'h3f42bbc7, 32'h00000000} /* (24, 17, 29) {real, imag} */,
  {32'h3f575622, 32'h00000000} /* (24, 17, 28) {real, imag} */,
  {32'h3f5d5a3f, 32'h00000000} /* (24, 17, 27) {real, imag} */,
  {32'h3eb32111, 32'h00000000} /* (24, 17, 26) {real, imag} */,
  {32'h3f52453f, 32'h00000000} /* (24, 17, 25) {real, imag} */,
  {32'h3f90ea97, 32'h00000000} /* (24, 17, 24) {real, imag} */,
  {32'h3f8b3323, 32'h00000000} /* (24, 17, 23) {real, imag} */,
  {32'h3f64630a, 32'h00000000} /* (24, 17, 22) {real, imag} */,
  {32'h3f380a08, 32'h00000000} /* (24, 17, 21) {real, imag} */,
  {32'hbf207d23, 32'h00000000} /* (24, 17, 20) {real, imag} */,
  {32'hbf63362c, 32'h00000000} /* (24, 17, 19) {real, imag} */,
  {32'hbf14ad49, 32'h00000000} /* (24, 17, 18) {real, imag} */,
  {32'hbf4fd54e, 32'h00000000} /* (24, 17, 17) {real, imag} */,
  {32'hbf063fae, 32'h00000000} /* (24, 17, 16) {real, imag} */,
  {32'hbf566b30, 32'h00000000} /* (24, 17, 15) {real, imag} */,
  {32'hbf8db4d2, 32'h00000000} /* (24, 17, 14) {real, imag} */,
  {32'hbf4537ca, 32'h00000000} /* (24, 17, 13) {real, imag} */,
  {32'hbf3f4182, 32'h00000000} /* (24, 17, 12) {real, imag} */,
  {32'hbf2a71f0, 32'h00000000} /* (24, 17, 11) {real, imag} */,
  {32'h3dc58199, 32'h00000000} /* (24, 17, 10) {real, imag} */,
  {32'h3f0f12b8, 32'h00000000} /* (24, 17, 9) {real, imag} */,
  {32'h3e3521a8, 32'h00000000} /* (24, 17, 8) {real, imag} */,
  {32'h3eeff6ac, 32'h00000000} /* (24, 17, 7) {real, imag} */,
  {32'h3f049ef4, 32'h00000000} /* (24, 17, 6) {real, imag} */,
  {32'h3ee68211, 32'h00000000} /* (24, 17, 5) {real, imag} */,
  {32'h3effb19a, 32'h00000000} /* (24, 17, 4) {real, imag} */,
  {32'h3f199d43, 32'h00000000} /* (24, 17, 3) {real, imag} */,
  {32'h3f1f501d, 32'h00000000} /* (24, 17, 2) {real, imag} */,
  {32'h3f97c296, 32'h00000000} /* (24, 17, 1) {real, imag} */,
  {32'h3fa927c7, 32'h00000000} /* (24, 17, 0) {real, imag} */,
  {32'h3f38050b, 32'h00000000} /* (24, 16, 31) {real, imag} */,
  {32'h3f9429a0, 32'h00000000} /* (24, 16, 30) {real, imag} */,
  {32'h3f5c68fc, 32'h00000000} /* (24, 16, 29) {real, imag} */,
  {32'h3f01b644, 32'h00000000} /* (24, 16, 28) {real, imag} */,
  {32'h3eca2b7d, 32'h00000000} /* (24, 16, 27) {real, imag} */,
  {32'h3e42a304, 32'h00000000} /* (24, 16, 26) {real, imag} */,
  {32'h3f15cbbe, 32'h00000000} /* (24, 16, 25) {real, imag} */,
  {32'h3f7b1f40, 32'h00000000} /* (24, 16, 24) {real, imag} */,
  {32'h3f9e52f8, 32'h00000000} /* (24, 16, 23) {real, imag} */,
  {32'h3f8637fc, 32'h00000000} /* (24, 16, 22) {real, imag} */,
  {32'h3ed02748, 32'h00000000} /* (24, 16, 21) {real, imag} */,
  {32'hbf79b91f, 32'h00000000} /* (24, 16, 20) {real, imag} */,
  {32'hbf928782, 32'h00000000} /* (24, 16, 19) {real, imag} */,
  {32'hbe88d4c7, 32'h00000000} /* (24, 16, 18) {real, imag} */,
  {32'hbe872afe, 32'h00000000} /* (24, 16, 17) {real, imag} */,
  {32'hbf380059, 32'h00000000} /* (24, 16, 16) {real, imag} */,
  {32'hbf1803c4, 32'h00000000} /* (24, 16, 15) {real, imag} */,
  {32'hbf70ad85, 32'h00000000} /* (24, 16, 14) {real, imag} */,
  {32'hbf898faf, 32'h00000000} /* (24, 16, 13) {real, imag} */,
  {32'hbfbdb29a, 32'h00000000} /* (24, 16, 12) {real, imag} */,
  {32'hbf5a654b, 32'h00000000} /* (24, 16, 11) {real, imag} */,
  {32'h3e2a8ec2, 32'h00000000} /* (24, 16, 10) {real, imag} */,
  {32'h3f13b42e, 32'h00000000} /* (24, 16, 9) {real, imag} */,
  {32'h3e729cd0, 32'h00000000} /* (24, 16, 8) {real, imag} */,
  {32'h3f3cc888, 32'h00000000} /* (24, 16, 7) {real, imag} */,
  {32'h3f738589, 32'h00000000} /* (24, 16, 6) {real, imag} */,
  {32'h3f86fdcb, 32'h00000000} /* (24, 16, 5) {real, imag} */,
  {32'h3f901a7b, 32'h00000000} /* (24, 16, 4) {real, imag} */,
  {32'h3f6c9bad, 32'h00000000} /* (24, 16, 3) {real, imag} */,
  {32'h3f8e00c5, 32'h00000000} /* (24, 16, 2) {real, imag} */,
  {32'h3fa412d7, 32'h00000000} /* (24, 16, 1) {real, imag} */,
  {32'h3f873e59, 32'h00000000} /* (24, 16, 0) {real, imag} */,
  {32'h3ef97f9b, 32'h00000000} /* (24, 15, 31) {real, imag} */,
  {32'h3f69242e, 32'h00000000} /* (24, 15, 30) {real, imag} */,
  {32'h3f472981, 32'h00000000} /* (24, 15, 29) {real, imag} */,
  {32'h3f3988bf, 32'h00000000} /* (24, 15, 28) {real, imag} */,
  {32'h3f2ef735, 32'h00000000} /* (24, 15, 27) {real, imag} */,
  {32'h3efad8bd, 32'h00000000} /* (24, 15, 26) {real, imag} */,
  {32'h3e5241ce, 32'h00000000} /* (24, 15, 25) {real, imag} */,
  {32'h3ee41ea3, 32'h00000000} /* (24, 15, 24) {real, imag} */,
  {32'h3f818bc7, 32'h00000000} /* (24, 15, 23) {real, imag} */,
  {32'h3f0ef8c3, 32'h00000000} /* (24, 15, 22) {real, imag} */,
  {32'h3dff0085, 32'h00000000} /* (24, 15, 21) {real, imag} */,
  {32'hbf2f036c, 32'h00000000} /* (24, 15, 20) {real, imag} */,
  {32'hbf790ce3, 32'h00000000} /* (24, 15, 19) {real, imag} */,
  {32'hbe67e1f7, 32'h00000000} /* (24, 15, 18) {real, imag} */,
  {32'hbea6a052, 32'h00000000} /* (24, 15, 17) {real, imag} */,
  {32'hbf43363f, 32'h00000000} /* (24, 15, 16) {real, imag} */,
  {32'hbf0f3f2b, 32'h00000000} /* (24, 15, 15) {real, imag} */,
  {32'hbf68959f, 32'h00000000} /* (24, 15, 14) {real, imag} */,
  {32'hbf69eb4a, 32'h00000000} /* (24, 15, 13) {real, imag} */,
  {32'hbf88315f, 32'h00000000} /* (24, 15, 12) {real, imag} */,
  {32'hbf00ceae, 32'h00000000} /* (24, 15, 11) {real, imag} */,
  {32'h3e9a0683, 32'h00000000} /* (24, 15, 10) {real, imag} */,
  {32'h3eb2ef6e, 32'h00000000} /* (24, 15, 9) {real, imag} */,
  {32'h3ea05af7, 32'h00000000} /* (24, 15, 8) {real, imag} */,
  {32'h3efa84d2, 32'h00000000} /* (24, 15, 7) {real, imag} */,
  {32'h3f12190f, 32'h00000000} /* (24, 15, 6) {real, imag} */,
  {32'h3f3dadf9, 32'h00000000} /* (24, 15, 5) {real, imag} */,
  {32'h3f4a117c, 32'h00000000} /* (24, 15, 4) {real, imag} */,
  {32'h3f89b475, 32'h00000000} /* (24, 15, 3) {real, imag} */,
  {32'h3f88838d, 32'h00000000} /* (24, 15, 2) {real, imag} */,
  {32'h3f454018, 32'h00000000} /* (24, 15, 1) {real, imag} */,
  {32'h3f05590e, 32'h00000000} /* (24, 15, 0) {real, imag} */,
  {32'h3f0e6333, 32'h00000000} /* (24, 14, 31) {real, imag} */,
  {32'h3f20412c, 32'h00000000} /* (24, 14, 30) {real, imag} */,
  {32'h3f0d0f5b, 32'h00000000} /* (24, 14, 29) {real, imag} */,
  {32'h3f48516e, 32'h00000000} /* (24, 14, 28) {real, imag} */,
  {32'h3f50b7c7, 32'h00000000} /* (24, 14, 27) {real, imag} */,
  {32'h3f445bb5, 32'h00000000} /* (24, 14, 26) {real, imag} */,
  {32'h3eeb1fc3, 32'h00000000} /* (24, 14, 25) {real, imag} */,
  {32'h3f758f58, 32'h00000000} /* (24, 14, 24) {real, imag} */,
  {32'h3fdb20fa, 32'h00000000} /* (24, 14, 23) {real, imag} */,
  {32'h3f74739b, 32'h00000000} /* (24, 14, 22) {real, imag} */,
  {32'h3e8963d4, 32'h00000000} /* (24, 14, 21) {real, imag} */,
  {32'hbed13874, 32'h00000000} /* (24, 14, 20) {real, imag} */,
  {32'hbf82b914, 32'h00000000} /* (24, 14, 19) {real, imag} */,
  {32'hbf28bf4d, 32'h00000000} /* (24, 14, 18) {real, imag} */,
  {32'hbf59cb16, 32'h00000000} /* (24, 14, 17) {real, imag} */,
  {32'hbf756230, 32'h00000000} /* (24, 14, 16) {real, imag} */,
  {32'hbf18c915, 32'h00000000} /* (24, 14, 15) {real, imag} */,
  {32'hbf2adebe, 32'h00000000} /* (24, 14, 14) {real, imag} */,
  {32'hbf4edecf, 32'h00000000} /* (24, 14, 13) {real, imag} */,
  {32'hbf2df915, 32'h00000000} /* (24, 14, 12) {real, imag} */,
  {32'hbf252e20, 32'h00000000} /* (24, 14, 11) {real, imag} */,
  {32'h3e0bc0c8, 32'h00000000} /* (24, 14, 10) {real, imag} */,
  {32'h3f1f9fef, 32'h00000000} /* (24, 14, 9) {real, imag} */,
  {32'h3f801f6f, 32'h00000000} /* (24, 14, 8) {real, imag} */,
  {32'h3f3a617e, 32'h00000000} /* (24, 14, 7) {real, imag} */,
  {32'h3f27dca6, 32'h00000000} /* (24, 14, 6) {real, imag} */,
  {32'h3f9b10a4, 32'h00000000} /* (24, 14, 5) {real, imag} */,
  {32'h3f999083, 32'h00000000} /* (24, 14, 4) {real, imag} */,
  {32'h3f6ffe7b, 32'h00000000} /* (24, 14, 3) {real, imag} */,
  {32'h3f0e8ce0, 32'h00000000} /* (24, 14, 2) {real, imag} */,
  {32'h3f0a1591, 32'h00000000} /* (24, 14, 1) {real, imag} */,
  {32'h3efc3110, 32'h00000000} /* (24, 14, 0) {real, imag} */,
  {32'h3ef72d9b, 32'h00000000} /* (24, 13, 31) {real, imag} */,
  {32'h3f207267, 32'h00000000} /* (24, 13, 30) {real, imag} */,
  {32'h3f44a968, 32'h00000000} /* (24, 13, 29) {real, imag} */,
  {32'h3fb01fb2, 32'h00000000} /* (24, 13, 28) {real, imag} */,
  {32'h3fa13752, 32'h00000000} /* (24, 13, 27) {real, imag} */,
  {32'h3f42d729, 32'h00000000} /* (24, 13, 26) {real, imag} */,
  {32'h3f05a5ad, 32'h00000000} /* (24, 13, 25) {real, imag} */,
  {32'h3f9fea19, 32'h00000000} /* (24, 13, 24) {real, imag} */,
  {32'h3fe3a46a, 32'h00000000} /* (24, 13, 23) {real, imag} */,
  {32'h3f53836b, 32'h00000000} /* (24, 13, 22) {real, imag} */,
  {32'h3eba5e36, 32'h00000000} /* (24, 13, 21) {real, imag} */,
  {32'hbee0d9dc, 32'h00000000} /* (24, 13, 20) {real, imag} */,
  {32'hbf91c2d1, 32'h00000000} /* (24, 13, 19) {real, imag} */,
  {32'hbf926132, 32'h00000000} /* (24, 13, 18) {real, imag} */,
  {32'hbf5b2d5d, 32'h00000000} /* (24, 13, 17) {real, imag} */,
  {32'hbf1db0e4, 32'h00000000} /* (24, 13, 16) {real, imag} */,
  {32'hbf279ab3, 32'h00000000} /* (24, 13, 15) {real, imag} */,
  {32'hbf102990, 32'h00000000} /* (24, 13, 14) {real, imag} */,
  {32'hbf49d190, 32'h00000000} /* (24, 13, 13) {real, imag} */,
  {32'hbf509094, 32'h00000000} /* (24, 13, 12) {real, imag} */,
  {32'hbf647e3b, 32'h00000000} /* (24, 13, 11) {real, imag} */,
  {32'h3ec66ff0, 32'h00000000} /* (24, 13, 10) {real, imag} */,
  {32'h3f44466f, 32'h00000000} /* (24, 13, 9) {real, imag} */,
  {32'h3f82ab18, 32'h00000000} /* (24, 13, 8) {real, imag} */,
  {32'h3f64d681, 32'h00000000} /* (24, 13, 7) {real, imag} */,
  {32'h3f8e3496, 32'h00000000} /* (24, 13, 6) {real, imag} */,
  {32'h3fd5d249, 32'h00000000} /* (24, 13, 5) {real, imag} */,
  {32'h3fb39294, 32'h00000000} /* (24, 13, 4) {real, imag} */,
  {32'h3f6a4d84, 32'h00000000} /* (24, 13, 3) {real, imag} */,
  {32'h3e84708a, 32'h00000000} /* (24, 13, 2) {real, imag} */,
  {32'h3ee8f040, 32'h00000000} /* (24, 13, 1) {real, imag} */,
  {32'h3ef15e0e, 32'h00000000} /* (24, 13, 0) {real, imag} */,
  {32'h3ef31127, 32'h00000000} /* (24, 12, 31) {real, imag} */,
  {32'h3f5fedc7, 32'h00000000} /* (24, 12, 30) {real, imag} */,
  {32'h3f0fb496, 32'h00000000} /* (24, 12, 29) {real, imag} */,
  {32'h3f90d4e9, 32'h00000000} /* (24, 12, 28) {real, imag} */,
  {32'h3fa70312, 32'h00000000} /* (24, 12, 27) {real, imag} */,
  {32'h3f957d21, 32'h00000000} /* (24, 12, 26) {real, imag} */,
  {32'h3f70d976, 32'h00000000} /* (24, 12, 25) {real, imag} */,
  {32'h3f93b61b, 32'h00000000} /* (24, 12, 24) {real, imag} */,
  {32'h3f800eb2, 32'h00000000} /* (24, 12, 23) {real, imag} */,
  {32'h3f0957c9, 32'h00000000} /* (24, 12, 22) {real, imag} */,
  {32'h3dc82c16, 32'h00000000} /* (24, 12, 21) {real, imag} */,
  {32'hbf3d8494, 32'h00000000} /* (24, 12, 20) {real, imag} */,
  {32'hbfc4775a, 32'h00000000} /* (24, 12, 19) {real, imag} */,
  {32'hbfef6abe, 32'h00000000} /* (24, 12, 18) {real, imag} */,
  {32'hbfc4d850, 32'h00000000} /* (24, 12, 17) {real, imag} */,
  {32'hbf8a849a, 32'h00000000} /* (24, 12, 16) {real, imag} */,
  {32'hbf9e23c2, 32'h00000000} /* (24, 12, 15) {real, imag} */,
  {32'hbeddd0fd, 32'h00000000} /* (24, 12, 14) {real, imag} */,
  {32'hbf13a561, 32'h00000000} /* (24, 12, 13) {real, imag} */,
  {32'hbf628c0d, 32'h00000000} /* (24, 12, 12) {real, imag} */,
  {32'hbf80ad24, 32'h00000000} /* (24, 12, 11) {real, imag} */,
  {32'h3f7125e3, 32'h00000000} /* (24, 12, 10) {real, imag} */,
  {32'h3f97abf9, 32'h00000000} /* (24, 12, 9) {real, imag} */,
  {32'h3fa203d7, 32'h00000000} /* (24, 12, 8) {real, imag} */,
  {32'h3f5dbc11, 32'h00000000} /* (24, 12, 7) {real, imag} */,
  {32'h3f9e5714, 32'h00000000} /* (24, 12, 6) {real, imag} */,
  {32'h3f9cb64d, 32'h00000000} /* (24, 12, 5) {real, imag} */,
  {32'h3f4a2cf6, 32'h00000000} /* (24, 12, 4) {real, imag} */,
  {32'h3f6d21fe, 32'h00000000} /* (24, 12, 3) {real, imag} */,
  {32'h3f70ea23, 32'h00000000} /* (24, 12, 2) {real, imag} */,
  {32'h3f973101, 32'h00000000} /* (24, 12, 1) {real, imag} */,
  {32'h3f34d63f, 32'h00000000} /* (24, 12, 0) {real, imag} */,
  {32'h3eedb9c3, 32'h00000000} /* (24, 11, 31) {real, imag} */,
  {32'h3f82915a, 32'h00000000} /* (24, 11, 30) {real, imag} */,
  {32'h3ecd2087, 32'h00000000} /* (24, 11, 29) {real, imag} */,
  {32'h3f10a2f5, 32'h00000000} /* (24, 11, 28) {real, imag} */,
  {32'h3f48c20c, 32'h00000000} /* (24, 11, 27) {real, imag} */,
  {32'h3f98ac81, 32'h00000000} /* (24, 11, 26) {real, imag} */,
  {32'h3f9400cf, 32'h00000000} /* (24, 11, 25) {real, imag} */,
  {32'h3fb0e002, 32'h00000000} /* (24, 11, 24) {real, imag} */,
  {32'h3fa0dcc7, 32'h00000000} /* (24, 11, 23) {real, imag} */,
  {32'h3fa01c72, 32'h00000000} /* (24, 11, 22) {real, imag} */,
  {32'h3cc06698, 32'h00000000} /* (24, 11, 21) {real, imag} */,
  {32'hbf4364d5, 32'h00000000} /* (24, 11, 20) {real, imag} */,
  {32'hbf860f6c, 32'h00000000} /* (24, 11, 19) {real, imag} */,
  {32'hbf9306ef, 32'h00000000} /* (24, 11, 18) {real, imag} */,
  {32'hbf88b28b, 32'h00000000} /* (24, 11, 17) {real, imag} */,
  {32'hbefba2d4, 32'h00000000} /* (24, 11, 16) {real, imag} */,
  {32'hbf3836e3, 32'h00000000} /* (24, 11, 15) {real, imag} */,
  {32'hbe64a9b7, 32'h00000000} /* (24, 11, 14) {real, imag} */,
  {32'hbe8de10e, 32'h00000000} /* (24, 11, 13) {real, imag} */,
  {32'hbecc1b57, 32'h00000000} /* (24, 11, 12) {real, imag} */,
  {32'hbef0baa0, 32'h00000000} /* (24, 11, 11) {real, imag} */,
  {32'h3de32f80, 32'h00000000} /* (24, 11, 10) {real, imag} */,
  {32'h3f63636c, 32'h00000000} /* (24, 11, 9) {real, imag} */,
  {32'h3f8b4d83, 32'h00000000} /* (24, 11, 8) {real, imag} */,
  {32'h3fcd0bc5, 32'h00000000} /* (24, 11, 7) {real, imag} */,
  {32'h3fc0802f, 32'h00000000} /* (24, 11, 6) {real, imag} */,
  {32'h3f3ad90e, 32'h00000000} /* (24, 11, 5) {real, imag} */,
  {32'h3e447510, 32'h00000000} /* (24, 11, 4) {real, imag} */,
  {32'h3e7632c2, 32'h00000000} /* (24, 11, 3) {real, imag} */,
  {32'h3f55f14e, 32'h00000000} /* (24, 11, 2) {real, imag} */,
  {32'h3f3861a2, 32'h00000000} /* (24, 11, 1) {real, imag} */,
  {32'h3ed2ddb2, 32'h00000000} /* (24, 11, 0) {real, imag} */,
  {32'hbe37ee8d, 32'h00000000} /* (24, 10, 31) {real, imag} */,
  {32'hbf05ae29, 32'h00000000} /* (24, 10, 30) {real, imag} */,
  {32'hbef0b8b0, 32'h00000000} /* (24, 10, 29) {real, imag} */,
  {32'hbea5cbac, 32'h00000000} /* (24, 10, 28) {real, imag} */,
  {32'hbee5a470, 32'h00000000} /* (24, 10, 27) {real, imag} */,
  {32'hbe8287cb, 32'h00000000} /* (24, 10, 26) {real, imag} */,
  {32'hbd5b5be0, 32'h00000000} /* (24, 10, 25) {real, imag} */,
  {32'h3dcd4f8f, 32'h00000000} /* (24, 10, 24) {real, imag} */,
  {32'hbe41925d, 32'h00000000} /* (24, 10, 23) {real, imag} */,
  {32'hbe1dcd1e, 32'h00000000} /* (24, 10, 22) {real, imag} */,
  {32'hbf019656, 32'h00000000} /* (24, 10, 21) {real, imag} */,
  {32'h3d7c9898, 32'h00000000} /* (24, 10, 20) {real, imag} */,
  {32'h3ef52189, 32'h00000000} /* (24, 10, 19) {real, imag} */,
  {32'h3eb38471, 32'h00000000} /* (24, 10, 18) {real, imag} */,
  {32'h3f2d2461, 32'h00000000} /* (24, 10, 17) {real, imag} */,
  {32'h3f75de3e, 32'h00000000} /* (24, 10, 16) {real, imag} */,
  {32'h3f80e35a, 32'h00000000} /* (24, 10, 15) {real, imag} */,
  {32'h3f5cebd0, 32'h00000000} /* (24, 10, 14) {real, imag} */,
  {32'h3eff42b4, 32'h00000000} /* (24, 10, 13) {real, imag} */,
  {32'h3f103c90, 32'h00000000} /* (24, 10, 12) {real, imag} */,
  {32'h3e9be4b3, 32'h00000000} /* (24, 10, 11) {real, imag} */,
  {32'hbe546531, 32'h00000000} /* (24, 10, 10) {real, imag} */,
  {32'hbe40b835, 32'h00000000} /* (24, 10, 9) {real, imag} */,
  {32'hbec4cead, 32'h00000000} /* (24, 10, 8) {real, imag} */,
  {32'h3eb1f061, 32'h00000000} /* (24, 10, 7) {real, imag} */,
  {32'h3c0d4511, 32'h00000000} /* (24, 10, 6) {real, imag} */,
  {32'h3df5d049, 32'h00000000} /* (24, 10, 5) {real, imag} */,
  {32'hbf1c9ac1, 32'h00000000} /* (24, 10, 4) {real, imag} */,
  {32'hbfb88fd7, 32'h00000000} /* (24, 10, 3) {real, imag} */,
  {32'hbed772d4, 32'h00000000} /* (24, 10, 2) {real, imag} */,
  {32'hbf0f7a6e, 32'h00000000} /* (24, 10, 1) {real, imag} */,
  {32'hbeebc59b, 32'h00000000} /* (24, 10, 0) {real, imag} */,
  {32'hbf203ca5, 32'h00000000} /* (24, 9, 31) {real, imag} */,
  {32'hbf75c621, 32'h00000000} /* (24, 9, 30) {real, imag} */,
  {32'hbf803f09, 32'h00000000} /* (24, 9, 29) {real, imag} */,
  {32'hbf71a718, 32'h00000000} /* (24, 9, 28) {real, imag} */,
  {32'hbfad3ddd, 32'h00000000} /* (24, 9, 27) {real, imag} */,
  {32'hbfa53392, 32'h00000000} /* (24, 9, 26) {real, imag} */,
  {32'hbf619a12, 32'h00000000} /* (24, 9, 25) {real, imag} */,
  {32'hbf93b4b8, 32'h00000000} /* (24, 9, 24) {real, imag} */,
  {32'hbf5d0d69, 32'h00000000} /* (24, 9, 23) {real, imag} */,
  {32'hbef1d3be, 32'h00000000} /* (24, 9, 22) {real, imag} */,
  {32'hbeea4a8e, 32'h00000000} /* (24, 9, 21) {real, imag} */,
  {32'h3e887e6f, 32'h00000000} /* (24, 9, 20) {real, imag} */,
  {32'h3f48191c, 32'h00000000} /* (24, 9, 19) {real, imag} */,
  {32'h3f49db4f, 32'h00000000} /* (24, 9, 18) {real, imag} */,
  {32'h3f7adc8d, 32'h00000000} /* (24, 9, 17) {real, imag} */,
  {32'h3f9cc0fc, 32'h00000000} /* (24, 9, 16) {real, imag} */,
  {32'h3f976fec, 32'h00000000} /* (24, 9, 15) {real, imag} */,
  {32'h3facb1cc, 32'h00000000} /* (24, 9, 14) {real, imag} */,
  {32'h3f8459fd, 32'h00000000} /* (24, 9, 13) {real, imag} */,
  {32'h3f9100b4, 32'h00000000} /* (24, 9, 12) {real, imag} */,
  {32'h3f1b45de, 32'h00000000} /* (24, 9, 11) {real, imag} */,
  {32'hbe99ee2d, 32'h00000000} /* (24, 9, 10) {real, imag} */,
  {32'hbf224a41, 32'h00000000} /* (24, 9, 9) {real, imag} */,
  {32'hbf881307, 32'h00000000} /* (24, 9, 8) {real, imag} */,
  {32'hbf4bd00f, 32'h00000000} /* (24, 9, 7) {real, imag} */,
  {32'hbf73d97f, 32'h00000000} /* (24, 9, 6) {real, imag} */,
  {32'hbf0ce352, 32'h00000000} /* (24, 9, 5) {real, imag} */,
  {32'hbf089c4b, 32'h00000000} /* (24, 9, 4) {real, imag} */,
  {32'hbfb9117a, 32'h00000000} /* (24, 9, 3) {real, imag} */,
  {32'hbf9ab133, 32'h00000000} /* (24, 9, 2) {real, imag} */,
  {32'hbf856b8d, 32'h00000000} /* (24, 9, 1) {real, imag} */,
  {32'hbf03e023, 32'h00000000} /* (24, 9, 0) {real, imag} */,
  {32'hbec46a4e, 32'h00000000} /* (24, 8, 31) {real, imag} */,
  {32'hbeecab0f, 32'h00000000} /* (24, 8, 30) {real, imag} */,
  {32'hbf973c87, 32'h00000000} /* (24, 8, 29) {real, imag} */,
  {32'hbf940f61, 32'h00000000} /* (24, 8, 28) {real, imag} */,
  {32'hbf723abc, 32'h00000000} /* (24, 8, 27) {real, imag} */,
  {32'hbf77b9bb, 32'h00000000} /* (24, 8, 26) {real, imag} */,
  {32'hbf936e0e, 32'h00000000} /* (24, 8, 25) {real, imag} */,
  {32'hbf968228, 32'h00000000} /* (24, 8, 24) {real, imag} */,
  {32'hbf2f3432, 32'h00000000} /* (24, 8, 23) {real, imag} */,
  {32'hbf37b121, 32'h00000000} /* (24, 8, 22) {real, imag} */,
  {32'hbebfaadc, 32'h00000000} /* (24, 8, 21) {real, imag} */,
  {32'h3f0a1ea3, 32'h00000000} /* (24, 8, 20) {real, imag} */,
  {32'h3f09e57d, 32'h00000000} /* (24, 8, 19) {real, imag} */,
  {32'h3f0a719b, 32'h00000000} /* (24, 8, 18) {real, imag} */,
  {32'h3f459cf7, 32'h00000000} /* (24, 8, 17) {real, imag} */,
  {32'h3fa05242, 32'h00000000} /* (24, 8, 16) {real, imag} */,
  {32'h3f909062, 32'h00000000} /* (24, 8, 15) {real, imag} */,
  {32'h3f437506, 32'h00000000} /* (24, 8, 14) {real, imag} */,
  {32'h3fa79526, 32'h00000000} /* (24, 8, 13) {real, imag} */,
  {32'h3fd2d81c, 32'h00000000} /* (24, 8, 12) {real, imag} */,
  {32'h3f84cc19, 32'h00000000} /* (24, 8, 11) {real, imag} */,
  {32'h3de61ef1, 32'h00000000} /* (24, 8, 10) {real, imag} */,
  {32'hbe998649, 32'h00000000} /* (24, 8, 9) {real, imag} */,
  {32'hbf9f4ade, 32'h00000000} /* (24, 8, 8) {real, imag} */,
  {32'hbfe2b101, 32'h00000000} /* (24, 8, 7) {real, imag} */,
  {32'hbfc74306, 32'h00000000} /* (24, 8, 6) {real, imag} */,
  {32'hbf514837, 32'h00000000} /* (24, 8, 5) {real, imag} */,
  {32'hbeaae46d, 32'h00000000} /* (24, 8, 4) {real, imag} */,
  {32'hbf267435, 32'h00000000} /* (24, 8, 3) {real, imag} */,
  {32'hbf99fa9e, 32'h00000000} /* (24, 8, 2) {real, imag} */,
  {32'hbf9976a7, 32'h00000000} /* (24, 8, 1) {real, imag} */,
  {32'hbebdd88a, 32'h00000000} /* (24, 8, 0) {real, imag} */,
  {32'hbeac31dc, 32'h00000000} /* (24, 7, 31) {real, imag} */,
  {32'hbf325706, 32'h00000000} /* (24, 7, 30) {real, imag} */,
  {32'hbf786f04, 32'h00000000} /* (24, 7, 29) {real, imag} */,
  {32'hbf8cdc21, 32'h00000000} /* (24, 7, 28) {real, imag} */,
  {32'hbf60a2b0, 32'h00000000} /* (24, 7, 27) {real, imag} */,
  {32'hbf366216, 32'h00000000} /* (24, 7, 26) {real, imag} */,
  {32'hbf822650, 32'h00000000} /* (24, 7, 25) {real, imag} */,
  {32'hbfac1795, 32'h00000000} /* (24, 7, 24) {real, imag} */,
  {32'hbf9509a1, 32'h00000000} /* (24, 7, 23) {real, imag} */,
  {32'hbf6eeba8, 32'h00000000} /* (24, 7, 22) {real, imag} */,
  {32'hbda27b8a, 32'h00000000} /* (24, 7, 21) {real, imag} */,
  {32'h3fb308e6, 32'h00000000} /* (24, 7, 20) {real, imag} */,
  {32'h3f44b507, 32'h00000000} /* (24, 7, 19) {real, imag} */,
  {32'h3e96ced0, 32'h00000000} /* (24, 7, 18) {real, imag} */,
  {32'h3f41b9d4, 32'h00000000} /* (24, 7, 17) {real, imag} */,
  {32'h3f65639c, 32'h00000000} /* (24, 7, 16) {real, imag} */,
  {32'h3f075ed2, 32'h00000000} /* (24, 7, 15) {real, imag} */,
  {32'h3ee39c97, 32'h00000000} /* (24, 7, 14) {real, imag} */,
  {32'h3f6d07ef, 32'h00000000} /* (24, 7, 13) {real, imag} */,
  {32'h3f8d9732, 32'h00000000} /* (24, 7, 12) {real, imag} */,
  {32'h3f1f21d9, 32'h00000000} /* (24, 7, 11) {real, imag} */,
  {32'hbe58e38a, 32'h00000000} /* (24, 7, 10) {real, imag} */,
  {32'hbf67ae49, 32'h00000000} /* (24, 7, 9) {real, imag} */,
  {32'hbfa6d441, 32'h00000000} /* (24, 7, 8) {real, imag} */,
  {32'hbf6c4e77, 32'h00000000} /* (24, 7, 7) {real, imag} */,
  {32'hbf854526, 32'h00000000} /* (24, 7, 6) {real, imag} */,
  {32'hbf70f85a, 32'h00000000} /* (24, 7, 5) {real, imag} */,
  {32'hbf2512cc, 32'h00000000} /* (24, 7, 4) {real, imag} */,
  {32'hbf2d2181, 32'h00000000} /* (24, 7, 3) {real, imag} */,
  {32'hbf926e68, 32'h00000000} /* (24, 7, 2) {real, imag} */,
  {32'hbfa4a248, 32'h00000000} /* (24, 7, 1) {real, imag} */,
  {32'hbf0c5894, 32'h00000000} /* (24, 7, 0) {real, imag} */,
  {32'hbe673570, 32'h00000000} /* (24, 6, 31) {real, imag} */,
  {32'hbee507b2, 32'h00000000} /* (24, 6, 30) {real, imag} */,
  {32'hbf6faff6, 32'h00000000} /* (24, 6, 29) {real, imag} */,
  {32'hbf8d08f2, 32'h00000000} /* (24, 6, 28) {real, imag} */,
  {32'hbf18e0ce, 32'h00000000} /* (24, 6, 27) {real, imag} */,
  {32'hbf317778, 32'h00000000} /* (24, 6, 26) {real, imag} */,
  {32'hbf634ac7, 32'h00000000} /* (24, 6, 25) {real, imag} */,
  {32'hbf9dd1eb, 32'h00000000} /* (24, 6, 24) {real, imag} */,
  {32'hbfba1b57, 32'h00000000} /* (24, 6, 23) {real, imag} */,
  {32'hbf9e08ba, 32'h00000000} /* (24, 6, 22) {real, imag} */,
  {32'hbf3232da, 32'h00000000} /* (24, 6, 21) {real, imag} */,
  {32'h3f179787, 32'h00000000} /* (24, 6, 20) {real, imag} */,
  {32'h3f192e93, 32'h00000000} /* (24, 6, 19) {real, imag} */,
  {32'h3f3d69f2, 32'h00000000} /* (24, 6, 18) {real, imag} */,
  {32'h3f382a6a, 32'h00000000} /* (24, 6, 17) {real, imag} */,
  {32'h3f366306, 32'h00000000} /* (24, 6, 16) {real, imag} */,
  {32'h3f40f6dd, 32'h00000000} /* (24, 6, 15) {real, imag} */,
  {32'h3f7b1a25, 32'h00000000} /* (24, 6, 14) {real, imag} */,
  {32'h3f8c510e, 32'h00000000} /* (24, 6, 13) {real, imag} */,
  {32'h3f7d1a43, 32'h00000000} /* (24, 6, 12) {real, imag} */,
  {32'h3e9cf2ec, 32'h00000000} /* (24, 6, 11) {real, imag} */,
  {32'hbf03cd15, 32'h00000000} /* (24, 6, 10) {real, imag} */,
  {32'hbf694074, 32'h00000000} /* (24, 6, 9) {real, imag} */,
  {32'hbfa2de17, 32'h00000000} /* (24, 6, 8) {real, imag} */,
  {32'hbf8fe7b2, 32'h00000000} /* (24, 6, 7) {real, imag} */,
  {32'hbf761b76, 32'h00000000} /* (24, 6, 6) {real, imag} */,
  {32'hbf1487f0, 32'h00000000} /* (24, 6, 5) {real, imag} */,
  {32'hbee5b86b, 32'h00000000} /* (24, 6, 4) {real, imag} */,
  {32'hbf5160d2, 32'h00000000} /* (24, 6, 3) {real, imag} */,
  {32'hbf7ae873, 32'h00000000} /* (24, 6, 2) {real, imag} */,
  {32'hbfa090da, 32'h00000000} /* (24, 6, 1) {real, imag} */,
  {32'hbf363fba, 32'h00000000} /* (24, 6, 0) {real, imag} */,
  {32'hbf13dd2a, 32'h00000000} /* (24, 5, 31) {real, imag} */,
  {32'hbf6a79f0, 32'h00000000} /* (24, 5, 30) {real, imag} */,
  {32'hbf9ba96d, 32'h00000000} /* (24, 5, 29) {real, imag} */,
  {32'hbf978300, 32'h00000000} /* (24, 5, 28) {real, imag} */,
  {32'hbf37f628, 32'h00000000} /* (24, 5, 27) {real, imag} */,
  {32'hbf42585d, 32'h00000000} /* (24, 5, 26) {real, imag} */,
  {32'hbf70561e, 32'h00000000} /* (24, 5, 25) {real, imag} */,
  {32'hbf4eac52, 32'h00000000} /* (24, 5, 24) {real, imag} */,
  {32'hbf5569e7, 32'h00000000} /* (24, 5, 23) {real, imag} */,
  {32'hbf6bb055, 32'h00000000} /* (24, 5, 22) {real, imag} */,
  {32'hbf9bebb3, 32'h00000000} /* (24, 5, 21) {real, imag} */,
  {32'hbf1a917b, 32'h00000000} /* (24, 5, 20) {real, imag} */,
  {32'hbebae5d7, 32'h00000000} /* (24, 5, 19) {real, imag} */,
  {32'hbefdae6a, 32'h00000000} /* (24, 5, 18) {real, imag} */,
  {32'hbf0f7982, 32'h00000000} /* (24, 5, 17) {real, imag} */,
  {32'h3e8ca216, 32'h00000000} /* (24, 5, 16) {real, imag} */,
  {32'h3fa0aefa, 32'h00000000} /* (24, 5, 15) {real, imag} */,
  {32'h3f8298ab, 32'h00000000} /* (24, 5, 14) {real, imag} */,
  {32'h3f56063d, 32'h00000000} /* (24, 5, 13) {real, imag} */,
  {32'h3f4757b1, 32'h00000000} /* (24, 5, 12) {real, imag} */,
  {32'h3f1905e1, 32'h00000000} /* (24, 5, 11) {real, imag} */,
  {32'h3f093212, 32'h00000000} /* (24, 5, 10) {real, imag} */,
  {32'h3e12fe38, 32'h00000000} /* (24, 5, 9) {real, imag} */,
  {32'hbd012eb6, 32'h00000000} /* (24, 5, 8) {real, imag} */,
  {32'hbe3135ce, 32'h00000000} /* (24, 5, 7) {real, imag} */,
  {32'hbd545f4b, 32'h00000000} /* (24, 5, 6) {real, imag} */,
  {32'hbeddb5f3, 32'h00000000} /* (24, 5, 5) {real, imag} */,
  {32'hbee53074, 32'h00000000} /* (24, 5, 4) {real, imag} */,
  {32'hbf7c052b, 32'h00000000} /* (24, 5, 3) {real, imag} */,
  {32'hbf2543c3, 32'h00000000} /* (24, 5, 2) {real, imag} */,
  {32'hbf7a5163, 32'h00000000} /* (24, 5, 1) {real, imag} */,
  {32'hbf37720d, 32'h00000000} /* (24, 5, 0) {real, imag} */,
  {32'hbf11b77c, 32'h00000000} /* (24, 4, 31) {real, imag} */,
  {32'hbf907bd9, 32'h00000000} /* (24, 4, 30) {real, imag} */,
  {32'hbf7c3e9b, 32'h00000000} /* (24, 4, 29) {real, imag} */,
  {32'hbf6b477e, 32'h00000000} /* (24, 4, 28) {real, imag} */,
  {32'hbf480752, 32'h00000000} /* (24, 4, 27) {real, imag} */,
  {32'hbf4b9d6d, 32'h00000000} /* (24, 4, 26) {real, imag} */,
  {32'hbf62e9aa, 32'h00000000} /* (24, 4, 25) {real, imag} */,
  {32'hbf853108, 32'h00000000} /* (24, 4, 24) {real, imag} */,
  {32'hbf5b712a, 32'h00000000} /* (24, 4, 23) {real, imag} */,
  {32'hbf89043a, 32'h00000000} /* (24, 4, 22) {real, imag} */,
  {32'hbfae35d1, 32'h00000000} /* (24, 4, 21) {real, imag} */,
  {32'hbfb95cc4, 32'h00000000} /* (24, 4, 20) {real, imag} */,
  {32'hbf99002d, 32'h00000000} /* (24, 4, 19) {real, imag} */,
  {32'hbf99a74b, 32'h00000000} /* (24, 4, 18) {real, imag} */,
  {32'hbf9f16de, 32'h00000000} /* (24, 4, 17) {real, imag} */,
  {32'hbf1c7df3, 32'h00000000} /* (24, 4, 16) {real, imag} */,
  {32'h3f7a1222, 32'h00000000} /* (24, 4, 15) {real, imag} */,
  {32'h3f3dea1e, 32'h00000000} /* (24, 4, 14) {real, imag} */,
  {32'h3f1ca4c3, 32'h00000000} /* (24, 4, 13) {real, imag} */,
  {32'h3f2d482b, 32'h00000000} /* (24, 4, 12) {real, imag} */,
  {32'h3ec85e5c, 32'h00000000} /* (24, 4, 11) {real, imag} */,
  {32'h3f597eae, 32'h00000000} /* (24, 4, 10) {real, imag} */,
  {32'h3f718e75, 32'h00000000} /* (24, 4, 9) {real, imag} */,
  {32'h3f706fb7, 32'h00000000} /* (24, 4, 8) {real, imag} */,
  {32'h3f4d8cbc, 32'h00000000} /* (24, 4, 7) {real, imag} */,
  {32'h3f4b51d4, 32'h00000000} /* (24, 4, 6) {real, imag} */,
  {32'hbe7584e0, 32'h00000000} /* (24, 4, 5) {real, imag} */,
  {32'hbf392370, 32'h00000000} /* (24, 4, 4) {real, imag} */,
  {32'hbf491e9b, 32'h00000000} /* (24, 4, 3) {real, imag} */,
  {32'hbf37e457, 32'h00000000} /* (24, 4, 2) {real, imag} */,
  {32'hbf411318, 32'h00000000} /* (24, 4, 1) {real, imag} */,
  {32'hbec4c835, 32'h00000000} /* (24, 4, 0) {real, imag} */,
  {32'hbed39b21, 32'h00000000} /* (24, 3, 31) {real, imag} */,
  {32'hbf487968, 32'h00000000} /* (24, 3, 30) {real, imag} */,
  {32'hbf771dec, 32'h00000000} /* (24, 3, 29) {real, imag} */,
  {32'hbfabd81b, 32'h00000000} /* (24, 3, 28) {real, imag} */,
  {32'hbf952df7, 32'h00000000} /* (24, 3, 27) {real, imag} */,
  {32'hbf16922c, 32'h00000000} /* (24, 3, 26) {real, imag} */,
  {32'hbef5cf4b, 32'h00000000} /* (24, 3, 25) {real, imag} */,
  {32'hbf73082d, 32'h00000000} /* (24, 3, 24) {real, imag} */,
  {32'hbf33ede2, 32'h00000000} /* (24, 3, 23) {real, imag} */,
  {32'hbf852e89, 32'h00000000} /* (24, 3, 22) {real, imag} */,
  {32'hbf8d0916, 32'h00000000} /* (24, 3, 21) {real, imag} */,
  {32'hbf90865d, 32'h00000000} /* (24, 3, 20) {real, imag} */,
  {32'hbf6eb503, 32'h00000000} /* (24, 3, 19) {real, imag} */,
  {32'hbf645e7a, 32'h00000000} /* (24, 3, 18) {real, imag} */,
  {32'hbf7d2966, 32'h00000000} /* (24, 3, 17) {real, imag} */,
  {32'hbf5ba70c, 32'h00000000} /* (24, 3, 16) {real, imag} */,
  {32'h3f0dcad6, 32'h00000000} /* (24, 3, 15) {real, imag} */,
  {32'h3f8352af, 32'h00000000} /* (24, 3, 14) {real, imag} */,
  {32'h3fdc0dac, 32'h00000000} /* (24, 3, 13) {real, imag} */,
  {32'h3fbaa28e, 32'h00000000} /* (24, 3, 12) {real, imag} */,
  {32'h3f283277, 32'h00000000} /* (24, 3, 11) {real, imag} */,
  {32'h3f584048, 32'h00000000} /* (24, 3, 10) {real, imag} */,
  {32'h3f6aafca, 32'h00000000} /* (24, 3, 9) {real, imag} */,
  {32'h3f6ab8d2, 32'h00000000} /* (24, 3, 8) {real, imag} */,
  {32'h3f7ae071, 32'h00000000} /* (24, 3, 7) {real, imag} */,
  {32'h3f4b9f10, 32'h00000000} /* (24, 3, 6) {real, imag} */,
  {32'hbea1110d, 32'h00000000} /* (24, 3, 5) {real, imag} */,
  {32'hbf9a4ecf, 32'h00000000} /* (24, 3, 4) {real, imag} */,
  {32'hbf21ebe3, 32'h00000000} /* (24, 3, 3) {real, imag} */,
  {32'hbf6236e1, 32'h00000000} /* (24, 3, 2) {real, imag} */,
  {32'hbf788c67, 32'h00000000} /* (24, 3, 1) {real, imag} */,
  {32'hbf0bb019, 32'h00000000} /* (24, 3, 0) {real, imag} */,
  {32'hbe7238d5, 32'h00000000} /* (24, 2, 31) {real, imag} */,
  {32'hbf1fdf42, 32'h00000000} /* (24, 2, 30) {real, imag} */,
  {32'hbf3216ec, 32'h00000000} /* (24, 2, 29) {real, imag} */,
  {32'hbf779f4f, 32'h00000000} /* (24, 2, 28) {real, imag} */,
  {32'hbf9d9c04, 32'h00000000} /* (24, 2, 27) {real, imag} */,
  {32'hbf7268a2, 32'h00000000} /* (24, 2, 26) {real, imag} */,
  {32'hbf2c8b2d, 32'h00000000} /* (24, 2, 25) {real, imag} */,
  {32'hbf33ecd1, 32'h00000000} /* (24, 2, 24) {real, imag} */,
  {32'hbf186d28, 32'h00000000} /* (24, 2, 23) {real, imag} */,
  {32'hbf5592e0, 32'h00000000} /* (24, 2, 22) {real, imag} */,
  {32'hbf8eb910, 32'h00000000} /* (24, 2, 21) {real, imag} */,
  {32'hbf9454a0, 32'h00000000} /* (24, 2, 20) {real, imag} */,
  {32'hbfd54796, 32'h00000000} /* (24, 2, 19) {real, imag} */,
  {32'hbfc1ee84, 32'h00000000} /* (24, 2, 18) {real, imag} */,
  {32'hbf93fa76, 32'h00000000} /* (24, 2, 17) {real, imag} */,
  {32'hbf340886, 32'h00000000} /* (24, 2, 16) {real, imag} */,
  {32'h3ea50190, 32'h00000000} /* (24, 2, 15) {real, imag} */,
  {32'h3f2111d7, 32'h00000000} /* (24, 2, 14) {real, imag} */,
  {32'h3fb11405, 32'h00000000} /* (24, 2, 13) {real, imag} */,
  {32'h3fd9b153, 32'h00000000} /* (24, 2, 12) {real, imag} */,
  {32'h3f979d06, 32'h00000000} /* (24, 2, 11) {real, imag} */,
  {32'h3f97f469, 32'h00000000} /* (24, 2, 10) {real, imag} */,
  {32'h3f981090, 32'h00000000} /* (24, 2, 9) {real, imag} */,
  {32'h3f47ffd1, 32'h00000000} /* (24, 2, 8) {real, imag} */,
  {32'h3f7fd6df, 32'h00000000} /* (24, 2, 7) {real, imag} */,
  {32'h3f9cb4d3, 32'h00000000} /* (24, 2, 6) {real, imag} */,
  {32'h3e2041b8, 32'h00000000} /* (24, 2, 5) {real, imag} */,
  {32'hbf7471bc, 32'h00000000} /* (24, 2, 4) {real, imag} */,
  {32'hbf60b8fa, 32'h00000000} /* (24, 2, 3) {real, imag} */,
  {32'hbf5c714d, 32'h00000000} /* (24, 2, 2) {real, imag} */,
  {32'hbf201ff0, 32'h00000000} /* (24, 2, 1) {real, imag} */,
  {32'hbe9429d5, 32'h00000000} /* (24, 2, 0) {real, imag} */,
  {32'hbdd94367, 32'h00000000} /* (24, 1, 31) {real, imag} */,
  {32'hbee602a3, 32'h00000000} /* (24, 1, 30) {real, imag} */,
  {32'hbf455ba9, 32'h00000000} /* (24, 1, 29) {real, imag} */,
  {32'hbf7daec8, 32'h00000000} /* (24, 1, 28) {real, imag} */,
  {32'hbfb60d51, 32'h00000000} /* (24, 1, 27) {real, imag} */,
  {32'hbfa0c38f, 32'h00000000} /* (24, 1, 26) {real, imag} */,
  {32'hbf379be2, 32'h00000000} /* (24, 1, 25) {real, imag} */,
  {32'hbefadcde, 32'h00000000} /* (24, 1, 24) {real, imag} */,
  {32'hbf1b8fae, 32'h00000000} /* (24, 1, 23) {real, imag} */,
  {32'hbf184cb1, 32'h00000000} /* (24, 1, 22) {real, imag} */,
  {32'hbf75877c, 32'h00000000} /* (24, 1, 21) {real, imag} */,
  {32'hbf29c37c, 32'h00000000} /* (24, 1, 20) {real, imag} */,
  {32'hbfbfbfac, 32'h00000000} /* (24, 1, 19) {real, imag} */,
  {32'hbfaef4c3, 32'h00000000} /* (24, 1, 18) {real, imag} */,
  {32'hbf8eac24, 32'h00000000} /* (24, 1, 17) {real, imag} */,
  {32'hbeff8222, 32'h00000000} /* (24, 1, 16) {real, imag} */,
  {32'h3f0f947d, 32'h00000000} /* (24, 1, 15) {real, imag} */,
  {32'h3f473645, 32'h00000000} /* (24, 1, 14) {real, imag} */,
  {32'h3f2e9e9e, 32'h00000000} /* (24, 1, 13) {real, imag} */,
  {32'h3f7f0e88, 32'h00000000} /* (24, 1, 12) {real, imag} */,
  {32'h3fbf1a94, 32'h00000000} /* (24, 1, 11) {real, imag} */,
  {32'h3f8e3610, 32'h00000000} /* (24, 1, 10) {real, imag} */,
  {32'h3f90bbb5, 32'h00000000} /* (24, 1, 9) {real, imag} */,
  {32'h3fa1717e, 32'h00000000} /* (24, 1, 8) {real, imag} */,
  {32'h3f8588bd, 32'h00000000} /* (24, 1, 7) {real, imag} */,
  {32'h3f32acc5, 32'h00000000} /* (24, 1, 6) {real, imag} */,
  {32'hbe459d4d, 32'h00000000} /* (24, 1, 5) {real, imag} */,
  {32'hbf2cec4e, 32'h00000000} /* (24, 1, 4) {real, imag} */,
  {32'hbf5e0d80, 32'h00000000} /* (24, 1, 3) {real, imag} */,
  {32'hbf40e0ae, 32'h00000000} /* (24, 1, 2) {real, imag} */,
  {32'hbf04ff6f, 32'h00000000} /* (24, 1, 1) {real, imag} */,
  {32'hbe314ae4, 32'h00000000} /* (24, 1, 0) {real, imag} */,
  {32'hbe51e556, 32'h00000000} /* (24, 0, 31) {real, imag} */,
  {32'hbf08f82a, 32'h00000000} /* (24, 0, 30) {real, imag} */,
  {32'hbf50f4b4, 32'h00000000} /* (24, 0, 29) {real, imag} */,
  {32'hbf4a0f9b, 32'h00000000} /* (24, 0, 28) {real, imag} */,
  {32'hbf8d4172, 32'h00000000} /* (24, 0, 27) {real, imag} */,
  {32'hbf7f497d, 32'h00000000} /* (24, 0, 26) {real, imag} */,
  {32'hbead3eed, 32'h00000000} /* (24, 0, 25) {real, imag} */,
  {32'hbe6d1638, 32'h00000000} /* (24, 0, 24) {real, imag} */,
  {32'hbebfb91b, 32'h00000000} /* (24, 0, 23) {real, imag} */,
  {32'hbe659c44, 32'h00000000} /* (24, 0, 22) {real, imag} */,
  {32'hbe410139, 32'h00000000} /* (24, 0, 21) {real, imag} */,
  {32'hbe16c666, 32'h00000000} /* (24, 0, 20) {real, imag} */,
  {32'hbf064b4f, 32'h00000000} /* (24, 0, 19) {real, imag} */,
  {32'hbeb71e71, 32'h00000000} /* (24, 0, 18) {real, imag} */,
  {32'hbeadf9b8, 32'h00000000} /* (24, 0, 17) {real, imag} */,
  {32'hbde14615, 32'h00000000} /* (24, 0, 16) {real, imag} */,
  {32'h3e98493c, 32'h00000000} /* (24, 0, 15) {real, imag} */,
  {32'h3f13b46a, 32'h00000000} /* (24, 0, 14) {real, imag} */,
  {32'h3e92d9a5, 32'h00000000} /* (24, 0, 13) {real, imag} */,
  {32'h3e96b922, 32'h00000000} /* (24, 0, 12) {real, imag} */,
  {32'h3ef1d55e, 32'h00000000} /* (24, 0, 11) {real, imag} */,
  {32'h3e5b5d86, 32'h00000000} /* (24, 0, 10) {real, imag} */,
  {32'h3eb85cac, 32'h00000000} /* (24, 0, 9) {real, imag} */,
  {32'h3f5b8735, 32'h00000000} /* (24, 0, 8) {real, imag} */,
  {32'h3f0d65d6, 32'h00000000} /* (24, 0, 7) {real, imag} */,
  {32'h3e2dea14, 32'h00000000} /* (24, 0, 6) {real, imag} */,
  {32'hbe80c2c4, 32'h00000000} /* (24, 0, 5) {real, imag} */,
  {32'hbedbe4d5, 32'h00000000} /* (24, 0, 4) {real, imag} */,
  {32'hbf0870c8, 32'h00000000} /* (24, 0, 3) {real, imag} */,
  {32'hbf1c8320, 32'h00000000} /* (24, 0, 2) {real, imag} */,
  {32'hbef367f6, 32'h00000000} /* (24, 0, 1) {real, imag} */,
  {32'hbe45cbd5, 32'h00000000} /* (24, 0, 0) {real, imag} */,
  {32'hbeb33d1f, 32'h00000000} /* (23, 31, 31) {real, imag} */,
  {32'hbf552e08, 32'h00000000} /* (23, 31, 30) {real, imag} */,
  {32'hbf22b9bb, 32'h00000000} /* (23, 31, 29) {real, imag} */,
  {32'hbebb715c, 32'h00000000} /* (23, 31, 28) {real, imag} */,
  {32'hbf07f4d1, 32'h00000000} /* (23, 31, 27) {real, imag} */,
  {32'hbf5155d7, 32'h00000000} /* (23, 31, 26) {real, imag} */,
  {32'hbf080054, 32'h00000000} /* (23, 31, 25) {real, imag} */,
  {32'hbf128ae8, 32'h00000000} /* (23, 31, 24) {real, imag} */,
  {32'hbedcfc09, 32'h00000000} /* (23, 31, 23) {real, imag} */,
  {32'hbf33998d, 32'h00000000} /* (23, 31, 22) {real, imag} */,
  {32'hbde5167a, 32'h00000000} /* (23, 31, 21) {real, imag} */,
  {32'h3f3bc656, 32'h00000000} /* (23, 31, 20) {real, imag} */,
  {32'h3e855376, 32'h00000000} /* (23, 31, 19) {real, imag} */,
  {32'h3e8e446b, 32'h00000000} /* (23, 31, 18) {real, imag} */,
  {32'h3eeb57cd, 32'h00000000} /* (23, 31, 17) {real, imag} */,
  {32'h3f150531, 32'h00000000} /* (23, 31, 16) {real, imag} */,
  {32'h3f0ef95a, 32'h00000000} /* (23, 31, 15) {real, imag} */,
  {32'h3eede70a, 32'h00000000} /* (23, 31, 14) {real, imag} */,
  {32'h3edf4729, 32'h00000000} /* (23, 31, 13) {real, imag} */,
  {32'h3ef7e07c, 32'h00000000} /* (23, 31, 12) {real, imag} */,
  {32'h3ecc8287, 32'h00000000} /* (23, 31, 11) {real, imag} */,
  {32'hbe9a34ad, 32'h00000000} /* (23, 31, 10) {real, imag} */,
  {32'hbf1d7781, 32'h00000000} /* (23, 31, 9) {real, imag} */,
  {32'hbf1a08b1, 32'h00000000} /* (23, 31, 8) {real, imag} */,
  {32'hbb111fe6, 32'h00000000} /* (23, 31, 7) {real, imag} */,
  {32'hbe994b57, 32'h00000000} /* (23, 31, 6) {real, imag} */,
  {32'hbf005be6, 32'h00000000} /* (23, 31, 5) {real, imag} */,
  {32'hbed8f597, 32'h00000000} /* (23, 31, 4) {real, imag} */,
  {32'hbea3246e, 32'h00000000} /* (23, 31, 3) {real, imag} */,
  {32'hbe0a8c50, 32'h00000000} /* (23, 31, 2) {real, imag} */,
  {32'hbe7b2cf2, 32'h00000000} /* (23, 31, 1) {real, imag} */,
  {32'hbe3fd5fc, 32'h00000000} /* (23, 31, 0) {real, imag} */,
  {32'hbe9fc230, 32'h00000000} /* (23, 30, 31) {real, imag} */,
  {32'hbf6fa71b, 32'h00000000} /* (23, 30, 30) {real, imag} */,
  {32'hbf755f0e, 32'h00000000} /* (23, 30, 29) {real, imag} */,
  {32'hbf33f65a, 32'h00000000} /* (23, 30, 28) {real, imag} */,
  {32'hbf455de6, 32'h00000000} /* (23, 30, 27) {real, imag} */,
  {32'hbf4f840f, 32'h00000000} /* (23, 30, 26) {real, imag} */,
  {32'hbf879fbc, 32'h00000000} /* (23, 30, 25) {real, imag} */,
  {32'hbfbcdd8d, 32'h00000000} /* (23, 30, 24) {real, imag} */,
  {32'hbf8792fb, 32'h00000000} /* (23, 30, 23) {real, imag} */,
  {32'hbf815649, 32'h00000000} /* (23, 30, 22) {real, imag} */,
  {32'hbf0dea87, 32'h00000000} /* (23, 30, 21) {real, imag} */,
  {32'h3f702c45, 32'h00000000} /* (23, 30, 20) {real, imag} */,
  {32'h3ee69ff4, 32'h00000000} /* (23, 30, 19) {real, imag} */,
  {32'h3f319fb5, 32'h00000000} /* (23, 30, 18) {real, imag} */,
  {32'h3f650f79, 32'h00000000} /* (23, 30, 17) {real, imag} */,
  {32'h3f9144e0, 32'h00000000} /* (23, 30, 16) {real, imag} */,
  {32'h3f14407e, 32'h00000000} /* (23, 30, 15) {real, imag} */,
  {32'h3ef53d0d, 32'h00000000} /* (23, 30, 14) {real, imag} */,
  {32'h3f0d2511, 32'h00000000} /* (23, 30, 13) {real, imag} */,
  {32'h3f87eb5c, 32'h00000000} /* (23, 30, 12) {real, imag} */,
  {32'h3fa452a1, 32'h00000000} /* (23, 30, 11) {real, imag} */,
  {32'hbe419deb, 32'h00000000} /* (23, 30, 10) {real, imag} */,
  {32'hbf8ede92, 32'h00000000} /* (23, 30, 9) {real, imag} */,
  {32'hbf8805d2, 32'h00000000} /* (23, 30, 8) {real, imag} */,
  {32'hbe6f7c89, 32'h00000000} /* (23, 30, 7) {real, imag} */,
  {32'hbee14417, 32'h00000000} /* (23, 30, 6) {real, imag} */,
  {32'hbf411bd4, 32'h00000000} /* (23, 30, 5) {real, imag} */,
  {32'hbf3e3646, 32'h00000000} /* (23, 30, 4) {real, imag} */,
  {32'hbf47a041, 32'h00000000} /* (23, 30, 3) {real, imag} */,
  {32'hbed3fe5d, 32'h00000000} /* (23, 30, 2) {real, imag} */,
  {32'hbeb91927, 32'h00000000} /* (23, 30, 1) {real, imag} */,
  {32'hbe8c69c9, 32'h00000000} /* (23, 30, 0) {real, imag} */,
  {32'hbeea0c38, 32'h00000000} /* (23, 29, 31) {real, imag} */,
  {32'hbf6268a5, 32'h00000000} /* (23, 29, 30) {real, imag} */,
  {32'hbf3e851c, 32'h00000000} /* (23, 29, 29) {real, imag} */,
  {32'hbf42af72, 32'h00000000} /* (23, 29, 28) {real, imag} */,
  {32'hbf4ce3c3, 32'h00000000} /* (23, 29, 27) {real, imag} */,
  {32'hbf4c9ce8, 32'h00000000} /* (23, 29, 26) {real, imag} */,
  {32'hbfc6a21b, 32'h00000000} /* (23, 29, 25) {real, imag} */,
  {32'hbfab80ef, 32'h00000000} /* (23, 29, 24) {real, imag} */,
  {32'hbf62c782, 32'h00000000} /* (23, 29, 23) {real, imag} */,
  {32'hbf227d2a, 32'h00000000} /* (23, 29, 22) {real, imag} */,
  {32'hbf3065ad, 32'h00000000} /* (23, 29, 21) {real, imag} */,
  {32'h3e955c75, 32'h00000000} /* (23, 29, 20) {real, imag} */,
  {32'h3f5e65a7, 32'h00000000} /* (23, 29, 19) {real, imag} */,
  {32'h3f8fd1ed, 32'h00000000} /* (23, 29, 18) {real, imag} */,
  {32'h3f95fa48, 32'h00000000} /* (23, 29, 17) {real, imag} */,
  {32'h3f8a9678, 32'h00000000} /* (23, 29, 16) {real, imag} */,
  {32'h3f3a27ee, 32'h00000000} /* (23, 29, 15) {real, imag} */,
  {32'h3efb4bd5, 32'h00000000} /* (23, 29, 14) {real, imag} */,
  {32'h3ed678e8, 32'h00000000} /* (23, 29, 13) {real, imag} */,
  {32'h3f6cbde5, 32'h00000000} /* (23, 29, 12) {real, imag} */,
  {32'h3f67997e, 32'h00000000} /* (23, 29, 11) {real, imag} */,
  {32'h3e3dab5e, 32'h00000000} /* (23, 29, 10) {real, imag} */,
  {32'hbf36f532, 32'h00000000} /* (23, 29, 9) {real, imag} */,
  {32'hbf9765c5, 32'h00000000} /* (23, 29, 8) {real, imag} */,
  {32'hbf77087f, 32'h00000000} /* (23, 29, 7) {real, imag} */,
  {32'hbf098b01, 32'h00000000} /* (23, 29, 6) {real, imag} */,
  {32'hbf031e52, 32'h00000000} /* (23, 29, 5) {real, imag} */,
  {32'hbe810ceb, 32'h00000000} /* (23, 29, 4) {real, imag} */,
  {32'hbeb0d39a, 32'h00000000} /* (23, 29, 3) {real, imag} */,
  {32'hbf5b49ea, 32'h00000000} /* (23, 29, 2) {real, imag} */,
  {32'hbf6d491b, 32'h00000000} /* (23, 29, 1) {real, imag} */,
  {32'hbebc87c0, 32'h00000000} /* (23, 29, 0) {real, imag} */,
  {32'hbf6f03cc, 32'h00000000} /* (23, 28, 31) {real, imag} */,
  {32'hbf946226, 32'h00000000} /* (23, 28, 30) {real, imag} */,
  {32'hbf5ee2b4, 32'h00000000} /* (23, 28, 29) {real, imag} */,
  {32'hbf1a68e9, 32'h00000000} /* (23, 28, 28) {real, imag} */,
  {32'hbf378751, 32'h00000000} /* (23, 28, 27) {real, imag} */,
  {32'hbf3134c3, 32'h00000000} /* (23, 28, 26) {real, imag} */,
  {32'hbfa23cb6, 32'h00000000} /* (23, 28, 25) {real, imag} */,
  {32'hbf9153cb, 32'h00000000} /* (23, 28, 24) {real, imag} */,
  {32'hbf40c63a, 32'h00000000} /* (23, 28, 23) {real, imag} */,
  {32'hbf3f0375, 32'h00000000} /* (23, 28, 22) {real, imag} */,
  {32'hbf187530, 32'h00000000} /* (23, 28, 21) {real, imag} */,
  {32'h3ee596f5, 32'h00000000} /* (23, 28, 20) {real, imag} */,
  {32'h3f8a84db, 32'h00000000} /* (23, 28, 19) {real, imag} */,
  {32'h3f88e40d, 32'h00000000} /* (23, 28, 18) {real, imag} */,
  {32'h3f71e9cd, 32'h00000000} /* (23, 28, 17) {real, imag} */,
  {32'h3fa91cbc, 32'h00000000} /* (23, 28, 16) {real, imag} */,
  {32'h3fba6aba, 32'h00000000} /* (23, 28, 15) {real, imag} */,
  {32'h3f6aa67b, 32'h00000000} /* (23, 28, 14) {real, imag} */,
  {32'h3f136b8f, 32'h00000000} /* (23, 28, 13) {real, imag} */,
  {32'h3f60bbc2, 32'h00000000} /* (23, 28, 12) {real, imag} */,
  {32'h3f532e6d, 32'h00000000} /* (23, 28, 11) {real, imag} */,
  {32'hbdab8e8e, 32'h00000000} /* (23, 28, 10) {real, imag} */,
  {32'hbf4d6787, 32'h00000000} /* (23, 28, 9) {real, imag} */,
  {32'hbfb2c5aa, 32'h00000000} /* (23, 28, 8) {real, imag} */,
  {32'hbfa35ff4, 32'h00000000} /* (23, 28, 7) {real, imag} */,
  {32'hbf6021c3, 32'h00000000} /* (23, 28, 6) {real, imag} */,
  {32'hbf2d13d1, 32'h00000000} /* (23, 28, 5) {real, imag} */,
  {32'hbf14c37e, 32'h00000000} /* (23, 28, 4) {real, imag} */,
  {32'hbf86bfda, 32'h00000000} /* (23, 28, 3) {real, imag} */,
  {32'hbfa3d32d, 32'h00000000} /* (23, 28, 2) {real, imag} */,
  {32'hbf51ceea, 32'h00000000} /* (23, 28, 1) {real, imag} */,
  {32'hbea4d86e, 32'h00000000} /* (23, 28, 0) {real, imag} */,
  {32'hbf0296ee, 32'h00000000} /* (23, 27, 31) {real, imag} */,
  {32'hbf970b38, 32'h00000000} /* (23, 27, 30) {real, imag} */,
  {32'hbf53c32b, 32'h00000000} /* (23, 27, 29) {real, imag} */,
  {32'hbf5521b9, 32'h00000000} /* (23, 27, 28) {real, imag} */,
  {32'hbfb79273, 32'h00000000} /* (23, 27, 27) {real, imag} */,
  {32'hbfb21631, 32'h00000000} /* (23, 27, 26) {real, imag} */,
  {32'hbf80de00, 32'h00000000} /* (23, 27, 25) {real, imag} */,
  {32'hbf4e9a01, 32'h00000000} /* (23, 27, 24) {real, imag} */,
  {32'hbf06796b, 32'h00000000} /* (23, 27, 23) {real, imag} */,
  {32'hbed737dd, 32'h00000000} /* (23, 27, 22) {real, imag} */,
  {32'hbe9208f3, 32'h00000000} /* (23, 27, 21) {real, imag} */,
  {32'h3e643ef2, 32'h00000000} /* (23, 27, 20) {real, imag} */,
  {32'h3f4d226b, 32'h00000000} /* (23, 27, 19) {real, imag} */,
  {32'h3f9b6b7a, 32'h00000000} /* (23, 27, 18) {real, imag} */,
  {32'h3f71a7bb, 32'h00000000} /* (23, 27, 17) {real, imag} */,
  {32'h3f4755d6, 32'h00000000} /* (23, 27, 16) {real, imag} */,
  {32'h3f3b49b6, 32'h00000000} /* (23, 27, 15) {real, imag} */,
  {32'h3f20dc3e, 32'h00000000} /* (23, 27, 14) {real, imag} */,
  {32'h3f5b49fa, 32'h00000000} /* (23, 27, 13) {real, imag} */,
  {32'h3f5e5e85, 32'h00000000} /* (23, 27, 12) {real, imag} */,
  {32'h3f6de2c3, 32'h00000000} /* (23, 27, 11) {real, imag} */,
  {32'hbe9cca87, 32'h00000000} /* (23, 27, 10) {real, imag} */,
  {32'hbf8a0366, 32'h00000000} /* (23, 27, 9) {real, imag} */,
  {32'hbf746463, 32'h00000000} /* (23, 27, 8) {real, imag} */,
  {32'hbf5bda25, 32'h00000000} /* (23, 27, 7) {real, imag} */,
  {32'hbf51b7b5, 32'h00000000} /* (23, 27, 6) {real, imag} */,
  {32'hbf83863c, 32'h00000000} /* (23, 27, 5) {real, imag} */,
  {32'hbfa3febc, 32'h00000000} /* (23, 27, 4) {real, imag} */,
  {32'hbfd57284, 32'h00000000} /* (23, 27, 3) {real, imag} */,
  {32'hbf9a47fc, 32'h00000000} /* (23, 27, 2) {real, imag} */,
  {32'hbead0bbe, 32'h00000000} /* (23, 27, 1) {real, imag} */,
  {32'hbe63fea5, 32'h00000000} /* (23, 27, 0) {real, imag} */,
  {32'hbebb4a23, 32'h00000000} /* (23, 26, 31) {real, imag} */,
  {32'hbf5b0670, 32'h00000000} /* (23, 26, 30) {real, imag} */,
  {32'hbf773a64, 32'h00000000} /* (23, 26, 29) {real, imag} */,
  {32'hbf903c43, 32'h00000000} /* (23, 26, 28) {real, imag} */,
  {32'hbfcb2db9, 32'h00000000} /* (23, 26, 27) {real, imag} */,
  {32'hbff34359, 32'h00000000} /* (23, 26, 26) {real, imag} */,
  {32'hbf95eb2e, 32'h00000000} /* (23, 26, 25) {real, imag} */,
  {32'hbf659192, 32'h00000000} /* (23, 26, 24) {real, imag} */,
  {32'hbf889c92, 32'h00000000} /* (23, 26, 23) {real, imag} */,
  {32'hbf571735, 32'h00000000} /* (23, 26, 22) {real, imag} */,
  {32'hbe199d06, 32'h00000000} /* (23, 26, 21) {real, imag} */,
  {32'h3eb28bf4, 32'h00000000} /* (23, 26, 20) {real, imag} */,
  {32'h3f4352c7, 32'h00000000} /* (23, 26, 19) {real, imag} */,
  {32'h3f8c7b12, 32'h00000000} /* (23, 26, 18) {real, imag} */,
  {32'h3f77e33a, 32'h00000000} /* (23, 26, 17) {real, imag} */,
  {32'h3ec3dca7, 32'h00000000} /* (23, 26, 16) {real, imag} */,
  {32'h3f19c25b, 32'h00000000} /* (23, 26, 15) {real, imag} */,
  {32'h3f2ddcb2, 32'h00000000} /* (23, 26, 14) {real, imag} */,
  {32'h3f14d86a, 32'h00000000} /* (23, 26, 13) {real, imag} */,
  {32'h3f1a371d, 32'h00000000} /* (23, 26, 12) {real, imag} */,
  {32'h3f0d6754, 32'h00000000} /* (23, 26, 11) {real, imag} */,
  {32'hbeed8ea3, 32'h00000000} /* (23, 26, 10) {real, imag} */,
  {32'hbf6ce518, 32'h00000000} /* (23, 26, 9) {real, imag} */,
  {32'hbefd740f, 32'h00000000} /* (23, 26, 8) {real, imag} */,
  {32'hbf2b3619, 32'h00000000} /* (23, 26, 7) {real, imag} */,
  {32'hbf297195, 32'h00000000} /* (23, 26, 6) {real, imag} */,
  {32'hbebcba65, 32'h00000000} /* (23, 26, 5) {real, imag} */,
  {32'hbf4e6e98, 32'h00000000} /* (23, 26, 4) {real, imag} */,
  {32'hbf7972f0, 32'h00000000} /* (23, 26, 3) {real, imag} */,
  {32'hbf6531c3, 32'h00000000} /* (23, 26, 2) {real, imag} */,
  {32'hbee7a80f, 32'h00000000} /* (23, 26, 1) {real, imag} */,
  {32'hbe95d60f, 32'h00000000} /* (23, 26, 0) {real, imag} */,
  {32'hbf15615c, 32'h00000000} /* (23, 25, 31) {real, imag} */,
  {32'hbfafa8ca, 32'h00000000} /* (23, 25, 30) {real, imag} */,
  {32'hbfad41a2, 32'h00000000} /* (23, 25, 29) {real, imag} */,
  {32'hbf7fb6f0, 32'h00000000} /* (23, 25, 28) {real, imag} */,
  {32'hbf7f1ecf, 32'h00000000} /* (23, 25, 27) {real, imag} */,
  {32'hbf89b2be, 32'h00000000} /* (23, 25, 26) {real, imag} */,
  {32'hbf9d1e05, 32'h00000000} /* (23, 25, 25) {real, imag} */,
  {32'hbf8c8b73, 32'h00000000} /* (23, 25, 24) {real, imag} */,
  {32'hbf8bd133, 32'h00000000} /* (23, 25, 23) {real, imag} */,
  {32'hbf594154, 32'h00000000} /* (23, 25, 22) {real, imag} */,
  {32'hbe9ba98e, 32'h00000000} /* (23, 25, 21) {real, imag} */,
  {32'h3f357502, 32'h00000000} /* (23, 25, 20) {real, imag} */,
  {32'h3f7bb1b5, 32'h00000000} /* (23, 25, 19) {real, imag} */,
  {32'h3f76cf21, 32'h00000000} /* (23, 25, 18) {real, imag} */,
  {32'h3f869851, 32'h00000000} /* (23, 25, 17) {real, imag} */,
  {32'h3f39f402, 32'h00000000} /* (23, 25, 16) {real, imag} */,
  {32'h3f478ffb, 32'h00000000} /* (23, 25, 15) {real, imag} */,
  {32'h3fa8262b, 32'h00000000} /* (23, 25, 14) {real, imag} */,
  {32'h3f8be880, 32'h00000000} /* (23, 25, 13) {real, imag} */,
  {32'h3f249417, 32'h00000000} /* (23, 25, 12) {real, imag} */,
  {32'h3dfca044, 32'h00000000} /* (23, 25, 11) {real, imag} */,
  {32'hbf98de6f, 32'h00000000} /* (23, 25, 10) {real, imag} */,
  {32'hbf92e402, 32'h00000000} /* (23, 25, 9) {real, imag} */,
  {32'hbf3d02d7, 32'h00000000} /* (23, 25, 8) {real, imag} */,
  {32'hbf4d53fd, 32'h00000000} /* (23, 25, 7) {real, imag} */,
  {32'hbf5559da, 32'h00000000} /* (23, 25, 6) {real, imag} */,
  {32'hbf1b212c, 32'h00000000} /* (23, 25, 5) {real, imag} */,
  {32'hbf7a0ea2, 32'h00000000} /* (23, 25, 4) {real, imag} */,
  {32'hbf96faf3, 32'h00000000} /* (23, 25, 3) {real, imag} */,
  {32'hbf8b4caf, 32'h00000000} /* (23, 25, 2) {real, imag} */,
  {32'hbec806aa, 32'h00000000} /* (23, 25, 1) {real, imag} */,
  {32'hbd0f5b81, 32'h00000000} /* (23, 25, 0) {real, imag} */,
  {32'hbee38085, 32'h00000000} /* (23, 24, 31) {real, imag} */,
  {32'hbf7a79ea, 32'h00000000} /* (23, 24, 30) {real, imag} */,
  {32'hbf86caf5, 32'h00000000} /* (23, 24, 29) {real, imag} */,
  {32'hbf9d5a0f, 32'h00000000} /* (23, 24, 28) {real, imag} */,
  {32'hbfa8e204, 32'h00000000} /* (23, 24, 27) {real, imag} */,
  {32'hbf158bf1, 32'h00000000} /* (23, 24, 26) {real, imag} */,
  {32'hbf42a166, 32'h00000000} /* (23, 24, 25) {real, imag} */,
  {32'hbf1997ae, 32'h00000000} /* (23, 24, 24) {real, imag} */,
  {32'hbf6106a5, 32'h00000000} /* (23, 24, 23) {real, imag} */,
  {32'hbf8785e6, 32'h00000000} /* (23, 24, 22) {real, imag} */,
  {32'hbf168f32, 32'h00000000} /* (23, 24, 21) {real, imag} */,
  {32'h3eb088b9, 32'h00000000} /* (23, 24, 20) {real, imag} */,
  {32'h3f24ebf0, 32'h00000000} /* (23, 24, 19) {real, imag} */,
  {32'h3f728766, 32'h00000000} /* (23, 24, 18) {real, imag} */,
  {32'h3fbd8850, 32'h00000000} /* (23, 24, 17) {real, imag} */,
  {32'h3fa605f5, 32'h00000000} /* (23, 24, 16) {real, imag} */,
  {32'h3f85050c, 32'h00000000} /* (23, 24, 15) {real, imag} */,
  {32'h3fd5fb30, 32'h00000000} /* (23, 24, 14) {real, imag} */,
  {32'h3f758889, 32'h00000000} /* (23, 24, 13) {real, imag} */,
  {32'h3f0dc013, 32'h00000000} /* (23, 24, 12) {real, imag} */,
  {32'h3dc04ea5, 32'h00000000} /* (23, 24, 11) {real, imag} */,
  {32'hbf42555c, 32'h00000000} /* (23, 24, 10) {real, imag} */,
  {32'hbf5eb05b, 32'h00000000} /* (23, 24, 9) {real, imag} */,
  {32'hbf9c1105, 32'h00000000} /* (23, 24, 8) {real, imag} */,
  {32'hbfb0c302, 32'h00000000} /* (23, 24, 7) {real, imag} */,
  {32'hbf60f514, 32'h00000000} /* (23, 24, 6) {real, imag} */,
  {32'hbf11af6b, 32'h00000000} /* (23, 24, 5) {real, imag} */,
  {32'hbf1fcb4b, 32'h00000000} /* (23, 24, 4) {real, imag} */,
  {32'hbfa0d5f8, 32'h00000000} /* (23, 24, 3) {real, imag} */,
  {32'hbf803859, 32'h00000000} /* (23, 24, 2) {real, imag} */,
  {32'hbea87c84, 32'h00000000} /* (23, 24, 1) {real, imag} */,
  {32'hbdd2ccf0, 32'h00000000} /* (23, 24, 0) {real, imag} */,
  {32'hbf2745a9, 32'h00000000} /* (23, 23, 31) {real, imag} */,
  {32'hbf45aaaa, 32'h00000000} /* (23, 23, 30) {real, imag} */,
  {32'hbf3ef453, 32'h00000000} /* (23, 23, 29) {real, imag} */,
  {32'hbf95141b, 32'h00000000} /* (23, 23, 28) {real, imag} */,
  {32'hbfaa13fe, 32'h00000000} /* (23, 23, 27) {real, imag} */,
  {32'hbf5c922d, 32'h00000000} /* (23, 23, 26) {real, imag} */,
  {32'hbf71e386, 32'h00000000} /* (23, 23, 25) {real, imag} */,
  {32'hbf2f2eef, 32'h00000000} /* (23, 23, 24) {real, imag} */,
  {32'hbf8b356b, 32'h00000000} /* (23, 23, 23) {real, imag} */,
  {32'hbf86aae0, 32'h00000000} /* (23, 23, 22) {real, imag} */,
  {32'hbeb8ea55, 32'h00000000} /* (23, 23, 21) {real, imag} */,
  {32'h3f14c129, 32'h00000000} /* (23, 23, 20) {real, imag} */,
  {32'h3f8b2453, 32'h00000000} /* (23, 23, 19) {real, imag} */,
  {32'h3fa640ae, 32'h00000000} /* (23, 23, 18) {real, imag} */,
  {32'h3fcfb6e8, 32'h00000000} /* (23, 23, 17) {real, imag} */,
  {32'h3f9152f8, 32'h00000000} /* (23, 23, 16) {real, imag} */,
  {32'h3f8024d7, 32'h00000000} /* (23, 23, 15) {real, imag} */,
  {32'h3fb95ee2, 32'h00000000} /* (23, 23, 14) {real, imag} */,
  {32'h3f4c0f1a, 32'h00000000} /* (23, 23, 13) {real, imag} */,
  {32'h3f52b543, 32'h00000000} /* (23, 23, 12) {real, imag} */,
  {32'h3eb34bf8, 32'h00000000} /* (23, 23, 11) {real, imag} */,
  {32'hbebc4200, 32'h00000000} /* (23, 23, 10) {real, imag} */,
  {32'hbeee649b, 32'h00000000} /* (23, 23, 9) {real, imag} */,
  {32'hbf807f1f, 32'h00000000} /* (23, 23, 8) {real, imag} */,
  {32'hbfa6c3ce, 32'h00000000} /* (23, 23, 7) {real, imag} */,
  {32'hbf48def4, 32'h00000000} /* (23, 23, 6) {real, imag} */,
  {32'hbf517d2b, 32'h00000000} /* (23, 23, 5) {real, imag} */,
  {32'hbf65343d, 32'h00000000} /* (23, 23, 4) {real, imag} */,
  {32'hbf4cdce7, 32'h00000000} /* (23, 23, 3) {real, imag} */,
  {32'hbec5a49f, 32'h00000000} /* (23, 23, 2) {real, imag} */,
  {32'hbee0c0cd, 32'h00000000} /* (23, 23, 1) {real, imag} */,
  {32'hbf1b4ef6, 32'h00000000} /* (23, 23, 0) {real, imag} */,
  {32'hbf0e5a1f, 32'h00000000} /* (23, 22, 31) {real, imag} */,
  {32'hbf333d4b, 32'h00000000} /* (23, 22, 30) {real, imag} */,
  {32'hbf6dc393, 32'h00000000} /* (23, 22, 29) {real, imag} */,
  {32'hbf72b53e, 32'h00000000} /* (23, 22, 28) {real, imag} */,
  {32'hbf2e76d8, 32'h00000000} /* (23, 22, 27) {real, imag} */,
  {32'hbefa2e5f, 32'h00000000} /* (23, 22, 26) {real, imag} */,
  {32'hbf2dea60, 32'h00000000} /* (23, 22, 25) {real, imag} */,
  {32'hbf4d3c2c, 32'h00000000} /* (23, 22, 24) {real, imag} */,
  {32'hbf65f797, 32'h00000000} /* (23, 22, 23) {real, imag} */,
  {32'hbf8b56ed, 32'h00000000} /* (23, 22, 22) {real, imag} */,
  {32'hbec3c71f, 32'h00000000} /* (23, 22, 21) {real, imag} */,
  {32'h3f68b116, 32'h00000000} /* (23, 22, 20) {real, imag} */,
  {32'h3fd4a7d3, 32'h00000000} /* (23, 22, 19) {real, imag} */,
  {32'h3fd635f4, 32'h00000000} /* (23, 22, 18) {real, imag} */,
  {32'h3f980c13, 32'h00000000} /* (23, 22, 17) {real, imag} */,
  {32'h3f91b89b, 32'h00000000} /* (23, 22, 16) {real, imag} */,
  {32'h3f394033, 32'h00000000} /* (23, 22, 15) {real, imag} */,
  {32'h3f672049, 32'h00000000} /* (23, 22, 14) {real, imag} */,
  {32'h3f5afb5b, 32'h00000000} /* (23, 22, 13) {real, imag} */,
  {32'h3f75528f, 32'h00000000} /* (23, 22, 12) {real, imag} */,
  {32'h3f1bc278, 32'h00000000} /* (23, 22, 11) {real, imag} */,
  {32'hbe826c5a, 32'h00000000} /* (23, 22, 10) {real, imag} */,
  {32'hbf1d7566, 32'h00000000} /* (23, 22, 9) {real, imag} */,
  {32'hbf4edf16, 32'h00000000} /* (23, 22, 8) {real, imag} */,
  {32'hbf4fce97, 32'h00000000} /* (23, 22, 7) {real, imag} */,
  {32'hbf2b679e, 32'h00000000} /* (23, 22, 6) {real, imag} */,
  {32'hbf454c9a, 32'h00000000} /* (23, 22, 5) {real, imag} */,
  {32'hbf58884b, 32'h00000000} /* (23, 22, 4) {real, imag} */,
  {32'hbf338e50, 32'h00000000} /* (23, 22, 3) {real, imag} */,
  {32'hbe75478e, 32'h00000000} /* (23, 22, 2) {real, imag} */,
  {32'hbf149bff, 32'h00000000} /* (23, 22, 1) {real, imag} */,
  {32'hbf37d90d, 32'h00000000} /* (23, 22, 0) {real, imag} */,
  {32'hbda52b67, 32'h00000000} /* (23, 21, 31) {real, imag} */,
  {32'hbeb2b57c, 32'h00000000} /* (23, 21, 30) {real, imag} */,
  {32'hbf8066ca, 32'h00000000} /* (23, 21, 29) {real, imag} */,
  {32'hbf68e7ce, 32'h00000000} /* (23, 21, 28) {real, imag} */,
  {32'hbe1cd3f4, 32'h00000000} /* (23, 21, 27) {real, imag} */,
  {32'h3ececd77, 32'h00000000} /* (23, 21, 26) {real, imag} */,
  {32'hbe3a24a8, 32'h00000000} /* (23, 21, 25) {real, imag} */,
  {32'hbea5761d, 32'h00000000} /* (23, 21, 24) {real, imag} */,
  {32'hbda5a9e0, 32'h00000000} /* (23, 21, 23) {real, imag} */,
  {32'hbf282320, 32'h00000000} /* (23, 21, 22) {real, imag} */,
  {32'hbf2e15af, 32'h00000000} /* (23, 21, 21) {real, imag} */,
  {32'hbe1bd488, 32'h00000000} /* (23, 21, 20) {real, imag} */,
  {32'h3ee1b2c1, 32'h00000000} /* (23, 21, 19) {real, imag} */,
  {32'h3f984d81, 32'h00000000} /* (23, 21, 18) {real, imag} */,
  {32'h3f352991, 32'h00000000} /* (23, 21, 17) {real, imag} */,
  {32'h3ea7bf71, 32'h00000000} /* (23, 21, 16) {real, imag} */,
  {32'h3e44ba32, 32'h00000000} /* (23, 21, 15) {real, imag} */,
  {32'h3f7eb8b9, 32'h00000000} /* (23, 21, 14) {real, imag} */,
  {32'h3f65564e, 32'h00000000} /* (23, 21, 13) {real, imag} */,
  {32'h3f12fe05, 32'h00000000} /* (23, 21, 12) {real, imag} */,
  {32'h3d289eff, 32'h00000000} /* (23, 21, 11) {real, imag} */,
  {32'hbea02f43, 32'h00000000} /* (23, 21, 10) {real, imag} */,
  {32'h3e4a0b8b, 32'h00000000} /* (23, 21, 9) {real, imag} */,
  {32'hbed19b38, 32'h00000000} /* (23, 21, 8) {real, imag} */,
  {32'hbf15049b, 32'h00000000} /* (23, 21, 7) {real, imag} */,
  {32'hbef53d23, 32'h00000000} /* (23, 21, 6) {real, imag} */,
  {32'hbf1e11c0, 32'h00000000} /* (23, 21, 5) {real, imag} */,
  {32'hbf47dea3, 32'h00000000} /* (23, 21, 4) {real, imag} */,
  {32'hbf01249e, 32'h00000000} /* (23, 21, 3) {real, imag} */,
  {32'hbe9899aa, 32'h00000000} /* (23, 21, 2) {real, imag} */,
  {32'hbec674fb, 32'h00000000} /* (23, 21, 1) {real, imag} */,
  {32'hbee5fbf6, 32'h00000000} /* (23, 21, 0) {real, imag} */,
  {32'h3f52c970, 32'h00000000} /* (23, 20, 31) {real, imag} */,
  {32'h3fafafec, 32'h00000000} /* (23, 20, 30) {real, imag} */,
  {32'h3f2e0c84, 32'h00000000} /* (23, 20, 29) {real, imag} */,
  {32'h3ebda233, 32'h00000000} /* (23, 20, 28) {real, imag} */,
  {32'h3f528da3, 32'h00000000} /* (23, 20, 27) {real, imag} */,
  {32'h3fc10053, 32'h00000000} /* (23, 20, 26) {real, imag} */,
  {32'h3fa2208b, 32'h00000000} /* (23, 20, 25) {real, imag} */,
  {32'h3f8e859d, 32'h00000000} /* (23, 20, 24) {real, imag} */,
  {32'h3fa5c62c, 32'h00000000} /* (23, 20, 23) {real, imag} */,
  {32'h3f1cd2ca, 32'h00000000} /* (23, 20, 22) {real, imag} */,
  {32'h3e0d2a93, 32'h00000000} /* (23, 20, 21) {real, imag} */,
  {32'hbf6f0c4e, 32'h00000000} /* (23, 20, 20) {real, imag} */,
  {32'hbf98868f, 32'h00000000} /* (23, 20, 19) {real, imag} */,
  {32'hbed6bf1b, 32'h00000000} /* (23, 20, 18) {real, imag} */,
  {32'hbf85560a, 32'h00000000} /* (23, 20, 17) {real, imag} */,
  {32'hbf9ffb44, 32'h00000000} /* (23, 20, 16) {real, imag} */,
  {32'hbe67f070, 32'h00000000} /* (23, 20, 15) {real, imag} */,
  {32'h3eaead69, 32'h00000000} /* (23, 20, 14) {real, imag} */,
  {32'hbe239082, 32'h00000000} /* (23, 20, 13) {real, imag} */,
  {32'hbe6c6048, 32'h00000000} /* (23, 20, 12) {real, imag} */,
  {32'hbef4815e, 32'h00000000} /* (23, 20, 11) {real, imag} */,
  {32'h3dacced7, 32'h00000000} /* (23, 20, 10) {real, imag} */,
  {32'h3f98de38, 32'h00000000} /* (23, 20, 9) {real, imag} */,
  {32'h3f3bb887, 32'h00000000} /* (23, 20, 8) {real, imag} */,
  {32'h3f05f65d, 32'h00000000} /* (23, 20, 7) {real, imag} */,
  {32'h3f3d81d4, 32'h00000000} /* (23, 20, 6) {real, imag} */,
  {32'h3f0b7c68, 32'h00000000} /* (23, 20, 5) {real, imag} */,
  {32'h3f133790, 32'h00000000} /* (23, 20, 4) {real, imag} */,
  {32'h3f2fd975, 32'h00000000} /* (23, 20, 3) {real, imag} */,
  {32'h3e955ab9, 32'h00000000} /* (23, 20, 2) {real, imag} */,
  {32'h3efe8976, 32'h00000000} /* (23, 20, 1) {real, imag} */,
  {32'h3e7b7d19, 32'h00000000} /* (23, 20, 0) {real, imag} */,
  {32'h3f6eb113, 32'h00000000} /* (23, 19, 31) {real, imag} */,
  {32'h3fb37c1b, 32'h00000000} /* (23, 19, 30) {real, imag} */,
  {32'h3f507505, 32'h00000000} /* (23, 19, 29) {real, imag} */,
  {32'h3f191d41, 32'h00000000} /* (23, 19, 28) {real, imag} */,
  {32'h3f4e7c01, 32'h00000000} /* (23, 19, 27) {real, imag} */,
  {32'h3f416b7d, 32'h00000000} /* (23, 19, 26) {real, imag} */,
  {32'h3f4558a8, 32'h00000000} /* (23, 19, 25) {real, imag} */,
  {32'h3f796675, 32'h00000000} /* (23, 19, 24) {real, imag} */,
  {32'h3fb6015a, 32'h00000000} /* (23, 19, 23) {real, imag} */,
  {32'h3fa60428, 32'h00000000} /* (23, 19, 22) {real, imag} */,
  {32'h3f0ce8b6, 32'h00000000} /* (23, 19, 21) {real, imag} */,
  {32'hbf0a090d, 32'h00000000} /* (23, 19, 20) {real, imag} */,
  {32'hbf70338c, 32'h00000000} /* (23, 19, 19) {real, imag} */,
  {32'hbf562dc5, 32'h00000000} /* (23, 19, 18) {real, imag} */,
  {32'hbf334058, 32'h00000000} /* (23, 19, 17) {real, imag} */,
  {32'hbf4e6130, 32'h00000000} /* (23, 19, 16) {real, imag} */,
  {32'hbe637d90, 32'h00000000} /* (23, 19, 15) {real, imag} */,
  {32'hbed13dfd, 32'h00000000} /* (23, 19, 14) {real, imag} */,
  {32'hbf66778e, 32'h00000000} /* (23, 19, 13) {real, imag} */,
  {32'hbf530402, 32'h00000000} /* (23, 19, 12) {real, imag} */,
  {32'hbf621837, 32'h00000000} /* (23, 19, 11) {real, imag} */,
  {32'hbe4c5825, 32'h00000000} /* (23, 19, 10) {real, imag} */,
  {32'h3f297a98, 32'h00000000} /* (23, 19, 9) {real, imag} */,
  {32'h3f175d18, 32'h00000000} /* (23, 19, 8) {real, imag} */,
  {32'h3f5426e5, 32'h00000000} /* (23, 19, 7) {real, imag} */,
  {32'h3f97d96e, 32'h00000000} /* (23, 19, 6) {real, imag} */,
  {32'h3faffa85, 32'h00000000} /* (23, 19, 5) {real, imag} */,
  {32'h3fa6b4ac, 32'h00000000} /* (23, 19, 4) {real, imag} */,
  {32'h3f3afb1d, 32'h00000000} /* (23, 19, 3) {real, imag} */,
  {32'h3f34f3c2, 32'h00000000} /* (23, 19, 2) {real, imag} */,
  {32'h3f7e895a, 32'h00000000} /* (23, 19, 1) {real, imag} */,
  {32'h3f082d64, 32'h00000000} /* (23, 19, 0) {real, imag} */,
  {32'h3f315915, 32'h00000000} /* (23, 18, 31) {real, imag} */,
  {32'h3faa3c51, 32'h00000000} /* (23, 18, 30) {real, imag} */,
  {32'h3f9d0352, 32'h00000000} /* (23, 18, 29) {real, imag} */,
  {32'h3f3fec98, 32'h00000000} /* (23, 18, 28) {real, imag} */,
  {32'h3ea2dc0b, 32'h00000000} /* (23, 18, 27) {real, imag} */,
  {32'h3d29b2b5, 32'h00000000} /* (23, 18, 26) {real, imag} */,
  {32'h3f08059a, 32'h00000000} /* (23, 18, 25) {real, imag} */,
  {32'h3f5177c1, 32'h00000000} /* (23, 18, 24) {real, imag} */,
  {32'h3f68fc0a, 32'h00000000} /* (23, 18, 23) {real, imag} */,
  {32'h3f69e92a, 32'h00000000} /* (23, 18, 22) {real, imag} */,
  {32'h3f2f6b63, 32'h00000000} /* (23, 18, 21) {real, imag} */,
  {32'hbf4c76ed, 32'h00000000} /* (23, 18, 20) {real, imag} */,
  {32'hbfc4fcf8, 32'h00000000} /* (23, 18, 19) {real, imag} */,
  {32'hbfa31122, 32'h00000000} /* (23, 18, 18) {real, imag} */,
  {32'hbee78d8c, 32'h00000000} /* (23, 18, 17) {real, imag} */,
  {32'hbe6d1768, 32'h00000000} /* (23, 18, 16) {real, imag} */,
  {32'hbf11d2bc, 32'h00000000} /* (23, 18, 15) {real, imag} */,
  {32'hbf8fac81, 32'h00000000} /* (23, 18, 14) {real, imag} */,
  {32'hbf8646e4, 32'h00000000} /* (23, 18, 13) {real, imag} */,
  {32'hbf6dd087, 32'h00000000} /* (23, 18, 12) {real, imag} */,
  {32'hbf6c6cbb, 32'h00000000} /* (23, 18, 11) {real, imag} */,
  {32'h3e796855, 32'h00000000} /* (23, 18, 10) {real, imag} */,
  {32'h3f560fbe, 32'h00000000} /* (23, 18, 9) {real, imag} */,
  {32'h3f7d4a38, 32'h00000000} /* (23, 18, 8) {real, imag} */,
  {32'h3f8bcf78, 32'h00000000} /* (23, 18, 7) {real, imag} */,
  {32'h3f81ed80, 32'h00000000} /* (23, 18, 6) {real, imag} */,
  {32'h3f894186, 32'h00000000} /* (23, 18, 5) {real, imag} */,
  {32'h3f681f69, 32'h00000000} /* (23, 18, 4) {real, imag} */,
  {32'h3f0eac6a, 32'h00000000} /* (23, 18, 3) {real, imag} */,
  {32'h3f4c994a, 32'h00000000} /* (23, 18, 2) {real, imag} */,
  {32'h3fb0d3c2, 32'h00000000} /* (23, 18, 1) {real, imag} */,
  {32'h3f3208d9, 32'h00000000} /* (23, 18, 0) {real, imag} */,
  {32'h3f81f391, 32'h00000000} /* (23, 17, 31) {real, imag} */,
  {32'h3f8686a8, 32'h00000000} /* (23, 17, 30) {real, imag} */,
  {32'h3f6fa6d0, 32'h00000000} /* (23, 17, 29) {real, imag} */,
  {32'h3f693960, 32'h00000000} /* (23, 17, 28) {real, imag} */,
  {32'h3deda694, 32'h00000000} /* (23, 17, 27) {real, imag} */,
  {32'hbdeab030, 32'h00000000} /* (23, 17, 26) {real, imag} */,
  {32'h3f36ca86, 32'h00000000} /* (23, 17, 25) {real, imag} */,
  {32'h3f7d5d11, 32'h00000000} /* (23, 17, 24) {real, imag} */,
  {32'h3f88f8ba, 32'h00000000} /* (23, 17, 23) {real, imag} */,
  {32'h3f483da7, 32'h00000000} /* (23, 17, 22) {real, imag} */,
  {32'h3e9e7e8d, 32'h00000000} /* (23, 17, 21) {real, imag} */,
  {32'hbf79c2d6, 32'h00000000} /* (23, 17, 20) {real, imag} */,
  {32'hbf9ca187, 32'h00000000} /* (23, 17, 19) {real, imag} */,
  {32'hbfa4d072, 32'h00000000} /* (23, 17, 18) {real, imag} */,
  {32'hbf73b180, 32'h00000000} /* (23, 17, 17) {real, imag} */,
  {32'hbf2fcace, 32'h00000000} /* (23, 17, 16) {real, imag} */,
  {32'hbf89cf34, 32'h00000000} /* (23, 17, 15) {real, imag} */,
  {32'hbfa3a085, 32'h00000000} /* (23, 17, 14) {real, imag} */,
  {32'hbf7dde9f, 32'h00000000} /* (23, 17, 13) {real, imag} */,
  {32'hbfa94e24, 32'h00000000} /* (23, 17, 12) {real, imag} */,
  {32'hbfabea2b, 32'h00000000} /* (23, 17, 11) {real, imag} */,
  {32'hbea28f1e, 32'h00000000} /* (23, 17, 10) {real, imag} */,
  {32'h3f82244d, 32'h00000000} /* (23, 17, 9) {real, imag} */,
  {32'h3f894427, 32'h00000000} /* (23, 17, 8) {real, imag} */,
  {32'h3f50bf10, 32'h00000000} /* (23, 17, 7) {real, imag} */,
  {32'h3f40133a, 32'h00000000} /* (23, 17, 6) {real, imag} */,
  {32'h3f2ce002, 32'h00000000} /* (23, 17, 5) {real, imag} */,
  {32'h3f1a7b1d, 32'h00000000} /* (23, 17, 4) {real, imag} */,
  {32'h3f096eae, 32'h00000000} /* (23, 17, 3) {real, imag} */,
  {32'h3f498293, 32'h00000000} /* (23, 17, 2) {real, imag} */,
  {32'h3f9c5571, 32'h00000000} /* (23, 17, 1) {real, imag} */,
  {32'h3f6ef2ec, 32'h00000000} /* (23, 17, 0) {real, imag} */,
  {32'h3f2c4105, 32'h00000000} /* (23, 16, 31) {real, imag} */,
  {32'h3f8d5cef, 32'h00000000} /* (23, 16, 30) {real, imag} */,
  {32'h3f87f7f1, 32'h00000000} /* (23, 16, 29) {real, imag} */,
  {32'h3eeeb433, 32'h00000000} /* (23, 16, 28) {real, imag} */,
  {32'h3f028605, 32'h00000000} /* (23, 16, 27) {real, imag} */,
  {32'h3f04c4a0, 32'h00000000} /* (23, 16, 26) {real, imag} */,
  {32'h3f831935, 32'h00000000} /* (23, 16, 25) {real, imag} */,
  {32'h3f904470, 32'h00000000} /* (23, 16, 24) {real, imag} */,
  {32'h3fc27ccc, 32'h00000000} /* (23, 16, 23) {real, imag} */,
  {32'h3f9ce170, 32'h00000000} /* (23, 16, 22) {real, imag} */,
  {32'h3d3bbd53, 32'h00000000} /* (23, 16, 21) {real, imag} */,
  {32'hbf8c350c, 32'h00000000} /* (23, 16, 20) {real, imag} */,
  {32'hbf5a50f4, 32'h00000000} /* (23, 16, 19) {real, imag} */,
  {32'hbf79d666, 32'h00000000} /* (23, 16, 18) {real, imag} */,
  {32'hbf69d479, 32'h00000000} /* (23, 16, 17) {real, imag} */,
  {32'hbf792f05, 32'h00000000} /* (23, 16, 16) {real, imag} */,
  {32'hbf414b41, 32'h00000000} /* (23, 16, 15) {real, imag} */,
  {32'hbf2e98f7, 32'h00000000} /* (23, 16, 14) {real, imag} */,
  {32'hbf65db43, 32'h00000000} /* (23, 16, 13) {real, imag} */,
  {32'hbfabba87, 32'h00000000} /* (23, 16, 12) {real, imag} */,
  {32'hbf7f9ba8, 32'h00000000} /* (23, 16, 11) {real, imag} */,
  {32'hbdcce2c9, 32'h00000000} /* (23, 16, 10) {real, imag} */,
  {32'h3f9b52e7, 32'h00000000} /* (23, 16, 9) {real, imag} */,
  {32'h3f44f5d3, 32'h00000000} /* (23, 16, 8) {real, imag} */,
  {32'h3f02f6b5, 32'h00000000} /* (23, 16, 7) {real, imag} */,
  {32'h3eca5165, 32'h00000000} /* (23, 16, 6) {real, imag} */,
  {32'h3f3e763c, 32'h00000000} /* (23, 16, 5) {real, imag} */,
  {32'h3f73a8b9, 32'h00000000} /* (23, 16, 4) {real, imag} */,
  {32'h3f4277f8, 32'h00000000} /* (23, 16, 3) {real, imag} */,
  {32'h3f92dd6e, 32'h00000000} /* (23, 16, 2) {real, imag} */,
  {32'h3f911655, 32'h00000000} /* (23, 16, 1) {real, imag} */,
  {32'h3f0efacc, 32'h00000000} /* (23, 16, 0) {real, imag} */,
  {32'h3efb3ab5, 32'h00000000} /* (23, 15, 31) {real, imag} */,
  {32'h3f7b2d8d, 32'h00000000} /* (23, 15, 30) {real, imag} */,
  {32'h3f8e7efe, 32'h00000000} /* (23, 15, 29) {real, imag} */,
  {32'h3f3d222e, 32'h00000000} /* (23, 15, 28) {real, imag} */,
  {32'h3fa54464, 32'h00000000} /* (23, 15, 27) {real, imag} */,
  {32'h3f9e0e3d, 32'h00000000} /* (23, 15, 26) {real, imag} */,
  {32'h3f30ae86, 32'h00000000} /* (23, 15, 25) {real, imag} */,
  {32'h3f590190, 32'h00000000} /* (23, 15, 24) {real, imag} */,
  {32'h3f96aa52, 32'h00000000} /* (23, 15, 23) {real, imag} */,
  {32'h3f1c3c2b, 32'h00000000} /* (23, 15, 22) {real, imag} */,
  {32'hbebf60e3, 32'h00000000} /* (23, 15, 21) {real, imag} */,
  {32'hbfac1661, 32'h00000000} /* (23, 15, 20) {real, imag} */,
  {32'hbf55d3e8, 32'h00000000} /* (23, 15, 19) {real, imag} */,
  {32'hbf653b72, 32'h00000000} /* (23, 15, 18) {real, imag} */,
  {32'hbf63d012, 32'h00000000} /* (23, 15, 17) {real, imag} */,
  {32'hbf5ed2cf, 32'h00000000} /* (23, 15, 16) {real, imag} */,
  {32'hbec8a174, 32'h00000000} /* (23, 15, 15) {real, imag} */,
  {32'hbec5dc3e, 32'h00000000} /* (23, 15, 14) {real, imag} */,
  {32'hbf886dfc, 32'h00000000} /* (23, 15, 13) {real, imag} */,
  {32'hbfafaf5e, 32'h00000000} /* (23, 15, 12) {real, imag} */,
  {32'hbf2d9c76, 32'h00000000} /* (23, 15, 11) {real, imag} */,
  {32'h3dca5ba7, 32'h00000000} /* (23, 15, 10) {real, imag} */,
  {32'h3f31f559, 32'h00000000} /* (23, 15, 9) {real, imag} */,
  {32'h3f54de25, 32'h00000000} /* (23, 15, 8) {real, imag} */,
  {32'h3f3c0951, 32'h00000000} /* (23, 15, 7) {real, imag} */,
  {32'h3f0cb706, 32'h00000000} /* (23, 15, 6) {real, imag} */,
  {32'h3f3a1ab6, 32'h00000000} /* (23, 15, 5) {real, imag} */,
  {32'h3f87e59b, 32'h00000000} /* (23, 15, 4) {real, imag} */,
  {32'h3f9d6054, 32'h00000000} /* (23, 15, 3) {real, imag} */,
  {32'h3f869df3, 32'h00000000} /* (23, 15, 2) {real, imag} */,
  {32'h3f43b50b, 32'h00000000} /* (23, 15, 1) {real, imag} */,
  {32'h3f09f03b, 32'h00000000} /* (23, 15, 0) {real, imag} */,
  {32'h3f27d8f8, 32'h00000000} /* (23, 14, 31) {real, imag} */,
  {32'h3f5db3ba, 32'h00000000} /* (23, 14, 30) {real, imag} */,
  {32'h3f5dd21b, 32'h00000000} /* (23, 14, 29) {real, imag} */,
  {32'h3f5248f7, 32'h00000000} /* (23, 14, 28) {real, imag} */,
  {32'h3f49e80a, 32'h00000000} /* (23, 14, 27) {real, imag} */,
  {32'h3f366404, 32'h00000000} /* (23, 14, 26) {real, imag} */,
  {32'h3f1f26b6, 32'h00000000} /* (23, 14, 25) {real, imag} */,
  {32'h3fbf8b22, 32'h00000000} /* (23, 14, 24) {real, imag} */,
  {32'h3fe2b3e7, 32'h00000000} /* (23, 14, 23) {real, imag} */,
  {32'h3f6e9ed5, 32'h00000000} /* (23, 14, 22) {real, imag} */,
  {32'hbd958fe7, 32'h00000000} /* (23, 14, 21) {real, imag} */,
  {32'hbf62447b, 32'h00000000} /* (23, 14, 20) {real, imag} */,
  {32'hbf629124, 32'h00000000} /* (23, 14, 19) {real, imag} */,
  {32'hbf38db39, 32'h00000000} /* (23, 14, 18) {real, imag} */,
  {32'hbf4a3402, 32'h00000000} /* (23, 14, 17) {real, imag} */,
  {32'hbf0bbbdb, 32'h00000000} /* (23, 14, 16) {real, imag} */,
  {32'hbe955671, 32'h00000000} /* (23, 14, 15) {real, imag} */,
  {32'hbec980c0, 32'h00000000} /* (23, 14, 14) {real, imag} */,
  {32'hbf33ba20, 32'h00000000} /* (23, 14, 13) {real, imag} */,
  {32'hbf60fa68, 32'h00000000} /* (23, 14, 12) {real, imag} */,
  {32'hbf1511e1, 32'h00000000} /* (23, 14, 11) {real, imag} */,
  {32'h3ef5145f, 32'h00000000} /* (23, 14, 10) {real, imag} */,
  {32'h3f8da9e0, 32'h00000000} /* (23, 14, 9) {real, imag} */,
  {32'h3fc5e34d, 32'h00000000} /* (23, 14, 8) {real, imag} */,
  {32'h3faa046e, 32'h00000000} /* (23, 14, 7) {real, imag} */,
  {32'h3f37dd1c, 32'h00000000} /* (23, 14, 6) {real, imag} */,
  {32'h3f5e2d71, 32'h00000000} /* (23, 14, 5) {real, imag} */,
  {32'h3f97f6c6, 32'h00000000} /* (23, 14, 4) {real, imag} */,
  {32'h3f81e090, 32'h00000000} /* (23, 14, 3) {real, imag} */,
  {32'h3eb6f680, 32'h00000000} /* (23, 14, 2) {real, imag} */,
  {32'h3f21eb4c, 32'h00000000} /* (23, 14, 1) {real, imag} */,
  {32'h3f718bf3, 32'h00000000} /* (23, 14, 0) {real, imag} */,
  {32'h3f0b3ae9, 32'h00000000} /* (23, 13, 31) {real, imag} */,
  {32'h3f0ed898, 32'h00000000} /* (23, 13, 30) {real, imag} */,
  {32'h3f7ea014, 32'h00000000} /* (23, 13, 29) {real, imag} */,
  {32'h3f9558bd, 32'h00000000} /* (23, 13, 28) {real, imag} */,
  {32'h3f62ae48, 32'h00000000} /* (23, 13, 27) {real, imag} */,
  {32'h3f1595a6, 32'h00000000} /* (23, 13, 26) {real, imag} */,
  {32'h3ec591bc, 32'h00000000} /* (23, 13, 25) {real, imag} */,
  {32'h3f9370c5, 32'h00000000} /* (23, 13, 24) {real, imag} */,
  {32'h3fd7b90a, 32'h00000000} /* (23, 13, 23) {real, imag} */,
  {32'h3fb52d7f, 32'h00000000} /* (23, 13, 22) {real, imag} */,
  {32'h3f0f79f1, 32'h00000000} /* (23, 13, 21) {real, imag} */,
  {32'hbf35d21a, 32'h00000000} /* (23, 13, 20) {real, imag} */,
  {32'hbfa0c06a, 32'h00000000} /* (23, 13, 19) {real, imag} */,
  {32'hbf764a3c, 32'h00000000} /* (23, 13, 18) {real, imag} */,
  {32'hbf835906, 32'h00000000} /* (23, 13, 17) {real, imag} */,
  {32'hbef38538, 32'h00000000} /* (23, 13, 16) {real, imag} */,
  {32'hbe02ab77, 32'h00000000} /* (23, 13, 15) {real, imag} */,
  {32'hbe6a036e, 32'h00000000} /* (23, 13, 14) {real, imag} */,
  {32'hbf80b0e8, 32'h00000000} /* (23, 13, 13) {real, imag} */,
  {32'hbf9144e7, 32'h00000000} /* (23, 13, 12) {real, imag} */,
  {32'hbf3e9408, 32'h00000000} /* (23, 13, 11) {real, imag} */,
  {32'h3f108289, 32'h00000000} /* (23, 13, 10) {real, imag} */,
  {32'h3facff19, 32'h00000000} /* (23, 13, 9) {real, imag} */,
  {32'h3fa723aa, 32'h00000000} /* (23, 13, 8) {real, imag} */,
  {32'h3fa4451f, 32'h00000000} /* (23, 13, 7) {real, imag} */,
  {32'h3f8edd46, 32'h00000000} /* (23, 13, 6) {real, imag} */,
  {32'h3f8fe6bf, 32'h00000000} /* (23, 13, 5) {real, imag} */,
  {32'h3f6bfb15, 32'h00000000} /* (23, 13, 4) {real, imag} */,
  {32'h3f04761d, 32'h00000000} /* (23, 13, 3) {real, imag} */,
  {32'hbdb56202, 32'h00000000} /* (23, 13, 2) {real, imag} */,
  {32'h3f0f06d8, 32'h00000000} /* (23, 13, 1) {real, imag} */,
  {32'h3f43cda9, 32'h00000000} /* (23, 13, 0) {real, imag} */,
  {32'h3f29695a, 32'h00000000} /* (23, 12, 31) {real, imag} */,
  {32'h3f46ebb0, 32'h00000000} /* (23, 12, 30) {real, imag} */,
  {32'h3f641c8b, 32'h00000000} /* (23, 12, 29) {real, imag} */,
  {32'h3faec288, 32'h00000000} /* (23, 12, 28) {real, imag} */,
  {32'h3f8f7f68, 32'h00000000} /* (23, 12, 27) {real, imag} */,
  {32'h3f91f1b0, 32'h00000000} /* (23, 12, 26) {real, imag} */,
  {32'h3f03e1ec, 32'h00000000} /* (23, 12, 25) {real, imag} */,
  {32'h3f2c3b0c, 32'h00000000} /* (23, 12, 24) {real, imag} */,
  {32'h3f8fa3e7, 32'h00000000} /* (23, 12, 23) {real, imag} */,
  {32'h3faec01a, 32'h00000000} /* (23, 12, 22) {real, imag} */,
  {32'h3ebb33ad, 32'h00000000} /* (23, 12, 21) {real, imag} */,
  {32'hbf4f8b24, 32'h00000000} /* (23, 12, 20) {real, imag} */,
  {32'hbfb7da8f, 32'h00000000} /* (23, 12, 19) {real, imag} */,
  {32'hbfc5e550, 32'h00000000} /* (23, 12, 18) {real, imag} */,
  {32'hbfdb680c, 32'h00000000} /* (23, 12, 17) {real, imag} */,
  {32'hbf84eb66, 32'h00000000} /* (23, 12, 16) {real, imag} */,
  {32'hbf070798, 32'h00000000} /* (23, 12, 15) {real, imag} */,
  {32'hbe8b47ca, 32'h00000000} /* (23, 12, 14) {real, imag} */,
  {32'hbf8a7920, 32'h00000000} /* (23, 12, 13) {real, imag} */,
  {32'hbfc4a1cd, 32'h00000000} /* (23, 12, 12) {real, imag} */,
  {32'hbfa3d282, 32'h00000000} /* (23, 12, 11) {real, imag} */,
  {32'h3f12fdb6, 32'h00000000} /* (23, 12, 10) {real, imag} */,
  {32'h3f9f8d66, 32'h00000000} /* (23, 12, 9) {real, imag} */,
  {32'h3fab3df1, 32'h00000000} /* (23, 12, 8) {real, imag} */,
  {32'h3f86cfd5, 32'h00000000} /* (23, 12, 7) {real, imag} */,
  {32'h3f8beabd, 32'h00000000} /* (23, 12, 6) {real, imag} */,
  {32'h3f93175c, 32'h00000000} /* (23, 12, 5) {real, imag} */,
  {32'h3f4e7907, 32'h00000000} /* (23, 12, 4) {real, imag} */,
  {32'h3f6a074e, 32'h00000000} /* (23, 12, 3) {real, imag} */,
  {32'h3f785f93, 32'h00000000} /* (23, 12, 2) {real, imag} */,
  {32'h3f776ee3, 32'h00000000} /* (23, 12, 1) {real, imag} */,
  {32'h3f1364cd, 32'h00000000} /* (23, 12, 0) {real, imag} */,
  {32'h3eb1d8e4, 32'h00000000} /* (23, 11, 31) {real, imag} */,
  {32'h3f584dbd, 32'h00000000} /* (23, 11, 30) {real, imag} */,
  {32'h3f681b99, 32'h00000000} /* (23, 11, 29) {real, imag} */,
  {32'h3fbb6085, 32'h00000000} /* (23, 11, 28) {real, imag} */,
  {32'h3f9f879b, 32'h00000000} /* (23, 11, 27) {real, imag} */,
  {32'h3fa4b6c5, 32'h00000000} /* (23, 11, 26) {real, imag} */,
  {32'h3f84a27b, 32'h00000000} /* (23, 11, 25) {real, imag} */,
  {32'h3f8e381f, 32'h00000000} /* (23, 11, 24) {real, imag} */,
  {32'h3f417d93, 32'h00000000} /* (23, 11, 23) {real, imag} */,
  {32'h3f577cd6, 32'h00000000} /* (23, 11, 22) {real, imag} */,
  {32'hbdab8ba1, 32'h00000000} /* (23, 11, 21) {real, imag} */,
  {32'hbf523f12, 32'h00000000} /* (23, 11, 20) {real, imag} */,
  {32'hbf7f3117, 32'h00000000} /* (23, 11, 19) {real, imag} */,
  {32'hbf007021, 32'h00000000} /* (23, 11, 18) {real, imag} */,
  {32'hbf50fa4e, 32'h00000000} /* (23, 11, 17) {real, imag} */,
  {32'hbf223784, 32'h00000000} /* (23, 11, 16) {real, imag} */,
  {32'hbf2b654e, 32'h00000000} /* (23, 11, 15) {real, imag} */,
  {32'hbf044c45, 32'h00000000} /* (23, 11, 14) {real, imag} */,
  {32'hbf5782f4, 32'h00000000} /* (23, 11, 13) {real, imag} */,
  {32'hbfa94621, 32'h00000000} /* (23, 11, 12) {real, imag} */,
  {32'hbf776c98, 32'h00000000} /* (23, 11, 11) {real, imag} */,
  {32'h3d20c053, 32'h00000000} /* (23, 11, 10) {real, imag} */,
  {32'h3f27b328, 32'h00000000} /* (23, 11, 9) {real, imag} */,
  {32'h3f4da7d3, 32'h00000000} /* (23, 11, 8) {real, imag} */,
  {32'h3f467b2a, 32'h00000000} /* (23, 11, 7) {real, imag} */,
  {32'h3f0f1d75, 32'h00000000} /* (23, 11, 6) {real, imag} */,
  {32'h3ea6a438, 32'h00000000} /* (23, 11, 5) {real, imag} */,
  {32'h3f07f4ab, 32'h00000000} /* (23, 11, 4) {real, imag} */,
  {32'h3f0204c1, 32'h00000000} /* (23, 11, 3) {real, imag} */,
  {32'h3f427a44, 32'h00000000} /* (23, 11, 2) {real, imag} */,
  {32'h3eca2823, 32'h00000000} /* (23, 11, 1) {real, imag} */,
  {32'h3e0dd496, 32'h00000000} /* (23, 11, 0) {real, imag} */,
  {32'hbebbf7bd, 32'h00000000} /* (23, 10, 31) {real, imag} */,
  {32'hbee5f1b3, 32'h00000000} /* (23, 10, 30) {real, imag} */,
  {32'hbe97197b, 32'h00000000} /* (23, 10, 29) {real, imag} */,
  {32'h3d1ad0cd, 32'h00000000} /* (23, 10, 28) {real, imag} */,
  {32'hbdc468ca, 32'h00000000} /* (23, 10, 27) {real, imag} */,
  {32'h3ea13bde, 32'h00000000} /* (23, 10, 26) {real, imag} */,
  {32'h3f25497e, 32'h00000000} /* (23, 10, 25) {real, imag} */,
  {32'h3eb75d7c, 32'h00000000} /* (23, 10, 24) {real, imag} */,
  {32'hbf771b68, 32'h00000000} /* (23, 10, 23) {real, imag} */,
  {32'hbf42bbbd, 32'h00000000} /* (23, 10, 22) {real, imag} */,
  {32'hbf393f60, 32'h00000000} /* (23, 10, 21) {real, imag} */,
  {32'hbe281597, 32'h00000000} /* (23, 10, 20) {real, imag} */,
  {32'h3e4eb003, 32'h00000000} /* (23, 10, 19) {real, imag} */,
  {32'h3f2577ac, 32'h00000000} /* (23, 10, 18) {real, imag} */,
  {32'h3f4ace77, 32'h00000000} /* (23, 10, 17) {real, imag} */,
  {32'h3f4d0655, 32'h00000000} /* (23, 10, 16) {real, imag} */,
  {32'h3f03c6fd, 32'h00000000} /* (23, 10, 15) {real, imag} */,
  {32'h3e79153a, 32'h00000000} /* (23, 10, 14) {real, imag} */,
  {32'h3e82cf13, 32'h00000000} /* (23, 10, 13) {real, imag} */,
  {32'h3e92c90e, 32'h00000000} /* (23, 10, 12) {real, imag} */,
  {32'h3db2f3dd, 32'h00000000} /* (23, 10, 11) {real, imag} */,
  {32'hbee244b9, 32'h00000000} /* (23, 10, 10) {real, imag} */,
  {32'hbe359a00, 32'h00000000} /* (23, 10, 9) {real, imag} */,
  {32'hbdebb4a4, 32'h00000000} /* (23, 10, 8) {real, imag} */,
  {32'hbe7c143a, 32'h00000000} /* (23, 10, 7) {real, imag} */,
  {32'hbf29af5d, 32'h00000000} /* (23, 10, 6) {real, imag} */,
  {32'hbef4bd99, 32'h00000000} /* (23, 10, 5) {real, imag} */,
  {32'hbf4e4a6b, 32'h00000000} /* (23, 10, 4) {real, imag} */,
  {32'hbfaba7ec, 32'h00000000} /* (23, 10, 3) {real, imag} */,
  {32'hbf13d961, 32'h00000000} /* (23, 10, 2) {real, imag} */,
  {32'hbec2c283, 32'h00000000} /* (23, 10, 1) {real, imag} */,
  {32'hbe528b72, 32'h00000000} /* (23, 10, 0) {real, imag} */,
  {32'hbf2e64d9, 32'h00000000} /* (23, 9, 31) {real, imag} */,
  {32'hbfa2c937, 32'h00000000} /* (23, 9, 30) {real, imag} */,
  {32'hbfb1a61e, 32'h00000000} /* (23, 9, 29) {real, imag} */,
  {32'hbf85db17, 32'h00000000} /* (23, 9, 28) {real, imag} */,
  {32'hbf7e2a6e, 32'h00000000} /* (23, 9, 27) {real, imag} */,
  {32'hbf309492, 32'h00000000} /* (23, 9, 26) {real, imag} */,
  {32'hbf197812, 32'h00000000} /* (23, 9, 25) {real, imag} */,
  {32'hbf80fb7a, 32'h00000000} /* (23, 9, 24) {real, imag} */,
  {32'hbf9c2d97, 32'h00000000} /* (23, 9, 23) {real, imag} */,
  {32'hbf90d2cf, 32'h00000000} /* (23, 9, 22) {real, imag} */,
  {32'hbf47224a, 32'h00000000} /* (23, 9, 21) {real, imag} */,
  {32'h3e33f4ea, 32'h00000000} /* (23, 9, 20) {real, imag} */,
  {32'h3f0ac5b2, 32'h00000000} /* (23, 9, 19) {real, imag} */,
  {32'h3f67860f, 32'h00000000} /* (23, 9, 18) {real, imag} */,
  {32'h3f871534, 32'h00000000} /* (23, 9, 17) {real, imag} */,
  {32'h3f810c16, 32'h00000000} /* (23, 9, 16) {real, imag} */,
  {32'h3f9cf9c1, 32'h00000000} /* (23, 9, 15) {real, imag} */,
  {32'h3f786c8b, 32'h00000000} /* (23, 9, 14) {real, imag} */,
  {32'h3f7ffddf, 32'h00000000} /* (23, 9, 13) {real, imag} */,
  {32'h3f9199b2, 32'h00000000} /* (23, 9, 12) {real, imag} */,
  {32'h3ee404ed, 32'h00000000} /* (23, 9, 11) {real, imag} */,
  {32'hbf4c7bb3, 32'h00000000} /* (23, 9, 10) {real, imag} */,
  {32'hbf670ff8, 32'h00000000} /* (23, 9, 9) {real, imag} */,
  {32'hbf9245f6, 32'h00000000} /* (23, 9, 8) {real, imag} */,
  {32'hbf8a49b2, 32'h00000000} /* (23, 9, 7) {real, imag} */,
  {32'hbf84ed04, 32'h00000000} /* (23, 9, 6) {real, imag} */,
  {32'hbf572b0a, 32'h00000000} /* (23, 9, 5) {real, imag} */,
  {32'hbf40a327, 32'h00000000} /* (23, 9, 4) {real, imag} */,
  {32'hbfa89549, 32'h00000000} /* (23, 9, 3) {real, imag} */,
  {32'hbf81616c, 32'h00000000} /* (23, 9, 2) {real, imag} */,
  {32'hbf160e2e, 32'h00000000} /* (23, 9, 1) {real, imag} */,
  {32'hbea1c77d, 32'h00000000} /* (23, 9, 0) {real, imag} */,
  {32'hbf1356d8, 32'h00000000} /* (23, 8, 31) {real, imag} */,
  {32'hbf805f11, 32'h00000000} /* (23, 8, 30) {real, imag} */,
  {32'hbfa39d40, 32'h00000000} /* (23, 8, 29) {real, imag} */,
  {32'hbfa04d43, 32'h00000000} /* (23, 8, 28) {real, imag} */,
  {32'hbfaafab6, 32'h00000000} /* (23, 8, 27) {real, imag} */,
  {32'hbf905d1d, 32'h00000000} /* (23, 8, 26) {real, imag} */,
  {32'hbf7ba8d6, 32'h00000000} /* (23, 8, 25) {real, imag} */,
  {32'hbfc01000, 32'h00000000} /* (23, 8, 24) {real, imag} */,
  {32'hbf9f9036, 32'h00000000} /* (23, 8, 23) {real, imag} */,
  {32'hbf841be7, 32'h00000000} /* (23, 8, 22) {real, imag} */,
  {32'hbef1d31e, 32'h00000000} /* (23, 8, 21) {real, imag} */,
  {32'h3f0db97f, 32'h00000000} /* (23, 8, 20) {real, imag} */,
  {32'h3efc2910, 32'h00000000} /* (23, 8, 19) {real, imag} */,
  {32'h3f1e29f8, 32'h00000000} /* (23, 8, 18) {real, imag} */,
  {32'h3f31c588, 32'h00000000} /* (23, 8, 17) {real, imag} */,
  {32'h3f6f7f89, 32'h00000000} /* (23, 8, 16) {real, imag} */,
  {32'h3fa23d4b, 32'h00000000} /* (23, 8, 15) {real, imag} */,
  {32'h3f25f474, 32'h00000000} /* (23, 8, 14) {real, imag} */,
  {32'h3f8d52ad, 32'h00000000} /* (23, 8, 13) {real, imag} */,
  {32'h3fe63527, 32'h00000000} /* (23, 8, 12) {real, imag} */,
  {32'h3f6efba7, 32'h00000000} /* (23, 8, 11) {real, imag} */,
  {32'hbdee5c91, 32'h00000000} /* (23, 8, 10) {real, imag} */,
  {32'hbf2d447d, 32'h00000000} /* (23, 8, 9) {real, imag} */,
  {32'hbfc68be3, 32'h00000000} /* (23, 8, 8) {real, imag} */,
  {32'hbfcb08d7, 32'h00000000} /* (23, 8, 7) {real, imag} */,
  {32'hbf8f5a8c, 32'h00000000} /* (23, 8, 6) {real, imag} */,
  {32'hbf650123, 32'h00000000} /* (23, 8, 5) {real, imag} */,
  {32'hbf5f7fec, 32'h00000000} /* (23, 8, 4) {real, imag} */,
  {32'hbf92227b, 32'h00000000} /* (23, 8, 3) {real, imag} */,
  {32'hbf667281, 32'h00000000} /* (23, 8, 2) {real, imag} */,
  {32'hbf11675c, 32'h00000000} /* (23, 8, 1) {real, imag} */,
  {32'hbe47f595, 32'h00000000} /* (23, 8, 0) {real, imag} */,
  {32'hbec1cd35, 32'h00000000} /* (23, 7, 31) {real, imag} */,
  {32'hbf18dd03, 32'h00000000} /* (23, 7, 30) {real, imag} */,
  {32'hbf28b8f0, 32'h00000000} /* (23, 7, 29) {real, imag} */,
  {32'hbf88d6d4, 32'h00000000} /* (23, 7, 28) {real, imag} */,
  {32'hbfa607c0, 32'h00000000} /* (23, 7, 27) {real, imag} */,
  {32'hbf9a9763, 32'h00000000} /* (23, 7, 26) {real, imag} */,
  {32'hbf8d4377, 32'h00000000} /* (23, 7, 25) {real, imag} */,
  {32'hbf8f1e86, 32'h00000000} /* (23, 7, 24) {real, imag} */,
  {32'hbfb6781d, 32'h00000000} /* (23, 7, 23) {real, imag} */,
  {32'hbf7ac19a, 32'h00000000} /* (23, 7, 22) {real, imag} */,
  {32'hbc5eee82, 32'h00000000} /* (23, 7, 21) {real, imag} */,
  {32'h3f725a19, 32'h00000000} /* (23, 7, 20) {real, imag} */,
  {32'h3f492599, 32'h00000000} /* (23, 7, 19) {real, imag} */,
  {32'h3eebd61c, 32'h00000000} /* (23, 7, 18) {real, imag} */,
  {32'h3f6f2358, 32'h00000000} /* (23, 7, 17) {real, imag} */,
  {32'h3f8e201d, 32'h00000000} /* (23, 7, 16) {real, imag} */,
  {32'h3f37b640, 32'h00000000} /* (23, 7, 15) {real, imag} */,
  {32'h3f0e1aa2, 32'h00000000} /* (23, 7, 14) {real, imag} */,
  {32'h3f31d1d8, 32'h00000000} /* (23, 7, 13) {real, imag} */,
  {32'h3f4ec413, 32'h00000000} /* (23, 7, 12) {real, imag} */,
  {32'h3f300137, 32'h00000000} /* (23, 7, 11) {real, imag} */,
  {32'hbebb72f6, 32'h00000000} /* (23, 7, 10) {real, imag} */,
  {32'hbf759df3, 32'h00000000} /* (23, 7, 9) {real, imag} */,
  {32'hbf9e6d9e, 32'h00000000} /* (23, 7, 8) {real, imag} */,
  {32'hbf534706, 32'h00000000} /* (23, 7, 7) {real, imag} */,
  {32'hbf9f6025, 32'h00000000} /* (23, 7, 6) {real, imag} */,
  {32'hbf7b26a7, 32'h00000000} /* (23, 7, 5) {real, imag} */,
  {32'hbf364193, 32'h00000000} /* (23, 7, 4) {real, imag} */,
  {32'hbf7cb43b, 32'h00000000} /* (23, 7, 3) {real, imag} */,
  {32'hbf9bfab6, 32'h00000000} /* (23, 7, 2) {real, imag} */,
  {32'hbf4f22df, 32'h00000000} /* (23, 7, 1) {real, imag} */,
  {32'hbe905516, 32'h00000000} /* (23, 7, 0) {real, imag} */,
  {32'hbea63b25, 32'h00000000} /* (23, 6, 31) {real, imag} */,
  {32'hbec2e777, 32'h00000000} /* (23, 6, 30) {real, imag} */,
  {32'hbf361abc, 32'h00000000} /* (23, 6, 29) {real, imag} */,
  {32'hbf634677, 32'h00000000} /* (23, 6, 28) {real, imag} */,
  {32'hbf468b55, 32'h00000000} /* (23, 6, 27) {real, imag} */,
  {32'hbf568abb, 32'h00000000} /* (23, 6, 26) {real, imag} */,
  {32'hbf324d44, 32'h00000000} /* (23, 6, 25) {real, imag} */,
  {32'hbf35bc85, 32'h00000000} /* (23, 6, 24) {real, imag} */,
  {32'hbf8caec4, 32'h00000000} /* (23, 6, 23) {real, imag} */,
  {32'hbf8c8f03, 32'h00000000} /* (23, 6, 22) {real, imag} */,
  {32'hbee5156d, 32'h00000000} /* (23, 6, 21) {real, imag} */,
  {32'h3ecbc98b, 32'h00000000} /* (23, 6, 20) {real, imag} */,
  {32'h3f082d1a, 32'h00000000} /* (23, 6, 19) {real, imag} */,
  {32'h3f2dc86f, 32'h00000000} /* (23, 6, 18) {real, imag} */,
  {32'h3f6f7325, 32'h00000000} /* (23, 6, 17) {real, imag} */,
  {32'h3f7ce345, 32'h00000000} /* (23, 6, 16) {real, imag} */,
  {32'h3f5867ab, 32'h00000000} /* (23, 6, 15) {real, imag} */,
  {32'h3f78e412, 32'h00000000} /* (23, 6, 14) {real, imag} */,
  {32'h3f82eb20, 32'h00000000} /* (23, 6, 13) {real, imag} */,
  {32'h3f824474, 32'h00000000} /* (23, 6, 12) {real, imag} */,
  {32'h3f6de936, 32'h00000000} /* (23, 6, 11) {real, imag} */,
  {32'hbea22ec6, 32'h00000000} /* (23, 6, 10) {real, imag} */,
  {32'hbf695548, 32'h00000000} /* (23, 6, 9) {real, imag} */,
  {32'hbf7d940b, 32'h00000000} /* (23, 6, 8) {real, imag} */,
  {32'hbf6e3926, 32'h00000000} /* (23, 6, 7) {real, imag} */,
  {32'hbf9e2eb5, 32'h00000000} /* (23, 6, 6) {real, imag} */,
  {32'hbf3000fb, 32'h00000000} /* (23, 6, 5) {real, imag} */,
  {32'hbef469e4, 32'h00000000} /* (23, 6, 4) {real, imag} */,
  {32'hbf216ced, 32'h00000000} /* (23, 6, 3) {real, imag} */,
  {32'hbf202db2, 32'h00000000} /* (23, 6, 2) {real, imag} */,
  {32'hbf55457f, 32'h00000000} /* (23, 6, 1) {real, imag} */,
  {32'hbf43573d, 32'h00000000} /* (23, 6, 0) {real, imag} */,
  {32'hbf2e31ec, 32'h00000000} /* (23, 5, 31) {real, imag} */,
  {32'hbf7f05a3, 32'h00000000} /* (23, 5, 30) {real, imag} */,
  {32'hbf9bfe2a, 32'h00000000} /* (23, 5, 29) {real, imag} */,
  {32'hbf8d535d, 32'h00000000} /* (23, 5, 28) {real, imag} */,
  {32'hbf642318, 32'h00000000} /* (23, 5, 27) {real, imag} */,
  {32'hbf7c2833, 32'h00000000} /* (23, 5, 26) {real, imag} */,
  {32'hbf6f265c, 32'h00000000} /* (23, 5, 25) {real, imag} */,
  {32'hbf88cbf2, 32'h00000000} /* (23, 5, 24) {real, imag} */,
  {32'hbf81b882, 32'h00000000} /* (23, 5, 23) {real, imag} */,
  {32'hbf79d2f5, 32'h00000000} /* (23, 5, 22) {real, imag} */,
  {32'hbf354dbe, 32'h00000000} /* (23, 5, 21) {real, imag} */,
  {32'hbf1dc57c, 32'h00000000} /* (23, 5, 20) {real, imag} */,
  {32'hbed55495, 32'h00000000} /* (23, 5, 19) {real, imag} */,
  {32'hbd8dfc59, 32'h00000000} /* (23, 5, 18) {real, imag} */,
  {32'hbde056f4, 32'h00000000} /* (23, 5, 17) {real, imag} */,
  {32'hbe8617f1, 32'h00000000} /* (23, 5, 16) {real, imag} */,
  {32'h3ef103b6, 32'h00000000} /* (23, 5, 15) {real, imag} */,
  {32'h3f5dcbde, 32'h00000000} /* (23, 5, 14) {real, imag} */,
  {32'h3f3aca73, 32'h00000000} /* (23, 5, 13) {real, imag} */,
  {32'h3f12b252, 32'h00000000} /* (23, 5, 12) {real, imag} */,
  {32'h3f61d6c4, 32'h00000000} /* (23, 5, 11) {real, imag} */,
  {32'h3f1f2538, 32'h00000000} /* (23, 5, 10) {real, imag} */,
  {32'h3e89bf31, 32'h00000000} /* (23, 5, 9) {real, imag} */,
  {32'h3e76ff83, 32'h00000000} /* (23, 5, 8) {real, imag} */,
  {32'hbdc15f4e, 32'h00000000} /* (23, 5, 7) {real, imag} */,
  {32'h3de1f452, 32'h00000000} /* (23, 5, 6) {real, imag} */,
  {32'hbef26378, 32'h00000000} /* (23, 5, 5) {real, imag} */,
  {32'hbf25d135, 32'h00000000} /* (23, 5, 4) {real, imag} */,
  {32'hbf677013, 32'h00000000} /* (23, 5, 3) {real, imag} */,
  {32'hbf055252, 32'h00000000} /* (23, 5, 2) {real, imag} */,
  {32'hbf2d9bcc, 32'h00000000} /* (23, 5, 1) {real, imag} */,
  {32'hbf3bac43, 32'h00000000} /* (23, 5, 0) {real, imag} */,
  {32'hbf45c1e6, 32'h00000000} /* (23, 4, 31) {real, imag} */,
  {32'hbfd48bca, 32'h00000000} /* (23, 4, 30) {real, imag} */,
  {32'hbfaa99a9, 32'h00000000} /* (23, 4, 29) {real, imag} */,
  {32'hbf86775f, 32'h00000000} /* (23, 4, 28) {real, imag} */,
  {32'hbf82e759, 32'h00000000} /* (23, 4, 27) {real, imag} */,
  {32'hbfa32bee, 32'h00000000} /* (23, 4, 26) {real, imag} */,
  {32'hbfc92ff5, 32'h00000000} /* (23, 4, 25) {real, imag} */,
  {32'hbfd07299, 32'h00000000} /* (23, 4, 24) {real, imag} */,
  {32'hbf885a6f, 32'h00000000} /* (23, 4, 23) {real, imag} */,
  {32'hbf561424, 32'h00000000} /* (23, 4, 22) {real, imag} */,
  {32'hbf19e05f, 32'h00000000} /* (23, 4, 21) {real, imag} */,
  {32'hbf9cfb69, 32'h00000000} /* (23, 4, 20) {real, imag} */,
  {32'hbf83f746, 32'h00000000} /* (23, 4, 19) {real, imag} */,
  {32'hbf07c334, 32'h00000000} /* (23, 4, 18) {real, imag} */,
  {32'hbf146715, 32'h00000000} /* (23, 4, 17) {real, imag} */,
  {32'hbf1f83fa, 32'h00000000} /* (23, 4, 16) {real, imag} */,
  {32'h3ebf14c2, 32'h00000000} /* (23, 4, 15) {real, imag} */,
  {32'h3f08d986, 32'h00000000} /* (23, 4, 14) {real, imag} */,
  {32'h3f246023, 32'h00000000} /* (23, 4, 13) {real, imag} */,
  {32'h3eceb881, 32'h00000000} /* (23, 4, 12) {real, imag} */,
  {32'h3ed7b41e, 32'h00000000} /* (23, 4, 11) {real, imag} */,
  {32'h3f6806ee, 32'h00000000} /* (23, 4, 10) {real, imag} */,
  {32'h3f6959e1, 32'h00000000} /* (23, 4, 9) {real, imag} */,
  {32'h3f5fe8ef, 32'h00000000} /* (23, 4, 8) {real, imag} */,
  {32'h3f66fd96, 32'h00000000} /* (23, 4, 7) {real, imag} */,
  {32'h3f89cc62, 32'h00000000} /* (23, 4, 6) {real, imag} */,
  {32'hbe7a2f20, 32'h00000000} /* (23, 4, 5) {real, imag} */,
  {32'hbf81149e, 32'h00000000} /* (23, 4, 4) {real, imag} */,
  {32'hbf930125, 32'h00000000} /* (23, 4, 3) {real, imag} */,
  {32'hbf3e1195, 32'h00000000} /* (23, 4, 2) {real, imag} */,
  {32'hbef3caee, 32'h00000000} /* (23, 4, 1) {real, imag} */,
  {32'hbebb1040, 32'h00000000} /* (23, 4, 0) {real, imag} */,
  {32'hbf6862f5, 32'h00000000} /* (23, 3, 31) {real, imag} */,
  {32'hbfd40d56, 32'h00000000} /* (23, 3, 30) {real, imag} */,
  {32'hbf9c68f8, 32'h00000000} /* (23, 3, 29) {real, imag} */,
  {32'hbf8eeb66, 32'h00000000} /* (23, 3, 28) {real, imag} */,
  {32'hbf6f9ed1, 32'h00000000} /* (23, 3, 27) {real, imag} */,
  {32'hbf628e88, 32'h00000000} /* (23, 3, 26) {real, imag} */,
  {32'hbf8974e4, 32'h00000000} /* (23, 3, 25) {real, imag} */,
  {32'hbf836832, 32'h00000000} /* (23, 3, 24) {real, imag} */,
  {32'hbf63f543, 32'h00000000} /* (23, 3, 23) {real, imag} */,
  {32'hbf5c17af, 32'h00000000} /* (23, 3, 22) {real, imag} */,
  {32'hbf0aec07, 32'h00000000} /* (23, 3, 21) {real, imag} */,
  {32'hbf510e85, 32'h00000000} /* (23, 3, 20) {real, imag} */,
  {32'hbf3af88b, 32'h00000000} /* (23, 3, 19) {real, imag} */,
  {32'hbf8f0514, 32'h00000000} /* (23, 3, 18) {real, imag} */,
  {32'hbf663802, 32'h00000000} /* (23, 3, 17) {real, imag} */,
  {32'hbf514c0e, 32'h00000000} /* (23, 3, 16) {real, imag} */,
  {32'h3f201608, 32'h00000000} /* (23, 3, 15) {real, imag} */,
  {32'h3fa4f4ea, 32'h00000000} /* (23, 3, 14) {real, imag} */,
  {32'h3f9255af, 32'h00000000} /* (23, 3, 13) {real, imag} */,
  {32'h3f654526, 32'h00000000} /* (23, 3, 12) {real, imag} */,
  {32'h3f6e1fe1, 32'h00000000} /* (23, 3, 11) {real, imag} */,
  {32'h3f83e8c3, 32'h00000000} /* (23, 3, 10) {real, imag} */,
  {32'h3f1109c3, 32'h00000000} /* (23, 3, 9) {real, imag} */,
  {32'h3eea635c, 32'h00000000} /* (23, 3, 8) {real, imag} */,
  {32'h3f646cc3, 32'h00000000} /* (23, 3, 7) {real, imag} */,
  {32'h3f911755, 32'h00000000} /* (23, 3, 6) {real, imag} */,
  {32'hbe05118a, 32'h00000000} /* (23, 3, 5) {real, imag} */,
  {32'hbfa5000c, 32'h00000000} /* (23, 3, 4) {real, imag} */,
  {32'hbfaded8d, 32'h00000000} /* (23, 3, 3) {real, imag} */,
  {32'hbfc6c57d, 32'h00000000} /* (23, 3, 2) {real, imag} */,
  {32'hbf53bbbb, 32'h00000000} /* (23, 3, 1) {real, imag} */,
  {32'hbf464a61, 32'h00000000} /* (23, 3, 0) {real, imag} */,
  {32'hbf10e20a, 32'h00000000} /* (23, 2, 31) {real, imag} */,
  {32'hbf4a0b78, 32'h00000000} /* (23, 2, 30) {real, imag} */,
  {32'hbf9c313a, 32'h00000000} /* (23, 2, 29) {real, imag} */,
  {32'hbf9b487a, 32'h00000000} /* (23, 2, 28) {real, imag} */,
  {32'hbf8d2513, 32'h00000000} /* (23, 2, 27) {real, imag} */,
  {32'hbfa9756e, 32'h00000000} /* (23, 2, 26) {real, imag} */,
  {32'hbf88885d, 32'h00000000} /* (23, 2, 25) {real, imag} */,
  {32'hbf5ba18b, 32'h00000000} /* (23, 2, 24) {real, imag} */,
  {32'hbf632aa0, 32'h00000000} /* (23, 2, 23) {real, imag} */,
  {32'hbfa3b897, 32'h00000000} /* (23, 2, 22) {real, imag} */,
  {32'hbf75c38b, 32'h00000000} /* (23, 2, 21) {real, imag} */,
  {32'hbf60ddfe, 32'h00000000} /* (23, 2, 20) {real, imag} */,
  {32'hbf9627af, 32'h00000000} /* (23, 2, 19) {real, imag} */,
  {32'hbf9a66b1, 32'h00000000} /* (23, 2, 18) {real, imag} */,
  {32'hbf9acb25, 32'h00000000} /* (23, 2, 17) {real, imag} */,
  {32'hbfb16cb2, 32'h00000000} /* (23, 2, 16) {real, imag} */,
  {32'hbdfc0f8d, 32'h00000000} /* (23, 2, 15) {real, imag} */,
  {32'h3f8e4b5b, 32'h00000000} /* (23, 2, 14) {real, imag} */,
  {32'h3f9ff24f, 32'h00000000} /* (23, 2, 13) {real, imag} */,
  {32'h3f6cdbd3, 32'h00000000} /* (23, 2, 12) {real, imag} */,
  {32'h3f7f692e, 32'h00000000} /* (23, 2, 11) {real, imag} */,
  {32'h3f10e5af, 32'h00000000} /* (23, 2, 10) {real, imag} */,
  {32'h3f00817d, 32'h00000000} /* (23, 2, 9) {real, imag} */,
  {32'h3ee8fcc0, 32'h00000000} /* (23, 2, 8) {real, imag} */,
  {32'h3f113aff, 32'h00000000} /* (23, 2, 7) {real, imag} */,
  {32'h3fa6d306, 32'h00000000} /* (23, 2, 6) {real, imag} */,
  {32'h3cac5349, 32'h00000000} /* (23, 2, 5) {real, imag} */,
  {32'hbf5d4617, 32'h00000000} /* (23, 2, 4) {real, imag} */,
  {32'hbf8c2c90, 32'h00000000} /* (23, 2, 3) {real, imag} */,
  {32'hbfa96e91, 32'h00000000} /* (23, 2, 2) {real, imag} */,
  {32'hbf28343b, 32'h00000000} /* (23, 2, 1) {real, imag} */,
  {32'hbf04cf40, 32'h00000000} /* (23, 2, 0) {real, imag} */,
  {32'hbe1056c7, 32'h00000000} /* (23, 1, 31) {real, imag} */,
  {32'hbec43208, 32'h00000000} /* (23, 1, 30) {real, imag} */,
  {32'hbf62e959, 32'h00000000} /* (23, 1, 29) {real, imag} */,
  {32'hbf5a24a0, 32'h00000000} /* (23, 1, 28) {real, imag} */,
  {32'hbfb53f59, 32'h00000000} /* (23, 1, 27) {real, imag} */,
  {32'hbfbf942b, 32'h00000000} /* (23, 1, 26) {real, imag} */,
  {32'hbf6252dc, 32'h00000000} /* (23, 1, 25) {real, imag} */,
  {32'hbf2eec9e, 32'h00000000} /* (23, 1, 24) {real, imag} */,
  {32'hbf306491, 32'h00000000} /* (23, 1, 23) {real, imag} */,
  {32'hbf1b2915, 32'h00000000} /* (23, 1, 22) {real, imag} */,
  {32'hbed96a10, 32'h00000000} /* (23, 1, 21) {real, imag} */,
  {32'hbf1602d8, 32'h00000000} /* (23, 1, 20) {real, imag} */,
  {32'hbf5e5d30, 32'h00000000} /* (23, 1, 19) {real, imag} */,
  {32'hbf5cd2fb, 32'h00000000} /* (23, 1, 18) {real, imag} */,
  {32'hbf95d06a, 32'h00000000} /* (23, 1, 17) {real, imag} */,
  {32'hbf85da29, 32'h00000000} /* (23, 1, 16) {real, imag} */,
  {32'h3e19a4ee, 32'h00000000} /* (23, 1, 15) {real, imag} */,
  {32'h3f6f389e, 32'h00000000} /* (23, 1, 14) {real, imag} */,
  {32'h3f8009b3, 32'h00000000} /* (23, 1, 13) {real, imag} */,
  {32'h3f8f433b, 32'h00000000} /* (23, 1, 12) {real, imag} */,
  {32'h3f838229, 32'h00000000} /* (23, 1, 11) {real, imag} */,
  {32'h3ed45291, 32'h00000000} /* (23, 1, 10) {real, imag} */,
  {32'h3f6a8cf1, 32'h00000000} /* (23, 1, 9) {real, imag} */,
  {32'h3fccf993, 32'h00000000} /* (23, 1, 8) {real, imag} */,
  {32'h3f812eba, 32'h00000000} /* (23, 1, 7) {real, imag} */,
  {32'h3f828052, 32'h00000000} /* (23, 1, 6) {real, imag} */,
  {32'hbdbbcd70, 32'h00000000} /* (23, 1, 5) {real, imag} */,
  {32'hbefa52ab, 32'h00000000} /* (23, 1, 4) {real, imag} */,
  {32'hbf367d41, 32'h00000000} /* (23, 1, 3) {real, imag} */,
  {32'hbf00e81f, 32'h00000000} /* (23, 1, 2) {real, imag} */,
  {32'hbeaccba2, 32'h00000000} /* (23, 1, 1) {real, imag} */,
  {32'hbe0f0114, 32'h00000000} /* (23, 1, 0) {real, imag} */,
  {32'hbe224a3d, 32'h00000000} /* (23, 0, 31) {real, imag} */,
  {32'hbf0170da, 32'h00000000} /* (23, 0, 30) {real, imag} */,
  {32'hbf1b0042, 32'h00000000} /* (23, 0, 29) {real, imag} */,
  {32'hbeb36992, 32'h00000000} /* (23, 0, 28) {real, imag} */,
  {32'hbf7556bb, 32'h00000000} /* (23, 0, 27) {real, imag} */,
  {32'hbf9e4c4c, 32'h00000000} /* (23, 0, 26) {real, imag} */,
  {32'hbefa9a88, 32'h00000000} /* (23, 0, 25) {real, imag} */,
  {32'hbedf1a82, 32'h00000000} /* (23, 0, 24) {real, imag} */,
  {32'hbedd82f2, 32'h00000000} /* (23, 0, 23) {real, imag} */,
  {32'hbd619bc7, 32'h00000000} /* (23, 0, 22) {real, imag} */,
  {32'h3d58fe67, 32'h00000000} /* (23, 0, 21) {real, imag} */,
  {32'hbeced71d, 32'h00000000} /* (23, 0, 20) {real, imag} */,
  {32'hbedec25e, 32'h00000000} /* (23, 0, 19) {real, imag} */,
  {32'hbedb6a8f, 32'h00000000} /* (23, 0, 18) {real, imag} */,
  {32'hbeece9ac, 32'h00000000} /* (23, 0, 17) {real, imag} */,
  {32'hbdb7f931, 32'h00000000} /* (23, 0, 16) {real, imag} */,
  {32'h3f022091, 32'h00000000} /* (23, 0, 15) {real, imag} */,
  {32'h3f339372, 32'h00000000} /* (23, 0, 14) {real, imag} */,
  {32'h3ebf95a9, 32'h00000000} /* (23, 0, 13) {real, imag} */,
  {32'h3eaaef9c, 32'h00000000} /* (23, 0, 12) {real, imag} */,
  {32'h3e84b49d, 32'h00000000} /* (23, 0, 11) {real, imag} */,
  {32'h3e2eb4f1, 32'h00000000} /* (23, 0, 10) {real, imag} */,
  {32'h3ec6e659, 32'h00000000} /* (23, 0, 9) {real, imag} */,
  {32'h3f7e8372, 32'h00000000} /* (23, 0, 8) {real, imag} */,
  {32'h3eebafd8, 32'h00000000} /* (23, 0, 7) {real, imag} */,
  {32'h3e95eaff, 32'h00000000} /* (23, 0, 6) {real, imag} */,
  {32'h3c6a65ee, 32'h00000000} /* (23, 0, 5) {real, imag} */,
  {32'hbdcc8d4f, 32'h00000000} /* (23, 0, 4) {real, imag} */,
  {32'hbea24250, 32'h00000000} /* (23, 0, 3) {real, imag} */,
  {32'hbe834db5, 32'h00000000} /* (23, 0, 2) {real, imag} */,
  {32'hbe8f0d91, 32'h00000000} /* (23, 0, 1) {real, imag} */,
  {32'hbe0afffc, 32'h00000000} /* (23, 0, 0) {real, imag} */,
  {32'hbeb4a27a, 32'h00000000} /* (22, 31, 31) {real, imag} */,
  {32'hbf12097d, 32'h00000000} /* (22, 31, 30) {real, imag} */,
  {32'hbecad0c4, 32'h00000000} /* (22, 31, 29) {real, imag} */,
  {32'hbec02d7c, 32'h00000000} /* (22, 31, 28) {real, imag} */,
  {32'hbeb7263d, 32'h00000000} /* (22, 31, 27) {real, imag} */,
  {32'hbeedf70e, 32'h00000000} /* (22, 31, 26) {real, imag} */,
  {32'hbeee3e96, 32'h00000000} /* (22, 31, 25) {real, imag} */,
  {32'hbf42e59f, 32'h00000000} /* (22, 31, 24) {real, imag} */,
  {32'hbec45943, 32'h00000000} /* (22, 31, 23) {real, imag} */,
  {32'hbef0276f, 32'h00000000} /* (22, 31, 22) {real, imag} */,
  {32'hbe5228d3, 32'h00000000} /* (22, 31, 21) {real, imag} */,
  {32'h3e9cbf34, 32'h00000000} /* (22, 31, 20) {real, imag} */,
  {32'h3e4ed715, 32'h00000000} /* (22, 31, 19) {real, imag} */,
  {32'h3e88ab24, 32'h00000000} /* (22, 31, 18) {real, imag} */,
  {32'h3dee1e8d, 32'h00000000} /* (22, 31, 17) {real, imag} */,
  {32'h3f05f01f, 32'h00000000} /* (22, 31, 16) {real, imag} */,
  {32'h3f2efa5b, 32'h00000000} /* (22, 31, 15) {real, imag} */,
  {32'h3ec4f599, 32'h00000000} /* (22, 31, 14) {real, imag} */,
  {32'h3f00bfd3, 32'h00000000} /* (22, 31, 13) {real, imag} */,
  {32'h3f188936, 32'h00000000} /* (22, 31, 12) {real, imag} */,
  {32'h3e5fb7b0, 32'h00000000} /* (22, 31, 11) {real, imag} */,
  {32'hbdaa5eba, 32'h00000000} /* (22, 31, 10) {real, imag} */,
  {32'hbefa1ac9, 32'h00000000} /* (22, 31, 9) {real, imag} */,
  {32'hbf19df3b, 32'h00000000} /* (22, 31, 8) {real, imag} */,
  {32'hbe8aed4b, 32'h00000000} /* (22, 31, 7) {real, imag} */,
  {32'hbe1beee4, 32'h00000000} /* (22, 31, 6) {real, imag} */,
  {32'hbe6bb8e3, 32'h00000000} /* (22, 31, 5) {real, imag} */,
  {32'hbe77ad83, 32'h00000000} /* (22, 31, 4) {real, imag} */,
  {32'hbd1236b5, 32'h00000000} /* (22, 31, 3) {real, imag} */,
  {32'hbe4d344b, 32'h00000000} /* (22, 31, 2) {real, imag} */,
  {32'hbf094b6e, 32'h00000000} /* (22, 31, 1) {real, imag} */,
  {32'hbe7a29a1, 32'h00000000} /* (22, 31, 0) {real, imag} */,
  {32'hbef6bcbc, 32'h00000000} /* (22, 30, 31) {real, imag} */,
  {32'hbf37adec, 32'h00000000} /* (22, 30, 30) {real, imag} */,
  {32'hbf58c401, 32'h00000000} /* (22, 30, 29) {real, imag} */,
  {32'hbf61c087, 32'h00000000} /* (22, 30, 28) {real, imag} */,
  {32'hbeb403e8, 32'h00000000} /* (22, 30, 27) {real, imag} */,
  {32'hbed8bfe2, 32'h00000000} /* (22, 30, 26) {real, imag} */,
  {32'hbf903c9b, 32'h00000000} /* (22, 30, 25) {real, imag} */,
  {32'hbfd66603, 32'h00000000} /* (22, 30, 24) {real, imag} */,
  {32'hbf91fc25, 32'h00000000} /* (22, 30, 23) {real, imag} */,
  {32'hbf8b3bcf, 32'h00000000} /* (22, 30, 22) {real, imag} */,
  {32'hbf11bd26, 32'h00000000} /* (22, 30, 21) {real, imag} */,
  {32'h3f79bed9, 32'h00000000} /* (22, 30, 20) {real, imag} */,
  {32'h3f3a88ab, 32'h00000000} /* (22, 30, 19) {real, imag} */,
  {32'h3ef266f6, 32'h00000000} /* (22, 30, 18) {real, imag} */,
  {32'h3ebb661a, 32'h00000000} /* (22, 30, 17) {real, imag} */,
  {32'h3f54a506, 32'h00000000} /* (22, 30, 16) {real, imag} */,
  {32'h3f3f834f, 32'h00000000} /* (22, 30, 15) {real, imag} */,
  {32'h3f412c45, 32'h00000000} /* (22, 30, 14) {real, imag} */,
  {32'h3f993180, 32'h00000000} /* (22, 30, 13) {real, imag} */,
  {32'h3f9d4188, 32'h00000000} /* (22, 30, 12) {real, imag} */,
  {32'h3eaf1b54, 32'h00000000} /* (22, 30, 11) {real, imag} */,
  {32'hbf09331c, 32'h00000000} /* (22, 30, 10) {real, imag} */,
  {32'hbf71f218, 32'h00000000} /* (22, 30, 9) {real, imag} */,
  {32'hbf72aaf2, 32'h00000000} /* (22, 30, 8) {real, imag} */,
  {32'hbee45373, 32'h00000000} /* (22, 30, 7) {real, imag} */,
  {32'hbe95e6de, 32'h00000000} /* (22, 30, 6) {real, imag} */,
  {32'hbf3892b7, 32'h00000000} /* (22, 30, 5) {real, imag} */,
  {32'hbef5e6fe, 32'h00000000} /* (22, 30, 4) {real, imag} */,
  {32'hbe826324, 32'h00000000} /* (22, 30, 3) {real, imag} */,
  {32'hbf17d72e, 32'h00000000} /* (22, 30, 2) {real, imag} */,
  {32'hbf8058eb, 32'h00000000} /* (22, 30, 1) {real, imag} */,
  {32'hbf01687f, 32'h00000000} /* (22, 30, 0) {real, imag} */,
  {32'hbea96902, 32'h00000000} /* (22, 29, 31) {real, imag} */,
  {32'hbf3c5b72, 32'h00000000} /* (22, 29, 30) {real, imag} */,
  {32'hbf4b3c49, 32'h00000000} /* (22, 29, 29) {real, imag} */,
  {32'hbf81b6b8, 32'h00000000} /* (22, 29, 28) {real, imag} */,
  {32'hbf546cf0, 32'h00000000} /* (22, 29, 27) {real, imag} */,
  {32'hbf006869, 32'h00000000} /* (22, 29, 26) {real, imag} */,
  {32'hbf974e6d, 32'h00000000} /* (22, 29, 25) {real, imag} */,
  {32'hbf8ddd39, 32'h00000000} /* (22, 29, 24) {real, imag} */,
  {32'hbf8a30fe, 32'h00000000} /* (22, 29, 23) {real, imag} */,
  {32'hbf8f0a40, 32'h00000000} /* (22, 29, 22) {real, imag} */,
  {32'hbf5e18b9, 32'h00000000} /* (22, 29, 21) {real, imag} */,
  {32'h3f3e053f, 32'h00000000} /* (22, 29, 20) {real, imag} */,
  {32'h3fdc9349, 32'h00000000} /* (22, 29, 19) {real, imag} */,
  {32'h3fa58d10, 32'h00000000} /* (22, 29, 18) {real, imag} */,
  {32'h3f8e2d8f, 32'h00000000} /* (22, 29, 17) {real, imag} */,
  {32'h3f988e58, 32'h00000000} /* (22, 29, 16) {real, imag} */,
  {32'h3f7b60a9, 32'h00000000} /* (22, 29, 15) {real, imag} */,
  {32'h3f46909d, 32'h00000000} /* (22, 29, 14) {real, imag} */,
  {32'h3f6c4128, 32'h00000000} /* (22, 29, 13) {real, imag} */,
  {32'h3fa471c3, 32'h00000000} /* (22, 29, 12) {real, imag} */,
  {32'h3f04f6aa, 32'h00000000} /* (22, 29, 11) {real, imag} */,
  {32'hbed6458e, 32'h00000000} /* (22, 29, 10) {real, imag} */,
  {32'hbf7902ec, 32'h00000000} /* (22, 29, 9) {real, imag} */,
  {32'hbf903ee3, 32'h00000000} /* (22, 29, 8) {real, imag} */,
  {32'hbf2d5864, 32'h00000000} /* (22, 29, 7) {real, imag} */,
  {32'hbf1c704d, 32'h00000000} /* (22, 29, 6) {real, imag} */,
  {32'hbf5f9bd1, 32'h00000000} /* (22, 29, 5) {real, imag} */,
  {32'hbf00c4e8, 32'h00000000} /* (22, 29, 4) {real, imag} */,
  {32'hbe327784, 32'h00000000} /* (22, 29, 3) {real, imag} */,
  {32'hbf82096f, 32'h00000000} /* (22, 29, 2) {real, imag} */,
  {32'hbfbe9598, 32'h00000000} /* (22, 29, 1) {real, imag} */,
  {32'hbf0217b3, 32'h00000000} /* (22, 29, 0) {real, imag} */,
  {32'hbee02f89, 32'h00000000} /* (22, 28, 31) {real, imag} */,
  {32'hbf49a350, 32'h00000000} /* (22, 28, 30) {real, imag} */,
  {32'hbf6ab271, 32'h00000000} /* (22, 28, 29) {real, imag} */,
  {32'hbf80ef65, 32'h00000000} /* (22, 28, 28) {real, imag} */,
  {32'hbf88592b, 32'h00000000} /* (22, 28, 27) {real, imag} */,
  {32'hbf1e5f56, 32'h00000000} /* (22, 28, 26) {real, imag} */,
  {32'hbfa7f7e1, 32'h00000000} /* (22, 28, 25) {real, imag} */,
  {32'hbf93f730, 32'h00000000} /* (22, 28, 24) {real, imag} */,
  {32'hbf933d50, 32'h00000000} /* (22, 28, 23) {real, imag} */,
  {32'hbfbc3b6f, 32'h00000000} /* (22, 28, 22) {real, imag} */,
  {32'hbf467ecc, 32'h00000000} /* (22, 28, 21) {real, imag} */,
  {32'h3f3fae3d, 32'h00000000} /* (22, 28, 20) {real, imag} */,
  {32'h3fe38a62, 32'h00000000} /* (22, 28, 19) {real, imag} */,
  {32'h3fccd4bc, 32'h00000000} /* (22, 28, 18) {real, imag} */,
  {32'h3f839428, 32'h00000000} /* (22, 28, 17) {real, imag} */,
  {32'h3fa56399, 32'h00000000} /* (22, 28, 16) {real, imag} */,
  {32'h3fd37d6d, 32'h00000000} /* (22, 28, 15) {real, imag} */,
  {32'h3f804a23, 32'h00000000} /* (22, 28, 14) {real, imag} */,
  {32'h3f2a080c, 32'h00000000} /* (22, 28, 13) {real, imag} */,
  {32'h3f8e0cbf, 32'h00000000} /* (22, 28, 12) {real, imag} */,
  {32'h3f3550de, 32'h00000000} /* (22, 28, 11) {real, imag} */,
  {32'hbea6dc8e, 32'h00000000} /* (22, 28, 10) {real, imag} */,
  {32'hbf94ab6f, 32'h00000000} /* (22, 28, 9) {real, imag} */,
  {32'hbfae405c, 32'h00000000} /* (22, 28, 8) {real, imag} */,
  {32'hbf84c82f, 32'h00000000} /* (22, 28, 7) {real, imag} */,
  {32'hbf8f7b0a, 32'h00000000} /* (22, 28, 6) {real, imag} */,
  {32'hbfa79ba3, 32'h00000000} /* (22, 28, 5) {real, imag} */,
  {32'hbf78edfa, 32'h00000000} /* (22, 28, 4) {real, imag} */,
  {32'hbf4fac3b, 32'h00000000} /* (22, 28, 3) {real, imag} */,
  {32'hbf87a0a5, 32'h00000000} /* (22, 28, 2) {real, imag} */,
  {32'hbf7b3092, 32'h00000000} /* (22, 28, 1) {real, imag} */,
  {32'hbee97632, 32'h00000000} /* (22, 28, 0) {real, imag} */,
  {32'hbe996012, 32'h00000000} /* (22, 27, 31) {real, imag} */,
  {32'hbf0c4854, 32'h00000000} /* (22, 27, 30) {real, imag} */,
  {32'hbefa97ac, 32'h00000000} /* (22, 27, 29) {real, imag} */,
  {32'hbf824f40, 32'h00000000} /* (22, 27, 28) {real, imag} */,
  {32'hbfc35080, 32'h00000000} /* (22, 27, 27) {real, imag} */,
  {32'hbf6cf635, 32'h00000000} /* (22, 27, 26) {real, imag} */,
  {32'hbf54c0ea, 32'h00000000} /* (22, 27, 25) {real, imag} */,
  {32'hbf77a820, 32'h00000000} /* (22, 27, 24) {real, imag} */,
  {32'hbf2bf700, 32'h00000000} /* (22, 27, 23) {real, imag} */,
  {32'hbf4a64d5, 32'h00000000} /* (22, 27, 22) {real, imag} */,
  {32'hbe436646, 32'h00000000} /* (22, 27, 21) {real, imag} */,
  {32'h3f31264b, 32'h00000000} /* (22, 27, 20) {real, imag} */,
  {32'h3f69d9cb, 32'h00000000} /* (22, 27, 19) {real, imag} */,
  {32'h3f876aad, 32'h00000000} /* (22, 27, 18) {real, imag} */,
  {32'h3f8ed2a0, 32'h00000000} /* (22, 27, 17) {real, imag} */,
  {32'h3f6486ec, 32'h00000000} /* (22, 27, 16) {real, imag} */,
  {32'h3f824df2, 32'h00000000} /* (22, 27, 15) {real, imag} */,
  {32'h3f6d8088, 32'h00000000} /* (22, 27, 14) {real, imag} */,
  {32'h3f8f0101, 32'h00000000} /* (22, 27, 13) {real, imag} */,
  {32'h3f788b7b, 32'h00000000} /* (22, 27, 12) {real, imag} */,
  {32'h3f3a3bc8, 32'h00000000} /* (22, 27, 11) {real, imag} */,
  {32'hbec524c4, 32'h00000000} /* (22, 27, 10) {real, imag} */,
  {32'hbfcc78ca, 32'h00000000} /* (22, 27, 9) {real, imag} */,
  {32'hbfd804ab, 32'h00000000} /* (22, 27, 8) {real, imag} */,
  {32'hbf8d5fd9, 32'h00000000} /* (22, 27, 7) {real, imag} */,
  {32'hbf8848b4, 32'h00000000} /* (22, 27, 6) {real, imag} */,
  {32'hbfd52e1a, 32'h00000000} /* (22, 27, 5) {real, imag} */,
  {32'hbfcf5db3, 32'h00000000} /* (22, 27, 4) {real, imag} */,
  {32'hbfa31abf, 32'h00000000} /* (22, 27, 3) {real, imag} */,
  {32'hbf7ee2fc, 32'h00000000} /* (22, 27, 2) {real, imag} */,
  {32'hbf7387ef, 32'h00000000} /* (22, 27, 1) {real, imag} */,
  {32'hbf35932e, 32'h00000000} /* (22, 27, 0) {real, imag} */,
  {32'hbe29ca43, 32'h00000000} /* (22, 26, 31) {real, imag} */,
  {32'hbef9624d, 32'h00000000} /* (22, 26, 30) {real, imag} */,
  {32'hbf1b434b, 32'h00000000} /* (22, 26, 29) {real, imag} */,
  {32'hbf4e7868, 32'h00000000} /* (22, 26, 28) {real, imag} */,
  {32'hbf8afb90, 32'h00000000} /* (22, 26, 27) {real, imag} */,
  {32'hbf82f957, 32'h00000000} /* (22, 26, 26) {real, imag} */,
  {32'hbf5b1d54, 32'h00000000} /* (22, 26, 25) {real, imag} */,
  {32'hbfb6bdaf, 32'h00000000} /* (22, 26, 24) {real, imag} */,
  {32'hbf9bb285, 32'h00000000} /* (22, 26, 23) {real, imag} */,
  {32'hbf8fcb45, 32'h00000000} /* (22, 26, 22) {real, imag} */,
  {32'hbed1ccfc, 32'h00000000} /* (22, 26, 21) {real, imag} */,
  {32'h3ec78740, 32'h00000000} /* (22, 26, 20) {real, imag} */,
  {32'h3f41c154, 32'h00000000} /* (22, 26, 19) {real, imag} */,
  {32'h3f4fddaa, 32'h00000000} /* (22, 26, 18) {real, imag} */,
  {32'h3f8b1645, 32'h00000000} /* (22, 26, 17) {real, imag} */,
  {32'h3f266f62, 32'h00000000} /* (22, 26, 16) {real, imag} */,
  {32'h3e9f7d65, 32'h00000000} /* (22, 26, 15) {real, imag} */,
  {32'h3f3ee8ed, 32'h00000000} /* (22, 26, 14) {real, imag} */,
  {32'h3f97f460, 32'h00000000} /* (22, 26, 13) {real, imag} */,
  {32'h3f8d32d7, 32'h00000000} /* (22, 26, 12) {real, imag} */,
  {32'h3f676eff, 32'h00000000} /* (22, 26, 11) {real, imag} */,
  {32'hbf18d7d0, 32'h00000000} /* (22, 26, 10) {real, imag} */,
  {32'hbfe5a64f, 32'h00000000} /* (22, 26, 9) {real, imag} */,
  {32'hbf8b2990, 32'h00000000} /* (22, 26, 8) {real, imag} */,
  {32'hbf305878, 32'h00000000} /* (22, 26, 7) {real, imag} */,
  {32'hbf682291, 32'h00000000} /* (22, 26, 6) {real, imag} */,
  {32'hbf3ecc87, 32'h00000000} /* (22, 26, 5) {real, imag} */,
  {32'hbf91be0d, 32'h00000000} /* (22, 26, 4) {real, imag} */,
  {32'hbf8b3e98, 32'h00000000} /* (22, 26, 3) {real, imag} */,
  {32'hbf83fdbf, 32'h00000000} /* (22, 26, 2) {real, imag} */,
  {32'hbf94d1fc, 32'h00000000} /* (22, 26, 1) {real, imag} */,
  {32'hbef6bb66, 32'h00000000} /* (22, 26, 0) {real, imag} */,
  {32'hbec16348, 32'h00000000} /* (22, 25, 31) {real, imag} */,
  {32'hbf46e946, 32'h00000000} /* (22, 25, 30) {real, imag} */,
  {32'hbf642c0a, 32'h00000000} /* (22, 25, 29) {real, imag} */,
  {32'hbf25c1b1, 32'h00000000} /* (22, 25, 28) {real, imag} */,
  {32'hbf3ed168, 32'h00000000} /* (22, 25, 27) {real, imag} */,
  {32'hbf5f71cc, 32'h00000000} /* (22, 25, 26) {real, imag} */,
  {32'hbf419087, 32'h00000000} /* (22, 25, 25) {real, imag} */,
  {32'hbfb9f5ab, 32'h00000000} /* (22, 25, 24) {real, imag} */,
  {32'hbfbd77fb, 32'h00000000} /* (22, 25, 23) {real, imag} */,
  {32'hbfafc380, 32'h00000000} /* (22, 25, 22) {real, imag} */,
  {32'hbf2e0417, 32'h00000000} /* (22, 25, 21) {real, imag} */,
  {32'h3ecb604e, 32'h00000000} /* (22, 25, 20) {real, imag} */,
  {32'h3f6f55aa, 32'h00000000} /* (22, 25, 19) {real, imag} */,
  {32'h3f8824c8, 32'h00000000} /* (22, 25, 18) {real, imag} */,
  {32'h3f92b7fd, 32'h00000000} /* (22, 25, 17) {real, imag} */,
  {32'h3f909d95, 32'h00000000} /* (22, 25, 16) {real, imag} */,
  {32'h3f4ff22a, 32'h00000000} /* (22, 25, 15) {real, imag} */,
  {32'h3f68a46f, 32'h00000000} /* (22, 25, 14) {real, imag} */,
  {32'h3f42e140, 32'h00000000} /* (22, 25, 13) {real, imag} */,
  {32'h3f44cf14, 32'h00000000} /* (22, 25, 12) {real, imag} */,
  {32'h3f053941, 32'h00000000} /* (22, 25, 11) {real, imag} */,
  {32'hbf817ea6, 32'h00000000} /* (22, 25, 10) {real, imag} */,
  {32'hbfaec7b1, 32'h00000000} /* (22, 25, 9) {real, imag} */,
  {32'hbf87f4d3, 32'h00000000} /* (22, 25, 8) {real, imag} */,
  {32'hbf1aea8b, 32'h00000000} /* (22, 25, 7) {real, imag} */,
  {32'hbf7b75b3, 32'h00000000} /* (22, 25, 6) {real, imag} */,
  {32'hbf5aa3e3, 32'h00000000} /* (22, 25, 5) {real, imag} */,
  {32'hbf57d25d, 32'h00000000} /* (22, 25, 4) {real, imag} */,
  {32'hbf52b3cb, 32'h00000000} /* (22, 25, 3) {real, imag} */,
  {32'hbf863965, 32'h00000000} /* (22, 25, 2) {real, imag} */,
  {32'hbf5a84d2, 32'h00000000} /* (22, 25, 1) {real, imag} */,
  {32'hbe5bc282, 32'h00000000} /* (22, 25, 0) {real, imag} */,
  {32'hbe9506bf, 32'h00000000} /* (22, 24, 31) {real, imag} */,
  {32'hbf881445, 32'h00000000} /* (22, 24, 30) {real, imag} */,
  {32'hbf89e2a0, 32'h00000000} /* (22, 24, 29) {real, imag} */,
  {32'hbf6c4082, 32'h00000000} /* (22, 24, 28) {real, imag} */,
  {32'hbf8b1b60, 32'h00000000} /* (22, 24, 27) {real, imag} */,
  {32'hbeff0819, 32'h00000000} /* (22, 24, 26) {real, imag} */,
  {32'hbf26240c, 32'h00000000} /* (22, 24, 25) {real, imag} */,
  {32'hbf2cbfcf, 32'h00000000} /* (22, 24, 24) {real, imag} */,
  {32'hbf6a853e, 32'h00000000} /* (22, 24, 23) {real, imag} */,
  {32'hbfafa4f9, 32'h00000000} /* (22, 24, 22) {real, imag} */,
  {32'hbf22144d, 32'h00000000} /* (22, 24, 21) {real, imag} */,
  {32'h3ed3aeee, 32'h00000000} /* (22, 24, 20) {real, imag} */,
  {32'h3f9bf6b6, 32'h00000000} /* (22, 24, 19) {real, imag} */,
  {32'h3fb1095a, 32'h00000000} /* (22, 24, 18) {real, imag} */,
  {32'h3fa2ffe0, 32'h00000000} /* (22, 24, 17) {real, imag} */,
  {32'h3fcb0a4d, 32'h00000000} /* (22, 24, 16) {real, imag} */,
  {32'h3fb58575, 32'h00000000} /* (22, 24, 15) {real, imag} */,
  {32'h3f74f617, 32'h00000000} /* (22, 24, 14) {real, imag} */,
  {32'h3f0cdc54, 32'h00000000} /* (22, 24, 13) {real, imag} */,
  {32'h3f114ca6, 32'h00000000} /* (22, 24, 12) {real, imag} */,
  {32'h3e9c3367, 32'h00000000} /* (22, 24, 11) {real, imag} */,
  {32'hbf1b446d, 32'h00000000} /* (22, 24, 10) {real, imag} */,
  {32'hbf1aa304, 32'h00000000} /* (22, 24, 9) {real, imag} */,
  {32'hbfa727f6, 32'h00000000} /* (22, 24, 8) {real, imag} */,
  {32'hbf9ab361, 32'h00000000} /* (22, 24, 7) {real, imag} */,
  {32'hbf7b3bfa, 32'h00000000} /* (22, 24, 6) {real, imag} */,
  {32'hbf34f200, 32'h00000000} /* (22, 24, 5) {real, imag} */,
  {32'hbf02ffaa, 32'h00000000} /* (22, 24, 4) {real, imag} */,
  {32'hbf4a358b, 32'h00000000} /* (22, 24, 3) {real, imag} */,
  {32'hbf375843, 32'h00000000} /* (22, 24, 2) {real, imag} */,
  {32'hbe3758f3, 32'h00000000} /* (22, 24, 1) {real, imag} */,
  {32'h3cfce057, 32'h00000000} /* (22, 24, 0) {real, imag} */,
  {32'hbe9ff8dc, 32'h00000000} /* (22, 23, 31) {real, imag} */,
  {32'hbf8c7244, 32'h00000000} /* (22, 23, 30) {real, imag} */,
  {32'hbfa0dba7, 32'h00000000} /* (22, 23, 29) {real, imag} */,
  {32'hbf9a6a12, 32'h00000000} /* (22, 23, 28) {real, imag} */,
  {32'hbf8e270f, 32'h00000000} /* (22, 23, 27) {real, imag} */,
  {32'hbf28a099, 32'h00000000} /* (22, 23, 26) {real, imag} */,
  {32'hbf3b2efe, 32'h00000000} /* (22, 23, 25) {real, imag} */,
  {32'hbf14af66, 32'h00000000} /* (22, 23, 24) {real, imag} */,
  {32'hbfb1b3da, 32'h00000000} /* (22, 23, 23) {real, imag} */,
  {32'hbfa1b43a, 32'h00000000} /* (22, 23, 22) {real, imag} */,
  {32'hbe7d8deb, 32'h00000000} /* (22, 23, 21) {real, imag} */,
  {32'h3f313e3e, 32'h00000000} /* (22, 23, 20) {real, imag} */,
  {32'h3f6fd52c, 32'h00000000} /* (22, 23, 19) {real, imag} */,
  {32'h3f55fbd5, 32'h00000000} /* (22, 23, 18) {real, imag} */,
  {32'h3f4e3366, 32'h00000000} /* (22, 23, 17) {real, imag} */,
  {32'h3f6fd723, 32'h00000000} /* (22, 23, 16) {real, imag} */,
  {32'h3f3c1eae, 32'h00000000} /* (22, 23, 15) {real, imag} */,
  {32'h3f2459ca, 32'h00000000} /* (22, 23, 14) {real, imag} */,
  {32'h3f07cefd, 32'h00000000} /* (22, 23, 13) {real, imag} */,
  {32'h3f303933, 32'h00000000} /* (22, 23, 12) {real, imag} */,
  {32'h3eb25179, 32'h00000000} /* (22, 23, 11) {real, imag} */,
  {32'hbdf7a7ec, 32'h00000000} /* (22, 23, 10) {real, imag} */,
  {32'hbe1eb87e, 32'h00000000} /* (22, 23, 9) {real, imag} */,
  {32'hbf5679c2, 32'h00000000} /* (22, 23, 8) {real, imag} */,
  {32'hbfb51802, 32'h00000000} /* (22, 23, 7) {real, imag} */,
  {32'hbf7b358d, 32'h00000000} /* (22, 23, 6) {real, imag} */,
  {32'hbf826333, 32'h00000000} /* (22, 23, 5) {real, imag} */,
  {32'hbf8b4cf9, 32'h00000000} /* (22, 23, 4) {real, imag} */,
  {32'hbfa5e6e2, 32'h00000000} /* (22, 23, 3) {real, imag} */,
  {32'hbf2fdb2f, 32'h00000000} /* (22, 23, 2) {real, imag} */,
  {32'hbef411a5, 32'h00000000} /* (22, 23, 1) {real, imag} */,
  {32'hbea15114, 32'h00000000} /* (22, 23, 0) {real, imag} */,
  {32'hbec8b615, 32'h00000000} /* (22, 22, 31) {real, imag} */,
  {32'hbf8f13e3, 32'h00000000} /* (22, 22, 30) {real, imag} */,
  {32'hbf929448, 32'h00000000} /* (22, 22, 29) {real, imag} */,
  {32'hbf98463b, 32'h00000000} /* (22, 22, 28) {real, imag} */,
  {32'hbf5f6313, 32'h00000000} /* (22, 22, 27) {real, imag} */,
  {32'hbebd71c7, 32'h00000000} /* (22, 22, 26) {real, imag} */,
  {32'hbef5bfb4, 32'h00000000} /* (22, 22, 25) {real, imag} */,
  {32'hbf15db39, 32'h00000000} /* (22, 22, 24) {real, imag} */,
  {32'hbf95dac5, 32'h00000000} /* (22, 22, 23) {real, imag} */,
  {32'hbf7e3945, 32'h00000000} /* (22, 22, 22) {real, imag} */,
  {32'hbec6fed3, 32'h00000000} /* (22, 22, 21) {real, imag} */,
  {32'h3f633b3a, 32'h00000000} /* (22, 22, 20) {real, imag} */,
  {32'h3f620782, 32'h00000000} /* (22, 22, 19) {real, imag} */,
  {32'h3f4cba49, 32'h00000000} /* (22, 22, 18) {real, imag} */,
  {32'h3f17dd9a, 32'h00000000} /* (22, 22, 17) {real, imag} */,
  {32'h3f34a7c5, 32'h00000000} /* (22, 22, 16) {real, imag} */,
  {32'h3efd7b9c, 32'h00000000} /* (22, 22, 15) {real, imag} */,
  {32'h3eb8668a, 32'h00000000} /* (22, 22, 14) {real, imag} */,
  {32'h3f3f5565, 32'h00000000} /* (22, 22, 13) {real, imag} */,
  {32'h3f8dd52f, 32'h00000000} /* (22, 22, 12) {real, imag} */,
  {32'h3f51904f, 32'h00000000} /* (22, 22, 11) {real, imag} */,
  {32'hbe270d47, 32'h00000000} /* (22, 22, 10) {real, imag} */,
  {32'hbef909b6, 32'h00000000} /* (22, 22, 9) {real, imag} */,
  {32'hbf00f93a, 32'h00000000} /* (22, 22, 8) {real, imag} */,
  {32'hbf6d5e81, 32'h00000000} /* (22, 22, 7) {real, imag} */,
  {32'hbf83fbe8, 32'h00000000} /* (22, 22, 6) {real, imag} */,
  {32'hbf5cc400, 32'h00000000} /* (22, 22, 5) {real, imag} */,
  {32'hbf4969a9, 32'h00000000} /* (22, 22, 4) {real, imag} */,
  {32'hbf62ad0a, 32'h00000000} /* (22, 22, 3) {real, imag} */,
  {32'hbefad8ff, 32'h00000000} /* (22, 22, 2) {real, imag} */,
  {32'hbf7334e0, 32'h00000000} /* (22, 22, 1) {real, imag} */,
  {32'hbf02aedf, 32'h00000000} /* (22, 22, 0) {real, imag} */,
  {32'hbe27fea4, 32'h00000000} /* (22, 21, 31) {real, imag} */,
  {32'hbef374e6, 32'h00000000} /* (22, 21, 30) {real, imag} */,
  {32'hbf13adea, 32'h00000000} /* (22, 21, 29) {real, imag} */,
  {32'hbf1dc412, 32'h00000000} /* (22, 21, 28) {real, imag} */,
  {32'hbe5946e2, 32'h00000000} /* (22, 21, 27) {real, imag} */,
  {32'hbdc2dfcb, 32'h00000000} /* (22, 21, 26) {real, imag} */,
  {32'hbe82b495, 32'h00000000} /* (22, 21, 25) {real, imag} */,
  {32'hbd956b66, 32'h00000000} /* (22, 21, 24) {real, imag} */,
  {32'hbebc78c9, 32'h00000000} /* (22, 21, 23) {real, imag} */,
  {32'hbece9e38, 32'h00000000} /* (22, 21, 22) {real, imag} */,
  {32'hbf0ea1d7, 32'h00000000} /* (22, 21, 21) {real, imag} */,
  {32'h3e80cdd5, 32'h00000000} /* (22, 21, 20) {real, imag} */,
  {32'h3f05610e, 32'h00000000} /* (22, 21, 19) {real, imag} */,
  {32'h3e478096, 32'h00000000} /* (22, 21, 18) {real, imag} */,
  {32'h3e04daf8, 32'h00000000} /* (22, 21, 17) {real, imag} */,
  {32'h3e02f868, 32'h00000000} /* (22, 21, 16) {real, imag} */,
  {32'h3e80f808, 32'h00000000} /* (22, 21, 15) {real, imag} */,
  {32'h3eb4f92c, 32'h00000000} /* (22, 21, 14) {real, imag} */,
  {32'h3f66b3e4, 32'h00000000} /* (22, 21, 13) {real, imag} */,
  {32'h3faa483e, 32'h00000000} /* (22, 21, 12) {real, imag} */,
  {32'h3f2ee549, 32'h00000000} /* (22, 21, 11) {real, imag} */,
  {32'hbed7dcf4, 32'h00000000} /* (22, 21, 10) {real, imag} */,
  {32'h3d223673, 32'h00000000} /* (22, 21, 9) {real, imag} */,
  {32'hbe711fa6, 32'h00000000} /* (22, 21, 8) {real, imag} */,
  {32'hbf236a6c, 32'h00000000} /* (22, 21, 7) {real, imag} */,
  {32'hbf04198a, 32'h00000000} /* (22, 21, 6) {real, imag} */,
  {32'hbed220ce, 32'h00000000} /* (22, 21, 5) {real, imag} */,
  {32'hbe903a12, 32'h00000000} /* (22, 21, 4) {real, imag} */,
  {32'hbe09554c, 32'h00000000} /* (22, 21, 3) {real, imag} */,
  {32'hbe92aaa4, 32'h00000000} /* (22, 21, 2) {real, imag} */,
  {32'hbf4e132c, 32'h00000000} /* (22, 21, 1) {real, imag} */,
  {32'hbeb25671, 32'h00000000} /* (22, 21, 0) {real, imag} */,
  {32'h3f1f7ed5, 32'h00000000} /* (22, 20, 31) {real, imag} */,
  {32'h3f982498, 32'h00000000} /* (22, 20, 30) {real, imag} */,
  {32'h3f8aa62a, 32'h00000000} /* (22, 20, 29) {real, imag} */,
  {32'h3f556d2c, 32'h00000000} /* (22, 20, 28) {real, imag} */,
  {32'h3f9731f6, 32'h00000000} /* (22, 20, 27) {real, imag} */,
  {32'h3f6dbee2, 32'h00000000} /* (22, 20, 26) {real, imag} */,
  {32'h3f77e115, 32'h00000000} /* (22, 20, 25) {real, imag} */,
  {32'h3fa3056a, 32'h00000000} /* (22, 20, 24) {real, imag} */,
  {32'h3f2bd7cc, 32'h00000000} /* (22, 20, 23) {real, imag} */,
  {32'h3e9892e5, 32'h00000000} /* (22, 20, 22) {real, imag} */,
  {32'hbd80a53f, 32'h00000000} /* (22, 20, 21) {real, imag} */,
  {32'hbf0a723c, 32'h00000000} /* (22, 20, 20) {real, imag} */,
  {32'hbf2b0514, 32'h00000000} /* (22, 20, 19) {real, imag} */,
  {32'hbf79aaa9, 32'h00000000} /* (22, 20, 18) {real, imag} */,
  {32'hbfb3184f, 32'h00000000} /* (22, 20, 17) {real, imag} */,
  {32'hbf867c76, 32'h00000000} /* (22, 20, 16) {real, imag} */,
  {32'hbe4ab462, 32'h00000000} /* (22, 20, 15) {real, imag} */,
  {32'hbe0530ca, 32'h00000000} /* (22, 20, 14) {real, imag} */,
  {32'hbf1b3ff6, 32'h00000000} /* (22, 20, 13) {real, imag} */,
  {32'hbe3cbd97, 32'h00000000} /* (22, 20, 12) {real, imag} */,
  {32'hbe0408c2, 32'h00000000} /* (22, 20, 11) {real, imag} */,
  {32'h3e2c8323, 32'h00000000} /* (22, 20, 10) {real, imag} */,
  {32'h3f79b72b, 32'h00000000} /* (22, 20, 9) {real, imag} */,
  {32'h3ed514c5, 32'h00000000} /* (22, 20, 8) {real, imag} */,
  {32'h3eaf69b9, 32'h00000000} /* (22, 20, 7) {real, imag} */,
  {32'h3f4989f3, 32'h00000000} /* (22, 20, 6) {real, imag} */,
  {32'h3f6ffe18, 32'h00000000} /* (22, 20, 5) {real, imag} */,
  {32'h3f8bcf1f, 32'h00000000} /* (22, 20, 4) {real, imag} */,
  {32'h3f81332b, 32'h00000000} /* (22, 20, 3) {real, imag} */,
  {32'h3ef94945, 32'h00000000} /* (22, 20, 2) {real, imag} */,
  {32'h3cf6ab30, 32'h00000000} /* (22, 20, 1) {real, imag} */,
  {32'h3d5d328d, 32'h00000000} /* (22, 20, 0) {real, imag} */,
  {32'h3f0c0ffd, 32'h00000000} /* (22, 19, 31) {real, imag} */,
  {32'h3f27c1f4, 32'h00000000} /* (22, 19, 30) {real, imag} */,
  {32'h3f249ad2, 32'h00000000} /* (22, 19, 29) {real, imag} */,
  {32'h3f6a128f, 32'h00000000} /* (22, 19, 28) {real, imag} */,
  {32'h3fafcf1c, 32'h00000000} /* (22, 19, 27) {real, imag} */,
  {32'h3f5135fe, 32'h00000000} /* (22, 19, 26) {real, imag} */,
  {32'h3f2dfdfc, 32'h00000000} /* (22, 19, 25) {real, imag} */,
  {32'h3f683f80, 32'h00000000} /* (22, 19, 24) {real, imag} */,
  {32'h3f71cbb8, 32'h00000000} /* (22, 19, 23) {real, imag} */,
  {32'h3f514f40, 32'h00000000} /* (22, 19, 22) {real, imag} */,
  {32'h3e122cf8, 32'h00000000} /* (22, 19, 21) {real, imag} */,
  {32'hbf030620, 32'h00000000} /* (22, 19, 20) {real, imag} */,
  {32'hbf01b54e, 32'h00000000} /* (22, 19, 19) {real, imag} */,
  {32'hbf479a52, 32'h00000000} /* (22, 19, 18) {real, imag} */,
  {32'hbf6bf342, 32'h00000000} /* (22, 19, 17) {real, imag} */,
  {32'hbf96a948, 32'h00000000} /* (22, 19, 16) {real, imag} */,
  {32'hbf54eccc, 32'h00000000} /* (22, 19, 15) {real, imag} */,
  {32'hbf6fefba, 32'h00000000} /* (22, 19, 14) {real, imag} */,
  {32'hbfcfac19, 32'h00000000} /* (22, 19, 13) {real, imag} */,
  {32'hbfce09ee, 32'h00000000} /* (22, 19, 12) {real, imag} */,
  {32'hbf4e4179, 32'h00000000} /* (22, 19, 11) {real, imag} */,
  {32'h3d0083f4, 32'h00000000} /* (22, 19, 10) {real, imag} */,
  {32'h3f16b452, 32'h00000000} /* (22, 19, 9) {real, imag} */,
  {32'h3ecebdbc, 32'h00000000} /* (22, 19, 8) {real, imag} */,
  {32'h3f477180, 32'h00000000} /* (22, 19, 7) {real, imag} */,
  {32'h3f9677af, 32'h00000000} /* (22, 19, 6) {real, imag} */,
  {32'h3f947145, 32'h00000000} /* (22, 19, 5) {real, imag} */,
  {32'h3f9b6d4b, 32'h00000000} /* (22, 19, 4) {real, imag} */,
  {32'h3f87f99d, 32'h00000000} /* (22, 19, 3) {real, imag} */,
  {32'h3f487a53, 32'h00000000} /* (22, 19, 2) {real, imag} */,
  {32'h3ea7a0b5, 32'h00000000} /* (22, 19, 1) {real, imag} */,
  {32'h3e115bd9, 32'h00000000} /* (22, 19, 0) {real, imag} */,
  {32'h3f233a71, 32'h00000000} /* (22, 18, 31) {real, imag} */,
  {32'h3f578eb7, 32'h00000000} /* (22, 18, 30) {real, imag} */,
  {32'h3f4d1626, 32'h00000000} /* (22, 18, 29) {real, imag} */,
  {32'h3f75a9e5, 32'h00000000} /* (22, 18, 28) {real, imag} */,
  {32'h3f50df9e, 32'h00000000} /* (22, 18, 27) {real, imag} */,
  {32'h3f20ad17, 32'h00000000} /* (22, 18, 26) {real, imag} */,
  {32'h3f4d9222, 32'h00000000} /* (22, 18, 25) {real, imag} */,
  {32'h3f3644b9, 32'h00000000} /* (22, 18, 24) {real, imag} */,
  {32'h3f280789, 32'h00000000} /* (22, 18, 23) {real, imag} */,
  {32'h3eba1a78, 32'h00000000} /* (22, 18, 22) {real, imag} */,
  {32'h3cb16769, 32'h00000000} /* (22, 18, 21) {real, imag} */,
  {32'hbe991e75, 32'h00000000} /* (22, 18, 20) {real, imag} */,
  {32'hbf4c1bc3, 32'h00000000} /* (22, 18, 19) {real, imag} */,
  {32'hbfa34968, 32'h00000000} /* (22, 18, 18) {real, imag} */,
  {32'hbf35f3c7, 32'h00000000} /* (22, 18, 17) {real, imag} */,
  {32'hbf8e6c5b, 32'h00000000} /* (22, 18, 16) {real, imag} */,
  {32'hbfaa8482, 32'h00000000} /* (22, 18, 15) {real, imag} */,
  {32'hbf9c1ff9, 32'h00000000} /* (22, 18, 14) {real, imag} */,
  {32'hbfa2b6aa, 32'h00000000} /* (22, 18, 13) {real, imag} */,
  {32'hbfc46eca, 32'h00000000} /* (22, 18, 12) {real, imag} */,
  {32'hbf9d8085, 32'h00000000} /* (22, 18, 11) {real, imag} */,
  {32'hbebc4a68, 32'h00000000} /* (22, 18, 10) {real, imag} */,
  {32'h3f42e69a, 32'h00000000} /* (22, 18, 9) {real, imag} */,
  {32'h3fa7d257, 32'h00000000} /* (22, 18, 8) {real, imag} */,
  {32'h3fbbdf89, 32'h00000000} /* (22, 18, 7) {real, imag} */,
  {32'h3f9076af, 32'h00000000} /* (22, 18, 6) {real, imag} */,
  {32'h3f40f11b, 32'h00000000} /* (22, 18, 5) {real, imag} */,
  {32'h3f24273b, 32'h00000000} /* (22, 18, 4) {real, imag} */,
  {32'h3edc30a6, 32'h00000000} /* (22, 18, 3) {real, imag} */,
  {32'h3f64867f, 32'h00000000} /* (22, 18, 2) {real, imag} */,
  {32'h3f809411, 32'h00000000} /* (22, 18, 1) {real, imag} */,
  {32'h3ebc0a2e, 32'h00000000} /* (22, 18, 0) {real, imag} */,
  {32'h3f3aeba8, 32'h00000000} /* (22, 17, 31) {real, imag} */,
  {32'h3f49889b, 32'h00000000} /* (22, 17, 30) {real, imag} */,
  {32'h3f5fc3ed, 32'h00000000} /* (22, 17, 29) {real, imag} */,
  {32'h3f572246, 32'h00000000} /* (22, 17, 28) {real, imag} */,
  {32'h3e6d9626, 32'h00000000} /* (22, 17, 27) {real, imag} */,
  {32'h3eaca1d6, 32'h00000000} /* (22, 17, 26) {real, imag} */,
  {32'h3f923a30, 32'h00000000} /* (22, 17, 25) {real, imag} */,
  {32'h3faf5647, 32'h00000000} /* (22, 17, 24) {real, imag} */,
  {32'h3fb5266b, 32'h00000000} /* (22, 17, 23) {real, imag} */,
  {32'h3f31b5fb, 32'h00000000} /* (22, 17, 22) {real, imag} */,
  {32'h3cd95d99, 32'h00000000} /* (22, 17, 21) {real, imag} */,
  {32'hbf0857f8, 32'h00000000} /* (22, 17, 20) {real, imag} */,
  {32'hbfb9994d, 32'h00000000} /* (22, 17, 19) {real, imag} */,
  {32'hbffa04e1, 32'h00000000} /* (22, 17, 18) {real, imag} */,
  {32'hbf8a78d6, 32'h00000000} /* (22, 17, 17) {real, imag} */,
  {32'hbf519bde, 32'h00000000} /* (22, 17, 16) {real, imag} */,
  {32'hbf7bf337, 32'h00000000} /* (22, 17, 15) {real, imag} */,
  {32'hbf82c4f2, 32'h00000000} /* (22, 17, 14) {real, imag} */,
  {32'hbf9c82a1, 32'h00000000} /* (22, 17, 13) {real, imag} */,
  {32'hbfe5252a, 32'h00000000} /* (22, 17, 12) {real, imag} */,
  {32'hbfa53ac0, 32'h00000000} /* (22, 17, 11) {real, imag} */,
  {32'hbe5648e4, 32'h00000000} /* (22, 17, 10) {real, imag} */,
  {32'h3f9edeb8, 32'h00000000} /* (22, 17, 9) {real, imag} */,
  {32'h3fbf4648, 32'h00000000} /* (22, 17, 8) {real, imag} */,
  {32'h3f9cd173, 32'h00000000} /* (22, 17, 7) {real, imag} */,
  {32'h3f7018d3, 32'h00000000} /* (22, 17, 6) {real, imag} */,
  {32'h3f613a8a, 32'h00000000} /* (22, 17, 5) {real, imag} */,
  {32'h3f66cfcb, 32'h00000000} /* (22, 17, 4) {real, imag} */,
  {32'h3f0bd3bc, 32'h00000000} /* (22, 17, 3) {real, imag} */,
  {32'h3f787f19, 32'h00000000} /* (22, 17, 2) {real, imag} */,
  {32'h3f9d3041, 32'h00000000} /* (22, 17, 1) {real, imag} */,
  {32'h3f26e204, 32'h00000000} /* (22, 17, 0) {real, imag} */,
  {32'h3f2dd883, 32'h00000000} /* (22, 16, 31) {real, imag} */,
  {32'h3f899814, 32'h00000000} /* (22, 16, 30) {real, imag} */,
  {32'h3f590425, 32'h00000000} /* (22, 16, 29) {real, imag} */,
  {32'h3efe60d9, 32'h00000000} /* (22, 16, 28) {real, imag} */,
  {32'h3ea9916c, 32'h00000000} /* (22, 16, 27) {real, imag} */,
  {32'h3f41b273, 32'h00000000} /* (22, 16, 26) {real, imag} */,
  {32'h3fa907b4, 32'h00000000} /* (22, 16, 25) {real, imag} */,
  {32'h3fa78a2f, 32'h00000000} /* (22, 16, 24) {real, imag} */,
  {32'h3fd9d38d, 32'h00000000} /* (22, 16, 23) {real, imag} */,
  {32'h3f9b292a, 32'h00000000} /* (22, 16, 22) {real, imag} */,
  {32'hbe17dd1f, 32'h00000000} /* (22, 16, 21) {real, imag} */,
  {32'hbf9cdf1a, 32'h00000000} /* (22, 16, 20) {real, imag} */,
  {32'hbfc900d0, 32'h00000000} /* (22, 16, 19) {real, imag} */,
  {32'hbfe9c51c, 32'h00000000} /* (22, 16, 18) {real, imag} */,
  {32'hbf81c02a, 32'h00000000} /* (22, 16, 17) {real, imag} */,
  {32'hbf2cf14d, 32'h00000000} /* (22, 16, 16) {real, imag} */,
  {32'hbf1934db, 32'h00000000} /* (22, 16, 15) {real, imag} */,
  {32'hbee5a59a, 32'h00000000} /* (22, 16, 14) {real, imag} */,
  {32'hbf6304ed, 32'h00000000} /* (22, 16, 13) {real, imag} */,
  {32'hbfa4c400, 32'h00000000} /* (22, 16, 12) {real, imag} */,
  {32'hbf9ee117, 32'h00000000} /* (22, 16, 11) {real, imag} */,
  {32'hbe6511cf, 32'h00000000} /* (22, 16, 10) {real, imag} */,
  {32'h3f95555b, 32'h00000000} /* (22, 16, 9) {real, imag} */,
  {32'h3f58df3a, 32'h00000000} /* (22, 16, 8) {real, imag} */,
  {32'h3f28204a, 32'h00000000} /* (22, 16, 7) {real, imag} */,
  {32'h3f3fe0a2, 32'h00000000} /* (22, 16, 6) {real, imag} */,
  {32'h3f5015e3, 32'h00000000} /* (22, 16, 5) {real, imag} */,
  {32'h3f883e92, 32'h00000000} /* (22, 16, 4) {real, imag} */,
  {32'h3f7a1b5a, 32'h00000000} /* (22, 16, 3) {real, imag} */,
  {32'h3f2910d2, 32'h00000000} /* (22, 16, 2) {real, imag} */,
  {32'h3f59c6cd, 32'h00000000} /* (22, 16, 1) {real, imag} */,
  {32'h3ed4a803, 32'h00000000} /* (22, 16, 0) {real, imag} */,
  {32'h3ed89784, 32'h00000000} /* (22, 15, 31) {real, imag} */,
  {32'h3f97cdd1, 32'h00000000} /* (22, 15, 30) {real, imag} */,
  {32'h3f90bdca, 32'h00000000} /* (22, 15, 29) {real, imag} */,
  {32'h3f6ff7f5, 32'h00000000} /* (22, 15, 28) {real, imag} */,
  {32'h3f53f227, 32'h00000000} /* (22, 15, 27) {real, imag} */,
  {32'h3f7e04de, 32'h00000000} /* (22, 15, 26) {real, imag} */,
  {32'h3f8c9d49, 32'h00000000} /* (22, 15, 25) {real, imag} */,
  {32'h3f83dda3, 32'h00000000} /* (22, 15, 24) {real, imag} */,
  {32'h3f9df594, 32'h00000000} /* (22, 15, 23) {real, imag} */,
  {32'h3f36d758, 32'h00000000} /* (22, 15, 22) {real, imag} */,
  {32'hbeacbc25, 32'h00000000} /* (22, 15, 21) {real, imag} */,
  {32'hbfb1e366, 32'h00000000} /* (22, 15, 20) {real, imag} */,
  {32'hbf91e388, 32'h00000000} /* (22, 15, 19) {real, imag} */,
  {32'hbf86ae75, 32'h00000000} /* (22, 15, 18) {real, imag} */,
  {32'hbf7fe54d, 32'h00000000} /* (22, 15, 17) {real, imag} */,
  {32'hbf6d7188, 32'h00000000} /* (22, 15, 16) {real, imag} */,
  {32'hbefd93af, 32'h00000000} /* (22, 15, 15) {real, imag} */,
  {32'hbe8a5948, 32'h00000000} /* (22, 15, 14) {real, imag} */,
  {32'hbf2e0467, 32'h00000000} /* (22, 15, 13) {real, imag} */,
  {32'hbfb8519a, 32'h00000000} /* (22, 15, 12) {real, imag} */,
  {32'hbfced5f8, 32'h00000000} /* (22, 15, 11) {real, imag} */,
  {32'hbec012b5, 32'h00000000} /* (22, 15, 10) {real, imag} */,
  {32'h3f381d05, 32'h00000000} /* (22, 15, 9) {real, imag} */,
  {32'h3f6da7b9, 32'h00000000} /* (22, 15, 8) {real, imag} */,
  {32'h3f4134cb, 32'h00000000} /* (22, 15, 7) {real, imag} */,
  {32'h3f044a0f, 32'h00000000} /* (22, 15, 6) {real, imag} */,
  {32'h3f1f6704, 32'h00000000} /* (22, 15, 5) {real, imag} */,
  {32'h3faf51fa, 32'h00000000} /* (22, 15, 4) {real, imag} */,
  {32'h3fb5766b, 32'h00000000} /* (22, 15, 3) {real, imag} */,
  {32'h3f450ce4, 32'h00000000} /* (22, 15, 2) {real, imag} */,
  {32'h3f4c228b, 32'h00000000} /* (22, 15, 1) {real, imag} */,
  {32'h3eaddab4, 32'h00000000} /* (22, 15, 0) {real, imag} */,
  {32'h3f152264, 32'h00000000} /* (22, 14, 31) {real, imag} */,
  {32'h3fad5c63, 32'h00000000} /* (22, 14, 30) {real, imag} */,
  {32'h3f9ceab7, 32'h00000000} /* (22, 14, 29) {real, imag} */,
  {32'h3f4bcc24, 32'h00000000} /* (22, 14, 28) {real, imag} */,
  {32'h3f44477b, 32'h00000000} /* (22, 14, 27) {real, imag} */,
  {32'h3faa19d4, 32'h00000000} /* (22, 14, 26) {real, imag} */,
  {32'h3fa7573b, 32'h00000000} /* (22, 14, 25) {real, imag} */,
  {32'h3f977fdb, 32'h00000000} /* (22, 14, 24) {real, imag} */,
  {32'h3fc4a4eb, 32'h00000000} /* (22, 14, 23) {real, imag} */,
  {32'h3fa1810a, 32'h00000000} /* (22, 14, 22) {real, imag} */,
  {32'hbd75c625, 32'h00000000} /* (22, 14, 21) {real, imag} */,
  {32'hbf6c15f0, 32'h00000000} /* (22, 14, 20) {real, imag} */,
  {32'hbf1e6414, 32'h00000000} /* (22, 14, 19) {real, imag} */,
  {32'hbf2c6cd9, 32'h00000000} /* (22, 14, 18) {real, imag} */,
  {32'hbf402fc8, 32'h00000000} /* (22, 14, 17) {real, imag} */,
  {32'hbf5b818b, 32'h00000000} /* (22, 14, 16) {real, imag} */,
  {32'hbf465398, 32'h00000000} /* (22, 14, 15) {real, imag} */,
  {32'hbe90f589, 32'h00000000} /* (22, 14, 14) {real, imag} */,
  {32'hbf3317cf, 32'h00000000} /* (22, 14, 13) {real, imag} */,
  {32'hbfa3eedb, 32'h00000000} /* (22, 14, 12) {real, imag} */,
  {32'hbf8f3aa6, 32'h00000000} /* (22, 14, 11) {real, imag} */,
  {32'h3e8e0338, 32'h00000000} /* (22, 14, 10) {real, imag} */,
  {32'h3f7aae74, 32'h00000000} /* (22, 14, 9) {real, imag} */,
  {32'h3fa322bf, 32'h00000000} /* (22, 14, 8) {real, imag} */,
  {32'h3f9d3a6f, 32'h00000000} /* (22, 14, 7) {real, imag} */,
  {32'h3f08f93d, 32'h00000000} /* (22, 14, 6) {real, imag} */,
  {32'h3f0e4081, 32'h00000000} /* (22, 14, 5) {real, imag} */,
  {32'h3f886fe4, 32'h00000000} /* (22, 14, 4) {real, imag} */,
  {32'h3f6ce771, 32'h00000000} /* (22, 14, 3) {real, imag} */,
  {32'h3f272559, 32'h00000000} /* (22, 14, 2) {real, imag} */,
  {32'h3f93a071, 32'h00000000} /* (22, 14, 1) {real, imag} */,
  {32'h3f8a954e, 32'h00000000} /* (22, 14, 0) {real, imag} */,
  {32'h3f205a43, 32'h00000000} /* (22, 13, 31) {real, imag} */,
  {32'h3f891004, 32'h00000000} /* (22, 13, 30) {real, imag} */,
  {32'h3f8d2632, 32'h00000000} /* (22, 13, 29) {real, imag} */,
  {32'h3f698802, 32'h00000000} /* (22, 13, 28) {real, imag} */,
  {32'h3f5211d2, 32'h00000000} /* (22, 13, 27) {real, imag} */,
  {32'h3f919daa, 32'h00000000} /* (22, 13, 26) {real, imag} */,
  {32'h3f506503, 32'h00000000} /* (22, 13, 25) {real, imag} */,
  {32'h3f17e294, 32'h00000000} /* (22, 13, 24) {real, imag} */,
  {32'h3f84a6b8, 32'h00000000} /* (22, 13, 23) {real, imag} */,
  {32'h3fd4032b, 32'h00000000} /* (22, 13, 22) {real, imag} */,
  {32'h3f0ba2fd, 32'h00000000} /* (22, 13, 21) {real, imag} */,
  {32'hbf420074, 32'h00000000} /* (22, 13, 20) {real, imag} */,
  {32'hbfbb2849, 32'h00000000} /* (22, 13, 19) {real, imag} */,
  {32'hbf8a684b, 32'h00000000} /* (22, 13, 18) {real, imag} */,
  {32'hbf587315, 32'h00000000} /* (22, 13, 17) {real, imag} */,
  {32'hbf56b8e7, 32'h00000000} /* (22, 13, 16) {real, imag} */,
  {32'hbeb8a74a, 32'h00000000} /* (22, 13, 15) {real, imag} */,
  {32'hbe270bed, 32'h00000000} /* (22, 13, 14) {real, imag} */,
  {32'hbf0289ae, 32'h00000000} /* (22, 13, 13) {real, imag} */,
  {32'hbf679492, 32'h00000000} /* (22, 13, 12) {real, imag} */,
  {32'hbf7b5041, 32'h00000000} /* (22, 13, 11) {real, imag} */,
  {32'h3f246f8d, 32'h00000000} /* (22, 13, 10) {real, imag} */,
  {32'h3fb0f8e7, 32'h00000000} /* (22, 13, 9) {real, imag} */,
  {32'h3fc63bed, 32'h00000000} /* (22, 13, 8) {real, imag} */,
  {32'h3fb6b1c0, 32'h00000000} /* (22, 13, 7) {real, imag} */,
  {32'h3f5dce74, 32'h00000000} /* (22, 13, 6) {real, imag} */,
  {32'h3f873394, 32'h00000000} /* (22, 13, 5) {real, imag} */,
  {32'h3f584a64, 32'h00000000} /* (22, 13, 4) {real, imag} */,
  {32'h3f10d648, 32'h00000000} /* (22, 13, 3) {real, imag} */,
  {32'h3eef9269, 32'h00000000} /* (22, 13, 2) {real, imag} */,
  {32'h3f87085a, 32'h00000000} /* (22, 13, 1) {real, imag} */,
  {32'h3f64d9fb, 32'h00000000} /* (22, 13, 0) {real, imag} */,
  {32'h3f01c18f, 32'h00000000} /* (22, 12, 31) {real, imag} */,
  {32'h3ef87f9e, 32'h00000000} /* (22, 12, 30) {real, imag} */,
  {32'h3f16c790, 32'h00000000} /* (22, 12, 29) {real, imag} */,
  {32'h3f98ddb5, 32'h00000000} /* (22, 12, 28) {real, imag} */,
  {32'h3f8c37a9, 32'h00000000} /* (22, 12, 27) {real, imag} */,
  {32'h3f3dc579, 32'h00000000} /* (22, 12, 26) {real, imag} */,
  {32'h3ed5461e, 32'h00000000} /* (22, 12, 25) {real, imag} */,
  {32'h3f598c4b, 32'h00000000} /* (22, 12, 24) {real, imag} */,
  {32'h3fd16be5, 32'h00000000} /* (22, 12, 23) {real, imag} */,
  {32'h3fdad285, 32'h00000000} /* (22, 12, 22) {real, imag} */,
  {32'h3ec36fc6, 32'h00000000} /* (22, 12, 21) {real, imag} */,
  {32'hbf7b08b8, 32'h00000000} /* (22, 12, 20) {real, imag} */,
  {32'hbff4a8e5, 32'h00000000} /* (22, 12, 19) {real, imag} */,
  {32'hbfc4ccdd, 32'h00000000} /* (22, 12, 18) {real, imag} */,
  {32'hbf86ea67, 32'h00000000} /* (22, 12, 17) {real, imag} */,
  {32'hbf4485b1, 32'h00000000} /* (22, 12, 16) {real, imag} */,
  {32'hbe7bb679, 32'h00000000} /* (22, 12, 15) {real, imag} */,
  {32'hbed0578d, 32'h00000000} /* (22, 12, 14) {real, imag} */,
  {32'hbf1ca309, 32'h00000000} /* (22, 12, 13) {real, imag} */,
  {32'hbf8d0934, 32'h00000000} /* (22, 12, 12) {real, imag} */,
  {32'hbf402b27, 32'h00000000} /* (22, 12, 11) {real, imag} */,
  {32'h3f6aa314, 32'h00000000} /* (22, 12, 10) {real, imag} */,
  {32'h3f4cf1ef, 32'h00000000} /* (22, 12, 9) {real, imag} */,
  {32'h3f8f3088, 32'h00000000} /* (22, 12, 8) {real, imag} */,
  {32'h3fa74d36, 32'h00000000} /* (22, 12, 7) {real, imag} */,
  {32'h3f83e3a8, 32'h00000000} /* (22, 12, 6) {real, imag} */,
  {32'h3fa8621b, 32'h00000000} /* (22, 12, 5) {real, imag} */,
  {32'h3f5209f0, 32'h00000000} /* (22, 12, 4) {real, imag} */,
  {32'h3f2291b3, 32'h00000000} /* (22, 12, 3) {real, imag} */,
  {32'h3f2b3c26, 32'h00000000} /* (22, 12, 2) {real, imag} */,
  {32'h3f4e59e9, 32'h00000000} /* (22, 12, 1) {real, imag} */,
  {32'h3e5e796a, 32'h00000000} /* (22, 12, 0) {real, imag} */,
  {32'h3e7d86c4, 32'h00000000} /* (22, 11, 31) {real, imag} */,
  {32'h3e5840db, 32'h00000000} /* (22, 11, 30) {real, imag} */,
  {32'h3e7f5c4c, 32'h00000000} /* (22, 11, 29) {real, imag} */,
  {32'h3f2b0973, 32'h00000000} /* (22, 11, 28) {real, imag} */,
  {32'h3f4ff436, 32'h00000000} /* (22, 11, 27) {real, imag} */,
  {32'h3f67a1aa, 32'h00000000} /* (22, 11, 26) {real, imag} */,
  {32'h3ef4910a, 32'h00000000} /* (22, 11, 25) {real, imag} */,
  {32'h3f64abac, 32'h00000000} /* (22, 11, 24) {real, imag} */,
  {32'h3f883a1e, 32'h00000000} /* (22, 11, 23) {real, imag} */,
  {32'h3f82b602, 32'h00000000} /* (22, 11, 22) {real, imag} */,
  {32'hbe990fd2, 32'h00000000} /* (22, 11, 21) {real, imag} */,
  {32'hbf872e30, 32'h00000000} /* (22, 11, 20) {real, imag} */,
  {32'hbf7b38a6, 32'h00000000} /* (22, 11, 19) {real, imag} */,
  {32'hbf161188, 32'h00000000} /* (22, 11, 18) {real, imag} */,
  {32'hbf146895, 32'h00000000} /* (22, 11, 17) {real, imag} */,
  {32'hbf239b41, 32'h00000000} /* (22, 11, 16) {real, imag} */,
  {32'hbf196a35, 32'h00000000} /* (22, 11, 15) {real, imag} */,
  {32'hbf0c92ad, 32'h00000000} /* (22, 11, 14) {real, imag} */,
  {32'hbf1f9f1f, 32'h00000000} /* (22, 11, 13) {real, imag} */,
  {32'hbf88d574, 32'h00000000} /* (22, 11, 12) {real, imag} */,
  {32'hbf118742, 32'h00000000} /* (22, 11, 11) {real, imag} */,
  {32'h3f20f8a5, 32'h00000000} /* (22, 11, 10) {real, imag} */,
  {32'h3f0455a5, 32'h00000000} /* (22, 11, 9) {real, imag} */,
  {32'h3fae57ad, 32'h00000000} /* (22, 11, 8) {real, imag} */,
  {32'h3faaf817, 32'h00000000} /* (22, 11, 7) {real, imag} */,
  {32'h3ef6de82, 32'h00000000} /* (22, 11, 6) {real, imag} */,
  {32'h3f29298f, 32'h00000000} /* (22, 11, 5) {real, imag} */,
  {32'h3f431abc, 32'h00000000} /* (22, 11, 4) {real, imag} */,
  {32'h3f1ec2b2, 32'h00000000} /* (22, 11, 3) {real, imag} */,
  {32'h3f0d3d03, 32'h00000000} /* (22, 11, 2) {real, imag} */,
  {32'h3f2bcd60, 32'h00000000} /* (22, 11, 1) {real, imag} */,
  {32'h3eac710c, 32'h00000000} /* (22, 11, 0) {real, imag} */,
  {32'hbeb1d7fa, 32'h00000000} /* (22, 10, 31) {real, imag} */,
  {32'hbf38d3b8, 32'h00000000} /* (22, 10, 30) {real, imag} */,
  {32'hbf4cb102, 32'h00000000} /* (22, 10, 29) {real, imag} */,
  {32'hbebe5fbd, 32'h00000000} /* (22, 10, 28) {real, imag} */,
  {32'hbe95dfb8, 32'h00000000} /* (22, 10, 27) {real, imag} */,
  {32'h3d590d78, 32'h00000000} /* (22, 10, 26) {real, imag} */,
  {32'hbe0b2613, 32'h00000000} /* (22, 10, 25) {real, imag} */,
  {32'hbe495963, 32'h00000000} /* (22, 10, 24) {real, imag} */,
  {32'hbf04c4ee, 32'h00000000} /* (22, 10, 23) {real, imag} */,
  {32'hbecbb697, 32'h00000000} /* (22, 10, 22) {real, imag} */,
  {32'hbf78cf4a, 32'h00000000} /* (22, 10, 21) {real, imag} */,
  {32'h3db7fff1, 32'h00000000} /* (22, 10, 20) {real, imag} */,
  {32'h3f1fd0eb, 32'h00000000} /* (22, 10, 19) {real, imag} */,
  {32'h3ef5434f, 32'h00000000} /* (22, 10, 18) {real, imag} */,
  {32'h3eeb2c70, 32'h00000000} /* (22, 10, 17) {real, imag} */,
  {32'h3edc9760, 32'h00000000} /* (22, 10, 16) {real, imag} */,
  {32'hbbf280f0, 32'h00000000} /* (22, 10, 15) {real, imag} */,
  {32'hbd7ba555, 32'h00000000} /* (22, 10, 14) {real, imag} */,
  {32'h3e25732d, 32'h00000000} /* (22, 10, 13) {real, imag} */,
  {32'h3eb73a67, 32'h00000000} /* (22, 10, 12) {real, imag} */,
  {32'h3ef8de4e, 32'h00000000} /* (22, 10, 11) {real, imag} */,
  {32'h3dee6c81, 32'h00000000} /* (22, 10, 10) {real, imag} */,
  {32'hbe85e81c, 32'h00000000} /* (22, 10, 9) {real, imag} */,
  {32'h3ec663c9, 32'h00000000} /* (22, 10, 8) {real, imag} */,
  {32'h3e229f92, 32'h00000000} /* (22, 10, 7) {real, imag} */,
  {32'hbec74bbe, 32'h00000000} /* (22, 10, 6) {real, imag} */,
  {32'hbeab9596, 32'h00000000} /* (22, 10, 5) {real, imag} */,
  {32'hbf171cb4, 32'h00000000} /* (22, 10, 4) {real, imag} */,
  {32'hbf12bc3c, 32'h00000000} /* (22, 10, 3) {real, imag} */,
  {32'hbe61de18, 32'h00000000} /* (22, 10, 2) {real, imag} */,
  {32'hbd2d3c63, 32'h00000000} /* (22, 10, 1) {real, imag} */,
  {32'hbd318d18, 32'h00000000} /* (22, 10, 0) {real, imag} */,
  {32'hbf1172fd, 32'h00000000} /* (22, 9, 31) {real, imag} */,
  {32'hbf9428a7, 32'h00000000} /* (22, 9, 30) {real, imag} */,
  {32'hbf9fbeea, 32'h00000000} /* (22, 9, 29) {real, imag} */,
  {32'hbf40293a, 32'h00000000} /* (22, 9, 28) {real, imag} */,
  {32'hbf33050d, 32'h00000000} /* (22, 9, 27) {real, imag} */,
  {32'hbf09a1c4, 32'h00000000} /* (22, 9, 26) {real, imag} */,
  {32'hbed0104d, 32'h00000000} /* (22, 9, 25) {real, imag} */,
  {32'hbf41279c, 32'h00000000} /* (22, 9, 24) {real, imag} */,
  {32'hbf66a8bf, 32'h00000000} /* (22, 9, 23) {real, imag} */,
  {32'hbf3bd571, 32'h00000000} /* (22, 9, 22) {real, imag} */,
  {32'hbf748a12, 32'h00000000} /* (22, 9, 21) {real, imag} */,
  {32'h3eaa1621, 32'h00000000} /* (22, 9, 20) {real, imag} */,
  {32'h3f3accd8, 32'h00000000} /* (22, 9, 19) {real, imag} */,
  {32'h3f91e97f, 32'h00000000} /* (22, 9, 18) {real, imag} */,
  {32'h3f802b42, 32'h00000000} /* (22, 9, 17) {real, imag} */,
  {32'h3f707686, 32'h00000000} /* (22, 9, 16) {real, imag} */,
  {32'h3f33e0ff, 32'h00000000} /* (22, 9, 15) {real, imag} */,
  {32'h3f023473, 32'h00000000} /* (22, 9, 14) {real, imag} */,
  {32'h3f4f53f6, 32'h00000000} /* (22, 9, 13) {real, imag} */,
  {32'h3f63a0a3, 32'h00000000} /* (22, 9, 12) {real, imag} */,
  {32'h3f6a5512, 32'h00000000} /* (22, 9, 11) {real, imag} */,
  {32'hbc256398, 32'h00000000} /* (22, 9, 10) {real, imag} */,
  {32'hbf2eddb1, 32'h00000000} /* (22, 9, 9) {real, imag} */,
  {32'hbf2888d1, 32'h00000000} /* (22, 9, 8) {real, imag} */,
  {32'hbf7ef4bf, 32'h00000000} /* (22, 9, 7) {real, imag} */,
  {32'hbf87316d, 32'h00000000} /* (22, 9, 6) {real, imag} */,
  {32'hbf48671a, 32'h00000000} /* (22, 9, 5) {real, imag} */,
  {32'hbfaa1db0, 32'h00000000} /* (22, 9, 4) {real, imag} */,
  {32'hbfba47fa, 32'h00000000} /* (22, 9, 3) {real, imag} */,
  {32'hbf70841a, 32'h00000000} /* (22, 9, 2) {real, imag} */,
  {32'hbf8a1060, 32'h00000000} /* (22, 9, 1) {real, imag} */,
  {32'hbf2b7076, 32'h00000000} /* (22, 9, 0) {real, imag} */,
  {32'hbee094fe, 32'h00000000} /* (22, 8, 31) {real, imag} */,
  {32'hbf92b994, 32'h00000000} /* (22, 8, 30) {real, imag} */,
  {32'hbf891ef6, 32'h00000000} /* (22, 8, 29) {real, imag} */,
  {32'hbf3ce0bb, 32'h00000000} /* (22, 8, 28) {real, imag} */,
  {32'hbf2745fd, 32'h00000000} /* (22, 8, 27) {real, imag} */,
  {32'hbf6046a8, 32'h00000000} /* (22, 8, 26) {real, imag} */,
  {32'hbf8340a1, 32'h00000000} /* (22, 8, 25) {real, imag} */,
  {32'hbfc5b572, 32'h00000000} /* (22, 8, 24) {real, imag} */,
  {32'hbfab095e, 32'h00000000} /* (22, 8, 23) {real, imag} */,
  {32'hbf576f6f, 32'h00000000} /* (22, 8, 22) {real, imag} */,
  {32'hbf333e08, 32'h00000000} /* (22, 8, 21) {real, imag} */,
  {32'h3ef68a75, 32'h00000000} /* (22, 8, 20) {real, imag} */,
  {32'h3f4cf923, 32'h00000000} /* (22, 8, 19) {real, imag} */,
  {32'h3f9e80cb, 32'h00000000} /* (22, 8, 18) {real, imag} */,
  {32'h3f980795, 32'h00000000} /* (22, 8, 17) {real, imag} */,
  {32'h3eeadb58, 32'h00000000} /* (22, 8, 16) {real, imag} */,
  {32'h3f459085, 32'h00000000} /* (22, 8, 15) {real, imag} */,
  {32'h3f87db93, 32'h00000000} /* (22, 8, 14) {real, imag} */,
  {32'h3f464e63, 32'h00000000} /* (22, 8, 13) {real, imag} */,
  {32'h3f4d3568, 32'h00000000} /* (22, 8, 12) {real, imag} */,
  {32'h3f3efe84, 32'h00000000} /* (22, 8, 11) {real, imag} */,
  {32'hbd8669db, 32'h00000000} /* (22, 8, 10) {real, imag} */,
  {32'hbf525e0e, 32'h00000000} /* (22, 8, 9) {real, imag} */,
  {32'hbf7f5e50, 32'h00000000} /* (22, 8, 8) {real, imag} */,
  {32'hbf535169, 32'h00000000} /* (22, 8, 7) {real, imag} */,
  {32'hbf60b1ac, 32'h00000000} /* (22, 8, 6) {real, imag} */,
  {32'hbf7eed4a, 32'h00000000} /* (22, 8, 5) {real, imag} */,
  {32'hbf827c3e, 32'h00000000} /* (22, 8, 4) {real, imag} */,
  {32'hbf6ed93b, 32'h00000000} /* (22, 8, 3) {real, imag} */,
  {32'hbf8e6ff4, 32'h00000000} /* (22, 8, 2) {real, imag} */,
  {32'hbf54bd49, 32'h00000000} /* (22, 8, 1) {real, imag} */,
  {32'h3c87ef38, 32'h00000000} /* (22, 8, 0) {real, imag} */,
  {32'hbebb66f3, 32'h00000000} /* (22, 7, 31) {real, imag} */,
  {32'hbf883111, 32'h00000000} /* (22, 7, 30) {real, imag} */,
  {32'hbf7bc699, 32'h00000000} /* (22, 7, 29) {real, imag} */,
  {32'hbf56ba51, 32'h00000000} /* (22, 7, 28) {real, imag} */,
  {32'hbf3735bd, 32'h00000000} /* (22, 7, 27) {real, imag} */,
  {32'hbf88d5bd, 32'h00000000} /* (22, 7, 26) {real, imag} */,
  {32'hbfd115c1, 32'h00000000} /* (22, 7, 25) {real, imag} */,
  {32'hbf951772, 32'h00000000} /* (22, 7, 24) {real, imag} */,
  {32'hbf9095d1, 32'h00000000} /* (22, 7, 23) {real, imag} */,
  {32'hbf836b47, 32'h00000000} /* (22, 7, 22) {real, imag} */,
  {32'hbf1f9cdc, 32'h00000000} /* (22, 7, 21) {real, imag} */,
  {32'h3f16605f, 32'h00000000} /* (22, 7, 20) {real, imag} */,
  {32'h3f5f9cd5, 32'h00000000} /* (22, 7, 19) {real, imag} */,
  {32'h3f4a5b5c, 32'h00000000} /* (22, 7, 18) {real, imag} */,
  {32'h3f83f718, 32'h00000000} /* (22, 7, 17) {real, imag} */,
  {32'h3f15a8dd, 32'h00000000} /* (22, 7, 16) {real, imag} */,
  {32'h3f1ca3ae, 32'h00000000} /* (22, 7, 15) {real, imag} */,
  {32'h3f6a0d5b, 32'h00000000} /* (22, 7, 14) {real, imag} */,
  {32'h3f5adbdf, 32'h00000000} /* (22, 7, 13) {real, imag} */,
  {32'h3f34f136, 32'h00000000} /* (22, 7, 12) {real, imag} */,
  {32'h3efa123a, 32'h00000000} /* (22, 7, 11) {real, imag} */,
  {32'hbe96fbf2, 32'h00000000} /* (22, 7, 10) {real, imag} */,
  {32'hbf11e5c4, 32'h00000000} /* (22, 7, 9) {real, imag} */,
  {32'hbf3db599, 32'h00000000} /* (22, 7, 8) {real, imag} */,
  {32'hbee96a44, 32'h00000000} /* (22, 7, 7) {real, imag} */,
  {32'hbf841b1a, 32'h00000000} /* (22, 7, 6) {real, imag} */,
  {32'hbfbee91e, 32'h00000000} /* (22, 7, 5) {real, imag} */,
  {32'hbf594f43, 32'h00000000} /* (22, 7, 4) {real, imag} */,
  {32'hbf74ebe8, 32'h00000000} /* (22, 7, 3) {real, imag} */,
  {32'hbfb64787, 32'h00000000} /* (22, 7, 2) {real, imag} */,
  {32'hbf35853c, 32'h00000000} /* (22, 7, 1) {real, imag} */,
  {32'hbdc4998f, 32'h00000000} /* (22, 7, 0) {real, imag} */,
  {32'hbe9d14d3, 32'h00000000} /* (22, 6, 31) {real, imag} */,
  {32'hbefd1af5, 32'h00000000} /* (22, 6, 30) {real, imag} */,
  {32'hbf1c0e8b, 32'h00000000} /* (22, 6, 29) {real, imag} */,
  {32'hbf7c9596, 32'h00000000} /* (22, 6, 28) {real, imag} */,
  {32'hbf7f105e, 32'h00000000} /* (22, 6, 27) {real, imag} */,
  {32'hbf82613e, 32'h00000000} /* (22, 6, 26) {real, imag} */,
  {32'hbf923208, 32'h00000000} /* (22, 6, 25) {real, imag} */,
  {32'hbf0b65be, 32'h00000000} /* (22, 6, 24) {real, imag} */,
  {32'hbf20d339, 32'h00000000} /* (22, 6, 23) {real, imag} */,
  {32'hbf6a6b3d, 32'h00000000} /* (22, 6, 22) {real, imag} */,
  {32'hbf032cc1, 32'h00000000} /* (22, 6, 21) {real, imag} */,
  {32'h3f0ee4f6, 32'h00000000} /* (22, 6, 20) {real, imag} */,
  {32'h3f118fdd, 32'h00000000} /* (22, 6, 19) {real, imag} */,
  {32'h3f19e23b, 32'h00000000} /* (22, 6, 18) {real, imag} */,
  {32'h3f3a8cf1, 32'h00000000} /* (22, 6, 17) {real, imag} */,
  {32'h3f2c0dee, 32'h00000000} /* (22, 6, 16) {real, imag} */,
  {32'h3f9033fe, 32'h00000000} /* (22, 6, 15) {real, imag} */,
  {32'h3f6fecb2, 32'h00000000} /* (22, 6, 14) {real, imag} */,
  {32'h3f807f3f, 32'h00000000} /* (22, 6, 13) {real, imag} */,
  {32'h3f6404a1, 32'h00000000} /* (22, 6, 12) {real, imag} */,
  {32'h3f1973ae, 32'h00000000} /* (22, 6, 11) {real, imag} */,
  {32'hbe51ba36, 32'h00000000} /* (22, 6, 10) {real, imag} */,
  {32'hbf50aaf1, 32'h00000000} /* (22, 6, 9) {real, imag} */,
  {32'hbf326f3e, 32'h00000000} /* (22, 6, 8) {real, imag} */,
  {32'hbe907966, 32'h00000000} /* (22, 6, 7) {real, imag} */,
  {32'hbf7eddbf, 32'h00000000} /* (22, 6, 6) {real, imag} */,
  {32'hbf2d382a, 32'h00000000} /* (22, 6, 5) {real, imag} */,
  {32'hbeea9a46, 32'h00000000} /* (22, 6, 4) {real, imag} */,
  {32'hbf568e39, 32'h00000000} /* (22, 6, 3) {real, imag} */,
  {32'hbf43998c, 32'h00000000} /* (22, 6, 2) {real, imag} */,
  {32'hbf1e9295, 32'h00000000} /* (22, 6, 1) {real, imag} */,
  {32'hbf07ec9d, 32'h00000000} /* (22, 6, 0) {real, imag} */,
  {32'hbf12f46d, 32'h00000000} /* (22, 5, 31) {real, imag} */,
  {32'hbf9c84e7, 32'h00000000} /* (22, 5, 30) {real, imag} */,
  {32'hbf88d3c3, 32'h00000000} /* (22, 5, 29) {real, imag} */,
  {32'hbf9a0893, 32'h00000000} /* (22, 5, 28) {real, imag} */,
  {32'hbfaae353, 32'h00000000} /* (22, 5, 27) {real, imag} */,
  {32'hbf95b226, 32'h00000000} /* (22, 5, 26) {real, imag} */,
  {32'hbf972854, 32'h00000000} /* (22, 5, 25) {real, imag} */,
  {32'hbf806cdc, 32'h00000000} /* (22, 5, 24) {real, imag} */,
  {32'hbf21efb0, 32'h00000000} /* (22, 5, 23) {real, imag} */,
  {32'hbf454fc9, 32'h00000000} /* (22, 5, 22) {real, imag} */,
  {32'hbf3d8481, 32'h00000000} /* (22, 5, 21) {real, imag} */,
  {32'hbed939fd, 32'h00000000} /* (22, 5, 20) {real, imag} */,
  {32'hbe81bd54, 32'h00000000} /* (22, 5, 19) {real, imag} */,
  {32'hbdb37588, 32'h00000000} /* (22, 5, 18) {real, imag} */,
  {32'hbeadcab9, 32'h00000000} /* (22, 5, 17) {real, imag} */,
  {32'hbf1f3c9a, 32'h00000000} /* (22, 5, 16) {real, imag} */,
  {32'h3f035108, 32'h00000000} /* (22, 5, 15) {real, imag} */,
  {32'h3f86c2da, 32'h00000000} /* (22, 5, 14) {real, imag} */,
  {32'h3f4b7752, 32'h00000000} /* (22, 5, 13) {real, imag} */,
  {32'h3f0f9af9, 32'h00000000} /* (22, 5, 12) {real, imag} */,
  {32'h3f8d6581, 32'h00000000} /* (22, 5, 11) {real, imag} */,
  {32'h3f861b50, 32'h00000000} /* (22, 5, 10) {real, imag} */,
  {32'h3e179d60, 32'h00000000} /* (22, 5, 9) {real, imag} */,
  {32'h3f1caa07, 32'h00000000} /* (22, 5, 8) {real, imag} */,
  {32'h3f57377d, 32'h00000000} /* (22, 5, 7) {real, imag} */,
  {32'h3ef62d0e, 32'h00000000} /* (22, 5, 6) {real, imag} */,
  {32'hbea2b6c9, 32'h00000000} /* (22, 5, 5) {real, imag} */,
  {32'hbf1cf188, 32'h00000000} /* (22, 5, 4) {real, imag} */,
  {32'hbfa4b7a6, 32'h00000000} /* (22, 5, 3) {real, imag} */,
  {32'hbf673d62, 32'h00000000} /* (22, 5, 2) {real, imag} */,
  {32'hbee25b9d, 32'h00000000} /* (22, 5, 1) {real, imag} */,
  {32'hbefd432d, 32'h00000000} /* (22, 5, 0) {real, imag} */,
  {32'hbf03387e, 32'h00000000} /* (22, 4, 31) {real, imag} */,
  {32'hbf9650bb, 32'h00000000} /* (22, 4, 30) {real, imag} */,
  {32'hbf952495, 32'h00000000} /* (22, 4, 29) {real, imag} */,
  {32'hbf9ac33d, 32'h00000000} /* (22, 4, 28) {real, imag} */,
  {32'hbfd8e66f, 32'h00000000} /* (22, 4, 27) {real, imag} */,
  {32'hbfb02591, 32'h00000000} /* (22, 4, 26) {real, imag} */,
  {32'hbfa4251b, 32'h00000000} /* (22, 4, 25) {real, imag} */,
  {32'hbfa0ee6d, 32'h00000000} /* (22, 4, 24) {real, imag} */,
  {32'hbf5322fd, 32'h00000000} /* (22, 4, 23) {real, imag} */,
  {32'hbee9646e, 32'h00000000} /* (22, 4, 22) {real, imag} */,
  {32'hbf0ee8af, 32'h00000000} /* (22, 4, 21) {real, imag} */,
  {32'hbf7caec0, 32'h00000000} /* (22, 4, 20) {real, imag} */,
  {32'hbf5c1565, 32'h00000000} /* (22, 4, 19) {real, imag} */,
  {32'hbf004bbe, 32'h00000000} /* (22, 4, 18) {real, imag} */,
  {32'hbf24a039, 32'h00000000} /* (22, 4, 17) {real, imag} */,
  {32'hbf5e79d5, 32'h00000000} /* (22, 4, 16) {real, imag} */,
  {32'h3e8de646, 32'h00000000} /* (22, 4, 15) {real, imag} */,
  {32'h3f7e1929, 32'h00000000} /* (22, 4, 14) {real, imag} */,
  {32'h3f54486d, 32'h00000000} /* (22, 4, 13) {real, imag} */,
  {32'h3f0d532b, 32'h00000000} /* (22, 4, 12) {real, imag} */,
  {32'h3f88bd12, 32'h00000000} /* (22, 4, 11) {real, imag} */,
  {32'h3fade0c1, 32'h00000000} /* (22, 4, 10) {real, imag} */,
  {32'h3fafcf03, 32'h00000000} /* (22, 4, 9) {real, imag} */,
  {32'h3fc6982c, 32'h00000000} /* (22, 4, 8) {real, imag} */,
  {32'h3fa00387, 32'h00000000} /* (22, 4, 7) {real, imag} */,
  {32'h3f8c247f, 32'h00000000} /* (22, 4, 6) {real, imag} */,
  {32'hbe8e1af2, 32'h00000000} /* (22, 4, 5) {real, imag} */,
  {32'hbf610201, 32'h00000000} /* (22, 4, 4) {real, imag} */,
  {32'hbf9828e8, 32'h00000000} /* (22, 4, 3) {real, imag} */,
  {32'hbf71d7de, 32'h00000000} /* (22, 4, 2) {real, imag} */,
  {32'hbefabfdf, 32'h00000000} /* (22, 4, 1) {real, imag} */,
  {32'hbef5e294, 32'h00000000} /* (22, 4, 0) {real, imag} */,
  {32'hbf065682, 32'h00000000} /* (22, 3, 31) {real, imag} */,
  {32'hbfa5edc3, 32'h00000000} /* (22, 3, 30) {real, imag} */,
  {32'hbf9511d9, 32'h00000000} /* (22, 3, 29) {real, imag} */,
  {32'hbfaafbb9, 32'h00000000} /* (22, 3, 28) {real, imag} */,
  {32'hbfd992e8, 32'h00000000} /* (22, 3, 27) {real, imag} */,
  {32'hbf924428, 32'h00000000} /* (22, 3, 26) {real, imag} */,
  {32'hbf98471f, 32'h00000000} /* (22, 3, 25) {real, imag} */,
  {32'hbf627df8, 32'h00000000} /* (22, 3, 24) {real, imag} */,
  {32'hbfb27b57, 32'h00000000} /* (22, 3, 23) {real, imag} */,
  {32'hbf5a86c5, 32'h00000000} /* (22, 3, 22) {real, imag} */,
  {32'hbf40f8c3, 32'h00000000} /* (22, 3, 21) {real, imag} */,
  {32'hbf301de1, 32'h00000000} /* (22, 3, 20) {real, imag} */,
  {32'hbe73078c, 32'h00000000} /* (22, 3, 19) {real, imag} */,
  {32'hbf1e17fe, 32'h00000000} /* (22, 3, 18) {real, imag} */,
  {32'hbf832665, 32'h00000000} /* (22, 3, 17) {real, imag} */,
  {32'hbf2efaa3, 32'h00000000} /* (22, 3, 16) {real, imag} */,
  {32'h3f0444b9, 32'h00000000} /* (22, 3, 15) {real, imag} */,
  {32'h3fba3146, 32'h00000000} /* (22, 3, 14) {real, imag} */,
  {32'h3f87bc5d, 32'h00000000} /* (22, 3, 13) {real, imag} */,
  {32'h3f385cc0, 32'h00000000} /* (22, 3, 12) {real, imag} */,
  {32'h3f9213c3, 32'h00000000} /* (22, 3, 11) {real, imag} */,
  {32'h3fa3c668, 32'h00000000} /* (22, 3, 10) {real, imag} */,
  {32'h3f71c00e, 32'h00000000} /* (22, 3, 9) {real, imag} */,
  {32'h3f732f12, 32'h00000000} /* (22, 3, 8) {real, imag} */,
  {32'h3f95e8ca, 32'h00000000} /* (22, 3, 7) {real, imag} */,
  {32'h3f83636f, 32'h00000000} /* (22, 3, 6) {real, imag} */,
  {32'hbef3bea0, 32'h00000000} /* (22, 3, 5) {real, imag} */,
  {32'hbfac27c3, 32'h00000000} /* (22, 3, 4) {real, imag} */,
  {32'hbfd41404, 32'h00000000} /* (22, 3, 3) {real, imag} */,
  {32'hbff68a74, 32'h00000000} /* (22, 3, 2) {real, imag} */,
  {32'hbf955cfd, 32'h00000000} /* (22, 3, 1) {real, imag} */,
  {32'hbf04ef78, 32'h00000000} /* (22, 3, 0) {real, imag} */,
  {32'hbf21f0ee, 32'h00000000} /* (22, 2, 31) {real, imag} */,
  {32'hbfabe053, 32'h00000000} /* (22, 2, 30) {real, imag} */,
  {32'hbfc49077, 32'h00000000} /* (22, 2, 29) {real, imag} */,
  {32'hbf811e21, 32'h00000000} /* (22, 2, 28) {real, imag} */,
  {32'hbf45afc2, 32'h00000000} /* (22, 2, 27) {real, imag} */,
  {32'hbf52c6d5, 32'h00000000} /* (22, 2, 26) {real, imag} */,
  {32'hbf7c1ab4, 32'h00000000} /* (22, 2, 25) {real, imag} */,
  {32'hbf55a066, 32'h00000000} /* (22, 2, 24) {real, imag} */,
  {32'hbfa671b4, 32'h00000000} /* (22, 2, 23) {real, imag} */,
  {32'hbf571033, 32'h00000000} /* (22, 2, 22) {real, imag} */,
  {32'hbf2f5a03, 32'h00000000} /* (22, 2, 21) {real, imag} */,
  {32'hbf12f7e7, 32'h00000000} /* (22, 2, 20) {real, imag} */,
  {32'hbf0a063b, 32'h00000000} /* (22, 2, 19) {real, imag} */,
  {32'hbf1256b1, 32'h00000000} /* (22, 2, 18) {real, imag} */,
  {32'hbf5c5c5e, 32'h00000000} /* (22, 2, 17) {real, imag} */,
  {32'hbf33bff3, 32'h00000000} /* (22, 2, 16) {real, imag} */,
  {32'h3e61de45, 32'h00000000} /* (22, 2, 15) {real, imag} */,
  {32'h3fac2418, 32'h00000000} /* (22, 2, 14) {real, imag} */,
  {32'h3f5be346, 32'h00000000} /* (22, 2, 13) {real, imag} */,
  {32'h3ef0a87a, 32'h00000000} /* (22, 2, 12) {real, imag} */,
  {32'h3f26d786, 32'h00000000} /* (22, 2, 11) {real, imag} */,
  {32'h3ef9b552, 32'h00000000} /* (22, 2, 10) {real, imag} */,
  {32'h3f46bc66, 32'h00000000} /* (22, 2, 9) {real, imag} */,
  {32'h3f81bf41, 32'h00000000} /* (22, 2, 8) {real, imag} */,
  {32'h3f4e6e8f, 32'h00000000} /* (22, 2, 7) {real, imag} */,
  {32'h3f5a723e, 32'h00000000} /* (22, 2, 6) {real, imag} */,
  {32'hbde25c28, 32'h00000000} /* (22, 2, 5) {real, imag} */,
  {32'hbf3bdf65, 32'h00000000} /* (22, 2, 4) {real, imag} */,
  {32'hbf7f1916, 32'h00000000} /* (22, 2, 3) {real, imag} */,
  {32'hbff36863, 32'h00000000} /* (22, 2, 2) {real, imag} */,
  {32'hbfbb8e29, 32'h00000000} /* (22, 2, 1) {real, imag} */,
  {32'hbed2a07a, 32'h00000000} /* (22, 2, 0) {real, imag} */,
  {32'hbea13db1, 32'h00000000} /* (22, 1, 31) {real, imag} */,
  {32'hbf1423e9, 32'h00000000} /* (22, 1, 30) {real, imag} */,
  {32'hbf5dcbc8, 32'h00000000} /* (22, 1, 29) {real, imag} */,
  {32'hbf0e3275, 32'h00000000} /* (22, 1, 28) {real, imag} */,
  {32'hbf255a6f, 32'h00000000} /* (22, 1, 27) {real, imag} */,
  {32'hbfad5153, 32'h00000000} /* (22, 1, 26) {real, imag} */,
  {32'hbf9ee515, 32'h00000000} /* (22, 1, 25) {real, imag} */,
  {32'hbf50bcae, 32'h00000000} /* (22, 1, 24) {real, imag} */,
  {32'hbf897364, 32'h00000000} /* (22, 1, 23) {real, imag} */,
  {32'hbf6243eb, 32'h00000000} /* (22, 1, 22) {real, imag} */,
  {32'hbeff0476, 32'h00000000} /* (22, 1, 21) {real, imag} */,
  {32'hbf450a93, 32'h00000000} /* (22, 1, 20) {real, imag} */,
  {32'hbf31337c, 32'h00000000} /* (22, 1, 19) {real, imag} */,
  {32'hbf368963, 32'h00000000} /* (22, 1, 18) {real, imag} */,
  {32'hbfa9674c, 32'h00000000} /* (22, 1, 17) {real, imag} */,
  {32'hbf70f718, 32'h00000000} /* (22, 1, 16) {real, imag} */,
  {32'h3e43d007, 32'h00000000} /* (22, 1, 15) {real, imag} */,
  {32'h3f998ad7, 32'h00000000} /* (22, 1, 14) {real, imag} */,
  {32'h3f5e9f98, 32'h00000000} /* (22, 1, 13) {real, imag} */,
  {32'h3f2dd02d, 32'h00000000} /* (22, 1, 12) {real, imag} */,
  {32'h3f0ba38b, 32'h00000000} /* (22, 1, 11) {real, imag} */,
  {32'h3ee7df7f, 32'h00000000} /* (22, 1, 10) {real, imag} */,
  {32'h3f6c54f2, 32'h00000000} /* (22, 1, 9) {real, imag} */,
  {32'h3fb03897, 32'h00000000} /* (22, 1, 8) {real, imag} */,
  {32'h3f661756, 32'h00000000} /* (22, 1, 7) {real, imag} */,
  {32'h3f49e1f8, 32'h00000000} /* (22, 1, 6) {real, imag} */,
  {32'h3d930cc8, 32'h00000000} /* (22, 1, 5) {real, imag} */,
  {32'hbf0bacf3, 32'h00000000} /* (22, 1, 4) {real, imag} */,
  {32'hbf580341, 32'h00000000} /* (22, 1, 3) {real, imag} */,
  {32'hbf97bf28, 32'h00000000} /* (22, 1, 2) {real, imag} */,
  {32'hbf5cbe86, 32'h00000000} /* (22, 1, 1) {real, imag} */,
  {32'hbeb95827, 32'h00000000} /* (22, 1, 0) {real, imag} */,
  {32'hbddf910b, 32'h00000000} /* (22, 0, 31) {real, imag} */,
  {32'hbe881640, 32'h00000000} /* (22, 0, 30) {real, imag} */,
  {32'hbe91ee15, 32'h00000000} /* (22, 0, 29) {real, imag} */,
  {32'hbdf9d92d, 32'h00000000} /* (22, 0, 28) {real, imag} */,
  {32'hbf203417, 32'h00000000} /* (22, 0, 27) {real, imag} */,
  {32'hbfbe3ba7, 32'h00000000} /* (22, 0, 26) {real, imag} */,
  {32'hbf341ebc, 32'h00000000} /* (22, 0, 25) {real, imag} */,
  {32'hbe3a41c3, 32'h00000000} /* (22, 0, 24) {real, imag} */,
  {32'hbeb6a2f4, 32'h00000000} /* (22, 0, 23) {real, imag} */,
  {32'hbec3dabf, 32'h00000000} /* (22, 0, 22) {real, imag} */,
  {32'hbd20c822, 32'h00000000} /* (22, 0, 21) {real, imag} */,
  {32'hbf376f4b, 32'h00000000} /* (22, 0, 20) {real, imag} */,
  {32'hbeb28d50, 32'h00000000} /* (22, 0, 19) {real, imag} */,
  {32'hbe9c1263, 32'h00000000} /* (22, 0, 18) {real, imag} */,
  {32'hbf4de59e, 32'h00000000} /* (22, 0, 17) {real, imag} */,
  {32'hbed87113, 32'h00000000} /* (22, 0, 16) {real, imag} */,
  {32'h3e8e6b2e, 32'h00000000} /* (22, 0, 15) {real, imag} */,
  {32'h3f338069, 32'h00000000} /* (22, 0, 14) {real, imag} */,
  {32'h3ee4e988, 32'h00000000} /* (22, 0, 13) {real, imag} */,
  {32'h3f0aebea, 32'h00000000} /* (22, 0, 12) {real, imag} */,
  {32'h3f0d66ac, 32'h00000000} /* (22, 0, 11) {real, imag} */,
  {32'h3ea64d3b, 32'h00000000} /* (22, 0, 10) {real, imag} */,
  {32'h3eb931f7, 32'h00000000} /* (22, 0, 9) {real, imag} */,
  {32'h3efa6976, 32'h00000000} /* (22, 0, 8) {real, imag} */,
  {32'h3e90759b, 32'h00000000} /* (22, 0, 7) {real, imag} */,
  {32'h3e4403e8, 32'h00000000} /* (22, 0, 6) {real, imag} */,
  {32'hba4fe6f8, 32'h00000000} /* (22, 0, 5) {real, imag} */,
  {32'hbe374469, 32'h00000000} /* (22, 0, 4) {real, imag} */,
  {32'hbe54154d, 32'h00000000} /* (22, 0, 3) {real, imag} */,
  {32'hbece258f, 32'h00000000} /* (22, 0, 2) {real, imag} */,
  {32'hbf3e5527, 32'h00000000} /* (22, 0, 1) {real, imag} */,
  {32'hbf018d8a, 32'h00000000} /* (22, 0, 0) {real, imag} */,
  {32'hbea59132, 32'h00000000} /* (21, 31, 31) {real, imag} */,
  {32'hbf0bebc4, 32'h00000000} /* (21, 31, 30) {real, imag} */,
  {32'hbe31fb9b, 32'h00000000} /* (21, 31, 29) {real, imag} */,
  {32'hbeba8300, 32'h00000000} /* (21, 31, 28) {real, imag} */,
  {32'hbee21f64, 32'h00000000} /* (21, 31, 27) {real, imag} */,
  {32'hbeb2dcb1, 32'h00000000} /* (21, 31, 26) {real, imag} */,
  {32'hbedd4ce9, 32'h00000000} /* (21, 31, 25) {real, imag} */,
  {32'hbec84703, 32'h00000000} /* (21, 31, 24) {real, imag} */,
  {32'hbe917d51, 32'h00000000} /* (21, 31, 23) {real, imag} */,
  {32'hbee08218, 32'h00000000} /* (21, 31, 22) {real, imag} */,
  {32'hbe773e78, 32'h00000000} /* (21, 31, 21) {real, imag} */,
  {32'h3c5c455c, 32'h00000000} /* (21, 31, 20) {real, imag} */,
  {32'h3e9f249e, 32'h00000000} /* (21, 31, 19) {real, imag} */,
  {32'h3e87a2b5, 32'h00000000} /* (21, 31, 18) {real, imag} */,
  {32'hbd19ac8b, 32'h00000000} /* (21, 31, 17) {real, imag} */,
  {32'h3ee233fe, 32'h00000000} /* (21, 31, 16) {real, imag} */,
  {32'h3f2451c5, 32'h00000000} /* (21, 31, 15) {real, imag} */,
  {32'h3f3085de, 32'h00000000} /* (21, 31, 14) {real, imag} */,
  {32'h3f33742a, 32'h00000000} /* (21, 31, 13) {real, imag} */,
  {32'h3ea6675e, 32'h00000000} /* (21, 31, 12) {real, imag} */,
  {32'h3e5ea477, 32'h00000000} /* (21, 31, 11) {real, imag} */,
  {32'h3ce103fb, 32'h00000000} /* (21, 31, 10) {real, imag} */,
  {32'hbeb8111a, 32'h00000000} /* (21, 31, 9) {real, imag} */,
  {32'hbedf8035, 32'h00000000} /* (21, 31, 8) {real, imag} */,
  {32'hbf3e81ed, 32'h00000000} /* (21, 31, 7) {real, imag} */,
  {32'hbf076a2d, 32'h00000000} /* (21, 31, 6) {real, imag} */,
  {32'hbe4c4570, 32'h00000000} /* (21, 31, 5) {real, imag} */,
  {32'hbd9ad980, 32'h00000000} /* (21, 31, 4) {real, imag} */,
  {32'hbe0e66cc, 32'h00000000} /* (21, 31, 3) {real, imag} */,
  {32'hbeb940bf, 32'h00000000} /* (21, 31, 2) {real, imag} */,
  {32'hbee08945, 32'h00000000} /* (21, 31, 1) {real, imag} */,
  {32'hbddebf71, 32'h00000000} /* (21, 31, 0) {real, imag} */,
  {32'hbf262422, 32'h00000000} /* (21, 30, 31) {real, imag} */,
  {32'hbf4e5d4d, 32'h00000000} /* (21, 30, 30) {real, imag} */,
  {32'hbefa70f2, 32'h00000000} /* (21, 30, 29) {real, imag} */,
  {32'hbf64f07b, 32'h00000000} /* (21, 30, 28) {real, imag} */,
  {32'hbf12781c, 32'h00000000} /* (21, 30, 27) {real, imag} */,
  {32'hbe73d280, 32'h00000000} /* (21, 30, 26) {real, imag} */,
  {32'hbf378596, 32'h00000000} /* (21, 30, 25) {real, imag} */,
  {32'hbf2b717b, 32'h00000000} /* (21, 30, 24) {real, imag} */,
  {32'hbf3b9afa, 32'h00000000} /* (21, 30, 23) {real, imag} */,
  {32'hbf99ec72, 32'h00000000} /* (21, 30, 22) {real, imag} */,
  {32'hbe87b9bc, 32'h00000000} /* (21, 30, 21) {real, imag} */,
  {32'h3f3eb50d, 32'h00000000} /* (21, 30, 20) {real, imag} */,
  {32'h3f91df0b, 32'h00000000} /* (21, 30, 19) {real, imag} */,
  {32'h3f52741b, 32'h00000000} /* (21, 30, 18) {real, imag} */,
  {32'h3df1d22a, 32'h00000000} /* (21, 30, 17) {real, imag} */,
  {32'h3f22cb3d, 32'h00000000} /* (21, 30, 16) {real, imag} */,
  {32'h3f653d9a, 32'h00000000} /* (21, 30, 15) {real, imag} */,
  {32'h3fb2b17a, 32'h00000000} /* (21, 30, 14) {real, imag} */,
  {32'h3fbbdddd, 32'h00000000} /* (21, 30, 13) {real, imag} */,
  {32'h3f6b3714, 32'h00000000} /* (21, 30, 12) {real, imag} */,
  {32'h3ef60f7e, 32'h00000000} /* (21, 30, 11) {real, imag} */,
  {32'hbdcbb19f, 32'h00000000} /* (21, 30, 10) {real, imag} */,
  {32'hbf144c6c, 32'h00000000} /* (21, 30, 9) {real, imag} */,
  {32'hbf00451a, 32'h00000000} /* (21, 30, 8) {real, imag} */,
  {32'hbf074c15, 32'h00000000} /* (21, 30, 7) {real, imag} */,
  {32'hbf2700af, 32'h00000000} /* (21, 30, 6) {real, imag} */,
  {32'hbef051b0, 32'h00000000} /* (21, 30, 5) {real, imag} */,
  {32'hbe19af09, 32'h00000000} /* (21, 30, 4) {real, imag} */,
  {32'hbe8da803, 32'h00000000} /* (21, 30, 3) {real, imag} */,
  {32'hbf524f27, 32'h00000000} /* (21, 30, 2) {real, imag} */,
  {32'hbf93b065, 32'h00000000} /* (21, 30, 1) {real, imag} */,
  {32'hbed12166, 32'h00000000} /* (21, 30, 0) {real, imag} */,
  {32'hbf6b700c, 32'h00000000} /* (21, 29, 31) {real, imag} */,
  {32'hbfb02ef2, 32'h00000000} /* (21, 29, 30) {real, imag} */,
  {32'hbf143a70, 32'h00000000} /* (21, 29, 29) {real, imag} */,
  {32'hbf4effa6, 32'h00000000} /* (21, 29, 28) {real, imag} */,
  {32'hbf3107dd, 32'h00000000} /* (21, 29, 27) {real, imag} */,
  {32'hbecc39eb, 32'h00000000} /* (21, 29, 26) {real, imag} */,
  {32'hbf7d4421, 32'h00000000} /* (21, 29, 25) {real, imag} */,
  {32'hbf14ed97, 32'h00000000} /* (21, 29, 24) {real, imag} */,
  {32'hbf3da8c7, 32'h00000000} /* (21, 29, 23) {real, imag} */,
  {32'hbf69c9b8, 32'h00000000} /* (21, 29, 22) {real, imag} */,
  {32'h3d4e7b38, 32'h00000000} /* (21, 29, 21) {real, imag} */,
  {32'h3fac81fd, 32'h00000000} /* (21, 29, 20) {real, imag} */,
  {32'h3fe25ae0, 32'h00000000} /* (21, 29, 19) {real, imag} */,
  {32'h3fd7b2b9, 32'h00000000} /* (21, 29, 18) {real, imag} */,
  {32'h3f784d22, 32'h00000000} /* (21, 29, 17) {real, imag} */,
  {32'h3f4db086, 32'h00000000} /* (21, 29, 16) {real, imag} */,
  {32'h3f3f505e, 32'h00000000} /* (21, 29, 15) {real, imag} */,
  {32'h3f5cb3cf, 32'h00000000} /* (21, 29, 14) {real, imag} */,
  {32'h3f8b2688, 32'h00000000} /* (21, 29, 13) {real, imag} */,
  {32'h3fa62bf3, 32'h00000000} /* (21, 29, 12) {real, imag} */,
  {32'h3f3f2ea9, 32'h00000000} /* (21, 29, 11) {real, imag} */,
  {32'hbe001770, 32'h00000000} /* (21, 29, 10) {real, imag} */,
  {32'hbf67d934, 32'h00000000} /* (21, 29, 9) {real, imag} */,
  {32'hbf3b6b07, 32'h00000000} /* (21, 29, 8) {real, imag} */,
  {32'hbee577e4, 32'h00000000} /* (21, 29, 7) {real, imag} */,
  {32'hbef404ef, 32'h00000000} /* (21, 29, 6) {real, imag} */,
  {32'hbee0b58f, 32'h00000000} /* (21, 29, 5) {real, imag} */,
  {32'hbf031209, 32'h00000000} /* (21, 29, 4) {real, imag} */,
  {32'hbef0eaa2, 32'h00000000} /* (21, 29, 3) {real, imag} */,
  {32'hbf4c2107, 32'h00000000} /* (21, 29, 2) {real, imag} */,
  {32'hbf922443, 32'h00000000} /* (21, 29, 1) {real, imag} */,
  {32'hbefa8c3a, 32'h00000000} /* (21, 29, 0) {real, imag} */,
  {32'hbf15b7c8, 32'h00000000} /* (21, 28, 31) {real, imag} */,
  {32'hbf6d1eb5, 32'h00000000} /* (21, 28, 30) {real, imag} */,
  {32'hbf1a2e5b, 32'h00000000} /* (21, 28, 29) {real, imag} */,
  {32'hbf8acfa5, 32'h00000000} /* (21, 28, 28) {real, imag} */,
  {32'hbf8b6f01, 32'h00000000} /* (21, 28, 27) {real, imag} */,
  {32'hbf07c6f7, 32'h00000000} /* (21, 28, 26) {real, imag} */,
  {32'hbf8a57c1, 32'h00000000} /* (21, 28, 25) {real, imag} */,
  {32'hbf632251, 32'h00000000} /* (21, 28, 24) {real, imag} */,
  {32'hbf9f749f, 32'h00000000} /* (21, 28, 23) {real, imag} */,
  {32'hbfb6e6cf, 32'h00000000} /* (21, 28, 22) {real, imag} */,
  {32'hbf3018ce, 32'h00000000} /* (21, 28, 21) {real, imag} */,
  {32'h3f0de996, 32'h00000000} /* (21, 28, 20) {real, imag} */,
  {32'h3fad0732, 32'h00000000} /* (21, 28, 19) {real, imag} */,
  {32'h3fb82533, 32'h00000000} /* (21, 28, 18) {real, imag} */,
  {32'h3f7aeb16, 32'h00000000} /* (21, 28, 17) {real, imag} */,
  {32'h3f70713d, 32'h00000000} /* (21, 28, 16) {real, imag} */,
  {32'h3f93ce5e, 32'h00000000} /* (21, 28, 15) {real, imag} */,
  {32'h3f5f8b79, 32'h00000000} /* (21, 28, 14) {real, imag} */,
  {32'h3f1c4d82, 32'h00000000} /* (21, 28, 13) {real, imag} */,
  {32'h3fb8c1b8, 32'h00000000} /* (21, 28, 12) {real, imag} */,
  {32'h3f896124, 32'h00000000} /* (21, 28, 11) {real, imag} */,
  {32'hbe84e39b, 32'h00000000} /* (21, 28, 10) {real, imag} */,
  {32'hbfb23ac2, 32'h00000000} /* (21, 28, 9) {real, imag} */,
  {32'hbfa0559f, 32'h00000000} /* (21, 28, 8) {real, imag} */,
  {32'hbf85dfff, 32'h00000000} /* (21, 28, 7) {real, imag} */,
  {32'hbf8801ad, 32'h00000000} /* (21, 28, 6) {real, imag} */,
  {32'hbf866c45, 32'h00000000} /* (21, 28, 5) {real, imag} */,
  {32'hbf93ad56, 32'h00000000} /* (21, 28, 4) {real, imag} */,
  {32'hbf5fc91b, 32'h00000000} /* (21, 28, 3) {real, imag} */,
  {32'hbf3ba045, 32'h00000000} /* (21, 28, 2) {real, imag} */,
  {32'hbf82b8ed, 32'h00000000} /* (21, 28, 1) {real, imag} */,
  {32'hbf7181eb, 32'h00000000} /* (21, 28, 0) {real, imag} */,
  {32'hbef4f3e0, 32'h00000000} /* (21, 27, 31) {real, imag} */,
  {32'hbf33b4a6, 32'h00000000} /* (21, 27, 30) {real, imag} */,
  {32'hbf5c20df, 32'h00000000} /* (21, 27, 29) {real, imag} */,
  {32'hbfb66f14, 32'h00000000} /* (21, 27, 28) {real, imag} */,
  {32'hbfc3bc15, 32'h00000000} /* (21, 27, 27) {real, imag} */,
  {32'hbf4f0974, 32'h00000000} /* (21, 27, 26) {real, imag} */,
  {32'hbf14a5ae, 32'h00000000} /* (21, 27, 25) {real, imag} */,
  {32'hbfaa103e, 32'h00000000} /* (21, 27, 24) {real, imag} */,
  {32'hbfbdc3f1, 32'h00000000} /* (21, 27, 23) {real, imag} */,
  {32'hbfab29ad, 32'h00000000} /* (21, 27, 22) {real, imag} */,
  {32'hbf1ae971, 32'h00000000} /* (21, 27, 21) {real, imag} */,
  {32'h3e3b2f2f, 32'h00000000} /* (21, 27, 20) {real, imag} */,
  {32'h3f0b70d9, 32'h00000000} /* (21, 27, 19) {real, imag} */,
  {32'h3f2e5e12, 32'h00000000} /* (21, 27, 18) {real, imag} */,
  {32'h3f389061, 32'h00000000} /* (21, 27, 17) {real, imag} */,
  {32'h3f1243b2, 32'h00000000} /* (21, 27, 16) {real, imag} */,
  {32'h3f8444a6, 32'h00000000} /* (21, 27, 15) {real, imag} */,
  {32'h3f6a7a33, 32'h00000000} /* (21, 27, 14) {real, imag} */,
  {32'h3f4c2e3e, 32'h00000000} /* (21, 27, 13) {real, imag} */,
  {32'h3f7a726e, 32'h00000000} /* (21, 27, 12) {real, imag} */,
  {32'h3f3debe9, 32'h00000000} /* (21, 27, 11) {real, imag} */,
  {32'hbeeb8f8e, 32'h00000000} /* (21, 27, 10) {real, imag} */,
  {32'hbf9ae54f, 32'h00000000} /* (21, 27, 9) {real, imag} */,
  {32'hbfb910ba, 32'h00000000} /* (21, 27, 8) {real, imag} */,
  {32'hbf979a0d, 32'h00000000} /* (21, 27, 7) {real, imag} */,
  {32'hbfb993c9, 32'h00000000} /* (21, 27, 6) {real, imag} */,
  {32'hbfb6b8be, 32'h00000000} /* (21, 27, 5) {real, imag} */,
  {32'hbf8fef87, 32'h00000000} /* (21, 27, 4) {real, imag} */,
  {32'hbf768718, 32'h00000000} /* (21, 27, 3) {real, imag} */,
  {32'hbfb35908, 32'h00000000} /* (21, 27, 2) {real, imag} */,
  {32'hbfa7852c, 32'h00000000} /* (21, 27, 1) {real, imag} */,
  {32'hbf77bafd, 32'h00000000} /* (21, 27, 0) {real, imag} */,
  {32'hbeaef8e8, 32'h00000000} /* (21, 26, 31) {real, imag} */,
  {32'hbf8451c5, 32'h00000000} /* (21, 26, 30) {real, imag} */,
  {32'hbf61c159, 32'h00000000} /* (21, 26, 29) {real, imag} */,
  {32'hbf6b0a55, 32'h00000000} /* (21, 26, 28) {real, imag} */,
  {32'hbfc65e44, 32'h00000000} /* (21, 26, 27) {real, imag} */,
  {32'hbf8a161a, 32'h00000000} /* (21, 26, 26) {real, imag} */,
  {32'hbf67f04d, 32'h00000000} /* (21, 26, 25) {real, imag} */,
  {32'hc004418e, 32'h00000000} /* (21, 26, 24) {real, imag} */,
  {32'hbfba4c68, 32'h00000000} /* (21, 26, 23) {real, imag} */,
  {32'hbf6e9abe, 32'h00000000} /* (21, 26, 22) {real, imag} */,
  {32'hbf10e242, 32'h00000000} /* (21, 26, 21) {real, imag} */,
  {32'h3e881ae9, 32'h00000000} /* (21, 26, 20) {real, imag} */,
  {32'h3f75ee95, 32'h00000000} /* (21, 26, 19) {real, imag} */,
  {32'h3f6778d9, 32'h00000000} /* (21, 26, 18) {real, imag} */,
  {32'h3f65e408, 32'h00000000} /* (21, 26, 17) {real, imag} */,
  {32'h3f3e78a3, 32'h00000000} /* (21, 26, 16) {real, imag} */,
  {32'h3f398e54, 32'h00000000} /* (21, 26, 15) {real, imag} */,
  {32'h3f7f865a, 32'h00000000} /* (21, 26, 14) {real, imag} */,
  {32'h3fa85eb1, 32'h00000000} /* (21, 26, 13) {real, imag} */,
  {32'h3fad0658, 32'h00000000} /* (21, 26, 12) {real, imag} */,
  {32'h3f427a62, 32'h00000000} /* (21, 26, 11) {real, imag} */,
  {32'hbf78b9f5, 32'h00000000} /* (21, 26, 10) {real, imag} */,
  {32'hbfd011b7, 32'h00000000} /* (21, 26, 9) {real, imag} */,
  {32'hbf9a500b, 32'h00000000} /* (21, 26, 8) {real, imag} */,
  {32'hbf8cd5ec, 32'h00000000} /* (21, 26, 7) {real, imag} */,
  {32'hbf8afa7f, 32'h00000000} /* (21, 26, 6) {real, imag} */,
  {32'hbf2cfbc4, 32'h00000000} /* (21, 26, 5) {real, imag} */,
  {32'hbf4be7b8, 32'h00000000} /* (21, 26, 4) {real, imag} */,
  {32'hbf7e3bee, 32'h00000000} /* (21, 26, 3) {real, imag} */,
  {32'hbf9cd453, 32'h00000000} /* (21, 26, 2) {real, imag} */,
  {32'hbf9cf1d2, 32'h00000000} /* (21, 26, 1) {real, imag} */,
  {32'hbf25ed46, 32'h00000000} /* (21, 26, 0) {real, imag} */,
  {32'hbef83f83, 32'h00000000} /* (21, 25, 31) {real, imag} */,
  {32'hbf2bc83b, 32'h00000000} /* (21, 25, 30) {real, imag} */,
  {32'hbf427a04, 32'h00000000} /* (21, 25, 29) {real, imag} */,
  {32'hbf77fca2, 32'h00000000} /* (21, 25, 28) {real, imag} */,
  {32'hbfc3aae4, 32'h00000000} /* (21, 25, 27) {real, imag} */,
  {32'hbfacf95a, 32'h00000000} /* (21, 25, 26) {real, imag} */,
  {32'hbf52f9b9, 32'h00000000} /* (21, 25, 25) {real, imag} */,
  {32'hbf9d8b12, 32'h00000000} /* (21, 25, 24) {real, imag} */,
  {32'hbf604b69, 32'h00000000} /* (21, 25, 23) {real, imag} */,
  {32'hbf968649, 32'h00000000} /* (21, 25, 22) {real, imag} */,
  {32'hbf5efdad, 32'h00000000} /* (21, 25, 21) {real, imag} */,
  {32'h3e92b4c8, 32'h00000000} /* (21, 25, 20) {real, imag} */,
  {32'h3f907433, 32'h00000000} /* (21, 25, 19) {real, imag} */,
  {32'h3fb2e208, 32'h00000000} /* (21, 25, 18) {real, imag} */,
  {32'h3f67213b, 32'h00000000} /* (21, 25, 17) {real, imag} */,
  {32'h3f83844b, 32'h00000000} /* (21, 25, 16) {real, imag} */,
  {32'h3f9e44e5, 32'h00000000} /* (21, 25, 15) {real, imag} */,
  {32'h3fbc42f1, 32'h00000000} /* (21, 25, 14) {real, imag} */,
  {32'h3f949ec9, 32'h00000000} /* (21, 25, 13) {real, imag} */,
  {32'h3fa6734e, 32'h00000000} /* (21, 25, 12) {real, imag} */,
  {32'h3f55ffe0, 32'h00000000} /* (21, 25, 11) {real, imag} */,
  {32'hbf678e47, 32'h00000000} /* (21, 25, 10) {real, imag} */,
  {32'hbfbbdfb0, 32'h00000000} /* (21, 25, 9) {real, imag} */,
  {32'hbf857444, 32'h00000000} /* (21, 25, 8) {real, imag} */,
  {32'hbf4488de, 32'h00000000} /* (21, 25, 7) {real, imag} */,
  {32'hbf5a0a4b, 32'h00000000} /* (21, 25, 6) {real, imag} */,
  {32'hbf49f6eb, 32'h00000000} /* (21, 25, 5) {real, imag} */,
  {32'hbf4b69a9, 32'h00000000} /* (21, 25, 4) {real, imag} */,
  {32'hbf81f787, 32'h00000000} /* (21, 25, 3) {real, imag} */,
  {32'hbfb54c60, 32'h00000000} /* (21, 25, 2) {real, imag} */,
  {32'hbf682567, 32'h00000000} /* (21, 25, 1) {real, imag} */,
  {32'hbefb02ed, 32'h00000000} /* (21, 25, 0) {real, imag} */,
  {32'hbe0b7760, 32'h00000000} /* (21, 24, 31) {real, imag} */,
  {32'hbed81e9c, 32'h00000000} /* (21, 24, 30) {real, imag} */,
  {32'hbeda521c, 32'h00000000} /* (21, 24, 29) {real, imag} */,
  {32'hbee29662, 32'h00000000} /* (21, 24, 28) {real, imag} */,
  {32'hbf2c36e3, 32'h00000000} /* (21, 24, 27) {real, imag} */,
  {32'hbf1f3b80, 32'h00000000} /* (21, 24, 26) {real, imag} */,
  {32'hbe7936b1, 32'h00000000} /* (21, 24, 25) {real, imag} */,
  {32'hbf30e0db, 32'h00000000} /* (21, 24, 24) {real, imag} */,
  {32'hbf4f967d, 32'h00000000} /* (21, 24, 23) {real, imag} */,
  {32'hbf8f3fa6, 32'h00000000} /* (21, 24, 22) {real, imag} */,
  {32'hbf2a9238, 32'h00000000} /* (21, 24, 21) {real, imag} */,
  {32'h3f29ecb0, 32'h00000000} /* (21, 24, 20) {real, imag} */,
  {32'h3fb6113b, 32'h00000000} /* (21, 24, 19) {real, imag} */,
  {32'h3fc44474, 32'h00000000} /* (21, 24, 18) {real, imag} */,
  {32'h3f2d354d, 32'h00000000} /* (21, 24, 17) {real, imag} */,
  {32'h3fada589, 32'h00000000} /* (21, 24, 16) {real, imag} */,
  {32'h3fb26635, 32'h00000000} /* (21, 24, 15) {real, imag} */,
  {32'h3f84ad63, 32'h00000000} /* (21, 24, 14) {real, imag} */,
  {32'h3f6bd798, 32'h00000000} /* (21, 24, 13) {real, imag} */,
  {32'h3fa2a44d, 32'h00000000} /* (21, 24, 12) {real, imag} */,
  {32'h3f754b96, 32'h00000000} /* (21, 24, 11) {real, imag} */,
  {32'hbe9a34ba, 32'h00000000} /* (21, 24, 10) {real, imag} */,
  {32'hbf500acf, 32'h00000000} /* (21, 24, 9) {real, imag} */,
  {32'hbf4c9112, 32'h00000000} /* (21, 24, 8) {real, imag} */,
  {32'hbf5bd657, 32'h00000000} /* (21, 24, 7) {real, imag} */,
  {32'hbf9907bd, 32'h00000000} /* (21, 24, 6) {real, imag} */,
  {32'hbf57f855, 32'h00000000} /* (21, 24, 5) {real, imag} */,
  {32'hbf298902, 32'h00000000} /* (21, 24, 4) {real, imag} */,
  {32'hbf724e96, 32'h00000000} /* (21, 24, 3) {real, imag} */,
  {32'hbf99f557, 32'h00000000} /* (21, 24, 2) {real, imag} */,
  {32'hbf43c7f7, 32'h00000000} /* (21, 24, 1) {real, imag} */,
  {32'hbe6a5a0c, 32'h00000000} /* (21, 24, 0) {real, imag} */,
  {32'hbe44dac1, 32'h00000000} /* (21, 23, 31) {real, imag} */,
  {32'hbf63a032, 32'h00000000} /* (21, 23, 30) {real, imag} */,
  {32'hbf8843ee, 32'h00000000} /* (21, 23, 29) {real, imag} */,
  {32'hbf4e4160, 32'h00000000} /* (21, 23, 28) {real, imag} */,
  {32'hbf177562, 32'h00000000} /* (21, 23, 27) {real, imag} */,
  {32'hbf099d8e, 32'h00000000} /* (21, 23, 26) {real, imag} */,
  {32'hbece7ed1, 32'h00000000} /* (21, 23, 25) {real, imag} */,
  {32'hbf339bab, 32'h00000000} /* (21, 23, 24) {real, imag} */,
  {32'hbf8fd042, 32'h00000000} /* (21, 23, 23) {real, imag} */,
  {32'hbf819268, 32'h00000000} /* (21, 23, 22) {real, imag} */,
  {32'hbf057348, 32'h00000000} /* (21, 23, 21) {real, imag} */,
  {32'h3f6cbe9b, 32'h00000000} /* (21, 23, 20) {real, imag} */,
  {32'h3f56b97e, 32'h00000000} /* (21, 23, 19) {real, imag} */,
  {32'h3f322e84, 32'h00000000} /* (21, 23, 18) {real, imag} */,
  {32'h3ef6f958, 32'h00000000} /* (21, 23, 17) {real, imag} */,
  {32'h3f9b21a5, 32'h00000000} /* (21, 23, 16) {real, imag} */,
  {32'h3f629392, 32'h00000000} /* (21, 23, 15) {real, imag} */,
  {32'h3f05fc1e, 32'h00000000} /* (21, 23, 14) {real, imag} */,
  {32'h3f678625, 32'h00000000} /* (21, 23, 13) {real, imag} */,
  {32'h3f8d2690, 32'h00000000} /* (21, 23, 12) {real, imag} */,
  {32'h3f06fa70, 32'h00000000} /* (21, 23, 11) {real, imag} */,
  {32'hbee89e5b, 32'h00000000} /* (21, 23, 10) {real, imag} */,
  {32'hbedc4213, 32'h00000000} /* (21, 23, 9) {real, imag} */,
  {32'hbef24859, 32'h00000000} /* (21, 23, 8) {real, imag} */,
  {32'hbf62f8e4, 32'h00000000} /* (21, 23, 7) {real, imag} */,
  {32'hbf6515b2, 32'h00000000} /* (21, 23, 6) {real, imag} */,
  {32'hbfa1cfb6, 32'h00000000} /* (21, 23, 5) {real, imag} */,
  {32'hbfaf57fe, 32'h00000000} /* (21, 23, 4) {real, imag} */,
  {32'hbfab3722, 32'h00000000} /* (21, 23, 3) {real, imag} */,
  {32'hbf43ce65, 32'h00000000} /* (21, 23, 2) {real, imag} */,
  {32'hbf685fde, 32'h00000000} /* (21, 23, 1) {real, imag} */,
  {32'hbec59472, 32'h00000000} /* (21, 23, 0) {real, imag} */,
  {32'hbee3b7ec, 32'h00000000} /* (21, 22, 31) {real, imag} */,
  {32'hbf7ce3b1, 32'h00000000} /* (21, 22, 30) {real, imag} */,
  {32'hbf63f466, 32'h00000000} /* (21, 22, 29) {real, imag} */,
  {32'hbf443039, 32'h00000000} /* (21, 22, 28) {real, imag} */,
  {32'hbf12f46b, 32'h00000000} /* (21, 22, 27) {real, imag} */,
  {32'hbe9caad5, 32'h00000000} /* (21, 22, 26) {real, imag} */,
  {32'hbe776649, 32'h00000000} /* (21, 22, 25) {real, imag} */,
  {32'hbf16d344, 32'h00000000} /* (21, 22, 24) {real, imag} */,
  {32'hbf7aedaa, 32'h00000000} /* (21, 22, 23) {real, imag} */,
  {32'hbf3f2a9d, 32'h00000000} /* (21, 22, 22) {real, imag} */,
  {32'hbeb3e7c9, 32'h00000000} /* (21, 22, 21) {real, imag} */,
  {32'h3f700221, 32'h00000000} /* (21, 22, 20) {real, imag} */,
  {32'h3f71239f, 32'h00000000} /* (21, 22, 19) {real, imag} */,
  {32'h3f52aebb, 32'h00000000} /* (21, 22, 18) {real, imag} */,
  {32'h3ebc4d04, 32'h00000000} /* (21, 22, 17) {real, imag} */,
  {32'h3f5b221d, 32'h00000000} /* (21, 22, 16) {real, imag} */,
  {32'h3f6738ba, 32'h00000000} /* (21, 22, 15) {real, imag} */,
  {32'h3f260b86, 32'h00000000} /* (21, 22, 14) {real, imag} */,
  {32'h3fa3ea18, 32'h00000000} /* (21, 22, 13) {real, imag} */,
  {32'h3fa40d9c, 32'h00000000} /* (21, 22, 12) {real, imag} */,
  {32'h3f230346, 32'h00000000} /* (21, 22, 11) {real, imag} */,
  {32'hbea8b1c3, 32'h00000000} /* (21, 22, 10) {real, imag} */,
  {32'hbe8c90b8, 32'h00000000} /* (21, 22, 9) {real, imag} */,
  {32'hbf02e6f7, 32'h00000000} /* (21, 22, 8) {real, imag} */,
  {32'hbf597d5c, 32'h00000000} /* (21, 22, 7) {real, imag} */,
  {32'hbf481834, 32'h00000000} /* (21, 22, 6) {real, imag} */,
  {32'hbf822369, 32'h00000000} /* (21, 22, 5) {real, imag} */,
  {32'hbfb9f18c, 32'h00000000} /* (21, 22, 4) {real, imag} */,
  {32'hbfd1084c, 32'h00000000} /* (21, 22, 3) {real, imag} */,
  {32'hbf6b286c, 32'h00000000} /* (21, 22, 2) {real, imag} */,
  {32'hbfbaaf61, 32'h00000000} /* (21, 22, 1) {real, imag} */,
  {32'hbf284f1c, 32'h00000000} /* (21, 22, 0) {real, imag} */,
  {32'hbe9b9cfc, 32'h00000000} /* (21, 21, 31) {real, imag} */,
  {32'hbe9a9881, 32'h00000000} /* (21, 21, 30) {real, imag} */,
  {32'hbd910307, 32'h00000000} /* (21, 21, 29) {real, imag} */,
  {32'hbdaf26ee, 32'h00000000} /* (21, 21, 28) {real, imag} */,
  {32'h3dd52c06, 32'h00000000} /* (21, 21, 27) {real, imag} */,
  {32'hbe1bba55, 32'h00000000} /* (21, 21, 26) {real, imag} */,
  {32'h3c68f803, 32'h00000000} /* (21, 21, 25) {real, imag} */,
  {32'h3e02c4ce, 32'h00000000} /* (21, 21, 24) {real, imag} */,
  {32'hbe5f6560, 32'h00000000} /* (21, 21, 23) {real, imag} */,
  {32'hbdd8aa97, 32'h00000000} /* (21, 21, 22) {real, imag} */,
  {32'hbbcad28a, 32'h00000000} /* (21, 21, 21) {real, imag} */,
  {32'h3d205500, 32'h00000000} /* (21, 21, 20) {real, imag} */,
  {32'h3ec04cdb, 32'h00000000} /* (21, 21, 19) {real, imag} */,
  {32'h3e39e91a, 32'h00000000} /* (21, 21, 18) {real, imag} */,
  {32'hbebc834c, 32'h00000000} /* (21, 21, 17) {real, imag} */,
  {32'hbcacbd3e, 32'h00000000} /* (21, 21, 16) {real, imag} */,
  {32'h3ef6cbe0, 32'h00000000} /* (21, 21, 15) {real, imag} */,
  {32'h3ecac803, 32'h00000000} /* (21, 21, 14) {real, imag} */,
  {32'h3f32f939, 32'h00000000} /* (21, 21, 13) {real, imag} */,
  {32'h3f6cc673, 32'h00000000} /* (21, 21, 12) {real, imag} */,
  {32'h3f116e7d, 32'h00000000} /* (21, 21, 11) {real, imag} */,
  {32'hbe9d5e94, 32'h00000000} /* (21, 21, 10) {real, imag} */,
  {32'h3e660a13, 32'h00000000} /* (21, 21, 9) {real, imag} */,
  {32'h3dd5d37d, 32'h00000000} /* (21, 21, 8) {real, imag} */,
  {32'hbe829d93, 32'h00000000} /* (21, 21, 7) {real, imag} */,
  {32'hbdb185dd, 32'h00000000} /* (21, 21, 6) {real, imag} */,
  {32'hbdbcc945, 32'h00000000} /* (21, 21, 5) {real, imag} */,
  {32'hbe4c1e11, 32'h00000000} /* (21, 21, 4) {real, imag} */,
  {32'hbe840064, 32'h00000000} /* (21, 21, 3) {real, imag} */,
  {32'hbe8ea157, 32'h00000000} /* (21, 21, 2) {real, imag} */,
  {32'hbf9095ef, 32'h00000000} /* (21, 21, 1) {real, imag} */,
  {32'hbf0b3c23, 32'h00000000} /* (21, 21, 0) {real, imag} */,
  {32'h3e68d07a, 32'h00000000} /* (21, 20, 31) {real, imag} */,
  {32'h3f497252, 32'h00000000} /* (21, 20, 30) {real, imag} */,
  {32'h3f8faac8, 32'h00000000} /* (21, 20, 29) {real, imag} */,
  {32'h3f4b6f80, 32'h00000000} /* (21, 20, 28) {real, imag} */,
  {32'h3f8c6599, 32'h00000000} /* (21, 20, 27) {real, imag} */,
  {32'h3f26692f, 32'h00000000} /* (21, 20, 26) {real, imag} */,
  {32'h3f5d14aa, 32'h00000000} /* (21, 20, 25) {real, imag} */,
  {32'h3f8b759d, 32'h00000000} /* (21, 20, 24) {real, imag} */,
  {32'h3ee6f629, 32'h00000000} /* (21, 20, 23) {real, imag} */,
  {32'h3eecfb72, 32'h00000000} /* (21, 20, 22) {real, imag} */,
  {32'h3e83060f, 32'h00000000} /* (21, 20, 21) {real, imag} */,
  {32'hbeeeb165, 32'h00000000} /* (21, 20, 20) {real, imag} */,
  {32'hbf0a1a0f, 32'h00000000} /* (21, 20, 19) {real, imag} */,
  {32'hbf6a2d97, 32'h00000000} /* (21, 20, 18) {real, imag} */,
  {32'hbffd5e3b, 32'h00000000} /* (21, 20, 17) {real, imag} */,
  {32'hbf9722a1, 32'h00000000} /* (21, 20, 16) {real, imag} */,
  {32'hbf06d4ad, 32'h00000000} /* (21, 20, 15) {real, imag} */,
  {32'hbf194ec4, 32'h00000000} /* (21, 20, 14) {real, imag} */,
  {32'hbf65bab9, 32'h00000000} /* (21, 20, 13) {real, imag} */,
  {32'hbe9d0e73, 32'h00000000} /* (21, 20, 12) {real, imag} */,
  {32'hbf150bfb, 32'h00000000} /* (21, 20, 11) {real, imag} */,
  {32'hbdb2f561, 32'h00000000} /* (21, 20, 10) {real, imag} */,
  {32'h3f6dd4a7, 32'h00000000} /* (21, 20, 9) {real, imag} */,
  {32'h3efcb9cd, 32'h00000000} /* (21, 20, 8) {real, imag} */,
  {32'h3e8feaa0, 32'h00000000} /* (21, 20, 7) {real, imag} */,
  {32'h3f6c07bf, 32'h00000000} /* (21, 20, 6) {real, imag} */,
  {32'h3f8039ba, 32'h00000000} /* (21, 20, 5) {real, imag} */,
  {32'h3f9a98bd, 32'h00000000} /* (21, 20, 4) {real, imag} */,
  {32'h3f97a958, 32'h00000000} /* (21, 20, 3) {real, imag} */,
  {32'h3f49f21d, 32'h00000000} /* (21, 20, 2) {real, imag} */,
  {32'hbdbacf1c, 32'h00000000} /* (21, 20, 1) {real, imag} */,
  {32'hbe2b6e9c, 32'h00000000} /* (21, 20, 0) {real, imag} */,
  {32'h3e987d8b, 32'h00000000} /* (21, 19, 31) {real, imag} */,
  {32'h3f3c2b68, 32'h00000000} /* (21, 19, 30) {real, imag} */,
  {32'h3fa90269, 32'h00000000} /* (21, 19, 29) {real, imag} */,
  {32'h3f94f657, 32'h00000000} /* (21, 19, 28) {real, imag} */,
  {32'h3f83cf19, 32'h00000000} /* (21, 19, 27) {real, imag} */,
  {32'h3f5a5693, 32'h00000000} /* (21, 19, 26) {real, imag} */,
  {32'h3f61b8a6, 32'h00000000} /* (21, 19, 25) {real, imag} */,
  {32'h3f91628c, 32'h00000000} /* (21, 19, 24) {real, imag} */,
  {32'h3f871548, 32'h00000000} /* (21, 19, 23) {real, imag} */,
  {32'h3f2a73f7, 32'h00000000} /* (21, 19, 22) {real, imag} */,
  {32'h3e0c46a9, 32'h00000000} /* (21, 19, 21) {real, imag} */,
  {32'hbf1c27aa, 32'h00000000} /* (21, 19, 20) {real, imag} */,
  {32'hbf10a324, 32'h00000000} /* (21, 19, 19) {real, imag} */,
  {32'hbf85c62e, 32'h00000000} /* (21, 19, 18) {real, imag} */,
  {32'hbfd377d8, 32'h00000000} /* (21, 19, 17) {real, imag} */,
  {32'hbfc439a3, 32'h00000000} /* (21, 19, 16) {real, imag} */,
  {32'hbfbad69f, 32'h00000000} /* (21, 19, 15) {real, imag} */,
  {32'hbfa58d57, 32'h00000000} /* (21, 19, 14) {real, imag} */,
  {32'hbfc84f66, 32'h00000000} /* (21, 19, 13) {real, imag} */,
  {32'hbfa4b3f0, 32'h00000000} /* (21, 19, 12) {real, imag} */,
  {32'hbf49ba9b, 32'h00000000} /* (21, 19, 11) {real, imag} */,
  {32'h3da050ea, 32'h00000000} /* (21, 19, 10) {real, imag} */,
  {32'h3f1ebdfb, 32'h00000000} /* (21, 19, 9) {real, imag} */,
  {32'h3eb9aad9, 32'h00000000} /* (21, 19, 8) {real, imag} */,
  {32'h3e9005c6, 32'h00000000} /* (21, 19, 7) {real, imag} */,
  {32'h3f7384cd, 32'h00000000} /* (21, 19, 6) {real, imag} */,
  {32'h3f383449, 32'h00000000} /* (21, 19, 5) {real, imag} */,
  {32'h3f082f94, 32'h00000000} /* (21, 19, 4) {real, imag} */,
  {32'h3f7cf90f, 32'h00000000} /* (21, 19, 3) {real, imag} */,
  {32'h3faf2c0f, 32'h00000000} /* (21, 19, 2) {real, imag} */,
  {32'h3f0d67ea, 32'h00000000} /* (21, 19, 1) {real, imag} */,
  {32'h3b5d8d1d, 32'h00000000} /* (21, 19, 0) {real, imag} */,
  {32'h3ead6f21, 32'h00000000} /* (21, 18, 31) {real, imag} */,
  {32'h3f1a30cb, 32'h00000000} /* (21, 18, 30) {real, imag} */,
  {32'h3fa1dd72, 32'h00000000} /* (21, 18, 29) {real, imag} */,
  {32'h3fa9a042, 32'h00000000} /* (21, 18, 28) {real, imag} */,
  {32'h3f8ceffc, 32'h00000000} /* (21, 18, 27) {real, imag} */,
  {32'h3f69459b, 32'h00000000} /* (21, 18, 26) {real, imag} */,
  {32'h3f8d897a, 32'h00000000} /* (21, 18, 25) {real, imag} */,
  {32'h3f909dd4, 32'h00000000} /* (21, 18, 24) {real, imag} */,
  {32'h3fa7052e, 32'h00000000} /* (21, 18, 23) {real, imag} */,
  {32'h3f11d3e4, 32'h00000000} /* (21, 18, 22) {real, imag} */,
  {32'hbd3cdaa5, 32'h00000000} /* (21, 18, 21) {real, imag} */,
  {32'hbd6aebaf, 32'h00000000} /* (21, 18, 20) {real, imag} */,
  {32'hbf14e37c, 32'h00000000} /* (21, 18, 19) {real, imag} */,
  {32'hbfc00dbe, 32'h00000000} /* (21, 18, 18) {real, imag} */,
  {32'hbfb5f3d6, 32'h00000000} /* (21, 18, 17) {real, imag} */,
  {32'hbfcfe1d1, 32'h00000000} /* (21, 18, 16) {real, imag} */,
  {32'hbfc8009d, 32'h00000000} /* (21, 18, 15) {real, imag} */,
  {32'hbf4d44bb, 32'h00000000} /* (21, 18, 14) {real, imag} */,
  {32'hbf4492f5, 32'h00000000} /* (21, 18, 13) {real, imag} */,
  {32'hbf636073, 32'h00000000} /* (21, 18, 12) {real, imag} */,
  {32'hbf02daaf, 32'h00000000} /* (21, 18, 11) {real, imag} */,
  {32'hbd6bb058, 32'h00000000} /* (21, 18, 10) {real, imag} */,
  {32'h3eb147fd, 32'h00000000} /* (21, 18, 9) {real, imag} */,
  {32'h3f5d8146, 32'h00000000} /* (21, 18, 8) {real, imag} */,
  {32'h3f6774dd, 32'h00000000} /* (21, 18, 7) {real, imag} */,
  {32'h3f84e7fa, 32'h00000000} /* (21, 18, 6) {real, imag} */,
  {32'h3f8ff91b, 32'h00000000} /* (21, 18, 5) {real, imag} */,
  {32'h3f204274, 32'h00000000} /* (21, 18, 4) {real, imag} */,
  {32'h3f18263b, 32'h00000000} /* (21, 18, 3) {real, imag} */,
  {32'h3fa252a5, 32'h00000000} /* (21, 18, 2) {real, imag} */,
  {32'h3fa4b236, 32'h00000000} /* (21, 18, 1) {real, imag} */,
  {32'h3edd48ed, 32'h00000000} /* (21, 18, 0) {real, imag} */,
  {32'h3db9219f, 32'h00000000} /* (21, 17, 31) {real, imag} */,
  {32'h3ee5bc91, 32'h00000000} /* (21, 17, 30) {real, imag} */,
  {32'h3f829683, 32'h00000000} /* (21, 17, 29) {real, imag} */,
  {32'h3fa63d88, 32'h00000000} /* (21, 17, 28) {real, imag} */,
  {32'h3fa0162b, 32'h00000000} /* (21, 17, 27) {real, imag} */,
  {32'h3f857f84, 32'h00000000} /* (21, 17, 26) {real, imag} */,
  {32'h3f987f51, 32'h00000000} /* (21, 17, 25) {real, imag} */,
  {32'h3fae71b3, 32'h00000000} /* (21, 17, 24) {real, imag} */,
  {32'h3fb9538b, 32'h00000000} /* (21, 17, 23) {real, imag} */,
  {32'h3f406f5b, 32'h00000000} /* (21, 17, 22) {real, imag} */,
  {32'h3e9ac219, 32'h00000000} /* (21, 17, 21) {real, imag} */,
  {32'hbe50806d, 32'h00000000} /* (21, 17, 20) {real, imag} */,
  {32'hbf9a5640, 32'h00000000} /* (21, 17, 19) {real, imag} */,
  {32'hbfeb0b8c, 32'h00000000} /* (21, 17, 18) {real, imag} */,
  {32'hbfc7069f, 32'h00000000} /* (21, 17, 17) {real, imag} */,
  {32'hbf8faea8, 32'h00000000} /* (21, 17, 16) {real, imag} */,
  {32'hbf699d3d, 32'h00000000} /* (21, 17, 15) {real, imag} */,
  {32'hbf5c3fa6, 32'h00000000} /* (21, 17, 14) {real, imag} */,
  {32'hbf649f6c, 32'h00000000} /* (21, 17, 13) {real, imag} */,
  {32'hbf547691, 32'h00000000} /* (21, 17, 12) {real, imag} */,
  {32'hbf4297c3, 32'h00000000} /* (21, 17, 11) {real, imag} */,
  {32'hbe204ddc, 32'h00000000} /* (21, 17, 10) {real, imag} */,
  {32'h3ebfa173, 32'h00000000} /* (21, 17, 9) {real, imag} */,
  {32'h3f27b55e, 32'h00000000} /* (21, 17, 8) {real, imag} */,
  {32'h3f336558, 32'h00000000} /* (21, 17, 7) {real, imag} */,
  {32'h3f46d1f9, 32'h00000000} /* (21, 17, 6) {real, imag} */,
  {32'h3fc7d24e, 32'h00000000} /* (21, 17, 5) {real, imag} */,
  {32'h3f91f819, 32'h00000000} /* (21, 17, 4) {real, imag} */,
  {32'h3f56a74d, 32'h00000000} /* (21, 17, 3) {real, imag} */,
  {32'h3fcca251, 32'h00000000} /* (21, 17, 2) {real, imag} */,
  {32'h3ffaed28, 32'h00000000} /* (21, 17, 1) {real, imag} */,
  {32'h3f10e82f, 32'h00000000} /* (21, 17, 0) {real, imag} */,
  {32'h3f0035be, 32'h00000000} /* (21, 16, 31) {real, imag} */,
  {32'h3f8005ac, 32'h00000000} /* (21, 16, 30) {real, imag} */,
  {32'h3f57186e, 32'h00000000} /* (21, 16, 29) {real, imag} */,
  {32'h3f6954a6, 32'h00000000} /* (21, 16, 28) {real, imag} */,
  {32'h3f4235ab, 32'h00000000} /* (21, 16, 27) {real, imag} */,
  {32'h3f8b9a2c, 32'h00000000} /* (21, 16, 26) {real, imag} */,
  {32'h3f883ca6, 32'h00000000} /* (21, 16, 25) {real, imag} */,
  {32'h3f717ac5, 32'h00000000} /* (21, 16, 24) {real, imag} */,
  {32'h3f85dac0, 32'h00000000} /* (21, 16, 23) {real, imag} */,
  {32'h3f4beee7, 32'h00000000} /* (21, 16, 22) {real, imag} */,
  {32'h3e6beafe, 32'h00000000} /* (21, 16, 21) {real, imag} */,
  {32'hbf95b992, 32'h00000000} /* (21, 16, 20) {real, imag} */,
  {32'hbfb9fb6e, 32'h00000000} /* (21, 16, 19) {real, imag} */,
  {32'hbf96280a, 32'h00000000} /* (21, 16, 18) {real, imag} */,
  {32'hbf26eb7a, 32'h00000000} /* (21, 16, 17) {real, imag} */,
  {32'hbe4c1343, 32'h00000000} /* (21, 16, 16) {real, imag} */,
  {32'hbf331962, 32'h00000000} /* (21, 16, 15) {real, imag} */,
  {32'hbfa89091, 32'h00000000} /* (21, 16, 14) {real, imag} */,
  {32'hbfaee716, 32'h00000000} /* (21, 16, 13) {real, imag} */,
  {32'hbf6fb288, 32'h00000000} /* (21, 16, 12) {real, imag} */,
  {32'hbf5994f3, 32'h00000000} /* (21, 16, 11) {real, imag} */,
  {32'h3e0387d3, 32'h00000000} /* (21, 16, 10) {real, imag} */,
  {32'h3f50eab8, 32'h00000000} /* (21, 16, 9) {real, imag} */,
  {32'h3efd7f78, 32'h00000000} /* (21, 16, 8) {real, imag} */,
  {32'h3eb1894e, 32'h00000000} /* (21, 16, 7) {real, imag} */,
  {32'h3f333e90, 32'h00000000} /* (21, 16, 6) {real, imag} */,
  {32'h3fb02a0f, 32'h00000000} /* (21, 16, 5) {real, imag} */,
  {32'h3f9926bd, 32'h00000000} /* (21, 16, 4) {real, imag} */,
  {32'h3f96cd17, 32'h00000000} /* (21, 16, 3) {real, imag} */,
  {32'h3f9905ce, 32'h00000000} /* (21, 16, 2) {real, imag} */,
  {32'h3fb7df5b, 32'h00000000} /* (21, 16, 1) {real, imag} */,
  {32'h3f24c574, 32'h00000000} /* (21, 16, 0) {real, imag} */,
  {32'h3f374fa6, 32'h00000000} /* (21, 15, 31) {real, imag} */,
  {32'h3fbe5a17, 32'h00000000} /* (21, 15, 30) {real, imag} */,
  {32'h3f96dae0, 32'h00000000} /* (21, 15, 29) {real, imag} */,
  {32'h3f732ae7, 32'h00000000} /* (21, 15, 28) {real, imag} */,
  {32'h3f206631, 32'h00000000} /* (21, 15, 27) {real, imag} */,
  {32'h3f9764f5, 32'h00000000} /* (21, 15, 26) {real, imag} */,
  {32'h3fc671c7, 32'h00000000} /* (21, 15, 25) {real, imag} */,
  {32'h3f269330, 32'h00000000} /* (21, 15, 24) {real, imag} */,
  {32'h3f2ed8d2, 32'h00000000} /* (21, 15, 23) {real, imag} */,
  {32'h3f0a775d, 32'h00000000} /* (21, 15, 22) {real, imag} */,
  {32'h3e406888, 32'h00000000} /* (21, 15, 21) {real, imag} */,
  {32'hbf9d1f7d, 32'h00000000} /* (21, 15, 20) {real, imag} */,
  {32'hbf7fb5f3, 32'h00000000} /* (21, 15, 19) {real, imag} */,
  {32'hbf3bfa62, 32'h00000000} /* (21, 15, 18) {real, imag} */,
  {32'hbf1c99cc, 32'h00000000} /* (21, 15, 17) {real, imag} */,
  {32'hbefcee46, 32'h00000000} /* (21, 15, 16) {real, imag} */,
  {32'hbf526309, 32'h00000000} /* (21, 15, 15) {real, imag} */,
  {32'hbf5959ca, 32'h00000000} /* (21, 15, 14) {real, imag} */,
  {32'hbf884aef, 32'h00000000} /* (21, 15, 13) {real, imag} */,
  {32'hbfacebd1, 32'h00000000} /* (21, 15, 12) {real, imag} */,
  {32'hbfa4d76e, 32'h00000000} /* (21, 15, 11) {real, imag} */,
  {32'hbc487a27, 32'h00000000} /* (21, 15, 10) {real, imag} */,
  {32'h3f30d421, 32'h00000000} /* (21, 15, 9) {real, imag} */,
  {32'h3ef6a75d, 32'h00000000} /* (21, 15, 8) {real, imag} */,
  {32'h3ed65b9c, 32'h00000000} /* (21, 15, 7) {real, imag} */,
  {32'h3ed9a91e, 32'h00000000} /* (21, 15, 6) {real, imag} */,
  {32'h3f870824, 32'h00000000} /* (21, 15, 5) {real, imag} */,
  {32'h3fd85eb2, 32'h00000000} /* (21, 15, 4) {real, imag} */,
  {32'h3fc4adbf, 32'h00000000} /* (21, 15, 3) {real, imag} */,
  {32'h3f84acfd, 32'h00000000} /* (21, 15, 2) {real, imag} */,
  {32'h3fab7c04, 32'h00000000} /* (21, 15, 1) {real, imag} */,
  {32'h3ef59fad, 32'h00000000} /* (21, 15, 0) {real, imag} */,
  {32'h3ef9927d, 32'h00000000} /* (21, 14, 31) {real, imag} */,
  {32'h3fb22bbf, 32'h00000000} /* (21, 14, 30) {real, imag} */,
  {32'h3fc94921, 32'h00000000} /* (21, 14, 29) {real, imag} */,
  {32'h3f8f1c6a, 32'h00000000} /* (21, 14, 28) {real, imag} */,
  {32'h3f87d305, 32'h00000000} /* (21, 14, 27) {real, imag} */,
  {32'h3fab9e20, 32'h00000000} /* (21, 14, 26) {real, imag} */,
  {32'h3fade721, 32'h00000000} /* (21, 14, 25) {real, imag} */,
  {32'h3f24f07a, 32'h00000000} /* (21, 14, 24) {real, imag} */,
  {32'h3f0d392a, 32'h00000000} /* (21, 14, 23) {real, imag} */,
  {32'h3f473173, 32'h00000000} /* (21, 14, 22) {real, imag} */,
  {32'h3ea572ac, 32'h00000000} /* (21, 14, 21) {real, imag} */,
  {32'hbf30ad08, 32'h00000000} /* (21, 14, 20) {real, imag} */,
  {32'hbf1086cf, 32'h00000000} /* (21, 14, 19) {real, imag} */,
  {32'hbef53d84, 32'h00000000} /* (21, 14, 18) {real, imag} */,
  {32'hbf433472, 32'h00000000} /* (21, 14, 17) {real, imag} */,
  {32'hbf531089, 32'h00000000} /* (21, 14, 16) {real, imag} */,
  {32'hbf837462, 32'h00000000} /* (21, 14, 15) {real, imag} */,
  {32'hbf21e587, 32'h00000000} /* (21, 14, 14) {real, imag} */,
  {32'hbf5ce9ef, 32'h00000000} /* (21, 14, 13) {real, imag} */,
  {32'hbfb112a0, 32'h00000000} /* (21, 14, 12) {real, imag} */,
  {32'hbfb8b513, 32'h00000000} /* (21, 14, 11) {real, imag} */,
  {32'hbe832061, 32'h00000000} /* (21, 14, 10) {real, imag} */,
  {32'h3f063ab3, 32'h00000000} /* (21, 14, 9) {real, imag} */,
  {32'h3f884cfc, 32'h00000000} /* (21, 14, 8) {real, imag} */,
  {32'h3f897512, 32'h00000000} /* (21, 14, 7) {real, imag} */,
  {32'h3f271679, 32'h00000000} /* (21, 14, 6) {real, imag} */,
  {32'h3f900f84, 32'h00000000} /* (21, 14, 5) {real, imag} */,
  {32'h3fa46b4e, 32'h00000000} /* (21, 14, 4) {real, imag} */,
  {32'h3f444380, 32'h00000000} /* (21, 14, 3) {real, imag} */,
  {32'h3f9b1924, 32'h00000000} /* (21, 14, 2) {real, imag} */,
  {32'h3ff15c2e, 32'h00000000} /* (21, 14, 1) {real, imag} */,
  {32'h3f3c5b22, 32'h00000000} /* (21, 14, 0) {real, imag} */,
  {32'h3ec62a07, 32'h00000000} /* (21, 13, 31) {real, imag} */,
  {32'h3f6c40b6, 32'h00000000} /* (21, 13, 30) {real, imag} */,
  {32'h3f94d18f, 32'h00000000} /* (21, 13, 29) {real, imag} */,
  {32'h3f86b776, 32'h00000000} /* (21, 13, 28) {real, imag} */,
  {32'h3fc8fd98, 32'h00000000} /* (21, 13, 27) {real, imag} */,
  {32'h3faa21d2, 32'h00000000} /* (21, 13, 26) {real, imag} */,
  {32'h3f02ff0e, 32'h00000000} /* (21, 13, 25) {real, imag} */,
  {32'h3f0268a8, 32'h00000000} /* (21, 13, 24) {real, imag} */,
  {32'h3f4671de, 32'h00000000} /* (21, 13, 23) {real, imag} */,
  {32'h3fd0f3ac, 32'h00000000} /* (21, 13, 22) {real, imag} */,
  {32'h3ed6f221, 32'h00000000} /* (21, 13, 21) {real, imag} */,
  {32'hbf1a221f, 32'h00000000} /* (21, 13, 20) {real, imag} */,
  {32'hbf99eea1, 32'h00000000} /* (21, 13, 19) {real, imag} */,
  {32'hbf631d69, 32'h00000000} /* (21, 13, 18) {real, imag} */,
  {32'hbf0d5697, 32'h00000000} /* (21, 13, 17) {real, imag} */,
  {32'hbf20b4de, 32'h00000000} /* (21, 13, 16) {real, imag} */,
  {32'hbf1e28b7, 32'h00000000} /* (21, 13, 15) {real, imag} */,
  {32'hbf5b5764, 32'h00000000} /* (21, 13, 14) {real, imag} */,
  {32'hbf84f59e, 32'h00000000} /* (21, 13, 13) {real, imag} */,
  {32'hbf887352, 32'h00000000} /* (21, 13, 12) {real, imag} */,
  {32'hbfba2243, 32'h00000000} /* (21, 13, 11) {real, imag} */,
  {32'hbdf84a47, 32'h00000000} /* (21, 13, 10) {real, imag} */,
  {32'h3f534029, 32'h00000000} /* (21, 13, 9) {real, imag} */,
  {32'h3fc3e1f4, 32'h00000000} /* (21, 13, 8) {real, imag} */,
  {32'h3f94e975, 32'h00000000} /* (21, 13, 7) {real, imag} */,
  {32'h3f1c04e1, 32'h00000000} /* (21, 13, 6) {real, imag} */,
  {32'h3f93f40a, 32'h00000000} /* (21, 13, 5) {real, imag} */,
  {32'h3f9067fa, 32'h00000000} /* (21, 13, 4) {real, imag} */,
  {32'h3ee72303, 32'h00000000} /* (21, 13, 3) {real, imag} */,
  {32'h3f69a84d, 32'h00000000} /* (21, 13, 2) {real, imag} */,
  {32'h3fd92590, 32'h00000000} /* (21, 13, 1) {real, imag} */,
  {32'h3f5c8ac5, 32'h00000000} /* (21, 13, 0) {real, imag} */,
  {32'h3ed3429e, 32'h00000000} /* (21, 12, 31) {real, imag} */,
  {32'h3f09a8e8, 32'h00000000} /* (21, 12, 30) {real, imag} */,
  {32'h3ea64fab, 32'h00000000} /* (21, 12, 29) {real, imag} */,
  {32'h3f3894cb, 32'h00000000} /* (21, 12, 28) {real, imag} */,
  {32'h3f952eea, 32'h00000000} /* (21, 12, 27) {real, imag} */,
  {32'h3f11e02d, 32'h00000000} /* (21, 12, 26) {real, imag} */,
  {32'h3e9995a7, 32'h00000000} /* (21, 12, 25) {real, imag} */,
  {32'h3f49b287, 32'h00000000} /* (21, 12, 24) {real, imag} */,
  {32'h3fb03085, 32'h00000000} /* (21, 12, 23) {real, imag} */,
  {32'h3ff942b1, 32'h00000000} /* (21, 12, 22) {real, imag} */,
  {32'h3eeb9894, 32'h00000000} /* (21, 12, 21) {real, imag} */,
  {32'hbf35accc, 32'h00000000} /* (21, 12, 20) {real, imag} */,
  {32'hbf8f0780, 32'h00000000} /* (21, 12, 19) {real, imag} */,
  {32'hbf9e5f1a, 32'h00000000} /* (21, 12, 18) {real, imag} */,
  {32'hbf64520c, 32'h00000000} /* (21, 12, 17) {real, imag} */,
  {32'hbf11621f, 32'h00000000} /* (21, 12, 16) {real, imag} */,
  {32'hbf0c3e98, 32'h00000000} /* (21, 12, 15) {real, imag} */,
  {32'hbfada47e, 32'h00000000} /* (21, 12, 14) {real, imag} */,
  {32'hbf8b6180, 32'h00000000} /* (21, 12, 13) {real, imag} */,
  {32'hbf0bb30e, 32'h00000000} /* (21, 12, 12) {real, imag} */,
  {32'hbf1b6f89, 32'h00000000} /* (21, 12, 11) {real, imag} */,
  {32'h3f67ab53, 32'h00000000} /* (21, 12, 10) {real, imag} */,
  {32'h3f880c12, 32'h00000000} /* (21, 12, 9) {real, imag} */,
  {32'h3f79f6f5, 32'h00000000} /* (21, 12, 8) {real, imag} */,
  {32'h3f73064c, 32'h00000000} /* (21, 12, 7) {real, imag} */,
  {32'h3f1ba82c, 32'h00000000} /* (21, 12, 6) {real, imag} */,
  {32'h3f6827c7, 32'h00000000} /* (21, 12, 5) {real, imag} */,
  {32'h3f7f6a1b, 32'h00000000} /* (21, 12, 4) {real, imag} */,
  {32'h3e8fc5f6, 32'h00000000} /* (21, 12, 3) {real, imag} */,
  {32'h3ed086f8, 32'h00000000} /* (21, 12, 2) {real, imag} */,
  {32'h3f722afe, 32'h00000000} /* (21, 12, 1) {real, imag} */,
  {32'h3ec2022a, 32'h00000000} /* (21, 12, 0) {real, imag} */,
  {32'h3f252327, 32'h00000000} /* (21, 11, 31) {real, imag} */,
  {32'h3f5b1343, 32'h00000000} /* (21, 11, 30) {real, imag} */,
  {32'h3efafe2c, 32'h00000000} /* (21, 11, 29) {real, imag} */,
  {32'h3f0eddde, 32'h00000000} /* (21, 11, 28) {real, imag} */,
  {32'h3f0573b8, 32'h00000000} /* (21, 11, 27) {real, imag} */,
  {32'h3efb29a8, 32'h00000000} /* (21, 11, 26) {real, imag} */,
  {32'h3f2efa59, 32'h00000000} /* (21, 11, 25) {real, imag} */,
  {32'h3f6402d6, 32'h00000000} /* (21, 11, 24) {real, imag} */,
  {32'h3f69352c, 32'h00000000} /* (21, 11, 23) {real, imag} */,
  {32'h3fa85ae8, 32'h00000000} /* (21, 11, 22) {real, imag} */,
  {32'hbd2bfcdc, 32'h00000000} /* (21, 11, 21) {real, imag} */,
  {32'hbf15e344, 32'h00000000} /* (21, 11, 20) {real, imag} */,
  {32'hbed8719c, 32'h00000000} /* (21, 11, 19) {real, imag} */,
  {32'hbf0050d7, 32'h00000000} /* (21, 11, 18) {real, imag} */,
  {32'hbf1b707e, 32'h00000000} /* (21, 11, 17) {real, imag} */,
  {32'hbeeebdad, 32'h00000000} /* (21, 11, 16) {real, imag} */,
  {32'hbee216dd, 32'h00000000} /* (21, 11, 15) {real, imag} */,
  {32'hbefed46f, 32'h00000000} /* (21, 11, 14) {real, imag} */,
  {32'hbe454db5, 32'h00000000} /* (21, 11, 13) {real, imag} */,
  {32'hbdcbb329, 32'h00000000} /* (21, 11, 12) {real, imag} */,
  {32'hbded9a4b, 32'h00000000} /* (21, 11, 11) {real, imag} */,
  {32'h3f890c16, 32'h00000000} /* (21, 11, 10) {real, imag} */,
  {32'h3f4ed7bf, 32'h00000000} /* (21, 11, 9) {real, imag} */,
  {32'h3f2e8e32, 32'h00000000} /* (21, 11, 8) {real, imag} */,
  {32'h3f9637b0, 32'h00000000} /* (21, 11, 7) {real, imag} */,
  {32'h3f92afb6, 32'h00000000} /* (21, 11, 6) {real, imag} */,
  {32'h3f6cee64, 32'h00000000} /* (21, 11, 5) {real, imag} */,
  {32'h3f2fb3a3, 32'h00000000} /* (21, 11, 4) {real, imag} */,
  {32'h3e75d761, 32'h00000000} /* (21, 11, 3) {real, imag} */,
  {32'h3f203e4c, 32'h00000000} /* (21, 11, 2) {real, imag} */,
  {32'h3f610a0d, 32'h00000000} /* (21, 11, 1) {real, imag} */,
  {32'h3f003142, 32'h00000000} /* (21, 11, 0) {real, imag} */,
  {32'h3e5fa24a, 32'h00000000} /* (21, 10, 31) {real, imag} */,
  {32'h3e1b80f7, 32'h00000000} /* (21, 10, 30) {real, imag} */,
  {32'hbebb11e2, 32'h00000000} /* (21, 10, 29) {real, imag} */,
  {32'hbebe7e31, 32'h00000000} /* (21, 10, 28) {real, imag} */,
  {32'hbf626c82, 32'h00000000} /* (21, 10, 27) {real, imag} */,
  {32'hbeec1589, 32'h00000000} /* (21, 10, 26) {real, imag} */,
  {32'hbe090670, 32'h00000000} /* (21, 10, 25) {real, imag} */,
  {32'hbd9e6b9a, 32'h00000000} /* (21, 10, 24) {real, imag} */,
  {32'hbe925c0a, 32'h00000000} /* (21, 10, 23) {real, imag} */,
  {32'hbf135a02, 32'h00000000} /* (21, 10, 22) {real, imag} */,
  {32'hbf0b622c, 32'h00000000} /* (21, 10, 21) {real, imag} */,
  {32'h3f2f6185, 32'h00000000} /* (21, 10, 20) {real, imag} */,
  {32'h3f0a7cea, 32'h00000000} /* (21, 10, 19) {real, imag} */,
  {32'h3dd602fe, 32'h00000000} /* (21, 10, 18) {real, imag} */,
  {32'h3e068a8a, 32'h00000000} /* (21, 10, 17) {real, imag} */,
  {32'h3f1a5410, 32'h00000000} /* (21, 10, 16) {real, imag} */,
  {32'h3ec05782, 32'h00000000} /* (21, 10, 15) {real, imag} */,
  {32'h3ebd3aa2, 32'h00000000} /* (21, 10, 14) {real, imag} */,
  {32'h3ecda4ca, 32'h00000000} /* (21, 10, 13) {real, imag} */,
  {32'h3f195752, 32'h00000000} /* (21, 10, 12) {real, imag} */,
  {32'h3ead01c6, 32'h00000000} /* (21, 10, 11) {real, imag} */,
  {32'h3cd39296, 32'h00000000} /* (21, 10, 10) {real, imag} */,
  {32'hbf317061, 32'h00000000} /* (21, 10, 9) {real, imag} */,
  {32'hbe76fc1e, 32'h00000000} /* (21, 10, 8) {real, imag} */,
  {32'h3e7695f2, 32'h00000000} /* (21, 10, 7) {real, imag} */,
  {32'hbcf9cd11, 32'h00000000} /* (21, 10, 6) {real, imag} */,
  {32'hbea9be90, 32'h00000000} /* (21, 10, 5) {real, imag} */,
  {32'hbf01e6d2, 32'h00000000} /* (21, 10, 4) {real, imag} */,
  {32'hbf05c835, 32'h00000000} /* (21, 10, 3) {real, imag} */,
  {32'hbd0569d6, 32'h00000000} /* (21, 10, 2) {real, imag} */,
  {32'hbd615ba4, 32'h00000000} /* (21, 10, 1) {real, imag} */,
  {32'hbdb5c6a3, 32'h00000000} /* (21, 10, 0) {real, imag} */,
  {32'hbda65cce, 32'h00000000} /* (21, 9, 31) {real, imag} */,
  {32'hbeeb78fc, 32'h00000000} /* (21, 9, 30) {real, imag} */,
  {32'hbf973887, 32'h00000000} /* (21, 9, 29) {real, imag} */,
  {32'hbf4ccce0, 32'h00000000} /* (21, 9, 28) {real, imag} */,
  {32'hbf61ed21, 32'h00000000} /* (21, 9, 27) {real, imag} */,
  {32'hbf535c14, 32'h00000000} /* (21, 9, 26) {real, imag} */,
  {32'hbf080807, 32'h00000000} /* (21, 9, 25) {real, imag} */,
  {32'hbf003a51, 32'h00000000} /* (21, 9, 24) {real, imag} */,
  {32'hbf5377c6, 32'h00000000} /* (21, 9, 23) {real, imag} */,
  {32'hbf603208, 32'h00000000} /* (21, 9, 22) {real, imag} */,
  {32'hbf41d6a0, 32'h00000000} /* (21, 9, 21) {real, imag} */,
  {32'h3f8a2e45, 32'h00000000} /* (21, 9, 20) {real, imag} */,
  {32'h3f6c252e, 32'h00000000} /* (21, 9, 19) {real, imag} */,
  {32'h3eff0ed6, 32'h00000000} /* (21, 9, 18) {real, imag} */,
  {32'h3f0f0c7f, 32'h00000000} /* (21, 9, 17) {real, imag} */,
  {32'h3f89191d, 32'h00000000} /* (21, 9, 16) {real, imag} */,
  {32'h3f6acb82, 32'h00000000} /* (21, 9, 15) {real, imag} */,
  {32'h3f3209bc, 32'h00000000} /* (21, 9, 14) {real, imag} */,
  {32'h3f0554cb, 32'h00000000} /* (21, 9, 13) {real, imag} */,
  {32'h3f1185e2, 32'h00000000} /* (21, 9, 12) {real, imag} */,
  {32'h3f4904c6, 32'h00000000} /* (21, 9, 11) {real, imag} */,
  {32'hbd309b71, 32'h00000000} /* (21, 9, 10) {real, imag} */,
  {32'hbf969769, 32'h00000000} /* (21, 9, 9) {real, imag} */,
  {32'hbf94f89d, 32'h00000000} /* (21, 9, 8) {real, imag} */,
  {32'hbf867340, 32'h00000000} /* (21, 9, 7) {real, imag} */,
  {32'hbfb43f7c, 32'h00000000} /* (21, 9, 6) {real, imag} */,
  {32'hbf91b9bf, 32'h00000000} /* (21, 9, 5) {real, imag} */,
  {32'hbfb02fed, 32'h00000000} /* (21, 9, 4) {real, imag} */,
  {32'hbf7de6fa, 32'h00000000} /* (21, 9, 3) {real, imag} */,
  {32'hbf15a722, 32'h00000000} /* (21, 9, 2) {real, imag} */,
  {32'hbf00e147, 32'h00000000} /* (21, 9, 1) {real, imag} */,
  {32'hbe90d129, 32'h00000000} /* (21, 9, 0) {real, imag} */,
  {32'hbe9b19ae, 32'h00000000} /* (21, 8, 31) {real, imag} */,
  {32'hbf6f43df, 32'h00000000} /* (21, 8, 30) {real, imag} */,
  {32'hbfb7a004, 32'h00000000} /* (21, 8, 29) {real, imag} */,
  {32'hbf80678d, 32'h00000000} /* (21, 8, 28) {real, imag} */,
  {32'hbf068e1f, 32'h00000000} /* (21, 8, 27) {real, imag} */,
  {32'hbf5c9c54, 32'h00000000} /* (21, 8, 26) {real, imag} */,
  {32'hbf77a4b7, 32'h00000000} /* (21, 8, 25) {real, imag} */,
  {32'hbf206271, 32'h00000000} /* (21, 8, 24) {real, imag} */,
  {32'hbf5dd309, 32'h00000000} /* (21, 8, 23) {real, imag} */,
  {32'hbf904e99, 32'h00000000} /* (21, 8, 22) {real, imag} */,
  {32'hbf82705b, 32'h00000000} /* (21, 8, 21) {real, imag} */,
  {32'h3f2b22a8, 32'h00000000} /* (21, 8, 20) {real, imag} */,
  {32'h3f894c20, 32'h00000000} /* (21, 8, 19) {real, imag} */,
  {32'h3f5cf128, 32'h00000000} /* (21, 8, 18) {real, imag} */,
  {32'h3f655488, 32'h00000000} /* (21, 8, 17) {real, imag} */,
  {32'h3f4b2f9b, 32'h00000000} /* (21, 8, 16) {real, imag} */,
  {32'h3fa92de3, 32'h00000000} /* (21, 8, 15) {real, imag} */,
  {32'h3f96685c, 32'h00000000} /* (21, 8, 14) {real, imag} */,
  {32'h3f096186, 32'h00000000} /* (21, 8, 13) {real, imag} */,
  {32'h3ee05284, 32'h00000000} /* (21, 8, 12) {real, imag} */,
  {32'h3f761526, 32'h00000000} /* (21, 8, 11) {real, imag} */,
  {32'h3e3031a0, 32'h00000000} /* (21, 8, 10) {real, imag} */,
  {32'hbf39b5d5, 32'h00000000} /* (21, 8, 9) {real, imag} */,
  {32'hbf59cf94, 32'h00000000} /* (21, 8, 8) {real, imag} */,
  {32'hbf1798b2, 32'h00000000} /* (21, 8, 7) {real, imag} */,
  {32'hbf75315f, 32'h00000000} /* (21, 8, 6) {real, imag} */,
  {32'hbf6acab9, 32'h00000000} /* (21, 8, 5) {real, imag} */,
  {32'hbf43f953, 32'h00000000} /* (21, 8, 4) {real, imag} */,
  {32'hbf22c924, 32'h00000000} /* (21, 8, 3) {real, imag} */,
  {32'hbf6737cc, 32'h00000000} /* (21, 8, 2) {real, imag} */,
  {32'hbf2b15da, 32'h00000000} /* (21, 8, 1) {real, imag} */,
  {32'h3e21cefe, 32'h00000000} /* (21, 8, 0) {real, imag} */,
  {32'hbf2684b3, 32'h00000000} /* (21, 7, 31) {real, imag} */,
  {32'hbfab3fb7, 32'h00000000} /* (21, 7, 30) {real, imag} */,
  {32'hbfc312e4, 32'h00000000} /* (21, 7, 29) {real, imag} */,
  {32'hbf491958, 32'h00000000} /* (21, 7, 28) {real, imag} */,
  {32'hbf1a5eea, 32'h00000000} /* (21, 7, 27) {real, imag} */,
  {32'hbf8b295b, 32'h00000000} /* (21, 7, 26) {real, imag} */,
  {32'hbfb721e4, 32'h00000000} /* (21, 7, 25) {real, imag} */,
  {32'hbf63486a, 32'h00000000} /* (21, 7, 24) {real, imag} */,
  {32'hbf22e39f, 32'h00000000} /* (21, 7, 23) {real, imag} */,
  {32'hbf694daf, 32'h00000000} /* (21, 7, 22) {real, imag} */,
  {32'hbf4a53fb, 32'h00000000} /* (21, 7, 21) {real, imag} */,
  {32'h3f08d9c4, 32'h00000000} /* (21, 7, 20) {real, imag} */,
  {32'h3f89934d, 32'h00000000} /* (21, 7, 19) {real, imag} */,
  {32'h3f742d6e, 32'h00000000} /* (21, 7, 18) {real, imag} */,
  {32'h3f3fa418, 32'h00000000} /* (21, 7, 17) {real, imag} */,
  {32'h3f83d93a, 32'h00000000} /* (21, 7, 16) {real, imag} */,
  {32'h3fa37824, 32'h00000000} /* (21, 7, 15) {real, imag} */,
  {32'h3f9c1fca, 32'h00000000} /* (21, 7, 14) {real, imag} */,
  {32'h3f51d97a, 32'h00000000} /* (21, 7, 13) {real, imag} */,
  {32'h3f4107ae, 32'h00000000} /* (21, 7, 12) {real, imag} */,
  {32'h3ec3ddbe, 32'h00000000} /* (21, 7, 11) {real, imag} */,
  {32'hbd3bf28e, 32'h00000000} /* (21, 7, 10) {real, imag} */,
  {32'hbec0a6cf, 32'h00000000} /* (21, 7, 9) {real, imag} */,
  {32'hbf1fc835, 32'h00000000} /* (21, 7, 8) {real, imag} */,
  {32'hbef2b0d7, 32'h00000000} /* (21, 7, 7) {real, imag} */,
  {32'hbf651181, 32'h00000000} /* (21, 7, 6) {real, imag} */,
  {32'hbfa3c248, 32'h00000000} /* (21, 7, 5) {real, imag} */,
  {32'hbf80ce15, 32'h00000000} /* (21, 7, 4) {real, imag} */,
  {32'hbf6d3d1f, 32'h00000000} /* (21, 7, 3) {real, imag} */,
  {32'hbfab719f, 32'h00000000} /* (21, 7, 2) {real, imag} */,
  {32'hbf666b38, 32'h00000000} /* (21, 7, 1) {real, imag} */,
  {32'hbe38f9ee, 32'h00000000} /* (21, 7, 0) {real, imag} */,
  {32'hbefcddcc, 32'h00000000} /* (21, 6, 31) {real, imag} */,
  {32'hbedf8598, 32'h00000000} /* (21, 6, 30) {real, imag} */,
  {32'hbeec0fab, 32'h00000000} /* (21, 6, 29) {real, imag} */,
  {32'hbf31def5, 32'h00000000} /* (21, 6, 28) {real, imag} */,
  {32'hbf750e6e, 32'h00000000} /* (21, 6, 27) {real, imag} */,
  {32'hbf5758e4, 32'h00000000} /* (21, 6, 26) {real, imag} */,
  {32'hbf8ebe5d, 32'h00000000} /* (21, 6, 25) {real, imag} */,
  {32'hbf1baa14, 32'h00000000} /* (21, 6, 24) {real, imag} */,
  {32'hbe9c2095, 32'h00000000} /* (21, 6, 23) {real, imag} */,
  {32'hbf198eb6, 32'h00000000} /* (21, 6, 22) {real, imag} */,
  {32'hbf1cb091, 32'h00000000} /* (21, 6, 21) {real, imag} */,
  {32'h3ed21cd5, 32'h00000000} /* (21, 6, 20) {real, imag} */,
  {32'h3f63dac6, 32'h00000000} /* (21, 6, 19) {real, imag} */,
  {32'h3f9137cd, 32'h00000000} /* (21, 6, 18) {real, imag} */,
  {32'h3f3370cb, 32'h00000000} /* (21, 6, 17) {real, imag} */,
  {32'h3f844ad6, 32'h00000000} /* (21, 6, 16) {real, imag} */,
  {32'h3fd35960, 32'h00000000} /* (21, 6, 15) {real, imag} */,
  {32'h3fc75c67, 32'h00000000} /* (21, 6, 14) {real, imag} */,
  {32'h3fc680ff, 32'h00000000} /* (21, 6, 13) {real, imag} */,
  {32'h3f4491f8, 32'h00000000} /* (21, 6, 12) {real, imag} */,
  {32'h3d7feaf8, 32'h00000000} /* (21, 6, 11) {real, imag} */,
  {32'hbeb2ba5c, 32'h00000000} /* (21, 6, 10) {real, imag} */,
  {32'hbf3c2b89, 32'h00000000} /* (21, 6, 9) {real, imag} */,
  {32'hbf3eb00c, 32'h00000000} /* (21, 6, 8) {real, imag} */,
  {32'hbe39ba3f, 32'h00000000} /* (21, 6, 7) {real, imag} */,
  {32'hbf7696a1, 32'h00000000} /* (21, 6, 6) {real, imag} */,
  {32'hbf685f3f, 32'h00000000} /* (21, 6, 5) {real, imag} */,
  {32'hbf2efbac, 32'h00000000} /* (21, 6, 4) {real, imag} */,
  {32'hbf990cf1, 32'h00000000} /* (21, 6, 3) {real, imag} */,
  {32'hbf956fce, 32'h00000000} /* (21, 6, 2) {real, imag} */,
  {32'hbf340d2c, 32'h00000000} /* (21, 6, 1) {real, imag} */,
  {32'hbebc298f, 32'h00000000} /* (21, 6, 0) {real, imag} */,
  {32'hbec0e70a, 32'h00000000} /* (21, 5, 31) {real, imag} */,
  {32'hbf3cf48e, 32'h00000000} /* (21, 5, 30) {real, imag} */,
  {32'hbf42f4b2, 32'h00000000} /* (21, 5, 29) {real, imag} */,
  {32'hbf2600a1, 32'h00000000} /* (21, 5, 28) {real, imag} */,
  {32'hbf9458c4, 32'h00000000} /* (21, 5, 27) {real, imag} */,
  {32'hbfa62c86, 32'h00000000} /* (21, 5, 26) {real, imag} */,
  {32'hbf84fa49, 32'h00000000} /* (21, 5, 25) {real, imag} */,
  {32'hbf394fbe, 32'h00000000} /* (21, 5, 24) {real, imag} */,
  {32'hbeb081c4, 32'h00000000} /* (21, 5, 23) {real, imag} */,
  {32'hbf097c06, 32'h00000000} /* (21, 5, 22) {real, imag} */,
  {32'hbf8a920e, 32'h00000000} /* (21, 5, 21) {real, imag} */,
  {32'hbf285dbb, 32'h00000000} /* (21, 5, 20) {real, imag} */,
  {32'h3be159f6, 32'h00000000} /* (21, 5, 19) {real, imag} */,
  {32'h3ec634e7, 32'h00000000} /* (21, 5, 18) {real, imag} */,
  {32'hbd78c8e0, 32'h00000000} /* (21, 5, 17) {real, imag} */,
  {32'h3e6e25b0, 32'h00000000} /* (21, 5, 16) {real, imag} */,
  {32'h3f93d622, 32'h00000000} /* (21, 5, 15) {real, imag} */,
  {32'h3fbf60b9, 32'h00000000} /* (21, 5, 14) {real, imag} */,
  {32'h3faf658e, 32'h00000000} /* (21, 5, 13) {real, imag} */,
  {32'h3f2291c4, 32'h00000000} /* (21, 5, 12) {real, imag} */,
  {32'h3f43d012, 32'h00000000} /* (21, 5, 11) {real, imag} */,
  {32'h3f4b441e, 32'h00000000} /* (21, 5, 10) {real, imag} */,
  {32'h3e8e5b0a, 32'h00000000} /* (21, 5, 9) {real, imag} */,
  {32'h3f5230b0, 32'h00000000} /* (21, 5, 8) {real, imag} */,
  {32'h3f952c13, 32'h00000000} /* (21, 5, 7) {real, imag} */,
  {32'h3e04d97d, 32'h00000000} /* (21, 5, 6) {real, imag} */,
  {32'hbf104123, 32'h00000000} /* (21, 5, 5) {real, imag} */,
  {32'hbf6794e1, 32'h00000000} /* (21, 5, 4) {real, imag} */,
  {32'hbfc45419, 32'h00000000} /* (21, 5, 3) {real, imag} */,
  {32'hbf7debb7, 32'h00000000} /* (21, 5, 2) {real, imag} */,
  {32'hbf220a24, 32'h00000000} /* (21, 5, 1) {real, imag} */,
  {32'hbf007fe5, 32'h00000000} /* (21, 5, 0) {real, imag} */,
  {32'hbe127784, 32'h00000000} /* (21, 4, 31) {real, imag} */,
  {32'hbed3a1bc, 32'h00000000} /* (21, 4, 30) {real, imag} */,
  {32'hbf00a13b, 32'h00000000} /* (21, 4, 29) {real, imag} */,
  {32'hbf0b6a4b, 32'h00000000} /* (21, 4, 28) {real, imag} */,
  {32'hbf9507bb, 32'h00000000} /* (21, 4, 27) {real, imag} */,
  {32'hbfb1fa45, 32'h00000000} /* (21, 4, 26) {real, imag} */,
  {32'hbf9adb4d, 32'h00000000} /* (21, 4, 25) {real, imag} */,
  {32'hbfc9b86e, 32'h00000000} /* (21, 4, 24) {real, imag} */,
  {32'hbf533d3c, 32'h00000000} /* (21, 4, 23) {real, imag} */,
  {32'hbe5eeb0c, 32'h00000000} /* (21, 4, 22) {real, imag} */,
  {32'hbf495ffc, 32'h00000000} /* (21, 4, 21) {real, imag} */,
  {32'hbfacb46e, 32'h00000000} /* (21, 4, 20) {real, imag} */,
  {32'hbf9a3759, 32'h00000000} /* (21, 4, 19) {real, imag} */,
  {32'hbf41289a, 32'h00000000} /* (21, 4, 18) {real, imag} */,
  {32'hbf2669b3, 32'h00000000} /* (21, 4, 17) {real, imag} */,
  {32'hbf114d33, 32'h00000000} /* (21, 4, 16) {real, imag} */,
  {32'h3edf318c, 32'h00000000} /* (21, 4, 15) {real, imag} */,
  {32'h3fa8d18b, 32'h00000000} /* (21, 4, 14) {real, imag} */,
  {32'h3f8d050e, 32'h00000000} /* (21, 4, 13) {real, imag} */,
  {32'h3ee1eb1b, 32'h00000000} /* (21, 4, 12) {real, imag} */,
  {32'h3f3377ea, 32'h00000000} /* (21, 4, 11) {real, imag} */,
  {32'h3f8f3761, 32'h00000000} /* (21, 4, 10) {real, imag} */,
  {32'h3f603772, 32'h00000000} /* (21, 4, 9) {real, imag} */,
  {32'h3f811154, 32'h00000000} /* (21, 4, 8) {real, imag} */,
  {32'h3fbb1042, 32'h00000000} /* (21, 4, 7) {real, imag} */,
  {32'h3f857424, 32'h00000000} /* (21, 4, 6) {real, imag} */,
  {32'hbe426d75, 32'h00000000} /* (21, 4, 5) {real, imag} */,
  {32'hbf10e533, 32'h00000000} /* (21, 4, 4) {real, imag} */,
  {32'hbfae4ac9, 32'h00000000} /* (21, 4, 3) {real, imag} */,
  {32'hbfa94f1a, 32'h00000000} /* (21, 4, 2) {real, imag} */,
  {32'hbf4e2f77, 32'h00000000} /* (21, 4, 1) {real, imag} */,
  {32'hbf010f75, 32'h00000000} /* (21, 4, 0) {real, imag} */,
  {32'hbf084662, 32'h00000000} /* (21, 3, 31) {real, imag} */,
  {32'hbf9b6915, 32'h00000000} /* (21, 3, 30) {real, imag} */,
  {32'hbf650571, 32'h00000000} /* (21, 3, 29) {real, imag} */,
  {32'hbf6fdc59, 32'h00000000} /* (21, 3, 28) {real, imag} */,
  {32'hbf92c2e0, 32'h00000000} /* (21, 3, 27) {real, imag} */,
  {32'hbf4abf54, 32'h00000000} /* (21, 3, 26) {real, imag} */,
  {32'hbf682309, 32'h00000000} /* (21, 3, 25) {real, imag} */,
  {32'hbfa52d5a, 32'h00000000} /* (21, 3, 24) {real, imag} */,
  {32'hbf96775b, 32'h00000000} /* (21, 3, 23) {real, imag} */,
  {32'hbf51164c, 32'h00000000} /* (21, 3, 22) {real, imag} */,
  {32'hbf822e0a, 32'h00000000} /* (21, 3, 21) {real, imag} */,
  {32'hbf6f34fc, 32'h00000000} /* (21, 3, 20) {real, imag} */,
  {32'hbf586358, 32'h00000000} /* (21, 3, 19) {real, imag} */,
  {32'hbf5b28e4, 32'h00000000} /* (21, 3, 18) {real, imag} */,
  {32'hbfa953eb, 32'h00000000} /* (21, 3, 17) {real, imag} */,
  {32'hbf3a681e, 32'h00000000} /* (21, 3, 16) {real, imag} */,
  {32'h3f33df9c, 32'h00000000} /* (21, 3, 15) {real, imag} */,
  {32'h3fa68032, 32'h00000000} /* (21, 3, 14) {real, imag} */,
  {32'h3f7dff3f, 32'h00000000} /* (21, 3, 13) {real, imag} */,
  {32'h3f2410bf, 32'h00000000} /* (21, 3, 12) {real, imag} */,
  {32'h3f1cd697, 32'h00000000} /* (21, 3, 11) {real, imag} */,
  {32'h3f17c858, 32'h00000000} /* (21, 3, 10) {real, imag} */,
  {32'h3f0f6564, 32'h00000000} /* (21, 3, 9) {real, imag} */,
  {32'h3f35d487, 32'h00000000} /* (21, 3, 8) {real, imag} */,
  {32'h3fd30ca1, 32'h00000000} /* (21, 3, 7) {real, imag} */,
  {32'h3f9ae231, 32'h00000000} /* (21, 3, 6) {real, imag} */,
  {32'hbdac3d08, 32'h00000000} /* (21, 3, 5) {real, imag} */,
  {32'hbf0b05a4, 32'h00000000} /* (21, 3, 4) {real, imag} */,
  {32'hbf9ffc6a, 32'h00000000} /* (21, 3, 3) {real, imag} */,
  {32'hbfc4d1ff, 32'h00000000} /* (21, 3, 2) {real, imag} */,
  {32'hbfbb230e, 32'h00000000} /* (21, 3, 1) {real, imag} */,
  {32'hbedd7d02, 32'h00000000} /* (21, 3, 0) {real, imag} */,
  {32'hbef88e84, 32'h00000000} /* (21, 2, 31) {real, imag} */,
  {32'hbf96c10b, 32'h00000000} /* (21, 2, 30) {real, imag} */,
  {32'hbf9715e8, 32'h00000000} /* (21, 2, 29) {real, imag} */,
  {32'hbf72da8a, 32'h00000000} /* (21, 2, 28) {real, imag} */,
  {32'hbf4b3f81, 32'h00000000} /* (21, 2, 27) {real, imag} */,
  {32'hbf21cb47, 32'h00000000} /* (21, 2, 26) {real, imag} */,
  {32'hbf7a9ff8, 32'h00000000} /* (21, 2, 25) {real, imag} */,
  {32'hbf890e95, 32'h00000000} /* (21, 2, 24) {real, imag} */,
  {32'hbf9a1d4b, 32'h00000000} /* (21, 2, 23) {real, imag} */,
  {32'hbf6bbab4, 32'h00000000} /* (21, 2, 22) {real, imag} */,
  {32'hbf8bde50, 32'h00000000} /* (21, 2, 21) {real, imag} */,
  {32'hbf3de72b, 32'h00000000} /* (21, 2, 20) {real, imag} */,
  {32'hbf0e0f56, 32'h00000000} /* (21, 2, 19) {real, imag} */,
  {32'hbec26631, 32'h00000000} /* (21, 2, 18) {real, imag} */,
  {32'hbeef74ea, 32'h00000000} /* (21, 2, 17) {real, imag} */,
  {32'hbeedb20c, 32'h00000000} /* (21, 2, 16) {real, imag} */,
  {32'h3ed5f958, 32'h00000000} /* (21, 2, 15) {real, imag} */,
  {32'h3f81671d, 32'h00000000} /* (21, 2, 14) {real, imag} */,
  {32'h3f4f7856, 32'h00000000} /* (21, 2, 13) {real, imag} */,
  {32'h3f1135f1, 32'h00000000} /* (21, 2, 12) {real, imag} */,
  {32'h3edcc496, 32'h00000000} /* (21, 2, 11) {real, imag} */,
  {32'h3f09a3dd, 32'h00000000} /* (21, 2, 10) {real, imag} */,
  {32'h3f2af8d5, 32'h00000000} /* (21, 2, 9) {real, imag} */,
  {32'h3f337466, 32'h00000000} /* (21, 2, 8) {real, imag} */,
  {32'h3f73f4d2, 32'h00000000} /* (21, 2, 7) {real, imag} */,
  {32'h3f83fb78, 32'h00000000} /* (21, 2, 6) {real, imag} */,
  {32'h3e47aa8e, 32'h00000000} /* (21, 2, 5) {real, imag} */,
  {32'hbf2ddc93, 32'h00000000} /* (21, 2, 4) {real, imag} */,
  {32'hbf5d9216, 32'h00000000} /* (21, 2, 3) {real, imag} */,
  {32'hbfbc5963, 32'h00000000} /* (21, 2, 2) {real, imag} */,
  {32'hbfa6a3c4, 32'h00000000} /* (21, 2, 1) {real, imag} */,
  {32'hbe39d0b8, 32'h00000000} /* (21, 2, 0) {real, imag} */,
  {32'hbdb8c8c7, 32'h00000000} /* (21, 1, 31) {real, imag} */,
  {32'hbf06da88, 32'h00000000} /* (21, 1, 30) {real, imag} */,
  {32'hbf948b4b, 32'h00000000} /* (21, 1, 29) {real, imag} */,
  {32'hbf9b1371, 32'h00000000} /* (21, 1, 28) {real, imag} */,
  {32'hbfa0c810, 32'h00000000} /* (21, 1, 27) {real, imag} */,
  {32'hbf99ea5a, 32'h00000000} /* (21, 1, 26) {real, imag} */,
  {32'hbf851fd1, 32'h00000000} /* (21, 1, 25) {real, imag} */,
  {32'hbf994bb3, 32'h00000000} /* (21, 1, 24) {real, imag} */,
  {32'hbfcee58d, 32'h00000000} /* (21, 1, 23) {real, imag} */,
  {32'hbf93745a, 32'h00000000} /* (21, 1, 22) {real, imag} */,
  {32'hbf8889f3, 32'h00000000} /* (21, 1, 21) {real, imag} */,
  {32'hbf96f4c0, 32'h00000000} /* (21, 1, 20) {real, imag} */,
  {32'hbf3197f5, 32'h00000000} /* (21, 1, 19) {real, imag} */,
  {32'hbf038864, 32'h00000000} /* (21, 1, 18) {real, imag} */,
  {32'hbf24f676, 32'h00000000} /* (21, 1, 17) {real, imag} */,
  {32'hbf0fa761, 32'h00000000} /* (21, 1, 16) {real, imag} */,
  {32'h3eb06f02, 32'h00000000} /* (21, 1, 15) {real, imag} */,
  {32'h3f669221, 32'h00000000} /* (21, 1, 14) {real, imag} */,
  {32'h3f508164, 32'h00000000} /* (21, 1, 13) {real, imag} */,
  {32'h3f6e3869, 32'h00000000} /* (21, 1, 12) {real, imag} */,
  {32'h3f2f384c, 32'h00000000} /* (21, 1, 11) {real, imag} */,
  {32'h3f76729f, 32'h00000000} /* (21, 1, 10) {real, imag} */,
  {32'h3f74232e, 32'h00000000} /* (21, 1, 9) {real, imag} */,
  {32'h3f25b844, 32'h00000000} /* (21, 1, 8) {real, imag} */,
  {32'h3ed01be5, 32'h00000000} /* (21, 1, 7) {real, imag} */,
  {32'h3f7076e5, 32'h00000000} /* (21, 1, 6) {real, imag} */,
  {32'h3dbd2a64, 32'h00000000} /* (21, 1, 5) {real, imag} */,
  {32'hbf6da30a, 32'h00000000} /* (21, 1, 4) {real, imag} */,
  {32'hbf8e4189, 32'h00000000} /* (21, 1, 3) {real, imag} */,
  {32'hbf9dce73, 32'h00000000} /* (21, 1, 2) {real, imag} */,
  {32'hbf1c757f, 32'h00000000} /* (21, 1, 1) {real, imag} */,
  {32'hbbdca484, 32'h00000000} /* (21, 1, 0) {real, imag} */,
  {32'hbd8e3229, 32'h00000000} /* (21, 0, 31) {real, imag} */,
  {32'hbe920d00, 32'h00000000} /* (21, 0, 30) {real, imag} */,
  {32'hbeb29b52, 32'h00000000} /* (21, 0, 29) {real, imag} */,
  {32'hbf1387af, 32'h00000000} /* (21, 0, 28) {real, imag} */,
  {32'hbf8f1f92, 32'h00000000} /* (21, 0, 27) {real, imag} */,
  {32'hbf98e0c5, 32'h00000000} /* (21, 0, 26) {real, imag} */,
  {32'hbefdcdfe, 32'h00000000} /* (21, 0, 25) {real, imag} */,
  {32'hbea9d5e2, 32'h00000000} /* (21, 0, 24) {real, imag} */,
  {32'hbf2d532e, 32'h00000000} /* (21, 0, 23) {real, imag} */,
  {32'hbf0dd3ae, 32'h00000000} /* (21, 0, 22) {real, imag} */,
  {32'hbebe594d, 32'h00000000} /* (21, 0, 21) {real, imag} */,
  {32'hbf6e3a08, 32'h00000000} /* (21, 0, 20) {real, imag} */,
  {32'hbed6ba44, 32'h00000000} /* (21, 0, 19) {real, imag} */,
  {32'hbeb15476, 32'h00000000} /* (21, 0, 18) {real, imag} */,
  {32'hbf7071e4, 32'h00000000} /* (21, 0, 17) {real, imag} */,
  {32'hbed4070c, 32'h00000000} /* (21, 0, 16) {real, imag} */,
  {32'h3ec9ec8d, 32'h00000000} /* (21, 0, 15) {real, imag} */,
  {32'h3ef834fe, 32'h00000000} /* (21, 0, 14) {real, imag} */,
  {32'h3f39b29b, 32'h00000000} /* (21, 0, 13) {real, imag} */,
  {32'h3f593cf8, 32'h00000000} /* (21, 0, 12) {real, imag} */,
  {32'h3f5a6fb6, 32'h00000000} /* (21, 0, 11) {real, imag} */,
  {32'h3f3d5801, 32'h00000000} /* (21, 0, 10) {real, imag} */,
  {32'h3f0b6708, 32'h00000000} /* (21, 0, 9) {real, imag} */,
  {32'h3e48a27a, 32'h00000000} /* (21, 0, 8) {real, imag} */,
  {32'hbbf60fc9, 32'h00000000} /* (21, 0, 7) {real, imag} */,
  {32'h3defaf35, 32'h00000000} /* (21, 0, 6) {real, imag} */,
  {32'hbddbdcdd, 32'h00000000} /* (21, 0, 5) {real, imag} */,
  {32'hbef5cd5e, 32'h00000000} /* (21, 0, 4) {real, imag} */,
  {32'hbea1bcdf, 32'h00000000} /* (21, 0, 3) {real, imag} */,
  {32'hbea9463d, 32'h00000000} /* (21, 0, 2) {real, imag} */,
  {32'hbef8b948, 32'h00000000} /* (21, 0, 1) {real, imag} */,
  {32'hbe952049, 32'h00000000} /* (21, 0, 0) {real, imag} */,
  {32'hbea34767, 32'h00000000} /* (20, 31, 31) {real, imag} */,
  {32'hbf1b3a49, 32'h00000000} /* (20, 31, 30) {real, imag} */,
  {32'hbea1c77a, 32'h00000000} /* (20, 31, 29) {real, imag} */,
  {32'hbef61300, 32'h00000000} /* (20, 31, 28) {real, imag} */,
  {32'hbeed3ab8, 32'h00000000} /* (20, 31, 27) {real, imag} */,
  {32'hbf1b4590, 32'h00000000} /* (20, 31, 26) {real, imag} */,
  {32'hbf27ab71, 32'h00000000} /* (20, 31, 25) {real, imag} */,
  {32'hbeea25be, 32'h00000000} /* (20, 31, 24) {real, imag} */,
  {32'hbf122003, 32'h00000000} /* (20, 31, 23) {real, imag} */,
  {32'hbef42786, 32'h00000000} /* (20, 31, 22) {real, imag} */,
  {32'hbe59a148, 32'h00000000} /* (20, 31, 21) {real, imag} */,
  {32'h3e0a7b16, 32'h00000000} /* (20, 31, 20) {real, imag} */,
  {32'h3eec0676, 32'h00000000} /* (20, 31, 19) {real, imag} */,
  {32'h3f22930a, 32'h00000000} /* (20, 31, 18) {real, imag} */,
  {32'h3e9c2d93, 32'h00000000} /* (20, 31, 17) {real, imag} */,
  {32'h3f28ea82, 32'h00000000} /* (20, 31, 16) {real, imag} */,
  {32'h3f0386b5, 32'h00000000} /* (20, 31, 15) {real, imag} */,
  {32'h3edd568b, 32'h00000000} /* (20, 31, 14) {real, imag} */,
  {32'h3ee9b025, 32'h00000000} /* (20, 31, 13) {real, imag} */,
  {32'h3e7d06f7, 32'h00000000} /* (20, 31, 12) {real, imag} */,
  {32'h3dadd993, 32'h00000000} /* (20, 31, 11) {real, imag} */,
  {32'hbe35cde5, 32'h00000000} /* (20, 31, 10) {real, imag} */,
  {32'hbe536f2a, 32'h00000000} /* (20, 31, 9) {real, imag} */,
  {32'hbf04ded7, 32'h00000000} /* (20, 31, 8) {real, imag} */,
  {32'hbf0b5a4c, 32'h00000000} /* (20, 31, 7) {real, imag} */,
  {32'hbf0fd71b, 32'h00000000} /* (20, 31, 6) {real, imag} */,
  {32'hbf741496, 32'h00000000} /* (20, 31, 5) {real, imag} */,
  {32'hbf234c01, 32'h00000000} /* (20, 31, 4) {real, imag} */,
  {32'hbeb85028, 32'h00000000} /* (20, 31, 3) {real, imag} */,
  {32'hbea53be0, 32'h00000000} /* (20, 31, 2) {real, imag} */,
  {32'hbea8e7e5, 32'h00000000} /* (20, 31, 1) {real, imag} */,
  {32'hbe67111e, 32'h00000000} /* (20, 31, 0) {real, imag} */,
  {32'hbf156f2e, 32'h00000000} /* (20, 30, 31) {real, imag} */,
  {32'hbf78e76f, 32'h00000000} /* (20, 30, 30) {real, imag} */,
  {32'hbf5f2901, 32'h00000000} /* (20, 30, 29) {real, imag} */,
  {32'hbf9b5a07, 32'h00000000} /* (20, 30, 28) {real, imag} */,
  {32'hbf8cb1c8, 32'h00000000} /* (20, 30, 27) {real, imag} */,
  {32'hbf4873ca, 32'h00000000} /* (20, 30, 26) {real, imag} */,
  {32'hbf7fbf3e, 32'h00000000} /* (20, 30, 25) {real, imag} */,
  {32'hbf87c989, 32'h00000000} /* (20, 30, 24) {real, imag} */,
  {32'hbf85615f, 32'h00000000} /* (20, 30, 23) {real, imag} */,
  {32'hbf8ccdf4, 32'h00000000} /* (20, 30, 22) {real, imag} */,
  {32'hbee8de40, 32'h00000000} /* (20, 30, 21) {real, imag} */,
  {32'h3f06c984, 32'h00000000} /* (20, 30, 20) {real, imag} */,
  {32'h3f815f0e, 32'h00000000} /* (20, 30, 19) {real, imag} */,
  {32'h3fb76acc, 32'h00000000} /* (20, 30, 18) {real, imag} */,
  {32'h3f7c259f, 32'h00000000} /* (20, 30, 17) {real, imag} */,
  {32'h3fb38441, 32'h00000000} /* (20, 30, 16) {real, imag} */,
  {32'h3f8f7206, 32'h00000000} /* (20, 30, 15) {real, imag} */,
  {32'h3fa4bc4f, 32'h00000000} /* (20, 30, 14) {real, imag} */,
  {32'h3f75cc8b, 32'h00000000} /* (20, 30, 13) {real, imag} */,
  {32'h3ed71a70, 32'h00000000} /* (20, 30, 12) {real, imag} */,
  {32'h3e85a0e1, 32'h00000000} /* (20, 30, 11) {real, imag} */,
  {32'hbe58701c, 32'h00000000} /* (20, 30, 10) {real, imag} */,
  {32'hbeb4dd43, 32'h00000000} /* (20, 30, 9) {real, imag} */,
  {32'hbf3eb884, 32'h00000000} /* (20, 30, 8) {real, imag} */,
  {32'hbf6b70b2, 32'h00000000} /* (20, 30, 7) {real, imag} */,
  {32'hbf80c9c3, 32'h00000000} /* (20, 30, 6) {real, imag} */,
  {32'hbf8d1569, 32'h00000000} /* (20, 30, 5) {real, imag} */,
  {32'hbf8110c4, 32'h00000000} /* (20, 30, 4) {real, imag} */,
  {32'hbf6033a2, 32'h00000000} /* (20, 30, 3) {real, imag} */,
  {32'hbf0f6d6f, 32'h00000000} /* (20, 30, 2) {real, imag} */,
  {32'hbf0b41f5, 32'h00000000} /* (20, 30, 1) {real, imag} */,
  {32'hbe91514b, 32'h00000000} /* (20, 30, 0) {real, imag} */,
  {32'hbf395c25, 32'h00000000} /* (20, 29, 31) {real, imag} */,
  {32'hbf67bbb4, 32'h00000000} /* (20, 29, 30) {real, imag} */,
  {32'hbf0c91cf, 32'h00000000} /* (20, 29, 29) {real, imag} */,
  {32'hbf5b1031, 32'h00000000} /* (20, 29, 28) {real, imag} */,
  {32'hbf5f11b9, 32'h00000000} /* (20, 29, 27) {real, imag} */,
  {32'hbf853750, 32'h00000000} /* (20, 29, 26) {real, imag} */,
  {32'hbfaa47eb, 32'h00000000} /* (20, 29, 25) {real, imag} */,
  {32'hbf92b717, 32'h00000000} /* (20, 29, 24) {real, imag} */,
  {32'hbf7b607f, 32'h00000000} /* (20, 29, 23) {real, imag} */,
  {32'hbf967ae3, 32'h00000000} /* (20, 29, 22) {real, imag} */,
  {32'h3b590ba0, 32'h00000000} /* (20, 29, 21) {real, imag} */,
  {32'h3f9d68ef, 32'h00000000} /* (20, 29, 20) {real, imag} */,
  {32'h3f70f846, 32'h00000000} /* (20, 29, 19) {real, imag} */,
  {32'h3f8619f2, 32'h00000000} /* (20, 29, 18) {real, imag} */,
  {32'h3f7d8382, 32'h00000000} /* (20, 29, 17) {real, imag} */,
  {32'h3f49a6af, 32'h00000000} /* (20, 29, 16) {real, imag} */,
  {32'h3f357f0f, 32'h00000000} /* (20, 29, 15) {real, imag} */,
  {32'h3f80170d, 32'h00000000} /* (20, 29, 14) {real, imag} */,
  {32'h3f7fe0c5, 32'h00000000} /* (20, 29, 13) {real, imag} */,
  {32'h3f39ec80, 32'h00000000} /* (20, 29, 12) {real, imag} */,
  {32'h3f2fc9c4, 32'h00000000} /* (20, 29, 11) {real, imag} */,
  {32'h3e45a1f5, 32'h00000000} /* (20, 29, 10) {real, imag} */,
  {32'hbed12551, 32'h00000000} /* (20, 29, 9) {real, imag} */,
  {32'hbf3c9bf8, 32'h00000000} /* (20, 29, 8) {real, imag} */,
  {32'hbf4c4444, 32'h00000000} /* (20, 29, 7) {real, imag} */,
  {32'hbf297c6c, 32'h00000000} /* (20, 29, 6) {real, imag} */,
  {32'hbe94d2a0, 32'h00000000} /* (20, 29, 5) {real, imag} */,
  {32'hbef0e0b8, 32'h00000000} /* (20, 29, 4) {real, imag} */,
  {32'hbee226a1, 32'h00000000} /* (20, 29, 3) {real, imag} */,
  {32'hbeb7f540, 32'h00000000} /* (20, 29, 2) {real, imag} */,
  {32'hbf2b0e3c, 32'h00000000} /* (20, 29, 1) {real, imag} */,
  {32'hbf1407af, 32'h00000000} /* (20, 29, 0) {real, imag} */,
  {32'hbee0b347, 32'h00000000} /* (20, 28, 31) {real, imag} */,
  {32'hbf11de42, 32'h00000000} /* (20, 28, 30) {real, imag} */,
  {32'hbf016999, 32'h00000000} /* (20, 28, 29) {real, imag} */,
  {32'hbf8fcb67, 32'h00000000} /* (20, 28, 28) {real, imag} */,
  {32'hbf42369d, 32'h00000000} /* (20, 28, 27) {real, imag} */,
  {32'hbf568f0d, 32'h00000000} /* (20, 28, 26) {real, imag} */,
  {32'hbfb5372e, 32'h00000000} /* (20, 28, 25) {real, imag} */,
  {32'hbfdc1258, 32'h00000000} /* (20, 28, 24) {real, imag} */,
  {32'hbfbb436e, 32'h00000000} /* (20, 28, 23) {real, imag} */,
  {32'hbf99bf0a, 32'h00000000} /* (20, 28, 22) {real, imag} */,
  {32'hbe9f1f1c, 32'h00000000} /* (20, 28, 21) {real, imag} */,
  {32'h3f2f0221, 32'h00000000} /* (20, 28, 20) {real, imag} */,
  {32'h3f1009a0, 32'h00000000} /* (20, 28, 19) {real, imag} */,
  {32'h3f1d61e0, 32'h00000000} /* (20, 28, 18) {real, imag} */,
  {32'h3f3eac54, 32'h00000000} /* (20, 28, 17) {real, imag} */,
  {32'h3f67ef78, 32'h00000000} /* (20, 28, 16) {real, imag} */,
  {32'h3f88b1e7, 32'h00000000} /* (20, 28, 15) {real, imag} */,
  {32'h3f40a560, 32'h00000000} /* (20, 28, 14) {real, imag} */,
  {32'h3f23b73a, 32'h00000000} /* (20, 28, 13) {real, imag} */,
  {32'h3f944f18, 32'h00000000} /* (20, 28, 12) {real, imag} */,
  {32'h3f94f831, 32'h00000000} /* (20, 28, 11) {real, imag} */,
  {32'h3eb5277f, 32'h00000000} /* (20, 28, 10) {real, imag} */,
  {32'hbf3dac82, 32'h00000000} /* (20, 28, 9) {real, imag} */,
  {32'hbf9688b7, 32'h00000000} /* (20, 28, 8) {real, imag} */,
  {32'hbf530a27, 32'h00000000} /* (20, 28, 7) {real, imag} */,
  {32'hbf31c1c3, 32'h00000000} /* (20, 28, 6) {real, imag} */,
  {32'hbf361c68, 32'h00000000} /* (20, 28, 5) {real, imag} */,
  {32'hbf4ebaca, 32'h00000000} /* (20, 28, 4) {real, imag} */,
  {32'hbeb46e2c, 32'h00000000} /* (20, 28, 3) {real, imag} */,
  {32'hbedd3b9d, 32'h00000000} /* (20, 28, 2) {real, imag} */,
  {32'hbf66b0bf, 32'h00000000} /* (20, 28, 1) {real, imag} */,
  {32'hbf422dd9, 32'h00000000} /* (20, 28, 0) {real, imag} */,
  {32'hbf0f02d6, 32'h00000000} /* (20, 27, 31) {real, imag} */,
  {32'hbf635f1c, 32'h00000000} /* (20, 27, 30) {real, imag} */,
  {32'hbf90a4a7, 32'h00000000} /* (20, 27, 29) {real, imag} */,
  {32'hbfc88ed1, 32'h00000000} /* (20, 27, 28) {real, imag} */,
  {32'hbf6ce124, 32'h00000000} /* (20, 27, 27) {real, imag} */,
  {32'hbed837a2, 32'h00000000} /* (20, 27, 26) {real, imag} */,
  {32'hbf35fdc2, 32'h00000000} /* (20, 27, 25) {real, imag} */,
  {32'hbfd452c6, 32'h00000000} /* (20, 27, 24) {real, imag} */,
  {32'hbfce49d3, 32'h00000000} /* (20, 27, 23) {real, imag} */,
  {32'hbf381aab, 32'h00000000} /* (20, 27, 22) {real, imag} */,
  {32'hbec613fc, 32'h00000000} /* (20, 27, 21) {real, imag} */,
  {32'h3e35d68f, 32'h00000000} /* (20, 27, 20) {real, imag} */,
  {32'h3ebc24b2, 32'h00000000} /* (20, 27, 19) {real, imag} */,
  {32'h3ed1c963, 32'h00000000} /* (20, 27, 18) {real, imag} */,
  {32'h3f354bff, 32'h00000000} /* (20, 27, 17) {real, imag} */,
  {32'h3f4e6046, 32'h00000000} /* (20, 27, 16) {real, imag} */,
  {32'h3f9aa2ee, 32'h00000000} /* (20, 27, 15) {real, imag} */,
  {32'h3f79356d, 32'h00000000} /* (20, 27, 14) {real, imag} */,
  {32'h3f4053d0, 32'h00000000} /* (20, 27, 13) {real, imag} */,
  {32'h3f7f6118, 32'h00000000} /* (20, 27, 12) {real, imag} */,
  {32'h3f5455ef, 32'h00000000} /* (20, 27, 11) {real, imag} */,
  {32'hbe1cc3db, 32'h00000000} /* (20, 27, 10) {real, imag} */,
  {32'hbf6b3ef9, 32'h00000000} /* (20, 27, 9) {real, imag} */,
  {32'hbf81d181, 32'h00000000} /* (20, 27, 8) {real, imag} */,
  {32'hbf62c0e5, 32'h00000000} /* (20, 27, 7) {real, imag} */,
  {32'hbf987e13, 32'h00000000} /* (20, 27, 6) {real, imag} */,
  {32'hbfb1d503, 32'h00000000} /* (20, 27, 5) {real, imag} */,
  {32'hbf7a7c69, 32'h00000000} /* (20, 27, 4) {real, imag} */,
  {32'hbf30c0e4, 32'h00000000} /* (20, 27, 3) {real, imag} */,
  {32'hbf8449f9, 32'h00000000} /* (20, 27, 2) {real, imag} */,
  {32'hbf67ec4c, 32'h00000000} /* (20, 27, 1) {real, imag} */,
  {32'hbf00994a, 32'h00000000} /* (20, 27, 0) {real, imag} */,
  {32'hbed135bd, 32'h00000000} /* (20, 26, 31) {real, imag} */,
  {32'hbf509b99, 32'h00000000} /* (20, 26, 30) {real, imag} */,
  {32'hbf8af95b, 32'h00000000} /* (20, 26, 29) {real, imag} */,
  {32'hbfc07270, 32'h00000000} /* (20, 26, 28) {real, imag} */,
  {32'hbf6adca7, 32'h00000000} /* (20, 26, 27) {real, imag} */,
  {32'hbefb0649, 32'h00000000} /* (20, 26, 26) {real, imag} */,
  {32'hbf326d18, 32'h00000000} /* (20, 26, 25) {real, imag} */,
  {32'hbf9841cc, 32'h00000000} /* (20, 26, 24) {real, imag} */,
  {32'hbfbbf5e5, 32'h00000000} /* (20, 26, 23) {real, imag} */,
  {32'hbf8b583e, 32'h00000000} /* (20, 26, 22) {real, imag} */,
  {32'hbebed1c5, 32'h00000000} /* (20, 26, 21) {real, imag} */,
  {32'h3f0c06f2, 32'h00000000} /* (20, 26, 20) {real, imag} */,
  {32'h3f5a2430, 32'h00000000} /* (20, 26, 19) {real, imag} */,
  {32'h3f737aba, 32'h00000000} /* (20, 26, 18) {real, imag} */,
  {32'h3f3a8c5c, 32'h00000000} /* (20, 26, 17) {real, imag} */,
  {32'h3ef966c3, 32'h00000000} /* (20, 26, 16) {real, imag} */,
  {32'h3fa8c54e, 32'h00000000} /* (20, 26, 15) {real, imag} */,
  {32'h3fb4dcbb, 32'h00000000} /* (20, 26, 14) {real, imag} */,
  {32'h3fa33a83, 32'h00000000} /* (20, 26, 13) {real, imag} */,
  {32'h3faa5a07, 32'h00000000} /* (20, 26, 12) {real, imag} */,
  {32'h3f4c21e3, 32'h00000000} /* (20, 26, 11) {real, imag} */,
  {32'hbf18f84f, 32'h00000000} /* (20, 26, 10) {real, imag} */,
  {32'hbf598e4a, 32'h00000000} /* (20, 26, 9) {real, imag} */,
  {32'hbf88d0e6, 32'h00000000} /* (20, 26, 8) {real, imag} */,
  {32'hbf926262, 32'h00000000} /* (20, 26, 7) {real, imag} */,
  {32'hbf7db20f, 32'h00000000} /* (20, 26, 6) {real, imag} */,
  {32'hbf24e39f, 32'h00000000} /* (20, 26, 5) {real, imag} */,
  {32'hbef6116f, 32'h00000000} /* (20, 26, 4) {real, imag} */,
  {32'hbf2856e6, 32'h00000000} /* (20, 26, 3) {real, imag} */,
  {32'hbf72daaa, 32'h00000000} /* (20, 26, 2) {real, imag} */,
  {32'hbf6676a9, 32'h00000000} /* (20, 26, 1) {real, imag} */,
  {32'hbf22e0d2, 32'h00000000} /* (20, 26, 0) {real, imag} */,
  {32'hbf128fa2, 32'h00000000} /* (20, 25, 31) {real, imag} */,
  {32'hbf5865aa, 32'h00000000} /* (20, 25, 30) {real, imag} */,
  {32'hbf72e393, 32'h00000000} /* (20, 25, 29) {real, imag} */,
  {32'hbfa778a0, 32'h00000000} /* (20, 25, 28) {real, imag} */,
  {32'hbf9cf104, 32'h00000000} /* (20, 25, 27) {real, imag} */,
  {32'hbf5bc026, 32'h00000000} /* (20, 25, 26) {real, imag} */,
  {32'hbf4431a5, 32'h00000000} /* (20, 25, 25) {real, imag} */,
  {32'hbecbd78c, 32'h00000000} /* (20, 25, 24) {real, imag} */,
  {32'hbf449a2c, 32'h00000000} /* (20, 25, 23) {real, imag} */,
  {32'hbfaf059b, 32'h00000000} /* (20, 25, 22) {real, imag} */,
  {32'hbf1371a2, 32'h00000000} /* (20, 25, 21) {real, imag} */,
  {32'h3f553b29, 32'h00000000} /* (20, 25, 20) {real, imag} */,
  {32'h3f5e2763, 32'h00000000} /* (20, 25, 19) {real, imag} */,
  {32'h3f93b343, 32'h00000000} /* (20, 25, 18) {real, imag} */,
  {32'h3f227dee, 32'h00000000} /* (20, 25, 17) {real, imag} */,
  {32'h3e93ebb6, 32'h00000000} /* (20, 25, 16) {real, imag} */,
  {32'h3f648d0e, 32'h00000000} /* (20, 25, 15) {real, imag} */,
  {32'h3fbdede4, 32'h00000000} /* (20, 25, 14) {real, imag} */,
  {32'h3fc04a79, 32'h00000000} /* (20, 25, 13) {real, imag} */,
  {32'h3fa9fa55, 32'h00000000} /* (20, 25, 12) {real, imag} */,
  {32'h3f4dab84, 32'h00000000} /* (20, 25, 11) {real, imag} */,
  {32'hbeed8052, 32'h00000000} /* (20, 25, 10) {real, imag} */,
  {32'hbf7879a0, 32'h00000000} /* (20, 25, 9) {real, imag} */,
  {32'hbfa70dd9, 32'h00000000} /* (20, 25, 8) {real, imag} */,
  {32'hbfa25747, 32'h00000000} /* (20, 25, 7) {real, imag} */,
  {32'hbfa36f71, 32'h00000000} /* (20, 25, 6) {real, imag} */,
  {32'hbefd0fbb, 32'h00000000} /* (20, 25, 5) {real, imag} */,
  {32'hbe5b68a4, 32'h00000000} /* (20, 25, 4) {real, imag} */,
  {32'hbf10e074, 32'h00000000} /* (20, 25, 3) {real, imag} */,
  {32'hbf8dfae1, 32'h00000000} /* (20, 25, 2) {real, imag} */,
  {32'hbf460816, 32'h00000000} /* (20, 25, 1) {real, imag} */,
  {32'hbf0e1d47, 32'h00000000} /* (20, 25, 0) {real, imag} */,
  {32'hbe161b23, 32'h00000000} /* (20, 24, 31) {real, imag} */,
  {32'hbec81206, 32'h00000000} /* (20, 24, 30) {real, imag} */,
  {32'hbea8c213, 32'h00000000} /* (20, 24, 29) {real, imag} */,
  {32'hbee897b4, 32'h00000000} /* (20, 24, 28) {real, imag} */,
  {32'hbf3adeed, 32'h00000000} /* (20, 24, 27) {real, imag} */,
  {32'hbedbea4d, 32'h00000000} /* (20, 24, 26) {real, imag} */,
  {32'hbf0e2fbe, 32'h00000000} /* (20, 24, 25) {real, imag} */,
  {32'hbf50b2e6, 32'h00000000} /* (20, 24, 24) {real, imag} */,
  {32'hbf896feb, 32'h00000000} /* (20, 24, 23) {real, imag} */,
  {32'hbf6b4a45, 32'h00000000} /* (20, 24, 22) {real, imag} */,
  {32'hbee2b609, 32'h00000000} /* (20, 24, 21) {real, imag} */,
  {32'h3f71380b, 32'h00000000} /* (20, 24, 20) {real, imag} */,
  {32'h3f5761c0, 32'h00000000} /* (20, 24, 19) {real, imag} */,
  {32'h3f42affa, 32'h00000000} /* (20, 24, 18) {real, imag} */,
  {32'h3f1b319b, 32'h00000000} /* (20, 24, 17) {real, imag} */,
  {32'h3f44a2fc, 32'h00000000} /* (20, 24, 16) {real, imag} */,
  {32'h3f7eb8ed, 32'h00000000} /* (20, 24, 15) {real, imag} */,
  {32'h3f9315ce, 32'h00000000} /* (20, 24, 14) {real, imag} */,
  {32'h3f3f4b28, 32'h00000000} /* (20, 24, 13) {real, imag} */,
  {32'h3f6d8713, 32'h00000000} /* (20, 24, 12) {real, imag} */,
  {32'h3f0f5da1, 32'h00000000} /* (20, 24, 11) {real, imag} */,
  {32'hbec898c8, 32'h00000000} /* (20, 24, 10) {real, imag} */,
  {32'hbfa224a3, 32'h00000000} /* (20, 24, 9) {real, imag} */,
  {32'hbfcde926, 32'h00000000} /* (20, 24, 8) {real, imag} */,
  {32'hbf8a5cb1, 32'h00000000} /* (20, 24, 7) {real, imag} */,
  {32'hbfc2e95d, 32'h00000000} /* (20, 24, 6) {real, imag} */,
  {32'hbf246ae8, 32'h00000000} /* (20, 24, 5) {real, imag} */,
  {32'hbf103dfb, 32'h00000000} /* (20, 24, 4) {real, imag} */,
  {32'hbf94fd93, 32'h00000000} /* (20, 24, 3) {real, imag} */,
  {32'hbfa2da1f, 32'h00000000} /* (20, 24, 2) {real, imag} */,
  {32'hbf4b1569, 32'h00000000} /* (20, 24, 1) {real, imag} */,
  {32'hbee68448, 32'h00000000} /* (20, 24, 0) {real, imag} */,
  {32'hbd19301c, 32'h00000000} /* (20, 23, 31) {real, imag} */,
  {32'hbe836528, 32'h00000000} /* (20, 23, 30) {real, imag} */,
  {32'hbed03936, 32'h00000000} /* (20, 23, 29) {real, imag} */,
  {32'hbf2e869e, 32'h00000000} /* (20, 23, 28) {real, imag} */,
  {32'hbf37427a, 32'h00000000} /* (20, 23, 27) {real, imag} */,
  {32'hbecf5c8c, 32'h00000000} /* (20, 23, 26) {real, imag} */,
  {32'hbf3748dd, 32'h00000000} /* (20, 23, 25) {real, imag} */,
  {32'hbfa3c088, 32'h00000000} /* (20, 23, 24) {real, imag} */,
  {32'hbfa1b506, 32'h00000000} /* (20, 23, 23) {real, imag} */,
  {32'hbf793bb2, 32'h00000000} /* (20, 23, 22) {real, imag} */,
  {32'hbf7fdb72, 32'h00000000} /* (20, 23, 21) {real, imag} */,
  {32'h3f3df6db, 32'h00000000} /* (20, 23, 20) {real, imag} */,
  {32'h3fb20a54, 32'h00000000} /* (20, 23, 19) {real, imag} */,
  {32'h3f464693, 32'h00000000} /* (20, 23, 18) {real, imag} */,
  {32'h3ea8af4a, 32'h00000000} /* (20, 23, 17) {real, imag} */,
  {32'h3f6bca35, 32'h00000000} /* (20, 23, 16) {real, imag} */,
  {32'h3f60ce1d, 32'h00000000} /* (20, 23, 15) {real, imag} */,
  {32'h3f810856, 32'h00000000} /* (20, 23, 14) {real, imag} */,
  {32'h3f857545, 32'h00000000} /* (20, 23, 13) {real, imag} */,
  {32'h3f876563, 32'h00000000} /* (20, 23, 12) {real, imag} */,
  {32'h3ecb4611, 32'h00000000} /* (20, 23, 11) {real, imag} */,
  {32'hbf63c37b, 32'h00000000} /* (20, 23, 10) {real, imag} */,
  {32'hbf8deed3, 32'h00000000} /* (20, 23, 9) {real, imag} */,
  {32'hbf828c23, 32'h00000000} /* (20, 23, 8) {real, imag} */,
  {32'hbf53a57d, 32'h00000000} /* (20, 23, 7) {real, imag} */,
  {32'hbf8c13c1, 32'h00000000} /* (20, 23, 6) {real, imag} */,
  {32'hbf820213, 32'h00000000} /* (20, 23, 5) {real, imag} */,
  {32'hbf8bc326, 32'h00000000} /* (20, 23, 4) {real, imag} */,
  {32'hbf9bcc4a, 32'h00000000} /* (20, 23, 3) {real, imag} */,
  {32'hbf7604f0, 32'h00000000} /* (20, 23, 2) {real, imag} */,
  {32'hbf9a7cd1, 32'h00000000} /* (20, 23, 1) {real, imag} */,
  {32'hbec84651, 32'h00000000} /* (20, 23, 0) {real, imag} */,
  {32'hbe76644a, 32'h00000000} /* (20, 22, 31) {real, imag} */,
  {32'hbf15b753, 32'h00000000} /* (20, 22, 30) {real, imag} */,
  {32'hbf602365, 32'h00000000} /* (20, 22, 29) {real, imag} */,
  {32'hbf828a9c, 32'h00000000} /* (20, 22, 28) {real, imag} */,
  {32'hbf525be1, 32'h00000000} /* (20, 22, 27) {real, imag} */,
  {32'hbf30ec67, 32'h00000000} /* (20, 22, 26) {real, imag} */,
  {32'hbf577a94, 32'h00000000} /* (20, 22, 25) {real, imag} */,
  {32'hbf829a23, 32'h00000000} /* (20, 22, 24) {real, imag} */,
  {32'hbf5b9c66, 32'h00000000} /* (20, 22, 23) {real, imag} */,
  {32'hbf3639b5, 32'h00000000} /* (20, 22, 22) {real, imag} */,
  {32'hbec52d99, 32'h00000000} /* (20, 22, 21) {real, imag} */,
  {32'h3f2aa28e, 32'h00000000} /* (20, 22, 20) {real, imag} */,
  {32'h3fbbf877, 32'h00000000} /* (20, 22, 19) {real, imag} */,
  {32'h3f8490f0, 32'h00000000} /* (20, 22, 18) {real, imag} */,
  {32'h3ee9cbbe, 32'h00000000} /* (20, 22, 17) {real, imag} */,
  {32'h3f449ab7, 32'h00000000} /* (20, 22, 16) {real, imag} */,
  {32'h3f5f25a8, 32'h00000000} /* (20, 22, 15) {real, imag} */,
  {32'h3fa86fde, 32'h00000000} /* (20, 22, 14) {real, imag} */,
  {32'h3fdba216, 32'h00000000} /* (20, 22, 13) {real, imag} */,
  {32'h3fca74a5, 32'h00000000} /* (20, 22, 12) {real, imag} */,
  {32'h3f66c623, 32'h00000000} /* (20, 22, 11) {real, imag} */,
  {32'hbf32121f, 32'h00000000} /* (20, 22, 10) {real, imag} */,
  {32'hbfab7d48, 32'h00000000} /* (20, 22, 9) {real, imag} */,
  {32'hbf832639, 32'h00000000} /* (20, 22, 8) {real, imag} */,
  {32'hbf92c668, 32'h00000000} /* (20, 22, 7) {real, imag} */,
  {32'hbf5d925f, 32'h00000000} /* (20, 22, 6) {real, imag} */,
  {32'hbf31c963, 32'h00000000} /* (20, 22, 5) {real, imag} */,
  {32'hbf990115, 32'h00000000} /* (20, 22, 4) {real, imag} */,
  {32'hbf97401b, 32'h00000000} /* (20, 22, 3) {real, imag} */,
  {32'hbf7ad2c6, 32'h00000000} /* (20, 22, 2) {real, imag} */,
  {32'hbfd0aecc, 32'h00000000} /* (20, 22, 1) {real, imag} */,
  {32'hbf1e0429, 32'h00000000} /* (20, 22, 0) {real, imag} */,
  {32'hbe9a7560, 32'h00000000} /* (20, 21, 31) {real, imag} */,
  {32'hbf0543ce, 32'h00000000} /* (20, 21, 30) {real, imag} */,
  {32'hbf357741, 32'h00000000} /* (20, 21, 29) {real, imag} */,
  {32'hbf239957, 32'h00000000} /* (20, 21, 28) {real, imag} */,
  {32'hbe18ffb0, 32'h00000000} /* (20, 21, 27) {real, imag} */,
  {32'hbe921209, 32'h00000000} /* (20, 21, 26) {real, imag} */,
  {32'hbec2dc64, 32'h00000000} /* (20, 21, 25) {real, imag} */,
  {32'hbeb6ac49, 32'h00000000} /* (20, 21, 24) {real, imag} */,
  {32'hbea2afab, 32'h00000000} /* (20, 21, 23) {real, imag} */,
  {32'hbd87303c, 32'h00000000} /* (20, 21, 22) {real, imag} */,
  {32'h3ef4b67a, 32'h00000000} /* (20, 21, 21) {real, imag} */,
  {32'hbea9e31b, 32'h00000000} /* (20, 21, 20) {real, imag} */,
  {32'h3e492c13, 32'h00000000} /* (20, 21, 19) {real, imag} */,
  {32'h3ee31f15, 32'h00000000} /* (20, 21, 18) {real, imag} */,
  {32'h3e2b32ad, 32'h00000000} /* (20, 21, 17) {real, imag} */,
  {32'h3e87e14e, 32'h00000000} /* (20, 21, 16) {real, imag} */,
  {32'h3f311241, 32'h00000000} /* (20, 21, 15) {real, imag} */,
  {32'h3f9c5f48, 32'h00000000} /* (20, 21, 14) {real, imag} */,
  {32'h3f7038c2, 32'h00000000} /* (20, 21, 13) {real, imag} */,
  {32'h3f4b113a, 32'h00000000} /* (20, 21, 12) {real, imag} */,
  {32'h3f101b68, 32'h00000000} /* (20, 21, 11) {real, imag} */,
  {32'hbf2a08bf, 32'h00000000} /* (20, 21, 10) {real, imag} */,
  {32'hbf2c8539, 32'h00000000} /* (20, 21, 9) {real, imag} */,
  {32'hbe5e4620, 32'h00000000} /* (20, 21, 8) {real, imag} */,
  {32'hbf2698ff, 32'h00000000} /* (20, 21, 7) {real, imag} */,
  {32'hbe944104, 32'h00000000} /* (20, 21, 6) {real, imag} */,
  {32'h3d31af45, 32'h00000000} /* (20, 21, 5) {real, imag} */,
  {32'hbf0ced3a, 32'h00000000} /* (20, 21, 4) {real, imag} */,
  {32'hbe13e03e, 32'h00000000} /* (20, 21, 3) {real, imag} */,
  {32'hbea4fb94, 32'h00000000} /* (20, 21, 2) {real, imag} */,
  {32'hbf47eceb, 32'h00000000} /* (20, 21, 1) {real, imag} */,
  {32'hbeab00d7, 32'h00000000} /* (20, 21, 0) {real, imag} */,
  {32'h3f250956, 32'h00000000} /* (20, 20, 31) {real, imag} */,
  {32'h3f972556, 32'h00000000} /* (20, 20, 30) {real, imag} */,
  {32'h3f4ad716, 32'h00000000} /* (20, 20, 29) {real, imag} */,
  {32'h3f322945, 32'h00000000} /* (20, 20, 28) {real, imag} */,
  {32'h3f9886e8, 32'h00000000} /* (20, 20, 27) {real, imag} */,
  {32'h3f512c87, 32'h00000000} /* (20, 20, 26) {real, imag} */,
  {32'h3f09e216, 32'h00000000} /* (20, 20, 25) {real, imag} */,
  {32'h3f0638be, 32'h00000000} /* (20, 20, 24) {real, imag} */,
  {32'h3f19f082, 32'h00000000} /* (20, 20, 23) {real, imag} */,
  {32'h3f88e0fa, 32'h00000000} /* (20, 20, 22) {real, imag} */,
  {32'h3f84ac7f, 32'h00000000} /* (20, 20, 21) {real, imag} */,
  {32'hbef2f5fc, 32'h00000000} /* (20, 20, 20) {real, imag} */,
  {32'hbf58c947, 32'h00000000} /* (20, 20, 19) {real, imag} */,
  {32'hbf0b7635, 32'h00000000} /* (20, 20, 18) {real, imag} */,
  {32'hbf66c9fe, 32'h00000000} /* (20, 20, 17) {real, imag} */,
  {32'hbf41e73d, 32'h00000000} /* (20, 20, 16) {real, imag} */,
  {32'hbf2082d1, 32'h00000000} /* (20, 20, 15) {real, imag} */,
  {32'hbebda3d9, 32'h00000000} /* (20, 20, 14) {real, imag} */,
  {32'hbf35201b, 32'h00000000} /* (20, 20, 13) {real, imag} */,
  {32'hbf30d503, 32'h00000000} /* (20, 20, 12) {real, imag} */,
  {32'hbf795401, 32'h00000000} /* (20, 20, 11) {real, imag} */,
  {32'hbe8c1959, 32'h00000000} /* (20, 20, 10) {real, imag} */,
  {32'h3ee56dcb, 32'h00000000} /* (20, 20, 9) {real, imag} */,
  {32'h3e4ba454, 32'h00000000} /* (20, 20, 8) {real, imag} */,
  {32'h3d7c27cd, 32'h00000000} /* (20, 20, 7) {real, imag} */,
  {32'h3f68e769, 32'h00000000} /* (20, 20, 6) {real, imag} */,
  {32'h3f5bd12f, 32'h00000000} /* (20, 20, 5) {real, imag} */,
  {32'h3e63b324, 32'h00000000} /* (20, 20, 4) {real, imag} */,
  {32'h3f07370e, 32'h00000000} /* (20, 20, 3) {real, imag} */,
  {32'h3f1fc0e1, 32'h00000000} /* (20, 20, 2) {real, imag} */,
  {32'h3ea4e40a, 32'h00000000} /* (20, 20, 1) {real, imag} */,
  {32'h3e1d9ef1, 32'h00000000} /* (20, 20, 0) {real, imag} */,
  {32'h3f0b5bcc, 32'h00000000} /* (20, 19, 31) {real, imag} */,
  {32'h3f8ba82f, 32'h00000000} /* (20, 19, 30) {real, imag} */,
  {32'h3fb305a6, 32'h00000000} /* (20, 19, 29) {real, imag} */,
  {32'h3fb6001b, 32'h00000000} /* (20, 19, 28) {real, imag} */,
  {32'h3f969582, 32'h00000000} /* (20, 19, 27) {real, imag} */,
  {32'h3f46093c, 32'h00000000} /* (20, 19, 26) {real, imag} */,
  {32'h3f5de428, 32'h00000000} /* (20, 19, 25) {real, imag} */,
  {32'h3fb9e989, 32'h00000000} /* (20, 19, 24) {real, imag} */,
  {32'h3fce1bf8, 32'h00000000} /* (20, 19, 23) {real, imag} */,
  {32'h3f9b0dd3, 32'h00000000} /* (20, 19, 22) {real, imag} */,
  {32'h3f2e49d1, 32'h00000000} /* (20, 19, 21) {real, imag} */,
  {32'hbf293d3a, 32'h00000000} /* (20, 19, 20) {real, imag} */,
  {32'hbf89bd8f, 32'h00000000} /* (20, 19, 19) {real, imag} */,
  {32'hbf9859e9, 32'h00000000} /* (20, 19, 18) {real, imag} */,
  {32'hbfa918cb, 32'h00000000} /* (20, 19, 17) {real, imag} */,
  {32'hbfbacdbd, 32'h00000000} /* (20, 19, 16) {real, imag} */,
  {32'hbfd337a7, 32'h00000000} /* (20, 19, 15) {real, imag} */,
  {32'hbfa3e3ff, 32'h00000000} /* (20, 19, 14) {real, imag} */,
  {32'hbf8d53c7, 32'h00000000} /* (20, 19, 13) {real, imag} */,
  {32'hbf53bb34, 32'h00000000} /* (20, 19, 12) {real, imag} */,
  {32'hbf7d425c, 32'h00000000} /* (20, 19, 11) {real, imag} */,
  {32'h3d5dff19, 32'h00000000} /* (20, 19, 10) {real, imag} */,
  {32'h3f5e0348, 32'h00000000} /* (20, 19, 9) {real, imag} */,
  {32'h3eabdd1b, 32'h00000000} /* (20, 19, 8) {real, imag} */,
  {32'h3cde1018, 32'h00000000} /* (20, 19, 7) {real, imag} */,
  {32'h3ed8df15, 32'h00000000} /* (20, 19, 6) {real, imag} */,
  {32'h3eeeff1a, 32'h00000000} /* (20, 19, 5) {real, imag} */,
  {32'h3f117a20, 32'h00000000} /* (20, 19, 4) {real, imag} */,
  {32'h3f0dcccf, 32'h00000000} /* (20, 19, 3) {real, imag} */,
  {32'h3f74309b, 32'h00000000} /* (20, 19, 2) {real, imag} */,
  {32'h3faa1443, 32'h00000000} /* (20, 19, 1) {real, imag} */,
  {32'h3f59355b, 32'h00000000} /* (20, 19, 0) {real, imag} */,
  {32'h3ec16931, 32'h00000000} /* (20, 18, 31) {real, imag} */,
  {32'h3f5a7242, 32'h00000000} /* (20, 18, 30) {real, imag} */,
  {32'h3f98ab5a, 32'h00000000} /* (20, 18, 29) {real, imag} */,
  {32'h3f8ee595, 32'h00000000} /* (20, 18, 28) {real, imag} */,
  {32'h3f7ab1d0, 32'h00000000} /* (20, 18, 27) {real, imag} */,
  {32'h3f4023f9, 32'h00000000} /* (20, 18, 26) {real, imag} */,
  {32'h3f764e8e, 32'h00000000} /* (20, 18, 25) {real, imag} */,
  {32'h3fc747d5, 32'h00000000} /* (20, 18, 24) {real, imag} */,
  {32'h3fc04166, 32'h00000000} /* (20, 18, 23) {real, imag} */,
  {32'h3f68d32e, 32'h00000000} /* (20, 18, 22) {real, imag} */,
  {32'h3f6ad02b, 32'h00000000} /* (20, 18, 21) {real, imag} */,
  {32'hbe233796, 32'h00000000} /* (20, 18, 20) {real, imag} */,
  {32'hbf518218, 32'h00000000} /* (20, 18, 19) {real, imag} */,
  {32'hbf9fae3c, 32'h00000000} /* (20, 18, 18) {real, imag} */,
  {32'hbfba370d, 32'h00000000} /* (20, 18, 17) {real, imag} */,
  {32'hbff4818e, 32'h00000000} /* (20, 18, 16) {real, imag} */,
  {32'hbfcd4082, 32'h00000000} /* (20, 18, 15) {real, imag} */,
  {32'hbf71288a, 32'h00000000} /* (20, 18, 14) {real, imag} */,
  {32'hbefebb38, 32'h00000000} /* (20, 18, 13) {real, imag} */,
  {32'hbf1f6e92, 32'h00000000} /* (20, 18, 12) {real, imag} */,
  {32'hbecc22b5, 32'h00000000} /* (20, 18, 11) {real, imag} */,
  {32'h3f1cf9b0, 32'h00000000} /* (20, 18, 10) {real, imag} */,
  {32'h3f38dfcc, 32'h00000000} /* (20, 18, 9) {real, imag} */,
  {32'h3f35094e, 32'h00000000} /* (20, 18, 8) {real, imag} */,
  {32'h3ecc18cf, 32'h00000000} /* (20, 18, 7) {real, imag} */,
  {32'h3f1664af, 32'h00000000} /* (20, 18, 6) {real, imag} */,
  {32'h3fa7181e, 32'h00000000} /* (20, 18, 5) {real, imag} */,
  {32'h3fa1999f, 32'h00000000} /* (20, 18, 4) {real, imag} */,
  {32'h3f3be97e, 32'h00000000} /* (20, 18, 3) {real, imag} */,
  {32'h3f6a8928, 32'h00000000} /* (20, 18, 2) {real, imag} */,
  {32'h3fe26d66, 32'h00000000} /* (20, 18, 1) {real, imag} */,
  {32'h3fc87e58, 32'h00000000} /* (20, 18, 0) {real, imag} */,
  {32'h3ed46255, 32'h00000000} /* (20, 17, 31) {real, imag} */,
  {32'h3f31c95b, 32'h00000000} /* (20, 17, 30) {real, imag} */,
  {32'h3f7840c1, 32'h00000000} /* (20, 17, 29) {real, imag} */,
  {32'h3f99d869, 32'h00000000} /* (20, 17, 28) {real, imag} */,
  {32'h3fae1453, 32'h00000000} /* (20, 17, 27) {real, imag} */,
  {32'h3faa211f, 32'h00000000} /* (20, 17, 26) {real, imag} */,
  {32'h3f95b905, 32'h00000000} /* (20, 17, 25) {real, imag} */,
  {32'h3f9b37f1, 32'h00000000} /* (20, 17, 24) {real, imag} */,
  {32'h3f758d0e, 32'h00000000} /* (20, 17, 23) {real, imag} */,
  {32'h3f3743d7, 32'h00000000} /* (20, 17, 22) {real, imag} */,
  {32'h3eaed750, 32'h00000000} /* (20, 17, 21) {real, imag} */,
  {32'hbe4f1468, 32'h00000000} /* (20, 17, 20) {real, imag} */,
  {32'hbf5fbfc6, 32'h00000000} /* (20, 17, 19) {real, imag} */,
  {32'hbf861d5b, 32'h00000000} /* (20, 17, 18) {real, imag} */,
  {32'hbf5c7e26, 32'h00000000} /* (20, 17, 17) {real, imag} */,
  {32'hbfd941a5, 32'h00000000} /* (20, 17, 16) {real, imag} */,
  {32'hbfafb99a, 32'h00000000} /* (20, 17, 15) {real, imag} */,
  {32'hbf4a8135, 32'h00000000} /* (20, 17, 14) {real, imag} */,
  {32'hbea7ee38, 32'h00000000} /* (20, 17, 13) {real, imag} */,
  {32'hbedf405a, 32'h00000000} /* (20, 17, 12) {real, imag} */,
  {32'hbf268ec8, 32'h00000000} /* (20, 17, 11) {real, imag} */,
  {32'h3e23f51c, 32'h00000000} /* (20, 17, 10) {real, imag} */,
  {32'h3f2a5343, 32'h00000000} /* (20, 17, 9) {real, imag} */,
  {32'h3f5c1001, 32'h00000000} /* (20, 17, 8) {real, imag} */,
  {32'h3f090596, 32'h00000000} /* (20, 17, 7) {real, imag} */,
  {32'h3f3980e9, 32'h00000000} /* (20, 17, 6) {real, imag} */,
  {32'h3fcc9671, 32'h00000000} /* (20, 17, 5) {real, imag} */,
  {32'h3fd0b543, 32'h00000000} /* (20, 17, 4) {real, imag} */,
  {32'h3f7cf1d8, 32'h00000000} /* (20, 17, 3) {real, imag} */,
  {32'h3fb80f5a, 32'h00000000} /* (20, 17, 2) {real, imag} */,
  {32'h3ffca7ac, 32'h00000000} /* (20, 17, 1) {real, imag} */,
  {32'h3f84c582, 32'h00000000} /* (20, 17, 0) {real, imag} */,
  {32'h3f5c5514, 32'h00000000} /* (20, 16, 31) {real, imag} */,
  {32'h3f80ec7e, 32'h00000000} /* (20, 16, 30) {real, imag} */,
  {32'h3f761c3e, 32'h00000000} /* (20, 16, 29) {real, imag} */,
  {32'h3f985a24, 32'h00000000} /* (20, 16, 28) {real, imag} */,
  {32'h3fa38632, 32'h00000000} /* (20, 16, 27) {real, imag} */,
  {32'h3f943072, 32'h00000000} /* (20, 16, 26) {real, imag} */,
  {32'h3f9d5c06, 32'h00000000} /* (20, 16, 25) {real, imag} */,
  {32'h3f88a65b, 32'h00000000} /* (20, 16, 24) {real, imag} */,
  {32'h3f152ce9, 32'h00000000} /* (20, 16, 23) {real, imag} */,
  {32'h3ec8f178, 32'h00000000} /* (20, 16, 22) {real, imag} */,
  {32'h3c96d3d4, 32'h00000000} /* (20, 16, 21) {real, imag} */,
  {32'hbf59854a, 32'h00000000} /* (20, 16, 20) {real, imag} */,
  {32'hbf7e8995, 32'h00000000} /* (20, 16, 19) {real, imag} */,
  {32'hbf3fcdf4, 32'h00000000} /* (20, 16, 18) {real, imag} */,
  {32'hbf4f8579, 32'h00000000} /* (20, 16, 17) {real, imag} */,
  {32'hbf7b8215, 32'h00000000} /* (20, 16, 16) {real, imag} */,
  {32'hbf4cdec8, 32'h00000000} /* (20, 16, 15) {real, imag} */,
  {32'hbf796b6f, 32'h00000000} /* (20, 16, 14) {real, imag} */,
  {32'hbf8ba667, 32'h00000000} /* (20, 16, 13) {real, imag} */,
  {32'hbf7dbf55, 32'h00000000} /* (20, 16, 12) {real, imag} */,
  {32'hbf8a7fa7, 32'h00000000} /* (20, 16, 11) {real, imag} */,
  {32'h3e496fa6, 32'h00000000} /* (20, 16, 10) {real, imag} */,
  {32'h3f8b70ec, 32'h00000000} /* (20, 16, 9) {real, imag} */,
  {32'h3f77df40, 32'h00000000} /* (20, 16, 8) {real, imag} */,
  {32'h3f06a7d5, 32'h00000000} /* (20, 16, 7) {real, imag} */,
  {32'h3f3e4b97, 32'h00000000} /* (20, 16, 6) {real, imag} */,
  {32'h3faab249, 32'h00000000} /* (20, 16, 5) {real, imag} */,
  {32'h3fa51fbe, 32'h00000000} /* (20, 16, 4) {real, imag} */,
  {32'h3fadc958, 32'h00000000} /* (20, 16, 3) {real, imag} */,
  {32'h3fa364e3, 32'h00000000} /* (20, 16, 2) {real, imag} */,
  {32'h3f839805, 32'h00000000} /* (20, 16, 1) {real, imag} */,
  {32'h3f446e68, 32'h00000000} /* (20, 16, 0) {real, imag} */,
  {32'h3f923772, 32'h00000000} /* (20, 15, 31) {real, imag} */,
  {32'h3fcdb897, 32'h00000000} /* (20, 15, 30) {real, imag} */,
  {32'h3fb66d15, 32'h00000000} /* (20, 15, 29) {real, imag} */,
  {32'h3f7dd784, 32'h00000000} /* (20, 15, 28) {real, imag} */,
  {32'h3f2fa976, 32'h00000000} /* (20, 15, 27) {real, imag} */,
  {32'h3f85921e, 32'h00000000} /* (20, 15, 26) {real, imag} */,
  {32'h3f84fe76, 32'h00000000} /* (20, 15, 25) {real, imag} */,
  {32'h3f4e3297, 32'h00000000} /* (20, 15, 24) {real, imag} */,
  {32'h3f197c49, 32'h00000000} /* (20, 15, 23) {real, imag} */,
  {32'h3f3e261b, 32'h00000000} /* (20, 15, 22) {real, imag} */,
  {32'h3f28a700, 32'h00000000} /* (20, 15, 21) {real, imag} */,
  {32'hbf64844c, 32'h00000000} /* (20, 15, 20) {real, imag} */,
  {32'hbfbe87c8, 32'h00000000} /* (20, 15, 19) {real, imag} */,
  {32'hbf48dd5b, 32'h00000000} /* (20, 15, 18) {real, imag} */,
  {32'hbf68b132, 32'h00000000} /* (20, 15, 17) {real, imag} */,
  {32'hbf72cd54, 32'h00000000} /* (20, 15, 16) {real, imag} */,
  {32'hbf82507e, 32'h00000000} /* (20, 15, 15) {real, imag} */,
  {32'hbf559b2b, 32'h00000000} /* (20, 15, 14) {real, imag} */,
  {32'hbfa3cc77, 32'h00000000} /* (20, 15, 13) {real, imag} */,
  {32'hbfc4c569, 32'h00000000} /* (20, 15, 12) {real, imag} */,
  {32'hbfb8d0cf, 32'h00000000} /* (20, 15, 11) {real, imag} */,
  {32'hbddadf3d, 32'h00000000} /* (20, 15, 10) {real, imag} */,
  {32'h3f38329a, 32'h00000000} /* (20, 15, 9) {real, imag} */,
  {32'h3f39e04c, 32'h00000000} /* (20, 15, 8) {real, imag} */,
  {32'h3f478471, 32'h00000000} /* (20, 15, 7) {real, imag} */,
  {32'h3f4ca1b2, 32'h00000000} /* (20, 15, 6) {real, imag} */,
  {32'h3fabf137, 32'h00000000} /* (20, 15, 5) {real, imag} */,
  {32'h3fb7b716, 32'h00000000} /* (20, 15, 4) {real, imag} */,
  {32'h3ff23490, 32'h00000000} /* (20, 15, 3) {real, imag} */,
  {32'h3faf7b0e, 32'h00000000} /* (20, 15, 2) {real, imag} */,
  {32'h3f39ae19, 32'h00000000} /* (20, 15, 1) {real, imag} */,
  {32'h3eb84f80, 32'h00000000} /* (20, 15, 0) {real, imag} */,
  {32'h3f00f52a, 32'h00000000} /* (20, 14, 31) {real, imag} */,
  {32'h3f6a04c0, 32'h00000000} /* (20, 14, 30) {real, imag} */,
  {32'h3f8b25df, 32'h00000000} /* (20, 14, 29) {real, imag} */,
  {32'h3f8f6c44, 32'h00000000} /* (20, 14, 28) {real, imag} */,
  {32'h3f3a25d5, 32'h00000000} /* (20, 14, 27) {real, imag} */,
  {32'h3f6424a9, 32'h00000000} /* (20, 14, 26) {real, imag} */,
  {32'h3f607a2a, 32'h00000000} /* (20, 14, 25) {real, imag} */,
  {32'h3f8246b4, 32'h00000000} /* (20, 14, 24) {real, imag} */,
  {32'h3f62618f, 32'h00000000} /* (20, 14, 23) {real, imag} */,
  {32'h3f834d12, 32'h00000000} /* (20, 14, 22) {real, imag} */,
  {32'h3f3861c6, 32'h00000000} /* (20, 14, 21) {real, imag} */,
  {32'hbf6c349f, 32'h00000000} /* (20, 14, 20) {real, imag} */,
  {32'hbf737e7e, 32'h00000000} /* (20, 14, 19) {real, imag} */,
  {32'hbed74315, 32'h00000000} /* (20, 14, 18) {real, imag} */,
  {32'hbf4ca0ea, 32'h00000000} /* (20, 14, 17) {real, imag} */,
  {32'hbf6904bb, 32'h00000000} /* (20, 14, 16) {real, imag} */,
  {32'hbf901c54, 32'h00000000} /* (20, 14, 15) {real, imag} */,
  {32'hbf7871a6, 32'h00000000} /* (20, 14, 14) {real, imag} */,
  {32'hbf83b053, 32'h00000000} /* (20, 14, 13) {real, imag} */,
  {32'hbfa89348, 32'h00000000} /* (20, 14, 12) {real, imag} */,
  {32'hbf66e3e2, 32'h00000000} /* (20, 14, 11) {real, imag} */,
  {32'hbd6639a2, 32'h00000000} /* (20, 14, 10) {real, imag} */,
  {32'h3f502309, 32'h00000000} /* (20, 14, 9) {real, imag} */,
  {32'h3f9cd114, 32'h00000000} /* (20, 14, 8) {real, imag} */,
  {32'h3f74a81d, 32'h00000000} /* (20, 14, 7) {real, imag} */,
  {32'h3f5182f7, 32'h00000000} /* (20, 14, 6) {real, imag} */,
  {32'h3f651be5, 32'h00000000} /* (20, 14, 5) {real, imag} */,
  {32'h3f4520d2, 32'h00000000} /* (20, 14, 4) {real, imag} */,
  {32'h3f32e53c, 32'h00000000} /* (20, 14, 3) {real, imag} */,
  {32'h3f5f3fd4, 32'h00000000} /* (20, 14, 2) {real, imag} */,
  {32'h3f855287, 32'h00000000} /* (20, 14, 1) {real, imag} */,
  {32'h3e78394d, 32'h00000000} /* (20, 14, 0) {real, imag} */,
  {32'h3e9b7c44, 32'h00000000} /* (20, 13, 31) {real, imag} */,
  {32'h3f36af7a, 32'h00000000} /* (20, 13, 30) {real, imag} */,
  {32'h3f5d62cf, 32'h00000000} /* (20, 13, 29) {real, imag} */,
  {32'h3f88577f, 32'h00000000} /* (20, 13, 28) {real, imag} */,
  {32'h3fa916eb, 32'h00000000} /* (20, 13, 27) {real, imag} */,
  {32'h3f815b97, 32'h00000000} /* (20, 13, 26) {real, imag} */,
  {32'h3ec3d10d, 32'h00000000} /* (20, 13, 25) {real, imag} */,
  {32'h3f46d2fa, 32'h00000000} /* (20, 13, 24) {real, imag} */,
  {32'h3f7b53d6, 32'h00000000} /* (20, 13, 23) {real, imag} */,
  {32'h3f965926, 32'h00000000} /* (20, 13, 22) {real, imag} */,
  {32'h3f3b3dc1, 32'h00000000} /* (20, 13, 21) {real, imag} */,
  {32'hbf14aae2, 32'h00000000} /* (20, 13, 20) {real, imag} */,
  {32'hbf251429, 32'h00000000} /* (20, 13, 19) {real, imag} */,
  {32'hbe52e10b, 32'h00000000} /* (20, 13, 18) {real, imag} */,
  {32'hbf149cbb, 32'h00000000} /* (20, 13, 17) {real, imag} */,
  {32'hbf0766a9, 32'h00000000} /* (20, 13, 16) {real, imag} */,
  {32'hbf2cc638, 32'h00000000} /* (20, 13, 15) {real, imag} */,
  {32'hbfa4b9b3, 32'h00000000} /* (20, 13, 14) {real, imag} */,
  {32'hbfd2ebe0, 32'h00000000} /* (20, 13, 13) {real, imag} */,
  {32'hbf958091, 32'h00000000} /* (20, 13, 12) {real, imag} */,
  {32'hbf4ad9f3, 32'h00000000} /* (20, 13, 11) {real, imag} */,
  {32'h3d9cbcfb, 32'h00000000} /* (20, 13, 10) {real, imag} */,
  {32'h3f90893e, 32'h00000000} /* (20, 13, 9) {real, imag} */,
  {32'h3fc488be, 32'h00000000} /* (20, 13, 8) {real, imag} */,
  {32'h3f4bb270, 32'h00000000} /* (20, 13, 7) {real, imag} */,
  {32'h3f0c6dc9, 32'h00000000} /* (20, 13, 6) {real, imag} */,
  {32'h3f560d9d, 32'h00000000} /* (20, 13, 5) {real, imag} */,
  {32'h3f69e717, 32'h00000000} /* (20, 13, 4) {real, imag} */,
  {32'h3ef5dbf2, 32'h00000000} /* (20, 13, 3) {real, imag} */,
  {32'h3f35c02c, 32'h00000000} /* (20, 13, 2) {real, imag} */,
  {32'h3f898ae8, 32'h00000000} /* (20, 13, 1) {real, imag} */,
  {32'h3f0ea370, 32'h00000000} /* (20, 13, 0) {real, imag} */,
  {32'h3edc6182, 32'h00000000} /* (20, 12, 31) {real, imag} */,
  {32'h3f5056be, 32'h00000000} /* (20, 12, 30) {real, imag} */,
  {32'h3ebc7114, 32'h00000000} /* (20, 12, 29) {real, imag} */,
  {32'h3f08cd8d, 32'h00000000} /* (20, 12, 28) {real, imag} */,
  {32'h3f8481e5, 32'h00000000} /* (20, 12, 27) {real, imag} */,
  {32'h3f44893c, 32'h00000000} /* (20, 12, 26) {real, imag} */,
  {32'h3e11cb7a, 32'h00000000} /* (20, 12, 25) {real, imag} */,
  {32'h3e8b8a9a, 32'h00000000} /* (20, 12, 24) {real, imag} */,
  {32'h3f79ff4c, 32'h00000000} /* (20, 12, 23) {real, imag} */,
  {32'h3fb68698, 32'h00000000} /* (20, 12, 22) {real, imag} */,
  {32'h3f6da05a, 32'h00000000} /* (20, 12, 21) {real, imag} */,
  {32'hbec8d311, 32'h00000000} /* (20, 12, 20) {real, imag} */,
  {32'hbf214e11, 32'h00000000} /* (20, 12, 19) {real, imag} */,
  {32'hbf010b16, 32'h00000000} /* (20, 12, 18) {real, imag} */,
  {32'hbf223354, 32'h00000000} /* (20, 12, 17) {real, imag} */,
  {32'hbef45c18, 32'h00000000} /* (20, 12, 16) {real, imag} */,
  {32'hbf5e02e9, 32'h00000000} /* (20, 12, 15) {real, imag} */,
  {32'hbfcb4eec, 32'h00000000} /* (20, 12, 14) {real, imag} */,
  {32'hbfdb42dd, 32'h00000000} /* (20, 12, 13) {real, imag} */,
  {32'hbf35bb80, 32'h00000000} /* (20, 12, 12) {real, imag} */,
  {32'hbe986f00, 32'h00000000} /* (20, 12, 11) {real, imag} */,
  {32'h3f3169c3, 32'h00000000} /* (20, 12, 10) {real, imag} */,
  {32'h3fb26c66, 32'h00000000} /* (20, 12, 9) {real, imag} */,
  {32'h3fafc257, 32'h00000000} /* (20, 12, 8) {real, imag} */,
  {32'h3f720262, 32'h00000000} /* (20, 12, 7) {real, imag} */,
  {32'h3eb2890b, 32'h00000000} /* (20, 12, 6) {real, imag} */,
  {32'h3ee280d6, 32'h00000000} /* (20, 12, 5) {real, imag} */,
  {32'h3f825905, 32'h00000000} /* (20, 12, 4) {real, imag} */,
  {32'h3f82e07b, 32'h00000000} /* (20, 12, 3) {real, imag} */,
  {32'h3f540b3e, 32'h00000000} /* (20, 12, 2) {real, imag} */,
  {32'h3f27d26c, 32'h00000000} /* (20, 12, 1) {real, imag} */,
  {32'h3e6a4f98, 32'h00000000} /* (20, 12, 0) {real, imag} */,
  {32'h3ee585ad, 32'h00000000} /* (20, 11, 31) {real, imag} */,
  {32'h3f85f14a, 32'h00000000} /* (20, 11, 30) {real, imag} */,
  {32'h3f36d213, 32'h00000000} /* (20, 11, 29) {real, imag} */,
  {32'h3f7cb881, 32'h00000000} /* (20, 11, 28) {real, imag} */,
  {32'h3f9163cc, 32'h00000000} /* (20, 11, 27) {real, imag} */,
  {32'h3f2f33bb, 32'h00000000} /* (20, 11, 26) {real, imag} */,
  {32'h3eb8242d, 32'h00000000} /* (20, 11, 25) {real, imag} */,
  {32'h3f2244aa, 32'h00000000} /* (20, 11, 24) {real, imag} */,
  {32'h3f6fab28, 32'h00000000} /* (20, 11, 23) {real, imag} */,
  {32'h3f6f299a, 32'h00000000} /* (20, 11, 22) {real, imag} */,
  {32'h3df776d9, 32'h00000000} /* (20, 11, 21) {real, imag} */,
  {32'hbf1945dd, 32'h00000000} /* (20, 11, 20) {real, imag} */,
  {32'hbef4a85c, 32'h00000000} /* (20, 11, 19) {real, imag} */,
  {32'hbf1496d4, 32'h00000000} /* (20, 11, 18) {real, imag} */,
  {32'hbf2fce06, 32'h00000000} /* (20, 11, 17) {real, imag} */,
  {32'hbdfc5702, 32'h00000000} /* (20, 11, 16) {real, imag} */,
  {32'hbe95ceb0, 32'h00000000} /* (20, 11, 15) {real, imag} */,
  {32'hbeeb2c9a, 32'h00000000} /* (20, 11, 14) {real, imag} */,
  {32'hbed4b03c, 32'h00000000} /* (20, 11, 13) {real, imag} */,
  {32'hbf0f3cb3, 32'h00000000} /* (20, 11, 12) {real, imag} */,
  {32'h3ca3209c, 32'h00000000} /* (20, 11, 11) {real, imag} */,
  {32'h3f85b558, 32'h00000000} /* (20, 11, 10) {real, imag} */,
  {32'h3f856fcb, 32'h00000000} /* (20, 11, 9) {real, imag} */,
  {32'h3f4d9a4b, 32'h00000000} /* (20, 11, 8) {real, imag} */,
  {32'h3f4f63bb, 32'h00000000} /* (20, 11, 7) {real, imag} */,
  {32'h3f30b5a6, 32'h00000000} /* (20, 11, 6) {real, imag} */,
  {32'h3e56b110, 32'h00000000} /* (20, 11, 5) {real, imag} */,
  {32'h3e8bc73f, 32'h00000000} /* (20, 11, 4) {real, imag} */,
  {32'h3f207d23, 32'h00000000} /* (20, 11, 3) {real, imag} */,
  {32'h3f2a70a6, 32'h00000000} /* (20, 11, 2) {real, imag} */,
  {32'h3ee648b0, 32'h00000000} /* (20, 11, 1) {real, imag} */,
  {32'h3db9e063, 32'h00000000} /* (20, 11, 0) {real, imag} */,
  {32'hbd2fb992, 32'h00000000} /* (20, 10, 31) {real, imag} */,
  {32'h3d009bc7, 32'h00000000} /* (20, 10, 30) {real, imag} */,
  {32'h3cecc381, 32'h00000000} /* (20, 10, 29) {real, imag} */,
  {32'hbe088300, 32'h00000000} /* (20, 10, 28) {real, imag} */,
  {32'hbf07f9a7, 32'h00000000} /* (20, 10, 27) {real, imag} */,
  {32'hbf0c2c2d, 32'h00000000} /* (20, 10, 26) {real, imag} */,
  {32'hbe438673, 32'h00000000} /* (20, 10, 25) {real, imag} */,
  {32'hbe684616, 32'h00000000} /* (20, 10, 24) {real, imag} */,
  {32'hbeb019f7, 32'h00000000} /* (20, 10, 23) {real, imag} */,
  {32'hbf1e7800, 32'h00000000} /* (20, 10, 22) {real, imag} */,
  {32'hbe94f1dd, 32'h00000000} /* (20, 10, 21) {real, imag} */,
  {32'h3e909b7b, 32'h00000000} /* (20, 10, 20) {real, imag} */,
  {32'h3eeff3bc, 32'h00000000} /* (20, 10, 19) {real, imag} */,
  {32'h3eb4ad79, 32'h00000000} /* (20, 10, 18) {real, imag} */,
  {32'h3e73a4b5, 32'h00000000} /* (20, 10, 17) {real, imag} */,
  {32'h3f84247b, 32'h00000000} /* (20, 10, 16) {real, imag} */,
  {32'h3f811fdf, 32'h00000000} /* (20, 10, 15) {real, imag} */,
  {32'h3f09b6ba, 32'h00000000} /* (20, 10, 14) {real, imag} */,
  {32'h3e83c7de, 32'h00000000} /* (20, 10, 13) {real, imag} */,
  {32'h3e008706, 32'h00000000} /* (20, 10, 12) {real, imag} */,
  {32'h3e093331, 32'h00000000} /* (20, 10, 11) {real, imag} */,
  {32'h3e98dbce, 32'h00000000} /* (20, 10, 10) {real, imag} */,
  {32'hbf19a4e0, 32'h00000000} /* (20, 10, 9) {real, imag} */,
  {32'hbecef898, 32'h00000000} /* (20, 10, 8) {real, imag} */,
  {32'h3d91bb1e, 32'h00000000} /* (20, 10, 7) {real, imag} */,
  {32'hbf05c0d9, 32'h00000000} /* (20, 10, 6) {real, imag} */,
  {32'hbf383d51, 32'h00000000} /* (20, 10, 5) {real, imag} */,
  {32'hbf020eef, 32'h00000000} /* (20, 10, 4) {real, imag} */,
  {32'hbf3a93d5, 32'h00000000} /* (20, 10, 3) {real, imag} */,
  {32'hbf6460dc, 32'h00000000} /* (20, 10, 2) {real, imag} */,
  {32'hbe9ccbaf, 32'h00000000} /* (20, 10, 1) {real, imag} */,
  {32'hbe6b3cc8, 32'h00000000} /* (20, 10, 0) {real, imag} */,
  {32'hbeac4dc8, 32'h00000000} /* (20, 9, 31) {real, imag} */,
  {32'hbef0111f, 32'h00000000} /* (20, 9, 30) {real, imag} */,
  {32'hbefbe1ea, 32'h00000000} /* (20, 9, 29) {real, imag} */,
  {32'hbf5e9d96, 32'h00000000} /* (20, 9, 28) {real, imag} */,
  {32'hbf88ab54, 32'h00000000} /* (20, 9, 27) {real, imag} */,
  {32'hbf7fbd4e, 32'h00000000} /* (20, 9, 26) {real, imag} */,
  {32'hbf0c1f48, 32'h00000000} /* (20, 9, 25) {real, imag} */,
  {32'hbf22722a, 32'h00000000} /* (20, 9, 24) {real, imag} */,
  {32'hbf4f7ba8, 32'h00000000} /* (20, 9, 23) {real, imag} */,
  {32'hbf726e10, 32'h00000000} /* (20, 9, 22) {real, imag} */,
  {32'hbf426cbd, 32'h00000000} /* (20, 9, 21) {real, imag} */,
  {32'h3f30ec27, 32'h00000000} /* (20, 9, 20) {real, imag} */,
  {32'h3f6c0074, 32'h00000000} /* (20, 9, 19) {real, imag} */,
  {32'h3f5cb408, 32'h00000000} /* (20, 9, 18) {real, imag} */,
  {32'h3f34e8fc, 32'h00000000} /* (20, 9, 17) {real, imag} */,
  {32'h3f82694b, 32'h00000000} /* (20, 9, 16) {real, imag} */,
  {32'h3fc66077, 32'h00000000} /* (20, 9, 15) {real, imag} */,
  {32'h3fa3b002, 32'h00000000} /* (20, 9, 14) {real, imag} */,
  {32'h3f049c08, 32'h00000000} /* (20, 9, 13) {real, imag} */,
  {32'h3f1aff80, 32'h00000000} /* (20, 9, 12) {real, imag} */,
  {32'h3ec08cde, 32'h00000000} /* (20, 9, 11) {real, imag} */,
  {32'hbec2fd5b, 32'h00000000} /* (20, 9, 10) {real, imag} */,
  {32'hbfa56003, 32'h00000000} /* (20, 9, 9) {real, imag} */,
  {32'hbf8ac850, 32'h00000000} /* (20, 9, 8) {real, imag} */,
  {32'hbf364380, 32'h00000000} /* (20, 9, 7) {real, imag} */,
  {32'hbf9983ba, 32'h00000000} /* (20, 9, 6) {real, imag} */,
  {32'hbf733dec, 32'h00000000} /* (20, 9, 5) {real, imag} */,
  {32'hbf50ad81, 32'h00000000} /* (20, 9, 4) {real, imag} */,
  {32'hbf35eef3, 32'h00000000} /* (20, 9, 3) {real, imag} */,
  {32'hbf299122, 32'h00000000} /* (20, 9, 2) {real, imag} */,
  {32'hbf387816, 32'h00000000} /* (20, 9, 1) {real, imag} */,
  {32'hbf26cde0, 32'h00000000} /* (20, 9, 0) {real, imag} */,
  {32'hbf01e4ad, 32'h00000000} /* (20, 8, 31) {real, imag} */,
  {32'hbf2979ae, 32'h00000000} /* (20, 8, 30) {real, imag} */,
  {32'hbf844348, 32'h00000000} /* (20, 8, 29) {real, imag} */,
  {32'hbf6e0712, 32'h00000000} /* (20, 8, 28) {real, imag} */,
  {32'hbf4e6d2d, 32'h00000000} /* (20, 8, 27) {real, imag} */,
  {32'hbfa12f5c, 32'h00000000} /* (20, 8, 26) {real, imag} */,
  {32'hbf7c94cc, 32'h00000000} /* (20, 8, 25) {real, imag} */,
  {32'hbf168e9b, 32'h00000000} /* (20, 8, 24) {real, imag} */,
  {32'hbf79de6a, 32'h00000000} /* (20, 8, 23) {real, imag} */,
  {32'hbfcb4f01, 32'h00000000} /* (20, 8, 22) {real, imag} */,
  {32'hbfa69ab9, 32'h00000000} /* (20, 8, 21) {real, imag} */,
  {32'h3f219686, 32'h00000000} /* (20, 8, 20) {real, imag} */,
  {32'h3f94e08b, 32'h00000000} /* (20, 8, 19) {real, imag} */,
  {32'h3f12b7b1, 32'h00000000} /* (20, 8, 18) {real, imag} */,
  {32'h3ef55fee, 32'h00000000} /* (20, 8, 17) {real, imag} */,
  {32'h3f4ddeab, 32'h00000000} /* (20, 8, 16) {real, imag} */,
  {32'h3ff012d8, 32'h00000000} /* (20, 8, 15) {real, imag} */,
  {32'h3fd15495, 32'h00000000} /* (20, 8, 14) {real, imag} */,
  {32'h3f32db08, 32'h00000000} /* (20, 8, 13) {real, imag} */,
  {32'h3eebf525, 32'h00000000} /* (20, 8, 12) {real, imag} */,
  {32'h3f1f945c, 32'h00000000} /* (20, 8, 11) {real, imag} */,
  {32'hbe2b962a, 32'h00000000} /* (20, 8, 10) {real, imag} */,
  {32'hbf3b5813, 32'h00000000} /* (20, 8, 9) {real, imag} */,
  {32'hbf42bb6a, 32'h00000000} /* (20, 8, 8) {real, imag} */,
  {32'hbf2e695e, 32'h00000000} /* (20, 8, 7) {real, imag} */,
  {32'hbf7cd5be, 32'h00000000} /* (20, 8, 6) {real, imag} */,
  {32'hbf2b7b8a, 32'h00000000} /* (20, 8, 5) {real, imag} */,
  {32'hbf545847, 32'h00000000} /* (20, 8, 4) {real, imag} */,
  {32'hbf44cde2, 32'h00000000} /* (20, 8, 3) {real, imag} */,
  {32'hbf1ab5a3, 32'h00000000} /* (20, 8, 2) {real, imag} */,
  {32'hbf832f79, 32'h00000000} /* (20, 8, 1) {real, imag} */,
  {32'hbf30d1aa, 32'h00000000} /* (20, 8, 0) {real, imag} */,
  {32'hbf149447, 32'h00000000} /* (20, 7, 31) {real, imag} */,
  {32'hbf719bb5, 32'h00000000} /* (20, 7, 30) {real, imag} */,
  {32'hbfb121a2, 32'h00000000} /* (20, 7, 29) {real, imag} */,
  {32'hbf7930b5, 32'h00000000} /* (20, 7, 28) {real, imag} */,
  {32'hbf31fb84, 32'h00000000} /* (20, 7, 27) {real, imag} */,
  {32'hbf6ee08a, 32'h00000000} /* (20, 7, 26) {real, imag} */,
  {32'hbf8fc0f2, 32'h00000000} /* (20, 7, 25) {real, imag} */,
  {32'hbf9924fd, 32'h00000000} /* (20, 7, 24) {real, imag} */,
  {32'hbf6cbaf2, 32'h00000000} /* (20, 7, 23) {real, imag} */,
  {32'hbfa41008, 32'h00000000} /* (20, 7, 22) {real, imag} */,
  {32'hbf808817, 32'h00000000} /* (20, 7, 21) {real, imag} */,
  {32'h3f332d7e, 32'h00000000} /* (20, 7, 20) {real, imag} */,
  {32'h3fceccbb, 32'h00000000} /* (20, 7, 19) {real, imag} */,
  {32'h3f353ca0, 32'h00000000} /* (20, 7, 18) {real, imag} */,
  {32'h3f2280c1, 32'h00000000} /* (20, 7, 17) {real, imag} */,
  {32'h3f7e0062, 32'h00000000} /* (20, 7, 16) {real, imag} */,
  {32'h3fb8e241, 32'h00000000} /* (20, 7, 15) {real, imag} */,
  {32'h3f97ded6, 32'h00000000} /* (20, 7, 14) {real, imag} */,
  {32'h3f0cc882, 32'h00000000} /* (20, 7, 13) {real, imag} */,
  {32'h3f83bc4c, 32'h00000000} /* (20, 7, 12) {real, imag} */,
  {32'h3f076a42, 32'h00000000} /* (20, 7, 11) {real, imag} */,
  {32'hbe770372, 32'h00000000} /* (20, 7, 10) {real, imag} */,
  {32'hbee70b06, 32'h00000000} /* (20, 7, 9) {real, imag} */,
  {32'hbf19f6f1, 32'h00000000} /* (20, 7, 8) {real, imag} */,
  {32'hbf350b40, 32'h00000000} /* (20, 7, 7) {real, imag} */,
  {32'hbf3ddf6a, 32'h00000000} /* (20, 7, 6) {real, imag} */,
  {32'hbf8175de, 32'h00000000} /* (20, 7, 5) {real, imag} */,
  {32'hbf984a44, 32'h00000000} /* (20, 7, 4) {real, imag} */,
  {32'hbf8e9ee6, 32'h00000000} /* (20, 7, 3) {real, imag} */,
  {32'hbf93b3f3, 32'h00000000} /* (20, 7, 2) {real, imag} */,
  {32'hbf759a20, 32'h00000000} /* (20, 7, 1) {real, imag} */,
  {32'hbed1776a, 32'h00000000} /* (20, 7, 0) {real, imag} */,
  {32'hbf1e6413, 32'h00000000} /* (20, 6, 31) {real, imag} */,
  {32'hbf23eaa9, 32'h00000000} /* (20, 6, 30) {real, imag} */,
  {32'hbf757228, 32'h00000000} /* (20, 6, 29) {real, imag} */,
  {32'hbf808262, 32'h00000000} /* (20, 6, 28) {real, imag} */,
  {32'hbf5f4b39, 32'h00000000} /* (20, 6, 27) {real, imag} */,
  {32'hbedc30b9, 32'h00000000} /* (20, 6, 26) {real, imag} */,
  {32'hbf2adc0e, 32'h00000000} /* (20, 6, 25) {real, imag} */,
  {32'hbf622c46, 32'h00000000} /* (20, 6, 24) {real, imag} */,
  {32'hbf1bb820, 32'h00000000} /* (20, 6, 23) {real, imag} */,
  {32'hbf2cd311, 32'h00000000} /* (20, 6, 22) {real, imag} */,
  {32'hbeab2e57, 32'h00000000} /* (20, 6, 21) {real, imag} */,
  {32'h3f02850d, 32'h00000000} /* (20, 6, 20) {real, imag} */,
  {32'h3f87f96c, 32'h00000000} /* (20, 6, 19) {real, imag} */,
  {32'h3f2e618a, 32'h00000000} /* (20, 6, 18) {real, imag} */,
  {32'h3ecee641, 32'h00000000} /* (20, 6, 17) {real, imag} */,
  {32'h3f89258e, 32'h00000000} /* (20, 6, 16) {real, imag} */,
  {32'h3fbe4409, 32'h00000000} /* (20, 6, 15) {real, imag} */,
  {32'h3fa39bff, 32'h00000000} /* (20, 6, 14) {real, imag} */,
  {32'h3f89c7b7, 32'h00000000} /* (20, 6, 13) {real, imag} */,
  {32'h3fae2570, 32'h00000000} /* (20, 6, 12) {real, imag} */,
  {32'h3ed48360, 32'h00000000} /* (20, 6, 11) {real, imag} */,
  {32'hbf01395e, 32'h00000000} /* (20, 6, 10) {real, imag} */,
  {32'hbf470230, 32'h00000000} /* (20, 6, 9) {real, imag} */,
  {32'hbf531058, 32'h00000000} /* (20, 6, 8) {real, imag} */,
  {32'hbedc97e1, 32'h00000000} /* (20, 6, 7) {real, imag} */,
  {32'hbf1d25b9, 32'h00000000} /* (20, 6, 6) {real, imag} */,
  {32'hbf3d0332, 32'h00000000} /* (20, 6, 5) {real, imag} */,
  {32'hbf6f225b, 32'h00000000} /* (20, 6, 4) {real, imag} */,
  {32'hbf84c849, 32'h00000000} /* (20, 6, 3) {real, imag} */,
  {32'hbf22edd3, 32'h00000000} /* (20, 6, 2) {real, imag} */,
  {32'hbf0a8e5b, 32'h00000000} /* (20, 6, 1) {real, imag} */,
  {32'hbe9f4cc7, 32'h00000000} /* (20, 6, 0) {real, imag} */,
  {32'hbf0be42a, 32'h00000000} /* (20, 5, 31) {real, imag} */,
  {32'hbf7c08b6, 32'h00000000} /* (20, 5, 30) {real, imag} */,
  {32'hbf9e30dc, 32'h00000000} /* (20, 5, 29) {real, imag} */,
  {32'hbf379e87, 32'h00000000} /* (20, 5, 28) {real, imag} */,
  {32'hbf8f3b4a, 32'h00000000} /* (20, 5, 27) {real, imag} */,
  {32'hbf81a810, 32'h00000000} /* (20, 5, 26) {real, imag} */,
  {32'hbf2fd9c6, 32'h00000000} /* (20, 5, 25) {real, imag} */,
  {32'hbf825053, 32'h00000000} /* (20, 5, 24) {real, imag} */,
  {32'hbf339948, 32'h00000000} /* (20, 5, 23) {real, imag} */,
  {32'hbec5296b, 32'h00000000} /* (20, 5, 22) {real, imag} */,
  {32'hbe77765b, 32'h00000000} /* (20, 5, 21) {real, imag} */,
  {32'hbe3e10fe, 32'h00000000} /* (20, 5, 20) {real, imag} */,
  {32'h3dad0157, 32'h00000000} /* (20, 5, 19) {real, imag} */,
  {32'h3e2483d6, 32'h00000000} /* (20, 5, 18) {real, imag} */,
  {32'hbd1e409b, 32'h00000000} /* (20, 5, 17) {real, imag} */,
  {32'h3f2e0134, 32'h00000000} /* (20, 5, 16) {real, imag} */,
  {32'h3f7341fb, 32'h00000000} /* (20, 5, 15) {real, imag} */,
  {32'h3f752835, 32'h00000000} /* (20, 5, 14) {real, imag} */,
  {32'h3f6e2cdc, 32'h00000000} /* (20, 5, 13) {real, imag} */,
  {32'h3f7f27eb, 32'h00000000} /* (20, 5, 12) {real, imag} */,
  {32'h3f82db1c, 32'h00000000} /* (20, 5, 11) {real, imag} */,
  {32'h3eb61806, 32'h00000000} /* (20, 5, 10) {real, imag} */,
  {32'h3bc4e34b, 32'h00000000} /* (20, 5, 9) {real, imag} */,
  {32'h3eff3417, 32'h00000000} /* (20, 5, 8) {real, imag} */,
  {32'h3f563097, 32'h00000000} /* (20, 5, 7) {real, imag} */,
  {32'h3ef91501, 32'h00000000} /* (20, 5, 6) {real, imag} */,
  {32'hbec5ee57, 32'h00000000} /* (20, 5, 5) {real, imag} */,
  {32'hbf7b2836, 32'h00000000} /* (20, 5, 4) {real, imag} */,
  {32'hbfb29ad0, 32'h00000000} /* (20, 5, 3) {real, imag} */,
  {32'hbf018b7f, 32'h00000000} /* (20, 5, 2) {real, imag} */,
  {32'hbf0ad680, 32'h00000000} /* (20, 5, 1) {real, imag} */,
  {32'hbeadaf07, 32'h00000000} /* (20, 5, 0) {real, imag} */,
  {32'hbf0b26a4, 32'h00000000} /* (20, 4, 31) {real, imag} */,
  {32'hbf53c684, 32'h00000000} /* (20, 4, 30) {real, imag} */,
  {32'hbf84abd8, 32'h00000000} /* (20, 4, 29) {real, imag} */,
  {32'hbf4a5d19, 32'h00000000} /* (20, 4, 28) {real, imag} */,
  {32'hbf7ae183, 32'h00000000} /* (20, 4, 27) {real, imag} */,
  {32'hbf7a6a8e, 32'h00000000} /* (20, 4, 26) {real, imag} */,
  {32'hbf50a4da, 32'h00000000} /* (20, 4, 25) {real, imag} */,
  {32'hbfcc2834, 32'h00000000} /* (20, 4, 24) {real, imag} */,
  {32'hbf7db540, 32'h00000000} /* (20, 4, 23) {real, imag} */,
  {32'hbf0ad745, 32'h00000000} /* (20, 4, 22) {real, imag} */,
  {32'hbf167267, 32'h00000000} /* (20, 4, 21) {real, imag} */,
  {32'hbf5981e8, 32'h00000000} /* (20, 4, 20) {real, imag} */,
  {32'hbf5048eb, 32'h00000000} /* (20, 4, 19) {real, imag} */,
  {32'hbf267e11, 32'h00000000} /* (20, 4, 18) {real, imag} */,
  {32'hbede7232, 32'h00000000} /* (20, 4, 17) {real, imag} */,
  {32'hbe0c709e, 32'h00000000} /* (20, 4, 16) {real, imag} */,
  {32'h3eae6152, 32'h00000000} /* (20, 4, 15) {real, imag} */,
  {32'h3f78a34c, 32'h00000000} /* (20, 4, 14) {real, imag} */,
  {32'h3f723e3c, 32'h00000000} /* (20, 4, 13) {real, imag} */,
  {32'h3f257fcf, 32'h00000000} /* (20, 4, 12) {real, imag} */,
  {32'h3f5572e7, 32'h00000000} /* (20, 4, 11) {real, imag} */,
  {32'h3f6d410a, 32'h00000000} /* (20, 4, 10) {real, imag} */,
  {32'h3f9108f5, 32'h00000000} /* (20, 4, 9) {real, imag} */,
  {32'h3fe55c5b, 32'h00000000} /* (20, 4, 8) {real, imag} */,
  {32'h3fd9ee59, 32'h00000000} /* (20, 4, 7) {real, imag} */,
  {32'h3f8e8ec6, 32'h00000000} /* (20, 4, 6) {real, imag} */,
  {32'hbec742d4, 32'h00000000} /* (20, 4, 5) {real, imag} */,
  {32'hbf361e75, 32'h00000000} /* (20, 4, 4) {real, imag} */,
  {32'hbf8cb450, 32'h00000000} /* (20, 4, 3) {real, imag} */,
  {32'hbf5480d8, 32'h00000000} /* (20, 4, 2) {real, imag} */,
  {32'hbf1ec67f, 32'h00000000} /* (20, 4, 1) {real, imag} */,
  {32'hbee49e98, 32'h00000000} /* (20, 4, 0) {real, imag} */,
  {32'hbf092877, 32'h00000000} /* (20, 3, 31) {real, imag} */,
  {32'hbf754943, 32'h00000000} /* (20, 3, 30) {real, imag} */,
  {32'hbf707212, 32'h00000000} /* (20, 3, 29) {real, imag} */,
  {32'hbf0b57a2, 32'h00000000} /* (20, 3, 28) {real, imag} */,
  {32'hbf06f6a7, 32'h00000000} /* (20, 3, 27) {real, imag} */,
  {32'hbf2fa5b6, 32'h00000000} /* (20, 3, 26) {real, imag} */,
  {32'hbf54fbc3, 32'h00000000} /* (20, 3, 25) {real, imag} */,
  {32'hbfb84b6c, 32'h00000000} /* (20, 3, 24) {real, imag} */,
  {32'hbf94e286, 32'h00000000} /* (20, 3, 23) {real, imag} */,
  {32'hbf898f7f, 32'h00000000} /* (20, 3, 22) {real, imag} */,
  {32'hbf941b53, 32'h00000000} /* (20, 3, 21) {real, imag} */,
  {32'hbfc3a557, 32'h00000000} /* (20, 3, 20) {real, imag} */,
  {32'hbfa01c25, 32'h00000000} /* (20, 3, 19) {real, imag} */,
  {32'hbf54ec28, 32'h00000000} /* (20, 3, 18) {real, imag} */,
  {32'hbf890747, 32'h00000000} /* (20, 3, 17) {real, imag} */,
  {32'hbf2280d9, 32'h00000000} /* (20, 3, 16) {real, imag} */,
  {32'h3ed92bb2, 32'h00000000} /* (20, 3, 15) {real, imag} */,
  {32'h3f410b4f, 32'h00000000} /* (20, 3, 14) {real, imag} */,
  {32'h3f613100, 32'h00000000} /* (20, 3, 13) {real, imag} */,
  {32'h3f7f3395, 32'h00000000} /* (20, 3, 12) {real, imag} */,
  {32'h3f362ff3, 32'h00000000} /* (20, 3, 11) {real, imag} */,
  {32'h3f51eaa3, 32'h00000000} /* (20, 3, 10) {real, imag} */,
  {32'h3fb0de59, 32'h00000000} /* (20, 3, 9) {real, imag} */,
  {32'h3fb46233, 32'h00000000} /* (20, 3, 8) {real, imag} */,
  {32'h3feda9be, 32'h00000000} /* (20, 3, 7) {real, imag} */,
  {32'h3f97dfcf, 32'h00000000} /* (20, 3, 6) {real, imag} */,
  {32'hbed842f2, 32'h00000000} /* (20, 3, 5) {real, imag} */,
  {32'hbf1ec1cf, 32'h00000000} /* (20, 3, 4) {real, imag} */,
  {32'hbf7c92e2, 32'h00000000} /* (20, 3, 3) {real, imag} */,
  {32'hbf96b040, 32'h00000000} /* (20, 3, 2) {real, imag} */,
  {32'hbfa6fa9b, 32'h00000000} /* (20, 3, 1) {real, imag} */,
  {32'hbed89b19, 32'h00000000} /* (20, 3, 0) {real, imag} */,
  {32'hbed737d5, 32'h00000000} /* (20, 2, 31) {real, imag} */,
  {32'hbf8cee44, 32'h00000000} /* (20, 2, 30) {real, imag} */,
  {32'hbf683e19, 32'h00000000} /* (20, 2, 29) {real, imag} */,
  {32'hbf729665, 32'h00000000} /* (20, 2, 28) {real, imag} */,
  {32'hbf844019, 32'h00000000} /* (20, 2, 27) {real, imag} */,
  {32'hbf42a1ee, 32'h00000000} /* (20, 2, 26) {real, imag} */,
  {32'hbf50e126, 32'h00000000} /* (20, 2, 25) {real, imag} */,
  {32'hbf9ab23b, 32'h00000000} /* (20, 2, 24) {real, imag} */,
  {32'hbfc2ea72, 32'h00000000} /* (20, 2, 23) {real, imag} */,
  {32'hbf948e2d, 32'h00000000} /* (20, 2, 22) {real, imag} */,
  {32'hbf4a58b3, 32'h00000000} /* (20, 2, 21) {real, imag} */,
  {32'hbf83492c, 32'h00000000} /* (20, 2, 20) {real, imag} */,
  {32'hbf70db8e, 32'h00000000} /* (20, 2, 19) {real, imag} */,
  {32'hbf4ae7a3, 32'h00000000} /* (20, 2, 18) {real, imag} */,
  {32'hbf3c6f75, 32'h00000000} /* (20, 2, 17) {real, imag} */,
  {32'hbef1f9d7, 32'h00000000} /* (20, 2, 16) {real, imag} */,
  {32'h3edf6cf9, 32'h00000000} /* (20, 2, 15) {real, imag} */,
  {32'h3f2b172c, 32'h00000000} /* (20, 2, 14) {real, imag} */,
  {32'h3f66a3dc, 32'h00000000} /* (20, 2, 13) {real, imag} */,
  {32'h3f749f7f, 32'h00000000} /* (20, 2, 12) {real, imag} */,
  {32'h3f0381b9, 32'h00000000} /* (20, 2, 11) {real, imag} */,
  {32'h3f178f64, 32'h00000000} /* (20, 2, 10) {real, imag} */,
  {32'h3f2d9b92, 32'h00000000} /* (20, 2, 9) {real, imag} */,
  {32'h3f044e3c, 32'h00000000} /* (20, 2, 8) {real, imag} */,
  {32'h3f648319, 32'h00000000} /* (20, 2, 7) {real, imag} */,
  {32'h3f834fd8, 32'h00000000} /* (20, 2, 6) {real, imag} */,
  {32'h3e637462, 32'h00000000} /* (20, 2, 5) {real, imag} */,
  {32'hbf46fd7d, 32'h00000000} /* (20, 2, 4) {real, imag} */,
  {32'hbfa35fde, 32'h00000000} /* (20, 2, 3) {real, imag} */,
  {32'hbf8cb8f5, 32'h00000000} /* (20, 2, 2) {real, imag} */,
  {32'hbf826db4, 32'h00000000} /* (20, 2, 1) {real, imag} */,
  {32'hbe9441a7, 32'h00000000} /* (20, 2, 0) {real, imag} */,
  {32'hbda471be, 32'h00000000} /* (20, 1, 31) {real, imag} */,
  {32'hbf08e345, 32'h00000000} /* (20, 1, 30) {real, imag} */,
  {32'hbf6fdae3, 32'h00000000} /* (20, 1, 29) {real, imag} */,
  {32'hbfbea006, 32'h00000000} /* (20, 1, 28) {real, imag} */,
  {32'hbfb2159a, 32'h00000000} /* (20, 1, 27) {real, imag} */,
  {32'hbf511c45, 32'h00000000} /* (20, 1, 26) {real, imag} */,
  {32'hbf053650, 32'h00000000} /* (20, 1, 25) {real, imag} */,
  {32'hbf820d8d, 32'h00000000} /* (20, 1, 24) {real, imag} */,
  {32'hbfac682f, 32'h00000000} /* (20, 1, 23) {real, imag} */,
  {32'hbf156d4c, 32'h00000000} /* (20, 1, 22) {real, imag} */,
  {32'hbedb3b72, 32'h00000000} /* (20, 1, 21) {real, imag} */,
  {32'hbf2882dd, 32'h00000000} /* (20, 1, 20) {real, imag} */,
  {32'hbf1dd175, 32'h00000000} /* (20, 1, 19) {real, imag} */,
  {32'hbf6a6615, 32'h00000000} /* (20, 1, 18) {real, imag} */,
  {32'hbf56860e, 32'h00000000} /* (20, 1, 17) {real, imag} */,
  {32'h3d890ec9, 32'h00000000} /* (20, 1, 16) {real, imag} */,
  {32'h3f5b8b64, 32'h00000000} /* (20, 1, 15) {real, imag} */,
  {32'h3f16b145, 32'h00000000} /* (20, 1, 14) {real, imag} */,
  {32'h3f032710, 32'h00000000} /* (20, 1, 13) {real, imag} */,
  {32'h3f78719a, 32'h00000000} /* (20, 1, 12) {real, imag} */,
  {32'h3f5c021f, 32'h00000000} /* (20, 1, 11) {real, imag} */,
  {32'h3f580fa3, 32'h00000000} /* (20, 1, 10) {real, imag} */,
  {32'h3f89d003, 32'h00000000} /* (20, 1, 9) {real, imag} */,
  {32'h3f3116e3, 32'h00000000} /* (20, 1, 8) {real, imag} */,
  {32'h3f15a092, 32'h00000000} /* (20, 1, 7) {real, imag} */,
  {32'h3f9bd79a, 32'h00000000} /* (20, 1, 6) {real, imag} */,
  {32'h3e804ebe, 32'h00000000} /* (20, 1, 5) {real, imag} */,
  {32'hbf9ddb23, 32'h00000000} /* (20, 1, 4) {real, imag} */,
  {32'hbfabf30f, 32'h00000000} /* (20, 1, 3) {real, imag} */,
  {32'hbf266a95, 32'h00000000} /* (20, 1, 2) {real, imag} */,
  {32'hbf20d975, 32'h00000000} /* (20, 1, 1) {real, imag} */,
  {32'hbec0d5df, 32'h00000000} /* (20, 1, 0) {real, imag} */,
  {32'hbdd774ff, 32'h00000000} /* (20, 0, 31) {real, imag} */,
  {32'hbe71161d, 32'h00000000} /* (20, 0, 30) {real, imag} */,
  {32'hbeab6830, 32'h00000000} /* (20, 0, 29) {real, imag} */,
  {32'hbf560962, 32'h00000000} /* (20, 0, 28) {real, imag} */,
  {32'hbf5819d4, 32'h00000000} /* (20, 0, 27) {real, imag} */,
  {32'hbf169b88, 32'h00000000} /* (20, 0, 26) {real, imag} */,
  {32'hbec9cce7, 32'h00000000} /* (20, 0, 25) {real, imag} */,
  {32'hbe8c6c0d, 32'h00000000} /* (20, 0, 24) {real, imag} */,
  {32'hbeb4a65c, 32'h00000000} /* (20, 0, 23) {real, imag} */,
  {32'hbdeaa106, 32'h00000000} /* (20, 0, 22) {real, imag} */,
  {32'hbe257d16, 32'h00000000} /* (20, 0, 21) {real, imag} */,
  {32'hbe9d04c0, 32'h00000000} /* (20, 0, 20) {real, imag} */,
  {32'hbe3e33cc, 32'h00000000} /* (20, 0, 19) {real, imag} */,
  {32'hbe82ff91, 32'h00000000} /* (20, 0, 18) {real, imag} */,
  {32'hbf17d209, 32'h00000000} /* (20, 0, 17) {real, imag} */,
  {32'h3e09b418, 32'h00000000} /* (20, 0, 16) {real, imag} */,
  {32'h3f38bd3e, 32'h00000000} /* (20, 0, 15) {real, imag} */,
  {32'h3e890598, 32'h00000000} /* (20, 0, 14) {real, imag} */,
  {32'h3eae381f, 32'h00000000} /* (20, 0, 13) {real, imag} */,
  {32'h3f39cd15, 32'h00000000} /* (20, 0, 12) {real, imag} */,
  {32'h3f4a9948, 32'h00000000} /* (20, 0, 11) {real, imag} */,
  {32'h3f122840, 32'h00000000} /* (20, 0, 10) {real, imag} */,
  {32'h3f3c4457, 32'h00000000} /* (20, 0, 9) {real, imag} */,
  {32'h3f014181, 32'h00000000} /* (20, 0, 8) {real, imag} */,
  {32'h3e8822ec, 32'h00000000} /* (20, 0, 7) {real, imag} */,
  {32'h3eb1a8a1, 32'h00000000} /* (20, 0, 6) {real, imag} */,
  {32'hbe403cc6, 32'h00000000} /* (20, 0, 5) {real, imag} */,
  {32'hbf0702e3, 32'h00000000} /* (20, 0, 4) {real, imag} */,
  {32'hbeb901f7, 32'h00000000} /* (20, 0, 3) {real, imag} */,
  {32'hbdf31fd3, 32'h00000000} /* (20, 0, 2) {real, imag} */,
  {32'hbf160a9d, 32'h00000000} /* (20, 0, 1) {real, imag} */,
  {32'hbf374dd8, 32'h00000000} /* (20, 0, 0) {real, imag} */,
  {32'hbf1e9364, 32'h00000000} /* (19, 31, 31) {real, imag} */,
  {32'hbf6ce0c0, 32'h00000000} /* (19, 31, 30) {real, imag} */,
  {32'hbf0953e7, 32'h00000000} /* (19, 31, 29) {real, imag} */,
  {32'hbf1a471b, 32'h00000000} /* (19, 31, 28) {real, imag} */,
  {32'hbf61e6a0, 32'h00000000} /* (19, 31, 27) {real, imag} */,
  {32'hbf79b4ea, 32'h00000000} /* (19, 31, 26) {real, imag} */,
  {32'hbecb0bac, 32'h00000000} /* (19, 31, 25) {real, imag} */,
  {32'hbe3f5444, 32'h00000000} /* (19, 31, 24) {real, imag} */,
  {32'hbeb89470, 32'h00000000} /* (19, 31, 23) {real, imag} */,
  {32'hbea1eb38, 32'h00000000} /* (19, 31, 22) {real, imag} */,
  {32'hbe39d873, 32'h00000000} /* (19, 31, 21) {real, imag} */,
  {32'h3d984700, 32'h00000000} /* (19, 31, 20) {real, imag} */,
  {32'h3ec38527, 32'h00000000} /* (19, 31, 19) {real, imag} */,
  {32'h3f5715d4, 32'h00000000} /* (19, 31, 18) {real, imag} */,
  {32'h3f0c508a, 32'h00000000} /* (19, 31, 17) {real, imag} */,
  {32'h3f094203, 32'h00000000} /* (19, 31, 16) {real, imag} */,
  {32'h3f1723b5, 32'h00000000} /* (19, 31, 15) {real, imag} */,
  {32'h3ea8a365, 32'h00000000} /* (19, 31, 14) {real, imag} */,
  {32'h3e57f131, 32'h00000000} /* (19, 31, 13) {real, imag} */,
  {32'h3ec1d293, 32'h00000000} /* (19, 31, 12) {real, imag} */,
  {32'h3eb86b1d, 32'h00000000} /* (19, 31, 11) {real, imag} */,
  {32'hbe370404, 32'h00000000} /* (19, 31, 10) {real, imag} */,
  {32'hbec98462, 32'h00000000} /* (19, 31, 9) {real, imag} */,
  {32'hbf0eff13, 32'h00000000} /* (19, 31, 8) {real, imag} */,
  {32'hbea9d5d5, 32'h00000000} /* (19, 31, 7) {real, imag} */,
  {32'hbeeaf7e7, 32'h00000000} /* (19, 31, 6) {real, imag} */,
  {32'hbf6c91f2, 32'h00000000} /* (19, 31, 5) {real, imag} */,
  {32'hbf11d93b, 32'h00000000} /* (19, 31, 4) {real, imag} */,
  {32'hbf08825c, 32'h00000000} /* (19, 31, 3) {real, imag} */,
  {32'hbf39244e, 32'h00000000} /* (19, 31, 2) {real, imag} */,
  {32'hbf4ba810, 32'h00000000} /* (19, 31, 1) {real, imag} */,
  {32'hbef995fb, 32'h00000000} /* (19, 31, 0) {real, imag} */,
  {32'hbf17100b, 32'h00000000} /* (19, 30, 31) {real, imag} */,
  {32'hbf9352e8, 32'h00000000} /* (19, 30, 30) {real, imag} */,
  {32'hbf774b26, 32'h00000000} /* (19, 30, 29) {real, imag} */,
  {32'hbf47ced9, 32'h00000000} /* (19, 30, 28) {real, imag} */,
  {32'hbfa6b9a1, 32'h00000000} /* (19, 30, 27) {real, imag} */,
  {32'hbfd92d8a, 32'h00000000} /* (19, 30, 26) {real, imag} */,
  {32'hbf2b8b80, 32'h00000000} /* (19, 30, 25) {real, imag} */,
  {32'hbf267112, 32'h00000000} /* (19, 30, 24) {real, imag} */,
  {32'hbf64bf44, 32'h00000000} /* (19, 30, 23) {real, imag} */,
  {32'hbf36d66c, 32'h00000000} /* (19, 30, 22) {real, imag} */,
  {32'hbec858db, 32'h00000000} /* (19, 30, 21) {real, imag} */,
  {32'h3f138292, 32'h00000000} /* (19, 30, 20) {real, imag} */,
  {32'h3f2187cf, 32'h00000000} /* (19, 30, 19) {real, imag} */,
  {32'h3f999e2d, 32'h00000000} /* (19, 30, 18) {real, imag} */,
  {32'h3fa59248, 32'h00000000} /* (19, 30, 17) {real, imag} */,
  {32'h3faf2dcc, 32'h00000000} /* (19, 30, 16) {real, imag} */,
  {32'h3f8fc68b, 32'h00000000} /* (19, 30, 15) {real, imag} */,
  {32'h3f9f457a, 32'h00000000} /* (19, 30, 14) {real, imag} */,
  {32'h3f660b34, 32'h00000000} /* (19, 30, 13) {real, imag} */,
  {32'h3f01c211, 32'h00000000} /* (19, 30, 12) {real, imag} */,
  {32'h3f12a5dc, 32'h00000000} /* (19, 30, 11) {real, imag} */,
  {32'h3e7bb404, 32'h00000000} /* (19, 30, 10) {real, imag} */,
  {32'hbf1e6cb1, 32'h00000000} /* (19, 30, 9) {real, imag} */,
  {32'hbf80e79f, 32'h00000000} /* (19, 30, 8) {real, imag} */,
  {32'hbf82da3e, 32'h00000000} /* (19, 30, 7) {real, imag} */,
  {32'hbf575067, 32'h00000000} /* (19, 30, 6) {real, imag} */,
  {32'hbf728dc4, 32'h00000000} /* (19, 30, 5) {real, imag} */,
  {32'hbf87347c, 32'h00000000} /* (19, 30, 4) {real, imag} */,
  {32'hbf84b775, 32'h00000000} /* (19, 30, 3) {real, imag} */,
  {32'hbf62a806, 32'h00000000} /* (19, 30, 2) {real, imag} */,
  {32'hbf490948, 32'h00000000} /* (19, 30, 1) {real, imag} */,
  {32'hbea4e4eb, 32'h00000000} /* (19, 30, 0) {real, imag} */,
  {32'hbf25e9cd, 32'h00000000} /* (19, 29, 31) {real, imag} */,
  {32'hbf310644, 32'h00000000} /* (19, 29, 30) {real, imag} */,
  {32'hbf09dabf, 32'h00000000} /* (19, 29, 29) {real, imag} */,
  {32'hbf1e8677, 32'h00000000} /* (19, 29, 28) {real, imag} */,
  {32'hbf1abb52, 32'h00000000} /* (19, 29, 27) {real, imag} */,
  {32'hbf66a570, 32'h00000000} /* (19, 29, 26) {real, imag} */,
  {32'hbf479a3a, 32'h00000000} /* (19, 29, 25) {real, imag} */,
  {32'hbfa23dc3, 32'h00000000} /* (19, 29, 24) {real, imag} */,
  {32'hbfab33cb, 32'h00000000} /* (19, 29, 23) {real, imag} */,
  {32'hbf54b7a3, 32'h00000000} /* (19, 29, 22) {real, imag} */,
  {32'h3e61fde0, 32'h00000000} /* (19, 29, 21) {real, imag} */,
  {32'h3fcd2d79, 32'h00000000} /* (19, 29, 20) {real, imag} */,
  {32'h3f4599b6, 32'h00000000} /* (19, 29, 19) {real, imag} */,
  {32'h3f8d6f00, 32'h00000000} /* (19, 29, 18) {real, imag} */,
  {32'h3fa8607c, 32'h00000000} /* (19, 29, 17) {real, imag} */,
  {32'h3f85bc10, 32'h00000000} /* (19, 29, 16) {real, imag} */,
  {32'h3f37e18e, 32'h00000000} /* (19, 29, 15) {real, imag} */,
  {32'h3f8f304d, 32'h00000000} /* (19, 29, 14) {real, imag} */,
  {32'h3f9e3022, 32'h00000000} /* (19, 29, 13) {real, imag} */,
  {32'h3f397912, 32'h00000000} /* (19, 29, 12) {real, imag} */,
  {32'h3ef9c788, 32'h00000000} /* (19, 29, 11) {real, imag} */,
  {32'h3e21c7f0, 32'h00000000} /* (19, 29, 10) {real, imag} */,
  {32'hbefe2d62, 32'h00000000} /* (19, 29, 9) {real, imag} */,
  {32'hbf83ddc0, 32'h00000000} /* (19, 29, 8) {real, imag} */,
  {32'hbf8ee679, 32'h00000000} /* (19, 29, 7) {real, imag} */,
  {32'hbf4e0324, 32'h00000000} /* (19, 29, 6) {real, imag} */,
  {32'hbf372434, 32'h00000000} /* (19, 29, 5) {real, imag} */,
  {32'hbf472ecd, 32'h00000000} /* (19, 29, 4) {real, imag} */,
  {32'hbf716abe, 32'h00000000} /* (19, 29, 3) {real, imag} */,
  {32'hbf2c3718, 32'h00000000} /* (19, 29, 2) {real, imag} */,
  {32'hbf732c6f, 32'h00000000} /* (19, 29, 1) {real, imag} */,
  {32'hbf347c7a, 32'h00000000} /* (19, 29, 0) {real, imag} */,
  {32'hbeddbac7, 32'h00000000} /* (19, 28, 31) {real, imag} */,
  {32'hbf136725, 32'h00000000} /* (19, 28, 30) {real, imag} */,
  {32'hbf684334, 32'h00000000} /* (19, 28, 29) {real, imag} */,
  {32'hbfb72a87, 32'h00000000} /* (19, 28, 28) {real, imag} */,
  {32'hbf2aee52, 32'h00000000} /* (19, 28, 27) {real, imag} */,
  {32'hbf5b11e5, 32'h00000000} /* (19, 28, 26) {real, imag} */,
  {32'hbfbec045, 32'h00000000} /* (19, 28, 25) {real, imag} */,
  {32'hc0107f2d, 32'h00000000} /* (19, 28, 24) {real, imag} */,
  {32'hbfbb4432, 32'h00000000} /* (19, 28, 23) {real, imag} */,
  {32'hbf40b6d3, 32'h00000000} /* (19, 28, 22) {real, imag} */,
  {32'h3e1decef, 32'h00000000} /* (19, 28, 21) {real, imag} */,
  {32'h3fd07586, 32'h00000000} /* (19, 28, 20) {real, imag} */,
  {32'h3f795de7, 32'h00000000} /* (19, 28, 19) {real, imag} */,
  {32'h3f8ad46d, 32'h00000000} /* (19, 28, 18) {real, imag} */,
  {32'h3f935d1d, 32'h00000000} /* (19, 28, 17) {real, imag} */,
  {32'h3f9f9ab2, 32'h00000000} /* (19, 28, 16) {real, imag} */,
  {32'h3f62f118, 32'h00000000} /* (19, 28, 15) {real, imag} */,
  {32'h3f69810f, 32'h00000000} /* (19, 28, 14) {real, imag} */,
  {32'h3f6429cb, 32'h00000000} /* (19, 28, 13) {real, imag} */,
  {32'h3f3c2ccd, 32'h00000000} /* (19, 28, 12) {real, imag} */,
  {32'h3f19a11a, 32'h00000000} /* (19, 28, 11) {real, imag} */,
  {32'hbd1ff73f, 32'h00000000} /* (19, 28, 10) {real, imag} */,
  {32'hbf1420bd, 32'h00000000} /* (19, 28, 9) {real, imag} */,
  {32'hbf216941, 32'h00000000} /* (19, 28, 8) {real, imag} */,
  {32'hbf148da2, 32'h00000000} /* (19, 28, 7) {real, imag} */,
  {32'hbf4a944f, 32'h00000000} /* (19, 28, 6) {real, imag} */,
  {32'hbf3712a8, 32'h00000000} /* (19, 28, 5) {real, imag} */,
  {32'hbf2d8c1e, 32'h00000000} /* (19, 28, 4) {real, imag} */,
  {32'hbf33591c, 32'h00000000} /* (19, 28, 3) {real, imag} */,
  {32'hbf451f34, 32'h00000000} /* (19, 28, 2) {real, imag} */,
  {32'hbf8d1ae1, 32'h00000000} /* (19, 28, 1) {real, imag} */,
  {32'hbf304104, 32'h00000000} /* (19, 28, 0) {real, imag} */,
  {32'hbf2e4e28, 32'h00000000} /* (19, 27, 31) {real, imag} */,
  {32'hbf7d0c5c, 32'h00000000} /* (19, 27, 30) {real, imag} */,
  {32'hbf79d56f, 32'h00000000} /* (19, 27, 29) {real, imag} */,
  {32'hbf5504a8, 32'h00000000} /* (19, 27, 28) {real, imag} */,
  {32'hbebc86ee, 32'h00000000} /* (19, 27, 27) {real, imag} */,
  {32'hbf42e9de, 32'h00000000} /* (19, 27, 26) {real, imag} */,
  {32'hbfdc0bc1, 32'h00000000} /* (19, 27, 25) {real, imag} */,
  {32'hbfdd66ea, 32'h00000000} /* (19, 27, 24) {real, imag} */,
  {32'hbf8b3ba8, 32'h00000000} /* (19, 27, 23) {real, imag} */,
  {32'hbe875998, 32'h00000000} /* (19, 27, 22) {real, imag} */,
  {32'hbd2d6b3c, 32'h00000000} /* (19, 27, 21) {real, imag} */,
  {32'h3f36340c, 32'h00000000} /* (19, 27, 20) {real, imag} */,
  {32'h3f2a7e37, 32'h00000000} /* (19, 27, 19) {real, imag} */,
  {32'h3f04ea4f, 32'h00000000} /* (19, 27, 18) {real, imag} */,
  {32'h3f7b0508, 32'h00000000} /* (19, 27, 17) {real, imag} */,
  {32'h3f8aa13c, 32'h00000000} /* (19, 27, 16) {real, imag} */,
  {32'h3f9b92bd, 32'h00000000} /* (19, 27, 15) {real, imag} */,
  {32'h3faa4f50, 32'h00000000} /* (19, 27, 14) {real, imag} */,
  {32'h3f550b62, 32'h00000000} /* (19, 27, 13) {real, imag} */,
  {32'h3f123ca1, 32'h00000000} /* (19, 27, 12) {real, imag} */,
  {32'h3e51e54f, 32'h00000000} /* (19, 27, 11) {real, imag} */,
  {32'hbef1c813, 32'h00000000} /* (19, 27, 10) {real, imag} */,
  {32'hbf9a3650, 32'h00000000} /* (19, 27, 9) {real, imag} */,
  {32'hbf614d35, 32'h00000000} /* (19, 27, 8) {real, imag} */,
  {32'hbf1a9a1c, 32'h00000000} /* (19, 27, 7) {real, imag} */,
  {32'hbf7e7232, 32'h00000000} /* (19, 27, 6) {real, imag} */,
  {32'hbfa8a171, 32'h00000000} /* (19, 27, 5) {real, imag} */,
  {32'hbf8902c2, 32'h00000000} /* (19, 27, 4) {real, imag} */,
  {32'hbf05eefc, 32'h00000000} /* (19, 27, 3) {real, imag} */,
  {32'hbf0277e0, 32'h00000000} /* (19, 27, 2) {real, imag} */,
  {32'hbf4e931b, 32'h00000000} /* (19, 27, 1) {real, imag} */,
  {32'hbed84ddb, 32'h00000000} /* (19, 27, 0) {real, imag} */,
  {32'hbf14d7c6, 32'h00000000} /* (19, 26, 31) {real, imag} */,
  {32'hbf357aa8, 32'h00000000} /* (19, 26, 30) {real, imag} */,
  {32'hbf4ffe4a, 32'h00000000} /* (19, 26, 29) {real, imag} */,
  {32'hbf8fb86d, 32'h00000000} /* (19, 26, 28) {real, imag} */,
  {32'hbf2cdf4e, 32'h00000000} /* (19, 26, 27) {real, imag} */,
  {32'hbf3b1f0f, 32'h00000000} /* (19, 26, 26) {real, imag} */,
  {32'hbf9c384e, 32'h00000000} /* (19, 26, 25) {real, imag} */,
  {32'hbf6c90a5, 32'h00000000} /* (19, 26, 24) {real, imag} */,
  {32'hbf819ef8, 32'h00000000} /* (19, 26, 23) {real, imag} */,
  {32'hbf463040, 32'h00000000} /* (19, 26, 22) {real, imag} */,
  {32'hbecfa152, 32'h00000000} /* (19, 26, 21) {real, imag} */,
  {32'h3e61fbb7, 32'h00000000} /* (19, 26, 20) {real, imag} */,
  {32'h3f042951, 32'h00000000} /* (19, 26, 19) {real, imag} */,
  {32'h3f025d81, 32'h00000000} /* (19, 26, 18) {real, imag} */,
  {32'h3f3803c6, 32'h00000000} /* (19, 26, 17) {real, imag} */,
  {32'h3ef6072d, 32'h00000000} /* (19, 26, 16) {real, imag} */,
  {32'h3f99314f, 32'h00000000} /* (19, 26, 15) {real, imag} */,
  {32'h3fbe47fd, 32'h00000000} /* (19, 26, 14) {real, imag} */,
  {32'h3fb91dc3, 32'h00000000} /* (19, 26, 13) {real, imag} */,
  {32'h3f7d412f, 32'h00000000} /* (19, 26, 12) {real, imag} */,
  {32'h3e9f34fb, 32'h00000000} /* (19, 26, 11) {real, imag} */,
  {32'hbe8a4ae6, 32'h00000000} /* (19, 26, 10) {real, imag} */,
  {32'hbf7be679, 32'h00000000} /* (19, 26, 9) {real, imag} */,
  {32'hbfc94afe, 32'h00000000} /* (19, 26, 8) {real, imag} */,
  {32'hbf854b27, 32'h00000000} /* (19, 26, 7) {real, imag} */,
  {32'hbf387d41, 32'h00000000} /* (19, 26, 6) {real, imag} */,
  {32'hbf803cc0, 32'h00000000} /* (19, 26, 5) {real, imag} */,
  {32'hbf4fc0ce, 32'h00000000} /* (19, 26, 4) {real, imag} */,
  {32'hbef13db8, 32'h00000000} /* (19, 26, 3) {real, imag} */,
  {32'hbf49ab06, 32'h00000000} /* (19, 26, 2) {real, imag} */,
  {32'hbfa01a0e, 32'h00000000} /* (19, 26, 1) {real, imag} */,
  {32'hbf490f42, 32'h00000000} /* (19, 26, 0) {real, imag} */,
  {32'hbf2dfee6, 32'h00000000} /* (19, 25, 31) {real, imag} */,
  {32'hbf7bcedc, 32'h00000000} /* (19, 25, 30) {real, imag} */,
  {32'hbf56d8e8, 32'h00000000} /* (19, 25, 29) {real, imag} */,
  {32'hbf717a42, 32'h00000000} /* (19, 25, 28) {real, imag} */,
  {32'hbfb3bb08, 32'h00000000} /* (19, 25, 27) {real, imag} */,
  {32'hbfc1974d, 32'h00000000} /* (19, 25, 26) {real, imag} */,
  {32'hbf8d9fd5, 32'h00000000} /* (19, 25, 25) {real, imag} */,
  {32'hbf112c6f, 32'h00000000} /* (19, 25, 24) {real, imag} */,
  {32'hbf94832a, 32'h00000000} /* (19, 25, 23) {real, imag} */,
  {32'hbfc00a6a, 32'h00000000} /* (19, 25, 22) {real, imag} */,
  {32'hbf7c3b6c, 32'h00000000} /* (19, 25, 21) {real, imag} */,
  {32'h3f48fea5, 32'h00000000} /* (19, 25, 20) {real, imag} */,
  {32'h3fa26c67, 32'h00000000} /* (19, 25, 19) {real, imag} */,
  {32'h3f5d6743, 32'h00000000} /* (19, 25, 18) {real, imag} */,
  {32'h3f21c5d4, 32'h00000000} /* (19, 25, 17) {real, imag} */,
  {32'h3e0a143a, 32'h00000000} /* (19, 25, 16) {real, imag} */,
  {32'h3f25ef8b, 32'h00000000} /* (19, 25, 15) {real, imag} */,
  {32'h3f9021ac, 32'h00000000} /* (19, 25, 14) {real, imag} */,
  {32'h3fcff5fe, 32'h00000000} /* (19, 25, 13) {real, imag} */,
  {32'h3f8536b2, 32'h00000000} /* (19, 25, 12) {real, imag} */,
  {32'h3ee6a1cc, 32'h00000000} /* (19, 25, 11) {real, imag} */,
  {32'hbe936ea3, 32'h00000000} /* (19, 25, 10) {real, imag} */,
  {32'hbf87cb4c, 32'h00000000} /* (19, 25, 9) {real, imag} */,
  {32'hbfe4acf4, 32'h00000000} /* (19, 25, 8) {real, imag} */,
  {32'hbfa4c0dc, 32'h00000000} /* (19, 25, 7) {real, imag} */,
  {32'hbf15986d, 32'h00000000} /* (19, 25, 6) {real, imag} */,
  {32'hbea41767, 32'h00000000} /* (19, 25, 5) {real, imag} */,
  {32'hbf019298, 32'h00000000} /* (19, 25, 4) {real, imag} */,
  {32'hbf0caf47, 32'h00000000} /* (19, 25, 3) {real, imag} */,
  {32'hbfa499ad, 32'h00000000} /* (19, 25, 2) {real, imag} */,
  {32'hbfd31f4e, 32'h00000000} /* (19, 25, 1) {real, imag} */,
  {32'hbf3f0994, 32'h00000000} /* (19, 25, 0) {real, imag} */,
  {32'hbee55c03, 32'h00000000} /* (19, 24, 31) {real, imag} */,
  {32'hbf17c40c, 32'h00000000} /* (19, 24, 30) {real, imag} */,
  {32'hbecb4ed8, 32'h00000000} /* (19, 24, 29) {real, imag} */,
  {32'hbeff2a8a, 32'h00000000} /* (19, 24, 28) {real, imag} */,
  {32'hbf6e3e94, 32'h00000000} /* (19, 24, 27) {real, imag} */,
  {32'hbf41bc11, 32'h00000000} /* (19, 24, 26) {real, imag} */,
  {32'hbf6155e5, 32'h00000000} /* (19, 24, 25) {real, imag} */,
  {32'hbf8ef3cf, 32'h00000000} /* (19, 24, 24) {real, imag} */,
  {32'hbff962e4, 32'h00000000} /* (19, 24, 23) {real, imag} */,
  {32'hbfb1b107, 32'h00000000} /* (19, 24, 22) {real, imag} */,
  {32'hbf0369eb, 32'h00000000} /* (19, 24, 21) {real, imag} */,
  {32'h3f8d5c87, 32'h00000000} /* (19, 24, 20) {real, imag} */,
  {32'h3fa3d14d, 32'h00000000} /* (19, 24, 19) {real, imag} */,
  {32'h3f900210, 32'h00000000} /* (19, 24, 18) {real, imag} */,
  {32'h3f4c9387, 32'h00000000} /* (19, 24, 17) {real, imag} */,
  {32'h3f1be16d, 32'h00000000} /* (19, 24, 16) {real, imag} */,
  {32'h3f7c4944, 32'h00000000} /* (19, 24, 15) {real, imag} */,
  {32'h3f9b6cee, 32'h00000000} /* (19, 24, 14) {real, imag} */,
  {32'h3f0a65f5, 32'h00000000} /* (19, 24, 13) {real, imag} */,
  {32'h3f17fca1, 32'h00000000} /* (19, 24, 12) {real, imag} */,
  {32'h3ee3ebc9, 32'h00000000} /* (19, 24, 11) {real, imag} */,
  {32'hbf33e2ea, 32'h00000000} /* (19, 24, 10) {real, imag} */,
  {32'hbfbae6ed, 32'h00000000} /* (19, 24, 9) {real, imag} */,
  {32'hbff5ae9f, 32'h00000000} /* (19, 24, 8) {real, imag} */,
  {32'hbfa28606, 32'h00000000} /* (19, 24, 7) {real, imag} */,
  {32'hbf4725f5, 32'h00000000} /* (19, 24, 6) {real, imag} */,
  {32'hbf0cafde, 32'h00000000} /* (19, 24, 5) {real, imag} */,
  {32'hbf32004f, 32'h00000000} /* (19, 24, 4) {real, imag} */,
  {32'hbf51a7c6, 32'h00000000} /* (19, 24, 3) {real, imag} */,
  {32'hbf920b22, 32'h00000000} /* (19, 24, 2) {real, imag} */,
  {32'hbf8a71d2, 32'h00000000} /* (19, 24, 1) {real, imag} */,
  {32'hbef4bc31, 32'h00000000} /* (19, 24, 0) {real, imag} */,
  {32'hbee06c24, 32'h00000000} /* (19, 23, 31) {real, imag} */,
  {32'hbf1bdfcc, 32'h00000000} /* (19, 23, 30) {real, imag} */,
  {32'hbeff168e, 32'h00000000} /* (19, 23, 29) {real, imag} */,
  {32'hbf40751b, 32'h00000000} /* (19, 23, 28) {real, imag} */,
  {32'hbf182554, 32'h00000000} /* (19, 23, 27) {real, imag} */,
  {32'hbecc80ed, 32'h00000000} /* (19, 23, 26) {real, imag} */,
  {32'hbf5290d8, 32'h00000000} /* (19, 23, 25) {real, imag} */,
  {32'hbfe152ab, 32'h00000000} /* (19, 23, 24) {real, imag} */,
  {32'hc0125676, 32'h00000000} /* (19, 23, 23) {real, imag} */,
  {32'hbffa32a6, 32'h00000000} /* (19, 23, 22) {real, imag} */,
  {32'hbf91810d, 32'h00000000} /* (19, 23, 21) {real, imag} */,
  {32'h3f3b5a41, 32'h00000000} /* (19, 23, 20) {real, imag} */,
  {32'h3fc72049, 32'h00000000} /* (19, 23, 19) {real, imag} */,
  {32'h3fcdd408, 32'h00000000} /* (19, 23, 18) {real, imag} */,
  {32'h3f634ae0, 32'h00000000} /* (19, 23, 17) {real, imag} */,
  {32'h3f862cde, 32'h00000000} /* (19, 23, 16) {real, imag} */,
  {32'h3f82f34a, 32'h00000000} /* (19, 23, 15) {real, imag} */,
  {32'h3f8c6143, 32'h00000000} /* (19, 23, 14) {real, imag} */,
  {32'h3f09a813, 32'h00000000} /* (19, 23, 13) {real, imag} */,
  {32'h3f504892, 32'h00000000} /* (19, 23, 12) {real, imag} */,
  {32'h3ed37dcc, 32'h00000000} /* (19, 23, 11) {real, imag} */,
  {32'hbf80ff48, 32'h00000000} /* (19, 23, 10) {real, imag} */,
  {32'hbf87b53c, 32'h00000000} /* (19, 23, 9) {real, imag} */,
  {32'hbf7c5452, 32'h00000000} /* (19, 23, 8) {real, imag} */,
  {32'hbf72691a, 32'h00000000} /* (19, 23, 7) {real, imag} */,
  {32'hbf97af17, 32'h00000000} /* (19, 23, 6) {real, imag} */,
  {32'hbfa1ad50, 32'h00000000} /* (19, 23, 5) {real, imag} */,
  {32'hbf8faccf, 32'h00000000} /* (19, 23, 4) {real, imag} */,
  {32'hbf72a6e8, 32'h00000000} /* (19, 23, 3) {real, imag} */,
  {32'hbf8c2cc3, 32'h00000000} /* (19, 23, 2) {real, imag} */,
  {32'hbf8bb75d, 32'h00000000} /* (19, 23, 1) {real, imag} */,
  {32'hbed619c3, 32'h00000000} /* (19, 23, 0) {real, imag} */,
  {32'hbeb063ed, 32'h00000000} /* (19, 22, 31) {real, imag} */,
  {32'hbf80ee7c, 32'h00000000} /* (19, 22, 30) {real, imag} */,
  {32'hbf9d1df6, 32'h00000000} /* (19, 22, 29) {real, imag} */,
  {32'hbfb147bb, 32'h00000000} /* (19, 22, 28) {real, imag} */,
  {32'hbfa7d3a7, 32'h00000000} /* (19, 22, 27) {real, imag} */,
  {32'hbf834a70, 32'h00000000} /* (19, 22, 26) {real, imag} */,
  {32'hbf109ba0, 32'h00000000} /* (19, 22, 25) {real, imag} */,
  {32'hbf7174c5, 32'h00000000} /* (19, 22, 24) {real, imag} */,
  {32'hbfb39c12, 32'h00000000} /* (19, 22, 23) {real, imag} */,
  {32'hbfafcba6, 32'h00000000} /* (19, 22, 22) {real, imag} */,
  {32'hbf3f2be5, 32'h00000000} /* (19, 22, 21) {real, imag} */,
  {32'h3ebd33ef, 32'h00000000} /* (19, 22, 20) {real, imag} */,
  {32'h3f80edae, 32'h00000000} /* (19, 22, 19) {real, imag} */,
  {32'h3f6b99d1, 32'h00000000} /* (19, 22, 18) {real, imag} */,
  {32'h3f5d7391, 32'h00000000} /* (19, 22, 17) {real, imag} */,
  {32'h3f91a585, 32'h00000000} /* (19, 22, 16) {real, imag} */,
  {32'h3f3dc4f5, 32'h00000000} /* (19, 22, 15) {real, imag} */,
  {32'h3f830dbf, 32'h00000000} /* (19, 22, 14) {real, imag} */,
  {32'h3f93b028, 32'h00000000} /* (19, 22, 13) {real, imag} */,
  {32'h3f346b70, 32'h00000000} /* (19, 22, 12) {real, imag} */,
  {32'h3ea6d9da, 32'h00000000} /* (19, 22, 11) {real, imag} */,
  {32'hbf78f9b1, 32'h00000000} /* (19, 22, 10) {real, imag} */,
  {32'hbfc66d38, 32'h00000000} /* (19, 22, 9) {real, imag} */,
  {32'hbf99f2c0, 32'h00000000} /* (19, 22, 8) {real, imag} */,
  {32'hbf9be299, 32'h00000000} /* (19, 22, 7) {real, imag} */,
  {32'hbf5b05dc, 32'h00000000} /* (19, 22, 6) {real, imag} */,
  {32'hbf0a1c31, 32'h00000000} /* (19, 22, 5) {real, imag} */,
  {32'hbf44b7e1, 32'h00000000} /* (19, 22, 4) {real, imag} */,
  {32'hbf351e09, 32'h00000000} /* (19, 22, 3) {real, imag} */,
  {32'hbfa0c24d, 32'h00000000} /* (19, 22, 2) {real, imag} */,
  {32'hbfd957ed, 32'h00000000} /* (19, 22, 1) {real, imag} */,
  {32'hbf5e59f5, 32'h00000000} /* (19, 22, 0) {real, imag} */,
  {32'hbea94c09, 32'h00000000} /* (19, 21, 31) {real, imag} */,
  {32'hbf42f241, 32'h00000000} /* (19, 21, 30) {real, imag} */,
  {32'hbf510b56, 32'h00000000} /* (19, 21, 29) {real, imag} */,
  {32'hbf08d52e, 32'h00000000} /* (19, 21, 28) {real, imag} */,
  {32'hbf1ab4d9, 32'h00000000} /* (19, 21, 27) {real, imag} */,
  {32'hbf5224a5, 32'h00000000} /* (19, 21, 26) {real, imag} */,
  {32'hbf11d62e, 32'h00000000} /* (19, 21, 25) {real, imag} */,
  {32'hbebc26dc, 32'h00000000} /* (19, 21, 24) {real, imag} */,
  {32'hbeed5dd3, 32'h00000000} /* (19, 21, 23) {real, imag} */,
  {32'hbe97cffe, 32'h00000000} /* (19, 21, 22) {real, imag} */,
  {32'hbdaeb0d6, 32'h00000000} /* (19, 21, 21) {real, imag} */,
  {32'hbeae84ac, 32'h00000000} /* (19, 21, 20) {real, imag} */,
  {32'h3e021584, 32'h00000000} /* (19, 21, 19) {real, imag} */,
  {32'h3e5d6f31, 32'h00000000} /* (19, 21, 18) {real, imag} */,
  {32'h3e843482, 32'h00000000} /* (19, 21, 17) {real, imag} */,
  {32'h3ecc2936, 32'h00000000} /* (19, 21, 16) {real, imag} */,
  {32'h3ef3d8aa, 32'h00000000} /* (19, 21, 15) {real, imag} */,
  {32'h3f3b784c, 32'h00000000} /* (19, 21, 14) {real, imag} */,
  {32'h3f31a56e, 32'h00000000} /* (19, 21, 13) {real, imag} */,
  {32'h3ea54197, 32'h00000000} /* (19, 21, 12) {real, imag} */,
  {32'h3dabd58e, 32'h00000000} /* (19, 21, 11) {real, imag} */,
  {32'hbf3ed12f, 32'h00000000} /* (19, 21, 10) {real, imag} */,
  {32'hbf8a321d, 32'h00000000} /* (19, 21, 9) {real, imag} */,
  {32'hbf33d91f, 32'h00000000} /* (19, 21, 8) {real, imag} */,
  {32'hbf451a13, 32'h00000000} /* (19, 21, 7) {real, imag} */,
  {32'hbe4dfd0b, 32'h00000000} /* (19, 21, 6) {real, imag} */,
  {32'h3e3cae3e, 32'h00000000} /* (19, 21, 5) {real, imag} */,
  {32'hbd00571f, 32'h00000000} /* (19, 21, 4) {real, imag} */,
  {32'h3d63dc02, 32'h00000000} /* (19, 21, 3) {real, imag} */,
  {32'hbec35aa4, 32'h00000000} /* (19, 21, 2) {real, imag} */,
  {32'hbf089954, 32'h00000000} /* (19, 21, 1) {real, imag} */,
  {32'hbe2283bf, 32'h00000000} /* (19, 21, 0) {real, imag} */,
  {32'h3ef6eb8c, 32'h00000000} /* (19, 20, 31) {real, imag} */,
  {32'h3f05c726, 32'h00000000} /* (19, 20, 30) {real, imag} */,
  {32'h3e96b0dd, 32'h00000000} /* (19, 20, 29) {real, imag} */,
  {32'h3f959512, 32'h00000000} /* (19, 20, 28) {real, imag} */,
  {32'h3fb3697a, 32'h00000000} /* (19, 20, 27) {real, imag} */,
  {32'h3f0d3be9, 32'h00000000} /* (19, 20, 26) {real, imag} */,
  {32'h3e3566d5, 32'h00000000} /* (19, 20, 25) {real, imag} */,
  {32'h3f3ce69a, 32'h00000000} /* (19, 20, 24) {real, imag} */,
  {32'h3f580393, 32'h00000000} /* (19, 20, 23) {real, imag} */,
  {32'h3f32307e, 32'h00000000} /* (19, 20, 22) {real, imag} */,
  {32'h3e8d967c, 32'h00000000} /* (19, 20, 21) {real, imag} */,
  {32'hbf3c88fa, 32'h00000000} /* (19, 20, 20) {real, imag} */,
  {32'hbf287b48, 32'h00000000} /* (19, 20, 19) {real, imag} */,
  {32'hbeb116a0, 32'h00000000} /* (19, 20, 18) {real, imag} */,
  {32'hbecddf3f, 32'h00000000} /* (19, 20, 17) {real, imag} */,
  {32'hbea8dcff, 32'h00000000} /* (19, 20, 16) {real, imag} */,
  {32'hbee260bb, 32'h00000000} /* (19, 20, 15) {real, imag} */,
  {32'hbec63cec, 32'h00000000} /* (19, 20, 14) {real, imag} */,
  {32'hbf6c144e, 32'h00000000} /* (19, 20, 13) {real, imag} */,
  {32'hbfae8974, 32'h00000000} /* (19, 20, 12) {real, imag} */,
  {32'hbf8c5986, 32'h00000000} /* (19, 20, 11) {real, imag} */,
  {32'h3d875f20, 32'h00000000} /* (19, 20, 10) {real, imag} */,
  {32'h3e808b3d, 32'h00000000} /* (19, 20, 9) {real, imag} */,
  {32'h3f056a64, 32'h00000000} /* (19, 20, 8) {real, imag} */,
  {32'h3ecebe6b, 32'h00000000} /* (19, 20, 7) {real, imag} */,
  {32'h3f2b4a3d, 32'h00000000} /* (19, 20, 6) {real, imag} */,
  {32'h3f31dcc8, 32'h00000000} /* (19, 20, 5) {real, imag} */,
  {32'h3eb3ea8e, 32'h00000000} /* (19, 20, 4) {real, imag} */,
  {32'h3f4ff6c0, 32'h00000000} /* (19, 20, 3) {real, imag} */,
  {32'h3f83256c, 32'h00000000} /* (19, 20, 2) {real, imag} */,
  {32'h3f492173, 32'h00000000} /* (19, 20, 1) {real, imag} */,
  {32'h3f13be89, 32'h00000000} /* (19, 20, 0) {real, imag} */,
  {32'h3f0899c6, 32'h00000000} /* (19, 19, 31) {real, imag} */,
  {32'h3f47c59f, 32'h00000000} /* (19, 19, 30) {real, imag} */,
  {32'h3f49b1c1, 32'h00000000} /* (19, 19, 29) {real, imag} */,
  {32'h3fdc9fa0, 32'h00000000} /* (19, 19, 28) {real, imag} */,
  {32'h3fcbe3a6, 32'h00000000} /* (19, 19, 27) {real, imag} */,
  {32'h3f5b76c6, 32'h00000000} /* (19, 19, 26) {real, imag} */,
  {32'h3f82a5de, 32'h00000000} /* (19, 19, 25) {real, imag} */,
  {32'h3fe4a669, 32'h00000000} /* (19, 19, 24) {real, imag} */,
  {32'h3f8a88a5, 32'h00000000} /* (19, 19, 23) {real, imag} */,
  {32'h3f539adf, 32'h00000000} /* (19, 19, 22) {real, imag} */,
  {32'h3eaf3ab4, 32'h00000000} /* (19, 19, 21) {real, imag} */,
  {32'hbf9aeb41, 32'h00000000} /* (19, 19, 20) {real, imag} */,
  {32'hbfbbf199, 32'h00000000} /* (19, 19, 19) {real, imag} */,
  {32'hbf8330a4, 32'h00000000} /* (19, 19, 18) {real, imag} */,
  {32'hbf441e1d, 32'h00000000} /* (19, 19, 17) {real, imag} */,
  {32'hbf56c7b9, 32'h00000000} /* (19, 19, 16) {real, imag} */,
  {32'hbf833a3a, 32'h00000000} /* (19, 19, 15) {real, imag} */,
  {32'hbf0d7d28, 32'h00000000} /* (19, 19, 14) {real, imag} */,
  {32'hbf31f059, 32'h00000000} /* (19, 19, 13) {real, imag} */,
  {32'hbf93e6f6, 32'h00000000} /* (19, 19, 12) {real, imag} */,
  {32'hbf8313d7, 32'h00000000} /* (19, 19, 11) {real, imag} */,
  {32'hbcdf6be0, 32'h00000000} /* (19, 19, 10) {real, imag} */,
  {32'h3f598ef9, 32'h00000000} /* (19, 19, 9) {real, imag} */,
  {32'h3f770e3b, 32'h00000000} /* (19, 19, 8) {real, imag} */,
  {32'h3f5b76fa, 32'h00000000} /* (19, 19, 7) {real, imag} */,
  {32'h3ed49489, 32'h00000000} /* (19, 19, 6) {real, imag} */,
  {32'h3ede1d39, 32'h00000000} /* (19, 19, 5) {real, imag} */,
  {32'h3f7297ab, 32'h00000000} /* (19, 19, 4) {real, imag} */,
  {32'h3f4a1030, 32'h00000000} /* (19, 19, 3) {real, imag} */,
  {32'h3f993782, 32'h00000000} /* (19, 19, 2) {real, imag} */,
  {32'h3fbf7ef3, 32'h00000000} /* (19, 19, 1) {real, imag} */,
  {32'h3f8df0ae, 32'h00000000} /* (19, 19, 0) {real, imag} */,
  {32'h3f2deaa2, 32'h00000000} /* (19, 18, 31) {real, imag} */,
  {32'h3f88a113, 32'h00000000} /* (19, 18, 30) {real, imag} */,
  {32'h3f091f59, 32'h00000000} /* (19, 18, 29) {real, imag} */,
  {32'h3f0d2df5, 32'h00000000} /* (19, 18, 28) {real, imag} */,
  {32'h3f0a467f, 32'h00000000} /* (19, 18, 27) {real, imag} */,
  {32'h3f23cdc6, 32'h00000000} /* (19, 18, 26) {real, imag} */,
  {32'h3fd0f7a8, 32'h00000000} /* (19, 18, 25) {real, imag} */,
  {32'h3fdd9ea0, 32'h00000000} /* (19, 18, 24) {real, imag} */,
  {32'h3f25afa3, 32'h00000000} /* (19, 18, 23) {real, imag} */,
  {32'h3ee5cb79, 32'h00000000} /* (19, 18, 22) {real, imag} */,
  {32'h3edf7cff, 32'h00000000} /* (19, 18, 21) {real, imag} */,
  {32'hbf3355bb, 32'h00000000} /* (19, 18, 20) {real, imag} */,
  {32'hbf7e951a, 32'h00000000} /* (19, 18, 19) {real, imag} */,
  {32'hbf8e54bd, 32'h00000000} /* (19, 18, 18) {real, imag} */,
  {32'hbf9c3761, 32'h00000000} /* (19, 18, 17) {real, imag} */,
  {32'hbfb5c9cd, 32'h00000000} /* (19, 18, 16) {real, imag} */,
  {32'hbf94673f, 32'h00000000} /* (19, 18, 15) {real, imag} */,
  {32'hbf262932, 32'h00000000} /* (19, 18, 14) {real, imag} */,
  {32'hbf009be3, 32'h00000000} /* (19, 18, 13) {real, imag} */,
  {32'hbf832ed7, 32'h00000000} /* (19, 18, 12) {real, imag} */,
  {32'hbf3a1a63, 32'h00000000} /* (19, 18, 11) {real, imag} */,
  {32'h3f2ca432, 32'h00000000} /* (19, 18, 10) {real, imag} */,
  {32'h3f8f2a6c, 32'h00000000} /* (19, 18, 9) {real, imag} */,
  {32'h3f5f4a0b, 32'h00000000} /* (19, 18, 8) {real, imag} */,
  {32'h3f7d5b01, 32'h00000000} /* (19, 18, 7) {real, imag} */,
  {32'h3f1347d3, 32'h00000000} /* (19, 18, 6) {real, imag} */,
  {32'h3f5208cb, 32'h00000000} /* (19, 18, 5) {real, imag} */,
  {32'h3fb460d9, 32'h00000000} /* (19, 18, 4) {real, imag} */,
  {32'h3f343611, 32'h00000000} /* (19, 18, 3) {real, imag} */,
  {32'h3f26d568, 32'h00000000} /* (19, 18, 2) {real, imag} */,
  {32'h3f9bb9d6, 32'h00000000} /* (19, 18, 1) {real, imag} */,
  {32'h3fb67c10, 32'h00000000} /* (19, 18, 0) {real, imag} */,
  {32'h3ee11651, 32'h00000000} /* (19, 17, 31) {real, imag} */,
  {32'h3f49eb68, 32'h00000000} /* (19, 17, 30) {real, imag} */,
  {32'h3f59f968, 32'h00000000} /* (19, 17, 29) {real, imag} */,
  {32'h3f437579, 32'h00000000} /* (19, 17, 28) {real, imag} */,
  {32'h3f927197, 32'h00000000} /* (19, 17, 27) {real, imag} */,
  {32'h3f6c41f1, 32'h00000000} /* (19, 17, 26) {real, imag} */,
  {32'h3f82c5c7, 32'h00000000} /* (19, 17, 25) {real, imag} */,
  {32'h3f5b5af9, 32'h00000000} /* (19, 17, 24) {real, imag} */,
  {32'h3f3096de, 32'h00000000} /* (19, 17, 23) {real, imag} */,
  {32'h3f49a907, 32'h00000000} /* (19, 17, 22) {real, imag} */,
  {32'h3e6b9ad0, 32'h00000000} /* (19, 17, 21) {real, imag} */,
  {32'hbf076453, 32'h00000000} /* (19, 17, 20) {real, imag} */,
  {32'hbf40e9a7, 32'h00000000} /* (19, 17, 19) {real, imag} */,
  {32'hbf3cf63d, 32'h00000000} /* (19, 17, 18) {real, imag} */,
  {32'hbf5359da, 32'h00000000} /* (19, 17, 17) {real, imag} */,
  {32'hbfc19ddc, 32'h00000000} /* (19, 17, 16) {real, imag} */,
  {32'hbf8b6006, 32'h00000000} /* (19, 17, 15) {real, imag} */,
  {32'hbece30dd, 32'h00000000} /* (19, 17, 14) {real, imag} */,
  {32'hbe77eb4a, 32'h00000000} /* (19, 17, 13) {real, imag} */,
  {32'hbf613bac, 32'h00000000} /* (19, 17, 12) {real, imag} */,
  {32'hbf520f3d, 32'h00000000} /* (19, 17, 11) {real, imag} */,
  {32'h3f0a33a9, 32'h00000000} /* (19, 17, 10) {real, imag} */,
  {32'h3f3c1b7c, 32'h00000000} /* (19, 17, 9) {real, imag} */,
  {32'h3f7efca9, 32'h00000000} /* (19, 17, 8) {real, imag} */,
  {32'h3f784a13, 32'h00000000} /* (19, 17, 7) {real, imag} */,
  {32'h3f6ca15b, 32'h00000000} /* (19, 17, 6) {real, imag} */,
  {32'h3f73c23a, 32'h00000000} /* (19, 17, 5) {real, imag} */,
  {32'h3fa94a4f, 32'h00000000} /* (19, 17, 4) {real, imag} */,
  {32'h3f2c373f, 32'h00000000} /* (19, 17, 3) {real, imag} */,
  {32'h3f64a15d, 32'h00000000} /* (19, 17, 2) {real, imag} */,
  {32'h3f61e226, 32'h00000000} /* (19, 17, 1) {real, imag} */,
  {32'h3f4b6a44, 32'h00000000} /* (19, 17, 0) {real, imag} */,
  {32'h3f113515, 32'h00000000} /* (19, 16, 31) {real, imag} */,
  {32'h3f455871, 32'h00000000} /* (19, 16, 30) {real, imag} */,
  {32'h3f6f8ba6, 32'h00000000} /* (19, 16, 29) {real, imag} */,
  {32'h3f9f7b0c, 32'h00000000} /* (19, 16, 28) {real, imag} */,
  {32'h3fc9be8a, 32'h00000000} /* (19, 16, 27) {real, imag} */,
  {32'h3f9c64f3, 32'h00000000} /* (19, 16, 26) {real, imag} */,
  {32'h3fa0da65, 32'h00000000} /* (19, 16, 25) {real, imag} */,
  {32'h3fa81134, 32'h00000000} /* (19, 16, 24) {real, imag} */,
  {32'h3f5196a4, 32'h00000000} /* (19, 16, 23) {real, imag} */,
  {32'h3f12b0b6, 32'h00000000} /* (19, 16, 22) {real, imag} */,
  {32'h3d73afee, 32'h00000000} /* (19, 16, 21) {real, imag} */,
  {32'hbf9dd69b, 32'h00000000} /* (19, 16, 20) {real, imag} */,
  {32'hbf96437e, 32'h00000000} /* (19, 16, 19) {real, imag} */,
  {32'hbf7ac9d3, 32'h00000000} /* (19, 16, 18) {real, imag} */,
  {32'hbf69b136, 32'h00000000} /* (19, 16, 17) {real, imag} */,
  {32'hbf79713f, 32'h00000000} /* (19, 16, 16) {real, imag} */,
  {32'hbf8429b5, 32'h00000000} /* (19, 16, 15) {real, imag} */,
  {32'hbf49869c, 32'h00000000} /* (19, 16, 14) {real, imag} */,
  {32'hbf4f334e, 32'h00000000} /* (19, 16, 13) {real, imag} */,
  {32'hbf4d8b2c, 32'h00000000} /* (19, 16, 12) {real, imag} */,
  {32'hbf83263d, 32'h00000000} /* (19, 16, 11) {real, imag} */,
  {32'h3eff6c95, 32'h00000000} /* (19, 16, 10) {real, imag} */,
  {32'h3fa546c3, 32'h00000000} /* (19, 16, 9) {real, imag} */,
  {32'h3fa4de97, 32'h00000000} /* (19, 16, 8) {real, imag} */,
  {32'h3f9b06af, 32'h00000000} /* (19, 16, 7) {real, imag} */,
  {32'h3f644f34, 32'h00000000} /* (19, 16, 6) {real, imag} */,
  {32'h3f1671c7, 32'h00000000} /* (19, 16, 5) {real, imag} */,
  {32'h3f2747d9, 32'h00000000} /* (19, 16, 4) {real, imag} */,
  {32'h3f2d9424, 32'h00000000} /* (19, 16, 3) {real, imag} */,
  {32'h3f2771cd, 32'h00000000} /* (19, 16, 2) {real, imag} */,
  {32'h3ee2350b, 32'h00000000} /* (19, 16, 1) {real, imag} */,
  {32'h3d93ac8f, 32'h00000000} /* (19, 16, 0) {real, imag} */,
  {32'h3f309ac4, 32'h00000000} /* (19, 15, 31) {real, imag} */,
  {32'h3f86cdd5, 32'h00000000} /* (19, 15, 30) {real, imag} */,
  {32'h3f6ea276, 32'h00000000} /* (19, 15, 29) {real, imag} */,
  {32'h3f99a006, 32'h00000000} /* (19, 15, 28) {real, imag} */,
  {32'h3f977841, 32'h00000000} /* (19, 15, 27) {real, imag} */,
  {32'h3fc5799a, 32'h00000000} /* (19, 15, 26) {real, imag} */,
  {32'h3fadf6eb, 32'h00000000} /* (19, 15, 25) {real, imag} */,
  {32'h3fd42aac, 32'h00000000} /* (19, 15, 24) {real, imag} */,
  {32'h3fa6b711, 32'h00000000} /* (19, 15, 23) {real, imag} */,
  {32'h3f88dbfa, 32'h00000000} /* (19, 15, 22) {real, imag} */,
  {32'h3f234096, 32'h00000000} /* (19, 15, 21) {real, imag} */,
  {32'hbf40ca43, 32'h00000000} /* (19, 15, 20) {real, imag} */,
  {32'hbfc947c5, 32'h00000000} /* (19, 15, 19) {real, imag} */,
  {32'hbf98378f, 32'h00000000} /* (19, 15, 18) {real, imag} */,
  {32'hbf6af88a, 32'h00000000} /* (19, 15, 17) {real, imag} */,
  {32'hbf55129c, 32'h00000000} /* (19, 15, 16) {real, imag} */,
  {32'hbf9aca71, 32'h00000000} /* (19, 15, 15) {real, imag} */,
  {32'hbf8ff22c, 32'h00000000} /* (19, 15, 14) {real, imag} */,
  {32'hbf77ce68, 32'h00000000} /* (19, 15, 13) {real, imag} */,
  {32'hbf426f88, 32'h00000000} /* (19, 15, 12) {real, imag} */,
  {32'hbf9a59c9, 32'h00000000} /* (19, 15, 11) {real, imag} */,
  {32'h3eb75079, 32'h00000000} /* (19, 15, 10) {real, imag} */,
  {32'h3f9ce4ba, 32'h00000000} /* (19, 15, 9) {real, imag} */,
  {32'h3fcc269a, 32'h00000000} /* (19, 15, 8) {real, imag} */,
  {32'h3fd505e5, 32'h00000000} /* (19, 15, 7) {real, imag} */,
  {32'h3f830374, 32'h00000000} /* (19, 15, 6) {real, imag} */,
  {32'h3f5b6f67, 32'h00000000} /* (19, 15, 5) {real, imag} */,
  {32'h3f512c72, 32'h00000000} /* (19, 15, 4) {real, imag} */,
  {32'h3f63f0e4, 32'h00000000} /* (19, 15, 3) {real, imag} */,
  {32'h3f1bf944, 32'h00000000} /* (19, 15, 2) {real, imag} */,
  {32'h3f1c9942, 32'h00000000} /* (19, 15, 1) {real, imag} */,
  {32'h3e6c7226, 32'h00000000} /* (19, 15, 0) {real, imag} */,
  {32'h3ea88795, 32'h00000000} /* (19, 14, 31) {real, imag} */,
  {32'h3f3544b7, 32'h00000000} /* (19, 14, 30) {real, imag} */,
  {32'h3f55da4b, 32'h00000000} /* (19, 14, 29) {real, imag} */,
  {32'h3fb338e3, 32'h00000000} /* (19, 14, 28) {real, imag} */,
  {32'h3f493970, 32'h00000000} /* (19, 14, 27) {real, imag} */,
  {32'h3f661f8d, 32'h00000000} /* (19, 14, 26) {real, imag} */,
  {32'h3f887559, 32'h00000000} /* (19, 14, 25) {real, imag} */,
  {32'h3fbcae4b, 32'h00000000} /* (19, 14, 24) {real, imag} */,
  {32'h3f8c6600, 32'h00000000} /* (19, 14, 23) {real, imag} */,
  {32'h3fa529a3, 32'h00000000} /* (19, 14, 22) {real, imag} */,
  {32'h3f3bc38a, 32'h00000000} /* (19, 14, 21) {real, imag} */,
  {32'hbf85245e, 32'h00000000} /* (19, 14, 20) {real, imag} */,
  {32'hbfa8a9fe, 32'h00000000} /* (19, 14, 19) {real, imag} */,
  {32'hbf3e11d8, 32'h00000000} /* (19, 14, 18) {real, imag} */,
  {32'hbf73bf0c, 32'h00000000} /* (19, 14, 17) {real, imag} */,
  {32'hbf9da3da, 32'h00000000} /* (19, 14, 16) {real, imag} */,
  {32'hbfbba841, 32'h00000000} /* (19, 14, 15) {real, imag} */,
  {32'hbfaf7458, 32'h00000000} /* (19, 14, 14) {real, imag} */,
  {32'hbf4f3dfe, 32'h00000000} /* (19, 14, 13) {real, imag} */,
  {32'hbf051f52, 32'h00000000} /* (19, 14, 12) {real, imag} */,
  {32'hbf1b9958, 32'h00000000} /* (19, 14, 11) {real, imag} */,
  {32'h3e0e83b2, 32'h00000000} /* (19, 14, 10) {real, imag} */,
  {32'h3f5c4306, 32'h00000000} /* (19, 14, 9) {real, imag} */,
  {32'h3f9caf40, 32'h00000000} /* (19, 14, 8) {real, imag} */,
  {32'h3f81d928, 32'h00000000} /* (19, 14, 7) {real, imag} */,
  {32'h3f58c588, 32'h00000000} /* (19, 14, 6) {real, imag} */,
  {32'h3f1d8917, 32'h00000000} /* (19, 14, 5) {real, imag} */,
  {32'h3f0fc9d8, 32'h00000000} /* (19, 14, 4) {real, imag} */,
  {32'h3f23cd6c, 32'h00000000} /* (19, 14, 3) {real, imag} */,
  {32'h3f1c8801, 32'h00000000} /* (19, 14, 2) {real, imag} */,
  {32'h3f115b09, 32'h00000000} /* (19, 14, 1) {real, imag} */,
  {32'h3e1783b4, 32'h00000000} /* (19, 14, 0) {real, imag} */,
  {32'h3e92f388, 32'h00000000} /* (19, 13, 31) {real, imag} */,
  {32'h3f806c18, 32'h00000000} /* (19, 13, 30) {real, imag} */,
  {32'h3f6f7cf2, 32'h00000000} /* (19, 13, 29) {real, imag} */,
  {32'h3fb3dbee, 32'h00000000} /* (19, 13, 28) {real, imag} */,
  {32'h3f5b645b, 32'h00000000} /* (19, 13, 27) {real, imag} */,
  {32'h3f2f9142, 32'h00000000} /* (19, 13, 26) {real, imag} */,
  {32'h3f3d28be, 32'h00000000} /* (19, 13, 25) {real, imag} */,
  {32'h3f4142c9, 32'h00000000} /* (19, 13, 24) {real, imag} */,
  {32'h3f288cfe, 32'h00000000} /* (19, 13, 23) {real, imag} */,
  {32'h3f41c776, 32'h00000000} /* (19, 13, 22) {real, imag} */,
  {32'h3f3cdca0, 32'h00000000} /* (19, 13, 21) {real, imag} */,
  {32'hbf8d4142, 32'h00000000} /* (19, 13, 20) {real, imag} */,
  {32'hbf762941, 32'h00000000} /* (19, 13, 19) {real, imag} */,
  {32'hbe936881, 32'h00000000} /* (19, 13, 18) {real, imag} */,
  {32'hbf8b417c, 32'h00000000} /* (19, 13, 17) {real, imag} */,
  {32'hbf86ebda, 32'h00000000} /* (19, 13, 16) {real, imag} */,
  {32'hbf9ec955, 32'h00000000} /* (19, 13, 15) {real, imag} */,
  {32'hbfdb4a4a, 32'h00000000} /* (19, 13, 14) {real, imag} */,
  {32'hbfd46056, 32'h00000000} /* (19, 13, 13) {real, imag} */,
  {32'hbf299429, 32'h00000000} /* (19, 13, 12) {real, imag} */,
  {32'hbe44c032, 32'h00000000} /* (19, 13, 11) {real, imag} */,
  {32'h3eb0e5f3, 32'h00000000} /* (19, 13, 10) {real, imag} */,
  {32'h3f34bc1b, 32'h00000000} /* (19, 13, 9) {real, imag} */,
  {32'h3f86609f, 32'h00000000} /* (19, 13, 8) {real, imag} */,
  {32'h3f57434a, 32'h00000000} /* (19, 13, 7) {real, imag} */,
  {32'h3f32eef0, 32'h00000000} /* (19, 13, 6) {real, imag} */,
  {32'h3f2e6d65, 32'h00000000} /* (19, 13, 5) {real, imag} */,
  {32'h3e862f05, 32'h00000000} /* (19, 13, 4) {real, imag} */,
  {32'h3ec14cfc, 32'h00000000} /* (19, 13, 3) {real, imag} */,
  {32'h3ec75f45, 32'h00000000} /* (19, 13, 2) {real, imag} */,
  {32'h3eb1c7d7, 32'h00000000} /* (19, 13, 1) {real, imag} */,
  {32'h3e915e0d, 32'h00000000} /* (19, 13, 0) {real, imag} */,
  {32'h3d2f0577, 32'h00000000} /* (19, 12, 31) {real, imag} */,
  {32'h3f30f0f6, 32'h00000000} /* (19, 12, 30) {real, imag} */,
  {32'h3f135d10, 32'h00000000} /* (19, 12, 29) {real, imag} */,
  {32'h3f3f4286, 32'h00000000} /* (19, 12, 28) {real, imag} */,
  {32'h3f4a32a6, 32'h00000000} /* (19, 12, 27) {real, imag} */,
  {32'h3f66a5f5, 32'h00000000} /* (19, 12, 26) {real, imag} */,
  {32'h3f073b40, 32'h00000000} /* (19, 12, 25) {real, imag} */,
  {32'h3e2a9de6, 32'h00000000} /* (19, 12, 24) {real, imag} */,
  {32'h3f6d5d46, 32'h00000000} /* (19, 12, 23) {real, imag} */,
  {32'h3fa8d335, 32'h00000000} /* (19, 12, 22) {real, imag} */,
  {32'h3f947458, 32'h00000000} /* (19, 12, 21) {real, imag} */,
  {32'hbeddefe8, 32'h00000000} /* (19, 12, 20) {real, imag} */,
  {32'hbf550495, 32'h00000000} /* (19, 12, 19) {real, imag} */,
  {32'hbf024042, 32'h00000000} /* (19, 12, 18) {real, imag} */,
  {32'hbfbd282d, 32'h00000000} /* (19, 12, 17) {real, imag} */,
  {32'hbf856504, 32'h00000000} /* (19, 12, 16) {real, imag} */,
  {32'hbf9605ed, 32'h00000000} /* (19, 12, 15) {real, imag} */,
  {32'hbfe825e7, 32'h00000000} /* (19, 12, 14) {real, imag} */,
  {32'hbff9452b, 32'h00000000} /* (19, 12, 13) {real, imag} */,
  {32'hbf82e634, 32'h00000000} /* (19, 12, 12) {real, imag} */,
  {32'hbe445536, 32'h00000000} /* (19, 12, 11) {real, imag} */,
  {32'h3f05cda4, 32'h00000000} /* (19, 12, 10) {real, imag} */,
  {32'h3f4f8393, 32'h00000000} /* (19, 12, 9) {real, imag} */,
  {32'h3f889063, 32'h00000000} /* (19, 12, 8) {real, imag} */,
  {32'h3f7d865a, 32'h00000000} /* (19, 12, 7) {real, imag} */,
  {32'h3f34ad47, 32'h00000000} /* (19, 12, 6) {real, imag} */,
  {32'h3f0f14d0, 32'h00000000} /* (19, 12, 5) {real, imag} */,
  {32'h3e91fde6, 32'h00000000} /* (19, 12, 4) {real, imag} */,
  {32'h3f2a4e71, 32'h00000000} /* (19, 12, 3) {real, imag} */,
  {32'h3ee73615, 32'h00000000} /* (19, 12, 2) {real, imag} */,
  {32'h3e9ae829, 32'h00000000} /* (19, 12, 1) {real, imag} */,
  {32'h3d7e250f, 32'h00000000} /* (19, 12, 0) {real, imag} */,
  {32'h3ded3832, 32'h00000000} /* (19, 11, 31) {real, imag} */,
  {32'h3f44a3de, 32'h00000000} /* (19, 11, 30) {real, imag} */,
  {32'h3f0705ae, 32'h00000000} /* (19, 11, 29) {real, imag} */,
  {32'h3f275d78, 32'h00000000} /* (19, 11, 28) {real, imag} */,
  {32'h3ec8d014, 32'h00000000} /* (19, 11, 27) {real, imag} */,
  {32'h3ee1807e, 32'h00000000} /* (19, 11, 26) {real, imag} */,
  {32'h3ef99201, 32'h00000000} /* (19, 11, 25) {real, imag} */,
  {32'h3e8d5b93, 32'h00000000} /* (19, 11, 24) {real, imag} */,
  {32'h3f10237f, 32'h00000000} /* (19, 11, 23) {real, imag} */,
  {32'h3f8d0328, 32'h00000000} /* (19, 11, 22) {real, imag} */,
  {32'h3f1a2936, 32'h00000000} /* (19, 11, 21) {real, imag} */,
  {32'hbee58867, 32'h00000000} /* (19, 11, 20) {real, imag} */,
  {32'hbf29bf68, 32'h00000000} /* (19, 11, 19) {real, imag} */,
  {32'hbf09bd36, 32'h00000000} /* (19, 11, 18) {real, imag} */,
  {32'hbf874409, 32'h00000000} /* (19, 11, 17) {real, imag} */,
  {32'hbe5b3376, 32'h00000000} /* (19, 11, 16) {real, imag} */,
  {32'hbed67c9a, 32'h00000000} /* (19, 11, 15) {real, imag} */,
  {32'hbfaa4cc1, 32'h00000000} /* (19, 11, 14) {real, imag} */,
  {32'hbfaff452, 32'h00000000} /* (19, 11, 13) {real, imag} */,
  {32'hbf31fa54, 32'h00000000} /* (19, 11, 12) {real, imag} */,
  {32'h3e95b351, 32'h00000000} /* (19, 11, 11) {real, imag} */,
  {32'h3f5033fa, 32'h00000000} /* (19, 11, 10) {real, imag} */,
  {32'h3ecb53bd, 32'h00000000} /* (19, 11, 9) {real, imag} */,
  {32'h3ed1d3d6, 32'h00000000} /* (19, 11, 8) {real, imag} */,
  {32'h3efdff57, 32'h00000000} /* (19, 11, 7) {real, imag} */,
  {32'h3f1cd38d, 32'h00000000} /* (19, 11, 6) {real, imag} */,
  {32'h3ea8dead, 32'h00000000} /* (19, 11, 5) {real, imag} */,
  {32'h3e345f6e, 32'h00000000} /* (19, 11, 4) {real, imag} */,
  {32'h3f0ca001, 32'h00000000} /* (19, 11, 3) {real, imag} */,
  {32'h3f339d5f, 32'h00000000} /* (19, 11, 2) {real, imag} */,
  {32'h3ec75fb9, 32'h00000000} /* (19, 11, 1) {real, imag} */,
  {32'h3d9f230f, 32'h00000000} /* (19, 11, 0) {real, imag} */,
  {32'hbeec0094, 32'h00000000} /* (19, 10, 31) {real, imag} */,
  {32'hbea2f488, 32'h00000000} /* (19, 10, 30) {real, imag} */,
  {32'hbe73dd82, 32'h00000000} /* (19, 10, 29) {real, imag} */,
  {32'hbf34b2dd, 32'h00000000} /* (19, 10, 28) {real, imag} */,
  {32'hbf6b7a20, 32'h00000000} /* (19, 10, 27) {real, imag} */,
  {32'hbf479117, 32'h00000000} /* (19, 10, 26) {real, imag} */,
  {32'hbf37c830, 32'h00000000} /* (19, 10, 25) {real, imag} */,
  {32'hbfa16899, 32'h00000000} /* (19, 10, 24) {real, imag} */,
  {32'hbf9900c8, 32'h00000000} /* (19, 10, 23) {real, imag} */,
  {32'hbf15dc1a, 32'h00000000} /* (19, 10, 22) {real, imag} */,
  {32'hbe053e6f, 32'h00000000} /* (19, 10, 21) {real, imag} */,
  {32'h3e915e0a, 32'h00000000} /* (19, 10, 20) {real, imag} */,
  {32'h3f0f121d, 32'h00000000} /* (19, 10, 19) {real, imag} */,
  {32'h3ed8947c, 32'h00000000} /* (19, 10, 18) {real, imag} */,
  {32'h3e826e39, 32'h00000000} /* (19, 10, 17) {real, imag} */,
  {32'h3f890060, 32'h00000000} /* (19, 10, 16) {real, imag} */,
  {32'h3fb495c7, 32'h00000000} /* (19, 10, 15) {real, imag} */,
  {32'h3ed68dd6, 32'h00000000} /* (19, 10, 14) {real, imag} */,
  {32'hbe0a1409, 32'h00000000} /* (19, 10, 13) {real, imag} */,
  {32'h3ef19071, 32'h00000000} /* (19, 10, 12) {real, imag} */,
  {32'h3f09a2f3, 32'h00000000} /* (19, 10, 11) {real, imag} */,
  {32'h3daf5185, 32'h00000000} /* (19, 10, 10) {real, imag} */,
  {32'hbf70ce00, 32'h00000000} /* (19, 10, 9) {real, imag} */,
  {32'hbf1cef49, 32'h00000000} /* (19, 10, 8) {real, imag} */,
  {32'hbea152ea, 32'h00000000} /* (19, 10, 7) {real, imag} */,
  {32'hbf0c2fe3, 32'h00000000} /* (19, 10, 6) {real, imag} */,
  {32'hbf2c3c96, 32'h00000000} /* (19, 10, 5) {real, imag} */,
  {32'hbf03b26d, 32'h00000000} /* (19, 10, 4) {real, imag} */,
  {32'hbed103cb, 32'h00000000} /* (19, 10, 3) {real, imag} */,
  {32'hbecead87, 32'h00000000} /* (19, 10, 2) {real, imag} */,
  {32'hbecff963, 32'h00000000} /* (19, 10, 1) {real, imag} */,
  {32'hbee3344a, 32'h00000000} /* (19, 10, 0) {real, imag} */,
  {32'hbef000da, 32'h00000000} /* (19, 9, 31) {real, imag} */,
  {32'hbf71ac63, 32'h00000000} /* (19, 9, 30) {real, imag} */,
  {32'hbf47ec92, 32'h00000000} /* (19, 9, 29) {real, imag} */,
  {32'hbfbc20b7, 32'h00000000} /* (19, 9, 28) {real, imag} */,
  {32'hbf98876b, 32'h00000000} /* (19, 9, 27) {real, imag} */,
  {32'hbf88c1fe, 32'h00000000} /* (19, 9, 26) {real, imag} */,
  {32'hbf83316d, 32'h00000000} /* (19, 9, 25) {real, imag} */,
  {32'hbfa2adaa, 32'h00000000} /* (19, 9, 24) {real, imag} */,
  {32'hbfab0b6d, 32'h00000000} /* (19, 9, 23) {real, imag} */,
  {32'hbf74b9a7, 32'h00000000} /* (19, 9, 22) {real, imag} */,
  {32'hbea8f4b4, 32'h00000000} /* (19, 9, 21) {real, imag} */,
  {32'h3f4fdfc2, 32'h00000000} /* (19, 9, 20) {real, imag} */,
  {32'h3f504d34, 32'h00000000} /* (19, 9, 19) {real, imag} */,
  {32'h3f900e53, 32'h00000000} /* (19, 9, 18) {real, imag} */,
  {32'h3fc16705, 32'h00000000} /* (19, 9, 17) {real, imag} */,
  {32'h3fc404c6, 32'h00000000} /* (19, 9, 16) {real, imag} */,
  {32'h401c4769, 32'h00000000} /* (19, 9, 15) {real, imag} */,
  {32'h3fc1f111, 32'h00000000} /* (19, 9, 14) {real, imag} */,
  {32'h3ec0cd64, 32'h00000000} /* (19, 9, 13) {real, imag} */,
  {32'h3f50544d, 32'h00000000} /* (19, 9, 12) {real, imag} */,
  {32'h3f13c609, 32'h00000000} /* (19, 9, 11) {real, imag} */,
  {32'hbf53935a, 32'h00000000} /* (19, 9, 10) {real, imag} */,
  {32'hbfd677d0, 32'h00000000} /* (19, 9, 9) {real, imag} */,
  {32'hbf27c162, 32'h00000000} /* (19, 9, 8) {real, imag} */,
  {32'hbf0d5976, 32'h00000000} /* (19, 9, 7) {real, imag} */,
  {32'hbf8eeee6, 32'h00000000} /* (19, 9, 6) {real, imag} */,
  {32'hbf74c43f, 32'h00000000} /* (19, 9, 5) {real, imag} */,
  {32'hbf81f4ab, 32'h00000000} /* (19, 9, 4) {real, imag} */,
  {32'hbf37a6dc, 32'h00000000} /* (19, 9, 3) {real, imag} */,
  {32'hbf26fd63, 32'h00000000} /* (19, 9, 2) {real, imag} */,
  {32'hbf77c58a, 32'h00000000} /* (19, 9, 1) {real, imag} */,
  {32'hbf5103ce, 32'h00000000} /* (19, 9, 0) {real, imag} */,
  {32'hbf2e4b5a, 32'h00000000} /* (19, 8, 31) {real, imag} */,
  {32'hbf8ff69d, 32'h00000000} /* (19, 8, 30) {real, imag} */,
  {32'hbfa1e5d8, 32'h00000000} /* (19, 8, 29) {real, imag} */,
  {32'hbf999360, 32'h00000000} /* (19, 8, 28) {real, imag} */,
  {32'hbf94f07a, 32'h00000000} /* (19, 8, 27) {real, imag} */,
  {32'hbf84f032, 32'h00000000} /* (19, 8, 26) {real, imag} */,
  {32'hbf52cc6e, 32'h00000000} /* (19, 8, 25) {real, imag} */,
  {32'hbf776288, 32'h00000000} /* (19, 8, 24) {real, imag} */,
  {32'hbf8207c0, 32'h00000000} /* (19, 8, 23) {real, imag} */,
  {32'hbf8c0c3f, 32'h00000000} /* (19, 8, 22) {real, imag} */,
  {32'hbf0613dc, 32'h00000000} /* (19, 8, 21) {real, imag} */,
  {32'h3f74ca2c, 32'h00000000} /* (19, 8, 20) {real, imag} */,
  {32'h3f853600, 32'h00000000} /* (19, 8, 19) {real, imag} */,
  {32'h3f849fdc, 32'h00000000} /* (19, 8, 18) {real, imag} */,
  {32'h3f825f67, 32'h00000000} /* (19, 8, 17) {real, imag} */,
  {32'h3f37a809, 32'h00000000} /* (19, 8, 16) {real, imag} */,
  {32'h3fc7baba, 32'h00000000} /* (19, 8, 15) {real, imag} */,
  {32'h3fab02b4, 32'h00000000} /* (19, 8, 14) {real, imag} */,
  {32'h3f13c946, 32'h00000000} /* (19, 8, 13) {real, imag} */,
  {32'h3f1bf3b9, 32'h00000000} /* (19, 8, 12) {real, imag} */,
  {32'h3f56ec8d, 32'h00000000} /* (19, 8, 11) {real, imag} */,
  {32'hbf5b3da2, 32'h00000000} /* (19, 8, 10) {real, imag} */,
  {32'hbf8fa134, 32'h00000000} /* (19, 8, 9) {real, imag} */,
  {32'hbeb7af5d, 32'h00000000} /* (19, 8, 8) {real, imag} */,
  {32'hbf316ff3, 32'h00000000} /* (19, 8, 7) {real, imag} */,
  {32'hbf8d929d, 32'h00000000} /* (19, 8, 6) {real, imag} */,
  {32'hbf0ce864, 32'h00000000} /* (19, 8, 5) {real, imag} */,
  {32'hbf164d0a, 32'h00000000} /* (19, 8, 4) {real, imag} */,
  {32'hbf64d30d, 32'h00000000} /* (19, 8, 3) {real, imag} */,
  {32'hbf3cb660, 32'h00000000} /* (19, 8, 2) {real, imag} */,
  {32'hbf7e3072, 32'h00000000} /* (19, 8, 1) {real, imag} */,
  {32'hbf708a69, 32'h00000000} /* (19, 8, 0) {real, imag} */,
  {32'hbf6fd916, 32'h00000000} /* (19, 7, 31) {real, imag} */,
  {32'hbf830f09, 32'h00000000} /* (19, 7, 30) {real, imag} */,
  {32'hbf91d47e, 32'h00000000} /* (19, 7, 29) {real, imag} */,
  {32'hbf4ff6d6, 32'h00000000} /* (19, 7, 28) {real, imag} */,
  {32'hbf482859, 32'h00000000} /* (19, 7, 27) {real, imag} */,
  {32'hbf5c461b, 32'h00000000} /* (19, 7, 26) {real, imag} */,
  {32'hbfb76a9d, 32'h00000000} /* (19, 7, 25) {real, imag} */,
  {32'hbfd430a2, 32'h00000000} /* (19, 7, 24) {real, imag} */,
  {32'hbf3fd586, 32'h00000000} /* (19, 7, 23) {real, imag} */,
  {32'hbfa11232, 32'h00000000} /* (19, 7, 22) {real, imag} */,
  {32'hbfc97d2a, 32'h00000000} /* (19, 7, 21) {real, imag} */,
  {32'h3eb1abbb, 32'h00000000} /* (19, 7, 20) {real, imag} */,
  {32'h3f95a5e4, 32'h00000000} /* (19, 7, 19) {real, imag} */,
  {32'h3f94f7c1, 32'h00000000} /* (19, 7, 18) {real, imag} */,
  {32'h3f978ebd, 32'h00000000} /* (19, 7, 17) {real, imag} */,
  {32'h3f511165, 32'h00000000} /* (19, 7, 16) {real, imag} */,
  {32'h3fa40a04, 32'h00000000} /* (19, 7, 15) {real, imag} */,
  {32'h3f990ce5, 32'h00000000} /* (19, 7, 14) {real, imag} */,
  {32'h3f0a38ef, 32'h00000000} /* (19, 7, 13) {real, imag} */,
  {32'h3f3abeaa, 32'h00000000} /* (19, 7, 12) {real, imag} */,
  {32'h3f5ca396, 32'h00000000} /* (19, 7, 11) {real, imag} */,
  {32'hbf072832, 32'h00000000} /* (19, 7, 10) {real, imag} */,
  {32'hbf4908a1, 32'h00000000} /* (19, 7, 9) {real, imag} */,
  {32'hbf58be7c, 32'h00000000} /* (19, 7, 8) {real, imag} */,
  {32'hbf83a5ab, 32'h00000000} /* (19, 7, 7) {real, imag} */,
  {32'hbf8c90fe, 32'h00000000} /* (19, 7, 6) {real, imag} */,
  {32'hbf589219, 32'h00000000} /* (19, 7, 5) {real, imag} */,
  {32'hbf34f0e1, 32'h00000000} /* (19, 7, 4) {real, imag} */,
  {32'hbf183848, 32'h00000000} /* (19, 7, 3) {real, imag} */,
  {32'hbf55911c, 32'h00000000} /* (19, 7, 2) {real, imag} */,
  {32'hbf4ca080, 32'h00000000} /* (19, 7, 1) {real, imag} */,
  {32'hbf1fc4e2, 32'h00000000} /* (19, 7, 0) {real, imag} */,
  {32'hbedb0463, 32'h00000000} /* (19, 6, 31) {real, imag} */,
  {32'hbf41f5c0, 32'h00000000} /* (19, 6, 30) {real, imag} */,
  {32'hbf717622, 32'h00000000} /* (19, 6, 29) {real, imag} */,
  {32'hbedd73ee, 32'h00000000} /* (19, 6, 28) {real, imag} */,
  {32'hbdd5ba0f, 32'h00000000} /* (19, 6, 27) {real, imag} */,
  {32'hbf2900f0, 32'h00000000} /* (19, 6, 26) {real, imag} */,
  {32'hbfa33ed6, 32'h00000000} /* (19, 6, 25) {real, imag} */,
  {32'hbf9dfbc0, 32'h00000000} /* (19, 6, 24) {real, imag} */,
  {32'hbee37cf3, 32'h00000000} /* (19, 6, 23) {real, imag} */,
  {32'hbf62cc3d, 32'h00000000} /* (19, 6, 22) {real, imag} */,
  {32'hbf76d29f, 32'h00000000} /* (19, 6, 21) {real, imag} */,
  {32'h3ebc7483, 32'h00000000} /* (19, 6, 20) {real, imag} */,
  {32'h3f61109c, 32'h00000000} /* (19, 6, 19) {real, imag} */,
  {32'h3f6e5286, 32'h00000000} /* (19, 6, 18) {real, imag} */,
  {32'h3f7561bb, 32'h00000000} /* (19, 6, 17) {real, imag} */,
  {32'h3f67e9b7, 32'h00000000} /* (19, 6, 16) {real, imag} */,
  {32'h3f961876, 32'h00000000} /* (19, 6, 15) {real, imag} */,
  {32'h3fbd57c3, 32'h00000000} /* (19, 6, 14) {real, imag} */,
  {32'h3f33b204, 32'h00000000} /* (19, 6, 13) {real, imag} */,
  {32'h3f51de4b, 32'h00000000} /* (19, 6, 12) {real, imag} */,
  {32'h3efd400b, 32'h00000000} /* (19, 6, 11) {real, imag} */,
  {32'hbdfc3a40, 32'h00000000} /* (19, 6, 10) {real, imag} */,
  {32'hbf07e63f, 32'h00000000} /* (19, 6, 9) {real, imag} */,
  {32'hbf6160d3, 32'h00000000} /* (19, 6, 8) {real, imag} */,
  {32'hbf365ab6, 32'h00000000} /* (19, 6, 7) {real, imag} */,
  {32'hbf830bb1, 32'h00000000} /* (19, 6, 6) {real, imag} */,
  {32'hbf76f929, 32'h00000000} /* (19, 6, 5) {real, imag} */,
  {32'hbf450ce2, 32'h00000000} /* (19, 6, 4) {real, imag} */,
  {32'hbf71efcd, 32'h00000000} /* (19, 6, 3) {real, imag} */,
  {32'hbf8f72ed, 32'h00000000} /* (19, 6, 2) {real, imag} */,
  {32'hbf778a7d, 32'h00000000} /* (19, 6, 1) {real, imag} */,
  {32'hbea74c3f, 32'h00000000} /* (19, 6, 0) {real, imag} */,
  {32'hbf275826, 32'h00000000} /* (19, 5, 31) {real, imag} */,
  {32'hbf94e2c6, 32'h00000000} /* (19, 5, 30) {real, imag} */,
  {32'hbfa6615e, 32'h00000000} /* (19, 5, 29) {real, imag} */,
  {32'hbf22ea6b, 32'h00000000} /* (19, 5, 28) {real, imag} */,
  {32'hbedd65d7, 32'h00000000} /* (19, 5, 27) {real, imag} */,
  {32'hbe3153e3, 32'h00000000} /* (19, 5, 26) {real, imag} */,
  {32'hbefcf3c3, 32'h00000000} /* (19, 5, 25) {real, imag} */,
  {32'hbf9e6edc, 32'h00000000} /* (19, 5, 24) {real, imag} */,
  {32'hbf67b2b8, 32'h00000000} /* (19, 5, 23) {real, imag} */,
  {32'hbf13e2b8, 32'h00000000} /* (19, 5, 22) {real, imag} */,
  {32'hbd90a8b8, 32'h00000000} /* (19, 5, 21) {real, imag} */,
  {32'h3e84f325, 32'h00000000} /* (19, 5, 20) {real, imag} */,
  {32'h3d7627cd, 32'h00000000} /* (19, 5, 19) {real, imag} */,
  {32'hbefba19f, 32'h00000000} /* (19, 5, 18) {real, imag} */,
  {32'hbe561fa9, 32'h00000000} /* (19, 5, 17) {real, imag} */,
  {32'h3eb48efd, 32'h00000000} /* (19, 5, 16) {real, imag} */,
  {32'h3f029efc, 32'h00000000} /* (19, 5, 15) {real, imag} */,
  {32'h3f4b74d4, 32'h00000000} /* (19, 5, 14) {real, imag} */,
  {32'h3ed6ad93, 32'h00000000} /* (19, 5, 13) {real, imag} */,
  {32'h3f6685e8, 32'h00000000} /* (19, 5, 12) {real, imag} */,
  {32'h3f8f7986, 32'h00000000} /* (19, 5, 11) {real, imag} */,
  {32'h3f89a492, 32'h00000000} /* (19, 5, 10) {real, imag} */,
  {32'h3ed73ad2, 32'h00000000} /* (19, 5, 9) {real, imag} */,
  {32'h3ec04629, 32'h00000000} /* (19, 5, 8) {real, imag} */,
  {32'h3e91ebf9, 32'h00000000} /* (19, 5, 7) {real, imag} */,
  {32'h3eb16e94, 32'h00000000} /* (19, 5, 6) {real, imag} */,
  {32'hbf26aa7e, 32'h00000000} /* (19, 5, 5) {real, imag} */,
  {32'hbf8727b7, 32'h00000000} /* (19, 5, 4) {real, imag} */,
  {32'hbf8b0b83, 32'h00000000} /* (19, 5, 3) {real, imag} */,
  {32'hbf994c1b, 32'h00000000} /* (19, 5, 2) {real, imag} */,
  {32'hbf8deff4, 32'h00000000} /* (19, 5, 1) {real, imag} */,
  {32'hbe8d5948, 32'h00000000} /* (19, 5, 0) {real, imag} */,
  {32'hbf6ba3f3, 32'h00000000} /* (19, 4, 31) {real, imag} */,
  {32'hbfa0d3e3, 32'h00000000} /* (19, 4, 30) {real, imag} */,
  {32'hbfb11f9c, 32'h00000000} /* (19, 4, 29) {real, imag} */,
  {32'hbf5e8d9f, 32'h00000000} /* (19, 4, 28) {real, imag} */,
  {32'hbf471c2d, 32'h00000000} /* (19, 4, 27) {real, imag} */,
  {32'hbe9f8005, 32'h00000000} /* (19, 4, 26) {real, imag} */,
  {32'hbe599f31, 32'h00000000} /* (19, 4, 25) {real, imag} */,
  {32'hbf8d99b9, 32'h00000000} /* (19, 4, 24) {real, imag} */,
  {32'hbf9effb5, 32'h00000000} /* (19, 4, 23) {real, imag} */,
  {32'hbf66bcdc, 32'h00000000} /* (19, 4, 22) {real, imag} */,
  {32'hbf8d7e34, 32'h00000000} /* (19, 4, 21) {real, imag} */,
  {32'hbf4df61d, 32'h00000000} /* (19, 4, 20) {real, imag} */,
  {32'hbf8267e7, 32'h00000000} /* (19, 4, 19) {real, imag} */,
  {32'hbf9a9f12, 32'h00000000} /* (19, 4, 18) {real, imag} */,
  {32'hbf833f1d, 32'h00000000} /* (19, 4, 17) {real, imag} */,
  {32'hbf084010, 32'h00000000} /* (19, 4, 16) {real, imag} */,
  {32'h3e3de1a2, 32'h00000000} /* (19, 4, 15) {real, imag} */,
  {32'h3f587263, 32'h00000000} /* (19, 4, 14) {real, imag} */,
  {32'h3f17430c, 32'h00000000} /* (19, 4, 13) {real, imag} */,
  {32'h3f51855c, 32'h00000000} /* (19, 4, 12) {real, imag} */,
  {32'h3f9a7e57, 32'h00000000} /* (19, 4, 11) {real, imag} */,
  {32'h3f9f7087, 32'h00000000} /* (19, 4, 10) {real, imag} */,
  {32'h3faf5327, 32'h00000000} /* (19, 4, 9) {real, imag} */,
  {32'h3fc502c1, 32'h00000000} /* (19, 4, 8) {real, imag} */,
  {32'h3f86e521, 32'h00000000} /* (19, 4, 7) {real, imag} */,
  {32'h3f6b7f32, 32'h00000000} /* (19, 4, 6) {real, imag} */,
  {32'hbf27b554, 32'h00000000} /* (19, 4, 5) {real, imag} */,
  {32'hbf99af18, 32'h00000000} /* (19, 4, 4) {real, imag} */,
  {32'hbf649215, 32'h00000000} /* (19, 4, 3) {real, imag} */,
  {32'hbf374fc9, 32'h00000000} /* (19, 4, 2) {real, imag} */,
  {32'hbf431d85, 32'h00000000} /* (19, 4, 1) {real, imag} */,
  {32'hbe7d4e09, 32'h00000000} /* (19, 4, 0) {real, imag} */,
  {32'hbedf697e, 32'h00000000} /* (19, 3, 31) {real, imag} */,
  {32'hbf39c69c, 32'h00000000} /* (19, 3, 30) {real, imag} */,
  {32'hbf248018, 32'h00000000} /* (19, 3, 29) {real, imag} */,
  {32'hbe795c62, 32'h00000000} /* (19, 3, 28) {real, imag} */,
  {32'hbecf3e5c, 32'h00000000} /* (19, 3, 27) {real, imag} */,
  {32'hbf03d31a, 32'h00000000} /* (19, 3, 26) {real, imag} */,
  {32'hbefd75da, 32'h00000000} /* (19, 3, 25) {real, imag} */,
  {32'hbf88da50, 32'h00000000} /* (19, 3, 24) {real, imag} */,
  {32'hbfd7a4b0, 32'h00000000} /* (19, 3, 23) {real, imag} */,
  {32'hbfd4f97e, 32'h00000000} /* (19, 3, 22) {real, imag} */,
  {32'hbf844931, 32'h00000000} /* (19, 3, 21) {real, imag} */,
  {32'hbfa08c8f, 32'h00000000} /* (19, 3, 20) {real, imag} */,
  {32'hbfcc4d8d, 32'h00000000} /* (19, 3, 19) {real, imag} */,
  {32'hbf78accd, 32'h00000000} /* (19, 3, 18) {real, imag} */,
  {32'hbf6ce2dd, 32'h00000000} /* (19, 3, 17) {real, imag} */,
  {32'hbf00ce05, 32'h00000000} /* (19, 3, 16) {real, imag} */,
  {32'h3e0fd3d9, 32'h00000000} /* (19, 3, 15) {real, imag} */,
  {32'h3f21b072, 32'h00000000} /* (19, 3, 14) {real, imag} */,
  {32'h3f6acb69, 32'h00000000} /* (19, 3, 13) {real, imag} */,
  {32'h3f88f6bd, 32'h00000000} /* (19, 3, 12) {real, imag} */,
  {32'h3f6a96f6, 32'h00000000} /* (19, 3, 11) {real, imag} */,
  {32'h3f6e8f51, 32'h00000000} /* (19, 3, 10) {real, imag} */,
  {32'h3fc9e3e6, 32'h00000000} /* (19, 3, 9) {real, imag} */,
  {32'h3fe72d22, 32'h00000000} /* (19, 3, 8) {real, imag} */,
  {32'h3fd49acf, 32'h00000000} /* (19, 3, 7) {real, imag} */,
  {32'h3f71a430, 32'h00000000} /* (19, 3, 6) {real, imag} */,
  {32'hbf005b2c, 32'h00000000} /* (19, 3, 5) {real, imag} */,
  {32'hbf769d13, 32'h00000000} /* (19, 3, 4) {real, imag} */,
  {32'hbf5461c7, 32'h00000000} /* (19, 3, 3) {real, imag} */,
  {32'hbf79adfa, 32'h00000000} /* (19, 3, 2) {real, imag} */,
  {32'hbf863f54, 32'h00000000} /* (19, 3, 1) {real, imag} */,
  {32'hbe7ac1e8, 32'h00000000} /* (19, 3, 0) {real, imag} */,
  {32'hbee1ae83, 32'h00000000} /* (19, 2, 31) {real, imag} */,
  {32'hbf8a970e, 32'h00000000} /* (19, 2, 30) {real, imag} */,
  {32'hbed6d493, 32'h00000000} /* (19, 2, 29) {real, imag} */,
  {32'hbe8558b5, 32'h00000000} /* (19, 2, 28) {real, imag} */,
  {32'hbf12f70e, 32'h00000000} /* (19, 2, 27) {real, imag} */,
  {32'hbeda0e8a, 32'h00000000} /* (19, 2, 26) {real, imag} */,
  {32'hbf08d341, 32'h00000000} /* (19, 2, 25) {real, imag} */,
  {32'hbf66ea04, 32'h00000000} /* (19, 2, 24) {real, imag} */,
  {32'hbffccf25, 32'h00000000} /* (19, 2, 23) {real, imag} */,
  {32'hbfbe3191, 32'h00000000} /* (19, 2, 22) {real, imag} */,
  {32'hbe19e171, 32'h00000000} /* (19, 2, 21) {real, imag} */,
  {32'hbf1fa64c, 32'h00000000} /* (19, 2, 20) {real, imag} */,
  {32'hbfbf30bf, 32'h00000000} /* (19, 2, 19) {real, imag} */,
  {32'hbfd318bd, 32'h00000000} /* (19, 2, 18) {real, imag} */,
  {32'hbf9a8bfb, 32'h00000000} /* (19, 2, 17) {real, imag} */,
  {32'hbeee2840, 32'h00000000} /* (19, 2, 16) {real, imag} */,
  {32'h3da432ee, 32'h00000000} /* (19, 2, 15) {real, imag} */,
  {32'h3ea54211, 32'h00000000} /* (19, 2, 14) {real, imag} */,
  {32'h3f37a3be, 32'h00000000} /* (19, 2, 13) {real, imag} */,
  {32'h3f30598e, 32'h00000000} /* (19, 2, 12) {real, imag} */,
  {32'h3ec3ce91, 32'h00000000} /* (19, 2, 11) {real, imag} */,
  {32'h3f161571, 32'h00000000} /* (19, 2, 10) {real, imag} */,
  {32'h3f9a3b99, 32'h00000000} /* (19, 2, 9) {real, imag} */,
  {32'h3fa1c3a7, 32'h00000000} /* (19, 2, 8) {real, imag} */,
  {32'h3fa2ee35, 32'h00000000} /* (19, 2, 7) {real, imag} */,
  {32'h3f4bf2ea, 32'h00000000} /* (19, 2, 6) {real, imag} */,
  {32'hbca2dabf, 32'h00000000} /* (19, 2, 5) {real, imag} */,
  {32'hbf411203, 32'h00000000} /* (19, 2, 4) {real, imag} */,
  {32'hbfb7d29d, 32'h00000000} /* (19, 2, 3) {real, imag} */,
  {32'hbfc20113, 32'h00000000} /* (19, 2, 2) {real, imag} */,
  {32'hbf9812b2, 32'h00000000} /* (19, 2, 1) {real, imag} */,
  {32'hbe3695fa, 32'h00000000} /* (19, 2, 0) {real, imag} */,
  {32'hbecb2daa, 32'h00000000} /* (19, 1, 31) {real, imag} */,
  {32'hbf33be6b, 32'h00000000} /* (19, 1, 30) {real, imag} */,
  {32'hbf6d3dae, 32'h00000000} /* (19, 1, 29) {real, imag} */,
  {32'hbf755272, 32'h00000000} /* (19, 1, 28) {real, imag} */,
  {32'hbf31e5b3, 32'h00000000} /* (19, 1, 27) {real, imag} */,
  {32'hbf04c5e5, 32'h00000000} /* (19, 1, 26) {real, imag} */,
  {32'hbf05d03f, 32'h00000000} /* (19, 1, 25) {real, imag} */,
  {32'hbf4830f5, 32'h00000000} /* (19, 1, 24) {real, imag} */,
  {32'hbfacaa3a, 32'h00000000} /* (19, 1, 23) {real, imag} */,
  {32'hbf58389e, 32'h00000000} /* (19, 1, 22) {real, imag} */,
  {32'hbeb80eb4, 32'h00000000} /* (19, 1, 21) {real, imag} */,
  {32'hbec95487, 32'h00000000} /* (19, 1, 20) {real, imag} */,
  {32'hbf5ef1ea, 32'h00000000} /* (19, 1, 19) {real, imag} */,
  {32'hbfce50dd, 32'h00000000} /* (19, 1, 18) {real, imag} */,
  {32'hbfd41ad4, 32'h00000000} /* (19, 1, 17) {real, imag} */,
  {32'hbe83c12e, 32'h00000000} /* (19, 1, 16) {real, imag} */,
  {32'h3f264775, 32'h00000000} /* (19, 1, 15) {real, imag} */,
  {32'h3ec86cc4, 32'h00000000} /* (19, 1, 14) {real, imag} */,
  {32'h3e8ac489, 32'h00000000} /* (19, 1, 13) {real, imag} */,
  {32'h3ef8c960, 32'h00000000} /* (19, 1, 12) {real, imag} */,
  {32'h3f48f280, 32'h00000000} /* (19, 1, 11) {real, imag} */,
  {32'h3f55a70a, 32'h00000000} /* (19, 1, 10) {real, imag} */,
  {32'h3f7783aa, 32'h00000000} /* (19, 1, 9) {real, imag} */,
  {32'h3f60778b, 32'h00000000} /* (19, 1, 8) {real, imag} */,
  {32'h3f5c207d, 32'h00000000} /* (19, 1, 7) {real, imag} */,
  {32'h3f4a6827, 32'h00000000} /* (19, 1, 6) {real, imag} */,
  {32'h3ec1dfd1, 32'h00000000} /* (19, 1, 5) {real, imag} */,
  {32'hbf535ad5, 32'h00000000} /* (19, 1, 4) {real, imag} */,
  {32'hbfdb798b, 32'h00000000} /* (19, 1, 3) {real, imag} */,
  {32'hbf9a231f, 32'h00000000} /* (19, 1, 2) {real, imag} */,
  {32'hbf87aac1, 32'h00000000} /* (19, 1, 1) {real, imag} */,
  {32'hbee2bb68, 32'h00000000} /* (19, 1, 0) {real, imag} */,
  {32'hbf1ba9b6, 32'h00000000} /* (19, 0, 31) {real, imag} */,
  {32'hbed186d8, 32'h00000000} /* (19, 0, 30) {real, imag} */,
  {32'hbed10c21, 32'h00000000} /* (19, 0, 29) {real, imag} */,
  {32'hbf2454a9, 32'h00000000} /* (19, 0, 28) {real, imag} */,
  {32'hbecb988f, 32'h00000000} /* (19, 0, 27) {real, imag} */,
  {32'hbed35589, 32'h00000000} /* (19, 0, 26) {real, imag} */,
  {32'hbee27312, 32'h00000000} /* (19, 0, 25) {real, imag} */,
  {32'hbec6bf87, 32'h00000000} /* (19, 0, 24) {real, imag} */,
  {32'hbea11e29, 32'h00000000} /* (19, 0, 23) {real, imag} */,
  {32'hbe8e519c, 32'h00000000} /* (19, 0, 22) {real, imag} */,
  {32'hbee11919, 32'h00000000} /* (19, 0, 21) {real, imag} */,
  {32'hbea88a8c, 32'h00000000} /* (19, 0, 20) {real, imag} */,
  {32'hbe6ccd17, 32'h00000000} /* (19, 0, 19) {real, imag} */,
  {32'hbe794577, 32'h00000000} /* (19, 0, 18) {real, imag} */,
  {32'hbf0ef822, 32'h00000000} /* (19, 0, 17) {real, imag} */,
  {32'h3cac897d, 32'h00000000} /* (19, 0, 16) {real, imag} */,
  {32'h3f09bebb, 32'h00000000} /* (19, 0, 15) {real, imag} */,
  {32'h3e29a1e0, 32'h00000000} /* (19, 0, 14) {real, imag} */,
  {32'h3de3dfec, 32'h00000000} /* (19, 0, 13) {real, imag} */,
  {32'h3ec675c0, 32'h00000000} /* (19, 0, 12) {real, imag} */,
  {32'h3f3126d3, 32'h00000000} /* (19, 0, 11) {real, imag} */,
  {32'h3f112c63, 32'h00000000} /* (19, 0, 10) {real, imag} */,
  {32'h3f164add, 32'h00000000} /* (19, 0, 9) {real, imag} */,
  {32'h3f0a95d8, 32'h00000000} /* (19, 0, 8) {real, imag} */,
  {32'h3f184141, 32'h00000000} /* (19, 0, 7) {real, imag} */,
  {32'h3f073bbc, 32'h00000000} /* (19, 0, 6) {real, imag} */,
  {32'hbd1c63a2, 32'h00000000} /* (19, 0, 5) {real, imag} */,
  {32'hbecd98a0, 32'h00000000} /* (19, 0, 4) {real, imag} */,
  {32'hbf276070, 32'h00000000} /* (19, 0, 3) {real, imag} */,
  {32'hbec9a51e, 32'h00000000} /* (19, 0, 2) {real, imag} */,
  {32'hbf5df0ee, 32'h00000000} /* (19, 0, 1) {real, imag} */,
  {32'hbf2e2825, 32'h00000000} /* (19, 0, 0) {real, imag} */,
  {32'hbee129f5, 32'h00000000} /* (18, 31, 31) {real, imag} */,
  {32'hbf385ac8, 32'h00000000} /* (18, 31, 30) {real, imag} */,
  {32'hbf71ab6d, 32'h00000000} /* (18, 31, 29) {real, imag} */,
  {32'hbf4e9c6f, 32'h00000000} /* (18, 31, 28) {real, imag} */,
  {32'hbf452f54, 32'h00000000} /* (18, 31, 27) {real, imag} */,
  {32'hbf6284e3, 32'h00000000} /* (18, 31, 26) {real, imag} */,
  {32'hbf2d8ffa, 32'h00000000} /* (18, 31, 25) {real, imag} */,
  {32'hbe99e421, 32'h00000000} /* (18, 31, 24) {real, imag} */,
  {32'hbe4a3ef7, 32'h00000000} /* (18, 31, 23) {real, imag} */,
  {32'hbea35b84, 32'h00000000} /* (18, 31, 22) {real, imag} */,
  {32'hbeafdae3, 32'h00000000} /* (18, 31, 21) {real, imag} */,
  {32'hbd3fbcd7, 32'h00000000} /* (18, 31, 20) {real, imag} */,
  {32'h3deffa12, 32'h00000000} /* (18, 31, 19) {real, imag} */,
  {32'h3ed2aa68, 32'h00000000} /* (18, 31, 18) {real, imag} */,
  {32'h3eda452f, 32'h00000000} /* (18, 31, 17) {real, imag} */,
  {32'h3e60d8df, 32'h00000000} /* (18, 31, 16) {real, imag} */,
  {32'h3f10cb14, 32'h00000000} /* (18, 31, 15) {real, imag} */,
  {32'h3f01215a, 32'h00000000} /* (18, 31, 14) {real, imag} */,
  {32'h3ea2ba00, 32'h00000000} /* (18, 31, 13) {real, imag} */,
  {32'h3e962017, 32'h00000000} /* (18, 31, 12) {real, imag} */,
  {32'h3f02da57, 32'h00000000} /* (18, 31, 11) {real, imag} */,
  {32'h3dfb0055, 32'h00000000} /* (18, 31, 10) {real, imag} */,
  {32'hbf18f5ad, 32'h00000000} /* (18, 31, 9) {real, imag} */,
  {32'hbf6c5e21, 32'h00000000} /* (18, 31, 8) {real, imag} */,
  {32'hbec6d58b, 32'h00000000} /* (18, 31, 7) {real, imag} */,
  {32'hbed6fc44, 32'h00000000} /* (18, 31, 6) {real, imag} */,
  {32'hbf149586, 32'h00000000} /* (18, 31, 5) {real, imag} */,
  {32'hbe90e872, 32'h00000000} /* (18, 31, 4) {real, imag} */,
  {32'hbf3c490e, 32'h00000000} /* (18, 31, 3) {real, imag} */,
  {32'hbf3f7da5, 32'h00000000} /* (18, 31, 2) {real, imag} */,
  {32'hbf0cd20c, 32'h00000000} /* (18, 31, 1) {real, imag} */,
  {32'hbe89aa35, 32'h00000000} /* (18, 31, 0) {real, imag} */,
  {32'hbf6a682d, 32'h00000000} /* (18, 30, 31) {real, imag} */,
  {32'hbfc99e43, 32'h00000000} /* (18, 30, 30) {real, imag} */,
  {32'hbff9d091, 32'h00000000} /* (18, 30, 29) {real, imag} */,
  {32'hbf999d12, 32'h00000000} /* (18, 30, 28) {real, imag} */,
  {32'hbfa1a688, 32'h00000000} /* (18, 30, 27) {real, imag} */,
  {32'hbfc4f1cf, 32'h00000000} /* (18, 30, 26) {real, imag} */,
  {32'hbf3c74c7, 32'h00000000} /* (18, 30, 25) {real, imag} */,
  {32'hbf205d09, 32'h00000000} /* (18, 30, 24) {real, imag} */,
  {32'hbec07584, 32'h00000000} /* (18, 30, 23) {real, imag} */,
  {32'hbf430946, 32'h00000000} /* (18, 30, 22) {real, imag} */,
  {32'hbf2ee1df, 32'h00000000} /* (18, 30, 21) {real, imag} */,
  {32'h3f22285f, 32'h00000000} /* (18, 30, 20) {real, imag} */,
  {32'h3f327eec, 32'h00000000} /* (18, 30, 19) {real, imag} */,
  {32'h3f18d596, 32'h00000000} /* (18, 30, 18) {real, imag} */,
  {32'h3f50121a, 32'h00000000} /* (18, 30, 17) {real, imag} */,
  {32'h3f53cc43, 32'h00000000} /* (18, 30, 16) {real, imag} */,
  {32'h3f966031, 32'h00000000} /* (18, 30, 15) {real, imag} */,
  {32'h3fac4ca7, 32'h00000000} /* (18, 30, 14) {real, imag} */,
  {32'h3f9b000d, 32'h00000000} /* (18, 30, 13) {real, imag} */,
  {32'h3f6d15cc, 32'h00000000} /* (18, 30, 12) {real, imag} */,
  {32'h3f62ab52, 32'h00000000} /* (18, 30, 11) {real, imag} */,
  {32'h3e866fce, 32'h00000000} /* (18, 30, 10) {real, imag} */,
  {32'hbf755440, 32'h00000000} /* (18, 30, 9) {real, imag} */,
  {32'hbfa5a30e, 32'h00000000} /* (18, 30, 8) {real, imag} */,
  {32'hbf4c2e28, 32'h00000000} /* (18, 30, 7) {real, imag} */,
  {32'hbf5e9cf7, 32'h00000000} /* (18, 30, 6) {real, imag} */,
  {32'hbf189788, 32'h00000000} /* (18, 30, 5) {real, imag} */,
  {32'hbf6fa05b, 32'h00000000} /* (18, 30, 4) {real, imag} */,
  {32'hbf85e327, 32'h00000000} /* (18, 30, 3) {real, imag} */,
  {32'hbf60566e, 32'h00000000} /* (18, 30, 2) {real, imag} */,
  {32'hbf145a17, 32'h00000000} /* (18, 30, 1) {real, imag} */,
  {32'hbeb87653, 32'h00000000} /* (18, 30, 0) {real, imag} */,
  {32'hbf6b5fce, 32'h00000000} /* (18, 29, 31) {real, imag} */,
  {32'hbfca497f, 32'h00000000} /* (18, 29, 30) {real, imag} */,
  {32'hbfb2d17a, 32'h00000000} /* (18, 29, 29) {real, imag} */,
  {32'hbf2c3270, 32'h00000000} /* (18, 29, 28) {real, imag} */,
  {32'hbf224e00, 32'h00000000} /* (18, 29, 27) {real, imag} */,
  {32'hbf661654, 32'h00000000} /* (18, 29, 26) {real, imag} */,
  {32'hbf803efd, 32'h00000000} /* (18, 29, 25) {real, imag} */,
  {32'hbfa808f9, 32'h00000000} /* (18, 29, 24) {real, imag} */,
  {32'hbf5824ca, 32'h00000000} /* (18, 29, 23) {real, imag} */,
  {32'hbf2d4ace, 32'h00000000} /* (18, 29, 22) {real, imag} */,
  {32'hbef918b5, 32'h00000000} /* (18, 29, 21) {real, imag} */,
  {32'h3f4d4863, 32'h00000000} /* (18, 29, 20) {real, imag} */,
  {32'h3f139a0d, 32'h00000000} /* (18, 29, 19) {real, imag} */,
  {32'h3f1b9939, 32'h00000000} /* (18, 29, 18) {real, imag} */,
  {32'h3f8c523d, 32'h00000000} /* (18, 29, 17) {real, imag} */,
  {32'h3fb5200c, 32'h00000000} /* (18, 29, 16) {real, imag} */,
  {32'h3f93204e, 32'h00000000} /* (18, 29, 15) {real, imag} */,
  {32'h3f5d6d6e, 32'h00000000} /* (18, 29, 14) {real, imag} */,
  {32'h3f8b6e48, 32'h00000000} /* (18, 29, 13) {real, imag} */,
  {32'h3f7a5b1c, 32'h00000000} /* (18, 29, 12) {real, imag} */,
  {32'h3f300445, 32'h00000000} /* (18, 29, 11) {real, imag} */,
  {32'h3d91094f, 32'h00000000} /* (18, 29, 10) {real, imag} */,
  {32'hbf12f0c2, 32'h00000000} /* (18, 29, 9) {real, imag} */,
  {32'hbf9ec12d, 32'h00000000} /* (18, 29, 8) {real, imag} */,
  {32'hbf970327, 32'h00000000} /* (18, 29, 7) {real, imag} */,
  {32'hbf4dd3be, 32'h00000000} /* (18, 29, 6) {real, imag} */,
  {32'hbf2a1d71, 32'h00000000} /* (18, 29, 5) {real, imag} */,
  {32'hbf9ba3f0, 32'h00000000} /* (18, 29, 4) {real, imag} */,
  {32'hbfa691c7, 32'h00000000} /* (18, 29, 3) {real, imag} */,
  {32'hbf01421c, 32'h00000000} /* (18, 29, 2) {real, imag} */,
  {32'hbf222e5d, 32'h00000000} /* (18, 29, 1) {real, imag} */,
  {32'hbf5f3c8b, 32'h00000000} /* (18, 29, 0) {real, imag} */,
  {32'hbeded7e2, 32'h00000000} /* (18, 28, 31) {real, imag} */,
  {32'hbf59341e, 32'h00000000} /* (18, 28, 30) {real, imag} */,
  {32'hbf80832f, 32'h00000000} /* (18, 28, 29) {real, imag} */,
  {32'hbf8dfec5, 32'h00000000} /* (18, 28, 28) {real, imag} */,
  {32'hbf2a8710, 32'h00000000} /* (18, 28, 27) {real, imag} */,
  {32'hbf4a3bbf, 32'h00000000} /* (18, 28, 26) {real, imag} */,
  {32'hbfd273e1, 32'h00000000} /* (18, 28, 25) {real, imag} */,
  {32'hbffd1cd5, 32'h00000000} /* (18, 28, 24) {real, imag} */,
  {32'hbf960608, 32'h00000000} /* (18, 28, 23) {real, imag} */,
  {32'hbf367a32, 32'h00000000} /* (18, 28, 22) {real, imag} */,
  {32'hbef22c25, 32'h00000000} /* (18, 28, 21) {real, imag} */,
  {32'h3eba5dfc, 32'h00000000} /* (18, 28, 20) {real, imag} */,
  {32'h3eeeb86c, 32'h00000000} /* (18, 28, 19) {real, imag} */,
  {32'h3f79ea55, 32'h00000000} /* (18, 28, 18) {real, imag} */,
  {32'h3f9cf740, 32'h00000000} /* (18, 28, 17) {real, imag} */,
  {32'h3fa4e88f, 32'h00000000} /* (18, 28, 16) {real, imag} */,
  {32'h3f866545, 32'h00000000} /* (18, 28, 15) {real, imag} */,
  {32'h3f73bd8a, 32'h00000000} /* (18, 28, 14) {real, imag} */,
  {32'h3f3cc422, 32'h00000000} /* (18, 28, 13) {real, imag} */,
  {32'h3f823352, 32'h00000000} /* (18, 28, 12) {real, imag} */,
  {32'h3f8cdeb0, 32'h00000000} /* (18, 28, 11) {real, imag} */,
  {32'hbe7618bc, 32'h00000000} /* (18, 28, 10) {real, imag} */,
  {32'hbf2dd696, 32'h00000000} /* (18, 28, 9) {real, imag} */,
  {32'hbf1597cf, 32'h00000000} /* (18, 28, 8) {real, imag} */,
  {32'hbf8b4d65, 32'h00000000} /* (18, 28, 7) {real, imag} */,
  {32'hbf983535, 32'h00000000} /* (18, 28, 6) {real, imag} */,
  {32'hbf801340, 32'h00000000} /* (18, 28, 5) {real, imag} */,
  {32'hbf8011c0, 32'h00000000} /* (18, 28, 4) {real, imag} */,
  {32'hbf7f12eb, 32'h00000000} /* (18, 28, 3) {real, imag} */,
  {32'hbf564f3f, 32'h00000000} /* (18, 28, 2) {real, imag} */,
  {32'hbf816c86, 32'h00000000} /* (18, 28, 1) {real, imag} */,
  {32'hbf3f3661, 32'h00000000} /* (18, 28, 0) {real, imag} */,
  {32'hbf1303eb, 32'h00000000} /* (18, 27, 31) {real, imag} */,
  {32'hbf55d4b8, 32'h00000000} /* (18, 27, 30) {real, imag} */,
  {32'hbf118f9f, 32'h00000000} /* (18, 27, 29) {real, imag} */,
  {32'hbef7c5e5, 32'h00000000} /* (18, 27, 28) {real, imag} */,
  {32'hbecd809a, 32'h00000000} /* (18, 27, 27) {real, imag} */,
  {32'hbf998163, 32'h00000000} /* (18, 27, 26) {real, imag} */,
  {32'hbfdeeb9c, 32'h00000000} /* (18, 27, 25) {real, imag} */,
  {32'hbf9c6b24, 32'h00000000} /* (18, 27, 24) {real, imag} */,
  {32'hbf53b0ae, 32'h00000000} /* (18, 27, 23) {real, imag} */,
  {32'hbf1483f5, 32'h00000000} /* (18, 27, 22) {real, imag} */,
  {32'hbef39f28, 32'h00000000} /* (18, 27, 21) {real, imag} */,
  {32'h3e52a451, 32'h00000000} /* (18, 27, 20) {real, imag} */,
  {32'h3f069ac8, 32'h00000000} /* (18, 27, 19) {real, imag} */,
  {32'h3f58ad47, 32'h00000000} /* (18, 27, 18) {real, imag} */,
  {32'h3f90230f, 32'h00000000} /* (18, 27, 17) {real, imag} */,
  {32'h3f89da8c, 32'h00000000} /* (18, 27, 16) {real, imag} */,
  {32'h3f69dc5f, 32'h00000000} /* (18, 27, 15) {real, imag} */,
  {32'h3fc1c150, 32'h00000000} /* (18, 27, 14) {real, imag} */,
  {32'h3f87a8fa, 32'h00000000} /* (18, 27, 13) {real, imag} */,
  {32'h3f47d627, 32'h00000000} /* (18, 27, 12) {real, imag} */,
  {32'h3f2e69e8, 32'h00000000} /* (18, 27, 11) {real, imag} */,
  {32'hbf1f0d7c, 32'h00000000} /* (18, 27, 10) {real, imag} */,
  {32'hbf874427, 32'h00000000} /* (18, 27, 9) {real, imag} */,
  {32'hbf6159d9, 32'h00000000} /* (18, 27, 8) {real, imag} */,
  {32'hbf8481a2, 32'h00000000} /* (18, 27, 7) {real, imag} */,
  {32'hbf9c1028, 32'h00000000} /* (18, 27, 6) {real, imag} */,
  {32'hbfe028ce, 32'h00000000} /* (18, 27, 5) {real, imag} */,
  {32'hbfd650f9, 32'h00000000} /* (18, 27, 4) {real, imag} */,
  {32'hbf5bae49, 32'h00000000} /* (18, 27, 3) {real, imag} */,
  {32'hbf468e2e, 32'h00000000} /* (18, 27, 2) {real, imag} */,
  {32'hbf983f5a, 32'h00000000} /* (18, 27, 1) {real, imag} */,
  {32'hbef65ad1, 32'h00000000} /* (18, 27, 0) {real, imag} */,
  {32'hbf1790e1, 32'h00000000} /* (18, 26, 31) {real, imag} */,
  {32'hbf3fc2a2, 32'h00000000} /* (18, 26, 30) {real, imag} */,
  {32'hbede6ed1, 32'h00000000} /* (18, 26, 29) {real, imag} */,
  {32'hbeb9ddb7, 32'h00000000} /* (18, 26, 28) {real, imag} */,
  {32'hbeeeeba7, 32'h00000000} /* (18, 26, 27) {real, imag} */,
  {32'hbf9dd3ba, 32'h00000000} /* (18, 26, 26) {real, imag} */,
  {32'hbfb4b8cf, 32'h00000000} /* (18, 26, 25) {real, imag} */,
  {32'hbf5e0d71, 32'h00000000} /* (18, 26, 24) {real, imag} */,
  {32'hbf39cfee, 32'h00000000} /* (18, 26, 23) {real, imag} */,
  {32'hbf2eb866, 32'h00000000} /* (18, 26, 22) {real, imag} */,
  {32'hbf285647, 32'h00000000} /* (18, 26, 21) {real, imag} */,
  {32'h3e1b70a2, 32'h00000000} /* (18, 26, 20) {real, imag} */,
  {32'h3f2384c9, 32'h00000000} /* (18, 26, 19) {real, imag} */,
  {32'h3eb6851b, 32'h00000000} /* (18, 26, 18) {real, imag} */,
  {32'h3efb204f, 32'h00000000} /* (18, 26, 17) {real, imag} */,
  {32'h3f83e2fe, 32'h00000000} /* (18, 26, 16) {real, imag} */,
  {32'h3f503269, 32'h00000000} /* (18, 26, 15) {real, imag} */,
  {32'h3fabce6e, 32'h00000000} /* (18, 26, 14) {real, imag} */,
  {32'h3f96f666, 32'h00000000} /* (18, 26, 13) {real, imag} */,
  {32'h3f808eae, 32'h00000000} /* (18, 26, 12) {real, imag} */,
  {32'h3f0dd10b, 32'h00000000} /* (18, 26, 11) {real, imag} */,
  {32'hbf17fb99, 32'h00000000} /* (18, 26, 10) {real, imag} */,
  {32'hbf4d016f, 32'h00000000} /* (18, 26, 9) {real, imag} */,
  {32'hbfb02b85, 32'h00000000} /* (18, 26, 8) {real, imag} */,
  {32'hbf88c3e8, 32'h00000000} /* (18, 26, 7) {real, imag} */,
  {32'hbf4e5900, 32'h00000000} /* (18, 26, 6) {real, imag} */,
  {32'hbfc48488, 32'h00000000} /* (18, 26, 5) {real, imag} */,
  {32'hbfbae3ce, 32'h00000000} /* (18, 26, 4) {real, imag} */,
  {32'hbf8471e2, 32'h00000000} /* (18, 26, 3) {real, imag} */,
  {32'hbf9d6bb4, 32'h00000000} /* (18, 26, 2) {real, imag} */,
  {32'hbfc47af8, 32'h00000000} /* (18, 26, 1) {real, imag} */,
  {32'hbf32659e, 32'h00000000} /* (18, 26, 0) {real, imag} */,
  {32'hbf02d9d0, 32'h00000000} /* (18, 25, 31) {real, imag} */,
  {32'hbf2e54b0, 32'h00000000} /* (18, 25, 30) {real, imag} */,
  {32'hbf16647d, 32'h00000000} /* (18, 25, 29) {real, imag} */,
  {32'hbf2979fe, 32'h00000000} /* (18, 25, 28) {real, imag} */,
  {32'hbfbd83a5, 32'h00000000} /* (18, 25, 27) {real, imag} */,
  {32'hbfecefc0, 32'h00000000} /* (18, 25, 26) {real, imag} */,
  {32'hbf65bf80, 32'h00000000} /* (18, 25, 25) {real, imag} */,
  {32'hbf117e75, 32'h00000000} /* (18, 25, 24) {real, imag} */,
  {32'hbf40be98, 32'h00000000} /* (18, 25, 23) {real, imag} */,
  {32'hbf35ca2d, 32'h00000000} /* (18, 25, 22) {real, imag} */,
  {32'hbf4ec311, 32'h00000000} /* (18, 25, 21) {real, imag} */,
  {32'h3fb0c87a, 32'h00000000} /* (18, 25, 20) {real, imag} */,
  {32'h4009a423, 32'h00000000} /* (18, 25, 19) {real, imag} */,
  {32'h3ee98384, 32'h00000000} /* (18, 25, 18) {real, imag} */,
  {32'h3e3cc4b7, 32'h00000000} /* (18, 25, 17) {real, imag} */,
  {32'h3f0f79f2, 32'h00000000} /* (18, 25, 16) {real, imag} */,
  {32'h3f0eb793, 32'h00000000} /* (18, 25, 15) {real, imag} */,
  {32'h3f2c06ad, 32'h00000000} /* (18, 25, 14) {real, imag} */,
  {32'h3f6a4960, 32'h00000000} /* (18, 25, 13) {real, imag} */,
  {32'h3fb150d6, 32'h00000000} /* (18, 25, 12) {real, imag} */,
  {32'h3f48fd79, 32'h00000000} /* (18, 25, 11) {real, imag} */,
  {32'hbf26672b, 32'h00000000} /* (18, 25, 10) {real, imag} */,
  {32'hbf6e42c5, 32'h00000000} /* (18, 25, 9) {real, imag} */,
  {32'hbfb8d55a, 32'h00000000} /* (18, 25, 8) {real, imag} */,
  {32'hbf99061a, 32'h00000000} /* (18, 25, 7) {real, imag} */,
  {32'hbef43fb1, 32'h00000000} /* (18, 25, 6) {real, imag} */,
  {32'hbf005d7e, 32'h00000000} /* (18, 25, 5) {real, imag} */,
  {32'hbf442e7c, 32'h00000000} /* (18, 25, 4) {real, imag} */,
  {32'hbf6363a2, 32'h00000000} /* (18, 25, 3) {real, imag} */,
  {32'hbf9b7e0a, 32'h00000000} /* (18, 25, 2) {real, imag} */,
  {32'hbfc96265, 32'h00000000} /* (18, 25, 1) {real, imag} */,
  {32'hbf158111, 32'h00000000} /* (18, 25, 0) {real, imag} */,
  {32'hbedf3716, 32'h00000000} /* (18, 24, 31) {real, imag} */,
  {32'hbefa9ef9, 32'h00000000} /* (18, 24, 30) {real, imag} */,
  {32'hbf0b83c2, 32'h00000000} /* (18, 24, 29) {real, imag} */,
  {32'hbf7215ed, 32'h00000000} /* (18, 24, 28) {real, imag} */,
  {32'hbf88a8e2, 32'h00000000} /* (18, 24, 27) {real, imag} */,
  {32'hbf9f8bac, 32'h00000000} /* (18, 24, 26) {real, imag} */,
  {32'hbf3d4160, 32'h00000000} /* (18, 24, 25) {real, imag} */,
  {32'hbf486037, 32'h00000000} /* (18, 24, 24) {real, imag} */,
  {32'hbf64e157, 32'h00000000} /* (18, 24, 23) {real, imag} */,
  {32'hbf834ddd, 32'h00000000} /* (18, 24, 22) {real, imag} */,
  {32'hbecf2f2d, 32'h00000000} /* (18, 24, 21) {real, imag} */,
  {32'h3fd85f6d, 32'h00000000} /* (18, 24, 20) {real, imag} */,
  {32'h3fecc858, 32'h00000000} /* (18, 24, 19) {real, imag} */,
  {32'h3f0f564e, 32'h00000000} /* (18, 24, 18) {real, imag} */,
  {32'h3f23326e, 32'h00000000} /* (18, 24, 17) {real, imag} */,
  {32'h3ef5013a, 32'h00000000} /* (18, 24, 16) {real, imag} */,
  {32'h3ed3c681, 32'h00000000} /* (18, 24, 15) {real, imag} */,
  {32'h3ee6a53d, 32'h00000000} /* (18, 24, 14) {real, imag} */,
  {32'h3f23d243, 32'h00000000} /* (18, 24, 13) {real, imag} */,
  {32'h3f1df034, 32'h00000000} /* (18, 24, 12) {real, imag} */,
  {32'h3ebaea64, 32'h00000000} /* (18, 24, 11) {real, imag} */,
  {32'hbf7738ce, 32'h00000000} /* (18, 24, 10) {real, imag} */,
  {32'hbf89ce69, 32'h00000000} /* (18, 24, 9) {real, imag} */,
  {32'hbf96c69b, 32'h00000000} /* (18, 24, 8) {real, imag} */,
  {32'hbf9bb590, 32'h00000000} /* (18, 24, 7) {real, imag} */,
  {32'hbf15ae37, 32'h00000000} /* (18, 24, 6) {real, imag} */,
  {32'hbe81b2ff, 32'h00000000} /* (18, 24, 5) {real, imag} */,
  {32'hbf3c14b8, 32'h00000000} /* (18, 24, 4) {real, imag} */,
  {32'hbf71fbdf, 32'h00000000} /* (18, 24, 3) {real, imag} */,
  {32'hbf8de834, 32'h00000000} /* (18, 24, 2) {real, imag} */,
  {32'hbf90ff35, 32'h00000000} /* (18, 24, 1) {real, imag} */,
  {32'hbec4e0f7, 32'h00000000} /* (18, 24, 0) {real, imag} */,
  {32'hbe4b3d80, 32'h00000000} /* (18, 23, 31) {real, imag} */,
  {32'hbea74e44, 32'h00000000} /* (18, 23, 30) {real, imag} */,
  {32'hbf29b504, 32'h00000000} /* (18, 23, 29) {real, imag} */,
  {32'hbfa04135, 32'h00000000} /* (18, 23, 28) {real, imag} */,
  {32'hbf39a2bf, 32'h00000000} /* (18, 23, 27) {real, imag} */,
  {32'hbf02de86, 32'h00000000} /* (18, 23, 26) {real, imag} */,
  {32'hbf13ca6b, 32'h00000000} /* (18, 23, 25) {real, imag} */,
  {32'hbf868c30, 32'h00000000} /* (18, 23, 24) {real, imag} */,
  {32'hbf8875f8, 32'h00000000} /* (18, 23, 23) {real, imag} */,
  {32'hbf8e892b, 32'h00000000} /* (18, 23, 22) {real, imag} */,
  {32'hbe843b65, 32'h00000000} /* (18, 23, 21) {real, imag} */,
  {32'h3f8ec15d, 32'h00000000} /* (18, 23, 20) {real, imag} */,
  {32'h3f84d015, 32'h00000000} /* (18, 23, 19) {real, imag} */,
  {32'h3f48f098, 32'h00000000} /* (18, 23, 18) {real, imag} */,
  {32'h3fa19a66, 32'h00000000} /* (18, 23, 17) {real, imag} */,
  {32'h3f9ca8e3, 32'h00000000} /* (18, 23, 16) {real, imag} */,
  {32'h3f5ef052, 32'h00000000} /* (18, 23, 15) {real, imag} */,
  {32'h3f1797b0, 32'h00000000} /* (18, 23, 14) {real, imag} */,
  {32'h3f281e18, 32'h00000000} /* (18, 23, 13) {real, imag} */,
  {32'h3f573463, 32'h00000000} /* (18, 23, 12) {real, imag} */,
  {32'h3e5e5d3f, 32'h00000000} /* (18, 23, 11) {real, imag} */,
  {32'hbf5e11e8, 32'h00000000} /* (18, 23, 10) {real, imag} */,
  {32'hbf4cbc90, 32'h00000000} /* (18, 23, 9) {real, imag} */,
  {32'hbf43f898, 32'h00000000} /* (18, 23, 8) {real, imag} */,
  {32'hbf5c43b6, 32'h00000000} /* (18, 23, 7) {real, imag} */,
  {32'hbf26a733, 32'h00000000} /* (18, 23, 6) {real, imag} */,
  {32'hbf1b69d0, 32'h00000000} /* (18, 23, 5) {real, imag} */,
  {32'hbf6e743d, 32'h00000000} /* (18, 23, 4) {real, imag} */,
  {32'hbf8ecc34, 32'h00000000} /* (18, 23, 3) {real, imag} */,
  {32'hbfa99e50, 32'h00000000} /* (18, 23, 2) {real, imag} */,
  {32'hbf5ad2e9, 32'h00000000} /* (18, 23, 1) {real, imag} */,
  {32'hbe6d8c2f, 32'h00000000} /* (18, 23, 0) {real, imag} */,
  {32'hbee5d132, 32'h00000000} /* (18, 22, 31) {real, imag} */,
  {32'hbf2bbde1, 32'h00000000} /* (18, 22, 30) {real, imag} */,
  {32'hbf597a83, 32'h00000000} /* (18, 22, 29) {real, imag} */,
  {32'hbfc488b6, 32'h00000000} /* (18, 22, 28) {real, imag} */,
  {32'hbfaccbdf, 32'h00000000} /* (18, 22, 27) {real, imag} */,
  {32'hbf2ae5ae, 32'h00000000} /* (18, 22, 26) {real, imag} */,
  {32'hbd2001ae, 32'h00000000} /* (18, 22, 25) {real, imag} */,
  {32'hbf1088a5, 32'h00000000} /* (18, 22, 24) {real, imag} */,
  {32'hbf92efaa, 32'h00000000} /* (18, 22, 23) {real, imag} */,
  {32'hbf84bb18, 32'h00000000} /* (18, 22, 22) {real, imag} */,
  {32'hbee50685, 32'h00000000} /* (18, 22, 21) {real, imag} */,
  {32'h3eb4e5ef, 32'h00000000} /* (18, 22, 20) {real, imag} */,
  {32'h3f2394eb, 32'h00000000} /* (18, 22, 19) {real, imag} */,
  {32'h3f6f1cd3, 32'h00000000} /* (18, 22, 18) {real, imag} */,
  {32'h3fc9401b, 32'h00000000} /* (18, 22, 17) {real, imag} */,
  {32'h3fbdb2f7, 32'h00000000} /* (18, 22, 16) {real, imag} */,
  {32'h3f7874d0, 32'h00000000} /* (18, 22, 15) {real, imag} */,
  {32'h3f3a0afa, 32'h00000000} /* (18, 22, 14) {real, imag} */,
  {32'h3f131a49, 32'h00000000} /* (18, 22, 13) {real, imag} */,
  {32'h3f27d198, 32'h00000000} /* (18, 22, 12) {real, imag} */,
  {32'h3e0aa592, 32'h00000000} /* (18, 22, 11) {real, imag} */,
  {32'hbf1ee09e, 32'h00000000} /* (18, 22, 10) {real, imag} */,
  {32'hbf50efb9, 32'h00000000} /* (18, 22, 9) {real, imag} */,
  {32'hbf767f77, 32'h00000000} /* (18, 22, 8) {real, imag} */,
  {32'hbf77c00f, 32'h00000000} /* (18, 22, 7) {real, imag} */,
  {32'hbf2bd950, 32'h00000000} /* (18, 22, 6) {real, imag} */,
  {32'hbf255d1f, 32'h00000000} /* (18, 22, 5) {real, imag} */,
  {32'hbf29566e, 32'h00000000} /* (18, 22, 4) {real, imag} */,
  {32'hbf144ac1, 32'h00000000} /* (18, 22, 3) {real, imag} */,
  {32'hbf6c9587, 32'h00000000} /* (18, 22, 2) {real, imag} */,
  {32'hbf95746e, 32'h00000000} /* (18, 22, 1) {real, imag} */,
  {32'hbf35101e, 32'h00000000} /* (18, 22, 0) {real, imag} */,
  {32'hbf162785, 32'h00000000} /* (18, 21, 31) {real, imag} */,
  {32'hbf9901d7, 32'h00000000} /* (18, 21, 30) {real, imag} */,
  {32'hbf53741b, 32'h00000000} /* (18, 21, 29) {real, imag} */,
  {32'hbf198507, 32'h00000000} /* (18, 21, 28) {real, imag} */,
  {32'hbf87e74c, 32'h00000000} /* (18, 21, 27) {real, imag} */,
  {32'hbf709c7e, 32'h00000000} /* (18, 21, 26) {real, imag} */,
  {32'hbeb086e7, 32'h00000000} /* (18, 21, 25) {real, imag} */,
  {32'hbe80084a, 32'h00000000} /* (18, 21, 24) {real, imag} */,
  {32'hbed06736, 32'h00000000} /* (18, 21, 23) {real, imag} */,
  {32'hbf00de31, 32'h00000000} /* (18, 21, 22) {real, imag} */,
  {32'hbf246ccc, 32'h00000000} /* (18, 21, 21) {real, imag} */,
  {32'hbbaa295c, 32'h00000000} /* (18, 21, 20) {real, imag} */,
  {32'h3f377cdd, 32'h00000000} /* (18, 21, 19) {real, imag} */,
  {32'h3f0c992c, 32'h00000000} /* (18, 21, 18) {real, imag} */,
  {32'h3f07799c, 32'h00000000} /* (18, 21, 17) {real, imag} */,
  {32'h3ebfea76, 32'h00000000} /* (18, 21, 16) {real, imag} */,
  {32'h3e9e9f63, 32'h00000000} /* (18, 21, 15) {real, imag} */,
  {32'h3e27b85a, 32'h00000000} /* (18, 21, 14) {real, imag} */,
  {32'h3e6f7a00, 32'h00000000} /* (18, 21, 13) {real, imag} */,
  {32'h3e522b9a, 32'h00000000} /* (18, 21, 12) {real, imag} */,
  {32'h3dd2fdc3, 32'h00000000} /* (18, 21, 11) {real, imag} */,
  {32'hbe4008ce, 32'h00000000} /* (18, 21, 10) {real, imag} */,
  {32'hbedea784, 32'h00000000} /* (18, 21, 9) {real, imag} */,
  {32'hbea9e890, 32'h00000000} /* (18, 21, 8) {real, imag} */,
  {32'hbec1d258, 32'h00000000} /* (18, 21, 7) {real, imag} */,
  {32'hbe160572, 32'h00000000} /* (18, 21, 6) {real, imag} */,
  {32'hbcd3cb4a, 32'h00000000} /* (18, 21, 5) {real, imag} */,
  {32'hbe2b7c4d, 32'h00000000} /* (18, 21, 4) {real, imag} */,
  {32'h3c7b3171, 32'h00000000} /* (18, 21, 3) {real, imag} */,
  {32'hbeb4e820, 32'h00000000} /* (18, 21, 2) {real, imag} */,
  {32'hbf3a95c2, 32'h00000000} /* (18, 21, 1) {real, imag} */,
  {32'hbe98156a, 32'h00000000} /* (18, 21, 0) {real, imag} */,
  {32'h3e4b94ba, 32'h00000000} /* (18, 20, 31) {real, imag} */,
  {32'hbcc71304, 32'h00000000} /* (18, 20, 30) {real, imag} */,
  {32'hbe5c975e, 32'h00000000} /* (18, 20, 29) {real, imag} */,
  {32'h3edc69f2, 32'h00000000} /* (18, 20, 28) {real, imag} */,
  {32'h3eb726f1, 32'h00000000} /* (18, 20, 27) {real, imag} */,
  {32'hbb1e4680, 32'h00000000} /* (18, 20, 26) {real, imag} */,
  {32'h3dc2d9f1, 32'h00000000} /* (18, 20, 25) {real, imag} */,
  {32'h3f2c4571, 32'h00000000} /* (18, 20, 24) {real, imag} */,
  {32'h3f6a2bdf, 32'h00000000} /* (18, 20, 23) {real, imag} */,
  {32'h3ef89f6f, 32'h00000000} /* (18, 20, 22) {real, imag} */,
  {32'hbeb4ab0c, 32'h00000000} /* (18, 20, 21) {real, imag} */,
  {32'hbf3163db, 32'h00000000} /* (18, 20, 20) {real, imag} */,
  {32'h3d9bb09c, 32'h00000000} /* (18, 20, 19) {real, imag} */,
  {32'hbdd064dd, 32'h00000000} /* (18, 20, 18) {real, imag} */,
  {32'hbea769f6, 32'h00000000} /* (18, 20, 17) {real, imag} */,
  {32'hbf1a76ed, 32'h00000000} /* (18, 20, 16) {real, imag} */,
  {32'hbf0eb522, 32'h00000000} /* (18, 20, 15) {real, imag} */,
  {32'hbf50bd4c, 32'h00000000} /* (18, 20, 14) {real, imag} */,
  {32'hbf57de30, 32'h00000000} /* (18, 20, 13) {real, imag} */,
  {32'hbf830726, 32'h00000000} /* (18, 20, 12) {real, imag} */,
  {32'hbf7ef387, 32'h00000000} /* (18, 20, 11) {real, imag} */,
  {32'h3e24d3d7, 32'h00000000} /* (18, 20, 10) {real, imag} */,
  {32'h3f3651b1, 32'h00000000} /* (18, 20, 9) {real, imag} */,
  {32'h3fa56bb8, 32'h00000000} /* (18, 20, 8) {real, imag} */,
  {32'h3f86ad48, 32'h00000000} /* (18, 20, 7) {real, imag} */,
  {32'h3ee425e3, 32'h00000000} /* (18, 20, 6) {real, imag} */,
  {32'h3f01cd0b, 32'h00000000} /* (18, 20, 5) {real, imag} */,
  {32'h3f22a710, 32'h00000000} /* (18, 20, 4) {real, imag} */,
  {32'h3f55551b, 32'h00000000} /* (18, 20, 3) {real, imag} */,
  {32'h3f675694, 32'h00000000} /* (18, 20, 2) {real, imag} */,
  {32'h3f09ef00, 32'h00000000} /* (18, 20, 1) {real, imag} */,
  {32'h3edc95c3, 32'h00000000} /* (18, 20, 0) {real, imag} */,
  {32'h3ed2ce4f, 32'h00000000} /* (18, 19, 31) {real, imag} */,
  {32'h3f44a68c, 32'h00000000} /* (18, 19, 30) {real, imag} */,
  {32'h3f0ffd05, 32'h00000000} /* (18, 19, 29) {real, imag} */,
  {32'h3f562c51, 32'h00000000} /* (18, 19, 28) {real, imag} */,
  {32'h3f2f02a7, 32'h00000000} /* (18, 19, 27) {real, imag} */,
  {32'h3ee6eb3c, 32'h00000000} /* (18, 19, 26) {real, imag} */,
  {32'h3f58c6d9, 32'h00000000} /* (18, 19, 25) {real, imag} */,
  {32'h3fc33df1, 32'h00000000} /* (18, 19, 24) {real, imag} */,
  {32'h3f88839f, 32'h00000000} /* (18, 19, 23) {real, imag} */,
  {32'h3f3d44fd, 32'h00000000} /* (18, 19, 22) {real, imag} */,
  {32'h3a7d1f00, 32'h00000000} /* (18, 19, 21) {real, imag} */,
  {32'hbf9dabd7, 32'h00000000} /* (18, 19, 20) {real, imag} */,
  {32'hbf48e9c4, 32'h00000000} /* (18, 19, 19) {real, imag} */,
  {32'hbf02fdcb, 32'h00000000} /* (18, 19, 18) {real, imag} */,
  {32'hbf3bc737, 32'h00000000} /* (18, 19, 17) {real, imag} */,
  {32'hbf1a8ac9, 32'h00000000} /* (18, 19, 16) {real, imag} */,
  {32'hbf3f3bbc, 32'h00000000} /* (18, 19, 15) {real, imag} */,
  {32'hbf376748, 32'h00000000} /* (18, 19, 14) {real, imag} */,
  {32'hbf387df4, 32'h00000000} /* (18, 19, 13) {real, imag} */,
  {32'hbf78ee52, 32'h00000000} /* (18, 19, 12) {real, imag} */,
  {32'hbf9d0747, 32'h00000000} /* (18, 19, 11) {real, imag} */,
  {32'hbe9f7f6f, 32'h00000000} /* (18, 19, 10) {real, imag} */,
  {32'h3f88f656, 32'h00000000} /* (18, 19, 9) {real, imag} */,
  {32'h3fdedf39, 32'h00000000} /* (18, 19, 8) {real, imag} */,
  {32'h3fc781b3, 32'h00000000} /* (18, 19, 7) {real, imag} */,
  {32'h3f28d1a7, 32'h00000000} /* (18, 19, 6) {real, imag} */,
  {32'h3f149c59, 32'h00000000} /* (18, 19, 5) {real, imag} */,
  {32'h3f738530, 32'h00000000} /* (18, 19, 4) {real, imag} */,
  {32'h3f40bafb, 32'h00000000} /* (18, 19, 3) {real, imag} */,
  {32'h3fa911c3, 32'h00000000} /* (18, 19, 2) {real, imag} */,
  {32'h3fae0d55, 32'h00000000} /* (18, 19, 1) {real, imag} */,
  {32'h3f18e021, 32'h00000000} /* (18, 19, 0) {real, imag} */,
  {32'h3f7d9f2f, 32'h00000000} /* (18, 18, 31) {real, imag} */,
  {32'h3fd010a6, 32'h00000000} /* (18, 18, 30) {real, imag} */,
  {32'h3f8296fd, 32'h00000000} /* (18, 18, 29) {real, imag} */,
  {32'h3f49bff5, 32'h00000000} /* (18, 18, 28) {real, imag} */,
  {32'h3f14619e, 32'h00000000} /* (18, 18, 27) {real, imag} */,
  {32'h3edc14ac, 32'h00000000} /* (18, 18, 26) {real, imag} */,
  {32'h3f8604a9, 32'h00000000} /* (18, 18, 25) {real, imag} */,
  {32'h3f99c98c, 32'h00000000} /* (18, 18, 24) {real, imag} */,
  {32'h3f66f679, 32'h00000000} /* (18, 18, 23) {real, imag} */,
  {32'h3f134e7d, 32'h00000000} /* (18, 18, 22) {real, imag} */,
  {32'h3d363aa6, 32'h00000000} /* (18, 18, 21) {real, imag} */,
  {32'hbf638c6e, 32'h00000000} /* (18, 18, 20) {real, imag} */,
  {32'hbf70cfb5, 32'h00000000} /* (18, 18, 19) {real, imag} */,
  {32'hbf54b88a, 32'h00000000} /* (18, 18, 18) {real, imag} */,
  {32'hbf70e58b, 32'h00000000} /* (18, 18, 17) {real, imag} */,
  {32'hbf3b0122, 32'h00000000} /* (18, 18, 16) {real, imag} */,
  {32'hbf430079, 32'h00000000} /* (18, 18, 15) {real, imag} */,
  {32'hbf459936, 32'h00000000} /* (18, 18, 14) {real, imag} */,
  {32'hbf7e91de, 32'h00000000} /* (18, 18, 13) {real, imag} */,
  {32'hbfa82c90, 32'h00000000} /* (18, 18, 12) {real, imag} */,
  {32'hbf90d82d, 32'h00000000} /* (18, 18, 11) {real, imag} */,
  {32'h3d3b8074, 32'h00000000} /* (18, 18, 10) {real, imag} */,
  {32'h3fb50405, 32'h00000000} /* (18, 18, 9) {real, imag} */,
  {32'h3fc802de, 32'h00000000} /* (18, 18, 8) {real, imag} */,
  {32'h3fa56dfc, 32'h00000000} /* (18, 18, 7) {real, imag} */,
  {32'h3f20c933, 32'h00000000} /* (18, 18, 6) {real, imag} */,
  {32'h3ebcb4c4, 32'h00000000} /* (18, 18, 5) {real, imag} */,
  {32'h3f31ba4b, 32'h00000000} /* (18, 18, 4) {real, imag} */,
  {32'h3edf7511, 32'h00000000} /* (18, 18, 3) {real, imag} */,
  {32'h3f3dcd52, 32'h00000000} /* (18, 18, 2) {real, imag} */,
  {32'h3f93ec66, 32'h00000000} /* (18, 18, 1) {real, imag} */,
  {32'h3f59fc8b, 32'h00000000} /* (18, 18, 0) {real, imag} */,
  {32'h3f5e43fc, 32'h00000000} /* (18, 17, 31) {real, imag} */,
  {32'h3fb3f266, 32'h00000000} /* (18, 17, 30) {real, imag} */,
  {32'h3f913edd, 32'h00000000} /* (18, 17, 29) {real, imag} */,
  {32'h3f797c5c, 32'h00000000} /* (18, 17, 28) {real, imag} */,
  {32'h3f81d8f5, 32'h00000000} /* (18, 17, 27) {real, imag} */,
  {32'h3f0764ce, 32'h00000000} /* (18, 17, 26) {real, imag} */,
  {32'h3f052f42, 32'h00000000} /* (18, 17, 25) {real, imag} */,
  {32'h3f469c79, 32'h00000000} /* (18, 17, 24) {real, imag} */,
  {32'h3f941da8, 32'h00000000} /* (18, 17, 23) {real, imag} */,
  {32'h3f2eed6a, 32'h00000000} /* (18, 17, 22) {real, imag} */,
  {32'h3d5c26b8, 32'h00000000} /* (18, 17, 21) {real, imag} */,
  {32'hbf798eb6, 32'h00000000} /* (18, 17, 20) {real, imag} */,
  {32'hbf7d1ee0, 32'h00000000} /* (18, 17, 19) {real, imag} */,
  {32'hbf1aa7a4, 32'h00000000} /* (18, 17, 18) {real, imag} */,
  {32'hbf4d9895, 32'h00000000} /* (18, 17, 17) {real, imag} */,
  {32'hbf638ec2, 32'h00000000} /* (18, 17, 16) {real, imag} */,
  {32'hbf5060c0, 32'h00000000} /* (18, 17, 15) {real, imag} */,
  {32'hbf3c1210, 32'h00000000} /* (18, 17, 14) {real, imag} */,
  {32'hbf59cf86, 32'h00000000} /* (18, 17, 13) {real, imag} */,
  {32'hbfcca2c8, 32'h00000000} /* (18, 17, 12) {real, imag} */,
  {32'hbf60af7c, 32'h00000000} /* (18, 17, 11) {real, imag} */,
  {32'h3f46c290, 32'h00000000} /* (18, 17, 10) {real, imag} */,
  {32'h3fb3d9b1, 32'h00000000} /* (18, 17, 9) {real, imag} */,
  {32'h3fa2b360, 32'h00000000} /* (18, 17, 8) {real, imag} */,
  {32'h3f5fbae9, 32'h00000000} /* (18, 17, 7) {real, imag} */,
  {32'h3f31f8f3, 32'h00000000} /* (18, 17, 6) {real, imag} */,
  {32'h3ee78d60, 32'h00000000} /* (18, 17, 5) {real, imag} */,
  {32'h3f1b0a90, 32'h00000000} /* (18, 17, 4) {real, imag} */,
  {32'h3f3047b1, 32'h00000000} /* (18, 17, 3) {real, imag} */,
  {32'h3f647eba, 32'h00000000} /* (18, 17, 2) {real, imag} */,
  {32'h3f4dad3b, 32'h00000000} /* (18, 17, 1) {real, imag} */,
  {32'h3f5baa3e, 32'h00000000} /* (18, 17, 0) {real, imag} */,
  {32'h3ee8a131, 32'h00000000} /* (18, 16, 31) {real, imag} */,
  {32'h3f9cd2ef, 32'h00000000} /* (18, 16, 30) {real, imag} */,
  {32'h3fbd3907, 32'h00000000} /* (18, 16, 29) {real, imag} */,
  {32'h3f8a4655, 32'h00000000} /* (18, 16, 28) {real, imag} */,
  {32'h3fc301cd, 32'h00000000} /* (18, 16, 27) {real, imag} */,
  {32'h3fa17197, 32'h00000000} /* (18, 16, 26) {real, imag} */,
  {32'h3f5d8b8b, 32'h00000000} /* (18, 16, 25) {real, imag} */,
  {32'h3faad503, 32'h00000000} /* (18, 16, 24) {real, imag} */,
  {32'h3fa1f269, 32'h00000000} /* (18, 16, 23) {real, imag} */,
  {32'h3f493ebf, 32'h00000000} /* (18, 16, 22) {real, imag} */,
  {32'h3eada49f, 32'h00000000} /* (18, 16, 21) {real, imag} */,
  {32'hbfaaae8d, 32'h00000000} /* (18, 16, 20) {real, imag} */,
  {32'hbfb41891, 32'h00000000} /* (18, 16, 19) {real, imag} */,
  {32'hbf7fefc9, 32'h00000000} /* (18, 16, 18) {real, imag} */,
  {32'hbf756581, 32'h00000000} /* (18, 16, 17) {real, imag} */,
  {32'hbf8238b8, 32'h00000000} /* (18, 16, 16) {real, imag} */,
  {32'hbf985be1, 32'h00000000} /* (18, 16, 15) {real, imag} */,
  {32'hbf82c048, 32'h00000000} /* (18, 16, 14) {real, imag} */,
  {32'hbf909711, 32'h00000000} /* (18, 16, 13) {real, imag} */,
  {32'hbfb260f7, 32'h00000000} /* (18, 16, 12) {real, imag} */,
  {32'hbef86cf5, 32'h00000000} /* (18, 16, 11) {real, imag} */,
  {32'h3f7588a2, 32'h00000000} /* (18, 16, 10) {real, imag} */,
  {32'h3fce9969, 32'h00000000} /* (18, 16, 9) {real, imag} */,
  {32'h3fca1dd9, 32'h00000000} /* (18, 16, 8) {real, imag} */,
  {32'h3f8829be, 32'h00000000} /* (18, 16, 7) {real, imag} */,
  {32'h3f0adaba, 32'h00000000} /* (18, 16, 6) {real, imag} */,
  {32'h3eeaaf03, 32'h00000000} /* (18, 16, 5) {real, imag} */,
  {32'h3f084eb7, 32'h00000000} /* (18, 16, 4) {real, imag} */,
  {32'h3f400934, 32'h00000000} /* (18, 16, 3) {real, imag} */,
  {32'h3f4da0b6, 32'h00000000} /* (18, 16, 2) {real, imag} */,
  {32'h3f8fbe31, 32'h00000000} /* (18, 16, 1) {real, imag} */,
  {32'h3f030dd4, 32'h00000000} /* (18, 16, 0) {real, imag} */,
  {32'h3e9ba400, 32'h00000000} /* (18, 15, 31) {real, imag} */,
  {32'h3f56dc2f, 32'h00000000} /* (18, 15, 30) {real, imag} */,
  {32'h3f8b5fd8, 32'h00000000} /* (18, 15, 29) {real, imag} */,
  {32'h3f6117f9, 32'h00000000} /* (18, 15, 28) {real, imag} */,
  {32'h3fac2ecd, 32'h00000000} /* (18, 15, 27) {real, imag} */,
  {32'h3fc0af1f, 32'h00000000} /* (18, 15, 26) {real, imag} */,
  {32'h3f5f21fc, 32'h00000000} /* (18, 15, 25) {real, imag} */,
  {32'h3f9e5d40, 32'h00000000} /* (18, 15, 24) {real, imag} */,
  {32'h3f7f3a9d, 32'h00000000} /* (18, 15, 23) {real, imag} */,
  {32'h3fa1ffff, 32'h00000000} /* (18, 15, 22) {real, imag} */,
  {32'h3f8d8c65, 32'h00000000} /* (18, 15, 21) {real, imag} */,
  {32'hbe47f2cc, 32'h00000000} /* (18, 15, 20) {real, imag} */,
  {32'hbf74f7c5, 32'h00000000} /* (18, 15, 19) {real, imag} */,
  {32'hbfa3e7de, 32'h00000000} /* (18, 15, 18) {real, imag} */,
  {32'hbfa6b8a7, 32'h00000000} /* (18, 15, 17) {real, imag} */,
  {32'hbf8d7e46, 32'h00000000} /* (18, 15, 16) {real, imag} */,
  {32'hbf9d7537, 32'h00000000} /* (18, 15, 15) {real, imag} */,
  {32'hbfb460fc, 32'h00000000} /* (18, 15, 14) {real, imag} */,
  {32'hbfa5797e, 32'h00000000} /* (18, 15, 13) {real, imag} */,
  {32'hbfab0ddb, 32'h00000000} /* (18, 15, 12) {real, imag} */,
  {32'hbf8f2fc2, 32'h00000000} /* (18, 15, 11) {real, imag} */,
  {32'h3f0dedf7, 32'h00000000} /* (18, 15, 10) {real, imag} */,
  {32'h3f9e773c, 32'h00000000} /* (18, 15, 9) {real, imag} */,
  {32'h3fb666f3, 32'h00000000} /* (18, 15, 8) {real, imag} */,
  {32'h3fbdbbea, 32'h00000000} /* (18, 15, 7) {real, imag} */,
  {32'h3f347a26, 32'h00000000} /* (18, 15, 6) {real, imag} */,
  {32'h3efaffd9, 32'h00000000} /* (18, 15, 5) {real, imag} */,
  {32'h3f7f2037, 32'h00000000} /* (18, 15, 4) {real, imag} */,
  {32'h3f8148e1, 32'h00000000} /* (18, 15, 3) {real, imag} */,
  {32'h3f395af5, 32'h00000000} /* (18, 15, 2) {real, imag} */,
  {32'h3fb71d96, 32'h00000000} /* (18, 15, 1) {real, imag} */,
  {32'h3f5feb24, 32'h00000000} /* (18, 15, 0) {real, imag} */,
  {32'h3ebddd1d, 32'h00000000} /* (18, 14, 31) {real, imag} */,
  {32'h3f149f55, 32'h00000000} /* (18, 14, 30) {real, imag} */,
  {32'h3f6af906, 32'h00000000} /* (18, 14, 29) {real, imag} */,
  {32'h3f663014, 32'h00000000} /* (18, 14, 28) {real, imag} */,
  {32'h3f359b19, 32'h00000000} /* (18, 14, 27) {real, imag} */,
  {32'h3f7b076f, 32'h00000000} /* (18, 14, 26) {real, imag} */,
  {32'h3f2ad6de, 32'h00000000} /* (18, 14, 25) {real, imag} */,
  {32'h3f2ee470, 32'h00000000} /* (18, 14, 24) {real, imag} */,
  {32'h3f4950b2, 32'h00000000} /* (18, 14, 23) {real, imag} */,
  {32'h3fe18fc6, 32'h00000000} /* (18, 14, 22) {real, imag} */,
  {32'h3fa4caef, 32'h00000000} /* (18, 14, 21) {real, imag} */,
  {32'hbe8b14c5, 32'h00000000} /* (18, 14, 20) {real, imag} */,
  {32'hbf8a0124, 32'h00000000} /* (18, 14, 19) {real, imag} */,
  {32'hbf9b15b3, 32'h00000000} /* (18, 14, 18) {real, imag} */,
  {32'hbf818f66, 32'h00000000} /* (18, 14, 17) {real, imag} */,
  {32'hbf6d8f33, 32'h00000000} /* (18, 14, 16) {real, imag} */,
  {32'hbf9221b6, 32'h00000000} /* (18, 14, 15) {real, imag} */,
  {32'hbfedc140, 32'h00000000} /* (18, 14, 14) {real, imag} */,
  {32'hbf9f17f2, 32'h00000000} /* (18, 14, 13) {real, imag} */,
  {32'hbf448578, 32'h00000000} /* (18, 14, 12) {real, imag} */,
  {32'hbf151332, 32'h00000000} /* (18, 14, 11) {real, imag} */,
  {32'h3eea5fa0, 32'h00000000} /* (18, 14, 10) {real, imag} */,
  {32'h3f8bef1a, 32'h00000000} /* (18, 14, 9) {real, imag} */,
  {32'h3f8c67e5, 32'h00000000} /* (18, 14, 8) {real, imag} */,
  {32'h3f75b2ba, 32'h00000000} /* (18, 14, 7) {real, imag} */,
  {32'h3f32cc29, 32'h00000000} /* (18, 14, 6) {real, imag} */,
  {32'h3ec407e8, 32'h00000000} /* (18, 14, 5) {real, imag} */,
  {32'h3f138239, 32'h00000000} /* (18, 14, 4) {real, imag} */,
  {32'h3f560262, 32'h00000000} /* (18, 14, 3) {real, imag} */,
  {32'h3f99a993, 32'h00000000} /* (18, 14, 2) {real, imag} */,
  {32'h3fb1af91, 32'h00000000} /* (18, 14, 1) {real, imag} */,
  {32'h3f4a2254, 32'h00000000} /* (18, 14, 0) {real, imag} */,
  {32'h3eb36f84, 32'h00000000} /* (18, 13, 31) {real, imag} */,
  {32'h3f47cf24, 32'h00000000} /* (18, 13, 30) {real, imag} */,
  {32'h3f648393, 32'h00000000} /* (18, 13, 29) {real, imag} */,
  {32'h3f86b5a7, 32'h00000000} /* (18, 13, 28) {real, imag} */,
  {32'h3f064ed0, 32'h00000000} /* (18, 13, 27) {real, imag} */,
  {32'h3f248a53, 32'h00000000} /* (18, 13, 26) {real, imag} */,
  {32'h3f2beb9c, 32'h00000000} /* (18, 13, 25) {real, imag} */,
  {32'h3ee39181, 32'h00000000} /* (18, 13, 24) {real, imag} */,
  {32'h3f0bda69, 32'h00000000} /* (18, 13, 23) {real, imag} */,
  {32'h3f73d622, 32'h00000000} /* (18, 13, 22) {real, imag} */,
  {32'h3f2ffd56, 32'h00000000} /* (18, 13, 21) {real, imag} */,
  {32'hbf13e926, 32'h00000000} /* (18, 13, 20) {real, imag} */,
  {32'hbf8030e1, 32'h00000000} /* (18, 13, 19) {real, imag} */,
  {32'hbf0d4495, 32'h00000000} /* (18, 13, 18) {real, imag} */,
  {32'hbf8ecb88, 32'h00000000} /* (18, 13, 17) {real, imag} */,
  {32'hbfa060d2, 32'h00000000} /* (18, 13, 16) {real, imag} */,
  {32'hbf8def26, 32'h00000000} /* (18, 13, 15) {real, imag} */,
  {32'hbfd5e2f8, 32'h00000000} /* (18, 13, 14) {real, imag} */,
  {32'hbf892a04, 32'h00000000} /* (18, 13, 13) {real, imag} */,
  {32'hbec74983, 32'h00000000} /* (18, 13, 12) {real, imag} */,
  {32'h3cf58432, 32'h00000000} /* (18, 13, 11) {real, imag} */,
  {32'h3f21d883, 32'h00000000} /* (18, 13, 10) {real, imag} */,
  {32'h3f4c150b, 32'h00000000} /* (18, 13, 9) {real, imag} */,
  {32'h3f8b52d8, 32'h00000000} /* (18, 13, 8) {real, imag} */,
  {32'h3f86839a, 32'h00000000} /* (18, 13, 7) {real, imag} */,
  {32'h3f513fe9, 32'h00000000} /* (18, 13, 6) {real, imag} */,
  {32'h3f54afe2, 32'h00000000} /* (18, 13, 5) {real, imag} */,
  {32'h3f035d6d, 32'h00000000} /* (18, 13, 4) {real, imag} */,
  {32'h3f88fe7c, 32'h00000000} /* (18, 13, 3) {real, imag} */,
  {32'h3f83af17, 32'h00000000} /* (18, 13, 2) {real, imag} */,
  {32'h3f81058c, 32'h00000000} /* (18, 13, 1) {real, imag} */,
  {32'h3f332205, 32'h00000000} /* (18, 13, 0) {real, imag} */,
  {32'h3eeb2c91, 32'h00000000} /* (18, 12, 31) {real, imag} */,
  {32'h3f37eaee, 32'h00000000} /* (18, 12, 30) {real, imag} */,
  {32'h3f27e78e, 32'h00000000} /* (18, 12, 29) {real, imag} */,
  {32'h3f51aba3, 32'h00000000} /* (18, 12, 28) {real, imag} */,
  {32'h3f3cfe4b, 32'h00000000} /* (18, 12, 27) {real, imag} */,
  {32'h3f443ce0, 32'h00000000} /* (18, 12, 26) {real, imag} */,
  {32'h3f23528f, 32'h00000000} /* (18, 12, 25) {real, imag} */,
  {32'h3e95ede6, 32'h00000000} /* (18, 12, 24) {real, imag} */,
  {32'h3f510256, 32'h00000000} /* (18, 12, 23) {real, imag} */,
  {32'h3f8cb213, 32'h00000000} /* (18, 12, 22) {real, imag} */,
  {32'h3f39353c, 32'h00000000} /* (18, 12, 21) {real, imag} */,
  {32'hbedee55a, 32'h00000000} /* (18, 12, 20) {real, imag} */,
  {32'hbf93dbe5, 32'h00000000} /* (18, 12, 19) {real, imag} */,
  {32'hbf15ee56, 32'h00000000} /* (18, 12, 18) {real, imag} */,
  {32'hbf967d38, 32'h00000000} /* (18, 12, 17) {real, imag} */,
  {32'hbfba9925, 32'h00000000} /* (18, 12, 16) {real, imag} */,
  {32'hbfa513a5, 32'h00000000} /* (18, 12, 15) {real, imag} */,
  {32'hbfbc7f72, 32'h00000000} /* (18, 12, 14) {real, imag} */,
  {32'hbf998b26, 32'h00000000} /* (18, 12, 13) {real, imag} */,
  {32'hbf5e10dc, 32'h00000000} /* (18, 12, 12) {real, imag} */,
  {32'hbf2a8702, 32'h00000000} /* (18, 12, 11) {real, imag} */,
  {32'h3ec7dd3c, 32'h00000000} /* (18, 12, 10) {real, imag} */,
  {32'h3f362a5c, 32'h00000000} /* (18, 12, 9) {real, imag} */,
  {32'h3f853b93, 32'h00000000} /* (18, 12, 8) {real, imag} */,
  {32'h3fbbac2c, 32'h00000000} /* (18, 12, 7) {real, imag} */,
  {32'h3f91b16d, 32'h00000000} /* (18, 12, 6) {real, imag} */,
  {32'h3f80fc91, 32'h00000000} /* (18, 12, 5) {real, imag} */,
  {32'h3f31ac3b, 32'h00000000} /* (18, 12, 4) {real, imag} */,
  {32'h3f89b054, 32'h00000000} /* (18, 12, 3) {real, imag} */,
  {32'h3f153217, 32'h00000000} /* (18, 12, 2) {real, imag} */,
  {32'h3f4b1d8e, 32'h00000000} /* (18, 12, 1) {real, imag} */,
  {32'h3f2cfb44, 32'h00000000} /* (18, 12, 0) {real, imag} */,
  {32'h3e9a28a3, 32'h00000000} /* (18, 11, 31) {real, imag} */,
  {32'h3f1cffd5, 32'h00000000} /* (18, 11, 30) {real, imag} */,
  {32'h3ed2bfd4, 32'h00000000} /* (18, 11, 29) {real, imag} */,
  {32'h3f199677, 32'h00000000} /* (18, 11, 28) {real, imag} */,
  {32'h3e118266, 32'h00000000} /* (18, 11, 27) {real, imag} */,
  {32'h3e82dacf, 32'h00000000} /* (18, 11, 26) {real, imag} */,
  {32'h3f19f78a, 32'h00000000} /* (18, 11, 25) {real, imag} */,
  {32'h3eb3349d, 32'h00000000} /* (18, 11, 24) {real, imag} */,
  {32'h3f3ea2d7, 32'h00000000} /* (18, 11, 23) {real, imag} */,
  {32'h3f87a501, 32'h00000000} /* (18, 11, 22) {real, imag} */,
  {32'h3f25ef65, 32'h00000000} /* (18, 11, 21) {real, imag} */,
  {32'hbf0685eb, 32'h00000000} /* (18, 11, 20) {real, imag} */,
  {32'hbf5c3091, 32'h00000000} /* (18, 11, 19) {real, imag} */,
  {32'hbf1f1cde, 32'h00000000} /* (18, 11, 18) {real, imag} */,
  {32'hbf5af733, 32'h00000000} /* (18, 11, 17) {real, imag} */,
  {32'hbf57d9f0, 32'h00000000} /* (18, 11, 16) {real, imag} */,
  {32'hbf45c41f, 32'h00000000} /* (18, 11, 15) {real, imag} */,
  {32'hbfac494d, 32'h00000000} /* (18, 11, 14) {real, imag} */,
  {32'hbf647622, 32'h00000000} /* (18, 11, 13) {real, imag} */,
  {32'hbea578d4, 32'h00000000} /* (18, 11, 12) {real, imag} */,
  {32'hbe548b91, 32'h00000000} /* (18, 11, 11) {real, imag} */,
  {32'h3ee03cdc, 32'h00000000} /* (18, 11, 10) {real, imag} */,
  {32'h3eedbd86, 32'h00000000} /* (18, 11, 9) {real, imag} */,
  {32'h3f0a22e8, 32'h00000000} /* (18, 11, 8) {real, imag} */,
  {32'h3f5fe2f0, 32'h00000000} /* (18, 11, 7) {real, imag} */,
  {32'h3f7d3394, 32'h00000000} /* (18, 11, 6) {real, imag} */,
  {32'h3f67e4d0, 32'h00000000} /* (18, 11, 5) {real, imag} */,
  {32'h3f09f619, 32'h00000000} /* (18, 11, 4) {real, imag} */,
  {32'h3f12d937, 32'h00000000} /* (18, 11, 3) {real, imag} */,
  {32'h3f8255b5, 32'h00000000} /* (18, 11, 2) {real, imag} */,
  {32'h3f817478, 32'h00000000} /* (18, 11, 1) {real, imag} */,
  {32'h3eab1cf2, 32'h00000000} /* (18, 11, 0) {real, imag} */,
  {32'hbea5c8ca, 32'h00000000} /* (18, 10, 31) {real, imag} */,
  {32'hbf028a34, 32'h00000000} /* (18, 10, 30) {real, imag} */,
  {32'hbf0e524c, 32'h00000000} /* (18, 10, 29) {real, imag} */,
  {32'hbf1306dd, 32'h00000000} /* (18, 10, 28) {real, imag} */,
  {32'hbf807e4f, 32'h00000000} /* (18, 10, 27) {real, imag} */,
  {32'hbf4fdf8b, 32'h00000000} /* (18, 10, 26) {real, imag} */,
  {32'hbf2d1fd8, 32'h00000000} /* (18, 10, 25) {real, imag} */,
  {32'hbf7b8098, 32'h00000000} /* (18, 10, 24) {real, imag} */,
  {32'hbf487218, 32'h00000000} /* (18, 10, 23) {real, imag} */,
  {32'hbed325c6, 32'h00000000} /* (18, 10, 22) {real, imag} */,
  {32'hbe41941f, 32'h00000000} /* (18, 10, 21) {real, imag} */,
  {32'h3c43394e, 32'h00000000} /* (18, 10, 20) {real, imag} */,
  {32'h3d625421, 32'h00000000} /* (18, 10, 19) {real, imag} */,
  {32'h3e47b4f0, 32'h00000000} /* (18, 10, 18) {real, imag} */,
  {32'h3e8c6004, 32'h00000000} /* (18, 10, 17) {real, imag} */,
  {32'h3eca8253, 32'h00000000} /* (18, 10, 16) {real, imag} */,
  {32'h3f30fd8c, 32'h00000000} /* (18, 10, 15) {real, imag} */,
  {32'h3ec9b9ed, 32'h00000000} /* (18, 10, 14) {real, imag} */,
  {32'h3f4d6ca8, 32'h00000000} /* (18, 10, 13) {real, imag} */,
  {32'h3f773f8c, 32'h00000000} /* (18, 10, 12) {real, imag} */,
  {32'h3f3720c7, 32'h00000000} /* (18, 10, 11) {real, imag} */,
  {32'hbed2e86f, 32'h00000000} /* (18, 10, 10) {real, imag} */,
  {32'hbf7a5106, 32'h00000000} /* (18, 10, 9) {real, imag} */,
  {32'hbf263d1d, 32'h00000000} /* (18, 10, 8) {real, imag} */,
  {32'hbf477a7f, 32'h00000000} /* (18, 10, 7) {real, imag} */,
  {32'hbf180295, 32'h00000000} /* (18, 10, 6) {real, imag} */,
  {32'hbf34628b, 32'h00000000} /* (18, 10, 5) {real, imag} */,
  {32'hbf60ef7a, 32'h00000000} /* (18, 10, 4) {real, imag} */,
  {32'hbe4d85c0, 32'h00000000} /* (18, 10, 3) {real, imag} */,
  {32'h3d7b8ba7, 32'h00000000} /* (18, 10, 2) {real, imag} */,
  {32'hbf0ab802, 32'h00000000} /* (18, 10, 1) {real, imag} */,
  {32'hbf2523ff, 32'h00000000} /* (18, 10, 0) {real, imag} */,
  {32'hbeba0639, 32'h00000000} /* (18, 9, 31) {real, imag} */,
  {32'hbf8a97a8, 32'h00000000} /* (18, 9, 30) {real, imag} */,
  {32'hbf8199fa, 32'h00000000} /* (18, 9, 29) {real, imag} */,
  {32'hbfb155c9, 32'h00000000} /* (18, 9, 28) {real, imag} */,
  {32'hbfa3e469, 32'h00000000} /* (18, 9, 27) {real, imag} */,
  {32'hbf98f943, 32'h00000000} /* (18, 9, 26) {real, imag} */,
  {32'hbfa58b42, 32'h00000000} /* (18, 9, 25) {real, imag} */,
  {32'hbfae88d7, 32'h00000000} /* (18, 9, 24) {real, imag} */,
  {32'hbf3bb954, 32'h00000000} /* (18, 9, 23) {real, imag} */,
  {32'hbf4a3858, 32'h00000000} /* (18, 9, 22) {real, imag} */,
  {32'hbedc8852, 32'h00000000} /* (18, 9, 21) {real, imag} */,
  {32'h3ea64109, 32'h00000000} /* (18, 9, 20) {real, imag} */,
  {32'h3ee2febc, 32'h00000000} /* (18, 9, 19) {real, imag} */,
  {32'h3f995569, 32'h00000000} /* (18, 9, 18) {real, imag} */,
  {32'h3fb1c6c5, 32'h00000000} /* (18, 9, 17) {real, imag} */,
  {32'h3fa9f239, 32'h00000000} /* (18, 9, 16) {real, imag} */,
  {32'h3fcd3e73, 32'h00000000} /* (18, 9, 15) {real, imag} */,
  {32'h3fa2bafe, 32'h00000000} /* (18, 9, 14) {real, imag} */,
  {32'h3f6fa7cb, 32'h00000000} /* (18, 9, 13) {real, imag} */,
  {32'h3f5d9e1c, 32'h00000000} /* (18, 9, 12) {real, imag} */,
  {32'h3f3320e7, 32'h00000000} /* (18, 9, 11) {real, imag} */,
  {32'hbf3ab08e, 32'h00000000} /* (18, 9, 10) {real, imag} */,
  {32'hbfd666ed, 32'h00000000} /* (18, 9, 9) {real, imag} */,
  {32'hbf965860, 32'h00000000} /* (18, 9, 8) {real, imag} */,
  {32'hbf85d2d6, 32'h00000000} /* (18, 9, 7) {real, imag} */,
  {32'hbf8b5a60, 32'h00000000} /* (18, 9, 6) {real, imag} */,
  {32'hbfc4721b, 32'h00000000} /* (18, 9, 5) {real, imag} */,
  {32'hbfdbf49f, 32'h00000000} /* (18, 9, 4) {real, imag} */,
  {32'hbf3ee7aa, 32'h00000000} /* (18, 9, 3) {real, imag} */,
  {32'hbf37179a, 32'h00000000} /* (18, 9, 2) {real, imag} */,
  {32'hbfadf851, 32'h00000000} /* (18, 9, 1) {real, imag} */,
  {32'hbf82785f, 32'h00000000} /* (18, 9, 0) {real, imag} */,
  {32'hbf2c08d3, 32'h00000000} /* (18, 8, 31) {real, imag} */,
  {32'hbf9e5d05, 32'h00000000} /* (18, 8, 30) {real, imag} */,
  {32'hbfc3f5f1, 32'h00000000} /* (18, 8, 29) {real, imag} */,
  {32'hbff9e985, 32'h00000000} /* (18, 8, 28) {real, imag} */,
  {32'hbfbc17a6, 32'h00000000} /* (18, 8, 27) {real, imag} */,
  {32'hbf9c1690, 32'h00000000} /* (18, 8, 26) {real, imag} */,
  {32'hbf9053e4, 32'h00000000} /* (18, 8, 25) {real, imag} */,
  {32'hbf0bb26e, 32'h00000000} /* (18, 8, 24) {real, imag} */,
  {32'hbec48816, 32'h00000000} /* (18, 8, 23) {real, imag} */,
  {32'hbf017a26, 32'h00000000} /* (18, 8, 22) {real, imag} */,
  {32'hbe7e14d2, 32'h00000000} /* (18, 8, 21) {real, imag} */,
  {32'h3f079bbd, 32'h00000000} /* (18, 8, 20) {real, imag} */,
  {32'h3ef2a1df, 32'h00000000} /* (18, 8, 19) {real, imag} */,
  {32'h3f7b0a1c, 32'h00000000} /* (18, 8, 18) {real, imag} */,
  {32'h3f6f682a, 32'h00000000} /* (18, 8, 17) {real, imag} */,
  {32'h3f87c43f, 32'h00000000} /* (18, 8, 16) {real, imag} */,
  {32'h3f8e63c2, 32'h00000000} /* (18, 8, 15) {real, imag} */,
  {32'h3f51a2a2, 32'h00000000} /* (18, 8, 14) {real, imag} */,
  {32'h3f16988d, 32'h00000000} /* (18, 8, 13) {real, imag} */,
  {32'h3f5606a9, 32'h00000000} /* (18, 8, 12) {real, imag} */,
  {32'h3f49f4c3, 32'h00000000} /* (18, 8, 11) {real, imag} */,
  {32'hbf1c680d, 32'h00000000} /* (18, 8, 10) {real, imag} */,
  {32'hbfa5b75d, 32'h00000000} /* (18, 8, 9) {real, imag} */,
  {32'hbf638c0a, 32'h00000000} /* (18, 8, 8) {real, imag} */,
  {32'hbf1c93a7, 32'h00000000} /* (18, 8, 7) {real, imag} */,
  {32'hbf8b6273, 32'h00000000} /* (18, 8, 6) {real, imag} */,
  {32'hbfafbb2d, 32'h00000000} /* (18, 8, 5) {real, imag} */,
  {32'hbf9952fc, 32'h00000000} /* (18, 8, 4) {real, imag} */,
  {32'hbf83738a, 32'h00000000} /* (18, 8, 3) {real, imag} */,
  {32'hbf899a4e, 32'h00000000} /* (18, 8, 2) {real, imag} */,
  {32'hbf6cbb65, 32'h00000000} /* (18, 8, 1) {real, imag} */,
  {32'hbf76f9b8, 32'h00000000} /* (18, 8, 0) {real, imag} */,
  {32'hbf57e15b, 32'h00000000} /* (18, 7, 31) {real, imag} */,
  {32'hbf92ddf5, 32'h00000000} /* (18, 7, 30) {real, imag} */,
  {32'hbf963aaf, 32'h00000000} /* (18, 7, 29) {real, imag} */,
  {32'hbf8a3335, 32'h00000000} /* (18, 7, 28) {real, imag} */,
  {32'hbf8a1f7c, 32'h00000000} /* (18, 7, 27) {real, imag} */,
  {32'hbfa8afa6, 32'h00000000} /* (18, 7, 26) {real, imag} */,
  {32'hbff899ed, 32'h00000000} /* (18, 7, 25) {real, imag} */,
  {32'hbf9a7721, 32'h00000000} /* (18, 7, 24) {real, imag} */,
  {32'hbf2fed43, 32'h00000000} /* (18, 7, 23) {real, imag} */,
  {32'hbf2dae61, 32'h00000000} /* (18, 7, 22) {real, imag} */,
  {32'hbf9747f2, 32'h00000000} /* (18, 7, 21) {real, imag} */,
  {32'h3eaccc86, 32'h00000000} /* (18, 7, 20) {real, imag} */,
  {32'h3f6d75df, 32'h00000000} /* (18, 7, 19) {real, imag} */,
  {32'h3fbe725b, 32'h00000000} /* (18, 7, 18) {real, imag} */,
  {32'h3f9d3296, 32'h00000000} /* (18, 7, 17) {real, imag} */,
  {32'h3f6b5929, 32'h00000000} /* (18, 7, 16) {real, imag} */,
  {32'h3f983927, 32'h00000000} /* (18, 7, 15) {real, imag} */,
  {32'h3f1ff803, 32'h00000000} /* (18, 7, 14) {real, imag} */,
  {32'h3efcea96, 32'h00000000} /* (18, 7, 13) {real, imag} */,
  {32'h3f914868, 32'h00000000} /* (18, 7, 12) {real, imag} */,
  {32'h3f96f5e7, 32'h00000000} /* (18, 7, 11) {real, imag} */,
  {32'hbf1a8732, 32'h00000000} /* (18, 7, 10) {real, imag} */,
  {32'hbfa391b9, 32'h00000000} /* (18, 7, 9) {real, imag} */,
  {32'hbf8b20c9, 32'h00000000} /* (18, 7, 8) {real, imag} */,
  {32'hbf3b6429, 32'h00000000} /* (18, 7, 7) {real, imag} */,
  {32'hbfb8ed26, 32'h00000000} /* (18, 7, 6) {real, imag} */,
  {32'hbfa53774, 32'h00000000} /* (18, 7, 5) {real, imag} */,
  {32'hbf464640, 32'h00000000} /* (18, 7, 4) {real, imag} */,
  {32'hbf0bdb89, 32'h00000000} /* (18, 7, 3) {real, imag} */,
  {32'hbf456670, 32'h00000000} /* (18, 7, 2) {real, imag} */,
  {32'hbf74d75e, 32'h00000000} /* (18, 7, 1) {real, imag} */,
  {32'hbf308bd5, 32'h00000000} /* (18, 7, 0) {real, imag} */,
  {32'hbef0d14d, 32'h00000000} /* (18, 6, 31) {real, imag} */,
  {32'hbf969143, 32'h00000000} /* (18, 6, 30) {real, imag} */,
  {32'hbf943c8a, 32'h00000000} /* (18, 6, 29) {real, imag} */,
  {32'hbe597d56, 32'h00000000} /* (18, 6, 28) {real, imag} */,
  {32'hbdb0c313, 32'h00000000} /* (18, 6, 27) {real, imag} */,
  {32'hbf80bd46, 32'h00000000} /* (18, 6, 26) {real, imag} */,
  {32'hbff785f4, 32'h00000000} /* (18, 6, 25) {real, imag} */,
  {32'hbfb125cc, 32'h00000000} /* (18, 6, 24) {real, imag} */,
  {32'hbf782bcb, 32'h00000000} /* (18, 6, 23) {real, imag} */,
  {32'hbf915faf, 32'h00000000} /* (18, 6, 22) {real, imag} */,
  {32'hbfa4dc3e, 32'h00000000} /* (18, 6, 21) {real, imag} */,
  {32'h3e9a8f4d, 32'h00000000} /* (18, 6, 20) {real, imag} */,
  {32'h3f7098c9, 32'h00000000} /* (18, 6, 19) {real, imag} */,
  {32'h3f99192d, 32'h00000000} /* (18, 6, 18) {real, imag} */,
  {32'h3fa35eee, 32'h00000000} /* (18, 6, 17) {real, imag} */,
  {32'h3f5dafec, 32'h00000000} /* (18, 6, 16) {real, imag} */,
  {32'h3f9870c6, 32'h00000000} /* (18, 6, 15) {real, imag} */,
  {32'h3f7c9402, 32'h00000000} /* (18, 6, 14) {real, imag} */,
  {32'h3f4c7f63, 32'h00000000} /* (18, 6, 13) {real, imag} */,
  {32'h3f88e985, 32'h00000000} /* (18, 6, 12) {real, imag} */,
  {32'h3f32d77f, 32'h00000000} /* (18, 6, 11) {real, imag} */,
  {32'hbba56ad5, 32'h00000000} /* (18, 6, 10) {real, imag} */,
  {32'hbf22b79d, 32'h00000000} /* (18, 6, 9) {real, imag} */,
  {32'hbf405ff5, 32'h00000000} /* (18, 6, 8) {real, imag} */,
  {32'hbf032dc3, 32'h00000000} /* (18, 6, 7) {real, imag} */,
  {32'hbf81263e, 32'h00000000} /* (18, 6, 6) {real, imag} */,
  {32'hbf813b47, 32'h00000000} /* (18, 6, 5) {real, imag} */,
  {32'hbf839371, 32'h00000000} /* (18, 6, 4) {real, imag} */,
  {32'hbfaf9005, 32'h00000000} /* (18, 6, 3) {real, imag} */,
  {32'hbfc82038, 32'h00000000} /* (18, 6, 2) {real, imag} */,
  {32'hbf7bfa22, 32'h00000000} /* (18, 6, 1) {real, imag} */,
  {32'hbecde31e, 32'h00000000} /* (18, 6, 0) {real, imag} */,
  {32'hbeda5640, 32'h00000000} /* (18, 5, 31) {real, imag} */,
  {32'hbf529161, 32'h00000000} /* (18, 5, 30) {real, imag} */,
  {32'hbfb49f5a, 32'h00000000} /* (18, 5, 29) {real, imag} */,
  {32'hbf3e7ad1, 32'h00000000} /* (18, 5, 28) {real, imag} */,
  {32'hbe996266, 32'h00000000} /* (18, 5, 27) {real, imag} */,
  {32'hbf0b8849, 32'h00000000} /* (18, 5, 26) {real, imag} */,
  {32'hbf95ffe2, 32'h00000000} /* (18, 5, 25) {real, imag} */,
  {32'hbf835fae, 32'h00000000} /* (18, 5, 24) {real, imag} */,
  {32'hbfa65d0a, 32'h00000000} /* (18, 5, 23) {real, imag} */,
  {32'hbfac4c6a, 32'h00000000} /* (18, 5, 22) {real, imag} */,
  {32'hbf26e3a7, 32'h00000000} /* (18, 5, 21) {real, imag} */,
  {32'hbeff8555, 32'h00000000} /* (18, 5, 20) {real, imag} */,
  {32'hbf434b86, 32'h00000000} /* (18, 5, 19) {real, imag} */,
  {32'hbef19f54, 32'h00000000} /* (18, 5, 18) {real, imag} */,
  {32'h3d41dd89, 32'h00000000} /* (18, 5, 17) {real, imag} */,
  {32'h3eaec070, 32'h00000000} /* (18, 5, 16) {real, imag} */,
  {32'h3ee2c783, 32'h00000000} /* (18, 5, 15) {real, imag} */,
  {32'h3ed65c11, 32'h00000000} /* (18, 5, 14) {real, imag} */,
  {32'h3f21f67c, 32'h00000000} /* (18, 5, 13) {real, imag} */,
  {32'h3f2836f8, 32'h00000000} /* (18, 5, 12) {real, imag} */,
  {32'h3f2e8a69, 32'h00000000} /* (18, 5, 11) {real, imag} */,
  {32'h3f54f9c7, 32'h00000000} /* (18, 5, 10) {real, imag} */,
  {32'h3e540105, 32'h00000000} /* (18, 5, 9) {real, imag} */,
  {32'h3db0f72d, 32'h00000000} /* (18, 5, 8) {real, imag} */,
  {32'h3dda59c3, 32'h00000000} /* (18, 5, 7) {real, imag} */,
  {32'hbe3e591a, 32'h00000000} /* (18, 5, 6) {real, imag} */,
  {32'hbeff2e06, 32'h00000000} /* (18, 5, 5) {real, imag} */,
  {32'hbf86064c, 32'h00000000} /* (18, 5, 4) {real, imag} */,
  {32'hbfa02b71, 32'h00000000} /* (18, 5, 3) {real, imag} */,
  {32'hbf9c87a0, 32'h00000000} /* (18, 5, 2) {real, imag} */,
  {32'hbf5a2c68, 32'h00000000} /* (18, 5, 1) {real, imag} */,
  {32'hbeac7917, 32'h00000000} /* (18, 5, 0) {real, imag} */,
  {32'hbedcec59, 32'h00000000} /* (18, 4, 31) {real, imag} */,
  {32'hbf8a6578, 32'h00000000} /* (18, 4, 30) {real, imag} */,
  {32'hbfbf2f07, 32'h00000000} /* (18, 4, 29) {real, imag} */,
  {32'hbf44e991, 32'h00000000} /* (18, 4, 28) {real, imag} */,
  {32'hbec03544, 32'h00000000} /* (18, 4, 27) {real, imag} */,
  {32'hbe8d73a1, 32'h00000000} /* (18, 4, 26) {real, imag} */,
  {32'hbed29409, 32'h00000000} /* (18, 4, 25) {real, imag} */,
  {32'hbf33ac20, 32'h00000000} /* (18, 4, 24) {real, imag} */,
  {32'hbfb55ca2, 32'h00000000} /* (18, 4, 23) {real, imag} */,
  {32'hbfb84458, 32'h00000000} /* (18, 4, 22) {real, imag} */,
  {32'hbfb5a379, 32'h00000000} /* (18, 4, 21) {real, imag} */,
  {32'hbf8eb7e3, 32'h00000000} /* (18, 4, 20) {real, imag} */,
  {32'hbfa911f1, 32'h00000000} /* (18, 4, 19) {real, imag} */,
  {32'hbf6fc1b1, 32'h00000000} /* (18, 4, 18) {real, imag} */,
  {32'hbf71bf9b, 32'h00000000} /* (18, 4, 17) {real, imag} */,
  {32'hbe442190, 32'h00000000} /* (18, 4, 16) {real, imag} */,
  {32'h3ea86345, 32'h00000000} /* (18, 4, 15) {real, imag} */,
  {32'h3ec0aff9, 32'h00000000} /* (18, 4, 14) {real, imag} */,
  {32'h3ed874f0, 32'h00000000} /* (18, 4, 13) {real, imag} */,
  {32'h3f3aae76, 32'h00000000} /* (18, 4, 12) {real, imag} */,
  {32'h3f904e5b, 32'h00000000} /* (18, 4, 11) {real, imag} */,
  {32'h3f90ecab, 32'h00000000} /* (18, 4, 10) {real, imag} */,
  {32'h3f8cf5c7, 32'h00000000} /* (18, 4, 9) {real, imag} */,
  {32'h3f691837, 32'h00000000} /* (18, 4, 8) {real, imag} */,
  {32'h3f511a54, 32'h00000000} /* (18, 4, 7) {real, imag} */,
  {32'h3f0246dd, 32'h00000000} /* (18, 4, 6) {real, imag} */,
  {32'hbf16d486, 32'h00000000} /* (18, 4, 5) {real, imag} */,
  {32'hbfbb96b5, 32'h00000000} /* (18, 4, 4) {real, imag} */,
  {32'hbf84432d, 32'h00000000} /* (18, 4, 3) {real, imag} */,
  {32'hbee84a7b, 32'h00000000} /* (18, 4, 2) {real, imag} */,
  {32'hbf212818, 32'h00000000} /* (18, 4, 1) {real, imag} */,
  {32'hbe192d33, 32'h00000000} /* (18, 4, 0) {real, imag} */,
  {32'hbe9bae5a, 32'h00000000} /* (18, 3, 31) {real, imag} */,
  {32'hbf6fea0d, 32'h00000000} /* (18, 3, 30) {real, imag} */,
  {32'hbf38ac28, 32'h00000000} /* (18, 3, 29) {real, imag} */,
  {32'hbe63f33b, 32'h00000000} /* (18, 3, 28) {real, imag} */,
  {32'hbeb0a2d5, 32'h00000000} /* (18, 3, 27) {real, imag} */,
  {32'hbe9e94f3, 32'h00000000} /* (18, 3, 26) {real, imag} */,
  {32'hbefce80a, 32'h00000000} /* (18, 3, 25) {real, imag} */,
  {32'hbf12c181, 32'h00000000} /* (18, 3, 24) {real, imag} */,
  {32'hbfade6b7, 32'h00000000} /* (18, 3, 23) {real, imag} */,
  {32'hbfdf62e2, 32'h00000000} /* (18, 3, 22) {real, imag} */,
  {32'hbf925cef, 32'h00000000} /* (18, 3, 21) {real, imag} */,
  {32'hbf307e5f, 32'h00000000} /* (18, 3, 20) {real, imag} */,
  {32'hbf8a21cd, 32'h00000000} /* (18, 3, 19) {real, imag} */,
  {32'hbf8a04c3, 32'h00000000} /* (18, 3, 18) {real, imag} */,
  {32'hbf742e2c, 32'h00000000} /* (18, 3, 17) {real, imag} */,
  {32'hbecfbdb0, 32'h00000000} /* (18, 3, 16) {real, imag} */,
  {32'h3f1b9a58, 32'h00000000} /* (18, 3, 15) {real, imag} */,
  {32'h3f471189, 32'h00000000} /* (18, 3, 14) {real, imag} */,
  {32'h3f777e8b, 32'h00000000} /* (18, 3, 13) {real, imag} */,
  {32'h3fa026c6, 32'h00000000} /* (18, 3, 12) {real, imag} */,
  {32'h3f9119c2, 32'h00000000} /* (18, 3, 11) {real, imag} */,
  {32'h3f6342f6, 32'h00000000} /* (18, 3, 10) {real, imag} */,
  {32'h3f8d38f9, 32'h00000000} /* (18, 3, 9) {real, imag} */,
  {32'h3f8a3a2d, 32'h00000000} /* (18, 3, 8) {real, imag} */,
  {32'h3f55a29b, 32'h00000000} /* (18, 3, 7) {real, imag} */,
  {32'h3f4286b4, 32'h00000000} /* (18, 3, 6) {real, imag} */,
  {32'hbeb5c0ed, 32'h00000000} /* (18, 3, 5) {real, imag} */,
  {32'hbf98098b, 32'h00000000} /* (18, 3, 4) {real, imag} */,
  {32'hbf584bf2, 32'h00000000} /* (18, 3, 3) {real, imag} */,
  {32'hbf3b246d, 32'h00000000} /* (18, 3, 2) {real, imag} */,
  {32'hbf6ded42, 32'h00000000} /* (18, 3, 1) {real, imag} */,
  {32'hbe4f54b2, 32'h00000000} /* (18, 3, 0) {real, imag} */,
  {32'hbecfd4f0, 32'h00000000} /* (18, 2, 31) {real, imag} */,
  {32'hbf83c34e, 32'h00000000} /* (18, 2, 30) {real, imag} */,
  {32'hbef5485e, 32'h00000000} /* (18, 2, 29) {real, imag} */,
  {32'hbe96a1b6, 32'h00000000} /* (18, 2, 28) {real, imag} */,
  {32'hbf316e78, 32'h00000000} /* (18, 2, 27) {real, imag} */,
  {32'hbf1bb284, 32'h00000000} /* (18, 2, 26) {real, imag} */,
  {32'hbf28367a, 32'h00000000} /* (18, 2, 25) {real, imag} */,
  {32'hbf0f36f3, 32'h00000000} /* (18, 2, 24) {real, imag} */,
  {32'hbf990508, 32'h00000000} /* (18, 2, 23) {real, imag} */,
  {32'hbf91a3b7, 32'h00000000} /* (18, 2, 22) {real, imag} */,
  {32'hbf0483d5, 32'h00000000} /* (18, 2, 21) {real, imag} */,
  {32'hbf162fca, 32'h00000000} /* (18, 2, 20) {real, imag} */,
  {32'hbfbd40b2, 32'h00000000} /* (18, 2, 19) {real, imag} */,
  {32'hbff127fc, 32'h00000000} /* (18, 2, 18) {real, imag} */,
  {32'hbfa04b72, 32'h00000000} /* (18, 2, 17) {real, imag} */,
  {32'hbf3f72fd, 32'h00000000} /* (18, 2, 16) {real, imag} */,
  {32'h3ec02bd0, 32'h00000000} /* (18, 2, 15) {real, imag} */,
  {32'h3ef14da8, 32'h00000000} /* (18, 2, 14) {real, imag} */,
  {32'h3f81b1bf, 32'h00000000} /* (18, 2, 13) {real, imag} */,
  {32'h3f57a744, 32'h00000000} /* (18, 2, 12) {real, imag} */,
  {32'h3f3aee8c, 32'h00000000} /* (18, 2, 11) {real, imag} */,
  {32'h3f3d39c8, 32'h00000000} /* (18, 2, 10) {real, imag} */,
  {32'h3f4f3636, 32'h00000000} /* (18, 2, 9) {real, imag} */,
  {32'h3f907fb3, 32'h00000000} /* (18, 2, 8) {real, imag} */,
  {32'h3f7125a5, 32'h00000000} /* (18, 2, 7) {real, imag} */,
  {32'h3f28b292, 32'h00000000} /* (18, 2, 6) {real, imag} */,
  {32'hbef4a8c4, 32'h00000000} /* (18, 2, 5) {real, imag} */,
  {32'hbf6bcd8c, 32'h00000000} /* (18, 2, 4) {real, imag} */,
  {32'hbf5abb91, 32'h00000000} /* (18, 2, 3) {real, imag} */,
  {32'hbf9ae261, 32'h00000000} /* (18, 2, 2) {real, imag} */,
  {32'hbf909f6e, 32'h00000000} /* (18, 2, 1) {real, imag} */,
  {32'hbe3e80ae, 32'h00000000} /* (18, 2, 0) {real, imag} */,
  {32'hbf135662, 32'h00000000} /* (18, 1, 31) {real, imag} */,
  {32'hbf778c0d, 32'h00000000} /* (18, 1, 30) {real, imag} */,
  {32'hbf82fc59, 32'h00000000} /* (18, 1, 29) {real, imag} */,
  {32'hbf1d5ee6, 32'h00000000} /* (18, 1, 28) {real, imag} */,
  {32'hbf120114, 32'h00000000} /* (18, 1, 27) {real, imag} */,
  {32'hbf182ae6, 32'h00000000} /* (18, 1, 26) {real, imag} */,
  {32'hbf4fdecd, 32'h00000000} /* (18, 1, 25) {real, imag} */,
  {32'hbf425ada, 32'h00000000} /* (18, 1, 24) {real, imag} */,
  {32'hbf72e94f, 32'h00000000} /* (18, 1, 23) {real, imag} */,
  {32'hbf476bd0, 32'h00000000} /* (18, 1, 22) {real, imag} */,
  {32'hbf15f2c5, 32'h00000000} /* (18, 1, 21) {real, imag} */,
  {32'hbf4c11ef, 32'h00000000} /* (18, 1, 20) {real, imag} */,
  {32'hbfb4b8bc, 32'h00000000} /* (18, 1, 19) {real, imag} */,
  {32'hc0038b1d, 32'h00000000} /* (18, 1, 18) {real, imag} */,
  {32'hbfcf0bf2, 32'h00000000} /* (18, 1, 17) {real, imag} */,
  {32'hbf16cc5c, 32'h00000000} /* (18, 1, 16) {real, imag} */,
  {32'h3edec1ec, 32'h00000000} /* (18, 1, 15) {real, imag} */,
  {32'h3f2716fa, 32'h00000000} /* (18, 1, 14) {real, imag} */,
  {32'h3f67d7a2, 32'h00000000} /* (18, 1, 13) {real, imag} */,
  {32'h3f56e6f4, 32'h00000000} /* (18, 1, 12) {real, imag} */,
  {32'h3f665c0d, 32'h00000000} /* (18, 1, 11) {real, imag} */,
  {32'h3f217fe9, 32'h00000000} /* (18, 1, 10) {real, imag} */,
  {32'h3f094701, 32'h00000000} /* (18, 1, 9) {real, imag} */,
  {32'h3f670013, 32'h00000000} /* (18, 1, 8) {real, imag} */,
  {32'h3f2e17e1, 32'h00000000} /* (18, 1, 7) {real, imag} */,
  {32'h3ede4ceb, 32'h00000000} /* (18, 1, 6) {real, imag} */,
  {32'hbd045559, 32'h00000000} /* (18, 1, 5) {real, imag} */,
  {32'hbf19c8fd, 32'h00000000} /* (18, 1, 4) {real, imag} */,
  {32'hbf878ab9, 32'h00000000} /* (18, 1, 3) {real, imag} */,
  {32'hbfb9045f, 32'h00000000} /* (18, 1, 2) {real, imag} */,
  {32'hbf857370, 32'h00000000} /* (18, 1, 1) {real, imag} */,
  {32'hbe83f363, 32'h00000000} /* (18, 1, 0) {real, imag} */,
  {32'hbf0e3063, 32'h00000000} /* (18, 0, 31) {real, imag} */,
  {32'hbf00218d, 32'h00000000} /* (18, 0, 30) {real, imag} */,
  {32'hbf136430, 32'h00000000} /* (18, 0, 29) {real, imag} */,
  {32'hbee436f4, 32'h00000000} /* (18, 0, 28) {real, imag} */,
  {32'hbea0283a, 32'h00000000} /* (18, 0, 27) {real, imag} */,
  {32'hbedc00b2, 32'h00000000} /* (18, 0, 26) {real, imag} */,
  {32'hbec0c07a, 32'h00000000} /* (18, 0, 25) {real, imag} */,
  {32'hbe8fbf87, 32'h00000000} /* (18, 0, 24) {real, imag} */,
  {32'hbe8f9602, 32'h00000000} /* (18, 0, 23) {real, imag} */,
  {32'hbee6cb3b, 32'h00000000} /* (18, 0, 22) {real, imag} */,
  {32'hbf2b4cc7, 32'h00000000} /* (18, 0, 21) {real, imag} */,
  {32'hbf1d6538, 32'h00000000} /* (18, 0, 20) {real, imag} */,
  {32'hbebd2f97, 32'h00000000} /* (18, 0, 19) {real, imag} */,
  {32'hbf0fcfa0, 32'h00000000} /* (18, 0, 18) {real, imag} */,
  {32'hbf1fe087, 32'h00000000} /* (18, 0, 17) {real, imag} */,
  {32'hbd9603ff, 32'h00000000} /* (18, 0, 16) {real, imag} */,
  {32'h3edda445, 32'h00000000} /* (18, 0, 15) {real, imag} */,
  {32'h3eb6f3c0, 32'h00000000} /* (18, 0, 14) {real, imag} */,
  {32'h3ee31e5a, 32'h00000000} /* (18, 0, 13) {real, imag} */,
  {32'h3f1b9566, 32'h00000000} /* (18, 0, 12) {real, imag} */,
  {32'h3f3e0542, 32'h00000000} /* (18, 0, 11) {real, imag} */,
  {32'h3ee8785c, 32'h00000000} /* (18, 0, 10) {real, imag} */,
  {32'h3e8c969c, 32'h00000000} /* (18, 0, 9) {real, imag} */,
  {32'h3f0b8c93, 32'h00000000} /* (18, 0, 8) {real, imag} */,
  {32'h3f0a1f16, 32'h00000000} /* (18, 0, 7) {real, imag} */,
  {32'h3ead554a, 32'h00000000} /* (18, 0, 6) {real, imag} */,
  {32'h3e9361b9, 32'h00000000} /* (18, 0, 5) {real, imag} */,
  {32'hbd327d54, 32'h00000000} /* (18, 0, 4) {real, imag} */,
  {32'hbeed1381, 32'h00000000} /* (18, 0, 3) {real, imag} */,
  {32'hbf459dfb, 32'h00000000} /* (18, 0, 2) {real, imag} */,
  {32'hbf5fc15d, 32'h00000000} /* (18, 0, 1) {real, imag} */,
  {32'hbeb3e596, 32'h00000000} /* (18, 0, 0) {real, imag} */,
  {32'hbe2f87ea, 32'h00000000} /* (17, 31, 31) {real, imag} */,
  {32'hbea12217, 32'h00000000} /* (17, 31, 30) {real, imag} */,
  {32'hbef5becf, 32'h00000000} /* (17, 31, 29) {real, imag} */,
  {32'hbeffc5e9, 32'h00000000} /* (17, 31, 28) {real, imag} */,
  {32'hbeb55e04, 32'h00000000} /* (17, 31, 27) {real, imag} */,
  {32'hbe832be9, 32'h00000000} /* (17, 31, 26) {real, imag} */,
  {32'hbf314415, 32'h00000000} /* (17, 31, 25) {real, imag} */,
  {32'hbf389dfc, 32'h00000000} /* (17, 31, 24) {real, imag} */,
  {32'hbf143938, 32'h00000000} /* (17, 31, 23) {real, imag} */,
  {32'hbf2de00c, 32'h00000000} /* (17, 31, 22) {real, imag} */,
  {32'hbf2b1bc3, 32'h00000000} /* (17, 31, 21) {real, imag} */,
  {32'hbe1d4426, 32'h00000000} /* (17, 31, 20) {real, imag} */,
  {32'h3e08993d, 32'h00000000} /* (17, 31, 19) {real, imag} */,
  {32'h3e521215, 32'h00000000} /* (17, 31, 18) {real, imag} */,
  {32'h3ef06759, 32'h00000000} /* (17, 31, 17) {real, imag} */,
  {32'h3e622140, 32'h00000000} /* (17, 31, 16) {real, imag} */,
  {32'h3ef3e912, 32'h00000000} /* (17, 31, 15) {real, imag} */,
  {32'h3ee6f5f9, 32'h00000000} /* (17, 31, 14) {real, imag} */,
  {32'h3eaaf78d, 32'h00000000} /* (17, 31, 13) {real, imag} */,
  {32'h3ee1f5da, 32'h00000000} /* (17, 31, 12) {real, imag} */,
  {32'h3f10176f, 32'h00000000} /* (17, 31, 11) {real, imag} */,
  {32'h3df18c75, 32'h00000000} /* (17, 31, 10) {real, imag} */,
  {32'hbeaaf8be, 32'h00000000} /* (17, 31, 9) {real, imag} */,
  {32'hbeeec4d4, 32'h00000000} /* (17, 31, 8) {real, imag} */,
  {32'hbf188845, 32'h00000000} /* (17, 31, 7) {real, imag} */,
  {32'hbed34f14, 32'h00000000} /* (17, 31, 6) {real, imag} */,
  {32'hbf1bb8cf, 32'h00000000} /* (17, 31, 5) {real, imag} */,
  {32'hbefc2361, 32'h00000000} /* (17, 31, 4) {real, imag} */,
  {32'hbf139d91, 32'h00000000} /* (17, 31, 3) {real, imag} */,
  {32'hbf159f00, 32'h00000000} /* (17, 31, 2) {real, imag} */,
  {32'hbea23e02, 32'h00000000} /* (17, 31, 1) {real, imag} */,
  {32'hbd9eb01b, 32'h00000000} /* (17, 31, 0) {real, imag} */,
  {32'hbed09724, 32'h00000000} /* (17, 30, 31) {real, imag} */,
  {32'hbf80bd03, 32'h00000000} /* (17, 30, 30) {real, imag} */,
  {32'hbfc222fa, 32'h00000000} /* (17, 30, 29) {real, imag} */,
  {32'hbf8ee182, 32'h00000000} /* (17, 30, 28) {real, imag} */,
  {32'hbf0f9044, 32'h00000000} /* (17, 30, 27) {real, imag} */,
  {32'hbea2bb5d, 32'h00000000} /* (17, 30, 26) {real, imag} */,
  {32'hbf25233e, 32'h00000000} /* (17, 30, 25) {real, imag} */,
  {32'hbf784bf5, 32'h00000000} /* (17, 30, 24) {real, imag} */,
  {32'hbf46f826, 32'h00000000} /* (17, 30, 23) {real, imag} */,
  {32'hbf84e806, 32'h00000000} /* (17, 30, 22) {real, imag} */,
  {32'hbf53aaf3, 32'h00000000} /* (17, 30, 21) {real, imag} */,
  {32'h3f47b375, 32'h00000000} /* (17, 30, 20) {real, imag} */,
  {32'h3f93c994, 32'h00000000} /* (17, 30, 19) {real, imag} */,
  {32'h3f2afe36, 32'h00000000} /* (17, 30, 18) {real, imag} */,
  {32'h3f4c03c2, 32'h00000000} /* (17, 30, 17) {real, imag} */,
  {32'h3f56139a, 32'h00000000} /* (17, 30, 16) {real, imag} */,
  {32'h3f939be1, 32'h00000000} /* (17, 30, 15) {real, imag} */,
  {32'h3f748818, 32'h00000000} /* (17, 30, 14) {real, imag} */,
  {32'h3f77601d, 32'h00000000} /* (17, 30, 13) {real, imag} */,
  {32'h3f6d59bd, 32'h00000000} /* (17, 30, 12) {real, imag} */,
  {32'h3f0486d2, 32'h00000000} /* (17, 30, 11) {real, imag} */,
  {32'hbebcbc36, 32'h00000000} /* (17, 30, 10) {real, imag} */,
  {32'hbf78cee4, 32'h00000000} /* (17, 30, 9) {real, imag} */,
  {32'hbf94c579, 32'h00000000} /* (17, 30, 8) {real, imag} */,
  {32'hbf967159, 32'h00000000} /* (17, 30, 7) {real, imag} */,
  {32'hbf8d517f, 32'h00000000} /* (17, 30, 6) {real, imag} */,
  {32'hbf7bb548, 32'h00000000} /* (17, 30, 5) {real, imag} */,
  {32'hbf86bf75, 32'h00000000} /* (17, 30, 4) {real, imag} */,
  {32'hbf717671, 32'h00000000} /* (17, 30, 3) {real, imag} */,
  {32'hbf9f1438, 32'h00000000} /* (17, 30, 2) {real, imag} */,
  {32'hbf147040, 32'h00000000} /* (17, 30, 1) {real, imag} */,
  {32'hbe88be67, 32'h00000000} /* (17, 30, 0) {real, imag} */,
  {32'hbf339d87, 32'h00000000} /* (17, 29, 31) {real, imag} */,
  {32'hbfba5b7a, 32'h00000000} /* (17, 29, 30) {real, imag} */,
  {32'hbfc9f86e, 32'h00000000} /* (17, 29, 29) {real, imag} */,
  {32'hbf8a3527, 32'h00000000} /* (17, 29, 28) {real, imag} */,
  {32'hbf3147a7, 32'h00000000} /* (17, 29, 27) {real, imag} */,
  {32'hbee6f06e, 32'h00000000} /* (17, 29, 26) {real, imag} */,
  {32'hbf537b00, 32'h00000000} /* (17, 29, 25) {real, imag} */,
  {32'hbfb7b931, 32'h00000000} /* (17, 29, 24) {real, imag} */,
  {32'hbf992831, 32'h00000000} /* (17, 29, 23) {real, imag} */,
  {32'hbf825bcd, 32'h00000000} /* (17, 29, 22) {real, imag} */,
  {32'hbefc24b2, 32'h00000000} /* (17, 29, 21) {real, imag} */,
  {32'h3f796563, 32'h00000000} /* (17, 29, 20) {real, imag} */,
  {32'h3f7cbe6e, 32'h00000000} /* (17, 29, 19) {real, imag} */,
  {32'h3f517b87, 32'h00000000} /* (17, 29, 18) {real, imag} */,
  {32'h3fc25f0c, 32'h00000000} /* (17, 29, 17) {real, imag} */,
  {32'h3fcf258f, 32'h00000000} /* (17, 29, 16) {real, imag} */,
  {32'h3fb151be, 32'h00000000} /* (17, 29, 15) {real, imag} */,
  {32'h3f718e6e, 32'h00000000} /* (17, 29, 14) {real, imag} */,
  {32'h3fab67e6, 32'h00000000} /* (17, 29, 13) {real, imag} */,
  {32'h3f8e7ebb, 32'h00000000} /* (17, 29, 12) {real, imag} */,
  {32'h3ef4dc96, 32'h00000000} /* (17, 29, 11) {real, imag} */,
  {32'hbe9d9132, 32'h00000000} /* (17, 29, 10) {real, imag} */,
  {32'hbf87f0f8, 32'h00000000} /* (17, 29, 9) {real, imag} */,
  {32'hbfcff0dc, 32'h00000000} /* (17, 29, 8) {real, imag} */,
  {32'hbf97b5cf, 32'h00000000} /* (17, 29, 7) {real, imag} */,
  {32'hbf7d36e4, 32'h00000000} /* (17, 29, 6) {real, imag} */,
  {32'hbf669699, 32'h00000000} /* (17, 29, 5) {real, imag} */,
  {32'hbf8fa725, 32'h00000000} /* (17, 29, 4) {real, imag} */,
  {32'hbf83373c, 32'h00000000} /* (17, 29, 3) {real, imag} */,
  {32'hbf8af19c, 32'h00000000} /* (17, 29, 2) {real, imag} */,
  {32'hbf4f394b, 32'h00000000} /* (17, 29, 1) {real, imag} */,
  {32'hbf583229, 32'h00000000} /* (17, 29, 0) {real, imag} */,
  {32'hbf45b4de, 32'h00000000} /* (17, 28, 31) {real, imag} */,
  {32'hbfb1dc2b, 32'h00000000} /* (17, 28, 30) {real, imag} */,
  {32'hbf88364a, 32'h00000000} /* (17, 28, 29) {real, imag} */,
  {32'hbf6814f3, 32'h00000000} /* (17, 28, 28) {real, imag} */,
  {32'hbf6a6ec0, 32'h00000000} /* (17, 28, 27) {real, imag} */,
  {32'hbf10d158, 32'h00000000} /* (17, 28, 26) {real, imag} */,
  {32'hbf987112, 32'h00000000} /* (17, 28, 25) {real, imag} */,
  {32'hbfc9d25e, 32'h00000000} /* (17, 28, 24) {real, imag} */,
  {32'hbfb13c31, 32'h00000000} /* (17, 28, 23) {real, imag} */,
  {32'hbf52da6a, 32'h00000000} /* (17, 28, 22) {real, imag} */,
  {32'hbea99612, 32'h00000000} /* (17, 28, 21) {real, imag} */,
  {32'h3e8274f5, 32'h00000000} /* (17, 28, 20) {real, imag} */,
  {32'h3f0cb0c9, 32'h00000000} /* (17, 28, 19) {real, imag} */,
  {32'h3f977018, 32'h00000000} /* (17, 28, 18) {real, imag} */,
  {32'h3fc01ffe, 32'h00000000} /* (17, 28, 17) {real, imag} */,
  {32'h3fa40682, 32'h00000000} /* (17, 28, 16) {real, imag} */,
  {32'h3f9aa413, 32'h00000000} /* (17, 28, 15) {real, imag} */,
  {32'h3f8468d1, 32'h00000000} /* (17, 28, 14) {real, imag} */,
  {32'h3f89a718, 32'h00000000} /* (17, 28, 13) {real, imag} */,
  {32'h3f88ec12, 32'h00000000} /* (17, 28, 12) {real, imag} */,
  {32'h3f83a08a, 32'h00000000} /* (17, 28, 11) {real, imag} */,
  {32'hbe28b727, 32'h00000000} /* (17, 28, 10) {real, imag} */,
  {32'hbf73ec99, 32'h00000000} /* (17, 28, 9) {real, imag} */,
  {32'hbf5e2dd7, 32'h00000000} /* (17, 28, 8) {real, imag} */,
  {32'hbf83bcc8, 32'h00000000} /* (17, 28, 7) {real, imag} */,
  {32'hbf8d24d7, 32'h00000000} /* (17, 28, 6) {real, imag} */,
  {32'hbf73b487, 32'h00000000} /* (17, 28, 5) {real, imag} */,
  {32'hbf93a39e, 32'h00000000} /* (17, 28, 4) {real, imag} */,
  {32'hbf999fea, 32'h00000000} /* (17, 28, 3) {real, imag} */,
  {32'hbfab7fe4, 32'h00000000} /* (17, 28, 2) {real, imag} */,
  {32'hbf8e7a47, 32'h00000000} /* (17, 28, 1) {real, imag} */,
  {32'hbf0c9baa, 32'h00000000} /* (17, 28, 0) {real, imag} */,
  {32'hbf7304a1, 32'h00000000} /* (17, 27, 31) {real, imag} */,
  {32'hbfb9ea70, 32'h00000000} /* (17, 27, 30) {real, imag} */,
  {32'hbf4a38ef, 32'h00000000} /* (17, 27, 29) {real, imag} */,
  {32'hbec0a354, 32'h00000000} /* (17, 27, 28) {real, imag} */,
  {32'hbefed619, 32'h00000000} /* (17, 27, 27) {real, imag} */,
  {32'hbf3539e7, 32'h00000000} /* (17, 27, 26) {real, imag} */,
  {32'hbf7136a2, 32'h00000000} /* (17, 27, 25) {real, imag} */,
  {32'hbf950cc0, 32'h00000000} /* (17, 27, 24) {real, imag} */,
  {32'hbfc9d1c4, 32'h00000000} /* (17, 27, 23) {real, imag} */,
  {32'hbf9d78b7, 32'h00000000} /* (17, 27, 22) {real, imag} */,
  {32'hbf270748, 32'h00000000} /* (17, 27, 21) {real, imag} */,
  {32'h3ebe3bf3, 32'h00000000} /* (17, 27, 20) {real, imag} */,
  {32'h3f421ae3, 32'h00000000} /* (17, 27, 19) {real, imag} */,
  {32'h3fa7223c, 32'h00000000} /* (17, 27, 18) {real, imag} */,
  {32'h3fc23680, 32'h00000000} /* (17, 27, 17) {real, imag} */,
  {32'h3f8cce85, 32'h00000000} /* (17, 27, 16) {real, imag} */,
  {32'h3f66eacf, 32'h00000000} /* (17, 27, 15) {real, imag} */,
  {32'h3f83340d, 32'h00000000} /* (17, 27, 14) {real, imag} */,
  {32'h3f7f0700, 32'h00000000} /* (17, 27, 13) {real, imag} */,
  {32'h3f65998f, 32'h00000000} /* (17, 27, 12) {real, imag} */,
  {32'h3f8e4bd7, 32'h00000000} /* (17, 27, 11) {real, imag} */,
  {32'hbeda4a37, 32'h00000000} /* (17, 27, 10) {real, imag} */,
  {32'hbf8a54f0, 32'h00000000} /* (17, 27, 9) {real, imag} */,
  {32'hbf84a8d4, 32'h00000000} /* (17, 27, 8) {real, imag} */,
  {32'hbfb388eb, 32'h00000000} /* (17, 27, 7) {real, imag} */,
  {32'hbfaf3c22, 32'h00000000} /* (17, 27, 6) {real, imag} */,
  {32'hbfbab606, 32'h00000000} /* (17, 27, 5) {real, imag} */,
  {32'hbfcb7e4e, 32'h00000000} /* (17, 27, 4) {real, imag} */,
  {32'hbf88093d, 32'h00000000} /* (17, 27, 3) {real, imag} */,
  {32'hbfa2fd5d, 32'h00000000} /* (17, 27, 2) {real, imag} */,
  {32'hbf97aca1, 32'h00000000} /* (17, 27, 1) {real, imag} */,
  {32'hbece70e6, 32'h00000000} /* (17, 27, 0) {real, imag} */,
  {32'hbf0e8728, 32'h00000000} /* (17, 26, 31) {real, imag} */,
  {32'hbf7c551e, 32'h00000000} /* (17, 26, 30) {real, imag} */,
  {32'hbee25cee, 32'h00000000} /* (17, 26, 29) {real, imag} */,
  {32'hbe531f58, 32'h00000000} /* (17, 26, 28) {real, imag} */,
  {32'hbedcd199, 32'h00000000} /* (17, 26, 27) {real, imag} */,
  {32'hbf6ca4cf, 32'h00000000} /* (17, 26, 26) {real, imag} */,
  {32'hbf530377, 32'h00000000} /* (17, 26, 25) {real, imag} */,
  {32'hbf38ec26, 32'h00000000} /* (17, 26, 24) {real, imag} */,
  {32'hbf6c744b, 32'h00000000} /* (17, 26, 23) {real, imag} */,
  {32'hbf6be251, 32'h00000000} /* (17, 26, 22) {real, imag} */,
  {32'hbed2452b, 32'h00000000} /* (17, 26, 21) {real, imag} */,
  {32'h3f12c840, 32'h00000000} /* (17, 26, 20) {real, imag} */,
  {32'h3f21c0f0, 32'h00000000} /* (17, 26, 19) {real, imag} */,
  {32'h3eb813f2, 32'h00000000} /* (17, 26, 18) {real, imag} */,
  {32'h3f3e3cee, 32'h00000000} /* (17, 26, 17) {real, imag} */,
  {32'h3f801893, 32'h00000000} /* (17, 26, 16) {real, imag} */,
  {32'h3f42e237, 32'h00000000} /* (17, 26, 15) {real, imag} */,
  {32'h3f91a89c, 32'h00000000} /* (17, 26, 14) {real, imag} */,
  {32'h3f865356, 32'h00000000} /* (17, 26, 13) {real, imag} */,
  {32'h3f45f74b, 32'h00000000} /* (17, 26, 12) {real, imag} */,
  {32'h3f3857f3, 32'h00000000} /* (17, 26, 11) {real, imag} */,
  {32'hbf6263ff, 32'h00000000} /* (17, 26, 10) {real, imag} */,
  {32'hbf95cf99, 32'h00000000} /* (17, 26, 9) {real, imag} */,
  {32'hbfb170cc, 32'h00000000} /* (17, 26, 8) {real, imag} */,
  {32'hbf9a12d2, 32'h00000000} /* (17, 26, 7) {real, imag} */,
  {32'hbf8ea6db, 32'h00000000} /* (17, 26, 6) {real, imag} */,
  {32'hbfa91af9, 32'h00000000} /* (17, 26, 5) {real, imag} */,
  {32'hbfa1921e, 32'h00000000} /* (17, 26, 4) {real, imag} */,
  {32'hbf86eea3, 32'h00000000} /* (17, 26, 3) {real, imag} */,
  {32'hbfa487c3, 32'h00000000} /* (17, 26, 2) {real, imag} */,
  {32'hbf9f67b0, 32'h00000000} /* (17, 26, 1) {real, imag} */,
  {32'hbf219fc7, 32'h00000000} /* (17, 26, 0) {real, imag} */,
  {32'hbee853ce, 32'h00000000} /* (17, 25, 31) {real, imag} */,
  {32'hbf90eebb, 32'h00000000} /* (17, 25, 30) {real, imag} */,
  {32'hbf52f586, 32'h00000000} /* (17, 25, 29) {real, imag} */,
  {32'hbf159a08, 32'h00000000} /* (17, 25, 28) {real, imag} */,
  {32'hbf36b035, 32'h00000000} /* (17, 25, 27) {real, imag} */,
  {32'hbf7044f0, 32'h00000000} /* (17, 25, 26) {real, imag} */,
  {32'hbf129cda, 32'h00000000} /* (17, 25, 25) {real, imag} */,
  {32'hbf1252c6, 32'h00000000} /* (17, 25, 24) {real, imag} */,
  {32'hbf3d3376, 32'h00000000} /* (17, 25, 23) {real, imag} */,
  {32'hbf4d2933, 32'h00000000} /* (17, 25, 22) {real, imag} */,
  {32'hbe009025, 32'h00000000} /* (17, 25, 21) {real, imag} */,
  {32'h3faa8bb8, 32'h00000000} /* (17, 25, 20) {real, imag} */,
  {32'h3fa138d6, 32'h00000000} /* (17, 25, 19) {real, imag} */,
  {32'h3e2eac90, 32'h00000000} /* (17, 25, 18) {real, imag} */,
  {32'h3ecf62cf, 32'h00000000} /* (17, 25, 17) {real, imag} */,
  {32'h3f7efd33, 32'h00000000} /* (17, 25, 16) {real, imag} */,
  {32'h3f6b3628, 32'h00000000} /* (17, 25, 15) {real, imag} */,
  {32'h3f1ad1cf, 32'h00000000} /* (17, 25, 14) {real, imag} */,
  {32'h3f5fee99, 32'h00000000} /* (17, 25, 13) {real, imag} */,
  {32'h3fa18b5f, 32'h00000000} /* (17, 25, 12) {real, imag} */,
  {32'h3f84684f, 32'h00000000} /* (17, 25, 11) {real, imag} */,
  {32'hbf783683, 32'h00000000} /* (17, 25, 10) {real, imag} */,
  {32'hbf9bd32c, 32'h00000000} /* (17, 25, 9) {real, imag} */,
  {32'hbf6cf520, 32'h00000000} /* (17, 25, 8) {real, imag} */,
  {32'hbf4127cd, 32'h00000000} /* (17, 25, 7) {real, imag} */,
  {32'hbf5bb9b4, 32'h00000000} /* (17, 25, 6) {real, imag} */,
  {32'hbf4ef32a, 32'h00000000} /* (17, 25, 5) {real, imag} */,
  {32'hbf34cf99, 32'h00000000} /* (17, 25, 4) {real, imag} */,
  {32'hbf96e038, 32'h00000000} /* (17, 25, 3) {real, imag} */,
  {32'hbfb28baa, 32'h00000000} /* (17, 25, 2) {real, imag} */,
  {32'hbfc5bc51, 32'h00000000} /* (17, 25, 1) {real, imag} */,
  {32'hbf23e5ae, 32'h00000000} /* (17, 25, 0) {real, imag} */,
  {32'hbf0f3122, 32'h00000000} /* (17, 24, 31) {real, imag} */,
  {32'hbf811143, 32'h00000000} /* (17, 24, 30) {real, imag} */,
  {32'hbf52d768, 32'h00000000} /* (17, 24, 29) {real, imag} */,
  {32'hbf8a6ac7, 32'h00000000} /* (17, 24, 28) {real, imag} */,
  {32'hbf8d64cf, 32'h00000000} /* (17, 24, 27) {real, imag} */,
  {32'hbfa29214, 32'h00000000} /* (17, 24, 26) {real, imag} */,
  {32'hbf25602c, 32'h00000000} /* (17, 24, 25) {real, imag} */,
  {32'hbf17a500, 32'h00000000} /* (17, 24, 24) {real, imag} */,
  {32'hbf60b92d, 32'h00000000} /* (17, 24, 23) {real, imag} */,
  {32'hbfa7f49e, 32'h00000000} /* (17, 24, 22) {real, imag} */,
  {32'hbe9305c6, 32'h00000000} /* (17, 24, 21) {real, imag} */,
  {32'h3fd06255, 32'h00000000} /* (17, 24, 20) {real, imag} */,
  {32'h3fafe7b5, 32'h00000000} /* (17, 24, 19) {real, imag} */,
  {32'h3ed0a2db, 32'h00000000} /* (17, 24, 18) {real, imag} */,
  {32'h3f6e11d6, 32'h00000000} /* (17, 24, 17) {real, imag} */,
  {32'h3f30cd33, 32'h00000000} /* (17, 24, 16) {real, imag} */,
  {32'h3ef3ef45, 32'h00000000} /* (17, 24, 15) {real, imag} */,
  {32'h3ebfd769, 32'h00000000} /* (17, 24, 14) {real, imag} */,
  {32'h3f8cb834, 32'h00000000} /* (17, 24, 13) {real, imag} */,
  {32'h3f94fc2b, 32'h00000000} /* (17, 24, 12) {real, imag} */,
  {32'h3f0360ec, 32'h00000000} /* (17, 24, 11) {real, imag} */,
  {32'hbfa2c0df, 32'h00000000} /* (17, 24, 10) {real, imag} */,
  {32'hbfafb9ee, 32'h00000000} /* (17, 24, 9) {real, imag} */,
  {32'hbf8e2440, 32'h00000000} /* (17, 24, 8) {real, imag} */,
  {32'hbf8408a2, 32'h00000000} /* (17, 24, 7) {real, imag} */,
  {32'hbf6f0f04, 32'h00000000} /* (17, 24, 6) {real, imag} */,
  {32'hbf193729, 32'h00000000} /* (17, 24, 5) {real, imag} */,
  {32'hbf00a030, 32'h00000000} /* (17, 24, 4) {real, imag} */,
  {32'hbf9c4290, 32'h00000000} /* (17, 24, 3) {real, imag} */,
  {32'hbfc34cf4, 32'h00000000} /* (17, 24, 2) {real, imag} */,
  {32'hbfc0804a, 32'h00000000} /* (17, 24, 1) {real, imag} */,
  {32'hbf172b50, 32'h00000000} /* (17, 24, 0) {real, imag} */,
  {32'hbea4028d, 32'h00000000} /* (17, 23, 31) {real, imag} */,
  {32'hbf067cf1, 32'h00000000} /* (17, 23, 30) {real, imag} */,
  {32'hbf8595e6, 32'h00000000} /* (17, 23, 29) {real, imag} */,
  {32'hbfc287a2, 32'h00000000} /* (17, 23, 28) {real, imag} */,
  {32'hbf933db1, 32'h00000000} /* (17, 23, 27) {real, imag} */,
  {32'hbf8d880c, 32'h00000000} /* (17, 23, 26) {real, imag} */,
  {32'hbf3e5653, 32'h00000000} /* (17, 23, 25) {real, imag} */,
  {32'hbe96e2f3, 32'h00000000} /* (17, 23, 24) {real, imag} */,
  {32'hbf48946e, 32'h00000000} /* (17, 23, 23) {real, imag} */,
  {32'hbf5f1d58, 32'h00000000} /* (17, 23, 22) {real, imag} */,
  {32'hbd25f971, 32'h00000000} /* (17, 23, 21) {real, imag} */,
  {32'h3f96c72c, 32'h00000000} /* (17, 23, 20) {real, imag} */,
  {32'h3f55cc48, 32'h00000000} /* (17, 23, 19) {real, imag} */,
  {32'h3f1a2d78, 32'h00000000} /* (17, 23, 18) {real, imag} */,
  {32'h3f590f64, 32'h00000000} /* (17, 23, 17) {real, imag} */,
  {32'h3f368450, 32'h00000000} /* (17, 23, 16) {real, imag} */,
  {32'h3f5bbf31, 32'h00000000} /* (17, 23, 15) {real, imag} */,
  {32'h3f35dcfd, 32'h00000000} /* (17, 23, 14) {real, imag} */,
  {32'h3f96e0c1, 32'h00000000} /* (17, 23, 13) {real, imag} */,
  {32'h3f6f4924, 32'h00000000} /* (17, 23, 12) {real, imag} */,
  {32'h3e96586e, 32'h00000000} /* (17, 23, 11) {real, imag} */,
  {32'hbf3ada27, 32'h00000000} /* (17, 23, 10) {real, imag} */,
  {32'hbf8bd8b8, 32'h00000000} /* (17, 23, 9) {real, imag} */,
  {32'hbf989a36, 32'h00000000} /* (17, 23, 8) {real, imag} */,
  {32'hbf6cb8b5, 32'h00000000} /* (17, 23, 7) {real, imag} */,
  {32'hbf7feb1b, 32'h00000000} /* (17, 23, 6) {real, imag} */,
  {32'hbf8a01af, 32'h00000000} /* (17, 23, 5) {real, imag} */,
  {32'hbf39f64f, 32'h00000000} /* (17, 23, 4) {real, imag} */,
  {32'hbf6b8438, 32'h00000000} /* (17, 23, 3) {real, imag} */,
  {32'hbfa7b1ec, 32'h00000000} /* (17, 23, 2) {real, imag} */,
  {32'hbf68634d, 32'h00000000} /* (17, 23, 1) {real, imag} */,
  {32'hbea0224c, 32'h00000000} /* (17, 23, 0) {real, imag} */,
  {32'hbf2ab7bc, 32'h00000000} /* (17, 22, 31) {real, imag} */,
  {32'hbf2d4b68, 32'h00000000} /* (17, 22, 30) {real, imag} */,
  {32'hbf16924d, 32'h00000000} /* (17, 22, 29) {real, imag} */,
  {32'hbf6cddd1, 32'h00000000} /* (17, 22, 28) {real, imag} */,
  {32'hbf3c294e, 32'h00000000} /* (17, 22, 27) {real, imag} */,
  {32'hbf18d5c6, 32'h00000000} /* (17, 22, 26) {real, imag} */,
  {32'hbf0097c6, 32'h00000000} /* (17, 22, 25) {real, imag} */,
  {32'hbecdf7b7, 32'h00000000} /* (17, 22, 24) {real, imag} */,
  {32'hbf4e265d, 32'h00000000} /* (17, 22, 23) {real, imag} */,
  {32'hbf82bb99, 32'h00000000} /* (17, 22, 22) {real, imag} */,
  {32'hbf011071, 32'h00000000} /* (17, 22, 21) {real, imag} */,
  {32'h3f021023, 32'h00000000} /* (17, 22, 20) {real, imag} */,
  {32'h3f0776dd, 32'h00000000} /* (17, 22, 19) {real, imag} */,
  {32'h3f3ab2ad, 32'h00000000} /* (17, 22, 18) {real, imag} */,
  {32'h3f8143b1, 32'h00000000} /* (17, 22, 17) {real, imag} */,
  {32'h3f3ae80b, 32'h00000000} /* (17, 22, 16) {real, imag} */,
  {32'h3f6f0113, 32'h00000000} /* (17, 22, 15) {real, imag} */,
  {32'h3f5e2c82, 32'h00000000} /* (17, 22, 14) {real, imag} */,
  {32'h3f4ba3d2, 32'h00000000} /* (17, 22, 13) {real, imag} */,
  {32'h3f483d34, 32'h00000000} /* (17, 22, 12) {real, imag} */,
  {32'h3f40435d, 32'h00000000} /* (17, 22, 11) {real, imag} */,
  {32'hbe95bdef, 32'h00000000} /* (17, 22, 10) {real, imag} */,
  {32'hbf52505a, 32'h00000000} /* (17, 22, 9) {real, imag} */,
  {32'hbf871356, 32'h00000000} /* (17, 22, 8) {real, imag} */,
  {32'hbf452a76, 32'h00000000} /* (17, 22, 7) {real, imag} */,
  {32'hbf44e5d3, 32'h00000000} /* (17, 22, 6) {real, imag} */,
  {32'hbf60042f, 32'h00000000} /* (17, 22, 5) {real, imag} */,
  {32'hbf5a3da0, 32'h00000000} /* (17, 22, 4) {real, imag} */,
  {32'hbf228a8a, 32'h00000000} /* (17, 22, 3) {real, imag} */,
  {32'hbf62b935, 32'h00000000} /* (17, 22, 2) {real, imag} */,
  {32'hbf62fee5, 32'h00000000} /* (17, 22, 1) {real, imag} */,
  {32'hbf12c9ad, 32'h00000000} /* (17, 22, 0) {real, imag} */,
  {32'hbeb01174, 32'h00000000} /* (17, 21, 31) {real, imag} */,
  {32'hbf5436cc, 32'h00000000} /* (17, 21, 30) {real, imag} */,
  {32'hbf29192b, 32'h00000000} /* (17, 21, 29) {real, imag} */,
  {32'hbee39dd4, 32'h00000000} /* (17, 21, 28) {real, imag} */,
  {32'hbf69b9cf, 32'h00000000} /* (17, 21, 27) {real, imag} */,
  {32'hbf3ebcd9, 32'h00000000} /* (17, 21, 26) {real, imag} */,
  {32'hbe5de718, 32'h00000000} /* (17, 21, 25) {real, imag} */,
  {32'hbe8be717, 32'h00000000} /* (17, 21, 24) {real, imag} */,
  {32'hbedddc96, 32'h00000000} /* (17, 21, 23) {real, imag} */,
  {32'hbf00a50e, 32'h00000000} /* (17, 21, 22) {real, imag} */,
  {32'hbec6ab73, 32'h00000000} /* (17, 21, 21) {real, imag} */,
  {32'h3e8406d2, 32'h00000000} /* (17, 21, 20) {real, imag} */,
  {32'h3f38c846, 32'h00000000} /* (17, 21, 19) {real, imag} */,
  {32'h3ecca770, 32'h00000000} /* (17, 21, 18) {real, imag} */,
  {32'h3ea90ef7, 32'h00000000} /* (17, 21, 17) {real, imag} */,
  {32'h3e2854f1, 32'h00000000} /* (17, 21, 16) {real, imag} */,
  {32'h3f14255d, 32'h00000000} /* (17, 21, 15) {real, imag} */,
  {32'h3ec3655c, 32'h00000000} /* (17, 21, 14) {real, imag} */,
  {32'h3e0a9495, 32'h00000000} /* (17, 21, 13) {real, imag} */,
  {32'h3e5e1759, 32'h00000000} /* (17, 21, 12) {real, imag} */,
  {32'h3ee8a054, 32'h00000000} /* (17, 21, 11) {real, imag} */,
  {32'h3de66b06, 32'h00000000} /* (17, 21, 10) {real, imag} */,
  {32'hbe663698, 32'h00000000} /* (17, 21, 9) {real, imag} */,
  {32'hbeb56654, 32'h00000000} /* (17, 21, 8) {real, imag} */,
  {32'hbe0b60de, 32'h00000000} /* (17, 21, 7) {real, imag} */,
  {32'h3cbee85a, 32'h00000000} /* (17, 21, 6) {real, imag} */,
  {32'h3e88f1e0, 32'h00000000} /* (17, 21, 5) {real, imag} */,
  {32'hbe44faa1, 32'h00000000} /* (17, 21, 4) {real, imag} */,
  {32'hbea1416f, 32'h00000000} /* (17, 21, 3) {real, imag} */,
  {32'hbe917a97, 32'h00000000} /* (17, 21, 2) {real, imag} */,
  {32'hbecbedd3, 32'h00000000} /* (17, 21, 1) {real, imag} */,
  {32'hbe8b719e, 32'h00000000} /* (17, 21, 0) {real, imag} */,
  {32'h3eee131e, 32'h00000000} /* (17, 20, 31) {real, imag} */,
  {32'h3f17b2c3, 32'h00000000} /* (17, 20, 30) {real, imag} */,
  {32'hbdc3482d, 32'h00000000} /* (17, 20, 29) {real, imag} */,
  {32'h3d52c8c9, 32'h00000000} /* (17, 20, 28) {real, imag} */,
  {32'hbde4815f, 32'h00000000} /* (17, 20, 27) {real, imag} */,
  {32'hbc6a7d9f, 32'h00000000} /* (17, 20, 26) {real, imag} */,
  {32'h3ebc0500, 32'h00000000} /* (17, 20, 25) {real, imag} */,
  {32'h3f2404ab, 32'h00000000} /* (17, 20, 24) {real, imag} */,
  {32'h3ee9d4e3, 32'h00000000} /* (17, 20, 23) {real, imag} */,
  {32'h3ef50679, 32'h00000000} /* (17, 20, 22) {real, imag} */,
  {32'h3e26067b, 32'h00000000} /* (17, 20, 21) {real, imag} */,
  {32'hbebdcb76, 32'h00000000} /* (17, 20, 20) {real, imag} */,
  {32'h3e667146, 32'h00000000} /* (17, 20, 19) {real, imag} */,
  {32'h3d427c38, 32'h00000000} /* (17, 20, 18) {real, imag} */,
  {32'hbe44f862, 32'h00000000} /* (17, 20, 17) {real, imag} */,
  {32'hbf0e936d, 32'h00000000} /* (17, 20, 16) {real, imag} */,
  {32'hbe89a171, 32'h00000000} /* (17, 20, 15) {real, imag} */,
  {32'hbf23aa5c, 32'h00000000} /* (17, 20, 14) {real, imag} */,
  {32'hbf44d247, 32'h00000000} /* (17, 20, 13) {real, imag} */,
  {32'hbf4b7b42, 32'h00000000} /* (17, 20, 12) {real, imag} */,
  {32'hbeef61a5, 32'h00000000} /* (17, 20, 11) {real, imag} */,
  {32'h3ec1e2e3, 32'h00000000} /* (17, 20, 10) {real, imag} */,
  {32'h3f6e855e, 32'h00000000} /* (17, 20, 9) {real, imag} */,
  {32'h3f550006, 32'h00000000} /* (17, 20, 8) {real, imag} */,
  {32'h3f372323, 32'h00000000} /* (17, 20, 7) {real, imag} */,
  {32'h3f7796c0, 32'h00000000} /* (17, 20, 6) {real, imag} */,
  {32'h3f848334, 32'h00000000} /* (17, 20, 5) {real, imag} */,
  {32'h3f00dbf9, 32'h00000000} /* (17, 20, 4) {real, imag} */,
  {32'h3ebe2d73, 32'h00000000} /* (17, 20, 3) {real, imag} */,
  {32'h3eeaef96, 32'h00000000} /* (17, 20, 2) {real, imag} */,
  {32'h3edacb38, 32'h00000000} /* (17, 20, 1) {real, imag} */,
  {32'h3ea43fc6, 32'h00000000} /* (17, 20, 0) {real, imag} */,
  {32'h3e7a317a, 32'h00000000} /* (17, 19, 31) {real, imag} */,
  {32'h3f2ae950, 32'h00000000} /* (17, 19, 30) {real, imag} */,
  {32'h3f1f5dd6, 32'h00000000} /* (17, 19, 29) {real, imag} */,
  {32'h3ea02ab9, 32'h00000000} /* (17, 19, 28) {real, imag} */,
  {32'h3ed73e5d, 32'h00000000} /* (17, 19, 27) {real, imag} */,
  {32'h3ef1e914, 32'h00000000} /* (17, 19, 26) {real, imag} */,
  {32'h3f4fc340, 32'h00000000} /* (17, 19, 25) {real, imag} */,
  {32'h3f8f34f1, 32'h00000000} /* (17, 19, 24) {real, imag} */,
  {32'h3fa645cc, 32'h00000000} /* (17, 19, 23) {real, imag} */,
  {32'h3f7a6f0a, 32'h00000000} /* (17, 19, 22) {real, imag} */,
  {32'h3eeae8c6, 32'h00000000} /* (17, 19, 21) {real, imag} */,
  {32'hbef1930c, 32'h00000000} /* (17, 19, 20) {real, imag} */,
  {32'hbf300eef, 32'h00000000} /* (17, 19, 19) {real, imag} */,
  {32'hbeda781a, 32'h00000000} /* (17, 19, 18) {real, imag} */,
  {32'hbec52138, 32'h00000000} /* (17, 19, 17) {real, imag} */,
  {32'hbf3da12c, 32'h00000000} /* (17, 19, 16) {real, imag} */,
  {32'hbf882f39, 32'h00000000} /* (17, 19, 15) {real, imag} */,
  {32'hbf6b7ab1, 32'h00000000} /* (17, 19, 14) {real, imag} */,
  {32'hbf0a8111, 32'h00000000} /* (17, 19, 13) {real, imag} */,
  {32'hbf22e4cc, 32'h00000000} /* (17, 19, 12) {real, imag} */,
  {32'hbf849a04, 32'h00000000} /* (17, 19, 11) {real, imag} */,
  {32'hbdb54c01, 32'h00000000} /* (17, 19, 10) {real, imag} */,
  {32'h3f6b5dac, 32'h00000000} /* (17, 19, 9) {real, imag} */,
  {32'h3f787851, 32'h00000000} /* (17, 19, 8) {real, imag} */,
  {32'h3f089657, 32'h00000000} /* (17, 19, 7) {real, imag} */,
  {32'h3f05c35a, 32'h00000000} /* (17, 19, 6) {real, imag} */,
  {32'h3f5a50a5, 32'h00000000} /* (17, 19, 5) {real, imag} */,
  {32'h3f7a7d51, 32'h00000000} /* (17, 19, 4) {real, imag} */,
  {32'h3f4b05c5, 32'h00000000} /* (17, 19, 3) {real, imag} */,
  {32'h3f8b9026, 32'h00000000} /* (17, 19, 2) {real, imag} */,
  {32'h3fa7abfd, 32'h00000000} /* (17, 19, 1) {real, imag} */,
  {32'h3f394520, 32'h00000000} /* (17, 19, 0) {real, imag} */,
  {32'h3ef0857b, 32'h00000000} /* (17, 18, 31) {real, imag} */,
  {32'h3f6c8b72, 32'h00000000} /* (17, 18, 30) {real, imag} */,
  {32'h3fa45903, 32'h00000000} /* (17, 18, 29) {real, imag} */,
  {32'h3f71a758, 32'h00000000} /* (17, 18, 28) {real, imag} */,
  {32'h3f40b057, 32'h00000000} /* (17, 18, 27) {real, imag} */,
  {32'h3f0841a6, 32'h00000000} /* (17, 18, 26) {real, imag} */,
  {32'h3f49570a, 32'h00000000} /* (17, 18, 25) {real, imag} */,
  {32'h3f942cff, 32'h00000000} /* (17, 18, 24) {real, imag} */,
  {32'h3facd3ec, 32'h00000000} /* (17, 18, 23) {real, imag} */,
  {32'h3f41e3dc, 32'h00000000} /* (17, 18, 22) {real, imag} */,
  {32'h3e8addc4, 32'h00000000} /* (17, 18, 21) {real, imag} */,
  {32'hbf102a14, 32'h00000000} /* (17, 18, 20) {real, imag} */,
  {32'hbf9e01d3, 32'h00000000} /* (17, 18, 19) {real, imag} */,
  {32'hbf6cc83c, 32'h00000000} /* (17, 18, 18) {real, imag} */,
  {32'hbf51ad31, 32'h00000000} /* (17, 18, 17) {real, imag} */,
  {32'hbf2bf201, 32'h00000000} /* (17, 18, 16) {real, imag} */,
  {32'hbf41fc23, 32'h00000000} /* (17, 18, 15) {real, imag} */,
  {32'hbf06733a, 32'h00000000} /* (17, 18, 14) {real, imag} */,
  {32'hbee8f6b9, 32'h00000000} /* (17, 18, 13) {real, imag} */,
  {32'hbec7acdd, 32'h00000000} /* (17, 18, 12) {real, imag} */,
  {32'hbf7e9981, 32'h00000000} /* (17, 18, 11) {real, imag} */,
  {32'h3f1c8752, 32'h00000000} /* (17, 18, 10) {real, imag} */,
  {32'h3fe80c9f, 32'h00000000} /* (17, 18, 9) {real, imag} */,
  {32'h3fb1709c, 32'h00000000} /* (17, 18, 8) {real, imag} */,
  {32'h3f2c90bd, 32'h00000000} /* (17, 18, 7) {real, imag} */,
  {32'h3f045abe, 32'h00000000} /* (17, 18, 6) {real, imag} */,
  {32'h3f0faad3, 32'h00000000} /* (17, 18, 5) {real, imag} */,
  {32'h3f85b991, 32'h00000000} /* (17, 18, 4) {real, imag} */,
  {32'h3f6fdef9, 32'h00000000} /* (17, 18, 3) {real, imag} */,
  {32'h3fb2c9c7, 32'h00000000} /* (17, 18, 2) {real, imag} */,
  {32'h3fbbd776, 32'h00000000} /* (17, 18, 1) {real, imag} */,
  {32'h3f4d92d0, 32'h00000000} /* (17, 18, 0) {real, imag} */,
  {32'h3f201098, 32'h00000000} /* (17, 17, 31) {real, imag} */,
  {32'h3f94c9e1, 32'h00000000} /* (17, 17, 30) {real, imag} */,
  {32'h3f975bfb, 32'h00000000} /* (17, 17, 29) {real, imag} */,
  {32'h3f8046ba, 32'h00000000} /* (17, 17, 28) {real, imag} */,
  {32'h3f2b6e1f, 32'h00000000} /* (17, 17, 27) {real, imag} */,
  {32'h3f12553d, 32'h00000000} /* (17, 17, 26) {real, imag} */,
  {32'h3f4606eb, 32'h00000000} /* (17, 17, 25) {real, imag} */,
  {32'h3faaf0c3, 32'h00000000} /* (17, 17, 24) {real, imag} */,
  {32'h3faed558, 32'h00000000} /* (17, 17, 23) {real, imag} */,
  {32'h3f6e5d23, 32'h00000000} /* (17, 17, 22) {real, imag} */,
  {32'h3ee05258, 32'h00000000} /* (17, 17, 21) {real, imag} */,
  {32'hbf0369e7, 32'h00000000} /* (17, 17, 20) {real, imag} */,
  {32'hbf893763, 32'h00000000} /* (17, 17, 19) {real, imag} */,
  {32'hbf659c67, 32'h00000000} /* (17, 17, 18) {real, imag} */,
  {32'hbf8ace75, 32'h00000000} /* (17, 17, 17) {real, imag} */,
  {32'hbf7aa0fd, 32'h00000000} /* (17, 17, 16) {real, imag} */,
  {32'hbf1ee4ae, 32'h00000000} /* (17, 17, 15) {real, imag} */,
  {32'hbf106cbc, 32'h00000000} /* (17, 17, 14) {real, imag} */,
  {32'hbf3cf0d5, 32'h00000000} /* (17, 17, 13) {real, imag} */,
  {32'hbf53cc9f, 32'h00000000} /* (17, 17, 12) {real, imag} */,
  {32'hbee5f63c, 32'h00000000} /* (17, 17, 11) {real, imag} */,
  {32'h3fd1fc82, 32'h00000000} /* (17, 17, 10) {real, imag} */,
  {32'h4005d940, 32'h00000000} /* (17, 17, 9) {real, imag} */,
  {32'h3fe97fb4, 32'h00000000} /* (17, 17, 8) {real, imag} */,
  {32'h3f844a66, 32'h00000000} /* (17, 17, 7) {real, imag} */,
  {32'h3ec2407f, 32'h00000000} /* (17, 17, 6) {real, imag} */,
  {32'h3f2bb042, 32'h00000000} /* (17, 17, 5) {real, imag} */,
  {32'h3f5d0f16, 32'h00000000} /* (17, 17, 4) {real, imag} */,
  {32'h3f509652, 32'h00000000} /* (17, 17, 3) {real, imag} */,
  {32'h3f6956b1, 32'h00000000} /* (17, 17, 2) {real, imag} */,
  {32'h3f579a13, 32'h00000000} /* (17, 17, 1) {real, imag} */,
  {32'h3f30677d, 32'h00000000} /* (17, 17, 0) {real, imag} */,
  {32'h3eab4b11, 32'h00000000} /* (17, 16, 31) {real, imag} */,
  {32'h3f599af4, 32'h00000000} /* (17, 16, 30) {real, imag} */,
  {32'h3f907e90, 32'h00000000} /* (17, 16, 29) {real, imag} */,
  {32'h3f5c766a, 32'h00000000} /* (17, 16, 28) {real, imag} */,
  {32'h3f6a0195, 32'h00000000} /* (17, 16, 27) {real, imag} */,
  {32'h3f59d0b4, 32'h00000000} /* (17, 16, 26) {real, imag} */,
  {32'h3f3374fd, 32'h00000000} /* (17, 16, 25) {real, imag} */,
  {32'h3f88b824, 32'h00000000} /* (17, 16, 24) {real, imag} */,
  {32'h3f956774, 32'h00000000} /* (17, 16, 23) {real, imag} */,
  {32'h3f5f91cf, 32'h00000000} /* (17, 16, 22) {real, imag} */,
  {32'h3efc7908, 32'h00000000} /* (17, 16, 21) {real, imag} */,
  {32'hbf0e1632, 32'h00000000} /* (17, 16, 20) {real, imag} */,
  {32'hbfb1a9dc, 32'h00000000} /* (17, 16, 19) {real, imag} */,
  {32'hbf878a71, 32'h00000000} /* (17, 16, 18) {real, imag} */,
  {32'hbf95315f, 32'h00000000} /* (17, 16, 17) {real, imag} */,
  {32'hbf806198, 32'h00000000} /* (17, 16, 16) {real, imag} */,
  {32'hbf626c68, 32'h00000000} /* (17, 16, 15) {real, imag} */,
  {32'hbf599cd2, 32'h00000000} /* (17, 16, 14) {real, imag} */,
  {32'hbfd89b7c, 32'h00000000} /* (17, 16, 13) {real, imag} */,
  {32'hbfddcfcb, 32'h00000000} /* (17, 16, 12) {real, imag} */,
  {32'hbf251306, 32'h00000000} /* (17, 16, 11) {real, imag} */,
  {32'h3f96b9b6, 32'h00000000} /* (17, 16, 10) {real, imag} */,
  {32'h3fe47be8, 32'h00000000} /* (17, 16, 9) {real, imag} */,
  {32'h3fbe2070, 32'h00000000} /* (17, 16, 8) {real, imag} */,
  {32'h3f6e6bd4, 32'h00000000} /* (17, 16, 7) {real, imag} */,
  {32'h3ecc3f6e, 32'h00000000} /* (17, 16, 6) {real, imag} */,
  {32'h3f1b0dfc, 32'h00000000} /* (17, 16, 5) {real, imag} */,
  {32'h3f0f7fa7, 32'h00000000} /* (17, 16, 4) {real, imag} */,
  {32'h3f231fef, 32'h00000000} /* (17, 16, 3) {real, imag} */,
  {32'h3f257907, 32'h00000000} /* (17, 16, 2) {real, imag} */,
  {32'h3f4fafe1, 32'h00000000} /* (17, 16, 1) {real, imag} */,
  {32'h3f035724, 32'h00000000} /* (17, 16, 0) {real, imag} */,
  {32'h3e21a601, 32'h00000000} /* (17, 15, 31) {real, imag} */,
  {32'h3f33823c, 32'h00000000} /* (17, 15, 30) {real, imag} */,
  {32'h3f8345e7, 32'h00000000} /* (17, 15, 29) {real, imag} */,
  {32'h3f0dba1c, 32'h00000000} /* (17, 15, 28) {real, imag} */,
  {32'h3f83d91f, 32'h00000000} /* (17, 15, 27) {real, imag} */,
  {32'h3f831914, 32'h00000000} /* (17, 15, 26) {real, imag} */,
  {32'h3f04d671, 32'h00000000} /* (17, 15, 25) {real, imag} */,
  {32'h3f05ad1d, 32'h00000000} /* (17, 15, 24) {real, imag} */,
  {32'h3f303cdb, 32'h00000000} /* (17, 15, 23) {real, imag} */,
  {32'h3f6981c9, 32'h00000000} /* (17, 15, 22) {real, imag} */,
  {32'h3f42f3b8, 32'h00000000} /* (17, 15, 21) {real, imag} */,
  {32'hbe81df2e, 32'h00000000} /* (17, 15, 20) {real, imag} */,
  {32'hbf6ae130, 32'h00000000} /* (17, 15, 19) {real, imag} */,
  {32'hbf86f046, 32'h00000000} /* (17, 15, 18) {real, imag} */,
  {32'hbf9458d4, 32'h00000000} /* (17, 15, 17) {real, imag} */,
  {32'hbf4575ce, 32'h00000000} /* (17, 15, 16) {real, imag} */,
  {32'hbf17cc4e, 32'h00000000} /* (17, 15, 15) {real, imag} */,
  {32'hbf305586, 32'h00000000} /* (17, 15, 14) {real, imag} */,
  {32'hbf937a86, 32'h00000000} /* (17, 15, 13) {real, imag} */,
  {32'hbfcce39d, 32'h00000000} /* (17, 15, 12) {real, imag} */,
  {32'hbf817c7a, 32'h00000000} /* (17, 15, 11) {real, imag} */,
  {32'h3fa387b1, 32'h00000000} /* (17, 15, 10) {real, imag} */,
  {32'h3ffeb8dd, 32'h00000000} /* (17, 15, 9) {real, imag} */,
  {32'h3f946612, 32'h00000000} /* (17, 15, 8) {real, imag} */,
  {32'h3f3c5d53, 32'h00000000} /* (17, 15, 7) {real, imag} */,
  {32'h3f1ad86b, 32'h00000000} /* (17, 15, 6) {real, imag} */,
  {32'h3f11bbb7, 32'h00000000} /* (17, 15, 5) {real, imag} */,
  {32'h3f868143, 32'h00000000} /* (17, 15, 4) {real, imag} */,
  {32'h3fa096ad, 32'h00000000} /* (17, 15, 3) {real, imag} */,
  {32'h3f8aff0f, 32'h00000000} /* (17, 15, 2) {real, imag} */,
  {32'h3f585d58, 32'h00000000} /* (17, 15, 1) {real, imag} */,
  {32'h3edd1fff, 32'h00000000} /* (17, 15, 0) {real, imag} */,
  {32'h3dce3a6f, 32'h00000000} /* (17, 14, 31) {real, imag} */,
  {32'h3f061ebd, 32'h00000000} /* (17, 14, 30) {real, imag} */,
  {32'h3fb6e751, 32'h00000000} /* (17, 14, 29) {real, imag} */,
  {32'h3f765f72, 32'h00000000} /* (17, 14, 28) {real, imag} */,
  {32'h3f5b5149, 32'h00000000} /* (17, 14, 27) {real, imag} */,
  {32'h3f33ac0a, 32'h00000000} /* (17, 14, 26) {real, imag} */,
  {32'h3ec8c651, 32'h00000000} /* (17, 14, 25) {real, imag} */,
  {32'h3e779701, 32'h00000000} /* (17, 14, 24) {real, imag} */,
  {32'h3f0c428b, 32'h00000000} /* (17, 14, 23) {real, imag} */,
  {32'h3fa4c0ad, 32'h00000000} /* (17, 14, 22) {real, imag} */,
  {32'h3f4b3b72, 32'h00000000} /* (17, 14, 21) {real, imag} */,
  {32'hbec9be2e, 32'h00000000} /* (17, 14, 20) {real, imag} */,
  {32'hbfd5be65, 32'h00000000} /* (17, 14, 19) {real, imag} */,
  {32'hbf9cd51e, 32'h00000000} /* (17, 14, 18) {real, imag} */,
  {32'hbf07797d, 32'h00000000} /* (17, 14, 17) {real, imag} */,
  {32'hbeec6d60, 32'h00000000} /* (17, 14, 16) {real, imag} */,
  {32'hbf052f51, 32'h00000000} /* (17, 14, 15) {real, imag} */,
  {32'hbf957871, 32'h00000000} /* (17, 14, 14) {real, imag} */,
  {32'hbf747f3b, 32'h00000000} /* (17, 14, 13) {real, imag} */,
  {32'hbf75bb32, 32'h00000000} /* (17, 14, 12) {real, imag} */,
  {32'hbeaf2c3f, 32'h00000000} /* (17, 14, 11) {real, imag} */,
  {32'h3f7a8842, 32'h00000000} /* (17, 14, 10) {real, imag} */,
  {32'h3fa32fc5, 32'h00000000} /* (17, 14, 9) {real, imag} */,
  {32'h3f4a9b74, 32'h00000000} /* (17, 14, 8) {real, imag} */,
  {32'h3f1ec596, 32'h00000000} /* (17, 14, 7) {real, imag} */,
  {32'h3ec97b5b, 32'h00000000} /* (17, 14, 6) {real, imag} */,
  {32'h3e05c24d, 32'h00000000} /* (17, 14, 5) {real, imag} */,
  {32'h3f618370, 32'h00000000} /* (17, 14, 4) {real, imag} */,
  {32'h3f9b6c2e, 32'h00000000} /* (17, 14, 3) {real, imag} */,
  {32'h3fabffd3, 32'h00000000} /* (17, 14, 2) {real, imag} */,
  {32'h3f7ae75e, 32'h00000000} /* (17, 14, 1) {real, imag} */,
  {32'h3ebe3050, 32'h00000000} /* (17, 14, 0) {real, imag} */,
  {32'h3e940671, 32'h00000000} /* (17, 13, 31) {real, imag} */,
  {32'h3f1ecef2, 32'h00000000} /* (17, 13, 30) {real, imag} */,
  {32'h3fa5696d, 32'h00000000} /* (17, 13, 29) {real, imag} */,
  {32'h3f82f91b, 32'h00000000} /* (17, 13, 28) {real, imag} */,
  {32'h3ef3068b, 32'h00000000} /* (17, 13, 27) {real, imag} */,
  {32'h3f3d4fda, 32'h00000000} /* (17, 13, 26) {real, imag} */,
  {32'h3f594998, 32'h00000000} /* (17, 13, 25) {real, imag} */,
  {32'h3ee7a15e, 32'h00000000} /* (17, 13, 24) {real, imag} */,
  {32'h3ed07d13, 32'h00000000} /* (17, 13, 23) {real, imag} */,
  {32'h3f918e86, 32'h00000000} /* (17, 13, 22) {real, imag} */,
  {32'h3f466d77, 32'h00000000} /* (17, 13, 21) {real, imag} */,
  {32'h3c2cc72f, 32'h00000000} /* (17, 13, 20) {real, imag} */,
  {32'hbf877ecb, 32'h00000000} /* (17, 13, 19) {real, imag} */,
  {32'hbf52e266, 32'h00000000} /* (17, 13, 18) {real, imag} */,
  {32'hbf35970c, 32'h00000000} /* (17, 13, 17) {real, imag} */,
  {32'hbf46c722, 32'h00000000} /* (17, 13, 16) {real, imag} */,
  {32'hbf4fcbdb, 32'h00000000} /* (17, 13, 15) {real, imag} */,
  {32'hbf8f6690, 32'h00000000} /* (17, 13, 14) {real, imag} */,
  {32'hbf22478d, 32'h00000000} /* (17, 13, 13) {real, imag} */,
  {32'hbea22b80, 32'h00000000} /* (17, 13, 12) {real, imag} */,
  {32'h3d3d42e8, 32'h00000000} /* (17, 13, 11) {real, imag} */,
  {32'h3f7a5223, 32'h00000000} /* (17, 13, 10) {real, imag} */,
  {32'h3fa7b537, 32'h00000000} /* (17, 13, 9) {real, imag} */,
  {32'h3fc5f955, 32'h00000000} /* (17, 13, 8) {real, imag} */,
  {32'h3f883b94, 32'h00000000} /* (17, 13, 7) {real, imag} */,
  {32'h3edf2b2c, 32'h00000000} /* (17, 13, 6) {real, imag} */,
  {32'h3eadf8ba, 32'h00000000} /* (17, 13, 5) {real, imag} */,
  {32'h3f5956d3, 32'h00000000} /* (17, 13, 4) {real, imag} */,
  {32'h3faa43d6, 32'h00000000} /* (17, 13, 3) {real, imag} */,
  {32'h3fa880c7, 32'h00000000} /* (17, 13, 2) {real, imag} */,
  {32'h3f5458b7, 32'h00000000} /* (17, 13, 1) {real, imag} */,
  {32'h3ef4f42d, 32'h00000000} /* (17, 13, 0) {real, imag} */,
  {32'h3f49f661, 32'h00000000} /* (17, 12, 31) {real, imag} */,
  {32'h3f829c9d, 32'h00000000} /* (17, 12, 30) {real, imag} */,
  {32'h3f94aa1e, 32'h00000000} /* (17, 12, 29) {real, imag} */,
  {32'h3f30b950, 32'h00000000} /* (17, 12, 28) {real, imag} */,
  {32'h3f00d8ef, 32'h00000000} /* (17, 12, 27) {real, imag} */,
  {32'h3f7ef686, 32'h00000000} /* (17, 12, 26) {real, imag} */,
  {32'h3fba90d2, 32'h00000000} /* (17, 12, 25) {real, imag} */,
  {32'h3f8be4db, 32'h00000000} /* (17, 12, 24) {real, imag} */,
  {32'h3f7a8507, 32'h00000000} /* (17, 12, 23) {real, imag} */,
  {32'h3fc0db3d, 32'h00000000} /* (17, 12, 22) {real, imag} */,
  {32'h3f6c2fd4, 32'h00000000} /* (17, 12, 21) {real, imag} */,
  {32'hbebfb745, 32'h00000000} /* (17, 12, 20) {real, imag} */,
  {32'hbfa7f0f8, 32'h00000000} /* (17, 12, 19) {real, imag} */,
  {32'hbf2de2d4, 32'h00000000} /* (17, 12, 18) {real, imag} */,
  {32'hbf2d243b, 32'h00000000} /* (17, 12, 17) {real, imag} */,
  {32'hbfbe405c, 32'h00000000} /* (17, 12, 16) {real, imag} */,
  {32'hbfc91ecc, 32'h00000000} /* (17, 12, 15) {real, imag} */,
  {32'hbf791054, 32'h00000000} /* (17, 12, 14) {real, imag} */,
  {32'hbec4e441, 32'h00000000} /* (17, 12, 13) {real, imag} */,
  {32'hbf145485, 32'h00000000} /* (17, 12, 12) {real, imag} */,
  {32'hbe9f1bd3, 32'h00000000} /* (17, 12, 11) {real, imag} */,
  {32'h3f3c124e, 32'h00000000} /* (17, 12, 10) {real, imag} */,
  {32'h3f9d021b, 32'h00000000} /* (17, 12, 9) {real, imag} */,
  {32'h3fa7b294, 32'h00000000} /* (17, 12, 8) {real, imag} */,
  {32'h3f8fb83b, 32'h00000000} /* (17, 12, 7) {real, imag} */,
  {32'h3f337f9f, 32'h00000000} /* (17, 12, 6) {real, imag} */,
  {32'h3f288a13, 32'h00000000} /* (17, 12, 5) {real, imag} */,
  {32'h3f530a21, 32'h00000000} /* (17, 12, 4) {real, imag} */,
  {32'h3fb20a62, 32'h00000000} /* (17, 12, 3) {real, imag} */,
  {32'h3faa1e2f, 32'h00000000} /* (17, 12, 2) {real, imag} */,
  {32'h3f945ff7, 32'h00000000} /* (17, 12, 1) {real, imag} */,
  {32'h3f37a123, 32'h00000000} /* (17, 12, 0) {real, imag} */,
  {32'h3ecd3a85, 32'h00000000} /* (17, 11, 31) {real, imag} */,
  {32'h3f4a5b7a, 32'h00000000} /* (17, 11, 30) {real, imag} */,
  {32'h3f5c4f60, 32'h00000000} /* (17, 11, 29) {real, imag} */,
  {32'h3f0a4b57, 32'h00000000} /* (17, 11, 28) {real, imag} */,
  {32'h3e7540bc, 32'h00000000} /* (17, 11, 27) {real, imag} */,
  {32'h3eb4869a, 32'h00000000} /* (17, 11, 26) {real, imag} */,
  {32'h3f6a02dc, 32'h00000000} /* (17, 11, 25) {real, imag} */,
  {32'h3f2169fb, 32'h00000000} /* (17, 11, 24) {real, imag} */,
  {32'h3f5efc3e, 32'h00000000} /* (17, 11, 23) {real, imag} */,
  {32'h3f740100, 32'h00000000} /* (17, 11, 22) {real, imag} */,
  {32'h3f87ec36, 32'h00000000} /* (17, 11, 21) {real, imag} */,
  {32'hbdf7ef1a, 32'h00000000} /* (17, 11, 20) {real, imag} */,
  {32'hbf89a94e, 32'h00000000} /* (17, 11, 19) {real, imag} */,
  {32'hbf578d70, 32'h00000000} /* (17, 11, 18) {real, imag} */,
  {32'hbf3089fe, 32'h00000000} /* (17, 11, 17) {real, imag} */,
  {32'hbfc36c13, 32'h00000000} /* (17, 11, 16) {real, imag} */,
  {32'hbfa00510, 32'h00000000} /* (17, 11, 15) {real, imag} */,
  {32'hbee34ccd, 32'h00000000} /* (17, 11, 14) {real, imag} */,
  {32'hbe88ae08, 32'h00000000} /* (17, 11, 13) {real, imag} */,
  {32'hbf1a62cb, 32'h00000000} /* (17, 11, 12) {real, imag} */,
  {32'hbee8d8d0, 32'h00000000} /* (17, 11, 11) {real, imag} */,
  {32'h3ea45a24, 32'h00000000} /* (17, 11, 10) {real, imag} */,
  {32'h3f8bcfbe, 32'h00000000} /* (17, 11, 9) {real, imag} */,
  {32'h3f8975a1, 32'h00000000} /* (17, 11, 8) {real, imag} */,
  {32'h3f23b794, 32'h00000000} /* (17, 11, 7) {real, imag} */,
  {32'h3f467da3, 32'h00000000} /* (17, 11, 6) {real, imag} */,
  {32'h3fb1d167, 32'h00000000} /* (17, 11, 5) {real, imag} */,
  {32'h3f57ac63, 32'h00000000} /* (17, 11, 4) {real, imag} */,
  {32'h3f37b3e6, 32'h00000000} /* (17, 11, 3) {real, imag} */,
  {32'h3f6a23e6, 32'h00000000} /* (17, 11, 2) {real, imag} */,
  {32'h3fb4dfa6, 32'h00000000} /* (17, 11, 1) {real, imag} */,
  {32'h3f373557, 32'h00000000} /* (17, 11, 0) {real, imag} */,
  {32'hbf011690, 32'h00000000} /* (17, 10, 31) {real, imag} */,
  {32'hbf26c74d, 32'h00000000} /* (17, 10, 30) {real, imag} */,
  {32'hbf3196ba, 32'h00000000} /* (17, 10, 29) {real, imag} */,
  {32'hbe9d4a3f, 32'h00000000} /* (17, 10, 28) {real, imag} */,
  {32'hbf15845f, 32'h00000000} /* (17, 10, 27) {real, imag} */,
  {32'hbf4358db, 32'h00000000} /* (17, 10, 26) {real, imag} */,
  {32'hbea5fc13, 32'h00000000} /* (17, 10, 25) {real, imag} */,
  {32'hbe65e786, 32'h00000000} /* (17, 10, 24) {real, imag} */,
  {32'h3d4b31fa, 32'h00000000} /* (17, 10, 23) {real, imag} */,
  {32'hbe495e07, 32'h00000000} /* (17, 10, 22) {real, imag} */,
  {32'hbc98d3c5, 32'h00000000} /* (17, 10, 21) {real, imag} */,
  {32'h3f021e9c, 32'h00000000} /* (17, 10, 20) {real, imag} */,
  {32'hbccf6b32, 32'h00000000} /* (17, 10, 19) {real, imag} */,
  {32'hbe62b7b0, 32'h00000000} /* (17, 10, 18) {real, imag} */,
  {32'hbd2af78c, 32'h00000000} /* (17, 10, 17) {real, imag} */,
  {32'hbbfef678, 32'h00000000} /* (17, 10, 16) {real, imag} */,
  {32'h3f19b406, 32'h00000000} /* (17, 10, 15) {real, imag} */,
  {32'h3ef75110, 32'h00000000} /* (17, 10, 14) {real, imag} */,
  {32'h3f58840f, 32'h00000000} /* (17, 10, 13) {real, imag} */,
  {32'h3f56818d, 32'h00000000} /* (17, 10, 12) {real, imag} */,
  {32'h3ec08d5e, 32'h00000000} /* (17, 10, 11) {real, imag} */,
  {32'hbd5a9710, 32'h00000000} /* (17, 10, 10) {real, imag} */,
  {32'hbe3fb6af, 32'h00000000} /* (17, 10, 9) {real, imag} */,
  {32'hbe00ab79, 32'h00000000} /* (17, 10, 8) {real, imag} */,
  {32'hbf0faaa4, 32'h00000000} /* (17, 10, 7) {real, imag} */,
  {32'hbe987759, 32'h00000000} /* (17, 10, 6) {real, imag} */,
  {32'hbd9facc4, 32'h00000000} /* (17, 10, 5) {real, imag} */,
  {32'hbe842103, 32'h00000000} /* (17, 10, 4) {real, imag} */,
  {32'hbe8e7779, 32'h00000000} /* (17, 10, 3) {real, imag} */,
  {32'hbf368d1d, 32'h00000000} /* (17, 10, 2) {real, imag} */,
  {32'hbe9b01a8, 32'h00000000} /* (17, 10, 1) {real, imag} */,
  {32'hbed4fb1a, 32'h00000000} /* (17, 10, 0) {real, imag} */,
  {32'hbf355c0f, 32'h00000000} /* (17, 9, 31) {real, imag} */,
  {32'hbf941a43, 32'h00000000} /* (17, 9, 30) {real, imag} */,
  {32'hbf319bcd, 32'h00000000} /* (17, 9, 29) {real, imag} */,
  {32'hbf2c0361, 32'h00000000} /* (17, 9, 28) {real, imag} */,
  {32'hbf812313, 32'h00000000} /* (17, 9, 27) {real, imag} */,
  {32'hbf5afcb7, 32'h00000000} /* (17, 9, 26) {real, imag} */,
  {32'hbee48959, 32'h00000000} /* (17, 9, 25) {real, imag} */,
  {32'hbece65f2, 32'h00000000} /* (17, 9, 24) {real, imag} */,
  {32'hbe3aaf8a, 32'h00000000} /* (17, 9, 23) {real, imag} */,
  {32'hbf70b965, 32'h00000000} /* (17, 9, 22) {real, imag} */,
  {32'hbf2adc78, 32'h00000000} /* (17, 9, 21) {real, imag} */,
  {32'h3f0ff79a, 32'h00000000} /* (17, 9, 20) {real, imag} */,
  {32'h3f1557ae, 32'h00000000} /* (17, 9, 19) {real, imag} */,
  {32'h3f11e034, 32'h00000000} /* (17, 9, 18) {real, imag} */,
  {32'h3f53bc3d, 32'h00000000} /* (17, 9, 17) {real, imag} */,
  {32'h3fa183e2, 32'h00000000} /* (17, 9, 16) {real, imag} */,
  {32'h3fc77a1e, 32'h00000000} /* (17, 9, 15) {real, imag} */,
  {32'h3f9ea845, 32'h00000000} /* (17, 9, 14) {real, imag} */,
  {32'h3f6394fe, 32'h00000000} /* (17, 9, 13) {real, imag} */,
  {32'h3f250f91, 32'h00000000} /* (17, 9, 12) {real, imag} */,
  {32'h3e7ca864, 32'h00000000} /* (17, 9, 11) {real, imag} */,
  {32'hbeb9e02e, 32'h00000000} /* (17, 9, 10) {real, imag} */,
  {32'hbf404c19, 32'h00000000} /* (17, 9, 9) {real, imag} */,
  {32'hbf375df6, 32'h00000000} /* (17, 9, 8) {real, imag} */,
  {32'hbf5a2efd, 32'h00000000} /* (17, 9, 7) {real, imag} */,
  {32'hbf2b2997, 32'h00000000} /* (17, 9, 6) {real, imag} */,
  {32'hbfb1a398, 32'h00000000} /* (17, 9, 5) {real, imag} */,
  {32'hbf85b764, 32'h00000000} /* (17, 9, 4) {real, imag} */,
  {32'hbee27942, 32'h00000000} /* (17, 9, 3) {real, imag} */,
  {32'hbf36a098, 32'h00000000} /* (17, 9, 2) {real, imag} */,
  {32'hbf71c244, 32'h00000000} /* (17, 9, 1) {real, imag} */,
  {32'hbf4cc0ef, 32'h00000000} /* (17, 9, 0) {real, imag} */,
  {32'hbf6deddf, 32'h00000000} /* (17, 8, 31) {real, imag} */,
  {32'hbf8eebde, 32'h00000000} /* (17, 8, 30) {real, imag} */,
  {32'hbf2863da, 32'h00000000} /* (17, 8, 29) {real, imag} */,
  {32'hbf66988b, 32'h00000000} /* (17, 8, 28) {real, imag} */,
  {32'hbf883dac, 32'h00000000} /* (17, 8, 27) {real, imag} */,
  {32'hbf83b6fc, 32'h00000000} /* (17, 8, 26) {real, imag} */,
  {32'hbf244f70, 32'h00000000} /* (17, 8, 25) {real, imag} */,
  {32'hbe4629bd, 32'h00000000} /* (17, 8, 24) {real, imag} */,
  {32'hbf14a2ad, 32'h00000000} /* (17, 8, 23) {real, imag} */,
  {32'hbf1983ea, 32'h00000000} /* (17, 8, 22) {real, imag} */,
  {32'hbeb7279d, 32'h00000000} /* (17, 8, 21) {real, imag} */,
  {32'h3de7f5c7, 32'h00000000} /* (17, 8, 20) {real, imag} */,
  {32'h3ee1647f, 32'h00000000} /* (17, 8, 19) {real, imag} */,
  {32'h3f04cd55, 32'h00000000} /* (17, 8, 18) {real, imag} */,
  {32'h3f32a8d1, 32'h00000000} /* (17, 8, 17) {real, imag} */,
  {32'h3fdd7d02, 32'h00000000} /* (17, 8, 16) {real, imag} */,
  {32'h3f98c547, 32'h00000000} /* (17, 8, 15) {real, imag} */,
  {32'h3f73ac60, 32'h00000000} /* (17, 8, 14) {real, imag} */,
  {32'h3f65a78b, 32'h00000000} /* (17, 8, 13) {real, imag} */,
  {32'h3f834140, 32'h00000000} /* (17, 8, 12) {real, imag} */,
  {32'h3e2d9d5d, 32'h00000000} /* (17, 8, 11) {real, imag} */,
  {32'hbf297311, 32'h00000000} /* (17, 8, 10) {real, imag} */,
  {32'hbf7a1ade, 32'h00000000} /* (17, 8, 9) {real, imag} */,
  {32'hbf52e61e, 32'h00000000} /* (17, 8, 8) {real, imag} */,
  {32'hbecd2c54, 32'h00000000} /* (17, 8, 7) {real, imag} */,
  {32'hbf1d4c42, 32'h00000000} /* (17, 8, 6) {real, imag} */,
  {32'hbfda4854, 32'h00000000} /* (17, 8, 5) {real, imag} */,
  {32'hbfc06156, 32'h00000000} /* (17, 8, 4) {real, imag} */,
  {32'hbf429c0a, 32'h00000000} /* (17, 8, 3) {real, imag} */,
  {32'hbf772659, 32'h00000000} /* (17, 8, 2) {real, imag} */,
  {32'hbf8387a7, 32'h00000000} /* (17, 8, 1) {real, imag} */,
  {32'hbf5f0f23, 32'h00000000} /* (17, 8, 0) {real, imag} */,
  {32'hbf985963, 32'h00000000} /* (17, 7, 31) {real, imag} */,
  {32'hbfc95d94, 32'h00000000} /* (17, 7, 30) {real, imag} */,
  {32'hbf933886, 32'h00000000} /* (17, 7, 29) {real, imag} */,
  {32'hbf43367d, 32'h00000000} /* (17, 7, 28) {real, imag} */,
  {32'hbf67ba9b, 32'h00000000} /* (17, 7, 27) {real, imag} */,
  {32'hbf86b094, 32'h00000000} /* (17, 7, 26) {real, imag} */,
  {32'hbf85884e, 32'h00000000} /* (17, 7, 25) {real, imag} */,
  {32'hbf44b988, 32'h00000000} /* (17, 7, 24) {real, imag} */,
  {32'hbfa80bbf, 32'h00000000} /* (17, 7, 23) {real, imag} */,
  {32'hbf556a33, 32'h00000000} /* (17, 7, 22) {real, imag} */,
  {32'hbf3b284d, 32'h00000000} /* (17, 7, 21) {real, imag} */,
  {32'h3ce93b3e, 32'h00000000} /* (17, 7, 20) {real, imag} */,
  {32'h3f138de0, 32'h00000000} /* (17, 7, 19) {real, imag} */,
  {32'h3f8b93e1, 32'h00000000} /* (17, 7, 18) {real, imag} */,
  {32'h3f6742e1, 32'h00000000} /* (17, 7, 17) {real, imag} */,
  {32'h3f4ecf50, 32'h00000000} /* (17, 7, 16) {real, imag} */,
  {32'h3f06f85e, 32'h00000000} /* (17, 7, 15) {real, imag} */,
  {32'h3f2c6237, 32'h00000000} /* (17, 7, 14) {real, imag} */,
  {32'h3f6bf248, 32'h00000000} /* (17, 7, 13) {real, imag} */,
  {32'h3fba7c56, 32'h00000000} /* (17, 7, 12) {real, imag} */,
  {32'h3f86d233, 32'h00000000} /* (17, 7, 11) {real, imag} */,
  {32'hbf3ccd7c, 32'h00000000} /* (17, 7, 10) {real, imag} */,
  {32'hbfc16676, 32'h00000000} /* (17, 7, 9) {real, imag} */,
  {32'hbf902508, 32'h00000000} /* (17, 7, 8) {real, imag} */,
  {32'hbf0a80d4, 32'h00000000} /* (17, 7, 7) {real, imag} */,
  {32'hbfa08c62, 32'h00000000} /* (17, 7, 6) {real, imag} */,
  {32'hbfac4a0e, 32'h00000000} /* (17, 7, 5) {real, imag} */,
  {32'hbfaea061, 32'h00000000} /* (17, 7, 4) {real, imag} */,
  {32'hbf876aa7, 32'h00000000} /* (17, 7, 3) {real, imag} */,
  {32'hbf7dbb9f, 32'h00000000} /* (17, 7, 2) {real, imag} */,
  {32'hbf6812d1, 32'h00000000} /* (17, 7, 1) {real, imag} */,
  {32'hbef43b90, 32'h00000000} /* (17, 7, 0) {real, imag} */,
  {32'hbf3d9076, 32'h00000000} /* (17, 6, 31) {real, imag} */,
  {32'hbfc09b54, 32'h00000000} /* (17, 6, 30) {real, imag} */,
  {32'hbfc45b53, 32'h00000000} /* (17, 6, 29) {real, imag} */,
  {32'hbf492f45, 32'h00000000} /* (17, 6, 28) {real, imag} */,
  {32'hbecb6112, 32'h00000000} /* (17, 6, 27) {real, imag} */,
  {32'hbf3b9d75, 32'h00000000} /* (17, 6, 26) {real, imag} */,
  {32'hbfb73d77, 32'h00000000} /* (17, 6, 25) {real, imag} */,
  {32'hbfb71cd9, 32'h00000000} /* (17, 6, 24) {real, imag} */,
  {32'hbf7fd89e, 32'h00000000} /* (17, 6, 23) {real, imag} */,
  {32'hbf6b0897, 32'h00000000} /* (17, 6, 22) {real, imag} */,
  {32'hbf85d144, 32'h00000000} /* (17, 6, 21) {real, imag} */,
  {32'h3ecf4a16, 32'h00000000} /* (17, 6, 20) {real, imag} */,
  {32'h3f4a37ef, 32'h00000000} /* (17, 6, 19) {real, imag} */,
  {32'h3f59785a, 32'h00000000} /* (17, 6, 18) {real, imag} */,
  {32'h3f7384af, 32'h00000000} /* (17, 6, 17) {real, imag} */,
  {32'h3f5f3996, 32'h00000000} /* (17, 6, 16) {real, imag} */,
  {32'h3f6effc6, 32'h00000000} /* (17, 6, 15) {real, imag} */,
  {32'h3f5298e1, 32'h00000000} /* (17, 6, 14) {real, imag} */,
  {32'h3f4efb60, 32'h00000000} /* (17, 6, 13) {real, imag} */,
  {32'h3f653b84, 32'h00000000} /* (17, 6, 12) {real, imag} */,
  {32'h3f470712, 32'h00000000} /* (17, 6, 11) {real, imag} */,
  {32'hbee9c716, 32'h00000000} /* (17, 6, 10) {real, imag} */,
  {32'hbfd64c3a, 32'h00000000} /* (17, 6, 9) {real, imag} */,
  {32'hbf7939dc, 32'h00000000} /* (17, 6, 8) {real, imag} */,
  {32'hbf0b902b, 32'h00000000} /* (17, 6, 7) {real, imag} */,
  {32'hbf84aa8b, 32'h00000000} /* (17, 6, 6) {real, imag} */,
  {32'hbf52b4a9, 32'h00000000} /* (17, 6, 5) {real, imag} */,
  {32'hbfaa3a04, 32'h00000000} /* (17, 6, 4) {real, imag} */,
  {32'hbfa176cb, 32'h00000000} /* (17, 6, 3) {real, imag} */,
  {32'hbf8f7443, 32'h00000000} /* (17, 6, 2) {real, imag} */,
  {32'hbf59f17d, 32'h00000000} /* (17, 6, 1) {real, imag} */,
  {32'hbeb60d4e, 32'h00000000} /* (17, 6, 0) {real, imag} */,
  {32'hbf100076, 32'h00000000} /* (17, 5, 31) {real, imag} */,
  {32'hbf8eabf1, 32'h00000000} /* (17, 5, 30) {real, imag} */,
  {32'hbfc6dc3e, 32'h00000000} /* (17, 5, 29) {real, imag} */,
  {32'hbf89a664, 32'h00000000} /* (17, 5, 28) {real, imag} */,
  {32'hbf0bc37b, 32'h00000000} /* (17, 5, 27) {real, imag} */,
  {32'hbef5d1c6, 32'h00000000} /* (17, 5, 26) {real, imag} */,
  {32'hbf92383f, 32'h00000000} /* (17, 5, 25) {real, imag} */,
  {32'hbf76da8f, 32'h00000000} /* (17, 5, 24) {real, imag} */,
  {32'hbf223e7d, 32'h00000000} /* (17, 5, 23) {real, imag} */,
  {32'hbf6d82ff, 32'h00000000} /* (17, 5, 22) {real, imag} */,
  {32'hbfa2d904, 32'h00000000} /* (17, 5, 21) {real, imag} */,
  {32'hbf6e916b, 32'h00000000} /* (17, 5, 20) {real, imag} */,
  {32'hbf20f884, 32'h00000000} /* (17, 5, 19) {real, imag} */,
  {32'hbe2caf98, 32'h00000000} /* (17, 5, 18) {real, imag} */,
  {32'h3ddb16ce, 32'h00000000} /* (17, 5, 17) {real, imag} */,
  {32'h3e395c27, 32'h00000000} /* (17, 5, 16) {real, imag} */,
  {32'h3f01082a, 32'h00000000} /* (17, 5, 15) {real, imag} */,
  {32'h3f434cbe, 32'h00000000} /* (17, 5, 14) {real, imag} */,
  {32'h3f1b3d76, 32'h00000000} /* (17, 5, 13) {real, imag} */,
  {32'h3e889dd5, 32'h00000000} /* (17, 5, 12) {real, imag} */,
  {32'h3f11743e, 32'h00000000} /* (17, 5, 11) {real, imag} */,
  {32'h3e90f92c, 32'h00000000} /* (17, 5, 10) {real, imag} */,
  {32'hbe082b8b, 32'h00000000} /* (17, 5, 9) {real, imag} */,
  {32'h3e9db0ad, 32'h00000000} /* (17, 5, 8) {real, imag} */,
  {32'h3e879a0b, 32'h00000000} /* (17, 5, 7) {real, imag} */,
  {32'hbe58ca25, 32'h00000000} /* (17, 5, 6) {real, imag} */,
  {32'hbf2db156, 32'h00000000} /* (17, 5, 5) {real, imag} */,
  {32'hbfac4a77, 32'h00000000} /* (17, 5, 4) {real, imag} */,
  {32'hbf7bb84d, 32'h00000000} /* (17, 5, 3) {real, imag} */,
  {32'hbf7b558b, 32'h00000000} /* (17, 5, 2) {real, imag} */,
  {32'hbf23a84c, 32'h00000000} /* (17, 5, 1) {real, imag} */,
  {32'hbeedd683, 32'h00000000} /* (17, 5, 0) {real, imag} */,
  {32'hbec5e125, 32'h00000000} /* (17, 4, 31) {real, imag} */,
  {32'hbf99523c, 32'h00000000} /* (17, 4, 30) {real, imag} */,
  {32'hbfbdce3a, 32'h00000000} /* (17, 4, 29) {real, imag} */,
  {32'hbf63338d, 32'h00000000} /* (17, 4, 28) {real, imag} */,
  {32'hbf180081, 32'h00000000} /* (17, 4, 27) {real, imag} */,
  {32'hbea8502c, 32'h00000000} /* (17, 4, 26) {real, imag} */,
  {32'hbee6c2db, 32'h00000000} /* (17, 4, 25) {real, imag} */,
  {32'hbed12edf, 32'h00000000} /* (17, 4, 24) {real, imag} */,
  {32'hbf2c4ad5, 32'h00000000} /* (17, 4, 23) {real, imag} */,
  {32'hbf48fd43, 32'h00000000} /* (17, 4, 22) {real, imag} */,
  {32'hbfa0faaf, 32'h00000000} /* (17, 4, 21) {real, imag} */,
  {32'hbfaf5bf2, 32'h00000000} /* (17, 4, 20) {real, imag} */,
  {32'hbf6e0e94, 32'h00000000} /* (17, 4, 19) {real, imag} */,
  {32'hbf2549f2, 32'h00000000} /* (17, 4, 18) {real, imag} */,
  {32'hbf8c84b0, 32'h00000000} /* (17, 4, 17) {real, imag} */,
  {32'hbf0ffd57, 32'h00000000} /* (17, 4, 16) {real, imag} */,
  {32'h3ed14abc, 32'h00000000} /* (17, 4, 15) {real, imag} */,
  {32'h3f86f961, 32'h00000000} /* (17, 4, 14) {real, imag} */,
  {32'h3f2b8348, 32'h00000000} /* (17, 4, 13) {real, imag} */,
  {32'h3e98770e, 32'h00000000} /* (17, 4, 12) {real, imag} */,
  {32'h3f58590a, 32'h00000000} /* (17, 4, 11) {real, imag} */,
  {32'h3f387d64, 32'h00000000} /* (17, 4, 10) {real, imag} */,
  {32'h3f8daa50, 32'h00000000} /* (17, 4, 9) {real, imag} */,
  {32'h3fd5e2ab, 32'h00000000} /* (17, 4, 8) {real, imag} */,
  {32'h3f9329ae, 32'h00000000} /* (17, 4, 7) {real, imag} */,
  {32'h3f0a921e, 32'h00000000} /* (17, 4, 6) {real, imag} */,
  {32'hbf08d511, 32'h00000000} /* (17, 4, 5) {real, imag} */,
  {32'hbfd24cb0, 32'h00000000} /* (17, 4, 4) {real, imag} */,
  {32'hbf5031f7, 32'h00000000} /* (17, 4, 3) {real, imag} */,
  {32'hbecd4eda, 32'h00000000} /* (17, 4, 2) {real, imag} */,
  {32'hbeda3e0d, 32'h00000000} /* (17, 4, 1) {real, imag} */,
  {32'hbeb96e2a, 32'h00000000} /* (17, 4, 0) {real, imag} */,
  {32'hbe8b7d9f, 32'h00000000} /* (17, 3, 31) {real, imag} */,
  {32'hbfcc57d7, 32'h00000000} /* (17, 3, 30) {real, imag} */,
  {32'hbfc35354, 32'h00000000} /* (17, 3, 29) {real, imag} */,
  {32'hbf241e11, 32'h00000000} /* (17, 3, 28) {real, imag} */,
  {32'hbf4f0853, 32'h00000000} /* (17, 3, 27) {real, imag} */,
  {32'hbf31b630, 32'h00000000} /* (17, 3, 26) {real, imag} */,
  {32'hbf21c6ce, 32'h00000000} /* (17, 3, 25) {real, imag} */,
  {32'hbf226374, 32'h00000000} /* (17, 3, 24) {real, imag} */,
  {32'hbf3c23fa, 32'h00000000} /* (17, 3, 23) {real, imag} */,
  {32'hbf773561, 32'h00000000} /* (17, 3, 22) {real, imag} */,
  {32'hbf70aac0, 32'h00000000} /* (17, 3, 21) {real, imag} */,
  {32'hbf3078dc, 32'h00000000} /* (17, 3, 20) {real, imag} */,
  {32'hbf64f474, 32'h00000000} /* (17, 3, 19) {real, imag} */,
  {32'hc001c1f1, 32'h00000000} /* (17, 3, 18) {real, imag} */,
  {32'hbfae1de0, 32'h00000000} /* (17, 3, 17) {real, imag} */,
  {32'hbe6c12cf, 32'h00000000} /* (17, 3, 16) {real, imag} */,
  {32'h3fac1cc7, 32'h00000000} /* (17, 3, 15) {real, imag} */,
  {32'h3fd2e629, 32'h00000000} /* (17, 3, 14) {real, imag} */,
  {32'h3fb70d4a, 32'h00000000} /* (17, 3, 13) {real, imag} */,
  {32'h3f97953a, 32'h00000000} /* (17, 3, 12) {real, imag} */,
  {32'h3fd39dca, 32'h00000000} /* (17, 3, 11) {real, imag} */,
  {32'h3f9d4eac, 32'h00000000} /* (17, 3, 10) {real, imag} */,
  {32'h3fa8fc57, 32'h00000000} /* (17, 3, 9) {real, imag} */,
  {32'h3fd2b3d7, 32'h00000000} /* (17, 3, 8) {real, imag} */,
  {32'h3f45ce32, 32'h00000000} /* (17, 3, 7) {real, imag} */,
  {32'h3ed5cddd, 32'h00000000} /* (17, 3, 6) {real, imag} */,
  {32'hbf2be92b, 32'h00000000} /* (17, 3, 5) {real, imag} */,
  {32'hbfadcebd, 32'h00000000} /* (17, 3, 4) {real, imag} */,
  {32'hbf1522d0, 32'h00000000} /* (17, 3, 3) {real, imag} */,
  {32'hbeaba0d5, 32'h00000000} /* (17, 3, 2) {real, imag} */,
  {32'hbee32afd, 32'h00000000} /* (17, 3, 1) {real, imag} */,
  {32'hbe5452cd, 32'h00000000} /* (17, 3, 0) {real, imag} */,
  {32'hbe510cd3, 32'h00000000} /* (17, 2, 31) {real, imag} */,
  {32'hbf68f8f8, 32'h00000000} /* (17, 2, 30) {real, imag} */,
  {32'hbf729eb6, 32'h00000000} /* (17, 2, 29) {real, imag} */,
  {32'hbefc5a3f, 32'h00000000} /* (17, 2, 28) {real, imag} */,
  {32'hbf4ea8b5, 32'h00000000} /* (17, 2, 27) {real, imag} */,
  {32'hbfa5bef7, 32'h00000000} /* (17, 2, 26) {real, imag} */,
  {32'hbf701491, 32'h00000000} /* (17, 2, 25) {real, imag} */,
  {32'hbefb467f, 32'h00000000} /* (17, 2, 24) {real, imag} */,
  {32'hbedc690e, 32'h00000000} /* (17, 2, 23) {real, imag} */,
  {32'hbf0a5ebe, 32'h00000000} /* (17, 2, 22) {real, imag} */,
  {32'hbeefc586, 32'h00000000} /* (17, 2, 21) {real, imag} */,
  {32'hbec135bc, 32'h00000000} /* (17, 2, 20) {real, imag} */,
  {32'hbf94de03, 32'h00000000} /* (17, 2, 19) {real, imag} */,
  {32'hc04488e9, 32'h00000000} /* (17, 2, 18) {real, imag} */,
  {32'hc00512a7, 32'h00000000} /* (17, 2, 17) {real, imag} */,
  {32'hbe963fe9, 32'h00000000} /* (17, 2, 16) {real, imag} */,
  {32'h3f9749f5, 32'h00000000} /* (17, 2, 15) {real, imag} */,
  {32'h3fb81a66, 32'h00000000} /* (17, 2, 14) {real, imag} */,
  {32'h3fdffe4e, 32'h00000000} /* (17, 2, 13) {real, imag} */,
  {32'h3f9a1987, 32'h00000000} /* (17, 2, 12) {real, imag} */,
  {32'h3fc91fb2, 32'h00000000} /* (17, 2, 11) {real, imag} */,
  {32'h3f862058, 32'h00000000} /* (17, 2, 10) {real, imag} */,
  {32'h3f48d406, 32'h00000000} /* (17, 2, 9) {real, imag} */,
  {32'h3f825188, 32'h00000000} /* (17, 2, 8) {real, imag} */,
  {32'h3f16455d, 32'h00000000} /* (17, 2, 7) {real, imag} */,
  {32'h3e98e3a2, 32'h00000000} /* (17, 2, 6) {real, imag} */,
  {32'hbf20db46, 32'h00000000} /* (17, 2, 5) {real, imag} */,
  {32'hbf8d8c03, 32'h00000000} /* (17, 2, 4) {real, imag} */,
  {32'hbf18b84f, 32'h00000000} /* (17, 2, 3) {real, imag} */,
  {32'hbf3ff6d1, 32'h00000000} /* (17, 2, 2) {real, imag} */,
  {32'hbf43b1f0, 32'h00000000} /* (17, 2, 1) {real, imag} */,
  {32'hbe94da72, 32'h00000000} /* (17, 2, 0) {real, imag} */,
  {32'hbe885e15, 32'h00000000} /* (17, 1, 31) {real, imag} */,
  {32'hbf1ba183, 32'h00000000} /* (17, 1, 30) {real, imag} */,
  {32'hbf67b4af, 32'h00000000} /* (17, 1, 29) {real, imag} */,
  {32'hbf35d214, 32'h00000000} /* (17, 1, 28) {real, imag} */,
  {32'hbf491025, 32'h00000000} /* (17, 1, 27) {real, imag} */,
  {32'hbf8e6acd, 32'h00000000} /* (17, 1, 26) {real, imag} */,
  {32'hbf8310d6, 32'h00000000} /* (17, 1, 25) {real, imag} */,
  {32'hbf1e34ba, 32'h00000000} /* (17, 1, 24) {real, imag} */,
  {32'hbf2dccaf, 32'h00000000} /* (17, 1, 23) {real, imag} */,
  {32'hbf5ccf4c, 32'h00000000} /* (17, 1, 22) {real, imag} */,
  {32'hbf138edf, 32'h00000000} /* (17, 1, 21) {real, imag} */,
  {32'hbf5894d3, 32'h00000000} /* (17, 1, 20) {real, imag} */,
  {32'hbfb131c7, 32'h00000000} /* (17, 1, 19) {real, imag} */,
  {32'hc027e9bd, 32'h00000000} /* (17, 1, 18) {real, imag} */,
  {32'hbffe628f, 32'h00000000} /* (17, 1, 17) {real, imag} */,
  {32'hbf173227, 32'h00000000} /* (17, 1, 16) {real, imag} */,
  {32'h3f4906f6, 32'h00000000} /* (17, 1, 15) {real, imag} */,
  {32'h3fca8b0f, 32'h00000000} /* (17, 1, 14) {real, imag} */,
  {32'h3fbd7f32, 32'h00000000} /* (17, 1, 13) {real, imag} */,
  {32'h3f8ec47f, 32'h00000000} /* (17, 1, 12) {real, imag} */,
  {32'h3f7df4b1, 32'h00000000} /* (17, 1, 11) {real, imag} */,
  {32'h3f26fa7c, 32'h00000000} /* (17, 1, 10) {real, imag} */,
  {32'h3ec2bcba, 32'h00000000} /* (17, 1, 9) {real, imag} */,
  {32'h3f50088c, 32'h00000000} /* (17, 1, 8) {real, imag} */,
  {32'h3f0e1911, 32'h00000000} /* (17, 1, 7) {real, imag} */,
  {32'h3e92be9f, 32'h00000000} /* (17, 1, 6) {real, imag} */,
  {32'hbf06e3b2, 32'h00000000} /* (17, 1, 5) {real, imag} */,
  {32'hbf89b0a8, 32'h00000000} /* (17, 1, 4) {real, imag} */,
  {32'hbf0c34a5, 32'h00000000} /* (17, 1, 3) {real, imag} */,
  {32'hbf418b73, 32'h00000000} /* (17, 1, 2) {real, imag} */,
  {32'hbf3c82b1, 32'h00000000} /* (17, 1, 1) {real, imag} */,
  {32'hbe9f8b55, 32'h00000000} /* (17, 1, 0) {real, imag} */,
  {32'hbea91bd3, 32'h00000000} /* (17, 0, 31) {real, imag} */,
  {32'hbe961460, 32'h00000000} /* (17, 0, 30) {real, imag} */,
  {32'hbef8cfac, 32'h00000000} /* (17, 0, 29) {real, imag} */,
  {32'hbee2a519, 32'h00000000} /* (17, 0, 28) {real, imag} */,
  {32'hbf0372bc, 32'h00000000} /* (17, 0, 27) {real, imag} */,
  {32'hbf29add8, 32'h00000000} /* (17, 0, 26) {real, imag} */,
  {32'hbf08bbb1, 32'h00000000} /* (17, 0, 25) {real, imag} */,
  {32'hbed486d9, 32'h00000000} /* (17, 0, 24) {real, imag} */,
  {32'hbf11b9aa, 32'h00000000} /* (17, 0, 23) {real, imag} */,
  {32'hbf589a22, 32'h00000000} /* (17, 0, 22) {real, imag} */,
  {32'hbf416f1c, 32'h00000000} /* (17, 0, 21) {real, imag} */,
  {32'hbf4b5eb7, 32'h00000000} /* (17, 0, 20) {real, imag} */,
  {32'hbf27a603, 32'h00000000} /* (17, 0, 19) {real, imag} */,
  {32'hbf6149b0, 32'h00000000} /* (17, 0, 18) {real, imag} */,
  {32'hbf1e4565, 32'h00000000} /* (17, 0, 17) {real, imag} */,
  {32'hbe21e509, 32'h00000000} /* (17, 0, 16) {real, imag} */,
  {32'h3eaba22f, 32'h00000000} /* (17, 0, 15) {real, imag} */,
  {32'h3f2d5354, 32'h00000000} /* (17, 0, 14) {real, imag} */,
  {32'h3f115fdd, 32'h00000000} /* (17, 0, 13) {real, imag} */,
  {32'h3f39eccd, 32'h00000000} /* (17, 0, 12) {real, imag} */,
  {32'h3f6f7c49, 32'h00000000} /* (17, 0, 11) {real, imag} */,
  {32'h3f0d9a63, 32'h00000000} /* (17, 0, 10) {real, imag} */,
  {32'h3e4099ab, 32'h00000000} /* (17, 0, 9) {real, imag} */,
  {32'h3eda0898, 32'h00000000} /* (17, 0, 8) {real, imag} */,
  {32'h3ea95bcc, 32'h00000000} /* (17, 0, 7) {real, imag} */,
  {32'h3e92c084, 32'h00000000} /* (17, 0, 6) {real, imag} */,
  {32'h3b89b68f, 32'h00000000} /* (17, 0, 5) {real, imag} */,
  {32'hbeafc1c4, 32'h00000000} /* (17, 0, 4) {real, imag} */,
  {32'hbe90cd14, 32'h00000000} /* (17, 0, 3) {real, imag} */,
  {32'hbee2b5a3, 32'h00000000} /* (17, 0, 2) {real, imag} */,
  {32'hbe865aa7, 32'h00000000} /* (17, 0, 1) {real, imag} */,
  {32'hbe187b99, 32'h00000000} /* (17, 0, 0) {real, imag} */,
  {32'hbe0cf9e0, 32'h00000000} /* (16, 31, 31) {real, imag} */,
  {32'hbe594e83, 32'h00000000} /* (16, 31, 30) {real, imag} */,
  {32'hbe737a66, 32'h00000000} /* (16, 31, 29) {real, imag} */,
  {32'hbe98ac1b, 32'h00000000} /* (16, 31, 28) {real, imag} */,
  {32'hbe770072, 32'h00000000} /* (16, 31, 27) {real, imag} */,
  {32'h3cb5372e, 32'h00000000} /* (16, 31, 26) {real, imag} */,
  {32'hbe5d73ce, 32'h00000000} /* (16, 31, 25) {real, imag} */,
  {32'hbeec3258, 32'h00000000} /* (16, 31, 24) {real, imag} */,
  {32'hbf230654, 32'h00000000} /* (16, 31, 23) {real, imag} */,
  {32'hbf2d3cfc, 32'h00000000} /* (16, 31, 22) {real, imag} */,
  {32'hbe8e4648, 32'h00000000} /* (16, 31, 21) {real, imag} */,
  {32'hbe2fd7f1, 32'h00000000} /* (16, 31, 20) {real, imag} */,
  {32'hbc975980, 32'h00000000} /* (16, 31, 19) {real, imag} */,
  {32'hbc0ab9e0, 32'h00000000} /* (16, 31, 18) {real, imag} */,
  {32'hbddc5d06, 32'h00000000} /* (16, 31, 17) {real, imag} */,
  {32'hbe0277f0, 32'h00000000} /* (16, 31, 16) {real, imag} */,
  {32'hbe87829f, 32'h00000000} /* (16, 31, 15) {real, imag} */,
  {32'h3d917104, 32'h00000000} /* (16, 31, 14) {real, imag} */,
  {32'h3d13a5ac, 32'h00000000} /* (16, 31, 13) {real, imag} */,
  {32'h3e51251e, 32'h00000000} /* (16, 31, 12) {real, imag} */,
  {32'h3e584e5e, 32'h00000000} /* (16, 31, 11) {real, imag} */,
  {32'hbdfdf004, 32'h00000000} /* (16, 31, 10) {real, imag} */,
  {32'hbe6a119e, 32'h00000000} /* (16, 31, 9) {real, imag} */,
  {32'hbf14e656, 32'h00000000} /* (16, 31, 8) {real, imag} */,
  {32'hbf2795ee, 32'h00000000} /* (16, 31, 7) {real, imag} */,
  {32'hbd74d3af, 32'h00000000} /* (16, 31, 6) {real, imag} */,
  {32'hbecbc9f3, 32'h00000000} /* (16, 31, 5) {real, imag} */,
  {32'hbebaacfe, 32'h00000000} /* (16, 31, 4) {real, imag} */,
  {32'hbedd0f67, 32'h00000000} /* (16, 31, 3) {real, imag} */,
  {32'hbdfa71f2, 32'h00000000} /* (16, 31, 2) {real, imag} */,
  {32'h3a5901fc, 32'h00000000} /* (16, 31, 1) {real, imag} */,
  {32'hbe0721f7, 32'h00000000} /* (16, 31, 0) {real, imag} */,
  {32'h3cf599e6, 32'h00000000} /* (16, 30, 31) {real, imag} */,
  {32'hbed476f4, 32'h00000000} /* (16, 30, 30) {real, imag} */,
  {32'hbf7abcc5, 32'h00000000} /* (16, 30, 29) {real, imag} */,
  {32'hbf5f92cc, 32'h00000000} /* (16, 30, 28) {real, imag} */,
  {32'hbf402512, 32'h00000000} /* (16, 30, 27) {real, imag} */,
  {32'hbdff5674, 32'h00000000} /* (16, 30, 26) {real, imag} */,
  {32'h3d107d7b, 32'h00000000} /* (16, 30, 25) {real, imag} */,
  {32'hbe48c741, 32'h00000000} /* (16, 30, 24) {real, imag} */,
  {32'hbefc99fa, 32'h00000000} /* (16, 30, 23) {real, imag} */,
  {32'hbef99ff5, 32'h00000000} /* (16, 30, 22) {real, imag} */,
  {32'hbd73104a, 32'h00000000} /* (16, 30, 21) {real, imag} */,
  {32'h3f0a3c2c, 32'h00000000} /* (16, 30, 20) {real, imag} */,
  {32'h3f356dd2, 32'h00000000} /* (16, 30, 19) {real, imag} */,
  {32'h3ea9e1dd, 32'h00000000} /* (16, 30, 18) {real, imag} */,
  {32'h3e35e9c7, 32'h00000000} /* (16, 30, 17) {real, imag} */,
  {32'h3df18115, 32'h00000000} /* (16, 30, 16) {real, imag} */,
  {32'h3f123e3a, 32'h00000000} /* (16, 30, 15) {real, imag} */,
  {32'h3f0b7825, 32'h00000000} /* (16, 30, 14) {real, imag} */,
  {32'h3e6fd4d2, 32'h00000000} /* (16, 30, 13) {real, imag} */,
  {32'h3e8c8446, 32'h00000000} /* (16, 30, 12) {real, imag} */,
  {32'h3eb95e24, 32'h00000000} /* (16, 30, 11) {real, imag} */,
  {32'hbd2814ea, 32'h00000000} /* (16, 30, 10) {real, imag} */,
  {32'hbf3bcfe5, 32'h00000000} /* (16, 30, 9) {real, imag} */,
  {32'hbf84f1d0, 32'h00000000} /* (16, 30, 8) {real, imag} */,
  {32'hbf938193, 32'h00000000} /* (16, 30, 7) {real, imag} */,
  {32'hbec1047e, 32'h00000000} /* (16, 30, 6) {real, imag} */,
  {32'hbe87e0cf, 32'h00000000} /* (16, 30, 5) {real, imag} */,
  {32'hbf5b79c9, 32'h00000000} /* (16, 30, 4) {real, imag} */,
  {32'hbf4393e3, 32'h00000000} /* (16, 30, 3) {real, imag} */,
  {32'hbf5b2145, 32'h00000000} /* (16, 30, 2) {real, imag} */,
  {32'hbc87e58e, 32'h00000000} /* (16, 30, 1) {real, imag} */,
  {32'h3d37ff68, 32'h00000000} /* (16, 30, 0) {real, imag} */,
  {32'hbca345ec, 32'h00000000} /* (16, 29, 31) {real, imag} */,
  {32'hbefe8f4b, 32'h00000000} /* (16, 29, 30) {real, imag} */,
  {32'hbf710ce6, 32'h00000000} /* (16, 29, 29) {real, imag} */,
  {32'hbf3f50a9, 32'h00000000} /* (16, 29, 28) {real, imag} */,
  {32'hbf1f94ff, 32'h00000000} /* (16, 29, 27) {real, imag} */,
  {32'hbda0af76, 32'h00000000} /* (16, 29, 26) {real, imag} */,
  {32'hbddd37cb, 32'h00000000} /* (16, 29, 25) {real, imag} */,
  {32'hbf2e1072, 32'h00000000} /* (16, 29, 24) {real, imag} */,
  {32'hbf737eff, 32'h00000000} /* (16, 29, 23) {real, imag} */,
  {32'hbd1f7679, 32'h00000000} /* (16, 29, 22) {real, imag} */,
  {32'h3f15b95a, 32'h00000000} /* (16, 29, 21) {real, imag} */,
  {32'h3f8a171f, 32'h00000000} /* (16, 29, 20) {real, imag} */,
  {32'h3f5051b6, 32'h00000000} /* (16, 29, 19) {real, imag} */,
  {32'h3f51ac22, 32'h00000000} /* (16, 29, 18) {real, imag} */,
  {32'h3f95d354, 32'h00000000} /* (16, 29, 17) {real, imag} */,
  {32'h3f3f3473, 32'h00000000} /* (16, 29, 16) {real, imag} */,
  {32'h3f881472, 32'h00000000} /* (16, 29, 15) {real, imag} */,
  {32'h3f7984b0, 32'h00000000} /* (16, 29, 14) {real, imag} */,
  {32'h3f74ef2b, 32'h00000000} /* (16, 29, 13) {real, imag} */,
  {32'h3f78c5a5, 32'h00000000} /* (16, 29, 12) {real, imag} */,
  {32'h3f696443, 32'h00000000} /* (16, 29, 11) {real, imag} */,
  {32'h3ed49db9, 32'h00000000} /* (16, 29, 10) {real, imag} */,
  {32'hbf4bbd4b, 32'h00000000} /* (16, 29, 9) {real, imag} */,
  {32'hbf8ecb12, 32'h00000000} /* (16, 29, 8) {real, imag} */,
  {32'hbf4c0e31, 32'h00000000} /* (16, 29, 7) {real, imag} */,
  {32'hbf476caf, 32'h00000000} /* (16, 29, 6) {real, imag} */,
  {32'hbe5886ac, 32'h00000000} /* (16, 29, 5) {real, imag} */,
  {32'hbf0a7ac5, 32'h00000000} /* (16, 29, 4) {real, imag} */,
  {32'hbf729d85, 32'h00000000} /* (16, 29, 3) {real, imag} */,
  {32'hbfaf9670, 32'h00000000} /* (16, 29, 2) {real, imag} */,
  {32'hbf56d460, 32'h00000000} /* (16, 29, 1) {real, imag} */,
  {32'hbe94d2ce, 32'h00000000} /* (16, 29, 0) {real, imag} */,
  {32'hbf048776, 32'h00000000} /* (16, 28, 31) {real, imag} */,
  {32'hbf30f5b8, 32'h00000000} /* (16, 28, 30) {real, imag} */,
  {32'hbea5b5f7, 32'h00000000} /* (16, 28, 29) {real, imag} */,
  {32'hbe90b256, 32'h00000000} /* (16, 28, 28) {real, imag} */,
  {32'hbf1c974f, 32'h00000000} /* (16, 28, 27) {real, imag} */,
  {32'hbe9b7f04, 32'h00000000} /* (16, 28, 26) {real, imag} */,
  {32'hbf275e15, 32'h00000000} /* (16, 28, 25) {real, imag} */,
  {32'hbf8f292c, 32'h00000000} /* (16, 28, 24) {real, imag} */,
  {32'hbf795fbb, 32'h00000000} /* (16, 28, 23) {real, imag} */,
  {32'h3e6d6a8e, 32'h00000000} /* (16, 28, 22) {real, imag} */,
  {32'h3f0cefad, 32'h00000000} /* (16, 28, 21) {real, imag} */,
  {32'h3e36ccd1, 32'h00000000} /* (16, 28, 20) {real, imag} */,
  {32'h3d70f9d0, 32'h00000000} /* (16, 28, 19) {real, imag} */,
  {32'h3f8dd91f, 32'h00000000} /* (16, 28, 18) {real, imag} */,
  {32'h3f48293d, 32'h00000000} /* (16, 28, 17) {real, imag} */,
  {32'h3f108c33, 32'h00000000} /* (16, 28, 16) {real, imag} */,
  {32'h3f8d6713, 32'h00000000} /* (16, 28, 15) {real, imag} */,
  {32'h3f98fbe4, 32'h00000000} /* (16, 28, 14) {real, imag} */,
  {32'h3f9c1438, 32'h00000000} /* (16, 28, 13) {real, imag} */,
  {32'h3f7cce44, 32'h00000000} /* (16, 28, 12) {real, imag} */,
  {32'h3f565dfb, 32'h00000000} /* (16, 28, 11) {real, imag} */,
  {32'h3e86d488, 32'h00000000} /* (16, 28, 10) {real, imag} */,
  {32'hbf59d6ef, 32'h00000000} /* (16, 28, 9) {real, imag} */,
  {32'hbf008ed2, 32'h00000000} /* (16, 28, 8) {real, imag} */,
  {32'hbedc68f1, 32'h00000000} /* (16, 28, 7) {real, imag} */,
  {32'hbf30d6a9, 32'h00000000} /* (16, 28, 6) {real, imag} */,
  {32'hbe88ca12, 32'h00000000} /* (16, 28, 5) {real, imag} */,
  {32'hbf0cd57d, 32'h00000000} /* (16, 28, 4) {real, imag} */,
  {32'hbf968e77, 32'h00000000} /* (16, 28, 3) {real, imag} */,
  {32'hbf9e5283, 32'h00000000} /* (16, 28, 2) {real, imag} */,
  {32'hbf8662fc, 32'h00000000} /* (16, 28, 1) {real, imag} */,
  {32'hbe9422c2, 32'h00000000} /* (16, 28, 0) {real, imag} */,
  {32'hbebe00bf, 32'h00000000} /* (16, 27, 31) {real, imag} */,
  {32'hbf03f4fc, 32'h00000000} /* (16, 27, 30) {real, imag} */,
  {32'hbec42d46, 32'h00000000} /* (16, 27, 29) {real, imag} */,
  {32'hbed84a3f, 32'h00000000} /* (16, 27, 28) {real, imag} */,
  {32'hbf10d20e, 32'h00000000} /* (16, 27, 27) {real, imag} */,
  {32'hbe25e9f5, 32'h00000000} /* (16, 27, 26) {real, imag} */,
  {32'hbe0dc50d, 32'h00000000} /* (16, 27, 25) {real, imag} */,
  {32'hbf6a3571, 32'h00000000} /* (16, 27, 24) {real, imag} */,
  {32'hbf3b95da, 32'h00000000} /* (16, 27, 23) {real, imag} */,
  {32'hbe03578f, 32'h00000000} /* (16, 27, 22) {real, imag} */,
  {32'h3eeec63a, 32'h00000000} /* (16, 27, 21) {real, imag} */,
  {32'h3efdb403, 32'h00000000} /* (16, 27, 20) {real, imag} */,
  {32'h3eae3cbb, 32'h00000000} /* (16, 27, 19) {real, imag} */,
  {32'h3f1f411d, 32'h00000000} /* (16, 27, 18) {real, imag} */,
  {32'h3e4d4344, 32'h00000000} /* (16, 27, 17) {real, imag} */,
  {32'h3e35a99c, 32'h00000000} /* (16, 27, 16) {real, imag} */,
  {32'h3f38bb22, 32'h00000000} /* (16, 27, 15) {real, imag} */,
  {32'h3f356d4b, 32'h00000000} /* (16, 27, 14) {real, imag} */,
  {32'h3f0698c4, 32'h00000000} /* (16, 27, 13) {real, imag} */,
  {32'h3f09eefa, 32'h00000000} /* (16, 27, 12) {real, imag} */,
  {32'h3f1b9044, 32'h00000000} /* (16, 27, 11) {real, imag} */,
  {32'h3d92a9eb, 32'h00000000} /* (16, 27, 10) {real, imag} */,
  {32'hbf3e2d47, 32'h00000000} /* (16, 27, 9) {real, imag} */,
  {32'hbf11d240, 32'h00000000} /* (16, 27, 8) {real, imag} */,
  {32'hbf42c1af, 32'h00000000} /* (16, 27, 7) {real, imag} */,
  {32'hbf10b2a6, 32'h00000000} /* (16, 27, 6) {real, imag} */,
  {32'hbe5abd33, 32'h00000000} /* (16, 27, 5) {real, imag} */,
  {32'hbf1eca76, 32'h00000000} /* (16, 27, 4) {real, imag} */,
  {32'hbf2d8691, 32'h00000000} /* (16, 27, 3) {real, imag} */,
  {32'hbf421787, 32'h00000000} /* (16, 27, 2) {real, imag} */,
  {32'hbf517a01, 32'h00000000} /* (16, 27, 1) {real, imag} */,
  {32'hbeb75030, 32'h00000000} /* (16, 27, 0) {real, imag} */,
  {32'hbeb39e52, 32'h00000000} /* (16, 26, 31) {real, imag} */,
  {32'hbf208ea8, 32'h00000000} /* (16, 26, 30) {real, imag} */,
  {32'hbe904b23, 32'h00000000} /* (16, 26, 29) {real, imag} */,
  {32'hbeab5f46, 32'h00000000} /* (16, 26, 28) {real, imag} */,
  {32'hbf265145, 32'h00000000} /* (16, 26, 27) {real, imag} */,
  {32'hbec49341, 32'h00000000} /* (16, 26, 26) {real, imag} */,
  {32'hbea4e0f1, 32'h00000000} /* (16, 26, 25) {real, imag} */,
  {32'hbf5e176b, 32'h00000000} /* (16, 26, 24) {real, imag} */,
  {32'hbec6f71f, 32'h00000000} /* (16, 26, 23) {real, imag} */,
  {32'hbe351f41, 32'h00000000} /* (16, 26, 22) {real, imag} */,
  {32'h3e674346, 32'h00000000} /* (16, 26, 21) {real, imag} */,
  {32'h3f2cabce, 32'h00000000} /* (16, 26, 20) {real, imag} */,
  {32'h3e98fe24, 32'h00000000} /* (16, 26, 19) {real, imag} */,
  {32'h3d715955, 32'h00000000} /* (16, 26, 18) {real, imag} */,
  {32'h3e4d10e7, 32'h00000000} /* (16, 26, 17) {real, imag} */,
  {32'h3e153ef4, 32'h00000000} /* (16, 26, 16) {real, imag} */,
  {32'h3eb609a6, 32'h00000000} /* (16, 26, 15) {real, imag} */,
  {32'h3eb44de0, 32'h00000000} /* (16, 26, 14) {real, imag} */,
  {32'h3e931a25, 32'h00000000} /* (16, 26, 13) {real, imag} */,
  {32'h3e88fe9c, 32'h00000000} /* (16, 26, 12) {real, imag} */,
  {32'h3eb4c14c, 32'h00000000} /* (16, 26, 11) {real, imag} */,
  {32'hbd981c0f, 32'h00000000} /* (16, 26, 10) {real, imag} */,
  {32'hbf40f092, 32'h00000000} /* (16, 26, 9) {real, imag} */,
  {32'hbf3dd4a2, 32'h00000000} /* (16, 26, 8) {real, imag} */,
  {32'hbf289556, 32'h00000000} /* (16, 26, 7) {real, imag} */,
  {32'hbf28f2b0, 32'h00000000} /* (16, 26, 6) {real, imag} */,
  {32'hbedabc89, 32'h00000000} /* (16, 26, 5) {real, imag} */,
  {32'hbecba50c, 32'h00000000} /* (16, 26, 4) {real, imag} */,
  {32'hbe9a9ee0, 32'h00000000} /* (16, 26, 3) {real, imag} */,
  {32'hbf6e1f75, 32'h00000000} /* (16, 26, 2) {real, imag} */,
  {32'hbf7bce25, 32'h00000000} /* (16, 26, 1) {real, imag} */,
  {32'hbee960d2, 32'h00000000} /* (16, 26, 0) {real, imag} */,
  {32'hbee798e5, 32'h00000000} /* (16, 25, 31) {real, imag} */,
  {32'hbf58582c, 32'h00000000} /* (16, 25, 30) {real, imag} */,
  {32'hbf38087c, 32'h00000000} /* (16, 25, 29) {real, imag} */,
  {32'hbebf983f, 32'h00000000} /* (16, 25, 28) {real, imag} */,
  {32'hbebd2f87, 32'h00000000} /* (16, 25, 27) {real, imag} */,
  {32'hbeb35bbc, 32'h00000000} /* (16, 25, 26) {real, imag} */,
  {32'hbf01e118, 32'h00000000} /* (16, 25, 25) {real, imag} */,
  {32'hbf4fb3bb, 32'h00000000} /* (16, 25, 24) {real, imag} */,
  {32'hbf3b4d62, 32'h00000000} /* (16, 25, 23) {real, imag} */,
  {32'hbf188bce, 32'h00000000} /* (16, 25, 22) {real, imag} */,
  {32'h3dfe70db, 32'h00000000} /* (16, 25, 21) {real, imag} */,
  {32'h3f51b9dd, 32'h00000000} /* (16, 25, 20) {real, imag} */,
  {32'h3f1d64f4, 32'h00000000} /* (16, 25, 19) {real, imag} */,
  {32'h3db490f0, 32'h00000000} /* (16, 25, 18) {real, imag} */,
  {32'h3edb3bf9, 32'h00000000} /* (16, 25, 17) {real, imag} */,
  {32'h3f0d15e2, 32'h00000000} /* (16, 25, 16) {real, imag} */,
  {32'h3f0fc698, 32'h00000000} /* (16, 25, 15) {real, imag} */,
  {32'h3e878d08, 32'h00000000} /* (16, 25, 14) {real, imag} */,
  {32'h3f154f91, 32'h00000000} /* (16, 25, 13) {real, imag} */,
  {32'h3f33e69d, 32'h00000000} /* (16, 25, 12) {real, imag} */,
  {32'h3f502c0e, 32'h00000000} /* (16, 25, 11) {real, imag} */,
  {32'hbe33a2e6, 32'h00000000} /* (16, 25, 10) {real, imag} */,
  {32'hbf4d4853, 32'h00000000} /* (16, 25, 9) {real, imag} */,
  {32'hbe60e8b4, 32'h00000000} /* (16, 25, 8) {real, imag} */,
  {32'hbdef2f82, 32'h00000000} /* (16, 25, 7) {real, imag} */,
  {32'hbeeab5eb, 32'h00000000} /* (16, 25, 6) {real, imag} */,
  {32'hbee94585, 32'h00000000} /* (16, 25, 5) {real, imag} */,
  {32'hbf030b26, 32'h00000000} /* (16, 25, 4) {real, imag} */,
  {32'hbf5906b3, 32'h00000000} /* (16, 25, 3) {real, imag} */,
  {32'hbf8901cc, 32'h00000000} /* (16, 25, 2) {real, imag} */,
  {32'hbf76b2b5, 32'h00000000} /* (16, 25, 1) {real, imag} */,
  {32'hbea4f81b, 32'h00000000} /* (16, 25, 0) {real, imag} */,
  {32'hbf0bd73d, 32'h00000000} /* (16, 24, 31) {real, imag} */,
  {32'hbed1964e, 32'h00000000} /* (16, 24, 30) {real, imag} */,
  {32'hbda35ec0, 32'h00000000} /* (16, 24, 29) {real, imag} */,
  {32'hbe1d9aa9, 32'h00000000} /* (16, 24, 28) {real, imag} */,
  {32'hbf1fed62, 32'h00000000} /* (16, 24, 27) {real, imag} */,
  {32'hbf49cd0c, 32'h00000000} /* (16, 24, 26) {real, imag} */,
  {32'hbf32deb6, 32'h00000000} /* (16, 24, 25) {real, imag} */,
  {32'hbf877ce5, 32'h00000000} /* (16, 24, 24) {real, imag} */,
  {32'hbf8f1dc3, 32'h00000000} /* (16, 24, 23) {real, imag} */,
  {32'hbf6f43ba, 32'h00000000} /* (16, 24, 22) {real, imag} */,
  {32'hbe7e8213, 32'h00000000} /* (16, 24, 21) {real, imag} */,
  {32'h3eef6795, 32'h00000000} /* (16, 24, 20) {real, imag} */,
  {32'h3f2c22c5, 32'h00000000} /* (16, 24, 19) {real, imag} */,
  {32'h3ee7513f, 32'h00000000} /* (16, 24, 18) {real, imag} */,
  {32'h3f5a7125, 32'h00000000} /* (16, 24, 17) {real, imag} */,
  {32'h3f38a5ec, 32'h00000000} /* (16, 24, 16) {real, imag} */,
  {32'h3eabecb9, 32'h00000000} /* (16, 24, 15) {real, imag} */,
  {32'h3ecd390f, 32'h00000000} /* (16, 24, 14) {real, imag} */,
  {32'h3f56b498, 32'h00000000} /* (16, 24, 13) {real, imag} */,
  {32'h3fb6e383, 32'h00000000} /* (16, 24, 12) {real, imag} */,
  {32'h3f46938a, 32'h00000000} /* (16, 24, 11) {real, imag} */,
  {32'hbf21a065, 32'h00000000} /* (16, 24, 10) {real, imag} */,
  {32'hbf86a8d6, 32'h00000000} /* (16, 24, 9) {real, imag} */,
  {32'hbf11afa3, 32'h00000000} /* (16, 24, 8) {real, imag} */,
  {32'hbe8ae611, 32'h00000000} /* (16, 24, 7) {real, imag} */,
  {32'hbecbbc60, 32'h00000000} /* (16, 24, 6) {real, imag} */,
  {32'hbf3a676c, 32'h00000000} /* (16, 24, 5) {real, imag} */,
  {32'hbee7573f, 32'h00000000} /* (16, 24, 4) {real, imag} */,
  {32'hbf7046f8, 32'h00000000} /* (16, 24, 3) {real, imag} */,
  {32'hbfb0cc1a, 32'h00000000} /* (16, 24, 2) {real, imag} */,
  {32'hbf842906, 32'h00000000} /* (16, 24, 1) {real, imag} */,
  {32'hbe955085, 32'h00000000} /* (16, 24, 0) {real, imag} */,
  {32'hbecb942a, 32'h00000000} /* (16, 23, 31) {real, imag} */,
  {32'hbdfa27c9, 32'h00000000} /* (16, 23, 30) {real, imag} */,
  {32'h3d3ea021, 32'h00000000} /* (16, 23, 29) {real, imag} */,
  {32'hbed5318d, 32'h00000000} /* (16, 23, 28) {real, imag} */,
  {32'hbf738a11, 32'h00000000} /* (16, 23, 27) {real, imag} */,
  {32'hbf99d5d6, 32'h00000000} /* (16, 23, 26) {real, imag} */,
  {32'hbf3be55c, 32'h00000000} /* (16, 23, 25) {real, imag} */,
  {32'hbf42c5ba, 32'h00000000} /* (16, 23, 24) {real, imag} */,
  {32'hbfaedc4c, 32'h00000000} /* (16, 23, 23) {real, imag} */,
  {32'hbf7a1ccb, 32'h00000000} /* (16, 23, 22) {real, imag} */,
  {32'hbeb4befc, 32'h00000000} /* (16, 23, 21) {real, imag} */,
  {32'h3f32d293, 32'h00000000} /* (16, 23, 20) {real, imag} */,
  {32'h3edff445, 32'h00000000} /* (16, 23, 19) {real, imag} */,
  {32'h3ec8ddd3, 32'h00000000} /* (16, 23, 18) {real, imag} */,
  {32'h3ec3ded0, 32'h00000000} /* (16, 23, 17) {real, imag} */,
  {32'h3f0fdbb7, 32'h00000000} /* (16, 23, 16) {real, imag} */,
  {32'h3f319d29, 32'h00000000} /* (16, 23, 15) {real, imag} */,
  {32'h3f1be58d, 32'h00000000} /* (16, 23, 14) {real, imag} */,
  {32'h3f53a8ff, 32'h00000000} /* (16, 23, 13) {real, imag} */,
  {32'h3f424bd7, 32'h00000000} /* (16, 23, 12) {real, imag} */,
  {32'h3e270230, 32'h00000000} /* (16, 23, 11) {real, imag} */,
  {32'hbf32fe47, 32'h00000000} /* (16, 23, 10) {real, imag} */,
  {32'hbf492bd3, 32'h00000000} /* (16, 23, 9) {real, imag} */,
  {32'hbf516132, 32'h00000000} /* (16, 23, 8) {real, imag} */,
  {32'hbe58a841, 32'h00000000} /* (16, 23, 7) {real, imag} */,
  {32'hbeea1988, 32'h00000000} /* (16, 23, 6) {real, imag} */,
  {32'hbf4d55ba, 32'h00000000} /* (16, 23, 5) {real, imag} */,
  {32'hbd4e6cc4, 32'h00000000} /* (16, 23, 4) {real, imag} */,
  {32'hbdd7db4b, 32'h00000000} /* (16, 23, 3) {real, imag} */,
  {32'hbf6f8173, 32'h00000000} /* (16, 23, 2) {real, imag} */,
  {32'hbf7364e7, 32'h00000000} /* (16, 23, 1) {real, imag} */,
  {32'hbec0e8eb, 32'h00000000} /* (16, 23, 0) {real, imag} */,
  {32'hbf0e9801, 32'h00000000} /* (16, 22, 31) {real, imag} */,
  {32'hbec2f322, 32'h00000000} /* (16, 22, 30) {real, imag} */,
  {32'hbea74d17, 32'h00000000} /* (16, 22, 29) {real, imag} */,
  {32'hbea86ab5, 32'h00000000} /* (16, 22, 28) {real, imag} */,
  {32'hbed1cd70, 32'h00000000} /* (16, 22, 27) {real, imag} */,
  {32'hbf381377, 32'h00000000} /* (16, 22, 26) {real, imag} */,
  {32'hbf5c2bb8, 32'h00000000} /* (16, 22, 25) {real, imag} */,
  {32'hbf4ac907, 32'h00000000} /* (16, 22, 24) {real, imag} */,
  {32'hbf5d2c89, 32'h00000000} /* (16, 22, 23) {real, imag} */,
  {32'hbf770297, 32'h00000000} /* (16, 22, 22) {real, imag} */,
  {32'hbf0dc79a, 32'h00000000} /* (16, 22, 21) {real, imag} */,
  {32'h3f1d7a8b, 32'h00000000} /* (16, 22, 20) {real, imag} */,
  {32'h3f01d620, 32'h00000000} /* (16, 22, 19) {real, imag} */,
  {32'h3e78eb0a, 32'h00000000} /* (16, 22, 18) {real, imag} */,
  {32'h3e8ad155, 32'h00000000} /* (16, 22, 17) {real, imag} */,
  {32'h3eb5a5c1, 32'h00000000} /* (16, 22, 16) {real, imag} */,
  {32'h3f22f60a, 32'h00000000} /* (16, 22, 15) {real, imag} */,
  {32'h3f49089c, 32'h00000000} /* (16, 22, 14) {real, imag} */,
  {32'h3f5556bd, 32'h00000000} /* (16, 22, 13) {real, imag} */,
  {32'h3e6b94b7, 32'h00000000} /* (16, 22, 12) {real, imag} */,
  {32'h3e65bf10, 32'h00000000} /* (16, 22, 11) {real, imag} */,
  {32'hbe6f889c, 32'h00000000} /* (16, 22, 10) {real, imag} */,
  {32'hbf47ca77, 32'h00000000} /* (16, 22, 9) {real, imag} */,
  {32'hbf793712, 32'h00000000} /* (16, 22, 8) {real, imag} */,
  {32'hbf3013ac, 32'h00000000} /* (16, 22, 7) {real, imag} */,
  {32'hbf368bbb, 32'h00000000} /* (16, 22, 6) {real, imag} */,
  {32'hbee2b6ee, 32'h00000000} /* (16, 22, 5) {real, imag} */,
  {32'hbea0137f, 32'h00000000} /* (16, 22, 4) {real, imag} */,
  {32'hbf048ce8, 32'h00000000} /* (16, 22, 3) {real, imag} */,
  {32'hbf250c8d, 32'h00000000} /* (16, 22, 2) {real, imag} */,
  {32'hbf597c9a, 32'h00000000} /* (16, 22, 1) {real, imag} */,
  {32'hbee41f2c, 32'h00000000} /* (16, 22, 0) {real, imag} */,
  {32'hbe0f5ef6, 32'h00000000} /* (16, 21, 31) {real, imag} */,
  {32'hbe356250, 32'h00000000} /* (16, 21, 30) {real, imag} */,
  {32'hbf0335f7, 32'h00000000} /* (16, 21, 29) {real, imag} */,
  {32'hbed1f98b, 32'h00000000} /* (16, 21, 28) {real, imag} */,
  {32'hbf116aeb, 32'h00000000} /* (16, 21, 27) {real, imag} */,
  {32'hbf2916d5, 32'h00000000} /* (16, 21, 26) {real, imag} */,
  {32'hbf199390, 32'h00000000} /* (16, 21, 25) {real, imag} */,
  {32'hbebd20a2, 32'h00000000} /* (16, 21, 24) {real, imag} */,
  {32'hbd3751ea, 32'h00000000} /* (16, 21, 23) {real, imag} */,
  {32'hbe3afd95, 32'h00000000} /* (16, 21, 22) {real, imag} */,
  {32'hbe9fea62, 32'h00000000} /* (16, 21, 21) {real, imag} */,
  {32'hbdf054c8, 32'h00000000} /* (16, 21, 20) {real, imag} */,
  {32'h3ea7e41e, 32'h00000000} /* (16, 21, 19) {real, imag} */,
  {32'hbd3c4a01, 32'h00000000} /* (16, 21, 18) {real, imag} */,
  {32'hbb28e0cc, 32'h00000000} /* (16, 21, 17) {real, imag} */,
  {32'h3d0c9ab8, 32'h00000000} /* (16, 21, 16) {real, imag} */,
  {32'h3f19e851, 32'h00000000} /* (16, 21, 15) {real, imag} */,
  {32'h3efc1b19, 32'h00000000} /* (16, 21, 14) {real, imag} */,
  {32'hbe074947, 32'h00000000} /* (16, 21, 13) {real, imag} */,
  {32'hbec7b7ad, 32'h00000000} /* (16, 21, 12) {real, imag} */,
  {32'hbe35ef64, 32'h00000000} /* (16, 21, 11) {real, imag} */,
  {32'hbdcdeb46, 32'h00000000} /* (16, 21, 10) {real, imag} */,
  {32'hbed52e74, 32'h00000000} /* (16, 21, 9) {real, imag} */,
  {32'hbf46e888, 32'h00000000} /* (16, 21, 8) {real, imag} */,
  {32'hbee70639, 32'h00000000} /* (16, 21, 7) {real, imag} */,
  {32'hbf1076a0, 32'h00000000} /* (16, 21, 6) {real, imag} */,
  {32'hbeb3103d, 32'h00000000} /* (16, 21, 5) {real, imag} */,
  {32'hbd8aa5db, 32'h00000000} /* (16, 21, 4) {real, imag} */,
  {32'hbf17e8c2, 32'h00000000} /* (16, 21, 3) {real, imag} */,
  {32'hbebc6f30, 32'h00000000} /* (16, 21, 2) {real, imag} */,
  {32'hbe2ab8f9, 32'h00000000} /* (16, 21, 1) {real, imag} */,
  {32'hbd72c206, 32'h00000000} /* (16, 21, 0) {real, imag} */,
  {32'h3ed6bfa3, 32'h00000000} /* (16, 20, 31) {real, imag} */,
  {32'h3f2da638, 32'h00000000} /* (16, 20, 30) {real, imag} */,
  {32'h3c4fc048, 32'h00000000} /* (16, 20, 29) {real, imag} */,
  {32'hbe95bd6b, 32'h00000000} /* (16, 20, 28) {real, imag} */,
  {32'hbf109600, 32'h00000000} /* (16, 20, 27) {real, imag} */,
  {32'hbd95318a, 32'h00000000} /* (16, 20, 26) {real, imag} */,
  {32'h3e48ebd4, 32'h00000000} /* (16, 20, 25) {real, imag} */,
  {32'h3f1b18a5, 32'h00000000} /* (16, 20, 24) {real, imag} */,
  {32'h3f0d19e0, 32'h00000000} /* (16, 20, 23) {real, imag} */,
  {32'h3eaa2ad4, 32'h00000000} /* (16, 20, 22) {real, imag} */,
  {32'hbd2ee2bc, 32'h00000000} /* (16, 20, 21) {real, imag} */,
  {32'hbf0ae082, 32'h00000000} /* (16, 20, 20) {real, imag} */,
  {32'hbe99c28a, 32'h00000000} /* (16, 20, 19) {real, imag} */,
  {32'hbe20716b, 32'h00000000} /* (16, 20, 18) {real, imag} */,
  {32'hbe7b6ea5, 32'h00000000} /* (16, 20, 17) {real, imag} */,
  {32'hbed00a12, 32'h00000000} /* (16, 20, 16) {real, imag} */,
  {32'h3eb2279e, 32'h00000000} /* (16, 20, 15) {real, imag} */,
  {32'h3eb932d3, 32'h00000000} /* (16, 20, 14) {real, imag} */,
  {32'hbef2185b, 32'h00000000} /* (16, 20, 13) {real, imag} */,
  {32'hbf70522a, 32'h00000000} /* (16, 20, 12) {real, imag} */,
  {32'hbf2882c5, 32'h00000000} /* (16, 20, 11) {real, imag} */,
  {32'hbe830e6e, 32'h00000000} /* (16, 20, 10) {real, imag} */,
  {32'h3eef151d, 32'h00000000} /* (16, 20, 9) {real, imag} */,
  {32'h3e879f6f, 32'h00000000} /* (16, 20, 8) {real, imag} */,
  {32'h3d8c052e, 32'h00000000} /* (16, 20, 7) {real, imag} */,
  {32'h3e32ea6e, 32'h00000000} /* (16, 20, 6) {real, imag} */,
  {32'h3e90dfa5, 32'h00000000} /* (16, 20, 5) {real, imag} */,
  {32'h3ed2311b, 32'h00000000} /* (16, 20, 4) {real, imag} */,
  {32'h3f17c825, 32'h00000000} /* (16, 20, 3) {real, imag} */,
  {32'h3f371794, 32'h00000000} /* (16, 20, 2) {real, imag} */,
  {32'h3e927e8d, 32'h00000000} /* (16, 20, 1) {real, imag} */,
  {32'h3e2695d2, 32'h00000000} /* (16, 20, 0) {real, imag} */,
  {32'h3e55c2ea, 32'h00000000} /* (16, 19, 31) {real, imag} */,
  {32'h3e913abd, 32'h00000000} /* (16, 19, 30) {real, imag} */,
  {32'h3dddd6f5, 32'h00000000} /* (16, 19, 29) {real, imag} */,
  {32'hbc39116c, 32'h00000000} /* (16, 19, 28) {real, imag} */,
  {32'hbd6a17d3, 32'h00000000} /* (16, 19, 27) {real, imag} */,
  {32'h3eaf24c3, 32'h00000000} /* (16, 19, 26) {real, imag} */,
  {32'h3e29fc35, 32'h00000000} /* (16, 19, 25) {real, imag} */,
  {32'h3f17b9e3, 32'h00000000} /* (16, 19, 24) {real, imag} */,
  {32'h3f95d83a, 32'h00000000} /* (16, 19, 23) {real, imag} */,
  {32'h3f9e8ed9, 32'h00000000} /* (16, 19, 22) {real, imag} */,
  {32'h3f1ff3c0, 32'h00000000} /* (16, 19, 21) {real, imag} */,
  {32'hbeb64f5a, 32'h00000000} /* (16, 19, 20) {real, imag} */,
  {32'hbf40cb52, 32'h00000000} /* (16, 19, 19) {real, imag} */,
  {32'hbe4c4052, 32'h00000000} /* (16, 19, 18) {real, imag} */,
  {32'hbdbeabdc, 32'h00000000} /* (16, 19, 17) {real, imag} */,
  {32'hbf14142d, 32'h00000000} /* (16, 19, 16) {real, imag} */,
  {32'hbf09ca47, 32'h00000000} /* (16, 19, 15) {real, imag} */,
  {32'hbe977968, 32'h00000000} /* (16, 19, 14) {real, imag} */,
  {32'hbeb7c9e5, 32'h00000000} /* (16, 19, 13) {real, imag} */,
  {32'hbed2870e, 32'h00000000} /* (16, 19, 12) {real, imag} */,
  {32'hbf331f24, 32'h00000000} /* (16, 19, 11) {real, imag} */,
  {32'h3e10d8ce, 32'h00000000} /* (16, 19, 10) {real, imag} */,
  {32'h3f4d6dbc, 32'h00000000} /* (16, 19, 9) {real, imag} */,
  {32'h3ec75d9e, 32'h00000000} /* (16, 19, 8) {real, imag} */,
  {32'h3d32bd28, 32'h00000000} /* (16, 19, 7) {real, imag} */,
  {32'h3ea81589, 32'h00000000} /* (16, 19, 6) {real, imag} */,
  {32'h3f413947, 32'h00000000} /* (16, 19, 5) {real, imag} */,
  {32'h3f2644f4, 32'h00000000} /* (16, 19, 4) {real, imag} */,
  {32'h3f1d9d92, 32'h00000000} /* (16, 19, 3) {real, imag} */,
  {32'h3f6cf443, 32'h00000000} /* (16, 19, 2) {real, imag} */,
  {32'h3f905734, 32'h00000000} /* (16, 19, 1) {real, imag} */,
  {32'h3efc588d, 32'h00000000} /* (16, 19, 0) {real, imag} */,
  {32'h3f060975, 32'h00000000} /* (16, 18, 31) {real, imag} */,
  {32'h3ea1e378, 32'h00000000} /* (16, 18, 30) {real, imag} */,
  {32'h3e4dc29c, 32'h00000000} /* (16, 18, 29) {real, imag} */,
  {32'h3e9b5be4, 32'h00000000} /* (16, 18, 28) {real, imag} */,
  {32'h3f42cc28, 32'h00000000} /* (16, 18, 27) {real, imag} */,
  {32'h3f742d91, 32'h00000000} /* (16, 18, 26) {real, imag} */,
  {32'h3f2e2b4d, 32'h00000000} /* (16, 18, 25) {real, imag} */,
  {32'h3fbab57f, 32'h00000000} /* (16, 18, 24) {real, imag} */,
  {32'h3fa81dd8, 32'h00000000} /* (16, 18, 23) {real, imag} */,
  {32'h3f37cf43, 32'h00000000} /* (16, 18, 22) {real, imag} */,
  {32'h3f3d447e, 32'h00000000} /* (16, 18, 21) {real, imag} */,
  {32'hbe057bc3, 32'h00000000} /* (16, 18, 20) {real, imag} */,
  {32'hbf2a9253, 32'h00000000} /* (16, 18, 19) {real, imag} */,
  {32'hbf39cb54, 32'h00000000} /* (16, 18, 18) {real, imag} */,
  {32'hbf65d30d, 32'h00000000} /* (16, 18, 17) {real, imag} */,
  {32'hbf445616, 32'h00000000} /* (16, 18, 16) {real, imag} */,
  {32'hbf3b5130, 32'h00000000} /* (16, 18, 15) {real, imag} */,
  {32'hbef10011, 32'h00000000} /* (16, 18, 14) {real, imag} */,
  {32'hbef9faf3, 32'h00000000} /* (16, 18, 13) {real, imag} */,
  {32'h3d0a55ac, 32'h00000000} /* (16, 18, 12) {real, imag} */,
  {32'hbe42c05d, 32'h00000000} /* (16, 18, 11) {real, imag} */,
  {32'h3f306757, 32'h00000000} /* (16, 18, 10) {real, imag} */,
  {32'h3f90def5, 32'h00000000} /* (16, 18, 9) {real, imag} */,
  {32'h3ef70ef4, 32'h00000000} /* (16, 18, 8) {real, imag} */,
  {32'h3dc08997, 32'h00000000} /* (16, 18, 7) {real, imag} */,
  {32'h3e972d17, 32'h00000000} /* (16, 18, 6) {real, imag} */,
  {32'h3f06f084, 32'h00000000} /* (16, 18, 5) {real, imag} */,
  {32'h3f81acd6, 32'h00000000} /* (16, 18, 4) {real, imag} */,
  {32'h3ec79512, 32'h00000000} /* (16, 18, 3) {real, imag} */,
  {32'h3f1a5fa2, 32'h00000000} /* (16, 18, 2) {real, imag} */,
  {32'h3f9b27c0, 32'h00000000} /* (16, 18, 1) {real, imag} */,
  {32'h3f3b3e2a, 32'h00000000} /* (16, 18, 0) {real, imag} */,
  {32'h3f43debd, 32'h00000000} /* (16, 17, 31) {real, imag} */,
  {32'h3f014dc6, 32'h00000000} /* (16, 17, 30) {real, imag} */,
  {32'h3eb62b84, 32'h00000000} /* (16, 17, 29) {real, imag} */,
  {32'h3f30d945, 32'h00000000} /* (16, 17, 28) {real, imag} */,
  {32'h3f0c99a1, 32'h00000000} /* (16, 17, 27) {real, imag} */,
  {32'h3f23178a, 32'h00000000} /* (16, 17, 26) {real, imag} */,
  {32'h3f88ca2f, 32'h00000000} /* (16, 17, 25) {real, imag} */,
  {32'h3fd1f6a0, 32'h00000000} /* (16, 17, 24) {real, imag} */,
  {32'h3f43308d, 32'h00000000} /* (16, 17, 23) {real, imag} */,
  {32'h3f597f58, 32'h00000000} /* (16, 17, 22) {real, imag} */,
  {32'h3f6e51c9, 32'h00000000} /* (16, 17, 21) {real, imag} */,
  {32'hbe9cc2bc, 32'h00000000} /* (16, 17, 20) {real, imag} */,
  {32'hbf021618, 32'h00000000} /* (16, 17, 19) {real, imag} */,
  {32'hbf24fa85, 32'h00000000} /* (16, 17, 18) {real, imag} */,
  {32'hbf70b067, 32'h00000000} /* (16, 17, 17) {real, imag} */,
  {32'hbf65ca54, 32'h00000000} /* (16, 17, 16) {real, imag} */,
  {32'hbf67e306, 32'h00000000} /* (16, 17, 15) {real, imag} */,
  {32'hbf98001c, 32'h00000000} /* (16, 17, 14) {real, imag} */,
  {32'hbf5f876c, 32'h00000000} /* (16, 17, 13) {real, imag} */,
  {32'hbec1c1a2, 32'h00000000} /* (16, 17, 12) {real, imag} */,
  {32'hbe8f72e8, 32'h00000000} /* (16, 17, 11) {real, imag} */,
  {32'h3f45058b, 32'h00000000} /* (16, 17, 10) {real, imag} */,
  {32'h3fa9e2d7, 32'h00000000} /* (16, 17, 9) {real, imag} */,
  {32'h3f91f31e, 32'h00000000} /* (16, 17, 8) {real, imag} */,
  {32'h3ef7ecd0, 32'h00000000} /* (16, 17, 7) {real, imag} */,
  {32'hbcf22810, 32'h00000000} /* (16, 17, 6) {real, imag} */,
  {32'h3e1054c0, 32'h00000000} /* (16, 17, 5) {real, imag} */,
  {32'h3f3bae7d, 32'h00000000} /* (16, 17, 4) {real, imag} */,
  {32'h3ee2958f, 32'h00000000} /* (16, 17, 3) {real, imag} */,
  {32'h3e019d67, 32'h00000000} /* (16, 17, 2) {real, imag} */,
  {32'h3f00c3ab, 32'h00000000} /* (16, 17, 1) {real, imag} */,
  {32'h3f348603, 32'h00000000} /* (16, 17, 0) {real, imag} */,
  {32'h3e8bdc45, 32'h00000000} /* (16, 16, 31) {real, imag} */,
  {32'h3db6efc2, 32'h00000000} /* (16, 16, 30) {real, imag} */,
  {32'h3f0dd198, 32'h00000000} /* (16, 16, 29) {real, imag} */,
  {32'h3f82f8cf, 32'h00000000} /* (16, 16, 28) {real, imag} */,
  {32'h3f31f3f9, 32'h00000000} /* (16, 16, 27) {real, imag} */,
  {32'h3ea1a4d5, 32'h00000000} /* (16, 16, 26) {real, imag} */,
  {32'h3e932ece, 32'h00000000} /* (16, 16, 25) {real, imag} */,
  {32'h3f33f90b, 32'h00000000} /* (16, 16, 24) {real, imag} */,
  {32'h3f0e8571, 32'h00000000} /* (16, 16, 23) {real, imag} */,
  {32'h3f2310e9, 32'h00000000} /* (16, 16, 22) {real, imag} */,
  {32'h3ebac6f8, 32'h00000000} /* (16, 16, 21) {real, imag} */,
  {32'hbf0e61d1, 32'h00000000} /* (16, 16, 20) {real, imag} */,
  {32'hbf4e825e, 32'h00000000} /* (16, 16, 19) {real, imag} */,
  {32'hbf12e252, 32'h00000000} /* (16, 16, 18) {real, imag} */,
  {32'hbf7f05c9, 32'h00000000} /* (16, 16, 17) {real, imag} */,
  {32'hbf833ffe, 32'h00000000} /* (16, 16, 16) {real, imag} */,
  {32'hbf55cc45, 32'h00000000} /* (16, 16, 15) {real, imag} */,
  {32'hbf938a4c, 32'h00000000} /* (16, 16, 14) {real, imag} */,
  {32'hbf52dd6b, 32'h00000000} /* (16, 16, 13) {real, imag} */,
  {32'hbf8c6c3c, 32'h00000000} /* (16, 16, 12) {real, imag} */,
  {32'hbf28641a, 32'h00000000} /* (16, 16, 11) {real, imag} */,
  {32'h3f01506a, 32'h00000000} /* (16, 16, 10) {real, imag} */,
  {32'h3f39cfbd, 32'h00000000} /* (16, 16, 9) {real, imag} */,
  {32'h3f538b58, 32'h00000000} /* (16, 16, 8) {real, imag} */,
  {32'h3ee74045, 32'h00000000} /* (16, 16, 7) {real, imag} */,
  {32'hbddac106, 32'h00000000} /* (16, 16, 6) {real, imag} */,
  {32'h3e2d9fc8, 32'h00000000} /* (16, 16, 5) {real, imag} */,
  {32'h3ed92e54, 32'h00000000} /* (16, 16, 4) {real, imag} */,
  {32'h3f28cb8c, 32'h00000000} /* (16, 16, 3) {real, imag} */,
  {32'h3f1cfdea, 32'h00000000} /* (16, 16, 2) {real, imag} */,
  {32'h3ecc266e, 32'h00000000} /* (16, 16, 1) {real, imag} */,
  {32'h3e9880a2, 32'h00000000} /* (16, 16, 0) {real, imag} */,
  {32'hbd49f5cf, 32'h00000000} /* (16, 15, 31) {real, imag} */,
  {32'h3d854e5f, 32'h00000000} /* (16, 15, 30) {real, imag} */,
  {32'h3f16167b, 32'h00000000} /* (16, 15, 29) {real, imag} */,
  {32'h3f57488b, 32'h00000000} /* (16, 15, 28) {real, imag} */,
  {32'h3f445247, 32'h00000000} /* (16, 15, 27) {real, imag} */,
  {32'h3ea27e6d, 32'h00000000} /* (16, 15, 26) {real, imag} */,
  {32'hbe265c14, 32'h00000000} /* (16, 15, 25) {real, imag} */,
  {32'hbdecb28d, 32'h00000000} /* (16, 15, 24) {real, imag} */,
  {32'h3ea387d1, 32'h00000000} /* (16, 15, 23) {real, imag} */,
  {32'h3f35f5ff, 32'h00000000} /* (16, 15, 22) {real, imag} */,
  {32'h3eafb6df, 32'h00000000} /* (16, 15, 21) {real, imag} */,
  {32'hbf0626ad, 32'h00000000} /* (16, 15, 20) {real, imag} */,
  {32'hbf3e2c02, 32'h00000000} /* (16, 15, 19) {real, imag} */,
  {32'hbeb9442e, 32'h00000000} /* (16, 15, 18) {real, imag} */,
  {32'hbf20e012, 32'h00000000} /* (16, 15, 17) {real, imag} */,
  {32'hbf1ced92, 32'h00000000} /* (16, 15, 16) {real, imag} */,
  {32'hbf2b7d40, 32'h00000000} /* (16, 15, 15) {real, imag} */,
  {32'hbf370f38, 32'h00000000} /* (16, 15, 14) {real, imag} */,
  {32'hbe8e8060, 32'h00000000} /* (16, 15, 13) {real, imag} */,
  {32'hbe9790ed, 32'h00000000} /* (16, 15, 12) {real, imag} */,
  {32'hbddfe4b9, 32'h00000000} /* (16, 15, 11) {real, imag} */,
  {32'h3f25f641, 32'h00000000} /* (16, 15, 10) {real, imag} */,
  {32'h3f6674e9, 32'h00000000} /* (16, 15, 9) {real, imag} */,
  {32'h3f09e294, 32'h00000000} /* (16, 15, 8) {real, imag} */,
  {32'h3f02ed2d, 32'h00000000} /* (16, 15, 7) {real, imag} */,
  {32'h3e678d43, 32'h00000000} /* (16, 15, 6) {real, imag} */,
  {32'h3e39067b, 32'h00000000} /* (16, 15, 5) {real, imag} */,
  {32'h3f1f89c5, 32'h00000000} /* (16, 15, 4) {real, imag} */,
  {32'h3f680a65, 32'h00000000} /* (16, 15, 3) {real, imag} */,
  {32'h3f35f19c, 32'h00000000} /* (16, 15, 2) {real, imag} */,
  {32'h3eb1c4de, 32'h00000000} /* (16, 15, 1) {real, imag} */,
  {32'h3d41ae22, 32'h00000000} /* (16, 15, 0) {real, imag} */,
  {32'h3d853594, 32'h00000000} /* (16, 14, 31) {real, imag} */,
  {32'h3e5bf74f, 32'h00000000} /* (16, 14, 30) {real, imag} */,
  {32'h3edcf9b0, 32'h00000000} /* (16, 14, 29) {real, imag} */,
  {32'hbc2f64e0, 32'h00000000} /* (16, 14, 28) {real, imag} */,
  {32'h3ed31aa1, 32'h00000000} /* (16, 14, 27) {real, imag} */,
  {32'h3e8536f4, 32'h00000000} /* (16, 14, 26) {real, imag} */,
  {32'hbe25d71b, 32'h00000000} /* (16, 14, 25) {real, imag} */,
  {32'h3ce51463, 32'h00000000} /* (16, 14, 24) {real, imag} */,
  {32'h3eecaa09, 32'h00000000} /* (16, 14, 23) {real, imag} */,
  {32'h3f4c7816, 32'h00000000} /* (16, 14, 22) {real, imag} */,
  {32'h3db0a3ec, 32'h00000000} /* (16, 14, 21) {real, imag} */,
  {32'hbf4bdc0a, 32'h00000000} /* (16, 14, 20) {real, imag} */,
  {32'hbfa31f39, 32'h00000000} /* (16, 14, 19) {real, imag} */,
  {32'hbebc4acb, 32'h00000000} /* (16, 14, 18) {real, imag} */,
  {32'h3d8d1b13, 32'h00000000} /* (16, 14, 17) {real, imag} */,
  {32'hbe1adab0, 32'h00000000} /* (16, 14, 16) {real, imag} */,
  {32'hbe34886a, 32'h00000000} /* (16, 14, 15) {real, imag} */,
  {32'hbef2e739, 32'h00000000} /* (16, 14, 14) {real, imag} */,
  {32'hbeed31a0, 32'h00000000} /* (16, 14, 13) {real, imag} */,
  {32'hbec19816, 32'h00000000} /* (16, 14, 12) {real, imag} */,
  {32'hbe1581b0, 32'h00000000} /* (16, 14, 11) {real, imag} */,
  {32'h3eec9244, 32'h00000000} /* (16, 14, 10) {real, imag} */,
  {32'h3f08c41f, 32'h00000000} /* (16, 14, 9) {real, imag} */,
  {32'h3eac3272, 32'h00000000} /* (16, 14, 8) {real, imag} */,
  {32'h3e661de1, 32'h00000000} /* (16, 14, 7) {real, imag} */,
  {32'h3dedad22, 32'h00000000} /* (16, 14, 6) {real, imag} */,
  {32'h3e4b72eb, 32'h00000000} /* (16, 14, 5) {real, imag} */,
  {32'h3f1ed703, 32'h00000000} /* (16, 14, 4) {real, imag} */,
  {32'h3f5c01e9, 32'h00000000} /* (16, 14, 3) {real, imag} */,
  {32'h3eba2a6e, 32'h00000000} /* (16, 14, 2) {real, imag} */,
  {32'h3daed59d, 32'h00000000} /* (16, 14, 1) {real, imag} */,
  {32'hbd6e768d, 32'h00000000} /* (16, 14, 0) {real, imag} */,
  {32'h3e73eb0c, 32'h00000000} /* (16, 13, 31) {real, imag} */,
  {32'h3ef1f0f9, 32'h00000000} /* (16, 13, 30) {real, imag} */,
  {32'h3f4488e4, 32'h00000000} /* (16, 13, 29) {real, imag} */,
  {32'h3e993e97, 32'h00000000} /* (16, 13, 28) {real, imag} */,
  {32'h3f00ac47, 32'h00000000} /* (16, 13, 27) {real, imag} */,
  {32'h3f58fd20, 32'h00000000} /* (16, 13, 26) {real, imag} */,
  {32'h3f3395ff, 32'h00000000} /* (16, 13, 25) {real, imag} */,
  {32'h3edf5aa2, 32'h00000000} /* (16, 13, 24) {real, imag} */,
  {32'h3e5612ce, 32'h00000000} /* (16, 13, 23) {real, imag} */,
  {32'h3e6bcae2, 32'h00000000} /* (16, 13, 22) {real, imag} */,
  {32'hbe371e82, 32'h00000000} /* (16, 13, 21) {real, imag} */,
  {32'hbf5dbcd6, 32'h00000000} /* (16, 13, 20) {real, imag} */,
  {32'hbf63b1fa, 32'h00000000} /* (16, 13, 19) {real, imag} */,
  {32'hbed96717, 32'h00000000} /* (16, 13, 18) {real, imag} */,
  {32'hbe30c872, 32'h00000000} /* (16, 13, 17) {real, imag} */,
  {32'hbda22afc, 32'h00000000} /* (16, 13, 16) {real, imag} */,
  {32'hbe58fb73, 32'h00000000} /* (16, 13, 15) {real, imag} */,
  {32'hbedb2069, 32'h00000000} /* (16, 13, 14) {real, imag} */,
  {32'hbef8566c, 32'h00000000} /* (16, 13, 13) {real, imag} */,
  {32'hbef63a47, 32'h00000000} /* (16, 13, 12) {real, imag} */,
  {32'hbef534d9, 32'h00000000} /* (16, 13, 11) {real, imag} */,
  {32'h3e6989da, 32'h00000000} /* (16, 13, 10) {real, imag} */,
  {32'h3f02949b, 32'h00000000} /* (16, 13, 9) {real, imag} */,
  {32'h3f4293e9, 32'h00000000} /* (16, 13, 8) {real, imag} */,
  {32'h3f006f2b, 32'h00000000} /* (16, 13, 7) {real, imag} */,
  {32'h3deded9c, 32'h00000000} /* (16, 13, 6) {real, imag} */,
  {32'h3e78347c, 32'h00000000} /* (16, 13, 5) {real, imag} */,
  {32'h3f3d6a62, 32'h00000000} /* (16, 13, 4) {real, imag} */,
  {32'h3fa04d33, 32'h00000000} /* (16, 13, 3) {real, imag} */,
  {32'h3f4e8d29, 32'h00000000} /* (16, 13, 2) {real, imag} */,
  {32'h3eb562a9, 32'h00000000} /* (16, 13, 1) {real, imag} */,
  {32'hbd048582, 32'h00000000} /* (16, 13, 0) {real, imag} */,
  {32'h3e8dbe48, 32'h00000000} /* (16, 12, 31) {real, imag} */,
  {32'h3eecf984, 32'h00000000} /* (16, 12, 30) {real, imag} */,
  {32'h3f5e01d0, 32'h00000000} /* (16, 12, 29) {real, imag} */,
  {32'h3f385a3e, 32'h00000000} /* (16, 12, 28) {real, imag} */,
  {32'h3f6c11dd, 32'h00000000} /* (16, 12, 27) {real, imag} */,
  {32'h3f86b6d9, 32'h00000000} /* (16, 12, 26) {real, imag} */,
  {32'h3f84c6f5, 32'h00000000} /* (16, 12, 25) {real, imag} */,
  {32'h3f6397d7, 32'h00000000} /* (16, 12, 24) {real, imag} */,
  {32'h3f1510fa, 32'h00000000} /* (16, 12, 23) {real, imag} */,
  {32'h3f1c8ffe, 32'h00000000} /* (16, 12, 22) {real, imag} */,
  {32'h3f4c7159, 32'h00000000} /* (16, 12, 21) {real, imag} */,
  {32'hbea12fdc, 32'h00000000} /* (16, 12, 20) {real, imag} */,
  {32'hbf84768d, 32'h00000000} /* (16, 12, 19) {real, imag} */,
  {32'hbf2fc025, 32'h00000000} /* (16, 12, 18) {real, imag} */,
  {32'hbe041776, 32'h00000000} /* (16, 12, 17) {real, imag} */,
  {32'hbee99dec, 32'h00000000} /* (16, 12, 16) {real, imag} */,
  {32'hbf822534, 32'h00000000} /* (16, 12, 15) {real, imag} */,
  {32'hbf3378ba, 32'h00000000} /* (16, 12, 14) {real, imag} */,
  {32'hbdf27ed7, 32'h00000000} /* (16, 12, 13) {real, imag} */,
  {32'hbe81837d, 32'h00000000} /* (16, 12, 12) {real, imag} */,
  {32'h3c82af28, 32'h00000000} /* (16, 12, 11) {real, imag} */,
  {32'h3ec76708, 32'h00000000} /* (16, 12, 10) {real, imag} */,
  {32'h3f14aaad, 32'h00000000} /* (16, 12, 9) {real, imag} */,
  {32'h3f099b10, 32'h00000000} /* (16, 12, 8) {real, imag} */,
  {32'h3f1d4e54, 32'h00000000} /* (16, 12, 7) {real, imag} */,
  {32'h3f4de33f, 32'h00000000} /* (16, 12, 6) {real, imag} */,
  {32'h3f0547a4, 32'h00000000} /* (16, 12, 5) {real, imag} */,
  {32'h3f30fb6c, 32'h00000000} /* (16, 12, 4) {real, imag} */,
  {32'h3f5db64b, 32'h00000000} /* (16, 12, 3) {real, imag} */,
  {32'h3f97c5b7, 32'h00000000} /* (16, 12, 2) {real, imag} */,
  {32'h3f64a372, 32'h00000000} /* (16, 12, 1) {real, imag} */,
  {32'h3ed62e8b, 32'h00000000} /* (16, 12, 0) {real, imag} */,
  {32'h3ec406b4, 32'h00000000} /* (16, 11, 31) {real, imag} */,
  {32'h3f54560a, 32'h00000000} /* (16, 11, 30) {real, imag} */,
  {32'h3f2ce4ae, 32'h00000000} /* (16, 11, 29) {real, imag} */,
  {32'h3f2bd4f0, 32'h00000000} /* (16, 11, 28) {real, imag} */,
  {32'h3f290364, 32'h00000000} /* (16, 11, 27) {real, imag} */,
  {32'h3e47f02c, 32'h00000000} /* (16, 11, 26) {real, imag} */,
  {32'h3e18f4be, 32'h00000000} /* (16, 11, 25) {real, imag} */,
  {32'h3ee59b5d, 32'h00000000} /* (16, 11, 24) {real, imag} */,
  {32'h3e8a110e, 32'h00000000} /* (16, 11, 23) {real, imag} */,
  {32'h3f16ca1a, 32'h00000000} /* (16, 11, 22) {real, imag} */,
  {32'h3f8d7f33, 32'h00000000} /* (16, 11, 21) {real, imag} */,
  {32'h3bfff469, 32'h00000000} /* (16, 11, 20) {real, imag} */,
  {32'hbf49a917, 32'h00000000} /* (16, 11, 19) {real, imag} */,
  {32'hbeacd162, 32'h00000000} /* (16, 11, 18) {real, imag} */,
  {32'h3d19bc44, 32'h00000000} /* (16, 11, 17) {real, imag} */,
  {32'hbee1355d, 32'h00000000} /* (16, 11, 16) {real, imag} */,
  {32'hbf37a16d, 32'h00000000} /* (16, 11, 15) {real, imag} */,
  {32'hbe3afb16, 32'h00000000} /* (16, 11, 14) {real, imag} */,
  {32'h3c9fe1eb, 32'h00000000} /* (16, 11, 13) {real, imag} */,
  {32'hbe626356, 32'h00000000} /* (16, 11, 12) {real, imag} */,
  {32'h3dd98083, 32'h00000000} /* (16, 11, 11) {real, imag} */,
  {32'h3e0d669a, 32'h00000000} /* (16, 11, 10) {real, imag} */,
  {32'h3f3433ca, 32'h00000000} /* (16, 11, 9) {real, imag} */,
  {32'h3f911aa2, 32'h00000000} /* (16, 11, 8) {real, imag} */,
  {32'h3f114b70, 32'h00000000} /* (16, 11, 7) {real, imag} */,
  {32'h3f9f245d, 32'h00000000} /* (16, 11, 6) {real, imag} */,
  {32'h3fab0db6, 32'h00000000} /* (16, 11, 5) {real, imag} */,
  {32'h3f3778ec, 32'h00000000} /* (16, 11, 4) {real, imag} */,
  {32'h3edaa7de, 32'h00000000} /* (16, 11, 3) {real, imag} */,
  {32'h3f079e91, 32'h00000000} /* (16, 11, 2) {real, imag} */,
  {32'h3f271e4b, 32'h00000000} /* (16, 11, 1) {real, imag} */,
  {32'h3f28f8cb, 32'h00000000} /* (16, 11, 0) {real, imag} */,
  {32'hbe894c22, 32'h00000000} /* (16, 10, 31) {real, imag} */,
  {32'h3d2d698a, 32'h00000000} /* (16, 10, 30) {real, imag} */,
  {32'h3e436a12, 32'h00000000} /* (16, 10, 29) {real, imag} */,
  {32'h3d5398a0, 32'h00000000} /* (16, 10, 28) {real, imag} */,
  {32'hbf074bab, 32'h00000000} /* (16, 10, 27) {real, imag} */,
  {32'hbf233040, 32'h00000000} /* (16, 10, 26) {real, imag} */,
  {32'hbec7e1aa, 32'h00000000} /* (16, 10, 25) {real, imag} */,
  {32'hbeac7bad, 32'h00000000} /* (16, 10, 24) {real, imag} */,
  {32'hbed27073, 32'h00000000} /* (16, 10, 23) {real, imag} */,
  {32'hbe1514b8, 32'h00000000} /* (16, 10, 22) {real, imag} */,
  {32'hbe064907, 32'h00000000} /* (16, 10, 21) {real, imag} */,
  {32'h3e4a8c17, 32'h00000000} /* (16, 10, 20) {real, imag} */,
  {32'h3e6f0281, 32'h00000000} /* (16, 10, 19) {real, imag} */,
  {32'h3f04053e, 32'h00000000} /* (16, 10, 18) {real, imag} */,
  {32'h3ecde400, 32'h00000000} /* (16, 10, 17) {real, imag} */,
  {32'h3ede743f, 32'h00000000} /* (16, 10, 16) {real, imag} */,
  {32'h3f423b76, 32'h00000000} /* (16, 10, 15) {real, imag} */,
  {32'h3e973067, 32'h00000000} /* (16, 10, 14) {real, imag} */,
  {32'h3e661a8b, 32'h00000000} /* (16, 10, 13) {real, imag} */,
  {32'h3e4435c3, 32'h00000000} /* (16, 10, 12) {real, imag} */,
  {32'h3d3e991b, 32'h00000000} /* (16, 10, 11) {real, imag} */,
  {32'hbdef557c, 32'h00000000} /* (16, 10, 10) {real, imag} */,
  {32'hbe0020ea, 32'h00000000} /* (16, 10, 9) {real, imag} */,
  {32'h3e37c83f, 32'h00000000} /* (16, 10, 8) {real, imag} */,
  {32'hbde9b9a8, 32'h00000000} /* (16, 10, 7) {real, imag} */,
  {32'h3f0718cc, 32'h00000000} /* (16, 10, 6) {real, imag} */,
  {32'h3ee2bd16, 32'h00000000} /* (16, 10, 5) {real, imag} */,
  {32'hbdbd7788, 32'h00000000} /* (16, 10, 4) {real, imag} */,
  {32'hbd2c03ea, 32'h00000000} /* (16, 10, 3) {real, imag} */,
  {32'hbdfcf430, 32'h00000000} /* (16, 10, 2) {real, imag} */,
  {32'hbd18686f, 32'h00000000} /* (16, 10, 1) {real, imag} */,
  {32'h3db0356c, 32'h00000000} /* (16, 10, 0) {real, imag} */,
  {32'hbebc9284, 32'h00000000} /* (16, 9, 31) {real, imag} */,
  {32'hbf375089, 32'h00000000} /* (16, 9, 30) {real, imag} */,
  {32'hbea57f66, 32'h00000000} /* (16, 9, 29) {real, imag} */,
  {32'hbe0f4de4, 32'h00000000} /* (16, 9, 28) {real, imag} */,
  {32'hbf513a0c, 32'h00000000} /* (16, 9, 27) {real, imag} */,
  {32'hbeb58b2e, 32'h00000000} /* (16, 9, 26) {real, imag} */,
  {32'hbe74ec9e, 32'h00000000} /* (16, 9, 25) {real, imag} */,
  {32'hbe8f0ad0, 32'h00000000} /* (16, 9, 24) {real, imag} */,
  {32'hbf24cda2, 32'h00000000} /* (16, 9, 23) {real, imag} */,
  {32'hbf645416, 32'h00000000} /* (16, 9, 22) {real, imag} */,
  {32'hbedf4533, 32'h00000000} /* (16, 9, 21) {real, imag} */,
  {32'h3e967473, 32'h00000000} /* (16, 9, 20) {real, imag} */,
  {32'h3f3c38ca, 32'h00000000} /* (16, 9, 19) {real, imag} */,
  {32'h3f341d8e, 32'h00000000} /* (16, 9, 18) {real, imag} */,
  {32'h3f758693, 32'h00000000} /* (16, 9, 17) {real, imag} */,
  {32'h3fa53d05, 32'h00000000} /* (16, 9, 16) {real, imag} */,
  {32'h3f9bfe67, 32'h00000000} /* (16, 9, 15) {real, imag} */,
  {32'h3f46d543, 32'h00000000} /* (16, 9, 14) {real, imag} */,
  {32'h3eb57c7e, 32'h00000000} /* (16, 9, 13) {real, imag} */,
  {32'h3eb78467, 32'h00000000} /* (16, 9, 12) {real, imag} */,
  {32'h3e30b034, 32'h00000000} /* (16, 9, 11) {real, imag} */,
  {32'hbeb46994, 32'h00000000} /* (16, 9, 10) {real, imag} */,
  {32'hbf24e006, 32'h00000000} /* (16, 9, 9) {real, imag} */,
  {32'hbf36a78e, 32'h00000000} /* (16, 9, 8) {real, imag} */,
  {32'hbf01b07c, 32'h00000000} /* (16, 9, 7) {real, imag} */,
  {32'hbbdce3b0, 32'h00000000} /* (16, 9, 6) {real, imag} */,
  {32'hbf4e294e, 32'h00000000} /* (16, 9, 5) {real, imag} */,
  {32'hbee3fe54, 32'h00000000} /* (16, 9, 4) {real, imag} */,
  {32'hbd35c1c4, 32'h00000000} /* (16, 9, 3) {real, imag} */,
  {32'hbe9633f6, 32'h00000000} /* (16, 9, 2) {real, imag} */,
  {32'hbeb3f1c3, 32'h00000000} /* (16, 9, 1) {real, imag} */,
  {32'hbebf530e, 32'h00000000} /* (16, 9, 0) {real, imag} */,
  {32'hbee38060, 32'h00000000} /* (16, 8, 31) {real, imag} */,
  {32'hbebdf1a4, 32'h00000000} /* (16, 8, 30) {real, imag} */,
  {32'hbe5ec9a2, 32'h00000000} /* (16, 8, 29) {real, imag} */,
  {32'h3d57c092, 32'h00000000} /* (16, 8, 28) {real, imag} */,
  {32'hbde5e083, 32'h00000000} /* (16, 8, 27) {real, imag} */,
  {32'hbe9ca662, 32'h00000000} /* (16, 8, 26) {real, imag} */,
  {32'hbede6fab, 32'h00000000} /* (16, 8, 25) {real, imag} */,
  {32'hbe3827a7, 32'h00000000} /* (16, 8, 24) {real, imag} */,
  {32'hbf2b3642, 32'h00000000} /* (16, 8, 23) {real, imag} */,
  {32'hbf29570d, 32'h00000000} /* (16, 8, 22) {real, imag} */,
  {32'hbe695c42, 32'h00000000} /* (16, 8, 21) {real, imag} */,
  {32'hbd352052, 32'h00000000} /* (16, 8, 20) {real, imag} */,
  {32'h3f47cf8e, 32'h00000000} /* (16, 8, 19) {real, imag} */,
  {32'h3f0288a3, 32'h00000000} /* (16, 8, 18) {real, imag} */,
  {32'h3f7991d2, 32'h00000000} /* (16, 8, 17) {real, imag} */,
  {32'h3fb15c8e, 32'h00000000} /* (16, 8, 16) {real, imag} */,
  {32'h3f222483, 32'h00000000} /* (16, 8, 15) {real, imag} */,
  {32'h3f69aa7c, 32'h00000000} /* (16, 8, 14) {real, imag} */,
  {32'h3f4cc550, 32'h00000000} /* (16, 8, 13) {real, imag} */,
  {32'h3ee18478, 32'h00000000} /* (16, 8, 12) {real, imag} */,
  {32'h3e0b9150, 32'h00000000} /* (16, 8, 11) {real, imag} */,
  {32'hbeecd5bb, 32'h00000000} /* (16, 8, 10) {real, imag} */,
  {32'hbf18fba4, 32'h00000000} /* (16, 8, 9) {real, imag} */,
  {32'hbe860a88, 32'h00000000} /* (16, 8, 8) {real, imag} */,
  {32'hbe431677, 32'h00000000} /* (16, 8, 7) {real, imag} */,
  {32'hbe4a8074, 32'h00000000} /* (16, 8, 6) {real, imag} */,
  {32'hbf8a8588, 32'h00000000} /* (16, 8, 5) {real, imag} */,
  {32'hbf284bde, 32'h00000000} /* (16, 8, 4) {real, imag} */,
  {32'hbc9f1950, 32'h00000000} /* (16, 8, 3) {real, imag} */,
  {32'hbf0f9434, 32'h00000000} /* (16, 8, 2) {real, imag} */,
  {32'hbf93d520, 32'h00000000} /* (16, 8, 1) {real, imag} */,
  {32'hbf8954b0, 32'h00000000} /* (16, 8, 0) {real, imag} */,
  {32'hbf059ca0, 32'h00000000} /* (16, 7, 31) {real, imag} */,
  {32'hbf0a0930, 32'h00000000} /* (16, 7, 30) {real, imag} */,
  {32'hbe84ce37, 32'h00000000} /* (16, 7, 29) {real, imag} */,
  {32'hbe5ad021, 32'h00000000} /* (16, 7, 28) {real, imag} */,
  {32'hbe9a2319, 32'h00000000} /* (16, 7, 27) {real, imag} */,
  {32'hbf105a96, 32'h00000000} /* (16, 7, 26) {real, imag} */,
  {32'hbf51aa7b, 32'h00000000} /* (16, 7, 25) {real, imag} */,
  {32'hbf030c8b, 32'h00000000} /* (16, 7, 24) {real, imag} */,
  {32'hbf218685, 32'h00000000} /* (16, 7, 23) {real, imag} */,
  {32'hbf2a9e95, 32'h00000000} /* (16, 7, 22) {real, imag} */,
  {32'hbefdc722, 32'h00000000} /* (16, 7, 21) {real, imag} */,
  {32'hbe3702f6, 32'h00000000} /* (16, 7, 20) {real, imag} */,
  {32'h3e9a57fc, 32'h00000000} /* (16, 7, 19) {real, imag} */,
  {32'h3ea1ceb3, 32'h00000000} /* (16, 7, 18) {real, imag} */,
  {32'h3f4a346e, 32'h00000000} /* (16, 7, 17) {real, imag} */,
  {32'h3eae630f, 32'h00000000} /* (16, 7, 16) {real, imag} */,
  {32'hbdb83b90, 32'h00000000} /* (16, 7, 15) {real, imag} */,
  {32'h3f4904bd, 32'h00000000} /* (16, 7, 14) {real, imag} */,
  {32'h3f84bff4, 32'h00000000} /* (16, 7, 13) {real, imag} */,
  {32'h3f0e84ef, 32'h00000000} /* (16, 7, 12) {real, imag} */,
  {32'h3f7e39b2, 32'h00000000} /* (16, 7, 11) {real, imag} */,
  {32'hbe8faa5f, 32'h00000000} /* (16, 7, 10) {real, imag} */,
  {32'hbf73b6a3, 32'h00000000} /* (16, 7, 9) {real, imag} */,
  {32'hbe9b1133, 32'h00000000} /* (16, 7, 8) {real, imag} */,
  {32'hbdb85dc8, 32'h00000000} /* (16, 7, 7) {real, imag} */,
  {32'hbf36c8aa, 32'h00000000} /* (16, 7, 6) {real, imag} */,
  {32'hbf181297, 32'h00000000} /* (16, 7, 5) {real, imag} */,
  {32'hbf6259d9, 32'h00000000} /* (16, 7, 4) {real, imag} */,
  {32'hbeef169c, 32'h00000000} /* (16, 7, 3) {real, imag} */,
  {32'hbf3dbe91, 32'h00000000} /* (16, 7, 2) {real, imag} */,
  {32'hbf5bf729, 32'h00000000} /* (16, 7, 1) {real, imag} */,
  {32'hbeed9b27, 32'h00000000} /* (16, 7, 0) {real, imag} */,
  {32'hbe5a30af, 32'h00000000} /* (16, 6, 31) {real, imag} */,
  {32'hbee85126, 32'h00000000} /* (16, 6, 30) {real, imag} */,
  {32'hbf5283ff, 32'h00000000} /* (16, 6, 29) {real, imag} */,
  {32'hbf315184, 32'h00000000} /* (16, 6, 28) {real, imag} */,
  {32'hbea84bfe, 32'h00000000} /* (16, 6, 27) {real, imag} */,
  {32'hbf2106d0, 32'h00000000} /* (16, 6, 26) {real, imag} */,
  {32'hbf4b94eb, 32'h00000000} /* (16, 6, 25) {real, imag} */,
  {32'hbef3ccb1, 32'h00000000} /* (16, 6, 24) {real, imag} */,
  {32'hbedfb88e, 32'h00000000} /* (16, 6, 23) {real, imag} */,
  {32'hbf1d572f, 32'h00000000} /* (16, 6, 22) {real, imag} */,
  {32'hbf1475d6, 32'h00000000} /* (16, 6, 21) {real, imag} */,
  {32'h3ea04609, 32'h00000000} /* (16, 6, 20) {real, imag} */,
  {32'h3f305120, 32'h00000000} /* (16, 6, 19) {real, imag} */,
  {32'h3ef182a7, 32'h00000000} /* (16, 6, 18) {real, imag} */,
  {32'h3f029fb3, 32'h00000000} /* (16, 6, 17) {real, imag} */,
  {32'h3f16101d, 32'h00000000} /* (16, 6, 16) {real, imag} */,
  {32'h3f11dd85, 32'h00000000} /* (16, 6, 15) {real, imag} */,
  {32'h3f222360, 32'h00000000} /* (16, 6, 14) {real, imag} */,
  {32'h3f51b3de, 32'h00000000} /* (16, 6, 13) {real, imag} */,
  {32'h3e960a27, 32'h00000000} /* (16, 6, 12) {real, imag} */,
  {32'h3f4d1251, 32'h00000000} /* (16, 6, 11) {real, imag} */,
  {32'h3db050d4, 32'h00000000} /* (16, 6, 10) {real, imag} */,
  {32'hbf672947, 32'h00000000} /* (16, 6, 9) {real, imag} */,
  {32'hbe81d088, 32'h00000000} /* (16, 6, 8) {real, imag} */,
  {32'hbe540046, 32'h00000000} /* (16, 6, 7) {real, imag} */,
  {32'hbf153850, 32'h00000000} /* (16, 6, 6) {real, imag} */,
  {32'hbdda264c, 32'h00000000} /* (16, 6, 5) {real, imag} */,
  {32'hbee8589e, 32'h00000000} /* (16, 6, 4) {real, imag} */,
  {32'hbf3e585e, 32'h00000000} /* (16, 6, 3) {real, imag} */,
  {32'hbf7d4714, 32'h00000000} /* (16, 6, 2) {real, imag} */,
  {32'hbf7f70de, 32'h00000000} /* (16, 6, 1) {real, imag} */,
  {32'hbe9091e8, 32'h00000000} /* (16, 6, 0) {real, imag} */,
  {32'hbe0b9900, 32'h00000000} /* (16, 5, 31) {real, imag} */,
  {32'hbf2dce46, 32'h00000000} /* (16, 5, 30) {real, imag} */,
  {32'hbf7f358b, 32'h00000000} /* (16, 5, 29) {real, imag} */,
  {32'hbf2f9a1a, 32'h00000000} /* (16, 5, 28) {real, imag} */,
  {32'hbed8d49d, 32'h00000000} /* (16, 5, 27) {real, imag} */,
  {32'hbf3768c8, 32'h00000000} /* (16, 5, 26) {real, imag} */,
  {32'hbed284ec, 32'h00000000} /* (16, 5, 25) {real, imag} */,
  {32'hbe1df807, 32'h00000000} /* (16, 5, 24) {real, imag} */,
  {32'hbee05813, 32'h00000000} /* (16, 5, 23) {real, imag} */,
  {32'hbf136c2a, 32'h00000000} /* (16, 5, 22) {real, imag} */,
  {32'hbf6f2a00, 32'h00000000} /* (16, 5, 21) {real, imag} */,
  {32'hbeb43d9a, 32'h00000000} /* (16, 5, 20) {real, imag} */,
  {32'h3e9ace19, 32'h00000000} /* (16, 5, 19) {real, imag} */,
  {32'h3df8c8af, 32'h00000000} /* (16, 5, 18) {real, imag} */,
  {32'hbd8cec10, 32'h00000000} /* (16, 5, 17) {real, imag} */,
  {32'h3dacdf79, 32'h00000000} /* (16, 5, 16) {real, imag} */,
  {32'h3ed2b564, 32'h00000000} /* (16, 5, 15) {real, imag} */,
  {32'h3f526d87, 32'h00000000} /* (16, 5, 14) {real, imag} */,
  {32'h3f36fc68, 32'h00000000} /* (16, 5, 13) {real, imag} */,
  {32'h3e6217a7, 32'h00000000} /* (16, 5, 12) {real, imag} */,
  {32'h3e4116ec, 32'h00000000} /* (16, 5, 11) {real, imag} */,
  {32'h3e9ea598, 32'h00000000} /* (16, 5, 10) {real, imag} */,
  {32'h3f011973, 32'h00000000} /* (16, 5, 9) {real, imag} */,
  {32'h3f37c4ce, 32'h00000000} /* (16, 5, 8) {real, imag} */,
  {32'h3ecb3ca0, 32'h00000000} /* (16, 5, 7) {real, imag} */,
  {32'h3ea93ab2, 32'h00000000} /* (16, 5, 6) {real, imag} */,
  {32'h3ccc6c80, 32'h00000000} /* (16, 5, 5) {real, imag} */,
  {32'hbef3c86b, 32'h00000000} /* (16, 5, 4) {real, imag} */,
  {32'hbf9301a6, 32'h00000000} /* (16, 5, 3) {real, imag} */,
  {32'hbfbbc8a8, 32'h00000000} /* (16, 5, 2) {real, imag} */,
  {32'hbf704fa2, 32'h00000000} /* (16, 5, 1) {real, imag} */,
  {32'hbeb74501, 32'h00000000} /* (16, 5, 0) {real, imag} */,
  {32'hbdbb3578, 32'h00000000} /* (16, 4, 31) {real, imag} */,
  {32'hbf2b51a2, 32'h00000000} /* (16, 4, 30) {real, imag} */,
  {32'hbf888f8f, 32'h00000000} /* (16, 4, 29) {real, imag} */,
  {32'hbf03a93d, 32'h00000000} /* (16, 4, 28) {real, imag} */,
  {32'hbe8eaf8d, 32'h00000000} /* (16, 4, 27) {real, imag} */,
  {32'hbe9030cd, 32'h00000000} /* (16, 4, 26) {real, imag} */,
  {32'hbe4d8cba, 32'h00000000} /* (16, 4, 25) {real, imag} */,
  {32'hbd6df900, 32'h00000000} /* (16, 4, 24) {real, imag} */,
  {32'hbd2d936e, 32'h00000000} /* (16, 4, 23) {real, imag} */,
  {32'hbcfd2ed0, 32'h00000000} /* (16, 4, 22) {real, imag} */,
  {32'hbf32d1ff, 32'h00000000} /* (16, 4, 21) {real, imag} */,
  {32'hbfa873bd, 32'h00000000} /* (16, 4, 20) {real, imag} */,
  {32'hbf0357f7, 32'h00000000} /* (16, 4, 19) {real, imag} */,
  {32'hbe7a7e32, 32'h00000000} /* (16, 4, 18) {real, imag} */,
  {32'hbf28a453, 32'h00000000} /* (16, 4, 17) {real, imag} */,
  {32'hbf714359, 32'h00000000} /* (16, 4, 16) {real, imag} */,
  {32'hbe8e9891, 32'h00000000} /* (16, 4, 15) {real, imag} */,
  {32'h3f5e823a, 32'h00000000} /* (16, 4, 14) {real, imag} */,
  {32'h3f1a6ca0, 32'h00000000} /* (16, 4, 13) {real, imag} */,
  {32'h3edcd6a0, 32'h00000000} /* (16, 4, 12) {real, imag} */,
  {32'h3f1035bb, 32'h00000000} /* (16, 4, 11) {real, imag} */,
  {32'h3ef15a14, 32'h00000000} /* (16, 4, 10) {real, imag} */,
  {32'h3f774317, 32'h00000000} /* (16, 4, 9) {real, imag} */,
  {32'h3f9daeca, 32'h00000000} /* (16, 4, 8) {real, imag} */,
  {32'h3f467c11, 32'h00000000} /* (16, 4, 7) {real, imag} */,
  {32'h3f87faa5, 32'h00000000} /* (16, 4, 6) {real, imag} */,
  {32'h3ec8a710, 32'h00000000} /* (16, 4, 5) {real, imag} */,
  {32'hbf4fae45, 32'h00000000} /* (16, 4, 4) {real, imag} */,
  {32'hbf744c62, 32'h00000000} /* (16, 4, 3) {real, imag} */,
  {32'hbf7793e4, 32'h00000000} /* (16, 4, 2) {real, imag} */,
  {32'hbeebe514, 32'h00000000} /* (16, 4, 1) {real, imag} */,
  {32'hbeb53151, 32'h00000000} /* (16, 4, 0) {real, imag} */,
  {32'hbdf56eb8, 32'h00000000} /* (16, 3, 31) {real, imag} */,
  {32'hbf66c983, 32'h00000000} /* (16, 3, 30) {real, imag} */,
  {32'hbf7d5344, 32'h00000000} /* (16, 3, 29) {real, imag} */,
  {32'hbe915f51, 32'h00000000} /* (16, 3, 28) {real, imag} */,
  {32'hbeda9bbb, 32'h00000000} /* (16, 3, 27) {real, imag} */,
  {32'hbecb3de2, 32'h00000000} /* (16, 3, 26) {real, imag} */,
  {32'hbeee50ae, 32'h00000000} /* (16, 3, 25) {real, imag} */,
  {32'hbf074ddd, 32'h00000000} /* (16, 3, 24) {real, imag} */,
  {32'hbeb3fedd, 32'h00000000} /* (16, 3, 23) {real, imag} */,
  {32'hbeec7f62, 32'h00000000} /* (16, 3, 22) {real, imag} */,
  {32'hbf3647e7, 32'h00000000} /* (16, 3, 21) {real, imag} */,
  {32'hbf2b9f4f, 32'h00000000} /* (16, 3, 20) {real, imag} */,
  {32'hbeaa34fa, 32'h00000000} /* (16, 3, 19) {real, imag} */,
  {32'hbf849031, 32'h00000000} /* (16, 3, 18) {real, imag} */,
  {32'hbf5f8277, 32'h00000000} /* (16, 3, 17) {real, imag} */,
  {32'hbedceb09, 32'h00000000} /* (16, 3, 16) {real, imag} */,
  {32'h3e2c6e7d, 32'h00000000} /* (16, 3, 15) {real, imag} */,
  {32'h3f4aa3bc, 32'h00000000} /* (16, 3, 14) {real, imag} */,
  {32'h3f077c98, 32'h00000000} /* (16, 3, 13) {real, imag} */,
  {32'h3ef3f6e4, 32'h00000000} /* (16, 3, 12) {real, imag} */,
  {32'h3f585350, 32'h00000000} /* (16, 3, 11) {real, imag} */,
  {32'h3f3149f5, 32'h00000000} /* (16, 3, 10) {real, imag} */,
  {32'h3f42c0f4, 32'h00000000} /* (16, 3, 9) {real, imag} */,
  {32'h3f814f53, 32'h00000000} /* (16, 3, 8) {real, imag} */,
  {32'h3f0a94b9, 32'h00000000} /* (16, 3, 7) {real, imag} */,
  {32'h3f3cc17e, 32'h00000000} /* (16, 3, 6) {real, imag} */,
  {32'h3e1b02d7, 32'h00000000} /* (16, 3, 5) {real, imag} */,
  {32'hbe915ddf, 32'h00000000} /* (16, 3, 4) {real, imag} */,
  {32'hbc09ad1c, 32'h00000000} /* (16, 3, 3) {real, imag} */,
  {32'hbe95d218, 32'h00000000} /* (16, 3, 2) {real, imag} */,
  {32'hbddaa1d1, 32'h00000000} /* (16, 3, 1) {real, imag} */,
  {32'hbce562a9, 32'h00000000} /* (16, 3, 0) {real, imag} */,
  {32'hbbe98523, 32'h00000000} /* (16, 2, 31) {real, imag} */,
  {32'hbe1bd207, 32'h00000000} /* (16, 2, 30) {real, imag} */,
  {32'hbeafdb30, 32'h00000000} /* (16, 2, 29) {real, imag} */,
  {32'hbee05180, 32'h00000000} /* (16, 2, 28) {real, imag} */,
  {32'hbf060e98, 32'h00000000} /* (16, 2, 27) {real, imag} */,
  {32'hbf7b5efd, 32'h00000000} /* (16, 2, 26) {real, imag} */,
  {32'hbf6e70c2, 32'h00000000} /* (16, 2, 25) {real, imag} */,
  {32'hbf137a0d, 32'h00000000} /* (16, 2, 24) {real, imag} */,
  {32'hbe54b7b5, 32'h00000000} /* (16, 2, 23) {real, imag} */,
  {32'hbef508ea, 32'h00000000} /* (16, 2, 22) {real, imag} */,
  {32'hbf2d54cd, 32'h00000000} /* (16, 2, 21) {real, imag} */,
  {32'hbe77c0be, 32'h00000000} /* (16, 2, 20) {real, imag} */,
  {32'hbee82489, 32'h00000000} /* (16, 2, 19) {real, imag} */,
  {32'hbfc16872, 32'h00000000} /* (16, 2, 18) {real, imag} */,
  {32'hbf872b1c, 32'h00000000} /* (16, 2, 17) {real, imag} */,
  {32'h3e8d80df, 32'h00000000} /* (16, 2, 16) {real, imag} */,
  {32'h3f14a911, 32'h00000000} /* (16, 2, 15) {real, imag} */,
  {32'h3f319df9, 32'h00000000} /* (16, 2, 14) {real, imag} */,
  {32'h3f7a0a84, 32'h00000000} /* (16, 2, 13) {real, imag} */,
  {32'h3f446865, 32'h00000000} /* (16, 2, 12) {real, imag} */,
  {32'h3f1434f6, 32'h00000000} /* (16, 2, 11) {real, imag} */,
  {32'h3f2fed00, 32'h00000000} /* (16, 2, 10) {real, imag} */,
  {32'h3f53a15b, 32'h00000000} /* (16, 2, 9) {real, imag} */,
  {32'h3f54c7ba, 32'h00000000} /* (16, 2, 8) {real, imag} */,
  {32'h3ed0e550, 32'h00000000} /* (16, 2, 7) {real, imag} */,
  {32'h3e06fd96, 32'h00000000} /* (16, 2, 6) {real, imag} */,
  {32'h3c07dbc5, 32'h00000000} /* (16, 2, 5) {real, imag} */,
  {32'hbe8a9272, 32'h00000000} /* (16, 2, 4) {real, imag} */,
  {32'hbe9bc233, 32'h00000000} /* (16, 2, 3) {real, imag} */,
  {32'hbf105521, 32'h00000000} /* (16, 2, 2) {real, imag} */,
  {32'hbea91d3b, 32'h00000000} /* (16, 2, 1) {real, imag} */,
  {32'hbe10a873, 32'h00000000} /* (16, 2, 0) {real, imag} */,
  {32'h3d94d406, 32'h00000000} /* (16, 1, 31) {real, imag} */,
  {32'hbe278916, 32'h00000000} /* (16, 1, 30) {real, imag} */,
  {32'hbeca588a, 32'h00000000} /* (16, 1, 29) {real, imag} */,
  {32'hbf55a41c, 32'h00000000} /* (16, 1, 28) {real, imag} */,
  {32'hbeb15941, 32'h00000000} /* (16, 1, 27) {real, imag} */,
  {32'hbf02852c, 32'h00000000} /* (16, 1, 26) {real, imag} */,
  {32'hbf1ecf97, 32'h00000000} /* (16, 1, 25) {real, imag} */,
  {32'hbf3e7fa5, 32'h00000000} /* (16, 1, 24) {real, imag} */,
  {32'hbe834eed, 32'h00000000} /* (16, 1, 23) {real, imag} */,
  {32'hbf31b8c3, 32'h00000000} /* (16, 1, 22) {real, imag} */,
  {32'hbf0a5429, 32'h00000000} /* (16, 1, 21) {real, imag} */,
  {32'hbe69f1a6, 32'h00000000} /* (16, 1, 20) {real, imag} */,
  {32'hbf008d5a, 32'h00000000} /* (16, 1, 19) {real, imag} */,
  {32'hbf8a954f, 32'h00000000} /* (16, 1, 18) {real, imag} */,
  {32'hbf13aa8b, 32'h00000000} /* (16, 1, 17) {real, imag} */,
  {32'h3dcc6518, 32'h00000000} /* (16, 1, 16) {real, imag} */,
  {32'h3ef82e65, 32'h00000000} /* (16, 1, 15) {real, imag} */,
  {32'h3f3c823b, 32'h00000000} /* (16, 1, 14) {real, imag} */,
  {32'h3f72638a, 32'h00000000} /* (16, 1, 13) {real, imag} */,
  {32'h3f84f37d, 32'h00000000} /* (16, 1, 12) {real, imag} */,
  {32'h3f05d94e, 32'h00000000} /* (16, 1, 11) {real, imag} */,
  {32'h3ec4ed07, 32'h00000000} /* (16, 1, 10) {real, imag} */,
  {32'h3e9e329c, 32'h00000000} /* (16, 1, 9) {real, imag} */,
  {32'h3f04e573, 32'h00000000} /* (16, 1, 8) {real, imag} */,
  {32'h3de7f103, 32'h00000000} /* (16, 1, 7) {real, imag} */,
  {32'hbdf3881a, 32'h00000000} /* (16, 1, 6) {real, imag} */,
  {32'hbe8808fa, 32'h00000000} /* (16, 1, 5) {real, imag} */,
  {32'hbf23f343, 32'h00000000} /* (16, 1, 4) {real, imag} */,
  {32'hbee194a1, 32'h00000000} /* (16, 1, 3) {real, imag} */,
  {32'hbea6a8cf, 32'h00000000} /* (16, 1, 2) {real, imag} */,
  {32'hbeab3779, 32'h00000000} /* (16, 1, 1) {real, imag} */,
  {32'hbee28564, 32'h00000000} /* (16, 1, 0) {real, imag} */,
  {32'hbd0d58ea, 32'h00000000} /* (16, 0, 31) {real, imag} */,
  {32'hbe4ccb60, 32'h00000000} /* (16, 0, 30) {real, imag} */,
  {32'hbe8a5677, 32'h00000000} /* (16, 0, 29) {real, imag} */,
  {32'hbe97d80e, 32'h00000000} /* (16, 0, 28) {real, imag} */,
  {32'hbe473574, 32'h00000000} /* (16, 0, 27) {real, imag} */,
  {32'hbe9c598c, 32'h00000000} /* (16, 0, 26) {real, imag} */,
  {32'hbed86afc, 32'h00000000} /* (16, 0, 25) {real, imag} */,
  {32'hbf37eaed, 32'h00000000} /* (16, 0, 24) {real, imag} */,
  {32'hbee8b780, 32'h00000000} /* (16, 0, 23) {real, imag} */,
  {32'hbf5724cc, 32'h00000000} /* (16, 0, 22) {real, imag} */,
  {32'hbf0d557b, 32'h00000000} /* (16, 0, 21) {real, imag} */,
  {32'hbeb5ab35, 32'h00000000} /* (16, 0, 20) {real, imag} */,
  {32'hbe983ad3, 32'h00000000} /* (16, 0, 19) {real, imag} */,
  {32'hbecdee77, 32'h00000000} /* (16, 0, 18) {real, imag} */,
  {32'hbda92b62, 32'h00000000} /* (16, 0, 17) {real, imag} */,
  {32'h3ced7421, 32'h00000000} /* (16, 0, 16) {real, imag} */,
  {32'h3e2043cd, 32'h00000000} /* (16, 0, 15) {real, imag} */,
  {32'h3ebdc3f5, 32'h00000000} /* (16, 0, 14) {real, imag} */,
  {32'h3e856f46, 32'h00000000} /* (16, 0, 13) {real, imag} */,
  {32'h3f1ac4e7, 32'h00000000} /* (16, 0, 12) {real, imag} */,
  {32'h3f4a43d9, 32'h00000000} /* (16, 0, 11) {real, imag} */,
  {32'h3eae7cdb, 32'h00000000} /* (16, 0, 10) {real, imag} */,
  {32'h3d72b5a6, 32'h00000000} /* (16, 0, 9) {real, imag} */,
  {32'h3ca13005, 32'h00000000} /* (16, 0, 8) {real, imag} */,
  {32'h3d73edfa, 32'h00000000} /* (16, 0, 7) {real, imag} */,
  {32'h3e1ad25b, 32'h00000000} /* (16, 0, 6) {real, imag} */,
  {32'hbe3a20f7, 32'h00000000} /* (16, 0, 5) {real, imag} */,
  {32'hbebde513, 32'h00000000} /* (16, 0, 4) {real, imag} */,
  {32'hbe1fa0f1, 32'h00000000} /* (16, 0, 3) {real, imag} */,
  {32'h3d089e8b, 32'h00000000} /* (16, 0, 2) {real, imag} */,
  {32'hbdb2f238, 32'h00000000} /* (16, 0, 1) {real, imag} */,
  {32'hbea16a5c, 32'h00000000} /* (16, 0, 0) {real, imag} */,
  {32'h3e1be867, 32'h00000000} /* (15, 31, 31) {real, imag} */,
  {32'h3f07e143, 32'h00000000} /* (15, 31, 30) {real, imag} */,
  {32'h3f10af8f, 32'h00000000} /* (15, 31, 29) {real, imag} */,
  {32'h3ecbfb53, 32'h00000000} /* (15, 31, 28) {real, imag} */,
  {32'h3e92a00d, 32'h00000000} /* (15, 31, 27) {real, imag} */,
  {32'h3e229798, 32'h00000000} /* (15, 31, 26) {real, imag} */,
  {32'h3dfef34e, 32'h00000000} /* (15, 31, 25) {real, imag} */,
  {32'h3e55e6f1, 32'h00000000} /* (15, 31, 24) {real, imag} */,
  {32'h3ef7f350, 32'h00000000} /* (15, 31, 23) {real, imag} */,
  {32'h3efe3881, 32'h00000000} /* (15, 31, 22) {real, imag} */,
  {32'h3aa674e3, 32'h00000000} /* (15, 31, 21) {real, imag} */,
  {32'hbebfd2a8, 32'h00000000} /* (15, 31, 20) {real, imag} */,
  {32'hbe1ad0b8, 32'h00000000} /* (15, 31, 19) {real, imag} */,
  {32'hbe25a270, 32'h00000000} /* (15, 31, 18) {real, imag} */,
  {32'hbf3a41e3, 32'h00000000} /* (15, 31, 17) {real, imag} */,
  {32'hbede2980, 32'h00000000} /* (15, 31, 16) {real, imag} */,
  {32'hbf22651b, 32'h00000000} /* (15, 31, 15) {real, imag} */,
  {32'hbf1e0996, 32'h00000000} /* (15, 31, 14) {real, imag} */,
  {32'hbf4ba2e1, 32'h00000000} /* (15, 31, 13) {real, imag} */,
  {32'hbf59d09a, 32'h00000000} /* (15, 31, 12) {real, imag} */,
  {32'hbf21c9aa, 32'h00000000} /* (15, 31, 11) {real, imag} */,
  {32'hbeb1e5c3, 32'h00000000} /* (15, 31, 10) {real, imag} */,
  {32'h3d04cdf1, 32'h00000000} /* (15, 31, 9) {real, imag} */,
  {32'h3e0536de, 32'h00000000} /* (15, 31, 8) {real, imag} */,
  {32'h3dcf746b, 32'h00000000} /* (15, 31, 7) {real, imag} */,
  {32'h3f4e9b72, 32'h00000000} /* (15, 31, 6) {real, imag} */,
  {32'h3f20dbaf, 32'h00000000} /* (15, 31, 5) {real, imag} */,
  {32'h3e64550a, 32'h00000000} /* (15, 31, 4) {real, imag} */,
  {32'h3ed940d5, 32'h00000000} /* (15, 31, 3) {real, imag} */,
  {32'h3f419998, 32'h00000000} /* (15, 31, 2) {real, imag} */,
  {32'h3f30f89d, 32'h00000000} /* (15, 31, 1) {real, imag} */,
  {32'h3e4799ec, 32'h00000000} /* (15, 31, 0) {real, imag} */,
  {32'h3e7c40fd, 32'h00000000} /* (15, 30, 31) {real, imag} */,
  {32'h3ec795b8, 32'h00000000} /* (15, 30, 30) {real, imag} */,
  {32'h3d806428, 32'h00000000} /* (15, 30, 29) {real, imag} */,
  {32'h3eba289a, 32'h00000000} /* (15, 30, 28) {real, imag} */,
  {32'h3eb0de30, 32'h00000000} /* (15, 30, 27) {real, imag} */,
  {32'h3e80c54a, 32'h00000000} /* (15, 30, 26) {real, imag} */,
  {32'h3f1e5d44, 32'h00000000} /* (15, 30, 25) {real, imag} */,
  {32'h3f47691f, 32'h00000000} /* (15, 30, 24) {real, imag} */,
  {32'h3f5b2b52, 32'h00000000} /* (15, 30, 23) {real, imag} */,
  {32'h3f5127f0, 32'h00000000} /* (15, 30, 22) {real, imag} */,
  {32'h3e84cfb7, 32'h00000000} /* (15, 30, 21) {real, imag} */,
  {32'hbe3a16e5, 32'h00000000} /* (15, 30, 20) {real, imag} */,
  {32'hbde9f5ed, 32'h00000000} /* (15, 30, 19) {real, imag} */,
  {32'hbf0b4280, 32'h00000000} /* (15, 30, 18) {real, imag} */,
  {32'hbf821ce0, 32'h00000000} /* (15, 30, 17) {real, imag} */,
  {32'hbf4ef6b6, 32'h00000000} /* (15, 30, 16) {real, imag} */,
  {32'hbeabd9a7, 32'h00000000} /* (15, 30, 15) {real, imag} */,
  {32'hbec478c2, 32'h00000000} /* (15, 30, 14) {real, imag} */,
  {32'hbf49f5f8, 32'h00000000} /* (15, 30, 13) {real, imag} */,
  {32'hbf9fa88f, 32'h00000000} /* (15, 30, 12) {real, imag} */,
  {32'hbeea30d2, 32'h00000000} /* (15, 30, 11) {real, imag} */,
  {32'h3da24614, 32'h00000000} /* (15, 30, 10) {real, imag} */,
  {32'h3e852ed3, 32'h00000000} /* (15, 30, 9) {real, imag} */,
  {32'h3ec7737d, 32'h00000000} /* (15, 30, 8) {real, imag} */,
  {32'h3e0cc49d, 32'h00000000} /* (15, 30, 7) {real, imag} */,
  {32'h3f6ffc9d, 32'h00000000} /* (15, 30, 6) {real, imag} */,
  {32'h3fa8fee9, 32'h00000000} /* (15, 30, 5) {real, imag} */,
  {32'h3e388354, 32'h00000000} /* (15, 30, 4) {real, imag} */,
  {32'h3e17f5eb, 32'h00000000} /* (15, 30, 3) {real, imag} */,
  {32'h3ee0cb2b, 32'h00000000} /* (15, 30, 2) {real, imag} */,
  {32'h3faa4f35, 32'h00000000} /* (15, 30, 1) {real, imag} */,
  {32'h3f6e385e, 32'h00000000} /* (15, 30, 0) {real, imag} */,
  {32'h3e51c439, 32'h00000000} /* (15, 29, 31) {real, imag} */,
  {32'h3e4dbe7b, 32'h00000000} /* (15, 29, 30) {real, imag} */,
  {32'hbe454e7b, 32'h00000000} /* (15, 29, 29) {real, imag} */,
  {32'h3f302523, 32'h00000000} /* (15, 29, 28) {real, imag} */,
  {32'h3f522ef8, 32'h00000000} /* (15, 29, 27) {real, imag} */,
  {32'h3e9a05d5, 32'h00000000} /* (15, 29, 26) {real, imag} */,
  {32'h3ee2d0d6, 32'h00000000} /* (15, 29, 25) {real, imag} */,
  {32'h3f1bc2b1, 32'h00000000} /* (15, 29, 24) {real, imag} */,
  {32'h3f2234f3, 32'h00000000} /* (15, 29, 23) {real, imag} */,
  {32'h3f7876e7, 32'h00000000} /* (15, 29, 22) {real, imag} */,
  {32'h3f51cf58, 32'h00000000} /* (15, 29, 21) {real, imag} */,
  {32'h3e419725, 32'h00000000} /* (15, 29, 20) {real, imag} */,
  {32'hbd06854a, 32'h00000000} /* (15, 29, 19) {real, imag} */,
  {32'hbdf72690, 32'h00000000} /* (15, 29, 18) {real, imag} */,
  {32'hbe367970, 32'h00000000} /* (15, 29, 17) {real, imag} */,
  {32'hbf374fac, 32'h00000000} /* (15, 29, 16) {real, imag} */,
  {32'hbeb9e8df, 32'h00000000} /* (15, 29, 15) {real, imag} */,
  {32'hbeafb3d5, 32'h00000000} /* (15, 29, 14) {real, imag} */,
  {32'hbddbf400, 32'h00000000} /* (15, 29, 13) {real, imag} */,
  {32'hbe4d6ce4, 32'h00000000} /* (15, 29, 12) {real, imag} */,
  {32'h3a946cdd, 32'h00000000} /* (15, 29, 11) {real, imag} */,
  {32'h3ec358fe, 32'h00000000} /* (15, 29, 10) {real, imag} */,
  {32'h3e98ebec, 32'h00000000} /* (15, 29, 9) {real, imag} */,
  {32'h3e94c84f, 32'h00000000} /* (15, 29, 8) {real, imag} */,
  {32'h3e9862e7, 32'h00000000} /* (15, 29, 7) {real, imag} */,
  {32'h3ed7e7c7, 32'h00000000} /* (15, 29, 6) {real, imag} */,
  {32'h3fa6a789, 32'h00000000} /* (15, 29, 5) {real, imag} */,
  {32'h3f131f0f, 32'h00000000} /* (15, 29, 4) {real, imag} */,
  {32'hbdc190e0, 32'h00000000} /* (15, 29, 3) {real, imag} */,
  {32'hbe8961ae, 32'h00000000} /* (15, 29, 2) {real, imag} */,
  {32'h3f0c6aad, 32'h00000000} /* (15, 29, 1) {real, imag} */,
  {32'h3f2f7682, 32'h00000000} /* (15, 29, 0) {real, imag} */,
  {32'h3df3f846, 32'h00000000} /* (15, 28, 31) {real, imag} */,
  {32'h3e6c4bcd, 32'h00000000} /* (15, 28, 30) {real, imag} */,
  {32'h3e4bc09c, 32'h00000000} /* (15, 28, 29) {real, imag} */,
  {32'h3f3e453b, 32'h00000000} /* (15, 28, 28) {real, imag} */,
  {32'h3f2bc4d1, 32'h00000000} /* (15, 28, 27) {real, imag} */,
  {32'h3f15862e, 32'h00000000} /* (15, 28, 26) {real, imag} */,
  {32'h3ed38607, 32'h00000000} /* (15, 28, 25) {real, imag} */,
  {32'h3eca5ade, 32'h00000000} /* (15, 28, 24) {real, imag} */,
  {32'h3f6354d6, 32'h00000000} /* (15, 28, 23) {real, imag} */,
  {32'h3fb5afe8, 32'h00000000} /* (15, 28, 22) {real, imag} */,
  {32'h3f7943f3, 32'h00000000} /* (15, 28, 21) {real, imag} */,
  {32'hbe95cf4e, 32'h00000000} /* (15, 28, 20) {real, imag} */,
  {32'hbedcca16, 32'h00000000} /* (15, 28, 19) {real, imag} */,
  {32'h3e1ad866, 32'h00000000} /* (15, 28, 18) {real, imag} */,
  {32'hbd8d7212, 32'h00000000} /* (15, 28, 17) {real, imag} */,
  {32'hbea8cd26, 32'h00000000} /* (15, 28, 16) {real, imag} */,
  {32'h3db517b1, 32'h00000000} /* (15, 28, 15) {real, imag} */,
  {32'h3df3abf4, 32'h00000000} /* (15, 28, 14) {real, imag} */,
  {32'h3e7c6907, 32'h00000000} /* (15, 28, 13) {real, imag} */,
  {32'h3e429823, 32'h00000000} /* (15, 28, 12) {real, imag} */,
  {32'h3e2f4aa8, 32'h00000000} /* (15, 28, 11) {real, imag} */,
  {32'h3f381468, 32'h00000000} /* (15, 28, 10) {real, imag} */,
  {32'h3f0d0837, 32'h00000000} /* (15, 28, 9) {real, imag} */,
  {32'h3f500661, 32'h00000000} /* (15, 28, 8) {real, imag} */,
  {32'h3e9c5c42, 32'h00000000} /* (15, 28, 7) {real, imag} */,
  {32'h3e66574f, 32'h00000000} /* (15, 28, 6) {real, imag} */,
  {32'h3f23d229, 32'h00000000} /* (15, 28, 5) {real, imag} */,
  {32'h3e6dbbaf, 32'h00000000} /* (15, 28, 4) {real, imag} */,
  {32'hbde25124, 32'h00000000} /* (15, 28, 3) {real, imag} */,
  {32'hbee378d8, 32'h00000000} /* (15, 28, 2) {real, imag} */,
  {32'hbd685d6c, 32'h00000000} /* (15, 28, 1) {real, imag} */,
  {32'h3ec3f43d, 32'h00000000} /* (15, 28, 0) {real, imag} */,
  {32'h3e5ecfb2, 32'h00000000} /* (15, 27, 31) {real, imag} */,
  {32'h3f243d87, 32'h00000000} /* (15, 27, 30) {real, imag} */,
  {32'h3eb126a5, 32'h00000000} /* (15, 27, 29) {real, imag} */,
  {32'h3e521154, 32'h00000000} /* (15, 27, 28) {real, imag} */,
  {32'h3d873559, 32'h00000000} /* (15, 27, 27) {real, imag} */,
  {32'h3f384416, 32'h00000000} /* (15, 27, 26) {real, imag} */,
  {32'h3f8aa9f4, 32'h00000000} /* (15, 27, 25) {real, imag} */,
  {32'h3eceb856, 32'h00000000} /* (15, 27, 24) {real, imag} */,
  {32'h3edb9260, 32'h00000000} /* (15, 27, 23) {real, imag} */,
  {32'h3f7e9bc1, 32'h00000000} /* (15, 27, 22) {real, imag} */,
  {32'h3fb66f0a, 32'h00000000} /* (15, 27, 21) {real, imag} */,
  {32'hbe9812d7, 32'h00000000} /* (15, 27, 20) {real, imag} */,
  {32'hbf135bf1, 32'h00000000} /* (15, 27, 19) {real, imag} */,
  {32'hbe457e50, 32'h00000000} /* (15, 27, 18) {real, imag} */,
  {32'hbf1abfb3, 32'h00000000} /* (15, 27, 17) {real, imag} */,
  {32'hbf44cfd2, 32'h00000000} /* (15, 27, 16) {real, imag} */,
  {32'hbec02f69, 32'h00000000} /* (15, 27, 15) {real, imag} */,
  {32'hbd29c406, 32'h00000000} /* (15, 27, 14) {real, imag} */,
  {32'hbdcd7f7c, 32'h00000000} /* (15, 27, 13) {real, imag} */,
  {32'hbd80c423, 32'h00000000} /* (15, 27, 12) {real, imag} */,
  {32'hbe22611b, 32'h00000000} /* (15, 27, 11) {real, imag} */,
  {32'h3f46e5a6, 32'h00000000} /* (15, 27, 10) {real, imag} */,
  {32'h3f2820e0, 32'h00000000} /* (15, 27, 9) {real, imag} */,
  {32'h3ee32d8f, 32'h00000000} /* (15, 27, 8) {real, imag} */,
  {32'h3e846cfc, 32'h00000000} /* (15, 27, 7) {real, imag} */,
  {32'h3f2769ae, 32'h00000000} /* (15, 27, 6) {real, imag} */,
  {32'h3f62c342, 32'h00000000} /* (15, 27, 5) {real, imag} */,
  {32'h3e40e960, 32'h00000000} /* (15, 27, 4) {real, imag} */,
  {32'h3e077b72, 32'h00000000} /* (15, 27, 3) {real, imag} */,
  {32'h3e2c1863, 32'h00000000} /* (15, 27, 2) {real, imag} */,
  {32'hbc5a84ae, 32'h00000000} /* (15, 27, 1) {real, imag} */,
  {32'h3e0cbce1, 32'h00000000} /* (15, 27, 0) {real, imag} */,
  {32'hbd4b51b8, 32'h00000000} /* (15, 26, 31) {real, imag} */,
  {32'h3e847fb1, 32'h00000000} /* (15, 26, 30) {real, imag} */,
  {32'h3ee596f0, 32'h00000000} /* (15, 26, 29) {real, imag} */,
  {32'h3f1390bb, 32'h00000000} /* (15, 26, 28) {real, imag} */,
  {32'h3e8c0738, 32'h00000000} /* (15, 26, 27) {real, imag} */,
  {32'h3ef24a41, 32'h00000000} /* (15, 26, 26) {real, imag} */,
  {32'h3f1de892, 32'h00000000} /* (15, 26, 25) {real, imag} */,
  {32'hbe099802, 32'h00000000} /* (15, 26, 24) {real, imag} */,
  {32'h3debdc79, 32'h00000000} /* (15, 26, 23) {real, imag} */,
  {32'h3f0490c1, 32'h00000000} /* (15, 26, 22) {real, imag} */,
  {32'h3f50d9f2, 32'h00000000} /* (15, 26, 21) {real, imag} */,
  {32'hbebd091c, 32'h00000000} /* (15, 26, 20) {real, imag} */,
  {32'hbf0f55e7, 32'h00000000} /* (15, 26, 19) {real, imag} */,
  {32'hbf2f2572, 32'h00000000} /* (15, 26, 18) {real, imag} */,
  {32'hbf966241, 32'h00000000} /* (15, 26, 17) {real, imag} */,
  {32'hbf8ec87d, 32'h00000000} /* (15, 26, 16) {real, imag} */,
  {32'hbe5abbac, 32'h00000000} /* (15, 26, 15) {real, imag} */,
  {32'hbe303855, 32'h00000000} /* (15, 26, 14) {real, imag} */,
  {32'hbf002c78, 32'h00000000} /* (15, 26, 13) {real, imag} */,
  {32'hbee1f2a8, 32'h00000000} /* (15, 26, 12) {real, imag} */,
  {32'hbe975f62, 32'h00000000} /* (15, 26, 11) {real, imag} */,
  {32'h3f231a75, 32'h00000000} /* (15, 26, 10) {real, imag} */,
  {32'h3eae7b15, 32'h00000000} /* (15, 26, 9) {real, imag} */,
  {32'h3e0cd31b, 32'h00000000} /* (15, 26, 8) {real, imag} */,
  {32'h3f23aed2, 32'h00000000} /* (15, 26, 7) {real, imag} */,
  {32'h3f2f85f5, 32'h00000000} /* (15, 26, 6) {real, imag} */,
  {32'h3ef53fd5, 32'h00000000} /* (15, 26, 5) {real, imag} */,
  {32'h3ecafc33, 32'h00000000} /* (15, 26, 4) {real, imag} */,
  {32'h3f779e03, 32'h00000000} /* (15, 26, 3) {real, imag} */,
  {32'h3f3b9585, 32'h00000000} /* (15, 26, 2) {real, imag} */,
  {32'h3e7ea1fa, 32'h00000000} /* (15, 26, 1) {real, imag} */,
  {32'h3e601710, 32'h00000000} /* (15, 26, 0) {real, imag} */,
  {32'h3dc09355, 32'h00000000} /* (15, 25, 31) {real, imag} */,
  {32'h3dfd25dd, 32'h00000000} /* (15, 25, 30) {real, imag} */,
  {32'h3e96b7ca, 32'h00000000} /* (15, 25, 29) {real, imag} */,
  {32'h3f39ed59, 32'h00000000} /* (15, 25, 28) {real, imag} */,
  {32'h3f10d4cf, 32'h00000000} /* (15, 25, 27) {real, imag} */,
  {32'h3ed4e071, 32'h00000000} /* (15, 25, 26) {real, imag} */,
  {32'h3e8b44f7, 32'h00000000} /* (15, 25, 25) {real, imag} */,
  {32'h3e73a9b0, 32'h00000000} /* (15, 25, 24) {real, imag} */,
  {32'h3ef24034, 32'h00000000} /* (15, 25, 23) {real, imag} */,
  {32'h3f16e79c, 32'h00000000} /* (15, 25, 22) {real, imag} */,
  {32'h3f10432d, 32'h00000000} /* (15, 25, 21) {real, imag} */,
  {32'hbe08a507, 32'h00000000} /* (15, 25, 20) {real, imag} */,
  {32'hbefbda26, 32'h00000000} /* (15, 25, 19) {real, imag} */,
  {32'hbf2257a1, 32'h00000000} /* (15, 25, 18) {real, imag} */,
  {32'hbf21d469, 32'h00000000} /* (15, 25, 17) {real, imag} */,
  {32'hbf588617, 32'h00000000} /* (15, 25, 16) {real, imag} */,
  {32'hbed3e4e3, 32'h00000000} /* (15, 25, 15) {real, imag} */,
  {32'hbeccb4d2, 32'h00000000} /* (15, 25, 14) {real, imag} */,
  {32'hbf4f41de, 32'h00000000} /* (15, 25, 13) {real, imag} */,
  {32'hbef76113, 32'h00000000} /* (15, 25, 12) {real, imag} */,
  {32'h3e4818e0, 32'h00000000} /* (15, 25, 11) {real, imag} */,
  {32'h3f1db9d2, 32'h00000000} /* (15, 25, 10) {real, imag} */,
  {32'h3f006754, 32'h00000000} /* (15, 25, 9) {real, imag} */,
  {32'h3f3e0237, 32'h00000000} /* (15, 25, 8) {real, imag} */,
  {32'h3f32c201, 32'h00000000} /* (15, 25, 7) {real, imag} */,
  {32'h3f18d9e8, 32'h00000000} /* (15, 25, 6) {real, imag} */,
  {32'h3f0e3334, 32'h00000000} /* (15, 25, 5) {real, imag} */,
  {32'h3eeacde2, 32'h00000000} /* (15, 25, 4) {real, imag} */,
  {32'h3f1cda24, 32'h00000000} /* (15, 25, 3) {real, imag} */,
  {32'h3f19ed22, 32'h00000000} /* (15, 25, 2) {real, imag} */,
  {32'h3f880499, 32'h00000000} /* (15, 25, 1) {real, imag} */,
  {32'h3f1def90, 32'h00000000} /* (15, 25, 0) {real, imag} */,
  {32'h3ea07cfc, 32'h00000000} /* (15, 24, 31) {real, imag} */,
  {32'h3f0e0ae7, 32'h00000000} /* (15, 24, 30) {real, imag} */,
  {32'h3f54b198, 32'h00000000} /* (15, 24, 29) {real, imag} */,
  {32'h3f7c1a0c, 32'h00000000} /* (15, 24, 28) {real, imag} */,
  {32'h3ebdaa39, 32'h00000000} /* (15, 24, 27) {real, imag} */,
  {32'hbdc5db4a, 32'h00000000} /* (15, 24, 26) {real, imag} */,
  {32'hbd9552e8, 32'h00000000} /* (15, 24, 25) {real, imag} */,
  {32'h3f062ef4, 32'h00000000} /* (15, 24, 24) {real, imag} */,
  {32'h3f55dcf2, 32'h00000000} /* (15, 24, 23) {real, imag} */,
  {32'h3f3f99ee, 32'h00000000} /* (15, 24, 22) {real, imag} */,
  {32'h3eafe878, 32'h00000000} /* (15, 24, 21) {real, imag} */,
  {32'hbe36d6ce, 32'h00000000} /* (15, 24, 20) {real, imag} */,
  {32'hbe9f5458, 32'h00000000} /* (15, 24, 19) {real, imag} */,
  {32'hbdee58ee, 32'h00000000} /* (15, 24, 18) {real, imag} */,
  {32'hbe874ba0, 32'h00000000} /* (15, 24, 17) {real, imag} */,
  {32'hbf3b68bb, 32'h00000000} /* (15, 24, 16) {real, imag} */,
  {32'hbf3a25b9, 32'h00000000} /* (15, 24, 15) {real, imag} */,
  {32'hbf1a0794, 32'h00000000} /* (15, 24, 14) {real, imag} */,
  {32'hbee2cfab, 32'h00000000} /* (15, 24, 13) {real, imag} */,
  {32'hbcee1900, 32'h00000000} /* (15, 24, 12) {real, imag} */,
  {32'hbee984a0, 32'h00000000} /* (15, 24, 11) {real, imag} */,
  {32'hbc324920, 32'h00000000} /* (15, 24, 10) {real, imag} */,
  {32'h3f1ca7fa, 32'h00000000} /* (15, 24, 9) {real, imag} */,
  {32'h3f5b5f12, 32'h00000000} /* (15, 24, 8) {real, imag} */,
  {32'h3f323e74, 32'h00000000} /* (15, 24, 7) {real, imag} */,
  {32'h3f0fc4ab, 32'h00000000} /* (15, 24, 6) {real, imag} */,
  {32'h3f080a3e, 32'h00000000} /* (15, 24, 5) {real, imag} */,
  {32'h3ee02bf5, 32'h00000000} /* (15, 24, 4) {real, imag} */,
  {32'h3ef00c85, 32'h00000000} /* (15, 24, 3) {real, imag} */,
  {32'h3e8aa640, 32'h00000000} /* (15, 24, 2) {real, imag} */,
  {32'h3f1cb242, 32'h00000000} /* (15, 24, 1) {real, imag} */,
  {32'h3ec391f1, 32'h00000000} /* (15, 24, 0) {real, imag} */,
  {32'h3e9904be, 32'h00000000} /* (15, 23, 31) {real, imag} */,
  {32'h3f71f85b, 32'h00000000} /* (15, 23, 30) {real, imag} */,
  {32'h3fb47564, 32'h00000000} /* (15, 23, 29) {real, imag} */,
  {32'h3f6c2c2c, 32'h00000000} /* (15, 23, 28) {real, imag} */,
  {32'h3e10f474, 32'h00000000} /* (15, 23, 27) {real, imag} */,
  {32'hbdb9ec1b, 32'h00000000} /* (15, 23, 26) {real, imag} */,
  {32'h3c86c602, 32'h00000000} /* (15, 23, 25) {real, imag} */,
  {32'h3ed304d9, 32'h00000000} /* (15, 23, 24) {real, imag} */,
  {32'h3ea5c53f, 32'h00000000} /* (15, 23, 23) {real, imag} */,
  {32'h3e988bb2, 32'h00000000} /* (15, 23, 22) {real, imag} */,
  {32'h3e8623ab, 32'h00000000} /* (15, 23, 21) {real, imag} */,
  {32'hbdec81dc, 32'h00000000} /* (15, 23, 20) {real, imag} */,
  {32'hbea87434, 32'h00000000} /* (15, 23, 19) {real, imag} */,
  {32'hbe98eab3, 32'h00000000} /* (15, 23, 18) {real, imag} */,
  {32'hbf48366c, 32'h00000000} /* (15, 23, 17) {real, imag} */,
  {32'hbf866f55, 32'h00000000} /* (15, 23, 16) {real, imag} */,
  {32'hbf1fbb37, 32'h00000000} /* (15, 23, 15) {real, imag} */,
  {32'hbeb2ccd9, 32'h00000000} /* (15, 23, 14) {real, imag} */,
  {32'hbee06439, 32'h00000000} /* (15, 23, 13) {real, imag} */,
  {32'hbf32cb84, 32'h00000000} /* (15, 23, 12) {real, imag} */,
  {32'hbf195105, 32'h00000000} /* (15, 23, 11) {real, imag} */,
  {32'h3d167b8b, 32'h00000000} /* (15, 23, 10) {real, imag} */,
  {32'h3f419b02, 32'h00000000} /* (15, 23, 9) {real, imag} */,
  {32'h3f2825f4, 32'h00000000} /* (15, 23, 8) {real, imag} */,
  {32'h3f42f1ab, 32'h00000000} /* (15, 23, 7) {real, imag} */,
  {32'h3f07d030, 32'h00000000} /* (15, 23, 6) {real, imag} */,
  {32'h3f8e719a, 32'h00000000} /* (15, 23, 5) {real, imag} */,
  {32'h3f45de4b, 32'h00000000} /* (15, 23, 4) {real, imag} */,
  {32'h3ebaaf8a, 32'h00000000} /* (15, 23, 3) {real, imag} */,
  {32'hbdb4cda9, 32'h00000000} /* (15, 23, 2) {real, imag} */,
  {32'hbe1b049f, 32'h00000000} /* (15, 23, 1) {real, imag} */,
  {32'hbda9eb5a, 32'h00000000} /* (15, 23, 0) {real, imag} */,
  {32'h3f255243, 32'h00000000} /* (15, 22, 31) {real, imag} */,
  {32'h3f8e57d7, 32'h00000000} /* (15, 22, 30) {real, imag} */,
  {32'h3f97902e, 32'h00000000} /* (15, 22, 29) {real, imag} */,
  {32'h3f86fd3e, 32'h00000000} /* (15, 22, 28) {real, imag} */,
  {32'h3f06d6e5, 32'h00000000} /* (15, 22, 27) {real, imag} */,
  {32'h3dd83516, 32'h00000000} /* (15, 22, 26) {real, imag} */,
  {32'h3d6a955a, 32'h00000000} /* (15, 22, 25) {real, imag} */,
  {32'h3ee23524, 32'h00000000} /* (15, 22, 24) {real, imag} */,
  {32'h3efdce85, 32'h00000000} /* (15, 22, 23) {real, imag} */,
  {32'h3e980993, 32'h00000000} /* (15, 22, 22) {real, imag} */,
  {32'h3df47e2e, 32'h00000000} /* (15, 22, 21) {real, imag} */,
  {32'h3cb72bd6, 32'h00000000} /* (15, 22, 20) {real, imag} */,
  {32'hbe0254bf, 32'h00000000} /* (15, 22, 19) {real, imag} */,
  {32'hbed551bf, 32'h00000000} /* (15, 22, 18) {real, imag} */,
  {32'hbf6c9601, 32'h00000000} /* (15, 22, 17) {real, imag} */,
  {32'hbfa70c4b, 32'h00000000} /* (15, 22, 16) {real, imag} */,
  {32'hbf314fe4, 32'h00000000} /* (15, 22, 15) {real, imag} */,
  {32'hbe962202, 32'h00000000} /* (15, 22, 14) {real, imag} */,
  {32'hbeb38675, 32'h00000000} /* (15, 22, 13) {real, imag} */,
  {32'hbf4964bf, 32'h00000000} /* (15, 22, 12) {real, imag} */,
  {32'hbf29526c, 32'h00000000} /* (15, 22, 11) {real, imag} */,
  {32'h3e356654, 32'h00000000} /* (15, 22, 10) {real, imag} */,
  {32'h3ef8b644, 32'h00000000} /* (15, 22, 9) {real, imag} */,
  {32'h3f48051d, 32'h00000000} /* (15, 22, 8) {real, imag} */,
  {32'h3eb1d38b, 32'h00000000} /* (15, 22, 7) {real, imag} */,
  {32'h3ec1cc86, 32'h00000000} /* (15, 22, 6) {real, imag} */,
  {32'h3f7768df, 32'h00000000} /* (15, 22, 5) {real, imag} */,
  {32'h3f4cb95e, 32'h00000000} /* (15, 22, 4) {real, imag} */,
  {32'h3e28f529, 32'h00000000} /* (15, 22, 3) {real, imag} */,
  {32'h3e8cd730, 32'h00000000} /* (15, 22, 2) {real, imag} */,
  {32'h3e284e9b, 32'h00000000} /* (15, 22, 1) {real, imag} */,
  {32'h3dcc7e2e, 32'h00000000} /* (15, 22, 0) {real, imag} */,
  {32'h3ed29ada, 32'h00000000} /* (15, 21, 31) {real, imag} */,
  {32'h3f36b8f2, 32'h00000000} /* (15, 21, 30) {real, imag} */,
  {32'h3e8cc01f, 32'h00000000} /* (15, 21, 29) {real, imag} */,
  {32'h3eb0e060, 32'h00000000} /* (15, 21, 28) {real, imag} */,
  {32'h3eaf22c8, 32'h00000000} /* (15, 21, 27) {real, imag} */,
  {32'hbd99e570, 32'h00000000} /* (15, 21, 26) {real, imag} */,
  {32'hbe3b80fe, 32'h00000000} /* (15, 21, 25) {real, imag} */,
  {32'h3e6e9241, 32'h00000000} /* (15, 21, 24) {real, imag} */,
  {32'h3ecf72da, 32'h00000000} /* (15, 21, 23) {real, imag} */,
  {32'h3f22571b, 32'h00000000} /* (15, 21, 22) {real, imag} */,
  {32'h3eb89fd5, 32'h00000000} /* (15, 21, 21) {real, imag} */,
  {32'h3b94b10a, 32'h00000000} /* (15, 21, 20) {real, imag} */,
  {32'h3c144331, 32'h00000000} /* (15, 21, 19) {real, imag} */,
  {32'hbebc33ad, 32'h00000000} /* (15, 21, 18) {real, imag} */,
  {32'hbec84aea, 32'h00000000} /* (15, 21, 17) {real, imag} */,
  {32'hbf096e10, 32'h00000000} /* (15, 21, 16) {real, imag} */,
  {32'hbda9e2cd, 32'h00000000} /* (15, 21, 15) {real, imag} */,
  {32'hbea1cb47, 32'h00000000} /* (15, 21, 14) {real, imag} */,
  {32'hbf12679c, 32'h00000000} /* (15, 21, 13) {real, imag} */,
  {32'hbf03bb80, 32'h00000000} /* (15, 21, 12) {real, imag} */,
  {32'hbe80550e, 32'h00000000} /* (15, 21, 11) {real, imag} */,
  {32'hbc925d94, 32'h00000000} /* (15, 21, 10) {real, imag} */,
  {32'h3e6de56c, 32'h00000000} /* (15, 21, 9) {real, imag} */,
  {32'h3d32deeb, 32'h00000000} /* (15, 21, 8) {real, imag} */,
  {32'h3e820f94, 32'h00000000} /* (15, 21, 7) {real, imag} */,
  {32'h3e9cff8b, 32'h00000000} /* (15, 21, 6) {real, imag} */,
  {32'h3b69b24e, 32'h00000000} /* (15, 21, 5) {real, imag} */,
  {32'h3ee14e56, 32'h00000000} /* (15, 21, 4) {real, imag} */,
  {32'h3d58c0e8, 32'h00000000} /* (15, 21, 3) {real, imag} */,
  {32'hbe7ac366, 32'h00000000} /* (15, 21, 2) {real, imag} */,
  {32'h3d41d739, 32'h00000000} /* (15, 21, 1) {real, imag} */,
  {32'h3e7bfe24, 32'h00000000} /* (15, 21, 0) {real, imag} */,
  {32'h3e0f720f, 32'h00000000} /* (15, 20, 31) {real, imag} */,
  {32'h3d66b256, 32'h00000000} /* (15, 20, 30) {real, imag} */,
  {32'hbf15f44e, 32'h00000000} /* (15, 20, 29) {real, imag} */,
  {32'hbf3c17d8, 32'h00000000} /* (15, 20, 28) {real, imag} */,
  {32'hbf482202, 32'h00000000} /* (15, 20, 27) {real, imag} */,
  {32'hbf0c8b92, 32'h00000000} /* (15, 20, 26) {real, imag} */,
  {32'hbf197b25, 32'h00000000} /* (15, 20, 25) {real, imag} */,
  {32'hbed8fc58, 32'h00000000} /* (15, 20, 24) {real, imag} */,
  {32'hbeefd35c, 32'h00000000} /* (15, 20, 23) {real, imag} */,
  {32'hbe9bd9b0, 32'h00000000} /* (15, 20, 22) {real, imag} */,
  {32'hbcbbcfa0, 32'h00000000} /* (15, 20, 21) {real, imag} */,
  {32'h3ea03be9, 32'h00000000} /* (15, 20, 20) {real, imag} */,
  {32'h3e8d2132, 32'h00000000} /* (15, 20, 19) {real, imag} */,
  {32'hbdc12108, 32'h00000000} /* (15, 20, 18) {real, imag} */,
  {32'h3dbfc5a7, 32'h00000000} /* (15, 20, 17) {real, imag} */,
  {32'h3f2090d2, 32'h00000000} /* (15, 20, 16) {real, imag} */,
  {32'h3f6282a6, 32'h00000000} /* (15, 20, 15) {real, imag} */,
  {32'h3f19ea7f, 32'h00000000} /* (15, 20, 14) {real, imag} */,
  {32'h3eacc155, 32'h00000000} /* (15, 20, 13) {real, imag} */,
  {32'h3f080152, 32'h00000000} /* (15, 20, 12) {real, imag} */,
  {32'h3f1d1726, 32'h00000000} /* (15, 20, 11) {real, imag} */,
  {32'hbe9f1436, 32'h00000000} /* (15, 20, 10) {real, imag} */,
  {32'hbe430dea, 32'h00000000} /* (15, 20, 9) {real, imag} */,
  {32'hbdda941f, 32'h00000000} /* (15, 20, 8) {real, imag} */,
  {32'hbdcd373b, 32'h00000000} /* (15, 20, 7) {real, imag} */,
  {32'hbecc1e81, 32'h00000000} /* (15, 20, 6) {real, imag} */,
  {32'hbf442376, 32'h00000000} /* (15, 20, 5) {real, imag} */,
  {32'hbe9df61f, 32'h00000000} /* (15, 20, 4) {real, imag} */,
  {32'hbe35d34c, 32'h00000000} /* (15, 20, 3) {real, imag} */,
  {32'hbed07cb0, 32'h00000000} /* (15, 20, 2) {real, imag} */,
  {32'hbf1cde40, 32'h00000000} /* (15, 20, 1) {real, imag} */,
  {32'hbeaef727, 32'h00000000} /* (15, 20, 0) {real, imag} */,
  {32'hbd152722, 32'h00000000} /* (15, 19, 31) {real, imag} */,
  {32'hbe66095b, 32'h00000000} /* (15, 19, 30) {real, imag} */,
  {32'hbefc7a54, 32'h00000000} /* (15, 19, 29) {real, imag} */,
  {32'hbf20bc22, 32'h00000000} /* (15, 19, 28) {real, imag} */,
  {32'hbf8ef1d1, 32'h00000000} /* (15, 19, 27) {real, imag} */,
  {32'hbf28031d, 32'h00000000} /* (15, 19, 26) {real, imag} */,
  {32'hbf3a61c0, 32'h00000000} /* (15, 19, 25) {real, imag} */,
  {32'hbeb3a92c, 32'h00000000} /* (15, 19, 24) {real, imag} */,
  {32'hbeac34ad, 32'h00000000} /* (15, 19, 23) {real, imag} */,
  {32'hbeb5958d, 32'h00000000} /* (15, 19, 22) {real, imag} */,
  {32'h3e39e112, 32'h00000000} /* (15, 19, 21) {real, imag} */,
  {32'h3eeef652, 32'h00000000} /* (15, 19, 20) {real, imag} */,
  {32'h3effa579, 32'h00000000} /* (15, 19, 19) {real, imag} */,
  {32'h3e86da06, 32'h00000000} /* (15, 19, 18) {real, imag} */,
  {32'h3e9ace37, 32'h00000000} /* (15, 19, 17) {real, imag} */,
  {32'h3f52921b, 32'h00000000} /* (15, 19, 16) {real, imag} */,
  {32'h3f6b7382, 32'h00000000} /* (15, 19, 15) {real, imag} */,
  {32'h3f5c5edb, 32'h00000000} /* (15, 19, 14) {real, imag} */,
  {32'h3f8d5d58, 32'h00000000} /* (15, 19, 13) {real, imag} */,
  {32'h3f821287, 32'h00000000} /* (15, 19, 12) {real, imag} */,
  {32'h3edefc68, 32'h00000000} /* (15, 19, 11) {real, imag} */,
  {32'hbe9fdbf4, 32'h00000000} /* (15, 19, 10) {real, imag} */,
  {32'hbe858797, 32'h00000000} /* (15, 19, 9) {real, imag} */,
  {32'hbd8fccd3, 32'h00000000} /* (15, 19, 8) {real, imag} */,
  {32'hbee86641, 32'h00000000} /* (15, 19, 7) {real, imag} */,
  {32'hbeed0541, 32'h00000000} /* (15, 19, 6) {real, imag} */,
  {32'hbe9da4c3, 32'h00000000} /* (15, 19, 5) {real, imag} */,
  {32'hbf5054eb, 32'h00000000} /* (15, 19, 4) {real, imag} */,
  {32'hbee78eef, 32'h00000000} /* (15, 19, 3) {real, imag} */,
  {32'hbde09286, 32'h00000000} /* (15, 19, 2) {real, imag} */,
  {32'hbe90f4e6, 32'h00000000} /* (15, 19, 1) {real, imag} */,
  {32'hbebce72b, 32'h00000000} /* (15, 19, 0) {real, imag} */,
  {32'hbe3d551f, 32'h00000000} /* (15, 18, 31) {real, imag} */,
  {32'hbf046266, 32'h00000000} /* (15, 18, 30) {real, imag} */,
  {32'hbec856e8, 32'h00000000} /* (15, 18, 29) {real, imag} */,
  {32'hbed510a1, 32'h00000000} /* (15, 18, 28) {real, imag} */,
  {32'hbe9d01ae, 32'h00000000} /* (15, 18, 27) {real, imag} */,
  {32'hbe00db8a, 32'h00000000} /* (15, 18, 26) {real, imag} */,
  {32'hbe2788c8, 32'h00000000} /* (15, 18, 25) {real, imag} */,
  {32'h3eb2bb1f, 32'h00000000} /* (15, 18, 24) {real, imag} */,
  {32'hbed3c4e7, 32'h00000000} /* (15, 18, 23) {real, imag} */,
  {32'hbf3603a0, 32'h00000000} /* (15, 18, 22) {real, imag} */,
  {32'h3e9751fd, 32'h00000000} /* (15, 18, 21) {real, imag} */,
  {32'h3f01b4a4, 32'h00000000} /* (15, 18, 20) {real, imag} */,
  {32'h3f2b9d9e, 32'h00000000} /* (15, 18, 19) {real, imag} */,
  {32'h3f4e359d, 32'h00000000} /* (15, 18, 18) {real, imag} */,
  {32'h3f12c505, 32'h00000000} /* (15, 18, 17) {real, imag} */,
  {32'h3f015269, 32'h00000000} /* (15, 18, 16) {real, imag} */,
  {32'h3e73c311, 32'h00000000} /* (15, 18, 15) {real, imag} */,
  {32'h3e8941c0, 32'h00000000} /* (15, 18, 14) {real, imag} */,
  {32'h3f535996, 32'h00000000} /* (15, 18, 13) {real, imag} */,
  {32'h3f725eaa, 32'h00000000} /* (15, 18, 12) {real, imag} */,
  {32'h3f0a8b37, 32'h00000000} /* (15, 18, 11) {real, imag} */,
  {32'hbe8330de, 32'h00000000} /* (15, 18, 10) {real, imag} */,
  {32'hbf06e75a, 32'h00000000} /* (15, 18, 9) {real, imag} */,
  {32'hbf2e0c9d, 32'h00000000} /* (15, 18, 8) {real, imag} */,
  {32'hbf81b8fa, 32'h00000000} /* (15, 18, 7) {real, imag} */,
  {32'hbf70a53c, 32'h00000000} /* (15, 18, 6) {real, imag} */,
  {32'hbec0a024, 32'h00000000} /* (15, 18, 5) {real, imag} */,
  {32'hbb6a87a2, 32'h00000000} /* (15, 18, 4) {real, imag} */,
  {32'hbebfe4a6, 32'h00000000} /* (15, 18, 3) {real, imag} */,
  {32'hbe3c489b, 32'h00000000} /* (15, 18, 2) {real, imag} */,
  {32'hbe1eaa42, 32'h00000000} /* (15, 18, 1) {real, imag} */,
  {32'hbecacfba, 32'h00000000} /* (15, 18, 0) {real, imag} */,
  {32'hbe0a9ff1, 32'h00000000} /* (15, 17, 31) {real, imag} */,
  {32'hbf1e47c3, 32'h00000000} /* (15, 17, 30) {real, imag} */,
  {32'hbed4da5b, 32'h00000000} /* (15, 17, 29) {real, imag} */,
  {32'hbe57481f, 32'h00000000} /* (15, 17, 28) {real, imag} */,
  {32'hbf391ca2, 32'h00000000} /* (15, 17, 27) {real, imag} */,
  {32'hbf0bf2a1, 32'h00000000} /* (15, 17, 26) {real, imag} */,
  {32'hbed142ed, 32'h00000000} /* (15, 17, 25) {real, imag} */,
  {32'h3dc194e2, 32'h00000000} /* (15, 17, 24) {real, imag} */,
  {32'hbede5865, 32'h00000000} /* (15, 17, 23) {real, imag} */,
  {32'hbf4af095, 32'h00000000} /* (15, 17, 22) {real, imag} */,
  {32'hbba2e9df, 32'h00000000} /* (15, 17, 21) {real, imag} */,
  {32'h3ed6bc92, 32'h00000000} /* (15, 17, 20) {real, imag} */,
  {32'h3f425479, 32'h00000000} /* (15, 17, 19) {real, imag} */,
  {32'h3f7b24aa, 32'h00000000} /* (15, 17, 18) {real, imag} */,
  {32'h3f5354ef, 32'h00000000} /* (15, 17, 17) {real, imag} */,
  {32'h3ed12a5c, 32'h00000000} /* (15, 17, 16) {real, imag} */,
  {32'h3e0c48fa, 32'h00000000} /* (15, 17, 15) {real, imag} */,
  {32'hbe6f1140, 32'h00000000} /* (15, 17, 14) {real, imag} */,
  {32'h3d3a31f5, 32'h00000000} /* (15, 17, 13) {real, imag} */,
  {32'h3ef56e9d, 32'h00000000} /* (15, 17, 12) {real, imag} */,
  {32'h3d6ce517, 32'h00000000} /* (15, 17, 11) {real, imag} */,
  {32'hbf6b83fc, 32'h00000000} /* (15, 17, 10) {real, imag} */,
  {32'hbf5615b2, 32'h00000000} /* (15, 17, 9) {real, imag} */,
  {32'hbf0b6d04, 32'h00000000} /* (15, 17, 8) {real, imag} */,
  {32'hbf39597d, 32'h00000000} /* (15, 17, 7) {real, imag} */,
  {32'hbfa8da1b, 32'h00000000} /* (15, 17, 6) {real, imag} */,
  {32'hbf873f5c, 32'h00000000} /* (15, 17, 5) {real, imag} */,
  {32'hbebd2448, 32'h00000000} /* (15, 17, 4) {real, imag} */,
  {32'hbe2e095a, 32'h00000000} /* (15, 17, 3) {real, imag} */,
  {32'hbe84cfd9, 32'h00000000} /* (15, 17, 2) {real, imag} */,
  {32'hbf019a98, 32'h00000000} /* (15, 17, 1) {real, imag} */,
  {32'hbef35665, 32'h00000000} /* (15, 17, 0) {real, imag} */,
  {32'hbe6ce2a4, 32'h00000000} /* (15, 16, 31) {real, imag} */,
  {32'hbf4215d1, 32'h00000000} /* (15, 16, 30) {real, imag} */,
  {32'hbed40f1b, 32'h00000000} /* (15, 16, 29) {real, imag} */,
  {32'h3cf62a53, 32'h00000000} /* (15, 16, 28) {real, imag} */,
  {32'hbf69a42b, 32'h00000000} /* (15, 16, 27) {real, imag} */,
  {32'hbf910567, 32'h00000000} /* (15, 16, 26) {real, imag} */,
  {32'hbf8c9e02, 32'h00000000} /* (15, 16, 25) {real, imag} */,
  {32'hbf3e0d37, 32'h00000000} /* (15, 16, 24) {real, imag} */,
  {32'hbf0a925e, 32'h00000000} /* (15, 16, 23) {real, imag} */,
  {32'hbf60f371, 32'h00000000} /* (15, 16, 22) {real, imag} */,
  {32'hbe245c38, 32'h00000000} /* (15, 16, 21) {real, imag} */,
  {32'h3ebf09b0, 32'h00000000} /* (15, 16, 20) {real, imag} */,
  {32'h3f5a2b33, 32'h00000000} /* (15, 16, 19) {real, imag} */,
  {32'h3f9df2c6, 32'h00000000} /* (15, 16, 18) {real, imag} */,
  {32'h3f3997fe, 32'h00000000} /* (15, 16, 17) {real, imag} */,
  {32'h3e591d33, 32'h00000000} /* (15, 16, 16) {real, imag} */,
  {32'h3d758cdc, 32'h00000000} /* (15, 16, 15) {real, imag} */,
  {32'h3d9f3158, 32'h00000000} /* (15, 16, 14) {real, imag} */,
  {32'h3eb9d244, 32'h00000000} /* (15, 16, 13) {real, imag} */,
  {32'h3e875441, 32'h00000000} /* (15, 16, 12) {real, imag} */,
  {32'h3e3332bd, 32'h00000000} /* (15, 16, 11) {real, imag} */,
  {32'hbe9c1b72, 32'h00000000} /* (15, 16, 10) {real, imag} */,
  {32'hbf1d9587, 32'h00000000} /* (15, 16, 9) {real, imag} */,
  {32'hbf3aa502, 32'h00000000} /* (15, 16, 8) {real, imag} */,
  {32'hbf8260c1, 32'h00000000} /* (15, 16, 7) {real, imag} */,
  {32'hbf8f36c2, 32'h00000000} /* (15, 16, 6) {real, imag} */,
  {32'hbf5e2f4f, 32'h00000000} /* (15, 16, 5) {real, imag} */,
  {32'hbeb31494, 32'h00000000} /* (15, 16, 4) {real, imag} */,
  {32'hbd3a19c2, 32'h00000000} /* (15, 16, 3) {real, imag} */,
  {32'hbe90afa1, 32'h00000000} /* (15, 16, 2) {real, imag} */,
  {32'hbec37b64, 32'h00000000} /* (15, 16, 1) {real, imag} */,
  {32'hbe0fa3d2, 32'h00000000} /* (15, 16, 0) {real, imag} */,
  {32'hbeb682fe, 32'h00000000} /* (15, 15, 31) {real, imag} */,
  {32'hbf2bfa58, 32'h00000000} /* (15, 15, 30) {real, imag} */,
  {32'hbef827b5, 32'h00000000} /* (15, 15, 29) {real, imag} */,
  {32'hbe8ff132, 32'h00000000} /* (15, 15, 28) {real, imag} */,
  {32'hbf496fc9, 32'h00000000} /* (15, 15, 27) {real, imag} */,
  {32'hbfb5c7d7, 32'h00000000} /* (15, 15, 26) {real, imag} */,
  {32'hbfc1cf30, 32'h00000000} /* (15, 15, 25) {real, imag} */,
  {32'hbf52a6a5, 32'h00000000} /* (15, 15, 24) {real, imag} */,
  {32'hbf1d9f24, 32'h00000000} /* (15, 15, 23) {real, imag} */,
  {32'hbf0d9954, 32'h00000000} /* (15, 15, 22) {real, imag} */,
  {32'h3e1bbe23, 32'h00000000} /* (15, 15, 21) {real, imag} */,
  {32'h3e8388a3, 32'h00000000} /* (15, 15, 20) {real, imag} */,
  {32'h3f43d525, 32'h00000000} /* (15, 15, 19) {real, imag} */,
  {32'h3fb39377, 32'h00000000} /* (15, 15, 18) {real, imag} */,
  {32'h3f525f76, 32'h00000000} /* (15, 15, 17) {real, imag} */,
  {32'h3f4e95dc, 32'h00000000} /* (15, 15, 16) {real, imag} */,
  {32'h3ed35b40, 32'h00000000} /* (15, 15, 15) {real, imag} */,
  {32'h3ef0e923, 32'h00000000} /* (15, 15, 14) {real, imag} */,
  {32'h3f3f165a, 32'h00000000} /* (15, 15, 13) {real, imag} */,
  {32'h3f0fdd53, 32'h00000000} /* (15, 15, 12) {real, imag} */,
  {32'h3f13290c, 32'h00000000} /* (15, 15, 11) {real, imag} */,
  {32'hbe434c1a, 32'h00000000} /* (15, 15, 10) {real, imag} */,
  {32'hbf1ff13b, 32'h00000000} /* (15, 15, 9) {real, imag} */,
  {32'hbf1377e4, 32'h00000000} /* (15, 15, 8) {real, imag} */,
  {32'hbf2c146f, 32'h00000000} /* (15, 15, 7) {real, imag} */,
  {32'hbf6b6a99, 32'h00000000} /* (15, 15, 6) {real, imag} */,
  {32'hbf602a2e, 32'h00000000} /* (15, 15, 5) {real, imag} */,
  {32'hbe638422, 32'h00000000} /* (15, 15, 4) {real, imag} */,
  {32'hbdbf1457, 32'h00000000} /* (15, 15, 3) {real, imag} */,
  {32'hbef8a084, 32'h00000000} /* (15, 15, 2) {real, imag} */,
  {32'hbedfe949, 32'h00000000} /* (15, 15, 1) {real, imag} */,
  {32'hbe865a66, 32'h00000000} /* (15, 15, 0) {real, imag} */,
  {32'hbe94719a, 32'h00000000} /* (15, 14, 31) {real, imag} */,
  {32'hbf2a03c4, 32'h00000000} /* (15, 14, 30) {real, imag} */,
  {32'hbfc4dc39, 32'h00000000} /* (15, 14, 29) {real, imag} */,
  {32'hbfcfd7f7, 32'h00000000} /* (15, 14, 28) {real, imag} */,
  {32'hbf8c4a35, 32'h00000000} /* (15, 14, 27) {real, imag} */,
  {32'hbf9639e6, 32'h00000000} /* (15, 14, 26) {real, imag} */,
  {32'hbfcc934b, 32'h00000000} /* (15, 14, 25) {real, imag} */,
  {32'hbf580bb1, 32'h00000000} /* (15, 14, 24) {real, imag} */,
  {32'hbf0f7880, 32'h00000000} /* (15, 14, 23) {real, imag} */,
  {32'hbf026c76, 32'h00000000} /* (15, 14, 22) {real, imag} */,
  {32'hbed5691e, 32'h00000000} /* (15, 14, 21) {real, imag} */,
  {32'h3e81e003, 32'h00000000} /* (15, 14, 20) {real, imag} */,
  {32'h3f19fbc5, 32'h00000000} /* (15, 14, 19) {real, imag} */,
  {32'h3fa0d900, 32'h00000000} /* (15, 14, 18) {real, imag} */,
  {32'h3f8cf69b, 32'h00000000} /* (15, 14, 17) {real, imag} */,
  {32'h3f46b3a6, 32'h00000000} /* (15, 14, 16) {real, imag} */,
  {32'h3f476ce5, 32'h00000000} /* (15, 14, 15) {real, imag} */,
  {32'h3f177970, 32'h00000000} /* (15, 14, 14) {real, imag} */,
  {32'h3f323800, 32'h00000000} /* (15, 14, 13) {real, imag} */,
  {32'h3f1a812a, 32'h00000000} /* (15, 14, 12) {real, imag} */,
  {32'h3f4877eb, 32'h00000000} /* (15, 14, 11) {real, imag} */,
  {32'h3daf26e9, 32'h00000000} /* (15, 14, 10) {real, imag} */,
  {32'hbed8b860, 32'h00000000} /* (15, 14, 9) {real, imag} */,
  {32'hbea37556, 32'h00000000} /* (15, 14, 8) {real, imag} */,
  {32'hbf30bf78, 32'h00000000} /* (15, 14, 7) {real, imag} */,
  {32'hbf73b35f, 32'h00000000} /* (15, 14, 6) {real, imag} */,
  {32'hbf012ac1, 32'h00000000} /* (15, 14, 5) {real, imag} */,
  {32'hbe98a3ce, 32'h00000000} /* (15, 14, 4) {real, imag} */,
  {32'hbe82b208, 32'h00000000} /* (15, 14, 3) {real, imag} */,
  {32'hbf1f1cbd, 32'h00000000} /* (15, 14, 2) {real, imag} */,
  {32'hbf2e5f7d, 32'h00000000} /* (15, 14, 1) {real, imag} */,
  {32'hbec7d794, 32'h00000000} /* (15, 14, 0) {real, imag} */,
  {32'hbe363048, 32'h00000000} /* (15, 13, 31) {real, imag} */,
  {32'hbf1d2269, 32'h00000000} /* (15, 13, 30) {real, imag} */,
  {32'hbf565061, 32'h00000000} /* (15, 13, 29) {real, imag} */,
  {32'hbf3bcb9f, 32'h00000000} /* (15, 13, 28) {real, imag} */,
  {32'hbf1f9b67, 32'h00000000} /* (15, 13, 27) {real, imag} */,
  {32'hbf0730a9, 32'h00000000} /* (15, 13, 26) {real, imag} */,
  {32'hbf577fbd, 32'h00000000} /* (15, 13, 25) {real, imag} */,
  {32'hbf7a6009, 32'h00000000} /* (15, 13, 24) {real, imag} */,
  {32'hbf6e7322, 32'h00000000} /* (15, 13, 23) {real, imag} */,
  {32'hbf6f99c6, 32'h00000000} /* (15, 13, 22) {real, imag} */,
  {32'hbf5d12ad, 32'h00000000} /* (15, 13, 21) {real, imag} */,
  {32'hbe0eca80, 32'h00000000} /* (15, 13, 20) {real, imag} */,
  {32'h3f092e8b, 32'h00000000} /* (15, 13, 19) {real, imag} */,
  {32'h3f4b5490, 32'h00000000} /* (15, 13, 18) {real, imag} */,
  {32'h3f00b7f3, 32'h00000000} /* (15, 13, 17) {real, imag} */,
  {32'h3efd9dde, 32'h00000000} /* (15, 13, 16) {real, imag} */,
  {32'h3f007bff, 32'h00000000} /* (15, 13, 15) {real, imag} */,
  {32'h3f1e017c, 32'h00000000} /* (15, 13, 14) {real, imag} */,
  {32'h3f0abcde, 32'h00000000} /* (15, 13, 13) {real, imag} */,
  {32'h3f228211, 32'h00000000} /* (15, 13, 12) {real, imag} */,
  {32'h3eba8dc8, 32'h00000000} /* (15, 13, 11) {real, imag} */,
  {32'hbe257f73, 32'h00000000} /* (15, 13, 10) {real, imag} */,
  {32'hbe1a6c7a, 32'h00000000} /* (15, 13, 9) {real, imag} */,
  {32'hbe772d4e, 32'h00000000} /* (15, 13, 8) {real, imag} */,
  {32'hbf643711, 32'h00000000} /* (15, 13, 7) {real, imag} */,
  {32'hbf8b8afb, 32'h00000000} /* (15, 13, 6) {real, imag} */,
  {32'hbe9fd642, 32'h00000000} /* (15, 13, 5) {real, imag} */,
  {32'hbeb99353, 32'h00000000} /* (15, 13, 4) {real, imag} */,
  {32'hbea96b13, 32'h00000000} /* (15, 13, 3) {real, imag} */,
  {32'hbe88516a, 32'h00000000} /* (15, 13, 2) {real, imag} */,
  {32'hbea9da98, 32'h00000000} /* (15, 13, 1) {real, imag} */,
  {32'hbf0d714d, 32'h00000000} /* (15, 13, 0) {real, imag} */,
  {32'hbeb40f92, 32'h00000000} /* (15, 12, 31) {real, imag} */,
  {32'hbf3ad027, 32'h00000000} /* (15, 12, 30) {real, imag} */,
  {32'hbf1dbacb, 32'h00000000} /* (15, 12, 29) {real, imag} */,
  {32'hbdfecf56, 32'h00000000} /* (15, 12, 28) {real, imag} */,
  {32'hbe52dc40, 32'h00000000} /* (15, 12, 27) {real, imag} */,
  {32'hbe9d0aaa, 32'h00000000} /* (15, 12, 26) {real, imag} */,
  {32'hbf0ef543, 32'h00000000} /* (15, 12, 25) {real, imag} */,
  {32'hbf298756, 32'h00000000} /* (15, 12, 24) {real, imag} */,
  {32'hbf320793, 32'h00000000} /* (15, 12, 23) {real, imag} */,
  {32'hbf2d9496, 32'h00000000} /* (15, 12, 22) {real, imag} */,
  {32'h3d1b3ddf, 32'h00000000} /* (15, 12, 21) {real, imag} */,
  {32'h3ef676d5, 32'h00000000} /* (15, 12, 20) {real, imag} */,
  {32'h3f1f7291, 32'h00000000} /* (15, 12, 19) {real, imag} */,
  {32'h3f28a857, 32'h00000000} /* (15, 12, 18) {real, imag} */,
  {32'h3f7d3a3e, 32'h00000000} /* (15, 12, 17) {real, imag} */,
  {32'h3f5bf2c3, 32'h00000000} /* (15, 12, 16) {real, imag} */,
  {32'h3c9c6252, 32'h00000000} /* (15, 12, 15) {real, imag} */,
  {32'h3de8232f, 32'h00000000} /* (15, 12, 14) {real, imag} */,
  {32'h3f3ec477, 32'h00000000} /* (15, 12, 13) {real, imag} */,
  {32'h3fab8664, 32'h00000000} /* (15, 12, 12) {real, imag} */,
  {32'h3f81dd96, 32'h00000000} /* (15, 12, 11) {real, imag} */,
  {32'hbe3d2bac, 32'h00000000} /* (15, 12, 10) {real, imag} */,
  {32'hbedb5bc0, 32'h00000000} /* (15, 12, 9) {real, imag} */,
  {32'hbf64b612, 32'h00000000} /* (15, 12, 8) {real, imag} */,
  {32'hbefeb54b, 32'h00000000} /* (15, 12, 7) {real, imag} */,
  {32'hbe386099, 32'h00000000} /* (15, 12, 6) {real, imag} */,
  {32'hbe3c43af, 32'h00000000} /* (15, 12, 5) {real, imag} */,
  {32'hbec3e677, 32'h00000000} /* (15, 12, 4) {real, imag} */,
  {32'hbefd3dc4, 32'h00000000} /* (15, 12, 3) {real, imag} */,
  {32'hbdff68b4, 32'h00000000} /* (15, 12, 2) {real, imag} */,
  {32'hbe547678, 32'h00000000} /* (15, 12, 1) {real, imag} */,
  {32'hbea55966, 32'h00000000} /* (15, 12, 0) {real, imag} */,
  {32'h3e4ea0e0, 32'h00000000} /* (15, 11, 31) {real, imag} */,
  {32'h3e2abe97, 32'h00000000} /* (15, 11, 30) {real, imag} */,
  {32'hbf07ef4e, 32'h00000000} /* (15, 11, 29) {real, imag} */,
  {32'hbecd54d0, 32'h00000000} /* (15, 11, 28) {real, imag} */,
  {32'hbe403fee, 32'h00000000} /* (15, 11, 27) {real, imag} */,
  {32'hbece7282, 32'h00000000} /* (15, 11, 26) {real, imag} */,
  {32'hbec56c46, 32'h00000000} /* (15, 11, 25) {real, imag} */,
  {32'hbe9728c2, 32'h00000000} /* (15, 11, 24) {real, imag} */,
  {32'hbfab82c7, 32'h00000000} /* (15, 11, 23) {real, imag} */,
  {32'hbe9f09fb, 32'h00000000} /* (15, 11, 22) {real, imag} */,
  {32'h3f119b9d, 32'h00000000} /* (15, 11, 21) {real, imag} */,
  {32'h3f3882c2, 32'h00000000} /* (15, 11, 20) {real, imag} */,
  {32'h3f1bbb79, 32'h00000000} /* (15, 11, 19) {real, imag} */,
  {32'h3f4d6fb8, 32'h00000000} /* (15, 11, 18) {real, imag} */,
  {32'h3f7fc0db, 32'h00000000} /* (15, 11, 17) {real, imag} */,
  {32'h3f5477f1, 32'h00000000} /* (15, 11, 16) {real, imag} */,
  {32'h3e92b57e, 32'h00000000} /* (15, 11, 15) {real, imag} */,
  {32'h3ef3baba, 32'h00000000} /* (15, 11, 14) {real, imag} */,
  {32'h3ef94fc1, 32'h00000000} /* (15, 11, 13) {real, imag} */,
  {32'h3f1dfca6, 32'h00000000} /* (15, 11, 12) {real, imag} */,
  {32'h3f7f3676, 32'h00000000} /* (15, 11, 11) {real, imag} */,
  {32'hbe401582, 32'h00000000} /* (15, 11, 10) {real, imag} */,
  {32'hbec175f9, 32'h00000000} /* (15, 11, 9) {real, imag} */,
  {32'hbf0cc7dc, 32'h00000000} /* (15, 11, 8) {real, imag} */,
  {32'hbea9ec24, 32'h00000000} /* (15, 11, 7) {real, imag} */,
  {32'h3dee40e8, 32'h00000000} /* (15, 11, 6) {real, imag} */,
  {32'h3d004e14, 32'h00000000} /* (15, 11, 5) {real, imag} */,
  {32'hbe88ea3e, 32'h00000000} /* (15, 11, 4) {real, imag} */,
  {32'hbd807e67, 32'h00000000} /* (15, 11, 3) {real, imag} */,
  {32'h3db5c9ed, 32'h00000000} /* (15, 11, 2) {real, imag} */,
  {32'hbe69f13d, 32'h00000000} /* (15, 11, 1) {real, imag} */,
  {32'hbd46fab9, 32'h00000000} /* (15, 11, 0) {real, imag} */,
  {32'h3ea778cd, 32'h00000000} /* (15, 10, 31) {real, imag} */,
  {32'h3f42a852, 32'h00000000} /* (15, 10, 30) {real, imag} */,
  {32'h3f764871, 32'h00000000} /* (15, 10, 29) {real, imag} */,
  {32'h3eea32a4, 32'h00000000} /* (15, 10, 28) {real, imag} */,
  {32'h3da8f6e0, 32'h00000000} /* (15, 10, 27) {real, imag} */,
  {32'h3e44c7f5, 32'h00000000} /* (15, 10, 26) {real, imag} */,
  {32'hbd92499f, 32'h00000000} /* (15, 10, 25) {real, imag} */,
  {32'hbeafd0b5, 32'h00000000} /* (15, 10, 24) {real, imag} */,
  {32'hbf5c73db, 32'h00000000} /* (15, 10, 23) {real, imag} */,
  {32'h3f2febcf, 32'h00000000} /* (15, 10, 22) {real, imag} */,
  {32'h3e9eee73, 32'h00000000} /* (15, 10, 21) {real, imag} */,
  {32'hbd165296, 32'h00000000} /* (15, 10, 20) {real, imag} */,
  {32'hbe6c6f0a, 32'h00000000} /* (15, 10, 19) {real, imag} */,
  {32'h3e6f0f84, 32'h00000000} /* (15, 10, 18) {real, imag} */,
  {32'h3e8c70b1, 32'h00000000} /* (15, 10, 17) {real, imag} */,
  {32'h3d43169d, 32'h00000000} /* (15, 10, 16) {real, imag} */,
  {32'hbeb03fb6, 32'h00000000} /* (15, 10, 15) {real, imag} */,
  {32'h3c1f39e6, 32'h00000000} /* (15, 10, 14) {real, imag} */,
  {32'hbe76fa93, 32'h00000000} /* (15, 10, 13) {real, imag} */,
  {32'hbe8a0cb9, 32'h00000000} /* (15, 10, 12) {real, imag} */,
  {32'hbd93e97b, 32'h00000000} /* (15, 10, 11) {real, imag} */,
  {32'hbe17e484, 32'h00000000} /* (15, 10, 10) {real, imag} */,
  {32'h3e22d14c, 32'h00000000} /* (15, 10, 9) {real, imag} */,
  {32'h3e9f8579, 32'h00000000} /* (15, 10, 8) {real, imag} */,
  {32'h3e768f22, 32'h00000000} /* (15, 10, 7) {real, imag} */,
  {32'h3eea7ee9, 32'h00000000} /* (15, 10, 6) {real, imag} */,
  {32'h3f44e86f, 32'h00000000} /* (15, 10, 5) {real, imag} */,
  {32'h3e511147, 32'h00000000} /* (15, 10, 4) {real, imag} */,
  {32'h3f1d3597, 32'h00000000} /* (15, 10, 3) {real, imag} */,
  {32'h3f6dd118, 32'h00000000} /* (15, 10, 2) {real, imag} */,
  {32'h3f070868, 32'h00000000} /* (15, 10, 1) {real, imag} */,
  {32'h3ed0a265, 32'h00000000} /* (15, 10, 0) {real, imag} */,
  {32'h3e3e8d05, 32'h00000000} /* (15, 9, 31) {real, imag} */,
  {32'h3eb486bf, 32'h00000000} /* (15, 9, 30) {real, imag} */,
  {32'h3f437b40, 32'h00000000} /* (15, 9, 29) {real, imag} */,
  {32'h3f80877b, 32'h00000000} /* (15, 9, 28) {real, imag} */,
  {32'h3f0d1cec, 32'h00000000} /* (15, 9, 27) {real, imag} */,
  {32'h3f4978ed, 32'h00000000} /* (15, 9, 26) {real, imag} */,
  {32'h3e4c6205, 32'h00000000} /* (15, 9, 25) {real, imag} */,
  {32'h3e24e3f3, 32'h00000000} /* (15, 9, 24) {real, imag} */,
  {32'h3e6276a8, 32'h00000000} /* (15, 9, 23) {real, imag} */,
  {32'h3f5eb49e, 32'h00000000} /* (15, 9, 22) {real, imag} */,
  {32'h3ecda20d, 32'h00000000} /* (15, 9, 21) {real, imag} */,
  {32'hbeb7c8c7, 32'h00000000} /* (15, 9, 20) {real, imag} */,
  {32'hbeadc538, 32'h00000000} /* (15, 9, 19) {real, imag} */,
  {32'hbeae4a6d, 32'h00000000} /* (15, 9, 18) {real, imag} */,
  {32'hbc7f82dc, 32'h00000000} /* (15, 9, 17) {real, imag} */,
  {32'h3e8e061f, 32'h00000000} /* (15, 9, 16) {real, imag} */,
  {32'hbf49b1d9, 32'h00000000} /* (15, 9, 15) {real, imag} */,
  {32'hbed8d92f, 32'h00000000} /* (15, 9, 14) {real, imag} */,
  {32'hbeb4d3e0, 32'h00000000} /* (15, 9, 13) {real, imag} */,
  {32'hbe6392fd, 32'h00000000} /* (15, 9, 12) {real, imag} */,
  {32'hbeb017f9, 32'h00000000} /* (15, 9, 11) {real, imag} */,
  {32'hbdf35f96, 32'h00000000} /* (15, 9, 10) {real, imag} */,
  {32'h3e8f79e9, 32'h00000000} /* (15, 9, 9) {real, imag} */,
  {32'h3dd4f4b7, 32'h00000000} /* (15, 9, 8) {real, imag} */,
  {32'h3e0bf3b8, 32'h00000000} /* (15, 9, 7) {real, imag} */,
  {32'h3f7b7a7c, 32'h00000000} /* (15, 9, 6) {real, imag} */,
  {32'h3f51caaa, 32'h00000000} /* (15, 9, 5) {real, imag} */,
  {32'h3f4f2ac8, 32'h00000000} /* (15, 9, 4) {real, imag} */,
  {32'h3f790bdf, 32'h00000000} /* (15, 9, 3) {real, imag} */,
  {32'h3f4828d3, 32'h00000000} /* (15, 9, 2) {real, imag} */,
  {32'h3f2972be, 32'h00000000} /* (15, 9, 1) {real, imag} */,
  {32'h3ecf2f36, 32'h00000000} /* (15, 9, 0) {real, imag} */,
  {32'h3c92ab82, 32'h00000000} /* (15, 8, 31) {real, imag} */,
  {32'h3f2ccae9, 32'h00000000} /* (15, 8, 30) {real, imag} */,
  {32'h3f2eb8b3, 32'h00000000} /* (15, 8, 29) {real, imag} */,
  {32'h3f219690, 32'h00000000} /* (15, 8, 28) {real, imag} */,
  {32'h3f300dfa, 32'h00000000} /* (15, 8, 27) {real, imag} */,
  {32'h3f4770c3, 32'h00000000} /* (15, 8, 26) {real, imag} */,
  {32'h3e90bfad, 32'h00000000} /* (15, 8, 25) {real, imag} */,
  {32'h3edf6e6a, 32'h00000000} /* (15, 8, 24) {real, imag} */,
  {32'h3ebb7dfc, 32'h00000000} /* (15, 8, 23) {real, imag} */,
  {32'h3f56e488, 32'h00000000} /* (15, 8, 22) {real, imag} */,
  {32'h3f6ad4aa, 32'h00000000} /* (15, 8, 21) {real, imag} */,
  {32'hbe1e7364, 32'h00000000} /* (15, 8, 20) {real, imag} */,
  {32'hbe572ba6, 32'h00000000} /* (15, 8, 19) {real, imag} */,
  {32'hbf012458, 32'h00000000} /* (15, 8, 18) {real, imag} */,
  {32'h3d274d4e, 32'h00000000} /* (15, 8, 17) {real, imag} */,
  {32'h3e2709e7, 32'h00000000} /* (15, 8, 16) {real, imag} */,
  {32'hbf1c2804, 32'h00000000} /* (15, 8, 15) {real, imag} */,
  {32'hbeaf6d71, 32'h00000000} /* (15, 8, 14) {real, imag} */,
  {32'hbedf4478, 32'h00000000} /* (15, 8, 13) {real, imag} */,
  {32'hbf3e9c20, 32'h00000000} /* (15, 8, 12) {real, imag} */,
  {32'hbf152a66, 32'h00000000} /* (15, 8, 11) {real, imag} */,
  {32'h3e27af9a, 32'h00000000} /* (15, 8, 10) {real, imag} */,
  {32'h3ed290a3, 32'h00000000} /* (15, 8, 9) {real, imag} */,
  {32'h3ead9564, 32'h00000000} /* (15, 8, 8) {real, imag} */,
  {32'h3ec69f15, 32'h00000000} /* (15, 8, 7) {real, imag} */,
  {32'h3fae8d84, 32'h00000000} /* (15, 8, 6) {real, imag} */,
  {32'h3f3ebf88, 32'h00000000} /* (15, 8, 5) {real, imag} */,
  {32'h3f106da2, 32'h00000000} /* (15, 8, 4) {real, imag} */,
  {32'h3f349384, 32'h00000000} /* (15, 8, 3) {real, imag} */,
  {32'h3e971940, 32'h00000000} /* (15, 8, 2) {real, imag} */,
  {32'h3e16111c, 32'h00000000} /* (15, 8, 1) {real, imag} */,
  {32'h3c4faa30, 32'h00000000} /* (15, 8, 0) {real, imag} */,
  {32'h3eee8e90, 32'h00000000} /* (15, 7, 31) {real, imag} */,
  {32'h3f60b843, 32'h00000000} /* (15, 7, 30) {real, imag} */,
  {32'h3f57dcec, 32'h00000000} /* (15, 7, 29) {real, imag} */,
  {32'h3ed4206a, 32'h00000000} /* (15, 7, 28) {real, imag} */,
  {32'h3e70f836, 32'h00000000} /* (15, 7, 27) {real, imag} */,
  {32'h3ee31180, 32'h00000000} /* (15, 7, 26) {real, imag} */,
  {32'h3e4b7e6b, 32'h00000000} /* (15, 7, 25) {real, imag} */,
  {32'h3e8f9abb, 32'h00000000} /* (15, 7, 24) {real, imag} */,
  {32'h3ef087db, 32'h00000000} /* (15, 7, 23) {real, imag} */,
  {32'h3f5d497d, 32'h00000000} /* (15, 7, 22) {real, imag} */,
  {32'h3f0d1f90, 32'h00000000} /* (15, 7, 21) {real, imag} */,
  {32'hbee4396c, 32'h00000000} /* (15, 7, 20) {real, imag} */,
  {32'hbefb78f9, 32'h00000000} /* (15, 7, 19) {real, imag} */,
  {32'hbf0ce455, 32'h00000000} /* (15, 7, 18) {real, imag} */,
  {32'hbdafbc17, 32'h00000000} /* (15, 7, 17) {real, imag} */,
  {32'hbea791e7, 32'h00000000} /* (15, 7, 16) {real, imag} */,
  {32'hbefd1497, 32'h00000000} /* (15, 7, 15) {real, imag} */,
  {32'hbeb16aa5, 32'h00000000} /* (15, 7, 14) {real, imag} */,
  {32'hbedfdd2d, 32'h00000000} /* (15, 7, 13) {real, imag} */,
  {32'hbf1ca727, 32'h00000000} /* (15, 7, 12) {real, imag} */,
  {32'h3e0e2398, 32'h00000000} /* (15, 7, 11) {real, imag} */,
  {32'h3f2fa7bf, 32'h00000000} /* (15, 7, 10) {real, imag} */,
  {32'h3eb68371, 32'h00000000} /* (15, 7, 9) {real, imag} */,
  {32'h3f63d18d, 32'h00000000} /* (15, 7, 8) {real, imag} */,
  {32'h3f590afc, 32'h00000000} /* (15, 7, 7) {real, imag} */,
  {32'h3f3f510d, 32'h00000000} /* (15, 7, 6) {real, imag} */,
  {32'h3f7dd506, 32'h00000000} /* (15, 7, 5) {real, imag} */,
  {32'h3f1bbe8a, 32'h00000000} /* (15, 7, 4) {real, imag} */,
  {32'h3f00385e, 32'h00000000} /* (15, 7, 3) {real, imag} */,
  {32'h3e1dd883, 32'h00000000} /* (15, 7, 2) {real, imag} */,
  {32'h3e9fe4bb, 32'h00000000} /* (15, 7, 1) {real, imag} */,
  {32'h3eb3989d, 32'h00000000} /* (15, 7, 0) {real, imag} */,
  {32'h3ea89323, 32'h00000000} /* (15, 6, 31) {real, imag} */,
  {32'h3f06a401, 32'h00000000} /* (15, 6, 30) {real, imag} */,
  {32'h3d13df4e, 32'h00000000} /* (15, 6, 29) {real, imag} */,
  {32'h3d8ef425, 32'h00000000} /* (15, 6, 28) {real, imag} */,
  {32'h3e906b7f, 32'h00000000} /* (15, 6, 27) {real, imag} */,
  {32'h3f0d4e0f, 32'h00000000} /* (15, 6, 26) {real, imag} */,
  {32'h3e7ea9e0, 32'h00000000} /* (15, 6, 25) {real, imag} */,
  {32'h3f0fca56, 32'h00000000} /* (15, 6, 24) {real, imag} */,
  {32'h3f28cef6, 32'h00000000} /* (15, 6, 23) {real, imag} */,
  {32'h3f30aa82, 32'h00000000} /* (15, 6, 22) {real, imag} */,
  {32'h3f06931d, 32'h00000000} /* (15, 6, 21) {real, imag} */,
  {32'hbe144979, 32'h00000000} /* (15, 6, 20) {real, imag} */,
  {32'hbece2bbc, 32'h00000000} /* (15, 6, 19) {real, imag} */,
  {32'hbf16308e, 32'h00000000} /* (15, 6, 18) {real, imag} */,
  {32'hbf231b66, 32'h00000000} /* (15, 6, 17) {real, imag} */,
  {32'hbe9b1c33, 32'h00000000} /* (15, 6, 16) {real, imag} */,
  {32'hbe279098, 32'h00000000} /* (15, 6, 15) {real, imag} */,
  {32'hbe913ed4, 32'h00000000} /* (15, 6, 14) {real, imag} */,
  {32'hbdc799ec, 32'h00000000} /* (15, 6, 13) {real, imag} */,
  {32'hbeed29a6, 32'h00000000} /* (15, 6, 12) {real, imag} */,
  {32'h3d7e1102, 32'h00000000} /* (15, 6, 11) {real, imag} */,
  {32'h3ee9c866, 32'h00000000} /* (15, 6, 10) {real, imag} */,
  {32'h3ec4ad1c, 32'h00000000} /* (15, 6, 9) {real, imag} */,
  {32'h3f3f57cb, 32'h00000000} /* (15, 6, 8) {real, imag} */,
  {32'h3e9873b2, 32'h00000000} /* (15, 6, 7) {real, imag} */,
  {32'h3ec4bf81, 32'h00000000} /* (15, 6, 6) {real, imag} */,
  {32'h3f692d0f, 32'h00000000} /* (15, 6, 5) {real, imag} */,
  {32'h3f84d9ab, 32'h00000000} /* (15, 6, 4) {real, imag} */,
  {32'h3efbc589, 32'h00000000} /* (15, 6, 3) {real, imag} */,
  {32'h3e4ea6d4, 32'h00000000} /* (15, 6, 2) {real, imag} */,
  {32'h3ec4c0c3, 32'h00000000} /* (15, 6, 1) {real, imag} */,
  {32'h3e903e7c, 32'h00000000} /* (15, 6, 0) {real, imag} */,
  {32'h3e7315ca, 32'h00000000} /* (15, 5, 31) {real, imag} */,
  {32'h3f286517, 32'h00000000} /* (15, 5, 30) {real, imag} */,
  {32'h3e8ebaca, 32'h00000000} /* (15, 5, 29) {real, imag} */,
  {32'h3f463fee, 32'h00000000} /* (15, 5, 28) {real, imag} */,
  {32'h3f320654, 32'h00000000} /* (15, 5, 27) {real, imag} */,
  {32'h3e9f0bcc, 32'h00000000} /* (15, 5, 26) {real, imag} */,
  {32'h3e76a9e9, 32'h00000000} /* (15, 5, 25) {real, imag} */,
  {32'h3f7a6cc2, 32'h00000000} /* (15, 5, 24) {real, imag} */,
  {32'h3f007fb0, 32'h00000000} /* (15, 5, 23) {real, imag} */,
  {32'h3ec0cbe4, 32'h00000000} /* (15, 5, 22) {real, imag} */,
  {32'h3e88ccff, 32'h00000000} /* (15, 5, 21) {real, imag} */,
  {32'h3eb6d8f7, 32'h00000000} /* (15, 5, 20) {real, imag} */,
  {32'hbdae7774, 32'h00000000} /* (15, 5, 19) {real, imag} */,
  {32'hbea933c6, 32'h00000000} /* (15, 5, 18) {real, imag} */,
  {32'hbf01e350, 32'h00000000} /* (15, 5, 17) {real, imag} */,
  {32'hbdc46260, 32'h00000000} /* (15, 5, 16) {real, imag} */,
  {32'hbe968f92, 32'h00000000} /* (15, 5, 15) {real, imag} */,
  {32'hbed6773e, 32'h00000000} /* (15, 5, 14) {real, imag} */,
  {32'hbe01ea66, 32'h00000000} /* (15, 5, 13) {real, imag} */,
  {32'hbf2d0ae8, 32'h00000000} /* (15, 5, 12) {real, imag} */,
  {32'hbf6e5224, 32'h00000000} /* (15, 5, 11) {real, imag} */,
  {32'hbf35d597, 32'h00000000} /* (15, 5, 10) {real, imag} */,
  {32'hbd7db128, 32'h00000000} /* (15, 5, 9) {real, imag} */,
  {32'hbe372700, 32'h00000000} /* (15, 5, 8) {real, imag} */,
  {32'hbf0f13de, 32'h00000000} /* (15, 5, 7) {real, imag} */,
  {32'h3e5001c5, 32'h00000000} /* (15, 5, 6) {real, imag} */,
  {32'h3f1f8003, 32'h00000000} /* (15, 5, 5) {real, imag} */,
  {32'h3f9844f5, 32'h00000000} /* (15, 5, 4) {real, imag} */,
  {32'h3eedac39, 32'h00000000} /* (15, 5, 3) {real, imag} */,
  {32'h3de7b59a, 32'h00000000} /* (15, 5, 2) {real, imag} */,
  {32'h3e4612ac, 32'h00000000} /* (15, 5, 1) {real, imag} */,
  {32'h3dcf8f8f, 32'h00000000} /* (15, 5, 0) {real, imag} */,
  {32'h3e6853b8, 32'h00000000} /* (15, 4, 31) {real, imag} */,
  {32'h3f0521b2, 32'h00000000} /* (15, 4, 30) {real, imag} */,
  {32'h3efce060, 32'h00000000} /* (15, 4, 29) {real, imag} */,
  {32'h3f5035ce, 32'h00000000} /* (15, 4, 28) {real, imag} */,
  {32'h3f3a16cb, 32'h00000000} /* (15, 4, 27) {real, imag} */,
  {32'h3efaf1c4, 32'h00000000} /* (15, 4, 26) {real, imag} */,
  {32'h3eb9abc4, 32'h00000000} /* (15, 4, 25) {real, imag} */,
  {32'h3f6fd750, 32'h00000000} /* (15, 4, 24) {real, imag} */,
  {32'h3f1f48f5, 32'h00000000} /* (15, 4, 23) {real, imag} */,
  {32'h3f5a4993, 32'h00000000} /* (15, 4, 22) {real, imag} */,
  {32'h3f40d6f1, 32'h00000000} /* (15, 4, 21) {real, imag} */,
  {32'h3f03afda, 32'h00000000} /* (15, 4, 20) {real, imag} */,
  {32'h3e098eea, 32'h00000000} /* (15, 4, 19) {real, imag} */,
  {32'h3e86614e, 32'h00000000} /* (15, 4, 18) {real, imag} */,
  {32'h3e564e89, 32'h00000000} /* (15, 4, 17) {real, imag} */,
  {32'h3d3b071b, 32'h00000000} /* (15, 4, 16) {real, imag} */,
  {32'hbf14af7d, 32'h00000000} /* (15, 4, 15) {real, imag} */,
  {32'hbea485e9, 32'h00000000} /* (15, 4, 14) {real, imag} */,
  {32'hbecfcb42, 32'h00000000} /* (15, 4, 13) {real, imag} */,
  {32'hbea1cd6c, 32'h00000000} /* (15, 4, 12) {real, imag} */,
  {32'hbf45e3c7, 32'h00000000} /* (15, 4, 11) {real, imag} */,
  {32'hbed7d920, 32'h00000000} /* (15, 4, 10) {real, imag} */,
  {32'hbefea817, 32'h00000000} /* (15, 4, 9) {real, imag} */,
  {32'hbf510989, 32'h00000000} /* (15, 4, 8) {real, imag} */,
  {32'hbf485680, 32'h00000000} /* (15, 4, 7) {real, imag} */,
  {32'hbe505707, 32'h00000000} /* (15, 4, 6) {real, imag} */,
  {32'h3e8ba2d1, 32'h00000000} /* (15, 4, 5) {real, imag} */,
  {32'h3f3aee2f, 32'h00000000} /* (15, 4, 4) {real, imag} */,
  {32'h3f521409, 32'h00000000} /* (15, 4, 3) {real, imag} */,
  {32'h3ec74da4, 32'h00000000} /* (15, 4, 2) {real, imag} */,
  {32'h3eae35c6, 32'h00000000} /* (15, 4, 1) {real, imag} */,
  {32'h3e81e202, 32'h00000000} /* (15, 4, 0) {real, imag} */,
  {32'h3f10ff5d, 32'h00000000} /* (15, 3, 31) {real, imag} */,
  {32'h3f032c46, 32'h00000000} /* (15, 3, 30) {real, imag} */,
  {32'h3ebb037b, 32'h00000000} /* (15, 3, 29) {real, imag} */,
  {32'h3f2a7fb3, 32'h00000000} /* (15, 3, 28) {real, imag} */,
  {32'h3f1f79ea, 32'h00000000} /* (15, 3, 27) {real, imag} */,
  {32'h3f319578, 32'h00000000} /* (15, 3, 26) {real, imag} */,
  {32'h3e8a2073, 32'h00000000} /* (15, 3, 25) {real, imag} */,
  {32'h3eee3332, 32'h00000000} /* (15, 3, 24) {real, imag} */,
  {32'h3ef0a4ce, 32'h00000000} /* (15, 3, 23) {real, imag} */,
  {32'h3f50849a, 32'h00000000} /* (15, 3, 22) {real, imag} */,
  {32'h3f15ae06, 32'h00000000} /* (15, 3, 21) {real, imag} */,
  {32'h3f07d795, 32'h00000000} /* (15, 3, 20) {real, imag} */,
  {32'h3f0465fe, 32'h00000000} /* (15, 3, 19) {real, imag} */,
  {32'h3f35bf28, 32'h00000000} /* (15, 3, 18) {real, imag} */,
  {32'h3ebbb98d, 32'h00000000} /* (15, 3, 17) {real, imag} */,
  {32'h3e8a04ac, 32'h00000000} /* (15, 3, 16) {real, imag} */,
  {32'hbf690551, 32'h00000000} /* (15, 3, 15) {real, imag} */,
  {32'hbf3b8a23, 32'h00000000} /* (15, 3, 14) {real, imag} */,
  {32'hbf24e47b, 32'h00000000} /* (15, 3, 13) {real, imag} */,
  {32'hbef0a09e, 32'h00000000} /* (15, 3, 12) {real, imag} */,
  {32'hbebe7f30, 32'h00000000} /* (15, 3, 11) {real, imag} */,
  {32'hbe219465, 32'h00000000} /* (15, 3, 10) {real, imag} */,
  {32'hbef17c8c, 32'h00000000} /* (15, 3, 9) {real, imag} */,
  {32'hbec9531b, 32'h00000000} /* (15, 3, 8) {real, imag} */,
  {32'hbeaabede, 32'h00000000} /* (15, 3, 7) {real, imag} */,
  {32'hbd13055a, 32'h00000000} /* (15, 3, 6) {real, imag} */,
  {32'h3f597e34, 32'h00000000} /* (15, 3, 5) {real, imag} */,
  {32'h3fb1cc5c, 32'h00000000} /* (15, 3, 4) {real, imag} */,
  {32'h3fad38b8, 32'h00000000} /* (15, 3, 3) {real, imag} */,
  {32'h3eaeeaeb, 32'h00000000} /* (15, 3, 2) {real, imag} */,
  {32'h3e888680, 32'h00000000} /* (15, 3, 1) {real, imag} */,
  {32'h3ef6a9bb, 32'h00000000} /* (15, 3, 0) {real, imag} */,
  {32'h3ef05c08, 32'h00000000} /* (15, 2, 31) {real, imag} */,
  {32'h3f82b97d, 32'h00000000} /* (15, 2, 30) {real, imag} */,
  {32'h3ef5a465, 32'h00000000} /* (15, 2, 29) {real, imag} */,
  {32'h3f16dd49, 32'h00000000} /* (15, 2, 28) {real, imag} */,
  {32'h3ee02e38, 32'h00000000} /* (15, 2, 27) {real, imag} */,
  {32'h3e9122d1, 32'h00000000} /* (15, 2, 26) {real, imag} */,
  {32'h3da027d1, 32'h00000000} /* (15, 2, 25) {real, imag} */,
  {32'h3ee19eb9, 32'h00000000} /* (15, 2, 24) {real, imag} */,
  {32'h3f0bc493, 32'h00000000} /* (15, 2, 23) {real, imag} */,
  {32'h3ed33801, 32'h00000000} /* (15, 2, 22) {real, imag} */,
  {32'h3e88f061, 32'h00000000} /* (15, 2, 21) {real, imag} */,
  {32'h3eb4ceb1, 32'h00000000} /* (15, 2, 20) {real, imag} */,
  {32'h3f27a7d9, 32'h00000000} /* (15, 2, 19) {real, imag} */,
  {32'h3ee52687, 32'h00000000} /* (15, 2, 18) {real, imag} */,
  {32'h3f345ea2, 32'h00000000} /* (15, 2, 17) {real, imag} */,
  {32'h3f79a144, 32'h00000000} /* (15, 2, 16) {real, imag} */,
  {32'hbefb25d0, 32'h00000000} /* (15, 2, 15) {real, imag} */,
  {32'hbf444f80, 32'h00000000} /* (15, 2, 14) {real, imag} */,
  {32'hbf1e5876, 32'h00000000} /* (15, 2, 13) {real, imag} */,
  {32'hbf19b450, 32'h00000000} /* (15, 2, 12) {real, imag} */,
  {32'hbf2f8c09, 32'h00000000} /* (15, 2, 11) {real, imag} */,
  {32'hbec08b95, 32'h00000000} /* (15, 2, 10) {real, imag} */,
  {32'hbebc7e1a, 32'h00000000} /* (15, 2, 9) {real, imag} */,
  {32'hbde35737, 32'h00000000} /* (15, 2, 8) {real, imag} */,
  {32'hbe525bd0, 32'h00000000} /* (15, 2, 7) {real, imag} */,
  {32'hbe95163c, 32'h00000000} /* (15, 2, 6) {real, imag} */,
  {32'h3f107604, 32'h00000000} /* (15, 2, 5) {real, imag} */,
  {32'h3f6c0a27, 32'h00000000} /* (15, 2, 4) {real, imag} */,
  {32'h3f7737e8, 32'h00000000} /* (15, 2, 3) {real, imag} */,
  {32'h3f27acd6, 32'h00000000} /* (15, 2, 2) {real, imag} */,
  {32'h3e94846b, 32'h00000000} /* (15, 2, 1) {real, imag} */,
  {32'h3e5c460f, 32'h00000000} /* (15, 2, 0) {real, imag} */,
  {32'h3dfbded8, 32'h00000000} /* (15, 1, 31) {real, imag} */,
  {32'h3f06df44, 32'h00000000} /* (15, 1, 30) {real, imag} */,
  {32'h3ebd6eb5, 32'h00000000} /* (15, 1, 29) {real, imag} */,
  {32'h3ee4c001, 32'h00000000} /* (15, 1, 28) {real, imag} */,
  {32'h3f02a64b, 32'h00000000} /* (15, 1, 27) {real, imag} */,
  {32'h3e45fff9, 32'h00000000} /* (15, 1, 26) {real, imag} */,
  {32'h3e7250c6, 32'h00000000} /* (15, 1, 25) {real, imag} */,
  {32'h3e749e81, 32'h00000000} /* (15, 1, 24) {real, imag} */,
  {32'h3f0f7a47, 32'h00000000} /* (15, 1, 23) {real, imag} */,
  {32'h3f25dd03, 32'h00000000} /* (15, 1, 22) {real, imag} */,
  {32'h3ebfb4a2, 32'h00000000} /* (15, 1, 21) {real, imag} */,
  {32'h3f0b8753, 32'h00000000} /* (15, 1, 20) {real, imag} */,
  {32'h3f23eea4, 32'h00000000} /* (15, 1, 19) {real, imag} */,
  {32'h3e14b741, 32'h00000000} /* (15, 1, 18) {real, imag} */,
  {32'h3f1cc51a, 32'h00000000} /* (15, 1, 17) {real, imag} */,
  {32'h3ef05477, 32'h00000000} /* (15, 1, 16) {real, imag} */,
  {32'hbf06be5e, 32'h00000000} /* (15, 1, 15) {real, imag} */,
  {32'hbf549966, 32'h00000000} /* (15, 1, 14) {real, imag} */,
  {32'hbf06157a, 32'h00000000} /* (15, 1, 13) {real, imag} */,
  {32'hbec6e7e0, 32'h00000000} /* (15, 1, 12) {real, imag} */,
  {32'hbf314d4c, 32'h00000000} /* (15, 1, 11) {real, imag} */,
  {32'hbf788f2b, 32'h00000000} /* (15, 1, 10) {real, imag} */,
  {32'hbf5b0756, 32'h00000000} /* (15, 1, 9) {real, imag} */,
  {32'hbf229436, 32'h00000000} /* (15, 1, 8) {real, imag} */,
  {32'hbf165605, 32'h00000000} /* (15, 1, 7) {real, imag} */,
  {32'hbf7bf4ad, 32'h00000000} /* (15, 1, 6) {real, imag} */,
  {32'hbf10a593, 32'h00000000} /* (15, 1, 5) {real, imag} */,
  {32'hbd5358e5, 32'h00000000} /* (15, 1, 4) {real, imag} */,
  {32'h3e9fb5ae, 32'h00000000} /* (15, 1, 3) {real, imag} */,
  {32'h3f2dd117, 32'h00000000} /* (15, 1, 2) {real, imag} */,
  {32'h3e8a12ec, 32'h00000000} /* (15, 1, 1) {real, imag} */,
  {32'hbe680fdd, 32'h00000000} /* (15, 1, 0) {real, imag} */,
  {32'h3c85e1eb, 32'h00000000} /* (15, 0, 31) {real, imag} */,
  {32'h3e0344ef, 32'h00000000} /* (15, 0, 30) {real, imag} */,
  {32'h3e39afbb, 32'h00000000} /* (15, 0, 29) {real, imag} */,
  {32'h3eac1dfc, 32'h00000000} /* (15, 0, 28) {real, imag} */,
  {32'h3e96b5b0, 32'h00000000} /* (15, 0, 27) {real, imag} */,
  {32'h3dc923ed, 32'h00000000} /* (15, 0, 26) {real, imag} */,
  {32'h3d3339c9, 32'h00000000} /* (15, 0, 25) {real, imag} */,
  {32'hbd0946cd, 32'h00000000} /* (15, 0, 24) {real, imag} */,
  {32'h3efa5e41, 32'h00000000} /* (15, 0, 23) {real, imag} */,
  {32'h3eb0349c, 32'h00000000} /* (15, 0, 22) {real, imag} */,
  {32'h3d1aafdf, 32'h00000000} /* (15, 0, 21) {real, imag} */,
  {32'h3d5faa17, 32'h00000000} /* (15, 0, 20) {real, imag} */,
  {32'h3de63809, 32'h00000000} /* (15, 0, 19) {real, imag} */,
  {32'h3d001a00, 32'h00000000} /* (15, 0, 18) {real, imag} */,
  {32'h3e4257e4, 32'h00000000} /* (15, 0, 17) {real, imag} */,
  {32'h3e43a55f, 32'h00000000} /* (15, 0, 16) {real, imag} */,
  {32'hbed0729c, 32'h00000000} /* (15, 0, 15) {real, imag} */,
  {32'hbf49f3ee, 32'h00000000} /* (15, 0, 14) {real, imag} */,
  {32'hbf3d20da, 32'h00000000} /* (15, 0, 13) {real, imag} */,
  {32'hbe8bf8a1, 32'h00000000} /* (15, 0, 12) {real, imag} */,
  {32'hbeb5d754, 32'h00000000} /* (15, 0, 11) {real, imag} */,
  {32'hbf196241, 32'h00000000} /* (15, 0, 10) {real, imag} */,
  {32'hbef1444a, 32'h00000000} /* (15, 0, 9) {real, imag} */,
  {32'hbedd4fad, 32'h00000000} /* (15, 0, 8) {real, imag} */,
  {32'hbeb9ecb3, 32'h00000000} /* (15, 0, 7) {real, imag} */,
  {32'hbeace204, 32'h00000000} /* (15, 0, 6) {real, imag} */,
  {32'hbe508197, 32'h00000000} /* (15, 0, 5) {real, imag} */,
  {32'hbb3369a8, 32'h00000000} /* (15, 0, 4) {real, imag} */,
  {32'h3ee4263f, 32'h00000000} /* (15, 0, 3) {real, imag} */,
  {32'h3f38870a, 32'h00000000} /* (15, 0, 2) {real, imag} */,
  {32'h3e1bc28a, 32'h00000000} /* (15, 0, 1) {real, imag} */,
  {32'hbe796f6d, 32'h00000000} /* (15, 0, 0) {real, imag} */,
  {32'h3e8c6e3f, 32'h00000000} /* (14, 31, 31) {real, imag} */,
  {32'h3f183f22, 32'h00000000} /* (14, 31, 30) {real, imag} */,
  {32'h3f2aaa04, 32'h00000000} /* (14, 31, 29) {real, imag} */,
  {32'h3f0ec80d, 32'h00000000} /* (14, 31, 28) {real, imag} */,
  {32'h3f0fc123, 32'h00000000} /* (14, 31, 27) {real, imag} */,
  {32'h3f4abb05, 32'h00000000} /* (14, 31, 26) {real, imag} */,
  {32'h3f2d45e8, 32'h00000000} /* (14, 31, 25) {real, imag} */,
  {32'h3f794f9a, 32'h00000000} /* (14, 31, 24) {real, imag} */,
  {32'h3f12c8e2, 32'h00000000} /* (14, 31, 23) {real, imag} */,
  {32'h3f17d53a, 32'h00000000} /* (14, 31, 22) {real, imag} */,
  {32'h3de20f6b, 32'h00000000} /* (14, 31, 21) {real, imag} */,
  {32'hbdc497dd, 32'h00000000} /* (14, 31, 20) {real, imag} */,
  {32'hbd94eb3a, 32'h00000000} /* (14, 31, 19) {real, imag} */,
  {32'hbedff9aa, 32'h00000000} /* (14, 31, 18) {real, imag} */,
  {32'hbf3cc164, 32'h00000000} /* (14, 31, 17) {real, imag} */,
  {32'hbe881119, 32'h00000000} /* (14, 31, 16) {real, imag} */,
  {32'hbee89e74, 32'h00000000} /* (14, 31, 15) {real, imag} */,
  {32'hbf18e329, 32'h00000000} /* (14, 31, 14) {real, imag} */,
  {32'hbf0c1552, 32'h00000000} /* (14, 31, 13) {real, imag} */,
  {32'hbee7ec12, 32'h00000000} /* (14, 31, 12) {real, imag} */,
  {32'hbf1681c6, 32'h00000000} /* (14, 31, 11) {real, imag} */,
  {32'hbe965d99, 32'h00000000} /* (14, 31, 10) {real, imag} */,
  {32'h3da0eff0, 32'h00000000} /* (14, 31, 9) {real, imag} */,
  {32'hbc7f62e9, 32'h00000000} /* (14, 31, 8) {real, imag} */,
  {32'h3db0638a, 32'h00000000} /* (14, 31, 7) {real, imag} */,
  {32'h3ed74285, 32'h00000000} /* (14, 31, 6) {real, imag} */,
  {32'h3eec7872, 32'h00000000} /* (14, 31, 5) {real, imag} */,
  {32'h3e64c2f0, 32'h00000000} /* (14, 31, 4) {real, imag} */,
  {32'h3e73971b, 32'h00000000} /* (14, 31, 3) {real, imag} */,
  {32'h3ee21369, 32'h00000000} /* (14, 31, 2) {real, imag} */,
  {32'h3f007987, 32'h00000000} /* (14, 31, 1) {real, imag} */,
  {32'h3e8e761b, 32'h00000000} /* (14, 31, 0) {real, imag} */,
  {32'h3ed737ca, 32'h00000000} /* (14, 30, 31) {real, imag} */,
  {32'h3f3d99d5, 32'h00000000} /* (14, 30, 30) {real, imag} */,
  {32'h3f274361, 32'h00000000} /* (14, 30, 29) {real, imag} */,
  {32'h3f2288d3, 32'h00000000} /* (14, 30, 28) {real, imag} */,
  {32'h3f529f53, 32'h00000000} /* (14, 30, 27) {real, imag} */,
  {32'h3fbfcb1e, 32'h00000000} /* (14, 30, 26) {real, imag} */,
  {32'h3fd47c5f, 32'h00000000} /* (14, 30, 25) {real, imag} */,
  {32'h3fe9c848, 32'h00000000} /* (14, 30, 24) {real, imag} */,
  {32'h3fa1e43b, 32'h00000000} /* (14, 30, 23) {real, imag} */,
  {32'h3f4443c0, 32'h00000000} /* (14, 30, 22) {real, imag} */,
  {32'h3dde919e, 32'h00000000} /* (14, 30, 21) {real, imag} */,
  {32'hbee21b82, 32'h00000000} /* (14, 30, 20) {real, imag} */,
  {32'hbf2b012b, 32'h00000000} /* (14, 30, 19) {real, imag} */,
  {32'hbfc1290a, 32'h00000000} /* (14, 30, 18) {real, imag} */,
  {32'hbfb0736e, 32'h00000000} /* (14, 30, 17) {real, imag} */,
  {32'hbf44f789, 32'h00000000} /* (14, 30, 16) {real, imag} */,
  {32'hbf979541, 32'h00000000} /* (14, 30, 15) {real, imag} */,
  {32'hbf999d49, 32'h00000000} /* (14, 30, 14) {real, imag} */,
  {32'hbf7e6e95, 32'h00000000} /* (14, 30, 13) {real, imag} */,
  {32'hbf94ce13, 32'h00000000} /* (14, 30, 12) {real, imag} */,
  {32'hbf4bcf31, 32'h00000000} /* (14, 30, 11) {real, imag} */,
  {32'h3e411b61, 32'h00000000} /* (14, 30, 10) {real, imag} */,
  {32'h3f4205b7, 32'h00000000} /* (14, 30, 9) {real, imag} */,
  {32'h3eb97be9, 32'h00000000} /* (14, 30, 8) {real, imag} */,
  {32'h3e77c240, 32'h00000000} /* (14, 30, 7) {real, imag} */,
  {32'h3f265df7, 32'h00000000} /* (14, 30, 6) {real, imag} */,
  {32'h3f2bdee7, 32'h00000000} /* (14, 30, 5) {real, imag} */,
  {32'h3eb6b129, 32'h00000000} /* (14, 30, 4) {real, imag} */,
  {32'h3e9aaf55, 32'h00000000} /* (14, 30, 3) {real, imag} */,
  {32'h3ebb41ed, 32'h00000000} /* (14, 30, 2) {real, imag} */,
  {32'h3f92b160, 32'h00000000} /* (14, 30, 1) {real, imag} */,
  {32'h3f770a43, 32'h00000000} /* (14, 30, 0) {real, imag} */,
  {32'h3edec036, 32'h00000000} /* (14, 29, 31) {real, imag} */,
  {32'h3f469c45, 32'h00000000} /* (14, 29, 30) {real, imag} */,
  {32'h3f012a6d, 32'h00000000} /* (14, 29, 29) {real, imag} */,
  {32'h3f3a1a98, 32'h00000000} /* (14, 29, 28) {real, imag} */,
  {32'h3f7e196b, 32'h00000000} /* (14, 29, 27) {real, imag} */,
  {32'h3f5c645f, 32'h00000000} /* (14, 29, 26) {real, imag} */,
  {32'h3f4a6bea, 32'h00000000} /* (14, 29, 25) {real, imag} */,
  {32'h3f5145d6, 32'h00000000} /* (14, 29, 24) {real, imag} */,
  {32'h3f67d9ea, 32'h00000000} /* (14, 29, 23) {real, imag} */,
  {32'h3eb0f93f, 32'h00000000} /* (14, 29, 22) {real, imag} */,
  {32'h3c5dfb89, 32'h00000000} /* (14, 29, 21) {real, imag} */,
  {32'hbf17dcbc, 32'h00000000} /* (14, 29, 20) {real, imag} */,
  {32'hbf2eca3b, 32'h00000000} /* (14, 29, 19) {real, imag} */,
  {32'hbf89e46d, 32'h00000000} /* (14, 29, 18) {real, imag} */,
  {32'hbf887874, 32'h00000000} /* (14, 29, 17) {real, imag} */,
  {32'hbf97e4b4, 32'h00000000} /* (14, 29, 16) {real, imag} */,
  {32'hbf90f4e9, 32'h00000000} /* (14, 29, 15) {real, imag} */,
  {32'hbf74b27e, 32'h00000000} /* (14, 29, 14) {real, imag} */,
  {32'hbf0e6983, 32'h00000000} /* (14, 29, 13) {real, imag} */,
  {32'hbf298055, 32'h00000000} /* (14, 29, 12) {real, imag} */,
  {32'hbf01076a, 32'h00000000} /* (14, 29, 11) {real, imag} */,
  {32'h3ee57bc3, 32'h00000000} /* (14, 29, 10) {real, imag} */,
  {32'h3f501d83, 32'h00000000} /* (14, 29, 9) {real, imag} */,
  {32'h3ee01848, 32'h00000000} /* (14, 29, 8) {real, imag} */,
  {32'h3e7557b8, 32'h00000000} /* (14, 29, 7) {real, imag} */,
  {32'h3f14e4ee, 32'h00000000} /* (14, 29, 6) {real, imag} */,
  {32'h3f9fb0e2, 32'h00000000} /* (14, 29, 5) {real, imag} */,
  {32'h3f42930b, 32'h00000000} /* (14, 29, 4) {real, imag} */,
  {32'h3eaf62a1, 32'h00000000} /* (14, 29, 3) {real, imag} */,
  {32'h3eddee4d, 32'h00000000} /* (14, 29, 2) {real, imag} */,
  {32'h3fc92c53, 32'h00000000} /* (14, 29, 1) {real, imag} */,
  {32'h3f85aca1, 32'h00000000} /* (14, 29, 0) {real, imag} */,
  {32'h3e8c3e7a, 32'h00000000} /* (14, 28, 31) {real, imag} */,
  {32'h3f2ea413, 32'h00000000} /* (14, 28, 30) {real, imag} */,
  {32'h3f21dba3, 32'h00000000} /* (14, 28, 29) {real, imag} */,
  {32'h3f7e9fd9, 32'h00000000} /* (14, 28, 28) {real, imag} */,
  {32'h3f813f09, 32'h00000000} /* (14, 28, 27) {real, imag} */,
  {32'h3f1b20d6, 32'h00000000} /* (14, 28, 26) {real, imag} */,
  {32'h3e97826c, 32'h00000000} /* (14, 28, 25) {real, imag} */,
  {32'h3f009d6f, 32'h00000000} /* (14, 28, 24) {real, imag} */,
  {32'h3f30a13a, 32'h00000000} /* (14, 28, 23) {real, imag} */,
  {32'h3f395c3a, 32'h00000000} /* (14, 28, 22) {real, imag} */,
  {32'h3f0e6310, 32'h00000000} /* (14, 28, 21) {real, imag} */,
  {32'hbe91b5fa, 32'h00000000} /* (14, 28, 20) {real, imag} */,
  {32'hbef1c36b, 32'h00000000} /* (14, 28, 19) {real, imag} */,
  {32'hbf5fb0cc, 32'h00000000} /* (14, 28, 18) {real, imag} */,
  {32'hbf88ea33, 32'h00000000} /* (14, 28, 17) {real, imag} */,
  {32'hbf988c89, 32'h00000000} /* (14, 28, 16) {real, imag} */,
  {32'hbf19d775, 32'h00000000} /* (14, 28, 15) {real, imag} */,
  {32'hbf25aa2d, 32'h00000000} /* (14, 28, 14) {real, imag} */,
  {32'hbe9aa45b, 32'h00000000} /* (14, 28, 13) {real, imag} */,
  {32'hbe634e1e, 32'h00000000} /* (14, 28, 12) {real, imag} */,
  {32'hbf44eda7, 32'h00000000} /* (14, 28, 11) {real, imag} */,
  {32'h3ea97db2, 32'h00000000} /* (14, 28, 10) {real, imag} */,
  {32'h3fa2b842, 32'h00000000} /* (14, 28, 9) {real, imag} */,
  {32'h3f861c2d, 32'h00000000} /* (14, 28, 8) {real, imag} */,
  {32'h3eff28d8, 32'h00000000} /* (14, 28, 7) {real, imag} */,
  {32'h3f51cf49, 32'h00000000} /* (14, 28, 6) {real, imag} */,
  {32'h3f938adc, 32'h00000000} /* (14, 28, 5) {real, imag} */,
  {32'h3f0754ef, 32'h00000000} /* (14, 28, 4) {real, imag} */,
  {32'h3ebc622c, 32'h00000000} /* (14, 28, 3) {real, imag} */,
  {32'h3eedeb09, 32'h00000000} /* (14, 28, 2) {real, imag} */,
  {32'h3f3c8894, 32'h00000000} /* (14, 28, 1) {real, imag} */,
  {32'h3f0a2dfb, 32'h00000000} /* (14, 28, 0) {real, imag} */,
  {32'h3e6a9621, 32'h00000000} /* (14, 27, 31) {real, imag} */,
  {32'h3f938d04, 32'h00000000} /* (14, 27, 30) {real, imag} */,
  {32'h3f9cd4f6, 32'h00000000} /* (14, 27, 29) {real, imag} */,
  {32'h3f843d7e, 32'h00000000} /* (14, 27, 28) {real, imag} */,
  {32'h3f1d764d, 32'h00000000} /* (14, 27, 27) {real, imag} */,
  {32'h3f0882c6, 32'h00000000} /* (14, 27, 26) {real, imag} */,
  {32'h3f33df63, 32'h00000000} /* (14, 27, 25) {real, imag} */,
  {32'h3f4dec7b, 32'h00000000} /* (14, 27, 24) {real, imag} */,
  {32'h3f29816a, 32'h00000000} /* (14, 27, 23) {real, imag} */,
  {32'h3faf0230, 32'h00000000} /* (14, 27, 22) {real, imag} */,
  {32'h3fa4a5f2, 32'h00000000} /* (14, 27, 21) {real, imag} */,
  {32'hbe0229f3, 32'h00000000} /* (14, 27, 20) {real, imag} */,
  {32'hbeea55b7, 32'h00000000} /* (14, 27, 19) {real, imag} */,
  {32'hbf2dc550, 32'h00000000} /* (14, 27, 18) {real, imag} */,
  {32'hbf35ce3c, 32'h00000000} /* (14, 27, 17) {real, imag} */,
  {32'hbf54b742, 32'h00000000} /* (14, 27, 16) {real, imag} */,
  {32'hbef9cdeb, 32'h00000000} /* (14, 27, 15) {real, imag} */,
  {32'hbf2035ce, 32'h00000000} /* (14, 27, 14) {real, imag} */,
  {32'hbec18ef3, 32'h00000000} /* (14, 27, 13) {real, imag} */,
  {32'hbf09ecd6, 32'h00000000} /* (14, 27, 12) {real, imag} */,
  {32'hbfd61788, 32'h00000000} /* (14, 27, 11) {real, imag} */,
  {32'h3b14881b, 32'h00000000} /* (14, 27, 10) {real, imag} */,
  {32'h3f897d52, 32'h00000000} /* (14, 27, 9) {real, imag} */,
  {32'h3f8eff81, 32'h00000000} /* (14, 27, 8) {real, imag} */,
  {32'h3f7f94bc, 32'h00000000} /* (14, 27, 7) {real, imag} */,
  {32'h3fb3588c, 32'h00000000} /* (14, 27, 6) {real, imag} */,
  {32'h3f88e295, 32'h00000000} /* (14, 27, 5) {real, imag} */,
  {32'h3ee6e94d, 32'h00000000} /* (14, 27, 4) {real, imag} */,
  {32'h3f04c595, 32'h00000000} /* (14, 27, 3) {real, imag} */,
  {32'h3f39c48b, 32'h00000000} /* (14, 27, 2) {real, imag} */,
  {32'h3eb38333, 32'h00000000} /* (14, 27, 1) {real, imag} */,
  {32'h3e3ee69e, 32'h00000000} /* (14, 27, 0) {real, imag} */,
  {32'hbca23250, 32'h00000000} /* (14, 26, 31) {real, imag} */,
  {32'h3f0f0ab0, 32'h00000000} /* (14, 26, 30) {real, imag} */,
  {32'h3f84c86c, 32'h00000000} /* (14, 26, 29) {real, imag} */,
  {32'h3fa506bc, 32'h00000000} /* (14, 26, 28) {real, imag} */,
  {32'h3f4d2eff, 32'h00000000} /* (14, 26, 27) {real, imag} */,
  {32'h3f2fba20, 32'h00000000} /* (14, 26, 26) {real, imag} */,
  {32'h3f9a1096, 32'h00000000} /* (14, 26, 25) {real, imag} */,
  {32'h3f2ac2dd, 32'h00000000} /* (14, 26, 24) {real, imag} */,
  {32'h3ec9b15e, 32'h00000000} /* (14, 26, 23) {real, imag} */,
  {32'h3f597e66, 32'h00000000} /* (14, 26, 22) {real, imag} */,
  {32'h3f24d6ee, 32'h00000000} /* (14, 26, 21) {real, imag} */,
  {32'hbf0907d2, 32'h00000000} /* (14, 26, 20) {real, imag} */,
  {32'hbf308fd2, 32'h00000000} /* (14, 26, 19) {real, imag} */,
  {32'hbf516532, 32'h00000000} /* (14, 26, 18) {real, imag} */,
  {32'hbf55eb3d, 32'h00000000} /* (14, 26, 17) {real, imag} */,
  {32'hbfa8ad2d, 32'h00000000} /* (14, 26, 16) {real, imag} */,
  {32'hbf149306, 32'h00000000} /* (14, 26, 15) {real, imag} */,
  {32'hbf2bc737, 32'h00000000} /* (14, 26, 14) {real, imag} */,
  {32'hbf6451b1, 32'h00000000} /* (14, 26, 13) {real, imag} */,
  {32'hbf6fc0d0, 32'h00000000} /* (14, 26, 12) {real, imag} */,
  {32'hbf7d1d99, 32'h00000000} /* (14, 26, 11) {real, imag} */,
  {32'h3df54849, 32'h00000000} /* (14, 26, 10) {real, imag} */,
  {32'h3ec123d5, 32'h00000000} /* (14, 26, 9) {real, imag} */,
  {32'h3f69ed1f, 32'h00000000} /* (14, 26, 8) {real, imag} */,
  {32'h3fd1c469, 32'h00000000} /* (14, 26, 7) {real, imag} */,
  {32'h3fd83582, 32'h00000000} /* (14, 26, 6) {real, imag} */,
  {32'h3f8ad1b6, 32'h00000000} /* (14, 26, 5) {real, imag} */,
  {32'h3f2f7131, 32'h00000000} /* (14, 26, 4) {real, imag} */,
  {32'h3f861413, 32'h00000000} /* (14, 26, 3) {real, imag} */,
  {32'h3f927e30, 32'h00000000} /* (14, 26, 2) {real, imag} */,
  {32'h3f2fcb0c, 32'h00000000} /* (14, 26, 1) {real, imag} */,
  {32'h3e87549e, 32'h00000000} /* (14, 26, 0) {real, imag} */,
  {32'h3ecc4a76, 32'h00000000} /* (14, 25, 31) {real, imag} */,
  {32'h3f3cc0db, 32'h00000000} /* (14, 25, 30) {real, imag} */,
  {32'h3f6600ad, 32'h00000000} /* (14, 25, 29) {real, imag} */,
  {32'h3fa5c8c2, 32'h00000000} /* (14, 25, 28) {real, imag} */,
  {32'h3f8a1124, 32'h00000000} /* (14, 25, 27) {real, imag} */,
  {32'h3f20c84f, 32'h00000000} /* (14, 25, 26) {real, imag} */,
  {32'h3f94dcde, 32'h00000000} /* (14, 25, 25) {real, imag} */,
  {32'h3f9bb341, 32'h00000000} /* (14, 25, 24) {real, imag} */,
  {32'h3f6db981, 32'h00000000} /* (14, 25, 23) {real, imag} */,
  {32'h3f9bd63e, 32'h00000000} /* (14, 25, 22) {real, imag} */,
  {32'h3f46ad96, 32'h00000000} /* (14, 25, 21) {real, imag} */,
  {32'hbf2ccc5f, 32'h00000000} /* (14, 25, 20) {real, imag} */,
  {32'hbfa31ec1, 32'h00000000} /* (14, 25, 19) {real, imag} */,
  {32'hbf853cff, 32'h00000000} /* (14, 25, 18) {real, imag} */,
  {32'hbf8cec94, 32'h00000000} /* (14, 25, 17) {real, imag} */,
  {32'hbfc0960c, 32'h00000000} /* (14, 25, 16) {real, imag} */,
  {32'hbf64b682, 32'h00000000} /* (14, 25, 15) {real, imag} */,
  {32'hbf75a9c5, 32'h00000000} /* (14, 25, 14) {real, imag} */,
  {32'hbfda500e, 32'h00000000} /* (14, 25, 13) {real, imag} */,
  {32'hbfb4d0d8, 32'h00000000} /* (14, 25, 12) {real, imag} */,
  {32'hbeae98a8, 32'h00000000} /* (14, 25, 11) {real, imag} */,
  {32'h3f052e3d, 32'h00000000} /* (14, 25, 10) {real, imag} */,
  {32'h3f5e15f2, 32'h00000000} /* (14, 25, 9) {real, imag} */,
  {32'h3f6b3d75, 32'h00000000} /* (14, 25, 8) {real, imag} */,
  {32'h3f7d2c56, 32'h00000000} /* (14, 25, 7) {real, imag} */,
  {32'h3f87febe, 32'h00000000} /* (14, 25, 6) {real, imag} */,
  {32'h3f9b67ea, 32'h00000000} /* (14, 25, 5) {real, imag} */,
  {32'h3f71c275, 32'h00000000} /* (14, 25, 4) {real, imag} */,
  {32'h3f906d68, 32'h00000000} /* (14, 25, 3) {real, imag} */,
  {32'h3f781c73, 32'h00000000} /* (14, 25, 2) {real, imag} */,
  {32'h3fa1d32c, 32'h00000000} /* (14, 25, 1) {real, imag} */,
  {32'h3eed4eef, 32'h00000000} /* (14, 25, 0) {real, imag} */,
  {32'h3f54dd81, 32'h00000000} /* (14, 24, 31) {real, imag} */,
  {32'h3f2d635e, 32'h00000000} /* (14, 24, 30) {real, imag} */,
  {32'h3f6514dc, 32'h00000000} /* (14, 24, 29) {real, imag} */,
  {32'h3fb49727, 32'h00000000} /* (14, 24, 28) {real, imag} */,
  {32'h3f4556e0, 32'h00000000} /* (14, 24, 27) {real, imag} */,
  {32'h3e5fd9d6, 32'h00000000} /* (14, 24, 26) {real, imag} */,
  {32'h3f000f31, 32'h00000000} /* (14, 24, 25) {real, imag} */,
  {32'h3fa996a0, 32'h00000000} /* (14, 24, 24) {real, imag} */,
  {32'h3fa2446f, 32'h00000000} /* (14, 24, 23) {real, imag} */,
  {32'h3fc20292, 32'h00000000} /* (14, 24, 22) {real, imag} */,
  {32'h3f22d008, 32'h00000000} /* (14, 24, 21) {real, imag} */,
  {32'hbeea1220, 32'h00000000} /* (14, 24, 20) {real, imag} */,
  {32'hbf51a2a5, 32'h00000000} /* (14, 24, 19) {real, imag} */,
  {32'hbf484568, 32'h00000000} /* (14, 24, 18) {real, imag} */,
  {32'hbf9bbb2a, 32'h00000000} /* (14, 24, 17) {real, imag} */,
  {32'hbfcdf799, 32'h00000000} /* (14, 24, 16) {real, imag} */,
  {32'hbf8c7a84, 32'h00000000} /* (14, 24, 15) {real, imag} */,
  {32'hbf9623a8, 32'h00000000} /* (14, 24, 14) {real, imag} */,
  {32'hbfe56312, 32'h00000000} /* (14, 24, 13) {real, imag} */,
  {32'hbfce30ad, 32'h00000000} /* (14, 24, 12) {real, imag} */,
  {32'hbf9af0a1, 32'h00000000} /* (14, 24, 11) {real, imag} */,
  {32'hbc9aaa11, 32'h00000000} /* (14, 24, 10) {real, imag} */,
  {32'h3fa637a3, 32'h00000000} /* (14, 24, 9) {real, imag} */,
  {32'h3fc7e449, 32'h00000000} /* (14, 24, 8) {real, imag} */,
  {32'h3f86466b, 32'h00000000} /* (14, 24, 7) {real, imag} */,
  {32'h3f2db3ce, 32'h00000000} /* (14, 24, 6) {real, imag} */,
  {32'h3f6ac94b, 32'h00000000} /* (14, 24, 5) {real, imag} */,
  {32'h3f8e72ec, 32'h00000000} /* (14, 24, 4) {real, imag} */,
  {32'h3f9f2035, 32'h00000000} /* (14, 24, 3) {real, imag} */,
  {32'h3f275be0, 32'h00000000} /* (14, 24, 2) {real, imag} */,
  {32'h3f7c087a, 32'h00000000} /* (14, 24, 1) {real, imag} */,
  {32'h3ef04ed8, 32'h00000000} /* (14, 24, 0) {real, imag} */,
  {32'h3f129f38, 32'h00000000} /* (14, 23, 31) {real, imag} */,
  {32'h3f67fec3, 32'h00000000} /* (14, 23, 30) {real, imag} */,
  {32'h3f7ecec7, 32'h00000000} /* (14, 23, 29) {real, imag} */,
  {32'h3f8f2906, 32'h00000000} /* (14, 23, 28) {real, imag} */,
  {32'h3f0a99f0, 32'h00000000} /* (14, 23, 27) {real, imag} */,
  {32'h3f064649, 32'h00000000} /* (14, 23, 26) {real, imag} */,
  {32'h3ee2e0cc, 32'h00000000} /* (14, 23, 25) {real, imag} */,
  {32'h3f53568c, 32'h00000000} /* (14, 23, 24) {real, imag} */,
  {32'h3f9584c6, 32'h00000000} /* (14, 23, 23) {real, imag} */,
  {32'h3f9b3b5e, 32'h00000000} /* (14, 23, 22) {real, imag} */,
  {32'h3ea78a48, 32'h00000000} /* (14, 23, 21) {real, imag} */,
  {32'hbf48ba18, 32'h00000000} /* (14, 23, 20) {real, imag} */,
  {32'hbf20c399, 32'h00000000} /* (14, 23, 19) {real, imag} */,
  {32'hbf5fbf08, 32'h00000000} /* (14, 23, 18) {real, imag} */,
  {32'hbfabcd7b, 32'h00000000} /* (14, 23, 17) {real, imag} */,
  {32'hbfbdc07e, 32'h00000000} /* (14, 23, 16) {real, imag} */,
  {32'hbf83a1f1, 32'h00000000} /* (14, 23, 15) {real, imag} */,
  {32'hbf8e2d2b, 32'h00000000} /* (14, 23, 14) {real, imag} */,
  {32'hbfbcc74a, 32'h00000000} /* (14, 23, 13) {real, imag} */,
  {32'hbfa05505, 32'h00000000} /* (14, 23, 12) {real, imag} */,
  {32'hbf4104e9, 32'h00000000} /* (14, 23, 11) {real, imag} */,
  {32'h3dea236f, 32'h00000000} /* (14, 23, 10) {real, imag} */,
  {32'h3f8e0a4f, 32'h00000000} /* (14, 23, 9) {real, imag} */,
  {32'h3fb781d5, 32'h00000000} /* (14, 23, 8) {real, imag} */,
  {32'h3f43e946, 32'h00000000} /* (14, 23, 7) {real, imag} */,
  {32'h3f4a72b5, 32'h00000000} /* (14, 23, 6) {real, imag} */,
  {32'h3fb6c5a6, 32'h00000000} /* (14, 23, 5) {real, imag} */,
  {32'h3f4ba5f3, 32'h00000000} /* (14, 23, 4) {real, imag} */,
  {32'h3f219bdc, 32'h00000000} /* (14, 23, 3) {real, imag} */,
  {32'h3f0f64cf, 32'h00000000} /* (14, 23, 2) {real, imag} */,
  {32'h3f38c2b7, 32'h00000000} /* (14, 23, 1) {real, imag} */,
  {32'h3f0c649d, 32'h00000000} /* (14, 23, 0) {real, imag} */,
  {32'h3f4170fa, 32'h00000000} /* (14, 22, 31) {real, imag} */,
  {32'h3fa5a345, 32'h00000000} /* (14, 22, 30) {real, imag} */,
  {32'h3fc3577a, 32'h00000000} /* (14, 22, 29) {real, imag} */,
  {32'h3fa7fa6d, 32'h00000000} /* (14, 22, 28) {real, imag} */,
  {32'h3f613c3d, 32'h00000000} /* (14, 22, 27) {real, imag} */,
  {32'h3f2c0c3c, 32'h00000000} /* (14, 22, 26) {real, imag} */,
  {32'h3f012062, 32'h00000000} /* (14, 22, 25) {real, imag} */,
  {32'h3f5da38b, 32'h00000000} /* (14, 22, 24) {real, imag} */,
  {32'h3fb8a515, 32'h00000000} /* (14, 22, 23) {real, imag} */,
  {32'h3fb13b63, 32'h00000000} /* (14, 22, 22) {real, imag} */,
  {32'h3e7c577c, 32'h00000000} /* (14, 22, 21) {real, imag} */,
  {32'hbf20e488, 32'h00000000} /* (14, 22, 20) {real, imag} */,
  {32'hbed4048c, 32'h00000000} /* (14, 22, 19) {real, imag} */,
  {32'hbf4b20ac, 32'h00000000} /* (14, 22, 18) {real, imag} */,
  {32'hbf6db221, 32'h00000000} /* (14, 22, 17) {real, imag} */,
  {32'hbf5366f1, 32'h00000000} /* (14, 22, 16) {real, imag} */,
  {32'hbf3bc638, 32'h00000000} /* (14, 22, 15) {real, imag} */,
  {32'hbf250aee, 32'h00000000} /* (14, 22, 14) {real, imag} */,
  {32'hbf4498c1, 32'h00000000} /* (14, 22, 13) {real, imag} */,
  {32'hbf59ce72, 32'h00000000} /* (14, 22, 12) {real, imag} */,
  {32'hbf467b25, 32'h00000000} /* (14, 22, 11) {real, imag} */,
  {32'h3e90d71b, 32'h00000000} /* (14, 22, 10) {real, imag} */,
  {32'h3f8479d1, 32'h00000000} /* (14, 22, 9) {real, imag} */,
  {32'h3fec8bb2, 32'h00000000} /* (14, 22, 8) {real, imag} */,
  {32'h3f81fa80, 32'h00000000} /* (14, 22, 7) {real, imag} */,
  {32'h3f61ee95, 32'h00000000} /* (14, 22, 6) {real, imag} */,
  {32'h3fc021c4, 32'h00000000} /* (14, 22, 5) {real, imag} */,
  {32'h3f696b18, 32'h00000000} /* (14, 22, 4) {real, imag} */,
  {32'h3eb250ce, 32'h00000000} /* (14, 22, 3) {real, imag} */,
  {32'h3f836c2b, 32'h00000000} /* (14, 22, 2) {real, imag} */,
  {32'h3f8682dc, 32'h00000000} /* (14, 22, 1) {real, imag} */,
  {32'h3f03e2f8, 32'h00000000} /* (14, 22, 0) {real, imag} */,
  {32'h3ef1d504, 32'h00000000} /* (14, 21, 31) {real, imag} */,
  {32'h3f1c80b4, 32'h00000000} /* (14, 21, 30) {real, imag} */,
  {32'h3ed26bb5, 32'h00000000} /* (14, 21, 29) {real, imag} */,
  {32'h3e1c51e8, 32'h00000000} /* (14, 21, 28) {real, imag} */,
  {32'h3ea0cf93, 32'h00000000} /* (14, 21, 27) {real, imag} */,
  {32'hbe2f8396, 32'h00000000} /* (14, 21, 26) {real, imag} */,
  {32'hbdd12374, 32'h00000000} /* (14, 21, 25) {real, imag} */,
  {32'h3f025246, 32'h00000000} /* (14, 21, 24) {real, imag} */,
  {32'h3f38810b, 32'h00000000} /* (14, 21, 23) {real, imag} */,
  {32'h3f900b16, 32'h00000000} /* (14, 21, 22) {real, imag} */,
  {32'h3ecbd9e8, 32'h00000000} /* (14, 21, 21) {real, imag} */,
  {32'h3e4c7938, 32'h00000000} /* (14, 21, 20) {real, imag} */,
  {32'hbd1eb7f0, 32'h00000000} /* (14, 21, 19) {real, imag} */,
  {32'hbe916fe8, 32'h00000000} /* (14, 21, 18) {real, imag} */,
  {32'hbe1b17ee, 32'h00000000} /* (14, 21, 17) {real, imag} */,
  {32'hbd986932, 32'h00000000} /* (14, 21, 16) {real, imag} */,
  {32'hbd996c91, 32'h00000000} /* (14, 21, 15) {real, imag} */,
  {32'hbe5aa826, 32'h00000000} /* (14, 21, 14) {real, imag} */,
  {32'hbe323520, 32'h00000000} /* (14, 21, 13) {real, imag} */,
  {32'hbda92c7d, 32'h00000000} /* (14, 21, 12) {real, imag} */,
  {32'hbd802eee, 32'h00000000} /* (14, 21, 11) {real, imag} */,
  {32'h3cb472fe, 32'h00000000} /* (14, 21, 10) {real, imag} */,
  {32'h3f96bd66, 32'h00000000} /* (14, 21, 9) {real, imag} */,
  {32'h3fbe5378, 32'h00000000} /* (14, 21, 8) {real, imag} */,
  {32'h3f465379, 32'h00000000} /* (14, 21, 7) {real, imag} */,
  {32'h3eaa1cb4, 32'h00000000} /* (14, 21, 6) {real, imag} */,
  {32'h3eba218a, 32'h00000000} /* (14, 21, 5) {real, imag} */,
  {32'h3f3ca5dc, 32'h00000000} /* (14, 21, 4) {real, imag} */,
  {32'h3f27ae79, 32'h00000000} /* (14, 21, 3) {real, imag} */,
  {32'h3e94902b, 32'h00000000} /* (14, 21, 2) {real, imag} */,
  {32'h3f024ad8, 32'h00000000} /* (14, 21, 1) {real, imag} */,
  {32'h3ec5f176, 32'h00000000} /* (14, 21, 0) {real, imag} */,
  {32'hbe59b1b4, 32'h00000000} /* (14, 20, 31) {real, imag} */,
  {32'hbe9c9ae9, 32'h00000000} /* (14, 20, 30) {real, imag} */,
  {32'hbf8d8a06, 32'h00000000} /* (14, 20, 29) {real, imag} */,
  {32'hbfc9d4ac, 32'h00000000} /* (14, 20, 28) {real, imag} */,
  {32'hbf83b5d5, 32'h00000000} /* (14, 20, 27) {real, imag} */,
  {32'hbf87a789, 32'h00000000} /* (14, 20, 26) {real, imag} */,
  {32'hbf86337b, 32'h00000000} /* (14, 20, 25) {real, imag} */,
  {32'hbef0c890, 32'h00000000} /* (14, 20, 24) {real, imag} */,
  {32'hbef1d844, 32'h00000000} /* (14, 20, 23) {real, imag} */,
  {32'hbf1334e3, 32'h00000000} /* (14, 20, 22) {real, imag} */,
  {32'hbd358b95, 32'h00000000} /* (14, 20, 21) {real, imag} */,
  {32'h3f3538a6, 32'h00000000} /* (14, 20, 20) {real, imag} */,
  {32'h3f0b3bc1, 32'h00000000} /* (14, 20, 19) {real, imag} */,
  {32'h3f34f86a, 32'h00000000} /* (14, 20, 18) {real, imag} */,
  {32'h3f33d665, 32'h00000000} /* (14, 20, 17) {real, imag} */,
  {32'h3f702765, 32'h00000000} /* (14, 20, 16) {real, imag} */,
  {32'h3f4d0239, 32'h00000000} /* (14, 20, 15) {real, imag} */,
  {32'h3f478b6f, 32'h00000000} /* (14, 20, 14) {real, imag} */,
  {32'h3f264934, 32'h00000000} /* (14, 20, 13) {real, imag} */,
  {32'h3f457f59, 32'h00000000} /* (14, 20, 12) {real, imag} */,
  {32'h3f8ac962, 32'h00000000} /* (14, 20, 11) {real, imag} */,
  {32'hbeaf0a02, 32'h00000000} /* (14, 20, 10) {real, imag} */,
  {32'hbd1e7bbf, 32'h00000000} /* (14, 20, 9) {real, imag} */,
  {32'hbea3dbca, 32'h00000000} /* (14, 20, 8) {real, imag} */,
  {32'hbf6b1446, 32'h00000000} /* (14, 20, 7) {real, imag} */,
  {32'hbf3ba599, 32'h00000000} /* (14, 20, 6) {real, imag} */,
  {32'hbf17a376, 32'h00000000} /* (14, 20, 5) {real, imag} */,
  {32'hbeb24f09, 32'h00000000} /* (14, 20, 4) {real, imag} */,
  {32'hbeff4169, 32'h00000000} /* (14, 20, 3) {real, imag} */,
  {32'hbf8a7de0, 32'h00000000} /* (14, 20, 2) {real, imag} */,
  {32'hbf4bbdbf, 32'h00000000} /* (14, 20, 1) {real, imag} */,
  {32'hbf083655, 32'h00000000} /* (14, 20, 0) {real, imag} */,
  {32'hbe844854, 32'h00000000} /* (14, 19, 31) {real, imag} */,
  {32'hbedaa29c, 32'h00000000} /* (14, 19, 30) {real, imag} */,
  {32'hbf3db81e, 32'h00000000} /* (14, 19, 29) {real, imag} */,
  {32'hbf6742a9, 32'h00000000} /* (14, 19, 28) {real, imag} */,
  {32'hbfbec628, 32'h00000000} /* (14, 19, 27) {real, imag} */,
  {32'hbfa07ed0, 32'h00000000} /* (14, 19, 26) {real, imag} */,
  {32'hbf4a0596, 32'h00000000} /* (14, 19, 25) {real, imag} */,
  {32'hbf1c41de, 32'h00000000} /* (14, 19, 24) {real, imag} */,
  {32'hbf47cd49, 32'h00000000} /* (14, 19, 23) {real, imag} */,
  {32'hbf7b29f1, 32'h00000000} /* (14, 19, 22) {real, imag} */,
  {32'hbd0e0dfc, 32'h00000000} /* (14, 19, 21) {real, imag} */,
  {32'h3f569611, 32'h00000000} /* (14, 19, 20) {real, imag} */,
  {32'h3f959b36, 32'h00000000} /* (14, 19, 19) {real, imag} */,
  {32'h3f7c0ddd, 32'h00000000} /* (14, 19, 18) {real, imag} */,
  {32'h3f1506cc, 32'h00000000} /* (14, 19, 17) {real, imag} */,
  {32'h3f5c73fe, 32'h00000000} /* (14, 19, 16) {real, imag} */,
  {32'h3f683ec8, 32'h00000000} /* (14, 19, 15) {real, imag} */,
  {32'h3f6d7d82, 32'h00000000} /* (14, 19, 14) {real, imag} */,
  {32'h3f8ed80b, 32'h00000000} /* (14, 19, 13) {real, imag} */,
  {32'h3faab35a, 32'h00000000} /* (14, 19, 12) {real, imag} */,
  {32'h3f984023, 32'h00000000} /* (14, 19, 11) {real, imag} */,
  {32'hbe3edfba, 32'h00000000} /* (14, 19, 10) {real, imag} */,
  {32'hbee19579, 32'h00000000} /* (14, 19, 9) {real, imag} */,
  {32'hbf114236, 32'h00000000} /* (14, 19, 8) {real, imag} */,
  {32'hbfbcd351, 32'h00000000} /* (14, 19, 7) {real, imag} */,
  {32'hbf7750ff, 32'h00000000} /* (14, 19, 6) {real, imag} */,
  {32'hbefd497a, 32'h00000000} /* (14, 19, 5) {real, imag} */,
  {32'hbf42295b, 32'h00000000} /* (14, 19, 4) {real, imag} */,
  {32'hbf401b50, 32'h00000000} /* (14, 19, 3) {real, imag} */,
  {32'hbf00f8d5, 32'h00000000} /* (14, 19, 2) {real, imag} */,
  {32'hbf1726fe, 32'h00000000} /* (14, 19, 1) {real, imag} */,
  {32'hbefac3ba, 32'h00000000} /* (14, 19, 0) {real, imag} */,
  {32'hbeb364f7, 32'h00000000} /* (14, 18, 31) {real, imag} */,
  {32'hbeec0b66, 32'h00000000} /* (14, 18, 30) {real, imag} */,
  {32'hbe8ff2b0, 32'h00000000} /* (14, 18, 29) {real, imag} */,
  {32'hbe86a9ca, 32'h00000000} /* (14, 18, 28) {real, imag} */,
  {32'hbf4165fc, 32'h00000000} /* (14, 18, 27) {real, imag} */,
  {32'hbf582a17, 32'h00000000} /* (14, 18, 26) {real, imag} */,
  {32'hbf147e6a, 32'h00000000} /* (14, 18, 25) {real, imag} */,
  {32'hbf34e8dd, 32'h00000000} /* (14, 18, 24) {real, imag} */,
  {32'hbf87f61c, 32'h00000000} /* (14, 18, 23) {real, imag} */,
  {32'hbf6f92c8, 32'h00000000} /* (14, 18, 22) {real, imag} */,
  {32'hbe009c56, 32'h00000000} /* (14, 18, 21) {real, imag} */,
  {32'h3f220633, 32'h00000000} /* (14, 18, 20) {real, imag} */,
  {32'h3f894fc5, 32'h00000000} /* (14, 18, 19) {real, imag} */,
  {32'h3f30bb9f, 32'h00000000} /* (14, 18, 18) {real, imag} */,
  {32'h3f0013b7, 32'h00000000} /* (14, 18, 17) {real, imag} */,
  {32'h3f701d8b, 32'h00000000} /* (14, 18, 16) {real, imag} */,
  {32'h3f2d4d92, 32'h00000000} /* (14, 18, 15) {real, imag} */,
  {32'h3f272ac4, 32'h00000000} /* (14, 18, 14) {real, imag} */,
  {32'h3f971c80, 32'h00000000} /* (14, 18, 13) {real, imag} */,
  {32'h3f7c3fdc, 32'h00000000} /* (14, 18, 12) {real, imag} */,
  {32'h3f760b43, 32'h00000000} /* (14, 18, 11) {real, imag} */,
  {32'hbd9a19d6, 32'h00000000} /* (14, 18, 10) {real, imag} */,
  {32'hbec494f9, 32'h00000000} /* (14, 18, 9) {real, imag} */,
  {32'hbf0fa657, 32'h00000000} /* (14, 18, 8) {real, imag} */,
  {32'hbf50506b, 32'h00000000} /* (14, 18, 7) {real, imag} */,
  {32'hbf9d4629, 32'h00000000} /* (14, 18, 6) {real, imag} */,
  {32'hbf8d873c, 32'h00000000} /* (14, 18, 5) {real, imag} */,
  {32'hbf59600b, 32'h00000000} /* (14, 18, 4) {real, imag} */,
  {32'hbf3640f1, 32'h00000000} /* (14, 18, 3) {real, imag} */,
  {32'hbe3a96c7, 32'h00000000} /* (14, 18, 2) {real, imag} */,
  {32'hbf74e675, 32'h00000000} /* (14, 18, 1) {real, imag} */,
  {32'hbf32e12a, 32'h00000000} /* (14, 18, 0) {real, imag} */,
  {32'hbe3fcccc, 32'h00000000} /* (14, 17, 31) {real, imag} */,
  {32'hbf0be0b4, 32'h00000000} /* (14, 17, 30) {real, imag} */,
  {32'hbee05d77, 32'h00000000} /* (14, 17, 29) {real, imag} */,
  {32'hbe949af1, 32'h00000000} /* (14, 17, 28) {real, imag} */,
  {32'hbf82a291, 32'h00000000} /* (14, 17, 27) {real, imag} */,
  {32'hbf5e77a2, 32'h00000000} /* (14, 17, 26) {real, imag} */,
  {32'hbf7cc806, 32'h00000000} /* (14, 17, 25) {real, imag} */,
  {32'hbf7615f6, 32'h00000000} /* (14, 17, 24) {real, imag} */,
  {32'hbfa81d02, 32'h00000000} /* (14, 17, 23) {real, imag} */,
  {32'hbfaa430e, 32'h00000000} /* (14, 17, 22) {real, imag} */,
  {32'hbe8b96b1, 32'h00000000} /* (14, 17, 21) {real, imag} */,
  {32'h3f3e049a, 32'h00000000} /* (14, 17, 20) {real, imag} */,
  {32'h3f994601, 32'h00000000} /* (14, 17, 19) {real, imag} */,
  {32'h3f69af98, 32'h00000000} /* (14, 17, 18) {real, imag} */,
  {32'h3f23ea69, 32'h00000000} /* (14, 17, 17) {real, imag} */,
  {32'h3f3a4ae7, 32'h00000000} /* (14, 17, 16) {real, imag} */,
  {32'h3f091ae2, 32'h00000000} /* (14, 17, 15) {real, imag} */,
  {32'h3ee42726, 32'h00000000} /* (14, 17, 14) {real, imag} */,
  {32'h3f2a671a, 32'h00000000} /* (14, 17, 13) {real, imag} */,
  {32'h3f258740, 32'h00000000} /* (14, 17, 12) {real, imag} */,
  {32'h3e38ce66, 32'h00000000} /* (14, 17, 11) {real, imag} */,
  {32'hbf64c4e3, 32'h00000000} /* (14, 17, 10) {real, imag} */,
  {32'hbf427a74, 32'h00000000} /* (14, 17, 9) {real, imag} */,
  {32'hbf2eeb0d, 32'h00000000} /* (14, 17, 8) {real, imag} */,
  {32'hbf57022e, 32'h00000000} /* (14, 17, 7) {real, imag} */,
  {32'hbfd51500, 32'h00000000} /* (14, 17, 6) {real, imag} */,
  {32'hbfeab188, 32'h00000000} /* (14, 17, 5) {real, imag} */,
  {32'hbf9d73df, 32'h00000000} /* (14, 17, 4) {real, imag} */,
  {32'hbf00c7c0, 32'h00000000} /* (14, 17, 3) {real, imag} */,
  {32'hbefc2260, 32'h00000000} /* (14, 17, 2) {real, imag} */,
  {32'hbf8db412, 32'h00000000} /* (14, 17, 1) {real, imag} */,
  {32'hbf22da75, 32'h00000000} /* (14, 17, 0) {real, imag} */,
  {32'hbe558c2f, 32'h00000000} /* (14, 16, 31) {real, imag} */,
  {32'hbf3b0d45, 32'h00000000} /* (14, 16, 30) {real, imag} */,
  {32'hbf300d36, 32'h00000000} /* (14, 16, 29) {real, imag} */,
  {32'hbea0fabe, 32'h00000000} /* (14, 16, 28) {real, imag} */,
  {32'hbf890c7f, 32'h00000000} /* (14, 16, 27) {real, imag} */,
  {32'hbf54e1de, 32'h00000000} /* (14, 16, 26) {real, imag} */,
  {32'hbf431598, 32'h00000000} /* (14, 16, 25) {real, imag} */,
  {32'hbfa507ab, 32'h00000000} /* (14, 16, 24) {real, imag} */,
  {32'hbff0a127, 32'h00000000} /* (14, 16, 23) {real, imag} */,
  {32'hbfe71933, 32'h00000000} /* (14, 16, 22) {real, imag} */,
  {32'hbe8d8056, 32'h00000000} /* (14, 16, 21) {real, imag} */,
  {32'h3f53e4af, 32'h00000000} /* (14, 16, 20) {real, imag} */,
  {32'h3f904c40, 32'h00000000} /* (14, 16, 19) {real, imag} */,
  {32'h3fa331cc, 32'h00000000} /* (14, 16, 18) {real, imag} */,
  {32'h3fb0d120, 32'h00000000} /* (14, 16, 17) {real, imag} */,
  {32'h3f94d07e, 32'h00000000} /* (14, 16, 16) {real, imag} */,
  {32'h3f56f8ef, 32'h00000000} /* (14, 16, 15) {real, imag} */,
  {32'h3f4f5eb0, 32'h00000000} /* (14, 16, 14) {real, imag} */,
  {32'h3f35aa59, 32'h00000000} /* (14, 16, 13) {real, imag} */,
  {32'h3f740b26, 32'h00000000} /* (14, 16, 12) {real, imag} */,
  {32'h3f7126e3, 32'h00000000} /* (14, 16, 11) {real, imag} */,
  {32'hbddf3b21, 32'h00000000} /* (14, 16, 10) {real, imag} */,
  {32'hbea54355, 32'h00000000} /* (14, 16, 9) {real, imag} */,
  {32'hbf3a761b, 32'h00000000} /* (14, 16, 8) {real, imag} */,
  {32'hbfa18769, 32'h00000000} /* (14, 16, 7) {real, imag} */,
  {32'hbf92249d, 32'h00000000} /* (14, 16, 6) {real, imag} */,
  {32'hbfa1f9ed, 32'h00000000} /* (14, 16, 5) {real, imag} */,
  {32'hbf796243, 32'h00000000} /* (14, 16, 4) {real, imag} */,
  {32'hbf1775d0, 32'h00000000} /* (14, 16, 3) {real, imag} */,
  {32'hbf6cd4c6, 32'h00000000} /* (14, 16, 2) {real, imag} */,
  {32'hbf34a4fe, 32'h00000000} /* (14, 16, 1) {real, imag} */,
  {32'hbe805261, 32'h00000000} /* (14, 16, 0) {real, imag} */,
  {32'hbed1fc92, 32'h00000000} /* (14, 15, 31) {real, imag} */,
  {32'hbf8ecef9, 32'h00000000} /* (14, 15, 30) {real, imag} */,
  {32'hbf9fe784, 32'h00000000} /* (14, 15, 29) {real, imag} */,
  {32'hbf74a984, 32'h00000000} /* (14, 15, 28) {real, imag} */,
  {32'hbf99dd63, 32'h00000000} /* (14, 15, 27) {real, imag} */,
  {32'hbf94d464, 32'h00000000} /* (14, 15, 26) {real, imag} */,
  {32'hbf3f45ba, 32'h00000000} /* (14, 15, 25) {real, imag} */,
  {32'hbf4da318, 32'h00000000} /* (14, 15, 24) {real, imag} */,
  {32'hc0147253, 32'h00000000} /* (14, 15, 23) {real, imag} */,
  {32'hbfefd51d, 32'h00000000} /* (14, 15, 22) {real, imag} */,
  {32'hbe4379a4, 32'h00000000} /* (14, 15, 21) {real, imag} */,
  {32'h3f1f4ab7, 32'h00000000} /* (14, 15, 20) {real, imag} */,
  {32'h3f80fb24, 32'h00000000} /* (14, 15, 19) {real, imag} */,
  {32'h3f6a7f6a, 32'h00000000} /* (14, 15, 18) {real, imag} */,
  {32'h3f822719, 32'h00000000} /* (14, 15, 17) {real, imag} */,
  {32'h3fbe84d1, 32'h00000000} /* (14, 15, 16) {real, imag} */,
  {32'h3f9c811e, 32'h00000000} /* (14, 15, 15) {real, imag} */,
  {32'h3f7b9ff9, 32'h00000000} /* (14, 15, 14) {real, imag} */,
  {32'h3f24d6f3, 32'h00000000} /* (14, 15, 13) {real, imag} */,
  {32'h3f478e53, 32'h00000000} /* (14, 15, 12) {real, imag} */,
  {32'h3f94b5a7, 32'h00000000} /* (14, 15, 11) {real, imag} */,
  {32'h3e1a35bc, 32'h00000000} /* (14, 15, 10) {real, imag} */,
  {32'hbe8d4ed2, 32'h00000000} /* (14, 15, 9) {real, imag} */,
  {32'hbf34f46e, 32'h00000000} /* (14, 15, 8) {real, imag} */,
  {32'hbfa4785b, 32'h00000000} /* (14, 15, 7) {real, imag} */,
  {32'hbfcd59bb, 32'h00000000} /* (14, 15, 6) {real, imag} */,
  {32'hbfa1aa7a, 32'h00000000} /* (14, 15, 5) {real, imag} */,
  {32'hbf0813f7, 32'h00000000} /* (14, 15, 4) {real, imag} */,
  {32'hbf322d4c, 32'h00000000} /* (14, 15, 3) {real, imag} */,
  {32'hbfa689e5, 32'h00000000} /* (14, 15, 2) {real, imag} */,
  {32'hbf828c1b, 32'h00000000} /* (14, 15, 1) {real, imag} */,
  {32'hbf21501b, 32'h00000000} /* (14, 15, 0) {real, imag} */,
  {32'hbef84157, 32'h00000000} /* (14, 14, 31) {real, imag} */,
  {32'hbf8fae87, 32'h00000000} /* (14, 14, 30) {real, imag} */,
  {32'hbfc6c79d, 32'h00000000} /* (14, 14, 29) {real, imag} */,
  {32'hbfb8f3b8, 32'h00000000} /* (14, 14, 28) {real, imag} */,
  {32'hbfb1a1e1, 32'h00000000} /* (14, 14, 27) {real, imag} */,
  {32'hbf1a33e9, 32'h00000000} /* (14, 14, 26) {real, imag} */,
  {32'hbec981db, 32'h00000000} /* (14, 14, 25) {real, imag} */,
  {32'hbef3393f, 32'h00000000} /* (14, 14, 24) {real, imag} */,
  {32'hbf988f84, 32'h00000000} /* (14, 14, 23) {real, imag} */,
  {32'hbf816d2b, 32'h00000000} /* (14, 14, 22) {real, imag} */,
  {32'hbe5671fe, 32'h00000000} /* (14, 14, 21) {real, imag} */,
  {32'h3f311d6f, 32'h00000000} /* (14, 14, 20) {real, imag} */,
  {32'h3f33ec0a, 32'h00000000} /* (14, 14, 19) {real, imag} */,
  {32'h3f34359c, 32'h00000000} /* (14, 14, 18) {real, imag} */,
  {32'h3f8736d5, 32'h00000000} /* (14, 14, 17) {real, imag} */,
  {32'h3fac0b3c, 32'h00000000} /* (14, 14, 16) {real, imag} */,
  {32'h3f939482, 32'h00000000} /* (14, 14, 15) {real, imag} */,
  {32'h3f4959e0, 32'h00000000} /* (14, 14, 14) {real, imag} */,
  {32'h3f6e5bf6, 32'h00000000} /* (14, 14, 13) {real, imag} */,
  {32'h3f4ac8ba, 32'h00000000} /* (14, 14, 12) {real, imag} */,
  {32'h3f7c51fe, 32'h00000000} /* (14, 14, 11) {real, imag} */,
  {32'hbd93e1ce, 32'h00000000} /* (14, 14, 10) {real, imag} */,
  {32'hbed12b55, 32'h00000000} /* (14, 14, 9) {real, imag} */,
  {32'hbeabbc1c, 32'h00000000} /* (14, 14, 8) {real, imag} */,
  {32'hbf6bcbd6, 32'h00000000} /* (14, 14, 7) {real, imag} */,
  {32'hbfabbb60, 32'h00000000} /* (14, 14, 6) {real, imag} */,
  {32'hbf692679, 32'h00000000} /* (14, 14, 5) {real, imag} */,
  {32'hbf732660, 32'h00000000} /* (14, 14, 4) {real, imag} */,
  {32'hbf9618ae, 32'h00000000} /* (14, 14, 3) {real, imag} */,
  {32'hbf96cade, 32'h00000000} /* (14, 14, 2) {real, imag} */,
  {32'hbf9183a0, 32'h00000000} /* (14, 14, 1) {real, imag} */,
  {32'hbf258dd0, 32'h00000000} /* (14, 14, 0) {real, imag} */,
  {32'hbed0c8bc, 32'h00000000} /* (14, 13, 31) {real, imag} */,
  {32'hbf9deb8e, 32'h00000000} /* (14, 13, 30) {real, imag} */,
  {32'hbf7e0f59, 32'h00000000} /* (14, 13, 29) {real, imag} */,
  {32'hbf899854, 32'h00000000} /* (14, 13, 28) {real, imag} */,
  {32'hbf97d1ac, 32'h00000000} /* (14, 13, 27) {real, imag} */,
  {32'hbe91c56c, 32'h00000000} /* (14, 13, 26) {real, imag} */,
  {32'hbe8b4e74, 32'h00000000} /* (14, 13, 25) {real, imag} */,
  {32'hbf384ad4, 32'h00000000} /* (14, 13, 24) {real, imag} */,
  {32'hbee9b586, 32'h00000000} /* (14, 13, 23) {real, imag} */,
  {32'hbf0585ce, 32'h00000000} /* (14, 13, 22) {real, imag} */,
  {32'hbeb80812, 32'h00000000} /* (14, 13, 21) {real, imag} */,
  {32'h3f551cfd, 32'h00000000} /* (14, 13, 20) {real, imag} */,
  {32'h3f809441, 32'h00000000} /* (14, 13, 19) {real, imag} */,
  {32'h3f6c5671, 32'h00000000} /* (14, 13, 18) {real, imag} */,
  {32'h3f6bfcec, 32'h00000000} /* (14, 13, 17) {real, imag} */,
  {32'h3f3aed63, 32'h00000000} /* (14, 13, 16) {real, imag} */,
  {32'h3f4b70d3, 32'h00000000} /* (14, 13, 15) {real, imag} */,
  {32'h3f22f06b, 32'h00000000} /* (14, 13, 14) {real, imag} */,
  {32'h3f50696e, 32'h00000000} /* (14, 13, 13) {real, imag} */,
  {32'h3f808064, 32'h00000000} /* (14, 13, 12) {real, imag} */,
  {32'h3f59c22b, 32'h00000000} /* (14, 13, 11) {real, imag} */,
  {32'hbce23520, 32'h00000000} /* (14, 13, 10) {real, imag} */,
  {32'hbec95182, 32'h00000000} /* (14, 13, 9) {real, imag} */,
  {32'hbf13c611, 32'h00000000} /* (14, 13, 8) {real, imag} */,
  {32'hbfb27cdf, 32'h00000000} /* (14, 13, 7) {real, imag} */,
  {32'hbf9f7577, 32'h00000000} /* (14, 13, 6) {real, imag} */,
  {32'hbefecac9, 32'h00000000} /* (14, 13, 5) {real, imag} */,
  {32'hbf3fa929, 32'h00000000} /* (14, 13, 4) {real, imag} */,
  {32'hbf952b16, 32'h00000000} /* (14, 13, 3) {real, imag} */,
  {32'hbf5e7daf, 32'h00000000} /* (14, 13, 2) {real, imag} */,
  {32'hbf69bb0b, 32'h00000000} /* (14, 13, 1) {real, imag} */,
  {32'hbf0063af, 32'h00000000} /* (14, 13, 0) {real, imag} */,
  {32'hbee76068, 32'h00000000} /* (14, 12, 31) {real, imag} */,
  {32'hbfb07cca, 32'h00000000} /* (14, 12, 30) {real, imag} */,
  {32'hbfc5f83a, 32'h00000000} /* (14, 12, 29) {real, imag} */,
  {32'hbf8d9666, 32'h00000000} /* (14, 12, 28) {real, imag} */,
  {32'hbf31365f, 32'h00000000} /* (14, 12, 27) {real, imag} */,
  {32'hbf191851, 32'h00000000} /* (14, 12, 26) {real, imag} */,
  {32'hbf069276, 32'h00000000} /* (14, 12, 25) {real, imag} */,
  {32'hbf78f6e6, 32'h00000000} /* (14, 12, 24) {real, imag} */,
  {32'hbf20a974, 32'h00000000} /* (14, 12, 23) {real, imag} */,
  {32'hbf50d118, 32'h00000000} /* (14, 12, 22) {real, imag} */,
  {32'hbe96acb3, 32'h00000000} /* (14, 12, 21) {real, imag} */,
  {32'h3f5ee4d4, 32'h00000000} /* (14, 12, 20) {real, imag} */,
  {32'h3fc3deff, 32'h00000000} /* (14, 12, 19) {real, imag} */,
  {32'h3fadc9c9, 32'h00000000} /* (14, 12, 18) {real, imag} */,
  {32'h3fa73919, 32'h00000000} /* (14, 12, 17) {real, imag} */,
  {32'h3f35b0d9, 32'h00000000} /* (14, 12, 16) {real, imag} */,
  {32'h3efa2def, 32'h00000000} /* (14, 12, 15) {real, imag} */,
  {32'h3ed3d968, 32'h00000000} /* (14, 12, 14) {real, imag} */,
  {32'h3f831d8e, 32'h00000000} /* (14, 12, 13) {real, imag} */,
  {32'h3fcb3d63, 32'h00000000} /* (14, 12, 12) {real, imag} */,
  {32'h3f8dae93, 32'h00000000} /* (14, 12, 11) {real, imag} */,
  {32'hbddc4fc9, 32'h00000000} /* (14, 12, 10) {real, imag} */,
  {32'hbee6c702, 32'h00000000} /* (14, 12, 9) {real, imag} */,
  {32'hbf2a1cf9, 32'h00000000} /* (14, 12, 8) {real, imag} */,
  {32'hbf725fa4, 32'h00000000} /* (14, 12, 7) {real, imag} */,
  {32'hbf235687, 32'h00000000} /* (14, 12, 6) {real, imag} */,
  {32'hbe3c777c, 32'h00000000} /* (14, 12, 5) {real, imag} */,
  {32'hbf0722fa, 32'h00000000} /* (14, 12, 4) {real, imag} */,
  {32'hbf7723e0, 32'h00000000} /* (14, 12, 3) {real, imag} */,
  {32'hbf767a3d, 32'h00000000} /* (14, 12, 2) {real, imag} */,
  {32'hbf727cb2, 32'h00000000} /* (14, 12, 1) {real, imag} */,
  {32'hbe96e27c, 32'h00000000} /* (14, 12, 0) {real, imag} */,
  {32'h3e19b932, 32'h00000000} /* (14, 11, 31) {real, imag} */,
  {32'hbe5fa60b, 32'h00000000} /* (14, 11, 30) {real, imag} */,
  {32'hbfa1d5cb, 32'h00000000} /* (14, 11, 29) {real, imag} */,
  {32'hbf941bd1, 32'h00000000} /* (14, 11, 28) {real, imag} */,
  {32'hbf1b56be, 32'h00000000} /* (14, 11, 27) {real, imag} */,
  {32'hbf91e36f, 32'h00000000} /* (14, 11, 26) {real, imag} */,
  {32'hbf1a9a64, 32'h00000000} /* (14, 11, 25) {real, imag} */,
  {32'hbf27ee5f, 32'h00000000} /* (14, 11, 24) {real, imag} */,
  {32'hbf7cea1c, 32'h00000000} /* (14, 11, 23) {real, imag} */,
  {32'hbedeb453, 32'h00000000} /* (14, 11, 22) {real, imag} */,
  {32'hbe74f8f1, 32'h00000000} /* (14, 11, 21) {real, imag} */,
  {32'h3eaea06b, 32'h00000000} /* (14, 11, 20) {real, imag} */,
  {32'h3f23ffda, 32'h00000000} /* (14, 11, 19) {real, imag} */,
  {32'h3f1c2f81, 32'h00000000} /* (14, 11, 18) {real, imag} */,
  {32'h3fb116df, 32'h00000000} /* (14, 11, 17) {real, imag} */,
  {32'h3f792848, 32'h00000000} /* (14, 11, 16) {real, imag} */,
  {32'h3ea88664, 32'h00000000} /* (14, 11, 15) {real, imag} */,
  {32'h3ead3e32, 32'h00000000} /* (14, 11, 14) {real, imag} */,
  {32'h3f38fa40, 32'h00000000} /* (14, 11, 13) {real, imag} */,
  {32'h3f899f3e, 32'h00000000} /* (14, 11, 12) {real, imag} */,
  {32'h3f557ed3, 32'h00000000} /* (14, 11, 11) {real, imag} */,
  {32'hbed0f1fc, 32'h00000000} /* (14, 11, 10) {real, imag} */,
  {32'hbf2afe95, 32'h00000000} /* (14, 11, 9) {real, imag} */,
  {32'hbf28f18a, 32'h00000000} /* (14, 11, 8) {real, imag} */,
  {32'hbf3d9ace, 32'h00000000} /* (14, 11, 7) {real, imag} */,
  {32'hbf2120c2, 32'h00000000} /* (14, 11, 6) {real, imag} */,
  {32'hbe3aeac1, 32'h00000000} /* (14, 11, 5) {real, imag} */,
  {32'hbed39c78, 32'h00000000} /* (14, 11, 4) {real, imag} */,
  {32'hbe7a55e6, 32'h00000000} /* (14, 11, 3) {real, imag} */,
  {32'hbdc5c2f4, 32'h00000000} /* (14, 11, 2) {real, imag} */,
  {32'hbed382bd, 32'h00000000} /* (14, 11, 1) {real, imag} */,
  {32'hbe2d47b3, 32'h00000000} /* (14, 11, 0) {real, imag} */,
  {32'h3f43c1cd, 32'h00000000} /* (14, 10, 31) {real, imag} */,
  {32'h3f7b0f39, 32'h00000000} /* (14, 10, 30) {real, imag} */,
  {32'h3fcf2188, 32'h00000000} /* (14, 10, 29) {real, imag} */,
  {32'h3f59fb66, 32'h00000000} /* (14, 10, 28) {real, imag} */,
  {32'h3ec64e87, 32'h00000000} /* (14, 10, 27) {real, imag} */,
  {32'h3e8bc728, 32'h00000000} /* (14, 10, 26) {real, imag} */,
  {32'h3dd67023, 32'h00000000} /* (14, 10, 25) {real, imag} */,
  {32'h3ea15c50, 32'h00000000} /* (14, 10, 24) {real, imag} */,
  {32'hbd283c74, 32'h00000000} /* (14, 10, 23) {real, imag} */,
  {32'h3f34b665, 32'h00000000} /* (14, 10, 22) {real, imag} */,
  {32'h3de8fde5, 32'h00000000} /* (14, 10, 21) {real, imag} */,
  {32'hbef1ac44, 32'h00000000} /* (14, 10, 20) {real, imag} */,
  {32'hbf1bc2c2, 32'h00000000} /* (14, 10, 19) {real, imag} */,
  {32'hbf78dec5, 32'h00000000} /* (14, 10, 18) {real, imag} */,
  {32'hbe882a69, 32'h00000000} /* (14, 10, 17) {real, imag} */,
  {32'hbe3e0d3f, 32'h00000000} /* (14, 10, 16) {real, imag} */,
  {32'hbf03c033, 32'h00000000} /* (14, 10, 15) {real, imag} */,
  {32'hbef26f9c, 32'h00000000} /* (14, 10, 14) {real, imag} */,
  {32'hbf119253, 32'h00000000} /* (14, 10, 13) {real, imag} */,
  {32'hbeb0c389, 32'h00000000} /* (14, 10, 12) {real, imag} */,
  {32'hbe9e0e5e, 32'h00000000} /* (14, 10, 11) {real, imag} */,
  {32'hbe503681, 32'h00000000} /* (14, 10, 10) {real, imag} */,
  {32'hbdcc1cc1, 32'h00000000} /* (14, 10, 9) {real, imag} */,
  {32'h3e99d2c9, 32'h00000000} /* (14, 10, 8) {real, imag} */,
  {32'h3d159014, 32'h00000000} /* (14, 10, 7) {real, imag} */,
  {32'hbde2f0e4, 32'h00000000} /* (14, 10, 6) {real, imag} */,
  {32'h3eda144e, 32'h00000000} /* (14, 10, 5) {real, imag} */,
  {32'h3f19d648, 32'h00000000} /* (14, 10, 4) {real, imag} */,
  {32'h3f8e3e04, 32'h00000000} /* (14, 10, 3) {real, imag} */,
  {32'h3fb97e40, 32'h00000000} /* (14, 10, 2) {real, imag} */,
  {32'h3f8f2625, 32'h00000000} /* (14, 10, 1) {real, imag} */,
  {32'h3f0e39e9, 32'h00000000} /* (14, 10, 0) {real, imag} */,
  {32'h3e796ac9, 32'h00000000} /* (14, 9, 31) {real, imag} */,
  {32'h3f44aaa2, 32'h00000000} /* (14, 9, 30) {real, imag} */,
  {32'h3fb39809, 32'h00000000} /* (14, 9, 29) {real, imag} */,
  {32'h3fab7bfa, 32'h00000000} /* (14, 9, 28) {real, imag} */,
  {32'h3f9d585e, 32'h00000000} /* (14, 9, 27) {real, imag} */,
  {32'h3fb97481, 32'h00000000} /* (14, 9, 26) {real, imag} */,
  {32'h3f6f9a6a, 32'h00000000} /* (14, 9, 25) {real, imag} */,
  {32'h3f99e443, 32'h00000000} /* (14, 9, 24) {real, imag} */,
  {32'h3f1da900, 32'h00000000} /* (14, 9, 23) {real, imag} */,
  {32'h3f8b303b, 32'h00000000} /* (14, 9, 22) {real, imag} */,
  {32'h3f8705fb, 32'h00000000} /* (14, 9, 21) {real, imag} */,
  {32'hbed3e6ea, 32'h00000000} /* (14, 9, 20) {real, imag} */,
  {32'hbf77c760, 32'h00000000} /* (14, 9, 19) {real, imag} */,
  {32'hbfe14b28, 32'h00000000} /* (14, 9, 18) {real, imag} */,
  {32'hbf98a4c0, 32'h00000000} /* (14, 9, 17) {real, imag} */,
  {32'hbf23e3ae, 32'h00000000} /* (14, 9, 16) {real, imag} */,
  {32'hbf63c8fc, 32'h00000000} /* (14, 9, 15) {real, imag} */,
  {32'hbf80224b, 32'h00000000} /* (14, 9, 14) {real, imag} */,
  {32'hbf48b01b, 32'h00000000} /* (14, 9, 13) {real, imag} */,
  {32'hbf0f02eb, 32'h00000000} /* (14, 9, 12) {real, imag} */,
  {32'hbf092a61, 32'h00000000} /* (14, 9, 11) {real, imag} */,
  {32'h3ec5f896, 32'h00000000} /* (14, 9, 10) {real, imag} */,
  {32'h3efdeffc, 32'h00000000} /* (14, 9, 9) {real, imag} */,
  {32'h3f253590, 32'h00000000} /* (14, 9, 8) {real, imag} */,
  {32'h3f13b05b, 32'h00000000} /* (14, 9, 7) {real, imag} */,
  {32'h3f10cd41, 32'h00000000} /* (14, 9, 6) {real, imag} */,
  {32'h3f831ee2, 32'h00000000} /* (14, 9, 5) {real, imag} */,
  {32'h3f948f95, 32'h00000000} /* (14, 9, 4) {real, imag} */,
  {32'h3fb82a9f, 32'h00000000} /* (14, 9, 3) {real, imag} */,
  {32'h3fd9f73a, 32'h00000000} /* (14, 9, 2) {real, imag} */,
  {32'h3fbe77b2, 32'h00000000} /* (14, 9, 1) {real, imag} */,
  {32'h3f35bdaf, 32'h00000000} /* (14, 9, 0) {real, imag} */,
  {32'h3ec574cc, 32'h00000000} /* (14, 8, 31) {real, imag} */,
  {32'h3f38548e, 32'h00000000} /* (14, 8, 30) {real, imag} */,
  {32'h3f0d481e, 32'h00000000} /* (14, 8, 29) {real, imag} */,
  {32'h3f31264b, 32'h00000000} /* (14, 8, 28) {real, imag} */,
  {32'h3f0ab450, 32'h00000000} /* (14, 8, 27) {real, imag} */,
  {32'h3f60cec1, 32'h00000000} /* (14, 8, 26) {real, imag} */,
  {32'h3f80ade5, 32'h00000000} /* (14, 8, 25) {real, imag} */,
  {32'h3fc3c20e, 32'h00000000} /* (14, 8, 24) {real, imag} */,
  {32'h3f5d15e6, 32'h00000000} /* (14, 8, 23) {real, imag} */,
  {32'h3f915002, 32'h00000000} /* (14, 8, 22) {real, imag} */,
  {32'h3f11bb85, 32'h00000000} /* (14, 8, 21) {real, imag} */,
  {32'hbee99d2c, 32'h00000000} /* (14, 8, 20) {real, imag} */,
  {32'hbf4d1915, 32'h00000000} /* (14, 8, 19) {real, imag} */,
  {32'hbf7367dd, 32'h00000000} /* (14, 8, 18) {real, imag} */,
  {32'hbf283be8, 32'h00000000} /* (14, 8, 17) {real, imag} */,
  {32'hbf2a88e5, 32'h00000000} /* (14, 8, 16) {real, imag} */,
  {32'hbf70b385, 32'h00000000} /* (14, 8, 15) {real, imag} */,
  {32'hbf7572a9, 32'h00000000} /* (14, 8, 14) {real, imag} */,
  {32'hbf57ceda, 32'h00000000} /* (14, 8, 13) {real, imag} */,
  {32'hbf00b1dd, 32'h00000000} /* (14, 8, 12) {real, imag} */,
  {32'hbf199915, 32'h00000000} /* (14, 8, 11) {real, imag} */,
  {32'h3ee3f5de, 32'h00000000} /* (14, 8, 10) {real, imag} */,
  {32'h3f2ddee6, 32'h00000000} /* (14, 8, 9) {real, imag} */,
  {32'h3f0e0cae, 32'h00000000} /* (14, 8, 8) {real, imag} */,
  {32'h3f88fdb1, 32'h00000000} /* (14, 8, 7) {real, imag} */,
  {32'h3fb8d042, 32'h00000000} /* (14, 8, 6) {real, imag} */,
  {32'h3fb4867c, 32'h00000000} /* (14, 8, 5) {real, imag} */,
  {32'h3eecc566, 32'h00000000} /* (14, 8, 4) {real, imag} */,
  {32'h3f6bc6cc, 32'h00000000} /* (14, 8, 3) {real, imag} */,
  {32'h3fc2e14f, 32'h00000000} /* (14, 8, 2) {real, imag} */,
  {32'h3fa0371b, 32'h00000000} /* (14, 8, 1) {real, imag} */,
  {32'h3ec5d586, 32'h00000000} /* (14, 8, 0) {real, imag} */,
  {32'h3f04132b, 32'h00000000} /* (14, 7, 31) {real, imag} */,
  {32'h3f3d856f, 32'h00000000} /* (14, 7, 30) {real, imag} */,
  {32'h3f0dc508, 32'h00000000} /* (14, 7, 29) {real, imag} */,
  {32'h3f059849, 32'h00000000} /* (14, 7, 28) {real, imag} */,
  {32'h3ef77ad2, 32'h00000000} /* (14, 7, 27) {real, imag} */,
  {32'h3f61ce30, 32'h00000000} /* (14, 7, 26) {real, imag} */,
  {32'h3f384011, 32'h00000000} /* (14, 7, 25) {real, imag} */,
  {32'h3f8298e4, 32'h00000000} /* (14, 7, 24) {real, imag} */,
  {32'h3f763362, 32'h00000000} /* (14, 7, 23) {real, imag} */,
  {32'h3fba8e4e, 32'h00000000} /* (14, 7, 22) {real, imag} */,
  {32'h3e252cc6, 32'h00000000} /* (14, 7, 21) {real, imag} */,
  {32'hbf94d323, 32'h00000000} /* (14, 7, 20) {real, imag} */,
  {32'hbf449921, 32'h00000000} /* (14, 7, 19) {real, imag} */,
  {32'hbf4e761f, 32'h00000000} /* (14, 7, 18) {real, imag} */,
  {32'hbf65145b, 32'h00000000} /* (14, 7, 17) {real, imag} */,
  {32'hbf1179c8, 32'h00000000} /* (14, 7, 16) {real, imag} */,
  {32'hbf399d57, 32'h00000000} /* (14, 7, 15) {real, imag} */,
  {32'hbf87916d, 32'h00000000} /* (14, 7, 14) {real, imag} */,
  {32'hbf80cfc1, 32'h00000000} /* (14, 7, 13) {real, imag} */,
  {32'hbf0aa48f, 32'h00000000} /* (14, 7, 12) {real, imag} */,
  {32'hbee3a3be, 32'h00000000} /* (14, 7, 11) {real, imag} */,
  {32'h3f1fe9ae, 32'h00000000} /* (14, 7, 10) {real, imag} */,
  {32'h3f3acc9e, 32'h00000000} /* (14, 7, 9) {real, imag} */,
  {32'h3f79fa6f, 32'h00000000} /* (14, 7, 8) {real, imag} */,
  {32'h3fc58b71, 32'h00000000} /* (14, 7, 7) {real, imag} */,
  {32'h3faf6ef6, 32'h00000000} /* (14, 7, 6) {real, imag} */,
  {32'h3f96096a, 32'h00000000} /* (14, 7, 5) {real, imag} */,
  {32'h3f2f3797, 32'h00000000} /* (14, 7, 4) {real, imag} */,
  {32'h3f4dd3a1, 32'h00000000} /* (14, 7, 3) {real, imag} */,
  {32'h3f8c263b, 32'h00000000} /* (14, 7, 2) {real, imag} */,
  {32'h3f75781c, 32'h00000000} /* (14, 7, 1) {real, imag} */,
  {32'h3ee98179, 32'h00000000} /* (14, 7, 0) {real, imag} */,
  {32'h3ea8231c, 32'h00000000} /* (14, 6, 31) {real, imag} */,
  {32'h3eb0a266, 32'h00000000} /* (14, 6, 30) {real, imag} */,
  {32'h3ed41060, 32'h00000000} /* (14, 6, 29) {real, imag} */,
  {32'h3f16d362, 32'h00000000} /* (14, 6, 28) {real, imag} */,
  {32'h3f950c37, 32'h00000000} /* (14, 6, 27) {real, imag} */,
  {32'h3f9168ba, 32'h00000000} /* (14, 6, 26) {real, imag} */,
  {32'h3f34e934, 32'h00000000} /* (14, 6, 25) {real, imag} */,
  {32'h3f1e6327, 32'h00000000} /* (14, 6, 24) {real, imag} */,
  {32'h3f5e93ca, 32'h00000000} /* (14, 6, 23) {real, imag} */,
  {32'h3fa44249, 32'h00000000} /* (14, 6, 22) {real, imag} */,
  {32'h3f15087a, 32'h00000000} /* (14, 6, 21) {real, imag} */,
  {32'hbf49346e, 32'h00000000} /* (14, 6, 20) {real, imag} */,
  {32'hbf5557e1, 32'h00000000} /* (14, 6, 19) {real, imag} */,
  {32'hbf82d746, 32'h00000000} /* (14, 6, 18) {real, imag} */,
  {32'hbf7c7474, 32'h00000000} /* (14, 6, 17) {real, imag} */,
  {32'hbecef5ec, 32'h00000000} /* (14, 6, 16) {real, imag} */,
  {32'hbf2cf07a, 32'h00000000} /* (14, 6, 15) {real, imag} */,
  {32'hbf913d18, 32'h00000000} /* (14, 6, 14) {real, imag} */,
  {32'hbf7566a7, 32'h00000000} /* (14, 6, 13) {real, imag} */,
  {32'hbf541149, 32'h00000000} /* (14, 6, 12) {real, imag} */,
  {32'hbf19d562, 32'h00000000} /* (14, 6, 11) {real, imag} */,
  {32'h3e1fd2ed, 32'h00000000} /* (14, 6, 10) {real, imag} */,
  {32'h3f38c29b, 32'h00000000} /* (14, 6, 9) {real, imag} */,
  {32'h3f8ac8da, 32'h00000000} /* (14, 6, 8) {real, imag} */,
  {32'h3f684983, 32'h00000000} /* (14, 6, 7) {real, imag} */,
  {32'h3f5dadd5, 32'h00000000} /* (14, 6, 6) {real, imag} */,
  {32'h3f3b2372, 32'h00000000} /* (14, 6, 5) {real, imag} */,
  {32'h3faebc52, 32'h00000000} /* (14, 6, 4) {real, imag} */,
  {32'h3f961c4a, 32'h00000000} /* (14, 6, 3) {real, imag} */,
  {32'h3f4db663, 32'h00000000} /* (14, 6, 2) {real, imag} */,
  {32'h3f98102d, 32'h00000000} /* (14, 6, 1) {real, imag} */,
  {32'h3f1a7360, 32'h00000000} /* (14, 6, 0) {real, imag} */,
  {32'h3eab3f5c, 32'h00000000} /* (14, 5, 31) {real, imag} */,
  {32'h3f43ab02, 32'h00000000} /* (14, 5, 30) {real, imag} */,
  {32'h3f4e2b10, 32'h00000000} /* (14, 5, 29) {real, imag} */,
  {32'h3f942e2b, 32'h00000000} /* (14, 5, 28) {real, imag} */,
  {32'h3f9e7c71, 32'h00000000} /* (14, 5, 27) {real, imag} */,
  {32'h3f2d4ba6, 32'h00000000} /* (14, 5, 26) {real, imag} */,
  {32'h3ea704a6, 32'h00000000} /* (14, 5, 25) {real, imag} */,
  {32'h3f423545, 32'h00000000} /* (14, 5, 24) {real, imag} */,
  {32'h3f24f740, 32'h00000000} /* (14, 5, 23) {real, imag} */,
  {32'h3f954372, 32'h00000000} /* (14, 5, 22) {real, imag} */,
  {32'h3f8fe9a1, 32'h00000000} /* (14, 5, 21) {real, imag} */,
  {32'h3ec11661, 32'h00000000} /* (14, 5, 20) {real, imag} */,
  {32'hbe8515f2, 32'h00000000} /* (14, 5, 19) {real, imag} */,
  {32'hbee835b3, 32'h00000000} /* (14, 5, 18) {real, imag} */,
  {32'hbdf8c550, 32'h00000000} /* (14, 5, 17) {real, imag} */,
  {32'h3e269318, 32'h00000000} /* (14, 5, 16) {real, imag} */,
  {32'hbf31e6ab, 32'h00000000} /* (14, 5, 15) {real, imag} */,
  {32'hbfb81b1c, 32'h00000000} /* (14, 5, 14) {real, imag} */,
  {32'hbf679e04, 32'h00000000} /* (14, 5, 13) {real, imag} */,
  {32'hbf3e1a43, 32'h00000000} /* (14, 5, 12) {real, imag} */,
  {32'hbf5d6dc4, 32'h00000000} /* (14, 5, 11) {real, imag} */,
  {32'hbf8ad534, 32'h00000000} /* (14, 5, 10) {real, imag} */,
  {32'hbf7d0b56, 32'h00000000} /* (14, 5, 9) {real, imag} */,
  {32'hbf42eb13, 32'h00000000} /* (14, 5, 8) {real, imag} */,
  {32'hbf20bdde, 32'h00000000} /* (14, 5, 7) {real, imag} */,
  {32'h3c9d5921, 32'h00000000} /* (14, 5, 6) {real, imag} */,
  {32'h3ef44035, 32'h00000000} /* (14, 5, 5) {real, imag} */,
  {32'h3f66d890, 32'h00000000} /* (14, 5, 4) {real, imag} */,
  {32'h3f9dcb2d, 32'h00000000} /* (14, 5, 3) {real, imag} */,
  {32'h3f8b7c8f, 32'h00000000} /* (14, 5, 2) {real, imag} */,
  {32'h3f499719, 32'h00000000} /* (14, 5, 1) {real, imag} */,
  {32'h3ec56cf3, 32'h00000000} /* (14, 5, 0) {real, imag} */,
  {32'h3f014bf4, 32'h00000000} /* (14, 4, 31) {real, imag} */,
  {32'h3f6124d8, 32'h00000000} /* (14, 4, 30) {real, imag} */,
  {32'h3f814b9f, 32'h00000000} /* (14, 4, 29) {real, imag} */,
  {32'h3f9e9073, 32'h00000000} /* (14, 4, 28) {real, imag} */,
  {32'h3f9cb7cc, 32'h00000000} /* (14, 4, 27) {real, imag} */,
  {32'h3f47866a, 32'h00000000} /* (14, 4, 26) {real, imag} */,
  {32'h3f18cce9, 32'h00000000} /* (14, 4, 25) {real, imag} */,
  {32'h3f84a8ec, 32'h00000000} /* (14, 4, 24) {real, imag} */,
  {32'h3f888802, 32'h00000000} /* (14, 4, 23) {real, imag} */,
  {32'h3fdf53bb, 32'h00000000} /* (14, 4, 22) {real, imag} */,
  {32'h3feb5efa, 32'h00000000} /* (14, 4, 21) {real, imag} */,
  {32'h3fa68ebb, 32'h00000000} /* (14, 4, 20) {real, imag} */,
  {32'h3ec31ff5, 32'h00000000} /* (14, 4, 19) {real, imag} */,
  {32'h3eefd9e5, 32'h00000000} /* (14, 4, 18) {real, imag} */,
  {32'h3f2ed119, 32'h00000000} /* (14, 4, 17) {real, imag} */,
  {32'h3f3d8700, 32'h00000000} /* (14, 4, 16) {real, imag} */,
  {32'hbe7a0ec9, 32'h00000000} /* (14, 4, 15) {real, imag} */,
  {32'hbf4623f5, 32'h00000000} /* (14, 4, 14) {real, imag} */,
  {32'hbf4084a9, 32'h00000000} /* (14, 4, 13) {real, imag} */,
  {32'hbef5c3a5, 32'h00000000} /* (14, 4, 12) {real, imag} */,
  {32'hbf29a188, 32'h00000000} /* (14, 4, 11) {real, imag} */,
  {32'hbf8aaf91, 32'h00000000} /* (14, 4, 10) {real, imag} */,
  {32'hbfdd35e0, 32'h00000000} /* (14, 4, 9) {real, imag} */,
  {32'hbfb059eb, 32'h00000000} /* (14, 4, 8) {real, imag} */,
  {32'hbf66fa0d, 32'h00000000} /* (14, 4, 7) {real, imag} */,
  {32'hbefcde92, 32'h00000000} /* (14, 4, 6) {real, imag} */,
  {32'h3e51d7fb, 32'h00000000} /* (14, 4, 5) {real, imag} */,
  {32'h3f2e8508, 32'h00000000} /* (14, 4, 4) {real, imag} */,
  {32'h3f9ccb79, 32'h00000000} /* (14, 4, 3) {real, imag} */,
  {32'h3fa73515, 32'h00000000} /* (14, 4, 2) {real, imag} */,
  {32'h3f3b2e35, 32'h00000000} /* (14, 4, 1) {real, imag} */,
  {32'h3ecae097, 32'h00000000} /* (14, 4, 0) {real, imag} */,
  {32'h3f88b304, 32'h00000000} /* (14, 3, 31) {real, imag} */,
  {32'h3f45519b, 32'h00000000} /* (14, 3, 30) {real, imag} */,
  {32'h3eecfb3e, 32'h00000000} /* (14, 3, 29) {real, imag} */,
  {32'h3f840efe, 32'h00000000} /* (14, 3, 28) {real, imag} */,
  {32'h3fc591ea, 32'h00000000} /* (14, 3, 27) {real, imag} */,
  {32'h3f7ac844, 32'h00000000} /* (14, 3, 26) {real, imag} */,
  {32'h3f2e2442, 32'h00000000} /* (14, 3, 25) {real, imag} */,
  {32'h3f98167a, 32'h00000000} /* (14, 3, 24) {real, imag} */,
  {32'h3f825ed7, 32'h00000000} /* (14, 3, 23) {real, imag} */,
  {32'h3fbd375b, 32'h00000000} /* (14, 3, 22) {real, imag} */,
  {32'h3faff7da, 32'h00000000} /* (14, 3, 21) {real, imag} */,
  {32'h3f88920a, 32'h00000000} /* (14, 3, 20) {real, imag} */,
  {32'h3f272be3, 32'h00000000} /* (14, 3, 19) {real, imag} */,
  {32'h3fa4b934, 32'h00000000} /* (14, 3, 18) {real, imag} */,
  {32'h3f57fe52, 32'h00000000} /* (14, 3, 17) {real, imag} */,
  {32'h3f1f4aa7, 32'h00000000} /* (14, 3, 16) {real, imag} */,
  {32'hbee17aea, 32'h00000000} /* (14, 3, 15) {real, imag} */,
  {32'hbf0b0700, 32'h00000000} /* (14, 3, 14) {real, imag} */,
  {32'hbf472885, 32'h00000000} /* (14, 3, 13) {real, imag} */,
  {32'hbf4ae164, 32'h00000000} /* (14, 3, 12) {real, imag} */,
  {32'hbf6443dd, 32'h00000000} /* (14, 3, 11) {real, imag} */,
  {32'hbf32665e, 32'h00000000} /* (14, 3, 10) {real, imag} */,
  {32'hbf7daeba, 32'h00000000} /* (14, 3, 9) {real, imag} */,
  {32'hbf439bf4, 32'h00000000} /* (14, 3, 8) {real, imag} */,
  {32'hbed3bef5, 32'h00000000} /* (14, 3, 7) {real, imag} */,
  {32'hbe9e82bc, 32'h00000000} /* (14, 3, 6) {real, imag} */,
  {32'h3f291eb1, 32'h00000000} /* (14, 3, 5) {real, imag} */,
  {32'h3fa485fb, 32'h00000000} /* (14, 3, 4) {real, imag} */,
  {32'h3fa20a77, 32'h00000000} /* (14, 3, 3) {real, imag} */,
  {32'h3f3ae4a8, 32'h00000000} /* (14, 3, 2) {real, imag} */,
  {32'h3ed1b7e1, 32'h00000000} /* (14, 3, 1) {real, imag} */,
  {32'h3f1e0fc7, 32'h00000000} /* (14, 3, 0) {real, imag} */,
  {32'h3f541c1f, 32'h00000000} /* (14, 2, 31) {real, imag} */,
  {32'h3f9557bf, 32'h00000000} /* (14, 2, 30) {real, imag} */,
  {32'h3f18c9e1, 32'h00000000} /* (14, 2, 29) {real, imag} */,
  {32'h3f690a66, 32'h00000000} /* (14, 2, 28) {real, imag} */,
  {32'h3f71154f, 32'h00000000} /* (14, 2, 27) {real, imag} */,
  {32'h3f38eab0, 32'h00000000} /* (14, 2, 26) {real, imag} */,
  {32'h3f1fd844, 32'h00000000} /* (14, 2, 25) {real, imag} */,
  {32'h3f941ddf, 32'h00000000} /* (14, 2, 24) {real, imag} */,
  {32'h3f512684, 32'h00000000} /* (14, 2, 23) {real, imag} */,
  {32'h3f4b276f, 32'h00000000} /* (14, 2, 22) {real, imag} */,
  {32'h3f64bda9, 32'h00000000} /* (14, 2, 21) {real, imag} */,
  {32'h3f085c6c, 32'h00000000} /* (14, 2, 20) {real, imag} */,
  {32'h3f320fae, 32'h00000000} /* (14, 2, 19) {real, imag} */,
  {32'h3f4ca4ac, 32'h00000000} /* (14, 2, 18) {real, imag} */,
  {32'h3f61e459, 32'h00000000} /* (14, 2, 17) {real, imag} */,
  {32'h3f3e33ff, 32'h00000000} /* (14, 2, 16) {real, imag} */,
  {32'hbf0425b8, 32'h00000000} /* (14, 2, 15) {real, imag} */,
  {32'hbeea53ac, 32'h00000000} /* (14, 2, 14) {real, imag} */,
  {32'hbf5593a3, 32'h00000000} /* (14, 2, 13) {real, imag} */,
  {32'hbf7a7b43, 32'h00000000} /* (14, 2, 12) {real, imag} */,
  {32'hbf2dd0b3, 32'h00000000} /* (14, 2, 11) {real, imag} */,
  {32'hbf189244, 32'h00000000} /* (14, 2, 10) {real, imag} */,
  {32'hbf67be00, 32'h00000000} /* (14, 2, 9) {real, imag} */,
  {32'hbf1b9a4c, 32'h00000000} /* (14, 2, 8) {real, imag} */,
  {32'hbf1a43da, 32'h00000000} /* (14, 2, 7) {real, imag} */,
  {32'hbf1cb2eb, 32'h00000000} /* (14, 2, 6) {real, imag} */,
  {32'h3e8db55b, 32'h00000000} /* (14, 2, 5) {real, imag} */,
  {32'h3f85f1ed, 32'h00000000} /* (14, 2, 4) {real, imag} */,
  {32'h3fc48e28, 32'h00000000} /* (14, 2, 3) {real, imag} */,
  {32'h3f9be975, 32'h00000000} /* (14, 2, 2) {real, imag} */,
  {32'h3ed1457a, 32'h00000000} /* (14, 2, 1) {real, imag} */,
  {32'h3e7a44ca, 32'h00000000} /* (14, 2, 0) {real, imag} */,
  {32'h3e591788, 32'h00000000} /* (14, 1, 31) {real, imag} */,
  {32'h3f5bae59, 32'h00000000} /* (14, 1, 30) {real, imag} */,
  {32'h3f70f373, 32'h00000000} /* (14, 1, 29) {real, imag} */,
  {32'h3f901a57, 32'h00000000} /* (14, 1, 28) {real, imag} */,
  {32'h3f6fb428, 32'h00000000} /* (14, 1, 27) {real, imag} */,
  {32'h3f163628, 32'h00000000} /* (14, 1, 26) {real, imag} */,
  {32'h3f3bfa84, 32'h00000000} /* (14, 1, 25) {real, imag} */,
  {32'h3f725d04, 32'h00000000} /* (14, 1, 24) {real, imag} */,
  {32'h3efb329f, 32'h00000000} /* (14, 1, 23) {real, imag} */,
  {32'h3f39b23a, 32'h00000000} /* (14, 1, 22) {real, imag} */,
  {32'h3f279cf0, 32'h00000000} /* (14, 1, 21) {real, imag} */,
  {32'h3f217845, 32'h00000000} /* (14, 1, 20) {real, imag} */,
  {32'h3f5380b0, 32'h00000000} /* (14, 1, 19) {real, imag} */,
  {32'h3f00c626, 32'h00000000} /* (14, 1, 18) {real, imag} */,
  {32'h3f270b5c, 32'h00000000} /* (14, 1, 17) {real, imag} */,
  {32'h3f0c4bb5, 32'h00000000} /* (14, 1, 16) {real, imag} */,
  {32'hbe78caf9, 32'h00000000} /* (14, 1, 15) {real, imag} */,
  {32'hbf18643e, 32'h00000000} /* (14, 1, 14) {real, imag} */,
  {32'hbf89c8c6, 32'h00000000} /* (14, 1, 13) {real, imag} */,
  {32'hbf706916, 32'h00000000} /* (14, 1, 12) {real, imag} */,
  {32'hbf44e243, 32'h00000000} /* (14, 1, 11) {real, imag} */,
  {32'hbfa3f226, 32'h00000000} /* (14, 1, 10) {real, imag} */,
  {32'hbf996238, 32'h00000000} /* (14, 1, 9) {real, imag} */,
  {32'hbf918732, 32'h00000000} /* (14, 1, 8) {real, imag} */,
  {32'hbf6efa39, 32'h00000000} /* (14, 1, 7) {real, imag} */,
  {32'hbf55959c, 32'h00000000} /* (14, 1, 6) {real, imag} */,
  {32'h3e22f0b9, 32'h00000000} /* (14, 1, 5) {real, imag} */,
  {32'h3ed3f5e8, 32'h00000000} /* (14, 1, 4) {real, imag} */,
  {32'h3f4732b7, 32'h00000000} /* (14, 1, 3) {real, imag} */,
  {32'h3f6f869c, 32'h00000000} /* (14, 1, 2) {real, imag} */,
  {32'h3e759a04, 32'h00000000} /* (14, 1, 1) {real, imag} */,
  {32'hbdbf6ce4, 32'h00000000} /* (14, 1, 0) {real, imag} */,
  {32'h3d154c3f, 32'h00000000} /* (14, 0, 31) {real, imag} */,
  {32'h3e9bbbdb, 32'h00000000} /* (14, 0, 30) {real, imag} */,
  {32'h3eff61ee, 32'h00000000} /* (14, 0, 29) {real, imag} */,
  {32'h3f3cb576, 32'h00000000} /* (14, 0, 28) {real, imag} */,
  {32'h3f75cde1, 32'h00000000} /* (14, 0, 27) {real, imag} */,
  {32'h3f1ccc8d, 32'h00000000} /* (14, 0, 26) {real, imag} */,
  {32'h3eb20349, 32'h00000000} /* (14, 0, 25) {real, imag} */,
  {32'h3eb70aec, 32'h00000000} /* (14, 0, 24) {real, imag} */,
  {32'h3eb96a8e, 32'h00000000} /* (14, 0, 23) {real, imag} */,
  {32'h3ec56bd0, 32'h00000000} /* (14, 0, 22) {real, imag} */,
  {32'h3e73a76f, 32'h00000000} /* (14, 0, 21) {real, imag} */,
  {32'h3ee227e1, 32'h00000000} /* (14, 0, 20) {real, imag} */,
  {32'h3ee74204, 32'h00000000} /* (14, 0, 19) {real, imag} */,
  {32'h3eeef61b, 32'h00000000} /* (14, 0, 18) {real, imag} */,
  {32'h3e6c00dd, 32'h00000000} /* (14, 0, 17) {real, imag} */,
  {32'h3e0c083e, 32'h00000000} /* (14, 0, 16) {real, imag} */,
  {32'hbe8361a9, 32'h00000000} /* (14, 0, 15) {real, imag} */,
  {32'hbf360db2, 32'h00000000} /* (14, 0, 14) {real, imag} */,
  {32'hbf5a84ac, 32'h00000000} /* (14, 0, 13) {real, imag} */,
  {32'hbf0d374f, 32'h00000000} /* (14, 0, 12) {real, imag} */,
  {32'hbf14df53, 32'h00000000} /* (14, 0, 11) {real, imag} */,
  {32'hbf4de882, 32'h00000000} /* (14, 0, 10) {real, imag} */,
  {32'hbef7072d, 32'h00000000} /* (14, 0, 9) {real, imag} */,
  {32'hbf47d8ab, 32'h00000000} /* (14, 0, 8) {real, imag} */,
  {32'hbf33518f, 32'h00000000} /* (14, 0, 7) {real, imag} */,
  {32'hbeef6481, 32'h00000000} /* (14, 0, 6) {real, imag} */,
  {32'h3d079ccb, 32'h00000000} /* (14, 0, 5) {real, imag} */,
  {32'h3e350e29, 32'h00000000} /* (14, 0, 4) {real, imag} */,
  {32'h3ee4546b, 32'h00000000} /* (14, 0, 3) {real, imag} */,
  {32'h3e924968, 32'h00000000} /* (14, 0, 2) {real, imag} */,
  {32'hbd1c2144, 32'h00000000} /* (14, 0, 1) {real, imag} */,
  {32'hbd9df948, 32'h00000000} /* (14, 0, 0) {real, imag} */,
  {32'h3ec6e8e0, 32'h00000000} /* (13, 31, 31) {real, imag} */,
  {32'h3f8e639f, 32'h00000000} /* (13, 31, 30) {real, imag} */,
  {32'h3f50fb88, 32'h00000000} /* (13, 31, 29) {real, imag} */,
  {32'h3f064c27, 32'h00000000} /* (13, 31, 28) {real, imag} */,
  {32'h3f1b6cab, 32'h00000000} /* (13, 31, 27) {real, imag} */,
  {32'h3f914c10, 32'h00000000} /* (13, 31, 26) {real, imag} */,
  {32'h3f28d03d, 32'h00000000} /* (13, 31, 25) {real, imag} */,
  {32'h3f23fc3a, 32'h00000000} /* (13, 31, 24) {real, imag} */,
  {32'h3efa978e, 32'h00000000} /* (13, 31, 23) {real, imag} */,
  {32'h3ece25b7, 32'h00000000} /* (13, 31, 22) {real, imag} */,
  {32'hbd5e38ef, 32'h00000000} /* (13, 31, 21) {real, imag} */,
  {32'hbe8e1d82, 32'h00000000} /* (13, 31, 20) {real, imag} */,
  {32'hbe99497b, 32'h00000000} /* (13, 31, 19) {real, imag} */,
  {32'hbf009c3b, 32'h00000000} /* (13, 31, 18) {real, imag} */,
  {32'hbef835ad, 32'h00000000} /* (13, 31, 17) {real, imag} */,
  {32'hbe87db24, 32'h00000000} /* (13, 31, 16) {real, imag} */,
  {32'hbedb82d3, 32'h00000000} /* (13, 31, 15) {real, imag} */,
  {32'hbf1661f2, 32'h00000000} /* (13, 31, 14) {real, imag} */,
  {32'hbf2843cb, 32'h00000000} /* (13, 31, 13) {real, imag} */,
  {32'hbe73c594, 32'h00000000} /* (13, 31, 12) {real, imag} */,
  {32'hbe2a78d1, 32'h00000000} /* (13, 31, 11) {real, imag} */,
  {32'h3df81b80, 32'h00000000} /* (13, 31, 10) {real, imag} */,
  {32'h3ed40f3a, 32'h00000000} /* (13, 31, 9) {real, imag} */,
  {32'hbd993998, 32'h00000000} /* (13, 31, 8) {real, imag} */,
  {32'h3dc3100e, 32'h00000000} /* (13, 31, 7) {real, imag} */,
  {32'h3f2ca6a4, 32'h00000000} /* (13, 31, 6) {real, imag} */,
  {32'h3f696814, 32'h00000000} /* (13, 31, 5) {real, imag} */,
  {32'h3f2b31cb, 32'h00000000} /* (13, 31, 4) {real, imag} */,
  {32'h3e47fac2, 32'h00000000} /* (13, 31, 3) {real, imag} */,
  {32'h3e0d0381, 32'h00000000} /* (13, 31, 2) {real, imag} */,
  {32'h3de71549, 32'h00000000} /* (13, 31, 1) {real, imag} */,
  {32'h3db19230, 32'h00000000} /* (13, 31, 0) {real, imag} */,
  {32'h3f1a6777, 32'h00000000} /* (13, 30, 31) {real, imag} */,
  {32'h3f8b15f7, 32'h00000000} /* (13, 30, 30) {real, imag} */,
  {32'h3f55efbc, 32'h00000000} /* (13, 30, 29) {real, imag} */,
  {32'h3ef51409, 32'h00000000} /* (13, 30, 28) {real, imag} */,
  {32'h3f0de034, 32'h00000000} /* (13, 30, 27) {real, imag} */,
  {32'h3f8e7605, 32'h00000000} /* (13, 30, 26) {real, imag} */,
  {32'h3fc229b8, 32'h00000000} /* (13, 30, 25) {real, imag} */,
  {32'h3fa46ecc, 32'h00000000} /* (13, 30, 24) {real, imag} */,
  {32'h3f9cac7e, 32'h00000000} /* (13, 30, 23) {real, imag} */,
  {32'h3fadd736, 32'h00000000} /* (13, 30, 22) {real, imag} */,
  {32'hbcbd358e, 32'h00000000} /* (13, 30, 21) {real, imag} */,
  {32'hbf7a5c59, 32'h00000000} /* (13, 30, 20) {real, imag} */,
  {32'hbf7a98fd, 32'h00000000} /* (13, 30, 19) {real, imag} */,
  {32'hbf991b25, 32'h00000000} /* (13, 30, 18) {real, imag} */,
  {32'hbf6b867c, 32'h00000000} /* (13, 30, 17) {real, imag} */,
  {32'hbf1c0586, 32'h00000000} /* (13, 30, 16) {real, imag} */,
  {32'hbf8c932a, 32'h00000000} /* (13, 30, 15) {real, imag} */,
  {32'hbf8a1d80, 32'h00000000} /* (13, 30, 14) {real, imag} */,
  {32'hbf6e816b, 32'h00000000} /* (13, 30, 13) {real, imag} */,
  {32'hbf0589f4, 32'h00000000} /* (13, 30, 12) {real, imag} */,
  {32'hbeac8269, 32'h00000000} /* (13, 30, 11) {real, imag} */,
  {32'h3f02a743, 32'h00000000} /* (13, 30, 10) {real, imag} */,
  {32'h3fada791, 32'h00000000} /* (13, 30, 9) {real, imag} */,
  {32'h3f03ec4a, 32'h00000000} /* (13, 30, 8) {real, imag} */,
  {32'h3eedacac, 32'h00000000} /* (13, 30, 7) {real, imag} */,
  {32'h3fb38195, 32'h00000000} /* (13, 30, 6) {real, imag} */,
  {32'h3f83ca96, 32'h00000000} /* (13, 30, 5) {real, imag} */,
  {32'h3f751b4f, 32'h00000000} /* (13, 30, 4) {real, imag} */,
  {32'h3f2ec5c8, 32'h00000000} /* (13, 30, 3) {real, imag} */,
  {32'h3ef52497, 32'h00000000} /* (13, 30, 2) {real, imag} */,
  {32'h3ed4e592, 32'h00000000} /* (13, 30, 1) {real, imag} */,
  {32'h3e560c0a, 32'h00000000} /* (13, 30, 0) {real, imag} */,
  {32'h3f22fcd6, 32'h00000000} /* (13, 29, 31) {real, imag} */,
  {32'h3fa174f9, 32'h00000000} /* (13, 29, 30) {real, imag} */,
  {32'h3f5b9170, 32'h00000000} /* (13, 29, 29) {real, imag} */,
  {32'h3db5bf53, 32'h00000000} /* (13, 29, 28) {real, imag} */,
  {32'h3eb0f6be, 32'h00000000} /* (13, 29, 27) {real, imag} */,
  {32'h3f7311c3, 32'h00000000} /* (13, 29, 26) {real, imag} */,
  {32'h3f90df3e, 32'h00000000} /* (13, 29, 25) {real, imag} */,
  {32'h3f1e635a, 32'h00000000} /* (13, 29, 24) {real, imag} */,
  {32'h3f94cffb, 32'h00000000} /* (13, 29, 23) {real, imag} */,
  {32'h3f946186, 32'h00000000} /* (13, 29, 22) {real, imag} */,
  {32'h3e6d76f2, 32'h00000000} /* (13, 29, 21) {real, imag} */,
  {32'hbf5ab000, 32'h00000000} /* (13, 29, 20) {real, imag} */,
  {32'hbf880e80, 32'h00000000} /* (13, 29, 19) {real, imag} */,
  {32'hbf7f3774, 32'h00000000} /* (13, 29, 18) {real, imag} */,
  {32'hbf8f06e3, 32'h00000000} /* (13, 29, 17) {real, imag} */,
  {32'hbf93f436, 32'h00000000} /* (13, 29, 16) {real, imag} */,
  {32'hbf9d8ba7, 32'h00000000} /* (13, 29, 15) {real, imag} */,
  {32'hbf73930c, 32'h00000000} /* (13, 29, 14) {real, imag} */,
  {32'hbf3d8f82, 32'h00000000} /* (13, 29, 13) {real, imag} */,
  {32'hbef37900, 32'h00000000} /* (13, 29, 12) {real, imag} */,
  {32'hbe8de4a2, 32'h00000000} /* (13, 29, 11) {real, imag} */,
  {32'h3f07b2bb, 32'h00000000} /* (13, 29, 10) {real, imag} */,
  {32'h3fa48efa, 32'h00000000} /* (13, 29, 9) {real, imag} */,
  {32'h3f1d5f14, 32'h00000000} /* (13, 29, 8) {real, imag} */,
  {32'h3f0c6e45, 32'h00000000} /* (13, 29, 7) {real, imag} */,
  {32'h3f92918d, 32'h00000000} /* (13, 29, 6) {real, imag} */,
  {32'h3f9f4168, 32'h00000000} /* (13, 29, 5) {real, imag} */,
  {32'h3f65529d, 32'h00000000} /* (13, 29, 4) {real, imag} */,
  {32'h3f42137a, 32'h00000000} /* (13, 29, 3) {real, imag} */,
  {32'h3f8e508f, 32'h00000000} /* (13, 29, 2) {real, imag} */,
  {32'h3fbc5da8, 32'h00000000} /* (13, 29, 1) {real, imag} */,
  {32'h3eeb3809, 32'h00000000} /* (13, 29, 0) {real, imag} */,
  {32'h3eac9c89, 32'h00000000} /* (13, 28, 31) {real, imag} */,
  {32'h3f85cd97, 32'h00000000} /* (13, 28, 30) {real, imag} */,
  {32'h3f6c0953, 32'h00000000} /* (13, 28, 29) {real, imag} */,
  {32'h3f466ac8, 32'h00000000} /* (13, 28, 28) {real, imag} */,
  {32'h3f8151a7, 32'h00000000} /* (13, 28, 27) {real, imag} */,
  {32'h3f5807fc, 32'h00000000} /* (13, 28, 26) {real, imag} */,
  {32'h3f281083, 32'h00000000} /* (13, 28, 25) {real, imag} */,
  {32'h3f35b261, 32'h00000000} /* (13, 28, 24) {real, imag} */,
  {32'h3f54e448, 32'h00000000} /* (13, 28, 23) {real, imag} */,
  {32'h3f144ea7, 32'h00000000} /* (13, 28, 22) {real, imag} */,
  {32'h3ee7f608, 32'h00000000} /* (13, 28, 21) {real, imag} */,
  {32'hbeba159f, 32'h00000000} /* (13, 28, 20) {real, imag} */,
  {32'hbf402427, 32'h00000000} /* (13, 28, 19) {real, imag} */,
  {32'hbf8da643, 32'h00000000} /* (13, 28, 18) {real, imag} */,
  {32'hbf922c65, 32'h00000000} /* (13, 28, 17) {real, imag} */,
  {32'hbf9868a3, 32'h00000000} /* (13, 28, 16) {real, imag} */,
  {32'hbf88189e, 32'h00000000} /* (13, 28, 15) {real, imag} */,
  {32'hbf482b4f, 32'h00000000} /* (13, 28, 14) {real, imag} */,
  {32'hbf1a395b, 32'h00000000} /* (13, 28, 13) {real, imag} */,
  {32'hbf2ffe22, 32'h00000000} /* (13, 28, 12) {real, imag} */,
  {32'hbf2daa43, 32'h00000000} /* (13, 28, 11) {real, imag} */,
  {32'h3de10838, 32'h00000000} /* (13, 28, 10) {real, imag} */,
  {32'h3f59d113, 32'h00000000} /* (13, 28, 9) {real, imag} */,
  {32'h3f4273d0, 32'h00000000} /* (13, 28, 8) {real, imag} */,
  {32'h3f4010bd, 32'h00000000} /* (13, 28, 7) {real, imag} */,
  {32'h3f89217e, 32'h00000000} /* (13, 28, 6) {real, imag} */,
  {32'h3fbd7b24, 32'h00000000} /* (13, 28, 5) {real, imag} */,
  {32'h3f252ba9, 32'h00000000} /* (13, 28, 4) {real, imag} */,
  {32'h3e7fcbc4, 32'h00000000} /* (13, 28, 3) {real, imag} */,
  {32'h3f3e988e, 32'h00000000} /* (13, 28, 2) {real, imag} */,
  {32'h3f69568f, 32'h00000000} /* (13, 28, 1) {real, imag} */,
  {32'h3ef3fbe7, 32'h00000000} /* (13, 28, 0) {real, imag} */,
  {32'h3ed8537a, 32'h00000000} /* (13, 27, 31) {real, imag} */,
  {32'h3f9a93bd, 32'h00000000} /* (13, 27, 30) {real, imag} */,
  {32'h3fb37d76, 32'h00000000} /* (13, 27, 29) {real, imag} */,
  {32'h3fc2e924, 32'h00000000} /* (13, 27, 28) {real, imag} */,
  {32'h3fae222d, 32'h00000000} /* (13, 27, 27) {real, imag} */,
  {32'h3f339521, 32'h00000000} /* (13, 27, 26) {real, imag} */,
  {32'h3f6453b8, 32'h00000000} /* (13, 27, 25) {real, imag} */,
  {32'h3f54b403, 32'h00000000} /* (13, 27, 24) {real, imag} */,
  {32'h3f4c2ba1, 32'h00000000} /* (13, 27, 23) {real, imag} */,
  {32'h3fa0ece0, 32'h00000000} /* (13, 27, 22) {real, imag} */,
  {32'h3f2506a1, 32'h00000000} /* (13, 27, 21) {real, imag} */,
  {32'hbd85dc2b, 32'h00000000} /* (13, 27, 20) {real, imag} */,
  {32'hbeddaed8, 32'h00000000} /* (13, 27, 19) {real, imag} */,
  {32'hbf888580, 32'h00000000} /* (13, 27, 18) {real, imag} */,
  {32'hbf6173d9, 32'h00000000} /* (13, 27, 17) {real, imag} */,
  {32'hbf5ff7c3, 32'h00000000} /* (13, 27, 16) {real, imag} */,
  {32'hbfaf93d1, 32'h00000000} /* (13, 27, 15) {real, imag} */,
  {32'hbf26d8b7, 32'h00000000} /* (13, 27, 14) {real, imag} */,
  {32'hbea28e36, 32'h00000000} /* (13, 27, 13) {real, imag} */,
  {32'hbf67b312, 32'h00000000} /* (13, 27, 12) {real, imag} */,
  {32'hbf8347fa, 32'h00000000} /* (13, 27, 11) {real, imag} */,
  {32'h3e09f04e, 32'h00000000} /* (13, 27, 10) {real, imag} */,
  {32'h3f712405, 32'h00000000} /* (13, 27, 9) {real, imag} */,
  {32'h3f8badc7, 32'h00000000} /* (13, 27, 8) {real, imag} */,
  {32'h3f875d45, 32'h00000000} /* (13, 27, 7) {real, imag} */,
  {32'h3f929209, 32'h00000000} /* (13, 27, 6) {real, imag} */,
  {32'h3f637d29, 32'h00000000} /* (13, 27, 5) {real, imag} */,
  {32'h3ee8baa1, 32'h00000000} /* (13, 27, 4) {real, imag} */,
  {32'h3f1cb22b, 32'h00000000} /* (13, 27, 3) {real, imag} */,
  {32'h3ef606ae, 32'h00000000} /* (13, 27, 2) {real, imag} */,
  {32'h3f1a4baa, 32'h00000000} /* (13, 27, 1) {real, imag} */,
  {32'h3f237170, 32'h00000000} /* (13, 27, 0) {real, imag} */,
  {32'h3f025504, 32'h00000000} /* (13, 26, 31) {real, imag} */,
  {32'h3f8812c5, 32'h00000000} /* (13, 26, 30) {real, imag} */,
  {32'h3faa9160, 32'h00000000} /* (13, 26, 29) {real, imag} */,
  {32'h3f8bbf7f, 32'h00000000} /* (13, 26, 28) {real, imag} */,
  {32'h3f634034, 32'h00000000} /* (13, 26, 27) {real, imag} */,
  {32'h3fb2cdbd, 32'h00000000} /* (13, 26, 26) {real, imag} */,
  {32'h3feb5faf, 32'h00000000} /* (13, 26, 25) {real, imag} */,
  {32'h3f2c9226, 32'h00000000} /* (13, 26, 24) {real, imag} */,
  {32'h3f5146cc, 32'h00000000} /* (13, 26, 23) {real, imag} */,
  {32'h3f93e2f1, 32'h00000000} /* (13, 26, 22) {real, imag} */,
  {32'h3e773808, 32'h00000000} /* (13, 26, 21) {real, imag} */,
  {32'hbece4b05, 32'h00000000} /* (13, 26, 20) {real, imag} */,
  {32'hbf1dc221, 32'h00000000} /* (13, 26, 19) {real, imag} */,
  {32'hbf7f5be2, 32'h00000000} /* (13, 26, 18) {real, imag} */,
  {32'hbf2d750e, 32'h00000000} /* (13, 26, 17) {real, imag} */,
  {32'hbf93f4a2, 32'h00000000} /* (13, 26, 16) {real, imag} */,
  {32'hbf891cc7, 32'h00000000} /* (13, 26, 15) {real, imag} */,
  {32'hbeea3afa, 32'h00000000} /* (13, 26, 14) {real, imag} */,
  {32'hbf126a1a, 32'h00000000} /* (13, 26, 13) {real, imag} */,
  {32'hbf83a58b, 32'h00000000} /* (13, 26, 12) {real, imag} */,
  {32'hbf240afb, 32'h00000000} /* (13, 26, 11) {real, imag} */,
  {32'h3e2f5e36, 32'h00000000} /* (13, 26, 10) {real, imag} */,
  {32'h3f64c1b2, 32'h00000000} /* (13, 26, 9) {real, imag} */,
  {32'h3fb66f32, 32'h00000000} /* (13, 26, 8) {real, imag} */,
  {32'h3fb8c305, 32'h00000000} /* (13, 26, 7) {real, imag} */,
  {32'h3f947aa9, 32'h00000000} /* (13, 26, 6) {real, imag} */,
  {32'h3f84906f, 32'h00000000} /* (13, 26, 5) {real, imag} */,
  {32'h3f2cce8a, 32'h00000000} /* (13, 26, 4) {real, imag} */,
  {32'h3f3b47e2, 32'h00000000} /* (13, 26, 3) {real, imag} */,
  {32'h3f38bbd3, 32'h00000000} /* (13, 26, 2) {real, imag} */,
  {32'h3f1123f2, 32'h00000000} /* (13, 26, 1) {real, imag} */,
  {32'h3e9daf5b, 32'h00000000} /* (13, 26, 0) {real, imag} */,
  {32'h3f356d23, 32'h00000000} /* (13, 25, 31) {real, imag} */,
  {32'h3f832e2c, 32'h00000000} /* (13, 25, 30) {real, imag} */,
  {32'h3fb1b460, 32'h00000000} /* (13, 25, 29) {real, imag} */,
  {32'h3f80d086, 32'h00000000} /* (13, 25, 28) {real, imag} */,
  {32'h3f672fa3, 32'h00000000} /* (13, 25, 27) {real, imag} */,
  {32'h3f99f006, 32'h00000000} /* (13, 25, 26) {real, imag} */,
  {32'h4000ff2a, 32'h00000000} /* (13, 25, 25) {real, imag} */,
  {32'h3fb61857, 32'h00000000} /* (13, 25, 24) {real, imag} */,
  {32'h3f5f0e36, 32'h00000000} /* (13, 25, 23) {real, imag} */,
  {32'h3f8f90c7, 32'h00000000} /* (13, 25, 22) {real, imag} */,
  {32'h3f4a2436, 32'h00000000} /* (13, 25, 21) {real, imag} */,
  {32'hbf0d0ee1, 32'h00000000} /* (13, 25, 20) {real, imag} */,
  {32'hbf7426ae, 32'h00000000} /* (13, 25, 19) {real, imag} */,
  {32'hbf6ac0c8, 32'h00000000} /* (13, 25, 18) {real, imag} */,
  {32'hbf6a1681, 32'h00000000} /* (13, 25, 17) {real, imag} */,
  {32'hbfabaf18, 32'h00000000} /* (13, 25, 16) {real, imag} */,
  {32'hbf3ad0b3, 32'h00000000} /* (13, 25, 15) {real, imag} */,
  {32'hbf3d4d80, 32'h00000000} /* (13, 25, 14) {real, imag} */,
  {32'hbfe8dc56, 32'h00000000} /* (13, 25, 13) {real, imag} */,
  {32'hbfa7fce0, 32'h00000000} /* (13, 25, 12) {real, imag} */,
  {32'hbf2efd6d, 32'h00000000} /* (13, 25, 11) {real, imag} */,
  {32'h3e9a92b7, 32'h00000000} /* (13, 25, 10) {real, imag} */,
  {32'h3fa5846c, 32'h00000000} /* (13, 25, 9) {real, imag} */,
  {32'h3fb7992b, 32'h00000000} /* (13, 25, 8) {real, imag} */,
  {32'h3f4a4888, 32'h00000000} /* (13, 25, 7) {real, imag} */,
  {32'h3f23832a, 32'h00000000} /* (13, 25, 6) {real, imag} */,
  {32'h3f9830ef, 32'h00000000} /* (13, 25, 5) {real, imag} */,
  {32'h3f6e28d1, 32'h00000000} /* (13, 25, 4) {real, imag} */,
  {32'h3f3c1281, 32'h00000000} /* (13, 25, 3) {real, imag} */,
  {32'h3f2332e0, 32'h00000000} /* (13, 25, 2) {real, imag} */,
  {32'h3f4a33df, 32'h00000000} /* (13, 25, 1) {real, imag} */,
  {32'h3f0c65df, 32'h00000000} /* (13, 25, 0) {real, imag} */,
  {32'h3f15177a, 32'h00000000} /* (13, 24, 31) {real, imag} */,
  {32'h3f1d41c0, 32'h00000000} /* (13, 24, 30) {real, imag} */,
  {32'h3f8b8fb3, 32'h00000000} /* (13, 24, 29) {real, imag} */,
  {32'h3f7fff60, 32'h00000000} /* (13, 24, 28) {real, imag} */,
  {32'h3f23b590, 32'h00000000} /* (13, 24, 27) {real, imag} */,
  {32'h3f72f8aa, 32'h00000000} /* (13, 24, 26) {real, imag} */,
  {32'h3fc08fff, 32'h00000000} /* (13, 24, 25) {real, imag} */,
  {32'h3fd12b35, 32'h00000000} /* (13, 24, 24) {real, imag} */,
  {32'h3f3b3f80, 32'h00000000} /* (13, 24, 23) {real, imag} */,
  {32'h3f8f4de5, 32'h00000000} /* (13, 24, 22) {real, imag} */,
  {32'h3f7fe995, 32'h00000000} /* (13, 24, 21) {real, imag} */,
  {32'hbe5354da, 32'h00000000} /* (13, 24, 20) {real, imag} */,
  {32'hbf12b66d, 32'h00000000} /* (13, 24, 19) {real, imag} */,
  {32'hbf55a303, 32'h00000000} /* (13, 24, 18) {real, imag} */,
  {32'hbf9d1deb, 32'h00000000} /* (13, 24, 17) {real, imag} */,
  {32'hbfd6a491, 32'h00000000} /* (13, 24, 16) {real, imag} */,
  {32'hbf8422cf, 32'h00000000} /* (13, 24, 15) {real, imag} */,
  {32'hbfa7a275, 32'h00000000} /* (13, 24, 14) {real, imag} */,
  {32'hc025eefd, 32'h00000000} /* (13, 24, 13) {real, imag} */,
  {32'hc004b8bb, 32'h00000000} /* (13, 24, 12) {real, imag} */,
  {32'hbfb09b34, 32'h00000000} /* (13, 24, 11) {real, imag} */,
  {32'h3d835014, 32'h00000000} /* (13, 24, 10) {real, imag} */,
  {32'h3faf23b0, 32'h00000000} /* (13, 24, 9) {real, imag} */,
  {32'h3fb47eaa, 32'h00000000} /* (13, 24, 8) {real, imag} */,
  {32'h3f593c79, 32'h00000000} /* (13, 24, 7) {real, imag} */,
  {32'h3eb08ec8, 32'h00000000} /* (13, 24, 6) {real, imag} */,
  {32'h3f2e6638, 32'h00000000} /* (13, 24, 5) {real, imag} */,
  {32'h3f707906, 32'h00000000} /* (13, 24, 4) {real, imag} */,
  {32'h3f1f1b2b, 32'h00000000} /* (13, 24, 3) {real, imag} */,
  {32'h3e99dfd4, 32'h00000000} /* (13, 24, 2) {real, imag} */,
  {32'h3f166487, 32'h00000000} /* (13, 24, 1) {real, imag} */,
  {32'h3f1ea03a, 32'h00000000} /* (13, 24, 0) {real, imag} */,
  {32'h3f06f271, 32'h00000000} /* (13, 23, 31) {real, imag} */,
  {32'h3f8fce8f, 32'h00000000} /* (13, 23, 30) {real, imag} */,
  {32'h3f614ad4, 32'h00000000} /* (13, 23, 29) {real, imag} */,
  {32'h3f5b27d3, 32'h00000000} /* (13, 23, 28) {real, imag} */,
  {32'h3f1088b2, 32'h00000000} /* (13, 23, 27) {real, imag} */,
  {32'h3f5f1343, 32'h00000000} /* (13, 23, 26) {real, imag} */,
  {32'h3f592630, 32'h00000000} /* (13, 23, 25) {real, imag} */,
  {32'h3f84a6e0, 32'h00000000} /* (13, 23, 24) {real, imag} */,
  {32'h3f881b7a, 32'h00000000} /* (13, 23, 23) {real, imag} */,
  {32'h3f81c649, 32'h00000000} /* (13, 23, 22) {real, imag} */,
  {32'h3ef027cb, 32'h00000000} /* (13, 23, 21) {real, imag} */,
  {32'hbf41fe6f, 32'h00000000} /* (13, 23, 20) {real, imag} */,
  {32'hbf1456f9, 32'h00000000} /* (13, 23, 19) {real, imag} */,
  {32'hbf4679ef, 32'h00000000} /* (13, 23, 18) {real, imag} */,
  {32'hbf5e1f32, 32'h00000000} /* (13, 23, 17) {real, imag} */,
  {32'hbf9d1996, 32'h00000000} /* (13, 23, 16) {real, imag} */,
  {32'hbf97ec61, 32'h00000000} /* (13, 23, 15) {real, imag} */,
  {32'hbfb13bcb, 32'h00000000} /* (13, 23, 14) {real, imag} */,
  {32'hbff4b58b, 32'h00000000} /* (13, 23, 13) {real, imag} */,
  {32'hbfdb1ca1, 32'h00000000} /* (13, 23, 12) {real, imag} */,
  {32'hbfa37fb7, 32'h00000000} /* (13, 23, 11) {real, imag} */,
  {32'hbec57669, 32'h00000000} /* (13, 23, 10) {real, imag} */,
  {32'h3f108b79, 32'h00000000} /* (13, 23, 9) {real, imag} */,
  {32'h3f96f82c, 32'h00000000} /* (13, 23, 8) {real, imag} */,
  {32'h3f806f06, 32'h00000000} /* (13, 23, 7) {real, imag} */,
  {32'h3f3e2fc5, 32'h00000000} /* (13, 23, 6) {real, imag} */,
  {32'h3f6335d4, 32'h00000000} /* (13, 23, 5) {real, imag} */,
  {32'h3f54e5e5, 32'h00000000} /* (13, 23, 4) {real, imag} */,
  {32'h3f215824, 32'h00000000} /* (13, 23, 3) {real, imag} */,
  {32'h3f1908fe, 32'h00000000} /* (13, 23, 2) {real, imag} */,
  {32'h3f222c1b, 32'h00000000} /* (13, 23, 1) {real, imag} */,
  {32'h3eec55d0, 32'h00000000} /* (13, 23, 0) {real, imag} */,
  {32'h3f4ceab2, 32'h00000000} /* (13, 22, 31) {real, imag} */,
  {32'h3fb2ac13, 32'h00000000} /* (13, 22, 30) {real, imag} */,
  {32'h3fa5d20f, 32'h00000000} /* (13, 22, 29) {real, imag} */,
  {32'h3f9aa223, 32'h00000000} /* (13, 22, 28) {real, imag} */,
  {32'h3f35ba1f, 32'h00000000} /* (13, 22, 27) {real, imag} */,
  {32'h3f47efe8, 32'h00000000} /* (13, 22, 26) {real, imag} */,
  {32'h3f0269a0, 32'h00000000} /* (13, 22, 25) {real, imag} */,
  {32'h3f5a745a, 32'h00000000} /* (13, 22, 24) {real, imag} */,
  {32'h3f9d433f, 32'h00000000} /* (13, 22, 23) {real, imag} */,
  {32'h3f921343, 32'h00000000} /* (13, 22, 22) {real, imag} */,
  {32'h3ca9a985, 32'h00000000} /* (13, 22, 21) {real, imag} */,
  {32'hbf80a2ea, 32'h00000000} /* (13, 22, 20) {real, imag} */,
  {32'hbf45ce88, 32'h00000000} /* (13, 22, 19) {real, imag} */,
  {32'hbf6fee9e, 32'h00000000} /* (13, 22, 18) {real, imag} */,
  {32'hbf4da88c, 32'h00000000} /* (13, 22, 17) {real, imag} */,
  {32'hbf053c0d, 32'h00000000} /* (13, 22, 16) {real, imag} */,
  {32'hbef4e1e0, 32'h00000000} /* (13, 22, 15) {real, imag} */,
  {32'hbf2b3cdd, 32'h00000000} /* (13, 22, 14) {real, imag} */,
  {32'hbf80a3ef, 32'h00000000} /* (13, 22, 13) {real, imag} */,
  {32'hbfaee06c, 32'h00000000} /* (13, 22, 12) {real, imag} */,
  {32'hbfad0ebb, 32'h00000000} /* (13, 22, 11) {real, imag} */,
  {32'hbedd9ed2, 32'h00000000} /* (13, 22, 10) {real, imag} */,
  {32'h3f5bb7df, 32'h00000000} /* (13, 22, 9) {real, imag} */,
  {32'h3f9856db, 32'h00000000} /* (13, 22, 8) {real, imag} */,
  {32'h3fac7b3c, 32'h00000000} /* (13, 22, 7) {real, imag} */,
  {32'h3f4ae0f3, 32'h00000000} /* (13, 22, 6) {real, imag} */,
  {32'h3f6fcdc3, 32'h00000000} /* (13, 22, 5) {real, imag} */,
  {32'h3f3f1aa8, 32'h00000000} /* (13, 22, 4) {real, imag} */,
  {32'h3f06f8e8, 32'h00000000} /* (13, 22, 3) {real, imag} */,
  {32'h3f8ca5e3, 32'h00000000} /* (13, 22, 2) {real, imag} */,
  {32'h3f4bb03e, 32'h00000000} /* (13, 22, 1) {real, imag} */,
  {32'h3ebadabf, 32'h00000000} /* (13, 22, 0) {real, imag} */,
  {32'h3e92d385, 32'h00000000} /* (13, 21, 31) {real, imag} */,
  {32'h3ea9d753, 32'h00000000} /* (13, 21, 30) {real, imag} */,
  {32'h3ed3225b, 32'h00000000} /* (13, 21, 29) {real, imag} */,
  {32'h3e668b81, 32'h00000000} /* (13, 21, 28) {real, imag} */,
  {32'h3dc403f5, 32'h00000000} /* (13, 21, 27) {real, imag} */,
  {32'hbda26aeb, 32'h00000000} /* (13, 21, 26) {real, imag} */,
  {32'hbe8f0a1b, 32'h00000000} /* (13, 21, 25) {real, imag} */,
  {32'h3f286ce0, 32'h00000000} /* (13, 21, 24) {real, imag} */,
  {32'h3ef728f6, 32'h00000000} /* (13, 21, 23) {real, imag} */,
  {32'h3f171575, 32'h00000000} /* (13, 21, 22) {real, imag} */,
  {32'h3e093770, 32'h00000000} /* (13, 21, 21) {real, imag} */,
  {32'h3de6913c, 32'h00000000} /* (13, 21, 20) {real, imag} */,
  {32'hbe9ea6e4, 32'h00000000} /* (13, 21, 19) {real, imag} */,
  {32'hbea5c61b, 32'h00000000} /* (13, 21, 18) {real, imag} */,
  {32'hbec299c7, 32'h00000000} /* (13, 21, 17) {real, imag} */,
  {32'hbdab9d52, 32'h00000000} /* (13, 21, 16) {real, imag} */,
  {32'h3b835b3a, 32'h00000000} /* (13, 21, 15) {real, imag} */,
  {32'h3cc70523, 32'h00000000} /* (13, 21, 14) {real, imag} */,
  {32'h3cad9c9e, 32'h00000000} /* (13, 21, 13) {real, imag} */,
  {32'hbd5d23ea, 32'h00000000} /* (13, 21, 12) {real, imag} */,
  {32'hbf0b16c1, 32'h00000000} /* (13, 21, 11) {real, imag} */,
  {32'hbe849535, 32'h00000000} /* (13, 21, 10) {real, imag} */,
  {32'h3f9366c5, 32'h00000000} /* (13, 21, 9) {real, imag} */,
  {32'h3fa9a657, 32'h00000000} /* (13, 21, 8) {real, imag} */,
  {32'h3f49c63f, 32'h00000000} /* (13, 21, 7) {real, imag} */,
  {32'hbe6086ab, 32'h00000000} /* (13, 21, 6) {real, imag} */,
  {32'h3e798537, 32'h00000000} /* (13, 21, 5) {real, imag} */,
  {32'h3eedb714, 32'h00000000} /* (13, 21, 4) {real, imag} */,
  {32'h3e951256, 32'h00000000} /* (13, 21, 3) {real, imag} */,
  {32'h3ea9c133, 32'h00000000} /* (13, 21, 2) {real, imag} */,
  {32'h3ea1cc44, 32'h00000000} /* (13, 21, 1) {real, imag} */,
  {32'h3e9e17e2, 32'h00000000} /* (13, 21, 0) {real, imag} */,
  {32'hbedaf1fe, 32'h00000000} /* (13, 20, 31) {real, imag} */,
  {32'hbf3fa8b7, 32'h00000000} /* (13, 20, 30) {real, imag} */,
  {32'hbf7cf6b5, 32'h00000000} /* (13, 20, 29) {real, imag} */,
  {32'hbfb44277, 32'h00000000} /* (13, 20, 28) {real, imag} */,
  {32'hbf8674f2, 32'h00000000} /* (13, 20, 27) {real, imag} */,
  {32'hbf36957d, 32'h00000000} /* (13, 20, 26) {real, imag} */,
  {32'hbf4991e0, 32'h00000000} /* (13, 20, 25) {real, imag} */,
  {32'hbe7a3a3c, 32'h00000000} /* (13, 20, 24) {real, imag} */,
  {32'hbf27cc2c, 32'h00000000} /* (13, 20, 23) {real, imag} */,
  {32'hbf638617, 32'h00000000} /* (13, 20, 22) {real, imag} */,
  {32'hbe9850dc, 32'h00000000} /* (13, 20, 21) {real, imag} */,
  {32'h3f15e5c0, 32'h00000000} /* (13, 20, 20) {real, imag} */,
  {32'h3f473b6c, 32'h00000000} /* (13, 20, 19) {real, imag} */,
  {32'h3f954496, 32'h00000000} /* (13, 20, 18) {real, imag} */,
  {32'h3f7714a4, 32'h00000000} /* (13, 20, 17) {real, imag} */,
  {32'h3f242ad0, 32'h00000000} /* (13, 20, 16) {real, imag} */,
  {32'h3f2fa970, 32'h00000000} /* (13, 20, 15) {real, imag} */,
  {32'h3f687426, 32'h00000000} /* (13, 20, 14) {real, imag} */,
  {32'h3f1f1c69, 32'h00000000} /* (13, 20, 13) {real, imag} */,
  {32'h3f71fad7, 32'h00000000} /* (13, 20, 12) {real, imag} */,
  {32'h3f185706, 32'h00000000} /* (13, 20, 11) {real, imag} */,
  {32'hbf1eccaf, 32'h00000000} /* (13, 20, 10) {real, imag} */,
  {32'hbe436d13, 32'h00000000} /* (13, 20, 9) {real, imag} */,
  {32'hbe949e61, 32'h00000000} /* (13, 20, 8) {real, imag} */,
  {32'hbf5c7dc2, 32'h00000000} /* (13, 20, 7) {real, imag} */,
  {32'hbf8021b7, 32'h00000000} /* (13, 20, 6) {real, imag} */,
  {32'hbf583c0c, 32'h00000000} /* (13, 20, 5) {real, imag} */,
  {32'hbf3ccd84, 32'h00000000} /* (13, 20, 4) {real, imag} */,
  {32'hbf62ef74, 32'h00000000} /* (13, 20, 3) {real, imag} */,
  {32'hbfb53327, 32'h00000000} /* (13, 20, 2) {real, imag} */,
  {32'hbf701460, 32'h00000000} /* (13, 20, 1) {real, imag} */,
  {32'hbf038807, 32'h00000000} /* (13, 20, 0) {real, imag} */,
  {32'hbe748a91, 32'h00000000} /* (13, 19, 31) {real, imag} */,
  {32'hbf4f5546, 32'h00000000} /* (13, 19, 30) {real, imag} */,
  {32'hbf984487, 32'h00000000} /* (13, 19, 29) {real, imag} */,
  {32'hbf8e4a14, 32'h00000000} /* (13, 19, 28) {real, imag} */,
  {32'hbf96553a, 32'h00000000} /* (13, 19, 27) {real, imag} */,
  {32'hbf383058, 32'h00000000} /* (13, 19, 26) {real, imag} */,
  {32'hbef4a701, 32'h00000000} /* (13, 19, 25) {real, imag} */,
  {32'hbf2d548f, 32'h00000000} /* (13, 19, 24) {real, imag} */,
  {32'hbf935ead, 32'h00000000} /* (13, 19, 23) {real, imag} */,
  {32'hbf87cae9, 32'h00000000} /* (13, 19, 22) {real, imag} */,
  {32'hbf074fe2, 32'h00000000} /* (13, 19, 21) {real, imag} */,
  {32'h3f36be49, 32'h00000000} /* (13, 19, 20) {real, imag} */,
  {32'h3fba1e74, 32'h00000000} /* (13, 19, 19) {real, imag} */,
  {32'h3fb28c7c, 32'h00000000} /* (13, 19, 18) {real, imag} */,
  {32'h3f4ebc43, 32'h00000000} /* (13, 19, 17) {real, imag} */,
  {32'h3f64cb20, 32'h00000000} /* (13, 19, 16) {real, imag} */,
  {32'h3f9304d2, 32'h00000000} /* (13, 19, 15) {real, imag} */,
  {32'h3f79b156, 32'h00000000} /* (13, 19, 14) {real, imag} */,
  {32'h3f09d7e5, 32'h00000000} /* (13, 19, 13) {real, imag} */,
  {32'h3f89b6e8, 32'h00000000} /* (13, 19, 12) {real, imag} */,
  {32'h3f77f081, 32'h00000000} /* (13, 19, 11) {real, imag} */,
  {32'hbf0adec4, 32'h00000000} /* (13, 19, 10) {real, imag} */,
  {32'hbf3a0e96, 32'h00000000} /* (13, 19, 9) {real, imag} */,
  {32'hbf426cd2, 32'h00000000} /* (13, 19, 8) {real, imag} */,
  {32'hbfb97f15, 32'h00000000} /* (13, 19, 7) {real, imag} */,
  {32'hbf58b02a, 32'h00000000} /* (13, 19, 6) {real, imag} */,
  {32'hbf513b51, 32'h00000000} /* (13, 19, 5) {real, imag} */,
  {32'hbf361b66, 32'h00000000} /* (13, 19, 4) {real, imag} */,
  {32'hbf575e77, 32'h00000000} /* (13, 19, 3) {real, imag} */,
  {32'hbf921dd4, 32'h00000000} /* (13, 19, 2) {real, imag} */,
  {32'hbf518289, 32'h00000000} /* (13, 19, 1) {real, imag} */,
  {32'hbedb8161, 32'h00000000} /* (13, 19, 0) {real, imag} */,
  {32'hbe4f66c5, 32'h00000000} /* (13, 18, 31) {real, imag} */,
  {32'hbf54c209, 32'h00000000} /* (13, 18, 30) {real, imag} */,
  {32'hbf703dfa, 32'h00000000} /* (13, 18, 29) {real, imag} */,
  {32'hbf18def1, 32'h00000000} /* (13, 18, 28) {real, imag} */,
  {32'hbf3e8ac1, 32'h00000000} /* (13, 18, 27) {real, imag} */,
  {32'hbf3735a4, 32'h00000000} /* (13, 18, 26) {real, imag} */,
  {32'hbef0f398, 32'h00000000} /* (13, 18, 25) {real, imag} */,
  {32'hbfa28b5c, 32'h00000000} /* (13, 18, 24) {real, imag} */,
  {32'hbfc8b815, 32'h00000000} /* (13, 18, 23) {real, imag} */,
  {32'hbf965584, 32'h00000000} /* (13, 18, 22) {real, imag} */,
  {32'hbf37d052, 32'h00000000} /* (13, 18, 21) {real, imag} */,
  {32'h3ecf6c13, 32'h00000000} /* (13, 18, 20) {real, imag} */,
  {32'h3f89afcc, 32'h00000000} /* (13, 18, 19) {real, imag} */,
  {32'h3f3b56b2, 32'h00000000} /* (13, 18, 18) {real, imag} */,
  {32'h3f094b99, 32'h00000000} /* (13, 18, 17) {real, imag} */,
  {32'h3f4828dd, 32'h00000000} /* (13, 18, 16) {real, imag} */,
  {32'h3f2d24ee, 32'h00000000} /* (13, 18, 15) {real, imag} */,
  {32'h3f501410, 32'h00000000} /* (13, 18, 14) {real, imag} */,
  {32'h3f5d309f, 32'h00000000} /* (13, 18, 13) {real, imag} */,
  {32'h3f55d62f, 32'h00000000} /* (13, 18, 12) {real, imag} */,
  {32'h3f8ed520, 32'h00000000} /* (13, 18, 11) {real, imag} */,
  {32'hbe8a9882, 32'h00000000} /* (13, 18, 10) {real, imag} */,
  {32'hbf48b69b, 32'h00000000} /* (13, 18, 9) {real, imag} */,
  {32'hbf6ea297, 32'h00000000} /* (13, 18, 8) {real, imag} */,
  {32'hbf45bc58, 32'h00000000} /* (13, 18, 7) {real, imag} */,
  {32'hbf8d9f58, 32'h00000000} /* (13, 18, 6) {real, imag} */,
  {32'hbfa4b788, 32'h00000000} /* (13, 18, 5) {real, imag} */,
  {32'hbf87328f, 32'h00000000} /* (13, 18, 4) {real, imag} */,
  {32'hbf70b5dd, 32'h00000000} /* (13, 18, 3) {real, imag} */,
  {32'hbf4a87c5, 32'h00000000} /* (13, 18, 2) {real, imag} */,
  {32'hbf3b29ce, 32'h00000000} /* (13, 18, 1) {real, imag} */,
  {32'hbeaf1293, 32'h00000000} /* (13, 18, 0) {real, imag} */,
  {32'hbda1a8c6, 32'h00000000} /* (13, 17, 31) {real, imag} */,
  {32'hbf41e523, 32'h00000000} /* (13, 17, 30) {real, imag} */,
  {32'hbfa34274, 32'h00000000} /* (13, 17, 29) {real, imag} */,
  {32'hbf5321c1, 32'h00000000} /* (13, 17, 28) {real, imag} */,
  {32'hbf7ff09c, 32'h00000000} /* (13, 17, 27) {real, imag} */,
  {32'hbf56e239, 32'h00000000} /* (13, 17, 26) {real, imag} */,
  {32'hbf23b7cd, 32'h00000000} /* (13, 17, 25) {real, imag} */,
  {32'hbfb4f79c, 32'h00000000} /* (13, 17, 24) {real, imag} */,
  {32'hbfe33999, 32'h00000000} /* (13, 17, 23) {real, imag} */,
  {32'hbfdd6042, 32'h00000000} /* (13, 17, 22) {real, imag} */,
  {32'hbea57252, 32'h00000000} /* (13, 17, 21) {real, imag} */,
  {32'h3f0fe49c, 32'h00000000} /* (13, 17, 20) {real, imag} */,
  {32'h3f465331, 32'h00000000} /* (13, 17, 19) {real, imag} */,
  {32'h3eeb51d8, 32'h00000000} /* (13, 17, 18) {real, imag} */,
  {32'h3f1d7468, 32'h00000000} /* (13, 17, 17) {real, imag} */,
  {32'h3f51b668, 32'h00000000} /* (13, 17, 16) {real, imag} */,
  {32'h3f5c22d3, 32'h00000000} /* (13, 17, 15) {real, imag} */,
  {32'h3efef20c, 32'h00000000} /* (13, 17, 14) {real, imag} */,
  {32'h3ef5efe0, 32'h00000000} /* (13, 17, 13) {real, imag} */,
  {32'h3f740c9c, 32'h00000000} /* (13, 17, 12) {real, imag} */,
  {32'h3f37dd14, 32'h00000000} /* (13, 17, 11) {real, imag} */,
  {32'hbea43991, 32'h00000000} /* (13, 17, 10) {real, imag} */,
  {32'hbf593084, 32'h00000000} /* (13, 17, 9) {real, imag} */,
  {32'hbf8981a6, 32'h00000000} /* (13, 17, 8) {real, imag} */,
  {32'hbf652fc2, 32'h00000000} /* (13, 17, 7) {real, imag} */,
  {32'hbfc295bf, 32'h00000000} /* (13, 17, 6) {real, imag} */,
  {32'hbfaa3a89, 32'h00000000} /* (13, 17, 5) {real, imag} */,
  {32'hbfa517e3, 32'h00000000} /* (13, 17, 4) {real, imag} */,
  {32'hbf768a30, 32'h00000000} /* (13, 17, 3) {real, imag} */,
  {32'hbee657cc, 32'h00000000} /* (13, 17, 2) {real, imag} */,
  {32'hbf43a4de, 32'h00000000} /* (13, 17, 1) {real, imag} */,
  {32'hbe988c9a, 32'h00000000} /* (13, 17, 0) {real, imag} */,
  {32'hbe641756, 32'h00000000} /* (13, 16, 31) {real, imag} */,
  {32'hbf1dd32e, 32'h00000000} /* (13, 16, 30) {real, imag} */,
  {32'hbf7a3d87, 32'h00000000} /* (13, 16, 29) {real, imag} */,
  {32'hbf50a3e7, 32'h00000000} /* (13, 16, 28) {real, imag} */,
  {32'hbf8c984a, 32'h00000000} /* (13, 16, 27) {real, imag} */,
  {32'hbf80c56d, 32'h00000000} /* (13, 16, 26) {real, imag} */,
  {32'hbf6b80bb, 32'h00000000} /* (13, 16, 25) {real, imag} */,
  {32'hbfa2f7c8, 32'h00000000} /* (13, 16, 24) {real, imag} */,
  {32'hbfcf5d46, 32'h00000000} /* (13, 16, 23) {real, imag} */,
  {32'hbfed1892, 32'h00000000} /* (13, 16, 22) {real, imag} */,
  {32'hbe3a5771, 32'h00000000} /* (13, 16, 21) {real, imag} */,
  {32'h3f81fd81, 32'h00000000} /* (13, 16, 20) {real, imag} */,
  {32'h3f4864ea, 32'h00000000} /* (13, 16, 19) {real, imag} */,
  {32'h3f54ff96, 32'h00000000} /* (13, 16, 18) {real, imag} */,
  {32'h3fb3561f, 32'h00000000} /* (13, 16, 17) {real, imag} */,
  {32'h3fa5e2d8, 32'h00000000} /* (13, 16, 16) {real, imag} */,
  {32'h3f92fca8, 32'h00000000} /* (13, 16, 15) {real, imag} */,
  {32'h3f25637f, 32'h00000000} /* (13, 16, 14) {real, imag} */,
  {32'h3f37e6e2, 32'h00000000} /* (13, 16, 13) {real, imag} */,
  {32'h3fc278a1, 32'h00000000} /* (13, 16, 12) {real, imag} */,
  {32'h3f8d19c4, 32'h00000000} /* (13, 16, 11) {real, imag} */,
  {32'h3e516f55, 32'h00000000} /* (13, 16, 10) {real, imag} */,
  {32'hbef782a1, 32'h00000000} /* (13, 16, 9) {real, imag} */,
  {32'hbef006af, 32'h00000000} /* (13, 16, 8) {real, imag} */,
  {32'hbf31cac4, 32'h00000000} /* (13, 16, 7) {real, imag} */,
  {32'hbf61d697, 32'h00000000} /* (13, 16, 6) {real, imag} */,
  {32'hbf5597ac, 32'h00000000} /* (13, 16, 5) {real, imag} */,
  {32'hbf3a2e70, 32'h00000000} /* (13, 16, 4) {real, imag} */,
  {32'hbf20cb9c, 32'h00000000} /* (13, 16, 3) {real, imag} */,
  {32'hbeff9a78, 32'h00000000} /* (13, 16, 2) {real, imag} */,
  {32'hbf6bdcb8, 32'h00000000} /* (13, 16, 1) {real, imag} */,
  {32'hbeec08a9, 32'h00000000} /* (13, 16, 0) {real, imag} */,
  {32'hbf01c29d, 32'h00000000} /* (13, 15, 31) {real, imag} */,
  {32'hbf286545, 32'h00000000} /* (13, 15, 30) {real, imag} */,
  {32'hbfa17da4, 32'h00000000} /* (13, 15, 29) {real, imag} */,
  {32'hbfbe610e, 32'h00000000} /* (13, 15, 28) {real, imag} */,
  {32'hbf964e24, 32'h00000000} /* (13, 15, 27) {real, imag} */,
  {32'hbf633122, 32'h00000000} /* (13, 15, 26) {real, imag} */,
  {32'hbf2e1357, 32'h00000000} /* (13, 15, 25) {real, imag} */,
  {32'hbf0813a2, 32'h00000000} /* (13, 15, 24) {real, imag} */,
  {32'hbfb96332, 32'h00000000} /* (13, 15, 23) {real, imag} */,
  {32'hbfaa439c, 32'h00000000} /* (13, 15, 22) {real, imag} */,
  {32'hbecc7271, 32'h00000000} /* (13, 15, 21) {real, imag} */,
  {32'h3f1a869c, 32'h00000000} /* (13, 15, 20) {real, imag} */,
  {32'h3f5a4a92, 32'h00000000} /* (13, 15, 19) {real, imag} */,
  {32'h3f615b28, 32'h00000000} /* (13, 15, 18) {real, imag} */,
  {32'h3f960d9c, 32'h00000000} /* (13, 15, 17) {real, imag} */,
  {32'h3f88c111, 32'h00000000} /* (13, 15, 16) {real, imag} */,
  {32'h3f789c4a, 32'h00000000} /* (13, 15, 15) {real, imag} */,
  {32'h3f2dec1e, 32'h00000000} /* (13, 15, 14) {real, imag} */,
  {32'h3f364362, 32'h00000000} /* (13, 15, 13) {real, imag} */,
  {32'h3f936df4, 32'h00000000} /* (13, 15, 12) {real, imag} */,
  {32'h3f8d0b27, 32'h00000000} /* (13, 15, 11) {real, imag} */,
  {32'h3e4d1e62, 32'h00000000} /* (13, 15, 10) {real, imag} */,
  {32'hbef94fd1, 32'h00000000} /* (13, 15, 9) {real, imag} */,
  {32'hbf26f3b0, 32'h00000000} /* (13, 15, 8) {real, imag} */,
  {32'hbf8b76ca, 32'h00000000} /* (13, 15, 7) {real, imag} */,
  {32'hbf9d06e7, 32'h00000000} /* (13, 15, 6) {real, imag} */,
  {32'hbf09b322, 32'h00000000} /* (13, 15, 5) {real, imag} */,
  {32'hbef94abe, 32'h00000000} /* (13, 15, 4) {real, imag} */,
  {32'hbf08a468, 32'h00000000} /* (13, 15, 3) {real, imag} */,
  {32'hbf74a293, 32'h00000000} /* (13, 15, 2) {real, imag} */,
  {32'hbfd4effb, 32'h00000000} /* (13, 15, 1) {real, imag} */,
  {32'hbfa217d4, 32'h00000000} /* (13, 15, 0) {real, imag} */,
  {32'hbe8a417e, 32'h00000000} /* (13, 14, 31) {real, imag} */,
  {32'hbedc412d, 32'h00000000} /* (13, 14, 30) {real, imag} */,
  {32'hbf6889ba, 32'h00000000} /* (13, 14, 29) {real, imag} */,
  {32'hbf98a0f7, 32'h00000000} /* (13, 14, 28) {real, imag} */,
  {32'hbf850e2c, 32'h00000000} /* (13, 14, 27) {real, imag} */,
  {32'hbed742c4, 32'h00000000} /* (13, 14, 26) {real, imag} */,
  {32'hbe540669, 32'h00000000} /* (13, 14, 25) {real, imag} */,
  {32'hbeaf1c46, 32'h00000000} /* (13, 14, 24) {real, imag} */,
  {32'hbf6562ad, 32'h00000000} /* (13, 14, 23) {real, imag} */,
  {32'hbed6f16f, 32'h00000000} /* (13, 14, 22) {real, imag} */,
  {32'h3e5d2653, 32'h00000000} /* (13, 14, 21) {real, imag} */,
  {32'h3f00c712, 32'h00000000} /* (13, 14, 20) {real, imag} */,
  {32'h3f2f4dbe, 32'h00000000} /* (13, 14, 19) {real, imag} */,
  {32'h3f09ff2b, 32'h00000000} /* (13, 14, 18) {real, imag} */,
  {32'h3f21a724, 32'h00000000} /* (13, 14, 17) {real, imag} */,
  {32'h3f7dd23d, 32'h00000000} /* (13, 14, 16) {real, imag} */,
  {32'h3f7be32d, 32'h00000000} /* (13, 14, 15) {real, imag} */,
  {32'h3f2fbfba, 32'h00000000} /* (13, 14, 14) {real, imag} */,
  {32'h3f20d08f, 32'h00000000} /* (13, 14, 13) {real, imag} */,
  {32'h3f055bf6, 32'h00000000} /* (13, 14, 12) {real, imag} */,
  {32'h3f1f7e5c, 32'h00000000} /* (13, 14, 11) {real, imag} */,
  {32'hbe769e6a, 32'h00000000} /* (13, 14, 10) {real, imag} */,
  {32'hbefdcf57, 32'h00000000} /* (13, 14, 9) {real, imag} */,
  {32'hbf006cd1, 32'h00000000} /* (13, 14, 8) {real, imag} */,
  {32'hbf934bea, 32'h00000000} /* (13, 14, 7) {real, imag} */,
  {32'hbf973392, 32'h00000000} /* (13, 14, 6) {real, imag} */,
  {32'hbf1333f6, 32'h00000000} /* (13, 14, 5) {real, imag} */,
  {32'hbf59570c, 32'h00000000} /* (13, 14, 4) {real, imag} */,
  {32'hbf5bd8c5, 32'h00000000} /* (13, 14, 3) {real, imag} */,
  {32'hbf906275, 32'h00000000} /* (13, 14, 2) {real, imag} */,
  {32'hbfe18328, 32'h00000000} /* (13, 14, 1) {real, imag} */,
  {32'hbfb244ca, 32'h00000000} /* (13, 14, 0) {real, imag} */,
  {32'hbe8b0c98, 32'h00000000} /* (13, 13, 31) {real, imag} */,
  {32'hbf6be3cf, 32'h00000000} /* (13, 13, 30) {real, imag} */,
  {32'hbf78ce95, 32'h00000000} /* (13, 13, 29) {real, imag} */,
  {32'hbf88ad30, 32'h00000000} /* (13, 13, 28) {real, imag} */,
  {32'hbf7c8aa4, 32'h00000000} /* (13, 13, 27) {real, imag} */,
  {32'hbe404044, 32'h00000000} /* (13, 13, 26) {real, imag} */,
  {32'hbeaa6820, 32'h00000000} /* (13, 13, 25) {real, imag} */,
  {32'hbf50ede7, 32'h00000000} /* (13, 13, 24) {real, imag} */,
  {32'hbeea3368, 32'h00000000} /* (13, 13, 23) {real, imag} */,
  {32'hbe96d6b0, 32'h00000000} /* (13, 13, 22) {real, imag} */,
  {32'hbd7e04df, 32'h00000000} /* (13, 13, 21) {real, imag} */,
  {32'h3efbe07e, 32'h00000000} /* (13, 13, 20) {real, imag} */,
  {32'h3f6f7707, 32'h00000000} /* (13, 13, 19) {real, imag} */,
  {32'h3f393c15, 32'h00000000} /* (13, 13, 18) {real, imag} */,
  {32'h3f01e337, 32'h00000000} /* (13, 13, 17) {real, imag} */,
  {32'h3edc73d2, 32'h00000000} /* (13, 13, 16) {real, imag} */,
  {32'h3f76abea, 32'h00000000} /* (13, 13, 15) {real, imag} */,
  {32'h3f6195a2, 32'h00000000} /* (13, 13, 14) {real, imag} */,
  {32'h3ec0c193, 32'h00000000} /* (13, 13, 13) {real, imag} */,
  {32'h3f0491c9, 32'h00000000} /* (13, 13, 12) {real, imag} */,
  {32'h3f44bf68, 32'h00000000} /* (13, 13, 11) {real, imag} */,
  {32'hbe436f6f, 32'h00000000} /* (13, 13, 10) {real, imag} */,
  {32'hbf15f51c, 32'h00000000} /* (13, 13, 9) {real, imag} */,
  {32'hbf209fa9, 32'h00000000} /* (13, 13, 8) {real, imag} */,
  {32'hbfbb8f5e, 32'h00000000} /* (13, 13, 7) {real, imag} */,
  {32'hbf77b832, 32'h00000000} /* (13, 13, 6) {real, imag} */,
  {32'hbf180b8c, 32'h00000000} /* (13, 13, 5) {real, imag} */,
  {32'hbf41a600, 32'h00000000} /* (13, 13, 4) {real, imag} */,
  {32'hbf4fa0e3, 32'h00000000} /* (13, 13, 3) {real, imag} */,
  {32'hbf55b24b, 32'h00000000} /* (13, 13, 2) {real, imag} */,
  {32'hbf802944, 32'h00000000} /* (13, 13, 1) {real, imag} */,
  {32'hbf232256, 32'h00000000} /* (13, 13, 0) {real, imag} */,
  {32'hbf0332b4, 32'h00000000} /* (13, 12, 31) {real, imag} */,
  {32'hbfa9cfb5, 32'h00000000} /* (13, 12, 30) {real, imag} */,
  {32'hbfe43d46, 32'h00000000} /* (13, 12, 29) {real, imag} */,
  {32'hbfd020f2, 32'h00000000} /* (13, 12, 28) {real, imag} */,
  {32'hbf2b8463, 32'h00000000} /* (13, 12, 27) {real, imag} */,
  {32'hbe9b929c, 32'h00000000} /* (13, 12, 26) {real, imag} */,
  {32'hbf041342, 32'h00000000} /* (13, 12, 25) {real, imag} */,
  {32'hbf5770d4, 32'h00000000} /* (13, 12, 24) {real, imag} */,
  {32'hbf0e1ad6, 32'h00000000} /* (13, 12, 23) {real, imag} */,
  {32'hbeee297f, 32'h00000000} /* (13, 12, 22) {real, imag} */,
  {32'hbd823ea8, 32'h00000000} /* (13, 12, 21) {real, imag} */,
  {32'h3f81fbae, 32'h00000000} /* (13, 12, 20) {real, imag} */,
  {32'h3ff04437, 32'h00000000} /* (13, 12, 19) {real, imag} */,
  {32'h3f90e973, 32'h00000000} /* (13, 12, 18) {real, imag} */,
  {32'h3f439963, 32'h00000000} /* (13, 12, 17) {real, imag} */,
  {32'h3f341fee, 32'h00000000} /* (13, 12, 16) {real, imag} */,
  {32'h3f521a1f, 32'h00000000} /* (13, 12, 15) {real, imag} */,
  {32'h3ecb9209, 32'h00000000} /* (13, 12, 14) {real, imag} */,
  {32'h3ea93c06, 32'h00000000} /* (13, 12, 13) {real, imag} */,
  {32'h3f940b6f, 32'h00000000} /* (13, 12, 12) {real, imag} */,
  {32'h3faf72b8, 32'h00000000} /* (13, 12, 11) {real, imag} */,
  {32'hbe28a202, 32'h00000000} /* (13, 12, 10) {real, imag} */,
  {32'hbf4be5cf, 32'h00000000} /* (13, 12, 9) {real, imag} */,
  {32'hbf24b73b, 32'h00000000} /* (13, 12, 8) {real, imag} */,
  {32'hbf9bc805, 32'h00000000} /* (13, 12, 7) {real, imag} */,
  {32'hbf9518b0, 32'h00000000} /* (13, 12, 6) {real, imag} */,
  {32'hbf72771f, 32'h00000000} /* (13, 12, 5) {real, imag} */,
  {32'hbf0eb9d3, 32'h00000000} /* (13, 12, 4) {real, imag} */,
  {32'hbf74fe6f, 32'h00000000} /* (13, 12, 3) {real, imag} */,
  {32'hbf7591a3, 32'h00000000} /* (13, 12, 2) {real, imag} */,
  {32'hbf30ba4c, 32'h00000000} /* (13, 12, 1) {real, imag} */,
  {32'hbe8d4ec8, 32'h00000000} /* (13, 12, 0) {real, imag} */,
  {32'hbe198f72, 32'h00000000} /* (13, 11, 31) {real, imag} */,
  {32'hbee7be3a, 32'h00000000} /* (13, 11, 30) {real, imag} */,
  {32'hbf49ba82, 32'h00000000} /* (13, 11, 29) {real, imag} */,
  {32'hbf942189, 32'h00000000} /* (13, 11, 28) {real, imag} */,
  {32'hbf111352, 32'h00000000} /* (13, 11, 27) {real, imag} */,
  {32'hbf2245eb, 32'h00000000} /* (13, 11, 26) {real, imag} */,
  {32'hbe901623, 32'h00000000} /* (13, 11, 25) {real, imag} */,
  {32'hbf090f43, 32'h00000000} /* (13, 11, 24) {real, imag} */,
  {32'hbf27bdbd, 32'h00000000} /* (13, 11, 23) {real, imag} */,
  {32'hbdbb4785, 32'h00000000} /* (13, 11, 22) {real, imag} */,
  {32'hbdc63dc6, 32'h00000000} /* (13, 11, 21) {real, imag} */,
  {32'h3eb7c349, 32'h00000000} /* (13, 11, 20) {real, imag} */,
  {32'h3f291af0, 32'h00000000} /* (13, 11, 19) {real, imag} */,
  {32'h3f30f4ed, 32'h00000000} /* (13, 11, 18) {real, imag} */,
  {32'h3faf1289, 32'h00000000} /* (13, 11, 17) {real, imag} */,
  {32'h3f4937c4, 32'h00000000} /* (13, 11, 16) {real, imag} */,
  {32'h3e4f0aed, 32'h00000000} /* (13, 11, 15) {real, imag} */,
  {32'h3e9b1f44, 32'h00000000} /* (13, 11, 14) {real, imag} */,
  {32'h3f36c967, 32'h00000000} /* (13, 11, 13) {real, imag} */,
  {32'h3f82cfc6, 32'h00000000} /* (13, 11, 12) {real, imag} */,
  {32'h3f7c8d5d, 32'h00000000} /* (13, 11, 11) {real, imag} */,
  {32'hbece87cb, 32'h00000000} /* (13, 11, 10) {real, imag} */,
  {32'hbf839463, 32'h00000000} /* (13, 11, 9) {real, imag} */,
  {32'hbf37a90f, 32'h00000000} /* (13, 11, 8) {real, imag} */,
  {32'hbf7e0174, 32'h00000000} /* (13, 11, 7) {real, imag} */,
  {32'hbfd2e96f, 32'h00000000} /* (13, 11, 6) {real, imag} */,
  {32'hbf4d4554, 32'h00000000} /* (13, 11, 5) {real, imag} */,
  {32'hbf0de39a, 32'h00000000} /* (13, 11, 4) {real, imag} */,
  {32'hbf35002f, 32'h00000000} /* (13, 11, 3) {real, imag} */,
  {32'hbf04b190, 32'h00000000} /* (13, 11, 2) {real, imag} */,
  {32'hbf0acbf3, 32'h00000000} /* (13, 11, 1) {real, imag} */,
  {32'hbeed8e51, 32'h00000000} /* (13, 11, 0) {real, imag} */,
  {32'h3f810adc, 32'h00000000} /* (13, 10, 31) {real, imag} */,
  {32'h3f8a0770, 32'h00000000} /* (13, 10, 30) {real, imag} */,
  {32'h3f88cfe6, 32'h00000000} /* (13, 10, 29) {real, imag} */,
  {32'h3f93fe82, 32'h00000000} /* (13, 10, 28) {real, imag} */,
  {32'h3f0fde12, 32'h00000000} /* (13, 10, 27) {real, imag} */,
  {32'h3e0ee294, 32'h00000000} /* (13, 10, 26) {real, imag} */,
  {32'h3e81939f, 32'h00000000} /* (13, 10, 25) {real, imag} */,
  {32'h3f0a39f4, 32'h00000000} /* (13, 10, 24) {real, imag} */,
  {32'hbc9e518b, 32'h00000000} /* (13, 10, 23) {real, imag} */,
  {32'h3e52c95c, 32'h00000000} /* (13, 10, 22) {real, imag} */,
  {32'hbef11f27, 32'h00000000} /* (13, 10, 21) {real, imag} */,
  {32'hbf4cff68, 32'h00000000} /* (13, 10, 20) {real, imag} */,
  {32'hbf1bb4a6, 32'h00000000} /* (13, 10, 19) {real, imag} */,
  {32'hbf2b203e, 32'h00000000} /* (13, 10, 18) {real, imag} */,
  {32'h3ec59897, 32'h00000000} /* (13, 10, 17) {real, imag} */,
  {32'hbec33183, 32'h00000000} /* (13, 10, 16) {real, imag} */,
  {32'hbf0675e6, 32'h00000000} /* (13, 10, 15) {real, imag} */,
  {32'hbe824602, 32'h00000000} /* (13, 10, 14) {real, imag} */,
  {32'h3b0a59c0, 32'h00000000} /* (13, 10, 13) {real, imag} */,
  {32'hbedbb007, 32'h00000000} /* (13, 10, 12) {real, imag} */,
  {32'hbf2d31c7, 32'h00000000} /* (13, 10, 11) {real, imag} */,
  {32'hbe27ac26, 32'h00000000} /* (13, 10, 10) {real, imag} */,
  {32'hbe0346bd, 32'h00000000} /* (13, 10, 9) {real, imag} */,
  {32'h3db12552, 32'h00000000} /* (13, 10, 8) {real, imag} */,
  {32'h3e580ec2, 32'h00000000} /* (13, 10, 7) {real, imag} */,
  {32'hbe54590c, 32'h00000000} /* (13, 10, 6) {real, imag} */,
  {32'h3ed25fc6, 32'h00000000} /* (13, 10, 5) {real, imag} */,
  {32'h3ec2b19e, 32'h00000000} /* (13, 10, 4) {real, imag} */,
  {32'h3ef2cefc, 32'h00000000} /* (13, 10, 3) {real, imag} */,
  {32'h3ef99eec, 32'h00000000} /* (13, 10, 2) {real, imag} */,
  {32'h3ef3e70c, 32'h00000000} /* (13, 10, 1) {real, imag} */,
  {32'h3ea292d7, 32'h00000000} /* (13, 10, 0) {real, imag} */,
  {32'h3eeabc8c, 32'h00000000} /* (13, 9, 31) {real, imag} */,
  {32'h3f1a64b8, 32'h00000000} /* (13, 9, 30) {real, imag} */,
  {32'h3f3175a5, 32'h00000000} /* (13, 9, 29) {real, imag} */,
  {32'h3fa9797a, 32'h00000000} /* (13, 9, 28) {real, imag} */,
  {32'h3f97f8c1, 32'h00000000} /* (13, 9, 27) {real, imag} */,
  {32'h3f68d4e2, 32'h00000000} /* (13, 9, 26) {real, imag} */,
  {32'h3f6827d3, 32'h00000000} /* (13, 9, 25) {real, imag} */,
  {32'h3fba4d35, 32'h00000000} /* (13, 9, 24) {real, imag} */,
  {32'h3ee10147, 32'h00000000} /* (13, 9, 23) {real, imag} */,
  {32'h3eca597d, 32'h00000000} /* (13, 9, 22) {real, imag} */,
  {32'h3e8aaf7e, 32'h00000000} /* (13, 9, 21) {real, imag} */,
  {32'hbf38904a, 32'h00000000} /* (13, 9, 20) {real, imag} */,
  {32'hbf2cd18e, 32'h00000000} /* (13, 9, 19) {real, imag} */,
  {32'hbf9d1286, 32'h00000000} /* (13, 9, 18) {real, imag} */,
  {32'hbf83ff4b, 32'h00000000} /* (13, 9, 17) {real, imag} */,
  {32'hbfa7da03, 32'h00000000} /* (13, 9, 16) {real, imag} */,
  {32'hbf6c658f, 32'h00000000} /* (13, 9, 15) {real, imag} */,
  {32'hbfbe969a, 32'h00000000} /* (13, 9, 14) {real, imag} */,
  {32'hbf5de63d, 32'h00000000} /* (13, 9, 13) {real, imag} */,
  {32'hbf5da746, 32'h00000000} /* (13, 9, 12) {real, imag} */,
  {32'hbf690e2d, 32'h00000000} /* (13, 9, 11) {real, imag} */,
  {32'h3eff320a, 32'h00000000} /* (13, 9, 10) {real, imag} */,
  {32'h3f2d466d, 32'h00000000} /* (13, 9, 9) {real, imag} */,
  {32'h3f4aa35d, 32'h00000000} /* (13, 9, 8) {real, imag} */,
  {32'h3f6d5fb2, 32'h00000000} /* (13, 9, 7) {real, imag} */,
  {32'h3efb366f, 32'h00000000} /* (13, 9, 6) {real, imag} */,
  {32'h3f9fbc90, 32'h00000000} /* (13, 9, 5) {real, imag} */,
  {32'h3f752bde, 32'h00000000} /* (13, 9, 4) {real, imag} */,
  {32'h3f4fd308, 32'h00000000} /* (13, 9, 3) {real, imag} */,
  {32'h3f5ad033, 32'h00000000} /* (13, 9, 2) {real, imag} */,
  {32'h3f5a2d8c, 32'h00000000} /* (13, 9, 1) {real, imag} */,
  {32'h3f091df6, 32'h00000000} /* (13, 9, 0) {real, imag} */,
  {32'h3ef87732, 32'h00000000} /* (13, 8, 31) {real, imag} */,
  {32'h3f08ae30, 32'h00000000} /* (13, 8, 30) {real, imag} */,
  {32'h3dedf438, 32'h00000000} /* (13, 8, 29) {real, imag} */,
  {32'h3f33f7b7, 32'h00000000} /* (13, 8, 28) {real, imag} */,
  {32'h3f50f5b9, 32'h00000000} /* (13, 8, 27) {real, imag} */,
  {32'h3f3297f2, 32'h00000000} /* (13, 8, 26) {real, imag} */,
  {32'h3f148ce3, 32'h00000000} /* (13, 8, 25) {real, imag} */,
  {32'h3fb60e81, 32'h00000000} /* (13, 8, 24) {real, imag} */,
  {32'h3f2adad2, 32'h00000000} /* (13, 8, 23) {real, imag} */,
  {32'h3ee2bea6, 32'h00000000} /* (13, 8, 22) {real, imag} */,
  {32'h3e52dd33, 32'h00000000} /* (13, 8, 21) {real, imag} */,
  {32'hbf503ac7, 32'h00000000} /* (13, 8, 20) {real, imag} */,
  {32'hbf803002, 32'h00000000} /* (13, 8, 19) {real, imag} */,
  {32'hbf32ac04, 32'h00000000} /* (13, 8, 18) {real, imag} */,
  {32'hbf367e9f, 32'h00000000} /* (13, 8, 17) {real, imag} */,
  {32'hbf88d5be, 32'h00000000} /* (13, 8, 16) {real, imag} */,
  {32'hbfaaa0bf, 32'h00000000} /* (13, 8, 15) {real, imag} */,
  {32'hbfaa7341, 32'h00000000} /* (13, 8, 14) {real, imag} */,
  {32'hbf30b1db, 32'h00000000} /* (13, 8, 13) {real, imag} */,
  {32'hbf36ec09, 32'h00000000} /* (13, 8, 12) {real, imag} */,
  {32'hbf82845a, 32'h00000000} /* (13, 8, 11) {real, imag} */,
  {32'h3e82bf7f, 32'h00000000} /* (13, 8, 10) {real, imag} */,
  {32'h3f5c326e, 32'h00000000} /* (13, 8, 9) {real, imag} */,
  {32'h3f5b58a3, 32'h00000000} /* (13, 8, 8) {real, imag} */,
  {32'h3fa1704f, 32'h00000000} /* (13, 8, 7) {real, imag} */,
  {32'h3f6581b1, 32'h00000000} /* (13, 8, 6) {real, imag} */,
  {32'h3f8cb1b6, 32'h00000000} /* (13, 8, 5) {real, imag} */,
  {32'h3f48f3c7, 32'h00000000} /* (13, 8, 4) {real, imag} */,
  {32'h3f532131, 32'h00000000} /* (13, 8, 3) {real, imag} */,
  {32'h3f9cfb3f, 32'h00000000} /* (13, 8, 2) {real, imag} */,
  {32'h3f5649a3, 32'h00000000} /* (13, 8, 1) {real, imag} */,
  {32'h3ea9f595, 32'h00000000} /* (13, 8, 0) {real, imag} */,
  {32'h3ea01fd5, 32'h00000000} /* (13, 7, 31) {real, imag} */,
  {32'h3f068b18, 32'h00000000} /* (13, 7, 30) {real, imag} */,
  {32'h3e584c43, 32'h00000000} /* (13, 7, 29) {real, imag} */,
  {32'h3ef19174, 32'h00000000} /* (13, 7, 28) {real, imag} */,
  {32'h3f1af1f5, 32'h00000000} /* (13, 7, 27) {real, imag} */,
  {32'h3f0a2167, 32'h00000000} /* (13, 7, 26) {real, imag} */,
  {32'h3e99fd88, 32'h00000000} /* (13, 7, 25) {real, imag} */,
  {32'h3f812dd1, 32'h00000000} /* (13, 7, 24) {real, imag} */,
  {32'h3f87bb50, 32'h00000000} /* (13, 7, 23) {real, imag} */,
  {32'h3fb018a6, 32'h00000000} /* (13, 7, 22) {real, imag} */,
  {32'h3df1aef2, 32'h00000000} /* (13, 7, 21) {real, imag} */,
  {32'hbfccaab3, 32'h00000000} /* (13, 7, 20) {real, imag} */,
  {32'hbfabdb84, 32'h00000000} /* (13, 7, 19) {real, imag} */,
  {32'hbf5ffacb, 32'h00000000} /* (13, 7, 18) {real, imag} */,
  {32'hbf7420c6, 32'h00000000} /* (13, 7, 17) {real, imag} */,
  {32'hbf41d0f2, 32'h00000000} /* (13, 7, 16) {real, imag} */,
  {32'hbf7d1ef1, 32'h00000000} /* (13, 7, 15) {real, imag} */,
  {32'hbf752b14, 32'h00000000} /* (13, 7, 14) {real, imag} */,
  {32'hbf34d500, 32'h00000000} /* (13, 7, 13) {real, imag} */,
  {32'hbf8d8107, 32'h00000000} /* (13, 7, 12) {real, imag} */,
  {32'hbfafe2b0, 32'h00000000} /* (13, 7, 11) {real, imag} */,
  {32'h3d61d893, 32'h00000000} /* (13, 7, 10) {real, imag} */,
  {32'h3f0daf40, 32'h00000000} /* (13, 7, 9) {real, imag} */,
  {32'h3f4a1719, 32'h00000000} /* (13, 7, 8) {real, imag} */,
  {32'h3fd07086, 32'h00000000} /* (13, 7, 7) {real, imag} */,
  {32'h3f8d64e0, 32'h00000000} /* (13, 7, 6) {real, imag} */,
  {32'h3f50f8ce, 32'h00000000} /* (13, 7, 5) {real, imag} */,
  {32'h3f98efc8, 32'h00000000} /* (13, 7, 4) {real, imag} */,
  {32'h3f6fe390, 32'h00000000} /* (13, 7, 3) {real, imag} */,
  {32'h3f88ed08, 32'h00000000} /* (13, 7, 2) {real, imag} */,
  {32'h3f4f3138, 32'h00000000} /* (13, 7, 1) {real, imag} */,
  {32'h3e45c1c0, 32'h00000000} /* (13, 7, 0) {real, imag} */,
  {32'h3e9b1062, 32'h00000000} /* (13, 6, 31) {real, imag} */,
  {32'h3e9310ed, 32'h00000000} /* (13, 6, 30) {real, imag} */,
  {32'h3edfa874, 32'h00000000} /* (13, 6, 29) {real, imag} */,
  {32'h3f4ef702, 32'h00000000} /* (13, 6, 28) {real, imag} */,
  {32'h3f83f27b, 32'h00000000} /* (13, 6, 27) {real, imag} */,
  {32'h3f1e5e01, 32'h00000000} /* (13, 6, 26) {real, imag} */,
  {32'h3f4aab36, 32'h00000000} /* (13, 6, 25) {real, imag} */,
  {32'h3f27f245, 32'h00000000} /* (13, 6, 24) {real, imag} */,
  {32'h3f474f59, 32'h00000000} /* (13, 6, 23) {real, imag} */,
  {32'h3faea077, 32'h00000000} /* (13, 6, 22) {real, imag} */,
  {32'h3f51a23f, 32'h00000000} /* (13, 6, 21) {real, imag} */,
  {32'hbf434628, 32'h00000000} /* (13, 6, 20) {real, imag} */,
  {32'hbf7b0ef7, 32'h00000000} /* (13, 6, 19) {real, imag} */,
  {32'hbf877f7f, 32'h00000000} /* (13, 6, 18) {real, imag} */,
  {32'hbf57867f, 32'h00000000} /* (13, 6, 17) {real, imag} */,
  {32'hbf2b4fbd, 32'h00000000} /* (13, 6, 16) {real, imag} */,
  {32'hbf089840, 32'h00000000} /* (13, 6, 15) {real, imag} */,
  {32'hbf3e4e0d, 32'h00000000} /* (13, 6, 14) {real, imag} */,
  {32'hbf661421, 32'h00000000} /* (13, 6, 13) {real, imag} */,
  {32'hbf80f42b, 32'h00000000} /* (13, 6, 12) {real, imag} */,
  {32'hbf5f3564, 32'h00000000} /* (13, 6, 11) {real, imag} */,
  {32'hbdafc13b, 32'h00000000} /* (13, 6, 10) {real, imag} */,
  {32'h3ebfe7be, 32'h00000000} /* (13, 6, 9) {real, imag} */,
  {32'h3f337f4c, 32'h00000000} /* (13, 6, 8) {real, imag} */,
  {32'h3f701bef, 32'h00000000} /* (13, 6, 7) {real, imag} */,
  {32'h3f6f088c, 32'h00000000} /* (13, 6, 6) {real, imag} */,
  {32'h3f24710c, 32'h00000000} /* (13, 6, 5) {real, imag} */,
  {32'h3f8b813d, 32'h00000000} /* (13, 6, 4) {real, imag} */,
  {32'h3f41b755, 32'h00000000} /* (13, 6, 3) {real, imag} */,
  {32'h3f27481f, 32'h00000000} /* (13, 6, 2) {real, imag} */,
  {32'h3f39c8c1, 32'h00000000} /* (13, 6, 1) {real, imag} */,
  {32'h3e95f736, 32'h00000000} /* (13, 6, 0) {real, imag} */,
  {32'h3f0837fe, 32'h00000000} /* (13, 5, 31) {real, imag} */,
  {32'h3f565225, 32'h00000000} /* (13, 5, 30) {real, imag} */,
  {32'h3f8464f9, 32'h00000000} /* (13, 5, 29) {real, imag} */,
  {32'h3f6940c1, 32'h00000000} /* (13, 5, 28) {real, imag} */,
  {32'h3f9b40e0, 32'h00000000} /* (13, 5, 27) {real, imag} */,
  {32'h3f3113f9, 32'h00000000} /* (13, 5, 26) {real, imag} */,
  {32'h3f0d242d, 32'h00000000} /* (13, 5, 25) {real, imag} */,
  {32'h3ed36cf0, 32'h00000000} /* (13, 5, 24) {real, imag} */,
  {32'h3f1022e4, 32'h00000000} /* (13, 5, 23) {real, imag} */,
  {32'h3f79ad54, 32'h00000000} /* (13, 5, 22) {real, imag} */,
  {32'h3fac3e9e, 32'h00000000} /* (13, 5, 21) {real, imag} */,
  {32'h3ed04ad6, 32'h00000000} /* (13, 5, 20) {real, imag} */,
  {32'hbd84fbbf, 32'h00000000} /* (13, 5, 19) {real, imag} */,
  {32'h3dbb01b8, 32'h00000000} /* (13, 5, 18) {real, imag} */,
  {32'h3f5c4509, 32'h00000000} /* (13, 5, 17) {real, imag} */,
  {32'h3eabd3ac, 32'h00000000} /* (13, 5, 16) {real, imag} */,
  {32'hbf1d4fd1, 32'h00000000} /* (13, 5, 15) {real, imag} */,
  {32'hbf8c81e5, 32'h00000000} /* (13, 5, 14) {real, imag} */,
  {32'hbf2cf28a, 32'h00000000} /* (13, 5, 13) {real, imag} */,
  {32'hbf47fa31, 32'h00000000} /* (13, 5, 12) {real, imag} */,
  {32'hbf40e5df, 32'h00000000} /* (13, 5, 11) {real, imag} */,
  {32'hbf296f35, 32'h00000000} /* (13, 5, 10) {real, imag} */,
  {32'hbf2d63ee, 32'h00000000} /* (13, 5, 9) {real, imag} */,
  {32'hbf4c1ca9, 32'h00000000} /* (13, 5, 8) {real, imag} */,
  {32'hbf59fbee, 32'h00000000} /* (13, 5, 7) {real, imag} */,
  {32'hbda45722, 32'h00000000} /* (13, 5, 6) {real, imag} */,
  {32'h3f30a136, 32'h00000000} /* (13, 5, 5) {real, imag} */,
  {32'h3f41bf56, 32'h00000000} /* (13, 5, 4) {real, imag} */,
  {32'h3f6add8a, 32'h00000000} /* (13, 5, 3) {real, imag} */,
  {32'h3f4d072b, 32'h00000000} /* (13, 5, 2) {real, imag} */,
  {32'h3f39bd0c, 32'h00000000} /* (13, 5, 1) {real, imag} */,
  {32'h3ecaec1b, 32'h00000000} /* (13, 5, 0) {real, imag} */,
  {32'h3f1e43b6, 32'h00000000} /* (13, 4, 31) {real, imag} */,
  {32'h3f7687c0, 32'h00000000} /* (13, 4, 30) {real, imag} */,
  {32'h3f88ea0e, 32'h00000000} /* (13, 4, 29) {real, imag} */,
  {32'h3f4928f2, 32'h00000000} /* (13, 4, 28) {real, imag} */,
  {32'h3f721bc6, 32'h00000000} /* (13, 4, 27) {real, imag} */,
  {32'h3f2e5625, 32'h00000000} /* (13, 4, 26) {real, imag} */,
  {32'h3f26db21, 32'h00000000} /* (13, 4, 25) {real, imag} */,
  {32'h3f5c1113, 32'h00000000} /* (13, 4, 24) {real, imag} */,
  {32'h3fa5710d, 32'h00000000} /* (13, 4, 23) {real, imag} */,
  {32'h3fe7e28f, 32'h00000000} /* (13, 4, 22) {real, imag} */,
  {32'h400b5878, 32'h00000000} /* (13, 4, 21) {real, imag} */,
  {32'h3fb4010b, 32'h00000000} /* (13, 4, 20) {real, imag} */,
  {32'h3f2aa736, 32'h00000000} /* (13, 4, 19) {real, imag} */,
  {32'h3f8ce921, 32'h00000000} /* (13, 4, 18) {real, imag} */,
  {32'h3fb5aa44, 32'h00000000} /* (13, 4, 17) {real, imag} */,
  {32'h3f836ee4, 32'h00000000} /* (13, 4, 16) {real, imag} */,
  {32'hbecd8e79, 32'h00000000} /* (13, 4, 15) {real, imag} */,
  {32'hbf89b498, 32'h00000000} /* (13, 4, 14) {real, imag} */,
  {32'hbf3e061f, 32'h00000000} /* (13, 4, 13) {real, imag} */,
  {32'hbf4d5560, 32'h00000000} /* (13, 4, 12) {real, imag} */,
  {32'hbf5460ad, 32'h00000000} /* (13, 4, 11) {real, imag} */,
  {32'hbfa2f3d1, 32'h00000000} /* (13, 4, 10) {real, imag} */,
  {32'hbfc2c5c0, 32'h00000000} /* (13, 4, 9) {real, imag} */,
  {32'hbfa39cea, 32'h00000000} /* (13, 4, 8) {real, imag} */,
  {32'hbf8b20a0, 32'h00000000} /* (13, 4, 7) {real, imag} */,
  {32'hbf2d4d25, 32'h00000000} /* (13, 4, 6) {real, imag} */,
  {32'h3ec77183, 32'h00000000} /* (13, 4, 5) {real, imag} */,
  {32'h3f5872ec, 32'h00000000} /* (13, 4, 4) {real, imag} */,
  {32'h3f74e013, 32'h00000000} /* (13, 4, 3) {real, imag} */,
  {32'h3f886e1c, 32'h00000000} /* (13, 4, 2) {real, imag} */,
  {32'h3f48aaf4, 32'h00000000} /* (13, 4, 1) {real, imag} */,
  {32'h3ef70692, 32'h00000000} /* (13, 4, 0) {real, imag} */,
  {32'h3f1a81d6, 32'h00000000} /* (13, 3, 31) {real, imag} */,
  {32'h3f221e59, 32'h00000000} /* (13, 3, 30) {real, imag} */,
  {32'h3f36e332, 32'h00000000} /* (13, 3, 29) {real, imag} */,
  {32'h3f85ecb5, 32'h00000000} /* (13, 3, 28) {real, imag} */,
  {32'h3f9f9aea, 32'h00000000} /* (13, 3, 27) {real, imag} */,
  {32'h3f771ecb, 32'h00000000} /* (13, 3, 26) {real, imag} */,
  {32'h3f81502b, 32'h00000000} /* (13, 3, 25) {real, imag} */,
  {32'h3fe52935, 32'h00000000} /* (13, 3, 24) {real, imag} */,
  {32'h3fa47ec4, 32'h00000000} /* (13, 3, 23) {real, imag} */,
  {32'h3fb596bc, 32'h00000000} /* (13, 3, 22) {real, imag} */,
  {32'h3faf28e6, 32'h00000000} /* (13, 3, 21) {real, imag} */,
  {32'h3f4f59c9, 32'h00000000} /* (13, 3, 20) {real, imag} */,
  {32'h3edd0688, 32'h00000000} /* (13, 3, 19) {real, imag} */,
  {32'h3f63431b, 32'h00000000} /* (13, 3, 18) {real, imag} */,
  {32'h3f621e08, 32'h00000000} /* (13, 3, 17) {real, imag} */,
  {32'h3efdc668, 32'h00000000} /* (13, 3, 16) {real, imag} */,
  {32'hbeea9aa1, 32'h00000000} /* (13, 3, 15) {real, imag} */,
  {32'hbf7095c0, 32'h00000000} /* (13, 3, 14) {real, imag} */,
  {32'hbf6930f9, 32'h00000000} /* (13, 3, 13) {real, imag} */,
  {32'hbf8441d1, 32'h00000000} /* (13, 3, 12) {real, imag} */,
  {32'hbfd6d5a9, 32'h00000000} /* (13, 3, 11) {real, imag} */,
  {32'hbf9ac4db, 32'h00000000} /* (13, 3, 10) {real, imag} */,
  {32'hbfafa0e2, 32'h00000000} /* (13, 3, 9) {real, imag} */,
  {32'hbf70779a, 32'h00000000} /* (13, 3, 8) {real, imag} */,
  {32'hbf12c7a7, 32'h00000000} /* (13, 3, 7) {real, imag} */,
  {32'hbf06a978, 32'h00000000} /* (13, 3, 6) {real, imag} */,
  {32'h3f26303a, 32'h00000000} /* (13, 3, 5) {real, imag} */,
  {32'h3fc13e6a, 32'h00000000} /* (13, 3, 4) {real, imag} */,
  {32'h3f4a5948, 32'h00000000} /* (13, 3, 3) {real, imag} */,
  {32'h3f22b9a4, 32'h00000000} /* (13, 3, 2) {real, imag} */,
  {32'h3f079cec, 32'h00000000} /* (13, 3, 1) {real, imag} */,
  {32'h3f1a0252, 32'h00000000} /* (13, 3, 0) {real, imag} */,
  {32'h3eca33f4, 32'h00000000} /* (13, 2, 31) {real, imag} */,
  {32'h3f49c839, 32'h00000000} /* (13, 2, 30) {real, imag} */,
  {32'h3fa26a5d, 32'h00000000} /* (13, 2, 29) {real, imag} */,
  {32'h3fb1e8fc, 32'h00000000} /* (13, 2, 28) {real, imag} */,
  {32'h3fb19f64, 32'h00000000} /* (13, 2, 27) {real, imag} */,
  {32'h3fbbbc22, 32'h00000000} /* (13, 2, 26) {real, imag} */,
  {32'h3fa383fc, 32'h00000000} /* (13, 2, 25) {real, imag} */,
  {32'h3ff1738b, 32'h00000000} /* (13, 2, 24) {real, imag} */,
  {32'h3f8d15e7, 32'h00000000} /* (13, 2, 23) {real, imag} */,
  {32'h3f24f48b, 32'h00000000} /* (13, 2, 22) {real, imag} */,
  {32'h3f301926, 32'h00000000} /* (13, 2, 21) {real, imag} */,
  {32'h3f31d1a6, 32'h00000000} /* (13, 2, 20) {real, imag} */,
  {32'h3f3d8880, 32'h00000000} /* (13, 2, 19) {real, imag} */,
  {32'h3f1071ad, 32'h00000000} /* (13, 2, 18) {real, imag} */,
  {32'h3f069059, 32'h00000000} /* (13, 2, 17) {real, imag} */,
  {32'h3f4da14f, 32'h00000000} /* (13, 2, 16) {real, imag} */,
  {32'hbe9a9174, 32'h00000000} /* (13, 2, 15) {real, imag} */,
  {32'hbf81580a, 32'h00000000} /* (13, 2, 14) {real, imag} */,
  {32'hbf62a750, 32'h00000000} /* (13, 2, 13) {real, imag} */,
  {32'hbf633ee6, 32'h00000000} /* (13, 2, 12) {real, imag} */,
  {32'hbf735833, 32'h00000000} /* (13, 2, 11) {real, imag} */,
  {32'hbf6b4aec, 32'h00000000} /* (13, 2, 10) {real, imag} */,
  {32'hbf8707a2, 32'h00000000} /* (13, 2, 9) {real, imag} */,
  {32'hbf7de625, 32'h00000000} /* (13, 2, 8) {real, imag} */,
  {32'hbf70dec9, 32'h00000000} /* (13, 2, 7) {real, imag} */,
  {32'hbf165269, 32'h00000000} /* (13, 2, 6) {real, imag} */,
  {32'h3f764f8c, 32'h00000000} /* (13, 2, 5) {real, imag} */,
  {32'h3fbcddf5, 32'h00000000} /* (13, 2, 4) {real, imag} */,
  {32'h3f424a90, 32'h00000000} /* (13, 2, 3) {real, imag} */,
  {32'h3f922cf3, 32'h00000000} /* (13, 2, 2) {real, imag} */,
  {32'h3f493c3c, 32'h00000000} /* (13, 2, 1) {real, imag} */,
  {32'h3ec9daf8, 32'h00000000} /* (13, 2, 0) {real, imag} */,
  {32'h3e6d35a3, 32'h00000000} /* (13, 1, 31) {real, imag} */,
  {32'h3f10101b, 32'h00000000} /* (13, 1, 30) {real, imag} */,
  {32'h3f737ca0, 32'h00000000} /* (13, 1, 29) {real, imag} */,
  {32'h3f73030a, 32'h00000000} /* (13, 1, 28) {real, imag} */,
  {32'h3f8b8aca, 32'h00000000} /* (13, 1, 27) {real, imag} */,
  {32'h3f6e9159, 32'h00000000} /* (13, 1, 26) {real, imag} */,
  {32'h3f217aff, 32'h00000000} /* (13, 1, 25) {real, imag} */,
  {32'h3f665de1, 32'h00000000} /* (13, 1, 24) {real, imag} */,
  {32'h3f7d20d0, 32'h00000000} /* (13, 1, 23) {real, imag} */,
  {32'h3f02d96f, 32'h00000000} /* (13, 1, 22) {real, imag} */,
  {32'h3f303a5f, 32'h00000000} /* (13, 1, 21) {real, imag} */,
  {32'h3f965f14, 32'h00000000} /* (13, 1, 20) {real, imag} */,
  {32'h3f708b62, 32'h00000000} /* (13, 1, 19) {real, imag} */,
  {32'h3f17d3bc, 32'h00000000} /* (13, 1, 18) {real, imag} */,
  {32'h3f51b875, 32'h00000000} /* (13, 1, 17) {real, imag} */,
  {32'h3f64cc8a, 32'h00000000} /* (13, 1, 16) {real, imag} */,
  {32'hbe4b374e, 32'h00000000} /* (13, 1, 15) {real, imag} */,
  {32'hbf40139b, 32'h00000000} /* (13, 1, 14) {real, imag} */,
  {32'hbf7f281d, 32'h00000000} /* (13, 1, 13) {real, imag} */,
  {32'hbf6ae7e4, 32'h00000000} /* (13, 1, 12) {real, imag} */,
  {32'hbf1f896a, 32'h00000000} /* (13, 1, 11) {real, imag} */,
  {32'hbf8fa946, 32'h00000000} /* (13, 1, 10) {real, imag} */,
  {32'hbf76659c, 32'h00000000} /* (13, 1, 9) {real, imag} */,
  {32'hbf7bf6db, 32'h00000000} /* (13, 1, 8) {real, imag} */,
  {32'hbfad9a19, 32'h00000000} /* (13, 1, 7) {real, imag} */,
  {32'hbfa4920e, 32'h00000000} /* (13, 1, 6) {real, imag} */,
  {32'h3f23bce1, 32'h00000000} /* (13, 1, 5) {real, imag} */,
  {32'h3f346f3d, 32'h00000000} /* (13, 1, 4) {real, imag} */,
  {32'h3ef7410e, 32'h00000000} /* (13, 1, 3) {real, imag} */,
  {32'h3f6790d6, 32'h00000000} /* (13, 1, 2) {real, imag} */,
  {32'h3f722418, 32'h00000000} /* (13, 1, 1) {real, imag} */,
  {32'h3f012116, 32'h00000000} /* (13, 1, 0) {real, imag} */,
  {32'h3e0d02a1, 32'h00000000} /* (13, 0, 31) {real, imag} */,
  {32'h3e88a23d, 32'h00000000} /* (13, 0, 30) {real, imag} */,
  {32'h3e9a3e61, 32'h00000000} /* (13, 0, 29) {real, imag} */,
  {32'h3f083e3b, 32'h00000000} /* (13, 0, 28) {real, imag} */,
  {32'h3f57fe0c, 32'h00000000} /* (13, 0, 27) {real, imag} */,
  {32'h3f4b3ebe, 32'h00000000} /* (13, 0, 26) {real, imag} */,
  {32'h3e764bb3, 32'h00000000} /* (13, 0, 25) {real, imag} */,
  {32'h3ec73d18, 32'h00000000} /* (13, 0, 24) {real, imag} */,
  {32'h3f1f4374, 32'h00000000} /* (13, 0, 23) {real, imag} */,
  {32'h3eac56bc, 32'h00000000} /* (13, 0, 22) {real, imag} */,
  {32'h3f0e399c, 32'h00000000} /* (13, 0, 21) {real, imag} */,
  {32'h3f818e0d, 32'h00000000} /* (13, 0, 20) {real, imag} */,
  {32'h3f442131, 32'h00000000} /* (13, 0, 19) {real, imag} */,
  {32'h3f32096e, 32'h00000000} /* (13, 0, 18) {real, imag} */,
  {32'h3f3cb760, 32'h00000000} /* (13, 0, 17) {real, imag} */,
  {32'h3d8f42fc, 32'h00000000} /* (13, 0, 16) {real, imag} */,
  {32'hbec0add7, 32'h00000000} /* (13, 0, 15) {real, imag} */,
  {32'hbee2609f, 32'h00000000} /* (13, 0, 14) {real, imag} */,
  {32'hbeee3ef1, 32'h00000000} /* (13, 0, 13) {real, imag} */,
  {32'hbed15332, 32'h00000000} /* (13, 0, 12) {real, imag} */,
  {32'hbf02fe8c, 32'h00000000} /* (13, 0, 11) {real, imag} */,
  {32'hbf69cd05, 32'h00000000} /* (13, 0, 10) {real, imag} */,
  {32'hbebeebe4, 32'h00000000} /* (13, 0, 9) {real, imag} */,
  {32'hbebefa64, 32'h00000000} /* (13, 0, 8) {real, imag} */,
  {32'hbf207552, 32'h00000000} /* (13, 0, 7) {real, imag} */,
  {32'hbf3e9c57, 32'h00000000} /* (13, 0, 6) {real, imag} */,
  {32'h3e029dc8, 32'h00000000} /* (13, 0, 5) {real, imag} */,
  {32'h3e9e4025, 32'h00000000} /* (13, 0, 4) {real, imag} */,
  {32'h3ede3eda, 32'h00000000} /* (13, 0, 3) {real, imag} */,
  {32'h3e1eede5, 32'h00000000} /* (13, 0, 2) {real, imag} */,
  {32'h3ec63e8b, 32'h00000000} /* (13, 0, 1) {real, imag} */,
  {32'h3f0ac704, 32'h00000000} /* (13, 0, 0) {real, imag} */,
  {32'h3ea3162b, 32'h00000000} /* (12, 31, 31) {real, imag} */,
  {32'h3f323cff, 32'h00000000} /* (12, 31, 30) {real, imag} */,
  {32'h3eda3a13, 32'h00000000} /* (12, 31, 29) {real, imag} */,
  {32'h3ed4970c, 32'h00000000} /* (12, 31, 28) {real, imag} */,
  {32'h3f21dd16, 32'h00000000} /* (12, 31, 27) {real, imag} */,
  {32'h3f806a0c, 32'h00000000} /* (12, 31, 26) {real, imag} */,
  {32'h3eda419c, 32'h00000000} /* (12, 31, 25) {real, imag} */,
  {32'h3ea37ea4, 32'h00000000} /* (12, 31, 24) {real, imag} */,
  {32'h3eeab7fd, 32'h00000000} /* (12, 31, 23) {real, imag} */,
  {32'h3f0d6c02, 32'h00000000} /* (12, 31, 22) {real, imag} */,
  {32'hbc2b979a, 32'h00000000} /* (12, 31, 21) {real, imag} */,
  {32'hbeeec814, 32'h00000000} /* (12, 31, 20) {real, imag} */,
  {32'hbf27bb1d, 32'h00000000} /* (12, 31, 19) {real, imag} */,
  {32'hbed56232, 32'h00000000} /* (12, 31, 18) {real, imag} */,
  {32'hbe66b2d0, 32'h00000000} /* (12, 31, 17) {real, imag} */,
  {32'hbe6a0dca, 32'h00000000} /* (12, 31, 16) {real, imag} */,
  {32'hbecf1e57, 32'h00000000} /* (12, 31, 15) {real, imag} */,
  {32'hbf1258a8, 32'h00000000} /* (12, 31, 14) {real, imag} */,
  {32'hbf0f8ad4, 32'h00000000} /* (12, 31, 13) {real, imag} */,
  {32'hbeb18c5e, 32'h00000000} /* (12, 31, 12) {real, imag} */,
  {32'hbe963b92, 32'h00000000} /* (12, 31, 11) {real, imag} */,
  {32'h3f01c05e, 32'h00000000} /* (12, 31, 10) {real, imag} */,
  {32'h3f1ae7f6, 32'h00000000} /* (12, 31, 9) {real, imag} */,
  {32'h3e4b5f16, 32'h00000000} /* (12, 31, 8) {real, imag} */,
  {32'h3e9c2150, 32'h00000000} /* (12, 31, 7) {real, imag} */,
  {32'h3f2fed6f, 32'h00000000} /* (12, 31, 6) {real, imag} */,
  {32'h3f308438, 32'h00000000} /* (12, 31, 5) {real, imag} */,
  {32'h3f3ea9ca, 32'h00000000} /* (12, 31, 4) {real, imag} */,
  {32'h3f241220, 32'h00000000} /* (12, 31, 3) {real, imag} */,
  {32'h3f597a23, 32'h00000000} /* (12, 31, 2) {real, imag} */,
  {32'h3e176143, 32'h00000000} /* (12, 31, 1) {real, imag} */,
  {32'h3df2ea4e, 32'h00000000} /* (12, 31, 0) {real, imag} */,
  {32'h3f171962, 32'h00000000} /* (12, 30, 31) {real, imag} */,
  {32'h3f8f4dd2, 32'h00000000} /* (12, 30, 30) {real, imag} */,
  {32'h3ede776c, 32'h00000000} /* (12, 30, 29) {real, imag} */,
  {32'h3ee88744, 32'h00000000} /* (12, 30, 28) {real, imag} */,
  {32'h3f37d252, 32'h00000000} /* (12, 30, 27) {real, imag} */,
  {32'h3f4bd095, 32'h00000000} /* (12, 30, 26) {real, imag} */,
  {32'h3f551f4b, 32'h00000000} /* (12, 30, 25) {real, imag} */,
  {32'h3f48fb5e, 32'h00000000} /* (12, 30, 24) {real, imag} */,
  {32'h3f8bb875, 32'h00000000} /* (12, 30, 23) {real, imag} */,
  {32'h3fb4acf2, 32'h00000000} /* (12, 30, 22) {real, imag} */,
  {32'h3e8ad802, 32'h00000000} /* (12, 30, 21) {real, imag} */,
  {32'hbf0fa6b6, 32'h00000000} /* (12, 30, 20) {real, imag} */,
  {32'hbf8acbb2, 32'h00000000} /* (12, 30, 19) {real, imag} */,
  {32'hbf690428, 32'h00000000} /* (12, 30, 18) {real, imag} */,
  {32'hbf221441, 32'h00000000} /* (12, 30, 17) {real, imag} */,
  {32'hbf04558d, 32'h00000000} /* (12, 30, 16) {real, imag} */,
  {32'hbf347524, 32'h00000000} /* (12, 30, 15) {real, imag} */,
  {32'hbf2ff96c, 32'h00000000} /* (12, 30, 14) {real, imag} */,
  {32'hbf1ef311, 32'h00000000} /* (12, 30, 13) {real, imag} */,
  {32'hbee45d86, 32'h00000000} /* (12, 30, 12) {real, imag} */,
  {32'h3cbc1868, 32'h00000000} /* (12, 30, 11) {real, imag} */,
  {32'h3f99241c, 32'h00000000} /* (12, 30, 10) {real, imag} */,
  {32'h3fa4096d, 32'h00000000} /* (12, 30, 9) {real, imag} */,
  {32'h3f565944, 32'h00000000} /* (12, 30, 8) {real, imag} */,
  {32'h3f6333e2, 32'h00000000} /* (12, 30, 7) {real, imag} */,
  {32'h3fa1d7b3, 32'h00000000} /* (12, 30, 6) {real, imag} */,
  {32'h3fa0adbe, 32'h00000000} /* (12, 30, 5) {real, imag} */,
  {32'h3fc36622, 32'h00000000} /* (12, 30, 4) {real, imag} */,
  {32'h3fabbfd6, 32'h00000000} /* (12, 30, 3) {real, imag} */,
  {32'h3f93ad8c, 32'h00000000} /* (12, 30, 2) {real, imag} */,
  {32'h3e991b88, 32'h00000000} /* (12, 30, 1) {real, imag} */,
  {32'h3daee026, 32'h00000000} /* (12, 30, 0) {real, imag} */,
  {32'h3f17d201, 32'h00000000} /* (12, 29, 31) {real, imag} */,
  {32'h3fcb0890, 32'h00000000} /* (12, 29, 30) {real, imag} */,
  {32'h3f66b1a8, 32'h00000000} /* (12, 29, 29) {real, imag} */,
  {32'h3efc1458, 32'h00000000} /* (12, 29, 28) {real, imag} */,
  {32'h3f04aa74, 32'h00000000} /* (12, 29, 27) {real, imag} */,
  {32'h3f44c1e6, 32'h00000000} /* (12, 29, 26) {real, imag} */,
  {32'h3f7c10b4, 32'h00000000} /* (12, 29, 25) {real, imag} */,
  {32'h3f4d3d7a, 32'h00000000} /* (12, 29, 24) {real, imag} */,
  {32'h3fcdce55, 32'h00000000} /* (12, 29, 23) {real, imag} */,
  {32'h3fb958b3, 32'h00000000} /* (12, 29, 22) {real, imag} */,
  {32'h3f00a251, 32'h00000000} /* (12, 29, 21) {real, imag} */,
  {32'hbf1c7286, 32'h00000000} /* (12, 29, 20) {real, imag} */,
  {32'hbf9c39b5, 32'h00000000} /* (12, 29, 19) {real, imag} */,
  {32'hbf84a23a, 32'h00000000} /* (12, 29, 18) {real, imag} */,
  {32'hbf4771de, 32'h00000000} /* (12, 29, 17) {real, imag} */,
  {32'hbf5a49f2, 32'h00000000} /* (12, 29, 16) {real, imag} */,
  {32'hbf37712a, 32'h00000000} /* (12, 29, 15) {real, imag} */,
  {32'hbf48aeb6, 32'h00000000} /* (12, 29, 14) {real, imag} */,
  {32'hbf8de53e, 32'h00000000} /* (12, 29, 13) {real, imag} */,
  {32'hbf1e0e4c, 32'h00000000} /* (12, 29, 12) {real, imag} */,
  {32'hbd265207, 32'h00000000} /* (12, 29, 11) {real, imag} */,
  {32'h3ef8420f, 32'h00000000} /* (12, 29, 10) {real, imag} */,
  {32'h3f4e7dd9, 32'h00000000} /* (12, 29, 9) {real, imag} */,
  {32'h3f4cfd3a, 32'h00000000} /* (12, 29, 8) {real, imag} */,
  {32'h3f9822d8, 32'h00000000} /* (12, 29, 7) {real, imag} */,
  {32'h3fc9ae44, 32'h00000000} /* (12, 29, 6) {real, imag} */,
  {32'h3fa361e1, 32'h00000000} /* (12, 29, 5) {real, imag} */,
  {32'h3f9dd020, 32'h00000000} /* (12, 29, 4) {real, imag} */,
  {32'h3faed201, 32'h00000000} /* (12, 29, 3) {real, imag} */,
  {32'h3f8b4852, 32'h00000000} /* (12, 29, 2) {real, imag} */,
  {32'h3f635ea4, 32'h00000000} /* (12, 29, 1) {real, imag} */,
  {32'h3e805ba3, 32'h00000000} /* (12, 29, 0) {real, imag} */,
  {32'h3eda87eb, 32'h00000000} /* (12, 28, 31) {real, imag} */,
  {32'h3fe371ad, 32'h00000000} /* (12, 28, 30) {real, imag} */,
  {32'h3fd01a43, 32'h00000000} /* (12, 28, 29) {real, imag} */,
  {32'h3f6bdfe0, 32'h00000000} /* (12, 28, 28) {real, imag} */,
  {32'h3f81d363, 32'h00000000} /* (12, 28, 27) {real, imag} */,
  {32'h3fa1fbd6, 32'h00000000} /* (12, 28, 26) {real, imag} */,
  {32'h3f60ded2, 32'h00000000} /* (12, 28, 25) {real, imag} */,
  {32'h3f441de3, 32'h00000000} /* (12, 28, 24) {real, imag} */,
  {32'h3fb9b9f9, 32'h00000000} /* (12, 28, 23) {real, imag} */,
  {32'h3f401f12, 32'h00000000} /* (12, 28, 22) {real, imag} */,
  {32'h3e7b2053, 32'h00000000} /* (12, 28, 21) {real, imag} */,
  {32'hbf71dcf5, 32'h00000000} /* (12, 28, 20) {real, imag} */,
  {32'hbfa90728, 32'h00000000} /* (12, 28, 19) {real, imag} */,
  {32'hbfc0169c, 32'h00000000} /* (12, 28, 18) {real, imag} */,
  {32'hbfa86c96, 32'h00000000} /* (12, 28, 17) {real, imag} */,
  {32'hbf93b3e6, 32'h00000000} /* (12, 28, 16) {real, imag} */,
  {32'hbf624028, 32'h00000000} /* (12, 28, 15) {real, imag} */,
  {32'hbf252dbb, 32'h00000000} /* (12, 28, 14) {real, imag} */,
  {32'hbf866e04, 32'h00000000} /* (12, 28, 13) {real, imag} */,
  {32'hbf8fa0fb, 32'h00000000} /* (12, 28, 12) {real, imag} */,
  {32'hbeb90794, 32'h00000000} /* (12, 28, 11) {real, imag} */,
  {32'hbcafee28, 32'h00000000} /* (12, 28, 10) {real, imag} */,
  {32'h3efbd73a, 32'h00000000} /* (12, 28, 9) {real, imag} */,
  {32'h3f3a2f13, 32'h00000000} /* (12, 28, 8) {real, imag} */,
  {32'h3f648fc0, 32'h00000000} /* (12, 28, 7) {real, imag} */,
  {32'h3fbc7113, 32'h00000000} /* (12, 28, 6) {real, imag} */,
  {32'h3fa02690, 32'h00000000} /* (12, 28, 5) {real, imag} */,
  {32'h3fa558b8, 32'h00000000} /* (12, 28, 4) {real, imag} */,
  {32'h3f3aa139, 32'h00000000} /* (12, 28, 3) {real, imag} */,
  {32'h3f758363, 32'h00000000} /* (12, 28, 2) {real, imag} */,
  {32'h3f8c0fcb, 32'h00000000} /* (12, 28, 1) {real, imag} */,
  {32'h3efb2220, 32'h00000000} /* (12, 28, 0) {real, imag} */,
  {32'h3f39064f, 32'h00000000} /* (12, 27, 31) {real, imag} */,
  {32'h3ffd1800, 32'h00000000} /* (12, 27, 30) {real, imag} */,
  {32'h40014991, 32'h00000000} /* (12, 27, 29) {real, imag} */,
  {32'h3fcd7c5c, 32'h00000000} /* (12, 27, 28) {real, imag} */,
  {32'h3fb292cc, 32'h00000000} /* (12, 27, 27) {real, imag} */,
  {32'h3f80e3fd, 32'h00000000} /* (12, 27, 26) {real, imag} */,
  {32'h3f4575b2, 32'h00000000} /* (12, 27, 25) {real, imag} */,
  {32'h3f2024c1, 32'h00000000} /* (12, 27, 24) {real, imag} */,
  {32'h3f818fae, 32'h00000000} /* (12, 27, 23) {real, imag} */,
  {32'h3f67349d, 32'h00000000} /* (12, 27, 22) {real, imag} */,
  {32'h3e64e54c, 32'h00000000} /* (12, 27, 21) {real, imag} */,
  {32'hbf2f0309, 32'h00000000} /* (12, 27, 20) {real, imag} */,
  {32'hbfaf91a1, 32'h00000000} /* (12, 27, 19) {real, imag} */,
  {32'hbfd892b6, 32'h00000000} /* (12, 27, 18) {real, imag} */,
  {32'hbf9212fe, 32'h00000000} /* (12, 27, 17) {real, imag} */,
  {32'hbf95a5c7, 32'h00000000} /* (12, 27, 16) {real, imag} */,
  {32'hbfd52aad, 32'h00000000} /* (12, 27, 15) {real, imag} */,
  {32'hbf85b1ba, 32'h00000000} /* (12, 27, 14) {real, imag} */,
  {32'hbe810d4b, 32'h00000000} /* (12, 27, 13) {real, imag} */,
  {32'hbf694fca, 32'h00000000} /* (12, 27, 12) {real, imag} */,
  {32'hbf33e1b1, 32'h00000000} /* (12, 27, 11) {real, imag} */,
  {32'hbd2b0f17, 32'h00000000} /* (12, 27, 10) {real, imag} */,
  {32'h3f31bfcc, 32'h00000000} /* (12, 27, 9) {real, imag} */,
  {32'h3f87b462, 32'h00000000} /* (12, 27, 8) {real, imag} */,
  {32'h3f51eb96, 32'h00000000} /* (12, 27, 7) {real, imag} */,
  {32'h3fb84c2e, 32'h00000000} /* (12, 27, 6) {real, imag} */,
  {32'h3f81b0db, 32'h00000000} /* (12, 27, 5) {real, imag} */,
  {32'h3f45833c, 32'h00000000} /* (12, 27, 4) {real, imag} */,
  {32'h3f2b7b95, 32'h00000000} /* (12, 27, 3) {real, imag} */,
  {32'h3f2b32af, 32'h00000000} /* (12, 27, 2) {real, imag} */,
  {32'h3f9273bf, 32'h00000000} /* (12, 27, 1) {real, imag} */,
  {32'h3f72e13d, 32'h00000000} /* (12, 27, 0) {real, imag} */,
  {32'h3f27edb1, 32'h00000000} /* (12, 26, 31) {real, imag} */,
  {32'h3fad25c7, 32'h00000000} /* (12, 26, 30) {real, imag} */,
  {32'h3facd938, 32'h00000000} /* (12, 26, 29) {real, imag} */,
  {32'h3f92fbab, 32'h00000000} /* (12, 26, 28) {real, imag} */,
  {32'h3f919f13, 32'h00000000} /* (12, 26, 27) {real, imag} */,
  {32'h3f88c8a4, 32'h00000000} /* (12, 26, 26) {real, imag} */,
  {32'h3fc7730f, 32'h00000000} /* (12, 26, 25) {real, imag} */,
  {32'h3f49acc9, 32'h00000000} /* (12, 26, 24) {real, imag} */,
  {32'h3f404eb9, 32'h00000000} /* (12, 26, 23) {real, imag} */,
  {32'h3f86441f, 32'h00000000} /* (12, 26, 22) {real, imag} */,
  {32'h3e962a8c, 32'h00000000} /* (12, 26, 21) {real, imag} */,
  {32'hbef1c486, 32'h00000000} /* (12, 26, 20) {real, imag} */,
  {32'hbf5c0436, 32'h00000000} /* (12, 26, 19) {real, imag} */,
  {32'hbf63c2c4, 32'h00000000} /* (12, 26, 18) {real, imag} */,
  {32'hbf402108, 32'h00000000} /* (12, 26, 17) {real, imag} */,
  {32'hbfa47678, 32'h00000000} /* (12, 26, 16) {real, imag} */,
  {32'hbfbd2f84, 32'h00000000} /* (12, 26, 15) {real, imag} */,
  {32'hbf8e7913, 32'h00000000} /* (12, 26, 14) {real, imag} */,
  {32'hbf011549, 32'h00000000} /* (12, 26, 13) {real, imag} */,
  {32'hbf20dd84, 32'h00000000} /* (12, 26, 12) {real, imag} */,
  {32'hbf3f20b3, 32'h00000000} /* (12, 26, 11) {real, imag} */,
  {32'h3e233775, 32'h00000000} /* (12, 26, 10) {real, imag} */,
  {32'h3fb2353e, 32'h00000000} /* (12, 26, 9) {real, imag} */,
  {32'h3fc71ea1, 32'h00000000} /* (12, 26, 8) {real, imag} */,
  {32'h3f2a921b, 32'h00000000} /* (12, 26, 7) {real, imag} */,
  {32'h3f041fa3, 32'h00000000} /* (12, 26, 6) {real, imag} */,
  {32'h3ec37d3b, 32'h00000000} /* (12, 26, 5) {real, imag} */,
  {32'h3f023220, 32'h00000000} /* (12, 26, 4) {real, imag} */,
  {32'h3f435dd7, 32'h00000000} /* (12, 26, 3) {real, imag} */,
  {32'h3f5a3df9, 32'h00000000} /* (12, 26, 2) {real, imag} */,
  {32'h3f8f4728, 32'h00000000} /* (12, 26, 1) {real, imag} */,
  {32'h3f4d28fa, 32'h00000000} /* (12, 26, 0) {real, imag} */,
  {32'h3f00ed10, 32'h00000000} /* (12, 25, 31) {real, imag} */,
  {32'h3f72fab0, 32'h00000000} /* (12, 25, 30) {real, imag} */,
  {32'h3f8cb579, 32'h00000000} /* (12, 25, 29) {real, imag} */,
  {32'h3f9ef82f, 32'h00000000} /* (12, 25, 28) {real, imag} */,
  {32'h3f80d87f, 32'h00000000} /* (12, 25, 27) {real, imag} */,
  {32'h3f5df67c, 32'h00000000} /* (12, 25, 26) {real, imag} */,
  {32'h40030b23, 32'h00000000} /* (12, 25, 25) {real, imag} */,
  {32'h3fa9a442, 32'h00000000} /* (12, 25, 24) {real, imag} */,
  {32'h3ec06f7b, 32'h00000000} /* (12, 25, 23) {real, imag} */,
  {32'h3f6da33a, 32'h00000000} /* (12, 25, 22) {real, imag} */,
  {32'h3efbd29d, 32'h00000000} /* (12, 25, 21) {real, imag} */,
  {32'hbf3c4ade, 32'h00000000} /* (12, 25, 20) {real, imag} */,
  {32'hbf2de8ab, 32'h00000000} /* (12, 25, 19) {real, imag} */,
  {32'hbf5fa8ea, 32'h00000000} /* (12, 25, 18) {real, imag} */,
  {32'hbfc01ace, 32'h00000000} /* (12, 25, 17) {real, imag} */,
  {32'hbfe16e29, 32'h00000000} /* (12, 25, 16) {real, imag} */,
  {32'hbf54208c, 32'h00000000} /* (12, 25, 15) {real, imag} */,
  {32'hbe88a74c, 32'h00000000} /* (12, 25, 14) {real, imag} */,
  {32'hbf426d73, 32'h00000000} /* (12, 25, 13) {real, imag} */,
  {32'hbf5a89f8, 32'h00000000} /* (12, 25, 12) {real, imag} */,
  {32'hbf7e8907, 32'h00000000} /* (12, 25, 11) {real, imag} */,
  {32'h3d931f35, 32'h00000000} /* (12, 25, 10) {real, imag} */,
  {32'h3faf8e23, 32'h00000000} /* (12, 25, 9) {real, imag} */,
  {32'h3fa4b778, 32'h00000000} /* (12, 25, 8) {real, imag} */,
  {32'h3eed21df, 32'h00000000} /* (12, 25, 7) {real, imag} */,
  {32'h3ea450fe, 32'h00000000} /* (12, 25, 6) {real, imag} */,
  {32'h3ee1aca6, 32'h00000000} /* (12, 25, 5) {real, imag} */,
  {32'h3f250026, 32'h00000000} /* (12, 25, 4) {real, imag} */,
  {32'h3f3bf71f, 32'h00000000} /* (12, 25, 3) {real, imag} */,
  {32'h3f9ed8ab, 32'h00000000} /* (12, 25, 2) {real, imag} */,
  {32'h3f849b73, 32'h00000000} /* (12, 25, 1) {real, imag} */,
  {32'h3f084b07, 32'h00000000} /* (12, 25, 0) {real, imag} */,
  {32'h3e9aeb31, 32'h00000000} /* (12, 24, 31) {real, imag} */,
  {32'h3f2a3d47, 32'h00000000} /* (12, 24, 30) {real, imag} */,
  {32'h3f965221, 32'h00000000} /* (12, 24, 29) {real, imag} */,
  {32'h3f8f8a09, 32'h00000000} /* (12, 24, 28) {real, imag} */,
  {32'h3f70571f, 32'h00000000} /* (12, 24, 27) {real, imag} */,
  {32'h3f8ab6a3, 32'h00000000} /* (12, 24, 26) {real, imag} */,
  {32'h3fd9ea11, 32'h00000000} /* (12, 24, 25) {real, imag} */,
  {32'h3f9b6361, 32'h00000000} /* (12, 24, 24) {real, imag} */,
  {32'h3e659844, 32'h00000000} /* (12, 24, 23) {real, imag} */,
  {32'h3f42e9e7, 32'h00000000} /* (12, 24, 22) {real, imag} */,
  {32'h3ecd8be1, 32'h00000000} /* (12, 24, 21) {real, imag} */,
  {32'hbf70cafe, 32'h00000000} /* (12, 24, 20) {real, imag} */,
  {32'hbf33e409, 32'h00000000} /* (12, 24, 19) {real, imag} */,
  {32'hbf3b941a, 32'h00000000} /* (12, 24, 18) {real, imag} */,
  {32'hbfb90bc9, 32'h00000000} /* (12, 24, 17) {real, imag} */,
  {32'hbfbc2365, 32'h00000000} /* (12, 24, 16) {real, imag} */,
  {32'hbf59cca3, 32'h00000000} /* (12, 24, 15) {real, imag} */,
  {32'hbf130a24, 32'h00000000} /* (12, 24, 14) {real, imag} */,
  {32'hbf727156, 32'h00000000} /* (12, 24, 13) {real, imag} */,
  {32'hbf8d1490, 32'h00000000} /* (12, 24, 12) {real, imag} */,
  {32'hbf9b20c5, 32'h00000000} /* (12, 24, 11) {real, imag} */,
  {32'hbd8c07ba, 32'h00000000} /* (12, 24, 10) {real, imag} */,
  {32'h3fb0ed75, 32'h00000000} /* (12, 24, 9) {real, imag} */,
  {32'h3f8289b8, 32'h00000000} /* (12, 24, 8) {real, imag} */,
  {32'h3f48d1b8, 32'h00000000} /* (12, 24, 7) {real, imag} */,
  {32'h3f0f26de, 32'h00000000} /* (12, 24, 6) {real, imag} */,
  {32'h3f1d31f9, 32'h00000000} /* (12, 24, 5) {real, imag} */,
  {32'h3f49b2c2, 32'h00000000} /* (12, 24, 4) {real, imag} */,
  {32'h3f27a564, 32'h00000000} /* (12, 24, 3) {real, imag} */,
  {32'h3f576559, 32'h00000000} /* (12, 24, 2) {real, imag} */,
  {32'h3f3c45b7, 32'h00000000} /* (12, 24, 1) {real, imag} */,
  {32'h3eff4258, 32'h00000000} /* (12, 24, 0) {real, imag} */,
  {32'h3eba6f5d, 32'h00000000} /* (12, 23, 31) {real, imag} */,
  {32'h3fb11c18, 32'h00000000} /* (12, 23, 30) {real, imag} */,
  {32'h3fb0fb9d, 32'h00000000} /* (12, 23, 29) {real, imag} */,
  {32'h3f682b8b, 32'h00000000} /* (12, 23, 28) {real, imag} */,
  {32'h3f78e64c, 32'h00000000} /* (12, 23, 27) {real, imag} */,
  {32'h3f802cbe, 32'h00000000} /* (12, 23, 26) {real, imag} */,
  {32'h3f6b171b, 32'h00000000} /* (12, 23, 25) {real, imag} */,
  {32'h3f5ca21c, 32'h00000000} /* (12, 23, 24) {real, imag} */,
  {32'h3f9a2200, 32'h00000000} /* (12, 23, 23) {real, imag} */,
  {32'h3f64b4cf, 32'h00000000} /* (12, 23, 22) {real, imag} */,
  {32'h3e3bcfde, 32'h00000000} /* (12, 23, 21) {real, imag} */,
  {32'hbf4238b0, 32'h00000000} /* (12, 23, 20) {real, imag} */,
  {32'hbf5d37e4, 32'h00000000} /* (12, 23, 19) {real, imag} */,
  {32'hbf849351, 32'h00000000} /* (12, 23, 18) {real, imag} */,
  {32'hbf56cd53, 32'h00000000} /* (12, 23, 17) {real, imag} */,
  {32'hbf685d2c, 32'h00000000} /* (12, 23, 16) {real, imag} */,
  {32'hbf43bfeb, 32'h00000000} /* (12, 23, 15) {real, imag} */,
  {32'hbf85a300, 32'h00000000} /* (12, 23, 14) {real, imag} */,
  {32'hbf86e3c1, 32'h00000000} /* (12, 23, 13) {real, imag} */,
  {32'hbf89d8b2, 32'h00000000} /* (12, 23, 12) {real, imag} */,
  {32'hbf9c962e, 32'h00000000} /* (12, 23, 11) {real, imag} */,
  {32'hbeca01f8, 32'h00000000} /* (12, 23, 10) {real, imag} */,
  {32'h3f24acb5, 32'h00000000} /* (12, 23, 9) {real, imag} */,
  {32'h3f0bf563, 32'h00000000} /* (12, 23, 8) {real, imag} */,
  {32'h3f1ad963, 32'h00000000} /* (12, 23, 7) {real, imag} */,
  {32'h3f1df4d0, 32'h00000000} /* (12, 23, 6) {real, imag} */,
  {32'h3f2af868, 32'h00000000} /* (12, 23, 5) {real, imag} */,
  {32'h3f6da995, 32'h00000000} /* (12, 23, 4) {real, imag} */,
  {32'h3f340757, 32'h00000000} /* (12, 23, 3) {real, imag} */,
  {32'h3f11ef03, 32'h00000000} /* (12, 23, 2) {real, imag} */,
  {32'h3f3692de, 32'h00000000} /* (12, 23, 1) {real, imag} */,
  {32'h3eaf5d4b, 32'h00000000} /* (12, 23, 0) {real, imag} */,
  {32'h3f207b1c, 32'h00000000} /* (12, 22, 31) {real, imag} */,
  {32'h3fbf5566, 32'h00000000} /* (12, 22, 30) {real, imag} */,
  {32'h3f94bd8b, 32'h00000000} /* (12, 22, 29) {real, imag} */,
  {32'h3f6df733, 32'h00000000} /* (12, 22, 28) {real, imag} */,
  {32'h3f2e63ba, 32'h00000000} /* (12, 22, 27) {real, imag} */,
  {32'h3f440330, 32'h00000000} /* (12, 22, 26) {real, imag} */,
  {32'h3f2e1a06, 32'h00000000} /* (12, 22, 25) {real, imag} */,
  {32'h3f4bdf39, 32'h00000000} /* (12, 22, 24) {real, imag} */,
  {32'h3fd5cc08, 32'h00000000} /* (12, 22, 23) {real, imag} */,
  {32'h3facf316, 32'h00000000} /* (12, 22, 22) {real, imag} */,
  {32'hbdfccf80, 32'h00000000} /* (12, 22, 21) {real, imag} */,
  {32'hbf8b0cff, 32'h00000000} /* (12, 22, 20) {real, imag} */,
  {32'hbf569797, 32'h00000000} /* (12, 22, 19) {real, imag} */,
  {32'hbf912277, 32'h00000000} /* (12, 22, 18) {real, imag} */,
  {32'hbf93f794, 32'h00000000} /* (12, 22, 17) {real, imag} */,
  {32'hbf7754ed, 32'h00000000} /* (12, 22, 16) {real, imag} */,
  {32'hbec83074, 32'h00000000} /* (12, 22, 15) {real, imag} */,
  {32'hbf408465, 32'h00000000} /* (12, 22, 14) {real, imag} */,
  {32'hbf939e71, 32'h00000000} /* (12, 22, 13) {real, imag} */,
  {32'hc0013616, 32'h00000000} /* (12, 22, 12) {real, imag} */,
  {32'hbfe4bb6c, 32'h00000000} /* (12, 22, 11) {real, imag} */,
  {32'hbe58dba2, 32'h00000000} /* (12, 22, 10) {real, imag} */,
  {32'h3f9d0fe7, 32'h00000000} /* (12, 22, 9) {real, imag} */,
  {32'h3f7cd6ca, 32'h00000000} /* (12, 22, 8) {real, imag} */,
  {32'h3f72e19e, 32'h00000000} /* (12, 22, 7) {real, imag} */,
  {32'h3f046836, 32'h00000000} /* (12, 22, 6) {real, imag} */,
  {32'h3efcc9c0, 32'h00000000} /* (12, 22, 5) {real, imag} */,
  {32'h3f482af9, 32'h00000000} /* (12, 22, 4) {real, imag} */,
  {32'h3f556b18, 32'h00000000} /* (12, 22, 3) {real, imag} */,
  {32'h3f9da969, 32'h00000000} /* (12, 22, 2) {real, imag} */,
  {32'h3f9c501b, 32'h00000000} /* (12, 22, 1) {real, imag} */,
  {32'h3f040648, 32'h00000000} /* (12, 22, 0) {real, imag} */,
  {32'h3e6038b7, 32'h00000000} /* (12, 21, 31) {real, imag} */,
  {32'h3e85d00b, 32'h00000000} /* (12, 21, 30) {real, imag} */,
  {32'h3ea646f6, 32'h00000000} /* (12, 21, 29) {real, imag} */,
  {32'h3f234256, 32'h00000000} /* (12, 21, 28) {real, imag} */,
  {32'h3e12396f, 32'h00000000} /* (12, 21, 27) {real, imag} */,
  {32'h3e629b91, 32'h00000000} /* (12, 21, 26) {real, imag} */,
  {32'h3e81da44, 32'h00000000} /* (12, 21, 25) {real, imag} */,
  {32'h3ef13c5b, 32'h00000000} /* (12, 21, 24) {real, imag} */,
  {32'h3e89899c, 32'h00000000} /* (12, 21, 23) {real, imag} */,
  {32'h3eb31e72, 32'h00000000} /* (12, 21, 22) {real, imag} */,
  {32'hbdf136bf, 32'h00000000} /* (12, 21, 21) {real, imag} */,
  {32'hbf33932f, 32'h00000000} /* (12, 21, 20) {real, imag} */,
  {32'hbf1c0a62, 32'h00000000} /* (12, 21, 19) {real, imag} */,
  {32'hbe76c6e5, 32'h00000000} /* (12, 21, 18) {real, imag} */,
  {32'hbf09bff0, 32'h00000000} /* (12, 21, 17) {real, imag} */,
  {32'hbee30508, 32'h00000000} /* (12, 21, 16) {real, imag} */,
  {32'hbd921006, 32'h00000000} /* (12, 21, 15) {real, imag} */,
  {32'hbe88403d, 32'h00000000} /* (12, 21, 14) {real, imag} */,
  {32'hbf1b942a, 32'h00000000} /* (12, 21, 13) {real, imag} */,
  {32'hbf288544, 32'h00000000} /* (12, 21, 12) {real, imag} */,
  {32'hbf23437a, 32'h00000000} /* (12, 21, 11) {real, imag} */,
  {32'h3e77e851, 32'h00000000} /* (12, 21, 10) {real, imag} */,
  {32'h3f32f850, 32'h00000000} /* (12, 21, 9) {real, imag} */,
  {32'h3f3faf78, 32'h00000000} /* (12, 21, 8) {real, imag} */,
  {32'h3f0aca0e, 32'h00000000} /* (12, 21, 7) {real, imag} */,
  {32'h3d9a75a6, 32'h00000000} /* (12, 21, 6) {real, imag} */,
  {32'h3dcc957c, 32'h00000000} /* (12, 21, 5) {real, imag} */,
  {32'h3ec75759, 32'h00000000} /* (12, 21, 4) {real, imag} */,
  {32'h3efa1495, 32'h00000000} /* (12, 21, 3) {real, imag} */,
  {32'h3f527711, 32'h00000000} /* (12, 21, 2) {real, imag} */,
  {32'h3f0dd0f0, 32'h00000000} /* (12, 21, 1) {real, imag} */,
  {32'h3d9dff09, 32'h00000000} /* (12, 21, 0) {real, imag} */,
  {32'hbf0a9382, 32'h00000000} /* (12, 20, 31) {real, imag} */,
  {32'hbfadf7f4, 32'h00000000} /* (12, 20, 30) {real, imag} */,
  {32'hbf76f9c6, 32'h00000000} /* (12, 20, 29) {real, imag} */,
  {32'hbf416cf3, 32'h00000000} /* (12, 20, 28) {real, imag} */,
  {32'hbee48ead, 32'h00000000} /* (12, 20, 27) {real, imag} */,
  {32'hbe812402, 32'h00000000} /* (12, 20, 26) {real, imag} */,
  {32'hbf1a1879, 32'h00000000} /* (12, 20, 25) {real, imag} */,
  {32'hbf1ff467, 32'h00000000} /* (12, 20, 24) {real, imag} */,
  {32'hbf9bb991, 32'h00000000} /* (12, 20, 23) {real, imag} */,
  {32'hbfcbeb35, 32'h00000000} /* (12, 20, 22) {real, imag} */,
  {32'hbf0d08a6, 32'h00000000} /* (12, 20, 21) {real, imag} */,
  {32'h3e5095fe, 32'h00000000} /* (12, 20, 20) {real, imag} */,
  {32'h3eff7dc4, 32'h00000000} /* (12, 20, 19) {real, imag} */,
  {32'h3f788d55, 32'h00000000} /* (12, 20, 18) {real, imag} */,
  {32'h3f8a581c, 32'h00000000} /* (12, 20, 17) {real, imag} */,
  {32'h3f06be6e, 32'h00000000} /* (12, 20, 16) {real, imag} */,
  {32'h3f41cb84, 32'h00000000} /* (12, 20, 15) {real, imag} */,
  {32'h3f089876, 32'h00000000} /* (12, 20, 14) {real, imag} */,
  {32'h3ea8ee4f, 32'h00000000} /* (12, 20, 13) {real, imag} */,
  {32'h3f597097, 32'h00000000} /* (12, 20, 12) {real, imag} */,
  {32'h3ee50d97, 32'h00000000} /* (12, 20, 11) {real, imag} */,
  {32'hbf0f8fb3, 32'h00000000} /* (12, 20, 10) {real, imag} */,
  {32'hbf84b0e9, 32'h00000000} /* (12, 20, 9) {real, imag} */,
  {32'hbeedfcb4, 32'h00000000} /* (12, 20, 8) {real, imag} */,
  {32'hbf25f25d, 32'h00000000} /* (12, 20, 7) {real, imag} */,
  {32'hbf3b0f9e, 32'h00000000} /* (12, 20, 6) {real, imag} */,
  {32'hbf7a8741, 32'h00000000} /* (12, 20, 5) {real, imag} */,
  {32'hbf2e020e, 32'h00000000} /* (12, 20, 4) {real, imag} */,
  {32'hbf11723a, 32'h00000000} /* (12, 20, 3) {real, imag} */,
  {32'hbf287a4c, 32'h00000000} /* (12, 20, 2) {real, imag} */,
  {32'hbf3f0c20, 32'h00000000} /* (12, 20, 1) {real, imag} */,
  {32'hbf0142e3, 32'h00000000} /* (12, 20, 0) {real, imag} */,
  {32'hbea26468, 32'h00000000} /* (12, 19, 31) {real, imag} */,
  {32'hbfa134ee, 32'h00000000} /* (12, 19, 30) {real, imag} */,
  {32'hbf7e8457, 32'h00000000} /* (12, 19, 29) {real, imag} */,
  {32'hbf351e35, 32'h00000000} /* (12, 19, 28) {real, imag} */,
  {32'hbf184238, 32'h00000000} /* (12, 19, 27) {real, imag} */,
  {32'hbf54b1dd, 32'h00000000} /* (12, 19, 26) {real, imag} */,
  {32'hbf3e46d7, 32'h00000000} /* (12, 19, 25) {real, imag} */,
  {32'hbf3e6c07, 32'h00000000} /* (12, 19, 24) {real, imag} */,
  {32'hbf914c30, 32'h00000000} /* (12, 19, 23) {real, imag} */,
  {32'hbfa0d0d0, 32'h00000000} /* (12, 19, 22) {real, imag} */,
  {32'hbf435923, 32'h00000000} /* (12, 19, 21) {real, imag} */,
  {32'h3f410d11, 32'h00000000} /* (12, 19, 20) {real, imag} */,
  {32'h3f68c00a, 32'h00000000} /* (12, 19, 19) {real, imag} */,
  {32'h3f6d916a, 32'h00000000} /* (12, 19, 18) {real, imag} */,
  {32'h3f305dd6, 32'h00000000} /* (12, 19, 17) {real, imag} */,
  {32'h3f5db321, 32'h00000000} /* (12, 19, 16) {real, imag} */,
  {32'h3fbf38f0, 32'h00000000} /* (12, 19, 15) {real, imag} */,
  {32'h3f6c1574, 32'h00000000} /* (12, 19, 14) {real, imag} */,
  {32'h3f03e9da, 32'h00000000} /* (12, 19, 13) {real, imag} */,
  {32'h3f2f2615, 32'h00000000} /* (12, 19, 12) {real, imag} */,
  {32'h3f03e79a, 32'h00000000} /* (12, 19, 11) {real, imag} */,
  {32'hbf84abf1, 32'h00000000} /* (12, 19, 10) {real, imag} */,
  {32'hbfb3f110, 32'h00000000} /* (12, 19, 9) {real, imag} */,
  {32'hbef4a099, 32'h00000000} /* (12, 19, 8) {real, imag} */,
  {32'hbf59977a, 32'h00000000} /* (12, 19, 7) {real, imag} */,
  {32'hbf0a1389, 32'h00000000} /* (12, 19, 6) {real, imag} */,
  {32'hbf910a30, 32'h00000000} /* (12, 19, 5) {real, imag} */,
  {32'hbf83e12e, 32'h00000000} /* (12, 19, 4) {real, imag} */,
  {32'hbefa08f8, 32'h00000000} /* (12, 19, 3) {real, imag} */,
  {32'hbf562a96, 32'h00000000} /* (12, 19, 2) {real, imag} */,
  {32'hbf7f9259, 32'h00000000} /* (12, 19, 1) {real, imag} */,
  {32'hbf288872, 32'h00000000} /* (12, 19, 0) {real, imag} */,
  {32'hbec1f441, 32'h00000000} /* (12, 18, 31) {real, imag} */,
  {32'hbf89a716, 32'h00000000} /* (12, 18, 30) {real, imag} */,
  {32'hbfbacb9f, 32'h00000000} /* (12, 18, 29) {real, imag} */,
  {32'hbfaaed12, 32'h00000000} /* (12, 18, 28) {real, imag} */,
  {32'hbf82cf7f, 32'h00000000} /* (12, 18, 27) {real, imag} */,
  {32'hbf70c304, 32'h00000000} /* (12, 18, 26) {real, imag} */,
  {32'hbf02b972, 32'h00000000} /* (12, 18, 25) {real, imag} */,
  {32'hbf625997, 32'h00000000} /* (12, 18, 24) {real, imag} */,
  {32'hbf9de3e4, 32'h00000000} /* (12, 18, 23) {real, imag} */,
  {32'hbf92396f, 32'h00000000} /* (12, 18, 22) {real, imag} */,
  {32'hbf953f42, 32'h00000000} /* (12, 18, 21) {real, imag} */,
  {32'h3ed6eb8a, 32'h00000000} /* (12, 18, 20) {real, imag} */,
  {32'h3f4bee01, 32'h00000000} /* (12, 18, 19) {real, imag} */,
  {32'h3f98cddd, 32'h00000000} /* (12, 18, 18) {real, imag} */,
  {32'h3f2b3ea0, 32'h00000000} /* (12, 18, 17) {real, imag} */,
  {32'h3ec805a9, 32'h00000000} /* (12, 18, 16) {real, imag} */,
  {32'h3f42bc77, 32'h00000000} /* (12, 18, 15) {real, imag} */,
  {32'h3f5f7e47, 32'h00000000} /* (12, 18, 14) {real, imag} */,
  {32'h3f5cf478, 32'h00000000} /* (12, 18, 13) {real, imag} */,
  {32'h3f29efaf, 32'h00000000} /* (12, 18, 12) {real, imag} */,
  {32'h3f3fd965, 32'h00000000} /* (12, 18, 11) {real, imag} */,
  {32'hbf4686fb, 32'h00000000} /* (12, 18, 10) {real, imag} */,
  {32'hbf923cc7, 32'h00000000} /* (12, 18, 9) {real, imag} */,
  {32'hbee3ec81, 32'h00000000} /* (12, 18, 8) {real, imag} */,
  {32'hbf142ebf, 32'h00000000} /* (12, 18, 7) {real, imag} */,
  {32'hbf37b31d, 32'h00000000} /* (12, 18, 6) {real, imag} */,
  {32'hbf6de4b2, 32'h00000000} /* (12, 18, 5) {real, imag} */,
  {32'hbf4e28a2, 32'h00000000} /* (12, 18, 4) {real, imag} */,
  {32'hbf5449ba, 32'h00000000} /* (12, 18, 3) {real, imag} */,
  {32'hbf7fab04, 32'h00000000} /* (12, 18, 2) {real, imag} */,
  {32'hbf151d20, 32'h00000000} /* (12, 18, 1) {real, imag} */,
  {32'hbebfebe2, 32'h00000000} /* (12, 18, 0) {real, imag} */,
  {32'hbd30f09a, 32'h00000000} /* (12, 17, 31) {real, imag} */,
  {32'hbf38b837, 32'h00000000} /* (12, 17, 30) {real, imag} */,
  {32'hbfb386b8, 32'h00000000} /* (12, 17, 29) {real, imag} */,
  {32'hbff81b61, 32'h00000000} /* (12, 17, 28) {real, imag} */,
  {32'hbfae7185, 32'h00000000} /* (12, 17, 27) {real, imag} */,
  {32'hbf447cce, 32'h00000000} /* (12, 17, 26) {real, imag} */,
  {32'hbeeb6768, 32'h00000000} /* (12, 17, 25) {real, imag} */,
  {32'hbf635830, 32'h00000000} /* (12, 17, 24) {real, imag} */,
  {32'hbfacc30e, 32'h00000000} /* (12, 17, 23) {real, imag} */,
  {32'hbf8b67b1, 32'h00000000} /* (12, 17, 22) {real, imag} */,
  {32'hbf0167aa, 32'h00000000} /* (12, 17, 21) {real, imag} */,
  {32'h3f2b6e92, 32'h00000000} /* (12, 17, 20) {real, imag} */,
  {32'h3f4b9db2, 32'h00000000} /* (12, 17, 19) {real, imag} */,
  {32'h3f7fe10e, 32'h00000000} /* (12, 17, 18) {real, imag} */,
  {32'h3f468fec, 32'h00000000} /* (12, 17, 17) {real, imag} */,
  {32'h3f4ab729, 32'h00000000} /* (12, 17, 16) {real, imag} */,
  {32'h3f894a81, 32'h00000000} /* (12, 17, 15) {real, imag} */,
  {32'h3f62a4df, 32'h00000000} /* (12, 17, 14) {real, imag} */,
  {32'h3f5ad48f, 32'h00000000} /* (12, 17, 13) {real, imag} */,
  {32'h3f839557, 32'h00000000} /* (12, 17, 12) {real, imag} */,
  {32'h3edbbdf6, 32'h00000000} /* (12, 17, 11) {real, imag} */,
  {32'hbf22c0a8, 32'h00000000} /* (12, 17, 10) {real, imag} */,
  {32'hbf0961fd, 32'h00000000} /* (12, 17, 9) {real, imag} */,
  {32'hbedff643, 32'h00000000} /* (12, 17, 8) {real, imag} */,
  {32'hbf1972c5, 32'h00000000} /* (12, 17, 7) {real, imag} */,
  {32'hbf59b107, 32'h00000000} /* (12, 17, 6) {real, imag} */,
  {32'hbf447799, 32'h00000000} /* (12, 17, 5) {real, imag} */,
  {32'hbfa0baee, 32'h00000000} /* (12, 17, 4) {real, imag} */,
  {32'hbfc1f65c, 32'h00000000} /* (12, 17, 3) {real, imag} */,
  {32'hbf19d6eb, 32'h00000000} /* (12, 17, 2) {real, imag} */,
  {32'hbe6d0bec, 32'h00000000} /* (12, 17, 1) {real, imag} */,
  {32'hbe5887af, 32'h00000000} /* (12, 17, 0) {real, imag} */,
  {32'hbedaa7fd, 32'h00000000} /* (12, 16, 31) {real, imag} */,
  {32'hbf5e1116, 32'h00000000} /* (12, 16, 30) {real, imag} */,
  {32'hbf658a9a, 32'h00000000} /* (12, 16, 29) {real, imag} */,
  {32'hbf8c7d8e, 32'h00000000} /* (12, 16, 28) {real, imag} */,
  {32'hbf7e06d1, 32'h00000000} /* (12, 16, 27) {real, imag} */,
  {32'hbf87ee66, 32'h00000000} /* (12, 16, 26) {real, imag} */,
  {32'hbf88e821, 32'h00000000} /* (12, 16, 25) {real, imag} */,
  {32'hbfa872d3, 32'h00000000} /* (12, 16, 24) {real, imag} */,
  {32'hbfae8133, 32'h00000000} /* (12, 16, 23) {real, imag} */,
  {32'hbf92211c, 32'h00000000} /* (12, 16, 22) {real, imag} */,
  {32'h3d83ace4, 32'h00000000} /* (12, 16, 21) {real, imag} */,
  {32'h3f955528, 32'h00000000} /* (12, 16, 20) {real, imag} */,
  {32'h3f841aa2, 32'h00000000} /* (12, 16, 19) {real, imag} */,
  {32'h3f76a5b8, 32'h00000000} /* (12, 16, 18) {real, imag} */,
  {32'h3f67faca, 32'h00000000} /* (12, 16, 17) {real, imag} */,
  {32'h3f89131c, 32'h00000000} /* (12, 16, 16) {real, imag} */,
  {32'h3f4f1e4b, 32'h00000000} /* (12, 16, 15) {real, imag} */,
  {32'h3f802624, 32'h00000000} /* (12, 16, 14) {real, imag} */,
  {32'h3fa36c5e, 32'h00000000} /* (12, 16, 13) {real, imag} */,
  {32'h3f971732, 32'h00000000} /* (12, 16, 12) {real, imag} */,
  {32'h3e7de835, 32'h00000000} /* (12, 16, 11) {real, imag} */,
  {32'hbf0f7c1c, 32'h00000000} /* (12, 16, 10) {real, imag} */,
  {32'hbf043937, 32'h00000000} /* (12, 16, 9) {real, imag} */,
  {32'hbe28e0d3, 32'h00000000} /* (12, 16, 8) {real, imag} */,
  {32'hbf11062c, 32'h00000000} /* (12, 16, 7) {real, imag} */,
  {32'hbf3040db, 32'h00000000} /* (12, 16, 6) {real, imag} */,
  {32'hbf1ddc55, 32'h00000000} /* (12, 16, 5) {real, imag} */,
  {32'hbf773ba2, 32'h00000000} /* (12, 16, 4) {real, imag} */,
  {32'hbf90db58, 32'h00000000} /* (12, 16, 3) {real, imag} */,
  {32'hbe3e3657, 32'h00000000} /* (12, 16, 2) {real, imag} */,
  {32'hbf2df6bc, 32'h00000000} /* (12, 16, 1) {real, imag} */,
  {32'hbf42ba6c, 32'h00000000} /* (12, 16, 0) {real, imag} */,
  {32'hbf02c3bb, 32'h00000000} /* (12, 15, 31) {real, imag} */,
  {32'hbf2c9c56, 32'h00000000} /* (12, 15, 30) {real, imag} */,
  {32'hbf4ef426, 32'h00000000} /* (12, 15, 29) {real, imag} */,
  {32'hbfb5676c, 32'h00000000} /* (12, 15, 28) {real, imag} */,
  {32'hbf8f959e, 32'h00000000} /* (12, 15, 27) {real, imag} */,
  {32'hbf8d6a21, 32'h00000000} /* (12, 15, 26) {real, imag} */,
  {32'hbf98ae96, 32'h00000000} /* (12, 15, 25) {real, imag} */,
  {32'hbf9927bf, 32'h00000000} /* (12, 15, 24) {real, imag} */,
  {32'hbf88147c, 32'h00000000} /* (12, 15, 23) {real, imag} */,
  {32'hbf37e33a, 32'h00000000} /* (12, 15, 22) {real, imag} */,
  {32'h3d555611, 32'h00000000} /* (12, 15, 21) {real, imag} */,
  {32'h3f3e4ec1, 32'h00000000} /* (12, 15, 20) {real, imag} */,
  {32'h3f35cf77, 32'h00000000} /* (12, 15, 19) {real, imag} */,
  {32'h3f584777, 32'h00000000} /* (12, 15, 18) {real, imag} */,
  {32'h3f59e917, 32'h00000000} /* (12, 15, 17) {real, imag} */,
  {32'h3f2c7185, 32'h00000000} /* (12, 15, 16) {real, imag} */,
  {32'h3f33a7d4, 32'h00000000} /* (12, 15, 15) {real, imag} */,
  {32'h3f3a29e6, 32'h00000000} /* (12, 15, 14) {real, imag} */,
  {32'h3f4e38c2, 32'h00000000} /* (12, 15, 13) {real, imag} */,
  {32'h3f4d8e74, 32'h00000000} /* (12, 15, 12) {real, imag} */,
  {32'h3ea4c1c1, 32'h00000000} /* (12, 15, 11) {real, imag} */,
  {32'hbeb3d2db, 32'h00000000} /* (12, 15, 10) {real, imag} */,
  {32'hbf05f806, 32'h00000000} /* (12, 15, 9) {real, imag} */,
  {32'hbf18b1c2, 32'h00000000} /* (12, 15, 8) {real, imag} */,
  {32'hbf941074, 32'h00000000} /* (12, 15, 7) {real, imag} */,
  {32'hbfa270c6, 32'h00000000} /* (12, 15, 6) {real, imag} */,
  {32'hbf0f249d, 32'h00000000} /* (12, 15, 5) {real, imag} */,
  {32'hbf3388d0, 32'h00000000} /* (12, 15, 4) {real, imag} */,
  {32'hbf2eae7b, 32'h00000000} /* (12, 15, 3) {real, imag} */,
  {32'hbef2370a, 32'h00000000} /* (12, 15, 2) {real, imag} */,
  {32'hbfa7140b, 32'h00000000} /* (12, 15, 1) {real, imag} */,
  {32'hbfb7f2e6, 32'h00000000} /* (12, 15, 0) {real, imag} */,
  {32'hbf2bb39b, 32'h00000000} /* (12, 14, 31) {real, imag} */,
  {32'hbf75bdda, 32'h00000000} /* (12, 14, 30) {real, imag} */,
  {32'hbf551621, 32'h00000000} /* (12, 14, 29) {real, imag} */,
  {32'hbf96c45c, 32'h00000000} /* (12, 14, 28) {real, imag} */,
  {32'hbfa31804, 32'h00000000} /* (12, 14, 27) {real, imag} */,
  {32'hbf81fdb7, 32'h00000000} /* (12, 14, 26) {real, imag} */,
  {32'hbf402c40, 32'h00000000} /* (12, 14, 25) {real, imag} */,
  {32'hbf5dc0ed, 32'h00000000} /* (12, 14, 24) {real, imag} */,
  {32'hbf84752e, 32'h00000000} /* (12, 14, 23) {real, imag} */,
  {32'hbf670ada, 32'h00000000} /* (12, 14, 22) {real, imag} */,
  {32'hbf078b73, 32'h00000000} /* (12, 14, 21) {real, imag} */,
  {32'h3ef5ce98, 32'h00000000} /* (12, 14, 20) {real, imag} */,
  {32'h3ef612d5, 32'h00000000} /* (12, 14, 19) {real, imag} */,
  {32'h3f2e664b, 32'h00000000} /* (12, 14, 18) {real, imag} */,
  {32'h3f3e121f, 32'h00000000} /* (12, 14, 17) {real, imag} */,
  {32'h3f29b909, 32'h00000000} /* (12, 14, 16) {real, imag} */,
  {32'h3f8c67c1, 32'h00000000} /* (12, 14, 15) {real, imag} */,
  {32'h3f816f4e, 32'h00000000} /* (12, 14, 14) {real, imag} */,
  {32'h3f178b9c, 32'h00000000} /* (12, 14, 13) {real, imag} */,
  {32'h3f4d04d8, 32'h00000000} /* (12, 14, 12) {real, imag} */,
  {32'h3f59f32a, 32'h00000000} /* (12, 14, 11) {real, imag} */,
  {32'h3d9d1dd4, 32'h00000000} /* (12, 14, 10) {real, imag} */,
  {32'hbec410b9, 32'h00000000} /* (12, 14, 9) {real, imag} */,
  {32'hbf487896, 32'h00000000} /* (12, 14, 8) {real, imag} */,
  {32'hbfe9b06d, 32'h00000000} /* (12, 14, 7) {real, imag} */,
  {32'hbfc52de4, 32'h00000000} /* (12, 14, 6) {real, imag} */,
  {32'hbeeaec97, 32'h00000000} /* (12, 14, 5) {real, imag} */,
  {32'hbf0f4ac0, 32'h00000000} /* (12, 14, 4) {real, imag} */,
  {32'hbef193e4, 32'h00000000} /* (12, 14, 3) {real, imag} */,
  {32'hbf5c5cf0, 32'h00000000} /* (12, 14, 2) {real, imag} */,
  {32'hbff1f651, 32'h00000000} /* (12, 14, 1) {real, imag} */,
  {32'hbfd26009, 32'h00000000} /* (12, 14, 0) {real, imag} */,
  {32'hbf6a2e1e, 32'h00000000} /* (12, 13, 31) {real, imag} */,
  {32'hbfde71c8, 32'h00000000} /* (12, 13, 30) {real, imag} */,
  {32'hbfa256a8, 32'h00000000} /* (12, 13, 29) {real, imag} */,
  {32'hbfb4c634, 32'h00000000} /* (12, 13, 28) {real, imag} */,
  {32'hbf77a7cb, 32'h00000000} /* (12, 13, 27) {real, imag} */,
  {32'hbe75c6fc, 32'h00000000} /* (12, 13, 26) {real, imag} */,
  {32'hbf39e11a, 32'h00000000} /* (12, 13, 25) {real, imag} */,
  {32'hbfa27a9c, 32'h00000000} /* (12, 13, 24) {real, imag} */,
  {32'hbf99db3d, 32'h00000000} /* (12, 13, 23) {real, imag} */,
  {32'hbfaf4e8e, 32'h00000000} /* (12, 13, 22) {real, imag} */,
  {32'hbf40e992, 32'h00000000} /* (12, 13, 21) {real, imag} */,
  {32'h3eaeaf0f, 32'h00000000} /* (12, 13, 20) {real, imag} */,
  {32'h3f3694a2, 32'h00000000} /* (12, 13, 19) {real, imag} */,
  {32'h3f931313, 32'h00000000} /* (12, 13, 18) {real, imag} */,
  {32'h3f74b67f, 32'h00000000} /* (12, 13, 17) {real, imag} */,
  {32'h3f2cc2b0, 32'h00000000} /* (12, 13, 16) {real, imag} */,
  {32'h3f788926, 32'h00000000} /* (12, 13, 15) {real, imag} */,
  {32'h3f9a0499, 32'h00000000} /* (12, 13, 14) {real, imag} */,
  {32'h3f06ee9e, 32'h00000000} /* (12, 13, 13) {real, imag} */,
  {32'h3f240286, 32'h00000000} /* (12, 13, 12) {real, imag} */,
  {32'h3f599d94, 32'h00000000} /* (12, 13, 11) {real, imag} */,
  {32'hbe680913, 32'h00000000} /* (12, 13, 10) {real, imag} */,
  {32'hbf20ae3c, 32'h00000000} /* (12, 13, 9) {real, imag} */,
  {32'hbf137aa8, 32'h00000000} /* (12, 13, 8) {real, imag} */,
  {32'hbf9c223c, 32'h00000000} /* (12, 13, 7) {real, imag} */,
  {32'hbf7df678, 32'h00000000} /* (12, 13, 6) {real, imag} */,
  {32'hbf16d95d, 32'h00000000} /* (12, 13, 5) {real, imag} */,
  {32'hbf3ca42d, 32'h00000000} /* (12, 13, 4) {real, imag} */,
  {32'hbf397dd4, 32'h00000000} /* (12, 13, 3) {real, imag} */,
  {32'hbf95f000, 32'h00000000} /* (12, 13, 2) {real, imag} */,
  {32'hbfbffdc1, 32'h00000000} /* (12, 13, 1) {real, imag} */,
  {32'hbf68e1d4, 32'h00000000} /* (12, 13, 0) {real, imag} */,
  {32'hbf837451, 32'h00000000} /* (12, 12, 31) {real, imag} */,
  {32'hbfcc8f7f, 32'h00000000} /* (12, 12, 30) {real, imag} */,
  {32'hbfaa883b, 32'h00000000} /* (12, 12, 29) {real, imag} */,
  {32'hbfbc314e, 32'h00000000} /* (12, 12, 28) {real, imag} */,
  {32'hbf61d262, 32'h00000000} /* (12, 12, 27) {real, imag} */,
  {32'hbe5c62ee, 32'h00000000} /* (12, 12, 26) {real, imag} */,
  {32'hbf19bea1, 32'h00000000} /* (12, 12, 25) {real, imag} */,
  {32'hbfa68475, 32'h00000000} /* (12, 12, 24) {real, imag} */,
  {32'hbf8597eb, 32'h00000000} /* (12, 12, 23) {real, imag} */,
  {32'hbf4fe080, 32'h00000000} /* (12, 12, 22) {real, imag} */,
  {32'hbefbe233, 32'h00000000} /* (12, 12, 21) {real, imag} */,
  {32'h3ee1ceb9, 32'h00000000} /* (12, 12, 20) {real, imag} */,
  {32'h3f8987ad, 32'h00000000} /* (12, 12, 19) {real, imag} */,
  {32'h3fb2ff67, 32'h00000000} /* (12, 12, 18) {real, imag} */,
  {32'h3faacdc0, 32'h00000000} /* (12, 12, 17) {real, imag} */,
  {32'h3fa47da5, 32'h00000000} /* (12, 12, 16) {real, imag} */,
  {32'h3f6d238d, 32'h00000000} /* (12, 12, 15) {real, imag} */,
  {32'h3f69eaba, 32'h00000000} /* (12, 12, 14) {real, imag} */,
  {32'h3f139953, 32'h00000000} /* (12, 12, 13) {real, imag} */,
  {32'h3f1c460a, 32'h00000000} /* (12, 12, 12) {real, imag} */,
  {32'h3f1181b9, 32'h00000000} /* (12, 12, 11) {real, imag} */,
  {32'hbf334cfc, 32'h00000000} /* (12, 12, 10) {real, imag} */,
  {32'hbf9a8383, 32'h00000000} /* (12, 12, 9) {real, imag} */,
  {32'hbf37914e, 32'h00000000} /* (12, 12, 8) {real, imag} */,
  {32'hbf8c1fd5, 32'h00000000} /* (12, 12, 7) {real, imag} */,
  {32'hbfd32292, 32'h00000000} /* (12, 12, 6) {real, imag} */,
  {32'hbfc4c249, 32'h00000000} /* (12, 12, 5) {real, imag} */,
  {32'hbf7a9c52, 32'h00000000} /* (12, 12, 4) {real, imag} */,
  {32'hbf8e8c3f, 32'h00000000} /* (12, 12, 3) {real, imag} */,
  {32'hbf8bd93d, 32'h00000000} /* (12, 12, 2) {real, imag} */,
  {32'hbf6aee71, 32'h00000000} /* (12, 12, 1) {real, imag} */,
  {32'hbec53d29, 32'h00000000} /* (12, 12, 0) {real, imag} */,
  {32'hbed317c0, 32'h00000000} /* (12, 11, 31) {real, imag} */,
  {32'hbf2f5898, 32'h00000000} /* (12, 11, 30) {real, imag} */,
  {32'hbe6fe3d6, 32'h00000000} /* (12, 11, 29) {real, imag} */,
  {32'hbf0ca382, 32'h00000000} /* (12, 11, 28) {real, imag} */,
  {32'hbec71284, 32'h00000000} /* (12, 11, 27) {real, imag} */,
  {32'hbe6ef6e6, 32'h00000000} /* (12, 11, 26) {real, imag} */,
  {32'hbe4be902, 32'h00000000} /* (12, 11, 25) {real, imag} */,
  {32'hbf7b81a1, 32'h00000000} /* (12, 11, 24) {real, imag} */,
  {32'hbf8c45ea, 32'h00000000} /* (12, 11, 23) {real, imag} */,
  {32'hbeff39ae, 32'h00000000} /* (12, 11, 22) {real, imag} */,
  {32'hbe25100e, 32'h00000000} /* (12, 11, 21) {real, imag} */,
  {32'h3eca144e, 32'h00000000} /* (12, 11, 20) {real, imag} */,
  {32'h3f269396, 32'h00000000} /* (12, 11, 19) {real, imag} */,
  {32'h3f2c6850, 32'h00000000} /* (12, 11, 18) {real, imag} */,
  {32'h3f5cfc9a, 32'h00000000} /* (12, 11, 17) {real, imag} */,
  {32'h3f304bc9, 32'h00000000} /* (12, 11, 16) {real, imag} */,
  {32'h3eca4544, 32'h00000000} /* (12, 11, 15) {real, imag} */,
  {32'h3f50a209, 32'h00000000} /* (12, 11, 14) {real, imag} */,
  {32'h3f485556, 32'h00000000} /* (12, 11, 13) {real, imag} */,
  {32'h3f228eee, 32'h00000000} /* (12, 11, 12) {real, imag} */,
  {32'h3ee0c8a9, 32'h00000000} /* (12, 11, 11) {real, imag} */,
  {32'hbf3510ab, 32'h00000000} /* (12, 11, 10) {real, imag} */,
  {32'hbfb444b1, 32'h00000000} /* (12, 11, 9) {real, imag} */,
  {32'hbf5fa11a, 32'h00000000} /* (12, 11, 8) {real, imag} */,
  {32'hbf7c8e06, 32'h00000000} /* (12, 11, 7) {real, imag} */,
  {32'hbfbfae70, 32'h00000000} /* (12, 11, 6) {real, imag} */,
  {32'hbf838d2a, 32'h00000000} /* (12, 11, 5) {real, imag} */,
  {32'hbf608142, 32'h00000000} /* (12, 11, 4) {real, imag} */,
  {32'hbf31778f, 32'h00000000} /* (12, 11, 3) {real, imag} */,
  {32'hbf0902a4, 32'h00000000} /* (12, 11, 2) {real, imag} */,
  {32'hbf248eea, 32'h00000000} /* (12, 11, 1) {real, imag} */,
  {32'hbed9bcdc, 32'h00000000} /* (12, 11, 0) {real, imag} */,
  {32'h3ece1655, 32'h00000000} /* (12, 10, 31) {real, imag} */,
  {32'h3f0880cb, 32'h00000000} /* (12, 10, 30) {real, imag} */,
  {32'h3f145cec, 32'h00000000} /* (12, 10, 29) {real, imag} */,
  {32'h3f880e5d, 32'h00000000} /* (12, 10, 28) {real, imag} */,
  {32'h3f84b845, 32'h00000000} /* (12, 10, 27) {real, imag} */,
  {32'h3eca18a3, 32'h00000000} /* (12, 10, 26) {real, imag} */,
  {32'h3f07d9be, 32'h00000000} /* (12, 10, 25) {real, imag} */,
  {32'h3edf0189, 32'h00000000} /* (12, 10, 24) {real, imag} */,
  {32'hbdaae059, 32'h00000000} /* (12, 10, 23) {real, imag} */,
  {32'h3c02b7ed, 32'h00000000} /* (12, 10, 22) {real, imag} */,
  {32'hbe033f37, 32'h00000000} /* (12, 10, 21) {real, imag} */,
  {32'hbee6c93a, 32'h00000000} /* (12, 10, 20) {real, imag} */,
  {32'hbef14121, 32'h00000000} /* (12, 10, 19) {real, imag} */,
  {32'hbf1da4a8, 32'h00000000} /* (12, 10, 18) {real, imag} */,
  {32'hbe03913a, 32'h00000000} /* (12, 10, 17) {real, imag} */,
  {32'hbf042aa6, 32'h00000000} /* (12, 10, 16) {real, imag} */,
  {32'hbecbcbde, 32'h00000000} /* (12, 10, 15) {real, imag} */,
  {32'h3cac21c1, 32'h00000000} /* (12, 10, 14) {real, imag} */,
  {32'hbe8a8d0e, 32'h00000000} /* (12, 10, 13) {real, imag} */,
  {32'hbe84081d, 32'h00000000} /* (12, 10, 12) {real, imag} */,
  {32'hbf05b851, 32'h00000000} /* (12, 10, 11) {real, imag} */,
  {32'hbead238e, 32'h00000000} /* (12, 10, 10) {real, imag} */,
  {32'hbe0f1738, 32'h00000000} /* (12, 10, 9) {real, imag} */,
  {32'h3e72c870, 32'h00000000} /* (12, 10, 8) {real, imag} */,
  {32'h3ed2bc71, 32'h00000000} /* (12, 10, 7) {real, imag} */,
  {32'h3e7319bd, 32'h00000000} /* (12, 10, 6) {real, imag} */,
  {32'h3f7da4a8, 32'h00000000} /* (12, 10, 5) {real, imag} */,
  {32'h3ef893d4, 32'h00000000} /* (12, 10, 4) {real, imag} */,
  {32'h3de47a6f, 32'h00000000} /* (12, 10, 3) {real, imag} */,
  {32'h3e3b8af5, 32'h00000000} /* (12, 10, 2) {real, imag} */,
  {32'h3f31caad, 32'h00000000} /* (12, 10, 1) {real, imag} */,
  {32'h3ee0aea2, 32'h00000000} /* (12, 10, 0) {real, imag} */,
  {32'h3ee9f524, 32'h00000000} /* (12, 9, 31) {real, imag} */,
  {32'h3f067747, 32'h00000000} /* (12, 9, 30) {real, imag} */,
  {32'h3f2439d5, 32'h00000000} /* (12, 9, 29) {real, imag} */,
  {32'h3fb4d049, 32'h00000000} /* (12, 9, 28) {real, imag} */,
  {32'h3f99a48f, 32'h00000000} /* (12, 9, 27) {real, imag} */,
  {32'h3f8285ff, 32'h00000000} /* (12, 9, 26) {real, imag} */,
  {32'h3f83e6e9, 32'h00000000} /* (12, 9, 25) {real, imag} */,
  {32'h3fb21d20, 32'h00000000} /* (12, 9, 24) {real, imag} */,
  {32'h3f49e9aa, 32'h00000000} /* (12, 9, 23) {real, imag} */,
  {32'h3ecb0e10, 32'h00000000} /* (12, 9, 22) {real, imag} */,
  {32'h3eadadfc, 32'h00000000} /* (12, 9, 21) {real, imag} */,
  {32'hbee79231, 32'h00000000} /* (12, 9, 20) {real, imag} */,
  {32'hbf192842, 32'h00000000} /* (12, 9, 19) {real, imag} */,
  {32'hbf47828f, 32'h00000000} /* (12, 9, 18) {real, imag} */,
  {32'hbf5141aa, 32'h00000000} /* (12, 9, 17) {real, imag} */,
  {32'hbf941eeb, 32'h00000000} /* (12, 9, 16) {real, imag} */,
  {32'hbf6ee522, 32'h00000000} /* (12, 9, 15) {real, imag} */,
  {32'hbf844cb4, 32'h00000000} /* (12, 9, 14) {real, imag} */,
  {32'hbf782164, 32'h00000000} /* (12, 9, 13) {real, imag} */,
  {32'hbf40f4a9, 32'h00000000} /* (12, 9, 12) {real, imag} */,
  {32'hbf21f2d5, 32'h00000000} /* (12, 9, 11) {real, imag} */,
  {32'h3eaca7b3, 32'h00000000} /* (12, 9, 10) {real, imag} */,
  {32'h3f3edc36, 32'h00000000} /* (12, 9, 9) {real, imag} */,
  {32'h3f857083, 32'h00000000} /* (12, 9, 8) {real, imag} */,
  {32'h3f63863b, 32'h00000000} /* (12, 9, 7) {real, imag} */,
  {32'h3f1aea96, 32'h00000000} /* (12, 9, 6) {real, imag} */,
  {32'h3f677aba, 32'h00000000} /* (12, 9, 5) {real, imag} */,
  {32'h3ed7e420, 32'h00000000} /* (12, 9, 4) {real, imag} */,
  {32'h3e860257, 32'h00000000} /* (12, 9, 3) {real, imag} */,
  {32'h3e59bf4c, 32'h00000000} /* (12, 9, 2) {real, imag} */,
  {32'h3f4521b9, 32'h00000000} /* (12, 9, 1) {real, imag} */,
  {32'h3ed4d7f9, 32'h00000000} /* (12, 9, 0) {real, imag} */,
  {32'h3eb7430b, 32'h00000000} /* (12, 8, 31) {real, imag} */,
  {32'h3efa4f81, 32'h00000000} /* (12, 8, 30) {real, imag} */,
  {32'h3f06cfb6, 32'h00000000} /* (12, 8, 29) {real, imag} */,
  {32'h3f98f887, 32'h00000000} /* (12, 8, 28) {real, imag} */,
  {32'h3f8d77a0, 32'h00000000} /* (12, 8, 27) {real, imag} */,
  {32'h3f983173, 32'h00000000} /* (12, 8, 26) {real, imag} */,
  {32'h3f583b01, 32'h00000000} /* (12, 8, 25) {real, imag} */,
  {32'h3ff38e83, 32'h00000000} /* (12, 8, 24) {real, imag} */,
  {32'h3fa04abf, 32'h00000000} /* (12, 8, 23) {real, imag} */,
  {32'h3f089fb2, 32'h00000000} /* (12, 8, 22) {real, imag} */,
  {32'h3f239874, 32'h00000000} /* (12, 8, 21) {real, imag} */,
  {32'hbef8af57, 32'h00000000} /* (12, 8, 20) {real, imag} */,
  {32'hbf174b65, 32'h00000000} /* (12, 8, 19) {real, imag} */,
  {32'hbf18fe86, 32'h00000000} /* (12, 8, 18) {real, imag} */,
  {32'hbf3c7fc0, 32'h00000000} /* (12, 8, 17) {real, imag} */,
  {32'hbf8bff74, 32'h00000000} /* (12, 8, 16) {real, imag} */,
  {32'hbfda2cc5, 32'h00000000} /* (12, 8, 15) {real, imag} */,
  {32'hbf8e4726, 32'h00000000} /* (12, 8, 14) {real, imag} */,
  {32'hbeb12e90, 32'h00000000} /* (12, 8, 13) {real, imag} */,
  {32'hbf04524f, 32'h00000000} /* (12, 8, 12) {real, imag} */,
  {32'hbeb9673a, 32'h00000000} /* (12, 8, 11) {real, imag} */,
  {32'h3f2162a0, 32'h00000000} /* (12, 8, 10) {real, imag} */,
  {32'h3f2d009b, 32'h00000000} /* (12, 8, 9) {real, imag} */,
  {32'h3f5708cd, 32'h00000000} /* (12, 8, 8) {real, imag} */,
  {32'h3f2402b2, 32'h00000000} /* (12, 8, 7) {real, imag} */,
  {32'h3eb3eef4, 32'h00000000} /* (12, 8, 6) {real, imag} */,
  {32'h3f105adf, 32'h00000000} /* (12, 8, 5) {real, imag} */,
  {32'h3f101394, 32'h00000000} /* (12, 8, 4) {real, imag} */,
  {32'h3e3e7016, 32'h00000000} /* (12, 8, 3) {real, imag} */,
  {32'h3df879f6, 32'h00000000} /* (12, 8, 2) {real, imag} */,
  {32'h3ef5b05f, 32'h00000000} /* (12, 8, 1) {real, imag} */,
  {32'h3e944382, 32'h00000000} /* (12, 8, 0) {real, imag} */,
  {32'h3e95978f, 32'h00000000} /* (12, 7, 31) {real, imag} */,
  {32'h3f138308, 32'h00000000} /* (12, 7, 30) {real, imag} */,
  {32'h3edb3dcc, 32'h00000000} /* (12, 7, 29) {real, imag} */,
  {32'h3f13ac69, 32'h00000000} /* (12, 7, 28) {real, imag} */,
  {32'h3f4f60a8, 32'h00000000} /* (12, 7, 27) {real, imag} */,
  {32'h3f37fdd7, 32'h00000000} /* (12, 7, 26) {real, imag} */,
  {32'h3ee4cb1e, 32'h00000000} /* (12, 7, 25) {real, imag} */,
  {32'h3f633a0d, 32'h00000000} /* (12, 7, 24) {real, imag} */,
  {32'h3f36ffaa, 32'h00000000} /* (12, 7, 23) {real, imag} */,
  {32'h3f5e4b21, 32'h00000000} /* (12, 7, 22) {real, imag} */,
  {32'h3f4c9dd7, 32'h00000000} /* (12, 7, 21) {real, imag} */,
  {32'hbf2e72ee, 32'h00000000} /* (12, 7, 20) {real, imag} */,
  {32'hbf8f2e19, 32'h00000000} /* (12, 7, 19) {real, imag} */,
  {32'hbf7cb213, 32'h00000000} /* (12, 7, 18) {real, imag} */,
  {32'hbf2e5174, 32'h00000000} /* (12, 7, 17) {real, imag} */,
  {32'hbf950e03, 32'h00000000} /* (12, 7, 16) {real, imag} */,
  {32'hbfcbf821, 32'h00000000} /* (12, 7, 15) {real, imag} */,
  {32'hbf88dd89, 32'h00000000} /* (12, 7, 14) {real, imag} */,
  {32'hbf13e2f2, 32'h00000000} /* (12, 7, 13) {real, imag} */,
  {32'hbf9a88e8, 32'h00000000} /* (12, 7, 12) {real, imag} */,
  {32'hbf5622b7, 32'h00000000} /* (12, 7, 11) {real, imag} */,
  {32'h3ed00cf9, 32'h00000000} /* (12, 7, 10) {real, imag} */,
  {32'h3eedf640, 32'h00000000} /* (12, 7, 9) {real, imag} */,
  {32'h3f801c0d, 32'h00000000} /* (12, 7, 8) {real, imag} */,
  {32'h3f6bf2fd, 32'h00000000} /* (12, 7, 7) {real, imag} */,
  {32'h3f01fa3b, 32'h00000000} /* (12, 7, 6) {real, imag} */,
  {32'h3f2829e7, 32'h00000000} /* (12, 7, 5) {real, imag} */,
  {32'h3fc2b1e3, 32'h00000000} /* (12, 7, 4) {real, imag} */,
  {32'h3f73341c, 32'h00000000} /* (12, 7, 3) {real, imag} */,
  {32'h3f388838, 32'h00000000} /* (12, 7, 2) {real, imag} */,
  {32'h3f1a8a9e, 32'h00000000} /* (12, 7, 1) {real, imag} */,
  {32'h3de5d0f3, 32'h00000000} /* (12, 7, 0) {real, imag} */,
  {32'h3e3a84d2, 32'h00000000} /* (12, 6, 31) {real, imag} */,
  {32'h3e73eee9, 32'h00000000} /* (12, 6, 30) {real, imag} */,
  {32'h3ec83dd3, 32'h00000000} /* (12, 6, 29) {real, imag} */,
  {32'h3f2717ea, 32'h00000000} /* (12, 6, 28) {real, imag} */,
  {32'h3f516126, 32'h00000000} /* (12, 6, 27) {real, imag} */,
  {32'h3f633818, 32'h00000000} /* (12, 6, 26) {real, imag} */,
  {32'h3f5a011f, 32'h00000000} /* (12, 6, 25) {real, imag} */,
  {32'h3f1a99c8, 32'h00000000} /* (12, 6, 24) {real, imag} */,
  {32'h3f11e8ce, 32'h00000000} /* (12, 6, 23) {real, imag} */,
  {32'h3f47979b, 32'h00000000} /* (12, 6, 22) {real, imag} */,
  {32'h3f61e5b7, 32'h00000000} /* (12, 6, 21) {real, imag} */,
  {32'hbe8442bc, 32'h00000000} /* (12, 6, 20) {real, imag} */,
  {32'hbf2c15e8, 32'h00000000} /* (12, 6, 19) {real, imag} */,
  {32'hbf7dd582, 32'h00000000} /* (12, 6, 18) {real, imag} */,
  {32'hbf59314d, 32'h00000000} /* (12, 6, 17) {real, imag} */,
  {32'hbfb2c950, 32'h00000000} /* (12, 6, 16) {real, imag} */,
  {32'hbf4f1935, 32'h00000000} /* (12, 6, 15) {real, imag} */,
  {32'hbf90458f, 32'h00000000} /* (12, 6, 14) {real, imag} */,
  {32'hbf7faedb, 32'h00000000} /* (12, 6, 13) {real, imag} */,
  {32'hbf84cb24, 32'h00000000} /* (12, 6, 12) {real, imag} */,
  {32'hbf61068d, 32'h00000000} /* (12, 6, 11) {real, imag} */,
  {32'hbe6a20a4, 32'h00000000} /* (12, 6, 10) {real, imag} */,
  {32'h3e8869f2, 32'h00000000} /* (12, 6, 9) {real, imag} */,
  {32'h3fa21b5c, 32'h00000000} /* (12, 6, 8) {real, imag} */,
  {32'h3f72b175, 32'h00000000} /* (12, 6, 7) {real, imag} */,
  {32'h3efe0d95, 32'h00000000} /* (12, 6, 6) {real, imag} */,
  {32'h3eff19be, 32'h00000000} /* (12, 6, 5) {real, imag} */,
  {32'h3f78f165, 32'h00000000} /* (12, 6, 4) {real, imag} */,
  {32'h3f848c34, 32'h00000000} /* (12, 6, 3) {real, imag} */,
  {32'h3f932216, 32'h00000000} /* (12, 6, 2) {real, imag} */,
  {32'h3f725fb2, 32'h00000000} /* (12, 6, 1) {real, imag} */,
  {32'h3e6fca78, 32'h00000000} /* (12, 6, 0) {real, imag} */,
  {32'h3e944a3f, 32'h00000000} /* (12, 5, 31) {real, imag} */,
  {32'h3f2fb5f8, 32'h00000000} /* (12, 5, 30) {real, imag} */,
  {32'h3f9311ce, 32'h00000000} /* (12, 5, 29) {real, imag} */,
  {32'h3f896d40, 32'h00000000} /* (12, 5, 28) {real, imag} */,
  {32'h3faa089f, 32'h00000000} /* (12, 5, 27) {real, imag} */,
  {32'h3f822232, 32'h00000000} /* (12, 5, 26) {real, imag} */,
  {32'h3f540e71, 32'h00000000} /* (12, 5, 25) {real, imag} */,
  {32'h3f2e01ce, 32'h00000000} /* (12, 5, 24) {real, imag} */,
  {32'h3f8b0e22, 32'h00000000} /* (12, 5, 23) {real, imag} */,
  {32'h3f18dd6c, 32'h00000000} /* (12, 5, 22) {real, imag} */,
  {32'h3f4690e8, 32'h00000000} /* (12, 5, 21) {real, imag} */,
  {32'h3ee3b417, 32'h00000000} /* (12, 5, 20) {real, imag} */,
  {32'h3eb7fee9, 32'h00000000} /* (12, 5, 19) {real, imag} */,
  {32'h3f457d7d, 32'h00000000} /* (12, 5, 18) {real, imag} */,
  {32'h3f58dce3, 32'h00000000} /* (12, 5, 17) {real, imag} */,
  {32'hbe349b96, 32'h00000000} /* (12, 5, 16) {real, imag} */,
  {32'hbf4a4731, 32'h00000000} /* (12, 5, 15) {real, imag} */,
  {32'hbf6e628d, 32'h00000000} /* (12, 5, 14) {real, imag} */,
  {32'hbf0c7d90, 32'h00000000} /* (12, 5, 13) {real, imag} */,
  {32'hbf489323, 32'h00000000} /* (12, 5, 12) {real, imag} */,
  {32'hbf8c7612, 32'h00000000} /* (12, 5, 11) {real, imag} */,
  {32'hbf003c38, 32'h00000000} /* (12, 5, 10) {real, imag} */,
  {32'hbe7a7a6d, 32'h00000000} /* (12, 5, 9) {real, imag} */,
  {32'h3cfbc168, 32'h00000000} /* (12, 5, 8) {real, imag} */,
  {32'hbeb89e3f, 32'h00000000} /* (12, 5, 7) {real, imag} */,
  {32'hbe9fe15c, 32'h00000000} /* (12, 5, 6) {real, imag} */,
  {32'h3e433f8e, 32'h00000000} /* (12, 5, 5) {real, imag} */,
  {32'h3f0b155a, 32'h00000000} /* (12, 5, 4) {real, imag} */,
  {32'h3f8dbf7d, 32'h00000000} /* (12, 5, 3) {real, imag} */,
  {32'h3f96150d, 32'h00000000} /* (12, 5, 2) {real, imag} */,
  {32'h3f807c4e, 32'h00000000} /* (12, 5, 1) {real, imag} */,
  {32'h3eac4a30, 32'h00000000} /* (12, 5, 0) {real, imag} */,
  {32'h3ee21fb6, 32'h00000000} /* (12, 4, 31) {real, imag} */,
  {32'h3fa1cc59, 32'h00000000} /* (12, 4, 30) {real, imag} */,
  {32'h3fa5f538, 32'h00000000} /* (12, 4, 29) {real, imag} */,
  {32'h3f34fd22, 32'h00000000} /* (12, 4, 28) {real, imag} */,
  {32'h3f8f3f1e, 32'h00000000} /* (12, 4, 27) {real, imag} */,
  {32'h3f64e3cb, 32'h00000000} /* (12, 4, 26) {real, imag} */,
  {32'h3f54314d, 32'h00000000} /* (12, 4, 25) {real, imag} */,
  {32'h3ee3c5b1, 32'h00000000} /* (12, 4, 24) {real, imag} */,
  {32'h3f8dff3f, 32'h00000000} /* (12, 4, 23) {real, imag} */,
  {32'h3fa645e8, 32'h00000000} /* (12, 4, 22) {real, imag} */,
  {32'h3fcf8c9f, 32'h00000000} /* (12, 4, 21) {real, imag} */,
  {32'h3fae5716, 32'h00000000} /* (12, 4, 20) {real, imag} */,
  {32'h3f80ae2b, 32'h00000000} /* (12, 4, 19) {real, imag} */,
  {32'h3fd1f656, 32'h00000000} /* (12, 4, 18) {real, imag} */,
  {32'h3fc4e340, 32'h00000000} /* (12, 4, 17) {real, imag} */,
  {32'h3f3d971b, 32'h00000000} /* (12, 4, 16) {real, imag} */,
  {32'hbf2eca60, 32'h00000000} /* (12, 4, 15) {real, imag} */,
  {32'hbf63ba49, 32'h00000000} /* (12, 4, 14) {real, imag} */,
  {32'hbf126df7, 32'h00000000} /* (12, 4, 13) {real, imag} */,
  {32'hbf327f18, 32'h00000000} /* (12, 4, 12) {real, imag} */,
  {32'hbf61e5d6, 32'h00000000} /* (12, 4, 11) {real, imag} */,
  {32'hbf77954f, 32'h00000000} /* (12, 4, 10) {real, imag} */,
  {32'hbf5e81ae, 32'h00000000} /* (12, 4, 9) {real, imag} */,
  {32'hbf5fb9cd, 32'h00000000} /* (12, 4, 8) {real, imag} */,
  {32'hbf54ac6f, 32'h00000000} /* (12, 4, 7) {real, imag} */,
  {32'hbf57bf62, 32'h00000000} /* (12, 4, 6) {real, imag} */,
  {32'h3c9cca65, 32'h00000000} /* (12, 4, 5) {real, imag} */,
  {32'h3f3d3a50, 32'h00000000} /* (12, 4, 4) {real, imag} */,
  {32'h3f438e69, 32'h00000000} /* (12, 4, 3) {real, imag} */,
  {32'h3f80b656, 32'h00000000} /* (12, 4, 2) {real, imag} */,
  {32'h3f5ac456, 32'h00000000} /* (12, 4, 1) {real, imag} */,
  {32'h3e898591, 32'h00000000} /* (12, 4, 0) {real, imag} */,
  {32'h3efac2f1, 32'h00000000} /* (12, 3, 31) {real, imag} */,
  {32'h3fa00cc1, 32'h00000000} /* (12, 3, 30) {real, imag} */,
  {32'h3fc7c220, 32'h00000000} /* (12, 3, 29) {real, imag} */,
  {32'h3f526109, 32'h00000000} /* (12, 3, 28) {real, imag} */,
  {32'h3f0913d4, 32'h00000000} /* (12, 3, 27) {real, imag} */,
  {32'h3ed073f3, 32'h00000000} /* (12, 3, 26) {real, imag} */,
  {32'h3f6c10a8, 32'h00000000} /* (12, 3, 25) {real, imag} */,
  {32'h3f86ddeb, 32'h00000000} /* (12, 3, 24) {real, imag} */,
  {32'h3fa22e94, 32'h00000000} /* (12, 3, 23) {real, imag} */,
  {32'h3fbc49f9, 32'h00000000} /* (12, 3, 22) {real, imag} */,
  {32'h3f82f60c, 32'h00000000} /* (12, 3, 21) {real, imag} */,
  {32'h3f65635c, 32'h00000000} /* (12, 3, 20) {real, imag} */,
  {32'h3f4916ef, 32'h00000000} /* (12, 3, 19) {real, imag} */,
  {32'h3f8a7da2, 32'h00000000} /* (12, 3, 18) {real, imag} */,
  {32'h3f728288, 32'h00000000} /* (12, 3, 17) {real, imag} */,
  {32'h3f0f9652, 32'h00000000} /* (12, 3, 16) {real, imag} */,
  {32'hbf2a9bba, 32'h00000000} /* (12, 3, 15) {real, imag} */,
  {32'hbf3df3c3, 32'h00000000} /* (12, 3, 14) {real, imag} */,
  {32'hbef5bf48, 32'h00000000} /* (12, 3, 13) {real, imag} */,
  {32'hbf257043, 32'h00000000} /* (12, 3, 12) {real, imag} */,
  {32'hbf60984d, 32'h00000000} /* (12, 3, 11) {real, imag} */,
  {32'hbf6d8ad8, 32'h00000000} /* (12, 3, 10) {real, imag} */,
  {32'hbf6b00be, 32'h00000000} /* (12, 3, 9) {real, imag} */,
  {32'hbf877333, 32'h00000000} /* (12, 3, 8) {real, imag} */,
  {32'hbf651c6a, 32'h00000000} /* (12, 3, 7) {real, imag} */,
  {32'hbfab9a41, 32'h00000000} /* (12, 3, 6) {real, imag} */,
  {32'h3eb0bcb8, 32'h00000000} /* (12, 3, 5) {real, imag} */,
  {32'h3fb5191f, 32'h00000000} /* (12, 3, 4) {real, imag} */,
  {32'h3eb468bf, 32'h00000000} /* (12, 3, 3) {real, imag} */,
  {32'h3f31bf53, 32'h00000000} /* (12, 3, 2) {real, imag} */,
  {32'h3f192504, 32'h00000000} /* (12, 3, 1) {real, imag} */,
  {32'h3e2e8a70, 32'h00000000} /* (12, 3, 0) {real, imag} */,
  {32'h3f31a860, 32'h00000000} /* (12, 2, 31) {real, imag} */,
  {32'h3f806efa, 32'h00000000} /* (12, 2, 30) {real, imag} */,
  {32'h3f8d4b69, 32'h00000000} /* (12, 2, 29) {real, imag} */,
  {32'h3f8577d4, 32'h00000000} /* (12, 2, 28) {real, imag} */,
  {32'h3f4160b8, 32'h00000000} /* (12, 2, 27) {real, imag} */,
  {32'h3f3a5517, 32'h00000000} /* (12, 2, 26) {real, imag} */,
  {32'h3fccd8f2, 32'h00000000} /* (12, 2, 25) {real, imag} */,
  {32'h3fef9419, 32'h00000000} /* (12, 2, 24) {real, imag} */,
  {32'h3fcaf855, 32'h00000000} /* (12, 2, 23) {real, imag} */,
  {32'h3f1a400c, 32'h00000000} /* (12, 2, 22) {real, imag} */,
  {32'h3e73d003, 32'h00000000} /* (12, 2, 21) {real, imag} */,
  {32'h3f8dcc35, 32'h00000000} /* (12, 2, 20) {real, imag} */,
  {32'h3f8b0f67, 32'h00000000} /* (12, 2, 19) {real, imag} */,
  {32'h3f8ff764, 32'h00000000} /* (12, 2, 18) {real, imag} */,
  {32'h3f206016, 32'h00000000} /* (12, 2, 17) {real, imag} */,
  {32'h3f4793a1, 32'h00000000} /* (12, 2, 16) {real, imag} */,
  {32'hbe2a4a6a, 32'h00000000} /* (12, 2, 15) {real, imag} */,
  {32'hbf4324e1, 32'h00000000} /* (12, 2, 14) {real, imag} */,
  {32'hbf8a1a16, 32'h00000000} /* (12, 2, 13) {real, imag} */,
  {32'hbf830f19, 32'h00000000} /* (12, 2, 12) {real, imag} */,
  {32'hbf16045c, 32'h00000000} /* (12, 2, 11) {real, imag} */,
  {32'hbf2e1568, 32'h00000000} /* (12, 2, 10) {real, imag} */,
  {32'hbf2c40bd, 32'h00000000} /* (12, 2, 9) {real, imag} */,
  {32'hbf920d62, 32'h00000000} /* (12, 2, 8) {real, imag} */,
  {32'hbf87f616, 32'h00000000} /* (12, 2, 7) {real, imag} */,
  {32'hbf94b61e, 32'h00000000} /* (12, 2, 6) {real, imag} */,
  {32'h3ed7b179, 32'h00000000} /* (12, 2, 5) {real, imag} */,
  {32'h3fe27051, 32'h00000000} /* (12, 2, 4) {real, imag} */,
  {32'h3f3922b9, 32'h00000000} /* (12, 2, 3) {real, imag} */,
  {32'h3f7c343f, 32'h00000000} /* (12, 2, 2) {real, imag} */,
  {32'h3f892112, 32'h00000000} /* (12, 2, 1) {real, imag} */,
  {32'h3efecef6, 32'h00000000} /* (12, 2, 0) {real, imag} */,
  {32'h3f4ddc17, 32'h00000000} /* (12, 1, 31) {real, imag} */,
  {32'h3f68c68d, 32'h00000000} /* (12, 1, 30) {real, imag} */,
  {32'h3f1ac02e, 32'h00000000} /* (12, 1, 29) {real, imag} */,
  {32'h3f19f674, 32'h00000000} /* (12, 1, 28) {real, imag} */,
  {32'h3f6ec24b, 32'h00000000} /* (12, 1, 27) {real, imag} */,
  {32'h3f47071d, 32'h00000000} /* (12, 1, 26) {real, imag} */,
  {32'h3f834d97, 32'h00000000} /* (12, 1, 25) {real, imag} */,
  {32'h3fbba4d3, 32'h00000000} /* (12, 1, 24) {real, imag} */,
  {32'h3fb7ceda, 32'h00000000} /* (12, 1, 23) {real, imag} */,
  {32'h3eb16b8a, 32'h00000000} /* (12, 1, 22) {real, imag} */,
  {32'h3f243f48, 32'h00000000} /* (12, 1, 21) {real, imag} */,
  {32'h3fb17bdf, 32'h00000000} /* (12, 1, 20) {real, imag} */,
  {32'h3f8a54ec, 32'h00000000} /* (12, 1, 19) {real, imag} */,
  {32'h3fa903ce, 32'h00000000} /* (12, 1, 18) {real, imag} */,
  {32'h3f5b6c2d, 32'h00000000} /* (12, 1, 17) {real, imag} */,
  {32'h3f391958, 32'h00000000} /* (12, 1, 16) {real, imag} */,
  {32'hbf222df7, 32'h00000000} /* (12, 1, 15) {real, imag} */,
  {32'hbfb2d932, 32'h00000000} /* (12, 1, 14) {real, imag} */,
  {32'hbf9225a3, 32'h00000000} /* (12, 1, 13) {real, imag} */,
  {32'hbf55748e, 32'h00000000} /* (12, 1, 12) {real, imag} */,
  {32'hbe2628df, 32'h00000000} /* (12, 1, 11) {real, imag} */,
  {32'hbf1a6506, 32'h00000000} /* (12, 1, 10) {real, imag} */,
  {32'hbf270d57, 32'h00000000} /* (12, 1, 9) {real, imag} */,
  {32'hbf8f2092, 32'h00000000} /* (12, 1, 8) {real, imag} */,
  {32'hbfadd2c3, 32'h00000000} /* (12, 1, 7) {real, imag} */,
  {32'hbf91df89, 32'h00000000} /* (12, 1, 6) {real, imag} */,
  {32'h3e227412, 32'h00000000} /* (12, 1, 5) {real, imag} */,
  {32'h3f85d673, 32'h00000000} /* (12, 1, 4) {real, imag} */,
  {32'h3f37d7e1, 32'h00000000} /* (12, 1, 3) {real, imag} */,
  {32'h3f29c89c, 32'h00000000} /* (12, 1, 2) {real, imag} */,
  {32'h3f9a3bc1, 32'h00000000} /* (12, 1, 1) {real, imag} */,
  {32'h3f673842, 32'h00000000} /* (12, 1, 0) {real, imag} */,
  {32'h3e9b5759, 32'h00000000} /* (12, 0, 31) {real, imag} */,
  {32'h3ef025fd, 32'h00000000} /* (12, 0, 30) {real, imag} */,
  {32'h3e89611c, 32'h00000000} /* (12, 0, 29) {real, imag} */,
  {32'h3ecf23d3, 32'h00000000} /* (12, 0, 28) {real, imag} */,
  {32'h3f21a0b4, 32'h00000000} /* (12, 0, 27) {real, imag} */,
  {32'h3f29dabe, 32'h00000000} /* (12, 0, 26) {real, imag} */,
  {32'h3ed475e6, 32'h00000000} /* (12, 0, 25) {real, imag} */,
  {32'h3f374c29, 32'h00000000} /* (12, 0, 24) {real, imag} */,
  {32'h3f88d988, 32'h00000000} /* (12, 0, 23) {real, imag} */,
  {32'h3f0c38e6, 32'h00000000} /* (12, 0, 22) {real, imag} */,
  {32'h3f185b19, 32'h00000000} /* (12, 0, 21) {real, imag} */,
  {32'h3f39692f, 32'h00000000} /* (12, 0, 20) {real, imag} */,
  {32'h3f2c8064, 32'h00000000} /* (12, 0, 19) {real, imag} */,
  {32'h3f326029, 32'h00000000} /* (12, 0, 18) {real, imag} */,
  {32'h3f0dbe8d, 32'h00000000} /* (12, 0, 17) {real, imag} */,
  {32'h3e4873cf, 32'h00000000} /* (12, 0, 16) {real, imag} */,
  {32'hbf104c32, 32'h00000000} /* (12, 0, 15) {real, imag} */,
  {32'hbf7e4fd1, 32'h00000000} /* (12, 0, 14) {real, imag} */,
  {32'hbec96f80, 32'h00000000} /* (12, 0, 13) {real, imag} */,
  {32'hbe713173, 32'h00000000} /* (12, 0, 12) {real, imag} */,
  {32'hbe3ead99, 32'h00000000} /* (12, 0, 11) {real, imag} */,
  {32'hbecafbd8, 32'h00000000} /* (12, 0, 10) {real, imag} */,
  {32'hbe3c78fa, 32'h00000000} /* (12, 0, 9) {real, imag} */,
  {32'hbeb61101, 32'h00000000} /* (12, 0, 8) {real, imag} */,
  {32'hbf05989d, 32'h00000000} /* (12, 0, 7) {real, imag} */,
  {32'hbedde569, 32'h00000000} /* (12, 0, 6) {real, imag} */,
  {32'h3e44e35c, 32'h00000000} /* (12, 0, 5) {real, imag} */,
  {32'h3f0ed0ea, 32'h00000000} /* (12, 0, 4) {real, imag} */,
  {32'h3f33c8c1, 32'h00000000} /* (12, 0, 3) {real, imag} */,
  {32'h3e9c2292, 32'h00000000} /* (12, 0, 2) {real, imag} */,
  {32'h3e9d0efa, 32'h00000000} /* (12, 0, 1) {real, imag} */,
  {32'h3ee55e1e, 32'h00000000} /* (12, 0, 0) {real, imag} */,
  {32'h3e4405da, 32'h00000000} /* (11, 31, 31) {real, imag} */,
  {32'h3eae6d09, 32'h00000000} /* (11, 31, 30) {real, imag} */,
  {32'h3ea76462, 32'h00000000} /* (11, 31, 29) {real, imag} */,
  {32'h3ec01762, 32'h00000000} /* (11, 31, 28) {real, imag} */,
  {32'h3f3710a1, 32'h00000000} /* (11, 31, 27) {real, imag} */,
  {32'h3f45ecf7, 32'h00000000} /* (11, 31, 26) {real, imag} */,
  {32'h3f199be7, 32'h00000000} /* (11, 31, 25) {real, imag} */,
  {32'h3f3329e4, 32'h00000000} /* (11, 31, 24) {real, imag} */,
  {32'h3f3f56bd, 32'h00000000} /* (11, 31, 23) {real, imag} */,
  {32'h3f337d5e, 32'h00000000} /* (11, 31, 22) {real, imag} */,
  {32'h3e8172b0, 32'h00000000} /* (11, 31, 21) {real, imag} */,
  {32'hbed9f081, 32'h00000000} /* (11, 31, 20) {real, imag} */,
  {32'hbecddfaf, 32'h00000000} /* (11, 31, 19) {real, imag} */,
  {32'hbe9be921, 32'h00000000} /* (11, 31, 18) {real, imag} */,
  {32'hbef11de2, 32'h00000000} /* (11, 31, 17) {real, imag} */,
  {32'hbf568f88, 32'h00000000} /* (11, 31, 16) {real, imag} */,
  {32'hbf6abf6d, 32'h00000000} /* (11, 31, 15) {real, imag} */,
  {32'hbf15f6d9, 32'h00000000} /* (11, 31, 14) {real, imag} */,
  {32'hbf4a8db0, 32'h00000000} /* (11, 31, 13) {real, imag} */,
  {32'hbf4bfe2f, 32'h00000000} /* (11, 31, 12) {real, imag} */,
  {32'hbf6992e5, 32'h00000000} /* (11, 31, 11) {real, imag} */,
  {32'h3ee1f9b3, 32'h00000000} /* (11, 31, 10) {real, imag} */,
  {32'h3f05c197, 32'h00000000} /* (11, 31, 9) {real, imag} */,
  {32'h3e9a49e6, 32'h00000000} /* (11, 31, 8) {real, imag} */,
  {32'h3e9a40b3, 32'h00000000} /* (11, 31, 7) {real, imag} */,
  {32'h3f21dece, 32'h00000000} /* (11, 31, 6) {real, imag} */,
  {32'h3f3876fa, 32'h00000000} /* (11, 31, 5) {real, imag} */,
  {32'h3f526f5b, 32'h00000000} /* (11, 31, 4) {real, imag} */,
  {32'h3f3646cc, 32'h00000000} /* (11, 31, 3) {real, imag} */,
  {32'h3f7da86d, 32'h00000000} /* (11, 31, 2) {real, imag} */,
  {32'h3ed8d5d6, 32'h00000000} /* (11, 31, 1) {real, imag} */,
  {32'h3f1a5a81, 32'h00000000} /* (11, 31, 0) {real, imag} */,
  {32'h3f094b4c, 32'h00000000} /* (11, 30, 31) {real, imag} */,
  {32'h3f0a4189, 32'h00000000} /* (11, 30, 30) {real, imag} */,
  {32'h3e27a829, 32'h00000000} /* (11, 30, 29) {real, imag} */,
  {32'h3ef8a35d, 32'h00000000} /* (11, 30, 28) {real, imag} */,
  {32'h3f144d2a, 32'h00000000} /* (11, 30, 27) {real, imag} */,
  {32'h3f5b8321, 32'h00000000} /* (11, 30, 26) {real, imag} */,
  {32'h3f88a8b5, 32'h00000000} /* (11, 30, 25) {real, imag} */,
  {32'h3fa4f0e6, 32'h00000000} /* (11, 30, 24) {real, imag} */,
  {32'h3f7431c2, 32'h00000000} /* (11, 30, 23) {real, imag} */,
  {32'h3f1fc2c8, 32'h00000000} /* (11, 30, 22) {real, imag} */,
  {32'h3e8cc6fa, 32'h00000000} /* (11, 30, 21) {real, imag} */,
  {32'hbe370981, 32'h00000000} /* (11, 30, 20) {real, imag} */,
  {32'hbef46111, 32'h00000000} /* (11, 30, 19) {real, imag} */,
  {32'hbf449745, 32'h00000000} /* (11, 30, 18) {real, imag} */,
  {32'hbf810432, 32'h00000000} /* (11, 30, 17) {real, imag} */,
  {32'hbf6cb1d6, 32'h00000000} /* (11, 30, 16) {real, imag} */,
  {32'hbf8abea6, 32'h00000000} /* (11, 30, 15) {real, imag} */,
  {32'hbf935b87, 32'h00000000} /* (11, 30, 14) {real, imag} */,
  {32'hbf87f3e1, 32'h00000000} /* (11, 30, 13) {real, imag} */,
  {32'hbf85910f, 32'h00000000} /* (11, 30, 12) {real, imag} */,
  {32'hbee77343, 32'h00000000} /* (11, 30, 11) {real, imag} */,
  {32'h3f99cfa1, 32'h00000000} /* (11, 30, 10) {real, imag} */,
  {32'h3f869a38, 32'h00000000} /* (11, 30, 9) {real, imag} */,
  {32'h3f365bb3, 32'h00000000} /* (11, 30, 8) {real, imag} */,
  {32'h3f4ce620, 32'h00000000} /* (11, 30, 7) {real, imag} */,
  {32'h3f8c8787, 32'h00000000} /* (11, 30, 6) {real, imag} */,
  {32'h3fb708ef, 32'h00000000} /* (11, 30, 5) {real, imag} */,
  {32'h3fde3c4f, 32'h00000000} /* (11, 30, 4) {real, imag} */,
  {32'h3f95e7d9, 32'h00000000} /* (11, 30, 3) {real, imag} */,
  {32'h3f93767a, 32'h00000000} /* (11, 30, 2) {real, imag} */,
  {32'h3ecb4e65, 32'h00000000} /* (11, 30, 1) {real, imag} */,
  {32'h3ea306c9, 32'h00000000} /* (11, 30, 0) {real, imag} */,
  {32'h3f208417, 32'h00000000} /* (11, 29, 31) {real, imag} */,
  {32'h3f868566, 32'h00000000} /* (11, 29, 30) {real, imag} */,
  {32'h3f2f4ce6, 32'h00000000} /* (11, 29, 29) {real, imag} */,
  {32'h3f170691, 32'h00000000} /* (11, 29, 28) {real, imag} */,
  {32'h3eaeb64c, 32'h00000000} /* (11, 29, 27) {real, imag} */,
  {32'h3f327e3c, 32'h00000000} /* (11, 29, 26) {real, imag} */,
  {32'h3f4ea7c2, 32'h00000000} /* (11, 29, 25) {real, imag} */,
  {32'h3f67ddf1, 32'h00000000} /* (11, 29, 24) {real, imag} */,
  {32'h3f91a01b, 32'h00000000} /* (11, 29, 23) {real, imag} */,
  {32'h3f5c99d8, 32'h00000000} /* (11, 29, 22) {real, imag} */,
  {32'h3ebd0f64, 32'h00000000} /* (11, 29, 21) {real, imag} */,
  {32'hbe9c8e79, 32'h00000000} /* (11, 29, 20) {real, imag} */,
  {32'hbf1f9010, 32'h00000000} /* (11, 29, 19) {real, imag} */,
  {32'hbf6bcd4c, 32'h00000000} /* (11, 29, 18) {real, imag} */,
  {32'hbf37d0be, 32'h00000000} /* (11, 29, 17) {real, imag} */,
  {32'hbeee3591, 32'h00000000} /* (11, 29, 16) {real, imag} */,
  {32'hbf47c4ad, 32'h00000000} /* (11, 29, 15) {real, imag} */,
  {32'hbf6cfdc6, 32'h00000000} /* (11, 29, 14) {real, imag} */,
  {32'hbf842777, 32'h00000000} /* (11, 29, 13) {real, imag} */,
  {32'hbf80fd8b, 32'h00000000} /* (11, 29, 12) {real, imag} */,
  {32'hbe5d81cf, 32'h00000000} /* (11, 29, 11) {real, imag} */,
  {32'h3f4302ba, 32'h00000000} /* (11, 29, 10) {real, imag} */,
  {32'h3f546c99, 32'h00000000} /* (11, 29, 9) {real, imag} */,
  {32'h3f42ab1c, 32'h00000000} /* (11, 29, 8) {real, imag} */,
  {32'h3f4098c7, 32'h00000000} /* (11, 29, 7) {real, imag} */,
  {32'h3f88315c, 32'h00000000} /* (11, 29, 6) {real, imag} */,
  {32'h3f6a2bb7, 32'h00000000} /* (11, 29, 5) {real, imag} */,
  {32'h3f8eff81, 32'h00000000} /* (11, 29, 4) {real, imag} */,
  {32'h3f812cb2, 32'h00000000} /* (11, 29, 3) {real, imag} */,
  {32'h3f59314b, 32'h00000000} /* (11, 29, 2) {real, imag} */,
  {32'h3f45c8ee, 32'h00000000} /* (11, 29, 1) {real, imag} */,
  {32'h3ec263f7, 32'h00000000} /* (11, 29, 0) {real, imag} */,
  {32'h3ee646dd, 32'h00000000} /* (11, 28, 31) {real, imag} */,
  {32'h3f8bbef3, 32'h00000000} /* (11, 28, 30) {real, imag} */,
  {32'h3f8bbf2f, 32'h00000000} /* (11, 28, 29) {real, imag} */,
  {32'h3f281767, 32'h00000000} /* (11, 28, 28) {real, imag} */,
  {32'h3f5ff8ec, 32'h00000000} /* (11, 28, 27) {real, imag} */,
  {32'h3f9c8ff7, 32'h00000000} /* (11, 28, 26) {real, imag} */,
  {32'h3f51498e, 32'h00000000} /* (11, 28, 25) {real, imag} */,
  {32'h3f225093, 32'h00000000} /* (11, 28, 24) {real, imag} */,
  {32'h3fb721bc, 32'h00000000} /* (11, 28, 23) {real, imag} */,
  {32'h3fa0f7f9, 32'h00000000} /* (11, 28, 22) {real, imag} */,
  {32'h3ec404e6, 32'h00000000} /* (11, 28, 21) {real, imag} */,
  {32'hbf79443e, 32'h00000000} /* (11, 28, 20) {real, imag} */,
  {32'hbf839b6f, 32'h00000000} /* (11, 28, 19) {real, imag} */,
  {32'hbf9b104c, 32'h00000000} /* (11, 28, 18) {real, imag} */,
  {32'hbf92fefe, 32'h00000000} /* (11, 28, 17) {real, imag} */,
  {32'hbf88e39e, 32'h00000000} /* (11, 28, 16) {real, imag} */,
  {32'hbf91fc9b, 32'h00000000} /* (11, 28, 15) {real, imag} */,
  {32'hbf508713, 32'h00000000} /* (11, 28, 14) {real, imag} */,
  {32'hbf49b2e0, 32'h00000000} /* (11, 28, 13) {real, imag} */,
  {32'hbf51c1bc, 32'h00000000} /* (11, 28, 12) {real, imag} */,
  {32'hbe549add, 32'h00000000} /* (11, 28, 11) {real, imag} */,
  {32'h3d8bb380, 32'h00000000} /* (11, 28, 10) {real, imag} */,
  {32'h3f0763bf, 32'h00000000} /* (11, 28, 9) {real, imag} */,
  {32'h3f277f60, 32'h00000000} /* (11, 28, 8) {real, imag} */,
  {32'h3f0a3254, 32'h00000000} /* (11, 28, 7) {real, imag} */,
  {32'h3f8685fe, 32'h00000000} /* (11, 28, 6) {real, imag} */,
  {32'h3f50ffcb, 32'h00000000} /* (11, 28, 5) {real, imag} */,
  {32'h3f9e8330, 32'h00000000} /* (11, 28, 4) {real, imag} */,
  {32'h3f6ff168, 32'h00000000} /* (11, 28, 3) {real, imag} */,
  {32'h3f8acf48, 32'h00000000} /* (11, 28, 2) {real, imag} */,
  {32'h3f903d8e, 32'h00000000} /* (11, 28, 1) {real, imag} */,
  {32'h3ee6cfc5, 32'h00000000} /* (11, 28, 0) {real, imag} */,
  {32'h3f2f9311, 32'h00000000} /* (11, 27, 31) {real, imag} */,
  {32'h3fa94c90, 32'h00000000} /* (11, 27, 30) {real, imag} */,
  {32'h3fda0284, 32'h00000000} /* (11, 27, 29) {real, imag} */,
  {32'h3f6ff9f2, 32'h00000000} /* (11, 27, 28) {real, imag} */,
  {32'h3f8196aa, 32'h00000000} /* (11, 27, 27) {real, imag} */,
  {32'h3fc6aee3, 32'h00000000} /* (11, 27, 26) {real, imag} */,
  {32'h3f8d57a0, 32'h00000000} /* (11, 27, 25) {real, imag} */,
  {32'h3f547aa9, 32'h00000000} /* (11, 27, 24) {real, imag} */,
  {32'h3fe421f5, 32'h00000000} /* (11, 27, 23) {real, imag} */,
  {32'h3fb61833, 32'h00000000} /* (11, 27, 22) {real, imag} */,
  {32'h3dd420ac, 32'h00000000} /* (11, 27, 21) {real, imag} */,
  {32'hbf78d5f4, 32'h00000000} /* (11, 27, 20) {real, imag} */,
  {32'hbfb8719c, 32'h00000000} /* (11, 27, 19) {real, imag} */,
  {32'hbfb06ede, 32'h00000000} /* (11, 27, 18) {real, imag} */,
  {32'hbf931954, 32'h00000000} /* (11, 27, 17) {real, imag} */,
  {32'hbfaa4228, 32'h00000000} /* (11, 27, 16) {real, imag} */,
  {32'hbfad6138, 32'h00000000} /* (11, 27, 15) {real, imag} */,
  {32'hbf996547, 32'h00000000} /* (11, 27, 14) {real, imag} */,
  {32'hbecdc410, 32'h00000000} /* (11, 27, 13) {real, imag} */,
  {32'hbef8674b, 32'h00000000} /* (11, 27, 12) {real, imag} */,
  {32'hbf388a6f, 32'h00000000} /* (11, 27, 11) {real, imag} */,
  {32'hbe685be3, 32'h00000000} /* (11, 27, 10) {real, imag} */,
  {32'h3ef2d2f7, 32'h00000000} /* (11, 27, 9) {real, imag} */,
  {32'h3f52de24, 32'h00000000} /* (11, 27, 8) {real, imag} */,
  {32'h3f83932e, 32'h00000000} /* (11, 27, 7) {real, imag} */,
  {32'h3fa2acde, 32'h00000000} /* (11, 27, 6) {real, imag} */,
  {32'h3f68d5fc, 32'h00000000} /* (11, 27, 5) {real, imag} */,
  {32'h3fb5f331, 32'h00000000} /* (11, 27, 4) {real, imag} */,
  {32'h3f57aac8, 32'h00000000} /* (11, 27, 3) {real, imag} */,
  {32'h3f305cc0, 32'h00000000} /* (11, 27, 2) {real, imag} */,
  {32'h3f6a4a8b, 32'h00000000} /* (11, 27, 1) {real, imag} */,
  {32'h3f429df8, 32'h00000000} /* (11, 27, 0) {real, imag} */,
  {32'h3f12a836, 32'h00000000} /* (11, 26, 31) {real, imag} */,
  {32'h3fabbaaf, 32'h00000000} /* (11, 26, 30) {real, imag} */,
  {32'h3fd2d58f, 32'h00000000} /* (11, 26, 29) {real, imag} */,
  {32'h3f814c79, 32'h00000000} /* (11, 26, 28) {real, imag} */,
  {32'h3f875c9c, 32'h00000000} /* (11, 26, 27) {real, imag} */,
  {32'h3f7632b0, 32'h00000000} /* (11, 26, 26) {real, imag} */,
  {32'h3fafcfa9, 32'h00000000} /* (11, 26, 25) {real, imag} */,
  {32'h3f937861, 32'h00000000} /* (11, 26, 24) {real, imag} */,
  {32'h3f8c4fe3, 32'h00000000} /* (11, 26, 23) {real, imag} */,
  {32'h3f7c6a4e, 32'h00000000} /* (11, 26, 22) {real, imag} */,
  {32'h3dc90255, 32'h00000000} /* (11, 26, 21) {real, imag} */,
  {32'hbf08d2f0, 32'h00000000} /* (11, 26, 20) {real, imag} */,
  {32'hbf58c630, 32'h00000000} /* (11, 26, 19) {real, imag} */,
  {32'hbf39d1bd, 32'h00000000} /* (11, 26, 18) {real, imag} */,
  {32'hbf840b9a, 32'h00000000} /* (11, 26, 17) {real, imag} */,
  {32'hbfbfc0ad, 32'h00000000} /* (11, 26, 16) {real, imag} */,
  {32'hbfb09cb6, 32'h00000000} /* (11, 26, 15) {real, imag} */,
  {32'hbf9a6df1, 32'h00000000} /* (11, 26, 14) {real, imag} */,
  {32'hbf2e236b, 32'h00000000} /* (11, 26, 13) {real, imag} */,
  {32'hbf1957ff, 32'h00000000} /* (11, 26, 12) {real, imag} */,
  {32'hbf10b015, 32'h00000000} /* (11, 26, 11) {real, imag} */,
  {32'h3dc52c7e, 32'h00000000} /* (11, 26, 10) {real, imag} */,
  {32'h3f7ced15, 32'h00000000} /* (11, 26, 9) {real, imag} */,
  {32'h3f992915, 32'h00000000} /* (11, 26, 8) {real, imag} */,
  {32'h3f8081c9, 32'h00000000} /* (11, 26, 7) {real, imag} */,
  {32'h3f11d92e, 32'h00000000} /* (11, 26, 6) {real, imag} */,
  {32'h3f2eeb66, 32'h00000000} /* (11, 26, 5) {real, imag} */,
  {32'h3f77a9bc, 32'h00000000} /* (11, 26, 4) {real, imag} */,
  {32'h3f5dd878, 32'h00000000} /* (11, 26, 3) {real, imag} */,
  {32'h3f50c63e, 32'h00000000} /* (11, 26, 2) {real, imag} */,
  {32'h3f686275, 32'h00000000} /* (11, 26, 1) {real, imag} */,
  {32'h3f67d1f9, 32'h00000000} /* (11, 26, 0) {real, imag} */,
  {32'h3e77deeb, 32'h00000000} /* (11, 25, 31) {real, imag} */,
  {32'h3f398f0d, 32'h00000000} /* (11, 25, 30) {real, imag} */,
  {32'h3f90e3a9, 32'h00000000} /* (11, 25, 29) {real, imag} */,
  {32'h3fa409ab, 32'h00000000} /* (11, 25, 28) {real, imag} */,
  {32'h3f6dd3e0, 32'h00000000} /* (11, 25, 27) {real, imag} */,
  {32'h3f1f3355, 32'h00000000} /* (11, 25, 26) {real, imag} */,
  {32'h3fe2efe0, 32'h00000000} /* (11, 25, 25) {real, imag} */,
  {32'h3f9bf60d, 32'h00000000} /* (11, 25, 24) {real, imag} */,
  {32'h3f04f172, 32'h00000000} /* (11, 25, 23) {real, imag} */,
  {32'h3f48731b, 32'h00000000} /* (11, 25, 22) {real, imag} */,
  {32'h3e4ce0d9, 32'h00000000} /* (11, 25, 21) {real, imag} */,
  {32'hbed20dc9, 32'h00000000} /* (11, 25, 20) {real, imag} */,
  {32'hbf182e15, 32'h00000000} /* (11, 25, 19) {real, imag} */,
  {32'hbf900404, 32'h00000000} /* (11, 25, 18) {real, imag} */,
  {32'hc007414a, 32'h00000000} /* (11, 25, 17) {real, imag} */,
  {32'hbfeeb34a, 32'h00000000} /* (11, 25, 16) {real, imag} */,
  {32'hbf31e91b, 32'h00000000} /* (11, 25, 15) {real, imag} */,
  {32'hbe595cbd, 32'h00000000} /* (11, 25, 14) {real, imag} */,
  {32'hbef090d4, 32'h00000000} /* (11, 25, 13) {real, imag} */,
  {32'hbf85f71a, 32'h00000000} /* (11, 25, 12) {real, imag} */,
  {32'hbf2227f2, 32'h00000000} /* (11, 25, 11) {real, imag} */,
  {32'h3e62cd5a, 32'h00000000} /* (11, 25, 10) {real, imag} */,
  {32'h3fa5ade7, 32'h00000000} /* (11, 25, 9) {real, imag} */,
  {32'h3fb7a590, 32'h00000000} /* (11, 25, 8) {real, imag} */,
  {32'h3f92691a, 32'h00000000} /* (11, 25, 7) {real, imag} */,
  {32'h3f3c6f02, 32'h00000000} /* (11, 25, 6) {real, imag} */,
  {32'h3f951e6a, 32'h00000000} /* (11, 25, 5) {real, imag} */,
  {32'h3fb8dd64, 32'h00000000} /* (11, 25, 4) {real, imag} */,
  {32'h3f9ccccb, 32'h00000000} /* (11, 25, 3) {real, imag} */,
  {32'h3f8de4e2, 32'h00000000} /* (11, 25, 2) {real, imag} */,
  {32'h3f16040a, 32'h00000000} /* (11, 25, 1) {real, imag} */,
  {32'h3e868771, 32'h00000000} /* (11, 25, 0) {real, imag} */,
  {32'h3e5340f6, 32'h00000000} /* (11, 24, 31) {real, imag} */,
  {32'h3f22e754, 32'h00000000} /* (11, 24, 30) {real, imag} */,
  {32'h3f54bd11, 32'h00000000} /* (11, 24, 29) {real, imag} */,
  {32'h3f974a0d, 32'h00000000} /* (11, 24, 28) {real, imag} */,
  {32'h3f9e1186, 32'h00000000} /* (11, 24, 27) {real, imag} */,
  {32'h3f304875, 32'h00000000} /* (11, 24, 26) {real, imag} */,
  {32'h3f9ae88d, 32'h00000000} /* (11, 24, 25) {real, imag} */,
  {32'h3f7f95e2, 32'h00000000} /* (11, 24, 24) {real, imag} */,
  {32'h3ec48a08, 32'h00000000} /* (11, 24, 23) {real, imag} */,
  {32'h3ef84eef, 32'h00000000} /* (11, 24, 22) {real, imag} */,
  {32'hbe2ff21f, 32'h00000000} /* (11, 24, 21) {real, imag} */,
  {32'hbfb8baf0, 32'h00000000} /* (11, 24, 20) {real, imag} */,
  {32'hbfa0695f, 32'h00000000} /* (11, 24, 19) {real, imag} */,
  {32'hbfc2afd4, 32'h00000000} /* (11, 24, 18) {real, imag} */,
  {32'hc005eed4, 32'h00000000} /* (11, 24, 17) {real, imag} */,
  {32'hbf85de0f, 32'h00000000} /* (11, 24, 16) {real, imag} */,
  {32'hbeef1f55, 32'h00000000} /* (11, 24, 15) {real, imag} */,
  {32'hbd8676a0, 32'h00000000} /* (11, 24, 14) {real, imag} */,
  {32'hbed1ed04, 32'h00000000} /* (11, 24, 13) {real, imag} */,
  {32'hbf5c37d5, 32'h00000000} /* (11, 24, 12) {real, imag} */,
  {32'hbe6ba921, 32'h00000000} /* (11, 24, 11) {real, imag} */,
  {32'h3f4201a8, 32'h00000000} /* (11, 24, 10) {real, imag} */,
  {32'h3fe0f5eb, 32'h00000000} /* (11, 24, 9) {real, imag} */,
  {32'h3fb16bbe, 32'h00000000} /* (11, 24, 8) {real, imag} */,
  {32'h3fc5a738, 32'h00000000} /* (11, 24, 7) {real, imag} */,
  {32'h3f9e5720, 32'h00000000} /* (11, 24, 6) {real, imag} */,
  {32'h3f7fd6aa, 32'h00000000} /* (11, 24, 5) {real, imag} */,
  {32'h3fa7400f, 32'h00000000} /* (11, 24, 4) {real, imag} */,
  {32'h3fd06451, 32'h00000000} /* (11, 24, 3) {real, imag} */,
  {32'h3f9f9751, 32'h00000000} /* (11, 24, 2) {real, imag} */,
  {32'h3ee7a59a, 32'h00000000} /* (11, 24, 1) {real, imag} */,
  {32'h3dc8c202, 32'h00000000} /* (11, 24, 0) {real, imag} */,
  {32'h3ee41de2, 32'h00000000} /* (11, 23, 31) {real, imag} */,
  {32'h3f85e3bb, 32'h00000000} /* (11, 23, 30) {real, imag} */,
  {32'h3f75450f, 32'h00000000} /* (11, 23, 29) {real, imag} */,
  {32'h3f5df6bf, 32'h00000000} /* (11, 23, 28) {real, imag} */,
  {32'h3f8067db, 32'h00000000} /* (11, 23, 27) {real, imag} */,
  {32'h3f53b13d, 32'h00000000} /* (11, 23, 26) {real, imag} */,
  {32'h3f16abbe, 32'h00000000} /* (11, 23, 25) {real, imag} */,
  {32'h3f280fa8, 32'h00000000} /* (11, 23, 24) {real, imag} */,
  {32'h3f138615, 32'h00000000} /* (11, 23, 23) {real, imag} */,
  {32'h3edf2c68, 32'h00000000} /* (11, 23, 22) {real, imag} */,
  {32'h3db0896e, 32'h00000000} /* (11, 23, 21) {real, imag} */,
  {32'hbfb1a5d7, 32'h00000000} /* (11, 23, 20) {real, imag} */,
  {32'hbfdef30b, 32'h00000000} /* (11, 23, 19) {real, imag} */,
  {32'hbfc92039, 32'h00000000} /* (11, 23, 18) {real, imag} */,
  {32'hbfb89e40, 32'h00000000} /* (11, 23, 17) {real, imag} */,
  {32'hbf5dfc99, 32'h00000000} /* (11, 23, 16) {real, imag} */,
  {32'hbeef5486, 32'h00000000} /* (11, 23, 15) {real, imag} */,
  {32'hbeca0d55, 32'h00000000} /* (11, 23, 14) {real, imag} */,
  {32'hbeeeacb5, 32'h00000000} /* (11, 23, 13) {real, imag} */,
  {32'hbf1e17f8, 32'h00000000} /* (11, 23, 12) {real, imag} */,
  {32'hbf114b49, 32'h00000000} /* (11, 23, 11) {real, imag} */,
  {32'h3ee5f013, 32'h00000000} /* (11, 23, 10) {real, imag} */,
  {32'h3fc5aa1e, 32'h00000000} /* (11, 23, 9) {real, imag} */,
  {32'h3f8a9cbc, 32'h00000000} /* (11, 23, 8) {real, imag} */,
  {32'h3f92d3c9, 32'h00000000} /* (11, 23, 7) {real, imag} */,
  {32'h3f91f8b2, 32'h00000000} /* (11, 23, 6) {real, imag} */,
  {32'h3f4e6e24, 32'h00000000} /* (11, 23, 5) {real, imag} */,
  {32'h3f8d21a1, 32'h00000000} /* (11, 23, 4) {real, imag} */,
  {32'h3f9dad5a, 32'h00000000} /* (11, 23, 3) {real, imag} */,
  {32'h3f55e322, 32'h00000000} /* (11, 23, 2) {real, imag} */,
  {32'h3f81271a, 32'h00000000} /* (11, 23, 1) {real, imag} */,
  {32'h3f11ccfe, 32'h00000000} /* (11, 23, 0) {real, imag} */,
  {32'h3ecf9537, 32'h00000000} /* (11, 22, 31) {real, imag} */,
  {32'h3f93b322, 32'h00000000} /* (11, 22, 30) {real, imag} */,
  {32'h3f8bfcce, 32'h00000000} /* (11, 22, 29) {real, imag} */,
  {32'h3f80555b, 32'h00000000} /* (11, 22, 28) {real, imag} */,
  {32'h3f25775a, 32'h00000000} /* (11, 22, 27) {real, imag} */,
  {32'h3f228f65, 32'h00000000} /* (11, 22, 26) {real, imag} */,
  {32'h3f0940d2, 32'h00000000} /* (11, 22, 25) {real, imag} */,
  {32'h3f295e1c, 32'h00000000} /* (11, 22, 24) {real, imag} */,
  {32'h3f81006e, 32'h00000000} /* (11, 22, 23) {real, imag} */,
  {32'h3f5585da, 32'h00000000} /* (11, 22, 22) {real, imag} */,
  {32'h3e6df42e, 32'h00000000} /* (11, 22, 21) {real, imag} */,
  {32'hbf997d3a, 32'h00000000} /* (11, 22, 20) {real, imag} */,
  {32'hbfd01e6a, 32'h00000000} /* (11, 22, 19) {real, imag} */,
  {32'hbf94be83, 32'h00000000} /* (11, 22, 18) {real, imag} */,
  {32'hbf75dfc5, 32'h00000000} /* (11, 22, 17) {real, imag} */,
  {32'hbf9d3e93, 32'h00000000} /* (11, 22, 16) {real, imag} */,
  {32'hbf238458, 32'h00000000} /* (11, 22, 15) {real, imag} */,
  {32'hbf3b6d6b, 32'h00000000} /* (11, 22, 14) {real, imag} */,
  {32'hbf6324bc, 32'h00000000} /* (11, 22, 13) {real, imag} */,
  {32'hbf8703d4, 32'h00000000} /* (11, 22, 12) {real, imag} */,
  {32'hbf9567ca, 32'h00000000} /* (11, 22, 11) {real, imag} */,
  {32'h3dcfb35a, 32'h00000000} /* (11, 22, 10) {real, imag} */,
  {32'h3f9080bf, 32'h00000000} /* (11, 22, 9) {real, imag} */,
  {32'h3f7e3e75, 32'h00000000} /* (11, 22, 8) {real, imag} */,
  {32'h3f46ad0f, 32'h00000000} /* (11, 22, 7) {real, imag} */,
  {32'h3f4c7a9a, 32'h00000000} /* (11, 22, 6) {real, imag} */,
  {32'h3edcfcbe, 32'h00000000} /* (11, 22, 5) {real, imag} */,
  {32'h3efd41b2, 32'h00000000} /* (11, 22, 4) {real, imag} */,
  {32'h3f252d4d, 32'h00000000} /* (11, 22, 3) {real, imag} */,
  {32'h3f84282f, 32'h00000000} /* (11, 22, 2) {real, imag} */,
  {32'h3fc6f710, 32'h00000000} /* (11, 22, 1) {real, imag} */,
  {32'h3f664b77, 32'h00000000} /* (11, 22, 0) {real, imag} */,
  {32'h3e3c634a, 32'h00000000} /* (11, 21, 31) {real, imag} */,
  {32'h3ed50935, 32'h00000000} /* (11, 21, 30) {real, imag} */,
  {32'h3f52ab89, 32'h00000000} /* (11, 21, 29) {real, imag} */,
  {32'h3fa029df, 32'h00000000} /* (11, 21, 28) {real, imag} */,
  {32'h3f04c932, 32'h00000000} /* (11, 21, 27) {real, imag} */,
  {32'h3e8ab7a5, 32'h00000000} /* (11, 21, 26) {real, imag} */,
  {32'h3e9fa7c9, 32'h00000000} /* (11, 21, 25) {real, imag} */,
  {32'h3ec543ff, 32'h00000000} /* (11, 21, 24) {real, imag} */,
  {32'h3d00ec38, 32'h00000000} /* (11, 21, 23) {real, imag} */,
  {32'h3d839d39, 32'h00000000} /* (11, 21, 22) {real, imag} */,
  {32'h3e86ad5c, 32'h00000000} /* (11, 21, 21) {real, imag} */,
  {32'hbf077034, 32'h00000000} /* (11, 21, 20) {real, imag} */,
  {32'hbf38ec54, 32'h00000000} /* (11, 21, 19) {real, imag} */,
  {32'hbeff1bf7, 32'h00000000} /* (11, 21, 18) {real, imag} */,
  {32'hbedb1eab, 32'h00000000} /* (11, 21, 17) {real, imag} */,
  {32'hbeb6bdd0, 32'h00000000} /* (11, 21, 16) {real, imag} */,
  {32'hbd848be5, 32'h00000000} /* (11, 21, 15) {real, imag} */,
  {32'hbf09fa30, 32'h00000000} /* (11, 21, 14) {real, imag} */,
  {32'hbf3486d0, 32'h00000000} /* (11, 21, 13) {real, imag} */,
  {32'hbe3e8a21, 32'h00000000} /* (11, 21, 12) {real, imag} */,
  {32'hbe66702c, 32'h00000000} /* (11, 21, 11) {real, imag} */,
  {32'hbd5b3922, 32'h00000000} /* (11, 21, 10) {real, imag} */,
  {32'h3e12060e, 32'h00000000} /* (11, 21, 9) {real, imag} */,
  {32'h3cf86ec2, 32'h00000000} /* (11, 21, 8) {real, imag} */,
  {32'h3c78ba49, 32'h00000000} /* (11, 21, 7) {real, imag} */,
  {32'h3ec3bd97, 32'h00000000} /* (11, 21, 6) {real, imag} */,
  {32'h3eade0f7, 32'h00000000} /* (11, 21, 5) {real, imag} */,
  {32'h3eee95a9, 32'h00000000} /* (11, 21, 4) {real, imag} */,
  {32'h3efa8096, 32'h00000000} /* (11, 21, 3) {real, imag} */,
  {32'h3f06d48a, 32'h00000000} /* (11, 21, 2) {real, imag} */,
  {32'h3f405cf0, 32'h00000000} /* (11, 21, 1) {real, imag} */,
  {32'h3eb5756f, 32'h00000000} /* (11, 21, 0) {real, imag} */,
  {32'hbe3172e3, 32'h00000000} /* (11, 20, 31) {real, imag} */,
  {32'hbf7e07a0, 32'h00000000} /* (11, 20, 30) {real, imag} */,
  {32'hbf1c67e8, 32'h00000000} /* (11, 20, 29) {real, imag} */,
  {32'hbc18dac8, 32'h00000000} /* (11, 20, 28) {real, imag} */,
  {32'h3e0d8886, 32'h00000000} /* (11, 20, 27) {real, imag} */,
  {32'h3d40f050, 32'h00000000} /* (11, 20, 26) {real, imag} */,
  {32'hbf2b9cc6, 32'h00000000} /* (11, 20, 25) {real, imag} */,
  {32'hbf6fcb74, 32'h00000000} /* (11, 20, 24) {real, imag} */,
  {32'hbf298486, 32'h00000000} /* (11, 20, 23) {real, imag} */,
  {32'hbf89696a, 32'h00000000} /* (11, 20, 22) {real, imag} */,
  {32'hbed5e6c9, 32'h00000000} /* (11, 20, 21) {real, imag} */,
  {32'h3e376c2b, 32'h00000000} /* (11, 20, 20) {real, imag} */,
  {32'h3f02d04b, 32'h00000000} /* (11, 20, 19) {real, imag} */,
  {32'h3f36b544, 32'h00000000} /* (11, 20, 18) {real, imag} */,
  {32'h3f5a78e1, 32'h00000000} /* (11, 20, 17) {real, imag} */,
  {32'h3f911a6f, 32'h00000000} /* (11, 20, 16) {real, imag} */,
  {32'h3f9646ff, 32'h00000000} /* (11, 20, 15) {real, imag} */,
  {32'h3f00e1ef, 32'h00000000} /* (11, 20, 14) {real, imag} */,
  {32'h3ed0717c, 32'h00000000} /* (11, 20, 13) {real, imag} */,
  {32'h3f743268, 32'h00000000} /* (11, 20, 12) {real, imag} */,
  {32'h3f1372a7, 32'h00000000} /* (11, 20, 11) {real, imag} */,
  {32'hbf38dfb1, 32'h00000000} /* (11, 20, 10) {real, imag} */,
  {32'hbf4ee677, 32'h00000000} /* (11, 20, 9) {real, imag} */,
  {32'hbf144347, 32'h00000000} /* (11, 20, 8) {real, imag} */,
  {32'hbf20d629, 32'h00000000} /* (11, 20, 7) {real, imag} */,
  {32'hbf174bde, 32'h00000000} /* (11, 20, 6) {real, imag} */,
  {32'hbf62efb7, 32'h00000000} /* (11, 20, 5) {real, imag} */,
  {32'hbed6fed3, 32'h00000000} /* (11, 20, 4) {real, imag} */,
  {32'hbeb79c85, 32'h00000000} /* (11, 20, 3) {real, imag} */,
  {32'hbf3f5d92, 32'h00000000} /* (11, 20, 2) {real, imag} */,
  {32'hbf5d9c21, 32'h00000000} /* (11, 20, 1) {real, imag} */,
  {32'hbe87c8f5, 32'h00000000} /* (11, 20, 0) {real, imag} */,
  {32'hbe9cdd7d, 32'h00000000} /* (11, 19, 31) {real, imag} */,
  {32'hbfb2fd76, 32'h00000000} /* (11, 19, 30) {real, imag} */,
  {32'hbfa9c00a, 32'h00000000} /* (11, 19, 29) {real, imag} */,
  {32'hbf2f178b, 32'h00000000} /* (11, 19, 28) {real, imag} */,
  {32'hbeb9deb0, 32'h00000000} /* (11, 19, 27) {real, imag} */,
  {32'hbf5340c0, 32'h00000000} /* (11, 19, 26) {real, imag} */,
  {32'hbf8b3a08, 32'h00000000} /* (11, 19, 25) {real, imag} */,
  {32'hbf8f04fe, 32'h00000000} /* (11, 19, 24) {real, imag} */,
  {32'hbf0196e4, 32'h00000000} /* (11, 19, 23) {real, imag} */,
  {32'hbf69aa8d, 32'h00000000} /* (11, 19, 22) {real, imag} */,
  {32'hbef1baad, 32'h00000000} /* (11, 19, 21) {real, imag} */,
  {32'h3f381e5b, 32'h00000000} /* (11, 19, 20) {real, imag} */,
  {32'h3f098ee5, 32'h00000000} /* (11, 19, 19) {real, imag} */,
  {32'h3ee97c30, 32'h00000000} /* (11, 19, 18) {real, imag} */,
  {32'h3f526b3a, 32'h00000000} /* (11, 19, 17) {real, imag} */,
  {32'h3fb1deda, 32'h00000000} /* (11, 19, 16) {real, imag} */,
  {32'h3ff5ca79, 32'h00000000} /* (11, 19, 15) {real, imag} */,
  {32'h3f569414, 32'h00000000} /* (11, 19, 14) {real, imag} */,
  {32'h3f204878, 32'h00000000} /* (11, 19, 13) {real, imag} */,
  {32'h3f3a992e, 32'h00000000} /* (11, 19, 12) {real, imag} */,
  {32'h3ea9ba1f, 32'h00000000} /* (11, 19, 11) {real, imag} */,
  {32'hbf56fbbe, 32'h00000000} /* (11, 19, 10) {real, imag} */,
  {32'hbf55fa0e, 32'h00000000} /* (11, 19, 9) {real, imag} */,
  {32'hbe9427b8, 32'h00000000} /* (11, 19, 8) {real, imag} */,
  {32'hbf2028af, 32'h00000000} /* (11, 19, 7) {real, imag} */,
  {32'hbef382e6, 32'h00000000} /* (11, 19, 6) {real, imag} */,
  {32'hbf71655a, 32'h00000000} /* (11, 19, 5) {real, imag} */,
  {32'hbf87feb7, 32'h00000000} /* (11, 19, 4) {real, imag} */,
  {32'hbf2d83d4, 32'h00000000} /* (11, 19, 3) {real, imag} */,
  {32'hbf48a825, 32'h00000000} /* (11, 19, 2) {real, imag} */,
  {32'hbf431947, 32'h00000000} /* (11, 19, 1) {real, imag} */,
  {32'hbedf3d25, 32'h00000000} /* (11, 19, 0) {real, imag} */,
  {32'hbf092be6, 32'h00000000} /* (11, 18, 31) {real, imag} */,
  {32'hbfafd4db, 32'h00000000} /* (11, 18, 30) {real, imag} */,
  {32'hbfb337f9, 32'h00000000} /* (11, 18, 29) {real, imag} */,
  {32'hbfb24339, 32'h00000000} /* (11, 18, 28) {real, imag} */,
  {32'hbf788fd6, 32'h00000000} /* (11, 18, 27) {real, imag} */,
  {32'hbf7ae304, 32'h00000000} /* (11, 18, 26) {real, imag} */,
  {32'hbf492c7f, 32'h00000000} /* (11, 18, 25) {real, imag} */,
  {32'hbf42d6a2, 32'h00000000} /* (11, 18, 24) {real, imag} */,
  {32'hbf66001e, 32'h00000000} /* (11, 18, 23) {real, imag} */,
  {32'hbf767ab9, 32'h00000000} /* (11, 18, 22) {real, imag} */,
  {32'hbf0f8ae6, 32'h00000000} /* (11, 18, 21) {real, imag} */,
  {32'h3f294a50, 32'h00000000} /* (11, 18, 20) {real, imag} */,
  {32'h3f52f1c9, 32'h00000000} /* (11, 18, 19) {real, imag} */,
  {32'h3f13d6c7, 32'h00000000} /* (11, 18, 18) {real, imag} */,
  {32'h3ec90969, 32'h00000000} /* (11, 18, 17) {real, imag} */,
  {32'h3efb62ef, 32'h00000000} /* (11, 18, 16) {real, imag} */,
  {32'h3f887fa8, 32'h00000000} /* (11, 18, 15) {real, imag} */,
  {32'h3f045c1c, 32'h00000000} /* (11, 18, 14) {real, imag} */,
  {32'h3f43fb4b, 32'h00000000} /* (11, 18, 13) {real, imag} */,
  {32'h3f22c4b5, 32'h00000000} /* (11, 18, 12) {real, imag} */,
  {32'h3e9899e2, 32'h00000000} /* (11, 18, 11) {real, imag} */,
  {32'hbf124727, 32'h00000000} /* (11, 18, 10) {real, imag} */,
  {32'hbeb9a9cd, 32'h00000000} /* (11, 18, 9) {real, imag} */,
  {32'hbedcf4b4, 32'h00000000} /* (11, 18, 8) {real, imag} */,
  {32'hbfaf7377, 32'h00000000} /* (11, 18, 7) {real, imag} */,
  {32'hbf933e8e, 32'h00000000} /* (11, 18, 6) {real, imag} */,
  {32'hbf73de63, 32'h00000000} /* (11, 18, 5) {real, imag} */,
  {32'hbf4a63f9, 32'h00000000} /* (11, 18, 4) {real, imag} */,
  {32'hbf37ad91, 32'h00000000} /* (11, 18, 3) {real, imag} */,
  {32'hbf58bd4f, 32'h00000000} /* (11, 18, 2) {real, imag} */,
  {32'hbef7e48c, 32'h00000000} /* (11, 18, 1) {real, imag} */,
  {32'hbe848918, 32'h00000000} /* (11, 18, 0) {real, imag} */,
  {32'hbc4f4c8c, 32'h00000000} /* (11, 17, 31) {real, imag} */,
  {32'hbef7bbc8, 32'h00000000} /* (11, 17, 30) {real, imag} */,
  {32'hbf3f4360, 32'h00000000} /* (11, 17, 29) {real, imag} */,
  {32'hbf9c7e33, 32'h00000000} /* (11, 17, 28) {real, imag} */,
  {32'hbf80c2d3, 32'h00000000} /* (11, 17, 27) {real, imag} */,
  {32'hbf3f3ef3, 32'h00000000} /* (11, 17, 26) {real, imag} */,
  {32'hbf135ed7, 32'h00000000} /* (11, 17, 25) {real, imag} */,
  {32'hbf3ef920, 32'h00000000} /* (11, 17, 24) {real, imag} */,
  {32'hbfa4a700, 32'h00000000} /* (11, 17, 23) {real, imag} */,
  {32'hbf777e4b, 32'h00000000} /* (11, 17, 22) {real, imag} */,
  {32'hbf315d47, 32'h00000000} /* (11, 17, 21) {real, imag} */,
  {32'h3f137571, 32'h00000000} /* (11, 17, 20) {real, imag} */,
  {32'h3f9bd831, 32'h00000000} /* (11, 17, 19) {real, imag} */,
  {32'h3fb93e09, 32'h00000000} /* (11, 17, 18) {real, imag} */,
  {32'h3f3852f9, 32'h00000000} /* (11, 17, 17) {real, imag} */,
  {32'h3ef466ed, 32'h00000000} /* (11, 17, 16) {real, imag} */,
  {32'h3f5f3753, 32'h00000000} /* (11, 17, 15) {real, imag} */,
  {32'h3f9392db, 32'h00000000} /* (11, 17, 14) {real, imag} */,
  {32'h3f8af8d9, 32'h00000000} /* (11, 17, 13) {real, imag} */,
  {32'h3f72fe9f, 32'h00000000} /* (11, 17, 12) {real, imag} */,
  {32'h3ec5109d, 32'h00000000} /* (11, 17, 11) {real, imag} */,
  {32'hbf1f56e1, 32'h00000000} /* (11, 17, 10) {real, imag} */,
  {32'hbea60b59, 32'h00000000} /* (11, 17, 9) {real, imag} */,
  {32'hbef2c664, 32'h00000000} /* (11, 17, 8) {real, imag} */,
  {32'hbf948b84, 32'h00000000} /* (11, 17, 7) {real, imag} */,
  {32'hbfc87692, 32'h00000000} /* (11, 17, 6) {real, imag} */,
  {32'hbf85e1c0, 32'h00000000} /* (11, 17, 5) {real, imag} */,
  {32'hbfb04618, 32'h00000000} /* (11, 17, 4) {real, imag} */,
  {32'hc007532c, 32'h00000000} /* (11, 17, 3) {real, imag} */,
  {32'hbfb516b2, 32'h00000000} /* (11, 17, 2) {real, imag} */,
  {32'hbeefbeac, 32'h00000000} /* (11, 17, 1) {real, imag} */,
  {32'hbe0b1a9d, 32'h00000000} /* (11, 17, 0) {real, imag} */,
  {32'hbeb99315, 32'h00000000} /* (11, 16, 31) {real, imag} */,
  {32'hbf60a547, 32'h00000000} /* (11, 16, 30) {real, imag} */,
  {32'hbf2e3945, 32'h00000000} /* (11, 16, 29) {real, imag} */,
  {32'hbf8ea347, 32'h00000000} /* (11, 16, 28) {real, imag} */,
  {32'hbf8cd74a, 32'h00000000} /* (11, 16, 27) {real, imag} */,
  {32'hbf5b1a41, 32'h00000000} /* (11, 16, 26) {real, imag} */,
  {32'hbf42d304, 32'h00000000} /* (11, 16, 25) {real, imag} */,
  {32'hbf85f8c4, 32'h00000000} /* (11, 16, 24) {real, imag} */,
  {32'hbf807176, 32'h00000000} /* (11, 16, 23) {real, imag} */,
  {32'hbef380fa, 32'h00000000} /* (11, 16, 22) {real, imag} */,
  {32'hbe018a77, 32'h00000000} /* (11, 16, 21) {real, imag} */,
  {32'h3f290fd7, 32'h00000000} /* (11, 16, 20) {real, imag} */,
  {32'h3f802168, 32'h00000000} /* (11, 16, 19) {real, imag} */,
  {32'h3f8320b2, 32'h00000000} /* (11, 16, 18) {real, imag} */,
  {32'h3f4a29de, 32'h00000000} /* (11, 16, 17) {real, imag} */,
  {32'h3f82a6cb, 32'h00000000} /* (11, 16, 16) {real, imag} */,
  {32'h3f5404f8, 32'h00000000} /* (11, 16, 15) {real, imag} */,
  {32'h3f97d021, 32'h00000000} /* (11, 16, 14) {real, imag} */,
  {32'h3fab3bd3, 32'h00000000} /* (11, 16, 13) {real, imag} */,
  {32'h3f74bf43, 32'h00000000} /* (11, 16, 12) {real, imag} */,
  {32'h3ea988b8, 32'h00000000} /* (11, 16, 11) {real, imag} */,
  {32'hbf7855cc, 32'h00000000} /* (11, 16, 10) {real, imag} */,
  {32'hbf9985a2, 32'h00000000} /* (11, 16, 9) {real, imag} */,
  {32'hbf90c103, 32'h00000000} /* (11, 16, 8) {real, imag} */,
  {32'hbf832cd5, 32'h00000000} /* (11, 16, 7) {real, imag} */,
  {32'hbf247788, 32'h00000000} /* (11, 16, 6) {real, imag} */,
  {32'hbf2efafa, 32'h00000000} /* (11, 16, 5) {real, imag} */,
  {32'hbf938349, 32'h00000000} /* (11, 16, 4) {real, imag} */,
  {32'hbffdef39, 32'h00000000} /* (11, 16, 3) {real, imag} */,
  {32'hbface347, 32'h00000000} /* (11, 16, 2) {real, imag} */,
  {32'hbf3b9feb, 32'h00000000} /* (11, 16, 1) {real, imag} */,
  {32'hbecc827e, 32'h00000000} /* (11, 16, 0) {real, imag} */,
  {32'hbec2e54b, 32'h00000000} /* (11, 15, 31) {real, imag} */,
  {32'hbfa87479, 32'h00000000} /* (11, 15, 30) {real, imag} */,
  {32'hbf997dfe, 32'h00000000} /* (11, 15, 29) {real, imag} */,
  {32'hbf867123, 32'h00000000} /* (11, 15, 28) {real, imag} */,
  {32'hbf6dfbef, 32'h00000000} /* (11, 15, 27) {real, imag} */,
  {32'hbf92e462, 32'h00000000} /* (11, 15, 26) {real, imag} */,
  {32'hbf67b65a, 32'h00000000} /* (11, 15, 25) {real, imag} */,
  {32'hbf813922, 32'h00000000} /* (11, 15, 24) {real, imag} */,
  {32'hbf61867a, 32'h00000000} /* (11, 15, 23) {real, imag} */,
  {32'hbdfc5201, 32'h00000000} /* (11, 15, 22) {real, imag} */,
  {32'h3f523ec6, 32'h00000000} /* (11, 15, 21) {real, imag} */,
  {32'h3f753f9b, 32'h00000000} /* (11, 15, 20) {real, imag} */,
  {32'h3f0da10c, 32'h00000000} /* (11, 15, 19) {real, imag} */,
  {32'h3f325ed0, 32'h00000000} /* (11, 15, 18) {real, imag} */,
  {32'h3f33c9b7, 32'h00000000} /* (11, 15, 17) {real, imag} */,
  {32'h3f6d4482, 32'h00000000} /* (11, 15, 16) {real, imag} */,
  {32'h3f87cb08, 32'h00000000} /* (11, 15, 15) {real, imag} */,
  {32'h3f4cca27, 32'h00000000} /* (11, 15, 14) {real, imag} */,
  {32'h3f4591c9, 32'h00000000} /* (11, 15, 13) {real, imag} */,
  {32'h3f524028, 32'h00000000} /* (11, 15, 12) {real, imag} */,
  {32'h3ee3403e, 32'h00000000} /* (11, 15, 11) {real, imag} */,
  {32'hbf4046e1, 32'h00000000} /* (11, 15, 10) {real, imag} */,
  {32'hbfb625cd, 32'h00000000} /* (11, 15, 9) {real, imag} */,
  {32'hbfc1cfdf, 32'h00000000} /* (11, 15, 8) {real, imag} */,
  {32'hbfbdcff7, 32'h00000000} /* (11, 15, 7) {real, imag} */,
  {32'hbf6ae1df, 32'h00000000} /* (11, 15, 6) {real, imag} */,
  {32'hbf436211, 32'h00000000} /* (11, 15, 5) {real, imag} */,
  {32'hbf9ccf42, 32'h00000000} /* (11, 15, 4) {real, imag} */,
  {32'hbfaf87e9, 32'h00000000} /* (11, 15, 3) {real, imag} */,
  {32'hbf90ef08, 32'h00000000} /* (11, 15, 2) {real, imag} */,
  {32'hbf8a6fca, 32'h00000000} /* (11, 15, 1) {real, imag} */,
  {32'hbf45989d, 32'h00000000} /* (11, 15, 0) {real, imag} */,
  {32'hbf1f5af7, 32'h00000000} /* (11, 14, 31) {real, imag} */,
  {32'hbfe2af4e, 32'h00000000} /* (11, 14, 30) {real, imag} */,
  {32'hbfc07d9d, 32'h00000000} /* (11, 14, 29) {real, imag} */,
  {32'hbf6e3749, 32'h00000000} /* (11, 14, 28) {real, imag} */,
  {32'hbf3f7b45, 32'h00000000} /* (11, 14, 27) {real, imag} */,
  {32'hbf8b5f6a, 32'h00000000} /* (11, 14, 26) {real, imag} */,
  {32'hbf64a8e8, 32'h00000000} /* (11, 14, 25) {real, imag} */,
  {32'hbf4e0a26, 32'h00000000} /* (11, 14, 24) {real, imag} */,
  {32'hbf6d8f13, 32'h00000000} /* (11, 14, 23) {real, imag} */,
  {32'hbf5696ee, 32'h00000000} /* (11, 14, 22) {real, imag} */,
  {32'hbf455356, 32'h00000000} /* (11, 14, 21) {real, imag} */,
  {32'h3f0b7648, 32'h00000000} /* (11, 14, 20) {real, imag} */,
  {32'h3f541572, 32'h00000000} /* (11, 14, 19) {real, imag} */,
  {32'h3f6533d9, 32'h00000000} /* (11, 14, 18) {real, imag} */,
  {32'h3f38386a, 32'h00000000} /* (11, 14, 17) {real, imag} */,
  {32'h3f1c53bf, 32'h00000000} /* (11, 14, 16) {real, imag} */,
  {32'h3f93c591, 32'h00000000} /* (11, 14, 15) {real, imag} */,
  {32'h3f95badd, 32'h00000000} /* (11, 14, 14) {real, imag} */,
  {32'h3f6c8a6f, 32'h00000000} /* (11, 14, 13) {real, imag} */,
  {32'h3fb8b0b6, 32'h00000000} /* (11, 14, 12) {real, imag} */,
  {32'h3f7ab52d, 32'h00000000} /* (11, 14, 11) {real, imag} */,
  {32'hbda03cc9, 32'h00000000} /* (11, 14, 10) {real, imag} */,
  {32'hbf515de9, 32'h00000000} /* (11, 14, 9) {real, imag} */,
  {32'hbf82349f, 32'h00000000} /* (11, 14, 8) {real, imag} */,
  {32'hbfa02918, 32'h00000000} /* (11, 14, 7) {real, imag} */,
  {32'hbf8db933, 32'h00000000} /* (11, 14, 6) {real, imag} */,
  {32'hbf0d197c, 32'h00000000} /* (11, 14, 5) {real, imag} */,
  {32'hbf63aba9, 32'h00000000} /* (11, 14, 4) {real, imag} */,
  {32'hbf85f4eb, 32'h00000000} /* (11, 14, 3) {real, imag} */,
  {32'hbf7e8045, 32'h00000000} /* (11, 14, 2) {real, imag} */,
  {32'hbfb445c4, 32'h00000000} /* (11, 14, 1) {real, imag} */,
  {32'hbf8c0771, 32'h00000000} /* (11, 14, 0) {real, imag} */,
  {32'hbf7b4044, 32'h00000000} /* (11, 13, 31) {real, imag} */,
  {32'hbfef60ae, 32'h00000000} /* (11, 13, 30) {real, imag} */,
  {32'hbf8ab058, 32'h00000000} /* (11, 13, 29) {real, imag} */,
  {32'hbf8ff7e5, 32'h00000000} /* (11, 13, 28) {real, imag} */,
  {32'hbf2d80c3, 32'h00000000} /* (11, 13, 27) {real, imag} */,
  {32'hbf324030, 32'h00000000} /* (11, 13, 26) {real, imag} */,
  {32'hbf974dc4, 32'h00000000} /* (11, 13, 25) {real, imag} */,
  {32'hbf7bcfe7, 32'h00000000} /* (11, 13, 24) {real, imag} */,
  {32'hbf92b9a6, 32'h00000000} /* (11, 13, 23) {real, imag} */,
  {32'hbf9dfc5c, 32'h00000000} /* (11, 13, 22) {real, imag} */,
  {32'hbf7a29ba, 32'h00000000} /* (11, 13, 21) {real, imag} */,
  {32'h3e9ec787, 32'h00000000} /* (11, 13, 20) {real, imag} */,
  {32'h3f93bcca, 32'h00000000} /* (11, 13, 19) {real, imag} */,
  {32'h3faa1bb7, 32'h00000000} /* (11, 13, 18) {real, imag} */,
  {32'h3f8ff81d, 32'h00000000} /* (11, 13, 17) {real, imag} */,
  {32'h3f82f30b, 32'h00000000} /* (11, 13, 16) {real, imag} */,
  {32'h3f910b22, 32'h00000000} /* (11, 13, 15) {real, imag} */,
  {32'h3f5eba07, 32'h00000000} /* (11, 13, 14) {real, imag} */,
  {32'h3f2ba1cd, 32'h00000000} /* (11, 13, 13) {real, imag} */,
  {32'h3f7e742a, 32'h00000000} /* (11, 13, 12) {real, imag} */,
  {32'h3f432c6e, 32'h00000000} /* (11, 13, 11) {real, imag} */,
  {32'hbe5a2f2a, 32'h00000000} /* (11, 13, 10) {real, imag} */,
  {32'hbf0e784b, 32'h00000000} /* (11, 13, 9) {real, imag} */,
  {32'hbf19a2cb, 32'h00000000} /* (11, 13, 8) {real, imag} */,
  {32'hbf27fc42, 32'h00000000} /* (11, 13, 7) {real, imag} */,
  {32'hbf9bd257, 32'h00000000} /* (11, 13, 6) {real, imag} */,
  {32'hbf1af997, 32'h00000000} /* (11, 13, 5) {real, imag} */,
  {32'hbee43b22, 32'h00000000} /* (11, 13, 4) {real, imag} */,
  {32'hbf2947f7, 32'h00000000} /* (11, 13, 3) {real, imag} */,
  {32'hbf1a5d10, 32'h00000000} /* (11, 13, 2) {real, imag} */,
  {32'hbf7a68d3, 32'h00000000} /* (11, 13, 1) {real, imag} */,
  {32'hbf3b542d, 32'h00000000} /* (11, 13, 0) {real, imag} */,
  {32'hbf4c0258, 32'h00000000} /* (11, 12, 31) {real, imag} */,
  {32'hbf962d07, 32'h00000000} /* (11, 12, 30) {real, imag} */,
  {32'hbf4f41e7, 32'h00000000} /* (11, 12, 29) {real, imag} */,
  {32'hbf4be347, 32'h00000000} /* (11, 12, 28) {real, imag} */,
  {32'hbef2fb36, 32'h00000000} /* (11, 12, 27) {real, imag} */,
  {32'hbea948ac, 32'h00000000} /* (11, 12, 26) {real, imag} */,
  {32'hbf1fa63b, 32'h00000000} /* (11, 12, 25) {real, imag} */,
  {32'hbf9f5652, 32'h00000000} /* (11, 12, 24) {real, imag} */,
  {32'hbfacc3e9, 32'h00000000} /* (11, 12, 23) {real, imag} */,
  {32'hbf8388be, 32'h00000000} /* (11, 12, 22) {real, imag} */,
  {32'hbf592c76, 32'h00000000} /* (11, 12, 21) {real, imag} */,
  {32'h3e594bad, 32'h00000000} /* (11, 12, 20) {real, imag} */,
  {32'h3f7e913a, 32'h00000000} /* (11, 12, 19) {real, imag} */,
  {32'h3facdde4, 32'h00000000} /* (11, 12, 18) {real, imag} */,
  {32'h3fb9131f, 32'h00000000} /* (11, 12, 17) {real, imag} */,
  {32'h3fd91961, 32'h00000000} /* (11, 12, 16) {real, imag} */,
  {32'h3f8f490d, 32'h00000000} /* (11, 12, 15) {real, imag} */,
  {32'h3f6dc159, 32'h00000000} /* (11, 12, 14) {real, imag} */,
  {32'h3f41b066, 32'h00000000} /* (11, 12, 13) {real, imag} */,
  {32'h3f37b16c, 32'h00000000} /* (11, 12, 12) {real, imag} */,
  {32'h3d3bca0e, 32'h00000000} /* (11, 12, 11) {real, imag} */,
  {32'hbf3b2cd4, 32'h00000000} /* (11, 12, 10) {real, imag} */,
  {32'hbf2d4785, 32'h00000000} /* (11, 12, 9) {real, imag} */,
  {32'hbf252bed, 32'h00000000} /* (11, 12, 8) {real, imag} */,
  {32'hbf38dc57, 32'h00000000} /* (11, 12, 7) {real, imag} */,
  {32'hbf9eb686, 32'h00000000} /* (11, 12, 6) {real, imag} */,
  {32'hbf8d1f39, 32'h00000000} /* (11, 12, 5) {real, imag} */,
  {32'hbf73d701, 32'h00000000} /* (11, 12, 4) {real, imag} */,
  {32'hbf3cf5dc, 32'h00000000} /* (11, 12, 3) {real, imag} */,
  {32'hbf20e852, 32'h00000000} /* (11, 12, 2) {real, imag} */,
  {32'hbf427161, 32'h00000000} /* (11, 12, 1) {real, imag} */,
  {32'hbeac140d, 32'h00000000} /* (11, 12, 0) {real, imag} */,
  {32'hbf0ca64a, 32'h00000000} /* (11, 11, 31) {real, imag} */,
  {32'hbf30f1e0, 32'h00000000} /* (11, 11, 30) {real, imag} */,
  {32'hbecdd708, 32'h00000000} /* (11, 11, 29) {real, imag} */,
  {32'hbeac05b0, 32'h00000000} /* (11, 11, 28) {real, imag} */,
  {32'hbead24f6, 32'h00000000} /* (11, 11, 27) {real, imag} */,
  {32'hbeb9084d, 32'h00000000} /* (11, 11, 26) {real, imag} */,
  {32'hbf2cd840, 32'h00000000} /* (11, 11, 25) {real, imag} */,
  {32'hbfb645c5, 32'h00000000} /* (11, 11, 24) {real, imag} */,
  {32'hbf89cb42, 32'h00000000} /* (11, 11, 23) {real, imag} */,
  {32'hbeebc2b6, 32'h00000000} /* (11, 11, 22) {real, imag} */,
  {32'hbe15bc84, 32'h00000000} /* (11, 11, 21) {real, imag} */,
  {32'h3ec0e77c, 32'h00000000} /* (11, 11, 20) {real, imag} */,
  {32'h3f41669f, 32'h00000000} /* (11, 11, 19) {real, imag} */,
  {32'h3f234240, 32'h00000000} /* (11, 11, 18) {real, imag} */,
  {32'h3f49e697, 32'h00000000} /* (11, 11, 17) {real, imag} */,
  {32'h3fdbdf6b, 32'h00000000} /* (11, 11, 16) {real, imag} */,
  {32'h3f808acf, 32'h00000000} /* (11, 11, 15) {real, imag} */,
  {32'h3f53719b, 32'h00000000} /* (11, 11, 14) {real, imag} */,
  {32'h3f69d9f7, 32'h00000000} /* (11, 11, 13) {real, imag} */,
  {32'h3f804f67, 32'h00000000} /* (11, 11, 12) {real, imag} */,
  {32'h3ed370f5, 32'h00000000} /* (11, 11, 11) {real, imag} */,
  {32'hbe238373, 32'h00000000} /* (11, 11, 10) {real, imag} */,
  {32'hbe826d0c, 32'h00000000} /* (11, 11, 9) {real, imag} */,
  {32'hbf324d14, 32'h00000000} /* (11, 11, 8) {real, imag} */,
  {32'hbf3e9533, 32'h00000000} /* (11, 11, 7) {real, imag} */,
  {32'hbf319b6e, 32'h00000000} /* (11, 11, 6) {real, imag} */,
  {32'hbef0cbef, 32'h00000000} /* (11, 11, 5) {real, imag} */,
  {32'hbf7b9589, 32'h00000000} /* (11, 11, 4) {real, imag} */,
  {32'hbf945c7b, 32'h00000000} /* (11, 11, 3) {real, imag} */,
  {32'hbf347b98, 32'h00000000} /* (11, 11, 2) {real, imag} */,
  {32'hbeba9970, 32'h00000000} /* (11, 11, 1) {real, imag} */,
  {32'hbe04dd94, 32'h00000000} /* (11, 11, 0) {real, imag} */,
  {32'h3e43aabe, 32'h00000000} /* (11, 10, 31) {real, imag} */,
  {32'h3f01d5ee, 32'h00000000} /* (11, 10, 30) {real, imag} */,
  {32'h3f278b81, 32'h00000000} /* (11, 10, 29) {real, imag} */,
  {32'h3f3bd0db, 32'h00000000} /* (11, 10, 28) {real, imag} */,
  {32'h3f2873a9, 32'h00000000} /* (11, 10, 27) {real, imag} */,
  {32'h3e8cdd26, 32'h00000000} /* (11, 10, 26) {real, imag} */,
  {32'h3eb6c690, 32'h00000000} /* (11, 10, 25) {real, imag} */,
  {32'h3dda8a99, 32'h00000000} /* (11, 10, 24) {real, imag} */,
  {32'h3efe4f2e, 32'h00000000} /* (11, 10, 23) {real, imag} */,
  {32'h3f8364a6, 32'h00000000} /* (11, 10, 22) {real, imag} */,
  {32'h3f986854, 32'h00000000} /* (11, 10, 21) {real, imag} */,
  {32'h3eb377d9, 32'h00000000} /* (11, 10, 20) {real, imag} */,
  {32'hbef6b254, 32'h00000000} /* (11, 10, 19) {real, imag} */,
  {32'hbf48c734, 32'h00000000} /* (11, 10, 18) {real, imag} */,
  {32'hbf15c61e, 32'h00000000} /* (11, 10, 17) {real, imag} */,
  {32'hbe26ed37, 32'h00000000} /* (11, 10, 16) {real, imag} */,
  {32'hbdddcbee, 32'h00000000} /* (11, 10, 15) {real, imag} */,
  {32'h3ce390a8, 32'h00000000} /* (11, 10, 14) {real, imag} */,
  {32'hbe4d0970, 32'h00000000} /* (11, 10, 13) {real, imag} */,
  {32'hbe621c54, 32'h00000000} /* (11, 10, 12) {real, imag} */,
  {32'hbe2a6a9b, 32'h00000000} /* (11, 10, 11) {real, imag} */,
  {32'h3dd12e42, 32'h00000000} /* (11, 10, 10) {real, imag} */,
  {32'h3f1455b2, 32'h00000000} /* (11, 10, 9) {real, imag} */,
  {32'h3eaeff87, 32'h00000000} /* (11, 10, 8) {real, imag} */,
  {32'h3f86371e, 32'h00000000} /* (11, 10, 7) {real, imag} */,
  {32'h3f6e8d69, 32'h00000000} /* (11, 10, 6) {real, imag} */,
  {32'h3f53ea40, 32'h00000000} /* (11, 10, 5) {real, imag} */,
  {32'h3efdd489, 32'h00000000} /* (11, 10, 4) {real, imag} */,
  {32'hbe81b185, 32'h00000000} /* (11, 10, 3) {real, imag} */,
  {32'hbe4e94c2, 32'h00000000} /* (11, 10, 2) {real, imag} */,
  {32'h3f23c2a3, 32'h00000000} /* (11, 10, 1) {real, imag} */,
  {32'h3eef981f, 32'h00000000} /* (11, 10, 0) {real, imag} */,
  {32'h3ea17e6d, 32'h00000000} /* (11, 9, 31) {real, imag} */,
  {32'h3f3bf8fc, 32'h00000000} /* (11, 9, 30) {real, imag} */,
  {32'h3fa9a1bc, 32'h00000000} /* (11, 9, 29) {real, imag} */,
  {32'h3fcc90ff, 32'h00000000} /* (11, 9, 28) {real, imag} */,
  {32'h3fa61519, 32'h00000000} /* (11, 9, 27) {real, imag} */,
  {32'h3f76ffab, 32'h00000000} /* (11, 9, 26) {real, imag} */,
  {32'h3f3c2a1a, 32'h00000000} /* (11, 9, 25) {real, imag} */,
  {32'h3f1ab4da, 32'h00000000} /* (11, 9, 24) {real, imag} */,
  {32'h3f90741b, 32'h00000000} /* (11, 9, 23) {real, imag} */,
  {32'h3f7d079f, 32'h00000000} /* (11, 9, 22) {real, imag} */,
  {32'h3f31d5f7, 32'h00000000} /* (11, 9, 21) {real, imag} */,
  {32'h3d83e34c, 32'h00000000} /* (11, 9, 20) {real, imag} */,
  {32'hbefff458, 32'h00000000} /* (11, 9, 19) {real, imag} */,
  {32'hbf16a8e3, 32'h00000000} /* (11, 9, 18) {real, imag} */,
  {32'hbf2a2ef7, 32'h00000000} /* (11, 9, 17) {real, imag} */,
  {32'hbf8c17be, 32'h00000000} /* (11, 9, 16) {real, imag} */,
  {32'hbf71ae34, 32'h00000000} /* (11, 9, 15) {real, imag} */,
  {32'hbefb908a, 32'h00000000} /* (11, 9, 14) {real, imag} */,
  {32'hbf10b795, 32'h00000000} /* (11, 9, 13) {real, imag} */,
  {32'hbf424df1, 32'h00000000} /* (11, 9, 12) {real, imag} */,
  {32'hbf11c24c, 32'h00000000} /* (11, 9, 11) {real, imag} */,
  {32'h3ec05492, 32'h00000000} /* (11, 9, 10) {real, imag} */,
  {32'h3f7026ff, 32'h00000000} /* (11, 9, 9) {real, imag} */,
  {32'h3f958c61, 32'h00000000} /* (11, 9, 8) {real, imag} */,
  {32'h3fbc61f2, 32'h00000000} /* (11, 9, 7) {real, imag} */,
  {32'h3f6b7018, 32'h00000000} /* (11, 9, 6) {real, imag} */,
  {32'h3eea6a44, 32'h00000000} /* (11, 9, 5) {real, imag} */,
  {32'h3f106176, 32'h00000000} /* (11, 9, 4) {real, imag} */,
  {32'h3f245240, 32'h00000000} /* (11, 9, 3) {real, imag} */,
  {32'h3ea19e58, 32'h00000000} /* (11, 9, 2) {real, imag} */,
  {32'h3f306351, 32'h00000000} /* (11, 9, 1) {real, imag} */,
  {32'h3efea9a5, 32'h00000000} /* (11, 9, 0) {real, imag} */,
  {32'h3cac7e3e, 32'h00000000} /* (11, 8, 31) {real, imag} */,
  {32'h3eeeff3a, 32'h00000000} /* (11, 8, 30) {real, imag} */,
  {32'h3f704fc7, 32'h00000000} /* (11, 8, 29) {real, imag} */,
  {32'h3fa21c23, 32'h00000000} /* (11, 8, 28) {real, imag} */,
  {32'h3fd8b268, 32'h00000000} /* (11, 8, 27) {real, imag} */,
  {32'h3fcaaeed, 32'h00000000} /* (11, 8, 26) {real, imag} */,
  {32'h3f503cee, 32'h00000000} /* (11, 8, 25) {real, imag} */,
  {32'h3f42b757, 32'h00000000} /* (11, 8, 24) {real, imag} */,
  {32'h3f929d54, 32'h00000000} /* (11, 8, 23) {real, imag} */,
  {32'h3f52501d, 32'h00000000} /* (11, 8, 22) {real, imag} */,
  {32'h3eb49493, 32'h00000000} /* (11, 8, 21) {real, imag} */,
  {32'hbd6c73f3, 32'h00000000} /* (11, 8, 20) {real, imag} */,
  {32'hbe657026, 32'h00000000} /* (11, 8, 19) {real, imag} */,
  {32'hbf2b8668, 32'h00000000} /* (11, 8, 18) {real, imag} */,
  {32'hbf45462a, 32'h00000000} /* (11, 8, 17) {real, imag} */,
  {32'hbf624da9, 32'h00000000} /* (11, 8, 16) {real, imag} */,
  {32'hbf938727, 32'h00000000} /* (11, 8, 15) {real, imag} */,
  {32'hbf0ce31d, 32'h00000000} /* (11, 8, 14) {real, imag} */,
  {32'hbced2503, 32'h00000000} /* (11, 8, 13) {real, imag} */,
  {32'hbec5afb1, 32'h00000000} /* (11, 8, 12) {real, imag} */,
  {32'hbecbaad5, 32'h00000000} /* (11, 8, 11) {real, imag} */,
  {32'h3ea36653, 32'h00000000} /* (11, 8, 10) {real, imag} */,
  {32'h3f09b53b, 32'h00000000} /* (11, 8, 9) {real, imag} */,
  {32'h3f7ca77d, 32'h00000000} /* (11, 8, 8) {real, imag} */,
  {32'h3f345ed5, 32'h00000000} /* (11, 8, 7) {real, imag} */,
  {32'h3f09aeb6, 32'h00000000} /* (11, 8, 6) {real, imag} */,
  {32'h3f2d5bbc, 32'h00000000} /* (11, 8, 5) {real, imag} */,
  {32'h3f04e197, 32'h00000000} /* (11, 8, 4) {real, imag} */,
  {32'h3f144205, 32'h00000000} /* (11, 8, 3) {real, imag} */,
  {32'h3f1e1b66, 32'h00000000} /* (11, 8, 2) {real, imag} */,
  {32'h3f503e26, 32'h00000000} /* (11, 8, 1) {real, imag} */,
  {32'h3ee3e1e4, 32'h00000000} /* (11, 8, 0) {real, imag} */,
  {32'h3eeed502, 32'h00000000} /* (11, 7, 31) {real, imag} */,
  {32'h3f045dae, 32'h00000000} /* (11, 7, 30) {real, imag} */,
  {32'h3f249c94, 32'h00000000} /* (11, 7, 29) {real, imag} */,
  {32'h3f2ce026, 32'h00000000} /* (11, 7, 28) {real, imag} */,
  {32'h3fae5821, 32'h00000000} /* (11, 7, 27) {real, imag} */,
  {32'h3fad8bca, 32'h00000000} /* (11, 7, 26) {real, imag} */,
  {32'h3f483c20, 32'h00000000} /* (11, 7, 25) {real, imag} */,
  {32'h3f3a934f, 32'h00000000} /* (11, 7, 24) {real, imag} */,
  {32'h3f1e6bbf, 32'h00000000} /* (11, 7, 23) {real, imag} */,
  {32'h3f679190, 32'h00000000} /* (11, 7, 22) {real, imag} */,
  {32'h3f82e9eb, 32'h00000000} /* (11, 7, 21) {real, imag} */,
  {32'h3cbcd876, 32'h00000000} /* (11, 7, 20) {real, imag} */,
  {32'hbf010835, 32'h00000000} /* (11, 7, 19) {real, imag} */,
  {32'hbf9166de, 32'h00000000} /* (11, 7, 18) {real, imag} */,
  {32'hbf36be8c, 32'h00000000} /* (11, 7, 17) {real, imag} */,
  {32'hbf73b697, 32'h00000000} /* (11, 7, 16) {real, imag} */,
  {32'hbf6cbbef, 32'h00000000} /* (11, 7, 15) {real, imag} */,
  {32'hbf3b76ce, 32'h00000000} /* (11, 7, 14) {real, imag} */,
  {32'hbed2907f, 32'h00000000} /* (11, 7, 13) {real, imag} */,
  {32'hbf64021e, 32'h00000000} /* (11, 7, 12) {real, imag} */,
  {32'hbf19027d, 32'h00000000} /* (11, 7, 11) {real, imag} */,
  {32'h3e303562, 32'h00000000} /* (11, 7, 10) {real, imag} */,
  {32'h3ef1636b, 32'h00000000} /* (11, 7, 9) {real, imag} */,
  {32'h3f8c77cc, 32'h00000000} /* (11, 7, 8) {real, imag} */,
  {32'h3fc46cb6, 32'h00000000} /* (11, 7, 7) {real, imag} */,
  {32'h3f9c4cce, 32'h00000000} /* (11, 7, 6) {real, imag} */,
  {32'h3f77dc59, 32'h00000000} /* (11, 7, 5) {real, imag} */,
  {32'h3f9736d4, 32'h00000000} /* (11, 7, 4) {real, imag} */,
  {32'h3fa7c07e, 32'h00000000} /* (11, 7, 3) {real, imag} */,
  {32'h3f705152, 32'h00000000} /* (11, 7, 2) {real, imag} */,
  {32'h3ef17358, 32'h00000000} /* (11, 7, 1) {real, imag} */,
  {32'h3e1b3c84, 32'h00000000} /* (11, 7, 0) {real, imag} */,
  {32'h3f0e6bfc, 32'h00000000} /* (11, 6, 31) {real, imag} */,
  {32'h3eef5ec4, 32'h00000000} /* (11, 6, 30) {real, imag} */,
  {32'h3ed22dd7, 32'h00000000} /* (11, 6, 29) {real, imag} */,
  {32'h3f448991, 32'h00000000} /* (11, 6, 28) {real, imag} */,
  {32'h3fa43264, 32'h00000000} /* (11, 6, 27) {real, imag} */,
  {32'h3fb1c865, 32'h00000000} /* (11, 6, 26) {real, imag} */,
  {32'h3f39b22d, 32'h00000000} /* (11, 6, 25) {real, imag} */,
  {32'h3f21849a, 32'h00000000} /* (11, 6, 24) {real, imag} */,
  {32'h3ede7837, 32'h00000000} /* (11, 6, 23) {real, imag} */,
  {32'h3ed1770c, 32'h00000000} /* (11, 6, 22) {real, imag} */,
  {32'h3f488d91, 32'h00000000} /* (11, 6, 21) {real, imag} */,
  {32'hbe75c6fa, 32'h00000000} /* (11, 6, 20) {real, imag} */,
  {32'hbee2cdbe, 32'h00000000} /* (11, 6, 19) {real, imag} */,
  {32'hbfc2c52e, 32'h00000000} /* (11, 6, 18) {real, imag} */,
  {32'hbf9baa04, 32'h00000000} /* (11, 6, 17) {real, imag} */,
  {32'hbfa1c39c, 32'h00000000} /* (11, 6, 16) {real, imag} */,
  {32'hbf394585, 32'h00000000} /* (11, 6, 15) {real, imag} */,
  {32'hbf8a70f5, 32'h00000000} /* (11, 6, 14) {real, imag} */,
  {32'hbf6e2db4, 32'h00000000} /* (11, 6, 13) {real, imag} */,
  {32'hbfa9bdb1, 32'h00000000} /* (11, 6, 12) {real, imag} */,
  {32'hbf865dc2, 32'h00000000} /* (11, 6, 11) {real, imag} */,
  {32'hbdcc132a, 32'h00000000} /* (11, 6, 10) {real, imag} */,
  {32'h3ed6edb7, 32'h00000000} /* (11, 6, 9) {real, imag} */,
  {32'h3fdb8e34, 32'h00000000} /* (11, 6, 8) {real, imag} */,
  {32'h3fdd9466, 32'h00000000} /* (11, 6, 7) {real, imag} */,
  {32'h3f61e054, 32'h00000000} /* (11, 6, 6) {real, imag} */,
  {32'h3ef44d77, 32'h00000000} /* (11, 6, 5) {real, imag} */,
  {32'h3f826730, 32'h00000000} /* (11, 6, 4) {real, imag} */,
  {32'h3f8d4fd3, 32'h00000000} /* (11, 6, 3) {real, imag} */,
  {32'h3f7fc47f, 32'h00000000} /* (11, 6, 2) {real, imag} */,
  {32'h3f94ebcf, 32'h00000000} /* (11, 6, 1) {real, imag} */,
  {32'h3f1bae8f, 32'h00000000} /* (11, 6, 0) {real, imag} */,
  {32'h3e5a3962, 32'h00000000} /* (11, 5, 31) {real, imag} */,
  {32'h3f1ea4b5, 32'h00000000} /* (11, 5, 30) {real, imag} */,
  {32'h3f597a6c, 32'h00000000} /* (11, 5, 29) {real, imag} */,
  {32'h3f514c81, 32'h00000000} /* (11, 5, 28) {real, imag} */,
  {32'h3fd3ff55, 32'h00000000} /* (11, 5, 27) {real, imag} */,
  {32'h3fac263c, 32'h00000000} /* (11, 5, 26) {real, imag} */,
  {32'h3f43b9ab, 32'h00000000} /* (11, 5, 25) {real, imag} */,
  {32'h3f02ed63, 32'h00000000} /* (11, 5, 24) {real, imag} */,
  {32'h3f8b1cec, 32'h00000000} /* (11, 5, 23) {real, imag} */,
  {32'h3f5cf124, 32'h00000000} /* (11, 5, 22) {real, imag} */,
  {32'h3ef8fbae, 32'h00000000} /* (11, 5, 21) {real, imag} */,
  {32'h3e6f6c6a, 32'h00000000} /* (11, 5, 20) {real, imag} */,
  {32'h3f3746ab, 32'h00000000} /* (11, 5, 19) {real, imag} */,
  {32'h3f0758d4, 32'h00000000} /* (11, 5, 18) {real, imag} */,
  {32'h3e30dd67, 32'h00000000} /* (11, 5, 17) {real, imag} */,
  {32'hbea1460e, 32'h00000000} /* (11, 5, 16) {real, imag} */,
  {32'hbf491617, 32'h00000000} /* (11, 5, 15) {real, imag} */,
  {32'hbf99727d, 32'h00000000} /* (11, 5, 14) {real, imag} */,
  {32'hbf165957, 32'h00000000} /* (11, 5, 13) {real, imag} */,
  {32'hbf6cd749, 32'h00000000} /* (11, 5, 12) {real, imag} */,
  {32'hbfbd189d, 32'h00000000} /* (11, 5, 11) {real, imag} */,
  {32'hbe9cecc2, 32'h00000000} /* (11, 5, 10) {real, imag} */,
  {32'hbc860964, 32'h00000000} /* (11, 5, 9) {real, imag} */,
  {32'h3ed13f6b, 32'h00000000} /* (11, 5, 8) {real, imag} */,
  {32'h3c1951a4, 32'h00000000} /* (11, 5, 7) {real, imag} */,
  {32'hbf0ee4fa, 32'h00000000} /* (11, 5, 6) {real, imag} */,
  {32'hbe167d94, 32'h00000000} /* (11, 5, 5) {real, imag} */,
  {32'h3f048ab3, 32'h00000000} /* (11, 5, 4) {real, imag} */,
  {32'h3f9b0791, 32'h00000000} /* (11, 5, 3) {real, imag} */,
  {32'h3fac496d, 32'h00000000} /* (11, 5, 2) {real, imag} */,
  {32'h3fb5f3b0, 32'h00000000} /* (11, 5, 1) {real, imag} */,
  {32'h3edafc6f, 32'h00000000} /* (11, 5, 0) {real, imag} */,
  {32'h3e3bca35, 32'h00000000} /* (11, 4, 31) {real, imag} */,
  {32'h3f66d448, 32'h00000000} /* (11, 4, 30) {real, imag} */,
  {32'h3f89ed56, 32'h00000000} /* (11, 4, 29) {real, imag} */,
  {32'h3f197705, 32'h00000000} /* (11, 4, 28) {real, imag} */,
  {32'h3f2e737d, 32'h00000000} /* (11, 4, 27) {real, imag} */,
  {32'h3f2c5bd1, 32'h00000000} /* (11, 4, 26) {real, imag} */,
  {32'h3f848850, 32'h00000000} /* (11, 4, 25) {real, imag} */,
  {32'h3ee81008, 32'h00000000} /* (11, 4, 24) {real, imag} */,
  {32'h3f8b66d0, 32'h00000000} /* (11, 4, 23) {real, imag} */,
  {32'h3fcd7c9d, 32'h00000000} /* (11, 4, 22) {real, imag} */,
  {32'h3fb82d42, 32'h00000000} /* (11, 4, 21) {real, imag} */,
  {32'h3fb0f1bf, 32'h00000000} /* (11, 4, 20) {real, imag} */,
  {32'h3faded82, 32'h00000000} /* (11, 4, 19) {real, imag} */,
  {32'h3fc4cc58, 32'h00000000} /* (11, 4, 18) {real, imag} */,
  {32'h3fe98e44, 32'h00000000} /* (11, 4, 17) {real, imag} */,
  {32'h3f91604f, 32'h00000000} /* (11, 4, 16) {real, imag} */,
  {32'hbf30c1d8, 32'h00000000} /* (11, 4, 15) {real, imag} */,
  {32'hbf24314d, 32'h00000000} /* (11, 4, 14) {real, imag} */,
  {32'hbef4bb92, 32'h00000000} /* (11, 4, 13) {real, imag} */,
  {32'hbf14677d, 32'h00000000} /* (11, 4, 12) {real, imag} */,
  {32'hbf8da697, 32'h00000000} /* (11, 4, 11) {real, imag} */,
  {32'hbf0bd762, 32'h00000000} /* (11, 4, 10) {real, imag} */,
  {32'hbf390a22, 32'h00000000} /* (11, 4, 9) {real, imag} */,
  {32'hbfac80ff, 32'h00000000} /* (11, 4, 8) {real, imag} */,
  {32'hbf6bea82, 32'h00000000} /* (11, 4, 7) {real, imag} */,
  {32'hbf2a097a, 32'h00000000} /* (11, 4, 6) {real, imag} */,
  {32'h3d8215fe, 32'h00000000} /* (11, 4, 5) {real, imag} */,
  {32'h3f22b0da, 32'h00000000} /* (11, 4, 4) {real, imag} */,
  {32'h3f7e2a16, 32'h00000000} /* (11, 4, 3) {real, imag} */,
  {32'h3f861507, 32'h00000000} /* (11, 4, 2) {real, imag} */,
  {32'h3f6d9ea0, 32'h00000000} /* (11, 4, 1) {real, imag} */,
  {32'h3e8472c8, 32'h00000000} /* (11, 4, 0) {real, imag} */,
  {32'h3e9a1464, 32'h00000000} /* (11, 3, 31) {real, imag} */,
  {32'h3f848374, 32'h00000000} /* (11, 3, 30) {real, imag} */,
  {32'h3fe18fdf, 32'h00000000} /* (11, 3, 29) {real, imag} */,
  {32'h3fa522ce, 32'h00000000} /* (11, 3, 28) {real, imag} */,
  {32'h3ef9f884, 32'h00000000} /* (11, 3, 27) {real, imag} */,
  {32'h3eb9ef93, 32'h00000000} /* (11, 3, 26) {real, imag} */,
  {32'h3f5cdaaa, 32'h00000000} /* (11, 3, 25) {real, imag} */,
  {32'h3f52efff, 32'h00000000} /* (11, 3, 24) {real, imag} */,
  {32'h3f7100b1, 32'h00000000} /* (11, 3, 23) {real, imag} */,
  {32'h3f988131, 32'h00000000} /* (11, 3, 22) {real, imag} */,
  {32'h3f8f9b9e, 32'h00000000} /* (11, 3, 21) {real, imag} */,
  {32'h3f87195c, 32'h00000000} /* (11, 3, 20) {real, imag} */,
  {32'h3f8c2520, 32'h00000000} /* (11, 3, 19) {real, imag} */,
  {32'h3f766d47, 32'h00000000} /* (11, 3, 18) {real, imag} */,
  {32'h3f8f61f2, 32'h00000000} /* (11, 3, 17) {real, imag} */,
  {32'h3f24d387, 32'h00000000} /* (11, 3, 16) {real, imag} */,
  {32'hbf76a31b, 32'h00000000} /* (11, 3, 15) {real, imag} */,
  {32'hbf494df8, 32'h00000000} /* (11, 3, 14) {real, imag} */,
  {32'hbf67998d, 32'h00000000} /* (11, 3, 13) {real, imag} */,
  {32'hbf37fa87, 32'h00000000} /* (11, 3, 12) {real, imag} */,
  {32'hbf5b25ba, 32'h00000000} /* (11, 3, 11) {real, imag} */,
  {32'hbf6a3335, 32'h00000000} /* (11, 3, 10) {real, imag} */,
  {32'hbf54bebe, 32'h00000000} /* (11, 3, 9) {real, imag} */,
  {32'hbfb5b089, 32'h00000000} /* (11, 3, 8) {real, imag} */,
  {32'hbf810f64, 32'h00000000} /* (11, 3, 7) {real, imag} */,
  {32'hbfa2cd4d, 32'h00000000} /* (11, 3, 6) {real, imag} */,
  {32'hbe3c0b8c, 32'h00000000} /* (11, 3, 5) {real, imag} */,
  {32'h3f637e7e, 32'h00000000} /* (11, 3, 4) {real, imag} */,
  {32'h3eed6d5e, 32'h00000000} /* (11, 3, 3) {real, imag} */,
  {32'h3f6d9533, 32'h00000000} /* (11, 3, 2) {real, imag} */,
  {32'h3f3a1668, 32'h00000000} /* (11, 3, 1) {real, imag} */,
  {32'h3e5d4894, 32'h00000000} /* (11, 3, 0) {real, imag} */,
  {32'h3ee60ad6, 32'h00000000} /* (11, 2, 31) {real, imag} */,
  {32'h3f58432c, 32'h00000000} /* (11, 2, 30) {real, imag} */,
  {32'h3fae6ca1, 32'h00000000} /* (11, 2, 29) {real, imag} */,
  {32'h3fc4de7b, 32'h00000000} /* (11, 2, 28) {real, imag} */,
  {32'h3f520596, 32'h00000000} /* (11, 2, 27) {real, imag} */,
  {32'h3ecc2aa2, 32'h00000000} /* (11, 2, 26) {real, imag} */,
  {32'h3f4296ea, 32'h00000000} /* (11, 2, 25) {real, imag} */,
  {32'h3f8205c7, 32'h00000000} /* (11, 2, 24) {real, imag} */,
  {32'h3f99a5a1, 32'h00000000} /* (11, 2, 23) {real, imag} */,
  {32'h3eda0173, 32'h00000000} /* (11, 2, 22) {real, imag} */,
  {32'h3f3b4e2f, 32'h00000000} /* (11, 2, 21) {real, imag} */,
  {32'h3fa62928, 32'h00000000} /* (11, 2, 20) {real, imag} */,
  {32'h3f986c88, 32'h00000000} /* (11, 2, 19) {real, imag} */,
  {32'h3f62f5bc, 32'h00000000} /* (11, 2, 18) {real, imag} */,
  {32'h3f22d411, 32'h00000000} /* (11, 2, 17) {real, imag} */,
  {32'h3dd7161c, 32'h00000000} /* (11, 2, 16) {real, imag} */,
  {32'hbf7923ba, 32'h00000000} /* (11, 2, 15) {real, imag} */,
  {32'hbf88c69c, 32'h00000000} /* (11, 2, 14) {real, imag} */,
  {32'hbf984cd2, 32'h00000000} /* (11, 2, 13) {real, imag} */,
  {32'hbf861448, 32'h00000000} /* (11, 2, 12) {real, imag} */,
  {32'hbf594f03, 32'h00000000} /* (11, 2, 11) {real, imag} */,
  {32'hbf81c7d6, 32'h00000000} /* (11, 2, 10) {real, imag} */,
  {32'hbf365e5e, 32'h00000000} /* (11, 2, 9) {real, imag} */,
  {32'hbf8b2df1, 32'h00000000} /* (11, 2, 8) {real, imag} */,
  {32'hbf9748b1, 32'h00000000} /* (11, 2, 7) {real, imag} */,
  {32'hbfc6248f, 32'h00000000} /* (11, 2, 6) {real, imag} */,
  {32'hbea02376, 32'h00000000} /* (11, 2, 5) {real, imag} */,
  {32'h3f924efa, 32'h00000000} /* (11, 2, 4) {real, imag} */,
  {32'h3f4f3a9e, 32'h00000000} /* (11, 2, 3) {real, imag} */,
  {32'h3f89b538, 32'h00000000} /* (11, 2, 2) {real, imag} */,
  {32'h3f62cdb7, 32'h00000000} /* (11, 2, 1) {real, imag} */,
  {32'h3e9682dc, 32'h00000000} /* (11, 2, 0) {real, imag} */,
  {32'h3efb2ae1, 32'h00000000} /* (11, 1, 31) {real, imag} */,
  {32'h3f804cda, 32'h00000000} /* (11, 1, 30) {real, imag} */,
  {32'h3fb16b91, 32'h00000000} /* (11, 1, 29) {real, imag} */,
  {32'h3fd21fa0, 32'h00000000} /* (11, 1, 28) {real, imag} */,
  {32'h3fc7ea0d, 32'h00000000} /* (11, 1, 27) {real, imag} */,
  {32'h3f5ac1d5, 32'h00000000} /* (11, 1, 26) {real, imag} */,
  {32'h3f26b65e, 32'h00000000} /* (11, 1, 25) {real, imag} */,
  {32'h3f96ef9d, 32'h00000000} /* (11, 1, 24) {real, imag} */,
  {32'h3f9aef2b, 32'h00000000} /* (11, 1, 23) {real, imag} */,
  {32'h3e9cea60, 32'h00000000} /* (11, 1, 22) {real, imag} */,
  {32'h3f294eaf, 32'h00000000} /* (11, 1, 21) {real, imag} */,
  {32'h3f97e7bd, 32'h00000000} /* (11, 1, 20) {real, imag} */,
  {32'h3f888470, 32'h00000000} /* (11, 1, 19) {real, imag} */,
  {32'h3f8c3f28, 32'h00000000} /* (11, 1, 18) {real, imag} */,
  {32'h3ed26fd9, 32'h00000000} /* (11, 1, 17) {real, imag} */,
  {32'h3e006001, 32'h00000000} /* (11, 1, 16) {real, imag} */,
  {32'hbf554ba0, 32'h00000000} /* (11, 1, 15) {real, imag} */,
  {32'hbf7da642, 32'h00000000} /* (11, 1, 14) {real, imag} */,
  {32'hbf8026e2, 32'h00000000} /* (11, 1, 13) {real, imag} */,
  {32'hbf86e16b, 32'h00000000} /* (11, 1, 12) {real, imag} */,
  {32'hbf0f40a7, 32'h00000000} /* (11, 1, 11) {real, imag} */,
  {32'hbf3a8817, 32'h00000000} /* (11, 1, 10) {real, imag} */,
  {32'hbeddf953, 32'h00000000} /* (11, 1, 9) {real, imag} */,
  {32'hbf4087d6, 32'h00000000} /* (11, 1, 8) {real, imag} */,
  {32'hbf9c47ac, 32'h00000000} /* (11, 1, 7) {real, imag} */,
  {32'hbf78e490, 32'h00000000} /* (11, 1, 6) {real, imag} */,
  {32'h3d7aaf90, 32'h00000000} /* (11, 1, 5) {real, imag} */,
  {32'h3f33828d, 32'h00000000} /* (11, 1, 4) {real, imag} */,
  {32'h3f0df71c, 32'h00000000} /* (11, 1, 3) {real, imag} */,
  {32'h3f073fae, 32'h00000000} /* (11, 1, 2) {real, imag} */,
  {32'h3f77076c, 32'h00000000} /* (11, 1, 1) {real, imag} */,
  {32'h3f188720, 32'h00000000} /* (11, 1, 0) {real, imag} */,
  {32'h3e6e8f46, 32'h00000000} /* (11, 0, 31) {real, imag} */,
  {32'h3f02cf11, 32'h00000000} /* (11, 0, 30) {real, imag} */,
  {32'h3f3f766f, 32'h00000000} /* (11, 0, 29) {real, imag} */,
  {32'h3f87c057, 32'h00000000} /* (11, 0, 28) {real, imag} */,
  {32'h3fa37f96, 32'h00000000} /* (11, 0, 27) {real, imag} */,
  {32'h3f28cc52, 32'h00000000} /* (11, 0, 26) {real, imag} */,
  {32'h3edb52f3, 32'h00000000} /* (11, 0, 25) {real, imag} */,
  {32'h3f32b141, 32'h00000000} /* (11, 0, 24) {real, imag} */,
  {32'h3f487237, 32'h00000000} /* (11, 0, 23) {real, imag} */,
  {32'h3ec66125, 32'h00000000} /* (11, 0, 22) {real, imag} */,
  {32'h3e7a0b46, 32'h00000000} /* (11, 0, 21) {real, imag} */,
  {32'h3e327438, 32'h00000000} /* (11, 0, 20) {real, imag} */,
  {32'h3f195dba, 32'h00000000} /* (11, 0, 19) {real, imag} */,
  {32'h3f28c4a1, 32'h00000000} /* (11, 0, 18) {real, imag} */,
  {32'h3e950132, 32'h00000000} /* (11, 0, 17) {real, imag} */,
  {32'h3e18182b, 32'h00000000} /* (11, 0, 16) {real, imag} */,
  {32'hbebd32b7, 32'h00000000} /* (11, 0, 15) {real, imag} */,
  {32'hbf11dc3e, 32'h00000000} /* (11, 0, 14) {real, imag} */,
  {32'hbeca4200, 32'h00000000} /* (11, 0, 13) {real, imag} */,
  {32'hbebbb9e0, 32'h00000000} /* (11, 0, 12) {real, imag} */,
  {32'hbe9f84dc, 32'h00000000} /* (11, 0, 11) {real, imag} */,
  {32'hbe0e9535, 32'h00000000} /* (11, 0, 10) {real, imag} */,
  {32'hbd81e5c5, 32'h00000000} /* (11, 0, 9) {real, imag} */,
  {32'hbeef4bba, 32'h00000000} /* (11, 0, 8) {real, imag} */,
  {32'hbf3b90b3, 32'h00000000} /* (11, 0, 7) {real, imag} */,
  {32'hbed76b32, 32'h00000000} /* (11, 0, 6) {real, imag} */,
  {32'h3e3d83ab, 32'h00000000} /* (11, 0, 5) {real, imag} */,
  {32'h3ea81459, 32'h00000000} /* (11, 0, 4) {real, imag} */,
  {32'h3f077351, 32'h00000000} /* (11, 0, 3) {real, imag} */,
  {32'h3f18461d, 32'h00000000} /* (11, 0, 2) {real, imag} */,
  {32'h3f2de68d, 32'h00000000} /* (11, 0, 1) {real, imag} */,
  {32'h3f06498a, 32'h00000000} /* (11, 0, 0) {real, imag} */,
  {32'h3dac3d72, 32'h00000000} /* (10, 31, 31) {real, imag} */,
  {32'h3eab9b3b, 32'h00000000} /* (10, 31, 30) {real, imag} */,
  {32'h3efba43c, 32'h00000000} /* (10, 31, 29) {real, imag} */,
  {32'h3f01090a, 32'h00000000} /* (10, 31, 28) {real, imag} */,
  {32'h3efa9646, 32'h00000000} /* (10, 31, 27) {real, imag} */,
  {32'h3e4796ac, 32'h00000000} /* (10, 31, 26) {real, imag} */,
  {32'h3f015137, 32'h00000000} /* (10, 31, 25) {real, imag} */,
  {32'h3f6098d3, 32'h00000000} /* (10, 31, 24) {real, imag} */,
  {32'h3f69d14d, 32'h00000000} /* (10, 31, 23) {real, imag} */,
  {32'h3f8fef68, 32'h00000000} /* (10, 31, 22) {real, imag} */,
  {32'h3f22be2a, 32'h00000000} /* (10, 31, 21) {real, imag} */,
  {32'hbe894c5c, 32'h00000000} /* (10, 31, 20) {real, imag} */,
  {32'hbe88b3ae, 32'h00000000} /* (10, 31, 19) {real, imag} */,
  {32'hbcf3415e, 32'h00000000} /* (10, 31, 18) {real, imag} */,
  {32'h3d619560, 32'h00000000} /* (10, 31, 17) {real, imag} */,
  {32'hbf34d7ad, 32'h00000000} /* (10, 31, 16) {real, imag} */,
  {32'hbf64fa91, 32'h00000000} /* (10, 31, 15) {real, imag} */,
  {32'hbf2400cd, 32'h00000000} /* (10, 31, 14) {real, imag} */,
  {32'hbf8e0e49, 32'h00000000} /* (10, 31, 13) {real, imag} */,
  {32'hbf55d9f4, 32'h00000000} /* (10, 31, 12) {real, imag} */,
  {32'hbed3a087, 32'h00000000} /* (10, 31, 11) {real, imag} */,
  {32'h3dae234c, 32'h00000000} /* (10, 31, 10) {real, imag} */,
  {32'h3e9950c6, 32'h00000000} /* (10, 31, 9) {real, imag} */,
  {32'h3f217811, 32'h00000000} /* (10, 31, 8) {real, imag} */,
  {32'h3f0d1a23, 32'h00000000} /* (10, 31, 7) {real, imag} */,
  {32'h3f2fcb24, 32'h00000000} /* (10, 31, 6) {real, imag} */,
  {32'h3eacc68f, 32'h00000000} /* (10, 31, 5) {real, imag} */,
  {32'h3eaae70f, 32'h00000000} /* (10, 31, 4) {real, imag} */,
  {32'h3e9254e9, 32'h00000000} /* (10, 31, 3) {real, imag} */,
  {32'h3ecce9b5, 32'h00000000} /* (10, 31, 2) {real, imag} */,
  {32'h3f3a6bc2, 32'h00000000} /* (10, 31, 1) {real, imag} */,
  {32'h3f082fc3, 32'h00000000} /* (10, 31, 0) {real, imag} */,
  {32'h3f1a00c1, 32'h00000000} /* (10, 30, 31) {real, imag} */,
  {32'h3f829ec4, 32'h00000000} /* (10, 30, 30) {real, imag} */,
  {32'h3f56cf98, 32'h00000000} /* (10, 30, 29) {real, imag} */,
  {32'h3f7093f9, 32'h00000000} /* (10, 30, 28) {real, imag} */,
  {32'h3f28b765, 32'h00000000} /* (10, 30, 27) {real, imag} */,
  {32'h3f06d999, 32'h00000000} /* (10, 30, 26) {real, imag} */,
  {32'h3f3a1b64, 32'h00000000} /* (10, 30, 25) {real, imag} */,
  {32'h3f8814c2, 32'h00000000} /* (10, 30, 24) {real, imag} */,
  {32'h3f421d90, 32'h00000000} /* (10, 30, 23) {real, imag} */,
  {32'h3f590ede, 32'h00000000} /* (10, 30, 22) {real, imag} */,
  {32'h3ef6a8b9, 32'h00000000} /* (10, 30, 21) {real, imag} */,
  {32'hbe9ba5f1, 32'h00000000} /* (10, 30, 20) {real, imag} */,
  {32'hbec97c06, 32'h00000000} /* (10, 30, 19) {real, imag} */,
  {32'hbf05ff85, 32'h00000000} /* (10, 30, 18) {real, imag} */,
  {32'hbe884824, 32'h00000000} /* (10, 30, 17) {real, imag} */,
  {32'hbf49652a, 32'h00000000} /* (10, 30, 16) {real, imag} */,
  {32'hbf771e09, 32'h00000000} /* (10, 30, 15) {real, imag} */,
  {32'hbf71afe1, 32'h00000000} /* (10, 30, 14) {real, imag} */,
  {32'hbfaf0539, 32'h00000000} /* (10, 30, 13) {real, imag} */,
  {32'hbfab485e, 32'h00000000} /* (10, 30, 12) {real, imag} */,
  {32'hbefb9219, 32'h00000000} /* (10, 30, 11) {real, imag} */,
  {32'h3ef7aa2c, 32'h00000000} /* (10, 30, 10) {real, imag} */,
  {32'h3f4565aa, 32'h00000000} /* (10, 30, 9) {real, imag} */,
  {32'h3fb22181, 32'h00000000} /* (10, 30, 8) {real, imag} */,
  {32'h3f8b4948, 32'h00000000} /* (10, 30, 7) {real, imag} */,
  {32'h3f2cc576, 32'h00000000} /* (10, 30, 6) {real, imag} */,
  {32'h3f4b6acc, 32'h00000000} /* (10, 30, 5) {real, imag} */,
  {32'h3f7fb399, 32'h00000000} /* (10, 30, 4) {real, imag} */,
  {32'h3f3272d9, 32'h00000000} /* (10, 30, 3) {real, imag} */,
  {32'h3f55de50, 32'h00000000} /* (10, 30, 2) {real, imag} */,
  {32'h3f77ca97, 32'h00000000} /* (10, 30, 1) {real, imag} */,
  {32'h3f0a3f86, 32'h00000000} /* (10, 30, 0) {real, imag} */,
  {32'h3f616a9a, 32'h00000000} /* (10, 29, 31) {real, imag} */,
  {32'h3f9ddd96, 32'h00000000} /* (10, 29, 30) {real, imag} */,
  {32'h3f3274b0, 32'h00000000} /* (10, 29, 29) {real, imag} */,
  {32'h3f2cf65e, 32'h00000000} /* (10, 29, 28) {real, imag} */,
  {32'h3f41817c, 32'h00000000} /* (10, 29, 27) {real, imag} */,
  {32'h3f7dc144, 32'h00000000} /* (10, 29, 26) {real, imag} */,
  {32'h3f25cb2b, 32'h00000000} /* (10, 29, 25) {real, imag} */,
  {32'h3f35a8d7, 32'h00000000} /* (10, 29, 24) {real, imag} */,
  {32'h3f0e2f8c, 32'h00000000} /* (10, 29, 23) {real, imag} */,
  {32'h3f19c323, 32'h00000000} /* (10, 29, 22) {real, imag} */,
  {32'h3eb55de5, 32'h00000000} /* (10, 29, 21) {real, imag} */,
  {32'hbed38509, 32'h00000000} /* (10, 29, 20) {real, imag} */,
  {32'hbf1da40d, 32'h00000000} /* (10, 29, 19) {real, imag} */,
  {32'hbf515abc, 32'h00000000} /* (10, 29, 18) {real, imag} */,
  {32'hbe8465cd, 32'h00000000} /* (10, 29, 17) {real, imag} */,
  {32'hbeada901, 32'h00000000} /* (10, 29, 16) {real, imag} */,
  {32'hbf794ce7, 32'h00000000} /* (10, 29, 15) {real, imag} */,
  {32'hbf197bb1, 32'h00000000} /* (10, 29, 14) {real, imag} */,
  {32'hbf1eb6df, 32'h00000000} /* (10, 29, 13) {real, imag} */,
  {32'hbf746d45, 32'h00000000} /* (10, 29, 12) {real, imag} */,
  {32'hbf16a1e8, 32'h00000000} /* (10, 29, 11) {real, imag} */,
  {32'h3f0b5374, 32'h00000000} /* (10, 29, 10) {real, imag} */,
  {32'h3f3b2fa9, 32'h00000000} /* (10, 29, 9) {real, imag} */,
  {32'h3f886232, 32'h00000000} /* (10, 29, 8) {real, imag} */,
  {32'h3f8528e4, 32'h00000000} /* (10, 29, 7) {real, imag} */,
  {32'h3f185f65, 32'h00000000} /* (10, 29, 6) {real, imag} */,
  {32'h3f132360, 32'h00000000} /* (10, 29, 5) {real, imag} */,
  {32'h3f9027c5, 32'h00000000} /* (10, 29, 4) {real, imag} */,
  {32'h3f877757, 32'h00000000} /* (10, 29, 3) {real, imag} */,
  {32'h3f1fb323, 32'h00000000} /* (10, 29, 2) {real, imag} */,
  {32'h3f70584e, 32'h00000000} /* (10, 29, 1) {real, imag} */,
  {32'h3f14f81d, 32'h00000000} /* (10, 29, 0) {real, imag} */,
  {32'h3f4207b1, 32'h00000000} /* (10, 28, 31) {real, imag} */,
  {32'h3f63278e, 32'h00000000} /* (10, 28, 30) {real, imag} */,
  {32'h3f18c36a, 32'h00000000} /* (10, 28, 29) {real, imag} */,
  {32'h3f11adcd, 32'h00000000} /* (10, 28, 28) {real, imag} */,
  {32'h3f8c5c68, 32'h00000000} /* (10, 28, 27) {real, imag} */,
  {32'h3f889be8, 32'h00000000} /* (10, 28, 26) {real, imag} */,
  {32'h3f31ff80, 32'h00000000} /* (10, 28, 25) {real, imag} */,
  {32'h3fa112d6, 32'h00000000} /* (10, 28, 24) {real, imag} */,
  {32'h3f94c563, 32'h00000000} /* (10, 28, 23) {real, imag} */,
  {32'h3f89505f, 32'h00000000} /* (10, 28, 22) {real, imag} */,
  {32'h3e0dc50d, 32'h00000000} /* (10, 28, 21) {real, imag} */,
  {32'hbf1a7e59, 32'h00000000} /* (10, 28, 20) {real, imag} */,
  {32'hbf62ba27, 32'h00000000} /* (10, 28, 19) {real, imag} */,
  {32'hbf6cb9b5, 32'h00000000} /* (10, 28, 18) {real, imag} */,
  {32'hbf1f85ba, 32'h00000000} /* (10, 28, 17) {real, imag} */,
  {32'hbf5f7401, 32'h00000000} /* (10, 28, 16) {real, imag} */,
  {32'hbfaf6a27, 32'h00000000} /* (10, 28, 15) {real, imag} */,
  {32'hbf4ea639, 32'h00000000} /* (10, 28, 14) {real, imag} */,
  {32'hbf08aa3d, 32'h00000000} /* (10, 28, 13) {real, imag} */,
  {32'hbf525ca1, 32'h00000000} /* (10, 28, 12) {real, imag} */,
  {32'hbf083bf0, 32'h00000000} /* (10, 28, 11) {real, imag} */,
  {32'h3eb5de11, 32'h00000000} /* (10, 28, 10) {real, imag} */,
  {32'h3f2e0e35, 32'h00000000} /* (10, 28, 9) {real, imag} */,
  {32'h3ec8b36f, 32'h00000000} /* (10, 28, 8) {real, imag} */,
  {32'h3f402725, 32'h00000000} /* (10, 28, 7) {real, imag} */,
  {32'h3f6eda87, 32'h00000000} /* (10, 28, 6) {real, imag} */,
  {32'h3f884bd9, 32'h00000000} /* (10, 28, 5) {real, imag} */,
  {32'h3fc92b48, 32'h00000000} /* (10, 28, 4) {real, imag} */,
  {32'h3f8c2bd8, 32'h00000000} /* (10, 28, 3) {real, imag} */,
  {32'h3f2afa63, 32'h00000000} /* (10, 28, 2) {real, imag} */,
  {32'h3f9b9d5c, 32'h00000000} /* (10, 28, 1) {real, imag} */,
  {32'h3f41c077, 32'h00000000} /* (10, 28, 0) {real, imag} */,
  {32'h3f268994, 32'h00000000} /* (10, 27, 31) {real, imag} */,
  {32'h3f72df1a, 32'h00000000} /* (10, 27, 30) {real, imag} */,
  {32'h3fc8b539, 32'h00000000} /* (10, 27, 29) {real, imag} */,
  {32'h3f5b06c0, 32'h00000000} /* (10, 27, 28) {real, imag} */,
  {32'h3fd7071e, 32'h00000000} /* (10, 27, 27) {real, imag} */,
  {32'h3fe37083, 32'h00000000} /* (10, 27, 26) {real, imag} */,
  {32'h3fb13aec, 32'h00000000} /* (10, 27, 25) {real, imag} */,
  {32'h3fcc42d5, 32'h00000000} /* (10, 27, 24) {real, imag} */,
  {32'h3fcbbeb6, 32'h00000000} /* (10, 27, 23) {real, imag} */,
  {32'h3fa4bfc8, 32'h00000000} /* (10, 27, 22) {real, imag} */,
  {32'hbdef6fd2, 32'h00000000} /* (10, 27, 21) {real, imag} */,
  {32'hbf82b21d, 32'h00000000} /* (10, 27, 20) {real, imag} */,
  {32'hbf9dd943, 32'h00000000} /* (10, 27, 19) {real, imag} */,
  {32'hbf843c51, 32'h00000000} /* (10, 27, 18) {real, imag} */,
  {32'hbfa910b8, 32'h00000000} /* (10, 27, 17) {real, imag} */,
  {32'hbfcb29d8, 32'h00000000} /* (10, 27, 16) {real, imag} */,
  {32'hbfa6b12e, 32'h00000000} /* (10, 27, 15) {real, imag} */,
  {32'hbf83ac30, 32'h00000000} /* (10, 27, 14) {real, imag} */,
  {32'hbf3a17fa, 32'h00000000} /* (10, 27, 13) {real, imag} */,
  {32'hbf1cd934, 32'h00000000} /* (10, 27, 12) {real, imag} */,
  {32'hbf5b87e1, 32'h00000000} /* (10, 27, 11) {real, imag} */,
  {32'hbd5e5a8e, 32'h00000000} /* (10, 27, 10) {real, imag} */,
  {32'h3f56548c, 32'h00000000} /* (10, 27, 9) {real, imag} */,
  {32'h3ef95f8e, 32'h00000000} /* (10, 27, 8) {real, imag} */,
  {32'h3f58fc48, 32'h00000000} /* (10, 27, 7) {real, imag} */,
  {32'h3f6c4ff1, 32'h00000000} /* (10, 27, 6) {real, imag} */,
  {32'h3fba35ab, 32'h00000000} /* (10, 27, 5) {real, imag} */,
  {32'h3fdd9506, 32'h00000000} /* (10, 27, 4) {real, imag} */,
  {32'h3f65642c, 32'h00000000} /* (10, 27, 3) {real, imag} */,
  {32'h3f46f575, 32'h00000000} /* (10, 27, 2) {real, imag} */,
  {32'h3f89d965, 32'h00000000} /* (10, 27, 1) {real, imag} */,
  {32'h3f7c0375, 32'h00000000} /* (10, 27, 0) {real, imag} */,
  {32'h3edd25d3, 32'h00000000} /* (10, 26, 31) {real, imag} */,
  {32'h3f615518, 32'h00000000} /* (10, 26, 30) {real, imag} */,
  {32'h3fde4ff0, 32'h00000000} /* (10, 26, 29) {real, imag} */,
  {32'h3f47b60c, 32'h00000000} /* (10, 26, 28) {real, imag} */,
  {32'h3f6996a2, 32'h00000000} /* (10, 26, 27) {real, imag} */,
  {32'h3f8614b7, 32'h00000000} /* (10, 26, 26) {real, imag} */,
  {32'h3fda562e, 32'h00000000} /* (10, 26, 25) {real, imag} */,
  {32'h3fbd7e23, 32'h00000000} /* (10, 26, 24) {real, imag} */,
  {32'h3f19dfb3, 32'h00000000} /* (10, 26, 23) {real, imag} */,
  {32'h3f5aedce, 32'h00000000} /* (10, 26, 22) {real, imag} */,
  {32'h3dbc2420, 32'h00000000} /* (10, 26, 21) {real, imag} */,
  {32'hbf63dfde, 32'h00000000} /* (10, 26, 20) {real, imag} */,
  {32'hbf93420f, 32'h00000000} /* (10, 26, 19) {real, imag} */,
  {32'hbf687c72, 32'h00000000} /* (10, 26, 18) {real, imag} */,
  {32'hbfc3b460, 32'h00000000} /* (10, 26, 17) {real, imag} */,
  {32'hbfda5db5, 32'h00000000} /* (10, 26, 16) {real, imag} */,
  {32'hbf6764e2, 32'h00000000} /* (10, 26, 15) {real, imag} */,
  {32'hbf155062, 32'h00000000} /* (10, 26, 14) {real, imag} */,
  {32'hbf48ffb4, 32'h00000000} /* (10, 26, 13) {real, imag} */,
  {32'hbf45bfa3, 32'h00000000} /* (10, 26, 12) {real, imag} */,
  {32'hbeb20b96, 32'h00000000} /* (10, 26, 11) {real, imag} */,
  {32'h3eaf43d9, 32'h00000000} /* (10, 26, 10) {real, imag} */,
  {32'h3fb56ad6, 32'h00000000} /* (10, 26, 9) {real, imag} */,
  {32'h3f964459, 32'h00000000} /* (10, 26, 8) {real, imag} */,
  {32'h3f97f8b9, 32'h00000000} /* (10, 26, 7) {real, imag} */,
  {32'h3f4a5568, 32'h00000000} /* (10, 26, 6) {real, imag} */,
  {32'h3f84953f, 32'h00000000} /* (10, 26, 5) {real, imag} */,
  {32'h3f7632ef, 32'h00000000} /* (10, 26, 4) {real, imag} */,
  {32'h3f63a071, 32'h00000000} /* (10, 26, 3) {real, imag} */,
  {32'h3fa322e2, 32'h00000000} /* (10, 26, 2) {real, imag} */,
  {32'h3f787ef9, 32'h00000000} /* (10, 26, 1) {real, imag} */,
  {32'h3f48f6b9, 32'h00000000} /* (10, 26, 0) {real, imag} */,
  {32'h3ebc45f9, 32'h00000000} /* (10, 25, 31) {real, imag} */,
  {32'h3edb28e6, 32'h00000000} /* (10, 25, 30) {real, imag} */,
  {32'h3f89d8b4, 32'h00000000} /* (10, 25, 29) {real, imag} */,
  {32'h3f84a13d, 32'h00000000} /* (10, 25, 28) {real, imag} */,
  {32'h3ec9712e, 32'h00000000} /* (10, 25, 27) {real, imag} */,
  {32'h3ee7e452, 32'h00000000} /* (10, 25, 26) {real, imag} */,
  {32'h3fbbc326, 32'h00000000} /* (10, 25, 25) {real, imag} */,
  {32'h3f7c0b06, 32'h00000000} /* (10, 25, 24) {real, imag} */,
  {32'h3e9fb3ab, 32'h00000000} /* (10, 25, 23) {real, imag} */,
  {32'h3f22402e, 32'h00000000} /* (10, 25, 22) {real, imag} */,
  {32'h3ebb6361, 32'h00000000} /* (10, 25, 21) {real, imag} */,
  {32'hbebc3ff2, 32'h00000000} /* (10, 25, 20) {real, imag} */,
  {32'hbf3a9dfa, 32'h00000000} /* (10, 25, 19) {real, imag} */,
  {32'hbf694d4b, 32'h00000000} /* (10, 25, 18) {real, imag} */,
  {32'hbfe4dc1a, 32'h00000000} /* (10, 25, 17) {real, imag} */,
  {32'hbfbc2d23, 32'h00000000} /* (10, 25, 16) {real, imag} */,
  {32'hbf37e860, 32'h00000000} /* (10, 25, 15) {real, imag} */,
  {32'hbf21b489, 32'h00000000} /* (10, 25, 14) {real, imag} */,
  {32'hbf1b8823, 32'h00000000} /* (10, 25, 13) {real, imag} */,
  {32'hbf3d7d19, 32'h00000000} /* (10, 25, 12) {real, imag} */,
  {32'hbeaa1fa8, 32'h00000000} /* (10, 25, 11) {real, imag} */,
  {32'h3f06a423, 32'h00000000} /* (10, 25, 10) {real, imag} */,
  {32'h3fa7a7f5, 32'h00000000} /* (10, 25, 9) {real, imag} */,
  {32'h3fa63ed2, 32'h00000000} /* (10, 25, 8) {real, imag} */,
  {32'h3fa42589, 32'h00000000} /* (10, 25, 7) {real, imag} */,
  {32'h3fa29ed8, 32'h00000000} /* (10, 25, 6) {real, imag} */,
  {32'h3fc37d98, 32'h00000000} /* (10, 25, 5) {real, imag} */,
  {32'h3fa59e5a, 32'h00000000} /* (10, 25, 4) {real, imag} */,
  {32'h3f6dc2bd, 32'h00000000} /* (10, 25, 3) {real, imag} */,
  {32'h3f874b86, 32'h00000000} /* (10, 25, 2) {real, imag} */,
  {32'h3f3e30e2, 32'h00000000} /* (10, 25, 1) {real, imag} */,
  {32'h3eef3145, 32'h00000000} /* (10, 25, 0) {real, imag} */,
  {32'h3e220912, 32'h00000000} /* (10, 24, 31) {real, imag} */,
  {32'h3ef154c9, 32'h00000000} /* (10, 24, 30) {real, imag} */,
  {32'h3f3e6919, 32'h00000000} /* (10, 24, 29) {real, imag} */,
  {32'h3f855ba1, 32'h00000000} /* (10, 24, 28) {real, imag} */,
  {32'h3f71ac4a, 32'h00000000} /* (10, 24, 27) {real, imag} */,
  {32'h3f1ff70c, 32'h00000000} /* (10, 24, 26) {real, imag} */,
  {32'h3f58a88e, 32'h00000000} /* (10, 24, 25) {real, imag} */,
  {32'h3f17ac59, 32'h00000000} /* (10, 24, 24) {real, imag} */,
  {32'h3e951a55, 32'h00000000} /* (10, 24, 23) {real, imag} */,
  {32'h3ebc3bd0, 32'h00000000} /* (10, 24, 22) {real, imag} */,
  {32'hbd98de32, 32'h00000000} /* (10, 24, 21) {real, imag} */,
  {32'hbfb885f4, 32'h00000000} /* (10, 24, 20) {real, imag} */,
  {32'hbf855ba7, 32'h00000000} /* (10, 24, 19) {real, imag} */,
  {32'hbf32ac1b, 32'h00000000} /* (10, 24, 18) {real, imag} */,
  {32'hbf82fbe5, 32'h00000000} /* (10, 24, 17) {real, imag} */,
  {32'hbf218f93, 32'h00000000} /* (10, 24, 16) {real, imag} */,
  {32'hbf17da06, 32'h00000000} /* (10, 24, 15) {real, imag} */,
  {32'hbec87c48, 32'h00000000} /* (10, 24, 14) {real, imag} */,
  {32'hbed81d40, 32'h00000000} /* (10, 24, 13) {real, imag} */,
  {32'hbf9bcda8, 32'h00000000} /* (10, 24, 12) {real, imag} */,
  {32'hbf70d889, 32'h00000000} /* (10, 24, 11) {real, imag} */,
  {32'h3f512815, 32'h00000000} /* (10, 24, 10) {real, imag} */,
  {32'h3fae136e, 32'h00000000} /* (10, 24, 9) {real, imag} */,
  {32'h3fa7a9c8, 32'h00000000} /* (10, 24, 8) {real, imag} */,
  {32'h3fd42f22, 32'h00000000} /* (10, 24, 7) {real, imag} */,
  {32'h3fb392b2, 32'h00000000} /* (10, 24, 6) {real, imag} */,
  {32'h3f647aac, 32'h00000000} /* (10, 24, 5) {real, imag} */,
  {32'h3f684a1e, 32'h00000000} /* (10, 24, 4) {real, imag} */,
  {32'h3f9a0168, 32'h00000000} /* (10, 24, 3) {real, imag} */,
  {32'h3fc4d68a, 32'h00000000} /* (10, 24, 2) {real, imag} */,
  {32'h3f4acce9, 32'h00000000} /* (10, 24, 1) {real, imag} */,
  {32'h3f11ca2a, 32'h00000000} /* (10, 24, 0) {real, imag} */,
  {32'h3bcf9544, 32'h00000000} /* (10, 23, 31) {real, imag} */,
  {32'h3ead148a, 32'h00000000} /* (10, 23, 30) {real, imag} */,
  {32'h3f114a9a, 32'h00000000} /* (10, 23, 29) {real, imag} */,
  {32'h3f3f953d, 32'h00000000} /* (10, 23, 28) {real, imag} */,
  {32'h3f33b582, 32'h00000000} /* (10, 23, 27) {real, imag} */,
  {32'h3f50150c, 32'h00000000} /* (10, 23, 26) {real, imag} */,
  {32'h3f369cfc, 32'h00000000} /* (10, 23, 25) {real, imag} */,
  {32'h3f20141c, 32'h00000000} /* (10, 23, 24) {real, imag} */,
  {32'h3e74cfcc, 32'h00000000} /* (10, 23, 23) {real, imag} */,
  {32'h3ee2d6a4, 32'h00000000} /* (10, 23, 22) {real, imag} */,
  {32'h3e4e889a, 32'h00000000} /* (10, 23, 21) {real, imag} */,
  {32'hbfd42330, 32'h00000000} /* (10, 23, 20) {real, imag} */,
  {32'hbfe31890, 32'h00000000} /* (10, 23, 19) {real, imag} */,
  {32'hbfb62a0e, 32'h00000000} /* (10, 23, 18) {real, imag} */,
  {32'hbf90316e, 32'h00000000} /* (10, 23, 17) {real, imag} */,
  {32'hbebc980b, 32'h00000000} /* (10, 23, 16) {real, imag} */,
  {32'hbe2ad179, 32'h00000000} /* (10, 23, 15) {real, imag} */,
  {32'hbe764bca, 32'h00000000} /* (10, 23, 14) {real, imag} */,
  {32'hbf059303, 32'h00000000} /* (10, 23, 13) {real, imag} */,
  {32'hbf7f8eca, 32'h00000000} /* (10, 23, 12) {real, imag} */,
  {32'hbf967d2e, 32'h00000000} /* (10, 23, 11) {real, imag} */,
  {32'h3edf5aa1, 32'h00000000} /* (10, 23, 10) {real, imag} */,
  {32'h3fb5e2f3, 32'h00000000} /* (10, 23, 9) {real, imag} */,
  {32'h3f9e5963, 32'h00000000} /* (10, 23, 8) {real, imag} */,
  {32'h3fc54b05, 32'h00000000} /* (10, 23, 7) {real, imag} */,
  {32'h3fc395f7, 32'h00000000} /* (10, 23, 6) {real, imag} */,
  {32'h3f3b69e8, 32'h00000000} /* (10, 23, 5) {real, imag} */,
  {32'h3f6a0c21, 32'h00000000} /* (10, 23, 4) {real, imag} */,
  {32'h3f9f112f, 32'h00000000} /* (10, 23, 3) {real, imag} */,
  {32'h3f98a457, 32'h00000000} /* (10, 23, 2) {real, imag} */,
  {32'h3f8aeda7, 32'h00000000} /* (10, 23, 1) {real, imag} */,
  {32'h3f0f1c66, 32'h00000000} /* (10, 23, 0) {real, imag} */,
  {32'h3e5b90cd, 32'h00000000} /* (10, 22, 31) {real, imag} */,
  {32'h3f52524c, 32'h00000000} /* (10, 22, 30) {real, imag} */,
  {32'h3f2edf16, 32'h00000000} /* (10, 22, 29) {real, imag} */,
  {32'h3f347c00, 32'h00000000} /* (10, 22, 28) {real, imag} */,
  {32'h3ee097d8, 32'h00000000} /* (10, 22, 27) {real, imag} */,
  {32'h3f762310, 32'h00000000} /* (10, 22, 26) {real, imag} */,
  {32'h3f766901, 32'h00000000} /* (10, 22, 25) {real, imag} */,
  {32'h3f22acfc, 32'h00000000} /* (10, 22, 24) {real, imag} */,
  {32'h3f1ade92, 32'h00000000} /* (10, 22, 23) {real, imag} */,
  {32'h3f1c2217, 32'h00000000} /* (10, 22, 22) {real, imag} */,
  {32'h3ed95dc2, 32'h00000000} /* (10, 22, 21) {real, imag} */,
  {32'hbfa1aa3f, 32'h00000000} /* (10, 22, 20) {real, imag} */,
  {32'hbfe05220, 32'h00000000} /* (10, 22, 19) {real, imag} */,
  {32'hbf9fa655, 32'h00000000} /* (10, 22, 18) {real, imag} */,
  {32'hbf4785eb, 32'h00000000} /* (10, 22, 17) {real, imag} */,
  {32'hbef5ef16, 32'h00000000} /* (10, 22, 16) {real, imag} */,
  {32'hbf005562, 32'h00000000} /* (10, 22, 15) {real, imag} */,
  {32'hbf9cd0ab, 32'h00000000} /* (10, 22, 14) {real, imag} */,
  {32'hbf9e12b5, 32'h00000000} /* (10, 22, 13) {real, imag} */,
  {32'hbf101e2e, 32'h00000000} /* (10, 22, 12) {real, imag} */,
  {32'hbf18f8c7, 32'h00000000} /* (10, 22, 11) {real, imag} */,
  {32'h3dd9a703, 32'h00000000} /* (10, 22, 10) {real, imag} */,
  {32'h3efe6fe9, 32'h00000000} /* (10, 22, 9) {real, imag} */,
  {32'h3eee8aba, 32'h00000000} /* (10, 22, 8) {real, imag} */,
  {32'h3f3cc867, 32'h00000000} /* (10, 22, 7) {real, imag} */,
  {32'h3f8874e9, 32'h00000000} /* (10, 22, 6) {real, imag} */,
  {32'h3f62b7f8, 32'h00000000} /* (10, 22, 5) {real, imag} */,
  {32'h3f33f93a, 32'h00000000} /* (10, 22, 4) {real, imag} */,
  {32'h3f9292ab, 32'h00000000} /* (10, 22, 3) {real, imag} */,
  {32'h3fcf9352, 32'h00000000} /* (10, 22, 2) {real, imag} */,
  {32'h3f83bd35, 32'h00000000} /* (10, 22, 1) {real, imag} */,
  {32'h3f0de10a, 32'h00000000} /* (10, 22, 0) {real, imag} */,
  {32'h3e17cdde, 32'h00000000} /* (10, 21, 31) {real, imag} */,
  {32'h3f1e340f, 32'h00000000} /* (10, 21, 30) {real, imag} */,
  {32'h3eb53a81, 32'h00000000} /* (10, 21, 29) {real, imag} */,
  {32'h3e5f51f3, 32'h00000000} /* (10, 21, 28) {real, imag} */,
  {32'h3e8abb0c, 32'h00000000} /* (10, 21, 27) {real, imag} */,
  {32'h3edae6b6, 32'h00000000} /* (10, 21, 26) {real, imag} */,
  {32'h3e60dd63, 32'h00000000} /* (10, 21, 25) {real, imag} */,
  {32'h3e34f811, 32'h00000000} /* (10, 21, 24) {real, imag} */,
  {32'h3eb78c0e, 32'h00000000} /* (10, 21, 23) {real, imag} */,
  {32'h3f2410bf, 32'h00000000} /* (10, 21, 22) {real, imag} */,
  {32'h3f5a812f, 32'h00000000} /* (10, 21, 21) {real, imag} */,
  {32'hbefe49b6, 32'h00000000} /* (10, 21, 20) {real, imag} */,
  {32'hbf46a787, 32'h00000000} /* (10, 21, 19) {real, imag} */,
  {32'hbea7fdc7, 32'h00000000} /* (10, 21, 18) {real, imag} */,
  {32'hbe49bd0a, 32'h00000000} /* (10, 21, 17) {real, imag} */,
  {32'h3e4a8c5b, 32'h00000000} /* (10, 21, 16) {real, imag} */,
  {32'h3d4435d1, 32'h00000000} /* (10, 21, 15) {real, imag} */,
  {32'hbf2f7485, 32'h00000000} /* (10, 21, 14) {real, imag} */,
  {32'hbf0eee1e, 32'h00000000} /* (10, 21, 13) {real, imag} */,
  {32'hbe3c22a0, 32'h00000000} /* (10, 21, 12) {real, imag} */,
  {32'hbe331a0a, 32'h00000000} /* (10, 21, 11) {real, imag} */,
  {32'hbc8355a4, 32'h00000000} /* (10, 21, 10) {real, imag} */,
  {32'h3e724057, 32'h00000000} /* (10, 21, 9) {real, imag} */,
  {32'hbcce6984, 32'h00000000} /* (10, 21, 8) {real, imag} */,
  {32'hbe216c73, 32'h00000000} /* (10, 21, 7) {real, imag} */,
  {32'h3e577972, 32'h00000000} /* (10, 21, 6) {real, imag} */,
  {32'h3f0ece17, 32'h00000000} /* (10, 21, 5) {real, imag} */,
  {32'h3eab59d5, 32'h00000000} /* (10, 21, 4) {real, imag} */,
  {32'h3e8b16b4, 32'h00000000} /* (10, 21, 3) {real, imag} */,
  {32'h3f3ca59e, 32'h00000000} /* (10, 21, 2) {real, imag} */,
  {32'h3ea1b752, 32'h00000000} /* (10, 21, 1) {real, imag} */,
  {32'h3e8b639f, 32'h00000000} /* (10, 21, 0) {real, imag} */,
  {32'hbe805d4c, 32'h00000000} /* (10, 20, 31) {real, imag} */,
  {32'hbf19430a, 32'h00000000} /* (10, 20, 30) {real, imag} */,
  {32'hbeeccc1e, 32'h00000000} /* (10, 20, 29) {real, imag} */,
  {32'hbea04f5b, 32'h00000000} /* (10, 20, 28) {real, imag} */,
  {32'hbe125e50, 32'h00000000} /* (10, 20, 27) {real, imag} */,
  {32'hbe8a8752, 32'h00000000} /* (10, 20, 26) {real, imag} */,
  {32'hbf5c8eeb, 32'h00000000} /* (10, 20, 25) {real, imag} */,
  {32'hbf8e6eaf, 32'h00000000} /* (10, 20, 24) {real, imag} */,
  {32'hbf430a3d, 32'h00000000} /* (10, 20, 23) {real, imag} */,
  {32'hbf202761, 32'h00000000} /* (10, 20, 22) {real, imag} */,
  {32'h3e2a3b5d, 32'h00000000} /* (10, 20, 21) {real, imag} */,
  {32'h3f334343, 32'h00000000} /* (10, 20, 20) {real, imag} */,
  {32'h3f4363fd, 32'h00000000} /* (10, 20, 19) {real, imag} */,
  {32'h3ea8a190, 32'h00000000} /* (10, 20, 18) {real, imag} */,
  {32'h3ebaabcb, 32'h00000000} /* (10, 20, 17) {real, imag} */,
  {32'h3f918690, 32'h00000000} /* (10, 20, 16) {real, imag} */,
  {32'h3f9441cb, 32'h00000000} /* (10, 20, 15) {real, imag} */,
  {32'h3f72812b, 32'h00000000} /* (10, 20, 14) {real, imag} */,
  {32'h3f5ac004, 32'h00000000} /* (10, 20, 13) {real, imag} */,
  {32'h3f44cdb8, 32'h00000000} /* (10, 20, 12) {real, imag} */,
  {32'h3f02e5f6, 32'h00000000} /* (10, 20, 11) {real, imag} */,
  {32'hbe8e50b2, 32'h00000000} /* (10, 20, 10) {real, imag} */,
  {32'hbe4451fc, 32'h00000000} /* (10, 20, 9) {real, imag} */,
  {32'hbf2bcb58, 32'h00000000} /* (10, 20, 8) {real, imag} */,
  {32'hbf7acc5e, 32'h00000000} /* (10, 20, 7) {real, imag} */,
  {32'hbf293c17, 32'h00000000} /* (10, 20, 6) {real, imag} */,
  {32'hbf1abf29, 32'h00000000} /* (10, 20, 5) {real, imag} */,
  {32'hbee2afb2, 32'h00000000} /* (10, 20, 4) {real, imag} */,
  {32'hbf564196, 32'h00000000} /* (10, 20, 3) {real, imag} */,
  {32'hbf3767d7, 32'h00000000} /* (10, 20, 2) {real, imag} */,
  {32'hbf914785, 32'h00000000} /* (10, 20, 1) {real, imag} */,
  {32'hbf0e5ba9, 32'h00000000} /* (10, 20, 0) {real, imag} */,
  {32'hbf3de97f, 32'h00000000} /* (10, 19, 31) {real, imag} */,
  {32'hbfb9249d, 32'h00000000} /* (10, 19, 30) {real, imag} */,
  {32'hbf8deae2, 32'h00000000} /* (10, 19, 29) {real, imag} */,
  {32'hbf5fc373, 32'h00000000} /* (10, 19, 28) {real, imag} */,
  {32'hbf29e108, 32'h00000000} /* (10, 19, 27) {real, imag} */,
  {32'hbf361bc3, 32'h00000000} /* (10, 19, 26) {real, imag} */,
  {32'hbf406929, 32'h00000000} /* (10, 19, 25) {real, imag} */,
  {32'hbf91401e, 32'h00000000} /* (10, 19, 24) {real, imag} */,
  {32'hbf6fc7bc, 32'h00000000} /* (10, 19, 23) {real, imag} */,
  {32'hbf9cc7c4, 32'h00000000} /* (10, 19, 22) {real, imag} */,
  {32'hbef7787e, 32'h00000000} /* (10, 19, 21) {real, imag} */,
  {32'h3eeb628f, 32'h00000000} /* (10, 19, 20) {real, imag} */,
  {32'h3ef5f598, 32'h00000000} /* (10, 19, 19) {real, imag} */,
  {32'h3e89b52d, 32'h00000000} /* (10, 19, 18) {real, imag} */,
  {32'h3f3c02a3, 32'h00000000} /* (10, 19, 17) {real, imag} */,
  {32'h3fb765b5, 32'h00000000} /* (10, 19, 16) {real, imag} */,
  {32'h3fbf0cd6, 32'h00000000} /* (10, 19, 15) {real, imag} */,
  {32'h3f992d03, 32'h00000000} /* (10, 19, 14) {real, imag} */,
  {32'h3f54e78f, 32'h00000000} /* (10, 19, 13) {real, imag} */,
  {32'h3f6dec54, 32'h00000000} /* (10, 19, 12) {real, imag} */,
  {32'h3f1e9f38, 32'h00000000} /* (10, 19, 11) {real, imag} */,
  {32'hbe35a147, 32'h00000000} /* (10, 19, 10) {real, imag} */,
  {32'hbe9cb7f0, 32'h00000000} /* (10, 19, 9) {real, imag} */,
  {32'hbf2761c4, 32'h00000000} /* (10, 19, 8) {real, imag} */,
  {32'hbf7be702, 32'h00000000} /* (10, 19, 7) {real, imag} */,
  {32'hbf22c02d, 32'h00000000} /* (10, 19, 6) {real, imag} */,
  {32'hbf835437, 32'h00000000} /* (10, 19, 5) {real, imag} */,
  {32'hbf73cef4, 32'h00000000} /* (10, 19, 4) {real, imag} */,
  {32'hbf33207f, 32'h00000000} /* (10, 19, 3) {real, imag} */,
  {32'hbf67cd27, 32'h00000000} /* (10, 19, 2) {real, imag} */,
  {32'hbf92407a, 32'h00000000} /* (10, 19, 1) {real, imag} */,
  {32'hbf4999b3, 32'h00000000} /* (10, 19, 0) {real, imag} */,
  {32'hbf3208fc, 32'h00000000} /* (10, 18, 31) {real, imag} */,
  {32'hbfad2f20, 32'h00000000} /* (10, 18, 30) {real, imag} */,
  {32'hbf622499, 32'h00000000} /* (10, 18, 29) {real, imag} */,
  {32'hbfb5f808, 32'h00000000} /* (10, 18, 28) {real, imag} */,
  {32'hbf990e9c, 32'h00000000} /* (10, 18, 27) {real, imag} */,
  {32'hbf447a28, 32'h00000000} /* (10, 18, 26) {real, imag} */,
  {32'hbf288878, 32'h00000000} /* (10, 18, 25) {real, imag} */,
  {32'hbf8b909c, 32'h00000000} /* (10, 18, 24) {real, imag} */,
  {32'hbf26c906, 32'h00000000} /* (10, 18, 23) {real, imag} */,
  {32'hbf39b00d, 32'h00000000} /* (10, 18, 22) {real, imag} */,
  {32'hbf1d78d0, 32'h00000000} /* (10, 18, 21) {real, imag} */,
  {32'h3ed82141, 32'h00000000} /* (10, 18, 20) {real, imag} */,
  {32'h3eb00b6d, 32'h00000000} /* (10, 18, 19) {real, imag} */,
  {32'h3e5089fd, 32'h00000000} /* (10, 18, 18) {real, imag} */,
  {32'h3eeddd65, 32'h00000000} /* (10, 18, 17) {real, imag} */,
  {32'h3f82d5b6, 32'h00000000} /* (10, 18, 16) {real, imag} */,
  {32'h3fab0371, 32'h00000000} /* (10, 18, 15) {real, imag} */,
  {32'h3f60d21c, 32'h00000000} /* (10, 18, 14) {real, imag} */,
  {32'h3f879a1f, 32'h00000000} /* (10, 18, 13) {real, imag} */,
  {32'h3fb95dc4, 32'h00000000} /* (10, 18, 12) {real, imag} */,
  {32'h3f70e861, 32'h00000000} /* (10, 18, 11) {real, imag} */,
  {32'hbefca91d, 32'h00000000} /* (10, 18, 10) {real, imag} */,
  {32'hbf2d3531, 32'h00000000} /* (10, 18, 9) {real, imag} */,
  {32'hbfaaafed, 32'h00000000} /* (10, 18, 8) {real, imag} */,
  {32'hbfe3b8e2, 32'h00000000} /* (10, 18, 7) {real, imag} */,
  {32'hbfa50cf3, 32'h00000000} /* (10, 18, 6) {real, imag} */,
  {32'hbf90c6e6, 32'h00000000} /* (10, 18, 5) {real, imag} */,
  {32'hbf8294a0, 32'h00000000} /* (10, 18, 4) {real, imag} */,
  {32'hbf82139a, 32'h00000000} /* (10, 18, 3) {real, imag} */,
  {32'hbf5ec2ff, 32'h00000000} /* (10, 18, 2) {real, imag} */,
  {32'hbf5af0e5, 32'h00000000} /* (10, 18, 1) {real, imag} */,
  {32'hbf32fa6c, 32'h00000000} /* (10, 18, 0) {real, imag} */,
  {32'hbe4c3b17, 32'h00000000} /* (10, 17, 31) {real, imag} */,
  {32'hbf2293bf, 32'h00000000} /* (10, 17, 30) {real, imag} */,
  {32'hbf41684d, 32'h00000000} /* (10, 17, 29) {real, imag} */,
  {32'hbf96670c, 32'h00000000} /* (10, 17, 28) {real, imag} */,
  {32'hbfb1f6c6, 32'h00000000} /* (10, 17, 27) {real, imag} */,
  {32'hbf8ab96a, 32'h00000000} /* (10, 17, 26) {real, imag} */,
  {32'hbf7bf891, 32'h00000000} /* (10, 17, 25) {real, imag} */,
  {32'hbf9db351, 32'h00000000} /* (10, 17, 24) {real, imag} */,
  {32'hbf7a478b, 32'h00000000} /* (10, 17, 23) {real, imag} */,
  {32'hbf8cd7de, 32'h00000000} /* (10, 17, 22) {real, imag} */,
  {32'hbf6bcfd4, 32'h00000000} /* (10, 17, 21) {real, imag} */,
  {32'h3eda6eb8, 32'h00000000} /* (10, 17, 20) {real, imag} */,
  {32'h3f5d5e0e, 32'h00000000} /* (10, 17, 19) {real, imag} */,
  {32'h3f9c183f, 32'h00000000} /* (10, 17, 18) {real, imag} */,
  {32'h3f60dad6, 32'h00000000} /* (10, 17, 17) {real, imag} */,
  {32'h3f28bab3, 32'h00000000} /* (10, 17, 16) {real, imag} */,
  {32'h3f676bd3, 32'h00000000} /* (10, 17, 15) {real, imag} */,
  {32'h3f992bb0, 32'h00000000} /* (10, 17, 14) {real, imag} */,
  {32'h3f967a58, 32'h00000000} /* (10, 17, 13) {real, imag} */,
  {32'h3fa32300, 32'h00000000} /* (10, 17, 12) {real, imag} */,
  {32'h3f40d708, 32'h00000000} /* (10, 17, 11) {real, imag} */,
  {32'hbf84e1d5, 32'h00000000} /* (10, 17, 10) {real, imag} */,
  {32'hbfa08551, 32'h00000000} /* (10, 17, 9) {real, imag} */,
  {32'hbfae1c6d, 32'h00000000} /* (10, 17, 8) {real, imag} */,
  {32'hbfb5c8ee, 32'h00000000} /* (10, 17, 7) {real, imag} */,
  {32'hbfdf58cf, 32'h00000000} /* (10, 17, 6) {real, imag} */,
  {32'hbf6be68b, 32'h00000000} /* (10, 17, 5) {real, imag} */,
  {32'hbf3a6e2a, 32'h00000000} /* (10, 17, 4) {real, imag} */,
  {32'hbfb0f5bd, 32'h00000000} /* (10, 17, 3) {real, imag} */,
  {32'hbfcc2fd7, 32'h00000000} /* (10, 17, 2) {real, imag} */,
  {32'hbf62528f, 32'h00000000} /* (10, 17, 1) {real, imag} */,
  {32'hbedde3b6, 32'h00000000} /* (10, 17, 0) {real, imag} */,
  {32'hbe4ba647, 32'h00000000} /* (10, 16, 31) {real, imag} */,
  {32'hbf65b3c7, 32'h00000000} /* (10, 16, 30) {real, imag} */,
  {32'hbf4f7679, 32'h00000000} /* (10, 16, 29) {real, imag} */,
  {32'hbf9b5652, 32'h00000000} /* (10, 16, 28) {real, imag} */,
  {32'hbfc016f0, 32'h00000000} /* (10, 16, 27) {real, imag} */,
  {32'hbf7c6420, 32'h00000000} /* (10, 16, 26) {real, imag} */,
  {32'hbf546fde, 32'h00000000} /* (10, 16, 25) {real, imag} */,
  {32'hbf7d4f26, 32'h00000000} /* (10, 16, 24) {real, imag} */,
  {32'hbf8181e8, 32'h00000000} /* (10, 16, 23) {real, imag} */,
  {32'hbf4c6b2a, 32'h00000000} /* (10, 16, 22) {real, imag} */,
  {32'hbd9febe8, 32'h00000000} /* (10, 16, 21) {real, imag} */,
  {32'h3f177bb0, 32'h00000000} /* (10, 16, 20) {real, imag} */,
  {32'h3f80743b, 32'h00000000} /* (10, 16, 19) {real, imag} */,
  {32'h3fa40d0f, 32'h00000000} /* (10, 16, 18) {real, imag} */,
  {32'h3f80d057, 32'h00000000} /* (10, 16, 17) {real, imag} */,
  {32'h3f901f2d, 32'h00000000} /* (10, 16, 16) {real, imag} */,
  {32'h3f58a3c8, 32'h00000000} /* (10, 16, 15) {real, imag} */,
  {32'h3f9fbfc9, 32'h00000000} /* (10, 16, 14) {real, imag} */,
  {32'h3fa7ab2c, 32'h00000000} /* (10, 16, 13) {real, imag} */,
  {32'h3f5243da, 32'h00000000} /* (10, 16, 12) {real, imag} */,
  {32'h3ec600a2, 32'h00000000} /* (10, 16, 11) {real, imag} */,
  {32'hbf771d9a, 32'h00000000} /* (10, 16, 10) {real, imag} */,
  {32'hbf9b4d3b, 32'h00000000} /* (10, 16, 9) {real, imag} */,
  {32'hbf9f78e4, 32'h00000000} /* (10, 16, 8) {real, imag} */,
  {32'hbf5f54c6, 32'h00000000} /* (10, 16, 7) {real, imag} */,
  {32'hbf36f36d, 32'h00000000} /* (10, 16, 6) {real, imag} */,
  {32'hbe98da97, 32'h00000000} /* (10, 16, 5) {real, imag} */,
  {32'hbef95793, 32'h00000000} /* (10, 16, 4) {real, imag} */,
  {32'hbf8adeb1, 32'h00000000} /* (10, 16, 3) {real, imag} */,
  {32'hbfc88c04, 32'h00000000} /* (10, 16, 2) {real, imag} */,
  {32'hbf63cb1f, 32'h00000000} /* (10, 16, 1) {real, imag} */,
  {32'hbe2b109d, 32'h00000000} /* (10, 16, 0) {real, imag} */,
  {32'hbecbfe39, 32'h00000000} /* (10, 15, 31) {real, imag} */,
  {32'hbf9207ff, 32'h00000000} /* (10, 15, 30) {real, imag} */,
  {32'hbf675af1, 32'h00000000} /* (10, 15, 29) {real, imag} */,
  {32'hbf60c3ca, 32'h00000000} /* (10, 15, 28) {real, imag} */,
  {32'hbf73c722, 32'h00000000} /* (10, 15, 27) {real, imag} */,
  {32'hbf88dcc3, 32'h00000000} /* (10, 15, 26) {real, imag} */,
  {32'hbf5e8f61, 32'h00000000} /* (10, 15, 25) {real, imag} */,
  {32'hbf7d3406, 32'h00000000} /* (10, 15, 24) {real, imag} */,
  {32'hbf5b0791, 32'h00000000} /* (10, 15, 23) {real, imag} */,
  {32'hbe8a3f34, 32'h00000000} /* (10, 15, 22) {real, imag} */,
  {32'h3f4e12ba, 32'h00000000} /* (10, 15, 21) {real, imag} */,
  {32'h3f912941, 32'h00000000} /* (10, 15, 20) {real, imag} */,
  {32'h3f3ef05d, 32'h00000000} /* (10, 15, 19) {real, imag} */,
  {32'h3f959ed8, 32'h00000000} /* (10, 15, 18) {real, imag} */,
  {32'h3f7d1639, 32'h00000000} /* (10, 15, 17) {real, imag} */,
  {32'h3f873bc2, 32'h00000000} /* (10, 15, 16) {real, imag} */,
  {32'h3f497e54, 32'h00000000} /* (10, 15, 15) {real, imag} */,
  {32'h3f3e114c, 32'h00000000} /* (10, 15, 14) {real, imag} */,
  {32'h3f591eea, 32'h00000000} /* (10, 15, 13) {real, imag} */,
  {32'h3f61a475, 32'h00000000} /* (10, 15, 12) {real, imag} */,
  {32'h3f065371, 32'h00000000} /* (10, 15, 11) {real, imag} */,
  {32'hbf1e890f, 32'h00000000} /* (10, 15, 10) {real, imag} */,
  {32'hbfa33f0a, 32'h00000000} /* (10, 15, 9) {real, imag} */,
  {32'hbfccd59a, 32'h00000000} /* (10, 15, 8) {real, imag} */,
  {32'hbf9456e4, 32'h00000000} /* (10, 15, 7) {real, imag} */,
  {32'hbf236d95, 32'h00000000} /* (10, 15, 6) {real, imag} */,
  {32'hbf22c61a, 32'h00000000} /* (10, 15, 5) {real, imag} */,
  {32'hbf9214ea, 32'h00000000} /* (10, 15, 4) {real, imag} */,
  {32'hbf8d834e, 32'h00000000} /* (10, 15, 3) {real, imag} */,
  {32'hbfa9705c, 32'h00000000} /* (10, 15, 2) {real, imag} */,
  {32'hbf9f0be9, 32'h00000000} /* (10, 15, 1) {real, imag} */,
  {32'hbf15e129, 32'h00000000} /* (10, 15, 0) {real, imag} */,
  {32'hbed41d03, 32'h00000000} /* (10, 14, 31) {real, imag} */,
  {32'hbf6e24ab, 32'h00000000} /* (10, 14, 30) {real, imag} */,
  {32'hbf4dfeb7, 32'h00000000} /* (10, 14, 29) {real, imag} */,
  {32'hbf5d5a8b, 32'h00000000} /* (10, 14, 28) {real, imag} */,
  {32'hbf3e9f50, 32'h00000000} /* (10, 14, 27) {real, imag} */,
  {32'hbf5fd253, 32'h00000000} /* (10, 14, 26) {real, imag} */,
  {32'hbf8b0200, 32'h00000000} /* (10, 14, 25) {real, imag} */,
  {32'hbf4273e3, 32'h00000000} /* (10, 14, 24) {real, imag} */,
  {32'hbed98e3c, 32'h00000000} /* (10, 14, 23) {real, imag} */,
  {32'hbe634fe8, 32'h00000000} /* (10, 14, 22) {real, imag} */,
  {32'hbe1e80ec, 32'h00000000} /* (10, 14, 21) {real, imag} */,
  {32'h3f15b285, 32'h00000000} /* (10, 14, 20) {real, imag} */,
  {32'h3f37abbb, 32'h00000000} /* (10, 14, 19) {real, imag} */,
  {32'h3f744166, 32'h00000000} /* (10, 14, 18) {real, imag} */,
  {32'h3f6a1d9a, 32'h00000000} /* (10, 14, 17) {real, imag} */,
  {32'h3f3746d3, 32'h00000000} /* (10, 14, 16) {real, imag} */,
  {32'h3f24fb53, 32'h00000000} /* (10, 14, 15) {real, imag} */,
  {32'h3f5995e8, 32'h00000000} /* (10, 14, 14) {real, imag} */,
  {32'h3f6519c3, 32'h00000000} /* (10, 14, 13) {real, imag} */,
  {32'h3f561bf5, 32'h00000000} /* (10, 14, 12) {real, imag} */,
  {32'h3f6e9795, 32'h00000000} /* (10, 14, 11) {real, imag} */,
  {32'hbd836e93, 32'h00000000} /* (10, 14, 10) {real, imag} */,
  {32'hbf8e6a28, 32'h00000000} /* (10, 14, 9) {real, imag} */,
  {32'hbf86d3a8, 32'h00000000} /* (10, 14, 8) {real, imag} */,
  {32'hbf421a74, 32'h00000000} /* (10, 14, 7) {real, imag} */,
  {32'hbf5bbcc3, 32'h00000000} /* (10, 14, 6) {real, imag} */,
  {32'hbf79210c, 32'h00000000} /* (10, 14, 5) {real, imag} */,
  {32'hbf803688, 32'h00000000} /* (10, 14, 4) {real, imag} */,
  {32'hbf61d568, 32'h00000000} /* (10, 14, 3) {real, imag} */,
  {32'hbf31dacb, 32'h00000000} /* (10, 14, 2) {real, imag} */,
  {32'hbfb087f0, 32'h00000000} /* (10, 14, 1) {real, imag} */,
  {32'hbf8f726c, 32'h00000000} /* (10, 14, 0) {real, imag} */,
  {32'hbed9be13, 32'h00000000} /* (10, 13, 31) {real, imag} */,
  {32'hbf3de2bf, 32'h00000000} /* (10, 13, 30) {real, imag} */,
  {32'hbf2a8ac0, 32'h00000000} /* (10, 13, 29) {real, imag} */,
  {32'hbf68343b, 32'h00000000} /* (10, 13, 28) {real, imag} */,
  {32'hbf4599b3, 32'h00000000} /* (10, 13, 27) {real, imag} */,
  {32'hbf4404e8, 32'h00000000} /* (10, 13, 26) {real, imag} */,
  {32'hbf7b428e, 32'h00000000} /* (10, 13, 25) {real, imag} */,
  {32'hbf6f2d95, 32'h00000000} /* (10, 13, 24) {real, imag} */,
  {32'hbf4eda99, 32'h00000000} /* (10, 13, 23) {real, imag} */,
  {32'hbf1c59b7, 32'h00000000} /* (10, 13, 22) {real, imag} */,
  {32'hbe06edfe, 32'h00000000} /* (10, 13, 21) {real, imag} */,
  {32'h3f0c013e, 32'h00000000} /* (10, 13, 20) {real, imag} */,
  {32'h3f75c1ac, 32'h00000000} /* (10, 13, 19) {real, imag} */,
  {32'h3f81a4ad, 32'h00000000} /* (10, 13, 18) {real, imag} */,
  {32'h3f37d606, 32'h00000000} /* (10, 13, 17) {real, imag} */,
  {32'h3f1be264, 32'h00000000} /* (10, 13, 16) {real, imag} */,
  {32'h3f0d0969, 32'h00000000} /* (10, 13, 15) {real, imag} */,
  {32'h3ec5d88a, 32'h00000000} /* (10, 13, 14) {real, imag} */,
  {32'h3f32f76d, 32'h00000000} /* (10, 13, 13) {real, imag} */,
  {32'h3f6075eb, 32'h00000000} /* (10, 13, 12) {real, imag} */,
  {32'h3f7b1498, 32'h00000000} /* (10, 13, 11) {real, imag} */,
  {32'hbd19e984, 32'h00000000} /* (10, 13, 10) {real, imag} */,
  {32'hbf629b44, 32'h00000000} /* (10, 13, 9) {real, imag} */,
  {32'hbf7d2f11, 32'h00000000} /* (10, 13, 8) {real, imag} */,
  {32'hbf93aa0a, 32'h00000000} /* (10, 13, 7) {real, imag} */,
  {32'hbf97f209, 32'h00000000} /* (10, 13, 6) {real, imag} */,
  {32'hbf78f40d, 32'h00000000} /* (10, 13, 5) {real, imag} */,
  {32'hbf38a625, 32'h00000000} /* (10, 13, 4) {real, imag} */,
  {32'hbf6d4378, 32'h00000000} /* (10, 13, 3) {real, imag} */,
  {32'hbecae27e, 32'h00000000} /* (10, 13, 2) {real, imag} */,
  {32'hbf8f3d94, 32'h00000000} /* (10, 13, 1) {real, imag} */,
  {32'hbf7d1474, 32'h00000000} /* (10, 13, 0) {real, imag} */,
  {32'hbf2dc563, 32'h00000000} /* (10, 12, 31) {real, imag} */,
  {32'hbf9107dd, 32'h00000000} /* (10, 12, 30) {real, imag} */,
  {32'hbf5beaff, 32'h00000000} /* (10, 12, 29) {real, imag} */,
  {32'hbf193403, 32'h00000000} /* (10, 12, 28) {real, imag} */,
  {32'hbf138cd1, 32'h00000000} /* (10, 12, 27) {real, imag} */,
  {32'hbf524a0c, 32'h00000000} /* (10, 12, 26) {real, imag} */,
  {32'hbf252108, 32'h00000000} /* (10, 12, 25) {real, imag} */,
  {32'hbf9e8c44, 32'h00000000} /* (10, 12, 24) {real, imag} */,
  {32'hbfa46f94, 32'h00000000} /* (10, 12, 23) {real, imag} */,
  {32'hbf5fcbbe, 32'h00000000} /* (10, 12, 22) {real, imag} */,
  {32'hbeff4c44, 32'h00000000} /* (10, 12, 21) {real, imag} */,
  {32'h3f0dca14, 32'h00000000} /* (10, 12, 20) {real, imag} */,
  {32'h3f9d4176, 32'h00000000} /* (10, 12, 19) {real, imag} */,
  {32'h3f559bd6, 32'h00000000} /* (10, 12, 18) {real, imag} */,
  {32'h3f78f6af, 32'h00000000} /* (10, 12, 17) {real, imag} */,
  {32'h3fa60a33, 32'h00000000} /* (10, 12, 16) {real, imag} */,
  {32'h3f44cb39, 32'h00000000} /* (10, 12, 15) {real, imag} */,
  {32'h3f0e45d7, 32'h00000000} /* (10, 12, 14) {real, imag} */,
  {32'h3f120abf, 32'h00000000} /* (10, 12, 13) {real, imag} */,
  {32'h3f369614, 32'h00000000} /* (10, 12, 12) {real, imag} */,
  {32'h3ea52956, 32'h00000000} /* (10, 12, 11) {real, imag} */,
  {32'hbf1763c1, 32'h00000000} /* (10, 12, 10) {real, imag} */,
  {32'hbf641549, 32'h00000000} /* (10, 12, 9) {real, imag} */,
  {32'hbf621943, 32'h00000000} /* (10, 12, 8) {real, imag} */,
  {32'hbf9dad9b, 32'h00000000} /* (10, 12, 7) {real, imag} */,
  {32'hbf9b7f23, 32'h00000000} /* (10, 12, 6) {real, imag} */,
  {32'hbf840c93, 32'h00000000} /* (10, 12, 5) {real, imag} */,
  {32'hbf6feaea, 32'h00000000} /* (10, 12, 4) {real, imag} */,
  {32'hbf1e1f3a, 32'h00000000} /* (10, 12, 3) {real, imag} */,
  {32'hbec1176f, 32'h00000000} /* (10, 12, 2) {real, imag} */,
  {32'hbf4614e3, 32'h00000000} /* (10, 12, 1) {real, imag} */,
  {32'hbf2a41c9, 32'h00000000} /* (10, 12, 0) {real, imag} */,
  {32'hbec37ccc, 32'h00000000} /* (10, 11, 31) {real, imag} */,
  {32'hbe886725, 32'h00000000} /* (10, 11, 30) {real, imag} */,
  {32'hbe501c58, 32'h00000000} /* (10, 11, 29) {real, imag} */,
  {32'hbf29c14d, 32'h00000000} /* (10, 11, 28) {real, imag} */,
  {32'hbf4e7c48, 32'h00000000} /* (10, 11, 27) {real, imag} */,
  {32'hbf2b753d, 32'h00000000} /* (10, 11, 26) {real, imag} */,
  {32'hbefd2576, 32'h00000000} /* (10, 11, 25) {real, imag} */,
  {32'hbf2f4cdf, 32'h00000000} /* (10, 11, 24) {real, imag} */,
  {32'hbf0ff653, 32'h00000000} /* (10, 11, 23) {real, imag} */,
  {32'hbef466c1, 32'h00000000} /* (10, 11, 22) {real, imag} */,
  {32'hbed3448c, 32'h00000000} /* (10, 11, 21) {real, imag} */,
  {32'h3ebeeb46, 32'h00000000} /* (10, 11, 20) {real, imag} */,
  {32'h3f85ce90, 32'h00000000} /* (10, 11, 19) {real, imag} */,
  {32'h3f83e9e5, 32'h00000000} /* (10, 11, 18) {real, imag} */,
  {32'h3f624b1a, 32'h00000000} /* (10, 11, 17) {real, imag} */,
  {32'h3fb80b59, 32'h00000000} /* (10, 11, 16) {real, imag} */,
  {32'h3fa0bad2, 32'h00000000} /* (10, 11, 15) {real, imag} */,
  {32'h3f6ef105, 32'h00000000} /* (10, 11, 14) {real, imag} */,
  {32'h3f3c3049, 32'h00000000} /* (10, 11, 13) {real, imag} */,
  {32'h3f397098, 32'h00000000} /* (10, 11, 12) {real, imag} */,
  {32'h3f0ced05, 32'h00000000} /* (10, 11, 11) {real, imag} */,
  {32'hbe2b35da, 32'h00000000} /* (10, 11, 10) {real, imag} */,
  {32'hbd98d9ff, 32'h00000000} /* (10, 11, 9) {real, imag} */,
  {32'hbe88fae4, 32'h00000000} /* (10, 11, 8) {real, imag} */,
  {32'hbecc85e1, 32'h00000000} /* (10, 11, 7) {real, imag} */,
  {32'hbeee8699, 32'h00000000} /* (10, 11, 6) {real, imag} */,
  {32'hbdf411b4, 32'h00000000} /* (10, 11, 5) {real, imag} */,
  {32'hbee726d6, 32'h00000000} /* (10, 11, 4) {real, imag} */,
  {32'hbf2cf898, 32'h00000000} /* (10, 11, 3) {real, imag} */,
  {32'hbf4eb987, 32'h00000000} /* (10, 11, 2) {real, imag} */,
  {32'hbefea56d, 32'h00000000} /* (10, 11, 1) {real, imag} */,
  {32'hbe2bacf2, 32'h00000000} /* (10, 11, 0) {real, imag} */,
  {32'h3e6ddcaf, 32'h00000000} /* (10, 10, 31) {real, imag} */,
  {32'h3f2f40d5, 32'h00000000} /* (10, 10, 30) {real, imag} */,
  {32'h3f923d60, 32'h00000000} /* (10, 10, 29) {real, imag} */,
  {32'h3eb5bc35, 32'h00000000} /* (10, 10, 28) {real, imag} */,
  {32'h3dabbeb0, 32'h00000000} /* (10, 10, 27) {real, imag} */,
  {32'h3edbe496, 32'h00000000} /* (10, 10, 26) {real, imag} */,
  {32'h3ef5c8f9, 32'h00000000} /* (10, 10, 25) {real, imag} */,
  {32'h3f02a97d, 32'h00000000} /* (10, 10, 24) {real, imag} */,
  {32'h3f32b79a, 32'h00000000} /* (10, 10, 23) {real, imag} */,
  {32'h3f2dbdca, 32'h00000000} /* (10, 10, 22) {real, imag} */,
  {32'h3f2a6b33, 32'h00000000} /* (10, 10, 21) {real, imag} */,
  {32'h3e4d49ec, 32'h00000000} /* (10, 10, 20) {real, imag} */,
  {32'hbf1b10a1, 32'h00000000} /* (10, 10, 19) {real, imag} */,
  {32'hbeb893b2, 32'h00000000} /* (10, 10, 18) {real, imag} */,
  {32'h3d20f4ca, 32'h00000000} /* (10, 10, 17) {real, imag} */,
  {32'hbe968f82, 32'h00000000} /* (10, 10, 16) {real, imag} */,
  {32'hbe30185c, 32'h00000000} /* (10, 10, 15) {real, imag} */,
  {32'hbdaec83f, 32'h00000000} /* (10, 10, 14) {real, imag} */,
  {32'hbe1fdede, 32'h00000000} /* (10, 10, 13) {real, imag} */,
  {32'hbf0625f7, 32'h00000000} /* (10, 10, 12) {real, imag} */,
  {32'hbe8eb32f, 32'h00000000} /* (10, 10, 11) {real, imag} */,
  {32'hbce739c8, 32'h00000000} /* (10, 10, 10) {real, imag} */,
  {32'h3eec05e7, 32'h00000000} /* (10, 10, 9) {real, imag} */,
  {32'h3ef47acf, 32'h00000000} /* (10, 10, 8) {real, imag} */,
  {32'h3faab8ab, 32'h00000000} /* (10, 10, 7) {real, imag} */,
  {32'h3fa9d456, 32'h00000000} /* (10, 10, 6) {real, imag} */,
  {32'h3fae1501, 32'h00000000} /* (10, 10, 5) {real, imag} */,
  {32'h3f895655, 32'h00000000} /* (10, 10, 4) {real, imag} */,
  {32'h3e4aee03, 32'h00000000} /* (10, 10, 3) {real, imag} */,
  {32'hbe6253e6, 32'h00000000} /* (10, 10, 2) {real, imag} */,
  {32'h3e7d32ca, 32'h00000000} /* (10, 10, 1) {real, imag} */,
  {32'h3eaa94dc, 32'h00000000} /* (10, 10, 0) {real, imag} */,
  {32'h3ee8fd83, 32'h00000000} /* (10, 9, 31) {real, imag} */,
  {32'h3f1a8969, 32'h00000000} /* (10, 9, 30) {real, imag} */,
  {32'h3faf04db, 32'h00000000} /* (10, 9, 29) {real, imag} */,
  {32'h3fd4fc62, 32'h00000000} /* (10, 9, 28) {real, imag} */,
  {32'h3fa5688b, 32'h00000000} /* (10, 9, 27) {real, imag} */,
  {32'h3f626e07, 32'h00000000} /* (10, 9, 26) {real, imag} */,
  {32'h3f4e9f43, 32'h00000000} /* (10, 9, 25) {real, imag} */,
  {32'h3f6626e6, 32'h00000000} /* (10, 9, 24) {real, imag} */,
  {32'h3f7b006f, 32'h00000000} /* (10, 9, 23) {real, imag} */,
  {32'h3f676397, 32'h00000000} /* (10, 9, 22) {real, imag} */,
  {32'h3f011bd6, 32'h00000000} /* (10, 9, 21) {real, imag} */,
  {32'hbd1713c2, 32'h00000000} /* (10, 9, 20) {real, imag} */,
  {32'hbf873317, 32'h00000000} /* (10, 9, 19) {real, imag} */,
  {32'hbf8bf340, 32'h00000000} /* (10, 9, 18) {real, imag} */,
  {32'hbf2f87e6, 32'h00000000} /* (10, 9, 17) {real, imag} */,
  {32'hbfac9451, 32'h00000000} /* (10, 9, 16) {real, imag} */,
  {32'hbf8cc004, 32'h00000000} /* (10, 9, 15) {real, imag} */,
  {32'hbef51f24, 32'h00000000} /* (10, 9, 14) {real, imag} */,
  {32'hbea96f4c, 32'h00000000} /* (10, 9, 13) {real, imag} */,
  {32'hbf56a887, 32'h00000000} /* (10, 9, 12) {real, imag} */,
  {32'hbf73eed0, 32'h00000000} /* (10, 9, 11) {real, imag} */,
  {32'h3de51e84, 32'h00000000} /* (10, 9, 10) {real, imag} */,
  {32'h3f853a72, 32'h00000000} /* (10, 9, 9) {real, imag} */,
  {32'h3f8ec3e3, 32'h00000000} /* (10, 9, 8) {real, imag} */,
  {32'h3fc0cd3f, 32'h00000000} /* (10, 9, 7) {real, imag} */,
  {32'h3f950be2, 32'h00000000} /* (10, 9, 6) {real, imag} */,
  {32'h3f6c5813, 32'h00000000} /* (10, 9, 5) {real, imag} */,
  {32'h3f8ac394, 32'h00000000} /* (10, 9, 4) {real, imag} */,
  {32'h3fa3b6b8, 32'h00000000} /* (10, 9, 3) {real, imag} */,
  {32'h3f07e19a, 32'h00000000} /* (10, 9, 2) {real, imag} */,
  {32'h3ef7f003, 32'h00000000} /* (10, 9, 1) {real, imag} */,
  {32'h3ec44bb4, 32'h00000000} /* (10, 9, 0) {real, imag} */,
  {32'h3d8aff55, 32'h00000000} /* (10, 8, 31) {real, imag} */,
  {32'h3e999bad, 32'h00000000} /* (10, 8, 30) {real, imag} */,
  {32'h3f95eba3, 32'h00000000} /* (10, 8, 29) {real, imag} */,
  {32'h3f8b75c6, 32'h00000000} /* (10, 8, 28) {real, imag} */,
  {32'h3fd9fa8f, 32'h00000000} /* (10, 8, 27) {real, imag} */,
  {32'h3fa80f76, 32'h00000000} /* (10, 8, 26) {real, imag} */,
  {32'h3f41a64d, 32'h00000000} /* (10, 8, 25) {real, imag} */,
  {32'h3f372ed4, 32'h00000000} /* (10, 8, 24) {real, imag} */,
  {32'h3f84b31d, 32'h00000000} /* (10, 8, 23) {real, imag} */,
  {32'h3f5ba4aa, 32'h00000000} /* (10, 8, 22) {real, imag} */,
  {32'h3e40b6ac, 32'h00000000} /* (10, 8, 21) {real, imag} */,
  {32'hbe5e0474, 32'h00000000} /* (10, 8, 20) {real, imag} */,
  {32'hbf0667ea, 32'h00000000} /* (10, 8, 19) {real, imag} */,
  {32'hbf7a7d57, 32'h00000000} /* (10, 8, 18) {real, imag} */,
  {32'hbf5d7af2, 32'h00000000} /* (10, 8, 17) {real, imag} */,
  {32'hbf66f4a0, 32'h00000000} /* (10, 8, 16) {real, imag} */,
  {32'hbf54638e, 32'h00000000} /* (10, 8, 15) {real, imag} */,
  {32'hbf2996e7, 32'h00000000} /* (10, 8, 14) {real, imag} */,
  {32'hbeeb0716, 32'h00000000} /* (10, 8, 13) {real, imag} */,
  {32'hbf523612, 32'h00000000} /* (10, 8, 12) {real, imag} */,
  {32'hbf9f514a, 32'h00000000} /* (10, 8, 11) {real, imag} */,
  {32'hbb6d0848, 32'h00000000} /* (10, 8, 10) {real, imag} */,
  {32'h3f91849b, 32'h00000000} /* (10, 8, 9) {real, imag} */,
  {32'h3fa73811, 32'h00000000} /* (10, 8, 8) {real, imag} */,
  {32'h3fd3cd16, 32'h00000000} /* (10, 8, 7) {real, imag} */,
  {32'h3f9f798c, 32'h00000000} /* (10, 8, 6) {real, imag} */,
  {32'h3f4a8efd, 32'h00000000} /* (10, 8, 5) {real, imag} */,
  {32'h3f851fb4, 32'h00000000} /* (10, 8, 4) {real, imag} */,
  {32'h3f94047e, 32'h00000000} /* (10, 8, 3) {real, imag} */,
  {32'h3f86c2d1, 32'h00000000} /* (10, 8, 2) {real, imag} */,
  {32'h3f82f7a0, 32'h00000000} /* (10, 8, 1) {real, imag} */,
  {32'h3ef771fd, 32'h00000000} /* (10, 8, 0) {real, imag} */,
  {32'h3ef6f410, 32'h00000000} /* (10, 7, 31) {real, imag} */,
  {32'h3f1068a9, 32'h00000000} /* (10, 7, 30) {real, imag} */,
  {32'h3fba5044, 32'h00000000} /* (10, 7, 29) {real, imag} */,
  {32'h3f7fcb30, 32'h00000000} /* (10, 7, 28) {real, imag} */,
  {32'h3f987b1a, 32'h00000000} /* (10, 7, 27) {real, imag} */,
  {32'h3f88ed9c, 32'h00000000} /* (10, 7, 26) {real, imag} */,
  {32'h3f1d3765, 32'h00000000} /* (10, 7, 25) {real, imag} */,
  {32'h3f4b8393, 32'h00000000} /* (10, 7, 24) {real, imag} */,
  {32'h3f7c8f7b, 32'h00000000} /* (10, 7, 23) {real, imag} */,
  {32'h3f91a03d, 32'h00000000} /* (10, 7, 22) {real, imag} */,
  {32'h3f25efa3, 32'h00000000} /* (10, 7, 21) {real, imag} */,
  {32'hbd4b9261, 32'h00000000} /* (10, 7, 20) {real, imag} */,
  {32'hbe367cb5, 32'h00000000} /* (10, 7, 19) {real, imag} */,
  {32'hbf618260, 32'h00000000} /* (10, 7, 18) {real, imag} */,
  {32'hbf4a5a8e, 32'h00000000} /* (10, 7, 17) {real, imag} */,
  {32'hbf6a3b05, 32'h00000000} /* (10, 7, 16) {real, imag} */,
  {32'hbf56a364, 32'h00000000} /* (10, 7, 15) {real, imag} */,
  {32'hbf51fe7c, 32'h00000000} /* (10, 7, 14) {real, imag} */,
  {32'hbf1f852d, 32'h00000000} /* (10, 7, 13) {real, imag} */,
  {32'hbf8c26c8, 32'h00000000} /* (10, 7, 12) {real, imag} */,
  {32'hbf898f3e, 32'h00000000} /* (10, 7, 11) {real, imag} */,
  {32'h3cdb52e5, 32'h00000000} /* (10, 7, 10) {real, imag} */,
  {32'h3f0c7595, 32'h00000000} /* (10, 7, 9) {real, imag} */,
  {32'h3f8efd2a, 32'h00000000} /* (10, 7, 8) {real, imag} */,
  {32'h3ff524d7, 32'h00000000} /* (10, 7, 7) {real, imag} */,
  {32'h3fb5fe8f, 32'h00000000} /* (10, 7, 6) {real, imag} */,
  {32'h3f6bac4f, 32'h00000000} /* (10, 7, 5) {real, imag} */,
  {32'h3fafd79c, 32'h00000000} /* (10, 7, 4) {real, imag} */,
  {32'h3fc6edba, 32'h00000000} /* (10, 7, 3) {real, imag} */,
  {32'h3f7ceb68, 32'h00000000} /* (10, 7, 2) {real, imag} */,
  {32'h3f8f17e5, 32'h00000000} /* (10, 7, 1) {real, imag} */,
  {32'h3f011a62, 32'h00000000} /* (10, 7, 0) {real, imag} */,
  {32'h3f37d7be, 32'h00000000} /* (10, 6, 31) {real, imag} */,
  {32'h3ee75c3d, 32'h00000000} /* (10, 6, 30) {real, imag} */,
  {32'h3f448293, 32'h00000000} /* (10, 6, 29) {real, imag} */,
  {32'h3f82add2, 32'h00000000} /* (10, 6, 28) {real, imag} */,
  {32'h3f899b77, 32'h00000000} /* (10, 6, 27) {real, imag} */,
  {32'h3f863e4b, 32'h00000000} /* (10, 6, 26) {real, imag} */,
  {32'h3f456559, 32'h00000000} /* (10, 6, 25) {real, imag} */,
  {32'h3f7e4a89, 32'h00000000} /* (10, 6, 24) {real, imag} */,
  {32'h3f811ff3, 32'h00000000} /* (10, 6, 23) {real, imag} */,
  {32'h3f6ed27e, 32'h00000000} /* (10, 6, 22) {real, imag} */,
  {32'h3f862563, 32'h00000000} /* (10, 6, 21) {real, imag} */,
  {32'h3e4bb555, 32'h00000000} /* (10, 6, 20) {real, imag} */,
  {32'hbd348ea1, 32'h00000000} /* (10, 6, 19) {real, imag} */,
  {32'hbf4644a8, 32'h00000000} /* (10, 6, 18) {real, imag} */,
  {32'hbf11f7cc, 32'h00000000} /* (10, 6, 17) {real, imag} */,
  {32'hbf61c169, 32'h00000000} /* (10, 6, 16) {real, imag} */,
  {32'hbf4dbc05, 32'h00000000} /* (10, 6, 15) {real, imag} */,
  {32'hbf6d1721, 32'h00000000} /* (10, 6, 14) {real, imag} */,
  {32'hbf415155, 32'h00000000} /* (10, 6, 13) {real, imag} */,
  {32'hbf8c5514, 32'h00000000} /* (10, 6, 12) {real, imag} */,
  {32'hbf4cb8c5, 32'h00000000} /* (10, 6, 11) {real, imag} */,
  {32'h3eb66ebb, 32'h00000000} /* (10, 6, 10) {real, imag} */,
  {32'h3e66e139, 32'h00000000} /* (10, 6, 9) {real, imag} */,
  {32'h3ee95944, 32'h00000000} /* (10, 6, 8) {real, imag} */,
  {32'h3f8663ad, 32'h00000000} /* (10, 6, 7) {real, imag} */,
  {32'h3f757ffd, 32'h00000000} /* (10, 6, 6) {real, imag} */,
  {32'h3f905245, 32'h00000000} /* (10, 6, 5) {real, imag} */,
  {32'h3fa67745, 32'h00000000} /* (10, 6, 4) {real, imag} */,
  {32'h3fb804b7, 32'h00000000} /* (10, 6, 3) {real, imag} */,
  {32'h3f804911, 32'h00000000} /* (10, 6, 2) {real, imag} */,
  {32'h3fa9ad5d, 32'h00000000} /* (10, 6, 1) {real, imag} */,
  {32'h3f595187, 32'h00000000} /* (10, 6, 0) {real, imag} */,
  {32'h3e327209, 32'h00000000} /* (10, 5, 31) {real, imag} */,
  {32'h3ed70ded, 32'h00000000} /* (10, 5, 30) {real, imag} */,
  {32'h3f179ca5, 32'h00000000} /* (10, 5, 29) {real, imag} */,
  {32'h3f5f5ee0, 32'h00000000} /* (10, 5, 28) {real, imag} */,
  {32'h3fc6e60b, 32'h00000000} /* (10, 5, 27) {real, imag} */,
  {32'h3fc46421, 32'h00000000} /* (10, 5, 26) {real, imag} */,
  {32'h3f8f4b02, 32'h00000000} /* (10, 5, 25) {real, imag} */,
  {32'h3f0a4aa2, 32'h00000000} /* (10, 5, 24) {real, imag} */,
  {32'h3f835760, 32'h00000000} /* (10, 5, 23) {real, imag} */,
  {32'h3f96808a, 32'h00000000} /* (10, 5, 22) {real, imag} */,
  {32'h3fa4ca89, 32'h00000000} /* (10, 5, 21) {real, imag} */,
  {32'h3f7d0296, 32'h00000000} /* (10, 5, 20) {real, imag} */,
  {32'h3f1d3b66, 32'h00000000} /* (10, 5, 19) {real, imag} */,
  {32'h3e6c7366, 32'h00000000} /* (10, 5, 18) {real, imag} */,
  {32'h3f29ee9f, 32'h00000000} /* (10, 5, 17) {real, imag} */,
  {32'h3df6658c, 32'h00000000} /* (10, 5, 16) {real, imag} */,
  {32'hbf2b1863, 32'h00000000} /* (10, 5, 15) {real, imag} */,
  {32'hbf2670d6, 32'h00000000} /* (10, 5, 14) {real, imag} */,
  {32'hbf058b1e, 32'h00000000} /* (10, 5, 13) {real, imag} */,
  {32'hbfa449ac, 32'h00000000} /* (10, 5, 12) {real, imag} */,
  {32'hbfb71799, 32'h00000000} /* (10, 5, 11) {real, imag} */,
  {32'h3dac49df, 32'h00000000} /* (10, 5, 10) {real, imag} */,
  {32'h3deda81b, 32'h00000000} /* (10, 5, 9) {real, imag} */,
  {32'hbbea4820, 32'h00000000} /* (10, 5, 8) {real, imag} */,
  {32'hbbd91006, 32'h00000000} /* (10, 5, 7) {real, imag} */,
  {32'h3d4606ae, 32'h00000000} /* (10, 5, 6) {real, imag} */,
  {32'h3f23a313, 32'h00000000} /* (10, 5, 5) {real, imag} */,
  {32'h3f0ef43f, 32'h00000000} /* (10, 5, 4) {real, imag} */,
  {32'h3f65594c, 32'h00000000} /* (10, 5, 3) {real, imag} */,
  {32'h3fa39d1e, 32'h00000000} /* (10, 5, 2) {real, imag} */,
  {32'h3fb59424, 32'h00000000} /* (10, 5, 1) {real, imag} */,
  {32'h3ef2fadc, 32'h00000000} /* (10, 5, 0) {real, imag} */,
  {32'h3e97605b, 32'h00000000} /* (10, 4, 31) {real, imag} */,
  {32'h3f2bd4b4, 32'h00000000} /* (10, 4, 30) {real, imag} */,
  {32'h3f5091c5, 32'h00000000} /* (10, 4, 29) {real, imag} */,
  {32'h3f85cbbf, 32'h00000000} /* (10, 4, 28) {real, imag} */,
  {32'h3fad9d7f, 32'h00000000} /* (10, 4, 27) {real, imag} */,
  {32'h3f9f9734, 32'h00000000} /* (10, 4, 26) {real, imag} */,
  {32'h3f7f8049, 32'h00000000} /* (10, 4, 25) {real, imag} */,
  {32'h3f0eb6e3, 32'h00000000} /* (10, 4, 24) {real, imag} */,
  {32'h3f3b1689, 32'h00000000} /* (10, 4, 23) {real, imag} */,
  {32'h3fa110b9, 32'h00000000} /* (10, 4, 22) {real, imag} */,
  {32'h3fabba5f, 32'h00000000} /* (10, 4, 21) {real, imag} */,
  {32'h3f92ef3a, 32'h00000000} /* (10, 4, 20) {real, imag} */,
  {32'h3f2891bd, 32'h00000000} /* (10, 4, 19) {real, imag} */,
  {32'h3f324104, 32'h00000000} /* (10, 4, 18) {real, imag} */,
  {32'h3fafd91a, 32'h00000000} /* (10, 4, 17) {real, imag} */,
  {32'h3eecf61d, 32'h00000000} /* (10, 4, 16) {real, imag} */,
  {32'hbf73e8e5, 32'h00000000} /* (10, 4, 15) {real, imag} */,
  {32'hbe40548b, 32'h00000000} /* (10, 4, 14) {real, imag} */,
  {32'hbea72667, 32'h00000000} /* (10, 4, 13) {real, imag} */,
  {32'hbf737c5d, 32'h00000000} /* (10, 4, 12) {real, imag} */,
  {32'hbf99a84c, 32'h00000000} /* (10, 4, 11) {real, imag} */,
  {32'hbe51de5c, 32'h00000000} /* (10, 4, 10) {real, imag} */,
  {32'hbdf0402c, 32'h00000000} /* (10, 4, 9) {real, imag} */,
  {32'hbf3bde9d, 32'h00000000} /* (10, 4, 8) {real, imag} */,
  {32'hbf15c53d, 32'h00000000} /* (10, 4, 7) {real, imag} */,
  {32'hbea7f001, 32'h00000000} /* (10, 4, 6) {real, imag} */,
  {32'h3eb294ab, 32'h00000000} /* (10, 4, 5) {real, imag} */,
  {32'h3f1c45ea, 32'h00000000} /* (10, 4, 4) {real, imag} */,
  {32'h3f465cd6, 32'h00000000} /* (10, 4, 3) {real, imag} */,
  {32'h3f95c27b, 32'h00000000} /* (10, 4, 2) {real, imag} */,
  {32'h3fa43add, 32'h00000000} /* (10, 4, 1) {real, imag} */,
  {32'h3f226669, 32'h00000000} /* (10, 4, 0) {real, imag} */,
  {32'h3e6fea83, 32'h00000000} /* (10, 3, 31) {real, imag} */,
  {32'h3f38aa2d, 32'h00000000} /* (10, 3, 30) {real, imag} */,
  {32'h3f8559ac, 32'h00000000} /* (10, 3, 29) {real, imag} */,
  {32'h3fabcef2, 32'h00000000} /* (10, 3, 28) {real, imag} */,
  {32'h3f2e7c66, 32'h00000000} /* (10, 3, 27) {real, imag} */,
  {32'h3f026825, 32'h00000000} /* (10, 3, 26) {real, imag} */,
  {32'h3f5c76f8, 32'h00000000} /* (10, 3, 25) {real, imag} */,
  {32'h3fb38a64, 32'h00000000} /* (10, 3, 24) {real, imag} */,
  {32'h3f62e0d6, 32'h00000000} /* (10, 3, 23) {real, imag} */,
  {32'h3f545689, 32'h00000000} /* (10, 3, 22) {real, imag} */,
  {32'h3fa4f40b, 32'h00000000} /* (10, 3, 21) {real, imag} */,
  {32'h3f9049d7, 32'h00000000} /* (10, 3, 20) {real, imag} */,
  {32'h3f59f90c, 32'h00000000} /* (10, 3, 19) {real, imag} */,
  {32'h3f2104ea, 32'h00000000} /* (10, 3, 18) {real, imag} */,
  {32'h3f703ceb, 32'h00000000} /* (10, 3, 17) {real, imag} */,
  {32'h3e4c02be, 32'h00000000} /* (10, 3, 16) {real, imag} */,
  {32'hbf8b9af4, 32'h00000000} /* (10, 3, 15) {real, imag} */,
  {32'hbf4254bc, 32'h00000000} /* (10, 3, 14) {real, imag} */,
  {32'hbf0ef750, 32'h00000000} /* (10, 3, 13) {real, imag} */,
  {32'hbf17e82c, 32'h00000000} /* (10, 3, 12) {real, imag} */,
  {32'hbf9862a2, 32'h00000000} /* (10, 3, 11) {real, imag} */,
  {32'hbf33b578, 32'h00000000} /* (10, 3, 10) {real, imag} */,
  {32'hbf162dcb, 32'h00000000} /* (10, 3, 9) {real, imag} */,
  {32'hbfb16bf2, 32'h00000000} /* (10, 3, 8) {real, imag} */,
  {32'hbf9fff01, 32'h00000000} /* (10, 3, 7) {real, imag} */,
  {32'hbf35e612, 32'h00000000} /* (10, 3, 6) {real, imag} */,
  {32'h3cd89c54, 32'h00000000} /* (10, 3, 5) {real, imag} */,
  {32'h3f69dcfe, 32'h00000000} /* (10, 3, 4) {real, imag} */,
  {32'h3f6d387b, 32'h00000000} /* (10, 3, 3) {real, imag} */,
  {32'h3fac0c20, 32'h00000000} /* (10, 3, 2) {real, imag} */,
  {32'h3fa49884, 32'h00000000} /* (10, 3, 1) {real, imag} */,
  {32'h3f42def1, 32'h00000000} /* (10, 3, 0) {real, imag} */,
  {32'h3e093711, 32'h00000000} /* (10, 2, 31) {real, imag} */,
  {32'h3efa26f7, 32'h00000000} /* (10, 2, 30) {real, imag} */,
  {32'h3f6adbcd, 32'h00000000} /* (10, 2, 29) {real, imag} */,
  {32'h3f91f46e, 32'h00000000} /* (10, 2, 28) {real, imag} */,
  {32'h3f306bc1, 32'h00000000} /* (10, 2, 27) {real, imag} */,
  {32'h3ec2018b, 32'h00000000} /* (10, 2, 26) {real, imag} */,
  {32'h3f5548d7, 32'h00000000} /* (10, 2, 25) {real, imag} */,
  {32'h3f889fb3, 32'h00000000} /* (10, 2, 24) {real, imag} */,
  {32'h3f665563, 32'h00000000} /* (10, 2, 23) {real, imag} */,
  {32'h3f07f3b5, 32'h00000000} /* (10, 2, 22) {real, imag} */,
  {32'h3f3ab804, 32'h00000000} /* (10, 2, 21) {real, imag} */,
  {32'h3f815ab2, 32'h00000000} /* (10, 2, 20) {real, imag} */,
  {32'h3fb2355d, 32'h00000000} /* (10, 2, 19) {real, imag} */,
  {32'h3f8958b7, 32'h00000000} /* (10, 2, 18) {real, imag} */,
  {32'h3f8b3a99, 32'h00000000} /* (10, 2, 17) {real, imag} */,
  {32'h3e45d8c4, 32'h00000000} /* (10, 2, 16) {real, imag} */,
  {32'hbf93c508, 32'h00000000} /* (10, 2, 15) {real, imag} */,
  {32'hbfb6eccc, 32'h00000000} /* (10, 2, 14) {real, imag} */,
  {32'hbf69e642, 32'h00000000} /* (10, 2, 13) {real, imag} */,
  {32'hbf63de35, 32'h00000000} /* (10, 2, 12) {real, imag} */,
  {32'hbf99b9db, 32'h00000000} /* (10, 2, 11) {real, imag} */,
  {32'hbf94478e, 32'h00000000} /* (10, 2, 10) {real, imag} */,
  {32'hbf5d112e, 32'h00000000} /* (10, 2, 9) {real, imag} */,
  {32'hbfa7f903, 32'h00000000} /* (10, 2, 8) {real, imag} */,
  {32'hbfad7c96, 32'h00000000} /* (10, 2, 7) {real, imag} */,
  {32'hbf66c1ca, 32'h00000000} /* (10, 2, 6) {real, imag} */,
  {32'hbd955540, 32'h00000000} /* (10, 2, 5) {real, imag} */,
  {32'h3f20afee, 32'h00000000} /* (10, 2, 4) {real, imag} */,
  {32'h3f547186, 32'h00000000} /* (10, 2, 3) {real, imag} */,
  {32'h3f7bb036, 32'h00000000} /* (10, 2, 2) {real, imag} */,
  {32'h3f42a4d8, 32'h00000000} /* (10, 2, 1) {real, imag} */,
  {32'h3ec03f7f, 32'h00000000} /* (10, 2, 0) {real, imag} */,
  {32'h3e24b87f, 32'h00000000} /* (10, 1, 31) {real, imag} */,
  {32'h3f18fc15, 32'h00000000} /* (10, 1, 30) {real, imag} */,
  {32'h3f9f6573, 32'h00000000} /* (10, 1, 29) {real, imag} */,
  {32'h3fc396c6, 32'h00000000} /* (10, 1, 28) {real, imag} */,
  {32'h3faec4a8, 32'h00000000} /* (10, 1, 27) {real, imag} */,
  {32'h3f3f11ee, 32'h00000000} /* (10, 1, 26) {real, imag} */,
  {32'h3f3553c9, 32'h00000000} /* (10, 1, 25) {real, imag} */,
  {32'h3f6d90c1, 32'h00000000} /* (10, 1, 24) {real, imag} */,
  {32'h3f199666, 32'h00000000} /* (10, 1, 23) {real, imag} */,
  {32'h3ea9f69a, 32'h00000000} /* (10, 1, 22) {real, imag} */,
  {32'h3efde3d1, 32'h00000000} /* (10, 1, 21) {real, imag} */,
  {32'h3f396ad3, 32'h00000000} /* (10, 1, 20) {real, imag} */,
  {32'h3f931454, 32'h00000000} /* (10, 1, 19) {real, imag} */,
  {32'h3fa7d9bf, 32'h00000000} /* (10, 1, 18) {real, imag} */,
  {32'h3f7e7e37, 32'h00000000} /* (10, 1, 17) {real, imag} */,
  {32'h3e2e53fc, 32'h00000000} /* (10, 1, 16) {real, imag} */,
  {32'hbf59fa78, 32'h00000000} /* (10, 1, 15) {real, imag} */,
  {32'hbf9e41fe, 32'h00000000} /* (10, 1, 14) {real, imag} */,
  {32'hbfd7b37c, 32'h00000000} /* (10, 1, 13) {real, imag} */,
  {32'hbfa66fec, 32'h00000000} /* (10, 1, 12) {real, imag} */,
  {32'hbf800308, 32'h00000000} /* (10, 1, 11) {real, imag} */,
  {32'hbf8b9123, 32'h00000000} /* (10, 1, 10) {real, imag} */,
  {32'hbf07f6d4, 32'h00000000} /* (10, 1, 9) {real, imag} */,
  {32'hbf114f28, 32'h00000000} /* (10, 1, 8) {real, imag} */,
  {32'hbf74c788, 32'h00000000} /* (10, 1, 7) {real, imag} */,
  {32'hbf4d80a9, 32'h00000000} /* (10, 1, 6) {real, imag} */,
  {32'hbcce0570, 32'h00000000} /* (10, 1, 5) {real, imag} */,
  {32'h3ef0a8b7, 32'h00000000} /* (10, 1, 4) {real, imag} */,
  {32'h3f25186c, 32'h00000000} /* (10, 1, 3) {real, imag} */,
  {32'h3f10de44, 32'h00000000} /* (10, 1, 2) {real, imag} */,
  {32'h3f189569, 32'h00000000} /* (10, 1, 1) {real, imag} */,
  {32'h3e462c43, 32'h00000000} /* (10, 1, 0) {real, imag} */,
  {32'h3e48df33, 32'h00000000} /* (10, 0, 31) {real, imag} */,
  {32'h3edcf8a8, 32'h00000000} /* (10, 0, 30) {real, imag} */,
  {32'h3f2cfb3c, 32'h00000000} /* (10, 0, 29) {real, imag} */,
  {32'h3f837d9f, 32'h00000000} /* (10, 0, 28) {real, imag} */,
  {32'h3f91cc24, 32'h00000000} /* (10, 0, 27) {real, imag} */,
  {32'h3ee23def, 32'h00000000} /* (10, 0, 26) {real, imag} */,
  {32'h3e885f7c, 32'h00000000} /* (10, 0, 25) {real, imag} */,
  {32'h3ef4c996, 32'h00000000} /* (10, 0, 24) {real, imag} */,
  {32'h3e9f7cda, 32'h00000000} /* (10, 0, 23) {real, imag} */,
  {32'h3e88472e, 32'h00000000} /* (10, 0, 22) {real, imag} */,
  {32'h3e68fb41, 32'h00000000} /* (10, 0, 21) {real, imag} */,
  {32'h3cb59c74, 32'h00000000} /* (10, 0, 20) {real, imag} */,
  {32'h3e8d3e78, 32'h00000000} /* (10, 0, 19) {real, imag} */,
  {32'h3f350893, 32'h00000000} /* (10, 0, 18) {real, imag} */,
  {32'h3eff9789, 32'h00000000} /* (10, 0, 17) {real, imag} */,
  {32'h3dac225e, 32'h00000000} /* (10, 0, 16) {real, imag} */,
  {32'hbe3e2f51, 32'h00000000} /* (10, 0, 15) {real, imag} */,
  {32'hbecec09a, 32'h00000000} /* (10, 0, 14) {real, imag} */,
  {32'hbf70708d, 32'h00000000} /* (10, 0, 13) {real, imag} */,
  {32'hbf0c47a5, 32'h00000000} /* (10, 0, 12) {real, imag} */,
  {32'hbecd8d18, 32'h00000000} /* (10, 0, 11) {real, imag} */,
  {32'hbe7d8bde, 32'h00000000} /* (10, 0, 10) {real, imag} */,
  {32'hbe413860, 32'h00000000} /* (10, 0, 9) {real, imag} */,
  {32'hbea656c7, 32'h00000000} /* (10, 0, 8) {real, imag} */,
  {32'hbf141f60, 32'h00000000} /* (10, 0, 7) {real, imag} */,
  {32'hbed9c911, 32'h00000000} /* (10, 0, 6) {real, imag} */,
  {32'h3c4ef4d4, 32'h00000000} /* (10, 0, 5) {real, imag} */,
  {32'h3eab0acc, 32'h00000000} /* (10, 0, 4) {real, imag} */,
  {32'h3f07fe44, 32'h00000000} /* (10, 0, 3) {real, imag} */,
  {32'h3ecbd57b, 32'h00000000} /* (10, 0, 2) {real, imag} */,
  {32'h3ee4aef4, 32'h00000000} /* (10, 0, 1) {real, imag} */,
  {32'h3e5fe19e, 32'h00000000} /* (10, 0, 0) {real, imag} */,
  {32'h3ae8afcb, 32'h00000000} /* (9, 31, 31) {real, imag} */,
  {32'h3e15abbf, 32'h00000000} /* (9, 31, 30) {real, imag} */,
  {32'h3f144f36, 32'h00000000} /* (9, 31, 29) {real, imag} */,
  {32'h3ea4fd88, 32'h00000000} /* (9, 31, 28) {real, imag} */,
  {32'h3ee9319c, 32'h00000000} /* (9, 31, 27) {real, imag} */,
  {32'h3f01dd89, 32'h00000000} /* (9, 31, 26) {real, imag} */,
  {32'h3f112784, 32'h00000000} /* (9, 31, 25) {real, imag} */,
  {32'h3f673b52, 32'h00000000} /* (9, 31, 24) {real, imag} */,
  {32'h3f36fb42, 32'h00000000} /* (9, 31, 23) {real, imag} */,
  {32'h3f6db93e, 32'h00000000} /* (9, 31, 22) {real, imag} */,
  {32'h3f247707, 32'h00000000} /* (9, 31, 21) {real, imag} */,
  {32'hbe17cb9e, 32'h00000000} /* (9, 31, 20) {real, imag} */,
  {32'hbe24423b, 32'h00000000} /* (9, 31, 19) {real, imag} */,
  {32'hbd0cccef, 32'h00000000} /* (9, 31, 18) {real, imag} */,
  {32'hbddfe0d4, 32'h00000000} /* (9, 31, 17) {real, imag} */,
  {32'hbf01eff5, 32'h00000000} /* (9, 31, 16) {real, imag} */,
  {32'hbf1d27f2, 32'h00000000} /* (9, 31, 15) {real, imag} */,
  {32'hbf54af39, 32'h00000000} /* (9, 31, 14) {real, imag} */,
  {32'hbf9f80d1, 32'h00000000} /* (9, 31, 13) {real, imag} */,
  {32'hbf640714, 32'h00000000} /* (9, 31, 12) {real, imag} */,
  {32'hbdd54342, 32'h00000000} /* (9, 31, 11) {real, imag} */,
  {32'h3f1e4b9e, 32'h00000000} /* (9, 31, 10) {real, imag} */,
  {32'h3eb03c0d, 32'h00000000} /* (9, 31, 9) {real, imag} */,
  {32'h3f22957f, 32'h00000000} /* (9, 31, 8) {real, imag} */,
  {32'h3f42a848, 32'h00000000} /* (9, 31, 7) {real, imag} */,
  {32'h3f166bf5, 32'h00000000} /* (9, 31, 6) {real, imag} */,
  {32'h3ebd7f50, 32'h00000000} /* (9, 31, 5) {real, imag} */,
  {32'h3eac836f, 32'h00000000} /* (9, 31, 4) {real, imag} */,
  {32'h3e9cb7d2, 32'h00000000} /* (9, 31, 3) {real, imag} */,
  {32'h3e3303af, 32'h00000000} /* (9, 31, 2) {real, imag} */,
  {32'h3e876340, 32'h00000000} /* (9, 31, 1) {real, imag} */,
  {32'h3e6b39a0, 32'h00000000} /* (9, 31, 0) {real, imag} */,
  {32'h3e92fe1e, 32'h00000000} /* (9, 30, 31) {real, imag} */,
  {32'h3f4c4182, 32'h00000000} /* (9, 30, 30) {real, imag} */,
  {32'h3f966b33, 32'h00000000} /* (9, 30, 29) {real, imag} */,
  {32'h3f591e1c, 32'h00000000} /* (9, 30, 28) {real, imag} */,
  {32'h3f88c312, 32'h00000000} /* (9, 30, 27) {real, imag} */,
  {32'h3f4d0a74, 32'h00000000} /* (9, 30, 26) {real, imag} */,
  {32'h3f4924b9, 32'h00000000} /* (9, 30, 25) {real, imag} */,
  {32'h3f9f3bef, 32'h00000000} /* (9, 30, 24) {real, imag} */,
  {32'h3f3dd2e4, 32'h00000000} /* (9, 30, 23) {real, imag} */,
  {32'h3f7b6e25, 32'h00000000} /* (9, 30, 22) {real, imag} */,
  {32'h3f369550, 32'h00000000} /* (9, 30, 21) {real, imag} */,
  {32'hbeb3dce2, 32'h00000000} /* (9, 30, 20) {real, imag} */,
  {32'hbeb2aed3, 32'h00000000} /* (9, 30, 19) {real, imag} */,
  {32'hbefa5c32, 32'h00000000} /* (9, 30, 18) {real, imag} */,
  {32'hbeb59ae2, 32'h00000000} /* (9, 30, 17) {real, imag} */,
  {32'hbf55c99b, 32'h00000000} /* (9, 30, 16) {real, imag} */,
  {32'hbf7c382d, 32'h00000000} /* (9, 30, 15) {real, imag} */,
  {32'hbf655efe, 32'h00000000} /* (9, 30, 14) {real, imag} */,
  {32'hbfb9d204, 32'h00000000} /* (9, 30, 13) {real, imag} */,
  {32'hbfa76851, 32'h00000000} /* (9, 30, 12) {real, imag} */,
  {32'hbe84edec, 32'h00000000} /* (9, 30, 11) {real, imag} */,
  {32'h3f6d6d86, 32'h00000000} /* (9, 30, 10) {real, imag} */,
  {32'h3f0f8b1c, 32'h00000000} /* (9, 30, 9) {real, imag} */,
  {32'h3f5c2de5, 32'h00000000} /* (9, 30, 8) {real, imag} */,
  {32'h3f912fe3, 32'h00000000} /* (9, 30, 7) {real, imag} */,
  {32'h3f0b89b6, 32'h00000000} /* (9, 30, 6) {real, imag} */,
  {32'h3f58f2ba, 32'h00000000} /* (9, 30, 5) {real, imag} */,
  {32'h3f7de5ce, 32'h00000000} /* (9, 30, 4) {real, imag} */,
  {32'h3f34e21f, 32'h00000000} /* (9, 30, 3) {real, imag} */,
  {32'h3eecf23e, 32'h00000000} /* (9, 30, 2) {real, imag} */,
  {32'h3f361d39, 32'h00000000} /* (9, 30, 1) {real, imag} */,
  {32'h3f09f2ae, 32'h00000000} /* (9, 30, 0) {real, imag} */,
  {32'h3f5f699f, 32'h00000000} /* (9, 29, 31) {real, imag} */,
  {32'h3fb349bd, 32'h00000000} /* (9, 29, 30) {real, imag} */,
  {32'h3f49ee8a, 32'h00000000} /* (9, 29, 29) {real, imag} */,
  {32'h3f2d9c06, 32'h00000000} /* (9, 29, 28) {real, imag} */,
  {32'h3f480483, 32'h00000000} /* (9, 29, 27) {real, imag} */,
  {32'h3f32f71b, 32'h00000000} /* (9, 29, 26) {real, imag} */,
  {32'h3f4f8a19, 32'h00000000} /* (9, 29, 25) {real, imag} */,
  {32'h3f83708c, 32'h00000000} /* (9, 29, 24) {real, imag} */,
  {32'h3f36c33a, 32'h00000000} /* (9, 29, 23) {real, imag} */,
  {32'h3f7a1cff, 32'h00000000} /* (9, 29, 22) {real, imag} */,
  {32'h3f36b3c7, 32'h00000000} /* (9, 29, 21) {real, imag} */,
  {32'hbe896b2e, 32'h00000000} /* (9, 29, 20) {real, imag} */,
  {32'hbeb98922, 32'h00000000} /* (9, 29, 19) {real, imag} */,
  {32'hbf080dcb, 32'h00000000} /* (9, 29, 18) {real, imag} */,
  {32'hbe888c68, 32'h00000000} /* (9, 29, 17) {real, imag} */,
  {32'hbf65b1bd, 32'h00000000} /* (9, 29, 16) {real, imag} */,
  {32'hbfe327c1, 32'h00000000} /* (9, 29, 15) {real, imag} */,
  {32'hbf8f0bb4, 32'h00000000} /* (9, 29, 14) {real, imag} */,
  {32'hbf791eac, 32'h00000000} /* (9, 29, 13) {real, imag} */,
  {32'hbf7190ad, 32'h00000000} /* (9, 29, 12) {real, imag} */,
  {32'hbf15f44b, 32'h00000000} /* (9, 29, 11) {real, imag} */,
  {32'h3ea79999, 32'h00000000} /* (9, 29, 10) {real, imag} */,
  {32'h3eba6edd, 32'h00000000} /* (9, 29, 9) {real, imag} */,
  {32'h3f33a04a, 32'h00000000} /* (9, 29, 8) {real, imag} */,
  {32'h3f338460, 32'h00000000} /* (9, 29, 7) {real, imag} */,
  {32'h3ea00269, 32'h00000000} /* (9, 29, 6) {real, imag} */,
  {32'h3ef94e02, 32'h00000000} /* (9, 29, 5) {real, imag} */,
  {32'h3f944c86, 32'h00000000} /* (9, 29, 4) {real, imag} */,
  {32'h3fa2bf75, 32'h00000000} /* (9, 29, 3) {real, imag} */,
  {32'h3f1964aa, 32'h00000000} /* (9, 29, 2) {real, imag} */,
  {32'h3f1dad70, 32'h00000000} /* (9, 29, 1) {real, imag} */,
  {32'h3e0fea6d, 32'h00000000} /* (9, 29, 0) {real, imag} */,
  {32'h3f863cc6, 32'h00000000} /* (9, 28, 31) {real, imag} */,
  {32'h3fa5fe3a, 32'h00000000} /* (9, 28, 30) {real, imag} */,
  {32'h3ec93b1f, 32'h00000000} /* (9, 28, 29) {real, imag} */,
  {32'h3e83912b, 32'h00000000} /* (9, 28, 28) {real, imag} */,
  {32'h3f0cf1fc, 32'h00000000} /* (9, 28, 27) {real, imag} */,
  {32'h3ecd2dae, 32'h00000000} /* (9, 28, 26) {real, imag} */,
  {32'h3f4aaddd, 32'h00000000} /* (9, 28, 25) {real, imag} */,
  {32'h3fba5ece, 32'h00000000} /* (9, 28, 24) {real, imag} */,
  {32'h3fa50eb6, 32'h00000000} /* (9, 28, 23) {real, imag} */,
  {32'h3fa20bf8, 32'h00000000} /* (9, 28, 22) {real, imag} */,
  {32'h3e829c5d, 32'h00000000} /* (9, 28, 21) {real, imag} */,
  {32'hbed40099, 32'h00000000} /* (9, 28, 20) {real, imag} */,
  {32'hbf2b9f37, 32'h00000000} /* (9, 28, 19) {real, imag} */,
  {32'hbf1fc841, 32'h00000000} /* (9, 28, 18) {real, imag} */,
  {32'hbf0c3ba1, 32'h00000000} /* (9, 28, 17) {real, imag} */,
  {32'hbf89b72f, 32'h00000000} /* (9, 28, 16) {real, imag} */,
  {32'hbfe8727d, 32'h00000000} /* (9, 28, 15) {real, imag} */,
  {32'hbf9d7746, 32'h00000000} /* (9, 28, 14) {real, imag} */,
  {32'hbf59816e, 32'h00000000} /* (9, 28, 13) {real, imag} */,
  {32'hbf59547c, 32'h00000000} /* (9, 28, 12) {real, imag} */,
  {32'hbf79b61c, 32'h00000000} /* (9, 28, 11) {real, imag} */,
  {32'h3f0f993b, 32'h00000000} /* (9, 28, 10) {real, imag} */,
  {32'h3f71eace, 32'h00000000} /* (9, 28, 9) {real, imag} */,
  {32'h3f70400e, 32'h00000000} /* (9, 28, 8) {real, imag} */,
  {32'h3f34affe, 32'h00000000} /* (9, 28, 7) {real, imag} */,
  {32'h3f017746, 32'h00000000} /* (9, 28, 6) {real, imag} */,
  {32'h3f6354df, 32'h00000000} /* (9, 28, 5) {real, imag} */,
  {32'h3fa660bf, 32'h00000000} /* (9, 28, 4) {real, imag} */,
  {32'h3faddc6f, 32'h00000000} /* (9, 28, 3) {real, imag} */,
  {32'h3f275195, 32'h00000000} /* (9, 28, 2) {real, imag} */,
  {32'h3f2a783a, 32'h00000000} /* (9, 28, 1) {real, imag} */,
  {32'h3eb0b4f3, 32'h00000000} /* (9, 28, 0) {real, imag} */,
  {32'h3f190bb3, 32'h00000000} /* (9, 27, 31) {real, imag} */,
  {32'h3f4f115b, 32'h00000000} /* (9, 27, 30) {real, imag} */,
  {32'h3f52ef32, 32'h00000000} /* (9, 27, 29) {real, imag} */,
  {32'h3ef3bf25, 32'h00000000} /* (9, 27, 28) {real, imag} */,
  {32'h3f400776, 32'h00000000} /* (9, 27, 27) {real, imag} */,
  {32'h3f8d5c13, 32'h00000000} /* (9, 27, 26) {real, imag} */,
  {32'h3fea9992, 32'h00000000} /* (9, 27, 25) {real, imag} */,
  {32'h3fca6ada, 32'h00000000} /* (9, 27, 24) {real, imag} */,
  {32'h3f9d4240, 32'h00000000} /* (9, 27, 23) {real, imag} */,
  {32'h3f3dcb74, 32'h00000000} /* (9, 27, 22) {real, imag} */,
  {32'hbe3e29f8, 32'h00000000} /* (9, 27, 21) {real, imag} */,
  {32'hbf865fd8, 32'h00000000} /* (9, 27, 20) {real, imag} */,
  {32'hbf6b1423, 32'h00000000} /* (9, 27, 19) {real, imag} */,
  {32'hbf1e6a54, 32'h00000000} /* (9, 27, 18) {real, imag} */,
  {32'hbf5a590e, 32'h00000000} /* (9, 27, 17) {real, imag} */,
  {32'hbfa8c49a, 32'h00000000} /* (9, 27, 16) {real, imag} */,
  {32'hbfa297f0, 32'h00000000} /* (9, 27, 15) {real, imag} */,
  {32'hbf4713af, 32'h00000000} /* (9, 27, 14) {real, imag} */,
  {32'hbf5eca42, 32'h00000000} /* (9, 27, 13) {real, imag} */,
  {32'hbf558e75, 32'h00000000} /* (9, 27, 12) {real, imag} */,
  {32'hbf80ab61, 32'h00000000} /* (9, 27, 11) {real, imag} */,
  {32'h3e6121ca, 32'h00000000} /* (9, 27, 10) {real, imag} */,
  {32'h3f7999a2, 32'h00000000} /* (9, 27, 9) {real, imag} */,
  {32'h3f8aec1e, 32'h00000000} /* (9, 27, 8) {real, imag} */,
  {32'h3fb476ef, 32'h00000000} /* (9, 27, 7) {real, imag} */,
  {32'h3f85c455, 32'h00000000} /* (9, 27, 6) {real, imag} */,
  {32'h3fb6da75, 32'h00000000} /* (9, 27, 5) {real, imag} */,
  {32'h3fbf88d7, 32'h00000000} /* (9, 27, 4) {real, imag} */,
  {32'h3f8144e3, 32'h00000000} /* (9, 27, 3) {real, imag} */,
  {32'h3f42b1a3, 32'h00000000} /* (9, 27, 2) {real, imag} */,
  {32'h3f81f04a, 32'h00000000} /* (9, 27, 1) {real, imag} */,
  {32'h3f375d98, 32'h00000000} /* (9, 27, 0) {real, imag} */,
  {32'h3f0759c2, 32'h00000000} /* (9, 26, 31) {real, imag} */,
  {32'h3f53e04f, 32'h00000000} /* (9, 26, 30) {real, imag} */,
  {32'h3fc1aaf6, 32'h00000000} /* (9, 26, 29) {real, imag} */,
  {32'h3f93e724, 32'h00000000} /* (9, 26, 28) {real, imag} */,
  {32'h3ede5ab6, 32'h00000000} /* (9, 26, 27) {real, imag} */,
  {32'h3f83e64f, 32'h00000000} /* (9, 26, 26) {real, imag} */,
  {32'h3fdef5ac, 32'h00000000} /* (9, 26, 25) {real, imag} */,
  {32'h3fbc4b13, 32'h00000000} /* (9, 26, 24) {real, imag} */,
  {32'h3f1af56e, 32'h00000000} /* (9, 26, 23) {real, imag} */,
  {32'h3f108fed, 32'h00000000} /* (9, 26, 22) {real, imag} */,
  {32'h3eaeb914, 32'h00000000} /* (9, 26, 21) {real, imag} */,
  {32'hbf80c830, 32'h00000000} /* (9, 26, 20) {real, imag} */,
  {32'hbfa911ab, 32'h00000000} /* (9, 26, 19) {real, imag} */,
  {32'hbf583e82, 32'h00000000} /* (9, 26, 18) {real, imag} */,
  {32'hbf6e1ccf, 32'h00000000} /* (9, 26, 17) {real, imag} */,
  {32'hbf948b5f, 32'h00000000} /* (9, 26, 16) {real, imag} */,
  {32'hbf5704c3, 32'h00000000} /* (9, 26, 15) {real, imag} */,
  {32'hbf10a1eb, 32'h00000000} /* (9, 26, 14) {real, imag} */,
  {32'hbf38e36a, 32'h00000000} /* (9, 26, 13) {real, imag} */,
  {32'hbedd9b9e, 32'h00000000} /* (9, 26, 12) {real, imag} */,
  {32'hbea7551d, 32'h00000000} /* (9, 26, 11) {real, imag} */,
  {32'h3e9dd0d7, 32'h00000000} /* (9, 26, 10) {real, imag} */,
  {32'h3fa424d8, 32'h00000000} /* (9, 26, 9) {real, imag} */,
  {32'h3f904332, 32'h00000000} /* (9, 26, 8) {real, imag} */,
  {32'h3f93949c, 32'h00000000} /* (9, 26, 7) {real, imag} */,
  {32'h3f8f3ba9, 32'h00000000} /* (9, 26, 6) {real, imag} */,
  {32'h3f956403, 32'h00000000} /* (9, 26, 5) {real, imag} */,
  {32'h3fa032ab, 32'h00000000} /* (9, 26, 4) {real, imag} */,
  {32'h3f7e1f5b, 32'h00000000} /* (9, 26, 3) {real, imag} */,
  {32'h3f900921, 32'h00000000} /* (9, 26, 2) {real, imag} */,
  {32'h3f974d8e, 32'h00000000} /* (9, 26, 1) {real, imag} */,
  {32'h3f3bf1e6, 32'h00000000} /* (9, 26, 0) {real, imag} */,
  {32'h3f2e4076, 32'h00000000} /* (9, 25, 31) {real, imag} */,
  {32'h3f8174ca, 32'h00000000} /* (9, 25, 30) {real, imag} */,
  {32'h3faa0271, 32'h00000000} /* (9, 25, 29) {real, imag} */,
  {32'h3fc8e4e8, 32'h00000000} /* (9, 25, 28) {real, imag} */,
  {32'h3e9ab506, 32'h00000000} /* (9, 25, 27) {real, imag} */,
  {32'h3eed2c61, 32'h00000000} /* (9, 25, 26) {real, imag} */,
  {32'h3f87c7ca, 32'h00000000} /* (9, 25, 25) {real, imag} */,
  {32'h3f6a693e, 32'h00000000} /* (9, 25, 24) {real, imag} */,
  {32'h3ec7531b, 32'h00000000} /* (9, 25, 23) {real, imag} */,
  {32'h3e90af14, 32'h00000000} /* (9, 25, 22) {real, imag} */,
  {32'h3eac3143, 32'h00000000} /* (9, 25, 21) {real, imag} */,
  {32'hbf2bdb47, 32'h00000000} /* (9, 25, 20) {real, imag} */,
  {32'hbf724635, 32'h00000000} /* (9, 25, 19) {real, imag} */,
  {32'hbf66f4cf, 32'h00000000} /* (9, 25, 18) {real, imag} */,
  {32'hbf84a531, 32'h00000000} /* (9, 25, 17) {real, imag} */,
  {32'hbf52fe79, 32'h00000000} /* (9, 25, 16) {real, imag} */,
  {32'hbf4265cd, 32'h00000000} /* (9, 25, 15) {real, imag} */,
  {32'hbf37d3a5, 32'h00000000} /* (9, 25, 14) {real, imag} */,
  {32'hbf36d35c, 32'h00000000} /* (9, 25, 13) {real, imag} */,
  {32'hbeb78723, 32'h00000000} /* (9, 25, 12) {real, imag} */,
  {32'hbf0b4d3c, 32'h00000000} /* (9, 25, 11) {real, imag} */,
  {32'h3f11d698, 32'h00000000} /* (9, 25, 10) {real, imag} */,
  {32'h3fb94be1, 32'h00000000} /* (9, 25, 9) {real, imag} */,
  {32'h3f5a4b6b, 32'h00000000} /* (9, 25, 8) {real, imag} */,
  {32'h3f713e9d, 32'h00000000} /* (9, 25, 7) {real, imag} */,
  {32'h3fba3743, 32'h00000000} /* (9, 25, 6) {real, imag} */,
  {32'h3fdf9c0b, 32'h00000000} /* (9, 25, 5) {real, imag} */,
  {32'h3fce14a7, 32'h00000000} /* (9, 25, 4) {real, imag} */,
  {32'h3f9fc377, 32'h00000000} /* (9, 25, 3) {real, imag} */,
  {32'h3f83da05, 32'h00000000} /* (9, 25, 2) {real, imag} */,
  {32'h3f90b9c7, 32'h00000000} /* (9, 25, 1) {real, imag} */,
  {32'h3f4a0a28, 32'h00000000} /* (9, 25, 0) {real, imag} */,
  {32'h3f1c817a, 32'h00000000} /* (9, 24, 31) {real, imag} */,
  {32'h3fa5f2cc, 32'h00000000} /* (9, 24, 30) {real, imag} */,
  {32'h3f0eacea, 32'h00000000} /* (9, 24, 29) {real, imag} */,
  {32'h3f1eae80, 32'h00000000} /* (9, 24, 28) {real, imag} */,
  {32'h3ee1dcb0, 32'h00000000} /* (9, 24, 27) {real, imag} */,
  {32'h3f127712, 32'h00000000} /* (9, 24, 26) {real, imag} */,
  {32'h3f1bfdda, 32'h00000000} /* (9, 24, 25) {real, imag} */,
  {32'h3ef617ce, 32'h00000000} /* (9, 24, 24) {real, imag} */,
  {32'h3ea514f2, 32'h00000000} /* (9, 24, 23) {real, imag} */,
  {32'h3c826edf, 32'h00000000} /* (9, 24, 22) {real, imag} */,
  {32'hbdedd6b9, 32'h00000000} /* (9, 24, 21) {real, imag} */,
  {32'hbf83a89d, 32'h00000000} /* (9, 24, 20) {real, imag} */,
  {32'hbf744ace, 32'h00000000} /* (9, 24, 19) {real, imag} */,
  {32'hbe6859b5, 32'h00000000} /* (9, 24, 18) {real, imag} */,
  {32'h3dbabab1, 32'h00000000} /* (9, 24, 17) {real, imag} */,
  {32'hbec6c522, 32'h00000000} /* (9, 24, 16) {real, imag} */,
  {32'hbf8fadc3, 32'h00000000} /* (9, 24, 15) {real, imag} */,
  {32'hbf1d0b61, 32'h00000000} /* (9, 24, 14) {real, imag} */,
  {32'hbf25570e, 32'h00000000} /* (9, 24, 13) {real, imag} */,
  {32'hbfa45f78, 32'h00000000} /* (9, 24, 12) {real, imag} */,
  {32'hbf8c5431, 32'h00000000} /* (9, 24, 11) {real, imag} */,
  {32'h3f9a73a1, 32'h00000000} /* (9, 24, 10) {real, imag} */,
  {32'h3fbdf12d, 32'h00000000} /* (9, 24, 9) {real, imag} */,
  {32'h3f8982bf, 32'h00000000} /* (9, 24, 8) {real, imag} */,
  {32'h3fa3abae, 32'h00000000} /* (9, 24, 7) {real, imag} */,
  {32'h3fa94254, 32'h00000000} /* (9, 24, 6) {real, imag} */,
  {32'h3fa7514b, 32'h00000000} /* (9, 24, 5) {real, imag} */,
  {32'h3fa158a7, 32'h00000000} /* (9, 24, 4) {real, imag} */,
  {32'h3f9282fb, 32'h00000000} /* (9, 24, 3) {real, imag} */,
  {32'h3f8da6a1, 32'h00000000} /* (9, 24, 2) {real, imag} */,
  {32'h3f57ff6c, 32'h00000000} /* (9, 24, 1) {real, imag} */,
  {32'h3efb5443, 32'h00000000} /* (9, 24, 0) {real, imag} */,
  {32'h3ea7fea4, 32'h00000000} /* (9, 23, 31) {real, imag} */,
  {32'h3f51cb90, 32'h00000000} /* (9, 23, 30) {real, imag} */,
  {32'h3f2edd7d, 32'h00000000} /* (9, 23, 29) {real, imag} */,
  {32'h3f30d67c, 32'h00000000} /* (9, 23, 28) {real, imag} */,
  {32'h3f0845b5, 32'h00000000} /* (9, 23, 27) {real, imag} */,
  {32'h3ed96321, 32'h00000000} /* (9, 23, 26) {real, imag} */,
  {32'h3e85d4a8, 32'h00000000} /* (9, 23, 25) {real, imag} */,
  {32'h3f2992b5, 32'h00000000} /* (9, 23, 24) {real, imag} */,
  {32'h3f8e9fa5, 32'h00000000} /* (9, 23, 23) {real, imag} */,
  {32'h3eee0ae0, 32'h00000000} /* (9, 23, 22) {real, imag} */,
  {32'h3e183475, 32'h00000000} /* (9, 23, 21) {real, imag} */,
  {32'hbf5f851e, 32'h00000000} /* (9, 23, 20) {real, imag} */,
  {32'hbf8e8e49, 32'h00000000} /* (9, 23, 19) {real, imag} */,
  {32'hbf47d93b, 32'h00000000} /* (9, 23, 18) {real, imag} */,
  {32'hbee8f359, 32'h00000000} /* (9, 23, 17) {real, imag} */,
  {32'hbecc489d, 32'h00000000} /* (9, 23, 16) {real, imag} */,
  {32'hbf1fb13c, 32'h00000000} /* (9, 23, 15) {real, imag} */,
  {32'hbf266468, 32'h00000000} /* (9, 23, 14) {real, imag} */,
  {32'hbf4650ec, 32'h00000000} /* (9, 23, 13) {real, imag} */,
  {32'hbf85ac3b, 32'h00000000} /* (9, 23, 12) {real, imag} */,
  {32'hbf91e600, 32'h00000000} /* (9, 23, 11) {real, imag} */,
  {32'h3f165803, 32'h00000000} /* (9, 23, 10) {real, imag} */,
  {32'h3f8f9054, 32'h00000000} /* (9, 23, 9) {real, imag} */,
  {32'h3f97f25b, 32'h00000000} /* (9, 23, 8) {real, imag} */,
  {32'h3fa46e22, 32'h00000000} /* (9, 23, 7) {real, imag} */,
  {32'h3f8a39fd, 32'h00000000} /* (9, 23, 6) {real, imag} */,
  {32'h3f565e0c, 32'h00000000} /* (9, 23, 5) {real, imag} */,
  {32'h3f864ffb, 32'h00000000} /* (9, 23, 4) {real, imag} */,
  {32'h3f8678e0, 32'h00000000} /* (9, 23, 3) {real, imag} */,
  {32'h3f6deb6f, 32'h00000000} /* (9, 23, 2) {real, imag} */,
  {32'h3f486f12, 32'h00000000} /* (9, 23, 1) {real, imag} */,
  {32'h3e9fb806, 32'h00000000} /* (9, 23, 0) {real, imag} */,
  {32'h3e9055f7, 32'h00000000} /* (9, 22, 31) {real, imag} */,
  {32'h3f7ce15d, 32'h00000000} /* (9, 22, 30) {real, imag} */,
  {32'h3fb0c5a8, 32'h00000000} /* (9, 22, 29) {real, imag} */,
  {32'h3f6af535, 32'h00000000} /* (9, 22, 28) {real, imag} */,
  {32'h3eb7c595, 32'h00000000} /* (9, 22, 27) {real, imag} */,
  {32'h3f40869f, 32'h00000000} /* (9, 22, 26) {real, imag} */,
  {32'h3f6833b2, 32'h00000000} /* (9, 22, 25) {real, imag} */,
  {32'h3f79904f, 32'h00000000} /* (9, 22, 24) {real, imag} */,
  {32'h3fb35e13, 32'h00000000} /* (9, 22, 23) {real, imag} */,
  {32'h3f443b94, 32'h00000000} /* (9, 22, 22) {real, imag} */,
  {32'h3f12cec8, 32'h00000000} /* (9, 22, 21) {real, imag} */,
  {32'hbf3b8fc5, 32'h00000000} /* (9, 22, 20) {real, imag} */,
  {32'hbf8708a7, 32'h00000000} /* (9, 22, 19) {real, imag} */,
  {32'hbfa9cdd5, 32'h00000000} /* (9, 22, 18) {real, imag} */,
  {32'hbf63a142, 32'h00000000} /* (9, 22, 17) {real, imag} */,
  {32'hbeb997c3, 32'h00000000} /* (9, 22, 16) {real, imag} */,
  {32'hbee64e6a, 32'h00000000} /* (9, 22, 15) {real, imag} */,
  {32'hbf76c539, 32'h00000000} /* (9, 22, 14) {real, imag} */,
  {32'hbf483a35, 32'h00000000} /* (9, 22, 13) {real, imag} */,
  {32'hbed8e5bb, 32'h00000000} /* (9, 22, 12) {real, imag} */,
  {32'hbe9eb8fd, 32'h00000000} /* (9, 22, 11) {real, imag} */,
  {32'h3eff0d92, 32'h00000000} /* (9, 22, 10) {real, imag} */,
  {32'h3f06dec5, 32'h00000000} /* (9, 22, 9) {real, imag} */,
  {32'h3ed048c2, 32'h00000000} /* (9, 22, 8) {real, imag} */,
  {32'h3f11dd57, 32'h00000000} /* (9, 22, 7) {real, imag} */,
  {32'h3f4214cc, 32'h00000000} /* (9, 22, 6) {real, imag} */,
  {32'h3f8335e5, 32'h00000000} /* (9, 22, 5) {real, imag} */,
  {32'h3f78317a, 32'h00000000} /* (9, 22, 4) {real, imag} */,
  {32'h3fb47f9a, 32'h00000000} /* (9, 22, 3) {real, imag} */,
  {32'h3fcdd56c, 32'h00000000} /* (9, 22, 2) {real, imag} */,
  {32'h3f40fe0f, 32'h00000000} /* (9, 22, 1) {real, imag} */,
  {32'h3e4a94d9, 32'h00000000} /* (9, 22, 0) {real, imag} */,
  {32'h3e6b29a3, 32'h00000000} /* (9, 21, 31) {real, imag} */,
  {32'h3ed21ad2, 32'h00000000} /* (9, 21, 30) {real, imag} */,
  {32'h3e6acc32, 32'h00000000} /* (9, 21, 29) {real, imag} */,
  {32'hbd118772, 32'h00000000} /* (9, 21, 28) {real, imag} */,
  {32'hbcd2bf52, 32'h00000000} /* (9, 21, 27) {real, imag} */,
  {32'h3eef61fa, 32'h00000000} /* (9, 21, 26) {real, imag} */,
  {32'h3f269a97, 32'h00000000} /* (9, 21, 25) {real, imag} */,
  {32'h3ee864df, 32'h00000000} /* (9, 21, 24) {real, imag} */,
  {32'h3ef8ba56, 32'h00000000} /* (9, 21, 23) {real, imag} */,
  {32'h3f107783, 32'h00000000} /* (9, 21, 22) {real, imag} */,
  {32'h3f6e5d93, 32'h00000000} /* (9, 21, 21) {real, imag} */,
  {32'hbf2849fa, 32'h00000000} /* (9, 21, 20) {real, imag} */,
  {32'hbf88690d, 32'h00000000} /* (9, 21, 19) {real, imag} */,
  {32'hbf1c51d5, 32'h00000000} /* (9, 21, 18) {real, imag} */,
  {32'hbead26b1, 32'h00000000} /* (9, 21, 17) {real, imag} */,
  {32'h3e1ea82e, 32'h00000000} /* (9, 21, 16) {real, imag} */,
  {32'hbe831877, 32'h00000000} /* (9, 21, 15) {real, imag} */,
  {32'hbed7c02c, 32'h00000000} /* (9, 21, 14) {real, imag} */,
  {32'hbd0cdaed, 32'h00000000} /* (9, 21, 13) {real, imag} */,
  {32'h3dd2e4fb, 32'h00000000} /* (9, 21, 12) {real, imag} */,
  {32'hbe4136c0, 32'h00000000} /* (9, 21, 11) {real, imag} */,
  {32'h3ebf1224, 32'h00000000} /* (9, 21, 10) {real, imag} */,
  {32'h3e908a0b, 32'h00000000} /* (9, 21, 9) {real, imag} */,
  {32'h3ce093d0, 32'h00000000} /* (9, 21, 8) {real, imag} */,
  {32'h3b4b0332, 32'h00000000} /* (9, 21, 7) {real, imag} */,
  {32'h3de93c6d, 32'h00000000} /* (9, 21, 6) {real, imag} */,
  {32'h3f1c7ddc, 32'h00000000} /* (9, 21, 5) {real, imag} */,
  {32'h3edc43d4, 32'h00000000} /* (9, 21, 4) {real, imag} */,
  {32'h3f194310, 32'h00000000} /* (9, 21, 3) {real, imag} */,
  {32'h3f9b8c8d, 32'h00000000} /* (9, 21, 2) {real, imag} */,
  {32'h3ea1447e, 32'h00000000} /* (9, 21, 1) {real, imag} */,
  {32'h3d82bd31, 32'h00000000} /* (9, 21, 0) {real, imag} */,
  {32'hbeb596a2, 32'h00000000} /* (9, 20, 31) {real, imag} */,
  {32'hbf5487e0, 32'h00000000} /* (9, 20, 30) {real, imag} */,
  {32'hbf5f50c3, 32'h00000000} /* (9, 20, 29) {real, imag} */,
  {32'hbf2b8e36, 32'h00000000} /* (9, 20, 28) {real, imag} */,
  {32'hbf0d43ba, 32'h00000000} /* (9, 20, 27) {real, imag} */,
  {32'hbf08f308, 32'h00000000} /* (9, 20, 26) {real, imag} */,
  {32'hbf1718b1, 32'h00000000} /* (9, 20, 25) {real, imag} */,
  {32'hbf32cced, 32'h00000000} /* (9, 20, 24) {real, imag} */,
  {32'hbf0327ee, 32'h00000000} /* (9, 20, 23) {real, imag} */,
  {32'hbe8d28c9, 32'h00000000} /* (9, 20, 22) {real, imag} */,
  {32'h3d8b58d0, 32'h00000000} /* (9, 20, 21) {real, imag} */,
  {32'h3f09b54c, 32'h00000000} /* (9, 20, 20) {real, imag} */,
  {32'h3d92e694, 32'h00000000} /* (9, 20, 19) {real, imag} */,
  {32'hbd2d1a55, 32'h00000000} /* (9, 20, 18) {real, imag} */,
  {32'h3e8de845, 32'h00000000} /* (9, 20, 17) {real, imag} */,
  {32'h3f36834c, 32'h00000000} /* (9, 20, 16) {real, imag} */,
  {32'h3f13e512, 32'h00000000} /* (9, 20, 15) {real, imag} */,
  {32'h3f3ecd25, 32'h00000000} /* (9, 20, 14) {real, imag} */,
  {32'h3f86e592, 32'h00000000} /* (9, 20, 13) {real, imag} */,
  {32'h3f84ed34, 32'h00000000} /* (9, 20, 12) {real, imag} */,
  {32'h3f257d50, 32'h00000000} /* (9, 20, 11) {real, imag} */,
  {32'hbdbd481e, 32'h00000000} /* (9, 20, 10) {real, imag} */,
  {32'hbf1e241a, 32'h00000000} /* (9, 20, 9) {real, imag} */,
  {32'hbf713d1b, 32'h00000000} /* (9, 20, 8) {real, imag} */,
  {32'hbf88612f, 32'h00000000} /* (9, 20, 7) {real, imag} */,
  {32'hbf431e66, 32'h00000000} /* (9, 20, 6) {real, imag} */,
  {32'hbeb44428, 32'h00000000} /* (9, 20, 5) {real, imag} */,
  {32'hbf0ffd26, 32'h00000000} /* (9, 20, 4) {real, imag} */,
  {32'hbf40c207, 32'h00000000} /* (9, 20, 3) {real, imag} */,
  {32'hbed8dd2d, 32'h00000000} /* (9, 20, 2) {real, imag} */,
  {32'hbf704e6d, 32'h00000000} /* (9, 20, 1) {real, imag} */,
  {32'hbebbb1ab, 32'h00000000} /* (9, 20, 0) {real, imag} */,
  {32'hbf40e88c, 32'h00000000} /* (9, 19, 31) {real, imag} */,
  {32'hbf9803ae, 32'h00000000} /* (9, 19, 30) {real, imag} */,
  {32'hbf66bb63, 32'h00000000} /* (9, 19, 29) {real, imag} */,
  {32'hbf26be6c, 32'h00000000} /* (9, 19, 28) {real, imag} */,
  {32'hbf3b87e3, 32'h00000000} /* (9, 19, 27) {real, imag} */,
  {32'hbf5b1fe8, 32'h00000000} /* (9, 19, 26) {real, imag} */,
  {32'hbf066be4, 32'h00000000} /* (9, 19, 25) {real, imag} */,
  {32'hbf7500c1, 32'h00000000} /* (9, 19, 24) {real, imag} */,
  {32'hbf82401b, 32'h00000000} /* (9, 19, 23) {real, imag} */,
  {32'hbf823e65, 32'h00000000} /* (9, 19, 22) {real, imag} */,
  {32'hbee4da3f, 32'h00000000} /* (9, 19, 21) {real, imag} */,
  {32'h3f538006, 32'h00000000} /* (9, 19, 20) {real, imag} */,
  {32'h3f19b4ff, 32'h00000000} /* (9, 19, 19) {real, imag} */,
  {32'h3dcabb10, 32'h00000000} /* (9, 19, 18) {real, imag} */,
  {32'h3ec1b50e, 32'h00000000} /* (9, 19, 17) {real, imag} */,
  {32'h3fa26a36, 32'h00000000} /* (9, 19, 16) {real, imag} */,
  {32'h3fa4d181, 32'h00000000} /* (9, 19, 15) {real, imag} */,
  {32'h3fc07553, 32'h00000000} /* (9, 19, 14) {real, imag} */,
  {32'h3f958be2, 32'h00000000} /* (9, 19, 13) {real, imag} */,
  {32'h3f557643, 32'h00000000} /* (9, 19, 12) {real, imag} */,
  {32'h3f4ce44e, 32'h00000000} /* (9, 19, 11) {real, imag} */,
  {32'hbe9c0044, 32'h00000000} /* (9, 19, 10) {real, imag} */,
  {32'hbf898958, 32'h00000000} /* (9, 19, 9) {real, imag} */,
  {32'hbfc0a0de, 32'h00000000} /* (9, 19, 8) {real, imag} */,
  {32'hbfb95000, 32'h00000000} /* (9, 19, 7) {real, imag} */,
  {32'hbf8fca91, 32'h00000000} /* (9, 19, 6) {real, imag} */,
  {32'hbf77be4e, 32'h00000000} /* (9, 19, 5) {real, imag} */,
  {32'hbf5f4019, 32'h00000000} /* (9, 19, 4) {real, imag} */,
  {32'hbf7c8dbe, 32'h00000000} /* (9, 19, 3) {real, imag} */,
  {32'hbf5273d7, 32'h00000000} /* (9, 19, 2) {real, imag} */,
  {32'hbf5a2ee7, 32'h00000000} /* (9, 19, 1) {real, imag} */,
  {32'hbeb8fab5, 32'h00000000} /* (9, 19, 0) {real, imag} */,
  {32'hbf88e0b9, 32'h00000000} /* (9, 18, 31) {real, imag} */,
  {32'hbfa86255, 32'h00000000} /* (9, 18, 30) {real, imag} */,
  {32'hbf700652, 32'h00000000} /* (9, 18, 29) {real, imag} */,
  {32'hbf6506c2, 32'h00000000} /* (9, 18, 28) {real, imag} */,
  {32'hbf54a776, 32'h00000000} /* (9, 18, 27) {real, imag} */,
  {32'hbf2381d8, 32'h00000000} /* (9, 18, 26) {real, imag} */,
  {32'hbf2ecd87, 32'h00000000} /* (9, 18, 25) {real, imag} */,
  {32'hbfb76ded, 32'h00000000} /* (9, 18, 24) {real, imag} */,
  {32'hbfa68c0b, 32'h00000000} /* (9, 18, 23) {real, imag} */,
  {32'hbf26d20a, 32'h00000000} /* (9, 18, 22) {real, imag} */,
  {32'hbe5ca900, 32'h00000000} /* (9, 18, 21) {real, imag} */,
  {32'h3f9fd3cb, 32'h00000000} /* (9, 18, 20) {real, imag} */,
  {32'h3f581aad, 32'h00000000} /* (9, 18, 19) {real, imag} */,
  {32'h3dcccf35, 32'h00000000} /* (9, 18, 18) {real, imag} */,
  {32'h3f03a09b, 32'h00000000} /* (9, 18, 17) {real, imag} */,
  {32'h3fc3ed01, 32'h00000000} /* (9, 18, 16) {real, imag} */,
  {32'h3fa882ff, 32'h00000000} /* (9, 18, 15) {real, imag} */,
  {32'h3f9d11a7, 32'h00000000} /* (9, 18, 14) {real, imag} */,
  {32'h3fb4a5fe, 32'h00000000} /* (9, 18, 13) {real, imag} */,
  {32'h3fac779d, 32'h00000000} /* (9, 18, 12) {real, imag} */,
  {32'h3f4dfb09, 32'h00000000} /* (9, 18, 11) {real, imag} */,
  {32'hbf014abe, 32'h00000000} /* (9, 18, 10) {real, imag} */,
  {32'hbf736d00, 32'h00000000} /* (9, 18, 9) {real, imag} */,
  {32'hbf89dbf0, 32'h00000000} /* (9, 18, 8) {real, imag} */,
  {32'hbf5f19e1, 32'h00000000} /* (9, 18, 7) {real, imag} */,
  {32'hbf5e5db9, 32'h00000000} /* (9, 18, 6) {real, imag} */,
  {32'hbf6497f9, 32'h00000000} /* (9, 18, 5) {real, imag} */,
  {32'hbf78079b, 32'h00000000} /* (9, 18, 4) {real, imag} */,
  {32'hbf9bb0c1, 32'h00000000} /* (9, 18, 3) {real, imag} */,
  {32'hbf5bbad1, 32'h00000000} /* (9, 18, 2) {real, imag} */,
  {32'hbf7a4420, 32'h00000000} /* (9, 18, 1) {real, imag} */,
  {32'hbf46958b, 32'h00000000} /* (9, 18, 0) {real, imag} */,
  {32'hbf6b4071, 32'h00000000} /* (9, 17, 31) {real, imag} */,
  {32'hbfd41af0, 32'h00000000} /* (9, 17, 30) {real, imag} */,
  {32'hbfbae76d, 32'h00000000} /* (9, 17, 29) {real, imag} */,
  {32'hbfc1f17d, 32'h00000000} /* (9, 17, 28) {real, imag} */,
  {32'hbfacb944, 32'h00000000} /* (9, 17, 27) {real, imag} */,
  {32'hbf632277, 32'h00000000} /* (9, 17, 26) {real, imag} */,
  {32'hbf5df5d6, 32'h00000000} /* (9, 17, 25) {real, imag} */,
  {32'hbfcfed25, 32'h00000000} /* (9, 17, 24) {real, imag} */,
  {32'hbfbf7f89, 32'h00000000} /* (9, 17, 23) {real, imag} */,
  {32'hbf341c3b, 32'h00000000} /* (9, 17, 22) {real, imag} */,
  {32'h3d1aeb66, 32'h00000000} /* (9, 17, 21) {real, imag} */,
  {32'h3fa0f94a, 32'h00000000} /* (9, 17, 20) {real, imag} */,
  {32'h3f5a8fd1, 32'h00000000} /* (9, 17, 19) {real, imag} */,
  {32'h3ee97f51, 32'h00000000} /* (9, 17, 18) {real, imag} */,
  {32'h3f56fa3c, 32'h00000000} /* (9, 17, 17) {real, imag} */,
  {32'h3f52fdfb, 32'h00000000} /* (9, 17, 16) {real, imag} */,
  {32'h3f1f5d68, 32'h00000000} /* (9, 17, 15) {real, imag} */,
  {32'h3f0d96e7, 32'h00000000} /* (9, 17, 14) {real, imag} */,
  {32'h3f4d9c00, 32'h00000000} /* (9, 17, 13) {real, imag} */,
  {32'h3f42d3a9, 32'h00000000} /* (9, 17, 12) {real, imag} */,
  {32'h3ed3ddce, 32'h00000000} /* (9, 17, 11) {real, imag} */,
  {32'hbf1c6f7e, 32'h00000000} /* (9, 17, 10) {real, imag} */,
  {32'hbf966641, 32'h00000000} /* (9, 17, 9) {real, imag} */,
  {32'hbfa4b575, 32'h00000000} /* (9, 17, 8) {real, imag} */,
  {32'hbf17dbec, 32'h00000000} /* (9, 17, 7) {real, imag} */,
  {32'hbf72703d, 32'h00000000} /* (9, 17, 6) {real, imag} */,
  {32'hbf8116d4, 32'h00000000} /* (9, 17, 5) {real, imag} */,
  {32'hbf5b123d, 32'h00000000} /* (9, 17, 4) {real, imag} */,
  {32'hbfb0128d, 32'h00000000} /* (9, 17, 3) {real, imag} */,
  {32'hbfb1176c, 32'h00000000} /* (9, 17, 2) {real, imag} */,
  {32'hbf47ed76, 32'h00000000} /* (9, 17, 1) {real, imag} */,
  {32'hbed508cd, 32'h00000000} /* (9, 17, 0) {real, imag} */,
  {32'hbf15c580, 32'h00000000} /* (9, 16, 31) {real, imag} */,
  {32'hbfd4c929, 32'h00000000} /* (9, 16, 30) {real, imag} */,
  {32'hbf97dfd9, 32'h00000000} /* (9, 16, 29) {real, imag} */,
  {32'hbfbab4a5, 32'h00000000} /* (9, 16, 28) {real, imag} */,
  {32'hbfa7ae63, 32'h00000000} /* (9, 16, 27) {real, imag} */,
  {32'hbf41daf4, 32'h00000000} /* (9, 16, 26) {real, imag} */,
  {32'hbf47fa13, 32'h00000000} /* (9, 16, 25) {real, imag} */,
  {32'hbf6d913f, 32'h00000000} /* (9, 16, 24) {real, imag} */,
  {32'hbf8ff4dd, 32'h00000000} /* (9, 16, 23) {real, imag} */,
  {32'hbf6a1c6e, 32'h00000000} /* (9, 16, 22) {real, imag} */,
  {32'hbcd9a434, 32'h00000000} /* (9, 16, 21) {real, imag} */,
  {32'h3f25936d, 32'h00000000} /* (9, 16, 20) {real, imag} */,
  {32'h3f25d142, 32'h00000000} /* (9, 16, 19) {real, imag} */,
  {32'h3f80a054, 32'h00000000} /* (9, 16, 18) {real, imag} */,
  {32'h3f904fef, 32'h00000000} /* (9, 16, 17) {real, imag} */,
  {32'h3f952fb6, 32'h00000000} /* (9, 16, 16) {real, imag} */,
  {32'h3f80b592, 32'h00000000} /* (9, 16, 15) {real, imag} */,
  {32'h3f346efe, 32'h00000000} /* (9, 16, 14) {real, imag} */,
  {32'h3f308501, 32'h00000000} /* (9, 16, 13) {real, imag} */,
  {32'h3f2195c5, 32'h00000000} /* (9, 16, 12) {real, imag} */,
  {32'h3e4b6702, 32'h00000000} /* (9, 16, 11) {real, imag} */,
  {32'hbf212217, 32'h00000000} /* (9, 16, 10) {real, imag} */,
  {32'hbf56aeae, 32'h00000000} /* (9, 16, 9) {real, imag} */,
  {32'hbf88d8bb, 32'h00000000} /* (9, 16, 8) {real, imag} */,
  {32'hbf111133, 32'h00000000} /* (9, 16, 7) {real, imag} */,
  {32'hbf185e66, 32'h00000000} /* (9, 16, 6) {real, imag} */,
  {32'hbf1f4acc, 32'h00000000} /* (9, 16, 5) {real, imag} */,
  {32'hbf3b2567, 32'h00000000} /* (9, 16, 4) {real, imag} */,
  {32'hbf9ecff0, 32'h00000000} /* (9, 16, 3) {real, imag} */,
  {32'hbf9ab1a6, 32'h00000000} /* (9, 16, 2) {real, imag} */,
  {32'hbf1608e2, 32'h00000000} /* (9, 16, 1) {real, imag} */,
  {32'hbda4098a, 32'h00000000} /* (9, 16, 0) {real, imag} */,
  {32'hbf10e219, 32'h00000000} /* (9, 15, 31) {real, imag} */,
  {32'hbfb2711c, 32'h00000000} /* (9, 15, 30) {real, imag} */,
  {32'hbf63aaf5, 32'h00000000} /* (9, 15, 29) {real, imag} */,
  {32'hbf4ddd71, 32'h00000000} /* (9, 15, 28) {real, imag} */,
  {32'hbf89b42c, 32'h00000000} /* (9, 15, 27) {real, imag} */,
  {32'hbf698b75, 32'h00000000} /* (9, 15, 26) {real, imag} */,
  {32'hbf794202, 32'h00000000} /* (9, 15, 25) {real, imag} */,
  {32'hbf8085f1, 32'h00000000} /* (9, 15, 24) {real, imag} */,
  {32'hbf6614f5, 32'h00000000} /* (9, 15, 23) {real, imag} */,
  {32'hbf393465, 32'h00000000} /* (9, 15, 22) {real, imag} */,
  {32'h3e117bb9, 32'h00000000} /* (9, 15, 21) {real, imag} */,
  {32'h3f4cd35b, 32'h00000000} /* (9, 15, 20) {real, imag} */,
  {32'h3f0f5f83, 32'h00000000} /* (9, 15, 19) {real, imag} */,
  {32'h3f8f00c8, 32'h00000000} /* (9, 15, 18) {real, imag} */,
  {32'h3f956106, 32'h00000000} /* (9, 15, 17) {real, imag} */,
  {32'h3f9edd7f, 32'h00000000} /* (9, 15, 16) {real, imag} */,
  {32'h3f5e479d, 32'h00000000} /* (9, 15, 15) {real, imag} */,
  {32'h3f2cca2b, 32'h00000000} /* (9, 15, 14) {real, imag} */,
  {32'h3f83691a, 32'h00000000} /* (9, 15, 13) {real, imag} */,
  {32'h3f95b1f3, 32'h00000000} /* (9, 15, 12) {real, imag} */,
  {32'h3f19823e, 32'h00000000} /* (9, 15, 11) {real, imag} */,
  {32'hbedd7bba, 32'h00000000} /* (9, 15, 10) {real, imag} */,
  {32'hbf266bfa, 32'h00000000} /* (9, 15, 9) {real, imag} */,
  {32'hbf84aa71, 32'h00000000} /* (9, 15, 8) {real, imag} */,
  {32'hbf791a52, 32'h00000000} /* (9, 15, 7) {real, imag} */,
  {32'hbf34f1e5, 32'h00000000} /* (9, 15, 6) {real, imag} */,
  {32'hbef4d2c4, 32'h00000000} /* (9, 15, 5) {real, imag} */,
  {32'hbf4b9e9a, 32'h00000000} /* (9, 15, 4) {real, imag} */,
  {32'hbf8070b9, 32'h00000000} /* (9, 15, 3) {real, imag} */,
  {32'hbf863817, 32'h00000000} /* (9, 15, 2) {real, imag} */,
  {32'hbf3ce95f, 32'h00000000} /* (9, 15, 1) {real, imag} */,
  {32'hbedadc76, 32'h00000000} /* (9, 15, 0) {real, imag} */,
  {32'hbf0d65d6, 32'h00000000} /* (9, 14, 31) {real, imag} */,
  {32'hbf832e9f, 32'h00000000} /* (9, 14, 30) {real, imag} */,
  {32'hbefa3605, 32'h00000000} /* (9, 14, 29) {real, imag} */,
  {32'hbf4ed1f8, 32'h00000000} /* (9, 14, 28) {real, imag} */,
  {32'hbfc19711, 32'h00000000} /* (9, 14, 27) {real, imag} */,
  {32'hbf980dd9, 32'h00000000} /* (9, 14, 26) {real, imag} */,
  {32'hbf9d9cc8, 32'h00000000} /* (9, 14, 25) {real, imag} */,
  {32'hbf341568, 32'h00000000} /* (9, 14, 24) {real, imag} */,
  {32'hbf254bdd, 32'h00000000} /* (9, 14, 23) {real, imag} */,
  {32'hbf3de941, 32'h00000000} /* (9, 14, 22) {real, imag} */,
  {32'hbe9b5783, 32'h00000000} /* (9, 14, 21) {real, imag} */,
  {32'h3f17335b, 32'h00000000} /* (9, 14, 20) {real, imag} */,
  {32'h3e80ef0b, 32'h00000000} /* (9, 14, 19) {real, imag} */,
  {32'h3f0b30d2, 32'h00000000} /* (9, 14, 18) {real, imag} */,
  {32'h3f2b8d90, 32'h00000000} /* (9, 14, 17) {real, imag} */,
  {32'h3f0f8217, 32'h00000000} /* (9, 14, 16) {real, imag} */,
  {32'h3eed3e61, 32'h00000000} /* (9, 14, 15) {real, imag} */,
  {32'h3f6aa6a9, 32'h00000000} /* (9, 14, 14) {real, imag} */,
  {32'h3fc5c5f3, 32'h00000000} /* (9, 14, 13) {real, imag} */,
  {32'h3f90a1cc, 32'h00000000} /* (9, 14, 12) {real, imag} */,
  {32'h3f50bae4, 32'h00000000} /* (9, 14, 11) {real, imag} */,
  {32'hbe0b649e, 32'h00000000} /* (9, 14, 10) {real, imag} */,
  {32'hbf850643, 32'h00000000} /* (9, 14, 9) {real, imag} */,
  {32'hbf7ceeea, 32'h00000000} /* (9, 14, 8) {real, imag} */,
  {32'hbf3e4cd1, 32'h00000000} /* (9, 14, 7) {real, imag} */,
  {32'hbee73338, 32'h00000000} /* (9, 14, 6) {real, imag} */,
  {32'hbef34d27, 32'h00000000} /* (9, 14, 5) {real, imag} */,
  {32'hbee25587, 32'h00000000} /* (9, 14, 4) {real, imag} */,
  {32'hbf02e974, 32'h00000000} /* (9, 14, 3) {real, imag} */,
  {32'hbf21cb99, 32'h00000000} /* (9, 14, 2) {real, imag} */,
  {32'hbf42e1d6, 32'h00000000} /* (9, 14, 1) {real, imag} */,
  {32'hbf00cdda, 32'h00000000} /* (9, 14, 0) {real, imag} */,
  {32'hbf037b89, 32'h00000000} /* (9, 13, 31) {real, imag} */,
  {32'hbf4121da, 32'h00000000} /* (9, 13, 30) {real, imag} */,
  {32'hbf2d0b40, 32'h00000000} /* (9, 13, 29) {real, imag} */,
  {32'hbf6d5f16, 32'h00000000} /* (9, 13, 28) {real, imag} */,
  {32'hbf3d4c1a, 32'h00000000} /* (9, 13, 27) {real, imag} */,
  {32'hbf33b1c8, 32'h00000000} /* (9, 13, 26) {real, imag} */,
  {32'hbf3f1371, 32'h00000000} /* (9, 13, 25) {real, imag} */,
  {32'hbf3b49f0, 32'h00000000} /* (9, 13, 24) {real, imag} */,
  {32'hbf4e9cda, 32'h00000000} /* (9, 13, 23) {real, imag} */,
  {32'hbf3fdde5, 32'h00000000} /* (9, 13, 22) {real, imag} */,
  {32'hbdb54e7a, 32'h00000000} /* (9, 13, 21) {real, imag} */,
  {32'h3f603dc6, 32'h00000000} /* (9, 13, 20) {real, imag} */,
  {32'h3f121f77, 32'h00000000} /* (9, 13, 19) {real, imag} */,
  {32'h3f408f49, 32'h00000000} /* (9, 13, 18) {real, imag} */,
  {32'h3f1179a2, 32'h00000000} /* (9, 13, 17) {real, imag} */,
  {32'h3e9e6103, 32'h00000000} /* (9, 13, 16) {real, imag} */,
  {32'h3eab797e, 32'h00000000} /* (9, 13, 15) {real, imag} */,
  {32'h3f0e9405, 32'h00000000} /* (9, 13, 14) {real, imag} */,
  {32'h3f969672, 32'h00000000} /* (9, 13, 13) {real, imag} */,
  {32'h3f81bfa1, 32'h00000000} /* (9, 13, 12) {real, imag} */,
  {32'h3f37fa42, 32'h00000000} /* (9, 13, 11) {real, imag} */,
  {32'hbf114756, 32'h00000000} /* (9, 13, 10) {real, imag} */,
  {32'hbfb2176a, 32'h00000000} /* (9, 13, 9) {real, imag} */,
  {32'hbf771802, 32'h00000000} /* (9, 13, 8) {real, imag} */,
  {32'hbf835192, 32'h00000000} /* (9, 13, 7) {real, imag} */,
  {32'hbf1ff62a, 32'h00000000} /* (9, 13, 6) {real, imag} */,
  {32'hbf3607b6, 32'h00000000} /* (9, 13, 5) {real, imag} */,
  {32'hbf2638cf, 32'h00000000} /* (9, 13, 4) {real, imag} */,
  {32'hbf516216, 32'h00000000} /* (9, 13, 3) {real, imag} */,
  {32'hbedd77c3, 32'h00000000} /* (9, 13, 2) {real, imag} */,
  {32'hbf41c88d, 32'h00000000} /* (9, 13, 1) {real, imag} */,
  {32'hbf509e4e, 32'h00000000} /* (9, 13, 0) {real, imag} */,
  {32'hbef960da, 32'h00000000} /* (9, 12, 31) {real, imag} */,
  {32'hbf89a49c, 32'h00000000} /* (9, 12, 30) {real, imag} */,
  {32'hbf7da554, 32'h00000000} /* (9, 12, 29) {real, imag} */,
  {32'hbf78d46f, 32'h00000000} /* (9, 12, 28) {real, imag} */,
  {32'hbf5f2e03, 32'h00000000} /* (9, 12, 27) {real, imag} */,
  {32'hbf44252f, 32'h00000000} /* (9, 12, 26) {real, imag} */,
  {32'hbf2c5d00, 32'h00000000} /* (9, 12, 25) {real, imag} */,
  {32'hbf6349d7, 32'h00000000} /* (9, 12, 24) {real, imag} */,
  {32'hbf3c37e7, 32'h00000000} /* (9, 12, 23) {real, imag} */,
  {32'hbf0a1310, 32'h00000000} /* (9, 12, 22) {real, imag} */,
  {32'hbac855df, 32'h00000000} /* (9, 12, 21) {real, imag} */,
  {32'h3f6fa2b4, 32'h00000000} /* (9, 12, 20) {real, imag} */,
  {32'h3f76e2b9, 32'h00000000} /* (9, 12, 19) {real, imag} */,
  {32'h3ed003b7, 32'h00000000} /* (9, 12, 18) {real, imag} */,
  {32'h3f14a451, 32'h00000000} /* (9, 12, 17) {real, imag} */,
  {32'h3f51b873, 32'h00000000} /* (9, 12, 16) {real, imag} */,
  {32'h3f2d7ae9, 32'h00000000} /* (9, 12, 15) {real, imag} */,
  {32'h3f2df9d3, 32'h00000000} /* (9, 12, 14) {real, imag} */,
  {32'h3eff6c92, 32'h00000000} /* (9, 12, 13) {real, imag} */,
  {32'h3f3b3198, 32'h00000000} /* (9, 12, 12) {real, imag} */,
  {32'h3e6853f0, 32'h00000000} /* (9, 12, 11) {real, imag} */,
  {32'hbf5e2bc8, 32'h00000000} /* (9, 12, 10) {real, imag} */,
  {32'hbfaf9104, 32'h00000000} /* (9, 12, 9) {real, imag} */,
  {32'hbf3575a6, 32'h00000000} /* (9, 12, 8) {real, imag} */,
  {32'hbf8348ea, 32'h00000000} /* (9, 12, 7) {real, imag} */,
  {32'hbf80eb02, 32'h00000000} /* (9, 12, 6) {real, imag} */,
  {32'hbf2961ac, 32'h00000000} /* (9, 12, 5) {real, imag} */,
  {32'hbf396e2c, 32'h00000000} /* (9, 12, 4) {real, imag} */,
  {32'hbf3a339a, 32'h00000000} /* (9, 12, 3) {real, imag} */,
  {32'hbed14c47, 32'h00000000} /* (9, 12, 2) {real, imag} */,
  {32'hbf048d9d, 32'h00000000} /* (9, 12, 1) {real, imag} */,
  {32'hbf0d4cb4, 32'h00000000} /* (9, 12, 0) {real, imag} */,
  {32'h3b12ba91, 32'h00000000} /* (9, 11, 31) {real, imag} */,
  {32'hbea4f8de, 32'h00000000} /* (9, 11, 30) {real, imag} */,
  {32'hbe83f7c7, 32'h00000000} /* (9, 11, 29) {real, imag} */,
  {32'hbf17b508, 32'h00000000} /* (9, 11, 28) {real, imag} */,
  {32'hbf615b4f, 32'h00000000} /* (9, 11, 27) {real, imag} */,
  {32'hbefe2f4b, 32'h00000000} /* (9, 11, 26) {real, imag} */,
  {32'hbf01f811, 32'h00000000} /* (9, 11, 25) {real, imag} */,
  {32'hbf65b89e, 32'h00000000} /* (9, 11, 24) {real, imag} */,
  {32'hbeea27e8, 32'h00000000} /* (9, 11, 23) {real, imag} */,
  {32'hbe3b58ea, 32'h00000000} /* (9, 11, 22) {real, imag} */,
  {32'hbe8e4b8a, 32'h00000000} /* (9, 11, 21) {real, imag} */,
  {32'h3ed4fe4b, 32'h00000000} /* (9, 11, 20) {real, imag} */,
  {32'h3eea058f, 32'h00000000} /* (9, 11, 19) {real, imag} */,
  {32'h3da28d2d, 32'h00000000} /* (9, 11, 18) {real, imag} */,
  {32'h3ea62136, 32'h00000000} /* (9, 11, 17) {real, imag} */,
  {32'h3f19b40d, 32'h00000000} /* (9, 11, 16) {real, imag} */,
  {32'h3f282efa, 32'h00000000} /* (9, 11, 15) {real, imag} */,
  {32'h3f48f7f5, 32'h00000000} /* (9, 11, 14) {real, imag} */,
  {32'h3f2da291, 32'h00000000} /* (9, 11, 13) {real, imag} */,
  {32'h3f021883, 32'h00000000} /* (9, 11, 12) {real, imag} */,
  {32'h3d51672c, 32'h00000000} /* (9, 11, 11) {real, imag} */,
  {32'hbf0b7726, 32'h00000000} /* (9, 11, 10) {real, imag} */,
  {32'hbebb2d09, 32'h00000000} /* (9, 11, 9) {real, imag} */,
  {32'hbee52ed4, 32'h00000000} /* (9, 11, 8) {real, imag} */,
  {32'hbf0c1b3c, 32'h00000000} /* (9, 11, 7) {real, imag} */,
  {32'hbee2673f, 32'h00000000} /* (9, 11, 6) {real, imag} */,
  {32'h3b968e27, 32'h00000000} /* (9, 11, 5) {real, imag} */,
  {32'hbde3331a, 32'h00000000} /* (9, 11, 4) {real, imag} */,
  {32'hbe3a9238, 32'h00000000} /* (9, 11, 3) {real, imag} */,
  {32'hbf29c5d5, 32'h00000000} /* (9, 11, 2) {real, imag} */,
  {32'hbf43fefc, 32'h00000000} /* (9, 11, 1) {real, imag} */,
  {32'hbd6675c7, 32'h00000000} /* (9, 11, 0) {real, imag} */,
  {32'h3ebc6713, 32'h00000000} /* (9, 10, 31) {real, imag} */,
  {32'h3eeb8f6d, 32'h00000000} /* (9, 10, 30) {real, imag} */,
  {32'h3f815214, 32'h00000000} /* (9, 10, 29) {real, imag} */,
  {32'h3f1c6dbb, 32'h00000000} /* (9, 10, 28) {real, imag} */,
  {32'h3f0deafa, 32'h00000000} /* (9, 10, 27) {real, imag} */,
  {32'h3e95f679, 32'h00000000} /* (9, 10, 26) {real, imag} */,
  {32'h3e6d1c61, 32'h00000000} /* (9, 10, 25) {real, imag} */,
  {32'h3dabd286, 32'h00000000} /* (9, 10, 24) {real, imag} */,
  {32'h3f0856fc, 32'h00000000} /* (9, 10, 23) {real, imag} */,
  {32'h3f5fd778, 32'h00000000} /* (9, 10, 22) {real, imag} */,
  {32'h3e9a3ec3, 32'h00000000} /* (9, 10, 21) {real, imag} */,
  {32'hbda83e34, 32'h00000000} /* (9, 10, 20) {real, imag} */,
  {32'hbf27947b, 32'h00000000} /* (9, 10, 19) {real, imag} */,
  {32'hbf8afaba, 32'h00000000} /* (9, 10, 18) {real, imag} */,
  {32'hbea2f777, 32'h00000000} /* (9, 10, 17) {real, imag} */,
  {32'hbf08d395, 32'h00000000} /* (9, 10, 16) {real, imag} */,
  {32'hbeee0519, 32'h00000000} /* (9, 10, 15) {real, imag} */,
  {32'hbedc82ab, 32'h00000000} /* (9, 10, 14) {real, imag} */,
  {32'hbeaf2f39, 32'h00000000} /* (9, 10, 13) {real, imag} */,
  {32'hbf175174, 32'h00000000} /* (9, 10, 12) {real, imag} */,
  {32'hbeb96304, 32'h00000000} /* (9, 10, 11) {real, imag} */,
  {32'hbe2ed651, 32'h00000000} /* (9, 10, 10) {real, imag} */,
  {32'h3e0ee5e1, 32'h00000000} /* (9, 10, 9) {real, imag} */,
  {32'hbcef596d, 32'h00000000} /* (9, 10, 8) {real, imag} */,
  {32'h3f03e58e, 32'h00000000} /* (9, 10, 7) {real, imag} */,
  {32'h3f52caca, 32'h00000000} /* (9, 10, 6) {real, imag} */,
  {32'h3f977ead, 32'h00000000} /* (9, 10, 5) {real, imag} */,
  {32'h3f5ac969, 32'h00000000} /* (9, 10, 4) {real, imag} */,
  {32'h3ec60ca9, 32'h00000000} /* (9, 10, 3) {real, imag} */,
  {32'hbe2d24e5, 32'h00000000} /* (9, 10, 2) {real, imag} */,
  {32'hbde97646, 32'h00000000} /* (9, 10, 1) {real, imag} */,
  {32'h3ece9513, 32'h00000000} /* (9, 10, 0) {real, imag} */,
  {32'h3ef1992f, 32'h00000000} /* (9, 9, 31) {real, imag} */,
  {32'h3f3fa17f, 32'h00000000} /* (9, 9, 30) {real, imag} */,
  {32'h3faf9e3e, 32'h00000000} /* (9, 9, 29) {real, imag} */,
  {32'h3fa74bcb, 32'h00000000} /* (9, 9, 28) {real, imag} */,
  {32'h3f9ef5da, 32'h00000000} /* (9, 9, 27) {real, imag} */,
  {32'h3f1a03a0, 32'h00000000} /* (9, 9, 26) {real, imag} */,
  {32'h3f2197e5, 32'h00000000} /* (9, 9, 25) {real, imag} */,
  {32'h3f588519, 32'h00000000} /* (9, 9, 24) {real, imag} */,
  {32'h3f634fa1, 32'h00000000} /* (9, 9, 23) {real, imag} */,
  {32'h3f35a9e9, 32'h00000000} /* (9, 9, 22) {real, imag} */,
  {32'h3ede826d, 32'h00000000} /* (9, 9, 21) {real, imag} */,
  {32'hbd99926c, 32'h00000000} /* (9, 9, 20) {real, imag} */,
  {32'hbf2cd7b1, 32'h00000000} /* (9, 9, 19) {real, imag} */,
  {32'hbfbd16e5, 32'h00000000} /* (9, 9, 18) {real, imag} */,
  {32'hbf8c69f3, 32'h00000000} /* (9, 9, 17) {real, imag} */,
  {32'hbf8bc202, 32'h00000000} /* (9, 9, 16) {real, imag} */,
  {32'hbf85457d, 32'h00000000} /* (9, 9, 15) {real, imag} */,
  {32'hbf8008f4, 32'h00000000} /* (9, 9, 14) {real, imag} */,
  {32'hbfa5af8b, 32'h00000000} /* (9, 9, 13) {real, imag} */,
  {32'hbfa1e714, 32'h00000000} /* (9, 9, 12) {real, imag} */,
  {32'hbf304fbf, 32'h00000000} /* (9, 9, 11) {real, imag} */,
  {32'hbc1a3f90, 32'h00000000} /* (9, 9, 10) {real, imag} */,
  {32'h3e148f03, 32'h00000000} /* (9, 9, 9) {real, imag} */,
  {32'h3e021ea3, 32'h00000000} /* (9, 9, 8) {real, imag} */,
  {32'h3f10ac6a, 32'h00000000} /* (9, 9, 7) {real, imag} */,
  {32'h3f64edf4, 32'h00000000} /* (9, 9, 6) {real, imag} */,
  {32'h3f903658, 32'h00000000} /* (9, 9, 5) {real, imag} */,
  {32'h3f4d1657, 32'h00000000} /* (9, 9, 4) {real, imag} */,
  {32'h3f3e22f7, 32'h00000000} /* (9, 9, 3) {real, imag} */,
  {32'h3ec48c65, 32'h00000000} /* (9, 9, 2) {real, imag} */,
  {32'h3e6e7f3c, 32'h00000000} /* (9, 9, 1) {real, imag} */,
  {32'h3e80704d, 32'h00000000} /* (9, 9, 0) {real, imag} */,
  {32'h3ed73105, 32'h00000000} /* (9, 8, 31) {real, imag} */,
  {32'h3f137b5d, 32'h00000000} /* (9, 8, 30) {real, imag} */,
  {32'h3fb7649f, 32'h00000000} /* (9, 8, 29) {real, imag} */,
  {32'h3f8e353c, 32'h00000000} /* (9, 8, 28) {real, imag} */,
  {32'h3f9f246f, 32'h00000000} /* (9, 8, 27) {real, imag} */,
  {32'h3f70cda3, 32'h00000000} /* (9, 8, 26) {real, imag} */,
  {32'h3f301c58, 32'h00000000} /* (9, 8, 25) {real, imag} */,
  {32'h3f8a635c, 32'h00000000} /* (9, 8, 24) {real, imag} */,
  {32'h3f9a27ca, 32'h00000000} /* (9, 8, 23) {real, imag} */,
  {32'h3f67d9ab, 32'h00000000} /* (9, 8, 22) {real, imag} */,
  {32'h3e55e05c, 32'h00000000} /* (9, 8, 21) {real, imag} */,
  {32'hbeb8c970, 32'h00000000} /* (9, 8, 20) {real, imag} */,
  {32'hbe892378, 32'h00000000} /* (9, 8, 19) {real, imag} */,
  {32'hbf56bcfb, 32'h00000000} /* (9, 8, 18) {real, imag} */,
  {32'hbf8f466b, 32'h00000000} /* (9, 8, 17) {real, imag} */,
  {32'hbf7f456e, 32'h00000000} /* (9, 8, 16) {real, imag} */,
  {32'hbf861e08, 32'h00000000} /* (9, 8, 15) {real, imag} */,
  {32'hbf827476, 32'h00000000} /* (9, 8, 14) {real, imag} */,
  {32'hbf86eee9, 32'h00000000} /* (9, 8, 13) {real, imag} */,
  {32'hbf844d67, 32'h00000000} /* (9, 8, 12) {real, imag} */,
  {32'hbf44a01e, 32'h00000000} /* (9, 8, 11) {real, imag} */,
  {32'h3e9a2cee, 32'h00000000} /* (9, 8, 10) {real, imag} */,
  {32'h3f1ba464, 32'h00000000} /* (9, 8, 9) {real, imag} */,
  {32'h3f4ef710, 32'h00000000} /* (9, 8, 8) {real, imag} */,
  {32'h3f9df3f8, 32'h00000000} /* (9, 8, 7) {real, imag} */,
  {32'h3fa74839, 32'h00000000} /* (9, 8, 6) {real, imag} */,
  {32'h3f605c72, 32'h00000000} /* (9, 8, 5) {real, imag} */,
  {32'h3f748337, 32'h00000000} /* (9, 8, 4) {real, imag} */,
  {32'h3f1bf957, 32'h00000000} /* (9, 8, 3) {real, imag} */,
  {32'h3f088d24, 32'h00000000} /* (9, 8, 2) {real, imag} */,
  {32'h3eefda84, 32'h00000000} /* (9, 8, 1) {real, imag} */,
  {32'h3e266c58, 32'h00000000} /* (9, 8, 0) {real, imag} */,
  {32'h3e27bba9, 32'h00000000} /* (9, 7, 31) {real, imag} */,
  {32'h3ea3f70d, 32'h00000000} /* (9, 7, 30) {real, imag} */,
  {32'h3fad3a67, 32'h00000000} /* (9, 7, 29) {real, imag} */,
  {32'h3f911a5a, 32'h00000000} /* (9, 7, 28) {real, imag} */,
  {32'h3f41ba2c, 32'h00000000} /* (9, 7, 27) {real, imag} */,
  {32'h3f16b3e6, 32'h00000000} /* (9, 7, 26) {real, imag} */,
  {32'h3ed9a069, 32'h00000000} /* (9, 7, 25) {real, imag} */,
  {32'h3f4a7b65, 32'h00000000} /* (9, 7, 24) {real, imag} */,
  {32'h3f924db3, 32'h00000000} /* (9, 7, 23) {real, imag} */,
  {32'h3f94a104, 32'h00000000} /* (9, 7, 22) {real, imag} */,
  {32'h3ee8ab9b, 32'h00000000} /* (9, 7, 21) {real, imag} */,
  {32'hbea20570, 32'h00000000} /* (9, 7, 20) {real, imag} */,
  {32'hbeeda6c7, 32'h00000000} /* (9, 7, 19) {real, imag} */,
  {32'hbf4affef, 32'h00000000} /* (9, 7, 18) {real, imag} */,
  {32'hbf8dc048, 32'h00000000} /* (9, 7, 17) {real, imag} */,
  {32'hbf5d18c9, 32'h00000000} /* (9, 7, 16) {real, imag} */,
  {32'hbf80e489, 32'h00000000} /* (9, 7, 15) {real, imag} */,
  {32'hbf7a96a0, 32'h00000000} /* (9, 7, 14) {real, imag} */,
  {32'hbf92f4c8, 32'h00000000} /* (9, 7, 13) {real, imag} */,
  {32'hbfa8f4ea, 32'h00000000} /* (9, 7, 12) {real, imag} */,
  {32'hbf7b0035, 32'h00000000} /* (9, 7, 11) {real, imag} */,
  {32'h3ebb4f3e, 32'h00000000} /* (9, 7, 10) {real, imag} */,
  {32'h3f857f49, 32'h00000000} /* (9, 7, 9) {real, imag} */,
  {32'h3f96f573, 32'h00000000} /* (9, 7, 8) {real, imag} */,
  {32'h3fa57b2c, 32'h00000000} /* (9, 7, 7) {real, imag} */,
  {32'h3f8063ae, 32'h00000000} /* (9, 7, 6) {real, imag} */,
  {32'h3f860034, 32'h00000000} /* (9, 7, 5) {real, imag} */,
  {32'h3f9a95fc, 32'h00000000} /* (9, 7, 4) {real, imag} */,
  {32'h3f40f02a, 32'h00000000} /* (9, 7, 3) {real, imag} */,
  {32'h3f338b2b, 32'h00000000} /* (9, 7, 2) {real, imag} */,
  {32'h3f6e7df8, 32'h00000000} /* (9, 7, 1) {real, imag} */,
  {32'h3edef1ad, 32'h00000000} /* (9, 7, 0) {real, imag} */,
  {32'h3e49d854, 32'h00000000} /* (9, 6, 31) {real, imag} */,
  {32'h3e0cbc54, 32'h00000000} /* (9, 6, 30) {real, imag} */,
  {32'h3f505706, 32'h00000000} /* (9, 6, 29) {real, imag} */,
  {32'h3f812e4f, 32'h00000000} /* (9, 6, 28) {real, imag} */,
  {32'h3ef70e42, 32'h00000000} /* (9, 6, 27) {real, imag} */,
  {32'h3edb7c2c, 32'h00000000} /* (9, 6, 26) {real, imag} */,
  {32'h3ed2d0a2, 32'h00000000} /* (9, 6, 25) {real, imag} */,
  {32'h3f897563, 32'h00000000} /* (9, 6, 24) {real, imag} */,
  {32'h3fc4abdc, 32'h00000000} /* (9, 6, 23) {real, imag} */,
  {32'h3f8dce91, 32'h00000000} /* (9, 6, 22) {real, imag} */,
  {32'h3f3114be, 32'h00000000} /* (9, 6, 21) {real, imag} */,
  {32'h3d287a00, 32'h00000000} /* (9, 6, 20) {real, imag} */,
  {32'hbef88ae9, 32'h00000000} /* (9, 6, 19) {real, imag} */,
  {32'hbf52a245, 32'h00000000} /* (9, 6, 18) {real, imag} */,
  {32'hbf145d8b, 32'h00000000} /* (9, 6, 17) {real, imag} */,
  {32'hbf5542b5, 32'h00000000} /* (9, 6, 16) {real, imag} */,
  {32'hbf92600d, 32'h00000000} /* (9, 6, 15) {real, imag} */,
  {32'hbf83577c, 32'h00000000} /* (9, 6, 14) {real, imag} */,
  {32'hbf9a92f8, 32'h00000000} /* (9, 6, 13) {real, imag} */,
  {32'hbf9dde41, 32'h00000000} /* (9, 6, 12) {real, imag} */,
  {32'hbf612d76, 32'h00000000} /* (9, 6, 11) {real, imag} */,
  {32'h3e2efaf0, 32'h00000000} /* (9, 6, 10) {real, imag} */,
  {32'h3ec5607c, 32'h00000000} /* (9, 6, 9) {real, imag} */,
  {32'h3ea302ec, 32'h00000000} /* (9, 6, 8) {real, imag} */,
  {32'h3f456f05, 32'h00000000} /* (9, 6, 7) {real, imag} */,
  {32'h3f8ad308, 32'h00000000} /* (9, 6, 6) {real, imag} */,
  {32'h3feaf4eb, 32'h00000000} /* (9, 6, 5) {real, imag} */,
  {32'h3f7a4933, 32'h00000000} /* (9, 6, 4) {real, imag} */,
  {32'h3f3c68f0, 32'h00000000} /* (9, 6, 3) {real, imag} */,
  {32'h3f3b4ec0, 32'h00000000} /* (9, 6, 2) {real, imag} */,
  {32'h3f7a82e0, 32'h00000000} /* (9, 6, 1) {real, imag} */,
  {32'h3f165c76, 32'h00000000} /* (9, 6, 0) {real, imag} */,
  {32'h3eda5698, 32'h00000000} /* (9, 5, 31) {real, imag} */,
  {32'h3e9bccaf, 32'h00000000} /* (9, 5, 30) {real, imag} */,
  {32'h3f1b0f72, 32'h00000000} /* (9, 5, 29) {real, imag} */,
  {32'h3f739d6d, 32'h00000000} /* (9, 5, 28) {real, imag} */,
  {32'h3f7225ec, 32'h00000000} /* (9, 5, 27) {real, imag} */,
  {32'h3f94b0ae, 32'h00000000} /* (9, 5, 26) {real, imag} */,
  {32'h3f2ec59f, 32'h00000000} /* (9, 5, 25) {real, imag} */,
  {32'h3f2c3ec1, 32'h00000000} /* (9, 5, 24) {real, imag} */,
  {32'h3fac0786, 32'h00000000} /* (9, 5, 23) {real, imag} */,
  {32'h3fb3d305, 32'h00000000} /* (9, 5, 22) {real, imag} */,
  {32'h3f86c1b0, 32'h00000000} /* (9, 5, 21) {real, imag} */,
  {32'h3f983fd0, 32'h00000000} /* (9, 5, 20) {real, imag} */,
  {32'h3efd42a2, 32'h00000000} /* (9, 5, 19) {real, imag} */,
  {32'h3cbc93ae, 32'h00000000} /* (9, 5, 18) {real, imag} */,
  {32'h3f45ad7f, 32'h00000000} /* (9, 5, 17) {real, imag} */,
  {32'h3d5a0912, 32'h00000000} /* (9, 5, 16) {real, imag} */,
  {32'hbf57a460, 32'h00000000} /* (9, 5, 15) {real, imag} */,
  {32'hbf477f80, 32'h00000000} /* (9, 5, 14) {real, imag} */,
  {32'hbf34c63e, 32'h00000000} /* (9, 5, 13) {real, imag} */,
  {32'hbfa7809a, 32'h00000000} /* (9, 5, 12) {real, imag} */,
  {32'hbfb7af92, 32'h00000000} /* (9, 5, 11) {real, imag} */,
  {32'hbecca7fc, 32'h00000000} /* (9, 5, 10) {real, imag} */,
  {32'hbec5a954, 32'h00000000} /* (9, 5, 9) {real, imag} */,
  {32'hbeafb66c, 32'h00000000} /* (9, 5, 8) {real, imag} */,
  {32'h3dc7d2ff, 32'h00000000} /* (9, 5, 7) {real, imag} */,
  {32'h3f1d544c, 32'h00000000} /* (9, 5, 6) {real, imag} */,
  {32'h3fb0e486, 32'h00000000} /* (9, 5, 5) {real, imag} */,
  {32'h3f19d6a1, 32'h00000000} /* (9, 5, 4) {real, imag} */,
  {32'h3f55e5da, 32'h00000000} /* (9, 5, 3) {real, imag} */,
  {32'h3f689319, 32'h00000000} /* (9, 5, 2) {real, imag} */,
  {32'h3fac78ea, 32'h00000000} /* (9, 5, 1) {real, imag} */,
  {32'h3f856531, 32'h00000000} /* (9, 5, 0) {real, imag} */,
  {32'h3f25b24f, 32'h00000000} /* (9, 4, 31) {real, imag} */,
  {32'h3f342d03, 32'h00000000} /* (9, 4, 30) {real, imag} */,
  {32'h3f56d95d, 32'h00000000} /* (9, 4, 29) {real, imag} */,
  {32'h3f83b337, 32'h00000000} /* (9, 4, 28) {real, imag} */,
  {32'h3fdf5e3a, 32'h00000000} /* (9, 4, 27) {real, imag} */,
  {32'h3fac224e, 32'h00000000} /* (9, 4, 26) {real, imag} */,
  {32'h3f1ada5b, 32'h00000000} /* (9, 4, 25) {real, imag} */,
  {32'h3f118b4a, 32'h00000000} /* (9, 4, 24) {real, imag} */,
  {32'h3f5a5921, 32'h00000000} /* (9, 4, 23) {real, imag} */,
  {32'h3f981ab5, 32'h00000000} /* (9, 4, 22) {real, imag} */,
  {32'h3f64fc0e, 32'h00000000} /* (9, 4, 21) {real, imag} */,
  {32'h3fa18029, 32'h00000000} /* (9, 4, 20) {real, imag} */,
  {32'h3f5a14ef, 32'h00000000} /* (9, 4, 19) {real, imag} */,
  {32'h3efd9bb9, 32'h00000000} /* (9, 4, 18) {real, imag} */,
  {32'h3f423044, 32'h00000000} /* (9, 4, 17) {real, imag} */,
  {32'h3ddc8312, 32'h00000000} /* (9, 4, 16) {real, imag} */,
  {32'hbf5c8364, 32'h00000000} /* (9, 4, 15) {real, imag} */,
  {32'hbea4e99d, 32'h00000000} /* (9, 4, 14) {real, imag} */,
  {32'hbf14438e, 32'h00000000} /* (9, 4, 13) {real, imag} */,
  {32'hbfd4f596, 32'h00000000} /* (9, 4, 12) {real, imag} */,
  {32'hbfc71136, 32'h00000000} /* (9, 4, 11) {real, imag} */,
  {32'hbf05dd70, 32'h00000000} /* (9, 4, 10) {real, imag} */,
  {32'hbea258d1, 32'h00000000} /* (9, 4, 9) {real, imag} */,
  {32'hbeec4375, 32'h00000000} /* (9, 4, 8) {real, imag} */,
  {32'hbef3e2ba, 32'h00000000} /* (9, 4, 7) {real, imag} */,
  {32'hbf29ba49, 32'h00000000} /* (9, 4, 6) {real, imag} */,
  {32'h3ebef204, 32'h00000000} /* (9, 4, 5) {real, imag} */,
  {32'h3f492250, 32'h00000000} /* (9, 4, 4) {real, imag} */,
  {32'h3f62cd87, 32'h00000000} /* (9, 4, 3) {real, imag} */,
  {32'h3f5e9329, 32'h00000000} /* (9, 4, 2) {real, imag} */,
  {32'h3f8bd82b, 32'h00000000} /* (9, 4, 1) {real, imag} */,
  {32'h3f802653, 32'h00000000} /* (9, 4, 0) {real, imag} */,
  {32'h3ec41692, 32'h00000000} /* (9, 3, 31) {real, imag} */,
  {32'h3f6c20b0, 32'h00000000} /* (9, 3, 30) {real, imag} */,
  {32'h3f871905, 32'h00000000} /* (9, 3, 29) {real, imag} */,
  {32'h3f576280, 32'h00000000} /* (9, 3, 28) {real, imag} */,
  {32'h3f885aa3, 32'h00000000} /* (9, 3, 27) {real, imag} */,
  {32'h3f8782a3, 32'h00000000} /* (9, 3, 26) {real, imag} */,
  {32'h3f94de26, 32'h00000000} /* (9, 3, 25) {real, imag} */,
  {32'h3fa55fec, 32'h00000000} /* (9, 3, 24) {real, imag} */,
  {32'h3f49e155, 32'h00000000} /* (9, 3, 23) {real, imag} */,
  {32'h3f296665, 32'h00000000} /* (9, 3, 22) {real, imag} */,
  {32'h3f5f3b4b, 32'h00000000} /* (9, 3, 21) {real, imag} */,
  {32'h3f8ad4ed, 32'h00000000} /* (9, 3, 20) {real, imag} */,
  {32'h3f82fbef, 32'h00000000} /* (9, 3, 19) {real, imag} */,
  {32'h3f37fba7, 32'h00000000} /* (9, 3, 18) {real, imag} */,
  {32'h3f2a1cab, 32'h00000000} /* (9, 3, 17) {real, imag} */,
  {32'h3e95dfb6, 32'h00000000} /* (9, 3, 16) {real, imag} */,
  {32'hbf218fd3, 32'h00000000} /* (9, 3, 15) {real, imag} */,
  {32'hbe4ac58c, 32'h00000000} /* (9, 3, 14) {real, imag} */,
  {32'hbf03cbc2, 32'h00000000} /* (9, 3, 13) {real, imag} */,
  {32'hbfb52e2c, 32'h00000000} /* (9, 3, 12) {real, imag} */,
  {32'hbfd6561e, 32'h00000000} /* (9, 3, 11) {real, imag} */,
  {32'hbf51f228, 32'h00000000} /* (9, 3, 10) {real, imag} */,
  {32'hbf423acb, 32'h00000000} /* (9, 3, 9) {real, imag} */,
  {32'hbf82e868, 32'h00000000} /* (9, 3, 8) {real, imag} */,
  {32'hbfb65ae7, 32'h00000000} /* (9, 3, 7) {real, imag} */,
  {32'hbf92d1f2, 32'h00000000} /* (9, 3, 6) {real, imag} */,
  {32'h3e1ef12d, 32'h00000000} /* (9, 3, 5) {real, imag} */,
  {32'h3f487121, 32'h00000000} /* (9, 3, 4) {real, imag} */,
  {32'h3f4fa118, 32'h00000000} /* (9, 3, 3) {real, imag} */,
  {32'h3f60ea5f, 32'h00000000} /* (9, 3, 2) {real, imag} */,
  {32'h3fb72e48, 32'h00000000} /* (9, 3, 1) {real, imag} */,
  {32'h3f786a8e, 32'h00000000} /* (9, 3, 0) {real, imag} */,
  {32'h3ef61611, 32'h00000000} /* (9, 2, 31) {real, imag} */,
  {32'h3f590981, 32'h00000000} /* (9, 2, 30) {real, imag} */,
  {32'h3f58e41b, 32'h00000000} /* (9, 2, 29) {real, imag} */,
  {32'h3f346b5a, 32'h00000000} /* (9, 2, 28) {real, imag} */,
  {32'h3f2f1ca1, 32'h00000000} /* (9, 2, 27) {real, imag} */,
  {32'h3f4e24ae, 32'h00000000} /* (9, 2, 26) {real, imag} */,
  {32'h3fcd6267, 32'h00000000} /* (9, 2, 25) {real, imag} */,
  {32'h3fef82d0, 32'h00000000} /* (9, 2, 24) {real, imag} */,
  {32'h3f610a3e, 32'h00000000} /* (9, 2, 23) {real, imag} */,
  {32'h3f1091a1, 32'h00000000} /* (9, 2, 22) {real, imag} */,
  {32'h3ee1668f, 32'h00000000} /* (9, 2, 21) {real, imag} */,
  {32'h3f477fb8, 32'h00000000} /* (9, 2, 20) {real, imag} */,
  {32'h3fb0b528, 32'h00000000} /* (9, 2, 19) {real, imag} */,
  {32'h3f962a8e, 32'h00000000} /* (9, 2, 18) {real, imag} */,
  {32'h3fd1b220, 32'h00000000} /* (9, 2, 17) {real, imag} */,
  {32'h3f62a73f, 32'h00000000} /* (9, 2, 16) {real, imag} */,
  {32'hbead060b, 32'h00000000} /* (9, 2, 15) {real, imag} */,
  {32'hbe73d93b, 32'h00000000} /* (9, 2, 14) {real, imag} */,
  {32'hbee9e471, 32'h00000000} /* (9, 2, 13) {real, imag} */,
  {32'hbf4ab3a2, 32'h00000000} /* (9, 2, 12) {real, imag} */,
  {32'hbf8cea87, 32'h00000000} /* (9, 2, 11) {real, imag} */,
  {32'hbf9bdcb3, 32'h00000000} /* (9, 2, 10) {real, imag} */,
  {32'hbfaca758, 32'h00000000} /* (9, 2, 9) {real, imag} */,
  {32'hbf90f184, 32'h00000000} /* (9, 2, 8) {real, imag} */,
  {32'hbfb4a49a, 32'h00000000} /* (9, 2, 7) {real, imag} */,
  {32'hbfa5f787, 32'h00000000} /* (9, 2, 6) {real, imag} */,
  {32'h3f05e974, 32'h00000000} /* (9, 2, 5) {real, imag} */,
  {32'h3f5c05d8, 32'h00000000} /* (9, 2, 4) {real, imag} */,
  {32'h3f15f037, 32'h00000000} /* (9, 2, 3) {real, imag} */,
  {32'h3f5cdb09, 32'h00000000} /* (9, 2, 2) {real, imag} */,
  {32'h3f630b4e, 32'h00000000} /* (9, 2, 1) {real, imag} */,
  {32'h3efb5d52, 32'h00000000} /* (9, 2, 0) {real, imag} */,
  {32'h3ef14a69, 32'h00000000} /* (9, 1, 31) {real, imag} */,
  {32'h3f2d08b7, 32'h00000000} /* (9, 1, 30) {real, imag} */,
  {32'h3f5dce3a, 32'h00000000} /* (9, 1, 29) {real, imag} */,
  {32'h3f824ff0, 32'h00000000} /* (9, 1, 28) {real, imag} */,
  {32'h3f8aec44, 32'h00000000} /* (9, 1, 27) {real, imag} */,
  {32'h3f29678f, 32'h00000000} /* (9, 1, 26) {real, imag} */,
  {32'h3fad0ede, 32'h00000000} /* (9, 1, 25) {real, imag} */,
  {32'h3fc6b519, 32'h00000000} /* (9, 1, 24) {real, imag} */,
  {32'h3f07215d, 32'h00000000} /* (9, 1, 23) {real, imag} */,
  {32'h3eb49f19, 32'h00000000} /* (9, 1, 22) {real, imag} */,
  {32'h3eaecbc8, 32'h00000000} /* (9, 1, 21) {real, imag} */,
  {32'h3ef8dc49, 32'h00000000} /* (9, 1, 20) {real, imag} */,
  {32'h3f8c7803, 32'h00000000} /* (9, 1, 19) {real, imag} */,
  {32'h3fa86d3c, 32'h00000000} /* (9, 1, 18) {real, imag} */,
  {32'h3fe0784e, 32'h00000000} /* (9, 1, 17) {real, imag} */,
  {32'h3f73cfec, 32'h00000000} /* (9, 1, 16) {real, imag} */,
  {32'hbe0d8bd3, 32'h00000000} /* (9, 1, 15) {real, imag} */,
  {32'hbf17338a, 32'h00000000} /* (9, 1, 14) {real, imag} */,
  {32'hbf974a28, 32'h00000000} /* (9, 1, 13) {real, imag} */,
  {32'hbf8a558b, 32'h00000000} /* (9, 1, 12) {real, imag} */,
  {32'hbf865c1e, 32'h00000000} /* (9, 1, 11) {real, imag} */,
  {32'hbf8de476, 32'h00000000} /* (9, 1, 10) {real, imag} */,
  {32'hbfab78d8, 32'h00000000} /* (9, 1, 9) {real, imag} */,
  {32'hbf88c242, 32'h00000000} /* (9, 1, 8) {real, imag} */,
  {32'hbf8d0ae8, 32'h00000000} /* (9, 1, 7) {real, imag} */,
  {32'hbf696b6d, 32'h00000000} /* (9, 1, 6) {real, imag} */,
  {32'h3e8329a9, 32'h00000000} /* (9, 1, 5) {real, imag} */,
  {32'h3f336211, 32'h00000000} /* (9, 1, 4) {real, imag} */,
  {32'h3f2aa078, 32'h00000000} /* (9, 1, 3) {real, imag} */,
  {32'h3f3d111a, 32'h00000000} /* (9, 1, 2) {real, imag} */,
  {32'h3f359238, 32'h00000000} /* (9, 1, 1) {real, imag} */,
  {32'h3eda2d01, 32'h00000000} /* (9, 1, 0) {real, imag} */,
  {32'h3ea09aba, 32'h00000000} /* (9, 0, 31) {real, imag} */,
  {32'h3e9dbf5e, 32'h00000000} /* (9, 0, 30) {real, imag} */,
  {32'h3deb12c5, 32'h00000000} /* (9, 0, 29) {real, imag} */,
  {32'h3ea9ccce, 32'h00000000} /* (9, 0, 28) {real, imag} */,
  {32'h3f069af7, 32'h00000000} /* (9, 0, 27) {real, imag} */,
  {32'h3e95880d, 32'h00000000} /* (9, 0, 26) {real, imag} */,
  {32'h3f07c9cb, 32'h00000000} /* (9, 0, 25) {real, imag} */,
  {32'h3f522e78, 32'h00000000} /* (9, 0, 24) {real, imag} */,
  {32'h3ea794e9, 32'h00000000} /* (9, 0, 23) {real, imag} */,
  {32'h3e6316e7, 32'h00000000} /* (9, 0, 22) {real, imag} */,
  {32'h3e79e338, 32'h00000000} /* (9, 0, 21) {real, imag} */,
  {32'h3c2ebfa4, 32'h00000000} /* (9, 0, 20) {real, imag} */,
  {32'h3e41f3f5, 32'h00000000} /* (9, 0, 19) {real, imag} */,
  {32'h3f1da2b3, 32'h00000000} /* (9, 0, 18) {real, imag} */,
  {32'h3f165500, 32'h00000000} /* (9, 0, 17) {real, imag} */,
  {32'h3ebf0894, 32'h00000000} /* (9, 0, 16) {real, imag} */,
  {32'hbb163468, 32'h00000000} /* (9, 0, 15) {real, imag} */,
  {32'hbedee189, 32'h00000000} /* (9, 0, 14) {real, imag} */,
  {32'hbf80db2f, 32'h00000000} /* (9, 0, 13) {real, imag} */,
  {32'hbf58e436, 32'h00000000} /* (9, 0, 12) {real, imag} */,
  {32'hbf3c0244, 32'h00000000} /* (9, 0, 11) {real, imag} */,
  {32'hbf1bf3f3, 32'h00000000} /* (9, 0, 10) {real, imag} */,
  {32'hbf56c862, 32'h00000000} /* (9, 0, 9) {real, imag} */,
  {32'hbf3494a5, 32'h00000000} /* (9, 0, 8) {real, imag} */,
  {32'hbf250fa0, 32'h00000000} /* (9, 0, 7) {real, imag} */,
  {32'hbe8640fd, 32'h00000000} /* (9, 0, 6) {real, imag} */,
  {32'h3d865339, 32'h00000000} /* (9, 0, 5) {real, imag} */,
  {32'h3ecec3bd, 32'h00000000} /* (9, 0, 4) {real, imag} */,
  {32'h3ef4b121, 32'h00000000} /* (9, 0, 3) {real, imag} */,
  {32'h3e97aa42, 32'h00000000} /* (9, 0, 2) {real, imag} */,
  {32'h3e93eeab, 32'h00000000} /* (9, 0, 1) {real, imag} */,
  {32'h3e438507, 32'h00000000} /* (9, 0, 0) {real, imag} */,
  {32'h3d0dfb3d, 32'h00000000} /* (8, 31, 31) {real, imag} */,
  {32'h3e3fc28b, 32'h00000000} /* (8, 31, 30) {real, imag} */,
  {32'h3f1edc34, 32'h00000000} /* (8, 31, 29) {real, imag} */,
  {32'h3f11d831, 32'h00000000} /* (8, 31, 28) {real, imag} */,
  {32'h3f354384, 32'h00000000} /* (8, 31, 27) {real, imag} */,
  {32'h3f3d8fbe, 32'h00000000} /* (8, 31, 26) {real, imag} */,
  {32'h3f3e567e, 32'h00000000} /* (8, 31, 25) {real, imag} */,
  {32'h3f1aae36, 32'h00000000} /* (8, 31, 24) {real, imag} */,
  {32'h3ed90d8b, 32'h00000000} /* (8, 31, 23) {real, imag} */,
  {32'h3f45b7a2, 32'h00000000} /* (8, 31, 22) {real, imag} */,
  {32'h3ed52484, 32'h00000000} /* (8, 31, 21) {real, imag} */,
  {32'hbeb78eca, 32'h00000000} /* (8, 31, 20) {real, imag} */,
  {32'hbe3500f2, 32'h00000000} /* (8, 31, 19) {real, imag} */,
  {32'hbdbb4389, 32'h00000000} /* (8, 31, 18) {real, imag} */,
  {32'hbeaff3f6, 32'h00000000} /* (8, 31, 17) {real, imag} */,
  {32'hbf40cfcf, 32'h00000000} /* (8, 31, 16) {real, imag} */,
  {32'hbf1c775f, 32'h00000000} /* (8, 31, 15) {real, imag} */,
  {32'hbf13a503, 32'h00000000} /* (8, 31, 14) {real, imag} */,
  {32'hbf006845, 32'h00000000} /* (8, 31, 13) {real, imag} */,
  {32'hbef13265, 32'h00000000} /* (8, 31, 12) {real, imag} */,
  {32'hbe8243e6, 32'h00000000} /* (8, 31, 11) {real, imag} */,
  {32'h3f8bd0e7, 32'h00000000} /* (8, 31, 10) {real, imag} */,
  {32'h3eefcc51, 32'h00000000} /* (8, 31, 9) {real, imag} */,
  {32'h3e94a6df, 32'h00000000} /* (8, 31, 8) {real, imag} */,
  {32'h3f35c657, 32'h00000000} /* (8, 31, 7) {real, imag} */,
  {32'h3f05fc52, 32'h00000000} /* (8, 31, 6) {real, imag} */,
  {32'h3eef3cac, 32'h00000000} /* (8, 31, 5) {real, imag} */,
  {32'h3f16c254, 32'h00000000} /* (8, 31, 4) {real, imag} */,
  {32'h3eefb9af, 32'h00000000} /* (8, 31, 3) {real, imag} */,
  {32'h3e9e8345, 32'h00000000} /* (8, 31, 2) {real, imag} */,
  {32'h3ecd339e, 32'h00000000} /* (8, 31, 1) {real, imag} */,
  {32'h3dc64fc0, 32'h00000000} /* (8, 31, 0) {real, imag} */,
  {32'h3eaa9111, 32'h00000000} /* (8, 30, 31) {real, imag} */,
  {32'h3f185eeb, 32'h00000000} /* (8, 30, 30) {real, imag} */,
  {32'h3f306db5, 32'h00000000} /* (8, 30, 29) {real, imag} */,
  {32'h3f886f51, 32'h00000000} /* (8, 30, 28) {real, imag} */,
  {32'h3f973da3, 32'h00000000} /* (8, 30, 27) {real, imag} */,
  {32'h3f48f4b4, 32'h00000000} /* (8, 30, 26) {real, imag} */,
  {32'h3f6d0d93, 32'h00000000} /* (8, 30, 25) {real, imag} */,
  {32'h3f538ccc, 32'h00000000} /* (8, 30, 24) {real, imag} */,
  {32'h3f247cf0, 32'h00000000} /* (8, 30, 23) {real, imag} */,
  {32'h3faca170, 32'h00000000} /* (8, 30, 22) {real, imag} */,
  {32'h3f611d01, 32'h00000000} /* (8, 30, 21) {real, imag} */,
  {32'hbf58e662, 32'h00000000} /* (8, 30, 20) {real, imag} */,
  {32'hbf7a5dd9, 32'h00000000} /* (8, 30, 19) {real, imag} */,
  {32'hbf533472, 32'h00000000} /* (8, 30, 18) {real, imag} */,
  {32'hbf2f9dc1, 32'h00000000} /* (8, 30, 17) {real, imag} */,
  {32'hbf9eea13, 32'h00000000} /* (8, 30, 16) {real, imag} */,
  {32'hbf722647, 32'h00000000} /* (8, 30, 15) {real, imag} */,
  {32'hbf167b80, 32'h00000000} /* (8, 30, 14) {real, imag} */,
  {32'hbf314527, 32'h00000000} /* (8, 30, 13) {real, imag} */,
  {32'hbf382cfd, 32'h00000000} /* (8, 30, 12) {real, imag} */,
  {32'hbef80599, 32'h00000000} /* (8, 30, 11) {real, imag} */,
  {32'h3f8d50b8, 32'h00000000} /* (8, 30, 10) {real, imag} */,
  {32'h3f1c0a8f, 32'h00000000} /* (8, 30, 9) {real, imag} */,
  {32'h3f245c88, 32'h00000000} /* (8, 30, 8) {real, imag} */,
  {32'h3f5d8e76, 32'h00000000} /* (8, 30, 7) {real, imag} */,
  {32'h3f2e970b, 32'h00000000} /* (8, 30, 6) {real, imag} */,
  {32'h3fae42e1, 32'h00000000} /* (8, 30, 5) {real, imag} */,
  {32'h3f94ee4c, 32'h00000000} /* (8, 30, 4) {real, imag} */,
  {32'h3f15e3a1, 32'h00000000} /* (8, 30, 3) {real, imag} */,
  {32'h3f6f0d2a, 32'h00000000} /* (8, 30, 2) {real, imag} */,
  {32'h3f9f90d4, 32'h00000000} /* (8, 30, 1) {real, imag} */,
  {32'h3ea421ea, 32'h00000000} /* (8, 30, 0) {real, imag} */,
  {32'h3f45a2e8, 32'h00000000} /* (8, 29, 31) {real, imag} */,
  {32'h3f8c1ed1, 32'h00000000} /* (8, 29, 30) {real, imag} */,
  {32'h3ec40b82, 32'h00000000} /* (8, 29, 29) {real, imag} */,
  {32'h3ee43a93, 32'h00000000} /* (8, 29, 28) {real, imag} */,
  {32'h3f0855b8, 32'h00000000} /* (8, 29, 27) {real, imag} */,
  {32'h3f0993bf, 32'h00000000} /* (8, 29, 26) {real, imag} */,
  {32'h3f23d4ac, 32'h00000000} /* (8, 29, 25) {real, imag} */,
  {32'h3ef329ea, 32'h00000000} /* (8, 29, 24) {real, imag} */,
  {32'h3f02f585, 32'h00000000} /* (8, 29, 23) {real, imag} */,
  {32'h3f8435e0, 32'h00000000} /* (8, 29, 22) {real, imag} */,
  {32'h3f2a1035, 32'h00000000} /* (8, 29, 21) {real, imag} */,
  {32'hbf9d590c, 32'h00000000} /* (8, 29, 20) {real, imag} */,
  {32'hbf8a4f43, 32'h00000000} /* (8, 29, 19) {real, imag} */,
  {32'hbf8813ee, 32'h00000000} /* (8, 29, 18) {real, imag} */,
  {32'hbf2ea95f, 32'h00000000} /* (8, 29, 17) {real, imag} */,
  {32'hbf5d620e, 32'h00000000} /* (8, 29, 16) {real, imag} */,
  {32'hbf87e1f4, 32'h00000000} /* (8, 29, 15) {real, imag} */,
  {32'hbf610356, 32'h00000000} /* (8, 29, 14) {real, imag} */,
  {32'hbf6bf65c, 32'h00000000} /* (8, 29, 13) {real, imag} */,
  {32'hbf4fb1a1, 32'h00000000} /* (8, 29, 12) {real, imag} */,
  {32'hbf5979f6, 32'h00000000} /* (8, 29, 11) {real, imag} */,
  {32'h3ed5b472, 32'h00000000} /* (8, 29, 10) {real, imag} */,
  {32'h3f13a7f9, 32'h00000000} /* (8, 29, 9) {real, imag} */,
  {32'h3f3a2f35, 32'h00000000} /* (8, 29, 8) {real, imag} */,
  {32'h3ee7786d, 32'h00000000} /* (8, 29, 7) {real, imag} */,
  {32'h3eb8b1fd, 32'h00000000} /* (8, 29, 6) {real, imag} */,
  {32'h3f7760bd, 32'h00000000} /* (8, 29, 5) {real, imag} */,
  {32'h3f88b6a3, 32'h00000000} /* (8, 29, 4) {real, imag} */,
  {32'h3f859f1a, 32'h00000000} /* (8, 29, 3) {real, imag} */,
  {32'h3fb56be3, 32'h00000000} /* (8, 29, 2) {real, imag} */,
  {32'h3fa9ae22, 32'h00000000} /* (8, 29, 1) {real, imag} */,
  {32'h3ebfd2c1, 32'h00000000} /* (8, 29, 0) {real, imag} */,
  {32'h3f1c4ba7, 32'h00000000} /* (8, 28, 31) {real, imag} */,
  {32'h3f8a6a7f, 32'h00000000} /* (8, 28, 30) {real, imag} */,
  {32'h3eb75d62, 32'h00000000} /* (8, 28, 29) {real, imag} */,
  {32'h3e30d2dd, 32'h00000000} /* (8, 28, 28) {real, imag} */,
  {32'h3e256c6c, 32'h00000000} /* (8, 28, 27) {real, imag} */,
  {32'h3f2b396c, 32'h00000000} /* (8, 28, 26) {real, imag} */,
  {32'h3f43e7a4, 32'h00000000} /* (8, 28, 25) {real, imag} */,
  {32'h3f29c667, 32'h00000000} /* (8, 28, 24) {real, imag} */,
  {32'h3f609777, 32'h00000000} /* (8, 28, 23) {real, imag} */,
  {32'h3f417ea5, 32'h00000000} /* (8, 28, 22) {real, imag} */,
  {32'h3f03d52f, 32'h00000000} /* (8, 28, 21) {real, imag} */,
  {32'hbefcd631, 32'h00000000} /* (8, 28, 20) {real, imag} */,
  {32'hbf27fdc9, 32'h00000000} /* (8, 28, 19) {real, imag} */,
  {32'hbf3b452a, 32'h00000000} /* (8, 28, 18) {real, imag} */,
  {32'hbefd5e88, 32'h00000000} /* (8, 28, 17) {real, imag} */,
  {32'hbf342793, 32'h00000000} /* (8, 28, 16) {real, imag} */,
  {32'hbf8599ca, 32'h00000000} /* (8, 28, 15) {real, imag} */,
  {32'hbfb4be6b, 32'h00000000} /* (8, 28, 14) {real, imag} */,
  {32'hbfa06bd1, 32'h00000000} /* (8, 28, 13) {real, imag} */,
  {32'hbf559055, 32'h00000000} /* (8, 28, 12) {real, imag} */,
  {32'hbf8eaa5f, 32'h00000000} /* (8, 28, 11) {real, imag} */,
  {32'h3d9e6bcd, 32'h00000000} /* (8, 28, 10) {real, imag} */,
  {32'h3f3e226f, 32'h00000000} /* (8, 28, 9) {real, imag} */,
  {32'h3f80531b, 32'h00000000} /* (8, 28, 8) {real, imag} */,
  {32'h3f099b4b, 32'h00000000} /* (8, 28, 7) {real, imag} */,
  {32'h3ea8ddcd, 32'h00000000} /* (8, 28, 6) {real, imag} */,
  {32'h3f3aa846, 32'h00000000} /* (8, 28, 5) {real, imag} */,
  {32'h3f9acd89, 32'h00000000} /* (8, 28, 4) {real, imag} */,
  {32'h3f85383a, 32'h00000000} /* (8, 28, 3) {real, imag} */,
  {32'h3f8bfb3a, 32'h00000000} /* (8, 28, 2) {real, imag} */,
  {32'h3f161f16, 32'h00000000} /* (8, 28, 1) {real, imag} */,
  {32'h3e4e4bd6, 32'h00000000} /* (8, 28, 0) {real, imag} */,
  {32'h3f4388a0, 32'h00000000} /* (8, 27, 31) {real, imag} */,
  {32'h3f4af15c, 32'h00000000} /* (8, 27, 30) {real, imag} */,
  {32'h3ed9065f, 32'h00000000} /* (8, 27, 29) {real, imag} */,
  {32'h3f1d096a, 32'h00000000} /* (8, 27, 28) {real, imag} */,
  {32'h3ec25028, 32'h00000000} /* (8, 27, 27) {real, imag} */,
  {32'h3f83e338, 32'h00000000} /* (8, 27, 26) {real, imag} */,
  {32'h3f872496, 32'h00000000} /* (8, 27, 25) {real, imag} */,
  {32'h3f846c0c, 32'h00000000} /* (8, 27, 24) {real, imag} */,
  {32'h3fb2d93e, 32'h00000000} /* (8, 27, 23) {real, imag} */,
  {32'h3f0d568d, 32'h00000000} /* (8, 27, 22) {real, imag} */,
  {32'h3ef398d4, 32'h00000000} /* (8, 27, 21) {real, imag} */,
  {32'hbea04dda, 32'h00000000} /* (8, 27, 20) {real, imag} */,
  {32'hbf3f535b, 32'h00000000} /* (8, 27, 19) {real, imag} */,
  {32'hbf511f45, 32'h00000000} /* (8, 27, 18) {real, imag} */,
  {32'hbf9ae0ab, 32'h00000000} /* (8, 27, 17) {real, imag} */,
  {32'hbfa487ab, 32'h00000000} /* (8, 27, 16) {real, imag} */,
  {32'hbf9de874, 32'h00000000} /* (8, 27, 15) {real, imag} */,
  {32'hbfa2e10d, 32'h00000000} /* (8, 27, 14) {real, imag} */,
  {32'hbf881b6f, 32'h00000000} /* (8, 27, 13) {real, imag} */,
  {32'hbf512d79, 32'h00000000} /* (8, 27, 12) {real, imag} */,
  {32'hbf595a07, 32'h00000000} /* (8, 27, 11) {real, imag} */,
  {32'h3e977589, 32'h00000000} /* (8, 27, 10) {real, imag} */,
  {32'h3f910c86, 32'h00000000} /* (8, 27, 9) {real, imag} */,
  {32'h3fa07e14, 32'h00000000} /* (8, 27, 8) {real, imag} */,
  {32'h3f91e932, 32'h00000000} /* (8, 27, 7) {real, imag} */,
  {32'h3ec5349f, 32'h00000000} /* (8, 27, 6) {real, imag} */,
  {32'h3f6e1b90, 32'h00000000} /* (8, 27, 5) {real, imag} */,
  {32'h3fe9b314, 32'h00000000} /* (8, 27, 4) {real, imag} */,
  {32'h3f61addf, 32'h00000000} /* (8, 27, 3) {real, imag} */,
  {32'h3f176eac, 32'h00000000} /* (8, 27, 2) {real, imag} */,
  {32'h3f4fff30, 32'h00000000} /* (8, 27, 1) {real, imag} */,
  {32'h3f3f64e1, 32'h00000000} /* (8, 27, 0) {real, imag} */,
  {32'h3f31c50a, 32'h00000000} /* (8, 26, 31) {real, imag} */,
  {32'h3f12cd02, 32'h00000000} /* (8, 26, 30) {real, imag} */,
  {32'h3f49b537, 32'h00000000} /* (8, 26, 29) {real, imag} */,
  {32'h3f82a902, 32'h00000000} /* (8, 26, 28) {real, imag} */,
  {32'h3f072e19, 32'h00000000} /* (8, 26, 27) {real, imag} */,
  {32'h3f934ec6, 32'h00000000} /* (8, 26, 26) {real, imag} */,
  {32'h3fa82195, 32'h00000000} /* (8, 26, 25) {real, imag} */,
  {32'h3f6fc320, 32'h00000000} /* (8, 26, 24) {real, imag} */,
  {32'h3f73f1e1, 32'h00000000} /* (8, 26, 23) {real, imag} */,
  {32'h3f17acd5, 32'h00000000} /* (8, 26, 22) {real, imag} */,
  {32'h3e51e4cb, 32'h00000000} /* (8, 26, 21) {real, imag} */,
  {32'hbf3cccf6, 32'h00000000} /* (8, 26, 20) {real, imag} */,
  {32'hbf8de108, 32'h00000000} /* (8, 26, 19) {real, imag} */,
  {32'hbf615531, 32'h00000000} /* (8, 26, 18) {real, imag} */,
  {32'hbf74d1d6, 32'h00000000} /* (8, 26, 17) {real, imag} */,
  {32'hbf89ae11, 32'h00000000} /* (8, 26, 16) {real, imag} */,
  {32'hbf97c2ba, 32'h00000000} /* (8, 26, 15) {real, imag} */,
  {32'hbfbc9b93, 32'h00000000} /* (8, 26, 14) {real, imag} */,
  {32'hbf903b26, 32'h00000000} /* (8, 26, 13) {real, imag} */,
  {32'hbeddfc15, 32'h00000000} /* (8, 26, 12) {real, imag} */,
  {32'hbf1048fa, 32'h00000000} /* (8, 26, 11) {real, imag} */,
  {32'h3ecc30be, 32'h00000000} /* (8, 26, 10) {real, imag} */,
  {32'h3fa4b168, 32'h00000000} /* (8, 26, 9) {real, imag} */,
  {32'h3fa98534, 32'h00000000} /* (8, 26, 8) {real, imag} */,
  {32'h3f9227e3, 32'h00000000} /* (8, 26, 7) {real, imag} */,
  {32'h3ea5f1e6, 32'h00000000} /* (8, 26, 6) {real, imag} */,
  {32'h3f2688b5, 32'h00000000} /* (8, 26, 5) {real, imag} */,
  {32'h3fc1d2bb, 32'h00000000} /* (8, 26, 4) {real, imag} */,
  {32'h3f3adedf, 32'h00000000} /* (8, 26, 3) {real, imag} */,
  {32'h3f289e83, 32'h00000000} /* (8, 26, 2) {real, imag} */,
  {32'h3f742def, 32'h00000000} /* (8, 26, 1) {real, imag} */,
  {32'h3f31a3b9, 32'h00000000} /* (8, 26, 0) {real, imag} */,
  {32'h3f2956cb, 32'h00000000} /* (8, 25, 31) {real, imag} */,
  {32'h3f5efeb4, 32'h00000000} /* (8, 25, 30) {real, imag} */,
  {32'h3f494845, 32'h00000000} /* (8, 25, 29) {real, imag} */,
  {32'h3f9c77c0, 32'h00000000} /* (8, 25, 28) {real, imag} */,
  {32'h3f4a5644, 32'h00000000} /* (8, 25, 27) {real, imag} */,
  {32'h3f5a1a81, 32'h00000000} /* (8, 25, 26) {real, imag} */,
  {32'h3f825af2, 32'h00000000} /* (8, 25, 25) {real, imag} */,
  {32'h3f43c2f0, 32'h00000000} /* (8, 25, 24) {real, imag} */,
  {32'h3f23e8b8, 32'h00000000} /* (8, 25, 23) {real, imag} */,
  {32'h3f1cb0e6, 32'h00000000} /* (8, 25, 22) {real, imag} */,
  {32'h3e31369f, 32'h00000000} /* (8, 25, 21) {real, imag} */,
  {32'hbf51cfd5, 32'h00000000} /* (8, 25, 20) {real, imag} */,
  {32'hbfb0e37c, 32'h00000000} /* (8, 25, 19) {real, imag} */,
  {32'hbf6b36e7, 32'h00000000} /* (8, 25, 18) {real, imag} */,
  {32'hbf183ad2, 32'h00000000} /* (8, 25, 17) {real, imag} */,
  {32'hbf0818a6, 32'h00000000} /* (8, 25, 16) {real, imag} */,
  {32'hbf8a6dfe, 32'h00000000} /* (8, 25, 15) {real, imag} */,
  {32'hbfc6540a, 32'h00000000} /* (8, 25, 14) {real, imag} */,
  {32'hbf90ea56, 32'h00000000} /* (8, 25, 13) {real, imag} */,
  {32'hbee13f7e, 32'h00000000} /* (8, 25, 12) {real, imag} */,
  {32'hbf071a26, 32'h00000000} /* (8, 25, 11) {real, imag} */,
  {32'h3ec93e23, 32'h00000000} /* (8, 25, 10) {real, imag} */,
  {32'h3f84bf8e, 32'h00000000} /* (8, 25, 9) {real, imag} */,
  {32'h3f6b41ee, 32'h00000000} /* (8, 25, 8) {real, imag} */,
  {32'h3f7ecd45, 32'h00000000} /* (8, 25, 7) {real, imag} */,
  {32'h3efb8c23, 32'h00000000} /* (8, 25, 6) {real, imag} */,
  {32'h3f535aa3, 32'h00000000} /* (8, 25, 5) {real, imag} */,
  {32'h3fa69380, 32'h00000000} /* (8, 25, 4) {real, imag} */,
  {32'h3f3cfe0f, 32'h00000000} /* (8, 25, 3) {real, imag} */,
  {32'h3f116895, 32'h00000000} /* (8, 25, 2) {real, imag} */,
  {32'h3f63ea65, 32'h00000000} /* (8, 25, 1) {real, imag} */,
  {32'h3f16b8b2, 32'h00000000} /* (8, 25, 0) {real, imag} */,
  {32'h3f21c37e, 32'h00000000} /* (8, 24, 31) {real, imag} */,
  {32'h3f8f841c, 32'h00000000} /* (8, 24, 30) {real, imag} */,
  {32'h3f1cfe61, 32'h00000000} /* (8, 24, 29) {real, imag} */,
  {32'h3fbf19d9, 32'h00000000} /* (8, 24, 28) {real, imag} */,
  {32'h3fb03814, 32'h00000000} /* (8, 24, 27) {real, imag} */,
  {32'h3fa32195, 32'h00000000} /* (8, 24, 26) {real, imag} */,
  {32'h3f90b09d, 32'h00000000} /* (8, 24, 25) {real, imag} */,
  {32'h3f2ee266, 32'h00000000} /* (8, 24, 24) {real, imag} */,
  {32'h3f00d0fd, 32'h00000000} /* (8, 24, 23) {real, imag} */,
  {32'h3f4c9711, 32'h00000000} /* (8, 24, 22) {real, imag} */,
  {32'h3ec596a3, 32'h00000000} /* (8, 24, 21) {real, imag} */,
  {32'hbf3e148c, 32'h00000000} /* (8, 24, 20) {real, imag} */,
  {32'hbfbe4a24, 32'h00000000} /* (8, 24, 19) {real, imag} */,
  {32'hbf5af9ad, 32'h00000000} /* (8, 24, 18) {real, imag} */,
  {32'hbeb8d635, 32'h00000000} /* (8, 24, 17) {real, imag} */,
  {32'hbf03b08b, 32'h00000000} /* (8, 24, 16) {real, imag} */,
  {32'hbfb91596, 32'h00000000} /* (8, 24, 15) {real, imag} */,
  {32'hbf9c3bd3, 32'h00000000} /* (8, 24, 14) {real, imag} */,
  {32'hbfa60180, 32'h00000000} /* (8, 24, 13) {real, imag} */,
  {32'hbf6e2ca0, 32'h00000000} /* (8, 24, 12) {real, imag} */,
  {32'hbeae5c54, 32'h00000000} /* (8, 24, 11) {real, imag} */,
  {32'h3f5b0d2a, 32'h00000000} /* (8, 24, 10) {real, imag} */,
  {32'h3fa6b651, 32'h00000000} /* (8, 24, 9) {real, imag} */,
  {32'h3f493ba2, 32'h00000000} /* (8, 24, 8) {real, imag} */,
  {32'h3f87f277, 32'h00000000} /* (8, 24, 7) {real, imag} */,
  {32'h3f7b0d10, 32'h00000000} /* (8, 24, 6) {real, imag} */,
  {32'h3f558146, 32'h00000000} /* (8, 24, 5) {real, imag} */,
  {32'h3f9039a5, 32'h00000000} /* (8, 24, 4) {real, imag} */,
  {32'h3f854ff2, 32'h00000000} /* (8, 24, 3) {real, imag} */,
  {32'h3f70ce6f, 32'h00000000} /* (8, 24, 2) {real, imag} */,
  {32'h3f81f5e5, 32'h00000000} /* (8, 24, 1) {real, imag} */,
  {32'h3ed1c10e, 32'h00000000} /* (8, 24, 0) {real, imag} */,
  {32'h3f0617f7, 32'h00000000} /* (8, 23, 31) {real, imag} */,
  {32'h3fafb432, 32'h00000000} /* (8, 23, 30) {real, imag} */,
  {32'h3f993a44, 32'h00000000} /* (8, 23, 29) {real, imag} */,
  {32'h3fab8169, 32'h00000000} /* (8, 23, 28) {real, imag} */,
  {32'h3f99fef0, 32'h00000000} /* (8, 23, 27) {real, imag} */,
  {32'h3f69537a, 32'h00000000} /* (8, 23, 26) {real, imag} */,
  {32'h3f197a8c, 32'h00000000} /* (8, 23, 25) {real, imag} */,
  {32'h3f111ac6, 32'h00000000} /* (8, 23, 24) {real, imag} */,
  {32'h3f5e829a, 32'h00000000} /* (8, 23, 23) {real, imag} */,
  {32'h3f45ec95, 32'h00000000} /* (8, 23, 22) {real, imag} */,
  {32'h3ef93541, 32'h00000000} /* (8, 23, 21) {real, imag} */,
  {32'hbf18fde1, 32'h00000000} /* (8, 23, 20) {real, imag} */,
  {32'hbf914fa3, 32'h00000000} /* (8, 23, 19) {real, imag} */,
  {32'hbf201c4a, 32'h00000000} /* (8, 23, 18) {real, imag} */,
  {32'hbeb7e924, 32'h00000000} /* (8, 23, 17) {real, imag} */,
  {32'hbf08651d, 32'h00000000} /* (8, 23, 16) {real, imag} */,
  {32'hbf54f3ba, 32'h00000000} /* (8, 23, 15) {real, imag} */,
  {32'hbf96f8f6, 32'h00000000} /* (8, 23, 14) {real, imag} */,
  {32'hbfcd08cd, 32'h00000000} /* (8, 23, 13) {real, imag} */,
  {32'hbfa255b7, 32'h00000000} /* (8, 23, 12) {real, imag} */,
  {32'hbf28a5c7, 32'h00000000} /* (8, 23, 11) {real, imag} */,
  {32'h3efd8ac3, 32'h00000000} /* (8, 23, 10) {real, imag} */,
  {32'h3fa1c84c, 32'h00000000} /* (8, 23, 9) {real, imag} */,
  {32'h3f653ada, 32'h00000000} /* (8, 23, 8) {real, imag} */,
  {32'h3fb54710, 32'h00000000} /* (8, 23, 7) {real, imag} */,
  {32'h3f87d312, 32'h00000000} /* (8, 23, 6) {real, imag} */,
  {32'h3f86984d, 32'h00000000} /* (8, 23, 5) {real, imag} */,
  {32'h3f84f14f, 32'h00000000} /* (8, 23, 4) {real, imag} */,
  {32'h3f926ffc, 32'h00000000} /* (8, 23, 3) {real, imag} */,
  {32'h3f7ad760, 32'h00000000} /* (8, 23, 2) {real, imag} */,
  {32'h3f02038b, 32'h00000000} /* (8, 23, 1) {real, imag} */,
  {32'h3dd3980f, 32'h00000000} /* (8, 23, 0) {real, imag} */,
  {32'h3e90768a, 32'h00000000} /* (8, 22, 31) {real, imag} */,
  {32'h3f79fb9f, 32'h00000000} /* (8, 22, 30) {real, imag} */,
  {32'h3fbd49bb, 32'h00000000} /* (8, 22, 29) {real, imag} */,
  {32'h3f2ccfb3, 32'h00000000} /* (8, 22, 28) {real, imag} */,
  {32'h3f333ead, 32'h00000000} /* (8, 22, 27) {real, imag} */,
  {32'h3f3aed09, 32'h00000000} /* (8, 22, 26) {real, imag} */,
  {32'h3f316d98, 32'h00000000} /* (8, 22, 25) {real, imag} */,
  {32'h3f59fa18, 32'h00000000} /* (8, 22, 24) {real, imag} */,
  {32'h3f9eb7e6, 32'h00000000} /* (8, 22, 23) {real, imag} */,
  {32'h3f78dc23, 32'h00000000} /* (8, 22, 22) {real, imag} */,
  {32'h3f4d6164, 32'h00000000} /* (8, 22, 21) {real, imag} */,
  {32'hbe56b0eb, 32'h00000000} /* (8, 22, 20) {real, imag} */,
  {32'hbf65ceef, 32'h00000000} /* (8, 22, 19) {real, imag} */,
  {32'hbf43a102, 32'h00000000} /* (8, 22, 18) {real, imag} */,
  {32'hbf2a1f0e, 32'h00000000} /* (8, 22, 17) {real, imag} */,
  {32'hbf1d18b1, 32'h00000000} /* (8, 22, 16) {real, imag} */,
  {32'hbefd1a04, 32'h00000000} /* (8, 22, 15) {real, imag} */,
  {32'hbf997798, 32'h00000000} /* (8, 22, 14) {real, imag} */,
  {32'hbf837b80, 32'h00000000} /* (8, 22, 13) {real, imag} */,
  {32'hbf5e09b7, 32'h00000000} /* (8, 22, 12) {real, imag} */,
  {32'hbefbf54b, 32'h00000000} /* (8, 22, 11) {real, imag} */,
  {32'h3f5e2cfe, 32'h00000000} /* (8, 22, 10) {real, imag} */,
  {32'h3f5cf977, 32'h00000000} /* (8, 22, 9) {real, imag} */,
  {32'h3f222ad7, 32'h00000000} /* (8, 22, 8) {real, imag} */,
  {32'h3f8c9c50, 32'h00000000} /* (8, 22, 7) {real, imag} */,
  {32'h3f476488, 32'h00000000} /* (8, 22, 6) {real, imag} */,
  {32'h3f78b56c, 32'h00000000} /* (8, 22, 5) {real, imag} */,
  {32'h3f26f609, 32'h00000000} /* (8, 22, 4) {real, imag} */,
  {32'h3f9cdc4c, 32'h00000000} /* (8, 22, 3) {real, imag} */,
  {32'h3f80e761, 32'h00000000} /* (8, 22, 2) {real, imag} */,
  {32'h3ed447d9, 32'h00000000} /* (8, 22, 1) {real, imag} */,
  {32'h3cbbaf20, 32'h00000000} /* (8, 22, 0) {real, imag} */,
  {32'h3e7bd814, 32'h00000000} /* (8, 21, 31) {real, imag} */,
  {32'h3ece2519, 32'h00000000} /* (8, 21, 30) {real, imag} */,
  {32'h3ed2decd, 32'h00000000} /* (8, 21, 29) {real, imag} */,
  {32'h3defb8ed, 32'h00000000} /* (8, 21, 28) {real, imag} */,
  {32'h3e1c4eb9, 32'h00000000} /* (8, 21, 27) {real, imag} */,
  {32'h3d8eef9e, 32'h00000000} /* (8, 21, 26) {real, imag} */,
  {32'h3ea399dd, 32'h00000000} /* (8, 21, 25) {real, imag} */,
  {32'h3df2b57a, 32'h00000000} /* (8, 21, 24) {real, imag} */,
  {32'h3e5005d6, 32'h00000000} /* (8, 21, 23) {real, imag} */,
  {32'h3e31da8b, 32'h00000000} /* (8, 21, 22) {real, imag} */,
  {32'h3ef17190, 32'h00000000} /* (8, 21, 21) {real, imag} */,
  {32'hbe9700ef, 32'h00000000} /* (8, 21, 20) {real, imag} */,
  {32'hbf6cd551, 32'h00000000} /* (8, 21, 19) {real, imag} */,
  {32'hbf0ba919, 32'h00000000} /* (8, 21, 18) {real, imag} */,
  {32'hbeca4106, 32'h00000000} /* (8, 21, 17) {real, imag} */,
  {32'hbea12f96, 32'h00000000} /* (8, 21, 16) {real, imag} */,
  {32'hbe916f99, 32'h00000000} /* (8, 21, 15) {real, imag} */,
  {32'hbf3b550c, 32'h00000000} /* (8, 21, 14) {real, imag} */,
  {32'hbdb6b741, 32'h00000000} /* (8, 21, 13) {real, imag} */,
  {32'h3d5aa9a0, 32'h00000000} /* (8, 21, 12) {real, imag} */,
  {32'hbdd7209c, 32'h00000000} /* (8, 21, 11) {real, imag} */,
  {32'h3f20e65d, 32'h00000000} /* (8, 21, 10) {real, imag} */,
  {32'h3ee6e31b, 32'h00000000} /* (8, 21, 9) {real, imag} */,
  {32'h3dc884cc, 32'h00000000} /* (8, 21, 8) {real, imag} */,
  {32'h3e066b5c, 32'h00000000} /* (8, 21, 7) {real, imag} */,
  {32'hbbefdf4f, 32'h00000000} /* (8, 21, 6) {real, imag} */,
  {32'h3ce8b92e, 32'h00000000} /* (8, 21, 5) {real, imag} */,
  {32'hbd8673cc, 32'h00000000} /* (8, 21, 4) {real, imag} */,
  {32'h3f2efba5, 32'h00000000} /* (8, 21, 3) {real, imag} */,
  {32'h3ee6a061, 32'h00000000} /* (8, 21, 2) {real, imag} */,
  {32'h3e0b77fb, 32'h00000000} /* (8, 21, 1) {real, imag} */,
  {32'hbddfceae, 32'h00000000} /* (8, 21, 0) {real, imag} */,
  {32'hbe8f9715, 32'h00000000} /* (8, 20, 31) {real, imag} */,
  {32'hbf7229d6, 32'h00000000} /* (8, 20, 30) {real, imag} */,
  {32'hbf45b399, 32'h00000000} /* (8, 20, 29) {real, imag} */,
  {32'hbf0f663d, 32'h00000000} /* (8, 20, 28) {real, imag} */,
  {32'hbf5af59a, 32'h00000000} /* (8, 20, 27) {real, imag} */,
  {32'hbf70f05d, 32'h00000000} /* (8, 20, 26) {real, imag} */,
  {32'hbf0cb41e, 32'h00000000} /* (8, 20, 25) {real, imag} */,
  {32'hbf1d506f, 32'h00000000} /* (8, 20, 24) {real, imag} */,
  {32'hbf4b1c9f, 32'h00000000} /* (8, 20, 23) {real, imag} */,
  {32'hbf312189, 32'h00000000} /* (8, 20, 22) {real, imag} */,
  {32'hbe8b5c18, 32'h00000000} /* (8, 20, 21) {real, imag} */,
  {32'h3e8997c0, 32'h00000000} /* (8, 20, 20) {real, imag} */,
  {32'h3e890b33, 32'h00000000} /* (8, 20, 19) {real, imag} */,
  {32'h3ee90fdc, 32'h00000000} /* (8, 20, 18) {real, imag} */,
  {32'h3f471d12, 32'h00000000} /* (8, 20, 17) {real, imag} */,
  {32'h3ef40447, 32'h00000000} /* (8, 20, 16) {real, imag} */,
  {32'h3eceefd2, 32'h00000000} /* (8, 20, 15) {real, imag} */,
  {32'h3ee33042, 32'h00000000} /* (8, 20, 14) {real, imag} */,
  {32'h3f85b8c7, 32'h00000000} /* (8, 20, 13) {real, imag} */,
  {32'h3f648f4d, 32'h00000000} /* (8, 20, 12) {real, imag} */,
  {32'h3effed08, 32'h00000000} /* (8, 20, 11) {real, imag} */,
  {32'hbdfc220c, 32'h00000000} /* (8, 20, 10) {real, imag} */,
  {32'hbf4636d5, 32'h00000000} /* (8, 20, 9) {real, imag} */,
  {32'hbfa07a19, 32'h00000000} /* (8, 20, 8) {real, imag} */,
  {32'hbf9da651, 32'h00000000} /* (8, 20, 7) {real, imag} */,
  {32'hbf735a53, 32'h00000000} /* (8, 20, 6) {real, imag} */,
  {32'hbf80a70b, 32'h00000000} /* (8, 20, 5) {real, imag} */,
  {32'hbfa1ce83, 32'h00000000} /* (8, 20, 4) {real, imag} */,
  {32'hbf4b1338, 32'h00000000} /* (8, 20, 3) {real, imag} */,
  {32'hbf4e2837, 32'h00000000} /* (8, 20, 2) {real, imag} */,
  {32'hbf5c6ace, 32'h00000000} /* (8, 20, 1) {real, imag} */,
  {32'hbeaf7292, 32'h00000000} /* (8, 20, 0) {real, imag} */,
  {32'hbeb24405, 32'h00000000} /* (8, 19, 31) {real, imag} */,
  {32'hbf2e7893, 32'h00000000} /* (8, 19, 30) {real, imag} */,
  {32'hbf3ae54d, 32'h00000000} /* (8, 19, 29) {real, imag} */,
  {32'hbf56c792, 32'h00000000} /* (8, 19, 28) {real, imag} */,
  {32'hbf520d7e, 32'h00000000} /* (8, 19, 27) {real, imag} */,
  {32'hbf9d6019, 32'h00000000} /* (8, 19, 26) {real, imag} */,
  {32'hbf66c999, 32'h00000000} /* (8, 19, 25) {real, imag} */,
  {32'hbf237d8e, 32'h00000000} /* (8, 19, 24) {real, imag} */,
  {32'hbf48d1a4, 32'h00000000} /* (8, 19, 23) {real, imag} */,
  {32'hbf387633, 32'h00000000} /* (8, 19, 22) {real, imag} */,
  {32'hbe2458a2, 32'h00000000} /* (8, 19, 21) {real, imag} */,
  {32'h3fa77ca7, 32'h00000000} /* (8, 19, 20) {real, imag} */,
  {32'h3fa2cd94, 32'h00000000} /* (8, 19, 19) {real, imag} */,
  {32'h3f1782ec, 32'h00000000} /* (8, 19, 18) {real, imag} */,
  {32'h3f5fec19, 32'h00000000} /* (8, 19, 17) {real, imag} */,
  {32'h3f6a7e8d, 32'h00000000} /* (8, 19, 16) {real, imag} */,
  {32'h3f82f70f, 32'h00000000} /* (8, 19, 15) {real, imag} */,
  {32'h3faa9b52, 32'h00000000} /* (8, 19, 14) {real, imag} */,
  {32'h3fc42368, 32'h00000000} /* (8, 19, 13) {real, imag} */,
  {32'h3f2e6ad0, 32'h00000000} /* (8, 19, 12) {real, imag} */,
  {32'h3ee90a14, 32'h00000000} /* (8, 19, 11) {real, imag} */,
  {32'hbec68266, 32'h00000000} /* (8, 19, 10) {real, imag} */,
  {32'hbfcc3cab, 32'h00000000} /* (8, 19, 9) {real, imag} */,
  {32'hbffbf4cf, 32'h00000000} /* (8, 19, 8) {real, imag} */,
  {32'hbfac13e0, 32'h00000000} /* (8, 19, 7) {real, imag} */,
  {32'hbf4f864f, 32'h00000000} /* (8, 19, 6) {real, imag} */,
  {32'hbf2c89c7, 32'h00000000} /* (8, 19, 5) {real, imag} */,
  {32'hbf8df5d7, 32'h00000000} /* (8, 19, 4) {real, imag} */,
  {32'hbfd04eb2, 32'h00000000} /* (8, 19, 3) {real, imag} */,
  {32'hbfac2821, 32'h00000000} /* (8, 19, 2) {real, imag} */,
  {32'hbf58bb9f, 32'h00000000} /* (8, 19, 1) {real, imag} */,
  {32'hbe99afc7, 32'h00000000} /* (8, 19, 0) {real, imag} */,
  {32'hbf8261bd, 32'h00000000} /* (8, 18, 31) {real, imag} */,
  {32'hbfb65467, 32'h00000000} /* (8, 18, 30) {real, imag} */,
  {32'hbf4b58ba, 32'h00000000} /* (8, 18, 29) {real, imag} */,
  {32'hbf0ca55e, 32'h00000000} /* (8, 18, 28) {real, imag} */,
  {32'hbf4b83dc, 32'h00000000} /* (8, 18, 27) {real, imag} */,
  {32'hbf727b52, 32'h00000000} /* (8, 18, 26) {real, imag} */,
  {32'hbf7413a2, 32'h00000000} /* (8, 18, 25) {real, imag} */,
  {32'hbfb4ba65, 32'h00000000} /* (8, 18, 24) {real, imag} */,
  {32'hbfd78b72, 32'h00000000} /* (8, 18, 23) {real, imag} */,
  {32'hbf6c044b, 32'h00000000} /* (8, 18, 22) {real, imag} */,
  {32'h3e49add0, 32'h00000000} /* (8, 18, 21) {real, imag} */,
  {32'h3fc97d94, 32'h00000000} /* (8, 18, 20) {real, imag} */,
  {32'h3f9ec785, 32'h00000000} /* (8, 18, 19) {real, imag} */,
  {32'h3ef88ab1, 32'h00000000} /* (8, 18, 18) {real, imag} */,
  {32'h3f5d28ab, 32'h00000000} /* (8, 18, 17) {real, imag} */,
  {32'h3fa40e62, 32'h00000000} /* (8, 18, 16) {real, imag} */,
  {32'h3f9f602e, 32'h00000000} /* (8, 18, 15) {real, imag} */,
  {32'h3fb87556, 32'h00000000} /* (8, 18, 14) {real, imag} */,
  {32'h3f9aaa47, 32'h00000000} /* (8, 18, 13) {real, imag} */,
  {32'h3f7163ff, 32'h00000000} /* (8, 18, 12) {real, imag} */,
  {32'h3ea93422, 32'h00000000} /* (8, 18, 11) {real, imag} */,
  {32'hbf2b3ad3, 32'h00000000} /* (8, 18, 10) {real, imag} */,
  {32'hbf3b0059, 32'h00000000} /* (8, 18, 9) {real, imag} */,
  {32'hbf8b2fd7, 32'h00000000} /* (8, 18, 8) {real, imag} */,
  {32'hbf5cc6e7, 32'h00000000} /* (8, 18, 7) {real, imag} */,
  {32'hbf41c689, 32'h00000000} /* (8, 18, 6) {real, imag} */,
  {32'hbee873ec, 32'h00000000} /* (8, 18, 5) {real, imag} */,
  {32'hbf71f959, 32'h00000000} /* (8, 18, 4) {real, imag} */,
  {32'hbfe62355, 32'h00000000} /* (8, 18, 3) {real, imag} */,
  {32'hbfae4035, 32'h00000000} /* (8, 18, 2) {real, imag} */,
  {32'hbf9ed573, 32'h00000000} /* (8, 18, 1) {real, imag} */,
  {32'hbf597fce, 32'h00000000} /* (8, 18, 0) {real, imag} */,
  {32'hbf96fc7f, 32'h00000000} /* (8, 17, 31) {real, imag} */,
  {32'hc018aa1f, 32'h00000000} /* (8, 17, 30) {real, imag} */,
  {32'hbfc53533, 32'h00000000} /* (8, 17, 29) {real, imag} */,
  {32'hbf89ab45, 32'h00000000} /* (8, 17, 28) {real, imag} */,
  {32'hbf8a32cc, 32'h00000000} /* (8, 17, 27) {real, imag} */,
  {32'hbf0d6e97, 32'h00000000} /* (8, 17, 26) {real, imag} */,
  {32'hbf3db485, 32'h00000000} /* (8, 17, 25) {real, imag} */,
  {32'hbfc74ab6, 32'h00000000} /* (8, 17, 24) {real, imag} */,
  {32'hbfec6074, 32'h00000000} /* (8, 17, 23) {real, imag} */,
  {32'hbf4fe785, 32'h00000000} /* (8, 17, 22) {real, imag} */,
  {32'h3ecdc867, 32'h00000000} /* (8, 17, 21) {real, imag} */,
  {32'h3f7455c5, 32'h00000000} /* (8, 17, 20) {real, imag} */,
  {32'h3eff6363, 32'h00000000} /* (8, 17, 19) {real, imag} */,
  {32'h3eadb120, 32'h00000000} /* (8, 17, 18) {real, imag} */,
  {32'h3f1960ab, 32'h00000000} /* (8, 17, 17) {real, imag} */,
  {32'h3f3c4d85, 32'h00000000} /* (8, 17, 16) {real, imag} */,
  {32'h3f3a8c04, 32'h00000000} /* (8, 17, 15) {real, imag} */,
  {32'h3f26f422, 32'h00000000} /* (8, 17, 14) {real, imag} */,
  {32'h3ef721fa, 32'h00000000} /* (8, 17, 13) {real, imag} */,
  {32'h3ed027a6, 32'h00000000} /* (8, 17, 12) {real, imag} */,
  {32'h3cde52d7, 32'h00000000} /* (8, 17, 11) {real, imag} */,
  {32'hbef2db0b, 32'h00000000} /* (8, 17, 10) {real, imag} */,
  {32'hbf1b67e1, 32'h00000000} /* (8, 17, 9) {real, imag} */,
  {32'hbf85a417, 32'h00000000} /* (8, 17, 8) {real, imag} */,
  {32'hbf26daf7, 32'h00000000} /* (8, 17, 7) {real, imag} */,
  {32'hbf896bf3, 32'h00000000} /* (8, 17, 6) {real, imag} */,
  {32'hbf80e6f7, 32'h00000000} /* (8, 17, 5) {real, imag} */,
  {32'hbfaf4f8f, 32'h00000000} /* (8, 17, 4) {real, imag} */,
  {32'hbfff6031, 32'h00000000} /* (8, 17, 3) {real, imag} */,
  {32'hbfb84e1a, 32'h00000000} /* (8, 17, 2) {real, imag} */,
  {32'hbf800b71, 32'h00000000} /* (8, 17, 1) {real, imag} */,
  {32'hbf058c3e, 32'h00000000} /* (8, 17, 0) {real, imag} */,
  {32'hbf5a63c9, 32'h00000000} /* (8, 16, 31) {real, imag} */,
  {32'hc0025314, 32'h00000000} /* (8, 16, 30) {real, imag} */,
  {32'hbf9984f6, 32'h00000000} /* (8, 16, 29) {real, imag} */,
  {32'hbf889496, 32'h00000000} /* (8, 16, 28) {real, imag} */,
  {32'hbf6a5f5e, 32'h00000000} /* (8, 16, 27) {real, imag} */,
  {32'hbea72cea, 32'h00000000} /* (8, 16, 26) {real, imag} */,
  {32'hbf208ba0, 32'h00000000} /* (8, 16, 25) {real, imag} */,
  {32'hbf7094d8, 32'h00000000} /* (8, 16, 24) {real, imag} */,
  {32'hbf8e16b1, 32'h00000000} /* (8, 16, 23) {real, imag} */,
  {32'hbf585ad4, 32'h00000000} /* (8, 16, 22) {real, imag} */,
  {32'h3e02541c, 32'h00000000} /* (8, 16, 21) {real, imag} */,
  {32'h3f3b64ee, 32'h00000000} /* (8, 16, 20) {real, imag} */,
  {32'h3f276a50, 32'h00000000} /* (8, 16, 19) {real, imag} */,
  {32'h3f8834a0, 32'h00000000} /* (8, 16, 18) {real, imag} */,
  {32'h3f943f5c, 32'h00000000} /* (8, 16, 17) {real, imag} */,
  {32'h3f69596e, 32'h00000000} /* (8, 16, 16) {real, imag} */,
  {32'h3f9505e8, 32'h00000000} /* (8, 16, 15) {real, imag} */,
  {32'h3f6cc6bc, 32'h00000000} /* (8, 16, 14) {real, imag} */,
  {32'h3f685956, 32'h00000000} /* (8, 16, 13) {real, imag} */,
  {32'h3f213c5a, 32'h00000000} /* (8, 16, 12) {real, imag} */,
  {32'h3e736990, 32'h00000000} /* (8, 16, 11) {real, imag} */,
  {32'hbe8d564d, 32'h00000000} /* (8, 16, 10) {real, imag} */,
  {32'hbf204ebb, 32'h00000000} /* (8, 16, 9) {real, imag} */,
  {32'hbf5d4f6a, 32'h00000000} /* (8, 16, 8) {real, imag} */,
  {32'hbf1bee3d, 32'h00000000} /* (8, 16, 7) {real, imag} */,
  {32'hbf683d47, 32'h00000000} /* (8, 16, 6) {real, imag} */,
  {32'hbf557fc7, 32'h00000000} /* (8, 16, 5) {real, imag} */,
  {32'hbf978055, 32'h00000000} /* (8, 16, 4) {real, imag} */,
  {32'hbfc20afc, 32'h00000000} /* (8, 16, 3) {real, imag} */,
  {32'hbfb85e83, 32'h00000000} /* (8, 16, 2) {real, imag} */,
  {32'hbf8c9745, 32'h00000000} /* (8, 16, 1) {real, imag} */,
  {32'hbebb58cf, 32'h00000000} /* (8, 16, 0) {real, imag} */,
  {32'hbf6a2b38, 32'h00000000} /* (8, 15, 31) {real, imag} */,
  {32'hbfd586c8, 32'h00000000} /* (8, 15, 30) {real, imag} */,
  {32'hbfab697b, 32'h00000000} /* (8, 15, 29) {real, imag} */,
  {32'hbf61a857, 32'h00000000} /* (8, 15, 28) {real, imag} */,
  {32'hbf2075c0, 32'h00000000} /* (8, 15, 27) {real, imag} */,
  {32'hbf367f82, 32'h00000000} /* (8, 15, 26) {real, imag} */,
  {32'hbf6f1b02, 32'h00000000} /* (8, 15, 25) {real, imag} */,
  {32'hbf882436, 32'h00000000} /* (8, 15, 24) {real, imag} */,
  {32'hbf5c4e2f, 32'h00000000} /* (8, 15, 23) {real, imag} */,
  {32'hbf3071ea, 32'h00000000} /* (8, 15, 22) {real, imag} */,
  {32'h3e54f6ba, 32'h00000000} /* (8, 15, 21) {real, imag} */,
  {32'h3f683e74, 32'h00000000} /* (8, 15, 20) {real, imag} */,
  {32'h3f0560d8, 32'h00000000} /* (8, 15, 19) {real, imag} */,
  {32'h3f93a72e, 32'h00000000} /* (8, 15, 18) {real, imag} */,
  {32'h3fc2274f, 32'h00000000} /* (8, 15, 17) {real, imag} */,
  {32'h3fa158e9, 32'h00000000} /* (8, 15, 16) {real, imag} */,
  {32'h3f854bc7, 32'h00000000} /* (8, 15, 15) {real, imag} */,
  {32'h3f8779bc, 32'h00000000} /* (8, 15, 14) {real, imag} */,
  {32'h3fa96548, 32'h00000000} /* (8, 15, 13) {real, imag} */,
  {32'h3f8f2f1c, 32'h00000000} /* (8, 15, 12) {real, imag} */,
  {32'h3f2701c2, 32'h00000000} /* (8, 15, 11) {real, imag} */,
  {32'hbe2d1320, 32'h00000000} /* (8, 15, 10) {real, imag} */,
  {32'hbf1215bd, 32'h00000000} /* (8, 15, 9) {real, imag} */,
  {32'hbf788aa5, 32'h00000000} /* (8, 15, 8) {real, imag} */,
  {32'hbfbafca9, 32'h00000000} /* (8, 15, 7) {real, imag} */,
  {32'hbf82be92, 32'h00000000} /* (8, 15, 6) {real, imag} */,
  {32'hbee969a2, 32'h00000000} /* (8, 15, 5) {real, imag} */,
  {32'hbf4dad2b, 32'h00000000} /* (8, 15, 4) {real, imag} */,
  {32'hbf85e9e7, 32'h00000000} /* (8, 15, 3) {real, imag} */,
  {32'hbf96c4a0, 32'h00000000} /* (8, 15, 2) {real, imag} */,
  {32'hbf82c304, 32'h00000000} /* (8, 15, 1) {real, imag} */,
  {32'hbf0f4f90, 32'h00000000} /* (8, 15, 0) {real, imag} */,
  {32'hbef5a169, 32'h00000000} /* (8, 14, 31) {real, imag} */,
  {32'hbf5cf1d5, 32'h00000000} /* (8, 14, 30) {real, imag} */,
  {32'hbf18d121, 32'h00000000} /* (8, 14, 29) {real, imag} */,
  {32'hbf58e3af, 32'h00000000} /* (8, 14, 28) {real, imag} */,
  {32'hbf87e100, 32'h00000000} /* (8, 14, 27) {real, imag} */,
  {32'hbf832f6b, 32'h00000000} /* (8, 14, 26) {real, imag} */,
  {32'hbf98cd55, 32'h00000000} /* (8, 14, 25) {real, imag} */,
  {32'hbf25fe11, 32'h00000000} /* (8, 14, 24) {real, imag} */,
  {32'hbf5d42cb, 32'h00000000} /* (8, 14, 23) {real, imag} */,
  {32'hbfa70fe5, 32'h00000000} /* (8, 14, 22) {real, imag} */,
  {32'hbf0d169f, 32'h00000000} /* (8, 14, 21) {real, imag} */,
  {32'h3f023b48, 32'h00000000} /* (8, 14, 20) {real, imag} */,
  {32'h3e7bfcd6, 32'h00000000} /* (8, 14, 19) {real, imag} */,
  {32'h3f11a73e, 32'h00000000} /* (8, 14, 18) {real, imag} */,
  {32'h3f560172, 32'h00000000} /* (8, 14, 17) {real, imag} */,
  {32'h3f2005fd, 32'h00000000} /* (8, 14, 16) {real, imag} */,
  {32'h3f09c936, 32'h00000000} /* (8, 14, 15) {real, imag} */,
  {32'h3f1ae5e5, 32'h00000000} /* (8, 14, 14) {real, imag} */,
  {32'h3f83b2d6, 32'h00000000} /* (8, 14, 13) {real, imag} */,
  {32'h3f5f9efa, 32'h00000000} /* (8, 14, 12) {real, imag} */,
  {32'h3f68e791, 32'h00000000} /* (8, 14, 11) {real, imag} */,
  {32'h3e1701fd, 32'h00000000} /* (8, 14, 10) {real, imag} */,
  {32'hbf84020c, 32'h00000000} /* (8, 14, 9) {real, imag} */,
  {32'hbfb3ef76, 32'h00000000} /* (8, 14, 8) {real, imag} */,
  {32'hbfc4895f, 32'h00000000} /* (8, 14, 7) {real, imag} */,
  {32'hbf5a50a0, 32'h00000000} /* (8, 14, 6) {real, imag} */,
  {32'hbf096ba2, 32'h00000000} /* (8, 14, 5) {real, imag} */,
  {32'hbf1cd8b1, 32'h00000000} /* (8, 14, 4) {real, imag} */,
  {32'hbf2de8cb, 32'h00000000} /* (8, 14, 3) {real, imag} */,
  {32'hbf5bb79c, 32'h00000000} /* (8, 14, 2) {real, imag} */,
  {32'hbf8fa194, 32'h00000000} /* (8, 14, 1) {real, imag} */,
  {32'hbf2dc39b, 32'h00000000} /* (8, 14, 0) {real, imag} */,
  {32'hbebfc9fa, 32'h00000000} /* (8, 13, 31) {real, imag} */,
  {32'hbf317e6b, 32'h00000000} /* (8, 13, 30) {real, imag} */,
  {32'hbee7731a, 32'h00000000} /* (8, 13, 29) {real, imag} */,
  {32'hbf495d7f, 32'h00000000} /* (8, 13, 28) {real, imag} */,
  {32'hbf6c5863, 32'h00000000} /* (8, 13, 27) {real, imag} */,
  {32'hbf506fba, 32'h00000000} /* (8, 13, 26) {real, imag} */,
  {32'hbf2d0c61, 32'h00000000} /* (8, 13, 25) {real, imag} */,
  {32'hbf2679dd, 32'h00000000} /* (8, 13, 24) {real, imag} */,
  {32'hbf6213ae, 32'h00000000} /* (8, 13, 23) {real, imag} */,
  {32'hbfbc42c4, 32'h00000000} /* (8, 13, 22) {real, imag} */,
  {32'hbf19d6f4, 32'h00000000} /* (8, 13, 21) {real, imag} */,
  {32'h3f539e3a, 32'h00000000} /* (8, 13, 20) {real, imag} */,
  {32'h3f0b25c0, 32'h00000000} /* (8, 13, 19) {real, imag} */,
  {32'h3f050998, 32'h00000000} /* (8, 13, 18) {real, imag} */,
  {32'h3f418575, 32'h00000000} /* (8, 13, 17) {real, imag} */,
  {32'h3f6c25c0, 32'h00000000} /* (8, 13, 16) {real, imag} */,
  {32'h3f7c7d52, 32'h00000000} /* (8, 13, 15) {real, imag} */,
  {32'h3f0de082, 32'h00000000} /* (8, 13, 14) {real, imag} */,
  {32'h3f4715a2, 32'h00000000} /* (8, 13, 13) {real, imag} */,
  {32'h3f93cace, 32'h00000000} /* (8, 13, 12) {real, imag} */,
  {32'h3f96fb77, 32'h00000000} /* (8, 13, 11) {real, imag} */,
  {32'hbe0d272e, 32'h00000000} /* (8, 13, 10) {real, imag} */,
  {32'hbf9e606d, 32'h00000000} /* (8, 13, 9) {real, imag} */,
  {32'hbf5ec573, 32'h00000000} /* (8, 13, 8) {real, imag} */,
  {32'hbf309132, 32'h00000000} /* (8, 13, 7) {real, imag} */,
  {32'hbf80f79b, 32'h00000000} /* (8, 13, 6) {real, imag} */,
  {32'hbfa8a3e3, 32'h00000000} /* (8, 13, 5) {real, imag} */,
  {32'hbf5733d4, 32'h00000000} /* (8, 13, 4) {real, imag} */,
  {32'hbf3cf304, 32'h00000000} /* (8, 13, 3) {real, imag} */,
  {32'hbf613b53, 32'h00000000} /* (8, 13, 2) {real, imag} */,
  {32'hbf84426b, 32'h00000000} /* (8, 13, 1) {real, imag} */,
  {32'hbf138fb9, 32'h00000000} /* (8, 13, 0) {real, imag} */,
  {32'h3dbd9d46, 32'h00000000} /* (8, 12, 31) {real, imag} */,
  {32'hbeafab64, 32'h00000000} /* (8, 12, 30) {real, imag} */,
  {32'hbf47f994, 32'h00000000} /* (8, 12, 29) {real, imag} */,
  {32'hbfcf6698, 32'h00000000} /* (8, 12, 28) {real, imag} */,
  {32'hbfbc9220, 32'h00000000} /* (8, 12, 27) {real, imag} */,
  {32'hbf8f1fb4, 32'h00000000} /* (8, 12, 26) {real, imag} */,
  {32'hbf94bec3, 32'h00000000} /* (8, 12, 25) {real, imag} */,
  {32'hbf877fe5, 32'h00000000} /* (8, 12, 24) {real, imag} */,
  {32'hbf0fa790, 32'h00000000} /* (8, 12, 23) {real, imag} */,
  {32'hbed61782, 32'h00000000} /* (8, 12, 22) {real, imag} */,
  {32'h3d8d3d11, 32'h00000000} /* (8, 12, 21) {real, imag} */,
  {32'h3f849a3a, 32'h00000000} /* (8, 12, 20) {real, imag} */,
  {32'h3f0f9180, 32'h00000000} /* (8, 12, 19) {real, imag} */,
  {32'h3e686922, 32'h00000000} /* (8, 12, 18) {real, imag} */,
  {32'h3f2a6956, 32'h00000000} /* (8, 12, 17) {real, imag} */,
  {32'h3f7a2b12, 32'h00000000} /* (8, 12, 16) {real, imag} */,
  {32'h3f991f84, 32'h00000000} /* (8, 12, 15) {real, imag} */,
  {32'h3f25a236, 32'h00000000} /* (8, 12, 14) {real, imag} */,
  {32'h3efe2221, 32'h00000000} /* (8, 12, 13) {real, imag} */,
  {32'h3f3dddff, 32'h00000000} /* (8, 12, 12) {real, imag} */,
  {32'h3f41a832, 32'h00000000} /* (8, 12, 11) {real, imag} */,
  {32'hbeb62d84, 32'h00000000} /* (8, 12, 10) {real, imag} */,
  {32'hbfa8721d, 32'h00000000} /* (8, 12, 9) {real, imag} */,
  {32'hbf2307c3, 32'h00000000} /* (8, 12, 8) {real, imag} */,
  {32'hbf1486a7, 32'h00000000} /* (8, 12, 7) {real, imag} */,
  {32'hbf8c57e1, 32'h00000000} /* (8, 12, 6) {real, imag} */,
  {32'hbf868895, 32'h00000000} /* (8, 12, 5) {real, imag} */,
  {32'hbf5037d2, 32'h00000000} /* (8, 12, 4) {real, imag} */,
  {32'hbf5cd779, 32'h00000000} /* (8, 12, 3) {real, imag} */,
  {32'hbf1d2b81, 32'h00000000} /* (8, 12, 2) {real, imag} */,
  {32'hbefb15dc, 32'h00000000} /* (8, 12, 1) {real, imag} */,
  {32'hbe66225e, 32'h00000000} /* (8, 12, 0) {real, imag} */,
  {32'h3e26041e, 32'h00000000} /* (8, 11, 31) {real, imag} */,
  {32'hbdf85f23, 32'h00000000} /* (8, 11, 30) {real, imag} */,
  {32'hbf10458d, 32'h00000000} /* (8, 11, 29) {real, imag} */,
  {32'hbf9d82be, 32'h00000000} /* (8, 11, 28) {real, imag} */,
  {32'hbf9a8977, 32'h00000000} /* (8, 11, 27) {real, imag} */,
  {32'hbf34d197, 32'h00000000} /* (8, 11, 26) {real, imag} */,
  {32'hbf6169d6, 32'h00000000} /* (8, 11, 25) {real, imag} */,
  {32'hbf9a57f9, 32'h00000000} /* (8, 11, 24) {real, imag} */,
  {32'hbe889a93, 32'h00000000} /* (8, 11, 23) {real, imag} */,
  {32'hbc981fe4, 32'h00000000} /* (8, 11, 22) {real, imag} */,
  {32'h3e1836ab, 32'h00000000} /* (8, 11, 21) {real, imag} */,
  {32'h3ed42aef, 32'h00000000} /* (8, 11, 20) {real, imag} */,
  {32'h3e03f6e2, 32'h00000000} /* (8, 11, 19) {real, imag} */,
  {32'hbe21d5b3, 32'h00000000} /* (8, 11, 18) {real, imag} */,
  {32'h3d02848e, 32'h00000000} /* (8, 11, 17) {real, imag} */,
  {32'h3f076813, 32'h00000000} /* (8, 11, 16) {real, imag} */,
  {32'h3f1fde6c, 32'h00000000} /* (8, 11, 15) {real, imag} */,
  {32'h3f024049, 32'h00000000} /* (8, 11, 14) {real, imag} */,
  {32'h3f3e19d9, 32'h00000000} /* (8, 11, 13) {real, imag} */,
  {32'h3f33abe4, 32'h00000000} /* (8, 11, 12) {real, imag} */,
  {32'h3f1fd2e9, 32'h00000000} /* (8, 11, 11) {real, imag} */,
  {32'hbec54cdc, 32'h00000000} /* (8, 11, 10) {real, imag} */,
  {32'hbf5d3d11, 32'h00000000} /* (8, 11, 9) {real, imag} */,
  {32'hbf2a5127, 32'h00000000} /* (8, 11, 8) {real, imag} */,
  {32'hbeed939e, 32'h00000000} /* (8, 11, 7) {real, imag} */,
  {32'hbf88464e, 32'h00000000} /* (8, 11, 6) {real, imag} */,
  {32'hbf82bf41, 32'h00000000} /* (8, 11, 5) {real, imag} */,
  {32'hbdc9abf0, 32'h00000000} /* (8, 11, 4) {real, imag} */,
  {32'hbdd1858b, 32'h00000000} /* (8, 11, 3) {real, imag} */,
  {32'hbf5951ae, 32'h00000000} /* (8, 11, 2) {real, imag} */,
  {32'hbf922285, 32'h00000000} /* (8, 11, 1) {real, imag} */,
  {32'hbecaab67, 32'h00000000} /* (8, 11, 0) {real, imag} */,
  {32'h3e400ea8, 32'h00000000} /* (8, 10, 31) {real, imag} */,
  {32'h3e6f4859, 32'h00000000} /* (8, 10, 30) {real, imag} */,
  {32'h3e488ac7, 32'h00000000} /* (8, 10, 29) {real, imag} */,
  {32'h3ed70b1a, 32'h00000000} /* (8, 10, 28) {real, imag} */,
  {32'h3f2b7847, 32'h00000000} /* (8, 10, 27) {real, imag} */,
  {32'h3e3d7fd8, 32'h00000000} /* (8, 10, 26) {real, imag} */,
  {32'h3e18187d, 32'h00000000} /* (8, 10, 25) {real, imag} */,
  {32'hbd01127c, 32'h00000000} /* (8, 10, 24) {real, imag} */,
  {32'h3f62d9c6, 32'h00000000} /* (8, 10, 23) {real, imag} */,
  {32'h3f32451d, 32'h00000000} /* (8, 10, 22) {real, imag} */,
  {32'h3efca37d, 32'h00000000} /* (8, 10, 21) {real, imag} */,
  {32'h3e42dcfa, 32'h00000000} /* (8, 10, 20) {real, imag} */,
  {32'hbf0ba232, 32'h00000000} /* (8, 10, 19) {real, imag} */,
  {32'hbf7d0639, 32'h00000000} /* (8, 10, 18) {real, imag} */,
  {32'hbf293d0b, 32'h00000000} /* (8, 10, 17) {real, imag} */,
  {32'hbf063d67, 32'h00000000} /* (8, 10, 16) {real, imag} */,
  {32'hbeffb5a7, 32'h00000000} /* (8, 10, 15) {real, imag} */,
  {32'hbec80a4f, 32'h00000000} /* (8, 10, 14) {real, imag} */,
  {32'hbea8727e, 32'h00000000} /* (8, 10, 13) {real, imag} */,
  {32'hbe91871f, 32'h00000000} /* (8, 10, 12) {real, imag} */,
  {32'hbe9f1519, 32'h00000000} /* (8, 10, 11) {real, imag} */,
  {32'hbd68af48, 32'h00000000} /* (8, 10, 10) {real, imag} */,
  {32'h3e842178, 32'h00000000} /* (8, 10, 9) {real, imag} */,
  {32'h3ef835c5, 32'h00000000} /* (8, 10, 8) {real, imag} */,
  {32'h3f0dc194, 32'h00000000} /* (8, 10, 7) {real, imag} */,
  {32'h3ba601d1, 32'h00000000} /* (8, 10, 6) {real, imag} */,
  {32'h3d50f1cb, 32'h00000000} /* (8, 10, 5) {real, imag} */,
  {32'h3f2d6d0c, 32'h00000000} /* (8, 10, 4) {real, imag} */,
  {32'h3f2b1cc7, 32'h00000000} /* (8, 10, 3) {real, imag} */,
  {32'hbd9a2b01, 32'h00000000} /* (8, 10, 2) {real, imag} */,
  {32'hbe31e30d, 32'h00000000} /* (8, 10, 1) {real, imag} */,
  {32'h3e3e1a13, 32'h00000000} /* (8, 10, 0) {real, imag} */,
  {32'h3f0a836a, 32'h00000000} /* (8, 9, 31) {real, imag} */,
  {32'h3f26d03a, 32'h00000000} /* (8, 9, 30) {real, imag} */,
  {32'h3f7f0019, 32'h00000000} /* (8, 9, 29) {real, imag} */,
  {32'h3f6d6643, 32'h00000000} /* (8, 9, 28) {real, imag} */,
  {32'h3f5ed9d3, 32'h00000000} /* (8, 9, 27) {real, imag} */,
  {32'h3f11473c, 32'h00000000} /* (8, 9, 26) {real, imag} */,
  {32'h3f768cb9, 32'h00000000} /* (8, 9, 25) {real, imag} */,
  {32'h3f6f4352, 32'h00000000} /* (8, 9, 24) {real, imag} */,
  {32'h3f6f7c84, 32'h00000000} /* (8, 9, 23) {real, imag} */,
  {32'h3f425068, 32'h00000000} /* (8, 9, 22) {real, imag} */,
  {32'h3f10b61a, 32'h00000000} /* (8, 9, 21) {real, imag} */,
  {32'h3df6de9a, 32'h00000000} /* (8, 9, 20) {real, imag} */,
  {32'hbf4375ec, 32'h00000000} /* (8, 9, 19) {real, imag} */,
  {32'hbfa193b5, 32'h00000000} /* (8, 9, 18) {real, imag} */,
  {32'hbf546659, 32'h00000000} /* (8, 9, 17) {real, imag} */,
  {32'hbf51f82b, 32'h00000000} /* (8, 9, 16) {real, imag} */,
  {32'hbf91912b, 32'h00000000} /* (8, 9, 15) {real, imag} */,
  {32'hbf9ec883, 32'h00000000} /* (8, 9, 14) {real, imag} */,
  {32'hbffe1769, 32'h00000000} /* (8, 9, 13) {real, imag} */,
  {32'hbf90d749, 32'h00000000} /* (8, 9, 12) {real, imag} */,
  {32'hbebbc6a7, 32'h00000000} /* (8, 9, 11) {real, imag} */,
  {32'h3de65223, 32'h00000000} /* (8, 9, 10) {real, imag} */,
  {32'h3f13be0d, 32'h00000000} /* (8, 9, 9) {real, imag} */,
  {32'h3f851d1a, 32'h00000000} /* (8, 9, 8) {real, imag} */,
  {32'h3f87f038, 32'h00000000} /* (8, 9, 7) {real, imag} */,
  {32'h3f313408, 32'h00000000} /* (8, 9, 6) {real, imag} */,
  {32'h3f56d4ec, 32'h00000000} /* (8, 9, 5) {real, imag} */,
  {32'h3f4790e0, 32'h00000000} /* (8, 9, 4) {real, imag} */,
  {32'h3f21accd, 32'h00000000} /* (8, 9, 3) {real, imag} */,
  {32'h3f0ae102, 32'h00000000} /* (8, 9, 2) {real, imag} */,
  {32'h3f345585, 32'h00000000} /* (8, 9, 1) {real, imag} */,
  {32'h3f292403, 32'h00000000} /* (8, 9, 0) {real, imag} */,
  {32'h3f4cbae2, 32'h00000000} /* (8, 8, 31) {real, imag} */,
  {32'h3f3bd424, 32'h00000000} /* (8, 8, 30) {real, imag} */,
  {32'h3f9b308b, 32'h00000000} /* (8, 8, 29) {real, imag} */,
  {32'h3f47ed56, 32'h00000000} /* (8, 8, 28) {real, imag} */,
  {32'h3f43a303, 32'h00000000} /* (8, 8, 27) {real, imag} */,
  {32'h3f86a835, 32'h00000000} /* (8, 8, 26) {real, imag} */,
  {32'h3f68654a, 32'h00000000} /* (8, 8, 25) {real, imag} */,
  {32'h3fb3ad6c, 32'h00000000} /* (8, 8, 24) {real, imag} */,
  {32'h3f9ee0e2, 32'h00000000} /* (8, 8, 23) {real, imag} */,
  {32'h3f8bc794, 32'h00000000} /* (8, 8, 22) {real, imag} */,
  {32'h3e233882, 32'h00000000} /* (8, 8, 21) {real, imag} */,
  {32'hbef86d13, 32'h00000000} /* (8, 8, 20) {real, imag} */,
  {32'hbf54a8d6, 32'h00000000} /* (8, 8, 19) {real, imag} */,
  {32'hbf9bb048, 32'h00000000} /* (8, 8, 18) {real, imag} */,
  {32'hbf905f5c, 32'h00000000} /* (8, 8, 17) {real, imag} */,
  {32'hbf74abd0, 32'h00000000} /* (8, 8, 16) {real, imag} */,
  {32'hbfb79c98, 32'h00000000} /* (8, 8, 15) {real, imag} */,
  {32'hbfbdca9e, 32'h00000000} /* (8, 8, 14) {real, imag} */,
  {32'hbfb3845e, 32'h00000000} /* (8, 8, 13) {real, imag} */,
  {32'hbf4e2c84, 32'h00000000} /* (8, 8, 12) {real, imag} */,
  {32'hbf06346a, 32'h00000000} /* (8, 8, 11) {real, imag} */,
  {32'h3f09a30c, 32'h00000000} /* (8, 8, 10) {real, imag} */,
  {32'h3f43e965, 32'h00000000} /* (8, 8, 9) {real, imag} */,
  {32'h3f69ca30, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'h3f39e95c, 32'h00000000} /* (8, 8, 7) {real, imag} */,
  {32'h3f7c29f5, 32'h00000000} /* (8, 8, 6) {real, imag} */,
  {32'h3f54ffb4, 32'h00000000} /* (8, 8, 5) {real, imag} */,
  {32'h3f730afb, 32'h00000000} /* (8, 8, 4) {real, imag} */,
  {32'h3f1e3414, 32'h00000000} /* (8, 8, 3) {real, imag} */,
  {32'h3ef99236, 32'h00000000} /* (8, 8, 2) {real, imag} */,
  {32'h3f1dd758, 32'h00000000} /* (8, 8, 1) {real, imag} */,
  {32'h3f1f5673, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h3ea3a890, 32'h00000000} /* (8, 7, 31) {real, imag} */,
  {32'h3f451ce8, 32'h00000000} /* (8, 7, 30) {real, imag} */,
  {32'h3fbaba1d, 32'h00000000} /* (8, 7, 29) {real, imag} */,
  {32'h3f68b98b, 32'h00000000} /* (8, 7, 28) {real, imag} */,
  {32'h3f3b0f89, 32'h00000000} /* (8, 7, 27) {real, imag} */,
  {32'h3ee9667f, 32'h00000000} /* (8, 7, 26) {real, imag} */,
  {32'h3ef89262, 32'h00000000} /* (8, 7, 25) {real, imag} */,
  {32'h3f9544b4, 32'h00000000} /* (8, 7, 24) {real, imag} */,
  {32'h3f891f28, 32'h00000000} /* (8, 7, 23) {real, imag} */,
  {32'h3f99552c, 32'h00000000} /* (8, 7, 22) {real, imag} */,
  {32'h3e9f3cbc, 32'h00000000} /* (8, 7, 21) {real, imag} */,
  {32'hbf51cdfc, 32'h00000000} /* (8, 7, 20) {real, imag} */,
  {32'hbfab0bea, 32'h00000000} /* (8, 7, 19) {real, imag} */,
  {32'hbfb6d931, 32'h00000000} /* (8, 7, 18) {real, imag} */,
  {32'hbfb3a625, 32'h00000000} /* (8, 7, 17) {real, imag} */,
  {32'hbfb85425, 32'h00000000} /* (8, 7, 16) {real, imag} */,
  {32'hbfcfb37c, 32'h00000000} /* (8, 7, 15) {real, imag} */,
  {32'hbfa7f1e1, 32'h00000000} /* (8, 7, 14) {real, imag} */,
  {32'hbf981ea6, 32'h00000000} /* (8, 7, 13) {real, imag} */,
  {32'hbf787179, 32'h00000000} /* (8, 7, 12) {real, imag} */,
  {32'hbf84f3a4, 32'h00000000} /* (8, 7, 11) {real, imag} */,
  {32'h3efac6bb, 32'h00000000} /* (8, 7, 10) {real, imag} */,
  {32'h3fa91fd7, 32'h00000000} /* (8, 7, 9) {real, imag} */,
  {32'h3fec4e08, 32'h00000000} /* (8, 7, 8) {real, imag} */,
  {32'h3f743970, 32'h00000000} /* (8, 7, 7) {real, imag} */,
  {32'h3f15bd46, 32'h00000000} /* (8, 7, 6) {real, imag} */,
  {32'h3f359c48, 32'h00000000} /* (8, 7, 5) {real, imag} */,
  {32'h3f7be2d0, 32'h00000000} /* (8, 7, 4) {real, imag} */,
  {32'h3f6dc514, 32'h00000000} /* (8, 7, 3) {real, imag} */,
  {32'h3f1ffd5f, 32'h00000000} /* (8, 7, 2) {real, imag} */,
  {32'h3f376471, 32'h00000000} /* (8, 7, 1) {real, imag} */,
  {32'h3f2056bd, 32'h00000000} /* (8, 7, 0) {real, imag} */,
  {32'h3e60621c, 32'h00000000} /* (8, 6, 31) {real, imag} */,
  {32'h3f112247, 32'h00000000} /* (8, 6, 30) {real, imag} */,
  {32'h3f7174c8, 32'h00000000} /* (8, 6, 29) {real, imag} */,
  {32'h3f6e59ee, 32'h00000000} /* (8, 6, 28) {real, imag} */,
  {32'h3f59b02f, 32'h00000000} /* (8, 6, 27) {real, imag} */,
  {32'h3f5ed4a1, 32'h00000000} /* (8, 6, 26) {real, imag} */,
  {32'h3f301caa, 32'h00000000} /* (8, 6, 25) {real, imag} */,
  {32'h3f6f931c, 32'h00000000} /* (8, 6, 24) {real, imag} */,
  {32'h3f6d18c1, 32'h00000000} /* (8, 6, 23) {real, imag} */,
  {32'h3f7b7f94, 32'h00000000} /* (8, 6, 22) {real, imag} */,
  {32'h3edf6d30, 32'h00000000} /* (8, 6, 21) {real, imag} */,
  {32'hbf321627, 32'h00000000} /* (8, 6, 20) {real, imag} */,
  {32'hbfa0dccd, 32'h00000000} /* (8, 6, 19) {real, imag} */,
  {32'hbf84c730, 32'h00000000} /* (8, 6, 18) {real, imag} */,
  {32'hbf83a059, 32'h00000000} /* (8, 6, 17) {real, imag} */,
  {32'hbfaf9612, 32'h00000000} /* (8, 6, 16) {real, imag} */,
  {32'hbfbf0529, 32'h00000000} /* (8, 6, 15) {real, imag} */,
  {32'hbfba9043, 32'h00000000} /* (8, 6, 14) {real, imag} */,
  {32'hbfbbcf08, 32'h00000000} /* (8, 6, 13) {real, imag} */,
  {32'hbf99f230, 32'h00000000} /* (8, 6, 12) {real, imag} */,
  {32'hbf781d97, 32'h00000000} /* (8, 6, 11) {real, imag} */,
  {32'h3d50bfba, 32'h00000000} /* (8, 6, 10) {real, imag} */,
  {32'h3f22ed67, 32'h00000000} /* (8, 6, 9) {real, imag} */,
  {32'h3f9264ee, 32'h00000000} /* (8, 6, 8) {real, imag} */,
  {32'h3f2d2d84, 32'h00000000} /* (8, 6, 7) {real, imag} */,
  {32'h3f2c031d, 32'h00000000} /* (8, 6, 6) {real, imag} */,
  {32'h3f88c8f0, 32'h00000000} /* (8, 6, 5) {real, imag} */,
  {32'h3f437a2d, 32'h00000000} /* (8, 6, 4) {real, imag} */,
  {32'h3f47052e, 32'h00000000} /* (8, 6, 3) {real, imag} */,
  {32'h3f92c984, 32'h00000000} /* (8, 6, 2) {real, imag} */,
  {32'h3f4ca922, 32'h00000000} /* (8, 6, 1) {real, imag} */,
  {32'h3ed3b445, 32'h00000000} /* (8, 6, 0) {real, imag} */,
  {32'h3f10003e, 32'h00000000} /* (8, 5, 31) {real, imag} */,
  {32'h3eb98180, 32'h00000000} /* (8, 5, 30) {real, imag} */,
  {32'h3f4eaead, 32'h00000000} /* (8, 5, 29) {real, imag} */,
  {32'h3f9d9479, 32'h00000000} /* (8, 5, 28) {real, imag} */,
  {32'h3fa80865, 32'h00000000} /* (8, 5, 27) {real, imag} */,
  {32'h3f90d43f, 32'h00000000} /* (8, 5, 26) {real, imag} */,
  {32'h3f70f2c9, 32'h00000000} /* (8, 5, 25) {real, imag} */,
  {32'h3f4e82ce, 32'h00000000} /* (8, 5, 24) {real, imag} */,
  {32'h3f8b3cd3, 32'h00000000} /* (8, 5, 23) {real, imag} */,
  {32'h3fc2ebaa, 32'h00000000} /* (8, 5, 22) {real, imag} */,
  {32'h3f681878, 32'h00000000} /* (8, 5, 21) {real, imag} */,
  {32'h3f50c099, 32'h00000000} /* (8, 5, 20) {real, imag} */,
  {32'h3f1922d6, 32'h00000000} /* (8, 5, 19) {real, imag} */,
  {32'h3e8d95e8, 32'h00000000} /* (8, 5, 18) {real, imag} */,
  {32'h3ebdeb66, 32'h00000000} /* (8, 5, 17) {real, imag} */,
  {32'hbe9347bf, 32'h00000000} /* (8, 5, 16) {real, imag} */,
  {32'hbf9c3364, 32'h00000000} /* (8, 5, 15) {real, imag} */,
  {32'hbfbd613c, 32'h00000000} /* (8, 5, 14) {real, imag} */,
  {32'hbf8d2d72, 32'h00000000} /* (8, 5, 13) {real, imag} */,
  {32'hbf8232d2, 32'h00000000} /* (8, 5, 12) {real, imag} */,
  {32'hbf6346c4, 32'h00000000} /* (8, 5, 11) {real, imag} */,
  {32'hbee3171f, 32'h00000000} /* (8, 5, 10) {real, imag} */,
  {32'hbebc2926, 32'h00000000} /* (8, 5, 9) {real, imag} */,
  {32'hbe76acf4, 32'h00000000} /* (8, 5, 8) {real, imag} */,
  {32'h3dacc222, 32'h00000000} /* (8, 5, 7) {real, imag} */,
  {32'hbe8a162f, 32'h00000000} /* (8, 5, 6) {real, imag} */,
  {32'h3f5a7310, 32'h00000000} /* (8, 5, 5) {real, imag} */,
  {32'h3f32b87e, 32'h00000000} /* (8, 5, 4) {real, imag} */,
  {32'h3ef239d6, 32'h00000000} /* (8, 5, 3) {real, imag} */,
  {32'h3f821cd3, 32'h00000000} /* (8, 5, 2) {real, imag} */,
  {32'h3fcc256a, 32'h00000000} /* (8, 5, 1) {real, imag} */,
  {32'h3f8bd305, 32'h00000000} /* (8, 5, 0) {real, imag} */,
  {32'h3ef91be8, 32'h00000000} /* (8, 4, 31) {real, imag} */,
  {32'h3f1a243b, 32'h00000000} /* (8, 4, 30) {real, imag} */,
  {32'h3ed30e26, 32'h00000000} /* (8, 4, 29) {real, imag} */,
  {32'h3f752a33, 32'h00000000} /* (8, 4, 28) {real, imag} */,
  {32'h3fd4a1c0, 32'h00000000} /* (8, 4, 27) {real, imag} */,
  {32'h3f5514c3, 32'h00000000} /* (8, 4, 26) {real, imag} */,
  {32'h3ef87dc9, 32'h00000000} /* (8, 4, 25) {real, imag} */,
  {32'h3f28bfad, 32'h00000000} /* (8, 4, 24) {real, imag} */,
  {32'h3f72c6b1, 32'h00000000} /* (8, 4, 23) {real, imag} */,
  {32'h3fbbec8a, 32'h00000000} /* (8, 4, 22) {real, imag} */,
  {32'h3fa7b90a, 32'h00000000} /* (8, 4, 21) {real, imag} */,
  {32'h3f9bd111, 32'h00000000} /* (8, 4, 20) {real, imag} */,
  {32'h3f7f55e9, 32'h00000000} /* (8, 4, 19) {real, imag} */,
  {32'h3f6b8feb, 32'h00000000} /* (8, 4, 18) {real, imag} */,
  {32'h3f8151ea, 32'h00000000} /* (8, 4, 17) {real, imag} */,
  {32'h3ee02ff0, 32'h00000000} /* (8, 4, 16) {real, imag} */,
  {32'hbf4ff23c, 32'h00000000} /* (8, 4, 15) {real, imag} */,
  {32'hbefc88c8, 32'h00000000} /* (8, 4, 14) {real, imag} */,
  {32'hbee33372, 32'h00000000} /* (8, 4, 13) {real, imag} */,
  {32'hbfa0d388, 32'h00000000} /* (8, 4, 12) {real, imag} */,
  {32'hbf830b95, 32'h00000000} /* (8, 4, 11) {real, imag} */,
  {32'hbf030d1e, 32'h00000000} /* (8, 4, 10) {real, imag} */,
  {32'hbf321c99, 32'h00000000} /* (8, 4, 9) {real, imag} */,
  {32'hbf1fbee8, 32'h00000000} /* (8, 4, 8) {real, imag} */,
  {32'hbe8865b6, 32'h00000000} /* (8, 4, 7) {real, imag} */,
  {32'hbf314249, 32'h00000000} /* (8, 4, 6) {real, imag} */,
  {32'h3e990104, 32'h00000000} /* (8, 4, 5) {real, imag} */,
  {32'h3f2a882a, 32'h00000000} /* (8, 4, 4) {real, imag} */,
  {32'h3f7770ca, 32'h00000000} /* (8, 4, 3) {real, imag} */,
  {32'h3f634c0e, 32'h00000000} /* (8, 4, 2) {real, imag} */,
  {32'h3f9307db, 32'h00000000} /* (8, 4, 1) {real, imag} */,
  {32'h3f2fd0ab, 32'h00000000} /* (8, 4, 0) {real, imag} */,
  {32'h3ec901cf, 32'h00000000} /* (8, 3, 31) {real, imag} */,
  {32'h3f5f99ef, 32'h00000000} /* (8, 3, 30) {real, imag} */,
  {32'h3f5a7881, 32'h00000000} /* (8, 3, 29) {real, imag} */,
  {32'h3f0c44f3, 32'h00000000} /* (8, 3, 28) {real, imag} */,
  {32'h3f5a027b, 32'h00000000} /* (8, 3, 27) {real, imag} */,
  {32'h3f854aed, 32'h00000000} /* (8, 3, 26) {real, imag} */,
  {32'h3f92a398, 32'h00000000} /* (8, 3, 25) {real, imag} */,
  {32'h3fb87ef1, 32'h00000000} /* (8, 3, 24) {real, imag} */,
  {32'h3f57b88b, 32'h00000000} /* (8, 3, 23) {real, imag} */,
  {32'h3f2880c4, 32'h00000000} /* (8, 3, 22) {real, imag} */,
  {32'h3f864dab, 32'h00000000} /* (8, 3, 21) {real, imag} */,
  {32'h3f624746, 32'h00000000} /* (8, 3, 20) {real, imag} */,
  {32'h3f98a52d, 32'h00000000} /* (8, 3, 19) {real, imag} */,
  {32'h3f6d8477, 32'h00000000} /* (8, 3, 18) {real, imag} */,
  {32'h3f0c1c56, 32'h00000000} /* (8, 3, 17) {real, imag} */,
  {32'h3eb1fcf9, 32'h00000000} /* (8, 3, 16) {real, imag} */,
  {32'hbec2871e, 32'h00000000} /* (8, 3, 15) {real, imag} */,
  {32'hbe767268, 32'h00000000} /* (8, 3, 14) {real, imag} */,
  {32'hbf67c5b9, 32'h00000000} /* (8, 3, 13) {real, imag} */,
  {32'hbfcfc2f5, 32'h00000000} /* (8, 3, 12) {real, imag} */,
  {32'hbf59509c, 32'h00000000} /* (8, 3, 11) {real, imag} */,
  {32'hbf043e1c, 32'h00000000} /* (8, 3, 10) {real, imag} */,
  {32'hbf7caa8b, 32'h00000000} /* (8, 3, 9) {real, imag} */,
  {32'hbf669dca, 32'h00000000} /* (8, 3, 8) {real, imag} */,
  {32'hbfa7065e, 32'h00000000} /* (8, 3, 7) {real, imag} */,
  {32'hbfaaeb5a, 32'h00000000} /* (8, 3, 6) {real, imag} */,
  {32'h3e80554e, 32'h00000000} /* (8, 3, 5) {real, imag} */,
  {32'h3f54193f, 32'h00000000} /* (8, 3, 4) {real, imag} */,
  {32'h3f931c69, 32'h00000000} /* (8, 3, 3) {real, imag} */,
  {32'h3f559986, 32'h00000000} /* (8, 3, 2) {real, imag} */,
  {32'h3f8438ea, 32'h00000000} /* (8, 3, 1) {real, imag} */,
  {32'h3ee1c926, 32'h00000000} /* (8, 3, 0) {real, imag} */,
  {32'h3ef607f0, 32'h00000000} /* (8, 2, 31) {real, imag} */,
  {32'h3f59a5cd, 32'h00000000} /* (8, 2, 30) {real, imag} */,
  {32'h3f8739bd, 32'h00000000} /* (8, 2, 29) {real, imag} */,
  {32'h3f439942, 32'h00000000} /* (8, 2, 28) {real, imag} */,
  {32'h3f371cf6, 32'h00000000} /* (8, 2, 27) {real, imag} */,
  {32'h3f9522dc, 32'h00000000} /* (8, 2, 26) {real, imag} */,
  {32'h3fbc7705, 32'h00000000} /* (8, 2, 25) {real, imag} */,
  {32'h3fe18373, 32'h00000000} /* (8, 2, 24) {real, imag} */,
  {32'h3fa4c936, 32'h00000000} /* (8, 2, 23) {real, imag} */,
  {32'h3f2db0e6, 32'h00000000} /* (8, 2, 22) {real, imag} */,
  {32'h3f3d676d, 32'h00000000} /* (8, 2, 21) {real, imag} */,
  {32'h3f73eafb, 32'h00000000} /* (8, 2, 20) {real, imag} */,
  {32'h3faf2fc8, 32'h00000000} /* (8, 2, 19) {real, imag} */,
  {32'h3f635707, 32'h00000000} /* (8, 2, 18) {real, imag} */,
  {32'h3f84f032, 32'h00000000} /* (8, 2, 17) {real, imag} */,
  {32'h3f52ac89, 32'h00000000} /* (8, 2, 16) {real, imag} */,
  {32'hbe09c7df, 32'h00000000} /* (8, 2, 15) {real, imag} */,
  {32'hbf08bb21, 32'h00000000} /* (8, 2, 14) {real, imag} */,
  {32'hbf6dd128, 32'h00000000} /* (8, 2, 13) {real, imag} */,
  {32'hbf844106, 32'h00000000} /* (8, 2, 12) {real, imag} */,
  {32'hbf59a0c3, 32'h00000000} /* (8, 2, 11) {real, imag} */,
  {32'hbf972167, 32'h00000000} /* (8, 2, 10) {real, imag} */,
  {32'hbfe61b64, 32'h00000000} /* (8, 2, 9) {real, imag} */,
  {32'hbfa963c0, 32'h00000000} /* (8, 2, 8) {real, imag} */,
  {32'hbfaedb23, 32'h00000000} /* (8, 2, 7) {real, imag} */,
  {32'hbfb64660, 32'h00000000} /* (8, 2, 6) {real, imag} */,
  {32'h3f812120, 32'h00000000} /* (8, 2, 5) {real, imag} */,
  {32'h3fc101c6, 32'h00000000} /* (8, 2, 4) {real, imag} */,
  {32'h3f9a10ee, 32'h00000000} /* (8, 2, 3) {real, imag} */,
  {32'h3fa8f1aa, 32'h00000000} /* (8, 2, 2) {real, imag} */,
  {32'h3fa7cc4c, 32'h00000000} /* (8, 2, 1) {real, imag} */,
  {32'h3f1a3fc2, 32'h00000000} /* (8, 2, 0) {real, imag} */,
  {32'h3ea0a2b7, 32'h00000000} /* (8, 1, 31) {real, imag} */,
  {32'h3f084a96, 32'h00000000} /* (8, 1, 30) {real, imag} */,
  {32'h3f5844d0, 32'h00000000} /* (8, 1, 29) {real, imag} */,
  {32'h3f570cc0, 32'h00000000} /* (8, 1, 28) {real, imag} */,
  {32'h3f90ae3a, 32'h00000000} /* (8, 1, 27) {real, imag} */,
  {32'h3f95b299, 32'h00000000} /* (8, 1, 26) {real, imag} */,
  {32'h3fc77170, 32'h00000000} /* (8, 1, 25) {real, imag} */,
  {32'h3fce884a, 32'h00000000} /* (8, 1, 24) {real, imag} */,
  {32'h3f60db25, 32'h00000000} /* (8, 1, 23) {real, imag} */,
  {32'h3e2a0b31, 32'h00000000} /* (8, 1, 22) {real, imag} */,
  {32'h3f131163, 32'h00000000} /* (8, 1, 21) {real, imag} */,
  {32'h3f660acf, 32'h00000000} /* (8, 1, 20) {real, imag} */,
  {32'h3f78a2d3, 32'h00000000} /* (8, 1, 19) {real, imag} */,
  {32'h3f722aad, 32'h00000000} /* (8, 1, 18) {real, imag} */,
  {32'h3f8275d4, 32'h00000000} /* (8, 1, 17) {real, imag} */,
  {32'h3f6bab8e, 32'h00000000} /* (8, 1, 16) {real, imag} */,
  {32'hbd3f9c4b, 32'h00000000} /* (8, 1, 15) {real, imag} */,
  {32'hbf4f51a8, 32'h00000000} /* (8, 1, 14) {real, imag} */,
  {32'hbf3afe5d, 32'h00000000} /* (8, 1, 13) {real, imag} */,
  {32'hbf6d5715, 32'h00000000} /* (8, 1, 12) {real, imag} */,
  {32'hbf4a3aa8, 32'h00000000} /* (8, 1, 11) {real, imag} */,
  {32'hbf6c1625, 32'h00000000} /* (8, 1, 10) {real, imag} */,
  {32'hbfdee0ab, 32'h00000000} /* (8, 1, 9) {real, imag} */,
  {32'hbfa99210, 32'h00000000} /* (8, 1, 8) {real, imag} */,
  {32'hbf849431, 32'h00000000} /* (8, 1, 7) {real, imag} */,
  {32'hbf606b81, 32'h00000000} /* (8, 1, 6) {real, imag} */,
  {32'h3e9143e5, 32'h00000000} /* (8, 1, 5) {real, imag} */,
  {32'h3f6d1a5a, 32'h00000000} /* (8, 1, 4) {real, imag} */,
  {32'h3f9c8883, 32'h00000000} /* (8, 1, 3) {real, imag} */,
  {32'h3f859c4b, 32'h00000000} /* (8, 1, 2) {real, imag} */,
  {32'h3f63a77e, 32'h00000000} /* (8, 1, 1) {real, imag} */,
  {32'h3f01dfcf, 32'h00000000} /* (8, 1, 0) {real, imag} */,
  {32'h3db78d27, 32'h00000000} /* (8, 0, 31) {real, imag} */,
  {32'h3e6cf447, 32'h00000000} /* (8, 0, 30) {real, imag} */,
  {32'h3ec9aeba, 32'h00000000} /* (8, 0, 29) {real, imag} */,
  {32'h3e72b806, 32'h00000000} /* (8, 0, 28) {real, imag} */,
  {32'h3f36980c, 32'h00000000} /* (8, 0, 27) {real, imag} */,
  {32'h3f4c6d7a, 32'h00000000} /* (8, 0, 26) {real, imag} */,
  {32'h3f61bfb2, 32'h00000000} /* (8, 0, 25) {real, imag} */,
  {32'h3f79207d, 32'h00000000} /* (8, 0, 24) {real, imag} */,
  {32'h3e7eb421, 32'h00000000} /* (8, 0, 23) {real, imag} */,
  {32'h3df561ab, 32'h00000000} /* (8, 0, 22) {real, imag} */,
  {32'h3e8dbaa0, 32'h00000000} /* (8, 0, 21) {real, imag} */,
  {32'h3e6ee694, 32'h00000000} /* (8, 0, 20) {real, imag} */,
  {32'h3f0d936c, 32'h00000000} /* (8, 0, 19) {real, imag} */,
  {32'h3f529294, 32'h00000000} /* (8, 0, 18) {real, imag} */,
  {32'h3f1c9964, 32'h00000000} /* (8, 0, 17) {real, imag} */,
  {32'h3ec87e4e, 32'h00000000} /* (8, 0, 16) {real, imag} */,
  {32'hbdc1f97b, 32'h00000000} /* (8, 0, 15) {real, imag} */,
  {32'hbf515984, 32'h00000000} /* (8, 0, 14) {real, imag} */,
  {32'hbf18f7a8, 32'h00000000} /* (8, 0, 13) {real, imag} */,
  {32'hbf29c1e8, 32'h00000000} /* (8, 0, 12) {real, imag} */,
  {32'hbf14e1bf, 32'h00000000} /* (8, 0, 11) {real, imag} */,
  {32'hbf1c4698, 32'h00000000} /* (8, 0, 10) {real, imag} */,
  {32'hbf7a1a82, 32'h00000000} /* (8, 0, 9) {real, imag} */,
  {32'hbf52cf9a, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'hbf22a95e, 32'h00000000} /* (8, 0, 7) {real, imag} */,
  {32'hbe61ef7c, 32'h00000000} /* (8, 0, 6) {real, imag} */,
  {32'hbc96c97a, 32'h00000000} /* (8, 0, 5) {real, imag} */,
  {32'h3e8e93e5, 32'h00000000} /* (8, 0, 4) {real, imag} */,
  {32'h3f4e3dbe, 32'h00000000} /* (8, 0, 3) {real, imag} */,
  {32'h3f03045c, 32'h00000000} /* (8, 0, 2) {real, imag} */,
  {32'h3e99b3a5, 32'h00000000} /* (8, 0, 1) {real, imag} */,
  {32'h3e10e319, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h3e9322cb, 32'h00000000} /* (7, 31, 31) {real, imag} */,
  {32'h3f076027, 32'h00000000} /* (7, 31, 30) {real, imag} */,
  {32'h3f28924a, 32'h00000000} /* (7, 31, 29) {real, imag} */,
  {32'h3f1d1b20, 32'h00000000} /* (7, 31, 28) {real, imag} */,
  {32'h3f15c73c, 32'h00000000} /* (7, 31, 27) {real, imag} */,
  {32'h3f25cdf7, 32'h00000000} /* (7, 31, 26) {real, imag} */,
  {32'h3f3d5693, 32'h00000000} /* (7, 31, 25) {real, imag} */,
  {32'h3ee6a2a9, 32'h00000000} /* (7, 31, 24) {real, imag} */,
  {32'h3f0d8607, 32'h00000000} /* (7, 31, 23) {real, imag} */,
  {32'h3ef4a3d2, 32'h00000000} /* (7, 31, 22) {real, imag} */,
  {32'hbc3a2180, 32'h00000000} /* (7, 31, 21) {real, imag} */,
  {32'hbf35b99f, 32'h00000000} /* (7, 31, 20) {real, imag} */,
  {32'hbeee95ee, 32'h00000000} /* (7, 31, 19) {real, imag} */,
  {32'hbe9cd266, 32'h00000000} /* (7, 31, 18) {real, imag} */,
  {32'hbe904861, 32'h00000000} /* (7, 31, 17) {real, imag} */,
  {32'hbeefc9a1, 32'h00000000} /* (7, 31, 16) {real, imag} */,
  {32'hbeb2f0cb, 32'h00000000} /* (7, 31, 15) {real, imag} */,
  {32'hbed363ba, 32'h00000000} /* (7, 31, 14) {real, imag} */,
  {32'hbebddef0, 32'h00000000} /* (7, 31, 13) {real, imag} */,
  {32'hbf667f7d, 32'h00000000} /* (7, 31, 12) {real, imag} */,
  {32'hbf332a10, 32'h00000000} /* (7, 31, 11) {real, imag} */,
  {32'h3f2eaacc, 32'h00000000} /* (7, 31, 10) {real, imag} */,
  {32'h3e891882, 32'h00000000} /* (7, 31, 9) {real, imag} */,
  {32'h3e395c08, 32'h00000000} /* (7, 31, 8) {real, imag} */,
  {32'h3f6388a0, 32'h00000000} /* (7, 31, 7) {real, imag} */,
  {32'h3f25512a, 32'h00000000} /* (7, 31, 6) {real, imag} */,
  {32'h3ebeef34, 32'h00000000} /* (7, 31, 5) {real, imag} */,
  {32'h3eae35b0, 32'h00000000} /* (7, 31, 4) {real, imag} */,
  {32'h3f03b01a, 32'h00000000} /* (7, 31, 3) {real, imag} */,
  {32'h3f0b27db, 32'h00000000} /* (7, 31, 2) {real, imag} */,
  {32'h3f4ac339, 32'h00000000} /* (7, 31, 1) {real, imag} */,
  {32'h3eaeeadc, 32'h00000000} /* (7, 31, 0) {real, imag} */,
  {32'h3ed1fdb2, 32'h00000000} /* (7, 30, 31) {real, imag} */,
  {32'h3f5e985e, 32'h00000000} /* (7, 30, 30) {real, imag} */,
  {32'h3f8d63bc, 32'h00000000} /* (7, 30, 29) {real, imag} */,
  {32'h3f96ddce, 32'h00000000} /* (7, 30, 28) {real, imag} */,
  {32'h3f5106b4, 32'h00000000} /* (7, 30, 27) {real, imag} */,
  {32'h3f12e556, 32'h00000000} /* (7, 30, 26) {real, imag} */,
  {32'h3f307ae8, 32'h00000000} /* (7, 30, 25) {real, imag} */,
  {32'h3f330cab, 32'h00000000} /* (7, 30, 24) {real, imag} */,
  {32'h3f9a92c8, 32'h00000000} /* (7, 30, 23) {real, imag} */,
  {32'h3fa6879d, 32'h00000000} /* (7, 30, 22) {real, imag} */,
  {32'h3d4f9553, 32'h00000000} /* (7, 30, 21) {real, imag} */,
  {32'hbff2a275, 32'h00000000} /* (7, 30, 20) {real, imag} */,
  {32'hbfbf3b90, 32'h00000000} /* (7, 30, 19) {real, imag} */,
  {32'hbf9243ff, 32'h00000000} /* (7, 30, 18) {real, imag} */,
  {32'hbf8b0a38, 32'h00000000} /* (7, 30, 17) {real, imag} */,
  {32'hbfa7385c, 32'h00000000} /* (7, 30, 16) {real, imag} */,
  {32'hbf838d2c, 32'h00000000} /* (7, 30, 15) {real, imag} */,
  {32'hbf8ee641, 32'h00000000} /* (7, 30, 14) {real, imag} */,
  {32'hbf654f67, 32'h00000000} /* (7, 30, 13) {real, imag} */,
  {32'hbf8c2e31, 32'h00000000} /* (7, 30, 12) {real, imag} */,
  {32'hbf8b65c4, 32'h00000000} /* (7, 30, 11) {real, imag} */,
  {32'h3ea073be, 32'h00000000} /* (7, 30, 10) {real, imag} */,
  {32'h3ecdccc0, 32'h00000000} /* (7, 30, 9) {real, imag} */,
  {32'h3f3c2962, 32'h00000000} /* (7, 30, 8) {real, imag} */,
  {32'h3f7f14db, 32'h00000000} /* (7, 30, 7) {real, imag} */,
  {32'h3f847472, 32'h00000000} /* (7, 30, 6) {real, imag} */,
  {32'h3f9cb5d9, 32'h00000000} /* (7, 30, 5) {real, imag} */,
  {32'h3f9dc30a, 32'h00000000} /* (7, 30, 4) {real, imag} */,
  {32'h3f66aa39, 32'h00000000} /* (7, 30, 3) {real, imag} */,
  {32'h3fc29a0e, 32'h00000000} /* (7, 30, 2) {real, imag} */,
  {32'h3fb2455d, 32'h00000000} /* (7, 30, 1) {real, imag} */,
  {32'h3ec7ef94, 32'h00000000} /* (7, 30, 0) {real, imag} */,
  {32'h3eef3b56, 32'h00000000} /* (7, 29, 31) {real, imag} */,
  {32'h3f41beb7, 32'h00000000} /* (7, 29, 30) {real, imag} */,
  {32'h3f452240, 32'h00000000} /* (7, 29, 29) {real, imag} */,
  {32'h3f5d848a, 32'h00000000} /* (7, 29, 28) {real, imag} */,
  {32'h3efde8ff, 32'h00000000} /* (7, 29, 27) {real, imag} */,
  {32'h3ef8e61c, 32'h00000000} /* (7, 29, 26) {real, imag} */,
  {32'h3ee4fb84, 32'h00000000} /* (7, 29, 25) {real, imag} */,
  {32'h3eb2c046, 32'h00000000} /* (7, 29, 24) {real, imag} */,
  {32'h3f0214ad, 32'h00000000} /* (7, 29, 23) {real, imag} */,
  {32'h3f32a026, 32'h00000000} /* (7, 29, 22) {real, imag} */,
  {32'h3e8a78ac, 32'h00000000} /* (7, 29, 21) {real, imag} */,
  {32'hbff66418, 32'h00000000} /* (7, 29, 20) {real, imag} */,
  {32'hbfadd218, 32'h00000000} /* (7, 29, 19) {real, imag} */,
  {32'hbf8801af, 32'h00000000} /* (7, 29, 18) {real, imag} */,
  {32'hbf756c1d, 32'h00000000} /* (7, 29, 17) {real, imag} */,
  {32'hbf5a114b, 32'h00000000} /* (7, 29, 16) {real, imag} */,
  {32'hbf78b94d, 32'h00000000} /* (7, 29, 15) {real, imag} */,
  {32'hbf8d4eac, 32'h00000000} /* (7, 29, 14) {real, imag} */,
  {32'hbf83fc1b, 32'h00000000} /* (7, 29, 13) {real, imag} */,
  {32'hbf726034, 32'h00000000} /* (7, 29, 12) {real, imag} */,
  {32'hbf7436ba, 32'h00000000} /* (7, 29, 11) {real, imag} */,
  {32'h3e99a11e, 32'h00000000} /* (7, 29, 10) {real, imag} */,
  {32'h3f7d5485, 32'h00000000} /* (7, 29, 9) {real, imag} */,
  {32'h3f968f22, 32'h00000000} /* (7, 29, 8) {real, imag} */,
  {32'h3f7ee61b, 32'h00000000} /* (7, 29, 7) {real, imag} */,
  {32'h3f91b82c, 32'h00000000} /* (7, 29, 6) {real, imag} */,
  {32'h3fcede75, 32'h00000000} /* (7, 29, 5) {real, imag} */,
  {32'h3fb6af5a, 32'h00000000} /* (7, 29, 4) {real, imag} */,
  {32'h3faaaeaf, 32'h00000000} /* (7, 29, 3) {real, imag} */,
  {32'h3fd054a6, 32'h00000000} /* (7, 29, 2) {real, imag} */,
  {32'h3f979efd, 32'h00000000} /* (7, 29, 1) {real, imag} */,
  {32'h3f06c561, 32'h00000000} /* (7, 29, 0) {real, imag} */,
  {32'h3efbb180, 32'h00000000} /* (7, 28, 31) {real, imag} */,
  {32'h3f329eab, 32'h00000000} /* (7, 28, 30) {real, imag} */,
  {32'h3f633296, 32'h00000000} /* (7, 28, 29) {real, imag} */,
  {32'h3f8ccef8, 32'h00000000} /* (7, 28, 28) {real, imag} */,
  {32'h3e94f38c, 32'h00000000} /* (7, 28, 27) {real, imag} */,
  {32'h3eb3d8bc, 32'h00000000} /* (7, 28, 26) {real, imag} */,
  {32'h3eb9d9d0, 32'h00000000} /* (7, 28, 25) {real, imag} */,
  {32'h3f0f3f9d, 32'h00000000} /* (7, 28, 24) {real, imag} */,
  {32'h3f150dad, 32'h00000000} /* (7, 28, 23) {real, imag} */,
  {32'h3ef722f4, 32'h00000000} /* (7, 28, 22) {real, imag} */,
  {32'h3ed54ac4, 32'h00000000} /* (7, 28, 21) {real, imag} */,
  {32'hbf3545bd, 32'h00000000} /* (7, 28, 20) {real, imag} */,
  {32'hbf0e6702, 32'h00000000} /* (7, 28, 19) {real, imag} */,
  {32'hbf4a1afe, 32'h00000000} /* (7, 28, 18) {real, imag} */,
  {32'hbf39f18b, 32'h00000000} /* (7, 28, 17) {real, imag} */,
  {32'hbedb0d17, 32'h00000000} /* (7, 28, 16) {real, imag} */,
  {32'hbf38edc8, 32'h00000000} /* (7, 28, 15) {real, imag} */,
  {32'hbf791000, 32'h00000000} /* (7, 28, 14) {real, imag} */,
  {32'hbf64a64f, 32'h00000000} /* (7, 28, 13) {real, imag} */,
  {32'hbf1fa03e, 32'h00000000} /* (7, 28, 12) {real, imag} */,
  {32'hbf466efd, 32'h00000000} /* (7, 28, 11) {real, imag} */,
  {32'h3de6b5ec, 32'h00000000} /* (7, 28, 10) {real, imag} */,
  {32'h3f6b3b30, 32'h00000000} /* (7, 28, 9) {real, imag} */,
  {32'h3f751ed2, 32'h00000000} /* (7, 28, 8) {real, imag} */,
  {32'h3fa99712, 32'h00000000} /* (7, 28, 7) {real, imag} */,
  {32'h3f62370c, 32'h00000000} /* (7, 28, 6) {real, imag} */,
  {32'h3f921424, 32'h00000000} /* (7, 28, 5) {real, imag} */,
  {32'h3f9b3251, 32'h00000000} /* (7, 28, 4) {real, imag} */,
  {32'h3fa765be, 32'h00000000} /* (7, 28, 3) {real, imag} */,
  {32'h3f720c02, 32'h00000000} /* (7, 28, 2) {real, imag} */,
  {32'h3eadd88b, 32'h00000000} /* (7, 28, 1) {real, imag} */,
  {32'h3e86dd7f, 32'h00000000} /* (7, 28, 0) {real, imag} */,
  {32'h3f40b7b1, 32'h00000000} /* (7, 27, 31) {real, imag} */,
  {32'h3f12ce73, 32'h00000000} /* (7, 27, 30) {real, imag} */,
  {32'h3f2cca2e, 32'h00000000} /* (7, 27, 29) {real, imag} */,
  {32'h3f895032, 32'h00000000} /* (7, 27, 28) {real, imag} */,
  {32'h3f236174, 32'h00000000} /* (7, 27, 27) {real, imag} */,
  {32'h3f2e41b5, 32'h00000000} /* (7, 27, 26) {real, imag} */,
  {32'h3ed51dd9, 32'h00000000} /* (7, 27, 25) {real, imag} */,
  {32'h3f8ee11b, 32'h00000000} /* (7, 27, 24) {real, imag} */,
  {32'h3f93f553, 32'h00000000} /* (7, 27, 23) {real, imag} */,
  {32'h3f49b2a8, 32'h00000000} /* (7, 27, 22) {real, imag} */,
  {32'h3f018c64, 32'h00000000} /* (7, 27, 21) {real, imag} */,
  {32'hbf42f428, 32'h00000000} /* (7, 27, 20) {real, imag} */,
  {32'hbf596e01, 32'h00000000} /* (7, 27, 19) {real, imag} */,
  {32'hbf6a11a6, 32'h00000000} /* (7, 27, 18) {real, imag} */,
  {32'hbf83ce8c, 32'h00000000} /* (7, 27, 17) {real, imag} */,
  {32'hbf89b171, 32'h00000000} /* (7, 27, 16) {real, imag} */,
  {32'hbf6514ad, 32'h00000000} /* (7, 27, 15) {real, imag} */,
  {32'hbf599c79, 32'h00000000} /* (7, 27, 14) {real, imag} */,
  {32'hbf7c1338, 32'h00000000} /* (7, 27, 13) {real, imag} */,
  {32'hbf7a054f, 32'h00000000} /* (7, 27, 12) {real, imag} */,
  {32'hbf80c4c3, 32'h00000000} /* (7, 27, 11) {real, imag} */,
  {32'h3e1c12ee, 32'h00000000} /* (7, 27, 10) {real, imag} */,
  {32'h3f4afb39, 32'h00000000} /* (7, 27, 9) {real, imag} */,
  {32'h3f4c8e2d, 32'h00000000} /* (7, 27, 8) {real, imag} */,
  {32'h3f90276d, 32'h00000000} /* (7, 27, 7) {real, imag} */,
  {32'h3f129cca, 32'h00000000} /* (7, 27, 6) {real, imag} */,
  {32'h3f70c002, 32'h00000000} /* (7, 27, 5) {real, imag} */,
  {32'h3f9d3e1d, 32'h00000000} /* (7, 27, 4) {real, imag} */,
  {32'h3f6b9687, 32'h00000000} /* (7, 27, 3) {real, imag} */,
  {32'h3ed4e758, 32'h00000000} /* (7, 27, 2) {real, imag} */,
  {32'h3f055a5f, 32'h00000000} /* (7, 27, 1) {real, imag} */,
  {32'h3f2377e4, 32'h00000000} /* (7, 27, 0) {real, imag} */,
  {32'h3eefa3d0, 32'h00000000} /* (7, 26, 31) {real, imag} */,
  {32'h3ed91870, 32'h00000000} /* (7, 26, 30) {real, imag} */,
  {32'h3f8c4c6a, 32'h00000000} /* (7, 26, 29) {real, imag} */,
  {32'h3fa496f1, 32'h00000000} /* (7, 26, 28) {real, imag} */,
  {32'h3f8dc525, 32'h00000000} /* (7, 26, 27) {real, imag} */,
  {32'h3f9c8e2a, 32'h00000000} /* (7, 26, 26) {real, imag} */,
  {32'h3f809210, 32'h00000000} /* (7, 26, 25) {real, imag} */,
  {32'h3f7edc7f, 32'h00000000} /* (7, 26, 24) {real, imag} */,
  {32'h3f755b80, 32'h00000000} /* (7, 26, 23) {real, imag} */,
  {32'h3f773281, 32'h00000000} /* (7, 26, 22) {real, imag} */,
  {32'h3f16090d, 32'h00000000} /* (7, 26, 21) {real, imag} */,
  {32'hbf23a784, 32'h00000000} /* (7, 26, 20) {real, imag} */,
  {32'hbf82cef1, 32'h00000000} /* (7, 26, 19) {real, imag} */,
  {32'hbf4323db, 32'h00000000} /* (7, 26, 18) {real, imag} */,
  {32'hbf6547ab, 32'h00000000} /* (7, 26, 17) {real, imag} */,
  {32'hbfa5becd, 32'h00000000} /* (7, 26, 16) {real, imag} */,
  {32'hbf90cdd1, 32'h00000000} /* (7, 26, 15) {real, imag} */,
  {32'hbfb52742, 32'h00000000} /* (7, 26, 14) {real, imag} */,
  {32'hbfa0bf86, 32'h00000000} /* (7, 26, 13) {real, imag} */,
  {32'hbf502b34, 32'h00000000} /* (7, 26, 12) {real, imag} */,
  {32'hbf17a6ef, 32'h00000000} /* (7, 26, 11) {real, imag} */,
  {32'h3f017f27, 32'h00000000} /* (7, 26, 10) {real, imag} */,
  {32'h3f902e24, 32'h00000000} /* (7, 26, 9) {real, imag} */,
  {32'h3f5ee64c, 32'h00000000} /* (7, 26, 8) {real, imag} */,
  {32'h3f2720b9, 32'h00000000} /* (7, 26, 7) {real, imag} */,
  {32'h3e4eac49, 32'h00000000} /* (7, 26, 6) {real, imag} */,
  {32'h3f184950, 32'h00000000} /* (7, 26, 5) {real, imag} */,
  {32'h3f610039, 32'h00000000} /* (7, 26, 4) {real, imag} */,
  {32'h3f139541, 32'h00000000} /* (7, 26, 3) {real, imag} */,
  {32'h3e99824b, 32'h00000000} /* (7, 26, 2) {real, imag} */,
  {32'h3f402766, 32'h00000000} /* (7, 26, 1) {real, imag} */,
  {32'h3f3c749b, 32'h00000000} /* (7, 26, 0) {real, imag} */,
  {32'h3f39d0b8, 32'h00000000} /* (7, 25, 31) {real, imag} */,
  {32'h3f5508d4, 32'h00000000} /* (7, 25, 30) {real, imag} */,
  {32'h3f50ecf7, 32'h00000000} /* (7, 25, 29) {real, imag} */,
  {32'h3f7e36bf, 32'h00000000} /* (7, 25, 28) {real, imag} */,
  {32'h3fa1db79, 32'h00000000} /* (7, 25, 27) {real, imag} */,
  {32'h3fb5343a, 32'h00000000} /* (7, 25, 26) {real, imag} */,
  {32'h3f8cf499, 32'h00000000} /* (7, 25, 25) {real, imag} */,
  {32'h3f851dcb, 32'h00000000} /* (7, 25, 24) {real, imag} */,
  {32'h3f905bf7, 32'h00000000} /* (7, 25, 23) {real, imag} */,
  {32'h3f8ef52a, 32'h00000000} /* (7, 25, 22) {real, imag} */,
  {32'h3f176747, 32'h00000000} /* (7, 25, 21) {real, imag} */,
  {32'hbeecdb40, 32'h00000000} /* (7, 25, 20) {real, imag} */,
  {32'hbf9dd1a1, 32'h00000000} /* (7, 25, 19) {real, imag} */,
  {32'hbf54ccf0, 32'h00000000} /* (7, 25, 18) {real, imag} */,
  {32'hbf62a479, 32'h00000000} /* (7, 25, 17) {real, imag} */,
  {32'hbf79800e, 32'h00000000} /* (7, 25, 16) {real, imag} */,
  {32'hbf8d9f01, 32'h00000000} /* (7, 25, 15) {real, imag} */,
  {32'hbfcdc9bb, 32'h00000000} /* (7, 25, 14) {real, imag} */,
  {32'hbf8c4017, 32'h00000000} /* (7, 25, 13) {real, imag} */,
  {32'hbf938dbc, 32'h00000000} /* (7, 25, 12) {real, imag} */,
  {32'hbf5990db, 32'h00000000} /* (7, 25, 11) {real, imag} */,
  {32'h3edd6789, 32'h00000000} /* (7, 25, 10) {real, imag} */,
  {32'h3f8bd547, 32'h00000000} /* (7, 25, 9) {real, imag} */,
  {32'h3f92b9a8, 32'h00000000} /* (7, 25, 8) {real, imag} */,
  {32'h3f51816e, 32'h00000000} /* (7, 25, 7) {real, imag} */,
  {32'h3eb24bfb, 32'h00000000} /* (7, 25, 6) {real, imag} */,
  {32'h3f022eb0, 32'h00000000} /* (7, 25, 5) {real, imag} */,
  {32'h3f263edc, 32'h00000000} /* (7, 25, 4) {real, imag} */,
  {32'h3f28da78, 32'h00000000} /* (7, 25, 3) {real, imag} */,
  {32'h3f1790ac, 32'h00000000} /* (7, 25, 2) {real, imag} */,
  {32'h3f06cdb2, 32'h00000000} /* (7, 25, 1) {real, imag} */,
  {32'h3e961559, 32'h00000000} /* (7, 25, 0) {real, imag} */,
  {32'h3f2e6b01, 32'h00000000} /* (7, 24, 31) {real, imag} */,
  {32'h3f857ae8, 32'h00000000} /* (7, 24, 30) {real, imag} */,
  {32'h3f1da62d, 32'h00000000} /* (7, 24, 29) {real, imag} */,
  {32'h3f92ff87, 32'h00000000} /* (7, 24, 28) {real, imag} */,
  {32'h3fbad0d1, 32'h00000000} /* (7, 24, 27) {real, imag} */,
  {32'h3fa43b60, 32'h00000000} /* (7, 24, 26) {real, imag} */,
  {32'h3fb78b09, 32'h00000000} /* (7, 24, 25) {real, imag} */,
  {32'h3fa5b059, 32'h00000000} /* (7, 24, 24) {real, imag} */,
  {32'h3fae1b80, 32'h00000000} /* (7, 24, 23) {real, imag} */,
  {32'h3fbec235, 32'h00000000} /* (7, 24, 22) {real, imag} */,
  {32'h3f337a0d, 32'h00000000} /* (7, 24, 21) {real, imag} */,
  {32'hbf26b135, 32'h00000000} /* (7, 24, 20) {real, imag} */,
  {32'hbf58d96e, 32'h00000000} /* (7, 24, 19) {real, imag} */,
  {32'hbf494438, 32'h00000000} /* (7, 24, 18) {real, imag} */,
  {32'hbf866fac, 32'h00000000} /* (7, 24, 17) {real, imag} */,
  {32'hbf95b823, 32'h00000000} /* (7, 24, 16) {real, imag} */,
  {32'hbfa9e8a2, 32'h00000000} /* (7, 24, 15) {real, imag} */,
  {32'hbfa366a4, 32'h00000000} /* (7, 24, 14) {real, imag} */,
  {32'hbfe12cc5, 32'h00000000} /* (7, 24, 13) {real, imag} */,
  {32'hbf9fe88d, 32'h00000000} /* (7, 24, 12) {real, imag} */,
  {32'hbf27b3e9, 32'h00000000} /* (7, 24, 11) {real, imag} */,
  {32'h3e4c80b4, 32'h00000000} /* (7, 24, 10) {real, imag} */,
  {32'h3fa18f09, 32'h00000000} /* (7, 24, 9) {real, imag} */,
  {32'h3f85efe6, 32'h00000000} /* (7, 24, 8) {real, imag} */,
  {32'h3f4ab441, 32'h00000000} /* (7, 24, 7) {real, imag} */,
  {32'h3f4106dc, 32'h00000000} /* (7, 24, 6) {real, imag} */,
  {32'h3f2866ce, 32'h00000000} /* (7, 24, 5) {real, imag} */,
  {32'h3f3444ba, 32'h00000000} /* (7, 24, 4) {real, imag} */,
  {32'h3f86dff5, 32'h00000000} /* (7, 24, 3) {real, imag} */,
  {32'h3f916374, 32'h00000000} /* (7, 24, 2) {real, imag} */,
  {32'h3f148b15, 32'h00000000} /* (7, 24, 1) {real, imag} */,
  {32'h3e764d46, 32'h00000000} /* (7, 24, 0) {real, imag} */,
  {32'h3efd9742, 32'h00000000} /* (7, 23, 31) {real, imag} */,
  {32'h3f86deb9, 32'h00000000} /* (7, 23, 30) {real, imag} */,
  {32'h3f65efe0, 32'h00000000} /* (7, 23, 29) {real, imag} */,
  {32'h3f8a70c8, 32'h00000000} /* (7, 23, 28) {real, imag} */,
  {32'h3fd8c2c8, 32'h00000000} /* (7, 23, 27) {real, imag} */,
  {32'h3fb486d7, 32'h00000000} /* (7, 23, 26) {real, imag} */,
  {32'h3f8efc27, 32'h00000000} /* (7, 23, 25) {real, imag} */,
  {32'h3f59510c, 32'h00000000} /* (7, 23, 24) {real, imag} */,
  {32'h3f9719d2, 32'h00000000} /* (7, 23, 23) {real, imag} */,
  {32'h3f99769c, 32'h00000000} /* (7, 23, 22) {real, imag} */,
  {32'h3f134de3, 32'h00000000} /* (7, 23, 21) {real, imag} */,
  {32'hbed3052d, 32'h00000000} /* (7, 23, 20) {real, imag} */,
  {32'hbf179473, 32'h00000000} /* (7, 23, 19) {real, imag} */,
  {32'hbf00b57b, 32'h00000000} /* (7, 23, 18) {real, imag} */,
  {32'hbf3eea8c, 32'h00000000} /* (7, 23, 17) {real, imag} */,
  {32'hbf5eba69, 32'h00000000} /* (7, 23, 16) {real, imag} */,
  {32'hbf3ccd97, 32'h00000000} /* (7, 23, 15) {real, imag} */,
  {32'hbf98216c, 32'h00000000} /* (7, 23, 14) {real, imag} */,
  {32'hbfe0de01, 32'h00000000} /* (7, 23, 13) {real, imag} */,
  {32'hbf903f17, 32'h00000000} /* (7, 23, 12) {real, imag} */,
  {32'hbf09d167, 32'h00000000} /* (7, 23, 11) {real, imag} */,
  {32'h3ce0efe5, 32'h00000000} /* (7, 23, 10) {real, imag} */,
  {32'h3f5dd33b, 32'h00000000} /* (7, 23, 9) {real, imag} */,
  {32'h3f910f13, 32'h00000000} /* (7, 23, 8) {real, imag} */,
  {32'h3f987cab, 32'h00000000} /* (7, 23, 7) {real, imag} */,
  {32'h3faaa108, 32'h00000000} /* (7, 23, 6) {real, imag} */,
  {32'h3f98aa68, 32'h00000000} /* (7, 23, 5) {real, imag} */,
  {32'h3f35ea31, 32'h00000000} /* (7, 23, 4) {real, imag} */,
  {32'h3f3c046c, 32'h00000000} /* (7, 23, 3) {real, imag} */,
  {32'h3f4d9b86, 32'h00000000} /* (7, 23, 2) {real, imag} */,
  {32'h3ec108ec, 32'h00000000} /* (7, 23, 1) {real, imag} */,
  {32'h3e587f5d, 32'h00000000} /* (7, 23, 0) {real, imag} */,
  {32'h3e4653e8, 32'h00000000} /* (7, 22, 31) {real, imag} */,
  {32'h3ef37bb1, 32'h00000000} /* (7, 22, 30) {real, imag} */,
  {32'h3f590779, 32'h00000000} /* (7, 22, 29) {real, imag} */,
  {32'h3f912df2, 32'h00000000} /* (7, 22, 28) {real, imag} */,
  {32'h3fe4792a, 32'h00000000} /* (7, 22, 27) {real, imag} */,
  {32'h3f9ccaff, 32'h00000000} /* (7, 22, 26) {real, imag} */,
  {32'h3f847921, 32'h00000000} /* (7, 22, 25) {real, imag} */,
  {32'h3f474379, 32'h00000000} /* (7, 22, 24) {real, imag} */,
  {32'h3faeb0bc, 32'h00000000} /* (7, 22, 23) {real, imag} */,
  {32'h3fb6716e, 32'h00000000} /* (7, 22, 22) {real, imag} */,
  {32'h3f079832, 32'h00000000} /* (7, 22, 21) {real, imag} */,
  {32'hbee629b1, 32'h00000000} /* (7, 22, 20) {real, imag} */,
  {32'hbf44359a, 32'h00000000} /* (7, 22, 19) {real, imag} */,
  {32'hbe8d56af, 32'h00000000} /* (7, 22, 18) {real, imag} */,
  {32'hbf104321, 32'h00000000} /* (7, 22, 17) {real, imag} */,
  {32'hbf7509fe, 32'h00000000} /* (7, 22, 16) {real, imag} */,
  {32'hbf2acd73, 32'h00000000} /* (7, 22, 15) {real, imag} */,
  {32'hbf8e0516, 32'h00000000} /* (7, 22, 14) {real, imag} */,
  {32'hbf983e5e, 32'h00000000} /* (7, 22, 13) {real, imag} */,
  {32'hbfb5a69c, 32'h00000000} /* (7, 22, 12) {real, imag} */,
  {32'hbf4e4f09, 32'h00000000} /* (7, 22, 11) {real, imag} */,
  {32'h3f0378ba, 32'h00000000} /* (7, 22, 10) {real, imag} */,
  {32'h3f8e40e4, 32'h00000000} /* (7, 22, 9) {real, imag} */,
  {32'h3fdff0e8, 32'h00000000} /* (7, 22, 8) {real, imag} */,
  {32'h3fd001bf, 32'h00000000} /* (7, 22, 7) {real, imag} */,
  {32'h3fa071f4, 32'h00000000} /* (7, 22, 6) {real, imag} */,
  {32'h3f960c7f, 32'h00000000} /* (7, 22, 5) {real, imag} */,
  {32'h3ef40208, 32'h00000000} /* (7, 22, 4) {real, imag} */,
  {32'h3f253580, 32'h00000000} /* (7, 22, 3) {real, imag} */,
  {32'h3f462489, 32'h00000000} /* (7, 22, 2) {real, imag} */,
  {32'h3e8a6807, 32'h00000000} /* (7, 22, 1) {real, imag} */,
  {32'h3dc266fa, 32'h00000000} /* (7, 22, 0) {real, imag} */,
  {32'h3e566be6, 32'h00000000} /* (7, 21, 31) {real, imag} */,
  {32'h3f18f3f9, 32'h00000000} /* (7, 21, 30) {real, imag} */,
  {32'h3ef2bead, 32'h00000000} /* (7, 21, 29) {real, imag} */,
  {32'h3f68f3e2, 32'h00000000} /* (7, 21, 28) {real, imag} */,
  {32'h3fc5e2e6, 32'h00000000} /* (7, 21, 27) {real, imag} */,
  {32'h3f401bc4, 32'h00000000} /* (7, 21, 26) {real, imag} */,
  {32'h3f21c46c, 32'h00000000} /* (7, 21, 25) {real, imag} */,
  {32'h3e2c5e74, 32'h00000000} /* (7, 21, 24) {real, imag} */,
  {32'h3f02fd1c, 32'h00000000} /* (7, 21, 23) {real, imag} */,
  {32'h3e9830ae, 32'h00000000} /* (7, 21, 22) {real, imag} */,
  {32'hbdcd1d3a, 32'h00000000} /* (7, 21, 21) {real, imag} */,
  {32'hbf40d7a9, 32'h00000000} /* (7, 21, 20) {real, imag} */,
  {32'hbf028964, 32'h00000000} /* (7, 21, 19) {real, imag} */,
  {32'hbdbe6ec7, 32'h00000000} /* (7, 21, 18) {real, imag} */,
  {32'hbe710434, 32'h00000000} /* (7, 21, 17) {real, imag} */,
  {32'hbe64776e, 32'h00000000} /* (7, 21, 16) {real, imag} */,
  {32'hbea98ea6, 32'h00000000} /* (7, 21, 15) {real, imag} */,
  {32'hbed31d61, 32'h00000000} /* (7, 21, 14) {real, imag} */,
  {32'hbe670e76, 32'h00000000} /* (7, 21, 13) {real, imag} */,
  {32'hbf0cde22, 32'h00000000} /* (7, 21, 12) {real, imag} */,
  {32'hbe38e4b9, 32'h00000000} /* (7, 21, 11) {real, imag} */,
  {32'h3f0ba204, 32'h00000000} /* (7, 21, 10) {real, imag} */,
  {32'h3f44557d, 32'h00000000} /* (7, 21, 9) {real, imag} */,
  {32'h3f73763e, 32'h00000000} /* (7, 21, 8) {real, imag} */,
  {32'h3f49bbbf, 32'h00000000} /* (7, 21, 7) {real, imag} */,
  {32'h3e00b8fd, 32'h00000000} /* (7, 21, 6) {real, imag} */,
  {32'hbdb9952b, 32'h00000000} /* (7, 21, 5) {real, imag} */,
  {32'hbd010149, 32'h00000000} /* (7, 21, 4) {real, imag} */,
  {32'h3e863f0b, 32'h00000000} /* (7, 21, 3) {real, imag} */,
  {32'h3ec91544, 32'h00000000} /* (7, 21, 2) {real, imag} */,
  {32'h3e6daa18, 32'h00000000} /* (7, 21, 1) {real, imag} */,
  {32'h3de4bab1, 32'h00000000} /* (7, 21, 0) {real, imag} */,
  {32'hbe182946, 32'h00000000} /* (7, 20, 31) {real, imag} */,
  {32'hbe962616, 32'h00000000} /* (7, 20, 30) {real, imag} */,
  {32'hbf388832, 32'h00000000} /* (7, 20, 29) {real, imag} */,
  {32'hbe74fdd2, 32'h00000000} /* (7, 20, 28) {real, imag} */,
  {32'h3cae5fa0, 32'h00000000} /* (7, 20, 27) {real, imag} */,
  {32'hbec42262, 32'h00000000} /* (7, 20, 26) {real, imag} */,
  {32'hbeeb4097, 32'h00000000} /* (7, 20, 25) {real, imag} */,
  {32'hbf4646d8, 32'h00000000} /* (7, 20, 24) {real, imag} */,
  {32'hbfa6e176, 32'h00000000} /* (7, 20, 23) {real, imag} */,
  {32'hbfb9ea64, 32'h00000000} /* (7, 20, 22) {real, imag} */,
  {32'hbf249436, 32'h00000000} /* (7, 20, 21) {real, imag} */,
  {32'hbe1eb641, 32'h00000000} /* (7, 20, 20) {real, imag} */,
  {32'h3ed41024, 32'h00000000} /* (7, 20, 19) {real, imag} */,
  {32'h3f6fb947, 32'h00000000} /* (7, 20, 18) {real, imag} */,
  {32'h3f575abe, 32'h00000000} /* (7, 20, 17) {real, imag} */,
  {32'h3ef6ba76, 32'h00000000} /* (7, 20, 16) {real, imag} */,
  {32'h3ed7f56f, 32'h00000000} /* (7, 20, 15) {real, imag} */,
  {32'h3f4f6409, 32'h00000000} /* (7, 20, 14) {real, imag} */,
  {32'h3f2e25e1, 32'h00000000} /* (7, 20, 13) {real, imag} */,
  {32'h3f10340a, 32'h00000000} /* (7, 20, 12) {real, imag} */,
  {32'h3eb86bfd, 32'h00000000} /* (7, 20, 11) {real, imag} */,
  {32'hbed67d66, 32'h00000000} /* (7, 20, 10) {real, imag} */,
  {32'hbf3796f0, 32'h00000000} /* (7, 20, 9) {real, imag} */,
  {32'hbf813241, 32'h00000000} /* (7, 20, 8) {real, imag} */,
  {32'hbf60a89a, 32'h00000000} /* (7, 20, 7) {real, imag} */,
  {32'hbf82aa5e, 32'h00000000} /* (7, 20, 6) {real, imag} */,
  {32'hbf4942cb, 32'h00000000} /* (7, 20, 5) {real, imag} */,
  {32'hbf71d8a0, 32'h00000000} /* (7, 20, 4) {real, imag} */,
  {32'hbf922062, 32'h00000000} /* (7, 20, 3) {real, imag} */,
  {32'hbf5d2ca2, 32'h00000000} /* (7, 20, 2) {real, imag} */,
  {32'hbf70ba90, 32'h00000000} /* (7, 20, 1) {real, imag} */,
  {32'hbec2b95a, 32'h00000000} /* (7, 20, 0) {real, imag} */,
  {32'hbe6b690d, 32'h00000000} /* (7, 19, 31) {real, imag} */,
  {32'hbec034b9, 32'h00000000} /* (7, 19, 30) {real, imag} */,
  {32'hbf145461, 32'h00000000} /* (7, 19, 29) {real, imag} */,
  {32'hbf353982, 32'h00000000} /* (7, 19, 28) {real, imag} */,
  {32'hbf1a2e40, 32'h00000000} /* (7, 19, 27) {real, imag} */,
  {32'hbf77e41f, 32'h00000000} /* (7, 19, 26) {real, imag} */,
  {32'hbf728db0, 32'h00000000} /* (7, 19, 25) {real, imag} */,
  {32'hbf806971, 32'h00000000} /* (7, 19, 24) {real, imag} */,
  {32'hbfc0788e, 32'h00000000} /* (7, 19, 23) {real, imag} */,
  {32'hbfc665c9, 32'h00000000} /* (7, 19, 22) {real, imag} */,
  {32'hbeeadc86, 32'h00000000} /* (7, 19, 21) {real, imag} */,
  {32'h3f06e303, 32'h00000000} /* (7, 19, 20) {real, imag} */,
  {32'h3f5cfd13, 32'h00000000} /* (7, 19, 19) {real, imag} */,
  {32'h3f96b463, 32'h00000000} /* (7, 19, 18) {real, imag} */,
  {32'h3fdcde78, 32'h00000000} /* (7, 19, 17) {real, imag} */,
  {32'h3fb2c943, 32'h00000000} /* (7, 19, 16) {real, imag} */,
  {32'h3fa10041, 32'h00000000} /* (7, 19, 15) {real, imag} */,
  {32'h3fbed7ba, 32'h00000000} /* (7, 19, 14) {real, imag} */,
  {32'h3fa10bf0, 32'h00000000} /* (7, 19, 13) {real, imag} */,
  {32'h3f4be39c, 32'h00000000} /* (7, 19, 12) {real, imag} */,
  {32'h3ebbc9bb, 32'h00000000} /* (7, 19, 11) {real, imag} */,
  {32'hbf312391, 32'h00000000} /* (7, 19, 10) {real, imag} */,
  {32'hbf75dd63, 32'h00000000} /* (7, 19, 9) {real, imag} */,
  {32'hbfcf9620, 32'h00000000} /* (7, 19, 8) {real, imag} */,
  {32'hbf3d95bd, 32'h00000000} /* (7, 19, 7) {real, imag} */,
  {32'hbec793f4, 32'h00000000} /* (7, 19, 6) {real, imag} */,
  {32'hbf126714, 32'h00000000} /* (7, 19, 5) {real, imag} */,
  {32'hbf827666, 32'h00000000} /* (7, 19, 4) {real, imag} */,
  {32'hbf9e2902, 32'h00000000} /* (7, 19, 3) {real, imag} */,
  {32'hbf937d6d, 32'h00000000} /* (7, 19, 2) {real, imag} */,
  {32'hbf8ed3b4, 32'h00000000} /* (7, 19, 1) {real, imag} */,
  {32'hbefc5c10, 32'h00000000} /* (7, 19, 0) {real, imag} */,
  {32'hbf246312, 32'h00000000} /* (7, 18, 31) {real, imag} */,
  {32'hbfa0d21a, 32'h00000000} /* (7, 18, 30) {real, imag} */,
  {32'hbf373845, 32'h00000000} /* (7, 18, 29) {real, imag} */,
  {32'hbf087a92, 32'h00000000} /* (7, 18, 28) {real, imag} */,
  {32'hbf6b90e4, 32'h00000000} /* (7, 18, 27) {real, imag} */,
  {32'hbf5496d4, 32'h00000000} /* (7, 18, 26) {real, imag} */,
  {32'hbf698e53, 32'h00000000} /* (7, 18, 25) {real, imag} */,
  {32'hbfc87f7e, 32'h00000000} /* (7, 18, 24) {real, imag} */,
  {32'hbfa817e6, 32'h00000000} /* (7, 18, 23) {real, imag} */,
  {32'hbf72d884, 32'h00000000} /* (7, 18, 22) {real, imag} */,
  {32'hbe859aac, 32'h00000000} /* (7, 18, 21) {real, imag} */,
  {32'h3f2628d9, 32'h00000000} /* (7, 18, 20) {real, imag} */,
  {32'h3f1e5380, 32'h00000000} /* (7, 18, 19) {real, imag} */,
  {32'h3f26df00, 32'h00000000} /* (7, 18, 18) {real, imag} */,
  {32'h40007939, 32'h00000000} /* (7, 18, 17) {real, imag} */,
  {32'h3fe5a0be, 32'h00000000} /* (7, 18, 16) {real, imag} */,
  {32'h3fbda73c, 32'h00000000} /* (7, 18, 15) {real, imag} */,
  {32'h3fe8ee8d, 32'h00000000} /* (7, 18, 14) {real, imag} */,
  {32'h3fadc9a4, 32'h00000000} /* (7, 18, 13) {real, imag} */,
  {32'h3f5bc14a, 32'h00000000} /* (7, 18, 12) {real, imag} */,
  {32'h3f3166a7, 32'h00000000} /* (7, 18, 11) {real, imag} */,
  {32'hbe7c46d6, 32'h00000000} /* (7, 18, 10) {real, imag} */,
  {32'hbf4836f9, 32'h00000000} /* (7, 18, 9) {real, imag} */,
  {32'hbf9a07ca, 32'h00000000} /* (7, 18, 8) {real, imag} */,
  {32'hbf26460d, 32'h00000000} /* (7, 18, 7) {real, imag} */,
  {32'hbf367ed5, 32'h00000000} /* (7, 18, 6) {real, imag} */,
  {32'hbf270571, 32'h00000000} /* (7, 18, 5) {real, imag} */,
  {32'hbf813da6, 32'h00000000} /* (7, 18, 4) {real, imag} */,
  {32'hbfad9a60, 32'h00000000} /* (7, 18, 3) {real, imag} */,
  {32'hbf7a4678, 32'h00000000} /* (7, 18, 2) {real, imag} */,
  {32'hbf720641, 32'h00000000} /* (7, 18, 1) {real, imag} */,
  {32'hbf18c08c, 32'h00000000} /* (7, 18, 0) {real, imag} */,
  {32'hbf538d81, 32'h00000000} /* (7, 17, 31) {real, imag} */,
  {32'hbfe68da8, 32'h00000000} /* (7, 17, 30) {real, imag} */,
  {32'hbf79cfe2, 32'h00000000} /* (7, 17, 29) {real, imag} */,
  {32'hbf06862f, 32'h00000000} /* (7, 17, 28) {real, imag} */,
  {32'hbf721d58, 32'h00000000} /* (7, 17, 27) {real, imag} */,
  {32'hbf23a308, 32'h00000000} /* (7, 17, 26) {real, imag} */,
  {32'hbfa0656f, 32'h00000000} /* (7, 17, 25) {real, imag} */,
  {32'hbfe0098c, 32'h00000000} /* (7, 17, 24) {real, imag} */,
  {32'hbf81ed59, 32'h00000000} /* (7, 17, 23) {real, imag} */,
  {32'hbf4ad213, 32'h00000000} /* (7, 17, 22) {real, imag} */,
  {32'hbe9a6abe, 32'h00000000} /* (7, 17, 21) {real, imag} */,
  {32'h3eb08e3e, 32'h00000000} /* (7, 17, 20) {real, imag} */,
  {32'h3f1c3838, 32'h00000000} /* (7, 17, 19) {real, imag} */,
  {32'h3f2dfad4, 32'h00000000} /* (7, 17, 18) {real, imag} */,
  {32'h3f874fab, 32'h00000000} /* (7, 17, 17) {real, imag} */,
  {32'h3f5350c0, 32'h00000000} /* (7, 17, 16) {real, imag} */,
  {32'h3fb455c2, 32'h00000000} /* (7, 17, 15) {real, imag} */,
  {32'h3fbcfaa8, 32'h00000000} /* (7, 17, 14) {real, imag} */,
  {32'h3f769bb6, 32'h00000000} /* (7, 17, 13) {real, imag} */,
  {32'h3f8f6d83, 32'h00000000} /* (7, 17, 12) {real, imag} */,
  {32'h3f1f4fa4, 32'h00000000} /* (7, 17, 11) {real, imag} */,
  {32'hbecace34, 32'h00000000} /* (7, 17, 10) {real, imag} */,
  {32'hbf33fff7, 32'h00000000} /* (7, 17, 9) {real, imag} */,
  {32'hbf2d2912, 32'h00000000} /* (7, 17, 8) {real, imag} */,
  {32'hbf2c4ef5, 32'h00000000} /* (7, 17, 7) {real, imag} */,
  {32'hbf9f6292, 32'h00000000} /* (7, 17, 6) {real, imag} */,
  {32'hbf83a1be, 32'h00000000} /* (7, 17, 5) {real, imag} */,
  {32'hbf98d91e, 32'h00000000} /* (7, 17, 4) {real, imag} */,
  {32'hbfcc6cfd, 32'h00000000} /* (7, 17, 3) {real, imag} */,
  {32'hbf91a98c, 32'h00000000} /* (7, 17, 2) {real, imag} */,
  {32'hbf40b811, 32'h00000000} /* (7, 17, 1) {real, imag} */,
  {32'hbebd09a2, 32'h00000000} /* (7, 17, 0) {real, imag} */,
  {32'hbed8bad0, 32'h00000000} /* (7, 16, 31) {real, imag} */,
  {32'hbfae42cf, 32'h00000000} /* (7, 16, 30) {real, imag} */,
  {32'hbf8357bd, 32'h00000000} /* (7, 16, 29) {real, imag} */,
  {32'hbf773dee, 32'h00000000} /* (7, 16, 28) {real, imag} */,
  {32'hbf86001f, 32'h00000000} /* (7, 16, 27) {real, imag} */,
  {32'hbf3d204d, 32'h00000000} /* (7, 16, 26) {real, imag} */,
  {32'hbfbd3da4, 32'h00000000} /* (7, 16, 25) {real, imag} */,
  {32'hbfb2c8e0, 32'h00000000} /* (7, 16, 24) {real, imag} */,
  {32'hbf6a157f, 32'h00000000} /* (7, 16, 23) {real, imag} */,
  {32'hbfa36041, 32'h00000000} /* (7, 16, 22) {real, imag} */,
  {32'hbe735596, 32'h00000000} /* (7, 16, 21) {real, imag} */,
  {32'h3f04f245, 32'h00000000} /* (7, 16, 20) {real, imag} */,
  {32'h3f72a9d5, 32'h00000000} /* (7, 16, 19) {real, imag} */,
  {32'h3fa3b1c0, 32'h00000000} /* (7, 16, 18) {real, imag} */,
  {32'h3f992b4b, 32'h00000000} /* (7, 16, 17) {real, imag} */,
  {32'h3f6c2b1d, 32'h00000000} /* (7, 16, 16) {real, imag} */,
  {32'h3f9b6fc7, 32'h00000000} /* (7, 16, 15) {real, imag} */,
  {32'h3f847346, 32'h00000000} /* (7, 16, 14) {real, imag} */,
  {32'h3f4278ea, 32'h00000000} /* (7, 16, 13) {real, imag} */,
  {32'h3f21eb0d, 32'h00000000} /* (7, 16, 12) {real, imag} */,
  {32'h3eea9a5d, 32'h00000000} /* (7, 16, 11) {real, imag} */,
  {32'hbe44eb1c, 32'h00000000} /* (7, 16, 10) {real, imag} */,
  {32'hbef6867a, 32'h00000000} /* (7, 16, 9) {real, imag} */,
  {32'hbf064ec5, 32'h00000000} /* (7, 16, 8) {real, imag} */,
  {32'hbf55b645, 32'h00000000} /* (7, 16, 7) {real, imag} */,
  {32'hbf99a974, 32'h00000000} /* (7, 16, 6) {real, imag} */,
  {32'hbf373298, 32'h00000000} /* (7, 16, 5) {real, imag} */,
  {32'hbf274189, 32'h00000000} /* (7, 16, 4) {real, imag} */,
  {32'hbf73d48c, 32'h00000000} /* (7, 16, 3) {real, imag} */,
  {32'hbfbb0e63, 32'h00000000} /* (7, 16, 2) {real, imag} */,
  {32'hbfb9bd24, 32'h00000000} /* (7, 16, 1) {real, imag} */,
  {32'hbeeb43cb, 32'h00000000} /* (7, 16, 0) {real, imag} */,
  {32'hbec98186, 32'h00000000} /* (7, 15, 31) {real, imag} */,
  {32'hbf59446d, 32'h00000000} /* (7, 15, 30) {real, imag} */,
  {32'hbfa33bd2, 32'h00000000} /* (7, 15, 29) {real, imag} */,
  {32'hbfce6076, 32'h00000000} /* (7, 15, 28) {real, imag} */,
  {32'hbfd18a98, 32'h00000000} /* (7, 15, 27) {real, imag} */,
  {32'hbfbd6a68, 32'h00000000} /* (7, 15, 26) {real, imag} */,
  {32'hbfde3f32, 32'h00000000} /* (7, 15, 25) {real, imag} */,
  {32'hbf9be536, 32'h00000000} /* (7, 15, 24) {real, imag} */,
  {32'hbf879077, 32'h00000000} /* (7, 15, 23) {real, imag} */,
  {32'hbfa56578, 32'h00000000} /* (7, 15, 22) {real, imag} */,
  {32'h3cf8726c, 32'h00000000} /* (7, 15, 21) {real, imag} */,
  {32'h3f690253, 32'h00000000} /* (7, 15, 20) {real, imag} */,
  {32'h3f3cc8b6, 32'h00000000} /* (7, 15, 19) {real, imag} */,
  {32'h3f677093, 32'h00000000} /* (7, 15, 18) {real, imag} */,
  {32'h3fa515a1, 32'h00000000} /* (7, 15, 17) {real, imag} */,
  {32'h3fc4f07e, 32'h00000000} /* (7, 15, 16) {real, imag} */,
  {32'h3f94877b, 32'h00000000} /* (7, 15, 15) {real, imag} */,
  {32'h3f64ec48, 32'h00000000} /* (7, 15, 14) {real, imag} */,
  {32'h3f992d06, 32'h00000000} /* (7, 15, 13) {real, imag} */,
  {32'h3f5de3db, 32'h00000000} /* (7, 15, 12) {real, imag} */,
  {32'h3ec732be, 32'h00000000} /* (7, 15, 11) {real, imag} */,
  {32'hbe27d08d, 32'h00000000} /* (7, 15, 10) {real, imag} */,
  {32'hbf597f44, 32'h00000000} /* (7, 15, 9) {real, imag} */,
  {32'hbf4dd409, 32'h00000000} /* (7, 15, 8) {real, imag} */,
  {32'hbf8848bd, 32'h00000000} /* (7, 15, 7) {real, imag} */,
  {32'hbf5023da, 32'h00000000} /* (7, 15, 6) {real, imag} */,
  {32'hbed84113, 32'h00000000} /* (7, 15, 5) {real, imag} */,
  {32'hbf367094, 32'h00000000} /* (7, 15, 4) {real, imag} */,
  {32'hbf814fdb, 32'h00000000} /* (7, 15, 3) {real, imag} */,
  {32'hbfcf04b2, 32'h00000000} /* (7, 15, 2) {real, imag} */,
  {32'hbffc8aa1, 32'h00000000} /* (7, 15, 1) {real, imag} */,
  {32'hbf33f50f, 32'h00000000} /* (7, 15, 0) {real, imag} */,
  {32'hbedb341d, 32'h00000000} /* (7, 14, 31) {real, imag} */,
  {32'hbf2650b0, 32'h00000000} /* (7, 14, 30) {real, imag} */,
  {32'hbf5653a0, 32'h00000000} /* (7, 14, 29) {real, imag} */,
  {32'hbfa62c37, 32'h00000000} /* (7, 14, 28) {real, imag} */,
  {32'hbfaae5a4, 32'h00000000} /* (7, 14, 27) {real, imag} */,
  {32'hbf8d4a74, 32'h00000000} /* (7, 14, 26) {real, imag} */,
  {32'hbfc3281e, 32'h00000000} /* (7, 14, 25) {real, imag} */,
  {32'hbf8430be, 32'h00000000} /* (7, 14, 24) {real, imag} */,
  {32'hbf99fb43, 32'h00000000} /* (7, 14, 23) {real, imag} */,
  {32'hbf8f4d9f, 32'h00000000} /* (7, 14, 22) {real, imag} */,
  {32'hbea41b49, 32'h00000000} /* (7, 14, 21) {real, imag} */,
  {32'h3f31853e, 32'h00000000} /* (7, 14, 20) {real, imag} */,
  {32'h3ef76231, 32'h00000000} /* (7, 14, 19) {real, imag} */,
  {32'h3f0584ff, 32'h00000000} /* (7, 14, 18) {real, imag} */,
  {32'h3f2a2ef6, 32'h00000000} /* (7, 14, 17) {real, imag} */,
  {32'h3f8baca7, 32'h00000000} /* (7, 14, 16) {real, imag} */,
  {32'h3f8e4f0b, 32'h00000000} /* (7, 14, 15) {real, imag} */,
  {32'h3f4b37c1, 32'h00000000} /* (7, 14, 14) {real, imag} */,
  {32'h3f90ca10, 32'h00000000} /* (7, 14, 13) {real, imag} */,
  {32'h3f497def, 32'h00000000} /* (7, 14, 12) {real, imag} */,
  {32'h3ec85fa7, 32'h00000000} /* (7, 14, 11) {real, imag} */,
  {32'hbed688d5, 32'h00000000} /* (7, 14, 10) {real, imag} */,
  {32'hbfb3cb5f, 32'h00000000} /* (7, 14, 9) {real, imag} */,
  {32'hbfa6a423, 32'h00000000} /* (7, 14, 8) {real, imag} */,
  {32'hbfb6ee13, 32'h00000000} /* (7, 14, 7) {real, imag} */,
  {32'hbf56ed7c, 32'h00000000} /* (7, 14, 6) {real, imag} */,
  {32'hbf525eb0, 32'h00000000} /* (7, 14, 5) {real, imag} */,
  {32'hbf8ab470, 32'h00000000} /* (7, 14, 4) {real, imag} */,
  {32'hbf8eb985, 32'h00000000} /* (7, 14, 3) {real, imag} */,
  {32'hbf8da42c, 32'h00000000} /* (7, 14, 2) {real, imag} */,
  {32'hbfb9107c, 32'h00000000} /* (7, 14, 1) {real, imag} */,
  {32'hbf05c3d7, 32'h00000000} /* (7, 14, 0) {real, imag} */,
  {32'hbf093cd0, 32'h00000000} /* (7, 13, 31) {real, imag} */,
  {32'hbf73ec99, 32'h00000000} /* (7, 13, 30) {real, imag} */,
  {32'hbf866d8a, 32'h00000000} /* (7, 13, 29) {real, imag} */,
  {32'hbf98bae4, 32'h00000000} /* (7, 13, 28) {real, imag} */,
  {32'hbf8e32bf, 32'h00000000} /* (7, 13, 27) {real, imag} */,
  {32'hbf5530e2, 32'h00000000} /* (7, 13, 26) {real, imag} */,
  {32'hbf862cf0, 32'h00000000} /* (7, 13, 25) {real, imag} */,
  {32'hbf974656, 32'h00000000} /* (7, 13, 24) {real, imag} */,
  {32'hbf9cb007, 32'h00000000} /* (7, 13, 23) {real, imag} */,
  {32'hbf9c77e0, 32'h00000000} /* (7, 13, 22) {real, imag} */,
  {32'hbebb44e7, 32'h00000000} /* (7, 13, 21) {real, imag} */,
  {32'h3f4a5eee, 32'h00000000} /* (7, 13, 20) {real, imag} */,
  {32'h3f5c8b9b, 32'h00000000} /* (7, 13, 19) {real, imag} */,
  {32'h3f56f106, 32'h00000000} /* (7, 13, 18) {real, imag} */,
  {32'h3f4032e5, 32'h00000000} /* (7, 13, 17) {real, imag} */,
  {32'h3f8656d0, 32'h00000000} /* (7, 13, 16) {real, imag} */,
  {32'h3f9059ef, 32'h00000000} /* (7, 13, 15) {real, imag} */,
  {32'h3f1180fd, 32'h00000000} /* (7, 13, 14) {real, imag} */,
  {32'h3eff5c5c, 32'h00000000} /* (7, 13, 13) {real, imag} */,
  {32'h3f2c64c4, 32'h00000000} /* (7, 13, 12) {real, imag} */,
  {32'h3f2f7811, 32'h00000000} /* (7, 13, 11) {real, imag} */,
  {32'hbef9bdc3, 32'h00000000} /* (7, 13, 10) {real, imag} */,
  {32'hbff9cf11, 32'h00000000} /* (7, 13, 9) {real, imag} */,
  {32'hbf7bac1d, 32'h00000000} /* (7, 13, 8) {real, imag} */,
  {32'hbf1ada59, 32'h00000000} /* (7, 13, 7) {real, imag} */,
  {32'hbf7cb391, 32'h00000000} /* (7, 13, 6) {real, imag} */,
  {32'hbfb08d04, 32'h00000000} /* (7, 13, 5) {real, imag} */,
  {32'hbf94f8ed, 32'h00000000} /* (7, 13, 4) {real, imag} */,
  {32'hbf989bd1, 32'h00000000} /* (7, 13, 3) {real, imag} */,
  {32'hbf6e06a4, 32'h00000000} /* (7, 13, 2) {real, imag} */,
  {32'hbf7ad9a6, 32'h00000000} /* (7, 13, 1) {real, imag} */,
  {32'hbeddb544, 32'h00000000} /* (7, 13, 0) {real, imag} */,
  {32'hbdcf2646, 32'h00000000} /* (7, 12, 31) {real, imag} */,
  {32'hbf1c33be, 32'h00000000} /* (7, 12, 30) {real, imag} */,
  {32'hbf9701d9, 32'h00000000} /* (7, 12, 29) {real, imag} */,
  {32'hbfdd8c17, 32'h00000000} /* (7, 12, 28) {real, imag} */,
  {32'hbfb738a2, 32'h00000000} /* (7, 12, 27) {real, imag} */,
  {32'hbf9447d8, 32'h00000000} /* (7, 12, 26) {real, imag} */,
  {32'hbfde9e31, 32'h00000000} /* (7, 12, 25) {real, imag} */,
  {32'hbfcb7674, 32'h00000000} /* (7, 12, 24) {real, imag} */,
  {32'hbf5d6d38, 32'h00000000} /* (7, 12, 23) {real, imag} */,
  {32'hbedc5cdb, 32'h00000000} /* (7, 12, 22) {real, imag} */,
  {32'hbe28d910, 32'h00000000} /* (7, 12, 21) {real, imag} */,
  {32'h3f2d629f, 32'h00000000} /* (7, 12, 20) {real, imag} */,
  {32'h3ed2ce51, 32'h00000000} /* (7, 12, 19) {real, imag} */,
  {32'h3edc057d, 32'h00000000} /* (7, 12, 18) {real, imag} */,
  {32'h3f2dc3bb, 32'h00000000} /* (7, 12, 17) {real, imag} */,
  {32'h3f3a8216, 32'h00000000} /* (7, 12, 16) {real, imag} */,
  {32'h3f718a68, 32'h00000000} /* (7, 12, 15) {real, imag} */,
  {32'h3f1ee98a, 32'h00000000} /* (7, 12, 14) {real, imag} */,
  {32'h3f32431e, 32'h00000000} /* (7, 12, 13) {real, imag} */,
  {32'h3f8b7bc3, 32'h00000000} /* (7, 12, 12) {real, imag} */,
  {32'h3f4fccc3, 32'h00000000} /* (7, 12, 11) {real, imag} */,
  {32'hbe82e0ef, 32'h00000000} /* (7, 12, 10) {real, imag} */,
  {32'hbf9b4b4d, 32'h00000000} /* (7, 12, 9) {real, imag} */,
  {32'hbf391989, 32'h00000000} /* (7, 12, 8) {real, imag} */,
  {32'hbf36c51e, 32'h00000000} /* (7, 12, 7) {real, imag} */,
  {32'hbfbe8d72, 32'h00000000} /* (7, 12, 6) {real, imag} */,
  {32'hbfa1fd3d, 32'h00000000} /* (7, 12, 5) {real, imag} */,
  {32'hbf2d572b, 32'h00000000} /* (7, 12, 4) {real, imag} */,
  {32'hbec2186a, 32'h00000000} /* (7, 12, 3) {real, imag} */,
  {32'hbef0129e, 32'h00000000} /* (7, 12, 2) {real, imag} */,
  {32'hbf3adc4a, 32'h00000000} /* (7, 12, 1) {real, imag} */,
  {32'hbec341bc, 32'h00000000} /* (7, 12, 0) {real, imag} */,
  {32'hbd2c9e89, 32'h00000000} /* (7, 11, 31) {real, imag} */,
  {32'hbed5d81a, 32'h00000000} /* (7, 11, 30) {real, imag} */,
  {32'hbf346762, 32'h00000000} /* (7, 11, 29) {real, imag} */,
  {32'hbf5115d8, 32'h00000000} /* (7, 11, 28) {real, imag} */,
  {32'hbf7e3789, 32'h00000000} /* (7, 11, 27) {real, imag} */,
  {32'hbf6b7150, 32'h00000000} /* (7, 11, 26) {real, imag} */,
  {32'hbfa40470, 32'h00000000} /* (7, 11, 25) {real, imag} */,
  {32'hbf40cdc8, 32'h00000000} /* (7, 11, 24) {real, imag} */,
  {32'hbea3849b, 32'h00000000} /* (7, 11, 23) {real, imag} */,
  {32'hbf039acd, 32'h00000000} /* (7, 11, 22) {real, imag} */,
  {32'hbe8c0cb7, 32'h00000000} /* (7, 11, 21) {real, imag} */,
  {32'h3edb53ec, 32'h00000000} /* (7, 11, 20) {real, imag} */,
  {32'h3e95dde2, 32'h00000000} /* (7, 11, 19) {real, imag} */,
  {32'h3e9ccf96, 32'h00000000} /* (7, 11, 18) {real, imag} */,
  {32'h3e5f208b, 32'h00000000} /* (7, 11, 17) {real, imag} */,
  {32'h3ec391de, 32'h00000000} /* (7, 11, 16) {real, imag} */,
  {32'h3f0c93b6, 32'h00000000} /* (7, 11, 15) {real, imag} */,
  {32'h3f335dd8, 32'h00000000} /* (7, 11, 14) {real, imag} */,
  {32'h3f5f67ee, 32'h00000000} /* (7, 11, 13) {real, imag} */,
  {32'h3f86106d, 32'h00000000} /* (7, 11, 12) {real, imag} */,
  {32'h3f376a8d, 32'h00000000} /* (7, 11, 11) {real, imag} */,
  {32'hbee96dbb, 32'h00000000} /* (7, 11, 10) {real, imag} */,
  {32'hbf4cda66, 32'h00000000} /* (7, 11, 9) {real, imag} */,
  {32'hbf288e49, 32'h00000000} /* (7, 11, 8) {real, imag} */,
  {32'hbf07505f, 32'h00000000} /* (7, 11, 7) {real, imag} */,
  {32'hbf978661, 32'h00000000} /* (7, 11, 6) {real, imag} */,
  {32'hbf97af89, 32'h00000000} /* (7, 11, 5) {real, imag} */,
  {32'hbeb700fd, 32'h00000000} /* (7, 11, 4) {real, imag} */,
  {32'hbe58dbb4, 32'h00000000} /* (7, 11, 3) {real, imag} */,
  {32'hbf1c9d43, 32'h00000000} /* (7, 11, 2) {real, imag} */,
  {32'hbf87d04a, 32'h00000000} /* (7, 11, 1) {real, imag} */,
  {32'hbf1307f5, 32'h00000000} /* (7, 11, 0) {real, imag} */,
  {32'h3eadf28a, 32'h00000000} /* (7, 10, 31) {real, imag} */,
  {32'h3e4c40be, 32'h00000000} /* (7, 10, 30) {real, imag} */,
  {32'h3d8f7c6b, 32'h00000000} /* (7, 10, 29) {real, imag} */,
  {32'h3f15ea89, 32'h00000000} /* (7, 10, 28) {real, imag} */,
  {32'h3f07926b, 32'h00000000} /* (7, 10, 27) {real, imag} */,
  {32'h3cb8d5ef, 32'h00000000} /* (7, 10, 26) {real, imag} */,
  {32'h3e83d87d, 32'h00000000} /* (7, 10, 25) {real, imag} */,
  {32'h3f171211, 32'h00000000} /* (7, 10, 24) {real, imag} */,
  {32'h3f1a9bcb, 32'h00000000} /* (7, 10, 23) {real, imag} */,
  {32'h3e4b1368, 32'h00000000} /* (7, 10, 22) {real, imag} */,
  {32'h3e954ea1, 32'h00000000} /* (7, 10, 21) {real, imag} */,
  {32'hbcc0819d, 32'h00000000} /* (7, 10, 20) {real, imag} */,
  {32'hbebdf332, 32'h00000000} /* (7, 10, 19) {real, imag} */,
  {32'hbeb56174, 32'h00000000} /* (7, 10, 18) {real, imag} */,
  {32'hbf7f6e7d, 32'h00000000} /* (7, 10, 17) {real, imag} */,
  {32'hbfbbb7b3, 32'h00000000} /* (7, 10, 16) {real, imag} */,
  {32'hbf446c24, 32'h00000000} /* (7, 10, 15) {real, imag} */,
  {32'hbe4284da, 32'h00000000} /* (7, 10, 14) {real, imag} */,
  {32'hbe3d6496, 32'h00000000} /* (7, 10, 13) {real, imag} */,
  {32'hbf056575, 32'h00000000} /* (7, 10, 12) {real, imag} */,
  {32'hbf423cca, 32'h00000000} /* (7, 10, 11) {real, imag} */,
  {32'hbca324c8, 32'h00000000} /* (7, 10, 10) {real, imag} */,
  {32'h3e920361, 32'h00000000} /* (7, 10, 9) {real, imag} */,
  {32'h3ed11b75, 32'h00000000} /* (7, 10, 8) {real, imag} */,
  {32'h3f4b4f87, 32'h00000000} /* (7, 10, 7) {real, imag} */,
  {32'h3ea97124, 32'h00000000} /* (7, 10, 6) {real, imag} */,
  {32'h3e8ab01d, 32'h00000000} /* (7, 10, 5) {real, imag} */,
  {32'h3e8fc597, 32'h00000000} /* (7, 10, 4) {real, imag} */,
  {32'h3e8f99a8, 32'h00000000} /* (7, 10, 3) {real, imag} */,
  {32'h3e866034, 32'h00000000} /* (7, 10, 2) {real, imag} */,
  {32'h3e97996f, 32'h00000000} /* (7, 10, 1) {real, imag} */,
  {32'h3ecfcb15, 32'h00000000} /* (7, 10, 0) {real, imag} */,
  {32'h3f62b110, 32'h00000000} /* (7, 9, 31) {real, imag} */,
  {32'h3f83ee32, 32'h00000000} /* (7, 9, 30) {real, imag} */,
  {32'h3f1eb1fa, 32'h00000000} /* (7, 9, 29) {real, imag} */,
  {32'h3f381402, 32'h00000000} /* (7, 9, 28) {real, imag} */,
  {32'h3f4b7ed5, 32'h00000000} /* (7, 9, 27) {real, imag} */,
  {32'h3f223457, 32'h00000000} /* (7, 9, 26) {real, imag} */,
  {32'h3fb0dd9d, 32'h00000000} /* (7, 9, 25) {real, imag} */,
  {32'h3fae2178, 32'h00000000} /* (7, 9, 24) {real, imag} */,
  {32'h3fa11b2c, 32'h00000000} /* (7, 9, 23) {real, imag} */,
  {32'h3fc174f4, 32'h00000000} /* (7, 9, 22) {real, imag} */,
  {32'h3f891a2e, 32'h00000000} /* (7, 9, 21) {real, imag} */,
  {32'hbe2233d0, 32'h00000000} /* (7, 9, 20) {real, imag} */,
  {32'hbf1976c5, 32'h00000000} /* (7, 9, 19) {real, imag} */,
  {32'hbf892cf6, 32'h00000000} /* (7, 9, 18) {real, imag} */,
  {32'hbfc9c737, 32'h00000000} /* (7, 9, 17) {real, imag} */,
  {32'hbfc5a0ec, 32'h00000000} /* (7, 9, 16) {real, imag} */,
  {32'hbf64b461, 32'h00000000} /* (7, 9, 15) {real, imag} */,
  {32'hbedd0d56, 32'h00000000} /* (7, 9, 14) {real, imag} */,
  {32'hbf81f217, 32'h00000000} /* (7, 9, 13) {real, imag} */,
  {32'hbf47132e, 32'h00000000} /* (7, 9, 12) {real, imag} */,
  {32'hbf2b8ad4, 32'h00000000} /* (7, 9, 11) {real, imag} */,
  {32'hbd4d80b5, 32'h00000000} /* (7, 9, 10) {real, imag} */,
  {32'h3ebdefc8, 32'h00000000} /* (7, 9, 9) {real, imag} */,
  {32'h3f997faf, 32'h00000000} /* (7, 9, 8) {real, imag} */,
  {32'h3fca824e, 32'h00000000} /* (7, 9, 7) {real, imag} */,
  {32'h3f2ef4d5, 32'h00000000} /* (7, 9, 6) {real, imag} */,
  {32'h3f0e7e71, 32'h00000000} /* (7, 9, 5) {real, imag} */,
  {32'h3f13f327, 32'h00000000} /* (7, 9, 4) {real, imag} */,
  {32'h3f664689, 32'h00000000} /* (7, 9, 3) {real, imag} */,
  {32'h3fa26a31, 32'h00000000} /* (7, 9, 2) {real, imag} */,
  {32'h3fbbf564, 32'h00000000} /* (7, 9, 1) {real, imag} */,
  {32'h3f76549f, 32'h00000000} /* (7, 9, 0) {real, imag} */,
  {32'h3f288305, 32'h00000000} /* (7, 8, 31) {real, imag} */,
  {32'h3f85edb6, 32'h00000000} /* (7, 8, 30) {real, imag} */,
  {32'h3f20f088, 32'h00000000} /* (7, 8, 29) {real, imag} */,
  {32'h3f096054, 32'h00000000} /* (7, 8, 28) {real, imag} */,
  {32'h3f02b674, 32'h00000000} /* (7, 8, 27) {real, imag} */,
  {32'h3f3ef65d, 32'h00000000} /* (7, 8, 26) {real, imag} */,
  {32'h3f4385b0, 32'h00000000} /* (7, 8, 25) {real, imag} */,
  {32'h3f7a6f96, 32'h00000000} /* (7, 8, 24) {real, imag} */,
  {32'h3fb685d8, 32'h00000000} /* (7, 8, 23) {real, imag} */,
  {32'h3fdb3ca6, 32'h00000000} /* (7, 8, 22) {real, imag} */,
  {32'h3e209093, 32'h00000000} /* (7, 8, 21) {real, imag} */,
  {32'hbf429d39, 32'h00000000} /* (7, 8, 20) {real, imag} */,
  {32'hbf628d71, 32'h00000000} /* (7, 8, 19) {real, imag} */,
  {32'hbfb561f6, 32'h00000000} /* (7, 8, 18) {real, imag} */,
  {32'hbfaf3b1f, 32'h00000000} /* (7, 8, 17) {real, imag} */,
  {32'hbf71b10d, 32'h00000000} /* (7, 8, 16) {real, imag} */,
  {32'hbf46c75d, 32'h00000000} /* (7, 8, 15) {real, imag} */,
  {32'hbf361f26, 32'h00000000} /* (7, 8, 14) {real, imag} */,
  {32'hbf474162, 32'h00000000} /* (7, 8, 13) {real, imag} */,
  {32'hbeeb8df3, 32'h00000000} /* (7, 8, 12) {real, imag} */,
  {32'hbf00daa4, 32'h00000000} /* (7, 8, 11) {real, imag} */,
  {32'h3e2f6264, 32'h00000000} /* (7, 8, 10) {real, imag} */,
  {32'h3ed0e3f6, 32'h00000000} /* (7, 8, 9) {real, imag} */,
  {32'h3f808acc, 32'h00000000} /* (7, 8, 8) {real, imag} */,
  {32'h3f88f1b4, 32'h00000000} /* (7, 8, 7) {real, imag} */,
  {32'h3edcab34, 32'h00000000} /* (7, 8, 6) {real, imag} */,
  {32'h3ee6a085, 32'h00000000} /* (7, 8, 5) {real, imag} */,
  {32'h3f6b2557, 32'h00000000} /* (7, 8, 4) {real, imag} */,
  {32'h3f86ae5c, 32'h00000000} /* (7, 8, 3) {real, imag} */,
  {32'h3f97bca0, 32'h00000000} /* (7, 8, 2) {real, imag} */,
  {32'h3f98fcdd, 32'h00000000} /* (7, 8, 1) {real, imag} */,
  {32'h3f404464, 32'h00000000} /* (7, 8, 0) {real, imag} */,
  {32'h3f4b6184, 32'h00000000} /* (7, 7, 31) {real, imag} */,
  {32'h3fbca222, 32'h00000000} /* (7, 7, 30) {real, imag} */,
  {32'h3f507eeb, 32'h00000000} /* (7, 7, 29) {real, imag} */,
  {32'h3ed215cb, 32'h00000000} /* (7, 7, 28) {real, imag} */,
  {32'h3f1ab142, 32'h00000000} /* (7, 7, 27) {real, imag} */,
  {32'h3ec7de56, 32'h00000000} /* (7, 7, 26) {real, imag} */,
  {32'h3eb639bd, 32'h00000000} /* (7, 7, 25) {real, imag} */,
  {32'h3f9b2200, 32'h00000000} /* (7, 7, 24) {real, imag} */,
  {32'h3f94133f, 32'h00000000} /* (7, 7, 23) {real, imag} */,
  {32'h3fba4b87, 32'h00000000} /* (7, 7, 22) {real, imag} */,
  {32'h3e990ea4, 32'h00000000} /* (7, 7, 21) {real, imag} */,
  {32'hbf5f21d5, 32'h00000000} /* (7, 7, 20) {real, imag} */,
  {32'hbf9881f6, 32'h00000000} /* (7, 7, 19) {real, imag} */,
  {32'hbfa4ddff, 32'h00000000} /* (7, 7, 18) {real, imag} */,
  {32'hbf937dbe, 32'h00000000} /* (7, 7, 17) {real, imag} */,
  {32'hbfaa79c1, 32'h00000000} /* (7, 7, 16) {real, imag} */,
  {32'hbfa699b0, 32'h00000000} /* (7, 7, 15) {real, imag} */,
  {32'hbf972aa5, 32'h00000000} /* (7, 7, 14) {real, imag} */,
  {32'hbf700b89, 32'h00000000} /* (7, 7, 13) {real, imag} */,
  {32'hbf49db53, 32'h00000000} /* (7, 7, 12) {real, imag} */,
  {32'hbf6c7c67, 32'h00000000} /* (7, 7, 11) {real, imag} */,
  {32'h3eda2312, 32'h00000000} /* (7, 7, 10) {real, imag} */,
  {32'h3f572356, 32'h00000000} /* (7, 7, 9) {real, imag} */,
  {32'h3fcd61c1, 32'h00000000} /* (7, 7, 8) {real, imag} */,
  {32'h3f3f1272, 32'h00000000} /* (7, 7, 7) {real, imag} */,
  {32'h3ebf0983, 32'h00000000} /* (7, 7, 6) {real, imag} */,
  {32'h3f0ca817, 32'h00000000} /* (7, 7, 5) {real, imag} */,
  {32'h3f8847a2, 32'h00000000} /* (7, 7, 4) {real, imag} */,
  {32'h3f9dd897, 32'h00000000} /* (7, 7, 3) {real, imag} */,
  {32'h3f4926b8, 32'h00000000} /* (7, 7, 2) {real, imag} */,
  {32'h3f310789, 32'h00000000} /* (7, 7, 1) {real, imag} */,
  {32'h3ed7b17f, 32'h00000000} /* (7, 7, 0) {real, imag} */,
  {32'h3f24594b, 32'h00000000} /* (7, 6, 31) {real, imag} */,
  {32'h3facca64, 32'h00000000} /* (7, 6, 30) {real, imag} */,
  {32'h3f8b683f, 32'h00000000} /* (7, 6, 29) {real, imag} */,
  {32'h3f5e16af, 32'h00000000} /* (7, 6, 28) {real, imag} */,
  {32'h3fa4c6c4, 32'h00000000} /* (7, 6, 27) {real, imag} */,
  {32'h3f924c37, 32'h00000000} /* (7, 6, 26) {real, imag} */,
  {32'h3f5fe15c, 32'h00000000} /* (7, 6, 25) {real, imag} */,
  {32'h3f842db7, 32'h00000000} /* (7, 6, 24) {real, imag} */,
  {32'h3f3ce6f6, 32'h00000000} /* (7, 6, 23) {real, imag} */,
  {32'h3fa0d942, 32'h00000000} /* (7, 6, 22) {real, imag} */,
  {32'h3ee46466, 32'h00000000} /* (7, 6, 21) {real, imag} */,
  {32'hbf9c9ee8, 32'h00000000} /* (7, 6, 20) {real, imag} */,
  {32'hbf859706, 32'h00000000} /* (7, 6, 19) {real, imag} */,
  {32'hbf314245, 32'h00000000} /* (7, 6, 18) {real, imag} */,
  {32'hbf7bd8fa, 32'h00000000} /* (7, 6, 17) {real, imag} */,
  {32'hbf924972, 32'h00000000} /* (7, 6, 16) {real, imag} */,
  {32'hbf8c0926, 32'h00000000} /* (7, 6, 15) {real, imag} */,
  {32'hbf7b30da, 32'h00000000} /* (7, 6, 14) {real, imag} */,
  {32'hbf57dbde, 32'h00000000} /* (7, 6, 13) {real, imag} */,
  {32'hbf7c0169, 32'h00000000} /* (7, 6, 12) {real, imag} */,
  {32'hbf9aadfb, 32'h00000000} /* (7, 6, 11) {real, imag} */,
  {32'h3ddadb03, 32'h00000000} /* (7, 6, 10) {real, imag} */,
  {32'h3f2eaf8a, 32'h00000000} /* (7, 6, 9) {real, imag} */,
  {32'h3fc68bb9, 32'h00000000} /* (7, 6, 8) {real, imag} */,
  {32'h3eb59c1f, 32'h00000000} /* (7, 6, 7) {real, imag} */,
  {32'h3f0fee20, 32'h00000000} /* (7, 6, 6) {real, imag} */,
  {32'h3fa9f999, 32'h00000000} /* (7, 6, 5) {real, imag} */,
  {32'h3f9942a2, 32'h00000000} /* (7, 6, 4) {real, imag} */,
  {32'h3f6695bd, 32'h00000000} /* (7, 6, 3) {real, imag} */,
  {32'h3fb37634, 32'h00000000} /* (7, 6, 2) {real, imag} */,
  {32'h3fbd0759, 32'h00000000} /* (7, 6, 1) {real, imag} */,
  {32'h3f0c7830, 32'h00000000} /* (7, 6, 0) {real, imag} */,
  {32'h3f235d4c, 32'h00000000} /* (7, 5, 31) {real, imag} */,
  {32'h3f030a11, 32'h00000000} /* (7, 5, 30) {real, imag} */,
  {32'h3f4753cf, 32'h00000000} /* (7, 5, 29) {real, imag} */,
  {32'h3fa2d161, 32'h00000000} /* (7, 5, 28) {real, imag} */,
  {32'h3fbf4f04, 32'h00000000} /* (7, 5, 27) {real, imag} */,
  {32'h3f7583e5, 32'h00000000} /* (7, 5, 26) {real, imag} */,
  {32'h3f8072d5, 32'h00000000} /* (7, 5, 25) {real, imag} */,
  {32'h3f532e90, 32'h00000000} /* (7, 5, 24) {real, imag} */,
  {32'h3f890f03, 32'h00000000} /* (7, 5, 23) {real, imag} */,
  {32'h3fa313f3, 32'h00000000} /* (7, 5, 22) {real, imag} */,
  {32'h3f2290d6, 32'h00000000} /* (7, 5, 21) {real, imag} */,
  {32'hbd81ea83, 32'h00000000} /* (7, 5, 20) {real, imag} */,
  {32'h3e90a80b, 32'h00000000} /* (7, 5, 19) {real, imag} */,
  {32'h3eabf10e, 32'h00000000} /* (7, 5, 18) {real, imag} */,
  {32'h3e75b0c3, 32'h00000000} /* (7, 5, 17) {real, imag} */,
  {32'hbe0c376a, 32'h00000000} /* (7, 5, 16) {real, imag} */,
  {32'hbfa041bb, 32'h00000000} /* (7, 5, 15) {real, imag} */,
  {32'hbfc3c429, 32'h00000000} /* (7, 5, 14) {real, imag} */,
  {32'hbf8276c6, 32'h00000000} /* (7, 5, 13) {real, imag} */,
  {32'hbf9b9c24, 32'h00000000} /* (7, 5, 12) {real, imag} */,
  {32'hbf8a308a, 32'h00000000} /* (7, 5, 11) {real, imag} */,
  {32'hbe86d06d, 32'h00000000} /* (7, 5, 10) {real, imag} */,
  {32'hbdedde0c, 32'h00000000} /* (7, 5, 9) {real, imag} */,
  {32'hbdf7ff23, 32'h00000000} /* (7, 5, 8) {real, imag} */,
  {32'hbed1960a, 32'h00000000} /* (7, 5, 7) {real, imag} */,
  {32'hbe4f2d80, 32'h00000000} /* (7, 5, 6) {real, imag} */,
  {32'h3f56275d, 32'h00000000} /* (7, 5, 5) {real, imag} */,
  {32'h3f8f6509, 32'h00000000} /* (7, 5, 4) {real, imag} */,
  {32'h3f235367, 32'h00000000} /* (7, 5, 3) {real, imag} */,
  {32'h3fa5c036, 32'h00000000} /* (7, 5, 2) {real, imag} */,
  {32'h3fe45e0c, 32'h00000000} /* (7, 5, 1) {real, imag} */,
  {32'h3f1af1b9, 32'h00000000} /* (7, 5, 0) {real, imag} */,
  {32'h3f171ae8, 32'h00000000} /* (7, 4, 31) {real, imag} */,
  {32'h3f5ea34d, 32'h00000000} /* (7, 4, 30) {real, imag} */,
  {32'h3eaa6e40, 32'h00000000} /* (7, 4, 29) {real, imag} */,
  {32'h3f40e25a, 32'h00000000} /* (7, 4, 28) {real, imag} */,
  {32'h3f92bfe7, 32'h00000000} /* (7, 4, 27) {real, imag} */,
  {32'h3f362531, 32'h00000000} /* (7, 4, 26) {real, imag} */,
  {32'h3f0be23d, 32'h00000000} /* (7, 4, 25) {real, imag} */,
  {32'h3f2f44b6, 32'h00000000} /* (7, 4, 24) {real, imag} */,
  {32'h3f9d223d, 32'h00000000} /* (7, 4, 23) {real, imag} */,
  {32'h3f97f481, 32'h00000000} /* (7, 4, 22) {real, imag} */,
  {32'h3f92f2d1, 32'h00000000} /* (7, 4, 21) {real, imag} */,
  {32'h3f4c1e03, 32'h00000000} /* (7, 4, 20) {real, imag} */,
  {32'h3f618362, 32'h00000000} /* (7, 4, 19) {real, imag} */,
  {32'h3fb73354, 32'h00000000} /* (7, 4, 18) {real, imag} */,
  {32'h3f9ff5d0, 32'h00000000} /* (7, 4, 17) {real, imag} */,
  {32'h3ed8c2e2, 32'h00000000} /* (7, 4, 16) {real, imag} */,
  {32'hbf9ff963, 32'h00000000} /* (7, 4, 15) {real, imag} */,
  {32'hbf8833a5, 32'h00000000} /* (7, 4, 14) {real, imag} */,
  {32'hbf222535, 32'h00000000} /* (7, 4, 13) {real, imag} */,
  {32'hbf883e23, 32'h00000000} /* (7, 4, 12) {real, imag} */,
  {32'hbf827f7e, 32'h00000000} /* (7, 4, 11) {real, imag} */,
  {32'hbf0060de, 32'h00000000} /* (7, 4, 10) {real, imag} */,
  {32'hbeeef3ec, 32'h00000000} /* (7, 4, 9) {real, imag} */,
  {32'hbf406472, 32'h00000000} /* (7, 4, 8) {real, imag} */,
  {32'hbf059b9e, 32'h00000000} /* (7, 4, 7) {real, imag} */,
  {32'hbf2f3e0e, 32'h00000000} /* (7, 4, 6) {real, imag} */,
  {32'hbe014799, 32'h00000000} /* (7, 4, 5) {real, imag} */,
  {32'h3efab26e, 32'h00000000} /* (7, 4, 4) {real, imag} */,
  {32'h3f8f0fbd, 32'h00000000} /* (7, 4, 3) {real, imag} */,
  {32'h3f7c477c, 32'h00000000} /* (7, 4, 2) {real, imag} */,
  {32'h3fae5716, 32'h00000000} /* (7, 4, 1) {real, imag} */,
  {32'h3f273966, 32'h00000000} /* (7, 4, 0) {real, imag} */,
  {32'h3ef8fa0f, 32'h00000000} /* (7, 3, 31) {real, imag} */,
  {32'h3f82736f, 32'h00000000} /* (7, 3, 30) {real, imag} */,
  {32'h3f1213a0, 32'h00000000} /* (7, 3, 29) {real, imag} */,
  {32'h3f0a4b1c, 32'h00000000} /* (7, 3, 28) {real, imag} */,
  {32'h3f508c7a, 32'h00000000} /* (7, 3, 27) {real, imag} */,
  {32'h3f6e0374, 32'h00000000} /* (7, 3, 26) {real, imag} */,
  {32'h3f563d84, 32'h00000000} /* (7, 3, 25) {real, imag} */,
  {32'h3fa11591, 32'h00000000} /* (7, 3, 24) {real, imag} */,
  {32'h3f6da0b2, 32'h00000000} /* (7, 3, 23) {real, imag} */,
  {32'h3f4df9f0, 32'h00000000} /* (7, 3, 22) {real, imag} */,
  {32'h3f9a7425, 32'h00000000} /* (7, 3, 21) {real, imag} */,
  {32'h3f29cf71, 32'h00000000} /* (7, 3, 20) {real, imag} */,
  {32'h3f43aaf5, 32'h00000000} /* (7, 3, 19) {real, imag} */,
  {32'h3fabb721, 32'h00000000} /* (7, 3, 18) {real, imag} */,
  {32'h3f6d9a34, 32'h00000000} /* (7, 3, 17) {real, imag} */,
  {32'h3ed99297, 32'h00000000} /* (7, 3, 16) {real, imag} */,
  {32'hbf0e2ff2, 32'h00000000} /* (7, 3, 15) {real, imag} */,
  {32'hbf3d947f, 32'h00000000} /* (7, 3, 14) {real, imag} */,
  {32'hbf492eef, 32'h00000000} /* (7, 3, 13) {real, imag} */,
  {32'hbf4c53d3, 32'h00000000} /* (7, 3, 12) {real, imag} */,
  {32'hbf21f4c6, 32'h00000000} /* (7, 3, 11) {real, imag} */,
  {32'hbedf3f09, 32'h00000000} /* (7, 3, 10) {real, imag} */,
  {32'hbf2c8935, 32'h00000000} /* (7, 3, 9) {real, imag} */,
  {32'hbf791d56, 32'h00000000} /* (7, 3, 8) {real, imag} */,
  {32'hbfcec15b, 32'h00000000} /* (7, 3, 7) {real, imag} */,
  {32'hbfb3bcb6, 32'h00000000} /* (7, 3, 6) {real, imag} */,
  {32'hbdf25990, 32'h00000000} /* (7, 3, 5) {real, imag} */,
  {32'h3f2e0e08, 32'h00000000} /* (7, 3, 4) {real, imag} */,
  {32'h3fcc54de, 32'h00000000} /* (7, 3, 3) {real, imag} */,
  {32'h3fa74ec4, 32'h00000000} /* (7, 3, 2) {real, imag} */,
  {32'h3f77fb6b, 32'h00000000} /* (7, 3, 1) {real, imag} */,
  {32'h3f186b2b, 32'h00000000} /* (7, 3, 0) {real, imag} */,
  {32'h3edab5bf, 32'h00000000} /* (7, 2, 31) {real, imag} */,
  {32'h3f6d2f2f, 32'h00000000} /* (7, 2, 30) {real, imag} */,
  {32'h3f8b9fa6, 32'h00000000} /* (7, 2, 29) {real, imag} */,
  {32'h3f713f7b, 32'h00000000} /* (7, 2, 28) {real, imag} */,
  {32'h3f50501c, 32'h00000000} /* (7, 2, 27) {real, imag} */,
  {32'h3f833d15, 32'h00000000} /* (7, 2, 26) {real, imag} */,
  {32'h3f8a21ab, 32'h00000000} /* (7, 2, 25) {real, imag} */,
  {32'h3f796cd7, 32'h00000000} /* (7, 2, 24) {real, imag} */,
  {32'h3f56a4bf, 32'h00000000} /* (7, 2, 23) {real, imag} */,
  {32'h3f9f3f6c, 32'h00000000} /* (7, 2, 22) {real, imag} */,
  {32'h3fe01039, 32'h00000000} /* (7, 2, 21) {real, imag} */,
  {32'h3fac44ba, 32'h00000000} /* (7, 2, 20) {real, imag} */,
  {32'h3f9ac7f1, 32'h00000000} /* (7, 2, 19) {real, imag} */,
  {32'h3fb4dbec, 32'h00000000} /* (7, 2, 18) {real, imag} */,
  {32'h3f9ca489, 32'h00000000} /* (7, 2, 17) {real, imag} */,
  {32'h3f41debf, 32'h00000000} /* (7, 2, 16) {real, imag} */,
  {32'hbe166ce1, 32'h00000000} /* (7, 2, 15) {real, imag} */,
  {32'hbf0487f6, 32'h00000000} /* (7, 2, 14) {real, imag} */,
  {32'hbf072b12, 32'h00000000} /* (7, 2, 13) {real, imag} */,
  {32'hbf0f282f, 32'h00000000} /* (7, 2, 12) {real, imag} */,
  {32'hbf486f20, 32'h00000000} /* (7, 2, 11) {real, imag} */,
  {32'hbf38e8cf, 32'h00000000} /* (7, 2, 10) {real, imag} */,
  {32'hbf6dfd52, 32'h00000000} /* (7, 2, 9) {real, imag} */,
  {32'hbf94b7f6, 32'h00000000} /* (7, 2, 8) {real, imag} */,
  {32'hbfc04e56, 32'h00000000} /* (7, 2, 7) {real, imag} */,
  {32'hbfa5a8db, 32'h00000000} /* (7, 2, 6) {real, imag} */,
  {32'h3ae31694, 32'h00000000} /* (7, 2, 5) {real, imag} */,
  {32'h3f8754ff, 32'h00000000} /* (7, 2, 4) {real, imag} */,
  {32'h3fa8cb99, 32'h00000000} /* (7, 2, 3) {real, imag} */,
  {32'h3fa49f9f, 32'h00000000} /* (7, 2, 2) {real, imag} */,
  {32'h3f9f605b, 32'h00000000} /* (7, 2, 1) {real, imag} */,
  {32'h3f667d87, 32'h00000000} /* (7, 2, 0) {real, imag} */,
  {32'h3e8fe972, 32'h00000000} /* (7, 1, 31) {real, imag} */,
  {32'h3f21e048, 32'h00000000} /* (7, 1, 30) {real, imag} */,
  {32'h3f68f3e5, 32'h00000000} /* (7, 1, 29) {real, imag} */,
  {32'h3f84b6f6, 32'h00000000} /* (7, 1, 28) {real, imag} */,
  {32'h3f6ac558, 32'h00000000} /* (7, 1, 27) {real, imag} */,
  {32'h3f38f8d3, 32'h00000000} /* (7, 1, 26) {real, imag} */,
  {32'h3f6d6cdb, 32'h00000000} /* (7, 1, 25) {real, imag} */,
  {32'h3f23aff4, 32'h00000000} /* (7, 1, 24) {real, imag} */,
  {32'h3f0eebb3, 32'h00000000} /* (7, 1, 23) {real, imag} */,
  {32'h3eef81c8, 32'h00000000} /* (7, 1, 22) {real, imag} */,
  {32'h3fa372e1, 32'h00000000} /* (7, 1, 21) {real, imag} */,
  {32'h3fa53769, 32'h00000000} /* (7, 1, 20) {real, imag} */,
  {32'h3f812337, 32'h00000000} /* (7, 1, 19) {real, imag} */,
  {32'h3fc84f44, 32'h00000000} /* (7, 1, 18) {real, imag} */,
  {32'h3fa49c19, 32'h00000000} /* (7, 1, 17) {real, imag} */,
  {32'h3f3c1529, 32'h00000000} /* (7, 1, 16) {real, imag} */,
  {32'hbd264155, 32'h00000000} /* (7, 1, 15) {real, imag} */,
  {32'hbe27981f, 32'h00000000} /* (7, 1, 14) {real, imag} */,
  {32'hbe26b547, 32'h00000000} /* (7, 1, 13) {real, imag} */,
  {32'hbf3483cb, 32'h00000000} /* (7, 1, 12) {real, imag} */,
  {32'hbfa927ef, 32'h00000000} /* (7, 1, 11) {real, imag} */,
  {32'hbf957404, 32'h00000000} /* (7, 1, 10) {real, imag} */,
  {32'hbf937dc0, 32'h00000000} /* (7, 1, 9) {real, imag} */,
  {32'hbf94df84, 32'h00000000} /* (7, 1, 8) {real, imag} */,
  {32'hbf4dae59, 32'h00000000} /* (7, 1, 7) {real, imag} */,
  {32'hbf244a86, 32'h00000000} /* (7, 1, 6) {real, imag} */,
  {32'hbede33fa, 32'h00000000} /* (7, 1, 5) {real, imag} */,
  {32'h3f23d2d5, 32'h00000000} /* (7, 1, 4) {real, imag} */,
  {32'h3fa4d0b1, 32'h00000000} /* (7, 1, 3) {real, imag} */,
  {32'h3f336038, 32'h00000000} /* (7, 1, 2) {real, imag} */,
  {32'h3f580678, 32'h00000000} /* (7, 1, 1) {real, imag} */,
  {32'h3f1bfd03, 32'h00000000} /* (7, 1, 0) {real, imag} */,
  {32'h3ed18cb3, 32'h00000000} /* (7, 0, 31) {real, imag} */,
  {32'h3ec92f39, 32'h00000000} /* (7, 0, 30) {real, imag} */,
  {32'h3e7090e6, 32'h00000000} /* (7, 0, 29) {real, imag} */,
  {32'h3e59896c, 32'h00000000} /* (7, 0, 28) {real, imag} */,
  {32'h3f2f2b38, 32'h00000000} /* (7, 0, 27) {real, imag} */,
  {32'h3f1bdd58, 32'h00000000} /* (7, 0, 26) {real, imag} */,
  {32'h3ed9ebed, 32'h00000000} /* (7, 0, 25) {real, imag} */,
  {32'h3cd06334, 32'h00000000} /* (7, 0, 24) {real, imag} */,
  {32'hbcbf6b39, 32'h00000000} /* (7, 0, 23) {real, imag} */,
  {32'h3d6459c9, 32'h00000000} /* (7, 0, 22) {real, imag} */,
  {32'h3ecc2820, 32'h00000000} /* (7, 0, 21) {real, imag} */,
  {32'h3f1e6ce4, 32'h00000000} /* (7, 0, 20) {real, imag} */,
  {32'h3f285a71, 32'h00000000} /* (7, 0, 19) {real, imag} */,
  {32'h3f6347de, 32'h00000000} /* (7, 0, 18) {real, imag} */,
  {32'h3f387634, 32'h00000000} /* (7, 0, 17) {real, imag} */,
  {32'h3e8acc89, 32'h00000000} /* (7, 0, 16) {real, imag} */,
  {32'hbdf22af5, 32'h00000000} /* (7, 0, 15) {real, imag} */,
  {32'hbf04d662, 32'h00000000} /* (7, 0, 14) {real, imag} */,
  {32'hbedcc153, 32'h00000000} /* (7, 0, 13) {real, imag} */,
  {32'hbf7137ff, 32'h00000000} /* (7, 0, 12) {real, imag} */,
  {32'hbf643fec, 32'h00000000} /* (7, 0, 11) {real, imag} */,
  {32'hbee9197b, 32'h00000000} /* (7, 0, 10) {real, imag} */,
  {32'hbf344922, 32'h00000000} /* (7, 0, 9) {real, imag} */,
  {32'hbf034b3a, 32'h00000000} /* (7, 0, 8) {real, imag} */,
  {32'hbe621a24, 32'h00000000} /* (7, 0, 7) {real, imag} */,
  {32'h3db8fcec, 32'h00000000} /* (7, 0, 6) {real, imag} */,
  {32'hbe186a97, 32'h00000000} /* (7, 0, 5) {real, imag} */,
  {32'h3c31f1ab, 32'h00000000} /* (7, 0, 4) {real, imag} */,
  {32'h3f489d3c, 32'h00000000} /* (7, 0, 3) {real, imag} */,
  {32'h3ea369bc, 32'h00000000} /* (7, 0, 2) {real, imag} */,
  {32'h3e8e9cb1, 32'h00000000} /* (7, 0, 1) {real, imag} */,
  {32'h3e8086d6, 32'h00000000} /* (7, 0, 0) {real, imag} */,
  {32'h3ec17d7f, 32'h00000000} /* (6, 31, 31) {real, imag} */,
  {32'h3f314da6, 32'h00000000} /* (6, 31, 30) {real, imag} */,
  {32'h3f0561d3, 32'h00000000} /* (6, 31, 29) {real, imag} */,
  {32'h3f36d242, 32'h00000000} /* (6, 31, 28) {real, imag} */,
  {32'h3f209699, 32'h00000000} /* (6, 31, 27) {real, imag} */,
  {32'h3f2384d4, 32'h00000000} /* (6, 31, 26) {real, imag} */,
  {32'h3f690a85, 32'h00000000} /* (6, 31, 25) {real, imag} */,
  {32'h3f1f4622, 32'h00000000} /* (6, 31, 24) {real, imag} */,
  {32'h3ed2cecf, 32'h00000000} /* (6, 31, 23) {real, imag} */,
  {32'h3e767b2d, 32'h00000000} /* (6, 31, 22) {real, imag} */,
  {32'h3dc5b7ce, 32'h00000000} /* (6, 31, 21) {real, imag} */,
  {32'hbef9f6c4, 32'h00000000} /* (6, 31, 20) {real, imag} */,
  {32'hbeeb94bf, 32'h00000000} /* (6, 31, 19) {real, imag} */,
  {32'hbe92a857, 32'h00000000} /* (6, 31, 18) {real, imag} */,
  {32'hbecb08c1, 32'h00000000} /* (6, 31, 17) {real, imag} */,
  {32'hbef9d3ea, 32'h00000000} /* (6, 31, 16) {real, imag} */,
  {32'hbea5695f, 32'h00000000} /* (6, 31, 15) {real, imag} */,
  {32'hbf2154a4, 32'h00000000} /* (6, 31, 14) {real, imag} */,
  {32'hbea1f9ac, 32'h00000000} /* (6, 31, 13) {real, imag} */,
  {32'hbec39d22, 32'h00000000} /* (6, 31, 12) {real, imag} */,
  {32'hbeb0b666, 32'h00000000} /* (6, 31, 11) {real, imag} */,
  {32'h3efea797, 32'h00000000} /* (6, 31, 10) {real, imag} */,
  {32'h3e55aae3, 32'h00000000} /* (6, 31, 9) {real, imag} */,
  {32'h3e3c8382, 32'h00000000} /* (6, 31, 8) {real, imag} */,
  {32'h3e3650b4, 32'h00000000} /* (6, 31, 7) {real, imag} */,
  {32'h3e1d1380, 32'h00000000} /* (6, 31, 6) {real, imag} */,
  {32'h3e8b165b, 32'h00000000} /* (6, 31, 5) {real, imag} */,
  {32'h3e46e013, 32'h00000000} /* (6, 31, 4) {real, imag} */,
  {32'h3ed07315, 32'h00000000} /* (6, 31, 3) {real, imag} */,
  {32'h3e76ab79, 32'h00000000} /* (6, 31, 2) {real, imag} */,
  {32'h3f281017, 32'h00000000} /* (6, 31, 1) {real, imag} */,
  {32'h3f1948e4, 32'h00000000} /* (6, 31, 0) {real, imag} */,
  {32'h3f49ef71, 32'h00000000} /* (6, 30, 31) {real, imag} */,
  {32'h3fc4ef4b, 32'h00000000} /* (6, 30, 30) {real, imag} */,
  {32'h3fb51f79, 32'h00000000} /* (6, 30, 29) {real, imag} */,
  {32'h3f9cbc7d, 32'h00000000} /* (6, 30, 28) {real, imag} */,
  {32'h3f62089d, 32'h00000000} /* (6, 30, 27) {real, imag} */,
  {32'h3f63c9a3, 32'h00000000} /* (6, 30, 26) {real, imag} */,
  {32'h3f4d9d24, 32'h00000000} /* (6, 30, 25) {real, imag} */,
  {32'h3f6119db, 32'h00000000} /* (6, 30, 24) {real, imag} */,
  {32'h3f627205, 32'h00000000} /* (6, 30, 23) {real, imag} */,
  {32'h3f75dcf5, 32'h00000000} /* (6, 30, 22) {real, imag} */,
  {32'h3dee7552, 32'h00000000} /* (6, 30, 21) {real, imag} */,
  {32'hbfabec4d, 32'h00000000} /* (6, 30, 20) {real, imag} */,
  {32'hbf85591b, 32'h00000000} /* (6, 30, 19) {real, imag} */,
  {32'hbf54bdaf, 32'h00000000} /* (6, 30, 18) {real, imag} */,
  {32'hbf6659b4, 32'h00000000} /* (6, 30, 17) {real, imag} */,
  {32'hbf4bf16e, 32'h00000000} /* (6, 30, 16) {real, imag} */,
  {32'hbf5eeaea, 32'h00000000} /* (6, 30, 15) {real, imag} */,
  {32'hbfe39f6e, 32'h00000000} /* (6, 30, 14) {real, imag} */,
  {32'hbf6f2c25, 32'h00000000} /* (6, 30, 13) {real, imag} */,
  {32'hbef59095, 32'h00000000} /* (6, 30, 12) {real, imag} */,
  {32'hbf13b60f, 32'h00000000} /* (6, 30, 11) {real, imag} */,
  {32'h3ea43fce, 32'h00000000} /* (6, 30, 10) {real, imag} */,
  {32'h3e49c9ff, 32'h00000000} /* (6, 30, 9) {real, imag} */,
  {32'h3ed928fd, 32'h00000000} /* (6, 30, 8) {real, imag} */,
  {32'h3f203049, 32'h00000000} /* (6, 30, 7) {real, imag} */,
  {32'h3eae0801, 32'h00000000} /* (6, 30, 6) {real, imag} */,
  {32'h3ece5f6d, 32'h00000000} /* (6, 30, 5) {real, imag} */,
  {32'h3f13a635, 32'h00000000} /* (6, 30, 4) {real, imag} */,
  {32'h3f554ce4, 32'h00000000} /* (6, 30, 3) {real, imag} */,
  {32'h3f8259f1, 32'h00000000} /* (6, 30, 2) {real, imag} */,
  {32'h3f981fc5, 32'h00000000} /* (6, 30, 1) {real, imag} */,
  {32'h3f30c140, 32'h00000000} /* (6, 30, 0) {real, imag} */,
  {32'h3f4cc81d, 32'h00000000} /* (6, 29, 31) {real, imag} */,
  {32'h3f957143, 32'h00000000} /* (6, 29, 30) {real, imag} */,
  {32'h3f61b22a, 32'h00000000} /* (6, 29, 29) {real, imag} */,
  {32'h3f7314e9, 32'h00000000} /* (6, 29, 28) {real, imag} */,
  {32'h3f34d26f, 32'h00000000} /* (6, 29, 27) {real, imag} */,
  {32'h3f08ba16, 32'h00000000} /* (6, 29, 26) {real, imag} */,
  {32'h3ddbc108, 32'h00000000} /* (6, 29, 25) {real, imag} */,
  {32'h3f3e00ee, 32'h00000000} /* (6, 29, 24) {real, imag} */,
  {32'h3f497fbe, 32'h00000000} /* (6, 29, 23) {real, imag} */,
  {32'h3f650afc, 32'h00000000} /* (6, 29, 22) {real, imag} */,
  {32'h3f1b50bb, 32'h00000000} /* (6, 29, 21) {real, imag} */,
  {32'hbf7715a5, 32'h00000000} /* (6, 29, 20) {real, imag} */,
  {32'hbf3e99dc, 32'h00000000} /* (6, 29, 19) {real, imag} */,
  {32'hbf51365b, 32'h00000000} /* (6, 29, 18) {real, imag} */,
  {32'hbf2c58dc, 32'h00000000} /* (6, 29, 17) {real, imag} */,
  {32'hbecf3393, 32'h00000000} /* (6, 29, 16) {real, imag} */,
  {32'hbef9c511, 32'h00000000} /* (6, 29, 15) {real, imag} */,
  {32'hbf85b616, 32'h00000000} /* (6, 29, 14) {real, imag} */,
  {32'hbf60c766, 32'h00000000} /* (6, 29, 13) {real, imag} */,
  {32'hbeedeee2, 32'h00000000} /* (6, 29, 12) {real, imag} */,
  {32'hbf16faa3, 32'h00000000} /* (6, 29, 11) {real, imag} */,
  {32'h3eea5703, 32'h00000000} /* (6, 29, 10) {real, imag} */,
  {32'h3f8a30cc, 32'h00000000} /* (6, 29, 9) {real, imag} */,
  {32'h3fba2e99, 32'h00000000} /* (6, 29, 8) {real, imag} */,
  {32'h3f93baf5, 32'h00000000} /* (6, 29, 7) {real, imag} */,
  {32'h3f525e10, 32'h00000000} /* (6, 29, 6) {real, imag} */,
  {32'h3f6639c3, 32'h00000000} /* (6, 29, 5) {real, imag} */,
  {32'h3f535ba6, 32'h00000000} /* (6, 29, 4) {real, imag} */,
  {32'h3f03dc66, 32'h00000000} /* (6, 29, 3) {real, imag} */,
  {32'h3ef06f1f, 32'h00000000} /* (6, 29, 2) {real, imag} */,
  {32'h3f490bee, 32'h00000000} /* (6, 29, 1) {real, imag} */,
  {32'h3f0c23f4, 32'h00000000} /* (6, 29, 0) {real, imag} */,
  {32'h3ef192cd, 32'h00000000} /* (6, 28, 31) {real, imag} */,
  {32'h3f2743a1, 32'h00000000} /* (6, 28, 30) {real, imag} */,
  {32'h3f2a73a1, 32'h00000000} /* (6, 28, 29) {real, imag} */,
  {32'h3f59351c, 32'h00000000} /* (6, 28, 28) {real, imag} */,
  {32'h3f118742, 32'h00000000} /* (6, 28, 27) {real, imag} */,
  {32'h3e6df54c, 32'h00000000} /* (6, 28, 26) {real, imag} */,
  {32'h3e24230a, 32'h00000000} /* (6, 28, 25) {real, imag} */,
  {32'h3f82058a, 32'h00000000} /* (6, 28, 24) {real, imag} */,
  {32'h3f81229c, 32'h00000000} /* (6, 28, 23) {real, imag} */,
  {32'h3f7e109b, 32'h00000000} /* (6, 28, 22) {real, imag} */,
  {32'h3f4a7bb6, 32'h00000000} /* (6, 28, 21) {real, imag} */,
  {32'hbf4d0410, 32'h00000000} /* (6, 28, 20) {real, imag} */,
  {32'hbf3b1c9d, 32'h00000000} /* (6, 28, 19) {real, imag} */,
  {32'hbf6901c3, 32'h00000000} /* (6, 28, 18) {real, imag} */,
  {32'hbf3ed0e3, 32'h00000000} /* (6, 28, 17) {real, imag} */,
  {32'hbeab5e88, 32'h00000000} /* (6, 28, 16) {real, imag} */,
  {32'hbf025fbe, 32'h00000000} /* (6, 28, 15) {real, imag} */,
  {32'hbf61705e, 32'h00000000} /* (6, 28, 14) {real, imag} */,
  {32'hbf3d5a03, 32'h00000000} /* (6, 28, 13) {real, imag} */,
  {32'hbedc1b87, 32'h00000000} /* (6, 28, 12) {real, imag} */,
  {32'hbecb9fc1, 32'h00000000} /* (6, 28, 11) {real, imag} */,
  {32'h3f89e1a4, 32'h00000000} /* (6, 28, 10) {real, imag} */,
  {32'h3fae9b0a, 32'h00000000} /* (6, 28, 9) {real, imag} */,
  {32'h3f98e8b5, 32'h00000000} /* (6, 28, 8) {real, imag} */,
  {32'h3f82f109, 32'h00000000} /* (6, 28, 7) {real, imag} */,
  {32'h3f54d5b8, 32'h00000000} /* (6, 28, 6) {real, imag} */,
  {32'h3f900e8c, 32'h00000000} /* (6, 28, 5) {real, imag} */,
  {32'h3f901353, 32'h00000000} /* (6, 28, 4) {real, imag} */,
  {32'h3f9c1938, 32'h00000000} /* (6, 28, 3) {real, imag} */,
  {32'h3f3d6e9a, 32'h00000000} /* (6, 28, 2) {real, imag} */,
  {32'h3e9cc3cb, 32'h00000000} /* (6, 28, 1) {real, imag} */,
  {32'h3e3fd2ae, 32'h00000000} /* (6, 28, 0) {real, imag} */,
  {32'h3f09c9f0, 32'h00000000} /* (6, 27, 31) {real, imag} */,
  {32'h3efde1f3, 32'h00000000} /* (6, 27, 30) {real, imag} */,
  {32'h3f2368ed, 32'h00000000} /* (6, 27, 29) {real, imag} */,
  {32'h3f29e8cd, 32'h00000000} /* (6, 27, 28) {real, imag} */,
  {32'h3f0206b0, 32'h00000000} /* (6, 27, 27) {real, imag} */,
  {32'h3f18c164, 32'h00000000} /* (6, 27, 26) {real, imag} */,
  {32'h3ec18f61, 32'h00000000} /* (6, 27, 25) {real, imag} */,
  {32'h3f918abe, 32'h00000000} /* (6, 27, 24) {real, imag} */,
  {32'h3fa8585e, 32'h00000000} /* (6, 27, 23) {real, imag} */,
  {32'h3fb3a41d, 32'h00000000} /* (6, 27, 22) {real, imag} */,
  {32'h3f53e23c, 32'h00000000} /* (6, 27, 21) {real, imag} */,
  {32'hbf4fff21, 32'h00000000} /* (6, 27, 20) {real, imag} */,
  {32'hbf7c909b, 32'h00000000} /* (6, 27, 19) {real, imag} */,
  {32'hbf9d482f, 32'h00000000} /* (6, 27, 18) {real, imag} */,
  {32'hbf550cee, 32'h00000000} /* (6, 27, 17) {real, imag} */,
  {32'hbf1da845, 32'h00000000} /* (6, 27, 16) {real, imag} */,
  {32'hbee6fa9e, 32'h00000000} /* (6, 27, 15) {real, imag} */,
  {32'hbf3717d2, 32'h00000000} /* (6, 27, 14) {real, imag} */,
  {32'hbf8e55b0, 32'h00000000} /* (6, 27, 13) {real, imag} */,
  {32'hbf4c737b, 32'h00000000} /* (6, 27, 12) {real, imag} */,
  {32'hbef890cc, 32'h00000000} /* (6, 27, 11) {real, imag} */,
  {32'h3f140657, 32'h00000000} /* (6, 27, 10) {real, imag} */,
  {32'h3f00cfdf, 32'h00000000} /* (6, 27, 9) {real, imag} */,
  {32'h3f5026d3, 32'h00000000} /* (6, 27, 8) {real, imag} */,
  {32'h3f7ae5de, 32'h00000000} /* (6, 27, 7) {real, imag} */,
  {32'h3f63ce4a, 32'h00000000} /* (6, 27, 6) {real, imag} */,
  {32'h3f82fe36, 32'h00000000} /* (6, 27, 5) {real, imag} */,
  {32'h3f3e4e79, 32'h00000000} /* (6, 27, 4) {real, imag} */,
  {32'h3f41da25, 32'h00000000} /* (6, 27, 3) {real, imag} */,
  {32'h3f0d65b4, 32'h00000000} /* (6, 27, 2) {real, imag} */,
  {32'h3f183679, 32'h00000000} /* (6, 27, 1) {real, imag} */,
  {32'h3eb84daa, 32'h00000000} /* (6, 27, 0) {real, imag} */,
  {32'h3ecb8a14, 32'h00000000} /* (6, 26, 31) {real, imag} */,
  {32'h3f03398f, 32'h00000000} /* (6, 26, 30) {real, imag} */,
  {32'h3f75578a, 32'h00000000} /* (6, 26, 29) {real, imag} */,
  {32'h3f55f6f6, 32'h00000000} /* (6, 26, 28) {real, imag} */,
  {32'h3f512f78, 32'h00000000} /* (6, 26, 27) {real, imag} */,
  {32'h3f84fed8, 32'h00000000} /* (6, 26, 26) {real, imag} */,
  {32'h3f07723b, 32'h00000000} /* (6, 26, 25) {real, imag} */,
  {32'h3f0c2ce6, 32'h00000000} /* (6, 26, 24) {real, imag} */,
  {32'h3f1e5301, 32'h00000000} /* (6, 26, 23) {real, imag} */,
  {32'h3f67f786, 32'h00000000} /* (6, 26, 22) {real, imag} */,
  {32'h3ef8b310, 32'h00000000} /* (6, 26, 21) {real, imag} */,
  {32'hbf2f46be, 32'h00000000} /* (6, 26, 20) {real, imag} */,
  {32'hbf7a8669, 32'h00000000} /* (6, 26, 19) {real, imag} */,
  {32'hbf91eaef, 32'h00000000} /* (6, 26, 18) {real, imag} */,
  {32'hbf8221d4, 32'h00000000} /* (6, 26, 17) {real, imag} */,
  {32'hbf205b04, 32'h00000000} /* (6, 26, 16) {real, imag} */,
  {32'hbeb5aeb6, 32'h00000000} /* (6, 26, 15) {real, imag} */,
  {32'hbf4898ea, 32'h00000000} /* (6, 26, 14) {real, imag} */,
  {32'hbfa66df7, 32'h00000000} /* (6, 26, 13) {real, imag} */,
  {32'hbf3ddf8a, 32'h00000000} /* (6, 26, 12) {real, imag} */,
  {32'hbf0d4091, 32'h00000000} /* (6, 26, 11) {real, imag} */,
  {32'h3f0a551f, 32'h00000000} /* (6, 26, 10) {real, imag} */,
  {32'h3f90d3a5, 32'h00000000} /* (6, 26, 9) {real, imag} */,
  {32'h3f6b3a70, 32'h00000000} /* (6, 26, 8) {real, imag} */,
  {32'h3f560a94, 32'h00000000} /* (6, 26, 7) {real, imag} */,
  {32'h3f47b7c0, 32'h00000000} /* (6, 26, 6) {real, imag} */,
  {32'h3f76e008, 32'h00000000} /* (6, 26, 5) {real, imag} */,
  {32'h3f139bdb, 32'h00000000} /* (6, 26, 4) {real, imag} */,
  {32'h3e5653b4, 32'h00000000} /* (6, 26, 3) {real, imag} */,
  {32'h3e91d018, 32'h00000000} /* (6, 26, 2) {real, imag} */,
  {32'h3f3cf673, 32'h00000000} /* (6, 26, 1) {real, imag} */,
  {32'h3e8709f7, 32'h00000000} /* (6, 26, 0) {real, imag} */,
  {32'h3f14c70d, 32'h00000000} /* (6, 25, 31) {real, imag} */,
  {32'h3f624fd6, 32'h00000000} /* (6, 25, 30) {real, imag} */,
  {32'h3f1e1279, 32'h00000000} /* (6, 25, 29) {real, imag} */,
  {32'h3f0bab28, 32'h00000000} /* (6, 25, 28) {real, imag} */,
  {32'h3f49b12e, 32'h00000000} /* (6, 25, 27) {real, imag} */,
  {32'h3f9ce84d, 32'h00000000} /* (6, 25, 26) {real, imag} */,
  {32'h3f2f24b3, 32'h00000000} /* (6, 25, 25) {real, imag} */,
  {32'h3ef1f52c, 32'h00000000} /* (6, 25, 24) {real, imag} */,
  {32'h3ef2b806, 32'h00000000} /* (6, 25, 23) {real, imag} */,
  {32'h3f0dca86, 32'h00000000} /* (6, 25, 22) {real, imag} */,
  {32'h3ec0b73a, 32'h00000000} /* (6, 25, 21) {real, imag} */,
  {32'hbeaf00ff, 32'h00000000} /* (6, 25, 20) {real, imag} */,
  {32'hbf3abb0b, 32'h00000000} /* (6, 25, 19) {real, imag} */,
  {32'hbf747652, 32'h00000000} /* (6, 25, 18) {real, imag} */,
  {32'hbfa16c8f, 32'h00000000} /* (6, 25, 17) {real, imag} */,
  {32'hbf4f962b, 32'h00000000} /* (6, 25, 16) {real, imag} */,
  {32'hbf187e1c, 32'h00000000} /* (6, 25, 15) {real, imag} */,
  {32'hbf2b01f2, 32'h00000000} /* (6, 25, 14) {real, imag} */,
  {32'hbf373157, 32'h00000000} /* (6, 25, 13) {real, imag} */,
  {32'hbf6782ed, 32'h00000000} /* (6, 25, 12) {real, imag} */,
  {32'hbeca5858, 32'h00000000} /* (6, 25, 11) {real, imag} */,
  {32'h3f499451, 32'h00000000} /* (6, 25, 10) {real, imag} */,
  {32'h3f8d5fa0, 32'h00000000} /* (6, 25, 9) {real, imag} */,
  {32'h3f0ff28e, 32'h00000000} /* (6, 25, 8) {real, imag} */,
  {32'h3f12bb30, 32'h00000000} /* (6, 25, 7) {real, imag} */,
  {32'h3f296f8b, 32'h00000000} /* (6, 25, 6) {real, imag} */,
  {32'h3f844d01, 32'h00000000} /* (6, 25, 5) {real, imag} */,
  {32'h3eeee53b, 32'h00000000} /* (6, 25, 4) {real, imag} */,
  {32'h3eaf8c18, 32'h00000000} /* (6, 25, 3) {real, imag} */,
  {32'h3f1e7a29, 32'h00000000} /* (6, 25, 2) {real, imag} */,
  {32'h3f4fdf2a, 32'h00000000} /* (6, 25, 1) {real, imag} */,
  {32'h3e36278a, 32'h00000000} /* (6, 25, 0) {real, imag} */,
  {32'h3f0eafe5, 32'h00000000} /* (6, 24, 31) {real, imag} */,
  {32'h3f8cee55, 32'h00000000} /* (6, 24, 30) {real, imag} */,
  {32'h3f1ee92c, 32'h00000000} /* (6, 24, 29) {real, imag} */,
  {32'h3f449b98, 32'h00000000} /* (6, 24, 28) {real, imag} */,
  {32'h3f631e77, 32'h00000000} /* (6, 24, 27) {real, imag} */,
  {32'h3f518320, 32'h00000000} /* (6, 24, 26) {real, imag} */,
  {32'h3f47fe7b, 32'h00000000} /* (6, 24, 25) {real, imag} */,
  {32'h3f6207f7, 32'h00000000} /* (6, 24, 24) {real, imag} */,
  {32'h3f610a28, 32'h00000000} /* (6, 24, 23) {real, imag} */,
  {32'h3f2ffafb, 32'h00000000} /* (6, 24, 22) {real, imag} */,
  {32'h3f1b3cae, 32'h00000000} /* (6, 24, 21) {real, imag} */,
  {32'hbebdf142, 32'h00000000} /* (6, 24, 20) {real, imag} */,
  {32'hbf30eb50, 32'h00000000} /* (6, 24, 19) {real, imag} */,
  {32'hbf07dd48, 32'h00000000} /* (6, 24, 18) {real, imag} */,
  {32'hbf9d9890, 32'h00000000} /* (6, 24, 17) {real, imag} */,
  {32'hbf98ec89, 32'h00000000} /* (6, 24, 16) {real, imag} */,
  {32'hbf297172, 32'h00000000} /* (6, 24, 15) {real, imag} */,
  {32'hbf2686f0, 32'h00000000} /* (6, 24, 14) {real, imag} */,
  {32'hbee62d16, 32'h00000000} /* (6, 24, 13) {real, imag} */,
  {32'hbf2481ce, 32'h00000000} /* (6, 24, 12) {real, imag} */,
  {32'hbe6075a0, 32'h00000000} /* (6, 24, 11) {real, imag} */,
  {32'h3f44675b, 32'h00000000} /* (6, 24, 10) {real, imag} */,
  {32'h3f32e09c, 32'h00000000} /* (6, 24, 9) {real, imag} */,
  {32'h3f1cb2f7, 32'h00000000} /* (6, 24, 8) {real, imag} */,
  {32'h3ecb6487, 32'h00000000} /* (6, 24, 7) {real, imag} */,
  {32'h3eeeb5af, 32'h00000000} /* (6, 24, 6) {real, imag} */,
  {32'h3f86f4f4, 32'h00000000} /* (6, 24, 5) {real, imag} */,
  {32'h3f31c6fc, 32'h00000000} /* (6, 24, 4) {real, imag} */,
  {32'h3f3eab65, 32'h00000000} /* (6, 24, 3) {real, imag} */,
  {32'h3f6a09ee, 32'h00000000} /* (6, 24, 2) {real, imag} */,
  {32'h3f35b706, 32'h00000000} /* (6, 24, 1) {real, imag} */,
  {32'h3ec735f1, 32'h00000000} /* (6, 24, 0) {real, imag} */,
  {32'h3f48b498, 32'h00000000} /* (6, 23, 31) {real, imag} */,
  {32'h3fa2a133, 32'h00000000} /* (6, 23, 30) {real, imag} */,
  {32'h3f36dd78, 32'h00000000} /* (6, 23, 29) {real, imag} */,
  {32'h3f092ec4, 32'h00000000} /* (6, 23, 28) {real, imag} */,
  {32'h3f80be4c, 32'h00000000} /* (6, 23, 27) {real, imag} */,
  {32'h3f894cac, 32'h00000000} /* (6, 23, 26) {real, imag} */,
  {32'h3f76b0ce, 32'h00000000} /* (6, 23, 25) {real, imag} */,
  {32'h3f594408, 32'h00000000} /* (6, 23, 24) {real, imag} */,
  {32'h3f780d07, 32'h00000000} /* (6, 23, 23) {real, imag} */,
  {32'h3f58c88f, 32'h00000000} /* (6, 23, 22) {real, imag} */,
  {32'h3f1bf421, 32'h00000000} /* (6, 23, 21) {real, imag} */,
  {32'hbe602f56, 32'h00000000} /* (6, 23, 20) {real, imag} */,
  {32'hbecf9b86, 32'h00000000} /* (6, 23, 19) {real, imag} */,
  {32'hbe960bda, 32'h00000000} /* (6, 23, 18) {real, imag} */,
  {32'hbf5bc9cd, 32'h00000000} /* (6, 23, 17) {real, imag} */,
  {32'hbf600db6, 32'h00000000} /* (6, 23, 16) {real, imag} */,
  {32'hbe948be2, 32'h00000000} /* (6, 23, 15) {real, imag} */,
  {32'hbf2a07df, 32'h00000000} /* (6, 23, 14) {real, imag} */,
  {32'hbf1721c5, 32'h00000000} /* (6, 23, 13) {real, imag} */,
  {32'hbef1026a, 32'h00000000} /* (6, 23, 12) {real, imag} */,
  {32'hbe182a14, 32'h00000000} /* (6, 23, 11) {real, imag} */,
  {32'h3ebf9787, 32'h00000000} /* (6, 23, 10) {real, imag} */,
  {32'h3edb9226, 32'h00000000} /* (6, 23, 9) {real, imag} */,
  {32'h3f53969b, 32'h00000000} /* (6, 23, 8) {real, imag} */,
  {32'h3ee0fa3a, 32'h00000000} /* (6, 23, 7) {real, imag} */,
  {32'h3ec75c8b, 32'h00000000} /* (6, 23, 6) {real, imag} */,
  {32'h3ee79973, 32'h00000000} /* (6, 23, 5) {real, imag} */,
  {32'h3ef1a1e1, 32'h00000000} /* (6, 23, 4) {real, imag} */,
  {32'h3ebdc849, 32'h00000000} /* (6, 23, 3) {real, imag} */,
  {32'h3ec89507, 32'h00000000} /* (6, 23, 2) {real, imag} */,
  {32'h3ebec3c7, 32'h00000000} /* (6, 23, 1) {real, imag} */,
  {32'h3ec33f68, 32'h00000000} /* (6, 23, 0) {real, imag} */,
  {32'h3eb21ccc, 32'h00000000} /* (6, 22, 31) {real, imag} */,
  {32'h3edd1264, 32'h00000000} /* (6, 22, 30) {real, imag} */,
  {32'h3eded580, 32'h00000000} /* (6, 22, 29) {real, imag} */,
  {32'h3f6d6622, 32'h00000000} /* (6, 22, 28) {real, imag} */,
  {32'h3fc4069d, 32'h00000000} /* (6, 22, 27) {real, imag} */,
  {32'h3fae73fc, 32'h00000000} /* (6, 22, 26) {real, imag} */,
  {32'h3f864f9f, 32'h00000000} /* (6, 22, 25) {real, imag} */,
  {32'h3f3b9de4, 32'h00000000} /* (6, 22, 24) {real, imag} */,
  {32'h3fb1d612, 32'h00000000} /* (6, 22, 23) {real, imag} */,
  {32'h3f93b6dc, 32'h00000000} /* (6, 22, 22) {real, imag} */,
  {32'h3ecb8f80, 32'h00000000} /* (6, 22, 21) {real, imag} */,
  {32'hbeb151b3, 32'h00000000} /* (6, 22, 20) {real, imag} */,
  {32'hbe8fbf6a, 32'h00000000} /* (6, 22, 19) {real, imag} */,
  {32'hbea396b4, 32'h00000000} /* (6, 22, 18) {real, imag} */,
  {32'hbf53fcc0, 32'h00000000} /* (6, 22, 17) {real, imag} */,
  {32'hbf2f5af4, 32'h00000000} /* (6, 22, 16) {real, imag} */,
  {32'hbf31cf10, 32'h00000000} /* (6, 22, 15) {real, imag} */,
  {32'hbf565a0b, 32'h00000000} /* (6, 22, 14) {real, imag} */,
  {32'hbf264955, 32'h00000000} /* (6, 22, 13) {real, imag} */,
  {32'hbf7114ef, 32'h00000000} /* (6, 22, 12) {real, imag} */,
  {32'hbf220779, 32'h00000000} /* (6, 22, 11) {real, imag} */,
  {32'h3f001995, 32'h00000000} /* (6, 22, 10) {real, imag} */,
  {32'h3f8d67a2, 32'h00000000} /* (6, 22, 9) {real, imag} */,
  {32'h3fab6663, 32'h00000000} /* (6, 22, 8) {real, imag} */,
  {32'h3f7bc2a6, 32'h00000000} /* (6, 22, 7) {real, imag} */,
  {32'h3f8779d8, 32'h00000000} /* (6, 22, 6) {real, imag} */,
  {32'h3f377a21, 32'h00000000} /* (6, 22, 5) {real, imag} */,
  {32'h3e105984, 32'h00000000} /* (6, 22, 4) {real, imag} */,
  {32'h3e4ba79e, 32'h00000000} /* (6, 22, 3) {real, imag} */,
  {32'h3e90d799, 32'h00000000} /* (6, 22, 2) {real, imag} */,
  {32'h3eca2724, 32'h00000000} /* (6, 22, 1) {real, imag} */,
  {32'h3e8c7bbd, 32'h00000000} /* (6, 22, 0) {real, imag} */,
  {32'hbe21b448, 32'h00000000} /* (6, 21, 31) {real, imag} */,
  {32'h3e9e1d28, 32'h00000000} /* (6, 21, 30) {real, imag} */,
  {32'h3f1593b2, 32'h00000000} /* (6, 21, 29) {real, imag} */,
  {32'h3fa8de6e, 32'h00000000} /* (6, 21, 28) {real, imag} */,
  {32'h3fc01473, 32'h00000000} /* (6, 21, 27) {real, imag} */,
  {32'h3f528ea0, 32'h00000000} /* (6, 21, 26) {real, imag} */,
  {32'h3f59806a, 32'h00000000} /* (6, 21, 25) {real, imag} */,
  {32'h3f0bd700, 32'h00000000} /* (6, 21, 24) {real, imag} */,
  {32'h3efb6b36, 32'h00000000} /* (6, 21, 23) {real, imag} */,
  {32'h3e825b60, 32'h00000000} /* (6, 21, 22) {real, imag} */,
  {32'hbe201a78, 32'h00000000} /* (6, 21, 21) {real, imag} */,
  {32'hbebeb5e6, 32'h00000000} /* (6, 21, 20) {real, imag} */,
  {32'h3e407e51, 32'h00000000} /* (6, 21, 19) {real, imag} */,
  {32'h3e0fd0ed, 32'h00000000} /* (6, 21, 18) {real, imag} */,
  {32'hbeec95e0, 32'h00000000} /* (6, 21, 17) {real, imag} */,
  {32'hbef16bb5, 32'h00000000} /* (6, 21, 16) {real, imag} */,
  {32'hbeb424e7, 32'h00000000} /* (6, 21, 15) {real, imag} */,
  {32'hbd272d15, 32'h00000000} /* (6, 21, 14) {real, imag} */,
  {32'hbe248a5c, 32'h00000000} /* (6, 21, 13) {real, imag} */,
  {32'hbe55fe88, 32'h00000000} /* (6, 21, 12) {real, imag} */,
  {32'hbd7670ce, 32'h00000000} /* (6, 21, 11) {real, imag} */,
  {32'h3ef7ed94, 32'h00000000} /* (6, 21, 10) {real, imag} */,
  {32'h3f122701, 32'h00000000} /* (6, 21, 9) {real, imag} */,
  {32'h3f8519f5, 32'h00000000} /* (6, 21, 8) {real, imag} */,
  {32'h3f39676c, 32'h00000000} /* (6, 21, 7) {real, imag} */,
  {32'h3f5bbbe9, 32'h00000000} /* (6, 21, 6) {real, imag} */,
  {32'h3ecfd9b8, 32'h00000000} /* (6, 21, 5) {real, imag} */,
  {32'hbdaad28e, 32'h00000000} /* (6, 21, 4) {real, imag} */,
  {32'hbc9c30ac, 32'h00000000} /* (6, 21, 3) {real, imag} */,
  {32'h3e9efb8d, 32'h00000000} /* (6, 21, 2) {real, imag} */,
  {32'h3eb73d80, 32'h00000000} /* (6, 21, 1) {real, imag} */,
  {32'h3db6606a, 32'h00000000} /* (6, 21, 0) {real, imag} */,
  {32'hbea05c5f, 32'h00000000} /* (6, 20, 31) {real, imag} */,
  {32'h3d4283db, 32'h00000000} /* (6, 20, 30) {real, imag} */,
  {32'hbe3c6e82, 32'h00000000} /* (6, 20, 29) {real, imag} */,
  {32'h3e8187e0, 32'h00000000} /* (6, 20, 28) {real, imag} */,
  {32'h3e3fdb66, 32'h00000000} /* (6, 20, 27) {real, imag} */,
  {32'hbe9a5f65, 32'h00000000} /* (6, 20, 26) {real, imag} */,
  {32'hbf258483, 32'h00000000} /* (6, 20, 25) {real, imag} */,
  {32'hbeef5712, 32'h00000000} /* (6, 20, 24) {real, imag} */,
  {32'hbf47b6bf, 32'h00000000} /* (6, 20, 23) {real, imag} */,
  {32'hbf313f65, 32'h00000000} /* (6, 20, 22) {real, imag} */,
  {32'hbe217cce, 32'h00000000} /* (6, 20, 21) {real, imag} */,
  {32'h3eade125, 32'h00000000} /* (6, 20, 20) {real, imag} */,
  {32'h3f377795, 32'h00000000} /* (6, 20, 19) {real, imag} */,
  {32'h3f749f21, 32'h00000000} /* (6, 20, 18) {real, imag} */,
  {32'h3f34a2b6, 32'h00000000} /* (6, 20, 17) {real, imag} */,
  {32'h3ef76244, 32'h00000000} /* (6, 20, 16) {real, imag} */,
  {32'h3f2a482c, 32'h00000000} /* (6, 20, 15) {real, imag} */,
  {32'h3f5e96f6, 32'h00000000} /* (6, 20, 14) {real, imag} */,
  {32'h3f0a92e2, 32'h00000000} /* (6, 20, 13) {real, imag} */,
  {32'h3f159f8e, 32'h00000000} /* (6, 20, 12) {real, imag} */,
  {32'h3d5a6022, 32'h00000000} /* (6, 20, 11) {real, imag} */,
  {32'hbf258933, 32'h00000000} /* (6, 20, 10) {real, imag} */,
  {32'hbf004fe5, 32'h00000000} /* (6, 20, 9) {real, imag} */,
  {32'hbedaf08d, 32'h00000000} /* (6, 20, 8) {real, imag} */,
  {32'hbf10cd6b, 32'h00000000} /* (6, 20, 7) {real, imag} */,
  {32'hbe91242d, 32'h00000000} /* (6, 20, 6) {real, imag} */,
  {32'hbe38a940, 32'h00000000} /* (6, 20, 5) {real, imag} */,
  {32'hbf2fac5c, 32'h00000000} /* (6, 20, 4) {real, imag} */,
  {32'hbf652d99, 32'h00000000} /* (6, 20, 3) {real, imag} */,
  {32'hbec81a78, 32'h00000000} /* (6, 20, 2) {real, imag} */,
  {32'hbf164256, 32'h00000000} /* (6, 20, 1) {real, imag} */,
  {32'hbec2b437, 32'h00000000} /* (6, 20, 0) {real, imag} */,
  {32'hbe7bdb44, 32'h00000000} /* (6, 19, 31) {real, imag} */,
  {32'hbe432610, 32'h00000000} /* (6, 19, 30) {real, imag} */,
  {32'hbf10d0a4, 32'h00000000} /* (6, 19, 29) {real, imag} */,
  {32'hbeba10ce, 32'h00000000} /* (6, 19, 28) {real, imag} */,
  {32'hbf0a3c59, 32'h00000000} /* (6, 19, 27) {real, imag} */,
  {32'hbf603986, 32'h00000000} /* (6, 19, 26) {real, imag} */,
  {32'hbfb3c2f3, 32'h00000000} /* (6, 19, 25) {real, imag} */,
  {32'hbfc2f2cd, 32'h00000000} /* (6, 19, 24) {real, imag} */,
  {32'hbfad0204, 32'h00000000} /* (6, 19, 23) {real, imag} */,
  {32'hbf8691f4, 32'h00000000} /* (6, 19, 22) {real, imag} */,
  {32'hbe94a807, 32'h00000000} /* (6, 19, 21) {real, imag} */,
  {32'h3f189ebc, 32'h00000000} /* (6, 19, 20) {real, imag} */,
  {32'h3f7cb503, 32'h00000000} /* (6, 19, 19) {real, imag} */,
  {32'h3fa73ea8, 32'h00000000} /* (6, 19, 18) {real, imag} */,
  {32'h3fc0ab01, 32'h00000000} /* (6, 19, 17) {real, imag} */,
  {32'h3f7a080c, 32'h00000000} /* (6, 19, 16) {real, imag} */,
  {32'h3f5a3a42, 32'h00000000} /* (6, 19, 15) {real, imag} */,
  {32'h3f630ca5, 32'h00000000} /* (6, 19, 14) {real, imag} */,
  {32'h3f5282c5, 32'h00000000} /* (6, 19, 13) {real, imag} */,
  {32'h3f4d4291, 32'h00000000} /* (6, 19, 12) {real, imag} */,
  {32'hbe1afc60, 32'h00000000} /* (6, 19, 11) {real, imag} */,
  {32'hbf2e5a38, 32'h00000000} /* (6, 19, 10) {real, imag} */,
  {32'h390a8c08, 32'h00000000} /* (6, 19, 9) {real, imag} */,
  {32'hbed868f8, 32'h00000000} /* (6, 19, 8) {real, imag} */,
  {32'hbde4f5fc, 32'h00000000} /* (6, 19, 7) {real, imag} */,
  {32'h3dd84a85, 32'h00000000} /* (6, 19, 6) {real, imag} */,
  {32'hbec1fb4b, 32'h00000000} /* (6, 19, 5) {real, imag} */,
  {32'hbf356267, 32'h00000000} /* (6, 19, 4) {real, imag} */,
  {32'hbf33700e, 32'h00000000} /* (6, 19, 3) {real, imag} */,
  {32'hbf358960, 32'h00000000} /* (6, 19, 2) {real, imag} */,
  {32'hbf785264, 32'h00000000} /* (6, 19, 1) {real, imag} */,
  {32'hbf2f9bfe, 32'h00000000} /* (6, 19, 0) {real, imag} */,
  {32'hbec37a21, 32'h00000000} /* (6, 18, 31) {real, imag} */,
  {32'hbf1b6c3b, 32'h00000000} /* (6, 18, 30) {real, imag} */,
  {32'hbf01190c, 32'h00000000} /* (6, 18, 29) {real, imag} */,
  {32'hbeda6f97, 32'h00000000} /* (6, 18, 28) {real, imag} */,
  {32'hbf49bfe9, 32'h00000000} /* (6, 18, 27) {real, imag} */,
  {32'hbf2cc587, 32'h00000000} /* (6, 18, 26) {real, imag} */,
  {32'hbf81c1c7, 32'h00000000} /* (6, 18, 25) {real, imag} */,
  {32'hbfe8e406, 32'h00000000} /* (6, 18, 24) {real, imag} */,
  {32'hbf718d73, 32'h00000000} /* (6, 18, 23) {real, imag} */,
  {32'hbec5d469, 32'h00000000} /* (6, 18, 22) {real, imag} */,
  {32'hbd800452, 32'h00000000} /* (6, 18, 21) {real, imag} */,
  {32'h3f78d8f3, 32'h00000000} /* (6, 18, 20) {real, imag} */,
  {32'h3f952411, 32'h00000000} /* (6, 18, 19) {real, imag} */,
  {32'h3f924149, 32'h00000000} /* (6, 18, 18) {real, imag} */,
  {32'h3fd32e20, 32'h00000000} /* (6, 18, 17) {real, imag} */,
  {32'h3f9137f1, 32'h00000000} /* (6, 18, 16) {real, imag} */,
  {32'h3f844373, 32'h00000000} /* (6, 18, 15) {real, imag} */,
  {32'h3f8dbc73, 32'h00000000} /* (6, 18, 14) {real, imag} */,
  {32'h3f8e01cf, 32'h00000000} /* (6, 18, 13) {real, imag} */,
  {32'h3f2b2c02, 32'h00000000} /* (6, 18, 12) {real, imag} */,
  {32'h3da1981c, 32'h00000000} /* (6, 18, 11) {real, imag} */,
  {32'hbeb18d88, 32'h00000000} /* (6, 18, 10) {real, imag} */,
  {32'hbf037695, 32'h00000000} /* (6, 18, 9) {real, imag} */,
  {32'hbf3d0423, 32'h00000000} /* (6, 18, 8) {real, imag} */,
  {32'hbe607cd9, 32'h00000000} /* (6, 18, 7) {real, imag} */,
  {32'hbd159b8c, 32'h00000000} /* (6, 18, 6) {real, imag} */,
  {32'hbdc1800a, 32'h00000000} /* (6, 18, 5) {real, imag} */,
  {32'hbf18d8f3, 32'h00000000} /* (6, 18, 4) {real, imag} */,
  {32'hbf31824d, 32'h00000000} /* (6, 18, 3) {real, imag} */,
  {32'hbeff164a, 32'h00000000} /* (6, 18, 2) {real, imag} */,
  {32'hbeb0fc3d, 32'h00000000} /* (6, 18, 1) {real, imag} */,
  {32'hbee1a4b2, 32'h00000000} /* (6, 18, 0) {real, imag} */,
  {32'hbeb355d7, 32'h00000000} /* (6, 17, 31) {real, imag} */,
  {32'hbf4c02e5, 32'h00000000} /* (6, 17, 30) {real, imag} */,
  {32'hbf3c4de7, 32'h00000000} /* (6, 17, 29) {real, imag} */,
  {32'hbef1646f, 32'h00000000} /* (6, 17, 28) {real, imag} */,
  {32'hbf20b4c2, 32'h00000000} /* (6, 17, 27) {real, imag} */,
  {32'hbf2c2dff, 32'h00000000} /* (6, 17, 26) {real, imag} */,
  {32'hbf902806, 32'h00000000} /* (6, 17, 25) {real, imag} */,
  {32'hbfa3edeb, 32'h00000000} /* (6, 17, 24) {real, imag} */,
  {32'hbec8a68a, 32'h00000000} /* (6, 17, 23) {real, imag} */,
  {32'hbedb48ba, 32'h00000000} /* (6, 17, 22) {real, imag} */,
  {32'hbe29ebc0, 32'h00000000} /* (6, 17, 21) {real, imag} */,
  {32'h3f3c2e98, 32'h00000000} /* (6, 17, 20) {real, imag} */,
  {32'h3f512648, 32'h00000000} /* (6, 17, 19) {real, imag} */,
  {32'h3f4f9e32, 32'h00000000} /* (6, 17, 18) {real, imag} */,
  {32'h3fa3851b, 32'h00000000} /* (6, 17, 17) {real, imag} */,
  {32'h3f952002, 32'h00000000} /* (6, 17, 16) {real, imag} */,
  {32'h3fb4fa07, 32'h00000000} /* (6, 17, 15) {real, imag} */,
  {32'h3fa353b6, 32'h00000000} /* (6, 17, 14) {real, imag} */,
  {32'h3f936add, 32'h00000000} /* (6, 17, 13) {real, imag} */,
  {32'h3f91d990, 32'h00000000} /* (6, 17, 12) {real, imag} */,
  {32'h3e2a4050, 32'h00000000} /* (6, 17, 11) {real, imag} */,
  {32'hbf2085a8, 32'h00000000} /* (6, 17, 10) {real, imag} */,
  {32'hbf711514, 32'h00000000} /* (6, 17, 9) {real, imag} */,
  {32'hbe94c705, 32'h00000000} /* (6, 17, 8) {real, imag} */,
  {32'hbf3579df, 32'h00000000} /* (6, 17, 7) {real, imag} */,
  {32'hbf77f8a9, 32'h00000000} /* (6, 17, 6) {real, imag} */,
  {32'hbf2a59e7, 32'h00000000} /* (6, 17, 5) {real, imag} */,
  {32'hbf3b2cf4, 32'h00000000} /* (6, 17, 4) {real, imag} */,
  {32'hbf211bb8, 32'h00000000} /* (6, 17, 3) {real, imag} */,
  {32'hbea58a50, 32'h00000000} /* (6, 17, 2) {real, imag} */,
  {32'hbe96a60d, 32'h00000000} /* (6, 17, 1) {real, imag} */,
  {32'hbe5e5193, 32'h00000000} /* (6, 17, 0) {real, imag} */,
  {32'hbe0a55de, 32'h00000000} /* (6, 16, 31) {real, imag} */,
  {32'hbf4b1176, 32'h00000000} /* (6, 16, 30) {real, imag} */,
  {32'hbf757be4, 32'h00000000} /* (6, 16, 29) {real, imag} */,
  {32'hbf05a441, 32'h00000000} /* (6, 16, 28) {real, imag} */,
  {32'hbf474ffc, 32'h00000000} /* (6, 16, 27) {real, imag} */,
  {32'hbf2be15c, 32'h00000000} /* (6, 16, 26) {real, imag} */,
  {32'hbf5986a0, 32'h00000000} /* (6, 16, 25) {real, imag} */,
  {32'hbf394853, 32'h00000000} /* (6, 16, 24) {real, imag} */,
  {32'hbe8a6954, 32'h00000000} /* (6, 16, 23) {real, imag} */,
  {32'hbf5f2326, 32'h00000000} /* (6, 16, 22) {real, imag} */,
  {32'hbeaeea81, 32'h00000000} /* (6, 16, 21) {real, imag} */,
  {32'h3f24235d, 32'h00000000} /* (6, 16, 20) {real, imag} */,
  {32'h3f500f8e, 32'h00000000} /* (6, 16, 19) {real, imag} */,
  {32'h3f3d7a13, 32'h00000000} /* (6, 16, 18) {real, imag} */,
  {32'h3f3ec8d0, 32'h00000000} /* (6, 16, 17) {real, imag} */,
  {32'h3f816eed, 32'h00000000} /* (6, 16, 16) {real, imag} */,
  {32'h3fc64787, 32'h00000000} /* (6, 16, 15) {real, imag} */,
  {32'h3fa5aa0b, 32'h00000000} /* (6, 16, 14) {real, imag} */,
  {32'h3f7d487a, 32'h00000000} /* (6, 16, 13) {real, imag} */,
  {32'h3f1b98d9, 32'h00000000} /* (6, 16, 12) {real, imag} */,
  {32'h3d9f9e8f, 32'h00000000} /* (6, 16, 11) {real, imag} */,
  {32'hbe8df286, 32'h00000000} /* (6, 16, 10) {real, imag} */,
  {32'hbf2d8bad, 32'h00000000} /* (6, 16, 9) {real, imag} */,
  {32'hbf494671, 32'h00000000} /* (6, 16, 8) {real, imag} */,
  {32'hbfa41632, 32'h00000000} /* (6, 16, 7) {real, imag} */,
  {32'hbf592924, 32'h00000000} /* (6, 16, 6) {real, imag} */,
  {32'hbf19a2c4, 32'h00000000} /* (6, 16, 5) {real, imag} */,
  {32'hbf63ee80, 32'h00000000} /* (6, 16, 4) {real, imag} */,
  {32'hbf8f4d00, 32'h00000000} /* (6, 16, 3) {real, imag} */,
  {32'hbfb9497d, 32'h00000000} /* (6, 16, 2) {real, imag} */,
  {32'hbfd8efde, 32'h00000000} /* (6, 16, 1) {real, imag} */,
  {32'hbf1f177d, 32'h00000000} /* (6, 16, 0) {real, imag} */,
  {32'hbd300461, 32'h00000000} /* (6, 15, 31) {real, imag} */,
  {32'hbf01eb1d, 32'h00000000} /* (6, 15, 30) {real, imag} */,
  {32'hbf3034bf, 32'h00000000} /* (6, 15, 29) {real, imag} */,
  {32'hbf7106df, 32'h00000000} /* (6, 15, 28) {real, imag} */,
  {32'hbf93d74b, 32'h00000000} /* (6, 15, 27) {real, imag} */,
  {32'hbf4dbccf, 32'h00000000} /* (6, 15, 26) {real, imag} */,
  {32'hbfaa40e8, 32'h00000000} /* (6, 15, 25) {real, imag} */,
  {32'hbf54902e, 32'h00000000} /* (6, 15, 24) {real, imag} */,
  {32'hbf2fc1e5, 32'h00000000} /* (6, 15, 23) {real, imag} */,
  {32'hbf4051cc, 32'h00000000} /* (6, 15, 22) {real, imag} */,
  {32'hbc73048f, 32'h00000000} /* (6, 15, 21) {real, imag} */,
  {32'h3f9011da, 32'h00000000} /* (6, 15, 20) {real, imag} */,
  {32'h3f7b63c4, 32'h00000000} /* (6, 15, 19) {real, imag} */,
  {32'h3f00f8d6, 32'h00000000} /* (6, 15, 18) {real, imag} */,
  {32'h3f06e589, 32'h00000000} /* (6, 15, 17) {real, imag} */,
  {32'h3fb14510, 32'h00000000} /* (6, 15, 16) {real, imag} */,
  {32'h3f8cc689, 32'h00000000} /* (6, 15, 15) {real, imag} */,
  {32'h3f6d1a46, 32'h00000000} /* (6, 15, 14) {real, imag} */,
  {32'h3f2342a3, 32'h00000000} /* (6, 15, 13) {real, imag} */,
  {32'h3e2fbb6e, 32'h00000000} /* (6, 15, 12) {real, imag} */,
  {32'h3db817e8, 32'h00000000} /* (6, 15, 11) {real, imag} */,
  {32'hbe9f0fa6, 32'h00000000} /* (6, 15, 10) {real, imag} */,
  {32'hbf335e0c, 32'h00000000} /* (6, 15, 9) {real, imag} */,
  {32'hbf78a23f, 32'h00000000} /* (6, 15, 8) {real, imag} */,
  {32'hbfa4e220, 32'h00000000} /* (6, 15, 7) {real, imag} */,
  {32'hbf3825c0, 32'h00000000} /* (6, 15, 6) {real, imag} */,
  {32'hbe877921, 32'h00000000} /* (6, 15, 5) {real, imag} */,
  {32'hbf2f85c4, 32'h00000000} /* (6, 15, 4) {real, imag} */,
  {32'hbfbec1af, 32'h00000000} /* (6, 15, 3) {real, imag} */,
  {32'hc006adea, 32'h00000000} /* (6, 15, 2) {real, imag} */,
  {32'hbfecb1a6, 32'h00000000} /* (6, 15, 1) {real, imag} */,
  {32'hbf2a81eb, 32'h00000000} /* (6, 15, 0) {real, imag} */,
  {32'hbe898673, 32'h00000000} /* (6, 14, 31) {real, imag} */,
  {32'hbf1a5a31, 32'h00000000} /* (6, 14, 30) {real, imag} */,
  {32'hbf3c84e2, 32'h00000000} /* (6, 14, 29) {real, imag} */,
  {32'hbf88fa69, 32'h00000000} /* (6, 14, 28) {real, imag} */,
  {32'hbf6fba6a, 32'h00000000} /* (6, 14, 27) {real, imag} */,
  {32'hbf831d3b, 32'h00000000} /* (6, 14, 26) {real, imag} */,
  {32'hbfcaf7c5, 32'h00000000} /* (6, 14, 25) {real, imag} */,
  {32'hbfacc21e, 32'h00000000} /* (6, 14, 24) {real, imag} */,
  {32'hbfbb10ba, 32'h00000000} /* (6, 14, 23) {real, imag} */,
  {32'hbf6bb391, 32'h00000000} /* (6, 14, 22) {real, imag} */,
  {32'hbdb80c62, 32'h00000000} /* (6, 14, 21) {real, imag} */,
  {32'h3f65af77, 32'h00000000} /* (6, 14, 20) {real, imag} */,
  {32'h3ec491c7, 32'h00000000} /* (6, 14, 19) {real, imag} */,
  {32'h3e9b7780, 32'h00000000} /* (6, 14, 18) {real, imag} */,
  {32'h3ea90dbd, 32'h00000000} /* (6, 14, 17) {real, imag} */,
  {32'h3f80e0bb, 32'h00000000} /* (6, 14, 16) {real, imag} */,
  {32'h3f693528, 32'h00000000} /* (6, 14, 15) {real, imag} */,
  {32'h3f7efc8d, 32'h00000000} /* (6, 14, 14) {real, imag} */,
  {32'h3f710244, 32'h00000000} /* (6, 14, 13) {real, imag} */,
  {32'h3ee8c3d2, 32'h00000000} /* (6, 14, 12) {real, imag} */,
  {32'h3e2a01f8, 32'h00000000} /* (6, 14, 11) {real, imag} */,
  {32'hbfa784a0, 32'h00000000} /* (6, 14, 10) {real, imag} */,
  {32'hbfa4cbe2, 32'h00000000} /* (6, 14, 9) {real, imag} */,
  {32'hbf06c935, 32'h00000000} /* (6, 14, 8) {real, imag} */,
  {32'hbf981323, 32'h00000000} /* (6, 14, 7) {real, imag} */,
  {32'hbf8771cf, 32'h00000000} /* (6, 14, 6) {real, imag} */,
  {32'hbf1a03f7, 32'h00000000} /* (6, 14, 5) {real, imag} */,
  {32'hbf2317cf, 32'h00000000} /* (6, 14, 4) {real, imag} */,
  {32'hbf8a710e, 32'h00000000} /* (6, 14, 3) {real, imag} */,
  {32'hbfb3a362, 32'h00000000} /* (6, 14, 2) {real, imag} */,
  {32'hbf5806ca, 32'h00000000} /* (6, 14, 1) {real, imag} */,
  {32'hbe1a00bd, 32'h00000000} /* (6, 14, 0) {real, imag} */,
  {32'hbee4af02, 32'h00000000} /* (6, 13, 31) {real, imag} */,
  {32'hbf7c7186, 32'h00000000} /* (6, 13, 30) {real, imag} */,
  {32'hbf696fbd, 32'h00000000} /* (6, 13, 29) {real, imag} */,
  {32'hbf637443, 32'h00000000} /* (6, 13, 28) {real, imag} */,
  {32'hbf5b0837, 32'h00000000} /* (6, 13, 27) {real, imag} */,
  {32'hbf31067e, 32'h00000000} /* (6, 13, 26) {real, imag} */,
  {32'hbfa34547, 32'h00000000} /* (6, 13, 25) {real, imag} */,
  {32'hbfe98cca, 32'h00000000} /* (6, 13, 24) {real, imag} */,
  {32'hbfa9dc62, 32'h00000000} /* (6, 13, 23) {real, imag} */,
  {32'hbf57cc28, 32'h00000000} /* (6, 13, 22) {real, imag} */,
  {32'hbed2926e, 32'h00000000} /* (6, 13, 21) {real, imag} */,
  {32'h3f0f8512, 32'h00000000} /* (6, 13, 20) {real, imag} */,
  {32'h3eb47f0f, 32'h00000000} /* (6, 13, 19) {real, imag} */,
  {32'h3ee353fe, 32'h00000000} /* (6, 13, 18) {real, imag} */,
  {32'h3f2f39a2, 32'h00000000} /* (6, 13, 17) {real, imag} */,
  {32'h3f51d308, 32'h00000000} /* (6, 13, 16) {real, imag} */,
  {32'h3f5cc69e, 32'h00000000} /* (6, 13, 15) {real, imag} */,
  {32'h3f08ac07, 32'h00000000} /* (6, 13, 14) {real, imag} */,
  {32'h3f7eb0cc, 32'h00000000} /* (6, 13, 13) {real, imag} */,
  {32'h3f564fa2, 32'h00000000} /* (6, 13, 12) {real, imag} */,
  {32'h3e9f2975, 32'h00000000} /* (6, 13, 11) {real, imag} */,
  {32'hbfbc5b31, 32'h00000000} /* (6, 13, 10) {real, imag} */,
  {32'hc0031ca6, 32'h00000000} /* (6, 13, 9) {real, imag} */,
  {32'hbf2412c9, 32'h00000000} /* (6, 13, 8) {real, imag} */,
  {32'hbf9993cf, 32'h00000000} /* (6, 13, 7) {real, imag} */,
  {32'hbf9ad8dc, 32'h00000000} /* (6, 13, 6) {real, imag} */,
  {32'hbf249905, 32'h00000000} /* (6, 13, 5) {real, imag} */,
  {32'hbf60b999, 32'h00000000} /* (6, 13, 4) {real, imag} */,
  {32'hbfb62b5f, 32'h00000000} /* (6, 13, 3) {real, imag} */,
  {32'hbf5bc02c, 32'h00000000} /* (6, 13, 2) {real, imag} */,
  {32'hbe9e9feb, 32'h00000000} /* (6, 13, 1) {real, imag} */,
  {32'h3c2cc74c, 32'h00000000} /* (6, 13, 0) {real, imag} */,
  {32'hbed32c83, 32'h00000000} /* (6, 12, 31) {real, imag} */,
  {32'hbf5ea0e2, 32'h00000000} /* (6, 12, 30) {real, imag} */,
  {32'hbf4dea4b, 32'h00000000} /* (6, 12, 29) {real, imag} */,
  {32'hbf367c47, 32'h00000000} /* (6, 12, 28) {real, imag} */,
  {32'hbf67882b, 32'h00000000} /* (6, 12, 27) {real, imag} */,
  {32'hbf8fe2cd, 32'h00000000} /* (6, 12, 26) {real, imag} */,
  {32'hbfa6f81b, 32'h00000000} /* (6, 12, 25) {real, imag} */,
  {32'hbfce3b98, 32'h00000000} /* (6, 12, 24) {real, imag} */,
  {32'hbf94ecb4, 32'h00000000} /* (6, 12, 23) {real, imag} */,
  {32'hbf0cd2bf, 32'h00000000} /* (6, 12, 22) {real, imag} */,
  {32'hbf1d8adb, 32'h00000000} /* (6, 12, 21) {real, imag} */,
  {32'h3e8586da, 32'h00000000} /* (6, 12, 20) {real, imag} */,
  {32'h3e43adf6, 32'h00000000} /* (6, 12, 19) {real, imag} */,
  {32'h3ec5740e, 32'h00000000} /* (6, 12, 18) {real, imag} */,
  {32'h3f8257b8, 32'h00000000} /* (6, 12, 17) {real, imag} */,
  {32'h3f578e83, 32'h00000000} /* (6, 12, 16) {real, imag} */,
  {32'h3f15ed5e, 32'h00000000} /* (6, 12, 15) {real, imag} */,
  {32'h3f126763, 32'h00000000} /* (6, 12, 14) {real, imag} */,
  {32'h3fa534de, 32'h00000000} /* (6, 12, 13) {real, imag} */,
  {32'h3fe30283, 32'h00000000} /* (6, 12, 12) {real, imag} */,
  {32'h3eee16d5, 32'h00000000} /* (6, 12, 11) {real, imag} */,
  {32'hbf03c5ed, 32'h00000000} /* (6, 12, 10) {real, imag} */,
  {32'hbf84bba2, 32'h00000000} /* (6, 12, 9) {real, imag} */,
  {32'hbf7f0a2c, 32'h00000000} /* (6, 12, 8) {real, imag} */,
  {32'hbf4e55e4, 32'h00000000} /* (6, 12, 7) {real, imag} */,
  {32'hbf8deebf, 32'h00000000} /* (6, 12, 6) {real, imag} */,
  {32'hbf58aeb0, 32'h00000000} /* (6, 12, 5) {real, imag} */,
  {32'hbf2fb4be, 32'h00000000} /* (6, 12, 4) {real, imag} */,
  {32'hbf135db7, 32'h00000000} /* (6, 12, 3) {real, imag} */,
  {32'hbf1dc9f5, 32'h00000000} /* (6, 12, 2) {real, imag} */,
  {32'hbef24a04, 32'h00000000} /* (6, 12, 1) {real, imag} */,
  {32'hbe5b764b, 32'h00000000} /* (6, 12, 0) {real, imag} */,
  {32'hbd450767, 32'h00000000} /* (6, 11, 31) {real, imag} */,
  {32'hbe850029, 32'h00000000} /* (6, 11, 30) {real, imag} */,
  {32'hbf615b2a, 32'h00000000} /* (6, 11, 29) {real, imag} */,
  {32'hbf2abbdf, 32'h00000000} /* (6, 11, 28) {real, imag} */,
  {32'hbf5a8ebb, 32'h00000000} /* (6, 11, 27) {real, imag} */,
  {32'hbf818f76, 32'h00000000} /* (6, 11, 26) {real, imag} */,
  {32'hbf550ebc, 32'h00000000} /* (6, 11, 25) {real, imag} */,
  {32'hbf1ed6e9, 32'h00000000} /* (6, 11, 24) {real, imag} */,
  {32'hbf02eeeb, 32'h00000000} /* (6, 11, 23) {real, imag} */,
  {32'hbeadf771, 32'h00000000} /* (6, 11, 22) {real, imag} */,
  {32'hbeeb52f5, 32'h00000000} /* (6, 11, 21) {real, imag} */,
  {32'h3dd6a18f, 32'h00000000} /* (6, 11, 20) {real, imag} */,
  {32'hbd4f47a5, 32'h00000000} /* (6, 11, 19) {real, imag} */,
  {32'h3ec90f57, 32'h00000000} /* (6, 11, 18) {real, imag} */,
  {32'h3f2ae717, 32'h00000000} /* (6, 11, 17) {real, imag} */,
  {32'h3f1829c3, 32'h00000000} /* (6, 11, 16) {real, imag} */,
  {32'h3ebb6607, 32'h00000000} /* (6, 11, 15) {real, imag} */,
  {32'h3f47da7d, 32'h00000000} /* (6, 11, 14) {real, imag} */,
  {32'h3f52ee1c, 32'h00000000} /* (6, 11, 13) {real, imag} */,
  {32'h3f4df6de, 32'h00000000} /* (6, 11, 12) {real, imag} */,
  {32'h3e96188b, 32'h00000000} /* (6, 11, 11) {real, imag} */,
  {32'hbed4394e, 32'h00000000} /* (6, 11, 10) {real, imag} */,
  {32'hbf7178d3, 32'h00000000} /* (6, 11, 9) {real, imag} */,
  {32'hbf7d86c5, 32'h00000000} /* (6, 11, 8) {real, imag} */,
  {32'hbf0b36c7, 32'h00000000} /* (6, 11, 7) {real, imag} */,
  {32'hbf89147d, 32'h00000000} /* (6, 11, 6) {real, imag} */,
  {32'hbfa27cb1, 32'h00000000} /* (6, 11, 5) {real, imag} */,
  {32'hbf67b2e9, 32'h00000000} /* (6, 11, 4) {real, imag} */,
  {32'hbf047179, 32'h00000000} /* (6, 11, 3) {real, imag} */,
  {32'hbf682d4b, 32'h00000000} /* (6, 11, 2) {real, imag} */,
  {32'hbf0a5e57, 32'h00000000} /* (6, 11, 1) {real, imag} */,
  {32'hbdab4c33, 32'h00000000} /* (6, 11, 0) {real, imag} */,
  {32'h3ea3f378, 32'h00000000} /* (6, 10, 31) {real, imag} */,
  {32'h3eeaa860, 32'h00000000} /* (6, 10, 30) {real, imag} */,
  {32'h3e8a1227, 32'h00000000} /* (6, 10, 29) {real, imag} */,
  {32'h3f3a8aee, 32'h00000000} /* (6, 10, 28) {real, imag} */,
  {32'h3f2990a3, 32'h00000000} /* (6, 10, 27) {real, imag} */,
  {32'h3ddd4123, 32'h00000000} /* (6, 10, 26) {real, imag} */,
  {32'h3ec9ac45, 32'h00000000} /* (6, 10, 25) {real, imag} */,
  {32'h3f1a2fdb, 32'h00000000} /* (6, 10, 24) {real, imag} */,
  {32'h3f2bf90c, 32'h00000000} /* (6, 10, 23) {real, imag} */,
  {32'h3f137e36, 32'h00000000} /* (6, 10, 22) {real, imag} */,
  {32'h3df698e4, 32'h00000000} /* (6, 10, 21) {real, imag} */,
  {32'hbefe2870, 32'h00000000} /* (6, 10, 20) {real, imag} */,
  {32'hbf2c1363, 32'h00000000} /* (6, 10, 19) {real, imag} */,
  {32'hbe669860, 32'h00000000} /* (6, 10, 18) {real, imag} */,
  {32'hbf22aec0, 32'h00000000} /* (6, 10, 17) {real, imag} */,
  {32'hbf03aa7f, 32'h00000000} /* (6, 10, 16) {real, imag} */,
  {32'hbc42b850, 32'h00000000} /* (6, 10, 15) {real, imag} */,
  {32'h3e18148a, 32'h00000000} /* (6, 10, 14) {real, imag} */,
  {32'hbcdea2a2, 32'h00000000} /* (6, 10, 13) {real, imag} */,
  {32'hbedd464a, 32'h00000000} /* (6, 10, 12) {real, imag} */,
  {32'hbf221cd8, 32'h00000000} /* (6, 10, 11) {real, imag} */,
  {32'hbed2b596, 32'h00000000} /* (6, 10, 10) {real, imag} */,
  {32'hbc8eec38, 32'h00000000} /* (6, 10, 9) {real, imag} */,
  {32'h3e240602, 32'h00000000} /* (6, 10, 8) {real, imag} */,
  {32'h3f3fc870, 32'h00000000} /* (6, 10, 7) {real, imag} */,
  {32'h3e61669c, 32'h00000000} /* (6, 10, 6) {real, imag} */,
  {32'h3e236729, 32'h00000000} /* (6, 10, 5) {real, imag} */,
  {32'h3e290a43, 32'h00000000} /* (6, 10, 4) {real, imag} */,
  {32'h3da33afb, 32'h00000000} /* (6, 10, 3) {real, imag} */,
  {32'hbe3aa8d2, 32'h00000000} /* (6, 10, 2) {real, imag} */,
  {32'h3ea2b0ba, 32'h00000000} /* (6, 10, 1) {real, imag} */,
  {32'h3efa7650, 32'h00000000} /* (6, 10, 0) {real, imag} */,
  {32'h3f1bebd4, 32'h00000000} /* (6, 9, 31) {real, imag} */,
  {32'h3f9eb0ed, 32'h00000000} /* (6, 9, 30) {real, imag} */,
  {32'h3f4c066f, 32'h00000000} /* (6, 9, 29) {real, imag} */,
  {32'h3f414eae, 32'h00000000} /* (6, 9, 28) {real, imag} */,
  {32'h3fb60cb1, 32'h00000000} /* (6, 9, 27) {real, imag} */,
  {32'h3f75e920, 32'h00000000} /* (6, 9, 26) {real, imag} */,
  {32'h3f5f64b4, 32'h00000000} /* (6, 9, 25) {real, imag} */,
  {32'h3f447003, 32'h00000000} /* (6, 9, 24) {real, imag} */,
  {32'h3fc0d7a6, 32'h00000000} /* (6, 9, 23) {real, imag} */,
  {32'h3fd51bc9, 32'h00000000} /* (6, 9, 22) {real, imag} */,
  {32'h3f596038, 32'h00000000} /* (6, 9, 21) {real, imag} */,
  {32'hbf6b7807, 32'h00000000} /* (6, 9, 20) {real, imag} */,
  {32'hbf5045f2, 32'h00000000} /* (6, 9, 19) {real, imag} */,
  {32'hbf02b463, 32'h00000000} /* (6, 9, 18) {real, imag} */,
  {32'hbfa1572c, 32'h00000000} /* (6, 9, 17) {real, imag} */,
  {32'hbf62550a, 32'h00000000} /* (6, 9, 16) {real, imag} */,
  {32'hbe17d7cd, 32'h00000000} /* (6, 9, 15) {real, imag} */,
  {32'hbea3f9f0, 32'h00000000} /* (6, 9, 14) {real, imag} */,
  {32'hbea40774, 32'h00000000} /* (6, 9, 13) {real, imag} */,
  {32'hbeb62bc2, 32'h00000000} /* (6, 9, 12) {real, imag} */,
  {32'hbf4ee40d, 32'h00000000} /* (6, 9, 11) {real, imag} */,
  {32'hbec71f3c, 32'h00000000} /* (6, 9, 10) {real, imag} */,
  {32'h3e6d1ac3, 32'h00000000} /* (6, 9, 9) {real, imag} */,
  {32'h3f80d8fd, 32'h00000000} /* (6, 9, 8) {real, imag} */,
  {32'h3fdb7161, 32'h00000000} /* (6, 9, 7) {real, imag} */,
  {32'h3f2f001e, 32'h00000000} /* (6, 9, 6) {real, imag} */,
  {32'h3eb8fb23, 32'h00000000} /* (6, 9, 5) {real, imag} */,
  {32'h3f192045, 32'h00000000} /* (6, 9, 4) {real, imag} */,
  {32'h3f65c041, 32'h00000000} /* (6, 9, 3) {real, imag} */,
  {32'h3f624219, 32'h00000000} /* (6, 9, 2) {real, imag} */,
  {32'h3f45b3c1, 32'h00000000} /* (6, 9, 1) {real, imag} */,
  {32'h3eee98ba, 32'h00000000} /* (6, 9, 0) {real, imag} */,
  {32'h3ef76735, 32'h00000000} /* (6, 8, 31) {real, imag} */,
  {32'h3f96f925, 32'h00000000} /* (6, 8, 30) {real, imag} */,
  {32'h3f267c82, 32'h00000000} /* (6, 8, 29) {real, imag} */,
  {32'h3e437d50, 32'h00000000} /* (6, 8, 28) {real, imag} */,
  {32'h3f18fda9, 32'h00000000} /* (6, 8, 27) {real, imag} */,
  {32'h3f1c07a5, 32'h00000000} /* (6, 8, 26) {real, imag} */,
  {32'h3d8a14ce, 32'h00000000} /* (6, 8, 25) {real, imag} */,
  {32'h3ec45a05, 32'h00000000} /* (6, 8, 24) {real, imag} */,
  {32'h3f901c2b, 32'h00000000} /* (6, 8, 23) {real, imag} */,
  {32'h3fa1976b, 32'h00000000} /* (6, 8, 22) {real, imag} */,
  {32'h3ef6a1d6, 32'h00000000} /* (6, 8, 21) {real, imag} */,
  {32'hbf0856e8, 32'h00000000} /* (6, 8, 20) {real, imag} */,
  {32'hbefe532d, 32'h00000000} /* (6, 8, 19) {real, imag} */,
  {32'hbed02b82, 32'h00000000} /* (6, 8, 18) {real, imag} */,
  {32'hbf54f502, 32'h00000000} /* (6, 8, 17) {real, imag} */,
  {32'hbf84953f, 32'h00000000} /* (6, 8, 16) {real, imag} */,
  {32'hbf0f287e, 32'h00000000} /* (6, 8, 15) {real, imag} */,
  {32'hbf4466d4, 32'h00000000} /* (6, 8, 14) {real, imag} */,
  {32'hbf5ad5fb, 32'h00000000} /* (6, 8, 13) {real, imag} */,
  {32'hbed1c8e9, 32'h00000000} /* (6, 8, 12) {real, imag} */,
  {32'hbeb9c8ba, 32'h00000000} /* (6, 8, 11) {real, imag} */,
  {32'h3c6db142, 32'h00000000} /* (6, 8, 10) {real, imag} */,
  {32'h3e31b258, 32'h00000000} /* (6, 8, 9) {real, imag} */,
  {32'h3f6fb1c6, 32'h00000000} /* (6, 8, 8) {real, imag} */,
  {32'h3f92dd6c, 32'h00000000} /* (6, 8, 7) {real, imag} */,
  {32'h3ef80999, 32'h00000000} /* (6, 8, 6) {real, imag} */,
  {32'h3e078645, 32'h00000000} /* (6, 8, 5) {real, imag} */,
  {32'h3f2048b1, 32'h00000000} /* (6, 8, 4) {real, imag} */,
  {32'h3fa2a212, 32'h00000000} /* (6, 8, 3) {real, imag} */,
  {32'h3f8f7e74, 32'h00000000} /* (6, 8, 2) {real, imag} */,
  {32'h3f47a21d, 32'h00000000} /* (6, 8, 1) {real, imag} */,
  {32'h3f074b19, 32'h00000000} /* (6, 8, 0) {real, imag} */,
  {32'h3f350624, 32'h00000000} /* (6, 7, 31) {real, imag} */,
  {32'h3f5e62e7, 32'h00000000} /* (6, 7, 30) {real, imag} */,
  {32'h3e8ebce5, 32'h00000000} /* (6, 7, 29) {real, imag} */,
  {32'h3dc8c838, 32'h00000000} /* (6, 7, 28) {real, imag} */,
  {32'h3ea671c7, 32'h00000000} /* (6, 7, 27) {real, imag} */,
  {32'h3ef33ee1, 32'h00000000} /* (6, 7, 26) {real, imag} */,
  {32'hbc50c2b2, 32'h00000000} /* (6, 7, 25) {real, imag} */,
  {32'h3f0076cd, 32'h00000000} /* (6, 7, 24) {real, imag} */,
  {32'h3f6ead00, 32'h00000000} /* (6, 7, 23) {real, imag} */,
  {32'h3f9520ac, 32'h00000000} /* (6, 7, 22) {real, imag} */,
  {32'h3f15c79a, 32'h00000000} /* (6, 7, 21) {real, imag} */,
  {32'hbe3481bb, 32'h00000000} /* (6, 7, 20) {real, imag} */,
  {32'hbece2bb8, 32'h00000000} /* (6, 7, 19) {real, imag} */,
  {32'hbedd63e7, 32'h00000000} /* (6, 7, 18) {real, imag} */,
  {32'hbf251516, 32'h00000000} /* (6, 7, 17) {real, imag} */,
  {32'hbf86c3bd, 32'h00000000} /* (6, 7, 16) {real, imag} */,
  {32'hbf9cd5ce, 32'h00000000} /* (6, 7, 15) {real, imag} */,
  {32'hbfa78e71, 32'h00000000} /* (6, 7, 14) {real, imag} */,
  {32'hbfade795, 32'h00000000} /* (6, 7, 13) {real, imag} */,
  {32'hbf5844a3, 32'h00000000} /* (6, 7, 12) {real, imag} */,
  {32'hbe9b955b, 32'h00000000} /* (6, 7, 11) {real, imag} */,
  {32'h3e56ab0a, 32'h00000000} /* (6, 7, 10) {real, imag} */,
  {32'h3ec4a263, 32'h00000000} /* (6, 7, 9) {real, imag} */,
  {32'h3f751df5, 32'h00000000} /* (6, 7, 8) {real, imag} */,
  {32'h3ece41a9, 32'h00000000} /* (6, 7, 7) {real, imag} */,
  {32'h3edf5a7d, 32'h00000000} /* (6, 7, 6) {real, imag} */,
  {32'h3f3e52c3, 32'h00000000} /* (6, 7, 5) {real, imag} */,
  {32'h3f5ae5cc, 32'h00000000} /* (6, 7, 4) {real, imag} */,
  {32'h3f8cdb80, 32'h00000000} /* (6, 7, 3) {real, imag} */,
  {32'h3f9a6ceb, 32'h00000000} /* (6, 7, 2) {real, imag} */,
  {32'h3f103a8b, 32'h00000000} /* (6, 7, 1) {real, imag} */,
  {32'h3eb16be2, 32'h00000000} /* (6, 7, 0) {real, imag} */,
  {32'h3f0e4740, 32'h00000000} /* (6, 6, 31) {real, imag} */,
  {32'h3f706a95, 32'h00000000} /* (6, 6, 30) {real, imag} */,
  {32'h3f1b0c96, 32'h00000000} /* (6, 6, 29) {real, imag} */,
  {32'h3ec16557, 32'h00000000} /* (6, 6, 28) {real, imag} */,
  {32'h3f63b5ca, 32'h00000000} /* (6, 6, 27) {real, imag} */,
  {32'h3f418845, 32'h00000000} /* (6, 6, 26) {real, imag} */,
  {32'h3efeee83, 32'h00000000} /* (6, 6, 25) {real, imag} */,
  {32'h3f48772c, 32'h00000000} /* (6, 6, 24) {real, imag} */,
  {32'h3f40b626, 32'h00000000} /* (6, 6, 23) {real, imag} */,
  {32'h3f7e3ee1, 32'h00000000} /* (6, 6, 22) {real, imag} */,
  {32'h3eddde0d, 32'h00000000} /* (6, 6, 21) {real, imag} */,
  {32'hbf3fe625, 32'h00000000} /* (6, 6, 20) {real, imag} */,
  {32'hbf121273, 32'h00000000} /* (6, 6, 19) {real, imag} */,
  {32'hbf28d84a, 32'h00000000} /* (6, 6, 18) {real, imag} */,
  {32'hbf3d50cf, 32'h00000000} /* (6, 6, 17) {real, imag} */,
  {32'hbf126309, 32'h00000000} /* (6, 6, 16) {real, imag} */,
  {32'hbf5af3f1, 32'h00000000} /* (6, 6, 15) {real, imag} */,
  {32'hbf11dbf7, 32'h00000000} /* (6, 6, 14) {real, imag} */,
  {32'hbf046658, 32'h00000000} /* (6, 6, 13) {real, imag} */,
  {32'hbf6f91e3, 32'h00000000} /* (6, 6, 12) {real, imag} */,
  {32'hbf088304, 32'h00000000} /* (6, 6, 11) {real, imag} */,
  {32'h3f29a52c, 32'h00000000} /* (6, 6, 10) {real, imag} */,
  {32'h3f45063c, 32'h00000000} /* (6, 6, 9) {real, imag} */,
  {32'h3f7714ad, 32'h00000000} /* (6, 6, 8) {real, imag} */,
  {32'h3f2356a0, 32'h00000000} /* (6, 6, 7) {real, imag} */,
  {32'h3fa0543c, 32'h00000000} /* (6, 6, 6) {real, imag} */,
  {32'h3ffb1886, 32'h00000000} /* (6, 6, 5) {real, imag} */,
  {32'h3fbc0023, 32'h00000000} /* (6, 6, 4) {real, imag} */,
  {32'h3f2a45fc, 32'h00000000} /* (6, 6, 3) {real, imag} */,
  {32'h3f68aa11, 32'h00000000} /* (6, 6, 2) {real, imag} */,
  {32'h3f48fc63, 32'h00000000} /* (6, 6, 1) {real, imag} */,
  {32'h3eb96759, 32'h00000000} /* (6, 6, 0) {real, imag} */,
  {32'h3f805387, 32'h00000000} /* (6, 5, 31) {real, imag} */,
  {32'h3f1d2af4, 32'h00000000} /* (6, 5, 30) {real, imag} */,
  {32'h3ed69439, 32'h00000000} /* (6, 5, 29) {real, imag} */,
  {32'h3f2f270b, 32'h00000000} /* (6, 5, 28) {real, imag} */,
  {32'h3f71e44e, 32'h00000000} /* (6, 5, 27) {real, imag} */,
  {32'h3f341f2d, 32'h00000000} /* (6, 5, 26) {real, imag} */,
  {32'h3f1f887c, 32'h00000000} /* (6, 5, 25) {real, imag} */,
  {32'h3f36f0ac, 32'h00000000} /* (6, 5, 24) {real, imag} */,
  {32'h3f84fdfb, 32'h00000000} /* (6, 5, 23) {real, imag} */,
  {32'h3f5fcf76, 32'h00000000} /* (6, 5, 22) {real, imag} */,
  {32'h3ec2ac84, 32'h00000000} /* (6, 5, 21) {real, imag} */,
  {32'hbd962fb2, 32'h00000000} /* (6, 5, 20) {real, imag} */,
  {32'h3e03ba24, 32'h00000000} /* (6, 5, 19) {real, imag} */,
  {32'h3be3c9f7, 32'h00000000} /* (6, 5, 18) {real, imag} */,
  {32'h3d3ebf81, 32'h00000000} /* (6, 5, 17) {real, imag} */,
  {32'h3e323827, 32'h00000000} /* (6, 5, 16) {real, imag} */,
  {32'hbf63f128, 32'h00000000} /* (6, 5, 15) {real, imag} */,
  {32'hbf80f01e, 32'h00000000} /* (6, 5, 14) {real, imag} */,
  {32'hbf0370e7, 32'h00000000} /* (6, 5, 13) {real, imag} */,
  {32'hbf4e848e, 32'h00000000} /* (6, 5, 12) {real, imag} */,
  {32'hbf96e6fa, 32'h00000000} /* (6, 5, 11) {real, imag} */,
  {32'hbdfbcb78, 32'h00000000} /* (6, 5, 10) {real, imag} */,
  {32'hbe2fbc28, 32'h00000000} /* (6, 5, 9) {real, imag} */,
  {32'hbf4717c1, 32'h00000000} /* (6, 5, 8) {real, imag} */,
  {32'hbeb7c5bf, 32'h00000000} /* (6, 5, 7) {real, imag} */,
  {32'h3e616db8, 32'h00000000} /* (6, 5, 6) {real, imag} */,
  {32'h3f447b00, 32'h00000000} /* (6, 5, 5) {real, imag} */,
  {32'h3f952ad3, 32'h00000000} /* (6, 5, 4) {real, imag} */,
  {32'h3f3c4c7a, 32'h00000000} /* (6, 5, 3) {real, imag} */,
  {32'h3f0d49af, 32'h00000000} /* (6, 5, 2) {real, imag} */,
  {32'h3f381bf9, 32'h00000000} /* (6, 5, 1) {real, imag} */,
  {32'h3ec2babe, 32'h00000000} /* (6, 5, 0) {real, imag} */,
  {32'h3f25782d, 32'h00000000} /* (6, 4, 31) {real, imag} */,
  {32'h3eac0ead, 32'h00000000} /* (6, 4, 30) {real, imag} */,
  {32'h3dc5a0bb, 32'h00000000} /* (6, 4, 29) {real, imag} */,
  {32'h3f0e304c, 32'h00000000} /* (6, 4, 28) {real, imag} */,
  {32'h3f2a532e, 32'h00000000} /* (6, 4, 27) {real, imag} */,
  {32'h3f20707f, 32'h00000000} /* (6, 4, 26) {real, imag} */,
  {32'h3ed82b40, 32'h00000000} /* (6, 4, 25) {real, imag} */,
  {32'h3ed9506a, 32'h00000000} /* (6, 4, 24) {real, imag} */,
  {32'h3f3f1e6f, 32'h00000000} /* (6, 4, 23) {real, imag} */,
  {32'h3f3a55c6, 32'h00000000} /* (6, 4, 22) {real, imag} */,
  {32'h3ef4bba6, 32'h00000000} /* (6, 4, 21) {real, imag} */,
  {32'h3f628211, 32'h00000000} /* (6, 4, 20) {real, imag} */,
  {32'h3f4132a3, 32'h00000000} /* (6, 4, 19) {real, imag} */,
  {32'h3f86ed18, 32'h00000000} /* (6, 4, 18) {real, imag} */,
  {32'h3f659eac, 32'h00000000} /* (6, 4, 17) {real, imag} */,
  {32'h3e34eb52, 32'h00000000} /* (6, 4, 16) {real, imag} */,
  {32'hbfda23a2, 32'h00000000} /* (6, 4, 15) {real, imag} */,
  {32'hbfd6624c, 32'h00000000} /* (6, 4, 14) {real, imag} */,
  {32'hbf3e5239, 32'h00000000} /* (6, 4, 13) {real, imag} */,
  {32'hbf865477, 32'h00000000} /* (6, 4, 12) {real, imag} */,
  {32'hbf8d4c3e, 32'h00000000} /* (6, 4, 11) {real, imag} */,
  {32'hbf2b6d06, 32'h00000000} /* (6, 4, 10) {real, imag} */,
  {32'hbf310f50, 32'h00000000} /* (6, 4, 9) {real, imag} */,
  {32'hbfb2b740, 32'h00000000} /* (6, 4, 8) {real, imag} */,
  {32'hbf934c4e, 32'h00000000} /* (6, 4, 7) {real, imag} */,
  {32'hbf667541, 32'h00000000} /* (6, 4, 6) {real, imag} */,
  {32'hbe381ac7, 32'h00000000} /* (6, 4, 5) {real, imag} */,
  {32'h3f4e85fa, 32'h00000000} /* (6, 4, 4) {real, imag} */,
  {32'h3f5167ec, 32'h00000000} /* (6, 4, 3) {real, imag} */,
  {32'h3f05673c, 32'h00000000} /* (6, 4, 2) {real, imag} */,
  {32'h3fb0761c, 32'h00000000} /* (6, 4, 1) {real, imag} */,
  {32'h3f5b330b, 32'h00000000} /* (6, 4, 0) {real, imag} */,
  {32'h3edd9048, 32'h00000000} /* (6, 3, 31) {real, imag} */,
  {32'h3f2702b5, 32'h00000000} /* (6, 3, 30) {real, imag} */,
  {32'h3ebec25c, 32'h00000000} /* (6, 3, 29) {real, imag} */,
  {32'h3f4d463e, 32'h00000000} /* (6, 3, 28) {real, imag} */,
  {32'h3f43beeb, 32'h00000000} /* (6, 3, 27) {real, imag} */,
  {32'h3f090eb6, 32'h00000000} /* (6, 3, 26) {real, imag} */,
  {32'h3f810081, 32'h00000000} /* (6, 3, 25) {real, imag} */,
  {32'h3f8a7035, 32'h00000000} /* (6, 3, 24) {real, imag} */,
  {32'h3f0d1c99, 32'h00000000} /* (6, 3, 23) {real, imag} */,
  {32'h3f54fce9, 32'h00000000} /* (6, 3, 22) {real, imag} */,
  {32'h3f303651, 32'h00000000} /* (6, 3, 21) {real, imag} */,
  {32'h3f303a6c, 32'h00000000} /* (6, 3, 20) {real, imag} */,
  {32'h3f388071, 32'h00000000} /* (6, 3, 19) {real, imag} */,
  {32'h3f8761a7, 32'h00000000} /* (6, 3, 18) {real, imag} */,
  {32'h3f6abd54, 32'h00000000} /* (6, 3, 17) {real, imag} */,
  {32'h3e9e6201, 32'h00000000} /* (6, 3, 16) {real, imag} */,
  {32'hbf345787, 32'h00000000} /* (6, 3, 15) {real, imag} */,
  {32'hbfa9698f, 32'h00000000} /* (6, 3, 14) {real, imag} */,
  {32'hbf40de38, 32'h00000000} /* (6, 3, 13) {real, imag} */,
  {32'hbf75b46e, 32'h00000000} /* (6, 3, 12) {real, imag} */,
  {32'hbf702372, 32'h00000000} /* (6, 3, 11) {real, imag} */,
  {32'hbf3c5c20, 32'h00000000} /* (6, 3, 10) {real, imag} */,
  {32'hbf5f96c7, 32'h00000000} /* (6, 3, 9) {real, imag} */,
  {32'hbf84208c, 32'h00000000} /* (6, 3, 8) {real, imag} */,
  {32'hbf88dcd5, 32'h00000000} /* (6, 3, 7) {real, imag} */,
  {32'hbf9b741a, 32'h00000000} /* (6, 3, 6) {real, imag} */,
  {32'hbecf2f33, 32'h00000000} /* (6, 3, 5) {real, imag} */,
  {32'h3f0a7b04, 32'h00000000} /* (6, 3, 4) {real, imag} */,
  {32'h3f2a7f4f, 32'h00000000} /* (6, 3, 3) {real, imag} */,
  {32'h3ebf25ce, 32'h00000000} /* (6, 3, 2) {real, imag} */,
  {32'h3f6a09f0, 32'h00000000} /* (6, 3, 1) {real, imag} */,
  {32'h3f5ce08d, 32'h00000000} /* (6, 3, 0) {real, imag} */,
  {32'h3eed5793, 32'h00000000} /* (6, 2, 31) {real, imag} */,
  {32'h3f6d03b2, 32'h00000000} /* (6, 2, 30) {real, imag} */,
  {32'h3f2c758d, 32'h00000000} /* (6, 2, 29) {real, imag} */,
  {32'h3f7428db, 32'h00000000} /* (6, 2, 28) {real, imag} */,
  {32'h3f6558f4, 32'h00000000} /* (6, 2, 27) {real, imag} */,
  {32'h3ed02c80, 32'h00000000} /* (6, 2, 26) {real, imag} */,
  {32'h3f8b591d, 32'h00000000} /* (6, 2, 25) {real, imag} */,
  {32'h3f94e669, 32'h00000000} /* (6, 2, 24) {real, imag} */,
  {32'h3f2cf7e6, 32'h00000000} /* (6, 2, 23) {real, imag} */,
  {32'h3fd6f927, 32'h00000000} /* (6, 2, 22) {real, imag} */,
  {32'h3fbf0eeb, 32'h00000000} /* (6, 2, 21) {real, imag} */,
  {32'h3f83c968, 32'h00000000} /* (6, 2, 20) {real, imag} */,
  {32'h3f589f9e, 32'h00000000} /* (6, 2, 19) {real, imag} */,
  {32'h3f90d632, 32'h00000000} /* (6, 2, 18) {real, imag} */,
  {32'h3fa5a457, 32'h00000000} /* (6, 2, 17) {real, imag} */,
  {32'h3f654dd6, 32'h00000000} /* (6, 2, 16) {real, imag} */,
  {32'h3b512a1e, 32'h00000000} /* (6, 2, 15) {real, imag} */,
  {32'hbf0f9db7, 32'h00000000} /* (6, 2, 14) {real, imag} */,
  {32'hbea6a309, 32'h00000000} /* (6, 2, 13) {real, imag} */,
  {32'hbefd0227, 32'h00000000} /* (6, 2, 12) {real, imag} */,
  {32'hbf4e662a, 32'h00000000} /* (6, 2, 11) {real, imag} */,
  {32'hbf4c9537, 32'h00000000} /* (6, 2, 10) {real, imag} */,
  {32'hbeb77143, 32'h00000000} /* (6, 2, 9) {real, imag} */,
  {32'hbf35b967, 32'h00000000} /* (6, 2, 8) {real, imag} */,
  {32'hbf58e2bb, 32'h00000000} /* (6, 2, 7) {real, imag} */,
  {32'hbf2baf93, 32'h00000000} /* (6, 2, 6) {real, imag} */,
  {32'hbdebc989, 32'h00000000} /* (6, 2, 5) {real, imag} */,
  {32'h3e34f44c, 32'h00000000} /* (6, 2, 4) {real, imag} */,
  {32'h3f2d231e, 32'h00000000} /* (6, 2, 3) {real, imag} */,
  {32'h3f5d42d4, 32'h00000000} /* (6, 2, 2) {real, imag} */,
  {32'h3f23458c, 32'h00000000} /* (6, 2, 1) {real, imag} */,
  {32'h3f2567e3, 32'h00000000} /* (6, 2, 0) {real, imag} */,
  {32'h3e792f01, 32'h00000000} /* (6, 1, 31) {real, imag} */,
  {32'h3efdabac, 32'h00000000} /* (6, 1, 30) {real, imag} */,
  {32'h3f1d61a0, 32'h00000000} /* (6, 1, 29) {real, imag} */,
  {32'h3f57b84f, 32'h00000000} /* (6, 1, 28) {real, imag} */,
  {32'h3f69c71a, 32'h00000000} /* (6, 1, 27) {real, imag} */,
  {32'h3e6a4647, 32'h00000000} /* (6, 1, 26) {real, imag} */,
  {32'h3f1ab254, 32'h00000000} /* (6, 1, 25) {real, imag} */,
  {32'h3f1e0f32, 32'h00000000} /* (6, 1, 24) {real, imag} */,
  {32'h3eed8fcc, 32'h00000000} /* (6, 1, 23) {real, imag} */,
  {32'h3f1d8d0c, 32'h00000000} /* (6, 1, 22) {real, imag} */,
  {32'h3f645e39, 32'h00000000} /* (6, 1, 21) {real, imag} */,
  {32'h3f1bb61a, 32'h00000000} /* (6, 1, 20) {real, imag} */,
  {32'h3e8d6ec0, 32'h00000000} /* (6, 1, 19) {real, imag} */,
  {32'h3f4af993, 32'h00000000} /* (6, 1, 18) {real, imag} */,
  {32'h3f5c5a50, 32'h00000000} /* (6, 1, 17) {real, imag} */,
  {32'h3f15fa3b, 32'h00000000} /* (6, 1, 16) {real, imag} */,
  {32'h3e1ba244, 32'h00000000} /* (6, 1, 15) {real, imag} */,
  {32'h3e81f132, 32'h00000000} /* (6, 1, 14) {real, imag} */,
  {32'hbea375f3, 32'h00000000} /* (6, 1, 13) {real, imag} */,
  {32'hbf25df06, 32'h00000000} /* (6, 1, 12) {real, imag} */,
  {32'hbf657f85, 32'h00000000} /* (6, 1, 11) {real, imag} */,
  {32'hbf32de93, 32'h00000000} /* (6, 1, 10) {real, imag} */,
  {32'hbed159d3, 32'h00000000} /* (6, 1, 9) {real, imag} */,
  {32'hbf1841dc, 32'h00000000} /* (6, 1, 8) {real, imag} */,
  {32'hbf247241, 32'h00000000} /* (6, 1, 7) {real, imag} */,
  {32'hbf0a3bdf, 32'h00000000} /* (6, 1, 6) {real, imag} */,
  {32'hbd8b4623, 32'h00000000} /* (6, 1, 5) {real, imag} */,
  {32'h3e64eba2, 32'h00000000} /* (6, 1, 4) {real, imag} */,
  {32'h3f11ffc0, 32'h00000000} /* (6, 1, 3) {real, imag} */,
  {32'h3e913385, 32'h00000000} /* (6, 1, 2) {real, imag} */,
  {32'h3ea6f798, 32'h00000000} /* (6, 1, 1) {real, imag} */,
  {32'h3e5c87b1, 32'h00000000} /* (6, 1, 0) {real, imag} */,
  {32'h3ecab1f4, 32'h00000000} /* (6, 0, 31) {real, imag} */,
  {32'h3ed558dd, 32'h00000000} /* (6, 0, 30) {real, imag} */,
  {32'h3e521ad1, 32'h00000000} /* (6, 0, 29) {real, imag} */,
  {32'h3eda4d28, 32'h00000000} /* (6, 0, 28) {real, imag} */,
  {32'h3f92e542, 32'h00000000} /* (6, 0, 27) {real, imag} */,
  {32'h3ee04029, 32'h00000000} /* (6, 0, 26) {real, imag} */,
  {32'h3ef889cd, 32'h00000000} /* (6, 0, 25) {real, imag} */,
  {32'h3e925ae0, 32'h00000000} /* (6, 0, 24) {real, imag} */,
  {32'h3e0e2f81, 32'h00000000} /* (6, 0, 23) {real, imag} */,
  {32'h3dd21b64, 32'h00000000} /* (6, 0, 22) {real, imag} */,
  {32'h3f0cf5af, 32'h00000000} /* (6, 0, 21) {real, imag} */,
  {32'h3ee9513b, 32'h00000000} /* (6, 0, 20) {real, imag} */,
  {32'h3dedbf06, 32'h00000000} /* (6, 0, 19) {real, imag} */,
  {32'h3e87374d, 32'h00000000} /* (6, 0, 18) {real, imag} */,
  {32'h3e86b83a, 32'h00000000} /* (6, 0, 17) {real, imag} */,
  {32'h3ca7998c, 32'h00000000} /* (6, 0, 16) {real, imag} */,
  {32'hbe1b0a7c, 32'h00000000} /* (6, 0, 15) {real, imag} */,
  {32'h3c1daf69, 32'h00000000} /* (6, 0, 14) {real, imag} */,
  {32'hbebab57e, 32'h00000000} /* (6, 0, 13) {real, imag} */,
  {32'hbf2440e7, 32'h00000000} /* (6, 0, 12) {real, imag} */,
  {32'hbef6782d, 32'h00000000} /* (6, 0, 11) {real, imag} */,
  {32'hbe03f6b4, 32'h00000000} /* (6, 0, 10) {real, imag} */,
  {32'hbea6d7d8, 32'h00000000} /* (6, 0, 9) {real, imag} */,
  {32'hbe9f981f, 32'h00000000} /* (6, 0, 8) {real, imag} */,
  {32'hbf0331da, 32'h00000000} /* (6, 0, 7) {real, imag} */,
  {32'hbeaf4f14, 32'h00000000} /* (6, 0, 6) {real, imag} */,
  {32'h3e5bac19, 32'h00000000} /* (6, 0, 5) {real, imag} */,
  {32'h3ec626d5, 32'h00000000} /* (6, 0, 4) {real, imag} */,
  {32'h3f12241d, 32'h00000000} /* (6, 0, 3) {real, imag} */,
  {32'h3e122d9e, 32'h00000000} /* (6, 0, 2) {real, imag} */,
  {32'h3df231d9, 32'h00000000} /* (6, 0, 1) {real, imag} */,
  {32'h3e1a5310, 32'h00000000} /* (6, 0, 0) {real, imag} */,
  {32'hbd90507f, 32'h00000000} /* (5, 31, 31) {real, imag} */,
  {32'h3e59d4d7, 32'h00000000} /* (5, 31, 30) {real, imag} */,
  {32'h3e2de9ac, 32'h00000000} /* (5, 31, 29) {real, imag} */,
  {32'h3e1a3de3, 32'h00000000} /* (5, 31, 28) {real, imag} */,
  {32'h3c0de180, 32'h00000000} /* (5, 31, 27) {real, imag} */,
  {32'hbe8acc13, 32'h00000000} /* (5, 31, 26) {real, imag} */,
  {32'h3d04f58c, 32'h00000000} /* (5, 31, 25) {real, imag} */,
  {32'hbd9913b0, 32'h00000000} /* (5, 31, 24) {real, imag} */,
  {32'hbde92b16, 32'h00000000} /* (5, 31, 23) {real, imag} */,
  {32'hbe4a5986, 32'h00000000} /* (5, 31, 22) {real, imag} */,
  {32'h3e0df30a, 32'h00000000} /* (5, 31, 21) {real, imag} */,
  {32'hbda95652, 32'h00000000} /* (5, 31, 20) {real, imag} */,
  {32'h3b5195a9, 32'h00000000} /* (5, 31, 19) {real, imag} */,
  {32'h3dd3d425, 32'h00000000} /* (5, 31, 18) {real, imag} */,
  {32'h3bf96670, 32'h00000000} /* (5, 31, 17) {real, imag} */,
  {32'hbb330207, 32'h00000000} /* (5, 31, 16) {real, imag} */,
  {32'h3d8e3a4e, 32'h00000000} /* (5, 31, 15) {real, imag} */,
  {32'hbe9e1034, 32'h00000000} /* (5, 31, 14) {real, imag} */,
  {32'h3e184709, 32'h00000000} /* (5, 31, 13) {real, imag} */,
  {32'h3e3b585a, 32'h00000000} /* (5, 31, 12) {real, imag} */,
  {32'h3e1cb724, 32'h00000000} /* (5, 31, 11) {real, imag} */,
  {32'h3e80e656, 32'h00000000} /* (5, 31, 10) {real, imag} */,
  {32'hbe0a637f, 32'h00000000} /* (5, 31, 9) {real, imag} */,
  {32'hbd857c43, 32'h00000000} /* (5, 31, 8) {real, imag} */,
  {32'hbcbc4501, 32'h00000000} /* (5, 31, 7) {real, imag} */,
  {32'hbeabec57, 32'h00000000} /* (5, 31, 6) {real, imag} */,
  {32'hbeb46b2d, 32'h00000000} /* (5, 31, 5) {real, imag} */,
  {32'hbf057ce5, 32'h00000000} /* (5, 31, 4) {real, imag} */,
  {32'hbf2000c3, 32'h00000000} /* (5, 31, 3) {real, imag} */,
  {32'hbee6753e, 32'h00000000} /* (5, 31, 2) {real, imag} */,
  {32'h3daf8a0b, 32'h00000000} /* (5, 31, 1) {real, imag} */,
  {32'h3df7caed, 32'h00000000} /* (5, 31, 0) {real, imag} */,
  {32'h3dd06bf9, 32'h00000000} /* (5, 30, 31) {real, imag} */,
  {32'h3ed49cef, 32'h00000000} /* (5, 30, 30) {real, imag} */,
  {32'h3e8e752d, 32'h00000000} /* (5, 30, 29) {real, imag} */,
  {32'h3e2b41d2, 32'h00000000} /* (5, 30, 28) {real, imag} */,
  {32'h3e07c6d8, 32'h00000000} /* (5, 30, 27) {real, imag} */,
  {32'hbed3ec17, 32'h00000000} /* (5, 30, 26) {real, imag} */,
  {32'hbebd8b13, 32'h00000000} /* (5, 30, 25) {real, imag} */,
  {32'h3d544292, 32'h00000000} /* (5, 30, 24) {real, imag} */,
  {32'hbe01283f, 32'h00000000} /* (5, 30, 23) {real, imag} */,
  {32'hbecbf801, 32'h00000000} /* (5, 30, 22) {real, imag} */,
  {32'h3eafa658, 32'h00000000} /* (5, 30, 21) {real, imag} */,
  {32'h3df3f870, 32'h00000000} /* (5, 30, 20) {real, imag} */,
  {32'hbdd785d0, 32'h00000000} /* (5, 30, 19) {real, imag} */,
  {32'h3d39207c, 32'h00000000} /* (5, 30, 18) {real, imag} */,
  {32'h3ed99f2d, 32'h00000000} /* (5, 30, 17) {real, imag} */,
  {32'h3e9ca970, 32'h00000000} /* (5, 30, 16) {real, imag} */,
  {32'h3ea2acab, 32'h00000000} /* (5, 30, 15) {real, imag} */,
  {32'hbe8de441, 32'h00000000} /* (5, 30, 14) {real, imag} */,
  {32'h3d38890c, 32'h00000000} /* (5, 30, 13) {real, imag} */,
  {32'h3e891fde, 32'h00000000} /* (5, 30, 12) {real, imag} */,
  {32'h3debc91f, 32'h00000000} /* (5, 30, 11) {real, imag} */,
  {32'hbdd2b8cd, 32'h00000000} /* (5, 30, 10) {real, imag} */,
  {32'hbeb9810f, 32'h00000000} /* (5, 30, 9) {real, imag} */,
  {32'h3e2f9dc4, 32'h00000000} /* (5, 30, 8) {real, imag} */,
  {32'h3e5f0e96, 32'h00000000} /* (5, 30, 7) {real, imag} */,
  {32'hbf81be52, 32'h00000000} /* (5, 30, 6) {real, imag} */,
  {32'hbf91f24f, 32'h00000000} /* (5, 30, 5) {real, imag} */,
  {32'hbf3aaa40, 32'h00000000} /* (5, 30, 4) {real, imag} */,
  {32'hbe058bd4, 32'h00000000} /* (5, 30, 3) {real, imag} */,
  {32'h3e0c4c56, 32'h00000000} /* (5, 30, 2) {real, imag} */,
  {32'h3ea36d0d, 32'h00000000} /* (5, 30, 1) {real, imag} */,
  {32'h3e67914f, 32'h00000000} /* (5, 30, 0) {real, imag} */,
  {32'h3e998f5a, 32'h00000000} /* (5, 29, 31) {real, imag} */,
  {32'hbe4c54ae, 32'h00000000} /* (5, 29, 30) {real, imag} */,
  {32'hbf4bdf84, 32'h00000000} /* (5, 29, 29) {real, imag} */,
  {32'h3d3d7944, 32'h00000000} /* (5, 29, 28) {real, imag} */,
  {32'hbd0dd9ce, 32'h00000000} /* (5, 29, 27) {real, imag} */,
  {32'hbf54576b, 32'h00000000} /* (5, 29, 26) {real, imag} */,
  {32'hbf7bab23, 32'h00000000} /* (5, 29, 25) {real, imag} */,
  {32'hbcc81917, 32'h00000000} /* (5, 29, 24) {real, imag} */,
  {32'hbed1c687, 32'h00000000} /* (5, 29, 23) {real, imag} */,
  {32'hbe9b4ca9, 32'h00000000} /* (5, 29, 22) {real, imag} */,
  {32'h3eae17c1, 32'h00000000} /* (5, 29, 21) {real, imag} */,
  {32'hbe180708, 32'h00000000} /* (5, 29, 20) {real, imag} */,
  {32'hbe8bebb8, 32'h00000000} /* (5, 29, 19) {real, imag} */,
  {32'hbe9c5004, 32'h00000000} /* (5, 29, 18) {real, imag} */,
  {32'h3ed05b72, 32'h00000000} /* (5, 29, 17) {real, imag} */,
  {32'h3f04d07b, 32'h00000000} /* (5, 29, 16) {real, imag} */,
  {32'h3f011700, 32'h00000000} /* (5, 29, 15) {real, imag} */,
  {32'h3e5747f2, 32'h00000000} /* (5, 29, 14) {real, imag} */,
  {32'h3e1570be, 32'h00000000} /* (5, 29, 13) {real, imag} */,
  {32'h3e94c7b5, 32'h00000000} /* (5, 29, 12) {real, imag} */,
  {32'hbe3f8fe3, 32'h00000000} /* (5, 29, 11) {real, imag} */,
  {32'hbeddf9ed, 32'h00000000} /* (5, 29, 10) {real, imag} */,
  {32'hbedf1671, 32'h00000000} /* (5, 29, 9) {real, imag} */,
  {32'h3ee66493, 32'h00000000} /* (5, 29, 8) {real, imag} */,
  {32'h3e3675fa, 32'h00000000} /* (5, 29, 7) {real, imag} */,
  {32'hbf778a75, 32'h00000000} /* (5, 29, 6) {real, imag} */,
  {32'hbf699347, 32'h00000000} /* (5, 29, 5) {real, imag} */,
  {32'hbf2b4a0a, 32'h00000000} /* (5, 29, 4) {real, imag} */,
  {32'hbd6402d1, 32'h00000000} /* (5, 29, 3) {real, imag} */,
  {32'h3d146df5, 32'h00000000} /* (5, 29, 2) {real, imag} */,
  {32'h3e0c9016, 32'h00000000} /* (5, 29, 1) {real, imag} */,
  {32'h3dbd6e42, 32'h00000000} /* (5, 29, 0) {real, imag} */,
  {32'h3e397a26, 32'h00000000} /* (5, 28, 31) {real, imag} */,
  {32'hbf2557f2, 32'h00000000} /* (5, 28, 30) {real, imag} */,
  {32'hbf43a28c, 32'h00000000} /* (5, 28, 29) {real, imag} */,
  {32'hbd47073f, 32'h00000000} /* (5, 28, 28) {real, imag} */,
  {32'hbe7d7db0, 32'h00000000} /* (5, 28, 27) {real, imag} */,
  {32'hbf4b87b1, 32'h00000000} /* (5, 28, 26) {real, imag} */,
  {32'hbf2de346, 32'h00000000} /* (5, 28, 25) {real, imag} */,
  {32'hbd12fca0, 32'h00000000} /* (5, 28, 24) {real, imag} */,
  {32'hbe981499, 32'h00000000} /* (5, 28, 23) {real, imag} */,
  {32'h3d011ad6, 32'h00000000} /* (5, 28, 22) {real, imag} */,
  {32'h3f1e087d, 32'h00000000} /* (5, 28, 21) {real, imag} */,
  {32'hbdcfb612, 32'h00000000} /* (5, 28, 20) {real, imag} */,
  {32'hbe92458a, 32'h00000000} /* (5, 28, 19) {real, imag} */,
  {32'hbe665a96, 32'h00000000} /* (5, 28, 18) {real, imag} */,
  {32'h3d74122f, 32'h00000000} /* (5, 28, 17) {real, imag} */,
  {32'h3e700d88, 32'h00000000} /* (5, 28, 16) {real, imag} */,
  {32'h3e582c07, 32'h00000000} /* (5, 28, 15) {real, imag} */,
  {32'hbd1adc91, 32'h00000000} /* (5, 28, 14) {real, imag} */,
  {32'h3eaf16b0, 32'h00000000} /* (5, 28, 13) {real, imag} */,
  {32'h3f2370b5, 32'h00000000} /* (5, 28, 12) {real, imag} */,
  {32'h3f18f3ae, 32'h00000000} /* (5, 28, 11) {real, imag} */,
  {32'h3f75fbc6, 32'h00000000} /* (5, 28, 10) {real, imag} */,
  {32'hbd0cd41a, 32'h00000000} /* (5, 28, 9) {real, imag} */,
  {32'hbed0dad5, 32'h00000000} /* (5, 28, 8) {real, imag} */,
  {32'hbefa173c, 32'h00000000} /* (5, 28, 7) {real, imag} */,
  {32'hbf150239, 32'h00000000} /* (5, 28, 6) {real, imag} */,
  {32'hbea648a8, 32'h00000000} /* (5, 28, 5) {real, imag} */,
  {32'hbdbd7f82, 32'h00000000} /* (5, 28, 4) {real, imag} */,
  {32'hbe53d173, 32'h00000000} /* (5, 28, 3) {real, imag} */,
  {32'hbe58cb65, 32'h00000000} /* (5, 28, 2) {real, imag} */,
  {32'hbe4dfec1, 32'h00000000} /* (5, 28, 1) {real, imag} */,
  {32'hbe564443, 32'h00000000} /* (5, 28, 0) {real, imag} */,
  {32'hbd9eed07, 32'h00000000} /* (5, 27, 31) {real, imag} */,
  {32'hbeecfbf4, 32'h00000000} /* (5, 27, 30) {real, imag} */,
  {32'hbe3f1496, 32'h00000000} /* (5, 27, 29) {real, imag} */,
  {32'hbef72f5c, 32'h00000000} /* (5, 27, 28) {real, imag} */,
  {32'hbf2c92f6, 32'h00000000} /* (5, 27, 27) {real, imag} */,
  {32'hbe7dc60d, 32'h00000000} /* (5, 27, 26) {real, imag} */,
  {32'hbf25d024, 32'h00000000} /* (5, 27, 25) {real, imag} */,
  {32'hbf8d9e77, 32'h00000000} /* (5, 27, 24) {real, imag} */,
  {32'hbef5c17c, 32'h00000000} /* (5, 27, 23) {real, imag} */,
  {32'h3c60ca00, 32'h00000000} /* (5, 27, 22) {real, imag} */,
  {32'h3eca7aca, 32'h00000000} /* (5, 27, 21) {real, imag} */,
  {32'h3e89ac94, 32'h00000000} /* (5, 27, 20) {real, imag} */,
  {32'h3dcebbee, 32'h00000000} /* (5, 27, 19) {real, imag} */,
  {32'h3d66fcc8, 32'h00000000} /* (5, 27, 18) {real, imag} */,
  {32'h3d834d26, 32'h00000000} /* (5, 27, 17) {real, imag} */,
  {32'h3e0f9deb, 32'h00000000} /* (5, 27, 16) {real, imag} */,
  {32'h3f0c2607, 32'h00000000} /* (5, 27, 15) {real, imag} */,
  {32'h3d975b0f, 32'h00000000} /* (5, 27, 14) {real, imag} */,
  {32'h3e74ffb2, 32'h00000000} /* (5, 27, 13) {real, imag} */,
  {32'h3f12ef30, 32'h00000000} /* (5, 27, 12) {real, imag} */,
  {32'h3f56e756, 32'h00000000} /* (5, 27, 11) {real, imag} */,
  {32'h3f05e62f, 32'h00000000} /* (5, 27, 10) {real, imag} */,
  {32'h3da89fda, 32'h00000000} /* (5, 27, 9) {real, imag} */,
  {32'h3d2302ae, 32'h00000000} /* (5, 27, 8) {real, imag} */,
  {32'h3be96c37, 32'h00000000} /* (5, 27, 7) {real, imag} */,
  {32'hbdba8d02, 32'h00000000} /* (5, 27, 6) {real, imag} */,
  {32'hbe0371eb, 32'h00000000} /* (5, 27, 5) {real, imag} */,
  {32'hbe375605, 32'h00000000} /* (5, 27, 4) {real, imag} */,
  {32'hbee65b94, 32'h00000000} /* (5, 27, 3) {real, imag} */,
  {32'hbe879318, 32'h00000000} /* (5, 27, 2) {real, imag} */,
  {32'hbe65ded4, 32'h00000000} /* (5, 27, 1) {real, imag} */,
  {32'hbf159e12, 32'h00000000} /* (5, 27, 0) {real, imag} */,
  {32'hbd845cc8, 32'h00000000} /* (5, 26, 31) {real, imag} */,
  {32'hbe37c38e, 32'h00000000} /* (5, 26, 30) {real, imag} */,
  {32'hbe2bd3f2, 32'h00000000} /* (5, 26, 29) {real, imag} */,
  {32'hbe766b1f, 32'h00000000} /* (5, 26, 28) {real, imag} */,
  {32'h3d41265e, 32'h00000000} /* (5, 26, 27) {real, imag} */,
  {32'h3e69a62e, 32'h00000000} /* (5, 26, 26) {real, imag} */,
  {32'hbefa54fc, 32'h00000000} /* (5, 26, 25) {real, imag} */,
  {32'hbf8f6b53, 32'h00000000} /* (5, 26, 24) {real, imag} */,
  {32'hbf1aef38, 32'h00000000} /* (5, 26, 23) {real, imag} */,
  {32'hbe6e74f4, 32'h00000000} /* (5, 26, 22) {real, imag} */,
  {32'hbe89b5a9, 32'h00000000} /* (5, 26, 21) {real, imag} */,
  {32'h3d9b3d86, 32'h00000000} /* (5, 26, 20) {real, imag} */,
  {32'h3e36bd50, 32'h00000000} /* (5, 26, 19) {real, imag} */,
  {32'h3ebc485e, 32'h00000000} /* (5, 26, 18) {real, imag} */,
  {32'h3e04cd47, 32'h00000000} /* (5, 26, 17) {real, imag} */,
  {32'h3ddb49be, 32'h00000000} /* (5, 26, 16) {real, imag} */,
  {32'h3f57a1ad, 32'h00000000} /* (5, 26, 15) {real, imag} */,
  {32'h3f09ee1a, 32'h00000000} /* (5, 26, 14) {real, imag} */,
  {32'hbd7f96b5, 32'h00000000} /* (5, 26, 13) {real, imag} */,
  {32'h3ec2698a, 32'h00000000} /* (5, 26, 12) {real, imag} */,
  {32'h3d041c12, 32'h00000000} /* (5, 26, 11) {real, imag} */,
  {32'hbe93dea2, 32'h00000000} /* (5, 26, 10) {real, imag} */,
  {32'h3e4a2870, 32'h00000000} /* (5, 26, 9) {real, imag} */,
  {32'h3eaf14be, 32'h00000000} /* (5, 26, 8) {real, imag} */,
  {32'h3ea1f3e5, 32'h00000000} /* (5, 26, 7) {real, imag} */,
  {32'h3e7d8db5, 32'h00000000} /* (5, 26, 6) {real, imag} */,
  {32'h3d57b25e, 32'h00000000} /* (5, 26, 5) {real, imag} */,
  {32'hbd9ae6c4, 32'h00000000} /* (5, 26, 4) {real, imag} */,
  {32'hbe966c24, 32'h00000000} /* (5, 26, 3) {real, imag} */,
  {32'hbdf57931, 32'h00000000} /* (5, 26, 2) {real, imag} */,
  {32'h3e142768, 32'h00000000} /* (5, 26, 1) {real, imag} */,
  {32'hbecd9d42, 32'h00000000} /* (5, 26, 0) {real, imag} */,
  {32'hbe0f775d, 32'h00000000} /* (5, 25, 31) {real, imag} */,
  {32'hbee3bfa2, 32'h00000000} /* (5, 25, 30) {real, imag} */,
  {32'hbf020699, 32'h00000000} /* (5, 25, 29) {real, imag} */,
  {32'hbe92c6d2, 32'h00000000} /* (5, 25, 28) {real, imag} */,
  {32'hbdb902c7, 32'h00000000} /* (5, 25, 27) {real, imag} */,
  {32'hbde85a7e, 32'h00000000} /* (5, 25, 26) {real, imag} */,
  {32'hbf08d341, 32'h00000000} /* (5, 25, 25) {real, imag} */,
  {32'hbf50f931, 32'h00000000} /* (5, 25, 24) {real, imag} */,
  {32'hbf0c99f3, 32'h00000000} /* (5, 25, 23) {real, imag} */,
  {32'hbf19213d, 32'h00000000} /* (5, 25, 22) {real, imag} */,
  {32'hbf008c55, 32'h00000000} /* (5, 25, 21) {real, imag} */,
  {32'h3f0507e5, 32'h00000000} /* (5, 25, 20) {real, imag} */,
  {32'h3f03e3f3, 32'h00000000} /* (5, 25, 19) {real, imag} */,
  {32'h3e93407c, 32'h00000000} /* (5, 25, 18) {real, imag} */,
  {32'h3ed17e16, 32'h00000000} /* (5, 25, 17) {real, imag} */,
  {32'h3e9ab19c, 32'h00000000} /* (5, 25, 16) {real, imag} */,
  {32'h3f30f456, 32'h00000000} /* (5, 25, 15) {real, imag} */,
  {32'h3efd5c8d, 32'h00000000} /* (5, 25, 14) {real, imag} */,
  {32'h3c8cea23, 32'h00000000} /* (5, 25, 13) {real, imag} */,
  {32'h3e6403de, 32'h00000000} /* (5, 25, 12) {real, imag} */,
  {32'h3ec89173, 32'h00000000} /* (5, 25, 11) {real, imag} */,
  {32'h3d0a4bb5, 32'h00000000} /* (5, 25, 10) {real, imag} */,
  {32'hbd367813, 32'h00000000} /* (5, 25, 9) {real, imag} */,
  {32'hbf194f62, 32'h00000000} /* (5, 25, 8) {real, imag} */,
  {32'hbe13c113, 32'h00000000} /* (5, 25, 7) {real, imag} */,
  {32'h3e91254b, 32'h00000000} /* (5, 25, 6) {real, imag} */,
  {32'h3e916de4, 32'h00000000} /* (5, 25, 5) {real, imag} */,
  {32'hbe0ff862, 32'h00000000} /* (5, 25, 4) {real, imag} */,
  {32'hbf06f892, 32'h00000000} /* (5, 25, 3) {real, imag} */,
  {32'hbf303ac7, 32'h00000000} /* (5, 25, 2) {real, imag} */,
  {32'h3e205a7d, 32'h00000000} /* (5, 25, 1) {real, imag} */,
  {32'hbe53cd4d, 32'h00000000} /* (5, 25, 0) {real, imag} */,
  {32'h3c290701, 32'h00000000} /* (5, 24, 31) {real, imag} */,
  {32'h3e05759a, 32'h00000000} /* (5, 24, 30) {real, imag} */,
  {32'hbee121dc, 32'h00000000} /* (5, 24, 29) {real, imag} */,
  {32'hbea80617, 32'h00000000} /* (5, 24, 28) {real, imag} */,
  {32'hbf0e431e, 32'h00000000} /* (5, 24, 27) {real, imag} */,
  {32'hbeeffdc7, 32'h00000000} /* (5, 24, 26) {real, imag} */,
  {32'hbe72b64c, 32'h00000000} /* (5, 24, 25) {real, imag} */,
  {32'hbe0cd245, 32'h00000000} /* (5, 24, 24) {real, imag} */,
  {32'hbe3ee8fd, 32'h00000000} /* (5, 24, 23) {real, imag} */,
  {32'hbecc2aec, 32'h00000000} /* (5, 24, 22) {real, imag} */,
  {32'h3e0c7bec, 32'h00000000} /* (5, 24, 21) {real, imag} */,
  {32'h3f2e7641, 32'h00000000} /* (5, 24, 20) {real, imag} */,
  {32'h3f12e3b3, 32'h00000000} /* (5, 24, 19) {real, imag} */,
  {32'h3ecd4ca5, 32'h00000000} /* (5, 24, 18) {real, imag} */,
  {32'h3e54cdcf, 32'h00000000} /* (5, 24, 17) {real, imag} */,
  {32'h3e7a7c08, 32'h00000000} /* (5, 24, 16) {real, imag} */,
  {32'h3ec12ec5, 32'h00000000} /* (5, 24, 15) {real, imag} */,
  {32'hbb31b5c5, 32'h00000000} /* (5, 24, 14) {real, imag} */,
  {32'h3e63cd42, 32'h00000000} /* (5, 24, 13) {real, imag} */,
  {32'h3e09b7d7, 32'h00000000} /* (5, 24, 12) {real, imag} */,
  {32'h3f35d745, 32'h00000000} /* (5, 24, 11) {real, imag} */,
  {32'h3ee20239, 32'h00000000} /* (5, 24, 10) {real, imag} */,
  {32'hbea9e2c9, 32'h00000000} /* (5, 24, 9) {real, imag} */,
  {32'hbf05d9c8, 32'h00000000} /* (5, 24, 8) {real, imag} */,
  {32'hbe0683ef, 32'h00000000} /* (5, 24, 7) {real, imag} */,
  {32'h3da23017, 32'h00000000} /* (5, 24, 6) {real, imag} */,
  {32'h3e4e9b30, 32'h00000000} /* (5, 24, 5) {real, imag} */,
  {32'h3db7d053, 32'h00000000} /* (5, 24, 4) {real, imag} */,
  {32'hbe046fa5, 32'h00000000} /* (5, 24, 3) {real, imag} */,
  {32'hbf389420, 32'h00000000} /* (5, 24, 2) {real, imag} */,
  {32'h3db30145, 32'h00000000} /* (5, 24, 1) {real, imag} */,
  {32'hbd150b4f, 32'h00000000} /* (5, 24, 0) {real, imag} */,
  {32'hbad8b620, 32'h00000000} /* (5, 23, 31) {real, imag} */,
  {32'h3ebc3b7e, 32'h00000000} /* (5, 23, 30) {real, imag} */,
  {32'hbe42ce7d, 32'h00000000} /* (5, 23, 29) {real, imag} */,
  {32'hbeca4074, 32'h00000000} /* (5, 23, 28) {real, imag} */,
  {32'hbef79398, 32'h00000000} /* (5, 23, 27) {real, imag} */,
  {32'hbe4ec56b, 32'h00000000} /* (5, 23, 26) {real, imag} */,
  {32'h3d50a5ac, 32'h00000000} /* (5, 23, 25) {real, imag} */,
  {32'h3d1dedc9, 32'h00000000} /* (5, 23, 24) {real, imag} */,
  {32'hbe7bcd99, 32'h00000000} /* (5, 23, 23) {real, imag} */,
  {32'hbed9c475, 32'h00000000} /* (5, 23, 22) {real, imag} */,
  {32'h3e6d8e1e, 32'h00000000} /* (5, 23, 21) {real, imag} */,
  {32'h3ed17e55, 32'h00000000} /* (5, 23, 20) {real, imag} */,
  {32'h3f0b9d80, 32'h00000000} /* (5, 23, 19) {real, imag} */,
  {32'h3f51a98d, 32'h00000000} /* (5, 23, 18) {real, imag} */,
  {32'h3f1b2aa6, 32'h00000000} /* (5, 23, 17) {real, imag} */,
  {32'h3eb4112b, 32'h00000000} /* (5, 23, 16) {real, imag} */,
  {32'h3f069e26, 32'h00000000} /* (5, 23, 15) {real, imag} */,
  {32'h3e89fd36, 32'h00000000} /* (5, 23, 14) {real, imag} */,
  {32'h3e570c06, 32'h00000000} /* (5, 23, 13) {real, imag} */,
  {32'h3dcd676a, 32'h00000000} /* (5, 23, 12) {real, imag} */,
  {32'h3e898f81, 32'h00000000} /* (5, 23, 11) {real, imag} */,
  {32'hbc449fa2, 32'h00000000} /* (5, 23, 10) {real, imag} */,
  {32'hbf0c7840, 32'h00000000} /* (5, 23, 9) {real, imag} */,
  {32'hbefbf86d, 32'h00000000} /* (5, 23, 8) {real, imag} */,
  {32'hbece2885, 32'h00000000} /* (5, 23, 7) {real, imag} */,
  {32'hbee739d9, 32'h00000000} /* (5, 23, 6) {real, imag} */,
  {32'hbea6ecc0, 32'h00000000} /* (5, 23, 5) {real, imag} */,
  {32'hbd976325, 32'h00000000} /* (5, 23, 4) {real, imag} */,
  {32'hbee322f1, 32'h00000000} /* (5, 23, 3) {real, imag} */,
  {32'hbf34a714, 32'h00000000} /* (5, 23, 2) {real, imag} */,
  {32'hbea37546, 32'h00000000} /* (5, 23, 1) {real, imag} */,
  {32'hbe5ab1af, 32'h00000000} /* (5, 23, 0) {real, imag} */,
  {32'hbe4b7068, 32'h00000000} /* (5, 22, 31) {real, imag} */,
  {32'hbe735596, 32'h00000000} /* (5, 22, 30) {real, imag} */,
  {32'hbec58ed9, 32'h00000000} /* (5, 22, 29) {real, imag} */,
  {32'hbeada070, 32'h00000000} /* (5, 22, 28) {real, imag} */,
  {32'h3ca91aeb, 32'h00000000} /* (5, 22, 27) {real, imag} */,
  {32'h3d90bb1d, 32'h00000000} /* (5, 22, 26) {real, imag} */,
  {32'hbe52cba4, 32'h00000000} /* (5, 22, 25) {real, imag} */,
  {32'hbefe7e1b, 32'h00000000} /* (5, 22, 24) {real, imag} */,
  {32'hbe534ee9, 32'h00000000} /* (5, 22, 23) {real, imag} */,
  {32'hbe46777e, 32'h00000000} /* (5, 22, 22) {real, imag} */,
  {32'hbe38d75e, 32'h00000000} /* (5, 22, 21) {real, imag} */,
  {32'h3efbce13, 32'h00000000} /* (5, 22, 20) {real, imag} */,
  {32'h3f8abcfa, 32'h00000000} /* (5, 22, 19) {real, imag} */,
  {32'h3f5e6b38, 32'h00000000} /* (5, 22, 18) {real, imag} */,
  {32'h3e66a04e, 32'h00000000} /* (5, 22, 17) {real, imag} */,
  {32'h3d7613e8, 32'h00000000} /* (5, 22, 16) {real, imag} */,
  {32'h3cae1584, 32'h00000000} /* (5, 22, 15) {real, imag} */,
  {32'hbc368553, 32'h00000000} /* (5, 22, 14) {real, imag} */,
  {32'hb9801c00, 32'h00000000} /* (5, 22, 13) {real, imag} */,
  {32'hbe642e42, 32'h00000000} /* (5, 22, 12) {real, imag} */,
  {32'h3b1bf120, 32'h00000000} /* (5, 22, 11) {real, imag} */,
  {32'hbe0df001, 32'h00000000} /* (5, 22, 10) {real, imag} */,
  {32'hbe9668bc, 32'h00000000} /* (5, 22, 9) {real, imag} */,
  {32'hbec0beb3, 32'h00000000} /* (5, 22, 8) {real, imag} */,
  {32'hbe5ffb26, 32'h00000000} /* (5, 22, 7) {real, imag} */,
  {32'hbee223ae, 32'h00000000} /* (5, 22, 6) {real, imag} */,
  {32'hbe4bd0a8, 32'h00000000} /* (5, 22, 5) {real, imag} */,
  {32'hbe66f852, 32'h00000000} /* (5, 22, 4) {real, imag} */,
  {32'hbefc45c0, 32'h00000000} /* (5, 22, 3) {real, imag} */,
  {32'hbf0e57d9, 32'h00000000} /* (5, 22, 2) {real, imag} */,
  {32'hbeb96966, 32'h00000000} /* (5, 22, 1) {real, imag} */,
  {32'hbe92a3ed, 32'h00000000} /* (5, 22, 0) {real, imag} */,
  {32'hbe389290, 32'h00000000} /* (5, 21, 31) {real, imag} */,
  {32'h3d893fe0, 32'h00000000} /* (5, 21, 30) {real, imag} */,
  {32'hbd98fd68, 32'h00000000} /* (5, 21, 29) {real, imag} */,
  {32'h3e228b0f, 32'h00000000} /* (5, 21, 28) {real, imag} */,
  {32'hbc42c954, 32'h00000000} /* (5, 21, 27) {real, imag} */,
  {32'hbeee2324, 32'h00000000} /* (5, 21, 26) {real, imag} */,
  {32'hbe8713b3, 32'h00000000} /* (5, 21, 25) {real, imag} */,
  {32'h3d707990, 32'h00000000} /* (5, 21, 24) {real, imag} */,
  {32'h3defa1bb, 32'h00000000} /* (5, 21, 23) {real, imag} */,
  {32'hbc3f935a, 32'h00000000} /* (5, 21, 22) {real, imag} */,
  {32'hbe8c3176, 32'h00000000} /* (5, 21, 21) {real, imag} */,
  {32'h3eb8ef2a, 32'h00000000} /* (5, 21, 20) {real, imag} */,
  {32'h3f836062, 32'h00000000} /* (5, 21, 19) {real, imag} */,
  {32'h3eb7b195, 32'h00000000} /* (5, 21, 18) {real, imag} */,
  {32'hbed03241, 32'h00000000} /* (5, 21, 17) {real, imag} */,
  {32'hbf167253, 32'h00000000} /* (5, 21, 16) {real, imag} */,
  {32'hbd48a81a, 32'h00000000} /* (5, 21, 15) {real, imag} */,
  {32'h3eb2a3d4, 32'h00000000} /* (5, 21, 14) {real, imag} */,
  {32'hbde0d636, 32'h00000000} /* (5, 21, 13) {real, imag} */,
  {32'hbe0e8800, 32'h00000000} /* (5, 21, 12) {real, imag} */,
  {32'h3ed96608, 32'h00000000} /* (5, 21, 11) {real, imag} */,
  {32'h3f121e26, 32'h00000000} /* (5, 21, 10) {real, imag} */,
  {32'h3e2f6dc0, 32'h00000000} /* (5, 21, 9) {real, imag} */,
  {32'h3e111851, 32'h00000000} /* (5, 21, 8) {real, imag} */,
  {32'h3bae26fc, 32'h00000000} /* (5, 21, 7) {real, imag} */,
  {32'hbe1eeed5, 32'h00000000} /* (5, 21, 6) {real, imag} */,
  {32'h3e4d1ba5, 32'h00000000} /* (5, 21, 5) {real, imag} */,
  {32'hbdbfc641, 32'h00000000} /* (5, 21, 4) {real, imag} */,
  {32'hbcf34217, 32'h00000000} /* (5, 21, 3) {real, imag} */,
  {32'h3e2eb934, 32'h00000000} /* (5, 21, 2) {real, imag} */,
  {32'hbc3c243e, 32'h00000000} /* (5, 21, 1) {real, imag} */,
  {32'hbe73d45e, 32'h00000000} /* (5, 21, 0) {real, imag} */,
  {32'h3e93dea6, 32'h00000000} /* (5, 20, 31) {real, imag} */,
  {32'h3f7563e3, 32'h00000000} /* (5, 20, 30) {real, imag} */,
  {32'h3ec4a54a, 32'h00000000} /* (5, 20, 29) {real, imag} */,
  {32'h3f0dfa8e, 32'h00000000} /* (5, 20, 28) {real, imag} */,
  {32'h3e60edc2, 32'h00000000} /* (5, 20, 27) {real, imag} */,
  {32'hbf015560, 32'h00000000} /* (5, 20, 26) {real, imag} */,
  {32'hbdb0e832, 32'h00000000} /* (5, 20, 25) {real, imag} */,
  {32'h3efd2d97, 32'h00000000} /* (5, 20, 24) {real, imag} */,
  {32'h3edbd1ab, 32'h00000000} /* (5, 20, 23) {real, imag} */,
  {32'h3e9cd03c, 32'h00000000} /* (5, 20, 22) {real, imag} */,
  {32'h3e9eee7a, 32'h00000000} /* (5, 20, 21) {real, imag} */,
  {32'h3e482b07, 32'h00000000} /* (5, 20, 20) {real, imag} */,
  {32'h3e850905, 32'h00000000} /* (5, 20, 19) {real, imag} */,
  {32'h3dbcea54, 32'h00000000} /* (5, 20, 18) {real, imag} */,
  {32'hbeeaa2ba, 32'h00000000} /* (5, 20, 17) {real, imag} */,
  {32'hbf1047f3, 32'h00000000} /* (5, 20, 16) {real, imag} */,
  {32'h3dae7bbe, 32'h00000000} /* (5, 20, 15) {real, imag} */,
  {32'h3d3d4d72, 32'h00000000} /* (5, 20, 14) {real, imag} */,
  {32'hbeb3a985, 32'h00000000} /* (5, 20, 13) {real, imag} */,
  {32'hbda4c1a5, 32'h00000000} /* (5, 20, 12) {real, imag} */,
  {32'h3ece4341, 32'h00000000} /* (5, 20, 11) {real, imag} */,
  {32'h3f819876, 32'h00000000} /* (5, 20, 10) {real, imag} */,
  {32'h3ef51835, 32'h00000000} /* (5, 20, 9) {real, imag} */,
  {32'hbdaf8ee3, 32'h00000000} /* (5, 20, 8) {real, imag} */,
  {32'h3e130e8c, 32'h00000000} /* (5, 20, 7) {real, imag} */,
  {32'h3f09796b, 32'h00000000} /* (5, 20, 6) {real, imag} */,
  {32'h3f700fcc, 32'h00000000} /* (5, 20, 5) {real, imag} */,
  {32'h3de860bf, 32'h00000000} /* (5, 20, 4) {real, imag} */,
  {32'hbcd2f665, 32'h00000000} /* (5, 20, 3) {real, imag} */,
  {32'h3f0b00d9, 32'h00000000} /* (5, 20, 2) {real, imag} */,
  {32'h3f031290, 32'h00000000} /* (5, 20, 1) {real, imag} */,
  {32'hbd1bbc89, 32'h00000000} /* (5, 20, 0) {real, imag} */,
  {32'h3e672d13, 32'h00000000} /* (5, 19, 31) {real, imag} */,
  {32'h3f2960f4, 32'h00000000} /* (5, 19, 30) {real, imag} */,
  {32'h3db55fd9, 32'h00000000} /* (5, 19, 29) {real, imag} */,
  {32'h3f0a9f34, 32'h00000000} /* (5, 19, 28) {real, imag} */,
  {32'h3e3ef689, 32'h00000000} /* (5, 19, 27) {real, imag} */,
  {32'hbe46fee9, 32'h00000000} /* (5, 19, 26) {real, imag} */,
  {32'hbeceeb58, 32'h00000000} /* (5, 19, 25) {real, imag} */,
  {32'hbe1b8917, 32'h00000000} /* (5, 19, 24) {real, imag} */,
  {32'h3de00f1b, 32'h00000000} /* (5, 19, 23) {real, imag} */,
  {32'h3e80ae0b, 32'h00000000} /* (5, 19, 22) {real, imag} */,
  {32'h3cd59519, 32'h00000000} /* (5, 19, 21) {real, imag} */,
  {32'hbe35b810, 32'h00000000} /* (5, 19, 20) {real, imag} */,
  {32'hbdf3b9ef, 32'h00000000} /* (5, 19, 19) {real, imag} */,
  {32'hbc8035a4, 32'h00000000} /* (5, 19, 18) {real, imag} */,
  {32'hbed9dd7d, 32'h00000000} /* (5, 19, 17) {real, imag} */,
  {32'hbf32c231, 32'h00000000} /* (5, 19, 16) {real, imag} */,
  {32'hbee637e9, 32'h00000000} /* (5, 19, 15) {real, imag} */,
  {32'hbeb71886, 32'h00000000} /* (5, 19, 14) {real, imag} */,
  {32'hbe29fd37, 32'h00000000} /* (5, 19, 13) {real, imag} */,
  {32'h3c4df3d0, 32'h00000000} /* (5, 19, 12) {real, imag} */,
  {32'hbce6c397, 32'h00000000} /* (5, 19, 11) {real, imag} */,
  {32'h3f08c60a, 32'h00000000} /* (5, 19, 10) {real, imag} */,
  {32'h3f295163, 32'h00000000} /* (5, 19, 9) {real, imag} */,
  {32'hbde8c350, 32'h00000000} /* (5, 19, 8) {real, imag} */,
  {32'h3e639ae8, 32'h00000000} /* (5, 19, 7) {real, imag} */,
  {32'h3ef613ff, 32'h00000000} /* (5, 19, 6) {real, imag} */,
  {32'h3f232938, 32'h00000000} /* (5, 19, 5) {real, imag} */,
  {32'h3e926ff5, 32'h00000000} /* (5, 19, 4) {real, imag} */,
  {32'hbe2000ca, 32'h00000000} /* (5, 19, 3) {real, imag} */,
  {32'hbd6201f0, 32'h00000000} /* (5, 19, 2) {real, imag} */,
  {32'h3e659334, 32'h00000000} /* (5, 19, 1) {real, imag} */,
  {32'hbea9445a, 32'h00000000} /* (5, 19, 0) {real, imag} */,
  {32'h3ded7723, 32'h00000000} /* (5, 18, 31) {real, imag} */,
  {32'h3e196006, 32'h00000000} /* (5, 18, 30) {real, imag} */,
  {32'h3e5dc94f, 32'h00000000} /* (5, 18, 29) {real, imag} */,
  {32'h3eb75b58, 32'h00000000} /* (5, 18, 28) {real, imag} */,
  {32'hbe489ce3, 32'h00000000} /* (5, 18, 27) {real, imag} */,
  {32'h3d8b3a2a, 32'h00000000} /* (5, 18, 26) {real, imag} */,
  {32'hbd97a0e1, 32'h00000000} /* (5, 18, 25) {real, imag} */,
  {32'hbeca6999, 32'h00000000} /* (5, 18, 24) {real, imag} */,
  {32'hbdb3bc75, 32'h00000000} /* (5, 18, 23) {real, imag} */,
  {32'h3e745dc2, 32'h00000000} /* (5, 18, 22) {real, imag} */,
  {32'h3e636210, 32'h00000000} /* (5, 18, 21) {real, imag} */,
  {32'h3ea63205, 32'h00000000} /* (5, 18, 20) {real, imag} */,
  {32'h3d9240bd, 32'h00000000} /* (5, 18, 19) {real, imag} */,
  {32'h3d9a0476, 32'h00000000} /* (5, 18, 18) {real, imag} */,
  {32'hbe7a7337, 32'h00000000} /* (5, 18, 17) {real, imag} */,
  {32'hbf3c685d, 32'h00000000} /* (5, 18, 16) {real, imag} */,
  {32'hbed48ccc, 32'h00000000} /* (5, 18, 15) {real, imag} */,
  {32'hbee0c026, 32'h00000000} /* (5, 18, 14) {real, imag} */,
  {32'hbe0d3d23, 32'h00000000} /* (5, 18, 13) {real, imag} */,
  {32'hbb015db4, 32'h00000000} /* (5, 18, 12) {real, imag} */,
  {32'hbe506923, 32'h00000000} /* (5, 18, 11) {real, imag} */,
  {32'h3c8c16b6, 32'h00000000} /* (5, 18, 10) {real, imag} */,
  {32'h3e1a13ca, 32'h00000000} /* (5, 18, 9) {real, imag} */,
  {32'h3d81634d, 32'h00000000} /* (5, 18, 8) {real, imag} */,
  {32'h3ea9d1ca, 32'h00000000} /* (5, 18, 7) {real, imag} */,
  {32'h3f3086e2, 32'h00000000} /* (5, 18, 6) {real, imag} */,
  {32'h3f616b7d, 32'h00000000} /* (5, 18, 5) {real, imag} */,
  {32'h3f05063b, 32'h00000000} /* (5, 18, 4) {real, imag} */,
  {32'h3dff0811, 32'h00000000} /* (5, 18, 3) {real, imag} */,
  {32'hbdd46b15, 32'h00000000} /* (5, 18, 2) {real, imag} */,
  {32'h3f17ffc1, 32'h00000000} /* (5, 18, 1) {real, imag} */,
  {32'hbdb5ddbd, 32'h00000000} /* (5, 18, 0) {real, imag} */,
  {32'h3d8c13ce, 32'h00000000} /* (5, 17, 31) {real, imag} */,
  {32'h3cd29143, 32'h00000000} /* (5, 17, 30) {real, imag} */,
  {32'hbe6c7950, 32'h00000000} /* (5, 17, 29) {real, imag} */,
  {32'hbe61e313, 32'h00000000} /* (5, 17, 28) {real, imag} */,
  {32'hbde79d19, 32'h00000000} /* (5, 17, 27) {real, imag} */,
  {32'h3e86eec2, 32'h00000000} /* (5, 17, 26) {real, imag} */,
  {32'h3ed3fc85, 32'h00000000} /* (5, 17, 25) {real, imag} */,
  {32'h3de158e4, 32'h00000000} /* (5, 17, 24) {real, imag} */,
  {32'h3ea7a9a2, 32'h00000000} /* (5, 17, 23) {real, imag} */,
  {32'h3e974d17, 32'h00000000} /* (5, 17, 22) {real, imag} */,
  {32'h3e9173fb, 32'h00000000} /* (5, 17, 21) {real, imag} */,
  {32'h3ef965e8, 32'h00000000} /* (5, 17, 20) {real, imag} */,
  {32'h3c2bea9e, 32'h00000000} /* (5, 17, 19) {real, imag} */,
  {32'hbe5b1337, 32'h00000000} /* (5, 17, 18) {real, imag} */,
  {32'hbe54076f, 32'h00000000} /* (5, 17, 17) {real, imag} */,
  {32'hbe249448, 32'h00000000} /* (5, 17, 16) {real, imag} */,
  {32'hbdc0bad8, 32'h00000000} /* (5, 17, 15) {real, imag} */,
  {32'h3da650b1, 32'h00000000} /* (5, 17, 14) {real, imag} */,
  {32'h3ce5361a, 32'h00000000} /* (5, 17, 13) {real, imag} */,
  {32'hbd11e2f6, 32'h00000000} /* (5, 17, 12) {real, imag} */,
  {32'hbe3d8815, 32'h00000000} /* (5, 17, 11) {real, imag} */,
  {32'h3e847cae, 32'h00000000} /* (5, 17, 10) {real, imag} */,
  {32'h3e04081c, 32'h00000000} /* (5, 17, 9) {real, imag} */,
  {32'h3efec785, 32'h00000000} /* (5, 17, 8) {real, imag} */,
  {32'h3e317d8d, 32'h00000000} /* (5, 17, 7) {real, imag} */,
  {32'h3e535f7f, 32'h00000000} /* (5, 17, 6) {real, imag} */,
  {32'h3f03cb82, 32'h00000000} /* (5, 17, 5) {real, imag} */,
  {32'h3eeb51b1, 32'h00000000} /* (5, 17, 4) {real, imag} */,
  {32'h3f092f9f, 32'h00000000} /* (5, 17, 3) {real, imag} */,
  {32'h3f30d6be, 32'h00000000} /* (5, 17, 2) {real, imag} */,
  {32'h3f5a8274, 32'h00000000} /* (5, 17, 1) {real, imag} */,
  {32'h3e792e29, 32'h00000000} /* (5, 17, 0) {real, imag} */,
  {32'h3e54f3b9, 32'h00000000} /* (5, 16, 31) {real, imag} */,
  {32'hbe02cd8d, 32'h00000000} /* (5, 16, 30) {real, imag} */,
  {32'hbe8102ad, 32'h00000000} /* (5, 16, 29) {real, imag} */,
  {32'h3de499a5, 32'h00000000} /* (5, 16, 28) {real, imag} */,
  {32'h3e1fabba, 32'h00000000} /* (5, 16, 27) {real, imag} */,
  {32'h3eca62bf, 32'h00000000} /* (5, 16, 26) {real, imag} */,
  {32'h3f185b2a, 32'h00000000} /* (5, 16, 25) {real, imag} */,
  {32'h3ee7ca34, 32'h00000000} /* (5, 16, 24) {real, imag} */,
  {32'h3f6a0477, 32'h00000000} /* (5, 16, 23) {real, imag} */,
  {32'h3ef91a8e, 32'h00000000} /* (5, 16, 22) {real, imag} */,
  {32'h3ec190e3, 32'h00000000} /* (5, 16, 21) {real, imag} */,
  {32'h3f0599a9, 32'h00000000} /* (5, 16, 20) {real, imag} */,
  {32'h3e59db6f, 32'h00000000} /* (5, 16, 19) {real, imag} */,
  {32'hbb21ca76, 32'h00000000} /* (5, 16, 18) {real, imag} */,
  {32'hbe22e8a0, 32'h00000000} /* (5, 16, 17) {real, imag} */,
  {32'hbf3eb50d, 32'h00000000} /* (5, 16, 16) {real, imag} */,
  {32'hbefa50a3, 32'h00000000} /* (5, 16, 15) {real, imag} */,
  {32'h3ed262e8, 32'h00000000} /* (5, 16, 14) {real, imag} */,
  {32'h3e7271c2, 32'h00000000} /* (5, 16, 13) {real, imag} */,
  {32'hbec11a61, 32'h00000000} /* (5, 16, 12) {real, imag} */,
  {32'hbe872177, 32'h00000000} /* (5, 16, 11) {real, imag} */,
  {32'h3e8ce430, 32'h00000000} /* (5, 16, 10) {real, imag} */,
  {32'h3e939b29, 32'h00000000} /* (5, 16, 9) {real, imag} */,
  {32'h3f0dd68a, 32'h00000000} /* (5, 16, 8) {real, imag} */,
  {32'h3eb1eec1, 32'h00000000} /* (5, 16, 7) {real, imag} */,
  {32'h3ecf1216, 32'h00000000} /* (5, 16, 6) {real, imag} */,
  {32'h3f068d9c, 32'h00000000} /* (5, 16, 5) {real, imag} */,
  {32'h3ea403eb, 32'h00000000} /* (5, 16, 4) {real, imag} */,
  {32'hbdc44d30, 32'h00000000} /* (5, 16, 3) {real, imag} */,
  {32'h3d99e81c, 32'h00000000} /* (5, 16, 2) {real, imag} */,
  {32'h3ea2f773, 32'h00000000} /* (5, 16, 1) {real, imag} */,
  {32'h3eb3f21c, 32'h00000000} /* (5, 16, 0) {real, imag} */,
  {32'h3ea115ab, 32'h00000000} /* (5, 15, 31) {real, imag} */,
  {32'h3e0e38b8, 32'h00000000} /* (5, 15, 30) {real, imag} */,
  {32'h3e721eaf, 32'h00000000} /* (5, 15, 29) {real, imag} */,
  {32'h3e685c23, 32'h00000000} /* (5, 15, 28) {real, imag} */,
  {32'h3e7bdbf4, 32'h00000000} /* (5, 15, 27) {real, imag} */,
  {32'h3eb55f51, 32'h00000000} /* (5, 15, 26) {real, imag} */,
  {32'hbd973690, 32'h00000000} /* (5, 15, 25) {real, imag} */,
  {32'h3e4b58db, 32'h00000000} /* (5, 15, 24) {real, imag} */,
  {32'h3f2c89a0, 32'h00000000} /* (5, 15, 23) {real, imag} */,
  {32'h3eb71b24, 32'h00000000} /* (5, 15, 22) {real, imag} */,
  {32'h3e4bd28e, 32'h00000000} /* (5, 15, 21) {real, imag} */,
  {32'h3efb14e0, 32'h00000000} /* (5, 15, 20) {real, imag} */,
  {32'h3edf2e79, 32'h00000000} /* (5, 15, 19) {real, imag} */,
  {32'h3dd171cc, 32'h00000000} /* (5, 15, 18) {real, imag} */,
  {32'hbdead0c5, 32'h00000000} /* (5, 15, 17) {real, imag} */,
  {32'hbd2ccde0, 32'h00000000} /* (5, 15, 16) {real, imag} */,
  {32'hbf3535e6, 32'h00000000} /* (5, 15, 15) {real, imag} */,
  {32'hbebecb08, 32'h00000000} /* (5, 15, 14) {real, imag} */,
  {32'hbf8e8d10, 32'h00000000} /* (5, 15, 13) {real, imag} */,
  {32'hbf7a533d, 32'h00000000} /* (5, 15, 12) {real, imag} */,
  {32'hbe7f155a, 32'h00000000} /* (5, 15, 11) {real, imag} */,
  {32'h3cae216f, 32'h00000000} /* (5, 15, 10) {real, imag} */,
  {32'h3f14f356, 32'h00000000} /* (5, 15, 9) {real, imag} */,
  {32'h3e5d8616, 32'h00000000} /* (5, 15, 8) {real, imag} */,
  {32'hbc597014, 32'h00000000} /* (5, 15, 7) {real, imag} */,
  {32'h3e7961a9, 32'h00000000} /* (5, 15, 6) {real, imag} */,
  {32'h3e708eef, 32'h00000000} /* (5, 15, 5) {real, imag} */,
  {32'h3cf522ae, 32'h00000000} /* (5, 15, 4) {real, imag} */,
  {32'hbef37827, 32'h00000000} /* (5, 15, 3) {real, imag} */,
  {32'hbf021d42, 32'h00000000} /* (5, 15, 2) {real, imag} */,
  {32'h3e809b57, 32'h00000000} /* (5, 15, 1) {real, imag} */,
  {32'h3e3002ff, 32'h00000000} /* (5, 15, 0) {real, imag} */,
  {32'h3e351aba, 32'h00000000} /* (5, 14, 31) {real, imag} */,
  {32'h3ddc9dc8, 32'h00000000} /* (5, 14, 30) {real, imag} */,
  {32'h3e8628d3, 32'h00000000} /* (5, 14, 29) {real, imag} */,
  {32'h3e89fbd5, 32'h00000000} /* (5, 14, 28) {real, imag} */,
  {32'h3eb7990a, 32'h00000000} /* (5, 14, 27) {real, imag} */,
  {32'h3d97e860, 32'h00000000} /* (5, 14, 26) {real, imag} */,
  {32'hbf0f1319, 32'h00000000} /* (5, 14, 25) {real, imag} */,
  {32'hbf047b9f, 32'h00000000} /* (5, 14, 24) {real, imag} */,
  {32'hbe0571fe, 32'h00000000} /* (5, 14, 23) {real, imag} */,
  {32'h3e34b172, 32'h00000000} /* (5, 14, 22) {real, imag} */,
  {32'h3d247c50, 32'h00000000} /* (5, 14, 21) {real, imag} */,
  {32'hbef320d0, 32'h00000000} /* (5, 14, 20) {real, imag} */,
  {32'hbe9b5136, 32'h00000000} /* (5, 14, 19) {real, imag} */,
  {32'hbe481f3e, 32'h00000000} /* (5, 14, 18) {real, imag} */,
  {32'hbf5ccaad, 32'h00000000} /* (5, 14, 17) {real, imag} */,
  {32'hbe603e01, 32'h00000000} /* (5, 14, 16) {real, imag} */,
  {32'hbec13039, 32'h00000000} /* (5, 14, 15) {real, imag} */,
  {32'hbe6bc8e1, 32'h00000000} /* (5, 14, 14) {real, imag} */,
  {32'hbf2acda0, 32'h00000000} /* (5, 14, 13) {real, imag} */,
  {32'hbe61969c, 32'h00000000} /* (5, 14, 12) {real, imag} */,
  {32'hbd787036, 32'h00000000} /* (5, 14, 11) {real, imag} */,
  {32'hbe8ff31e, 32'h00000000} /* (5, 14, 10) {real, imag} */,
  {32'h3ecc95c9, 32'h00000000} /* (5, 14, 9) {real, imag} */,
  {32'h3f079d11, 32'h00000000} /* (5, 14, 8) {real, imag} */,
  {32'h3df03499, 32'h00000000} /* (5, 14, 7) {real, imag} */,
  {32'h3d4d6f9f, 32'h00000000} /* (5, 14, 6) {real, imag} */,
  {32'hbddec66b, 32'h00000000} /* (5, 14, 5) {real, imag} */,
  {32'hbe24bf18, 32'h00000000} /* (5, 14, 4) {real, imag} */,
  {32'hbec58b66, 32'h00000000} /* (5, 14, 3) {real, imag} */,
  {32'hbf2b989d, 32'h00000000} /* (5, 14, 2) {real, imag} */,
  {32'hbdb6af9f, 32'h00000000} /* (5, 14, 1) {real, imag} */,
  {32'h3e154c9e, 32'h00000000} /* (5, 14, 0) {real, imag} */,
  {32'hbc2a6358, 32'h00000000} /* (5, 13, 31) {real, imag} */,
  {32'hbe4f42a4, 32'h00000000} /* (5, 13, 30) {real, imag} */,
  {32'h3eed8ba0, 32'h00000000} /* (5, 13, 29) {real, imag} */,
  {32'h3f69e84c, 32'h00000000} /* (5, 13, 28) {real, imag} */,
  {32'h3f57cc70, 32'h00000000} /* (5, 13, 27) {real, imag} */,
  {32'h3f00ea27, 32'h00000000} /* (5, 13, 26) {real, imag} */,
  {32'hbea69e69, 32'h00000000} /* (5, 13, 25) {real, imag} */,
  {32'hbf443aa5, 32'h00000000} /* (5, 13, 24) {real, imag} */,
  {32'hbe61388c, 32'h00000000} /* (5, 13, 23) {real, imag} */,
  {32'h3f47813e, 32'h00000000} /* (5, 13, 22) {real, imag} */,
  {32'h3f097717, 32'h00000000} /* (5, 13, 21) {real, imag} */,
  {32'hbf880329, 32'h00000000} /* (5, 13, 20) {real, imag} */,
  {32'hbf7bfe5f, 32'h00000000} /* (5, 13, 19) {real, imag} */,
  {32'hbf5f0a5c, 32'h00000000} /* (5, 13, 18) {real, imag} */,
  {32'hbf771992, 32'h00000000} /* (5, 13, 17) {real, imag} */,
  {32'hbee4a493, 32'h00000000} /* (5, 13, 16) {real, imag} */,
  {32'hbe3a552a, 32'h00000000} /* (5, 13, 15) {real, imag} */,
  {32'hbec46ed3, 32'h00000000} /* (5, 13, 14) {real, imag} */,
  {32'hbeb12b84, 32'h00000000} /* (5, 13, 13) {real, imag} */,
  {32'hbd28ed50, 32'h00000000} /* (5, 13, 12) {real, imag} */,
  {32'hbd061a5e, 32'h00000000} /* (5, 13, 11) {real, imag} */,
  {32'hbe4a540e, 32'h00000000} /* (5, 13, 10) {real, imag} */,
  {32'hbe54f6da, 32'h00000000} /* (5, 13, 9) {real, imag} */,
  {32'h3e0bf257, 32'h00000000} /* (5, 13, 8) {real, imag} */,
  {32'hbddc18ab, 32'h00000000} /* (5, 13, 7) {real, imag} */,
  {32'hbcd30b54, 32'h00000000} /* (5, 13, 6) {real, imag} */,
  {32'hbd2cce76, 32'h00000000} /* (5, 13, 5) {real, imag} */,
  {32'hbea236aa, 32'h00000000} /* (5, 13, 4) {real, imag} */,
  {32'hbf09a4d2, 32'h00000000} /* (5, 13, 3) {real, imag} */,
  {32'hbc2899cd, 32'h00000000} /* (5, 13, 2) {real, imag} */,
  {32'h3e3e5eeb, 32'h00000000} /* (5, 13, 1) {real, imag} */,
  {32'h3e3ec059, 32'h00000000} /* (5, 13, 0) {real, imag} */,
  {32'hbdadf5b2, 32'h00000000} /* (5, 12, 31) {real, imag} */,
  {32'hbe002e02, 32'h00000000} /* (5, 12, 30) {real, imag} */,
  {32'h3efc0428, 32'h00000000} /* (5, 12, 29) {real, imag} */,
  {32'h3f55abc0, 32'h00000000} /* (5, 12, 28) {real, imag} */,
  {32'h3edd501e, 32'h00000000} /* (5, 12, 27) {real, imag} */,
  {32'hbe206c30, 32'h00000000} /* (5, 12, 26) {real, imag} */,
  {32'hbd79bd5d, 32'h00000000} /* (5, 12, 25) {real, imag} */,
  {32'hbf00c9df, 32'h00000000} /* (5, 12, 24) {real, imag} */,
  {32'hbe815230, 32'h00000000} /* (5, 12, 23) {real, imag} */,
  {32'h3edacd8b, 32'h00000000} /* (5, 12, 22) {real, imag} */,
  {32'h3ed061d3, 32'h00000000} /* (5, 12, 21) {real, imag} */,
  {32'hbf09f386, 32'h00000000} /* (5, 12, 20) {real, imag} */,
  {32'hbf8eea11, 32'h00000000} /* (5, 12, 19) {real, imag} */,
  {32'hbf0ce64c, 32'h00000000} /* (5, 12, 18) {real, imag} */,
  {32'hbe855883, 32'h00000000} /* (5, 12, 17) {real, imag} */,
  {32'hbd66a98c, 32'h00000000} /* (5, 12, 16) {real, imag} */,
  {32'hbce9ef11, 32'h00000000} /* (5, 12, 15) {real, imag} */,
  {32'hbedd2491, 32'h00000000} /* (5, 12, 14) {real, imag} */,
  {32'hbda04241, 32'h00000000} /* (5, 12, 13) {real, imag} */,
  {32'h3ee46814, 32'h00000000} /* (5, 12, 12) {real, imag} */,
  {32'h3e5f7737, 32'h00000000} /* (5, 12, 11) {real, imag} */,
  {32'h3e8526ad, 32'h00000000} /* (5, 12, 10) {real, imag} */,
  {32'hbe0745a2, 32'h00000000} /* (5, 12, 9) {real, imag} */,
  {32'hbdc53062, 32'h00000000} /* (5, 12, 8) {real, imag} */,
  {32'h3bda03ce, 32'h00000000} /* (5, 12, 7) {real, imag} */,
  {32'hbdc4781a, 32'h00000000} /* (5, 12, 6) {real, imag} */,
  {32'h3dbbe1f7, 32'h00000000} /* (5, 12, 5) {real, imag} */,
  {32'h3e62fdfd, 32'h00000000} /* (5, 12, 4) {real, imag} */,
  {32'h3e776214, 32'h00000000} /* (5, 12, 3) {real, imag} */,
  {32'h3f2385db, 32'h00000000} /* (5, 12, 2) {real, imag} */,
  {32'h3f386569, 32'h00000000} /* (5, 12, 1) {real, imag} */,
  {32'h3e83247d, 32'h00000000} /* (5, 12, 0) {real, imag} */,
  {32'h3e2fbafc, 32'h00000000} /* (5, 11, 31) {real, imag} */,
  {32'h3ec6aef3, 32'h00000000} /* (5, 11, 30) {real, imag} */,
  {32'h3d0b3ad7, 32'h00000000} /* (5, 11, 29) {real, imag} */,
  {32'h3ed83778, 32'h00000000} /* (5, 11, 28) {real, imag} */,
  {32'h3e83bd83, 32'h00000000} /* (5, 11, 27) {real, imag} */,
  {32'h3d1a93ee, 32'h00000000} /* (5, 11, 26) {real, imag} */,
  {32'h3e991bcc, 32'h00000000} /* (5, 11, 25) {real, imag} */,
  {32'hbe0a3ba9, 32'h00000000} /* (5, 11, 24) {real, imag} */,
  {32'h3de6f08a, 32'h00000000} /* (5, 11, 23) {real, imag} */,
  {32'h3f3d98b0, 32'h00000000} /* (5, 11, 22) {real, imag} */,
  {32'h3e7280c4, 32'h00000000} /* (5, 11, 21) {real, imag} */,
  {32'h3de0a819, 32'h00000000} /* (5, 11, 20) {real, imag} */,
  {32'hbf078bcd, 32'h00000000} /* (5, 11, 19) {real, imag} */,
  {32'hbea8dc13, 32'h00000000} /* (5, 11, 18) {real, imag} */,
  {32'hbe9a1fff, 32'h00000000} /* (5, 11, 17) {real, imag} */,
  {32'h3dc99822, 32'h00000000} /* (5, 11, 16) {real, imag} */,
  {32'h3d97c857, 32'h00000000} /* (5, 11, 15) {real, imag} */,
  {32'hbd65a9fd, 32'h00000000} /* (5, 11, 14) {real, imag} */,
  {32'hbf039c56, 32'h00000000} /* (5, 11, 13) {real, imag} */,
  {32'hbe1a6d3f, 32'h00000000} /* (5, 11, 12) {real, imag} */,
  {32'h3de12d58, 32'h00000000} /* (5, 11, 11) {real, imag} */,
  {32'h3e916499, 32'h00000000} /* (5, 11, 10) {real, imag} */,
  {32'hbe44659d, 32'h00000000} /* (5, 11, 9) {real, imag} */,
  {32'hbe15e494, 32'h00000000} /* (5, 11, 8) {real, imag} */,
  {32'h3e19aefa, 32'h00000000} /* (5, 11, 7) {real, imag} */,
  {32'hbebfbc1b, 32'h00000000} /* (5, 11, 6) {real, imag} */,
  {32'hbe3b8ab6, 32'h00000000} /* (5, 11, 5) {real, imag} */,
  {32'h3d9b360c, 32'h00000000} /* (5, 11, 4) {real, imag} */,
  {32'hbd90126e, 32'h00000000} /* (5, 11, 3) {real, imag} */,
  {32'hbd66fd29, 32'h00000000} /* (5, 11, 2) {real, imag} */,
  {32'h3f8002bb, 32'h00000000} /* (5, 11, 1) {real, imag} */,
  {32'h3f21d0b6, 32'h00000000} /* (5, 11, 0) {real, imag} */,
  {32'h3d985049, 32'h00000000} /* (5, 10, 31) {real, imag} */,
  {32'h3ecb14e8, 32'h00000000} /* (5, 10, 30) {real, imag} */,
  {32'h3d849f21, 32'h00000000} /* (5, 10, 29) {real, imag} */,
  {32'hbd0934f5, 32'h00000000} /* (5, 10, 28) {real, imag} */,
  {32'h3d971732, 32'h00000000} /* (5, 10, 27) {real, imag} */,
  {32'h3e2f1421, 32'h00000000} /* (5, 10, 26) {real, imag} */,
  {32'hbdfad87d, 32'h00000000} /* (5, 10, 25) {real, imag} */,
  {32'hbe78d9a9, 32'h00000000} /* (5, 10, 24) {real, imag} */,
  {32'h3eb5cef4, 32'h00000000} /* (5, 10, 23) {real, imag} */,
  {32'h3e992b25, 32'h00000000} /* (5, 10, 22) {real, imag} */,
  {32'hbf3ea6fc, 32'h00000000} /* (5, 10, 21) {real, imag} */,
  {32'h3ca36f52, 32'h00000000} /* (5, 10, 20) {real, imag} */,
  {32'h3f01758b, 32'h00000000} /* (5, 10, 19) {real, imag} */,
  {32'hbe8b3abb, 32'h00000000} /* (5, 10, 18) {real, imag} */,
  {32'hbe8a7922, 32'h00000000} /* (5, 10, 17) {real, imag} */,
  {32'h3ee84269, 32'h00000000} /* (5, 10, 16) {real, imag} */,
  {32'h3f1f5ba3, 32'h00000000} /* (5, 10, 15) {real, imag} */,
  {32'h3e45b507, 32'h00000000} /* (5, 10, 14) {real, imag} */,
  {32'hbe68a81e, 32'h00000000} /* (5, 10, 13) {real, imag} */,
  {32'hbdfe4b5a, 32'h00000000} /* (5, 10, 12) {real, imag} */,
  {32'h3e900c99, 32'h00000000} /* (5, 10, 11) {real, imag} */,
  {32'hbebc1a49, 32'h00000000} /* (5, 10, 10) {real, imag} */,
  {32'hbf0dc4f4, 32'h00000000} /* (5, 10, 9) {real, imag} */,
  {32'hbcb96ecb, 32'h00000000} /* (5, 10, 8) {real, imag} */,
  {32'h3d82ac7b, 32'h00000000} /* (5, 10, 7) {real, imag} */,
  {32'hbf1dc78d, 32'h00000000} /* (5, 10, 6) {real, imag} */,
  {32'hbe7a23c7, 32'h00000000} /* (5, 10, 5) {real, imag} */,
  {32'hbe3ecd66, 32'h00000000} /* (5, 10, 4) {real, imag} */,
  {32'hbe19235a, 32'h00000000} /* (5, 10, 3) {real, imag} */,
  {32'hbf1d8ce5, 32'h00000000} /* (5, 10, 2) {real, imag} */,
  {32'h3d983e19, 32'h00000000} /* (5, 10, 1) {real, imag} */,
  {32'h3df7ccd4, 32'h00000000} /* (5, 10, 0) {real, imag} */,
  {32'hbe08ccd6, 32'h00000000} /* (5, 9, 31) {real, imag} */,
  {32'hbe8321a3, 32'h00000000} /* (5, 9, 30) {real, imag} */,
  {32'hbe6de67d, 32'h00000000} /* (5, 9, 29) {real, imag} */,
  {32'hbe615929, 32'h00000000} /* (5, 9, 28) {real, imag} */,
  {32'hbbb25cec, 32'h00000000} /* (5, 9, 27) {real, imag} */,
  {32'h3e0eea67, 32'h00000000} /* (5, 9, 26) {real, imag} */,
  {32'hbe28ae87, 32'h00000000} /* (5, 9, 25) {real, imag} */,
  {32'hbed2e821, 32'h00000000} /* (5, 9, 24) {real, imag} */,
  {32'h3e97ff39, 32'h00000000} /* (5, 9, 23) {real, imag} */,
  {32'h3dc17347, 32'h00000000} /* (5, 9, 22) {real, imag} */,
  {32'hbeaf506d, 32'h00000000} /* (5, 9, 21) {real, imag} */,
  {32'h3ab31434, 32'h00000000} /* (5, 9, 20) {real, imag} */,
  {32'h3e6a212f, 32'h00000000} /* (5, 9, 19) {real, imag} */,
  {32'h3e787b06, 32'h00000000} /* (5, 9, 18) {real, imag} */,
  {32'h3e58540c, 32'h00000000} /* (5, 9, 17) {real, imag} */,
  {32'h3f49a929, 32'h00000000} /* (5, 9, 16) {real, imag} */,
  {32'h3f7a619a, 32'h00000000} /* (5, 9, 15) {real, imag} */,
  {32'hba8192dc, 32'h00000000} /* (5, 9, 14) {real, imag} */,
  {32'h3d13d765, 32'h00000000} /* (5, 9, 13) {real, imag} */,
  {32'h3ec6fd67, 32'h00000000} /* (5, 9, 12) {real, imag} */,
  {32'h3f27b012, 32'h00000000} /* (5, 9, 11) {real, imag} */,
  {32'hbccac09c, 32'h00000000} /* (5, 9, 10) {real, imag} */,
  {32'hbe9613fb, 32'h00000000} /* (5, 9, 9) {real, imag} */,
  {32'hbea89f9a, 32'h00000000} /* (5, 9, 8) {real, imag} */,
  {32'h3e3ccae6, 32'h00000000} /* (5, 9, 7) {real, imag} */,
  {32'hbe2cf759, 32'h00000000} /* (5, 9, 6) {real, imag} */,
  {32'hbe9b8270, 32'h00000000} /* (5, 9, 5) {real, imag} */,
  {32'hbe03022f, 32'h00000000} /* (5, 9, 4) {real, imag} */,
  {32'hbdcce089, 32'h00000000} /* (5, 9, 3) {real, imag} */,
  {32'hbf02cbdd, 32'h00000000} /* (5, 9, 2) {real, imag} */,
  {32'hbdf2df84, 32'h00000000} /* (5, 9, 1) {real, imag} */,
  {32'hbd5a2f01, 32'h00000000} /* (5, 9, 0) {real, imag} */,
  {32'hbd8b2099, 32'h00000000} /* (5, 8, 31) {real, imag} */,
  {32'hbeb42363, 32'h00000000} /* (5, 8, 30) {real, imag} */,
  {32'hbea956ed, 32'h00000000} /* (5, 8, 29) {real, imag} */,
  {32'hbf2f9e2b, 32'h00000000} /* (5, 8, 28) {real, imag} */,
  {32'hbee41fca, 32'h00000000} /* (5, 8, 27) {real, imag} */,
  {32'hbee6fb34, 32'h00000000} /* (5, 8, 26) {real, imag} */,
  {32'hbf861cb8, 32'h00000000} /* (5, 8, 25) {real, imag} */,
  {32'hbed79147, 32'h00000000} /* (5, 8, 24) {real, imag} */,
  {32'h3e82322f, 32'h00000000} /* (5, 8, 23) {real, imag} */,
  {32'hbe20fe51, 32'h00000000} /* (5, 8, 22) {real, imag} */,
  {32'h3e0219ce, 32'h00000000} /* (5, 8, 21) {real, imag} */,
  {32'h3f1212ed, 32'h00000000} /* (5, 8, 20) {real, imag} */,
  {32'h3f0d30cd, 32'h00000000} /* (5, 8, 19) {real, imag} */,
  {32'h3f442d45, 32'h00000000} /* (5, 8, 18) {real, imag} */,
  {32'h3f317ae9, 32'h00000000} /* (5, 8, 17) {real, imag} */,
  {32'h3ef966c5, 32'h00000000} /* (5, 8, 16) {real, imag} */,
  {32'h3f2f5aca, 32'h00000000} /* (5, 8, 15) {real, imag} */,
  {32'hbebdc019, 32'h00000000} /* (5, 8, 14) {real, imag} */,
  {32'hbf34adf3, 32'h00000000} /* (5, 8, 13) {real, imag} */,
  {32'h3ddca051, 32'h00000000} /* (5, 8, 12) {real, imag} */,
  {32'h3f2aa0d4, 32'h00000000} /* (5, 8, 11) {real, imag} */,
  {32'h3d853580, 32'h00000000} /* (5, 8, 10) {real, imag} */,
  {32'hbeacad10, 32'h00000000} /* (5, 8, 9) {real, imag} */,
  {32'hbe06c013, 32'h00000000} /* (5, 8, 8) {real, imag} */,
  {32'h3d35152e, 32'h00000000} /* (5, 8, 7) {real, imag} */,
  {32'hbf08d48d, 32'h00000000} /* (5, 8, 6) {real, imag} */,
  {32'hbf3f07ae, 32'h00000000} /* (5, 8, 5) {real, imag} */,
  {32'hbee8d59f, 32'h00000000} /* (5, 8, 4) {real, imag} */,
  {32'h3d5f4aac, 32'h00000000} /* (5, 8, 3) {real, imag} */,
  {32'h3d94bb34, 32'h00000000} /* (5, 8, 2) {real, imag} */,
  {32'h3bc4f83b, 32'h00000000} /* (5, 8, 1) {real, imag} */,
  {32'hbde35e4f, 32'h00000000} /* (5, 8, 0) {real, imag} */,
  {32'h3d47cda4, 32'h00000000} /* (5, 7, 31) {real, imag} */,
  {32'hbe8d8d7f, 32'h00000000} /* (5, 7, 30) {real, imag} */,
  {32'hbf04fbbd, 32'h00000000} /* (5, 7, 29) {real, imag} */,
  {32'hbf08b603, 32'h00000000} /* (5, 7, 28) {real, imag} */,
  {32'hbef528b7, 32'h00000000} /* (5, 7, 27) {real, imag} */,
  {32'hbed455d2, 32'h00000000} /* (5, 7, 26) {real, imag} */,
  {32'hbfa25ec6, 32'h00000000} /* (5, 7, 25) {real, imag} */,
  {32'hbf87e7a7, 32'h00000000} /* (5, 7, 24) {real, imag} */,
  {32'h3e983855, 32'h00000000} /* (5, 7, 23) {real, imag} */,
  {32'h3e7902c4, 32'h00000000} /* (5, 7, 22) {real, imag} */,
  {32'h3ccb8377, 32'h00000000} /* (5, 7, 21) {real, imag} */,
  {32'h3f3f4d4e, 32'h00000000} /* (5, 7, 20) {real, imag} */,
  {32'h3f1f54d8, 32'h00000000} /* (5, 7, 19) {real, imag} */,
  {32'h3f4626df, 32'h00000000} /* (5, 7, 18) {real, imag} */,
  {32'h3f617285, 32'h00000000} /* (5, 7, 17) {real, imag} */,
  {32'h3f25be08, 32'h00000000} /* (5, 7, 16) {real, imag} */,
  {32'h3e096953, 32'h00000000} /* (5, 7, 15) {real, imag} */,
  {32'hbf241c7a, 32'h00000000} /* (5, 7, 14) {real, imag} */,
  {32'hbf3b6b91, 32'h00000000} /* (5, 7, 13) {real, imag} */,
  {32'h3e4ec7bb, 32'h00000000} /* (5, 7, 12) {real, imag} */,
  {32'h3f33611d, 32'h00000000} /* (5, 7, 11) {real, imag} */,
  {32'hbe2842ae, 32'h00000000} /* (5, 7, 10) {real, imag} */,
  {32'hbe35e686, 32'h00000000} /* (5, 7, 9) {real, imag} */,
  {32'h3ea2d9b4, 32'h00000000} /* (5, 7, 8) {real, imag} */,
  {32'h3cbf643f, 32'h00000000} /* (5, 7, 7) {real, imag} */,
  {32'hbf59400d, 32'h00000000} /* (5, 7, 6) {real, imag} */,
  {32'hbf261b26, 32'h00000000} /* (5, 7, 5) {real, imag} */,
  {32'hbf1f2ac5, 32'h00000000} /* (5, 7, 4) {real, imag} */,
  {32'h3ccea4f0, 32'h00000000} /* (5, 7, 3) {real, imag} */,
  {32'h3f33d690, 32'h00000000} /* (5, 7, 2) {real, imag} */,
  {32'h3c04e3a6, 32'h00000000} /* (5, 7, 1) {real, imag} */,
  {32'hbe6e5c68, 32'h00000000} /* (5, 7, 0) {real, imag} */,
  {32'hbe073412, 32'h00000000} /* (5, 6, 31) {real, imag} */,
  {32'h3d09ddd0, 32'h00000000} /* (5, 6, 30) {real, imag} */,
  {32'hbf701487, 32'h00000000} /* (5, 6, 29) {real, imag} */,
  {32'hbf237d74, 32'h00000000} /* (5, 6, 28) {real, imag} */,
  {32'hbd21f94e, 32'h00000000} /* (5, 6, 27) {real, imag} */,
  {32'hbdd5b884, 32'h00000000} /* (5, 6, 26) {real, imag} */,
  {32'hbe7209b2, 32'h00000000} /* (5, 6, 25) {real, imag} */,
  {32'hbe8b96f2, 32'h00000000} /* (5, 6, 24) {real, imag} */,
  {32'h3eba4324, 32'h00000000} /* (5, 6, 23) {real, imag} */,
  {32'h3f0ac02e, 32'h00000000} /* (5, 6, 22) {real, imag} */,
  {32'h3cfde7b2, 32'h00000000} /* (5, 6, 21) {real, imag} */,
  {32'hbe5ccdec, 32'h00000000} /* (5, 6, 20) {real, imag} */,
  {32'hbcb33090, 32'h00000000} /* (5, 6, 19) {real, imag} */,
  {32'h3e37658f, 32'h00000000} /* (5, 6, 18) {real, imag} */,
  {32'h3e13a050, 32'h00000000} /* (5, 6, 17) {real, imag} */,
  {32'h3e9a6256, 32'h00000000} /* (5, 6, 16) {real, imag} */,
  {32'hbd539d7a, 32'h00000000} /* (5, 6, 15) {real, imag} */,
  {32'h3ebac332, 32'h00000000} /* (5, 6, 14) {real, imag} */,
  {32'h3e33fc2f, 32'h00000000} /* (5, 6, 13) {real, imag} */,
  {32'h3e3246d1, 32'h00000000} /* (5, 6, 12) {real, imag} */,
  {32'h3f025bf8, 32'h00000000} /* (5, 6, 11) {real, imag} */,
  {32'h3edf3a98, 32'h00000000} /* (5, 6, 10) {real, imag} */,
  {32'h3eb3ca91, 32'h00000000} /* (5, 6, 9) {real, imag} */,
  {32'h3eae696c, 32'h00000000} /* (5, 6, 8) {real, imag} */,
  {32'hbd359d68, 32'h00000000} /* (5, 6, 7) {real, imag} */,
  {32'hbe83350a, 32'h00000000} /* (5, 6, 6) {real, imag} */,
  {32'h3eb628ba, 32'h00000000} /* (5, 6, 5) {real, imag} */,
  {32'hbda00d5a, 32'h00000000} /* (5, 6, 4) {real, imag} */,
  {32'hbe4a2475, 32'h00000000} /* (5, 6, 3) {real, imag} */,
  {32'h3dc1bbc8, 32'h00000000} /* (5, 6, 2) {real, imag} */,
  {32'hbe74ee80, 32'h00000000} /* (5, 6, 1) {real, imag} */,
  {32'hbe94fabd, 32'h00000000} /* (5, 6, 0) {real, imag} */,
  {32'h3e8586bc, 32'h00000000} /* (5, 5, 31) {real, imag} */,
  {32'h3e2154d5, 32'h00000000} /* (5, 5, 30) {real, imag} */,
  {32'hbf1252e1, 32'h00000000} /* (5, 5, 29) {real, imag} */,
  {32'hbf1eadcb, 32'h00000000} /* (5, 5, 28) {real, imag} */,
  {32'hbd5ad7db, 32'h00000000} /* (5, 5, 27) {real, imag} */,
  {32'hbdd0cb00, 32'h00000000} /* (5, 5, 26) {real, imag} */,
  {32'hbef475a6, 32'h00000000} /* (5, 5, 25) {real, imag} */,
  {32'hbe8fa70b, 32'h00000000} /* (5, 5, 24) {real, imag} */,
  {32'h3def1819, 32'h00000000} /* (5, 5, 23) {real, imag} */,
  {32'h3e0c10e0, 32'h00000000} /* (5, 5, 22) {real, imag} */,
  {32'hbe848ca1, 32'h00000000} /* (5, 5, 21) {real, imag} */,
  {32'hbf4cafd2, 32'h00000000} /* (5, 5, 20) {real, imag} */,
  {32'hbf207ad5, 32'h00000000} /* (5, 5, 19) {real, imag} */,
  {32'hbe8f7e30, 32'h00000000} /* (5, 5, 18) {real, imag} */,
  {32'hbf12b3f0, 32'h00000000} /* (5, 5, 17) {real, imag} */,
  {32'hbdc9c290, 32'h00000000} /* (5, 5, 16) {real, imag} */,
  {32'hbd988914, 32'h00000000} /* (5, 5, 15) {real, imag} */,
  {32'h3ec4c79b, 32'h00000000} /* (5, 5, 14) {real, imag} */,
  {32'h3dd2e0f2, 32'h00000000} /* (5, 5, 13) {real, imag} */,
  {32'h3eae45a0, 32'h00000000} /* (5, 5, 12) {real, imag} */,
  {32'hbe3056e2, 32'h00000000} /* (5, 5, 11) {real, imag} */,
  {32'h3e4f7efa, 32'h00000000} /* (5, 5, 10) {real, imag} */,
  {32'h3d883ed9, 32'h00000000} /* (5, 5, 9) {real, imag} */,
  {32'hbd5b5216, 32'h00000000} /* (5, 5, 8) {real, imag} */,
  {32'h3e1d17d3, 32'h00000000} /* (5, 5, 7) {real, imag} */,
  {32'h3dadcce2, 32'h00000000} /* (5, 5, 6) {real, imag} */,
  {32'h3f0c9cf5, 32'h00000000} /* (5, 5, 5) {real, imag} */,
  {32'h3e895816, 32'h00000000} /* (5, 5, 4) {real, imag} */,
  {32'hbad0b1fa, 32'h00000000} /* (5, 5, 3) {real, imag} */,
  {32'hbe5759b0, 32'h00000000} /* (5, 5, 2) {real, imag} */,
  {32'hbe9399b9, 32'h00000000} /* (5, 5, 1) {real, imag} */,
  {32'hbe221ee2, 32'h00000000} /* (5, 5, 0) {real, imag} */,
  {32'hbd46bb38, 32'h00000000} /* (5, 4, 31) {real, imag} */,
  {32'hbe422d0d, 32'h00000000} /* (5, 4, 30) {real, imag} */,
  {32'hbf19653a, 32'h00000000} /* (5, 4, 29) {real, imag} */,
  {32'hbf34b6ba, 32'h00000000} /* (5, 4, 28) {real, imag} */,
  {32'hbe43b5b0, 32'h00000000} /* (5, 4, 27) {real, imag} */,
  {32'hbd9775ad, 32'h00000000} /* (5, 4, 26) {real, imag} */,
  {32'hbec299e7, 32'h00000000} /* (5, 4, 25) {real, imag} */,
  {32'hbf2be870, 32'h00000000} /* (5, 4, 24) {real, imag} */,
  {32'hbe4c4f20, 32'h00000000} /* (5, 4, 23) {real, imag} */,
  {32'hbcf5b479, 32'h00000000} /* (5, 4, 22) {real, imag} */,
  {32'hbeff51cf, 32'h00000000} /* (5, 4, 21) {real, imag} */,
  {32'hbe5e7049, 32'h00000000} /* (5, 4, 20) {real, imag} */,
  {32'hbf196443, 32'h00000000} /* (5, 4, 19) {real, imag} */,
  {32'hbefe12b9, 32'h00000000} /* (5, 4, 18) {real, imag} */,
  {32'hbe80485a, 32'h00000000} /* (5, 4, 17) {real, imag} */,
  {32'hbea889aa, 32'h00000000} /* (5, 4, 16) {real, imag} */,
  {32'hbf2d457c, 32'h00000000} /* (5, 4, 15) {real, imag} */,
  {32'hbe3ad003, 32'h00000000} /* (5, 4, 14) {real, imag} */,
  {32'hbd32e500, 32'h00000000} /* (5, 4, 13) {real, imag} */,
  {32'hbdb0329b, 32'h00000000} /* (5, 4, 12) {real, imag} */,
  {32'hbe783c01, 32'h00000000} /* (5, 4, 11) {real, imag} */,
  {32'hbc0bac91, 32'h00000000} /* (5, 4, 10) {real, imag} */,
  {32'h3d0af70e, 32'h00000000} /* (5, 4, 9) {real, imag} */,
  {32'hbe5782a5, 32'h00000000} /* (5, 4, 8) {real, imag} */,
  {32'h3d38165f, 32'h00000000} /* (5, 4, 7) {real, imag} */,
  {32'h3e426aaf, 32'h00000000} /* (5, 4, 6) {real, imag} */,
  {32'h3df84bda, 32'h00000000} /* (5, 4, 5) {real, imag} */,
  {32'hbc3d6544, 32'h00000000} /* (5, 4, 4) {real, imag} */,
  {32'hbeebd331, 32'h00000000} /* (5, 4, 3) {real, imag} */,
  {32'hbec726e8, 32'h00000000} /* (5, 4, 2) {real, imag} */,
  {32'h3e0e30ba, 32'h00000000} /* (5, 4, 1) {real, imag} */,
  {32'h3e4ab7c4, 32'h00000000} /* (5, 4, 0) {real, imag} */,
  {32'hbe8967a8, 32'h00000000} /* (5, 3, 31) {real, imag} */,
  {32'hbde9e6c0, 32'h00000000} /* (5, 3, 30) {real, imag} */,
  {32'hbeda6876, 32'h00000000} /* (5, 3, 29) {real, imag} */,
  {32'hbf1fa6a3, 32'h00000000} /* (5, 3, 28) {real, imag} */,
  {32'hbdadf8b8, 32'h00000000} /* (5, 3, 27) {real, imag} */,
  {32'h3d41d4c9, 32'h00000000} /* (5, 3, 26) {real, imag} */,
  {32'h3e848caa, 32'h00000000} /* (5, 3, 25) {real, imag} */,
  {32'hbec93305, 32'h00000000} /* (5, 3, 24) {real, imag} */,
  {32'hbf180c56, 32'h00000000} /* (5, 3, 23) {real, imag} */,
  {32'hbe3da261, 32'h00000000} /* (5, 3, 22) {real, imag} */,
  {32'hbe64137b, 32'h00000000} /* (5, 3, 21) {real, imag} */,
  {32'h3dbc917b, 32'h00000000} /* (5, 3, 20) {real, imag} */,
  {32'hbe7432fd, 32'h00000000} /* (5, 3, 19) {real, imag} */,
  {32'hbeda160c, 32'h00000000} /* (5, 3, 18) {real, imag} */,
  {32'hbe73d0e5, 32'h00000000} /* (5, 3, 17) {real, imag} */,
  {32'hbf14190c, 32'h00000000} /* (5, 3, 16) {real, imag} */,
  {32'hbe91c4d3, 32'h00000000} /* (5, 3, 15) {real, imag} */,
  {32'hbda7c055, 32'h00000000} /* (5, 3, 14) {real, imag} */,
  {32'h3cbd340a, 32'h00000000} /* (5, 3, 13) {real, imag} */,
  {32'hbe06a741, 32'h00000000} /* (5, 3, 12) {real, imag} */,
  {32'hbda612d2, 32'h00000000} /* (5, 3, 11) {real, imag} */,
  {32'hbd7e6846, 32'h00000000} /* (5, 3, 10) {real, imag} */,
  {32'hbd805632, 32'h00000000} /* (5, 3, 9) {real, imag} */,
  {32'hbe694cb3, 32'h00000000} /* (5, 3, 8) {real, imag} */,
  {32'hbbf49dd4, 32'h00000000} /* (5, 3, 7) {real, imag} */,
  {32'hbe9e087f, 32'h00000000} /* (5, 3, 6) {real, imag} */,
  {32'hbea69c43, 32'h00000000} /* (5, 3, 5) {real, imag} */,
  {32'hbc9ce244, 32'h00000000} /* (5, 3, 4) {real, imag} */,
  {32'hbf391829, 32'h00000000} /* (5, 3, 3) {real, imag} */,
  {32'hbf34d2eb, 32'h00000000} /* (5, 3, 2) {real, imag} */,
  {32'hbc94ec4b, 32'h00000000} /* (5, 3, 1) {real, imag} */,
  {32'h3e67b864, 32'h00000000} /* (5, 3, 0) {real, imag} */,
  {32'h3d72c788, 32'h00000000} /* (5, 2, 31) {real, imag} */,
  {32'h3eb47f00, 32'h00000000} /* (5, 2, 30) {real, imag} */,
  {32'hbe27e48b, 32'h00000000} /* (5, 2, 29) {real, imag} */,
  {32'hbf1b6266, 32'h00000000} /* (5, 2, 28) {real, imag} */,
  {32'hbe8bb91a, 32'h00000000} /* (5, 2, 27) {real, imag} */,
  {32'hbea98404, 32'h00000000} /* (5, 2, 26) {real, imag} */,
  {32'hbdc0372e, 32'h00000000} /* (5, 2, 25) {real, imag} */,
  {32'h3d0112b4, 32'h00000000} /* (5, 2, 24) {real, imag} */,
  {32'hbf077178, 32'h00000000} /* (5, 2, 23) {real, imag} */,
  {32'h3cf127aa, 32'h00000000} /* (5, 2, 22) {real, imag} */,
  {32'h3a86a6cc, 32'h00000000} /* (5, 2, 21) {real, imag} */,
  {32'hbe712c76, 32'h00000000} /* (5, 2, 20) {real, imag} */,
  {32'hbeac8e40, 32'h00000000} /* (5, 2, 19) {real, imag} */,
  {32'hbed55977, 32'h00000000} /* (5, 2, 18) {real, imag} */,
  {32'hbea1f5b6, 32'h00000000} /* (5, 2, 17) {real, imag} */,
  {32'h3d8e6f73, 32'h00000000} /* (5, 2, 16) {real, imag} */,
  {32'h3ed19388, 32'h00000000} /* (5, 2, 15) {real, imag} */,
  {32'hbc6afed4, 32'h00000000} /* (5, 2, 14) {real, imag} */,
  {32'h3e52550b, 32'h00000000} /* (5, 2, 13) {real, imag} */,
  {32'h3f182a34, 32'h00000000} /* (5, 2, 12) {real, imag} */,
  {32'h3ea816cd, 32'h00000000} /* (5, 2, 11) {real, imag} */,
  {32'hbe7bbada, 32'h00000000} /* (5, 2, 10) {real, imag} */,
  {32'h3e1a4165, 32'h00000000} /* (5, 2, 9) {real, imag} */,
  {32'h3d86898e, 32'h00000000} /* (5, 2, 8) {real, imag} */,
  {32'h3da71b2c, 32'h00000000} /* (5, 2, 7) {real, imag} */,
  {32'hbe0ed9cb, 32'h00000000} /* (5, 2, 6) {real, imag} */,
  {32'hbed30c4c, 32'h00000000} /* (5, 2, 5) {real, imag} */,
  {32'hbeff6a1b, 32'h00000000} /* (5, 2, 4) {real, imag} */,
  {32'hbed96c20, 32'h00000000} /* (5, 2, 3) {real, imag} */,
  {32'hbe1d5cef, 32'h00000000} /* (5, 2, 2) {real, imag} */,
  {32'hbec13361, 32'h00000000} /* (5, 2, 1) {real, imag} */,
  {32'hbea81383, 32'h00000000} /* (5, 2, 0) {real, imag} */,
  {32'h3c4c767c, 32'h00000000} /* (5, 1, 31) {real, imag} */,
  {32'h3e4112f8, 32'h00000000} /* (5, 1, 30) {real, imag} */,
  {32'h3e41d060, 32'h00000000} /* (5, 1, 29) {real, imag} */,
  {32'h3c9423f9, 32'h00000000} /* (5, 1, 28) {real, imag} */,
  {32'hbeb02fc7, 32'h00000000} /* (5, 1, 27) {real, imag} */,
  {32'hbf62dc73, 32'h00000000} /* (5, 1, 26) {real, imag} */,
  {32'hbf0dbd4c, 32'h00000000} /* (5, 1, 25) {real, imag} */,
  {32'h3e44a85a, 32'h00000000} /* (5, 1, 24) {real, imag} */,
  {32'hbe58479b, 32'h00000000} /* (5, 1, 23) {real, imag} */,
  {32'hbf1bdd9d, 32'h00000000} /* (5, 1, 22) {real, imag} */,
  {32'hbef875ba, 32'h00000000} /* (5, 1, 21) {real, imag} */,
  {32'hbecadd34, 32'h00000000} /* (5, 1, 20) {real, imag} */,
  {32'hbeea280a, 32'h00000000} /* (5, 1, 19) {real, imag} */,
  {32'hbf79c5e1, 32'h00000000} /* (5, 1, 18) {real, imag} */,
  {32'hbf34cd3b, 32'h00000000} /* (5, 1, 17) {real, imag} */,
  {32'h3e90deca, 32'h00000000} /* (5, 1, 16) {real, imag} */,
  {32'h3edef159, 32'h00000000} /* (5, 1, 15) {real, imag} */,
  {32'h3edfed62, 32'h00000000} /* (5, 1, 14) {real, imag} */,
  {32'h3ddad820, 32'h00000000} /* (5, 1, 13) {real, imag} */,
  {32'h3e79d0ab, 32'h00000000} /* (5, 1, 12) {real, imag} */,
  {32'h3f02da69, 32'h00000000} /* (5, 1, 11) {real, imag} */,
  {32'h3ed72654, 32'h00000000} /* (5, 1, 10) {real, imag} */,
  {32'h3edfa4e7, 32'h00000000} /* (5, 1, 9) {real, imag} */,
  {32'h3e967f51, 32'h00000000} /* (5, 1, 8) {real, imag} */,
  {32'h3e5afc8c, 32'h00000000} /* (5, 1, 7) {real, imag} */,
  {32'hbd515934, 32'h00000000} /* (5, 1, 6) {real, imag} */,
  {32'hbf1a4132, 32'h00000000} /* (5, 1, 5) {real, imag} */,
  {32'hbf1c5cd7, 32'h00000000} /* (5, 1, 4) {real, imag} */,
  {32'hbebb72a5, 32'h00000000} /* (5, 1, 3) {real, imag} */,
  {32'hbe323454, 32'h00000000} /* (5, 1, 2) {real, imag} */,
  {32'hbe79ce77, 32'h00000000} /* (5, 1, 1) {real, imag} */,
  {32'hbe9c6cdf, 32'h00000000} /* (5, 1, 0) {real, imag} */,
  {32'h3d51a943, 32'h00000000} /* (5, 0, 31) {real, imag} */,
  {32'h3e9313fa, 32'h00000000} /* (5, 0, 30) {real, imag} */,
  {32'h3e2171f9, 32'h00000000} /* (5, 0, 29) {real, imag} */,
  {32'h3e3fac4b, 32'h00000000} /* (5, 0, 28) {real, imag} */,
  {32'h3dbefd89, 32'h00000000} /* (5, 0, 27) {real, imag} */,
  {32'hbee1dd99, 32'h00000000} /* (5, 0, 26) {real, imag} */,
  {32'hbdf5767e, 32'h00000000} /* (5, 0, 25) {real, imag} */,
  {32'h3e9b4970, 32'h00000000} /* (5, 0, 24) {real, imag} */,
  {32'hbd0cb8e3, 32'h00000000} /* (5, 0, 23) {real, imag} */,
  {32'hbe87ae32, 32'h00000000} /* (5, 0, 22) {real, imag} */,
  {32'hbd4e66f2, 32'h00000000} /* (5, 0, 21) {real, imag} */,
  {32'hbdba69d4, 32'h00000000} /* (5, 0, 20) {real, imag} */,
  {32'hbe47ec88, 32'h00000000} /* (5, 0, 19) {real, imag} */,
  {32'hbef48588, 32'h00000000} /* (5, 0, 18) {real, imag} */,
  {32'hbe8d403b, 32'h00000000} /* (5, 0, 17) {real, imag} */,
  {32'h3dbc56c1, 32'h00000000} /* (5, 0, 16) {real, imag} */,
  {32'h3c723a45, 32'h00000000} /* (5, 0, 15) {real, imag} */,
  {32'h3e8ce7ad, 32'h00000000} /* (5, 0, 14) {real, imag} */,
  {32'h3e6680df, 32'h00000000} /* (5, 0, 13) {real, imag} */,
  {32'h3e8c154d, 32'h00000000} /* (5, 0, 12) {real, imag} */,
  {32'h3e73e5b2, 32'h00000000} /* (5, 0, 11) {real, imag} */,
  {32'h3e57e84f, 32'h00000000} /* (5, 0, 10) {real, imag} */,
  {32'hbe1670c5, 32'h00000000} /* (5, 0, 9) {real, imag} */,
  {32'hbe188528, 32'h00000000} /* (5, 0, 8) {real, imag} */,
  {32'hbe921cf8, 32'h00000000} /* (5, 0, 7) {real, imag} */,
  {32'hbeb1f6dc, 32'h00000000} /* (5, 0, 6) {real, imag} */,
  {32'hbeb827a6, 32'h00000000} /* (5, 0, 5) {real, imag} */,
  {32'hbec54be9, 32'h00000000} /* (5, 0, 4) {real, imag} */,
  {32'hbdefdeac, 32'h00000000} /* (5, 0, 3) {real, imag} */,
  {32'hbdbc20dd, 32'h00000000} /* (5, 0, 2) {real, imag} */,
  {32'hbdff8623, 32'h00000000} /* (5, 0, 1) {real, imag} */,
  {32'hbe4fdb58, 32'h00000000} /* (5, 0, 0) {real, imag} */,
  {32'hbe8e35bf, 32'h00000000} /* (4, 31, 31) {real, imag} */,
  {32'hbe457aaf, 32'h00000000} /* (4, 31, 30) {real, imag} */,
  {32'hbe808c10, 32'h00000000} /* (4, 31, 29) {real, imag} */,
  {32'hbf020f35, 32'h00000000} /* (4, 31, 28) {real, imag} */,
  {32'hbf4ad84e, 32'h00000000} /* (4, 31, 27) {real, imag} */,
  {32'hbf8e2cc7, 32'h00000000} /* (4, 31, 26) {real, imag} */,
  {32'hbf6af369, 32'h00000000} /* (4, 31, 25) {real, imag} */,
  {32'hbf81f318, 32'h00000000} /* (4, 31, 24) {real, imag} */,
  {32'hbf0df28c, 32'h00000000} /* (4, 31, 23) {real, imag} */,
  {32'hbe97a779, 32'h00000000} /* (4, 31, 22) {real, imag} */,
  {32'hbd1f27c5, 32'h00000000} /* (4, 31, 21) {real, imag} */,
  {32'h3e90fee8, 32'h00000000} /* (4, 31, 20) {real, imag} */,
  {32'h3f22d22e, 32'h00000000} /* (4, 31, 19) {real, imag} */,
  {32'h3ec8791f, 32'h00000000} /* (4, 31, 18) {real, imag} */,
  {32'h3ec28dc4, 32'h00000000} /* (4, 31, 17) {real, imag} */,
  {32'h3e3a361a, 32'h00000000} /* (4, 31, 16) {real, imag} */,
  {32'h3e740c8d, 32'h00000000} /* (4, 31, 15) {real, imag} */,
  {32'h3ebeba07, 32'h00000000} /* (4, 31, 14) {real, imag} */,
  {32'h3f84fad1, 32'h00000000} /* (4, 31, 13) {real, imag} */,
  {32'h3f154ee7, 32'h00000000} /* (4, 31, 12) {real, imag} */,
  {32'h3e8cec1e, 32'h00000000} /* (4, 31, 11) {real, imag} */,
  {32'hbea97b65, 32'h00000000} /* (4, 31, 10) {real, imag} */,
  {32'hbeefe633, 32'h00000000} /* (4, 31, 9) {real, imag} */,
  {32'hbed676c7, 32'h00000000} /* (4, 31, 8) {real, imag} */,
  {32'hbecf043d, 32'h00000000} /* (4, 31, 7) {real, imag} */,
  {32'hbf188e22, 32'h00000000} /* (4, 31, 6) {real, imag} */,
  {32'hbf0bd5fe, 32'h00000000} /* (4, 31, 5) {real, imag} */,
  {32'hbecd67bc, 32'h00000000} /* (4, 31, 4) {real, imag} */,
  {32'hbf025801, 32'h00000000} /* (4, 31, 3) {real, imag} */,
  {32'hbeaaee41, 32'h00000000} /* (4, 31, 2) {real, imag} */,
  {32'hbe86b408, 32'h00000000} /* (4, 31, 1) {real, imag} */,
  {32'hbe99d071, 32'h00000000} /* (4, 31, 0) {real, imag} */,
  {32'hbf2609f0, 32'h00000000} /* (4, 30, 31) {real, imag} */,
  {32'hbf5131c1, 32'h00000000} /* (4, 30, 30) {real, imag} */,
  {32'hbeecfa88, 32'h00000000} /* (4, 30, 29) {real, imag} */,
  {32'hbf31d516, 32'h00000000} /* (4, 30, 28) {real, imag} */,
  {32'hbf81bc75, 32'h00000000} /* (4, 30, 27) {real, imag} */,
  {32'hbfc69432, 32'h00000000} /* (4, 30, 26) {real, imag} */,
  {32'hbf9e4c0f, 32'h00000000} /* (4, 30, 25) {real, imag} */,
  {32'hbf8ce2a7, 32'h00000000} /* (4, 30, 24) {real, imag} */,
  {32'hbf689b52, 32'h00000000} /* (4, 30, 23) {real, imag} */,
  {32'hbf30d8dd, 32'h00000000} /* (4, 30, 22) {real, imag} */,
  {32'hbe4a3aca, 32'h00000000} /* (4, 30, 21) {real, imag} */,
  {32'h3eca4e04, 32'h00000000} /* (4, 30, 20) {real, imag} */,
  {32'h3f5f1366, 32'h00000000} /* (4, 30, 19) {real, imag} */,
  {32'h3f258660, 32'h00000000} /* (4, 30, 18) {real, imag} */,
  {32'h3f6b570d, 32'h00000000} /* (4, 30, 17) {real, imag} */,
  {32'h3f37812d, 32'h00000000} /* (4, 30, 16) {real, imag} */,
  {32'h3f58b243, 32'h00000000} /* (4, 30, 15) {real, imag} */,
  {32'h3f18d376, 32'h00000000} /* (4, 30, 14) {real, imag} */,
  {32'h3f886cde, 32'h00000000} /* (4, 30, 13) {real, imag} */,
  {32'h3f8c6280, 32'h00000000} /* (4, 30, 12) {real, imag} */,
  {32'h3f410c51, 32'h00000000} /* (4, 30, 11) {real, imag} */,
  {32'hbf106ce7, 32'h00000000} /* (4, 30, 10) {real, imag} */,
  {32'hbf65663a, 32'h00000000} /* (4, 30, 9) {real, imag} */,
  {32'hbf24227d, 32'h00000000} /* (4, 30, 8) {real, imag} */,
  {32'hbf826bed, 32'h00000000} /* (4, 30, 7) {real, imag} */,
  {32'hbfa98055, 32'h00000000} /* (4, 30, 6) {real, imag} */,
  {32'hbf8c2d5b, 32'h00000000} /* (4, 30, 5) {real, imag} */,
  {32'hbf6244f3, 32'h00000000} /* (4, 30, 4) {real, imag} */,
  {32'hbf15ad52, 32'h00000000} /* (4, 30, 3) {real, imag} */,
  {32'hbee54d80, 32'h00000000} /* (4, 30, 2) {real, imag} */,
  {32'hbf20e1cc, 32'h00000000} /* (4, 30, 1) {real, imag} */,
  {32'hbee4c0ca, 32'h00000000} /* (4, 30, 0) {real, imag} */,
  {32'hbf27efe4, 32'h00000000} /* (4, 29, 31) {real, imag} */,
  {32'hbfa4417c, 32'h00000000} /* (4, 29, 30) {real, imag} */,
  {32'hbf96f0ba, 32'h00000000} /* (4, 29, 29) {real, imag} */,
  {32'hbf07611f, 32'h00000000} /* (4, 29, 28) {real, imag} */,
  {32'hbf166ad2, 32'h00000000} /* (4, 29, 27) {real, imag} */,
  {32'hbf934ad4, 32'h00000000} /* (4, 29, 26) {real, imag} */,
  {32'hbfaa1837, 32'h00000000} /* (4, 29, 25) {real, imag} */,
  {32'hbf90d4df, 32'h00000000} /* (4, 29, 24) {real, imag} */,
  {32'hbf9f91aa, 32'h00000000} /* (4, 29, 23) {real, imag} */,
  {32'hbf64805e, 32'h00000000} /* (4, 29, 22) {real, imag} */,
  {32'hbe46ece2, 32'h00000000} /* (4, 29, 21) {real, imag} */,
  {32'h3ef8b430, 32'h00000000} /* (4, 29, 20) {real, imag} */,
  {32'h3f6eebf5, 32'h00000000} /* (4, 29, 19) {real, imag} */,
  {32'h3ef121ca, 32'h00000000} /* (4, 29, 18) {real, imag} */,
  {32'h3fab5bd0, 32'h00000000} /* (4, 29, 17) {real, imag} */,
  {32'h3fb96a88, 32'h00000000} /* (4, 29, 16) {real, imag} */,
  {32'h3f887153, 32'h00000000} /* (4, 29, 15) {real, imag} */,
  {32'h3eed6db5, 32'h00000000} /* (4, 29, 14) {real, imag} */,
  {32'h3f01f33f, 32'h00000000} /* (4, 29, 13) {real, imag} */,
  {32'h3f8cfc2d, 32'h00000000} /* (4, 29, 12) {real, imag} */,
  {32'h3f405ef4, 32'h00000000} /* (4, 29, 11) {real, imag} */,
  {32'hbf72d2cc, 32'h00000000} /* (4, 29, 10) {real, imag} */,
  {32'hbfa2a484, 32'h00000000} /* (4, 29, 9) {real, imag} */,
  {32'hbf530780, 32'h00000000} /* (4, 29, 8) {real, imag} */,
  {32'hbf82f96a, 32'h00000000} /* (4, 29, 7) {real, imag} */,
  {32'hbf7ca12d, 32'h00000000} /* (4, 29, 6) {real, imag} */,
  {32'hbf843d31, 32'h00000000} /* (4, 29, 5) {real, imag} */,
  {32'hbf9a187b, 32'h00000000} /* (4, 29, 4) {real, imag} */,
  {32'hbf086d89, 32'h00000000} /* (4, 29, 3) {real, imag} */,
  {32'hbe91d3fd, 32'h00000000} /* (4, 29, 2) {real, imag} */,
  {32'hbf4a6dea, 32'h00000000} /* (4, 29, 1) {real, imag} */,
  {32'hbf3e9594, 32'h00000000} /* (4, 29, 0) {real, imag} */,
  {32'hbe286fcf, 32'h00000000} /* (4, 28, 31) {real, imag} */,
  {32'hbf74eeff, 32'h00000000} /* (4, 28, 30) {real, imag} */,
  {32'hbfa2fe2d, 32'h00000000} /* (4, 28, 29) {real, imag} */,
  {32'hbf380a63, 32'h00000000} /* (4, 28, 28) {real, imag} */,
  {32'hbf429ade, 32'h00000000} /* (4, 28, 27) {real, imag} */,
  {32'hbf58d969, 32'h00000000} /* (4, 28, 26) {real, imag} */,
  {32'hbf6892e3, 32'h00000000} /* (4, 28, 25) {real, imag} */,
  {32'hbf75ac10, 32'h00000000} /* (4, 28, 24) {real, imag} */,
  {32'hbf58e834, 32'h00000000} /* (4, 28, 23) {real, imag} */,
  {32'hbf154bf6, 32'h00000000} /* (4, 28, 22) {real, imag} */,
  {32'h3ed313a3, 32'h00000000} /* (4, 28, 21) {real, imag} */,
  {32'h3f7d6c0b, 32'h00000000} /* (4, 28, 20) {real, imag} */,
  {32'h3f4f82d8, 32'h00000000} /* (4, 28, 19) {real, imag} */,
  {32'h3ea3438f, 32'h00000000} /* (4, 28, 18) {real, imag} */,
  {32'h3f2e6f33, 32'h00000000} /* (4, 28, 17) {real, imag} */,
  {32'h3f4f5b5c, 32'h00000000} /* (4, 28, 16) {real, imag} */,
  {32'h3f1486f9, 32'h00000000} /* (4, 28, 15) {real, imag} */,
  {32'h3e73028a, 32'h00000000} /* (4, 28, 14) {real, imag} */,
  {32'h3f09296b, 32'h00000000} /* (4, 28, 13) {real, imag} */,
  {32'h3f7d6697, 32'h00000000} /* (4, 28, 12) {real, imag} */,
  {32'h3f9429b7, 32'h00000000} /* (4, 28, 11) {real, imag} */,
  {32'hbd45ab9e, 32'h00000000} /* (4, 28, 10) {real, imag} */,
  {32'hbfa24158, 32'h00000000} /* (4, 28, 9) {real, imag} */,
  {32'hbfaa9de0, 32'h00000000} /* (4, 28, 8) {real, imag} */,
  {32'hbf57985e, 32'h00000000} /* (4, 28, 7) {real, imag} */,
  {32'hbf39fe1e, 32'h00000000} /* (4, 28, 6) {real, imag} */,
  {32'hbf3803f7, 32'h00000000} /* (4, 28, 5) {real, imag} */,
  {32'hbf62b7a6, 32'h00000000} /* (4, 28, 4) {real, imag} */,
  {32'hbf820de7, 32'h00000000} /* (4, 28, 3) {real, imag} */,
  {32'hbf453791, 32'h00000000} /* (4, 28, 2) {real, imag} */,
  {32'hbf4a2059, 32'h00000000} /* (4, 28, 1) {real, imag} */,
  {32'hbf10319a, 32'h00000000} /* (4, 28, 0) {real, imag} */,
  {32'hbe951164, 32'h00000000} /* (4, 27, 31) {real, imag} */,
  {32'hbf3c6a98, 32'h00000000} /* (4, 27, 30) {real, imag} */,
  {32'hbf204bc3, 32'h00000000} /* (4, 27, 29) {real, imag} */,
  {32'hbf6e3662, 32'h00000000} /* (4, 27, 28) {real, imag} */,
  {32'hbf73ff8a, 32'h00000000} /* (4, 27, 27) {real, imag} */,
  {32'hbf564f72, 32'h00000000} /* (4, 27, 26) {real, imag} */,
  {32'hbf8cccb1, 32'h00000000} /* (4, 27, 25) {real, imag} */,
  {32'hbfbfdc76, 32'h00000000} /* (4, 27, 24) {real, imag} */,
  {32'hbf6f1855, 32'h00000000} /* (4, 27, 23) {real, imag} */,
  {32'hbf659129, 32'h00000000} /* (4, 27, 22) {real, imag} */,
  {32'hbda043b6, 32'h00000000} /* (4, 27, 21) {real, imag} */,
  {32'h3f8b6c3a, 32'h00000000} /* (4, 27, 20) {real, imag} */,
  {32'h3f87df0d, 32'h00000000} /* (4, 27, 19) {real, imag} */,
  {32'h3f8597b4, 32'h00000000} /* (4, 27, 18) {real, imag} */,
  {32'h3f2750e4, 32'h00000000} /* (4, 27, 17) {real, imag} */,
  {32'h3ecb57bd, 32'h00000000} /* (4, 27, 16) {real, imag} */,
  {32'h3f9c0789, 32'h00000000} /* (4, 27, 15) {real, imag} */,
  {32'h3f280a2d, 32'h00000000} /* (4, 27, 14) {real, imag} */,
  {32'h3f4da19f, 32'h00000000} /* (4, 27, 13) {real, imag} */,
  {32'h3f9cb4f9, 32'h00000000} /* (4, 27, 12) {real, imag} */,
  {32'h3f9cf984, 32'h00000000} /* (4, 27, 11) {real, imag} */,
  {32'hbec27f6d, 32'h00000000} /* (4, 27, 10) {real, imag} */,
  {32'hbf6f1096, 32'h00000000} /* (4, 27, 9) {real, imag} */,
  {32'hbf532882, 32'h00000000} /* (4, 27, 8) {real, imag} */,
  {32'hbf0410d8, 32'h00000000} /* (4, 27, 7) {real, imag} */,
  {32'hbf5ad3fa, 32'h00000000} /* (4, 27, 6) {real, imag} */,
  {32'hbf25931d, 32'h00000000} /* (4, 27, 5) {real, imag} */,
  {32'hbeff497b, 32'h00000000} /* (4, 27, 4) {real, imag} */,
  {32'hbf639c67, 32'h00000000} /* (4, 27, 3) {real, imag} */,
  {32'hbf54ce1b, 32'h00000000} /* (4, 27, 2) {real, imag} */,
  {32'hbf768e75, 32'h00000000} /* (4, 27, 1) {real, imag} */,
  {32'hbf39cf9f, 32'h00000000} /* (4, 27, 0) {real, imag} */,
  {32'hbe74f6be, 32'h00000000} /* (4, 26, 31) {real, imag} */,
  {32'hbf34ebff, 32'h00000000} /* (4, 26, 30) {real, imag} */,
  {32'hbf398dfd, 32'h00000000} /* (4, 26, 29) {real, imag} */,
  {32'hbf2e4f63, 32'h00000000} /* (4, 26, 28) {real, imag} */,
  {32'hbf13d6f8, 32'h00000000} /* (4, 26, 27) {real, imag} */,
  {32'hbf6e5f05, 32'h00000000} /* (4, 26, 26) {real, imag} */,
  {32'hbfa233c4, 32'h00000000} /* (4, 26, 25) {real, imag} */,
  {32'hbfdfa7d3, 32'h00000000} /* (4, 26, 24) {real, imag} */,
  {32'hbfb8c016, 32'h00000000} /* (4, 26, 23) {real, imag} */,
  {32'hbf74227a, 32'h00000000} /* (4, 26, 22) {real, imag} */,
  {32'hbee1c1df, 32'h00000000} /* (4, 26, 21) {real, imag} */,
  {32'h3f0fd8da, 32'h00000000} /* (4, 26, 20) {real, imag} */,
  {32'h3f231fa0, 32'h00000000} /* (4, 26, 19) {real, imag} */,
  {32'h3f59d14e, 32'h00000000} /* (4, 26, 18) {real, imag} */,
  {32'h3f57c1bc, 32'h00000000} /* (4, 26, 17) {real, imag} */,
  {32'h3f087477, 32'h00000000} /* (4, 26, 16) {real, imag} */,
  {32'h3fb9739d, 32'h00000000} /* (4, 26, 15) {real, imag} */,
  {32'h3f9cb70d, 32'h00000000} /* (4, 26, 14) {real, imag} */,
  {32'h3f435122, 32'h00000000} /* (4, 26, 13) {real, imag} */,
  {32'h3f77e91e, 32'h00000000} /* (4, 26, 12) {real, imag} */,
  {32'h3efd8198, 32'h00000000} /* (4, 26, 11) {real, imag} */,
  {32'hbf0a58e4, 32'h00000000} /* (4, 26, 10) {real, imag} */,
  {32'hbf411cc9, 32'h00000000} /* (4, 26, 9) {real, imag} */,
  {32'hbf25d6ff, 32'h00000000} /* (4, 26, 8) {real, imag} */,
  {32'hbe9d90c3, 32'h00000000} /* (4, 26, 7) {real, imag} */,
  {32'hbedb9b35, 32'h00000000} /* (4, 26, 6) {real, imag} */,
  {32'hbf4ee434, 32'h00000000} /* (4, 26, 5) {real, imag} */,
  {32'hbf274bd4, 32'h00000000} /* (4, 26, 4) {real, imag} */,
  {32'hbed7d9e4, 32'h00000000} /* (4, 26, 3) {real, imag} */,
  {32'hbf38d04c, 32'h00000000} /* (4, 26, 2) {real, imag} */,
  {32'hbf0ced0a, 32'h00000000} /* (4, 26, 1) {real, imag} */,
  {32'hbe9edf35, 32'h00000000} /* (4, 26, 0) {real, imag} */,
  {32'hbef06293, 32'h00000000} /* (4, 25, 31) {real, imag} */,
  {32'hbf7ecf2c, 32'h00000000} /* (4, 25, 30) {real, imag} */,
  {32'hbf86f17c, 32'h00000000} /* (4, 25, 29) {real, imag} */,
  {32'hbf914bca, 32'h00000000} /* (4, 25, 28) {real, imag} */,
  {32'hbf8fbe89, 32'h00000000} /* (4, 25, 27) {real, imag} */,
  {32'hbfb7e9f3, 32'h00000000} /* (4, 25, 26) {real, imag} */,
  {32'hbfccf238, 32'h00000000} /* (4, 25, 25) {real, imag} */,
  {32'hbfb3c158, 32'h00000000} /* (4, 25, 24) {real, imag} */,
  {32'hbfb7ffdc, 32'h00000000} /* (4, 25, 23) {real, imag} */,
  {32'hbfb81913, 32'h00000000} /* (4, 25, 22) {real, imag} */,
  {32'hbf546472, 32'h00000000} /* (4, 25, 21) {real, imag} */,
  {32'h3f74840b, 32'h00000000} /* (4, 25, 20) {real, imag} */,
  {32'h3f796ed4, 32'h00000000} /* (4, 25, 19) {real, imag} */,
  {32'h3f3a6f8e, 32'h00000000} /* (4, 25, 18) {real, imag} */,
  {32'h3f540ce6, 32'h00000000} /* (4, 25, 17) {real, imag} */,
  {32'h3f435768, 32'h00000000} /* (4, 25, 16) {real, imag} */,
  {32'h3f936f0a, 32'h00000000} /* (4, 25, 15) {real, imag} */,
  {32'h3f5301e6, 32'h00000000} /* (4, 25, 14) {real, imag} */,
  {32'h3f1f4b0a, 32'h00000000} /* (4, 25, 13) {real, imag} */,
  {32'h3f17e47e, 32'h00000000} /* (4, 25, 12) {real, imag} */,
  {32'h3f3133ea, 32'h00000000} /* (4, 25, 11) {real, imag} */,
  {32'hbeb4c8a7, 32'h00000000} /* (4, 25, 10) {real, imag} */,
  {32'hbf54a3b1, 32'h00000000} /* (4, 25, 9) {real, imag} */,
  {32'hbfb5839a, 32'h00000000} /* (4, 25, 8) {real, imag} */,
  {32'hbf4a7773, 32'h00000000} /* (4, 25, 7) {real, imag} */,
  {32'hbf2e7382, 32'h00000000} /* (4, 25, 6) {real, imag} */,
  {32'hbfb6a8f3, 32'h00000000} /* (4, 25, 5) {real, imag} */,
  {32'hbf9adc48, 32'h00000000} /* (4, 25, 4) {real, imag} */,
  {32'hbf33a1fa, 32'h00000000} /* (4, 25, 3) {real, imag} */,
  {32'hbf9d2d96, 32'h00000000} /* (4, 25, 2) {real, imag} */,
  {32'hbf36723c, 32'h00000000} /* (4, 25, 1) {real, imag} */,
  {32'hbed72c2f, 32'h00000000} /* (4, 25, 0) {real, imag} */,
  {32'hbee2fa97, 32'h00000000} /* (4, 24, 31) {real, imag} */,
  {32'hbf86ac0d, 32'h00000000} /* (4, 24, 30) {real, imag} */,
  {32'hbfb082e1, 32'h00000000} /* (4, 24, 29) {real, imag} */,
  {32'hbfb6dcdf, 32'h00000000} /* (4, 24, 28) {real, imag} */,
  {32'hbf963044, 32'h00000000} /* (4, 24, 27) {real, imag} */,
  {32'hbfa91aa4, 32'h00000000} /* (4, 24, 26) {real, imag} */,
  {32'hbfa8b60b, 32'h00000000} /* (4, 24, 25) {real, imag} */,
  {32'hbf6e60f5, 32'h00000000} /* (4, 24, 24) {real, imag} */,
  {32'hbf732871, 32'h00000000} /* (4, 24, 23) {real, imag} */,
  {32'hbf728f6e, 32'h00000000} /* (4, 24, 22) {real, imag} */,
  {32'hbea99334, 32'h00000000} /* (4, 24, 21) {real, imag} */,
  {32'h3f9e0c5c, 32'h00000000} /* (4, 24, 20) {real, imag} */,
  {32'h3faa147c, 32'h00000000} /* (4, 24, 19) {real, imag} */,
  {32'h3fa0baaa, 32'h00000000} /* (4, 24, 18) {real, imag} */,
  {32'h3f7d3dc3, 32'h00000000} /* (4, 24, 17) {real, imag} */,
  {32'h3f932007, 32'h00000000} /* (4, 24, 16) {real, imag} */,
  {32'h3fb93ded, 32'h00000000} /* (4, 24, 15) {real, imag} */,
  {32'h3f8a9083, 32'h00000000} /* (4, 24, 14) {real, imag} */,
  {32'h3f3baf86, 32'h00000000} /* (4, 24, 13) {real, imag} */,
  {32'h3f15b86b, 32'h00000000} /* (4, 24, 12) {real, imag} */,
  {32'h3f48bd1f, 32'h00000000} /* (4, 24, 11) {real, imag} */,
  {32'hbeef76d1, 32'h00000000} /* (4, 24, 10) {real, imag} */,
  {32'hbf81ae60, 32'h00000000} /* (4, 24, 9) {real, imag} */,
  {32'hbf9d507e, 32'h00000000} /* (4, 24, 8) {real, imag} */,
  {32'hbf1d0871, 32'h00000000} /* (4, 24, 7) {real, imag} */,
  {32'hbf33745b, 32'h00000000} /* (4, 24, 6) {real, imag} */,
  {32'hbf52b063, 32'h00000000} /* (4, 24, 5) {real, imag} */,
  {32'hbefc092a, 32'h00000000} /* (4, 24, 4) {real, imag} */,
  {32'hbef35ec0, 32'h00000000} /* (4, 24, 3) {real, imag} */,
  {32'hbfa7ce79, 32'h00000000} /* (4, 24, 2) {real, imag} */,
  {32'hbfa47f8e, 32'h00000000} /* (4, 24, 1) {real, imag} */,
  {32'hbf4917e2, 32'h00000000} /* (4, 24, 0) {real, imag} */,
  {32'hbf43835c, 32'h00000000} /* (4, 23, 31) {real, imag} */,
  {32'hbf91c995, 32'h00000000} /* (4, 23, 30) {real, imag} */,
  {32'hbf9635ce, 32'h00000000} /* (4, 23, 29) {real, imag} */,
  {32'hbfb523fb, 32'h00000000} /* (4, 23, 28) {real, imag} */,
  {32'hbfbc6206, 32'h00000000} /* (4, 23, 27) {real, imag} */,
  {32'hbf800b61, 32'h00000000} /* (4, 23, 26) {real, imag} */,
  {32'hbf894120, 32'h00000000} /* (4, 23, 25) {real, imag} */,
  {32'hbf8ce0b9, 32'h00000000} /* (4, 23, 24) {real, imag} */,
  {32'hbf69d79b, 32'h00000000} /* (4, 23, 23) {real, imag} */,
  {32'hbf4008bf, 32'h00000000} /* (4, 23, 22) {real, imag} */,
  {32'h3bb97e96, 32'h00000000} /* (4, 23, 21) {real, imag} */,
  {32'h3f998a1a, 32'h00000000} /* (4, 23, 20) {real, imag} */,
  {32'h3f9a5750, 32'h00000000} /* (4, 23, 19) {real, imag} */,
  {32'h3fcbffcf, 32'h00000000} /* (4, 23, 18) {real, imag} */,
  {32'h3fc6e5d9, 32'h00000000} /* (4, 23, 17) {real, imag} */,
  {32'h3f84b6eb, 32'h00000000} /* (4, 23, 16) {real, imag} */,
  {32'h3f90c506, 32'h00000000} /* (4, 23, 15) {real, imag} */,
  {32'h3fa9ac83, 32'h00000000} /* (4, 23, 14) {real, imag} */,
  {32'h3f494b5c, 32'h00000000} /* (4, 23, 13) {real, imag} */,
  {32'h3eed5b7c, 32'h00000000} /* (4, 23, 12) {real, imag} */,
  {32'h3f36213c, 32'h00000000} /* (4, 23, 11) {real, imag} */,
  {32'hbf16e1e5, 32'h00000000} /* (4, 23, 10) {real, imag} */,
  {32'hbfb90eab, 32'h00000000} /* (4, 23, 9) {real, imag} */,
  {32'hbfbe5f21, 32'h00000000} /* (4, 23, 8) {real, imag} */,
  {32'hbf7c25a0, 32'h00000000} /* (4, 23, 7) {real, imag} */,
  {32'hbf4c2c82, 32'h00000000} /* (4, 23, 6) {real, imag} */,
  {32'hbf25df35, 32'h00000000} /* (4, 23, 5) {real, imag} */,
  {32'hbec07dc6, 32'h00000000} /* (4, 23, 4) {real, imag} */,
  {32'hbf621bb6, 32'h00000000} /* (4, 23, 3) {real, imag} */,
  {32'hbf585a7f, 32'h00000000} /* (4, 23, 2) {real, imag} */,
  {32'hbf93f722, 32'h00000000} /* (4, 23, 1) {real, imag} */,
  {32'hbf54e068, 32'h00000000} /* (4, 23, 0) {real, imag} */,
  {32'hbf10788b, 32'h00000000} /* (4, 22, 31) {real, imag} */,
  {32'hbfad0c9d, 32'h00000000} /* (4, 22, 30) {real, imag} */,
  {32'hbfa17fb1, 32'h00000000} /* (4, 22, 29) {real, imag} */,
  {32'hbf99acf0, 32'h00000000} /* (4, 22, 28) {real, imag} */,
  {32'hbf924572, 32'h00000000} /* (4, 22, 27) {real, imag} */,
  {32'hbf723610, 32'h00000000} /* (4, 22, 26) {real, imag} */,
  {32'hbf85d3ba, 32'h00000000} /* (4, 22, 25) {real, imag} */,
  {32'hbfb1849b, 32'h00000000} /* (4, 22, 24) {real, imag} */,
  {32'hbfac512c, 32'h00000000} /* (4, 22, 23) {real, imag} */,
  {32'hbf12b30b, 32'h00000000} /* (4, 22, 22) {real, imag} */,
  {32'hbe0a76b9, 32'h00000000} /* (4, 22, 21) {real, imag} */,
  {32'h3f8e4ce0, 32'h00000000} /* (4, 22, 20) {real, imag} */,
  {32'h3fa96602, 32'h00000000} /* (4, 22, 19) {real, imag} */,
  {32'h3fad9782, 32'h00000000} /* (4, 22, 18) {real, imag} */,
  {32'h3fabccd3, 32'h00000000} /* (4, 22, 17) {real, imag} */,
  {32'h3eebd216, 32'h00000000} /* (4, 22, 16) {real, imag} */,
  {32'h3f174f03, 32'h00000000} /* (4, 22, 15) {real, imag} */,
  {32'h3f91d3d6, 32'h00000000} /* (4, 22, 14) {real, imag} */,
  {32'h3f470a4b, 32'h00000000} /* (4, 22, 13) {real, imag} */,
  {32'h3ea6b3bd, 32'h00000000} /* (4, 22, 12) {real, imag} */,
  {32'h3e91e633, 32'h00000000} /* (4, 22, 11) {real, imag} */,
  {32'hbf4a2575, 32'h00000000} /* (4, 22, 10) {real, imag} */,
  {32'hbfad8a8f, 32'h00000000} /* (4, 22, 9) {real, imag} */,
  {32'hbf8f01b3, 32'h00000000} /* (4, 22, 8) {real, imag} */,
  {32'hbf5ded3f, 32'h00000000} /* (4, 22, 7) {real, imag} */,
  {32'hbf8ae083, 32'h00000000} /* (4, 22, 6) {real, imag} */,
  {32'hbf74934f, 32'h00000000} /* (4, 22, 5) {real, imag} */,
  {32'hbf32af5d, 32'h00000000} /* (4, 22, 4) {real, imag} */,
  {32'hbf5673cf, 32'h00000000} /* (4, 22, 3) {real, imag} */,
  {32'hbf11246b, 32'h00000000} /* (4, 22, 2) {real, imag} */,
  {32'hbf8a21ba, 32'h00000000} /* (4, 22, 1) {real, imag} */,
  {32'hbf2efc66, 32'h00000000} /* (4, 22, 0) {real, imag} */,
  {32'h3d0657f4, 32'h00000000} /* (4, 21, 31) {real, imag} */,
  {32'hbd303d0a, 32'h00000000} /* (4, 21, 30) {real, imag} */,
  {32'hbf023281, 32'h00000000} /* (4, 21, 29) {real, imag} */,
  {32'hbea4b643, 32'h00000000} /* (4, 21, 28) {real, imag} */,
  {32'hbec53bea, 32'h00000000} /* (4, 21, 27) {real, imag} */,
  {32'hbf7f017d, 32'h00000000} /* (4, 21, 26) {real, imag} */,
  {32'hbcc11a20, 32'h00000000} /* (4, 21, 25) {real, imag} */,
  {32'hbd519c83, 32'h00000000} /* (4, 21, 24) {real, imag} */,
  {32'hbedd1ffc, 32'h00000000} /* (4, 21, 23) {real, imag} */,
  {32'hbe4cf3a5, 32'h00000000} /* (4, 21, 22) {real, imag} */,
  {32'hbd8e9fc8, 32'h00000000} /* (4, 21, 21) {real, imag} */,
  {32'h3ebdb3cb, 32'h00000000} /* (4, 21, 20) {real, imag} */,
  {32'h3f5f3906, 32'h00000000} /* (4, 21, 19) {real, imag} */,
  {32'h3f070a01, 32'h00000000} /* (4, 21, 18) {real, imag} */,
  {32'h3edc2577, 32'h00000000} /* (4, 21, 17) {real, imag} */,
  {32'hbdd52b27, 32'h00000000} /* (4, 21, 16) {real, imag} */,
  {32'h3e469bb2, 32'h00000000} /* (4, 21, 15) {real, imag} */,
  {32'h3f4dca89, 32'h00000000} /* (4, 21, 14) {real, imag} */,
  {32'h3eec6304, 32'h00000000} /* (4, 21, 13) {real, imag} */,
  {32'hbd5b0d5e, 32'h00000000} /* (4, 21, 12) {real, imag} */,
  {32'h3ea6e702, 32'h00000000} /* (4, 21, 11) {real, imag} */,
  {32'h3e6730ac, 32'h00000000} /* (4, 21, 10) {real, imag} */,
  {32'hbe7f1ccd, 32'h00000000} /* (4, 21, 9) {real, imag} */,
  {32'hbe58b0a3, 32'h00000000} /* (4, 21, 8) {real, imag} */,
  {32'hbeb17e41, 32'h00000000} /* (4, 21, 7) {real, imag} */,
  {32'hbf1bd285, 32'h00000000} /* (4, 21, 6) {real, imag} */,
  {32'hbe49d44e, 32'h00000000} /* (4, 21, 5) {real, imag} */,
  {32'hbeb67044, 32'h00000000} /* (4, 21, 4) {real, imag} */,
  {32'hbf1c6184, 32'h00000000} /* (4, 21, 3) {real, imag} */,
  {32'h3d914a24, 32'h00000000} /* (4, 21, 2) {real, imag} */,
  {32'hbe9f4b21, 32'h00000000} /* (4, 21, 1) {real, imag} */,
  {32'hbebc10ae, 32'h00000000} /* (4, 21, 0) {real, imag} */,
  {32'h3f817ea3, 32'h00000000} /* (4, 20, 31) {real, imag} */,
  {32'h3fd247e2, 32'h00000000} /* (4, 20, 30) {real, imag} */,
  {32'h3f82e1ea, 32'h00000000} /* (4, 20, 29) {real, imag} */,
  {32'h3fab4ed7, 32'h00000000} /* (4, 20, 28) {real, imag} */,
  {32'h3f7ad7b3, 32'h00000000} /* (4, 20, 27) {real, imag} */,
  {32'h3ed5f40d, 32'h00000000} /* (4, 20, 26) {real, imag} */,
  {32'h3fb47c0e, 32'h00000000} /* (4, 20, 25) {real, imag} */,
  {32'h3fc12535, 32'h00000000} /* (4, 20, 24) {real, imag} */,
  {32'h3fa591ab, 32'h00000000} /* (4, 20, 23) {real, imag} */,
  {32'h3efb6a2d, 32'h00000000} /* (4, 20, 22) {real, imag} */,
  {32'h3e6cb1bb, 32'h00000000} /* (4, 20, 21) {real, imag} */,
  {32'hbef67905, 32'h00000000} /* (4, 20, 20) {real, imag} */,
  {32'hbe75bb9f, 32'h00000000} /* (4, 20, 19) {real, imag} */,
  {32'hbee1c670, 32'h00000000} /* (4, 20, 18) {real, imag} */,
  {32'hbf4e4fc0, 32'h00000000} /* (4, 20, 17) {real, imag} */,
  {32'hbf3ddb68, 32'h00000000} /* (4, 20, 16) {real, imag} */,
  {32'hbedad388, 32'h00000000} /* (4, 20, 15) {real, imag} */,
  {32'hbecbf85e, 32'h00000000} /* (4, 20, 14) {real, imag} */,
  {32'hbf2712ab, 32'h00000000} /* (4, 20, 13) {real, imag} */,
  {32'hbf56c01c, 32'h00000000} /* (4, 20, 12) {real, imag} */,
  {32'h3e0b7c6e, 32'h00000000} /* (4, 20, 11) {real, imag} */,
  {32'h3f94715e, 32'h00000000} /* (4, 20, 10) {real, imag} */,
  {32'h3f2bf76d, 32'h00000000} /* (4, 20, 9) {real, imag} */,
  {32'h3ea19fbf, 32'h00000000} /* (4, 20, 8) {real, imag} */,
  {32'h3f0a03eb, 32'h00000000} /* (4, 20, 7) {real, imag} */,
  {32'h3f35d44a, 32'h00000000} /* (4, 20, 6) {real, imag} */,
  {32'h3f92e618, 32'h00000000} /* (4, 20, 5) {real, imag} */,
  {32'h3f094308, 32'h00000000} /* (4, 20, 4) {real, imag} */,
  {32'h3e243d3d, 32'h00000000} /* (4, 20, 3) {real, imag} */,
  {32'h3f397d1b, 32'h00000000} /* (4, 20, 2) {real, imag} */,
  {32'h3f14bd02, 32'h00000000} /* (4, 20, 1) {real, imag} */,
  {32'h3e27868a, 32'h00000000} /* (4, 20, 0) {real, imag} */,
  {32'h3f372953, 32'h00000000} /* (4, 19, 31) {real, imag} */,
  {32'h3fb20002, 32'h00000000} /* (4, 19, 30) {real, imag} */,
  {32'h3f4a09a4, 32'h00000000} /* (4, 19, 29) {real, imag} */,
  {32'h3f92b3f9, 32'h00000000} /* (4, 19, 28) {real, imag} */,
  {32'h3f334142, 32'h00000000} /* (4, 19, 27) {real, imag} */,
  {32'h3f0e49e7, 32'h00000000} /* (4, 19, 26) {real, imag} */,
  {32'h3f84a34c, 32'h00000000} /* (4, 19, 25) {real, imag} */,
  {32'h3f8ed981, 32'h00000000} /* (4, 19, 24) {real, imag} */,
  {32'h3f56220a, 32'h00000000} /* (4, 19, 23) {real, imag} */,
  {32'h3f20aa15, 32'h00000000} /* (4, 19, 22) {real, imag} */,
  {32'h3e338f17, 32'h00000000} /* (4, 19, 21) {real, imag} */,
  {32'hbf6af24e, 32'h00000000} /* (4, 19, 20) {real, imag} */,
  {32'hbf797ba3, 32'h00000000} /* (4, 19, 19) {real, imag} */,
  {32'hbf60dae4, 32'h00000000} /* (4, 19, 18) {real, imag} */,
  {32'hbfc1bb0f, 32'h00000000} /* (4, 19, 17) {real, imag} */,
  {32'hbf8076f8, 32'h00000000} /* (4, 19, 16) {real, imag} */,
  {32'hbf65de6d, 32'h00000000} /* (4, 19, 15) {real, imag} */,
  {32'hbf3735da, 32'h00000000} /* (4, 19, 14) {real, imag} */,
  {32'hbf38512e, 32'h00000000} /* (4, 19, 13) {real, imag} */,
  {32'hbf56d919, 32'h00000000} /* (4, 19, 12) {real, imag} */,
  {32'hbf0aa479, 32'h00000000} /* (4, 19, 11) {real, imag} */,
  {32'h3f273517, 32'h00000000} /* (4, 19, 10) {real, imag} */,
  {32'h3f543a6c, 32'h00000000} /* (4, 19, 9) {real, imag} */,
  {32'h3ee62993, 32'h00000000} /* (4, 19, 8) {real, imag} */,
  {32'h3f530170, 32'h00000000} /* (4, 19, 7) {real, imag} */,
  {32'h3f351041, 32'h00000000} /* (4, 19, 6) {real, imag} */,
  {32'h3f991a55, 32'h00000000} /* (4, 19, 5) {real, imag} */,
  {32'h3f96fc97, 32'h00000000} /* (4, 19, 4) {real, imag} */,
  {32'h3f2c5942, 32'h00000000} /* (4, 19, 3) {real, imag} */,
  {32'h3e5c148b, 32'h00000000} /* (4, 19, 2) {real, imag} */,
  {32'h3f1277b1, 32'h00000000} /* (4, 19, 1) {real, imag} */,
  {32'h3eddfd4f, 32'h00000000} /* (4, 19, 0) {real, imag} */,
  {32'h3f142e64, 32'h00000000} /* (4, 18, 31) {real, imag} */,
  {32'h3f8276a7, 32'h00000000} /* (4, 18, 30) {real, imag} */,
  {32'h3f42c218, 32'h00000000} /* (4, 18, 29) {real, imag} */,
  {32'h3f5a974c, 32'h00000000} /* (4, 18, 28) {real, imag} */,
  {32'h3ea77abf, 32'h00000000} /* (4, 18, 27) {real, imag} */,
  {32'h3ed2c694, 32'h00000000} /* (4, 18, 26) {real, imag} */,
  {32'h3ef80d5f, 32'h00000000} /* (4, 18, 25) {real, imag} */,
  {32'h3f467be0, 32'h00000000} /* (4, 18, 24) {real, imag} */,
  {32'h3f251752, 32'h00000000} /* (4, 18, 23) {real, imag} */,
  {32'h3f340c6e, 32'h00000000} /* (4, 18, 22) {real, imag} */,
  {32'h3f212089, 32'h00000000} /* (4, 18, 21) {real, imag} */,
  {32'hbf394ca8, 32'h00000000} /* (4, 18, 20) {real, imag} */,
  {32'hbf506a6a, 32'h00000000} /* (4, 18, 19) {real, imag} */,
  {32'hbec9e4a3, 32'h00000000} /* (4, 18, 18) {real, imag} */,
  {32'hbf55f85a, 32'h00000000} /* (4, 18, 17) {real, imag} */,
  {32'hbf42c575, 32'h00000000} /* (4, 18, 16) {real, imag} */,
  {32'hbf79ff42, 32'h00000000} /* (4, 18, 15) {real, imag} */,
  {32'hbf7660f8, 32'h00000000} /* (4, 18, 14) {real, imag} */,
  {32'hbf847b4d, 32'h00000000} /* (4, 18, 13) {real, imag} */,
  {32'hbf44e8eb, 32'h00000000} /* (4, 18, 12) {real, imag} */,
  {32'hbf79cfc6, 32'h00000000} /* (4, 18, 11) {real, imag} */,
  {32'h3e5ac122, 32'h00000000} /* (4, 18, 10) {real, imag} */,
  {32'h3f663207, 32'h00000000} /* (4, 18, 9) {real, imag} */,
  {32'h3f3528e0, 32'h00000000} /* (4, 18, 8) {real, imag} */,
  {32'h3f58bb50, 32'h00000000} /* (4, 18, 7) {real, imag} */,
  {32'h3f9ae613, 32'h00000000} /* (4, 18, 6) {real, imag} */,
  {32'h3fc98d53, 32'h00000000} /* (4, 18, 5) {real, imag} */,
  {32'h3fb69ad7, 32'h00000000} /* (4, 18, 4) {real, imag} */,
  {32'h3f51b3b2, 32'h00000000} /* (4, 18, 3) {real, imag} */,
  {32'h3ee9e325, 32'h00000000} /* (4, 18, 2) {real, imag} */,
  {32'h3f504d75, 32'h00000000} /* (4, 18, 1) {real, imag} */,
  {32'h3ebe9bba, 32'h00000000} /* (4, 18, 0) {real, imag} */,
  {32'h3f08a171, 32'h00000000} /* (4, 17, 31) {real, imag} */,
  {32'h3f7a785e, 32'h00000000} /* (4, 17, 30) {real, imag} */,
  {32'h3f33b565, 32'h00000000} /* (4, 17, 29) {real, imag} */,
  {32'h3f1cbe88, 32'h00000000} /* (4, 17, 28) {real, imag} */,
  {32'h3f3fb599, 32'h00000000} /* (4, 17, 27) {real, imag} */,
  {32'h3f72b415, 32'h00000000} /* (4, 17, 26) {real, imag} */,
  {32'h3f1f9784, 32'h00000000} /* (4, 17, 25) {real, imag} */,
  {32'h3efb7b96, 32'h00000000} /* (4, 17, 24) {real, imag} */,
  {32'h3f3aa056, 32'h00000000} /* (4, 17, 23) {real, imag} */,
  {32'h3f28c705, 32'h00000000} /* (4, 17, 22) {real, imag} */,
  {32'h3ebf44a4, 32'h00000000} /* (4, 17, 21) {real, imag} */,
  {32'hbf3b5f3d, 32'h00000000} /* (4, 17, 20) {real, imag} */,
  {32'hbf79f838, 32'h00000000} /* (4, 17, 19) {real, imag} */,
  {32'hbee33bf3, 32'h00000000} /* (4, 17, 18) {real, imag} */,
  {32'hbf226dc9, 32'h00000000} /* (4, 17, 17) {real, imag} */,
  {32'hbf84f3b0, 32'h00000000} /* (4, 17, 16) {real, imag} */,
  {32'hbf8efb3b, 32'h00000000} /* (4, 17, 15) {real, imag} */,
  {32'hbf241fa9, 32'h00000000} /* (4, 17, 14) {real, imag} */,
  {32'hbf3c8fed, 32'h00000000} /* (4, 17, 13) {real, imag} */,
  {32'hbf441cc6, 32'h00000000} /* (4, 17, 12) {real, imag} */,
  {32'hbf68d83f, 32'h00000000} /* (4, 17, 11) {real, imag} */,
  {32'h3f1fde4d, 32'h00000000} /* (4, 17, 10) {real, imag} */,
  {32'h3f507730, 32'h00000000} /* (4, 17, 9) {real, imag} */,
  {32'h3f243c53, 32'h00000000} /* (4, 17, 8) {real, imag} */,
  {32'h3f2a29f1, 32'h00000000} /* (4, 17, 7) {real, imag} */,
  {32'h3f763045, 32'h00000000} /* (4, 17, 6) {real, imag} */,
  {32'h3fe24614, 32'h00000000} /* (4, 17, 5) {real, imag} */,
  {32'h3fcd8279, 32'h00000000} /* (4, 17, 4) {real, imag} */,
  {32'h3fab665f, 32'h00000000} /* (4, 17, 3) {real, imag} */,
  {32'h3f94b4f7, 32'h00000000} /* (4, 17, 2) {real, imag} */,
  {32'h3f585e15, 32'h00000000} /* (4, 17, 1) {real, imag} */,
  {32'h3e96060f, 32'h00000000} /* (4, 17, 0) {real, imag} */,
  {32'h3ed3bb56, 32'h00000000} /* (4, 16, 31) {real, imag} */,
  {32'h3f5cf7a0, 32'h00000000} /* (4, 16, 30) {real, imag} */,
  {32'h3f6b10e0, 32'h00000000} /* (4, 16, 29) {real, imag} */,
  {32'h3f0b455e, 32'h00000000} /* (4, 16, 28) {real, imag} */,
  {32'h3f5198ad, 32'h00000000} /* (4, 16, 27) {real, imag} */,
  {32'h3f8f299f, 32'h00000000} /* (4, 16, 26) {real, imag} */,
  {32'h3f889fba, 32'h00000000} /* (4, 16, 25) {real, imag} */,
  {32'h3f11f2e4, 32'h00000000} /* (4, 16, 24) {real, imag} */,
  {32'h3f799828, 32'h00000000} /* (4, 16, 23) {real, imag} */,
  {32'h3f669ef8, 32'h00000000} /* (4, 16, 22) {real, imag} */,
  {32'h3f17d4e7, 32'h00000000} /* (4, 16, 21) {real, imag} */,
  {32'hbf1c84f7, 32'h00000000} /* (4, 16, 20) {real, imag} */,
  {32'hbf93587b, 32'h00000000} /* (4, 16, 19) {real, imag} */,
  {32'hbf5cf2e3, 32'h00000000} /* (4, 16, 18) {real, imag} */,
  {32'hbf44e0f4, 32'h00000000} /* (4, 16, 17) {real, imag} */,
  {32'hbfaf1d1c, 32'h00000000} /* (4, 16, 16) {real, imag} */,
  {32'hbfb44db2, 32'h00000000} /* (4, 16, 15) {real, imag} */,
  {32'hbee92da8, 32'h00000000} /* (4, 16, 14) {real, imag} */,
  {32'hbf5197c5, 32'h00000000} /* (4, 16, 13) {real, imag} */,
  {32'hbf99828d, 32'h00000000} /* (4, 16, 12) {real, imag} */,
  {32'hbf8b4b42, 32'h00000000} /* (4, 16, 11) {real, imag} */,
  {32'h3e5c2c45, 32'h00000000} /* (4, 16, 10) {real, imag} */,
  {32'h3f3ddbd5, 32'h00000000} /* (4, 16, 9) {real, imag} */,
  {32'h3f8cf1ed, 32'h00000000} /* (4, 16, 8) {real, imag} */,
  {32'h3f89c3ea, 32'h00000000} /* (4, 16, 7) {real, imag} */,
  {32'h3f3183cc, 32'h00000000} /* (4, 16, 6) {real, imag} */,
  {32'h3f86c5b7, 32'h00000000} /* (4, 16, 5) {real, imag} */,
  {32'h3f86b7da, 32'h00000000} /* (4, 16, 4) {real, imag} */,
  {32'h3f885aff, 32'h00000000} /* (4, 16, 3) {real, imag} */,
  {32'h3f8b5cc8, 32'h00000000} /* (4, 16, 2) {real, imag} */,
  {32'h3f5eb172, 32'h00000000} /* (4, 16, 1) {real, imag} */,
  {32'h3f3b61b4, 32'h00000000} /* (4, 16, 0) {real, imag} */,
  {32'h3ecfd52d, 32'h00000000} /* (4, 15, 31) {real, imag} */,
  {32'h3f87d010, 32'h00000000} /* (4, 15, 30) {real, imag} */,
  {32'h3fa4a1a4, 32'h00000000} /* (4, 15, 29) {real, imag} */,
  {32'h3f982597, 32'h00000000} /* (4, 15, 28) {real, imag} */,
  {32'h3f914c04, 32'h00000000} /* (4, 15, 27) {real, imag} */,
  {32'h3f844221, 32'h00000000} /* (4, 15, 26) {real, imag} */,
  {32'h3f758082, 32'h00000000} /* (4, 15, 25) {real, imag} */,
  {32'h3f4eb2bd, 32'h00000000} /* (4, 15, 24) {real, imag} */,
  {32'h3fb6310a, 32'h00000000} /* (4, 15, 23) {real, imag} */,
  {32'h3fae04fb, 32'h00000000} /* (4, 15, 22) {real, imag} */,
  {32'h3f2e8887, 32'h00000000} /* (4, 15, 21) {real, imag} */,
  {32'hbf16e6f4, 32'h00000000} /* (4, 15, 20) {real, imag} */,
  {32'hbf21cd09, 32'h00000000} /* (4, 15, 19) {real, imag} */,
  {32'hbf186052, 32'h00000000} /* (4, 15, 18) {real, imag} */,
  {32'hbf0eb868, 32'h00000000} /* (4, 15, 17) {real, imag} */,
  {32'hbf016642, 32'h00000000} /* (4, 15, 16) {real, imag} */,
  {32'hbf90e114, 32'h00000000} /* (4, 15, 15) {real, imag} */,
  {32'hbf6f9da5, 32'h00000000} /* (4, 15, 14) {real, imag} */,
  {32'hbfd43299, 32'h00000000} /* (4, 15, 13) {real, imag} */,
  {32'hbfaae329, 32'h00000000} /* (4, 15, 12) {real, imag} */,
  {32'hbf203a0d, 32'h00000000} /* (4, 15, 11) {real, imag} */,
  {32'h3ef0b6a3, 32'h00000000} /* (4, 15, 10) {real, imag} */,
  {32'h3f7d246d, 32'h00000000} /* (4, 15, 9) {real, imag} */,
  {32'h3f69c276, 32'h00000000} /* (4, 15, 8) {real, imag} */,
  {32'h3f48ee1b, 32'h00000000} /* (4, 15, 7) {real, imag} */,
  {32'h3ed940fd, 32'h00000000} /* (4, 15, 6) {real, imag} */,
  {32'h3eccf012, 32'h00000000} /* (4, 15, 5) {real, imag} */,
  {32'h3efb7f0c, 32'h00000000} /* (4, 15, 4) {real, imag} */,
  {32'h3f080c8f, 32'h00000000} /* (4, 15, 3) {real, imag} */,
  {32'h3f1f44ae, 32'h00000000} /* (4, 15, 2) {real, imag} */,
  {32'h3f8f5019, 32'h00000000} /* (4, 15, 1) {real, imag} */,
  {32'h3f45d47a, 32'h00000000} /* (4, 15, 0) {real, imag} */,
  {32'h3f4a4ddf, 32'h00000000} /* (4, 14, 31) {real, imag} */,
  {32'h3f3fe13b, 32'h00000000} /* (4, 14, 30) {real, imag} */,
  {32'h3f8114a0, 32'h00000000} /* (4, 14, 29) {real, imag} */,
  {32'h3fbc1bcd, 32'h00000000} /* (4, 14, 28) {real, imag} */,
  {32'h3f98572a, 32'h00000000} /* (4, 14, 27) {real, imag} */,
  {32'h3f5d0128, 32'h00000000} /* (4, 14, 26) {real, imag} */,
  {32'h3efcd276, 32'h00000000} /* (4, 14, 25) {real, imag} */,
  {32'h3eb12a5b, 32'h00000000} /* (4, 14, 24) {real, imag} */,
  {32'h3f3f5d79, 32'h00000000} /* (4, 14, 23) {real, imag} */,
  {32'h3f9b602c, 32'h00000000} /* (4, 14, 22) {real, imag} */,
  {32'h3f3053cf, 32'h00000000} /* (4, 14, 21) {real, imag} */,
  {32'hbf38b4ae, 32'h00000000} /* (4, 14, 20) {real, imag} */,
  {32'hbf14a4f0, 32'h00000000} /* (4, 14, 19) {real, imag} */,
  {32'hbf066868, 32'h00000000} /* (4, 14, 18) {real, imag} */,
  {32'hbf7e775b, 32'h00000000} /* (4, 14, 17) {real, imag} */,
  {32'hbf308b16, 32'h00000000} /* (4, 14, 16) {real, imag} */,
  {32'hbf7e5d48, 32'h00000000} /* (4, 14, 15) {real, imag} */,
  {32'hbf272d80, 32'h00000000} /* (4, 14, 14) {real, imag} */,
  {32'hbf717529, 32'h00000000} /* (4, 14, 13) {real, imag} */,
  {32'hbf1faaaa, 32'h00000000} /* (4, 14, 12) {real, imag} */,
  {32'hbe4a2ac1, 32'h00000000} /* (4, 14, 11) {real, imag} */,
  {32'h3f0a925e, 32'h00000000} /* (4, 14, 10) {real, imag} */,
  {32'h3f853697, 32'h00000000} /* (4, 14, 9) {real, imag} */,
  {32'h3f8e47b9, 32'h00000000} /* (4, 14, 8) {real, imag} */,
  {32'h3f9d9aab, 32'h00000000} /* (4, 14, 7) {real, imag} */,
  {32'h3f4f0a4b, 32'h00000000} /* (4, 14, 6) {real, imag} */,
  {32'h3f132637, 32'h00000000} /* (4, 14, 5) {real, imag} */,
  {32'h3ec982f5, 32'h00000000} /* (4, 14, 4) {real, imag} */,
  {32'h3e5bcb25, 32'h00000000} /* (4, 14, 3) {real, imag} */,
  {32'h3e75678c, 32'h00000000} /* (4, 14, 2) {real, imag} */,
  {32'h3f92c4d4, 32'h00000000} /* (4, 14, 1) {real, imag} */,
  {32'h3f6a3461, 32'h00000000} /* (4, 14, 0) {real, imag} */,
  {32'h3ee9c94c, 32'h00000000} /* (4, 13, 31) {real, imag} */,
  {32'h3ed210c1, 32'h00000000} /* (4, 13, 30) {real, imag} */,
  {32'h3f5d0d66, 32'h00000000} /* (4, 13, 29) {real, imag} */,
  {32'h3f9b0817, 32'h00000000} /* (4, 13, 28) {real, imag} */,
  {32'h3fa36257, 32'h00000000} /* (4, 13, 27) {real, imag} */,
  {32'h3f87320e, 32'h00000000} /* (4, 13, 26) {real, imag} */,
  {32'h3f058a59, 32'h00000000} /* (4, 13, 25) {real, imag} */,
  {32'h3ed04c74, 32'h00000000} /* (4, 13, 24) {real, imag} */,
  {32'h3eedb520, 32'h00000000} /* (4, 13, 23) {real, imag} */,
  {32'h3fa832f2, 32'h00000000} /* (4, 13, 22) {real, imag} */,
  {32'h3f7fe1ad, 32'h00000000} /* (4, 13, 21) {real, imag} */,
  {32'hbf86e6fb, 32'h00000000} /* (4, 13, 20) {real, imag} */,
  {32'hbfb0c7ea, 32'h00000000} /* (4, 13, 19) {real, imag} */,
  {32'hbf62576b, 32'h00000000} /* (4, 13, 18) {real, imag} */,
  {32'hbfa12052, 32'h00000000} /* (4, 13, 17) {real, imag} */,
  {32'hbf3c264b, 32'h00000000} /* (4, 13, 16) {real, imag} */,
  {32'hbee3f303, 32'h00000000} /* (4, 13, 15) {real, imag} */,
  {32'hbf1f8130, 32'h00000000} /* (4, 13, 14) {real, imag} */,
  {32'hbf47c124, 32'h00000000} /* (4, 13, 13) {real, imag} */,
  {32'hbedaf90b, 32'h00000000} /* (4, 13, 12) {real, imag} */,
  {32'hbe1e0bfd, 32'h00000000} /* (4, 13, 11) {real, imag} */,
  {32'h3f1a0eaa, 32'h00000000} /* (4, 13, 10) {real, imag} */,
  {32'h3f1b356f, 32'h00000000} /* (4, 13, 9) {real, imag} */,
  {32'h3f05909c, 32'h00000000} /* (4, 13, 8) {real, imag} */,
  {32'h3f56f514, 32'h00000000} /* (4, 13, 7) {real, imag} */,
  {32'h3f325737, 32'h00000000} /* (4, 13, 6) {real, imag} */,
  {32'h3eeb55cb, 32'h00000000} /* (4, 13, 5) {real, imag} */,
  {32'h3e9a540c, 32'h00000000} /* (4, 13, 4) {real, imag} */,
  {32'h3ed77340, 32'h00000000} /* (4, 13, 3) {real, imag} */,
  {32'h3f839670, 32'h00000000} /* (4, 13, 2) {real, imag} */,
  {32'h3fb1717a, 32'h00000000} /* (4, 13, 1) {real, imag} */,
  {32'h3f8558ef, 32'h00000000} /* (4, 13, 0) {real, imag} */,
  {32'h3db74475, 32'h00000000} /* (4, 12, 31) {real, imag} */,
  {32'h3eff04d6, 32'h00000000} /* (4, 12, 30) {real, imag} */,
  {32'h3f723535, 32'h00000000} /* (4, 12, 29) {real, imag} */,
  {32'h3f867c5f, 32'h00000000} /* (4, 12, 28) {real, imag} */,
  {32'h3f67981a, 32'h00000000} /* (4, 12, 27) {real, imag} */,
  {32'h3f1899df, 32'h00000000} /* (4, 12, 26) {real, imag} */,
  {32'h3f298c86, 32'h00000000} /* (4, 12, 25) {real, imag} */,
  {32'h3f7a28d0, 32'h00000000} /* (4, 12, 24) {real, imag} */,
  {32'h3f6485fc, 32'h00000000} /* (4, 12, 23) {real, imag} */,
  {32'h3fadcff3, 32'h00000000} /* (4, 12, 22) {real, imag} */,
  {32'h3f38e1b6, 32'h00000000} /* (4, 12, 21) {real, imag} */,
  {32'hbf40d88f, 32'h00000000} /* (4, 12, 20) {real, imag} */,
  {32'hbfa6cc50, 32'h00000000} /* (4, 12, 19) {real, imag} */,
  {32'hbf43e103, 32'h00000000} /* (4, 12, 18) {real, imag} */,
  {32'hbf4c64b8, 32'h00000000} /* (4, 12, 17) {real, imag} */,
  {32'hbf0c8e00, 32'h00000000} /* (4, 12, 16) {real, imag} */,
  {32'hbf06c241, 32'h00000000} /* (4, 12, 15) {real, imag} */,
  {32'hbf4f163c, 32'h00000000} /* (4, 12, 14) {real, imag} */,
  {32'hbf301cf5, 32'h00000000} /* (4, 12, 13) {real, imag} */,
  {32'hbe9a1161, 32'h00000000} /* (4, 12, 12) {real, imag} */,
  {32'h3d873a10, 32'h00000000} /* (4, 12, 11) {real, imag} */,
  {32'h3f895905, 32'h00000000} /* (4, 12, 10) {real, imag} */,
  {32'h3f42cd13, 32'h00000000} /* (4, 12, 9) {real, imag} */,
  {32'h3ebf3452, 32'h00000000} /* (4, 12, 8) {real, imag} */,
  {32'h3f3df672, 32'h00000000} /* (4, 12, 7) {real, imag} */,
  {32'h3f42fdb2, 32'h00000000} /* (4, 12, 6) {real, imag} */,
  {32'h3f1df1b7, 32'h00000000} /* (4, 12, 5) {real, imag} */,
  {32'h3f5745ea, 32'h00000000} /* (4, 12, 4) {real, imag} */,
  {32'h3f45fbf7, 32'h00000000} /* (4, 12, 3) {real, imag} */,
  {32'h3f8c70c4, 32'h00000000} /* (4, 12, 2) {real, imag} */,
  {32'h3fa72b34, 32'h00000000} /* (4, 12, 1) {real, imag} */,
  {32'h3f376872, 32'h00000000} /* (4, 12, 0) {real, imag} */,
  {32'h3e6aa43d, 32'h00000000} /* (4, 11, 31) {real, imag} */,
  {32'h3f27d5a6, 32'h00000000} /* (4, 11, 30) {real, imag} */,
  {32'h3f1d697b, 32'h00000000} /* (4, 11, 29) {real, imag} */,
  {32'h3f80f8aa, 32'h00000000} /* (4, 11, 28) {real, imag} */,
  {32'h3f544569, 32'h00000000} /* (4, 11, 27) {real, imag} */,
  {32'h3f18e741, 32'h00000000} /* (4, 11, 26) {real, imag} */,
  {32'h3efe84aa, 32'h00000000} /* (4, 11, 25) {real, imag} */,
  {32'h3efb7c04, 32'h00000000} /* (4, 11, 24) {real, imag} */,
  {32'h3f5e1cd4, 32'h00000000} /* (4, 11, 23) {real, imag} */,
  {32'h3f98f85e, 32'h00000000} /* (4, 11, 22) {real, imag} */,
  {32'h3ef8e10b, 32'h00000000} /* (4, 11, 21) {real, imag} */,
  {32'hbe6426a9, 32'h00000000} /* (4, 11, 20) {real, imag} */,
  {32'hbf68f9e2, 32'h00000000} /* (4, 11, 19) {real, imag} */,
  {32'hbf92765f, 32'h00000000} /* (4, 11, 18) {real, imag} */,
  {32'hbf43ff55, 32'h00000000} /* (4, 11, 17) {real, imag} */,
  {32'hbe93085d, 32'h00000000} /* (4, 11, 16) {real, imag} */,
  {32'hbf332591, 32'h00000000} /* (4, 11, 15) {real, imag} */,
  {32'hbf60dd10, 32'h00000000} /* (4, 11, 14) {real, imag} */,
  {32'hbf6a9e60, 32'h00000000} /* (4, 11, 13) {real, imag} */,
  {32'hbf0547b1, 32'h00000000} /* (4, 11, 12) {real, imag} */,
  {32'hbb35d9de, 32'h00000000} /* (4, 11, 11) {real, imag} */,
  {32'h3f9bca3a, 32'h00000000} /* (4, 11, 10) {real, imag} */,
  {32'h3f58f21f, 32'h00000000} /* (4, 11, 9) {real, imag} */,
  {32'h3e8cfce8, 32'h00000000} /* (4, 11, 8) {real, imag} */,
  {32'h3f10876d, 32'h00000000} /* (4, 11, 7) {real, imag} */,
  {32'h3f2dc644, 32'h00000000} /* (4, 11, 6) {real, imag} */,
  {32'h3f315e5c, 32'h00000000} /* (4, 11, 5) {real, imag} */,
  {32'h3f1ee646, 32'h00000000} /* (4, 11, 4) {real, imag} */,
  {32'h3f11e1be, 32'h00000000} /* (4, 11, 3) {real, imag} */,
  {32'h3f0316c1, 32'h00000000} /* (4, 11, 2) {real, imag} */,
  {32'h3f8b0020, 32'h00000000} /* (4, 11, 1) {real, imag} */,
  {32'h3f1620a2, 32'h00000000} /* (4, 11, 0) {real, imag} */,
  {32'hbdb1fcaa, 32'h00000000} /* (4, 10, 31) {real, imag} */,
  {32'hbcd7ab72, 32'h00000000} /* (4, 10, 30) {real, imag} */,
  {32'hbeb6b83a, 32'h00000000} /* (4, 10, 29) {real, imag} */,
  {32'hbf027ecb, 32'h00000000} /* (4, 10, 28) {real, imag} */,
  {32'hbf0677a1, 32'h00000000} /* (4, 10, 27) {real, imag} */,
  {32'hbec76313, 32'h00000000} /* (4, 10, 26) {real, imag} */,
  {32'hbee0f0e7, 32'h00000000} /* (4, 10, 25) {real, imag} */,
  {32'hbf2ce950, 32'h00000000} /* (4, 10, 24) {real, imag} */,
  {32'hbf26e28d, 32'h00000000} /* (4, 10, 23) {real, imag} */,
  {32'hbea75b8b, 32'h00000000} /* (4, 10, 22) {real, imag} */,
  {32'hbf1b05e3, 32'h00000000} /* (4, 10, 21) {real, imag} */,
  {32'h3ebda763, 32'h00000000} /* (4, 10, 20) {real, imag} */,
  {32'h3f0d1118, 32'h00000000} /* (4, 10, 19) {real, imag} */,
  {32'hbef2c57c, 32'h00000000} /* (4, 10, 18) {real, imag} */,
  {32'hbdb5d65f, 32'h00000000} /* (4, 10, 17) {real, imag} */,
  {32'h3f16bf1a, 32'h00000000} /* (4, 10, 16) {real, imag} */,
  {32'h3e97ef38, 32'h00000000} /* (4, 10, 15) {real, imag} */,
  {32'hbdb9e189, 32'h00000000} /* (4, 10, 14) {real, imag} */,
  {32'hbe3ea714, 32'h00000000} /* (4, 10, 13) {real, imag} */,
  {32'h3ef05e01, 32'h00000000} /* (4, 10, 12) {real, imag} */,
  {32'h3f594e8a, 32'h00000000} /* (4, 10, 11) {real, imag} */,
  {32'h3a3b9b04, 32'h00000000} /* (4, 10, 10) {real, imag} */,
  {32'hbf233cd4, 32'h00000000} /* (4, 10, 9) {real, imag} */,
  {32'hbf431714, 32'h00000000} /* (4, 10, 8) {real, imag} */,
  {32'hbf33a346, 32'h00000000} /* (4, 10, 7) {real, imag} */,
  {32'hbece42fc, 32'h00000000} /* (4, 10, 6) {real, imag} */,
  {32'hbe0369d4, 32'h00000000} /* (4, 10, 5) {real, imag} */,
  {32'hbf00bfed, 32'h00000000} /* (4, 10, 4) {real, imag} */,
  {32'hbf12e1dd, 32'h00000000} /* (4, 10, 3) {real, imag} */,
  {32'hbf126f26, 32'h00000000} /* (4, 10, 2) {real, imag} */,
  {32'hbd3cbc1a, 32'h00000000} /* (4, 10, 1) {real, imag} */,
  {32'hbe859e7e, 32'h00000000} /* (4, 10, 0) {real, imag} */,
  {32'hbea605cb, 32'h00000000} /* (4, 9, 31) {real, imag} */,
  {32'hbf60450c, 32'h00000000} /* (4, 9, 30) {real, imag} */,
  {32'hbf8d6329, 32'h00000000} /* (4, 9, 29) {real, imag} */,
  {32'hbf8df061, 32'h00000000} /* (4, 9, 28) {real, imag} */,
  {32'hbf56b46d, 32'h00000000} /* (4, 9, 27) {real, imag} */,
  {32'hbf2cbd11, 32'h00000000} /* (4, 9, 26) {real, imag} */,
  {32'hbefd566d, 32'h00000000} /* (4, 9, 25) {real, imag} */,
  {32'hbf512e97, 32'h00000000} /* (4, 9, 24) {real, imag} */,
  {32'hbf90f9d6, 32'h00000000} /* (4, 9, 23) {real, imag} */,
  {32'hbf696e93, 32'h00000000} /* (4, 9, 22) {real, imag} */,
  {32'hbf2a1e94, 32'h00000000} /* (4, 9, 21) {real, imag} */,
  {32'h3f457624, 32'h00000000} /* (4, 9, 20) {real, imag} */,
  {32'h3f6884cc, 32'h00000000} /* (4, 9, 19) {real, imag} */,
  {32'h3f3eec89, 32'h00000000} /* (4, 9, 18) {real, imag} */,
  {32'h3f33c0f6, 32'h00000000} /* (4, 9, 17) {real, imag} */,
  {32'h3f724650, 32'h00000000} /* (4, 9, 16) {real, imag} */,
  {32'h3f60b8b6, 32'h00000000} /* (4, 9, 15) {real, imag} */,
  {32'h3ec10d3c, 32'h00000000} /* (4, 9, 14) {real, imag} */,
  {32'h3ed573d0, 32'h00000000} /* (4, 9, 13) {real, imag} */,
  {32'h3fa3f070, 32'h00000000} /* (4, 9, 12) {real, imag} */,
  {32'h3f8efb72, 32'h00000000} /* (4, 9, 11) {real, imag} */,
  {32'hbe2aea12, 32'h00000000} /* (4, 9, 10) {real, imag} */,
  {32'hbf8e6fef, 32'h00000000} /* (4, 9, 9) {real, imag} */,
  {32'hbf9f475b, 32'h00000000} /* (4, 9, 8) {real, imag} */,
  {32'hbf32941f, 32'h00000000} /* (4, 9, 7) {real, imag} */,
  {32'hbefe06e7, 32'h00000000} /* (4, 9, 6) {real, imag} */,
  {32'hbf070cc5, 32'h00000000} /* (4, 9, 5) {real, imag} */,
  {32'hbf34d0a9, 32'h00000000} /* (4, 9, 4) {real, imag} */,
  {32'hbf547829, 32'h00000000} /* (4, 9, 3) {real, imag} */,
  {32'hbf928290, 32'h00000000} /* (4, 9, 2) {real, imag} */,
  {32'hbf1f4392, 32'h00000000} /* (4, 9, 1) {real, imag} */,
  {32'hbeb526d5, 32'h00000000} /* (4, 9, 0) {real, imag} */,
  {32'hbe405fc7, 32'h00000000} /* (4, 8, 31) {real, imag} */,
  {32'hbf2eb127, 32'h00000000} /* (4, 8, 30) {real, imag} */,
  {32'hbf6aec91, 32'h00000000} /* (4, 8, 29) {real, imag} */,
  {32'hbf926018, 32'h00000000} /* (4, 8, 28) {real, imag} */,
  {32'hbf7a7806, 32'h00000000} /* (4, 8, 27) {real, imag} */,
  {32'hbf957a36, 32'h00000000} /* (4, 8, 26) {real, imag} */,
  {32'hbf6549b0, 32'h00000000} /* (4, 8, 25) {real, imag} */,
  {32'hbf0eb4af, 32'h00000000} /* (4, 8, 24) {real, imag} */,
  {32'hbf043a4b, 32'h00000000} /* (4, 8, 23) {real, imag} */,
  {32'hbf26e4e8, 32'h00000000} /* (4, 8, 22) {real, imag} */,
  {32'hbdbf913e, 32'h00000000} /* (4, 8, 21) {real, imag} */,
  {32'h3f4d7778, 32'h00000000} /* (4, 8, 20) {real, imag} */,
  {32'h3f853fb8, 32'h00000000} /* (4, 8, 19) {real, imag} */,
  {32'h3fa32297, 32'h00000000} /* (4, 8, 18) {real, imag} */,
  {32'h3f7a86dd, 32'h00000000} /* (4, 8, 17) {real, imag} */,
  {32'h3f6e09a7, 32'h00000000} /* (4, 8, 16) {real, imag} */,
  {32'h3fa6b4d0, 32'h00000000} /* (4, 8, 15) {real, imag} */,
  {32'h3e9da007, 32'h00000000} /* (4, 8, 14) {real, imag} */,
  {32'h3e3e8922, 32'h00000000} /* (4, 8, 13) {real, imag} */,
  {32'h3f96b911, 32'h00000000} /* (4, 8, 12) {real, imag} */,
  {32'h3f2ac321, 32'h00000000} /* (4, 8, 11) {real, imag} */,
  {32'hbeda6999, 32'h00000000} /* (4, 8, 10) {real, imag} */,
  {32'hbf5a9432, 32'h00000000} /* (4, 8, 9) {real, imag} */,
  {32'hbf8c682e, 32'h00000000} /* (4, 8, 8) {real, imag} */,
  {32'hbeca63dc, 32'h00000000} /* (4, 8, 7) {real, imag} */,
  {32'hbf36b3df, 32'h00000000} /* (4, 8, 6) {real, imag} */,
  {32'hbf7c1bf3, 32'h00000000} /* (4, 8, 5) {real, imag} */,
  {32'hbf8ff70e, 32'h00000000} /* (4, 8, 4) {real, imag} */,
  {32'hbf4a67a4, 32'h00000000} /* (4, 8, 3) {real, imag} */,
  {32'hbf1bee02, 32'h00000000} /* (4, 8, 2) {real, imag} */,
  {32'hbf25db06, 32'h00000000} /* (4, 8, 1) {real, imag} */,
  {32'hbec18e00, 32'h00000000} /* (4, 8, 0) {real, imag} */,
  {32'hbd8d1ace, 32'h00000000} /* (4, 7, 31) {real, imag} */,
  {32'hbe9739a9, 32'h00000000} /* (4, 7, 30) {real, imag} */,
  {32'hbf17d2e1, 32'h00000000} /* (4, 7, 29) {real, imag} */,
  {32'hbf4be536, 32'h00000000} /* (4, 7, 28) {real, imag} */,
  {32'hbf7cd9e8, 32'h00000000} /* (4, 7, 27) {real, imag} */,
  {32'hbfc28bc9, 32'h00000000} /* (4, 7, 26) {real, imag} */,
  {32'hbf968c43, 32'h00000000} /* (4, 7, 25) {real, imag} */,
  {32'hbf81829c, 32'h00000000} /* (4, 7, 24) {real, imag} */,
  {32'hbe7bfd07, 32'h00000000} /* (4, 7, 23) {real, imag} */,
  {32'hbe905437, 32'h00000000} /* (4, 7, 22) {real, imag} */,
  {32'hbcae3791, 32'h00000000} /* (4, 7, 21) {real, imag} */,
  {32'h3f2b101b, 32'h00000000} /* (4, 7, 20) {real, imag} */,
  {32'h3f5a4f0a, 32'h00000000} /* (4, 7, 19) {real, imag} */,
  {32'h3f9ae964, 32'h00000000} /* (4, 7, 18) {real, imag} */,
  {32'h3fd17d0f, 32'h00000000} /* (4, 7, 17) {real, imag} */,
  {32'h3fa67004, 32'h00000000} /* (4, 7, 16) {real, imag} */,
  {32'h3fb35bff, 32'h00000000} /* (4, 7, 15) {real, imag} */,
  {32'h3f8d7e36, 32'h00000000} /* (4, 7, 14) {real, imag} */,
  {32'h3f110d44, 32'h00000000} /* (4, 7, 13) {real, imag} */,
  {32'h3f815d7a, 32'h00000000} /* (4, 7, 12) {real, imag} */,
  {32'h3f6adcb2, 32'h00000000} /* (4, 7, 11) {real, imag} */,
  {32'hbe6013a6, 32'h00000000} /* (4, 7, 10) {real, imag} */,
  {32'hbe011121, 32'h00000000} /* (4, 7, 9) {real, imag} */,
  {32'hbeacece9, 32'h00000000} /* (4, 7, 8) {real, imag} */,
  {32'hbe9b0fe1, 32'h00000000} /* (4, 7, 7) {real, imag} */,
  {32'hbf6de4e3, 32'h00000000} /* (4, 7, 6) {real, imag} */,
  {32'hbf8b63ac, 32'h00000000} /* (4, 7, 5) {real, imag} */,
  {32'hbfb277f1, 32'h00000000} /* (4, 7, 4) {real, imag} */,
  {32'hbf4d9f29, 32'h00000000} /* (4, 7, 3) {real, imag} */,
  {32'hbe39d50c, 32'h00000000} /* (4, 7, 2) {real, imag} */,
  {32'hbdcbc9c7, 32'h00000000} /* (4, 7, 1) {real, imag} */,
  {32'hbe105101, 32'h00000000} /* (4, 7, 0) {real, imag} */,
  {32'hbdd3db13, 32'h00000000} /* (4, 6, 31) {real, imag} */,
  {32'hbe593ee8, 32'h00000000} /* (4, 6, 30) {real, imag} */,
  {32'hbfb1f02c, 32'h00000000} /* (4, 6, 29) {real, imag} */,
  {32'hbf488cc8, 32'h00000000} /* (4, 6, 28) {real, imag} */,
  {32'hbf0ac3c7, 32'h00000000} /* (4, 6, 27) {real, imag} */,
  {32'hbf791f65, 32'h00000000} /* (4, 6, 26) {real, imag} */,
  {32'hbf574739, 32'h00000000} /* (4, 6, 25) {real, imag} */,
  {32'hbf3880c3, 32'h00000000} /* (4, 6, 24) {real, imag} */,
  {32'h3ccea4cb, 32'h00000000} /* (4, 6, 23) {real, imag} */,
  {32'h3d3ee425, 32'h00000000} /* (4, 6, 22) {real, imag} */,
  {32'hbe3f89b9, 32'h00000000} /* (4, 6, 21) {real, imag} */,
  {32'hbe19d453, 32'h00000000} /* (4, 6, 20) {real, imag} */,
  {32'h3e8f06de, 32'h00000000} /* (4, 6, 19) {real, imag} */,
  {32'h3f55077c, 32'h00000000} /* (4, 6, 18) {real, imag} */,
  {32'h3f98a2db, 32'h00000000} /* (4, 6, 17) {real, imag} */,
  {32'h3f76ed6a, 32'h00000000} /* (4, 6, 16) {real, imag} */,
  {32'h3f53e1d5, 32'h00000000} /* (4, 6, 15) {real, imag} */,
  {32'h3fa2a251, 32'h00000000} /* (4, 6, 14) {real, imag} */,
  {32'h3f701cd4, 32'h00000000} /* (4, 6, 13) {real, imag} */,
  {32'h3f45336a, 32'h00000000} /* (4, 6, 12) {real, imag} */,
  {32'h3f0ccf92, 32'h00000000} /* (4, 6, 11) {real, imag} */,
  {32'h3c8c942a, 32'h00000000} /* (4, 6, 10) {real, imag} */,
  {32'hbde9956b, 32'h00000000} /* (4, 6, 9) {real, imag} */,
  {32'hbec0310c, 32'h00000000} /* (4, 6, 8) {real, imag} */,
  {32'hbf020aa4, 32'h00000000} /* (4, 6, 7) {real, imag} */,
  {32'hbf9184cd, 32'h00000000} /* (4, 6, 6) {real, imag} */,
  {32'hbf19ec6e, 32'h00000000} /* (4, 6, 5) {real, imag} */,
  {32'hbf54abde, 32'h00000000} /* (4, 6, 4) {real, imag} */,
  {32'hbf4083b3, 32'h00000000} /* (4, 6, 3) {real, imag} */,
  {32'hbf161705, 32'h00000000} /* (4, 6, 2) {real, imag} */,
  {32'hbef5cef8, 32'h00000000} /* (4, 6, 1) {real, imag} */,
  {32'hbe9964a8, 32'h00000000} /* (4, 6, 0) {real, imag} */,
  {32'h3d01f658, 32'h00000000} /* (4, 5, 31) {real, imag} */,
  {32'hbe5ab08d, 32'h00000000} /* (4, 5, 30) {real, imag} */,
  {32'hbf9eca41, 32'h00000000} /* (4, 5, 29) {real, imag} */,
  {32'hbf7df4d4, 32'h00000000} /* (4, 5, 28) {real, imag} */,
  {32'hbf984bb7, 32'h00000000} /* (4, 5, 27) {real, imag} */,
  {32'hbfc414ea, 32'h00000000} /* (4, 5, 26) {real, imag} */,
  {32'hbfd451ad, 32'h00000000} /* (4, 5, 25) {real, imag} */,
  {32'hbfba3d62, 32'h00000000} /* (4, 5, 24) {real, imag} */,
  {32'hbf4bc1dd, 32'h00000000} /* (4, 5, 23) {real, imag} */,
  {32'hbeb68918, 32'h00000000} /* (4, 5, 22) {real, imag} */,
  {32'hbf2d958e, 32'h00000000} /* (4, 5, 21) {real, imag} */,
  {32'hbf7290bd, 32'h00000000} /* (4, 5, 20) {real, imag} */,
  {32'hbedd2b40, 32'h00000000} /* (4, 5, 19) {real, imag} */,
  {32'h3d739590, 32'h00000000} /* (4, 5, 18) {real, imag} */,
  {32'hbed1a8ec, 32'h00000000} /* (4, 5, 17) {real, imag} */,
  {32'hbe39072a, 32'h00000000} /* (4, 5, 16) {real, imag} */,
  {32'h3e7953cd, 32'h00000000} /* (4, 5, 15) {real, imag} */,
  {32'h3f6da383, 32'h00000000} /* (4, 5, 14) {real, imag} */,
  {32'h3f5ac5e6, 32'h00000000} /* (4, 5, 13) {real, imag} */,
  {32'h3f8ee8d4, 32'h00000000} /* (4, 5, 12) {real, imag} */,
  {32'h3ee96ddc, 32'h00000000} /* (4, 5, 11) {real, imag} */,
  {32'h3eabf5d2, 32'h00000000} /* (4, 5, 10) {real, imag} */,
  {32'h3e86c8e3, 32'h00000000} /* (4, 5, 9) {real, imag} */,
  {32'h3ec44310, 32'h00000000} /* (4, 5, 8) {real, imag} */,
  {32'h3f555229, 32'h00000000} /* (4, 5, 7) {real, imag} */,
  {32'h3e96b9c1, 32'h00000000} /* (4, 5, 6) {real, imag} */,
  {32'hbd42dcfd, 32'h00000000} /* (4, 5, 5) {real, imag} */,
  {32'hbf11c4bc, 32'h00000000} /* (4, 5, 4) {real, imag} */,
  {32'hbf24ee0f, 32'h00000000} /* (4, 5, 3) {real, imag} */,
  {32'hbf03cb0b, 32'h00000000} /* (4, 5, 2) {real, imag} */,
  {32'hbf245ad4, 32'h00000000} /* (4, 5, 1) {real, imag} */,
  {32'hbeb3f793, 32'h00000000} /* (4, 5, 0) {real, imag} */,
  {32'hbdffd43c, 32'h00000000} /* (4, 4, 31) {real, imag} */,
  {32'hbee3ceca, 32'h00000000} /* (4, 4, 30) {real, imag} */,
  {32'hbfb991e9, 32'h00000000} /* (4, 4, 29) {real, imag} */,
  {32'hbfeaf2fe, 32'h00000000} /* (4, 4, 28) {real, imag} */,
  {32'hbf89b6dd, 32'h00000000} /* (4, 4, 27) {real, imag} */,
  {32'hbf36173f, 32'h00000000} /* (4, 4, 26) {real, imag} */,
  {32'hbf8b0064, 32'h00000000} /* (4, 4, 25) {real, imag} */,
  {32'hbfe1d786, 32'h00000000} /* (4, 4, 24) {real, imag} */,
  {32'hbfb661de, 32'h00000000} /* (4, 4, 23) {real, imag} */,
  {32'hbf121fa0, 32'h00000000} /* (4, 4, 22) {real, imag} */,
  {32'hbf458777, 32'h00000000} /* (4, 4, 21) {real, imag} */,
  {32'hbf3c7d82, 32'h00000000} /* (4, 4, 20) {real, imag} */,
  {32'hbf69840a, 32'h00000000} /* (4, 4, 19) {real, imag} */,
  {32'hbf4c6ebf, 32'h00000000} /* (4, 4, 18) {real, imag} */,
  {32'hbf5090d8, 32'h00000000} /* (4, 4, 17) {real, imag} */,
  {32'hbf12ab8e, 32'h00000000} /* (4, 4, 16) {real, imag} */,
  {32'h3ec7d291, 32'h00000000} /* (4, 4, 15) {real, imag} */,
  {32'h3f894d76, 32'h00000000} /* (4, 4, 14) {real, imag} */,
  {32'h3f9d4152, 32'h00000000} /* (4, 4, 13) {real, imag} */,
  {32'h3f611dca, 32'h00000000} /* (4, 4, 12) {real, imag} */,
  {32'h3f201388, 32'h00000000} /* (4, 4, 11) {real, imag} */,
  {32'h3f183c4a, 32'h00000000} /* (4, 4, 10) {real, imag} */,
  {32'h3f0e9887, 32'h00000000} /* (4, 4, 9) {real, imag} */,
  {32'h3f78453d, 32'h00000000} /* (4, 4, 8) {real, imag} */,
  {32'h3f84b9a4, 32'h00000000} /* (4, 4, 7) {real, imag} */,
  {32'h3f9ace40, 32'h00000000} /* (4, 4, 6) {real, imag} */,
  {32'h3ea3b72e, 32'h00000000} /* (4, 4, 5) {real, imag} */,
  {32'hbf5f24e3, 32'h00000000} /* (4, 4, 4) {real, imag} */,
  {32'hbf9da2d4, 32'h00000000} /* (4, 4, 3) {real, imag} */,
  {32'hbf7030e8, 32'h00000000} /* (4, 4, 2) {real, imag} */,
  {32'hbf6c6193, 32'h00000000} /* (4, 4, 1) {real, imag} */,
  {32'hbee80387, 32'h00000000} /* (4, 4, 0) {real, imag} */,
  {32'hbecb5a32, 32'h00000000} /* (4, 3, 31) {real, imag} */,
  {32'hbf3b2341, 32'h00000000} /* (4, 3, 30) {real, imag} */,
  {32'hbfa48716, 32'h00000000} /* (4, 3, 29) {real, imag} */,
  {32'hbfc399ca, 32'h00000000} /* (4, 3, 28) {real, imag} */,
  {32'hbf0cc35e, 32'h00000000} /* (4, 3, 27) {real, imag} */,
  {32'hbe806154, 32'h00000000} /* (4, 3, 26) {real, imag} */,
  {32'hbef148f3, 32'h00000000} /* (4, 3, 25) {real, imag} */,
  {32'hbf7f6523, 32'h00000000} /* (4, 3, 24) {real, imag} */,
  {32'hbf820e80, 32'h00000000} /* (4, 3, 23) {real, imag} */,
  {32'hbf39779f, 32'h00000000} /* (4, 3, 22) {real, imag} */,
  {32'hbf0a2013, 32'h00000000} /* (4, 3, 21) {real, imag} */,
  {32'hbf168e60, 32'h00000000} /* (4, 3, 20) {real, imag} */,
  {32'hbf8056da, 32'h00000000} /* (4, 3, 19) {real, imag} */,
  {32'hbfa5f84b, 32'h00000000} /* (4, 3, 18) {real, imag} */,
  {32'hbf91b9e8, 32'h00000000} /* (4, 3, 17) {real, imag} */,
  {32'hbf7a1d62, 32'h00000000} /* (4, 3, 16) {real, imag} */,
  {32'h3edb71c3, 32'h00000000} /* (4, 3, 15) {real, imag} */,
  {32'h3f9dd21f, 32'h00000000} /* (4, 3, 14) {real, imag} */,
  {32'h3fa2dd31, 32'h00000000} /* (4, 3, 13) {real, imag} */,
  {32'h3f34d89a, 32'h00000000} /* (4, 3, 12) {real, imag} */,
  {32'h3f116709, 32'h00000000} /* (4, 3, 11) {real, imag} */,
  {32'h3f5d25f0, 32'h00000000} /* (4, 3, 10) {real, imag} */,
  {32'h3f1ecac8, 32'h00000000} /* (4, 3, 9) {real, imag} */,
  {32'h3f3138ed, 32'h00000000} /* (4, 3, 8) {real, imag} */,
  {32'h3f5ba80e, 32'h00000000} /* (4, 3, 7) {real, imag} */,
  {32'h3fa10846, 32'h00000000} /* (4, 3, 6) {real, imag} */,
  {32'h3f1f2e9f, 32'h00000000} /* (4, 3, 5) {real, imag} */,
  {32'hbf15cbf1, 32'h00000000} /* (4, 3, 4) {real, imag} */,
  {32'hbfcd2333, 32'h00000000} /* (4, 3, 3) {real, imag} */,
  {32'hbf9e3f7c, 32'h00000000} /* (4, 3, 2) {real, imag} */,
  {32'hbf6c35e8, 32'h00000000} /* (4, 3, 1) {real, imag} */,
  {32'hbe8907f6, 32'h00000000} /* (4, 3, 0) {real, imag} */,
  {32'hbec649f5, 32'h00000000} /* (4, 2, 31) {real, imag} */,
  {32'hbf23ace0, 32'h00000000} /* (4, 2, 30) {real, imag} */,
  {32'hbf54bf9c, 32'h00000000} /* (4, 2, 29) {real, imag} */,
  {32'hbf9ac144, 32'h00000000} /* (4, 2, 28) {real, imag} */,
  {32'hbf78e2b8, 32'h00000000} /* (4, 2, 27) {real, imag} */,
  {32'hbf712bfc, 32'h00000000} /* (4, 2, 26) {real, imag} */,
  {32'hbf14de83, 32'h00000000} /* (4, 2, 25) {real, imag} */,
  {32'hbe1eb284, 32'h00000000} /* (4, 2, 24) {real, imag} */,
  {32'hbf004f23, 32'h00000000} /* (4, 2, 23) {real, imag} */,
  {32'hbeb995a9, 32'h00000000} /* (4, 2, 22) {real, imag} */,
  {32'hbf4eb2cd, 32'h00000000} /* (4, 2, 21) {real, imag} */,
  {32'hbfadf5f8, 32'h00000000} /* (4, 2, 20) {real, imag} */,
  {32'hbf9ecbad, 32'h00000000} /* (4, 2, 19) {real, imag} */,
  {32'hbf8b13dc, 32'h00000000} /* (4, 2, 18) {real, imag} */,
  {32'hbf5dd1c7, 32'h00000000} /* (4, 2, 17) {real, imag} */,
  {32'hbec87a60, 32'h00000000} /* (4, 2, 16) {real, imag} */,
  {32'h3f5a8e1f, 32'h00000000} /* (4, 2, 15) {real, imag} */,
  {32'h3f456edf, 32'h00000000} /* (4, 2, 14) {real, imag} */,
  {32'h3f2cc3c0, 32'h00000000} /* (4, 2, 13) {real, imag} */,
  {32'h3f9ae015, 32'h00000000} /* (4, 2, 12) {real, imag} */,
  {32'h3f24e1fa, 32'h00000000} /* (4, 2, 11) {real, imag} */,
  {32'h3f1d5b5f, 32'h00000000} /* (4, 2, 10) {real, imag} */,
  {32'h3f4e6495, 32'h00000000} /* (4, 2, 9) {real, imag} */,
  {32'h3f52c7e4, 32'h00000000} /* (4, 2, 8) {real, imag} */,
  {32'h3f7b0c40, 32'h00000000} /* (4, 2, 7) {real, imag} */,
  {32'h3f8eaaab, 32'h00000000} /* (4, 2, 6) {real, imag} */,
  {32'h3e7edf5d, 32'h00000000} /* (4, 2, 5) {real, imag} */,
  {32'hbf588003, 32'h00000000} /* (4, 2, 4) {real, imag} */,
  {32'hbfa426d1, 32'h00000000} /* (4, 2, 3) {real, imag} */,
  {32'hbf6cdb36, 32'h00000000} /* (4, 2, 2) {real, imag} */,
  {32'hbf69fc9b, 32'h00000000} /* (4, 2, 1) {real, imag} */,
  {32'hbedd4e97, 32'h00000000} /* (4, 2, 0) {real, imag} */,
  {32'hbe02aa11, 32'h00000000} /* (4, 1, 31) {real, imag} */,
  {32'hbf00de9b, 32'h00000000} /* (4, 1, 30) {real, imag} */,
  {32'hbf6d8992, 32'h00000000} /* (4, 1, 29) {real, imag} */,
  {32'hbf53f576, 32'h00000000} /* (4, 1, 28) {real, imag} */,
  {32'hbf63de0a, 32'h00000000} /* (4, 1, 27) {real, imag} */,
  {32'hbf47a89f, 32'h00000000} /* (4, 1, 26) {real, imag} */,
  {32'hbf320f14, 32'h00000000} /* (4, 1, 25) {real, imag} */,
  {32'hbee51682, 32'h00000000} /* (4, 1, 24) {real, imag} */,
  {32'hbf6ee6f0, 32'h00000000} /* (4, 1, 23) {real, imag} */,
  {32'hbf49744e, 32'h00000000} /* (4, 1, 22) {real, imag} */,
  {32'hbf8b71fe, 32'h00000000} /* (4, 1, 21) {real, imag} */,
  {32'hbf8087f0, 32'h00000000} /* (4, 1, 20) {real, imag} */,
  {32'hbf475679, 32'h00000000} /* (4, 1, 19) {real, imag} */,
  {32'hbf8390b6, 32'h00000000} /* (4, 1, 18) {real, imag} */,
  {32'hbf532646, 32'h00000000} /* (4, 1, 17) {real, imag} */,
  {32'hbe7ced64, 32'h00000000} /* (4, 1, 16) {real, imag} */,
  {32'h3efd69b8, 32'h00000000} /* (4, 1, 15) {real, imag} */,
  {32'h3f5aea76, 32'h00000000} /* (4, 1, 14) {real, imag} */,
  {32'h3f8beab5, 32'h00000000} /* (4, 1, 13) {real, imag} */,
  {32'h3f342dcf, 32'h00000000} /* (4, 1, 12) {real, imag} */,
  {32'h3ee655a2, 32'h00000000} /* (4, 1, 11) {real, imag} */,
  {32'h3f815ef5, 32'h00000000} /* (4, 1, 10) {real, imag} */,
  {32'h3f96a286, 32'h00000000} /* (4, 1, 9) {real, imag} */,
  {32'h3f5638cf, 32'h00000000} /* (4, 1, 8) {real, imag} */,
  {32'h3fac79e8, 32'h00000000} /* (4, 1, 7) {real, imag} */,
  {32'h3fa96545, 32'h00000000} /* (4, 1, 6) {real, imag} */,
  {32'hbee635d3, 32'h00000000} /* (4, 1, 5) {real, imag} */,
  {32'hbfabd73b, 32'h00000000} /* (4, 1, 4) {real, imag} */,
  {32'hbf821119, 32'h00000000} /* (4, 1, 3) {real, imag} */,
  {32'hbed20f8f, 32'h00000000} /* (4, 1, 2) {real, imag} */,
  {32'hbf0f2e20, 32'h00000000} /* (4, 1, 1) {real, imag} */,
  {32'hbe9f60c7, 32'h00000000} /* (4, 1, 0) {real, imag} */,
  {32'hbd29fa10, 32'h00000000} /* (4, 0, 31) {real, imag} */,
  {32'hbe385d3f, 32'h00000000} /* (4, 0, 30) {real, imag} */,
  {32'hbf58ae4d, 32'h00000000} /* (4, 0, 29) {real, imag} */,
  {32'hbf10449e, 32'h00000000} /* (4, 0, 28) {real, imag} */,
  {32'hbe8831fc, 32'h00000000} /* (4, 0, 27) {real, imag} */,
  {32'hbee06553, 32'h00000000} /* (4, 0, 26) {real, imag} */,
  {32'hbefd49e1, 32'h00000000} /* (4, 0, 25) {real, imag} */,
  {32'hbeff7503, 32'h00000000} /* (4, 0, 24) {real, imag} */,
  {32'hbf646320, 32'h00000000} /* (4, 0, 23) {real, imag} */,
  {32'hbf11c1b6, 32'h00000000} /* (4, 0, 22) {real, imag} */,
  {32'hbec8819b, 32'h00000000} /* (4, 0, 21) {real, imag} */,
  {32'hbec11479, 32'h00000000} /* (4, 0, 20) {real, imag} */,
  {32'hbe8395f5, 32'h00000000} /* (4, 0, 19) {real, imag} */,
  {32'hbece6369, 32'h00000000} /* (4, 0, 18) {real, imag} */,
  {32'hbebdf873, 32'h00000000} /* (4, 0, 17) {real, imag} */,
  {32'hbd1075bc, 32'h00000000} /* (4, 0, 16) {real, imag} */,
  {32'h3e660c28, 32'h00000000} /* (4, 0, 15) {real, imag} */,
  {32'h3f31e38c, 32'h00000000} /* (4, 0, 14) {real, imag} */,
  {32'h3f991e33, 32'h00000000} /* (4, 0, 13) {real, imag} */,
  {32'h3ef134ec, 32'h00000000} /* (4, 0, 12) {real, imag} */,
  {32'h3e1a2b0f, 32'h00000000} /* (4, 0, 11) {real, imag} */,
  {32'h3e970789, 32'h00000000} /* (4, 0, 10) {real, imag} */,
  {32'h3eef9e9a, 32'h00000000} /* (4, 0, 9) {real, imag} */,
  {32'h3ea2482e, 32'h00000000} /* (4, 0, 8) {real, imag} */,
  {32'h3f3b6c0c, 32'h00000000} /* (4, 0, 7) {real, imag} */,
  {32'h3f47b4b1, 32'h00000000} /* (4, 0, 6) {real, imag} */,
  {32'hbec940ac, 32'h00000000} /* (4, 0, 5) {real, imag} */,
  {32'hbf628d20, 32'h00000000} /* (4, 0, 4) {real, imag} */,
  {32'hbf2d660a, 32'h00000000} /* (4, 0, 3) {real, imag} */,
  {32'hbe7de941, 32'h00000000} /* (4, 0, 2) {real, imag} */,
  {32'hbebbc97c, 32'h00000000} /* (4, 0, 1) {real, imag} */,
  {32'hbec28f78, 32'h00000000} /* (4, 0, 0) {real, imag} */,
  {32'hbdce2f80, 32'h00000000} /* (3, 31, 31) {real, imag} */,
  {32'hbe52a309, 32'h00000000} /* (3, 31, 30) {real, imag} */,
  {32'hbf020770, 32'h00000000} /* (3, 31, 29) {real, imag} */,
  {32'hbf56b134, 32'h00000000} /* (3, 31, 28) {real, imag} */,
  {32'hbf86e7f9, 32'h00000000} /* (3, 31, 27) {real, imag} */,
  {32'hbf4b4057, 32'h00000000} /* (3, 31, 26) {real, imag} */,
  {32'hbf3c3d64, 32'h00000000} /* (3, 31, 25) {real, imag} */,
  {32'hbf51b940, 32'h00000000} /* (3, 31, 24) {real, imag} */,
  {32'hbf314e69, 32'h00000000} /* (3, 31, 23) {real, imag} */,
  {32'hbef5241c, 32'h00000000} /* (3, 31, 22) {real, imag} */,
  {32'hbe8a29c6, 32'h00000000} /* (3, 31, 21) {real, imag} */,
  {32'h3e63dc4e, 32'h00000000} /* (3, 31, 20) {real, imag} */,
  {32'h3f3381e3, 32'h00000000} /* (3, 31, 19) {real, imag} */,
  {32'h3ea190f8, 32'h00000000} /* (3, 31, 18) {real, imag} */,
  {32'h3e69f368, 32'h00000000} /* (3, 31, 17) {real, imag} */,
  {32'h3e2cfb51, 32'h00000000} /* (3, 31, 16) {real, imag} */,
  {32'h3ec9c1a7, 32'h00000000} /* (3, 31, 15) {real, imag} */,
  {32'h3f84f46c, 32'h00000000} /* (3, 31, 14) {real, imag} */,
  {32'h3f808ab2, 32'h00000000} /* (3, 31, 13) {real, imag} */,
  {32'h3ee4e699, 32'h00000000} /* (3, 31, 12) {real, imag} */,
  {32'h3f05f8d6, 32'h00000000} /* (3, 31, 11) {real, imag} */,
  {32'hbe8dae61, 32'h00000000} /* (3, 31, 10) {real, imag} */,
  {32'hbf3b46fa, 32'h00000000} /* (3, 31, 9) {real, imag} */,
  {32'hbf39b9c2, 32'h00000000} /* (3, 31, 8) {real, imag} */,
  {32'hbf045796, 32'h00000000} /* (3, 31, 7) {real, imag} */,
  {32'hbee38fdc, 32'h00000000} /* (3, 31, 6) {real, imag} */,
  {32'hbe7f2c3e, 32'h00000000} /* (3, 31, 5) {real, imag} */,
  {32'hbe570207, 32'h00000000} /* (3, 31, 4) {real, imag} */,
  {32'hbf284746, 32'h00000000} /* (3, 31, 3) {real, imag} */,
  {32'hbf6d0bf7, 32'h00000000} /* (3, 31, 2) {real, imag} */,
  {32'hbf45f437, 32'h00000000} /* (3, 31, 1) {real, imag} */,
  {32'hbea4ecd8, 32'h00000000} /* (3, 31, 0) {real, imag} */,
  {32'hbeb52cb4, 32'h00000000} /* (3, 30, 31) {real, imag} */,
  {32'hbf156d9e, 32'h00000000} /* (3, 30, 30) {real, imag} */,
  {32'hbf055393, 32'h00000000} /* (3, 30, 29) {real, imag} */,
  {32'hbf98442e, 32'h00000000} /* (3, 30, 28) {real, imag} */,
  {32'hbfcbe236, 32'h00000000} /* (3, 30, 27) {real, imag} */,
  {32'hbfae3528, 32'h00000000} /* (3, 30, 26) {real, imag} */,
  {32'hbf855cff, 32'h00000000} /* (3, 30, 25) {real, imag} */,
  {32'hbf89651b, 32'h00000000} /* (3, 30, 24) {real, imag} */,
  {32'hbf71fbc4, 32'h00000000} /* (3, 30, 23) {real, imag} */,
  {32'hbf5a9942, 32'h00000000} /* (3, 30, 22) {real, imag} */,
  {32'hbf1878a1, 32'h00000000} /* (3, 30, 21) {real, imag} */,
  {32'h3ef55bd4, 32'h00000000} /* (3, 30, 20) {real, imag} */,
  {32'h3fa5bbac, 32'h00000000} /* (3, 30, 19) {real, imag} */,
  {32'h3f4382e6, 32'h00000000} /* (3, 30, 18) {real, imag} */,
  {32'h3f1ff338, 32'h00000000} /* (3, 30, 17) {real, imag} */,
  {32'h3f1b2131, 32'h00000000} /* (3, 30, 16) {real, imag} */,
  {32'h3f4de2f4, 32'h00000000} /* (3, 30, 15) {real, imag} */,
  {32'h3f61c758, 32'h00000000} /* (3, 30, 14) {real, imag} */,
  {32'h3f87965c, 32'h00000000} /* (3, 30, 13) {real, imag} */,
  {32'h3fb01704, 32'h00000000} /* (3, 30, 12) {real, imag} */,
  {32'h3f9311f9, 32'h00000000} /* (3, 30, 11) {real, imag} */,
  {32'hbf246e7d, 32'h00000000} /* (3, 30, 10) {real, imag} */,
  {32'hbfb1e667, 32'h00000000} /* (3, 30, 9) {real, imag} */,
  {32'hbf7a4b12, 32'h00000000} /* (3, 30, 8) {real, imag} */,
  {32'hbf940f39, 32'h00000000} /* (3, 30, 7) {real, imag} */,
  {32'hbf8fb300, 32'h00000000} /* (3, 30, 6) {real, imag} */,
  {32'hbecb081c, 32'h00000000} /* (3, 30, 5) {real, imag} */,
  {32'hbf60fc4a, 32'h00000000} /* (3, 30, 4) {real, imag} */,
  {32'hbf8161e9, 32'h00000000} /* (3, 30, 3) {real, imag} */,
  {32'hbf9a03ed, 32'h00000000} /* (3, 30, 2) {real, imag} */,
  {32'hbf11581d, 32'h00000000} /* (3, 30, 1) {real, imag} */,
  {32'h3d8fac6a, 32'h00000000} /* (3, 30, 0) {real, imag} */,
  {32'hbf1f14c1, 32'h00000000} /* (3, 29, 31) {real, imag} */,
  {32'hbf887b00, 32'h00000000} /* (3, 29, 30) {real, imag} */,
  {32'hbf525ca6, 32'h00000000} /* (3, 29, 29) {real, imag} */,
  {32'hbf85cf8a, 32'h00000000} /* (3, 29, 28) {real, imag} */,
  {32'hbfb88183, 32'h00000000} /* (3, 29, 27) {real, imag} */,
  {32'hbf94f524, 32'h00000000} /* (3, 29, 26) {real, imag} */,
  {32'hbfb3ded0, 32'h00000000} /* (3, 29, 25) {real, imag} */,
  {32'hbfaafb85, 32'h00000000} /* (3, 29, 24) {real, imag} */,
  {32'hbf63f514, 32'h00000000} /* (3, 29, 23) {real, imag} */,
  {32'hbf6c8b5c, 32'h00000000} /* (3, 29, 22) {real, imag} */,
  {32'hbed1fc96, 32'h00000000} /* (3, 29, 21) {real, imag} */,
  {32'h3f7b17b8, 32'h00000000} /* (3, 29, 20) {real, imag} */,
  {32'h400018bf, 32'h00000000} /* (3, 29, 19) {real, imag} */,
  {32'h3f9c7303, 32'h00000000} /* (3, 29, 18) {real, imag} */,
  {32'h3f9c4936, 32'h00000000} /* (3, 29, 17) {real, imag} */,
  {32'h3f98704a, 32'h00000000} /* (3, 29, 16) {real, imag} */,
  {32'h3f4e2b16, 32'h00000000} /* (3, 29, 15) {real, imag} */,
  {32'h3e9bba74, 32'h00000000} /* (3, 29, 14) {real, imag} */,
  {32'h3efe0366, 32'h00000000} /* (3, 29, 13) {real, imag} */,
  {32'h3ffdef99, 32'h00000000} /* (3, 29, 12) {real, imag} */,
  {32'h3fb81665, 32'h00000000} /* (3, 29, 11) {real, imag} */,
  {32'hbf1ef4b9, 32'h00000000} /* (3, 29, 10) {real, imag} */,
  {32'hbf95f461, 32'h00000000} /* (3, 29, 9) {real, imag} */,
  {32'hbf36e160, 32'h00000000} /* (3, 29, 8) {real, imag} */,
  {32'hbf75817e, 32'h00000000} /* (3, 29, 7) {real, imag} */,
  {32'hbf1f491e, 32'h00000000} /* (3, 29, 6) {real, imag} */,
  {32'hbee61f15, 32'h00000000} /* (3, 29, 5) {real, imag} */,
  {32'hbfa7c962, 32'h00000000} /* (3, 29, 4) {real, imag} */,
  {32'hbf8bd596, 32'h00000000} /* (3, 29, 3) {real, imag} */,
  {32'hbf0fc4ba, 32'h00000000} /* (3, 29, 2) {real, imag} */,
  {32'hbea94ed2, 32'h00000000} /* (3, 29, 1) {real, imag} */,
  {32'hbdb4ab8c, 32'h00000000} /* (3, 29, 0) {real, imag} */,
  {32'hbe9a50be, 32'h00000000} /* (3, 28, 31) {real, imag} */,
  {32'hbf3fc8a9, 32'h00000000} /* (3, 28, 30) {real, imag} */,
  {32'hbf70b8e0, 32'h00000000} /* (3, 28, 29) {real, imag} */,
  {32'hbfa73010, 32'h00000000} /* (3, 28, 28) {real, imag} */,
  {32'hbfd1d862, 32'h00000000} /* (3, 28, 27) {real, imag} */,
  {32'hbf50a844, 32'h00000000} /* (3, 28, 26) {real, imag} */,
  {32'hbf3dcf50, 32'h00000000} /* (3, 28, 25) {real, imag} */,
  {32'hbf56e713, 32'h00000000} /* (3, 28, 24) {real, imag} */,
  {32'hbf588036, 32'h00000000} /* (3, 28, 23) {real, imag} */,
  {32'hbf9d6b46, 32'h00000000} /* (3, 28, 22) {real, imag} */,
  {32'hbeb9c351, 32'h00000000} /* (3, 28, 21) {real, imag} */,
  {32'h3f7db685, 32'h00000000} /* (3, 28, 20) {real, imag} */,
  {32'h3fb663f9, 32'h00000000} /* (3, 28, 19) {real, imag} */,
  {32'h3f28370e, 32'h00000000} /* (3, 28, 18) {real, imag} */,
  {32'h3f809066, 32'h00000000} /* (3, 28, 17) {real, imag} */,
  {32'h3f9c7a87, 32'h00000000} /* (3, 28, 16) {real, imag} */,
  {32'h3f3aafed, 32'h00000000} /* (3, 28, 15) {real, imag} */,
  {32'h3f0ad610, 32'h00000000} /* (3, 28, 14) {real, imag} */,
  {32'h3f13a27d, 32'h00000000} /* (3, 28, 13) {real, imag} */,
  {32'h3fba7640, 32'h00000000} /* (3, 28, 12) {real, imag} */,
  {32'h3f6c1bcf, 32'h00000000} /* (3, 28, 11) {real, imag} */,
  {32'hbed8cdac, 32'h00000000} /* (3, 28, 10) {real, imag} */,
  {32'hbf759801, 32'h00000000} /* (3, 28, 9) {real, imag} */,
  {32'hbf6fccec, 32'h00000000} /* (3, 28, 8) {real, imag} */,
  {32'hbf6798f1, 32'h00000000} /* (3, 28, 7) {real, imag} */,
  {32'hbeb22ffc, 32'h00000000} /* (3, 28, 6) {real, imag} */,
  {32'hbf15b453, 32'h00000000} /* (3, 28, 5) {real, imag} */,
  {32'hbf8d4eb8, 32'h00000000} /* (3, 28, 4) {real, imag} */,
  {32'hbf972e8b, 32'h00000000} /* (3, 28, 3) {real, imag} */,
  {32'hbf3c1707, 32'h00000000} /* (3, 28, 2) {real, imag} */,
  {32'hbf06a7b7, 32'h00000000} /* (3, 28, 1) {real, imag} */,
  {32'hbe780309, 32'h00000000} /* (3, 28, 0) {real, imag} */,
  {32'hbe5ebc11, 32'h00000000} /* (3, 27, 31) {real, imag} */,
  {32'hbef97069, 32'h00000000} /* (3, 27, 30) {real, imag} */,
  {32'hbf161879, 32'h00000000} /* (3, 27, 29) {real, imag} */,
  {32'hbf2f6c85, 32'h00000000} /* (3, 27, 28) {real, imag} */,
  {32'hbf846b36, 32'h00000000} /* (3, 27, 27) {real, imag} */,
  {32'hbf7f2e3e, 32'h00000000} /* (3, 27, 26) {real, imag} */,
  {32'hbf66e805, 32'h00000000} /* (3, 27, 25) {real, imag} */,
  {32'hbf7375fd, 32'h00000000} /* (3, 27, 24) {real, imag} */,
  {32'hbfa30b0e, 32'h00000000} /* (3, 27, 23) {real, imag} */,
  {32'hbfa9efd0, 32'h00000000} /* (3, 27, 22) {real, imag} */,
  {32'hbea9f740, 32'h00000000} /* (3, 27, 21) {real, imag} */,
  {32'h3f5771a2, 32'h00000000} /* (3, 27, 20) {real, imag} */,
  {32'h3fa59250, 32'h00000000} /* (3, 27, 19) {real, imag} */,
  {32'h3f50a7d9, 32'h00000000} /* (3, 27, 18) {real, imag} */,
  {32'h3f313ae8, 32'h00000000} /* (3, 27, 17) {real, imag} */,
  {32'h3eaf170a, 32'h00000000} /* (3, 27, 16) {real, imag} */,
  {32'h3f335b3d, 32'h00000000} /* (3, 27, 15) {real, imag} */,
  {32'h3f3b446f, 32'h00000000} /* (3, 27, 14) {real, imag} */,
  {32'h3f9a41b1, 32'h00000000} /* (3, 27, 13) {real, imag} */,
  {32'h3fa6bc9e, 32'h00000000} /* (3, 27, 12) {real, imag} */,
  {32'h3f4b7a43, 32'h00000000} /* (3, 27, 11) {real, imag} */,
  {32'hbf398d91, 32'h00000000} /* (3, 27, 10) {real, imag} */,
  {32'hbf36631c, 32'h00000000} /* (3, 27, 9) {real, imag} */,
  {32'hbf0f1ce2, 32'h00000000} /* (3, 27, 8) {real, imag} */,
  {32'hbf1bd869, 32'h00000000} /* (3, 27, 7) {real, imag} */,
  {32'hbf51f8df, 32'h00000000} /* (3, 27, 6) {real, imag} */,
  {32'hbf6ebc74, 32'h00000000} /* (3, 27, 5) {real, imag} */,
  {32'hbf64d5bc, 32'h00000000} /* (3, 27, 4) {real, imag} */,
  {32'hbf8b2a41, 32'h00000000} /* (3, 27, 3) {real, imag} */,
  {32'hbf8eec4b, 32'h00000000} /* (3, 27, 2) {real, imag} */,
  {32'hbf8205c4, 32'h00000000} /* (3, 27, 1) {real, imag} */,
  {32'hbe880813, 32'h00000000} /* (3, 27, 0) {real, imag} */,
  {32'hbe04e444, 32'h00000000} /* (3, 26, 31) {real, imag} */,
  {32'hbeeba839, 32'h00000000} /* (3, 26, 30) {real, imag} */,
  {32'hbf395313, 32'h00000000} /* (3, 26, 29) {real, imag} */,
  {32'hbf1a21c6, 32'h00000000} /* (3, 26, 28) {real, imag} */,
  {32'hbf451a42, 32'h00000000} /* (3, 26, 27) {real, imag} */,
  {32'hbf6b6459, 32'h00000000} /* (3, 26, 26) {real, imag} */,
  {32'hbf8acc2f, 32'h00000000} /* (3, 26, 25) {real, imag} */,
  {32'hbfb725d4, 32'h00000000} /* (3, 26, 24) {real, imag} */,
  {32'hbfc1c9b1, 32'h00000000} /* (3, 26, 23) {real, imag} */,
  {32'hbf7fc1b2, 32'h00000000} /* (3, 26, 22) {real, imag} */,
  {32'h3ded210d, 32'h00000000} /* (3, 26, 21) {real, imag} */,
  {32'h3fa2f74b, 32'h00000000} /* (3, 26, 20) {real, imag} */,
  {32'h3f84051e, 32'h00000000} /* (3, 26, 19) {real, imag} */,
  {32'h3f649e92, 32'h00000000} /* (3, 26, 18) {real, imag} */,
  {32'h3f7aa8d4, 32'h00000000} /* (3, 26, 17) {real, imag} */,
  {32'h3efb578d, 32'h00000000} /* (3, 26, 16) {real, imag} */,
  {32'h3f97617f, 32'h00000000} /* (3, 26, 15) {real, imag} */,
  {32'h3f8dec86, 32'h00000000} /* (3, 26, 14) {real, imag} */,
  {32'h3f65102d, 32'h00000000} /* (3, 26, 13) {real, imag} */,
  {32'h3f941015, 32'h00000000} /* (3, 26, 12) {real, imag} */,
  {32'h3f3028b2, 32'h00000000} /* (3, 26, 11) {real, imag} */,
  {32'hbdfeb2d0, 32'h00000000} /* (3, 26, 10) {real, imag} */,
  {32'hbf381714, 32'h00000000} /* (3, 26, 9) {real, imag} */,
  {32'hbf511670, 32'h00000000} /* (3, 26, 8) {real, imag} */,
  {32'hbf0fd65a, 32'h00000000} /* (3, 26, 7) {real, imag} */,
  {32'hbf2dca86, 32'h00000000} /* (3, 26, 6) {real, imag} */,
  {32'hbf8346a7, 32'h00000000} /* (3, 26, 5) {real, imag} */,
  {32'hbf0a407d, 32'h00000000} /* (3, 26, 4) {real, imag} */,
  {32'hbece1100, 32'h00000000} /* (3, 26, 3) {real, imag} */,
  {32'hbf874e94, 32'h00000000} /* (3, 26, 2) {real, imag} */,
  {32'hbf4f3904, 32'h00000000} /* (3, 26, 1) {real, imag} */,
  {32'hbe4e16a7, 32'h00000000} /* (3, 26, 0) {real, imag} */,
  {32'hbe4a8414, 32'h00000000} /* (3, 25, 31) {real, imag} */,
  {32'hbf200c3e, 32'h00000000} /* (3, 25, 30) {real, imag} */,
  {32'hbf592196, 32'h00000000} /* (3, 25, 29) {real, imag} */,
  {32'hbfabc5d7, 32'h00000000} /* (3, 25, 28) {real, imag} */,
  {32'hbfb4c88b, 32'h00000000} /* (3, 25, 27) {real, imag} */,
  {32'hbfb085e2, 32'h00000000} /* (3, 25, 26) {real, imag} */,
  {32'hbf98f8df, 32'h00000000} /* (3, 25, 25) {real, imag} */,
  {32'hbf9d9603, 32'h00000000} /* (3, 25, 24) {real, imag} */,
  {32'hbfa39fd2, 32'h00000000} /* (3, 25, 23) {real, imag} */,
  {32'hbf960ec9, 32'h00000000} /* (3, 25, 22) {real, imag} */,
  {32'hbd6e6e84, 32'h00000000} /* (3, 25, 21) {real, imag} */,
  {32'h3f99318d, 32'h00000000} /* (3, 25, 20) {real, imag} */,
  {32'h3f8f4048, 32'h00000000} /* (3, 25, 19) {real, imag} */,
  {32'h3f9a204b, 32'h00000000} /* (3, 25, 18) {real, imag} */,
  {32'h3f9c694a, 32'h00000000} /* (3, 25, 17) {real, imag} */,
  {32'h3f6bdf28, 32'h00000000} /* (3, 25, 16) {real, imag} */,
  {32'h3faf8bd9, 32'h00000000} /* (3, 25, 15) {real, imag} */,
  {32'h3f9caf6f, 32'h00000000} /* (3, 25, 14) {real, imag} */,
  {32'h3f00be4b, 32'h00000000} /* (3, 25, 13) {real, imag} */,
  {32'h3f88dce7, 32'h00000000} /* (3, 25, 12) {real, imag} */,
  {32'h3f791115, 32'h00000000} /* (3, 25, 11) {real, imag} */,
  {32'h3b986c0c, 32'h00000000} /* (3, 25, 10) {real, imag} */,
  {32'hbf813022, 32'h00000000} /* (3, 25, 9) {real, imag} */,
  {32'hbf9b96a4, 32'h00000000} /* (3, 25, 8) {real, imag} */,
  {32'hbf6e0519, 32'h00000000} /* (3, 25, 7) {real, imag} */,
  {32'hbf6fb8fa, 32'h00000000} /* (3, 25, 6) {real, imag} */,
  {32'hbf9ffcce, 32'h00000000} /* (3, 25, 5) {real, imag} */,
  {32'hbf5d4799, 32'h00000000} /* (3, 25, 4) {real, imag} */,
  {32'hbf008188, 32'h00000000} /* (3, 25, 3) {real, imag} */,
  {32'hbf8dbae4, 32'h00000000} /* (3, 25, 2) {real, imag} */,
  {32'hbf63895c, 32'h00000000} /* (3, 25, 1) {real, imag} */,
  {32'hbef12110, 32'h00000000} /* (3, 25, 0) {real, imag} */,
  {32'hbee42a18, 32'h00000000} /* (3, 24, 31) {real, imag} */,
  {32'hbf8ee1db, 32'h00000000} /* (3, 24, 30) {real, imag} */,
  {32'hbf86bbaf, 32'h00000000} /* (3, 24, 29) {real, imag} */,
  {32'hbfdabc48, 32'h00000000} /* (3, 24, 28) {real, imag} */,
  {32'hbf931cc1, 32'h00000000} /* (3, 24, 27) {real, imag} */,
  {32'hbf8ea363, 32'h00000000} /* (3, 24, 26) {real, imag} */,
  {32'hbfc0e558, 32'h00000000} /* (3, 24, 25) {real, imag} */,
  {32'hbf8608f5, 32'h00000000} /* (3, 24, 24) {real, imag} */,
  {32'hbf938cea, 32'h00000000} /* (3, 24, 23) {real, imag} */,
  {32'hbf882257, 32'h00000000} /* (3, 24, 22) {real, imag} */,
  {32'hbd6351e3, 32'h00000000} /* (3, 24, 21) {real, imag} */,
  {32'h3f5ea509, 32'h00000000} /* (3, 24, 20) {real, imag} */,
  {32'h3f59a99c, 32'h00000000} /* (3, 24, 19) {real, imag} */,
  {32'h3f8ec12c, 32'h00000000} /* (3, 24, 18) {real, imag} */,
  {32'h3f88618e, 32'h00000000} /* (3, 24, 17) {real, imag} */,
  {32'h3f66df55, 32'h00000000} /* (3, 24, 16) {real, imag} */,
  {32'h3f9b1a6b, 32'h00000000} /* (3, 24, 15) {real, imag} */,
  {32'h3fbf1879, 32'h00000000} /* (3, 24, 14) {real, imag} */,
  {32'h3f371612, 32'h00000000} /* (3, 24, 13) {real, imag} */,
  {32'h3fa0bbc0, 32'h00000000} /* (3, 24, 12) {real, imag} */,
  {32'h3f7c19ed, 32'h00000000} /* (3, 24, 11) {real, imag} */,
  {32'hbef13d75, 32'h00000000} /* (3, 24, 10) {real, imag} */,
  {32'hbf8ce866, 32'h00000000} /* (3, 24, 9) {real, imag} */,
  {32'hbf82c692, 32'h00000000} /* (3, 24, 8) {real, imag} */,
  {32'hbf470d87, 32'h00000000} /* (3, 24, 7) {real, imag} */,
  {32'hbf66098e, 32'h00000000} /* (3, 24, 6) {real, imag} */,
  {32'hbf64b793, 32'h00000000} /* (3, 24, 5) {real, imag} */,
  {32'hbf117d99, 32'h00000000} /* (3, 24, 4) {real, imag} */,
  {32'hbf686583, 32'h00000000} /* (3, 24, 3) {real, imag} */,
  {32'hbf94b934, 32'h00000000} /* (3, 24, 2) {real, imag} */,
  {32'hbf89b9de, 32'h00000000} /* (3, 24, 1) {real, imag} */,
  {32'hbf3a07e9, 32'h00000000} /* (3, 24, 0) {real, imag} */,
  {32'hbf1db606, 32'h00000000} /* (3, 23, 31) {real, imag} */,
  {32'hbf882901, 32'h00000000} /* (3, 23, 30) {real, imag} */,
  {32'hbf96b65c, 32'h00000000} /* (3, 23, 29) {real, imag} */,
  {32'hbfb96561, 32'h00000000} /* (3, 23, 28) {real, imag} */,
  {32'hbfc6b26b, 32'h00000000} /* (3, 23, 27) {real, imag} */,
  {32'hbf904e7c, 32'h00000000} /* (3, 23, 26) {real, imag} */,
  {32'hbf8ad2f3, 32'h00000000} /* (3, 23, 25) {real, imag} */,
  {32'hbf5c1efa, 32'h00000000} /* (3, 23, 24) {real, imag} */,
  {32'hbf2643f2, 32'h00000000} /* (3, 23, 23) {real, imag} */,
  {32'hbf635f95, 32'h00000000} /* (3, 23, 22) {real, imag} */,
  {32'hbe13a043, 32'h00000000} /* (3, 23, 21) {real, imag} */,
  {32'h3f48ff36, 32'h00000000} /* (3, 23, 20) {real, imag} */,
  {32'h3f27125a, 32'h00000000} /* (3, 23, 19) {real, imag} */,
  {32'h3f47b98b, 32'h00000000} /* (3, 23, 18) {real, imag} */,
  {32'h3f6d0864, 32'h00000000} /* (3, 23, 17) {real, imag} */,
  {32'h3f027f53, 32'h00000000} /* (3, 23, 16) {real, imag} */,
  {32'h3f26be43, 32'h00000000} /* (3, 23, 15) {real, imag} */,
  {32'h3fbaa649, 32'h00000000} /* (3, 23, 14) {real, imag} */,
  {32'h3fa54263, 32'h00000000} /* (3, 23, 13) {real, imag} */,
  {32'h3f9b3acb, 32'h00000000} /* (3, 23, 12) {real, imag} */,
  {32'h3f8cdbbd, 32'h00000000} /* (3, 23, 11) {real, imag} */,
  {32'hbeb541da, 32'h00000000} /* (3, 23, 10) {real, imag} */,
  {32'hbf7f390a, 32'h00000000} /* (3, 23, 9) {real, imag} */,
  {32'hbf6bf4d0, 32'h00000000} /* (3, 23, 8) {real, imag} */,
  {32'hbf5f337b, 32'h00000000} /* (3, 23, 7) {real, imag} */,
  {32'hbf2b8b74, 32'h00000000} /* (3, 23, 6) {real, imag} */,
  {32'hbf5af462, 32'h00000000} /* (3, 23, 5) {real, imag} */,
  {32'hbf151a6e, 32'h00000000} /* (3, 23, 4) {real, imag} */,
  {32'hbfbfe5a3, 32'h00000000} /* (3, 23, 3) {real, imag} */,
  {32'hbfa71142, 32'h00000000} /* (3, 23, 2) {real, imag} */,
  {32'hbf8081ab, 32'h00000000} /* (3, 23, 1) {real, imag} */,
  {32'hbf0764d8, 32'h00000000} /* (3, 23, 0) {real, imag} */,
  {32'hbf017f06, 32'h00000000} /* (3, 22, 31) {real, imag} */,
  {32'hbfae9c68, 32'h00000000} /* (3, 22, 30) {real, imag} */,
  {32'hbfb67373, 32'h00000000} /* (3, 22, 29) {real, imag} */,
  {32'hbfae82e6, 32'h00000000} /* (3, 22, 28) {real, imag} */,
  {32'hbfe23012, 32'h00000000} /* (3, 22, 27) {real, imag} */,
  {32'hbfb01476, 32'h00000000} /* (3, 22, 26) {real, imag} */,
  {32'hbf28b4d5, 32'h00000000} /* (3, 22, 25) {real, imag} */,
  {32'hbf564b9a, 32'h00000000} /* (3, 22, 24) {real, imag} */,
  {32'hbf38511a, 32'h00000000} /* (3, 22, 23) {real, imag} */,
  {32'hbe87d73d, 32'h00000000} /* (3, 22, 22) {real, imag} */,
  {32'hbe3567b5, 32'h00000000} /* (3, 22, 21) {real, imag} */,
  {32'h3ef26ee3, 32'h00000000} /* (3, 22, 20) {real, imag} */,
  {32'h3f008df1, 32'h00000000} /* (3, 22, 19) {real, imag} */,
  {32'h3f124979, 32'h00000000} /* (3, 22, 18) {real, imag} */,
  {32'h3f61e7a7, 32'h00000000} /* (3, 22, 17) {real, imag} */,
  {32'h3ea914a0, 32'h00000000} /* (3, 22, 16) {real, imag} */,
  {32'h3e8b79b7, 32'h00000000} /* (3, 22, 15) {real, imag} */,
  {32'h3fa5a0ce, 32'h00000000} /* (3, 22, 14) {real, imag} */,
  {32'h3fb9a230, 32'h00000000} /* (3, 22, 13) {real, imag} */,
  {32'h3f382f96, 32'h00000000} /* (3, 22, 12) {real, imag} */,
  {32'h3eafa398, 32'h00000000} /* (3, 22, 11) {real, imag} */,
  {32'hbefa9837, 32'h00000000} /* (3, 22, 10) {real, imag} */,
  {32'hbf8feeea, 32'h00000000} /* (3, 22, 9) {real, imag} */,
  {32'hbf805669, 32'h00000000} /* (3, 22, 8) {real, imag} */,
  {32'hbf85e5a6, 32'h00000000} /* (3, 22, 7) {real, imag} */,
  {32'hbf4ec8ee, 32'h00000000} /* (3, 22, 6) {real, imag} */,
  {32'hbf9b5451, 32'h00000000} /* (3, 22, 5) {real, imag} */,
  {32'hbf47bd59, 32'h00000000} /* (3, 22, 4) {real, imag} */,
  {32'hbf8bcfd4, 32'h00000000} /* (3, 22, 3) {real, imag} */,
  {32'hbf9ab181, 32'h00000000} /* (3, 22, 2) {real, imag} */,
  {32'hbf74909c, 32'h00000000} /* (3, 22, 1) {real, imag} */,
  {32'hbecc793c, 32'h00000000} /* (3, 22, 0) {real, imag} */,
  {32'h3bd131c4, 32'h00000000} /* (3, 21, 31) {real, imag} */,
  {32'hbdae9d44, 32'h00000000} /* (3, 21, 30) {real, imag} */,
  {32'h3e00d236, 32'h00000000} /* (3, 21, 29) {real, imag} */,
  {32'hbe91229b, 32'h00000000} /* (3, 21, 28) {real, imag} */,
  {32'hbf549482, 32'h00000000} /* (3, 21, 27) {real, imag} */,
  {32'hbf34901d, 32'h00000000} /* (3, 21, 26) {real, imag} */,
  {32'h3e9c9fcb, 32'h00000000} /* (3, 21, 25) {real, imag} */,
  {32'h3dddf5cc, 32'h00000000} /* (3, 21, 24) {real, imag} */,
  {32'hbec55a4b, 32'h00000000} /* (3, 21, 23) {real, imag} */,
  {32'hbe516f94, 32'h00000000} /* (3, 21, 22) {real, imag} */,
  {32'hbe81b9ae, 32'h00000000} /* (3, 21, 21) {real, imag} */,
  {32'hbe3511ce, 32'h00000000} /* (3, 21, 20) {real, imag} */,
  {32'h3e2fcb1b, 32'h00000000} /* (3, 21, 19) {real, imag} */,
  {32'h3e92faa8, 32'h00000000} /* (3, 21, 18) {real, imag} */,
  {32'h3f271c48, 32'h00000000} /* (3, 21, 17) {real, imag} */,
  {32'h3f198f6a, 32'h00000000} /* (3, 21, 16) {real, imag} */,
  {32'h3d0c7485, 32'h00000000} /* (3, 21, 15) {real, imag} */,
  {32'h3ed6be21, 32'h00000000} /* (3, 21, 14) {real, imag} */,
  {32'h3f01742f, 32'h00000000} /* (3, 21, 13) {real, imag} */,
  {32'hbe1e0ce2, 32'h00000000} /* (3, 21, 12) {real, imag} */,
  {32'h3d7e4e6e, 32'h00000000} /* (3, 21, 11) {real, imag} */,
  {32'hbd32f34f, 32'h00000000} /* (3, 21, 10) {real, imag} */,
  {32'hbf426d0b, 32'h00000000} /* (3, 21, 9) {real, imag} */,
  {32'hbf163407, 32'h00000000} /* (3, 21, 8) {real, imag} */,
  {32'h3d88ba7f, 32'h00000000} /* (3, 21, 7) {real, imag} */,
  {32'hbe0a68ca, 32'h00000000} /* (3, 21, 6) {real, imag} */,
  {32'hbeda3a07, 32'h00000000} /* (3, 21, 5) {real, imag} */,
  {32'hbf1b7445, 32'h00000000} /* (3, 21, 4) {real, imag} */,
  {32'hbf646dee, 32'h00000000} /* (3, 21, 3) {real, imag} */,
  {32'hbf027038, 32'h00000000} /* (3, 21, 2) {real, imag} */,
  {32'hbe96e108, 32'h00000000} /* (3, 21, 1) {real, imag} */,
  {32'hbdf1a6dd, 32'h00000000} /* (3, 21, 0) {real, imag} */,
  {32'h3f2c1271, 32'h00000000} /* (3, 20, 31) {real, imag} */,
  {32'h3f80f3de, 32'h00000000} /* (3, 20, 30) {real, imag} */,
  {32'h3f9d726a, 32'h00000000} /* (3, 20, 29) {real, imag} */,
  {32'h3fa6c108, 32'h00000000} /* (3, 20, 28) {real, imag} */,
  {32'h3f7d9887, 32'h00000000} /* (3, 20, 27) {real, imag} */,
  {32'h3f34e6db, 32'h00000000} /* (3, 20, 26) {real, imag} */,
  {32'h3ff3c150, 32'h00000000} /* (3, 20, 25) {real, imag} */,
  {32'h3fcfe5d3, 32'h00000000} /* (3, 20, 24) {real, imag} */,
  {32'h3f78ebd7, 32'h00000000} /* (3, 20, 23) {real, imag} */,
  {32'h3ebe28c7, 32'h00000000} /* (3, 20, 22) {real, imag} */,
  {32'hbe38059d, 32'h00000000} /* (3, 20, 21) {real, imag} */,
  {32'hbf948699, 32'h00000000} /* (3, 20, 20) {real, imag} */,
  {32'hbf1d3db9, 32'h00000000} /* (3, 20, 19) {real, imag} */,
  {32'hbee1f060, 32'h00000000} /* (3, 20, 18) {real, imag} */,
  {32'hbea9ca06, 32'h00000000} /* (3, 20, 17) {real, imag} */,
  {32'hbe268ee6, 32'h00000000} /* (3, 20, 16) {real, imag} */,
  {32'hbf069ad1, 32'h00000000} /* (3, 20, 15) {real, imag} */,
  {32'hbf3e73d5, 32'h00000000} /* (3, 20, 14) {real, imag} */,
  {32'hbf476866, 32'h00000000} /* (3, 20, 13) {real, imag} */,
  {32'hbfa9e8d5, 32'h00000000} /* (3, 20, 12) {real, imag} */,
  {32'hbec5cbf0, 32'h00000000} /* (3, 20, 11) {real, imag} */,
  {32'h3f291406, 32'h00000000} /* (3, 20, 10) {real, imag} */,
  {32'h3e1e7d2c, 32'h00000000} /* (3, 20, 9) {real, imag} */,
  {32'h3ce742fd, 32'h00000000} /* (3, 20, 8) {real, imag} */,
  {32'h3f8e393a, 32'h00000000} /* (3, 20, 7) {real, imag} */,
  {32'h3f5a9161, 32'h00000000} /* (3, 20, 6) {real, imag} */,
  {32'h3f91c6ce, 32'h00000000} /* (3, 20, 5) {real, imag} */,
  {32'h3f1a8299, 32'h00000000} /* (3, 20, 4) {real, imag} */,
  {32'h3e1ec605, 32'h00000000} /* (3, 20, 3) {real, imag} */,
  {32'h3f0277a8, 32'h00000000} /* (3, 20, 2) {real, imag} */,
  {32'h3edd76c6, 32'h00000000} /* (3, 20, 1) {real, imag} */,
  {32'h3e2a134f, 32'h00000000} /* (3, 20, 0) {real, imag} */,
  {32'h3f14ddf0, 32'h00000000} /* (3, 19, 31) {real, imag} */,
  {32'h3f47754f, 32'h00000000} /* (3, 19, 30) {real, imag} */,
  {32'h3f4ba212, 32'h00000000} /* (3, 19, 29) {real, imag} */,
  {32'h3fa5205d, 32'h00000000} /* (3, 19, 28) {real, imag} */,
  {32'h3f87f951, 32'h00000000} /* (3, 19, 27) {real, imag} */,
  {32'h3f6254af, 32'h00000000} /* (3, 19, 26) {real, imag} */,
  {32'h3fe71176, 32'h00000000} /* (3, 19, 25) {real, imag} */,
  {32'h3fdaea8d, 32'h00000000} /* (3, 19, 24) {real, imag} */,
  {32'h3f560b47, 32'h00000000} /* (3, 19, 23) {real, imag} */,
  {32'h3f0a317d, 32'h00000000} /* (3, 19, 22) {real, imag} */,
  {32'hbe851c00, 32'h00000000} /* (3, 19, 21) {real, imag} */,
  {32'hbfcd853d, 32'h00000000} /* (3, 19, 20) {real, imag} */,
  {32'hbf6b246a, 32'h00000000} /* (3, 19, 19) {real, imag} */,
  {32'hbf7f35ec, 32'h00000000} /* (3, 19, 18) {real, imag} */,
  {32'hbf8ef362, 32'h00000000} /* (3, 19, 17) {real, imag} */,
  {32'hbf016ba5, 32'h00000000} /* (3, 19, 16) {real, imag} */,
  {32'hbf5e33af, 32'h00000000} /* (3, 19, 15) {real, imag} */,
  {32'hbf45ecd3, 32'h00000000} /* (3, 19, 14) {real, imag} */,
  {32'hbf73f006, 32'h00000000} /* (3, 19, 13) {real, imag} */,
  {32'hbfd33bd9, 32'h00000000} /* (3, 19, 12) {real, imag} */,
  {32'hbf8f5026, 32'h00000000} /* (3, 19, 11) {real, imag} */,
  {32'h3f2cfba6, 32'h00000000} /* (3, 19, 10) {real, imag} */,
  {32'h3f483d4f, 32'h00000000} /* (3, 19, 9) {real, imag} */,
  {32'h3f40a5f7, 32'h00000000} /* (3, 19, 8) {real, imag} */,
  {32'h3f994012, 32'h00000000} /* (3, 19, 7) {real, imag} */,
  {32'h3ec11a95, 32'h00000000} /* (3, 19, 6) {real, imag} */,
  {32'h3f7099c1, 32'h00000000} /* (3, 19, 5) {real, imag} */,
  {32'h3f831aaf, 32'h00000000} /* (3, 19, 4) {real, imag} */,
  {32'h3f259dcc, 32'h00000000} /* (3, 19, 3) {real, imag} */,
  {32'h3f0e567f, 32'h00000000} /* (3, 19, 2) {real, imag} */,
  {32'h3f55ab07, 32'h00000000} /* (3, 19, 1) {real, imag} */,
  {32'h3ef5c685, 32'h00000000} /* (3, 19, 0) {real, imag} */,
  {32'h3ea38c5e, 32'h00000000} /* (3, 18, 31) {real, imag} */,
  {32'h3f296a4b, 32'h00000000} /* (3, 18, 30) {real, imag} */,
  {32'h3f3a2059, 32'h00000000} /* (3, 18, 29) {real, imag} */,
  {32'h3f8e5547, 32'h00000000} /* (3, 18, 28) {real, imag} */,
  {32'h3f2cd5f8, 32'h00000000} /* (3, 18, 27) {real, imag} */,
  {32'h3f98f040, 32'h00000000} /* (3, 18, 26) {real, imag} */,
  {32'h3f92e588, 32'h00000000} /* (3, 18, 25) {real, imag} */,
  {32'h3fb39cf7, 32'h00000000} /* (3, 18, 24) {real, imag} */,
  {32'h3f4165c3, 32'h00000000} /* (3, 18, 23) {real, imag} */,
  {32'h3f1c3a4a, 32'h00000000} /* (3, 18, 22) {real, imag} */,
  {32'h3e4c7fde, 32'h00000000} /* (3, 18, 21) {real, imag} */,
  {32'hbfc332eb, 32'h00000000} /* (3, 18, 20) {real, imag} */,
  {32'hbf4a2d47, 32'h00000000} /* (3, 18, 19) {real, imag} */,
  {32'hbf97ce4f, 32'h00000000} /* (3, 18, 18) {real, imag} */,
  {32'hbfb2e124, 32'h00000000} /* (3, 18, 17) {real, imag} */,
  {32'hbef5d37f, 32'h00000000} /* (3, 18, 16) {real, imag} */,
  {32'hbf8904ee, 32'h00000000} /* (3, 18, 15) {real, imag} */,
  {32'hbf968e31, 32'h00000000} /* (3, 18, 14) {real, imag} */,
  {32'hbfadf64c, 32'h00000000} /* (3, 18, 13) {real, imag} */,
  {32'hbfda51dd, 32'h00000000} /* (3, 18, 12) {real, imag} */,
  {32'hbfe7d214, 32'h00000000} /* (3, 18, 11) {real, imag} */,
  {32'hbd527630, 32'h00000000} /* (3, 18, 10) {real, imag} */,
  {32'h3f654b09, 32'h00000000} /* (3, 18, 9) {real, imag} */,
  {32'h3fabc5c0, 32'h00000000} /* (3, 18, 8) {real, imag} */,
  {32'h3f9b5a4f, 32'h00000000} /* (3, 18, 7) {real, imag} */,
  {32'h3f078b8e, 32'h00000000} /* (3, 18, 6) {real, imag} */,
  {32'h3f5545e1, 32'h00000000} /* (3, 18, 5) {real, imag} */,
  {32'h3f82e0fd, 32'h00000000} /* (3, 18, 4) {real, imag} */,
  {32'h3f4112fa, 32'h00000000} /* (3, 18, 3) {real, imag} */,
  {32'h3f1f2328, 32'h00000000} /* (3, 18, 2) {real, imag} */,
  {32'h3f28f1bb, 32'h00000000} /* (3, 18, 1) {real, imag} */,
  {32'h3ea3c655, 32'h00000000} /* (3, 18, 0) {real, imag} */,
  {32'h3f1852d1, 32'h00000000} /* (3, 17, 31) {real, imag} */,
  {32'h3f748f99, 32'h00000000} /* (3, 17, 30) {real, imag} */,
  {32'h3f5bf995, 32'h00000000} /* (3, 17, 29) {real, imag} */,
  {32'h3f662aa3, 32'h00000000} /* (3, 17, 28) {real, imag} */,
  {32'h3f61d262, 32'h00000000} /* (3, 17, 27) {real, imag} */,
  {32'h3fa827e4, 32'h00000000} /* (3, 17, 26) {real, imag} */,
  {32'h3f68fc35, 32'h00000000} /* (3, 17, 25) {real, imag} */,
  {32'h3f2bf7a7, 32'h00000000} /* (3, 17, 24) {real, imag} */,
  {32'h3f3bec6d, 32'h00000000} /* (3, 17, 23) {real, imag} */,
  {32'h3f295210, 32'h00000000} /* (3, 17, 22) {real, imag} */,
  {32'h3c922604, 32'h00000000} /* (3, 17, 21) {real, imag} */,
  {32'hbfacf376, 32'h00000000} /* (3, 17, 20) {real, imag} */,
  {32'hbf74f091, 32'h00000000} /* (3, 17, 19) {real, imag} */,
  {32'hbf81ee3b, 32'h00000000} /* (3, 17, 18) {real, imag} */,
  {32'hbfb003f3, 32'h00000000} /* (3, 17, 17) {real, imag} */,
  {32'hbfa50223, 32'h00000000} /* (3, 17, 16) {real, imag} */,
  {32'hbf9a4eea, 32'h00000000} /* (3, 17, 15) {real, imag} */,
  {32'hbf800d02, 32'h00000000} /* (3, 17, 14) {real, imag} */,
  {32'hbf77e717, 32'h00000000} /* (3, 17, 13) {real, imag} */,
  {32'hbf338c38, 32'h00000000} /* (3, 17, 12) {real, imag} */,
  {32'hbf8a5d8a, 32'h00000000} /* (3, 17, 11) {real, imag} */,
  {32'h3e167cb5, 32'h00000000} /* (3, 17, 10) {real, imag} */,
  {32'h3f3ea851, 32'h00000000} /* (3, 17, 9) {real, imag} */,
  {32'h3f222208, 32'h00000000} /* (3, 17, 8) {real, imag} */,
  {32'h3f380140, 32'h00000000} /* (3, 17, 7) {real, imag} */,
  {32'h3f3d3b24, 32'h00000000} /* (3, 17, 6) {real, imag} */,
  {32'h3f8388dc, 32'h00000000} /* (3, 17, 5) {real, imag} */,
  {32'h3fa89fc6, 32'h00000000} /* (3, 17, 4) {real, imag} */,
  {32'h3f64f6af, 32'h00000000} /* (3, 17, 3) {real, imag} */,
  {32'h3f009f38, 32'h00000000} /* (3, 17, 2) {real, imag} */,
  {32'h3eb9a7fd, 32'h00000000} /* (3, 17, 1) {real, imag} */,
  {32'h3ef36bce, 32'h00000000} /* (3, 17, 0) {real, imag} */,
  {32'h3f4f3128, 32'h00000000} /* (3, 16, 31) {real, imag} */,
  {32'h3fabf6b8, 32'h00000000} /* (3, 16, 30) {real, imag} */,
  {32'h3f52fbb5, 32'h00000000} /* (3, 16, 29) {real, imag} */,
  {32'h3ed62418, 32'h00000000} /* (3, 16, 28) {real, imag} */,
  {32'h3f012dfe, 32'h00000000} /* (3, 16, 27) {real, imag} */,
  {32'h3f402580, 32'h00000000} /* (3, 16, 26) {real, imag} */,
  {32'h3f7512ae, 32'h00000000} /* (3, 16, 25) {real, imag} */,
  {32'h3f25ef32, 32'h00000000} /* (3, 16, 24) {real, imag} */,
  {32'h3f308faf, 32'h00000000} /* (3, 16, 23) {real, imag} */,
  {32'h3f43541e, 32'h00000000} /* (3, 16, 22) {real, imag} */,
  {32'h3e4f3994, 32'h00000000} /* (3, 16, 21) {real, imag} */,
  {32'hbfa7d4cc, 32'h00000000} /* (3, 16, 20) {real, imag} */,
  {32'hbfa9f9d9, 32'h00000000} /* (3, 16, 19) {real, imag} */,
  {32'hbf8fc386, 32'h00000000} /* (3, 16, 18) {real, imag} */,
  {32'hbfac1de4, 32'h00000000} /* (3, 16, 17) {real, imag} */,
  {32'hbfcee735, 32'h00000000} /* (3, 16, 16) {real, imag} */,
  {32'hbfc43d08, 32'h00000000} /* (3, 16, 15) {real, imag} */,
  {32'hbf564654, 32'h00000000} /* (3, 16, 14) {real, imag} */,
  {32'hbf98f67b, 32'h00000000} /* (3, 16, 13) {real, imag} */,
  {32'hbf7b2664, 32'h00000000} /* (3, 16, 12) {real, imag} */,
  {32'hbf671390, 32'h00000000} /* (3, 16, 11) {real, imag} */,
  {32'h3e90a680, 32'h00000000} /* (3, 16, 10) {real, imag} */,
  {32'h3f724498, 32'h00000000} /* (3, 16, 9) {real, imag} */,
  {32'h3f3b6070, 32'h00000000} /* (3, 16, 8) {real, imag} */,
  {32'h3f511789, 32'h00000000} /* (3, 16, 7) {real, imag} */,
  {32'h3f0c25c9, 32'h00000000} /* (3, 16, 6) {real, imag} */,
  {32'h3f4e7f37, 32'h00000000} /* (3, 16, 5) {real, imag} */,
  {32'h3f6f8347, 32'h00000000} /* (3, 16, 4) {real, imag} */,
  {32'h3f9fb25d, 32'h00000000} /* (3, 16, 3) {real, imag} */,
  {32'h3f9b07b4, 32'h00000000} /* (3, 16, 2) {real, imag} */,
  {32'h3f70d38f, 32'h00000000} /* (3, 16, 1) {real, imag} */,
  {32'h3f7d1376, 32'h00000000} /* (3, 16, 0) {real, imag} */,
  {32'h3f2c8616, 32'h00000000} /* (3, 15, 31) {real, imag} */,
  {32'h3f863ea5, 32'h00000000} /* (3, 15, 30) {real, imag} */,
  {32'h3f20a07e, 32'h00000000} /* (3, 15, 29) {real, imag} */,
  {32'h3f0be66d, 32'h00000000} /* (3, 15, 28) {real, imag} */,
  {32'h3f616ff1, 32'h00000000} /* (3, 15, 27) {real, imag} */,
  {32'h3f52c15b, 32'h00000000} /* (3, 15, 26) {real, imag} */,
  {32'h3f54abc5, 32'h00000000} /* (3, 15, 25) {real, imag} */,
  {32'h3f5f5d36, 32'h00000000} /* (3, 15, 24) {real, imag} */,
  {32'h3f9d76f8, 32'h00000000} /* (3, 15, 23) {real, imag} */,
  {32'h3fbeb9cf, 32'h00000000} /* (3, 15, 22) {real, imag} */,
  {32'h3f29b625, 32'h00000000} /* (3, 15, 21) {real, imag} */,
  {32'hbf644b10, 32'h00000000} /* (3, 15, 20) {real, imag} */,
  {32'hbf57a874, 32'h00000000} /* (3, 15, 19) {real, imag} */,
  {32'hbf3414bc, 32'h00000000} /* (3, 15, 18) {real, imag} */,
  {32'hbf49f7b5, 32'h00000000} /* (3, 15, 17) {real, imag} */,
  {32'hbf39cba9, 32'h00000000} /* (3, 15, 16) {real, imag} */,
  {32'hbf5c34bd, 32'h00000000} /* (3, 15, 15) {real, imag} */,
  {32'hbf32dcb6, 32'h00000000} /* (3, 15, 14) {real, imag} */,
  {32'hbf790f13, 32'h00000000} /* (3, 15, 13) {real, imag} */,
  {32'hbf8bd01f, 32'h00000000} /* (3, 15, 12) {real, imag} */,
  {32'hbf2a68a7, 32'h00000000} /* (3, 15, 11) {real, imag} */,
  {32'h3ef618b7, 32'h00000000} /* (3, 15, 10) {real, imag} */,
  {32'h3f752aa9, 32'h00000000} /* (3, 15, 9) {real, imag} */,
  {32'h3f3ba5f0, 32'h00000000} /* (3, 15, 8) {real, imag} */,
  {32'h3f598195, 32'h00000000} /* (3, 15, 7) {real, imag} */,
  {32'h3ef4b39f, 32'h00000000} /* (3, 15, 6) {real, imag} */,
  {32'h3f623921, 32'h00000000} /* (3, 15, 5) {real, imag} */,
  {32'h3f4188f3, 32'h00000000} /* (3, 15, 4) {real, imag} */,
  {32'h3f8e5199, 32'h00000000} /* (3, 15, 3) {real, imag} */,
  {32'h3f9d5641, 32'h00000000} /* (3, 15, 2) {real, imag} */,
  {32'h3f705b5c, 32'h00000000} /* (3, 15, 1) {real, imag} */,
  {32'h3f536193, 32'h00000000} /* (3, 15, 0) {real, imag} */,
  {32'h3f18f74c, 32'h00000000} /* (3, 14, 31) {real, imag} */,
  {32'h3f410d32, 32'h00000000} /* (3, 14, 30) {real, imag} */,
  {32'h3f30a376, 32'h00000000} /* (3, 14, 29) {real, imag} */,
  {32'h3f770d61, 32'h00000000} /* (3, 14, 28) {real, imag} */,
  {32'h3f781682, 32'h00000000} /* (3, 14, 27) {real, imag} */,
  {32'h3f5d9a38, 32'h00000000} /* (3, 14, 26) {real, imag} */,
  {32'h3edbe85b, 32'h00000000} /* (3, 14, 25) {real, imag} */,
  {32'h3f151fc0, 32'h00000000} /* (3, 14, 24) {real, imag} */,
  {32'h3f99c9f6, 32'h00000000} /* (3, 14, 23) {real, imag} */,
  {32'h3fe89479, 32'h00000000} /* (3, 14, 22) {real, imag} */,
  {32'h3f995ca6, 32'h00000000} /* (3, 14, 21) {real, imag} */,
  {32'hbf26e3aa, 32'h00000000} /* (3, 14, 20) {real, imag} */,
  {32'hbf833444, 32'h00000000} /* (3, 14, 19) {real, imag} */,
  {32'hbf66dac5, 32'h00000000} /* (3, 14, 18) {real, imag} */,
  {32'hbf6257b0, 32'h00000000} /* (3, 14, 17) {real, imag} */,
  {32'hbf908480, 32'h00000000} /* (3, 14, 16) {real, imag} */,
  {32'hbf3a5f2d, 32'h00000000} /* (3, 14, 15) {real, imag} */,
  {32'hbe9af26e, 32'h00000000} /* (3, 14, 14) {real, imag} */,
  {32'hbf16693e, 32'h00000000} /* (3, 14, 13) {real, imag} */,
  {32'hbf34da9e, 32'h00000000} /* (3, 14, 12) {real, imag} */,
  {32'hbedf1ebc, 32'h00000000} /* (3, 14, 11) {real, imag} */,
  {32'h3f217fad, 32'h00000000} /* (3, 14, 10) {real, imag} */,
  {32'h3f943bcf, 32'h00000000} /* (3, 14, 9) {real, imag} */,
  {32'h3f9cac46, 32'h00000000} /* (3, 14, 8) {real, imag} */,
  {32'h3f748587, 32'h00000000} /* (3, 14, 7) {real, imag} */,
  {32'h3f4877e2, 32'h00000000} /* (3, 14, 6) {real, imag} */,
  {32'h3f709329, 32'h00000000} /* (3, 14, 5) {real, imag} */,
  {32'h3f28eb20, 32'h00000000} /* (3, 14, 4) {real, imag} */,
  {32'h3f6b1aab, 32'h00000000} /* (3, 14, 3) {real, imag} */,
  {32'h3f8ee27c, 32'h00000000} /* (3, 14, 2) {real, imag} */,
  {32'h3fa0d340, 32'h00000000} /* (3, 14, 1) {real, imag} */,
  {32'h3f5b3968, 32'h00000000} /* (3, 14, 0) {real, imag} */,
  {32'h3f08f53f, 32'h00000000} /* (3, 13, 31) {real, imag} */,
  {32'h3f90676c, 32'h00000000} /* (3, 13, 30) {real, imag} */,
  {32'h3fb98e12, 32'h00000000} /* (3, 13, 29) {real, imag} */,
  {32'h3fb3a7fc, 32'h00000000} /* (3, 13, 28) {real, imag} */,
  {32'h3f0f21c6, 32'h00000000} /* (3, 13, 27) {real, imag} */,
  {32'h3f5158cf, 32'h00000000} /* (3, 13, 26) {real, imag} */,
  {32'h3f6a4424, 32'h00000000} /* (3, 13, 25) {real, imag} */,
  {32'h3f76db0b, 32'h00000000} /* (3, 13, 24) {real, imag} */,
  {32'h3f91bec8, 32'h00000000} /* (3, 13, 23) {real, imag} */,
  {32'h3fbebec7, 32'h00000000} /* (3, 13, 22) {real, imag} */,
  {32'h3f45ca1a, 32'h00000000} /* (3, 13, 21) {real, imag} */,
  {32'hbf4c5408, 32'h00000000} /* (3, 13, 20) {real, imag} */,
  {32'hbf8fe3b3, 32'h00000000} /* (3, 13, 19) {real, imag} */,
  {32'hbf07e3e0, 32'h00000000} /* (3, 13, 18) {real, imag} */,
  {32'hbf95ced4, 32'h00000000} /* (3, 13, 17) {real, imag} */,
  {32'hbf9ccc82, 32'h00000000} /* (3, 13, 16) {real, imag} */,
  {32'hbefb86a8, 32'h00000000} /* (3, 13, 15) {real, imag} */,
  {32'hbf27ec56, 32'h00000000} /* (3, 13, 14) {real, imag} */,
  {32'hbf3ab246, 32'h00000000} /* (3, 13, 13) {real, imag} */,
  {32'hbf189e46, 32'h00000000} /* (3, 13, 12) {real, imag} */,
  {32'hbefd4a54, 32'h00000000} /* (3, 13, 11) {real, imag} */,
  {32'h3edb2945, 32'h00000000} /* (3, 13, 10) {real, imag} */,
  {32'h3f1ebe4f, 32'h00000000} /* (3, 13, 9) {real, imag} */,
  {32'h3f44444a, 32'h00000000} /* (3, 13, 8) {real, imag} */,
  {32'h3f7f8106, 32'h00000000} /* (3, 13, 7) {real, imag} */,
  {32'h3f41e9ff, 32'h00000000} /* (3, 13, 6) {real, imag} */,
  {32'h3f313c70, 32'h00000000} /* (3, 13, 5) {real, imag} */,
  {32'h3ea893aa, 32'h00000000} /* (3, 13, 4) {real, imag} */,
  {32'h3f21325d, 32'h00000000} /* (3, 13, 3) {real, imag} */,
  {32'h3f945c13, 32'h00000000} /* (3, 13, 2) {real, imag} */,
  {32'h3ff1fce7, 32'h00000000} /* (3, 13, 1) {real, imag} */,
  {32'h3f72f921, 32'h00000000} /* (3, 13, 0) {real, imag} */,
  {32'h3e905e04, 32'h00000000} /* (3, 12, 31) {real, imag} */,
  {32'h3f82e635, 32'h00000000} /* (3, 12, 30) {real, imag} */,
  {32'h3fb1d680, 32'h00000000} /* (3, 12, 29) {real, imag} */,
  {32'h3f97eb7a, 32'h00000000} /* (3, 12, 28) {real, imag} */,
  {32'h3f21525f, 32'h00000000} /* (3, 12, 27) {real, imag} */,
  {32'h3ec21762, 32'h00000000} /* (3, 12, 26) {real, imag} */,
  {32'h3f706e89, 32'h00000000} /* (3, 12, 25) {real, imag} */,
  {32'h3fb6f5c9, 32'h00000000} /* (3, 12, 24) {real, imag} */,
  {32'h3f730288, 32'h00000000} /* (3, 12, 23) {real, imag} */,
  {32'h3f7ee209, 32'h00000000} /* (3, 12, 22) {real, imag} */,
  {32'h3e681011, 32'h00000000} /* (3, 12, 21) {real, imag} */,
  {32'hbf4ea55b, 32'h00000000} /* (3, 12, 20) {real, imag} */,
  {32'hbf4333a2, 32'h00000000} /* (3, 12, 19) {real, imag} */,
  {32'hbf20d7a1, 32'h00000000} /* (3, 12, 18) {real, imag} */,
  {32'hbf5d1b99, 32'h00000000} /* (3, 12, 17) {real, imag} */,
  {32'hbf8ca4a5, 32'h00000000} /* (3, 12, 16) {real, imag} */,
  {32'hbf625ed3, 32'h00000000} /* (3, 12, 15) {real, imag} */,
  {32'hbf65f42d, 32'h00000000} /* (3, 12, 14) {real, imag} */,
  {32'hbf284e6e, 32'h00000000} /* (3, 12, 13) {real, imag} */,
  {32'hbed9eeed, 32'h00000000} /* (3, 12, 12) {real, imag} */,
  {32'hbebda857, 32'h00000000} /* (3, 12, 11) {real, imag} */,
  {32'h3ed856e7, 32'h00000000} /* (3, 12, 10) {real, imag} */,
  {32'h3f20e1e6, 32'h00000000} /* (3, 12, 9) {real, imag} */,
  {32'h3f3076cd, 32'h00000000} /* (3, 12, 8) {real, imag} */,
  {32'h3f983ad2, 32'h00000000} /* (3, 12, 7) {real, imag} */,
  {32'h3f8c4da4, 32'h00000000} /* (3, 12, 6) {real, imag} */,
  {32'h3f137cc1, 32'h00000000} /* (3, 12, 5) {real, imag} */,
  {32'h3f0e71e0, 32'h00000000} /* (3, 12, 4) {real, imag} */,
  {32'h3f668870, 32'h00000000} /* (3, 12, 3) {real, imag} */,
  {32'h3f84acf4, 32'h00000000} /* (3, 12, 2) {real, imag} */,
  {32'h3ffe2104, 32'h00000000} /* (3, 12, 1) {real, imag} */,
  {32'h3f6e7e7b, 32'h00000000} /* (3, 12, 0) {real, imag} */,
  {32'h3eb03a78, 32'h00000000} /* (3, 11, 31) {real, imag} */,
  {32'h3f57d6f3, 32'h00000000} /* (3, 11, 30) {real, imag} */,
  {32'h3f6e45f6, 32'h00000000} /* (3, 11, 29) {real, imag} */,
  {32'h3f4b5e80, 32'h00000000} /* (3, 11, 28) {real, imag} */,
  {32'h3f4d080a, 32'h00000000} /* (3, 11, 27) {real, imag} */,
  {32'h3e971e27, 32'h00000000} /* (3, 11, 26) {real, imag} */,
  {32'h3ec944e7, 32'h00000000} /* (3, 11, 25) {real, imag} */,
  {32'h3f202208, 32'h00000000} /* (3, 11, 24) {real, imag} */,
  {32'h3ed664ce, 32'h00000000} /* (3, 11, 23) {real, imag} */,
  {32'h3ee77531, 32'h00000000} /* (3, 11, 22) {real, imag} */,
  {32'h3e8ec91a, 32'h00000000} /* (3, 11, 21) {real, imag} */,
  {32'hbf2fc4ba, 32'h00000000} /* (3, 11, 20) {real, imag} */,
  {32'hbfb2681c, 32'h00000000} /* (3, 11, 19) {real, imag} */,
  {32'hbf88b645, 32'h00000000} /* (3, 11, 18) {real, imag} */,
  {32'hbf09f897, 32'h00000000} /* (3, 11, 17) {real, imag} */,
  {32'hbf2fbb50, 32'h00000000} /* (3, 11, 16) {real, imag} */,
  {32'hbf7c146d, 32'h00000000} /* (3, 11, 15) {real, imag} */,
  {32'hbf3a318a, 32'h00000000} /* (3, 11, 14) {real, imag} */,
  {32'hbf2ffb7d, 32'h00000000} /* (3, 11, 13) {real, imag} */,
  {32'hbf36ae4c, 32'h00000000} /* (3, 11, 12) {real, imag} */,
  {32'hbf001712, 32'h00000000} /* (3, 11, 11) {real, imag} */,
  {32'h3f409206, 32'h00000000} /* (3, 11, 10) {real, imag} */,
  {32'h3fb04868, 32'h00000000} /* (3, 11, 9) {real, imag} */,
  {32'h3f8d2de6, 32'h00000000} /* (3, 11, 8) {real, imag} */,
  {32'h3f99a443, 32'h00000000} /* (3, 11, 7) {real, imag} */,
  {32'h3f6c9936, 32'h00000000} /* (3, 11, 6) {real, imag} */,
  {32'h3f1647fb, 32'h00000000} /* (3, 11, 5) {real, imag} */,
  {32'h3f5f36aa, 32'h00000000} /* (3, 11, 4) {real, imag} */,
  {32'h3f6c75f9, 32'h00000000} /* (3, 11, 3) {real, imag} */,
  {32'h3f110d81, 32'h00000000} /* (3, 11, 2) {real, imag} */,
  {32'h3f5ca9f6, 32'h00000000} /* (3, 11, 1) {real, imag} */,
  {32'h3eec077d, 32'h00000000} /* (3, 11, 0) {real, imag} */,
  {32'hbe885aed, 32'h00000000} /* (3, 10, 31) {real, imag} */,
  {32'hbeafb659, 32'h00000000} /* (3, 10, 30) {real, imag} */,
  {32'hbe1b1277, 32'h00000000} /* (3, 10, 29) {real, imag} */,
  {32'hbe810c85, 32'h00000000} /* (3, 10, 28) {real, imag} */,
  {32'hbe4f6011, 32'h00000000} /* (3, 10, 27) {real, imag} */,
  {32'hbf363a60, 32'h00000000} /* (3, 10, 26) {real, imag} */,
  {32'hbebc32e7, 32'h00000000} /* (3, 10, 25) {real, imag} */,
  {32'hbf4f4194, 32'h00000000} /* (3, 10, 24) {real, imag} */,
  {32'hbf45abb3, 32'h00000000} /* (3, 10, 23) {real, imag} */,
  {32'hbf2bf5dc, 32'h00000000} /* (3, 10, 22) {real, imag} */,
  {32'hbe8d0f86, 32'h00000000} /* (3, 10, 21) {real, imag} */,
  {32'h3bc597d1, 32'h00000000} /* (3, 10, 20) {real, imag} */,
  {32'hbdd908aa, 32'h00000000} /* (3, 10, 19) {real, imag} */,
  {32'h3e20ba17, 32'h00000000} /* (3, 10, 18) {real, imag} */,
  {32'h3f0ba61e, 32'h00000000} /* (3, 10, 17) {real, imag} */,
  {32'h3f297002, 32'h00000000} /* (3, 10, 16) {real, imag} */,
  {32'h3d504264, 32'h00000000} /* (3, 10, 15) {real, imag} */,
  {32'h3dcda627, 32'h00000000} /* (3, 10, 14) {real, imag} */,
  {32'h3baefcd6, 32'h00000000} /* (3, 10, 13) {real, imag} */,
  {32'h3ee81468, 32'h00000000} /* (3, 10, 12) {real, imag} */,
  {32'h3f3fba2b, 32'h00000000} /* (3, 10, 11) {real, imag} */,
  {32'h3ee92bef, 32'h00000000} /* (3, 10, 10) {real, imag} */,
  {32'h3e7114dd, 32'h00000000} /* (3, 10, 9) {real, imag} */,
  {32'hbe31105d, 32'h00000000} /* (3, 10, 8) {real, imag} */,
  {32'hbc73123c, 32'h00000000} /* (3, 10, 7) {real, imag} */,
  {32'hbe844875, 32'h00000000} /* (3, 10, 6) {real, imag} */,
  {32'hbe9596fb, 32'h00000000} /* (3, 10, 5) {real, imag} */,
  {32'hbebe5e10, 32'h00000000} /* (3, 10, 4) {real, imag} */,
  {32'hbf328f7d, 32'h00000000} /* (3, 10, 3) {real, imag} */,
  {32'hbf11256a, 32'h00000000} /* (3, 10, 2) {real, imag} */,
  {32'hbeecf2d9, 32'h00000000} /* (3, 10, 1) {real, imag} */,
  {32'hbf0cfe64, 32'h00000000} /* (3, 10, 0) {real, imag} */,
  {32'hbf20ae67, 32'h00000000} /* (3, 9, 31) {real, imag} */,
  {32'hbf977e4b, 32'h00000000} /* (3, 9, 30) {real, imag} */,
  {32'hbf3df107, 32'h00000000} /* (3, 9, 29) {real, imag} */,
  {32'hbf463285, 32'h00000000} /* (3, 9, 28) {real, imag} */,
  {32'hbf235b4d, 32'h00000000} /* (3, 9, 27) {real, imag} */,
  {32'hbf515027, 32'h00000000} /* (3, 9, 26) {real, imag} */,
  {32'hbea217a7, 32'h00000000} /* (3, 9, 25) {real, imag} */,
  {32'hbf1349dd, 32'h00000000} /* (3, 9, 24) {real, imag} */,
  {32'hbf85c2cd, 32'h00000000} /* (3, 9, 23) {real, imag} */,
  {32'hbf96b01e, 32'h00000000} /* (3, 9, 22) {real, imag} */,
  {32'hbf1624fa, 32'h00000000} /* (3, 9, 21) {real, imag} */,
  {32'h3e760185, 32'h00000000} /* (3, 9, 20) {real, imag} */,
  {32'h3f4fd6af, 32'h00000000} /* (3, 9, 19) {real, imag} */,
  {32'h3f5b8f24, 32'h00000000} /* (3, 9, 18) {real, imag} */,
  {32'h3f7bc234, 32'h00000000} /* (3, 9, 17) {real, imag} */,
  {32'h3f745501, 32'h00000000} /* (3, 9, 16) {real, imag} */,
  {32'h3f4f39d9, 32'h00000000} /* (3, 9, 15) {real, imag} */,
  {32'h3f31a884, 32'h00000000} /* (3, 9, 14) {real, imag} */,
  {32'h3f17a498, 32'h00000000} /* (3, 9, 13) {real, imag} */,
  {32'h3ff279bf, 32'h00000000} /* (3, 9, 12) {real, imag} */,
  {32'h3fa98208, 32'h00000000} /* (3, 9, 11) {real, imag} */,
  {32'hbe10b7c6, 32'h00000000} /* (3, 9, 10) {real, imag} */,
  {32'hbf3fe374, 32'h00000000} /* (3, 9, 9) {real, imag} */,
  {32'hbf52703a, 32'h00000000} /* (3, 9, 8) {real, imag} */,
  {32'hbeabef92, 32'h00000000} /* (3, 9, 7) {real, imag} */,
  {32'hbf58d019, 32'h00000000} /* (3, 9, 6) {real, imag} */,
  {32'hbf513b1d, 32'h00000000} /* (3, 9, 5) {real, imag} */,
  {32'hbf84d52a, 32'h00000000} /* (3, 9, 4) {real, imag} */,
  {32'hbfb29cee, 32'h00000000} /* (3, 9, 3) {real, imag} */,
  {32'hbf8197f2, 32'h00000000} /* (3, 9, 2) {real, imag} */,
  {32'hbf5069d6, 32'h00000000} /* (3, 9, 1) {real, imag} */,
  {32'hbeef61bc, 32'h00000000} /* (3, 9, 0) {real, imag} */,
  {32'hbee8e180, 32'h00000000} /* (3, 8, 31) {real, imag} */,
  {32'hbf517eb7, 32'h00000000} /* (3, 8, 30) {real, imag} */,
  {32'hbf43473e, 32'h00000000} /* (3, 8, 29) {real, imag} */,
  {32'hbf86c033, 32'h00000000} /* (3, 8, 28) {real, imag} */,
  {32'hbf887007, 32'h00000000} /* (3, 8, 27) {real, imag} */,
  {32'hbf9b5c4c, 32'h00000000} /* (3, 8, 26) {real, imag} */,
  {32'hbefced92, 32'h00000000} /* (3, 8, 25) {real, imag} */,
  {32'hbeee849e, 32'h00000000} /* (3, 8, 24) {real, imag} */,
  {32'hbf4b1511, 32'h00000000} /* (3, 8, 23) {real, imag} */,
  {32'hbf1a4bfd, 32'h00000000} /* (3, 8, 22) {real, imag} */,
  {32'hbe116e6f, 32'h00000000} /* (3, 8, 21) {real, imag} */,
  {32'h3efe046f, 32'h00000000} /* (3, 8, 20) {real, imag} */,
  {32'h3f9b2152, 32'h00000000} /* (3, 8, 19) {real, imag} */,
  {32'h3fa14c46, 32'h00000000} /* (3, 8, 18) {real, imag} */,
  {32'h3f47aed5, 32'h00000000} /* (3, 8, 17) {real, imag} */,
  {32'h3f10f0c5, 32'h00000000} /* (3, 8, 16) {real, imag} */,
  {32'h3f76ec37, 32'h00000000} /* (3, 8, 15) {real, imag} */,
  {32'h3f12eadb, 32'h00000000} /* (3, 8, 14) {real, imag} */,
  {32'h3e9481cf, 32'h00000000} /* (3, 8, 13) {real, imag} */,
  {32'h3fbf0953, 32'h00000000} /* (3, 8, 12) {real, imag} */,
  {32'h3f01f608, 32'h00000000} /* (3, 8, 11) {real, imag} */,
  {32'hbfa34e1a, 32'h00000000} /* (3, 8, 10) {real, imag} */,
  {32'hbfcc2afe, 32'h00000000} /* (3, 8, 9) {real, imag} */,
  {32'hbfb0221c, 32'h00000000} /* (3, 8, 8) {real, imag} */,
  {32'hbf2da8b2, 32'h00000000} /* (3, 8, 7) {real, imag} */,
  {32'hbf50a79e, 32'h00000000} /* (3, 8, 6) {real, imag} */,
  {32'hbf4cb72c, 32'h00000000} /* (3, 8, 5) {real, imag} */,
  {32'hbf7ae172, 32'h00000000} /* (3, 8, 4) {real, imag} */,
  {32'hbfaf971d, 32'h00000000} /* (3, 8, 3) {real, imag} */,
  {32'hbf35a026, 32'h00000000} /* (3, 8, 2) {real, imag} */,
  {32'hbf420c12, 32'h00000000} /* (3, 8, 1) {real, imag} */,
  {32'hbede5046, 32'h00000000} /* (3, 8, 0) {real, imag} */,
  {32'hbe728b23, 32'h00000000} /* (3, 7, 31) {real, imag} */,
  {32'hbec7041a, 32'h00000000} /* (3, 7, 30) {real, imag} */,
  {32'hbf81a7f2, 32'h00000000} /* (3, 7, 29) {real, imag} */,
  {32'hbfcb1ef1, 32'h00000000} /* (3, 7, 28) {real, imag} */,
  {32'hbfbfbfe9, 32'h00000000} /* (3, 7, 27) {real, imag} */,
  {32'hbfe4d347, 32'h00000000} /* (3, 7, 26) {real, imag} */,
  {32'hbf59c7b6, 32'h00000000} /* (3, 7, 25) {real, imag} */,
  {32'hbf57713d, 32'h00000000} /* (3, 7, 24) {real, imag} */,
  {32'hbf2b3433, 32'h00000000} /* (3, 7, 23) {real, imag} */,
  {32'hbecf4290, 32'h00000000} /* (3, 7, 22) {real, imag} */,
  {32'hbdd1d626, 32'h00000000} /* (3, 7, 21) {real, imag} */,
  {32'h3f53aa4b, 32'h00000000} /* (3, 7, 20) {real, imag} */,
  {32'h3f51cf0f, 32'h00000000} /* (3, 7, 19) {real, imag} */,
  {32'h3f6a07d4, 32'h00000000} /* (3, 7, 18) {real, imag} */,
  {32'h3fbfe1bc, 32'h00000000} /* (3, 7, 17) {real, imag} */,
  {32'h3f80144d, 32'h00000000} /* (3, 7, 16) {real, imag} */,
  {32'h3f5e7233, 32'h00000000} /* (3, 7, 15) {real, imag} */,
  {32'h3f83dda6, 32'h00000000} /* (3, 7, 14) {real, imag} */,
  {32'h3ed122ac, 32'h00000000} /* (3, 7, 13) {real, imag} */,
  {32'h3f4d7ba7, 32'h00000000} /* (3, 7, 12) {real, imag} */,
  {32'h3eaa9dec, 32'h00000000} /* (3, 7, 11) {real, imag} */,
  {32'hbf8f83d3, 32'h00000000} /* (3, 7, 10) {real, imag} */,
  {32'hbfaa7eca, 32'h00000000} /* (3, 7, 9) {real, imag} */,
  {32'hbf39549b, 32'h00000000} /* (3, 7, 8) {real, imag} */,
  {32'hbf2a2160, 32'h00000000} /* (3, 7, 7) {real, imag} */,
  {32'hbf2a50b7, 32'h00000000} /* (3, 7, 6) {real, imag} */,
  {32'hbf611162, 32'h00000000} /* (3, 7, 5) {real, imag} */,
  {32'hbf928cea, 32'h00000000} /* (3, 7, 4) {real, imag} */,
  {32'hbfcaf2fd, 32'h00000000} /* (3, 7, 3) {real, imag} */,
  {32'hbf5c1865, 32'h00000000} /* (3, 7, 2) {real, imag} */,
  {32'hbf294646, 32'h00000000} /* (3, 7, 1) {real, imag} */,
  {32'hbebd51f8, 32'h00000000} /* (3, 7, 0) {real, imag} */,
  {32'hbe399a5f, 32'h00000000} /* (3, 6, 31) {real, imag} */,
  {32'hbf13efaa, 32'h00000000} /* (3, 6, 30) {real, imag} */,
  {32'hbf89675a, 32'h00000000} /* (3, 6, 29) {real, imag} */,
  {32'hbf9063e8, 32'h00000000} /* (3, 6, 28) {real, imag} */,
  {32'hbfa0e321, 32'h00000000} /* (3, 6, 27) {real, imag} */,
  {32'hbf99cb37, 32'h00000000} /* (3, 6, 26) {real, imag} */,
  {32'hbf7ac5fe, 32'h00000000} /* (3, 6, 25) {real, imag} */,
  {32'hbf6ca345, 32'h00000000} /* (3, 6, 24) {real, imag} */,
  {32'hbef28836, 32'h00000000} /* (3, 6, 23) {real, imag} */,
  {32'hbe73b003, 32'h00000000} /* (3, 6, 22) {real, imag} */,
  {32'hbd263f50, 32'h00000000} /* (3, 6, 21) {real, imag} */,
  {32'h3ed1c54b, 32'h00000000} /* (3, 6, 20) {real, imag} */,
  {32'h3f018ce3, 32'h00000000} /* (3, 6, 19) {real, imag} */,
  {32'h3ee51bcd, 32'h00000000} /* (3, 6, 18) {real, imag} */,
  {32'h3f5d87ef, 32'h00000000} /* (3, 6, 17) {real, imag} */,
  {32'h3f55123f, 32'h00000000} /* (3, 6, 16) {real, imag} */,
  {32'h3f56c404, 32'h00000000} /* (3, 6, 15) {real, imag} */,
  {32'h3f92ace5, 32'h00000000} /* (3, 6, 14) {real, imag} */,
  {32'h3f15a733, 32'h00000000} /* (3, 6, 13) {real, imag} */,
  {32'h3f2b5af0, 32'h00000000} /* (3, 6, 12) {real, imag} */,
  {32'h3f269f4a, 32'h00000000} /* (3, 6, 11) {real, imag} */,
  {32'hbed64160, 32'h00000000} /* (3, 6, 10) {real, imag} */,
  {32'hbf3c2ffb, 32'h00000000} /* (3, 6, 9) {real, imag} */,
  {32'hbee1dd1c, 32'h00000000} /* (3, 6, 8) {real, imag} */,
  {32'hbf0d6f2a, 32'h00000000} /* (3, 6, 7) {real, imag} */,
  {32'hbf9152cd, 32'h00000000} /* (3, 6, 6) {real, imag} */,
  {32'hbf4f0f3a, 32'h00000000} /* (3, 6, 5) {real, imag} */,
  {32'hbf09a878, 32'h00000000} /* (3, 6, 4) {real, imag} */,
  {32'hbf68946e, 32'h00000000} /* (3, 6, 3) {real, imag} */,
  {32'hbfad33c3, 32'h00000000} /* (3, 6, 2) {real, imag} */,
  {32'hbf80cfaa, 32'h00000000} /* (3, 6, 1) {real, imag} */,
  {32'hbee7aa5f, 32'h00000000} /* (3, 6, 0) {real, imag} */,
  {32'hbec9705e, 32'h00000000} /* (3, 5, 31) {real, imag} */,
  {32'hbf24354e, 32'h00000000} /* (3, 5, 30) {real, imag} */,
  {32'hbf67e8d3, 32'h00000000} /* (3, 5, 29) {real, imag} */,
  {32'hbf4f29b4, 32'h00000000} /* (3, 5, 28) {real, imag} */,
  {32'hbf8edfdb, 32'h00000000} /* (3, 5, 27) {real, imag} */,
  {32'hbf97b63d, 32'h00000000} /* (3, 5, 26) {real, imag} */,
  {32'hbfa8a339, 32'h00000000} /* (3, 5, 25) {real, imag} */,
  {32'hbfb0d37a, 32'h00000000} /* (3, 5, 24) {real, imag} */,
  {32'hbf2fc236, 32'h00000000} /* (3, 5, 23) {real, imag} */,
  {32'hbe2bf8df, 32'h00000000} /* (3, 5, 22) {real, imag} */,
  {32'hbd8b8355, 32'h00000000} /* (3, 5, 21) {real, imag} */,
  {32'hbec34d14, 32'h00000000} /* (3, 5, 20) {real, imag} */,
  {32'hbd6132d6, 32'h00000000} /* (3, 5, 19) {real, imag} */,
  {32'hbcff74b0, 32'h00000000} /* (3, 5, 18) {real, imag} */,
  {32'hbe950b70, 32'h00000000} /* (3, 5, 17) {real, imag} */,
  {32'hbd9744cb, 32'h00000000} /* (3, 5, 16) {real, imag} */,
  {32'h3edfb766, 32'h00000000} /* (3, 5, 15) {real, imag} */,
  {32'h3f3bcd1a, 32'h00000000} /* (3, 5, 14) {real, imag} */,
  {32'h3f6f2a83, 32'h00000000} /* (3, 5, 13) {real, imag} */,
  {32'h3f9a0384, 32'h00000000} /* (3, 5, 12) {real, imag} */,
  {32'h3f64a04f, 32'h00000000} /* (3, 5, 11) {real, imag} */,
  {32'h3f618da3, 32'h00000000} /* (3, 5, 10) {real, imag} */,
  {32'h3e2c0cec, 32'h00000000} /* (3, 5, 9) {real, imag} */,
  {32'h3e4d5d35, 32'h00000000} /* (3, 5, 8) {real, imag} */,
  {32'h3ea5f74b, 32'h00000000} /* (3, 5, 7) {real, imag} */,
  {32'hbe089943, 32'h00000000} /* (3, 5, 6) {real, imag} */,
  {32'hbe93eaa5, 32'h00000000} /* (3, 5, 5) {real, imag} */,
  {32'hbf011f81, 32'h00000000} /* (3, 5, 4) {real, imag} */,
  {32'hbf0f72be, 32'h00000000} /* (3, 5, 3) {real, imag} */,
  {32'hbf417fb9, 32'h00000000} /* (3, 5, 2) {real, imag} */,
  {32'hbf2c26c3, 32'h00000000} /* (3, 5, 1) {real, imag} */,
  {32'hbee248bc, 32'h00000000} /* (3, 5, 0) {real, imag} */,
  {32'hbf29e009, 32'h00000000} /* (3, 4, 31) {real, imag} */,
  {32'hbf9d955a, 32'h00000000} /* (3, 4, 30) {real, imag} */,
  {32'hbfc03f56, 32'h00000000} /* (3, 4, 29) {real, imag} */,
  {32'hbfb1afdd, 32'h00000000} /* (3, 4, 28) {real, imag} */,
  {32'hbfb79f9a, 32'h00000000} /* (3, 4, 27) {real, imag} */,
  {32'hbfa1db70, 32'h00000000} /* (3, 4, 26) {real, imag} */,
  {32'hbf7b560e, 32'h00000000} /* (3, 4, 25) {real, imag} */,
  {32'hbf8fc8fa, 32'h00000000} /* (3, 4, 24) {real, imag} */,
  {32'hbf8ce71b, 32'h00000000} /* (3, 4, 23) {real, imag} */,
  {32'hbf15bbcf, 32'h00000000} /* (3, 4, 22) {real, imag} */,
  {32'hbe8e4539, 32'h00000000} /* (3, 4, 21) {real, imag} */,
  {32'hbf278fd6, 32'h00000000} /* (3, 4, 20) {real, imag} */,
  {32'hbf42139f, 32'h00000000} /* (3, 4, 19) {real, imag} */,
  {32'hbf0c51ef, 32'h00000000} /* (3, 4, 18) {real, imag} */,
  {32'hbf13614d, 32'h00000000} /* (3, 4, 17) {real, imag} */,
  {32'hbe608679, 32'h00000000} /* (3, 4, 16) {real, imag} */,
  {32'h3f5b2a50, 32'h00000000} /* (3, 4, 15) {real, imag} */,
  {32'h3f747440, 32'h00000000} /* (3, 4, 14) {real, imag} */,
  {32'h3fa7b9b0, 32'h00000000} /* (3, 4, 13) {real, imag} */,
  {32'h3fa0b30a, 32'h00000000} /* (3, 4, 12) {real, imag} */,
  {32'h3f69db24, 32'h00000000} /* (3, 4, 11) {real, imag} */,
  {32'h3fa35790, 32'h00000000} /* (3, 4, 10) {real, imag} */,
  {32'h3f5ad88c, 32'h00000000} /* (3, 4, 9) {real, imag} */,
  {32'h3f89ed85, 32'h00000000} /* (3, 4, 8) {real, imag} */,
  {32'h3f79ede4, 32'h00000000} /* (3, 4, 7) {real, imag} */,
  {32'h3f8daee2, 32'h00000000} /* (3, 4, 6) {real, imag} */,
  {32'h3ea75905, 32'h00000000} /* (3, 4, 5) {real, imag} */,
  {32'hbea1f5a1, 32'h00000000} /* (3, 4, 4) {real, imag} */,
  {32'hbf08fa5a, 32'h00000000} /* (3, 4, 3) {real, imag} */,
  {32'hbf0704c8, 32'h00000000} /* (3, 4, 2) {real, imag} */,
  {32'hbf360913, 32'h00000000} /* (3, 4, 1) {real, imag} */,
  {32'hbea8474a, 32'h00000000} /* (3, 4, 0) {real, imag} */,
  {32'hbf007524, 32'h00000000} /* (3, 3, 31) {real, imag} */,
  {32'hbfb9fa4e, 32'h00000000} /* (3, 3, 30) {real, imag} */,
  {32'hbfe32a53, 32'h00000000} /* (3, 3, 29) {real, imag} */,
  {32'hbf9d7928, 32'h00000000} /* (3, 3, 28) {real, imag} */,
  {32'hbf892a17, 32'h00000000} /* (3, 3, 27) {real, imag} */,
  {32'hbf6cd324, 32'h00000000} /* (3, 3, 26) {real, imag} */,
  {32'hbf7ee6aa, 32'h00000000} /* (3, 3, 25) {real, imag} */,
  {32'hbf873b17, 32'h00000000} /* (3, 3, 24) {real, imag} */,
  {32'hbf746144, 32'h00000000} /* (3, 3, 23) {real, imag} */,
  {32'hbf570f65, 32'h00000000} /* (3, 3, 22) {real, imag} */,
  {32'hbf21071c, 32'h00000000} /* (3, 3, 21) {real, imag} */,
  {32'hbf606258, 32'h00000000} /* (3, 3, 20) {real, imag} */,
  {32'hbf6e1056, 32'h00000000} /* (3, 3, 19) {real, imag} */,
  {32'hbf600356, 32'h00000000} /* (3, 3, 18) {real, imag} */,
  {32'hbf58dc00, 32'h00000000} /* (3, 3, 17) {real, imag} */,
  {32'hbf526fd7, 32'h00000000} /* (3, 3, 16) {real, imag} */,
  {32'h3f004c20, 32'h00000000} /* (3, 3, 15) {real, imag} */,
  {32'h3f84b046, 32'h00000000} /* (3, 3, 14) {real, imag} */,
  {32'h3fa24a1b, 32'h00000000} /* (3, 3, 13) {real, imag} */,
  {32'h3f97f17d, 32'h00000000} /* (3, 3, 12) {real, imag} */,
  {32'h3f856c38, 32'h00000000} /* (3, 3, 11) {real, imag} */,
  {32'h3fa0f851, 32'h00000000} /* (3, 3, 10) {real, imag} */,
  {32'h3f43fee4, 32'h00000000} /* (3, 3, 9) {real, imag} */,
  {32'h3f491111, 32'h00000000} /* (3, 3, 8) {real, imag} */,
  {32'h3f35cc72, 32'h00000000} /* (3, 3, 7) {real, imag} */,
  {32'h3f8894d8, 32'h00000000} /* (3, 3, 6) {real, imag} */,
  {32'h3d7e7f66, 32'h00000000} /* (3, 3, 5) {real, imag} */,
  {32'hbf097b07, 32'h00000000} /* (3, 3, 4) {real, imag} */,
  {32'hbf7b60a2, 32'h00000000} /* (3, 3, 3) {real, imag} */,
  {32'hbf51913d, 32'h00000000} /* (3, 3, 2) {real, imag} */,
  {32'hbf8063fa, 32'h00000000} /* (3, 3, 1) {real, imag} */,
  {32'hbe92be1c, 32'h00000000} /* (3, 3, 0) {real, imag} */,
  {32'hbee63346, 32'h00000000} /* (3, 2, 31) {real, imag} */,
  {32'hbf95c235, 32'h00000000} /* (3, 2, 30) {real, imag} */,
  {32'hbfb02ed0, 32'h00000000} /* (3, 2, 29) {real, imag} */,
  {32'hbf821bc9, 32'h00000000} /* (3, 2, 28) {real, imag} */,
  {32'hbf7a5712, 32'h00000000} /* (3, 2, 27) {real, imag} */,
  {32'hbf6756b1, 32'h00000000} /* (3, 2, 26) {real, imag} */,
  {32'hbf8b6a3e, 32'h00000000} /* (3, 2, 25) {real, imag} */,
  {32'hbf10df0d, 32'h00000000} /* (3, 2, 24) {real, imag} */,
  {32'hbebc8f03, 32'h00000000} /* (3, 2, 23) {real, imag} */,
  {32'hbf11a240, 32'h00000000} /* (3, 2, 22) {real, imag} */,
  {32'hbf84c1b4, 32'h00000000} /* (3, 2, 21) {real, imag} */,
  {32'hbfc9aa9e, 32'h00000000} /* (3, 2, 20) {real, imag} */,
  {32'hbfa35f5e, 32'h00000000} /* (3, 2, 19) {real, imag} */,
  {32'hbf7aa41b, 32'h00000000} /* (3, 2, 18) {real, imag} */,
  {32'hbf550301, 32'h00000000} /* (3, 2, 17) {real, imag} */,
  {32'hbec5dd31, 32'h00000000} /* (3, 2, 16) {real, imag} */,
  {32'h3f426cea, 32'h00000000} /* (3, 2, 15) {real, imag} */,
  {32'h3f851efd, 32'h00000000} /* (3, 2, 14) {real, imag} */,
  {32'h3f2b2fb6, 32'h00000000} /* (3, 2, 13) {real, imag} */,
  {32'h3f5af4eb, 32'h00000000} /* (3, 2, 12) {real, imag} */,
  {32'h3f872312, 32'h00000000} /* (3, 2, 11) {real, imag} */,
  {32'h3f9312ff, 32'h00000000} /* (3, 2, 10) {real, imag} */,
  {32'h3f8749cb, 32'h00000000} /* (3, 2, 9) {real, imag} */,
  {32'h3f029907, 32'h00000000} /* (3, 2, 8) {real, imag} */,
  {32'h3f4657f0, 32'h00000000} /* (3, 2, 7) {real, imag} */,
  {32'h3f94f4a5, 32'h00000000} /* (3, 2, 6) {real, imag} */,
  {32'hbe04fa1d, 32'h00000000} /* (3, 2, 5) {real, imag} */,
  {32'hbf4d38dc, 32'h00000000} /* (3, 2, 4) {real, imag} */,
  {32'hbf47594e, 32'h00000000} /* (3, 2, 3) {real, imag} */,
  {32'hbf414e96, 32'h00000000} /* (3, 2, 2) {real, imag} */,
  {32'hbf633300, 32'h00000000} /* (3, 2, 1) {real, imag} */,
  {32'hbe9f36a4, 32'h00000000} /* (3, 2, 0) {real, imag} */,
  {32'hbe9c4bd6, 32'h00000000} /* (3, 1, 31) {real, imag} */,
  {32'hbf4cca5a, 32'h00000000} /* (3, 1, 30) {real, imag} */,
  {32'hbf80e2d2, 32'h00000000} /* (3, 1, 29) {real, imag} */,
  {32'hbf381159, 32'h00000000} /* (3, 1, 28) {real, imag} */,
  {32'hbf60e40e, 32'h00000000} /* (3, 1, 27) {real, imag} */,
  {32'hbf6a13c1, 32'h00000000} /* (3, 1, 26) {real, imag} */,
  {32'hbf6f020a, 32'h00000000} /* (3, 1, 25) {real, imag} */,
  {32'hbeffa9c9, 32'h00000000} /* (3, 1, 24) {real, imag} */,
  {32'hbea78cd3, 32'h00000000} /* (3, 1, 23) {real, imag} */,
  {32'hbf15270b, 32'h00000000} /* (3, 1, 22) {real, imag} */,
  {32'hbf940d90, 32'h00000000} /* (3, 1, 21) {real, imag} */,
  {32'hbf894c09, 32'h00000000} /* (3, 1, 20) {real, imag} */,
  {32'hbf4b268a, 32'h00000000} /* (3, 1, 19) {real, imag} */,
  {32'hbf35da64, 32'h00000000} /* (3, 1, 18) {real, imag} */,
  {32'hbf05bfaf, 32'h00000000} /* (3, 1, 17) {real, imag} */,
  {32'hbeb4dc2c, 32'h00000000} /* (3, 1, 16) {real, imag} */,
  {32'h3ed7160b, 32'h00000000} /* (3, 1, 15) {real, imag} */,
  {32'h3f2300d4, 32'h00000000} /* (3, 1, 14) {real, imag} */,
  {32'h3f5ed780, 32'h00000000} /* (3, 1, 13) {real, imag} */,
  {32'h3f5448e2, 32'h00000000} /* (3, 1, 12) {real, imag} */,
  {32'h3f743808, 32'h00000000} /* (3, 1, 11) {real, imag} */,
  {32'h3fa53832, 32'h00000000} /* (3, 1, 10) {real, imag} */,
  {32'h3f892a15, 32'h00000000} /* (3, 1, 9) {real, imag} */,
  {32'h3f3aa894, 32'h00000000} /* (3, 1, 8) {real, imag} */,
  {32'h3fbfbc53, 32'h00000000} /* (3, 1, 7) {real, imag} */,
  {32'h3fed8244, 32'h00000000} /* (3, 1, 6) {real, imag} */,
  {32'h3e0fe784, 32'h00000000} /* (3, 1, 5) {real, imag} */,
  {32'hbf4435cf, 32'h00000000} /* (3, 1, 4) {real, imag} */,
  {32'hbf2c10bc, 32'h00000000} /* (3, 1, 3) {real, imag} */,
  {32'hbf278fcf, 32'h00000000} /* (3, 1, 2) {real, imag} */,
  {32'hbf8cf9a9, 32'h00000000} /* (3, 1, 1) {real, imag} */,
  {32'hbef3c245, 32'h00000000} /* (3, 1, 0) {real, imag} */,
  {32'hbe681f82, 32'h00000000} /* (3, 0, 31) {real, imag} */,
  {32'hbef11048, 32'h00000000} /* (3, 0, 30) {real, imag} */,
  {32'hbf5b6b6d, 32'h00000000} /* (3, 0, 29) {real, imag} */,
  {32'hbf17875a, 32'h00000000} /* (3, 0, 28) {real, imag} */,
  {32'hbe934ac5, 32'h00000000} /* (3, 0, 27) {real, imag} */,
  {32'hbecb4eb0, 32'h00000000} /* (3, 0, 26) {real, imag} */,
  {32'hbef9e2b4, 32'h00000000} /* (3, 0, 25) {real, imag} */,
  {32'hbee5602a, 32'h00000000} /* (3, 0, 24) {real, imag} */,
  {32'hbee51114, 32'h00000000} /* (3, 0, 23) {real, imag} */,
  {32'hbea9dd80, 32'h00000000} /* (3, 0, 22) {real, imag} */,
  {32'hbed1977e, 32'h00000000} /* (3, 0, 21) {real, imag} */,
  {32'hbed1bc53, 32'h00000000} /* (3, 0, 20) {real, imag} */,
  {32'hbead2225, 32'h00000000} /* (3, 0, 19) {real, imag} */,
  {32'hbf03b53f, 32'h00000000} /* (3, 0, 18) {real, imag} */,
  {32'hbed28cff, 32'h00000000} /* (3, 0, 17) {real, imag} */,
  {32'hbe4e62f4, 32'h00000000} /* (3, 0, 16) {real, imag} */,
  {32'h3e200393, 32'h00000000} /* (3, 0, 15) {real, imag} */,
  {32'h3ef405a1, 32'h00000000} /* (3, 0, 14) {real, imag} */,
  {32'h3f6a6cd8, 32'h00000000} /* (3, 0, 13) {real, imag} */,
  {32'h3eef2e88, 32'h00000000} /* (3, 0, 12) {real, imag} */,
  {32'h3ec063d6, 32'h00000000} /* (3, 0, 11) {real, imag} */,
  {32'h3efb0fe2, 32'h00000000} /* (3, 0, 10) {real, imag} */,
  {32'h3f3a9663, 32'h00000000} /* (3, 0, 9) {real, imag} */,
  {32'h3f12a3cb, 32'h00000000} /* (3, 0, 8) {real, imag} */,
  {32'h3f81245b, 32'h00000000} /* (3, 0, 7) {real, imag} */,
  {32'h3fb39eea, 32'h00000000} /* (3, 0, 6) {real, imag} */,
  {32'h3e63ca4d, 32'h00000000} /* (3, 0, 5) {real, imag} */,
  {32'hbeb3e687, 32'h00000000} /* (3, 0, 4) {real, imag} */,
  {32'hbf3d9230, 32'h00000000} /* (3, 0, 3) {real, imag} */,
  {32'hbf132133, 32'h00000000} /* (3, 0, 2) {real, imag} */,
  {32'hbf1d8621, 32'h00000000} /* (3, 0, 1) {real, imag} */,
  {32'hbedac841, 32'h00000000} /* (3, 0, 0) {real, imag} */,
  {32'hbddd0597, 32'h00000000} /* (2, 31, 31) {real, imag} */,
  {32'hbebc60a4, 32'h00000000} /* (2, 31, 30) {real, imag} */,
  {32'hbe8ecdf5, 32'h00000000} /* (2, 31, 29) {real, imag} */,
  {32'hbf1d8d5f, 32'h00000000} /* (2, 31, 28) {real, imag} */,
  {32'hbf3f3de2, 32'h00000000} /* (2, 31, 27) {real, imag} */,
  {32'hbebf22a3, 32'h00000000} /* (2, 31, 26) {real, imag} */,
  {32'hbe9beb75, 32'h00000000} /* (2, 31, 25) {real, imag} */,
  {32'hbed5dc76, 32'h00000000} /* (2, 31, 24) {real, imag} */,
  {32'hbef1b57c, 32'h00000000} /* (2, 31, 23) {real, imag} */,
  {32'hbf03087e, 32'h00000000} /* (2, 31, 22) {real, imag} */,
  {32'hbef3318f, 32'h00000000} /* (2, 31, 21) {real, imag} */,
  {32'h3ecfb4e5, 32'h00000000} /* (2, 31, 20) {real, imag} */,
  {32'h3f15e189, 32'h00000000} /* (2, 31, 19) {real, imag} */,
  {32'h3dc97f18, 32'h00000000} /* (2, 31, 18) {real, imag} */,
  {32'h3e7556aa, 32'h00000000} /* (2, 31, 17) {real, imag} */,
  {32'h3ee62c8f, 32'h00000000} /* (2, 31, 16) {real, imag} */,
  {32'h3f429737, 32'h00000000} /* (2, 31, 15) {real, imag} */,
  {32'h3f72f105, 32'h00000000} /* (2, 31, 14) {real, imag} */,
  {32'h3f3ab9cf, 32'h00000000} /* (2, 31, 13) {real, imag} */,
  {32'h3e8497df, 32'h00000000} /* (2, 31, 12) {real, imag} */,
  {32'h3e7802bc, 32'h00000000} /* (2, 31, 11) {real, imag} */,
  {32'hbebcada9, 32'h00000000} /* (2, 31, 10) {real, imag} */,
  {32'hbf584ea4, 32'h00000000} /* (2, 31, 9) {real, imag} */,
  {32'hbf291ccd, 32'h00000000} /* (2, 31, 8) {real, imag} */,
  {32'hbf63e80a, 32'h00000000} /* (2, 31, 7) {real, imag} */,
  {32'hbf39face, 32'h00000000} /* (2, 31, 6) {real, imag} */,
  {32'hbf1251fb, 32'h00000000} /* (2, 31, 5) {real, imag} */,
  {32'hbe9a1e88, 32'h00000000} /* (2, 31, 4) {real, imag} */,
  {32'hbea657ca, 32'h00000000} /* (2, 31, 3) {real, imag} */,
  {32'hbf868442, 32'h00000000} /* (2, 31, 2) {real, imag} */,
  {32'hbf7312d9, 32'h00000000} /* (2, 31, 1) {real, imag} */,
  {32'hbe200497, 32'h00000000} /* (2, 31, 0) {real, imag} */,
  {32'hbe51e951, 32'h00000000} /* (2, 30, 31) {real, imag} */,
  {32'hbf04fbc4, 32'h00000000} /* (2, 30, 30) {real, imag} */,
  {32'hbee5cd88, 32'h00000000} /* (2, 30, 29) {real, imag} */,
  {32'hbf9d078b, 32'h00000000} /* (2, 30, 28) {real, imag} */,
  {32'hbf872b2f, 32'h00000000} /* (2, 30, 27) {real, imag} */,
  {32'hbf45ddff, 32'h00000000} /* (2, 30, 26) {real, imag} */,
  {32'hbf3e8c61, 32'h00000000} /* (2, 30, 25) {real, imag} */,
  {32'hbf0c470c, 32'h00000000} /* (2, 30, 24) {real, imag} */,
  {32'hbeddb39d, 32'h00000000} /* (2, 30, 23) {real, imag} */,
  {32'hbf867816, 32'h00000000} /* (2, 30, 22) {real, imag} */,
  {32'hbf139eb3, 32'h00000000} /* (2, 30, 21) {real, imag} */,
  {32'h3f806fee, 32'h00000000} /* (2, 30, 20) {real, imag} */,
  {32'h3f9f9d24, 32'h00000000} /* (2, 30, 19) {real, imag} */,
  {32'h3eeaca19, 32'h00000000} /* (2, 30, 18) {real, imag} */,
  {32'h3f25c904, 32'h00000000} /* (2, 30, 17) {real, imag} */,
  {32'h3f67ef7e, 32'h00000000} /* (2, 30, 16) {real, imag} */,
  {32'h3f81fb61, 32'h00000000} /* (2, 30, 15) {real, imag} */,
  {32'h3f86df86, 32'h00000000} /* (2, 30, 14) {real, imag} */,
  {32'h3f50bf48, 32'h00000000} /* (2, 30, 13) {real, imag} */,
  {32'h3f2c715e, 32'h00000000} /* (2, 30, 12) {real, imag} */,
  {32'h3f061ae7, 32'h00000000} /* (2, 30, 11) {real, imag} */,
  {32'hbf336a6e, 32'h00000000} /* (2, 30, 10) {real, imag} */,
  {32'hbf8cfe4c, 32'h00000000} /* (2, 30, 9) {real, imag} */,
  {32'hbf25f879, 32'h00000000} /* (2, 30, 8) {real, imag} */,
  {32'hbf84e020, 32'h00000000} /* (2, 30, 7) {real, imag} */,
  {32'hbf8f2786, 32'h00000000} /* (2, 30, 6) {real, imag} */,
  {32'hbf2ff341, 32'h00000000} /* (2, 30, 5) {real, imag} */,
  {32'hbf6b4308, 32'h00000000} /* (2, 30, 4) {real, imag} */,
  {32'hbf2f4b06, 32'h00000000} /* (2, 30, 3) {real, imag} */,
  {32'hbfd26d4d, 32'h00000000} /* (2, 30, 2) {real, imag} */,
  {32'hbf23f1bf, 32'h00000000} /* (2, 30, 1) {real, imag} */,
  {32'h3d268fb8, 32'h00000000} /* (2, 30, 0) {real, imag} */,
  {32'hbeb49966, 32'h00000000} /* (2, 29, 31) {real, imag} */,
  {32'hbf32d679, 32'h00000000} /* (2, 29, 30) {real, imag} */,
  {32'hbf6a5c25, 32'h00000000} /* (2, 29, 29) {real, imag} */,
  {32'hbf8bb11e, 32'h00000000} /* (2, 29, 28) {real, imag} */,
  {32'hbf99d466, 32'h00000000} /* (2, 29, 27) {real, imag} */,
  {32'hbfaf4902, 32'h00000000} /* (2, 29, 26) {real, imag} */,
  {32'hbf9a4daa, 32'h00000000} /* (2, 29, 25) {real, imag} */,
  {32'hbfaa2374, 32'h00000000} /* (2, 29, 24) {real, imag} */,
  {32'hbf4ca2c2, 32'h00000000} /* (2, 29, 23) {real, imag} */,
  {32'hbfa3a389, 32'h00000000} /* (2, 29, 22) {real, imag} */,
  {32'hbeccab49, 32'h00000000} /* (2, 29, 21) {real, imag} */,
  {32'h3fa64029, 32'h00000000} /* (2, 29, 20) {real, imag} */,
  {32'h3ffc42c9, 32'h00000000} /* (2, 29, 19) {real, imag} */,
  {32'h3fb01c25, 32'h00000000} /* (2, 29, 18) {real, imag} */,
  {32'h3f841081, 32'h00000000} /* (2, 29, 17) {real, imag} */,
  {32'h3f954ba5, 32'h00000000} /* (2, 29, 16) {real, imag} */,
  {32'h3f3db24c, 32'h00000000} /* (2, 29, 15) {real, imag} */,
  {32'h3f224c1e, 32'h00000000} /* (2, 29, 14) {real, imag} */,
  {32'h3f2453fd, 32'h00000000} /* (2, 29, 13) {real, imag} */,
  {32'h3f5ceee9, 32'h00000000} /* (2, 29, 12) {real, imag} */,
  {32'h3efa6c1e, 32'h00000000} /* (2, 29, 11) {real, imag} */,
  {32'hbf4d29c3, 32'h00000000} /* (2, 29, 10) {real, imag} */,
  {32'hbf825dac, 32'h00000000} /* (2, 29, 9) {real, imag} */,
  {32'hbef0b4b9, 32'h00000000} /* (2, 29, 8) {real, imag} */,
  {32'hbf2c239c, 32'h00000000} /* (2, 29, 7) {real, imag} */,
  {32'hbf2e29ec, 32'h00000000} /* (2, 29, 6) {real, imag} */,
  {32'hbf1a9ea3, 32'h00000000} /* (2, 29, 5) {real, imag} */,
  {32'hbfa97eee, 32'h00000000} /* (2, 29, 4) {real, imag} */,
  {32'hbf8dc595, 32'h00000000} /* (2, 29, 3) {real, imag} */,
  {32'hbfa91cd2, 32'h00000000} /* (2, 29, 2) {real, imag} */,
  {32'hbebcc365, 32'h00000000} /* (2, 29, 1) {real, imag} */,
  {32'h3d3a936e, 32'h00000000} /* (2, 29, 0) {real, imag} */,
  {32'hbf04362e, 32'h00000000} /* (2, 28, 31) {real, imag} */,
  {32'hbf5c43e4, 32'h00000000} /* (2, 28, 30) {real, imag} */,
  {32'hbf80b7c5, 32'h00000000} /* (2, 28, 29) {real, imag} */,
  {32'hbf9d8cf2, 32'h00000000} /* (2, 28, 28) {real, imag} */,
  {32'hbfba2e80, 32'h00000000} /* (2, 28, 27) {real, imag} */,
  {32'hbfb21083, 32'h00000000} /* (2, 28, 26) {real, imag} */,
  {32'hbf551b48, 32'h00000000} /* (2, 28, 25) {real, imag} */,
  {32'hbf52a93e, 32'h00000000} /* (2, 28, 24) {real, imag} */,
  {32'hbf8e2124, 32'h00000000} /* (2, 28, 23) {real, imag} */,
  {32'hbfd2b9c8, 32'h00000000} /* (2, 28, 22) {real, imag} */,
  {32'hbef4b110, 32'h00000000} /* (2, 28, 21) {real, imag} */,
  {32'h3fad23b9, 32'h00000000} /* (2, 28, 20) {real, imag} */,
  {32'h3fefcb10, 32'h00000000} /* (2, 28, 19) {real, imag} */,
  {32'h3facd44d, 32'h00000000} /* (2, 28, 18) {real, imag} */,
  {32'h3fa4b82f, 32'h00000000} /* (2, 28, 17) {real, imag} */,
  {32'h3fb597c1, 32'h00000000} /* (2, 28, 16) {real, imag} */,
  {32'h3f29ff9c, 32'h00000000} /* (2, 28, 15) {real, imag} */,
  {32'h3f2863af, 32'h00000000} /* (2, 28, 14) {real, imag} */,
  {32'h3f237e30, 32'h00000000} /* (2, 28, 13) {real, imag} */,
  {32'h3f4ec887, 32'h00000000} /* (2, 28, 12) {real, imag} */,
  {32'h3e98e2cd, 32'h00000000} /* (2, 28, 11) {real, imag} */,
  {32'hbf452266, 32'h00000000} /* (2, 28, 10) {real, imag} */,
  {32'hbfa22863, 32'h00000000} /* (2, 28, 9) {real, imag} */,
  {32'hbf977c08, 32'h00000000} /* (2, 28, 8) {real, imag} */,
  {32'hbfb6343a, 32'h00000000} /* (2, 28, 7) {real, imag} */,
  {32'hbef18784, 32'h00000000} /* (2, 28, 6) {real, imag} */,
  {32'hbf22dfd8, 32'h00000000} /* (2, 28, 5) {real, imag} */,
  {32'hbfa7b71c, 32'h00000000} /* (2, 28, 4) {real, imag} */,
  {32'hbf8f9367, 32'h00000000} /* (2, 28, 3) {real, imag} */,
  {32'hbf69fc55, 32'h00000000} /* (2, 28, 2) {real, imag} */,
  {32'hbead3c00, 32'h00000000} /* (2, 28, 1) {real, imag} */,
  {32'hbe380995, 32'h00000000} /* (2, 28, 0) {real, imag} */,
  {32'hbe3a5713, 32'h00000000} /* (2, 27, 31) {real, imag} */,
  {32'hbf3563dc, 32'h00000000} /* (2, 27, 30) {real, imag} */,
  {32'hbf253617, 32'h00000000} /* (2, 27, 29) {real, imag} */,
  {32'hbf568f4e, 32'h00000000} /* (2, 27, 28) {real, imag} */,
  {32'hbf97eefb, 32'h00000000} /* (2, 27, 27) {real, imag} */,
  {32'hbf8c7a3f, 32'h00000000} /* (2, 27, 26) {real, imag} */,
  {32'hbf5b53e4, 32'h00000000} /* (2, 27, 25) {real, imag} */,
  {32'hbf1abebb, 32'h00000000} /* (2, 27, 24) {real, imag} */,
  {32'hbf795105, 32'h00000000} /* (2, 27, 23) {real, imag} */,
  {32'hbf81c78f, 32'h00000000} /* (2, 27, 22) {real, imag} */,
  {32'hbe9f33ad, 32'h00000000} /* (2, 27, 21) {real, imag} */,
  {32'h3f900d1b, 32'h00000000} /* (2, 27, 20) {real, imag} */,
  {32'h3fcc481d, 32'h00000000} /* (2, 27, 19) {real, imag} */,
  {32'h3f6db61f, 32'h00000000} /* (2, 27, 18) {real, imag} */,
  {32'h3f8a253d, 32'h00000000} /* (2, 27, 17) {real, imag} */,
  {32'h3f76c8e6, 32'h00000000} /* (2, 27, 16) {real, imag} */,
  {32'h3f1bd984, 32'h00000000} /* (2, 27, 15) {real, imag} */,
  {32'h3f40c4f6, 32'h00000000} /* (2, 27, 14) {real, imag} */,
  {32'h3f904998, 32'h00000000} /* (2, 27, 13) {real, imag} */,
  {32'h3f8cf93a, 32'h00000000} /* (2, 27, 12) {real, imag} */,
  {32'h3f35310e, 32'h00000000} /* (2, 27, 11) {real, imag} */,
  {32'hbf0b069c, 32'h00000000} /* (2, 27, 10) {real, imag} */,
  {32'hbf3dd36c, 32'h00000000} /* (2, 27, 9) {real, imag} */,
  {32'hbf347049, 32'h00000000} /* (2, 27, 8) {real, imag} */,
  {32'hbf955ac9, 32'h00000000} /* (2, 27, 7) {real, imag} */,
  {32'hbf77dc20, 32'h00000000} /* (2, 27, 6) {real, imag} */,
  {32'hbf840783, 32'h00000000} /* (2, 27, 5) {real, imag} */,
  {32'hbf53c290, 32'h00000000} /* (2, 27, 4) {real, imag} */,
  {32'hbf8efea3, 32'h00000000} /* (2, 27, 3) {real, imag} */,
  {32'hbfd45487, 32'h00000000} /* (2, 27, 2) {real, imag} */,
  {32'hbf2f490a, 32'h00000000} /* (2, 27, 1) {real, imag} */,
  {32'hbdea2d97, 32'h00000000} /* (2, 27, 0) {real, imag} */,
  {32'hbe99126e, 32'h00000000} /* (2, 26, 31) {real, imag} */,
  {32'hbf3b878c, 32'h00000000} /* (2, 26, 30) {real, imag} */,
  {32'hbf1deb6b, 32'h00000000} /* (2, 26, 29) {real, imag} */,
  {32'hbf6d9f01, 32'h00000000} /* (2, 26, 28) {real, imag} */,
  {32'hbf617c42, 32'h00000000} /* (2, 26, 27) {real, imag} */,
  {32'hbf0547fa, 32'h00000000} /* (2, 26, 26) {real, imag} */,
  {32'hbf59e148, 32'h00000000} /* (2, 26, 25) {real, imag} */,
  {32'hbf568799, 32'h00000000} /* (2, 26, 24) {real, imag} */,
  {32'hbf7779d5, 32'h00000000} /* (2, 26, 23) {real, imag} */,
  {32'hbf360a62, 32'h00000000} /* (2, 26, 22) {real, imag} */,
  {32'h3d8b84f6, 32'h00000000} /* (2, 26, 21) {real, imag} */,
  {32'h3fa3aaa1, 32'h00000000} /* (2, 26, 20) {real, imag} */,
  {32'h3f763db7, 32'h00000000} /* (2, 26, 19) {real, imag} */,
  {32'h3effabef, 32'h00000000} /* (2, 26, 18) {real, imag} */,
  {32'h3f7ab073, 32'h00000000} /* (2, 26, 17) {real, imag} */,
  {32'h3f3c1b59, 32'h00000000} /* (2, 26, 16) {real, imag} */,
  {32'h3f156ab1, 32'h00000000} /* (2, 26, 15) {real, imag} */,
  {32'h3f83aadb, 32'h00000000} /* (2, 26, 14) {real, imag} */,
  {32'h3f8247bc, 32'h00000000} /* (2, 26, 13) {real, imag} */,
  {32'h3fb69e8a, 32'h00000000} /* (2, 26, 12) {real, imag} */,
  {32'h3f77890c, 32'h00000000} /* (2, 26, 11) {real, imag} */,
  {32'h3e0f8e73, 32'h00000000} /* (2, 26, 10) {real, imag} */,
  {32'hbf1a73be, 32'h00000000} /* (2, 26, 9) {real, imag} */,
  {32'hbf00351c, 32'h00000000} /* (2, 26, 8) {real, imag} */,
  {32'hbf13cac6, 32'h00000000} /* (2, 26, 7) {real, imag} */,
  {32'hbf774ff2, 32'h00000000} /* (2, 26, 6) {real, imag} */,
  {32'hbf1e52ea, 32'h00000000} /* (2, 26, 5) {real, imag} */,
  {32'hbe8cd58b, 32'h00000000} /* (2, 26, 4) {real, imag} */,
  {32'hbf43238d, 32'h00000000} /* (2, 26, 3) {real, imag} */,
  {32'hbfb0f7fc, 32'h00000000} /* (2, 26, 2) {real, imag} */,
  {32'hbf6080a5, 32'h00000000} /* (2, 26, 1) {real, imag} */,
  {32'hbe99109b, 32'h00000000} /* (2, 26, 0) {real, imag} */,
  {32'hbf02a2cc, 32'h00000000} /* (2, 25, 31) {real, imag} */,
  {32'hbf687750, 32'h00000000} /* (2, 25, 30) {real, imag} */,
  {32'hbf0d070e, 32'h00000000} /* (2, 25, 29) {real, imag} */,
  {32'hbf3689bd, 32'h00000000} /* (2, 25, 28) {real, imag} */,
  {32'hbf7c1420, 32'h00000000} /* (2, 25, 27) {real, imag} */,
  {32'hbf6a0965, 32'h00000000} /* (2, 25, 26) {real, imag} */,
  {32'hbf9c3166, 32'h00000000} /* (2, 25, 25) {real, imag} */,
  {32'hbf94dc04, 32'h00000000} /* (2, 25, 24) {real, imag} */,
  {32'hbf6ad18e, 32'h00000000} /* (2, 25, 23) {real, imag} */,
  {32'hbf8161d5, 32'h00000000} /* (2, 25, 22) {real, imag} */,
  {32'h3e02a27e, 32'h00000000} /* (2, 25, 21) {real, imag} */,
  {32'h3fa5fc96, 32'h00000000} /* (2, 25, 20) {real, imag} */,
  {32'h3f79a235, 32'h00000000} /* (2, 25, 19) {real, imag} */,
  {32'h3f78345c, 32'h00000000} /* (2, 25, 18) {real, imag} */,
  {32'h3f53d5e4, 32'h00000000} /* (2, 25, 17) {real, imag} */,
  {32'h3f2ea5f1, 32'h00000000} /* (2, 25, 16) {real, imag} */,
  {32'h3f85704b, 32'h00000000} /* (2, 25, 15) {real, imag} */,
  {32'h3f96bcc9, 32'h00000000} /* (2, 25, 14) {real, imag} */,
  {32'h3eff54fc, 32'h00000000} /* (2, 25, 13) {real, imag} */,
  {32'h3f7722cd, 32'h00000000} /* (2, 25, 12) {real, imag} */,
  {32'h3fac3a7a, 32'h00000000} /* (2, 25, 11) {real, imag} */,
  {32'h3e7cd61b, 32'h00000000} /* (2, 25, 10) {real, imag} */,
  {32'hbf731a90, 32'h00000000} /* (2, 25, 9) {real, imag} */,
  {32'hbf57496c, 32'h00000000} /* (2, 25, 8) {real, imag} */,
  {32'hbf720c36, 32'h00000000} /* (2, 25, 7) {real, imag} */,
  {32'hbf9c511a, 32'h00000000} /* (2, 25, 6) {real, imag} */,
  {32'hbf73cb43, 32'h00000000} /* (2, 25, 5) {real, imag} */,
  {32'hbf10176a, 32'h00000000} /* (2, 25, 4) {real, imag} */,
  {32'hbf3e7d21, 32'h00000000} /* (2, 25, 3) {real, imag} */,
  {32'hbf871e93, 32'h00000000} /* (2, 25, 2) {real, imag} */,
  {32'hbf847888, 32'h00000000} /* (2, 25, 1) {real, imag} */,
  {32'hbf5ce8da, 32'h00000000} /* (2, 25, 0) {real, imag} */,
  {32'hbf36c6ba, 32'h00000000} /* (2, 24, 31) {real, imag} */,
  {32'hbf6dcd16, 32'h00000000} /* (2, 24, 30) {real, imag} */,
  {32'hbf0ba9e7, 32'h00000000} /* (2, 24, 29) {real, imag} */,
  {32'hbf15becf, 32'h00000000} /* (2, 24, 28) {real, imag} */,
  {32'hbf69f08a, 32'h00000000} /* (2, 24, 27) {real, imag} */,
  {32'hbfa5a944, 32'h00000000} /* (2, 24, 26) {real, imag} */,
  {32'hbfab305b, 32'h00000000} /* (2, 24, 25) {real, imag} */,
  {32'hbf71e073, 32'h00000000} /* (2, 24, 24) {real, imag} */,
  {32'hbf5e344a, 32'h00000000} /* (2, 24, 23) {real, imag} */,
  {32'hbf8a5a57, 32'h00000000} /* (2, 24, 22) {real, imag} */,
  {32'h3d927eea, 32'h00000000} /* (2, 24, 21) {real, imag} */,
  {32'h3f8cb522, 32'h00000000} /* (2, 24, 20) {real, imag} */,
  {32'h3f6b3626, 32'h00000000} /* (2, 24, 19) {real, imag} */,
  {32'h3fa1cab5, 32'h00000000} /* (2, 24, 18) {real, imag} */,
  {32'h3f954590, 32'h00000000} /* (2, 24, 17) {real, imag} */,
  {32'h3f36b2c7, 32'h00000000} /* (2, 24, 16) {real, imag} */,
  {32'h3f2dca69, 32'h00000000} /* (2, 24, 15) {real, imag} */,
  {32'h3f223ede, 32'h00000000} /* (2, 24, 14) {real, imag} */,
  {32'h3ed4bc68, 32'h00000000} /* (2, 24, 13) {real, imag} */,
  {32'h3f3d1687, 32'h00000000} /* (2, 24, 12) {real, imag} */,
  {32'h3f33d012, 32'h00000000} /* (2, 24, 11) {real, imag} */,
  {32'hbf70a754, 32'h00000000} /* (2, 24, 10) {real, imag} */,
  {32'hbfa09a2e, 32'h00000000} /* (2, 24, 9) {real, imag} */,
  {32'hbef49a90, 32'h00000000} /* (2, 24, 8) {real, imag} */,
  {32'hbf6fbdbc, 32'h00000000} /* (2, 24, 7) {real, imag} */,
  {32'hbf845e89, 32'h00000000} /* (2, 24, 6) {real, imag} */,
  {32'hbf8f22ba, 32'h00000000} /* (2, 24, 5) {real, imag} */,
  {32'hbf487c25, 32'h00000000} /* (2, 24, 4) {real, imag} */,
  {32'hbf838eae, 32'h00000000} /* (2, 24, 3) {real, imag} */,
  {32'hbf9f1ced, 32'h00000000} /* (2, 24, 2) {real, imag} */,
  {32'hbfb6704c, 32'h00000000} /* (2, 24, 1) {real, imag} */,
  {32'hbf62d84e, 32'h00000000} /* (2, 24, 0) {real, imag} */,
  {32'hbf13d308, 32'h00000000} /* (2, 23, 31) {real, imag} */,
  {32'hbf41ee9a, 32'h00000000} /* (2, 23, 30) {real, imag} */,
  {32'hbf85bf1a, 32'h00000000} /* (2, 23, 29) {real, imag} */,
  {32'hbf19d0b8, 32'h00000000} /* (2, 23, 28) {real, imag} */,
  {32'hbf6f6958, 32'h00000000} /* (2, 23, 27) {real, imag} */,
  {32'hbf81acdf, 32'h00000000} /* (2, 23, 26) {real, imag} */,
  {32'hbf67fdce, 32'h00000000} /* (2, 23, 25) {real, imag} */,
  {32'hbf1a83ca, 32'h00000000} /* (2, 23, 24) {real, imag} */,
  {32'hbf0c3651, 32'h00000000} /* (2, 23, 23) {real, imag} */,
  {32'hbf52712e, 32'h00000000} /* (2, 23, 22) {real, imag} */,
  {32'hbecd9025, 32'h00000000} /* (2, 23, 21) {real, imag} */,
  {32'h3f5bc811, 32'h00000000} /* (2, 23, 20) {real, imag} */,
  {32'h3f841c9a, 32'h00000000} /* (2, 23, 19) {real, imag} */,
  {32'h3f8cb76d, 32'h00000000} /* (2, 23, 18) {real, imag} */,
  {32'h3fb7ea9a, 32'h00000000} /* (2, 23, 17) {real, imag} */,
  {32'h3f32274d, 32'h00000000} /* (2, 23, 16) {real, imag} */,
  {32'h3ec217d3, 32'h00000000} /* (2, 23, 15) {real, imag} */,
  {32'h3f3f7c0c, 32'h00000000} /* (2, 23, 14) {real, imag} */,
  {32'h3f3be26e, 32'h00000000} /* (2, 23, 13) {real, imag} */,
  {32'h3f20e17d, 32'h00000000} /* (2, 23, 12) {real, imag} */,
  {32'h3f689808, 32'h00000000} /* (2, 23, 11) {real, imag} */,
  {32'hbeec81af, 32'h00000000} /* (2, 23, 10) {real, imag} */,
  {32'hbf8a69b7, 32'h00000000} /* (2, 23, 9) {real, imag} */,
  {32'hbf3f6506, 32'h00000000} /* (2, 23, 8) {real, imag} */,
  {32'hbf4def88, 32'h00000000} /* (2, 23, 7) {real, imag} */,
  {32'hbefb50c8, 32'h00000000} /* (2, 23, 6) {real, imag} */,
  {32'hbf4397ea, 32'h00000000} /* (2, 23, 5) {real, imag} */,
  {32'hbf296f78, 32'h00000000} /* (2, 23, 4) {real, imag} */,
  {32'hbf52383e, 32'h00000000} /* (2, 23, 3) {real, imag} */,
  {32'hbfa4392d, 32'h00000000} /* (2, 23, 2) {real, imag} */,
  {32'hbfe9186a, 32'h00000000} /* (2, 23, 1) {real, imag} */,
  {32'hbf468c96, 32'h00000000} /* (2, 23, 0) {real, imag} */,
  {32'hbf2904fb, 32'h00000000} /* (2, 22, 31) {real, imag} */,
  {32'hbf531529, 32'h00000000} /* (2, 22, 30) {real, imag} */,
  {32'hbf8add92, 32'h00000000} /* (2, 22, 29) {real, imag} */,
  {32'hbf6b60ad, 32'h00000000} /* (2, 22, 28) {real, imag} */,
  {32'hbf9d2455, 32'h00000000} /* (2, 22, 27) {real, imag} */,
  {32'hbf43a409, 32'h00000000} /* (2, 22, 26) {real, imag} */,
  {32'hbf02ca23, 32'h00000000} /* (2, 22, 25) {real, imag} */,
  {32'hbf49aa84, 32'h00000000} /* (2, 22, 24) {real, imag} */,
  {32'hbef409d6, 32'h00000000} /* (2, 22, 23) {real, imag} */,
  {32'hbf01ade1, 32'h00000000} /* (2, 22, 22) {real, imag} */,
  {32'hbf86e2c9, 32'h00000000} /* (2, 22, 21) {real, imag} */,
  {32'h3ee655e8, 32'h00000000} /* (2, 22, 20) {real, imag} */,
  {32'h3f89eacc, 32'h00000000} /* (2, 22, 19) {real, imag} */,
  {32'h3f57a5e8, 32'h00000000} /* (2, 22, 18) {real, imag} */,
  {32'h3f5cf612, 32'h00000000} /* (2, 22, 17) {real, imag} */,
  {32'h3f5ae373, 32'h00000000} /* (2, 22, 16) {real, imag} */,
  {32'h3f11799a, 32'h00000000} /* (2, 22, 15) {real, imag} */,
  {32'h3faccf93, 32'h00000000} /* (2, 22, 14) {real, imag} */,
  {32'h3fad3b90, 32'h00000000} /* (2, 22, 13) {real, imag} */,
  {32'h3f548274, 32'h00000000} /* (2, 22, 12) {real, imag} */,
  {32'h3efd60ad, 32'h00000000} /* (2, 22, 11) {real, imag} */,
  {32'hbf0fbd52, 32'h00000000} /* (2, 22, 10) {real, imag} */,
  {32'hbf9d1f46, 32'h00000000} /* (2, 22, 9) {real, imag} */,
  {32'hbfbfb10b, 32'h00000000} /* (2, 22, 8) {real, imag} */,
  {32'hbf7d1bf2, 32'h00000000} /* (2, 22, 7) {real, imag} */,
  {32'hbf0cde3e, 32'h00000000} /* (2, 22, 6) {real, imag} */,
  {32'hbf50edef, 32'h00000000} /* (2, 22, 5) {real, imag} */,
  {32'hbf107d0b, 32'h00000000} /* (2, 22, 4) {real, imag} */,
  {32'hbf4b657f, 32'h00000000} /* (2, 22, 3) {real, imag} */,
  {32'hbf889159, 32'h00000000} /* (2, 22, 2) {real, imag} */,
  {32'hbf874e7e, 32'h00000000} /* (2, 22, 1) {real, imag} */,
  {32'hbf5d2ea6, 32'h00000000} /* (2, 22, 0) {real, imag} */,
  {32'hbf23c5e6, 32'h00000000} /* (2, 21, 31) {real, imag} */,
  {32'hbeca3865, 32'h00000000} /* (2, 21, 30) {real, imag} */,
  {32'hbccbb7af, 32'h00000000} /* (2, 21, 29) {real, imag} */,
  {32'hbec7de5e, 32'h00000000} /* (2, 21, 28) {real, imag} */,
  {32'hbf29257d, 32'h00000000} /* (2, 21, 27) {real, imag} */,
  {32'hbe61e10f, 32'h00000000} /* (2, 21, 26) {real, imag} */,
  {32'h3e2b8525, 32'h00000000} /* (2, 21, 25) {real, imag} */,
  {32'hbe6b60da, 32'h00000000} /* (2, 21, 24) {real, imag} */,
  {32'hbe590fde, 32'h00000000} /* (2, 21, 23) {real, imag} */,
  {32'hbedd243e, 32'h00000000} /* (2, 21, 22) {real, imag} */,
  {32'hbf5542ef, 32'h00000000} /* (2, 21, 21) {real, imag} */,
  {32'h3d60c9ab, 32'h00000000} /* (2, 21, 20) {real, imag} */,
  {32'h3efc78f6, 32'h00000000} /* (2, 21, 19) {real, imag} */,
  {32'h3f0e3b0d, 32'h00000000} /* (2, 21, 18) {real, imag} */,
  {32'h3f1073a0, 32'h00000000} /* (2, 21, 17) {real, imag} */,
  {32'h3f5e13e5, 32'h00000000} /* (2, 21, 16) {real, imag} */,
  {32'h3e128dd9, 32'h00000000} /* (2, 21, 15) {real, imag} */,
  {32'h3e8881e3, 32'h00000000} /* (2, 21, 14) {real, imag} */,
  {32'h3ed5a7db, 32'h00000000} /* (2, 21, 13) {real, imag} */,
  {32'h3dd6b792, 32'h00000000} /* (2, 21, 12) {real, imag} */,
  {32'h3ec7ad9c, 32'h00000000} /* (2, 21, 11) {real, imag} */,
  {32'h3dbf990a, 32'h00000000} /* (2, 21, 10) {real, imag} */,
  {32'hbeebd941, 32'h00000000} /* (2, 21, 9) {real, imag} */,
  {32'hbf648176, 32'h00000000} /* (2, 21, 8) {real, imag} */,
  {32'hbedff4be, 32'h00000000} /* (2, 21, 7) {real, imag} */,
  {32'h3c43d2bb, 32'h00000000} /* (2, 21, 6) {real, imag} */,
  {32'hbe6843a3, 32'h00000000} /* (2, 21, 5) {real, imag} */,
  {32'hbf0a7e08, 32'h00000000} /* (2, 21, 4) {real, imag} */,
  {32'hbf2adf4c, 32'h00000000} /* (2, 21, 3) {real, imag} */,
  {32'hbf2c01ec, 32'h00000000} /* (2, 21, 2) {real, imag} */,
  {32'hbf2454ac, 32'h00000000} /* (2, 21, 1) {real, imag} */,
  {32'hbf0e7834, 32'h00000000} /* (2, 21, 0) {real, imag} */,
  {32'h3d923734, 32'h00000000} /* (2, 20, 31) {real, imag} */,
  {32'h3f215db1, 32'h00000000} /* (2, 20, 30) {real, imag} */,
  {32'h3f8d91d5, 32'h00000000} /* (2, 20, 29) {real, imag} */,
  {32'h3fbcbc21, 32'h00000000} /* (2, 20, 28) {real, imag} */,
  {32'h3f8160c7, 32'h00000000} /* (2, 20, 27) {real, imag} */,
  {32'h3eef9fec, 32'h00000000} /* (2, 20, 26) {real, imag} */,
  {32'h3fc493ca, 32'h00000000} /* (2, 20, 25) {real, imag} */,
  {32'h3fa1b60e, 32'h00000000} /* (2, 20, 24) {real, imag} */,
  {32'h3f30ee76, 32'h00000000} /* (2, 20, 23) {real, imag} */,
  {32'h3f2e2bbc, 32'h00000000} /* (2, 20, 22) {real, imag} */,
  {32'h3ce4a8ec, 32'h00000000} /* (2, 20, 21) {real, imag} */,
  {32'hbf31df47, 32'h00000000} /* (2, 20, 20) {real, imag} */,
  {32'hbf15f789, 32'h00000000} /* (2, 20, 19) {real, imag} */,
  {32'hbee5a2c5, 32'h00000000} /* (2, 20, 18) {real, imag} */,
  {32'hbf065767, 32'h00000000} /* (2, 20, 17) {real, imag} */,
  {32'hbe9b722d, 32'h00000000} /* (2, 20, 16) {real, imag} */,
  {32'hbf57068e, 32'h00000000} /* (2, 20, 15) {real, imag} */,
  {32'hbfa2c970, 32'h00000000} /* (2, 20, 14) {real, imag} */,
  {32'hbf659b8b, 32'h00000000} /* (2, 20, 13) {real, imag} */,
  {32'hbf532c38, 32'h00000000} /* (2, 20, 12) {real, imag} */,
  {32'hbf066bac, 32'h00000000} /* (2, 20, 11) {real, imag} */,
  {32'h3e016005, 32'h00000000} /* (2, 20, 10) {real, imag} */,
  {32'h3eef18f7, 32'h00000000} /* (2, 20, 9) {real, imag} */,
  {32'h3d96d417, 32'h00000000} /* (2, 20, 8) {real, imag} */,
  {32'h3efd2a15, 32'h00000000} /* (2, 20, 7) {real, imag} */,
  {32'h3f7fcd43, 32'h00000000} /* (2, 20, 6) {real, imag} */,
  {32'h3f821ac5, 32'h00000000} /* (2, 20, 5) {real, imag} */,
  {32'h3efb15ef, 32'h00000000} /* (2, 20, 4) {real, imag} */,
  {32'h3ecd28a6, 32'h00000000} /* (2, 20, 3) {real, imag} */,
  {32'h3f308f35, 32'h00000000} /* (2, 20, 2) {real, imag} */,
  {32'h3e94d3c1, 32'h00000000} /* (2, 20, 1) {real, imag} */,
  {32'hbd771674, 32'h00000000} /* (2, 20, 0) {real, imag} */,
  {32'h3f20ba3f, 32'h00000000} /* (2, 19, 31) {real, imag} */,
  {32'h3f48c085, 32'h00000000} /* (2, 19, 30) {real, imag} */,
  {32'h3f539792, 32'h00000000} /* (2, 19, 29) {real, imag} */,
  {32'h3fce7f55, 32'h00000000} /* (2, 19, 28) {real, imag} */,
  {32'h3fb17ad9, 32'h00000000} /* (2, 19, 27) {real, imag} */,
  {32'h3f486838, 32'h00000000} /* (2, 19, 26) {real, imag} */,
  {32'h3fbea4b3, 32'h00000000} /* (2, 19, 25) {real, imag} */,
  {32'h3fe0c735, 32'h00000000} /* (2, 19, 24) {real, imag} */,
  {32'h3f8b1b31, 32'h00000000} /* (2, 19, 23) {real, imag} */,
  {32'h3f86bccd, 32'h00000000} /* (2, 19, 22) {real, imag} */,
  {32'h3e1c251d, 32'h00000000} /* (2, 19, 21) {real, imag} */,
  {32'hbf89893e, 32'h00000000} /* (2, 19, 20) {real, imag} */,
  {32'hbf6f2318, 32'h00000000} /* (2, 19, 19) {real, imag} */,
  {32'hbfae0f73, 32'h00000000} /* (2, 19, 18) {real, imag} */,
  {32'hbf817e7d, 32'h00000000} /* (2, 19, 17) {real, imag} */,
  {32'hbf15bcb1, 32'h00000000} /* (2, 19, 16) {real, imag} */,
  {32'hbf5d42d2, 32'h00000000} /* (2, 19, 15) {real, imag} */,
  {32'hbf41a82b, 32'h00000000} /* (2, 19, 14) {real, imag} */,
  {32'hbf4b5775, 32'h00000000} /* (2, 19, 13) {real, imag} */,
  {32'hbf8385e7, 32'h00000000} /* (2, 19, 12) {real, imag} */,
  {32'hbf5432c4, 32'h00000000} /* (2, 19, 11) {real, imag} */,
  {32'h3ef5ba93, 32'h00000000} /* (2, 19, 10) {real, imag} */,
  {32'h3f2a9668, 32'h00000000} /* (2, 19, 9) {real, imag} */,
  {32'h3f1d3cf5, 32'h00000000} /* (2, 19, 8) {real, imag} */,
  {32'h3f74c2f8, 32'h00000000} /* (2, 19, 7) {real, imag} */,
  {32'h3f089b6a, 32'h00000000} /* (2, 19, 6) {real, imag} */,
  {32'h3f39121a, 32'h00000000} /* (2, 19, 5) {real, imag} */,
  {32'h3f3a822c, 32'h00000000} /* (2, 19, 4) {real, imag} */,
  {32'h3f639432, 32'h00000000} /* (2, 19, 3) {real, imag} */,
  {32'h3f8f3e35, 32'h00000000} /* (2, 19, 2) {real, imag} */,
  {32'h3f579f1c, 32'h00000000} /* (2, 19, 1) {real, imag} */,
  {32'h3e933d08, 32'h00000000} /* (2, 19, 0) {real, imag} */,
  {32'h3eb47aa2, 32'h00000000} /* (2, 18, 31) {real, imag} */,
  {32'h3f4d4916, 32'h00000000} /* (2, 18, 30) {real, imag} */,
  {32'h3f3a5de3, 32'h00000000} /* (2, 18, 29) {real, imag} */,
  {32'h3f90a8de, 32'h00000000} /* (2, 18, 28) {real, imag} */,
  {32'h3f962a5d, 32'h00000000} /* (2, 18, 27) {real, imag} */,
  {32'h3fa46dd1, 32'h00000000} /* (2, 18, 26) {real, imag} */,
  {32'h3f9a1293, 32'h00000000} /* (2, 18, 25) {real, imag} */,
  {32'h3f6b16eb, 32'h00000000} /* (2, 18, 24) {real, imag} */,
  {32'h3f226fdd, 32'h00000000} /* (2, 18, 23) {real, imag} */,
  {32'h3f2483f7, 32'h00000000} /* (2, 18, 22) {real, imag} */,
  {32'hbd8d5327, 32'h00000000} /* (2, 18, 21) {real, imag} */,
  {32'hbf976946, 32'h00000000} /* (2, 18, 20) {real, imag} */,
  {32'hbf8bdcdc, 32'h00000000} /* (2, 18, 19) {real, imag} */,
  {32'hbfbe8628, 32'h00000000} /* (2, 18, 18) {real, imag} */,
  {32'hbf9c929c, 32'h00000000} /* (2, 18, 17) {real, imag} */,
  {32'hbf12b45f, 32'h00000000} /* (2, 18, 16) {real, imag} */,
  {32'hbf1bc04c, 32'h00000000} /* (2, 18, 15) {real, imag} */,
  {32'hbf14c1bf, 32'h00000000} /* (2, 18, 14) {real, imag} */,
  {32'hbf496400, 32'h00000000} /* (2, 18, 13) {real, imag} */,
  {32'hbf84ce6e, 32'h00000000} /* (2, 18, 12) {real, imag} */,
  {32'hbf8f6cb1, 32'h00000000} /* (2, 18, 11) {real, imag} */,
  {32'h3e941b46, 32'h00000000} /* (2, 18, 10) {real, imag} */,
  {32'h3f3f93a8, 32'h00000000} /* (2, 18, 9) {real, imag} */,
  {32'h3f7a90bb, 32'h00000000} /* (2, 18, 8) {real, imag} */,
  {32'h3fa09b9c, 32'h00000000} /* (2, 18, 7) {real, imag} */,
  {32'h3ecfb1fa, 32'h00000000} /* (2, 18, 6) {real, imag} */,
  {32'h3eefaa20, 32'h00000000} /* (2, 18, 5) {real, imag} */,
  {32'h3f11550f, 32'h00000000} /* (2, 18, 4) {real, imag} */,
  {32'h3f07f971, 32'h00000000} /* (2, 18, 3) {real, imag} */,
  {32'h3f7b6e53, 32'h00000000} /* (2, 18, 2) {real, imag} */,
  {32'h3f3544b3, 32'h00000000} /* (2, 18, 1) {real, imag} */,
  {32'h3e9e3593, 32'h00000000} /* (2, 18, 0) {real, imag} */,
  {32'h3ef8c06a, 32'h00000000} /* (2, 17, 31) {real, imag} */,
  {32'h3f4be85a, 32'h00000000} /* (2, 17, 30) {real, imag} */,
  {32'h3f61a1df, 32'h00000000} /* (2, 17, 29) {real, imag} */,
  {32'h3f3e1b08, 32'h00000000} /* (2, 17, 28) {real, imag} */,
  {32'h3f4f3c9a, 32'h00000000} /* (2, 17, 27) {real, imag} */,
  {32'h3f67bb1f, 32'h00000000} /* (2, 17, 26) {real, imag} */,
  {32'h3f300788, 32'h00000000} /* (2, 17, 25) {real, imag} */,
  {32'h3eaeaf80, 32'h00000000} /* (2, 17, 24) {real, imag} */,
  {32'h3f65c5b0, 32'h00000000} /* (2, 17, 23) {real, imag} */,
  {32'h3f841914, 32'h00000000} /* (2, 17, 22) {real, imag} */,
  {32'h3dd782c2, 32'h00000000} /* (2, 17, 21) {real, imag} */,
  {32'hbf3b8d4c, 32'h00000000} /* (2, 17, 20) {real, imag} */,
  {32'hbf5eafb3, 32'h00000000} /* (2, 17, 19) {real, imag} */,
  {32'hbf9cb094, 32'h00000000} /* (2, 17, 18) {real, imag} */,
  {32'hbfe9e607, 32'h00000000} /* (2, 17, 17) {real, imag} */,
  {32'hbf990c64, 32'h00000000} /* (2, 17, 16) {real, imag} */,
  {32'hbf18ba58, 32'h00000000} /* (2, 17, 15) {real, imag} */,
  {32'hbf298964, 32'h00000000} /* (2, 17, 14) {real, imag} */,
  {32'hbf46d713, 32'h00000000} /* (2, 17, 13) {real, imag} */,
  {32'hbf00eec9, 32'h00000000} /* (2, 17, 12) {real, imag} */,
  {32'hbf203bfa, 32'h00000000} /* (2, 17, 11) {real, imag} */,
  {32'h3e1e4329, 32'h00000000} /* (2, 17, 10) {real, imag} */,
  {32'h3f3ba54a, 32'h00000000} /* (2, 17, 9) {real, imag} */,
  {32'h3f341188, 32'h00000000} /* (2, 17, 8) {real, imag} */,
  {32'h3f7d4fa5, 32'h00000000} /* (2, 17, 7) {real, imag} */,
  {32'h3faf7f86, 32'h00000000} /* (2, 17, 6) {real, imag} */,
  {32'h3f3b5aee, 32'h00000000} /* (2, 17, 5) {real, imag} */,
  {32'h3ef5802b, 32'h00000000} /* (2, 17, 4) {real, imag} */,
  {32'h3f026e03, 32'h00000000} /* (2, 17, 3) {real, imag} */,
  {32'h3efcda08, 32'h00000000} /* (2, 17, 2) {real, imag} */,
  {32'h3eb64b84, 32'h00000000} /* (2, 17, 1) {real, imag} */,
  {32'h3f0ce834, 32'h00000000} /* (2, 17, 0) {real, imag} */,
  {32'h3f4c9027, 32'h00000000} /* (2, 16, 31) {real, imag} */,
  {32'h3f5ea6ed, 32'h00000000} /* (2, 16, 30) {real, imag} */,
  {32'h3f02fb3e, 32'h00000000} /* (2, 16, 29) {real, imag} */,
  {32'h3eecabbd, 32'h00000000} /* (2, 16, 28) {real, imag} */,
  {32'h3eab40e4, 32'h00000000} /* (2, 16, 27) {real, imag} */,
  {32'h3f1c9240, 32'h00000000} /* (2, 16, 26) {real, imag} */,
  {32'h3f26cdec, 32'h00000000} /* (2, 16, 25) {real, imag} */,
  {32'h3f165fa9, 32'h00000000} /* (2, 16, 24) {real, imag} */,
  {32'h3f73471a, 32'h00000000} /* (2, 16, 23) {real, imag} */,
  {32'h3fa036ef, 32'h00000000} /* (2, 16, 22) {real, imag} */,
  {32'h3ef5ecbe, 32'h00000000} /* (2, 16, 21) {real, imag} */,
  {32'hbf852448, 32'h00000000} /* (2, 16, 20) {real, imag} */,
  {32'hbf8f6369, 32'h00000000} /* (2, 16, 19) {real, imag} */,
  {32'hbf5c50be, 32'h00000000} /* (2, 16, 18) {real, imag} */,
  {32'hbf8e07c4, 32'h00000000} /* (2, 16, 17) {real, imag} */,
  {32'hbf8557b0, 32'h00000000} /* (2, 16, 16) {real, imag} */,
  {32'hbf6777bf, 32'h00000000} /* (2, 16, 15) {real, imag} */,
  {32'hbf178acb, 32'h00000000} /* (2, 16, 14) {real, imag} */,
  {32'hbef7e120, 32'h00000000} /* (2, 16, 13) {real, imag} */,
  {32'hbf0962cc, 32'h00000000} /* (2, 16, 12) {real, imag} */,
  {32'hbf158dba, 32'h00000000} /* (2, 16, 11) {real, imag} */,
  {32'h3ed39c2b, 32'h00000000} /* (2, 16, 10) {real, imag} */,
  {32'h3f57dc8f, 32'h00000000} /* (2, 16, 9) {real, imag} */,
  {32'h3f5623ee, 32'h00000000} /* (2, 16, 8) {real, imag} */,
  {32'h3f790edb, 32'h00000000} /* (2, 16, 7) {real, imag} */,
  {32'h3f83f8f7, 32'h00000000} /* (2, 16, 6) {real, imag} */,
  {32'h3f19a5bf, 32'h00000000} /* (2, 16, 5) {real, imag} */,
  {32'h3ebdcda0, 32'h00000000} /* (2, 16, 4) {real, imag} */,
  {32'h3f8e8b72, 32'h00000000} /* (2, 16, 3) {real, imag} */,
  {32'h3f8d2164, 32'h00000000} /* (2, 16, 2) {real, imag} */,
  {32'h3f2a06f4, 32'h00000000} /* (2, 16, 1) {real, imag} */,
  {32'h3f45276b, 32'h00000000} /* (2, 16, 0) {real, imag} */,
  {32'h3f559b95, 32'h00000000} /* (2, 15, 31) {real, imag} */,
  {32'h3f670022, 32'h00000000} /* (2, 15, 30) {real, imag} */,
  {32'h3f308f59, 32'h00000000} /* (2, 15, 29) {real, imag} */,
  {32'h3f4afbe5, 32'h00000000} /* (2, 15, 28) {real, imag} */,
  {32'h3f037cd3, 32'h00000000} /* (2, 15, 27) {real, imag} */,
  {32'h3f0ed362, 32'h00000000} /* (2, 15, 26) {real, imag} */,
  {32'h3f04cf1e, 32'h00000000} /* (2, 15, 25) {real, imag} */,
  {32'h3f396016, 32'h00000000} /* (2, 15, 24) {real, imag} */,
  {32'h3f204c82, 32'h00000000} /* (2, 15, 23) {real, imag} */,
  {32'h3f7261af, 32'h00000000} /* (2, 15, 22) {real, imag} */,
  {32'h3efc4437, 32'h00000000} /* (2, 15, 21) {real, imag} */,
  {32'hbf446df3, 32'h00000000} /* (2, 15, 20) {real, imag} */,
  {32'hbf3e7721, 32'h00000000} /* (2, 15, 19) {real, imag} */,
  {32'hbef0ec37, 32'h00000000} /* (2, 15, 18) {real, imag} */,
  {32'hbf5375f0, 32'h00000000} /* (2, 15, 17) {real, imag} */,
  {32'hbf329f93, 32'h00000000} /* (2, 15, 16) {real, imag} */,
  {32'hbee36dae, 32'h00000000} /* (2, 15, 15) {real, imag} */,
  {32'hbf1476cd, 32'h00000000} /* (2, 15, 14) {real, imag} */,
  {32'hbf10088d, 32'h00000000} /* (2, 15, 13) {real, imag} */,
  {32'hbf3d7575, 32'h00000000} /* (2, 15, 12) {real, imag} */,
  {32'hbf2641a0, 32'h00000000} /* (2, 15, 11) {real, imag} */,
  {32'h3eaf5c4d, 32'h00000000} /* (2, 15, 10) {real, imag} */,
  {32'h3f3f2cff, 32'h00000000} /* (2, 15, 9) {real, imag} */,
  {32'h3f8acdbd, 32'h00000000} /* (2, 15, 8) {real, imag} */,
  {32'h3f90855a, 32'h00000000} /* (2, 15, 7) {real, imag} */,
  {32'h3ebf168c, 32'h00000000} /* (2, 15, 6) {real, imag} */,
  {32'h3eec1f60, 32'h00000000} /* (2, 15, 5) {real, imag} */,
  {32'h3f3eb45b, 32'h00000000} /* (2, 15, 4) {real, imag} */,
  {32'h3f882690, 32'h00000000} /* (2, 15, 3) {real, imag} */,
  {32'h3fa11eef, 32'h00000000} /* (2, 15, 2) {real, imag} */,
  {32'h3f4bfb1c, 32'h00000000} /* (2, 15, 1) {real, imag} */,
  {32'h3ecd107c, 32'h00000000} /* (2, 15, 0) {real, imag} */,
  {32'h3f52065a, 32'h00000000} /* (2, 14, 31) {real, imag} */,
  {32'h3f9210c8, 32'h00000000} /* (2, 14, 30) {real, imag} */,
  {32'h3f973d4a, 32'h00000000} /* (2, 14, 29) {real, imag} */,
  {32'h3f823193, 32'h00000000} /* (2, 14, 28) {real, imag} */,
  {32'h3f587772, 32'h00000000} /* (2, 14, 27) {real, imag} */,
  {32'h3f6b641a, 32'h00000000} /* (2, 14, 26) {real, imag} */,
  {32'h3f10f414, 32'h00000000} /* (2, 14, 25) {real, imag} */,
  {32'h3f060bd1, 32'h00000000} /* (2, 14, 24) {real, imag} */,
  {32'h3f3220fa, 32'h00000000} /* (2, 14, 23) {real, imag} */,
  {32'h3f86b8a3, 32'h00000000} /* (2, 14, 22) {real, imag} */,
  {32'h3f113f6d, 32'h00000000} /* (2, 14, 21) {real, imag} */,
  {32'hbf0b7491, 32'h00000000} /* (2, 14, 20) {real, imag} */,
  {32'hbf72e9b5, 32'h00000000} /* (2, 14, 19) {real, imag} */,
  {32'hbf3f7595, 32'h00000000} /* (2, 14, 18) {real, imag} */,
  {32'hbf738839, 32'h00000000} /* (2, 14, 17) {real, imag} */,
  {32'hbf81d9b8, 32'h00000000} /* (2, 14, 16) {real, imag} */,
  {32'hbf01c202, 32'h00000000} /* (2, 14, 15) {real, imag} */,
  {32'hbf8062ec, 32'h00000000} /* (2, 14, 14) {real, imag} */,
  {32'hbf813b3a, 32'h00000000} /* (2, 14, 13) {real, imag} */,
  {32'hbf2f35c7, 32'h00000000} /* (2, 14, 12) {real, imag} */,
  {32'hbf0368ab, 32'h00000000} /* (2, 14, 11) {real, imag} */,
  {32'h3f580682, 32'h00000000} /* (2, 14, 10) {real, imag} */,
  {32'h3f9caeef, 32'h00000000} /* (2, 14, 9) {real, imag} */,
  {32'h3fb7af82, 32'h00000000} /* (2, 14, 8) {real, imag} */,
  {32'h3f7a648b, 32'h00000000} /* (2, 14, 7) {real, imag} */,
  {32'h3f0fcb3a, 32'h00000000} /* (2, 14, 6) {real, imag} */,
  {32'h3f322ab4, 32'h00000000} /* (2, 14, 5) {real, imag} */,
  {32'h3f2b7233, 32'h00000000} /* (2, 14, 4) {real, imag} */,
  {32'h3fa8d3e4, 32'h00000000} /* (2, 14, 3) {real, imag} */,
  {32'h3fd0f1ec, 32'h00000000} /* (2, 14, 2) {real, imag} */,
  {32'h3f80f421, 32'h00000000} /* (2, 14, 1) {real, imag} */,
  {32'h3ecfd6d9, 32'h00000000} /* (2, 14, 0) {real, imag} */,
  {32'h3f2517d4, 32'h00000000} /* (2, 13, 31) {real, imag} */,
  {32'h3fc2f24a, 32'h00000000} /* (2, 13, 30) {real, imag} */,
  {32'h4009a759, 32'h00000000} /* (2, 13, 29) {real, imag} */,
  {32'h3fede251, 32'h00000000} /* (2, 13, 28) {real, imag} */,
  {32'h3f78c5ac, 32'h00000000} /* (2, 13, 27) {real, imag} */,
  {32'h3fa048da, 32'h00000000} /* (2, 13, 26) {real, imag} */,
  {32'h3f9010d1, 32'h00000000} /* (2, 13, 25) {real, imag} */,
  {32'h3f8ba350, 32'h00000000} /* (2, 13, 24) {real, imag} */,
  {32'h3fa437f2, 32'h00000000} /* (2, 13, 23) {real, imag} */,
  {32'h3fb19e04, 32'h00000000} /* (2, 13, 22) {real, imag} */,
  {32'h3e96614c, 32'h00000000} /* (2, 13, 21) {real, imag} */,
  {32'hbf41bb39, 32'h00000000} /* (2, 13, 20) {real, imag} */,
  {32'hbf60ea48, 32'h00000000} /* (2, 13, 19) {real, imag} */,
  {32'hbf216a75, 32'h00000000} /* (2, 13, 18) {real, imag} */,
  {32'hbf778196, 32'h00000000} /* (2, 13, 17) {real, imag} */,
  {32'hbf9ffcae, 32'h00000000} /* (2, 13, 16) {real, imag} */,
  {32'hbf2c2af8, 32'h00000000} /* (2, 13, 15) {real, imag} */,
  {32'hbf927f03, 32'h00000000} /* (2, 13, 14) {real, imag} */,
  {32'hbf70b2d4, 32'h00000000} /* (2, 13, 13) {real, imag} */,
  {32'hbf23eeeb, 32'h00000000} /* (2, 13, 12) {real, imag} */,
  {32'hbf273e60, 32'h00000000} /* (2, 13, 11) {real, imag} */,
  {32'h3f147ecf, 32'h00000000} /* (2, 13, 10) {real, imag} */,
  {32'h3f4c7024, 32'h00000000} /* (2, 13, 9) {real, imag} */,
  {32'h3f8101dd, 32'h00000000} /* (2, 13, 8) {real, imag} */,
  {32'h3f615f6b, 32'h00000000} /* (2, 13, 7) {real, imag} */,
  {32'h3f3c255f, 32'h00000000} /* (2, 13, 6) {real, imag} */,
  {32'h3f5cf670, 32'h00000000} /* (2, 13, 5) {real, imag} */,
  {32'h3ec41ca9, 32'h00000000} /* (2, 13, 4) {real, imag} */,
  {32'h3f3de3c9, 32'h00000000} /* (2, 13, 3) {real, imag} */,
  {32'h3f83eea3, 32'h00000000} /* (2, 13, 2) {real, imag} */,
  {32'h3f904861, 32'h00000000} /* (2, 13, 1) {real, imag} */,
  {32'h3f3277c4, 32'h00000000} /* (2, 13, 0) {real, imag} */,
  {32'h3ebf7ac9, 32'h00000000} /* (2, 12, 31) {real, imag} */,
  {32'h3f7d8303, 32'h00000000} /* (2, 12, 30) {real, imag} */,
  {32'h3fc6f69a, 32'h00000000} /* (2, 12, 29) {real, imag} */,
  {32'h3fd53ec7, 32'h00000000} /* (2, 12, 28) {real, imag} */,
  {32'h3f6ffebf, 32'h00000000} /* (2, 12, 27) {real, imag} */,
  {32'h3f1d5865, 32'h00000000} /* (2, 12, 26) {real, imag} */,
  {32'h3f9e9859, 32'h00000000} /* (2, 12, 25) {real, imag} */,
  {32'h3fcfa33a, 32'h00000000} /* (2, 12, 24) {real, imag} */,
  {32'h3fc28a47, 32'h00000000} /* (2, 12, 23) {real, imag} */,
  {32'h3f7efdbc, 32'h00000000} /* (2, 12, 22) {real, imag} */,
  {32'h3d3a7874, 32'h00000000} /* (2, 12, 21) {real, imag} */,
  {32'hbf5e5786, 32'h00000000} /* (2, 12, 20) {real, imag} */,
  {32'hbf53169c, 32'h00000000} /* (2, 12, 19) {real, imag} */,
  {32'hbf33f49a, 32'h00000000} /* (2, 12, 18) {real, imag} */,
  {32'hbf624cb0, 32'h00000000} /* (2, 12, 17) {real, imag} */,
  {32'hbf8873ad, 32'h00000000} /* (2, 12, 16) {real, imag} */,
  {32'hbf8546b1, 32'h00000000} /* (2, 12, 15) {real, imag} */,
  {32'hbf8970c5, 32'h00000000} /* (2, 12, 14) {real, imag} */,
  {32'hbf1bd7e9, 32'h00000000} /* (2, 12, 13) {real, imag} */,
  {32'hbf7e3086, 32'h00000000} /* (2, 12, 12) {real, imag} */,
  {32'hbf805751, 32'h00000000} /* (2, 12, 11) {real, imag} */,
  {32'h3d1e15e3, 32'h00000000} /* (2, 12, 10) {real, imag} */,
  {32'h3f05f787, 32'h00000000} /* (2, 12, 9) {real, imag} */,
  {32'h3f5a3d0a, 32'h00000000} /* (2, 12, 8) {real, imag} */,
  {32'h3f8bd97e, 32'h00000000} /* (2, 12, 7) {real, imag} */,
  {32'h3f87b4c3, 32'h00000000} /* (2, 12, 6) {real, imag} */,
  {32'h3f5aa80f, 32'h00000000} /* (2, 12, 5) {real, imag} */,
  {32'h3f49f748, 32'h00000000} /* (2, 12, 4) {real, imag} */,
  {32'h3f9ee0d6, 32'h00000000} /* (2, 12, 3) {real, imag} */,
  {32'h3fa33949, 32'h00000000} /* (2, 12, 2) {real, imag} */,
  {32'h3fc235c7, 32'h00000000} /* (2, 12, 1) {real, imag} */,
  {32'h3f64ef2d, 32'h00000000} /* (2, 12, 0) {real, imag} */,
  {32'h3f0ac16e, 32'h00000000} /* (2, 11, 31) {real, imag} */,
  {32'h3f50d095, 32'h00000000} /* (2, 11, 30) {real, imag} */,
  {32'h3f84ddab, 32'h00000000} /* (2, 11, 29) {real, imag} */,
  {32'h3f7fddd0, 32'h00000000} /* (2, 11, 28) {real, imag} */,
  {32'h3f2cf944, 32'h00000000} /* (2, 11, 27) {real, imag} */,
  {32'h3e233412, 32'h00000000} /* (2, 11, 26) {real, imag} */,
  {32'h3f268e04, 32'h00000000} /* (2, 11, 25) {real, imag} */,
  {32'h3f5c4019, 32'h00000000} /* (2, 11, 24) {real, imag} */,
  {32'h3f23cd3d, 32'h00000000} /* (2, 11, 23) {real, imag} */,
  {32'h3ecaf722, 32'h00000000} /* (2, 11, 22) {real, imag} */,
  {32'h3e4e0529, 32'h00000000} /* (2, 11, 21) {real, imag} */,
  {32'hbf14fc58, 32'h00000000} /* (2, 11, 20) {real, imag} */,
  {32'hbf53be81, 32'h00000000} /* (2, 11, 19) {real, imag} */,
  {32'hbf3531f1, 32'h00000000} /* (2, 11, 18) {real, imag} */,
  {32'hbf1a5d0b, 32'h00000000} /* (2, 11, 17) {real, imag} */,
  {32'hbf6a000a, 32'h00000000} /* (2, 11, 16) {real, imag} */,
  {32'hbf8a2628, 32'h00000000} /* (2, 11, 15) {real, imag} */,
  {32'hbf83d834, 32'h00000000} /* (2, 11, 14) {real, imag} */,
  {32'hbf6209a6, 32'h00000000} /* (2, 11, 13) {real, imag} */,
  {32'hbfa8befc, 32'h00000000} /* (2, 11, 12) {real, imag} */,
  {32'hbfa9a370, 32'h00000000} /* (2, 11, 11) {real, imag} */,
  {32'hbc5a4f57, 32'h00000000} /* (2, 11, 10) {real, imag} */,
  {32'h3f8a452b, 32'h00000000} /* (2, 11, 9) {real, imag} */,
  {32'h3fa83614, 32'h00000000} /* (2, 11, 8) {real, imag} */,
  {32'h3fb76c8b, 32'h00000000} /* (2, 11, 7) {real, imag} */,
  {32'h3f9ac1c1, 32'h00000000} /* (2, 11, 6) {real, imag} */,
  {32'h3f3bc440, 32'h00000000} /* (2, 11, 5) {real, imag} */,
  {32'h3f915e89, 32'h00000000} /* (2, 11, 4) {real, imag} */,
  {32'h3f735d4c, 32'h00000000} /* (2, 11, 3) {real, imag} */,
  {32'h3ec7c805, 32'h00000000} /* (2, 11, 2) {real, imag} */,
  {32'h3f15bb6e, 32'h00000000} /* (2, 11, 1) {real, imag} */,
  {32'h3f1f9e99, 32'h00000000} /* (2, 11, 0) {real, imag} */,
  {32'hbe9b4fce, 32'h00000000} /* (2, 10, 31) {real, imag} */,
  {32'hbe137655, 32'h00000000} /* (2, 10, 30) {real, imag} */,
  {32'h3e37c7ce, 32'h00000000} /* (2, 10, 29) {real, imag} */,
  {32'hbd7c73de, 32'h00000000} /* (2, 10, 28) {real, imag} */,
  {32'hbdb954ad, 32'h00000000} /* (2, 10, 27) {real, imag} */,
  {32'hbf804766, 32'h00000000} /* (2, 10, 26) {real, imag} */,
  {32'hbf187ef2, 32'h00000000} /* (2, 10, 25) {real, imag} */,
  {32'hbe9db486, 32'h00000000} /* (2, 10, 24) {real, imag} */,
  {32'hbe6ecb99, 32'h00000000} /* (2, 10, 23) {real, imag} */,
  {32'hbeb34dd9, 32'h00000000} /* (2, 10, 22) {real, imag} */,
  {32'hbd8a3e8a, 32'h00000000} /* (2, 10, 21) {real, imag} */,
  {32'h3e87756f, 32'h00000000} /* (2, 10, 20) {real, imag} */,
  {32'h3e30b4d2, 32'h00000000} /* (2, 10, 19) {real, imag} */,
  {32'h3eb59a34, 32'h00000000} /* (2, 10, 18) {real, imag} */,
  {32'h3f12f600, 32'h00000000} /* (2, 10, 17) {real, imag} */,
  {32'h3e9795b7, 32'h00000000} /* (2, 10, 16) {real, imag} */,
  {32'h3e93b331, 32'h00000000} /* (2, 10, 15) {real, imag} */,
  {32'h3e71c246, 32'h00000000} /* (2, 10, 14) {real, imag} */,
  {32'h3eb20f03, 32'h00000000} /* (2, 10, 13) {real, imag} */,
  {32'h3df6064e, 32'h00000000} /* (2, 10, 12) {real, imag} */,
  {32'h3e776215, 32'h00000000} /* (2, 10, 11) {real, imag} */,
  {32'h3e62aafe, 32'h00000000} /* (2, 10, 10) {real, imag} */,
  {32'h3e5486e4, 32'h00000000} /* (2, 10, 9) {real, imag} */,
  {32'hbe35d5a3, 32'h00000000} /* (2, 10, 8) {real, imag} */,
  {32'h3c9637c9, 32'h00000000} /* (2, 10, 7) {real, imag} */,
  {32'hbc4509c4, 32'h00000000} /* (2, 10, 6) {real, imag} */,
  {32'hbe4a2f67, 32'h00000000} /* (2, 10, 5) {real, imag} */,
  {32'hbe891209, 32'h00000000} /* (2, 10, 4) {real, imag} */,
  {32'hbf577b65, 32'h00000000} /* (2, 10, 3) {real, imag} */,
  {32'hbf9a3d8e, 32'h00000000} /* (2, 10, 2) {real, imag} */,
  {32'hbfbb2053, 32'h00000000} /* (2, 10, 1) {real, imag} */,
  {32'hbf42ab62, 32'h00000000} /* (2, 10, 0) {real, imag} */,
  {32'hbf98d168, 32'h00000000} /* (2, 9, 31) {real, imag} */,
  {32'hbf9b375a, 32'h00000000} /* (2, 9, 30) {real, imag} */,
  {32'hbeacc60b, 32'h00000000} /* (2, 9, 29) {real, imag} */,
  {32'hbf0920cd, 32'h00000000} /* (2, 9, 28) {real, imag} */,
  {32'hbf0904e6, 32'h00000000} /* (2, 9, 27) {real, imag} */,
  {32'hbf9a4b45, 32'h00000000} /* (2, 9, 26) {real, imag} */,
  {32'hbf8de3aa, 32'h00000000} /* (2, 9, 25) {real, imag} */,
  {32'hbf502fda, 32'h00000000} /* (2, 9, 24) {real, imag} */,
  {32'hbf3b3e3f, 32'h00000000} /* (2, 9, 23) {real, imag} */,
  {32'hbf9587d4, 32'h00000000} /* (2, 9, 22) {real, imag} */,
  {32'hbf365f9c, 32'h00000000} /* (2, 9, 21) {real, imag} */,
  {32'h3eb89146, 32'h00000000} /* (2, 9, 20) {real, imag} */,
  {32'h3f7d6b0f, 32'h00000000} /* (2, 9, 19) {real, imag} */,
  {32'h3ed2cd1c, 32'h00000000} /* (2, 9, 18) {real, imag} */,
  {32'h3ed2bd52, 32'h00000000} /* (2, 9, 17) {real, imag} */,
  {32'h3f3bfc36, 32'h00000000} /* (2, 9, 16) {real, imag} */,
  {32'h3f950031, 32'h00000000} /* (2, 9, 15) {real, imag} */,
  {32'h3f2ad8f4, 32'h00000000} /* (2, 9, 14) {real, imag} */,
  {32'h3f378934, 32'h00000000} /* (2, 9, 13) {real, imag} */,
  {32'h3f936507, 32'h00000000} /* (2, 9, 12) {real, imag} */,
  {32'h3f8dab9d, 32'h00000000} /* (2, 9, 11) {real, imag} */,
  {32'h3cb95bdd, 32'h00000000} /* (2, 9, 10) {real, imag} */,
  {32'hbeb37a21, 32'h00000000} /* (2, 9, 9) {real, imag} */,
  {32'hbefe1361, 32'h00000000} /* (2, 9, 8) {real, imag} */,
  {32'hbeda81a0, 32'h00000000} /* (2, 9, 7) {real, imag} */,
  {32'hbf373360, 32'h00000000} /* (2, 9, 6) {real, imag} */,
  {32'hbf771a66, 32'h00000000} /* (2, 9, 5) {real, imag} */,
  {32'hbfa143a3, 32'h00000000} /* (2, 9, 4) {real, imag} */,
  {32'hbfeea1cf, 32'h00000000} /* (2, 9, 3) {real, imag} */,
  {32'hbfdf69ab, 32'h00000000} /* (2, 9, 2) {real, imag} */,
  {32'hbf93739e, 32'h00000000} /* (2, 9, 1) {real, imag} */,
  {32'hbf394a2a, 32'h00000000} /* (2, 9, 0) {real, imag} */,
  {32'hbf99f55e, 32'h00000000} /* (2, 8, 31) {real, imag} */,
  {32'hbfc5df6e, 32'h00000000} /* (2, 8, 30) {real, imag} */,
  {32'hbf595677, 32'h00000000} /* (2, 8, 29) {real, imag} */,
  {32'hbf41e6e8, 32'h00000000} /* (2, 8, 28) {real, imag} */,
  {32'hbf3dcadc, 32'h00000000} /* (2, 8, 27) {real, imag} */,
  {32'hbf7b93e9, 32'h00000000} /* (2, 8, 26) {real, imag} */,
  {32'hbf682dbe, 32'h00000000} /* (2, 8, 25) {real, imag} */,
  {32'hbf81f080, 32'h00000000} /* (2, 8, 24) {real, imag} */,
  {32'hbf8bd57d, 32'h00000000} /* (2, 8, 23) {real, imag} */,
  {32'hbf8b9cd6, 32'h00000000} /* (2, 8, 22) {real, imag} */,
  {32'hbf1123bb, 32'h00000000} /* (2, 8, 21) {real, imag} */,
  {32'h3f0250c6, 32'h00000000} /* (2, 8, 20) {real, imag} */,
  {32'h3f9f2b57, 32'h00000000} /* (2, 8, 19) {real, imag} */,
  {32'h3f4ff5bc, 32'h00000000} /* (2, 8, 18) {real, imag} */,
  {32'h3f456bef, 32'h00000000} /* (2, 8, 17) {real, imag} */,
  {32'h3f8569aa, 32'h00000000} /* (2, 8, 16) {real, imag} */,
  {32'h3f6ca024, 32'h00000000} /* (2, 8, 15) {real, imag} */,
  {32'h3f3261d3, 32'h00000000} /* (2, 8, 14) {real, imag} */,
  {32'h3e94e178, 32'h00000000} /* (2, 8, 13) {real, imag} */,
  {32'h3f2bdefa, 32'h00000000} /* (2, 8, 12) {real, imag} */,
  {32'h3eef08dc, 32'h00000000} /* (2, 8, 11) {real, imag} */,
  {32'hbf4b8be5, 32'h00000000} /* (2, 8, 10) {real, imag} */,
  {32'hbfbc14bc, 32'h00000000} /* (2, 8, 9) {real, imag} */,
  {32'hbf8c6288, 32'h00000000} /* (2, 8, 8) {real, imag} */,
  {32'hbf62d2d5, 32'h00000000} /* (2, 8, 7) {real, imag} */,
  {32'hbf538c26, 32'h00000000} /* (2, 8, 6) {real, imag} */,
  {32'hbf583c4c, 32'h00000000} /* (2, 8, 5) {real, imag} */,
  {32'hbf98a6f4, 32'h00000000} /* (2, 8, 4) {real, imag} */,
  {32'hbfcb77dd, 32'h00000000} /* (2, 8, 3) {real, imag} */,
  {32'hbf91ba7a, 32'h00000000} /* (2, 8, 2) {real, imag} */,
  {32'hbf2d408a, 32'h00000000} /* (2, 8, 1) {real, imag} */,
  {32'hbee6c03f, 32'h00000000} /* (2, 8, 0) {real, imag} */,
  {32'hbf020e10, 32'h00000000} /* (2, 7, 31) {real, imag} */,
  {32'hbf7ac502, 32'h00000000} /* (2, 7, 30) {real, imag} */,
  {32'hbfc44e6d, 32'h00000000} /* (2, 7, 29) {real, imag} */,
  {32'hbfb4c86f, 32'h00000000} /* (2, 7, 28) {real, imag} */,
  {32'hbfa3dd8e, 32'h00000000} /* (2, 7, 27) {real, imag} */,
  {32'hbfc8c5d2, 32'h00000000} /* (2, 7, 26) {real, imag} */,
  {32'hbfb59084, 32'h00000000} /* (2, 7, 25) {real, imag} */,
  {32'hbfe4427f, 32'h00000000} /* (2, 7, 24) {real, imag} */,
  {32'hbf90f278, 32'h00000000} /* (2, 7, 23) {real, imag} */,
  {32'hbf311b40, 32'h00000000} /* (2, 7, 22) {real, imag} */,
  {32'hbe64d4a0, 32'h00000000} /* (2, 7, 21) {real, imag} */,
  {32'h3fa0a1e0, 32'h00000000} /* (2, 7, 20) {real, imag} */,
  {32'h3f100dce, 32'h00000000} /* (2, 7, 19) {real, imag} */,
  {32'h3f0068f4, 32'h00000000} /* (2, 7, 18) {real, imag} */,
  {32'h3f8e718b, 32'h00000000} /* (2, 7, 17) {real, imag} */,
  {32'h3f9834c2, 32'h00000000} /* (2, 7, 16) {real, imag} */,
  {32'h3fa588d2, 32'h00000000} /* (2, 7, 15) {real, imag} */,
  {32'h3f94ad9a, 32'h00000000} /* (2, 7, 14) {real, imag} */,
  {32'h3efbd1c3, 32'h00000000} /* (2, 7, 13) {real, imag} */,
  {32'h3f13f8db, 32'h00000000} /* (2, 7, 12) {real, imag} */,
  {32'h3bdc82a3, 32'h00000000} /* (2, 7, 11) {real, imag} */,
  {32'hbf667917, 32'h00000000} /* (2, 7, 10) {real, imag} */,
  {32'hbfb7943e, 32'h00000000} /* (2, 7, 9) {real, imag} */,
  {32'hbf4fb84d, 32'h00000000} /* (2, 7, 8) {real, imag} */,
  {32'hbf88e12c, 32'h00000000} /* (2, 7, 7) {real, imag} */,
  {32'hbf8aa1c7, 32'h00000000} /* (2, 7, 6) {real, imag} */,
  {32'hbf84793d, 32'h00000000} /* (2, 7, 5) {real, imag} */,
  {32'hbfa59981, 32'h00000000} /* (2, 7, 4) {real, imag} */,
  {32'hbfc9c972, 32'h00000000} /* (2, 7, 3) {real, imag} */,
  {32'hbfa4e2be, 32'h00000000} /* (2, 7, 2) {real, imag} */,
  {32'hbfa8b6a4, 32'h00000000} /* (2, 7, 1) {real, imag} */,
  {32'hbf1ab2ed, 32'h00000000} /* (2, 7, 0) {real, imag} */,
  {32'hbecfee39, 32'h00000000} /* (2, 6, 31) {real, imag} */,
  {32'hbf57d248, 32'h00000000} /* (2, 6, 30) {real, imag} */,
  {32'hbf993560, 32'h00000000} /* (2, 6, 29) {real, imag} */,
  {32'hbfb29055, 32'h00000000} /* (2, 6, 28) {real, imag} */,
  {32'hbfd15034, 32'h00000000} /* (2, 6, 27) {real, imag} */,
  {32'hbfcb9018, 32'h00000000} /* (2, 6, 26) {real, imag} */,
  {32'hbfb63858, 32'h00000000} /* (2, 6, 25) {real, imag} */,
  {32'hbfb0ad42, 32'h00000000} /* (2, 6, 24) {real, imag} */,
  {32'hbf343ed6, 32'h00000000} /* (2, 6, 23) {real, imag} */,
  {32'hbecbdf65, 32'h00000000} /* (2, 6, 22) {real, imag} */,
  {32'hbe94a029, 32'h00000000} /* (2, 6, 21) {real, imag} */,
  {32'h3f5e5a4a, 32'h00000000} /* (2, 6, 20) {real, imag} */,
  {32'h3ee869a2, 32'h00000000} /* (2, 6, 19) {real, imag} */,
  {32'h3e149a53, 32'h00000000} /* (2, 6, 18) {real, imag} */,
  {32'h3f320834, 32'h00000000} /* (2, 6, 17) {real, imag} */,
  {32'h3f811a1a, 32'h00000000} /* (2, 6, 16) {real, imag} */,
  {32'h3f701698, 32'h00000000} /* (2, 6, 15) {real, imag} */,
  {32'h3f796391, 32'h00000000} /* (2, 6, 14) {real, imag} */,
  {32'h3f7039f1, 32'h00000000} /* (2, 6, 13) {real, imag} */,
  {32'h3fcbf722, 32'h00000000} /* (2, 6, 12) {real, imag} */,
  {32'h3f721f55, 32'h00000000} /* (2, 6, 11) {real, imag} */,
  {32'hbe566623, 32'h00000000} /* (2, 6, 10) {real, imag} */,
  {32'hbf6e44bd, 32'h00000000} /* (2, 6, 9) {real, imag} */,
  {32'hbf6114ab, 32'h00000000} /* (2, 6, 8) {real, imag} */,
  {32'hbf5b3eed, 32'h00000000} /* (2, 6, 7) {real, imag} */,
  {32'hbf566916, 32'h00000000} /* (2, 6, 6) {real, imag} */,
  {32'hbf442e30, 32'h00000000} /* (2, 6, 5) {real, imag} */,
  {32'hbf388a87, 32'h00000000} /* (2, 6, 4) {real, imag} */,
  {32'hbf6eea8f, 32'h00000000} /* (2, 6, 3) {real, imag} */,
  {32'hbf8f7e86, 32'h00000000} /* (2, 6, 2) {real, imag} */,
  {32'hbf4120a0, 32'h00000000} /* (2, 6, 1) {real, imag} */,
  {32'hbebfb2da, 32'h00000000} /* (2, 6, 0) {real, imag} */,
  {32'hbf834495, 32'h00000000} /* (2, 5, 31) {real, imag} */,
  {32'hbf806007, 32'h00000000} /* (2, 5, 30) {real, imag} */,
  {32'hbf481661, 32'h00000000} /* (2, 5, 29) {real, imag} */,
  {32'hbf50c166, 32'h00000000} /* (2, 5, 28) {real, imag} */,
  {32'hbfa67a7c, 32'h00000000} /* (2, 5, 27) {real, imag} */,
  {32'hbfafce94, 32'h00000000} /* (2, 5, 26) {real, imag} */,
  {32'hbface730, 32'h00000000} /* (2, 5, 25) {real, imag} */,
  {32'hbf90514b, 32'h00000000} /* (2, 5, 24) {real, imag} */,
  {32'hbf51377b, 32'h00000000} /* (2, 5, 23) {real, imag} */,
  {32'hbf18bc6d, 32'h00000000} /* (2, 5, 22) {real, imag} */,
  {32'hbe7ecff0, 32'h00000000} /* (2, 5, 21) {real, imag} */,
  {32'hbcf51120, 32'h00000000} /* (2, 5, 20) {real, imag} */,
  {32'h3d0e3f26, 32'h00000000} /* (2, 5, 19) {real, imag} */,
  {32'hbe792f99, 32'h00000000} /* (2, 5, 18) {real, imag} */,
  {32'hbe9c3611, 32'h00000000} /* (2, 5, 17) {real, imag} */,
  {32'hbf0a43a6, 32'h00000000} /* (2, 5, 16) {real, imag} */,
  {32'h3e58c681, 32'h00000000} /* (2, 5, 15) {real, imag} */,
  {32'h3e68e431, 32'h00000000} /* (2, 5, 14) {real, imag} */,
  {32'h3f861ba4, 32'h00000000} /* (2, 5, 13) {real, imag} */,
  {32'h3ff2afac, 32'h00000000} /* (2, 5, 12) {real, imag} */,
  {32'h3fafa362, 32'h00000000} /* (2, 5, 11) {real, imag} */,
  {32'h3f1d719c, 32'h00000000} /* (2, 5, 10) {real, imag} */,
  {32'h3e6d45a4, 32'h00000000} /* (2, 5, 9) {real, imag} */,
  {32'h3e0e594c, 32'h00000000} /* (2, 5, 8) {real, imag} */,
  {32'hbd12317c, 32'h00000000} /* (2, 5, 7) {real, imag} */,
  {32'hbe13a678, 32'h00000000} /* (2, 5, 6) {real, imag} */,
  {32'hbe905efb, 32'h00000000} /* (2, 5, 5) {real, imag} */,
  {32'hbf5c7b77, 32'h00000000} /* (2, 5, 4) {real, imag} */,
  {32'hbf3b231c, 32'h00000000} /* (2, 5, 3) {real, imag} */,
  {32'hbf1cc6d6, 32'h00000000} /* (2, 5, 2) {real, imag} */,
  {32'hbf0f17cc, 32'h00000000} /* (2, 5, 1) {real, imag} */,
  {32'hbf2864ad, 32'h00000000} /* (2, 5, 0) {real, imag} */,
  {32'hbfa88751, 32'h00000000} /* (2, 4, 31) {real, imag} */,
  {32'hbffff300, 32'h00000000} /* (2, 4, 30) {real, imag} */,
  {32'hbfbae494, 32'h00000000} /* (2, 4, 29) {real, imag} */,
  {32'hbf49c887, 32'h00000000} /* (2, 4, 28) {real, imag} */,
  {32'hbfc2bb5e, 32'h00000000} /* (2, 4, 27) {real, imag} */,
  {32'hbff16eb7, 32'h00000000} /* (2, 4, 26) {real, imag} */,
  {32'hbfc58618, 32'h00000000} /* (2, 4, 25) {real, imag} */,
  {32'hbf9e59fc, 32'h00000000} /* (2, 4, 24) {real, imag} */,
  {32'hbf645996, 32'h00000000} /* (2, 4, 23) {real, imag} */,
  {32'hbf37e70f, 32'h00000000} /* (2, 4, 22) {real, imag} */,
  {32'hbf45c7d2, 32'h00000000} /* (2, 4, 21) {real, imag} */,
  {32'hbf8e8600, 32'h00000000} /* (2, 4, 20) {real, imag} */,
  {32'hbf1b8e91, 32'h00000000} /* (2, 4, 19) {real, imag} */,
  {32'hbedcfcf6, 32'h00000000} /* (2, 4, 18) {real, imag} */,
  {32'hbf5b1b45, 32'h00000000} /* (2, 4, 17) {real, imag} */,
  {32'hbf93699d, 32'h00000000} /* (2, 4, 16) {real, imag} */,
  {32'h3ee0ecd2, 32'h00000000} /* (2, 4, 15) {real, imag} */,
  {32'h3ef3dc1e, 32'h00000000} /* (2, 4, 14) {real, imag} */,
  {32'h3f30aff3, 32'h00000000} /* (2, 4, 13) {real, imag} */,
  {32'h3f8de516, 32'h00000000} /* (2, 4, 12) {real, imag} */,
  {32'h3f9545eb, 32'h00000000} /* (2, 4, 11) {real, imag} */,
  {32'h3fb36dc4, 32'h00000000} /* (2, 4, 10) {real, imag} */,
  {32'h3f96afb8, 32'h00000000} /* (2, 4, 9) {real, imag} */,
  {32'h3f8cde35, 32'h00000000} /* (2, 4, 8) {real, imag} */,
  {32'h3f8f301b, 32'h00000000} /* (2, 4, 7) {real, imag} */,
  {32'h3f7fcf86, 32'h00000000} /* (2, 4, 6) {real, imag} */,
  {32'h3e87cff5, 32'h00000000} /* (2, 4, 5) {real, imag} */,
  {32'hbe9852d7, 32'h00000000} /* (2, 4, 4) {real, imag} */,
  {32'hbf216272, 32'h00000000} /* (2, 4, 3) {real, imag} */,
  {32'hbf29e6c1, 32'h00000000} /* (2, 4, 2) {real, imag} */,
  {32'hbf66ec0a, 32'h00000000} /* (2, 4, 1) {real, imag} */,
  {32'hbf2f863f, 32'h00000000} /* (2, 4, 0) {real, imag} */,
  {32'hbf5322a9, 32'h00000000} /* (2, 3, 31) {real, imag} */,
  {32'hbfe4bd17, 32'h00000000} /* (2, 3, 30) {real, imag} */,
  {32'hbfafe7f3, 32'h00000000} /* (2, 3, 29) {real, imag} */,
  {32'hbf42fc61, 32'h00000000} /* (2, 3, 28) {real, imag} */,
  {32'hbf9e822f, 32'h00000000} /* (2, 3, 27) {real, imag} */,
  {32'hbfa8e9d4, 32'h00000000} /* (2, 3, 26) {real, imag} */,
  {32'hbf9bbf6b, 32'h00000000} /* (2, 3, 25) {real, imag} */,
  {32'hbf8d2fc6, 32'h00000000} /* (2, 3, 24) {real, imag} */,
  {32'hbf64dcd2, 32'h00000000} /* (2, 3, 23) {real, imag} */,
  {32'hbf41000d, 32'h00000000} /* (2, 3, 22) {real, imag} */,
  {32'hbf532769, 32'h00000000} /* (2, 3, 21) {real, imag} */,
  {32'hbf924d14, 32'h00000000} /* (2, 3, 20) {real, imag} */,
  {32'hbf94a1a8, 32'h00000000} /* (2, 3, 19) {real, imag} */,
  {32'hbf212122, 32'h00000000} /* (2, 3, 18) {real, imag} */,
  {32'hbf825656, 32'h00000000} /* (2, 3, 17) {real, imag} */,
  {32'hbf8b813f, 32'h00000000} /* (2, 3, 16) {real, imag} */,
  {32'h3e904def, 32'h00000000} /* (2, 3, 15) {real, imag} */,
  {32'h3f4f1ab4, 32'h00000000} /* (2, 3, 14) {real, imag} */,
  {32'h3f6b0930, 32'h00000000} /* (2, 3, 13) {real, imag} */,
  {32'h3f7819e0, 32'h00000000} /* (2, 3, 12) {real, imag} */,
  {32'h3fb867e3, 32'h00000000} /* (2, 3, 11) {real, imag} */,
  {32'h3faa18e0, 32'h00000000} /* (2, 3, 10) {real, imag} */,
  {32'h3f5ded9d, 32'h00000000} /* (2, 3, 9) {real, imag} */,
  {32'h3f6694cf, 32'h00000000} /* (2, 3, 8) {real, imag} */,
  {32'h3f87bc9f, 32'h00000000} /* (2, 3, 7) {real, imag} */,
  {32'h3f6ddbbd, 32'h00000000} /* (2, 3, 6) {real, imag} */,
  {32'hbedcf660, 32'h00000000} /* (2, 3, 5) {real, imag} */,
  {32'hbf0c5fd6, 32'h00000000} /* (2, 3, 4) {real, imag} */,
  {32'hbf83a0a3, 32'h00000000} /* (2, 3, 3) {real, imag} */,
  {32'hbf4e883d, 32'h00000000} /* (2, 3, 2) {real, imag} */,
  {32'hbf64b10a, 32'h00000000} /* (2, 3, 1) {real, imag} */,
  {32'hbec390a4, 32'h00000000} /* (2, 3, 0) {real, imag} */,
  {32'hbf03e517, 32'h00000000} /* (2, 2, 31) {real, imag} */,
  {32'hbf8d7332, 32'h00000000} /* (2, 2, 30) {real, imag} */,
  {32'hbf960046, 32'h00000000} /* (2, 2, 29) {real, imag} */,
  {32'hbf86aa74, 32'h00000000} /* (2, 2, 28) {real, imag} */,
  {32'hbf772971, 32'h00000000} /* (2, 2, 27) {real, imag} */,
  {32'hbf78faea, 32'h00000000} /* (2, 2, 26) {real, imag} */,
  {32'hbfa3c0fe, 32'h00000000} /* (2, 2, 25) {real, imag} */,
  {32'hbf3c5bb7, 32'h00000000} /* (2, 2, 24) {real, imag} */,
  {32'hbed18532, 32'h00000000} /* (2, 2, 23) {real, imag} */,
  {32'hbf2a1c93, 32'h00000000} /* (2, 2, 22) {real, imag} */,
  {32'hbf9c5cad, 32'h00000000} /* (2, 2, 21) {real, imag} */,
  {32'hbfe09885, 32'h00000000} /* (2, 2, 20) {real, imag} */,
  {32'hbfd5dd2f, 32'h00000000} /* (2, 2, 19) {real, imag} */,
  {32'hbfaa0036, 32'h00000000} /* (2, 2, 18) {real, imag} */,
  {32'hbf9a857a, 32'h00000000} /* (2, 2, 17) {real, imag} */,
  {32'hbed42468, 32'h00000000} /* (2, 2, 16) {real, imag} */,
  {32'h3f444507, 32'h00000000} /* (2, 2, 15) {real, imag} */,
  {32'h3f8b79dc, 32'h00000000} /* (2, 2, 14) {real, imag} */,
  {32'h3faa4f8c, 32'h00000000} /* (2, 2, 13) {real, imag} */,
  {32'h3f89e38f, 32'h00000000} /* (2, 2, 12) {real, imag} */,
  {32'h3fc0aeb3, 32'h00000000} /* (2, 2, 11) {real, imag} */,
  {32'h3f88270d, 32'h00000000} /* (2, 2, 10) {real, imag} */,
  {32'h3fa65808, 32'h00000000} /* (2, 2, 9) {real, imag} */,
  {32'h3f5304e7, 32'h00000000} /* (2, 2, 8) {real, imag} */,
  {32'h3f37b2e3, 32'h00000000} /* (2, 2, 7) {real, imag} */,
  {32'h3f5daef1, 32'h00000000} /* (2, 2, 6) {real, imag} */,
  {32'hbf3344e0, 32'h00000000} /* (2, 2, 5) {real, imag} */,
  {32'hbfb24a20, 32'h00000000} /* (2, 2, 4) {real, imag} */,
  {32'hbfbd9fe9, 32'h00000000} /* (2, 2, 3) {real, imag} */,
  {32'hbf80a4c6, 32'h00000000} /* (2, 2, 2) {real, imag} */,
  {32'hbfbdd15a, 32'h00000000} /* (2, 2, 1) {real, imag} */,
  {32'hbf2ca7a3, 32'h00000000} /* (2, 2, 0) {real, imag} */,
  {32'hbf21263a, 32'h00000000} /* (2, 1, 31) {real, imag} */,
  {32'hbf49864f, 32'h00000000} /* (2, 1, 30) {real, imag} */,
  {32'hbf08c4df, 32'h00000000} /* (2, 1, 29) {real, imag} */,
  {32'hbf11ef55, 32'h00000000} /* (2, 1, 28) {real, imag} */,
  {32'hbf284400, 32'h00000000} /* (2, 1, 27) {real, imag} */,
  {32'hbf7d6c47, 32'h00000000} /* (2, 1, 26) {real, imag} */,
  {32'hbf7d5d2b, 32'h00000000} /* (2, 1, 25) {real, imag} */,
  {32'hbf267287, 32'h00000000} /* (2, 1, 24) {real, imag} */,
  {32'hbf13d70d, 32'h00000000} /* (2, 1, 23) {real, imag} */,
  {32'hbf216f76, 32'h00000000} /* (2, 1, 22) {real, imag} */,
  {32'hbf1181aa, 32'h00000000} /* (2, 1, 21) {real, imag} */,
  {32'hbf734562, 32'h00000000} /* (2, 1, 20) {real, imag} */,
  {32'hbf89f5ac, 32'h00000000} /* (2, 1, 19) {real, imag} */,
  {32'hbf953818, 32'h00000000} /* (2, 1, 18) {real, imag} */,
  {32'hbf081e7c, 32'h00000000} /* (2, 1, 17) {real, imag} */,
  {32'hbc2cb938, 32'h00000000} /* (2, 1, 16) {real, imag} */,
  {32'h3f4bb44b, 32'h00000000} /* (2, 1, 15) {real, imag} */,
  {32'h3f836623, 32'h00000000} /* (2, 1, 14) {real, imag} */,
  {32'h3fb829ef, 32'h00000000} /* (2, 1, 13) {real, imag} */,
  {32'h3fb118d8, 32'h00000000} /* (2, 1, 12) {real, imag} */,
  {32'h3fa5a4b7, 32'h00000000} /* (2, 1, 11) {real, imag} */,
  {32'h3f8eebd4, 32'h00000000} /* (2, 1, 10) {real, imag} */,
  {32'h3fadbff5, 32'h00000000} /* (2, 1, 9) {real, imag} */,
  {32'h3f4fb891, 32'h00000000} /* (2, 1, 8) {real, imag} */,
  {32'h3f793d0d, 32'h00000000} /* (2, 1, 7) {real, imag} */,
  {32'h3fcff82f, 32'h00000000} /* (2, 1, 6) {real, imag} */,
  {32'hbe444621, 32'h00000000} /* (2, 1, 5) {real, imag} */,
  {32'hbfcdea84, 32'h00000000} /* (2, 1, 4) {real, imag} */,
  {32'hbf783fd8, 32'h00000000} /* (2, 1, 3) {real, imag} */,
  {32'hbf32baa7, 32'h00000000} /* (2, 1, 2) {real, imag} */,
  {32'hbfacc5cd, 32'h00000000} /* (2, 1, 1) {real, imag} */,
  {32'hbf627b67, 32'h00000000} /* (2, 1, 0) {real, imag} */,
  {32'hbef3810e, 32'h00000000} /* (2, 0, 31) {real, imag} */,
  {32'hbef106d1, 32'h00000000} /* (2, 0, 30) {real, imag} */,
  {32'hbe7f65e3, 32'h00000000} /* (2, 0, 29) {real, imag} */,
  {32'hbea01f23, 32'h00000000} /* (2, 0, 28) {real, imag} */,
  {32'hbea02d90, 32'h00000000} /* (2, 0, 27) {real, imag} */,
  {32'hbec55ce1, 32'h00000000} /* (2, 0, 26) {real, imag} */,
  {32'hbe9abc3a, 32'h00000000} /* (2, 0, 25) {real, imag} */,
  {32'hbeef27bb, 32'h00000000} /* (2, 0, 24) {real, imag} */,
  {32'hbf6e8272, 32'h00000000} /* (2, 0, 23) {real, imag} */,
  {32'hbf1088c5, 32'h00000000} /* (2, 0, 22) {real, imag} */,
  {32'hbdcafbc3, 32'h00000000} /* (2, 0, 21) {real, imag} */,
  {32'hbe8a6791, 32'h00000000} /* (2, 0, 20) {real, imag} */,
  {32'hbed4c5d2, 32'h00000000} /* (2, 0, 19) {real, imag} */,
  {32'hbf279cf4, 32'h00000000} /* (2, 0, 18) {real, imag} */,
  {32'hbe555775, 32'h00000000} /* (2, 0, 17) {real, imag} */,
  {32'h3dc132d3, 32'h00000000} /* (2, 0, 16) {real, imag} */,
  {32'h3eae41ef, 32'h00000000} /* (2, 0, 15) {real, imag} */,
  {32'h3ed60b3a, 32'h00000000} /* (2, 0, 14) {real, imag} */,
  {32'h3f4897e5, 32'h00000000} /* (2, 0, 13) {real, imag} */,
  {32'h3f2d92ba, 32'h00000000} /* (2, 0, 12) {real, imag} */,
  {32'h3ee903c6, 32'h00000000} /* (2, 0, 11) {real, imag} */,
  {32'h3f143db2, 32'h00000000} /* (2, 0, 10) {real, imag} */,
  {32'h3f048167, 32'h00000000} /* (2, 0, 9) {real, imag} */,
  {32'h3e401266, 32'h00000000} /* (2, 0, 8) {real, imag} */,
  {32'h3f17790b, 32'h00000000} /* (2, 0, 7) {real, imag} */,
  {32'h3fb17966, 32'h00000000} /* (2, 0, 6) {real, imag} */,
  {32'hbce423db, 32'h00000000} /* (2, 0, 5) {real, imag} */,
  {32'hbf4054bd, 32'h00000000} /* (2, 0, 4) {real, imag} */,
  {32'hbf04cd65, 32'h00000000} /* (2, 0, 3) {real, imag} */,
  {32'hbf33ccaa, 32'h00000000} /* (2, 0, 2) {real, imag} */,
  {32'hbf6533d2, 32'h00000000} /* (2, 0, 1) {real, imag} */,
  {32'hbf2b207a, 32'h00000000} /* (2, 0, 0) {real, imag} */,
  {32'hbde9cb0a, 32'h00000000} /* (1, 31, 31) {real, imag} */,
  {32'hbea1742d, 32'h00000000} /* (1, 31, 30) {real, imag} */,
  {32'hbf043706, 32'h00000000} /* (1, 31, 29) {real, imag} */,
  {32'hbf8544bc, 32'h00000000} /* (1, 31, 28) {real, imag} */,
  {32'hbf14604f, 32'h00000000} /* (1, 31, 27) {real, imag} */,
  {32'hbe428e43, 32'h00000000} /* (1, 31, 26) {real, imag} */,
  {32'hbe5ddcfe, 32'h00000000} /* (1, 31, 25) {real, imag} */,
  {32'hbefd87c0, 32'h00000000} /* (1, 31, 24) {real, imag} */,
  {32'hbf33dd45, 32'h00000000} /* (1, 31, 23) {real, imag} */,
  {32'hbf5e7371, 32'h00000000} /* (1, 31, 22) {real, imag} */,
  {32'hbf328160, 32'h00000000} /* (1, 31, 21) {real, imag} */,
  {32'h3e25451c, 32'h00000000} /* (1, 31, 20) {real, imag} */,
  {32'h3ec0414f, 32'h00000000} /* (1, 31, 19) {real, imag} */,
  {32'h3e8a6349, 32'h00000000} /* (1, 31, 18) {real, imag} */,
  {32'h3d04dc18, 32'h00000000} /* (1, 31, 17) {real, imag} */,
  {32'h3ea64f8d, 32'h00000000} /* (1, 31, 16) {real, imag} */,
  {32'h3f22361e, 32'h00000000} /* (1, 31, 15) {real, imag} */,
  {32'h3f4c6b2a, 32'h00000000} /* (1, 31, 14) {real, imag} */,
  {32'h3ece8ee6, 32'h00000000} /* (1, 31, 13) {real, imag} */,
  {32'h3e8761a5, 32'h00000000} /* (1, 31, 12) {real, imag} */,
  {32'h3f08ee42, 32'h00000000} /* (1, 31, 11) {real, imag} */,
  {32'hbd1f43b6, 32'h00000000} /* (1, 31, 10) {real, imag} */,
  {32'hbedbf431, 32'h00000000} /* (1, 31, 9) {real, imag} */,
  {32'hbebc7f13, 32'h00000000} /* (1, 31, 8) {real, imag} */,
  {32'hbf02e25d, 32'h00000000} /* (1, 31, 7) {real, imag} */,
  {32'hbee527a0, 32'h00000000} /* (1, 31, 6) {real, imag} */,
  {32'hbf33b3cf, 32'h00000000} /* (1, 31, 5) {real, imag} */,
  {32'hbef13055, 32'h00000000} /* (1, 31, 4) {real, imag} */,
  {32'hbe58324a, 32'h00000000} /* (1, 31, 3) {real, imag} */,
  {32'hbee19316, 32'h00000000} /* (1, 31, 2) {real, imag} */,
  {32'hbec2f691, 32'h00000000} /* (1, 31, 1) {real, imag} */,
  {32'hbda4b544, 32'h00000000} /* (1, 31, 0) {real, imag} */,
  {32'hbe11dced, 32'h00000000} /* (1, 30, 31) {real, imag} */,
  {32'hbca95de8, 32'h00000000} /* (1, 30, 30) {real, imag} */,
  {32'hbf0d3a0c, 32'h00000000} /* (1, 30, 29) {real, imag} */,
  {32'hbfc1c6b9, 32'h00000000} /* (1, 30, 28) {real, imag} */,
  {32'hbf496583, 32'h00000000} /* (1, 30, 27) {real, imag} */,
  {32'hbeaefc00, 32'h00000000} /* (1, 30, 26) {real, imag} */,
  {32'hbede2305, 32'h00000000} /* (1, 30, 25) {real, imag} */,
  {32'hbeeb2636, 32'h00000000} /* (1, 30, 24) {real, imag} */,
  {32'hbf265953, 32'h00000000} /* (1, 30, 23) {real, imag} */,
  {32'hbf99dbda, 32'h00000000} /* (1, 30, 22) {real, imag} */,
  {32'hbf3f8045, 32'h00000000} /* (1, 30, 21) {real, imag} */,
  {32'h3f293dcc, 32'h00000000} /* (1, 30, 20) {real, imag} */,
  {32'h3eda4fa8, 32'h00000000} /* (1, 30, 19) {real, imag} */,
  {32'h3e8abbfe, 32'h00000000} /* (1, 30, 18) {real, imag} */,
  {32'h3f048b5a, 32'h00000000} /* (1, 30, 17) {real, imag} */,
  {32'h3f89eeb4, 32'h00000000} /* (1, 30, 16) {real, imag} */,
  {32'h3f6c0457, 32'h00000000} /* (1, 30, 15) {real, imag} */,
  {32'h3f3dbd0a, 32'h00000000} /* (1, 30, 14) {real, imag} */,
  {32'h3e98f816, 32'h00000000} /* (1, 30, 13) {real, imag} */,
  {32'h3eb781c7, 32'h00000000} /* (1, 30, 12) {real, imag} */,
  {32'h3f37ae7d, 32'h00000000} /* (1, 30, 11) {real, imag} */,
  {32'hbe45ff25, 32'h00000000} /* (1, 30, 10) {real, imag} */,
  {32'hbf598e16, 32'h00000000} /* (1, 30, 9) {real, imag} */,
  {32'hbf3a5e98, 32'h00000000} /* (1, 30, 8) {real, imag} */,
  {32'hbf75a24e, 32'h00000000} /* (1, 30, 7) {real, imag} */,
  {32'hbf880adc, 32'h00000000} /* (1, 30, 6) {real, imag} */,
  {32'hbf867187, 32'h00000000} /* (1, 30, 5) {real, imag} */,
  {32'hbf8dd41a, 32'h00000000} /* (1, 30, 4) {real, imag} */,
  {32'hbf6b3a3f, 32'h00000000} /* (1, 30, 3) {real, imag} */,
  {32'hbf5c6e55, 32'h00000000} /* (1, 30, 2) {real, imag} */,
  {32'hbe4ee3ee, 32'h00000000} /* (1, 30, 1) {real, imag} */,
  {32'hbe6e7e35, 32'h00000000} /* (1, 30, 0) {real, imag} */,
  {32'hbecf935e, 32'h00000000} /* (1, 29, 31) {real, imag} */,
  {32'hbef7de07, 32'h00000000} /* (1, 29, 30) {real, imag} */,
  {32'hbf7e2995, 32'h00000000} /* (1, 29, 29) {real, imag} */,
  {32'hbf6921e3, 32'h00000000} /* (1, 29, 28) {real, imag} */,
  {32'hbeee04a5, 32'h00000000} /* (1, 29, 27) {real, imag} */,
  {32'hbf30e975, 32'h00000000} /* (1, 29, 26) {real, imag} */,
  {32'hbf2154aa, 32'h00000000} /* (1, 29, 25) {real, imag} */,
  {32'hbf302a92, 32'h00000000} /* (1, 29, 24) {real, imag} */,
  {32'hbf80d7e8, 32'h00000000} /* (1, 29, 23) {real, imag} */,
  {32'hbfb3d5d0, 32'h00000000} /* (1, 29, 22) {real, imag} */,
  {32'hbf0c1896, 32'h00000000} /* (1, 29, 21) {real, imag} */,
  {32'h3f424abc, 32'h00000000} /* (1, 29, 20) {real, imag} */,
  {32'h3f3d6a37, 32'h00000000} /* (1, 29, 19) {real, imag} */,
  {32'h3f17bc92, 32'h00000000} /* (1, 29, 18) {real, imag} */,
  {32'h3f4f30c8, 32'h00000000} /* (1, 29, 17) {real, imag} */,
  {32'h3f85c062, 32'h00000000} /* (1, 29, 16) {real, imag} */,
  {32'h3f5a9431, 32'h00000000} /* (1, 29, 15) {real, imag} */,
  {32'h3f81a4d5, 32'h00000000} /* (1, 29, 14) {real, imag} */,
  {32'h3f321e8e, 32'h00000000} /* (1, 29, 13) {real, imag} */,
  {32'h3f1e9b61, 32'h00000000} /* (1, 29, 12) {real, imag} */,
  {32'h3f024637, 32'h00000000} /* (1, 29, 11) {real, imag} */,
  {32'hbf3add88, 32'h00000000} /* (1, 29, 10) {real, imag} */,
  {32'hbfa1ace3, 32'h00000000} /* (1, 29, 9) {real, imag} */,
  {32'hbf7905ab, 32'h00000000} /* (1, 29, 8) {real, imag} */,
  {32'hbf62fbff, 32'h00000000} /* (1, 29, 7) {real, imag} */,
  {32'hbf787b04, 32'h00000000} /* (1, 29, 6) {real, imag} */,
  {32'hbfb89292, 32'h00000000} /* (1, 29, 5) {real, imag} */,
  {32'hbfed08ee, 32'h00000000} /* (1, 29, 4) {real, imag} */,
  {32'hbfac2541, 32'h00000000} /* (1, 29, 3) {real, imag} */,
  {32'hbf808057, 32'h00000000} /* (1, 29, 2) {real, imag} */,
  {32'hbeeca358, 32'h00000000} /* (1, 29, 1) {real, imag} */,
  {32'hbec7f02f, 32'h00000000} /* (1, 29, 0) {real, imag} */,
  {32'hbf24fa8e, 32'h00000000} /* (1, 28, 31) {real, imag} */,
  {32'hbf97238b, 32'h00000000} /* (1, 28, 30) {real, imag} */,
  {32'hbfbdc968, 32'h00000000} /* (1, 28, 29) {real, imag} */,
  {32'hbf40dfb8, 32'h00000000} /* (1, 28, 28) {real, imag} */,
  {32'hbf03eb2c, 32'h00000000} /* (1, 28, 27) {real, imag} */,
  {32'hbf8836b5, 32'h00000000} /* (1, 28, 26) {real, imag} */,
  {32'hbf5a518c, 32'h00000000} /* (1, 28, 25) {real, imag} */,
  {32'hbf2a907f, 32'h00000000} /* (1, 28, 24) {real, imag} */,
  {32'hbf8c2b6d, 32'h00000000} /* (1, 28, 23) {real, imag} */,
  {32'hbfa6a922, 32'h00000000} /* (1, 28, 22) {real, imag} */,
  {32'hbf199133, 32'h00000000} /* (1, 28, 21) {real, imag} */,
  {32'h3f6c85ab, 32'h00000000} /* (1, 28, 20) {real, imag} */,
  {32'h3fb27abb, 32'h00000000} /* (1, 28, 19) {real, imag} */,
  {32'h3f64eebe, 32'h00000000} /* (1, 28, 18) {real, imag} */,
  {32'h3f3bda4b, 32'h00000000} /* (1, 28, 17) {real, imag} */,
  {32'h3f4ff6f7, 32'h00000000} /* (1, 28, 16) {real, imag} */,
  {32'h3f18e216, 32'h00000000} /* (1, 28, 15) {real, imag} */,
  {32'h3f32b293, 32'h00000000} /* (1, 28, 14) {real, imag} */,
  {32'h3f43c5e8, 32'h00000000} /* (1, 28, 13) {real, imag} */,
  {32'h3f781f25, 32'h00000000} /* (1, 28, 12) {real, imag} */,
  {32'h3f0996d1, 32'h00000000} /* (1, 28, 11) {real, imag} */,
  {32'hbf367a0a, 32'h00000000} /* (1, 28, 10) {real, imag} */,
  {32'hbf743c60, 32'h00000000} /* (1, 28, 9) {real, imag} */,
  {32'hbf6f6128, 32'h00000000} /* (1, 28, 8) {real, imag} */,
  {32'hbf93ce55, 32'h00000000} /* (1, 28, 7) {real, imag} */,
  {32'hbf27a568, 32'h00000000} /* (1, 28, 6) {real, imag} */,
  {32'hbf78b85f, 32'h00000000} /* (1, 28, 5) {real, imag} */,
  {32'hbf93741f, 32'h00000000} /* (1, 28, 4) {real, imag} */,
  {32'hbf61a221, 32'h00000000} /* (1, 28, 3) {real, imag} */,
  {32'hbf36b718, 32'h00000000} /* (1, 28, 2) {real, imag} */,
  {32'hbf2081f8, 32'h00000000} /* (1, 28, 1) {real, imag} */,
  {32'hbf2c99f7, 32'h00000000} /* (1, 28, 0) {real, imag} */,
  {32'hbe8a62e7, 32'h00000000} /* (1, 27, 31) {real, imag} */,
  {32'hbfa8250a, 32'h00000000} /* (1, 27, 30) {real, imag} */,
  {32'hbfe560b0, 32'h00000000} /* (1, 27, 29) {real, imag} */,
  {32'hbf8f2f3a, 32'h00000000} /* (1, 27, 28) {real, imag} */,
  {32'hbeecaf05, 32'h00000000} /* (1, 27, 27) {real, imag} */,
  {32'hbefddf8c, 32'h00000000} /* (1, 27, 26) {real, imag} */,
  {32'hbf41dbbc, 32'h00000000} /* (1, 27, 25) {real, imag} */,
  {32'hbf0f8ce2, 32'h00000000} /* (1, 27, 24) {real, imag} */,
  {32'hbf8c680d, 32'h00000000} /* (1, 27, 23) {real, imag} */,
  {32'hbf57433c, 32'h00000000} /* (1, 27, 22) {real, imag} */,
  {32'hbe75644a, 32'h00000000} /* (1, 27, 21) {real, imag} */,
  {32'h3f90d143, 32'h00000000} /* (1, 27, 20) {real, imag} */,
  {32'h3fb865e7, 32'h00000000} /* (1, 27, 19) {real, imag} */,
  {32'h3f7a8b87, 32'h00000000} /* (1, 27, 18) {real, imag} */,
  {32'h3f62fce9, 32'h00000000} /* (1, 27, 17) {real, imag} */,
  {32'h3f3882b0, 32'h00000000} /* (1, 27, 16) {real, imag} */,
  {32'h3f1cf993, 32'h00000000} /* (1, 27, 15) {real, imag} */,
  {32'h3f303df1, 32'h00000000} /* (1, 27, 14) {real, imag} */,
  {32'h3f3b0829, 32'h00000000} /* (1, 27, 13) {real, imag} */,
  {32'h3f57bf04, 32'h00000000} /* (1, 27, 12) {real, imag} */,
  {32'h3f4555de, 32'h00000000} /* (1, 27, 11) {real, imag} */,
  {32'hbe187d82, 32'h00000000} /* (1, 27, 10) {real, imag} */,
  {32'hbeeefdbe, 32'h00000000} /* (1, 27, 9) {real, imag} */,
  {32'hbf31cf94, 32'h00000000} /* (1, 27, 8) {real, imag} */,
  {32'hbf3d5262, 32'h00000000} /* (1, 27, 7) {real, imag} */,
  {32'hbf0cfa5e, 32'h00000000} /* (1, 27, 6) {real, imag} */,
  {32'hbf5e0b37, 32'h00000000} /* (1, 27, 5) {real, imag} */,
  {32'hbf3a136f, 32'h00000000} /* (1, 27, 4) {real, imag} */,
  {32'hbf512dfd, 32'h00000000} /* (1, 27, 3) {real, imag} */,
  {32'hbf96b0f7, 32'h00000000} /* (1, 27, 2) {real, imag} */,
  {32'hbf2b781f, 32'h00000000} /* (1, 27, 1) {real, imag} */,
  {32'hbea7d549, 32'h00000000} /* (1, 27, 0) {real, imag} */,
  {32'hbeea5b9a, 32'h00000000} /* (1, 26, 31) {real, imag} */,
  {32'hbfabb60e, 32'h00000000} /* (1, 26, 30) {real, imag} */,
  {32'hbfb60a0d, 32'h00000000} /* (1, 26, 29) {real, imag} */,
  {32'hbf48e208, 32'h00000000} /* (1, 26, 28) {real, imag} */,
  {32'hbedcc81b, 32'h00000000} /* (1, 26, 27) {real, imag} */,
  {32'hbefd6ad9, 32'h00000000} /* (1, 26, 26) {real, imag} */,
  {32'hbf31902a, 32'h00000000} /* (1, 26, 25) {real, imag} */,
  {32'hbf156c33, 32'h00000000} /* (1, 26, 24) {real, imag} */,
  {32'hbf639bfa, 32'h00000000} /* (1, 26, 23) {real, imag} */,
  {32'hbf5ae47a, 32'h00000000} /* (1, 26, 22) {real, imag} */,
  {32'hbea70384, 32'h00000000} /* (1, 26, 21) {real, imag} */,
  {32'h3f1aaa87, 32'h00000000} /* (1, 26, 20) {real, imag} */,
  {32'h3f58a0ce, 32'h00000000} /* (1, 26, 19) {real, imag} */,
  {32'h3f082969, 32'h00000000} /* (1, 26, 18) {real, imag} */,
  {32'h3f48fccb, 32'h00000000} /* (1, 26, 17) {real, imag} */,
  {32'h3f41794d, 32'h00000000} /* (1, 26, 16) {real, imag} */,
  {32'h3ed52ca5, 32'h00000000} /* (1, 26, 15) {real, imag} */,
  {32'h3f03088f, 32'h00000000} /* (1, 26, 14) {real, imag} */,
  {32'h3eb159e6, 32'h00000000} /* (1, 26, 13) {real, imag} */,
  {32'h3f297ce4, 32'h00000000} /* (1, 26, 12) {real, imag} */,
  {32'h3f5ec77f, 32'h00000000} /* (1, 26, 11) {real, imag} */,
  {32'h3d846a9b, 32'h00000000} /* (1, 26, 10) {real, imag} */,
  {32'hbf9116f7, 32'h00000000} /* (1, 26, 9) {real, imag} */,
  {32'hbf42e569, 32'h00000000} /* (1, 26, 8) {real, imag} */,
  {32'hbe52eda6, 32'h00000000} /* (1, 26, 7) {real, imag} */,
  {32'hbf03dbb1, 32'h00000000} /* (1, 26, 6) {real, imag} */,
  {32'hbf0745ed, 32'h00000000} /* (1, 26, 5) {real, imag} */,
  {32'hbf4c307c, 32'h00000000} /* (1, 26, 4) {real, imag} */,
  {32'hbf8dd5da, 32'h00000000} /* (1, 26, 3) {real, imag} */,
  {32'hbfaf2d0e, 32'h00000000} /* (1, 26, 2) {real, imag} */,
  {32'hbf9766c0, 32'h00000000} /* (1, 26, 1) {real, imag} */,
  {32'hbf17f9f1, 32'h00000000} /* (1, 26, 0) {real, imag} */,
  {32'hbf3d8949, 32'h00000000} /* (1, 25, 31) {real, imag} */,
  {32'hbfa76e7e, 32'h00000000} /* (1, 25, 30) {real, imag} */,
  {32'hbf9054f8, 32'h00000000} /* (1, 25, 29) {real, imag} */,
  {32'hbf126ae2, 32'h00000000} /* (1, 25, 28) {real, imag} */,
  {32'hbf2498ce, 32'h00000000} /* (1, 25, 27) {real, imag} */,
  {32'hbf5b1ce1, 32'h00000000} /* (1, 25, 26) {real, imag} */,
  {32'hbf730e99, 32'h00000000} /* (1, 25, 25) {real, imag} */,
  {32'hbf45f0ce, 32'h00000000} /* (1, 25, 24) {real, imag} */,
  {32'hbf2df76e, 32'h00000000} /* (1, 25, 23) {real, imag} */,
  {32'hbf433738, 32'h00000000} /* (1, 25, 22) {real, imag} */,
  {32'hba881e22, 32'h00000000} /* (1, 25, 21) {real, imag} */,
  {32'h3fb70985, 32'h00000000} /* (1, 25, 20) {real, imag} */,
  {32'h3fb39415, 32'h00000000} /* (1, 25, 19) {real, imag} */,
  {32'h3f626b73, 32'h00000000} /* (1, 25, 18) {real, imag} */,
  {32'h3ef02c00, 32'h00000000} /* (1, 25, 17) {real, imag} */,
  {32'h3f3e3956, 32'h00000000} /* (1, 25, 16) {real, imag} */,
  {32'h3f72ed4f, 32'h00000000} /* (1, 25, 15) {real, imag} */,
  {32'h3f369646, 32'h00000000} /* (1, 25, 14) {real, imag} */,
  {32'h3e361ad6, 32'h00000000} /* (1, 25, 13) {real, imag} */,
  {32'h3ee84259, 32'h00000000} /* (1, 25, 12) {real, imag} */,
  {32'h3f4b1242, 32'h00000000} /* (1, 25, 11) {real, imag} */,
  {32'hbdea423c, 32'h00000000} /* (1, 25, 10) {real, imag} */,
  {32'hbfdf9a08, 32'h00000000} /* (1, 25, 9) {real, imag} */,
  {32'hbfb654fb, 32'h00000000} /* (1, 25, 8) {real, imag} */,
  {32'hbf553972, 32'h00000000} /* (1, 25, 7) {real, imag} */,
  {32'hbf259ec6, 32'h00000000} /* (1, 25, 6) {real, imag} */,
  {32'hbf11b653, 32'h00000000} /* (1, 25, 5) {real, imag} */,
  {32'hbf8332fe, 32'h00000000} /* (1, 25, 4) {real, imag} */,
  {32'hbf76737b, 32'h00000000} /* (1, 25, 3) {real, imag} */,
  {32'hbf40825a, 32'h00000000} /* (1, 25, 2) {real, imag} */,
  {32'hbfad1987, 32'h00000000} /* (1, 25, 1) {real, imag} */,
  {32'hbf843c5f, 32'h00000000} /* (1, 25, 0) {real, imag} */,
  {32'hbf3b8673, 32'h00000000} /* (1, 24, 31) {real, imag} */,
  {32'hbf57e1af, 32'h00000000} /* (1, 24, 30) {real, imag} */,
  {32'hbef397c2, 32'h00000000} /* (1, 24, 29) {real, imag} */,
  {32'hbe5f6bd0, 32'h00000000} /* (1, 24, 28) {real, imag} */,
  {32'hbf160f82, 32'h00000000} /* (1, 24, 27) {real, imag} */,
  {32'hbf86b61a, 32'h00000000} /* (1, 24, 26) {real, imag} */,
  {32'hbf5d045c, 32'h00000000} /* (1, 24, 25) {real, imag} */,
  {32'hbf69a369, 32'h00000000} /* (1, 24, 24) {real, imag} */,
  {32'hbf362bc2, 32'h00000000} /* (1, 24, 23) {real, imag} */,
  {32'hbf236523, 32'h00000000} /* (1, 24, 22) {real, imag} */,
  {32'h3e1e1b2c, 32'h00000000} /* (1, 24, 21) {real, imag} */,
  {32'h3fe45d84, 32'h00000000} /* (1, 24, 20) {real, imag} */,
  {32'h3fa6711f, 32'h00000000} /* (1, 24, 19) {real, imag} */,
  {32'h3f91aeab, 32'h00000000} /* (1, 24, 18) {real, imag} */,
  {32'h3f5029b2, 32'h00000000} /* (1, 24, 17) {real, imag} */,
  {32'h3f05097c, 32'h00000000} /* (1, 24, 16) {real, imag} */,
  {32'h3f43db05, 32'h00000000} /* (1, 24, 15) {real, imag} */,
  {32'h3f828b65, 32'h00000000} /* (1, 24, 14) {real, imag} */,
  {32'h3f25a74b, 32'h00000000} /* (1, 24, 13) {real, imag} */,
  {32'h3ec65b49, 32'h00000000} /* (1, 24, 12) {real, imag} */,
  {32'h3ef32b1b, 32'h00000000} /* (1, 24, 11) {real, imag} */,
  {32'hbf7df8d5, 32'h00000000} /* (1, 24, 10) {real, imag} */,
  {32'hbfc384cb, 32'h00000000} /* (1, 24, 9) {real, imag} */,
  {32'hbf98fa04, 32'h00000000} /* (1, 24, 8) {real, imag} */,
  {32'hbf4fd3d0, 32'h00000000} /* (1, 24, 7) {real, imag} */,
  {32'hbf0d33da, 32'h00000000} /* (1, 24, 6) {real, imag} */,
  {32'hbf55cba5, 32'h00000000} /* (1, 24, 5) {real, imag} */,
  {32'hbf3e1a60, 32'h00000000} /* (1, 24, 4) {real, imag} */,
  {32'hbf2c9aed, 32'h00000000} /* (1, 24, 3) {real, imag} */,
  {32'hbf248c28, 32'h00000000} /* (1, 24, 2) {real, imag} */,
  {32'hbf42f581, 32'h00000000} /* (1, 24, 1) {real, imag} */,
  {32'hbf2799e1, 32'h00000000} /* (1, 24, 0) {real, imag} */,
  {32'hbf1f3c6c, 32'h00000000} /* (1, 23, 31) {real, imag} */,
  {32'hbf3797cb, 32'h00000000} /* (1, 23, 30) {real, imag} */,
  {32'hbf25ee35, 32'h00000000} /* (1, 23, 29) {real, imag} */,
  {32'hbf01bd32, 32'h00000000} /* (1, 23, 28) {real, imag} */,
  {32'hbf4e0894, 32'h00000000} /* (1, 23, 27) {real, imag} */,
  {32'hbf8124b0, 32'h00000000} /* (1, 23, 26) {real, imag} */,
  {32'hbf3f4190, 32'h00000000} /* (1, 23, 25) {real, imag} */,
  {32'hbefdf4a4, 32'h00000000} /* (1, 23, 24) {real, imag} */,
  {32'hbea189dd, 32'h00000000} /* (1, 23, 23) {real, imag} */,
  {32'hbe3e62e4, 32'h00000000} /* (1, 23, 22) {real, imag} */,
  {32'hba110900, 32'h00000000} /* (1, 23, 21) {real, imag} */,
  {32'h3f9cf4a9, 32'h00000000} /* (1, 23, 20) {real, imag} */,
  {32'h3f6d1ff7, 32'h00000000} /* (1, 23, 19) {real, imag} */,
  {32'h3f478a7c, 32'h00000000} /* (1, 23, 18) {real, imag} */,
  {32'h3f57c419, 32'h00000000} /* (1, 23, 17) {real, imag} */,
  {32'h3f307d44, 32'h00000000} /* (1, 23, 16) {real, imag} */,
  {32'h3f062ee0, 32'h00000000} /* (1, 23, 15) {real, imag} */,
  {32'h3f25d204, 32'h00000000} /* (1, 23, 14) {real, imag} */,
  {32'h3f424380, 32'h00000000} /* (1, 23, 13) {real, imag} */,
  {32'h3f324655, 32'h00000000} /* (1, 23, 12) {real, imag} */,
  {32'h3f931714, 32'h00000000} /* (1, 23, 11) {real, imag} */,
  {32'hbe7c42e2, 32'h00000000} /* (1, 23, 10) {real, imag} */,
  {32'hbf3d4405, 32'h00000000} /* (1, 23, 9) {real, imag} */,
  {32'hbf73d6ef, 32'h00000000} /* (1, 23, 8) {real, imag} */,
  {32'hbf377913, 32'h00000000} /* (1, 23, 7) {real, imag} */,
  {32'hbe64eecc, 32'h00000000} /* (1, 23, 6) {real, imag} */,
  {32'hbf183443, 32'h00000000} /* (1, 23, 5) {real, imag} */,
  {32'hbf2b58a7, 32'h00000000} /* (1, 23, 4) {real, imag} */,
  {32'hbeb5bef7, 32'h00000000} /* (1, 23, 3) {real, imag} */,
  {32'hbf0e9baf, 32'h00000000} /* (1, 23, 2) {real, imag} */,
  {32'hbf6cac9e, 32'h00000000} /* (1, 23, 1) {real, imag} */,
  {32'hbec9e07b, 32'h00000000} /* (1, 23, 0) {real, imag} */,
  {32'hbf1754c1, 32'h00000000} /* (1, 22, 31) {real, imag} */,
  {32'hbe8ba1c7, 32'h00000000} /* (1, 22, 30) {real, imag} */,
  {32'hbee2a9d1, 32'h00000000} /* (1, 22, 29) {real, imag} */,
  {32'hbfa5d7ca, 32'h00000000} /* (1, 22, 28) {real, imag} */,
  {32'hbfb59d50, 32'h00000000} /* (1, 22, 27) {real, imag} */,
  {32'hbf7266c8, 32'h00000000} /* (1, 22, 26) {real, imag} */,
  {32'hbf560691, 32'h00000000} /* (1, 22, 25) {real, imag} */,
  {32'hbf21d9cf, 32'h00000000} /* (1, 22, 24) {real, imag} */,
  {32'hbeb47e0f, 32'h00000000} /* (1, 22, 23) {real, imag} */,
  {32'hbecf075c, 32'h00000000} /* (1, 22, 22) {real, imag} */,
  {32'hbef7e6ce, 32'h00000000} /* (1, 22, 21) {real, imag} */,
  {32'h3f635127, 32'h00000000} /* (1, 22, 20) {real, imag} */,
  {32'h3f58f939, 32'h00000000} /* (1, 22, 19) {real, imag} */,
  {32'h3edd8f2d, 32'h00000000} /* (1, 22, 18) {real, imag} */,
  {32'h3f1bf6ff, 32'h00000000} /* (1, 22, 17) {real, imag} */,
  {32'h3f8a0264, 32'h00000000} /* (1, 22, 16) {real, imag} */,
  {32'h3f3218b2, 32'h00000000} /* (1, 22, 15) {real, imag} */,
  {32'h3f4f0c4c, 32'h00000000} /* (1, 22, 14) {real, imag} */,
  {32'h3f8aee3e, 32'h00000000} /* (1, 22, 13) {real, imag} */,
  {32'h3f827f73, 32'h00000000} /* (1, 22, 12) {real, imag} */,
  {32'h3f60e1bb, 32'h00000000} /* (1, 22, 11) {real, imag} */,
  {32'hbe77fee9, 32'h00000000} /* (1, 22, 10) {real, imag} */,
  {32'hbf801c02, 32'h00000000} /* (1, 22, 9) {real, imag} */,
  {32'hbf81dfba, 32'h00000000} /* (1, 22, 8) {real, imag} */,
  {32'hbf1394a9, 32'h00000000} /* (1, 22, 7) {real, imag} */,
  {32'hbecaf800, 32'h00000000} /* (1, 22, 6) {real, imag} */,
  {32'hbf2094ba, 32'h00000000} /* (1, 22, 5) {real, imag} */,
  {32'hbf0dc85c, 32'h00000000} /* (1, 22, 4) {real, imag} */,
  {32'hbed2fa24, 32'h00000000} /* (1, 22, 3) {real, imag} */,
  {32'hbf1cabd2, 32'h00000000} /* (1, 22, 2) {real, imag} */,
  {32'hbf160987, 32'h00000000} /* (1, 22, 1) {real, imag} */,
  {32'hbed59326, 32'h00000000} /* (1, 22, 0) {real, imag} */,
  {32'hbf3c81dc, 32'h00000000} /* (1, 21, 31) {real, imag} */,
  {32'hbea85180, 32'h00000000} /* (1, 21, 30) {real, imag} */,
  {32'h3d88ed43, 32'h00000000} /* (1, 21, 29) {real, imag} */,
  {32'hbf71811e, 32'h00000000} /* (1, 21, 28) {real, imag} */,
  {32'hbf20c4b9, 32'h00000000} /* (1, 21, 27) {real, imag} */,
  {32'hbe68ad5e, 32'h00000000} /* (1, 21, 26) {real, imag} */,
  {32'hbe8dc8fa, 32'h00000000} /* (1, 21, 25) {real, imag} */,
  {32'hbf0be70d, 32'h00000000} /* (1, 21, 24) {real, imag} */,
  {32'hbec75b0c, 32'h00000000} /* (1, 21, 23) {real, imag} */,
  {32'hbebd6ed9, 32'h00000000} /* (1, 21, 22) {real, imag} */,
  {32'hbeed66e7, 32'h00000000} /* (1, 21, 21) {real, imag} */,
  {32'h3d16e15d, 32'h00000000} /* (1, 21, 20) {real, imag} */,
  {32'h3e7dac37, 32'h00000000} /* (1, 21, 19) {real, imag} */,
  {32'h3ed2cd1b, 32'h00000000} /* (1, 21, 18) {real, imag} */,
  {32'h3c8265a4, 32'h00000000} /* (1, 21, 17) {real, imag} */,
  {32'h3e85c37c, 32'h00000000} /* (1, 21, 16) {real, imag} */,
  {32'h3ebb541a, 32'h00000000} /* (1, 21, 15) {real, imag} */,
  {32'h3ec4cdb4, 32'h00000000} /* (1, 21, 14) {real, imag} */,
  {32'h3f069f5e, 32'h00000000} /* (1, 21, 13) {real, imag} */,
  {32'h3ecb2441, 32'h00000000} /* (1, 21, 12) {real, imag} */,
  {32'h3edb3f1b, 32'h00000000} /* (1, 21, 11) {real, imag} */,
  {32'hbd82075b, 32'h00000000} /* (1, 21, 10) {real, imag} */,
  {32'hbf10090f, 32'h00000000} /* (1, 21, 9) {real, imag} */,
  {32'hbf185f14, 32'h00000000} /* (1, 21, 8) {real, imag} */,
  {32'hbec0a410, 32'h00000000} /* (1, 21, 7) {real, imag} */,
  {32'hbe8bf769, 32'h00000000} /* (1, 21, 6) {real, imag} */,
  {32'hbec60432, 32'h00000000} /* (1, 21, 5) {real, imag} */,
  {32'hbea990d9, 32'h00000000} /* (1, 21, 4) {real, imag} */,
  {32'hbd4e02c5, 32'h00000000} /* (1, 21, 3) {real, imag} */,
  {32'hbe234801, 32'h00000000} /* (1, 21, 2) {real, imag} */,
  {32'hbe9b0cd1, 32'h00000000} /* (1, 21, 1) {real, imag} */,
  {32'hbec60adb, 32'h00000000} /* (1, 21, 0) {real, imag} */,
  {32'h3e384afb, 32'h00000000} /* (1, 20, 31) {real, imag} */,
  {32'h3f1738d7, 32'h00000000} /* (1, 20, 30) {real, imag} */,
  {32'h3f86dc2e, 32'h00000000} /* (1, 20, 29) {real, imag} */,
  {32'h3f395aa4, 32'h00000000} /* (1, 20, 28) {real, imag} */,
  {32'h3f01cbb5, 32'h00000000} /* (1, 20, 27) {real, imag} */,
  {32'h3e811703, 32'h00000000} /* (1, 20, 26) {real, imag} */,
  {32'h3f96bd31, 32'h00000000} /* (1, 20, 25) {real, imag} */,
  {32'h3f760766, 32'h00000000} /* (1, 20, 24) {real, imag} */,
  {32'h3f2a3a5e, 32'h00000000} /* (1, 20, 23) {real, imag} */,
  {32'h3f76277e, 32'h00000000} /* (1, 20, 22) {real, imag} */,
  {32'h3eebf2aa, 32'h00000000} /* (1, 20, 21) {real, imag} */,
  {32'hbebcb279, 32'h00000000} /* (1, 20, 20) {real, imag} */,
  {32'hbf524606, 32'h00000000} /* (1, 20, 19) {real, imag} */,
  {32'hbf44963a, 32'h00000000} /* (1, 20, 18) {real, imag} */,
  {32'hbf4a87d9, 32'h00000000} /* (1, 20, 17) {real, imag} */,
  {32'hbf572135, 32'h00000000} /* (1, 20, 16) {real, imag} */,
  {32'hbf8ce733, 32'h00000000} /* (1, 20, 15) {real, imag} */,
  {32'hbf3a1d4f, 32'h00000000} /* (1, 20, 14) {real, imag} */,
  {32'hbf07f6e2, 32'h00000000} /* (1, 20, 13) {real, imag} */,
  {32'hbf03bd6a, 32'h00000000} /* (1, 20, 12) {real, imag} */,
  {32'hbee3fd0d, 32'h00000000} /* (1, 20, 11) {real, imag} */,
  {32'hbe4c873c, 32'h00000000} /* (1, 20, 10) {real, imag} */,
  {32'h3e8cffdc, 32'h00000000} /* (1, 20, 9) {real, imag} */,
  {32'h3e87f5f3, 32'h00000000} /* (1, 20, 8) {real, imag} */,
  {32'h3ebd896e, 32'h00000000} /* (1, 20, 7) {real, imag} */,
  {32'h3f03a821, 32'h00000000} /* (1, 20, 6) {real, imag} */,
  {32'h3ec86b73, 32'h00000000} /* (1, 20, 5) {real, imag} */,
  {32'h3efae826, 32'h00000000} /* (1, 20, 4) {real, imag} */,
  {32'h3f657769, 32'h00000000} /* (1, 20, 3) {real, imag} */,
  {32'h3f8d4008, 32'h00000000} /* (1, 20, 2) {real, imag} */,
  {32'h3f00e6e2, 32'h00000000} /* (1, 20, 1) {real, imag} */,
  {32'h3b515894, 32'h00000000} /* (1, 20, 0) {real, imag} */,
  {32'h3f4fdcdf, 32'h00000000} /* (1, 19, 31) {real, imag} */,
  {32'h3f752f82, 32'h00000000} /* (1, 19, 30) {real, imag} */,
  {32'h3f4465a2, 32'h00000000} /* (1, 19, 29) {real, imag} */,
  {32'h3f136c8b, 32'h00000000} /* (1, 19, 28) {real, imag} */,
  {32'h3f421b0d, 32'h00000000} /* (1, 19, 27) {real, imag} */,
  {32'h3f07979a, 32'h00000000} /* (1, 19, 26) {real, imag} */,
  {32'h3f8557af, 32'h00000000} /* (1, 19, 25) {real, imag} */,
  {32'h3f8ff15a, 32'h00000000} /* (1, 19, 24) {real, imag} */,
  {32'h3fa09a7f, 32'h00000000} /* (1, 19, 23) {real, imag} */,
  {32'h3fb1b75e, 32'h00000000} /* (1, 19, 22) {real, imag} */,
  {32'h3f304b15, 32'h00000000} /* (1, 19, 21) {real, imag} */,
  {32'hbeb55881, 32'h00000000} /* (1, 19, 20) {real, imag} */,
  {32'hbf160a99, 32'h00000000} /* (1, 19, 19) {real, imag} */,
  {32'hbf73f356, 32'h00000000} /* (1, 19, 18) {real, imag} */,
  {32'hbf600819, 32'h00000000} /* (1, 19, 17) {real, imag} */,
  {32'hbf501f46, 32'h00000000} /* (1, 19, 16) {real, imag} */,
  {32'hbf5b23d9, 32'h00000000} /* (1, 19, 15) {real, imag} */,
  {32'hbf3d41a8, 32'h00000000} /* (1, 19, 14) {real, imag} */,
  {32'hbf5875f7, 32'h00000000} /* (1, 19, 13) {real, imag} */,
  {32'hbf805218, 32'h00000000} /* (1, 19, 12) {real, imag} */,
  {32'hbf5e9954, 32'h00000000} /* (1, 19, 11) {real, imag} */,
  {32'hbdca824c, 32'h00000000} /* (1, 19, 10) {real, imag} */,
  {32'h3ee04db5, 32'h00000000} /* (1, 19, 9) {real, imag} */,
  {32'h3f23a81d, 32'h00000000} /* (1, 19, 8) {real, imag} */,
  {32'h3f81af9c, 32'h00000000} /* (1, 19, 7) {real, imag} */,
  {32'h3f297639, 32'h00000000} /* (1, 19, 6) {real, imag} */,
  {32'h3f4764c5, 32'h00000000} /* (1, 19, 5) {real, imag} */,
  {32'h3f983eb8, 32'h00000000} /* (1, 19, 4) {real, imag} */,
  {32'h3fc6def1, 32'h00000000} /* (1, 19, 3) {real, imag} */,
  {32'h3f8dddff, 32'h00000000} /* (1, 19, 2) {real, imag} */,
  {32'h3f7c70f1, 32'h00000000} /* (1, 19, 1) {real, imag} */,
  {32'h3f208d09, 32'h00000000} /* (1, 19, 0) {real, imag} */,
  {32'h3f0d9aff, 32'h00000000} /* (1, 18, 31) {real, imag} */,
  {32'h3f46a5f0, 32'h00000000} /* (1, 18, 30) {real, imag} */,
  {32'h3e767443, 32'h00000000} /* (1, 18, 29) {real, imag} */,
  {32'h3e96bc6a, 32'h00000000} /* (1, 18, 28) {real, imag} */,
  {32'h3f772307, 32'h00000000} /* (1, 18, 27) {real, imag} */,
  {32'h3f8c58e7, 32'h00000000} /* (1, 18, 26) {real, imag} */,
  {32'h3f5b5923, 32'h00000000} /* (1, 18, 25) {real, imag} */,
  {32'h3f4d9749, 32'h00000000} /* (1, 18, 24) {real, imag} */,
  {32'h3f6ed5c2, 32'h00000000} /* (1, 18, 23) {real, imag} */,
  {32'h3f689054, 32'h00000000} /* (1, 18, 22) {real, imag} */,
  {32'hbd00fcea, 32'h00000000} /* (1, 18, 21) {real, imag} */,
  {32'hbf01e96c, 32'h00000000} /* (1, 18, 20) {real, imag} */,
  {32'hbf089030, 32'h00000000} /* (1, 18, 19) {real, imag} */,
  {32'hbf32de0f, 32'h00000000} /* (1, 18, 18) {real, imag} */,
  {32'hbf287835, 32'h00000000} /* (1, 18, 17) {real, imag} */,
  {32'hbede1aca, 32'h00000000} /* (1, 18, 16) {real, imag} */,
  {32'hbee5b104, 32'h00000000} /* (1, 18, 15) {real, imag} */,
  {32'hbf501580, 32'h00000000} /* (1, 18, 14) {real, imag} */,
  {32'hbf95398b, 32'h00000000} /* (1, 18, 13) {real, imag} */,
  {32'hbf486243, 32'h00000000} /* (1, 18, 12) {real, imag} */,
  {32'hbed80058, 32'h00000000} /* (1, 18, 11) {real, imag} */,
  {32'h3f17232a, 32'h00000000} /* (1, 18, 10) {real, imag} */,
  {32'h3f36a42b, 32'h00000000} /* (1, 18, 9) {real, imag} */,
  {32'h3f4d3698, 32'h00000000} /* (1, 18, 8) {real, imag} */,
  {32'h3fb38443, 32'h00000000} /* (1, 18, 7) {real, imag} */,
  {32'h3f42cb62, 32'h00000000} /* (1, 18, 6) {real, imag} */,
  {32'h3f2e5768, 32'h00000000} /* (1, 18, 5) {real, imag} */,
  {32'h3f366abd, 32'h00000000} /* (1, 18, 4) {real, imag} */,
  {32'h3f7a468a, 32'h00000000} /* (1, 18, 3) {real, imag} */,
  {32'h3f7acf56, 32'h00000000} /* (1, 18, 2) {real, imag} */,
  {32'h3f1eb9d4, 32'h00000000} /* (1, 18, 1) {real, imag} */,
  {32'h3f230b15, 32'h00000000} /* (1, 18, 0) {real, imag} */,
  {32'h3f2e4750, 32'h00000000} /* (1, 17, 31) {real, imag} */,
  {32'h3f5e30c0, 32'h00000000} /* (1, 17, 30) {real, imag} */,
  {32'h3f14fa54, 32'h00000000} /* (1, 17, 29) {real, imag} */,
  {32'h3f546fe6, 32'h00000000} /* (1, 17, 28) {real, imag} */,
  {32'h3f819dcd, 32'h00000000} /* (1, 17, 27) {real, imag} */,
  {32'h3f8333f0, 32'h00000000} /* (1, 17, 26) {real, imag} */,
  {32'h3f811264, 32'h00000000} /* (1, 17, 25) {real, imag} */,
  {32'h3f0e811f, 32'h00000000} /* (1, 17, 24) {real, imag} */,
  {32'h3f973f22, 32'h00000000} /* (1, 17, 23) {real, imag} */,
  {32'h3fa73fce, 32'h00000000} /* (1, 17, 22) {real, imag} */,
  {32'hbb2a3501, 32'h00000000} /* (1, 17, 21) {real, imag} */,
  {32'hbebfc93f, 32'h00000000} /* (1, 17, 20) {real, imag} */,
  {32'hbf07cf24, 32'h00000000} /* (1, 17, 19) {real, imag} */,
  {32'hbf36ead1, 32'h00000000} /* (1, 17, 18) {real, imag} */,
  {32'hbf816d52, 32'h00000000} /* (1, 17, 17) {real, imag} */,
  {32'hbf4e4391, 32'h00000000} /* (1, 17, 16) {real, imag} */,
  {32'hbf080dc4, 32'h00000000} /* (1, 17, 15) {real, imag} */,
  {32'hbef476b5, 32'h00000000} /* (1, 17, 14) {real, imag} */,
  {32'hbf55dd93, 32'h00000000} /* (1, 17, 13) {real, imag} */,
  {32'hbf3a91fc, 32'h00000000} /* (1, 17, 12) {real, imag} */,
  {32'hbebb297a, 32'h00000000} /* (1, 17, 11) {real, imag} */,
  {32'h3f5143df, 32'h00000000} /* (1, 17, 10) {real, imag} */,
  {32'h3f9f578b, 32'h00000000} /* (1, 17, 9) {real, imag} */,
  {32'h3f7a3d49, 32'h00000000} /* (1, 17, 8) {real, imag} */,
  {32'h3f6f8f55, 32'h00000000} /* (1, 17, 7) {real, imag} */,
  {32'h3fcbf015, 32'h00000000} /* (1, 17, 6) {real, imag} */,
  {32'h3f552859, 32'h00000000} /* (1, 17, 5) {real, imag} */,
  {32'h3e95823a, 32'h00000000} /* (1, 17, 4) {real, imag} */,
  {32'h3e92c54f, 32'h00000000} /* (1, 17, 3) {real, imag} */,
  {32'h3ec5c78f, 32'h00000000} /* (1, 17, 2) {real, imag} */,
  {32'h3f0227c6, 32'h00000000} /* (1, 17, 1) {real, imag} */,
  {32'h3f0ff425, 32'h00000000} /* (1, 17, 0) {real, imag} */,
  {32'h3e956f57, 32'h00000000} /* (1, 16, 31) {real, imag} */,
  {32'h3f1c9073, 32'h00000000} /* (1, 16, 30) {real, imag} */,
  {32'h3f60347f, 32'h00000000} /* (1, 16, 29) {real, imag} */,
  {32'h3f665d04, 32'h00000000} /* (1, 16, 28) {real, imag} */,
  {32'h3f52a1ed, 32'h00000000} /* (1, 16, 27) {real, imag} */,
  {32'h3f3a752a, 32'h00000000} /* (1, 16, 26) {real, imag} */,
  {32'h3f3faabd, 32'h00000000} /* (1, 16, 25) {real, imag} */,
  {32'h3ea5ae95, 32'h00000000} /* (1, 16, 24) {real, imag} */,
  {32'h3f6ccb20, 32'h00000000} /* (1, 16, 23) {real, imag} */,
  {32'h3fca962e, 32'h00000000} /* (1, 16, 22) {real, imag} */,
  {32'h3f46a399, 32'h00000000} /* (1, 16, 21) {real, imag} */,
  {32'hbedea625, 32'h00000000} /* (1, 16, 20) {real, imag} */,
  {32'hbf36ea5e, 32'h00000000} /* (1, 16, 19) {real, imag} */,
  {32'hbf0c6ca6, 32'h00000000} /* (1, 16, 18) {real, imag} */,
  {32'hbf563bb8, 32'h00000000} /* (1, 16, 17) {real, imag} */,
  {32'hbf569de2, 32'h00000000} /* (1, 16, 16) {real, imag} */,
  {32'hbf494f84, 32'h00000000} /* (1, 16, 15) {real, imag} */,
  {32'hbf23e515, 32'h00000000} /* (1, 16, 14) {real, imag} */,
  {32'hbf1681fe, 32'h00000000} /* (1, 16, 13) {real, imag} */,
  {32'hbf368feb, 32'h00000000} /* (1, 16, 12) {real, imag} */,
  {32'hbf019eda, 32'h00000000} /* (1, 16, 11) {real, imag} */,
  {32'h3f1b666e, 32'h00000000} /* (1, 16, 10) {real, imag} */,
  {32'h3fd31338, 32'h00000000} /* (1, 16, 9) {real, imag} */,
  {32'h3f9f7b73, 32'h00000000} /* (1, 16, 8) {real, imag} */,
  {32'h3f8f40d4, 32'h00000000} /* (1, 16, 7) {real, imag} */,
  {32'h3fbf6056, 32'h00000000} /* (1, 16, 6) {real, imag} */,
  {32'h3f2c6c52, 32'h00000000} /* (1, 16, 5) {real, imag} */,
  {32'h3e8b832a, 32'h00000000} /* (1, 16, 4) {real, imag} */,
  {32'h3e7fb248, 32'h00000000} /* (1, 16, 3) {real, imag} */,
  {32'h3edb80a9, 32'h00000000} /* (1, 16, 2) {real, imag} */,
  {32'h3f745cd5, 32'h00000000} /* (1, 16, 1) {real, imag} */,
  {32'h3f2b00ed, 32'h00000000} /* (1, 16, 0) {real, imag} */,
  {32'h3ecbc114, 32'h00000000} /* (1, 15, 31) {real, imag} */,
  {32'h3f5d77da, 32'h00000000} /* (1, 15, 30) {real, imag} */,
  {32'h3fa49cf4, 32'h00000000} /* (1, 15, 29) {real, imag} */,
  {32'h3f77c3d2, 32'h00000000} /* (1, 15, 28) {real, imag} */,
  {32'h3f4d2785, 32'h00000000} /* (1, 15, 27) {real, imag} */,
  {32'h3f3e635f, 32'h00000000} /* (1, 15, 26) {real, imag} */,
  {32'h3f08af18, 32'h00000000} /* (1, 15, 25) {real, imag} */,
  {32'h3edd9186, 32'h00000000} /* (1, 15, 24) {real, imag} */,
  {32'h3ebeb6aa, 32'h00000000} /* (1, 15, 23) {real, imag} */,
  {32'h3f5ef00f, 32'h00000000} /* (1, 15, 22) {real, imag} */,
  {32'h3f213875, 32'h00000000} /* (1, 15, 21) {real, imag} */,
  {32'hbf26c984, 32'h00000000} /* (1, 15, 20) {real, imag} */,
  {32'hbf55f671, 32'h00000000} /* (1, 15, 19) {real, imag} */,
  {32'hbed6b41d, 32'h00000000} /* (1, 15, 18) {real, imag} */,
  {32'hbf049a22, 32'h00000000} /* (1, 15, 17) {real, imag} */,
  {32'hbf182aec, 32'h00000000} /* (1, 15, 16) {real, imag} */,
  {32'hbf13df09, 32'h00000000} /* (1, 15, 15) {real, imag} */,
  {32'hbf35287f, 32'h00000000} /* (1, 15, 14) {real, imag} */,
  {32'hbf88cbe7, 32'h00000000} /* (1, 15, 13) {real, imag} */,
  {32'hbf99f0e1, 32'h00000000} /* (1, 15, 12) {real, imag} */,
  {32'hbf380f95, 32'h00000000} /* (1, 15, 11) {real, imag} */,
  {32'h3e4e8a39, 32'h00000000} /* (1, 15, 10) {real, imag} */,
  {32'h3f7941ce, 32'h00000000} /* (1, 15, 9) {real, imag} */,
  {32'h3f634209, 32'h00000000} /* (1, 15, 8) {real, imag} */,
  {32'h3f86189e, 32'h00000000} /* (1, 15, 7) {real, imag} */,
  {32'h3f956fd3, 32'h00000000} /* (1, 15, 6) {real, imag} */,
  {32'h3f71cf8b, 32'h00000000} /* (1, 15, 5) {real, imag} */,
  {32'h3f878e2a, 32'h00000000} /* (1, 15, 4) {real, imag} */,
  {32'h3f318b58, 32'h00000000} /* (1, 15, 3) {real, imag} */,
  {32'h3f837eac, 32'h00000000} /* (1, 15, 2) {real, imag} */,
  {32'h3fa42661, 32'h00000000} /* (1, 15, 1) {real, imag} */,
  {32'h3ee3e499, 32'h00000000} /* (1, 15, 0) {real, imag} */,
  {32'h3f1881ca, 32'h00000000} /* (1, 14, 31) {real, imag} */,
  {32'h3fa3460b, 32'h00000000} /* (1, 14, 30) {real, imag} */,
  {32'h3fa73a9a, 32'h00000000} /* (1, 14, 29) {real, imag} */,
  {32'h3f5ec119, 32'h00000000} /* (1, 14, 28) {real, imag} */,
  {32'h3f8b0f48, 32'h00000000} /* (1, 14, 27) {real, imag} */,
  {32'h3f9777ef, 32'h00000000} /* (1, 14, 26) {real, imag} */,
  {32'h3f4a98a4, 32'h00000000} /* (1, 14, 25) {real, imag} */,
  {32'h3ef3eaf2, 32'h00000000} /* (1, 14, 24) {real, imag} */,
  {32'h3ed0daa8, 32'h00000000} /* (1, 14, 23) {real, imag} */,
  {32'h3f3d6b4c, 32'h00000000} /* (1, 14, 22) {real, imag} */,
  {32'h3e544f17, 32'h00000000} /* (1, 14, 21) {real, imag} */,
  {32'hbf24e659, 32'h00000000} /* (1, 14, 20) {real, imag} */,
  {32'hbf8f2506, 32'h00000000} /* (1, 14, 19) {real, imag} */,
  {32'hbf94d93f, 32'h00000000} /* (1, 14, 18) {real, imag} */,
  {32'hbfa35b5a, 32'h00000000} /* (1, 14, 17) {real, imag} */,
  {32'hbf1ff0ab, 32'h00000000} /* (1, 14, 16) {real, imag} */,
  {32'hbf26a933, 32'h00000000} /* (1, 14, 15) {real, imag} */,
  {32'hbf8a0fa9, 32'h00000000} /* (1, 14, 14) {real, imag} */,
  {32'hbfb27fc1, 32'h00000000} /* (1, 14, 13) {real, imag} */,
  {32'hbf88b463, 32'h00000000} /* (1, 14, 12) {real, imag} */,
  {32'hbf113ed4, 32'h00000000} /* (1, 14, 11) {real, imag} */,
  {32'h3eefc655, 32'h00000000} /* (1, 14, 10) {real, imag} */,
  {32'h3f599f5e, 32'h00000000} /* (1, 14, 9) {real, imag} */,
  {32'h3f808f9f, 32'h00000000} /* (1, 14, 8) {real, imag} */,
  {32'h3f444b76, 32'h00000000} /* (1, 14, 7) {real, imag} */,
  {32'h3f33d510, 32'h00000000} /* (1, 14, 6) {real, imag} */,
  {32'h3f74ef0c, 32'h00000000} /* (1, 14, 5) {real, imag} */,
  {32'h3f6f93ca, 32'h00000000} /* (1, 14, 4) {real, imag} */,
  {32'h3f8a17bf, 32'h00000000} /* (1, 14, 3) {real, imag} */,
  {32'h3f9a56da, 32'h00000000} /* (1, 14, 2) {real, imag} */,
  {32'h3f42ef89, 32'h00000000} /* (1, 14, 1) {real, imag} */,
  {32'h3e4cf495, 32'h00000000} /* (1, 14, 0) {real, imag} */,
  {32'h3e9fa62a, 32'h00000000} /* (1, 13, 31) {real, imag} */,
  {32'h3f6f67aa, 32'h00000000} /* (1, 13, 30) {real, imag} */,
  {32'h3fcd51f3, 32'h00000000} /* (1, 13, 29) {real, imag} */,
  {32'h3fa0ff03, 32'h00000000} /* (1, 13, 28) {real, imag} */,
  {32'h3fadee20, 32'h00000000} /* (1, 13, 27) {real, imag} */,
  {32'h3fcac4bc, 32'h00000000} /* (1, 13, 26) {real, imag} */,
  {32'h3f94ecf6, 32'h00000000} /* (1, 13, 25) {real, imag} */,
  {32'h3f2a51f7, 32'h00000000} /* (1, 13, 24) {real, imag} */,
  {32'h3f2e856d, 32'h00000000} /* (1, 13, 23) {real, imag} */,
  {32'h3f7ba619, 32'h00000000} /* (1, 13, 22) {real, imag} */,
  {32'h3e1da1f6, 32'h00000000} /* (1, 13, 21) {real, imag} */,
  {32'hbf686654, 32'h00000000} /* (1, 13, 20) {real, imag} */,
  {32'hbfbe0c12, 32'h00000000} /* (1, 13, 19) {real, imag} */,
  {32'hbfa529f6, 32'h00000000} /* (1, 13, 18) {real, imag} */,
  {32'hbfd0f5f6, 32'h00000000} /* (1, 13, 17) {real, imag} */,
  {32'hbfd3c11a, 32'h00000000} /* (1, 13, 16) {real, imag} */,
  {32'hbf1cc1ba, 32'h00000000} /* (1, 13, 15) {real, imag} */,
  {32'hbf2576a7, 32'h00000000} /* (1, 13, 14) {real, imag} */,
  {32'hbf3dbb00, 32'h00000000} /* (1, 13, 13) {real, imag} */,
  {32'hbf7265d0, 32'h00000000} /* (1, 13, 12) {real, imag} */,
  {32'hbf847217, 32'h00000000} /* (1, 13, 11) {real, imag} */,
  {32'h3e3e9e37, 32'h00000000} /* (1, 13, 10) {real, imag} */,
  {32'h3f5de0d5, 32'h00000000} /* (1, 13, 9) {real, imag} */,
  {32'h3fa46fd1, 32'h00000000} /* (1, 13, 8) {real, imag} */,
  {32'h3f80da31, 32'h00000000} /* (1, 13, 7) {real, imag} */,
  {32'h3ecb0678, 32'h00000000} /* (1, 13, 6) {real, imag} */,
  {32'h3f4ff11f, 32'h00000000} /* (1, 13, 5) {real, imag} */,
  {32'h3f0f49c1, 32'h00000000} /* (1, 13, 4) {real, imag} */,
  {32'h3f65eaa2, 32'h00000000} /* (1, 13, 3) {real, imag} */,
  {32'h3f93f968, 32'h00000000} /* (1, 13, 2) {real, imag} */,
  {32'h3f4425ad, 32'h00000000} /* (1, 13, 1) {real, imag} */,
  {32'h3f07271d, 32'h00000000} /* (1, 13, 0) {real, imag} */,
  {32'h3e6794fd, 32'h00000000} /* (1, 12, 31) {real, imag} */,
  {32'h3f0c27dd, 32'h00000000} /* (1, 12, 30) {real, imag} */,
  {32'h3f7095c8, 32'h00000000} /* (1, 12, 29) {real, imag} */,
  {32'h3f93c6bd, 32'h00000000} /* (1, 12, 28) {real, imag} */,
  {32'h3f8813c9, 32'h00000000} /* (1, 12, 27) {real, imag} */,
  {32'h3f70e027, 32'h00000000} /* (1, 12, 26) {real, imag} */,
  {32'h3f65e7c8, 32'h00000000} /* (1, 12, 25) {real, imag} */,
  {32'h3fb79ee2, 32'h00000000} /* (1, 12, 24) {real, imag} */,
  {32'h3fec571f, 32'h00000000} /* (1, 12, 23) {real, imag} */,
  {32'h3fb675ec, 32'h00000000} /* (1, 12, 22) {real, imag} */,
  {32'h3f219106, 32'h00000000} /* (1, 12, 21) {real, imag} */,
  {32'hbf4cb5f0, 32'h00000000} /* (1, 12, 20) {real, imag} */,
  {32'hbfa87562, 32'h00000000} /* (1, 12, 19) {real, imag} */,
  {32'hbf6cb2c1, 32'h00000000} /* (1, 12, 18) {real, imag} */,
  {32'hbfbdfa8f, 32'h00000000} /* (1, 12, 17) {real, imag} */,
  {32'hbfb489f8, 32'h00000000} /* (1, 12, 16) {real, imag} */,
  {32'hbf021cd8, 32'h00000000} /* (1, 12, 15) {real, imag} */,
  {32'hbefac53b, 32'h00000000} /* (1, 12, 14) {real, imag} */,
  {32'hbeb3b2c7, 32'h00000000} /* (1, 12, 13) {real, imag} */,
  {32'hbf554c34, 32'h00000000} /* (1, 12, 12) {real, imag} */,
  {32'hbf81b150, 32'h00000000} /* (1, 12, 11) {real, imag} */,
  {32'h3e5b8227, 32'h00000000} /* (1, 12, 10) {real, imag} */,
  {32'h3f329673, 32'h00000000} /* (1, 12, 9) {real, imag} */,
  {32'h3f4e3f87, 32'h00000000} /* (1, 12, 8) {real, imag} */,
  {32'h3f826d34, 32'h00000000} /* (1, 12, 7) {real, imag} */,
  {32'h3f6fd7d4, 32'h00000000} /* (1, 12, 6) {real, imag} */,
  {32'h3f8abdea, 32'h00000000} /* (1, 12, 5) {real, imag} */,
  {32'h3f5efd2d, 32'h00000000} /* (1, 12, 4) {real, imag} */,
  {32'h3f7c7eb8, 32'h00000000} /* (1, 12, 3) {real, imag} */,
  {32'h3f757504, 32'h00000000} /* (1, 12, 2) {real, imag} */,
  {32'h3f827f5f, 32'h00000000} /* (1, 12, 1) {real, imag} */,
  {32'h3f35c80b, 32'h00000000} /* (1, 12, 0) {real, imag} */,
  {32'h3ec5c1d0, 32'h00000000} /* (1, 11, 31) {real, imag} */,
  {32'h3eefee9d, 32'h00000000} /* (1, 11, 30) {real, imag} */,
  {32'h3f116c81, 32'h00000000} /* (1, 11, 29) {real, imag} */,
  {32'h3f2d7364, 32'h00000000} /* (1, 11, 28) {real, imag} */,
  {32'h3f31b1ab, 32'h00000000} /* (1, 11, 27) {real, imag} */,
  {32'h3ed50f5c, 32'h00000000} /* (1, 11, 26) {real, imag} */,
  {32'h3efd31e5, 32'h00000000} /* (1, 11, 25) {real, imag} */,
  {32'h3f981c5c, 32'h00000000} /* (1, 11, 24) {real, imag} */,
  {32'h3fabdff7, 32'h00000000} /* (1, 11, 23) {real, imag} */,
  {32'h3f54b8b9, 32'h00000000} /* (1, 11, 22) {real, imag} */,
  {32'h3ef1bc72, 32'h00000000} /* (1, 11, 21) {real, imag} */,
  {32'hbed8489c, 32'h00000000} /* (1, 11, 20) {real, imag} */,
  {32'hbee1f59b, 32'h00000000} /* (1, 11, 19) {real, imag} */,
  {32'hbf1a7d0b, 32'h00000000} /* (1, 11, 18) {real, imag} */,
  {32'hbf9457a4, 32'h00000000} /* (1, 11, 17) {real, imag} */,
  {32'hbf3f44d5, 32'h00000000} /* (1, 11, 16) {real, imag} */,
  {32'hbf5b62c0, 32'h00000000} /* (1, 11, 15) {real, imag} */,
  {32'hbf551f1c, 32'h00000000} /* (1, 11, 14) {real, imag} */,
  {32'hbf04d0a0, 32'h00000000} /* (1, 11, 13) {real, imag} */,
  {32'hbf920f34, 32'h00000000} /* (1, 11, 12) {real, imag} */,
  {32'hbf7861dc, 32'h00000000} /* (1, 11, 11) {real, imag} */,
  {32'hbd249656, 32'h00000000} /* (1, 11, 10) {real, imag} */,
  {32'h3e7cb36e, 32'h00000000} /* (1, 11, 9) {real, imag} */,
  {32'h3f1cacad, 32'h00000000} /* (1, 11, 8) {real, imag} */,
  {32'h3f6e0184, 32'h00000000} /* (1, 11, 7) {real, imag} */,
  {32'h3f96aaf2, 32'h00000000} /* (1, 11, 6) {real, imag} */,
  {32'h3f74bde8, 32'h00000000} /* (1, 11, 5) {real, imag} */,
  {32'h3f399626, 32'h00000000} /* (1, 11, 4) {real, imag} */,
  {32'h3ed6e4c2, 32'h00000000} /* (1, 11, 3) {real, imag} */,
  {32'h3e846472, 32'h00000000} /* (1, 11, 2) {real, imag} */,
  {32'h3ec9d3b6, 32'h00000000} /* (1, 11, 1) {real, imag} */,
  {32'h3ec340a1, 32'h00000000} /* (1, 11, 0) {real, imag} */,
  {32'hbd6ae9d0, 32'h00000000} /* (1, 10, 31) {real, imag} */,
  {32'hbe106550, 32'h00000000} /* (1, 10, 30) {real, imag} */,
  {32'h3e075606, 32'h00000000} /* (1, 10, 29) {real, imag} */,
  {32'hbe414652, 32'h00000000} /* (1, 10, 28) {real, imag} */,
  {32'hbf25318d, 32'h00000000} /* (1, 10, 27) {real, imag} */,
  {32'hbf33ade7, 32'h00000000} /* (1, 10, 26) {real, imag} */,
  {32'hbe8a6779, 32'h00000000} /* (1, 10, 25) {real, imag} */,
  {32'h3da4ec63, 32'h00000000} /* (1, 10, 24) {real, imag} */,
  {32'h3d8af5e1, 32'h00000000} /* (1, 10, 23) {real, imag} */,
  {32'hbe711d06, 32'h00000000} /* (1, 10, 22) {real, imag} */,
  {32'hbeba0d8c, 32'h00000000} /* (1, 10, 21) {real, imag} */,
  {32'h3ecf3dc1, 32'h00000000} /* (1, 10, 20) {real, imag} */,
  {32'h3f31cc14, 32'h00000000} /* (1, 10, 19) {real, imag} */,
  {32'h3e8fe033, 32'h00000000} /* (1, 10, 18) {real, imag} */,
  {32'hbdb71a84, 32'h00000000} /* (1, 10, 17) {real, imag} */,
  {32'h3de2f158, 32'h00000000} /* (1, 10, 16) {real, imag} */,
  {32'hbe064bc9, 32'h00000000} /* (1, 10, 15) {real, imag} */,
  {32'h3be0d440, 32'h00000000} /* (1, 10, 14) {real, imag} */,
  {32'h3ea9cae5, 32'h00000000} /* (1, 10, 13) {real, imag} */,
  {32'hbdff88e4, 32'h00000000} /* (1, 10, 12) {real, imag} */,
  {32'hbd9d3ddd, 32'h00000000} /* (1, 10, 11) {real, imag} */,
  {32'hbe25cb71, 32'h00000000} /* (1, 10, 10) {real, imag} */,
  {32'hbf3075c0, 32'h00000000} /* (1, 10, 9) {real, imag} */,
  {32'hbed19cb8, 32'h00000000} /* (1, 10, 8) {real, imag} */,
  {32'hbe984903, 32'h00000000} /* (1, 10, 7) {real, imag} */,
  {32'h3e66df33, 32'h00000000} /* (1, 10, 6) {real, imag} */,
  {32'hbbe5c39c, 32'h00000000} /* (1, 10, 5) {real, imag} */,
  {32'h3da8bfbb, 32'h00000000} /* (1, 10, 4) {real, imag} */,
  {32'hbe539064, 32'h00000000} /* (1, 10, 3) {real, imag} */,
  {32'hbf38d9ee, 32'h00000000} /* (1, 10, 2) {real, imag} */,
  {32'hbf22b1ac, 32'h00000000} /* (1, 10, 1) {real, imag} */,
  {32'hbe5c8fad, 32'h00000000} /* (1, 10, 0) {real, imag} */,
  {32'hbf2e123b, 32'h00000000} /* (1, 9, 31) {real, imag} */,
  {32'hbf568314, 32'h00000000} /* (1, 9, 30) {real, imag} */,
  {32'hbeb4ebd0, 32'h00000000} /* (1, 9, 29) {real, imag} */,
  {32'hbf16c12e, 32'h00000000} /* (1, 9, 28) {real, imag} */,
  {32'hbf3693e2, 32'h00000000} /* (1, 9, 27) {real, imag} */,
  {32'hbf720168, 32'h00000000} /* (1, 9, 26) {real, imag} */,
  {32'hbf57a004, 32'h00000000} /* (1, 9, 25) {real, imag} */,
  {32'hbf53f50d, 32'h00000000} /* (1, 9, 24) {real, imag} */,
  {32'hbf6b9f96, 32'h00000000} /* (1, 9, 23) {real, imag} */,
  {32'hbf960f77, 32'h00000000} /* (1, 9, 22) {real, imag} */,
  {32'hbf616594, 32'h00000000} /* (1, 9, 21) {real, imag} */,
  {32'h3eed5015, 32'h00000000} /* (1, 9, 20) {real, imag} */,
  {32'h3f8e1401, 32'h00000000} /* (1, 9, 19) {real, imag} */,
  {32'h3e986a31, 32'h00000000} /* (1, 9, 18) {real, imag} */,
  {32'h3dea52fb, 32'h00000000} /* (1, 9, 17) {real, imag} */,
  {32'h3eecbe2e, 32'h00000000} /* (1, 9, 16) {real, imag} */,
  {32'h3f7fa8f5, 32'h00000000} /* (1, 9, 15) {real, imag} */,
  {32'h3f27f7cc, 32'h00000000} /* (1, 9, 14) {real, imag} */,
  {32'h3eeb3f12, 32'h00000000} /* (1, 9, 13) {real, imag} */,
  {32'h3f637b00, 32'h00000000} /* (1, 9, 12) {real, imag} */,
  {32'h3f7ae177, 32'h00000000} /* (1, 9, 11) {real, imag} */,
  {32'hbe8d7968, 32'h00000000} /* (1, 9, 10) {real, imag} */,
  {32'hbf564b5b, 32'h00000000} /* (1, 9, 9) {real, imag} */,
  {32'hbf2eb135, 32'h00000000} /* (1, 9, 8) {real, imag} */,
  {32'hbf6023f5, 32'h00000000} /* (1, 9, 7) {real, imag} */,
  {32'hbea10bc5, 32'h00000000} /* (1, 9, 6) {real, imag} */,
  {32'hbf4ce0b4, 32'h00000000} /* (1, 9, 5) {real, imag} */,
  {32'hbf2b6686, 32'h00000000} /* (1, 9, 4) {real, imag} */,
  {32'hbf5affc1, 32'h00000000} /* (1, 9, 3) {real, imag} */,
  {32'hbfc117b7, 32'h00000000} /* (1, 9, 2) {real, imag} */,
  {32'hbf62296e, 32'h00000000} /* (1, 9, 1) {real, imag} */,
  {32'hbee6345b, 32'h00000000} /* (1, 9, 0) {real, imag} */,
  {32'hbf0d67f2, 32'h00000000} /* (1, 8, 31) {real, imag} */,
  {32'hbf27df5e, 32'h00000000} /* (1, 8, 30) {real, imag} */,
  {32'hbf0c323c, 32'h00000000} /* (1, 8, 29) {real, imag} */,
  {32'hbee95dcb, 32'h00000000} /* (1, 8, 28) {real, imag} */,
  {32'hbe9ecfbb, 32'h00000000} /* (1, 8, 27) {real, imag} */,
  {32'hbf0008a5, 32'h00000000} /* (1, 8, 26) {real, imag} */,
  {32'hbf683495, 32'h00000000} /* (1, 8, 25) {real, imag} */,
  {32'hbfa170da, 32'h00000000} /* (1, 8, 24) {real, imag} */,
  {32'hbfa70783, 32'h00000000} /* (1, 8, 23) {real, imag} */,
  {32'hbfabc7b8, 32'h00000000} /* (1, 8, 22) {real, imag} */,
  {32'hbf03c5a8, 32'h00000000} /* (1, 8, 21) {real, imag} */,
  {32'h3f129ce0, 32'h00000000} /* (1, 8, 20) {real, imag} */,
  {32'h3f520f06, 32'h00000000} /* (1, 8, 19) {real, imag} */,
  {32'h3e92699c, 32'h00000000} /* (1, 8, 18) {real, imag} */,
  {32'h3f283264, 32'h00000000} /* (1, 8, 17) {real, imag} */,
  {32'h3f725a82, 32'h00000000} /* (1, 8, 16) {real, imag} */,
  {32'h3f785c96, 32'h00000000} /* (1, 8, 15) {real, imag} */,
  {32'h3f79173d, 32'h00000000} /* (1, 8, 14) {real, imag} */,
  {32'h3f07234c, 32'h00000000} /* (1, 8, 13) {real, imag} */,
  {32'h3f2e7137, 32'h00000000} /* (1, 8, 12) {real, imag} */,
  {32'h3f0b8638, 32'h00000000} /* (1, 8, 11) {real, imag} */,
  {32'hbf2b60e2, 32'h00000000} /* (1, 8, 10) {real, imag} */,
  {32'hbf487349, 32'h00000000} /* (1, 8, 9) {real, imag} */,
  {32'hbed7ef1d, 32'h00000000} /* (1, 8, 8) {real, imag} */,
  {32'hbf2c01e8, 32'h00000000} /* (1, 8, 7) {real, imag} */,
  {32'hbecabaa1, 32'h00000000} /* (1, 8, 6) {real, imag} */,
  {32'hbf4e72dc, 32'h00000000} /* (1, 8, 5) {real, imag} */,
  {32'hbf789541, 32'h00000000} /* (1, 8, 4) {real, imag} */,
  {32'hbf35f2c2, 32'h00000000} /* (1, 8, 3) {real, imag} */,
  {32'hbfbedffd, 32'h00000000} /* (1, 8, 2) {real, imag} */,
  {32'hbf5ace61, 32'h00000000} /* (1, 8, 1) {real, imag} */,
  {32'hbe0b2dd0, 32'h00000000} /* (1, 8, 0) {real, imag} */,
  {32'hbedb5851, 32'h00000000} /* (1, 7, 31) {real, imag} */,
  {32'hbf29db35, 32'h00000000} /* (1, 7, 30) {real, imag} */,
  {32'hbf2bf656, 32'h00000000} /* (1, 7, 29) {real, imag} */,
  {32'hbf473d4b, 32'h00000000} /* (1, 7, 28) {real, imag} */,
  {32'hbf3493b8, 32'h00000000} /* (1, 7, 27) {real, imag} */,
  {32'hbf937614, 32'h00000000} /* (1, 7, 26) {real, imag} */,
  {32'hbfb27f4c, 32'h00000000} /* (1, 7, 25) {real, imag} */,
  {32'hbfae5c28, 32'h00000000} /* (1, 7, 24) {real, imag} */,
  {32'hbf8e3656, 32'h00000000} /* (1, 7, 23) {real, imag} */,
  {32'hbf830821, 32'h00000000} /* (1, 7, 22) {real, imag} */,
  {32'hbe062408, 32'h00000000} /* (1, 7, 21) {real, imag} */,
  {32'h3f95dfdd, 32'h00000000} /* (1, 7, 20) {real, imag} */,
  {32'h3f1b835e, 32'h00000000} /* (1, 7, 19) {real, imag} */,
  {32'h3f0b06c4, 32'h00000000} /* (1, 7, 18) {real, imag} */,
  {32'h3f856242, 32'h00000000} /* (1, 7, 17) {real, imag} */,
  {32'h3f97a238, 32'h00000000} /* (1, 7, 16) {real, imag} */,
  {32'h3fbba7ca, 32'h00000000} /* (1, 7, 15) {real, imag} */,
  {32'h3fbeba92, 32'h00000000} /* (1, 7, 14) {real, imag} */,
  {32'h3f828b3b, 32'h00000000} /* (1, 7, 13) {real, imag} */,
  {32'h3f34dbc6, 32'h00000000} /* (1, 7, 12) {real, imag} */,
  {32'hbe3c22d0, 32'h00000000} /* (1, 7, 11) {real, imag} */,
  {32'hbf5e150f, 32'h00000000} /* (1, 7, 10) {real, imag} */,
  {32'hbf82dd11, 32'h00000000} /* (1, 7, 9) {real, imag} */,
  {32'hbef32aab, 32'h00000000} /* (1, 7, 8) {real, imag} */,
  {32'hbf2dceab, 32'h00000000} /* (1, 7, 7) {real, imag} */,
  {32'hbf724736, 32'h00000000} /* (1, 7, 6) {real, imag} */,
  {32'hbf9ed858, 32'h00000000} /* (1, 7, 5) {real, imag} */,
  {32'hbfb53397, 32'h00000000} /* (1, 7, 4) {real, imag} */,
  {32'hbf78de15, 32'h00000000} /* (1, 7, 3) {real, imag} */,
  {32'hbfd10298, 32'h00000000} /* (1, 7, 2) {real, imag} */,
  {32'hbf9afc82, 32'h00000000} /* (1, 7, 1) {real, imag} */,
  {32'hbe26847d, 32'h00000000} /* (1, 7, 0) {real, imag} */,
  {32'hbe8cc5ff, 32'h00000000} /* (1, 6, 31) {real, imag} */,
  {32'hbed12a3a, 32'h00000000} /* (1, 6, 30) {real, imag} */,
  {32'hbf17bf82, 32'h00000000} /* (1, 6, 29) {real, imag} */,
  {32'hbf404bfc, 32'h00000000} /* (1, 6, 28) {real, imag} */,
  {32'hbf245f4f, 32'h00000000} /* (1, 6, 27) {real, imag} */,
  {32'hbfbad310, 32'h00000000} /* (1, 6, 26) {real, imag} */,
  {32'hbfb3e3e1, 32'h00000000} /* (1, 6, 25) {real, imag} */,
  {32'hbf73a296, 32'h00000000} /* (1, 6, 24) {real, imag} */,
  {32'hbf0d9b62, 32'h00000000} /* (1, 6, 23) {real, imag} */,
  {32'hbf7cfddb, 32'h00000000} /* (1, 6, 22) {real, imag} */,
  {32'hbf586f79, 32'h00000000} /* (1, 6, 21) {real, imag} */,
  {32'h3fa9f549, 32'h00000000} /* (1, 6, 20) {real, imag} */,
  {32'h3f2147e2, 32'h00000000} /* (1, 6, 19) {real, imag} */,
  {32'h3e918502, 32'h00000000} /* (1, 6, 18) {real, imag} */,
  {32'h3f427f36, 32'h00000000} /* (1, 6, 17) {real, imag} */,
  {32'h3f952c71, 32'h00000000} /* (1, 6, 16) {real, imag} */,
  {32'h3f9fd41d, 32'h00000000} /* (1, 6, 15) {real, imag} */,
  {32'h3f86678b, 32'h00000000} /* (1, 6, 14) {real, imag} */,
  {32'h3f82e7ab, 32'h00000000} /* (1, 6, 13) {real, imag} */,
  {32'h3f930ea5, 32'h00000000} /* (1, 6, 12) {real, imag} */,
  {32'h3ecbc4dc, 32'h00000000} /* (1, 6, 11) {real, imag} */,
  {32'hbee1f626, 32'h00000000} /* (1, 6, 10) {real, imag} */,
  {32'hbfb96043, 32'h00000000} /* (1, 6, 9) {real, imag} */,
  {32'hbf87ed5b, 32'h00000000} /* (1, 6, 8) {real, imag} */,
  {32'hbf30899b, 32'h00000000} /* (1, 6, 7) {real, imag} */,
  {32'hbf3b69d9, 32'h00000000} /* (1, 6, 6) {real, imag} */,
  {32'hbf609827, 32'h00000000} /* (1, 6, 5) {real, imag} */,
  {32'hbf6c65a5, 32'h00000000} /* (1, 6, 4) {real, imag} */,
  {32'hbf473ad7, 32'h00000000} /* (1, 6, 3) {real, imag} */,
  {32'hbf2b7f31, 32'h00000000} /* (1, 6, 2) {real, imag} */,
  {32'hbeb5f408, 32'h00000000} /* (1, 6, 1) {real, imag} */,
  {32'hbe25a6ec, 32'h00000000} /* (1, 6, 0) {real, imag} */,
  {32'hbf3e273a, 32'h00000000} /* (1, 5, 31) {real, imag} */,
  {32'hbf6f6d10, 32'h00000000} /* (1, 5, 30) {real, imag} */,
  {32'hbf4e5179, 32'h00000000} /* (1, 5, 29) {real, imag} */,
  {32'hbf5092f8, 32'h00000000} /* (1, 5, 28) {real, imag} */,
  {32'hbf330567, 32'h00000000} /* (1, 5, 27) {real, imag} */,
  {32'hbfa60250, 32'h00000000} /* (1, 5, 26) {real, imag} */,
  {32'hbf7148ce, 32'h00000000} /* (1, 5, 25) {real, imag} */,
  {32'hbf24d730, 32'h00000000} /* (1, 5, 24) {real, imag} */,
  {32'hbf82757a, 32'h00000000} /* (1, 5, 23) {real, imag} */,
  {32'hbfaea46a, 32'h00000000} /* (1, 5, 22) {real, imag} */,
  {32'hbf63935f, 32'h00000000} /* (1, 5, 21) {real, imag} */,
  {32'h3e7894ec, 32'h00000000} /* (1, 5, 20) {real, imag} */,
  {32'hbd2214c0, 32'h00000000} /* (1, 5, 19) {real, imag} */,
  {32'hbea56b42, 32'h00000000} /* (1, 5, 18) {real, imag} */,
  {32'hbf2384fb, 32'h00000000} /* (1, 5, 17) {real, imag} */,
  {32'hbec51f00, 32'h00000000} /* (1, 5, 16) {real, imag} */,
  {32'h3d57974b, 32'h00000000} /* (1, 5, 15) {real, imag} */,
  {32'h3db1441d, 32'h00000000} /* (1, 5, 14) {real, imag} */,
  {32'h3f21509a, 32'h00000000} /* (1, 5, 13) {real, imag} */,
  {32'h3f927a5a, 32'h00000000} /* (1, 5, 12) {real, imag} */,
  {32'h3f72f179, 32'h00000000} /* (1, 5, 11) {real, imag} */,
  {32'h3e7a0323, 32'h00000000} /* (1, 5, 10) {real, imag} */,
  {32'h3d3be55f, 32'h00000000} /* (1, 5, 9) {real, imag} */,
  {32'hbdc7f8ef, 32'h00000000} /* (1, 5, 8) {real, imag} */,
  {32'hbdb5da34, 32'h00000000} /* (1, 5, 7) {real, imag} */,
  {32'hbe36e2cd, 32'h00000000} /* (1, 5, 6) {real, imag} */,
  {32'hbe7e11fb, 32'h00000000} /* (1, 5, 5) {real, imag} */,
  {32'hbf3bcd60, 32'h00000000} /* (1, 5, 4) {real, imag} */,
  {32'hbf508a84, 32'h00000000} /* (1, 5, 3) {real, imag} */,
  {32'hbf52a695, 32'h00000000} /* (1, 5, 2) {real, imag} */,
  {32'hbf3f337e, 32'h00000000} /* (1, 5, 1) {real, imag} */,
  {32'hbec6f73b, 32'h00000000} /* (1, 5, 0) {real, imag} */,
  {32'hbf461fca, 32'h00000000} /* (1, 4, 31) {real, imag} */,
  {32'hbf86f855, 32'h00000000} /* (1, 4, 30) {real, imag} */,
  {32'hbf7f5458, 32'h00000000} /* (1, 4, 29) {real, imag} */,
  {32'hbf6f3137, 32'h00000000} /* (1, 4, 28) {real, imag} */,
  {32'hbf94574c, 32'h00000000} /* (1, 4, 27) {real, imag} */,
  {32'hbfadc77b, 32'h00000000} /* (1, 4, 26) {real, imag} */,
  {32'hbf9ed57a, 32'h00000000} /* (1, 4, 25) {real, imag} */,
  {32'hbf8e76b7, 32'h00000000} /* (1, 4, 24) {real, imag} */,
  {32'hbf6e42cc, 32'h00000000} /* (1, 4, 23) {real, imag} */,
  {32'hbf33fb9d, 32'h00000000} /* (1, 4, 22) {real, imag} */,
  {32'hbefec7d3, 32'h00000000} /* (1, 4, 21) {real, imag} */,
  {32'hbf6ab936, 32'h00000000} /* (1, 4, 20) {real, imag} */,
  {32'hbf77feb3, 32'h00000000} /* (1, 4, 19) {real, imag} */,
  {32'hbf1619e6, 32'h00000000} /* (1, 4, 18) {real, imag} */,
  {32'hbf861fdb, 32'h00000000} /* (1, 4, 17) {real, imag} */,
  {32'hbf837c3d, 32'h00000000} /* (1, 4, 16) {real, imag} */,
  {32'h3bcc19ce, 32'h00000000} /* (1, 4, 15) {real, imag} */,
  {32'h3e982678, 32'h00000000} /* (1, 4, 14) {real, imag} */,
  {32'h3e551f2f, 32'h00000000} /* (1, 4, 13) {real, imag} */,
  {32'h3ee07adb, 32'h00000000} /* (1, 4, 12) {real, imag} */,
  {32'h3f341e0c, 32'h00000000} /* (1, 4, 11) {real, imag} */,
  {32'h3f65771b, 32'h00000000} /* (1, 4, 10) {real, imag} */,
  {32'h3f8c0103, 32'h00000000} /* (1, 4, 9) {real, imag} */,
  {32'h3f33c077, 32'h00000000} /* (1, 4, 8) {real, imag} */,
  {32'h3f633253, 32'h00000000} /* (1, 4, 7) {real, imag} */,
  {32'h3f17b8a0, 32'h00000000} /* (1, 4, 6) {real, imag} */,
  {32'hbe2967ac, 32'h00000000} /* (1, 4, 5) {real, imag} */,
  {32'hbf1196a6, 32'h00000000} /* (1, 4, 4) {real, imag} */,
  {32'hbf91a6fc, 32'h00000000} /* (1, 4, 3) {real, imag} */,
  {32'hbfaa4e1d, 32'h00000000} /* (1, 4, 2) {real, imag} */,
  {32'hbfa03dfd, 32'h00000000} /* (1, 4, 1) {real, imag} */,
  {32'hbf04a544, 32'h00000000} /* (1, 4, 0) {real, imag} */,
  {32'hbf038719, 32'h00000000} /* (1, 3, 31) {real, imag} */,
  {32'hbf73a70a, 32'h00000000} /* (1, 3, 30) {real, imag} */,
  {32'hbf682969, 32'h00000000} /* (1, 3, 29) {real, imag} */,
  {32'hbf6189dd, 32'h00000000} /* (1, 3, 28) {real, imag} */,
  {32'hbf884f09, 32'h00000000} /* (1, 3, 27) {real, imag} */,
  {32'hbf7ce380, 32'h00000000} /* (1, 3, 26) {real, imag} */,
  {32'hbf90f3b0, 32'h00000000} /* (1, 3, 25) {real, imag} */,
  {32'hbfb9b8b9, 32'h00000000} /* (1, 3, 24) {real, imag} */,
  {32'hbfa52d1c, 32'h00000000} /* (1, 3, 23) {real, imag} */,
  {32'hbf4dddc5, 32'h00000000} /* (1, 3, 22) {real, imag} */,
  {32'hbf12b2b9, 32'h00000000} /* (1, 3, 21) {real, imag} */,
  {32'hbf505493, 32'h00000000} /* (1, 3, 20) {real, imag} */,
  {32'hbfc31876, 32'h00000000} /* (1, 3, 19) {real, imag} */,
  {32'hbfafd472, 32'h00000000} /* (1, 3, 18) {real, imag} */,
  {32'hbf8462a5, 32'h00000000} /* (1, 3, 17) {real, imag} */,
  {32'hbf1ec698, 32'h00000000} /* (1, 3, 16) {real, imag} */,
  {32'h3e58ca0e, 32'h00000000} /* (1, 3, 15) {real, imag} */,
  {32'h3f21ff0c, 32'h00000000} /* (1, 3, 14) {real, imag} */,
  {32'h3f4d0a45, 32'h00000000} /* (1, 3, 13) {real, imag} */,
  {32'h3f140e45, 32'h00000000} /* (1, 3, 12) {real, imag} */,
  {32'h3f6a86d3, 32'h00000000} /* (1, 3, 11) {real, imag} */,
  {32'h3fa4c4d8, 32'h00000000} /* (1, 3, 10) {real, imag} */,
  {32'h3f632941, 32'h00000000} /* (1, 3, 9) {real, imag} */,
  {32'h3f0c79f2, 32'h00000000} /* (1, 3, 8) {real, imag} */,
  {32'h3f2e8ae7, 32'h00000000} /* (1, 3, 7) {real, imag} */,
  {32'h3ece6b64, 32'h00000000} /* (1, 3, 6) {real, imag} */,
  {32'hbf4a1e68, 32'h00000000} /* (1, 3, 5) {real, imag} */,
  {32'hbf31dc7a, 32'h00000000} /* (1, 3, 4) {real, imag} */,
  {32'hbf881b88, 32'h00000000} /* (1, 3, 3) {real, imag} */,
  {32'hbf5eece5, 32'h00000000} /* (1, 3, 2) {real, imag} */,
  {32'hbf3ac35c, 32'h00000000} /* (1, 3, 1) {real, imag} */,
  {32'hbec3e004, 32'h00000000} /* (1, 3, 0) {real, imag} */,
  {32'hbf28a0c4, 32'h00000000} /* (1, 2, 31) {real, imag} */,
  {32'hbf850512, 32'h00000000} /* (1, 2, 30) {real, imag} */,
  {32'hbf84e52e, 32'h00000000} /* (1, 2, 29) {real, imag} */,
  {32'hbfb36ef7, 32'h00000000} /* (1, 2, 28) {real, imag} */,
  {32'hbf735079, 32'h00000000} /* (1, 2, 27) {real, imag} */,
  {32'hbf383592, 32'h00000000} /* (1, 2, 26) {real, imag} */,
  {32'hbf88279a, 32'h00000000} /* (1, 2, 25) {real, imag} */,
  {32'hbf4b9783, 32'h00000000} /* (1, 2, 24) {real, imag} */,
  {32'hbf3783d5, 32'h00000000} /* (1, 2, 23) {real, imag} */,
  {32'hbf2b8049, 32'h00000000} /* (1, 2, 22) {real, imag} */,
  {32'hbee7aab6, 32'h00000000} /* (1, 2, 21) {real, imag} */,
  {32'hbef0eda8, 32'h00000000} /* (1, 2, 20) {real, imag} */,
  {32'hbf842c6c, 32'h00000000} /* (1, 2, 19) {real, imag} */,
  {32'hbfb75c4e, 32'h00000000} /* (1, 2, 18) {real, imag} */,
  {32'hbf961862, 32'h00000000} /* (1, 2, 17) {real, imag} */,
  {32'hbeff4611, 32'h00000000} /* (1, 2, 16) {real, imag} */,
  {32'h3ea6590d, 32'h00000000} /* (1, 2, 15) {real, imag} */,
  {32'h3f62d714, 32'h00000000} /* (1, 2, 14) {real, imag} */,
  {32'h3feb113c, 32'h00000000} /* (1, 2, 13) {real, imag} */,
  {32'h3f9177d6, 32'h00000000} /* (1, 2, 12) {real, imag} */,
  {32'h3f9d82ed, 32'h00000000} /* (1, 2, 11) {real, imag} */,
  {32'h3f9d9ee6, 32'h00000000} /* (1, 2, 10) {real, imag} */,
  {32'h3f9958fd, 32'h00000000} /* (1, 2, 9) {real, imag} */,
  {32'h3f38551f, 32'h00000000} /* (1, 2, 8) {real, imag} */,
  {32'h3eee366a, 32'h00000000} /* (1, 2, 7) {real, imag} */,
  {32'h3f694fdb, 32'h00000000} /* (1, 2, 6) {real, imag} */,
  {32'hbf214fb2, 32'h00000000} /* (1, 2, 5) {real, imag} */,
  {32'hbfd01212, 32'h00000000} /* (1, 2, 4) {real, imag} */,
  {32'hbfae7b5b, 32'h00000000} /* (1, 2, 3) {real, imag} */,
  {32'hbf6f0229, 32'h00000000} /* (1, 2, 2) {real, imag} */,
  {32'hbfbd4455, 32'h00000000} /* (1, 2, 1) {real, imag} */,
  {32'hbf80f043, 32'h00000000} /* (1, 2, 0) {real, imag} */,
  {32'hbf07377e, 32'h00000000} /* (1, 1, 31) {real, imag} */,
  {32'hbf4fbda5, 32'h00000000} /* (1, 1, 30) {real, imag} */,
  {32'hbf21aefc, 32'h00000000} /* (1, 1, 29) {real, imag} */,
  {32'hbf211728, 32'h00000000} /* (1, 1, 28) {real, imag} */,
  {32'hbed06b96, 32'h00000000} /* (1, 1, 27) {real, imag} */,
  {32'hbf1d2883, 32'h00000000} /* (1, 1, 26) {real, imag} */,
  {32'hbf38e77d, 32'h00000000} /* (1, 1, 25) {real, imag} */,
  {32'hbf21a8f7, 32'h00000000} /* (1, 1, 24) {real, imag} */,
  {32'hbf5dda19, 32'h00000000} /* (1, 1, 23) {real, imag} */,
  {32'hbf1840ac, 32'h00000000} /* (1, 1, 22) {real, imag} */,
  {32'hbde22841, 32'h00000000} /* (1, 1, 21) {real, imag} */,
  {32'hbe928925, 32'h00000000} /* (1, 1, 20) {real, imag} */,
  {32'hbf39723f, 32'h00000000} /* (1, 1, 19) {real, imag} */,
  {32'hbf9ca8d5, 32'h00000000} /* (1, 1, 18) {real, imag} */,
  {32'hbf407d85, 32'h00000000} /* (1, 1, 17) {real, imag} */,
  {32'hbed902b4, 32'h00000000} /* (1, 1, 16) {real, imag} */,
  {32'h3ea55fcb, 32'h00000000} /* (1, 1, 15) {real, imag} */,
  {32'h3f90f49a, 32'h00000000} /* (1, 1, 14) {real, imag} */,
  {32'h3fe714d9, 32'h00000000} /* (1, 1, 13) {real, imag} */,
  {32'h3fac4dc5, 32'h00000000} /* (1, 1, 12) {real, imag} */,
  {32'h3fa7d4fb, 32'h00000000} /* (1, 1, 11) {real, imag} */,
  {32'h3f72190b, 32'h00000000} /* (1, 1, 10) {real, imag} */,
  {32'h3f8b8f51, 32'h00000000} /* (1, 1, 9) {real, imag} */,
  {32'h3f7dfe58, 32'h00000000} /* (1, 1, 8) {real, imag} */,
  {32'h3f7c7d3b, 32'h00000000} /* (1, 1, 7) {real, imag} */,
  {32'h3f881903, 32'h00000000} /* (1, 1, 6) {real, imag} */,
  {32'hbf163ed2, 32'h00000000} /* (1, 1, 5) {real, imag} */,
  {32'hc0054996, 32'h00000000} /* (1, 1, 4) {real, imag} */,
  {32'hbfb5408a, 32'h00000000} /* (1, 1, 3) {real, imag} */,
  {32'hbf48e4c8, 32'h00000000} /* (1, 1, 2) {real, imag} */,
  {32'hbf66fd0f, 32'h00000000} /* (1, 1, 1) {real, imag} */,
  {32'hbf26f575, 32'h00000000} /* (1, 1, 0) {real, imag} */,
  {32'hbecf602e, 32'h00000000} /* (1, 0, 31) {real, imag} */,
  {32'hbecbe4f9, 32'h00000000} /* (1, 0, 30) {real, imag} */,
  {32'hbe809869, 32'h00000000} /* (1, 0, 29) {real, imag} */,
  {32'hbe5d0099, 32'h00000000} /* (1, 0, 28) {real, imag} */,
  {32'hbe7ceebe, 32'h00000000} /* (1, 0, 27) {real, imag} */,
  {32'hbec069a9, 32'h00000000} /* (1, 0, 26) {real, imag} */,
  {32'hbdf1647f, 32'h00000000} /* (1, 0, 25) {real, imag} */,
  {32'hbe6033c9, 32'h00000000} /* (1, 0, 24) {real, imag} */,
  {32'hbf8b0a19, 32'h00000000} /* (1, 0, 23) {real, imag} */,
  {32'hbf4aced6, 32'h00000000} /* (1, 0, 22) {real, imag} */,
  {32'hbdf6293e, 32'h00000000} /* (1, 0, 21) {real, imag} */,
  {32'hbe3271dd, 32'h00000000} /* (1, 0, 20) {real, imag} */,
  {32'hbee65d3e, 32'h00000000} /* (1, 0, 19) {real, imag} */,
  {32'hbf109b71, 32'h00000000} /* (1, 0, 18) {real, imag} */,
  {32'hbe500183, 32'h00000000} /* (1, 0, 17) {real, imag} */,
  {32'hbe592c53, 32'h00000000} /* (1, 0, 16) {real, imag} */,
  {32'h3e39e8d3, 32'h00000000} /* (1, 0, 15) {real, imag} */,
  {32'h3f346e9e, 32'h00000000} /* (1, 0, 14) {real, imag} */,
  {32'h3f2c2f1a, 32'h00000000} /* (1, 0, 13) {real, imag} */,
  {32'h3edc1238, 32'h00000000} /* (1, 0, 12) {real, imag} */,
  {32'h3f20ef15, 32'h00000000} /* (1, 0, 11) {real, imag} */,
  {32'h3f222d0b, 32'h00000000} /* (1, 0, 10) {real, imag} */,
  {32'h3eb960c9, 32'h00000000} /* (1, 0, 9) {real, imag} */,
  {32'h3ea5e791, 32'h00000000} /* (1, 0, 8) {real, imag} */,
  {32'h3f1d6cfc, 32'h00000000} /* (1, 0, 7) {real, imag} */,
  {32'h3f0f7030, 32'h00000000} /* (1, 0, 6) {real, imag} */,
  {32'hbeab60eb, 32'h00000000} /* (1, 0, 5) {real, imag} */,
  {32'hbf30afea, 32'h00000000} /* (1, 0, 4) {real, imag} */,
  {32'hbf22c1cc, 32'h00000000} /* (1, 0, 3) {real, imag} */,
  {32'hbf335594, 32'h00000000} /* (1, 0, 2) {real, imag} */,
  {32'hbf11b1ef, 32'h00000000} /* (1, 0, 1) {real, imag} */,
  {32'hbed10649, 32'h00000000} /* (1, 0, 0) {real, imag} */,
  {32'hbd87055d, 32'h00000000} /* (0, 31, 31) {real, imag} */,
  {32'hbdd7bb82, 32'h00000000} /* (0, 31, 30) {real, imag} */,
  {32'hbf4b7326, 32'h00000000} /* (0, 31, 29) {real, imag} */,
  {32'hbf7d7ff4, 32'h00000000} /* (0, 31, 28) {real, imag} */,
  {32'hbe74afad, 32'h00000000} /* (0, 31, 27) {real, imag} */,
  {32'hbd06df04, 32'h00000000} /* (0, 31, 26) {real, imag} */,
  {32'hbc5f2ed1, 32'h00000000} /* (0, 31, 25) {real, imag} */,
  {32'hbe159a94, 32'h00000000} /* (0, 31, 24) {real, imag} */,
  {32'hbe74d139, 32'h00000000} /* (0, 31, 23) {real, imag} */,
  {32'hbe73a809, 32'h00000000} /* (0, 31, 22) {real, imag} */,
  {32'hbe0ca029, 32'h00000000} /* (0, 31, 21) {real, imag} */,
  {32'h3d43dbf5, 32'h00000000} /* (0, 31, 20) {real, imag} */,
  {32'h3d8451cb, 32'h00000000} /* (0, 31, 19) {real, imag} */,
  {32'hbda23c08, 32'h00000000} /* (0, 31, 18) {real, imag} */,
  {32'hbe0df703, 32'h00000000} /* (0, 31, 17) {real, imag} */,
  {32'hbc84e35c, 32'h00000000} /* (0, 31, 16) {real, imag} */,
  {32'h3e057069, 32'h00000000} /* (0, 31, 15) {real, imag} */,
  {32'h3ed960cf, 32'h00000000} /* (0, 31, 14) {real, imag} */,
  {32'h3e3c4edc, 32'h00000000} /* (0, 31, 13) {real, imag} */,
  {32'h3e0282ec, 32'h00000000} /* (0, 31, 12) {real, imag} */,
  {32'h3ec68f33, 32'h00000000} /* (0, 31, 11) {real, imag} */,
  {32'h3df62d8e, 32'h00000000} /* (0, 31, 10) {real, imag} */,
  {32'h3d063932, 32'h00000000} /* (0, 31, 9) {real, imag} */,
  {32'hbcc029c0, 32'h00000000} /* (0, 31, 8) {real, imag} */,
  {32'hbd2c9312, 32'h00000000} /* (0, 31, 7) {real, imag} */,
  {32'hbd881107, 32'h00000000} /* (0, 31, 6) {real, imag} */,
  {32'hbeaccfe1, 32'h00000000} /* (0, 31, 5) {real, imag} */,
  {32'hbeb99293, 32'h00000000} /* (0, 31, 4) {real, imag} */,
  {32'hbe59f497, 32'h00000000} /* (0, 31, 3) {real, imag} */,
  {32'hbd9b9227, 32'h00000000} /* (0, 31, 2) {real, imag} */,
  {32'hbc192d82, 32'h00000000} /* (0, 31, 1) {real, imag} */,
  {32'hbc77d5cb, 32'h00000000} /* (0, 31, 0) {real, imag} */,
  {32'hbeae23fc, 32'h00000000} /* (0, 30, 31) {real, imag} */,
  {32'hbc51feb0, 32'h00000000} /* (0, 30, 30) {real, imag} */,
  {32'hbf22ff0b, 32'h00000000} /* (0, 30, 29) {real, imag} */,
  {32'hbf81cbbe, 32'h00000000} /* (0, 30, 28) {real, imag} */,
  {32'hbeaade16, 32'h00000000} /* (0, 30, 27) {real, imag} */,
  {32'hbde53b9c, 32'h00000000} /* (0, 30, 26) {real, imag} */,
  {32'hbe8afc5e, 32'h00000000} /* (0, 30, 25) {real, imag} */,
  {32'hbf083d84, 32'h00000000} /* (0, 30, 24) {real, imag} */,
  {32'hbec9b637, 32'h00000000} /* (0, 30, 23) {real, imag} */,
  {32'hbe586710, 32'h00000000} /* (0, 30, 22) {real, imag} */,
  {32'hbd8486ad, 32'h00000000} /* (0, 30, 21) {real, imag} */,
  {32'h3ea4ed67, 32'h00000000} /* (0, 30, 20) {real, imag} */,
  {32'h3bfa7740, 32'h00000000} /* (0, 30, 19) {real, imag} */,
  {32'hbe2ec77d, 32'h00000000} /* (0, 30, 18) {real, imag} */,
  {32'h3e1ca67e, 32'h00000000} /* (0, 30, 17) {real, imag} */,
  {32'h3f091743, 32'h00000000} /* (0, 30, 16) {real, imag} */,
  {32'h3e1f353e, 32'h00000000} /* (0, 30, 15) {real, imag} */,
  {32'h3ea7d688, 32'h00000000} /* (0, 30, 14) {real, imag} */,
  {32'h3dbda3cf, 32'h00000000} /* (0, 30, 13) {real, imag} */,
  {32'h3db82b38, 32'h00000000} /* (0, 30, 12) {real, imag} */,
  {32'h3e9e3fa6, 32'h00000000} /* (0, 30, 11) {real, imag} */,
  {32'hbdae3f8b, 32'h00000000} /* (0, 30, 10) {real, imag} */,
  {32'hbe2b09c4, 32'h00000000} /* (0, 30, 9) {real, imag} */,
  {32'hbe9ac7a3, 32'h00000000} /* (0, 30, 8) {real, imag} */,
  {32'hbea070f5, 32'h00000000} /* (0, 30, 7) {real, imag} */,
  {32'hbebbb41e, 32'h00000000} /* (0, 30, 6) {real, imag} */,
  {32'hbf3adc8c, 32'h00000000} /* (0, 30, 5) {real, imag} */,
  {32'hbf31b779, 32'h00000000} /* (0, 30, 4) {real, imag} */,
  {32'hbf1d05ce, 32'h00000000} /* (0, 30, 3) {real, imag} */,
  {32'hbedbbebf, 32'h00000000} /* (0, 30, 2) {real, imag} */,
  {32'h3daadc8f, 32'h00000000} /* (0, 30, 1) {real, imag} */,
  {32'hbda66e63, 32'h00000000} /* (0, 30, 0) {real, imag} */,
  {32'hbf0835a7, 32'h00000000} /* (0, 29, 31) {real, imag} */,
  {32'hbe94d856, 32'h00000000} /* (0, 29, 30) {real, imag} */,
  {32'hbf228925, 32'h00000000} /* (0, 29, 29) {real, imag} */,
  {32'hbf21b880, 32'h00000000} /* (0, 29, 28) {real, imag} */,
  {32'hbe0c8ae8, 32'h00000000} /* (0, 29, 27) {real, imag} */,
  {32'hbe908808, 32'h00000000} /* (0, 29, 26) {real, imag} */,
  {32'hbeedac05, 32'h00000000} /* (0, 29, 25) {real, imag} */,
  {32'hbf19fafe, 32'h00000000} /* (0, 29, 24) {real, imag} */,
  {32'hbf099fe9, 32'h00000000} /* (0, 29, 23) {real, imag} */,
  {32'hbe8161c7, 32'h00000000} /* (0, 29, 22) {real, imag} */,
  {32'hbe862a53, 32'h00000000} /* (0, 29, 21) {real, imag} */,
  {32'h3dd2806b, 32'h00000000} /* (0, 29, 20) {real, imag} */,
  {32'h3d3b3206, 32'h00000000} /* (0, 29, 19) {real, imag} */,
  {32'h3d72c698, 32'h00000000} /* (0, 29, 18) {real, imag} */,
  {32'h3ed4f29f, 32'h00000000} /* (0, 29, 17) {real, imag} */,
  {32'h3f24cf6b, 32'h00000000} /* (0, 29, 16) {real, imag} */,
  {32'h3ea1bf28, 32'h00000000} /* (0, 29, 15) {real, imag} */,
  {32'h3f36c9b3, 32'h00000000} /* (0, 29, 14) {real, imag} */,
  {32'h3f01cfe9, 32'h00000000} /* (0, 29, 13) {real, imag} */,
  {32'h3ee7dd1e, 32'h00000000} /* (0, 29, 12) {real, imag} */,
  {32'h3ed7f9e9, 32'h00000000} /* (0, 29, 11) {real, imag} */,
  {32'hbeb36a19, 32'h00000000} /* (0, 29, 10) {real, imag} */,
  {32'hbf23bc2a, 32'h00000000} /* (0, 29, 9) {real, imag} */,
  {32'hbf022f17, 32'h00000000} /* (0, 29, 8) {real, imag} */,
  {32'hbefd7ca5, 32'h00000000} /* (0, 29, 7) {real, imag} */,
  {32'hbef83131, 32'h00000000} /* (0, 29, 6) {real, imag} */,
  {32'hbf49ed15, 32'h00000000} /* (0, 29, 5) {real, imag} */,
  {32'hbf1071cd, 32'h00000000} /* (0, 29, 4) {real, imag} */,
  {32'hbf0448c2, 32'h00000000} /* (0, 29, 3) {real, imag} */,
  {32'hbed9c0f5, 32'h00000000} /* (0, 29, 2) {real, imag} */,
  {32'hbe05aff2, 32'h00000000} /* (0, 29, 1) {real, imag} */,
  {32'hbea63862, 32'h00000000} /* (0, 29, 0) {real, imag} */,
  {32'hbeca1ff2, 32'h00000000} /* (0, 28, 31) {real, imag} */,
  {32'hbf19aa38, 32'h00000000} /* (0, 28, 30) {real, imag} */,
  {32'hbf489358, 32'h00000000} /* (0, 28, 29) {real, imag} */,
  {32'hbed7c108, 32'h00000000} /* (0, 28, 28) {real, imag} */,
  {32'h3d4e24cc, 32'h00000000} /* (0, 28, 27) {real, imag} */,
  {32'hbe94efb6, 32'h00000000} /* (0, 28, 26) {real, imag} */,
  {32'hbe8be512, 32'h00000000} /* (0, 28, 25) {real, imag} */,
  {32'hbe2ce58d, 32'h00000000} /* (0, 28, 24) {real, imag} */,
  {32'hbee3da44, 32'h00000000} /* (0, 28, 23) {real, imag} */,
  {32'hbed34ec6, 32'h00000000} /* (0, 28, 22) {real, imag} */,
  {32'hbe9e94d5, 32'h00000000} /* (0, 28, 21) {real, imag} */,
  {32'h3de89ece, 32'h00000000} /* (0, 28, 20) {real, imag} */,
  {32'h3efce3a8, 32'h00000000} /* (0, 28, 19) {real, imag} */,
  {32'h3f076b86, 32'h00000000} /* (0, 28, 18) {real, imag} */,
  {32'h3eee1419, 32'h00000000} /* (0, 28, 17) {real, imag} */,
  {32'h3eac82dd, 32'h00000000} /* (0, 28, 16) {real, imag} */,
  {32'h3e5d0bad, 32'h00000000} /* (0, 28, 15) {real, imag} */,
  {32'h3ebafd9e, 32'h00000000} /* (0, 28, 14) {real, imag} */,
  {32'h3ef7ab63, 32'h00000000} /* (0, 28, 13) {real, imag} */,
  {32'h3f2962ca, 32'h00000000} /* (0, 28, 12) {real, imag} */,
  {32'h3f0110f0, 32'h00000000} /* (0, 28, 11) {real, imag} */,
  {32'hbe9ca15a, 32'h00000000} /* (0, 28, 10) {real, imag} */,
  {32'hbf020e2d, 32'h00000000} /* (0, 28, 9) {real, imag} */,
  {32'hbed51bf1, 32'h00000000} /* (0, 28, 8) {real, imag} */,
  {32'hbe9d8fac, 32'h00000000} /* (0, 28, 7) {real, imag} */,
  {32'hbea9a1a6, 32'h00000000} /* (0, 28, 6) {real, imag} */,
  {32'hbf377937, 32'h00000000} /* (0, 28, 5) {real, imag} */,
  {32'hbedc0a87, 32'h00000000} /* (0, 28, 4) {real, imag} */,
  {32'hbec8ae5e, 32'h00000000} /* (0, 28, 3) {real, imag} */,
  {32'hbe99b507, 32'h00000000} /* (0, 28, 2) {real, imag} */,
  {32'hbe818b41, 32'h00000000} /* (0, 28, 1) {real, imag} */,
  {32'hbecc83bc, 32'h00000000} /* (0, 28, 0) {real, imag} */,
  {32'hbe32b32a, 32'h00000000} /* (0, 27, 31) {real, imag} */,
  {32'hbf270295, 32'h00000000} /* (0, 27, 30) {real, imag} */,
  {32'hbf526c18, 32'h00000000} /* (0, 27, 29) {real, imag} */,
  {32'hbf058505, 32'h00000000} /* (0, 27, 28) {real, imag} */,
  {32'hbddfa386, 32'h00000000} /* (0, 27, 27) {real, imag} */,
  {32'hbe89603a, 32'h00000000} /* (0, 27, 26) {real, imag} */,
  {32'hbe9b3268, 32'h00000000} /* (0, 27, 25) {real, imag} */,
  {32'hbe845839, 32'h00000000} /* (0, 27, 24) {real, imag} */,
  {32'hbf2a6183, 32'h00000000} /* (0, 27, 23) {real, imag} */,
  {32'hbf01ddc4, 32'h00000000} /* (0, 27, 22) {real, imag} */,
  {32'hbdab0b7a, 32'h00000000} /* (0, 27, 21) {real, imag} */,
  {32'h3e8b3514, 32'h00000000} /* (0, 27, 20) {real, imag} */,
  {32'h3ec4b206, 32'h00000000} /* (0, 27, 19) {real, imag} */,
  {32'h3eff9426, 32'h00000000} /* (0, 27, 18) {real, imag} */,
  {32'h3f0f9526, 32'h00000000} /* (0, 27, 17) {real, imag} */,
  {32'h3e19610d, 32'h00000000} /* (0, 27, 16) {real, imag} */,
  {32'h3e3f763c, 32'h00000000} /* (0, 27, 15) {real, imag} */,
  {32'h3e87b266, 32'h00000000} /* (0, 27, 14) {real, imag} */,
  {32'h3e85c7f3, 32'h00000000} /* (0, 27, 13) {real, imag} */,
  {32'h3ec41dbd, 32'h00000000} /* (0, 27, 12) {real, imag} */,
  {32'h3ef7854a, 32'h00000000} /* (0, 27, 11) {real, imag} */,
  {32'h3ca7dd23, 32'h00000000} /* (0, 27, 10) {real, imag} */,
  {32'hbe130f53, 32'h00000000} /* (0, 27, 9) {real, imag} */,
  {32'hbe903c46, 32'h00000000} /* (0, 27, 8) {real, imag} */,
  {32'hbe160ea9, 32'h00000000} /* (0, 27, 7) {real, imag} */,
  {32'hbe7f4570, 32'h00000000} /* (0, 27, 6) {real, imag} */,
  {32'hbf021e05, 32'h00000000} /* (0, 27, 5) {real, imag} */,
  {32'hbee8d6e1, 32'h00000000} /* (0, 27, 4) {real, imag} */,
  {32'hbe60a91c, 32'h00000000} /* (0, 27, 3) {real, imag} */,
  {32'hbe595d56, 32'h00000000} /* (0, 27, 2) {real, imag} */,
  {32'hbe9b9d76, 32'h00000000} /* (0, 27, 1) {real, imag} */,
  {32'hbe98b845, 32'h00000000} /* (0, 27, 0) {real, imag} */,
  {32'hbeaf53d1, 32'h00000000} /* (0, 26, 31) {real, imag} */,
  {32'hbf85fad8, 32'h00000000} /* (0, 26, 30) {real, imag} */,
  {32'hbf748198, 32'h00000000} /* (0, 26, 29) {real, imag} */,
  {32'hbeb60b5c, 32'h00000000} /* (0, 26, 28) {real, imag} */,
  {32'hbe1158af, 32'h00000000} /* (0, 26, 27) {real, imag} */,
  {32'hbeef0969, 32'h00000000} /* (0, 26, 26) {real, imag} */,
  {32'hbed7cadb, 32'h00000000} /* (0, 26, 25) {real, imag} */,
  {32'hbe51329c, 32'h00000000} /* (0, 26, 24) {real, imag} */,
  {32'hbf247589, 32'h00000000} /* (0, 26, 23) {real, imag} */,
  {32'hbf24203d, 32'h00000000} /* (0, 26, 22) {real, imag} */,
  {32'hbe61028e, 32'h00000000} /* (0, 26, 21) {real, imag} */,
  {32'h3e8f5a06, 32'h00000000} /* (0, 26, 20) {real, imag} */,
  {32'h3f321ed7, 32'h00000000} /* (0, 26, 19) {real, imag} */,
  {32'h3ef18fba, 32'h00000000} /* (0, 26, 18) {real, imag} */,
  {32'h3ec27530, 32'h00000000} /* (0, 26, 17) {real, imag} */,
  {32'h3ea4bd76, 32'h00000000} /* (0, 26, 16) {real, imag} */,
  {32'h3ea60986, 32'h00000000} /* (0, 26, 15) {real, imag} */,
  {32'h3ee260b6, 32'h00000000} /* (0, 26, 14) {real, imag} */,
  {32'h3e4ca492, 32'h00000000} /* (0, 26, 13) {real, imag} */,
  {32'h3ea07daf, 32'h00000000} /* (0, 26, 12) {real, imag} */,
  {32'h3f0a51b4, 32'h00000000} /* (0, 26, 11) {real, imag} */,
  {32'hbd7c2b08, 32'h00000000} /* (0, 26, 10) {real, imag} */,
  {32'hbf42ea23, 32'h00000000} /* (0, 26, 9) {real, imag} */,
  {32'hbf04a7f2, 32'h00000000} /* (0, 26, 8) {real, imag} */,
  {32'hbe4b5c7b, 32'h00000000} /* (0, 26, 7) {real, imag} */,
  {32'hbeb785a9, 32'h00000000} /* (0, 26, 6) {real, imag} */,
  {32'hbea9c318, 32'h00000000} /* (0, 26, 5) {real, imag} */,
  {32'hbefe96de, 32'h00000000} /* (0, 26, 4) {real, imag} */,
  {32'hbf15b061, 32'h00000000} /* (0, 26, 3) {real, imag} */,
  {32'hbf02f512, 32'h00000000} /* (0, 26, 2) {real, imag} */,
  {32'hbf1a4c69, 32'h00000000} /* (0, 26, 1) {real, imag} */,
  {32'hbec2cc30, 32'h00000000} /* (0, 26, 0) {real, imag} */,
  {32'hbe93b497, 32'h00000000} /* (0, 25, 31) {real, imag} */,
  {32'hbf7a9215, 32'h00000000} /* (0, 25, 30) {real, imag} */,
  {32'hbf90f507, 32'h00000000} /* (0, 25, 29) {real, imag} */,
  {32'hbf009e86, 32'h00000000} /* (0, 25, 28) {real, imag} */,
  {32'hbddf4f2f, 32'h00000000} /* (0, 25, 27) {real, imag} */,
  {32'hbe949d61, 32'h00000000} /* (0, 25, 26) {real, imag} */,
  {32'hbe86f2e7, 32'h00000000} /* (0, 25, 25) {real, imag} */,
  {32'hbcd61d38, 32'h00000000} /* (0, 25, 24) {real, imag} */,
  {32'hbe656635, 32'h00000000} /* (0, 25, 23) {real, imag} */,
  {32'hbead0a8b, 32'h00000000} /* (0, 25, 22) {real, imag} */,
  {32'hbe29939c, 32'h00000000} /* (0, 25, 21) {real, imag} */,
  {32'h3f457b83, 32'h00000000} /* (0, 25, 20) {real, imag} */,
  {32'h3fa63896, 32'h00000000} /* (0, 25, 19) {real, imag} */,
  {32'h3f467903, 32'h00000000} /* (0, 25, 18) {real, imag} */,
  {32'h3e8b5287, 32'h00000000} /* (0, 25, 17) {real, imag} */,
  {32'h3f619552, 32'h00000000} /* (0, 25, 16) {real, imag} */,
  {32'h3f359a2b, 32'h00000000} /* (0, 25, 15) {real, imag} */,
  {32'h3eda83ec, 32'h00000000} /* (0, 25, 14) {real, imag} */,
  {32'h3e7b2552, 32'h00000000} /* (0, 25, 13) {real, imag} */,
  {32'h3e18b255, 32'h00000000} /* (0, 25, 12) {real, imag} */,
  {32'h3d9a0be3, 32'h00000000} /* (0, 25, 11) {real, imag} */,
  {32'hbeafdbc9, 32'h00000000} /* (0, 25, 10) {real, imag} */,
  {32'hbfca5c68, 32'h00000000} /* (0, 25, 9) {real, imag} */,
  {32'hbfc09e58, 32'h00000000} /* (0, 25, 8) {real, imag} */,
  {32'hbf3a81e1, 32'h00000000} /* (0, 25, 7) {real, imag} */,
  {32'hbe89136e, 32'h00000000} /* (0, 25, 6) {real, imag} */,
  {32'hbe6232b0, 32'h00000000} /* (0, 25, 5) {real, imag} */,
  {32'hbf3624d9, 32'h00000000} /* (0, 25, 4) {real, imag} */,
  {32'hbf55095a, 32'h00000000} /* (0, 25, 3) {real, imag} */,
  {32'hbf2f467c, 32'h00000000} /* (0, 25, 2) {real, imag} */,
  {32'hbf67a700, 32'h00000000} /* (0, 25, 1) {real, imag} */,
  {32'hbf0cb674, 32'h00000000} /* (0, 25, 0) {real, imag} */,
  {32'hbe238b48, 32'h00000000} /* (0, 24, 31) {real, imag} */,
  {32'hbe607455, 32'h00000000} /* (0, 24, 30) {real, imag} */,
  {32'hbe2647d5, 32'h00000000} /* (0, 24, 29) {real, imag} */,
  {32'hbdcc090f, 32'h00000000} /* (0, 24, 28) {real, imag} */,
  {32'hbe0a2cab, 32'h00000000} /* (0, 24, 27) {real, imag} */,
  {32'hbe65c767, 32'h00000000} /* (0, 24, 26) {real, imag} */,
  {32'hbd324917, 32'h00000000} /* (0, 24, 25) {real, imag} */,
  {32'hbde4b090, 32'h00000000} /* (0, 24, 24) {real, imag} */,
  {32'hbe0c5243, 32'h00000000} /* (0, 24, 23) {real, imag} */,
  {32'hbe97c478, 32'h00000000} /* (0, 24, 22) {real, imag} */,
  {32'hbe6f025d, 32'h00000000} /* (0, 24, 21) {real, imag} */,
  {32'h3f3ea593, 32'h00000000} /* (0, 24, 20) {real, imag} */,
  {32'h3f344995, 32'h00000000} /* (0, 24, 19) {real, imag} */,
  {32'h3f12a025, 32'h00000000} /* (0, 24, 18) {real, imag} */,
  {32'h3e5d9da6, 32'h00000000} /* (0, 24, 17) {real, imag} */,
  {32'h3ed0b717, 32'h00000000} /* (0, 24, 16) {real, imag} */,
  {32'h3ea91564, 32'h00000000} /* (0, 24, 15) {real, imag} */,
  {32'h3f27cf0d, 32'h00000000} /* (0, 24, 14) {real, imag} */,
  {32'h3f33d79c, 32'h00000000} /* (0, 24, 13) {real, imag} */,
  {32'h3e0b1413, 32'h00000000} /* (0, 24, 12) {real, imag} */,
  {32'h3e174f0e, 32'h00000000} /* (0, 24, 11) {real, imag} */,
  {32'hbe9e869a, 32'h00000000} /* (0, 24, 10) {real, imag} */,
  {32'hbf53911b, 32'h00000000} /* (0, 24, 9) {real, imag} */,
  {32'hbf848622, 32'h00000000} /* (0, 24, 8) {real, imag} */,
  {32'hbec43f80, 32'h00000000} /* (0, 24, 7) {real, imag} */,
  {32'hbdee68d0, 32'h00000000} /* (0, 24, 6) {real, imag} */,
  {32'hbe62bd4e, 32'h00000000} /* (0, 24, 5) {real, imag} */,
  {32'hbea8d748, 32'h00000000} /* (0, 24, 4) {real, imag} */,
  {32'hbeccf0dd, 32'h00000000} /* (0, 24, 3) {real, imag} */,
  {32'hbeeefe9a, 32'h00000000} /* (0, 24, 2) {real, imag} */,
  {32'hbed5c89d, 32'h00000000} /* (0, 24, 1) {real, imag} */,
  {32'hbeb03883, 32'h00000000} /* (0, 24, 0) {real, imag} */,
  {32'hbe30daf3, 32'h00000000} /* (0, 23, 31) {real, imag} */,
  {32'hbe8193b2, 32'h00000000} /* (0, 23, 30) {real, imag} */,
  {32'hbe3605d7, 32'h00000000} /* (0, 23, 29) {real, imag} */,
  {32'hbedbd6bb, 32'h00000000} /* (0, 23, 28) {real, imag} */,
  {32'hbee90690, 32'h00000000} /* (0, 23, 27) {real, imag} */,
  {32'hbed93246, 32'h00000000} /* (0, 23, 26) {real, imag} */,
  {32'h3cde46c6, 32'h00000000} /* (0, 23, 25) {real, imag} */,
  {32'hbc96cb9e, 32'h00000000} /* (0, 23, 24) {real, imag} */,
  {32'hbdfe2995, 32'h00000000} /* (0, 23, 23) {real, imag} */,
  {32'hbea2a6a8, 32'h00000000} /* (0, 23, 22) {real, imag} */,
  {32'hbbd88190, 32'h00000000} /* (0, 23, 21) {real, imag} */,
  {32'h3f23d6c4, 32'h00000000} /* (0, 23, 20) {real, imag} */,
  {32'h3e979a20, 32'h00000000} /* (0, 23, 19) {real, imag} */,
  {32'h3e48a069, 32'h00000000} /* (0, 23, 18) {real, imag} */,
  {32'h3de9b9e1, 32'h00000000} /* (0, 23, 17) {real, imag} */,
  {32'h3e65c3bc, 32'h00000000} /* (0, 23, 16) {real, imag} */,
  {32'h3de7f70a, 32'h00000000} /* (0, 23, 15) {real, imag} */,
  {32'h3e3fc103, 32'h00000000} /* (0, 23, 14) {real, imag} */,
  {32'h3f0b2d71, 32'h00000000} /* (0, 23, 13) {real, imag} */,
  {32'h3f0a3f02, 32'h00000000} /* (0, 23, 12) {real, imag} */,
  {32'h3f02cbf7, 32'h00000000} /* (0, 23, 11) {real, imag} */,
  {32'hbdea0a79, 32'h00000000} /* (0, 23, 10) {real, imag} */,
  {32'hbe05a000, 32'h00000000} /* (0, 23, 9) {real, imag} */,
  {32'hbea0faac, 32'h00000000} /* (0, 23, 8) {real, imag} */,
  {32'hbe61df8c, 32'h00000000} /* (0, 23, 7) {real, imag} */,
  {32'hbd7003a0, 32'h00000000} /* (0, 23, 6) {real, imag} */,
  {32'hbea380e8, 32'h00000000} /* (0, 23, 5) {real, imag} */,
  {32'hbf055b77, 32'h00000000} /* (0, 23, 4) {real, imag} */,
  {32'hbe216348, 32'h00000000} /* (0, 23, 3) {real, imag} */,
  {32'hbe5e1f4f, 32'h00000000} /* (0, 23, 2) {real, imag} */,
  {32'hbe539842, 32'h00000000} /* (0, 23, 1) {real, imag} */,
  {32'hbc989282, 32'h00000000} /* (0, 23, 0) {real, imag} */,
  {32'hbe1176e7, 32'h00000000} /* (0, 22, 31) {real, imag} */,
  {32'hbd8f58e3, 32'h00000000} /* (0, 22, 30) {real, imag} */,
  {32'hbe8f7687, 32'h00000000} /* (0, 22, 29) {real, imag} */,
  {32'hbf61f683, 32'h00000000} /* (0, 22, 28) {real, imag} */,
  {32'hbf5c72fb, 32'h00000000} /* (0, 22, 27) {real, imag} */,
  {32'hbf033fec, 32'h00000000} /* (0, 22, 26) {real, imag} */,
  {32'hbea7f953, 32'h00000000} /* (0, 22, 25) {real, imag} */,
  {32'hbeb40bf8, 32'h00000000} /* (0, 22, 24) {real, imag} */,
  {32'hbe94105d, 32'h00000000} /* (0, 22, 23) {real, imag} */,
  {32'hbe9dd6a9, 32'h00000000} /* (0, 22, 22) {real, imag} */,
  {32'hbd9757a9, 32'h00000000} /* (0, 22, 21) {real, imag} */,
  {32'h3ebd2cec, 32'h00000000} /* (0, 22, 20) {real, imag} */,
  {32'h3e299975, 32'h00000000} /* (0, 22, 19) {real, imag} */,
  {32'h3b8974bc, 32'h00000000} /* (0, 22, 18) {real, imag} */,
  {32'h3be45546, 32'h00000000} /* (0, 22, 17) {real, imag} */,
  {32'h3e735d40, 32'h00000000} /* (0, 22, 16) {real, imag} */,
  {32'h3e39e5ac, 32'h00000000} /* (0, 22, 15) {real, imag} */,
  {32'h3da87e0a, 32'h00000000} /* (0, 22, 14) {real, imag} */,
  {32'h3f587287, 32'h00000000} /* (0, 22, 13) {real, imag} */,
  {32'h3f548da8, 32'h00000000} /* (0, 22, 12) {real, imag} */,
  {32'h3f142e39, 32'h00000000} /* (0, 22, 11) {real, imag} */,
  {32'hbd5fc3b8, 32'h00000000} /* (0, 22, 10) {real, imag} */,
  {32'hbe94b062, 32'h00000000} /* (0, 22, 9) {real, imag} */,
  {32'hbd0844d8, 32'h00000000} /* (0, 22, 8) {real, imag} */,
  {32'hbe3daf93, 32'h00000000} /* (0, 22, 7) {real, imag} */,
  {32'hbe604e84, 32'h00000000} /* (0, 22, 6) {real, imag} */,
  {32'hbe905df6, 32'h00000000} /* (0, 22, 5) {real, imag} */,
  {32'hbe9bed5c, 32'h00000000} /* (0, 22, 4) {real, imag} */,
  {32'hbd489a16, 32'h00000000} /* (0, 22, 3) {real, imag} */,
  {32'hbe64ee8e, 32'h00000000} /* (0, 22, 2) {real, imag} */,
  {32'hbe078bea, 32'h00000000} /* (0, 22, 1) {real, imag} */,
  {32'hbcb41770, 32'h00000000} /* (0, 22, 0) {real, imag} */,
  {32'hbe56c078, 32'h00000000} /* (0, 21, 31) {real, imag} */,
  {32'hbda2545c, 32'h00000000} /* (0, 21, 30) {real, imag} */,
  {32'hbd79b4e9, 32'h00000000} /* (0, 21, 29) {real, imag} */,
  {32'hbf4b3c77, 32'h00000000} /* (0, 21, 28) {real, imag} */,
  {32'hbecda548, 32'h00000000} /* (0, 21, 27) {real, imag} */,
  {32'h3cbe1f21, 32'h00000000} /* (0, 21, 26) {real, imag} */,
  {32'hbe30de7b, 32'h00000000} /* (0, 21, 25) {real, imag} */,
  {32'hbed47dba, 32'h00000000} /* (0, 21, 24) {real, imag} */,
  {32'hbe03ec7b, 32'h00000000} /* (0, 21, 23) {real, imag} */,
  {32'hbe095bba, 32'h00000000} /* (0, 21, 22) {real, imag} */,
  {32'hbe5dcb5b, 32'h00000000} /* (0, 21, 21) {real, imag} */,
  {32'hbe4a353a, 32'h00000000} /* (0, 21, 20) {real, imag} */,
  {32'hbde82d2d, 32'h00000000} /* (0, 21, 19) {real, imag} */,
  {32'h3e5ac72c, 32'h00000000} /* (0, 21, 18) {real, imag} */,
  {32'hbd007cb7, 32'h00000000} /* (0, 21, 17) {real, imag} */,
  {32'h3cd5ac4c, 32'h00000000} /* (0, 21, 16) {real, imag} */,
  {32'hbb79c010, 32'h00000000} /* (0, 21, 15) {real, imag} */,
  {32'hbd184858, 32'h00000000} /* (0, 21, 14) {real, imag} */,
  {32'h3f10b804, 32'h00000000} /* (0, 21, 13) {real, imag} */,
  {32'h3ef2289d, 32'h00000000} /* (0, 21, 12) {real, imag} */,
  {32'h3ebfae96, 32'h00000000} /* (0, 21, 11) {real, imag} */,
  {32'hbe74eeeb, 32'h00000000} /* (0, 21, 10) {real, imag} */,
  {32'hbe501da2, 32'h00000000} /* (0, 21, 9) {real, imag} */,
  {32'h3e8a144a, 32'h00000000} /* (0, 21, 8) {real, imag} */,
  {32'hbe171fa9, 32'h00000000} /* (0, 21, 7) {real, imag} */,
  {32'hbe19791e, 32'h00000000} /* (0, 21, 6) {real, imag} */,
  {32'hbdbf6f7a, 32'h00000000} /* (0, 21, 5) {real, imag} */,
  {32'h3d02465b, 32'h00000000} /* (0, 21, 4) {real, imag} */,
  {32'h3d59b10b, 32'h00000000} /* (0, 21, 3) {real, imag} */,
  {32'hbda59c30, 32'h00000000} /* (0, 21, 2) {real, imag} */,
  {32'hbe7fcb73, 32'h00000000} /* (0, 21, 1) {real, imag} */,
  {32'hbe6d48a5, 32'h00000000} /* (0, 21, 0) {real, imag} */,
  {32'h3df3caef, 32'h00000000} /* (0, 20, 31) {real, imag} */,
  {32'h3e8f1909, 32'h00000000} /* (0, 20, 30) {real, imag} */,
  {32'h3ed7ee96, 32'h00000000} /* (0, 20, 29) {real, imag} */,
  {32'h3dffd6db, 32'h00000000} /* (0, 20, 28) {real, imag} */,
  {32'h3e703126, 32'h00000000} /* (0, 20, 27) {real, imag} */,
  {32'h3eb79e95, 32'h00000000} /* (0, 20, 26) {real, imag} */,
  {32'h3f610dbc, 32'h00000000} /* (0, 20, 25) {real, imag} */,
  {32'h3f22f7ee, 32'h00000000} /* (0, 20, 24) {real, imag} */,
  {32'h3ea00ad4, 32'h00000000} /* (0, 20, 23) {real, imag} */,
  {32'h3ea4966e, 32'h00000000} /* (0, 20, 22) {real, imag} */,
  {32'h3e238be3, 32'h00000000} /* (0, 20, 21) {real, imag} */,
  {32'hbec5912c, 32'h00000000} /* (0, 20, 20) {real, imag} */,
  {32'hbf1747c6, 32'h00000000} /* (0, 20, 19) {real, imag} */,
  {32'hbe1deb82, 32'h00000000} /* (0, 20, 18) {real, imag} */,
  {32'hbe68ed1a, 32'h00000000} /* (0, 20, 17) {real, imag} */,
  {32'hbdd04dac, 32'h00000000} /* (0, 20, 16) {real, imag} */,
  {32'hbf0b2b14, 32'h00000000} /* (0, 20, 15) {real, imag} */,
  {32'hbef1a4a8, 32'h00000000} /* (0, 20, 14) {real, imag} */,
  {32'hbdb4891b, 32'h00000000} /* (0, 20, 13) {real, imag} */,
  {32'h3d62b5e1, 32'h00000000} /* (0, 20, 12) {real, imag} */,
  {32'hbc7be15c, 32'h00000000} /* (0, 20, 11) {real, imag} */,
  {32'hbe9be110, 32'h00000000} /* (0, 20, 10) {real, imag} */,
  {32'h3e4890c6, 32'h00000000} /* (0, 20, 9) {real, imag} */,
  {32'h3ee05d83, 32'h00000000} /* (0, 20, 8) {real, imag} */,
  {32'h3e978540, 32'h00000000} /* (0, 20, 7) {real, imag} */,
  {32'h3ea69478, 32'h00000000} /* (0, 20, 6) {real, imag} */,
  {32'h3e8b3e70, 32'h00000000} /* (0, 20, 5) {real, imag} */,
  {32'h3ecc6b65, 32'h00000000} /* (0, 20, 4) {real, imag} */,
  {32'h3ea4586a, 32'h00000000} /* (0, 20, 3) {real, imag} */,
  {32'h3e952316, 32'h00000000} /* (0, 20, 2) {real, imag} */,
  {32'h3d41694d, 32'h00000000} /* (0, 20, 1) {real, imag} */,
  {32'hbdac4efb, 32'h00000000} /* (0, 20, 0) {real, imag} */,
  {32'h3ed19bfc, 32'h00000000} /* (0, 19, 31) {real, imag} */,
  {32'h3f5b0890, 32'h00000000} /* (0, 19, 30) {real, imag} */,
  {32'h3f2da6e5, 32'h00000000} /* (0, 19, 29) {real, imag} */,
  {32'h3e15f797, 32'h00000000} /* (0, 19, 28) {real, imag} */,
  {32'h3eadce1e, 32'h00000000} /* (0, 19, 27) {real, imag} */,
  {32'h3ebf11c6, 32'h00000000} /* (0, 19, 26) {real, imag} */,
  {32'h3f1f0b2b, 32'h00000000} /* (0, 19, 25) {real, imag} */,
  {32'h3f16344d, 32'h00000000} /* (0, 19, 24) {real, imag} */,
  {32'h3e61d6b8, 32'h00000000} /* (0, 19, 23) {real, imag} */,
  {32'h3e8993ae, 32'h00000000} /* (0, 19, 22) {real, imag} */,
  {32'h3e9fde5f, 32'h00000000} /* (0, 19, 21) {real, imag} */,
  {32'hbd521d4c, 32'h00000000} /* (0, 19, 20) {real, imag} */,
  {32'hbe4c0b42, 32'h00000000} /* (0, 19, 19) {real, imag} */,
  {32'hbe58c782, 32'h00000000} /* (0, 19, 18) {real, imag} */,
  {32'hbeb12dc1, 32'h00000000} /* (0, 19, 17) {real, imag} */,
  {32'hbdec2ff3, 32'h00000000} /* (0, 19, 16) {real, imag} */,
  {32'hbe43ff43, 32'h00000000} /* (0, 19, 15) {real, imag} */,
  {32'hbe940045, 32'h00000000} /* (0, 19, 14) {real, imag} */,
  {32'hbdc70798, 32'h00000000} /* (0, 19, 13) {real, imag} */,
  {32'hbe80449e, 32'h00000000} /* (0, 19, 12) {real, imag} */,
  {32'hbf000f71, 32'h00000000} /* (0, 19, 11) {real, imag} */,
  {32'hbe2b437c, 32'h00000000} /* (0, 19, 10) {real, imag} */,
  {32'h3ea38e85, 32'h00000000} /* (0, 19, 9) {real, imag} */,
  {32'h3ec4c432, 32'h00000000} /* (0, 19, 8) {real, imag} */,
  {32'h3f33ec97, 32'h00000000} /* (0, 19, 7) {real, imag} */,
  {32'h3f075d6c, 32'h00000000} /* (0, 19, 6) {real, imag} */,
  {32'h3f1bbbd1, 32'h00000000} /* (0, 19, 5) {real, imag} */,
  {32'h3f567876, 32'h00000000} /* (0, 19, 4) {real, imag} */,
  {32'h3f0701e6, 32'h00000000} /* (0, 19, 3) {real, imag} */,
  {32'h3eb0535e, 32'h00000000} /* (0, 19, 2) {real, imag} */,
  {32'h3ed202f4, 32'h00000000} /* (0, 19, 1) {real, imag} */,
  {32'h3e224598, 32'h00000000} /* (0, 19, 0) {real, imag} */,
  {32'h3e684c8b, 32'h00000000} /* (0, 18, 31) {real, imag} */,
  {32'h3f14a8c4, 32'h00000000} /* (0, 18, 30) {real, imag} */,
  {32'h3eb35f21, 32'h00000000} /* (0, 18, 29) {real, imag} */,
  {32'h3d3730c6, 32'h00000000} /* (0, 18, 28) {real, imag} */,
  {32'h3e8cb912, 32'h00000000} /* (0, 18, 27) {real, imag} */,
  {32'h3f009479, 32'h00000000} /* (0, 18, 26) {real, imag} */,
  {32'h3ed9b6c0, 32'h00000000} /* (0, 18, 25) {real, imag} */,
  {32'h3f374d4e, 32'h00000000} /* (0, 18, 24) {real, imag} */,
  {32'h3eb12a89, 32'h00000000} /* (0, 18, 23) {real, imag} */,
  {32'h3e43fed5, 32'h00000000} /* (0, 18, 22) {real, imag} */,
  {32'h3dbbf345, 32'h00000000} /* (0, 18, 21) {real, imag} */,
  {32'hbcc51208, 32'h00000000} /* (0, 18, 20) {real, imag} */,
  {32'hbe380a97, 32'h00000000} /* (0, 18, 19) {real, imag} */,
  {32'hbeff975a, 32'h00000000} /* (0, 18, 18) {real, imag} */,
  {32'hbf0baf75, 32'h00000000} /* (0, 18, 17) {real, imag} */,
  {32'hbcf2399e, 32'h00000000} /* (0, 18, 16) {real, imag} */,
  {32'hbcc29e3d, 32'h00000000} /* (0, 18, 15) {real, imag} */,
  {32'hbebf88dc, 32'h00000000} /* (0, 18, 14) {real, imag} */,
  {32'hbf391fe9, 32'h00000000} /* (0, 18, 13) {real, imag} */,
  {32'hbf3680b5, 32'h00000000} /* (0, 18, 12) {real, imag} */,
  {32'hbefc59c3, 32'h00000000} /* (0, 18, 11) {real, imag} */,
  {32'h3df2365d, 32'h00000000} /* (0, 18, 10) {real, imag} */,
  {32'h3dec8016, 32'h00000000} /* (0, 18, 9) {real, imag} */,
  {32'h3e7d7eb9, 32'h00000000} /* (0, 18, 8) {real, imag} */,
  {32'h3f3555d0, 32'h00000000} /* (0, 18, 7) {real, imag} */,
  {32'h3f1fdf3e, 32'h00000000} /* (0, 18, 6) {real, imag} */,
  {32'h3f36c826, 32'h00000000} /* (0, 18, 5) {real, imag} */,
  {32'h3f22ebb5, 32'h00000000} /* (0, 18, 4) {real, imag} */,
  {32'h3f1965cb, 32'h00000000} /* (0, 18, 3) {real, imag} */,
  {32'h3f028193, 32'h00000000} /* (0, 18, 2) {real, imag} */,
  {32'h3eeb3cc4, 32'h00000000} /* (0, 18, 1) {real, imag} */,
  {32'h3e3f119b, 32'h00000000} /* (0, 18, 0) {real, imag} */,
  {32'h3e8b6423, 32'h00000000} /* (0, 17, 31) {real, imag} */,
  {32'h3ed3acc9, 32'h00000000} /* (0, 17, 30) {real, imag} */,
  {32'h3eadc8d5, 32'h00000000} /* (0, 17, 29) {real, imag} */,
  {32'h3f1c20aa, 32'h00000000} /* (0, 17, 28) {real, imag} */,
  {32'h3f028559, 32'h00000000} /* (0, 17, 27) {real, imag} */,
  {32'h3f094bbf, 32'h00000000} /* (0, 17, 26) {real, imag} */,
  {32'h3f1eea44, 32'h00000000} /* (0, 17, 25) {real, imag} */,
  {32'h3f0fb9e6, 32'h00000000} /* (0, 17, 24) {real, imag} */,
  {32'h3eb7cee9, 32'h00000000} /* (0, 17, 23) {real, imag} */,
  {32'h3ec4bd16, 32'h00000000} /* (0, 17, 22) {real, imag} */,
  {32'h3d526da4, 32'h00000000} /* (0, 17, 21) {real, imag} */,
  {32'h3d88c430, 32'h00000000} /* (0, 17, 20) {real, imag} */,
  {32'hbd945ced, 32'h00000000} /* (0, 17, 19) {real, imag} */,
  {32'hbee2b8c7, 32'h00000000} /* (0, 17, 18) {real, imag} */,
  {32'hbf34c3ca, 32'h00000000} /* (0, 17, 17) {real, imag} */,
  {32'hbe8d8515, 32'h00000000} /* (0, 17, 16) {real, imag} */,
  {32'hbea13aea, 32'h00000000} /* (0, 17, 15) {real, imag} */,
  {32'hbe79ed87, 32'h00000000} /* (0, 17, 14) {real, imag} */,
  {32'hbf02329c, 32'h00000000} /* (0, 17, 13) {real, imag} */,
  {32'hbf19e9c9, 32'h00000000} /* (0, 17, 12) {real, imag} */,
  {32'hbe712dc3, 32'h00000000} /* (0, 17, 11) {real, imag} */,
  {32'h3f0d2180, 32'h00000000} /* (0, 17, 10) {real, imag} */,
  {32'h3f1d50f7, 32'h00000000} /* (0, 17, 9) {real, imag} */,
  {32'h3ebf566f, 32'h00000000} /* (0, 17, 8) {real, imag} */,
  {32'h3f03c9d6, 32'h00000000} /* (0, 17, 7) {real, imag} */,
  {32'h3f2b39d7, 32'h00000000} /* (0, 17, 6) {real, imag} */,
  {32'h3e96d09f, 32'h00000000} /* (0, 17, 5) {real, imag} */,
  {32'h3e0f0b53, 32'h00000000} /* (0, 17, 4) {real, imag} */,
  {32'h3de113dd, 32'h00000000} /* (0, 17, 3) {real, imag} */,
  {32'h3e070b0b, 32'h00000000} /* (0, 17, 2) {real, imag} */,
  {32'h3e7fc19d, 32'h00000000} /* (0, 17, 1) {real, imag} */,
  {32'h3e745c6d, 32'h00000000} /* (0, 17, 0) {real, imag} */,
  {32'h3d7e5f1d, 32'h00000000} /* (0, 16, 31) {real, imag} */,
  {32'h3ee344fc, 32'h00000000} /* (0, 16, 30) {real, imag} */,
  {32'h3f384abc, 32'h00000000} /* (0, 16, 29) {real, imag} */,
  {32'h3f5de899, 32'h00000000} /* (0, 16, 28) {real, imag} */,
  {32'h3f4cfc21, 32'h00000000} /* (0, 16, 27) {real, imag} */,
  {32'h3ee509e8, 32'h00000000} /* (0, 16, 26) {real, imag} */,
  {32'h3f06d398, 32'h00000000} /* (0, 16, 25) {real, imag} */,
  {32'h3e93d66b, 32'h00000000} /* (0, 16, 24) {real, imag} */,
  {32'h3e93b668, 32'h00000000} /* (0, 16, 23) {real, imag} */,
  {32'h3f1a3aee, 32'h00000000} /* (0, 16, 22) {real, imag} */,
  {32'h3e811515, 32'h00000000} /* (0, 16, 21) {real, imag} */,
  {32'h3d4b5ba4, 32'h00000000} /* (0, 16, 20) {real, imag} */,
  {32'hbd64ce23, 32'h00000000} /* (0, 16, 19) {real, imag} */,
  {32'h3c58ed52, 32'h00000000} /* (0, 16, 18) {real, imag} */,
  {32'hbf00923d, 32'h00000000} /* (0, 16, 17) {real, imag} */,
  {32'hbee5d164, 32'h00000000} /* (0, 16, 16) {real, imag} */,
  {32'hbf0d3129, 32'h00000000} /* (0, 16, 15) {real, imag} */,
  {32'hbef3c4a3, 32'h00000000} /* (0, 16, 14) {real, imag} */,
  {32'hbf2c1961, 32'h00000000} /* (0, 16, 13) {real, imag} */,
  {32'hbf3cd4ae, 32'h00000000} /* (0, 16, 12) {real, imag} */,
  {32'hbe9da5a0, 32'h00000000} /* (0, 16, 11) {real, imag} */,
  {32'h3eedf4b5, 32'h00000000} /* (0, 16, 10) {real, imag} */,
  {32'h3fb70842, 32'h00000000} /* (0, 16, 9) {real, imag} */,
  {32'h3f814c5f, 32'h00000000} /* (0, 16, 8) {real, imag} */,
  {32'h3f41904e, 32'h00000000} /* (0, 16, 7) {real, imag} */,
  {32'h3f3de1f1, 32'h00000000} /* (0, 16, 6) {real, imag} */,
  {32'h3e913242, 32'h00000000} /* (0, 16, 5) {real, imag} */,
  {32'h3de94a5c, 32'h00000000} /* (0, 16, 4) {real, imag} */,
  {32'h3d3a4150, 32'h00000000} /* (0, 16, 3) {real, imag} */,
  {32'h3e0a33a6, 32'h00000000} /* (0, 16, 2) {real, imag} */,
  {32'h3e9b9f03, 32'h00000000} /* (0, 16, 1) {real, imag} */,
  {32'h3e5417b6, 32'h00000000} /* (0, 16, 0) {real, imag} */,
  {32'h3e2af295, 32'h00000000} /* (0, 15, 31) {real, imag} */,
  {32'h3ecf8a53, 32'h00000000} /* (0, 15, 30) {real, imag} */,
  {32'h3f370bec, 32'h00000000} /* (0, 15, 29) {real, imag} */,
  {32'h3f194cb9, 32'h00000000} /* (0, 15, 28) {real, imag} */,
  {32'h3f01ae6f, 32'h00000000} /* (0, 15, 27) {real, imag} */,
  {32'h3ea6b419, 32'h00000000} /* (0, 15, 26) {real, imag} */,
  {32'h3e30d31a, 32'h00000000} /* (0, 15, 25) {real, imag} */,
  {32'h3d8333eb, 32'h00000000} /* (0, 15, 24) {real, imag} */,
  {32'h3e0ccc68, 32'h00000000} /* (0, 15, 23) {real, imag} */,
  {32'h3e52c456, 32'h00000000} /* (0, 15, 22) {real, imag} */,
  {32'h3e243e7b, 32'h00000000} /* (0, 15, 21) {real, imag} */,
  {32'hbdc9b20d, 32'h00000000} /* (0, 15, 20) {real, imag} */,
  {32'hbe2043f4, 32'h00000000} /* (0, 15, 19) {real, imag} */,
  {32'hbd26777f, 32'h00000000} /* (0, 15, 18) {real, imag} */,
  {32'hbe5e89ee, 32'h00000000} /* (0, 15, 17) {real, imag} */,
  {32'hbe8a58bd, 32'h00000000} /* (0, 15, 16) {real, imag} */,
  {32'hbf1b7ec6, 32'h00000000} /* (0, 15, 15) {real, imag} */,
  {32'hbf32b010, 32'h00000000} /* (0, 15, 14) {real, imag} */,
  {32'hbf846b78, 32'h00000000} /* (0, 15, 13) {real, imag} */,
  {32'hbfb8c6b3, 32'h00000000} /* (0, 15, 12) {real, imag} */,
  {32'hbf4bd456, 32'h00000000} /* (0, 15, 11) {real, imag} */,
  {32'hbdbfca88, 32'h00000000} /* (0, 15, 10) {real, imag} */,
  {32'h3f0da8fb, 32'h00000000} /* (0, 15, 9) {real, imag} */,
  {32'h3e530010, 32'h00000000} /* (0, 15, 8) {real, imag} */,
  {32'h3e9ab263, 32'h00000000} /* (0, 15, 7) {real, imag} */,
  {32'h3f4b52e1, 32'h00000000} /* (0, 15, 6) {real, imag} */,
  {32'h3f4d7279, 32'h00000000} /* (0, 15, 5) {real, imag} */,
  {32'h3f4723ce, 32'h00000000} /* (0, 15, 4) {real, imag} */,
  {32'h3ef62282, 32'h00000000} /* (0, 15, 3) {real, imag} */,
  {32'h3f3ecf0b, 32'h00000000} /* (0, 15, 2) {real, imag} */,
  {32'h3f17688a, 32'h00000000} /* (0, 15, 1) {real, imag} */,
  {32'h3e00c81d, 32'h00000000} /* (0, 15, 0) {real, imag} */,
  {32'h3dfa0f39, 32'h00000000} /* (0, 14, 31) {real, imag} */,
  {32'h3e92e9d5, 32'h00000000} /* (0, 14, 30) {real, imag} */,
  {32'h3ed3129a, 32'h00000000} /* (0, 14, 29) {real, imag} */,
  {32'h3eacbab2, 32'h00000000} /* (0, 14, 28) {real, imag} */,
  {32'h3eb9a138, 32'h00000000} /* (0, 14, 27) {real, imag} */,
  {32'h3ee6571a, 32'h00000000} /* (0, 14, 26) {real, imag} */,
  {32'h3e84062d, 32'h00000000} /* (0, 14, 25) {real, imag} */,
  {32'h3df99e31, 32'h00000000} /* (0, 14, 24) {real, imag} */,
  {32'h3e964745, 32'h00000000} /* (0, 14, 23) {real, imag} */,
  {32'h3e632958, 32'h00000000} /* (0, 14, 22) {real, imag} */,
  {32'hbd946b42, 32'h00000000} /* (0, 14, 21) {real, imag} */,
  {32'hbea76b12, 32'h00000000} /* (0, 14, 20) {real, imag} */,
  {32'hbec60d13, 32'h00000000} /* (0, 14, 19) {real, imag} */,
  {32'hbf09ec53, 32'h00000000} /* (0, 14, 18) {real, imag} */,
  {32'hbf3538fe, 32'h00000000} /* (0, 14, 17) {real, imag} */,
  {32'hbe526055, 32'h00000000} /* (0, 14, 16) {real, imag} */,
  {32'hbe8f9c7b, 32'h00000000} /* (0, 14, 15) {real, imag} */,
  {32'hbec7de49, 32'h00000000} /* (0, 14, 14) {real, imag} */,
  {32'hbf1254f2, 32'h00000000} /* (0, 14, 13) {real, imag} */,
  {32'hbf2e154d, 32'h00000000} /* (0, 14, 12) {real, imag} */,
  {32'hbebb5e6a, 32'h00000000} /* (0, 14, 11) {real, imag} */,
  {32'hbd8e1759, 32'h00000000} /* (0, 14, 10) {real, imag} */,
  {32'h3da14797, 32'h00000000} /* (0, 14, 9) {real, imag} */,
  {32'h3db7d6d8, 32'h00000000} /* (0, 14, 8) {real, imag} */,
  {32'h3e8188c1, 32'h00000000} /* (0, 14, 7) {real, imag} */,
  {32'h3ec8647e, 32'h00000000} /* (0, 14, 6) {real, imag} */,
  {32'h3f42b890, 32'h00000000} /* (0, 14, 5) {real, imag} */,
  {32'h3f60360d, 32'h00000000} /* (0, 14, 4) {real, imag} */,
  {32'h3f3b5967, 32'h00000000} /* (0, 14, 3) {real, imag} */,
  {32'h3f24fa4e, 32'h00000000} /* (0, 14, 2) {real, imag} */,
  {32'h3eea4a4a, 32'h00000000} /* (0, 14, 1) {real, imag} */,
  {32'h3ddd5f08, 32'h00000000} /* (0, 14, 0) {real, imag} */,
  {32'h3d0ddc0a, 32'h00000000} /* (0, 13, 31) {real, imag} */,
  {32'h3e7748f3, 32'h00000000} /* (0, 13, 30) {real, imag} */,
  {32'h3ef9144f, 32'h00000000} /* (0, 13, 29) {real, imag} */,
  {32'h3ed8f224, 32'h00000000} /* (0, 13, 28) {real, imag} */,
  {32'h3f097e25, 32'h00000000} /* (0, 13, 27) {real, imag} */,
  {32'h3f145d28, 32'h00000000} /* (0, 13, 26) {real, imag} */,
  {32'h3f059e24, 32'h00000000} /* (0, 13, 25) {real, imag} */,
  {32'h3df52e47, 32'h00000000} /* (0, 13, 24) {real, imag} */,
  {32'h3e4dce0e, 32'h00000000} /* (0, 13, 23) {real, imag} */,
  {32'h3ed3fc03, 32'h00000000} /* (0, 13, 22) {real, imag} */,
  {32'hbe0cbb75, 32'h00000000} /* (0, 13, 21) {real, imag} */,
  {32'hbf27df2e, 32'h00000000} /* (0, 13, 20) {real, imag} */,
  {32'hbf31e191, 32'h00000000} /* (0, 13, 19) {real, imag} */,
  {32'hbf331036, 32'h00000000} /* (0, 13, 18) {real, imag} */,
  {32'hbf32ffe7, 32'h00000000} /* (0, 13, 17) {real, imag} */,
  {32'hbf1ed6c7, 32'h00000000} /* (0, 13, 16) {real, imag} */,
  {32'hbd7a1c89, 32'h00000000} /* (0, 13, 15) {real, imag} */,
  {32'hbc5453af, 32'h00000000} /* (0, 13, 14) {real, imag} */,
  {32'hbe1819d8, 32'h00000000} /* (0, 13, 13) {real, imag} */,
  {32'hbeb8bac2, 32'h00000000} /* (0, 13, 12) {real, imag} */,
  {32'hbee9a508, 32'h00000000} /* (0, 13, 11) {real, imag} */,
  {32'hbe6298c4, 32'h00000000} /* (0, 13, 10) {real, imag} */,
  {32'h3d8a30d8, 32'h00000000} /* (0, 13, 9) {real, imag} */,
  {32'h3ea1a029, 32'h00000000} /* (0, 13, 8) {real, imag} */,
  {32'h3f44a6a6, 32'h00000000} /* (0, 13, 7) {real, imag} */,
  {32'h3e93a64f, 32'h00000000} /* (0, 13, 6) {real, imag} */,
  {32'h3ecee577, 32'h00000000} /* (0, 13, 5) {real, imag} */,
  {32'h3ed21a55, 32'h00000000} /* (0, 13, 4) {real, imag} */,
  {32'h3ed1a26e, 32'h00000000} /* (0, 13, 3) {real, imag} */,
  {32'h3ef89b15, 32'h00000000} /* (0, 13, 2) {real, imag} */,
  {32'h3f01ccc5, 32'h00000000} /* (0, 13, 1) {real, imag} */,
  {32'h3e3583ed, 32'h00000000} /* (0, 13, 0) {real, imag} */,
  {32'h3dc87ae6, 32'h00000000} /* (0, 12, 31) {real, imag} */,
  {32'h3e4f5667, 32'h00000000} /* (0, 12, 30) {real, imag} */,
  {32'h3e3a47a8, 32'h00000000} /* (0, 12, 29) {real, imag} */,
  {32'h3ee4e82c, 32'h00000000} /* (0, 12, 28) {real, imag} */,
  {32'h3ec1c51b, 32'h00000000} /* (0, 12, 27) {real, imag} */,
  {32'h3e81ea7a, 32'h00000000} /* (0, 12, 26) {real, imag} */,
  {32'h3eeaf943, 32'h00000000} /* (0, 12, 25) {real, imag} */,
  {32'h3ed3139b, 32'h00000000} /* (0, 12, 24) {real, imag} */,
  {32'h3eb62f9e, 32'h00000000} /* (0, 12, 23) {real, imag} */,
  {32'h3f07262f, 32'h00000000} /* (0, 12, 22) {real, imag} */,
  {32'h3f07e92f, 32'h00000000} /* (0, 12, 21) {real, imag} */,
  {32'hbe5db915, 32'h00000000} /* (0, 12, 20) {real, imag} */,
  {32'hbf00043e, 32'h00000000} /* (0, 12, 19) {real, imag} */,
  {32'hbeb49a07, 32'h00000000} /* (0, 12, 18) {real, imag} */,
  {32'hbef920de, 32'h00000000} /* (0, 12, 17) {real, imag} */,
  {32'hbf139b9c, 32'h00000000} /* (0, 12, 16) {real, imag} */,
  {32'h3c848309, 32'h00000000} /* (0, 12, 15) {real, imag} */,
  {32'hbdfa4a94, 32'h00000000} /* (0, 12, 14) {real, imag} */,
  {32'hbe1a2d0e, 32'h00000000} /* (0, 12, 13) {real, imag} */,
  {32'hbda25ae7, 32'h00000000} /* (0, 12, 12) {real, imag} */,
  {32'hbe6ccc0f, 32'h00000000} /* (0, 12, 11) {real, imag} */,
  {32'hbd9b5792, 32'h00000000} /* (0, 12, 10) {real, imag} */,
  {32'h3cdb7186, 32'h00000000} /* (0, 12, 9) {real, imag} */,
  {32'h3e5e003e, 32'h00000000} /* (0, 12, 8) {real, imag} */,
  {32'h3f443e90, 32'h00000000} /* (0, 12, 7) {real, imag} */,
  {32'h3ef2ac11, 32'h00000000} /* (0, 12, 6) {real, imag} */,
  {32'h3f1f02af, 32'h00000000} /* (0, 12, 5) {real, imag} */,
  {32'h3ee2a8bc, 32'h00000000} /* (0, 12, 4) {real, imag} */,
  {32'h3e0649b8, 32'h00000000} /* (0, 12, 3) {real, imag} */,
  {32'h3e9b7010, 32'h00000000} /* (0, 12, 2) {real, imag} */,
  {32'h3efbd5ad, 32'h00000000} /* (0, 12, 1) {real, imag} */,
  {32'h3e11c008, 32'h00000000} /* (0, 12, 0) {real, imag} */,
  {32'h3daee46c, 32'h00000000} /* (0, 11, 31) {real, imag} */,
  {32'h3d3922a7, 32'h00000000} /* (0, 11, 30) {real, imag} */,
  {32'h3e4eb9c7, 32'h00000000} /* (0, 11, 29) {real, imag} */,
  {32'h3e930f34, 32'h00000000} /* (0, 11, 28) {real, imag} */,
  {32'h3df942c6, 32'h00000000} /* (0, 11, 27) {real, imag} */,
  {32'hbc9f46ef, 32'h00000000} /* (0, 11, 26) {real, imag} */,
  {32'h3e647ea0, 32'h00000000} /* (0, 11, 25) {real, imag} */,
  {32'h3eec21b8, 32'h00000000} /* (0, 11, 24) {real, imag} */,
  {32'h3e1e21aa, 32'h00000000} /* (0, 11, 23) {real, imag} */,
  {32'h3eabf29d, 32'h00000000} /* (0, 11, 22) {real, imag} */,
  {32'h3ef16577, 32'h00000000} /* (0, 11, 21) {real, imag} */,
  {32'hbd3d691c, 32'h00000000} /* (0, 11, 20) {real, imag} */,
  {32'hbdfbd1ec, 32'h00000000} /* (0, 11, 19) {real, imag} */,
  {32'hbea32c1f, 32'h00000000} /* (0, 11, 18) {real, imag} */,
  {32'hbf3a6ea2, 32'h00000000} /* (0, 11, 17) {real, imag} */,
  {32'hbead3349, 32'h00000000} /* (0, 11, 16) {real, imag} */,
  {32'hbe629801, 32'h00000000} /* (0, 11, 15) {real, imag} */,
  {32'hbea69594, 32'h00000000} /* (0, 11, 14) {real, imag} */,
  {32'hbe7ae88c, 32'h00000000} /* (0, 11, 13) {real, imag} */,
  {32'hbe378ce9, 32'h00000000} /* (0, 11, 12) {real, imag} */,
  {32'hbe6eb37d, 32'h00000000} /* (0, 11, 11) {real, imag} */,
  {32'hbdfd515c, 32'h00000000} /* (0, 11, 10) {real, imag} */,
  {32'hbd9fd2f4, 32'h00000000} /* (0, 11, 9) {real, imag} */,
  {32'h3e2ed12a, 32'h00000000} /* (0, 11, 8) {real, imag} */,
  {32'h3ef632e1, 32'h00000000} /* (0, 11, 7) {real, imag} */,
  {32'h3eff8afc, 32'h00000000} /* (0, 11, 6) {real, imag} */,
  {32'h3f051675, 32'h00000000} /* (0, 11, 5) {real, imag} */,
  {32'h3eaf30af, 32'h00000000} /* (0, 11, 4) {real, imag} */,
  {32'hbcd7bc9a, 32'h00000000} /* (0, 11, 3) {real, imag} */,
  {32'h3bc16eca, 32'h00000000} /* (0, 11, 2) {real, imag} */,
  {32'h3dcf3384, 32'h00000000} /* (0, 11, 1) {real, imag} */,
  {32'h3d06a74a, 32'h00000000} /* (0, 11, 0) {real, imag} */,
  {32'h3ba48e58, 32'h00000000} /* (0, 10, 31) {real, imag} */,
  {32'hbe96b6c2, 32'h00000000} /* (0, 10, 30) {real, imag} */,
  {32'h3d345daf, 32'h00000000} /* (0, 10, 29) {real, imag} */,
  {32'hbe048017, 32'h00000000} /* (0, 10, 28) {real, imag} */,
  {32'hbf370ddd, 32'h00000000} /* (0, 10, 27) {real, imag} */,
  {32'hbefcd066, 32'h00000000} /* (0, 10, 26) {real, imag} */,
  {32'hbde021ff, 32'h00000000} /* (0, 10, 25) {real, imag} */,
  {32'hbd50c68a, 32'h00000000} /* (0, 10, 24) {real, imag} */,
  {32'hbece8089, 32'h00000000} /* (0, 10, 23) {real, imag} */,
  {32'hbefc958e, 32'h00000000} /* (0, 10, 22) {real, imag} */,
  {32'hbf015b83, 32'h00000000} /* (0, 10, 21) {real, imag} */,
  {32'h3ea54e0f, 32'h00000000} /* (0, 10, 20) {real, imag} */,
  {32'h3ecb2853, 32'h00000000} /* (0, 10, 19) {real, imag} */,
  {32'h3d34d847, 32'h00000000} /* (0, 10, 18) {real, imag} */,
  {32'h3cf25d20, 32'h00000000} /* (0, 10, 17) {real, imag} */,
  {32'h3e4f9dd0, 32'h00000000} /* (0, 10, 16) {real, imag} */,
  {32'hbe994287, 32'h00000000} /* (0, 10, 15) {real, imag} */,
  {32'hbdca28bc, 32'h00000000} /* (0, 10, 14) {real, imag} */,
  {32'hbd312edc, 32'h00000000} /* (0, 10, 13) {real, imag} */,
  {32'h3d13f0a6, 32'h00000000} /* (0, 10, 12) {real, imag} */,
  {32'hbd4446de, 32'h00000000} /* (0, 10, 11) {real, imag} */,
  {32'hbe7520ad, 32'h00000000} /* (0, 10, 10) {real, imag} */,
  {32'hbf004421, 32'h00000000} /* (0, 10, 9) {real, imag} */,
  {32'hbe8535fc, 32'h00000000} /* (0, 10, 8) {real, imag} */,
  {32'hbe9b935a, 32'h00000000} /* (0, 10, 7) {real, imag} */,
  {32'h3d703524, 32'h00000000} /* (0, 10, 6) {real, imag} */,
  {32'hbe2b5161, 32'h00000000} /* (0, 10, 5) {real, imag} */,
  {32'h3e1f1f6a, 32'h00000000} /* (0, 10, 4) {real, imag} */,
  {32'h3c613e57, 32'h00000000} /* (0, 10, 3) {real, imag} */,
  {32'hbe8f8f54, 32'h00000000} /* (0, 10, 2) {real, imag} */,
  {32'hbe641331, 32'h00000000} /* (0, 10, 1) {real, imag} */,
  {32'hbd027368, 32'h00000000} /* (0, 10, 0) {real, imag} */,
  {32'hbe19b605, 32'h00000000} /* (0, 9, 31) {real, imag} */,
  {32'hbecb52aa, 32'h00000000} /* (0, 9, 30) {real, imag} */,
  {32'hbea66717, 32'h00000000} /* (0, 9, 29) {real, imag} */,
  {32'hbef6f9f3, 32'h00000000} /* (0, 9, 28) {real, imag} */,
  {32'hbf0c6678, 32'h00000000} /* (0, 9, 27) {real, imag} */,
  {32'hbed87c0a, 32'h00000000} /* (0, 9, 26) {real, imag} */,
  {32'hbe695b3a, 32'h00000000} /* (0, 9, 25) {real, imag} */,
  {32'hbe3ae216, 32'h00000000} /* (0, 9, 24) {real, imag} */,
  {32'hbed024ef, 32'h00000000} /* (0, 9, 23) {real, imag} */,
  {32'hbf32fcd2, 32'h00000000} /* (0, 9, 22) {real, imag} */,
  {32'hbf06b202, 32'h00000000} /* (0, 9, 21) {real, imag} */,
  {32'h3dacbc00, 32'h00000000} /* (0, 9, 20) {real, imag} */,
  {32'h3e978d93, 32'h00000000} /* (0, 9, 19) {real, imag} */,
  {32'h3e463ed4, 32'h00000000} /* (0, 9, 18) {real, imag} */,
  {32'h3e3db0a7, 32'h00000000} /* (0, 9, 17) {real, imag} */,
  {32'h3e83b018, 32'h00000000} /* (0, 9, 16) {real, imag} */,
  {32'h3e0a66d7, 32'h00000000} /* (0, 9, 15) {real, imag} */,
  {32'h3e8b5136, 32'h00000000} /* (0, 9, 14) {real, imag} */,
  {32'h3e21d7f2, 32'h00000000} /* (0, 9, 13) {real, imag} */,
  {32'h3f394aff, 32'h00000000} /* (0, 9, 12) {real, imag} */,
  {32'h3f3ce8dc, 32'h00000000} /* (0, 9, 11) {real, imag} */,
  {32'hbda24449, 32'h00000000} /* (0, 9, 10) {real, imag} */,
  {32'hbe8b6f87, 32'h00000000} /* (0, 9, 9) {real, imag} */,
  {32'hbe7afc87, 32'h00000000} /* (0, 9, 8) {real, imag} */,
  {32'hbf0da3b7, 32'h00000000} /* (0, 9, 7) {real, imag} */,
  {32'hbe586a3e, 32'h00000000} /* (0, 9, 6) {real, imag} */,
  {32'hbed374d1, 32'h00000000} /* (0, 9, 5) {real, imag} */,
  {32'hbdccb694, 32'h00000000} /* (0, 9, 4) {real, imag} */,
  {32'hbc627c4b, 32'h00000000} /* (0, 9, 3) {real, imag} */,
  {32'hbea5a171, 32'h00000000} /* (0, 9, 2) {real, imag} */,
  {32'hbed3421a, 32'h00000000} /* (0, 9, 1) {real, imag} */,
  {32'hbe8be06d, 32'h00000000} /* (0, 9, 0) {real, imag} */,
  {32'hbe1430e1, 32'h00000000} /* (0, 8, 31) {real, imag} */,
  {32'hbddcf502, 32'h00000000} /* (0, 8, 30) {real, imag} */,
  {32'hbe9edf1a, 32'h00000000} /* (0, 8, 29) {real, imag} */,
  {32'hbebcba06, 32'h00000000} /* (0, 8, 28) {real, imag} */,
  {32'hbe0a04eb, 32'h00000000} /* (0, 8, 27) {real, imag} */,
  {32'hbe86e251, 32'h00000000} /* (0, 8, 26) {real, imag} */,
  {32'hbe873c35, 32'h00000000} /* (0, 8, 25) {real, imag} */,
  {32'hbeadda11, 32'h00000000} /* (0, 8, 24) {real, imag} */,
  {32'hbf07972f, 32'h00000000} /* (0, 8, 23) {real, imag} */,
  {32'hbf206260, 32'h00000000} /* (0, 8, 22) {real, imag} */,
  {32'hbe27ee2f, 32'h00000000} /* (0, 8, 21) {real, imag} */,
  {32'h3e2ac2fd, 32'h00000000} /* (0, 8, 20) {real, imag} */,
  {32'h3e920fda, 32'h00000000} /* (0, 8, 19) {real, imag} */,
  {32'h3e1c459e, 32'h00000000} /* (0, 8, 18) {real, imag} */,
  {32'h3e3e9f81, 32'h00000000} /* (0, 8, 17) {real, imag} */,
  {32'h3ed01f29, 32'h00000000} /* (0, 8, 16) {real, imag} */,
  {32'h3f1bb16b, 32'h00000000} /* (0, 8, 15) {real, imag} */,
  {32'h3f25e6e9, 32'h00000000} /* (0, 8, 14) {real, imag} */,
  {32'h3eb402b7, 32'h00000000} /* (0, 8, 13) {real, imag} */,
  {32'h3f08d089, 32'h00000000} /* (0, 8, 12) {real, imag} */,
  {32'h3ed6647a, 32'h00000000} /* (0, 8, 11) {real, imag} */,
  {32'hbdae4804, 32'h00000000} /* (0, 8, 10) {real, imag} */,
  {32'hbcd819bc, 32'h00000000} /* (0, 8, 9) {real, imag} */,
  {32'h3d0ca767, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hbe0c9a72, 32'h00000000} /* (0, 8, 7) {real, imag} */,
  {32'hbe291c63, 32'h00000000} /* (0, 8, 6) {real, imag} */,
  {32'hbe82b3fb, 32'h00000000} /* (0, 8, 5) {real, imag} */,
  {32'hbe0741d5, 32'h00000000} /* (0, 8, 4) {real, imag} */,
  {32'hbd8a5963, 32'h00000000} /* (0, 8, 3) {real, imag} */,
  {32'hbf0a49e9, 32'h00000000} /* (0, 8, 2) {real, imag} */,
  {32'hbf074f4f, 32'h00000000} /* (0, 8, 1) {real, imag} */,
  {32'hbe55e940, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'hbe5576d2, 32'h00000000} /* (0, 7, 31) {real, imag} */,
  {32'hbe62dd7f, 32'h00000000} /* (0, 7, 30) {real, imag} */,
  {32'hbe5d45b3, 32'h00000000} /* (0, 7, 29) {real, imag} */,
  {32'hbed53938, 32'h00000000} /* (0, 7, 28) {real, imag} */,
  {32'hbe754d43, 32'h00000000} /* (0, 7, 27) {real, imag} */,
  {32'hbeeda699, 32'h00000000} /* (0, 7, 26) {real, imag} */,
  {32'hbee67503, 32'h00000000} /* (0, 7, 25) {real, imag} */,
  {32'hbeea9122, 32'h00000000} /* (0, 7, 24) {real, imag} */,
  {32'hbed647b1, 32'h00000000} /* (0, 7, 23) {real, imag} */,
  {32'hbe6c9e40, 32'h00000000} /* (0, 7, 22) {real, imag} */,
  {32'h3d2481f2, 32'h00000000} /* (0, 7, 21) {real, imag} */,
  {32'h3ee43bd4, 32'h00000000} /* (0, 7, 20) {real, imag} */,
  {32'h3f03de9e, 32'h00000000} /* (0, 7, 19) {real, imag} */,
  {32'h3e9e271c, 32'h00000000} /* (0, 7, 18) {real, imag} */,
  {32'h3e9c0cd7, 32'h00000000} /* (0, 7, 17) {real, imag} */,
  {32'h3e990851, 32'h00000000} /* (0, 7, 16) {real, imag} */,
  {32'h3f20e6c7, 32'h00000000} /* (0, 7, 15) {real, imag} */,
  {32'h3f81f512, 32'h00000000} /* (0, 7, 14) {real, imag} */,
  {32'h3f21faa9, 32'h00000000} /* (0, 7, 13) {real, imag} */,
  {32'h3ef9f3cf, 32'h00000000} /* (0, 7, 12) {real, imag} */,
  {32'hbd81bbaf, 32'h00000000} /* (0, 7, 11) {real, imag} */,
  {32'hbebedecc, 32'h00000000} /* (0, 7, 10) {real, imag} */,
  {32'hbe4e889c, 32'h00000000} /* (0, 7, 9) {real, imag} */,
  {32'hbc76dae9, 32'h00000000} /* (0, 7, 8) {real, imag} */,
  {32'hbda9ff64, 32'h00000000} /* (0, 7, 7) {real, imag} */,
  {32'hbf1768b6, 32'h00000000} /* (0, 7, 6) {real, imag} */,
  {32'hbf14189c, 32'h00000000} /* (0, 7, 5) {real, imag} */,
  {32'hbea5b53e, 32'h00000000} /* (0, 7, 4) {real, imag} */,
  {32'hbe1c81b1, 32'h00000000} /* (0, 7, 3) {real, imag} */,
  {32'hbf44cb5b, 32'h00000000} /* (0, 7, 2) {real, imag} */,
  {32'hbf2e434c, 32'h00000000} /* (0, 7, 1) {real, imag} */,
  {32'hbd7f2180, 32'h00000000} /* (0, 7, 0) {real, imag} */,
  {32'hbdb7c614, 32'h00000000} /* (0, 6, 31) {real, imag} */,
  {32'hbdeb3a89, 32'h00000000} /* (0, 6, 30) {real, imag} */,
  {32'hbe8da89b, 32'h00000000} /* (0, 6, 29) {real, imag} */,
  {32'hbf1e3dd5, 32'h00000000} /* (0, 6, 28) {real, imag} */,
  {32'hbedb8fb0, 32'h00000000} /* (0, 6, 27) {real, imag} */,
  {32'hbf17f480, 32'h00000000} /* (0, 6, 26) {real, imag} */,
  {32'hbf10bc67, 32'h00000000} /* (0, 6, 25) {real, imag} */,
  {32'hbf2a6d46, 32'h00000000} /* (0, 6, 24) {real, imag} */,
  {32'hbea7e1f9, 32'h00000000} /* (0, 6, 23) {real, imag} */,
  {32'hbefe0cd6, 32'h00000000} /* (0, 6, 22) {real, imag} */,
  {32'hbe551fd1, 32'h00000000} /* (0, 6, 21) {real, imag} */,
  {32'h3f4941aa, 32'h00000000} /* (0, 6, 20) {real, imag} */,
  {32'h3f09014d, 32'h00000000} /* (0, 6, 19) {real, imag} */,
  {32'h3eb0b45d, 32'h00000000} /* (0, 6, 18) {real, imag} */,
  {32'h3e761ac6, 32'h00000000} /* (0, 6, 17) {real, imag} */,
  {32'h3e6d3d25, 32'h00000000} /* (0, 6, 16) {real, imag} */,
  {32'h3ef63060, 32'h00000000} /* (0, 6, 15) {real, imag} */,
  {32'h3f3068ed, 32'h00000000} /* (0, 6, 14) {real, imag} */,
  {32'h3e6058b1, 32'h00000000} /* (0, 6, 13) {real, imag} */,
  {32'h3eac45b5, 32'h00000000} /* (0, 6, 12) {real, imag} */,
  {32'h3df7cd8d, 32'h00000000} /* (0, 6, 11) {real, imag} */,
  {32'hbe49af0d, 32'h00000000} /* (0, 6, 10) {real, imag} */,
  {32'hbf371308, 32'h00000000} /* (0, 6, 9) {real, imag} */,
  {32'hbf0fbfc9, 32'h00000000} /* (0, 6, 8) {real, imag} */,
  {32'hbe820199, 32'h00000000} /* (0, 6, 7) {real, imag} */,
  {32'hbf092dd1, 32'h00000000} /* (0, 6, 6) {real, imag} */,
  {32'hbf029f58, 32'h00000000} /* (0, 6, 5) {real, imag} */,
  {32'hbe784ed9, 32'h00000000} /* (0, 6, 4) {real, imag} */,
  {32'hbcf98c27, 32'h00000000} /* (0, 6, 3) {real, imag} */,
  {32'hbe34476f, 32'h00000000} /* (0, 6, 2) {real, imag} */,
  {32'h3c220e07, 32'h00000000} /* (0, 6, 1) {real, imag} */,
  {32'h3d049355, 32'h00000000} /* (0, 6, 0) {real, imag} */,
  {32'hbec758d0, 32'h00000000} /* (0, 5, 31) {real, imag} */,
  {32'hbf19e679, 32'h00000000} /* (0, 5, 30) {real, imag} */,
  {32'hbf19d066, 32'h00000000} /* (0, 5, 29) {real, imag} */,
  {32'hbf7ecb8b, 32'h00000000} /* (0, 5, 28) {real, imag} */,
  {32'hbf5cc603, 32'h00000000} /* (0, 5, 27) {real, imag} */,
  {32'hbebdc19d, 32'h00000000} /* (0, 5, 26) {real, imag} */,
  {32'hbea1fdd9, 32'h00000000} /* (0, 5, 25) {real, imag} */,
  {32'hbf1ca674, 32'h00000000} /* (0, 5, 24) {real, imag} */,
  {32'hbf2e7465, 32'h00000000} /* (0, 5, 23) {real, imag} */,
  {32'hbf26da76, 32'h00000000} /* (0, 5, 22) {real, imag} */,
  {32'hbeb1f957, 32'h00000000} /* (0, 5, 21) {real, imag} */,
  {32'hbdbd05e0, 32'h00000000} /* (0, 5, 20) {real, imag} */,
  {32'hbd93a79a, 32'h00000000} /* (0, 5, 19) {real, imag} */,
  {32'hbd255e46, 32'h00000000} /* (0, 5, 18) {real, imag} */,
  {32'hbf22f0d5, 32'h00000000} /* (0, 5, 17) {real, imag} */,
  {32'hbef4a218, 32'h00000000} /* (0, 5, 16) {real, imag} */,
  {32'hbdd2b574, 32'h00000000} /* (0, 5, 15) {real, imag} */,
  {32'h3e68d349, 32'h00000000} /* (0, 5, 14) {real, imag} */,
  {32'hbc5c6f86, 32'h00000000} /* (0, 5, 13) {real, imag} */,
  {32'h3dc8436f, 32'h00000000} /* (0, 5, 12) {real, imag} */,
  {32'h3df0d27e, 32'h00000000} /* (0, 5, 11) {real, imag} */,
  {32'h3c1e566e, 32'h00000000} /* (0, 5, 10) {real, imag} */,
  {32'hbca3cdda, 32'h00000000} /* (0, 5, 9) {real, imag} */,
  {32'h392c1b80, 32'h00000000} /* (0, 5, 8) {real, imag} */,
  {32'hbde7f0bd, 32'h00000000} /* (0, 5, 7) {real, imag} */,
  {32'hbebc879a, 32'h00000000} /* (0, 5, 6) {real, imag} */,
  {32'hbe5a26d4, 32'h00000000} /* (0, 5, 5) {real, imag} */,
  {32'hbe124d5f, 32'h00000000} /* (0, 5, 4) {real, imag} */,
  {32'hbe6222c7, 32'h00000000} /* (0, 5, 3) {real, imag} */,
  {32'hbeaf258a, 32'h00000000} /* (0, 5, 2) {real, imag} */,
  {32'hbecd3685, 32'h00000000} /* (0, 5, 1) {real, imag} */,
  {32'hbe0dec4b, 32'h00000000} /* (0, 5, 0) {real, imag} */,
  {32'hbedc825f, 32'h00000000} /* (0, 4, 31) {real, imag} */,
  {32'hbf108ba2, 32'h00000000} /* (0, 4, 30) {real, imag} */,
  {32'hbf313c96, 32'h00000000} /* (0, 4, 29) {real, imag} */,
  {32'hbf8aa427, 32'h00000000} /* (0, 4, 28) {real, imag} */,
  {32'hbf33810e, 32'h00000000} /* (0, 4, 27) {real, imag} */,
  {32'hbeb21f26, 32'h00000000} /* (0, 4, 26) {real, imag} */,
  {32'hbeb691d2, 32'h00000000} /* (0, 4, 25) {real, imag} */,
  {32'hbf307aea, 32'h00000000} /* (0, 4, 24) {real, imag} */,
  {32'hbf17262f, 32'h00000000} /* (0, 4, 23) {real, imag} */,
  {32'hbeef7462, 32'h00000000} /* (0, 4, 22) {real, imag} */,
  {32'hbe609e50, 32'h00000000} /* (0, 4, 21) {real, imag} */,
  {32'hbf0debc0, 32'h00000000} /* (0, 4, 20) {real, imag} */,
  {32'hbf42e395, 32'h00000000} /* (0, 4, 19) {real, imag} */,
  {32'hbea85820, 32'h00000000} /* (0, 4, 18) {real, imag} */,
  {32'hbf1a973a, 32'h00000000} /* (0, 4, 17) {real, imag} */,
  {32'hbf1b133a, 32'h00000000} /* (0, 4, 16) {real, imag} */,
  {32'h3e6e3891, 32'h00000000} /* (0, 4, 15) {real, imag} */,
  {32'h3f3757a7, 32'h00000000} /* (0, 4, 14) {real, imag} */,
  {32'h3e367c85, 32'h00000000} /* (0, 4, 13) {real, imag} */,
  {32'h3d882947, 32'h00000000} /* (0, 4, 12) {real, imag} */,
  {32'h3e1208db, 32'h00000000} /* (0, 4, 11) {real, imag} */,
  {32'h3e270650, 32'h00000000} /* (0, 4, 10) {real, imag} */,
  {32'h3f00275b, 32'h00000000} /* (0, 4, 9) {real, imag} */,
  {32'h3eac2bdf, 32'h00000000} /* (0, 4, 8) {real, imag} */,
  {32'h3ed4f50e, 32'h00000000} /* (0, 4, 7) {real, imag} */,
  {32'h3e4d2a29, 32'h00000000} /* (0, 4, 6) {real, imag} */,
  {32'hbe34b9c7, 32'h00000000} /* (0, 4, 5) {real, imag} */,
  {32'hbe5f965b, 32'h00000000} /* (0, 4, 4) {real, imag} */,
  {32'hbed4c45a, 32'h00000000} /* (0, 4, 3) {real, imag} */,
  {32'hbf03d9a3, 32'h00000000} /* (0, 4, 2) {real, imag} */,
  {32'hbf0e4d59, 32'h00000000} /* (0, 4, 1) {real, imag} */,
  {32'hbe10e82b, 32'h00000000} /* (0, 4, 0) {real, imag} */,
  {32'hbe5cc56b, 32'h00000000} /* (0, 3, 31) {real, imag} */,
  {32'hbe65d5e9, 32'h00000000} /* (0, 3, 30) {real, imag} */,
  {32'hbe4298d5, 32'h00000000} /* (0, 3, 29) {real, imag} */,
  {32'hbed6a706, 32'h00000000} /* (0, 3, 28) {real, imag} */,
  {32'hbec220c1, 32'h00000000} /* (0, 3, 27) {real, imag} */,
  {32'hbec0db8b, 32'h00000000} /* (0, 3, 26) {real, imag} */,
  {32'hbf30e50b, 32'h00000000} /* (0, 3, 25) {real, imag} */,
  {32'hbf768c44, 32'h00000000} /* (0, 3, 24) {real, imag} */,
  {32'hbf399e05, 32'h00000000} /* (0, 3, 23) {real, imag} */,
  {32'hbf157f7a, 32'h00000000} /* (0, 3, 22) {real, imag} */,
  {32'hbe986cc6, 32'h00000000} /* (0, 3, 21) {real, imag} */,
  {32'hbec5f0bf, 32'h00000000} /* (0, 3, 20) {real, imag} */,
  {32'hbf43b1f4, 32'h00000000} /* (0, 3, 19) {real, imag} */,
  {32'hbf7e62a7, 32'h00000000} /* (0, 3, 18) {real, imag} */,
  {32'hbf27daba, 32'h00000000} /* (0, 3, 17) {real, imag} */,
  {32'hbeb5d84b, 32'h00000000} /* (0, 3, 16) {real, imag} */,
  {32'h3e4bc44b, 32'h00000000} /* (0, 3, 15) {real, imag} */,
  {32'h3f0a9671, 32'h00000000} /* (0, 3, 14) {real, imag} */,
  {32'h3ed99913, 32'h00000000} /* (0, 3, 13) {real, imag} */,
  {32'h3ee075e9, 32'h00000000} /* (0, 3, 12) {real, imag} */,
  {32'h3ee5a10e, 32'h00000000} /* (0, 3, 11) {real, imag} */,
  {32'h3e40a352, 32'h00000000} /* (0, 3, 10) {real, imag} */,
  {32'h3dae23b3, 32'h00000000} /* (0, 3, 9) {real, imag} */,
  {32'h3dd0a2a9, 32'h00000000} /* (0, 3, 8) {real, imag} */,
  {32'h3e6b88c0, 32'h00000000} /* (0, 3, 7) {real, imag} */,
  {32'h3e1c5619, 32'h00000000} /* (0, 3, 6) {real, imag} */,
  {32'hbe55ae31, 32'h00000000} /* (0, 3, 5) {real, imag} */,
  {32'hbe7c7208, 32'h00000000} /* (0, 3, 4) {real, imag} */,
  {32'hbea5886b, 32'h00000000} /* (0, 3, 3) {real, imag} */,
  {32'hbe8d2076, 32'h00000000} /* (0, 3, 2) {real, imag} */,
  {32'hbe636093, 32'h00000000} /* (0, 3, 1) {real, imag} */,
  {32'hbd954eba, 32'h00000000} /* (0, 3, 0) {real, imag} */,
  {32'hbeaf17c7, 32'h00000000} /* (0, 2, 31) {real, imag} */,
  {32'hbe802cb1, 32'h00000000} /* (0, 2, 30) {real, imag} */,
  {32'hbe0099af, 32'h00000000} /* (0, 2, 29) {real, imag} */,
  {32'hbe9a2581, 32'h00000000} /* (0, 2, 28) {real, imag} */,
  {32'hbed6ac2e, 32'h00000000} /* (0, 2, 27) {real, imag} */,
  {32'hbede942d, 32'h00000000} /* (0, 2, 26) {real, imag} */,
  {32'hbf08b933, 32'h00000000} /* (0, 2, 25) {real, imag} */,
  {32'hbea84618, 32'h00000000} /* (0, 2, 24) {real, imag} */,
  {32'hbec6530a, 32'h00000000} /* (0, 2, 23) {real, imag} */,
  {32'hbee5657a, 32'h00000000} /* (0, 2, 22) {real, imag} */,
  {32'h3c0e3280, 32'h00000000} /* (0, 2, 21) {real, imag} */,
  {32'h3dba7928, 32'h00000000} /* (0, 2, 20) {real, imag} */,
  {32'hbe93488e, 32'h00000000} /* (0, 2, 19) {real, imag} */,
  {32'hbf532a6d, 32'h00000000} /* (0, 2, 18) {real, imag} */,
  {32'hbf2ad166, 32'h00000000} /* (0, 2, 17) {real, imag} */,
  {32'hbed62457, 32'h00000000} /* (0, 2, 16) {real, imag} */,
  {32'hbbb3fd68, 32'h00000000} /* (0, 2, 15) {real, imag} */,
  {32'h3ec3f0b7, 32'h00000000} /* (0, 2, 14) {real, imag} */,
  {32'h3f20305d, 32'h00000000} /* (0, 2, 13) {real, imag} */,
  {32'h3ef1c71c, 32'h00000000} /* (0, 2, 12) {real, imag} */,
  {32'h3f5c99fe, 32'h00000000} /* (0, 2, 11) {real, imag} */,
  {32'h3f178f38, 32'h00000000} /* (0, 2, 10) {real, imag} */,
  {32'h3e8989f3, 32'h00000000} /* (0, 2, 9) {real, imag} */,
  {32'h3e967bab, 32'h00000000} /* (0, 2, 8) {real, imag} */,
  {32'h3e580c32, 32'h00000000} /* (0, 2, 7) {real, imag} */,
  {32'h3ee58361, 32'h00000000} /* (0, 2, 6) {real, imag} */,
  {32'hbe0aeaad, 32'h00000000} /* (0, 2, 5) {real, imag} */,
  {32'hbedf88ec, 32'h00000000} /* (0, 2, 4) {real, imag} */,
  {32'hbe4ab141, 32'h00000000} /* (0, 2, 3) {real, imag} */,
  {32'hbdcb684f, 32'h00000000} /* (0, 2, 2) {real, imag} */,
  {32'hbe40fe08, 32'h00000000} /* (0, 2, 1) {real, imag} */,
  {32'hbe9d2a34, 32'h00000000} /* (0, 2, 0) {real, imag} */,
  {32'hbe54e78d, 32'h00000000} /* (0, 1, 31) {real, imag} */,
  {32'hbeac3a8e, 32'h00000000} /* (0, 1, 30) {real, imag} */,
  {32'hbec575b3, 32'h00000000} /* (0, 1, 29) {real, imag} */,
  {32'hbe900032, 32'h00000000} /* (0, 1, 28) {real, imag} */,
  {32'hbe98c323, 32'h00000000} /* (0, 1, 27) {real, imag} */,
  {32'hbec43cb8, 32'h00000000} /* (0, 1, 26) {real, imag} */,
  {32'hbea0689a, 32'h00000000} /* (0, 1, 25) {real, imag} */,
  {32'hb8e55280, 32'h00000000} /* (0, 1, 24) {real, imag} */,
  {32'hbe4c23ae, 32'h00000000} /* (0, 1, 23) {real, imag} */,
  {32'hbea6ceca, 32'h00000000} /* (0, 1, 22) {real, imag} */,
  {32'hbd943cf8, 32'h00000000} /* (0, 1, 21) {real, imag} */,
  {32'h3d87c7c8, 32'h00000000} /* (0, 1, 20) {real, imag} */,
  {32'hbe315819, 32'h00000000} /* (0, 1, 19) {real, imag} */,
  {32'hbf14c9ea, 32'h00000000} /* (0, 1, 18) {real, imag} */,
  {32'hbf042972, 32'h00000000} /* (0, 1, 17) {real, imag} */,
  {32'hbf08849b, 32'h00000000} /* (0, 1, 16) {real, imag} */,
  {32'h3da70c6d, 32'h00000000} /* (0, 1, 15) {real, imag} */,
  {32'h3efcf8d6, 32'h00000000} /* (0, 1, 14) {real, imag} */,
  {32'h3f0e75d7, 32'h00000000} /* (0, 1, 13) {real, imag} */,
  {32'h3f1572fd, 32'h00000000} /* (0, 1, 12) {real, imag} */,
  {32'h3f68a8f8, 32'h00000000} /* (0, 1, 11) {real, imag} */,
  {32'h3ee60ced, 32'h00000000} /* (0, 1, 10) {real, imag} */,
  {32'h3f088d73, 32'h00000000} /* (0, 1, 9) {real, imag} */,
  {32'h3f769bc8, 32'h00000000} /* (0, 1, 8) {real, imag} */,
  {32'h3f764aaa, 32'h00000000} /* (0, 1, 7) {real, imag} */,
  {32'h3f5ec90c, 32'h00000000} /* (0, 1, 6) {real, imag} */,
  {32'hbe2c27dc, 32'h00000000} /* (0, 1, 5) {real, imag} */,
  {32'hbf129fa8, 32'h00000000} /* (0, 1, 4) {real, imag} */,
  {32'hbf0ac8b1, 32'h00000000} /* (0, 1, 3) {real, imag} */,
  {32'hbe85c3c6, 32'h00000000} /* (0, 1, 2) {real, imag} */,
  {32'hbdd756cd, 32'h00000000} /* (0, 1, 1) {real, imag} */,
  {32'hbe139f86, 32'h00000000} /* (0, 1, 0) {real, imag} */,
  {32'hbe53a89c, 32'h00000000} /* (0, 0, 31) {real, imag} */,
  {32'hbec76961, 32'h00000000} /* (0, 0, 30) {real, imag} */,
  {32'hbf27731a, 32'h00000000} /* (0, 0, 29) {real, imag} */,
  {32'hbec109cf, 32'h00000000} /* (0, 0, 28) {real, imag} */,
  {32'hbeb5e633, 32'h00000000} /* (0, 0, 27) {real, imag} */,
  {32'hbeb50601, 32'h00000000} /* (0, 0, 26) {real, imag} */,
  {32'hbcb83de8, 32'h00000000} /* (0, 0, 25) {real, imag} */,
  {32'h3d530409, 32'h00000000} /* (0, 0, 24) {real, imag} */,
  {32'hbe4e608d, 32'h00000000} /* (0, 0, 23) {real, imag} */,
  {32'hbe5dd8b9, 32'h00000000} /* (0, 0, 22) {real, imag} */,
  {32'hbdc19b0e, 32'h00000000} /* (0, 0, 21) {real, imag} */,
  {32'hbd3609c5, 32'h00000000} /* (0, 0, 20) {real, imag} */,
  {32'hbde4db85, 32'h00000000} /* (0, 0, 19) {real, imag} */,
  {32'hbe2db9dc, 32'h00000000} /* (0, 0, 18) {real, imag} */,
  {32'hbe275cba, 32'h00000000} /* (0, 0, 17) {real, imag} */,
  {32'hbec473ab, 32'h00000000} /* (0, 0, 16) {real, imag} */,
  {32'h3e0cc667, 32'h00000000} /* (0, 0, 15) {real, imag} */,
  {32'h3effcb1f, 32'h00000000} /* (0, 0, 14) {real, imag} */,
  {32'h3e91eaf8, 32'h00000000} /* (0, 0, 13) {real, imag} */,
  {32'h3e7cf596, 32'h00000000} /* (0, 0, 12) {real, imag} */,
  {32'h3ec280f5, 32'h00000000} /* (0, 0, 11) {real, imag} */,
  {32'h3e09426e, 32'h00000000} /* (0, 0, 10) {real, imag} */,
  {32'h3e1f5424, 32'h00000000} /* (0, 0, 9) {real, imag} */,
  {32'h3efe988f, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h3f0cb0c1, 32'h00000000} /* (0, 0, 7) {real, imag} */,
  {32'h3ef7bbfb, 32'h00000000} /* (0, 0, 6) {real, imag} */,
  {32'h3dbdc04d, 32'h00000000} /* (0, 0, 5) {real, imag} */,
  {32'hbe1ad2ad, 32'h00000000} /* (0, 0, 4) {real, imag} */,
  {32'hbe97e14b, 32'h00000000} /* (0, 0, 3) {real, imag} */,
  {32'hbe954d3d, 32'h00000000} /* (0, 0, 2) {real, imag} */,
  {32'hbd766893, 32'h00000000} /* (0, 0, 1) {real, imag} */,
  {32'hbd112ca7, 32'h00000000} /* (0, 0, 0) {real, imag} */};
