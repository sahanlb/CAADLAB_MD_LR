-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ukZaEuyLkuKdQRqz/gttc1kOym3xvV+JFSIf2Hna5i1Hcgy3eq6x/rC0It5cBJa28pPkx12i7DL4
/T414pUFRHYaJbGwq0XYHmUTbPZ1WqCiS04wrxZPjMcDa1Pgk02cBZnB9IoRzQc0ji9NXwNEnwd7
xR9ejnUYHXzG4hdOIQXywplF7AV4MtF7j6AwrS5aPt3NvjxM/T8dv4IOh88Yi8irBF2oqkT/vS8H
wzoveiFMatz0cMctVWC2rGp8J+OSdGKQlEwb17n2GcE+70eC9KeSH2YjGoHmDsqQUU1OFDTvpEym
KJAqTUEoR6XotjRuPYYEqaZvyCconGAavsbOjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11536)
`protect data_block
z3kUqlsqcjF0bAXIhSvh/X0pgsevYfJsehXRlZft7JPxpCmPoyjQO/Q+qkylpk5VF2MpmeRh0awX
hVVdiKhtksU/T4h8483Gi66bbhmXq3Tqg2sgUb1dLnFI8btigTD6wGdJVnKg9ry3Qo96UjGrtUeZ
HtHdtG78o643zbDGR8bzCaTpidpnC5dBoy7jzag6C1gUA9LCdXJx3YTNhAupq1ovC7biycPFSNyO
vzteIvFzdwEHwwKNtJ3PGN38aqd+dKFjn82zGGC/LcEYCgLsDprMoLxSxkE2sLxXLCJsNz6JCFGq
8bYMVWcLnpstPfQcU2aVapNfy1bwRNuNbAMbJFIh8jBkexgUgPw0Jh/EsJN9NI+Tbhs/4I6VC519
9Nl2Q2WRAWgzeP1CDFP7zonHphIqusk5g/TgJEC5gODwQTrWmbnNlzmxtall9BGbExUyBT33MZoh
jv9DobpIlz0lbgkzCgIFDe+Z8AE+LWOJL+VaVtgwXnjiJasxMYT7wv9lHOAHpFfio1zkGn705Lb6
XbFBSB0kSbqJFgBnYZOVo7MoJrVDjSPq3QHkrFWu095q08l7OfbhZmqfJZ90n5tLe1jbvjNwppkI
nOf4+3+W3QlolSBNvy7o7JI0S2bi4WWKVlnIjVf7BXZ+XCbz4B5OzjQr/dJc4q/k+LBnbnBTqVpE
ycaHd8/nWX9FYn3gt8Kvn4GczQ8TPg7ILR5tN3VN29EJobMZP1u7RKAQ8mVItmghblM1Yjg1h0ne
hjDrtiif8IkaBDeLEV1yRHbQyFmPAIC+Z7I4Malbmn1174egibrl6nWouf9x9LvzlxDGG92bteG7
bpeDIx7VGI5DhD5RjoKdE6cOWuFbHSWqdCWio2szhOwQweA0oLJxp4IFyQDRgPI29D9OWO/9gXSL
1W32c6RFaV9gk/rgX5k2EwSmtt5HLfSG4en/uL/aIJkVI/dONCW363UqQoymBLRkW2/OVzXk3w56
cdd0yPUsIZXh4NR9exAVxoCspJpZY+JVgMFLOutDYWANCU8EXl5h5EwhV3mBDd+Cx3Bcqg82c1to
DyBcJQRHc3zBAs2v0VmW9BOhbXiBv3XIRnH5/3d0LhgOvSPWJdbM5yvB/xWgLZF1m1CXbgoi8XYr
kt59aiVdMK8ykobmY772hqRNQxv4lcScvQJzKfRf2mQuMlSPPyoa+s31cb1etvgcYnuJgEvrZm04
uGN6lvUw7+xBxfbS4eXUxJncgm8ZcF+4PhSHzwVp59yB84g5igfZP6qgLQSM5mRbMAfCtxFcBBDB
/3pRscGwh3fStHPwXl72y++6jyt1refWFwHBCMOu5EfPlP09I2JfSsQAmau6UrQT1wyA5LRSMuhf
FKvoWcP/vOsiC7gmab8ovYMqulnxaTqcCoE+3+zCWShu+HiU5vHDOx9k1gHcR3PMLnDjYcUc0mUk
GxauFqktNjfZD/9w9r49Q9ZfztODu/4zzPwNSyWgWfWENMVUjVvHtNTMX5mUNCW/wF9wcCy3JEQV
3FIFwokk28PRXpsfOzNwBqNhUK/yezfhVbSJYXL4fQRkURMUdELtMpjQXn1CVjfZHm+RvkKd4mBU
FrcnY4C+1kokEzq5hPclx5LwGLvbFezgU94H4sDLvgFZ3bdIstMwigmYGEJHfhBvVBdBobQ9F9ap
v9hm6OVtGlO7L4AGHSLy9hRUqIv6ZfZCUuMsTfP3Seb0DqzDUxnifNWRgFfULycL9CcLDgFKujxc
WfiTiV9wPkftE8OmGfQq2W/DGlh5FuNywXRDjUMxFtijextVQmi8KMe9dygRtXCJu01jUz3Ey76+
s1cWWRnPX6xz5XawUMYR15NJqQMSzdLQP82SB3fmbXM7XKLkm5aU6jwhn20x7TXJ6gGZLM8G8Y1+
rbFuHrAcqjYDau4AoqvEf5BRwUszj1A2ie8NCRm+cXUq9O3+nAhcqAMjRvsIwInLW4HDXfhdEFo9
QyW+XOigO7q+4O5SunA+weS1sxfEbf/HBVO1xv0hs78iI0tiX44Nd57bczdV1q149VE0tB1r5z6K
x6Et8uZYzwsndByUhAA/hw4NaNRkfiJBdWCUPwq226cNWqX18hoMjvDyP5qNUl6dWTggxz0Yn6/P
/dVEWIj4RcjNdqoAT/rQOAVH9mPmyiJUkR4UuMVkUpY/geQ35IF+6BL16F5d989Q0DkS8bGyuFXq
6Ogy43hqCgp1uuP3tECFOe9xZrc8JGc9VshuPvku4JXbtZ3u6me1S2vomEKG3ODeNVTeX3bR68+N
4ps/fHAO4N2sXx9jPO0Yi9OWvR4t+u2ZD78ym+m3B42wKYuQAwqkAffGyYyQxfACVXTiUEkEoLXP
oLg3klisx5T8FvweRD9E6w+WfeiA5WGCF9tH7E7AtQevankr+CU7N/SxI/l/KWHkCys+dtmm2AM6
PDQfhdYpWtxcRCRu1OoR4ddPlT2UWUc87SnpKyWqPhPx9aGKaqPi0S05CIRD1YIFvhNEuRGZDfP/
EYey6I+DTB5jlO+5kXT2T4ILCBJzg8kLPriI6K52t02nVr/mxxhU1TMPpkEz9L487QsMMm6MyHn4
FMV5O3Upgbhxtd7uCYKlicgsnwcv8L5sdToneQiocYQcZsnZ3A2xHwAgs4WktbaWaHhc5Zku71Fz
GOB/z3KZ39dY/Lc+2F7h1pI+/Zj/p9TUB+UTGbL33BfRELZCkAhbr/L3+z+BM6zZTstEKr1QS7Ru
aEXWgPQ3rmbpbyDctppZbQfkriDmfyohle0RsGE5LSSUsQ3+ycS1h3/mBo885nlFRovlr9MkQLgx
nDBtDtCfKzkVu8a8oh3D6avcntqNKW7QstTheY0AoEVzrFtxi8qT/tBgX7FxmFksMwiX4iLkhRO2
NqrH1zdceN9/aA5tFAU5dDQA+hPJPuGxpwjkXm/wV1pbRCXO51mObSJViQpDCEbBcxdOoK6/pf9o
/9uMguXDWZlmvjp2dYjD6ymvVKjI3tEoYDWuJUS/6XRghrFakv9ay/+BqqlV9jKQ2qEU55TEh10Z
V20wF5raUSK8pi2jxHJBMbhGLP5USLTDWhiM2VW6zGYXZXukkvCUPDXqFEemsC5wi8/x3bnLsFD0
4DDO3/El3/CI3BQVbY/F6vZjiGC2lCJfVK/+VWM0QPnilsx3JYngsSxT+MTtjXQXQ44NCe3hJXoX
uPFPAdzMLkTaTpiQuNy4auRbgl1k8I5XGrLJky1Uta4z9CFygMH2GSogjdsv7kgWPITXiPx2RDD5
nkuTx6PTBDftR2botjvtalRF3bv+NkAgINqAYq9e6i+KQ5YFxVeG6UqFhtj/GCDiPBZ8O9uX3UXj
47IovrHjqKvkhKjIvvYX62KYG2bceWDiiGtffYkYioTwxzs2ewSlVHwBUPCpGb8TO+K14xRzE59D
OUjnxItIkknqOKkV/IjNUs17Xwn0d9oZl8LIsVcBRSI3q2RcW+5BKqJNElO4F1WkI8AIOomfI6zG
HU8TC3an6mJq7hsu6r31uG7FIiOaGYXcXtKaAPG3bDsxwkOW8+XWku800H6116hVhhzrWyxBat2w
agGFn9OX3kyG/JEHEGudNDBAHUK6XpyJoqjn/DURtBf+u0ibNxtAfTkeJsdFNAIK9SSJw0GnK0u2
9vaynSsdU53cpqbT3EPoXKREEPrhK93GruI7UYDIZBM4nyERRlBhZlWLNlweaeqbjm7PabUVcTM7
DYm1c0NQlYYYRrhBtsJU5/zUmgpGMYWjxH8KHvnWOoxx+D1ETUL15C8QDF8VFQEop7kAKjYgIbtJ
jh/xDgxXEKb3/dfX8rlOuS6vdscVi5As4E5eHDELUE17BwE8MwP3x0AxTNwlYhaeDSaed8h+L2GD
TlfOQVZHo+61j5AOXsnPJI3R1kVQv24iBpDBeOopTR/JRnqtNuAne7sftlaeYQBFigc1sAggM2Z0
9hNpHpQT+qr2n38Ot4TC2CBUgDTlVQOS36JzloAimyE0jJTYdWAfG7XbUMzlNnccWhXn2gl11Bde
vkD7oPHnUoaei5pWReYK/BKypgJgiCkjcLPO3qj9NFULSgeVQAdCtcct7gU9StP+YfkxbzfyiPSg
IOcTqyZFScngRBKqwkInmUScwsxsU1lEH/1vBIBv4OS5FsTwGKy4zdwDPwT7ZkH/mEX8hGevMD7e
e7OhAjPe6jnjxC5f57FY1F93Nf3expvJAqwLvsz3+I4MEtu8KSKbn63ydR9K0zo3A7IIyVVCeuSK
HeR1BnGGRYxWYmgGMjCG/BX1j3Ves7oJVcSR8zYNNAoqghNFvMcb45yQccJPI/OcAvD8gzt+HITb
PxeOl+CXFnkh9WUtUUhBvVRdeG7yUoLyJrQgf8k3IkdGJuk2vLdjDikpmlHRNj959oLO1HSDe7XY
9frhEsgpOl9fA2EJG7TgATQEXx7jx370xALSF0usRQbjxIIA9rJGjNicaOEKqwf6RZ8Yi8eJJDMw
j14z4LG8HgDC1E90YJOKFeHhIvyC/pV18vk6+y58scrCU9XxExA/oIm13MbX436gC2czXtT3BzC+
mVAvLz4U51kL1SA2Gy3xHIAJ/uQLbO+mbnC5ClKzV6qlKOdZDsvkP0jV9W9stPR40R4/6aESodkc
9jvunJOHY0dlPG7YbhB1IqpyydLSNGvQ1PaVtH5qZZbzt/uIYC0hdZwKIHzby5Dfq2fWhkSUIbEu
SOC+4x3HyQpABgvf33QPmZMkq8h0vb0jbW2bLq/3+eaOxwHpcLi/j8t7PL9LUGdteBVuyCDe43j9
yha6bOzR2bXgK2DGvN0SH4DlmCofKQFRxl8a/A5UCCNfszy7Qd5Z2u6BhRZmM+uYolFesR0PrH49
dCES5aKgNo+LFaZEsbCafCdejIJhiCdoCmAmh0Jt5dUrb37jXZtcYg1LpyxI+T8A4+vdfTH1tp/A
PwkDzXRtc/nVywRcB7VT5+n90zHXDNWhRbhc1aJxW2KzuKBiit63weOJnc91WT63JxJJ50xX4qZN
IFIgz8nnWXJyRNXkIET9AuyX+vqTb2qHHE0aane5iTv5VUuhLPot1FCrml3a0mddCjE+LabCL8ty
eTUm1bOVL6uBrkU0VVZvJsM1o+PF3pkIhuNOBZaFqbV69tGpqCa9I49w1IbI796hR2/huECS1sIY
2vWEwmqpequROo0X6y9vbe4CBFH6BwY0bBXJEmemPk5XSGc9BuCjgeOgumHae4M30G1k0fUZcVbr
lsbm8ebzxTwppKwquWZgeCS6i/wmdD6ib7gv/ivM5Kdx4m++QAE/xJ8AAw9sMuy2gSH+2GrbS/JJ
2tXyRAmxVeXBVqv2gtMzhgwvVa8MmpRlUfuD9CYtauzmuh3vk/E4CmTiDjvb+dQqwm+yBs9Y2hQi
4Xxp29C33x3kVRNT79146HfnU82RSRF95UeYAuemMVUHqmwLNSyaMhq4BSIWoXcWoohAL5/0IL3G
elmEZlvff+DHwRbondEts2785KqS0a3KXlOVKhxtQgQFOVf98iF7AcX4gKhzPgjGPbS9VWRBpUE1
xHEP7G3UVLZ9KQexlvbejfKCYxWGg6s9bvGZT6Xk93K+xJsPHdZb5mwOvkbOSDyjekSevzDf4zk+
QQg6BUiKONteSnW6vlOo4gvlG6Ii/76jpKe2iZWbIuzSrErAJOoCeVbzyYCyIjUDDsltzjHSq75l
25DrqnGpD2ly3Qu6rrvmZDjyk7Dp6e2BdnJJ4C1oiHW3f/QY0jDCQokZbs9kl2SfzpI488F6SDOM
1LtIg6cZ+MuZqYGPoRkELu0BfuKfMEDU5U5VDHZfS4lugzrj6J4RJgo64RA78UPqpCbT2FJiwFCc
+rbKf3B+SpMsyJJnOMlVyxOGXIlHBrY2nmqfpwm9E4tgCWeOF6PKdqPQvl6tJsGbQL2G3mJwYgMQ
VC1wgcsWXnGx49+9dJVxRFFKZSWHWAZjT9sDOHvHW9gsWGCGCjDnLarHPO6JUfuz8kcs5WJ39I34
3Maq7kjci8BSPr0hmdewgBFhg+ZYg+b+PW3zc8YYUrWJdJ2YTR7A5Q1cZZlCsz7swrONgD0LLfxd
DKqS4Ipdc4xcnn5E+tiI0v7xwKt9naZSK1+E7HH5RB8K20xjv55CRmYNR6mDUeDgWeDlvOYZS/1N
VsNTxKjuFLqOsonLuhYtPbs3opxsj/fWP9BWppBi/KXId1s6ntBVpl3bizFdtTy6O5V7BmmGCVEn
UfIOTLcKaBdfRVwVHhze9F7+Sb4gYQy7KrhaGM3MeHUok+Bui5UlUsI3FQpa5JXenuKq5V+iXTcO
hYhC3iWNwFnLQcdcD+3gABZF9QrDGqz8XUeoLfaWZ+hFcMFTyN3K9jmUj8OXLhviAa3tY0fN7VBI
4EqVAbug31U1PL+JUoFsOV4ATmRfOZtAyLqB84q+bqAY+v53uMpM1wpZKsJJnx7mAC314cbC5cgP
ojF+3INxdrLtfot67MS/it/msP26U/ywlI85l+hHMkoGjUz/rgWivFSzXZrf3XY/4pho8rJs+l7L
34q/H9UjgsvqaFRv1XEL/6gNQNDQXFZtCHFGvEadY4OZeqsw/KxacdK8D1hEs2/mws6r+sk3GF27
FlddX1D9F65AeMohv83DNA9MzAu5MsI4dMWcr5OcPGm0Cmfu966NLyK4Ot/icTsrTVcoOOZovEcq
hh3Ak45YBrlNQSLHuZ63DI6XkEk9ypVaIGgEtngRzE1rfCuJ2ZLBu3Da54Aa9QB5b4lxALRxXTKZ
Ly9Sld1egdXQEIAeVlnsiCcoXFq4IYaDJnyWwctI+3mlnd9BHZuz+SMiiH47y1mCt/vwI7GG6rFj
L3OKwraVtHfMZOaUTPxoNnSm2HSe7DoT4HEWWCPtRuMqANB22iQi10JmehQi/v2yD/kEupOwXZ7s
ypwWuCRc6VY7sHMp7Zq/Gb9IKOl9phSOncAyaZc7JXohP68T7r1wbF/3Sy6vywJipn87d/teRO80
E2WCaXv/ZzrP84YuZOSx3RUXhaHF/+R4BMNrzucqDU8kEkMcEDSeyfMvTnG/ex5XYM2G/A61NSCj
mZfLs+MxC3dyCd3fy8G8M4TWAQilPsP/bcgkej0zN2+ZCpUCOU7gLiUtyWq7IcTvDZO559bc4tDr
E5hfH4uhucU3YfHAWm4SZzELTIqaba3Ta9bauJbe4NYAWYFjDOtoH17W3LUVSJbahbFw1onzjvtL
SP0jn79v/HRb5MgjXVN58JbtNuKAxoYam3Adkku0dFZxmVw/ctCROon80otEaYl73IOL3hroNmpJ
ucGcu8erT7yKGGgFv07bhNOW5V9K0+EzWvCO4XhUoZk2umjHEtDEUa4bF0L7wAMQGo4tqKBl1E0v
yqWyAjkgzUmqdFjBmHvRd8DB0WhwiY2kZGrBNMaAz/2JpNIEgEnc9CpbEh0r6m6pEWSyWEQ5Rnz2
zLY+MHOPrjAi6rbIW64zfp6ZifaJz1pOgboBDC7bAyDZVGmW/42BkSHs7lo0SUbrThnRlJr+uZCn
86kY8vvBS3cYlyAL623t1gdhIBwpst8MOF2j/Rw3L0Qs1kiGjCMYQ2vTWtDdsMfuzHMZcFPJOado
U9tx7p4lqyp/PYvmkqDll+LJC1c/fce7I6905fwMTH9XXYhTEhUR2t0/HdzGhjB56kNM2wYYSrR0
1roAS8CBjvjlveYWwuTiysRqmVPZ/xOqKgWx/s13OkXVm/MBXDx9a6uFAgWj8+qxJWQNCNT01mSy
5V4C9zMhOrVw3t01qLYSON1mxxQ6lVKMxff7RKQHTg/gf979JK6yLT5wlaQDlyo/pJ3Nu2X7uuc4
QxEvMiCWVwJ2EJjYAsMcinwanbfiJddZhLRT0kMeRX87WTmY0JN+d1Qy5RL83HUItRj29iA8/Zxd
QIwpW+OnPJdhu2GxJSFNW2kh6SKS38KnvEjSXlBekXbfIp1zJIog7P3lPHhZKZhOltZ9Ke54EDcl
GHaZCSKZVRC1KFI6q8kicCyy6PpYBzVakLH+1LpoXY/eRGJQ1FFq2v3jlItZmsuCRJWR41OWfd/T
uwvzD9QLMf3OIxEylar8Sf5dlWFgNgiQcXK5FsgDfOOiA0jSgw2gpwy9BwjyZ8defiavUjh6fepX
f2NveewNN7oQlI3R28+6MZr4sw7zUG2wbku5cD4lmk1q3KnQStBL0llCpusPYAUlSOuzTfa8H5S2
poGwuWNqPsx+8VvlMOtHVD/OGkB7exoNB2l+rUtaMoEaI7MQxZjjaony/Hp/3Q7e+bIGXZdLj0UH
f0OGxpY7pdFVJDXw/5IiOnHut11gMvA2hrD1zn3yL3V6aGa1OTq/h7VHGRxJnqCsIwK0Rnrnnw92
kQZnTdh4F1OOJPVjS2Xy2QHH/VtvFqjmluTmoRzVqNC3tChQzpQMhoyJud1AYgozP+v4LXhLjsYk
BuSjjWNLyNss/gAOPYBfPxPs8BQVhGBg+NgcG1DgcY+niXLUasEALcmIEKZQpTpxWfcktxZTKBnx
tALIlpF6dm+TYUrEo77hupIdto4/o7uGiKPleAODubj1dIgpo1VUEYoeAOOl43tGguml4/OIQy4q
P01kGb6OUSpWkukW406BdKS1szvgvleTaV1E1M4iWJkigiL+qgLDJ2droouezL3Hi0IsSEnsmBQb
MqTeUfe/qMSTwBGi7ngphPu0yg1GXRVPBfvcT4JTNTdw/1Zf/mtxyIeThq/eYdH3FlgOaJ2UbzLL
HqZtFi9z8kFisw6CTfl5UIg2C2A7BYttcQGQDOk7C5FMZ+/q5mw1yn+u/r1AXvTNNCUI+nzfzhXE
KLozY3JMVPX5gSYjZqPVSsxhdSWUPCzZNYM94Lw+oo+fyrTPlY3C4mdjjTdpzkg5ToVFbMhjkL4l
BMhtrItnaAliP2ajB0rAKOJpaRUG0AXtLlJi/wEzJ6txLYhRfTAnWAGuXrS07ptQ7Nd7Vuoc9KIc
mXa5fcj4m0QJ1vU6Hk5oP8qIqYLp3Dja44OR5Plua6Us+sPGtmxbd1/1xUUsQFDJM7yGpF3HhZcJ
YSAXDYMkNzTwI0nNCBw/rC2Y+rShNfFDHtimEVVCphUH0EjaorbTKluuA3E186zz/T9mwW7ochC8
jrl/A9tcup709Xri68xd05tZl96s9w/qrhP1dUrEezgQlNVdkvwgUcMO5wtevrApozKMoQuRkTe0
QwtsZF2iNX57GmCjFWO6ZSrqhdbuM80RsHely1xYQtmRIfSXik8b/EEqsPGb89Nk8BQ0XND+iA9b
GpF+gRajEd7r3D5ueC15xVHn++QKCF8Xhz9ZCoShohC+NbdU6/pDYN1eHmFgLtHn2nx6yS00rFDs
G2nTOBd+HADWfE4Cyj/kssjQ3DfcuMT1iACC2Q1F+kKTafb1fF5R54B/iPjN+hLh1PTxey12m+7G
ynD7kbqWppsrCZ3/bRC6amiM6hlDmiz+4T3Qw91XcW/JKDWbX1jyePy/oT1SRWHrIRvkAOIXwqGj
o1ivsGMLMh5waORvEGvNFSuOG93691Ta6rWThxWIMEhKPQolo8/K0xLnjXG8A6/XUDYbVKtDGn5G
inpIFzimtWprF9HBoOhbkzepLPsG2Jjm1UyWVOIQCvvlcn6yt/3m4+mEF3RhCUFzaMgkfGV+dqQV
Zsj2OCkN4PUMCY6QJT6jzu40ZaZopJ2Pv6S96SIEHDFmYBHqrjInvcdTmgiFdeQP0nGoWuVR+5iU
Uvq5URzWxBiBRMjtx0l16yS0RJy2ewhC1nyVKnTAU/jq1cgHSr63XIpLy5f7/GEMVat5SzsCVyyT
TD6p3aKBP9TZHLBi2KypXtGmbMbwQa1hPldXKcqytwlQWMK3Q3eQBdC3lV0FZ7hiIhohstYagwzp
2JZGChmNNOiXI7fmckobHOyZoVCH8Vwc5qDoxO9OkMioFWSfxyZKK+zxDGb6ch8VR+KvG4EuUBbd
YZDQCe9KjE1q5mhNshkMYPj/4pfpSm+FeM0AssIgm6vInSdA5suqfkfjNcTGxXwRCUyKzwhqWyeo
+ZEAMGS+StUiokr6fnz7dRukdgYhuT9jL7bDaYkGm0VFbmzaBr+E2b/ODjfQSycw4qSPRhTOnfWt
OFI32mqEZLHLRCnypKsA6HNuAl4rKQTbChuCyjFiC6+pn5Sy9pmInF2iAxNPyTYH3HFoxziSUEsU
xgfepfLHgpbUsXwD0GO96cGrVwQWC6U0SCoxXmyWkzm0wNbeJlbm1Ik26uRaX0C01krqHkOp3w6s
fdNDgU7FLMwJ9he7ECbWLTo9c87CYPvak4SBd48LQgfpu1MAZQHvHS3DpMsMlmPXnxuDjdmAf7GI
4W6ceUbSKci2VkYJ+TY3tQyvllBvdu4PscEXV01HECNxJW+AosIyFphOgPXcWv+NHTq8qtnYlEQC
LBeT/kXACbKkXERtYD+aYqxQBDRsk0Mn0m4g1e0XdM+cLtxkTdGi5p1ne3SDv5nA2DvM1jIaH89K
PQn7ynoSAqj7Blyg7wmOOUbz0IJYwcmDMcwDNZcbKgkkjigyBVfjZbIT1ksx0qD9oTTywl8s01s+
PS50iM4LmgWnnf98SDxK/xMArVz/yQ3tHguKhJsLxaqMnUNTlcd4mQrG4gejY+5GdP3i3NtZkSWS
2QaVTVExPid5ubkZoYmVFks0oh7tFiClW20SpJ7LekAbLgTnhllX9MLb/Jzfln3zs0UeOXY7sRWT
1BfCCvmjk8sZcVO1+D8+bM7M4wjyhdSaM2526x21vi6WRTLhU999c5XX0OBx75JbKjTeOPByph9H
F+NDMfn0/OYNjAV9eLVUQUSzzHzy7O2QNZQTbgnYhv90G/iBnZCcVB3EGhjDq33MABj+Y4VwORWa
fEMFSSsIm4SvzaxS2kagRyP+XQS29dvYeOhxkUJUYS95vS7YRvda6fOba0tx2u4vuEen4JAp0vtL
9bmMiTeFNFXrLuS0xEzAM0UKlQYGDnDXhU6ayACmEVmu7edBmOzDlwiXepLA0ABDmDSVXUKS8t6P
8Jtf2qOamRsNnnv+2rVRM2+j4NGQbTfe1s4Fwhvu9LMAtZlhtw/SkidQskachQ+4pDaCYJneO13T
Arm/OcthnU76l8geoOukMmoNA85SZlR3BpNwRsrQ4ap3c3sDPjigcUw/Jg4/gdkrvlQ7+z+svYxM
5BZwYc4OHgFC1ezlinj53D9Zi4QKPvcDW3iY74Bv238GHteim5xkJQOLTFgI5kp1lPdwtkdWv5eI
U0WkFalbPt+2KLiZZz2Wr43W1R/sE5f1sGYfmOzWT2JImhyAIgGjdbi87l1ucxWFUp9UWth9e0iY
dvMBMZCBfRW5S20BUxWpEA5oOpNEIysOJDTm+qtuZz+act0lPr4vqU9xUx8diU/735LJKDXV4GPO
Dc3E0X4DWwp6Krr4OCww6Q6RGz7WvrtyYiPJ1RCtvHdPiMXPnZVRK8c92Mc9ucOArCtfivCKud+q
zBDyCMRTP9D/E03vtQfeKFFzrBNslzpfz1YGtk+NzHyct1jMBczDV6S3a4UTZDZCr7mYi4wpj8CR
r4675EHFyQizJc1k+LiCwhmfahXxQxJSkYCyZFKYdqbiCpMgpkRF21vDRR1fi7okkTxFjrVZYuZk
hGxnpXzOQzE7iOqHk5Bev098w1r23G1Rjngkgf/Jihh+42kQTx4HXNvlwYv8sUD4XfgkvlXDYRn6
EHG/DUdLOMhd11zFyBND4fwO69OKdXNSu2VLrQ+YZCI4ROD5YDEFI18+rMj0TYmk6EI9Hj46d7xo
9ow10p4EKl+zDygJiVm2WiI8MdmQJW7yd3La/I+NKF4aMCUflBLj3nOWqN9kfb/NEfQ4hpkZ65AY
UO54JMUBQV7UQGh3gMWZjQuMBoNsBjSl1hY3TlX4Wy+hyowXfH4ZpPEx/Hg4RUV6aBkjWvSf1ZFc
FSzxALE4p4hmKiRNMjfVssw2WUMSzJWr1nltNoFpiCxDTGlmjxNIIsA5o4QyYWQAU1wO1MSnui72
yB9gCBSxcEuqczLHOqjUAz46xojrUgDwpNxwN/e17gKM4wsUJ1njBLf/YOUX+tV0woy6Gnvs3Ax7
8+1wQw1lSN5e4+on9eRDQcrqbpOD9UmSOmNkqPTKHbuOAEZ0UXWvpYuPNZpYNpWBXZVPaZSgBQM7
xSLSfr/fRBVHFyPY4npP9ljj0j1PFGF5pwzFx6uJQFGYKHWDX0MJeDtLgKsGeg8VJRzF01tnmcKL
wEWIAASpRfS/tvtLSR62izCNQzwXx66ru0YEgO6ORmGmzlfVDansRW++PmQBdPjxS/Y7vTQzb/HL
OvfrhHYSN33rX4J2oYU3fcosajWmYH/lRxkpoHovBU3w9kJfZOfYCxK6bHEokYgduBYrGzRJvBte
xOHeD94VEVOPLOOW7LvMl0VV8tjs8Pd7u1ztVe6K9CZOiVWxrCErUFOHq0Jh6OdwcITKPDa+mK+M
5EAOGu2QmIqm+GkYJrZnR5J2Fk3xsAODUMwtKRsvU9hgML6osghnZ711h3RVvvpoCZleiBQNu/J6
4iE5/lvmV9oUDYwg8VahppJCR9jCNdS20QZVau9am1GJuC21Wo5Ylw4KY9A1Pw045wzc/Qwt3A3i
1BnmtTuz2zDyuknYC3V8gaBKB1KGsZJVu+L7biL7b5JjkVd1/6yNHjSb4YwDSzwv5JfvBGUoqUSZ
8TiZwId9rXnBlNLPWWmOb4CZ/KldvNipBo+Ve43dSLK/1EmaVU+fKK4V9fnbT4vbNW03wnGogRfX
4uOZ/4NtwLaGLP8PzslI8gpEkcoe3Js7ZA3icW5euKnZZ+fZzninIawmFeLJVukvBbOKzrDevCdP
pnksbS/m/s8BV74kQoOnciFQ+mLQGcB3Pp2f6+dmQ/+4oFsAiLTsawvKBZEZjGUEoIGs2ySkotOe
WXqnsR7Dzn2MPF8XeMIeyJVCor7ODyk32QMxQ1ukZvjOITmheO0Qq+4jMqL8+EqpBLHvz2iFui01
dHCREjfogpvLjs8KIuhQzmiBhSxZCQlnaHGEEtFO6Qif7zNmm58rxVdRj6znME0hS0rU43NPqXbS
O08PWRgRd5sjbPlthwbO4JnLPwGw9130SiezH5AnKme3uM946NGmvyTKXbBTp0rc+SgFxYEt/HBu
d/fx8XOf/XcOrsd28g7X6s8AD5NFyPIBBKvYcBzelPKVwBE4FOWbYIyWIQYIlIhDVc+buH6bnGwe
aVInibbGXQ1iB+2jtXXk7qoxJ9Aae0x3hJgu9GqTUu5iHo0L5caqgVytT/EOG93cxpgiuIezhPfH
pEuCTOdvjinp34zubeR6WzXr1rpkgWLvWr94GlD86/iyb8XbLTe9ns2QEN8aXZcmHSDRARDkPTCC
cLfcYIeUXyytN+61sxMmsf1uKLA5sV/PFROETTnRRnfrWped9uSe4/suRdBrftuB2R8nc7cMrQSw
LRMXP5eb/SEXOuZv8MXLcVDqtkOVgJxc9nljf7GM8kQdGeEmmnq2BGmAW72NiQokVBcDS104147i
cf93GqCpKVIkuow26B6BSVpGAGHNQpAivOJOQUl3oe6Brxx2y9bDLOA5mAKWxOwqh3AW6KNAS+gl
Np3J+xOr95baOscH+zStUMiEi6QXcpySU6ujS/XbbVqX+RoqNqSfohZ4xvWRn0dpnFYBYwXA3GB8
vnEQPsZI8z8ZSLZZSpTn0Wdq+8pkCrPDJl89J3YfhHMUWaHAnHCXjpOH8D2o6AEYUqoK0dTU5NrP
fqsnYTgUyW3IsGQBwxisHPRw3CzZgKjaxSt19UYma1eZrtNEoq8MCSA0harcGUcnS5uwG46fhn4j
J1I2WBO+c/zTM7MINyVcCq5H2f8Tfp5/8DNnfE9Ee2c0zz95goW4Md/z3KL1MfWecwSYRJkS2JXg
6vw0IiHiMhs6USBeITLWk35Av4UvmeIH+o27nDdLQC3/i1PeXJoyOl/6TySNr2G9y0/EOL9uq/or
NntvJow3/uEGzqKGbtS3m3zttjfDf1IMDXFhsUqE4Pc/TCONSOmeeaQs/usxiDDel951Mx0zbRhK
7KXAcoj7Q7D2DX7yOmA49aoEpp0pMaOrEdRkHSi3gjSu9jo5xaf0A9LWeDlIqLOlM1OOvkAZHaGm
HNP7gUp+6AOMSxFFU9E3KaCPMnyrMAJbc690pdcnXmhYD903ehTLtQuVbymBKo+NlXWAjunEKFes
4fofqcydy/eJGLBgD6NlTTf695zmEyTJkA64fH3lmMhqVNKauLYoFSOS5LT4rS0YJPcib6bC9epa
WntfZuEcPb0J9dXa1wCxZQeSCcossTz277KYBMUzchzXqyA8ezimN0TWrHuyMPbhR0KDKqdCYfwG
ZpQno5eS2qYN8EOZxhcjsuJ4MJX48OCZSvUJu8tGaMUyQO7NMJjd/Zr0fSjCXdQDFvwuz/5t8tiW
6dc13+VCH4LD8qUWioTzkYEOehtLk4qYARrorVnvCTC/OSOmjUGxuJw2dohlLzSwk2EVlFH5M+TF
qBz8PY3me3nQzgENvU8ASLFaXV3eyzRlvp2ySoMbnjcpSeBeWRrj1l+N4MW6om2qpxtbK9VEUPYq
1C4A16UK3k6grVAf4oTDuUR/xuOsJ8oVv3Q1UPaYTdVZsNJf+gvelfx+xIGrgE0M8gvOJ4h7Hir0
58fQvqe5WLj21SASqOBxuMDFIbXnGy9h6G4JtjELhocybCdQZox1woXz8ZOW3peVN5Nml3Jhaxnf
kqNXj+eO1vPObjoZyl6I6DrzTf5cbxhrN2DH7tfP+mac1IHFzwSF45aikV51Fj1hXI71UDHnus4l
lGvMxwvrJjK0LXU/ioo+/BzWEBVs+hjyZ61xEtLdIDVUOMPiC7Uex+QSol52++qhSYGRzH5fRvrz
LjhCd8xPpnF7f8D3N3OyU/bF/79gWvuwjlujq6CctvYPmQKHGtd8Yz3vNLnc4MWUZPy//T+1mx5W
SQMiLSeTPBOIhgRL1MNFI/zHEJBSknpaQ21knYF+LL4xBF+XBVSaoPOFTIwSzF0WSJ6Py6kXkGAh
EeyRsRyHwvchdcSxwul020h5BJb0vGuquyuJo/Z1UZIt52ykhWM1O3ZCDV0EuzcFAuqiZlftfg+j
IZLcz64cwl8u0X4nTe6uS/HgOVcSRlN2xiV7rwDmqdHqU4ri1BtU3j9JtJwR3Fy/qQdRdyTdJRkU
pj7tfpIv2xiRsXv1bOtHvdAIV9b9Zs4eyiG4Qa2ifrbx//i5mF5j7Q4mhZL4JqFCRGtJG4Oe4kh6
s+3NwxX4mAy/3hz78GEdrkZLW3SF5jEhkrz29hgVNPHyG/3CdfR7naAIjciyR9cb333EFBtiwjHX
y6tBgAYneVR/Wmop767nDG65vlq6gg==
`protect end_protected
