-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SnNtSIWYyEb17LFNwB2v/ZEMp6kXXjzGN0InTtPHBYawq7VTlX3KpEQd7BIYWb1oJYuWUmNgTRr6
GMptRDQFEqRBh83BPaDfW07jcJVeSWNkfeUug3HbETLXV9fOXYenY90OcJEYNAIisuaBg0E6EQNp
xrt1X0dkjuJEdCbf4uUDSyOkl653F86LkwiAZoGQg0zcfQxshdJyHNUB6wvYgn8oghtnRtsUR3Q2
TflTkeii98jSfSnrydYkflippIujzASkFjokID/fw+HQuumE3D2phNsi/yhAyoJXyITsMRLJYa7U
NnW9YTNXeCO43tL1lqB4O1pv/dPvYeTCpQHiig==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13856)
`protect data_block
HEf9ihXNxOmwdEMpkVQnFOiAuBcoFhE5fTdxnWZWki8QDyNO4+kLRswMIqnb01hrlaPwYVmT0Cg7
ntNY2FiH2RG8IMk3wDWZcGmqqcNnlnxnUR2mzvjlYjj0L3LIHuJ0aVOs8y09QbbQ78+uD2tNrnBK
n47FX51On9luBF/+nne23GgzpSKBW3gHGHMoovpHc9e1bf2sWKWCk88DD1jR7VDFvKV+jBuBPygh
3kCK3rdyhkA2e5XvxLtC10tP+PU+kFenILVE8Ro08qtHdavslaKXsfgm8xCSEa3SDq6V41smwHjg
wXtGDrYmv+8+oV9pmAlNqr2Led1MFDseAwOoiv20MtEe08tQUaADJqm00H4OB7YaG218MXnHfwPB
H2IGxk05GzKFF4t8ztPRgNW8w7FucfxKTJsNWfR1vLZLA/QUBpo21O0GBCxZj6I+tYho7Ks8zJzC
tqEn8KUIMNVQqej39o+BcWIzrMGqZO3jnDtLpTyb6HwIEC6d0PVGJGhNzZSo9AIQmht8bBTpgI64
eq0bRHhLKK8TDXQq78wtxBXF71a+iO6G7bPZ4QW3QrffL9GHJrC7Y33XiY1Fp/vjBh4fPN0zpsnY
zJ7ZaF+JTrqnjxIrfU+qmFcXqF9dGJggmCJmbd2jVTz7SBV+dsOtG04k/kFjcale13bIwj5DhSIQ
2Y7Z9xACb9R/6nPMO8e25SNdQNZge1K82VJrMFROxODRgQ0dtvstNbklVXBWqcgAwNSXziJXtgFg
j1Fzay4d/JaLRjq2vSktpeEv2+GrWZ1gPTZsALwE08OGLs25sl4kQ+AcyNF8qjlp/kF+SbZB+qO/
q00g9sETUydMngFHSnHxpRn3lVvM+L9qudnm9s2ZdgXBkFKPaPXr4DZIgHZjfXMVFJtKDvex5GYT
k+IQUEWY53jPoU8tyHVmAda1wJ9jtJ4bUp/6SHwlQ1eA6RJO4GenxQjH7+aBPIwRaUM5/sHMTkMU
2QJJwxWVujPxlZBoxu8yXcIvvIsaQ2/ZbJ8yGCfmpfXaaWS23sXR62+sSQ/jmcyhZQpju1nuLS+c
mOalSJXrjkKxd4BvihrM0jEOmgg46GX61eI0cjzFJXG//hRiQmfg377QplC3sYhrI+597qmFRTXA
rPldOKcLKD7Bwp07CpSEID+cKbDcxUSNQ9o+/vLNyXof2BXbPlHzhwOB8fWD1C5TXK9PPKuOFs+w
WYKNyFyVDMnmVkzL8KbtUZy1NJzhXS+sHV/ovsSypFES+vvsjPqg3AQE5UDbTEZo/eyrnpC6qM3k
3oCbrBNtkol6fR5zxQn/wRtA9MAY9oufcRgBoCZ1aGrChH3cJQ4wn6oxGBCRyyT/m6xGg5rei/Dk
YkFYTrsGLq2tUta5c+jW1RxE6dgn0UC74etE0yxq9OMveubfVIBGaC5EDbfzaU0+d2Ci2Xji/s6i
jQQDRyh56+x17kaUFCbr2Gz0B3U9EQHYdovck5b4XLz7AdTcg4iwJnTe4u0eTr4ADM/FKxpfImHD
WtjW5MbW2neKkCZQjILcrpRM16w7Dp69czMkJ/lqFtgXsuIBbWrZyemUAqHbZ697B5+Yc5BqUzGk
eDFLXNyeK61xf6UJxOcYOAoOvAsW4lU9Ubx3XHf2EN7MGDmDSDaIWqwkZvza1rYqLXWKVxH2XKdV
YUXC0SXQo6bytDfUvlDsfYdrQbxHhsuJbOUfUG7GQ8O7BsZ+4kme95yyrStoflwZawRgxB0lD7Wd
2UR2M1cKg7RW6Br/Rg5ILcQfcPL5TLPKvHEjSW2l0yRr49LbuZ0xvTSsGUZJQvXC0gH8SVnHh5N9
apdXG8ZBzOWGbPzQrT6XG6SulnSCusnBB94rsyslmVVAHx1yGYczpNv0/urFGhyewCeT4Zc9zkcz
AK3EUoEt+tXnnebCZQXYLifbn6+uCg7CqWC+UkYn/D7uoE/pUaxcZxL6iY0AGT6jc/hkiHJHw0Lu
+CxCe+Yo6Q4C48zDbM+sq6zgT8r0O5HixKAJMvg4IRSIa+ZiLL8xrmT7jTHLkjOxoDAR9A3hzpa6
ejXL+NKtPeQK0/PCypTrYaEh0oayWnS4z9qyxdg7X6HgrENB8VrcrtNgpwtMfwuRWrR4YZ6VqwlU
S7dH1TyOJt+eCBNgpaKCjIyMW33tX9ZjNXZ58BRcNApgFs7c35+t05Gib7wVmNtc+kecVFguNzUd
i1ZiC4WmzwMlTQA9O75fSZy+r7re/FqOvH7DOOhVjuUAoQvMrDhQacBymd8EEK/NQ5ZQeg8wBXdZ
CITZMUmdyE0qfHuGrYnNIBs4RLjb+G2kr3Zm0+Dv2sbRphvRjRnOIMzNfq3PxVp5YgjBWYZN+Yk+
qSExvJs3EssnUZH9/Wcm1FtUHa+apth9Bt/AYSVcZ0X4ej32uINaANNO+tNTpQWz25umlLkapwk1
ZZCQOqQs9FlIdysJmB1vDELdQU2w1syjJvYuX1xlgSDO+MOuNXpLWD2sORr96Bi7cuqQtebNY9qM
EyIXGgbZDQoAs8MTm0/XmMQjBmKP+FskvSmWOnlZ51v2FjdufH8NWpy5zW3iJyPrNQDz/SzBPzfx
MahM8pr9rsH6e7i5VNEU25mAEamwZ75aLVfznaxn+/mA52BKUkgRUG7SBkB2io2giSGBDwMKa3Vb
EzEP+b5oQNx5eoepT6AQyg6UlbK4NEjt/2FcgY854H385bw7wbsxxRR+moCqRHkNDoLnc8++VbaM
jE4PZQrgbYaExLlyH9wHrxL86G+jzR2bPJ1XDauevKvN6y59dqer2LuXSce8/FQwkBgWJ4bxuRLR
2CHNWko4LFCvfL4Ezf33xkEmpT+YmslmOg+OAUO692TYiakaHI46KY6qqhdfv4BMnfxzPL3wpQ/Q
BAKOQamo37cbN5XvrZI9WyuWWRvRxjhqLiML4XuiVU4m16Ha933FvdBG46GQC1ujZ/b3igIouFP+
sb4rfki14tWv6eSgU3e3HSkQuGozyDtP7Uc0QzErnL1ym9SxW0ZCfdv1DQ+MmTyuM2a3xcY/gTIZ
9m5JWCoCPiT7H7zUQMqOrmabURcaSxDCwtNrWABLTtpl2iT+EMVbeXRd/z4yTqcMGSg4u7/eLs1l
9uz8aFRQxdEn449YbNRBu2GnzSI040BuobfySH/e6JCIRHgF3jgTj4qaZgUW/0rQelRyECeTR0T9
bffW74WKju3svd5sWgmTcv3llde26iJzQwCz6oEAH5E3vMR5OBlZhlfL782jWi1sm4n2Q8s+EC2P
6ZmbyE6ICwUjyeSREPhSV05f/dKB6LThmAf/WNq40RZUECuGAyfHNDEQCJ+Gs0Eid/oePFfsu2I9
34EbY8mRUktUk6oCTJ+PDTt1xE2txrd72k79vRYs9XiyO/VAWoFr4NT9xo90JT3pPMYB4uvrtXO8
5WBRPKu0As1Y3q61y1JXoyDba3isE1E/f922XLCiMWMl3ZxSdIjYUCm64TRE85twMzSuVgMinxvQ
n9PuMYx9goXld2Z/JG4CXcNXohTlJOfkvueXcxijvJo7pFOIiF7gQ6OII/YoboPcLm9Wuef9/Wgi
Tf0qHZ23W9f7vpXN1uK3wCE8t+45zteXwAMUX1N2vTLTab7Hz0xHWmzi18eWLaphXq4WJ5x5TiIA
DoiyKqgmQhjjT7n8PeZaZ3eXVIRcz6n/Zx/0qLkxWoNjCAMAvkpXryKguUu8Bxul1vv47XV23LTC
3T6kYO8I7OYE6Ueo46/yEnlg4BdwfxPqL0JE42g/vTAT06fNn0jIBX7gacj9YOEa7HsPrtdlV6Bv
UuiZUvJTfZ5Eyo3D9rzoOcp1jYNUweZIDx/D3ppenGkupxcvcFyoBuwqixFTpsDbsdB3NAmv2R85
ZUJUwQULYdw3aeq1/LEt7KuQZjeNIKpPnXojZnm8ZNr22kncwQgwBsUd1P/CRnYNYW4qRcAjiEJ1
+n+FF/1fD8vWpvcGP4OCeIrBB4JNncQTsTDzdwfVRgFBcZSkUoa95fFbKiq/JgNcxPwYqcS3tp9Q
OQ+V+fsKwJfhKFDmdxI0HEPAGLa/ZTG5dSK2JJQQHfNP2UzTLHkNf2hHKaux/G/D6q6GqSAaQ3jo
jlrQjB6qdy8rUoeSuBiMiZWklsRm+oqbORVcronPWvuf76yBjl8Y2m9jiUDZm2y1laXLYsfqbuEE
hA8B0OIUl5HJd+GxxkccO6D9Ql3gROyZPIe7VK6P4thq3+zFb/VjaHg7cootBGBDHHmlVbnvigeF
06ykWyfD4hqlFkNJBvXViu6Fe6bISXpw2C8170f7qtH8LoR8V91XuLqiwBI1FS08fr+OrPG3jwWX
4cNAfXbOJx/ektE/+0PSC394E5JndCaZGskWP908/LyXviOifCj1STEpbrHYe2hFgn7rw+n76jt7
yLorIQCulhNbTVFeuy+RusEFBa/jzI3DDc6Jj/kE8SBczcIS5yrHVaSagmsxawtyg0dKKmmOEf7/
NG1v34u0F9pViPsac5fc8q5RdU/6zM+vUVsCNW/cD8kwKLpN/294c/PHwi5vahjHwRgtObPBW9TR
eqebBpIG+VWQg2+h5LSd1J+E3zDh3M+bHxuSyRwY9hvL2d/uT6aHTE4HYdSqeeSUF5cIoIgUn3dx
G7r2UguMF2tOumOSf8DBVn9nxQBHhgnzhzzSycAintB0Hu5cUg7ty7LmknR6oqRYeoXH2CMOLSnR
uYTn908IbGzZXZ/2RteBFDNx854hdQ8/tv8v4JOChguP8rcXFME/zE7jp5uOOS2sYj6fKi/zYpG0
nmeobUu3T6NscwjJTFMqHCl9mMLmG0drCMwIAU9bBga4DzDrYme4ghcQFVjP2K+u6qvBujnZGEoM
RSeeYT/cxkepwR3/0JiDu+Py4S4OER5qp7m/WJL967UBHFAKQQYPafI75aFaXGFsfYdYmGEWDI+O
tAZa+RMrpIf6y8ks1L/teo/Ur7ZkpoLsSRdITulKXyZUoFCWkIsWEKYpecsey25faUP7A0JQ1BBc
pUAcV5yCRt/3hVj7XEXcwCucXE4U54KEQS15Z5u3bmMbajxKGNW0OxljN32Af6jDv5YuZlzJcWTE
rurY/Q0xbmkOuOw0RXdDkUlNfttCvTPll07wuEftcaPts8H3zX+SYfZVBklbjzvl6iba73z97bCE
oTYoeSbCMwoSfz65G2SeTI30fRYKukcVVdxpDh7oPFza14dN2Pn6POIzi76P2QQrkuzlwc0PRXHj
gc/VGBUZjFV7egoqg7ZnbT7aVuOy7r9BgKK3iTu7lzWsegSV8OTZtwUUOjvpNMdj0tpOCOjZ54Ff
Tyv6Djj1pGDRgpiRaLXgTmCTerYAtg2DcERR2L7O6TaKu8Poeg/zEPpy6o2ileFI2wpZSh5/bHvH
WviAAmCOqKn4DF2LpB79o+UP6XbzVZxHWpiAQz94vW3Jlh48oqIZzts3aWdPnCCRQj9j7A3lR61q
ixk2AD478OkAFsUskfnQfx3n3QLgnUB+Nz1WzkOX4VBIbrofSK7Rk5EQ/HUXFxn4D7FqGsjFIpf1
MJH8pBr3aFghvhQDP8Ftv2kUNbrhvoS8BWdW8kUa4G3v6wpY5AQVTA7LtLM7OZqfductO4WpTgP5
3zRVFJjagbbYkJYUMuI5mMKYjSpsFAdW8wBmwtndA7b33rxutmRcfMRJEWfH3pSVT3SGFQOUZaLV
76Tm6Woy43o/Pcggy6yYDOEiuk+pupDaq0E7Y3BI0dYUVvHEhqpm/2WS0v22HoOgfT0BphRSNt+s
Trww2y2mHt++m6jt8BOwZIHo7GAdpyYEO6zZcEC+AD1KVEPcxM2Ie5V9UoPXCU/Eb3qwCKms/lYK
OCKN7QsGMD8vw1Ile3oNasl5jLS/ylBSI++lzegCjGE3EhI+384q+gNmHTBIJif0KmnIWcl7MHpd
rCyooZ3MyhvmDZTRCWdJQOT6cIheIEXFwhGtlHtCmkuSNpZHqYiAc6+Czwn1gKWd0qtJBzBNNHYE
cYIc+xW4JpSOGGK+zNito46eRibnXcokOFgn9DRZnPOPa4bONdfAdVUkTVQOyzjaYd2dBC5xTq5a
+IvHl5+IDDbC4AjUDxq/+KeyQysv+o6An9NNHQUJ0mrltVoemRZG7PU2bobFSh7QnAxqYo9icofr
F8xb1CGYDlRlGkN9xr6GeTLdZ7vm+Y8LeEPDnhOkRUa6KCUI79E38HSXEpFvGu6KQsMiSsEgnI7v
1O8l5s88pvq8MXiGRMoiohZFaRaGhL5HO46XkxYD19Y66y6gegH/Hb70gD2ALqZqfZF67Vq4vfzF
V3cR/zCfnlbGbYTCBBbOq3sEMNTvDRH6q7Hdaxkr/XOolBzXa/o1RYMhZFVXX3jVv/Exul3pGvPK
di8xh9/bzJLw4+clDCtbSJU6RuQflL/RUWuX4G8T2LtnX9WzBATz1YHQizPtJfKFh83BP9osgaDV
7k7VdLk6Y8ea1yt0DizG/Aw7ZcsoPBzTQtsVY9Ks2bjMjPlCWwkF0JvY/ynUmGMkTus/dSLYzwWN
zYu+z24OKpqkMyNsezh8WBj5LMIXJlFPavaFZZAaY+xp1bDNVq9hjpsOkm+hmWajxd6NJwLui5jb
/9/bFMulMqLMoRLr/kga5QSq3d70Hgb663KLpgmiRcgqgWFFbskuopCg+n/YjFbWLuDEnkL4URad
dTbcvDRDbsettRJi+3xw7rHejhv15C+9MUdOEysTiwXlujiQ08r8JCkKjYSNxIY7B7w93Z0yZwsB
hRnh4ScAwsJyswRGSzqFloNRuXKsWiA9QRl6Qb7YiIZjmfppAKn1FI3AoQ3WIozYOJ3qZCBG3+fJ
QSiLOHecCnbzh1wJA2GCNwwCIU6nO04zAt4tefHjbHRi/YhgpKfWJhYxi2oDZzgD5468O4SvS5iP
VN7wvXr6uyvW6t+cm9F4LUp/z4jkuqXo46XrxOOvDnFwzqhfjOlGpo5+vbpIAZf33jx8uFEbkdol
Wugi9/AxD6oZT8RC+Lg/2Hfp//9pLg6CxgLYruMu9eUU5qkJZFzdQm1Au08bEG7ar3y1qG4TzAaC
PiWDiv1vzi2gjq35lLVfy+BrQtT4HdQ16tL4KM4CYiq7Wll0AO5JU7a3MgcEdTPbjcb+g/x8kcLS
q6QhCNm6piTC2K5sKPV2un7v73eomfL1hb9/c+tvkGPuy/X0abnZ5FHUzXm43CXvyHM7oonVV54n
vgfKenchE0KjUS2etR+VyyAX6RJ4XsMvJ+hEKTUSw5gvdBKuhcWBJZbEEdAYje8FpRjgE+mEgWl1
LJD/NApKvnr4fid9bSBIRAnNFsctph12/frTET1/OW7in1bApFHo9/Do8B01ZzNSkLTgoFRSXzPJ
wZGKLtIrfpVi85XLdJeVu6XWjpGBsLFxsZx14NIjsmDfF29j32xFLQm2agzUjcXfoiQsWi5NtD9O
SVmECOr6O69vVvXHzEvvLPUCTicGPcNPwSnJ+w1wbLmYAV0xDpSBCu7eZEScrC99xGSpqHpxgm3y
1JJD6ANiCKCXvZ9oXLHE4ADvwpKwJCH0OUv6cfZ2ShHI8NrCxkfpD7Zp0Hkw59xv2k1mYbkE2+eD
okyD6s0qJLdnZRwr2lqMgay1NE0Tn0P2uV/kQkYuUiCkLL4DFOMBMJtO8PMyOAClgYV4+aEoimJ9
vpY9wkocm5FPRD8thH7mJYqx9NLgQNxv5x0nC3B8ZI0tG+1Ry4Ge6jrOLUjoNg3C8XlMNxaZvt6n
sMPUK2s+CDKwu7+V1QXJfofasarv3KlALwx5Ws4UBtoKXZu6Tgz3kLzI4gMFDe9RlK3ubTmeMl+y
UKoPxoaRlr7E+TlsHsgLAHTBY/obRfPOOsSWEfllEfwfaBOeFuYA+HJSgPe5EBZdzFD7GVkH9iTb
ihgpmQkxWouJrYCoUDpQGW2PC0BhbPI4P98CMQrgK+bj9BPeSoNZu1+MySVyKPrcq4mm0Du7Z1Qc
596lO9QyUZO7qnQDS5xwRHmelfWZ7KegJCyuO1dXWYVA2S6yYjrzGme+1DhxNsNdipoj38m+SxRE
G4G3acbT4YTTn2kQBS4Do8qJHvjAilv9aCHeYhbFcZZb0sq88Nrd5909iXQPhgsj9gqP6UL1JTT9
Rk/LLprlMRxc2uwE2oct2rAusSQcX0sPupd5WtiXe2OlJXSRcDXsuSEW+qmUNHUlJoy1ZuwmE6Pt
k6TRcziGLzWLpcIyf4P96eMeLOaZTV4r7Xy9sNT/snrHl/7doBm+pY3WFeObj/hDeUF5y8fD8APz
LzVeTJDZcPQdxzJbCcXEnmrKKCZFcpt8VyKnV18gmUgz+b7DqI95fQ1ZlaH2BJz7QRi1vh4PF9f+
Fug/wtf7pYM2tJOr8s0uLK4Pak0o6K8D9c8xJ2m+4l8KSF3nQcVU5rKpVXfvpYbjifb/rKfoeIfW
9NbU3wA51J84ZZTGaMLrBXFMe7aANuJFndhVOYb1K9dqtRiXpYJFgKPZMXBHXuEy1IH4IMQ5HmbE
Y86smnTqUdtPGGUvdzVb8lMvEpIgJn4MyBAQ0iyVI0IDJVrtjfKY2pMajsm23Z0IB6wyRVswZkxr
nOErC9PqCI+VmIWQh9xdHhbgzQT7YN+6kNRm+gt6gZvjL4V57uA4ORHrm2Fp0GII3qLNHQHgLP7L
gRXNlRxPfT9FGodcMRKR6r8NuW/RCPTAzJORV5cbz2FJKj6CDsAkCXtj/CvpdEIMLwaTIY56dm+O
EedWOOw6SSpwLuHYCuJ4rerRI9j9fxlJd6HIPNWDhWf4c1xL2HCL0yEngKXdGy//3oSlQv5zdKa7
tak9QemnLl4s27ThYoanZe9nIuVIdSscddyFcGKVm4WVIFWoab1marDbX3d60k2vKiP9V/6z7/dz
YNUwLz8j1U58YqBNFRxb2qUdxSko1Z/q9Hwhw/l5Yod231xXmGa+PUiKWNKa1l73bG1VczU88O1h
M0W9CR2eCPlAfIrL6O+MaB/uBp9NEHeXMw5FZKTEeQ4Q7UbYa+6dZY5LZOROXbfA/E45dkjGXFB8
jUyn0wBhehBAIGBPgpOyr4GzFC04uFhgHBqXq9w/3F4J/cVTePWDzuSxuFhX2Zv3rA0m/1FUgYGa
JxaspOsTarcWceppEw6knZ8dU4rkdgE6rsfXM7p9oQ2gjqS3RTaRAd5jvii+bAantwP9duedHhM7
a9tuO48qcfGIHJeKO6ww/Wmu8cWWa+/AZaNXe9xxIEu00nsvquwK346P80ANMLFDI0i2/3kF+bKL
D6tapjlkvgUKnraIuDd55uaOiOXhsncb1o8bSSWON/MFDlb35dc8eJ7ShQtyxeZIYOWUMQ7M+qnR
5NZ0UL+8wc/yHWGVoMTgo4mVgj96JV106ffAIHCjCzOlbaveSs4CQtwtbU76b17KY75RF5BtTD2U
yJlk4dA+lVW3+83/qMRAaEEJjD8DS8JdIiVyjgWs0R0x2ODXchDFaeqX8FE8pm8ARkIFHDU+/Ggp
6qZDeZGM34U79gguy8iIlXSCzusKC2l8eRpbXbMhLiHteekoSuhNzye6vmo8+w6epVrgaeobw+aQ
Pv2UwLh0M0AdMUG7vw2b5L9+A8A/Iczz+rHBGwLYuGuNic5GGQxcX9GnljfbJrn4STQ3OeJiGwXR
cmCbFWA8y3Vs6d5e/rQl7DPaQx+Q40vzNHXnium3qUxas2u/0yaMSqaY7d3SPF01bPzXNcFn2tUZ
JV0RIbh+OpdWR7Q2/AneT1XLXCFlZx1KksiJ6lzq2T1y4S5knfDGoz5wo4TW20L/yeFJ2x61e7D4
Ju8toyA11+fqB7UsiIuXa9hrgRZrIz87XJ8tXQQqxTyGnBPs9cDERVqrawuJBHYtY7agsCX8zVss
RmYGFHIS6KrK5E7Enolv16AZWrCvGdYzo677YGQu0chrF0bvXAUvuhBsrOJx7YoO7x+fS821xj9I
ml5lw6jAHsdNuqOSFEAk+7ZN/DeEqqLvcZopgDxS11b0FpbbphkZN/j2h7Wn76SQBKp7UHygC48w
tK2RbksDCTMXsDPYyOHDwX/aRVId52hu7GvQXFiDqz342x28kcc/L4BlO8nu+Vo6Eoi9rQ/iG4KO
KokXo9TEmayhNTR3ODqSeL1Oc/nZkM4ArB42lcbOTN2JeMG6ffIbNKqoN1534aQzbzRuJEPp8Fhz
n0+690Dki4YkIH+BfxwfmNG5aAMscym3f/iWxZx0f6mcelh1MHt3jRKX9mDwf74B8dF7BgskHyDS
qlMAs7E4K6T+V4pwOgOROfI7AkB9iEbzKEHSQVgk5Dl1tLUDmGvyFUOa51hcERBUFYwP7d1iiquc
7sdXPCHC6vKF1qD2iuxsZYtmBpGYuNKpPmKboRHZ+959FhOATBP4BksFeQlu0LB33UbInG7gGsCf
uxIDmM0ckKp3t+9SPZskGQlNGz0Sof73aCGbh65eHERuU+sdCzLXT3JzLM92YKFbSWkDnKuVCxGj
r2QsJv0hMfBlCTJXIPT1oVV9qaidU5vapOvcuVyV1QPJ2O1HACmf5ubvBBdSscyBXcDmebF4yjg3
kQkAIveOCNYoEBQGDYNHZ2BtumDUc8vp3ELEeCtbDr4KXANYa2ocf81IcvgwtZsV/tTLtUe85uyS
573+GjYy5UJaylmYgOm0jrDf5UjRxih1pw4ElU0C3dbzk4sY3WcLGEHGhRU4GEDmVE8YfBETMe2C
LVytHZ7lgOTwcAHBsOyoHJNshYZeMT1dNE1O94rhOnifN3XFkzqwy9pZpzct3LI9TnOlG7Nahz34
R0i1qlwu1qm0Yl3g+3i8G4wTML4MdvnRoOLL7RCcCD0Go2Q0H5sZP7Fs5TDsB2u5pdSd/OKD2RcN
hhThDasA9MNFoX/0DGvECbMevtwgEB2pd3/xme/L86jt6CMLA0fjvrJcWaeXkJHWTRjnOi0NwX3Z
cTOwgkKHcBnaEUUmv9yBmZs/VRdFi23XUOuZ7TKjzQObUsbtxil139JxWTi5gW2AgpI9zYTEjIZO
aLQ752VL26FZJgot6c6BX8kQclNGZmBq3c+gjOGh2KKcXY1i2dxUO4ETUILmkCwMlvKm9nl1p1Hd
6nd8weKQJ3tDV9wZ20H/KG2bws1yS1TH8U0JtUcMgx20SOblHhYVE5wczroM6rN/bj2GTMSXj7Ku
iYXlvUvpx2grUtHVJYrAW8nB7WChRFX5lcSoCvCY0563beLQiVzn9uui9aQ/P1mZ5WC+ic6bfa+H
YHkjsvy/7tSWYB6lF9CL5SXEzsejGh2ssAiujRNVh7xDMoPIVHGlnOqB3LPan9j31iGib24kkTCn
SBBc4VmH96EM5KQW08R9AQdGiU7OneXVCnRuE5WP7zKzFpReGUiZ2cBoz/zFcFqbOZWAiYuZHNHj
Ei0hl41IDJ+dBC1RRaSVk2AhB8KSBrRI44vSZMDuaf2XDsy1SoH2/iycg7boTWl3fZS7I+6F5xOx
w7LbmCWGR93rc21l0f3/jScxAZH9uCRLtINz9EKacjbtJKXiBdmH1uyu/DrAszGs4jU7qwfLNiKo
CH5K6TS1xOoxsfXeYLir0YDcRxI2sB0uTg5JHYpYHoyzKw/zFVEAvf3ygoxRIoIY5eA8M2YUQZ9A
1r5+bTWZL/B2hXD1snsEjO1wCvknvY9VtAO/xvpz0jaEA20ic4FgCN0cq2LoczzK7H+dEIeWZcWj
c52AzGsYJtWXu3coRn4VSh7OKSBtjKJcAgP5IpRazOf/Gx/iECejnaOeF6wkitGsWqYH0Mcmi1Up
grTwF02+4pUMmfGUXWFJYpLu/EQz7TbnmWmi8ByR+I5M9LdQ4tVODGvh7QIaF4cEICzxNZCSheZG
vUbZAbQU5hw0oFNly9Pv0OMTzn7ucldW5wMHbXRpvRunzfVHlA5ZDzlJIW+vrL7jeehoaTRIi2CZ
4Sw7Kj9I38Xbkf1l+EbTa7zhaz0GImk6zThB+5Q2XD276Ikn37gceM59naHHPjD2I255Vr96i4UP
b7hjdXXtXUsZinGxwvqDUNOJdM/wVL90yHsM856jPxKu3QpzWruQkeL936sqS6e0K7+mjBmzVhpx
X4g5FnPrSYOqGbHehx1Q+wCw9WGb0DYQZcCjh+YB+HmBWbaYnbLQJ4pdOmUFXCYwz728UISJRXA3
5au13SpX0hhrHc0f0hmpTUea29FHHjv9THAGwijIiyOKjIxgrP/Je6iW/ofPN6I77Ih4xb6O0ZAT
s1Pb8WsuDVL6FQGNiDToEBuEFc8EJkCcP5LInj4C2erVVvtSsN4whWCh8/0d1yLJauB7jIuok2Rd
vVZXQWPzgBO6r+pqWXezPoUFt84kcXejYjHd1di+5r2/jkSripU3AS4RTOSRIbwJTgu8+SygUApH
7paH0NoDSPbkyjkafQSDaJ03uCkET366FZN3R2HmXQLn4eBCggch4uX605QSYBCcv0GCDVVWH1vp
XNW7B3mGDLyBRKp/C4Y6gQMfFaD5VeIEfDo15R/x6+7OD9EUpiSJ61xHKesw9zMR5a3HL975eyD3
fBc/Qz3vld5IHaftw4jS+QGQHJTyH+w4UoYIlCPa1nMx5X08Jdyo8m4s7W+AYvLdzBWaJVX2KXIm
d1Yl8aTKUPLLYwgLhtsSeG1UW23ryS6cL5mHXskHv1x0Rcf/FDe/mcOi7bkQGBjqgo7xC3owVVfN
YFLowD8m2MlmuseJj4JuO+0e5oqEFAvzZ2CzbLukzTGDhruswrPPckil1MyWSfsYnG/QzTmz0Gby
O3Yr4s2Q1WuucuXekSfRxdXXTxy4+AKRWflpjR52R10E9klpYwVMyTIL6SWFEhpRTHy2FE4u1LUu
sO+E3dUc1tAgxTkrzCBMjmlVkLKG89ywfoDxUx2jNYM3gjQfW6HU3Zt1M+6KTMd1gmetONG05DK2
QWsaDQuieCJx12IX/AAIWytClKQXsrSgQ5k34v1CTUHr17QuGDjVYc7xwnnzvBLaZbohcVjrvvxt
RzGN1MeKrQM+r3TICaAfcesCSaRYHvjEfPKaM4beU6Pl3aoEGlDEuvLdXe9LX07za/TkqQcVmyTf
k1r77eU/jalR60Xe7XLsOz4e5vqS0uDKBRjN6pBLNQ13az5Gk8Fl3yZp37ZS0eTxvxwPA3Enf5M0
MfUTjnm1xQT0A1YvyPggyvSMSY/xIL6vBCKUHEYBmDuHQo1Ow1jgyDRU3ZsNhBPlwe7ON+FVHwie
PevWG1C8KWWPLHQoK508MLAXPVDVYCivnGcVH5t3V6s7Vf5yQugl+QBuYO3nLIZtEYDGsVKXLu1X
M/MZzgOr5yQtx98dg0HpaVcZx24Vk48cWY4gisRAH2Xfxo2OcB4K96mnj9POuWVvifahQ4E2NSPq
sawO1Qm2k1NihBUng4rI38H1ZE7On0gibm/gAS2v57S4eWG0EQZfMuiotO8p9m047NE3l2esgwtJ
uJTT/+m4UUfr2xIsGIvts5PhYXxbEfFHmumGVp5S2w13LZ0Qgy/TrpIRUGz2fcOq71CDsh0OKDWB
f8gzgUlx3aBw7jj3DwOOk7X059F8Asf7FGbIk468iOaXRI39h3gLPJJfiveG/BtSjrNLds7qc4ZP
VgfWUyxWtg6xOi3sTir8sUJaRQvXJErcId/fMRGn/MVcdj0bXmaiqW70CRYGuOKcwXy2S/xAMGUV
QiuHyZWqNcnUcKWgF0O3Tqc+KCLX+bxqBRnJMbwU3e7HIF5xVyZJbYSY3jN/iu2n8ulFGvKwTYVb
TLhu2aQcePZegCJjJyVSOiE8hMYjxr29FhUJiEyuAsHU9BgbmZSQE9Nf1lngaf5T8kOf/6/VZRiR
2sdMVVpqr5Z5zKFIqQDPiVo/yV/N7J5HBB1pMDy/JyfYB3CQExewyew/olrnRgRQHampi72v+icd
nGyVggOpKO1j0FteGQxNAATjFhtEDTOxwZBVl6xFnix2Ns8WbxmsBMqTmlGqpap2tpW8Cazg41Hq
KrYV2+a0VRkSJOUQR5apdpbIEG2Jp757huohUPwntqh3yBx8D3PtvgMp8CWKBYLUyFk7g/dy9p4T
zd0qXs7XF8D7OfBtVMrVVCq8cWBERZYmhBriAOZyNadVs+ajnHZ2xims9cMTGDsoK9jj8/AM2L9p
r6r/+Nb5H0hco10pPeyK5q+Ekvov/l1zjsnh3xSZgqSb7ycpeuXCQIiv5CRbRFaoo8B9JPH5/QxE
gRhGN/ceGj34V1+HYmtY7q74PZoAQOrX7DC4wtBVqjQ2EcMh19/+z3fFsRIuUwUCraLjeBm/D9a3
QFhFyDEdYGGcYAeLqT6Gu5ShuGh6E2EheHV8RXPoQPogBkDPcmTzSWeqsCjfmBqDHZDFwfz7okuo
bb5VUN5DX7MlI29vYbnthVrx6Ff88CYXKliHhLzd4qIS4Crk/yNPLVcvjZjCgtvToZsn3+FXcl28
eXzAu3Sc3ic8x/bXWB40BwA8/n8LywC46g1nB1Ju/03IimRz0shu7Dw9AkD2cxOp7xtXm7GtIIxE
ljGRMjBFvxvER8YPm8B3M0s4fxG9v19AWpXlEIhi/Qr550MoioV+T//bmTn6edfgvNH/bhsOpU3G
es34Grj5G3j9ACj9z61yCZhSzpK1PCDKvdLzQHptxSaAxsjlfS6xJ1PAo565TyqPMeZipj/4EJeS
yRNu9aTNFAJQUhK2onjvmpzTA0vpGqQYwJHekmEgFW5n3VhPzaPyh0p9nzcNG/Me9nVQzSCWaEgK
9gzCia1PdbYPWAG5rr8m5b44N6C8L+s9JYNlp9N08dfXtZc1nrcq3cUMwImbsL44ZLY77Go8UWOb
bK3n50PkN0xUxjKFbXIgH9icczu8KKqHk/UZQjwsR5Ss7Oabd60Vqhjb6aOFqv1l1kSHagYsOaMN
Px5UKnv400ep+E+Xvdjg6kVEx3zeeTTWWiHs/F+AgXcRXUvc8SOhKF+8rfu7dudkAb9dQV0gg+J/
dzuw1NOyXD5t18T+tbDtD3chleWREmIF54nrehTY5gVq70+uRsusH3YnYdk5eTlzYPeIyK2/+hkl
WHeZ6NzNGbUs2ydK/B7wGKj63sKurSjvtmEByjo6plcBtalVBVn9hRtBfjdNkTqR5gRBEtmixcPw
LG1GJtugLewf9BB0MieLpay5QeuKv45U6zU6tNfrXVPQPQxfON6YFArn7dKTYKuSkbmj3vD59Egs
bIw28si1azUqiXVmAGjKzMg6D0KuYQa9X5KAW24c5ND1KLxn6GUVDP9WS+3R8d14RNlcQLvOu+Ez
EOyMwvE8HMQpgErMA4dMBV0mDsbxCAIFLkn2S7A7c75Z7MH0ObRpuZGaI41XLpXG6kvAxBDp1dRc
YMlw+nZ6lQf+EMbqNJ1abyNBhvMU1F7RLfgdkfH8XHspkXmju1HueR854FTFvW2Ty7VqzI+gkYLA
OuZsKAOk7vHWbN1jCWqey7J2//xncN5AFcZp6lCR1n+LE2ASa/ei+oAu+cZJCN9E0wZ0OFFJwnI0
kMTlaOdISFpotA+J93RSYbrMQif+KwSARmYC+cwjWyJqNaKXbJfDxzc6Xre8NQGXlCx36zDAgmP3
3Nc1URgaG62pW1r/Kjrjo2itGdqRN3fuYvpoV3fU3Sm8AYLAs8GpbVAcUGWZTmX76zZrQXyVs/NP
tyhbzrT1VyttMshN23KC4q/9An/t9jqyLTofzyDz1Bxojk5VGcCldMvLot2KR7WKnb041GfNtk/C
l9A6mw4hXIy53S3ZdYARAlorb6jwr0G3Uo+MSqUgvNh3jwV9Lhy3S/CVnlqWgWvsJUKBI8//UL51
Bhs3AKJ9QLaN8FFxEUTkoIiDF1qC3PXtTn4teNOMnVsb02oAaC9wX4HUJG1eqmtfTUWg1j9jtOdx
Hr18mX9rNiNeKLL1kqh6LuHRD1jB/NpoYZIRWX20XtyZdXc1rjnFMWVzgohKIAnl7l5bYZMj/1Vi
cE3jTZeUiB+Qf7o0OaHux1ziTVLxceEIex1bER+xgpFXk0gVl5KPNRFZ8rW8gOxj2ggF4LuOfPP4
oqvpkTUwGRsqnZSDLMbUdyrJ4qe1GXDe3l/Tu41iYbrnTj93hQCIFY21kNIyogzTIrJBq37ztS8R
kqi0/bkAqltXWG5qEype25e4csNGiCg2G8tiX9bc7Gqzgyka/VzscQ5J9uDp/6CHvzTrP+vw5poh
bUuaom+YD8UwpwD49XrqoHZ28I8M/wuANl3rKo5PYV9b0+XQ/A4jOYeQ/F/nKMj3lUngZY0fMl+u
M/ptDS0Kgi8vvbr9ydPvqCmCJ1E+XO+tmnZP8LOORBQvsqGmidcn4PLflykYxcZ7Y80oj/CE2XtJ
o66uE3cB0RA6yLXTbBCG9IAek1954dgN0Nmaie0zCD5YixmKODhKRpedCV5zR74qOBcNyrhdrSdK
ZLYsplq+K0nPHiq0Ka8e4AX5jv9YAlxhMp0j0iLRM7v8xfpVxLG2Ir4JoxHU+TNHLgpkzpd1nHHi
MG4MCXhOaU5yDsDmW7ADDTbjRa40riFKFJZhq7DoY2eU2UTcuxRkXJHgQ4/0C1wPZLA9dBw/EN8u
cTdMGWIjzl+HdNeiLw6RULiisI2HHSo0rOiiPIrRoklmmC5j/KLsCD8HZk6q2ruq92mf0ATgTn46
g8sY/ig6Gw/o8lKm23qEqqAfittvON50jtsU9NCVP3CZgghFVJC0g15fT+pq62bmadb1TguNNYsp
WQD17dU4JA1opruK5LBCxR4ZhelSIhUd05mBMRaJNHsWG7JP1UZun9rDPAt6onNNU6s6THT9Okc2
BihedfR4JDDL5E6p9PK5+4EycJ8dP3SqFuKY5JJUgLwpROzIsPDBLv7rgMgGGDfHatdAoiNBgl20
fmKqb9AVWDSbZC8YDI5iA0vCkKN8onoApPRqxxm+cWW31/LEwac9NQXUjV9jmhVHd95WzEA7bxGA
6c/6fY3THcTqKWAbc63HAzN+KzKjP18fvqY6h9llrsJWSd2ClJutJQJQASpj1l5Q/0WRL79xH67v
3bj73tDFlAAe1M5bLNKirwFvyrKfZBip602gIFUhSfxI+Q/1loxCrHB1V7d38X0OYE4jv5jCzlo2
uLa9CD5ADynVpznfUk/aEEyEGAWsU1bE2M73OuMtKkEhZOKsaohOqcwJuKQamshweC0JDJeNQeiK
IUql6RjQ5S3D6dIW7Z3NhOcI22PcvviXIt2C5J4xjdaJzm39yXyu5rxTnpYBjsKEqhZ1d/O++85L
dznxcn/aqdfrXzeb0bw9cyo1j6gZ0a4Him8Kd6BvHDGOMcsMH0w5xg7pVwn5Nop/kKkToYrgh7UW
6zr0mZ+Ho1avoC8vQRf4FXMTC6OTPkEbRIpjFg9hh0N0sJwTaagpLOAgrqzAyb5aor/IFsVd9/y0
YwyYQukL3/k7Upwnfj/+IsJxyRb51hViVORW27snEiizaB93+FcxtzW27Yq5tqRevcIWJuftuv5F
d2OC1LM1u+4YQwpoclDjxy72VXWRrsj/Ioyp0xy1sV0dSang38mK/fK7AZKkTvjUAgWvjKDynLHN
iX//wws43/l19fRR1gwTRoPR2BohDrE6i89ZYl7teEpILApMsn4/cG8bwOLvXhAhDnEVt9yvJaDU
qfjF+6el9LKChoQvkykYTMZm2SoMiyaMU1Yzy0EDkeqa/q176O0QOuz5wXKG/Q1nlj5hJIl35545
RYG2ovdAdr9QrDvzFUX0mZdCKjfS7gvXGnFg8rgUqCVASR+Ag1AwtGAbdkCoY/Dss5oWXgAGZvDH
LCDHn7/EUfp5b0ifhF3h8hY3weL/CkDhupsMuf2dib+LfI8ex7CfgpVspXpzCx3Q4Tm63VmqcyFf
HfZGjPfUaE0+EGdePdeUDxKu3osfMyMFieoL+AWi2WaQ03icBfzG/hKGiNEhBWNAIhft786n4JiX
I6CH/BFE0fQq2uo1RNaq8s1yduAy7J70Wl/HFNdBLheLM6EqhSFJfd20I3WZ/0xP+2ZG5sRDmsm0
/tW5JjaegmcGNzJ31K8TBRGfatLH9cYjFNxPuFCjIWcPHsfsT9ftkTfL2whsH40zGhIlLjByqDwj
y665TTMcqq/gVPdn8C9XXjG9GivI7K4XXhxztaMEicw5NmvQJtsMPxuQ98OTRU7JCa04wafdnu8q
/lvoE+iCvE5/wZwXhToNQF43IAF8xlyHzfPYPpUOKc9kbpEe8sm5mUe+FHz/EtEO/ZUqU8Xw3+TQ
vo9aMNMg5fWbnR/HbW35FJsvsOZ69zaitqLhU8wgTXx8XHN8EFkLPXGQ5WBA4nB2FFEbqlQVwsf6
SJljcC4qQel0gzjrXovWoHvAdTln8fhvx9OBuV/9I5nHL1j2lI8pb3EHAsTAa7j8qPfhl6OWsCwf
FntcKunuP9XLkQSamrkDlS7XpbaEHbuU0sL3hcYVWsyinrAbjdx4qr2XeS+0nDGZgnq2ibin957P
32/537g=
`protect end_protected
