-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
EIwanltF+Fj+8yUCh4uasy45a2lkCZdSRfdC0Ua29tkU5rO0HI2YJVpQrGQvFfE3
/pJ1m8B//UpqFs0jse8PJWDQIiHdLiO9yef5lndAvf1yes5B9OX2uRzMEsZTrEBX
CCyAmqs9pvVNINWCltZnCP0sruHAIJSy5yxoXsQYSLDWjy3YC8H9Bw==
--pragma protect end_key_block
--pragma protect digest_block
JjVNlEWsGR00jMtqMzaK9iOeRKQ=
--pragma protect end_digest_block
--pragma protect data_block
NxZSI30D7mq1zSoh3n2H0ZqDscUkymq0GF5xxqJbDTlMvry/iCw+lEUzD1g8QLqO
9QYnrmlzUu+wYoB3M4hBapWuoM2D7/JwxJNYX48XH34F/zhdgHQ+svNfxKEcS9E/
p+RRXc8WpOudSFbIE4CzkCsgDg6tXNq7YJcrSUcRIB2EVMBcsHgv4qg9JpQIKHvs
/ZeuVULi2XHYlDTTfDQc2GP+7P+FAVMV1e2udHNCMzx76Iih7nr09vZLwpOkKYsh
JeovteJulsugMZ1TZf2qEdAYOJUWG1NBdyfcEz6koUHdmJEh0VXjnOKkJhhhGmfY
XKtyXC5aImZMJffKTcVr7b0ylWfRi2z02KtXzMRl1/ZuU9qJgj1JSTCgA13akpJu
7SW5dAoPjy60rGYipFjp72W8FEhYAceXIzlkgZ5K1Fj2XNP5xrrF0BDayPiys2QY
hBXvotuOEOwb4ps6AUfGyDyEpNdxUHi1nMCI9qESfR3M14UEHAT/ECbwUpNNJ0yA
onB1lHOTD2S1UMEp+brTn8oUb5MCknXRv3SO4vhyq3U77s8nvPY3C4P7/ffL1jDa
4BUMQPA57tO+XVzzC5YNnKoXA6YtXzParRiDZhrkvvc3QxSVBVcRdkIOx9LuWk/M
V9tAKweBtujfh8eNbnF1rJcCfrjEsWwFqsr3bQBWDM74yyO/rkdGbIbGwmWTt6KY
0JsTYJMbSlT/XNg4a9/tFYfBt7Ptt4nQ9bxE+tu+8haXkCJMt937fBwql/mtxHGM
ZF3O8tuWGtAzEZwOMchnAreE8/lFelOaivhb5va0cc3KHtxBni0rX192bJQ2pEWb
R85ohbgDBR1HfpNHuQwRszeE6O0MltttjebGldW+hyEKmj7aSv7bcECE0fb8PI6I
WEuvKI64bOuj9SRgAEReJxXhsWqLuhTIV1T1ywMFhtdQLj6kI1nXF+eptYC+ykkx
BdUvBWNExtHDLYJBTz0q5Hef8uQ6ovTI1eBsaOc4L7ax9tF5FtR0cTazLydOMce0
bw0sHFGmGl1Un/hdHZo64M7dPXSNGjX0nrnpmfhrZnBWwTvr5OQXpvyq3INHT3Il
16dSzMK8IAjSoDswOJ3CDLi4dFk+GCji3QzaFwTO4cejNAzlTHtOsTDpnConkZEu
MVq0VafdYqC603E3fW1ReGBPhB8zFDh3iBdMVmyG/tuoQkhfcbbZN1qtX0StXZk8
ciNCCZBqFFqFkL7qXEojtTU8zuWN8PlLe4jKChcsgG49PBtaw7T1cakIIrsNGxeD
dWVpZbqq38nk7i1jpj+L6sv8zIPhBwXYDkt9Ytds9ccb0HKTz98PaBu/jDNSoCm9
hNZeorx3lEYzrdPjcBzTKuZBajgLKGg/XAUou4YyWzVLNgWTTFZ1mUt5EieMa7jg
sfyuYq00S37lgt04o2CbyoRY9R/zAtv75xU4FHD+RZQDoqw0pnr8ZZpUD8vIQvXt
hxzJs39i0DDn+GENseVXvXTpny5pSTk7Qkou2LTnrRF1QoeT6k24DgVKSxeh9l7G
3MwvDEmY674CvPFUBmzGj0T1iYaqXpwHB6gLT1ewq1s5HO2Blh8W8AqcnmUVX6cU
xVg/HhP65AhVTAjuwFl1NbrQTzFQi+Isb6bt9ukCWlS/bQMruf5tqd7Xti7oQCvV
gkj8SmjIBaf7QakQmg5mYtZOnYUdTKZxSYViJOtlrBIuKFscQywm5YJV4QLw9nT/
UKGgTvOKTaEKTCEYmp3DlOpVENXu8i9PLN91zGwx0G6FBQ2GKVudbH1gtCR5VQMX
UNAwTwuq5sjTYsUD5+bFODYgkRwDdQUGrdgMPcl7lS7nAP34JGaSQ/vj/wC7QlNV
2q8dXY+PUYqlvnYA3HWiuap/B65maEwQQGShezy/347ySNiZtJXzYGLRXJoXh9xx
PjEKqaI07NNzHBp1VDnOPObVIxT3tSSWBmHX6y2E85t3M2lC0/zbUKXZNEJFjQxF
nzGZaGcOisVoR2QTfagscB9vFuj5fMRYfB5EzLlGnEV8KFfHfXhtpl9mauwHWk1s
B/NaBAEsKdC8YFhTscM/ZK/hTd66nmqkV7gf7cAIL7xmWrqiCiVMdo+uGXHkGBts
Cb18sSXtHGyo6YIuR7UBCzgmuKD2RrzTIFIdlWHYmKpU2oRFe2Glf89UKOh4BhsI
HzQolPdb71bzoZT1EUEFEpNgGT1ZId+x8sjl1ZCNYO/xl+Q4jIUGg95MCN2FduKv
Dw6DLnroZ+qH9AlNUYCHTCAZ4kHsfLVDbhazXP5LDsdzt7yTdzfp8eg7MAZKvh8H
tTUCybqb9XmIjGILp4kVfHRH2g5cQGPHaDOQIrc+t8+IoQWU5/nSTk+Q2888haUx
3tGOQb3PF+9muzRcsHnsQJU4lo8wZzQrusgyXTABKbkOs5oOHSvJgCSm6XtplNu3
K5bLcH1ydmfrgu64y3zRH3NY23q+H4ymBFs2RipiLO9RvETYZN79/11ZbJkukULz
XVsyK2BfxphrqfFrFAlOg6YEb7E08fAVzy8NBaU1nN/UZfISK37cWXtLAatysgrP
PHWnrlyZFbJ3tiY8gOM1cIUJN3DsC3CnpoQH6axHDMwYY05v7qefk5L+eg03meCx
MFy7n4I70onJFl8EhRGN8HFOMixQT8rR+HYU1M7ubnfLbsdsMZrZ07IMAYEhCH44
lGKGDNpkce4deq4/Xkj4DSDooL/qauSBJ/IqFCb98PlAyVD5F2Q7dGyMg82bPH5k
756kb7GTLJkkMUCqIWwZPU79QwmvpO+pGlSsAaPhOmom0lrCrHJXoSSL0Dc5jLyB
Z/0/3kL2WMZE6VTc39fq/8KtrIXKuHZ1dX8LvNBchAr2PENZaxncq/z6rdoYwTfP
MHO3u6BZx4v6N1Y8CXLgLu8jiNp2Sosid0nrZAuU4uEcetnIiTW9Pf45Vkur8gt9
rKnk9m1agHzoxyas7gMkJTJgaKMANiRXBe6OcxzxoXj4fAvefKlj6guEXsSjK3Br
q8+q7j5kMHf7xNKnNFXBdUwSL3uZm5V9kw8Hhfo/Uh/+jT1N8V8oUjCMu+05WUaG
NS+dnAusy/wvs4s+ZdMcX8EwElkTQnayXRUN2D294HDzAiR6FDWFUEllFxWNBpFd
+Q15GaNjYhkR2FMU2fTr1sX6E0z+icDyT3Q7WEPNfiUiRf1FTwP8N1JdL2v/j3ln
DEwVRpQSAB9/Eus1wUQblIBNrZCsiih6Z4aYw7RD4htTlWMmUI/hM8Qe3fCc/Oo5
Mrely6t7bm8TAeOl+Jjs5Wsnb1WMfbyjIEgeglPFRXevGwylgRK8PMbLHcJIgeYx
vDc39/kuz1eJlASF8HLaFfrjSxjJcBZkcLpw6p12lNFjNx5bqmUPA/tPSEwHsCXv
ypbkORUIHD5AmvCwz9GLDjfvU5hwGNHgxKD0WTgiP8GsfW8IkBPDHd+vqusZkZlR
7pg8G/W3qZ+lTEMNZe3i+frpVd5vZKkVpOWelRdeDYfVdlXDYKFngvmkvfHcXD7a
hsgoNbvmx8yibQl7iHWuGWzSDEXnpliSibT5O2y6i5aSK768ucaytLAOMetiC+To
mCsXOfOc/2r7rczTbX2kFgmBgX35dvcskq1PFTWg15ME8bpV1yFEZt7Ne0evs+XR
uH9UDX/ZSbP6ucpGuCqxerTRIilahdp0DAwtafHaDJd3xfAbYawpim9X/dDaOpJf
c8b6BpZxJLXM+lJoPyTAgl1g696nFDmKzd6dIlEPvZQnO4P+jjoeML6AtRv2YFyT
7hcQuscLlmDOxVZNwW7SdxIC3qxp4/x16JAayJKc8rPY89ve2a0a4XgPjHcQjvDt
MJTnQKMDzukUEu9/GBtEfEcSPn/x7E49SQQatYSXsVQSb8UmQ2MQdaesu8PsR5tf
oD/Jn13oen8CzdrP0w8/TIgsIlimlVCeqnq2muglm9w+HDTYKjbEYOi0NTeZWlhV
IfUGhGdhYen7sOpAcTrs9vc3984BM+RxapXdtFo3CB3/Sw7I3rYeaZc+YD9Ji2JV
/flXBQh8LbCMoIOvQq7f6JTlb7i8SZvTZrgJZ+SelOIJMWhyRoOniMiKbZ0qWTBi
/N3PeOE65e1AdPB4ptYzSJxK2ahmLJnnpzoD/EibUOku05uyMQl6r+PEFATq41h/
9LR6raSGcmiSbCLKXzPdZixkBg5J8Tr6N5J0Ldmwft4oQVRtHyYIeZC2LKp3R3/u
ZEQvBLo9zENWAvaUAKU3gE9DSOmeCrwX62o2QOJlQJxPwm338ZhqM5CfyZs874dt
CN0XM/8zxMWjvwpsJbkmIyal88PPwodZtAB22qU2Ck9mGjZqYO7walBSpoHvvUfB
ZIBv8VmZDnFfc2m78EuW2y806z4mPNOLKN0H+9WpIJbd1DEhIlmnrozlbK37n2jC
Na7iSONS3kZlYkwnuVxoFmKV4i9U/Z1XxtPgG6VI1VLdR5AYpi2X0NherqcO4ux7
mOXoyQNubMYcnMZrUn+yiiN1X9Vs36lG1NNUQ0rjU/aWJFY+onpJnng1S8A9UMv7
gQVPjaXncSbcLu/BvtFGbd/9idaD/Ei7R+EraW3kkeSOYHbCktmkIjijupr64ODA
hGtpkMlYTVv/pSt+pDfKvpjiw+0DFqdt6Z8Zo3rxVBDPslcxrJf/Cx04lCMKgkFA
4E44AHHAoF1DrR28mj90m1q3vE6JQB7sHIy45LlvFqazeDo2GwDtHy96+NKrFUJ4
H2XQvVzo7kjmkkYzTxEh9fG81c/oVBF9h3jaJpoY+6SuRvoDix1YOh90tYhtpUuR
7Tp6L5Ja9kB4uMz6CDlIMcvTtuvFgQAIwPWqtgJQ6pty22jsm7b4bwVgHku/0FK5
k+DrP7hEtcp/1XPfs0EBH12WcLY30ivRMUepbBRNi1Z9PWd7hzS48FRr5jWMejSQ
fOf13reTlif/Bz/0Va+ZXMXCOnCTqt8rWUuXGl1nkRvMTXHcuihLLSHarEH1JyCf
NXp1M+orMMXSXRH8O5wZMJs4ihMLxMko05A2NONqXMMQrQ8BKNUVO4Bo9+UHauK3
L/wvKRekXdYR5475KeYDUMQINWyEp2Y2pMTM1b7RcaAg6AN3t5djzdQgwF3qNcOW
MVz/M+Rzss/c6PbOxdsqHTTbIYrl24Zd5GHdJz8chPwecp9R/SC4eRGN23jrdC5W
kocv+JRHNeZMI6p4wLTabfjHaDloJMtRaakW82bjKPBN/VTipwURMvbV1sCNVDoE
yJdOH1Kw9ke83msfpUXY9x8XqeppZZ3mZXzKhbWrkIxGGrmQQ7FBQ7Bni1FT+i0l
TMfzVOwDxYPqdId51YxcwDwEPMJVoralayC8GmnjK90GVkrs582zxCky/buL4CIk
9hOEfEEKXYelozfmvClJctPbn8nxn72TnlpN73Y6EeYn4ltpEZ75p0/aA8YkLnrg
vBWQmi9hEv7S7pdtNNQ9cG4uvTWpTmSws7rO+ikAuebxKxRkbzFQocgCaiQMKrhZ
lfOyWwCAlpsMk7xhFKW7T/rzlMk4bRuNwE7cCMDboOMMuWK5IzrIxS8M7rTYcwdY
JRUUHOjUZdwa3qT6co1pejiOZ7BwXfU1SmcWrwewQ2UmMhObZwg3roKBoOw2ZtfA
ifIdQreiGDKZIl6OHuloFEhpPNSJIC5tYOvPxRukW7DzSqwTg1L8xGlK8FBE/bJT
yqwXD8vKvhN6F7kEpinoW/yns71cbKhOQplGWqnBZEymRO9Jh+0vrDCfgRb1EwKx
oBdG2IA2JkOS2Vkypj+8F62H8Gk7VVEk7iFXEXasOMgtbMfbJVIZqiw9ibVotNGH
dic3A6vZ5tqdrWPcRI7CUgfr+QxEBoXlPqvQIWFn1Gm7r4RVISZBUMFBqzwwiAcc
+mmzyqsjZRs+3k77+48FqEQLupPpU5lZ+ceA5bwEr3gG0l118PwU0hEmaxT+up+T
66H6N80xPqUt2xePf6KMe0INWU4G5OJnosa1S/tZISfEWVGoD+cNFy2YjdXpiVBg
xb5FxN6WLJsxZpLviCsQbr0mpF3jzBPS9KKXxe+IzenI6iRTlKe25N91ns8mfoFl
+4sRdMqwuG96zLgDjO7vQfplIb7wXHJ9t85dDvE0x/WUC6XpByejgeElPyq7YTm5
3NZ9TnKu2buc6Vw6fVDOpdJIZGraEWLtfL0Zlb6BKLGVFLBVM8s0wZ4vqwRGeTfx
lgPPPXjZqCzqqG1CYFXYo9vgGI+YW1X8W9RLbV8QTq0AnLrTU2EHus3ZbBuAyRII
WaN8CiBvRniuvFsKPl5teu3Ulre2SjUu08AF/Bec6OATyLz1VQTHKoPnYzBycm7c
CMY7czoegtW42Qz2+LLZsvk8eUr26JDqbehhKd+6NZ8jTllsK80XU8C9IjeCr5iJ
iZOCHPfr1r52GvqgvMnSSBM0rrNIRust90Zm0fhXSr136De0sHHgUydsssOqMm7o
LiXERZwCp8Z7LWfmUL0VUTe9ode0c/JtuuBK2VjgqWL27cxh/ixr9sdd4eXW8LwB
C+EQcx/EXCyg34UJ/vVeTsJpICsxYmYaB5UKfbTxvWhdQJXXHPJVuzZWUt1WbrPl
bT+gTI+SB96kGDgYUmNJpgE8b3mCDw1zHUOQtTJyXR+jpr8e0LAuC+Z3v56gNoBP
Gu/FO7aj30PyYqksTqdH7AVyDN1wYhLDZgQ6piJrqJX5m/dwZzuttJMENuzZF8bo
xL6XVdY9CbYKHM+UhYf5DTKFbH5qSMp8RVAdT4VfvXzU8qKvHTzI0iNSUrPW0TVg
Z0Teg5OxB6uSb9MZUy4t23ojST3T2jd3X6bog54EFrADqJQZ8qd1YP015laSbfSG
HcwvbQCJfqQMDtzB335HIpplnTot38HjOtl+r3CjRMg5L4xuMFzH6RQH28azsud5
3ea0sQQwZFp5yZh1VNMuAmHHcJtPcfzirU1ueqsaYJJAliH6uRdT1dlxjIatohle
bzy5vGxU9omCsRBjbFhWCdsmkMP14F6OTzvEoTDvJRINA2NeX7hiDU9KGafAkV+8
3EZ8nipYWdlAkhK15WYpGd6B+07gU9MoPMnuGTmgIqNORN/daCS+JiltgRfdN5D1
BIL2UofCLmGsRCUNPwIu9Xou2NBwmANR13v8FfE4kpEa7mdajKaJlL6+9wVa9asp
a6PxlIlF4X8dLMd/VwJ0/v+zEXkYqmIPvnmEqSbEac/IV/3lqJ4lkcJpmefBT/tN
rxCEycc+RL16kNfiXrDSeR8e9f6baiD5CNoKCw6WFR4MVJQ5zGq5ht4GWVmG2kNf
wA7ta6KEZ4hQHfU7/nFkNwsRR1mvsJJCaUsBFkqym6Tp4biJIhSo77bMtRYM9d2D
E80fQbz2ij4QCzWMym4ZC627nDcV5Cgb02NqeYoxdlwcWcuNuLrIYbwJBqCVqGO2
J4JPf7tUn4CdWntAIHSDV3/hwaKOZuW1cF60FL2yAGNbt/vAWxLSutw2XClZQCet
c+Q6agrXD6JosxhDP5qMMWON9wS578ntBetrndPsHc4FVZnIMk5P1i9amfHCQQfc
LDVBStk7se9uo6CMGx3F8s2/NzY5aeFc6R/0GYeMhZUBCmAFcm1ylmice9vv3iDr
qpjm6hegbPtKGcsMjKNu3ADs6ec3NoWesmLKCZ3JvMSoB4Uiyb2/828NAw4+NMtN
OJVmhw4LCUZ21k5qlHYR9v49p84/neo+P0yKJas1vvb+MCStM5hm+DQB93YPBxsR
44pUxlzwXBKZcmtejeZWRLbYibtRXDzLGE1C52xk0V465I54aJZdGzfQHkqnxiKu
PcdfafLx0l3eFAVHRorF1vKs9cN+MY90lg/9+WwrgIv3xFFTixKRfjCtAXZoVZXZ
Vvtxmd0THKKSQ2PNwfQGBHZXdlriMJEHzZk1iWwIj6CONWf8KS6aactgYvRC3KRr
dLsSfgNeqSyreTSMqD+FBAhCw22i9avbMyiQpUecP7INZQeaMJo3MJxUrxe4dpXZ
a6GgyVP78KeaUwWQEp9M3mXL4mPgoZ0Ptha9GB5f7mNj5W2WiDN5PCAxwDp1sMMH
jH+Y5GyW56zehCwbCVrDL7nSmXzK623LHVCjKK4qAwubU7bPS2cRlbG8QOZtgkO+
GejL5C5xVUO2B02+oqxM+r8Ekl/RveOQiBInCxi7lWgfQzLLxlNYLzIGeMQ90fLo
Xd7zZLIuaaSXlJNHpybP2iqGlFnF5X5JOmrF0j5SfYCQDv1HHCO3NvcYtNuZfIEP
AAy+5lcoITxjEo0o+wjr61MsMsVz0Fu4TRYxKTPbnVEL1E59mQ/R1lKdVRhbPr62
B+zLc4k4YeNseIAJYiTo9iB4lUdMDAHoU9VDrdvrzP5lMxSamMu4rJ2+XD2ke1Qj
p9c4Cmsix5z7BMaLAmAEYq13HBS+VPHlV8isvjEYlCzmHlRTFUODcn84uNFUF2bE
4hl6HVANdNUvvC1MDNoUaxR0LJi+pPr7GocHSbzZSaE9WiwatTB/FNA/qtCUsxNW
y4O2gWD4AR4+QMyEVYKNzvdVRooWQCdKl+jEd9mJHVPU+bOO1Cb2h3H9ReO+RA8x
NBe8peTukxdjzScxJTwQRgmPPOuJRoWTMt1XniSDJtvEGHejlkWICItbrwG9bBau
T+mY+uyEJr+WNDmqbIdWz7whv83zhN5m7FNB97577QgNpTjvhtCkvms0IvbdRiGK
QTaoAZTXYxqN6cPgqzJqnJiYvEFcDhaI5Tgd2ZxL2DpzkNjnOhvuWSpp1p+4zJfW
pFqd0TKB5YxUEWD4UcapubI8l4daMPkH35TbgroMJUzUz7ouCbG1CFUoOULe2st8
kwzTzsBHIvb/nVv7MYkIH4qMfMGMiXSnvuDMgDprzGH0TQRmCzXQNblu/wUtZpBI
A1hsdM1ufryUNulgd9h0vrNDuVvFkc+aDbkHCmLD7mMxXvxz/wUyZoeNCnweYu3n
D2UjePydz7bEJyOr3BNEcKJno33aVJXCfJ9UvgWMYhi5f31H+HwzyKxDLW4OhHLb
Z1RYu/UfKIRwhs41i+Az67nECbsyvfsB+McThloJ7T5A0nQKLx+cSFCz3EeVmgFC
D0DQJdz5/w36msjqwTTRDuMlTjQXxJemKLd0yMa+ts5UsVK7xe0/6x1eBoPC+54h
IfYRInigiJywx9Dq2h0faiPGXcWuJeonsiIyByypd9MQDZiOA7QucOhmQZrTclef
7xMEYCAqJ6y3JE5pAnJsWJh+GdTdcSst5xKwMqBnQ34wM29RDCokrY2nkkfCToKj
l5DPDcTrKWnyR01fGAYvdTrrw6Vw1b7apYf/YNyAMY9WLPZtmGnWcBZ2kwd2Z1MG
M5GgpCUsLOnXG7bjjYFZBmUTcWz38IJ3V+1G1bXaNBW6b/YSu8BhElSdsD2Lbf97
0ULNHcwLwDocT+8bN07Up3Tn2BLDkDdxSEaQmtv6MQr4nUBlxnlpu0zOZ3rPWssq
kpzWpCMMGNRgQez0NVlsmqz89ve3Tmu6Clotrs8+3aHeOO5w8w7k4MIKR/NtfYLH
AzdHxBvBs+U1eK78A0xyczVqUEmc7a4RauzCyMkFNQPCEGqBg4tuSnDCDapPOZUz
EWxpcr3ljjXQAAE+hSfohbxnA2pL1pX46Dt2OCcjAdkg48XUzUq0Po1fOIsz+22B
x6z8QO1Vb0cKBgprd9SV0tyz7SzoEPL7AneeF3P/7v5EkEJAfsaTXDS0LwUQYvhv
6wyeUDu9MiqJ2V1F8WgY2dSSMP9jV2ZhLTQTyKrckiXMjjBBzFvBJGxXDHZySh60
fSpdNttzII6QPRK30FKiWsM2mImkgS+LOZS1HO0mxow1zmQEzX+pkeHpwkYvfGVJ
cWoipUbeYds30/abwPUyB3zRmuSbwvPDuj/T+wvUx4CBqVnIwK5LPVEiB46SsxFP
3qglURuUPogUgGQ9syfNKf8leJLGHvQIoU8E9BdE0RWjY3+mxXUxFPGSTuCgWvlB
ihPCEiVzSRM2pYgoGd95T0zHA2BacRpvfg/vsTH8eQKZRdurnR3SWKIJB3Udj8nK
K9rOKO+ke5h4XzDSQr/361GA9GQXydwm0B6XYqjtQO7BE7d1nmqWShIuoZ1r5owa
bAFNKTegd/VWuKY8ML2/xzhQwwXbo7cfX9LHPwQ8OHJA2B0px16MZPPhZIXFhgey
A2+s1S+Ad9oK8seZSUDeRwiX31pyQfQfEt3/wVwSS32GNZc4L3kSm60WifRVLqtW
gQ8NKCNqv0FefAn8vYMrkDnXMV+W3X8IDP4vgl2oW8WUIoKW1SO3WgORs1d1fJYP
7AyOLFBFwGN9pfG0gXENnlckt/xhDO3WQz0V+VYSyXR0z/jixxar15Wp35fmm+fe
AuixxVdsdPgPEsGG8DlbV7I787tuA+cTYPkgYK2ymqP7qxrt7Sh/PZhX55dAh/WY
mkO29jxP3Xuh3H63Zj+JnZxO+vdIqJ3XBT0l+JoFTe6P/B3tuv2WufyXrgdVPUiX
Ey3kE6gwb6oJ8toU4HHXRtxk1hLWllGbKTNU1SWKsg9FOEN6OLFOWfJ5TgCypK//
Lq8fNElna+fmPViXYblqFpqmtetdkUFuxiv7Kb/3gNP1QG81pU456fINBwjhcuIg
yXm3rQFenKf/1KE5oV2g0ROIYZT3EMJu+1FK6C5jlP/hzZK0qL4+lt6h5tu3qYrv
TkYhHbGQzCiJv8mxjPHk9PIgaOZ1/tt/IrQ0Yo+qbfHGpOYRll6sIVmtdt5hziEj
LYuA8mMuMn9faVkXu6VKsAiH55hFVb29W473JrgYUxzg+Kl5aH4IuSRxCjQ+O0bM
u43IDkvLkWCYueD1c9uSZc5x/VpXnZohhPCJUgWugUxh9G56fTpxRioTJg/5eU32
oaKmpmW3VSOvflC720SDaDjSPaZHXr5NjCQwNbG+gH8bsKS41GeeuqE7D6ndaexT
b8TgiwXvXGPTrS7XOm7u8yGcY2XstBnbxZV3VniZQEpqC7ZKlSzTLObOdHvDyn9D
Sg9WqKd2AZnPD9QVO4Fa/u7JzmOtImj99pzyHzWY5LHl+2b96E7Qdth85h99x6T9
eFVp+eEXyH6WFZRMztFkllwn2Iv5PoMeYg1Rb3umYaS1eN37UK4JohdqGKjLUvGL
cNV4i2n7xBatexbNPfRVDpy5C1tuzU6TgTPuzD/K8u5BoMQui+NuG1qf101Uiy10
cnwDlIv3GdGR4gwJJrVtUkAwNnYK/sdS3zeoivq1JRs2Xd2b6RdvsNYnpnl/YcRz
y8kQcwiXLBwxU4QY8zCM/ehuqBkCgRfXnt6LSCdmGU8xpVZ9rXj5ImOlI3rjjCn5
uHQeJt+eoySXFf1va9F1sVNCqa9MKsjrGhiC/aCWjnWCtK/HA2lvCVB4IdMvcM7h
8GvS8YSSejTDmwIF5FU0tdn+BBH4QOsOeRlfN9N5rThRZlerCL+u0Yu7aXjOTng5
ATXugafz7sg8Jg4CAVX3Db95qsQjOLCdXTqEwJuj+GSw4m2Bc89m3gdRl4+DReq7
7rZrTXIvSypL2DlwOFeOOd02xYg45/cR1kY0MRKLuQOtIF664G1oJHsYWvCu2cYy
TBiylFpKXZ0skmGccN4X5zKMnwMs99C8lz6ouj92V8CCkrAg+Qzb+gL+Z9wQkQUA
T/B77cIE7+RgOJDtwF1N/FQtvMeh8Y3zJQbxxmPKTRlff94/5G+sY9Q/7d7WcSvJ
K7TQaRhuRct/BKi+zDqcAEe7ApKgTXYjHMIeVjBlS42jTeuFVJvBOvI0kSBjfd2h
u6Vb/OgGhIFiREuv6hGxv4SJ2ECsIx1yLEC2vrk305+EiD0NyJR7wT4lniTzFT8Z
2mp5dEXhaLhCG8XhibQnxYH9Y78V3uLWeCx9cskX6iDnnvzJDXKRY3/eUrxwSKmF
lhYj+Xi0xqKv9z1BeguhvXtRwJJpqCLfmMonnHmcEfK/OyI3HkyqIf1RolAcA1lB
MSBUjkHHm/sL+6/Mrt99lF4dimKgj4dmM33qsxLLCHbed5JjJ9HkVX8Uq43RzvlM
cLuHXYkNzOf/47Qf81D0uX/2aERWTOSlRcTZmf4/P0dRqZMoMZtkwlxgNxFRm1AF
VDVX3uBweO9VlWK1jDT/HQjePgvAZFsCbY3phVedl5a+1y19CtGlOxjKjUoiGG0q
eHqTcXB2ZznTmS3gWNa+BFIg5t1I+orytAPmEXwyqoBkYuwemMia5bsy100fDztF
C+CIB0Yy3nlraFocEb0tCKO7DQV11kllI/d+uIT0QyuTtnBqrx/6pvfB6GZW9UKh
9RKKDpRaLXx08Qbe+12inKLeQTB0/k3Y9Q0AeCG6Eq1JD9EYmsQREPLjmf3CjyqO
ILumlBTORJVCIfD7wyGNGtUVS+J0x3ZQhK9Q8naWEbueDWw/fNMEtW0hU7mcwM6h
j7R95/CnoqyZk3siev5JHgE909ZT68iC+X2jEx4STZIltAZKiMVGvIY28DG44iYB
pfPXWvDlUqeBSDKeBl5IHfa60O3UQmq/G1CWUlbSqS2FTh0IuHb0ANtmdwZRQwSE
JnrvIL1ytN51hztPJuXYZEju26ct866YviwfxwLLLYBcioY67Hl0COzC9seK8Vo4
i/zruZ96rfJSQXocJexuBgHwuOBDAOGTdW/r2kFIO1udfoh/guO9B4QMmuuyslDE
2XvNPKwpwNnY4Ycrpyo4xZGf7AFE7Vnlii9B5YntOtM1lXDZMIaate40dhPtZKjM
2gb7UewGcTswA7tHcr7Ao0rx5B0CuJGIasV8zrEMw4Yqfr1zoJvVMf+hkEc3W1hE
Kk5MYyKqD5QhOI5qXM2hW45g66H2MkWjaaOABIfEb0PXzNTGobFfLSaO7W5g539Q
CXItO0dOGZv41S5z2mzeNGiKX/527jD3LduvHm4ZljKiVVMCj3aNN+qj2nLQYAeh
KK29UTHaOXYaRcuKar8+SxyD12slh25ar9kGb6KiNO7LdfMss66R4Cv9F4H+qXCY
z8Mm6abed7+H4C3miJ3If74XCb5RNeSI1h5PqbVr6w56y2ABYkZSPFIah5ImNXBS
jgCkL+zZajWdLjxT4V8ErVtqQKZlvhlmnwdLJXgF4W1e8uzeOvdbiJF8aAeJcZUW
VWJwanmRsHAOcLdc2ixzQZxKR3kYPtge+ykqngfMbTQyns31PBDFeAK54aOXWIDu
ZunXXVWgh4HzzJtFBqjeeeaSaejWY+jEy4z26go3/70pL1ZnN+gySWnjAg+9zPp2
21wWc6ut/6UnF7OecWjsDt/s32e/PRWb5CFzoMuJbYbu6P7A2jL1r9OhACVb4fAb
p2O6iOrut7rPyHROIeOEXqvHRJ11clzvlXElkdVSiVrsYGaQBkXLUM8qdVK7R/IG
/0D+IMcJPp1CnvfTLT0hhimKb37bub4n2l2NdLjXKWRGCxHL+qXZ/0j0yeP4kCFI
Cp9jnsHr5W9J7FOh5m1UWZMFCIQ/p49DXcoG/H+iru44kQ2Gq02I+fn7/zKcDK31
AVTDCr1v9/nHwkOreV0dALJSu2U6Hka8vbSbb4fq72ydm67hffpDOXVxmyyLiJfF
tpKLesorI/KLjPWUbSPfRFDvCnCpGA1Tjju55dAz3sAkYYabYa/XVasazDop3anG
0ZvGDJm34HTcCPZtpNlPjvZXtc2aYO7sTzpJlTfszuivfYViBFasopHjFfuUtRFk
EBCMdYySnd+yzAhGYSkXyY20JZBXCO8awOZjxDkY8dU1P2jNxAMtsJ/aYdzTUHPJ
NPSR1D/jrvVTSmogKKFpJ0HYo5Anp8igjbAUbRHvZ4QgjGeYcIIwotIGbJkZNN9L
utAEwTtURLwSL+dS4KrKo8QWZmTB/9FwilqsxvypuiyN5LvIeCsYbL7kDdfY7D+S
kb7d1Yt7KGMSewRvdVLQGAS01mGLp5N/5+ySV2/Moc+pQ6IROT55ePcGQw7Ukm8w
CTmfsCzWs8auewraB1D0a/qOy0vATqix7uUykT8A2Pr+hCqNSXrV7qsJBgu1OEkK
mIumhO6M1DOtXAE/oakCyFb26gxKeeNx9aVOMB3sSsrxNusHJBeQRAInginMnNv7
LpAKkD6y7bmLaL278oDP6ikhQKdaA63goG4PbqmUTXB5SqiJIRudKe+4v2xvrzWC
ERLIf0MUXPS3eLG1bOurDUBTY7VHfRoBo5hktKy/SWYWAGS5bImERzuH4EGVKOyb
tBO4nyORg8+8tS4IaCn3qYJ9GIksw6Mk/xDYw0Ah6Q67X+/K28qpsJc3VVuvi6dr
al3/7RX3YEVr69qQni/lZmPyjjWKJf/jMm4eBH977Qvzt2xkf5E74ya18ghG5jKE
5bWc0QVkLWWNTsmpz0WM7rnEB4h5+vyfebsLqUaopapuK+FkotoeNxhdMvBPg5Fg
0PNaImsJhEx4ZxLANJZabQBDpx1/hz7xEcBEsAOd7YDFXHB0MxxKZmxPbjgudLg8
n7NV5e+K/j5epIKav8Urk2qNkz69nsENJN3MxxRgAWxgVEsBOrl3XHUjgyD5sZ74
v4DRbPtMdtNzlb5zMO4msFPYgIDXEy5u/MLZEita3WTfbA3rY55+8EGg5gX69Jpo
8p/z3sve3G6VhQFBRr4FriZaU/M4DNx12I2HCwbilwPq1sNTk3zoYBdkY1/rW7i8
tByM7nx/7xytqELa4xCtXS3NayyMKbAFhykpoZyYvsDYOn5mwVsYbmuaeGYy23rT
z2q1XcegPA+B9nYLFVWlEDYx1u24ub0O7+g2U0VjmuBBH5VPqgQ66+2FGzYM0pq7
7YsL8X3qyWmC7nTfrdvsejX3QRsdCybL1nOvUbjEdIfmk/HT9yNphGnbK3CzTfH6
5ZTLjwmMfq8ZgxJz6qyNYxWV1ghooYLekmtWRkuMs67CU3islMZpJFCSfS0n3Ych
BkX9pD00jE5jHm58+KC6NeyPlh4PfPnR3aHPDYe8eawyk1rwGx/QUf8kmy4iKSNT
2CdKLBIF4a9k7sTsgLHthpUEdncgd20DhsxBOQ5oIYa3evv1UtGgwh3Tg59kVbiC
hrbfkjvPIgy9nI8J7RxwzfUJA2H6N4swQRxW0grmmQ7utb5bdxgaAS+AblTJxinG
HqucZmBA2CImR7pSAsE0CLs0RAjSRGP1/lMX6gKTv9RLBUmcFgf6zbVeAg1xVIwK
lMxsOQNGTgGJXVfBR985V5bf/pf1kCV5m7D9SXbSty4xBLP6+62/SJMytcpfZ+qo
dEAXKtl5sMYvF3GOchP/1kkkYc3DMYB5SfS7dG5Is/nXyGV2MXWEhBb1mtgPk8BQ
ta5zyKZ6lkRGlZ+cgSm+RtoNW7HAnDfxawaV4fVH6V6C35YPGC3d56ieNY7XZ26e
fIq2OHOgbRHki/U19uqJ1MtAu/fLd01/DZemTUBDZoZ9zH0sMwt11jY+qGsOxsbV
XG+VOMecEiMI3kWvcvNTBbgbG98ObBSkL347MLWcmI8sbasDguMWFDaTa1tCRn1X
iJ3cOlVy/T1x4ZzR0tyoZFPj0H97FMAInLhHSYuoKGprd4Np5R+eRWcrk+pTsnhx
Kgpac8DnKv5w0VDZ8g4WQDi6GRk4Ad2b0A5aTAPIV+xjVaP6M0UHFk20zzuO48rp
jiZ9ufAc6nZrPkAgahcCkdVUdutN7NapmqFKfkXjacQal8wotexla/mvjH5krECM
wmgF3GgFy/u+xCyr59Uld9CKAhyL8gPm5wD8k2r/uxdFucJpu69/Y2WZUe3d3tbF
gBHql7O9EnWD1LgIwJ9EaaaA9aJyJnvMVsnwmaGAq63QUOaGrjRe1pmMOOf/XzLb
qhw+12gu9URb8Dr3wk2H8t8gt5mXAucfo91vjr+HWRdp1zD0pxVaZ6T4bZmTxSEU
qdIuHJtotx8oway+II/ZdvMJlOkFY5WbyjTlhcXuVa54h0vepZ4Gq3ZC85j6GDd/
E7bE9GGgyPAQf1x2MkX81ZEdKmQ2G5NdumvbRlc0fhKpETTyPsMLfVgKqb6co6a0
50GRJEI2sdGS6ImVpBx4gRW0ssuIZkf16dn9QNwrzpasU+jxeFM8tmNo9dAxxuT6
TR4XMVl+oGFgAsmend+AIgle4wMAseIawGLXT3IFbuztywx6jwDKqxPxwLybOOir
mI4GM5+WWgRqsxfwROgoZxurFDUXaYbxq5C0r1CemjMJD4oMO7VcAin77zFWa1qX
QiAp32bjiVFrMUhlqIW4pX9jDfHkDPNt8DvF/2pWkghufnsTCsSX3Tnnn4t6seWD
SVqowe50kpchP7PBLYN8VSstD7bnfYHNQuW/X10TqPOn/5eeDzEi9buHbvQjCSUv
vhKDOMUjQPMpLYYf5sygAIn8G+oHGc3RsnZ+gHL2rNgcW7Y/eRIYb0tyDzQxz9Is
YMCie6zRliKdBLsD1MtDqgPU34vy4mdLVWs8fPu6p4+znNuL6HSKuKcbk4ErbC5E
QjKF2vfNCi8gG2daUp5y9CeYYKqo83PktNKS8NmZYE8QtVUQ+LtysPH6EZpIaz8B
vm/u1x9JmgkE+eQxz2hu++AI9RjXxquZt9c77uQxFGAA/WyMkAeQ5+qSg0b9O/hp
lAhiyk2GPwojlnmiBQlNmbRYfIbkoBrOT3jm8jBb9meFh6wLWe5dw1gXmE4CyPKo
A5ZDWeHzvMi7IS97B26USO1Si9/kI3QrZVYyEvV3lE8hUr6lYzzymnYlZk4KCyKf
IaQKS/8hqwVswRsCBw2I8xAzUw/PPbj4X82+W0ak79dLzJ9xtLKAXV9Pb7AVGRbS
+tHB4mTpGHPhVnHO6/rdGmWsuRJ1CsjLxHDyG4ZX74B9e6Q+7mm1YBHXuhGARh/I
gX9CDaiI+OoBDDXlUT7Bhhyfq1owQ1vutT6v2nD3gtqsdURcWFyMeThl57+aIago
ebJLJ8rmuNFaxAXqqW+KV+8ipxy8/01vuDM/zvafbIIFGxO/D1zjck3+9jS1I7Zk
CXoCnMxbqRrwMFuJVSnGSGlwrhBdifFiWR2T7nC+VpH+THm/P/dFxmHdr8IIFqWw
2xcJ6kSUNuPLQrKzsF5BKfE47TAbr+/vkxj3yR7smSxU4AAsBB+IKEBAyzXP+cLR
7/35ND0+h6XYfkAYu26EAXKY21Vs+SfqA20aLndkF2jbzvtZH9e21U74Vi+vXwYL
A3VjkIBj8YzU75XqD9dvzK37sNL6q00oCub1MdXp0x6BShdxGLUij0g61HD4Toiz
FYMDq+2PzqxQlFLlG6+KkBJZZG/HmJQ37iwQ7xzctQ59hbVCU+CUC9OnMPfsPuhk
Aif9cLnMLVWImApCo+cu50Hx/JtLz3MR1cSXuD+g9esyaDwKvD6vj3FiW0y3FHJb
wj9Tantip3pG4e2576xrrb2/k/TyrLLMfC1h12vzwShGdttP5PtRiZcFpjXfST61
LLiuZeA/waABgRAGyfkLSCcqJ9qVzhpNFfkAU4p/HKhdzUPDfxysf+hMEToi+462
nIX8BZw6+tU8HMDQcdycSUt/wvrKoQTD7N5jNRobBpR8E2OtrAW1h/nuyOuQHRl4
q5/5IYnhYWuvp6gniVY6ot24jMWFP+kR9/+LDs8i8ijRfrWoVfQqriVqNOUAcOZe
8Pfmatx4c/gd78YJreOZx8+o9IAu5BiHGagy+Y+lDD27HSRfrxs+V3Zdm/D8kpl+
jn0k//kzPsv5pQP49Fc63dAC7qVjMRa5wExnkD+ZW2oQb8pgzO4lS08BC9HLOc2T
FmZrxdNWbEm0dU4jV4GsR7Oy0TINMSGPb52Bk8XYFeum8QWrprWT7nzI5ytaiipd
X+SzamBOZWbHaWDz6kFbnKevplert/+X0p4LpjM4AQup42XvSuIjjtJ/XfweZ4Qk
t/tY1ype/jbciDb9HX7mqMB9ImNgegBLsOWLEmDKCfrPbRe5FRaJ09D3fBlitKWF
ms4+pQCHxyOJcYW5SgnY0YxNbrlyBBA8EE3sE60se7LOSIZ6dfSGdeObvQAQzDQx
7t+2OjbNNGky0PztYzed0aWoanS92AoPFeZibdU34LT7YdF5Ryg2VmO0CT+8i3yD
6idHDk4IgY1B9uOGE6ZPHumFb1bUG61VD1JrOBRk6gD/fSICUyfpTq5WhdSjaDOm
Jr3glRrWw1PCaF3lIPUuKmRuJ29+JVCb83FJbyGwbePwHMxHbeDyENMihT7cb4sr
qgl9Mg6Ni15k3IhXkk5/Ak61MhdCpZSYoJ0+LPpsGExSyMwTQ9imGF/GmZlJPSJx
yg94JsDkkYmMgMJwxH5zqyJOwLN55XPIn7bhJ9yXNN9bj2Ls0kZ46kd/PXaCuEhM
smHkbehdVaJbYTxqR9IIbvqCAgJeEL2pz3m6naf/CsxNyTDf13sW5ggLhS9gCDze
LZZg8SpqccnK7h3G+r5J9DuIFiyvbDfgbp3TEsVSac9FiAjkLhz6uERd9xyP1z1b
VbbpG3Rhnjwu638fqzu2qaymHXgWxMGt75z//LzNnIKW1Hemm5X5ivgqmuUdsSuL
THWZlAkoxW+kiafk5jMgOoo1WLIaIeNwCMSToBXxv9ilvhdydZWEPw8NF691IU8k
RbnwxEmxYs5t7ovzYLIteJdjgG7FOTajUXxipnUtm7JU+XC6zlsENlUdHZ82Vgxn
AJeiPaHMU58ImBMUGEfVmfizUfAD6mcKjgiCvB3QbVYl85pv6n+7umF3+QJhmFId
TY+vzqVu3K+fSPQYq0ujkOo9W7UKByp2C7J57sR2a50fj+CqSXuWoi/LgnU3Nusj
1x0X3yu1j3F37+LaX2LHmQj/fHkfqb3NErQE6uf2fMQCyLFpZXz1Uwzrr86znJFu
4QWTC+F84ai4MYU5E16nv+H867EC4KRJvPEv2zW4FsjqZE+oI9K1mfxpEKnjMSBO
l49DSIamy7CoyPL2ul3W+NTKUCySPCBB1Cf0Oacvr4N+Mb6Jmwxo3AvgzIdX180u
pdvsDNMBSj90lN4NzXs3iVJTro/FST8qvLuIRMm5G2TK3Lr4xjnLU78LHyuc1DvC
lOYaGflPOZA0N2CkLq1tnokiEebgFGYh1V0ue65BKbPZeXrxundxz0dIgSCkbvfu
ujZrgQiZeeY0SPKfoieyMtCgitb1YlTeBZIvu55FvPgSAYvSKPVrzcLYQJQBeweD
y5b3uE0Tf6ZheNiZkc94VXqO6kPJWDb8zBFEv1+34V5B3qKzdDUZ2XIYZ/JrrnhN
BdUdnLL8NEpFXQ45Yy6MADVbKyh8UDaQjEA4A2Bm8/I/54ioZuzK7wZ93u/f5bnN
rRKG+VGqWdfuMi1WNd94gn6FzTn1xV4rWE1lBRoBrFpDm3rG791FaZlryv1yfXT4
uSuIKLq2x9sWvHlwxKb5zAO8nI8psDEOH13cosLqgTlzNGbWnVjIMG1kXo8YMMjj
a64ylFCFoYpOH/dd5UXYaUGcwfooFUnd3eADPU/oIny1rAdqjCDBqMYMixtBfOQj
vHsWcLtYJfowkRFx0ludRvXYF/bgrqoViz/KrNJnmZ0JUeAHPPb4P39D+J8gsFyl
TRylsIeuQeRYRUzEEgrkQAgZ6Io94dnwuoAIMQsU0PEOK0OSIVlS9Q2krkG3aXtM
z5G0+Nc2cyh62u5MpHF8p+gANLZkBNxFymTBtLwTVvw+ZwRrOQMyPzyfug9cz2xM
pQjmX+euHhs1Wc7TgG6iQxNYJRrFHQRvz6EsI22uMYugRWKEfJvqawu4sUcvwjjl
BfSKma3tEJXXJHXZg1pEPuMMoN+dOAvV1PB1FGJiSHX8D3PDPkG/RLrVdkImiag8
j6vX5VE7tqYlfcdjtIwlCVIzhHF915rQ9BCxqoiWbtr2fWuiUxikeD2HDyTYFrYl
3WUo0WcUmiQ9Rm1DlxX2EY37/c5OjWy0oqTKYop4DKXf0ZvxOsJA50tZo5iUj6tL
v/VqX/tWhJkBpBI76T/b4Kxug3aI5rmDxYXGDYoi+OFeyzhIszy3d1wj5prKYPtZ
PhEDktOa1GgWsDYahHhP2PgLCSnCmpwl3rilCHDYcgaRmdH0coPAIsVhRdjggMvx
fKD/XS3WKR7oZ79MBmAC3vkqtDWqsSDbbv10Zn9FLnSIZ8yG6IKxSRmwxnew0KyY
dKc4gfv4oK17GoTJXvfN7ELDMuG2kBtrLU5Qic7IqV22rOKJipV1T37CBNbyo6c2
c0QlwNMiD5iVdChFIaoQ6twOwWbFxq2emIopW5fhNdYw0Dj2+HVikzlGt03Sywg4
9Z6aG89vltw6u8Nlu1IUTkYza9Oa2jZVfYv97UXTNNmWhYs13PpWJ/RE1lN/sA5Z
vE/DpkgHNtFlsBBHGDDMB4eER5B2W+1gO8bMmV+UD9Gu91aNJuWPC+MtZtlhpFFw
a5LAl7xJC5cXSf3iUHntmyA+PkYxuUxwosIg9HuxvUC4Xepy62ZUjZEIJNYaN49P
91AoZgsFMqQ2tHFo9nqSmwF/jvjrOZvPTkeokXZEpQ0msJpD2SdtSMUOquxyJuTb
8WQuOaE2Gp3hc4vlCsnCSy3/5FTngVtwsFN/ZkNIVIpIxCnssQjoaxInU9dBxqdu
CxIBnvv4UuI9yuDoYX9CC4qUCxY4V5U0pMy3sin8Mz/aOG7xcnoXo9XpUnTPyT9K
JjvjEVmkxtJ3Ef+SUzoJiJhCW4WSd3/dOv+Q8ND965tqn8lsCXpyymyGsW8b/HFB
m/Z5ZJEcEZftRXaB3OmwhprS0ul1+0PT7SA0QJPwSVoQV6PWCGklfr+twQQEVIej
Xnx7Qh3Zs1oaq2D7Zh1ciKGfjrEHwo3jI79GBmz67Pvpkm/HLc/8WDn8Eh6SwJhb
dTJl/wN+G/nznYOBLaKoelfsjLjg80ItfoJJjghwIay+YCoci8q2dl62aVX/Pdxu
oTcn78sWRxFRICrMP8EXYUWTbHmCEu18uLj2SnLMW/4p4uYqVk4BFvHxJOM36OI9
PAM6bwMVrDX0fELGkE/1lQ22r/ilLje9k6WUs7mjv5khs6/Ws4f2dGuC1O75QM2m
GQIt8tGnGzurduIxK6qAMiJr4nhwg6JqMd4CvfspxjzqPHu9lcIQwoj66p+qKfyP
nuU1Mp+vrBJaaJUbk8ZfdT5W8WSVuQKRVrz+nlp3cm6XHrigrGtahxrpzB1mWpeL
a605W84wj8cDKDZ/Cpz1PKkH9JCfigHl0ZOaN9et4r6vK7rWHuTbsQYi29jurByB
zM3pZe58O4lm+WCJ1oFNj6gtKQa/8uTiE6EErLz2mNGkxGalVuXpc5Rl3ljdgAIl
4S+6uwFpVSVX6Ad+lvX3aHFFxjzRt1MiKgMLEIZhhN51fFQgA+1bt79h0yW+cO/z
LLI+kW2UV3hgILg2Nsj9yr5HJwlz4lKs9S1M4Nnpo6V37FoXoJpyCldGWcU9wJCg
xLTg3er2VjLXsiMzdYe8GwTHBSGTrch0zv+EdfCUfSDB+zabX9AUgYT7beYCZrBP
Z5O9Py24/jheKuicgGyM3DoSb1vyqJjyVlSw++5aHK8iX/bqblyK6HjOd4bgONiq
FQvYG7iRc369ZFxbdGFyn9X3t86rwhynJhLUlSFUdmiQL/n9WCVSFxmeCehKXs74
xtnHRMxWJrU4jpfkhIHkD98TJvFr6Vb3wwGn2wuxNA6wiPi6Lv+YIXjt4jfrfDQP
CZ03k78c+j1xzCC7uhyXqCeXdtaZRz29rS1qB0DCh6ynpEGicO3wLzKiAtTB5dJ/
1oO2DwWI7UzQLa4C3EZd+B2ywMTZa84JJuuYZVs9oOUDbimh6z1wh6nPFA/cKREz
OYeAOgAZViMyM99yjqz/+EAxHbnCkSfc3dgdHIAOFy9OxN4GXdJqKy989+QEGpcZ
ICRlwJ+9PRMIkPhL06Xmf7aJUNfgDBY/UdRaxCc7v4iUBYj8rxdcxpC+WWjo6gyJ
6RG8gm1gmGMH3aSJtVp9eD1LdwQaMzFBkcS37OrDYWEzy1lryeAgHtj0JGnS6KCa
+AMeaUakgulC1t1WiTebVIEsG3DcZxIU0VeQ15NjFbjlmY9qEQIk+v5v9VdRMOzz
HqHZR4fdnt+XbrwiRLujWJOvgX7s21wniyiuaTkcZ9eRmcVQ4cFqaCKRK5fbYv/e
B7RmLL7QrLJzet1Eb0bn0cUumwzfeZh0trddLvqrOpdA548jMO9gbEBi6VEeYMkC
SEvkE5Bdzp2eoX31zLRFwu71S4TvBy0AK1Qc2avyIFFPpzqr1vYS1IeymyYPUr4w
gqzALD5An4sF+nUvrVaba12W7ATdaQXee4+aGeZX3Rjd7MqXaeuvrvCtzc4bUQtR
9JeepZgvSJ3pNAXZ1bMWaZBsscogAo7geBNmbMdapGy7SjgmyGczLfLUBsj7HpRL
Mb0nwVzfGiLfJfx4dFTufbf3mLotEco4JHkEHpvLdcU8i5ejGcPF7zrIPAP8e6ws
bZmTsie3Y7jiCQS8Yuf8YhLAk/kT/fu7pQo2Zrcu4q3s5UwxlchP9WZUzRDKivq7
Uk0vaVRrNbwVcyZ+UTqvFyKcDYWizaMPVjZUxBFnJv8yhm1YK4NjIgfFBaCajF3G
HpN2W+Y2yJ+wb6eqhXyBHKxFpGubx9MzuGXxpfjkTg1bin+CvfjGT6GYvPHvS0SS
xRQVivObEdEjHpTWPGuJdMgLabKhYz/quKdl8fEACXT8oqwQaO5kF7r3W62bPxFa
VwE+sNy+Dfc5zj5CYhb4W59+AgXiQG/QlmhLvkvspsySSJMT1bXLRLYgc2YR0B37
W1JY/FfL8k4Xjf0PvP1OofnU9GlFpWMwXuqVN6LmJaQw8gNYAfuPVng0xVePRWo5
ptL8UyXqbegkmbEODzmqVV+gC2TzjxXBS3kJpR5ADeldUeFczYw9nXy8Xs8yx/ur
JZJJ0vnHXR3pqC5s6Gh9hNfg8c3Fu5zspITUBIfIvS+vQLKIjBmR6IeP/z+b2PrC
AmuWvnFYrhCzrNEbNzPVkQ++1HELhV3y8G5XkVdP9uRBRFqoh2Ta70WZrMB+meN1
UtkQvAraITpWa2sZ2STspBOcgREeHDJOIbWflw0n9Ji9feADJrVQGG0lE3UVxXNE
93V53jKgduJP3heG6eCeLGtps3gDhYjhdLA1DxUQ0eq3ki/qK4aw2mL4xtU8JEpn
7XBwEpPFX3C03K+o97XsK/sSwSgObwCqXUmHl31gi9D58ctL+IizQ00R1FieFzlC
HwFSO+Xsn9jhQOFANVf+wEqt/CL0/in+MTwQjR0imV9sx60Xf+8iRSV2lJP+J/Qb
4BVV1XPclJ+eELxFkq0lizfd+Gidz9izJHMHDyjApADaQLtcIiAnSS12iXZpj7Fj
vV/h9C3nqJhr4J1Ms2FIlCvEASeY/ctWHHy5w06dwqVd8ah65VU3IXTf1iOfERY1
/PZgGX56WieFZzHn+yU1ifhrwb7HXS+3/2ynJ8OTnmWWFl3h+jnn8Ts/VvziKufy
yFe+uT7tfM6OlBmv3ADP+a+MciRhgdN5lWoYVAhC4LZJ2aQ4T4Tq4iC2lWN89/UD
8z6HQtYeLB4vnfv0k7HaghIMK3q9AKSFYeyXMxSh399dVFIbVWeWEs0lQZ0OozSI
HD+bD9gwMR/qgP4sJN0Cg4uJUvbIdQDriaot0SQwnqBY0FMMShkBCsyBSfi8+km3
OZLjezvpv5ua2Yp+hdaw3e53pZjR/xmXwxhknKyBQRBPiXPgZpnRlIY87MOoyoGz
CZiXZbszPhUq0MvV2ZoN1Dn2Qze+xFAT3VlOs9iG7YGt+SJBIRgzMrx4p7cH1R8O
XaU3fzsl3TSiesTqniMCaknwgituRxGiC4ChksdRXSoLxO/+AnPZXgmFrgGqPLuz
SPRj3V8ZxygoAh3XzqcgsOh+J7Al8Ci0KUtADvFUI9cHXKoCQCjWY68/llpNDtf8
zeRjeIeJwn8B0YSIGmsIfRszuWbHFxeBUbwNR/RqwA4Cn5Zr/Y7PDank+w4iNKX4
37mKwZKiSF0Ek6tbS19okhl+V57kOLriuFlsC1uDV5mAwo6mjHq70YvYSTUT66my
ud6uekQxJn1+kzQxwQ8dU7fja9uwHPzm3TsMicKgjaeqISakDfgAWTR5qtXOJ39J
6eog4k/+EIG10aKv0d4W56kgN5wSaqcD/Z33a9DY4tuw7Ono29Yfvvlsb52dYFCK
BH+lu7B2Mkrz2bgpVIxh+yDKU6J5LX5pAv+/A8ODQbwDxrxS+eZkKzW6tOxv4efM
wHxeXuDIJ3JjvDbUh78WVF9NL8wKMqx8BQVchAMyUf/P4HFxrVsQIRizVW450ahI
TG5NGAanRQI6P99tlJCzXKc4tUAiRsfjmwBecmuLuDdDmT82TjeJji71StUpZZRv
Px5feFj85dCSRnGTb+988pFd3IphlLFA9sjhRh3OZwxC7mNKgEw61xPS5dJ9C9Mf
4uG69/045R2VnIcOsQTsHlDwxKinZbmpUGASNV7VOGHzwnLKDG4VfutE474xuIvd
yU4FfVINW+evDaHMbYeBVzJDdwyOzzf+4tqwFI2+P29Ca7HaHnVpOhKE5Lyjnom/
7ldQYY2VPpQO8EjuFgRvmTBHYLLoXdFqHn7DB9hCrIXwuW1/agqyutI5GvpD2n+s
Sj4bZc1wNWJsyXDM2Hy8IPYk0KxaKTUSF95m9YgkpLxnisadhdK+kZOfVWBUPU4+
BlvrJs/RPH3JCAimpMRxsT2stLQkZUzHdUKHjwflkCos/THEbpLpaxDKaGnwFcev
6RcxHKS12xETaiqbw3So65RS4H7tb7U3CujO+YhDmaDdjaqLMcl3bwZ1DL2AP3LA
kSzF6weLch+uNhmkdYWA2lWk9tYFhHGFkpPy5wzmz7OuZMYfDZAlWtCAdGzKf308
tETXlt5+IM+gdO2Bie+dsrrA8IwiTjievMa0Kl1EZzppRR5fFLcd0/YOLpgpYDqi
ek3Do8tGzs9c2gRmgiYUC5OiOWFtlyLZciEIfT+ylQbfXkQp0sTSQuYl093X5aHv
lHUoIFkY3AcAOCB11hbSm5HuVvI5g+NkDaNZh7hTqoWiC7iT3HWZQfmy/XJADQuo
mp9UZYh0sJ18DPcU8bWJRAE5L+73CGaC5I1u/rFeA16oANdpdJwGmPZfkPcRozjQ
3t2WkQaHl3OYND8dWLSYfVaCHD/R2KGRSYIUEhiMfCq1wCox1K5uGwYVFZNyH0dM
OKvNKRAzXIESVEGAS3wGg24F8PSjpuqJ4bjX37Fa7d+re7AcjEKgx3ml0lY4lsz+
KPOlAxm/1HGRWO4iO+KqSvgWcQpTHh3mLmCddccoy1EbImPOVQ5fViXlJze6Fke/
+3K49xTxc27npKD10pBgSzMEdbbWJNtAcsWvpABbyup13xA2BcXdApoXg45NNZvl
xDtWW7i063vnxC7H0wCLUisoM48H2Bd/fYKffrJRvs0jXmzMANy2hIvvYvcJhDXP
MgKgaZR089Qd8UGSRhSuvc0fCh3YlGvR5JXsRD010Hk012AuoxFg9fZJp3gFj630
wAFKcwwaDLRogJGFWpUYnpnEc7gIT5BhPXm27nI/tlofHDfGUuVDxdktV/gP6Q0n
PgsvrNrEcz7N4jfBDoHBSnshn4YVnyQcgR2joDtUVFuRAiwElVPiTTvLhgY/gY4E
0DTBTYAa2WG/EBD8yr6wFekgC79wbq4G3zcMi5EQ8JGryfllyVRkwyMWPXvIIE0D
v0kEFtUCLf0lQpd+osQgbBmusR3T2Wr2Kl1DxYVjtDYxW7cCMsXYZc8EPaJ+Y6sI
Yh5hIM4ARvfFobgdExob4GQgbod9hE5HM5P0qctDwUDEnEDk2It0HdaZsAXO+IUv
DZTIeson4VONDwYHNtMe9336ISUOTL55SlUY+A8hGayegVJbIY0yyDDA/wD6DbRE
VzhEz9ifBICl4NzNv0HlXEcTX69vfkVSII+VM5bGEfcQstNBt6i5HOV15ZYXcnUU
Q+V9T/rJXqbZtX5KzZKGN7c/BguBbAcduF/E68iMrwqOZPbVfzEnqHyklZaJpOwA
S1cJsE0jZR3lhWcJkgxliqt7psoCYGRR8HK4EtILi0Hoa2EC/Vfydeepaf770eH6
wH63wDwpR56k6PbCbykl4PgT35fdeym7rE1f2Z0j7TZTfBDT/ChfPgOyds14+oVK
YCdR63LClS6TyAebwwZS7PUTPZ0uaQoodwXKdpDPFP7qXg9egv00ym7szAYKNr9M
nh41o5/1aq0sdth7WU8ph2LjKrjBLtBvQaeVer76+nmgLlzFsoD0cpBVCvrHPqep
WgAbnUEn8CUBXm1O9npPfRcvu1/VZNuXjnIlQrLQE0FF/In8Ae25ievUBg/XWLSS
HtD86+YOsHIUL1TzlLZ6hx2dFnKkxP6xmC5Mrx2AzqOSmJMTBUebWRymE545fbsp
QJuPPEBHkAbaUXcnA7TlY5nnhucpRL97yIGKTo9y0Wx3p8H80pNlyyVgpCZZHKdD
FR9Ov/Qi9RLQPlG+7JLeVCaBJH+fFK8BlCfLKIo+yqmA99eHMr7QJX1Y140CxXov
I83TfA3Tb9gSs3p5M/waRNObx9ihv93M4FSImm29fsFQ8P5MAwliYZeUhKjcFliL
sSUxh1Y0Te+hHpWmbhbeuNM3Gu+VN4Pcbpzf2xJ1uQN+ma34ss5N3rF7Mj4e18dk
GnvvJ7hAKm/00buAo8MeyiEd8olWedgp8Xp34Tb3v3JW2flW7ZYQtF7P2rtQ30bR
DIpP9C/UdexKlUaeqshidiZhSPSEG8fSsw68RWiJv6qybRghAiYe/i/yxZnXAZO5
mLjT3IQdp2iYXptENhzHrtrFBhZokhGzzRgNxFcyyXmJgFRrFXi/7Hp4Toe0wrs6
+aNPp5L6TaYJ8qdYLHytxU8bLHMZx6KFiwqEGWC0EPE/tNUFbqWulX1qEPOcHnBL
xDQXAHhfWZEuY2T0FdHyxaPo8+Nf1yB3z5u9PSoIstFF5CdC1HvtBY2Zca4LH18I
uCfeAJ3HzUkF0TcugcR6BhcXRqT4HslvxznU/YOVKsey7285n3MPWlQEVCRtvQ0p
/bu16JG9i88YVoxzS9T6PVIuAbYyU31J67NxE+/Y4FmZXavUquWSDSkTEifI9Oea
iXZLENozYM+5yHQy0cdc+2OPifaI6zuw3LeTa5et7wCZD2V2TzMQn+/9S17bt8dB
NYz/teAKx88qHhjYprz21ENpzjrOs1WbwehePFVTgx9akA7d2GelQV8PCLvUzNzN
i0z4k3CLZLxGyhr+Ccpc5FHYcFXS/A1YWZug6v6yF0Dg/e1gQDY2jOTJn4cXkyVU
iC/slEk1HNzKW044nZcni/X8k2XwfnwT/6mUsftKflWW6oBcHLEYIWlxhZl7eXsC
/il0dMd4cPnUEF+OMxbJIua/iUXN0R+OGx8NguaYsDCr/J0XSJ3F8UqeV8Ihg56u
kQUNIzcDuKOLYC+3Qe9RX0gTTgdrJdvlsRmqwI2ZK4VgOa2Rk1EBVNELvDQhynaL
JKlvr5BOMf5VExqQN5DdXvRFE6Le/lMv9GzhUUEY0z3C/F2/Hf+eTqS7thmoOgJ2
KahXjXGtzsvIwhsCJfIufxndjsugevckpe4yin1ozhO2waLoRPaJiFOwXLoYdPfE
0+jMi47Bv02gokLe+VOr80z0XsewsFsM7WFM4JqjJKIT7fzJwo0jedO2gKHLeuz6
cS7hMnMvfssd5+5W83uJsbim5FhAwgYeryiUl5dx16nvABXn7L1Hqj0bvs14Pyzo
2aftoA530G0d2R1lKq/RSJ4EXkug1MvWFqc1nDxjVcYoAuw6r6v6eU7X9SKXMwHL
b+rqXYLIfhM3AeUwtPVqypXfsaIlXuq8E71BorHrbGk36aennMe4mQNITqrwvT3R
ZM0lbGUOOkJh8eB9HJIwpAf41AKR/2WbQqgFy+8KJe0U7NlAzd0KwNsGaIWac0Fz
HJUDoJH0ykiRLFiLj6km/Kh+2+0mtv8fc1QTE7vM1YzocZggWdRB0C5d1KB5HrAb
J0fyzpgtxNH/SSlfnNRWJRkFUe0zk5r/qi8WOm0Bv1T1nKwocbdrYM/7ldKXfiZc
qbhuBw5idE/gD4iZ9fC/mvBq0v6JlPkVpn5dtP2Tk9lUAwOBvEmEESoODM8w1fqi
IrcHZwKR8dNCptXGC8tPVo4WA7+MfvizKY6JrrpIvIs7YDjJ++ymDIDTjTj4CVUY
PJqG0xz0CQ7qgM9GyMXFxEEGURhMsKTfvBd12b3jD1vXXTucHBexktZo8mJxUI83
GOZmn9K8hbz4L39yEIT/E3gO/0TaHCvqO/sISkPyJW9asiYbo2+i/1lXTvFCttIp
kUmBo09YkZ6TpW89EOC9ipa2WHOai8ZnHc/CWcI4BlNQVd4TT0RVDh9vKociDU29
efHXdn3RLqQsPPfkeCwwJJlHWJJGXI5MCQEvyXRKu/ngYbNENl07RFzlypRFCuIn
geu8nimFZT3mo9PZ7DWf1B5n2Oehxckq48BjOZDKW8pkyZ8tjTRJgOLJkNR7hs+r
JzCk8dU9zpfCZW2Mp40QxPbYr9EeYFAVSKlXSZ29cvhx5BttPvL8RzU1mYRcR73s
+GqryzwTWRS5IfSQIm4Ck7hl3mgFrciW5ODcQ05fUNNyWVbO1YLO195w+rSSfJ44
i9SN4Cst45wGoKK66wZ4FuYdcgAxC1mAlFR2txo+OsyKFU8pTRNJin7tm6RfsI3h
92Qi+O7O2w94RBopg+Hrchjy3tgL4cy+gGKWzEl2HWmvOdaqvbmYOc4jyoodvO2v
PzKSb/7s1uB7YlWSC3LzwQts6tYWKGbPJcHyC63CCWemtreUBJV/QNpj/464bEsk
fYP7R0eCjBTzdzOXzRPwfLQSsVkEBfwS0EH19xbOH0ywe1RlhKXZ1e8Zp+xyKPz9
NLEug/OylXAxWyJcM5pA/tJVmGY9YQutw9n+T+m5aV3dEOczUYMsU/oHV33BgaLn
qqyUGB7vcwDyzUyABnmHkeEH9N1U9GsgwjO2BOld1BD8SgxNU9YbyMaUq5YFpi7m
V5kg7F2ZnI6BEs04dzBQxkC0TDiT7r0+X/IeC2p90y3Ux0mOBr46cW0k7oLpIbR0
dV0rfWiC7JY7ataxTZFIzTDkDCPsV/zu1aCLOcIm7+SnwnIJtYOnQ/8RcVJ91xf9
RdLfYp84PKq0/AykaucBq618bwfpxYD77ZGQDCpBSqY6Xsb5a6HBs3EpB+TF5bK0
7ydME9MmVBNHPoclJERrb1VDYHg8wcJ8VnWzHL6tvBJM3gdgK8dKB5zzgNGpbdvk
eoKFvQmB5jfAme030x2dTZ7JXC9bFSKTcsRfeFL7tfu/Sk4Jt3lbsvySnqxSk3kt
udHo1h49AI9mNZ3Nd2flEDok9dpw2JfMMp+4+2U6nMPs9mIhySN++7vGZgmNpu3H
acTd64kwe0DrDgcaGIrZwvDOWFWaKE/TTB3XbXwM+yIp3KCy/LNSQ7rhRwq6g8n2
oc47xfSdegxYityM/cSYAFF3UQItDDj0U1e/82T6m8fg+N54WhR/4ESYX6543T73
ishFKmT1AAVLF6q4N5sMQrapVAwAjzX3Cu67lZfTuX9hV4dno28uvU1tadWLDIFI
b1nSK5p+zBZiss203TATB/hEy0JMb8OGbM1QOnjfVYDoOuOfMiIqKBErICt9K9Gq
R1rsm93wIRYgWkh1HSjnJtG+oJ/1RFpnUWbOHHyKYiPuLXAKCYY1H0Y/WW556R3x
/2xAKz+pmQE00kkEiVNIQNvlTkX9cJhnbrXov5bvfLk7AexKUbUWiG4CIKO9lCdI
bETJrJU0lzQZikhtyHPzGCRplD3L5sC/SlxgSFG/vGo8AIH8I0KtZvIAK0HBH1Mm
OA902uOT9xjHDxXjIMOG4i7P4IC8PdUmB5c9HT6pyxGQx+l7AjGcaGR0fyINFomT
ztkfrmVePFdO3+mGqDUA4JsDzukqtO+t6wrn78KqdGeAY1F0v2RbQiGlFQpJBuNo
GtO+rJ5MRNMFCyuuptMY8b5ZDKxXiYrw63ytGu/GnzZHGJ2h+rbq2Hj3MqN0TZtk
IddwvhCUqsRZ7Vh1ygTHicqGuElzE1rBnkvGoaW93g8p2el3ybwoaIpxQFnvyjVJ
Th8wCwxDcKjRd5sR6G6Ii6w5SxifFfjXc3bK51sfbAf0mECb5xAm9kqGdrLXmowZ
j0OS2FxDIct6QggXVF6bbic70YaYupcuksagr94OnJ2QSP4NIp0uysD2WkVPs8WY
QG9Nnzd+juShKz/Cc6Evy65wIuMxGMz/4BjhHOkAUO716J0c2oIwg4iZ10mN5pXa
KX+8mDCLRa/EMqWh+G9t7EdO6c0eYhCsUCRJh8mCXFi3a3uHYJnRpzVssD0kNQik
HnWvnul+RJoi+vLgNiUFW6/5ucxqwoGGIyQI3jZNG+kLP2jGDLTL4czqdg6t8XLf
c9aNKlaAKTRpoHKcKkHWcokbgUqJ97tsQc6NazDU/hkYDaZ0ZD8RJtr6AMSJgdX4
HCBjMnilqK/jVFnCFlVg+iujSGItEWZgZAQnudnnAesfy0r6DlffxwW2PrfrKLOK
8YmcQK/MZiSP4d2qgdAD9dFAob05xFnReP57xYSIzTddoIX5vkpYGmKFxSsxi88q
W5w+SzjU6w8a3vwJY9mj+axYBQRJBTntOyC+2l7ciBL8A2LK6fg20TwHfvXdrgp9
NizhB3Efw2xLp5xFSzv9eToXrpNiRkaVYac4AEJqCG2xA5R7IQjtc7didhPZkM2+
pznTz/w2TYNu1rB69Cvkwx5HaAMrpEjUuf/7+n/Y3gJBRxIxpdhUhlARMw3jUapa
9Gu4fv4p27qt8Y63CPdOYNAmJ+G9DuNQLbR4CZUAbcvqTvQaeBrrOaZ2inGARP8o
y9LNtXfqOwmq59jeJGFZZOhs+jfc1SpTjc86sPxc2ywcxxX1yd7Eakx1YDdEHupH
IOqZ29/2w0T57KezNuEpk2eZ9uz1bZVl/x83xFz6saVnae6H6H3QHVS9t4HdaiB3
bDO66V9x0fzOsX2Egh0GQRnPZCB/VzKVwyXqRUt25h+EOQlE/n3Jqn7QpNEBLI9c
Msx+GUyNtw5qtnZy65++AY6h5c8O5pX+SPQ67DiFW2Tq9R4GeOU9vPHlpQtYq4OL
1DynBjqJ8OUR6GnABXbJkpArasUxUQX8nYul8wuOsgFdUrn/Igq3tzrbQ2RI6gG/
CNBeVz4kRks6ws5AjFrb2Sm8Z29bYcPedo9XPNi8qgsW3F3qIl+PhLyNFbuSJ7UW
ToA3XJA7lmKmbJSNfu6iwzhwuoMcFwvtDiD5/YG71bR2NvYJDXYs0pSTqmfZnq4n
ZOyhDgRXdhFjV7O5vTe1ObqqFi+WxJu6iok8L8k3iPM+0U0rpe8DYzw3MA+O3BIB
sBBEGtu04utkx3PpAT9R+UZwexCSIP0WjHVzS3fYdXaqKaNFpEVFc4Ge+Qm0esZv
+iwDeRdUuZkI5ubyyNVBJ3Irvt7KbcDgzRlWAUTv9tUKV+rujuUQ07+7m5Bw7dCV
f6XU2VXYUiAM6Iu4ltj8eYidzdTu0qR437ZFM01zn/tF8Ni+SJp9iOdcY1WUsaCQ
7b247fCKVR1z7NXrzTtO9xCB0XUa13q2Ox4NzWtOihjDdEPikx6hKVdDb2Fzb8QG
qE4l1KCS2CwwwJFBtT4ghok+oOPeHTm27N81Y3LN1LsrtLiEG64TFnNDyg2rv32m
YFy4oSyL6YBhyDRDQzx7kgDF6yumSAX8oOVbxIrS8CMhc9xavD+28yZJVqW4FjXK
SePbxNZJ0KlnckyuBF7Qs50ZFcXznMgp06DBoZDGcsVys7ZWj29z1RB+391kFjxP
aapNjHjbcp6xTYI+WlLu3tLG+doGSCFpXk3Acs0drBYGVO3JjQVBFYioDIBQftGc
qtewu0x4rrHVF0+50BBDVMby48/6FwdFuw8cEvvReu1nAR5IilHWB+zN1O9bJ77U
oilwINLnMVL+JINzs8sUm0NFZWIFWdKEkS2TjriJhzvfth6tJdqYxWwR6B3qlxh5
hqciNNEYItmMhCHIUC0v5kQslXGtGY40mK++tR2cZYLPucBywNCQvjedU960t/oE
sMlquPq2zkBpY0REUSnk8/hUOjQp7FubRENCk2uoujyUKcCCLPVEw/Kkkll9OaG7
c2emuYy1bnAIJnuS1bQdCu3luxlD6jdvqQK8ygFJ5Zwl5VWXhER18oh+UkLCS4y5
E0x1RBmc3FNKQx+z9cADU30rJ0iabov6XsfG30H/2ECW+3s7E2IsuJ8lFRizFNfu
Di6Mt68tIsjgZc+z8DjTRjHo5iKO9iQmYtS4nKp1cBhibqCDslAUCvDFB9zK3xsL
pEk2FfYJc9dnhjxcO7193/KaCWgI9fUbj6o4GUUGQbHIZ+JS6DR3JSqt/FmaA1mD
9PUNGCowE0TGEWCzuXkQHVxYiEdSDDFA0X1l/1lzfU3AWgoKCRE6cZhAZ+8dEroL
0IYgIGSqv4ZwS/oLfIuwFqwTeoFwHOQ4lqbw7YD2IKYlMObBqV+NwVnIjom2dTRG
d3x1Vij07QAQcl5wtEXBX5vKtPQo4/RFLieyK8pvHdYEZjDeBJAKZFRij93PvvrG
Q+OAItKaNJpTRHzosVG+2dkDEFPMleqLt15kVcFKEApBB+SltS19vpk7X8sXNXXq
Q5j56/hoJ1j0wx359POk+Uyd4M0OJfjjpeOlo4yCdlqSXA/SvyY9eHdDfbrR+CMb
kHFx1Yj1Qn9sbH68MWSRJkNWOURbS0UiECp0Wa386h9pneUN/jvDCU2vRa/X2Jp2
p5lKH498Hb9iAnvd2bEo1m+UO9xV4UqNdQ1+QQlDQWfmRrLHexrNkv0x1Jkd3mTX
I0Obe+CIvm+aSCs34+/9fxff9ow++3tRbQA0V4raZfL2fRdOK4UrsWG1d4u6q/X9
c3F3pRSfe8/ze1iYBGxIBgtHKJnP7slRpICT32sHF8EF5liTZtJ9aOpk5Nr0jXBA
vBTN+NHvPuqxGQP83rg5eTmHmMxfxhFb2wWo0Eq3SLL6Np8kblgHGNRW5JBhhWZt
cBF7EL7xo5bhGmRSNu8+ac3xU8ZqHtWlh8bqhSyxZDBvvXtAfloHiF/XHD85K4DY
LnbvUrcyaR2jWG3ELLgYgmyfBq6Pw2nLSUVmrh/Qr+lVbGvcHT/LOB5WKDK7pg1f
y6WYMqi5qtNijrWSFz+3dbYjSKh4Ib6I1YlieVI7LF4EAaFAEbvtBRsPf8QkdLYy
XzNVHGL6lhRNUsMIOOkYSJZW+0J9ud5TU2irJHG+4OkFjnLrLFqqQrr8GGF/FYyt
LTw66LZ5FXAEFGGmrqDI88UAexeuaPLRafgD8w08sqH0lUpUGK/GrzXHsjYu8ZTI
gTqi1odIUTW5+tfaPO/Z/9dJtvwMjCzsA/1F5g9Z9fMXDlWiTRHt/vaVlOylWFgs
PXpTrT8vMxZhiyIaNfiDr5HRCsrWYE7CQPaPswQX2Yiy6UUaJpKyUBY4oX+n3KLa
AvnbjJz6MqD5vAybmaiTzjnya2Tx976QL4kA57isksgniMmpz7v4ZcY8wvEiRK/s
qX0aNH4Nsd+N2uSZDKVDWw==
--pragma protect end_data_block
--pragma protect digest_block
pj7QcqCfLicHwLtlWHjy00jo2RQ=
--pragma protect end_digest_block
--pragma protect end_protected
