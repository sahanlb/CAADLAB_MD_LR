-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vgq7xrsxfkIi2ZfEPsJlGqlaSeX/LNsxdxHQ9G91ENl/+FGM9TBycXKoDKQmmutX
v+58EOwEr6MLKBHZsQciqYnoc+/AkQU3esfIiR9gFCFVxvSlsF0EBXXbXRuhKcfF
XZgycD/GqT+whAC7HFm4Vtu6npoutVT3LwptnoIjJN/K8WMFVKcidw==
--pragma protect end_key_block
--pragma protect digest_block
nlh+CgyzAbkvZYKptg6aTZtjN9A=
--pragma protect end_digest_block
--pragma protect data_block
yrIf7QdQURPlyjWaPvkFrN8W1P5wdGchcUEVKxznesoL88jhvDAoIlLqPX/e+kZW
Dh+msMBRacViwp66cC89YeOQWNFLFKI7q2GK1ylsOEgBDU4qYzIq9W80P+NFBGdF
Qk5N/MZ9hbeuBNO5jDFAEyv4WFgXpC5b6aHZKVK9LbO+xj6aWrIeLSG40+Hqyoao
l2X3ykIlvN4xjYmb1/ahBL4ixLIIeRYSQesE4tOzGl1OKXMgzDCz1CM+osuAQgzH
L+wWre4XQV7wNw1xIiik16ZSEPUU9FqRod8GHNicy0XqnOBe4YkOcN28JQ2abIuy
F4xMAlNyyDgli8fSuS5yqN3TgeWEf1BZ8nJ1Zf5dYBiI1C/qzeoHLU8PsE8GguQA
3srrFa3QqHodWaTDEYBo3yxPgoHRCW3AEQKrUwykFHlEi8WrTpwLPBaW7SxJJiH/
PKsIIVhSR+sBZqqKspMj9NBCsRUTU6Aw0HPVI6UilfpWwF97yrT+N0xCJSTbf0mu
2R6klvy9lBlAkKudyj4velaiZH/9FDNE+Y7VOeAKTiu75WYJw9++VeCxnOsEtYiC
IaXWFdOyS8rp8ZoQqRQ7pIVgU3aS6T4lrjGhwe3TbIl4vpH+HRUXW3CLfUZOKixp
bPZFnFR07y72R0SLZJWjij/R7MyTrbRC26SGBCW5PjL9nkViTeED9isN1ivKgswj
VuyFqYWqNgZruGuYzq80sXBLDhZIRdLzQfMTCu7E3wXzq3N4BS1L0A5IR88LrK3n
qrDblAXIcJKIR1rOHxDlxt5okKa/+LwtXG+WDIKKhXKv3ges3DzF46ggzYeE4yh7
C19GSncFv9Y07BKLQKd9N6JawohCc2wm+831tYTR4waMFrIRouh2gCGoHKCRyZFP
CjLpB9LrRpQjmRdcCN8m3kmfWI2Dqn5NY1UksOOXxM9F0Hd56R8f76RjvRNJ9Tlm
+cS1Pz00xmM2rkeRsc0n6y1yQpI3gzZioCiz62kvSP0UFanABcYF2v1ZWxkKL7sh
4XVuylD3VLbDpJZ8TKWgPR9CP+a0rtrfzAUyNqbKMc2RC+aZRz3a7VQJKJc/U0KF
60KO0K6Gn5jZCkjAoQIm6kkw93jNppB1ORzZk8KkGLjM38UmqMvXz6n1ODCptJN2
5scMyAVX6On+Sh4Oqy9kwvSRR7dHtC9j4R/vg1uRKfjsboHTgmqeMwXtLcAclHyF
50MMqETaY4J102urnhx+JqI5HkHfrDs+MhoMA2vqBrOwCDUrkpJsgFuKSeKdgUbg
+Dl4grabyXXc/4sv26PJuTf8iVjJY9QPSIWl1TRQBJAq8EjmLwfLk1cKLCC9T25E
NQzskosh3tv5LYYV4INRew31mmJBzR5wNi16HD0AGP1Jo8P3wW0/4OUZkF9O0epp
GOlB4wUOaOMRD7wN8CD7aBq7JjqGOjmsjuV4ELl9IkbjWO2yWgANI9JWmdIEekAZ
dp6FxRpTKyoHtpAuIX91xAaWTrtkIyxJ3jrze5OEnwFyfsEWy3SgpyTEV0VBcTXY
a/5x9eMjDMJ9v6z0BF5j3nwkcKZUltNMbs/muK0h3EzkBgcRTRsz7hr18ghLIzEG
X1TEAA+azw82D2VareKyQFXyOsjyBagJ4ocHlvt0osl8ZjSUNeVTT3BcOPHrrDj1
eL+02Vv5afN9m+6cHMo5ZD2nwm04H69U3PLi1IMtRhQnFN1iYDOLcm60MlG5T/UH
CuP7RLrAJGN2wRy+VoVfgZ8LIEl2mKFljBgVz/gKxawDhcL3ua7h/MhG/G/b0zPT
y1FmI8dSubJIO/pa9GCByrv6ykmpCCckv8Fn6mrXxE2lmA8mJgbr06aMwvVXE2Eg
nBTMmyq2DTsEtuTy+2XL2RhK+Q4CX8rp7pxOj87aSygdUmxsbc8W3VCmqhG7UkE3
LjlptSpdGUP/SN/l4dkIt1zBs+32DTdTP3UJfh2KuO/hvObz5YJQKq/+ARfsKmDQ
YobBZBfoJCJkE/PDazIP4jktoisyhejNvz0cLjHCCoF95Ighyn9Y5vcVzSK5yBYh
Uj1lWRuOKsqmmKOsXrkVsKPB0hetH+s3gGbqZxX9/8b5WYAUCWU1i8XRs7w/71Rj
YoapPfD92DvvagrqJ0NKfoqAaecFJ+uSnKHpnOsrSMjN3wcqX414hzTyVeWJTdbE
eJd66YlI9Md4OO3EQe8zBrfvxHt1J1t+YgJF7kMtQpvOFtsQbhEhuz8b1/+o9JAM
ro3GvbiBZpIjuHOdo/rOCGULRCLd81ZcZJFvXSWaH/wyXWy1oGxLioZ9VjEIVF2k
TS70U4wkpscYscGn1PCgDrz1gv6nzEmQa/BDNQsTWdGN926700oZwn+d0B5YGBS6
/S9WEPk2FYuneM3R7IQrTBqivL6zqDRZyazRJN92/Ts4vrY9S48cygIuB5h45poC
FB3u3m688d36oY3w7HDZ97vj/IkElPaS3leW/RTwb+HgtPy1z9RUs9VM2GjlPaA2
EQYNd37LnSdwuMeYGj3+FgS9T9rMmxX39uyRSQxaPmAWvTWKgQDcZ/8EyqPkLwBm
LoAzDGPvWxUuoPQhtYj8QWiDxssF5Cdb5TxE+6sQKTZaCMgwR2+HtH8Jb2yv5qbz
U/GkYDZfpnkdZOOtAXnAI1O2O8ktiPZ274De6dqdLAQN8GL6m6/Ed2vPmqSTnkO3
93mkLAvNbAu8u+uOiMpt8Iqoth9J1+u/nHoHh1HqfAvFtBqFEkS7AktRyXSjPthW
qhSeZAsHlAmHvqVqt9B5guctrAhXBpKMlzhLzHuN0imkz4Fsj4v4KoS9I5er6htH
yGO3psZSvJb7k6Rwue08i5/dLYFp4yZlui5PjwFUiBF5oYslBIEr8rb/gE73lpyA
juUCR/KxUBnLLdN1LK0s5bD0PniRcoSgokynkGAKeNPMGGoLcAhus3NASHTBqcTY
Ij0B+Uz3qhB0hxe/ABxEBU08j/Np1d7wuUoT4Gh+0YdUmD5rXDOIreU/bY8o0oKW
bDea1arYBt0UvVtMnZM6N8regkBRNP573NGmKfW4rcdT4s/ELOsOWzoTo3Apttfl
uZhxZhFY8GntilMTCEcd7WOD4lpAtyGQUyDiWNYtT9V5tBD60D9y8Ka//oT640hm
deMLIKWf1r6rvb4S6d05hBl3GwUQj8Oj/EvyuTcr96yXTwM3VQgiz/0ACjrvIGuF
UWjtZcGtdnI02VHyOJqlNsPsuHnwL6v1ZxF0RGOVEcoNuLOk4YUoIgl9dA5wZDGM
3Mxan0MYpGCp7bvjIfafKlZP/HZ3LROV8fAgwUU1dCWIau0y43HqaagkglsmV3Gx
Z8a8oxvNj/Yrt7y8quY+ADSMLAY/5QXWSwCiUZL217c3b8blWy5GClbNqYOVFdMN
9/Z57pWrE7UPV6jMkCdE34arNykGNM10uujD9lWiC2p6vSvD3q9v0HChBzHeWyJX
GvsxxMbBhsssd1Ze6d2v2Hhv5Y24+wsB3Dpl/94X+5BlTGpaO2ws3Mprnye1fdqs
oQ6+S0RfE8FGvtVQ65NyS6RP2h9ZD+o5gxOmkqrf/0ttsaqAWEx7NSNEHhtobXpB
icTaShHR8NJdS5KmzDced4HmleFCCd1+5/obeYbOvUfeOGl3RJ+DcPL8/MgEqIw0
j+F5hm3gjIDW7OGxZ7CiwOlod63WlRn2e+p4eyMpoXIGccItXJ4VTSH5peLCCq1f
BD81puV3D/pzAnLHpzHbOrFNY3Cn/olrsdySZPPiOM7Z7gL5ByhuQTsX93MOSiJI
xvP0VGalLqb232Er5U+ikiX1aD4cxYDugtnspB4cLCRp7+T7RD9QZ2f/E9/PssnH
lVWlUZk/dgDsGFMEFT0V3X5yKaN8FFx2hFuE+K+V7RHBxG4lWCvgLExQNoOtotMz
HZfLcHbvt/hp+AeOdFcNu/AtqIb75Uiwl8X1qVCdW6Qx8nlECCQJ6/J7Or4mOhex
2e31szXiwuGYgYekfm6RkHLjqVSBIH84u3gnqhJXUIIJFTZdOOvox2cYpmyZayn6
Iot3qe2JnpaKQz/VoFeQZRukPTGepk0aIwGeUOGcfdSepj0de+UEe6dDgE6T+EBP
QSPo2AFLY9kHPu8A7IS3iL/oHl3aSS+9JxNDtAXdT2mmg9oN6s18s4T9dfqzwnf4
ij6BoYgj4HCOYYhkslCHSRhsvejG0UK2ulZQFu1hYU9i7PhTyQ+rvDEC2yj1AAE8
62URXegJaNTfO9Hu6gViqE1QycARw2ADwZqeZldLF/vhIakwfEoQuThVsmvsTkWh
nXMcuspO2ileN3daWwXlWyTfQ89ScyE5/C0XXp0Bk5iOHMpTiDEsKrmlUX5Pq8h1
8107nHYLu2t3AReFiPApTFp15ddJR4U0oz0ogSDi7UcNgjgO551F+sronR3q7CjY
U4fDQbM4qXmlDTAROzAhhMAgFae0rFbxNrriqCKzBBflsPvUVX0z5RZA/EMKu9ML
91XQn2/1jQvYU0kRwwwxGcVACWxwgv7iWeHtpq7mfytMCYFTp1FYzjciNc27fyCf
MrEOip1SbEDArCF8xjFfzMjbS7wYncGo6xDeMqFlCfELdnSt5IQgl0TzverrW/YL
qj91wXgsHI6vOaQ8MZVIZOrgUrdurNAHTlbKV6dFhZjPATiF4FAYPUto0z+O5DVi
smZyjjRCfSkxi2RsnZ0Ack3c0FVgWPId3QVIXMOou5L8uTsQNEO4cP+2JRscapnj
Zk/1yFryoKkjhXcNCa8iYqc79XqQFplYN7u3Rusb8JLJuAZ20/kVZ3IzqCIdwlMj
muQGy1IEmqfjtu2/pZal8ljOAX70DooAv+d6Bm494D5Idk+2vXcqHoTssigACzLq
YQu3u5PcoWys9043LUnO/66ZCYAephl9GIUphxmhgzagcb3QLU1KyNLi0CxciPJx
/rBYkm0hfEaEnvFjtUUeeEVYA0kkjvwtiFm1gTGWIIeDG3C5U2v1i/mJGksr9ZTl
3r7jPW+L+XR78dxFECf8LZeW3MGBj4hawyLzQTS+6lpPLGq6izvF4ZtxqOhM/I9K
SHb9pidZ+jLH7FvjaFuuY9cVFuQ1oChQ4pq7p5c2vaNLIm22pE8V+7q4EVQRSTli
o/K/39dmblUfj78rK32yjCesQbd0NRrbLLmszhlUFYkqLsXYRnhCJGcTrRdROuNc
C3fgSAVcqMTawVI7ZHlqqGVm+sxF75V0LofYYN7vAobTerHGTZ9w1yM8hdivFsnH
6j7+zLzct5nLAeg9CP95IIEIi59rpS2L22DzNfc1FUjvDyhFKFtw48giFOY4Mqx7
jesqTdN9H+CoQKXTFNFOjyUa5U0/iIBtBdukEGTONeuGHZ2ZplqhNWR6sOdngdpv
P7BRh1xfVwPU4jDeHlxNfQi17fR8IMuRXbnx/Zvd3YneXDrFy2YBe5D01H5tAAPz
gnNMIWLmBvYrg54h4UU1utx4BPgPyuWm8snhX0X2VYfBqE8WsCDMWfpN6LVQdqJm
ikaEPatiVP/OdbVdHKVs9V1kmJ1Ex5Luyq0pGyfPSXOLYij8PHaOhLKMrn7M6Hx+
jOc0tACEus95nz7461lBTeMR8GpctHGRL/rpUr9RkwSRIkrveM98Ju2r9ljZrwTp
MaQ0l347kWdQ+CjZFOGzX0kByxNpFsknZhlQGsWCy5Ylj3rpszYDx1La1C+ReHMk
5rMZshGSG49Y+9W+DVa+7BVHgwFv/7SPFQtVUXRPTloSvCo87RftfTGnv6fg4J4Y
f8QXvmikItzgAdWYV47RGgNOnMN1jOkH/+e3lvSePnv+gmoX+f+WoyGm+i7R48t9
ZkQTtmHMus23E6j1MnkD4CS44xrajJoUfMUySM3ZVvxd9glxIhCTa90QZj8kDvOP
f/yJI5v2ni7sqIGODOi/H4Tg/YAISSL8x1fDMK7ctrGeoR3T5HCCDQ224bHnH7HT
DMCbT+KRLUtyZ3Z+XYXnv54BMDJGwEZ72VXNzXD/gSLCkXb/SVeuJgqlDEdHD0Hv
udxpPhyWUWHvoy/1Ff2O1+0S62SBjTRe1z6nQ+NPv5kjQA5pEioaTPoodijT0zmc
sL3JfJriGxlbHXUAdYkS32g/iuh8p9MsY37jHjJloVcoQkS+w/YepNNbPT0dJTDo
Lp1Ww4FeBTKzFOmAcl3BcTkJHdz+d7fkNJP9ENU23M8Ml7a68r39Ed6sT3ATDhIV
1b8qvoBEzfTUl4kzArtfqVy+Zj1kPbrxTPOxjUrM/PsWlrEIgsytRkP1QeEydY+h
6Y9XF2a0ZwUEKN6kx2Byeo4YoQDRofTw0sBzBMJM4pZlvrZFT6BSGsihOI0ZLht1
siw12n/Ub0WFT7apc1tj/Vu2weO7+2TQIE37sVLVQB9eAcqAM7wulAxby+IKGmJf
xXn7qGH1SThg1k/3cFaiiWFgMy/U4LS83e55OLAfnchoKTtANkjR8Qyoem/ybVCo
Tq8ST0lOVXhI5/F/7GAoQTrBoieSFoTAxztohom+PVRnyC1r8q8xlpkmor88aTOL
cURk4EMH/UnFLxSZfVDivJLJNGyVLpmMMZwpiXzzJBBsL+baQB/A8FzZfdCaeXTJ
DrNmwVx1FZmp5WCHq5ub7wYMruKpIeRWEXAw9cepUTpLIFvzp84oOjmESax1/LQQ
rBychhpKnc+zrofCeNB9zZB43SBZsPfo2cxgAfGtzxPA289+BvZlQKxPcU9rziyu
DWbJc0kafbVCyFyRo5n99cPjdwxfeaSVTHma73FWnlL2ufk1diTeXmw042Yg6L3m
vyu+itfHKRs/+K8IHqiqj9WgkY9WBBq6+BQR8uJ5mYadICOgU8Dq8w1TQWizVDa5
9zaj34UaKXpuTPjL6482kM8uEIdnZGagcvn0N1844Y2/vqSznYE7h9C1UQe7qSpr
5GaX2jkADFtB0BcBSlN7cpJdt7N9ttHhuKGs5+ZcqDcQuJCrE7juphJZvUiyd8Xy
R7IuEZyxhAdLGPnv95vyvINHmDiE3i5BT82v8JQNlFzl5O8oiqRirj2/HoLco7Qu
g3peXKzoj2OOtCy7oImjCF0/cSSFAb1SZ96ZxUW8Kz0sL5APkgJx1JvQzk0dnOcE
8M4e8bhoybgWXcitQ3RP1dnFIsBHfN0BytaqaVbPLr8Bhz3NaQqRUj1haUtqFxJF
I96Es+MWmWav0gRxh0kLaB3n5oivlkBD7Ucp7mktLkeV66wQ6f4+LcU/m1AYty6O
MR4obKzZ7udLn42Z381rvGjrLfyFd9Do41WYVahYa16zErF8YTQzedNXc7Kc/uvI
AaENFdw1k9r47osT0TXEkIADTN6tsuLfH+t1qGxpm8IAABmn4XkRvmu1Nzc22OnB
VNZ/pXycjJD3xSgZ3kqKklNYMDGPTIprnDSE73YIvfpjB7cdS4uk99SYfCQoLTw6
z5d5HfaiexCW9VdUVqa+xpVwboytzsfa7v/lPG6KLSxR29uyD9FuzbELrdgmIH+E
+StyhoY8lA8QZsTRRxW4eP8S+HiafTie1PDfjKsQHq0xgSlRquGgVhDoL1yVxjVk
CWskGunpnU6oDPV0rGnzgh0++JbnfjFB/7j3nELwtqoxzAO8wVJJmTf2al4EFIRL
jCRyZmTn3Mb59DmGoUXSpWOtsVcGwbXfEj7Yqf7KfsGmYVpQDVzFbVq1nyzRBFhA
nFyWt4EXnTw8jFXrBwIRc0xUkP2fvIoV5wd9RSCpW9N+ZF5wu3+AgNNMeIPf2Alf
tvyQ+tdWXTO2+PLJ6hLMusHg/V8YtdicurHvltS2Mia3GxI4wTbn9qr63PR6kgn7
gi5xs2+XqirBc4z/8/sAeYH1AjGAcAYRE2BxFYy/dj43eXuOx2HNcxWiaxoCIQi6
WEY5uxhpz6CO8dBBpib8i9hrvWCkkWjx+tgeyiZStnOo6wfaLIm4gSDueJ/btpiB
NDSCibhyoHkePpKylNYuOSDk9ulwjVSAWrwmTELGDRGWFo3yDhAcye6wjxGXjnKf
1x1RC6DXea93f1WhuM8sJnaCPJr528UTFqw50xL4pei9xf5PHbMBms707U70/2Sc
D3JcOhnV7K0WZfDqrmaFueNQ5FbkCZ7Azkw+T/XjJsFz8fnIDUB9cjyGcPLWHJiw
1tkDry4YQw6FMgVZlRkEycARWLBiBAAbE3QKQ/V5D7TyWN1YVfqXKX5/ZcEt7axb
pw6fE6FQhXslpD00dQ8mzUoFrRhhyRxMxe1asXI2sUD6+2lUhJyJfNaqK/Rl+SaD
s7g2FCGcV6JkBlz2Upji2cJoJxGbSuDgforNnBtqJ8i95z32QseKFIBan2LmpIRJ
0MXP98/GRnwl807feJXn4ZcetAI1wdfm55fcpuEzo73BzrBYjkMeEJljUp12hcYH
SFwOupODJAqw5H5NFTRMPsyvCgE0XC1JtkR6L3CSZ0MvBJFKqFZMtVhzM0ZRyMNw
nUaXpezgONA5WIz6NA+crgITJprz/5C6Coj6y/neL6fdc3XH9DGuTmo5+pLcrwB3
UtuDK4qSdEu2Z9BzrTEfH6ukJuxNQ+zObmxb0VgpZEFT/dIBST+gpAbu31MSM375
kHYDRMvV1/rjONRI8CHUPcqqbJtTgXVkKaebWe2ODQHBkPVEndwzZ9qXuyJ1ii7R
1GLAb3G6egg9ts1nzdTk9xAbpahCn7LpfdFK+TjTe3YSVHy3BeVyREixTi5YWZfN
NzDm4eflT1z8pTf8ZLj86dmKZyPhL4+pWeZMd47QKzdmbf6EB/PyAfE+Vhliu+/H
w8f52XYXggY4FobHJBd/djnYTw6pOOGc5B0QqIbJWUviqBNP+gtCnWB+0VC8Nh+/
kz3BG704caw+D/itYMv/GzHpGV0jNEJwof8FFKBaCLjPFcePIES6d5VEQ2mqRkc8
P/cYE3dhkAgvEDBNZExQYWDYuuuALKGJUoa/jSLOLQDLY+6Dro78R5zi6noqfncv
6Gw1Zbib/2ciEYeuuQOAxfhEccJw4a/ugeSHCKhRpc5+hl63qm91MLZoU1IlHuHz
8oKLeFLNTMyZ+HW65NDZrKwCD7YWQoSFMOj2gECtyrHBEB8tDjxKooyZFvpRfKV0
zjxeJa2VV3ALDIrr1pSLIF+9vS2L43B1zPljGvvfZMnMaClF6vQAju6S5qwX/lwz
YN4KbrFu/S07xs2CREvG0Y2KAMNVFEeSIkls2MZloQaIaQUM//nVQ41f1i/WtGW6
2a5WYJdxeAFKU6T7oRQKZKTCscII7P+JRbIpQFGKQ1DxsOm1DPM24YFJHXkwMcbJ
abqYYR3TVm/Wjv7SR+MoV7H8QhrlJLiGHXHSID/bhN4vGZMBzeOcAD6qe3PQuPXc
1KZCQDhoCS9J9JkGKFpih4dP6ta+rPH/bPNxj+0zo0c/0MFf02A8xdMHGTyYlb4F
p3xGNGqTrHZThNs22h9kpDpZ/fj0Dct5QiH6rzh5/+tS7LRVC6zVmvCIIfMwSZ/c
/hefwhybZJA0avdm+rqJzQhu/TMpgYcf4R5TlwfsRK77QrUQI1amd9/6Yfxj3jjq
tRXW9l1M2y/Ge0KB/9ISbOJwY8rj7tC24RCPfTxLBkg4z4lF9mTW2TPteh3Dtxd6
ajmonWfc1daa1zn+90O/TbPkZw8OmurTWTHNYzVVezgaLtAAfMk2RZMOQQOsz2v4
GgkwJb+HAp4VAS3D6+R8fhUmk7OFT2QLpbkYB33S5jbLEWB1beSADbiC0iA5lR0j
cBOGa/Puh3lpOzVoErjlYv8vk4cMY4yJgBu2apO7xKD5sHvocWDPbBBaFP6hMj7j
rVTUOx3b2PjxMIN9piLyhzHM+PLRRF6fOvnmpS/My5dvUJHnldva5hZ9Fazoran1
pzn6cuZ49QBI/KyRQiaTxg5C8X/MN1i5VmnqXFKKUEJDyNWLI19MGrYWvZgEd3i8
qfm5s1lOhlrzizuH+cxY1+gptelRtuzJCOs36vi+kCDWwIcAvVW4uIScFCLenCYh
OSoRXqOhaMkHABMb5EM/YmVDEvN3sf2I+j/+kr4A8LGXkTEOib2UZ+wQweNCMj7q
4+49ezLS8ZOOi+HADvm5r1otbKIl5ASydBtRzR2IIqGCian6N09kYxwUJFyg+jJA
Y/RTrDL2cKcKeKDvJHORIT22QvufsND3/KRjhKKgeHPLq8BbyBWBwSsV0VqGSi2t
JB6dyvt3sFHUgEJa3qSbhPHQGBT7dLzGfhhfRZEcki4V8d/ewsrtBILBplzGbCfi
NgwTBLebNuiYz2FNdP3OWaPSuNwEehPQwrFnzkFHPbQYhW07v8z2uF7qeAZuQimx
3XZyiCJTHH/s7373ICL2jDL2wnZjK8TddOp1aoMvyE2q/T7TuI4WIaIlDVTOaXVr
2hHmELcXy6gxGmyC3u0PQ37lXHK0cdpr+FPoSCOXBhI4spF1iVtp0khqq9UhrWS5
Zt/pOFFNCoSn+POEpHaWuuoMejmjceHer08Kwvdq9URUsk/TAHZ3aKV1YsM1AK14
uEvn7UqCd+0jOVQSfulptwJcJYWDh1JAsqh0AFqqvOwxi6VEKQSC9SuKvCx0nhGN
WBkEuHFcAZ1ZdFMoQSmj1lnZRgeAHUbzvC72hZz9lThdxygK86bEvNLeBW6apnxx
77HpAPMv3yBYl7PcH8v4291Cr2cdiTRkAgdT3xKfJtUoIcLjMUN9qeZ0R52EmOH+
aA+FUbyyRsBJ/Qffm7UsH7iQjyNSnH9/sGCQa0RNFENmP976ZGxsLzPbDRHM4vHx
hX7awJ+4HYMcS/UWgmK3HaKrWCzQfIlMs0O3ctUL1SvGg7IeLd8QWtb+/QUBHX3E
TAzi+MG3sbqCaX77MIQScWoR2a1GBk+3SLWB8ZCVgU2vGelJuaWpm9tYTkcqeyq6
E66O71ZnNA5nO9Qp6NnjOc3OB7uj4Ldwjy3foMCT9sQOiEFwDhyEFRAl5UKbtQaF
mXTzrJT6a8Kqx0DgxX6hHbc3JNAVxMcsl7dDyCuyTnMXtSsxdhn8dwCmi8XrZPZY
tww2YWVegw34pEi7SpFFqMU3AQq1qEjUG6iq5+XxYGRjbjtQbFO4a7iVYYMqCOvY
ey1/ESQZ/ratkpDQC7fmFFfaRWsdrYS+0BQx4KgLrguLOA5weVpUxYZPsdh3XsOm
1oPz3T5nZTfZ8jmOUxUJGfQqCNztafTfV3/EnR39MVcODh4j7GwjjwS/BHy6N3HU
xb0qlFLdRJrqzcBOQz13XJL+WOKpOcNYk7RhqSKrU0PEqNvtbLA9f6kmYvoVmCsV
J02S8umCoIW7/ItlHEhWVXnI9H9OBfR2wz4dDXLWblhwaumHN8lwbYvdn6v2GZDS
q6lvUwtn54IiuYdDFbYKHBJ+BqCjzfHldRRwvLgQdOAhF5QHn9Ipl/UVe0cULFBr
p2uyrRuVlTlEkm267lo8s49Jk716WF04FPaFSqxpsMRp1LqZpjzcryd3AJ3HythE
K1hkykEIEDBZMvB71DJFUsuDGPM2iwVVoR+PmFwrUXQoBe7W4yAng5womXR+fGwK
e0UgOl77y8a6Rmtq/nPtSDmLzFpVRsFTZ4hwHRF+b9V6d0k3wuElfthsBvOkPhOD
QCxTV7HL3A4jvZl7M4MxXho07aK8KhkaqETMoAt9hHyWpmrHhDVAahxTfe7Mw66r
9u9Bqi4MhkDu2HUqmYEmQLZRGMeWrjO+bOo9VSwSdrSBXB9XAHiUw7vqvXJmh4R0
5MWsFexlHg8Q2ENbmGdhpsj1zgBFDSlcRaANfikSl5Ljc+IKhUdXiNk7msnIgatP
21z0dZur/XRESl9jPO9KowagDHffG/I1THSHHrM3DQ8oRKTmCuQYRkYHTEOfykLp
feSWZl0X+MplyA0i8OHNiitnbrhZK5aL4Yl6TePr1uF1lLqxUK4axlJgA4R31ZFB
OeDbvsFuSEvSoNNFz3lsLdDnXTAC6nEIH1QRS36dGpu689iCocm/3Hu5O++YgiUO
XuiQaL1ibfrC2Qq2KqJaXP6YTqhIbDjVSQckX1auKbaDswInyqibll5fkg0pHnu/
abcdK56DgniV/hro390lZCrj6SFB58hhKx+8/L2YB4FrFrSIseMs4dm+owgzk+rd
sJtACVYwQ8q9h+cXtFLdWUTT/NNhgLbnP20vhi3VVOBOyVAOIet7sJnPJEsK5jyk
sKH/xsvi8gbIfno1hd+TFyt9+QsB+aXKjExDgmk9Ao2J9purilZl6ki4L/KzGMH0
jqquuFIdSQBC41OsLSXdslpcwoQxmiGy9tbD3JREQvE10XYg+MCH4iJex3kqqtQ7
nxTbsU2T7CiDoCENS/wEN8sxtIaa08j0zPw7rVcmHVd3hHs1YnICb6ZB67coa+nU
OWHkpaJOK3jPa2YZI8k0n0aZHFsttdI7kaQ5Dovh+ow/1p77+VkEmrD+mX//ou6a
mZR03P5guaacrOj2JXb2MZ5bq44vjl0opCtbw/zHESyevFBdukhRXDH1hcVoe37j
zzqy3JjDeU27l6o0UQUrYpelVn8Vmn+z0d6/oucsqaVMk0cIzdYaATuh18SpEidv
3Qh0Wf2kHmpW8rn8/m9grEVNRPqt/UuNxKcfRFb3YLd1HFKbPQZS4RW9cQ3/uPft
mMAkv2dket1216GuUKu3TVuanALTBI3Ija+IVy0NfeNsb/h6t25j1OZEwMuMkXK+
k3IvS294GVKVo7iybF9iPji+gu8koh83H+dH0x/brLPQXGB1X2uRkufc+POUy+LI
fakyHWOrrM1DAiv7jL6UvxeT5i9N8LntyZR3zzMrCmStbhJXgYpv2zZ1iUErcCYa
su31KwrZHQ6uqjbKt/K+7IIW0UcXF4/qyUXJEHrcQy57IRrBZEqQdFoPEgGGBLrr
RacstweCPvORiEEHSozNp/JeAZr352Z7oFsM9JY3lmPqfCWU0GpHATGA/5a+mIHr
tXJPm2fByKChGkol4ACSV4XtUz18YJkaNKd7KTj/hc7mvfeTHSbSZ2HlYKDsVeFK
YONmGNvOHWYUFTXVfqJmDFJ4MEsc9GEUATLj59eH3U1qsZjvHsPIsLGtmEBmmd+n
ajCuhT1yGwEaLVD6zJ5iLenq9Q4/qi5JJjy/20JV8fefBR/ZqDqhCC/mrWvDUCmx
Dl7AXB+IY+fBAA4jp3guKSZuynAuK2mNArFpfcXYhCGnfz8nerqYY4T4LBktn0ut
IepuEugp+IRRP8XllOJHb5InzLuDLfS2eeHjKIsKLdpw2yiVPERZ2/pDhNkcfeJ9
HP4VGYyMAqyDS4SnhIruf9Rd65XU064A8JLYO3+0ZlGcZmLhvE8b4VjmU3ZI3WAB
rk95RQugWOIxeR+UzlIOZ50wmcJJpiJyEhrUn7rp3ohl2CojpFTnXOApJYHzbd6L
5Om++Oun0+fCY+hGGE9WLEG9JWBNzA57UulLWvO+Lvub4i1ipKeIFD8nAEmPA1Jj
ONJWNHuhDAu7K0gVfW0Rfg5i5s2s5Mj6HGx7IRajzG+ggju1GWz4HejDHucRlRjb
utw+CfhV9kbFrNPGOkznmgxByYsqOygoqjOItxIqwxwI6m94jWVJC5SLttae2P+v
2ZYrYi12eJbZMPPLjmZ+5J6VhHTjr4nZ+RQCd5rN7GxzuzECrcVRKCMAp+NaNMtZ
PW8X0Jw4gTTQm/6iwr27HeeGjXGYoFta4uRTycU57O55lq+xlVQCzbHF0zQ8s8F9
ALnwZXaIbV34JZnDyLJX93TRV6wUAFHGxhbBL4oCKv57q3OxkoCCE6HMcQ1xQd5R
F9mxzBP1hWHK6dI+XHpOLPPltmNirTIlTOaWWbzHr9tiRh3nE/oaXnhY4RFRNAMH
H49reI0t/uxl00RsFgUHbS4tLqbEU26haYIfyAE3H4bvq7ewmyg3tr5Xs9LmCBMT
kSlRpOIAUfxICGXOubwqmXJ3AqgBzkPaxl7Pszw/NlqXsE9+0mXu6e8vV8hXwLm6
3oruAy2S3FYTL+N/ETk8XHpgChKnn6OV7t5UsVs2eTXoNdjPjkeXxz818BvE+JjG
AbSjeMQRWTWcC7XyscoqW8VyWcrY+rqXhuUie6ysN3w6S5eDbrqbljsaR9FU/OaV
93Vjk6zCicuA8DPKON4JYQxwGJUlrluaLFy+QV83sNbEoi/xaITdwaPV0aKXcmHA
zYoT9vkh2rca1cEMzOIIfnzvohKHNNOeKRUY6yF+OPbGOvzVbmdikUCIySGUCWrc
5dkN8ZZ9kiYpR7aM+r4+i+inngPEjRO7kF8xVtsKWBGgbhSm9A9Pd+DZOiekPwka
PlqIgGju9DdmXIw9rkDtRYgw4W7MhbmYLforPWejKdv6wsDzCH7+FkP8tdxRKBwP
xU+XhQXN4egB/58VQ246OZCz60XA4xJaSru1i+IJMNmA4t7IJ50mU+BIXkdVy80Z
kWR2FFA2TDtNfm1X0fCUGzeFHtJ16ucTOObHzZHCvM1er4Qll8i2wzXHxIHISHip
xGHMqxf+3N0+3n1D+LZk5tidgkA9K9LTaOhdMIzmwsne31o1toJ4DSn6J1fJj8HZ
zEypFqlzqaxXE3siWbAue5Ai9RTvm5BCnifEgdeQJsU+13jTcU0WYLz9OCsAAD7i
Kz4kF1+rBMU9holOpWpz5gCHvwtEe7UB7ra1i4ypsBcr6tV/ZAKVlAWIwqvTSnWt
v85d0kds4SB9dcVf9KA5G3V5vWm6Px9yiYg33IL/59EgDmQRM8PfqmZE/QA5+q2e
kuBh8iP/icyUQZBDlw7WHZQZ1d/aYzDYJQKLJdNuKOK4q/5Yd1jjYlMbAkI6YMLZ
tIX0SsKPbtrk/9Zg0Tk5ARWKhi7MeqbhSzYrLMZCMCzzRoiVJWJZMfankSTk1fLx
41yJy4LmZJvccqMPbykWSkdhx5TTDHpQB2rQTt5pxhRMThgfNLFDJYRUmi/83vq/
MKY4z0EbpZhd2qbI3GF9X266hmLLeW8uaIJ2/Z4Htd69R/+XOOTip87XEd/n38j1
k9njbpZiKz353IQVCCs2HNzw04bdNm4nbZsF1dsJfcjrAfT4qJwvVktpHrx3HS9I
X/Qc0czQzNY1DtIEjXlL+/W+RO7kXk0fnDWCD0e2IVHy3iJeQfTRzLXuSQ6PuALo
kQMkQbxcde6VrpHvrcD5NfLdc3asWZaA8PMs70U/hFNw7QschL5kOGlCC5gagM3t
ssNHPI/XNyQfADckepMB6GBd5bZHH3EGrV/Dj++RJF9CXeARnEWaBvMgytNZO9Tm
kE7cpNbpwhKtz9Do2vNeUbaPhy9/lWoGjWT/Dv7fgyZNl3NrNY+knr8BV00uzWNr
uAv3IiIVZO+JYVTGIf5D5Zve5dxu138wUzYDjqyXWxi50/uTQ13BHwAQXMSyIAG3
LE2Uyobg2dUpyBtaixUZowt4rliKyWJBbFtM/tIVdj2RsnExv93PNDETHN9oXwGE
A3krbCe5IDMAZQfjFv3mKNFkoq2PlTKard7quoVG2b9MvIYvkMOvnNmraWpvlEmI
J7Eu4oSXErgWELAu5g4sF4wpxsGAnQs1OhezObRrmKCUFiFsws+Pc3uzRzKTIM6c
Z/P9YzM+wxWxju/xNIyC4hHxQdltgMLzAL/m5GB+wMLyGBzaMDwmiNjVQS5Fvgja
g2F8DuDOMYH1mq53FcmMLiiI/iS7nog9bZPxv0T5UQi74Cvr3L/TiLj5NBGpksXq
OqxFDfrbR5I67troOBl07Misk70DxIjMFJe2wgcybd2yFZLmzP3KoCGcneDGf2/D
c2okXYVllVyPf15ZUesJR4Bb1Gvs+2DFCVHCVnUJ618CIVsi3u5/+RFB1pKg3+By
BoeyIYm/LMfTgdOkUPBbJuzIHZqjkhdqOS8Tvxp/GmxlbshJdIT/qBeZQwJMKVVL
6kahFfIkefXveTAO/Lx7YKUepVVg7OHDrLgaXKjIDf0AxHrr1VjoPgwhULEsd2cw
4KB3Xh+fKSYmcTDuduQVdxGTTh70FVIG6PurQkYselMlgLwrqY7zAGWFtMgFUiWL
P+n2VwOhy+gTArKFBAA+xoZb9Woi+9IEJIQtxCQwK+s75OXb7hFFOcEMUUKe6TpO
+b1nzdrRT777Lq+9ZljOVzN0YjrHEdEvzx3ONLr1YD1nZ66pv7KFy4zDV7B51ZEi
PbTAbP0KMDHMtsccdahu48PHQvPRMlKPry4UOijAkz7b1bYSW5fjypBPGJFhaO59
DUTxa2DJqMKkPwCLLx4yXiPQ8f42OK4PumkBQPLXhA842PzAdHTl+6OlaBVMeOjo
H2UkhcSNMJdeqMAqiopWv8zr/HJefBqD5Oy09mPkaRrmCGAO5kU41L8ZwxFWOmCO
lv1g5e/GES6wAa06naCnsxP4ocJlWhO6yiwc7Gc6OBFTwZWQeZ7ezTP7gMCTriHY
DqM8AbSmb1A1nePcpqWr6iaM2Kt7HdPo6QLDP72Ei5F65RvgL5J5ukzek2QaiJCv
5kdiGZL+MB8mu4qXRaPeIyWGT8IZO5+0PQ0vxzHV6/Wl54J7oeHlsn06rFIZPDUY
I5DS6I5S326LdvEic8KobU1N0cJUYuGWej+tJFzhpeznv4eKht5hNvnN5HhVw7Vm
u03191Q0MKDlwFoG40jOmkSbkH7xnHgh37Bm9ZbsLZupGbB8iu7Pnq5x4dKWj/IK
lKXqjRthYhGxQIIONaj5JN7Ok4fZRRQUm1X+heo38GvHyhUTcoTTMqXiKkRG2QYt
NtlUm3JYcCBqK2K25iS/iAtAtnecaFEq2CApigMSmBlcRXf9QyU81IzzdpmnMGKC
JDrAcI7lt/yWkLIFs0eO7KmFybK9v5YkzrkU3sqA/uZeiPWJ3VY3/zLThCwsComw
t8yx+uqAWHxdqjHMYWElvX8TO2ZyJB7py5YD1bgVxDC3pWxZ4vbrLpq5Qbnil6DK
ScmwNS1N9z0KeNd61UXXsKkXI34LQP0wV85EbrLfnoHGQVk60e7EiJxaYaca06fW
6rJ8+eYt5tYsKs/4Nvf2CU36CpMJyuYAEtV7cL2aUdTL9WPT8GEstXJ6bnIsjqsQ
+A6M1jk02Be0XiLwJbG+B+cBMZhA3m7xth4bCo3NJ8AfpZKXuJ4bIK5izAfPMkZ7
+PMMIKGc88xgpGrYQv2SYL3bLVK7Rlm0atEpE1Yec85KWAm1h6t81ldwowZyE46C
HVs5lQy8B9JwqPgrH+ggjNkmsyxpghckbZ8ZG5ebzPyeP5poVaHOu3Uci4Utao/G
zcT7OgUmeMFqSMwvQJq9NCbDM1k7SiO//2IObsCMi6yzAZi61PFOobHcEbK+pEs5
FzMvxeMlbb+ETpZgVwQKlIEeX9qZ8Yk/injbOjmBfmIEy7r89d5BViO5qSZ4Lfnx
GwZhOfqMmPqgxsxmu9GBgg/0YXq2ypwSpkADnptP2wmGKuERpuOaZQyIzKBCj44g
CnvCxNHosgtXrYLSBuEj5xuZrs7sBFjVfOMY09xLpdQ3nbWqDh1ZRS7Ir12rFOmd
eZRHQFDPiatV8sTM0WfBXcapJKUN2aPaWRBU2W2dmmxflZTKTei2a9QaQXFcr27Q
e7MGJzyvzJ7vDWeiaYJZ6fUsyaiPbk3VcOb1ffeCr3RABofhpV+761nyA7oikp4q
5mcaEMPZVuQd/wBlX6JWGcRbkEQjr4j8iXIMzASiiSQI84XMiWWRKoDfrCiI3ER+
ss4AI7z5aAB+Aq54Yw7xl9RvFz5SZVDBaDvvKNjVc/go9lL63SIkPbvNdo1mPQRu
iPltPtlrwPLKlq9YWzKCCzm6134W3RJ+FK1/+Qd4S39ObNx59hzDYMY18mwOU40m
pilCBjpQfDvc1/vvvPlRBxP3xxiJBxVw53uZM8xnR2J7TMOExqzM5+KBkkJlgGUr
um43yc4Zqf7+r5m5DF+hXdxDCmfu1oe3Ujiubw4+lJpYFWl07FUzdB762YJOF49z
uwyjFbsZfeXIZ9NffL1YFxaBP0XhAZ5M1wrCNjXmpAhyghYx79YXddFjhVqsWqU9
AIFYTau20IqK3YENaj+IQnBBhNIYvYkjAXNav3P2nkKTI4Z1zIy7CnH44wbWqDHi
jQG2U+IFB/Agwe5a+XG7dA1Dk8/Dg1ElBXpVTrB+DC/J9Q2m132UIfyXUXgsdiO4
VXaXSXowucZAR8PYq3n4CLn0jUcm7FuevOInFf4t4YBFbHZdkmesTdCXTXKJ9XSj
ZG0oezZO602aNzHNzhyD+mO6xEZxUKsu+awlVo5U13u4X6oMFWX7I/DM0iD+Pz47
vuuQ53AAjT5bsLJkVobHHC+I3GSYt2enj1QNApCspTB+7IPi+B5GmxmuZT2TDNXV
f9VEtR8sAJzwPiQn18O/dvofaUEFBrgSEF6ZLgdfRD3QL1gzopwzy4jtGm5oMiF5
PNA+pvPisELmpT5tQbHR4risN5K4QL47BsM9q92Ub461+b+H58jUx/SXdGH8QhBV
uMDuyREvB8TlPb7L4fmKnaT8JX4CuH/7YZrNLBFhGEEk2tp2nkzC0Jo2gt2ll4/T
CkYqByNbMoHWI+UvJEiNZl49ZQhW6yfNX/SBQ7ksf/+r+jbo42I3wUqnxjkeFEl/
Egjge79YV96oaKjt6m6eNrGMOwoRwS5Gl2a60HdE+s6FtxI+GtCDL3NejHc7fmIi
2YPbOpClrLzhSG9YtMU+GUZd4H+Ni9mHGcmgk9B+9439QJoC8KumiyClPD4KpItl
dW6wDEa4ptHZvDPgeLO7r5Nbstr+Ld+jV/4mNQau++iDVTdzlM8/WUuuKWL3I66u
sGsKHhQzMCNoLHPV1Xt63LRCWh3M2UZsF8jk0Ttu1yXwiTDMZwhaZ9SDOev9sE7c
ojH4N+PwMw682OjSbj1X6Fz6fdbIBsWy3puL5ZHdkYrHdGIN3wo1xnAZIdiEPe/8
CsyIfeQhnPf1SIsKZY2fextxXMgLSGysO3bAGDE6SNTBrMn7YATMto1RNrNySEAV
bbhfusp6e0PsA67e8d0Auev1KZ0kKIx/8RkdFRj0pvJDfVHiK/sZclIH/gxLs0Hq
sP1ecKiDOEQp1eiFzcQKldy0GxloL8O2UDu82gB68HEpIbX9w5jPKuC/xV42GE//
jcECSpOA6gZ6/iek48Ia4M853ffAeCqCaK/7BSsVS5I2ZBSGMDvix+O1qZFj6Kc1
rwaVPnUkPnCsLyMz9EAHFPkkJ3B5uHhykuzH7azm3sFUG4u4RgiFQDY2p/Z/2Qdb
t/Flx7n6UYtAw4gQMWTzJc1l2ua/4XUIvApaTG3U/pu3bs3ciO6UWprcjGdY5ItR
R81pqqXdNfsCuGkL3DxS92VLwetQFfUl8ZXh8cRsZCIfM+ZzZFw/e6frmM8s8RbK
zHnn1LpAXeM0n9iNgeaqO88w+OAALMfv2glEFBd+MQPIxCvEmB8Z5ULaxQZFj37s
GKT2rVlm9CKw/mJzjTvAplbWWoz4um/2XrvXmBmmpS6hKVl5zT3T+qcj6TYLLOxB
SxEMulhnBt0ZEi4NrmJClE3HN8MRanIaaVZiPFe63QqcSJl+b+K4MLrtA0CcZAXC
zIyIu5PIn63TXnvrXNKe2LDuXR/DK1TdRs1W21P7MMsj1cvRQWssNlWrK1NXCbS0
6rC/o7G+TqRphqudBP/GN9Y/sACx6HMMC9N9+6sLRUB5rhUAWYTE3WEmW30fHkn+
r+7UVAmPXXs/HCycXWlstUOApV1ZKlZNefUTMW2QqIAtI0tqwJUnvb8/JqZ/AK75
X1eP2QyzvBgJtj6w6bk7jwdybLA3Cs/WSYkZIrKhsXHQlwDVcHRnxWVBMfK4tBSA
qWhQpj54wZihJ3Y8sD2hIqbVZ/A6274SVOYZsmhlWWpk35bl0maU1FIrbgKHojky
2O1aTPG8h9qd4yRIMIlDoehOMar01KHAbj9S1iYg7+j3LXfX2dqNm7ihKY2rup7f
deMDsyrbwVrj49e6tZyNj5qRaDWzbpKVf39D713Y0M5lFw1emHiuUs3MJRrQ7uOk
A57l3e0GJ/To6FClBIoNQHZLrGc9b4EnzPNa5evFty5JHM2AopugC4zYu/xJrWPr
mm3rOv/B6EN0CDHXQGrHZRo+/SiGqJ5bEu35+/F3AX4Gz3dmoCdod5oP4pr+XzVl
TehWC/ac+95X58nOrU+xGEsSFZBp+cLtQ2YI4+BAZ7c+QMyzLmSTSbE8Zd5jQ4Ma
QGeVQnAQiHLCGMusBdKaXKQTBGYJ5y8RdRfjSZuZgD7oNPUMoBWxgk7w0XvxWNA0
8ihOK8TGer79s2NItjbF5NjHU3tCIoCIEwl3o+VGBdJCTFEZVyqeq4gq6bcztyAQ
PRpcvNQ5JD9gsxiP+AimyKdMHdpP+KRA+igdI5HwbYiR28sm+h/Aiurfep7eQi2V
gdSRnaUL4hJPxGOszLyKj6zPY2mNX0OHUplFOG/U0AwX1sUlfo6YvEo0ixwgcb/H
sc+l2qu/0OcntV7pGe3ZgBRkE+HgSssxMjVato7AlRCu/f5LFTAQrvI2yX0kFgpW
DFApropKzxi2H+ASKIKcHR1VkKVd4xRQXaOoG2YEJA1grJyL8CiEI1XnVDS26yXx
8X1XlhzhDTmlwcDwgRWJa1wAnFDgjpBvvFASv+K8PEKI9usARbrBTWCi5B+KW8cK
2lnwmZlbcglaqf/qOyy1rWOsPqsXLlj6B2aknhv6HLEBxHXaHS66l6lwnMT5yUUP
V3FfWx1qekPoG53JPW+RpxfLOtDGXnllZaa/3GsYvRzSZ++eRhKWCmLDQZ2sGQkV
umM0qdDFwDpzeW3aPkCfozUYnsrkcnCQ3LLIi3O4JZHZDNnA8qOgWK3Pz6QSLHOO
5Ddmv+WvNJHgfehZEL3s709h9IzsQzx03jjAYhHI63v+dM3m4csEaYUUZIimkYPx
jQOUJzbKKo4aopP3sLAWE5hA3GiSuy+BVvZIrZkLIdIDr59D4fbZ/N9s9JNVc0L4
zp/KqxVJ/kmQ8YqNjVW1j+a49j7yWQoZtp8yaKpdOvijVQqAfybZaq0QsVYm98Th
94VRaN8zhCdZ5q/4n7npnyzQBvODHIovFwigE2GiPS/u+G6fXrRAzT+IlRlz4Shy
0EZdsodUJYmCUC8708Mo2tAPX8RYsunOoro59gihm/V03kTemfF9V1ExWocSiEtU
zEdSDps5K3E0RJjBGnokD3WphYPQO7g92AZaER4t1E+jdXrtWvWeJ3AAR+M67cJK
e2GkXe7gP4fPY0Kc6RYNtrdOZsQU1pZo7n0kF+fzwfi85TwvjueSByjU7RJtmZMN
/ss8blpm1ZVoWZT/hYkl2bFmOnBwsHBUO2peKjkSXN9LTc8Qd8+U6orp1VH1JvYN
l3VRq2rEzQjI1m6uqnjZtgcISUwCUz52lfLsrIaY+IMGRuhuU5W9pTQagQm4UWA4
Fp/NZLdWHcp8Z9TmxFhyhQ0Wi9ZTQCoAreTaNXoD1SyoxbQhpqrKOIAzNbhuV9Hv
NDKakajlDuCsDFIY5P/NxoAaPN3g83YkVl/tVB+awKmFcCg9c5SvmqxagBiCutjL
KvAhCYss9/AQ1kjlyI33P9NLqzCnzfWLQaxhnyuJuOeQ2h69nxH4//07rI0Vw/uF
oFWS5Ua8ziXhIypPS6KQ0RCr1dWXgsp2ZTwHxAmMKkHPjt5pYH8vEgc63TgRk1Mc
W0xUCZlrWXliy6LZpqyGCp36qVBdulMSg2U94LA+bq1s56KQApojCyu3Jt67MCOI
Cgz+zEaNkkdFHB385tbUB9NQVf0Lfpl8MbSHIs0LXxJLCzjZRU9wgJtoDqEDpjf/
rfCs5L60k4VNaY1SDhs+4ph3ZfeCCOydkYB2XQw7ccynEkfLZFaKniuTGL8PySP9
JzwsbOoyiIdCXgasvUnTWfxgjpncEscTwRQIGlbDQiB32NmnsL9HgCZ9ZM/yHe0v
EdiQXuYn+H0LMv87fcrEAMWAClEHI6xCqZUPlgpomOnXQ60VhjhpK1v5bW39ncQA
SrDVrgoTmUfwjSVg6T4KfhtuoA/QZJK5Wy//J2RFDIhacJMgVMizG6dVUW1brM/q
I2Il4wKbKDRtTmMBvDkA8UKGR7DEes2+B5y1noV3wYTNGh65Lk2q5s3ciqZim69o
ImeOn3+INRuRI4XseHuFBHo9ger8vkdFMEfWTckKlqnSb0Lxdfvx20DSpnB1gbjt
UqIEsje70KtNZnfx5gdvDBlqHir2NsfgeAqa+cbgs8aDv8QppiDBpwjY0hPiFYzl
AZIrvbR+eFFI3UZhkPukUtruRlM/Zbc1mQ2avz+my0u8Vg19jaPwJejstg/9xlkE
bETzg73sunb+r9srL/1pcbPkpI8YKXOTT95Epl8t/JZ+VUEGSRjXQDurI4O9H+sZ
LrOmRjZJ3xQaVzeNb22uM3oVJR7WNcVrt0Kn1ETaQfPamDS2qBidXB/rN033waW8
eroP4ySnc7be/eek8XM8bmoLAkHtjcediD7Wj45n+DWsuPdQ2x4W13awoa7o7fhr
IMjk/xbwDd64x0HxsZm4zxmuIUN3iRGWLiGf/8YE7e+a5hj1Y+YfjJhxYWoKDxvb
Po+ODFr3rJWnGjc9fyKTPaPzYOv5AiYGKW+E7wFtSTfg5O3y4wHyqDnq0aILi+gc
dfNLIVpM3tnVN2E1MX5B6XxncEBS+7yMHa+ovwpGB3YBsqxbfnEuC1vEb/CMDczL
n5k758ilMkcj7ReWd5ldXUJ+09AUqq1jse9Q1v45HcDHHD3jY3NPRv0A+VT0dHRq
WfypVgBYocNK61kD4ankeuirjMGZrLQ3HchWUA+2Pqqe4r/qIPVRhEu3g6otCBR/
OiRxHiiz/QOC8qBQD0CZYAWObBZJFXNLK4o+4OqUvx7NrrXUwb7v0OOX1vZSj5tO
OzItRcfc3mKHOIxen5x2dtb2CH+fsIb/wALHr4kJEC1HlZtl3SN0QivkpytTnEtA
z4EMj7nQLrxbnjFy37rqGK7Ur/P8OYPPNHGkUPQ+Y1YvOp5yZo6Aw0DZM7ay9GBt
tGAoG/1cCUmneknjnMzfxl3Al41Wmwk0dMUM5w+hIjJKhS2nzp6fOmO+tDaWa8Cb
5OEoBst2lPrIEjnI40buaMkKs0+JVcbOUdZYFfJbHrOYK+/IffUtrdbMwZoG4uCf
xz3KKpfbMAzPLbpZgj4hEt0KNWO8v0cO6bDJ5JfXX4jqODfuihyZjxbCydX5KEnf
ruDbmytW2NfeM6/8vDDeqV5ow9/UJSpW8aQsoq1B523L70jSxYlxO4gpQXLSmHXU
x8S5AGM35j61NzxMMqFgAaqydMW7pnUYHk4G1d5OxiGiOatLJol4eJ4aF3TjpP8p
m3qLFEu0nXPhCzO4qBhK8wZmcGDSWchIj6Y3gG/JNz3e1GJGkfXuUhFSJWG+sbQW
im8c091QmnCA5kbQCR2bki5WprTK1u/tg514oq9WTcncbPjkmLPxXFMhjJSTQgpn
MEc1uBZECttozFAtNMEPNNsvnHgC3beeUbycLXo2fu72TNd073resqrzMdmaFutI
LHGMjQMAvIuoXqE4nGyEyMcxStFFLdEWHxBeDNSl2HrWbJQ/14K9t/xXr31w0cwK
hWqbTWKcb839qBEty/0O+MDqBx3d6lBWKABrRGL/KAGx45ozacNl48LcSjNagbcc
dUsz0T5rZ+ep0vA08vhvw61psyQwanI6e2zarMzw25V4c40D25eMz9+LditWPXlV
KUD0U/WHmrOk1dpzUfdZrNOSngsPUpfQ0bsvmXxeBFdTAVZMDNFfiQJRLTEZ3TN+
IYT+9qkdKDxuj99CvK5byB3XVArvOI0p/OHXkPKGFAhAa23gjQd/bwE+Nhlf8fQl
MyJX0s/ylXTxNvWdbOVO7km8Z2AJ7/YZ0mytX/pKRt2h3UJ2+UCyQ/z362IiB35A
R56Xhzdf1hY/CdvyRz49x/cj/xvgWzoX6wGfUDLRJhg66FEec3BEtK6zRBd+ZPek
P5tXzEnYSvfce2SuptMkNIUNvdSrEQZaSyG+mGuBdFq9PA1JBbNEAWxYKb0mqyKM
dKz76bVz6x/xphR5mNQckF0yxLQKP6VqSW3HU5YCiwSf8VEoLcnoqvCwDX2ZaKEL
/8L4eB2c1B5XMW7AJthxqP4ecndEgYSriRBa+HdrRkhv8R1QsH9SKtMJyP2BVseH
wYfvPo+1h4inImvHZIKrIhYwAiYbAg8LrTog1co+Tsw8IUGQfYH7ABzvREC27G7E
o0RMztZIObioO9oZStoKXgIl3+4qmBj4qT5/pXvrC6xonWkei7ruZcBSnyQL2rxJ
tAnucEnrz1BeJjDTu7uk1tWErsQmWf3B8v3FErjv4GXaq2qjljLVJEEZp51m1sHt
jtTuH84pfHx4fd2vR5kjvjzo3c/+4WzD1ueu/SeTmTR50HccfuRUqiMbWUouiFlb
UIpI8TtiqEW3hXthWJcBhdmW846v/qoEuN3ojSek9rjur+54CGUazoho7NT3cMlk
NKAB/loqcS8+HI21sURwaLtU75V79FqtyJ5WdiQj0FVbi4uQrvvvHCbaVdMOop8h
3HHUTrVrUuhqTBprn75abIGxGMmk87uU6jg4joGlU88YxP4XvMjNYTz27QTIgpKW
hAYBwzM3EsS9wb6/imIlrAH85A+f4SyR8hbA4+ZzgWLL14lvN4n07rVJEiypfgqB
SbZp+GaI0OEq31MGhSAaXpxSOx/GHBzVvHkKV8cE0+cP1WdVDciPekXUOTeWz8Ie
9SUY7GMgmg2G1EkzUKyFnwP/eGraH2Cc8b+XYMJnYZ9Uf2T9k1ZO2VKjSPETMECW
pKjhtV987gSJL3ANARcBO8/G1y4zWzzNYsRYluZYuSFJnT6dC219o8y6L0qI1sc5
zZ20v/qyUpAaS/ztyq2lABxaiyBoqJAuabS7wK+gE7/ka7vSHOxYjPQrqq7K6B2Z
5d4vrjn2ZeH6n0Xj3Z0WitwSfWsTjW4T7pUzPGpYBOW8ujY3f/BVqvMdrcsyegq2
5l43O+H5GWIquWyz1I7uMYsowCIa3cAsQLyRea6c0DhSmhivDlI3YwIK0gMt1Kri
3uQPkN8TvKrhklocPspKoaJLgY+u3g1MqdMK2wv2pNK9RSgu740ZPjg7sZc0PvqM
2BTwDWtkMY2/bp7uxphh/1rtq2fKZDeVZg/j8znmnacyRvuj0QieivotxsV5Pktf
VIxSe8SZKbFSF87nFKK0V3K+LCyNttqd89MTAPlz8yukTtYmxIsz3i9Dz7oeXAjG
JOrs4IHrg1kI/O+ywHSCLUO9Ie+QyfzOP4mnWVoT++7RRc2FfNsGWcz8b6tZ+719
LkbuPdJEYGN0ihnOPQSdPBjr8ypWmw+CD2ivanGM81M9K6E1gMKoicwMggSXkk0j
UAzd9M7UEclpnNDidBtBo81pcXojAS9lyQZjRFjU39/MvdnlUzb/EJk72sp14uUv
hm3t8W9sU/XaEAeCWpvvNuVEJTF0HmhTuQ0z/4PV7ygYFVCbgTfIPE/4O+21f69L
p0hv42qHz8gu6TX0fk4pQi8LCYScOXiYkLw5QLuvsO/Y9qbbbS+5NStv/PcNJGmr
tzBloEx1y3qcKpRkhfaGQH9JKKPCIHibI5cET6KKRLgDL+1qTW5iR9N4lH7c/UGV
/4T4hwRCV7p1ijgw1l58FMLYwM+L817EoonwHItdHo5F23w9O5IeY8ltmxTSRlVe
pQxU1vgbwfrxBekTPjoeUMEskhuahWbzCG0uS7fXOFLLdGOo070+OqwPZrN3oWVy
W3DSYD3+ALpgPicMrfNN4SK9PJrndGIUkLfWtKSSjA0iN3zLr2XKlntNjrgLntIP
OdlAOaS7l303KkCq4tMUjPn+J6vmoJ3qBCivhlCigLaptFJk9JBbLq2V7h+PQ4ec
FyMHhBThQv+CMKRXX0q+gLeU7p/yNfn7jxCaZLJw5mf4LJFqWfXHXSBXjBy9QZCb
K4r+Z5A8LZ/JTHJOGEeqR363wUHoFPnW8NZFU3qHdkc3UPAbLwF73B0EXvzD4V7w
QeiAr4x10m6NcUG6vriu/pOuTmF/h5E8GzSmt86Z9+fnU2ZRxVJZHQZueu86wKKJ
8PGFFL/KIazmqmwaUHes2zqp/h9OnLtnrQcyw60d0pqSHNC9H27sDLxEIYYOCe8f
yoe5BFN5RBY8C3s6neRAsG9A+7WYO2j2r+6l+ic1NJH5kunrEdGJC4barAJfysso
6rsHIfTN2b9FKI1NZL4//NIsJTtNsu0xjdgXQ3/6DlvIdZINqAME9rvM1uNfoQHn
oCHVl8BwRLn8ngsCzx70OLEO43xs6MKFdtolat9C0/tUafR8uDXmMafRnFOrbr7a
ZLEdPbkS7EPl8RZeodLOL7l0cefyv1aJ7Xbg1Et/gqyqL1wWjMIQ4eC8exaSQt1E
6pwdqn1/9CdBTMfWPdM737zr96/96mYazvub99M6BpxPMZbddnvCn868WBqB2BfT
tYAM/2vJ/+YafDyDcHQSXxEhoB+/bgrxRz7tJPBhf2uk3Tjlflg2T5G43XtqwG6c
5drl19DAsRWa7rwt8N+GY7ddsNw92vgifbrkqO6FYz7wqCdFWPdm0NELg8QyaRir
3gAw4AgDwx5kqq0bTdchITeUGLs3hGOLUis86dVU5TRecaDybdQvm0188z6fZyv4

--pragma protect end_data_block
--pragma protect digest_block
2cRBd6a4IbDg889kp6jUkYnEEeM=
--pragma protect end_digest_block
--pragma protect end_protected
