-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
myO7W82JkmkTzsn76l4o4q2rsil5X/KbIFBzRJkPSDjZ9lKjQd1CBs7Xdi48Oyrf
um6zU3jGHUfbZrKOf40JguQImD0FKPcQSJ7uTFo6EMOVHWll2LClbiAAYxxqtzGD
PNmMN14McWUKEGu7Wtil6HIJqXiBR6h5BNMsc+5Jh0o=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 21381)

`protect DATA_BLOCK
xoeYYy9TG4CiT3z3oH8tGvbWdl+e7U54O3tpMsmBP6wBwKlGZkLTitL/Cd0j7uAl
VDD9bxHGpGR7Bm5e+/N8UoKWzFO7KASf9F+/1VldffSEZJFf0q2TF8lptVLIDUqc
ghMifwFjRme5INHvgC0Fl97B994wST88UzIUO9Lc2HZZ5wiGBLHcdJY4SvTOlj1K
SVgUx5itj+cEQIVt+AwNPAz1EWzJHioQ/miE1xpLpBalBU8Gm2bzyvADNqgihDfk
b8ngg8lX5T4J9CdzC/hKXU+DkAC0mJfpqygQaDHX42b0s3oBD4e9kjq+lQamilaj
kxnY88TCZTRHpwvhMItYC4ClfngPyejMiCuDvOC3YPZcHahS80kP9kZrgDIhNaU9
tcIn2aqSJBy0Ueimivhi6GS+5cY3DZIlZexVdIaGsEFai6KVOKfT3AjwY94uAEGP
+cOGw2bZnNIa4drsPX8LpLelt+mLzwM/e+ohyOnALomL7NkmlXpbY314r2ocflfE
FD7uo02K9kPH1XUOVpdW4vCVoNMvO8GTSwbaXLCaLyyYGFKSJAntI6lM/nFtDAKu
RBse7s1skai9Y2nBGN526ZusOJZRpxR/deWwzCttPf1Okyeae+KRKk1jgQ3Rag9K
jiCYADHDcm9prrtGfchkHrvOXKyBtpGvS+/XVZkxDcYmrnVCDBkZmCMsKjgsFxw5
tomfQ3NEnelfLf4FrBSXRFD2hz1d7B4ZDRh0HjytKG0WankQi1jwup90qlAMLjAs
XQhzwBnPQNMwtmSM8H2ig429nXXnRwQ1uYczbU0iumGbxhC/h1HtXqalu0vzJLsl
j9UOsOMI2T5r8lF8Oz5g/P0H4Slx5FknF17EQoENbZ6MohII4JZVhA5rCoinn0hz
PKk1kCNziR+KN+/4AhWrZA2Ve7dMiWlDdctvtGc1zAEGdiX1yk+v585JQOCGyx4Z
Vx9nEbnaDgmryRqrXbJgoE0b0TCYi5Ho9CHdVSG+lX4VwVtGsrfzSbd6JWzqfDAw
JIFUmN29lNXEEjqGHh8e7ufMEqkjqhAKjudEN0pmvJwUc+LzOBN4rE2QQjGaO6bN
lv7iuFUVMDtdel6gs9ViRKXqpk3MpGldoKaGbyjw/jPEtBZYnwmKWWZMKAeFUmbl
UQ1OXSDk5nD4EiSnVYAaN+eDbyWiLh1ELaoMbQ8oUfyvzxz3moVu8iUBCfKUE/kQ
+qDe/c1c9I8FzedZMkOKSg1NSuNAc4DT4mBz6Dxb6k9f8WLkMvudgQglMn5k+uEY
ALbeWeke7QKVKmLAZEJyfm7yozY8NWoUiKLQRXk0UNExSlTAEm0GU79FpgHA4Qdh
QDB9+tod8oAUVooFTCNnTGWTNEZ7WCOKTguf50DyX9OLbLXaldccIF95bUcE36XG
MtAx/gh+PA8XPS50CFshlq7NoCD5rMg3/lx6Gm72B0cvxAnpP9D8OwLYpMnQ+Suh
T5DA84Tr7pIgK8b8AK6EaMubK4uWkobz1tLaHwP3XRAVHHJExHfaCQT63nuAmfdB
605CWX6WwbLltsNLYt7ZGnTQCX2W6mcBDniu4iAwiuDzQcauakb34IGFc+rcwBwK
ZQHIUZmJDP1GDJ/bEW3cEjdvRrpabxTT/wTpGqDYBRr3yjQ3jHQJYkeuueJovi5U
pw/anjzogtmwLpGKjCvuL6SkIRhO4QfGLBVEvP/YBZ6KLsMYJmkeP688c8/zlkem
Oyq4JlIlU7kG6P6u0U/6d5Adeki2g8Q6O4rwh/EgkUrQWz2Mv0lAayoJfVHzw9Xv
h3LBJPJ8i3Ri/SRej/LDJaE63NZrxYW/sgRnwG/P3ZjWP8fWSTKNpbknnr19xydt
dB4ctaf8+q2HTiE/xaChJrSb7ew0V/PaC+acH4Hmz6u2WjjN58UZ+4gos9psVtPh
sxPPv738sB50B/dIaMN4B0fCIqdIOtfDGUXQ6AGJu/vuk4fc8WRH7N7wWJGU8RT/
TgQaGrtDv9O2pA7xkSwBhxQTlZm6ePJ+8Dm0g23hQSatwTAfDBO4zcx8Pj84xviD
VBLDIZO2urFA3Dh9LEbpBT2SdmVAaOyVY88MN2yCK768vdqnVi/l/oP8dcCQbBXl
GYfURX+ha9BWc0sG2jqAFb+gAHKCiD4urrEaCHr9ClwlsdqYcv+LAd+XDiC7HKG4
tqpwc0HUgVFqRXZlM/a53aPyl+byidbIv1cUY9OCiP7P/9+NhenDD4r8DuAEUVt6
yzyhH8A+jPbzjhucM4dedQE8HxpgvsmHRVZNoqe5YhtpTDuYYS4L1cGMZrLY/3vH
2fFhIXA++tNK+F6wxYGx9htda9NmDW3SU8gWKBpkNtrGr07JTw2cki3XzszzXGUp
A7OvQSWrMsWaTliwhN9zJ/kRzWY7Nwm51pAPiuy5E4VYaCyATS2Zg2ErJH9tt8VE
6xT2S+MttRJrKxn3Qe6IraQJ278Isj7OL269yblEA2gyhmRjqV+OoaXUfhdmFOmY
zEAmCav8fsuoLcXf6G+g4VipE8qu4WZ8OD7da4dAhqWxqRiWhk/QCVd3D3C0B1aG
ZBfZ+G+ZxmLNYJazXb5PXYmGoHQ6iFxhhP/Hxwq2m0+DXKGuNxpKClCMXfI39iEf
jqjlzLCJrHxvyaoFHt5MewxbpIiQQWlaFJfc2L2g244gwxn35nAyGfmqKawOyHN8
NF2PEykMjSQm3wqHtx27wk2JGupKjLhLjWqVr97BX4cmitvrIVxVHru5tFnjrEcp
/X3Z/QPD2sebrYnJG6iSub0bZwT2H9FxYNj62n/Hy0nevTO58DUGdHdIqNJ5pknq
4vl7nWeQOCiyq3W9qN9XR/plyovcL5rsle7rUQfUq7MUks/emZ60e0M2UpenxDWP
G1A5dGgfGprHBAqr2egO7+g3zzaC2vfabEmmpwqqJijsZ3gn8CINlB+ZzD/8WE/4
hlJDl65KCfdG34gCOp892+iutCPuo2o/3lj1Awy65DXzhpRfVbm+pD0LDaibwt5x
fj4h5sEmHJZUgE41X2DwwLtKbI/DtV6eVsr9C675/uhIlhKV+TiP5qy7JniKBQax
bd43UG6XcVvX8W7qFv3uOKnvODAZ/6RnV6uh/eDrX7lUCq2KroMIaGU8lXolm4vz
FLOWDDy9fbNbg5NJ++g2LEvWZWkQtE3J05sq2X+YF03UIvutWTJXPncqT1rH2+6v
UCP/v5MqNEm09dFWf9W5wMIJIw4xut//sGDx7fZ0vDmelZQxLkpkp3Pcn+zcQIEL
Y+B4RO5hKj67uSkXZydKCzbzSBmHXzW0IdU/35gH3dITMCi3g7FDO69i6NqFUlnF
IIy/jZOT4mVhQwG9tC22mZ98VPsqj8or0hAKO810y9E025DZVEntwCSzIpQtDYy7
Zvq5axEHXy8PDj9Nk+22n1GuklPvqgGb1Pj87y3bIENcRhnZO5AQxNUltqKjY+cL
xA4MWdFK0wqKPmnLSiyZCDmqyhnugnbH2rBCIUB7LKh5Oh5+k6ReVRf5emgpdEiT
FhW2CGCy1AydJGa5aABrtR70JClTDP5h0NgcXzuYzfu2uWbXpZr5DC48wL1/ktpP
6mk7gy9SFKDaxwllu1BhZNUA+9Ls4egAvvZEY0oVTcgBEJKMhUVRCjwbKKOEB11b
LeL4t/kDISKmgvUq6C6eN/XOJRlzDKdvgKanVvwH1dJ1YtBK3aijdB9WvcpGAsBl
yEO1/jggh4S/wz1zdkofGlBNAnAuJUN58wBjt70QUtTrhLIbEps8mQzfgjjB+No/
VSEZSL+qAZIWjpoSpvAPECSinlyu7D0UBo8dMmFiOuqTpOmX2EQSFZcOB6CL5cSV
U5oyVDGA/lRzyocciKVM9C51tIy5DiT9f+1zwnvCBc3WPfVm8nYawDzk1Vz9B79T
oyzRTAyGFzMYPjdqYrkOfTZi/1XI4k6YMJtchnybhNJqImfb8x0ZhE/LMtGHb4si
/M3PxNJzFu0uVSieeLZqquAU+/u3KMXmOG8DyZ0M5MjHknvYx1jeTm/BLeA4jN4v
7Y9l7EMP3JizYmBuL/HTYRZdJabJcU7g6HNMn4gflwKx8EgtyypSF8m828JzxR7K
Jl7+uuPTByu5W9zIvo4AuKu/BC7CaxJRieiendcVFXcO16qMyBsyO8Skr8biR3MI
E9Pzg96k4lLVdhXnY7VO8SkQBFHv802fe1w9hTvVrcMAFC1EydURcUqfQiZOceOQ
BW50jDCiRVFYtl7mdiEl/b/ZIwESw1tm3+6kltfdGaN5UXOh/PUa9xB5+AkUhrMQ
uiALyp5N5N7zG6lKd/CvRYeFV54ZZvY3zET/Ht4CJNQ6RlXJ9TYXQubPZ8iA6iFy
xPvccW5Jfykzsv8B5n6cLptbIkJdkSv9knAtR8Lmsi5sihSNtRF/2qpNJy413if1
WSSFOHPzgbHmifWwSz5787L4JpU8BUJRNktaYHBdjuw37Zd7/MfEEqEHoUIWbb44
AzprFN2jERYGMc+T7fIfxPh3lqySUGBBlSTLnhptR83eC9PwVnY4SzkhHQU2ubmX
u7z6iq/6LwWFjdgO5LA9GK+fYdWfDHTugNDcoI3BGck5th0IGU136IaiMZI9AEQx
uCB8/geJvBoZNJsJlyXvOkMi1/58dIcDguFeIFy8stPwgaO92KShERyYIeEMThyk
e5qs4bb7yvUTIKleGELcgnwFur4cHnrZXoVKbHXNMqzWWkgjGWn01WKoUm8Pm9p3
/KNlY0ZHoRSWKGKVdV7mNBdQzWGKVe1dlL5QGqJorAgwJR3boMq7Ez9Iz3zl+XrD
23LplZz749mtk6OCOeUOuhXzTmeiYP+RFnJgFxiWiXY/9b1V9QPyYp8NI0IoHLnQ
nH9m/n/BoiAciIBZ3zWTPMfvSQcGzll+ciyhht9Lw2o4XVSQr+AkpT3tvGqK2lz5
hZ70hckXDMAxU50ms8c1KRJZlpABg0vRmzCn/5wJCyzw2+VHDsOlVyy2DNsJ60Uh
uTGnP4IJyaSyXprVJvTPnGpGX2LvPuvxGO7prfLCXnUvNpeeEjVi0NLvatkDJH2r
/MXcY17aB2OGyje6dJ4VR/ZlmwQ3c5oUehv3eFUi9NIzvQ0PK+PY6dfWtYUswhBt
uJASBAOFTkD1qBEDAr8/G3hCdHDsuSF6m7JmYlwlZanPJwznripwF8bXLHZu8FOI
6+vS1eYYvHM09mk2YVIPZkIhlgotNAecfTeazJzFy5amGn9aVpj+V+bZDTzSK/I1
hN6zo8vp2vLhkO60AojmR474WLx8DlK5EbAba/bwMcVU4wX066s+zXPo/7ArUitw
/8Vx/sfBsqOEdsOUhiqnIJYqSJveo14P1zd5TuoaUzfv2UCsI6H4bCUsw8K9KvQ0
GVJY3iTfG+tF8NjgrCCA2ZZWdlDoSNv5FY2afXKtbjkNxCBdcWcyo52156Ry4MLJ
ZB6PlEvAWnTkxl84AszSx0YfRbH/Q4kET/zzHMAJ2tDVI15hKewD2LOi6Rwa7KzC
nf32b4+IhXS8IIYkR74NKE8hyDDj1dFBzqoIIaeDlyV7vyUVpYEPv085yW4Rgb2l
vfkjQ0skLXo6JFlPeq1m/BwWuRODWH6/7UTt+REBDNuzzDylenCgciygxZ1dNI+z
HMI6H4NFE2hmhVxgdQWzMzeHKGRJ1o9d96i+aAPAnl8BNc9+cUSieV1K7pIKsY7M
YJnljbDtP0RVyGs5RLOEqrT8gzKBGeSFmcSy/DjraM2Ww7oG8TK0tjvvpXlVfZS4
nVOsGOXvweyYVHNb574RLhsK4EVwvlT+Q0BCMp/31jrpn6e4CYhzAHCjtrRucC4y
k6YXFNVDNt2DxjUuAu/S9cbDqVNPMLKwiqWQNLiau5E55f1j87fZCyRftUmjaAP6
bRSheqDY6YO/D1B12RXz9U3LBz85LqfYrbLX23iSAzJxTFKbR3s/R8wlY6ZYiRaY
OJqDLhlkfgxU7jlWBDfc7Tkvgax3Xp7RmgMNczFrEvi4C+3gG8jHwnua+lQWqu5T
ouVJfFxlvk/Aabvs2r+A9sGaShERQIbX7Fq4C+3FJ2AUPbtseM8AmHhwrcsUWycu
d6qKNyR7LY3vdjnW49WEIfm3vFhfWSAhJY6b920wDZ2uzbsugTaLbaXEku2pK5Kl
P9oJlzhKfz2cYiXYTkAt3E6RhOXFH0E6Nk/hKwJg35fbt649GZd+hkoZ7uncdUM6
dG4IvG513pbE03UEZgs3PMi4RIRBGhM+hbOUF1MrsURX5QA8nrlyy1PGKCcBDqir
YGJmjkDWcM39ZjQzBGS0/9Gry+PPDD4wHuW+mJxmuNsnD8sn7FpRpLtgMnixHtDJ
JpZFvMuZ6sAhXwPRq4xEP9kYom3WEAO4Zy8AIp2jHD/aPQW0gfOLB6rihHCs/n1K
nouwHWKG6D9OPUtR21aMDv4fc2MJ7XHC7683Ct1fowcO4I4Mx0nw2vSYSN07IxkZ
P1gM6TSQmoUVAL31wMAd2V7UW40eKWs+E2xm8cFm2EyD+yuzNUpSQipYBKZKATD0
wNSK/o/9SYwSToGWIXgfgIoEsem+3mhVwt35OH9rUzMscTCdSvxSafzP5CB22nLw
lcc1ad2K1SdS94Mg4jubDRmqyLUObcB27+nyJFJtarIaezsdwrnBzue8VdNKGZMv
Py+9/uVJAYlyHxIejW3ZPk92O5GnVEAVipLRRVnKoFeRbplL7bFyQoXGfIAh8RHU
xoO6w+cw85WPB1oChiqslU0fozY1+GNHDC7Q7t1QGjBrIKY9asuiDZsde4Il9xNm
Efa4YJfj9mruoGvdk5iOWLEZFHp0YIshY7bboQLQ786ctJ3UbpdQp+rPNijdXTmB
u9p9Sva+05flrCxOcNegl7mh6NMnku5hPX3BNjZiJxM/J3Vi0mAykjq1/7LbCL1I
HI3hmID2QsJrzti6KCdPpS5d8Etyu1zFxIu/o95NOLU13U2b7AZhsKYzo3JiGqlC
oPR4lIaUEmZfZLCcEXgEedHyZc9d0XyZW9sMVj7Ztl1gPfEKMuj5CasptlmjAd+L
d4a6GdRnAAGx5LPyQjzcTinkLdb5ZGpXAebabDL1UoSVRbD//SNbundIt+pjTX3Y
t1Z/lqTNMzqMMSFBAlYCMrG9g+InqX/UCUVjbjhFZM0B+WLdmN8xbWG3SE5ZPsVl
FFc8gb7di+MbU5d+324MWYzKFeR+kOknGRxGmd1KOR77297fqH8Qo/G4g+jjb5Xd
x1thCUXyA6ju2++NnAHDTNJtWlVMsNh5rMYzXkNCBewh/yDTE6EkfBmTycs5Z1Qr
x3iG7/1+9weWpObUOXsNUk5f/DX+JiQwLYS3cZNW0IazoXI2YPKfUbaUc2OZocf9
LPUkzgX5PnLWIYSiVxpDgQV5fUSg6m1msxNO7UybeQIbylJX5vYhEUZ3kgBGslBT
tDAKBiKQD5ZdXFBx4c7VC2qunRfXU0oGJP2Nb8KHli+2AozKMEdHqMepeL9O0Zln
0GjfJB3m6t00VmV1hObhGqupZesbo7pjdV0C97s35Z3uCJUCDjlCf+8+lYbp6cIi
rSvTxGfR0ozQza4GaaHnQFdVcj8p0ccjUooEoCudjBLx2yPTmd64LJlmm1fhs2Eu
W9kJsuRwNU7cJh9H3DutwpMJBeuRjRinqRMixYxqabU+Q4efw0tELAWF/J+s6Jkq
QUbedYOmAFEPoGsfFB9sOpf8hUcIafMepeVFsLsJFkWXQdnSwLu8OZR6uLzPGwik
V8cbVLifWnobz6zacEciBTyqRwCYWcJJmc2mYbnyMzyDP/IRSmBGpe8JWwU1DbaE
cbmClJWjt3swdL/Qs0vn8glCLFm9o8eTVGVFBpKTKNCRZUWb9VaqRo//Qv+2Ecp/
NwrAq54QlTKwMyInA9bpc9N1O2I5g+/q54gwTOWWvCmGuhZTm+Gsl2K1fIj8L/qj
jBjs2L48WQK/gc8x9poS8NuhBGzDLhk3A6U7FyisNwSnm9bM/jfgCWsZSbbGWDu8
C88SN3SPGSfDq/GHWjaI0l3Lwu0n04LwC+pK5GuMqwX5URZx2WjmPvIkr3Ohu5fL
bEB6S3HZpHk+vq7WZSsT4z9I7xKLGbCrTgCtVjc0+xXbwKbdrKJucPM15c27Cia0
XxgMp2ok1cfMV6ZiegdrU1y0CqTVgdVo+66vkGXXawk+gAcDBPseRptPdnvKlXx0
iBJywlmOR08t8Yho3m2DwZOHghQxmyFN/RXXHlxgkVNWu5/q+AcqesSXgjEKF7x6
dY9C3/mp7UGf9UjIoH8d4jjh++H1as+lVU57o1thdyrg6tfn15XGtaOM+mwB2llj
yhMRm0lTr4begCV3lBkW2UpWawLQEpj6162XuYPUl1D0inwC+e0/BYW70Y6qdHlN
OGcifu0UZcFLDiWwQbNiEQTMx+auCZ+c5XLnXY72hW4LIVMADwc0+6FH+KeHnBXc
V1Kvz43gvC4P9BZnF87YlVCy9Gc/MWVChwL98d97jqUXl0nXddM//MB7LQg+G4zT
nepm2Tf/tXnktClgkY4hi9KgCZ9HjhBqkWyFESAEzjr41kEXb7NcEq9zHIwV4/nX
0vAYsWXhYfMbevsqAlE8MTd0njH0NzrPIMydX1XMfXi9VRYouda2VQfx85L71/JZ
AqAjHOT6YInUH4CCVRxOo53dVPHQiIBnm9y8NDEzfoYEzDjf4jZnO7cvUSHZUzLW
EgjxeLUQdVdqPZHwgOwIGs2zfLZJ9EpSVObC7O65q6Rgt/efjrNimMv3rSwJyThj
rAeUsHyeBWkT+XwUfuX0X39g2DXRkDRkX8oQp3SguOZNdKjW1TB7e2H++oxwgc/u
M74j6Sd/ych1JiFpbh/fvgv6xTpJV/vXLw3//AOaBztuMF+SHrdwY77DBUvbqOtN
rCb0V0JRtEYuE/h9m3WYQzkGPwWdcE6vN9hcvPNgyzNa7e8QAeY1hfOm7B2LTuOS
nYk/T+fjbB/nHlaj8ScymGgZcEGbrJq+x+4gpD70Jbr4jEM9iCNI+EoR7y79VJ5J
KgVhcjjQXHzn6m1LfF56peuXTHoXWd8XJR8SwODk/Evc+Z2o3haeDaJdq6gFpNfX
U3oe1itgXczTF6Lpa21WRlYdVSNW7tWai5Cw6qsrFTZVtss5c0kK2jpjIvJuUwIV
zdAeSrsW0ja7SItI2DPePkEgQuyfnIPVtUvqzXU66sjazoI18rKNcr+KjZWzXwxg
6dSvdRh38cxpJJ6EvNIU6OOG73yz9c8rK+w/NB0ukKWuKiwxFkdwkiXczNMp0Yu9
9x4Cog1rqzVCCq6GwqUWo3IDK+y7QBpzMtBNZlYYI3hRaYMXDRAIyjeuxgnMOqFz
a8nyKGm0iyyVTpVcpVRrFoeBhTOMnZ9GvgCD3Fd2l4bDt1y1Y+Zf7grUv6afK0xx
OONkTmlqHo1FarzRIjhYRH8QUEnZ6Z2vIVi2Z9HS3peA+kR2hi7yB1dLxsxWMPIw
FMWMd6uTeNaZsp6TkU6tTrDSNel/SZTzOFEEd5DB3lAS1fcFjKay2CL2SBGOKYRG
AEoVkHJ5ld2EtwMuVGzkSlfAoPw0VQHNmXzNMP3UtOa6a1XJnarfX68jGNbdOqod
fk6eUqO55QmPUbA+iPdFVeK4l5ZaCQCxILgHsDVw2sobvGAmRViW+eaXjHVHncfZ
8UgLiKzvFhgCY5f0rdRHMHCKRrD5r3W9QRcT30EOzRNdhSUWhN2V7OIgKJfE7PAv
5Go3tCXEzBjkj5g/Ofel3vs3RcyfCLgpR6Jsc71qf83Q9h0W/ffNAMFV/E2r5hel
/JJo48cwOg2qB4Xkegp3zamMkgZJZpj9wNeP5LfmWTabyaZkRFcuv0dBZeerMH+w
/tULH6RJwaJpqY5jbsiT+I3ogxwXiBv6DlNwCGMKFV2vNq0wrTIeKYMK6qd71n5q
RUJ3y6bry4vyJX94abk6IO2G0mmrk6O2vDpOWvutkJarGKly8IYXbO6SapcvX8cE
Mg9IB74EQbGzzZY8UN71gURZB5L3z0PUHhNCOpiCNOBYxKnj0r05nEnfl3fgv8QB
M5zA/pTLwsk0/9vK2AiKopEryGp+hHpmcRrhosT0nyUBNCh8eGcLqhQpurMG7JOZ
EeItBPYUUXvehK5t7G0cAF19itGTt0/ZMg9LPWr/E0vgXoFiYQggEv9IO1l7y0XT
gCzoRzz764JDbxBOKRNLu9Y+MGnJH9x1u2aT0PYyeomd7FGLR1D+idJvbbFHy9mx
BlUf98f++6WOi0a0SPq01cla8BsCOyFhbNJFlVIV10LXKygEwaQA90s4rQNo44p+
BNFXtzuLPfa6hI1ekSBc3HfmTSmvHn9KQYAfRuN9C8/mPlF+FnHZhK1+WGYzLEui
4SINKLANrf/kShmwBorsKM45EYmFDsDK8H9UWQMLUwKrT0qWHoF0H29u3gfVc7O/
LU/BgMFE95ZZYYCHBAB2qQletA9EN2sFILdE3XTpdnd40clxX1blG5Cfp+LTNAL9
huIq21iGL7Bwc45ZPVTcUFqyvaqqA8c1TNgEhFupSVVOPDgIkjM6hcx0Jf1pW3Dx
/kFdiKydN5cArlbIv6+jHQ/E7LSTWIfbF+HpwTIzzktoc9Oy7INCny6Zk63/MmNZ
N6keZPtviWe4jOKS0Xx2JKpZt+zETdbI+2mYrAYItNx/3Tg3otUrvW4EKLoztDeX
RSzA4iw/v3fp/0aiS5c0f7LGbx1+TkWmnoa4YnH+qpCoRBD7oa3GWjIc/xVcr3Lj
Up65FjUxKHFEWMkunyevJ6jTMFgT7IkVWSod5c3QaXOJLensHYofcEWcRe6i+bON
QXjSzDHB9pmvTZxjGY8IE7ugpkeNo6McYQc+VWSxyP3xwBcLZJKybTbim0Ye3iXk
8Qahxw2xE4SDMFe+j9Ltv+5tDdBOiCvyvlhhhAoEpoDfCyDbMwBdctgo8sBOXLVg
WpXRZqwOjwbCnv79euJTp0/nFAoM2oOfAxVVsTeE66HOLcBbiwh4GYauZJEaeryJ
HuweTXWuWitJaPf3q/Zrvwwp5WHY1gkMnvNif9k8hk/ty0UTVJ9VIB9BACCt+w4G
WBHZ5pOxC8Ffu6ej+9zl9ed6sW/BFXZ5iQZDVSQsRlrYAGEFnfpPp7szkFek4eLr
+aQptWZNu2hRSfvK3As2k/R338x3HNUegvNNT7d27kGOn5nCgGRqvqM7MiwxyXC4
yGysc3y92wYiylD3btaZU8aURmuj4uJQ0E0xHpLxrodzgSdbB8UelZV4ZHUP+S7Z
lg+GiXhwktdVxMYBjaixWnZOBDjbH6JEfqsJerq+AxGkvDRbLn/Gd1122k8WXBT2
04lXLin2qGtJMC/ByedE04TCIkUpJpNUNU0Wd23e4aKjZKrEkU9wcuEvCLxMDuc1
PFmP6tauXUSta3PN63QahivQDadU/qEb+k46vMUBd6RgwcBqvE9vbCeqAwusgBGh
fSYSRAVlsVBJW75nntsv91Ip0NVLT3W82wWE+BtsAQPP+APWwjLonn9CiFD37eJe
VumlOvLbhrFXHoQ6lywzHLX1bvKcOQ7iJZH4K5PS/tiHYOo9+IAl097WPps5457F
5/TBErDBMKVxJeFvYTDW/DIx19eYYFZET+oLp/nmriUQqfQWbPLtZSgXQS3Tof4v
QD3INIg6fj5aPXjb65AeqtV22r5XavFXBxpSho/GltcTvx6VKRcdSal9tMwDuArD
3XotiehmgWMgcsJXzbfAur2nh9EP9VGUt6ZtVH/T1OQPMcwENXrga2ycOcgflsvQ
TKsQ5qE2fDlApE7f2/XwxHpyIKNDvc4wrgc6HxlCZcQxTXaiNYwO3O5TGECr8Fk0
o+R+btKM28bSvVpVwKfO5PQi1WTl9JhZgJxkTwZcEcgwkzq5b/kuD+g/o/k7zpcW
I8/A8p1HFN5hfrrGUtO7w3Y0aMOMRQ2AAox7fIMkhl0pneqF9uV5qJhB8HOXhM36
2YTFD5ax/bxLbeTTVbzVdiajNS4sudGKnDV6K/6FPDpb5Hs7ck35Jq4+Nwk/IOde
yT5YXQcpa8icU1pLYIZ+gVsoG2JnWGiHJ8PoP+e8lmptWfBMDnolSGiDldBAxh6z
WHD+cKwMZc5nx7YfOAHQFqIBg4XZSIPqsZCOef2GjhnpdHKo80w6r76RLhOhWdeY
S7I4yJMyDoldPLWtR8pmUFB99NRkvcDP0827a8UtsE81e/A/BkwnAOsIzuh6sEjq
V2nliRbatn/55eoKN8rko8tBUv0uiI9RVSsXyf4AhXFinIvWDTfh2Z41i6uNjgnh
oafzbCY1tAboRGjF5LLLAAi5VEFsjmmoBFGHv9altScKYe2bVf+aSJhpIPvpJVnN
dGsIdMXQnYTR8usuSLzn89KCz8W5y1o8v9ACVvuov7QgiXHNJPrdZEyotY35D6xH
P0JGM9xpXcHa9j4Qb9fK6f3v6J45PSTUzeOuNj4R9HhP7igetOJQcHCEUF5PdRZA
gSz1GtGn3rRaraN95+ximHpZNRvcWLhQvAlUc/RT2tFu0V5JsgfUkeYLtCBCBvj/
FLEuFReakt7ywTP7kKeK7FE7WwB++x3fbu+QIgeEb9mzPDjc65BP9YWvOLf+hXYw
XoKeAyQ3fh1vcMnPaqMnSTrcrGSBiOVJ9vSecdCO9HlWhOVJzHV5t4iAGeAYYktY
IvuEjmINBrZ/NZb82kxMw2kUcke3azi98WBHXmFanslHJsMsqrT5FFttEKV4NLew
BnEuxaRMRNpN4XZVzatamiwxzzi/txPgOKQ+9QzdMcPeNZl/U0UMN+xxaKFhIOcf
qTG9iD/4YS4Be31iuApZkjrNzu5FMvUDPWH+PR7G3uqKl1kmGQFPsIDHt68YmX/V
YdZXAuX6Z9swMMvjnrgCtcRa7tzj+EM0LT14tXJmkPtFnx/QRV5girkJq2pf8lb6
gxL5D4uKzetmCzzE1ymrbnszm3Ac3HXHo+acyVZSmRhaf8jUQhn71sdHs0YsY7SP
ZxJxb/xEvS8DpTW4PyjEz1KSQJTs4UGKOQ77aXA5OSyjtSEcN23i75OHBTXux1+c
IdGFViHkq/DSlW+q/Odfpu6z9gF1EHMpuoClpAchO3R25CAWEqCU0Jw8GamSF5S/
1hPsWaKrskZQKKDy5+X0WJ4oGD33hAgu7vc0zjbO7Gel10/0Vpg+byssMs7nTARG
6Q03B1v66nRUFYZu5PgFibHFFBS5TdTzHyaXc0mecGCCNtnI/kMNutiNWP0+PNwm
BkNciVTyb7qEpi7EuKK+SaWvILD8mJLizAMgTZGor7V6npM8kZx8U45trSPZdq/s
c4TmuLxtKK0+K1BFP8yGqQENPScjMk8GLqsIzXEVhoaf6gZdRjycS+9D46Io+ISL
ti0dx60irctfpAsFXC/Wy+sfLrPIn8wvSsDJIPzVJQJM75kqgxzPrYIZz5cY08Jk
KzXC3YwppodVezVzETBQcitS+iYBploRRgOLWUD4GBOXdguBOkY08mkbyy8Oo9I/
n+ALAB5VYcKwnXzP6INvD0gEzqiYrfqsIC5/48SdGboifwpL7pnO3cGb9T9477+c
c709rExe7wVsmSxKpi3yvkSVb0rsUPxx746I/7q7qNFKo4LgHh6D5RrGYEolUmBq
DrMuFCIztXQmCVR7hA35jAZ2otNp6EwfvLvT38EsUoc7V93qvN5wxDF0VRUViqf+
dzctg4Vx5o/9XYTyJunXq0Bi+Ok5Bi5nON19vXAMNF/K+6Ij7LrHlCJhEPBA9RgL
ShJPvJeuk4oaOQvD5Arb64qktBe3Ct9t7In0s23a7loB12WjgLW6IblkEIBRQozd
xYS6+BtSAZsxNwKO9DTGSK2fHpOYsmlTrqII8XKsgaYZLL5F30CfnAF5xLJu58GA
MOku6TFMwB362p0O17FrQoc7oYadWlep5GgKXsY0ugVmfqlo0XrkZ65w5jmt3e+G
miZatpxmXMH3CyCU4J975/I2ZGBi9fBXKZjWya+0R0Zv+PucSWjRPvegWbN/FRjN
Cr4MrtCI/pWGIPwKWfPIXgj3bhPdT0CiCPLhSXSMfKUF2IpetVPZUUpljNNe5KsE
GaRUMS8KsTxMj2cfgSj6B1abNpXpf6TnjRN/muhAo7INs46DrXE+MRh2584LeM1M
os+WmbvnpQLL5MQBCWsDhQtnv0Eb8gf3XPU0qjsd/KXuuY2p3pRhvv1MAnoZBwpi
2lJXvgTzXMGdcYAdVjajx23FIpzLB5Xd8Z5tlZ/ZuroKhCxhI1uRAPzt7sRMHSla
mjKz/McWiVF+PVyMZ/l2RiJgn+tST+41DIaTAfQpT7hZ3e6gwXKsbe55usucDdLK
zHQ5imknothq0JGol3VMHC3VMITtornoZghk5wBAwPfs9Ub885j9zRnL09bkePxZ
uavf0QqzsW69JvDNShGyLKbB49eHbu2CaIMz+pddaMC0HPyMMXmJsEoipFkstwO6
HwYRkqkNrVm2pi/4oOIzzq6meSOYzoKVZS7SUszQDxXcRI4Hpypu/y2QTQRCeLMa
TZkH0U9uphPsagj9anefthmZy0gT+qP+AN6wr07jNuQA/GJd6w5MDCJJLOAF+UJI
LSoV/Hk23zwfKRkdDSBzUHdEEzYFE5rIkGYX2DCbcbc3OK9PHFImlPon19uysaXT
NUyEa3yA6V+W3I/1jjlL8gvVAyBWsWvPMvne4S2P68KBWSagtS4SpfVg5R7qbAoY
ELzV9VpekyFR1b6mbYgmMRd+/xicXj+SsXrmLBns4ysBQFtwXK8BYTGst4N9VTCD
FY0bG3pKgCUmMC5A5DZHE7PBB94vdDjPSJhj01VpX/GdRBY+9BI/BvGvaqzZwNpi
dJQ25szyBaqIO//7f1Wkz8yORruTMokqAqGn7CoAETn6azivMi/YNFoVRH5l2h77
i64bNXh2ufCpHKG7zXlE6+6Hhpbr7cFNSJ3nSU5yREqErq9e2GqxcSS7HZx5FFk/
EiSBLFeLN6syqa/MpCyiJdC+nMnQs8G07DTY/Mt5ousd2BuYgBb9p7oMXqrvDLPC
1Yd3tUYy+Yd1458JQD4sI/ewAFIPW+Bs61AIsetv2a09Dpjvi5d4uQ9z/SeSHDEA
h3hUPI3PGSBSJVjUXNIpkl0i7OLqqbO1j5ZImGKRsT/lGpLloa4HrqcoY1b08t2e
PpoLw+bz/wYxlmHwVKCcNUNU03cn+/0j5KHdD6CvFco1cBZBcRB9iq6b8uTsbgOs
ljnNcXTxHcl49hlxOEBX0WVjvbCloGLzRHY5tflgz3X8HWgK4rG1Ju3wX/NXwlaP
Vgw84v1VqHoNHJDnIDDeJxAwqjQmMT7s13XKqv3406FhZ9V/utrjZy55nrC9+YYJ
wNKzr674lDonT9CIbFvbTT4LEjUvPEFjIrgPwRqSOS3I/EMdUM9PzYm4VfXt3wgi
Vv6ru3MB8iMXnQSYoTdi676GSDR77canhRk4LZ9nVoNBjHNcmubL1QkysO0ZdKKg
lgO65/o1AV1R1Wx5yzVqZhxvwSvxxaap/2eQ+iLEEJXXTYfli6Mk0SbmZSlPymDH
/x9eP9JUDALx8KOe7prymwmhPcHbM9FWG8u5Lv/ZGHdMvTDQjzI4H0lEjbp8l4rD
9J3FaYMENo3WhHW0gEH2TjD3rpiOOJvth/cz5PzXP02VoR3M68+ctM/3phCiNjMQ
JHUVhhv0dVXGOdHqr8q4XbZ70JWqkqVOB5lutlJdLke045e2IBaEXUiGOsG5UdaZ
XDsqGI4tayme2cQyh0ZN0zPYqvrkK5DYdZJc6/ryZFY1qI4Llpt+e+oaL6QxO3CT
Rr5N/W5pGkkyB0FnwaJiVTDe3cGO5JzDDY1FwVgtid+tkpL7xi22k2zG+zDw12i7
eypgRQJfqKbWZQRJCDiBfhGP2nBn8M1/57N9UWiACXi42avTiJ3K62qorOssmPvQ
dXz9LUhMl4yhLiiJMymB4IzoJcA6+FiZj6VKD29AB8rOjYJj5VPeaHPb32UuXZsv
+tE0UUuUkQihIyaJiC6uXr+dueP36At+T7Gsoc3LgnpvQd4+NTHlUBEhRGdbEAPO
MfvTOXIBSdJCVVIdqZ6CcrcVA2pbWVrSvzoXgW3krAVlzoeFYZoiRFJG0Rj1QhUO
zLWIId4s9EIa5LU+8jZdbJ058AQaRFpq0BV02gjwovWPWGdZPu/21MkSX/Q542rI
PWXLEKcW8Kd2pkGZPNIbZmVRC5zBVYnf5HPRI1m0DrOsK1YDZlu3jW48ToXSqDe+
VE68KlIYLpc+oWMjYgFYOYGfXK186+jj+URPdRZTD616gqbI/woV4Z9LmeGcfllP
7Fhwzu55Bb3uHaFR9KmXR16wVN/fuh31TkMe0Q+YTsp/bn7XRHEXgWAd1YYRhRxg
6rsM/mVMQtx+RaGPW6CZtkmio/x22rBnJDE5klRuveDcDD3SU1L6mt+Tm3wwL1Ca
RLeVHs1AnMtzwwjPl7qf0Oo57axEuqZDDBVRMC4Pnb7ZtcIo/t+DTsDJKMbSBrdd
4knMVPE0eKh52NM053MmWfOGZOJO0OX7t5WUeLm0H1b8+KsLt269XxdC7da67pQI
E0xBJYAnZwHLqjKHQGeFraUZSLhge1copY5n/KOilfs4GRm+dm7ozABFfTCnhq3l
T2u6vlcBmYCL4COQq+oosb+jaogj21vFNqhb4A5AiYgcEtMu4RRc8b8Jnj81MZTK
rq+ZbP5hOoeeCKhc95HL0yMZQHHB+z91dNHIxIN8damFjGybWU37znWmKtUZIHl8
i81Ph8+c5DLfMKTWMbkxHnj+Zij5vBvXmuYYCxCW7fOY0c4CBfb3gHzHs8svM9Rt
1uceGbCmel178j/5gFfnh4CnnyetDzlb8z/wiMLmtH2mDeXTE2FrJIe8hQJGM95B
B+/aTFN/1B0TiCn/rpqOPdJwDKQtJ43YZF2w2jzUspE1tXgOce0oBsSPW/Mo2W4/
9lHEwpiiFa/kA3Jf3orDbV+cg7qdS7yje59Zt6vXR3DsBqp1izxy+QCg0X6EQxYs
Xituh2J3AaYHZIAHRaE69HwBVRDTLGpZEPS4EgA2FIw5Zu99zLACkFwDJoWRgZsw
XRluAV3MLoxkWIJ9hJjdbA9p1efqjLDnFUc2M2s+tQH+bXnd+1dzjpmpCi8K0fEw
nAF7sqytGFuz3DaISc/wJod9k8ZLB91f1vXVkmbWAoMNwBnz5BkKR3RZZI6HWmbY
tW1xuGgGnk2gxhucVeWuKFkQWpwNGbEcNSukIqPa51JmyJhLdwsq6sTyz+v4Y6f0
lSfix3w6ZmXVG7StT+J3BjXVzwPDUxZ9+gP8inV/kU4v79RPpAs33eIWHo6twi8f
rkxjatKrR9vTAJ1k8uVoh7XBBmYZC/0qBiGlaib095nG5U67t6INTqpDI0mx3aAC
9XBD0PWeHnbt/HcmrVdQpXEZUDosJ7i3yxJHRns39SoLWCX2xsa0UGc+1xfSY0C1
CIDdhIqxhx01i7lPp1xzbITNCPBZcAlQ/8TsNgppRAI68sFnEot3Jug/ADj2cU3p
5E8Bw9bL5opVzViUY4F5jsk2t/oEjqiwMZdXPcR7QbtXUYCKdzBbNCGwKsxm0YVF
LYi2aJHGt7TntZEZgd5vk8KQhAKscT+tg+KIGa4a/BrKiPlTHUrJBJh5bLrOS7NV
Ta5IkqPmmf/rXerHVbF3ytbEpTp6SsjSwhIfjTS++a9HJRcJb8W7X8DRxl9RAROI
oyjGxLBr0EiwBW2Ji3u4cpE5nTkIVat6HMmmKcbON7DT6BcQdV07T9Mnnr7An/s3
lF7T1byasRz21ulr09VrNqpqift3s16DhRpZMo21ORHv/j/Oi+4rYYB/iI27oSx+
iZ8u5BrviO7+fHDPQ5Vp2RKCbxjf4t7KPkXS4pl6Hu4d+cDAOILQMz4ZahBvxHbx
5r1+Hlq+/X4v3sXV/GICrN+2HlFAjbUZsFJCOYl9lbvsYpg5yCmcNaNqG6U9aR1Q
oirjvJneQTTkKiKzxFYW9NWCO0c8qxmTITuB4xSNvvNAMRxE5Xdipcw7faE0Li6k
pxdfwXt1LAhdk2HGfFFyD1WIYdo86hsUxFC33xsBcQT84Brlmsl4r+rojf46mwTi
y/6f+KxhFeEKTM66sXemkj4RyJxBAbQXfkkw/rDgcjhwt5bx8eAkxo8hdfl7/OzO
5GAPbbqEBBfVtwR4Y+QtYEjxbkzJsunsxE+NWCNoFwPkU0EKhdwNkAeEgpoMoJAX
vcY3wIvCAkjDbWs33xIsCYy8GvDiJbLbqzEI5yvj2PbsqJ3rf+qI4PDhTje9iaHu
ioQaNeAyEqPNxlWgwNGiiYFvAu3ZhFEXWb6UbD3xUnC88zwZtoyYV09o3Om5PeRg
3RiNnbZbnyuvMytqz+mHZfIZi07mtw8Yxj0LOikZ5aFY+X7oaUNHZK8CtXLMUGwa
Yr7F0Xod5FQPo4pxDnQG70sJTw5XDyYLtKanjuYwNo+FErQ+CSTRE+uGOrSS9+ry
JIWN4Fd6jbTyC/6pQ9s0pnIA5rtS9Sj1RPN+WJmJQXMIrzI+wWiyxfE4oJWYvs2Q
jrv4M2eWLkWTKG2ODlvI6z48KQM6m5E9/6m4YdKxxcwfu0boGf4pIPLWvFFF63lb
biHUNSUfQXaifbOkkxACUnPZ4Bei+aIk9irJovBG+hnrs4crUyrv7tn2/cOCihZP
hoAmjPyDX5cWDVKZmxhL2TftXRKG/FqJR6A4mubR+N9isAa3To7RWdHNM9bIuhQx
GklPYMTGcqfVGv/OYDh2HWDiulpFvJpmtHVfkKNAnskUHjXv6SuDqYDyU5+NAP+X
fX3/Jp14gMwP3tUbu5l7NmBgVgrwCfJqlcy3B17wFjj2Ffy5ndMh44bFLKRbSzHx
VtwA5dFMP7fNLiEDT/jKvFkBA35OeWL1bsLkHzi++N1+LvnPxSL3G6kKkr5Ds2xn
V0BaRmMVYLcdJ7R2MMKnCznOXr0tTiBOoSUrfUwLFyWYZBbP/SHIovuL5JlIxAP1
14YQfNfDyT3Kg+Lk3ia1E9Ixgx90mYPthjPbPvbE6QM17KCDf4+fAI/xBiuj3wRm
BzmN9KkEyFGIiJ+N7iQyQIyhjY7H/87+iwIspLSLmtuI9YJf2q2wtGldfXN46/9V
WMCsyR1JPtZZbF47o4wfBV9rjSsJLK13yP9GlJSJ9Ndq5HufHYcQ04hHs4RpgspU
EE99E+VR8yoTYsYMZ+tN7KlB4LOPUei0/P6ysRnstNA0f3djn0sehYCW3ObrPpwX
83IRvqNNz0lfsPulEbRIPz6jW4cFccgglJQ/eWix/KlTMT/x+/GTWisXra+DrNO4
p7Srgkvgbf1NupcBiBNoI8yrByZdA5XXacCDUCIWnzdtc0ep1+bR2DwkjjFStQeP
vdFh7stcL92/EzVJ6vfRhahYopl0FZSXBvb4RE/objwd6G95iyhmDS0lQiKeLH6H
fgtSrZpzfD2U+uVsptxegioC9ZdhBn4rBL4my9t3YKPEAJrAZ5XTpV69er3EzXvH
UV9YNBeg4fF0CHUv069BS7Sr5NsK1wKdDzH61/xF8ffxd6FKSfjdRqLSOjFDh7/K
3CnhqVo1fLdXhuJh08RMcfNaMTqL5FmdJ9t4reGjnBlmnawkCf/cUblZzcGmCJ9L
ROkoNfzP57fcsX55sngiVyh3ycMZUD04zHBHb0kMiYmLxL1HG03heyLcjMMhj4En
livtHtBR2cUH/42ygqfPAD3AZ9wz2QiHJaGyh3nyz0MAotamVQ89ZJyceAqTM+KO
HXsfTtvHx05+feVv7BuOSx7t0qgpU9TSb2D1GKvtbgk/QvHqY2ASlrnolCnEwPuS
ulUUylXLgVsnoUT2B4FZbRU42jTtpPzDTq2vt45HylAKRmocXl6WcTLPGgABL3TF
m0q9jg1pfkl5O+DMu8Jg8AGdvmF/isyegWvFyEZgTEOyZ0dp9AyYkizzsVNVdNOO
siZiYaTn6HL01kLF52Msco2KR9aHVB1dab2R+aPTo6LEl5rwykYoB+1J7i5B8nUp
qajgW0Yf1SMbKxecDwIbWjRD48ezkK7DHYD4zdgDNdylHKt9VO/qTHSDIVCgm0Pz
I1QHYol8fDcgDfdGVIseg7mEnw1gXg/VmrDd8c9TG7qtB0XuYg9CBDsAWr53qlPw
twSkAGD1PPGenlRPNXQUGlEQbkHxhOhvtQ1+xrIkuLxmbUIXB0cJsuJlIxV2/Egv
Kmd+vO4PeGzM5qwgd/la4k6vBNpaSz8KYwklBfZtF+cxWYi103V4mc+DsxMj4k8r
vTCe91ikVurI1bRya6C+7MC2ZlapjNc2vcBVu5FHDhmRJXbhUbiGqLzkg6mq7cj5
8Q4OZkFglB3krqNf8xBz8HbKMCxXbeZNUkPWQjNCzXJjkP7NiylFBipWlnbNJRNw
p4FhYLNScduWVpfOYJGx8FnuOoP10xP2r4jJF/6wxbIZ7Bl2/zWCprGczh8Ln3Vc
hTZJLmHWWN29TKbd5tvqTWnpR7B971dwCfzy3Jak8JelKDHHEFDcvWhgR++mHwTL
ZTVz4aShP73FDpUtwbQrts8I+lYIl8ZI/jpkGYOlBimGtQFteDn/tYy3HB3qEcQC
F3JdvAzek1Iy3O26DfQX+6VldRVj+U+X5HNAfW/Y4RMeBf9B6wX6G1jgXRXC1PdZ
zG3yNCrbnvTtw2baK59uu7iFIR5fU3gMotNTzOx1YE/e9xRfETPQaScrB95/AuHU
6OzyivTVnLf372Fx3KQ1+OTVtYTFwAAU9S2lnvEEpPSA9OR/EAgSo7TPrzu9OyjO
Z62K3K5jFqguw6MtpIBqFhrwtkpotGpfnxr3e1NSXbfhVdiyVXJTO0RuewJJ1yUM
hf0fBx9xinNobhJwibK0nhEy1joa7FUp7JkOkwNeUFt958nnFgZWQ4rtoEjh5avo
7zra1XVVuVjX3DUwXzZoxTHt5P/Rd1co4w9R5npGc5uOF5bC5dVHRY9Txrkybioo
8061qg+APaCvQowM3A/ul7d6yTorEHNj0XAX2HQXGbEwdZqH50M1R0KkVUGPQdrG
sok36WGs7J7PLiqzjZ9wlnfowqa4ob0Ljqm41LQfta1nP6AqxtWQ7V1abMKD30nX
shKRLqAZ2DLMs5kWVvlZz4l3adHTxdjIKNz5Kcv1zRUiVHQyesIf4dY+fQ/vmIK2
aHdQ1CU7Y+g/JvK8lbiScMFnQ4w1frVCv0UNs5IZoaviTQlS+aZazdpqXoys6taC
scsNjBP4UWreOSa1wP/pd6SKGv+Cef9kQPdQ0Z4hlztjDWpiGoSzRcUanGd5q5My
NtD46VWv5qNefNWFwkhSjbEIZhBzjTdywkwkpkwdLboW5Lhh3u6U/P7l2xyL3C4s
F8sl6ojF6FFLRheEPuVKOOc0lHmeeFPIC65mo89fxgETFTNsR5V9voqfqkfF1u0x
5+JaKfnC8LUAvdGaJiY3AuQrJvjv6X3KGNeGTuDavm6GvBJrOMouyffdpanZd19K
kWJ0yDK/VwFcXsgxYJfo3kbqKHAzlqMNC3xXtXnje2q4P8ETsJfnOJu4Bjt3n2hw
G4V9kqNwvhFF2ED4+u7kGlTfBDUBTG0ZQD5CoVrPtr21/OWmlcJOzyY0XE/lvmVu
nsfowlg9QgfISnCtwTpTH4EoHCIitLQU9nvQJR9WeN+wQUrqWbZvUZIorVcVCD5K
1QnY9L5iUYyOmvcM0iqGjbpibiPwQXkFqB1sFDBmEjCzXfO37TCVuB7WFSGPkU7z
IM12pF3adjTuKFQVUsPU+wnTYFDo5FbZKZ2fp2B7pOGYZkqY1DtDhBI7TIXheLH5
vGfdxfHO08ErS3AthxnqgUuHJs/ocRKqdLiiBrsugQYlD4ngo2JB7DZLL+AXKKAE
dTJL89eQAJRaFISqXpGiF3kH6nw4a+kV2heiHXG81OuDbRFflKS7NSG/szfNSwXP
W8Y3uapWGaT3ipJUE142O7Tz8kqXTyZIkhK5eyjoSlk/6JB7+BWX6ZmoDWFWR7ou
o7YbRvlVaM7y8q0qpXBpXGCHapJmYArpUU8ZgeC+bvOLU9wurGk7isCwkTvKWGxO
nN6FQP7AEgKfWDaiU9gWZA/MumBvwMos2LoNJgOII//x0YIsyiglstb6L/VlZSaF
JYLz8Dh+RkD8qX5hdxgS/5+9CBKvTamUuaMsYq99IU3vY5oCNrPg952TGgPK93ia
ebuFeN57LOZ9wTjjAfhNubjYZa+bTwvWx9U0SohEBsHf7s5n5z3omuz59NPOurCr
TdurhHxRhWZ/aMXgk1r95Xekc/NRkVHfm7EEvDRYC9CBOG+Qvaj208m+GQuKdjkd
n6CZcenchRFeDrfiEVLBDNsPwBaBcSjdf2/ShewoYvOsq0gVs4fijR5emUMwZSGf
rqETlANEZiro283RFVoUB96JnWQ/oxa7P4EtTUx90t91umXmsHjjQVRU5szRBwfn
SRRP5jopST/1hKCU85POIIq/gQ15fSYc4DP0rs7seXi7nbWpe7w7ZdUDNNo6d8wR
+XurSDz2BXeC+qNRHjQLUKh3+oIgso2bgd6xIQOETJ2fWAa6jOtUt9mQmf1qvAXD
L7zcqC7aDw+w67QFmq50DY/zWhgo6I717r94CglQaETdCScLVMsQQYFqwG3HepbW
3vItjNZdpgBHTHKX+a4zevUhJO1WVPgMSqn7/qaFarAsVt3RHcK4LemN6iqZCXOA
f19Rl0Xd4pQE8wvB1Um6ts0LZYSN/qvpmHgR0pA2d8McCJmdPnaV5Mr47pkgLTjM
KTSNBnHJGOEPUl8jdSZDgKusX47oIjLskFbB/R8KplqoIo+EpG/zTBceoqR6GfrX
RvXaslZL71E0X4DJ7eTPgR36rkNkOfO9C4AxIKca+O/b0R5oztdCINICzyXLNJII
xD+vMwvBrnGIKlqIF5sW8tnGl7bVF3pW3Mw1Un23ysNdCIIHSd1CVFN5z6VeDfaD
KIbJd4yBYkEPw0KnJEpMuFL6zNXpuNlH2bHJ2tM0YwkQH2PnYnYKw/CvzE+G8MgF
Uui8fLXbT8Z4P0Nm0nTPEvIDuVfTHgkebjLTZ2Eg9EgGprmwTKEyCvjNLy899Inz
WLLV338/hcGJXD76zGpWWAUi5yi4lvCTxpQkolnzujT4z/elMTKRDtoLyCfqWfBZ
JsDSnZ9xP3Tlnbw9shgm6nx8QhA0+YZxeDCB2/mymVIlJwkVBkZy5jpPNvejD0lZ
yHKhDndr3RvNm1sKt55vFdSD1uvHpLDG5ufNoLZr6z9wUOFgnn7p1RLPDqHSptCk
4/H6vBkAJkLQ6dsI3MLBJToToL/L53ETHxkV+qQRMqcqwJ64jLrwgsC3gnMGVIwZ
wXYPJKmzuux31BXAZU/j9PeDYTCTiBqZ9p87IG1JPdwHVOlj67foSAsoCLceZ2Rf
NCGVM5x1m9Jz2nePN8/snmkuzo4Gx7GaN0ls/AHnBPTR7tmP/Oet2FNXrNZ/iaQS
WRaMNuDsmACCglkKorUrcqBRzzxri7eIxxc5btOUAnx915PDlXnoofoWC37hYSgS
YUybdzheq0dI59bw40NrzY75NLnSDx/g89QEnELCSloZte0mLetI1xTwG+qvZ+iG
VpkqxltTE4Aca5AHO4SX7FTKDnit9AYJTs38RkxOSLwY1ggZMjHTVGuTtPJYT25p
CfzEDtDDjsWKSmn3ru7iBhjZ28wjji63ivGk96o1yjc8H1C2KVp1Fo9v8yXgLvVJ
L/XGgKwncPXNxArrXMJxdfSzUpBNLAVxNvubZPGpwDANG/xJRIKP1403yuJy4hFV
0il3RHJ3Bs1tsdQBZUg3dUO7K2SbNUtTX/iqRqVkLSxFpWYFFt0DW+YnQcdKGwjz
833zVz1ijCBxTEAtn3NJXQai4KEgHxjviw+x2s6YCLV8m/zT9PgI+QlO6tHMLLGt
R8c8qCPqONHjmGx5tKHeSHO9vleZwQLSeiIq1fIqI9XT4VoOCwl6ZFEFJLCe9Uaw
ctkBr+Mpwrf5FwicbRpRcV56rneef9VsSa3WcF6fK+LqocwTKQie3vlBJhOH3Gun
LClcz/Rimd86Lz4EcR6mG+wxrIx6m6TB3kFYypmqi9mO+xbQFmj+1YbEQ0GCid46
bDG3VxANECtTOxFpCUcg7Opk5FKn4j3g12QAXFtgMCyoFfMuUi5p49hh5O0RU1Vx
dyc1YMzpZB553s5KLmQjJ9wUWacSfgTfubJURuOjwlbzMFAuhUHnFQZ4xAh1fAhT
Eo0xnaxaA2U9TODhxgD9eRSDhy4vTGKZHfpbgtp+8+XXIfpbomwvGiHde+eSBzRE
bohIGtBZ264v1yb6dPHQybgcWbf2wXtPCz/vvNQaiDaYeLTwDyU5aJWfWBVAlSs9
CtikYzefBed//+PoNR/VmNESGcBzVqLWw7GwaRbvxCMmlwV8rkBioevWQaF5MmZ/
rPLdoXsbuYgriJ5N3Q3VJUPf50UZksmRpNt0ScJ3qG/5+Bxj0Tlg68C5WYQyrxZ4
V9w5m34h19ePeU5IhVjrvVg+BZfX5XmQQ5AvcXtN0SHMHItpbMdvhzpJmnJI0hy/
BCc8KNvtLOWfrDmmhYuMqddT68ze6/i4xqCT9FI5PzKB+kAITQHujrDQPNW/wuKF
qAM3BMOL5jaV8yCO/1vGVdpB4SqDp3+yXzVV7Wl0zbkb01yfTanyALZavW+dTbLq
ejIHwC2WQj8omBX52n0s0v1SNMtDryTQ3Y3erKRPftpisHnmGMB8fDs0UuRlJUom
7Ag5lfataUmgx5kkwmQ0rW2t7IKX8sKf2ShUAyb4j1VXhk9gXIry0BiATimvMyDC
ss5cnGuK/ZuZUg/kw7oTMKrwcFF/VTaqjhyR9KHTtHsberxF0PgeoQ9ThA5cmhU4
gMn2dlclXLfnkcAjoT3CG27/cPz6MAh7xHeLdAO04skOPo/BhJT5zxjzJEu7wx20
fRxAcP1km3kwGkffZ94149v5tvJbHxp5sUvxzRQoK6uVoqkvVJo9GflHzhTZA/34
t3pp/NP0LJ6DAymYuXiMav1mzjW0r00cd3aH83W2NajtZfX799PBOQesXhBteXzY
VZ8ecO3fYvkbTYvNlpIsbW+w4pl2YbFjRSpeqKut4ZwDyhOPckBZLkM+a71iEjw5
rmlYIfizPl8jCjQYVqr/eFU+KXJ1+9BSyct0079LJMEiqS7+jjKwKSvqTwzSD1gt
zbXjClZ5cej6tlWM9Mv3BZSSuBVWNFDr2lSPcn1BRmAU8IR26paevRNnfMeug/HO
hQ+5ASIP3EVcj/D+lrWwCBlu62b5L1OnmCm/PV5I/YJc3Om9KN7LxiNpqcjQYX6O
npSuA7JHS1Xmosn+tUDq+NdXUGDinp5OIhJrhyOXYhzLdGLAKAgG25tUNPPdxuQn
ddbzZvmhuSPgZ1HTdKWoIElAmEkPm34WfhJXZHHyQZyxtQLGNDMIxzIqfAtkrGtu
FPv4mz3ZodbKGGwc8qeRXpgI7bZaTUm4fnEiCAmIj7b/quixVEBfuOdi4nzpdRea
wPzFtyG0AIXZ38yVUOzMU7Gw5vy/o3fCWfmEbWKHuGLJChNOh72T1JYMp4llmU5G
qGhtJRa2Ygup2j3x1UL07j7mbljk6H/m/Azf1vvP7AX0wqSsC4jY9Sfeec8tNxm7
Zb1h527UVT8usk86as06LHkKH+cWNdOQQQ75rSnCGOikmPX+TWNGh0lJaxNUd0lM
6oP0VipKXyOghBzjdoWNQF9o/7uISvfuB4kZaSfeYpbb511PTds1j5CPjXOw7cLm
qrg0Rr77m2BfNQnJcbB2GR63qBURQ7iqz0OoNu2ydloFgBLkc7lyWBdWAzm5WUP/
bi4RedNH0B3m22hmi1HLWQll1hUFLX2AW0g7ut3iXBkRD2NLlWo/1Fn8IJQSz/Bj
VV/cb+AliyzIkoqzIWJQ8AXWVF3b4C/SaEIoPXe2B8p52lG37TNRv0R19PdjBhi3
At3g3+Pw473oKJftLbzt3CG70Vl7DWPHd46I9TfkfZHto2jSO82olcsqWAyCWtel
crdrKzMT/N5lOfQLspy1gdk1dBSM4UXdv3mwfTBjVxFl0moIcuWrLVgJGRIllL7H
ZEKCaNsLdt7sT+1rSL/OwUsPqe7nr6TfhWCo3TdUfFjtLRrDNBQTjx5QBPGDIxsb
xkiNO7KUEp31jHQ/GQU8+dpZCr8DtSiUnab+jgMM52JygrNW6K39LQ0ORycObsEl
C5FL8+jWzCemnllHMKig2QKkpfY4S2Ss0H0vyf8Ync56Y1dm6AkV9k73MQ5ARWuf
owa4UNBdBo6IzFpaU1rsU4G4PftkcJ6V5HtjV9c0xca/rXgaQzYYFWwOVQdP3CZ4
gKBwQOkmaVocYGzrkASbvQ+kb8ZSMSQQgBlypChty21ytvcFOPfaHnq33jS/a6QU
nqz4fYW3BTR/6s1Hiw1+CGkW7OCRWZiiq5uTfslQSOK9LNJ0AykIgp56MS8I8sVa
XtrrFgkzOWNJtuZAMN7MDzgjc99bXXM2opyoFw968adj5maGDsjMVA4Ae099Wk4b
keGiqOoCTTEFkrbYrNqr1KpFmuf0CL94wgMM2+lZ3OIGFzU4Lce1biCX17IsUmSF
oXBM3y3x/s9TmgzMo2D3F34oSw3x8yu/6PYB0HPwDnxfTAu4p6tfvhh3U9Ok4V+k
lt6gpz3hAcuQ4VFF5538wqE5ilQPngdZhfvYTWeRBQPeygSwpcD6DejErrQFsYaq
SX8GbNoWdE6FkbHGB91Jt8DN1esbj3sC4RMm1Q/fKGuVEHo1WeIcA9C92COYo9um
EHsEyRC2ToJ7DPtVquQgW2DDTeAGBN5hQmIyak6uGSVnQNLqzXC+nAtIW47R1+BR
QLypJH/81WDr23M0KN+6dP7qo5IPCHzweURtzAP0YaLAptJeWAjeJkmwTXfz376I
1MHMmhvehgTWSVQKG1SZFzgXaB+scbgls0zhQSxd9T3lSEDzQRmaFJiPsld6A1Iy
DhtysaFfaCxYxYRYfHLS8KgAsnSoG1Rl8dOclmgPlBEAC91J67cPqoMHdrFx7b9y
k1GB2g54VGmJO7JWWJH2zKVliKL84IqQ2sQXBT1l7Ph8QNL6bh4i4VfwFpkVypdY
6HsX/5NCp0zWcyV6k6R8PL0ldtz/lx8+gE0oTAz3HPiqCUgucX3R0j21BIdzKBpU
uNR1QHrzLyzgsOjrY0YBiyMCmY0bLEKBb7ahxAl/9/phJXiWaC98Hju6TyOQVv1i
ok87JtH0sW6mLsEU/Z2X6Uz+0xicQk2nVlY8+gp7A7d57p5BWI6j82seYYiuF89R
k2y8yciaKnvMQgS2wr/XNcJFmfDxw2jwSqsU4N2871mXJPc4u31yWccfCcXDMKCf
PcvqUk1Aaa51tRBizjemTzS1BNBDyMrgxgYCJYvKv3CMAMoh/8UJ1lLGZNphv+a5
QN7f5dRr6pLMcgx/2ZE6R5b34495HaNy1Jlx1X38ow1RWJNuwYrIRSLbd/0QAQNe
jW5+K9/N+VMo14kys0IxLt00S14qtgeyUedISCo1VJrXGw+60gNCwOAZsD/fUyXp
i0iDnGGkMTZ/VSnq0GVgKqG2G+m2KviUXYAwkYgpOrXG4QoEJ6GBx+FDJaY++GT9
mODFVkmWUe0F/wZmiJQJcpTLXi7UScU7pXOgBaRsVlJodxl92JerTWdVXdldKzMd
DMAgXUOxUR8JCl6czMnJtZVfmiKUZvEFDApS8+XyjYd7dai1Ci6mWoGT4z68FMx5
XYTHi464zoCUBp7dg8lIZc3EkQN97ErzZVb4+I3uoKaKcQTcDmlBciYKUZE6B9r+
qMiLnJjKRmurtSprmzlufXt0f+xXTTWB09NAl4Jl17/q8Fd7mz/tTqyE0F/gwF9k
feYXhj+Vqh9DViv/oIv7vJDeJpBCpcNKiRQ3/TMTmj7iXk3bJ4c5M+dwqZvSI4Ww
M/JW5cA5l+5/XQfgEl3x+vg2b+TSjealqtJx7cxBT1ovGaSsUPIYg+C/83uClZhO
gOgNWjF+JhuQWTmNjSaypfstH/OlypnTXm02Tc2HeRDSn96/BCVlaGINcAjJ16Tx
8c2GmahHwbazroS23QzqmXS59HvJrqu3aIK9QHIu4WOpZ27zjQe9cQLv16t2uzUj
D+hw4ZgCb3/tKaOK+qY1tEzZtllH7K2fnQcG1KvY0E5KlOn710zwSMjdG2komLDl
jvQJRAP8bbZmSWFqevgYDizCRdPGoPu+X7yztxLYRu64D9W/9tEO5oqAeozRBQWl
gU1u4ZjeYeMXobT8Q+XZYR33ZoQ+f3VohT8jRI5PMtBxa/+fxNinvk3PAQzT7zsT
mFJKTYvQgwZ9T3G4OdU4P6wC7eyji1/PCD/SRups0OAs8rLuYQS1lIo4Dl3TH5xf
YnRI4RH9xsIQcKg0m/EcIDz7V8kHFSjionJxARrqjvhR3lmW7W3wcx2/qYy6hMsp
XcQawuL+/RntAV0MnnOfaHGsZ+47Me0/AeF433h/keeHvGg6ADW3CmdFhMb8ufXn
`protect END_PROTECTED