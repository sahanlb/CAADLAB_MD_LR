-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hDeoatANJcswzLNAkQuNURCfnmbf1KBAp/jAkRfmaDC8b/9sUm10Oun8I2599Ml4sdI0WiurD0q1
J4lsZGsRw2Xgf6vJlMQ204NjxiSOPk+feJKvAY7PVP2vMWvidn9VBeLh7+424k/UZ7HSSMQvbKNr
GMGEbHJ8lpdNEa4DyZ42ofJk2DIr7cCXTNCilULA1XpEmovGkbFk5feHzIk6ikW2AjU7IAgwO60o
PMdzm+8xAAfWA0mL8PwDe1zrFHpPeBY/HD3OFhk1KebBrOwM31xtd9txatHCF72MYQDyP3Q4j4vZ
Kf4dIcbNFHFY3xbTVVgTZh3lqLHa5EaQRoJFIQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
HZuPPLlzu2WY2AbUvB1ET+BvJm6lje2x4EkWlip/FoWJsh79XvyIRTSIULqa9bmuApQm7xaBDnWa
v4yGv7qGgAk7Zwd31gVAudGVKVVrW/R9lq+K+v6la+tcqfpBTmT9SRY8eSUtskcbG4H9DkclU8mF
GO4suKBa0nnwDWwpAxI9zJAcRuPA3xvDoapKamW6k5b74FSdoXKoutqlxoa1173vFMKk/kxethCZ
EBFZsXHorfWUwxCCZhE2sKwm58H6DhCkRqJL6plAOQBnRydSAODUqBrIHKLaGuQYApbqfFEivbfB
+fqEKX6A8B37j/Mao3ELNkpnuYqdoT2xRtbyFWael4cUIiWqaGcPwQwSjDoYy4SRG1RhFMFOiKB7
ltCdCucPsryY/RqZjYpendbyfFfRNZPYZtBtjJLBLHPuDhBAR4uVvDNg+z4AYoL1AdhP+833Y+vr
dRduv5ftF68mssJzgDJNbcRVI2tG0yk3Mj0QQPzu6uF0C4i802SXCScf62b0QxnNzh+rQvlJKi64
BScfY5l0t2F8P0dJg+o2BYl7fHdjqq0xv4N457ogWNI3g/rzIesppN69sg7kj0dV2gnU8p1ak1vu
rtuBjuPTySUh6mCFU+UITgL4mRjlJNZjEr1wHsUWNUQxYsrWeRDUT3x9mFUgS/hmQCLKppfSleK9
xtH/CjFdCXSpkdyFVn4l7V2VWHJfkTpMp8l14f80cSYwrfExm3kQ9169RzXe0CTbjZfoV0FHwedo
ppaW0eXf0qrKp5Eao2DkecSlNDcME8RlgNenlubPD9SZCjlcAEg4bfwxiBbTxUYOajOru59O/HSk
FQ2ojm+H6pHY9KNvrZq34+2djO0gVwsMYgJZnxmgsyQStWaqDfNsv+uV8zvKYR4WicwGChv6Ijwq
SfqE+s8DVxkmgby/u3kUNXwhytrGBUw8hW1t5v/Vq1RiOsd84aO8taB7f/aiSHH8wEmiOc3qnbWg
xx9OJBM8RWyD7+4nsYpNbzOQEOj6yhvjrrb3TEgOgS9y5bCPfAhBaNwAKtYeob6z2fypnq/LI/9e
Ed7FRsJCh+cO3ufiA4p5uJ5NQBOde90j7Lvo23BCDXG0m5AesHULPWYlPuo7VgFW38aimcLsyHbQ
CjuNh96Rpn3E8QDGTu8Io0X2M1+QGB04jIX5FtFaQa+6z1ELqPlHOf8JQVOUiS8o+S8vk4NfQ57F
UvlA7P/RU3Lazay3+o9cY+hNHF3qaBbY3KbiiPHtW45OiFiGhyf8qQcDnG2c0A/c2ysQoqz/iFdB
X0H51T2Zs6KLci7N9e6yrhA/sHKRVh5DB+jG8ORBzzWlmlXfHXIVO4XCiSyLs7uj97wvoCFPlqPL
SoUv/SJi0iJiHB4cTStVmsJj3krEQHMf93Ym3d15PtMgI5FyRlIWi8SeivKw6IyqIv8DYZetjKei
t4KCUzMRgljl7FygJLAdECWSGom81VFPWpT4qv2FoNL5nJCf6gMuYlZJT7/qtA/xxObhfBans5vX
/p9XXgqYBHOFeP6TAKojZqhJS/w+ZLx+R00GfpNoljFqoGq/P5QipsmBv1a5Ij6RyqtF8iJ3QOtx
IJmBAW9QZUSIevkXXW9qdRO1yOAb1ItnYAJBnNx3V7WCXhJZMQUGvnxr2G8YFVh2KKHaamB7z3WF
MD2qUr04ZmI1q+sV3UXe/YmJN28vQ/WVY+ignUeJ9RDuz/jpwxVikXPFPpGhUwc3sHW6k8J3eho9
7byUBdt52PJ44sX0KpL3QY7rhCert3yyRUtZ2+6fP6lAN4SChGSlU5lTAG3WqCOhsL3Eg22tNeUt
2fwzMLe+P1qa7T51NVblMEQdnZTNCvTxP1oP+OEKC8Eby3Jgpavv8r6ekrjC/MOrIof2F+aOxNjA
IgzMsWElp0zYqGqqvJJdxyMmajdKKB8dlEKJTeQvtoVjOuxYxI0YnOKMvlrk2TK2AIW5iVhIHf1m
AcR/Gtpt8XVjbkLa82v1J1w5ClZuBWteC62VONMRASfG4dtPntSe1ERYlBU3yRsDUqH0wXBhaHSt
EjZ5TjY7Wb89KwwklUHtYLRoLZRcQDNP61AZQ/CKCqEY3mX8oQ1hqRKSu71u5JBCfPDVR43QAcIM
Df4+N7VpaUgByOlPh5sYqpHGMRcG53lkNduR70k4/bb05MsN3JYX20MyTPS8Ai0yp++IboU7vGHi
FUkZjtmz1VIzEEXpSmWE18jFLrKM4ZrDT9+fN/sbABAEvouWDEXap+H3WabyYmYKztf0BYVojhlJ
crnmqBJbz3yjmhsgQZ2EVd8GVQd9+L2wbbMUewv0ySBy5Ms9r0Az613wekAGPvCGwIhnF67gTadT
s60W+RtqjkRowDCrmSBCJAe2SRhs4Hh3ipfjYzzwCUxfOw7bUnBT56WnahGp2R/58uJ5eLHBMeBw
/AObNhhuCFur5pBxDCIGzMs+fyV8l4wRHeiuzHYYQrhncVIF1aKbhsOL4UU8h1KvZwBg09qMQIjE
Nsn0iJ1KYizZKH4MwwuVwC3J5SaaKwznq7xMZkkl9EdipD8+DycPtj9L0c+l8UJLi25fYVK4CtVb
IjFhz4QdcsKdbolONhLy+SuIk2UQxJ0veMNdgo4BGQ0oJt0YMpNJt2wRtm4UKYuTGMtByCxgzdxQ
HRwsJkt66oLydQd66HczIrjwkARNmUuqfZf1qbp+TrwD3wzlNcksGS95QNZKtaAI6/Hm7s06VOI0
8SNzbjzxdj9aOvhlNd+ekrJhSXXTtEVs53HL42NJf9kh7ZSG4F/4Pc0AMfb1AnTX5btRm4+vlbQQ
Epds9Xvi649qqUQqrEmED+ot4Ov1GYuxNnhO9JgjYytYbBKYINL6YDrwJuDJIMZapGxY92pDrYQL
2gXJ62gXEPlRgUKzI2/jvtVUjraKUosYgxKBuQKyBCJ5yK2XLTanM66CXnjyqI3594O+pBPGRa00
VNAJf45JysZlsKexM8/aDSdYshvCB089uKxnRW5NgiYY0MlQZb6hGoCtsCmAcbEU668F0mYhJgBX
PRWDD5fqwXZ/0cbE7mn3csk5LACTzTtz7d3ny6ZCgMuz0Ut0kTlQ1Dz5y0QE7vzzBamQv1S0OaP/
xfPoGBU6YblvfEnlyeZyF0YFlc94DKC5SQAB2V63SX5JCYtoLeT+MacLIIILa/fJnYMjNmUI3TmG
cOrJ5JbxR3tm9J2pojT9UxZsdiiuampvHjglY7SnwhSCdDXT+w394M32ErhvM+ZWeisNinjP/U9X
jFRDDhGauUiMR2zJ7kLQ1fFW8QpBrBNyA87Z3EkLdDR7VeOjbYvqg23+DUwtl40Q9R/Xgqae6ImT
/UOJ9OSN65Z5Xyl6+KJHpj4qT1JHlFTfKRIKppoZQYE9e1qNaw2hpZoK7oRwHocN/n8gd9p4tpoX
hP3ppjyZHNDEzSNg4gJwRt7FagqZ3g3XgvU8MQzdvYMcI3racPtk7/8Q5wtVefHqiwDvDoWR8BcO
I7DGk0q/cHRK8AO+LbFAd4pDwNvo+wwvVZvrtZbNqNeiedN8e9jGkGUgdgsoKAMWfvaocF9txYSQ
I1ymktVTiW/AvTdxbVgZuXLStYDhi2pAVouVLwcRXVN4ohJsxXBk+bbCKvDqJUd6AHxGf+GCtKR1
0W96tCtaXtwA+mSuvU2RsHE9QbRbUwopXJH4eCuCrN4SWAN3cIyYktpc4bbc8BE9cF07t4av+KB9
LG9ghA54ZubydqAGheKWRfX03ZFAJNpd0UIvMwQhJfcGbHahDYXrGM2sqJJgukAUKTve0T1N6E6A
q4QzlEl89FXLnbsPSzJSgCFc2WhgCduPCyszZmScgqyP4dzsvaIY1V6539H5E5b1BA6bV5Hs9b5Z
ndWMsIzueB6Ps56cCCG28UlclzbslrVZ9ApqCJxs3XFvBsTPVwPUvysxfEeoQvTbfW0wDfsKcXom
T5SyZZaE6mj7T1IlzrrGZofUsHL2NT8Bqyq5IJCAibwQlem2rI60zJXeOW7w/rWpRHR3RKMHFOry
4Fay8volwi+NumOp48ZjhtGAuQX2h8fjUw0Qjsm3Lq9F/MdfPRzicvlCYW8QElwuW4zY0IELRdAA
ugamB1C0otVqZLuAX2bKjpD2pZp+bk5lc+rOfbMhfq/2ovTdgek+7Gz1Q4TRMUOZNWK190nEVIL+
TuFWNWWKwIa3stndy7BXYMVW4Rz4lrd731+TXMk77YAO2PwaQ8HZL4BOdRrkRaVwfYm68BGkXK2H
xDOZmiVo/n+a/CUHqUZPCrQSts6YMbEjEabvCT6Gr6576ir8qE9d+pPfgu1etzDFpaEDw1XxwVqk
+Pqwm8awcswMGlWKfVDmoabJRwlOdpPcZpRIVOB3f7cBRt5n1HOHQ8kZ5sKezDUMb2JAN/1MtM4o
ptqh+sdQmc6QCxpSCIUaZS5Tpbbc4gszc+xlLo1GVdE2+miuAI+xtYugNkU8+VaSbDvxA+6KO6Ef
zIvJm509+Q8Nt8COzbTUpTDdYhJlg/0t5HI79Hun2W7qXezTxaGDZP+LCYCOAJxGLRNuNwi4c0sg
KL2IRjU4rJ8kh6H6OcNFfZBasBEM4B+QSw7mnEfHTZ+zGPopUN6XkgE1+y5pJuf4GYCuDebRKpYU
rW9A/+/KMSenWCoALJFElniiHeyIRskuufFm9c2fKE6Uyyy0rCCJq+aFBuWFH+yoEQO889LHoTUz
tYUgiRVEz1rEFswq1lm6wJ5JCgVSOJi1ymnWwOHRuf4CFXuptJqs6I1hxwnNc6c1hMwQ/aQE16ej
u6QV/2sU9Znjl571ONGnJ6YzzQb00aSt7hIME1Zg4ZQR9dTAyNOkzI0aDc6qwprilMhnmDLioKUd
U1+i4nl9xMvO9z4nDWXOayq01oYozEXZyGU9G7q4fORWSY5vqyB1m6gZ1L5/im72B71/u6//7Mph
tPD8fi3irHwj2+piel560mPKoK45F2Sa72Qw0aRAjnej9CpBV18WHjYuahjla3ViRSibK1mCqq4R
56ppfrnT9tce1y8gnQrupsOwkjiIBr8CQMZVeuTHIfk15IMHT5lyJWT7aKRBLogN1/wOCuLMhuHM
rFE4ahCfvDhseeeJABVPpBl1YvZlNk8CWKMZqCfJXhCIA0QYQv2inJ7ZJA6/y0QDVT0i7X+txm6t
B4Gc5E56uMvJfWu+G6UHqKOmVvrx5cd0KjCUtYg8MhOpV+L1J22bTh/EUlD1Yc2MhCiqr+brKvoQ
oq9bc4ljNCyuUsLQGfl9rT+f89kfMxz5Id7TQP8wrt40FnHA0KLGdqip35KSsbZDA+eA20vAT23J
Mo/O9QrMOhUmDQfdUN2TTAGq52hnCAwZ2zjxXncYYnvVcYFEVysb2ttC90BZzQMARl/Dtgmx8wDH
FUtqR1PmCTP2HnmOYDVF9pdeb2KZlh1iJAxHduwhjdveu6s09Wn4GThcSNCI3GKRGoVbJwglOBXr
6nn7pFnrFrXAC0V4Eqin7Gy+Br68W6lQAwKAFyQ4LHrOekTCeATgILvkOQb8aWFCb79uHYXP6Fqx
rVF9IGy4HAhk3/zzFcEbiq8Bvs3gOfkGCiozgacAL+0mFHVo6GUrDebNCZAqficRPvoqR54hpZcm
dz1QiMSzPGWe7pZPGkJcVBCBwQ62T1BsQgaHODeFhtz+ogmo8Ab8kJmIecVc5i9KsFZIsTyx44gk
YztWh+ZPJ4+dntpwdw==
`protect end_protected
