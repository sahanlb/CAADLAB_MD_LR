// (C) 2001-2018 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
P89TBaMmHh0f2L/gKiqgq5htduYuZifOW/tkjD/qPY9CFGCqflVkSnRY6G+NQbwVtHPCs3SEw6O9
piu83UolTFzryPY3S4n63eC7LxGvtz0pT5Fsir7/JQAO2/Gv4HxVHqSfYbnHES/vxDWg3R5hFhBJ
zRKxlJWD6Kn14ZIYiHYI+3ezlvNqwxO5KPAEuDL0jqeJMaoyAmmUE4jkQXy14JUnp1Tq9eVkdsrj
YdyPJbE7DvluLdyVpi+6RKDhKD0eqUtszRfcH1Smn5qy9PWF2gU59eNQPU5/fkMaYc5bn5i4s5tW
1bPqr+Ozum5tNEET+luqaax9EZH9SmXz77Er/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11008)
sPkuSWidHB5vb4BEQ7/gkyVAqOJN9WV+RINk3nPWP+qzP54YhG7ioGRWSY1S32S9mo9Qn4Hpp3Ba
QxvtOO9Xu3pPbfctXU4luccjBUt0HgUkDahYTj9ZcoZ5w0HlOgNh25oO1njZzOPVl2KxPaAeTr2y
G8X/1EgrxxHMtQ1DWaDu+/P6AlTqqI18aVFwgpRm+Z87fT6DqqATy/tj5r6cSO2215quvgPN8Xlb
JX19u5iR4QqqpDO8LTUbOjJJhL4LyYEyig9DBCZ5v6TSL7LQW9IjlBypnUaTSoOMok055CLO5vxS
0rIWaBrcXLmQ9hksZZ65uslsrG7gMVYudxuTmS5EplgtqTiNeyQlEzVVXRjJCAxvq6sjPmYrK5w2
k4ah5qRyuMD/0H38SART7Wlf4PqWsnYjTVv2TCEv31CDL/jXpWUrQGpBg1nyzARakyOXh1CJXGdw
ees1VY7wWip5AnRXt8jW5a/8681RNFhCwdOExXD5cN1lwjpbNFf2BVKiH9ybwkLx9c7pyBM+UPYZ
XuAG00bzSi1T6SV9nZcAgigK4qSJksePoLrMSF2gTUS9DnmPq4dZbatcmwHjWMMpIa2YCnckRm1K
Duzk5XU4Q7ptsPGvUG2X3mhRjxMY+emC9BlhO8nizuAoskYl5dpVPeU3ZuUrwRxHLZy+scvNSPKr
Yym0LzrdCoP1yoQ4RowZfGrtSzDEhMa10AlrT0YANBcKmLYn0uXapqYP2jY2ODknBzJbo/MGoxGa
8qUH1i8AlM/NqIkbvkqw/+fogRZ5n6rty7GX7AubZFBdL3BzmqtmkbeTl/B9y8iNsDvqNI3btLiI
FE1vXYfWswLzBr5bBYUh3HbgD/PKKpy4yeiSswt1cWttIIwfCLARVRXbZf6pA/izrpPGc+XWrUop
AUoCbJM6B5va0cFqBbLGZPoOB4+kGzSZaCLxg21lSWHvI7ptaEM3a+i+35EGhnnuZYfgfKv9qGuI
bRs+mjEYsL70P6QoRoUww+eWSpGkcomNoB7ajmqLhlM2wea/bXEd2yYvlxjUdDlxqBSKk1YCrDtk
fhsGJDSjC69NdIyvazXQNbEIlK2P8pnWDTJoPxnUQxHIWvaXG53PoHTqkU0IVeNjldE2danBI6F4
LwT3gjg10N/WZHhEkyuCE+7//zob4epmD6oaM2sCtxMhCGXXOVcuZe9rVRkFH+Yen4GDrxa0khop
0lqTrZ2Y2Vwf3uCI/hTmgPUU0HmhGeBUsKEZ8Jyck0apWjA0bwPgC/UqFzlBHFDW7Xv4TLyI3ieU
l6XU0iGsnDQgKXd6TW3Rtb02rH8k1rhjCzORNz1kQx2m/XLUy0B/+8QFcEhf9RGyu9ORKIxBxgyw
pyS84Vh5a0n21NShtBO+22qAKxKkklwlBQpooIXmGjOhO+LqoJvtIKsCtdJD85qOzkxdUA+8UM/g
wotV+y347XeDlQjm2LuY2lfhoVmi2LoKySo7IAXrwqPqyzr8QsxP/XkVxBeOzfk3P9JLI67PK2tT
gvxajb8vjvgIa8h6URhLr58f/lt6JNcAYHI8ji976i8hCI6g5EFyfATDXuweVTJbLpEd9P7RqR7t
k1t3JmCfpJcSyr93B2t/sw3nkTyNUXHiuNt7LSQAr3ynEMgyYAuA7johWhXXuoFnyufLNkDJKdg/
E7k+dAo+3lm9S4vn/8gc/TuvzOz1mES1oLKvVvwFlRcB/3X/6eMUL6poKwWuUO0y2A+jlrtQ4eG+
bvyLOWLILEkd7O3PeSZSqsdG+EgAIJpWlCQcdP9Oeha7sZfCO1o9qiH7u1oy9zc+xHqtgrZUdcsF
P57AHPIcmi8b1/Qr0HJoeQSoRQEuLYArqvbjbP1dUdVnZxQK670365yNYYBVVu6JRTeNDh5vbw/U
piCJ8ZY0v+twlrQ/HCgx6uMsNRBjn09dccVHVJCcUplZZ6MJJ0LnLrqnYtFeZ/IZlxDC6WBNCQAD
27VDclqk8f8WKOtUANgRsJksqWPqIG0PLcFRf1jS3WqqKc+zvbj0n72FNjV5GDMyM85+kS6gWPLq
/1xZ1nVzMwuXTE+WcmguK97YFZmbBel3gGSzTUnwPvcVWFWEA+KNhHONJm+TS1yWR8hSTIy1DAlw
TbnRemG1FyyS1Zg+U673JKvrxM1WrLmXmZL4R5wqpkEJo5HfDzwDa0lbKuYdVrb4EqrQMyRPJSAo
891A4ksVEqlO8oBaBVmchlfbsh9/5BKkWOaJP+C+AlgPwyrDk3wdwCpYyEeQ5kJsJTu/Egg4NheF
68qxvd9brITlH1dxgZZCB1MHqjt+ILPBoPwinOiz2kJM90Lv73kVyIZTXVJJ5u1t9aLBJTc8OEq3
1URZN55FHdk8Fev07qYPP8HPWrI4WnCSlXkUS6AVtWXvfqWZo4ojZa2c8L5kVSTlxdbXS8tkUHcN
KYWIAXtqHA+4g4Ok8DInO7xFhUa8+VzfH8JkVdEfx5YYBnKrNUhNvL17qkLlVaBO4gejCRp2WmDn
qR+oNfCKBEM8v8ea1Y7MVDUQoZQsAmmIwkUWnRoGCCoFxFkm0vZwoknPy87dwc2RkGtCg1t98FjY
iCIN3f/NAznHlitth1uC/gEplOt4udQ3l0tI5U9Zip37OXbIp2G7XdfZHS04XnIe6wxtOBGFT++M
GbUx7SVfAQmY2nIJvMqe6If+oHut3YastcaWQtRMpZj1NmVd82Jaxz2X/D2DWBYAgrQHKQfs/Jgz
Y4pzBEz5selir8uITMojlQyQ/iU/tAQ6hI49vsoHsu34Z3Eulrmvg0zGngTRIwEG0vMgAWfbHC+D
HTpbw3PhCOHVYXMYKXYDFCNHD1Yc0fas1/L5HGtxd4AfudEu+YX3glY9uX2HzObL0fKM3WCNMCdY
3rRdV+XIn09d45vxAY/zdPURszXlZwTbEHa5Nyfl3EGdOPz1MOTDg0lfZiaHVIAKoHFOKQWvG8Bj
s2wTomcWIn+AKOM9aiPHPl3AqEP+r77d5WMR/Lh3HakquY85WLErPb9owIBt7qxp5kfbKceuIojC
f/xPSxfcvt6BVf+6g/79NjLHqZeGghsvXhzOOV4hIO+GVMmTWN/DGyiDXCEaiVPfsMAidl+DAaeL
rBMlhZhLowF6d1GpwSVn2QLdqAgQgHks/7aadGlceIfh/ibMRKo6k+w/m4wQ6KCIKdpXkONeifg3
0rdXEFvvFZqA9y/kk7NNEoM9eLvFw1KFIzQrToJgm0yBEu04SqFR7G9W2/8Lh5/sCOUhiXzqASaX
nCpfdxCWy2+AqAj6wf73CvNVS50knfXvqpZaQCfuTIab1lU/G4r8xuF7o3jIxIv8IeN3HBpvdM/u
V1nIFj2CEyU390i42EuSqhazPaZHXHC2QG1pv8owC2nKm+28D3BB0PzW4bT4R39+UCI9L82amnVQ
Hv9UgF3nq4s+FI5Yt3LGPPh1/5Ul+n39QKwOXAZPdzu6vL7F0hErOw91ZqvMc0xE1OTcLRw7upTQ
e6qvjsh2ist2rBFKWN47s2guSl3Y85/0bqYYeptHJwW8dcUTUaz7S2te3M6mGgmg0tUKGl7LIpnh
+VaS+Vmg0IEdWuWrDimTp4aNLO346Ht1FS/JLSnQHsbCsQfh02CksV3aFVeTYxe3J18z/3GRydQ8
dnud9Cmzm2dRixEish24l9NkgPfaIWlBt2EAH6Cr452FsAnFPQM0srZqZkonwe/uhsT7jnUBGwZL
Y/yU4YnlrisUuL3oHve0pqEP3ggPWRgkenFuCv2dm3Clv7HyAEtzwoYzO1LqFC4DyWq5F7yyOIil
1M/cbKR8+1Kb+FbNXlPVSWjmkDkOnieQipgNcrtvuhjKdaBbjkZRu5rj5TTkxIF6VcaG4pTKfD3F
xaPf5z8FA2FVyg3I8tv+IZQ9OrwPfPvnFvuSszCcHG6zfnM8BrBmg/Ez72WNIH/tHsj+NoOmwH5D
C1gx8Kk54JR5EaPK9sU5Q0DfXhJJsKzRB3xtJAVCIhxx1OCsJe3BSroy0pM9+iW7ciCJhi4H3xCd
4PPqtWMQ2hpofW0e5LjNF5z6weHhjfPY8TtGY/t90LrJDV9oq3aKeF6X/+1MfI4BJi2TioOd6BCE
KUXu9cQyvz6eUwo/1s1T1E9gR1QhOZCtfN+V2t+Ox7E6K4itsqHFuOiMyyrj+G6YmvtjninvH6CK
KeHN/dq1W6+Ub7wi/8wb60wuKm0qaZILIOcmDVtHCrbwWvjWf9HnUwv7XLMgjeAxEdgHmfVn8XJj
2RblvmKARwm+zdksG7LrVqvy3YNR65U51YnuqKgg1oCMiUP6FPeeb70AGtTtyA27EFEonepFliQN
z3/X0Z8jVL8gE4dS8DMT9xjgUwEEekG16AFRM6xDpwYK7X1OxfYEJdT4btSi/6yzppkIkIU3qahb
P1/f/jjztv1VFdMhL8bMgwoPL8mmJB5XrBi5IhhNXbxZbDdz0rj8N2vLQ46WL+SsWgs4ZIt7n3jn
T7CVXtQx3qqOyyR2Cx+Bl8YZuLZtIN7tNVRlxeTFnluGqNkWeIrD03RkETHQdwWD0cAbmzMdRpkc
TuuJpHKqZ3cUOB5vwNcnkJVRkDxsutCTjUTpHeN1lcODsF6eeReCVYiNB+//cAst9w3Qi+fwb7/Y
/Em++eBgXaHS1pVZe+wiGd0ZKnw6eQ9qRdQTDGWs6c4/K8m2FqbO29k68EYEH63OzTxjSTUNKScf
R4RC3IlGGJNRBBcnJAhvflFInRaqWcA+4Yb+pYly/xEA6k3JsPma3tF1feMbBhSOg+xBSyE2299T
sD1+gOOFP9lCz29Tx4HpbbpqRHREigHVl3toVKoKkw3rwEwiv630UIJHvvcQaFwL6w12q4o9hBdp
p1Dp0uQWLUQdteVyCb/rlJFXMMpcfkT+3PPPdY6I5G7d+LvCukwCT1+PqHTbPbId8XPNn5Va3RUM
wLOdP4cwf1Jp/JYsz1hRbJ662Bu9fV9FiKov+JYLvOnF1TBBZzEY0i2qhg1joiPmBnzikU91XZAd
oWCTuy0GaBDyFwK5dElNBy3UQpgP5iZAYyoZsmE6oO0eMMet7TF89u8S78JFtUgpinUVOp60QbTN
Wo2EDVZcgSI5owIKocyE0Bj5yQi5GoPTCq7zrTuCdjES80BM8Pu0McwrJ781cwHnBJzJWM84I/Fq
bA98iXaEgI4O8AIvXz/ybR7KOA7oGYG0m3zg8hx4v9mrv9sfceEY0Y04vGeE3eSakHK+v5tRqxI+
89ThIhiY/p07sn663Nkyh3dP98CbX7t4I1NUHdwEWH++rJmPGofnVKUEk0OzngwDp50EG9WeurxM
UJfqQMJF7EB8ANE54Zx4TB7Si+VuguKiXiN0ILXDIGzFXN1goNVIkHIABw4QHhIT6ZRKvMpHwiVb
oINzZWUtCRkh4oBWzJ4pZWtgl4En2369oYlRP0IMjNYkWrTsN5m4mx4SdxlhQIn3GmXzDYY387QJ
jzbPenUOEqb29M57ZCE+s61clmQHi5zr61slav2ZKcnZVa3XIWbW+sYvrHzjIo9Czbqo+o76b7wI
Cx7w0Hdt6LC6Om2J7Y7aT/S7Bm4W+m9y6/i4VlvjxKUIi2EExE4oxzCcCjeWB+LU1ccWrTSGTJcS
u9gV2+9eOFmsn8IH0EmyDivoyZW0xu6K1DO2ATpPa0Ezu6lA/HeoLh1NdQNEovuF16uu510nQD8K
Vl/QwPMhk93yAJEV2h478zvPDvVa+kBjSEc++3eJ2oPt4AruYB8BT5zFklF/H2Rsf5dJDhfBx1lp
jW3yW++Jj6Mr941Gm857zm+srXX2iUTSff8D57OSpf/uFwOmJMlBG2iRIpG7hyl+H4FqWKI0PbQs
45QM47Kc0Cv2sKaLHBK82QcDSVb1fqpHmNjG7HMzMUGrQJ7mEq3AsUYDg///x05C7GkW39piqsdQ
N3avWMZ35P+WYseSmb9vR9ZkwXzauy0/g7kp6NuDgEcgZCb2ivp0/D8aXbhGrzNM1ijtIVARN/Xg
l7qmgYGtcpTxRj+tVhPKQUKjAI6B3hxvXIQC5J+HK2nCJVPu076DyySSx2cUF51qrjkiW+Rs5prU
KTvq07ygWkTcPnKAz7/CWEcUYNjgcfMTTNrdj6Gl1myp7FijnjpjBkJKOo2U1eqxliBFNJzEe4ip
F5v2K8QhFmmmpGGazTVILaxuAny/AtHy7fQlUKJQzljtXlKTdsZZiuhrvuoTzKMteiremZXB5lhv
76thRgmdMIZ6ldiD1vEN75YwCezLaXjuoit3pNI67oV8ZXxMdc6plLDcOp9nmXOfIyibJn6DNSWt
s7K8ts859BeZqKt7rsNFFsjcxcyQKPmjJHOUyCFsHjiRJUeAODtVvG/bK67nOgXpcYj9NNKR6Rme
ldQCc6qniJ8M8MAnI9MbDxTOs6izvZBZygpGtrxACFuGrvit2b6wxPZnevIjLRRa/M1oSdAFeqYC
bADxtPBMGOG+3q15PvKirRRgF917QWjbfqKJ4enMMMGEv0gpUHrUyuRLfM08VU9LNFHrV0TMl/q1
eZJ2cVLBuKs7gP7TfPIj8JmYPH3/iVQqtCrOhjnTqmke2dG3mRou4D9zLq7KF7cu8FJ4doaP2ZCD
D3vCiOM7ZewxHtKx5HUOxGTLnEgxzbGp3Gzhdb96cz9k9jdVG9RMI9hr/eB8Y1JKcu622+lbjhLA
uWBu6bS+ULVGDHXRj76rpcGY8WYZ315DaJI3eHAylI8bqs2Rr8wpu9j5TmD/mXRrWqvbfQZu3i0I
ES8YG9QDFkpUhf2qC1XkbmZ9qmp4fJoiM85SKrj56i8kmUD07dac70tEAiWJXPnvpHuObemlBJz0
bjwPOaOLdTpHH3IIWL134HXnV/TJwqYLCqu7QvgcFZmKgHRm/IumpJE+XVjHGt5LVA+BZg1422Ci
MwCv64XIFnnCK7vas80BFZPOW9vXYDgdhhmQ1uDMCN9n0DpYv66LtVqlBY2hI7PrHnvP0AZctmC8
C+zT+ROo+XXT1QvhnUVX6pQDvAAOIjCnSQJZrueX+S8r/KBRz3J4sxBMrHORktp27KyoTjzoF5ei
B9PpE1z29IQv7Wc22Pfg5Dq5YuG6tBwirA9eimAFsZYrkdqm/vSwIG++9HuPF3oU38QTCNJwHoCc
VjwZ+8rx5wrTR1/fGmaRhfhfqARw3ZWL3zdpl8mHTOo+eeSDSZ2apNaESfRBCTyJb5YxSI4HK5Yb
3Vgs2Fg33X4q0Ixo53j91Wzor8NqS0Bbh9RfNkAfcd1Do+uFOl33Myu9dhIpKtNeT0YwyjcoDppn
oaRAWq6QVOo1ZrB964jx8O+22vKR4723my9HptxgQRFT5aTUSWAXRCtFm+87/vLB0g9pU2eUIAV4
byaM3B0at8Xt5yq1GLt3J6XV2HmaepbB0wgNArdrFh7ppkZldStZ2ZwlAsP13PNd/eXeoffvs02r
h8oZ4D4J+RNMOmkEmRW5GA+0geJIoKF18i/a0TErSiFdMVNEQLluW1N344ZqeNLSm6Pytv1nXFIS
8z/WfnQexrI73xtOkPCyWdcj7NYnbt8bNIxWJFd9CqFXPueWm0AO6F0H/OAvjjVUDJykanN8YH+s
EJbD/bU4rlWeAXO9UYasUsvvAUZnPmx44X89Z+QemkbO0pDRD0szC1H8uoOPtjaZZBYbuv6A0/EZ
XLcpYJthonfPKd8QpV7FxvZyR4T0jMIukrEv4wYACuc1LjkYVdPM8I8f5huXWtXGLs2FaPhmXalP
Kb1Ffd07/wCw4BKZHl6m25hmtuuy9pwpf4w54mWGiNMobLN6j9nguy9AjCbB5o1MdwjXcvAs2by6
a92qr9cx53O94lNYVO0ZBlNsdBBUyeC7U40z+iuj4ZMRix1ivkxHlhKjPlle56tQnJuQYBE4DArK
Pf6J1uePCAzdrydrk/o/9+TedDOiAAkyI1r9lkKmvt6s3EdjKV/943SS1O4IFbVdPes43fhGRFaz
nvVXgv6LEpArSjcPUiS4tN/Emy3weiCLNM83eF97MPXKobLujzHcFR8CBvj7D3qZkex5Mq5Ed8az
F80A0iVjsOnhB6pdntPiwpNABkiDv95NMBJca89nqzTSdUvCUKmASU43XV+Tyx0Lm8+z/KyMy9zR
ZMLYpt1Eogba+eep9ExpHe6jP8YANcS7PTIh55+/PAvybaaazziBdiHUBd8UqTiYej02eZTT2d+w
7IK15TgZp7bvJ9xIi/FIPf9gqkmDW+JUOZANp9XEboUHhQvk/YzBoE3scuya/HqibfwNy5fdAU2/
C8o4JM2Y5qmwvnWxcYLinNqj8+IiLqD5sdlE64TrbFtp1Twde7U/5PYEunOOssEvbtqALINWM6aH
EMGbcKwEbdNcBYdtVmaDR1oyVrUqR4SatM1tjCTxe8xtk95z5vxDwBxAAmzrVGEV6XFzrVbJeG4n
6ZH39YBPibzs3OmFOyRSZmyi0yJL1wqf2GLfBy+5oU/Ocyb/TQ41OjxMKy/9z8pjE+j2WJxMnKpG
tuc0U7uqeC3conknRsf7DvPvoFCGfofkkkBsKzm38popSbzuVXAtHDQKdyPdpN8fHO2RUGZ+nZw1
mwZfs2SCqpsj18iT3v5eQkruv2M0fMItSqEuqkR/M6z2xd8fKKpG6XWMSxbNr6leexLf02p8HU46
U4eASbzsSjsBYWP7sVvx4tUdFu6Wg1DSSsjzmsSEXI9ObsLBm9cDFx1yP2ITLhfdFNjnbeWlBlJD
CdbJ3Bju63mNsypvN1X/3xQNCLfoYWxkPFel0vmbA2sdT1VBRjZBUdSe+lBYiumfvQM5aKmJkZQ9
tUG0tKpxitEXAop1resgtzTm/s/QXVytLhyVaDsurszXlDP5imJoTa0UTmSeGV4VaGlyAliGEQDz
d+fvCnQ5WmkYUUxWb9gSq06DjLfiHSdN5/gBVgT3rGAmSD+SKxv8704i742c8/TMD91pmFKwhS07
UTsqe7hTAEAO355j6WVrdi1kKe0cycfQw4n58UvupNYVKaWX8fazNHnqRtlwE7CTztBSD2PKQJUy
f4AyhTaLgyd51oMwCRGQanfRjfS0SrWOLqoITkpZkLeoTZLbv6NWDyWxgmBcFd4GgUfZWLs3+4dM
zpqdBKW1qzMBlRah1p4waF3lP8IU5c/hmzazrysiyrpbsqEOABvviaz6zhYnh7G9yntE8ai0sZAg
qPcoH2EYVlkVJEj9l6p5Bkgam57UhzEE99vrp41lLTx7V0IttQofzMdiI1YMEv4NQOoPS/LOP3g4
VO4a7wKnJuXzlZ13EzoLVkMyvM6RpvASNtPpD63Cz6JMZTsXtVurOyhzjHSo9kMWHxvRC8WXMfeQ
wtMhubaOseN1WP8vPHWeXFU09YXo0246YC4tvJcwYDrED0sY5vvg2HbIfFZVNKeSsXUeN3v7BaqZ
8gzpYcXRx7yM+m0KL33dp3xxhcnJ+VClb+i4h1o1gz5NTgyviPXrxirMQr6Py6oqTWnt7sKAHPiR
kYDZeYaMsa8f95qVf2uV01zynYrCQK6o3kt8NP5DjzDvnp3wqU35SssC1z+cW70RYa0q8MC4lQiK
DrjX5zxUHwxKYXooJzbHnOf2EJ9mVIiiUzzqG/5Qz1DAZRulaMTL3amurXjQNm4oxtP9bvu4F7N+
tKTSfRwRLNm/TTc/8zDF9tZC+jk7ltDYVrnk8XI5ITul6m55PxeJbsIOGW/IVfTErjaSJU/hkQbW
ihT87yQYv8DNw1tvThJ+AK/DcDikxgMsW9GeTFA7zc5yBBmJnc8xBZbSOb/JYLOFJ37KZBvtqLsE
+dh+X0kFIBfDrkoSh54S0a5J+RkNQJ067sJxe0LZi/VYqi5cXTbs1Gv/dIS/fzoPFVDEgtXaYmEg
SingeLmd6TQIBnuXHM9O914K5OFm+dH6M/GHjsqmkp4JonwoIqco4BZl4w/jwiCVy2tirvnmzpD6
mse2l/wXq1NLAEuBTtCNmp8zf4elVAuA3u8bNlInP4CvTtESUcVoO1WiMtipTR3oi+brk5O2rdtA
BOOQu+BP5tjCUshWDDIV2k2LuVQfLzr56EK5Wf4fnLfU9hAAYpTwIMXjNDLiCR4meKObTGlw8plN
pGalr/TA9Y5pzc4Dx1uzgaXmXOLXBMeRv5BqM32ByMSDNdHhgzmfo7xio2WDNA8Upnis/hxFwhP/
dnIN2zzC/BlapmoQNJaY/ooyCGTIFl8f1cU1M/VlRHA3sw7tYwAUaOlg/2gsVzzllJ7QF0F8DJEE
3Q1JiJEaT/tXAOCMxg5stwtwwErbUol0u6/ToVY6TR/dtlBCIgSNQnCkhZ0avkBko0PwQdHJdO7k
d/yvUGzz3otXLSBDwVA/iZQGUEOps7XTo8OWhPG4RGm81iGYejQ3cxGb8jOl5bF2fzDdzdGyKtF6
HVn2VH1alK3mCz4wSSSlaRxdDu9EZdX0jTNxpiWn2/zSPMI8DcfDtIMGpVtxLl1v5ChUAGxlJXiA
zYI93Y3JoZkgdy5GvBXkH6+3OYQmmkqFfxeAq8QLqC6NAu79FuZFp0JUErRIL6kZuEUY9ztq/hUF
DN99rbfvMQde1JHXDzbI41AG7lABav8tFYSka+Q15xwIaOMf3xCybS5nFLdg8Ob1L7bcnQVR/u40
Jkx2WADQvkUass++vhNL2286gxwLTz5DZxDqEWYwPSKuhIvY8cmHlsCTbS430PcZo2JQpkZlGEfZ
d8kSlU8ro6Y0Cfz4NhmeR44HSZ5jFLfsPKZ40Tt8/9Y/5ROOEQjrchsfCobUZIpCQ/QK3w+bhqOU
TUoJ8+MBT/6vU74a+LE/foZF36hRdArP98btnvXoUYeQqiPgS9lupVtQqu+4x+uLcVi3o3T4BArE
cZ5h3DExOVicXrx+foyZY389R81CyBSRVY6QpQwUYeg7k8FSq3HEOY+NUdkxf4OvGGCg5uL7Bhid
j5KA65TetAqeLCgh6qU85laaAoToy88z0npXrMQvT23udnMwTeXxWUkqdepCODDg6A3wRojRN7uc
vBS27sY6nbbNq0msls4q5/EERoxwo4xjxsNBVkY6DzH8zZ3cqFtqClg4PJ/EGKpdUYeF2xyOn7GM
bMc97+b0Z0WvyEKMsuAKKkR6zYjgP79JPpglHyJh9Zq2NMF4wA+WS1CPwIG1YF01DBHy2TiBeXoA
HH3Y7BFRXmz/yaJp2ywjSm8DfvXFcAIDQkGT2OsUarbbdDkRaiBos7TRz6GnhNHb3tzqp6dJryWq
/DnhdUsL75R33vGxN6oVvS5nfHiH97S/KkQ34KCu4/BaI+efMY6p+W381RvuP4Df4DaYq5GT9NOz
OMb8ppmEPBRMZxcYz75EK81UcMiMWhtus4Za0uIG4yPUwaYyDtymzqKKJ48G4peKCe8bn/c6rEdW
Ve9h7Giev2bQTlE4WRlLNlJh8kvKvZOAQjkSA1gLcJmaI6NFMhR7eDOvoweoFwidUqNtfGuhKYSd
BZ76r3ekx+wjYup31ZSqZi7H+zocq4oIJCWkSTT+ScQOpDEwRWpI5sd6ud20wZt7XMkNrGg73972
9vahGZ62rlmwKsG8Pd/0iDxpyFc33MAZVZztwWRxM11QhfyMA1BvyCCj4U8tKh7YNgk63OjAWowQ
V1bhqsOeh/VcVvJZSoOz4SJ5NrhdovoH1rpk+MW6E36v0Pny58vGEOTP7+AFeUA8uH9g7Yfjo4ag
3AnV8fgFCDH+505cvBmMuj13eaAmYpY25AQ9WpBq61uA7FbsJbzd8gx8lonaCHdlMcOzUOfcw6rB
Fr60k/DjinpOe2n4jIAhSCE3JzXV6gGmIy7BYrKDA0CsRW2y8MiJPiY0U1BGzRf8dKVWyaud6D5B
nOO3yjV9CAIuiyKkk622pTKw0sLYrfzKIPyrtStKhSjYrcCuoUUIjTFNusL5RyuAH82dxjPnPFVE
g0v01a5h+Ial4Zl7ilP6nz2a/35FcLtnLZefZu9hSCv4lhV7s01r1F3WXV88p0Hj/M5DxRokrdac
WvAa5J+XdEc/sF5fvSPiTJBkHV6vRt3KvSQUjtD+oIm9roRWpgK0I+TDYpIYVkXN2W3PATM4C571
pjPWHyfMGQztHbySUC0I5iauYeqkeJ4muZ8ajPU1OiHxyXMC4q4wa0i4GtT76SaYxqmhEs+/fyda
kmDRfOqnbz4zHWkTOhfe6RmIgccN32+l4pMeHVXjfiUudy31BYYeiR7tbK4rvnugnLGAuCGKlDjM
LFmuUjlnwzaaLu0hZ7FNsGf/oADnc3OgLHGSxz2EJRSwZeFN+OduSV/Ztr4jSu40qpjLMGSr+pB5
CjX3hf14+YmmxI/GV63traB4kWGVwA4bChd/4Ku7cQxjsb/G/Yk6pMPmNsdPjvNZvzkUokpnQ8jP
cR/sdtFv2Hn55eVZk6xtfFIs5ej+WLVpL9gr9OYdGjJHqfxeqJgQ9J6j3XNByEhwrXdKTdZzB+ma
A7llbYzmAsQAW5r13moZmbgRW2B5ZBWhI2X9XPZm/M25zqxjMU3UWqmAUZCvYbmF22m+9Pr7NaPP
Rz1CANg04aGxR59ebQSTvr/8qInaTE8qGV7+l/siw5YDiQOg1kewtHdSntviMmyyvas2luAMaqsG
iyhs2dkmt4mF7tptA/bkYbQ+7AnIb70wXNuq2bm/Ih6EgBXTBKuZ5nGbKxL1PWJTCu0nHJYFCOKy
uONlkiSAW86gpPp2tMya9hftqgNFP2fhPVbh0uTj9k48QzPmIehDKXQkMMCS9ZhhxPIXDw/0w3BB
sjLt01j7o7S4AL4AnulSTga3bZ1fmYA1m4o+floCZnf1iRnuxWRhLzxl5blY+e/JIQzPB/bJj2+j
kefY91CNmMsfDQFMJvvc8mR7ekag3CqAfvnfq61pk6RkB4RDz3zbghFmpDZP1GfmIWb2jgsjQBXd
5+FZOtJ6hWkB3DxTN1MGK3N4dQnTOl7pzgcsCmlEDAj1dwd/9wHGstTNZJRI0K92gAouVBwKOLiM
v4gxxdM34ETHC/czfUhctE8g4sUp1TVBBaQa4G7EHzralmvi2aXmjUGiTPe9z8wRbOipte1xufVB
bXoHczJksk8qInjIsUcfVFNx7ybdSl5Wf1odJIQ8oX131fLqSZG3FpdzAlcKYPf27DClvEewCu9W
44XmtrR6lW6DiNGJlQqCVPEjWgI48miE+LMHFoPrI0pbYjRY2Nr7qylg2amytcTVYF+0elaTzX5/
mAedDh6iHBQnWO91KQifiidzWSien+/EMiUIyD0RBACTE1Au39f5PWCh8Gqi/Kgfam3C+bx8gZLJ
BPzHoXFlk4MtN8ufPdfAgB9/bDs8hLDeTOaIQnRtjSle87uq+8T2ane4EpN4O+PZeuXrsTly5MEQ
CPwT3lxLxxkK+yFYXRB9pq1OPZWX5hdhfircTSAn4EUpdxa1zlbYiytmaL1rQzIz52J2uRFWh3kc
Y9klhEv+LYjFjoy7PypoeJpSK8Kvv/nWgF6KCXczHbhjkP/sn2WcDMJU4uriDzItus+DqDflM7GP
3wKddwXLplcQEhQ4zvMHPLjrOqCH15kYqKxfyUXZRPpRX92BihPaiVD5LtOf0q3m97o812nlu8OL
bs7V/uOxV6cDRzAlpdOz5AYHY+S/xiOzhSuaFkh+hEl/2Gd6KAjCU7m+u6Fpqh+J1J/VL1Oowt+X
Ul1PrD9KZ+kkBNpBc8E1FMzQN3EPwdJ4K4uO5DkdmVUz3xnx9edYRcmrAT5j+KihUgoSz/ZV5dXl
8fBtMX/JH8BcLekVzglTDlBbUaOIOlyivs0Cq8TDDdWwSSUOJsGzGMXpZdnpc2yYhq6lWPVxleCI
CIaQSxMspIgY8XXhC5SstDoc2qjXgbnLJk0P0sBqlBu/eo253hhAHHNnoh+n1XsE7LINfo0QseBV
FnxMzcIG+y8AjEm4bXXPNHgK8ZLfb4TvfIMd/JqNBvpNt2HMnni2TbKHMZ1c7jhgFm62PYKNaKTZ
VbrAt6bSpc7RngL1WjrQS3l+nGGwXWgXbbvfvUobu01k1Ssywnx/7T/pGvN0Lrdc8kclHI9DGbpz
MdiA7hDx/fUsWsTZ1QMZMYOKTlM1jDAZPkiypG9KWHuTAS1+9F4cpBWQx3VYWHu3VHmHEWWT1sm2
TkpU7m+xMI8DpSa6/afhUilV6AU0yjFew7PNe66zSNDf09QpyJX5bsm5udoyXgpJRn9QWsvBpAE9
sLpku6cVCHrupSGZ20sYb6V04hjq9AUDEH+0/+3JtCxGEVfFvkmg4t46pHTFMxOiYYJ5hg3pjRkI
D1kKMOBx9KVMytrPRjKGszf6ynz7QodZDFY0Mw7qOzBG7kZSq6CCXqunb2WpX9QEHgs0Rl6kiVr/
xJerCSxCMjx2VvClxMeVESS8+ZrhEti1jMORLWV9xM9NTd+012WkzaBzO/nrfWeHzYQmLX6y/TwD
rh0+ShvX3VzMNTu8XErEnD9SzHFXdrDwQmwxVtJx5pSh6aSWcv7EOAcji4LXFQxyQ93xHgNPkwCb
Px2Ts8bkXV2TB4OZCuIoLDu8F5xfKO4/MoXX+wmEpzhdmXym4zkYe8XhD/eyPD3Hke/SWd6R2Yzp
UlOdo57t9d0VID02vnSW+bwpSKjJyBpR8GscXVOTUubogLNDe5bagoA/rj6N3Vxy45AezcQM/eFn
/rvYno1YBw==
`pragma protect end_protected
