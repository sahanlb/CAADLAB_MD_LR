localparam [GSIZE1DX-1:0][GSIZE1DY-1:0][GSIZE1DZ-1:0][1:0][31:0] GMEM_FFTZNG_CHK = {
  {32'h41bde247, 32'hc0321e23} /* (15, 15, 15) {real, imag} */,
  {32'hc1df0ca3, 32'h40cbe9b7} /* (15, 15, 14) {real, imag} */,
  {32'hc1dc5023, 32'hc047d6e7} /* (15, 15, 13) {real, imag} */,
  {32'h3f510b61, 32'hc0ae5903} /* (15, 15, 12) {real, imag} */,
  {32'hc04118ea, 32'hc0ea1cad} /* (15, 15, 11) {real, imag} */,
  {32'h405c9995, 32'hbf9c4a4a} /* (15, 15, 10) {real, imag} */,
  {32'hc08b8b18, 32'h409deee8} /* (15, 15, 9) {real, imag} */,
  {32'hbf261c20, 32'h3f49637c} /* (15, 15, 8) {real, imag} */,
  {32'hbf88dc7d, 32'h40598e5c} /* (15, 15, 7) {real, imag} */,
  {32'h400eb278, 32'h4087b00e} /* (15, 15, 6) {real, imag} */,
  {32'h3eb94449, 32'h40c7560b} /* (15, 15, 5) {real, imag} */,
  {32'h403ab2e6, 32'h40490cee} /* (15, 15, 4) {real, imag} */,
  {32'hc013c98b, 32'hc18b5f4a} /* (15, 15, 3) {real, imag} */,
  {32'h41deecc4, 32'h410c5e8b} /* (15, 15, 2) {real, imag} */,
  {32'hc0cf05d6, 32'hc20592d9} /* (15, 15, 1) {real, imag} */,
  {32'h41707117, 32'h411c5a46} /* (15, 15, 0) {real, imag} */,
  {32'h40b96ba7, 32'hbf974c27} /* (15, 14, 15) {real, imag} */,
  {32'h41d44b9a, 32'hbe00e7e5} /* (15, 14, 14) {real, imag} */,
  {32'h40b46c87, 32'hbf357254} /* (15, 14, 13) {real, imag} */,
  {32'hc01ca732, 32'hc03cc774} /* (15, 14, 12) {real, imag} */,
  {32'h40d192f5, 32'h40888162} /* (15, 14, 11) {real, imag} */,
  {32'hbfc5b821, 32'h3f97e5ea} /* (15, 14, 10) {real, imag} */,
  {32'hc0a30357, 32'h4023bb01} /* (15, 14, 9) {real, imag} */,
  {32'h4073e89b, 32'h3f1884a4} /* (15, 14, 8) {real, imag} */,
  {32'h3fccc00d, 32'h4041d99c} /* (15, 14, 7) {real, imag} */,
  {32'h405cc1cc, 32'hc05c16f3} /* (15, 14, 6) {real, imag} */,
  {32'hc05eb9c6, 32'h4045362a} /* (15, 14, 5) {real, imag} */,
  {32'h410369cd, 32'hc02a8b22} /* (15, 14, 4) {real, imag} */,
  {32'hc063679a, 32'hbf3aa381} /* (15, 14, 3) {real, imag} */,
  {32'hc0bd7b2b, 32'hc0a6208a} /* (15, 14, 2) {real, imag} */,
  {32'hc17f7e0f, 32'hbff85c38} /* (15, 14, 1) {real, imag} */,
  {32'hc0f14c72, 32'h41b222f3} /* (15, 14, 0) {real, imag} */,
  {32'hc12586f1, 32'hc0e42c79} /* (15, 13, 15) {real, imag} */,
  {32'h41267575, 32'h40279acc} /* (15, 13, 14) {real, imag} */,
  {32'h40a26de8, 32'h408ce1fa} /* (15, 13, 13) {real, imag} */,
  {32'hc129a6d0, 32'h40d282e5} /* (15, 13, 12) {real, imag} */,
  {32'hc0b8be13, 32'h3f003f84} /* (15, 13, 11) {real, imag} */,
  {32'hbf172679, 32'h409e840a} /* (15, 13, 10) {real, imag} */,
  {32'hc00c4cae, 32'hc0132ba4} /* (15, 13, 9) {real, imag} */,
  {32'hbfd1de4b, 32'hc04fa946} /* (15, 13, 8) {real, imag} */,
  {32'hc044f5f1, 32'hc03f0733} /* (15, 13, 7) {real, imag} */,
  {32'h3fe4a302, 32'h3f6d9f09} /* (15, 13, 6) {real, imag} */,
  {32'hc0c397f4, 32'hc0808795} /* (15, 13, 5) {real, imag} */,
  {32'h411e427b, 32'hc0909893} /* (15, 13, 4) {real, imag} */,
  {32'h40dc9bca, 32'hc08c2f64} /* (15, 13, 3) {real, imag} */,
  {32'h40331f45, 32'hc1203c61} /* (15, 13, 2) {real, imag} */,
  {32'hc15b4b0a, 32'h41ba5cb3} /* (15, 13, 1) {real, imag} */,
  {32'hc0477230, 32'hc0d3282f} /* (15, 13, 0) {real, imag} */,
  {32'h4114d7f1, 32'h40c58b5c} /* (15, 12, 15) {real, imag} */,
  {32'h4037b09f, 32'hbfc730c1} /* (15, 12, 14) {real, imag} */,
  {32'hc0b5ac32, 32'hbf328b6c} /* (15, 12, 13) {real, imag} */,
  {32'hc0c9541d, 32'hc02348c2} /* (15, 12, 12) {real, imag} */,
  {32'hbfb3a4b4, 32'h4011e30d} /* (15, 12, 11) {real, imag} */,
  {32'h408af906, 32'hbf909b46} /* (15, 12, 10) {real, imag} */,
  {32'hc080e49a, 32'h3fe1273b} /* (15, 12, 9) {real, imag} */,
  {32'hbf5491a9, 32'hc076813c} /* (15, 12, 8) {real, imag} */,
  {32'h40b87411, 32'h40320f21} /* (15, 12, 7) {real, imag} */,
  {32'hc081cdfc, 32'h4061ec00} /* (15, 12, 6) {real, imag} */,
  {32'hc0e83509, 32'h401ac7c7} /* (15, 12, 5) {real, imag} */,
  {32'hc10690d4, 32'hc185f5b1} /* (15, 12, 4) {real, imag} */,
  {32'h402844a0, 32'h40ce9738} /* (15, 12, 3) {real, imag} */,
  {32'hc0a1aacb, 32'hc0603e81} /* (15, 12, 2) {real, imag} */,
  {32'h41375898, 32'hc0065711} /* (15, 12, 1) {real, imag} */,
  {32'hbfbf33fa, 32'h4108ac90} /* (15, 12, 0) {real, imag} */,
  {32'h3fe5ab1b, 32'h4018ebe2} /* (15, 11, 15) {real, imag} */,
  {32'hc0e401fd, 32'hc00abb44} /* (15, 11, 14) {real, imag} */,
  {32'hc004c169, 32'h408aede6} /* (15, 11, 13) {real, imag} */,
  {32'hbf803fa6, 32'hc04900a2} /* (15, 11, 12) {real, imag} */,
  {32'hbf458b22, 32'hc0d27050} /* (15, 11, 11) {real, imag} */,
  {32'h40379a7f, 32'h407a05e0} /* (15, 11, 10) {real, imag} */,
  {32'h40a9b909, 32'hc0b3a25f} /* (15, 11, 9) {real, imag} */,
  {32'hc03fd695, 32'hc06f41e5} /* (15, 11, 8) {real, imag} */,
  {32'hc0bfeef9, 32'hc048d11f} /* (15, 11, 7) {real, imag} */,
  {32'hc045b7de, 32'hbeaf6185} /* (15, 11, 6) {real, imag} */,
  {32'h408cf11c, 32'hc110dcbe} /* (15, 11, 5) {real, imag} */,
  {32'h3e644b44, 32'h3fff9367} /* (15, 11, 4) {real, imag} */,
  {32'hbfdce858, 32'hbe95db80} /* (15, 11, 3) {real, imag} */,
  {32'h41278eb7, 32'h41567416} /* (15, 11, 2) {real, imag} */,
  {32'hc0b27248, 32'hbf0fe108} /* (15, 11, 1) {real, imag} */,
  {32'hc03703ad, 32'hc167ef7d} /* (15, 11, 0) {real, imag} */,
  {32'hc0cd2b2e, 32'hc009f0aa} /* (15, 10, 15) {real, imag} */,
  {32'hc095906e, 32'h3f296fec} /* (15, 10, 14) {real, imag} */,
  {32'hc119ce31, 32'h402ea9d9} /* (15, 10, 13) {real, imag} */,
  {32'h41676393, 32'hbfcb1dbe} /* (15, 10, 12) {real, imag} */,
  {32'h4110fda0, 32'h3dcd2d7f} /* (15, 10, 11) {real, imag} */,
  {32'hbf64d309, 32'hbf9e8efe} /* (15, 10, 10) {real, imag} */,
  {32'hbf5f3723, 32'hc09163a8} /* (15, 10, 9) {real, imag} */,
  {32'h40294b3e, 32'h40bd2d8e} /* (15, 10, 8) {real, imag} */,
  {32'h409028ba, 32'h40761289} /* (15, 10, 7) {real, imag} */,
  {32'h3f8b9687, 32'hc1120e4a} /* (15, 10, 6) {real, imag} */,
  {32'hbf5d2a26, 32'h409eb4e2} /* (15, 10, 5) {real, imag} */,
  {32'hbfa0d6d4, 32'h40af63ec} /* (15, 10, 4) {real, imag} */,
  {32'hbf072e2c, 32'h408fac98} /* (15, 10, 3) {real, imag} */,
  {32'hc06fc600, 32'hc053e090} /* (15, 10, 2) {real, imag} */,
  {32'h3f5d9414, 32'h4009d5a8} /* (15, 10, 1) {real, imag} */,
  {32'h40bc13d8, 32'hbef5e5e2} /* (15, 10, 0) {real, imag} */,
  {32'hbf18370b, 32'h40a24c45} /* (15, 9, 15) {real, imag} */,
  {32'hc00812b6, 32'h3eaf119f} /* (15, 9, 14) {real, imag} */,
  {32'h3f58b232, 32'hc0211ffb} /* (15, 9, 13) {real, imag} */,
  {32'hc074784e, 32'h3faa6967} /* (15, 9, 12) {real, imag} */,
  {32'hbfe2038d, 32'h3fb4ad1e} /* (15, 9, 11) {real, imag} */,
  {32'hc0fef844, 32'h40227cf1} /* (15, 9, 10) {real, imag} */,
  {32'h4020733d, 32'h3fc844eb} /* (15, 9, 9) {real, imag} */,
  {32'hbe2edcee, 32'hc0014a8c} /* (15, 9, 8) {real, imag} */,
  {32'hc10abbc6, 32'hbf83f683} /* (15, 9, 7) {real, imag} */,
  {32'h3fe93910, 32'hbfaef098} /* (15, 9, 6) {real, imag} */,
  {32'h3f991fba, 32'hbe9aca32} /* (15, 9, 5) {real, imag} */,
  {32'h41200e55, 32'hc0061b25} /* (15, 9, 4) {real, imag} */,
  {32'h3fa0142b, 32'hbfbdbf81} /* (15, 9, 3) {real, imag} */,
  {32'hbf55c174, 32'h40018b11} /* (15, 9, 2) {real, imag} */,
  {32'h3f9b5826, 32'hbee69659} /* (15, 9, 1) {real, imag} */,
  {32'h40517ede, 32'hbf949bee} /* (15, 9, 0) {real, imag} */,
  {32'hc03d7005, 32'h3e893fc2} /* (15, 8, 15) {real, imag} */,
  {32'hc02837db, 32'hc02207d6} /* (15, 8, 14) {real, imag} */,
  {32'h4018435a, 32'h401304e9} /* (15, 8, 13) {real, imag} */,
  {32'hc08b1518, 32'hc051cd39} /* (15, 8, 12) {real, imag} */,
  {32'h3f88a884, 32'hc01cd6cc} /* (15, 8, 11) {real, imag} */,
  {32'hc0d59027, 32'h401ca943} /* (15, 8, 10) {real, imag} */,
  {32'h408d5388, 32'h405b11a5} /* (15, 8, 9) {real, imag} */,
  {32'h40162360, 32'h40573852} /* (15, 8, 8) {real, imag} */,
  {32'hbea5f3e2, 32'hc060494b} /* (15, 8, 7) {real, imag} */,
  {32'hc010951c, 32'h3e7f02a7} /* (15, 8, 6) {real, imag} */,
  {32'h3f641087, 32'hc0b06acb} /* (15, 8, 5) {real, imag} */,
  {32'hc0457b78, 32'h3fddc49e} /* (15, 8, 4) {real, imag} */,
  {32'hbf72ae23, 32'h40bef5c1} /* (15, 8, 3) {real, imag} */,
  {32'hbfba2c1c, 32'hc00fb3de} /* (15, 8, 2) {real, imag} */,
  {32'h3fcb1a54, 32'h40236276} /* (15, 8, 1) {real, imag} */,
  {32'hbffcb177, 32'h3f1d66e1} /* (15, 8, 0) {real, imag} */,
  {32'h405b3ac7, 32'hc086f4ba} /* (15, 7, 15) {real, imag} */,
  {32'h40823ccd, 32'h40925735} /* (15, 7, 14) {real, imag} */,
  {32'hbf96780f, 32'hc011f99b} /* (15, 7, 13) {real, imag} */,
  {32'hc00b9d4f, 32'h4123b09d} /* (15, 7, 12) {real, imag} */,
  {32'hc0473e50, 32'h40a281eb} /* (15, 7, 11) {real, imag} */,
  {32'h409c42d7, 32'h406ab150} /* (15, 7, 10) {real, imag} */,
  {32'hbf3866f2, 32'hbeee0ac6} /* (15, 7, 9) {real, imag} */,
  {32'h401e7118, 32'hbffb3e92} /* (15, 7, 8) {real, imag} */,
  {32'h3e82a052, 32'h40da7b01} /* (15, 7, 7) {real, imag} */,
  {32'hbfda9d01, 32'h40344056} /* (15, 7, 6) {real, imag} */,
  {32'h40504dc4, 32'hc0a58469} /* (15, 7, 5) {real, imag} */,
  {32'h3fdb716e, 32'h3f9767a5} /* (15, 7, 4) {real, imag} */,
  {32'hbf903a25, 32'hc0d81fdc} /* (15, 7, 3) {real, imag} */,
  {32'hc03b033e, 32'h400fbe16} /* (15, 7, 2) {real, imag} */,
  {32'h40242b69, 32'hc0180647} /* (15, 7, 1) {real, imag} */,
  {32'h408970fa, 32'h402b9f8c} /* (15, 7, 0) {real, imag} */,
  {32'h409e8ea0, 32'h4102bb7e} /* (15, 6, 15) {real, imag} */,
  {32'hbf11342a, 32'h403fcda4} /* (15, 6, 14) {real, imag} */,
  {32'hbea088e6, 32'h3f3392c0} /* (15, 6, 13) {real, imag} */,
  {32'h40f64f95, 32'hbf9e82a9} /* (15, 6, 12) {real, imag} */,
  {32'hc061bb61, 32'hbf2564c5} /* (15, 6, 11) {real, imag} */,
  {32'hc10f43df, 32'h410478a5} /* (15, 6, 10) {real, imag} */,
  {32'hc098b84a, 32'hc0b0a5ad} /* (15, 6, 9) {real, imag} */,
  {32'h4094ebcc, 32'h3fd94971} /* (15, 6, 8) {real, imag} */,
  {32'h3ff4aec4, 32'h4078e20d} /* (15, 6, 7) {real, imag} */,
  {32'h40641174, 32'hc0b9c4b4} /* (15, 6, 6) {real, imag} */,
  {32'hbf5a5287, 32'hc1122c94} /* (15, 6, 5) {real, imag} */,
  {32'hc0ea0a2f, 32'h406b8147} /* (15, 6, 4) {real, imag} */,
  {32'hc01f44cb, 32'h41138482} /* (15, 6, 3) {real, imag} */,
  {32'hc0714624, 32'h3f593dc9} /* (15, 6, 2) {real, imag} */,
  {32'h40da0d27, 32'h408cd47c} /* (15, 6, 1) {real, imag} */,
  {32'h4062734c, 32'hbb75e187} /* (15, 6, 0) {real, imag} */,
  {32'h40ed19c4, 32'h4087b427} /* (15, 5, 15) {real, imag} */,
  {32'hbf5d1fd1, 32'hc0c9c918} /* (15, 5, 14) {real, imag} */,
  {32'h41534b80, 32'hc0d0aab3} /* (15, 5, 13) {real, imag} */,
  {32'hbe676ef6, 32'hc0d375e0} /* (15, 5, 12) {real, imag} */,
  {32'h40bd7e27, 32'hbfad10bc} /* (15, 5, 11) {real, imag} */,
  {32'h4004948e, 32'hc094776e} /* (15, 5, 10) {real, imag} */,
  {32'h3f5aca9c, 32'h40c23cea} /* (15, 5, 9) {real, imag} */,
  {32'h3fd751d4, 32'hc0097d71} /* (15, 5, 8) {real, imag} */,
  {32'h4094e041, 32'hc0aa1eeb} /* (15, 5, 7) {real, imag} */,
  {32'hc0a249f5, 32'hc0c29dcb} /* (15, 5, 6) {real, imag} */,
  {32'h4057c435, 32'h40d1dd6a} /* (15, 5, 5) {real, imag} */,
  {32'h40141083, 32'h3e8687c0} /* (15, 5, 4) {real, imag} */,
  {32'h409bb0c2, 32'h402bf1e9} /* (15, 5, 3) {real, imag} */,
  {32'hc07f7777, 32'hc02decec} /* (15, 5, 2) {real, imag} */,
  {32'h40200a48, 32'h40cc41f6} /* (15, 5, 1) {real, imag} */,
  {32'hc0a6826a, 32'hbea823d1} /* (15, 5, 0) {real, imag} */,
  {32'h403fed67, 32'h40a0cfa2} /* (15, 4, 15) {real, imag} */,
  {32'h3fdd00fa, 32'hbe86a062} /* (15, 4, 14) {real, imag} */,
  {32'h3fb2dcd1, 32'h3ffa6ae3} /* (15, 4, 13) {real, imag} */,
  {32'hc052d8af, 32'h3f2acc81} /* (15, 4, 12) {real, imag} */,
  {32'hc08a5e39, 32'hc07e8457} /* (15, 4, 11) {real, imag} */,
  {32'h4052b2da, 32'hc011c2eb} /* (15, 4, 10) {real, imag} */,
  {32'hc0006ae3, 32'h410d3b68} /* (15, 4, 9) {real, imag} */,
  {32'h3f919c30, 32'hc01fcc31} /* (15, 4, 8) {real, imag} */,
  {32'hc1138209, 32'h40268790} /* (15, 4, 7) {real, imag} */,
  {32'hbf81e017, 32'h3f0b8d06} /* (15, 4, 6) {real, imag} */,
  {32'hbed09a51, 32'h410d8a4f} /* (15, 4, 5) {real, imag} */,
  {32'h40aa60a0, 32'hc01406d6} /* (15, 4, 4) {real, imag} */,
  {32'hc0513a4f, 32'hc13e8a88} /* (15, 4, 3) {real, imag} */,
  {32'hc17fe5b6, 32'hc10ebc4e} /* (15, 4, 2) {real, imag} */,
  {32'h3e3e22be, 32'hc1bc2cb8} /* (15, 4, 1) {real, imag} */,
  {32'hbfb3db82, 32'h4145ad77} /* (15, 4, 0) {real, imag} */,
  {32'h415ce201, 32'hc0195597} /* (15, 3, 15) {real, imag} */,
  {32'hc0cfa381, 32'hc1689415} /* (15, 3, 14) {real, imag} */,
  {32'hc085eba1, 32'h41894841} /* (15, 3, 13) {real, imag} */,
  {32'h408c5cd5, 32'hc04992f4} /* (15, 3, 12) {real, imag} */,
  {32'hc08ffeba, 32'hc01353e8} /* (15, 3, 11) {real, imag} */,
  {32'h401b734c, 32'h3ee665d5} /* (15, 3, 10) {real, imag} */,
  {32'h3eb4cd7c, 32'hc0c516ee} /* (15, 3, 9) {real, imag} */,
  {32'hc0187793, 32'h40c9bf22} /* (15, 3, 8) {real, imag} */,
  {32'hc06ee97c, 32'hc13e67d7} /* (15, 3, 7) {real, imag} */,
  {32'hbf023d0b, 32'hc040f249} /* (15, 3, 6) {real, imag} */,
  {32'h4009a0dc, 32'h40d8a038} /* (15, 3, 5) {real, imag} */,
  {32'hc11e07fb, 32'hc0233346} /* (15, 3, 4) {real, imag} */,
  {32'hc05f091e, 32'hc1752b0b} /* (15, 3, 3) {real, imag} */,
  {32'hbe693de8, 32'h410fe12e} /* (15, 3, 2) {real, imag} */,
  {32'h4135f285, 32'hc035eecb} /* (15, 3, 1) {real, imag} */,
  {32'hc1206f34, 32'hc1821d47} /* (15, 3, 0) {real, imag} */,
  {32'hc2398330, 32'h40fadc0c} /* (15, 2, 15) {real, imag} */,
  {32'hc1b973aa, 32'h3d65dcb1} /* (15, 2, 14) {real, imag} */,
  {32'h413e86a7, 32'hc1652d93} /* (15, 2, 13) {real, imag} */,
  {32'hc08ae559, 32'h40d1a150} /* (15, 2, 12) {real, imag} */,
  {32'hc08dc219, 32'hc0353925} /* (15, 2, 11) {real, imag} */,
  {32'hc08ebf62, 32'hc01ba486} /* (15, 2, 10) {real, imag} */,
  {32'h4116d5bf, 32'hc0eccc2c} /* (15, 2, 9) {real, imag} */,
  {32'hc02b7db1, 32'hbf7d2119} /* (15, 2, 8) {real, imag} */,
  {32'h41268b1a, 32'h3febc4e1} /* (15, 2, 7) {real, imag} */,
  {32'h4016eb31, 32'hc0e67d5d} /* (15, 2, 6) {real, imag} */,
  {32'h3ffb74a9, 32'h41027f09} /* (15, 2, 5) {real, imag} */,
  {32'hc10e6733, 32'hc0550d16} /* (15, 2, 4) {real, imag} */,
  {32'hc08a4217, 32'h40d3f94c} /* (15, 2, 3) {real, imag} */,
  {32'hc18443a9, 32'h41d189af} /* (15, 2, 2) {real, imag} */,
  {32'h41dfff9d, 32'hc194c48c} /* (15, 2, 1) {real, imag} */,
  {32'h4105e123, 32'h41bba2c6} /* (15, 2, 0) {real, imag} */,
  {32'hc174eee3, 32'hc217a280} /* (15, 1, 15) {real, imag} */,
  {32'h41c14442, 32'hc1a2ed52} /* (15, 1, 14) {real, imag} */,
  {32'hc0dc6e39, 32'h40e0b850} /* (15, 1, 13) {real, imag} */,
  {32'hc0801ab5, 32'h40b95c54} /* (15, 1, 12) {real, imag} */,
  {32'hc063903a, 32'hc0b84dab} /* (15, 1, 11) {real, imag} */,
  {32'hc082fd01, 32'h40c2b7b4} /* (15, 1, 10) {real, imag} */,
  {32'h405eb8f1, 32'hbfa3cc8c} /* (15, 1, 9) {real, imag} */,
  {32'hc074933f, 32'h3fc49775} /* (15, 1, 8) {real, imag} */,
  {32'hbe254606, 32'h40f72b59} /* (15, 1, 7) {real, imag} */,
  {32'h401c393d, 32'h4038d6f7} /* (15, 1, 6) {real, imag} */,
  {32'hc12f0083, 32'hc10d2ab0} /* (15, 1, 5) {real, imag} */,
  {32'hbe1cf784, 32'hc0addc6a} /* (15, 1, 4) {real, imag} */,
  {32'h4107c53a, 32'h404e7503} /* (15, 1, 3) {real, imag} */,
  {32'hc03d76d1, 32'hc196b22e} /* (15, 1, 2) {real, imag} */,
  {32'hc0f281fe, 32'h41056a1c} /* (15, 1, 1) {real, imag} */,
  {32'hc1c7ee53, 32'hc1aabbde} /* (15, 1, 0) {real, imag} */,
  {32'h4114ee81, 32'hc2ce4ee9} /* (15, 0, 15) {real, imag} */,
  {32'h418b1860, 32'h41d832a9} /* (15, 0, 14) {real, imag} */,
  {32'hbe47a2dd, 32'h41b9de55} /* (15, 0, 13) {real, imag} */,
  {32'hc063855d, 32'hc1009e33} /* (15, 0, 12) {real, imag} */,
  {32'h410e07e8, 32'h4084e3a0} /* (15, 0, 11) {real, imag} */,
  {32'h40f31cb1, 32'h400f7172} /* (15, 0, 10) {real, imag} */,
  {32'hc0f52ed5, 32'h3ef2501c} /* (15, 0, 9) {real, imag} */,
  {32'h409139b0, 32'h3f8d36c2} /* (15, 0, 8) {real, imag} */,
  {32'hc00264c0, 32'hc1077297} /* (15, 0, 7) {real, imag} */,
  {32'hc060875d, 32'h4185a6dc} /* (15, 0, 6) {real, imag} */,
  {32'h404fd7ee, 32'hc081d444} /* (15, 0, 5) {real, imag} */,
  {32'h41b13766, 32'h410662c3} /* (15, 0, 4) {real, imag} */,
  {32'hc0540f9c, 32'h401a4456} /* (15, 0, 3) {real, imag} */,
  {32'hc1072dcd, 32'hc20a5b8d} /* (15, 0, 2) {real, imag} */,
  {32'h420a9b30, 32'h424fd7ab} /* (15, 0, 1) {real, imag} */,
  {32'hc2395ed2, 32'hc2dd263a} /* (15, 0, 0) {real, imag} */,
  {32'hc23327f3, 32'hc19ade10} /* (14, 15, 15) {real, imag} */,
  {32'h3d23688c, 32'hc19e2294} /* (14, 15, 14) {real, imag} */,
  {32'hbfaac18a, 32'h414c955f} /* (14, 15, 13) {real, imag} */,
  {32'h402cf484, 32'h40c0a7c8} /* (14, 15, 12) {real, imag} */,
  {32'hc13b2cb5, 32'hc0327736} /* (14, 15, 11) {real, imag} */,
  {32'hc01aae7a, 32'h3e50bfef} /* (14, 15, 10) {real, imag} */,
  {32'h40b84a73, 32'hbfbc64ab} /* (14, 15, 9) {real, imag} */,
  {32'h3e2c0d4a, 32'h3e5d82e4} /* (14, 15, 8) {real, imag} */,
  {32'h4037dd78, 32'hc09f430d} /* (14, 15, 7) {real, imag} */,
  {32'hc100b4f7, 32'hbfc537ea} /* (14, 15, 6) {real, imag} */,
  {32'h404ac1c8, 32'h3f93e8ae} /* (14, 15, 5) {real, imag} */,
  {32'hc158b11b, 32'hc04ee17f} /* (14, 15, 4) {real, imag} */,
  {32'h413badbe, 32'h41a49a44} /* (14, 15, 3) {real, imag} */,
  {32'h411508b0, 32'hc06d83c3} /* (14, 15, 2) {real, imag} */,
  {32'hc03698a7, 32'h407e8863} /* (14, 15, 1) {real, imag} */,
  {32'h41aae521, 32'hc07ed176} /* (14, 15, 0) {real, imag} */,
  {32'hbff67419, 32'hc15149a8} /* (14, 14, 15) {real, imag} */,
  {32'hc0fde47a, 32'hc105ddd6} /* (14, 14, 14) {real, imag} */,
  {32'h4125e688, 32'hc08e49bf} /* (14, 14, 13) {real, imag} */,
  {32'h41844830, 32'hc149dc2a} /* (14, 14, 12) {real, imag} */,
  {32'hc08cc4ba, 32'hc02e9de6} /* (14, 14, 11) {real, imag} */,
  {32'hc110827b, 32'hc0c0f788} /* (14, 14, 10) {real, imag} */,
  {32'h3efcd575, 32'h413d4aca} /* (14, 14, 9) {real, imag} */,
  {32'hc040a2b6, 32'hbf338b3e} /* (14, 14, 8) {real, imag} */,
  {32'hc02c4d2f, 32'hc05b002d} /* (14, 14, 7) {real, imag} */,
  {32'h4084f3ac, 32'h3ddad7dc} /* (14, 14, 6) {real, imag} */,
  {32'h40563996, 32'h4129effb} /* (14, 14, 5) {real, imag} */,
  {32'h3f0ecb42, 32'hc02bf287} /* (14, 14, 4) {real, imag} */,
  {32'hc14ce3a8, 32'hc15ddf6c} /* (14, 14, 3) {real, imag} */,
  {32'hc1bbaff9, 32'h41722424} /* (14, 14, 2) {real, imag} */,
  {32'h413a6e0e, 32'h40990c4d} /* (14, 14, 1) {real, imag} */,
  {32'h40a9e51d, 32'h408f1ccb} /* (14, 14, 0) {real, imag} */,
  {32'h40ac54ec, 32'h3fa01c65} /* (14, 13, 15) {real, imag} */,
  {32'hbf05e791, 32'h3f821a99} /* (14, 13, 14) {real, imag} */,
  {32'hc13519e1, 32'h40127b39} /* (14, 13, 13) {real, imag} */,
  {32'hc10c95d0, 32'h40d1bb36} /* (14, 13, 12) {real, imag} */,
  {32'h3ff0fb35, 32'h40bd7de0} /* (14, 13, 11) {real, imag} */,
  {32'hbfe4c6b1, 32'hc0bb16b4} /* (14, 13, 10) {real, imag} */,
  {32'hc060afa7, 32'hbff20b64} /* (14, 13, 9) {real, imag} */,
  {32'hc0245e41, 32'h4013a146} /* (14, 13, 8) {real, imag} */,
  {32'hc0ad0563, 32'h3f716673} /* (14, 13, 7) {real, imag} */,
  {32'hc10dee0f, 32'hc0c32137} /* (14, 13, 6) {real, imag} */,
  {32'hc075c5ef, 32'h407a6488} /* (14, 13, 5) {real, imag} */,
  {32'hc0e98d0c, 32'h4073d71c} /* (14, 13, 4) {real, imag} */,
  {32'hbff17a90, 32'h4150cb25} /* (14, 13, 3) {real, imag} */,
  {32'h4145100c, 32'hc08b98a0} /* (14, 13, 2) {real, imag} */,
  {32'h40b47ad8, 32'h410538cc} /* (14, 13, 1) {real, imag} */,
  {32'hc15ebb3a, 32'h3e25193d} /* (14, 13, 0) {real, imag} */,
  {32'hc11ad0c1, 32'h400af0e4} /* (14, 12, 15) {real, imag} */,
  {32'hc138f5bc, 32'h3fc59c6a} /* (14, 12, 14) {real, imag} */,
  {32'hc1367c70, 32'h410a42d2} /* (14, 12, 13) {real, imag} */,
  {32'h40000b1b, 32'h3fb1696d} /* (14, 12, 12) {real, imag} */,
  {32'h40f4ad67, 32'hc064eae9} /* (14, 12, 11) {real, imag} */,
  {32'hc0dc2dfd, 32'hbe97332f} /* (14, 12, 10) {real, imag} */,
  {32'h40db856f, 32'hc03f5506} /* (14, 12, 9) {real, imag} */,
  {32'h3e06ccf4, 32'hc01d96cc} /* (14, 12, 8) {real, imag} */,
  {32'h40a61242, 32'h40849214} /* (14, 12, 7) {real, imag} */,
  {32'h4077456a, 32'h40f6e070} /* (14, 12, 6) {real, imag} */,
  {32'h4023fada, 32'h4070922b} /* (14, 12, 5) {real, imag} */,
  {32'hbfc66537, 32'h40dc84a5} /* (14, 12, 4) {real, imag} */,
  {32'hbf483ae3, 32'h405f6ec5} /* (14, 12, 3) {real, imag} */,
  {32'h3ff9ac31, 32'hc10f674e} /* (14, 12, 2) {real, imag} */,
  {32'h41192742, 32'hbf958c90} /* (14, 12, 1) {real, imag} */,
  {32'hc1259084, 32'h40370775} /* (14, 12, 0) {real, imag} */,
  {32'hc03d0a00, 32'h40fbae05} /* (14, 11, 15) {real, imag} */,
  {32'h41096033, 32'hbe986b2b} /* (14, 11, 14) {real, imag} */,
  {32'hbead2021, 32'hc105bae4} /* (14, 11, 13) {real, imag} */,
  {32'h40bbda2c, 32'h4108872e} /* (14, 11, 12) {real, imag} */,
  {32'h40454948, 32'h3fa8d4a0} /* (14, 11, 11) {real, imag} */,
  {32'hc131ffb6, 32'h3f8eac4c} /* (14, 11, 10) {real, imag} */,
  {32'hc0245a35, 32'hbfba9350} /* (14, 11, 9) {real, imag} */,
  {32'h3f9605c9, 32'hbef58fc4} /* (14, 11, 8) {real, imag} */,
  {32'h3ffbaef3, 32'h40da8be0} /* (14, 11, 7) {real, imag} */,
  {32'hc10b0155, 32'hc1839231} /* (14, 11, 6) {real, imag} */,
  {32'hbfa38739, 32'h41139ebc} /* (14, 11, 5) {real, imag} */,
  {32'hbfe21dc8, 32'h3fac9415} /* (14, 11, 4) {real, imag} */,
  {32'h406cb527, 32'hc123fc25} /* (14, 11, 3) {real, imag} */,
  {32'h403f209c, 32'hc019f228} /* (14, 11, 2) {real, imag} */,
  {32'hc0953ac1, 32'h3f83b58b} /* (14, 11, 1) {real, imag} */,
  {32'hc07dc4e3, 32'hc0f3d682} /* (14, 11, 0) {real, imag} */,
  {32'h3e456cc9, 32'hc0f8d03b} /* (14, 10, 15) {real, imag} */,
  {32'h402e219b, 32'h3f15aa2d} /* (14, 10, 14) {real, imag} */,
  {32'h40b9c3ea, 32'h3fa6edb3} /* (14, 10, 13) {real, imag} */,
  {32'hc0c1f600, 32'h3ff8ac2c} /* (14, 10, 12) {real, imag} */,
  {32'hc11d37a8, 32'h3f87fb3b} /* (14, 10, 11) {real, imag} */,
  {32'hc0841881, 32'hc1527f70} /* (14, 10, 10) {real, imag} */,
  {32'h3fd2c0c9, 32'h405a5adb} /* (14, 10, 9) {real, imag} */,
  {32'h40736640, 32'h3f8227f5} /* (14, 10, 8) {real, imag} */,
  {32'h3fe901f3, 32'hc1270ea1} /* (14, 10, 7) {real, imag} */,
  {32'h40ce4b51, 32'hc0b97903} /* (14, 10, 6) {real, imag} */,
  {32'hc13fcfc6, 32'h3ef2e0d6} /* (14, 10, 5) {real, imag} */,
  {32'h40d0bddb, 32'hbdd20eaa} /* (14, 10, 4) {real, imag} */,
  {32'hbf8a732a, 32'hbf9ac8a2} /* (14, 10, 3) {real, imag} */,
  {32'hbe547e19, 32'hbf92a118} /* (14, 10, 2) {real, imag} */,
  {32'hbff6766e, 32'h41028c7c} /* (14, 10, 1) {real, imag} */,
  {32'hc003b8ce, 32'hc021c4c6} /* (14, 10, 0) {real, imag} */,
  {32'h40157e41, 32'hbea30eb5} /* (14, 9, 15) {real, imag} */,
  {32'hc100a3ce, 32'hbe39d365} /* (14, 9, 14) {real, imag} */,
  {32'h3f4828f9, 32'hc0b8630f} /* (14, 9, 13) {real, imag} */,
  {32'h3f3891db, 32'hbfb7e398} /* (14, 9, 12) {real, imag} */,
  {32'h40ad562a, 32'h3f8af25b} /* (14, 9, 11) {real, imag} */,
  {32'h41557e2c, 32'hc01873bb} /* (14, 9, 10) {real, imag} */,
  {32'hbf47d0f7, 32'h40ab5173} /* (14, 9, 9) {real, imag} */,
  {32'hbf366e86, 32'hbe2988d8} /* (14, 9, 8) {real, imag} */,
  {32'h402aaf2c, 32'h4081d30e} /* (14, 9, 7) {real, imag} */,
  {32'h40aeecbb, 32'h40dc9d30} /* (14, 9, 6) {real, imag} */,
  {32'h409d43bd, 32'hbfd8ccb6} /* (14, 9, 5) {real, imag} */,
  {32'hc0915673, 32'hbfa139af} /* (14, 9, 4) {real, imag} */,
  {32'h4024ae04, 32'hc0458f0c} /* (14, 9, 3) {real, imag} */,
  {32'hbfd0b663, 32'h4031c66b} /* (14, 9, 2) {real, imag} */,
  {32'hc0157bcf, 32'h4014e742} /* (14, 9, 1) {real, imag} */,
  {32'h4032c568, 32'h3f7007e6} /* (14, 9, 0) {real, imag} */,
  {32'h409d51d2, 32'hbf035c99} /* (14, 8, 15) {real, imag} */,
  {32'h3fd40658, 32'h3fc011cc} /* (14, 8, 14) {real, imag} */,
  {32'hc08e87f2, 32'h4053c7cd} /* (14, 8, 13) {real, imag} */,
  {32'hc059c57a, 32'hc0ed0f35} /* (14, 8, 12) {real, imag} */,
  {32'h40b7a983, 32'hc037c623} /* (14, 8, 11) {real, imag} */,
  {32'h4045ebc0, 32'hbfab078e} /* (14, 8, 10) {real, imag} */,
  {32'h3e1b04c2, 32'hbfd6f9bd} /* (14, 8, 9) {real, imag} */,
  {32'hbf48663f, 32'h4011baf3} /* (14, 8, 8) {real, imag} */,
  {32'h40264bd0, 32'hc0258f28} /* (14, 8, 7) {real, imag} */,
  {32'h3f636953, 32'h3f2ed44f} /* (14, 8, 6) {real, imag} */,
  {32'hc086cd8e, 32'hbf94e677} /* (14, 8, 5) {real, imag} */,
  {32'hc073dd27, 32'hc07b31a8} /* (14, 8, 4) {real, imag} */,
  {32'hc093aea1, 32'h3fc49fdc} /* (14, 8, 3) {real, imag} */,
  {32'hc0bc83c4, 32'hc0b34c7c} /* (14, 8, 2) {real, imag} */,
  {32'hc03fc1fc, 32'h3f4b5b57} /* (14, 8, 1) {real, imag} */,
  {32'h3e293d05, 32'hc0821a1a} /* (14, 8, 0) {real, imag} */,
  {32'hc03b6914, 32'h3e82e22c} /* (14, 7, 15) {real, imag} */,
  {32'hbf72932a, 32'hc06ca6a1} /* (14, 7, 14) {real, imag} */,
  {32'h40ea6a50, 32'hbfe42b44} /* (14, 7, 13) {real, imag} */,
  {32'hc0d50817, 32'hbf9875f3} /* (14, 7, 12) {real, imag} */,
  {32'hc0fc0bb5, 32'h3e01af94} /* (14, 7, 11) {real, imag} */,
  {32'hc0b036fc, 32'hbf5f7700} /* (14, 7, 10) {real, imag} */,
  {32'hbfc52e81, 32'h3f465da7} /* (14, 7, 9) {real, imag} */,
  {32'h40987881, 32'h4039a288} /* (14, 7, 8) {real, imag} */,
  {32'h3e6d8c8b, 32'h3ea54dfe} /* (14, 7, 7) {real, imag} */,
  {32'hc0c4d6e1, 32'h404242d0} /* (14, 7, 6) {real, imag} */,
  {32'h3f24acec, 32'h40d7227c} /* (14, 7, 5) {real, imag} */,
  {32'h40533f1b, 32'h4090d775} /* (14, 7, 4) {real, imag} */,
  {32'h3f308496, 32'h40941ead} /* (14, 7, 3) {real, imag} */,
  {32'hbd243917, 32'h4015f72b} /* (14, 7, 2) {real, imag} */,
  {32'hc0192c87, 32'h3ea5b609} /* (14, 7, 1) {real, imag} */,
  {32'h40140570, 32'h3ff8d9c3} /* (14, 7, 0) {real, imag} */,
  {32'h4098ea72, 32'hbec30641} /* (14, 6, 15) {real, imag} */,
  {32'hc01897f7, 32'h3eb7610b} /* (14, 6, 14) {real, imag} */,
  {32'h40cb5ad6, 32'hc00b27a9} /* (14, 6, 13) {real, imag} */,
  {32'hc0adcf76, 32'h40ac93f9} /* (14, 6, 12) {real, imag} */,
  {32'h408b9dda, 32'hc03e00be} /* (14, 6, 11) {real, imag} */,
  {32'h40868d5a, 32'hbf5959ba} /* (14, 6, 10) {real, imag} */,
  {32'hbfaeeb97, 32'h407b192e} /* (14, 6, 9) {real, imag} */,
  {32'hc01f7e74, 32'h40183c3a} /* (14, 6, 8) {real, imag} */,
  {32'hc03b87d8, 32'h3fc0a318} /* (14, 6, 7) {real, imag} */,
  {32'hc08a9599, 32'hbe9e162d} /* (14, 6, 6) {real, imag} */,
  {32'hbfa816d0, 32'h3ff53f7e} /* (14, 6, 5) {real, imag} */,
  {32'h3fc1d7d2, 32'hc0ff572c} /* (14, 6, 4) {real, imag} */,
  {32'hc069a39b, 32'h3f178c19} /* (14, 6, 3) {real, imag} */,
  {32'hc0f7fdd4, 32'h3fabab6b} /* (14, 6, 2) {real, imag} */,
  {32'hc01b54d5, 32'hc0683223} /* (14, 6, 1) {real, imag} */,
  {32'h4084b32d, 32'hbffc07d8} /* (14, 6, 0) {real, imag} */,
  {32'hbefc3636, 32'h40360225} /* (14, 5, 15) {real, imag} */,
  {32'hc0f90562, 32'hc047fa30} /* (14, 5, 14) {real, imag} */,
  {32'hbf7b7280, 32'h406c52d2} /* (14, 5, 13) {real, imag} */,
  {32'h40ae469b, 32'h4042a6e7} /* (14, 5, 12) {real, imag} */,
  {32'hc038acfe, 32'hbf8a6a84} /* (14, 5, 11) {real, imag} */,
  {32'h40e7d599, 32'hbfb47b4a} /* (14, 5, 10) {real, imag} */,
  {32'h40bc9882, 32'hc0eee966} /* (14, 5, 9) {real, imag} */,
  {32'h3e82620a, 32'h40147c60} /* (14, 5, 8) {real, imag} */,
  {32'h4069025e, 32'h409f1a35} /* (14, 5, 7) {real, imag} */,
  {32'h40ce4e3f, 32'hc0f7ee37} /* (14, 5, 6) {real, imag} */,
  {32'hc059bf02, 32'hc095db76} /* (14, 5, 5) {real, imag} */,
  {32'hc081dd4d, 32'h405de783} /* (14, 5, 4) {real, imag} */,
  {32'hbf8f2576, 32'hc09085f3} /* (14, 5, 3) {real, imag} */,
  {32'h3fd8f2ec, 32'h40cfafcc} /* (14, 5, 2) {real, imag} */,
  {32'h41097fba, 32'h413cc050} /* (14, 5, 1) {real, imag} */,
  {32'h4063fc9b, 32'hc0f3f917} /* (14, 5, 0) {real, imag} */,
  {32'h4097d034, 32'h415ddda8} /* (14, 4, 15) {real, imag} */,
  {32'hbf446ceb, 32'h404bc527} /* (14, 4, 14) {real, imag} */,
  {32'h40923a15, 32'h40d27e62} /* (14, 4, 13) {real, imag} */,
  {32'h410cd4e7, 32'hc1742529} /* (14, 4, 12) {real, imag} */,
  {32'hbf164d62, 32'h41210048} /* (14, 4, 11) {real, imag} */,
  {32'h4065aeaf, 32'h404734a9} /* (14, 4, 10) {real, imag} */,
  {32'h40824ca3, 32'h40a2cdb0} /* (14, 4, 9) {real, imag} */,
  {32'hc0ad7333, 32'hbfd02556} /* (14, 4, 8) {real, imag} */,
  {32'h3f324b8f, 32'hbfe87114} /* (14, 4, 7) {real, imag} */,
  {32'hc0520f5c, 32'hbfdc15d9} /* (14, 4, 6) {real, imag} */,
  {32'h4187b5f5, 32'h40978c8b} /* (14, 4, 5) {real, imag} */,
  {32'hbf086fdb, 32'h3fb4033d} /* (14, 4, 4) {real, imag} */,
  {32'h3fce97af, 32'hc1af75bc} /* (14, 4, 3) {real, imag} */,
  {32'hc023ce29, 32'h407a3f90} /* (14, 4, 2) {real, imag} */,
  {32'hbf8469e9, 32'hbfc0d386} /* (14, 4, 1) {real, imag} */,
  {32'h3ff4fb9c, 32'hc059948d} /* (14, 4, 0) {real, imag} */,
  {32'h40a463b1, 32'hc15c557f} /* (14, 3, 15) {real, imag} */,
  {32'h3f96623c, 32'hc095dc9e} /* (14, 3, 14) {real, imag} */,
  {32'h3ee7df85, 32'h409a2027} /* (14, 3, 13) {real, imag} */,
  {32'h3f84c106, 32'hc1372222} /* (14, 3, 12) {real, imag} */,
  {32'h40af1ba5, 32'h40ab52f6} /* (14, 3, 11) {real, imag} */,
  {32'h403fc84a, 32'h40bf8cc6} /* (14, 3, 10) {real, imag} */,
  {32'h4039f606, 32'hc0a44caf} /* (14, 3, 9) {real, imag} */,
  {32'hc00c117e, 32'hbf45db82} /* (14, 3, 8) {real, imag} */,
  {32'hc0c0ea1b, 32'hbff3751b} /* (14, 3, 7) {real, imag} */,
  {32'hc02bb1a3, 32'hc0008202} /* (14, 3, 6) {real, imag} */,
  {32'hc09f1e13, 32'h3ebed3f1} /* (14, 3, 5) {real, imag} */,
  {32'h4158f9a1, 32'hc053dfb6} /* (14, 3, 4) {real, imag} */,
  {32'h41411bf8, 32'hc0053ae8} /* (14, 3, 3) {real, imag} */,
  {32'h3fce6a09, 32'hbfbbdd37} /* (14, 3, 2) {real, imag} */,
  {32'hc09d956e, 32'h3d9db9ac} /* (14, 3, 1) {real, imag} */,
  {32'hc007c99a, 32'h4002f782} /* (14, 3, 0) {real, imag} */,
  {32'h418be2e3, 32'h41d1baeb} /* (14, 2, 15) {real, imag} */,
  {32'h416fe832, 32'h410e11a0} /* (14, 2, 14) {real, imag} */,
  {32'h3fe8c321, 32'h41257ee3} /* (14, 2, 13) {real, imag} */,
  {32'hbf942ca6, 32'hc11874ce} /* (14, 2, 12) {real, imag} */,
  {32'hbff0f5e5, 32'hc00585de} /* (14, 2, 11) {real, imag} */,
  {32'h3dc9f830, 32'hbf7b5986} /* (14, 2, 10) {real, imag} */,
  {32'hbf99f8bf, 32'h3fbb4d32} /* (14, 2, 9) {real, imag} */,
  {32'h3d42c9a2, 32'h3ec3d88c} /* (14, 2, 8) {real, imag} */,
  {32'hbf15797c, 32'hc01ed5dd} /* (14, 2, 7) {real, imag} */,
  {32'h3f83cf4d, 32'hc014e5c4} /* (14, 2, 6) {real, imag} */,
  {32'h40914d03, 32'hc049dc03} /* (14, 2, 5) {real, imag} */,
  {32'hbfe57f63, 32'h409ce21d} /* (14, 2, 4) {real, imag} */,
  {32'h41992c98, 32'hc051db31} /* (14, 2, 3) {real, imag} */,
  {32'h3fd81f60, 32'hc136b930} /* (14, 2, 2) {real, imag} */,
  {32'hc235186c, 32'hc08e37ab} /* (14, 2, 1) {real, imag} */,
  {32'hc0d2f493, 32'h4082ff3c} /* (14, 2, 0) {real, imag} */,
  {32'hc14e7e58, 32'hc11be58a} /* (14, 1, 15) {real, imag} */,
  {32'hc08dbc97, 32'h4103dc3f} /* (14, 1, 14) {real, imag} */,
  {32'hbc852c80, 32'h40b6397f} /* (14, 1, 13) {real, imag} */,
  {32'h3f99241a, 32'hc19dc948} /* (14, 1, 12) {real, imag} */,
  {32'hbf74c4a1, 32'hbfe00257} /* (14, 1, 11) {real, imag} */,
  {32'h3ef349d2, 32'h405816c7} /* (14, 1, 10) {real, imag} */,
  {32'hc015ac1d, 32'hc0b3f5cf} /* (14, 1, 9) {real, imag} */,
  {32'hbfb0acd3, 32'hbee18cbc} /* (14, 1, 8) {real, imag} */,
  {32'hbaae89b8, 32'hc0787b64} /* (14, 1, 7) {real, imag} */,
  {32'hbfbc9772, 32'hbe0be238} /* (14, 1, 6) {real, imag} */,
  {32'hbf3ca61f, 32'hbf2c5a03} /* (14, 1, 5) {real, imag} */,
  {32'hc0a43f19, 32'hbf8281cc} /* (14, 1, 4) {real, imag} */,
  {32'h409c195e, 32'h41063807} /* (14, 1, 3) {real, imag} */,
  {32'h41d59e36, 32'h3fb8114f} /* (14, 1, 2) {real, imag} */,
  {32'h3dd853e8, 32'hc19ff426} /* (14, 1, 1) {real, imag} */,
  {32'hc22204cb, 32'h408b92c8} /* (14, 1, 0) {real, imag} */,
  {32'h415e4540, 32'hc0a94fff} /* (14, 0, 15) {real, imag} */,
  {32'hbe9ffd8a, 32'hbd348ce6} /* (14, 0, 14) {real, imag} */,
  {32'hc1241861, 32'h4097f0ae} /* (14, 0, 13) {real, imag} */,
  {32'hbf2b74a2, 32'h415ca590} /* (14, 0, 12) {real, imag} */,
  {32'hc14951d7, 32'h3f72251f} /* (14, 0, 11) {real, imag} */,
  {32'hbfdbc11b, 32'h3f1685b0} /* (14, 0, 10) {real, imag} */,
  {32'h3d43bced, 32'h3f32687b} /* (14, 0, 9) {real, imag} */,
  {32'h40c816bf, 32'hc0285e06} /* (14, 0, 8) {real, imag} */,
  {32'hbf6dd62f, 32'h40816368} /* (14, 0, 7) {real, imag} */,
  {32'hbfcc3abe, 32'hc101a282} /* (14, 0, 6) {real, imag} */,
  {32'h40d044b4, 32'h401c8ebf} /* (14, 0, 5) {real, imag} */,
  {32'hc0af23fd, 32'h3fba7dfa} /* (14, 0, 4) {real, imag} */,
  {32'h41641223, 32'h4072da92} /* (14, 0, 3) {real, imag} */,
  {32'hc1165c31, 32'hc03c94c7} /* (14, 0, 2) {real, imag} */,
  {32'h4096977f, 32'h40ed4fe7} /* (14, 0, 1) {real, imag} */,
  {32'h41e91fb8, 32'h4281efb1} /* (14, 0, 0) {real, imag} */,
  {32'hc168b51b, 32'hc1350bdf} /* (13, 15, 15) {real, imag} */,
  {32'h40ce0335, 32'h408fc691} /* (13, 15, 14) {real, imag} */,
  {32'h41567895, 32'hc11ad06b} /* (13, 15, 13) {real, imag} */,
  {32'hbfec2936, 32'hbfd0dcd2} /* (13, 15, 12) {real, imag} */,
  {32'h3f469aef, 32'hc00e0e90} /* (13, 15, 11) {real, imag} */,
  {32'h409d18b5, 32'h411fd03f} /* (13, 15, 10) {real, imag} */,
  {32'h3ee0d7d7, 32'h3fc1168f} /* (13, 15, 9) {real, imag} */,
  {32'hbf41b865, 32'hc038e5ba} /* (13, 15, 8) {real, imag} */,
  {32'hc10ee7db, 32'h3fc2bca1} /* (13, 15, 7) {real, imag} */,
  {32'hbfdceed1, 32'hc051424e} /* (13, 15, 6) {real, imag} */,
  {32'hc0370230, 32'hbf9bf946} /* (13, 15, 5) {real, imag} */,
  {32'h4039dea8, 32'h3ce733c4} /* (13, 15, 4) {real, imag} */,
  {32'hc0bd0339, 32'h40e51bd2} /* (13, 15, 3) {real, imag} */,
  {32'hc176b20b, 32'h407d95bb} /* (13, 15, 2) {real, imag} */,
  {32'h40cbfdf3, 32'h40d4d676} /* (13, 15, 1) {real, imag} */,
  {32'hc10b97b3, 32'hc15deff9} /* (13, 15, 0) {real, imag} */,
  {32'hc0be9944, 32'hbda352c8} /* (13, 14, 15) {real, imag} */,
  {32'h41268ded, 32'h4132ba34} /* (13, 14, 14) {real, imag} */,
  {32'hc043824e, 32'h404320b1} /* (13, 14, 13) {real, imag} */,
  {32'h40fb43d7, 32'hbff96528} /* (13, 14, 12) {real, imag} */,
  {32'h40c7b596, 32'h3faf841a} /* (13, 14, 11) {real, imag} */,
  {32'hc023c7e0, 32'hbfa7411a} /* (13, 14, 10) {real, imag} */,
  {32'h3f2429d1, 32'hbead63eb} /* (13, 14, 9) {real, imag} */,
  {32'h3fc0a641, 32'hbfc4c810} /* (13, 14, 8) {real, imag} */,
  {32'h3f08bd30, 32'h3ef8f386} /* (13, 14, 7) {real, imag} */,
  {32'h3fd19c46, 32'hc00b1517} /* (13, 14, 6) {real, imag} */,
  {32'hc03852b5, 32'hc12b6247} /* (13, 14, 5) {real, imag} */,
  {32'h40c72054, 32'h3e167928} /* (13, 14, 4) {real, imag} */,
  {32'h4081740b, 32'h41395947} /* (13, 14, 3) {real, imag} */,
  {32'h416502a6, 32'hc145e652} /* (13, 14, 2) {real, imag} */,
  {32'h41196145, 32'hc195dca1} /* (13, 14, 1) {real, imag} */,
  {32'hc1321b7a, 32'h4068041f} /* (13, 14, 0) {real, imag} */,
  {32'hc0e6a322, 32'h40bbcf5c} /* (13, 13, 15) {real, imag} */,
  {32'h3de1edf4, 32'hc112a104} /* (13, 13, 14) {real, imag} */,
  {32'hc09b6d32, 32'h401b422c} /* (13, 13, 13) {real, imag} */,
  {32'h3fc03f17, 32'h4104bbf6} /* (13, 13, 12) {real, imag} */,
  {32'hc14bc7cd, 32'hc04d2dbd} /* (13, 13, 11) {real, imag} */,
  {32'hbeb28a1b, 32'h412abf9e} /* (13, 13, 10) {real, imag} */,
  {32'hc0bea61c, 32'h40b51a63} /* (13, 13, 9) {real, imag} */,
  {32'h408ff864, 32'hbe75af3c} /* (13, 13, 8) {real, imag} */,
  {32'hbf1ab9a9, 32'hbfacfb63} /* (13, 13, 7) {real, imag} */,
  {32'hc0b21d97, 32'h404c0830} /* (13, 13, 6) {real, imag} */,
  {32'h407270da, 32'h4106dcfc} /* (13, 13, 5) {real, imag} */,
  {32'hbf15a8d7, 32'h40d0dc40} /* (13, 13, 4) {real, imag} */,
  {32'h40a5e74a, 32'hbe7db0fb} /* (13, 13, 3) {real, imag} */,
  {32'h408e5a08, 32'h41203f02} /* (13, 13, 2) {real, imag} */,
  {32'h3f44a88f, 32'h3f372a1f} /* (13, 13, 1) {real, imag} */,
  {32'h40e2426b, 32'hc07ebd59} /* (13, 13, 0) {real, imag} */,
  {32'h4186a8d5, 32'hc11937c2} /* (13, 12, 15) {real, imag} */,
  {32'h3d873785, 32'h40962575} /* (13, 12, 14) {real, imag} */,
  {32'hc0082f29, 32'hc00f72bf} /* (13, 12, 13) {real, imag} */,
  {32'hc0e55523, 32'hc00d2ef8} /* (13, 12, 12) {real, imag} */,
  {32'hc0cd594e, 32'h3f643428} /* (13, 12, 11) {real, imag} */,
  {32'h411427b1, 32'hbfeb3138} /* (13, 12, 10) {real, imag} */,
  {32'hbfa56c8f, 32'h409fd571} /* (13, 12, 9) {real, imag} */,
  {32'h402d0dc5, 32'hbfbbf4df} /* (13, 12, 8) {real, imag} */,
  {32'hbf6eb275, 32'h3fab3e2c} /* (13, 12, 7) {real, imag} */,
  {32'h3fb863f3, 32'h3f8f4fd4} /* (13, 12, 6) {real, imag} */,
  {32'hbe8d501a, 32'hc07d6b39} /* (13, 12, 5) {real, imag} */,
  {32'hbe43cb71, 32'h417af258} /* (13, 12, 4) {real, imag} */,
  {32'hbfe5a5aa, 32'hc1152ce6} /* (13, 12, 3) {real, imag} */,
  {32'h41172118, 32'hc090676f} /* (13, 12, 2) {real, imag} */,
  {32'h405c37b6, 32'h3e83de9f} /* (13, 12, 1) {real, imag} */,
  {32'hc10fc4eb, 32'h40eb8788} /* (13, 12, 0) {real, imag} */,
  {32'h3ff0f7f6, 32'hc087000e} /* (13, 11, 15) {real, imag} */,
  {32'hbfd52d96, 32'hc03d0219} /* (13, 11, 14) {real, imag} */,
  {32'hc00137fe, 32'h40124cb9} /* (13, 11, 13) {real, imag} */,
  {32'hc17d29da, 32'hc131803f} /* (13, 11, 12) {real, imag} */,
  {32'hc017407c, 32'h4009664c} /* (13, 11, 11) {real, imag} */,
  {32'h401ab879, 32'hc092439e} /* (13, 11, 10) {real, imag} */,
  {32'hc0538a82, 32'hbeb2a171} /* (13, 11, 9) {real, imag} */,
  {32'h3f2d7f8a, 32'h40089a23} /* (13, 11, 8) {real, imag} */,
  {32'h40c7355e, 32'hc01fb972} /* (13, 11, 7) {real, imag} */,
  {32'hc0878cf5, 32'hc0c0586b} /* (13, 11, 6) {real, imag} */,
  {32'hbdfba962, 32'hc121dc85} /* (13, 11, 5) {real, imag} */,
  {32'hbef0b576, 32'hbffb9a33} /* (13, 11, 4) {real, imag} */,
  {32'hc0cf045e, 32'h416e4f75} /* (13, 11, 3) {real, imag} */,
  {32'h3f95ae03, 32'hbfc9fcc5} /* (13, 11, 2) {real, imag} */,
  {32'h40ed12f0, 32'h40d5f56b} /* (13, 11, 1) {real, imag} */,
  {32'hbf83407c, 32'h4146487f} /* (13, 11, 0) {real, imag} */,
  {32'h3fe620fe, 32'hc0ba14f1} /* (13, 10, 15) {real, imag} */,
  {32'h401a0df5, 32'h40297e31} /* (13, 10, 14) {real, imag} */,
  {32'h3f594405, 32'h3df56372} /* (13, 10, 13) {real, imag} */,
  {32'hc0c25638, 32'hc1186162} /* (13, 10, 12) {real, imag} */,
  {32'h40a6abc0, 32'h3ea68ae0} /* (13, 10, 11) {real, imag} */,
  {32'h3f378b44, 32'h3f99c232} /* (13, 10, 10) {real, imag} */,
  {32'h40cd4e91, 32'hc018f79a} /* (13, 10, 9) {real, imag} */,
  {32'hc012398a, 32'h409c753f} /* (13, 10, 8) {real, imag} */,
  {32'hc009f839, 32'hc06b4d32} /* (13, 10, 7) {real, imag} */,
  {32'h3f397839, 32'hc06dda49} /* (13, 10, 6) {real, imag} */,
  {32'h40c2cadb, 32'h40d30ae8} /* (13, 10, 5) {real, imag} */,
  {32'hbf1bda83, 32'h403ece04} /* (13, 10, 4) {real, imag} */,
  {32'hbed95429, 32'h3f88606e} /* (13, 10, 3) {real, imag} */,
  {32'h3ed074c2, 32'h3fa81e5d} /* (13, 10, 2) {real, imag} */,
  {32'hc106e226, 32'h40bad9eb} /* (13, 10, 1) {real, imag} */,
  {32'hc102a751, 32'h3eef19d4} /* (13, 10, 0) {real, imag} */,
  {32'hc0a13a6b, 32'h403440de} /* (13, 9, 15) {real, imag} */,
  {32'h3e832974, 32'hbfbb4492} /* (13, 9, 14) {real, imag} */,
  {32'h40395c9b, 32'h40e47c83} /* (13, 9, 13) {real, imag} */,
  {32'h405a2646, 32'h402244e6} /* (13, 9, 12) {real, imag} */,
  {32'hbff339d1, 32'hbffddd0a} /* (13, 9, 11) {real, imag} */,
  {32'hc095e7fe, 32'h402efae2} /* (13, 9, 10) {real, imag} */,
  {32'h40d7700a, 32'hc0292b14} /* (13, 9, 9) {real, imag} */,
  {32'hc0bc2cfb, 32'hbe646c6e} /* (13, 9, 8) {real, imag} */,
  {32'hbf15def7, 32'hc0140267} /* (13, 9, 7) {real, imag} */,
  {32'h409280fc, 32'hbf02879f} /* (13, 9, 6) {real, imag} */,
  {32'hbf2244a5, 32'h3f29c9c1} /* (13, 9, 5) {real, imag} */,
  {32'hbffa67f3, 32'h3dc68f36} /* (13, 9, 4) {real, imag} */,
  {32'h407729fe, 32'hc06c9928} /* (13, 9, 3) {real, imag} */,
  {32'h410248c1, 32'hbfe5b85a} /* (13, 9, 2) {real, imag} */,
  {32'hbf923c8f, 32'h4097a4c2} /* (13, 9, 1) {real, imag} */,
  {32'h3d2f77b8, 32'hbec03d59} /* (13, 9, 0) {real, imag} */,
  {32'hbfdc52a0, 32'h3fc9fd44} /* (13, 8, 15) {real, imag} */,
  {32'hbf9c24f7, 32'h404f9548} /* (13, 8, 14) {real, imag} */,
  {32'h40211c30, 32'hc0b44a42} /* (13, 8, 13) {real, imag} */,
  {32'h408ce177, 32'hc01837d0} /* (13, 8, 12) {real, imag} */,
  {32'h3ffa0eb6, 32'h3f3bfd0c} /* (13, 8, 11) {real, imag} */,
  {32'hc0394820, 32'hbf34e83c} /* (13, 8, 10) {real, imag} */,
  {32'h401dd922, 32'hbf0f4c43} /* (13, 8, 9) {real, imag} */,
  {32'hc065abe1, 32'h3e9dd167} /* (13, 8, 8) {real, imag} */,
  {32'h40d0e74e, 32'h4112cb63} /* (13, 8, 7) {real, imag} */,
  {32'h4063fd5c, 32'h40764f28} /* (13, 8, 6) {real, imag} */,
  {32'hc0d5e0c2, 32'h407d7bbc} /* (13, 8, 5) {real, imag} */,
  {32'h3fa6788e, 32'hbeb0d96f} /* (13, 8, 4) {real, imag} */,
  {32'hbf13f980, 32'hc0077ef2} /* (13, 8, 3) {real, imag} */,
  {32'hbf6ad8b4, 32'hbea3daf3} /* (13, 8, 2) {real, imag} */,
  {32'h40204646, 32'hc02f0a2a} /* (13, 8, 1) {real, imag} */,
  {32'h3f263e4e, 32'h3fd33e7e} /* (13, 8, 0) {real, imag} */,
  {32'h40013783, 32'h40421f63} /* (13, 7, 15) {real, imag} */,
  {32'hc07f5764, 32'h406b6262} /* (13, 7, 14) {real, imag} */,
  {32'hc05c660c, 32'h40d6150c} /* (13, 7, 13) {real, imag} */,
  {32'hbfa95b6e, 32'hc09128dc} /* (13, 7, 12) {real, imag} */,
  {32'h40f9caf8, 32'hc048366e} /* (13, 7, 11) {real, imag} */,
  {32'h3f85a97c, 32'hc10597a8} /* (13, 7, 10) {real, imag} */,
  {32'hbf25f186, 32'hc095a269} /* (13, 7, 9) {real, imag} */,
  {32'hbfbc8ce5, 32'hc03f027e} /* (13, 7, 8) {real, imag} */,
  {32'hbf02f407, 32'h40ddfe11} /* (13, 7, 7) {real, imag} */,
  {32'h402752a7, 32'hc04cc238} /* (13, 7, 6) {real, imag} */,
  {32'hbfef949a, 32'h402dd992} /* (13, 7, 5) {real, imag} */,
  {32'hbf914ba5, 32'h407d706e} /* (13, 7, 4) {real, imag} */,
  {32'h409e535c, 32'hbe003e7c} /* (13, 7, 3) {real, imag} */,
  {32'h40635030, 32'hc03f0e12} /* (13, 7, 2) {real, imag} */,
  {32'h3fa99d43, 32'hc09f6b97} /* (13, 7, 1) {real, imag} */,
  {32'hc08cf8dd, 32'h3f407e88} /* (13, 7, 0) {real, imag} */,
  {32'hbff1ec04, 32'hc099db5c} /* (13, 6, 15) {real, imag} */,
  {32'h405dfe67, 32'hc0e8a374} /* (13, 6, 14) {real, imag} */,
  {32'h3eb243f7, 32'hc11472fc} /* (13, 6, 13) {real, imag} */,
  {32'hbff9a097, 32'h4008c207} /* (13, 6, 12) {real, imag} */,
  {32'hc090cb8d, 32'hc0caf30e} /* (13, 6, 11) {real, imag} */,
  {32'h40b480d5, 32'h3fb2dde8} /* (13, 6, 10) {real, imag} */,
  {32'h3f1a4b39, 32'h4117e1ce} /* (13, 6, 9) {real, imag} */,
  {32'hbff35e8b, 32'h3f4dd9f7} /* (13, 6, 8) {real, imag} */,
  {32'h402994b7, 32'h3ed31afd} /* (13, 6, 7) {real, imag} */,
  {32'hc0769945, 32'h410428b4} /* (13, 6, 6) {real, imag} */,
  {32'hc014e170, 32'hc08c07cd} /* (13, 6, 5) {real, imag} */,
  {32'hc0c34141, 32'h407aa1b3} /* (13, 6, 4) {real, imag} */,
  {32'hbfdf99e1, 32'hc11e7909} /* (13, 6, 3) {real, imag} */,
  {32'h3e7570bc, 32'h40892b7b} /* (13, 6, 2) {real, imag} */,
  {32'hc053ea6a, 32'h406dc09b} /* (13, 6, 1) {real, imag} */,
  {32'h3e3b1d3a, 32'hc0156d47} /* (13, 6, 0) {real, imag} */,
  {32'h411d40f9, 32'hc10689b8} /* (13, 5, 15) {real, imag} */,
  {32'h3daf42b8, 32'hc091b8cd} /* (13, 5, 14) {real, imag} */,
  {32'hc0dac0eb, 32'h40013127} /* (13, 5, 13) {real, imag} */,
  {32'hc08a431a, 32'h3e80e5aa} /* (13, 5, 12) {real, imag} */,
  {32'h40102f8c, 32'h4108f8d9} /* (13, 5, 11) {real, imag} */,
  {32'h40f77f0d, 32'h408529c1} /* (13, 5, 10) {real, imag} */,
  {32'h40c50664, 32'h409e092b} /* (13, 5, 9) {real, imag} */,
  {32'h3de34415, 32'h3f95eaea} /* (13, 5, 8) {real, imag} */,
  {32'hc0fa7d30, 32'hc0b36edb} /* (13, 5, 7) {real, imag} */,
  {32'h3f027575, 32'h40f549ae} /* (13, 5, 6) {real, imag} */,
  {32'hbfefc6da, 32'hc0758d08} /* (13, 5, 5) {real, imag} */,
  {32'hc0cf7c72, 32'h409fcaa3} /* (13, 5, 4) {real, imag} */,
  {32'hbec8c493, 32'hbeebdef8} /* (13, 5, 3) {real, imag} */,
  {32'h413c9d40, 32'hc0529213} /* (13, 5, 2) {real, imag} */,
  {32'hc0ad6570, 32'hc0d160cd} /* (13, 5, 1) {real, imag} */,
  {32'hc0a20fdc, 32'hbf465326} /* (13, 5, 0) {real, imag} */,
  {32'h401e4f54, 32'h41709db4} /* (13, 4, 15) {real, imag} */,
  {32'h402c0509, 32'hbf9c6fba} /* (13, 4, 14) {real, imag} */,
  {32'h4123ce63, 32'hbfb536d0} /* (13, 4, 13) {real, imag} */,
  {32'hc127348c, 32'h3e4f7ad2} /* (13, 4, 12) {real, imag} */,
  {32'h3dcb041b, 32'hc0c0d862} /* (13, 4, 11) {real, imag} */,
  {32'hc125cb36, 32'hc0d7ae6c} /* (13, 4, 10) {real, imag} */,
  {32'hbf946963, 32'hbf4cd93b} /* (13, 4, 9) {real, imag} */,
  {32'hbee19fd7, 32'h408b1196} /* (13, 4, 8) {real, imag} */,
  {32'h4107ecf5, 32'h3fd9e0c0} /* (13, 4, 7) {real, imag} */,
  {32'hc0e600fd, 32'hc046430d} /* (13, 4, 6) {real, imag} */,
  {32'hc0e32e40, 32'h411f6120} /* (13, 4, 5) {real, imag} */,
  {32'hbec3b00d, 32'hbf93e289} /* (13, 4, 4) {real, imag} */,
  {32'h40c5fe03, 32'h40a276a8} /* (13, 4, 3) {real, imag} */,
  {32'hbf1b5009, 32'hc0521288} /* (13, 4, 2) {real, imag} */,
  {32'h40e1b520, 32'hbf7f6a88} /* (13, 4, 1) {real, imag} */,
  {32'hc005b869, 32'hbfa77930} /* (13, 4, 0) {real, imag} */,
  {32'h40cabf61, 32'h3fb94b3f} /* (13, 3, 15) {real, imag} */,
  {32'hc10e7ea2, 32'h401e27f7} /* (13, 3, 14) {real, imag} */,
  {32'h40046fcd, 32'h4102b5d9} /* (13, 3, 13) {real, imag} */,
  {32'hbe3dd80c, 32'hc01bebac} /* (13, 3, 12) {real, imag} */,
  {32'h40b0071a, 32'hc019c010} /* (13, 3, 11) {real, imag} */,
  {32'h4112cf9d, 32'hc0b4cde1} /* (13, 3, 10) {real, imag} */,
  {32'h3ff176f6, 32'h3fab3c40} /* (13, 3, 9) {real, imag} */,
  {32'h410305d8, 32'h3f27347a} /* (13, 3, 8) {real, imag} */,
  {32'h403034c4, 32'hc01e185c} /* (13, 3, 7) {real, imag} */,
  {32'h3fdb58b4, 32'hc00bef70} /* (13, 3, 6) {real, imag} */,
  {32'hc094859f, 32'h4093d643} /* (13, 3, 5) {real, imag} */,
  {32'h4183b1f9, 32'h40b77d9d} /* (13, 3, 4) {real, imag} */,
  {32'h41170ee1, 32'hc0b06c79} /* (13, 3, 3) {real, imag} */,
  {32'hc0865bea, 32'h40f0bbfe} /* (13, 3, 2) {real, imag} */,
  {32'hc0a68d4a, 32'hc093d175} /* (13, 3, 1) {real, imag} */,
  {32'hc0fa605a, 32'hbe373c99} /* (13, 3, 0) {real, imag} */,
  {32'hc064695f, 32'h3f36361d} /* (13, 2, 15) {real, imag} */,
  {32'hc08f4a3f, 32'h3f11eb9a} /* (13, 2, 14) {real, imag} */,
  {32'h3e4f19d7, 32'hc0976fa3} /* (13, 2, 13) {real, imag} */,
  {32'h40983997, 32'hbeb2b301} /* (13, 2, 12) {real, imag} */,
  {32'h409b8671, 32'hbfe1774b} /* (13, 2, 11) {real, imag} */,
  {32'hc12cee8a, 32'hc0098fa1} /* (13, 2, 10) {real, imag} */,
  {32'hc0ce2ce8, 32'h40ba90a8} /* (13, 2, 9) {real, imag} */,
  {32'hc01a9e68, 32'h408247a5} /* (13, 2, 8) {real, imag} */,
  {32'h3d33c78e, 32'hbfee92a3} /* (13, 2, 7) {real, imag} */,
  {32'hc03dc734, 32'h3e7efe97} /* (13, 2, 6) {real, imag} */,
  {32'h3f3d068d, 32'h401b332f} /* (13, 2, 5) {real, imag} */,
  {32'hbccfd9ff, 32'hc0d23980} /* (13, 2, 4) {real, imag} */,
  {32'h3f90bf40, 32'h411ee0ec} /* (13, 2, 3) {real, imag} */,
  {32'hc108b1c8, 32'h406b6835} /* (13, 2, 2) {real, imag} */,
  {32'h4067553f, 32'h41153fef} /* (13, 2, 1) {real, imag} */,
  {32'h410565ac, 32'hc01870c9} /* (13, 2, 0) {real, imag} */,
  {32'hc18f4955, 32'h4106844e} /* (13, 1, 15) {real, imag} */,
  {32'hc01a3ac1, 32'hc0be817f} /* (13, 1, 14) {real, imag} */,
  {32'hc0a23499, 32'h40ed8f71} /* (13, 1, 13) {real, imag} */,
  {32'h40cadd20, 32'hbd38b123} /* (13, 1, 12) {real, imag} */,
  {32'h40babda3, 32'h415b25a8} /* (13, 1, 11) {real, imag} */,
  {32'hc00dfe53, 32'hc0dec1cd} /* (13, 1, 10) {real, imag} */,
  {32'hc048a66d, 32'hc0244f47} /* (13, 1, 9) {real, imag} */,
  {32'hc01fdfc3, 32'hbfcb49dc} /* (13, 1, 8) {real, imag} */,
  {32'h3f5478f5, 32'h4016478f} /* (13, 1, 7) {real, imag} */,
  {32'h41109528, 32'hc0b7f3bf} /* (13, 1, 6) {real, imag} */,
  {32'h40b92e08, 32'hc13e5efe} /* (13, 1, 5) {real, imag} */,
  {32'h3f6ee909, 32'hc1374b37} /* (13, 1, 4) {real, imag} */,
  {32'h40a47e77, 32'hc0c4b74e} /* (13, 1, 3) {real, imag} */,
  {32'hc18512af, 32'h40dc2428} /* (13, 1, 2) {real, imag} */,
  {32'h3fcebb0e, 32'hbf5b732f} /* (13, 1, 1) {real, imag} */,
  {32'h40afa5cd, 32'h40568109} /* (13, 1, 0) {real, imag} */,
  {32'h40ef830a, 32'h41483ce9} /* (13, 0, 15) {real, imag} */,
  {32'h3f64746d, 32'hbfe660f7} /* (13, 0, 14) {real, imag} */,
  {32'hc021cf7b, 32'hc109dd2c} /* (13, 0, 13) {real, imag} */,
  {32'hc000b965, 32'hc0815f00} /* (13, 0, 12) {real, imag} */,
  {32'hbf873a03, 32'h418b2a03} /* (13, 0, 11) {real, imag} */,
  {32'hc0435496, 32'hc045e56f} /* (13, 0, 10) {real, imag} */,
  {32'h40f5adba, 32'hbc78ef12} /* (13, 0, 9) {real, imag} */,
  {32'hbfce924b, 32'hc0a3e63e} /* (13, 0, 8) {real, imag} */,
  {32'h3fb46335, 32'h3fe8d137} /* (13, 0, 7) {real, imag} */,
  {32'hbedd6488, 32'hbe899dc5} /* (13, 0, 6) {real, imag} */,
  {32'h3faf6c44, 32'hc148daa6} /* (13, 0, 5) {real, imag} */,
  {32'hc164d78d, 32'h4132f946} /* (13, 0, 4) {real, imag} */,
  {32'h40be77de, 32'h4029f4ef} /* (13, 0, 3) {real, imag} */,
  {32'h4188093d, 32'hc0dcd2c6} /* (13, 0, 2) {real, imag} */,
  {32'hbf9f9ed1, 32'hc19d68de} /* (13, 0, 1) {real, imag} */,
  {32'h4123be88, 32'h41a2eb87} /* (13, 0, 0) {real, imag} */,
  {32'hc0e932b1, 32'hc0aa44c0} /* (12, 15, 15) {real, imag} */,
  {32'h410fc737, 32'hbe807443} /* (12, 15, 14) {real, imag} */,
  {32'hc02b52a1, 32'hc10dcf84} /* (12, 15, 13) {real, imag} */,
  {32'h403f5101, 32'hbf17386a} /* (12, 15, 12) {real, imag} */,
  {32'hc0a089b1, 32'hc08afeee} /* (12, 15, 11) {real, imag} */,
  {32'hc037db01, 32'h3e3abca9} /* (12, 15, 10) {real, imag} */,
  {32'hbf790f31, 32'hbf7a4538} /* (12, 15, 9) {real, imag} */,
  {32'hc06e501c, 32'hbfbb5d84} /* (12, 15, 8) {real, imag} */,
  {32'h3fc6afc5, 32'h3f19db58} /* (12, 15, 7) {real, imag} */,
  {32'h4074f888, 32'hc1053dc1} /* (12, 15, 6) {real, imag} */,
  {32'hc074643f, 32'h3e628677} /* (12, 15, 5) {real, imag} */,
  {32'h3fe8c785, 32'h40e545f1} /* (12, 15, 4) {real, imag} */,
  {32'hc0993e60, 32'h41325d64} /* (12, 15, 3) {real, imag} */,
  {32'hc0efc3d8, 32'hbf9daba5} /* (12, 15, 2) {real, imag} */,
  {32'h3e0e403e, 32'hc17e5fe9} /* (12, 15, 1) {real, imag} */,
  {32'hc06d1897, 32'h400b483b} /* (12, 15, 0) {real, imag} */,
  {32'h4030c5d2, 32'hc0528983} /* (12, 14, 15) {real, imag} */,
  {32'h405ec1b6, 32'h405ce535} /* (12, 14, 14) {real, imag} */,
  {32'h40b081ef, 32'h409a82b1} /* (12, 14, 13) {real, imag} */,
  {32'hbf70fcee, 32'h4102bd59} /* (12, 14, 12) {real, imag} */,
  {32'hbf95a8cf, 32'h40607e30} /* (12, 14, 11) {real, imag} */,
  {32'h40f9282c, 32'hc0cb8cc5} /* (12, 14, 10) {real, imag} */,
  {32'hc093cd77, 32'h3fc7280f} /* (12, 14, 9) {real, imag} */,
  {32'h40e3fd98, 32'hbfb7934c} /* (12, 14, 8) {real, imag} */,
  {32'hbf64a094, 32'hbfa6876f} /* (12, 14, 7) {real, imag} */,
  {32'hbeddd4fc, 32'h3fee4509} /* (12, 14, 6) {real, imag} */,
  {32'h40b05a00, 32'hc0346391} /* (12, 14, 5) {real, imag} */,
  {32'h3fc4af1a, 32'hc081436c} /* (12, 14, 4) {real, imag} */,
  {32'h413487d1, 32'hc0a03e53} /* (12, 14, 3) {real, imag} */,
  {32'hc00eed5d, 32'h41171dc9} /* (12, 14, 2) {real, imag} */,
  {32'h40a41d99, 32'hc0fb52d9} /* (12, 14, 1) {real, imag} */,
  {32'hc12baba7, 32'h40d9c1e4} /* (12, 14, 0) {real, imag} */,
  {32'hc00a594b, 32'hc0d74b8d} /* (12, 13, 15) {real, imag} */,
  {32'h4055943c, 32'hc04a858c} /* (12, 13, 14) {real, imag} */,
  {32'hbe46ca70, 32'h4085d0f6} /* (12, 13, 13) {real, imag} */,
  {32'hc1276831, 32'hc04efd52} /* (12, 13, 12) {real, imag} */,
  {32'h4118eb86, 32'hc0f3b68e} /* (12, 13, 11) {real, imag} */,
  {32'h40e82b87, 32'hbf89771f} /* (12, 13, 10) {real, imag} */,
  {32'hc012a630, 32'hc0b5dfb6} /* (12, 13, 9) {real, imag} */,
  {32'h4043d872, 32'h3f0d72e8} /* (12, 13, 8) {real, imag} */,
  {32'h4094c30c, 32'hbf8f7eab} /* (12, 13, 7) {real, imag} */,
  {32'h40f3c561, 32'h40ee8d46} /* (12, 13, 6) {real, imag} */,
  {32'h409c9222, 32'hc06265c5} /* (12, 13, 5) {real, imag} */,
  {32'hc0426572, 32'h407f93ab} /* (12, 13, 4) {real, imag} */,
  {32'hc09d302a, 32'h40a589ce} /* (12, 13, 3) {real, imag} */,
  {32'h3fa8b7d6, 32'h3fec6341} /* (12, 13, 2) {real, imag} */,
  {32'hc0dd0425, 32'hc015ce32} /* (12, 13, 1) {real, imag} */,
  {32'h4079fb3a, 32'hbfb731a9} /* (12, 13, 0) {real, imag} */,
  {32'h4084893f, 32'hc014fc4b} /* (12, 12, 15) {real, imag} */,
  {32'hc00e9eb3, 32'hc08021ed} /* (12, 12, 14) {real, imag} */,
  {32'hc0a8dd8e, 32'h4073b27b} /* (12, 12, 13) {real, imag} */,
  {32'h4073f26c, 32'hbf1c6210} /* (12, 12, 12) {real, imag} */,
  {32'h40e36815, 32'hbee8dc0a} /* (12, 12, 11) {real, imag} */,
  {32'h40163af5, 32'h40c3edb9} /* (12, 12, 10) {real, imag} */,
  {32'h4053c391, 32'h4018b5d3} /* (12, 12, 9) {real, imag} */,
  {32'h40502110, 32'h3c7e881f} /* (12, 12, 8) {real, imag} */,
  {32'hbe14dbf8, 32'hc11e2092} /* (12, 12, 7) {real, imag} */,
  {32'hc173743b, 32'h4098905e} /* (12, 12, 6) {real, imag} */,
  {32'h3f82b094, 32'hc09d4efa} /* (12, 12, 5) {real, imag} */,
  {32'h4082e17d, 32'hc07f8c39} /* (12, 12, 4) {real, imag} */,
  {32'hc028cd08, 32'hc1129296} /* (12, 12, 3) {real, imag} */,
  {32'h405396a3, 32'hc092dce8} /* (12, 12, 2) {real, imag} */,
  {32'h41249b5e, 32'h406a3393} /* (12, 12, 1) {real, imag} */,
  {32'h409930ee, 32'hc000c00a} /* (12, 12, 0) {real, imag} */,
  {32'h3ea1056b, 32'hc0b15b09} /* (12, 11, 15) {real, imag} */,
  {32'hbde1c001, 32'h40ab5568} /* (12, 11, 14) {real, imag} */,
  {32'hc1598ee7, 32'hc16729ae} /* (12, 11, 13) {real, imag} */,
  {32'h403706b9, 32'hc0bc2daf} /* (12, 11, 12) {real, imag} */,
  {32'h40d6ebfc, 32'h40edf348} /* (12, 11, 11) {real, imag} */,
  {32'h40207a74, 32'hc01d251f} /* (12, 11, 10) {real, imag} */,
  {32'h40b5f5ac, 32'hbfe37f5e} /* (12, 11, 9) {real, imag} */,
  {32'h404dab87, 32'hc060e9c1} /* (12, 11, 8) {real, imag} */,
  {32'h40ad004b, 32'h3fc21685} /* (12, 11, 7) {real, imag} */,
  {32'hc0421138, 32'h410c7ad3} /* (12, 11, 6) {real, imag} */,
  {32'hc12f8c24, 32'hbfb38bcf} /* (12, 11, 5) {real, imag} */,
  {32'h40402017, 32'h40c57d01} /* (12, 11, 4) {real, imag} */,
  {32'hc02225c2, 32'h40d1c1db} /* (12, 11, 3) {real, imag} */,
  {32'hc00faf28, 32'h40ca6d71} /* (12, 11, 2) {real, imag} */,
  {32'hc170194a, 32'hc07d05f9} /* (12, 11, 1) {real, imag} */,
  {32'hbd802de5, 32'hbfe57e79} /* (12, 11, 0) {real, imag} */,
  {32'hbf48c932, 32'h410fd874} /* (12, 10, 15) {real, imag} */,
  {32'h411357af, 32'h405c4569} /* (12, 10, 14) {real, imag} */,
  {32'hc08fc80e, 32'h410ed02e} /* (12, 10, 13) {real, imag} */,
  {32'h4106237c, 32'hc15de5db} /* (12, 10, 12) {real, imag} */,
  {32'hc05f3abf, 32'hc099c131} /* (12, 10, 11) {real, imag} */,
  {32'h40b26166, 32'hc020f0ec} /* (12, 10, 10) {real, imag} */,
  {32'hbfc34536, 32'h3d2735be} /* (12, 10, 9) {real, imag} */,
  {32'h40beba6b, 32'hc06c6f5c} /* (12, 10, 8) {real, imag} */,
  {32'hc07ec43d, 32'h4104a325} /* (12, 10, 7) {real, imag} */,
  {32'h402797bf, 32'hbf0adb9c} /* (12, 10, 6) {real, imag} */,
  {32'hc00119a0, 32'h3fe104dd} /* (12, 10, 5) {real, imag} */,
  {32'hc12450f2, 32'h40466804} /* (12, 10, 4) {real, imag} */,
  {32'hbf03fbc1, 32'hbf372b57} /* (12, 10, 3) {real, imag} */,
  {32'hbf1cee19, 32'h40965762} /* (12, 10, 2) {real, imag} */,
  {32'hbf9245c6, 32'hc162144a} /* (12, 10, 1) {real, imag} */,
  {32'hc0b394b5, 32'hc15263cf} /* (12, 10, 0) {real, imag} */,
  {32'h3fdeab87, 32'h40c16ea8} /* (12, 9, 15) {real, imag} */,
  {32'h40ac21e5, 32'hbfc0f621} /* (12, 9, 14) {real, imag} */,
  {32'hbff8deea, 32'hc06ca059} /* (12, 9, 13) {real, imag} */,
  {32'hbf5d5b3b, 32'hc083ba4f} /* (12, 9, 12) {real, imag} */,
  {32'h40b6b4f3, 32'h404a73eb} /* (12, 9, 11) {real, imag} */,
  {32'hc127d04b, 32'hc07c6b0f} /* (12, 9, 10) {real, imag} */,
  {32'hbfb520d2, 32'hc07fb937} /* (12, 9, 9) {real, imag} */,
  {32'h3feec3ba, 32'hbf2e2ba9} /* (12, 9, 8) {real, imag} */,
  {32'h40e43883, 32'hc0442a7b} /* (12, 9, 7) {real, imag} */,
  {32'h3f0f759d, 32'h40b7f154} /* (12, 9, 6) {real, imag} */,
  {32'hbf82ac79, 32'hbf84d7c7} /* (12, 9, 5) {real, imag} */,
  {32'hc151c892, 32'h3e1ff026} /* (12, 9, 4) {real, imag} */,
  {32'h4045d73e, 32'h3f602a10} /* (12, 9, 3) {real, imag} */,
  {32'hc0914026, 32'hc05d6458} /* (12, 9, 2) {real, imag} */,
  {32'hbecd39f8, 32'hc0d3b745} /* (12, 9, 1) {real, imag} */,
  {32'h3fde0eba, 32'h4105c267} /* (12, 9, 0) {real, imag} */,
  {32'h406002ad, 32'h3f1bf36c} /* (12, 8, 15) {real, imag} */,
  {32'h404aece7, 32'h405764a8} /* (12, 8, 14) {real, imag} */,
  {32'hbf717e49, 32'hc03b7886} /* (12, 8, 13) {real, imag} */,
  {32'h4032bcd2, 32'h3f7fa7a6} /* (12, 8, 12) {real, imag} */,
  {32'hc0bc4ead, 32'h40a88f17} /* (12, 8, 11) {real, imag} */,
  {32'h40ebff79, 32'hc08d38fd} /* (12, 8, 10) {real, imag} */,
  {32'hbf41b754, 32'hbe9da841} /* (12, 8, 9) {real, imag} */,
  {32'hc04a6665, 32'hc01353a1} /* (12, 8, 8) {real, imag} */,
  {32'h3f193052, 32'h403336a9} /* (12, 8, 7) {real, imag} */,
  {32'h41264451, 32'hc0a60dd5} /* (12, 8, 6) {real, imag} */,
  {32'hbfdc28ec, 32'hc05f550c} /* (12, 8, 5) {real, imag} */,
  {32'hc06ee6b0, 32'hc0e1e6f6} /* (12, 8, 4) {real, imag} */,
  {32'hbf5509ba, 32'h3faad099} /* (12, 8, 3) {real, imag} */,
  {32'hc026fe1d, 32'hbe63ce1a} /* (12, 8, 2) {real, imag} */,
  {32'h40d6081b, 32'hbe23cbda} /* (12, 8, 1) {real, imag} */,
  {32'hc0bb3ab9, 32'hbf826da2} /* (12, 8, 0) {real, imag} */,
  {32'hc1300528, 32'hc0519843} /* (12, 7, 15) {real, imag} */,
  {32'h405b57c7, 32'h40370c66} /* (12, 7, 14) {real, imag} */,
  {32'hbea7f3dc, 32'h4023d62a} /* (12, 7, 13) {real, imag} */,
  {32'hc00f7bb6, 32'h3d5118a5} /* (12, 7, 12) {real, imag} */,
  {32'hbfe46f45, 32'hc04a8c5c} /* (12, 7, 11) {real, imag} */,
  {32'h407e81b3, 32'h4119a977} /* (12, 7, 10) {real, imag} */,
  {32'hbfcf93d2, 32'hbf8b9aac} /* (12, 7, 9) {real, imag} */,
  {32'h3fa2f7c1, 32'hc07aec84} /* (12, 7, 8) {real, imag} */,
  {32'hbee2b952, 32'h3d53c2e3} /* (12, 7, 7) {real, imag} */,
  {32'hbff73308, 32'hc0eeba0f} /* (12, 7, 6) {real, imag} */,
  {32'h409751f0, 32'h3ff8eedb} /* (12, 7, 5) {real, imag} */,
  {32'h4044dded, 32'hc0011e57} /* (12, 7, 4) {real, imag} */,
  {32'hc08dc826, 32'h3f17e050} /* (12, 7, 3) {real, imag} */,
  {32'hc001d18d, 32'hc0668a33} /* (12, 7, 2) {real, imag} */,
  {32'h40553337, 32'h3f9ee217} /* (12, 7, 1) {real, imag} */,
  {32'h3cad9d20, 32'h3fc58c74} /* (12, 7, 0) {real, imag} */,
  {32'h40917842, 32'hc074a5ee} /* (12, 6, 15) {real, imag} */,
  {32'h4023bdf6, 32'hc12fbd85} /* (12, 6, 14) {real, imag} */,
  {32'h40e59d2e, 32'hbf71bae1} /* (12, 6, 13) {real, imag} */,
  {32'h401c7126, 32'h40baf6fb} /* (12, 6, 12) {real, imag} */,
  {32'h411b36d4, 32'h40d1b3f1} /* (12, 6, 11) {real, imag} */,
  {32'hc09cea2b, 32'hbfd9f200} /* (12, 6, 10) {real, imag} */,
  {32'hbfec99e0, 32'hbfa3c271} /* (12, 6, 9) {real, imag} */,
  {32'hbfa39fc0, 32'h4065c839} /* (12, 6, 8) {real, imag} */,
  {32'h3f8d1502, 32'hbffad29a} /* (12, 6, 7) {real, imag} */,
  {32'hc128819f, 32'h400d8a0e} /* (12, 6, 6) {real, imag} */,
  {32'hc06c0b76, 32'hc04cbd92} /* (12, 6, 5) {real, imag} */,
  {32'hc08b06f0, 32'hc0831b1e} /* (12, 6, 4) {real, imag} */,
  {32'h4064a9fc, 32'h3e37b243} /* (12, 6, 3) {real, imag} */,
  {32'h415ae054, 32'h40252f59} /* (12, 6, 2) {real, imag} */,
  {32'hc149af2e, 32'hbf58aada} /* (12, 6, 1) {real, imag} */,
  {32'hc004c443, 32'h402c14c0} /* (12, 6, 0) {real, imag} */,
  {32'hc0eb0c47, 32'h3b365898} /* (12, 5, 15) {real, imag} */,
  {32'h4054e032, 32'hc0a2325b} /* (12, 5, 14) {real, imag} */,
  {32'h3f8934b3, 32'h3f49c05b} /* (12, 5, 13) {real, imag} */,
  {32'h40963d83, 32'h4053d8ca} /* (12, 5, 12) {real, imag} */,
  {32'h3feb6c61, 32'hc02e0221} /* (12, 5, 11) {real, imag} */,
  {32'hc0eb1962, 32'h401733f8} /* (12, 5, 10) {real, imag} */,
  {32'hbfc29454, 32'hbf4847aa} /* (12, 5, 9) {real, imag} */,
  {32'h3f5c5b55, 32'hc092b50c} /* (12, 5, 8) {real, imag} */,
  {32'hc0d7d0ae, 32'h3eef032e} /* (12, 5, 7) {real, imag} */,
  {32'h3f6663e9, 32'hc059922b} /* (12, 5, 6) {real, imag} */,
  {32'h3f4ac918, 32'h409f6531} /* (12, 5, 5) {real, imag} */,
  {32'h40a8db77, 32'hc0f18ae0} /* (12, 5, 4) {real, imag} */,
  {32'hc0ff1239, 32'hc06314e5} /* (12, 5, 3) {real, imag} */,
  {32'hbf08b9c4, 32'h40f5845e} /* (12, 5, 2) {real, imag} */,
  {32'hc16b65cb, 32'h410c76eb} /* (12, 5, 1) {real, imag} */,
  {32'hc0c4b502, 32'hc101c0ad} /* (12, 5, 0) {real, imag} */,
  {32'h40ba0f28, 32'hc0c7bce7} /* (12, 4, 15) {real, imag} */,
  {32'hc10c3286, 32'hc09cb6f2} /* (12, 4, 14) {real, imag} */,
  {32'h4059edbc, 32'hc0a75371} /* (12, 4, 13) {real, imag} */,
  {32'h3eedd483, 32'hc0134704} /* (12, 4, 12) {real, imag} */,
  {32'h407ff0ff, 32'hc074cda8} /* (12, 4, 11) {real, imag} */,
  {32'h411f013c, 32'hc0b07849} /* (12, 4, 10) {real, imag} */,
  {32'hbf3c7360, 32'h40a01d0e} /* (12, 4, 9) {real, imag} */,
  {32'h40aa5658, 32'hbfc82d1f} /* (12, 4, 8) {real, imag} */,
  {32'h409f7b31, 32'hc0c2278e} /* (12, 4, 7) {real, imag} */,
  {32'hbe8122f3, 32'h3f905af1} /* (12, 4, 6) {real, imag} */,
  {32'h404d8202, 32'h3f8b5d2c} /* (12, 4, 5) {real, imag} */,
  {32'hc1781de9, 32'hbe14c422} /* (12, 4, 4) {real, imag} */,
  {32'h4006ed3b, 32'h3f7b4046} /* (12, 4, 3) {real, imag} */,
  {32'hc0225711, 32'h41025d6a} /* (12, 4, 2) {real, imag} */,
  {32'hbef7055e, 32'h3f95d681} /* (12, 4, 1) {real, imag} */,
  {32'hbfe1f851, 32'hc08d263d} /* (12, 4, 0) {real, imag} */,
  {32'hc099a64c, 32'h4082d468} /* (12, 3, 15) {real, imag} */,
  {32'h40641d61, 32'hc020e8f7} /* (12, 3, 14) {real, imag} */,
  {32'hbeda50f9, 32'hc0095ce8} /* (12, 3, 13) {real, imag} */,
  {32'h40550532, 32'h3ed76676} /* (12, 3, 12) {real, imag} */,
  {32'h406b6c04, 32'h412a73cd} /* (12, 3, 11) {real, imag} */,
  {32'hc028d546, 32'hc0841ab9} /* (12, 3, 10) {real, imag} */,
  {32'hbf93e6a3, 32'hc0d727ec} /* (12, 3, 9) {real, imag} */,
  {32'hc09fd0d4, 32'h3f10f477} /* (12, 3, 8) {real, imag} */,
  {32'hc0bc8dfe, 32'hc11c1fbf} /* (12, 3, 7) {real, imag} */,
  {32'h411f938f, 32'h40aedd1d} /* (12, 3, 6) {real, imag} */,
  {32'hc08137dd, 32'hc03f85de} /* (12, 3, 5) {real, imag} */,
  {32'hc0b09723, 32'hc01d4549} /* (12, 3, 4) {real, imag} */,
  {32'hc05d5d4c, 32'h40928ed1} /* (12, 3, 3) {real, imag} */,
  {32'hc0688499, 32'hc0f23a05} /* (12, 3, 2) {real, imag} */,
  {32'hc09f6713, 32'hbdb3eee1} /* (12, 3, 1) {real, imag} */,
  {32'h4046d5dd, 32'hbf9def25} /* (12, 3, 0) {real, imag} */,
  {32'hc1706c22, 32'h40be7fd2} /* (12, 2, 15) {real, imag} */,
  {32'h4128a820, 32'hbfc9445a} /* (12, 2, 14) {real, imag} */,
  {32'hc039fa94, 32'hbfa40105} /* (12, 2, 13) {real, imag} */,
  {32'hbe55a7f0, 32'h41025359} /* (12, 2, 12) {real, imag} */,
  {32'hc03c079c, 32'hc0ba282e} /* (12, 2, 11) {real, imag} */,
  {32'h3fa70be7, 32'h40f70abf} /* (12, 2, 10) {real, imag} */,
  {32'hc0efda8e, 32'hbfb7e5a1} /* (12, 2, 9) {real, imag} */,
  {32'hc0181c93, 32'h40840e77} /* (12, 2, 8) {real, imag} */,
  {32'hc01b773d, 32'h40c44475} /* (12, 2, 7) {real, imag} */,
  {32'h40c55617, 32'hc0c85853} /* (12, 2, 6) {real, imag} */,
  {32'hc0af87a9, 32'hc0c0f41c} /* (12, 2, 5) {real, imag} */,
  {32'h3f74a3ff, 32'h3d696fe4} /* (12, 2, 4) {real, imag} */,
  {32'hc02c7e37, 32'hc0d5630a} /* (12, 2, 3) {real, imag} */,
  {32'h410162a9, 32'hc0b9f213} /* (12, 2, 2) {real, imag} */,
  {32'h4123b580, 32'h402ec640} /* (12, 2, 1) {real, imag} */,
  {32'hc0bb6c3f, 32'h417f07f4} /* (12, 2, 0) {real, imag} */,
  {32'h411eac5a, 32'h4123923e} /* (12, 1, 15) {real, imag} */,
  {32'hc14644eb, 32'h3f5b85af} /* (12, 1, 14) {real, imag} */,
  {32'hc0accb95, 32'h3f9c7c5b} /* (12, 1, 13) {real, imag} */,
  {32'h3eb76200, 32'hc0070ca2} /* (12, 1, 12) {real, imag} */,
  {32'hc0ea133a, 32'h4085f286} /* (12, 1, 11) {real, imag} */,
  {32'hc0208ffa, 32'h4013878f} /* (12, 1, 10) {real, imag} */,
  {32'h40bdfde9, 32'h3e9ee513} /* (12, 1, 9) {real, imag} */,
  {32'hc04e39b8, 32'hc06d3bec} /* (12, 1, 8) {real, imag} */,
  {32'hbfde8912, 32'hc056b39d} /* (12, 1, 7) {real, imag} */,
  {32'h3f405a77, 32'h40c7e617} /* (12, 1, 6) {real, imag} */,
  {32'hc085e830, 32'h3f87ab15} /* (12, 1, 5) {real, imag} */,
  {32'h40ef9260, 32'h40c8f8aa} /* (12, 1, 4) {real, imag} */,
  {32'hbea38287, 32'hbebb89bd} /* (12, 1, 3) {real, imag} */,
  {32'h40a78c59, 32'h3ff970b9} /* (12, 1, 2) {real, imag} */,
  {32'h3f3effd0, 32'hc05432d4} /* (12, 1, 1) {real, imag} */,
  {32'h41b49cd3, 32'hc15712b2} /* (12, 1, 0) {real, imag} */,
  {32'h3e3a7b45, 32'h412710ed} /* (12, 0, 15) {real, imag} */,
  {32'hc0179f0f, 32'h3ed144bf} /* (12, 0, 14) {real, imag} */,
  {32'h3f8cc2c5, 32'h40b7cb53} /* (12, 0, 13) {real, imag} */,
  {32'hc0d777a2, 32'h41078757} /* (12, 0, 12) {real, imag} */,
  {32'hbf8abf98, 32'hc124a1dc} /* (12, 0, 11) {real, imag} */,
  {32'hc071f363, 32'h3ee508da} /* (12, 0, 10) {real, imag} */,
  {32'hbfab6815, 32'h406e3bbb} /* (12, 0, 9) {real, imag} */,
  {32'hbefcd082, 32'h3f07f3ed} /* (12, 0, 8) {real, imag} */,
  {32'h40a9fc38, 32'h3ffd70a0} /* (12, 0, 7) {real, imag} */,
  {32'hc017d6bd, 32'h3f3096e4} /* (12, 0, 6) {real, imag} */,
  {32'h40a49e35, 32'h40efd47b} /* (12, 0, 5) {real, imag} */,
  {32'h407aecb7, 32'hc03c805b} /* (12, 0, 4) {real, imag} */,
  {32'h40f4f089, 32'hc134f737} /* (12, 0, 3) {real, imag} */,
  {32'hc11c76bc, 32'h401b958b} /* (12, 0, 2) {real, imag} */,
  {32'hc1525390, 32'h405b795c} /* (12, 0, 1) {real, imag} */,
  {32'hc0b6046b, 32'hbf4872f1} /* (12, 0, 0) {real, imag} */,
  {32'h406a695a, 32'h402a22e1} /* (11, 15, 15) {real, imag} */,
  {32'h405bc194, 32'hc1181ead} /* (11, 15, 14) {real, imag} */,
  {32'hbff6f9be, 32'h412defa8} /* (11, 15, 13) {real, imag} */,
  {32'h3ff49d29, 32'h3fdec1a5} /* (11, 15, 12) {real, imag} */,
  {32'hbfb49d06, 32'h41314697} /* (11, 15, 11) {real, imag} */,
  {32'h40b8ee23, 32'hc06d587e} /* (11, 15, 10) {real, imag} */,
  {32'h3f92e928, 32'hbc84df57} /* (11, 15, 9) {real, imag} */,
  {32'hbfc968da, 32'hbf86304a} /* (11, 15, 8) {real, imag} */,
  {32'hc0be4b8e, 32'hc0a1a1fa} /* (11, 15, 7) {real, imag} */,
  {32'hbf7571e3, 32'h40931eae} /* (11, 15, 6) {real, imag} */,
  {32'hc0108e0e, 32'hc0361d33} /* (11, 15, 5) {real, imag} */,
  {32'h404595cc, 32'hc1039a2b} /* (11, 15, 4) {real, imag} */,
  {32'h4074e298, 32'hc04c31b4} /* (11, 15, 3) {real, imag} */,
  {32'hc162305a, 32'h40fbbc02} /* (11, 15, 2) {real, imag} */,
  {32'h41002885, 32'hc031b43c} /* (11, 15, 1) {real, imag} */,
  {32'h409d6d34, 32'hc1025c39} /* (11, 15, 0) {real, imag} */,
  {32'h415567aa, 32'h409e2c1d} /* (11, 14, 15) {real, imag} */,
  {32'h413825d3, 32'h40a7d5d6} /* (11, 14, 14) {real, imag} */,
  {32'h410a46f9, 32'h3ef1ff30} /* (11, 14, 13) {real, imag} */,
  {32'hc0ccd9f6, 32'hc0183a4f} /* (11, 14, 12) {real, imag} */,
  {32'hc0ae4c74, 32'hbf19cad3} /* (11, 14, 11) {real, imag} */,
  {32'h403b2521, 32'h40904956} /* (11, 14, 10) {real, imag} */,
  {32'hc09b92f6, 32'hbfada953} /* (11, 14, 9) {real, imag} */,
  {32'hbf43ed65, 32'h3df29da4} /* (11, 14, 8) {real, imag} */,
  {32'h3ed9b0e0, 32'h40965d27} /* (11, 14, 7) {real, imag} */,
  {32'hc1167f26, 32'hc107406c} /* (11, 14, 6) {real, imag} */,
  {32'h3fed8916, 32'hc0ccc265} /* (11, 14, 5) {real, imag} */,
  {32'hc07712ed, 32'h41334e83} /* (11, 14, 4) {real, imag} */,
  {32'hc0ece269, 32'hc0254d90} /* (11, 14, 3) {real, imag} */,
  {32'hbfdb03de, 32'hc0ca0af1} /* (11, 14, 2) {real, imag} */,
  {32'h40eb73a5, 32'hc0b56247} /* (11, 14, 1) {real, imag} */,
  {32'h3fcb00f7, 32'h3f4bcbf8} /* (11, 14, 0) {real, imag} */,
  {32'hc0a9de95, 32'h3f04773c} /* (11, 13, 15) {real, imag} */,
  {32'hbf48bb72, 32'hc01c4ed5} /* (11, 13, 14) {real, imag} */,
  {32'h41071e5c, 32'hc0e444fb} /* (11, 13, 13) {real, imag} */,
  {32'hc0b6a924, 32'hbfa875ef} /* (11, 13, 12) {real, imag} */,
  {32'hbfe0ef54, 32'h414fd879} /* (11, 13, 11) {real, imag} */,
  {32'h409c5db5, 32'h3e31ab7f} /* (11, 13, 10) {real, imag} */,
  {32'hbfe3051e, 32'hc00acb31} /* (11, 13, 9) {real, imag} */,
  {32'hbee74252, 32'hc07c03ef} /* (11, 13, 8) {real, imag} */,
  {32'hc048b807, 32'hc05fd6f6} /* (11, 13, 7) {real, imag} */,
  {32'h4117b350, 32'h3f5a1f06} /* (11, 13, 6) {real, imag} */,
  {32'h412244cc, 32'hc03304de} /* (11, 13, 5) {real, imag} */,
  {32'h40e04968, 32'hbfdc6f4e} /* (11, 13, 4) {real, imag} */,
  {32'h40a9b4a1, 32'h401715b2} /* (11, 13, 3) {real, imag} */,
  {32'h3f65cc58, 32'h3ddb704b} /* (11, 13, 2) {real, imag} */,
  {32'h4082d4e2, 32'hc087fbf7} /* (11, 13, 1) {real, imag} */,
  {32'h3ff10c26, 32'h403c6c81} /* (11, 13, 0) {real, imag} */,
  {32'hc0ff5b38, 32'h408118a2} /* (11, 12, 15) {real, imag} */,
  {32'hc10294ac, 32'hc0547d64} /* (11, 12, 14) {real, imag} */,
  {32'hbf409ff6, 32'h409fd414} /* (11, 12, 13) {real, imag} */,
  {32'hc0d0e4fc, 32'h3dd33688} /* (11, 12, 12) {real, imag} */,
  {32'h40a2159a, 32'h3eb65a2f} /* (11, 12, 11) {real, imag} */,
  {32'hbf94d24d, 32'h3d878350} /* (11, 12, 10) {real, imag} */,
  {32'h409163c0, 32'hc0dc1794} /* (11, 12, 9) {real, imag} */,
  {32'hbf7654d3, 32'hbc4b4563} /* (11, 12, 8) {real, imag} */,
  {32'h3fa863e3, 32'h4016ffae} /* (11, 12, 7) {real, imag} */,
  {32'h4136c3cc, 32'hc0263f62} /* (11, 12, 6) {real, imag} */,
  {32'hc09ff3e9, 32'h4092ce8a} /* (11, 12, 5) {real, imag} */,
  {32'h3f58eae4, 32'hc08d3511} /* (11, 12, 4) {real, imag} */,
  {32'h40345fa0, 32'h40c6fe6e} /* (11, 12, 3) {real, imag} */,
  {32'h3f14940f, 32'h402a81ec} /* (11, 12, 2) {real, imag} */,
  {32'hbec49070, 32'h4148c74a} /* (11, 12, 1) {real, imag} */,
  {32'hc0217bf6, 32'hbf8d81ba} /* (11, 12, 0) {real, imag} */,
  {32'h412aa69b, 32'hc05e9b15} /* (11, 11, 15) {real, imag} */,
  {32'hc0c263a2, 32'h403f63a2} /* (11, 11, 14) {real, imag} */,
  {32'hbfe564d0, 32'hc0dc4322} /* (11, 11, 13) {real, imag} */,
  {32'h40cd99ab, 32'h40e12b05} /* (11, 11, 12) {real, imag} */,
  {32'h40d86de2, 32'h3f75315d} /* (11, 11, 11) {real, imag} */,
  {32'hc0fe860d, 32'h401e3ce3} /* (11, 11, 10) {real, imag} */,
  {32'hc0b324f5, 32'hbfb68a4a} /* (11, 11, 9) {real, imag} */,
  {32'hbb2bd2e5, 32'h409f7f1a} /* (11, 11, 8) {real, imag} */,
  {32'h3fa8fe07, 32'h409457a3} /* (11, 11, 7) {real, imag} */,
  {32'h40112cdc, 32'h40b0278d} /* (11, 11, 6) {real, imag} */,
  {32'h3f64839e, 32'h40d34a59} /* (11, 11, 5) {real, imag} */,
  {32'hc02fd0a6, 32'h404a6f17} /* (11, 11, 4) {real, imag} */,
  {32'hc0501efd, 32'hc11ad6c6} /* (11, 11, 3) {real, imag} */,
  {32'hbf9774a6, 32'hc12c7114} /* (11, 11, 2) {real, imag} */,
  {32'hbf0e9128, 32'h40ea2645} /* (11, 11, 1) {real, imag} */,
  {32'hc0a04e9f, 32'h3ebf80e7} /* (11, 11, 0) {real, imag} */,
  {32'hc13fd900, 32'hc05c8b34} /* (11, 10, 15) {real, imag} */,
  {32'hbf3372ef, 32'hbe2a11f2} /* (11, 10, 14) {real, imag} */,
  {32'h408c8bed, 32'hc05d9219} /* (11, 10, 13) {real, imag} */,
  {32'h400b6ba9, 32'h4118da98} /* (11, 10, 12) {real, imag} */,
  {32'hc10e9611, 32'hc00a270f} /* (11, 10, 11) {real, imag} */,
  {32'hc10438bb, 32'hbf9ef9da} /* (11, 10, 10) {real, imag} */,
  {32'h40182ea0, 32'hbf477673} /* (11, 10, 9) {real, imag} */,
  {32'hbf1e7162, 32'h40bbe68d} /* (11, 10, 8) {real, imag} */,
  {32'hc097c033, 32'hc0799482} /* (11, 10, 7) {real, imag} */,
  {32'hbfe109f4, 32'h408484b1} /* (11, 10, 6) {real, imag} */,
  {32'h3f888182, 32'hc10200af} /* (11, 10, 5) {real, imag} */,
  {32'h4010e7c2, 32'h4077d62a} /* (11, 10, 4) {real, imag} */,
  {32'hc0a7495f, 32'h406f4ce0} /* (11, 10, 3) {real, imag} */,
  {32'hc139c713, 32'hbd61a7af} /* (11, 10, 2) {real, imag} */,
  {32'hc085940c, 32'hc0157d81} /* (11, 10, 1) {real, imag} */,
  {32'h40e9a601, 32'h402dcd49} /* (11, 10, 0) {real, imag} */,
  {32'hc0938435, 32'hc0b660d1} /* (11, 9, 15) {real, imag} */,
  {32'h401a3054, 32'hc076bdd9} /* (11, 9, 14) {real, imag} */,
  {32'h40c92d4b, 32'hc00822e2} /* (11, 9, 13) {real, imag} */,
  {32'h40abbad0, 32'h410cbbad} /* (11, 9, 12) {real, imag} */,
  {32'hbfb85363, 32'h3f7f4644} /* (11, 9, 11) {real, imag} */,
  {32'hc0c06ccb, 32'h40c325a3} /* (11, 9, 10) {real, imag} */,
  {32'h40c827f3, 32'hc028f6a5} /* (11, 9, 9) {real, imag} */,
  {32'h4094aec0, 32'hc05b8b1a} /* (11, 9, 8) {real, imag} */,
  {32'hc030e8e8, 32'h40815776} /* (11, 9, 7) {real, imag} */,
  {32'hc0802a35, 32'hc069bb1b} /* (11, 9, 6) {real, imag} */,
  {32'h406928e3, 32'hc08ec0c7} /* (11, 9, 5) {real, imag} */,
  {32'hc00d2178, 32'h3f59ccb7} /* (11, 9, 4) {real, imag} */,
  {32'h40781707, 32'h40c32605} /* (11, 9, 3) {real, imag} */,
  {32'hc014c713, 32'hc0113621} /* (11, 9, 2) {real, imag} */,
  {32'hc01e7d24, 32'h3eaa6fe8} /* (11, 9, 1) {real, imag} */,
  {32'h3f293aef, 32'hc0791faf} /* (11, 9, 0) {real, imag} */,
  {32'h400b462a, 32'hc08cd555} /* (11, 8, 15) {real, imag} */,
  {32'hc08163f1, 32'h4010adc1} /* (11, 8, 14) {real, imag} */,
  {32'h4058cf91, 32'hbf890541} /* (11, 8, 13) {real, imag} */,
  {32'hbfd7312d, 32'h402707bf} /* (11, 8, 12) {real, imag} */,
  {32'h3a88daf7, 32'h4022c0b7} /* (11, 8, 11) {real, imag} */,
  {32'hbfe4af93, 32'hbda3e51b} /* (11, 8, 10) {real, imag} */,
  {32'h409539bd, 32'h4000d86f} /* (11, 8, 9) {real, imag} */,
  {32'h3d058620, 32'hc011c020} /* (11, 8, 8) {real, imag} */,
  {32'hc08ca80b, 32'hc0a9bc9c} /* (11, 8, 7) {real, imag} */,
  {32'hc05b201a, 32'h4038b552} /* (11, 8, 6) {real, imag} */,
  {32'h40e19ccb, 32'h406bcee1} /* (11, 8, 5) {real, imag} */,
  {32'h40ef33ff, 32'hbe6bbe05} /* (11, 8, 4) {real, imag} */,
  {32'h40b6d0e3, 32'hc073e0ef} /* (11, 8, 3) {real, imag} */,
  {32'h40057087, 32'h3f37e4de} /* (11, 8, 2) {real, imag} */,
  {32'hbf73edbf, 32'h40e02ec9} /* (11, 8, 1) {real, imag} */,
  {32'hc053f04c, 32'hc07417de} /* (11, 8, 0) {real, imag} */,
  {32'h40d2e79b, 32'h40a1e8fd} /* (11, 7, 15) {real, imag} */,
  {32'hc0db1d13, 32'hc00de8c2} /* (11, 7, 14) {real, imag} */,
  {32'hbee6990a, 32'h3fb276b9} /* (11, 7, 13) {real, imag} */,
  {32'h3ef0cdca, 32'hc0350b72} /* (11, 7, 12) {real, imag} */,
  {32'hc09707c6, 32'h3fedba5e} /* (11, 7, 11) {real, imag} */,
  {32'h402ca0af, 32'hc04fb022} /* (11, 7, 10) {real, imag} */,
  {32'hc0c69534, 32'h3fbad0e0} /* (11, 7, 9) {real, imag} */,
  {32'hc04b440c, 32'h40f0ab3d} /* (11, 7, 8) {real, imag} */,
  {32'h4010eb51, 32'h401d9459} /* (11, 7, 7) {real, imag} */,
  {32'h3facb8b0, 32'h40df4759} /* (11, 7, 6) {real, imag} */,
  {32'hbfa85070, 32'hc079dd28} /* (11, 7, 5) {real, imag} */,
  {32'hc04ed7a6, 32'hc10b4a74} /* (11, 7, 4) {real, imag} */,
  {32'h3fe8e818, 32'h40a7fd9f} /* (11, 7, 3) {real, imag} */,
  {32'h3ffe536e, 32'h3fb8f510} /* (11, 7, 2) {real, imag} */,
  {32'h3f8bdc33, 32'h4005c69c} /* (11, 7, 1) {real, imag} */,
  {32'h3e9a8d38, 32'hc0a6e2c2} /* (11, 7, 0) {real, imag} */,
  {32'hbf0a301a, 32'hc11ddbfe} /* (11, 6, 15) {real, imag} */,
  {32'h40100b48, 32'hc05f959b} /* (11, 6, 14) {real, imag} */,
  {32'h3fa2780a, 32'hc0f0053a} /* (11, 6, 13) {real, imag} */,
  {32'h40a96624, 32'h408e6083} /* (11, 6, 12) {real, imag} */,
  {32'h40a3c469, 32'h4127cab8} /* (11, 6, 11) {real, imag} */,
  {32'hc099c31d, 32'hc01c5f65} /* (11, 6, 10) {real, imag} */,
  {32'h3f50e12d, 32'h404b0a6c} /* (11, 6, 9) {real, imag} */,
  {32'h3e80d6b8, 32'hc051d688} /* (11, 6, 8) {real, imag} */,
  {32'hc062346d, 32'h3ff40115} /* (11, 6, 7) {real, imag} */,
  {32'h3fe71f5c, 32'h3ecbfd8b} /* (11, 6, 6) {real, imag} */,
  {32'h40cbde19, 32'hc057811c} /* (11, 6, 5) {real, imag} */,
  {32'hc0456fca, 32'hc06c6797} /* (11, 6, 4) {real, imag} */,
  {32'h4047c6c9, 32'hc09fd691} /* (11, 6, 3) {real, imag} */,
  {32'h4035916d, 32'hc0c126a5} /* (11, 6, 2) {real, imag} */,
  {32'hc08b212e, 32'hc05cf036} /* (11, 6, 1) {real, imag} */,
  {32'hc0c804f2, 32'h4081374b} /* (11, 6, 0) {real, imag} */,
  {32'h3fb02741, 32'hc083a9e7} /* (11, 5, 15) {real, imag} */,
  {32'hbfda8f36, 32'h416bc2dc} /* (11, 5, 14) {real, imag} */,
  {32'h3f2263f8, 32'hc0d1f1e8} /* (11, 5, 13) {real, imag} */,
  {32'h3f70ff71, 32'hc0810eaf} /* (11, 5, 12) {real, imag} */,
  {32'h40e6beac, 32'h40607d44} /* (11, 5, 11) {real, imag} */,
  {32'hc109e2c9, 32'hbf4c1972} /* (11, 5, 10) {real, imag} */,
  {32'hbf1fd540, 32'h40c166c0} /* (11, 5, 9) {real, imag} */,
  {32'hc0841f8c, 32'h40328ca8} /* (11, 5, 8) {real, imag} */,
  {32'h3fea5039, 32'h40ad34c7} /* (11, 5, 7) {real, imag} */,
  {32'h3eddb8b3, 32'hbf0f833a} /* (11, 5, 6) {real, imag} */,
  {32'hbfc6c6e1, 32'hc0984d9c} /* (11, 5, 5) {real, imag} */,
  {32'hc06df3a4, 32'hc0d419d3} /* (11, 5, 4) {real, imag} */,
  {32'hbf09d576, 32'hbfc5851f} /* (11, 5, 3) {real, imag} */,
  {32'hc0b2eec9, 32'h40efb792} /* (11, 5, 2) {real, imag} */,
  {32'h3f477123, 32'hc04a9503} /* (11, 5, 1) {real, imag} */,
  {32'h4097f439, 32'h405931a8} /* (11, 5, 0) {real, imag} */,
  {32'hc054154a, 32'h3f5f838e} /* (11, 4, 15) {real, imag} */,
  {32'hc10b0939, 32'h3f2879f1} /* (11, 4, 14) {real, imag} */,
  {32'h40048715, 32'hc06379c3} /* (11, 4, 13) {real, imag} */,
  {32'hc0176d8c, 32'h4068baf8} /* (11, 4, 12) {real, imag} */,
  {32'hc0d29ed5, 32'hc10539da} /* (11, 4, 11) {real, imag} */,
  {32'h40be17d1, 32'h40fab5c7} /* (11, 4, 10) {real, imag} */,
  {32'hc09e5a25, 32'h40b3466f} /* (11, 4, 9) {real, imag} */,
  {32'h4028b071, 32'hc0afe22c} /* (11, 4, 8) {real, imag} */,
  {32'hc0f29573, 32'hc04b553a} /* (11, 4, 7) {real, imag} */,
  {32'h3ff4ed63, 32'hc10110b6} /* (11, 4, 6) {real, imag} */,
  {32'hbfbebc3b, 32'h40c5e84f} /* (11, 4, 5) {real, imag} */,
  {32'h40bf9708, 32'hbe12c02b} /* (11, 4, 4) {real, imag} */,
  {32'h400ad92e, 32'hc082242a} /* (11, 4, 3) {real, imag} */,
  {32'h41084e61, 32'h40990be5} /* (11, 4, 2) {real, imag} */,
  {32'h3faba832, 32'h3f3884d4} /* (11, 4, 1) {real, imag} */,
  {32'h4096f19a, 32'hc0477501} /* (11, 4, 0) {real, imag} */,
  {32'hc00c28c6, 32'hbf18be7b} /* (11, 3, 15) {real, imag} */,
  {32'h40dbced6, 32'h411de712} /* (11, 3, 14) {real, imag} */,
  {32'h402ea681, 32'hc0a65c7c} /* (11, 3, 13) {real, imag} */,
  {32'hbfb1b785, 32'h40ca569e} /* (11, 3, 12) {real, imag} */,
  {32'h4085ba9b, 32'hc09f02f8} /* (11, 3, 11) {real, imag} */,
  {32'hc0f12eba, 32'hbfb2476a} /* (11, 3, 10) {real, imag} */,
  {32'hbea92559, 32'h3f18009f} /* (11, 3, 9) {real, imag} */,
  {32'h3f28e9cd, 32'hbf0492e4} /* (11, 3, 8) {real, imag} */,
  {32'h3fa8279c, 32'hc022ab8c} /* (11, 3, 7) {real, imag} */,
  {32'hbff8f681, 32'h406186fc} /* (11, 3, 6) {real, imag} */,
  {32'h41017e70, 32'hc03d2c1d} /* (11, 3, 5) {real, imag} */,
  {32'h4033b9d4, 32'h40a2e666} /* (11, 3, 4) {real, imag} */,
  {32'h403b45a1, 32'h40a34135} /* (11, 3, 3) {real, imag} */,
  {32'hc09bd049, 32'h4020ced7} /* (11, 3, 2) {real, imag} */,
  {32'h40633218, 32'hc0803132} /* (11, 3, 1) {real, imag} */,
  {32'hbffd7526, 32'hbf75d0ff} /* (11, 3, 0) {real, imag} */,
  {32'h4093710e, 32'h3fd16966} /* (11, 2, 15) {real, imag} */,
  {32'h3f410110, 32'hc0c62d31} /* (11, 2, 14) {real, imag} */,
  {32'hc0cc2f25, 32'h411bc6d2} /* (11, 2, 13) {real, imag} */,
  {32'hbf526e52, 32'hc0b49eec} /* (11, 2, 12) {real, imag} */,
  {32'h40ab8a81, 32'hc10da436} /* (11, 2, 11) {real, imag} */,
  {32'h412846b4, 32'hc0bcb93a} /* (11, 2, 10) {real, imag} */,
  {32'hbf6f163c, 32'h403f6ada} /* (11, 2, 9) {real, imag} */,
  {32'h4084c774, 32'h3fc8508b} /* (11, 2, 8) {real, imag} */,
  {32'h410c6495, 32'hc14b85cc} /* (11, 2, 7) {real, imag} */,
  {32'hc1068bdd, 32'h408b3115} /* (11, 2, 6) {real, imag} */,
  {32'hbf808fae, 32'hc02cada2} /* (11, 2, 5) {real, imag} */,
  {32'h3ffd5a57, 32'hc1004f77} /* (11, 2, 4) {real, imag} */,
  {32'hc086cfcd, 32'h41009aa4} /* (11, 2, 3) {real, imag} */,
  {32'hc0a5ade9, 32'h408f00cc} /* (11, 2, 2) {real, imag} */,
  {32'h3f1368d2, 32'h40aead62} /* (11, 2, 1) {real, imag} */,
  {32'hbefa3045, 32'hc08800db} /* (11, 2, 0) {real, imag} */,
  {32'h40bf30e4, 32'hbfcd10d9} /* (11, 1, 15) {real, imag} */,
  {32'h40e9010e, 32'h3f724221} /* (11, 1, 14) {real, imag} */,
  {32'hbfcc3d28, 32'h409be3b5} /* (11, 1, 13) {real, imag} */,
  {32'h40f4e93c, 32'hc0d41d91} /* (11, 1, 12) {real, imag} */,
  {32'hbe71d7a3, 32'h40a4cef8} /* (11, 1, 11) {real, imag} */,
  {32'hbfc79da7, 32'hbfa37064} /* (11, 1, 10) {real, imag} */,
  {32'h3fb34c25, 32'hc01a3ff6} /* (11, 1, 9) {real, imag} */,
  {32'hbe9df1f0, 32'h3f8c4fd9} /* (11, 1, 8) {real, imag} */,
  {32'h4049016e, 32'h3f8ebf44} /* (11, 1, 7) {real, imag} */,
  {32'h414f3a39, 32'h40052813} /* (11, 1, 6) {real, imag} */,
  {32'hc1355d6f, 32'hc0c7b7ec} /* (11, 1, 5) {real, imag} */,
  {32'h3f37e4ae, 32'h3fbe09f6} /* (11, 1, 4) {real, imag} */,
  {32'h40526b80, 32'h3ff8ee83} /* (11, 1, 3) {real, imag} */,
  {32'hbf9b97af, 32'h3ef5ffc1} /* (11, 1, 2) {real, imag} */,
  {32'h404f2d57, 32'h40a56c76} /* (11, 1, 1) {real, imag} */,
  {32'h40642f82, 32'h40153326} /* (11, 1, 0) {real, imag} */,
  {32'h400ec935, 32'h3f7390a3} /* (11, 0, 15) {real, imag} */,
  {32'hc0adac02, 32'hbcf343c1} /* (11, 0, 14) {real, imag} */,
  {32'hc0580aa9, 32'h406727ab} /* (11, 0, 13) {real, imag} */,
  {32'h404cd604, 32'h4123382d} /* (11, 0, 12) {real, imag} */,
  {32'hc03f9a9e, 32'hc0975821} /* (11, 0, 11) {real, imag} */,
  {32'h406258f2, 32'h40899bc1} /* (11, 0, 10) {real, imag} */,
  {32'hc08deaec, 32'h3fbf8dda} /* (11, 0, 9) {real, imag} */,
  {32'hbfc396e1, 32'h3d263c72} /* (11, 0, 8) {real, imag} */,
  {32'h4021485b, 32'h40ad2af5} /* (11, 0, 7) {real, imag} */,
  {32'hbf2860fa, 32'h4088569a} /* (11, 0, 6) {real, imag} */,
  {32'hbfaa2128, 32'h41586b54} /* (11, 0, 5) {real, imag} */,
  {32'h40a10d96, 32'h3fff9b4f} /* (11, 0, 4) {real, imag} */,
  {32'hc0437b52, 32'hc031bb74} /* (11, 0, 3) {real, imag} */,
  {32'hc09b9369, 32'hc0110a1b} /* (11, 0, 2) {real, imag} */,
  {32'hc07395a1, 32'hc0a55cec} /* (11, 0, 1) {real, imag} */,
  {32'h410516d2, 32'h413222bc} /* (11, 0, 0) {real, imag} */,
  {32'h4020ac32, 32'h402bffcf} /* (10, 15, 15) {real, imag} */,
  {32'hc00fc011, 32'hbf62af50} /* (10, 15, 14) {real, imag} */,
  {32'h3fab0424, 32'hc149d60c} /* (10, 15, 13) {real, imag} */,
  {32'h3f31ed04, 32'h3fc3fcc3} /* (10, 15, 12) {real, imag} */,
  {32'h404732de, 32'hc0d80a35} /* (10, 15, 11) {real, imag} */,
  {32'h411cf580, 32'hc05cf0d8} /* (10, 15, 10) {real, imag} */,
  {32'hbf8a062c, 32'hbfd5d2d3} /* (10, 15, 9) {real, imag} */,
  {32'hc009c4a2, 32'h402f33dd} /* (10, 15, 8) {real, imag} */,
  {32'h4042edd5, 32'hc049572e} /* (10, 15, 7) {real, imag} */,
  {32'hc082a46b, 32'h40a6714e} /* (10, 15, 6) {real, imag} */,
  {32'hc0016147, 32'hc02718a7} /* (10, 15, 5) {real, imag} */,
  {32'h41178f86, 32'hc12d5c8a} /* (10, 15, 4) {real, imag} */,
  {32'hc0aebe51, 32'hc0ff6b9b} /* (10, 15, 3) {real, imag} */,
  {32'hc11f946e, 32'hbfa6ee4a} /* (10, 15, 2) {real, imag} */,
  {32'hc06a8b5d, 32'hc04afcf2} /* (10, 15, 1) {real, imag} */,
  {32'h411d7d8b, 32'h4020db05} /* (10, 15, 0) {real, imag} */,
  {32'hc17eef01, 32'hc0548105} /* (10, 14, 15) {real, imag} */,
  {32'hc0077d63, 32'hc010def7} /* (10, 14, 14) {real, imag} */,
  {32'h40c9a0a7, 32'h3fdfe6ea} /* (10, 14, 13) {real, imag} */,
  {32'hc088c6d3, 32'h4134f836} /* (10, 14, 12) {real, imag} */,
  {32'h40f170f1, 32'hc0e6ce79} /* (10, 14, 11) {real, imag} */,
  {32'hbf79f3c6, 32'h3fe6f805} /* (10, 14, 10) {real, imag} */,
  {32'h4092ef2c, 32'hc00e2791} /* (10, 14, 9) {real, imag} */,
  {32'h3fce58d7, 32'hc006b15c} /* (10, 14, 8) {real, imag} */,
  {32'hc008346d, 32'hbe7c28ca} /* (10, 14, 7) {real, imag} */,
  {32'h3ff591b9, 32'h404adb02} /* (10, 14, 6) {real, imag} */,
  {32'hc09fcbfb, 32'h3f3ef20b} /* (10, 14, 5) {real, imag} */,
  {32'h3f691606, 32'hc0cc3b25} /* (10, 14, 4) {real, imag} */,
  {32'h4070c678, 32'hbeabdb06} /* (10, 14, 3) {real, imag} */,
  {32'hc105fa01, 32'h3f90b79b} /* (10, 14, 2) {real, imag} */,
  {32'h40e4dd0d, 32'hc0b1d8a1} /* (10, 14, 1) {real, imag} */,
  {32'h4110ae5d, 32'hc0dafafe} /* (10, 14, 0) {real, imag} */,
  {32'hbf2300ed, 32'h409a6b0c} /* (10, 13, 15) {real, imag} */,
  {32'h3f10b93f, 32'hc0a5471f} /* (10, 13, 14) {real, imag} */,
  {32'hc0ba0199, 32'hc06b0e0e} /* (10, 13, 13) {real, imag} */,
  {32'h409b2498, 32'hc0521712} /* (10, 13, 12) {real, imag} */,
  {32'h3fc02dce, 32'hbfec1fb9} /* (10, 13, 11) {real, imag} */,
  {32'hc093c5b1, 32'h3e5760b1} /* (10, 13, 10) {real, imag} */,
  {32'h407188c1, 32'hc0503a8d} /* (10, 13, 9) {real, imag} */,
  {32'hbf41f644, 32'hc0179977} /* (10, 13, 8) {real, imag} */,
  {32'hbfa34486, 32'hc06de7ab} /* (10, 13, 7) {real, imag} */,
  {32'hbfe5dd5f, 32'hc020d6d4} /* (10, 13, 6) {real, imag} */,
  {32'h3f4f2d02, 32'h4026650d} /* (10, 13, 5) {real, imag} */,
  {32'h40a00933, 32'hc00015a9} /* (10, 13, 4) {real, imag} */,
  {32'h40415d2f, 32'hc10a73d3} /* (10, 13, 3) {real, imag} */,
  {32'hbe289dc3, 32'hbf575d38} /* (10, 13, 2) {real, imag} */,
  {32'hc04810f6, 32'h400d4d95} /* (10, 13, 1) {real, imag} */,
  {32'hbd23c333, 32'h40e95153} /* (10, 13, 0) {real, imag} */,
  {32'h40bec05e, 32'hbfd35f61} /* (10, 12, 15) {real, imag} */,
  {32'h40f4a8dd, 32'hc0e7248c} /* (10, 12, 14) {real, imag} */,
  {32'hc008fbb8, 32'h40634149} /* (10, 12, 13) {real, imag} */,
  {32'hc148a072, 32'h3f1fd9d8} /* (10, 12, 12) {real, imag} */,
  {32'h3fe201ab, 32'h3fd55aaa} /* (10, 12, 11) {real, imag} */,
  {32'h4090276d, 32'hc01d197d} /* (10, 12, 10) {real, imag} */,
  {32'hc081119e, 32'h4043de81} /* (10, 12, 9) {real, imag} */,
  {32'h3f7022d0, 32'h41269ce6} /* (10, 12, 8) {real, imag} */,
  {32'h3e780501, 32'h408e76f5} /* (10, 12, 7) {real, imag} */,
  {32'hc0eece7c, 32'hbfe3a78a} /* (10, 12, 6) {real, imag} */,
  {32'hc06236ec, 32'hbeb19665} /* (10, 12, 5) {real, imag} */,
  {32'h405ac727, 32'hbf2da4da} /* (10, 12, 4) {real, imag} */,
  {32'hbfe5b401, 32'hbf725c54} /* (10, 12, 3) {real, imag} */,
  {32'hc0e994a1, 32'hc0361171} /* (10, 12, 2) {real, imag} */,
  {32'h40d4f4d2, 32'h40d05cff} /* (10, 12, 1) {real, imag} */,
  {32'hc0900b90, 32'hc062129d} /* (10, 12, 0) {real, imag} */,
  {32'h40f6a19c, 32'hbe872390} /* (10, 11, 15) {real, imag} */,
  {32'hbf055506, 32'h412c5fae} /* (10, 11, 14) {real, imag} */,
  {32'h40fbb959, 32'h40add896} /* (10, 11, 13) {real, imag} */,
  {32'hc10480d6, 32'hc0195d59} /* (10, 11, 12) {real, imag} */,
  {32'h3e730f2f, 32'hc13d8962} /* (10, 11, 11) {real, imag} */,
  {32'hc0ea8c1b, 32'hc0969eb0} /* (10, 11, 10) {real, imag} */,
  {32'hc0eff9ff, 32'h41341868} /* (10, 11, 9) {real, imag} */,
  {32'hc07bf31f, 32'hc0844e97} /* (10, 11, 8) {real, imag} */,
  {32'hc0340a47, 32'h40822b20} /* (10, 11, 7) {real, imag} */,
  {32'h40426323, 32'hc015bad8} /* (10, 11, 6) {real, imag} */,
  {32'h3ff9bde9, 32'hbf72b9a5} /* (10, 11, 5) {real, imag} */,
  {32'hc037697d, 32'h410acf09} /* (10, 11, 4) {real, imag} */,
  {32'hbf60f8ec, 32'hc152a809} /* (10, 11, 3) {real, imag} */,
  {32'h3f16184d, 32'h40c11994} /* (10, 11, 2) {real, imag} */,
  {32'h3f072f72, 32'h3f14322f} /* (10, 11, 1) {real, imag} */,
  {32'h40299827, 32'hc0eb0c45} /* (10, 11, 0) {real, imag} */,
  {32'h404ffc42, 32'h404d87a2} /* (10, 10, 15) {real, imag} */,
  {32'h40dd7d5b, 32'h40c99a6b} /* (10, 10, 14) {real, imag} */,
  {32'hbe84ca8d, 32'hbf442bb0} /* (10, 10, 13) {real, imag} */,
  {32'hc0128c2b, 32'hc0ea59f5} /* (10, 10, 12) {real, imag} */,
  {32'h4064af94, 32'hbf16ee70} /* (10, 10, 11) {real, imag} */,
  {32'h41002cd9, 32'hc07b7514} /* (10, 10, 10) {real, imag} */,
  {32'hbf306a9f, 32'h403f020d} /* (10, 10, 9) {real, imag} */,
  {32'h3fe5bfd5, 32'hc035a36e} /* (10, 10, 8) {real, imag} */,
  {32'h40d249de, 32'hbfe5e92f} /* (10, 10, 7) {real, imag} */,
  {32'h40850aab, 32'h409ed226} /* (10, 10, 6) {real, imag} */,
  {32'hbf8351c8, 32'hc0df1d2a} /* (10, 10, 5) {real, imag} */,
  {32'h40bff674, 32'hc105d851} /* (10, 10, 4) {real, imag} */,
  {32'hc0454066, 32'h3fd93ff6} /* (10, 10, 3) {real, imag} */,
  {32'hc074a9d0, 32'hbfe1050d} /* (10, 10, 2) {real, imag} */,
  {32'hc089bdf5, 32'h40aa1d6d} /* (10, 10, 1) {real, imag} */,
  {32'hc1109b5c, 32'h404d597d} /* (10, 10, 0) {real, imag} */,
  {32'hc09e519e, 32'hbe133e13} /* (10, 9, 15) {real, imag} */,
  {32'hc09557a6, 32'hc0876579} /* (10, 9, 14) {real, imag} */,
  {32'hc0d21769, 32'h3fd09199} /* (10, 9, 13) {real, imag} */,
  {32'hc081f871, 32'hc00ccc1f} /* (10, 9, 12) {real, imag} */,
  {32'h402723fa, 32'h414d4e2d} /* (10, 9, 11) {real, imag} */,
  {32'h40785883, 32'hbfe9ab22} /* (10, 9, 10) {real, imag} */,
  {32'hbf7c5da0, 32'hc0964a06} /* (10, 9, 9) {real, imag} */,
  {32'h40f39702, 32'h40cc3dec} /* (10, 9, 8) {real, imag} */,
  {32'hc0ae1e76, 32'h405cac02} /* (10, 9, 7) {real, imag} */,
  {32'hc088b411, 32'hc0417572} /* (10, 9, 6) {real, imag} */,
  {32'h40448fcc, 32'hc0a6b9c4} /* (10, 9, 5) {real, imag} */,
  {32'h3e63f6d8, 32'h405bbc13} /* (10, 9, 4) {real, imag} */,
  {32'h410f00ba, 32'h413194f1} /* (10, 9, 3) {real, imag} */,
  {32'hbf40858b, 32'h3f70eb2a} /* (10, 9, 2) {real, imag} */,
  {32'hbee5cae5, 32'h3f871604} /* (10, 9, 1) {real, imag} */,
  {32'h40b7ab4d, 32'h3fd99b01} /* (10, 9, 0) {real, imag} */,
  {32'h40b55f5f, 32'hbfb82a33} /* (10, 8, 15) {real, imag} */,
  {32'hc0516d77, 32'hc0c50c65} /* (10, 8, 14) {real, imag} */,
  {32'hc002f77a, 32'h40b5a370} /* (10, 8, 13) {real, imag} */,
  {32'h3fa3bfa7, 32'hc07d7899} /* (10, 8, 12) {real, imag} */,
  {32'hc0999cb0, 32'h40e0aa41} /* (10, 8, 11) {real, imag} */,
  {32'h410a590b, 32'hc05efde6} /* (10, 8, 10) {real, imag} */,
  {32'h4095afef, 32'hc00cf2c2} /* (10, 8, 9) {real, imag} */,
  {32'hbf4b2f46, 32'h4003acfa} /* (10, 8, 8) {real, imag} */,
  {32'h3d87c7b7, 32'hc07d4c80} /* (10, 8, 7) {real, imag} */,
  {32'h3ffefe22, 32'h408f5871} /* (10, 8, 6) {real, imag} */,
  {32'h40c680d8, 32'h3fe309a0} /* (10, 8, 5) {real, imag} */,
  {32'hbfbb8f20, 32'h4003cb26} /* (10, 8, 4) {real, imag} */,
  {32'h3d10eef0, 32'hbfed7a44} /* (10, 8, 3) {real, imag} */,
  {32'h3fc95f0c, 32'hbffe14bb} /* (10, 8, 2) {real, imag} */,
  {32'hc05963d9, 32'h3f11e4e1} /* (10, 8, 1) {real, imag} */,
  {32'h400fc950, 32'hc0535aa0} /* (10, 8, 0) {real, imag} */,
  {32'h3fc7c5f5, 32'hc0596035} /* (10, 7, 15) {real, imag} */,
  {32'hc05e8412, 32'h410603a7} /* (10, 7, 14) {real, imag} */,
  {32'h3e7556d0, 32'hbf6f89c9} /* (10, 7, 13) {real, imag} */,
  {32'h3ea47289, 32'hc1280341} /* (10, 7, 12) {real, imag} */,
  {32'hc056ee7b, 32'hc000250b} /* (10, 7, 11) {real, imag} */,
  {32'hbeb2ae6f, 32'hbec3dd7a} /* (10, 7, 10) {real, imag} */,
  {32'h3cdfba8c, 32'hbff481a3} /* (10, 7, 9) {real, imag} */,
  {32'h3f6e30fa, 32'h407bb9c0} /* (10, 7, 8) {real, imag} */,
  {32'hc0566b02, 32'hbfa5f9f7} /* (10, 7, 7) {real, imag} */,
  {32'h407fdc1b, 32'hc11d9d10} /* (10, 7, 6) {real, imag} */,
  {32'h4068ccf1, 32'h3f3b67e4} /* (10, 7, 5) {real, imag} */,
  {32'h4028de5f, 32'h403abb36} /* (10, 7, 4) {real, imag} */,
  {32'hc0dc43a2, 32'h4129a71f} /* (10, 7, 3) {real, imag} */,
  {32'h3f026290, 32'h3fc0263a} /* (10, 7, 2) {real, imag} */,
  {32'hc0a2efc5, 32'hbfd577f3} /* (10, 7, 1) {real, imag} */,
  {32'h4090f1bc, 32'hc03d83f0} /* (10, 7, 0) {real, imag} */,
  {32'hc0c576bb, 32'hbc68b3dd} /* (10, 6, 15) {real, imag} */,
  {32'hc0ac6f6d, 32'h402e0190} /* (10, 6, 14) {real, imag} */,
  {32'h4081e3a7, 32'h40c30b97} /* (10, 6, 13) {real, imag} */,
  {32'hbf6cc1da, 32'hc09d7f41} /* (10, 6, 12) {real, imag} */,
  {32'hc1490523, 32'hbfb7e5e6} /* (10, 6, 11) {real, imag} */,
  {32'h406ae90e, 32'hc10ad77e} /* (10, 6, 10) {real, imag} */,
  {32'h411cfeba, 32'hc0554832} /* (10, 6, 9) {real, imag} */,
  {32'hc0ca6727, 32'hc0963ef1} /* (10, 6, 8) {real, imag} */,
  {32'hc0a9a438, 32'h413cb3db} /* (10, 6, 7) {real, imag} */,
  {32'h4138093e, 32'hbf858ed5} /* (10, 6, 6) {real, imag} */,
  {32'hc0a688c8, 32'h3f4c4813} /* (10, 6, 5) {real, imag} */,
  {32'h418fb3aa, 32'h3efad31e} /* (10, 6, 4) {real, imag} */,
  {32'hc07e6d2f, 32'hc07cd2ba} /* (10, 6, 3) {real, imag} */,
  {32'hc11ef296, 32'h3fb89451} /* (10, 6, 2) {real, imag} */,
  {32'h40a7ed10, 32'hbe55eb90} /* (10, 6, 1) {real, imag} */,
  {32'hbf94544c, 32'h3fe2953b} /* (10, 6, 0) {real, imag} */,
  {32'hbf83fe8d, 32'h40b258f5} /* (10, 5, 15) {real, imag} */,
  {32'hbfa4d48c, 32'hc054525c} /* (10, 5, 14) {real, imag} */,
  {32'hc11d5bb4, 32'hbf87edd8} /* (10, 5, 13) {real, imag} */,
  {32'h402eb955, 32'h413d9594} /* (10, 5, 12) {real, imag} */,
  {32'hc03e5615, 32'hc09bd9e1} /* (10, 5, 11) {real, imag} */,
  {32'hc02c62ff, 32'hc1237358} /* (10, 5, 10) {real, imag} */,
  {32'h40992b93, 32'h4155a805} /* (10, 5, 9) {real, imag} */,
  {32'hc05f6828, 32'hc0a7b217} /* (10, 5, 8) {real, imag} */,
  {32'hc04e2ffe, 32'h40153634} /* (10, 5, 7) {real, imag} */,
  {32'hc0d88da6, 32'h407b8e30} /* (10, 5, 6) {real, imag} */,
  {32'h40b71305, 32'hc06a9ebb} /* (10, 5, 5) {real, imag} */,
  {32'hbfa13528, 32'hc08a2d4e} /* (10, 5, 4) {real, imag} */,
  {32'hc061a4fb, 32'hc0c5ba15} /* (10, 5, 3) {real, imag} */,
  {32'hc04092f2, 32'hbf27db32} /* (10, 5, 2) {real, imag} */,
  {32'h3f849b31, 32'hc03635f0} /* (10, 5, 1) {real, imag} */,
  {32'h40a18ba8, 32'hc085364f} /* (10, 5, 0) {real, imag} */,
  {32'hc12bb27a, 32'h4065bec6} /* (10, 4, 15) {real, imag} */,
  {32'h3f9918c2, 32'hc0ab5284} /* (10, 4, 14) {real, imag} */,
  {32'hc151a381, 32'h40c4c954} /* (10, 4, 13) {real, imag} */,
  {32'h40d49f8a, 32'h41071164} /* (10, 4, 12) {real, imag} */,
  {32'hbed51383, 32'h405c9194} /* (10, 4, 11) {real, imag} */,
  {32'h40436d01, 32'hbe471bac} /* (10, 4, 10) {real, imag} */,
  {32'hc0b65c60, 32'hc0b21c9b} /* (10, 4, 9) {real, imag} */,
  {32'h40c1f875, 32'h402350e3} /* (10, 4, 8) {real, imag} */,
  {32'h403036dd, 32'hc06bd83b} /* (10, 4, 7) {real, imag} */,
  {32'hc07a23f5, 32'h410c4d02} /* (10, 4, 6) {real, imag} */,
  {32'h40cf4d76, 32'hc153eecc} /* (10, 4, 5) {real, imag} */,
  {32'hbf004fa1, 32'h40e40fb4} /* (10, 4, 4) {real, imag} */,
  {32'hc0beaee5, 32'h4033aba1} /* (10, 4, 3) {real, imag} */,
  {32'h3f2c41f9, 32'hbe4f6db8} /* (10, 4, 2) {real, imag} */,
  {32'hbf5737f0, 32'h40b11624} /* (10, 4, 1) {real, imag} */,
  {32'h407e74bf, 32'hc0eed3c0} /* (10, 4, 0) {real, imag} */,
  {32'h40a96420, 32'h3f7dde2d} /* (10, 3, 15) {real, imag} */,
  {32'h40d96efc, 32'h40bde833} /* (10, 3, 14) {real, imag} */,
  {32'h40580cfe, 32'hc0468f54} /* (10, 3, 13) {real, imag} */,
  {32'hbf899a44, 32'h41206777} /* (10, 3, 12) {real, imag} */,
  {32'h3fac0524, 32'h400fb32f} /* (10, 3, 11) {real, imag} */,
  {32'h40396642, 32'h40ab6f82} /* (10, 3, 10) {real, imag} */,
  {32'hc084d83a, 32'hbfc63f90} /* (10, 3, 9) {real, imag} */,
  {32'h3e1ba08b, 32'hbf63510f} /* (10, 3, 8) {real, imag} */,
  {32'h3f8d924b, 32'hc0856e99} /* (10, 3, 7) {real, imag} */,
  {32'h4020db58, 32'h40393438} /* (10, 3, 6) {real, imag} */,
  {32'h41515cf5, 32'hbfd181b5} /* (10, 3, 5) {real, imag} */,
  {32'hc06c771f, 32'hc024c8d9} /* (10, 3, 4) {real, imag} */,
  {32'hc0392c66, 32'hc114ae3f} /* (10, 3, 3) {real, imag} */,
  {32'hc01a4dec, 32'hc05933f1} /* (10, 3, 2) {real, imag} */,
  {32'h40ff9bd4, 32'h40656826} /* (10, 3, 1) {real, imag} */,
  {32'hc0c8a0a6, 32'h40e48bbd} /* (10, 3, 0) {real, imag} */,
  {32'h40accc07, 32'hbfc97fd3} /* (10, 2, 15) {real, imag} */,
  {32'hbf44fd32, 32'hc002d7ba} /* (10, 2, 14) {real, imag} */,
  {32'h404f2e16, 32'h3e7716ff} /* (10, 2, 13) {real, imag} */,
  {32'h40bbaaf7, 32'h40ae9293} /* (10, 2, 12) {real, imag} */,
  {32'hc012e1cf, 32'hc0516074} /* (10, 2, 11) {real, imag} */,
  {32'hbfca91a9, 32'h40eeb14c} /* (10, 2, 10) {real, imag} */,
  {32'hc0ee1057, 32'h3ddbd59f} /* (10, 2, 9) {real, imag} */,
  {32'h40ee1498, 32'h400cb7cf} /* (10, 2, 8) {real, imag} */,
  {32'h4010b239, 32'hc079028a} /* (10, 2, 7) {real, imag} */,
  {32'hc0ae81c0, 32'hbeb76558} /* (10, 2, 6) {real, imag} */,
  {32'hc0e753a3, 32'hc01b48d1} /* (10, 2, 5) {real, imag} */,
  {32'h400c9b4e, 32'hc08ee483} /* (10, 2, 4) {real, imag} */,
  {32'hbecaf886, 32'h406613c5} /* (10, 2, 3) {real, imag} */,
  {32'hc02c631d, 32'h40f9dc37} /* (10, 2, 2) {real, imag} */,
  {32'hc02ba22b, 32'hc030439b} /* (10, 2, 1) {real, imag} */,
  {32'h3febfa15, 32'hc01fa633} /* (10, 2, 0) {real, imag} */,
  {32'h40ffdb88, 32'h3f6890cc} /* (10, 1, 15) {real, imag} */,
  {32'h3f384640, 32'hc111b0f2} /* (10, 1, 14) {real, imag} */,
  {32'h3e5cdbf5, 32'h4047d464} /* (10, 1, 13) {real, imag} */,
  {32'hc02ef38e, 32'h3fce023c} /* (10, 1, 12) {real, imag} */,
  {32'h3f921c0b, 32'hc001440e} /* (10, 1, 11) {real, imag} */,
  {32'h4051de29, 32'h3edc5013} /* (10, 1, 10) {real, imag} */,
  {32'h4152f439, 32'hbfad7fda} /* (10, 1, 9) {real, imag} */,
  {32'hbfa40643, 32'h40416a22} /* (10, 1, 8) {real, imag} */,
  {32'h403abe91, 32'h40bd5a66} /* (10, 1, 7) {real, imag} */,
  {32'hbf3c7541, 32'hbf1dd2d4} /* (10, 1, 6) {real, imag} */,
  {32'h3fdab7cf, 32'h403b250d} /* (10, 1, 5) {real, imag} */,
  {32'hc01fc859, 32'h3e3988ae} /* (10, 1, 4) {real, imag} */,
  {32'hc0bede06, 32'hc0cbf17a} /* (10, 1, 3) {real, imag} */,
  {32'h40e0a593, 32'hc0d6f6f8} /* (10, 1, 2) {real, imag} */,
  {32'hbfec3d3c, 32'h3fd49a6f} /* (10, 1, 1) {real, imag} */,
  {32'hc11b4135, 32'hc0a3b381} /* (10, 1, 0) {real, imag} */,
  {32'h3f5f6514, 32'h40264903} /* (10, 0, 15) {real, imag} */,
  {32'hc10c4f85, 32'h40bacf57} /* (10, 0, 14) {real, imag} */,
  {32'hc027a5c5, 32'hbf55525f} /* (10, 0, 13) {real, imag} */,
  {32'h40083a22, 32'hbfbfc246} /* (10, 0, 12) {real, imag} */,
  {32'hc0a6258d, 32'h3f33b50a} /* (10, 0, 11) {real, imag} */,
  {32'hc06862da, 32'hbfdf273b} /* (10, 0, 10) {real, imag} */,
  {32'hbff6f7fa, 32'hbf99c1b5} /* (10, 0, 9) {real, imag} */,
  {32'hc036a137, 32'h4011727e} /* (10, 0, 8) {real, imag} */,
  {32'hbeef7dc4, 32'hbfbed9ba} /* (10, 0, 7) {real, imag} */,
  {32'h40a1c530, 32'hbf3821c3} /* (10, 0, 6) {real, imag} */,
  {32'hc0725f66, 32'hbf9ab391} /* (10, 0, 5) {real, imag} */,
  {32'hc0b42b44, 32'h40ac0006} /* (10, 0, 4) {real, imag} */,
  {32'hc02ed998, 32'h40aab37c} /* (10, 0, 3) {real, imag} */,
  {32'h411ddfd9, 32'hc00d9f7b} /* (10, 0, 2) {real, imag} */,
  {32'h40483413, 32'h409376e5} /* (10, 0, 1) {real, imag} */,
  {32'h3f3dcb7f, 32'hc00488f1} /* (10, 0, 0) {real, imag} */,
  {32'h4101135a, 32'hc02d3f08} /* (9, 15, 15) {real, imag} */,
  {32'h3eddcd7e, 32'hbe59444c} /* (9, 15, 14) {real, imag} */,
  {32'hc0bd4cfe, 32'h401484ac} /* (9, 15, 13) {real, imag} */,
  {32'h3f58ba4a, 32'hc0e7cca3} /* (9, 15, 12) {real, imag} */,
  {32'h410549bd, 32'hc10445d9} /* (9, 15, 11) {real, imag} */,
  {32'hc0f92ba0, 32'hbfc7b229} /* (9, 15, 10) {real, imag} */,
  {32'h3ef7b049, 32'hc0888078} /* (9, 15, 9) {real, imag} */,
  {32'h400dabdb, 32'hc056e7f8} /* (9, 15, 8) {real, imag} */,
  {32'hbf380436, 32'hc048e755} /* (9, 15, 7) {real, imag} */,
  {32'h3f9288df, 32'hbfacdaab} /* (9, 15, 6) {real, imag} */,
  {32'hc0c79ce1, 32'h3f8f1163} /* (9, 15, 5) {real, imag} */,
  {32'hc02588d0, 32'h403669a9} /* (9, 15, 4) {real, imag} */,
  {32'hc09e2b3b, 32'hbfc06208} /* (9, 15, 3) {real, imag} */,
  {32'h3f13acf4, 32'hbf21e3fa} /* (9, 15, 2) {real, imag} */,
  {32'hbf882ad3, 32'h3f9d32bc} /* (9, 15, 1) {real, imag} */,
  {32'hbef1e514, 32'h40727ba6} /* (9, 15, 0) {real, imag} */,
  {32'h402e2766, 32'h408dbc34} /* (9, 14, 15) {real, imag} */,
  {32'hc0da8731, 32'hc060b4c3} /* (9, 14, 14) {real, imag} */,
  {32'hbfc3c26c, 32'hbd3a9327} /* (9, 14, 13) {real, imag} */,
  {32'h3f465ddb, 32'h40069e1d} /* (9, 14, 12) {real, imag} */,
  {32'hc0eaf60b, 32'h40267e63} /* (9, 14, 11) {real, imag} */,
  {32'h4102966c, 32'h408a0951} /* (9, 14, 10) {real, imag} */,
  {32'h4002d012, 32'hbf5288fb} /* (9, 14, 9) {real, imag} */,
  {32'h3fcf9302, 32'h4040d707} /* (9, 14, 8) {real, imag} */,
  {32'hc031276f, 32'hc056e18e} /* (9, 14, 7) {real, imag} */,
  {32'h401a59a1, 32'h3e76545a} /* (9, 14, 6) {real, imag} */,
  {32'h40d5e4fe, 32'h3f27560d} /* (9, 14, 5) {real, imag} */,
  {32'hbf14a44b, 32'h409fae46} /* (9, 14, 4) {real, imag} */,
  {32'h40365d31, 32'h4047a3d7} /* (9, 14, 3) {real, imag} */,
  {32'h3fb5cd7a, 32'hbe4da5a6} /* (9, 14, 2) {real, imag} */,
  {32'hbf6219d4, 32'hc029cbf7} /* (9, 14, 1) {real, imag} */,
  {32'hbff960a2, 32'hbf9c6d46} /* (9, 14, 0) {real, imag} */,
  {32'h404f4009, 32'h3fbbb82f} /* (9, 13, 15) {real, imag} */,
  {32'hc00565bd, 32'h3f0efb89} /* (9, 13, 14) {real, imag} */,
  {32'h3f6f5d0d, 32'h4021b7ea} /* (9, 13, 13) {real, imag} */,
  {32'h40b5fc94, 32'h3fa197f4} /* (9, 13, 12) {real, imag} */,
  {32'hbf121573, 32'h3f764ee5} /* (9, 13, 11) {real, imag} */,
  {32'hc0a94ba7, 32'hbf859152} /* (9, 13, 10) {real, imag} */,
  {32'h3f9b0c86, 32'hbff7cf3d} /* (9, 13, 9) {real, imag} */,
  {32'h3f660fda, 32'h3f9c9939} /* (9, 13, 8) {real, imag} */,
  {32'h3fb1b512, 32'h40c913a7} /* (9, 13, 7) {real, imag} */,
  {32'hc10026ba, 32'hc01a537b} /* (9, 13, 6) {real, imag} */,
  {32'h3f2d1d8e, 32'h3f296441} /* (9, 13, 5) {real, imag} */,
  {32'hc00b431e, 32'h40e361e0} /* (9, 13, 4) {real, imag} */,
  {32'h40556148, 32'hc0909178} /* (9, 13, 3) {real, imag} */,
  {32'h407136b8, 32'hc071c8c8} /* (9, 13, 2) {real, imag} */,
  {32'hc0e6906d, 32'h3f6c0388} /* (9, 13, 1) {real, imag} */,
  {32'hc06117ce, 32'hc09db10e} /* (9, 13, 0) {real, imag} */,
  {32'hc064d1a7, 32'h410927ca} /* (9, 12, 15) {real, imag} */,
  {32'h3fcb6b66, 32'h4053fbf1} /* (9, 12, 14) {real, imag} */,
  {32'hc0366f7c, 32'hc0b62040} /* (9, 12, 13) {real, imag} */,
  {32'h3fddd06f, 32'hc0ad5887} /* (9, 12, 12) {real, imag} */,
  {32'hc0aa246d, 32'h40821627} /* (9, 12, 11) {real, imag} */,
  {32'hc09b4d4a, 32'h3df4a12e} /* (9, 12, 10) {real, imag} */,
  {32'hbff7e7ea, 32'h3f79634b} /* (9, 12, 9) {real, imag} */,
  {32'h400d774e, 32'h4040dd61} /* (9, 12, 8) {real, imag} */,
  {32'hbd47589b, 32'h3fd07b6b} /* (9, 12, 7) {real, imag} */,
  {32'h4046be6a, 32'h3f61f04c} /* (9, 12, 6) {real, imag} */,
  {32'h3fdb7c48, 32'h409a3d47} /* (9, 12, 5) {real, imag} */,
  {32'hbfaaf86b, 32'h4006c8ba} /* (9, 12, 4) {real, imag} */,
  {32'h3fccaddf, 32'hc00bdef9} /* (9, 12, 3) {real, imag} */,
  {32'h3fca0afb, 32'h4057323f} /* (9, 12, 2) {real, imag} */,
  {32'hc1214886, 32'hc02e1db0} /* (9, 12, 1) {real, imag} */,
  {32'h400cfbb2, 32'h3f3e0589} /* (9, 12, 0) {real, imag} */,
  {32'h40bb7f30, 32'hbfbe18ad} /* (9, 11, 15) {real, imag} */,
  {32'hbf659556, 32'hc097dec0} /* (9, 11, 14) {real, imag} */,
  {32'h3fb04b02, 32'h40997073} /* (9, 11, 13) {real, imag} */,
  {32'hbf66764b, 32'h3f001319} /* (9, 11, 12) {real, imag} */,
  {32'h4088b8be, 32'hc065dcd4} /* (9, 11, 11) {real, imag} */,
  {32'hbfca932a, 32'h40886d11} /* (9, 11, 10) {real, imag} */,
  {32'h4103e0a5, 32'hc08a81c9} /* (9, 11, 9) {real, imag} */,
  {32'hbffc1900, 32'hc009f87e} /* (9, 11, 8) {real, imag} */,
  {32'h4027729f, 32'hc003a442} /* (9, 11, 7) {real, imag} */,
  {32'h3fb9ea64, 32'hc064b9bb} /* (9, 11, 6) {real, imag} */,
  {32'h40ca91f5, 32'h402dd03a} /* (9, 11, 5) {real, imag} */,
  {32'h40392297, 32'hc10b83f9} /* (9, 11, 4) {real, imag} */,
  {32'hc0d316eb, 32'h40a78cae} /* (9, 11, 3) {real, imag} */,
  {32'hbf9ab1ce, 32'h406fa800} /* (9, 11, 2) {real, imag} */,
  {32'h3f88ef14, 32'h405ccca0} /* (9, 11, 1) {real, imag} */,
  {32'hc10c8167, 32'h3ffb126a} /* (9, 11, 0) {real, imag} */,
  {32'h401d07dd, 32'h40a2cd54} /* (9, 10, 15) {real, imag} */,
  {32'h4066926c, 32'h404b1f23} /* (9, 10, 14) {real, imag} */,
  {32'hc0d18296, 32'h3f0857f7} /* (9, 10, 13) {real, imag} */,
  {32'hc08f5de4, 32'h40c39517} /* (9, 10, 12) {real, imag} */,
  {32'h402cdd66, 32'hbe648838} /* (9, 10, 11) {real, imag} */,
  {32'hc119ef67, 32'hbfc3c523} /* (9, 10, 10) {real, imag} */,
  {32'hc01373c5, 32'hbfe4f24d} /* (9, 10, 9) {real, imag} */,
  {32'h3f5a6bed, 32'hc0ab2a5b} /* (9, 10, 8) {real, imag} */,
  {32'h3f9cbdc1, 32'h3ec7bb41} /* (9, 10, 7) {real, imag} */,
  {32'h4170e741, 32'h41461b5e} /* (9, 10, 6) {real, imag} */,
  {32'h404b76ce, 32'h40062f78} /* (9, 10, 5) {real, imag} */,
  {32'hc104bf65, 32'h3e65a044} /* (9, 10, 4) {real, imag} */,
  {32'hc0dc0c4b, 32'h409efbe9} /* (9, 10, 3) {real, imag} */,
  {32'h40db68fa, 32'hc0a4f364} /* (9, 10, 2) {real, imag} */,
  {32'hbf7ab9d1, 32'hbfcae520} /* (9, 10, 1) {real, imag} */,
  {32'h3fa10601, 32'h40f3390f} /* (9, 10, 0) {real, imag} */,
  {32'hbfd22499, 32'h402f02c8} /* (9, 9, 15) {real, imag} */,
  {32'hc01b1346, 32'h4102704e} /* (9, 9, 14) {real, imag} */,
  {32'h40fb32be, 32'hbdbdb0e5} /* (9, 9, 13) {real, imag} */,
  {32'h40807d27, 32'hc082ed68} /* (9, 9, 12) {real, imag} */,
  {32'hc1127c9b, 32'hc02c4ca0} /* (9, 9, 11) {real, imag} */,
  {32'h411ce0f4, 32'hc0991c91} /* (9, 9, 10) {real, imag} */,
  {32'hc088da08, 32'h4100dad1} /* (9, 9, 9) {real, imag} */,
  {32'hbf8cce15, 32'hc0032300} /* (9, 9, 8) {real, imag} */,
  {32'hc095e6f6, 32'h4112d930} /* (9, 9, 7) {real, imag} */,
  {32'h406f8a8b, 32'h404a6ca8} /* (9, 9, 6) {real, imag} */,
  {32'hbfcdce51, 32'h4112e270} /* (9, 9, 5) {real, imag} */,
  {32'h40d9627c, 32'hc0b98589} /* (9, 9, 4) {real, imag} */,
  {32'h3fac6fd1, 32'h3fc86ac4} /* (9, 9, 3) {real, imag} */,
  {32'hc0f1b0fe, 32'hc0d09af3} /* (9, 9, 2) {real, imag} */,
  {32'hc0c1be00, 32'hbe26e2f0} /* (9, 9, 1) {real, imag} */,
  {32'h408a9d03, 32'hc03ad60c} /* (9, 9, 0) {real, imag} */,
  {32'hbf3c14ef, 32'hbf353ec4} /* (9, 8, 15) {real, imag} */,
  {32'h406f2d9a, 32'h3fbc346c} /* (9, 8, 14) {real, imag} */,
  {32'h403c9130, 32'hc093a4dc} /* (9, 8, 13) {real, imag} */,
  {32'h3fde5948, 32'h40c326d8} /* (9, 8, 12) {real, imag} */,
  {32'hc096fdb0, 32'hc08e2f59} /* (9, 8, 11) {real, imag} */,
  {32'h3e396329, 32'hbf48f3aa} /* (9, 8, 10) {real, imag} */,
  {32'h3f25c345, 32'h409dd412} /* (9, 8, 9) {real, imag} */,
  {32'hbe553ef0, 32'h40423d07} /* (9, 8, 8) {real, imag} */,
  {32'hbfb16f8a, 32'hc053b18c} /* (9, 8, 7) {real, imag} */,
  {32'hc0b764ab, 32'h3f4ff82e} /* (9, 8, 6) {real, imag} */,
  {32'h40aa9f72, 32'hc067d252} /* (9, 8, 5) {real, imag} */,
  {32'h404feba2, 32'h40b1936e} /* (9, 8, 4) {real, imag} */,
  {32'hbf2781f5, 32'hc0687f5c} /* (9, 8, 3) {real, imag} */,
  {32'h4000299b, 32'hc001eaae} /* (9, 8, 2) {real, imag} */,
  {32'h40b57c67, 32'h3fade9d0} /* (9, 8, 1) {real, imag} */,
  {32'h3fc8dbe6, 32'h3fdac877} /* (9, 8, 0) {real, imag} */,
  {32'h40c45ed4, 32'h401536a8} /* (9, 7, 15) {real, imag} */,
  {32'h40ff0c7e, 32'hbe8a28fc} /* (9, 7, 14) {real, imag} */,
  {32'h3f51652e, 32'h3ffbbceb} /* (9, 7, 13) {real, imag} */,
  {32'hc1170ca8, 32'h3f18071b} /* (9, 7, 12) {real, imag} */,
  {32'hc01e3155, 32'hc024a23e} /* (9, 7, 11) {real, imag} */,
  {32'hbe5fcfb7, 32'hc0256498} /* (9, 7, 10) {real, imag} */,
  {32'hbfac25dd, 32'h3f4bc95f} /* (9, 7, 9) {real, imag} */,
  {32'h3f0c9a88, 32'hbfd318f4} /* (9, 7, 8) {real, imag} */,
  {32'hc0b6a59b, 32'hc07df880} /* (9, 7, 7) {real, imag} */,
  {32'h3fe3ad74, 32'hbf0baeb4} /* (9, 7, 6) {real, imag} */,
  {32'hc0801c4a, 32'hbf238cf2} /* (9, 7, 5) {real, imag} */,
  {32'hc0383acc, 32'hbf13d7b8} /* (9, 7, 4) {real, imag} */,
  {32'h3fb44909, 32'hc069160e} /* (9, 7, 3) {real, imag} */,
  {32'h401ef6ba, 32'hbfb7ce6c} /* (9, 7, 2) {real, imag} */,
  {32'h4008f173, 32'h4083a825} /* (9, 7, 1) {real, imag} */,
  {32'hc05d2f7b, 32'hbfb7b71b} /* (9, 7, 0) {real, imag} */,
  {32'h40ba3b39, 32'hbfff7e5e} /* (9, 6, 15) {real, imag} */,
  {32'hbfc65ed4, 32'h408d077d} /* (9, 6, 14) {real, imag} */,
  {32'h40626405, 32'h3f2d3159} /* (9, 6, 13) {real, imag} */,
  {32'h3f8df11c, 32'h3f78bccc} /* (9, 6, 12) {real, imag} */,
  {32'hc0ad6944, 32'h4031a6d8} /* (9, 6, 11) {real, imag} */,
  {32'hc0dab354, 32'hbf2b0e26} /* (9, 6, 10) {real, imag} */,
  {32'h403e00fb, 32'hc0a4765b} /* (9, 6, 9) {real, imag} */,
  {32'h408ee152, 32'h4081fe62} /* (9, 6, 8) {real, imag} */,
  {32'h3eb237f6, 32'hc0f78634} /* (9, 6, 7) {real, imag} */,
  {32'h40adf51c, 32'hc0c88a18} /* (9, 6, 6) {real, imag} */,
  {32'h3f91dccc, 32'hc0f3891b} /* (9, 6, 5) {real, imag} */,
  {32'h3fd35bf1, 32'h40db67f2} /* (9, 6, 4) {real, imag} */,
  {32'hc01fbc23, 32'hc0cd754e} /* (9, 6, 3) {real, imag} */,
  {32'h40249209, 32'hc08c5564} /* (9, 6, 2) {real, imag} */,
  {32'h3f951478, 32'hc050caea} /* (9, 6, 1) {real, imag} */,
  {32'h4015ca50, 32'h40cf4cc9} /* (9, 6, 0) {real, imag} */,
  {32'hc0863532, 32'h40a33db0} /* (9, 5, 15) {real, imag} */,
  {32'h3f79056e, 32'h3f3f503f} /* (9, 5, 14) {real, imag} */,
  {32'hc07b15af, 32'h408b18dd} /* (9, 5, 13) {real, imag} */,
  {32'h3c826fa2, 32'h3f454c96} /* (9, 5, 12) {real, imag} */,
  {32'hc09eb404, 32'hc079ebf6} /* (9, 5, 11) {real, imag} */,
  {32'h3f2599a1, 32'hbd4d6cac} /* (9, 5, 10) {real, imag} */,
  {32'hc0d5651b, 32'hc123e9ce} /* (9, 5, 9) {real, imag} */,
  {32'hc0094ab0, 32'hbfee7737} /* (9, 5, 8) {real, imag} */,
  {32'h404a3936, 32'hbf0df615} /* (9, 5, 7) {real, imag} */,
  {32'h404e05ec, 32'h3d4105e3} /* (9, 5, 6) {real, imag} */,
  {32'h3f70cccb, 32'hbda8ab71} /* (9, 5, 5) {real, imag} */,
  {32'h4110620c, 32'hc006a244} /* (9, 5, 4) {real, imag} */,
  {32'hbf9baa8e, 32'hbe06d77f} /* (9, 5, 3) {real, imag} */,
  {32'hbf06a267, 32'hc0ca6647} /* (9, 5, 2) {real, imag} */,
  {32'hc10a6c59, 32'h412807d9} /* (9, 5, 1) {real, imag} */,
  {32'hbcdb2dc5, 32'h401812fd} /* (9, 5, 0) {real, imag} */,
  {32'h40621147, 32'h409bc352} /* (9, 4, 15) {real, imag} */,
  {32'h3fbf70d1, 32'h4051ca37} /* (9, 4, 14) {real, imag} */,
  {32'hc05b5625, 32'h3f9fcd11} /* (9, 4, 13) {real, imag} */,
  {32'h402e8a36, 32'hc0ec3f6e} /* (9, 4, 12) {real, imag} */,
  {32'h405bdf03, 32'hc0cb59e8} /* (9, 4, 11) {real, imag} */,
  {32'h40a837c9, 32'h4102c6a8} /* (9, 4, 10) {real, imag} */,
  {32'h403e1ea5, 32'h3e686c91} /* (9, 4, 9) {real, imag} */,
  {32'h4004b0b9, 32'hbfe09c12} /* (9, 4, 8) {real, imag} */,
  {32'h402f8da6, 32'h3f879f06} /* (9, 4, 7) {real, imag} */,
  {32'h3f4b6d42, 32'hc0117889} /* (9, 4, 6) {real, imag} */,
  {32'hbf8e2248, 32'h400deed5} /* (9, 4, 5) {real, imag} */,
  {32'hbf014628, 32'h401e2d7d} /* (9, 4, 4) {real, imag} */,
  {32'h40f45f2a, 32'hc08c387b} /* (9, 4, 3) {real, imag} */,
  {32'hc05df299, 32'hc0be1c8c} /* (9, 4, 2) {real, imag} */,
  {32'h40fa4326, 32'h4102328a} /* (9, 4, 1) {real, imag} */,
  {32'hbf3406e9, 32'hbfb589ac} /* (9, 4, 0) {real, imag} */,
  {32'hc083ecff, 32'h3e84a54c} /* (9, 3, 15) {real, imag} */,
  {32'h3e819bd1, 32'hbfb4f295} /* (9, 3, 14) {real, imag} */,
  {32'hc0263166, 32'h3f889fb3} /* (9, 3, 13) {real, imag} */,
  {32'h407e6017, 32'hbde3f9fd} /* (9, 3, 12) {real, imag} */,
  {32'h40d530c9, 32'hc09271b1} /* (9, 3, 11) {real, imag} */,
  {32'hc0052e4b, 32'h3fcdc611} /* (9, 3, 10) {real, imag} */,
  {32'hbfbff146, 32'h402b41a0} /* (9, 3, 9) {real, imag} */,
  {32'h40544907, 32'hbf68561a} /* (9, 3, 8) {real, imag} */,
  {32'hbf5a099d, 32'h40d1bfe4} /* (9, 3, 7) {real, imag} */,
  {32'h3fa36114, 32'h4040bbc5} /* (9, 3, 6) {real, imag} */,
  {32'hbff51f6d, 32'hc0250227} /* (9, 3, 5) {real, imag} */,
  {32'hbff0b52f, 32'h40bd7452} /* (9, 3, 4) {real, imag} */,
  {32'h3f884222, 32'h3fa89575} /* (9, 3, 3) {real, imag} */,
  {32'h3f89d2ae, 32'hc0faa1b3} /* (9, 3, 2) {real, imag} */,
  {32'h3f5f6c16, 32'hbf8b9115} /* (9, 3, 1) {real, imag} */,
  {32'hc03c433f, 32'hc05c7952} /* (9, 3, 0) {real, imag} */,
  {32'hc04bfd4d, 32'hc07faa7c} /* (9, 2, 15) {real, imag} */,
  {32'hc02f3545, 32'h41081825} /* (9, 2, 14) {real, imag} */,
  {32'hc02ef342, 32'h3ffb1fee} /* (9, 2, 13) {real, imag} */,
  {32'hc0d7f14c, 32'hbe84780c} /* (9, 2, 12) {real, imag} */,
  {32'h4105e3c5, 32'hc05cec75} /* (9, 2, 11) {real, imag} */,
  {32'h3e3706ab, 32'h3fbdf71b} /* (9, 2, 10) {real, imag} */,
  {32'h4031c1fa, 32'hc0c1e573} /* (9, 2, 9) {real, imag} */,
  {32'h408cf9a3, 32'h3f466d81} /* (9, 2, 8) {real, imag} */,
  {32'hbfe7b955, 32'hc0465ca2} /* (9, 2, 7) {real, imag} */,
  {32'hbf94f29d, 32'h3eb76a21} /* (9, 2, 6) {real, imag} */,
  {32'hbfb498f6, 32'h406d93c1} /* (9, 2, 5) {real, imag} */,
  {32'h40060871, 32'h40f46aea} /* (9, 2, 4) {real, imag} */,
  {32'hbca2d274, 32'hc0a81e70} /* (9, 2, 3) {real, imag} */,
  {32'h4091bbf5, 32'hbfc349b1} /* (9, 2, 2) {real, imag} */,
  {32'hc01383b8, 32'hc0aca95d} /* (9, 2, 1) {real, imag} */,
  {32'h4040cf01, 32'h400772bc} /* (9, 2, 0) {real, imag} */,
  {32'hc09bde59, 32'h40b342c7} /* (9, 1, 15) {real, imag} */,
  {32'hbf51de21, 32'hc0f094ee} /* (9, 1, 14) {real, imag} */,
  {32'hc059a2c0, 32'hbeddff66} /* (9, 1, 13) {real, imag} */,
  {32'h40712001, 32'hc041ef3d} /* (9, 1, 12) {real, imag} */,
  {32'hbf2b8a0b, 32'h4013dc1e} /* (9, 1, 11) {real, imag} */,
  {32'hbd68bbc7, 32'hc019abe9} /* (9, 1, 10) {real, imag} */,
  {32'hbf2916ec, 32'h411fa465} /* (9, 1, 9) {real, imag} */,
  {32'h3e85dfd6, 32'h4011e83d} /* (9, 1, 8) {real, imag} */,
  {32'hbf1955e6, 32'hbf0a22fd} /* (9, 1, 7) {real, imag} */,
  {32'hc08ad8ac, 32'h40e9c2e5} /* (9, 1, 6) {real, imag} */,
  {32'h3fe905a8, 32'hc10772e0} /* (9, 1, 5) {real, imag} */,
  {32'hbf104e75, 32'hc0196062} /* (9, 1, 4) {real, imag} */,
  {32'h410cd867, 32'h3e8c5e08} /* (9, 1, 3) {real, imag} */,
  {32'hc0985f6e, 32'h4011b739} /* (9, 1, 2) {real, imag} */,
  {32'h40ca9fb8, 32'h40675333} /* (9, 1, 1) {real, imag} */,
  {32'h3f31fe42, 32'h4008de34} /* (9, 1, 0) {real, imag} */,
  {32'h40a86f65, 32'hc04e0e48} /* (9, 0, 15) {real, imag} */,
  {32'hc069b9b0, 32'hc080708b} /* (9, 0, 14) {real, imag} */,
  {32'h40e4bde7, 32'hbce995a5} /* (9, 0, 13) {real, imag} */,
  {32'hc0085af5, 32'h3ec3269f} /* (9, 0, 12) {real, imag} */,
  {32'hc0c6ec1c, 32'h3f888e05} /* (9, 0, 11) {real, imag} */,
  {32'h3fe4ff35, 32'h411b2b0d} /* (9, 0, 10) {real, imag} */,
  {32'h40b0aeed, 32'hbf9446f0} /* (9, 0, 9) {real, imag} */,
  {32'hc0d0ebdd, 32'h408ef88b} /* (9, 0, 8) {real, imag} */,
  {32'h4016428c, 32'hbf512c4d} /* (9, 0, 7) {real, imag} */,
  {32'hbe1642db, 32'h3fc83b9e} /* (9, 0, 6) {real, imag} */,
  {32'h3e936454, 32'hc0c84235} /* (9, 0, 5) {real, imag} */,
  {32'hbe7566c1, 32'hc00f9993} /* (9, 0, 4) {real, imag} */,
  {32'hbfd7eca2, 32'h40d4cf1d} /* (9, 0, 3) {real, imag} */,
  {32'h40148df2, 32'h3e8a5b58} /* (9, 0, 2) {real, imag} */,
  {32'hc0603ac3, 32'hc09351de} /* (9, 0, 1) {real, imag} */,
  {32'h3faf7242, 32'hc0bcc546} /* (9, 0, 0) {real, imag} */,
  {32'h3f1a286a, 32'hbde9f465} /* (8, 15, 15) {real, imag} */,
  {32'hc08c85a4, 32'hbf30e2d8} /* (8, 15, 14) {real, imag} */,
  {32'h3fc3adbd, 32'h3d206b88} /* (8, 15, 13) {real, imag} */,
  {32'hc08d7f3d, 32'h3d85d151} /* (8, 15, 12) {real, imag} */,
  {32'h3f9ec775, 32'hc02b1c06} /* (8, 15, 11) {real, imag} */,
  {32'hc0a676b0, 32'hbfecc20a} /* (8, 15, 10) {real, imag} */,
  {32'h402f5752, 32'h40553b9a} /* (8, 15, 9) {real, imag} */,
  {32'hbf3cc9c4, 32'h40038b6f} /* (8, 15, 8) {real, imag} */,
  {32'hc02c6cc5, 32'hbf02def3} /* (8, 15, 7) {real, imag} */,
  {32'hc029219a, 32'hbe799fa7} /* (8, 15, 6) {real, imag} */,
  {32'h403e3003, 32'h3fc41db7} /* (8, 15, 5) {real, imag} */,
  {32'h3f9783da, 32'hbf23e785} /* (8, 15, 4) {real, imag} */,
  {32'hbf9bdf2f, 32'h406898ba} /* (8, 15, 3) {real, imag} */,
  {32'h3eace800, 32'hc0799a92} /* (8, 15, 2) {real, imag} */,
  {32'hc0084728, 32'hc097efb8} /* (8, 15, 1) {real, imag} */,
  {32'hbf48c257, 32'h3f58cac9} /* (8, 15, 0) {real, imag} */,
  {32'hbfb09032, 32'hc0fb55ca} /* (8, 14, 15) {real, imag} */,
  {32'hbf2e8fbc, 32'h40a7b849} /* (8, 14, 14) {real, imag} */,
  {32'hc0218250, 32'hbfca07ff} /* (8, 14, 13) {real, imag} */,
  {32'hbf8a3178, 32'hc0926569} /* (8, 14, 12) {real, imag} */,
  {32'h3f773374, 32'h40b2affa} /* (8, 14, 11) {real, imag} */,
  {32'h3f69efff, 32'hc016d2b0} /* (8, 14, 10) {real, imag} */,
  {32'h3e2bb16f, 32'hbf4c93f2} /* (8, 14, 9) {real, imag} */,
  {32'hbf55d3f1, 32'h4091adcd} /* (8, 14, 8) {real, imag} */,
  {32'h40b1b11e, 32'h409f4a87} /* (8, 14, 7) {real, imag} */,
  {32'h4061a1ae, 32'hbe9a121d} /* (8, 14, 6) {real, imag} */,
  {32'hbf199ec8, 32'h40d4c219} /* (8, 14, 5) {real, imag} */,
  {32'h40917d64, 32'h40632195} /* (8, 14, 4) {real, imag} */,
  {32'hc009a3f9, 32'hbfb748ed} /* (8, 14, 3) {real, imag} */,
  {32'hbe3d3be1, 32'h3fb3bcc2} /* (8, 14, 2) {real, imag} */,
  {32'h3beb754f, 32'hbe4fabe1} /* (8, 14, 1) {real, imag} */,
  {32'hbf4b1ed6, 32'h404de68b} /* (8, 14, 0) {real, imag} */,
  {32'hc08c180f, 32'h3f926af5} /* (8, 13, 15) {real, imag} */,
  {32'hbf5ba29d, 32'hbefc837d} /* (8, 13, 14) {real, imag} */,
  {32'h3fc4e28f, 32'hc0308128} /* (8, 13, 13) {real, imag} */,
  {32'h3fe9521d, 32'h40308037} /* (8, 13, 12) {real, imag} */,
  {32'hc0af6895, 32'h3f4aea00} /* (8, 13, 11) {real, imag} */,
  {32'h3f7c57c5, 32'h409bba52} /* (8, 13, 10) {real, imag} */,
  {32'h409ac016, 32'h40afa951} /* (8, 13, 9) {real, imag} */,
  {32'hc01bb076, 32'hc02e963c} /* (8, 13, 8) {real, imag} */,
  {32'h3f7b63da, 32'h4079b464} /* (8, 13, 7) {real, imag} */,
  {32'h4063513c, 32'hc09efbf2} /* (8, 13, 6) {real, imag} */,
  {32'hbfdc7f5f, 32'h4087ef1f} /* (8, 13, 5) {real, imag} */,
  {32'h3ff5adc1, 32'hc0497148} /* (8, 13, 4) {real, imag} */,
  {32'hc0b8e7f5, 32'h3fcf5bfa} /* (8, 13, 3) {real, imag} */,
  {32'hbe217bbc, 32'h3fd89068} /* (8, 13, 2) {real, imag} */,
  {32'h3f94481c, 32'hc0786f7f} /* (8, 13, 1) {real, imag} */,
  {32'hc012ca11, 32'h3f2030b6} /* (8, 13, 0) {real, imag} */,
  {32'hc0786613, 32'hc033fe43} /* (8, 12, 15) {real, imag} */,
  {32'h3f01b52f, 32'hc01b4fc4} /* (8, 12, 14) {real, imag} */,
  {32'hbf57df62, 32'h409c2da4} /* (8, 12, 13) {real, imag} */,
  {32'h3f6e01f1, 32'h407978b7} /* (8, 12, 12) {real, imag} */,
  {32'h3fd6631c, 32'h3e6391bc} /* (8, 12, 11) {real, imag} */,
  {32'hbf53fc1b, 32'hc01a11a0} /* (8, 12, 10) {real, imag} */,
  {32'h3e08f9c4, 32'h40364a41} /* (8, 12, 9) {real, imag} */,
  {32'hc0aa4609, 32'hc021d61d} /* (8, 12, 8) {real, imag} */,
  {32'h40bc194c, 32'hc0ba1be7} /* (8, 12, 7) {real, imag} */,
  {32'h3f9475d5, 32'hbf97b1f5} /* (8, 12, 6) {real, imag} */,
  {32'h3ff47cb8, 32'h3f88aa40} /* (8, 12, 5) {real, imag} */,
  {32'hbe5d2fe7, 32'hc09b2270} /* (8, 12, 4) {real, imag} */,
  {32'h3e97bb89, 32'h401f1d7a} /* (8, 12, 3) {real, imag} */,
  {32'h40bf6101, 32'hbf8019da} /* (8, 12, 2) {real, imag} */,
  {32'hc088b986, 32'h40bfab45} /* (8, 12, 1) {real, imag} */,
  {32'h3fed5585, 32'hc0a4b496} /* (8, 12, 0) {real, imag} */,
  {32'h4054b6bb, 32'h408f636f} /* (8, 11, 15) {real, imag} */,
  {32'hc09b5c7e, 32'h40830e65} /* (8, 11, 14) {real, imag} */,
  {32'h40e9bb7a, 32'hc088f43b} /* (8, 11, 13) {real, imag} */,
  {32'h40601161, 32'h40229427} /* (8, 11, 12) {real, imag} */,
  {32'hbfc5f847, 32'hbfca5bea} /* (8, 11, 11) {real, imag} */,
  {32'h3ef454ce, 32'h3ef818c4} /* (8, 11, 10) {real, imag} */,
  {32'hbebed9d7, 32'h3f833808} /* (8, 11, 9) {real, imag} */,
  {32'h408277d5, 32'hc048730e} /* (8, 11, 8) {real, imag} */,
  {32'hbfef94b4, 32'h40a12513} /* (8, 11, 7) {real, imag} */,
  {32'h4035c6b2, 32'h4028fd77} /* (8, 11, 6) {real, imag} */,
  {32'h408b3a2a, 32'h404775a1} /* (8, 11, 5) {real, imag} */,
  {32'h404680b3, 32'h3fe61999} /* (8, 11, 4) {real, imag} */,
  {32'h4088306b, 32'hbfc5e667} /* (8, 11, 3) {real, imag} */,
  {32'hc03f6346, 32'h409af10b} /* (8, 11, 2) {real, imag} */,
  {32'hc047a695, 32'h3f7f3d40} /* (8, 11, 1) {real, imag} */,
  {32'h40631eef, 32'hc029301a} /* (8, 11, 0) {real, imag} */,
  {32'hc02f9191, 32'hbf99414b} /* (8, 10, 15) {real, imag} */,
  {32'hc0a41c80, 32'hc093c8c5} /* (8, 10, 14) {real, imag} */,
  {32'hc04337b4, 32'hc0147e48} /* (8, 10, 13) {real, imag} */,
  {32'h3fbc2327, 32'hc035d7ed} /* (8, 10, 12) {real, imag} */,
  {32'h40a0803d, 32'h3f906a3d} /* (8, 10, 11) {real, imag} */,
  {32'hc0ae0fe2, 32'hc04d6790} /* (8, 10, 10) {real, imag} */,
  {32'h3f816a7c, 32'h409b64e0} /* (8, 10, 9) {real, imag} */,
  {32'h4000f496, 32'h3fe68cb7} /* (8, 10, 8) {real, imag} */,
  {32'hc095f442, 32'h3e9ceeda} /* (8, 10, 7) {real, imag} */,
  {32'hbfb76c3d, 32'h406e1c7a} /* (8, 10, 6) {real, imag} */,
  {32'hc09f73ad, 32'hbfea4449} /* (8, 10, 5) {real, imag} */,
  {32'h400e0cad, 32'h4084f86b} /* (8, 10, 4) {real, imag} */,
  {32'h3eb533cd, 32'hc0688c03} /* (8, 10, 3) {real, imag} */,
  {32'hbfc098b8, 32'h3e8eccba} /* (8, 10, 2) {real, imag} */,
  {32'h40a83aa4, 32'hbf647f5b} /* (8, 10, 1) {real, imag} */,
  {32'hbfcd010a, 32'h4006691b} /* (8, 10, 0) {real, imag} */,
  {32'hc07bcff5, 32'hbef23af8} /* (8, 9, 15) {real, imag} */,
  {32'h40a087ec, 32'h4081a912} /* (8, 9, 14) {real, imag} */,
  {32'hc01aa65b, 32'h40b3f897} /* (8, 9, 13) {real, imag} */,
  {32'hc00be884, 32'hc09b1bff} /* (8, 9, 12) {real, imag} */,
  {32'h404874b2, 32'h40a6677c} /* (8, 9, 11) {real, imag} */,
  {32'hc0027312, 32'h4079102f} /* (8, 9, 10) {real, imag} */,
  {32'h40884181, 32'hbf717fae} /* (8, 9, 9) {real, imag} */,
  {32'hc038c87e, 32'h3f98c385} /* (8, 9, 8) {real, imag} */,
  {32'h3e8f843a, 32'hc0eeb880} /* (8, 9, 7) {real, imag} */,
  {32'h408a08c6, 32'h405ed675} /* (8, 9, 6) {real, imag} */,
  {32'h4082cb14, 32'hbf630d43} /* (8, 9, 5) {real, imag} */,
  {32'h3ea737c1, 32'h3ec576f6} /* (8, 9, 4) {real, imag} */,
  {32'hbe958650, 32'hbf0552d3} /* (8, 9, 3) {real, imag} */,
  {32'hbfcf163a, 32'hc0616cb3} /* (8, 9, 2) {real, imag} */,
  {32'h3fce8745, 32'h3fe17c46} /* (8, 9, 1) {real, imag} */,
  {32'h4009f6bd, 32'hc0844df1} /* (8, 9, 0) {real, imag} */,
  {32'h40cd226f, 32'h3f5fcf42} /* (8, 8, 15) {real, imag} */,
  {32'hbe509d80, 32'hbdba0055} /* (8, 8, 14) {real, imag} */,
  {32'hbf0b18c6, 32'h40217d6a} /* (8, 8, 13) {real, imag} */,
  {32'hbff193ec, 32'hc0248739} /* (8, 8, 12) {real, imag} */,
  {32'hc08403e7, 32'hbeb025c6} /* (8, 8, 11) {real, imag} */,
  {32'h4077cb33, 32'h3f8567d4} /* (8, 8, 10) {real, imag} */,
  {32'hc1034577, 32'h402fdaf2} /* (8, 8, 9) {real, imag} */,
  {32'h40553028, 32'h00000000} /* (8, 8, 8) {real, imag} */,
  {32'hc1034577, 32'hc02fdaf2} /* (8, 8, 7) {real, imag} */,
  {32'h4077cb33, 32'hbf8567d4} /* (8, 8, 6) {real, imag} */,
  {32'hc08403e7, 32'h3eb025c6} /* (8, 8, 5) {real, imag} */,
  {32'hbff193ec, 32'h40248739} /* (8, 8, 4) {real, imag} */,
  {32'hbf0b18c6, 32'hc0217d6a} /* (8, 8, 3) {real, imag} */,
  {32'hbe509d80, 32'h3dba0055} /* (8, 8, 2) {real, imag} */,
  {32'h40cd226f, 32'hbf5fcf42} /* (8, 8, 1) {real, imag} */,
  {32'hbee5c348, 32'h00000000} /* (8, 8, 0) {real, imag} */,
  {32'h3fce8745, 32'hbfe17c46} /* (8, 7, 15) {real, imag} */,
  {32'hbfcf163a, 32'h40616cb3} /* (8, 7, 14) {real, imag} */,
  {32'hbe958650, 32'h3f0552d3} /* (8, 7, 13) {real, imag} */,
  {32'h3ea737c1, 32'hbec576f6} /* (8, 7, 12) {real, imag} */,
  {32'h4082cb14, 32'h3f630d43} /* (8, 7, 11) {real, imag} */,
  {32'h408a08c6, 32'hc05ed675} /* (8, 7, 10) {real, imag} */,
  {32'h3e8f843a, 32'h40eeb880} /* (8, 7, 9) {real, imag} */,
  {32'hc038c87e, 32'hbf98c385} /* (8, 7, 8) {real, imag} */,
  {32'h40884181, 32'h3f717fae} /* (8, 7, 7) {real, imag} */,
  {32'hc0027312, 32'hc079102f} /* (8, 7, 6) {real, imag} */,
  {32'h404874b2, 32'hc0a6677c} /* (8, 7, 5) {real, imag} */,
  {32'hc00be884, 32'h409b1bff} /* (8, 7, 4) {real, imag} */,
  {32'hc01aa65b, 32'hc0b3f897} /* (8, 7, 3) {real, imag} */,
  {32'h40a087ec, 32'hc081a912} /* (8, 7, 2) {real, imag} */,
  {32'hc07bcff5, 32'h3ef23af8} /* (8, 7, 1) {real, imag} */,
  {32'h4009f6bd, 32'h40844df1} /* (8, 7, 0) {real, imag} */,
  {32'h40a83aa4, 32'h3f647f5b} /* (8, 6, 15) {real, imag} */,
  {32'hbfc098b8, 32'hbe8eccba} /* (8, 6, 14) {real, imag} */,
  {32'h3eb533cd, 32'h40688c03} /* (8, 6, 13) {real, imag} */,
  {32'h400e0cad, 32'hc084f86b} /* (8, 6, 12) {real, imag} */,
  {32'hc09f73ad, 32'h3fea4449} /* (8, 6, 11) {real, imag} */,
  {32'hbfb76c3d, 32'hc06e1c7a} /* (8, 6, 10) {real, imag} */,
  {32'hc095f442, 32'hbe9ceeda} /* (8, 6, 9) {real, imag} */,
  {32'h4000f496, 32'hbfe68cb7} /* (8, 6, 8) {real, imag} */,
  {32'h3f816a7c, 32'hc09b64e0} /* (8, 6, 7) {real, imag} */,
  {32'hc0ae0fe2, 32'h404d6790} /* (8, 6, 6) {real, imag} */,
  {32'h40a0803d, 32'hbf906a3d} /* (8, 6, 5) {real, imag} */,
  {32'h3fbc2327, 32'h4035d7ed} /* (8, 6, 4) {real, imag} */,
  {32'hc04337b4, 32'h40147e48} /* (8, 6, 3) {real, imag} */,
  {32'hc0a41c80, 32'h4093c8c5} /* (8, 6, 2) {real, imag} */,
  {32'hc02f9191, 32'h3f99414b} /* (8, 6, 1) {real, imag} */,
  {32'hbfcd010a, 32'hc006691b} /* (8, 6, 0) {real, imag} */,
  {32'hc047a695, 32'hbf7f3d40} /* (8, 5, 15) {real, imag} */,
  {32'hc03f6346, 32'hc09af10b} /* (8, 5, 14) {real, imag} */,
  {32'h4088306b, 32'h3fc5e667} /* (8, 5, 13) {real, imag} */,
  {32'h404680b3, 32'hbfe61999} /* (8, 5, 12) {real, imag} */,
  {32'h408b3a2a, 32'hc04775a1} /* (8, 5, 11) {real, imag} */,
  {32'h4035c6b2, 32'hc028fd77} /* (8, 5, 10) {real, imag} */,
  {32'hbfef94b4, 32'hc0a12513} /* (8, 5, 9) {real, imag} */,
  {32'h408277d5, 32'h4048730e} /* (8, 5, 8) {real, imag} */,
  {32'hbebed9d7, 32'hbf833808} /* (8, 5, 7) {real, imag} */,
  {32'h3ef454ce, 32'hbef818c4} /* (8, 5, 6) {real, imag} */,
  {32'hbfc5f847, 32'h3fca5bea} /* (8, 5, 5) {real, imag} */,
  {32'h40601161, 32'hc0229427} /* (8, 5, 4) {real, imag} */,
  {32'h40e9bb7a, 32'h4088f43b} /* (8, 5, 3) {real, imag} */,
  {32'hc09b5c7e, 32'hc0830e65} /* (8, 5, 2) {real, imag} */,
  {32'h4054b6bb, 32'hc08f636f} /* (8, 5, 1) {real, imag} */,
  {32'h40631eef, 32'h4029301a} /* (8, 5, 0) {real, imag} */,
  {32'hc088b986, 32'hc0bfab45} /* (8, 4, 15) {real, imag} */,
  {32'h40bf6101, 32'h3f8019da} /* (8, 4, 14) {real, imag} */,
  {32'h3e97bb89, 32'hc01f1d7a} /* (8, 4, 13) {real, imag} */,
  {32'hbe5d2fe7, 32'h409b2270} /* (8, 4, 12) {real, imag} */,
  {32'h3ff47cb8, 32'hbf88aa40} /* (8, 4, 11) {real, imag} */,
  {32'h3f9475d5, 32'h3f97b1f5} /* (8, 4, 10) {real, imag} */,
  {32'h40bc194c, 32'h40ba1be7} /* (8, 4, 9) {real, imag} */,
  {32'hc0aa4609, 32'h4021d61d} /* (8, 4, 8) {real, imag} */,
  {32'h3e08f9c4, 32'hc0364a41} /* (8, 4, 7) {real, imag} */,
  {32'hbf53fc1b, 32'h401a11a0} /* (8, 4, 6) {real, imag} */,
  {32'h3fd6631c, 32'hbe6391bc} /* (8, 4, 5) {real, imag} */,
  {32'h3f6e01f1, 32'hc07978b7} /* (8, 4, 4) {real, imag} */,
  {32'hbf57df62, 32'hc09c2da4} /* (8, 4, 3) {real, imag} */,
  {32'h3f01b52f, 32'h401b4fc4} /* (8, 4, 2) {real, imag} */,
  {32'hc0786613, 32'h4033fe43} /* (8, 4, 1) {real, imag} */,
  {32'h3fed5585, 32'h40a4b496} /* (8, 4, 0) {real, imag} */,
  {32'h3f94481c, 32'h40786f7f} /* (8, 3, 15) {real, imag} */,
  {32'hbe217bbc, 32'hbfd89068} /* (8, 3, 14) {real, imag} */,
  {32'hc0b8e7f5, 32'hbfcf5bfa} /* (8, 3, 13) {real, imag} */,
  {32'h3ff5adc1, 32'h40497148} /* (8, 3, 12) {real, imag} */,
  {32'hbfdc7f5f, 32'hc087ef1f} /* (8, 3, 11) {real, imag} */,
  {32'h4063513c, 32'h409efbf2} /* (8, 3, 10) {real, imag} */,
  {32'h3f7b63da, 32'hc079b464} /* (8, 3, 9) {real, imag} */,
  {32'hc01bb076, 32'h402e963c} /* (8, 3, 8) {real, imag} */,
  {32'h409ac016, 32'hc0afa951} /* (8, 3, 7) {real, imag} */,
  {32'h3f7c57c5, 32'hc09bba52} /* (8, 3, 6) {real, imag} */,
  {32'hc0af6895, 32'hbf4aea00} /* (8, 3, 5) {real, imag} */,
  {32'h3fe9521d, 32'hc0308037} /* (8, 3, 4) {real, imag} */,
  {32'h3fc4e28f, 32'h40308128} /* (8, 3, 3) {real, imag} */,
  {32'hbf5ba29d, 32'h3efc837d} /* (8, 3, 2) {real, imag} */,
  {32'hc08c180f, 32'hbf926af5} /* (8, 3, 1) {real, imag} */,
  {32'hc012ca11, 32'hbf2030b6} /* (8, 3, 0) {real, imag} */,
  {32'h3beb754f, 32'h3e4fabe1} /* (8, 2, 15) {real, imag} */,
  {32'hbe3d3be1, 32'hbfb3bcc2} /* (8, 2, 14) {real, imag} */,
  {32'hc009a3f9, 32'h3fb748ed} /* (8, 2, 13) {real, imag} */,
  {32'h40917d64, 32'hc0632195} /* (8, 2, 12) {real, imag} */,
  {32'hbf199ec8, 32'hc0d4c219} /* (8, 2, 11) {real, imag} */,
  {32'h4061a1ae, 32'h3e9a121d} /* (8, 2, 10) {real, imag} */,
  {32'h40b1b11e, 32'hc09f4a87} /* (8, 2, 9) {real, imag} */,
  {32'hbf55d3f1, 32'hc091adcd} /* (8, 2, 8) {real, imag} */,
  {32'h3e2bb16f, 32'h3f4c93f2} /* (8, 2, 7) {real, imag} */,
  {32'h3f69efff, 32'h4016d2b0} /* (8, 2, 6) {real, imag} */,
  {32'h3f773374, 32'hc0b2affa} /* (8, 2, 5) {real, imag} */,
  {32'hbf8a3178, 32'h40926569} /* (8, 2, 4) {real, imag} */,
  {32'hc0218250, 32'h3fca07ff} /* (8, 2, 3) {real, imag} */,
  {32'hbf2e8fbc, 32'hc0a7b849} /* (8, 2, 2) {real, imag} */,
  {32'hbfb09032, 32'h40fb55ca} /* (8, 2, 1) {real, imag} */,
  {32'hbf4b1ed6, 32'hc04de68b} /* (8, 2, 0) {real, imag} */,
  {32'hc0084728, 32'h4097efb8} /* (8, 1, 15) {real, imag} */,
  {32'h3eace800, 32'h40799a92} /* (8, 1, 14) {real, imag} */,
  {32'hbf9bdf2f, 32'hc06898ba} /* (8, 1, 13) {real, imag} */,
  {32'h3f9783da, 32'h3f23e785} /* (8, 1, 12) {real, imag} */,
  {32'h403e3003, 32'hbfc41db7} /* (8, 1, 11) {real, imag} */,
  {32'hc029219a, 32'h3e799fa7} /* (8, 1, 10) {real, imag} */,
  {32'hc02c6cc5, 32'h3f02def3} /* (8, 1, 9) {real, imag} */,
  {32'hbf3cc9c4, 32'hc0038b6f} /* (8, 1, 8) {real, imag} */,
  {32'h402f5752, 32'hc0553b9a} /* (8, 1, 7) {real, imag} */,
  {32'hc0a676b0, 32'h3fecc20a} /* (8, 1, 6) {real, imag} */,
  {32'h3f9ec775, 32'h402b1c06} /* (8, 1, 5) {real, imag} */,
  {32'hc08d7f3d, 32'hbd85d151} /* (8, 1, 4) {real, imag} */,
  {32'h3fc3adbd, 32'hbd206b88} /* (8, 1, 3) {real, imag} */,
  {32'hc08c85a4, 32'h3f30e2d8} /* (8, 1, 2) {real, imag} */,
  {32'h3f1a286a, 32'h3de9f465} /* (8, 1, 1) {real, imag} */,
  {32'hbf48c257, 32'hbf58cac9} /* (8, 1, 0) {real, imag} */,
  {32'h3fb36ca1, 32'hbf8db8ef} /* (8, 0, 15) {real, imag} */,
  {32'h3f5790da, 32'hbecfc14e} /* (8, 0, 14) {real, imag} */,
  {32'h3fa94e74, 32'hbf49ce54} /* (8, 0, 13) {real, imag} */,
  {32'hbfe56e29, 32'hbfa012c7} /* (8, 0, 12) {real, imag} */,
  {32'hbecc0e46, 32'hbf7615e6} /* (8, 0, 11) {real, imag} */,
  {32'h3f98ccf1, 32'h3fa3b223} /* (8, 0, 10) {real, imag} */,
  {32'hc0480726, 32'hc011cb4a} /* (8, 0, 9) {real, imag} */,
  {32'h4062579b, 32'h00000000} /* (8, 0, 8) {real, imag} */,
  {32'hc0480726, 32'h4011cb4a} /* (8, 0, 7) {real, imag} */,
  {32'h3f98ccf1, 32'hbfa3b223} /* (8, 0, 6) {real, imag} */,
  {32'hbecc0e46, 32'h3f7615e6} /* (8, 0, 5) {real, imag} */,
  {32'hbfe56e29, 32'h3fa012c7} /* (8, 0, 4) {real, imag} */,
  {32'h3fa94e74, 32'h3f49ce54} /* (8, 0, 3) {real, imag} */,
  {32'h3f5790da, 32'h3ecfc14e} /* (8, 0, 2) {real, imag} */,
  {32'h3fb36ca1, 32'h3f8db8ef} /* (8, 0, 1) {real, imag} */,
  {32'h3f88e7d7, 32'h00000000} /* (8, 0, 0) {real, imag} */,
  {32'h40ca9fb8, 32'hc0675333} /* (7, 15, 15) {real, imag} */,
  {32'hc0985f6e, 32'hc011b739} /* (7, 15, 14) {real, imag} */,
  {32'h410cd867, 32'hbe8c5e08} /* (7, 15, 13) {real, imag} */,
  {32'hbf104e75, 32'h40196062} /* (7, 15, 12) {real, imag} */,
  {32'h3fe905a8, 32'h410772e0} /* (7, 15, 11) {real, imag} */,
  {32'hc08ad8ac, 32'hc0e9c2e5} /* (7, 15, 10) {real, imag} */,
  {32'hbf1955e6, 32'h3f0a22fd} /* (7, 15, 9) {real, imag} */,
  {32'h3e85dfd6, 32'hc011e83d} /* (7, 15, 8) {real, imag} */,
  {32'hbf2916ec, 32'hc11fa465} /* (7, 15, 7) {real, imag} */,
  {32'hbd68bbc7, 32'h4019abe9} /* (7, 15, 6) {real, imag} */,
  {32'hbf2b8a0b, 32'hc013dc1e} /* (7, 15, 5) {real, imag} */,
  {32'h40712001, 32'h4041ef3d} /* (7, 15, 4) {real, imag} */,
  {32'hc059a2c0, 32'h3eddff66} /* (7, 15, 3) {real, imag} */,
  {32'hbf51de21, 32'h40f094ee} /* (7, 15, 2) {real, imag} */,
  {32'hc09bde59, 32'hc0b342c7} /* (7, 15, 1) {real, imag} */,
  {32'h3f31fe42, 32'hc008de34} /* (7, 15, 0) {real, imag} */,
  {32'hc01383b8, 32'h40aca95d} /* (7, 14, 15) {real, imag} */,
  {32'h4091bbf5, 32'h3fc349b1} /* (7, 14, 14) {real, imag} */,
  {32'hbca2d274, 32'h40a81e70} /* (7, 14, 13) {real, imag} */,
  {32'h40060871, 32'hc0f46aea} /* (7, 14, 12) {real, imag} */,
  {32'hbfb498f6, 32'hc06d93c1} /* (7, 14, 11) {real, imag} */,
  {32'hbf94f29d, 32'hbeb76a21} /* (7, 14, 10) {real, imag} */,
  {32'hbfe7b955, 32'h40465ca2} /* (7, 14, 9) {real, imag} */,
  {32'h408cf9a3, 32'hbf466d81} /* (7, 14, 8) {real, imag} */,
  {32'h4031c1fa, 32'h40c1e573} /* (7, 14, 7) {real, imag} */,
  {32'h3e3706ab, 32'hbfbdf71b} /* (7, 14, 6) {real, imag} */,
  {32'h4105e3c5, 32'h405cec75} /* (7, 14, 5) {real, imag} */,
  {32'hc0d7f14c, 32'h3e84780c} /* (7, 14, 4) {real, imag} */,
  {32'hc02ef342, 32'hbffb1fee} /* (7, 14, 3) {real, imag} */,
  {32'hc02f3545, 32'hc1081825} /* (7, 14, 2) {real, imag} */,
  {32'hc04bfd4d, 32'h407faa7c} /* (7, 14, 1) {real, imag} */,
  {32'h4040cf01, 32'hc00772bc} /* (7, 14, 0) {real, imag} */,
  {32'h3f5f6c16, 32'h3f8b9115} /* (7, 13, 15) {real, imag} */,
  {32'h3f89d2ae, 32'h40faa1b3} /* (7, 13, 14) {real, imag} */,
  {32'h3f884222, 32'hbfa89575} /* (7, 13, 13) {real, imag} */,
  {32'hbff0b52f, 32'hc0bd7452} /* (7, 13, 12) {real, imag} */,
  {32'hbff51f6d, 32'h40250227} /* (7, 13, 11) {real, imag} */,
  {32'h3fa36114, 32'hc040bbc5} /* (7, 13, 10) {real, imag} */,
  {32'hbf5a099d, 32'hc0d1bfe4} /* (7, 13, 9) {real, imag} */,
  {32'h40544907, 32'h3f68561a} /* (7, 13, 8) {real, imag} */,
  {32'hbfbff146, 32'hc02b41a0} /* (7, 13, 7) {real, imag} */,
  {32'hc0052e4b, 32'hbfcdc611} /* (7, 13, 6) {real, imag} */,
  {32'h40d530c9, 32'h409271b1} /* (7, 13, 5) {real, imag} */,
  {32'h407e6017, 32'h3de3f9fd} /* (7, 13, 4) {real, imag} */,
  {32'hc0263166, 32'hbf889fb3} /* (7, 13, 3) {real, imag} */,
  {32'h3e819bd1, 32'h3fb4f295} /* (7, 13, 2) {real, imag} */,
  {32'hc083ecff, 32'hbe84a54c} /* (7, 13, 1) {real, imag} */,
  {32'hc03c433f, 32'h405c7952} /* (7, 13, 0) {real, imag} */,
  {32'h40fa4326, 32'hc102328a} /* (7, 12, 15) {real, imag} */,
  {32'hc05df299, 32'h40be1c8c} /* (7, 12, 14) {real, imag} */,
  {32'h40f45f2a, 32'h408c387b} /* (7, 12, 13) {real, imag} */,
  {32'hbf014628, 32'hc01e2d7d} /* (7, 12, 12) {real, imag} */,
  {32'hbf8e2248, 32'hc00deed5} /* (7, 12, 11) {real, imag} */,
  {32'h3f4b6d42, 32'h40117889} /* (7, 12, 10) {real, imag} */,
  {32'h402f8da6, 32'hbf879f06} /* (7, 12, 9) {real, imag} */,
  {32'h4004b0b9, 32'h3fe09c12} /* (7, 12, 8) {real, imag} */,
  {32'h403e1ea5, 32'hbe686c91} /* (7, 12, 7) {real, imag} */,
  {32'h40a837c9, 32'hc102c6a8} /* (7, 12, 6) {real, imag} */,
  {32'h405bdf03, 32'h40cb59e8} /* (7, 12, 5) {real, imag} */,
  {32'h402e8a36, 32'h40ec3f6e} /* (7, 12, 4) {real, imag} */,
  {32'hc05b5625, 32'hbf9fcd11} /* (7, 12, 3) {real, imag} */,
  {32'h3fbf70d1, 32'hc051ca37} /* (7, 12, 2) {real, imag} */,
  {32'h40621147, 32'hc09bc352} /* (7, 12, 1) {real, imag} */,
  {32'hbf3406e9, 32'h3fb589ac} /* (7, 12, 0) {real, imag} */,
  {32'hc10a6c59, 32'hc12807d9} /* (7, 11, 15) {real, imag} */,
  {32'hbf06a267, 32'h40ca6647} /* (7, 11, 14) {real, imag} */,
  {32'hbf9baa8e, 32'h3e06d77f} /* (7, 11, 13) {real, imag} */,
  {32'h4110620c, 32'h4006a244} /* (7, 11, 12) {real, imag} */,
  {32'h3f70cccb, 32'h3da8ab71} /* (7, 11, 11) {real, imag} */,
  {32'h404e05ec, 32'hbd4105e3} /* (7, 11, 10) {real, imag} */,
  {32'h404a3936, 32'h3f0df615} /* (7, 11, 9) {real, imag} */,
  {32'hc0094ab0, 32'h3fee7737} /* (7, 11, 8) {real, imag} */,
  {32'hc0d5651b, 32'h4123e9ce} /* (7, 11, 7) {real, imag} */,
  {32'h3f2599a1, 32'h3d4d6cac} /* (7, 11, 6) {real, imag} */,
  {32'hc09eb404, 32'h4079ebf6} /* (7, 11, 5) {real, imag} */,
  {32'h3c826fa2, 32'hbf454c96} /* (7, 11, 4) {real, imag} */,
  {32'hc07b15af, 32'hc08b18dd} /* (7, 11, 3) {real, imag} */,
  {32'h3f79056e, 32'hbf3f503f} /* (7, 11, 2) {real, imag} */,
  {32'hc0863532, 32'hc0a33db0} /* (7, 11, 1) {real, imag} */,
  {32'hbcdb2dc5, 32'hc01812fd} /* (7, 11, 0) {real, imag} */,
  {32'h3f951478, 32'h4050caea} /* (7, 10, 15) {real, imag} */,
  {32'h40249209, 32'h408c5564} /* (7, 10, 14) {real, imag} */,
  {32'hc01fbc23, 32'h40cd754e} /* (7, 10, 13) {real, imag} */,
  {32'h3fd35bf1, 32'hc0db67f2} /* (7, 10, 12) {real, imag} */,
  {32'h3f91dccc, 32'h40f3891b} /* (7, 10, 11) {real, imag} */,
  {32'h40adf51c, 32'h40c88a18} /* (7, 10, 10) {real, imag} */,
  {32'h3eb237f6, 32'h40f78634} /* (7, 10, 9) {real, imag} */,
  {32'h408ee152, 32'hc081fe62} /* (7, 10, 8) {real, imag} */,
  {32'h403e00fb, 32'h40a4765b} /* (7, 10, 7) {real, imag} */,
  {32'hc0dab354, 32'h3f2b0e26} /* (7, 10, 6) {real, imag} */,
  {32'hc0ad6944, 32'hc031a6d8} /* (7, 10, 5) {real, imag} */,
  {32'h3f8df11c, 32'hbf78bccc} /* (7, 10, 4) {real, imag} */,
  {32'h40626405, 32'hbf2d3159} /* (7, 10, 3) {real, imag} */,
  {32'hbfc65ed4, 32'hc08d077d} /* (7, 10, 2) {real, imag} */,
  {32'h40ba3b39, 32'h3fff7e5e} /* (7, 10, 1) {real, imag} */,
  {32'h4015ca50, 32'hc0cf4cc9} /* (7, 10, 0) {real, imag} */,
  {32'h4008f173, 32'hc083a825} /* (7, 9, 15) {real, imag} */,
  {32'h401ef6ba, 32'h3fb7ce6c} /* (7, 9, 14) {real, imag} */,
  {32'h3fb44909, 32'h4069160e} /* (7, 9, 13) {real, imag} */,
  {32'hc0383acc, 32'h3f13d7b8} /* (7, 9, 12) {real, imag} */,
  {32'hc0801c4a, 32'h3f238cf2} /* (7, 9, 11) {real, imag} */,
  {32'h3fe3ad74, 32'h3f0baeb4} /* (7, 9, 10) {real, imag} */,
  {32'hc0b6a59b, 32'h407df880} /* (7, 9, 9) {real, imag} */,
  {32'h3f0c9a88, 32'h3fd318f4} /* (7, 9, 8) {real, imag} */,
  {32'hbfac25dd, 32'hbf4bc95f} /* (7, 9, 7) {real, imag} */,
  {32'hbe5fcfb7, 32'h40256498} /* (7, 9, 6) {real, imag} */,
  {32'hc01e3155, 32'h4024a23e} /* (7, 9, 5) {real, imag} */,
  {32'hc1170ca8, 32'hbf18071b} /* (7, 9, 4) {real, imag} */,
  {32'h3f51652e, 32'hbffbbceb} /* (7, 9, 3) {real, imag} */,
  {32'h40ff0c7e, 32'h3e8a28fc} /* (7, 9, 2) {real, imag} */,
  {32'h40c45ed4, 32'hc01536a8} /* (7, 9, 1) {real, imag} */,
  {32'hc05d2f7b, 32'h3fb7b71b} /* (7, 9, 0) {real, imag} */,
  {32'h40b57c67, 32'hbfade9d0} /* (7, 8, 15) {real, imag} */,
  {32'h4000299b, 32'h4001eaae} /* (7, 8, 14) {real, imag} */,
  {32'hbf2781f5, 32'h40687f5c} /* (7, 8, 13) {real, imag} */,
  {32'h404feba2, 32'hc0b1936e} /* (7, 8, 12) {real, imag} */,
  {32'h40aa9f72, 32'h4067d252} /* (7, 8, 11) {real, imag} */,
  {32'hc0b764ab, 32'hbf4ff82e} /* (7, 8, 10) {real, imag} */,
  {32'hbfb16f8a, 32'h4053b18c} /* (7, 8, 9) {real, imag} */,
  {32'hbe553ef0, 32'hc0423d07} /* (7, 8, 8) {real, imag} */,
  {32'h3f25c345, 32'hc09dd412} /* (7, 8, 7) {real, imag} */,
  {32'h3e396329, 32'h3f48f3aa} /* (7, 8, 6) {real, imag} */,
  {32'hc096fdb0, 32'h408e2f59} /* (7, 8, 5) {real, imag} */,
  {32'h3fde5948, 32'hc0c326d8} /* (7, 8, 4) {real, imag} */,
  {32'h403c9130, 32'h4093a4dc} /* (7, 8, 3) {real, imag} */,
  {32'h406f2d9a, 32'hbfbc346c} /* (7, 8, 2) {real, imag} */,
  {32'hbf3c14ef, 32'h3f353ec4} /* (7, 8, 1) {real, imag} */,
  {32'h3fc8dbe6, 32'hbfdac877} /* (7, 8, 0) {real, imag} */,
  {32'hc0c1be00, 32'h3e26e2f0} /* (7, 7, 15) {real, imag} */,
  {32'hc0f1b0fe, 32'h40d09af3} /* (7, 7, 14) {real, imag} */,
  {32'h3fac6fd1, 32'hbfc86ac4} /* (7, 7, 13) {real, imag} */,
  {32'h40d9627c, 32'h40b98589} /* (7, 7, 12) {real, imag} */,
  {32'hbfcdce51, 32'hc112e270} /* (7, 7, 11) {real, imag} */,
  {32'h406f8a8b, 32'hc04a6ca8} /* (7, 7, 10) {real, imag} */,
  {32'hc095e6f6, 32'hc112d930} /* (7, 7, 9) {real, imag} */,
  {32'hbf8cce15, 32'h40032300} /* (7, 7, 8) {real, imag} */,
  {32'hc088da08, 32'hc100dad1} /* (7, 7, 7) {real, imag} */,
  {32'h411ce0f4, 32'h40991c91} /* (7, 7, 6) {real, imag} */,
  {32'hc1127c9b, 32'h402c4ca0} /* (7, 7, 5) {real, imag} */,
  {32'h40807d27, 32'h4082ed68} /* (7, 7, 4) {real, imag} */,
  {32'h40fb32be, 32'h3dbdb0e5} /* (7, 7, 3) {real, imag} */,
  {32'hc01b1346, 32'hc102704e} /* (7, 7, 2) {real, imag} */,
  {32'hbfd22499, 32'hc02f02c8} /* (7, 7, 1) {real, imag} */,
  {32'h408a9d03, 32'h403ad60c} /* (7, 7, 0) {real, imag} */,
  {32'hbf7ab9d1, 32'h3fcae520} /* (7, 6, 15) {real, imag} */,
  {32'h40db68fa, 32'h40a4f364} /* (7, 6, 14) {real, imag} */,
  {32'hc0dc0c4b, 32'hc09efbe9} /* (7, 6, 13) {real, imag} */,
  {32'hc104bf65, 32'hbe65a044} /* (7, 6, 12) {real, imag} */,
  {32'h404b76ce, 32'hc0062f78} /* (7, 6, 11) {real, imag} */,
  {32'h4170e741, 32'hc1461b5e} /* (7, 6, 10) {real, imag} */,
  {32'h3f9cbdc1, 32'hbec7bb41} /* (7, 6, 9) {real, imag} */,
  {32'h3f5a6bed, 32'h40ab2a5b} /* (7, 6, 8) {real, imag} */,
  {32'hc01373c5, 32'h3fe4f24d} /* (7, 6, 7) {real, imag} */,
  {32'hc119ef67, 32'h3fc3c523} /* (7, 6, 6) {real, imag} */,
  {32'h402cdd66, 32'h3e648838} /* (7, 6, 5) {real, imag} */,
  {32'hc08f5de4, 32'hc0c39517} /* (7, 6, 4) {real, imag} */,
  {32'hc0d18296, 32'hbf0857f7} /* (7, 6, 3) {real, imag} */,
  {32'h4066926c, 32'hc04b1f23} /* (7, 6, 2) {real, imag} */,
  {32'h401d07dd, 32'hc0a2cd54} /* (7, 6, 1) {real, imag} */,
  {32'h3fa10601, 32'hc0f3390f} /* (7, 6, 0) {real, imag} */,
  {32'h3f88ef14, 32'hc05ccca0} /* (7, 5, 15) {real, imag} */,
  {32'hbf9ab1ce, 32'hc06fa800} /* (7, 5, 14) {real, imag} */,
  {32'hc0d316eb, 32'hc0a78cae} /* (7, 5, 13) {real, imag} */,
  {32'h40392297, 32'h410b83f9} /* (7, 5, 12) {real, imag} */,
  {32'h40ca91f5, 32'hc02dd03a} /* (7, 5, 11) {real, imag} */,
  {32'h3fb9ea64, 32'h4064b9bb} /* (7, 5, 10) {real, imag} */,
  {32'h4027729f, 32'h4003a442} /* (7, 5, 9) {real, imag} */,
  {32'hbffc1900, 32'h4009f87e} /* (7, 5, 8) {real, imag} */,
  {32'h4103e0a5, 32'h408a81c9} /* (7, 5, 7) {real, imag} */,
  {32'hbfca932a, 32'hc0886d11} /* (7, 5, 6) {real, imag} */,
  {32'h4088b8be, 32'h4065dcd4} /* (7, 5, 5) {real, imag} */,
  {32'hbf66764b, 32'hbf001319} /* (7, 5, 4) {real, imag} */,
  {32'h3fb04b02, 32'hc0997073} /* (7, 5, 3) {real, imag} */,
  {32'hbf659556, 32'h4097dec0} /* (7, 5, 2) {real, imag} */,
  {32'h40bb7f30, 32'h3fbe18ad} /* (7, 5, 1) {real, imag} */,
  {32'hc10c8167, 32'hbffb126a} /* (7, 5, 0) {real, imag} */,
  {32'hc1214886, 32'h402e1db0} /* (7, 4, 15) {real, imag} */,
  {32'h3fca0afb, 32'hc057323f} /* (7, 4, 14) {real, imag} */,
  {32'h3fccaddf, 32'h400bdef9} /* (7, 4, 13) {real, imag} */,
  {32'hbfaaf86b, 32'hc006c8ba} /* (7, 4, 12) {real, imag} */,
  {32'h3fdb7c48, 32'hc09a3d47} /* (7, 4, 11) {real, imag} */,
  {32'h4046be6a, 32'hbf61f04c} /* (7, 4, 10) {real, imag} */,
  {32'hbd47589b, 32'hbfd07b6b} /* (7, 4, 9) {real, imag} */,
  {32'h400d774e, 32'hc040dd61} /* (7, 4, 8) {real, imag} */,
  {32'hbff7e7ea, 32'hbf79634b} /* (7, 4, 7) {real, imag} */,
  {32'hc09b4d4a, 32'hbdf4a12e} /* (7, 4, 6) {real, imag} */,
  {32'hc0aa246d, 32'hc0821627} /* (7, 4, 5) {real, imag} */,
  {32'h3fddd06f, 32'h40ad5887} /* (7, 4, 4) {real, imag} */,
  {32'hc0366f7c, 32'h40b62040} /* (7, 4, 3) {real, imag} */,
  {32'h3fcb6b66, 32'hc053fbf1} /* (7, 4, 2) {real, imag} */,
  {32'hc064d1a7, 32'hc10927ca} /* (7, 4, 1) {real, imag} */,
  {32'h400cfbb2, 32'hbf3e0589} /* (7, 4, 0) {real, imag} */,
  {32'hc0e6906d, 32'hbf6c0388} /* (7, 3, 15) {real, imag} */,
  {32'h407136b8, 32'h4071c8c8} /* (7, 3, 14) {real, imag} */,
  {32'h40556148, 32'h40909178} /* (7, 3, 13) {real, imag} */,
  {32'hc00b431e, 32'hc0e361e0} /* (7, 3, 12) {real, imag} */,
  {32'h3f2d1d8e, 32'hbf296441} /* (7, 3, 11) {real, imag} */,
  {32'hc10026ba, 32'h401a537b} /* (7, 3, 10) {real, imag} */,
  {32'h3fb1b512, 32'hc0c913a7} /* (7, 3, 9) {real, imag} */,
  {32'h3f660fda, 32'hbf9c9939} /* (7, 3, 8) {real, imag} */,
  {32'h3f9b0c86, 32'h3ff7cf3d} /* (7, 3, 7) {real, imag} */,
  {32'hc0a94ba7, 32'h3f859152} /* (7, 3, 6) {real, imag} */,
  {32'hbf121573, 32'hbf764ee5} /* (7, 3, 5) {real, imag} */,
  {32'h40b5fc94, 32'hbfa197f4} /* (7, 3, 4) {real, imag} */,
  {32'h3f6f5d0d, 32'hc021b7ea} /* (7, 3, 3) {real, imag} */,
  {32'hc00565bd, 32'hbf0efb89} /* (7, 3, 2) {real, imag} */,
  {32'h404f4009, 32'hbfbbb82f} /* (7, 3, 1) {real, imag} */,
  {32'hc06117ce, 32'h409db10e} /* (7, 3, 0) {real, imag} */,
  {32'hbf6219d4, 32'h4029cbf7} /* (7, 2, 15) {real, imag} */,
  {32'h3fb5cd7a, 32'h3e4da5a6} /* (7, 2, 14) {real, imag} */,
  {32'h40365d31, 32'hc047a3d7} /* (7, 2, 13) {real, imag} */,
  {32'hbf14a44b, 32'hc09fae46} /* (7, 2, 12) {real, imag} */,
  {32'h40d5e4fe, 32'hbf27560d} /* (7, 2, 11) {real, imag} */,
  {32'h401a59a1, 32'hbe76545a} /* (7, 2, 10) {real, imag} */,
  {32'hc031276f, 32'h4056e18e} /* (7, 2, 9) {real, imag} */,
  {32'h3fcf9302, 32'hc040d707} /* (7, 2, 8) {real, imag} */,
  {32'h4002d012, 32'h3f5288fb} /* (7, 2, 7) {real, imag} */,
  {32'h4102966c, 32'hc08a0951} /* (7, 2, 6) {real, imag} */,
  {32'hc0eaf60b, 32'hc0267e63} /* (7, 2, 5) {real, imag} */,
  {32'h3f465ddb, 32'hc0069e1d} /* (7, 2, 4) {real, imag} */,
  {32'hbfc3c26c, 32'h3d3a9327} /* (7, 2, 3) {real, imag} */,
  {32'hc0da8731, 32'h4060b4c3} /* (7, 2, 2) {real, imag} */,
  {32'h402e2766, 32'hc08dbc34} /* (7, 2, 1) {real, imag} */,
  {32'hbff960a2, 32'h3f9c6d46} /* (7, 2, 0) {real, imag} */,
  {32'hbf882ad3, 32'hbf9d32bc} /* (7, 1, 15) {real, imag} */,
  {32'h3f13acf4, 32'h3f21e3fa} /* (7, 1, 14) {real, imag} */,
  {32'hc09e2b3b, 32'h3fc06208} /* (7, 1, 13) {real, imag} */,
  {32'hc02588d0, 32'hc03669a9} /* (7, 1, 12) {real, imag} */,
  {32'hc0c79ce1, 32'hbf8f1163} /* (7, 1, 11) {real, imag} */,
  {32'h3f9288df, 32'h3facdaab} /* (7, 1, 10) {real, imag} */,
  {32'hbf380436, 32'h4048e755} /* (7, 1, 9) {real, imag} */,
  {32'h400dabdb, 32'h4056e7f8} /* (7, 1, 8) {real, imag} */,
  {32'h3ef7b049, 32'h40888078} /* (7, 1, 7) {real, imag} */,
  {32'hc0f92ba0, 32'h3fc7b229} /* (7, 1, 6) {real, imag} */,
  {32'h410549bd, 32'h410445d9} /* (7, 1, 5) {real, imag} */,
  {32'h3f58ba4a, 32'h40e7cca3} /* (7, 1, 4) {real, imag} */,
  {32'hc0bd4cfe, 32'hc01484ac} /* (7, 1, 3) {real, imag} */,
  {32'h3eddcd7e, 32'h3e59444c} /* (7, 1, 2) {real, imag} */,
  {32'h4101135a, 32'h402d3f08} /* (7, 1, 1) {real, imag} */,
  {32'hbef1e514, 32'hc0727ba6} /* (7, 1, 0) {real, imag} */,
  {32'hc0603ac3, 32'h409351de} /* (7, 0, 15) {real, imag} */,
  {32'h40148df2, 32'hbe8a5b58} /* (7, 0, 14) {real, imag} */,
  {32'hbfd7eca2, 32'hc0d4cf1d} /* (7, 0, 13) {real, imag} */,
  {32'hbe7566c1, 32'h400f9993} /* (7, 0, 12) {real, imag} */,
  {32'h3e936454, 32'h40c84235} /* (7, 0, 11) {real, imag} */,
  {32'hbe1642db, 32'hbfc83b9e} /* (7, 0, 10) {real, imag} */,
  {32'h4016428c, 32'h3f512c4d} /* (7, 0, 9) {real, imag} */,
  {32'hc0d0ebdd, 32'hc08ef88b} /* (7, 0, 8) {real, imag} */,
  {32'h40b0aeed, 32'h3f9446f0} /* (7, 0, 7) {real, imag} */,
  {32'h3fe4ff35, 32'hc11b2b0d} /* (7, 0, 6) {real, imag} */,
  {32'hc0c6ec1c, 32'hbf888e05} /* (7, 0, 5) {real, imag} */,
  {32'hc0085af5, 32'hbec3269f} /* (7, 0, 4) {real, imag} */,
  {32'h40e4bde7, 32'h3ce995a5} /* (7, 0, 3) {real, imag} */,
  {32'hc069b9b0, 32'h4080708b} /* (7, 0, 2) {real, imag} */,
  {32'h40a86f65, 32'h404e0e48} /* (7, 0, 1) {real, imag} */,
  {32'h3faf7242, 32'h40bcc546} /* (7, 0, 0) {real, imag} */,
  {32'hbfec3d3c, 32'hbfd49a6f} /* (6, 15, 15) {real, imag} */,
  {32'h40e0a593, 32'h40d6f6f8} /* (6, 15, 14) {real, imag} */,
  {32'hc0bede06, 32'h40cbf17a} /* (6, 15, 13) {real, imag} */,
  {32'hc01fc859, 32'hbe3988ae} /* (6, 15, 12) {real, imag} */,
  {32'h3fdab7cf, 32'hc03b250d} /* (6, 15, 11) {real, imag} */,
  {32'hbf3c7541, 32'h3f1dd2d4} /* (6, 15, 10) {real, imag} */,
  {32'h403abe91, 32'hc0bd5a66} /* (6, 15, 9) {real, imag} */,
  {32'hbfa40643, 32'hc0416a22} /* (6, 15, 8) {real, imag} */,
  {32'h4152f439, 32'h3fad7fda} /* (6, 15, 7) {real, imag} */,
  {32'h4051de29, 32'hbedc5013} /* (6, 15, 6) {real, imag} */,
  {32'h3f921c0b, 32'h4001440e} /* (6, 15, 5) {real, imag} */,
  {32'hc02ef38e, 32'hbfce023c} /* (6, 15, 4) {real, imag} */,
  {32'h3e5cdbf5, 32'hc047d464} /* (6, 15, 3) {real, imag} */,
  {32'h3f384640, 32'h4111b0f2} /* (6, 15, 2) {real, imag} */,
  {32'h40ffdb88, 32'hbf6890cc} /* (6, 15, 1) {real, imag} */,
  {32'hc11b4135, 32'h40a3b381} /* (6, 15, 0) {real, imag} */,
  {32'hc02ba22b, 32'h4030439b} /* (6, 14, 15) {real, imag} */,
  {32'hc02c631d, 32'hc0f9dc37} /* (6, 14, 14) {real, imag} */,
  {32'hbecaf886, 32'hc06613c5} /* (6, 14, 13) {real, imag} */,
  {32'h400c9b4e, 32'h408ee483} /* (6, 14, 12) {real, imag} */,
  {32'hc0e753a3, 32'h401b48d1} /* (6, 14, 11) {real, imag} */,
  {32'hc0ae81c0, 32'h3eb76558} /* (6, 14, 10) {real, imag} */,
  {32'h4010b239, 32'h4079028a} /* (6, 14, 9) {real, imag} */,
  {32'h40ee1498, 32'hc00cb7cf} /* (6, 14, 8) {real, imag} */,
  {32'hc0ee1057, 32'hbddbd59f} /* (6, 14, 7) {real, imag} */,
  {32'hbfca91a9, 32'hc0eeb14c} /* (6, 14, 6) {real, imag} */,
  {32'hc012e1cf, 32'h40516074} /* (6, 14, 5) {real, imag} */,
  {32'h40bbaaf7, 32'hc0ae9293} /* (6, 14, 4) {real, imag} */,
  {32'h404f2e16, 32'hbe7716ff} /* (6, 14, 3) {real, imag} */,
  {32'hbf44fd32, 32'h4002d7ba} /* (6, 14, 2) {real, imag} */,
  {32'h40accc07, 32'h3fc97fd3} /* (6, 14, 1) {real, imag} */,
  {32'h3febfa15, 32'h401fa633} /* (6, 14, 0) {real, imag} */,
  {32'h40ff9bd4, 32'hc0656826} /* (6, 13, 15) {real, imag} */,
  {32'hc01a4dec, 32'h405933f1} /* (6, 13, 14) {real, imag} */,
  {32'hc0392c66, 32'h4114ae3f} /* (6, 13, 13) {real, imag} */,
  {32'hc06c771f, 32'h4024c8d9} /* (6, 13, 12) {real, imag} */,
  {32'h41515cf5, 32'h3fd181b5} /* (6, 13, 11) {real, imag} */,
  {32'h4020db58, 32'hc0393438} /* (6, 13, 10) {real, imag} */,
  {32'h3f8d924b, 32'h40856e99} /* (6, 13, 9) {real, imag} */,
  {32'h3e1ba08b, 32'h3f63510f} /* (6, 13, 8) {real, imag} */,
  {32'hc084d83a, 32'h3fc63f90} /* (6, 13, 7) {real, imag} */,
  {32'h40396642, 32'hc0ab6f82} /* (6, 13, 6) {real, imag} */,
  {32'h3fac0524, 32'hc00fb32f} /* (6, 13, 5) {real, imag} */,
  {32'hbf899a44, 32'hc1206777} /* (6, 13, 4) {real, imag} */,
  {32'h40580cfe, 32'h40468f54} /* (6, 13, 3) {real, imag} */,
  {32'h40d96efc, 32'hc0bde833} /* (6, 13, 2) {real, imag} */,
  {32'h40a96420, 32'hbf7dde2d} /* (6, 13, 1) {real, imag} */,
  {32'hc0c8a0a6, 32'hc0e48bbd} /* (6, 13, 0) {real, imag} */,
  {32'hbf5737f0, 32'hc0b11624} /* (6, 12, 15) {real, imag} */,
  {32'h3f2c41f9, 32'h3e4f6db8} /* (6, 12, 14) {real, imag} */,
  {32'hc0beaee5, 32'hc033aba1} /* (6, 12, 13) {real, imag} */,
  {32'hbf004fa1, 32'hc0e40fb4} /* (6, 12, 12) {real, imag} */,
  {32'h40cf4d76, 32'h4153eecc} /* (6, 12, 11) {real, imag} */,
  {32'hc07a23f5, 32'hc10c4d02} /* (6, 12, 10) {real, imag} */,
  {32'h403036dd, 32'h406bd83b} /* (6, 12, 9) {real, imag} */,
  {32'h40c1f875, 32'hc02350e3} /* (6, 12, 8) {real, imag} */,
  {32'hc0b65c60, 32'h40b21c9b} /* (6, 12, 7) {real, imag} */,
  {32'h40436d01, 32'h3e471bac} /* (6, 12, 6) {real, imag} */,
  {32'hbed51383, 32'hc05c9194} /* (6, 12, 5) {real, imag} */,
  {32'h40d49f8a, 32'hc1071164} /* (6, 12, 4) {real, imag} */,
  {32'hc151a381, 32'hc0c4c954} /* (6, 12, 3) {real, imag} */,
  {32'h3f9918c2, 32'h40ab5284} /* (6, 12, 2) {real, imag} */,
  {32'hc12bb27a, 32'hc065bec6} /* (6, 12, 1) {real, imag} */,
  {32'h407e74bf, 32'h40eed3c0} /* (6, 12, 0) {real, imag} */,
  {32'h3f849b31, 32'h403635f0} /* (6, 11, 15) {real, imag} */,
  {32'hc04092f2, 32'h3f27db32} /* (6, 11, 14) {real, imag} */,
  {32'hc061a4fb, 32'h40c5ba15} /* (6, 11, 13) {real, imag} */,
  {32'hbfa13528, 32'h408a2d4e} /* (6, 11, 12) {real, imag} */,
  {32'h40b71305, 32'h406a9ebb} /* (6, 11, 11) {real, imag} */,
  {32'hc0d88da6, 32'hc07b8e30} /* (6, 11, 10) {real, imag} */,
  {32'hc04e2ffe, 32'hc0153634} /* (6, 11, 9) {real, imag} */,
  {32'hc05f6828, 32'h40a7b217} /* (6, 11, 8) {real, imag} */,
  {32'h40992b93, 32'hc155a805} /* (6, 11, 7) {real, imag} */,
  {32'hc02c62ff, 32'h41237358} /* (6, 11, 6) {real, imag} */,
  {32'hc03e5615, 32'h409bd9e1} /* (6, 11, 5) {real, imag} */,
  {32'h402eb955, 32'hc13d9594} /* (6, 11, 4) {real, imag} */,
  {32'hc11d5bb4, 32'h3f87edd8} /* (6, 11, 3) {real, imag} */,
  {32'hbfa4d48c, 32'h4054525c} /* (6, 11, 2) {real, imag} */,
  {32'hbf83fe8d, 32'hc0b258f5} /* (6, 11, 1) {real, imag} */,
  {32'h40a18ba8, 32'h4085364f} /* (6, 11, 0) {real, imag} */,
  {32'h40a7ed10, 32'h3e55eb90} /* (6, 10, 15) {real, imag} */,
  {32'hc11ef296, 32'hbfb89451} /* (6, 10, 14) {real, imag} */,
  {32'hc07e6d2f, 32'h407cd2ba} /* (6, 10, 13) {real, imag} */,
  {32'h418fb3aa, 32'hbefad31e} /* (6, 10, 12) {real, imag} */,
  {32'hc0a688c8, 32'hbf4c4813} /* (6, 10, 11) {real, imag} */,
  {32'h4138093e, 32'h3f858ed5} /* (6, 10, 10) {real, imag} */,
  {32'hc0a9a438, 32'hc13cb3db} /* (6, 10, 9) {real, imag} */,
  {32'hc0ca6727, 32'h40963ef1} /* (6, 10, 8) {real, imag} */,
  {32'h411cfeba, 32'h40554832} /* (6, 10, 7) {real, imag} */,
  {32'h406ae90e, 32'h410ad77e} /* (6, 10, 6) {real, imag} */,
  {32'hc1490523, 32'h3fb7e5e6} /* (6, 10, 5) {real, imag} */,
  {32'hbf6cc1da, 32'h409d7f41} /* (6, 10, 4) {real, imag} */,
  {32'h4081e3a7, 32'hc0c30b97} /* (6, 10, 3) {real, imag} */,
  {32'hc0ac6f6d, 32'hc02e0190} /* (6, 10, 2) {real, imag} */,
  {32'hc0c576bb, 32'h3c68b3dd} /* (6, 10, 1) {real, imag} */,
  {32'hbf94544c, 32'hbfe2953b} /* (6, 10, 0) {real, imag} */,
  {32'hc0a2efc5, 32'h3fd577f3} /* (6, 9, 15) {real, imag} */,
  {32'h3f026290, 32'hbfc0263a} /* (6, 9, 14) {real, imag} */,
  {32'hc0dc43a2, 32'hc129a71f} /* (6, 9, 13) {real, imag} */,
  {32'h4028de5f, 32'hc03abb36} /* (6, 9, 12) {real, imag} */,
  {32'h4068ccf1, 32'hbf3b67e4} /* (6, 9, 11) {real, imag} */,
  {32'h407fdc1b, 32'h411d9d10} /* (6, 9, 10) {real, imag} */,
  {32'hc0566b02, 32'h3fa5f9f7} /* (6, 9, 9) {real, imag} */,
  {32'h3f6e30fa, 32'hc07bb9c0} /* (6, 9, 8) {real, imag} */,
  {32'h3cdfba8c, 32'h3ff481a3} /* (6, 9, 7) {real, imag} */,
  {32'hbeb2ae6f, 32'h3ec3dd7a} /* (6, 9, 6) {real, imag} */,
  {32'hc056ee7b, 32'h4000250b} /* (6, 9, 5) {real, imag} */,
  {32'h3ea47289, 32'h41280341} /* (6, 9, 4) {real, imag} */,
  {32'h3e7556d0, 32'h3f6f89c9} /* (6, 9, 3) {real, imag} */,
  {32'hc05e8412, 32'hc10603a7} /* (6, 9, 2) {real, imag} */,
  {32'h3fc7c5f5, 32'h40596035} /* (6, 9, 1) {real, imag} */,
  {32'h4090f1bc, 32'h403d83f0} /* (6, 9, 0) {real, imag} */,
  {32'hc05963d9, 32'hbf11e4e1} /* (6, 8, 15) {real, imag} */,
  {32'h3fc95f0c, 32'h3ffe14bb} /* (6, 8, 14) {real, imag} */,
  {32'h3d10eef0, 32'h3fed7a44} /* (6, 8, 13) {real, imag} */,
  {32'hbfbb8f20, 32'hc003cb26} /* (6, 8, 12) {real, imag} */,
  {32'h40c680d8, 32'hbfe309a0} /* (6, 8, 11) {real, imag} */,
  {32'h3ffefe22, 32'hc08f5871} /* (6, 8, 10) {real, imag} */,
  {32'h3d87c7b7, 32'h407d4c80} /* (6, 8, 9) {real, imag} */,
  {32'hbf4b2f46, 32'hc003acfa} /* (6, 8, 8) {real, imag} */,
  {32'h4095afef, 32'h400cf2c2} /* (6, 8, 7) {real, imag} */,
  {32'h410a590b, 32'h405efde6} /* (6, 8, 6) {real, imag} */,
  {32'hc0999cb0, 32'hc0e0aa41} /* (6, 8, 5) {real, imag} */,
  {32'h3fa3bfa7, 32'h407d7899} /* (6, 8, 4) {real, imag} */,
  {32'hc002f77a, 32'hc0b5a370} /* (6, 8, 3) {real, imag} */,
  {32'hc0516d77, 32'h40c50c65} /* (6, 8, 2) {real, imag} */,
  {32'h40b55f5f, 32'h3fb82a33} /* (6, 8, 1) {real, imag} */,
  {32'h400fc950, 32'h40535aa0} /* (6, 8, 0) {real, imag} */,
  {32'hbee5cae5, 32'hbf871604} /* (6, 7, 15) {real, imag} */,
  {32'hbf40858b, 32'hbf70eb2a} /* (6, 7, 14) {real, imag} */,
  {32'h410f00ba, 32'hc13194f1} /* (6, 7, 13) {real, imag} */,
  {32'h3e63f6d8, 32'hc05bbc13} /* (6, 7, 12) {real, imag} */,
  {32'h40448fcc, 32'h40a6b9c4} /* (6, 7, 11) {real, imag} */,
  {32'hc088b411, 32'h40417572} /* (6, 7, 10) {real, imag} */,
  {32'hc0ae1e76, 32'hc05cac02} /* (6, 7, 9) {real, imag} */,
  {32'h40f39702, 32'hc0cc3dec} /* (6, 7, 8) {real, imag} */,
  {32'hbf7c5da0, 32'h40964a06} /* (6, 7, 7) {real, imag} */,
  {32'h40785883, 32'h3fe9ab22} /* (6, 7, 6) {real, imag} */,
  {32'h402723fa, 32'hc14d4e2d} /* (6, 7, 5) {real, imag} */,
  {32'hc081f871, 32'h400ccc1f} /* (6, 7, 4) {real, imag} */,
  {32'hc0d21769, 32'hbfd09199} /* (6, 7, 3) {real, imag} */,
  {32'hc09557a6, 32'h40876579} /* (6, 7, 2) {real, imag} */,
  {32'hc09e519e, 32'h3e133e13} /* (6, 7, 1) {real, imag} */,
  {32'h40b7ab4d, 32'hbfd99b01} /* (6, 7, 0) {real, imag} */,
  {32'hc089bdf5, 32'hc0aa1d6d} /* (6, 6, 15) {real, imag} */,
  {32'hc074a9d0, 32'h3fe1050d} /* (6, 6, 14) {real, imag} */,
  {32'hc0454066, 32'hbfd93ff6} /* (6, 6, 13) {real, imag} */,
  {32'h40bff674, 32'h4105d851} /* (6, 6, 12) {real, imag} */,
  {32'hbf8351c8, 32'h40df1d2a} /* (6, 6, 11) {real, imag} */,
  {32'h40850aab, 32'hc09ed226} /* (6, 6, 10) {real, imag} */,
  {32'h40d249de, 32'h3fe5e92f} /* (6, 6, 9) {real, imag} */,
  {32'h3fe5bfd5, 32'h4035a36e} /* (6, 6, 8) {real, imag} */,
  {32'hbf306a9f, 32'hc03f020d} /* (6, 6, 7) {real, imag} */,
  {32'h41002cd9, 32'h407b7514} /* (6, 6, 6) {real, imag} */,
  {32'h4064af94, 32'h3f16ee70} /* (6, 6, 5) {real, imag} */,
  {32'hc0128c2b, 32'h40ea59f5} /* (6, 6, 4) {real, imag} */,
  {32'hbe84ca8d, 32'h3f442bb0} /* (6, 6, 3) {real, imag} */,
  {32'h40dd7d5b, 32'hc0c99a6b} /* (6, 6, 2) {real, imag} */,
  {32'h404ffc42, 32'hc04d87a2} /* (6, 6, 1) {real, imag} */,
  {32'hc1109b5c, 32'hc04d597d} /* (6, 6, 0) {real, imag} */,
  {32'h3f072f72, 32'hbf14322f} /* (6, 5, 15) {real, imag} */,
  {32'h3f16184d, 32'hc0c11994} /* (6, 5, 14) {real, imag} */,
  {32'hbf60f8ec, 32'h4152a809} /* (6, 5, 13) {real, imag} */,
  {32'hc037697d, 32'hc10acf09} /* (6, 5, 12) {real, imag} */,
  {32'h3ff9bde9, 32'h3f72b9a5} /* (6, 5, 11) {real, imag} */,
  {32'h40426323, 32'h4015bad8} /* (6, 5, 10) {real, imag} */,
  {32'hc0340a47, 32'hc0822b20} /* (6, 5, 9) {real, imag} */,
  {32'hc07bf31f, 32'h40844e97} /* (6, 5, 8) {real, imag} */,
  {32'hc0eff9ff, 32'hc1341868} /* (6, 5, 7) {real, imag} */,
  {32'hc0ea8c1b, 32'h40969eb0} /* (6, 5, 6) {real, imag} */,
  {32'h3e730f2f, 32'h413d8962} /* (6, 5, 5) {real, imag} */,
  {32'hc10480d6, 32'h40195d59} /* (6, 5, 4) {real, imag} */,
  {32'h40fbb959, 32'hc0add896} /* (6, 5, 3) {real, imag} */,
  {32'hbf055506, 32'hc12c5fae} /* (6, 5, 2) {real, imag} */,
  {32'h40f6a19c, 32'h3e872390} /* (6, 5, 1) {real, imag} */,
  {32'h40299827, 32'h40eb0c45} /* (6, 5, 0) {real, imag} */,
  {32'h40d4f4d2, 32'hc0d05cff} /* (6, 4, 15) {real, imag} */,
  {32'hc0e994a1, 32'h40361171} /* (6, 4, 14) {real, imag} */,
  {32'hbfe5b401, 32'h3f725c54} /* (6, 4, 13) {real, imag} */,
  {32'h405ac727, 32'h3f2da4da} /* (6, 4, 12) {real, imag} */,
  {32'hc06236ec, 32'h3eb19665} /* (6, 4, 11) {real, imag} */,
  {32'hc0eece7c, 32'h3fe3a78a} /* (6, 4, 10) {real, imag} */,
  {32'h3e780501, 32'hc08e76f5} /* (6, 4, 9) {real, imag} */,
  {32'h3f7022d0, 32'hc1269ce6} /* (6, 4, 8) {real, imag} */,
  {32'hc081119e, 32'hc043de81} /* (6, 4, 7) {real, imag} */,
  {32'h4090276d, 32'h401d197d} /* (6, 4, 6) {real, imag} */,
  {32'h3fe201ab, 32'hbfd55aaa} /* (6, 4, 5) {real, imag} */,
  {32'hc148a072, 32'hbf1fd9d8} /* (6, 4, 4) {real, imag} */,
  {32'hc008fbb8, 32'hc0634149} /* (6, 4, 3) {real, imag} */,
  {32'h40f4a8dd, 32'h40e7248c} /* (6, 4, 2) {real, imag} */,
  {32'h40bec05e, 32'h3fd35f61} /* (6, 4, 1) {real, imag} */,
  {32'hc0900b90, 32'h4062129d} /* (6, 4, 0) {real, imag} */,
  {32'hc04810f6, 32'hc00d4d95} /* (6, 3, 15) {real, imag} */,
  {32'hbe289dc3, 32'h3f575d38} /* (6, 3, 14) {real, imag} */,
  {32'h40415d2f, 32'h410a73d3} /* (6, 3, 13) {real, imag} */,
  {32'h40a00933, 32'h400015a9} /* (6, 3, 12) {real, imag} */,
  {32'h3f4f2d02, 32'hc026650d} /* (6, 3, 11) {real, imag} */,
  {32'hbfe5dd5f, 32'h4020d6d4} /* (6, 3, 10) {real, imag} */,
  {32'hbfa34486, 32'h406de7ab} /* (6, 3, 9) {real, imag} */,
  {32'hbf41f644, 32'h40179977} /* (6, 3, 8) {real, imag} */,
  {32'h407188c1, 32'h40503a8d} /* (6, 3, 7) {real, imag} */,
  {32'hc093c5b1, 32'hbe5760b1} /* (6, 3, 6) {real, imag} */,
  {32'h3fc02dce, 32'h3fec1fb9} /* (6, 3, 5) {real, imag} */,
  {32'h409b2498, 32'h40521712} /* (6, 3, 4) {real, imag} */,
  {32'hc0ba0199, 32'h406b0e0e} /* (6, 3, 3) {real, imag} */,
  {32'h3f10b93f, 32'h40a5471f} /* (6, 3, 2) {real, imag} */,
  {32'hbf2300ed, 32'hc09a6b0c} /* (6, 3, 1) {real, imag} */,
  {32'hbd23c333, 32'hc0e95153} /* (6, 3, 0) {real, imag} */,
  {32'h40e4dd0d, 32'h40b1d8a1} /* (6, 2, 15) {real, imag} */,
  {32'hc105fa01, 32'hbf90b79b} /* (6, 2, 14) {real, imag} */,
  {32'h4070c678, 32'h3eabdb06} /* (6, 2, 13) {real, imag} */,
  {32'h3f691606, 32'h40cc3b25} /* (6, 2, 12) {real, imag} */,
  {32'hc09fcbfb, 32'hbf3ef20b} /* (6, 2, 11) {real, imag} */,
  {32'h3ff591b9, 32'hc04adb02} /* (6, 2, 10) {real, imag} */,
  {32'hc008346d, 32'h3e7c28ca} /* (6, 2, 9) {real, imag} */,
  {32'h3fce58d7, 32'h4006b15c} /* (6, 2, 8) {real, imag} */,
  {32'h4092ef2c, 32'h400e2791} /* (6, 2, 7) {real, imag} */,
  {32'hbf79f3c6, 32'hbfe6f805} /* (6, 2, 6) {real, imag} */,
  {32'h40f170f1, 32'h40e6ce79} /* (6, 2, 5) {real, imag} */,
  {32'hc088c6d3, 32'hc134f836} /* (6, 2, 4) {real, imag} */,
  {32'h40c9a0a7, 32'hbfdfe6ea} /* (6, 2, 3) {real, imag} */,
  {32'hc0077d63, 32'h4010def7} /* (6, 2, 2) {real, imag} */,
  {32'hc17eef01, 32'h40548105} /* (6, 2, 1) {real, imag} */,
  {32'h4110ae5d, 32'h40dafafe} /* (6, 2, 0) {real, imag} */,
  {32'hc06a8b5d, 32'h404afcf2} /* (6, 1, 15) {real, imag} */,
  {32'hc11f946e, 32'h3fa6ee4a} /* (6, 1, 14) {real, imag} */,
  {32'hc0aebe51, 32'h40ff6b9b} /* (6, 1, 13) {real, imag} */,
  {32'h41178f86, 32'h412d5c8a} /* (6, 1, 12) {real, imag} */,
  {32'hc0016147, 32'h402718a7} /* (6, 1, 11) {real, imag} */,
  {32'hc082a46b, 32'hc0a6714e} /* (6, 1, 10) {real, imag} */,
  {32'h4042edd5, 32'h4049572e} /* (6, 1, 9) {real, imag} */,
  {32'hc009c4a2, 32'hc02f33dd} /* (6, 1, 8) {real, imag} */,
  {32'hbf8a062c, 32'h3fd5d2d3} /* (6, 1, 7) {real, imag} */,
  {32'h411cf580, 32'h405cf0d8} /* (6, 1, 6) {real, imag} */,
  {32'h404732de, 32'h40d80a35} /* (6, 1, 5) {real, imag} */,
  {32'h3f31ed04, 32'hbfc3fcc3} /* (6, 1, 4) {real, imag} */,
  {32'h3fab0424, 32'h4149d60c} /* (6, 1, 3) {real, imag} */,
  {32'hc00fc011, 32'h3f62af50} /* (6, 1, 2) {real, imag} */,
  {32'h4020ac32, 32'hc02bffcf} /* (6, 1, 1) {real, imag} */,
  {32'h411d7d8b, 32'hc020db05} /* (6, 1, 0) {real, imag} */,
  {32'h40483413, 32'hc09376e5} /* (6, 0, 15) {real, imag} */,
  {32'h411ddfd9, 32'h400d9f7b} /* (6, 0, 14) {real, imag} */,
  {32'hc02ed998, 32'hc0aab37c} /* (6, 0, 13) {real, imag} */,
  {32'hc0b42b44, 32'hc0ac0006} /* (6, 0, 12) {real, imag} */,
  {32'hc0725f66, 32'h3f9ab391} /* (6, 0, 11) {real, imag} */,
  {32'h40a1c530, 32'h3f3821c3} /* (6, 0, 10) {real, imag} */,
  {32'hbeef7dc4, 32'h3fbed9ba} /* (6, 0, 9) {real, imag} */,
  {32'hc036a137, 32'hc011727e} /* (6, 0, 8) {real, imag} */,
  {32'hbff6f7fa, 32'h3f99c1b5} /* (6, 0, 7) {real, imag} */,
  {32'hc06862da, 32'h3fdf273b} /* (6, 0, 6) {real, imag} */,
  {32'hc0a6258d, 32'hbf33b50a} /* (6, 0, 5) {real, imag} */,
  {32'h40083a22, 32'h3fbfc246} /* (6, 0, 4) {real, imag} */,
  {32'hc027a5c5, 32'h3f55525f} /* (6, 0, 3) {real, imag} */,
  {32'hc10c4f85, 32'hc0bacf57} /* (6, 0, 2) {real, imag} */,
  {32'h3f5f6514, 32'hc0264903} /* (6, 0, 1) {real, imag} */,
  {32'h3f3dcb7f, 32'h400488f1} /* (6, 0, 0) {real, imag} */,
  {32'h404f2d57, 32'hc0a56c76} /* (5, 15, 15) {real, imag} */,
  {32'hbf9b97af, 32'hbef5ffc1} /* (5, 15, 14) {real, imag} */,
  {32'h40526b80, 32'hbff8ee83} /* (5, 15, 13) {real, imag} */,
  {32'h3f37e4ae, 32'hbfbe09f6} /* (5, 15, 12) {real, imag} */,
  {32'hc1355d6f, 32'h40c7b7ec} /* (5, 15, 11) {real, imag} */,
  {32'h414f3a39, 32'hc0052813} /* (5, 15, 10) {real, imag} */,
  {32'h4049016e, 32'hbf8ebf44} /* (5, 15, 9) {real, imag} */,
  {32'hbe9df1f0, 32'hbf8c4fd9} /* (5, 15, 8) {real, imag} */,
  {32'h3fb34c25, 32'h401a3ff6} /* (5, 15, 7) {real, imag} */,
  {32'hbfc79da7, 32'h3fa37064} /* (5, 15, 6) {real, imag} */,
  {32'hbe71d7a3, 32'hc0a4cef8} /* (5, 15, 5) {real, imag} */,
  {32'h40f4e93c, 32'h40d41d91} /* (5, 15, 4) {real, imag} */,
  {32'hbfcc3d28, 32'hc09be3b5} /* (5, 15, 3) {real, imag} */,
  {32'h40e9010e, 32'hbf724221} /* (5, 15, 2) {real, imag} */,
  {32'h40bf30e4, 32'h3fcd10d9} /* (5, 15, 1) {real, imag} */,
  {32'h40642f82, 32'hc0153326} /* (5, 15, 0) {real, imag} */,
  {32'h3f1368d2, 32'hc0aead62} /* (5, 14, 15) {real, imag} */,
  {32'hc0a5ade9, 32'hc08f00cc} /* (5, 14, 14) {real, imag} */,
  {32'hc086cfcd, 32'hc1009aa4} /* (5, 14, 13) {real, imag} */,
  {32'h3ffd5a57, 32'h41004f77} /* (5, 14, 12) {real, imag} */,
  {32'hbf808fae, 32'h402cada2} /* (5, 14, 11) {real, imag} */,
  {32'hc1068bdd, 32'hc08b3115} /* (5, 14, 10) {real, imag} */,
  {32'h410c6495, 32'h414b85cc} /* (5, 14, 9) {real, imag} */,
  {32'h4084c774, 32'hbfc8508b} /* (5, 14, 8) {real, imag} */,
  {32'hbf6f163c, 32'hc03f6ada} /* (5, 14, 7) {real, imag} */,
  {32'h412846b4, 32'h40bcb93a} /* (5, 14, 6) {real, imag} */,
  {32'h40ab8a81, 32'h410da436} /* (5, 14, 5) {real, imag} */,
  {32'hbf526e52, 32'h40b49eec} /* (5, 14, 4) {real, imag} */,
  {32'hc0cc2f25, 32'hc11bc6d2} /* (5, 14, 3) {real, imag} */,
  {32'h3f410110, 32'h40c62d31} /* (5, 14, 2) {real, imag} */,
  {32'h4093710e, 32'hbfd16966} /* (5, 14, 1) {real, imag} */,
  {32'hbefa3045, 32'h408800db} /* (5, 14, 0) {real, imag} */,
  {32'h40633218, 32'h40803132} /* (5, 13, 15) {real, imag} */,
  {32'hc09bd049, 32'hc020ced7} /* (5, 13, 14) {real, imag} */,
  {32'h403b45a1, 32'hc0a34135} /* (5, 13, 13) {real, imag} */,
  {32'h4033b9d4, 32'hc0a2e666} /* (5, 13, 12) {real, imag} */,
  {32'h41017e70, 32'h403d2c1d} /* (5, 13, 11) {real, imag} */,
  {32'hbff8f681, 32'hc06186fc} /* (5, 13, 10) {real, imag} */,
  {32'h3fa8279c, 32'h4022ab8c} /* (5, 13, 9) {real, imag} */,
  {32'h3f28e9cd, 32'h3f0492e4} /* (5, 13, 8) {real, imag} */,
  {32'hbea92559, 32'hbf18009f} /* (5, 13, 7) {real, imag} */,
  {32'hc0f12eba, 32'h3fb2476a} /* (5, 13, 6) {real, imag} */,
  {32'h4085ba9b, 32'h409f02f8} /* (5, 13, 5) {real, imag} */,
  {32'hbfb1b785, 32'hc0ca569e} /* (5, 13, 4) {real, imag} */,
  {32'h402ea681, 32'h40a65c7c} /* (5, 13, 3) {real, imag} */,
  {32'h40dbced6, 32'hc11de712} /* (5, 13, 2) {real, imag} */,
  {32'hc00c28c6, 32'h3f18be7b} /* (5, 13, 1) {real, imag} */,
  {32'hbffd7526, 32'h3f75d0ff} /* (5, 13, 0) {real, imag} */,
  {32'h3faba832, 32'hbf3884d4} /* (5, 12, 15) {real, imag} */,
  {32'h41084e61, 32'hc0990be5} /* (5, 12, 14) {real, imag} */,
  {32'h400ad92e, 32'h4082242a} /* (5, 12, 13) {real, imag} */,
  {32'h40bf9708, 32'h3e12c02b} /* (5, 12, 12) {real, imag} */,
  {32'hbfbebc3b, 32'hc0c5e84f} /* (5, 12, 11) {real, imag} */,
  {32'h3ff4ed63, 32'h410110b6} /* (5, 12, 10) {real, imag} */,
  {32'hc0f29573, 32'h404b553a} /* (5, 12, 9) {real, imag} */,
  {32'h4028b071, 32'h40afe22c} /* (5, 12, 8) {real, imag} */,
  {32'hc09e5a25, 32'hc0b3466f} /* (5, 12, 7) {real, imag} */,
  {32'h40be17d1, 32'hc0fab5c7} /* (5, 12, 6) {real, imag} */,
  {32'hc0d29ed5, 32'h410539da} /* (5, 12, 5) {real, imag} */,
  {32'hc0176d8c, 32'hc068baf8} /* (5, 12, 4) {real, imag} */,
  {32'h40048715, 32'h406379c3} /* (5, 12, 3) {real, imag} */,
  {32'hc10b0939, 32'hbf2879f1} /* (5, 12, 2) {real, imag} */,
  {32'hc054154a, 32'hbf5f838e} /* (5, 12, 1) {real, imag} */,
  {32'h4096f19a, 32'h40477501} /* (5, 12, 0) {real, imag} */,
  {32'h3f477123, 32'h404a9503} /* (5, 11, 15) {real, imag} */,
  {32'hc0b2eec9, 32'hc0efb792} /* (5, 11, 14) {real, imag} */,
  {32'hbf09d576, 32'h3fc5851f} /* (5, 11, 13) {real, imag} */,
  {32'hc06df3a4, 32'h40d419d3} /* (5, 11, 12) {real, imag} */,
  {32'hbfc6c6e1, 32'h40984d9c} /* (5, 11, 11) {real, imag} */,
  {32'h3eddb8b3, 32'h3f0f833a} /* (5, 11, 10) {real, imag} */,
  {32'h3fea5039, 32'hc0ad34c7} /* (5, 11, 9) {real, imag} */,
  {32'hc0841f8c, 32'hc0328ca8} /* (5, 11, 8) {real, imag} */,
  {32'hbf1fd540, 32'hc0c166c0} /* (5, 11, 7) {real, imag} */,
  {32'hc109e2c9, 32'h3f4c1972} /* (5, 11, 6) {real, imag} */,
  {32'h40e6beac, 32'hc0607d44} /* (5, 11, 5) {real, imag} */,
  {32'h3f70ff71, 32'h40810eaf} /* (5, 11, 4) {real, imag} */,
  {32'h3f2263f8, 32'h40d1f1e8} /* (5, 11, 3) {real, imag} */,
  {32'hbfda8f36, 32'hc16bc2dc} /* (5, 11, 2) {real, imag} */,
  {32'h3fb02741, 32'h4083a9e7} /* (5, 11, 1) {real, imag} */,
  {32'h4097f439, 32'hc05931a8} /* (5, 11, 0) {real, imag} */,
  {32'hc08b212e, 32'h405cf036} /* (5, 10, 15) {real, imag} */,
  {32'h4035916d, 32'h40c126a5} /* (5, 10, 14) {real, imag} */,
  {32'h4047c6c9, 32'h409fd691} /* (5, 10, 13) {real, imag} */,
  {32'hc0456fca, 32'h406c6797} /* (5, 10, 12) {real, imag} */,
  {32'h40cbde19, 32'h4057811c} /* (5, 10, 11) {real, imag} */,
  {32'h3fe71f5c, 32'hbecbfd8b} /* (5, 10, 10) {real, imag} */,
  {32'hc062346d, 32'hbff40115} /* (5, 10, 9) {real, imag} */,
  {32'h3e80d6b8, 32'h4051d688} /* (5, 10, 8) {real, imag} */,
  {32'h3f50e12d, 32'hc04b0a6c} /* (5, 10, 7) {real, imag} */,
  {32'hc099c31d, 32'h401c5f65} /* (5, 10, 6) {real, imag} */,
  {32'h40a3c469, 32'hc127cab8} /* (5, 10, 5) {real, imag} */,
  {32'h40a96624, 32'hc08e6083} /* (5, 10, 4) {real, imag} */,
  {32'h3fa2780a, 32'h40f0053a} /* (5, 10, 3) {real, imag} */,
  {32'h40100b48, 32'h405f959b} /* (5, 10, 2) {real, imag} */,
  {32'hbf0a301a, 32'h411ddbfe} /* (5, 10, 1) {real, imag} */,
  {32'hc0c804f2, 32'hc081374b} /* (5, 10, 0) {real, imag} */,
  {32'h3f8bdc33, 32'hc005c69c} /* (5, 9, 15) {real, imag} */,
  {32'h3ffe536e, 32'hbfb8f510} /* (5, 9, 14) {real, imag} */,
  {32'h3fe8e818, 32'hc0a7fd9f} /* (5, 9, 13) {real, imag} */,
  {32'hc04ed7a6, 32'h410b4a74} /* (5, 9, 12) {real, imag} */,
  {32'hbfa85070, 32'h4079dd28} /* (5, 9, 11) {real, imag} */,
  {32'h3facb8b0, 32'hc0df4759} /* (5, 9, 10) {real, imag} */,
  {32'h4010eb51, 32'hc01d9459} /* (5, 9, 9) {real, imag} */,
  {32'hc04b440c, 32'hc0f0ab3d} /* (5, 9, 8) {real, imag} */,
  {32'hc0c69534, 32'hbfbad0e0} /* (5, 9, 7) {real, imag} */,
  {32'h402ca0af, 32'h404fb022} /* (5, 9, 6) {real, imag} */,
  {32'hc09707c6, 32'hbfedba5e} /* (5, 9, 5) {real, imag} */,
  {32'h3ef0cdca, 32'h40350b72} /* (5, 9, 4) {real, imag} */,
  {32'hbee6990a, 32'hbfb276b9} /* (5, 9, 3) {real, imag} */,
  {32'hc0db1d13, 32'h400de8c2} /* (5, 9, 2) {real, imag} */,
  {32'h40d2e79b, 32'hc0a1e8fd} /* (5, 9, 1) {real, imag} */,
  {32'h3e9a8d38, 32'h40a6e2c2} /* (5, 9, 0) {real, imag} */,
  {32'hbf73edbf, 32'hc0e02ec9} /* (5, 8, 15) {real, imag} */,
  {32'h40057087, 32'hbf37e4de} /* (5, 8, 14) {real, imag} */,
  {32'h40b6d0e3, 32'h4073e0ef} /* (5, 8, 13) {real, imag} */,
  {32'h40ef33ff, 32'h3e6bbe05} /* (5, 8, 12) {real, imag} */,
  {32'h40e19ccb, 32'hc06bcee1} /* (5, 8, 11) {real, imag} */,
  {32'hc05b201a, 32'hc038b552} /* (5, 8, 10) {real, imag} */,
  {32'hc08ca80b, 32'h40a9bc9c} /* (5, 8, 9) {real, imag} */,
  {32'h3d058620, 32'h4011c020} /* (5, 8, 8) {real, imag} */,
  {32'h409539bd, 32'hc000d86f} /* (5, 8, 7) {real, imag} */,
  {32'hbfe4af93, 32'h3da3e51b} /* (5, 8, 6) {real, imag} */,
  {32'h3a88daf7, 32'hc022c0b7} /* (5, 8, 5) {real, imag} */,
  {32'hbfd7312d, 32'hc02707bf} /* (5, 8, 4) {real, imag} */,
  {32'h4058cf91, 32'h3f890541} /* (5, 8, 3) {real, imag} */,
  {32'hc08163f1, 32'hc010adc1} /* (5, 8, 2) {real, imag} */,
  {32'h400b462a, 32'h408cd555} /* (5, 8, 1) {real, imag} */,
  {32'hc053f04c, 32'h407417de} /* (5, 8, 0) {real, imag} */,
  {32'hc01e7d24, 32'hbeaa6fe8} /* (5, 7, 15) {real, imag} */,
  {32'hc014c713, 32'h40113621} /* (5, 7, 14) {real, imag} */,
  {32'h40781707, 32'hc0c32605} /* (5, 7, 13) {real, imag} */,
  {32'hc00d2178, 32'hbf59ccb7} /* (5, 7, 12) {real, imag} */,
  {32'h406928e3, 32'h408ec0c7} /* (5, 7, 11) {real, imag} */,
  {32'hc0802a35, 32'h4069bb1b} /* (5, 7, 10) {real, imag} */,
  {32'hc030e8e8, 32'hc0815776} /* (5, 7, 9) {real, imag} */,
  {32'h4094aec0, 32'h405b8b1a} /* (5, 7, 8) {real, imag} */,
  {32'h40c827f3, 32'h4028f6a5} /* (5, 7, 7) {real, imag} */,
  {32'hc0c06ccb, 32'hc0c325a3} /* (5, 7, 6) {real, imag} */,
  {32'hbfb85363, 32'hbf7f4644} /* (5, 7, 5) {real, imag} */,
  {32'h40abbad0, 32'hc10cbbad} /* (5, 7, 4) {real, imag} */,
  {32'h40c92d4b, 32'h400822e2} /* (5, 7, 3) {real, imag} */,
  {32'h401a3054, 32'h4076bdd9} /* (5, 7, 2) {real, imag} */,
  {32'hc0938435, 32'h40b660d1} /* (5, 7, 1) {real, imag} */,
  {32'h3f293aef, 32'h40791faf} /* (5, 7, 0) {real, imag} */,
  {32'hc085940c, 32'h40157d81} /* (5, 6, 15) {real, imag} */,
  {32'hc139c713, 32'h3d61a7af} /* (5, 6, 14) {real, imag} */,
  {32'hc0a7495f, 32'hc06f4ce0} /* (5, 6, 13) {real, imag} */,
  {32'h4010e7c2, 32'hc077d62a} /* (5, 6, 12) {real, imag} */,
  {32'h3f888182, 32'h410200af} /* (5, 6, 11) {real, imag} */,
  {32'hbfe109f4, 32'hc08484b1} /* (5, 6, 10) {real, imag} */,
  {32'hc097c033, 32'h40799482} /* (5, 6, 9) {real, imag} */,
  {32'hbf1e7162, 32'hc0bbe68d} /* (5, 6, 8) {real, imag} */,
  {32'h40182ea0, 32'h3f477673} /* (5, 6, 7) {real, imag} */,
  {32'hc10438bb, 32'h3f9ef9da} /* (5, 6, 6) {real, imag} */,
  {32'hc10e9611, 32'h400a270f} /* (5, 6, 5) {real, imag} */,
  {32'h400b6ba9, 32'hc118da98} /* (5, 6, 4) {real, imag} */,
  {32'h408c8bed, 32'h405d9219} /* (5, 6, 3) {real, imag} */,
  {32'hbf3372ef, 32'h3e2a11f2} /* (5, 6, 2) {real, imag} */,
  {32'hc13fd900, 32'h405c8b34} /* (5, 6, 1) {real, imag} */,
  {32'h40e9a601, 32'hc02dcd49} /* (5, 6, 0) {real, imag} */,
  {32'hbf0e9128, 32'hc0ea2645} /* (5, 5, 15) {real, imag} */,
  {32'hbf9774a6, 32'h412c7114} /* (5, 5, 14) {real, imag} */,
  {32'hc0501efd, 32'h411ad6c6} /* (5, 5, 13) {real, imag} */,
  {32'hc02fd0a6, 32'hc04a6f17} /* (5, 5, 12) {real, imag} */,
  {32'h3f64839e, 32'hc0d34a59} /* (5, 5, 11) {real, imag} */,
  {32'h40112cdc, 32'hc0b0278d} /* (5, 5, 10) {real, imag} */,
  {32'h3fa8fe07, 32'hc09457a3} /* (5, 5, 9) {real, imag} */,
  {32'hbb2bd2e5, 32'hc09f7f1a} /* (5, 5, 8) {real, imag} */,
  {32'hc0b324f5, 32'h3fb68a4a} /* (5, 5, 7) {real, imag} */,
  {32'hc0fe860d, 32'hc01e3ce3} /* (5, 5, 6) {real, imag} */,
  {32'h40d86de2, 32'hbf75315d} /* (5, 5, 5) {real, imag} */,
  {32'h40cd99ab, 32'hc0e12b05} /* (5, 5, 4) {real, imag} */,
  {32'hbfe564d0, 32'h40dc4322} /* (5, 5, 3) {real, imag} */,
  {32'hc0c263a2, 32'hc03f63a2} /* (5, 5, 2) {real, imag} */,
  {32'h412aa69b, 32'h405e9b15} /* (5, 5, 1) {real, imag} */,
  {32'hc0a04e9f, 32'hbebf80e7} /* (5, 5, 0) {real, imag} */,
  {32'hbec49070, 32'hc148c74a} /* (5, 4, 15) {real, imag} */,
  {32'h3f14940f, 32'hc02a81ec} /* (5, 4, 14) {real, imag} */,
  {32'h40345fa0, 32'hc0c6fe6e} /* (5, 4, 13) {real, imag} */,
  {32'h3f58eae4, 32'h408d3511} /* (5, 4, 12) {real, imag} */,
  {32'hc09ff3e9, 32'hc092ce8a} /* (5, 4, 11) {real, imag} */,
  {32'h4136c3cc, 32'h40263f62} /* (5, 4, 10) {real, imag} */,
  {32'h3fa863e3, 32'hc016ffae} /* (5, 4, 9) {real, imag} */,
  {32'hbf7654d3, 32'h3c4b4563} /* (5, 4, 8) {real, imag} */,
  {32'h409163c0, 32'h40dc1794} /* (5, 4, 7) {real, imag} */,
  {32'hbf94d24d, 32'hbd878350} /* (5, 4, 6) {real, imag} */,
  {32'h40a2159a, 32'hbeb65a2f} /* (5, 4, 5) {real, imag} */,
  {32'hc0d0e4fc, 32'hbdd33688} /* (5, 4, 4) {real, imag} */,
  {32'hbf409ff6, 32'hc09fd414} /* (5, 4, 3) {real, imag} */,
  {32'hc10294ac, 32'h40547d64} /* (5, 4, 2) {real, imag} */,
  {32'hc0ff5b38, 32'hc08118a2} /* (5, 4, 1) {real, imag} */,
  {32'hc0217bf6, 32'h3f8d81ba} /* (5, 4, 0) {real, imag} */,
  {32'h4082d4e2, 32'h4087fbf7} /* (5, 3, 15) {real, imag} */,
  {32'h3f65cc58, 32'hbddb704b} /* (5, 3, 14) {real, imag} */,
  {32'h40a9b4a1, 32'hc01715b2} /* (5, 3, 13) {real, imag} */,
  {32'h40e04968, 32'h3fdc6f4e} /* (5, 3, 12) {real, imag} */,
  {32'h412244cc, 32'h403304de} /* (5, 3, 11) {real, imag} */,
  {32'h4117b350, 32'hbf5a1f06} /* (5, 3, 10) {real, imag} */,
  {32'hc048b807, 32'h405fd6f6} /* (5, 3, 9) {real, imag} */,
  {32'hbee74252, 32'h407c03ef} /* (5, 3, 8) {real, imag} */,
  {32'hbfe3051e, 32'h400acb31} /* (5, 3, 7) {real, imag} */,
  {32'h409c5db5, 32'hbe31ab7f} /* (5, 3, 6) {real, imag} */,
  {32'hbfe0ef54, 32'hc14fd879} /* (5, 3, 5) {real, imag} */,
  {32'hc0b6a924, 32'h3fa875ef} /* (5, 3, 4) {real, imag} */,
  {32'h41071e5c, 32'h40e444fb} /* (5, 3, 3) {real, imag} */,
  {32'hbf48bb72, 32'h401c4ed5} /* (5, 3, 2) {real, imag} */,
  {32'hc0a9de95, 32'hbf04773c} /* (5, 3, 1) {real, imag} */,
  {32'h3ff10c26, 32'hc03c6c81} /* (5, 3, 0) {real, imag} */,
  {32'h40eb73a5, 32'h40b56247} /* (5, 2, 15) {real, imag} */,
  {32'hbfdb03de, 32'h40ca0af1} /* (5, 2, 14) {real, imag} */,
  {32'hc0ece269, 32'h40254d90} /* (5, 2, 13) {real, imag} */,
  {32'hc07712ed, 32'hc1334e83} /* (5, 2, 12) {real, imag} */,
  {32'h3fed8916, 32'h40ccc265} /* (5, 2, 11) {real, imag} */,
  {32'hc1167f26, 32'h4107406c} /* (5, 2, 10) {real, imag} */,
  {32'h3ed9b0e0, 32'hc0965d27} /* (5, 2, 9) {real, imag} */,
  {32'hbf43ed65, 32'hbdf29da4} /* (5, 2, 8) {real, imag} */,
  {32'hc09b92f6, 32'h3fada953} /* (5, 2, 7) {real, imag} */,
  {32'h403b2521, 32'hc0904956} /* (5, 2, 6) {real, imag} */,
  {32'hc0ae4c74, 32'h3f19cad3} /* (5, 2, 5) {real, imag} */,
  {32'hc0ccd9f6, 32'h40183a4f} /* (5, 2, 4) {real, imag} */,
  {32'h410a46f9, 32'hbef1ff30} /* (5, 2, 3) {real, imag} */,
  {32'h413825d3, 32'hc0a7d5d6} /* (5, 2, 2) {real, imag} */,
  {32'h415567aa, 32'hc09e2c1d} /* (5, 2, 1) {real, imag} */,
  {32'h3fcb00f7, 32'hbf4bcbf8} /* (5, 2, 0) {real, imag} */,
  {32'h41002885, 32'h4031b43c} /* (5, 1, 15) {real, imag} */,
  {32'hc162305a, 32'hc0fbbc02} /* (5, 1, 14) {real, imag} */,
  {32'h4074e298, 32'h404c31b4} /* (5, 1, 13) {real, imag} */,
  {32'h404595cc, 32'h41039a2b} /* (5, 1, 12) {real, imag} */,
  {32'hc0108e0e, 32'h40361d33} /* (5, 1, 11) {real, imag} */,
  {32'hbf7571e3, 32'hc0931eae} /* (5, 1, 10) {real, imag} */,
  {32'hc0be4b8e, 32'h40a1a1fa} /* (5, 1, 9) {real, imag} */,
  {32'hbfc968da, 32'h3f86304a} /* (5, 1, 8) {real, imag} */,
  {32'h3f92e928, 32'h3c84df57} /* (5, 1, 7) {real, imag} */,
  {32'h40b8ee23, 32'h406d587e} /* (5, 1, 6) {real, imag} */,
  {32'hbfb49d06, 32'hc1314697} /* (5, 1, 5) {real, imag} */,
  {32'h3ff49d29, 32'hbfdec1a5} /* (5, 1, 4) {real, imag} */,
  {32'hbff6f9be, 32'hc12defa8} /* (5, 1, 3) {real, imag} */,
  {32'h405bc194, 32'h41181ead} /* (5, 1, 2) {real, imag} */,
  {32'h406a695a, 32'hc02a22e1} /* (5, 1, 1) {real, imag} */,
  {32'h409d6d34, 32'h41025c39} /* (5, 1, 0) {real, imag} */,
  {32'hc07395a1, 32'h40a55cec} /* (5, 0, 15) {real, imag} */,
  {32'hc09b9369, 32'h40110a1b} /* (5, 0, 14) {real, imag} */,
  {32'hc0437b52, 32'h4031bb74} /* (5, 0, 13) {real, imag} */,
  {32'h40a10d96, 32'hbfff9b4f} /* (5, 0, 12) {real, imag} */,
  {32'hbfaa2128, 32'hc1586b54} /* (5, 0, 11) {real, imag} */,
  {32'hbf2860fa, 32'hc088569a} /* (5, 0, 10) {real, imag} */,
  {32'h4021485b, 32'hc0ad2af5} /* (5, 0, 9) {real, imag} */,
  {32'hbfc396e1, 32'hbd263c72} /* (5, 0, 8) {real, imag} */,
  {32'hc08deaec, 32'hbfbf8dda} /* (5, 0, 7) {real, imag} */,
  {32'h406258f2, 32'hc0899bc1} /* (5, 0, 6) {real, imag} */,
  {32'hc03f9a9e, 32'h40975821} /* (5, 0, 5) {real, imag} */,
  {32'h404cd604, 32'hc123382d} /* (5, 0, 4) {real, imag} */,
  {32'hc0580aa9, 32'hc06727ab} /* (5, 0, 3) {real, imag} */,
  {32'hc0adac02, 32'h3cf343c1} /* (5, 0, 2) {real, imag} */,
  {32'h400ec935, 32'hbf7390a3} /* (5, 0, 1) {real, imag} */,
  {32'h410516d2, 32'hc13222bc} /* (5, 0, 0) {real, imag} */,
  {32'h3f3effd0, 32'h405432d4} /* (4, 15, 15) {real, imag} */,
  {32'h40a78c59, 32'hbff970b9} /* (4, 15, 14) {real, imag} */,
  {32'hbea38287, 32'h3ebb89bd} /* (4, 15, 13) {real, imag} */,
  {32'h40ef9260, 32'hc0c8f8aa} /* (4, 15, 12) {real, imag} */,
  {32'hc085e830, 32'hbf87ab15} /* (4, 15, 11) {real, imag} */,
  {32'h3f405a77, 32'hc0c7e617} /* (4, 15, 10) {real, imag} */,
  {32'hbfde8912, 32'h4056b39d} /* (4, 15, 9) {real, imag} */,
  {32'hc04e39b8, 32'h406d3bec} /* (4, 15, 8) {real, imag} */,
  {32'h40bdfde9, 32'hbe9ee513} /* (4, 15, 7) {real, imag} */,
  {32'hc0208ffa, 32'hc013878f} /* (4, 15, 6) {real, imag} */,
  {32'hc0ea133a, 32'hc085f286} /* (4, 15, 5) {real, imag} */,
  {32'h3eb76200, 32'h40070ca2} /* (4, 15, 4) {real, imag} */,
  {32'hc0accb95, 32'hbf9c7c5b} /* (4, 15, 3) {real, imag} */,
  {32'hc14644eb, 32'hbf5b85af} /* (4, 15, 2) {real, imag} */,
  {32'h411eac5a, 32'hc123923e} /* (4, 15, 1) {real, imag} */,
  {32'h41b49cd3, 32'h415712b2} /* (4, 15, 0) {real, imag} */,
  {32'h4123b580, 32'hc02ec640} /* (4, 14, 15) {real, imag} */,
  {32'h410162a9, 32'h40b9f213} /* (4, 14, 14) {real, imag} */,
  {32'hc02c7e37, 32'h40d5630a} /* (4, 14, 13) {real, imag} */,
  {32'h3f74a3ff, 32'hbd696fe4} /* (4, 14, 12) {real, imag} */,
  {32'hc0af87a9, 32'h40c0f41c} /* (4, 14, 11) {real, imag} */,
  {32'h40c55617, 32'h40c85853} /* (4, 14, 10) {real, imag} */,
  {32'hc01b773d, 32'hc0c44475} /* (4, 14, 9) {real, imag} */,
  {32'hc0181c93, 32'hc0840e77} /* (4, 14, 8) {real, imag} */,
  {32'hc0efda8e, 32'h3fb7e5a1} /* (4, 14, 7) {real, imag} */,
  {32'h3fa70be7, 32'hc0f70abf} /* (4, 14, 6) {real, imag} */,
  {32'hc03c079c, 32'h40ba282e} /* (4, 14, 5) {real, imag} */,
  {32'hbe55a7f0, 32'hc1025359} /* (4, 14, 4) {real, imag} */,
  {32'hc039fa94, 32'h3fa40105} /* (4, 14, 3) {real, imag} */,
  {32'h4128a820, 32'h3fc9445a} /* (4, 14, 2) {real, imag} */,
  {32'hc1706c22, 32'hc0be7fd2} /* (4, 14, 1) {real, imag} */,
  {32'hc0bb6c3f, 32'hc17f07f4} /* (4, 14, 0) {real, imag} */,
  {32'hc09f6713, 32'h3db3eee1} /* (4, 13, 15) {real, imag} */,
  {32'hc0688499, 32'h40f23a05} /* (4, 13, 14) {real, imag} */,
  {32'hc05d5d4c, 32'hc0928ed1} /* (4, 13, 13) {real, imag} */,
  {32'hc0b09723, 32'h401d4549} /* (4, 13, 12) {real, imag} */,
  {32'hc08137dd, 32'h403f85de} /* (4, 13, 11) {real, imag} */,
  {32'h411f938f, 32'hc0aedd1d} /* (4, 13, 10) {real, imag} */,
  {32'hc0bc8dfe, 32'h411c1fbf} /* (4, 13, 9) {real, imag} */,
  {32'hc09fd0d4, 32'hbf10f477} /* (4, 13, 8) {real, imag} */,
  {32'hbf93e6a3, 32'h40d727ec} /* (4, 13, 7) {real, imag} */,
  {32'hc028d546, 32'h40841ab9} /* (4, 13, 6) {real, imag} */,
  {32'h406b6c04, 32'hc12a73cd} /* (4, 13, 5) {real, imag} */,
  {32'h40550532, 32'hbed76676} /* (4, 13, 4) {real, imag} */,
  {32'hbeda50f9, 32'h40095ce8} /* (4, 13, 3) {real, imag} */,
  {32'h40641d61, 32'h4020e8f7} /* (4, 13, 2) {real, imag} */,
  {32'hc099a64c, 32'hc082d468} /* (4, 13, 1) {real, imag} */,
  {32'h4046d5dd, 32'h3f9def25} /* (4, 13, 0) {real, imag} */,
  {32'hbef7055e, 32'hbf95d681} /* (4, 12, 15) {real, imag} */,
  {32'hc0225711, 32'hc1025d6a} /* (4, 12, 14) {real, imag} */,
  {32'h4006ed3b, 32'hbf7b4046} /* (4, 12, 13) {real, imag} */,
  {32'hc1781de9, 32'h3e14c422} /* (4, 12, 12) {real, imag} */,
  {32'h404d8202, 32'hbf8b5d2c} /* (4, 12, 11) {real, imag} */,
  {32'hbe8122f3, 32'hbf905af1} /* (4, 12, 10) {real, imag} */,
  {32'h409f7b31, 32'h40c2278e} /* (4, 12, 9) {real, imag} */,
  {32'h40aa5658, 32'h3fc82d1f} /* (4, 12, 8) {real, imag} */,
  {32'hbf3c7360, 32'hc0a01d0e} /* (4, 12, 7) {real, imag} */,
  {32'h411f013c, 32'h40b07849} /* (4, 12, 6) {real, imag} */,
  {32'h407ff0ff, 32'h4074cda8} /* (4, 12, 5) {real, imag} */,
  {32'h3eedd483, 32'h40134704} /* (4, 12, 4) {real, imag} */,
  {32'h4059edbc, 32'h40a75371} /* (4, 12, 3) {real, imag} */,
  {32'hc10c3286, 32'h409cb6f2} /* (4, 12, 2) {real, imag} */,
  {32'h40ba0f28, 32'h40c7bce7} /* (4, 12, 1) {real, imag} */,
  {32'hbfe1f851, 32'h408d263d} /* (4, 12, 0) {real, imag} */,
  {32'hc16b65cb, 32'hc10c76eb} /* (4, 11, 15) {real, imag} */,
  {32'hbf08b9c4, 32'hc0f5845e} /* (4, 11, 14) {real, imag} */,
  {32'hc0ff1239, 32'h406314e5} /* (4, 11, 13) {real, imag} */,
  {32'h40a8db77, 32'h40f18ae0} /* (4, 11, 12) {real, imag} */,
  {32'h3f4ac918, 32'hc09f6531} /* (4, 11, 11) {real, imag} */,
  {32'h3f6663e9, 32'h4059922b} /* (4, 11, 10) {real, imag} */,
  {32'hc0d7d0ae, 32'hbeef032e} /* (4, 11, 9) {real, imag} */,
  {32'h3f5c5b55, 32'h4092b50c} /* (4, 11, 8) {real, imag} */,
  {32'hbfc29454, 32'h3f4847aa} /* (4, 11, 7) {real, imag} */,
  {32'hc0eb1962, 32'hc01733f8} /* (4, 11, 6) {real, imag} */,
  {32'h3feb6c61, 32'h402e0221} /* (4, 11, 5) {real, imag} */,
  {32'h40963d83, 32'hc053d8ca} /* (4, 11, 4) {real, imag} */,
  {32'h3f8934b3, 32'hbf49c05b} /* (4, 11, 3) {real, imag} */,
  {32'h4054e032, 32'h40a2325b} /* (4, 11, 2) {real, imag} */,
  {32'hc0eb0c47, 32'hbb365898} /* (4, 11, 1) {real, imag} */,
  {32'hc0c4b502, 32'h4101c0ad} /* (4, 11, 0) {real, imag} */,
  {32'hc149af2e, 32'h3f58aada} /* (4, 10, 15) {real, imag} */,
  {32'h415ae054, 32'hc0252f59} /* (4, 10, 14) {real, imag} */,
  {32'h4064a9fc, 32'hbe37b243} /* (4, 10, 13) {real, imag} */,
  {32'hc08b06f0, 32'h40831b1e} /* (4, 10, 12) {real, imag} */,
  {32'hc06c0b76, 32'h404cbd92} /* (4, 10, 11) {real, imag} */,
  {32'hc128819f, 32'hc00d8a0e} /* (4, 10, 10) {real, imag} */,
  {32'h3f8d1502, 32'h3ffad29a} /* (4, 10, 9) {real, imag} */,
  {32'hbfa39fc0, 32'hc065c839} /* (4, 10, 8) {real, imag} */,
  {32'hbfec99e0, 32'h3fa3c271} /* (4, 10, 7) {real, imag} */,
  {32'hc09cea2b, 32'h3fd9f200} /* (4, 10, 6) {real, imag} */,
  {32'h411b36d4, 32'hc0d1b3f1} /* (4, 10, 5) {real, imag} */,
  {32'h401c7126, 32'hc0baf6fb} /* (4, 10, 4) {real, imag} */,
  {32'h40e59d2e, 32'h3f71bae1} /* (4, 10, 3) {real, imag} */,
  {32'h4023bdf6, 32'h412fbd85} /* (4, 10, 2) {real, imag} */,
  {32'h40917842, 32'h4074a5ee} /* (4, 10, 1) {real, imag} */,
  {32'hc004c443, 32'hc02c14c0} /* (4, 10, 0) {real, imag} */,
  {32'h40553337, 32'hbf9ee217} /* (4, 9, 15) {real, imag} */,
  {32'hc001d18d, 32'h40668a33} /* (4, 9, 14) {real, imag} */,
  {32'hc08dc826, 32'hbf17e050} /* (4, 9, 13) {real, imag} */,
  {32'h4044dded, 32'h40011e57} /* (4, 9, 12) {real, imag} */,
  {32'h409751f0, 32'hbff8eedb} /* (4, 9, 11) {real, imag} */,
  {32'hbff73308, 32'h40eeba0f} /* (4, 9, 10) {real, imag} */,
  {32'hbee2b952, 32'hbd53c2e3} /* (4, 9, 9) {real, imag} */,
  {32'h3fa2f7c1, 32'h407aec84} /* (4, 9, 8) {real, imag} */,
  {32'hbfcf93d2, 32'h3f8b9aac} /* (4, 9, 7) {real, imag} */,
  {32'h407e81b3, 32'hc119a977} /* (4, 9, 6) {real, imag} */,
  {32'hbfe46f45, 32'h404a8c5c} /* (4, 9, 5) {real, imag} */,
  {32'hc00f7bb6, 32'hbd5118a5} /* (4, 9, 4) {real, imag} */,
  {32'hbea7f3dc, 32'hc023d62a} /* (4, 9, 3) {real, imag} */,
  {32'h405b57c7, 32'hc0370c66} /* (4, 9, 2) {real, imag} */,
  {32'hc1300528, 32'h40519843} /* (4, 9, 1) {real, imag} */,
  {32'h3cad9d20, 32'hbfc58c74} /* (4, 9, 0) {real, imag} */,
  {32'h40d6081b, 32'h3e23cbda} /* (4, 8, 15) {real, imag} */,
  {32'hc026fe1d, 32'h3e63ce1a} /* (4, 8, 14) {real, imag} */,
  {32'hbf5509ba, 32'hbfaad099} /* (4, 8, 13) {real, imag} */,
  {32'hc06ee6b0, 32'h40e1e6f6} /* (4, 8, 12) {real, imag} */,
  {32'hbfdc28ec, 32'h405f550c} /* (4, 8, 11) {real, imag} */,
  {32'h41264451, 32'h40a60dd5} /* (4, 8, 10) {real, imag} */,
  {32'h3f193052, 32'hc03336a9} /* (4, 8, 9) {real, imag} */,
  {32'hc04a6665, 32'h401353a1} /* (4, 8, 8) {real, imag} */,
  {32'hbf41b754, 32'h3e9da841} /* (4, 8, 7) {real, imag} */,
  {32'h40ebff79, 32'h408d38fd} /* (4, 8, 6) {real, imag} */,
  {32'hc0bc4ead, 32'hc0a88f17} /* (4, 8, 5) {real, imag} */,
  {32'h4032bcd2, 32'hbf7fa7a6} /* (4, 8, 4) {real, imag} */,
  {32'hbf717e49, 32'h403b7886} /* (4, 8, 3) {real, imag} */,
  {32'h404aece7, 32'hc05764a8} /* (4, 8, 2) {real, imag} */,
  {32'h406002ad, 32'hbf1bf36c} /* (4, 8, 1) {real, imag} */,
  {32'hc0bb3ab9, 32'h3f826da2} /* (4, 8, 0) {real, imag} */,
  {32'hbecd39f8, 32'h40d3b745} /* (4, 7, 15) {real, imag} */,
  {32'hc0914026, 32'h405d6458} /* (4, 7, 14) {real, imag} */,
  {32'h4045d73e, 32'hbf602a10} /* (4, 7, 13) {real, imag} */,
  {32'hc151c892, 32'hbe1ff026} /* (4, 7, 12) {real, imag} */,
  {32'hbf82ac79, 32'h3f84d7c7} /* (4, 7, 11) {real, imag} */,
  {32'h3f0f759d, 32'hc0b7f154} /* (4, 7, 10) {real, imag} */,
  {32'h40e43883, 32'h40442a7b} /* (4, 7, 9) {real, imag} */,
  {32'h3feec3ba, 32'h3f2e2ba9} /* (4, 7, 8) {real, imag} */,
  {32'hbfb520d2, 32'h407fb937} /* (4, 7, 7) {real, imag} */,
  {32'hc127d04b, 32'h407c6b0f} /* (4, 7, 6) {real, imag} */,
  {32'h40b6b4f3, 32'hc04a73eb} /* (4, 7, 5) {real, imag} */,
  {32'hbf5d5b3b, 32'h4083ba4f} /* (4, 7, 4) {real, imag} */,
  {32'hbff8deea, 32'h406ca059} /* (4, 7, 3) {real, imag} */,
  {32'h40ac21e5, 32'h3fc0f621} /* (4, 7, 2) {real, imag} */,
  {32'h3fdeab87, 32'hc0c16ea8} /* (4, 7, 1) {real, imag} */,
  {32'h3fde0eba, 32'hc105c267} /* (4, 7, 0) {real, imag} */,
  {32'hbf9245c6, 32'h4162144a} /* (4, 6, 15) {real, imag} */,
  {32'hbf1cee19, 32'hc0965762} /* (4, 6, 14) {real, imag} */,
  {32'hbf03fbc1, 32'h3f372b57} /* (4, 6, 13) {real, imag} */,
  {32'hc12450f2, 32'hc0466804} /* (4, 6, 12) {real, imag} */,
  {32'hc00119a0, 32'hbfe104dd} /* (4, 6, 11) {real, imag} */,
  {32'h402797bf, 32'h3f0adb9c} /* (4, 6, 10) {real, imag} */,
  {32'hc07ec43d, 32'hc104a325} /* (4, 6, 9) {real, imag} */,
  {32'h40beba6b, 32'h406c6f5c} /* (4, 6, 8) {real, imag} */,
  {32'hbfc34536, 32'hbd2735be} /* (4, 6, 7) {real, imag} */,
  {32'h40b26166, 32'h4020f0ec} /* (4, 6, 6) {real, imag} */,
  {32'hc05f3abf, 32'h4099c131} /* (4, 6, 5) {real, imag} */,
  {32'h4106237c, 32'h415de5db} /* (4, 6, 4) {real, imag} */,
  {32'hc08fc80e, 32'hc10ed02e} /* (4, 6, 3) {real, imag} */,
  {32'h411357af, 32'hc05c4569} /* (4, 6, 2) {real, imag} */,
  {32'hbf48c932, 32'hc10fd874} /* (4, 6, 1) {real, imag} */,
  {32'hc0b394b5, 32'h415263cf} /* (4, 6, 0) {real, imag} */,
  {32'hc170194a, 32'h407d05f9} /* (4, 5, 15) {real, imag} */,
  {32'hc00faf28, 32'hc0ca6d71} /* (4, 5, 14) {real, imag} */,
  {32'hc02225c2, 32'hc0d1c1db} /* (4, 5, 13) {real, imag} */,
  {32'h40402017, 32'hc0c57d01} /* (4, 5, 12) {real, imag} */,
  {32'hc12f8c24, 32'h3fb38bcf} /* (4, 5, 11) {real, imag} */,
  {32'hc0421138, 32'hc10c7ad3} /* (4, 5, 10) {real, imag} */,
  {32'h40ad004b, 32'hbfc21685} /* (4, 5, 9) {real, imag} */,
  {32'h404dab87, 32'h4060e9c1} /* (4, 5, 8) {real, imag} */,
  {32'h40b5f5ac, 32'h3fe37f5e} /* (4, 5, 7) {real, imag} */,
  {32'h40207a74, 32'h401d251f} /* (4, 5, 6) {real, imag} */,
  {32'h40d6ebfc, 32'hc0edf348} /* (4, 5, 5) {real, imag} */,
  {32'h403706b9, 32'h40bc2daf} /* (4, 5, 4) {real, imag} */,
  {32'hc1598ee7, 32'h416729ae} /* (4, 5, 3) {real, imag} */,
  {32'hbde1c001, 32'hc0ab5568} /* (4, 5, 2) {real, imag} */,
  {32'h3ea1056b, 32'h40b15b09} /* (4, 5, 1) {real, imag} */,
  {32'hbd802de5, 32'h3fe57e79} /* (4, 5, 0) {real, imag} */,
  {32'h41249b5e, 32'hc06a3393} /* (4, 4, 15) {real, imag} */,
  {32'h405396a3, 32'h4092dce8} /* (4, 4, 14) {real, imag} */,
  {32'hc028cd08, 32'h41129296} /* (4, 4, 13) {real, imag} */,
  {32'h4082e17d, 32'h407f8c39} /* (4, 4, 12) {real, imag} */,
  {32'h3f82b094, 32'h409d4efa} /* (4, 4, 11) {real, imag} */,
  {32'hc173743b, 32'hc098905e} /* (4, 4, 10) {real, imag} */,
  {32'hbe14dbf8, 32'h411e2092} /* (4, 4, 9) {real, imag} */,
  {32'h40502110, 32'hbc7e881f} /* (4, 4, 8) {real, imag} */,
  {32'h4053c391, 32'hc018b5d3} /* (4, 4, 7) {real, imag} */,
  {32'h40163af5, 32'hc0c3edb9} /* (4, 4, 6) {real, imag} */,
  {32'h40e36815, 32'h3ee8dc0a} /* (4, 4, 5) {real, imag} */,
  {32'h4073f26c, 32'h3f1c6210} /* (4, 4, 4) {real, imag} */,
  {32'hc0a8dd8e, 32'hc073b27b} /* (4, 4, 3) {real, imag} */,
  {32'hc00e9eb3, 32'h408021ed} /* (4, 4, 2) {real, imag} */,
  {32'h4084893f, 32'h4014fc4b} /* (4, 4, 1) {real, imag} */,
  {32'h409930ee, 32'h4000c00a} /* (4, 4, 0) {real, imag} */,
  {32'hc0dd0425, 32'h4015ce32} /* (4, 3, 15) {real, imag} */,
  {32'h3fa8b7d6, 32'hbfec6341} /* (4, 3, 14) {real, imag} */,
  {32'hc09d302a, 32'hc0a589ce} /* (4, 3, 13) {real, imag} */,
  {32'hc0426572, 32'hc07f93ab} /* (4, 3, 12) {real, imag} */,
  {32'h409c9222, 32'h406265c5} /* (4, 3, 11) {real, imag} */,
  {32'h40f3c561, 32'hc0ee8d46} /* (4, 3, 10) {real, imag} */,
  {32'h4094c30c, 32'h3f8f7eab} /* (4, 3, 9) {real, imag} */,
  {32'h4043d872, 32'hbf0d72e8} /* (4, 3, 8) {real, imag} */,
  {32'hc012a630, 32'h40b5dfb6} /* (4, 3, 7) {real, imag} */,
  {32'h40e82b87, 32'h3f89771f} /* (4, 3, 6) {real, imag} */,
  {32'h4118eb86, 32'h40f3b68e} /* (4, 3, 5) {real, imag} */,
  {32'hc1276831, 32'h404efd52} /* (4, 3, 4) {real, imag} */,
  {32'hbe46ca70, 32'hc085d0f6} /* (4, 3, 3) {real, imag} */,
  {32'h4055943c, 32'h404a858c} /* (4, 3, 2) {real, imag} */,
  {32'hc00a594b, 32'h40d74b8d} /* (4, 3, 1) {real, imag} */,
  {32'h4079fb3a, 32'h3fb731a9} /* (4, 3, 0) {real, imag} */,
  {32'h40a41d99, 32'h40fb52d9} /* (4, 2, 15) {real, imag} */,
  {32'hc00eed5d, 32'hc1171dc9} /* (4, 2, 14) {real, imag} */,
  {32'h413487d1, 32'h40a03e53} /* (4, 2, 13) {real, imag} */,
  {32'h3fc4af1a, 32'h4081436c} /* (4, 2, 12) {real, imag} */,
  {32'h40b05a00, 32'h40346391} /* (4, 2, 11) {real, imag} */,
  {32'hbeddd4fc, 32'hbfee4509} /* (4, 2, 10) {real, imag} */,
  {32'hbf64a094, 32'h3fa6876f} /* (4, 2, 9) {real, imag} */,
  {32'h40e3fd98, 32'h3fb7934c} /* (4, 2, 8) {real, imag} */,
  {32'hc093cd77, 32'hbfc7280f} /* (4, 2, 7) {real, imag} */,
  {32'h40f9282c, 32'h40cb8cc5} /* (4, 2, 6) {real, imag} */,
  {32'hbf95a8cf, 32'hc0607e30} /* (4, 2, 5) {real, imag} */,
  {32'hbf70fcee, 32'hc102bd59} /* (4, 2, 4) {real, imag} */,
  {32'h40b081ef, 32'hc09a82b1} /* (4, 2, 3) {real, imag} */,
  {32'h405ec1b6, 32'hc05ce535} /* (4, 2, 2) {real, imag} */,
  {32'h4030c5d2, 32'h40528983} /* (4, 2, 1) {real, imag} */,
  {32'hc12baba7, 32'hc0d9c1e4} /* (4, 2, 0) {real, imag} */,
  {32'h3e0e403e, 32'h417e5fe9} /* (4, 1, 15) {real, imag} */,
  {32'hc0efc3d8, 32'h3f9daba5} /* (4, 1, 14) {real, imag} */,
  {32'hc0993e60, 32'hc1325d64} /* (4, 1, 13) {real, imag} */,
  {32'h3fe8c785, 32'hc0e545f1} /* (4, 1, 12) {real, imag} */,
  {32'hc074643f, 32'hbe628677} /* (4, 1, 11) {real, imag} */,
  {32'h4074f888, 32'h41053dc1} /* (4, 1, 10) {real, imag} */,
  {32'h3fc6afc5, 32'hbf19db58} /* (4, 1, 9) {real, imag} */,
  {32'hc06e501c, 32'h3fbb5d84} /* (4, 1, 8) {real, imag} */,
  {32'hbf790f31, 32'h3f7a4538} /* (4, 1, 7) {real, imag} */,
  {32'hc037db01, 32'hbe3abca9} /* (4, 1, 6) {real, imag} */,
  {32'hc0a089b1, 32'h408afeee} /* (4, 1, 5) {real, imag} */,
  {32'h403f5101, 32'h3f17386a} /* (4, 1, 4) {real, imag} */,
  {32'hc02b52a1, 32'h410dcf84} /* (4, 1, 3) {real, imag} */,
  {32'h410fc737, 32'h3e807443} /* (4, 1, 2) {real, imag} */,
  {32'hc0e932b1, 32'h40aa44c0} /* (4, 1, 1) {real, imag} */,
  {32'hc06d1897, 32'hc00b483b} /* (4, 1, 0) {real, imag} */,
  {32'hc1525390, 32'hc05b795c} /* (4, 0, 15) {real, imag} */,
  {32'hc11c76bc, 32'hc01b958b} /* (4, 0, 14) {real, imag} */,
  {32'h40f4f089, 32'h4134f737} /* (4, 0, 13) {real, imag} */,
  {32'h407aecb7, 32'h403c805b} /* (4, 0, 12) {real, imag} */,
  {32'h40a49e35, 32'hc0efd47b} /* (4, 0, 11) {real, imag} */,
  {32'hc017d6bd, 32'hbf3096e4} /* (4, 0, 10) {real, imag} */,
  {32'h40a9fc38, 32'hbffd70a0} /* (4, 0, 9) {real, imag} */,
  {32'hbefcd082, 32'hbf07f3ed} /* (4, 0, 8) {real, imag} */,
  {32'hbfab6815, 32'hc06e3bbb} /* (4, 0, 7) {real, imag} */,
  {32'hc071f363, 32'hbee508da} /* (4, 0, 6) {real, imag} */,
  {32'hbf8abf98, 32'h4124a1dc} /* (4, 0, 5) {real, imag} */,
  {32'hc0d777a2, 32'hc1078757} /* (4, 0, 4) {real, imag} */,
  {32'h3f8cc2c5, 32'hc0b7cb53} /* (4, 0, 3) {real, imag} */,
  {32'hc0179f0f, 32'hbed144bf} /* (4, 0, 2) {real, imag} */,
  {32'h3e3a7b45, 32'hc12710ed} /* (4, 0, 1) {real, imag} */,
  {32'hc0b6046b, 32'h3f4872f1} /* (4, 0, 0) {real, imag} */,
  {32'h3fcebb0e, 32'h3f5b732f} /* (3, 15, 15) {real, imag} */,
  {32'hc18512af, 32'hc0dc2428} /* (3, 15, 14) {real, imag} */,
  {32'h40a47e77, 32'h40c4b74e} /* (3, 15, 13) {real, imag} */,
  {32'h3f6ee909, 32'h41374b37} /* (3, 15, 12) {real, imag} */,
  {32'h40b92e08, 32'h413e5efe} /* (3, 15, 11) {real, imag} */,
  {32'h41109528, 32'h40b7f3bf} /* (3, 15, 10) {real, imag} */,
  {32'h3f5478f5, 32'hc016478f} /* (3, 15, 9) {real, imag} */,
  {32'hc01fdfc3, 32'h3fcb49dc} /* (3, 15, 8) {real, imag} */,
  {32'hc048a66d, 32'h40244f47} /* (3, 15, 7) {real, imag} */,
  {32'hc00dfe53, 32'h40dec1cd} /* (3, 15, 6) {real, imag} */,
  {32'h40babda3, 32'hc15b25a8} /* (3, 15, 5) {real, imag} */,
  {32'h40cadd20, 32'h3d38b123} /* (3, 15, 4) {real, imag} */,
  {32'hc0a23499, 32'hc0ed8f71} /* (3, 15, 3) {real, imag} */,
  {32'hc01a3ac1, 32'h40be817f} /* (3, 15, 2) {real, imag} */,
  {32'hc18f4955, 32'hc106844e} /* (3, 15, 1) {real, imag} */,
  {32'h40afa5cd, 32'hc0568109} /* (3, 15, 0) {real, imag} */,
  {32'h4067553f, 32'hc1153fef} /* (3, 14, 15) {real, imag} */,
  {32'hc108b1c8, 32'hc06b6835} /* (3, 14, 14) {real, imag} */,
  {32'h3f90bf40, 32'hc11ee0ec} /* (3, 14, 13) {real, imag} */,
  {32'hbccfd9ff, 32'h40d23980} /* (3, 14, 12) {real, imag} */,
  {32'h3f3d068d, 32'hc01b332f} /* (3, 14, 11) {real, imag} */,
  {32'hc03dc734, 32'hbe7efe97} /* (3, 14, 10) {real, imag} */,
  {32'h3d33c78e, 32'h3fee92a3} /* (3, 14, 9) {real, imag} */,
  {32'hc01a9e68, 32'hc08247a5} /* (3, 14, 8) {real, imag} */,
  {32'hc0ce2ce8, 32'hc0ba90a8} /* (3, 14, 7) {real, imag} */,
  {32'hc12cee8a, 32'h40098fa1} /* (3, 14, 6) {real, imag} */,
  {32'h409b8671, 32'h3fe1774b} /* (3, 14, 5) {real, imag} */,
  {32'h40983997, 32'h3eb2b301} /* (3, 14, 4) {real, imag} */,
  {32'h3e4f19d7, 32'h40976fa3} /* (3, 14, 3) {real, imag} */,
  {32'hc08f4a3f, 32'hbf11eb9a} /* (3, 14, 2) {real, imag} */,
  {32'hc064695f, 32'hbf36361d} /* (3, 14, 1) {real, imag} */,
  {32'h410565ac, 32'h401870c9} /* (3, 14, 0) {real, imag} */,
  {32'hc0a68d4a, 32'h4093d175} /* (3, 13, 15) {real, imag} */,
  {32'hc0865bea, 32'hc0f0bbfe} /* (3, 13, 14) {real, imag} */,
  {32'h41170ee1, 32'h40b06c79} /* (3, 13, 13) {real, imag} */,
  {32'h4183b1f9, 32'hc0b77d9d} /* (3, 13, 12) {real, imag} */,
  {32'hc094859f, 32'hc093d643} /* (3, 13, 11) {real, imag} */,
  {32'h3fdb58b4, 32'h400bef70} /* (3, 13, 10) {real, imag} */,
  {32'h403034c4, 32'h401e185c} /* (3, 13, 9) {real, imag} */,
  {32'h410305d8, 32'hbf27347a} /* (3, 13, 8) {real, imag} */,
  {32'h3ff176f6, 32'hbfab3c40} /* (3, 13, 7) {real, imag} */,
  {32'h4112cf9d, 32'h40b4cde1} /* (3, 13, 6) {real, imag} */,
  {32'h40b0071a, 32'h4019c010} /* (3, 13, 5) {real, imag} */,
  {32'hbe3dd80c, 32'h401bebac} /* (3, 13, 4) {real, imag} */,
  {32'h40046fcd, 32'hc102b5d9} /* (3, 13, 3) {real, imag} */,
  {32'hc10e7ea2, 32'hc01e27f7} /* (3, 13, 2) {real, imag} */,
  {32'h40cabf61, 32'hbfb94b3f} /* (3, 13, 1) {real, imag} */,
  {32'hc0fa605a, 32'h3e373c99} /* (3, 13, 0) {real, imag} */,
  {32'h40e1b520, 32'h3f7f6a88} /* (3, 12, 15) {real, imag} */,
  {32'hbf1b5009, 32'h40521288} /* (3, 12, 14) {real, imag} */,
  {32'h40c5fe03, 32'hc0a276a8} /* (3, 12, 13) {real, imag} */,
  {32'hbec3b00d, 32'h3f93e289} /* (3, 12, 12) {real, imag} */,
  {32'hc0e32e40, 32'hc11f6120} /* (3, 12, 11) {real, imag} */,
  {32'hc0e600fd, 32'h4046430d} /* (3, 12, 10) {real, imag} */,
  {32'h4107ecf5, 32'hbfd9e0c0} /* (3, 12, 9) {real, imag} */,
  {32'hbee19fd7, 32'hc08b1196} /* (3, 12, 8) {real, imag} */,
  {32'hbf946963, 32'h3f4cd93b} /* (3, 12, 7) {real, imag} */,
  {32'hc125cb36, 32'h40d7ae6c} /* (3, 12, 6) {real, imag} */,
  {32'h3dcb041b, 32'h40c0d862} /* (3, 12, 5) {real, imag} */,
  {32'hc127348c, 32'hbe4f7ad2} /* (3, 12, 4) {real, imag} */,
  {32'h4123ce63, 32'h3fb536d0} /* (3, 12, 3) {real, imag} */,
  {32'h402c0509, 32'h3f9c6fba} /* (3, 12, 2) {real, imag} */,
  {32'h401e4f54, 32'hc1709db4} /* (3, 12, 1) {real, imag} */,
  {32'hc005b869, 32'h3fa77930} /* (3, 12, 0) {real, imag} */,
  {32'hc0ad6570, 32'h40d160cd} /* (3, 11, 15) {real, imag} */,
  {32'h413c9d40, 32'h40529213} /* (3, 11, 14) {real, imag} */,
  {32'hbec8c493, 32'h3eebdef8} /* (3, 11, 13) {real, imag} */,
  {32'hc0cf7c72, 32'hc09fcaa3} /* (3, 11, 12) {real, imag} */,
  {32'hbfefc6da, 32'h40758d08} /* (3, 11, 11) {real, imag} */,
  {32'h3f027575, 32'hc0f549ae} /* (3, 11, 10) {real, imag} */,
  {32'hc0fa7d30, 32'h40b36edb} /* (3, 11, 9) {real, imag} */,
  {32'h3de34415, 32'hbf95eaea} /* (3, 11, 8) {real, imag} */,
  {32'h40c50664, 32'hc09e092b} /* (3, 11, 7) {real, imag} */,
  {32'h40f77f0d, 32'hc08529c1} /* (3, 11, 6) {real, imag} */,
  {32'h40102f8c, 32'hc108f8d9} /* (3, 11, 5) {real, imag} */,
  {32'hc08a431a, 32'hbe80e5aa} /* (3, 11, 4) {real, imag} */,
  {32'hc0dac0eb, 32'hc0013127} /* (3, 11, 3) {real, imag} */,
  {32'h3daf42b8, 32'h4091b8cd} /* (3, 11, 2) {real, imag} */,
  {32'h411d40f9, 32'h410689b8} /* (3, 11, 1) {real, imag} */,
  {32'hc0a20fdc, 32'h3f465326} /* (3, 11, 0) {real, imag} */,
  {32'hc053ea6a, 32'hc06dc09b} /* (3, 10, 15) {real, imag} */,
  {32'h3e7570bc, 32'hc0892b7b} /* (3, 10, 14) {real, imag} */,
  {32'hbfdf99e1, 32'h411e7909} /* (3, 10, 13) {real, imag} */,
  {32'hc0c34141, 32'hc07aa1b3} /* (3, 10, 12) {real, imag} */,
  {32'hc014e170, 32'h408c07cd} /* (3, 10, 11) {real, imag} */,
  {32'hc0769945, 32'hc10428b4} /* (3, 10, 10) {real, imag} */,
  {32'h402994b7, 32'hbed31afd} /* (3, 10, 9) {real, imag} */,
  {32'hbff35e8b, 32'hbf4dd9f7} /* (3, 10, 8) {real, imag} */,
  {32'h3f1a4b39, 32'hc117e1ce} /* (3, 10, 7) {real, imag} */,
  {32'h40b480d5, 32'hbfb2dde8} /* (3, 10, 6) {real, imag} */,
  {32'hc090cb8d, 32'h40caf30e} /* (3, 10, 5) {real, imag} */,
  {32'hbff9a097, 32'hc008c207} /* (3, 10, 4) {real, imag} */,
  {32'h3eb243f7, 32'h411472fc} /* (3, 10, 3) {real, imag} */,
  {32'h405dfe67, 32'h40e8a374} /* (3, 10, 2) {real, imag} */,
  {32'hbff1ec04, 32'h4099db5c} /* (3, 10, 1) {real, imag} */,
  {32'h3e3b1d3a, 32'h40156d47} /* (3, 10, 0) {real, imag} */,
  {32'h3fa99d43, 32'h409f6b97} /* (3, 9, 15) {real, imag} */,
  {32'h40635030, 32'h403f0e12} /* (3, 9, 14) {real, imag} */,
  {32'h409e535c, 32'h3e003e7c} /* (3, 9, 13) {real, imag} */,
  {32'hbf914ba5, 32'hc07d706e} /* (3, 9, 12) {real, imag} */,
  {32'hbfef949a, 32'hc02dd992} /* (3, 9, 11) {real, imag} */,
  {32'h402752a7, 32'h404cc238} /* (3, 9, 10) {real, imag} */,
  {32'hbf02f407, 32'hc0ddfe11} /* (3, 9, 9) {real, imag} */,
  {32'hbfbc8ce5, 32'h403f027e} /* (3, 9, 8) {real, imag} */,
  {32'hbf25f186, 32'h4095a269} /* (3, 9, 7) {real, imag} */,
  {32'h3f85a97c, 32'h410597a8} /* (3, 9, 6) {real, imag} */,
  {32'h40f9caf8, 32'h4048366e} /* (3, 9, 5) {real, imag} */,
  {32'hbfa95b6e, 32'h409128dc} /* (3, 9, 4) {real, imag} */,
  {32'hc05c660c, 32'hc0d6150c} /* (3, 9, 3) {real, imag} */,
  {32'hc07f5764, 32'hc06b6262} /* (3, 9, 2) {real, imag} */,
  {32'h40013783, 32'hc0421f63} /* (3, 9, 1) {real, imag} */,
  {32'hc08cf8dd, 32'hbf407e88} /* (3, 9, 0) {real, imag} */,
  {32'h40204646, 32'h402f0a2a} /* (3, 8, 15) {real, imag} */,
  {32'hbf6ad8b4, 32'h3ea3daf3} /* (3, 8, 14) {real, imag} */,
  {32'hbf13f980, 32'h40077ef2} /* (3, 8, 13) {real, imag} */,
  {32'h3fa6788e, 32'h3eb0d96f} /* (3, 8, 12) {real, imag} */,
  {32'hc0d5e0c2, 32'hc07d7bbc} /* (3, 8, 11) {real, imag} */,
  {32'h4063fd5c, 32'hc0764f28} /* (3, 8, 10) {real, imag} */,
  {32'h40d0e74e, 32'hc112cb63} /* (3, 8, 9) {real, imag} */,
  {32'hc065abe1, 32'hbe9dd167} /* (3, 8, 8) {real, imag} */,
  {32'h401dd922, 32'h3f0f4c43} /* (3, 8, 7) {real, imag} */,
  {32'hc0394820, 32'h3f34e83c} /* (3, 8, 6) {real, imag} */,
  {32'h3ffa0eb6, 32'hbf3bfd0c} /* (3, 8, 5) {real, imag} */,
  {32'h408ce177, 32'h401837d0} /* (3, 8, 4) {real, imag} */,
  {32'h40211c30, 32'h40b44a42} /* (3, 8, 3) {real, imag} */,
  {32'hbf9c24f7, 32'hc04f9548} /* (3, 8, 2) {real, imag} */,
  {32'hbfdc52a0, 32'hbfc9fd44} /* (3, 8, 1) {real, imag} */,
  {32'h3f263e4e, 32'hbfd33e7e} /* (3, 8, 0) {real, imag} */,
  {32'hbf923c8f, 32'hc097a4c2} /* (3, 7, 15) {real, imag} */,
  {32'h410248c1, 32'h3fe5b85a} /* (3, 7, 14) {real, imag} */,
  {32'h407729fe, 32'h406c9928} /* (3, 7, 13) {real, imag} */,
  {32'hbffa67f3, 32'hbdc68f36} /* (3, 7, 12) {real, imag} */,
  {32'hbf2244a5, 32'hbf29c9c1} /* (3, 7, 11) {real, imag} */,
  {32'h409280fc, 32'h3f02879f} /* (3, 7, 10) {real, imag} */,
  {32'hbf15def7, 32'h40140267} /* (3, 7, 9) {real, imag} */,
  {32'hc0bc2cfb, 32'h3e646c6e} /* (3, 7, 8) {real, imag} */,
  {32'h40d7700a, 32'h40292b14} /* (3, 7, 7) {real, imag} */,
  {32'hc095e7fe, 32'hc02efae2} /* (3, 7, 6) {real, imag} */,
  {32'hbff339d1, 32'h3ffddd0a} /* (3, 7, 5) {real, imag} */,
  {32'h405a2646, 32'hc02244e6} /* (3, 7, 4) {real, imag} */,
  {32'h40395c9b, 32'hc0e47c83} /* (3, 7, 3) {real, imag} */,
  {32'h3e832974, 32'h3fbb4492} /* (3, 7, 2) {real, imag} */,
  {32'hc0a13a6b, 32'hc03440de} /* (3, 7, 1) {real, imag} */,
  {32'h3d2f77b8, 32'h3ec03d59} /* (3, 7, 0) {real, imag} */,
  {32'hc106e226, 32'hc0bad9eb} /* (3, 6, 15) {real, imag} */,
  {32'h3ed074c2, 32'hbfa81e5d} /* (3, 6, 14) {real, imag} */,
  {32'hbed95429, 32'hbf88606e} /* (3, 6, 13) {real, imag} */,
  {32'hbf1bda83, 32'hc03ece04} /* (3, 6, 12) {real, imag} */,
  {32'h40c2cadb, 32'hc0d30ae8} /* (3, 6, 11) {real, imag} */,
  {32'h3f397839, 32'h406dda49} /* (3, 6, 10) {real, imag} */,
  {32'hc009f839, 32'h406b4d32} /* (3, 6, 9) {real, imag} */,
  {32'hc012398a, 32'hc09c753f} /* (3, 6, 8) {real, imag} */,
  {32'h40cd4e91, 32'h4018f79a} /* (3, 6, 7) {real, imag} */,
  {32'h3f378b44, 32'hbf99c232} /* (3, 6, 6) {real, imag} */,
  {32'h40a6abc0, 32'hbea68ae0} /* (3, 6, 5) {real, imag} */,
  {32'hc0c25638, 32'h41186162} /* (3, 6, 4) {real, imag} */,
  {32'h3f594405, 32'hbdf56372} /* (3, 6, 3) {real, imag} */,
  {32'h401a0df5, 32'hc0297e31} /* (3, 6, 2) {real, imag} */,
  {32'h3fe620fe, 32'h40ba14f1} /* (3, 6, 1) {real, imag} */,
  {32'hc102a751, 32'hbeef19d4} /* (3, 6, 0) {real, imag} */,
  {32'h40ed12f0, 32'hc0d5f56b} /* (3, 5, 15) {real, imag} */,
  {32'h3f95ae03, 32'h3fc9fcc5} /* (3, 5, 14) {real, imag} */,
  {32'hc0cf045e, 32'hc16e4f75} /* (3, 5, 13) {real, imag} */,
  {32'hbef0b576, 32'h3ffb9a33} /* (3, 5, 12) {real, imag} */,
  {32'hbdfba962, 32'h4121dc85} /* (3, 5, 11) {real, imag} */,
  {32'hc0878cf5, 32'h40c0586b} /* (3, 5, 10) {real, imag} */,
  {32'h40c7355e, 32'h401fb972} /* (3, 5, 9) {real, imag} */,
  {32'h3f2d7f8a, 32'hc0089a23} /* (3, 5, 8) {real, imag} */,
  {32'hc0538a82, 32'h3eb2a171} /* (3, 5, 7) {real, imag} */,
  {32'h401ab879, 32'h4092439e} /* (3, 5, 6) {real, imag} */,
  {32'hc017407c, 32'hc009664c} /* (3, 5, 5) {real, imag} */,
  {32'hc17d29da, 32'h4131803f} /* (3, 5, 4) {real, imag} */,
  {32'hc00137fe, 32'hc0124cb9} /* (3, 5, 3) {real, imag} */,
  {32'hbfd52d96, 32'h403d0219} /* (3, 5, 2) {real, imag} */,
  {32'h3ff0f7f6, 32'h4087000e} /* (3, 5, 1) {real, imag} */,
  {32'hbf83407c, 32'hc146487f} /* (3, 5, 0) {real, imag} */,
  {32'h405c37b6, 32'hbe83de9f} /* (3, 4, 15) {real, imag} */,
  {32'h41172118, 32'h4090676f} /* (3, 4, 14) {real, imag} */,
  {32'hbfe5a5aa, 32'h41152ce6} /* (3, 4, 13) {real, imag} */,
  {32'hbe43cb71, 32'hc17af258} /* (3, 4, 12) {real, imag} */,
  {32'hbe8d501a, 32'h407d6b39} /* (3, 4, 11) {real, imag} */,
  {32'h3fb863f3, 32'hbf8f4fd4} /* (3, 4, 10) {real, imag} */,
  {32'hbf6eb275, 32'hbfab3e2c} /* (3, 4, 9) {real, imag} */,
  {32'h402d0dc5, 32'h3fbbf4df} /* (3, 4, 8) {real, imag} */,
  {32'hbfa56c8f, 32'hc09fd571} /* (3, 4, 7) {real, imag} */,
  {32'h411427b1, 32'h3feb3138} /* (3, 4, 6) {real, imag} */,
  {32'hc0cd594e, 32'hbf643428} /* (3, 4, 5) {real, imag} */,
  {32'hc0e55523, 32'h400d2ef8} /* (3, 4, 4) {real, imag} */,
  {32'hc0082f29, 32'h400f72bf} /* (3, 4, 3) {real, imag} */,
  {32'h3d873785, 32'hc0962575} /* (3, 4, 2) {real, imag} */,
  {32'h4186a8d5, 32'h411937c2} /* (3, 4, 1) {real, imag} */,
  {32'hc10fc4eb, 32'hc0eb8788} /* (3, 4, 0) {real, imag} */,
  {32'h3f44a88f, 32'hbf372a1f} /* (3, 3, 15) {real, imag} */,
  {32'h408e5a08, 32'hc1203f02} /* (3, 3, 14) {real, imag} */,
  {32'h40a5e74a, 32'h3e7db0fb} /* (3, 3, 13) {real, imag} */,
  {32'hbf15a8d7, 32'hc0d0dc40} /* (3, 3, 12) {real, imag} */,
  {32'h407270da, 32'hc106dcfc} /* (3, 3, 11) {real, imag} */,
  {32'hc0b21d97, 32'hc04c0830} /* (3, 3, 10) {real, imag} */,
  {32'hbf1ab9a9, 32'h3facfb63} /* (3, 3, 9) {real, imag} */,
  {32'h408ff864, 32'h3e75af3c} /* (3, 3, 8) {real, imag} */,
  {32'hc0bea61c, 32'hc0b51a63} /* (3, 3, 7) {real, imag} */,
  {32'hbeb28a1b, 32'hc12abf9e} /* (3, 3, 6) {real, imag} */,
  {32'hc14bc7cd, 32'h404d2dbd} /* (3, 3, 5) {real, imag} */,
  {32'h3fc03f17, 32'hc104bbf6} /* (3, 3, 4) {real, imag} */,
  {32'hc09b6d32, 32'hc01b422c} /* (3, 3, 3) {real, imag} */,
  {32'h3de1edf4, 32'h4112a104} /* (3, 3, 2) {real, imag} */,
  {32'hc0e6a322, 32'hc0bbcf5c} /* (3, 3, 1) {real, imag} */,
  {32'h40e2426b, 32'h407ebd59} /* (3, 3, 0) {real, imag} */,
  {32'h41196145, 32'h4195dca1} /* (3, 2, 15) {real, imag} */,
  {32'h416502a6, 32'h4145e652} /* (3, 2, 14) {real, imag} */,
  {32'h4081740b, 32'hc1395947} /* (3, 2, 13) {real, imag} */,
  {32'h40c72054, 32'hbe167928} /* (3, 2, 12) {real, imag} */,
  {32'hc03852b5, 32'h412b6247} /* (3, 2, 11) {real, imag} */,
  {32'h3fd19c46, 32'h400b1517} /* (3, 2, 10) {real, imag} */,
  {32'h3f08bd30, 32'hbef8f386} /* (3, 2, 9) {real, imag} */,
  {32'h3fc0a641, 32'h3fc4c810} /* (3, 2, 8) {real, imag} */,
  {32'h3f2429d1, 32'h3ead63eb} /* (3, 2, 7) {real, imag} */,
  {32'hc023c7e0, 32'h3fa7411a} /* (3, 2, 6) {real, imag} */,
  {32'h40c7b596, 32'hbfaf841a} /* (3, 2, 5) {real, imag} */,
  {32'h40fb43d7, 32'h3ff96528} /* (3, 2, 4) {real, imag} */,
  {32'hc043824e, 32'hc04320b1} /* (3, 2, 3) {real, imag} */,
  {32'h41268ded, 32'hc132ba34} /* (3, 2, 2) {real, imag} */,
  {32'hc0be9944, 32'h3da352c8} /* (3, 2, 1) {real, imag} */,
  {32'hc1321b7a, 32'hc068041f} /* (3, 2, 0) {real, imag} */,
  {32'h40cbfdf3, 32'hc0d4d676} /* (3, 1, 15) {real, imag} */,
  {32'hc176b20b, 32'hc07d95bb} /* (3, 1, 14) {real, imag} */,
  {32'hc0bd0339, 32'hc0e51bd2} /* (3, 1, 13) {real, imag} */,
  {32'h4039dea8, 32'hbce733c4} /* (3, 1, 12) {real, imag} */,
  {32'hc0370230, 32'h3f9bf946} /* (3, 1, 11) {real, imag} */,
  {32'hbfdceed1, 32'h4051424e} /* (3, 1, 10) {real, imag} */,
  {32'hc10ee7db, 32'hbfc2bca1} /* (3, 1, 9) {real, imag} */,
  {32'hbf41b865, 32'h4038e5ba} /* (3, 1, 8) {real, imag} */,
  {32'h3ee0d7d7, 32'hbfc1168f} /* (3, 1, 7) {real, imag} */,
  {32'h409d18b5, 32'hc11fd03f} /* (3, 1, 6) {real, imag} */,
  {32'h3f469aef, 32'h400e0e90} /* (3, 1, 5) {real, imag} */,
  {32'hbfec2936, 32'h3fd0dcd2} /* (3, 1, 4) {real, imag} */,
  {32'h41567895, 32'h411ad06b} /* (3, 1, 3) {real, imag} */,
  {32'h40ce0335, 32'hc08fc691} /* (3, 1, 2) {real, imag} */,
  {32'hc168b51b, 32'h41350bdf} /* (3, 1, 1) {real, imag} */,
  {32'hc10b97b3, 32'h415deff9} /* (3, 1, 0) {real, imag} */,
  {32'hbf9f9ed1, 32'h419d68de} /* (3, 0, 15) {real, imag} */,
  {32'h4188093d, 32'h40dcd2c6} /* (3, 0, 14) {real, imag} */,
  {32'h40be77de, 32'hc029f4ef} /* (3, 0, 13) {real, imag} */,
  {32'hc164d78d, 32'hc132f946} /* (3, 0, 12) {real, imag} */,
  {32'h3faf6c44, 32'h4148daa6} /* (3, 0, 11) {real, imag} */,
  {32'hbedd6488, 32'h3e899dc5} /* (3, 0, 10) {real, imag} */,
  {32'h3fb46335, 32'hbfe8d137} /* (3, 0, 9) {real, imag} */,
  {32'hbfce924b, 32'h40a3e63e} /* (3, 0, 8) {real, imag} */,
  {32'h40f5adba, 32'h3c78ef12} /* (3, 0, 7) {real, imag} */,
  {32'hc0435496, 32'h4045e56f} /* (3, 0, 6) {real, imag} */,
  {32'hbf873a03, 32'hc18b2a03} /* (3, 0, 5) {real, imag} */,
  {32'hc000b965, 32'h40815f00} /* (3, 0, 4) {real, imag} */,
  {32'hc021cf7b, 32'h4109dd2c} /* (3, 0, 3) {real, imag} */,
  {32'h3f64746d, 32'h3fe660f7} /* (3, 0, 2) {real, imag} */,
  {32'h40ef830a, 32'hc1483ce9} /* (3, 0, 1) {real, imag} */,
  {32'h4123be88, 32'hc1a2eb87} /* (3, 0, 0) {real, imag} */,
  {32'h3dd853e8, 32'h419ff426} /* (2, 15, 15) {real, imag} */,
  {32'h41d59e36, 32'hbfb8114f} /* (2, 15, 14) {real, imag} */,
  {32'h409c195e, 32'hc1063807} /* (2, 15, 13) {real, imag} */,
  {32'hc0a43f19, 32'h3f8281cc} /* (2, 15, 12) {real, imag} */,
  {32'hbf3ca61f, 32'h3f2c5a03} /* (2, 15, 11) {real, imag} */,
  {32'hbfbc9772, 32'h3e0be238} /* (2, 15, 10) {real, imag} */,
  {32'hbaae89b8, 32'h40787b64} /* (2, 15, 9) {real, imag} */,
  {32'hbfb0acd3, 32'h3ee18cbc} /* (2, 15, 8) {real, imag} */,
  {32'hc015ac1d, 32'h40b3f5cf} /* (2, 15, 7) {real, imag} */,
  {32'h3ef349d2, 32'hc05816c7} /* (2, 15, 6) {real, imag} */,
  {32'hbf74c4a1, 32'h3fe00257} /* (2, 15, 5) {real, imag} */,
  {32'h3f99241a, 32'h419dc948} /* (2, 15, 4) {real, imag} */,
  {32'hbc852c80, 32'hc0b6397f} /* (2, 15, 3) {real, imag} */,
  {32'hc08dbc97, 32'hc103dc3f} /* (2, 15, 2) {real, imag} */,
  {32'hc14e7e58, 32'h411be58a} /* (2, 15, 1) {real, imag} */,
  {32'hc22204cb, 32'hc08b92c8} /* (2, 15, 0) {real, imag} */,
  {32'hc235186c, 32'h408e37ab} /* (2, 14, 15) {real, imag} */,
  {32'h3fd81f60, 32'h4136b930} /* (2, 14, 14) {real, imag} */,
  {32'h41992c98, 32'h4051db31} /* (2, 14, 13) {real, imag} */,
  {32'hbfe57f63, 32'hc09ce21d} /* (2, 14, 12) {real, imag} */,
  {32'h40914d03, 32'h4049dc03} /* (2, 14, 11) {real, imag} */,
  {32'h3f83cf4d, 32'h4014e5c4} /* (2, 14, 10) {real, imag} */,
  {32'hbf15797c, 32'h401ed5dd} /* (2, 14, 9) {real, imag} */,
  {32'h3d42c9a2, 32'hbec3d88c} /* (2, 14, 8) {real, imag} */,
  {32'hbf99f8bf, 32'hbfbb4d32} /* (2, 14, 7) {real, imag} */,
  {32'h3dc9f830, 32'h3f7b5986} /* (2, 14, 6) {real, imag} */,
  {32'hbff0f5e5, 32'h400585de} /* (2, 14, 5) {real, imag} */,
  {32'hbf942ca6, 32'h411874ce} /* (2, 14, 4) {real, imag} */,
  {32'h3fe8c321, 32'hc1257ee3} /* (2, 14, 3) {real, imag} */,
  {32'h416fe832, 32'hc10e11a0} /* (2, 14, 2) {real, imag} */,
  {32'h418be2e3, 32'hc1d1baeb} /* (2, 14, 1) {real, imag} */,
  {32'hc0d2f493, 32'hc082ff3c} /* (2, 14, 0) {real, imag} */,
  {32'hc09d956e, 32'hbd9db9ac} /* (2, 13, 15) {real, imag} */,
  {32'h3fce6a09, 32'h3fbbdd37} /* (2, 13, 14) {real, imag} */,
  {32'h41411bf8, 32'h40053ae8} /* (2, 13, 13) {real, imag} */,
  {32'h4158f9a1, 32'h4053dfb6} /* (2, 13, 12) {real, imag} */,
  {32'hc09f1e13, 32'hbebed3f1} /* (2, 13, 11) {real, imag} */,
  {32'hc02bb1a3, 32'h40008202} /* (2, 13, 10) {real, imag} */,
  {32'hc0c0ea1b, 32'h3ff3751b} /* (2, 13, 9) {real, imag} */,
  {32'hc00c117e, 32'h3f45db82} /* (2, 13, 8) {real, imag} */,
  {32'h4039f606, 32'h40a44caf} /* (2, 13, 7) {real, imag} */,
  {32'h403fc84a, 32'hc0bf8cc6} /* (2, 13, 6) {real, imag} */,
  {32'h40af1ba5, 32'hc0ab52f6} /* (2, 13, 5) {real, imag} */,
  {32'h3f84c106, 32'h41372222} /* (2, 13, 4) {real, imag} */,
  {32'h3ee7df85, 32'hc09a2027} /* (2, 13, 3) {real, imag} */,
  {32'h3f96623c, 32'h4095dc9e} /* (2, 13, 2) {real, imag} */,
  {32'h40a463b1, 32'h415c557f} /* (2, 13, 1) {real, imag} */,
  {32'hc007c99a, 32'hc002f782} /* (2, 13, 0) {real, imag} */,
  {32'hbf8469e9, 32'h3fc0d386} /* (2, 12, 15) {real, imag} */,
  {32'hc023ce29, 32'hc07a3f90} /* (2, 12, 14) {real, imag} */,
  {32'h3fce97af, 32'h41af75bc} /* (2, 12, 13) {real, imag} */,
  {32'hbf086fdb, 32'hbfb4033d} /* (2, 12, 12) {real, imag} */,
  {32'h4187b5f5, 32'hc0978c8b} /* (2, 12, 11) {real, imag} */,
  {32'hc0520f5c, 32'h3fdc15d9} /* (2, 12, 10) {real, imag} */,
  {32'h3f324b8f, 32'h3fe87114} /* (2, 12, 9) {real, imag} */,
  {32'hc0ad7333, 32'h3fd02556} /* (2, 12, 8) {real, imag} */,
  {32'h40824ca3, 32'hc0a2cdb0} /* (2, 12, 7) {real, imag} */,
  {32'h4065aeaf, 32'hc04734a9} /* (2, 12, 6) {real, imag} */,
  {32'hbf164d62, 32'hc1210048} /* (2, 12, 5) {real, imag} */,
  {32'h410cd4e7, 32'h41742529} /* (2, 12, 4) {real, imag} */,
  {32'h40923a15, 32'hc0d27e62} /* (2, 12, 3) {real, imag} */,
  {32'hbf446ceb, 32'hc04bc527} /* (2, 12, 2) {real, imag} */,
  {32'h4097d034, 32'hc15ddda8} /* (2, 12, 1) {real, imag} */,
  {32'h3ff4fb9c, 32'h4059948d} /* (2, 12, 0) {real, imag} */,
  {32'h41097fba, 32'hc13cc050} /* (2, 11, 15) {real, imag} */,
  {32'h3fd8f2ec, 32'hc0cfafcc} /* (2, 11, 14) {real, imag} */,
  {32'hbf8f2576, 32'h409085f3} /* (2, 11, 13) {real, imag} */,
  {32'hc081dd4d, 32'hc05de783} /* (2, 11, 12) {real, imag} */,
  {32'hc059bf02, 32'h4095db76} /* (2, 11, 11) {real, imag} */,
  {32'h40ce4e3f, 32'h40f7ee37} /* (2, 11, 10) {real, imag} */,
  {32'h4069025e, 32'hc09f1a35} /* (2, 11, 9) {real, imag} */,
  {32'h3e82620a, 32'hc0147c60} /* (2, 11, 8) {real, imag} */,
  {32'h40bc9882, 32'h40eee966} /* (2, 11, 7) {real, imag} */,
  {32'h40e7d599, 32'h3fb47b4a} /* (2, 11, 6) {real, imag} */,
  {32'hc038acfe, 32'h3f8a6a84} /* (2, 11, 5) {real, imag} */,
  {32'h40ae469b, 32'hc042a6e7} /* (2, 11, 4) {real, imag} */,
  {32'hbf7b7280, 32'hc06c52d2} /* (2, 11, 3) {real, imag} */,
  {32'hc0f90562, 32'h4047fa30} /* (2, 11, 2) {real, imag} */,
  {32'hbefc3636, 32'hc0360225} /* (2, 11, 1) {real, imag} */,
  {32'h4063fc9b, 32'h40f3f917} /* (2, 11, 0) {real, imag} */,
  {32'hc01b54d5, 32'h40683223} /* (2, 10, 15) {real, imag} */,
  {32'hc0f7fdd4, 32'hbfabab6b} /* (2, 10, 14) {real, imag} */,
  {32'hc069a39b, 32'hbf178c19} /* (2, 10, 13) {real, imag} */,
  {32'h3fc1d7d2, 32'h40ff572c} /* (2, 10, 12) {real, imag} */,
  {32'hbfa816d0, 32'hbff53f7e} /* (2, 10, 11) {real, imag} */,
  {32'hc08a9599, 32'h3e9e162d} /* (2, 10, 10) {real, imag} */,
  {32'hc03b87d8, 32'hbfc0a318} /* (2, 10, 9) {real, imag} */,
  {32'hc01f7e74, 32'hc0183c3a} /* (2, 10, 8) {real, imag} */,
  {32'hbfaeeb97, 32'hc07b192e} /* (2, 10, 7) {real, imag} */,
  {32'h40868d5a, 32'h3f5959ba} /* (2, 10, 6) {real, imag} */,
  {32'h408b9dda, 32'h403e00be} /* (2, 10, 5) {real, imag} */,
  {32'hc0adcf76, 32'hc0ac93f9} /* (2, 10, 4) {real, imag} */,
  {32'h40cb5ad6, 32'h400b27a9} /* (2, 10, 3) {real, imag} */,
  {32'hc01897f7, 32'hbeb7610b} /* (2, 10, 2) {real, imag} */,
  {32'h4098ea72, 32'h3ec30641} /* (2, 10, 1) {real, imag} */,
  {32'h4084b32d, 32'h3ffc07d8} /* (2, 10, 0) {real, imag} */,
  {32'hc0192c87, 32'hbea5b609} /* (2, 9, 15) {real, imag} */,
  {32'hbd243917, 32'hc015f72b} /* (2, 9, 14) {real, imag} */,
  {32'h3f308496, 32'hc0941ead} /* (2, 9, 13) {real, imag} */,
  {32'h40533f1b, 32'hc090d775} /* (2, 9, 12) {real, imag} */,
  {32'h3f24acec, 32'hc0d7227c} /* (2, 9, 11) {real, imag} */,
  {32'hc0c4d6e1, 32'hc04242d0} /* (2, 9, 10) {real, imag} */,
  {32'h3e6d8c8b, 32'hbea54dfe} /* (2, 9, 9) {real, imag} */,
  {32'h40987881, 32'hc039a288} /* (2, 9, 8) {real, imag} */,
  {32'hbfc52e81, 32'hbf465da7} /* (2, 9, 7) {real, imag} */,
  {32'hc0b036fc, 32'h3f5f7700} /* (2, 9, 6) {real, imag} */,
  {32'hc0fc0bb5, 32'hbe01af94} /* (2, 9, 5) {real, imag} */,
  {32'hc0d50817, 32'h3f9875f3} /* (2, 9, 4) {real, imag} */,
  {32'h40ea6a50, 32'h3fe42b44} /* (2, 9, 3) {real, imag} */,
  {32'hbf72932a, 32'h406ca6a1} /* (2, 9, 2) {real, imag} */,
  {32'hc03b6914, 32'hbe82e22c} /* (2, 9, 1) {real, imag} */,
  {32'h40140570, 32'hbff8d9c3} /* (2, 9, 0) {real, imag} */,
  {32'hc03fc1fc, 32'hbf4b5b57} /* (2, 8, 15) {real, imag} */,
  {32'hc0bc83c4, 32'h40b34c7c} /* (2, 8, 14) {real, imag} */,
  {32'hc093aea1, 32'hbfc49fdc} /* (2, 8, 13) {real, imag} */,
  {32'hc073dd27, 32'h407b31a8} /* (2, 8, 12) {real, imag} */,
  {32'hc086cd8e, 32'h3f94e677} /* (2, 8, 11) {real, imag} */,
  {32'h3f636953, 32'hbf2ed44f} /* (2, 8, 10) {real, imag} */,
  {32'h40264bd0, 32'h40258f28} /* (2, 8, 9) {real, imag} */,
  {32'hbf48663f, 32'hc011baf3} /* (2, 8, 8) {real, imag} */,
  {32'h3e1b04c2, 32'h3fd6f9bd} /* (2, 8, 7) {real, imag} */,
  {32'h4045ebc0, 32'h3fab078e} /* (2, 8, 6) {real, imag} */,
  {32'h40b7a983, 32'h4037c623} /* (2, 8, 5) {real, imag} */,
  {32'hc059c57a, 32'h40ed0f35} /* (2, 8, 4) {real, imag} */,
  {32'hc08e87f2, 32'hc053c7cd} /* (2, 8, 3) {real, imag} */,
  {32'h3fd40658, 32'hbfc011cc} /* (2, 8, 2) {real, imag} */,
  {32'h409d51d2, 32'h3f035c99} /* (2, 8, 1) {real, imag} */,
  {32'h3e293d05, 32'h40821a1a} /* (2, 8, 0) {real, imag} */,
  {32'hc0157bcf, 32'hc014e742} /* (2, 7, 15) {real, imag} */,
  {32'hbfd0b663, 32'hc031c66b} /* (2, 7, 14) {real, imag} */,
  {32'h4024ae04, 32'h40458f0c} /* (2, 7, 13) {real, imag} */,
  {32'hc0915673, 32'h3fa139af} /* (2, 7, 12) {real, imag} */,
  {32'h409d43bd, 32'h3fd8ccb6} /* (2, 7, 11) {real, imag} */,
  {32'h40aeecbb, 32'hc0dc9d30} /* (2, 7, 10) {real, imag} */,
  {32'h402aaf2c, 32'hc081d30e} /* (2, 7, 9) {real, imag} */,
  {32'hbf366e86, 32'h3e2988d8} /* (2, 7, 8) {real, imag} */,
  {32'hbf47d0f7, 32'hc0ab5173} /* (2, 7, 7) {real, imag} */,
  {32'h41557e2c, 32'h401873bb} /* (2, 7, 6) {real, imag} */,
  {32'h40ad562a, 32'hbf8af25b} /* (2, 7, 5) {real, imag} */,
  {32'h3f3891db, 32'h3fb7e398} /* (2, 7, 4) {real, imag} */,
  {32'h3f4828f9, 32'h40b8630f} /* (2, 7, 3) {real, imag} */,
  {32'hc100a3ce, 32'h3e39d365} /* (2, 7, 2) {real, imag} */,
  {32'h40157e41, 32'h3ea30eb5} /* (2, 7, 1) {real, imag} */,
  {32'h4032c568, 32'hbf7007e6} /* (2, 7, 0) {real, imag} */,
  {32'hbff6766e, 32'hc1028c7c} /* (2, 6, 15) {real, imag} */,
  {32'hbe547e19, 32'h3f92a118} /* (2, 6, 14) {real, imag} */,
  {32'hbf8a732a, 32'h3f9ac8a2} /* (2, 6, 13) {real, imag} */,
  {32'h40d0bddb, 32'h3dd20eaa} /* (2, 6, 12) {real, imag} */,
  {32'hc13fcfc6, 32'hbef2e0d6} /* (2, 6, 11) {real, imag} */,
  {32'h40ce4b51, 32'h40b97903} /* (2, 6, 10) {real, imag} */,
  {32'h3fe901f3, 32'h41270ea1} /* (2, 6, 9) {real, imag} */,
  {32'h40736640, 32'hbf8227f5} /* (2, 6, 8) {real, imag} */,
  {32'h3fd2c0c9, 32'hc05a5adb} /* (2, 6, 7) {real, imag} */,
  {32'hc0841881, 32'h41527f70} /* (2, 6, 6) {real, imag} */,
  {32'hc11d37a8, 32'hbf87fb3b} /* (2, 6, 5) {real, imag} */,
  {32'hc0c1f600, 32'hbff8ac2c} /* (2, 6, 4) {real, imag} */,
  {32'h40b9c3ea, 32'hbfa6edb3} /* (2, 6, 3) {real, imag} */,
  {32'h402e219b, 32'hbf15aa2d} /* (2, 6, 2) {real, imag} */,
  {32'h3e456cc9, 32'h40f8d03b} /* (2, 6, 1) {real, imag} */,
  {32'hc003b8ce, 32'h4021c4c6} /* (2, 6, 0) {real, imag} */,
  {32'hc0953ac1, 32'hbf83b58b} /* (2, 5, 15) {real, imag} */,
  {32'h403f209c, 32'h4019f228} /* (2, 5, 14) {real, imag} */,
  {32'h406cb527, 32'h4123fc25} /* (2, 5, 13) {real, imag} */,
  {32'hbfe21dc8, 32'hbfac9415} /* (2, 5, 12) {real, imag} */,
  {32'hbfa38739, 32'hc1139ebc} /* (2, 5, 11) {real, imag} */,
  {32'hc10b0155, 32'h41839231} /* (2, 5, 10) {real, imag} */,
  {32'h3ffbaef3, 32'hc0da8be0} /* (2, 5, 9) {real, imag} */,
  {32'h3f9605c9, 32'h3ef58fc4} /* (2, 5, 8) {real, imag} */,
  {32'hc0245a35, 32'h3fba9350} /* (2, 5, 7) {real, imag} */,
  {32'hc131ffb6, 32'hbf8eac4c} /* (2, 5, 6) {real, imag} */,
  {32'h40454948, 32'hbfa8d4a0} /* (2, 5, 5) {real, imag} */,
  {32'h40bbda2c, 32'hc108872e} /* (2, 5, 4) {real, imag} */,
  {32'hbead2021, 32'h4105bae4} /* (2, 5, 3) {real, imag} */,
  {32'h41096033, 32'h3e986b2b} /* (2, 5, 2) {real, imag} */,
  {32'hc03d0a00, 32'hc0fbae05} /* (2, 5, 1) {real, imag} */,
  {32'hc07dc4e3, 32'h40f3d682} /* (2, 5, 0) {real, imag} */,
  {32'h41192742, 32'h3f958c90} /* (2, 4, 15) {real, imag} */,
  {32'h3ff9ac31, 32'h410f674e} /* (2, 4, 14) {real, imag} */,
  {32'hbf483ae3, 32'hc05f6ec5} /* (2, 4, 13) {real, imag} */,
  {32'hbfc66537, 32'hc0dc84a5} /* (2, 4, 12) {real, imag} */,
  {32'h4023fada, 32'hc070922b} /* (2, 4, 11) {real, imag} */,
  {32'h4077456a, 32'hc0f6e070} /* (2, 4, 10) {real, imag} */,
  {32'h40a61242, 32'hc0849214} /* (2, 4, 9) {real, imag} */,
  {32'h3e06ccf4, 32'h401d96cc} /* (2, 4, 8) {real, imag} */,
  {32'h40db856f, 32'h403f5506} /* (2, 4, 7) {real, imag} */,
  {32'hc0dc2dfd, 32'h3e97332f} /* (2, 4, 6) {real, imag} */,
  {32'h40f4ad67, 32'h4064eae9} /* (2, 4, 5) {real, imag} */,
  {32'h40000b1b, 32'hbfb1696d} /* (2, 4, 4) {real, imag} */,
  {32'hc1367c70, 32'hc10a42d2} /* (2, 4, 3) {real, imag} */,
  {32'hc138f5bc, 32'hbfc59c6a} /* (2, 4, 2) {real, imag} */,
  {32'hc11ad0c1, 32'hc00af0e4} /* (2, 4, 1) {real, imag} */,
  {32'hc1259084, 32'hc0370775} /* (2, 4, 0) {real, imag} */,
  {32'h40b47ad8, 32'hc10538cc} /* (2, 3, 15) {real, imag} */,
  {32'h4145100c, 32'h408b98a0} /* (2, 3, 14) {real, imag} */,
  {32'hbff17a90, 32'hc150cb25} /* (2, 3, 13) {real, imag} */,
  {32'hc0e98d0c, 32'hc073d71c} /* (2, 3, 12) {real, imag} */,
  {32'hc075c5ef, 32'hc07a6488} /* (2, 3, 11) {real, imag} */,
  {32'hc10dee0f, 32'h40c32137} /* (2, 3, 10) {real, imag} */,
  {32'hc0ad0563, 32'hbf716673} /* (2, 3, 9) {real, imag} */,
  {32'hc0245e41, 32'hc013a146} /* (2, 3, 8) {real, imag} */,
  {32'hc060afa7, 32'h3ff20b64} /* (2, 3, 7) {real, imag} */,
  {32'hbfe4c6b1, 32'h40bb16b4} /* (2, 3, 6) {real, imag} */,
  {32'h3ff0fb35, 32'hc0bd7de0} /* (2, 3, 5) {real, imag} */,
  {32'hc10c95d0, 32'hc0d1bb36} /* (2, 3, 4) {real, imag} */,
  {32'hc13519e1, 32'hc0127b39} /* (2, 3, 3) {real, imag} */,
  {32'hbf05e791, 32'hbf821a99} /* (2, 3, 2) {real, imag} */,
  {32'h40ac54ec, 32'hbfa01c65} /* (2, 3, 1) {real, imag} */,
  {32'hc15ebb3a, 32'hbe25193d} /* (2, 3, 0) {real, imag} */,
  {32'h413a6e0e, 32'hc0990c4d} /* (2, 2, 15) {real, imag} */,
  {32'hc1bbaff9, 32'hc1722424} /* (2, 2, 14) {real, imag} */,
  {32'hc14ce3a8, 32'h415ddf6c} /* (2, 2, 13) {real, imag} */,
  {32'h3f0ecb42, 32'h402bf287} /* (2, 2, 12) {real, imag} */,
  {32'h40563996, 32'hc129effb} /* (2, 2, 11) {real, imag} */,
  {32'h4084f3ac, 32'hbddad7dc} /* (2, 2, 10) {real, imag} */,
  {32'hc02c4d2f, 32'h405b002d} /* (2, 2, 9) {real, imag} */,
  {32'hc040a2b6, 32'h3f338b3e} /* (2, 2, 8) {real, imag} */,
  {32'h3efcd575, 32'hc13d4aca} /* (2, 2, 7) {real, imag} */,
  {32'hc110827b, 32'h40c0f788} /* (2, 2, 6) {real, imag} */,
  {32'hc08cc4ba, 32'h402e9de6} /* (2, 2, 5) {real, imag} */,
  {32'h41844830, 32'h4149dc2a} /* (2, 2, 4) {real, imag} */,
  {32'h4125e688, 32'h408e49bf} /* (2, 2, 3) {real, imag} */,
  {32'hc0fde47a, 32'h4105ddd6} /* (2, 2, 2) {real, imag} */,
  {32'hbff67419, 32'h415149a8} /* (2, 2, 1) {real, imag} */,
  {32'h40a9e51d, 32'hc08f1ccb} /* (2, 2, 0) {real, imag} */,
  {32'hc03698a7, 32'hc07e8863} /* (2, 1, 15) {real, imag} */,
  {32'h411508b0, 32'h406d83c3} /* (2, 1, 14) {real, imag} */,
  {32'h413badbe, 32'hc1a49a44} /* (2, 1, 13) {real, imag} */,
  {32'hc158b11b, 32'h404ee17f} /* (2, 1, 12) {real, imag} */,
  {32'h404ac1c8, 32'hbf93e8ae} /* (2, 1, 11) {real, imag} */,
  {32'hc100b4f7, 32'h3fc537ea} /* (2, 1, 10) {real, imag} */,
  {32'h4037dd78, 32'h409f430d} /* (2, 1, 9) {real, imag} */,
  {32'h3e2c0d4a, 32'hbe5d82e4} /* (2, 1, 8) {real, imag} */,
  {32'h40b84a73, 32'h3fbc64ab} /* (2, 1, 7) {real, imag} */,
  {32'hc01aae7a, 32'hbe50bfef} /* (2, 1, 6) {real, imag} */,
  {32'hc13b2cb5, 32'h40327736} /* (2, 1, 5) {real, imag} */,
  {32'h402cf484, 32'hc0c0a7c8} /* (2, 1, 4) {real, imag} */,
  {32'hbfaac18a, 32'hc14c955f} /* (2, 1, 3) {real, imag} */,
  {32'h3d23688c, 32'h419e2294} /* (2, 1, 2) {real, imag} */,
  {32'hc23327f3, 32'h419ade10} /* (2, 1, 1) {real, imag} */,
  {32'h41aae521, 32'h407ed176} /* (2, 1, 0) {real, imag} */,
  {32'h4096977f, 32'hc0ed4fe7} /* (2, 0, 15) {real, imag} */,
  {32'hc1165c31, 32'h403c94c7} /* (2, 0, 14) {real, imag} */,
  {32'h41641223, 32'hc072da92} /* (2, 0, 13) {real, imag} */,
  {32'hc0af23fd, 32'hbfba7dfa} /* (2, 0, 12) {real, imag} */,
  {32'h40d044b4, 32'hc01c8ebf} /* (2, 0, 11) {real, imag} */,
  {32'hbfcc3abe, 32'h4101a282} /* (2, 0, 10) {real, imag} */,
  {32'hbf6dd62f, 32'hc0816368} /* (2, 0, 9) {real, imag} */,
  {32'h40c816bf, 32'h40285e06} /* (2, 0, 8) {real, imag} */,
  {32'h3d43bced, 32'hbf32687b} /* (2, 0, 7) {real, imag} */,
  {32'hbfdbc11b, 32'hbf1685b0} /* (2, 0, 6) {real, imag} */,
  {32'hc14951d7, 32'hbf72251f} /* (2, 0, 5) {real, imag} */,
  {32'hbf2b74a2, 32'hc15ca590} /* (2, 0, 4) {real, imag} */,
  {32'hc1241861, 32'hc097f0ae} /* (2, 0, 3) {real, imag} */,
  {32'hbe9ffd8a, 32'h3d348ce6} /* (2, 0, 2) {real, imag} */,
  {32'h415e4540, 32'h40a94fff} /* (2, 0, 1) {real, imag} */,
  {32'h41e91fb8, 32'hc281efb1} /* (2, 0, 0) {real, imag} */,
  {32'hc0f281fe, 32'hc1056a1c} /* (1, 15, 15) {real, imag} */,
  {32'hc03d76d1, 32'h4196b22e} /* (1, 15, 14) {real, imag} */,
  {32'h4107c53a, 32'hc04e7503} /* (1, 15, 13) {real, imag} */,
  {32'hbe1cf784, 32'h40addc6a} /* (1, 15, 12) {real, imag} */,
  {32'hc12f0083, 32'h410d2ab0} /* (1, 15, 11) {real, imag} */,
  {32'h401c393d, 32'hc038d6f7} /* (1, 15, 10) {real, imag} */,
  {32'hbe254606, 32'hc0f72b59} /* (1, 15, 9) {real, imag} */,
  {32'hc074933f, 32'hbfc49775} /* (1, 15, 8) {real, imag} */,
  {32'h405eb8f1, 32'h3fa3cc8c} /* (1, 15, 7) {real, imag} */,
  {32'hc082fd01, 32'hc0c2b7b4} /* (1, 15, 6) {real, imag} */,
  {32'hc063903a, 32'h40b84dab} /* (1, 15, 5) {real, imag} */,
  {32'hc0801ab5, 32'hc0b95c54} /* (1, 15, 4) {real, imag} */,
  {32'hc0dc6e39, 32'hc0e0b850} /* (1, 15, 3) {real, imag} */,
  {32'h41c14442, 32'h41a2ed52} /* (1, 15, 2) {real, imag} */,
  {32'hc174eee3, 32'h4217a280} /* (1, 15, 1) {real, imag} */,
  {32'hc1c7ee53, 32'h41aabbde} /* (1, 15, 0) {real, imag} */,
  {32'h41dfff9d, 32'h4194c48c} /* (1, 14, 15) {real, imag} */,
  {32'hc18443a9, 32'hc1d189af} /* (1, 14, 14) {real, imag} */,
  {32'hc08a4217, 32'hc0d3f94c} /* (1, 14, 13) {real, imag} */,
  {32'hc10e6733, 32'h40550d16} /* (1, 14, 12) {real, imag} */,
  {32'h3ffb74a9, 32'hc1027f09} /* (1, 14, 11) {real, imag} */,
  {32'h4016eb31, 32'h40e67d5d} /* (1, 14, 10) {real, imag} */,
  {32'h41268b1a, 32'hbfebc4e1} /* (1, 14, 9) {real, imag} */,
  {32'hc02b7db1, 32'h3f7d2119} /* (1, 14, 8) {real, imag} */,
  {32'h4116d5bf, 32'h40eccc2c} /* (1, 14, 7) {real, imag} */,
  {32'hc08ebf62, 32'h401ba486} /* (1, 14, 6) {real, imag} */,
  {32'hc08dc219, 32'h40353925} /* (1, 14, 5) {real, imag} */,
  {32'hc08ae559, 32'hc0d1a150} /* (1, 14, 4) {real, imag} */,
  {32'h413e86a7, 32'h41652d93} /* (1, 14, 3) {real, imag} */,
  {32'hc1b973aa, 32'hbd65dcb1} /* (1, 14, 2) {real, imag} */,
  {32'hc2398330, 32'hc0fadc0c} /* (1, 14, 1) {real, imag} */,
  {32'h4105e123, 32'hc1bba2c6} /* (1, 14, 0) {real, imag} */,
  {32'h4135f285, 32'h4035eecb} /* (1, 13, 15) {real, imag} */,
  {32'hbe693de8, 32'hc10fe12e} /* (1, 13, 14) {real, imag} */,
  {32'hc05f091e, 32'h41752b0b} /* (1, 13, 13) {real, imag} */,
  {32'hc11e07fb, 32'h40233346} /* (1, 13, 12) {real, imag} */,
  {32'h4009a0dc, 32'hc0d8a038} /* (1, 13, 11) {real, imag} */,
  {32'hbf023d0b, 32'h4040f249} /* (1, 13, 10) {real, imag} */,
  {32'hc06ee97c, 32'h413e67d7} /* (1, 13, 9) {real, imag} */,
  {32'hc0187793, 32'hc0c9bf22} /* (1, 13, 8) {real, imag} */,
  {32'h3eb4cd7c, 32'h40c516ee} /* (1, 13, 7) {real, imag} */,
  {32'h401b734c, 32'hbee665d5} /* (1, 13, 6) {real, imag} */,
  {32'hc08ffeba, 32'h401353e8} /* (1, 13, 5) {real, imag} */,
  {32'h408c5cd5, 32'h404992f4} /* (1, 13, 4) {real, imag} */,
  {32'hc085eba1, 32'hc1894841} /* (1, 13, 3) {real, imag} */,
  {32'hc0cfa381, 32'h41689415} /* (1, 13, 2) {real, imag} */,
  {32'h415ce201, 32'h40195597} /* (1, 13, 1) {real, imag} */,
  {32'hc1206f34, 32'h41821d47} /* (1, 13, 0) {real, imag} */,
  {32'h3e3e22be, 32'h41bc2cb8} /* (1, 12, 15) {real, imag} */,
  {32'hc17fe5b6, 32'h410ebc4e} /* (1, 12, 14) {real, imag} */,
  {32'hc0513a4f, 32'h413e8a88} /* (1, 12, 13) {real, imag} */,
  {32'h40aa60a0, 32'h401406d6} /* (1, 12, 12) {real, imag} */,
  {32'hbed09a51, 32'hc10d8a4f} /* (1, 12, 11) {real, imag} */,
  {32'hbf81e017, 32'hbf0b8d06} /* (1, 12, 10) {real, imag} */,
  {32'hc1138209, 32'hc0268790} /* (1, 12, 9) {real, imag} */,
  {32'h3f919c30, 32'h401fcc31} /* (1, 12, 8) {real, imag} */,
  {32'hc0006ae3, 32'hc10d3b68} /* (1, 12, 7) {real, imag} */,
  {32'h4052b2da, 32'h4011c2eb} /* (1, 12, 6) {real, imag} */,
  {32'hc08a5e39, 32'h407e8457} /* (1, 12, 5) {real, imag} */,
  {32'hc052d8af, 32'hbf2acc81} /* (1, 12, 4) {real, imag} */,
  {32'h3fb2dcd1, 32'hbffa6ae3} /* (1, 12, 3) {real, imag} */,
  {32'h3fdd00fa, 32'h3e86a062} /* (1, 12, 2) {real, imag} */,
  {32'h403fed67, 32'hc0a0cfa2} /* (1, 12, 1) {real, imag} */,
  {32'hbfb3db82, 32'hc145ad77} /* (1, 12, 0) {real, imag} */,
  {32'h40200a48, 32'hc0cc41f6} /* (1, 11, 15) {real, imag} */,
  {32'hc07f7777, 32'h402decec} /* (1, 11, 14) {real, imag} */,
  {32'h409bb0c2, 32'hc02bf1e9} /* (1, 11, 13) {real, imag} */,
  {32'h40141083, 32'hbe8687c0} /* (1, 11, 12) {real, imag} */,
  {32'h4057c435, 32'hc0d1dd6a} /* (1, 11, 11) {real, imag} */,
  {32'hc0a249f5, 32'h40c29dcb} /* (1, 11, 10) {real, imag} */,
  {32'h4094e041, 32'h40aa1eeb} /* (1, 11, 9) {real, imag} */,
  {32'h3fd751d4, 32'h40097d71} /* (1, 11, 8) {real, imag} */,
  {32'h3f5aca9c, 32'hc0c23cea} /* (1, 11, 7) {real, imag} */,
  {32'h4004948e, 32'h4094776e} /* (1, 11, 6) {real, imag} */,
  {32'h40bd7e27, 32'h3fad10bc} /* (1, 11, 5) {real, imag} */,
  {32'hbe676ef6, 32'h40d375e0} /* (1, 11, 4) {real, imag} */,
  {32'h41534b80, 32'h40d0aab3} /* (1, 11, 3) {real, imag} */,
  {32'hbf5d1fd1, 32'h40c9c918} /* (1, 11, 2) {real, imag} */,
  {32'h40ed19c4, 32'hc087b427} /* (1, 11, 1) {real, imag} */,
  {32'hc0a6826a, 32'h3ea823d1} /* (1, 11, 0) {real, imag} */,
  {32'h40da0d27, 32'hc08cd47c} /* (1, 10, 15) {real, imag} */,
  {32'hc0714624, 32'hbf593dc9} /* (1, 10, 14) {real, imag} */,
  {32'hc01f44cb, 32'hc1138482} /* (1, 10, 13) {real, imag} */,
  {32'hc0ea0a2f, 32'hc06b8147} /* (1, 10, 12) {real, imag} */,
  {32'hbf5a5287, 32'h41122c94} /* (1, 10, 11) {real, imag} */,
  {32'h40641174, 32'h40b9c4b4} /* (1, 10, 10) {real, imag} */,
  {32'h3ff4aec4, 32'hc078e20d} /* (1, 10, 9) {real, imag} */,
  {32'h4094ebcc, 32'hbfd94971} /* (1, 10, 8) {real, imag} */,
  {32'hc098b84a, 32'h40b0a5ad} /* (1, 10, 7) {real, imag} */,
  {32'hc10f43df, 32'hc10478a5} /* (1, 10, 6) {real, imag} */,
  {32'hc061bb61, 32'h3f2564c5} /* (1, 10, 5) {real, imag} */,
  {32'h40f64f95, 32'h3f9e82a9} /* (1, 10, 4) {real, imag} */,
  {32'hbea088e6, 32'hbf3392c0} /* (1, 10, 3) {real, imag} */,
  {32'hbf11342a, 32'hc03fcda4} /* (1, 10, 2) {real, imag} */,
  {32'h409e8ea0, 32'hc102bb7e} /* (1, 10, 1) {real, imag} */,
  {32'h4062734c, 32'h3b75e187} /* (1, 10, 0) {real, imag} */,
  {32'h40242b69, 32'h40180647} /* (1, 9, 15) {real, imag} */,
  {32'hc03b033e, 32'hc00fbe16} /* (1, 9, 14) {real, imag} */,
  {32'hbf903a25, 32'h40d81fdc} /* (1, 9, 13) {real, imag} */,
  {32'h3fdb716e, 32'hbf9767a5} /* (1, 9, 12) {real, imag} */,
  {32'h40504dc4, 32'h40a58469} /* (1, 9, 11) {real, imag} */,
  {32'hbfda9d01, 32'hc0344056} /* (1, 9, 10) {real, imag} */,
  {32'h3e82a052, 32'hc0da7b01} /* (1, 9, 9) {real, imag} */,
  {32'h401e7118, 32'h3ffb3e92} /* (1, 9, 8) {real, imag} */,
  {32'hbf3866f2, 32'h3eee0ac6} /* (1, 9, 7) {real, imag} */,
  {32'h409c42d7, 32'hc06ab150} /* (1, 9, 6) {real, imag} */,
  {32'hc0473e50, 32'hc0a281eb} /* (1, 9, 5) {real, imag} */,
  {32'hc00b9d4f, 32'hc123b09d} /* (1, 9, 4) {real, imag} */,
  {32'hbf96780f, 32'h4011f99b} /* (1, 9, 3) {real, imag} */,
  {32'h40823ccd, 32'hc0925735} /* (1, 9, 2) {real, imag} */,
  {32'h405b3ac7, 32'h4086f4ba} /* (1, 9, 1) {real, imag} */,
  {32'h408970fa, 32'hc02b9f8c} /* (1, 9, 0) {real, imag} */,
  {32'h3fcb1a54, 32'hc0236276} /* (1, 8, 15) {real, imag} */,
  {32'hbfba2c1c, 32'h400fb3de} /* (1, 8, 14) {real, imag} */,
  {32'hbf72ae23, 32'hc0bef5c1} /* (1, 8, 13) {real, imag} */,
  {32'hc0457b78, 32'hbfddc49e} /* (1, 8, 12) {real, imag} */,
  {32'h3f641087, 32'h40b06acb} /* (1, 8, 11) {real, imag} */,
  {32'hc010951c, 32'hbe7f02a7} /* (1, 8, 10) {real, imag} */,
  {32'hbea5f3e2, 32'h4060494b} /* (1, 8, 9) {real, imag} */,
  {32'h40162360, 32'hc0573852} /* (1, 8, 8) {real, imag} */,
  {32'h408d5388, 32'hc05b11a5} /* (1, 8, 7) {real, imag} */,
  {32'hc0d59027, 32'hc01ca943} /* (1, 8, 6) {real, imag} */,
  {32'h3f88a884, 32'h401cd6cc} /* (1, 8, 5) {real, imag} */,
  {32'hc08b1518, 32'h4051cd39} /* (1, 8, 4) {real, imag} */,
  {32'h4018435a, 32'hc01304e9} /* (1, 8, 3) {real, imag} */,
  {32'hc02837db, 32'h402207d6} /* (1, 8, 2) {real, imag} */,
  {32'hc03d7005, 32'hbe893fc2} /* (1, 8, 1) {real, imag} */,
  {32'hbffcb177, 32'hbf1d66e1} /* (1, 8, 0) {real, imag} */,
  {32'h3f9b5826, 32'h3ee69659} /* (1, 7, 15) {real, imag} */,
  {32'hbf55c174, 32'hc0018b11} /* (1, 7, 14) {real, imag} */,
  {32'h3fa0142b, 32'h3fbdbf81} /* (1, 7, 13) {real, imag} */,
  {32'h41200e55, 32'h40061b25} /* (1, 7, 12) {real, imag} */,
  {32'h3f991fba, 32'h3e9aca32} /* (1, 7, 11) {real, imag} */,
  {32'h3fe93910, 32'h3faef098} /* (1, 7, 10) {real, imag} */,
  {32'hc10abbc6, 32'h3f83f683} /* (1, 7, 9) {real, imag} */,
  {32'hbe2edcee, 32'h40014a8c} /* (1, 7, 8) {real, imag} */,
  {32'h4020733d, 32'hbfc844eb} /* (1, 7, 7) {real, imag} */,
  {32'hc0fef844, 32'hc0227cf1} /* (1, 7, 6) {real, imag} */,
  {32'hbfe2038d, 32'hbfb4ad1e} /* (1, 7, 5) {real, imag} */,
  {32'hc074784e, 32'hbfaa6967} /* (1, 7, 4) {real, imag} */,
  {32'h3f58b232, 32'h40211ffb} /* (1, 7, 3) {real, imag} */,
  {32'hc00812b6, 32'hbeaf119f} /* (1, 7, 2) {real, imag} */,
  {32'hbf18370b, 32'hc0a24c45} /* (1, 7, 1) {real, imag} */,
  {32'h40517ede, 32'h3f949bee} /* (1, 7, 0) {real, imag} */,
  {32'h3f5d9414, 32'hc009d5a8} /* (1, 6, 15) {real, imag} */,
  {32'hc06fc600, 32'h4053e090} /* (1, 6, 14) {real, imag} */,
  {32'hbf072e2c, 32'hc08fac98} /* (1, 6, 13) {real, imag} */,
  {32'hbfa0d6d4, 32'hc0af63ec} /* (1, 6, 12) {real, imag} */,
  {32'hbf5d2a26, 32'hc09eb4e2} /* (1, 6, 11) {real, imag} */,
  {32'h3f8b9687, 32'h41120e4a} /* (1, 6, 10) {real, imag} */,
  {32'h409028ba, 32'hc0761289} /* (1, 6, 9) {real, imag} */,
  {32'h40294b3e, 32'hc0bd2d8e} /* (1, 6, 8) {real, imag} */,
  {32'hbf5f3723, 32'h409163a8} /* (1, 6, 7) {real, imag} */,
  {32'hbf64d309, 32'h3f9e8efe} /* (1, 6, 6) {real, imag} */,
  {32'h4110fda0, 32'hbdcd2d7f} /* (1, 6, 5) {real, imag} */,
  {32'h41676393, 32'h3fcb1dbe} /* (1, 6, 4) {real, imag} */,
  {32'hc119ce31, 32'hc02ea9d9} /* (1, 6, 3) {real, imag} */,
  {32'hc095906e, 32'hbf296fec} /* (1, 6, 2) {real, imag} */,
  {32'hc0cd2b2e, 32'h4009f0aa} /* (1, 6, 1) {real, imag} */,
  {32'h40bc13d8, 32'h3ef5e5e2} /* (1, 6, 0) {real, imag} */,
  {32'hc0b27248, 32'h3f0fe108} /* (1, 5, 15) {real, imag} */,
  {32'h41278eb7, 32'hc1567416} /* (1, 5, 14) {real, imag} */,
  {32'hbfdce858, 32'h3e95db80} /* (1, 5, 13) {real, imag} */,
  {32'h3e644b44, 32'hbfff9367} /* (1, 5, 12) {real, imag} */,
  {32'h408cf11c, 32'h4110dcbe} /* (1, 5, 11) {real, imag} */,
  {32'hc045b7de, 32'h3eaf6185} /* (1, 5, 10) {real, imag} */,
  {32'hc0bfeef9, 32'h4048d11f} /* (1, 5, 9) {real, imag} */,
  {32'hc03fd695, 32'h406f41e5} /* (1, 5, 8) {real, imag} */,
  {32'h40a9b909, 32'h40b3a25f} /* (1, 5, 7) {real, imag} */,
  {32'h40379a7f, 32'hc07a05e0} /* (1, 5, 6) {real, imag} */,
  {32'hbf458b22, 32'h40d27050} /* (1, 5, 5) {real, imag} */,
  {32'hbf803fa6, 32'h404900a2} /* (1, 5, 4) {real, imag} */,
  {32'hc004c169, 32'hc08aede6} /* (1, 5, 3) {real, imag} */,
  {32'hc0e401fd, 32'h400abb44} /* (1, 5, 2) {real, imag} */,
  {32'h3fe5ab1b, 32'hc018ebe2} /* (1, 5, 1) {real, imag} */,
  {32'hc03703ad, 32'h4167ef7d} /* (1, 5, 0) {real, imag} */,
  {32'h41375898, 32'h40065711} /* (1, 4, 15) {real, imag} */,
  {32'hc0a1aacb, 32'h40603e81} /* (1, 4, 14) {real, imag} */,
  {32'h402844a0, 32'hc0ce9738} /* (1, 4, 13) {real, imag} */,
  {32'hc10690d4, 32'h4185f5b1} /* (1, 4, 12) {real, imag} */,
  {32'hc0e83509, 32'hc01ac7c7} /* (1, 4, 11) {real, imag} */,
  {32'hc081cdfc, 32'hc061ec00} /* (1, 4, 10) {real, imag} */,
  {32'h40b87411, 32'hc0320f21} /* (1, 4, 9) {real, imag} */,
  {32'hbf5491a9, 32'h4076813c} /* (1, 4, 8) {real, imag} */,
  {32'hc080e49a, 32'hbfe1273b} /* (1, 4, 7) {real, imag} */,
  {32'h408af906, 32'h3f909b46} /* (1, 4, 6) {real, imag} */,
  {32'hbfb3a4b4, 32'hc011e30d} /* (1, 4, 5) {real, imag} */,
  {32'hc0c9541d, 32'h402348c2} /* (1, 4, 4) {real, imag} */,
  {32'hc0b5ac32, 32'h3f328b6c} /* (1, 4, 3) {real, imag} */,
  {32'h4037b09f, 32'h3fc730c1} /* (1, 4, 2) {real, imag} */,
  {32'h4114d7f1, 32'hc0c58b5c} /* (1, 4, 1) {real, imag} */,
  {32'hbfbf33fa, 32'hc108ac90} /* (1, 4, 0) {real, imag} */,
  {32'hc15b4b0a, 32'hc1ba5cb3} /* (1, 3, 15) {real, imag} */,
  {32'h40331f45, 32'h41203c61} /* (1, 3, 14) {real, imag} */,
  {32'h40dc9bca, 32'h408c2f64} /* (1, 3, 13) {real, imag} */,
  {32'h411e427b, 32'h40909893} /* (1, 3, 12) {real, imag} */,
  {32'hc0c397f4, 32'h40808795} /* (1, 3, 11) {real, imag} */,
  {32'h3fe4a302, 32'hbf6d9f09} /* (1, 3, 10) {real, imag} */,
  {32'hc044f5f1, 32'h403f0733} /* (1, 3, 9) {real, imag} */,
  {32'hbfd1de4b, 32'h404fa946} /* (1, 3, 8) {real, imag} */,
  {32'hc00c4cae, 32'h40132ba4} /* (1, 3, 7) {real, imag} */,
  {32'hbf172679, 32'hc09e840a} /* (1, 3, 6) {real, imag} */,
  {32'hc0b8be13, 32'hbf003f84} /* (1, 3, 5) {real, imag} */,
  {32'hc129a6d0, 32'hc0d282e5} /* (1, 3, 4) {real, imag} */,
  {32'h40a26de8, 32'hc08ce1fa} /* (1, 3, 3) {real, imag} */,
  {32'h41267575, 32'hc0279acc} /* (1, 3, 2) {real, imag} */,
  {32'hc12586f1, 32'h40e42c79} /* (1, 3, 1) {real, imag} */,
  {32'hc0477230, 32'h40d3282f} /* (1, 3, 0) {real, imag} */,
  {32'hc17f7e0f, 32'h3ff85c38} /* (1, 2, 15) {real, imag} */,
  {32'hc0bd7b2b, 32'h40a6208a} /* (1, 2, 14) {real, imag} */,
  {32'hc063679a, 32'h3f3aa381} /* (1, 2, 13) {real, imag} */,
  {32'h410369cd, 32'h402a8b22} /* (1, 2, 12) {real, imag} */,
  {32'hc05eb9c6, 32'hc045362a} /* (1, 2, 11) {real, imag} */,
  {32'h405cc1cc, 32'h405c16f3} /* (1, 2, 10) {real, imag} */,
  {32'h3fccc00d, 32'hc041d99c} /* (1, 2, 9) {real, imag} */,
  {32'h4073e89b, 32'hbf1884a4} /* (1, 2, 8) {real, imag} */,
  {32'hc0a30357, 32'hc023bb01} /* (1, 2, 7) {real, imag} */,
  {32'hbfc5b821, 32'hbf97e5ea} /* (1, 2, 6) {real, imag} */,
  {32'h40d192f5, 32'hc0888162} /* (1, 2, 5) {real, imag} */,
  {32'hc01ca732, 32'h403cc774} /* (1, 2, 4) {real, imag} */,
  {32'h40b46c87, 32'h3f357254} /* (1, 2, 3) {real, imag} */,
  {32'h41d44b9a, 32'h3e00e7e5} /* (1, 2, 2) {real, imag} */,
  {32'h40b96ba7, 32'h3f974c27} /* (1, 2, 1) {real, imag} */,
  {32'hc0f14c72, 32'hc1b222f3} /* (1, 2, 0) {real, imag} */,
  {32'hc0cf05d6, 32'h420592d9} /* (1, 1, 15) {real, imag} */,
  {32'h41deecc4, 32'hc10c5e8b} /* (1, 1, 14) {real, imag} */,
  {32'hc013c98b, 32'h418b5f4a} /* (1, 1, 13) {real, imag} */,
  {32'h403ab2e6, 32'hc0490cee} /* (1, 1, 12) {real, imag} */,
  {32'h3eb94449, 32'hc0c7560b} /* (1, 1, 11) {real, imag} */,
  {32'h400eb278, 32'hc087b00e} /* (1, 1, 10) {real, imag} */,
  {32'hbf88dc7d, 32'hc0598e5c} /* (1, 1, 9) {real, imag} */,
  {32'hbf261c20, 32'hbf49637c} /* (1, 1, 8) {real, imag} */,
  {32'hc08b8b18, 32'hc09deee8} /* (1, 1, 7) {real, imag} */,
  {32'h405c9995, 32'h3f9c4a4a} /* (1, 1, 6) {real, imag} */,
  {32'hc04118ea, 32'h40ea1cad} /* (1, 1, 5) {real, imag} */,
  {32'h3f510b61, 32'h40ae5903} /* (1, 1, 4) {real, imag} */,
  {32'hc1dc5023, 32'h4047d6e7} /* (1, 1, 3) {real, imag} */,
  {32'hc1df0ca3, 32'hc0cbe9b7} /* (1, 1, 2) {real, imag} */,
  {32'h41bde247, 32'h40321e23} /* (1, 1, 1) {real, imag} */,
  {32'h41707117, 32'hc11c5a46} /* (1, 1, 0) {real, imag} */,
  {32'h420a9b30, 32'hc24fd7ab} /* (1, 0, 15) {real, imag} */,
  {32'hc1072dcd, 32'h420a5b8d} /* (1, 0, 14) {real, imag} */,
  {32'hc0540f9c, 32'hc01a4456} /* (1, 0, 13) {real, imag} */,
  {32'h41b13766, 32'hc10662c3} /* (1, 0, 12) {real, imag} */,
  {32'h404fd7ee, 32'h4081d444} /* (1, 0, 11) {real, imag} */,
  {32'hc060875d, 32'hc185a6dc} /* (1, 0, 10) {real, imag} */,
  {32'hc00264c0, 32'h41077297} /* (1, 0, 9) {real, imag} */,
  {32'h409139b0, 32'hbf8d36c2} /* (1, 0, 8) {real, imag} */,
  {32'hc0f52ed5, 32'hbef2501c} /* (1, 0, 7) {real, imag} */,
  {32'h40f31cb1, 32'hc00f7172} /* (1, 0, 6) {real, imag} */,
  {32'h410e07e8, 32'hc084e3a0} /* (1, 0, 5) {real, imag} */,
  {32'hc063855d, 32'h41009e33} /* (1, 0, 4) {real, imag} */,
  {32'hbe47a2dd, 32'hc1b9de55} /* (1, 0, 3) {real, imag} */,
  {32'h418b1860, 32'hc1d832a9} /* (1, 0, 2) {real, imag} */,
  {32'h4114ee81, 32'h42ce4ee9} /* (1, 0, 1) {real, imag} */,
  {32'hc2395ed2, 32'h42dd263a} /* (1, 0, 0) {real, imag} */,
  {32'h414e7da6, 32'hc2459d0e} /* (0, 15, 15) {real, imag} */,
  {32'hc1c97f9c, 32'hc143a71d} /* (0, 15, 14) {real, imag} */,
  {32'hc08656d3, 32'h40c34713} /* (0, 15, 13) {real, imag} */,
  {32'h4120fa47, 32'h400830d4} /* (0, 15, 12) {real, imag} */,
  {32'h4006794c, 32'h40559b1b} /* (0, 15, 11) {real, imag} */,
  {32'h40a35ba4, 32'h3eec7782} /* (0, 15, 10) {real, imag} */,
  {32'hbe0f6f25, 32'h3ff88f81} /* (0, 15, 9) {real, imag} */,
  {32'h4060b7f3, 32'h4081847d} /* (0, 15, 8) {real, imag} */,
  {32'hc0453a42, 32'h40d5f3da} /* (0, 15, 7) {real, imag} */,
  {32'h40ee9b28, 32'h4060a726} /* (0, 15, 6) {real, imag} */,
  {32'h3f6c0a01, 32'h41344466} /* (0, 15, 5) {real, imag} */,
  {32'h4066f500, 32'hbfdc6c4b} /* (0, 15, 4) {real, imag} */,
  {32'h407b917f, 32'hc1a895b1} /* (0, 15, 3) {real, imag} */,
  {32'hc18a9125, 32'h40f04b6a} /* (0, 15, 2) {real, imag} */,
  {32'hc22c0133, 32'hc1644de9} /* (0, 15, 1) {real, imag} */,
  {32'hc288beac, 32'hc2616ac3} /* (0, 15, 0) {real, imag} */,
  {32'h416058b5, 32'hc0a36f98} /* (0, 14, 15) {real, imag} */,
  {32'hc1825bdf, 32'hc09aab45} /* (0, 14, 14) {real, imag} */,
  {32'h3da5db4e, 32'hc18a4c9b} /* (0, 14, 13) {real, imag} */,
  {32'hc0a77922, 32'hc0255ce2} /* (0, 14, 12) {real, imag} */,
  {32'hc0a1259c, 32'h3fde0f4a} /* (0, 14, 11) {real, imag} */,
  {32'h40155c64, 32'hc0cd8625} /* (0, 14, 10) {real, imag} */,
  {32'h3f41df83, 32'hbee9c514} /* (0, 14, 9) {real, imag} */,
  {32'hbfbe8c4f, 32'hbf02f15e} /* (0, 14, 8) {real, imag} */,
  {32'h3ecefabb, 32'hbf41b514} /* (0, 14, 7) {real, imag} */,
  {32'hc0f1f842, 32'h40f9610b} /* (0, 14, 6) {real, imag} */,
  {32'h40097ef3, 32'hc01aa938} /* (0, 14, 5) {real, imag} */,
  {32'hbf1685e0, 32'h411ada2f} /* (0, 14, 4) {real, imag} */,
  {32'h3f7bb7ed, 32'hc122a316} /* (0, 14, 3) {real, imag} */,
  {32'h417cc82e, 32'hc1884012} /* (0, 14, 2) {real, imag} */,
  {32'hc0c8f354, 32'h41990969} /* (0, 14, 1) {real, imag} */,
  {32'hc047f81d, 32'h41e95d99} /* (0, 14, 0) {real, imag} */,
  {32'h3e8fa9aa, 32'h400fbe9a} /* (0, 13, 15) {real, imag} */,
  {32'hc089cf5b, 32'h3f9a1a8b} /* (0, 13, 14) {real, imag} */,
  {32'h3f063e12, 32'hc151fd8c} /* (0, 13, 13) {real, imag} */,
  {32'hbf84b245, 32'h417fed27} /* (0, 13, 12) {real, imag} */,
  {32'h410e78b2, 32'h408b99b5} /* (0, 13, 11) {real, imag} */,
  {32'hc0b1a7d5, 32'h400c13b3} /* (0, 13, 10) {real, imag} */,
  {32'hbf191ba3, 32'hbffce45e} /* (0, 13, 9) {real, imag} */,
  {32'h4065a34e, 32'h3f06e864} /* (0, 13, 8) {real, imag} */,
  {32'h3ecd09f1, 32'h401d900b} /* (0, 13, 7) {real, imag} */,
  {32'hc11722a5, 32'hbfe2239e} /* (0, 13, 6) {real, imag} */,
  {32'hc06c7f07, 32'h413c5efb} /* (0, 13, 5) {real, imag} */,
  {32'h414658fa, 32'hc0809c53} /* (0, 13, 4) {real, imag} */,
  {32'hc139d44a, 32'h3ffcfb23} /* (0, 13, 3) {real, imag} */,
  {32'hc1199d85, 32'hbeccbcb9} /* (0, 13, 2) {real, imag} */,
  {32'hc1214594, 32'hc1c26a44} /* (0, 13, 1) {real, imag} */,
  {32'h41870b14, 32'hc19d8ad0} /* (0, 13, 0) {real, imag} */,
  {32'h400a9f06, 32'hc0841129} /* (0, 12, 15) {real, imag} */,
  {32'h3fa72601, 32'h40e2988c} /* (0, 12, 14) {real, imag} */,
  {32'hc10104ea, 32'h4008fa91} /* (0, 12, 13) {real, imag} */,
  {32'hc0d1f681, 32'h4160d27b} /* (0, 12, 12) {real, imag} */,
  {32'hc0c0b45d, 32'h40abac8c} /* (0, 12, 11) {real, imag} */,
  {32'hbf73c2ec, 32'hc14e2731} /* (0, 12, 10) {real, imag} */,
  {32'hbfba8fa1, 32'h3f4ac924} /* (0, 12, 9) {real, imag} */,
  {32'h3fdf096f, 32'h408e4f28} /* (0, 12, 8) {real, imag} */,
  {32'hc03ba4b0, 32'hc0bf4dc9} /* (0, 12, 7) {real, imag} */,
  {32'h3fb5d91d, 32'hbff733f9} /* (0, 12, 6) {real, imag} */,
  {32'hbfbc6c4d, 32'h3fcfffe5} /* (0, 12, 5) {real, imag} */,
  {32'hbd99637f, 32'hc11efcbc} /* (0, 12, 4) {real, imag} */,
  {32'hc11e9cf0, 32'h413078a0} /* (0, 12, 3) {real, imag} */,
  {32'hc00b9ef3, 32'hc01b0e50} /* (0, 12, 2) {real, imag} */,
  {32'h419196c8, 32'hc0c72742} /* (0, 12, 1) {real, imag} */,
  {32'h40dc0c6f, 32'h41186820} /* (0, 12, 0) {real, imag} */,
  {32'hc0ad0e61, 32'hc048fe8c} /* (0, 11, 15) {real, imag} */,
  {32'h40939216, 32'h41131673} /* (0, 11, 14) {real, imag} */,
  {32'h40439411, 32'hbfde851c} /* (0, 11, 13) {real, imag} */,
  {32'hbf304506, 32'h3f7ccc5b} /* (0, 11, 12) {real, imag} */,
  {32'h40caf102, 32'hc0b1431e} /* (0, 11, 11) {real, imag} */,
  {32'h400f72cd, 32'h3f819a68} /* (0, 11, 10) {real, imag} */,
  {32'h3fc12ea5, 32'h3fd60560} /* (0, 11, 9) {real, imag} */,
  {32'h40cf1f57, 32'h40dedaf0} /* (0, 11, 8) {real, imag} */,
  {32'hc0219709, 32'hc0892e9f} /* (0, 11, 7) {real, imag} */,
  {32'h4104b0b9, 32'hbffd1d09} /* (0, 11, 6) {real, imag} */,
  {32'hc01cb420, 32'hbe224e43} /* (0, 11, 5) {real, imag} */,
  {32'h4028ddbb, 32'hbeb449be} /* (0, 11, 4) {real, imag} */,
  {32'hc100fd4c, 32'hc11b4672} /* (0, 11, 3) {real, imag} */,
  {32'h3e32d3c4, 32'hc13787d2} /* (0, 11, 2) {real, imag} */,
  {32'h409422ea, 32'h3c305820} /* (0, 11, 1) {real, imag} */,
  {32'h40e843f3, 32'h40cd2708} /* (0, 11, 0) {real, imag} */,
  {32'h40b1826b, 32'h3fddc0b2} /* (0, 10, 15) {real, imag} */,
  {32'h40a3bff6, 32'hc0aaa759} /* (0, 10, 14) {real, imag} */,
  {32'h402401c8, 32'h409b2ad2} /* (0, 10, 13) {real, imag} */,
  {32'hc0ae6d2c, 32'h40bc5da0} /* (0, 10, 12) {real, imag} */,
  {32'hc0a44f13, 32'h3e1a6c2e} /* (0, 10, 11) {real, imag} */,
  {32'h3fe6c76d, 32'h40d08ad0} /* (0, 10, 10) {real, imag} */,
  {32'h3fa0507c, 32'hc02be93f} /* (0, 10, 9) {real, imag} */,
  {32'h3d872bde, 32'hc1123437} /* (0, 10, 8) {real, imag} */,
  {32'h408066e6, 32'h40aee23b} /* (0, 10, 7) {real, imag} */,
  {32'h406a3ddf, 32'h404dafc6} /* (0, 10, 6) {real, imag} */,
  {32'hc09c85e6, 32'hbff8a3c1} /* (0, 10, 5) {real, imag} */,
  {32'h4082b716, 32'h40b195b4} /* (0, 10, 4) {real, imag} */,
  {32'hc01a0291, 32'h409ceb89} /* (0, 10, 3) {real, imag} */,
  {32'h3f97f5b0, 32'h40676453} /* (0, 10, 2) {real, imag} */,
  {32'hc10ee2ac, 32'hc00b5bc4} /* (0, 10, 1) {real, imag} */,
  {32'h40d2a7fb, 32'h3eb55138} /* (0, 10, 0) {real, imag} */,
  {32'h40b54cf5, 32'h40d6ec0d} /* (0, 9, 15) {real, imag} */,
  {32'hc02e4a74, 32'h3fc2429a} /* (0, 9, 14) {real, imag} */,
  {32'hc0abc4be, 32'h3f16fe71} /* (0, 9, 13) {real, imag} */,
  {32'h3ea9e17b, 32'hc0a737c9} /* (0, 9, 12) {real, imag} */,
  {32'h3d96670a, 32'h3f9f5cb7} /* (0, 9, 11) {real, imag} */,
  {32'h405cb694, 32'hbfac243a} /* (0, 9, 10) {real, imag} */,
  {32'h400d2124, 32'h4029dfb4} /* (0, 9, 9) {real, imag} */,
  {32'h3e8df1e5, 32'hbf9204d0} /* (0, 9, 8) {real, imag} */,
  {32'hc00c5604, 32'h3fe8e0c2} /* (0, 9, 7) {real, imag} */,
  {32'h409b0e5c, 32'h40102208} /* (0, 9, 6) {real, imag} */,
  {32'hc0aa02ba, 32'hc047220f} /* (0, 9, 5) {real, imag} */,
  {32'h3fb5b7ab, 32'h404e5f22} /* (0, 9, 4) {real, imag} */,
  {32'hbeac8bb5, 32'hc0c9ee9e} /* (0, 9, 3) {real, imag} */,
  {32'h4026df70, 32'hbf7ffd87} /* (0, 9, 2) {real, imag} */,
  {32'h4096ca87, 32'hbfec464b} /* (0, 9, 1) {real, imag} */,
  {32'h3f8d2e1c, 32'h3f169282} /* (0, 9, 0) {real, imag} */,
  {32'h3f0703d8, 32'hbe9e2191} /* (0, 8, 15) {real, imag} */,
  {32'hbee7337e, 32'hc0c49a0d} /* (0, 8, 14) {real, imag} */,
  {32'h402e8dd3, 32'hc068a689} /* (0, 8, 13) {real, imag} */,
  {32'h4095afc6, 32'hbf0dd740} /* (0, 8, 12) {real, imag} */,
  {32'h3ed754ad, 32'h3f562912} /* (0, 8, 11) {real, imag} */,
  {32'hbfd363da, 32'h3e920a5d} /* (0, 8, 10) {real, imag} */,
  {32'hc015ec21, 32'h3f9ed7a5} /* (0, 8, 9) {real, imag} */,
  {32'hbe9023e6, 32'h00000000} /* (0, 8, 8) {real, imag} */,
  {32'hc015ec21, 32'hbf9ed7a5} /* (0, 8, 7) {real, imag} */,
  {32'hbfd363da, 32'hbe920a5d} /* (0, 8, 6) {real, imag} */,
  {32'h3ed754ad, 32'hbf562912} /* (0, 8, 5) {real, imag} */,
  {32'h4095afc6, 32'h3f0dd740} /* (0, 8, 4) {real, imag} */,
  {32'h402e8dd3, 32'h4068a689} /* (0, 8, 3) {real, imag} */,
  {32'hbee7337e, 32'h40c49a0d} /* (0, 8, 2) {real, imag} */,
  {32'h3f0703d8, 32'h3e9e2191} /* (0, 8, 1) {real, imag} */,
  {32'hc0da7ea8, 32'h00000000} /* (0, 8, 0) {real, imag} */,
  {32'h4096ca87, 32'h3fec464b} /* (0, 7, 15) {real, imag} */,
  {32'h4026df70, 32'h3f7ffd87} /* (0, 7, 14) {real, imag} */,
  {32'hbeac8bb5, 32'h40c9ee9e} /* (0, 7, 13) {real, imag} */,
  {32'h3fb5b7ab, 32'hc04e5f22} /* (0, 7, 12) {real, imag} */,
  {32'hc0aa02ba, 32'h4047220f} /* (0, 7, 11) {real, imag} */,
  {32'h409b0e5c, 32'hc0102208} /* (0, 7, 10) {real, imag} */,
  {32'hc00c5604, 32'hbfe8e0c2} /* (0, 7, 9) {real, imag} */,
  {32'h3e8df1e5, 32'h3f9204d0} /* (0, 7, 8) {real, imag} */,
  {32'h400d2124, 32'hc029dfb4} /* (0, 7, 7) {real, imag} */,
  {32'h405cb694, 32'h3fac243a} /* (0, 7, 6) {real, imag} */,
  {32'h3d96670a, 32'hbf9f5cb7} /* (0, 7, 5) {real, imag} */,
  {32'h3ea9e17b, 32'h40a737c9} /* (0, 7, 4) {real, imag} */,
  {32'hc0abc4be, 32'hbf16fe71} /* (0, 7, 3) {real, imag} */,
  {32'hc02e4a74, 32'hbfc2429a} /* (0, 7, 2) {real, imag} */,
  {32'h40b54cf5, 32'hc0d6ec0d} /* (0, 7, 1) {real, imag} */,
  {32'h3f8d2e1c, 32'hbf169282} /* (0, 7, 0) {real, imag} */,
  {32'hc10ee2ac, 32'h400b5bc4} /* (0, 6, 15) {real, imag} */,
  {32'h3f97f5b0, 32'hc0676453} /* (0, 6, 14) {real, imag} */,
  {32'hc01a0291, 32'hc09ceb89} /* (0, 6, 13) {real, imag} */,
  {32'h4082b716, 32'hc0b195b4} /* (0, 6, 12) {real, imag} */,
  {32'hc09c85e6, 32'h3ff8a3c1} /* (0, 6, 11) {real, imag} */,
  {32'h406a3ddf, 32'hc04dafc6} /* (0, 6, 10) {real, imag} */,
  {32'h408066e6, 32'hc0aee23b} /* (0, 6, 9) {real, imag} */,
  {32'h3d872bde, 32'h41123437} /* (0, 6, 8) {real, imag} */,
  {32'h3fa0507c, 32'h402be93f} /* (0, 6, 7) {real, imag} */,
  {32'h3fe6c76d, 32'hc0d08ad0} /* (0, 6, 6) {real, imag} */,
  {32'hc0a44f13, 32'hbe1a6c2e} /* (0, 6, 5) {real, imag} */,
  {32'hc0ae6d2c, 32'hc0bc5da0} /* (0, 6, 4) {real, imag} */,
  {32'h402401c8, 32'hc09b2ad2} /* (0, 6, 3) {real, imag} */,
  {32'h40a3bff6, 32'h40aaa759} /* (0, 6, 2) {real, imag} */,
  {32'h40b1826b, 32'hbfddc0b2} /* (0, 6, 1) {real, imag} */,
  {32'h40d2a7fb, 32'hbeb55138} /* (0, 6, 0) {real, imag} */,
  {32'h409422ea, 32'hbc305820} /* (0, 5, 15) {real, imag} */,
  {32'h3e32d3c4, 32'h413787d2} /* (0, 5, 14) {real, imag} */,
  {32'hc100fd4c, 32'h411b4672} /* (0, 5, 13) {real, imag} */,
  {32'h4028ddbb, 32'h3eb449be} /* (0, 5, 12) {real, imag} */,
  {32'hc01cb420, 32'h3e224e43} /* (0, 5, 11) {real, imag} */,
  {32'h4104b0b9, 32'h3ffd1d09} /* (0, 5, 10) {real, imag} */,
  {32'hc0219709, 32'h40892e9f} /* (0, 5, 9) {real, imag} */,
  {32'h40cf1f57, 32'hc0dedaf0} /* (0, 5, 8) {real, imag} */,
  {32'h3fc12ea5, 32'hbfd60560} /* (0, 5, 7) {real, imag} */,
  {32'h400f72cd, 32'hbf819a68} /* (0, 5, 6) {real, imag} */,
  {32'h40caf102, 32'h40b1431e} /* (0, 5, 5) {real, imag} */,
  {32'hbf304506, 32'hbf7ccc5b} /* (0, 5, 4) {real, imag} */,
  {32'h40439411, 32'h3fde851c} /* (0, 5, 3) {real, imag} */,
  {32'h40939216, 32'hc1131673} /* (0, 5, 2) {real, imag} */,
  {32'hc0ad0e61, 32'h4048fe8c} /* (0, 5, 1) {real, imag} */,
  {32'h40e843f3, 32'hc0cd2708} /* (0, 5, 0) {real, imag} */,
  {32'h419196c8, 32'h40c72742} /* (0, 4, 15) {real, imag} */,
  {32'hc00b9ef3, 32'h401b0e50} /* (0, 4, 14) {real, imag} */,
  {32'hc11e9cf0, 32'hc13078a0} /* (0, 4, 13) {real, imag} */,
  {32'hbd99637f, 32'h411efcbc} /* (0, 4, 12) {real, imag} */,
  {32'hbfbc6c4d, 32'hbfcfffe5} /* (0, 4, 11) {real, imag} */,
  {32'h3fb5d91d, 32'h3ff733f9} /* (0, 4, 10) {real, imag} */,
  {32'hc03ba4b0, 32'h40bf4dc9} /* (0, 4, 9) {real, imag} */,
  {32'h3fdf096f, 32'hc08e4f28} /* (0, 4, 8) {real, imag} */,
  {32'hbfba8fa1, 32'hbf4ac924} /* (0, 4, 7) {real, imag} */,
  {32'hbf73c2ec, 32'h414e2731} /* (0, 4, 6) {real, imag} */,
  {32'hc0c0b45d, 32'hc0abac8c} /* (0, 4, 5) {real, imag} */,
  {32'hc0d1f681, 32'hc160d27b} /* (0, 4, 4) {real, imag} */,
  {32'hc10104ea, 32'hc008fa91} /* (0, 4, 3) {real, imag} */,
  {32'h3fa72601, 32'hc0e2988c} /* (0, 4, 2) {real, imag} */,
  {32'h400a9f06, 32'h40841129} /* (0, 4, 1) {real, imag} */,
  {32'h40dc0c6f, 32'hc1186820} /* (0, 4, 0) {real, imag} */,
  {32'hc1214594, 32'h41c26a44} /* (0, 3, 15) {real, imag} */,
  {32'hc1199d85, 32'h3eccbcb9} /* (0, 3, 14) {real, imag} */,
  {32'hc139d44a, 32'hbffcfb23} /* (0, 3, 13) {real, imag} */,
  {32'h414658fa, 32'h40809c53} /* (0, 3, 12) {real, imag} */,
  {32'hc06c7f07, 32'hc13c5efb} /* (0, 3, 11) {real, imag} */,
  {32'hc11722a5, 32'h3fe2239e} /* (0, 3, 10) {real, imag} */,
  {32'h3ecd09f1, 32'hc01d900b} /* (0, 3, 9) {real, imag} */,
  {32'h4065a34e, 32'hbf06e864} /* (0, 3, 8) {real, imag} */,
  {32'hbf191ba3, 32'h3ffce45e} /* (0, 3, 7) {real, imag} */,
  {32'hc0b1a7d5, 32'hc00c13b3} /* (0, 3, 6) {real, imag} */,
  {32'h410e78b2, 32'hc08b99b5} /* (0, 3, 5) {real, imag} */,
  {32'hbf84b245, 32'hc17fed27} /* (0, 3, 4) {real, imag} */,
  {32'h3f063e12, 32'h4151fd8c} /* (0, 3, 3) {real, imag} */,
  {32'hc089cf5b, 32'hbf9a1a8b} /* (0, 3, 2) {real, imag} */,
  {32'h3e8fa9aa, 32'hc00fbe9a} /* (0, 3, 1) {real, imag} */,
  {32'h41870b14, 32'h419d8ad0} /* (0, 3, 0) {real, imag} */,
  {32'hc0c8f354, 32'hc1990969} /* (0, 2, 15) {real, imag} */,
  {32'h417cc82e, 32'h41884012} /* (0, 2, 14) {real, imag} */,
  {32'h3f7bb7ed, 32'h4122a316} /* (0, 2, 13) {real, imag} */,
  {32'hbf1685e0, 32'hc11ada2f} /* (0, 2, 12) {real, imag} */,
  {32'h40097ef3, 32'h401aa938} /* (0, 2, 11) {real, imag} */,
  {32'hc0f1f842, 32'hc0f9610b} /* (0, 2, 10) {real, imag} */,
  {32'h3ecefabb, 32'h3f41b514} /* (0, 2, 9) {real, imag} */,
  {32'hbfbe8c4f, 32'h3f02f15e} /* (0, 2, 8) {real, imag} */,
  {32'h3f41df83, 32'h3ee9c514} /* (0, 2, 7) {real, imag} */,
  {32'h40155c64, 32'h40cd8625} /* (0, 2, 6) {real, imag} */,
  {32'hc0a1259c, 32'hbfde0f4a} /* (0, 2, 5) {real, imag} */,
  {32'hc0a77922, 32'h40255ce2} /* (0, 2, 4) {real, imag} */,
  {32'h3da5db4e, 32'h418a4c9b} /* (0, 2, 3) {real, imag} */,
  {32'hc1825bdf, 32'h409aab45} /* (0, 2, 2) {real, imag} */,
  {32'h416058b5, 32'h40a36f98} /* (0, 2, 1) {real, imag} */,
  {32'hc047f81d, 32'hc1e95d99} /* (0, 2, 0) {real, imag} */,
  {32'hc22c0133, 32'h41644de9} /* (0, 1, 15) {real, imag} */,
  {32'hc18a9125, 32'hc0f04b6a} /* (0, 1, 14) {real, imag} */,
  {32'h407b917f, 32'h41a895b1} /* (0, 1, 13) {real, imag} */,
  {32'h4066f500, 32'h3fdc6c4b} /* (0, 1, 12) {real, imag} */,
  {32'h3f6c0a01, 32'hc1344466} /* (0, 1, 11) {real, imag} */,
  {32'h40ee9b28, 32'hc060a726} /* (0, 1, 10) {real, imag} */,
  {32'hc0453a42, 32'hc0d5f3da} /* (0, 1, 9) {real, imag} */,
  {32'h4060b7f3, 32'hc081847d} /* (0, 1, 8) {real, imag} */,
  {32'hbe0f6f25, 32'hbff88f81} /* (0, 1, 7) {real, imag} */,
  {32'h40a35ba4, 32'hbeec7782} /* (0, 1, 6) {real, imag} */,
  {32'h4006794c, 32'hc0559b1b} /* (0, 1, 5) {real, imag} */,
  {32'h4120fa47, 32'hc00830d4} /* (0, 1, 4) {real, imag} */,
  {32'hc08656d3, 32'hc0c34713} /* (0, 1, 3) {real, imag} */,
  {32'hc1c97f9c, 32'h4143a71d} /* (0, 1, 2) {real, imag} */,
  {32'h414e7da6, 32'h42459d0e} /* (0, 1, 1) {real, imag} */,
  {32'hc288beac, 32'h42616ac3} /* (0, 1, 0) {real, imag} */,
  {32'hc1e478c9, 32'hc14d6cdf} /* (0, 0, 15) {real, imag} */,
  {32'h4108dc85, 32'hc20e117a} /* (0, 0, 14) {real, imag} */,
  {32'h41b7c081, 32'h407e1633} /* (0, 0, 13) {real, imag} */,
  {32'h419201fb, 32'hc083ffdd} /* (0, 0, 12) {real, imag} */,
  {32'h411c2bdc, 32'h40824ded} /* (0, 0, 11) {real, imag} */,
  {32'hc03f0de7, 32'h4160eb69} /* (0, 0, 10) {real, imag} */,
  {32'h40d19163, 32'hc014a5af} /* (0, 0, 9) {real, imag} */,
  {32'hc103e6a0, 32'h00000000} /* (0, 0, 8) {real, imag} */,
  {32'h40d19163, 32'h4014a5af} /* (0, 0, 7) {real, imag} */,
  {32'hc03f0de7, 32'hc160eb69} /* (0, 0, 6) {real, imag} */,
  {32'h411c2bdc, 32'hc0824ded} /* (0, 0, 5) {real, imag} */,
  {32'h419201fb, 32'h4083ffdd} /* (0, 0, 4) {real, imag} */,
  {32'h41b7c081, 32'hc07e1633} /* (0, 0, 3) {real, imag} */,
  {32'h4108dc85, 32'h420e117a} /* (0, 0, 2) {real, imag} */,
  {32'hc1e478c9, 32'h414d6cdf} /* (0, 0, 1) {real, imag} */,
  {32'hbe13431d, 32'h00000000} /* (0, 0, 0) {real, imag} */};
