-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
KS5u/riiaqld4ES5Cy0t/0WGFvYVezdVXUqeWxaqyFeIFconIec1v9MX78JYRVzz
LxELv1iW0o7dppKi+7nU6daohikH493BPoq4NMPLpx1gLGDT8zhIqu99+kFAmvHY
KZv6BxnaRwKB4kbGuEf0T17U5WMbSssdfiiybZhTSSQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 4832)
`protect data_block
TvM8f15tPd3TjjDQIvJfpDrYZHbTa1WKvZzLhmtVGDU3Sr+p6vMJeQw6XkqoKG1x
L6nJa/8zfJlWyMYbkf4JcbkntAceCYwlax0wE1s4kDhnCYfORASsznJTMZLKHN21
RtIiAXrd/9qHTmifAiWc571eYfZRDbP17jE70PPOxfWChTVIYeYKJCAVmzoIImqH
13EHmC14t/5ZpXzCHh0c9oPuEb2qA9OLgHzjeNxqLEKWlr05Vymv69iAvL0WVl3m
wHyeeFl4KTcjAYdxJfsNhFZTGqUkQ68xPSvnhWLEzSM9jprLVaNtA3ATVT7d2MKR
u0iY+9DUZ5+ugEwysqiNv1bKXVgxU1LiQv4RPAzfOPSCm+K7xoJyogrNO9Pw9oce
BhKhYKItu1q/dWWhxcZedZJxWJQT7SiKdXDdInH1DlThntkfme+H+3GbW7gCVOld
MOxDBNT8UxD58dX/v3wQnZhm8L4f8EDJtP6F7Lfj+LlZfU/qpr4boJ7E/FkwvpBL
KUEiS1MDLrOBBa6El0nR8G1iRJdIkcn+9QY4n/GBQzlF8VIs/T/0/hJdCklCjAXu
eMizrZU8dUu8hB147M3BUMNQVgzmkCL+kcMd1KTLtflh2mSlgf8LrhYhpKrn3/gI
/jmBp0mNQJ7JvuJyyu9PVrLL2err3MzYflW/GxeI6kBW5j4nUACBAXz5I+gIeb7j
6d+2CQYL8a9MAl+t4EHNYOLCSLhJxW94aA1mZ24gIui6BABC6V5QYD+wK+9JFJjF
2TUdW4DGHy74EL554UvNVjQc/4fmVHdbDxq2nzwOSmWwV0H1Je6fpW3BRCRxHQTg
xiS0+lVqFVsU7cedqMN5Zm8J8Y535YhGCJSWYEsJVXqmMfkqg3UxdW7P18UDrx9K
TKXaTYQgqaX1n0TBMK1PzbjAvKBJxxc4KE2xHvXS42npEfCbtUvbc2s1i/O/idXX
0qvKyi4KoFVjwwClCaaolTo62sMsCUEAKP2OyqO9DB28ES6M53RmYHb53Nhn524v
Kx/L6Mkx3A9ZDgNkmhUPI2+Wf11rzJcKA/V8WmmaZNMzX085MsyJjycPCH1H3i3s
pI+///MX7l2ifZZ9XJHMojikBvE4iQv7kh3bUDdU1jclwSedkbb8ft3hjg2ncICC
GL3Q1K2Tw5Pi9DSvcdJc2H7Ocg48FAFbikg2XNcvKBPwQdVPbiNWl528e7YKZnd/
1hUpgO7l6w8FZLZdzdukaERKEklJkIrIizF55Cy1EVZSfKfMu4Plnhea8bMkn9vB
VlmijCz4YwqyaT0Nc97XCupUVfrVWEaj7g+lD+fZXQ1OmThp6uTLjHAja6jiIBR9
ljDV+JzjcYX3Elgt96IqfIz/7ULpvQ+vekF/eD8P4CLyLr3phjozIq31qiQqv/7C
qw9CydHvjzyRr/j+E+0v4uexd0eKaFR35dRTMzqM+qUzXcwTsI8T55Fk/zGbGRrI
7KP5ttGE2aVoqovLNJqlh6M5CtgAqJaatBZqoXI+UyBvSgCW59tqTLM0CvLNQpGe
3pbiWofqVf/R3erDfK6+VusVMEsrslUzPaQC8Dhi/I1juh8/pNNF8T31/xnEPhu1
1hXgBH7YuyENbugIMjC5pyZbI0nMwGZF5kMKrlgxeG9CEOLxgE6yOQVV+5FOWwGQ
MByF7kqS7lsJeNibE2Jy6uWOn3qFDvaoidPpcRr68sIYIMPsweiOIiNvvu5S8ZUv
4DNBwuRFULTVow2+Zm0H6Ad54IuDxuU1fst3MQQ07VaFyTP4ZTqCiYJBVYCeIreP
j9K7aeNBMFDdzqU8OKxLPWak4CBILZ67mcs0itxc7qvEEN4DKnir9/POiysRAiaY
/FFDe8ZfyoKl168EnJQE3eD6qPmMuLfyzOWNUMQFxSQrwEGE/oyZ2M4RoifzDOYd
nPGYfQQaQ7uhJCOokeYo8Xlx9CZojItnu3USqcKxGsusTdxVI3CnI9yQeJH3iN5l
Hnv5BXZIeMwcNxGPuco+iRu2lT8FB9z+dUWCsqwjQxUuvhD+tCMzUtPun7zW8xjT
r2h679gVa8wzPSsh5W2y//LyPVz79n4jEP4SF3DODfxPAPssmMkqP5B2HQDfA1Wn
7HR1MhIgJUPu0s9lS/qZq6x41ZG8o6di1ktEJUqTBIIwYGmb+p9qUwb+IXzRFgMU
yTGgl34KmW2FjnJ84ShJeTz7yInD3Q8lYWuWnSRN1DHAVoBC8LU4/LOHYZxyg9/K
o60UxNeMeMl67GyITcXPn90V+avKJgnzA4oUXwhyDJOEsGcCFZUC5gWPNJmVCYnU
IKQ2UMcL3rmADvLNAy6nJLMUvie0PKMqXDgfBAuSCTnzvsgTTR7wy7peLC75lQNU
TfnYLTgZlsnnWKNvw1prHbhytwtBvx4Ych2jSBE8CUgsCCEdmI8zvAHPdqgOcW/P
r0BLW5J41kGCO8xBfcXgl0kO75n38g3guUTlFk7hk0Idt4ZdxEEsscF8CwJe0BDN
yac3IR+aTU9U3e1f+oGcTe5tCibfJ7gaphMDmrTX1dod9ZvsOVEJOQvYVZGfaDBv
VUzGPST6LnSc5kuEeco0xXhI3O7ls02+5XaXDbit4pfTN9Y+EmuUJJrjllj4xMus
0+68nhlBISBJ8RXVq2/bDt93Fe2vKXWqO28viucr9atauPJcoewSUA2Vt6NhKcOB
ohyEQaSj+xiaI7hgq5UMBx+NxK+gGRAkP16k00kJAhO/11SWag0lk18Ebpncf8vA
19QPSk7oqS+lxTlTly0CJKlsXr1bI6eO5cRoJKjpLCq09MzaSmmUqXold8z/oyCY
f5KrwaXMLuIieaj15XqK41xYa0rsjat4VRMHCHh2fEBbdRW7b1pL4jo2t4OAwwYj
obpImMGw06xJ2Jl6RlfijrZP7c07jlD+lf172rTHRt9RhWNtJqbOypdvtwPyoy6E
lrvgcN31e+x2rEGuFuiO2TPoHy+idTa2wRnnTOM5LMZZO1Lpp54l/NlB51yo6apD
EzlWxqA3AK/nL2NJOUnuVMrviIEA8HELOOH+rIUAz2hgG7AEnDOpZMV6B0YpPKDV
NPf3qY5IpbM4TnNmydU6/qVLZq+ZdjHnClnMNshZlfr8VPrHt7xptGyHZUbqtRhw
jsOMMEi+FbEHtalKcrc46KrC+IRHVDoSlBuNILWSrtlieN/msLmov4XYC6OdulUq
8m5emfIVkIDjACkEsjFXVi1PKZTM4uJMHRhLNrKwmTfNQDzQX86n6FD+orT9qnXz
GpBp4xIG+Lvg5rJhusQlWq5L5l9SNgJYQpXigDeJLgA7bDZz702GpVfrMxsjuRez
xrmlwjkPeyxQIr86jaC/029sRPU/Z0Uq9jHM0RL7+nnKSxuQtPH2wjPFVpwQbCKd
KpmrV4qTTXIYUJ74AK1AN3p9QXSnHiiIbfF64cllWrIzcpGmftiTEXlHsIzOJlls
WmM73+GV+fp3xiH1t91jg10XX7sqh+vfIgxJ2yVAgHiVHsaatSa0E/QUK/gqUSiX
QX3FCpbS1g1OaDVnir8p49ZxSdn517LVJlR+aDDEpcdUoMVxRtg6KjgCfoO2aAyd
0zwy81yQej1EJiHkuQ/ceQxXRuVAXky5oT8uk3DRkZX5TuPLDmPsT3T7Rhrf+3DH
cTQnr697ReW8MLzF0PUSf6iR7KhAVYIkhdolLR/FVoBLY7LmDBmX4PKCOSsvZJwl
hMYkmkB8oiZDLBXAUFl1L3o+pBigTKqY9oHzLFk0FPwZciSPnrGGF+I7FEMNEya3
Zz+hyclb3hFccqFKy30l6Ts1P3fSfdOmVnMDE9lKvhKxQWuKTh4EzIRhbelJ9MVc
H57ORkN/WcJXNG7vbTgt36IT/G2iF9i7YqJv05raW6DLVKpyx8uAEpW+gP/a2K9f
tyH6PcAN8bSZL5ZuuycRw/2Izjr8+yFnWwXQmU/PB0beu2/nsnTkY9DsRY3+9KON
mI68KsL52DMGxQJ/hRWeoFZ7tgK/B3Z64yVYWfmFSmu5qSgNPUyFjqNmdMGRtlw8
c387Rsq+Rw0EIYh1tJcHNjOlBWo0k2Kx3Y7hkdtzveCzfqlWP5m0vi/qYXttSf+T
q8g8Z2FXdutegN41yJWEWMlwZCILhZ2H1KoFmWSARwOnOpLL2q9oxlkIuvwYIQNF
CFsXH6dW0kP78vp2HEYjJ3CheSpugrrL7M0jrdixrVZrXoRHzCAN7XR4Ls6C2J9k
HZ9UmxIyv7xCpJmamLqJD5PeZW/kR5z/3o4xMPbGDAWQ7fb3Gd38k/wRmxWZlKHX
gXz7hLJhYb5pWC2ddMd5hyuKgGi00gSIOb1fXDX+vnWWB0If+1w8tPCq0yGeekTU
xzfUs9UXBeCb+8/VKPAgiPRExxSW7OH3SBAkpDkNp3SBO3lbm56JLZU66jNdFh9E
n+FuXT+YVCJ3BREire75NBGHbmEsKRubO3+PL/rQm3Q6WGj5Th1M78R+PSu/uoid
zEFL8SHLFPdpRRRP0PuwWt7AeDVNide8H8UzSX93YIrZmwy30S3JvN12WBTHEERC
qQ8r8GOCglchiG1G9zVSstpnqttZpF9Uk9KJXLeqRHxfqho5TUAVI7CkGmG5dhac
wu3cwvXT5GMwy5pp3nEPXNfDRiraUwWpXInHWAJPWDM+Hh6+ObekEj7wycCBuULA
9FwcjGKFQBzDFJ39d14ELxNmBtaxH+KsSsvjNgsEskY0ADtoqgCO016CA34iLbSd
lpcqGZlQew0sBgijaO/ZfVbkzChIcdOcRV4nt0CpZOrjpENnVQZ2a/LKweh3EeqD
0PuO5qeCSEsalxdfG5sTLDJ1PqT2cUBIS0oQxw5Ll2zGpRrbPXq726mJtHmCPh62
HT+BgiV4XBCFnpyO/bclqrhTRgeHi2TS3QrBOURznr1G91stAKpGk+cowWH7Pbwg
KmTBnlRMlV9KQdgPeXYaG1WQ2OfkWLfBfkozOimaMO9vyMxdxhM5rb6tmEzAUvGB
bgAIBq8fkJZKYcDecgJPpcNBT84CEoT7mwaD/x5d7WkKHIvyA7JrYzSVMZnScYfO
fJeynT5on79w1/BlICeDtiEo29X2l+roa2AeCGtYgZX8sDgU+hHoElSX3O514T5x
w0KhOQSjJkmxYK0pKk+0xYs+eDVxIvZleDaE9FQ8nyWlIt+Lvtqyi9CMNNU6isU6
6k54tqbQ+xB07HiOstVY+R2NpDpwP7fkFmXqi0WWAHkMsentRNt1Vcchp/RsaS/v
CjctXnxkzsZVWySetEsyoXND8DXgAHbgzc3p3C5nhbPxy1IquvRbLVFeUcbWOwK6
ECz8HuWbCpziHi5mO6wz37uB6U4R95DGRTDley0j0pMBTNtbkQREfULhb29IyGXq
5w1hdyteOESkqrrdSa+jK8dZTjg+BVOxORArJFsMWTfgqDPUdm3JBHlssnN6dh94
Xe3L08ZXRTWPJNfGGos+juGGEkD/MPsuJMjUUTtd/RV4FJApTeZLv9N2baB9bEGj
AQAYDpRcQ8dJAtj+3O9ihX42te1Jht5Se8k0c3PIhiUhuEAZUHp4eJ86SV2SkTRX
Mr8n+sjLcbk9aIcsL0WpAt/6Xz+7HujYmlAxDJ8hlhQ2yrbOKGX0oAx1muD31wS3
IKRJ5MTbFBkqEIb3teSWCEDGFvvevdlndZZNQ/GdDVFZ0XmESg1fX/4ztNMTll+u
bRckDlnHd2cQSymemWdBSrqq71pmxSdFpuhoI8RzAOEkEArOX+HDN9sQWaYzzD5Z
8jDq65iMBBYiTBYohvVcw70L5yLGwMTnRW+XB1E1ebIVtOWxKKCcgZoslnU2OY+O
o4K7PTEWPcUswdzHbpa7YAFey/OHS4DxXL7I8JfWPNRLNvC12wH6FRoln6IV6jlh
/BgubrurC/oLSENzcTpJ4hcGttgOq1I0ycacXSq8J6vH7ejJqUr05su/l8e1Vtu5
49HXk8FLdgzKj/YeLO47v3K1erTqSsWr/AuLOW5rAeDHpB5jxsD6cASe5y34Hqzl
iM0VzOY1upUW1B5shW6Jl7IbrifatE171QyPXH1D6qSMSpfTQCHknnJ0SNjVx7Lm
8DbJR8AlRp4WFFDo7hUYsd9rMfpyAS5c9D4MId+Z8FmoKXUzpy7QXSbyrY5SzTAK
h/gOZoaeH3Qoc+cl+eR9TtOaxYPIT2HLIHrPTw9FQMBvxyYPUpnQADic9O7HsAqu
EsabSSU2ipbgXzjuxWz8wPb0BBItVvCZUqZoYA/AEupDQ6DkRb+1y74BfGEWM/r2
frz02Qh4fLtvSGvy/dyUEm/bqE6+WT8izrfuY5VR6NA98cyPSwlRBrWZDt13u/gv
l10xl+iT9ilC8ptuqn/VS/bY2C1jK3u2ATTgse07bNVM/ZGoVAfNkYyNrFADRNK7
YjPplFRjdOvqTQtJp0OGAgncHUApJewIu1Vanjf+bIk=
`protect end_protected
