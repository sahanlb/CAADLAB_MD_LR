-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
CqM9lhPPNZaKe/vxKIhdqE4SjrnjtQslEC4nzsuKsBU7Y+y4T7BImUM/xMPVZIw2
jSYceu8mRS/n+oVheQl3GBpxdxGOSyV6pfzFw03vwQ24HfslPfa7Nx+g1v4SrWVp
dg4+pHBFLFFyHgHNuFcjMbawQ8Q2V19akrWp/8wFC8s=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7920)

`protect DATA_BLOCK
5hKNtOAdXEnhuHDsunKuJpRYw/+/LrI5SsRntZu7ILdhLxA4Ew6iyCf3gX69QbPr
5l7lEypu7EeG7v/w30qbo/b4/8dQ4sX41s1fTDg+Y6y3K24xVD3uwYR0vyTKyHpP
brE+bMTvu74b0wmUrKneTveyC7SkuBNWqggYb7cDlBxNJZaL8r69yXZFWOmqKT1J
iOPK0xkuGEKjvMR0+OMt7b6zNM2nVBviVdpERWxOFnmt4J314YrkDXaiqc7R81X9
YmWk5FWiSa2d85GLHlozVHs43Jd5gMBG6M5JsU9zCgIQqcytgLWUDJoW+b0pyAD7
/Ij+RjfPKOenZMJlOH9WCLz+1PPkWoCmYc7o2bhoOBqtmnp4mShulQ5SjXTFBbat
MANzwLRXbdoJJYtiJiHNIIsMEhIeg7tKWwtWPdQy/H7FTNdi7GRzYlYLDdb8uVPp
PdbXt4V/86uY42mtw3ZFMOFEcfM2qVrQFIL0ruds8LJN7O2+STl/IMTJr5aXnBUo
d86GQRjZ/Ql/cFJs1R/Ej+X8dthDtv9m1I/nnQ+Mv0zIuyNXf4kTkPQnmhubpxee
IIJ+WgqfvnRN/Km5Szh0voVwDRAgMsxn4Z2zdB7D3nCKV8xdg5R2HLzh+BKG9EoS
d3fac2q4fxEVoW+cxfsJFslK+dM/GwK48qEIrQuY7w/jViShLcLInSfuw8maKHkG
isN3LV7vq1PQE/9AIT+niSdysQVPJh3Pw8J7UZIyyDmcH0se59CpQUfgykazqUjC
QtFfho4emCHLI12PPIS+Xo0UUQcyfs5xoRzNN2kIzYOUBI/ojPYaRew9aJgM6X4J
i9zziggEt4I4/JxX8gixV3vljSUykXdJ9tY6efTg68jtQdKHHgdaZbrhRIaLx6cc
lTIn8yQnaY/Ksk1G689nNOqtC619r7pMpIdImDct+7KenWlg4QhLAd6m+IPfiCiB
1cSt1LqZyLCuR2Tur0b3hsj7EcbhGI3l2vfcaZmhORKBZsTM8A3uo9xFmM6FpWPp
IAZiPmNfDGZk2lp62FFBteQyN3P//IGmbjWZ96xTIQdTkUuSTdbWngXx9WxSOtXb
iTFyU/8prwx7skfoF96O0sSaqLn6Us0kAZSzkqyiDOVVW9OBfvQLRrLiY/VNznLg
CvDnLYit4IHDnaOF+YfFM6yTgZwucxQGendyMESZbpkJaWd6lTElWs7xum9q+7Ft
LhH4VgZiYDeXYu5EIYqVLiR67UwwprkRUNOy8CRbMrt0i67jZ7uR/LNgxi2uzKAs
r53RrjFotCM1ZgqKb61WecN293Zk8ltpmg/mxGyd2puRxrsfeicimTiQpVo9RUzN
UQkuInB/zhXLCGEr85ZTRX2Lhul6KvdludvREEwQXpLqXtpzq25BVwSxJozS+yjY
cB/RPQ/iOyjQpM8qjJhPka7mUqppHYr1f8DG0r+pBlBebus8Ju4dbzOWflANRKqx
YkhdEviqk8STajZykly8qPO76da6bfnuMgz+1POakfWf8wgC1E1IG76PJmlKin8Y
5lMxyknQaKWmm1uS8dz19J8uwYklU2weEJ7ewhYjrn9Vg8GkiilVJ0pQJafYOBek
is+813JcAT6RCXifcRAoiKlHGZPKoTL1t8FLsIbas9VF+6UimS8H2zLgl3i4kUJ1
R3gzI0WsV17UjQd/fqJEhN9gMYjMNnaGvqCBtWsXDLTikbfrOGm0JW5AxZgMWBRj
Zy4a0AYZ6kb7fyOudIFQnTGLXm5TjVooNTq40E2AG/pxZ9fnIN0a6KGH6Ls/LWrH
Jn+3s3iDYTByENUP0QNXfBKrooNn+/l8nhAWyv8lh0HHtQw3Sm0ydhk2EZXqWd7H
W1YtU+PPUNwZWQVwUErDldQDn1cLAMHoorCSDpRMsPTYPwECvL4oFXNbZlpO7LGm
8nMty4QrY5eXfaw+OgmabHLKY22ILfcbBsu999iICG+feQAtX9aSNMuN9ixpmSE/
8F3/ROqUra5lJoIa90h1RHRov3MqEK4jvwOVu89kd9vkbwSxW3ckm/Z0wXjvDo03
1LFhFMlJTH8pdveQ8wSiP6IIcwF5Vg/VezbohAMzX5cehGh0eGiGHtZe23FRjKkN
xVveUKX973ytv72jAvtrsR+jOTn1fEqt6W1PTAKv6VJvvrOTycspsAr5qPZm1Qk6
VOMcRWBFIFfJX6jH2sd2KVwn5TiUtPcb+M9DLbt9Q4P46hwHo2v7VuDkU6colt83
9U+7ZECuWVJjo0+NMS7ayanm7hIcVmXISq+t6mk5HxOEj9Y1019Rfm8IW1Z0H0QR
RjO2eAPzhdXBo1KhaISbTwSlnTV/A8KNnA8vDmaT3al799oO4PTXtvEGnHtAsGLd
H7FKQhjP5FkXP99oZlqOIU+gg133hg1ctzfY4D141d8P1ZtzHZQKKsNOaHHh5axr
nrdfWcNn6XMsEkY46JXKkdSXbiCnOqgHI6TMIxU0sDdRTGb/IKKtRGbVl41dW1Ty
OEnQU0DQTn6Gx/LWZj/GUVR9++Plp+80XBnNSW3wIGeVPqMZjbDD7gKxnvddUapz
Mfhr5r+T54DO7CAS8CYeNeFXo0Qbbx+IOZhWuH7/CI6gloFRFoh7P2G/T48nkQw5
bv8iw6kLZxSQgRzRHTqFDprCVkIBiXKobI5gKzC+ZWvXy8qRthbgEi7bMBU5xIgO
huz+ZE18A9CjWZIKW8dnRinDPUB/3WQVVvqMKLOdcKDxJG4KZHmQsIDYnCPQ8p8P
+WtuhqaULO0M/jywESrc5VLiAG/uxKFtVwYQehEXZxUGDO2VCiVd/udQtraLegqZ
dTzVD/HOaFBUZYgiOVCf1UA5oIUTGtzudfusaDgJBQ/W53wUj+y4qHfqFC9JWvIw
LIrWlOyntoLWjl3RbF3Wy1ONMg7dvQlcYsyhnl6WyUmWHGMTA2W0m7qclBI5N1z4
bvH56wFawbnDf4555b5VNYrS8i0zTGKgLkmwCcNem3PXsi7JPWIGENQh/GO/gxbT
LiiTDn89k/gT/8CBsztSwOmTNQk9MGVHIkT9XnZ+ugyuudD/tC/v3UEe1EGH6rZP
jFPlPynkA9wwHGGEgao9YOZ9Pbkq+uAUrRl0IpUVk1/VLUowPggwpIsPmQwhKpPV
CGvXsdnLFpejnz3y5C27LZY6d9jDZHZJ9P8BCTSWxMPQa8zHOujkhzp7W8K1X1vE
yinwCGqLkVO1B/LHeZHqFkcYObJY8zGnanDXyQcLOFTn2aFfr8bi1fRa2S/lZOFz
TsRncWV/LxDpb4f00XD9iE7BdQdASMAvgqQIQVV8AZwJRtwDYHC8HpXoTRSWuwXU
aYUEuJVFYg1zD9zm23PwWJMYII7BxxxL9oHAnM3bb5SoLJIr6YDn6SkI40Plswdf
VPePiGX4pEb56LQAhhV2LIUIXFyd4cRNDI3qWHxiEXmM8G6miyjdr4ItX1wGPGyk
BwY63J/lHbdMXknUjrwwUtK9G3AHxb80f0L+Ui/nSDgIgsecsgYcoPc2KMgCepcW
zdjpNQ6yETvcSREduRpORzn6LYDVfnFAcRJU0Ejdg/JrmOn2YY+AQI3gH2ey9Q4U
Kr0jx8VmCscksP+nXfHI9VkCjfFIzPkYKgNy+vWSSeoddoaky468Wv+jfJ41DSf/
F1eycE9V9HAKbFdZz8wPDGLOe2REkW4xJ9XlsnIwvb+QhOBbpr47B0BXlNhPenms
sFhmQBez3qnus/xRIGbf1gB/oFEQ73JwQZkHlBotfvBZKVSSpVxVYgIgBuAl/XHz
1jVevKyi0voE7jhpCsKFQEV5d/nr7oBalln5BE5c2WR20PrcWkUXVmaUq4wcZo3J
7mgfP58QKYVolgzx5MH6uEPU4Y8TKhtC09Tv2cSt+S85Rv7jgT+yvBvVT0ufLzpj
Vx2+1zPMsBxc1BkWcLTQH8kzNr07Sn9jVtNu5EICiTuVC9NzJ3QunEz1htC7UK0g
pyU9OZurSp2t/2w4OS2sUU2wIEEt7qfrMTcpDFSB4yeBIokiZR1kqLnuy4HiajtF
61c0BbxRAWIbYzjL9gKtFnwUZ2pAys9v5/ht/EzOlHtrmyJft5VIDWLVcCjlRO1G
gT/19uQ3G/pzJPDquCVXAyaPAmaE41ejOxpMnTTmLWYAjT9UdnrC43u0W3x4Lncj
6/ziQPj/mmtgBi+e+9urJ+lV0LagkK1H9pqwfGTioILELgmYoYj4TSvUWTesqrfE
9AvbgW/fw7gOr1JYwxMLUQb2/nkItXEfeIbo8B++eDEcVNDYzzjyqARXRku/SP/a
LnplJ0zPM+itEMBX2XLfHG8kNsGEK0ifHhhscMvyhB/FdQxbtF6yPzFDj3snnQ67
pPH9G22SGqxtWtPI3gPKNTleslKZ2OyfcBo1VsdVDvMQNuFFbDEmPKog7FURQhFj
KzA5KvU1xVQ19wXFQ8ujrA57a1wt/GHNrooXH+YS1rm8EJ+v5FBJJjR9Qk52Mqnl
r5N3999muKIKkyyYq/rUwpFMk+smCeAtYneJY2OqRNVaX67HNSqg4HH/F68H75a8
7p0F2B+LPhAxzQu7s1ybu7J5F0GGJYIzwZ0Vb6SBAiXUVstrV0mTEuGbk7yjZnmY
PuBc4Qqi3wlNi9MB0Tc5N7frowRKWbmSBPqiv2s5XMwKnJ3Nnr+PQmGFb45xTh2G
n7eIVz8Z1lzgh4rTbH/m9D86uyOaNsh/ZqSXaV9V8TSVlx0W0DRkRfhhFa0NTzUZ
owaGaugX8h5u0SHRa3d4xxbiO/mzKM9zQ4AbyM1R+VB8R5aQmAdQdRXSFqpaz+Mo
D65n6PH3MNk5gesTYRttA4ADdjjhZmJyzzV8apQ/6u3t4qnY7VdCpcjlK+3+PBUc
2HgUCON/D1hbHakxRtTfXkK4OFUJT00IzxkOsUKAK1croYkmF15cyc7SMcknM/Bx
sJSg/FztehtPPbCCUGDYeJBBd7nkJ4/IwN9q0LwwmyCnVQdrzdvf702eF3RD2oX7
SfXS4AuSerSqOWJKYvkcxkiR/OBIgWMv9yJE7aClzFyFz0/DSjyEh965zT5HRj0+
fduVzyARmPPdT6FXv9/K1h11mxWLpRZkG+ZmsFA4WfaNARipoEoIqjtVGe9ldeTL
HhXLGgnf/iKRPbTrZAwJvSRtpXy0SDFNmrQbSbZyP5DxHIDsOAdRKqBjJaK6V5Fs
gtp4UHh8GrpfOyhO3p9DiP1O6yP5ja+iXwD3EzFHS4OgVCyv+2FZALi5eX2fPisV
1wQZuzzxA+GdxU5j3b3aQELhDKFI6xQQvUt5/ouLTOX9jKinwoR5sK427Q7rseW7
tmIE0rvHt7x9VkUXknzUOjy5eNjxVL287D9oaMnIx+UnhDbjxnEZhgN+GsJ5veuR
MqA0U0c9knnz0EDkbHgo6WDdjoMFniD6/a5TVh1hqU8Ha7gwSJeIDHpu3yTIsaIr
MsUJxqRz95DlqKhgaR9AhA5b2nBRGTMCOsUC9TbPP+Bp7sMFFWUUZVsK8f4Mg2DL
KUX7h7eqSr6TOfLKaaenFfdWgHn4AxWshWgfJ+VsllaVAEXvuRZsMv+cxndtOaUR
QsJUjE5i7xVhIVHdHmzp19ztGdnu9h9/8/IzBb8uIXTvy47Vsqa3UUm6u1bqDNb1
hTXM8hMRA/H4b5hajyRFZ1yAMV1WLkeyesBLQgg6SzDCy+ftzWpk32hd0RLpGIiF
FQed5IjP2D2BVhm/QTL50xBV+jzpki5McCIQKovA3tpCREweZOiSlrSIvUidsBzY
8ahFFFonPJP2KkZk2v/I8SERv+AvkBVqrwKa2u/7BA3tq+JesViGrj0VvSozuN+6
D8xcOLis6EiH/UoFtqptSY7HGWcjxgMBG6TDOx9etsvdKTfqCUNnEj+Yc2LtcZQU
3SDAC3tRn71L3GCnupJORlPqJ20bm9y+cn4tg8HJTRUiwYwGYpC7mfgoLn6aqWx+
5qLDhReZzucpp43DS/qYsPEUK9cDZ27UUHHoFJVHAwtRAU4/lf7G6V8oXgBmB0nh
cXwenMuXlyZjT6+N9rOwzojI5vbfLe/OoTtfIKfiQ1tzT6d4MUnUx0vmfIlyvhDC
gUFBvbQQ0kYbBxZ+Olwde81B8qiER6FvLsFxFsy3w3pY/tFf6eBRsWgrvVRhvEFx
bz3oLk/4KUtELED5Ou1iOyUXu1XgHxbU+saIAuO9RJkmf2cj8O9tEji5kNgob4tg
bIMem6lhDolb0SZImhsrGEGZL9bjtQe50pQG22j+JxbJfAdKb6Od8ZCL6KafGGVx
iGM4fqKMW/57k4qUyGJxH5EK9JEYCuKnaY6cx/uGaP1kOQYUzKlNekSAM/4vx+eR
nnFE4JSHtwyVpVZpKoArBm84NByHhcK4viyMXf7T5GE7RCJe8OE+VpbENs19LSmx
6kXE1f4aI31nITbQSLymSXiJKiWwoewQa0/B+erSyVRlP2kQ3BZeEt6NUGGQJg5P
Vx8w/P3bEmVmhquueL1qUJWPuiuhvRU74izsmxk6wKkznkYZlJTfS46RDKBNLwO+
pnoKu2cI/3zz5jcvQhGaDrLTBv2LWrFuoYWgRNPmSTi9o2ERRc4jHjmZH2Yrj+6H
JAcMSBphSMxzMFU3ZpjZQlKTGh66X+RkS/baqoEN8QSo18RpWFgOj8xnmpzDY7Iz
F9ppvDLmJigBhGDKKR2PRoGQQZVqOVXS9l8T6Wa73SCKPlxbrky/FU8PWI6bUavP
6M1bvfcHdZzsdx2MWwBows8UgZ7vvX0NEFvfoys+ULtOLlnUgXWcFZk1VjMxA/3T
asc04jdCnGdjVAc9608cbYVmlNhvq3rtTPbNpZgPF9hFy2cjZNcfALj+lPaTY4Jz
saI0lDaRhmqTcySE4LKcywkkMegJlHbb3EJmBAvdm4Tte0yl3Y/RG44zZNKp/cfB
rXxU7Id7TD3jjbIBA0GMWZR2/hzuDxOy7Ektj343AX4UfSa2262BbsyV5+42abFV
B12UbiU60X4/YGGvVHUUS/dTHbGQk4qQ1l71K5RzaL2TculovdfftCsHW6elgx30
q79cN4No9KvIvweGGvjFkhHwqkuPUIsaHPH7/1Oq/p6TZeT5EHwX/YLJyI97MaA3
zqRYLj9HWNEGoOqRJPqF5ErpCwhI2IgHr+3UF0BnFbj2NlYyQgXktEPYfVIjexy6
BGGoKbPZ9Oaz1symxljg+YMuykgASHA/6P4KoyB5QU79l6oZdeywgG0hIuvz3Qc5
kuPp7cSgpcb92rhDkgNlKz7fCK9yKXkraCo5hZNtyLjNJjwYlQo0HmOS3ys99A99
wHix5Cx/V4VXAvdExb1tC2XsrAUkkG2T2mL/anuQMAtghw2fBRiiYyv4S2ZN6//w
LcJEC53kAwjQMqPg0nsUNB0G4uhu/w28KLYaJ3k09PPm6Jw+jmhMpjjBugHbOUR6
xNTElyrt0upZLCdXNpPIa5RJeANqDmsylXYcfh9sGYIbqBtMwjWW+jhYrqX5khTM
XqbBbAz/pcu7KfZ4J70nPDvtvCy1ydryuU84V8biTBAOO0X5xiikKbCIrdJVBEwS
slTsG4i4Ng5Zaj6NLZecT9c+GrzQ+fJYcT8mLYLQc192+D4wUcVMiXITu2AlqmEz
0QuT5CPUHw+NtxkEy88e1Oa4UIMzz6VKKrJgeopZ8UMwuRGZ/W24/kd6LosejB0O
9PDRaowLibk/9XjbyCZMWCWHEuAveLE53YLeoY8CV8EwMyS8NVLtygMHzO3I2UmQ
5BnvVP18Y6y5cut2T+DYdvV3wdsZD+Q+oD5T7tCtOdmv7Te+TKfZ4YMr/piW+dHd
7ZQRt7mIGlTIi7hhMxotO/OLsmtm4Ib5QJCZT25QCIWr/4m9qnKgtlVx/N+AISpa
7lWP4BLJh2n/5u3bmZg416sFXNFc7viaUe2onN7o6GGwXz0W5ZOzQ9/pEoX6sbTR
pehzlT4+cevXh/8wmQywa2/nbt1pnEyWowjSIp58vAvYLxPUnoZ7fy9a7x3Iyspw
wIr+pk5QE8PA1wV6WiAx7zG7oqcICCMJcK4r4Eo8TnKp00ydszSTIVmojtF0zDlM
HjS8uEoGr5n6gSFELXX3zLlFs9yA8WEjsuRHDBbxAZ4lnkMnfUUHoG9SmGvEDyjc
OfcG2OLSKZlUk+bGxf6hprb5EBzjdSmPdrfeLg1mgBmeD1RDR3QE5vDnPxOdOQ0T
CFE/vZpfUPA5KKe/i/LOj8C6sK54KyB0aOerL97tZd7xG7daIlTK8fnUaJ62Z1Wp
zOu/Fj5cfhJOYZfklra2OCjLq3bRJt3JBKGoovn4CcsBZW1e47QfavUw4bMyLOOa
oGwLtEWiXMN8qnrxHrMTCNhCfJ7qIx3Iw40PkTl1SxtMFv2eBY5zKnSZfjs05Hw6
Ks+ew03xbrTIS8DM2G/eWnDZsVUNMhw+XDVw9swZfx4Q2jGNbr4FNlbpZ7XXcoGI
fhPJoH9ZPJLHi6z6zvu4Ch+OkH4HMy6NY4pJClSGhzW56zlTSrx0SNlw983yoDEv
2D2vl4rPadaa0+fFVuEgALlPpw8tVidIxn9Mzjt2dDrx8f+/t3Mvn/uGB809qy30
w8pthi+GMgjNrev4XPLK9ZMtlpWV8W/3Cb43RAySwkdblE58Yf7SMQxhTT2y4R+Q
TCQibI4GkQ45SqBq791nAxxveLYwDES6iC0+SMs29ZAu2XFTCXa5BjMJHamnnbGQ
ERD9lRUh0LkzYWzADdZLYuJfxwD9MULjMDXaEm/UuG9/gsBrXJIrwQvHP7TJ4QG7
TS/qieQLST6y9UxZ6EnwzJkfZiyfZDLzg83LQQHAE0hYVBKSj7GKMgf+zJJG/Lhg
E8yOp54saRdk5MhVbxbM3K6TfX6vXoVS6e9vgC20/NnnAGbaddDiVM30UOK2w6uj
bdIgNgIcrdUB9DVHLmXMjHffBPAZHfzQzwz1vtIuqLQ6ywwdj2N48Nc7j3rGpnfo
EFlUHN6nOGQlQLC5chshMxKov9//QhnBMJi3I4L8osIA6iNLbM/AsiOIiw267WVw
BTXlZiOrOg7b7JGAz1eQow4Ne7OkBDbgSlmcJfiPF+/j+WWk3V77iB/g47Qp5flE
jDqke/gNkbKGfv8VR8vB+yMiyxA6UKla/hSAV98ZHpc8HTD37Ho8vifQAlclN6fN
Fu8CxhN0SU7GhYoK4hJREgFz+ti1olwjMzPyMnuSBiWwZNVIOHZiPBUvI4jFE4zy
5PIi0wEwi0Y6sLrvdYu/jrBT/LuJ5URd1p7ZjwvY1sh+A65LTm1HxyFCdUo7e75a
kfPQJU2ovlfkcqxjonhd0j9EaLhN6PcVgDFXZ4K/yn4LWDLgVs3J/i44MiXy2UYC
Mtea4AzWSuXyj4YUZHxj4/sJ/rU6qgPsGK2ygSiKZiGUaoi9gMG/NdO5n2hhRYuG
htRHZo2Yu/A1aJAhOG3N/z52zSi3bk1f32kuvYZj9W4VDqu+8FHXPuiP3I8tFD71
htP6XhCFQOpYH1V50hOgUpSkh5tyeDkyOj5Q6tqR1NcMwrxSgIpb7Ev4k5bg3hMc
ANur+dlR+RyusZA81XJ3Uqtiu40z0aqJMNxi3igtoDHRNa5uuLque1mO+1vEoCkJ
2piYM1d0M7E/XdXWJ5kWA/LxqRx7n3dw+gBurhqLWqpejWSuJjLBryfw00R5eHX+
h9kqrFvFDR+dPmYZ8eKms5pW66/7JldnqtofEQQSSC/Zg6qISJJTA2HQW6vGaptQ
E3tZYLhM9GIBGH0pnuelCxO/NatAL2l2fQlnKYAQDGoArqGSnRxD9V3FgWmFx/BP
NeddDS1JKBl30MVygXnHucamX/yiDZrSYLhVO4p6SZ/YwBUp786JYg2dNMO49I6+
9eaHyHiku7TnbXfRI+ZhHtv2p91ultjgd5OmLyFNK8d35mixTooxOCkRraukf4F6
JsCvc7k5ypfwfE1NrTnb/3kZg+nkVilPYne8o1qLNapCQxAZPtbn0hviiwwoQXU3
bDShQC4fQA+YgvTJIK7dEwWYGALEDKVk7PdHS7f9DHXHBm7zKwkPLSzWTo7JJvXH
F7Ry+Bj5EenoyfUCjVDw5Vnr2mbkHiyB5Is2U/Nu71T25NIgfpM1UDkESLEKUSaX
FY7iNsK9d8rL8CbV4dp+K5xIoV3Zrh6MP9VqUFrRKdeRc+iDO0X+uNd+pCQwpIlp
RC8F3Y2Thlktjkr7rtW6aGtIG4qdzsH9kzaI3I62zeH4gbIjpxw+zxpd3u1NdwgX
BHkpFOF8wvuq+ZVT5wR+ADLAdPLIShQNf+TsULhIOPyOqGLXmgLVb59+XhX0qRHY
ZPScy5ntQ4wsmDYAA0Dd8OIHOdCutisD2PuMrl6+2/N7c++jFqc6Y5WjYN0rKEoQ
VhNiCxeYMO/XV4QY3NsK6ir1T4rTNUnVDFjAGbcN+Nace20FDxSLNBXt1cuDg1Ky
ZyzN2b5Pqw1cqD1UFPMwYaT1qe+5CfK677ixwB2eA0gWZa8QZdfApf+P1GqK+W6N
3EpCL2t7UWKnOjGP9ZyOunMs0Zaa2SFS5naC+DVQiuKqcPhmd1DL/W0uCXJLj0gO
machO6wwjbWWt2IKk20TEUk0yK0FAUfUQ6FVFXgh4HY=
`protect END_PROTECTED