-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
NKE3RV0yFVr9j4O5QLl+JtW/WTi/4srrQEXyCPNEM/hhpAZ6i4fXLF5w1aKNJl/R
VPNLYkS0hVAkyNrKWmRs/oVGvBVWjDVXZ1ftgcBoWPuMWHC2qgv2LqyRnkT9Hz4u
CnStgYpBIO8P5txHH5S0ZvHIksXwd38yOfmIEFiuNiM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 23287)

`protect DATA_BLOCK
MTTio6YSPGmTDi2TcgRKUcWGPdczmXFVOKEu1N/efpkCpdV+es8tD21pjA8u1hs5
RTxk09DStiI3KAZYM0D4A6gYLSA0WYUMSNkEB440KIdTZwh0Ammc+BffRorndjE8
x5SaOxokhxJC03BBB4N4GbyIG36BhBqhFJAiXjAokAsI9UYilqY7C/aNi2iiDB9m
0ZC7WHYmzWrtC/qXKpbVT0Rr4QQzuZERAJd8Q4edujYEryWkUx74kVHFq1nxD1ju
KUWeoLlblg6zmm5LvQY98Du14VHxewtBTCSMi4jJpwDDzINZCcZ2Rz90q0TX1E7/
4GoAT8yNT3vzv8cGmudkzPMf3er4JUmkAo0MMLbMXGSrXjRjJMIKGiSnRfOwZX2O
pv6Av7KT0RX3S4PVFYKKan7vKmQ+qHhfZobrnkpduzUvuC1lAD46gwc5KLJoi/Ed
pPXpEUFQrEsEFysa6du12PVaiS5MhC5hXXpsG+BUHmseJGf++Hie7K1ZIDKHDsal
uVvTyXrxNINBVoQgxvt5/pcUvNDfKHONBsJAwqHLuZRgrueMZomsklhALnFko8QU
jhBp2u4YqJut3pYGOf+zKfPOtrJIug2mFgfPheCofXN+DvUbLhg9+YzvBpxNN8uC
JgADmx9YX7sV0Apkj2+A0UyYI/RCvICDAfVgp9cc29hH0V278NOe28Rrr+3KPE31
/KpvZQmHHJUCGMalqr8J9+w4IiyJzuEUJyDzpwV2WTSYblpZqywk7WsffjTq6Db2
yxQ+G+TXdXumnLS176I+RG6jEXCvNE6bQe7CibVvtrAEi3moTdOBcFsvD01xlxyC
C8qZEpb0zSZwhwgNJuG7j14v0IvupEQY8Y2Bt5va+30ljsxcDVdX0TAmZCyXq1lL
DtwMbduVQ/iFJc/O9Yv8vYdhbpYOC5L7nZF4ZSUZMCQvZc18JZTF9ILyeXLo+hiA
0Tkbj+1WbP7ne7LGdqYBc35JiHjJHjMaLXQs2r9ORoVV9yEK1lOBPIVWKZl940fA
dDsZDDYpEESGiPgKJY3YBMbjNUfInNBO8ve1lliHQY+I57eL/bKuoko2So2jS9cQ
nn1/QKuaZSoKRi9ktTkEbAs+YFJn9KHv15rRArK2Xx1eJhKbj+8RaK9J4syO7x/z
31L2LN3rZdGMgoF2VexOImITsK2dy78zovZTujw/CYOsqF8i2rjZkarUlywjWF5N
IdV00gK3Mwo9JaxylRps4nQ1zOHEyUlB1QNSRiOgkB1RJPDAphUyvy4sO6R8oc1H
eCt9+ppeyIVMcP2Yn+pfdJ2660CZyBrFDKVzRoLpS1f0WTSsvqs4bBsalocVCvzg
0gURY9IOvltgVTzMEwidiUuqB88H/KEMoVeomGJDbOfuZUNtDZfA4UrGKFRHx4x7
AlWUjHsZida3iAJErgtiGHNFGtsrWCi/X/CACmHyRZADhW2p9yabxqdKc+bHf/2m
eAFRb6awLwPYz2nIiUzTJlefNcq1uhjhnIRjeoLTicjXB1PFn0TtU036M9c+CNMc
G10D8pPiQ/42DE8GiexHCd63ZLnY5Hwce4tnSpTpQhhQuS0/XGEduu3r86DnlezK
y8ldgsG7z2mwEZStR5657+tnUKa6+ml8ELczRwZ9wD8xOXyYpOCRfXAU+h0YNjsx
B67OC2JrKZbFYdI1iEiOC0PyIR445Uxhj7WIwA9gVijz9e5ldJdQi9iXtbc8lwaP
Wk08Y5h5IN1ZV4f8KtBVJwaOP14+puoaFRRbiGFfnZgrtDDXc1exeLfQvgRvPN2j
1En8XCl8zo3Qonha7CN840AwU8qroIj0P5l9/zNYyw6bPgqX5uqpR8XS3594Ze9U
wCx1qDav5cwZGYgPMdGfIx3s0La23CW1QXNcDIlU20MHA5xLv6m2NzhzW3IlKNgu
bUUigocb+pGe6zi0Z7osYWx+xJ011g0xU23Fu2kJ2nmJSqzeHme2H0J/D+Sbc0pk
d8THRat0dsCGa5I1zIARDPcj3I4uEcj3aYR3GCSdDziYHiPHNYFLqLaPGb++hiv9
WGCX7XobQ6Z+lz4LxDeqfAUn7AQSLdQy3uf3dPYq9JDEYbjUTWp3fLmbMyIwKm+R
RH80hJmnLHpszYXBGkMS3AakgQ1PDSYndyf+B+/36lsqZ1vXIdi2Q0ZtGyjF32+j
rzNX/2aFsuP3Ze9oakFgVJeYndyHzysSFbCeutYXOxJm/Ng8l/jPamERI+Ws/0Yc
wkpYf97Lci56DSGJLnNoXdqWqnX5FSZTRBCl+yrGSxr/nj8EzBXMpSk9k7aaXRVh
4ZKo74p7CszDrvaXm9upxxN95FaXMGnPKc5I9sPT5iTJa7FPDZLtLb0RWalun9eW
2GdO25eC5HwaspXgddkCX6zBFpZ+GK18BPijTnVC0K65/uhwBMOQi7+QzlZN5VVH
Yv3DL1WTWqfB+HgcajDVBIVlKpg5rpHvrTkiDNOj810X+D2fH8e3qZLAlPK27D5C
bKbefRfLbPXoqi+7Vctn23fPwYgiSGDpovNMU+SNwbWiADY6DBj5bk5/4e72DabX
qEvlvCeZOeubT4htble1d8/FM4xfsWewun5LUcwHgYN24v/hx1FU9NXerLTe5NN7
0laMfXm8Emvj7hqWpTOPgyeG+MDMFqBCmH2eLIjPtGL+tkvgANfAggn65tnKNJJB
ci21vbx9oNsR/+2ahCkBSpCaBixgn9FEwYOQuqbWhu0dYM2dFvUwBsoYHNkRXSE0
G5+Hwji7ADTumA7Yzr0YtJOPwNJqU4q1KWyUP3VfpYJYPjRuwHnhYHZIUtlIkQDJ
em0nLlsEUazPSoEH+kII6ACX/jRdgHsIOuXmYLKeHTFMJ0PSD4FK4V/R3Go+42RK
Tshh3k7/4vpwNdFjl3Gtu8DbuT5XTnySl0ziBQ4bSUG4aNt8Cyl+Wi8oOWEEKfT7
NA/Nx/kqPMAnWOhWy7/qoBN4mg5zvKqNOyIKknRAM8U449mJAZd9s1vapWsKVgnN
2qdyBYfDvU3rBlH+/BI08hoXbncEQenSDM12REfVhGAIIWfrG6Vsw75vpDA4MRA0
N0oqmNYVS2GQhkQ4Q8Sc5DKbXjdftITVK3k7HFCRXo9avRCxFS3H95qTp9eayXtz
n4JH/glcT3evUlrzURUiynkR0wOUtNVe495nOwXVtmamWxiupw6IvlQ1CEhYbiJd
V2T0idzto7N/lsR+59UwKdQ1Cx7sKS+7QIJ8OB9cQ09mwtIl9jBVRgqdUbBN64+7
vhiSrbTsMqiiiUFYh3ObEWCC6oTvnje8Mqq303tc7xU15j5XmBsmFte60YacjXCC
Xx8e1sJNEJk0gBBNFRBQB7zFZdwf5FcpO7eM5FP6He4OpmwjL8J8Xy3BHQUgOx2p
kWcUbdjTcQAqmSHxBRV530k0hRfwVfKBRasOoQUt52eQ5HOE9oAxhLbAuq1ACPpo
vG8KK3feDRqATamLFzQoUXLgFN5jwZqO4+qjLOdlXLsCjWEPumPWxCqRqdTECOKp
KC7lMYP2dGpWz8ZIANxUziPz3VhkcT3O5Uhets0NkjdHjgPF8tXGAbmNzJ659CWu
YkZ7xmiiXhoUnoecAp6l0b8GloDIXK2jHdF+W5UFu2dZvA4OIdMRtP4R1G9B7i7U
104nWmTJtH8+5qgy1KbVXROuR4+9phjTFp84kgPTNPTgb1Rw92XBn/YWsrUPnj11
K+O+OQLW8T7K1bIrycjhm3fi7DikEXvJPcJhso8bkVL4WNIM1mwxzw8JOBJ3DBC4
Sf/OFJR0jLpK6AN29PWr1kTOF3ctPpKyNsFPEfh4gbiCcn9nd4Q3W0cFlC6ij60/
fuZy2ck9x0M4l/OG36Xuh3BOVblSndZB28AkehBH/qTGYu94TpQpdugR7rrW/WMW
og/zr/jML+6itUArLRJeam4InkiNC3YfPeBx14tKar/dchCKE48PLnOqiU0pA7bu
ZNIBaSKm1dDb7t9S7TZNSv7T5MU98z0ETic/LasZ6ic/rvvGV3lJpnNsV1YGwSj1
9PfhmAdEqSvy9l3uBAjcXuWQS7NwMMtHySM84x8MAtk8R2tpDX6Iolo7LA4r71K8
1inZuToC663cDAKv3p3uekqbmMAvnGP1r9oDimlKSXuvqwF+1ggysVW/nJjBW7c+
mGLZOc1Z0Zjn8CEPn75CQL10hb3qGmnwf8fNIhrKNMyo4I4koLjA/UGiCkJJxnoX
KLGJlY2xmA5+gMqdVUAGLg8E2ajxx3E1nR9J1uU5THWYUAIJWTGxy78rUU8zO2pF
IfRdEO63MNMFYUGhT9hew226t0nzo49uCQvrgy9TpR1FBv9Y85rhoZVaHpGKFCt8
4yvJAUImfBJ0giquzBz+tyMBh1YBd+ItRZzI4zcMS24Hk247fIMylsbrnoosFAZn
A6aKcnQcnwGdGpvD/m6OGYzSu+E7TuOGKgOAfrkyisChT9N24BnZRl/PNgsOXv4v
6j7E4Qtco8P+wBZ8KXVh6b89epy9TP5A9WOCVcNBMyMN7a0h4ywh61ktXJOgSleB
xrNBpvdaO+k/cyilE0fCV3mkF7PxMkXgzj7U08/vm10BWQuQaf0KF+68MvxitEbZ
fhgladkGrodm57tlHDQumjwUHbVx3CoBicNc5vK2zcK35gzLhTDcwhN8gU1Kr7Al
fzd5f8AT1Nt6q3q7TmF4BU5KCfyhCZpoOwsIPp4YjsqPj7GzzXCfN6l4Q+VI8vl7
53ZzxI7qrRoo7SzTHx9v+MGBsY9VbJmjI7I5OIAyrQWqPSCqFn92K22AM0Vo1720
rg+bW2vZq7H/GNRFHf3yZZXSEIQI3d++WNIphSCN8sFsSHFNxPLMGJZDchYKVal6
JYyAeCLOPLelrQC3OgpmrLahylLEva/e2JMrXXi9qWN17nvHb/d3brdGSLd7o4jo
h7Lj2k78UEE2xuUmuOH4u8RyVWzexGWRE6KccSahKVyl/gjJAKhRfcEBgZjFCAn5
8ZQKU/oV4PK8Tbc7cxde1eLZcF4HnthnzztS/YZh3gqttqWslTm/Kz2qe8t8bA5u
LhSOYNuYtn9OUtqzcuMV8wSzdre5tYI+phLZZIGaef5x8VzuMboDWkEA3lqq64ip
/nenOhOthyrBkVdvDdY0i3U9yphhilxuMNXesa0XZdMHH4/D33M+oW/vjIkbxsjW
E7LPjncMR8M/Lc0H0taBDxmkiTaPzpbU8oc++XxRM7tPzeWTFViwRHGrh8Ow7ReH
TjXMl6xvAtaGyqAS5CRc+jAsle6Y66IU0b+MX5iQtDpHjElePIH271Ex6wVkNBX0
3P1vx1fp8Ozy/P5+8zl5iVJ7lS7wVRxBDb0OxteFUQFYmbW+rpw3+SjvcJWhAz7S
JjmVgYAqXnPHqyTeq02PS0XFRdwGbBGY4nImYZiG8yfHSb0JEeWZBdTZebc3B1fd
zRrU2iA0+S3REU4aeX76PB6bWY18+mpIc5IAm+PEnvdcCku4KM4p2liCVb1wYRze
UPmeV9QnECp9YO83GGXOwECcLZnT6TOqjgINb9H4UbfN8HkoKipKevW6ZMweI4wZ
gA/BjK0iPMm5RE99aDBc1yVHboRIQCbW7BKQPCL3/0Hf/YJxZlTJxHLuwKHDCnbJ
iYTwIlcfQbYGUlQmnvr+0o7wdsv3u1bTE+OwHqT9neFFLUL4GCGGnpFk1eFlVPUM
K18Wb10z53pkTjbJDYHoKOFJS1pje3puF61isd4Qa5xHRduwa8mwYmNvQFy2XqXi
RC6JJlKjV7oVyTjdTJii2TWXeST/6Wi19Q3i1hwc9pc9Yml+BFa1FX5H3T6RcMkh
2giqGlobgs/38Nmj9vg89Gh8vMa4YQebz6RnjIuU70EYE/8juhCE1avrYg9yAwNH
VBlcnqMF7qaPLdpwbOGMqjKludk8gYZmHOwAwkWgLTVw187ISIyCe7YNzoWHtS/5
HWqcS9G7ZStdBvGiN1a2cvbQ/WsYYVzs14QQ68XoaIW1haKD6DlDtfpr16fjH9sA
1Hg3J6UdqtkR6siDQjVIMPXlHNWNKU5GUJVZ3uC1WkbmjvIbaSZe8QMB8eYuKm7q
lVkXIih5qycEqQDDAz01OnEjtRDgqfscYrKrlr7NXWT6vg1sC6pMk/hRxgxeeh9I
OviBDLI2FDqVaTln/uFeXh/X0vxUMf46yTjqMd8swuWiOQ+SF54bDiBYX6TVk+al
RWvEqtnsaOkhH6XR92Qm3Sy05Mqt4+DVEEApzsSDsOHiRPoo8dlKL0EUMUWScjNi
6WTEoaxMeqvQBzkiXMeyqbGHfgQgIAVVq+T4SpDTLVckEUD21eHTpuXjtG9wtNjk
BvyGt1AJ37Y0qlyxgThSPOX6/lloMWEBcgl9FvwF7syaA84qqqLMwBEeBlgitEI/
KAzAobBR6h2dO9pmVkivaPU25Crf5nMNcs5oYl8m1iJCZ7pZoT3W7q17XqC59k8u
aGw23YXz/yUS8G/csKxQO1mvgUSCf6Bo8pqaf/yLzjJD1vsoBQLC81zRQ8eC2IQw
IY/Ux4U8oysYzRVzpxcaC1dwWNsKo8iC3fLeVw1BIiWpUGN/wdwYFrfT+bWEjVQ3
XJSUs2h3MUsGnI6Lqr/UiUDyBeL0H++j0jK/ctU9X5Ru3bCPjAgfPkyvbJlvofrE
E1J76WsWNhVtyJ1gkwQMYAbJRJH+Due9nfX+RDTQtgSQ/aWTWBzogV77hHUquG2J
FGRg7urqPE4z4z3d7jiVJYQkuokgI5zEgSKCTDWiPIannaB//klHtPKIGM6Q+WhM
QhVpoFoKXDvU9TKchOnQtZQyAZSGpD9Y74VibCDLUoYEZZTqJ5reolR07uE1S55J
xVyqGMmFdWmxMpWHRvqoqwUY4pYEGgLS5nbPyXZWjV2CpTu0nNyCnrTdrUaTwFtu
aKfv15qzhJAZfSij9wu7/YDe0og86cLMfcy1FQbxgxlpZpsj771hdVb0/X6NXEvu
d/t8jYecvahzKizTGZXHoZAg0+GmwVt5eOP78YizAYFYL4Mrd1EAasjr07gHFmnK
/4LecjlJ1lHj8S8WUcVgX0QP2ApCfCdYiWL/ipbUG1GP8744u1PVAXVmIwKa+Fdp
TiwDY+u6urJ14uievrzh7Nu1BMYoT4nu2x7eWgC9oZ16NtbxzFXLELkBpRraCkeI
dAK6H61Vwus9CltMZEZabvJRUYJn53wu39cNGNftfg/mFN2yjfdYfjRhwaUXwk5m
qJHbd7nZIiuLw+EEZsRsSBLKGKoIQhWr8WX6+568h4CcJQqva3Sk7ep9d5yAUg7z
yvByVpYjxnAJuJUtcdx8enaQhSScaZwVU5kvc2B2k63OPK6FhdW87z3Sw/nfazqk
kOIpKgpjii/HIxS05+BUrzJXfQN31rqItUmKQEo9J4j2Dy5zDZ8MiXGxil80FhJL
aLiA9UMsCHyrX5xq63fM4RWP5a0WruBbk57AwNlv3vaFSF9VaJ1kRZMudyrSt0i+
5U7JALtx5nlLxVxuZ8UDIyVfIsj2+I0SUl1BJJ1hPbZAd/8TU6GLP+lxdg2vHovS
EpvVlyRNvxuCXL3zN/O1anFVNKU4qDcdttdryvlkjXCS/F5o2sh1BRt5trXF+wg/
7RK5ZdY5WHux/8Sx9BkyitWDi64IZC9slPK/IkWgV10fdWxSWEVxYYHWThFiIuRI
QvboVwLZfofUe8UAeSSAIfz85p4o4GyG6VU1NI01+jCuMEU32jkRFWK950fT7YAd
8W1HPhu3ahW2xTlUZe4i2VpFi8Az67v87vtYayRzYTWo77ovyOijc2UFE7dvy2U+
PbRcxfKt5Mq2cAiYn+FOkQ1KNcmurk22D7a/Nra/qnflRBvhtJssKQWZMFPwPaBv
FFqky9Syv3csy4aDL16ay2yfNevmc+jEqmzlBk6Op/RlsDirMcaFmXZF8/NkJjVv
3s7kkwx3b0DT8mUgFUy6oilp+Ac9bvlEDwFyHYKDpxTrT+fizaeeCMe5jK8FURqo
SSiSyzWM9oqrjykC8RjfNpHLJPGXK67AzMk+P8pS2/R8VINKTnZhbLddL4jEwO1U
OzinkpuTYOyrgnTMqWY5UcDUXH5uTHaHVtrsDamGtMA88QtzGUyKf+qa6NxwVlNq
czWB+p1U9v7nEZV8zZtoU/gXLxxkDhxN6w4742HJEMl/+Or4nyoHm/bnjyl88IDY
EUxcPO5FEtCXo99RzOM0HdindjK1GMIFa5gzqGFlzMRbzZOvdqBqextzp4bc3ax/
vfsrFT6jxiWoHTsG2qTJh8wIGxa1ofi34KGIXn4DqTjHSbTlfkT1fsY22WzWK1BL
FW2yo6F3JB1+If11pewOyNsGBa8uNiXA+PMcvM+QMS6rAbt8C7sPyGHcrFUCJ8uv
GjlZmhpmtePfrK9wC/aW2MmY5NPOYZHOPy5Hu6CuKm0++vFZyZnlc1eFjCiqKXhQ
7gWddZAFjzDufVlUhKqpnHkheNG4LDGETCjbna4CRiEXwBTR8FPAxD8BNrXKHjp+
zCUfQ3zmLXx6xiwqBrA2TCADfSaolDlIdiWbBg0MdhcS/mRK08U5L+bvv2yRTEpf
BwFzboNkyBmycEJ1sEySVLpKF+OMf3nqCxayHfY8jzyJOhE9UQMrAw2hmtB6pYPG
eUUg1Bq6l2K+7SdxCSMcOOmPtxrsy3/re02B/SdnqBEhcowawVifbcxSOp/9qcau
OSW2NONK7R23EMUbJPGtmeL33JAnY1LuToWVAt9rAY81hAt3/LsGk6iAMi6NGWOh
2D7fCSR9GbGiw58zauviqAtF2gMASYZIzZdQldks6v1lFkjlyzWfT0IqxVSmLubR
dJhb0CSMHeb7NYnRhyBIfWdY4k7jtlcSW9tCoVBZT4DWE1wD6W7GTTziqSNdjuV/
HGSqq/14BcEBpgjBddyfhTOvKQIa21q2enzN1qwJ2pCC/oYoRYuGS0GdMGW9rchz
GjXA1nzadd5M2p2PvNpEpwbXoFTh/SfRcMoLD5QS8DCwd71ekZQ+Z9dg3w2tZrRi
yVD+mAr70eNbXpuU48JFVmuteo/T4cl4j/s5lJrtIbiMxugnBtItHHqf0tNWXZoW
LJzCEWog9HAJO8BeXuSb7R9ivXOlhmUeS9xKPJ5TmsTGeA6HqgPfo+fjKr4S3hRU
7IjuBqv4QKkO0ZICqm4RsgdZuSFNn4nFWMQhXNVzlikqM9lQS6GFPnlKvOinFq32
JBhEyeI2xaQYh+qLwZmq0yX0e4CWR2B8wZurSBmoyq42XpwTVpz9H8cbV38LZO7c
TjzC2W3WEDWQNxuKuwzDGSgfuvtnA+UCZZqpoCRKHpMZ2gAjbIrXYVAwwv5KhNpg
ywUpw1Rzg9UAEBELBfNu0OhuNARaMAMslu+1MKIWKuhsPcrJ/pyR0mKgCy0BiXWW
zTQ0hZfO9bm0gcG2DCE0aP3G70YIehlJM8dEZa9jMCedIBqX3Jb1U7v7uxSeqMdN
bDFT/WMhLBw4+KbcQ7xA7zm9V22lFlpSkHTWLZPqmrGvuR5vlJQ0ILffkN/g/0HO
dUTH6d23DpNGFpUHgkib1V8wgaeSn2jFAbBQ3eeErr3H4Zkv9C7MWYuYYt1SlrZx
8Zr5NtkeJ9QJ9Ir8noWFY62HzviA2U4tpgGnkBs3nTItfmlzIqTo3hBgBAexpAGi
55T7E+ek0Pm9iXXgHusuVJBhGqMWUyLbDDedqiOIeIfve1/Nx3vvJuFaCMkGRwQB
VHEZrg2guyJ/c6rpNbSMVmR3Aovg5eLCU8Kq5hIYXopYkMT3vhVksJ4JgKk4/o/R
x8ULqxMChsQ2z0wL2I9r90GU3lpt9TqLer6L7NXEO0KJssPRGJ0/nYXqCqugAHAO
lxeBQIth5cIjaRmEhSPQw7qr5BrpFoukY2erdIYwgmA7Fqo+as66pauBz8ArO9pE
iRNo0MmHXzWjTthEbwnD/0IZohjSBl+tGs3vk6F6snmXr81qhY67FB44R7LE6BFx
GXYqbBEcjNSpUFIyRLVoy80+JQupOO58iZZThhjROBoaxAvBcYDGIQxdrclShwpw
0RoKMiyidValfJpKaKlH5lYqioph/rkWZzJUre5dKnhhbJtWTn8/I9DfKoJxyy3k
P4RNNnwa6DQdyV9FrM+HKEPDZq8WHTaqLg9/m/BwfVilx73jZNallHCkeZb6z2+c
CM7oxn23bogKZN2y/G60bbbjABYIc+ZXzQo7W9AgUVocpDL9vWnSuP+MtMhIu4nQ
G5Ss4N63kjAw2Gi8l1bcV8FvC7thcVMXKEOYlsnD2EP+0JglLzm7qNYSMaGAkLlD
ajv29wu/m+IxgighRkg73fJbiqNuBFOnSzybDoNSwOaYKlewFi/ha/IY3mQTLmqe
eGqjZbB/UeX/3dZ/awxv+6eEWG/vZOk5oNs8gwKeJayEubjid2mVTxEoPKrz3fbs
FECNbc2vMoNI2uUwyc683BnLT1aYzv9MDf/3HbwbpYrW5pNa+bNLl2MitXP5yiSW
iWEdi+vrOAoXUATRRZocHjaVNe983Dbbm84cophbI5Q38Hv/ZAw8s+ehsoxW5W0f
aW2i5vXx4bj2TTiSsytVyGoKzE6nR54hmueh6DYvkQjiE4Te/9szg0r3YPiwDksA
loCTQMv8LAFuEScEdgBL3nQq4GJ4KndSXBKRRyeuM4432ehLrxAsU5X39KZAnhdP
JDdIxMAiDt6/Lt/IiTka4GL7Nfth0jOte/Uhz5XnleHboyisRG7V30oCkWep/mWu
TyMzHaL2iVSBdfj2q1yICmXSRktX1oMlYBLKAHDDsa7NVs04VopfW+JUUGrIlPDD
ChS+LMxzwllmphQ3Tj80ZoblRzryGOfTuVD0Ph4qMzs5Yj2DsHssANB5upGf5k0X
bnPW1hN0QXgCLon3wlH1ZA2rAClPuAm8d0F5p/80LQeGr0Upu00lur/+RX9vsXUI
IFdtVE+VqY0zf/Hxfke/PnrBROfj8h7jN+2MHxv/I1ZcRDL4GNAnIPsBU1bWdiL7
7vrL4Xa/imr7LtqWyIC845yutj2CTkYJHBMu8becr2n4hqmhh69IcZ/dJlC7n0Bx
kN+nYtI11PeH9OvI59o/G8MMwNxzB1wyN/ouumXgoDOpqvFTF3Gfr0j7MxKtlV+3
uTRnGzHN8COaYemr2hzYMPbdk0RxO+3V2HbI7sMxLz4xMkQBo2zZkphOCNVrqFph
wB5i0J82G4JLsvKwXqe1LQwez1CleW69QBvFylfh476BR/rS+DPQsNQEMpXPqwnA
8xGd0peIGjafg7Xx8gCKpKoQslBDnNL1xkBlmEkiip9eY9MpPBXfZHqzTUrgeFv3
EUR/+i0TOvLsKqgp1IQSuS9U8iwcqzso7G+VXs4qLDlY1DeuMwJu3162re9phNn2
B4i78mwPMfSOOIHBji/zpppLD6MjISV2QBvFAwc3k8hcfsplJwYMgSwF689TYutI
Smt8HnQBnVhSIFhEjpGw50Jhmofdxahd+U4BBEnZVA/9BLRHV98XTIBkaVO27pIb
NAFfxW1jam1WxL0ojGH32WiAGfFzPWH8Cn3ufrAB93bp6cK155Wb1BfE7p8ESYRi
ggeUsekRgwmms5PSEFMfuSKTH2chluvzOHdyOr6wHns5sWQ27jChms2SRawF4faF
SH5HNo/mnRJ3Ja0sEOhzarwhqo8V8XTsZ0gOlbUt5z4pDl5cFoWiDzPsU+aPiQhC
UUulfLramiRa5ZezbbY4BitnZiJXMQUjLI/BOal4OAOp7aUGNbW7+2gopcpAHQ/M
jO2WAFJ4NFsqPVucAl+h37caXdk1ePQR96z6yjwYLkZJQQg0KsM4Z78geWh//5iW
xfVJDQPni1NFrkua4M7Ipkw6x76rQmfd5PP/8q8XuMB8W5sH5lVIlWqV9pEqcKYX
D/M0Gggom+d1YMEPEBktB81l5vDVJeR1P/aYE/E+dTYGr0SvWXsib6RYzgkiZp7A
PNnCDsaw3Y5l7clC8QZTYf2P193G2mJUm0hPgxG3YLikfdV/k3XXNzJt6/sbqGEr
YWifMAC54OKpnEZeBH+kYgcWB4lI7lls5iAN8nL0f2Wx60z2Eqom5RNwCDIHuv4I
DJQ5LWeBsTMpZ0Yf9TTaRvRQfNH7fJq7Q4xM9QJTpbQLFFuw6KuY0F+gsIXWQ6ia
xMhlKPqSlsv8VwwaHGhD6gpZYZRVSleGZaIRuhjnJD4/kQYimhs92mxbYp7E8wDK
cHFK5nAXMSJmZpk3a/WM0SFMOIYKOe6Jqs78fMpTp88t8UgDBYnYFDmGOjCrGGjb
Kt23/U+rC0tfbzNQQLfnpfOAo4NTPP/u5h7s/rqFH/xEJ7eTsgqK6IEEoVh/OtMD
8od56pi1E5fOD2yLRCZZvqn4pIGSz5bLcd7eS5vWI3ORjV3I8AbxnGxqgScLERsH
EFcl0pmPtzVL0F8u/b0fOjYXf3lzoujxLBXZLhzWHUZu4QzCwyhYEFocLyhJrHdm
ZRNVxPKfLyQg7fAP13p4nRtXAhdiXV99RnyHKPyLdwYLFVUP4CM3lGAnHAfd/TXR
YukC7XBHAsh5GPXoWjYWJRPAsO/YhchyfEEzSztVW1bB1tehr2LqeRFa6vTFFmHv
5WfdD2MVUO0vDjC4p3+kxjAJOmPuyHn93Z/mlJUP9odR79+t3CVRk6A+yFau3aJr
LxD1w1Ok1lbYetmWUqPovJFW62vKp8I43zPdohwq08OBJucFdGKaHTPm0UBkSwBb
tAeBGm0ENT91iylxzQeKwymABJVrut+ixTDwJ5H8lVIfpkb3StOX3krwilfUg8os
X2S/LJ/c6YEsK27oLNwQ26TiE2iYN2s10Wj6KzhWRJ9SAVd0iQiHdp2rXQ0fEplN
Un01+AhNN+nyWQWM1R57sNDJ5vLkwELWZj70ssBLPPI9Q+T03javNSgxPtOCpPiX
csQiyolGqGQ0lM8vpnhhl2eJU5HLPkE7HBIkoLTzdHzoZN93zOJ08EXt4pY3zUJ5
kGHmoilz3xhqKbxVfTQMtO7p9Kw0bhekikkoFgzvvtFUTL67u5v8cDhjTmQoorua
yRBex5ocw/hiVjHsF6wmL2l3GpO4xPkSBGPcCIoGvmhZB2MwzYiRdVxKTQpakRD5
2JfST3FYGvoX+O9bMOWCUrudwmY2cQg7neTCUgSK4WEKtXl6CAcdmmkiOWTK/lkF
PDVg4+S4uUXh8iVoeFSpBewA7hKs00T60b48GYXJxbveYmShxLzMgH9t+OvhDiLI
kwO32EYvVYxr/+I6SUm0+2pNnP0IeCbuDkkHTxib3jWEZpYDRjJOLmksUPYxzT+6
UYcYh01ZdfI7lTij0jmxGIlycJURFA1K+IyFapu5WhD7HSS/qDEfFF/UU1zhWlcJ
ArLVeVxc3ov43d7Yh4YNj/C4bL9yX6y7xo4LWcQXeU9Cw07BY/hpgR9DtJ0+f6CK
Mkcehy81dbWGcxe3QAreRuJF2qPS32gqnco3ChNYGpjrwKHkMTXcvLeCvZRnXvC3
TdHCmzPncsXgt0tDZbXh5SoHhq9o7QsMALqvBozv3wCryN4k0yRZFnHaCX1u2ejq
kdyfMBHjtbrBun5rnFy07LN7WWQ2mfVrTGcSjMo/XyZ9lqrz4MVioHFHpVxtXQhr
zVAaPpMmzOvHpWDAn1HyxMALcZJmCNfqEP1BAGZgVOPB8SE/E/h6+K39YjaEc5qy
QT9arVmqRMnHAH/hQ50Y+PVy6UzNXhecns+UvqBx7HmaCF35Fdj9L73jcli6AjBg
GUUdalDTtxh2J1eDQw93d5/aIHTkEYIv7jpCp7JkKC4grr8e+4Wp8TDsvk6wgCgw
zgXJonUYzsf9KPssnvcvvxWfzsxtgRYrtZmIRLekYoCSP0GxDj0e2q+1AIxZV8lV
KHAtcGo/1+J9CtrWzoPe7kEwVC4rth/+cIuxb3p46Amrq3I89ki1jI/uJZ81zqqI
qPCdA4KnhDuSNU9eRFEyTx9TlDE/wnPaVmmKkbxrKU01tV7gTOJUb5vTjsukgyEW
DR/6j0DFo3ibfTEOyX+tSPhjBNHhJHTkqeqf/HP9yCfIw08vdfutajpyJhc5aj5n
+F2G1ssjQdxh+JDCauFwVXLXDnf1abrsCRukKm2QctsXVX1YLCz4zOkskchRSuT0
csKxbtH+14LoKptLoMvIXRAsURC5c4bLgR/adKL7Bsn61iz7m7YgXChoszt6U4LN
KLHo/mWfVNIZ4i3a1cNVH/+FQXrQHqiD0eGKFSxNcwaJaSAH4mSEn78IQhvVSRwM
VBt128+qcSPUxPoCe3jOH5jocAZPepARA3FbyESetbnYpLDiHSgDVpEQj7zZdB+8
qHfFVL7oZU97OlN5XV0tdT43s4nzMuz9uR87rNwwc6sXmY4zMtr2FtoP6BSL9dpC
5d1fkhRzk401xGdbciRo25w24g6txRzSxnnLR8OFbbgXyVIYtp9ZL5sd2sgu1snL
Ejf+1Xipf4e+B+UDwpAek2+PtlYQf1u9rs3MAkikvS5iRyPShIIi1IvBXMyq/LnY
XhldHlUmfy7PHo1tf3YfG/X4aNyOB/Pp8DS/tU6kdS5Z55hARIl19yMtfTmOQ5ji
oeLS9jSOx3ArEe2N/l2I87WTkLbvOzFDHYEwz4DD7yCxgfZaZKsCROsXgjzjmbYD
nSikmxe847QxftGNBBbCrQIQsFzB19ggcP11dq2CPQYoudCc9vpWz8pyWRIy+3XB
Z1+YR9FMzKQYgM9pBsv/yhfadq7nflQSa6bnuWPFDy1zxzuE2F0imdOUJt1LLQ8G
wByJcxe4c94nNyL4kFVgzefJKVRAzht7TkoByXqzn1TNOojtdwdQ9BJmiIMIjbHq
42ffW+t02zX8VlSsAPAuU8UjODIjmPJ5dakV28VXd+Ykf4lZbr0OqhN3VOaU/C5p
WPca11uNLlHJ0BtE8MHFFCmVWZp23ZAu/ReVsFMEOHQqldKCezMVqlvaGy4yjcq8
HMgX0r6u1Ce6yju/vCm16StYSvtdnnQoVGsoqu1oEe0zuyWKyK5cfIpOP9DCoEiD
zeBkefKVuM8WwLVS8XSEmorm0ppb78g6tHV/qASYvc6wRp3X8VdCU0yGVat843a2
Sy/mwM/6gA9qFYRtiDm9Qm5/WDSK0cnAZMyj0jVRKjcuq96fYSJkFzWRp2EYxPa8
oyY8L2C+eUMH2kPp235gYewCmMi/k9ZnBNbvtKdROJEJciAaFytoPm2Y+52/E38i
flWp5mVM4lcAhz27c0Zub8oTxYkTjsTt7UligAtKA4hzStF3IqRYWmhcld2VL9KH
e1ddKN7s5Ze3sU7uReIRRmZmbmGhAaUKNq3l6ZdG+VUXzORTmpQn7sCmmggNYiLW
hJI6u04ou6934WLTQgFzybTMTzCxwq/si3GLU+3WaK2i9MwdqqyqAS+Zv76BmJZ6
7NinDt54X58l1H8ylwBC3umDq9GJBJgrkzzxxjnr867R4mQ2b2awEkemdFsHxqkO
kzpnOb86BbmdHM6+Om2mS623DmRDZGZqLy+FH9ynAaUpCh1f+5pvNmZjqKHFNPTn
iTTLsZpDKYGM0DuOUkF+hN9/6zAhtyar4SL+2UD71xCbQnQl9UBdVRgixDCuZ6iK
0v1fGGtaN6I5aPBRcVu5zZWKjB+oyKsKZOOdlc4JmJWX5bQq3YX+gfGmP8MMeQ/N
bjuwLl/o86MotQq8o91t1G7/Ar2+Rz4PCvfs+KR+pkZj0E92j5pvwD1xogDIAGfo
0/niAkHCXmjvQFsspGdikKlqCN7hkB0xwNhrbC9JH7nD7kJ1EY4obeMIvvn+EDBa
Lc7O+rOZx/E9GrxoCr5qXzbvETp2ZBg2ofPsmBjvdJ4WcQ7UD6YcvNotSBd/ciEG
xu06MlFTxwu1J9BJ164AzY8VuRhJnTBhRo39nbL3mN6enKwUoGR6RZFgU22U0hIA
qZx/tUUR9HyXLDZt8N/B2PZexaZQBEzG3pdWUL+pzwvd0KXkUl3x85btf20kkcGJ
nbqgS7DqkbiRyB3H19PemTpvp7OIjZ/vfQb2MlW6ThbblzCZzejInOGLY3yZNTad
LOpy40rTbjkmd/uOkPSCFk6WG/gdoklXIurBUMLfz5aoiqJMDlcKK6v5YcRY+FDS
upQdj955gwoGELQ1milgSa9OHi/tBsXSvyN3IjhYqe2/mCaHIdjhvCf0Su+ot5q9
7prkdw57agJm9jLsKdrN+eVM20TWayTizzTUVbh7z/6pb4hkg4DV0YQS7m9GbMdt
5guVXQpcNprkPO4ptVg4YSmSDfl3rvvMPIdONCXEJadYtXBFxwqTL81YfxVp8lIp
CF30Gh2xf+s1st0YNbEEofOAJCQWaMym6n9CiyVhoz0jhBefSsczP44Gikm+piSf
y3kMgR4Acqr/mzYG9hAHowMyWGLkQvkxlY4xYPlVkkaLpibr2f/XS6hEjROp0Cms
uM/gViYdITAlscpMD4V+g6MSNLYxjsnGebn7SMzJP23YIE3kVVeUqTutskfkzEb3
d4cwP6jdKVpb3FzAt91pjt8sromCOnxCIWbBkBirQKji7bP3xj4achd/sP7gcPwR
JypVvT2mI+Ombwix3K0MYjuyqdUFQJ4bpbHGDzBQuNJADJgqqBiZTmy2gtlYzfdz
IvwvzXdfWH0K8hAakfgn6p6WNKM/hTon0TLNwzzStxFFEHDg5mtQ0lrkMX6FO1lp
EbeVTQWCsaug5bY3JBPc1dlEbgP/vi7M3v+Vsvwh58gyUY/kQK6U82UUmzeBE81C
ARLvGaE98NIMDHhCJG4iMpdl90fPjFlsVZA18aMloFoljNRS25et0onMkQzFwt6W
UttqZGF3aaU34DItWdatlvGUP5+gzxzdqd3M0yU+k9i3g0oJXm/xlJhsar9ZH25Q
hCROMydSVnSdJbxHq6wP0GBE8HHEjVB/JZu5LLwiQ+ajjOWnkG9cyZsacDjjk3JO
JEz/WvUQTvZ+Ic6p2XjNij/BHbDPMIE3uPW4KCNzGZITf9o6UkZr3nbRWWAyUvhz
UHtGUOolAzu1U7T+ZMeUppLvQx9c4AF20HSvOvzw2oVgM33eKNdjpQdP3MY8hR0u
0Yvg7zna6duT+ArBlzgqSQ+BtMLb5PIFtEXYXjUfE/5BbMHCoDPIrAnF8wAcitxE
0kh2mMTj+nGpvqmoyA5Q+Xg3Lp336gJTVVVSwHXwU4wEZNqNhq59M+MPvTL6Jkuu
csXPFCBP+Q4SYHfYQVMPgy5JHtqhwO5Ol4W4W5fzJE4c22sTvZ9uteKPmkfozjm3
aMZ+f8qZAI0a/aUCjLS+Bf8vZLHEkLNRO2RuutWpaeWbTJ6rfI2vGRQ2I/d7hquq
VUd4vyZUDXfiekpm5Mla3eQ9bYZfAV6jWdKdKlLQtpkZ4LgESs8ga/GG3cbxVww7
6xcoFAri8Dp6sj03tsz7+/PI4W/9ZJPrZy4kM8vDZd3UKM7wDNkwye1owxXgAVgn
QQJjH8xf4wMftTJP05TjhD7LCR7FAOR+FtDNBJjvPrMXT+mUqvkSxG9aP7pMf0kL
VdMaVtCop4Z8qkcgqmA9IyQjgdefJPEApIxNj4NyXFGrPcbAeNJShsgeXQRaNEvj
ivZiHlstM2SvIdVqCBo9g0HzlARv3a3FquFFticvLIwlybnnlm10CO4l+sxyZ+56
3hQxRlVXm1MxUE7aL4QeOsFVepoAJENEbVPf3qNCZpiZ28YZOAhIeRXxgkLomZJR
5LmtYhu1+Kudwz9y5IlWq3vBipTlAZP37Fq/szM1vp3v/j/Sz/688ENJ00zDunlk
jfuGhpaRT+Dw4fbScM31oNz28Lh9KvdZMUVYe+5qB9hZbM4P/YIMAlC2MldVRqDF
EJ5B4v8SEya2cjiVVtbVU1obaMRSXvw46ljyAeOvgXiynFIVthEGCg5b5hZhhJNg
zXho1TDjHmYsSRbefdZKr+n01NRyCobWIB/RyKVKgCzU16KB5OrCsXqBCyf9UJaj
yRPmYD1PC4rMbkzWS/dvDdoawPY7dL/QOhVb3kCCpIlLu5QTQyP4aBGzvvnAFVDx
cv6fj4CHU35hD2QU6fKngOWyI/Iy95r40JNAdLl/QGu1nWxXgLkfCnw+79woAlrd
6f6JV+ATEk46jDfHA3U16yUbKEOp89FzzYh8d7xu04JY2aBD/raDERuPPFCeRXWO
MRVd+ruwMAjA1AIKW6ZFvzgAD0ctetEN9YpGgf4wKEziKidYtR98LsuvLdojXQ/s
hDTWiCErTTAevkVT4cUMMOpSdL8fkGmkM0oBrejK+b9TgxXkrEGtMD2EWcO/gGGq
wKxkGDgMr/sVYBJooWHbDC9L3nHOmB1Kl184EbJNE/mpzgoi7MbV5d8nG+pzq/3q
FsYkP1IiHzfGuUiGlwkYiL2VPHVAykWiCf4vM9YAocEyKyuUUM/ghelaA3E4cBp2
eZaAjVJia+SQKPvWik6pq8aWCIN0gwM5deOQRRTXwVi/tX8rv8nDIPvHYOY1+Zsh
t/AUZwUFG5S4nFRB8FJhkN2FVahVMp97ry3wjR3gEQE35ztHMBHyEfwwhLsdtGQu
G420K5CyGZyCZl/GiGsgLE6BQsZyKLFOP29aHfMuTmgiocU88FBz5DYT92gBZ1sM
JiNMrSRsiE6RSVfsLJeCfgEau52fSkaRLq+uJ0qzs/LSJDAwyq0snWe+58gAvluN
4BWRkt/LkZRcfFqdFrQjvVmw+F2LytNPiq55DwsxUCmbJnyf544kiJkUonQJ+dh6
+IjccOpnabaPwLks0hROy+f9S0Kywn3F0pZrBZG9gj8cVn4P7OJD614XDPVUe04J
aXGXIbplRif2MvzJ+Bgq80p5ChkT1MAL/S8HNpHwWsgaB0dRFOV6eePNVJKBZzWv
ZiEZqvc1b/PyvxmOyWcEqURZ2ksXFGRjw7twQvB69oMVT87Ukjhng5RnOxfRHmRx
w+kfMS7cLMp5YUKHRZ+S8YbtS6vWsM9L5yP6TNO+aVXqr/bMyy0hEjQvI7IIyUlE
G6p/rbV0Hc0cj+vOhNJ2mTgXiwxR7mD2/mb9CxukwXhmv1DJrGF7cRTMp2pmkHDT
YBTBcvUQTgCjZK6dXd0lvB1SZ5Jwkv2TyyJosG2QGMPjLQNyWwgLrfAyNuEvVb+O
dNNjNfTgI/FTM/g8phdsUkdsjDSCvbCYAtXm0Hw+JYBVk5mylYs6weVWX9/gO5BI
eVjgQRqKAyVVQfF+vJox7EqYmk6JoBMviotOtUqYEPbwoDDMrUnGp4hKB7Rw2N6w
WUKtdOoSu2GuXlsDTbNJUtkcoVTLWsdDl8N65ynypcDypiCc8ZoHUMd/QGZQp8lK
8UkLJifJxArOjgtI//C8Qb10k0jTb/pqPG621cft/z+LzflGPS0hvzr/zAbkMLbS
YpkytgvP468FzRIIC1AA5Bu0ZF3m8WPO0AITZtbxd1QQ+uUjY44O6M7qD7PMIU0z
CHa2BTPVRlFY/7vHA1vdYTkjALeAWswlMimWe7WaSlpDhOUzH00rT8Z860HogZp8
vreiFurtUsI+3AryrwdUAbeheScz64sZZifxetY5/frCpebL14l1bqSGX0nr/iZF
qOBfIjzZT9PqUFTLo9rtQdy3OI6WJt+YxiAioBSEpA1x7QAAFH28ppyr5nqFyi87
O5zl+PpAfM9sJEu/mM5UlrNmLYxIkAA5GYDGsIx4q9oa8ltV+txZ8TKshsmll4Hl
BvMDJHhg2Nh4qQX8woVKS+CF8IPA0w0iPd4RZcdvqTbwxKIVXFc8cNWZTvU6oWBA
mUZOF/6QR6v+pTS13i6BdvAozH1hPZucdDP5AZ9WHG3hcX+IYDwySjBRy+0XxTHy
B58SqzUkelv4bSPI7Lrj0UuO5xfidSEdEep4Ejtkya19szeG1qRIXrhTUhYI/r3g
k5hmyhsEj3J22d+i2WgQqA2v3Wb3EOrQY526uX/xUkmuFibggs9SofJpIdGUd7sX
Y5BfA3H3xgL+9egJhQ3b15ZZKAqi4qU3j+vY0KwztHEjaB7IaVsU/w+aDo6/+Xuu
FBNkTEw8V8tIygoWxC5c+DuH8P/h8oEmTLGWrjeYXhAX7RCXlXEFZKAgJFZlzWGD
xJNQeqnubx1lK28KFWOJCTdhWmDyMMRR9wcFzuIr9v1LIfhQaN7u+pcPfFuOUMLr
Q+MSHzMqTXcDhkKSXqneeKbNDG6bChrBKTW+BI3fmUvge57SQ7hx3Xcc4+uHXN24
k+1Vmo5riGmC434yTx2g/9Dcjdz433oYDSOpvsGCqVUXDaxAiJdIbu3I+opCIQxv
HZl6K7h/Xakf6gZo3Lcra4rwYvL36pDAVI9PTWw8+bOehvulWGyPhoOIvnrbxdGR
He22FD85Sd36oWlp1JDKxJi0k7gOZLrVc16wD8LiTbxlSPLkx+FWLMrkEnOBke18
gM0jn+9EYSRhgQmHZKuktKkdPSz+iqF+p0ErjvDXulFBd/OHkTZVpVj+WqvVOVUg
20gS+BCJn9KJunfpaLmVOPENY8Ji2czasFZhsd3Mk0+rvdZIJLJJ4eQNtpAlxATS
ut0F2xEeaGrskgT8ovQ+6Y/bY1EvdAqj4EFdrllxsLhSmaLaGnhfIiXBVnLutogA
fxIPoL2K3bBMdwet1zdZfejDRioivh0Mge+L/xfavg17ywHLJoaeA36ZXWU3Oj0B
ABSiosSwdUiRzEw3ftuAY2wFcwHU0XJjApPjpWM65KEbmd8Nw+xb2zaNret/s0gh
hrFUJAWdP4jk7qkHw11EXACovb2iaO/yowCYVDSCJDP0GzpssnhqTmkpFyHNI95G
yAU0kEHQsJzKSmHVj3LeZQW5ogEvCOWMOT+4Z1TBAvg10cAGx/tFAnfMpaQAtkki
SBQTfRhfbq4jnRXl2C84On8b4DHLF6kYdKqoVf1W6YDMPhPRZ8kD/Ixb6p1TB97E
H6KoTNAist3rq2KA7Mcm12sDpPpbQiUMdrl7dA92wHqGQ2PMV3UggWiZvJ19lyMJ
1on/SKPlIL5Nd1rMvpCg8AGIpew0SK2M9PrPY00mp4mFh0mJHvnbcqpD7+cPMQwl
sLJ7j+kVvZ9MvD08KYnxwu7kbvvDA9mkbDnzPwj+nhng8VnWCSMniXd1805hRZP0
ZSTD0pZM0nYIluMjbySIZtmxi0i9T6fCO6nTbbZwkjQ69GItMSuv0r6ZaeoR0S3L
9Y1e1wubPikv8GdWBVZutgYuZyw41zAQx5NlqnoSpSxKyDWRzOkOGuO1tC7L/vxu
oQuMd4KVfEYaaQ9xhwi3dWp4kxmFGMK4c/cJ7u3QoNZSL+gFUop9w1EFK/6nj78u
vcz/mdvrMzAiIQ55feAtm8NZ8QqdkbPsmltou9RfKPy86SLvp2m48fgi4GKihuy2
89tKUq19JM985E9T0tTxtDkbB8CvwUcqHlTMtqdOr2z9GsU3oHSERCtokciGMuVc
5w20Ph1FD/WiyzCp+eWt/xUPas+fJU/1r85XxETCO2gKcSa3LjDqTAUtr0D+KuJV
0IAh/ebEEtSNxkcBssl+2iMjfxNh8gxbU9A27OuPiIkNGM86VVO5JAE87fLmiP4g
sPNckbLpZH6bad5FFIuwz4LXMbaphV9c+o0WoSvCDqExBMv0XoDRUbeDfGtLCIuV
XcqWOaEIb2SrIASAPxSSCeMvkjZ/oRvp9C3G77yGf9oCwf//D5StmTARTTTftoSl
oFwrQ9GPSAMg22WEUrqMw+22/B4nFL/90HxvNzEg6aq3qTqn/SUFedqBGsHWR/Rn
Tp1uQwP3qviQ949ON7RiC3IwOCgA5+pXyU+fFJFzA3JhnsjOy4gQ/J4jp/b4hFgR
M2R75LwVNoxmLc10TkUK5rj+9cgtWB24JygCCu/fIQVDFW5TDlQwbkBxNsRyDVzb
iGz6wOCMh3KyyIN4xNMQnl3QZf3x8SGfM/K1N+YI59g1d2bIENYjWvlYjdqXM08I
QLEyMUoVxhxgK60SSnZP5sWH5zWhvq8HzuKcyDkbHCVdtamUZTyIYmQhhC2L3wsI
XDUrqWF3hgZ9aaMULZVxK5aiQmz5QpYqHrJtlICon2G2ky6ctfESbNvCQCKMnOXJ
dE/2IbAM8EuyEhrV7aXgn5zP+6YMpHyCAFhnVTNNwOiLtFJVvu7orMSiG/lop6NL
Q32lonu3pDj2tFlTVy9BG1Lo520DxgGonDyTozGhc/wlDRUx8xid46iUbtonyvvl
zEf+8I5VEF4y/MhWfwWwlgNwSc8K5/s3B9HVvmZOHSD3sGdxfVyu80VvWa93T0J/
Zb3jdncueQBF4iXnS0E9o4/gug+kAvZubEQyCya7pvXnm6a2kIUQbcAaAaqz/ZFn
S6ltqsTK+aNRmpXwmu3SYEtCuvxLmDWIzECs7Hfx8rEfkKyxUcH5UGzxoTDbdKYi
1WtS2M9/b6/g+XFAju752eTAUOh+xSc4q8DP3PMlCB9x3IUIAcrxnWLj+1jmEGTy
w5nhdKzvriwAqfe1QqoGrezKIEEUOxj7vCzV6an2AdUvTTS6bA78+xCKXNXirgXS
085sH10rbNPwfGPX6/pbsrOwdsMZOUzkBWIuMjDlI22B50MPXCU6aYqGvilqlPrI
LfxjfjM4A5Pibt/6Fi2wt4ufhRNYYxA/ZEKM6jFLN0YMHygnmiW7ylza+Z1pRbm5
jIw0SV3ADL/oFTWFMf9w/wn6MSOs2jRIAsbqeI1i6z12NGB7JjLJb3REVx0spocm
6i26aFsaH4uy1s/zlLx7SrYexTQDoslBasSMHxtXlg3X+01C2VpAyKhfp4BMw0KA
eTxq+ZdTGiMDwR9b4jrxzD9sBIN2+BDVaj8sy1XKKj25GqKsdDu4ZdvTugcIXMgQ
sKnlwes6XFdwEAH+OPWQPBg8vmchCzuYL/Ny9x1vn5Hp5NBaiTOUHruJUtlUqRHn
SWF/YJiL7aU9kvf+KR2jlWKEWGEiDEPajc+NmDggDC9NYmjzuBKJVhM12HXZlD18
MGN0i46ItQzENK3NqKMdTCgrOzcYDzj6Em3Kcwwpra9+d4nmfVGrukDdImlCPtTt
ismo0EbvjOK0x2ixmouFp3tuI9QBW7WNUJCV4rF2/vyepUIdoINkS4pH1ICXTunV
jwan9ruf546Qml0LhNrqL360vMzViqRwIl+IBzEAhNu4oG+kqauv5M54glD8hXMI
7U9T9jdMyrfkEJOUxuRaRABalQpdmRy6jKOUFlnfg6L1MGeTYL4WhprlnD0llVQo
KwPC7IoDM3LtelFuUkMxmii6cO+lE3R0AsbbveqxNZEFikzKSNpFP4BZnmuXPX7U
VbICMEB9Pilah5cqhmrrcid0jUtOFdtMavjNpcXsXvZNBsceZR6AKTN3Jx4SkGNx
f/4fLXeaIwtNRB71gExjbNjr7HLiyE+lVU9T5fi4gwq8pbJxZZs7kPHpHmX/B2lP
BHFjRbGRhxDtCxNWN4QIEP0N1gS5nI581KXg7f5Ommwfk1+dqOXF1iZZTzEIXQWl
9rrx8QgFUr7MIW0q3lzzBC2GClTVW7YF+b3kwbaMcub2yUhDnPNQINg17RBKUuL9
TIuWsjYMtyQZUivFYPWpzbcCOHLUBDsLcW8KCckl5X+nFYkdUajaf4/fdwZNY3J6
pss0gBlhKEA6cehJS8pLn/QMaMDXXeQaOblwOyGnpQZn12epcfLlihMCrXXyuP8A
LATyvtGYEaSjx5zvRWoigViiobaT9T6By3Qeqx4w4xVttbbXe2gcWEobbrjgbO3c
Iq9tH9DFXcK7VgZzY19muycUpI5KKWxRzfFGEZChYzlLxKMHei0fLE4n5GBJkVZw
n6LjLYIkR9qOMIjpY5+DmOpA1o0zx4JrjCdqTN9tlRxwJn3n/cSbggwGsWBGTE4F
Ieu8qlJ4IinqcGulBJ8a8O9dDZS8ZuRubu0XD0Eg2946hsJYh+ZwI2dBVaxmPVZr
O4f3FkJem3qNPmirMwwkXYawry/XLO4R51+vPHL+1Bfx2klhk29DXz1vimA7owbO
iZ2Jfc5CvY9Wwa3nes9KWbww/Z5mLR24qDlW2tXVLTUv/hx1+xkA6RPJ8cDYLFWu
1mgyMxlx4pQZg7iwn1pJG5H3wK+oKQq8fk1JmYCNSWd29snUVquoaYpCNvJRahPh
DlwTrcxh0p+tjeVbPoZZIiByavk3GGsV0i4h0CGQ2++CTPLCdEfHv0oEZLKP/UIm
lWvngxhRySUKBrpGFdYQugESlCuJP5HzEegYQT5k5U7GScbV4B5UfAtWgP1hBz99
E6DMRP5vQHq/kB80eIRlbn4tTDPhFeYgO+qOH5tqrjPXjWJ5JeCNbpXmpC1cgWAX
pnLjejIQbgvD7a68B3J/Mre7xKDeh8yL3Ex73A+qSU7TLknoA86mXfHbJ0d8+6tK
Scipt51RNOq+EAIpxNBdgru00nVKWuLqSrjlbDfMvd8hqpNawNKH6yW0++Nn0wf3
MoqO0NPJh2rckmQiVj6CwGnBWoAgDe8y5PT/NEVYtAxiRj6iNk7sjYKEL0Wi8Lk9
RoJ3e44rHXDeXL5laGRvG+pttP7dLCyC3zrIVT3L8EcgMfiKs52qxJAIW00lNIW8
vnaZmrEMJH5DFT4/P0jZFbOxEiBfzJI6jjAj7MIEzGePyahQF9phM0PnM69uD81R
gdULcodLjMVgmE/iihgbHD+zj3d7A3ZynZHV2HXx/yxbPt8wzEQCKSvDnIqvQ5e/
1qPM1tBAuSBjstPdVLxfckx7hf1izJVfHfLzv/RQtHkj/xEU1CG7nyeG+sE4t5pG
e4OZWNKp81uGuocNbS2feko/yINheBlbWUkaZHLnKSdEgk6LQ4zVkoET5xMWW/aH
HvMUbCWEvDk7jqviP+eMtauhEqT8FnDFY9Y3T5oF3ZZE+rhct3WrP1qfI3BIiixz
pr3IN5x80vMV1K6eotoA+0fb+vKaFxXPBZ1W55Pdru4Lryqo5AIDO8amusVM2gRr
WYDPkWwtoOpiFhWS65D5NoAM/K2UTzHmpHnVI+lpQtaBlAD5EwyyG14nCYqakII4
r04SaCbRNSXMCbWcqkYtOHGairijIxqEuEWs9z8Gk0piUva3SpssViUkSl1tqcfd
t8pe8utzs1mTm+3r6KKl4cRWuJCGxujcf8dYsvZdTiiCGZGt//wE2h9QfgwPj+eT
tu4N2j+ZtHmURTsxpTdo/2CzlWp8SrB+c5ZePlNKloEy58pEDUc1yas/PBiofwP0
39epZTvAndb7B1UyPbYL6o239vnzNb7a16xfBh0YxOW7buIN2/TFNMmC4ACs4LdL
YIPIpH6MGXSqMezlI9Tf/DIkWDyDBWsG3IVUWUh55Jtt7nP+7tL/hqiAtEj6aqII
nqg2HEfM2zxTXrh6l3qWjtYiRtvnm9YYq/bsm3Li+JpqdFIttJjmbt5DhxsRmnzr
cRggbsSLMb1K1DQPTFUnL5fwLhjpMnh8/Hb7IFJkc/bkP/69bbmuG/mmEZn4hGjW
8kYJdHU3lBPxpOki0BQZDKukeCK050T8B2g5jzYyxl7rlFmB4DJ6mjHrgNtn06wQ
mx8bEnrPzGk262gF1XxZ4DP6W/6t2v+QmMIn8rCewBCmbAof3YU9SNvG9KhCbWUK
52mA1w0hREqHrmoqGHq/SCyLRdXrzZVblwpW9rZwxU0Jv080V8ksAq7Wc7fr1t+1
Lr6mYELfYY0RIRwt+sONBFPSw+PCYOyAFHqV2H5Jxs/Z86mugDd2dvLsq3H0sX0E
sK4Gy6eK/uL0h1Yx36rlisUVrw8b+EtahGb7TrFRd2YflzSs2I36oFbLlR6kxIHP
KFSslr7f90sh8zSLhfHn13bIggwOY40/7d4jDBYs+LQHKnDxd7pmk4/Ur5aCKIlt
J4kPwWz74wAakaWk+D/SKuU98qaifMhnngXCDRS/P1ukhqw5Qg+2MH+r0qL1XWqZ
eA/sjH2Q8jrrPON6cghWiTxiZS+ioNdu3QUOVEz9lIX5o2zihI6MeIIrrAvcAP2m
huEZfbvUJN/YRJI38L2k/NtgdIS/6lS5ZRRZM70BMnOiZvW10oj2L1MU8FJGne7N
WPjC/k52y1vWFxVBbIJf3UipA/r+2ZPXQ4uXetahLL7394+C5Syv98clVAfJYOVz
TmK4O8tUkONqxxpqTE6EaBhYUlhVB7sY9nIJA4Hw14x/92w3XkH0cMbn/C5YKg9i
1qn0tUbcwObi/3KBFnMkNXoypO/7i0DEmxfTV62SEFt9FhbxGtthyQB7uYgx72fW
uAjebZd8t1j2kC30EUTCQ3ES2gSyjxbn1TDMyYUDWbVy/Z2IjFCtS82ahpT4unFg
tsy9g3HJD74BOAsTQcY9hzc7DYHHGJMaWsRzBaKsH3+efABSMmVFxycFYD7VZzai
X9GGIqSQYYm7CQf1DKSKMAbCw8Yclw0+PioO1WuKPSm/4sacRo/PNsiJjYpJGzZf
P+7ND7wZsKxlibyP4twW/XsDBl3R4wpAhP9GN6U+L1l6UsRFBGveHlQOsRPPrgD3
2ogAs0hdFSKW8W+7tLoL4hD+nfYqiqOEE8zFn7ki6OGedVbJo18l+PJLRkAlFJb2
ierhy6EUN7Geq5Vq0zM3j4OUN1ezGDyhBWheGYI8FVK8J1NMvUBsryFa1Vs4TCvi
GZyi6d8Qo+OIdwQG5mJhu6BPmJ0eh2XHpeiiViwy+knHSpyeQIw6fLqpU5mf08W3
EWsZuk6bFR82rXsrloI8Kp8xf+4L18fxnRWqIufCM4DbN7T4H5EgJGUnTN/15MKS
hXQXUmCagxWkxZIyOPbojVemY95lnq4Qq3UttwAOymBO/gIvFCoAsoM2F4DYVsxj
b2ymxUGKvODjD1FuWkRvQk5G5QK9Z+odwcMDjlR9zRFZPflyJceTaTSvC3xBibH6
q0sPJu3qOkuDxBiuO/hqvo0nWvWvYI4veLjeRNY9QRVam6EaJ6jN4HQzxYu908hG
LEfNUkrg0sE3Tf1lswIbwmDEPlbsn1ASJDzEohIRBKBsc7KEHpAjk77a3ofDYqmB
8C+eVZk4Hj2FndptrHfGI5p/0gWfUmz6rWamLvu0EZKn1eThe/UEkFSCPsVj7BO3
/vroP1lofwE7iDMFx9tDfezYv/JPmjtLIUill7gWPzE7QNNQ9hPFUj3fAq6JLSO5
DdSFaiSnvae5od2I5goDLEJSg/EAbnvbF1CB8WHjBdQXu4/QtSzOixnTF7lrsATl
/F5kFM09hqaIwhdSAiphmmZAMTnYX0t8bzOgJp3Kbcl2awEtxh2jVGOPgIVgrIZ0
RdKqa9hd3x7eNM+874G4Q2JpRAIoCVuEgnoI2zZarvR36ZXHGCjBs3YXTNPOuE5R
9NSpw4N7EswByLq4/nUJzExu7aWpA6QwqsffSwSc2ivc3rP0QXIuHypj26sP5Rn4
mX/zIHzPsaMqM2wOhSxw+Fjf3toxh7AFOrdQhxRw9EWnw82rd7l3n7npchcQFCZZ
4rAhf5GcyvXygVn+hd8OGoS3HYVC8tiTTQ6KTYR+bfgCdGT3HGPfNI4OMBwooxto
6AJM7saSOu5BX/RxUxzowdmyJZq1rI19Wlx0q3bGuaSfEIu/bKZh9SWyfoBIsWFo
P1AyeBsPRhMbUZuy4QiqJzKybzg/VG4cd5pa2AEqaze/HYOF1s1bz562an1z/TME
7vtRhadwRD58cJT/ioD/2DVDI4PbXwErTWakG8PFI1F+VUXpJZI7ORs7T9uFAB98
vr9Z/a71l6vt3uaK4jRu+HmnDik/kFkKDFHeeVv2xTWjF0tU9jLV6BwzbDWcxRJL
6r1Fh1Bb6+GggnvC88rAjP5jcNn3VbZgkVYtay0Y+iE/pDbT9gc13KmJm9XTTttT
JiFrpqZAbOU7hAkxkAqis32kMP5M6E9IpB+laEb8RibU4fBc5DPoLClOMQ7iGsDu
DDkKtf5s+uA4TRr59QwJ2JLyWUsotm7K/LbcOoWpouXYRKsYiF9vF/ZsFSeSp5em
VC1YNyPP+9aXjuishqWjyaZQonhsVbjz0ZtVkrKoC0aep3vEIEdHiFme6lxXOw7u
pl2bo1fb1UxCjZYHRoeC6x4duFclGeh6g0FfZaBjJDBr05z76LAeVZdSRK93eQaK
vpj+MTqP4ty2EEOamVb9owOh9XQROWEdhLbN7Msfl0KKJ+Eu7sx6Bl5BCwUG+evN
b9u6Gr8gk83gEPaX2ypjki1gmEl2qqc7JsxxRHGJK+ybtXZOloPiLbKDK2zQGOC/
XufhgOu+0nj6lWkTwmxFIlb2twxe8nL8f4WqmkPuMkikI4P1l0fVnBkHTh2bRl90
TeajAJ3gIK/7OPeg+YzkWbWWBnyZKj1smhxQy5X9QfqQ9XHQwBN0HbmLgu8cUww9
kEM7sn0ZbPHDyD21xkHOvHQB90AU0ud4s2SlEl1h7lisueGss8ilYDyNjto0w6Ri
VqU2E+8nEqVN/Wx4U85vnvE2+ysUm10PXs/XqbJ3OKGoWK8KRYJHiIBD0RoASUk4
IzzvSHuFgoaMdcX5lvbKBOfitOvzCaS8ShhciJdPNbz/lhRo2W/2bF6RuhRFfjST
0PYksTVeuE+ODtDqnQDPa/NT38zNReq/or12uxYaYc+ybz8Y+kd/2xN0JQKBp/Bs
O0doCRVW9/AzdmrzQ5G3N2yRS60V5QceooZbGD1b8AaA+mIeyyuvqsXsSrlM1lmZ
SMEP6/CxkH+jjmnvpZ/YWnjDivPmjBDfazGcp8pdHdzJo97dlzX6aeStw+dsAM8D
/hVoGB/4PgiRuFKWSEYJZjCzdv1UJ33J/hQpwxQ2/G/a9gRgYIfTEjQGXfo9AQyI
aZKmVsG8LeOud/OsBBEcCfNoTCWSEbgguqXuBPYqJ8k3pto2d2egFoYECbzace1u
WhXJWxCX/9t4+LfFqk+Kv6tJv6eHFXBcWz4x5QrfAVkV7M8KlZuCpw1iVyt6pNNX
SGXQdSAsVD1IJ937pnVY4e0LX78e7sN4MwhQYcP454+VlqnBNozXBmP2ODLO3Suu
/FhK+Tu6U82ItmyhtqPpdWDG+H75eJ9+l0F+k/I5e9hXNr7Q89dx3TYjuyfCIviw
ec+avxo0mBXBCCn6c1opFj1LPoJd6z8bf7Odv/F61y//OrmRWXr7y/VKwVPMDoiU
LIK7PGvQ+zO4fSsEXvlMyq6kZyK/Tmld/qejB8GS1iA5X0OnGw5+Ul2MSnU9HFWh
i1yvhGc1bRvP6tcyqso09TxlvYFKub8jJ6bSV0Mq+RIAc6F6hzGNKn04TLoosuNh
iBzPUsdfLTOwz9kyjqZ1jLFEuoxW+pFKjDSxenXiX2AJ2rCdFkPAqbsckgUVLcSe
wFoe5Jx1uGwJlLNJ29+gMiKUU1Gl16cDC3gxIOUM3ntn7EMoU8zUTgoR/pEtGhM0
y4/nkHaHGRg41DGpd1O6aTekuWng5kOdWi/4xo9iviatKBcntPzhRWSglB1RzgIz
xzWwz8JwLld4dTbGif38cnJ6JYpfAHaZjx+XVuuXSICvZYlHEAYW7e0dWwkjf5yr
W3XOO/JEp2RYna+Nd4Dc6/XwUEVbe1DtsJkPESRCZEvfjosjPGn5noIzhKkBc7B4
x7SixKAHNGBQi/faqA+YcP5Q37aO2FA3yItigyUm2/EVL602euwEBvlcElPEi229
5k8SeM8SPG/Be5WYLsQVMON70lsQrkK8tEBBPjJK+bWlNWFv8luqWSjQ35yLnQmi
UPdLLU9SEMDed1lgjuv6PD5U5sFzJjQ+iDb9ETzhJm8Ynbh/4aslUNKCqf01bmDY
xk0aVD2CXPtd9GhKxKmWeMCduinIb2dr0PsgYmzx74W45QVCnfF5SMrz4dkH2qR0
YlytGFjYTesHfIykKRqJMb5yOYFBGsGuTsnmbSHk0Bm/DDSLymY2TV7WAp970wfU
KqEBuIGbm13ApN6bbBnVl/sF8JQJ/7mg9DhhfVBXdfeVqOZErzpPmubzNU/kfZxn
cKI7Zfufwopb8ZZp14ml2mz97UYCXNxYJd90O5RO5BmyRPWuuN/eafQmjk6bg3F7
mAS3S1sgmENEf8kwP6fM04TA3oF4NAz2usY5X/0K5ot5zdeaMwGzuChncOoIgD7t
9x7Vk3UbSx9I4W56rJTD3LjXunvxlW948IXqkjvBNBpW8Z5oLZif73cg/OMfvGof
TNoCzKy29SJKUrKj/PUB4qgnUhYyqaLZn2kvWiu8PXbEzXeQIpInYXfmS7t2V0Oy
veS13s94L6Izdl+PTM07GS5VBsMh8bKFtoDs0MdfpWJv4BoNYOoPaXBNWzr8qnSy
jCS6E53LEO90qi/Bc5lAT9UNdUqdarHu+Z3h4fFQHjVJ+TkTQdSX437lb1rN9sQR
aHB0XI/d5aBiZK7XQIvIWBorQAnY1pg6d0A1DzMGAAVm8Qsq88T60nGMRkeKLXOt
ZrNmjG0EIV2DB0SFGuRWxGlbEE2HY05AOcaNsvvKiS8hANKlVw7m7ZAZvN4XkI8b
dFmDTEfEzPZcXk8r0d6PMxqrAqTwBVWqsraL0+mk4AQQedmyWAPzKBM4xLtXkHeg
6npUOppZFBltwtJoIbq6tcNG4+Q1c7H2BcomaJcCAK6WRGroIfsqsi4j8nRhDmoZ
ckCAyN+kvVkVAsIMK4vy1PjadtdrzVjGSgZFFrdMkdd/rM6yQ3tdtpCDr1biux7y
cVN6pyF5V36hHfr6A2g5P+MsoEDkXM/Dr+AHTUrm7GLhS+gg/r/4x8O0XinvhRQW
A9gBb7yhNLKubpergePYzr/tO6jSkfObzgntftUHNFG8HOGYhpfBEjnFSyp14Qm7
Ad3W72OWe4RR1hZddvnxBO2KcOSnhtOJSkiiRyjA7HoG0YXL6Zh5u7t67DTRDMSB
fspT6bozOesb6KJrH8hvitbxA9flUmGkJBPrKqkJLfU2HW3JNNZ9QNGProJcOZa1
xpcy3ugIj8l9lRqSwOaY1GX5SSujYHPOHGCMCReuNQKfEyEOPY+b3R7D9Ej/zEdO
m9QzTdV0mkOzmY34yUr0/wzLtfgcxxdA4zPYzp7yv3NLV4LOea44d4zItqkebG54
uyAabC77h/uhC5ViVxEmGpa6giC1JlrEtZHKbT9FJss=
`protect END_PROTECTED