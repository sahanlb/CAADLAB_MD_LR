-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dnefGXF38bWZeDItqT0l0jLll2pkT9wdtidJEMWk1N9yNPZYuAV0YE8JqL32er0DARNyjOiMlids
qeI3lLWy7EuPtNQyFzQDJRnoNWZFqnWH1icYGrogY1QqooolBH4d0oaq4FB1Kp1AdbH4cMErPm3D
UUMPx70reZfC/FPEjl4Jku5M7ACGGhxwmPDtKGX2QHu5eU5dYxA7f+43kZUv4hPaw5pG1apNo1VL
8a5BfT4vFanQeGKMIt0iXD8JDBe0J57wNDWNWALE9AH5wQcj/TAojqn3es9YCpLavqLuqyLdRcOG
QQf6ZhyGOmbH1S6b1LWKeLMHc/CcMe0msswSNg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
esuCpBmYR4qPf8tKKaP9L+Bpy27N+sSjuO5Q1smOToO+TgNgc9Kl3L328p1cIH+c9ULCxB0xZ4yn
rPyPcwM0cMq0IeU0DYaPEFFmOVzT6I81uSBT2d7r9XhGSQmaxnA6vMwXkaBzrSAVyUzBEley9ghr
ODaIWxEPTTzy6SPnuxqbCTk1eY4Vpk4Ro7QBjaLFrdIFA5VuCzUzgHDo1a9g+fzEYQwpJ6dp5eYr
wkD8ON9CDiluu0bQrA9tRIZ8NKMEz7rf700e8jm3I9El9Hh83qOOFhkex8uzuo7u3otxu4J8cAKr
hoq7OrUUponzoaP2muSwkD3VcmiYotnU3QPwgYG5K8zZ5RXrhePXuv3oSgx/Etye2K+1/IvL4zj3
s9+STTFsg0GNJ4ya0wsk3etx9cGCmTzdfAV2Q5+3+jTGlOwefIDApdxfVPnw/1ztkVHBJud+lADC
j+ekZnJp2QxTg2nWOD4/N9l700s7KlUiyAYZXVRZtUILxm0pMni6BHP+54aSagAQC/2qGY2VHC51
RRI/qaobmIeqSeM9xqAqQcwBmRx+hGv0hkpDGkt2yaBtsG3FjVyeTOwVOZjAffRcdLZe3zi94dBy
6VQZ+F+RtH7N3zx4+n5yoWW7UChQ+HJoj6FuL/Ryaz5+fE7rFxlIebtJvE9k0GraKaxG4ddbmFoA
UXaIEZ0UBSxWg6iS+3DmHP/DyYCysUQxsJRL5/UipTXfuTyukvtPQ7RjZnpHDMeviCgoEwEcwBC5
ezsWmjmyp+wuV9TuCq689fDUKG8ARsbXuGNfuTpauuH51AQXU//ZfxnzDSUmE0nXG9DjVbBFBBZw
zwmKQBz+dkWS1DeKqelwk7ibRU10RwTQVFQ3b0CtC7B4x2lzQ8XB7NG4GVO9LbdFaj9SFF1mSlat
8fDopyK32BDXGGrtBMPjTjKZO06x2ZfzJZUuC4uKc/6cLBueToAn7JdwjS3aQWs4NaNkuWhqa3iW
OBnyk1AQj97zF0ZCrnEW4waHGoMJqlTNMNtPC2Wm0lve7ZbJISdgHVt/4SdAjGvg2az013Ha5wsz
/ZavHzNQUDDkutL2tZwqUo3QjGXJbbxRqgPI5MJyo/x9Kk93mm2KEDV2jqEn+a/iA7dqq0Bbksyo
arrbl6dV9kdw/flzjbKtg3Tnm2r0Cm5+Vkyxj2IDOR/Bqm0Ku2Yl8IimsQ40kPPXN5JcndWRkswV
uQ2Z3Emijv/wEmkF/JIcz2XmsHZgCKYxpqnvd1WtUwUbs2f6FNFHHsq7ABh1GJkfcbx0BX8BZfBq
u3/qN4RA2jV4Vux7R1Uo+zQPaRf97HFhFQPbQiNMwRagLXaQGj02YyetFtMVq1EdNbsru0VY2AJn
poibuRv7SRhzXzY9fVV5dL1N8CKspfrAue8zyAsqRGbirBLs/tG6HUmqLqXyNaYGyABMzh+vdiTp
b5uQ67wAle5v3kyn9UZM96TZ3e3m6MlbKary2j4bCTmgazu/60fyM+g2iOl8WPL65XT8XlOfVEl3
PXqMmW3DR6Imcr6u3LnmpQokrBRwAbO/gr1AM6dE8pjEqUJEy4z8QbcofCNljCLAnenZS+pVyQND
PPhzJ+XB/y8/fp7tryxMV+KN7wQI0VYZ+HBDCFPEPhPYMbXqLCrwVDq512En31J8kL2kP2BpCyaS
mH5WrZPmIs33M67w0sxgwkD9jQPgWi9p7ShPRzOCPI/DL9Y9NrQwXsqH0HQhUJ+wQhsSg7ZB3VTn
g9gVw6pXGRY6yQk4K0f2YJFNyEMLHU/pCDFmWsjdFUSRbVWG4mPoQK2fgdOBBIer4+BIX2q5qOMG
9atdPuCUWRYHz3ltf9KUbu8LAJQqgbxl54u/JWeicLGrLJ59+YuWOu7R/Iw5rXo7ExyYEt0WR7uQ
H1RT2IdSZ0RHjX8CdGU2ZKk0xwiNQ4Olyc3lexHXFU1JKYfoGmVesHungYG89Pg37Qg6ndR4e++n
Ne23BeE4i5GzEM6mcdBi4BT2mSifNx+oVCPV93p7JHXXMKrhkMKH8vqGWLdaafhYyxSJSRoXNp7s
uV0GpkYBaYVAmJsIvTr6q2OZFqYmh9uEgOgTfAFTz745b4dq5Ei9BwRLv0XaYdLO/9SzEQGPRJuC
0SpGewKRmRbiXU1q5R4HLmcWNUUS8Cx87M6cbKU3vwlxziPGdbs/5i/P5ngK5veba75qcsPKPLCV
nkxUmwBd9fFX55c9QzJvQBFICkPG1aEBVSCYIG6wuBzPOT4rGiG3Hjuk0hUmN8ndEZZ3ZjW4Lsqo
Y9/wk8lAk+GmO6zQ5hATnoTIPTiAJSyWQLzF12s794crLhnCqoRSt4a32uauxjf5SszztVaefSB5
YdkzeN7h833J0cGVcXvknn7rw+3uOZ4f5ZnjwPjizXrfHRLDl4vqU+i20cE9cG82qFclslFMViDr
VRoENuCcw9eSao59TxQBB8RM59ZxBB/mpHArKZ1EZ04JKMgNrgNjIFtq2Sm+aUWBqARUu47tcg5V
Ow340LWkvWx/FrHvCdcr2vLK9vKrJHvX2hIJEFKSm+KHiArw3KZFrL7O+PsPOKZr9Chz1yI8kJdF
6B9DCX3Y/ATE2xI2u8D+a/Ktx7s8cPLHg9uuYgZwfxSsqE86FlFaT5atiUP6D6FWqoFu68BByWYU
l3HPlxHgnDRFHuXqkmuPPDUHJzpzxC7/BLX5rD4eHAH8u1oGTvuoXyAKlO2p7Q9zYeRI8ka7z1La
H3p0nqvdNwFPv76AuNKbcpKB4FKdx7XPxII+Q/fQRcw1p6lm6gkhHihYYVwZHLdx5TQrRcZ2JbEG
4+EwekayW6y75rfu6kPIpy0DIRY3ola1UWW0hhdRyj0Ih3fSzhUPOhPAkGHGg4VIRK4S8eN7SdlP
qXX2DnoEKz/WgebSlCH6aM+PuW1WWCaHnFbdqNi/GBMa1x88kmLy2/Zq3kyiL0OdxHvbGPfNVDnz
96ri/OBsI8oMDuXZq92YUY1E/Dk/EG9E/B+XvcljK0WtLxVwLNa98vXe4QFt2ndcH9uMFtOWs7Wn
iTeAtmEgd0jWReANpM+GhVuvcgFdM5eTF5ZAGWzZFASXqc4OdDU4PGJ3PaQsW9a2evc086k/tgK5
i77HE1wnn4YQgD+GEkVeKbwVnE3uylUfv2URkJN3c+vfPRQi8gmBGqp4tvLMduCLJ4jo9k41R9HR
HYYipxat6UjdQOtC/HItIr1c0RoW822QM22GC7PURjmmL0xU53Vvza7ABM5VWocO5FGRN/E5G7dc
Oj6gps8sDcYdfZcD1EL3oHbMTrSKTed4dzka3K7MYC7U1mO0Y4aWGkkXyN7Cyrvj0m0aT1nQkq3E
LPZxqTyGYuSE2POLsL8pvJY5k6SC/BUMUv4AnWTd92HFo5KXDbcrmjV1jF6pmPLizlYTZIUphHYC
UlbNL67qPaoF3h1HIJ6ZXGURzoVqF1M5k0JE48hLIcnGj9gp4vWm8d3YLWwcGX1yitysrKGkep7Q
oilEurdFHbxGeKwe3BmRYOTSJ8bQoU7QwPOtuf5mqPu9hMRU37JMUpjmYvKX6n9tEhmnT1n++Vo4
r4m99ZKPClkJTXa+nhsqA0PTDMqtx7AYQQP3UBQ4be8VCCjujK8ZxHXHX3hYXy2rhxpax9zf5KMd
cAoSSUDf/aIsSOoW2cWMobIjBbv/jmrchW1viLbhdnCr9hBBOWP5tbxW37k5mgmMYalcglghW94x
9Q6I/XBZLgFPnHtmR7gjs304GIqjBc6NpQEDE6XQSHPIiagwMfdkSHPZJPxrbOdHx32ZCqP+6Yb7
mGWUUnQ7PHd2s8/epfA9ZqnGmjmJ/KZvT1GzMOOvzjlqULvzj7LcLeWwt7CcN/f1UiHVWu21Qlba
jxoI9tgCAsWtOsMJjzwb1OyHkCaaLNopuJEc7sgsqAknPQj6ArziibqroGD6RJ6mii+1P3ddie0l
SJouDGCz0jWSEeORVqoMobOh0RuRJML8hl7ElR1f6HHr2cBZo/3U+BTn6vuecYZ8i2uWN+XTP459
3CwD6SsTNpqgwHecTz8w8q4p96X1+UaV613QNWUIyhAXvVOxzv2EQVXB+Icz9hRWfeEyQZIiqIMp
ZD4pOnPgGGqbp+t6fqQkKZLic3/2qfoPsjLqO21P8djmuVMwdGr31HVTU2UjvFXMTMKdJUymmJUl
UwnL1BvNuyp3W+AdAKhA3SnuteeJTUQmziyZETfKvTo3CaXg/XlH/NkMDku+AcLEduwwC0oHq7TR
HWPWfJnEPn7C44y6J0KDts/ky0k2YcZnY/d88rz0eT3irPaNwN1RWM57P5gueKen3wdCqNsQt+ke
Z12ue3J5S0cFOtr132JJ7/RH4/qdNc9M4eg0xO5/EZtbkQ+Q8fgh4ubX7Rq0Dlfkalo3i1A3GkF+
zh13Ap18rgylzTtH4BT1ZNUBSy7qOLsVxEBjFv0Q0obMdu5zJX81c/Rz5J/6Kr1gSF3j7VQ3lQ2c
YpVsulFbRUQfkfl8taY0f8LqybhiT75t+t4fY9LtP+i+CZ8DXdgofZyoAlMi2VHghWX9UsghpzpY
IRuQ1sA9eaAlW0SNQ5/X6nhILFxUPHEgqFWgbBFKbIgDm71YDMapB0yWsZzrKw7eC4FPSnY2EE7i
DkyNwO/tneD1TsnFfgi9ZuEYs+5/bPObq7bTWz4wGF7Nf3pwvsjFU3gRwcO/TcGeAh2ljogPSdPB
iO+1GPnoS/QiPdnRALEpeLp7kxFGxL2WSukORraliNwvbzz3FttG3kbXJGQDi2EyxvNnl5kS/buD
ssJGdNU6eCDvwZ47Bu71ahd1oF6avgGRj3aFmIRlH44DamlpGy8izwaHw8U+Ci43mjYcEou28900
Y/XOZJN6qPr/Jm+mgmhffOVtcnEj4L7Kj/UOknO8kK56NukjZqhdMw+9KYDF05h7pRstR1vclzwk
Pz/8OZZLDCHKd0+Omi3ipeIIcYrCL5jdqSql2u1ac5SBuSKW+md//XoRXsO6EJxX4i2eVFRa7NT2
j2gnAIR++0NWSlkjCypZJJAFzer0z91kRkrjG08fEMX55uLNrw+jTRMXWeU/Z/M9P14KNd/ng4F8
OU8zPT6+GOHpKR9Ujmn5jsgJicDK15jHHUosD7FZZBr+NT7JrnjtNWBCxSN1U+fA78uA2Ral8fQc
wnF2tdb+JLFDY+2sDOo2rcfd/oNGYD4hgelQ5/JhfYi2SWywi3ebPzKQyKT/Q2JE7fWJ01fMO4IR
1+zgc6JZzlXFCdIMJgubIF8b9qOch5frFTTG7ueBL+RTFil9NmklBVu6JheJnydsMLIBAcVD4Q73
fajUt698v1t9cv56LuF2C60jDQ5itFZHjOSUya28MRmcerz3cHSGdar/HSgciJ1gFbYG6KRbWV4L
rYdA39xSpE14mWtR/6J6EdllHsPLnej7AgJSiLKnoZkNuEdAt+SXFO/BdoP/Ft/bYy2ED6xQP2rt
HjCEYZdVIluZJ+hWUgoZPbByVV6H68Kwm5E2XYaPpolncemzOl5jvq+QR3xE7dAwixim1XpB1q4S
FEctWBY9vubXC1nXPXMo8Wks/Hyoyo0gqTXiwX7qpG1/PeEzfnOZLPmOI9wYWTit5hrDkmwRYIrZ
zmk+xgD+1gg/YA91yi6eZ3LP71UJqK+W87ZxkOKxz/iYi14YqaobIo6IimkMv0He+sgbnMczXCIJ
p6PSkqjUqHSA23bcl/LMrY13XQlba12P7gk98EQPFmH2FTXrPobOL3HZaEqlQsEF8S06FBBU2QKF
cRk7I+8aTf6DJZ33k0YxEXCoq7he7PlLpZyAfQ858x5xRSLpBAMRLDNZCHED9L2POHQRNSX+u2Zt
50JzvBDV6HQf09FrpW7OprLdnHRH6TFE6+PjgYla318p+oNYWRGrZh5+XSnRxBO7eUXrxk3/Jddp
loc7vCBjPvsafO2O1S4ag9TawDmNn3uKqfvBUawnxC53aSgeP64sidl71UpYTP9CWshiSrpBffI4
xk8jIgAYuQ0LBRgMKU9SHxBWajd+MCIuLo4rotzPgadFzzFUkK+7uaROHBOtsBorfsgnHiRZ8SHl
KYYLQRqRegPiFAg1H6JNOBqx3KbeRU6v3wEhleAlKbR8N150NSxXYl1r3k8kfIxgIcb/HguhJCwf
h/U+8Z+irmYWK0g8RBT7DvcrWmm8DObEbD9kxswGyBvR+ABMXVl5Jc7tpvhZksQ10QRc3kEaI66R
qaqMjCqf8uAOavVol348p2tB9Kq0X7ZGKeb1IurW1p3x44GuTzm74lEgwDvQAQFGjqHMhAbhOmH4
jT4jD3KaK4V5udHl63ApI6biAqNanhKXPlD6W8sgoexUJMpZ1K6xvqMrZa3+6v+5anPinmChmmbn
5K+V1OOeZKElRhbQyFrlh1DQ68lDNepJJAk7ZOxvdboKx8CKtNr/jL2gX/giAjisWUCsRPe0myKR
OPlw5tBRXUoM82Xdy1gsuNCFY69nrW6fB641U03sSFt9yABA7GnmJ94p9bER2YKWs7bTKh3W2KW/
EeYxUuWb/RllbXvxHEUzzEdPPgmRBLZtU0pzkcA6KKGxn6FIx8sV+0adr0wJ20cBPBZ4cxTYN5n7
+79ot+tg+D8HDrkzRDPxFC5HZMcEhhuuU/SaSHyMoHHlqL3hU9rkh0+cz0JENdnGkSJEsUv0qGRq
sUoN/oRaWetSb/oVhvjM0H2Kx9rSA+5NJOCCWw3x2b2of+9iufoigYWGLpFJ68C0asn2j3rCBwTN
qb6NbjF/PPcv1zU/8W14ZbHCZtnqqtmGrVSbS4k6so65inFBo4YzJscKCtnp72eYOGirNpmt+bZg
kYB0aVX+8NkG2kGoyQKmPH4wJ7sCKeeCJQIrNrJR7B8Xk46Cv1UcyWFFV5TWp5nm5MguJmYHgbvp
VDlVshMZYqWUtJjaY+imRYfcc6lhzABpT0tiDpPC6OqA5TWc0vro7su93PlzJXIHPojg8oJV3Xw7
INrJX+SBkX9GrNvBwN2DwSQlWLNQO1Q78c7pz0OhnmVrz/OL/e+rJW9BA49opweKYiUMy2y9l/dE
uzlFUBZ7ye9iETFNEIL3r74uhQ3zntnqaccYBZe1Q0PE1veeLie+s9ieDmAfHJMpLiry1kA2/gbF
V2rXr2hr73adicKex3XskoKbvfrZ4mWNjG/vyGnocy+ETQQGBkF/O6oEmg/ha7Y7D8Rxbwq8Ki7/
8vCg5fnOSOCLupatDEYQb9Ql3tF04SCc99BDFHjNwuvrRziF/ziPiagCND3fxjw1VaJlj+cdyrgP
Y9SRfnvTodBY4UXfk4RacXu5czoKq3ylu3JuXyZ1KtRW0gmNr7fc2NBPHYIDz1d0BElLlPByGZ/p
MvQ01dmiDPLE2iCqJHWFdl7W1FcEiP0ovn0nXn/U174F4lmgpW3Um2RLNiAjQxg+ZkiriB/4074d
UIZoOEjbSzqwbkB55vbvAmTllzhASAQ8hVBqjbCcrFFV1+AaVtExBts4gwy4M24MXn5O1icjjyO+
Okzc3y1H7NyZU2/1ZrA9h2MsVWvE5I87LR4xWr6c9P831T0v/aOyKzZfl2JQXhd2ZXIOHbtmDl/C
1Ha0JtxYkSabmi5DI6U/hk8iREtk2OdIun3zEJRRSqNGJ61wIeWxjSCfi+l+groseSVm9hX3FDf2
DQ+CaKyTBtzwsIPQaeSujqgDsQtCBZoqT+d9kizSqX87Wd8wjcSpVqdvbe82oQ9kn/VhpBQ9xXm3
4CQMLgzXFhLVe7EiXzthZBUqrJU6U7Ws46km+FGY8Yj60IbqNlxOgM+4TJxpqNB4JUficINSDIxE
hUzc1wKXtuIEW59A7R6BPPif/y7MWEuhToxBLEk8O4nu6R3ZPD3HYLdmsbB5olat3LKIJY1hspoa
3AL/Wf81wuHhrKL41Ul4bjOBM3lxoMgvmQa/I84La9UtRb48tXVYIZHCsiDgWTnwkMtQjkGlFDhk
ck7kRTD4OEeixnLs/zLB9Si9CKOqLssE9FCfL941HJvGyMJJz9lLCrrrfMKfvb7FXJOXfe4kT9Kd
sdrJBd4LZ/onFk9tttQLqElFcp2ocrkz4T18TezBf7d3PHUmd9LgSTLpfxXhRwnmJusyOvlQIxga
vu59rFLKDKGVfxaoRqz26BmNob9dXMbB/1vLKqGMRqA7WS6Rz5YLllAkI2OWgKtUHWg0aBXcTqpf
gmzNrq561LHthMV6OT2bgTDYX7Cyht3VVs0azjsiwCNxlI/+d70kU+3biiAu7jbzJOeYXMSUUOzN
q1lKMh0xHQQ/lFf9LeZhW6mvNpvbBdZLhCklHvy0nB0kzQBnq+JpAUa3TDZI02iqE9866gi+Unin
Y2gs5wFBnAuXbSU4ccV9mQuLlNGg9hLlW8l1KnvvO8DAPIamnGzUpjgaVLVN6dSVlLsnrITzbWcZ
9+Yp1R2ggJHUR9z3tl8o4+xw9y8ebFNOqnRtmaCV3DCf5f9fcbg+ebhdimcuJ3MfrCNa+X/sXORW
fRgkHx/r0ytAwVlkff/D1Kn8bsg4QvquQiKyN4vaER/SH+oDA0jiZTf5DSPpy2uG4QzjY2zxWdap
4Ptz8d3mj3J2NQOuvVRLz8MMgkhYfKaEISXIipRo0UpBnh51L/Lupp8tJ8uJR5I82Y5FTKMYIg9s
lKEooevcT3cW//tvK5eLr7wPO3gFnyTm8TtNLwN9xKe57SrgjfSfVqxWsAHms/iuwVrEmp4Agnnj
7JUFcTjjHfKv/nZqAOmCFq2GPuYlbU4GB1NtDu04zmBwqBZDYcBUKUnDYKFbXNUzH/uuioJHc2ga
Isx4Td/AcDcXazHSPch48ISJ5DCOEGVgNhnjXZBORdlp4ggjOehJdsvgGjON5FCGAhPxF9j9AUwq
qUX6xNqt+l9m6V05tYbH0ajoJHuC4BuClOfAJhb60sn1sy2fwwEIktB9hBQ6rJ1Xa31ggs4LfFmv
y6wzJ1K/lvudiCWO3N/KteFZaKcKZxH0vE8vEW4dUKwu3nVqmOaJz2SG4G5ylsqHwEZx1m25CQpJ
cygDJz7ru2sQKiQvO9jJIGmAva2Om1qdGTVtsehzZYx48jg3i91+fvS0nMMxnLAJNkuYUWOuZLdx
gATliCllhCU9RxYJQ34GD+SVKidoXV5T8QN0XBokcUNamWT425eaAuiTIbapJtcVqteSHDveAOjN
yty0NGyk3E0WlJrzT6/1k5RLbgqEyzxdCBesIPSpneLHeP4XQCiL4iCc8VWFxnatSJFqEH+3uXFI
BrXllvHWbTFfai8b6++FIOyBJmGMjfC4+QphPwjnGQ0Xt7nfCtPGugpWkyJ3V+4rJwhg+2X0MMYX
wo6J7bqm6EizbEgN/Po2mmSk6EQJZYaF5a8BVA6o7rjPeIq8gT/BtF7mrW7+apt2FBKSKuNFVkBh
7LlASHb9gBkCDVbSJ+gU4a/dOfMX1f4jeZ1W32gKhIGrQ3TB4gFO+XXcGZ83YLLxO0vfYSlIsNw2
od3wEI+A6LtDqTbTR3tdWqnhFNfCeuuNkbxeYeHzfzepB93U1fYiLOdubcF2s+D9lrDUi0t2Iz3s
Bht+Fuu0K4lqKmTy25kaNlcH709YyGsIHLHc9RJGn6PF9kXuTpvWghZYp8eTZK10FL6ns68fcKEu
wvVF+bEbwVcwmIYIWPSAv00UY2ZdGVa/5Dmdah9RKa035BFKrzN+gCjs5GaJNwUdIpLd6eakdXKD
vcalY82c57Qp61g8PVEBiiQFdFcrCjG2S56ZrnWqLlE/FCTcki02TEiQ2WZMM8ZWSi1MUw9JpJAx
5Xi02i5Tcpm3Lqmw9MurA5Vxyo0dSf77Zzske82CoxjoNSIz+qskB5SdElwp/Pqzt7MuSgDxsJI1
D1oywBn361j4ztrV+GI+Tzh+4owL6JKzkNR/3fgdKmJkLDZ0Vuv3YWh9eQzoX+UopAk7ZA+Qovvx
Lf4TrRPXKSF0KpPPMQwz0WmoBOLRarJIFStV8vZusEcNQaCtI4kaTkSGa99P5/O5nWJmweGRVHkO
xMVykmh5spqEsOOF7GaofIjY3RKEJDiS0HduMzwXdfzG60DLs8/QvW6EtYxgVJZujXiZESI+st96
l8Awf7N5VwVXIu4SnC6XuDbUcIc6G9FWgNW7svj7Wd/fhi5RW2SjLipQav/ECtIJNiE5OV02Cj1U
JHTiMtovhkCc5KhnxNAD3JDBsSngDRaLquyW6fHzNOYyKgAqwdcKsytaG8R5eLXK+5cJ5MYDARGc
jdOJNrI8wXNcsXyn8v1Y0CeDbsdcHSj584S3hBAXb8R//kkgQrLaR9WDy5fKq4bEds12RFO8Uvv1
0nCi52riAjcrnAiPuA9kVMdV9BeOoadMOjMCUYa2yoORx8y0SV+UzlnxEjWSxhuPy5nGSpi6SUIK
xFmdBT5F+qViBOuXyopBkSAmBwGdVVLUGsBfxBDrePYAM/M7w6rNZgOAJwwpnCzarU+b++HRIlB1
xw+j8LhZgL6plkoHSRvVUoT6rB+07QUMlAf6KIOES6d8G7pxl8U+S5UXJsGktRsm/86aJUgmg/ii
o3Er8LPnBsGKLhH0WfCtZ3tExXvzlcTJ92L6swBosK8NtrQKdLVjMEFh5JJ6BeF7uyZlof7DvSoS
CB689eqe7uxPNgdjDMZEedsewmM1Oz7aBnc2hhcy0WCbJkh8GIGNxCHd9G4dcQY8YpqvMzpeF/Yx
3xpCdeBxhpdcWF8K0YIOgR14ex4/+dCqrZ3HvxvISegWhlRLSmzCzY/YfsW9AqCdAZSHTaLAtlZ3
sG6KETnyilnX7bla5UjUsl09zoLn+GfC6TMHY8mGKU5m8gab7fGb9KuU0f1mwxkOGn3EP3dR2P4A
3JS4Agm9WMltGXOyrnYrLMS89xFCPB0Ngs+tWrmYJ6NNwnIrMmCuuqLdMDD+wtNLkzAq2lZLqtre
8aEdnJxsqekx3SzbRuLfJBOAUhnalIZbKmc8OuJt6bjX3lr/0AYsXnshEq3Sb3fN4RdtXTvlooea
tIYrPvq4XuGr5gmaLBUplyeAtEAhyqbEbSAWnZl7l80a+5keYyk+BJwuoZDY88bH+5sihb67OCJR
J8v5CAY7Rey3hsuH/hrW2AV4GSNI1ATexvv/UE303o6sE2Cbfp9TXbsqsllc2wgEP/t/B72oY5Oh
FWndRITkkCW/XSIis55Wlsp6qZHF33DIrcP9kbITZNI0pbtb7njEkoedUUlKBYhAWBKwlJHQ62qs
GtU6tdq/5/Xo0pSQqoSNGzX4eawIBGRLrmQzuk6l0yWT2eDyHlGf/h1kfTvUQzEx7DgE1ZV6jVg9
bGTdogHj598ZbsAtJ/cLxhuagzp0KiiqQJkLf9lQXhus/S9BECGsrgUwEcu8ZJ7cM045zeiTXfDb
Ff4dM7gYnlu4Wc5fbudZ0p/nVpV4ccYE+JKCZ9g/Vj34/S2MaCXz58OYSPM9Gxp5EGopD+MNXK/G
gXExhqCB1af8L+bJK/5DInaCOMGLu62wom52SiCyoPoTo3bGTeALEU1eXLHyFGQhIO5fOT8NAsYu
hS2MdVL9eFuFiJqRmt0EDT+m5chVYxS6QcqejaiP4ryE/1BLz+NZqcQeKcWaUyfL5re+O0lxzLGB
AkrMW1+PTtz1olrEkOHcYFmbOwWw3PX99oTzqMnakhP83o6TsfpK4nYx8JkgfJf/rgcXi4aNACRf
S49veQ+Qgx1UdDPgXh9pbeAC7Pc9rik8JfSVHQpNq9xh9NeBXmYmgx3+P3QdePub3NHl/f8Sj/Nv
7N5YuJXZsqp0XCbwFQ==
`protect end_protected
