-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "ModelSim", encrypt_agent_info = "10.4d"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
EG6BSpo6wAx2OTIiXAfUyEna23ZkZuxg/r72v0cxdnsNeHgYklNU9oX8UJl8xpcn
L/Mra82DPUUKA259OQFgzsfFOR6jz74YDvGRzMX78nPq1bloTQQ8wO6WaAr0WAYw
H9weTglO7n9bmTa65uXNwlk+xKLXdjCj6VoGSYPUmTM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13828)

`protect DATA_BLOCK
Ha1vZ3YB2hHfWzXJJPDARqmQHiqdvqDNRiGpRMPcHtUzpcyN901R5OKXZwk9Vjoe
u4YlnTuxkPm0j0z1nT7WrDf2Ka2wDk9vtKdn0qM1Pt+rgWoUEMVjyGbCQAZlu1ya
pBWytE/NrrbfpP+hOtQ/jya0mXTP3Kif830+NQdQs2mfM0vbNPUim4qh6N48AYaR
1u/xDaHfCMlSK0ZfXbvTc9oieX4F9wG0m4+8jF6SLaFk5VL+MUUVoG8QLKa4l4r2
sG2Xt4+sE2+O4DzptX9yJfxnUBXjxuGCqEm+PrR/T+znS85uJ5Pimi1TNAO4/9yV
oHB6yw2aLKgi2mJfJD4IQWdwubWkmrV6mmvHsxcG03DeVnyvkk3eHWDKjbmpU0C1
w+zOM9rhmSwyFzhUQ7SCum39qUX5u/SUKgpgo+Z4pl+LDtLjjWfpa1Ap0N9U/GZR
oqWjcXjvnZOQAPER9tTbg+U+1pRizOhJMbBNkRcAVfbSebfheFwmDonOsjtjnGKL
X+g57kDgPVNdPw5gzppG6PC9IwhWYVPVdnVGiR9D6TXSosW/Hp/qe2UmfKKCMCp0
0Es9KgBlab26m6sbCmA5c4nmaIMje4pcsyq1P2oZ/sHDw6awEhzUqkE8HXull0/q
PHWgZJHmFkLNf1a3Vsgtn7AgMtQeKCr6kDvB/16/xyFpwwpVMMHSCQqfB3k6SGWN
cXJdTGYTB5N1Vuvk4exGe66Eiv1laaOXcx7zpP+khAZ4Y0JgFoiYegj4AZ5ajn72
YNLuDjI+ZwtHBL6KJ+czxQReuSyMD5lboEnfTS6ysyOPyAVv0FKBuYsurdS1CmcB
9YjJxRbYWFgl3AqGARwnrwTnC2Fqjuy+If1ZsVV76HZcaB7qlZADjhe3i9wZEUyx
uENP5x3C33mq2rTYyeMAKlCKPYrr86lGX/H07ssl63F+GeI/nVY5a5cGOEuNHgDe
ZyLd/xqyS3sPR471b8AdLX5LvhGaVlbIze0N36S7lwdgxkl+Mx7dFsxyU54j22CZ
8Os3t9hzJvQ5rniMqkgkcPDmb7YntNnGdfJuLDrszafXoqFFAJx0fXrpYgl4hrD6
7V9wl1Z5GGDazwSzehlYzJd33/eq4mKDmU7OtX202qIuREfaHVEQyM1JRj8KMExg
dya6lTUZFtM1KIaH9J+HlBC72W9g3l4N7q6YOWMg4b1Cf/KktFNZmCemOAHyEII0
Le9t4hskJqs+9sSzsAFTTtRdS6TzHqwRZ4iLsNCGy0QO+qPZ2mP1hPHxlF2OMhSX
YwtzOlpGOiaJvB5iKc/7Tlv60HoT3N1bMlB/pIva0GWwQw1+00dR/QdIoJZFrj6l
LlFYq/ipvxT672mt0ITO5qTA3ULj9vOJNtKCDsEnBDDYxnE3BUFE7c5yGNIRefea
iBMIDwdboWd92rcIA+dNTXbXP1Bt/UrCsP7PFhcReq0Dp9Z2kog/XcrSQ2u18fVQ
bGZ9EGxkbu6BxDcmucbyslqK41/I3SUGJHVjwljakCi+sbJlK9cotsb5TtLgTaL6
PWpambtobx65SNiraOFj62Du5bOqx54wUQMRi0SrJ6EYY14u1rvDFk5GG0n2Nu0l
Jih09DtFWtQ+ZeHid4knSN8p2ez0RE/+DyXCtf7SLsNX3TvjOerEraDO8qW7eZuX
efXA9lco7y5v5HlFRAe47iUXk8sDXz6ND25lzo0jO86lDOz2V3rY2tBwaVDr//tf
fZ2/hY+pU/yA9c5LNj9KxFDbVBLzOOkNqeIxQ2+F9/7as/unz08slOghqEyySe5Y
cT+Q8qkMdPVjQQZTgvqhNU4RKW9V7rAnxWjLYtvNw2BG+QULLtY9rSOUaWFbrxRS
peQq+eoDG7oOpOg8KHdu9cuBNTKGlUaj1QHso/3dYf0io0WP4/XnJcv7r3iyd3Bq
SuZQG6QJ4f8CEm6YwiiXhSH5zU7jejKd3HvuYDY9fP/DlmMeUTArXr+LDkCKc78V
MSOnpZT36f9R5AJQuVf9zA9BOcdAnKSNZzgM8u80uUgus3uv5240jVM4bOAIRIHR
kJ4gKQIPlroIsgFcn9fInafeFq+RnIurJCAqrDz2ubO3LW0nLojlqeKzwNUX363L
u/6552dJiSR7Vy+V9gFsj8u/HQwaWfpugL1606OpDXZL08Hkvic7W4wwSKZTIKTb
5FkQ2osUNcoPhPMhZFkEQIb4n6pZNb3hhzJ60v60QcZp81/DelxTvZ4xUV5CgX3y
ml/Ti0tk+NWJY9QcbBw3Lkptj2QrBbeh//QCQzJVrir6ZIzbaLTi1kr6Gd5MTlmO
gMqqnYFth7D1tVJNaIfs5c02djmZ1gZCM0uJb+3knr32XYEhjbeNo6aGAFpShXTo
CUpKOSNfoZA1CeVjRBNtofFk0cHFtaPt5JWDSkmkkTr+RyGVEJiVM2bJmZyeoGfG
s+Cyxl6Kh9D3LWiIarAEuwtlfZhiLx8oX5xVUFwsAnV/pci68DdC/+c2rYDqmRdF
Zat8llAwEikS5LYfqkHR3PnCu/n3oiR1H+64yl1EN22/S11l1gN8+YlM1RnBvt74
NEOzlEVzr8/pdd+aBiXYrIZ0/Vq1Qidq/81fBbFEfFYqj7JjCzmff05ifkwxkMfI
U6Vk0FeUGE6TSKINiIJo3JFY1cYt24HyxqLKahUtk8USpBGItG6Sc419twiZlq/f
Zz5r/K4Kx/Qj4VmMs57VKt3ctTF91mGrF3VUTbQqjKu/7B7PmtIX3CtQnVCfLapq
xxTjx4p/BltJ2uhDVjX/qCvuH31ZvvIc1g8FKXiHLnY2Tak/IUBBlHLc2V9L5pom
hCKbhvu3HrlncUEjBSvbzfzxKB3RH81S9KzJnNxdoVHECr1oCz7W87IoCNH3fQ3Q
PRWjd/1RD0Hc3+CB+lZ1kFvRVV0TmrowOB7Z/HOWIdshGSWuvf8bvsHAslp+yFBV
ECMTkj+i5Cb0d/9vqACHDqyl0acP/S1okjM50D8a/AMSFXjrJDZNWHV3f4NRX0AQ
od0ymScD7LL4hLoUOL6xXUI20mEND+M964ixJ1Ec7pssUB2gkzMUqf9RHOt0eUs9
7arV0iHZNvdVkSt7i2AQvx9arS0CQV/bX22z+BKZjapHC6rWCCKkzyLl6ud2AVv6
GfigOfUtKfSpcI52E0ac3aOitrRUU2XdoKkq3CUBJfGi3lzwgWd9NitWy+4XWm/t
YGEPjCP4xAoRHO2WiX+XQXPa526cXt1AKnESUjRktAbB7Y9jI2DhXL5h6oy/+DE3
hEYr+z35WiWGXIDmkDoPckHDVbU1uElZ/P8DBa0ttGdgInTro+QEHuwO3TfX3Ey/
+fXFt7xDS+q1mNojKrErSFGeasbI6wc4Om969l6jJrtD7n0JySln3PFXh6MwZC9X
/SqQJpvzP/Goc3uGtMPS1U5al58jeglytwjg2Jp9mkZDvc0imKbILG3kODYF0jZI
bXHnBD2Z0OWCbICSUlMwhaVn3R0EN+01z/vmEg4tQiecfHoCTec+2+x5VWPOBRM+
okTNogpClOOvVTVni0HTd3N8XIGc+kgpW0VKY3t/LbiJwHZbsWwwFR8xQ0eJSEo8
ymw9ceK5aGQqg0Kl+vGjqTp4NYaGIkvBrYkIFoZV2LfyCfmbYR28zzrMSumKnMj+
ikH8SQZRK++rEyq4QEPZXuC/qvFmaoTnZdNZUtKObqUPf1x988BZDYFkTtwBpP6s
/NMdwAx32KM+18+nWbGcl3XDuzjAm7wWR3FhpbOcu9YiuFbvgd2+0FE1qZ7+WQ7B
frVkG/euwTF6EOz7Pfl3KcIEH/qEWSUplOI9IvOR3FQS4IJh0b/qtMb2GB8DFlRk
Flod18wug8c4+3tXkbaBaY7TD7zvpS7xRwMUS7lpI/gLM9U5WhvILLCNF3kHMofz
z2U1urdOb7ej0LZ/UhNv0RzHOWY8SZ3Z4TKtJyJJ3DiTpBS3zZJFLLzX6gwvsdRO
ilEMKpxvIF/P8aJacEINH8DS5qDzxq29uplnC8dUhhWts+Gqldzd7RW/BUNc78ol
DQXCKtCVb2FItXQNHSFCqMJ+Pq7foOTIRt9dwbVXxhJLI1QsMQngXJHGsxoUoAYC
SvblF60sUAx9jH/Gj1otfd4/05ZdeMMg0Gu4Bcn3c7y35H7DCPdTMb3P7lHWKtSB
bQ/qACGcKZn809aKSDN5nPWu+gOezmf09A+j3EYZ9u3HBEGCZkDoUGdxjqcPlWzP
JGuVwOvBGI1uD9HtUlGnAqT7EcKGdjEyRGF3Wzl+FoEI7DYgVkfhudswa6O0BGNJ
y39XUe58yL47NhDcm8heiTJk1uBXOrhHk7O88wGlmxO17Bu9ANUAPxXHvaaYuR3I
oP/hNHZ3x4mthHaPCFDoh9FwqY/2tBzHcWJak2ZbfxTw2R+UTr93eoKIhJoj6mmn
t/RjfNFqEiYxWCojOzEPF7XJGfl5U23Bb3con1RgnK9R8CjIZdZjZBcMq/yj3F7N
jpd5sifiHnYES+kR1poOogm7/6tF4BIC/OUGhcgZL+SoURkLTJRxyaetUOqetenu
F8/GUs4mreKw1BSjp6GdQoXDhYl4QXhg+3t0a3WIoAX8HpT/BbXEHzbJQ+8EzpDa
c7u2GMb0xl41rhzoz6INUpGq1RlXatMWeJ0K/fbFmbmlTufrs7GqtIeRh6c6Mf8I
gf2/2QTDefNzb4bGMBaQ9uI3hJrj95EUKQi1DYxBZcLMfyTqATJeR3Znvh+b7N0E
0fXUrh1VDv/aHvjhvvj5xeJ2/ga9b/Sviahw6QRxBcg7nx7b+v5FMTrevMmC9Rhm
XUAbPQ1qT4XnpHEaj6W4HM4MYfUjcIya3TSlCGWrkXHPxTP4scV+r9OHL44l54SU
HBkv5iXXQr4yr4i8OW4Nwh0mYTTxfFLsW9ME+TiKtqwPtahxIwQhLJEZpnUiWyqk
pNaJXOGQ1Q3XX2JMvzsqlB60VxXYyqNhKi+14MZAgF1E2OOboUrrc8hbYSwwz4tE
S2AaHk+T2qrtStWWayrcimhGXvR+6CpgIhvyHQtjn26bbSflmk4SPfB82VQWkC0o
6UEtpAogEZicFjR80AwBv1F3olz/QOK85n5CbDE9ID+ocTz6DXnKFLXc/IB8z+8d
Qqt4FXVQ/lIM0b+N1gqAy2DN8fA5rtSbPPxPjoyZUEnkOQtt1Sw4jCBLiJV5YsEZ
tImZ+KLEKrjpjqAv+X3QcGiShTQoezOotpOPNjcDgFAASnNB+HqhoQs8DIGwEOB2
juEwpz7JqegbAzVtQKLuXwOBYHZis7rTnt5Hu0A18nO0kOfyqMeamzvNW+B1A9pL
DmI/4k1Z5pO3+27RrYcU7UgLAcvggUKA8Mc8yXrafNerTU9nBtBTJtQIYwrFXmYq
03XUYBwNS5UpZp642HOQW+BfJQJByn/zjMMK6bCIJatkB6ptq4DwejDW6D08I7FJ
vzk634D7xgy4F2ORN7f6GjpJmsLe7CJaIrTT3Yr9fEVm5pNiTSQnjkCAYsF/iwPV
ltC+ZHLjtM9CS/8N/CGJJ8y0NhrJgs4IpuWAgzmDfBdxaJqyaz4PHb4zlkFG7LCv
TLRtwyVnO8ukNHWFYV5uXVHSIxu0enCij7pGQgv2UGMreEs4y691BegXAPCwiOxb
I9JJGQAcBIkhtUSQdS65s7bEmf40qgX52MgP/hx3O0Qs4a5hPhLKo6i5y0ATG4EG
SL1NCNOjKLClVuGKFQnM+0ak6hXcZlPbK5pkxtA1CrMKcP6MU2qg5GnTex8E3KF4
jlIoUSPkdPThoPCmYacEoxp5afTqC1AdxEG5HCs/6gZuShnBHilx6Zsqn5P3bZ2k
xlZ+EwVnA9C6gtysijGu2N7XLLntFfXQcTuJ5jMA+Me5BGPcrbHU1ZDtzS2uke32
3q4hLcuvVqylU66KwJH4zy6Ic+qtKk4SsTTaogobQpSjA/gFbYeiIZ6nRIBpSDJC
U89oDyfYQ9nVmg8ub/sXE8LI+4JTaQPX1BLC2HxMiAbz3vSq7kcPdkFp+vpZ5czW
Tcmc7NNlzAg9YAXzXYQtd+HNqY2I9pUoEgFIjurjIH1+jbvIB8h/YJKtiJfut/5f
Ww+HZZ8bV8MVFNj9YoDtZlsFqxw9YWQo07hbHEgle9j/na1VsPlqbUmtjH/OFPpx
nEQ8lGvy/f7PfhNaTXwF7UeBJ1Eu3l6V0X7YOi36bYiLtWX8EV2GkUJxZFrbYjW8
q4gyoJGWiH1DFVEcbWFjDp00LfuNbt/Bnc3Zum2j5KRKWa5hBBeGYFQ6Isq5ZNKJ
7o7M/ZYmXcrDdgU88FTP4fGi4vsWHHTq2F7xnPWS9pijVctE7I3qxZeulXk3p+GC
wAcwajiVgFefa5fmMFYyFBSs72c3JrZ4eblJnzkKlLUw7Ly4rK7pO0VoMlb05A38
zXWHqbaJ5H9GW7SjQFGMy7SoQZQuIzELuAevGFDcMJW1Q6/V6KNyKNFLC5e/eKsP
tPb4wDd/4a968YS4WXXK8Yopc/h5Zit3cEeM+zCa5ajCT3am/S8Zz8yQArMMMzC9
y7aJTi7XDKnbCPKUpgPHqxKjGiu3sEGjthEYYZi7kHGsNCzhScOLSsx8cilCbYPA
RtbTD+U1AaD4aNUTxqIhoqv3hCYL8Dz0u3m91uanCLIV1axrhTmIAFeHexB3TYhp
gOtPrUuLvv4UINaRvbx1brwZyg7Vb4qeRX5ccHbN1tR80YdMtAmq88JLOkHQQ5FX
pOpoLfriYcWq2qJ9G01UA4YakP9F4MGxfxt8jkfbjRmWJ4Bk0BJ5FKP36xmnluni
o/EM2ecqNH3qygfLEoJjaX+dzAE40JmZNDCXnLaR1ZTTe3fdZ7LH5EiqW4B3CPjc
oM8HGT0kBhjzPWytL7jdF4eaOI5U3ARoFrMRrQ7mqz30MiS/FPmKa7OZ7UtVulGL
GOC4BXyGxA57Ef8h13Ty3hwRScha6uHffM9TfX6wwOrTKTQdbbaCuksTIhjujFRl
J6xjFi2i6jS2LjplOnKGU5setsPUfr36jLj/3ZQHq5O/8V8csmgwoccf/zXvxrXk
0M6OE1DCmWzRizVaV9dVduucCwXeSUM0aWPhZ5P0FbbVDv/jiW+Su69DZhXQloNj
JxRr8gz6CxnhMgX2ZDwm7dOsQoY321bitlGTG5/9infXbGIoNSxN741rXHMl6mJ8
YmFA+hgUWN39Pz7BPlQxsLLIopkeFe+x97Zid8GtQtBajrSmxa/KJM+wbLx3TXzQ
ugbzDv7bwmnA/6okUf5fdWymXGR1YmiprVDjB72Y4Sx1xL2a1uAUjodz+AtdphcB
Wy8ICy/t+BCAVcjDVvJeqLQj6XyxOrjFU8Glj4VgZEjvwv5NfgwA4cCZgQldSQzT
MtYszV2b9Zeih9uDiVyNaMt7T+cEnxESwGnOpSO6QSsgQCpCRaMP5iGl2WYlkiHO
VqiYqSw9AeD3UJZVWuB+TPN3HqU1SDVV7Wej+4rQ19YMn14jSwhK/TK+xMNWQdBG
xpSSuAGLDr3g0dJ2SX8uw7RM3RSfPTXjgq+gFC1Hmr2tvZNf9Mn6ktx5gcauyY37
CdyGX6jPtZ3BHDd3/zDjgAej9kLowVxo/6QCYvFen5bMcTChnlTY5BsDBLk66dZp
bv99/UzFaZ9iH2yvH9dAyE+bAPH+FRHixT/l6QDr/VEK3LvpGCQwEr3Ss+PI1cZ8
OFWT+0JrH+RXtWmTNSgV6lsfTvi2/NEYUxgdRPlKcjkxX7wUmtui/WTJ3OSydTsX
YUT3TuCpmN/M7oSM7g46leN6v/O+m4SlPACZ9kOJAyNgmqAejYhZaS6o+mecOlE2
RURLVWK1+CuGfewbveIsuEYPm4YPKs1XhUreDM2XLPD/8A3JzkiHX3Ws94N+m8Ip
X/eTBzqdA2ooxKR/rabGGF1fDcVOboRvPVuzVKHIbbVBJNmUxQXvLEqF8h922WZs
ESttcLY2OYwl61RybwtZOpsVIxMXH1cPRt53VrOSCM42iLagOq7vHFwEjiaY5tSj
i9K+yyJ/6/fRo6F1w4IG5F7ZxS7S2rDUfQ5lPGPP0T0lyzyzkVl0lEFgcmoCWGbJ
hFdQVPWnH24RpiG8d5oM1Vu7IjDLFQbSQnMRo2p2XrIkpREaoZGcuQ/Rd5rNMAlf
5wM31KYglW8l7itkL8jdkeF1KIVcxRyI3reQ2PIL/BaVYOSlzd8mfZ+m/FDWoMZm
5iRfDBGho0J7RRKoNL1KiKkFM6C5F4fNKcLEocKO7hz6lNYOjUiaoyX0sTl3cYx5
k2PTvm7ue4gPD2S9qQgVrl85hJvuW4zGP1fK4J8n7tAUIVwHqfw9S8AJ6fpIbfXf
7ymq2zfpQHM0Awce7Nbqms4i6Y3TKHmX6rijQCzIjLe3rB+s2G0RrGNe6jw6M9Xl
QZpGGIEJ1F6WqwI6ixVwaFuiPYfwppn27pyOR03Xf0TQvGksTxSi9Sf0e2skmFYE
+7qTfb7QmnXwbufW1XAqcKR+Cm1uoqxtvo1zt9RJa8deQcs4mb9c5RK+M4SdnG5f
Hq2DCmkJhAmZrHOxD1jQ+q9lE8ybUk6f1kwSh5ctvG16kPXEr12ZR3jDg86d3tUz
NRXJIKYNs8ufx+vDY0zX1natuXxaI7agi/ptg8cg1Kcwcf9tajGpuxzSdt+ZLXMA
GkiRzyoLd69uzkNWM+VN7rlfMIAhc4HioXjDsnxzktgHTCGYO55HOetiCyA3Jorx
UAhKCJekaaBaGvN34wr++T8S7jWWEN6ot3pHCaURCgTvN1/UWGaPIUofG+Y3E/tT
/iLqj3N1KjlhkF6JMzzQRYh6wTDj5thhHe8B+R+YQjZluepzzPItw9djDQD2dCeW
8m0mKoP98eeC4FLs8EXUr3PEOae8fegOvLDsARCKWY0w3dNw3f7Yj9Vp1RBXEz/i
DCI3Dus/rx2IYWZc00PqPNUxHNSx0V1zX3sX9naKh3l1NOW2kHhjrB/MHj9fJG58
ak9Qnkcno4ZxzLnD3/+TWqYTRNdaVe44+e08j5Kh835bevzkA6XsNMv/chp7kVM4
sJg+uPrLYzq5BCvYqRk9wj76GJej+MHtMfSNXV7BAPP+rGEYCvvrcgIS+kUP4CLz
B4GaBh0baee1Q4l2jTFbh4eTlcAzxZa6pV4RrgxHH1vtcNmE9vPxzKWoZ7w57h0p
Y1db0LpdR3bVKPltyQA9Uh8asTkGcSKkjXHBF1B3SuJ3papqfcFbusoYfIgeWOtF
CS+Yq7RboJMfhM7v/L+WlCbU01HpeOFeO1J32nmL/uam12m9Mn+YnuaG1S5J5IgL
Hd27g8nWs9e2/HF1Zw0SwF5P5f/wV9AChfeeqfIg2nNRr083RkLi1Ivk6WeZuwWb
tpUqCZ8U8XTSZpLb7Jpmn7eRlpM+itbRV5tbPYg3akWjwttXnbFeGrBVWdAQyBYL
prFCMKG4SE/TEN+1hSo4w8g2zsXiIYpVzPf1QjWkf2S1lj/HLzITm3pc85GujYra
uaTgh6V6fNqw8rR4xdLD+Uu7AaBYqX3vjy2JT/s8UOeAitOxIwdSPeCcKB99mjD4
1xFvLQPUi9/uY02sPOqTGfDo042tTMYN1qWvCCW2b4r6mGzqLY6RbwOTYiFzKy9X
55RRWwHFqjX0dsv5Nt9uCsEuNOxkl3a1GIIl6vXlQb+KvvBYNggrLNIwVb507Ar9
yOBoCql3CXuBNCorgLNi4h/x1fYJDFf7o342eU1xPIDEI7debbZoqwIG5Wp+/DD7
Yyt4ALoEaDVbS6tok47x5xSK7mi9fKWuTvtal6tDS0GvpdVv3xKiz3eB63+k6S9P
jOjFsxHLzO6FDGPFdMKyaO0pptjUqD2/cDtzCaEvbWiqKKm+XBqhf1s/d+s4l8/e
8wHu+hpnrUAhuZKCZHHfhmZPtP/BWd2tEnU0VUj6EbBjAksifGH/i8coWXNtvniM
J7a747NADD30aoka7Amq7i9nSB2AeyIFkRVvxSWWb7+L5cPugPBSF5sR9wC5BRdH
UPJpi6bNAm87SiqggwwaTL3Pwda7itBdh6iLqVQeyTpw8pWUThWdZ4V1SBEYPWFy
uDvKoJt6+Li/jKTdHzalhlA+hvTncB2xR+Bv+/OHeFkChJhH112pwLJl8hh3qVXj
TYJ+QJtoZLI+3+bToz4c6RRjHTCh5bvvA63m+NQ8cDDrTaZugKyFLZpNwJXOVJUL
75Cc2wk3fXvGQbY2Nd1/kMHSp5lPoezAKlbP13tIV1b61ggbMDhqU9HBPJeQZH+8
7pn+uUPosLBqHdDeBpid3oIf9YIbMFhGpxbcL9noAIP2N8iL3KEm5ETekjj/Ouil
b1W5Zsg8sBNFSZ8wfHXyj2tn05rbqG3J/ZKhS8mPUGiUOEaU/+SL9i5p1zwqLOFZ
CYFwI5joDTFsK65ZCcDeiajp62moKnflNQWplYPbnSQXrAeMCYoZavXyevTEccYi
aDs9CqIk08ikzaMStZHIgDKFIGVEjXCVZr4nZMDIdKh1j3a1FibJFDvQ3+9yrF30
pF+v+3ez3IuxQF2jMXXEeM0FGGlTOhHokupdiRJ6GDPGRRfJISDlgB/RaQjh9lx/
TApijRvDHdYmMALacgjkQ95PpwtZzN8HURsJotjrUzVJArKSL26msItV9Dt2YepX
kDNSYY/n0YAHsIQeQY5LLogQlVKNPL5mI6jhflqXPNcctyqLu73Oelpsh4hkB03g
b3lSFf8cyxs0rUWr3lEPXXwrUooBwIUrtzfnjU5zqq+OdV7DM+tIhiRgJ6oqQdXB
DcGWx4sN5vHtz11bIOozQaouR1eVRT+NGNI789OHbfVh1RVtYeT4B4fmiWaICQE2
BgKaKC/W3lFOrboDMhtTzJsfD/6C2nTUp7h8LGayNxN4VfbGaHq6pd2V/r2n9sgr
XQDS7sCEQYxYlRRWIAoo7sSBRnJvD4m7Av+JjQuq81c69HKtj96TOT3H8puJIw9y
ANBi8EvOVEtUk6geaMQsrwuKryrInBPwaT6be2aAmKWocDfOLfLhV1d2EhGY4V+i
yqWQBN0AclFg2CXLr5XI1tsyfO8+KTI02XpHt4xpOokVsHcrFWusHNRWj/FNW0Qw
SkaxtsqHXcWkTNRKsWaBripbTXjllRuCSAPOKyLwh7uHkBQWMrZrKz+Llj6tmPXl
YTgYjH7IiEH6MLEmTygtIqIKjXVCQJnqGrTwm0syJMPrJ6maX//v/4lS1+3EJyR7
njeoXHpiGSXMbKDC79oRn3SmhrxEOnfK8F8Vzow8rT0uBaYkqkjlpHcP6iYo2YQs
TdWyMnONv2dl2Mf0SNwQ0JqVFF5HiHCgnhDqPiQSv32S1ohDt8sN37Kmc+Jm4h/n
3OmrRfS0ecVlC0+WJxt5049hs2nYbClsWOfTi7FGiBG7IWQ/zG/bVf4cqMYttuII
fEhPC+UCh19wGBYdwF3I8cdOSQRSzNpf1R5W9YFPiaj3V5yKj5bPii1Yo/2GpugK
RGbumyGp+MY2AKZBeoTBhka7WMVQWaiT+vs22qT6sOiLuLnpMgbN4EmlRWwlkRCs
acWrfTYl9XEy3ceNgUI2QN6rdgsj+grihSCcQm+Axbq68ee+kUFxuWSa8x4hdv4H
BtiUFoyTyP9r70EFE0ra9o4kwZxoY7z0m0B5PNThzUDneRVZjW5AZm8sLfxPBpuy
lXvj3Mf1f/hqjyqxz9ybwt8i41d6zB41n8JWpDvDq0wJdeD9BPKktmtTkGWJBc06
yDcsInPh2NXCe8z7AHzuHKP9E0HFb1A/kMr1+baDCJwbo4wK7zHyxsE8Uikqjfma
wfQ2qhhPdA0u85SKhXhinXVdkdPMmMbsXUMmy5xDU9/hofGNlmDlrRJytZebACfx
Idcx3hXqYqdtesZETXyfs4qqp4OcyDdluvrMdBVkn8t0wmRDNk/xE3yClgRLEkhQ
vOj8WiWC4F7L8eyrWCvgTKPTbDYUPjIiiXd7iesK3ICpgLmsSgI1ibOOdMNa5wZo
ksxSMSMC6mPpngG9XLoziTLOjzQfSuBet6MBgXIr8qWevyO5zkV8KKxYYLF5pQIH
DBImV43fcYlyIfk8IXA3NxhivarTuVmg+0cMpjD7D8PxuoWYeT9/IQjrTE8UAcfz
hUtEasEJy8lrQNde3c4SFuah1UI+h5wtvkTswyD9WR4ylaGMGFNaj6mhLhfgGAxY
5eN++MCDjVGwGjDuAkxcwv22sFhylRObVPUSH/9ZF2iVw62/QW3gVaKkSmP15GFH
RpyL3XZUIUHYrA3Z18Jnksy6bpNBgrzaJPWp5ZxMixXAMWxC2j75Okeqds/C+WVp
c0ZuMPHebnaxLnMpKpfmFL+Gjql+t+/JcoBXna8HYIY3XDkFGeRmPoY+9x2bLTtL
n4OyzQTBlAehyw4qPcBc+TgC9DOq9FkhAGtDH7fDcxIXxA9H7mnW7ulzqMvAUjhA
q8YRN0IcMWkebvA0tEtbWT/DDbjMS7oVRdtoLwoLxWtR5umB+iQW/AaeckkxuwMs
4XOdp9dWCaX0ofPMowJfvJDrUcZlXGZt3R0baP0v0FPPbjIZksqFBXmn55cyN1sG
uCkzf0eaBxEVodV2HRyTOJt/qGBOfTTnbWCSJL0wDXNV4uBpUugLs/wnAeNs+q9G
zB6rXkTTqxS1P24CEbnObmYGb1pIj7NPFNE2dpFrNdPLMqAlzu3GjuJy4BfZUBgE
ObNtMmSIJuRGqc6eCIFoWeDoZBWd2MaxRhb7mYtI1Uw2TGNPvsaC6qj3n5wht90r
YSsPOnLfOW3h8eHONQ4Qxhnbwfpo7fT2HiweSfeukHxEU28wVTQGWOfvN1hY/20x
gACUNTZUSz1TKnpE8To1xgLl3Td59Mte1DvXNlCN1QVPKcTGv5gRcgeK6c2mbiFK
xOAZNM1gYTBt2r18/UNYXuO5L8VVhQNLD7Q2jybaureZ+L1jaPWtwjs43EvXRtq7
aMrsb+WqQepTemB3NUrS0ZSuXdFRJG8aLxeumOoh0tSXSWewJm4dPEWJlEwZ7a4N
5tKKdjPiJOZHwfZpIvF2KPBMixhCfxOxCgArKS2iyRsKVEPNADFwrAwq8LRj7jdo
J3s94DPbKdFJVX2dm5Yhe/aV4pRR+v2dGZvq36MripVF5FX5nsLDMBafprsyFzyY
SkVpZ+jnW0g/z7xrey1GfzRZYTTWP6tlnuqm6ozoKTi/OBl0BPMm0m8Isy/X5W2U
YeqTMrjP+MpjHzgdsxhS3iBsRr3TtFd/sgtC8/ceyBUawyKm/Fgroj1yXVxvQJCu
Cm+wpkqgirymW+PukbnSvCDccCBxfaPTNeQGKXQjx0LAlCogByei8EyM2iTGjGzb
sUu70o31289L2CnCM8P6mVWUobMMmDjJ7LGDPHNVfA3r4rWP2i+sKhmXiSLoFsg+
qwkM4YOaTfV7BmZ/OCZkUk8bOSKXgamfs0viMp8vN85t3IKaSq3lzzJAdJEw4/29
hnI4xH4+bOHP9mdgnlVVDpJBrMsWdUpzt7hRKeN4riw1p8rvgB14iOzXCWMqesNH
GOqWNQO50bnmlYAwSrMbh+3h8cDAel5me5sdhzymswnARQSe4Mf6h2EYO0MqM2rI
2TNwYV5zXtX45x289ybIWClbWoMYy1gi5tZxbV7ZrIdT4/yDuYgnx+kozde71kjP
2Fh4eEhrydZRlsoRjBWzLyHUsHnsmCr09VsvVlczyA0cFnhjfF+y1N3fO9XZutb3
vFs7xUhGMqMw0tuvBt7SGpa985NYB80WmRn68sX4Cwxq16O09adf2SqwEMnul7Qr
RRbdyIr88gm3TO0OHsVQpuqu1QSFTvT/v1GN6jF8ir6G4LtgEGBSOxscKK0khjLY
fG4pGmYpnrQSwOYV531YnsWfyW0Kvs4KhFnLaMKqjPPA/3UUVO5hRQlrjBLM+tlZ
2J2x2TymEtB9mMcBFxRRUdC6qjVqEeHDoqKNwml21DB5RLEOkSQEUDhz4ymEILQj
TiklBhV4p2Wt7lCHzHwLH0uGjoMWiKrAKb/1ZsgRS4VjFhZuyqxuy/BY0K1qkdww
BKibwLcurF+L5+a9R/WPa57PzlUhT4yO3cZ2BVGMni+cIGOU5zR3LJ8otU238DTp
dIVBlf66GUPET9/8zUQSbK48jKQFTgv/aa4XlofE4j4/qzbngA02rJkI0s34nk+Y
bIEhe1IE+K9T4gXkx4vbhrFk0seNE5XTF1gZ6rGAqhIFdh+wjinb8LLoL2zOutJ9
Mga0AvRNwjlADNfQWsah3v0+G6NfOrL0dKysgyMDQpg8sf1CWktAp5jqSbdlZGyN
OZtkf1LbYe2wAi/rEXbmWQcEDYXR7eCLEFi9cnDu4vlzPEXADBpcoYkRpLH/q2tX
m3XkmLb4IZENzHlzzSfAbd/3f/zSrrXcY4wQydf6q2SZloXOmU6U5+A7VmnqdDF/
qF/b8km/knCKqvAPiS2sPkRuiGnm2XP7mBuTb5pH0z0cllVxRVZSjumXaA6BbRPt
Qm6idw8FTergoGarFHP6leOIt0mzt/1xInmCSzAuKmrmWbJ0/tJKqCUgw8mO0eNx
tbIfiulHkkx0ffhm0/RaHOZTX1KPJKHrNAHhmVIane1YObAd+KUI7/jlva6mgTzE
aWI5jOQD0bTf2TD2yshhhulGmyhqHNKAli7chQxLe2h1yC37rhjNJBnqRnIcC77b
XOA7qBOilqDbNq2VXc3RJGVeBbSUQ68FlYwAUOPr2swkp2tbhxuT9zG3VPs+UJP1
RLNbbWSkZo7J9lrSi9nWLOKnWHwY7GZ0hcfUe16Nu+CxE8t9WmZNLjTNtEVKjRjQ
S46XPR21qhNQszO2nx2SxlA1kiMwTPqHCmgv1K2sgsjngIxx67ow33fpvnSzkqrn
i0vDPPz4j9KSTX7qrjmF18jkN9k6dEU6fUvlmNXgB2AqWttktSg6Jv1m17kqVk+f
NNkVzYBCKBfD0e20rxDntaVQ/0IGM2x21PtOwmChKqqdVuvcVMkiZgKYux8flgmI
xoG9VfDQvTyj0Z/uluyX/N06FW65M1DAO4YJoW/fcPZ1FxIR479O/yL2ecU5xB/8
whjJfL7nN5K6VUOm022o+SN6UunFDlayYpTXNt8uEctBm47S99dGAvnfVqJThD+R
AX/BRKQ62rD2puoOG9JMbGJ3P+k4N0ceX8GP+uMLiOKmFCnkDG8a4lZ5ik1qI6r9
rOZYfjXTbGTC+OWWrg01vlMbSlNiN6M2GTpNq5/yINkKJ32YEGCpPJCAQnkTEkDl
BMLXsSh6FXMlwevFNiqTl+0d7xBozUiykn3koZejaakZhcAqSGYKy6MSUkW7HfbQ
OvmXr+87FWYrpC3XlVLKK0+JsEKmDHZQT/g4Az3Rof7bD71Lixh90cFyXn4y1LdC
a5BeI4TUMXTKUW/7csFol2W+xQ39a0Q54O9PHDeWejJ/ousaKygvnfOgQSnVDuaC
6zYsimZjhX8HqXSSGpF0iefkixDf3oVDYidHWcq+BC9rPS9SPs5+79tg8FxkK1fj
sHrWW0lmEFwI7+1/L6HsGmHQL2ElsZmDYiEOMhAxmgej7mD1LpV7tGFpLsmC/nG7
rdR66MtgOjAZnxIDf31Qw9qfADBX5c63JbFwSaAupnE8qbNbmhms4vJW9OmAGNaG
Nm6M9tJE1Ix6J+VoVbNhapgmZNHM/SZKZbskiGWN9910F/8B/wy22kq2Qde69WPh
7x9pZG4nkzubOQu2X70wsd9mb+/nS4bG+zkggjrI8rSK1r8j2eWzKwY6mng5u68K
BZ5yuLRFaybOciXZ0Ufw4bBa2S2mrL3PBZ8alXEupCH1DoQMkZ87uHs3z1TV32pW
Cl8sQzQNgc8l4dAZ00wsCJclcVzmR43UlrbZ9DrgRRmSH9uHh13pp/KEeZYUX97s
zSo4i6qzyaenFhpsrIGeB+Lo3z6tw16uqKP6EjKZIs3I1PbYEMfZaHjQz2mAm03K
ONLfztkwoOIlhY3lJmTexPrt4GxdXLkM386bIZOw2rdZtu9BHwx8Gzo2kV+rz6jN
Kj7+DetBOCiuNrZH4EzFPtDtgwgjIGTFN6iZ88CMhrg00KfHnzs8nFSGWfceA4Yl
PpW1ed7rs/CTn6TbPVH5qQHT1Wr2EsDcKWvhe7BoJIDc+mpobaOuWtOo1BZ+xyVh
AJ9JvQd63BOVaJPH/ViMuObnfTkg1a+5Hbr1yfP89FouhYa9Df4vUKmgc1M8M1V0
JULk+jP00cqERdub3Mv10oclRun6lLM0Gm4spvnLdmykH6NPv5n3MXwS2N+4oII0
NS+lDYynw7FfXqgJcBwdf0nXCp660LzdjiFM3N04R1b30U8RbQRzjgGUy++zMMgN
EnwlrhqWouL62U1VzDgGJu3mKE7v7cRPNEpwTwOKNoh1aajhl5GFx0/wE5xjQqCM
UU9mBo29n4KmjF88wBkzk/Ip8XYieqyTOsbYs5ybImBbkDZ6cupWdI61Mq6+iG0U
ijzJUsKcc7dQmd/0xLKywh28AW83r4lQKn3Kl0ZXWM/7DrRJKnpeeD6wOVWaZ0At
74/IVQo5WPRl5vDtuKlGxhQShRLQXRZNiLsdZ8KOdE3wWWzusDjD4ucjbTzIevu7
D7BtnOeDSGH+GezChkGYIxqfhpJ/2wg5+TLlIn6dniePVmNdJBKS1wdUDrXZZxLT
3UpuHKfb64cBWVHXCi+96LdfRHZyDeMtY0LR0b5/UpSZC57FKt7oXdWuPghyC+dB
2+/aNnq1D05aUVbWmm8NlbdzV60q/ku10EQBNcTPgg3N2vqvCt4weAUD4riMvWE2
2ONraNdmxsod/l5Z2ObYAlk/qdQMnnEKxD7wULXswG+fVff+C2MQ5/CO/BziuOeU
FrWuLiej/SUqGxKo3YiisL7TZbvavfDTGBRjtOmQMUpa0BuaFL7cJSvjR6HyEds4
MBeoecxcpjr+K6fcrpbFuF2LvqXWyS3iJ59vMjytgxlJh1P0f7pZL5sKQfgKgccG
Rzt0e20B/HZ/DaI7hCvcHQObgx8HRvVLI4nA7chnXvRi5w60VQuJOmCs9X5+HW+T
c4w4XLQOHmWK6/rzFHCXpraaaR56tk/RgcaGt7+QOgu7RhKTapLCeWCE7oTX9/0a
QJCFmZVIVsjtdXkcJkqKH3Z/NTuj0fy3j9eO0H0Dl7LXm2Fws+uv/kVeMRv5MjAe
1238Fr1Miy4lypXIkymMTvxXS+i9pcpM+XNwMua/F/awyoSAR52zrljNKnAmXSJg
Fi06ExiP3nQyqnLZQHsPWFjsfiKuvn4FCf8ulz5tx03yRGSNZ4v4DxX5Q4cmE5iA
vFmGFYBLreMqUfJeq5LNUviaXEcRU2o008NxRyZZfUeoxYmuYgBjwzYPzMabpJZk
c1MslWp68xffNOLA0UrX/LODt3eDDeBPAvoanxOVk5KsagVqf0nMBtv9NvNOj0u0
NgbVFTw3dIUAZ25jmeZVocZM8HcEEMf2YhmH7Cs2FTRv0jB+w09u3BnhqukeVuHO
nzcIU/ISnCAti1CczTdTbJUD6jTeIzExw23SGCf8q3Fnxam2C47pPvj0I13ML7mC
skM/3BMozyo0HBWy0SY6bVXhx+nrb9Ak9pJWsxyT2aLowqXmlclSU8Ex33M9OCaH
U9OO62JdD0YbKSszz78aYrilGV81i28hO7Kb2KGP9kjQeikjnvsIEEvKowdi0pSA
JavPINe0LqgJeL+b3gs/11rdEnaRlzVJCCsVKNz/CAfLyAL3yNEeDJLmsMU9SXEo
GLlffm9RlWNYU3dLxJK8a3/DEcoKXd4BqoG2OqRmVBCB6RmAht6qmqI2qNFNT93p
yXInShSmTiFXBEc/tbXj3k7Mzi6NyK7Uby+9p1dgZkp+etNs+DC7kemNQl6qPrQr
cIh3dnHjb5G8V+duBTJhlcbayj5fSNrCCTbn/gzfW2x8rAo2xB73lXOmKROmw+cr
4W9QQrXmKnIG3DdxiPgO8p5Szcpeab3ufDDxdob1K3TwC4GwCiDvzmZ9fIZ0FgXk
tVtmGjwlY4QLdP+2XB60WbShvvyXdKqkJUsqMs/1aV9CujG+I9msWe7WHa2d1HWs
HpHnacaqjko3eceG5Jv3IoByFyrJEOIPSWzLlVzIkpNY7JWt1Ry+R6uCUBOwHwOb
1MFCfw+4gInadpeCPjfcGwS6d39Uu4bKwUnMjHKOssjA+ctZtRGlnNRH2xyyQYlw
GwZx0Sf97KVVwc2bC2QYiYtsd2LRta+KjD6kTurkjlOV6oI/Ct6SrQv4hu+VaR+I
SWtWzMZ9hlFqk/s9qaxDbvbsIAODcx04pdwRzW5VCjYnroGWDs+a65xm78AcQNTd
1Yaj7NyIDO/HybGoqAICLXhQEqDr3kdbSP9dAvSxl3eCguiPuO2vtVnn3j3trwvQ
zErSzhbAelDPXuRo5lja9I9SwZf8F/Brl7xK4yx2eO/J+dYT8XMs9RI0+txtsBuK
A/iyIVlVMz7uVv2VPeBJv9mWZI4x9boGONX0UVTq4qs=
`protect END_PROTECTED