-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OkoFsxvB6rUJfD96+IoP0kejVHq7RtatvkHDKSnrsGoTSxjRST86BtJqTPVNqVVEc5gnJkr3nCES
sc+Pl/Fh5R4iIUtCCqKaxvPgzvhiOzK+hgYRNQeX/wJea64JWYdfRKd6PGnlkZrx7F5FNAcoLPPa
7zEDBOrtdPXJfEiVUMeRADxEmClq2pbS7dbezn8KdTzYg546v78tCRlT5l3i4ytbWkdCRGZdAVdi
4gkzC++lzFBXVmothq5IquNQQqSUbodKc+zOjEUfnX5H9SS62U5ygwQKU/eq1tKE1cpedO7eQvma
2fytRRLFIOpRtTZd99XEfX2S/fmDKa7hX5BD/Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 36336)
`protect data_block
eoz0f2guJT1vwtdjPyUjiMfMOnPMOHRi+Z2p7HXYhm0y/x2UyffFFt6+RIKoqhgTB8TVW3iSJ6Lf
Oq4438LiQBop8+WS8NFVBN4zW89qANrPBC5YmgBhP+mjIoaNC7rXV+sOJ7zg/5eU5ZmOARdQCxsx
AXwGJU8dmR8RmiOcMg8GUA1D1GxQxLlcsz2wvwdg/3bQx1cFiF8un5/4opvhusAY3p5777cinRyg
gisKhCxuEWAkFN19XpeawWadsNGrE2K2rj/N7dAQPPV8YsWu1OrYOkKi0Lw+85bWfB79sZmDvdIz
TwGvQKzqK4hlzke9z2QQWEYsIFDI97sajzF4BMUEc9msMb1jXCHtRAijwcZLwCY1iNkQX3aZsdy9
jUX3HtazK8fBQhVN7lDVniYfYP3FixwLRsjlAma3HHAIfzcmCzBKSu4ZKHi0pUj2Wwqbw8ZZwhoH
XpJPOo8XsByW0Je2brAtHkXEjQhC5YNFInyVAmT/yiV5R4Tt+FZREi9ZDBKpMjfY/1E2zCsYRKUY
J9JSLmJe1jeS6s7C38gRKvZtDA0eQfnM+q5qK/qhLcTBQFHOd8CpywJj7uuvPuG1G92y/S2bM3TQ
c8RhNEuKzL2Svfe9n6hbkt1Lg6xTa9WorW26zM7p3ti1BWenBtjFvYoL7pUft7lLmGETksB6iHBe
7OBLmRoubZNOoEN2vPqw3MwC/oqswoLP2BGNQAM1z/txBKbisIXGENUpkZABdcp3Xggck6Fwy++j
OswUXa6JKH3hODdiBfSwB21WtV/cmX4HzIC4KjSnjCiDeHk27/vxPFrKpkf1zpm+xMS8qyka2ni5
H+V9k1FS0gWAgT2K2KLhsucenlbOrA+xaPPyvj84G9S73tDBy+/p3T4phbIKFaljcALu+YYdfOav
CrRFjELmD6ej3r2tOqdkhjXvx1dYPaKMcxIMkhasMSCCqihl6LEXay1nmnSJ0vMi32V0v7k4FSZR
QDJRI/JgOeSR4J4U3ciGIAseJMBqv9uiZdGdxCs9m8690BKjKs6rJDhmw3mzfJVzeMrn1vKbWGxI
ScAeCShx238+EtuyYdZeKeZT+L5GimnuEh6UYw+APPj7j/vJjOIx5mkI5tE8JU+vAZg/zs0EsJ26
KuoYVt5qGxIK1Mta0NX8Db5T39857SvFuysXiqRyi6Z83XquuSkwOaDCGkUK7DVCLIkCHFlPMEH7
yQD32ZblAvwZcZP02Aqn07Vn6K63U2C5cRKVM2DIVkMXqWf170gjsDXKm+kGnztsbiPfZllzh/7/
If5+HcxEFJc65kmrseQJhuniPxt/okPdYsN6iINlSr566Ln06buRqR70NjetViec2JOQ04I/Z1z+
3qmtxNNyja5CsGkgFZbYXMMWMWsNi/Mae7+v1L2ceCOUvefOrLaEE2vA1oLnwMLCbA//pWil+x07
6wOcwhjSeERGiyDBimYb9XongfnHs9LLdrYnouDAxbBI5YItzZJ4tuU/JdyeNPyDN2ngsIzZkmg0
dxarhFpc8r/hGVCBzBy18HKrK+3qPVSe407RvXLpiQA5NMzAeSzfL0W+d2YzLVHdDF9GEIAx/tuJ
aG0LX0lLMuTK3FLWoso3L3F17m2NvuV/w0pkLOtHmFRLc/cRVYN6U33jnwxF22C7vneSY+M9sR39
Ve3WORn/spc/wlzksWQ/x2d38Jl5vgDWGYx9lV7+YrYa2MvkyQTi4lVbPMFEouX2X00YwtVaqa+B
YL5t6MXNt9tEdM4W9o+muu1yWXhgpSVg29IzVV8BdtiweRoPmbGFvFP7XwMbpKWGrxwRiqglKBte
/Op5JivgDCKnsvsmRL/zB8R8J/EB91in7ergXO6pqyqZ1lASxF0LQR+1QdQujLhT3bsHtXSTGQ3r
fe93dxztb6U0pES6QF1S9l8a3v2TAMwkqEf2F0S1egphcBV2zcSHKUvYkh0OBKpUeSIut/hQrelW
efMySeTmpceRHPiewzoiQ3R+sDmimpXecAlfHcFjmu24/M0W5nvPbODtGlCYQawGvLTeg4PB5o7m
ErxUKCRZpOlYCz7YbHH1yoKaCZiVAjPsXwq7XblefqlsSEfQ8Ds/oJvBbe0vcE9CFDysbIyxjfh+
b4hjWrer2NhRMQ0h6Qe8DYfAxNQilnZbfpdrTjpBEWP7cMUK8kGXC5BvjR3BoHDPeMLcXwYG1pmx
Y/maLAv5Kz1bP/VpzUstgJrinihRqXV0kJdsRCcx/0tpgCOirm+sFCYCFahmzR24/lgNSCkQrEcW
i7PXB/2czNCSCm5+JwT8asIpRzOTbmF8tNP3IE3bExlOWtcwFPUATnefDsLPMmZdnEbvBTXAEuor
a6z7jRHOgtacRSMG/m8qi1u0GX/R4PyYHXXD9f07KRTbeyRj1il7UnkYxIzTf7dR89sR0DA7YYFF
tKFaORQY4ASYQn/wNFIKqznqvcH//qvq/y55q+o+F49HEtdVmszx5PBacu+BwKyN4mo6y6poRKU6
PzgWJ59pSTAezpF4Kp/xygkQaLRZuhici5FkTED2W00PoSSNj91k/MNFgtPcGqk08Bz4PS1qatYd
CLVzI6U5cUHHC3WltPbys+v1Ql1ZtDtV1bkWl5rp7PNDTNxNv4IwPVYtChu67CR2Yw9F18wxBG4K
jeuMulRKiLAK877yZhIjt1ndd9mpRWgjlytJzOJcY7ytviZqruzmbImsNKyAwRlXOeKgc5mDu6Nb
81IgSMgj6mrd4IbR3L+fMKE4d5o+6xU4uRIAMsB2SwpgYqBnSuVNwhrQ1PnSoAtNXyObp8767SQ+
/UcnewmfH6QBLRNoKRQDhmMqIT5Emp00Z58bMp5lre6VBVjMjd50Z42NRDVs+njHghUfU2OiCOKK
iBE2eOm53NLVxzkpIblc0IqVuwyDIB9IPTkQ31uhql4R0MravzfhC6fxy2UULvPAISrFmj6KlPqz
H2O/tXNZ68l6B2TXjGaf3eLdkWS4VqYmhjxQqD6rjtpQxC9blNsgEa+SKjYYCSWH4JcQ3OQHCp68
jm03RJqG3K3s6aKWesmhgtSZ2aDYGTE/05/Hd5WXnV62jCJvyn3L/FdtCCaHMQXkpaZNpiHW9SYh
Mb6OkRlWmbhxqImkBZJc1vhrgAi5SuAknjraiSR6nABx4oe8LaHJUSHejkOgI7OIPY80ulfjnvK8
EdYXBPJ7Fj1it5netmtlY1nIWBVJohuiZmiovfaf3abP+0TPnDnE98ikLPnauEuNYoUKZUNItEF1
2LGjYs7g2NXqthKaNfv8MwfwC7LhFqhAAuw1/hCKW6rsitSD6UcJI9QFcV04k8MuDgk8elbqwsW0
K2ji6AIi0/C7DY7bur8n3KjHzhYzM4mFNuPp3p9sZA27KloxXDqnfVWVqv7kLewtcDjc6JYLTZjE
bvjrtOSvptP8EC1kc3P8RPlNkdg/6tfkFC3QcAeuscXHqFuTRRBcdxDHByxMYl2uCzcpcc20lb7o
evQecgtoAwWx3/LPnVDZqQBWqToyHZrt6Ux5inpSoiht+XUDN6vr6vtkyc6rLYxmnwpX7Tdx1YpE
lVVp57sGBz8LzgNOLv838ElX5pUDDM7gfYt/oDuuUIduWVLN4+uH1TDebqE+2KnO9LoM9yQUUKUc
h6rM35MdZiw5H4O8gp+aFu74tDDWq3TM8sLXc+9aFfGxykDOX4MEHDzR+44MzCceU4dL/REfWp3j
SjlyesAi05H8YaUrW85G70IQzgU93bvUPCvzPKytTpLr74ptNxMlyemPnpJKZ3kLbIgXbVN6V9AV
ozYvGZ39+IcPcOk6ZNTQsS6eQVziuMn/QamRtcaC30Qo16evkioUHWbtSIszJZH4RAxY9H5+a0lF
kgvWz//eYm8mT1ZlM6rnoXbpKYTXHb9NELp4YS+4s6R/U4QFMvbZMaM55Eld7QyIyrGJPj+h0wz3
LsOpQ4uGeV8BGjDDfSf2zCFJOG9N8xPhOGTBW3mgAFbBufwfwxwMl+DcBXYp0gUjU588dZ3xF8/J
OZGzU/hfzYitDh1JGrgBfQRZYGF2KHBWYe68ngpY/ssBk32YZ8325IRRpQSdq2Ok9nYKNBorZvjR
pYRF6za4xcIW7VaVK4V0wLcp0InYvKCC+eLm3mDrfyk18t+rgdNIMDbOqfZEzvXW82JONfPygQa7
+WAzNPQQ2ttQlPSzGrpcJpgbdhTzBgTLwpRI3Q+O7N2fmc99EzLo00MpQjnI8AqUd4kBDudHIpC7
j+r9CT5XqfRcHVH4GwXMEi+TInGUBr0A8dxWzkYgLXyMOYojynMfXtSDpLky75upgvfQ5PRb2Xka
HZQzvmoUJrvDmQjvDCRxX3Etmzf8X5Lh43xTBv90RbN+e/Hlpil/wQQ4Ai/vHWkkZ2QX1+mK8Pfo
V/fVSb5gGEhmilEyF5tzJkXJI6yWpvn016Jp1CHte+umAd7thbR1umOPXnYVKQJfuamFEU44vAsq
Kp+C3nbDIHBfBgTwMrJXqgagTUZiwpN1fv/BDzDMb0E9RpjL7P0s20gCwnNLCbBC3pepRzBvUxpG
lGUx9Jw5poOuARIpaOAEb35qHcOkbl9zPrUNr3tQ/Oiht4b2p7YvLykAVSwvKRw1HyRBTyw5++oB
aTY/PMPKajTTWOB32YJT3u8Y7smmx0iPhI1P1/Y4nvck2ZD1JUYWN/VFpsX/Fo1bSWb8Q9vk4y8f
EJ4LbrA7deBltl1maWZE/YbFt0cQXby9tC1BcZ8qDKe1xP1dVIBFiJNm+IgH9THlEz7RLsXZd9hD
2kYUyP38g1XO8U6aCKxccDeOes1pGB2T4oYvcAMAtMflHQjjAhDi82DIqt+8UC2ZsVVsxf75i70Y
25mYYt/ul23TopDjevJMgnZ4sUIwTZ8Wk89kWl7gBfnsDQdNnjqJhn82+Mfh3nJODDmwDtHjPJB7
uMZdU2Aiakp8WbNsERaPDI7Vt2sR/PcwRmXaaVjWNJX7qgSVjvIQSeMF2ltxvAzqsy/floy8OXAL
cnrS7A2PFR4+1kCemiwLuFx6y9EN1G3wRx3FgaKIM8nN5YYDlQmdz19lIy9+aOWbzV1GPPuq19r2
ttNKWpD4jJEwIc2qNBZcyHN3yCl9876RSA5p9G+JF5fBF1z5c1DShhZmIC6sEkEFrdvdBaasZOqA
IR8nWP205AZiZMJvaOnTAE1O7O+fys3kQsZWnLu5S9xP0bdrj6CwGjRSifpA2Vf9ub1sz3v4isxC
0Hlz0HK+H6UK4XdILISYnnt+fNbM397GlTs3BFcoMJDbIB5Xen6zjPb77JXcqVORwaPZTCkM6hhR
0QiBBNXwFztnz/r6GpXhH5PToUCsfhqv28f2I5x730bIibnXT9NA/dFFzJ+KxPsmSL22D6cEMDui
qcl7JapYOf4+XK8VzLNriwsx6Nx51q5rjBOyx/ReV24vB4uASltOn3svoEmHo8J3EJ50bPzsCr/T
vi0dBRudMj1sgDzXirnhGOOotvHttjAQg/h3ImWiJ52Y67XgCANv+xjCOPiYEQLrhleHJJBhkeYv
nt6DMokL9+wkjdKxtEV8RGL2U++Uj/NFtnMYqndP++p7lGh20hFzEEiBW3+MIqOCeD+q871oBnIR
KTNuGhfOW/CVDat6zgfYO+xblTiZFypGnCvsUZ7vpIySKCNBVvB/OImnHey8BDfWURnVt9J6Iclq
Wi1RTDLxM24nfyG41Mc4AbX1hv+B/lvvLQlgwI9flmLQBTJlyXt4uLRLydd9VVj4ofMnVYlYGiLR
sN5V4IBgxQ5lIzQ85o8BmCvdiCZxel1v0EBTsXeUpsE1ACCmfA86RsCaqNrvlpl5wz/rypJSp2TI
uGV9OXdtkWdnND7pOdJ9oiz2+bANaHTQeD36dI9QY8paot2jyukhKDFPxmTEOKXpX8B9KslYDe/E
jBcqm/JepMH2K+vF8Zi5hvekvJuyRUBD3v9Md3myM6AL7zS0GHqXiYLRaIn7gzgj1xJfeEZ/AO5g
cBs5wxbW6tAZ8MV55pohG37ON9ZOlEGQNha/298ggSKKd6gEObKiw3Uty3jAj5sWIPzQ5If3E3LC
1s7yCcexY1mBcF0ifdgRZqrr76HUMVMuJUQwkI3BfKfDf3REQG5eP2K1qB1JLk8p33vMe9GCxSTU
lpRaw1qjLyCLcBAN90mIlIT1STO+CKjJ84WJ7ipyPdJpDG8bloYtFeWyLtlziRF3G0txDr1Gj6Mj
CMKvsV7yv35ezpP3Zx3HZHHT7uuASlUFolXXcVDTyhAjpidZ7s6FY/VRxJxCwdjIA5+v2zrJKn6d
WiLuz66uMkHt/VJG/plQ8FT3lJ28JmHUbGQrvZsoVg/3fjdOBmuVskfXydQWK+3sL9Ig+HRQkJ1B
RtC6Fj3kkZvqA8ZeXVI7gj+0nw2b9b568wDzjpqs4Yo/eQIg3ibai+69WZv64O/tqTsjoiq/TrAd
OEqrtd7CjDztQ+abyaAHLKURJfBQ5yBjdxtZAI5ENLIVF6SjBfExKEZ8LTLdf30QxJ9H3TJdptGu
FZi5P2k2wgsvshEVbKta7iKQgl5uhAr1P/m2xmC1+zkfD2Hp9BgQhMf/nO2L6qiAu66efDmWFksy
7N28XTDVINARHYV+E6BapW8y9xNsdxsUg7gwuw5xAKN29FojH9lwkzq4sfiwznGSS7qxA12RI9HS
P08AAjjC/m4meEa3oherEe2J8TLhSur+2YYeJoIeYGelnYTq3jKBTPo127jmrPqmwdaXkGytgltX
KCWg5V7sKLvwmU+YV/JlAKr+cJ5WXBC1y4ITZQ8Gdl673iXQDtJJomy+wKnVueJbSaI0H08xrr4D
6TFZbSFgjBnh6QocUM8rGydOhDba7CSqxJPma7MrBNUSYS8qXebgl/tUg2a25cDjwK4QOh9oBIV4
zZaib0jOlrmDvS0YUzsuON8p/UNccMr6W9MpfgC5C2utei+o8hLxf3vBV/hhvZddnj+8TArUaxxz
oWD1ev8m3tR3b+UqMQuCzisLBkl1eRdCkOkE6boe1F0jqNNG2L11aNY9G+JZkhAmVMFb8qRADkOy
44bVgYcoZSLj2GVBLkMm96BaX1E7ex5myHwpQYTIUZGHNatRxiYyUyMNnRhuHD6luergRdQ6DccA
66/S1U0HBSWLDGRebGoeL4xlrBXqWSRqy7x4qyemmnvWj4zoxSNxEse+Lzvl0/6WK2oSD0Zw7/vW
VZcYkxEU8ok9Q7bcNpTTPpLR/Clg5Ayy+Cl/iCElJuI84DN4NqiPZKdWSd2zOwGBj/+kvDTnBBob
5oJVIqKu77TMaYqzudWRow7OX+VAFWtlZH3R4K6LA+n2LquPi06ijWqHb6aFV0oCjCFFaRLGMC2s
BxbCD25mRbTYumv6DyUhwKuSEr8+9rZW04aPpAhcMODkpLhGc4GdxjyOS4d3u7j2GP87PmtPYdCv
hFrH92dT9v6Lj9XtYCLQXstEDKYCjTwUVvLbD6wCz8b1ddsNhp8mwD0ABUnlYUH1TFxNDHpk6q1R
NBueE/4exOcFz5N4dRIpWh1ivwt9BDoy9dP1CtBazNmN1r3J9j/M6dVBkXpJsaghCNnrLeBEwKAK
T6w5BTNVcW8w/B4wKB0odDIBM/KlyarOQYYnvB8Mb16lq2VPqca8pfyvL5YsBen5rwCpFg5kmAHM
5n/1oFXwLdKrkD2pcUx95H256AGhL8w7YZo3d+JdRLiLUJjGRu0FnHLB3GNOuIPqmM1VWfDQMKut
xgHY/iqPlnA+Z9B/S2nkAaScAv11S9Lmc1c51/PPfx4HpLbZl4LD+0zQBEN9m/Gby8Z2M0ofI4YL
ttaDeymlpnnBQEQYjL8kC86fsn6J8etZH4Zj15D3PMmMxCzDLQ/8ezdKLTZBU8GO4TVokdGYNQIq
zJStH6FP19jxsBvXPCbesiG190TB/3kC3mU0NVY5dzTU16ea0MjanHDEySd1M7nYj9iSSO9x65uL
uMg415/7gm9yDADpUvJkuqEoSdHTZblwMo+lXOhxz0uVARCF/Baw58usc6NLF5avKIqS9f0Nf1QG
fBnA2ogNh/4TMqg1OTS84neG3Ww0DXnWXuKCyD7FJ0HrYOFMxZ7j4TkaB/ZlAO/msUL+hipcTMdp
Emjxx4qXKqIjMqPrkJKquR6mcuMs+aNszSLDa4SWHRC2I+KSMx7r7JvdEz9sutP7WTQZCTiM9rDG
yFUqGb8RUKH6gbQ+f48/kFd6VvRfqomsyMAyhkfu2nN8Pu/m7BDYa2V1qkqUs6hZADmAugaOquaY
YxC9cU5/NpgKGlV+U2JYeKNgivqC/bE7Ux2uBVVbmP34BhS9qePJbU1SeXZJ7QPFScgEaD0Uyjdb
7enL6VGBT8GeggxLAIzSgPZqrFGMn0yXxFjXh/LJtDunOwARarSJfh8c2IGpR4PsHii+bVBkmQ4/
mjTwyaaoFoRkxMZ5RnYUEBdEFSKuNRiHKK8VfS0qx6iAQuYkZMGHs3ebkgvNLGFcAYsmWOp/oRch
G1HE+bm+jpNcCUyE45koMztxOYXaf5bSliYBlPEExAoWenJG6gYgVgar58vPQ1AcW/kqA97Ve14i
Q3u7eEdLQxqjJH2eVufEkyeDNf3zIg4bf7lRBVSPmBXSU9z1gbH9znKagnnjB2Lwv6WWoSCtZQvj
lXLC/rJJ6Hn5IWYYwFNJUGr73jFLwDRWKofIEK8fifjtnYbYXvREzbvJuzq6KkcrHgsAv/COyB0K
bUq7OFQPtcE5KlSXr2t1IXNSq7yXAyl+EV8+ROHBVs9qdK3wSZJRnvThjD+atDsFK8Ubl4cBxRWM
w4TZuOQRpUs04SBbAPvdKtRA4JK/K/DUc5SApBm9fLnHJzHeXcE1aJamGpJXJXvfAgxWrgl9s18B
UOO9TuvC9TRQ4QTg9SJG5c3Bg9OiRJeSWNro5dibf/z6xF0O1inm6ptUnZjJvEOCi/4JMCeVZPoI
EIn0r+VONG5P3Y1H6BuAUlEW54En+OzaZjES2qlrSwsJTfZeEp1h1SGbTllqeX8sYbx54xR8pGv0
ThdTrU2zVy8NiIaIN/bv6dJ/EQfIZ7tYjJQ17e/zrspKDUQfIsOh6kZH96xnQ1ksGUuY82PCvJOt
ZEs6LhLRq8SwzVYBGNiNjq61IemQl7VO+CmFFLP/L/pj1tZg912cGAsFgT5VkXq3dI/RIS9v89dE
DFaJS7160AE68VIQVdIpyHM7DF9rbw7RJKkYCTiwIG6X/zYFvTbw392SFDEVNmeZAA8mkuPTQP82
0Z+Hqh3Kg6geJFg0ce3Z3XawYoRvbsjNp6hT9uM9rNSmPTeWldd6k3pHZMaMvQ0YUlJZ2+l71TDE
KHsC4KA5hMTLKdCGgClJLWAB2dfLF6CqbXM9AxuM1zFfHUNSgwpcHbz+/brGsAbtT/PQ/11wbP+N
pSDKfiTpBEerbhCQvfeNrLWCN4ZhKErLu4HXs5lOIGvpqTmfbl6/JGbgSfSByx4zSL0R7laRt9U8
HwZPLX4LzKGVackoSx2e7bmbd/ZYK0h+5oma5U5YnHhaRCrA3MlqYOk8KMZaCWHqH4zmMtWXGYKG
Ri/J82NG1cjX9OzO6UGStZnFwmIUfZF6HQE/bzRGT6g24gpg543cQjXsOkrAUbYoJ7iousCmOkRK
ZA6hYu3JEZBJQnZY/mxiZv4UKrtraHzIqfsSlfP/g2QSTbN9xhgOGGmTWs2m4KAJZdqJf+qc8BIf
nyF2ej5ISzHYq19Hv51FkndZY6WfsN36MveljaWBPXT30A5aYsflbO5eQHFA2JcDu1Jb9tT77bnE
zgwHV4pzo9TyipNNiDYn6A+b9aELNh89k42aaaN/le3kKyKZMpAdGls7addiQwTW0bFV6SBMbSVl
6sRx/heoHKhUUpLlfep8JOwjObPAf4xpdNOOOK/iCLQBO+N6870UmMw7Jev5v8hWsgyQSKZz6GjB
Rtp13A4ZuBg/kKetlOBEJKvsyvPcVwcBAumBD1Whz/xQWdz5zP2Vs7Mj4rfxNSUZMx5j8gelHN3G
i7Gq17FXa3uSayildDNFrND3OlpcnO/EUxBAdjDNm0f6UJVxkl34KnGPDzQKBnW3Lv5RsRst2K1d
+sG0r/LHpHXtui3dAH7+sO9exM06SwYrAhYHHCBWAub/MYMDpQkmBSM/CCytuvEpEAY/v0qewb8R
YC/Toj4uzWjzEfp80acJ8VZy47WWzN9sVC6w1Bez5u5YCNaY0IloGShLslm79oh47+WtTbwJd+Kc
y0Cr56+Mb6Tk8L1ABS8k6WyV2JvUzrRAg4abO6Rta+REeqg++6kepmBeRANaMrPIwZvR10xkdmRo
MAN6fHy1BTug/K5NG+bq+hXA5/APjum6+aEsBOtu2qG4TZDiOIU7/cRBGIpJWJEAFdfn82DmmF7A
Utrpt8b0KEu3cJZ2ynGWoWVf7CnfTL8b2tnlcF3cCeX/sF/iDYGYzOs5jg0Gl/ZlT6t+bNDIBeF7
ww+7mGqkOW6fkBFUukc9/KHDcCt5y4q65iOoZ2ZhumaZkrV9tdrx2avf68j6TlT+HpA8WsP79rg5
IjUpoQUTQCw1jY7xxF3XBPUcXPnnU8EGWaO6mpXNQVsX2iJEecoZ4+kp+5R6Pt836FDgXwbwuJnn
1+JUIrZGJLkgIsunuqqn5r/04roJlHCCZWECuAQjfgzPWXO534+0JAn2+LEUHTtkYNIBDfcu0xyQ
FTp1n5FT9TwvHvY3SWaa/VNq32cCfN+dZTyJUSef2SkgCpCiDi46GdUFvqbDTSoSM7IpNGQ15nI4
P0+DeR/cqWfKl1RZGlc5hhWEaqXQdU14dzLdY5arU6bV+rvnh4LYzZleNo17je2iMZ/PEDtYqIRK
UrVCO54ic2U25dYV/LIpBym2IbiyiWAXWWATbrnZSfwArE+wAFp/GSyjUmwpDYkdswP0eyjuOK98
2ZjMuul0aRoVU+58HYRH5Nl7Bcqu/kcZGJiYIhUoD47WNgq1UnISUiHq7H3duIHmpmBYpXrwcepU
//+ixfFXg6dRwFdZQ3S7xXb0EEv8itYRgLME0R1WC7D4Fg81pzrm28gAMEtmbW/MM4C1d+gyROFn
x/YSgJjYRD5NC9FLhA76nY00uMa73/5YEpK/SndM5nqdL38F2vLsGyzKX/1Ou3F92lei9XbuJpcR
Ux5FgGdiIna/tjYt752uIM62yJga8fP4XaWPpCRFYoR+czudXcUBMK721H+7vQ00MXIHdxLzApNu
x0lLAlj8fOuX6m6P6U5NMHTG3D7WGTvjKzrSArYw7TRytrpsOQ6PhluIJZ38TdjW/SUL6yPBTSNN
KuITA3aWGCPh0QjPks4lB/2j3bkt0YMJcc7X3h/lTLkSnVOg7ZpuNhjJX11ylH4WBduE2Gu0DyMr
ZJuFVHwjrOePCLTHt6FgnnsSu12+iZeakdKl22LfMLaXDrXKd1OaEgx+Kv2w+KxhT6G8ixFfTutW
MGnKYOioXOYphrzxgGlYu8qYM3OsDcfsiJwJG5pMOaaFhVFM/6GZBqUVCK6WODPJ8mJ5P+dA4tWa
LVkeAOYtiOJFxIKNaL8FUnJWmx8Sr2SGq6luLXNh60sOkoqq9XDiQEa/1gul0EBObAxZkDt9a/MH
vxJOik9qHd1BVKsX32CQs04+LlVq9rIX2MHxzdSwQ83h7xX02Z1PtTVJPGIBQ1Y5DcTLF0kQXSFb
IwQrMv/TuhQ9ER+p+1ffXgs0scoqcJ8Pcva2kOaGXD/CJ0y8whdHr637pRdYv+8D7ztpHHZsuGKR
2eSx4m9gsg64EQ06bG/yqttF+PxDLXLeKneFNjx2E3uyv4lqzlLfp/FY++H0cm8cgVO05Njgbg9s
WLdRqL0SIvuTco2df/tOSi08Z363AgioUefAqeDtKIvo3K5GfTYCN+D58kHP/XitHLyPQ9BKe3ts
WwTADCaZ0Mqe1hpqOdc2WTTkQzMFKOREXXlLX9rIoPC8vaHGzoCDpCPMhGvKDg6OxaqHxlPuXVwl
AhZvFhnbj3siz8F+emupFerG6INoXN1he9hpYs8m2jNhIbxbAw7tOfLXcxFbWPxer2xJasDqJ11C
6urOaXh4RVomh0og2LGhXAIZ0eR4jVqHokZjdvbEWRn7jA38tRWdIeQ8QCgx6dDP51EgV5T6seX2
HMPxVPlbkgDv5F+0AJGzrozk3uQvKnIhc7Er3UWdgKi5/vkgn5PoJXvHQSKw1Zs3nuTXP7huIgHZ
yZ2EYXLXQYh9mCZ1xdVuOZhs6qTCZoclMWEYDOhnZssm9isPU1xFUh6llekXrgcYH/6Dtw3ec0vv
LN+ytvr8xagHJinPO6pxOp7ZF3z/Y6E0z1jME66nEhWPDiUZKDdIaYs2spcTEZOljR632Wip1jl9
rs7+j4xmhhLEvv9BRDZ+aAEG/ZVubOLBKvDww4Um09aonuDBsBsgVMabfKYd1i1YBxDNgJDZgiIJ
qhnRPm8N1fFIkchOp01clgpFrNRYxBfpqen25E5nFIrlwSgFzxP2if9Bx4Yu8vb4xNme2TFVDLE9
vzvgRNAdswCNEnUFSjw0VDza9Vu3tqhaAss90fOBxLpYYqe2+DS7eCuXhLJY2ZgekO9m1PZCTy25
ekeKAPBFoZ98Pm3fESAl0ElTsdxcaTkL8Rge3LuVmwlYkFaPxEHX8syxRQszzsLh9JaDdOcHo5WY
hEBFwgVNXRgx/qa8tqDfKcCGjEFbrG+p8clRQRYgGXx0E3hXORPet+dcAMh9L00Bhi7Q+Br6hW0C
2ELCJOa/M5uAmumlVVepZoEN/cBw1y07Dk/v6Dtn7sNP3W1EQdGV3laatcN7MPyHjJ5PQKFkkhlo
1G8ZECIRfZ9vyjX6uofuSlXOeT7b0ss/CaRsKiXD3iB6w6IDuS6nABrAGhfCL/xw5TDF/e9xtH7+
tQhssK6SlZL/IYbgh4FXJIc5yDamorEwNRUV4GtHVJdQk4J4WWcbFFdcrrceirYZadPt06hgb0vF
dmYjCYOg/ngvSh4B07kwxzfcFKohear/9hOZ9upM+YC7IG3aA19eM2nEZdjSiHCutoxMwuK+sYzP
OPtmDPiGi9co3KHVmfiffgBO/ojMUHTsTbXzroYQe9N29mtOdyZAQkR+g5ihgn9Tf/y0j1WH8nZw
uHDRhMysqG/CZyt7Heyg8OYQgiKXCQSNChIRk9mm/jZnk47US9OVgainYw+qFCwW41O7P/IJwPpc
Vj4OWZVzXRGA8+tsDjfpTQSsqvP1yYFIcNJ9D/spBIIikeso1eA2K5TBDzxBCJWENbcJGULxyeCV
w2JacC39jKQOm7vxqMg3hMce5wZEyXmaBdp0vsCTWinT5oMftA3jLwajMN1zw/nE0ZEGVLNgn+cw
XEQNWKe9FXUi1wv5nQxR6/xGReTL8FZLs5cLpmyw4ufGfjIDI/VgqrgMeBzMAVJkTjlwvFHKzjFw
GLYnljaMnnuGJAWrXuORdnIylX+5T5fs4gcKBYUoLNA4U1U+m06IePMv7S3qovUbiymw5yKswufs
FPgJh5TbmLSH6ZebxwbhtjKHonvVvahTpBgJZwC7X/9s4Q9C/pPVqU1ADnISKWkiLDdpH35Kwnei
ffraB3gn94Z454VItt6p+cWak3LTQIulIKn6eJKNson/xh+GVdPRq9G9GmwLakCRZLq9mDTx8MXW
GCz8+PEhnfibxg33QqCURSod8EWtBwafkgwcMTu3CEnbfhnB9RA9b1AmuDdLCjMt6iN+SCtihCQv
RG0OzgJ1d88YMJvrV/KmEbe7z+M/FsivJdi5K9FIu69vRmolPPiRv1n2/Y2TvQaYTNVaNz+UIlRr
KDTex/W34ou97OOJ3zPioRSpbuUHX0FSbwJ9qi0rxuypY6T9WhNEvUtt14JYL8AHwIA24ttvygt6
UWrRYeEgD1FLj6iEOWPqvRt4FJfCARjM7h+LI3rOKoYsZ3ww2T/GSL913Qa+wYExmvkm5wb4qp6N
MtX22G3Ab36dibOMb/xch/KlUg7OIhJ/0qUdMMhWwFAtAk3SFt1LtpRn1zAHNVFKVwpgWaB/++0Q
C26UgrF6cc1jTI2KaJ9vWGTW8u5qXFT9rw+U5wXdpraFUmxQi6ucjiVgVMqBFz4180chExdkVUko
Ng1S1sJtgzEHVJXUwvkwQsQmZ0hLePzWVD9amOhFPRo+nRAtl7X9zLtd87JDJLIwoOn7HTkhnoYB
VV+qVJEMqPKgB3/HCOlcIWIP40UWu0SCsDEVkz8smqh1/r0cQJSeDxIvYjzt+iOsgT9O9KunmInk
bey7DHYPIHnBrf+4npoYQK6mPAZee8ULwMBWE72dDTS/8TK3p7K2FBsg68bbCKWDkgnqf90d3P8C
YNrPQF688Ueju4njVPPZlpj8HFuL/7wvhRml2Ko5YzgZo7B2/JjcrxePkFzg2QQraQurbwbn5H3/
yB0gnmq/D0ypLK8y+Pt56fGk1WG/yp4q7mhJMc+GJzhswYfIaDqyYjE6YdaVJhvfhtl99GVUEWLg
PWshuIJ4n6AyttTZeRaLFXe366eGSeWEE1YLMcYG/3drLq1AztRLztFI0N5OT/NwQYtzQW+54Lel
PLFe7Fil9n+56kogZrLx6UeJlYNW0o4x9XA+wKD/0Cp1TQA501mSYJyOTeqIqjI3zE/GkaEfrg8q
6tNovzUYicxBTIAaB8nX3RW2Osvd36i9VMVNWN4CLc/XdTwu4BDnqHiIkrauVg5NAeQKcFDxWfNH
NOvW5w4SDsjDo0jDzt+/WW7I6pG1uZt5SyxxnN0HjRDhB9z2vBUT1REhOa/pCdwvm9q1d29hNdIJ
nDF1Mnx1y0j1vn/JHqcO2Pv2BrBhZwd1kplATrgpHsm3uy+lhYINFbwVhI2lJvK5+naQ/+KMa9Tv
QRWL5aeGBKCmUrEo5YVnmnTxEegFzYCbWj45FOGt/AUh3iQoBmNfPgAajnLRuTfIi2rHNrRNx116
Kixs0Y+0qtiXffXzGYuCbKGNz+akPli+lqpTg8rKvL0zbJ/E1iItnMtBclU1C5y/U4gUlT0Drlax
i3aqJY6VeDeh8qeSuYvHAkcc3R7mPppsXQzngw9LOW3O5Lrqxr8kqgyzDgucRfREldFeYjh6YfMF
adM4SZ87pcQzfWOKI4dW83U/O8DRjL6hYN/5T0SkgzypOpZ1s3gkeYCIm9BB1RJgg7iWbLsn21k5
pfQGpY7AavXsQG2r35Si1vv8+qjVmbuL/6Yv+tRtOmm10SQ8Kkivxlz8auTN7cyUuvyIRZlGNbUN
bILt1RudhPgmLu4shThCim7d+WdMfEo1AhNL2uFDt1URn9/yLUVPzRT+GYFapJv6F6nUC0GMk5cH
Cc8f/4DqqMBmZ2ZHAZ0gDrJdsgR15eC9NmdeZHx6PUc4vsOYlqkmYGXNdxOa986foxHuhiGUA6J2
s/VAtWBKoAIc8LQSUoVpEP23bzVbLqA6MU7GApBx0i4vKr51GNiCcOfAl/jVzKffxZUYnMTroxur
moq/BLi6tL6NRpNejEekqBxTDaDJo7xutwVzLs1HzoJtzmFFnO4W2noFcuul/+nzbIOjR0WL5QvA
MN47ORVs2pgwA30U5yh8F3xPCPoS2GhwkNKjDoYrFkbyLSAfRgxH77qXyqe1aLd1ANgjTNqyR8dB
8OOLHIpPPo9scho/krX8KFnSGC1+cVIRu/jQnrfGfiyH1UVVCOiiFjgcjbgSnDvO4F+LjXHsdeuB
rjBM2GdDUcosChwFAqijsvWQLW7jUAgOd6A/I1oGkcp8B0Furt0ObozmwMef2++jOeMyxqYhUUGD
B0suJHPvgusS6LuIXUgrnpSpr+3tRINH6q4X8vI9FlgkOZtpw/3UZi1KeINUOBzSPJmYtKwL7bo6
vc7NuosaZ8wd9r3m8GOgWFguuxpgDrWdFLKLhCAfETAr7MrmHPJtPxdntcvrA3ze2tCow/AMUsxI
cLBZHw0Kl6qKaCxxVAKcvWxxpuX+t+yI/I2FMJT5XLeX13DmbhyunR44fVYckTF1j7jN4bhY9KIQ
gofDaE4w0l+cGE6Wi3HnlxRGhdjKlA4tMNifIb2SFKAP9ac8a9oH3g0ZYJ1QB5j87F9m1ky3Cx+j
rGMmMiG1PZMUuiL51HYAJxI17K1pUZ83AqSKBBS3pCK5gDB31WPqz8MGPk1Nc/nqCr+zJOw0lGF2
bMvpawsrAKBuhpt+4TSF4tShIs1ET0Ep2J8e3k+UqaBWKIWFkJgle1kWlZ2zwLouzRBA+5QML+h1
JXzEkkMidUl2p1B+v9dzDtJ7oTIcYXt0JQ31US1dlrt1ZQoszmRsj2B8o2Da6WgqunKUuTx66dXM
nc9++4H6/Z5LfizMCi7GbzbihG6jWwoXbDAlcU1i53THSnPtIC39sYF/hBAmK7/ahPvqpdSMsgZQ
gZ0e+cV0FNiTCGKxcIGjqYJsDf06teMMmaRYMrtjMuGtDA8Zohui34SdGaj7jzZ4gY1hJeTpW+ES
cxdyM6LRPN14CUddjZl52weRmw/CodFNFkmcQOzHbmuV3wH1sVeVP8EKbnbCujlxPtoBr2gfPpdt
hZQMMjYubPIMORaj+H3WlpmAqjTV1AgL3c29uDHSx/aJUJltNsr9kSy3ZtN05rDaRRsQdzN99BHf
6S5K+glSMOyxjtuNx3L+ATi4mTh3lhHFu0WOFsb/9+/9vWFj5zZ95Ba1f9F+jqqIXdSuIpFIIL4B
SQ+1PT+slLUQs002c3tA4JBjwG9H+W6UW/MFWMXdH8U10mC4xX+eGrWn1ZRR2KjRYUfUlBUtdQ3H
bkxTTobhL+KzU8YJj1LGoQT7JHCG116w1hvu+kJEYxLHvbU7ftCgpP37Qd56J17E8FStsX6xSSrq
wlnio5xsq/S8GVGJ/Z39wpdtnuWckYGHG1YgT3hnF8SKbyA3vn8a+hsmJaHP6L7N4oVpVHJTc2Ra
YvyeX4YZLqHBwdjgT296sy9RDuVy0M/rW4mqf+SNvnw2m1eR9Y+gwlKN8tq4LuH6dSbupiXeZT1R
Jx5hwJyCkaNa0NUfte3FmheYJ25T2wBYDIzW4WayTXFh0yoMqeN3m2sKQLuSJIYTrnjxICPeMmm4
dN/bcfD1RYFx0FySqHez6rl9js61TimXJpI4cns4duQKHSiENkxQGLMZwAzGJVD79osNvRR43CWv
mOWUj/jURy4bE+yj3m5SXXy6Xp0SCALbffk72fuTX1fyJQSlqCacFqXfXF47RYezwY4cniS07dvF
F2Mrzh0nGpCkvituzXLulvWMLiBC4VkWltSjzi47OTdl3leTU2jUpdtris2nGG0c82lTlL26k6t4
EFVn/TjYuGOXkzenHgY4vmkISdDphUw8h/IuZc5auD1BiXk/agRHCxcXQpC4na5xTsBqNkuHPAdT
IPqu53YjHdaE5i/muC+bHkQLMmKQvopf7Wog9q2qNvNZ1u4iQNW0TwSBsdNgGjDTir/s4GApPDhi
hg0aYy9liWRJX6w9YEfLO2TOaQa6DTOLtEo2cXKs5ti/dI26tsSyrUl5QpB00DgDwxuxBRP0+PN6
9fEFazstHi+psmaaAT51Uu73Vriv+mBq+grbpcbMuOlDJNGV4MHKa18oHvw/KFp6wZE7ijlZzbhA
zuryDMTh5PsKI/dyqzsHZA4aV611W9roixiSbfY4+M4GvWBdAMfTLCz8WBvJ3z2vYHzYNJos0oF3
DtrdJkU0tXNYxBxxEejDTdaDPi+Wgqoyb7yuRnHqh4yVvgcN6NuJeLnqddKvS7xq89Rbg/6ggFxH
6tduVVdWCLuA+lPM+u9SzS9zkPQPUlsIJwGf5ot1+XFBDWGmXPitNIBJL/t4E7NVve4r0DIGvMAM
zL6ugMqFmozYW0FQK/Zv457uUM11DdCbkicwtUchAreVofXkyqmuY0DMAs4aAYVnWVTCF5rRiA2S
RDMEzh7jCWJABxJj1WpESegHBkvwLkW5j7vsN56paKkYq87C4ZE8MSlj2iBjIGxk8oTGApVHUKhl
XDtF4vWJdcP6r3aMVkVL9kJr179xam+QndfrHWSB3oTr1irthp1pF06rzloTcmfoy0n3cGObq43a
wrbtdX+OcmRIFhGnvAuVQOy8MPmMeEBbTKy66SO6M8WBYWm+SXAnqlSmHwdw55rpIUOvUc5pAAjc
AlXWRzOt5LgOCKTtwWOPNNlGStaB0PjORsujL6vVmVnZu5FraiHTtbm1Y9d4NC/Sybb29SmvEtzP
jIFAErtgO0+p7HlW3fALZmDov5TdH+AT0PVXgxKD3Cjkq/g02ZVAvNfo2KrgVwWxo0XvttmgNrxb
3U/NPWqTBaHur3NgnQzM4sGxn1aRn3v3amItD41iV55GKopib6iqETBdOkYaOozfboUdivN6JSa7
wkhMl2G0fjhv67HzdRyeq6A584nBmCWnJxi7ZRZzkhrH0a0z62JqMi9dqWUF04T99yBCuXe2w771
qlNfpLL8fOHAFgxKm/ajJiCwA7LyFo4YpRTPNG3UNZ1QISizF7I4smbQAYWC9n9LN2oNxOvIZ/xM
KNs9FqRQdCKOrJprtKebUwlxHUcPV1Vjvmjv8KSiIcJqyXVlL4o2uPqPsARknpvkMwNLNCO3EWTi
wz6g5k8X9LGYJnXmYpCUNMdwwkYsTKV6BgqPluouZMvNTYN4vFdJNSosgQscaHl8zAoJ9FlG0Hpe
1GQ4zZrfKghGk1Gst0ytpY9l85DNYxgdTm0PhMHqIRk0Z+9LswXSbXKaihJqjDp2umfLtNvlyPQT
+c9zqghjBWqQVZCdd4pox/aVXYre+LxJEFdhTx/C4fhfnwtdIbLemONNmdgCWbBuLanMhg4tNZ6z
E47DDIt76veCZBB5yjv+l8H4hzT5IjrxE3sUA/h9b2FuXRJC5YfXIaI7Z3VxoVkWSr/cGUE+vBH8
q58Z6hyROr0T/mBHJEHJPz7qsi6GekvkQfT1AytP5tG03BODfAhph6M0gGbRm1/LumyV4CNocQxU
tO8EDvP5HUJ2XFKhAwUX9+Xeg3YAUUctd1J4pWWrBA0IJeS6XJGA/FXk1zUuZqExs6p0j4AP96o5
HY4wzrvFEBwGFdzI9PpU0oZN0m8ZlweZT+vGizoZ412jSw+GOaaN6p5zHPFY025OmbxJ3X9GQj4o
il8fQz2zVsMS45MPmP5CCLAdpyWyhw0aAf908ojtRfONbQ/VmYMCnFmWk83v5b741ITeCeouTbC0
j05Qe8SYieABzf+xNkijQ2E30O6ykWdKiOSPC1zvXn5vWxEiyLf1V00Z4pKJzxB6ibOHI60O/wAN
1bBSuAOX5dT4CUr2B1LeweLF0JLk8B/1+Nbplo9fLLyDN75cU/KBn/Wtqjb8TXWF+n5GQMwHWpwJ
88eIgnLBJnSZ5qlgFFr66wEk/j7k41+wIgoBUqK1+Dz8oM1GHm2WHeQFb3ZqnhYNQvK98n1RZady
N46iP4A0mrD69/JNA2yzhTKdD3Yjwx12zAEwrOEZS/zmisacpNtqdUaBYqNJ8Qvepg+sUjCqVK7T
c5junnXPZp6lBI6wKiBTB/DvjchnnGTdSU5EKCTozBbuuJ9quArkOCt5NyK2/OIc1TV1u0jUDNZH
XSvS5N0N8SoOqHcCbDwCcz7ZtphpMnZwtJODjkzgYYb7WRIaVGCo2DR4vd6N1noH0hAcgKIOqWDy
x7j95uoMW1vQfuxOXQ16xg2KqldZFH/JjfzC+p5bSp78WIRVnA7AxWPX1UkaIfKjcEzPAuHR99Do
saYBUT1HrCl3EFAVJmTyOYyWvlhUa9YrRYsNTbXSKONfpZaOL8LjngBBlz4n1uoYx7EEOBWgf1TI
mO1leKvTvhDd37XV+UT8d7Aq2w2q8YCE7tWV61kNSYr5f/F8KTAYsGfZnzESOM+nHZxYZv6coL4p
RiIe7q+pQT/GoRDqg6JioUOBlpOGxaLm5UoaWDiKQy/6Zpdtg2sI/EQA8xGhDGL0qzC4MUOyoOce
LC/VUTEfXpaMDcoSGq+5kO91L6NJIOXES3gyJ8OJuAtJa9AcBr1pj0QRKkBN3kw9oFwy8yGRJVlK
gvm0oJA/xsyw5KrcYwL6Sr0AEBkJsuvu76Ps8TnjIxnl1NDsiWMQFPs3mx7vrPNLqyZer8xZKywx
NlrGVAp8lNnuRCiigVkzYFyvaForz7TvgGuyj3RA04J+cpNPOreV3NgegaB6MhNhlRn6MpLXiieO
IbIbbsGekaJ+FJLYjlAqVFPyaQDRwEsxF5pDn4qVDwNgdWmooIL6kiFNMOpEMXazkCIQdykKRT6i
1MOtt78GNvJhUx63bEKdX9xMg9uKcw98ICyVLg7tXrnzEDffZsdwh4jmR36PiRAGtqjDfgQSW4rj
K4BUS6VruZCYAcGs3b7L0y1G7W1fE9R8///+H3xQfAoEvYovOpdw2Xv01Z22A//kU7WI5EIwIahV
qIvTRTh30UQuvStss70T43eIKCwt+e4laY4EPSpDmrdEkqohuYGgYuVSERVBD5b3pDUl+mSIkv1C
LLkEHknW4/rkKaEOFD+XlTuTckVTpS6dYWqx/5H3tcK6cMArQlpDwe5gZLioagCRJ2PN67twJSrD
qBycXPeeds2XTFY47+IMAZn6nPWdj+2cc+jAH2HxEav+OwQrPW4W4skGlAlMTCxndSr+qvjbhc/I
matPclWvsqhKD0UGf3HtEBxzOIgNGOJAfjCUAyN+vgGhVDum+6gyItZGR2i/naCTV8mjSXvixHfs
NHrnjbUlvg4l4kRkwnE4ngRVAAcbVdsFz/WZ3nzFwEzMcCdVFpK5SiIF6HRrb/VaHZInz9/PjVDV
nWN+Qu+lz2SWMNLmfOFEZYDPa3EdptVNciHz1jZisqnvSwhPznKKixCwuuAlc3HEuNJoSTyMkmA1
BAmWCQjTImRz4RtdOcg8sm5fJuE9Rv7WmvPYXpXXa35Xa6BF6IG39gfnJUE33O4Pkg6KhA6iQFHy
DY2CTwyMqVewrYcTyTVp3oR/aH7d5bOIpC5QWx9ge8Pol0qY0Vz/RPLiUIGEzo09sK8Nk+Vz4BR6
skbz7c+k2j/L50gqTNdGrFvezGkyVb2Zfk/80hxOu7WYozkQ76dsaCwkG1dBGGAG4Og9Vn+y0yVh
9ABP3F7mps0G+BbwYYBlDpAFwYtOEnQcS6DcI81GtwWxLoycjIFN/IS0JnoTTCmh1sChBRKB2xzg
gr+JFejz6KcsILEY+RXQdSkaE8ma91qwCNAEvT8udPWQSTQTepuLs9H1efdNtKZsTkEjivYEyV/1
V+4MfQ51BIkzVsohnqOEShnqsB+oiH7qqqJ6Ck0ej47jY/PvowcjgkxCPipgWf3u3qBJfPvXEnPb
Nk4Jx7a++kQLNEAj8a4Mag39iIPdwn/12GhuEHVBxD98xdlnH0MChAP7mGyg0IBm0Nx12C4kfJ38
5xxh0ofybw6QDiab8bvEWQ1p7DSEn9PRG/j7RXwFZXzSxUfDz6MNB7060eX+3eXB5n4mo/IpsoZH
59/T9u7nvGajsUl4+th7uXu5bPr8svlwdyibPDFAaMg+Bj0KPQkoEt22rCZoHQRKArJbGXbL9+Gw
Y7uHepT6UoWZy+VUHeYLrFmzB9A+GSDt8N9Ey5BfBtGu54pSMJmy/cZj/dS3EZ0DR1jenxLNXspE
voGN8z2ZY008ACtDZroYB9cTv+0Jwi70uDrlv1RfgNd6s21aI3EJH1H3irlUBZbiOb1gfsD10It4
lpd9hXS4XYhY5M2NqiFTvyjWrfYL/N2PQhPBOxADfbOq36eOyhueVZKIIWZcg2Z/G0pC3z88rZac
TBRRwUbZyH6GCasTu4lp9Lk0EVqpbzszGBWmmm4FnOn8K+ZWbcC2hzsdZVgDxRFuvKXOmOzspKAo
0rf8w71iuWfhIH6ccXtvqCiA2GyjViBYIWm33s/zmOYGNQ3v2A3L9990bbAldqZbwqH8dCFb/bQK
s1qYcY8FkxoManrb0DVVbceOtmnTsET1AVypXatXJI+tUeltaOVs24FXLCZvr9jALTfrb0tKL5P+
Gf8618HpxOY6UTUMy8HMhEGRFtcRwsGvYMGqvWkZ9KAQYx7i7vdnTsgpZygjEjbcd0PIYEkoB4oO
dYnmm2EOGkLMejLD3i0z5NJ84OSA5NA/NTNAx8H9pw43/ivjUoNAj1A0S0Bj5Oqt/pUVI020yxwd
X91+3LgMKzeqm9Oz4Hv+Whh8EGR04tmdggzPqLRif7C7Iudy650n+Qrk8Db1BYLJQwlbeeE1ytUU
M3ehXK6Loy7arxiDPBTEkQ4XWzJkR2+Ajvj5XzOGorgWqtCSVPT/X97peAWpvlPDlxbqYixGJ0kw
w1LE15trnVJm3cuglIRg8XBZ6mmlaRpWFV/tt7x1WKrg11xQvCtw897ObTZnDd/etEqTUnXe9nIg
yXPHg2UfeQG5p9BrnW9OXyDorXCXbAVPpxMd2dHpxf/u0sHW7fQCbJwiCMpcSfClTUHKrY4IQTDM
5Dh5T6uEUJ/zWcF0g9acSoWSJhQZxs6v6hdquSORmJjsc9oprBftENoZqk1qUHaONoZ6fWx8hmEr
oY4PBzEjUm5kVb7DPhzXJjK4gG1J4g4Cn6ehinNJV1/NBEh/1OUn6zkrasO4iF5Dxa+bWyYgExjj
ccWqILnAUwNjJSMXD60CiEjTep8HiulYvQInz+1+ptEqf+YC9Eh/qcphb8rXNW8NCdPcNhHLv8Zs
N2gW4zwXNrW5PK6zuWJBoSxj8PgsMTx+LLPhSU0fPBvEcVoR4rFSA1kAgkIGRQc/zVgZ33Uoo/xM
U2jD0DepKnKG0GQTyobeAGHyj5//JZaow2xbQSbl6XLAL8RXqDzR/liG6ZC7tmrhkgPvI9r4QMF3
Gj5oReHXdCdDaP38ANQZKO4OACYlPy8k4onahTlHV5F7LQUYUDTGEXeUiepw5zDuEGGLNDck1vOv
6kq5l10Qoochgi9vK4a3Zo3qqnvanaQrUjmwrjOLQGolM1/AGIl2Zc0Iah6Vq5FT39PinZR2xaNN
orO6OQopYELpEmNf9A52vK1mIH6j1PF0OJHyZTPAezGL+HPs+WBViJWW8ca0uaYYfB4ey848k4yb
+qxImN/+yzRfPiHMqeJXHCHKe3gLKRhUm/BvSKc8oNDfTVephTxDx0NDfSPtd5sxInuCCyzlSNIj
J1uve7ai4qsRsNPb+IYHZ+Q25DEHoQl0LUeRT6rVvr2IO8HRD0pol+I+WPMO4yZV9hdqQ56S/fC5
Ku7qf4RJKrcuPbIPqTWENabvjeZ8eJG+uXfh2ziCNVLhfsGsIng/sXt/MFT9/1qcpOxr5QXpn4fZ
Q7pJSNGDWvDLcdO0Zr/yAUiR7j03jvuKWJr+Una5m19aPRz9wJJnrlZaxSKW7gdftl2H0PKI4EOM
0QJCivI6p4ivva6+LxsdOEThJj+vvOI+RCmL5abL403CTLtwNK3qKeV5EgqQeWyQFfDJOdvb1ok9
Fz577lKMdwAnf43xx61wv3oNXKN0V81v+fyGZ8qusp4nv8FemEctCdoW3BKmG6zdRZZ/LaUKW9MY
jLK1auVARIuKd4A0MEQy2eARmDMimWSMJRpmtPFHqr5pyrc32W7WiB94dL611usFv/on2lSHIixS
1owDGvSp0FcTNoNH7scZv6zDm/uyvyqMu7FViCc0CqjVRZh8jMf5IdOW0vFnDvkJOscRDzCLGxdr
ofJ+6cMhw990bFAbs3e+s0R3A4TQgnrlz1bE0HeLIUGzn3gGJC13ow7hdRl83PPjRhAhTjwPWDpt
U77Cfi/3D6MDRHMcxG3KEH19X+6Kx+JRYmEqSGrsdnJZVTH12DqvJb1rZijuQgWLmBLMSmrvGIUY
vKjcWLkULL+QUFKiP+Ast+BMSxUdpOt52nphAqeY+pYYY5zF+oKgLf0adB9s67W1UwMvOxsigrax
LIE8VDUKGKTMz3F4IOI2NahZF7RQVXyROuxvxVBZIgyStI3fHW2NO65AabyL/ITq5fXrT/mKoOU0
TWuoM6qUXcvAUiJX21ul13GJrd5ubyfVoeF6YL/Evs+zszKUmEih9ncKaElVxaSM/pFL8DkCbsMn
Gtx7hNsCSG19cyIER9gnurIUCwT39kR3TSgWAZaI4/CSkpgzYWr+xY1EtXSJUDqyWtv2DkRUuND3
qcgF31Q0bMMks0btDBUdqLMfdwg31UcMM7UsTN/c85ayYlrcfN35bkXYYq+msBI73ldAJkrz9MNQ
5ZD1dFE+wqCVuoDewJTmXY4Lr5rq00IbYWU075LFqo+dW/fMjhv9LKkHBe+kOlrAiRVSQaqIozpM
MM6XqHw3fHiudwVRfruGHjbBqWgFlVsbO//2n/gAXpzVX9MoAbtBaXRkJKnW5RmEXJ/2Bpbkjb2Z
MG0dDD/J0Rn1t2HKP10H5xu1/i84vLCmVNrpj7G6eKeeUD62CY/aESoz78HkDV+9uflNCXSf5Y/M
bh1OTsX91KDniKTbLqhr9bCO+Wd8Yp7Gb/PX91QcXOIiHsQBsGHQHsN4vQmKrz/t/mhSnLKbccZJ
xQl0LA4gNTBnb40QaLPBb8Xr6oxJ3yeHdInrzLq3TWfM9giWXT5II0iawvM2RHgKfXpHvsWIv8MZ
Lzi7Ej9eFyDYC0LR6TnW+92tuxwDduMzXkcAMUpRvpUwbXdthuI6VexbwXAsMNg6r5QqY98eTH9S
1QIBiK6steOzIAciaK4DypmOm/8zfjfU9G2nvxZ2vC92LH5yfSojFVsz8jlcdn0FTwgSRZRzuN2X
U3Xgof91q2Uev7OV4nZuqj4aTVnA/XCXW9BdRSp0Aji70KAM+bF0KME4VCGfiNs8YKdIlaEKoV8e
e00Ra2iOF7eWhQm8cx/2KjJIJYCB3kWH09gugDU+mktJmS73l+j6xReH6lfP/HHPUGg/mHKuiPKk
bsrnb66BNniXGxTiPEI5DoS52kJsj00ILGr6EPV6Q69EK/TFxxLLX9YfmTpsQ3PoJalntkSHtHKV
ybNA5RMbVb15aVoTSOmfe7XYqN0zqyUUpKSGed4R8OT+e8mFfboObb06NHCBvNqmC/q+e428wRxS
GB378dMS0czH16cmDNQJ6wXorqXM10Z/yaPBjsZwoRzyx4/5M2o3iuJ1DexhOm6hzKUAcmXHCBX6
w0rb16iHqJTKLQwDlOWHqOMc4fxQ4Jij9aB/Tmp4YZDvoJTaFIJZ7ZpCULIiJTQnHDYQ3EoMLW3I
gxTaJ2vGIzIIwI7onYE5viBHkhEJnpwhOgQKE5mJmg5gBJsjdyIRittzJFacDY2X65UP3B16rpXd
LrAFi26F5iahz3ixHM6t+OQtrsfcZJ6XQrs8/gg/uFoHOFbgBmwybBar3XpGaUNTgVqS8fcVzYdi
pwu1DROnB55E1mLQ//tm9/LmPVmPWIFYRIkmMn1ewggztEWSSsWLYFdAOd2G22NuNgfpxyTVCpd+
yC9NmX2b5Ues++2luNwdPew+KfsiKlor9p/sXnySC8/hfD9mxjSHwrYFi2afMtVAc2sVhU1T3EAZ
N/fllItTOz/iUB6nqceBj2ZW1GdysNYmK+h9Nf80qPDyXtm+GHr8UUsEdNyelpZKZD8KYI24bWPg
mFABfZMTsda8DGw0nmb2sG0F8ip9wrz84xUBesFfVEL4alRjXP1roqsYZxBWIlPxYpnXK/geYrbp
DPoXOt6tOy/bDqAVzpkSq6IkQIKRZJpg/q8a+LHxqYO7hVvBUobWasahJyIHf19NdvEZ7OtzVmvP
GoHok8iGmFXM5twgCo0ZT/Y5XPYvSunxDfor3M7uQZyI4Sx7RPi+JHRsOEy++Z+ote6Y/zOI/NY9
CEmpdUuqSo21aeS2zttARcs/hM6o0h2RwjMOBY8PoOrH3XLPes//+jU9MVMcXa8IHLdshbPjwqLO
BApVp9+v+3rclPek3FGe81lMdCnLfGUdHaMLtO92bH10zKSbTDTE2QQeuiCuIdlWLF46b8Ypo8Ev
1vu+xJ7ttCpR8eURuHbq4Cy4Y8vQa2InVt24mCm4C2RANVd/d4spBtf+mGnDlKm802pabPYFp9p+
SuKccwiJGuQ/jfZ2GTNLa6DDRaIYZVDdz+Izhvt/2khfBX0Xa0E1Q55KzrE/4drxyeiKLpMT1/TD
BzNzLM44/LDIUY6f33miJf4HJZl6X8LJwFn5RkVJgWvL2nXl45rnybRFHJGXUiAaVEX5nWWO8eq5
4MunJO7zw2kUSMRYiPT3Zm8/tyM/Bmv0rDvTKhbaSmPvBgGfhlcauygsuSMs4T51cAtjDa6jcP/w
Mi1emKsHy1m+gzWIoergAdjObXZzoo1m73scQwqXh/r84oscluu49mvo7y7BzPQaX9LI042RSRhy
c0YdctnRXFUk6aaIS9v+y3qFgcQ/aHKjacth3SbVbjYn8QX99WKg3GHLUBhHPsaOe2gmDbptpSQ1
/8PkTEJ9dfKa4CIW5yR5ml3gfeCCCu5hjXgC/ch6EIShr8bWCPC+VGLObIkbGJVAuscUdXPa53gj
jJcNvQxkrv7um1wxLA7Trtb2uBTdpYcZx+xQmx3T70dHXVX9kgCC9cJtJWGE7DOvaU7TEZCXosuo
G/ghPCl2QH4E3gtvUYhv3uGemY6uLHYfiULDv3sijJNImpnj2rYuhSHZ/CpTV8tbesB47P1k54Nu
RXKx65zDnbCu38VtEIZk9N9gUzF1Zb1J0qM5+G5fHUTGhdocLDih/1829cQS3qInWXC6+DU9dB2r
yMxDIsKjklBd+G6p44pRApkKsNOBFOjQNtJ4pzy0YKDwzpu+5ukK1VTF8+7fm6FqQNzwKR3hdFtf
OJerffEQLrKIbodzcIbEOq2FVY4qyvOKwuV+YRlNn1/oZhLIEBjhoLvHiSmpywVg1CsTtJ1qbf9m
y0dIh4wCLWf+Ycelb63yTpJKIOjgvwBDawlNY0AvhTUXuoesX/4Hw4oZJ93RKQPGtmtetysN8mey
PyDTeqY4yYr/SLRTu9ER0hrud0wBD0Au3ydNrbrc1HWFDglgIYoLZjE5nT/9FCUbfpuEdXnU5s5C
2yahyA569/PmhF90TZ0QdiSHnAu0h0+LWldLniEoM8BUvIsy1fb/eh6cOBuyhnyHVb3LG2cJjLWi
G7bgqUbB2z/TFBoq5shTY9UDTXqdiRsMJhtvdHHb2bn2S4w5bnFkpEn+tSke/izhQ56T2hwIYgpB
xPLqGeAHjAqMW3SFEbHcmbWokLkkjR6PkIivu2JXpjwl3u7pLM87E5jMEpPR4eFanFQY/jyJGfil
wzABb6uX7xSh6wXZlbta8Cw2ogDA72fmiKKL8QUNmoA0ebR1X6mkDdbItsUE/K5ZfqmlTRtsq6zf
aGNhdeBKun0IVQu6tpGRoFh49VWAhCK2zpPVtZTX2qIFzEbfkEv57gVrhUvjNc1hotzpt61ffhBF
MqcXAkw2aUWzCWunH8TJfTUzx7FR9henVBFX0DdpNIMFk1RFtKMss2Ye+wqGoWf9rzgL3yDVpntO
1afM4AZvC9R6WC6wi7+wNXI3Nts+qCwCzqHLhgDblIM2m9SP23sAFGbaeELRhdSA5RQ6e2qE1BBu
UurW4BqgorDEDTiusRFsI6Z2Plpvh5uLRxVePxfC8aUNxJwH8GxEtYrDxk+DeUlStgJiHqmoZhb/
MlSu9E0rcuNWhp3IVAHumNojhrWVRpUIFGMBBBK5WVPXBL4dzAwaMr1cFkofwQnP5cImQ1vFfiPO
8+qoQ0AmfYQzmaJK1p+14Hvjpk3lg7nauTC5cI+Zys+03MACwS7YgWT2HgN07xoC/l+0mZ/I/VOd
gzuL7Y5tpGJ5nlrnmzVhdPx7iog23eKpfk4K6TUe8r4q7dF7Qw8GMlzkyyWGjQhQoZrpJX8v6H0B
U5fQH/fswXxY3SSYWmOJyJDtLaELQijdeU3d4HIRiTVsMhWVxJIX1xhVzpcm5pwDuTwxQo5+gK3z
iNKpPnDi3/X60KzId02BGF9y5m6q4z4j1CYFt2Fimsah0voJKK5iBGep6fNxmy+ETnKF43OpSsGM
vZ+a50JTeo0li+uLG36M7kyQM9aQBddKTRJKRWex8IR0J8K94PsmdmRbxiXaxmf721ITg3a7yEvF
pNOhrSEFCJE0BEJ1/isV8nHjefedjKuNmwYO9UIejry1gzg9okwe16OnB9nGvShC/HJvTOHfItbd
fDFHT0mSQ+DB2v2qT27HSmcp45tbEAIcPB5TtjuJtwG4eaOvnhdVJMu6xiHVND9ZzkjOV5eVD8/H
G4X9EnrwoWZPScZogZSsX97euh+CK+h3wM59kI78+e+4iJ/3N3SYB9SjrponlnHxVPatxGSaG5a+
TZmqdLdewUAbawtJY/wWbW/rW/Pkaa/taVC6ftDfxjTyHyhw0rJim8O7ZDKeibOweRoONhUO1BM2
XHx6SajSQF6cwiXYs3WvF4KFV2Qnon9dfsgpXw2if/ZdNKE7xDpVzNYggLIyFrg5dSPxB9HfsU9E
XvawD1Pea53khU6EuaXkD4CQJezbKSMsXR5kFeR4s9P0tyFa5+c1z+FwqYbvX0EKVnLyRumD5E7q
qvhgfJ2tol7JyQzgGfCd9/zBIlTxOtfe8iDehHHhf+ZRrK66pXuEngtTgDjkKdBAYuc1gmmAyMRx
IfZbk4WqubHyaowP5t/JdFEAr99M85Nh9C/IO67YBTSQwkOncVMZo7coxylH5GTC4EAo6xON/V0H
/d31MJc3mF3CQUPpQSofl0kGjc061DSLuq9CSVFDKuDkj5cIvIcZKkzoDx5a9paB2NkXzM2fXS+e
UuTF3qf1kO6OPlq+575H3kb/E9zgYzH2qnIqqctpATDVGqNKZJZXjEtTHaFGHmwaIubQWITQnfxH
NWekObrZNpTlsKyBwrRUCDc6YbbOaDX1B7I6Q3M1ADJ9i6rB44Rorj2YRrTGmdmpehxFocaWU+oK
5TJ88pyvJZ9XDAw9N3bjlHsER4aBxMkO8Wflv4ZP/F8Prq31AtQUvwJctRMgTxu/qNYG/gbZK/ns
koJylK+0U/TE8CgIaXEsJPnrcJbaKIN+X4NSi1KR3vr06ap3159+HwUPqlq+aw7V/y1BTyk+jtHU
hn/9pCi8SFvvGmlyNncDvieqHjkEcW21zs7Vo8MmyO5l3jDBRWx3SnxaZGEISSvao3eLNB598a1m
LNutNQudahMXDU7ySo+WroIRf0NAdwhqkp7uwXQCUHqne5GwgSkrhqWUGWOQxWdGLtaEK+ibpW0c
1OPTyI6AZJsL/J4UUikPLLZUtySPj9OglkuSfHWzH1NB4j8cH0lJCoWmVK5xsrsmGySdnZVx5GAX
6EeYSeD45ZKLnFUr11gQ6pJ5JRHkrNGiVVGM64SSfVdstWbHP7S84CcsJsme5o6FhyKhEGvswnBC
ASbTlHgGO+58KkUAVabGw0eXxY3MdsnNiZJKv4AR9/TE2Bc8w8ToQ+7vp28/q00S4UmmgbM4i6+5
Y2K703gHogcMFShE5Nqc4LtfNZmvU6nvMfEsXUMwE2rh4DliI/XSE1/C6GkHeOkWPCobdK+pbfBJ
Fe+De0WlyinijdW+fkZhaJveIfA216cGNF9eQ9vkwcks0IhFV8U++MbNySDuwoPB3fOnOByf49+c
g8ENJaSUYfSclMiPjArd3B/1sOqnniiWZB+Izpc+Ewaxd+RwzPGEPsCiyHmBhrU/XMfsDHrUg0KY
yJxgF/7TLrlHDtm/necemcsS8JhMI5teqP8ZreVTITUWAyuRQzy42xTacLO40WqgJEYpGGJzxqlT
MG4nKq627Ft1innRF5EJ/dsZoH5JMKK/h04vgNcPdHn6mgD3Uf613iD3S9P7reZAxZG6n/GeWMQA
bS4YN+h4vecafflFoPXfTPm+yh4xIukHMdIY2Cmbg1PUVzIeT+N3wf9K8HjsnmApgLpqVn2QYKH9
m8yMxXH3ZRAyERgM2Mxsb3NA4+E7A1XO1pmxo39ix4b9oOawyuNWIIiH8gK/NECe+2a6A0prAtrr
BnTBouptCTaS6ABUxE/XidE08S+F8k8Y9ZUoMXP0bwbUitf7lpqqKr7GUDaYCv/sUS/OoVJP9Tqo
a8vy7x0xYNuns0pU/DvqZxWBqN+i6s3nWAONbamJ9JkTixQmNJNI1dar4nw3w4ERPEZcU8HUnIkC
rMRZ3kgosSLd6r7m9KNqpx8OMk9GGBmRI9y5clF9f69JQMch+yp6IeRBUovYtnm45BLIRaYI+m/l
wO113Xp71fhuBuXwekHxj97vtIEqWOqcdyR4hH0h6qT3tojZEAERxJHIX1TjQTZgBOWB462oWvGR
oOJlxPY9f1VIu2uOsTqiFGDkDvrCOjTdG2jeobZh8HZEusaUM+41N/CvnLJNczpHjcF3yhS9xer1
HQNvob+R14gwKPjGILg5ulnkdFeadO12KCVVXAeIcPXqnXw3bGRi2Zk/Cy3E9ONDb81m/zID4GJc
EtjKxHmJA0x1RLr2GSspPq87u5hztWMkaQ8EO89Lbvq9+rEQWyxxOQFsvx8KCUOr7HZ0Aj3UCW1y
Q0u9i2h+itW1HDm9QZ5F4e8CtlvyEKx+kvXJYLlA5XZm/u6Ne4S2BXTrTwP42/0N8IlWXHufHyz9
wQ7kj1QgMeDFIGMH/IVnCvwJT0qBxn+bUHcZjU0RXbIiDeDqhvb41P3nW1FVcnF9W9DkZaDcw77U
VwiUvLZBm/vZcY98efhfUbz1AanMW1lJxyCWM0rtlYEcyj0ksvDvRX94p/X9v81HvQMx+39jgSe3
d3+8+f5mmrlf8jXLgXw12UGu7pAtQGy5rbzitQ/JETnKqBxyKkogaAxaXohOiYTG6xaBFFhYGe5p
XwxDqcnKBR+yZFGg0n0S2uvyc+aIngJ1HcXiqdB5gaEFHF/OkvNN+tpcCcX2SAgJ3eVaOa2aAbEv
eLqVx2cgF8wTgh6tXbbJfoPPS2EOmrM6qkQnGJCPRq0IsIYftIlZkJav5YzLLLo6BUXUrH9CVVe6
gBXtMCVfCJsL2DvQjplxXa0UthIcaBXGcS4isKxycVvkAsvMtzU45N5h4ajl15+q0Tl1H2agvE9B
PlSQeJTZk/vW/w+d7VAadRgiCMStxQS2+pXl9ZtJfQSI8zBqVf9xtn1ZHMtuJ05xrkjIA2sDF693
O+NujDs/iUFyHwm0FAhpIjiBEnevGTvdT+uAv5ob+Re6ysk2T7dusrA/maJMaBZW4I9yd0Kx79lE
LaBDh4GKGl+6rBuPrxtugeWVyBgWhIsYCtJMEQeh+APC7BkJCYhykdKBRWag6k6skKeRzhhBtGKS
pXX99WRaHQyPKt0/LO22+TXllgjFhclg+kXiiNDYU7YBp82ip05D9SKCToLQG/c7pFnfLeTye7LD
Vjf3VpWsAUbS40yAC1164kR9vI/2mFNF8W7SkWeqlHw3lc4F6kZlzyfyKBLKalOs9wCwEVfxLRAI
ET60ooByuKCn8IFgowhMqqpnmWpd8Y8yp+DrLy5Wm8zsGPMC7Cct5mhYQbbti09/yAXEZkgTiwCp
C0qcXfffP/3ebOPdVi3Pp9K9bfnyKw4xGwXVXGc0IiqWkOEpKjnf5m0iFD0cLTvZ06CqoTbvszZ2
X3hBCWZFI6p7uIWtZZrAnG1Ia2KrR3vo9nVvCPVj2FKSsr5BIpfx6Kt0/KZvVhFwut04zgxIFfSO
DKYCxjYDRcbwy/tht/jDcGhcvOFPhPDm7FJSCcgvJbV8OyULi3xo/BtorLutV5RkAQp5KkLKD2Ci
XsS1FecqcMbBjkjDEh5fRQbD/zG/tqWYtDcPC8soWLje7OpwxtuM1zBZq6yGT986s/2hBhef3C11
fyrA4HSjNJA5zM31wNjkk/mQCl4iO3T3IEf/Sejl32pRn7jN/Q9KfzPCM61Ldbc4wsu8GIqT4sek
jMxu6IegA6VIvjEGN6HUYUsGVHdevv5Qjsma+Wf8cSEmky/9VpIwHOxn590R+jpaaidLbuVUddj2
jS9F7InOJXWEAIx1aAElFGNic6jUVrI+19K0lR3v9AsD0I0tqK6NMecAJcjt7FxOBRPnFCdZfKyc
KrPRl7a6JemAbC6UOu7ArIcuG9tQIAT9rx7OpehwScGCjtdBUYr21gWCtp7eez0b8BnVYcMeU8Gz
DvnTppGqyyWz7dVPTuvoHKv0m97zWYUGmZ51ZPpSieeznIxgldAbCpQeIoA4mAoPEJghRGcpCByM
6DI5ISa1+5vzLVRS9vpT75kvpDLVifi4QTgKiYRl6/+excIeIxt9z49uFsiJIP9926Dox6/W04yi
nYMW3tjz50Q4D8ikHzLfZsDKmqA/DMS++jNka8IBBR4SdujZ/E09VJHk1sxECpwI+YKmvYpqybMd
lB6mcJepvOLJstE/3/jV24bdbZ5e+Tu2x1WLhkNEERJg1U47Uhfc8XLEfpHv57twuA2XIJ5PK0W5
mZuceSJ8lImKZ4t+Dv7hsGz82v5l+MjnyfJDnIxvLT35KeSuh7zFQDTxui44TxDM59f+pE/aaFU4
/cGvsLVuZiK1Rm6EFpcv/8XPXJhhJ24FtowkUtGZhiD/jJsNKjr4bt0FRUSoPUqmXCoR96FF8B0v
i3kFh+QcNKqPuNVbvgb7WLt9/4bvLP6feCPGr7dH0l4xpTRV6Hyjhd51oBAzJo64SkA6GaHr+Fy1
AxfcGRmsocw8J5N/In8Ik5aXl2rGcuuGhXIOiP6w1eSi0rWDIHju3BAa57s2y8O00tN/yrgiGOgC
lPS6dbBxN94NaeOiCClUjzPnavqUw6GcHKEH7csKukBzuRYH5aDCXxRxecNdD9BGszP88G9teimh
GjEYPGPBNeIRvNfrx5/cwyVHagM0ib9DnWoYyN8uN+ekIuOdwQho4byWrpgUGukGxyCOkwch+oSn
PR7qRTWbgx2WUScuz+uCx8iAV+ovBu5jme+4TPZ+vgMaYBQdGKDE4y24a/HddMjbBcIqzd63tc4f
gXbIU2DkSLTgR9w2+hcdWu4iVELiUJ+/Ix7iqHi81tjEBBUthYc4R5wLgxdmVZWY4csZBmZNG2qW
f5oCwHoan6wVO58kcZpQoNKknaYvzJu1YoRZgLcDJCTtFq0YdAkE6+EOsIY+VqiRe6haGhgzQ1y7
2LXjqisJx1iw9Bo4GzRh5BLBUZJ7ZSVU+naPPz6/obZuMhMJLLDXWoT5xrkhQPtNjXM7xqP+6CtN
jvdLmfHHdvKWhFg3XB4Az1D46QT/0SlLkc7bgmQkSuaHtRjnZ01hrzCen3/0LiAd61BhcPZlOc1P
K51AI0y0gfQqMTiG/EfYYdeT0R8iaXBZZMSwNy+jM3kyyZ3MQuAzVHfhGf3kzlgjeN9iu7V74+S2
iEx3+r94IWkVqft+KrU4qqYDtoOvPfdVGjE5PNrq+bKz6Tz4cx8Tba6r771/FgQJnGCg7IvOarci
RU37bs5DHYZ0+h2jW++dtAW34tvuqL7YitSFa6+HlMlADaEBa0KGityHZODG4SVJDUVCGCnAgDgt
ZMkUEV4FZCO8g6Xij2s3e3KQo5ni+xDuU1t9qCsLKKDz65Jn8sFI4GnXqtaXkskSya6bFBOsCZnn
76AIxpd82s0ChvgVIrvkw9p2EKntRMpIbC/yQx9TTaCvJqiuUESipuWkt2a4Pb5IfdwaJ7E52I1y
113WC0aacODRG87qwt9GHeoojEPOkbw92d9s712qfG8mSapL6VEPoV3IJbJK/9siLMvkMv0z+Ie7
nFYb3UqYL6EuveCcADJsAWd43kE/tgQdtY5gnxmXT997q+tqkDTPGHosXoGzsQNyPzd9PTnH06HG
V8jbnFJ51dVYWzcRR299Zs8FycFW3yNJYL42Fhw2CvqcO8wj/hclFbe4yG8REKIuX0rdzPCwGIpM
StT1tuPhHzRA9InCUE+xl7XVNxI9cgORM2wG0J0dAyHiwvDzK0ZCsDefH7dOlYQ6B1yFwwAJb+jr
xY9fCbSBe+MJeNyqx5wjkELjbLa8NYk8tcDgVpij4Qq6OIXDGOsjBWB5GjcrmyljoeVraVTOdlQL
zslzQbc4Rr+2UGWIptzoz6+ALQQZ+7Cn5+IhtJVL+4//cZ88XfTPrMbh1zI+UNdvHjHNWa9Yp/EV
Pde0b5+MKv7eNXSs5kucis/M9i8yErsItCO0N3XCGqZknNbvvRdB7tUK2L7wwGa54yl4o/JqQrO4
4QCSBrCNPAAF8lIgLI2F951H00xuYt11NnWn8dfyG0X3qbgxwpn11qJ9V6sq3PLvaCc3NIEM0LKo
j47v3ba3TZ63tmmn0D3kI+luU7Ch4BiHypMRUbqCa9TQ5s4+xfDqz1FG1EFvqkM3QupuVS9oR+ao
RLm8Svp1jHdLnQD7Q3j0jX5yB9SIz3C//E2Ud/dBYYKtjCWeEVXhZzHYN0NgAKgSQN8+fNk3j7MX
R28HjejHcoC+clo1wdFY9pwAyOhMKQzbEqcsnB3pHBh+4geyKegyVxm2tssAhCJtisxa7jmUE1k+
kPZu3jKO+qs4VzDpQmla4j/XYvwa8CGyzIP9HOh7RNF5wzD+pSfc2eka7NgbRk9KjDKQ1Hbm9bFO
VJTxE1jU5A9PWyxJs3Ep+pTrK9OEQMm6FeGDe11xF/2dDTVl8+QV0TTsOFf0905ZCE+/OR5hHgp/
F1oPk6rvXD8f6O3vr6gXg75XRfrREIZJMiGG6XF/TPyF3YGET3v0mzFrM7WAddlWcCOIoBErsDDC
uVB98iBOuh9rRjBYNbSIUtaHxn4Z7tzPodZAmbh64aswHgZoPR1cgulIIoyzHDBdzem4eDmVErg/
Vis7xq+7gx/WUowakmsf9pt+rGtVCyG4MyiP4ivK7wl9WQEININqN6ZivN9sV0IsWsD3vB1/MlcG
9TQMwiYLIiJu19eYdrKjHGWfnUH9PeflhrMKXP/3tBIdOxDKeg4wvuV0gc1iSKoY+hjRpdTcdBGy
vaZomK78cghnrVxvnN2S0b80sjq9rVwItVTsvG/Tq/waTkIcnNYRNuomMz8R3KJdO52aHWxV19yc
/SC+FdFuAW59/3iqQyDeGHdP8h0OhFnUO/wNj4fSrSWUw9BVPcqQgBt70fFfAd3uzX/Md1Jbdpfy
GZ7a+iwPUw8O65UN9zckc3NhLWyBPqeEFyZO32kIB+zLUleA3/v+Lyk4aJHa5bIv6mJF61A9Sh6n
+X4C9oelmXRflfI0bUGSKPURy/qVkZ+ocz4KF14Klt/jiHij1dwXblCctXYPdBXY5qtsWX9iPQ9U
Rm5fAsgKLkVtksgnk7nIVNY2QqGsDFkmi9ShUXlL3uwPMNWttC8QEjum8qt+lJyKGdvuFV31PsVU
HyhT8uEH/kefrDOnhL5F96v3bP9CbHurwQxN7uyJnxvql69Hi2r5LSOdmxh91iFFnmn8FVGCWzzT
3x4SaAQo8EItdl6affmT5zoZ5MQ539xNi6o3aI8sKD6Z8JWXhBhUPBwzYj8jBIgRZxjoOBQJS9Lu
KWi4vyEAHpmnOO6OHfms15MQ9DTXLOU1evFgqCKXG2xjp8CIu5e8f0oDS98/fwktY+8BToHGAfEs
qnOKm4ic/oxbZ0v7jse9QG4AY3zVxp3uQt1hQDuMexYiSdardR+AI3UeXhgIpLVBSNnBlP8dHlyY
r+FUdqI7xc2UPGFUBvmO78N1NEtAUl+BBtSdSPCGyUKPMOKkvj55q0V+xWK0FMyr6nGcRbXcXUQD
hEDUv0XnlJteS9+uNKau8Vg6VHkSl1mE9Qh4KtOFluwxAkM0njAdxh2+f5+REY3nTU7U9rr7iTfO
fWIK43Nf4KnwQZZvQJknB44YdzHpyOA10mLBlT3+j1+rKGi+3Js4zk8c6qYQCQXajac+k4Qg3NWe
yvyu9sBHFK8u1aAI86qtVq9QCXdwGUNtnO0w2a/EHgFiMqdjansaL4zwdKkygva4rN4c0h41JYf1
adi64c74XPpKHBLulvB0bkYOoz5OFt819H2yFQ7vXlXTr/7fd1dBIsMkE5lP2hquGJbYXrJqKVsS
IBxONOjv0IjEfc/lSBD+YxtVmw5T5tLNBsY4+wo7Fgar3TrfVzYlVZFPRsISkTPk7ZLHxARRSvRu
Ihxh89eotLWw7wZ4tx9m/ABsk7o8odEc0lZaqrvh6ezJFydmcsyGutFMwSpBsXMvkFsKu5m5SWJ3
M9pkETKHYZHJXTEfa3D4aKMj3GL5Jpj/d4GR20ltTaurX4LIMvRs+nF9WnOjAzLhEN+qRbHIa79Z
5E4X1C7Uy9FL3LenOPNKXCj6oZ4TVP0JWM/3Kess+F1PsEPZ+uVnXJGaTIWC0Ju1AOWvM+ptgNT9
GaK0y4iN40Ma1g6hmKxpFc1zWMWuBU46VZMtPJExsujelMAH++z6ORk6Hxb3BE+T0VSlzKdUeKPd
xdqVGKgiq69EhRvF5PX5RzuEK2BVivkE67FPXfoL3onEfZgCsDEDPA/V/k6YfhM3Ol3GS50eHIR8
bxmAhLZsThBSyQ0L20Lr2S58qtlSrPsluhPWfa3MFUqhAIZL/hpP6cVJhLW+aOJzV8Pz4DXVhYaM
SoD/SxnuOsLlg642x+qqrA02GRj3EE+u2Z9ZyfH7KkpgVSiV3OdpXY7AA5TepqfoHBujBBPvv6ir
qxv8waiUDwSFsRPFdGdcxLBHHdopJd6qyDWPIBsk0FrnosM7bphk1y7roO+LT+tTkpnNCQaNSAZu
TX073mFbb7n+DgaBH0IVoKVisG2zUxF6b41WAre+98eZzFyxcdzR23NDrRdi54fescx7JviEDgxE
/USrnLEwUKKfKMENjxFwrNNOrsvmisdcMwY0yt9+mu8fiVQ1MxRS9KzGW4y8iZmZKXtrMdMs7EtJ
RqroUeIO8QLZhGslafPtQzGd21SDFXlLwcuqoSYslVSB6En4v3Jo53hCn6EJ1CDDnsD50chbkUz4
MSd9CDib8lj/X4evqlbE6a0VienOhCNrvrnpxISCrduVhIJ+vuZtVZf2NL+UQ7CiAZ52gX+PAPYq
Pyn2ysF/L5QoeD1fUEBXD4wwb7HLt1KYjb+VLw+VHDzTPtUMWO5HWmtoCyu+YDG+P4XMvwYX+BeI
1rYTbtdDs/FA9tYn+OH/fkNdD6h1a//poRmZCIYj1VmoCPM6Z2draF1oeAdfNd6amsWdvM09pmhw
YhnCOgeVZ+bY5yHXd/lEkf/e8Pg79Wi/Q8FevJQ1XRhUeZgLe3uYmjhsXqYcSBIJyidKA8UUM54g
YULlo1LYQQk1oEF5nRpYk1m7ieDcsQtXpbWMc/dq2G16fjHIU2zBQVvYwrEHKqNjB8jUGN4QpXbP
awXOsC33Sn+1BICT6xHq4AvBMFCfkTMo8ky9qyq4llFqY28syUSlUYMBewZsN9bkoD9/TeHg2fXQ
uOx/eK2UwP0DI7BVEWwt4phIZFfpltHR2MEZUoAn2zj/MUigu8c2/age018hoqkETOSf0m7oWG+k
GpQVT/orR0dvogO6/uQFWP8ZoYU2RAaI7+ugNNOlr7ORl9ler5PtfCyYfd678BecceEPFfe21Lh/
WN/9d7DuaDmB+ftZQcHXH+AJv0UwlV1+7S38qAXY7dNIif1CY1s34tTyM5u3DRQ0tIdZUdNmtSNd
RDz+JEZyLHXIZuOcLeYcd1ij6Y5Q9vUjChPDsQzQTI4BffTOqI3GBdF8dp9uWF0H0XLwWazujEZ7
a9q3x1X57LgHpQ8Vo3014TCZMNQHAUynjapr2tcPCqY90NxVNwFtlFEIblf91/fnUwq1ccm0I3bW
Qz3wE6/UohgjIkgeRsvAJUhKa4ezZqaoQq5SpaIupRmyeu6htOW7XBH0IyFkFj9KE4PFUDBGHRz4
fOVPyOOKtTbkwEjvn15+kPXWiv9d08Y9FYcS0ZYuLZjv7fdaSAL5fM1obWSFCrY2eCAu89Ghn5QF
R5XshRg6wz+soEzKgkRh3J3ZLx0SJI4az2i4Amf1Z0VG3UCbDvpfgQwcin/3xibeHQ/L0lXTYyeM
6Ldg3Ph69rTALdjG7OSZVH8LN0CSefIT9nB8glaEcCirv8BCJnLN/EESuWe8cDqGOMYLJu325mMA
sqJfb7HdzRhgABLQAFMiTP95ugDvp4MrQ7szrYQxSds8wqW5lZCpcDOy9PkfWX155l3+Jzfqx0PP
qB7jG40WA3VhkL7JFhJ429FB9wLQn0AcBnFZBGstro9RQYTyU70DYlaYSb7N6eSdAh0CVHUbWAn3
AK6wH2/9qRABWV471vBrQGFl5nKN4N0BdjcBfSU7mIPg+KsXsN9cCi519uEWMGnNT2MGKCho9zjs
583MqOGda1jkPCusU1Ux/1iBqfAGC4CPdvTN80zUER9lqRy6Jnk+aHaQUpvuG2HCXPOpCiNKpNoi
rIkazaquurkmWw9dqaVfPSGcrw90JegwKYPSjdmSVGwb0QBB0iTRvL6Yq2Rw95rze3klKDexcVjS
ntMJGibtiKz4erXDxWs2++lyz0VyXZekFR0Y/ZTZndZzTeMsHXbSa4Qkcmyu6ctPLL2hjqx+tUez
W7rMkupAX/jr5jXV8OEB9Y0ojtYJHVwWm8t5NaRbhaVpkF01qNKROJQFC33UuSj3H/JkPwaP+A7n
jUGcG/AxX+s+uxwya5hSl1wFB9KVBCaRk3E9ZF7VDZsFjnEhzSV2Gv4XxNWCsScY9Lw+INUjgraa
w8Bf/zMw1tckaJnn+fN+QCl93kPc32eLlfnDdeK+/lzgpxtq0yzrMXmYmhUYOLgcQyRMA8urS+HD
/RjP0HHC0aI5HJeIws83l7/K3Qdnj9sDm2HeOe1J+yKWOGdWP3srtmIMEHGUnSipNCxQdLrJ2+/n
PjJT2p58VMkwTLvKrjDcxV1nyiBuMf+1ZCPwMeXsDCkaC3mLRJJ74MM5zGr9rmyxud+2AB+MDA7g
mw9jkh6pwa+n2UK+1+fF2UQ9P3ro62csiqPtPup2DdzXpDTvCnnMkNb55aoiEK7ayMJFcSV+J7GJ
DCsMo5u05mAhWo1Tlo1v1PzRKNgf3t1tTYuoWYBlo/7C+bkgfupllMHqoYBUHia0PCQAe5rB0bnN
mBAIjIVrLZQGdlI1x4XMNtymDYNfLBaEFtzvjtwuaAvwWDV07bfKD+fff15ltHqpIspfkp2DMF1j
CAwUgg21YcGpie5NtSbIDOp5B26I+MGqgs9ybHHoIRLswvhNyzPf+s3uSSyt/QhyaIBmv56pYfIn
DFuDdhf4K/gAh64HjqzKugzJFmkI5ZJ+ErWac7lRombxNgA3u0U3rLS0dgm8rLUGp2iczCU9FAMt
Is4hVfxP1DlfyzvOQDkZSZlR0zcemStteKz2ni5JotAuGlWXPsxKXzoQwfDbM8nwRE5muX9kSwK2
sJYC8nV+UmLoTP9I647CTLb7EtCuqHlYIiqSz5dV/3SkTN2xmgLWKHxItMnYnIK2Muc69h99OqDl
JuLRnIdFhBl7NxY6QzAlwlKAM6Ku6/w87LhtRvG0h3/24ozuwX9ui7K9wmfR7RSvs11M8YXn2lKs
l13IVqhYTZRVJTcBqsSPBX+FWVv3hbzKt7hB5lvIbZuZqu3hjS8zSqzu3X3cbC7fTcy/fbCaMAPT
qarnZqSAMu5KxFCHYyS9hRwyBQB5VzoNoBFKuukcHO61tKIZ/We026ll5P91QeQ0fVltshjRHeHS
J/KpP7GtJpo9PPDC1mJqCDUySSzidKUEgAGC7cg+b5CS5FuTr+x0g7sA07Yao4T5zkjkMK2V1jaY
FLoLupuUett1ur0gJETHsWYY6LQKjVcphzWMmjduUGBeaSG3auMtaW10E2LbHuWoGH8j1YjJ9++5
LNptmeDnP+VHTco5Hy/mwSiOxhy4eEP13GtcsMCtcYboWHR9a9VBAD4kRwWOlL0ttrVmtV67/tz8
IYmBxvxgCUR9f4FbDbp5MkyOlP7ugtTe1svpIy+f1rVx29irWa/2zihc/h+oxhYtzCPsifVhqVzR
XgTU/WENXpvbgzFsyJ9JSWa9tk1XkmtXkp+PN20Uq58ejR1r/QbxmURxdcOCMQ/PWiOMlz5/j1wZ
gdxrrOsHm7nVDiV6w8oc0uwaeK9PX0POXuYfnvqKgJ2EHX2DiVjmRL1kXa9bMuwcoaSix/4ViUtX
TVjnw1QBjOv6AqIqedmJHDvmcrwNuls70XOTA07KacPwvOKt05IuknYAXY8X+98+Ay987kgT+bTw
ybC/b7h3WcBOb/IvoXI5iTltsJXUGcbF+Jtf5YAj3t7mS5QAnPEtqznsS6xnzE/JSmFbohVcP5ai
+r7jIl2moP1M0F3XhiDZ93gCVcTQOMOMSAeZCCzL9pFqywa2vFmrzrtzNBXC0JWQ3i/D91vAwzQR
Wd3z8ymt1jdbTNcfSX6rRD7FME47w/0ASRA3Ey5tKFqM++wFiHL7gCxeKLcti2WWi/vzetwZSSeB
nUYbMReA7ErlEXgYDY8GNHsJJjq32Uhz2w+yzA6JSi134Z3FnFM7uKlwWFKw0bzr6SpcUFMUXckQ
fgKkndxm4ZvR1b591/ixZyfuBtTJY/QamG8OdIK5gay+5zSJXApySZ29hHlUs6Ah0MSW+6eOkXwc
IXh4EdDIbgEl5VuWQEJsaFwFBAc2Q+CEQ4f6YSdRXFdBq7xlNOckSCEkoKXGUVa/NPUOnLJId3Ui
vd0AAFwVzObMKbJowv2jIDgU5qWnebJmKwYm37pzj70tUAFRakq4VhiZ3W0JGfBA1s9KECQQd+1b
jBfQcvkjD48hkZet48vUsKG7hBmsSKEN+UyrfUYKJQ67nT1aLc4178oONXDGJ2vvORp7wGaWtBIS
3vxqD+iUAOr7lAK3siWjmhYdOFe0WBCULe61EU7LstKgrSxwpXwxWyW07O9nq3VF/8lZYX+Szxqr
EJQZx24bw6JYwgOakW1PNRYiLyhcIzwJmxBxbOlIDEF1YroaNVuJLVV1U0uKq76AwxMOKFLdClcK
dqmsieggnlQwTIAObnNXRyi2RWdNASgsEVbEyBTPXenpBwg/+3A/Pbp78FITsg1KlAMLebPHMw1o
V9mU/SfWIIsyn/9ODmjoPfK8lWQP+cU2WY3atOAFWImu+FWs+YYZwLw09fHiNMZUrvOLPpm6CGRa
OUA/8cfdcN7rJh6Vt+a+EFjSOmhZr9EMAD33yoX4A9waS6AJflLAEyX8VGOVGxzmY5f17+pT26x6
qAigVnAIMjKbxReZYzr2MNuRAOGn4DxY2fM4LEtC1bFJ+vlmPHxG/QldYq1xXdjLSN6yZ531DKax
bILMxKUjF0SLxyhGDpWZ91Dblyyj1cD/BggtexkncDsM/7ufYos190jxA1uiQ99oIZJekgKKH7CH
xmZ4kDmmaQDpInbCgFCerAhsJq7NQS1+oPSEfGd7M2aPRGlfHXhzZjaElbzWqUtaWTku5/yZ+8lZ
ZDZsom6rDbYSz/dBgWyovBJDLRr0iIxPWqJK9HkQRRmwsnPqBE5VY5ZknSVLr+MXHVDmIlrNmcSK
f7GU3Jr3e7vJ/vBfH5+IZXnhRjwEb4yAMInBlsFRg3zCKxV2mBJsAU/vnO04zkIKElfi/gb+gFO4
h0EBYizcfS74SijgKQqrzBzvzTT+PN7C5cCPIRHMfpapKgPuAlMKmfuF3RUZxBEmPPJfXKiXXrNz
z0dFvOToxCoV3i6BibwRNnHA39iB4Zp9dZliCMU9+AqBlzMWfNYPwlDtixqBARw59Gv5nUsFKkpS
hLRSfRsaIigC9rdLxc556B6+9jqDoUAmSd/LZ3YcsH4+yuiqve1k//YF74UiyKDFzFgfJsVKKh11
SuKu8sDqj2IpNRxkec+rHm/UeqzAZJUCYfqSmDt+d+QGKJwfcJVOVD7+gDww5kQ7vg2IQL/XrwKu
KiewmKGDEEf5GpUqhhrLzX3KL4VMG3ylYK/sh8yFp+h7HdTEdUV+OECA3y9OlFjJslfoVdLgo8ns
8JyWIHIDJHLBfYjh6Or8cObWYHGs1lTxyaFPjMbL95CWGJCvbrLsqefQ8h0QpljBXdWQFtDaDo9+
XwLyB/awIQIfq57TwavA5sqIj6kO2ZhKXUZfwwCSOAJZVLBCLjjOqf6Lz/2/GgkOT5pWnTdMH5U7
ceAU3CZT4OamLPem7BV1CNnggTCxuw0qOMlxn9Vm4KBONl6Qn3IJex31CYdkXfgwwW1SdOAeJ4k7
/trKnhVreAXBQdqAQVFBGvTrA8RvmC/f6DeDIQAZTc7r4mXxl+27zW/Fm9dhE1x4vFgDSlkwI5Fd
JuumD4CCuQyD/G7SURFC5BMPga8dKC+NQIUTgVZczAug4i85qD2VQIRUFfhweH1nxvUpVpUWwkf8
GniL8M5fURzK+fRcnM6TB+CUT7vU/aL9AzOEr1bcDmPvwUKs0AoMBC+0L7XMLQ7HGRJUBDT5Cyos
NYJrkYKXxFcLSkWOlSJjCehJ+7v0k2/y8Dug4Adsnx3G8GMH75llw7CUGwXEOsyqQ5zXAgp4FeEX
jTadR1DYNBTr2O/lO4OBZx8gcWS6j55TRCS33/U6zl5j0wieZ8VC/nkbbYVRr95+A8ATWR43ejSq
EScsa1dTZZ/gZNkdB8246V5VlZrbFLc2Av7KPAM5SQc+3IjIzJNSaOu3rOYgOFlga54u2Y7WeXFh
Q0wqOZ2czL40gd4JdWHGMLoYyL9z8MKzPa9nEOuR3i3T6w3I05yXWscTDagG1L/1XeaiJJZp8Frz
o/Q0Bm9tZfZXJ8lDciKtp6CENKwx84Xp92eC4p+dtZJW4eS8RGaZiHsPwL1DLJrgxJvS6yfK45kh
/7QAQxKKPGkLBKVpx70u749LBZWDxdQTqpZjHOGqObki6WqbQo+ijVSdX7VZd7abZJ/t3LKGL4ud
4Cb1b21eBRXEz6Mhp2YdfBXuaoUwmgVwZXi3b8Oj5shEBom6n7bN+yB3fcpvYlHuSuSb49e7RTWa
LYWN1+1jMn/urzvNKz9uDgU1SpeFv9BtpTJ4NIdN8qhaMWmNPyjrz4XNZiBLgmr4E8yEPxtEAEon
Ac/wXjMqhS4x1ER43QncpCempf/xdeI6jaDn0agYut1PX5ZqSjq8XRCHBMXT0DGhSswYq+GL1yln
rX2hPPUxy5yIHE4DJVjq5TKFYMF3wnysgu5QgBpCesZ4QkJkTR9Ajp8ilRVu+C98j+qADU8ssfVC
soCryf9otAGMl7yo6A/tl+CqOMUjUEhVwwoEIuE/nigiSq9gr813r2zZhsHweEhpFiTTQN6vaovg
cXuUaSJKwx6PV45uNvDET9X9jd1LQkUBx7vKQjFXru0Apu1kjN7wvLq6Uo8Zu3WbTcSYeGSljv21
8x3pznP561Pv+aDf5pYNGsCjDmtu/7cm5RA6XemIohLsFQCGLSSAyDbULrTSlUzyeYXKMBrNQsQH
y77Yclp0a8RgN51v1LX1bXl6KlLNYg8PqNbzakPBqjHSFJgCEzaz0SJ0rVjme2M91DPA1kgb9uLa
LfM9fRQVp3VFofhCTupWTS+6oLvjpP0HDuJpJZF+uUujIqITHcjwBWE5GstZ8XYEEy4ZOKaW49Oe
QIayi2N1nO0T9iRFj2j0eZZMQYYn5PhqZPYLaSPrT9nf6zFoecufkhz/7PY5LHAf9oyARBmpfq8j
LpkhpJ3qJa4B+z2V7aWoS0nRaF7rZ/V1lWd65IR1+B5x6R4EextgMKIP0TACbX6xXkHnJJQ1oMyY
upzBJzfC4FBWp34eDky2DCoLBtVcilBckZaLFT4kXUYN6ptwy3Xchd3FZHd4JZ39L+ab9LkVArFH
ISvn+Yqdn/Ynf3Zv+QuWP+vVPC4FDluTOrlPecWfyPFG4C3TFWV2fiKjwO2Ld3bGJYywALAe0vv3
RkKRsFwD53YW4c+Y3Z96+DgTQtcKpn0rm9cPqJlyG7iZLEJG1hu/S66AoAWprBCLqy/gj8Ay8IBd
q7R+eg/bumEg98oDhfPB9nNeOxPNOKsflOd+jgJ2S55a9MD6gEqB50DctOamJeyCs2qVYJaubOCQ
qc2dy8eY3x/Oa4csQS6NFkv/cOnyfglyqnZP8j00ziZGdZ/ki5RfNfoBYxR96ekFKVK0cbuaKbvQ
WIIWFDba4UbPp8l6xcSKJqBWtvpQ9MWovklxWbn43Qhexq8uvRZEB1wAl/xuQ1J2d1MosapiZyxf
Aktr+qV/1ZrsYgxFhMkYVZGlIEUz2bYAYbh9vNASklm4ZIX6VqqOGX9++JQrU/aA/gC6ZD37Y4UU
lUTuXHBvEGkUdTg82wlb45CQIZfwprPy41Q3wvGcm/9JKxKT4ptofheatipapSDGcY+DCICaLiv3
TlagGosj9Q3JGxn+4teC+4mQvUjWnInmUq+5UbVa2NK+KVwuLV7+hYZ5pMHhhYtoj1icRtuUuDkA
b3OALxKBNkqgIRA0ok5hvH3RQyGyzNFYZLzuhfqOtNUG6vq7u907PP8Bh6ADLe3IO8ivCHRjOavb
LtwGwEla+5lJcd7txKX7ao5AI1GLkKN8/TX8kkVhE5xdPBY/Pv814vEnSLfNm3LF4NUL66lfO2bL
wDsHuwnaGlPaRAgVQQIH2Mjh/PIl1vuFK9dawMtizmxeOsr5WLGvf8stKvYFRiXIx/GbAzvwiu/k
PoVADTgBFJDDIjHJQQYsv9prZwHsC4O16qS6x8geDGLlDYUTO2ITcr+TMl5g+PvUmxFGVOABZmCO
CvNu9MlMgPqEj0lo9jxGa4H+rp0jMBufCU/fs8C9/9enR2IyOa7N1JsCr7O5e63a73PS+yTpLqtF
0Qc6MVydQfcgLjwsPpG2yZVtkLRKVwFEEsyMCUZy/BDgciUMcg2P1WepIAozHgoZUQYIe4zjXoaR
2sZIAeKvfC0c+KWAdBgM9tGOXMq04xP89JJpsI89VprmKJSzw/CScAAT+L24xh2OKTYGMpP+qvz2
T1ihYCdkaQl4nfJBcNBxl+tS/C2VBqSwJLA0C3T9OfWaKJCGLpxbAnhXd2XjOgsXSJs8t9edRmW+
TjYli7IHC2txpDOOpi0copsRZCquMim9yIQqJC1u01b1WGoeCvnr5notuUwwd3XPMtc/cyT+tQ5a
XFjc+7+palHsVr02Qla3PPXjFEuWf5EwiiGdbP6/NWZfLMKdVgG/LeK5sc8dELYvW914z5WIfaH5
zOfgdFFUJffMcjIZtEyc90OYLTf0rD2QFRuJMMm4u/5bBjWZ6lLReCXIqa895T5BZJ285AAmgxzD
RbmmcAweqHkwxTZxfSFLJYLHA1uW4eh4HWRVaVf3XazIeVI3X4QRejZYc4m/Hy9HMMCQFZ3R5/Pd
pCWSJWidZwSTyxmQiuD6OdgYb1NrZgh6L9EqjcErzcPcYn0NjSoomE48UTvZo+llk1WEQfzHOuAi
YEjfOVSyILfywZFg8NLKxr2hxgBcVc1gTfCDgPrmCvZq5EXlwi6Hkqg2UtUf0y0zSiaAvuUVRNVu
yPc5ySflQznPrKErNcSbVe23drKNmSetIHumtsd83TKH9QK4fPhjQ6hi/XozQcvSe0nIuHNd+G2o
obLVETMT2mmWG2n6hJWtCOZI524gMWC98PBnIpdizVOkTdn5OIJy2srXlzvScRkBiQ5kNQ4pWSHY
g/b8t4oznYODaAFTKn41IVwFq0McxPYGDAlxjPvryIz88yGIMNmft+4jaicDa5GW7xEkmucR2a/v
4RdPnLz3jSSgGF+E7s/A3SKAIMfEDx40YW5crOdOF8OqwasgsJUnPssaWfCLv6iem2RYz4im2J7r
Szg0hnvwTmTpDOvOTfQ80PIlpkBvFo0QBzNQd8I/5G0WYW6locqpRXreMsdPA32l2bwGp3gHILCZ
0SjnzaLQbLAb/7u+zqu2TREuXZAAhHmOOEKO2r9iW4Ouui9iAdKtGeFLxIYw62Ahz4KO0BODiOSc
/9w6RZWbwz3p8sTfYzjwMNUNIKmfrbGL/NWitalA8jRVtGmqwJWoP4yXQWHmEx2+voah2YwRE3gN
jlbOPLDAv+Rn2dTVMV9oEYCWpu0bbKP4tZI7jtsZgTwquoglSzAo5U0v2vlcQmS6btS5BLwZ+RBC
06lcNCrEXg6Baw4Nhy1W9gAnJzXnBsDgkEtjhXIlRfssba7QZFu8PXJUSdwMeEXV8fnJxbKGqr2y
Eak4MeRBzUX+FKAFyVzsW0zgUyidLSeRsOIV53Uo9aJD/I2bHlXjprCq9WZ+y/cG0Fjd5IQ2uuQn
0cGN00K7VY8lnnJeb/vWh8qqihCFrAR3hSq5/4dfDhIGASdSeWMf/VUeKLjK4dSdOGLTIcTydRVN
DMMtPmCVPyqbV0cuLwTMqJRNgv+U1yeJi3oqKU8EbnSzn2nJgF1dfN4kY7XURlS+ty4c2sNqohn/
twHUW3XqGgYogMlwF+qZwsMZb/2Mv53znhX5wbsgziOu/dIt6O64xmjhy7QFuA8Uo29ApHRFqCW4
6yec1PW3aWFXv4Ifhm1DDZUjw3Lv+X0xJoPk/OX8WzDJOMvswAXcVsUnYt3b60g5mek0zqSTALxb
TgvUvz4ltOQypGrnnWSGIYYLzaYOHt+SHJv4T/AMsNCfRuMfk/hKtILqqIKRqrs7vnee5fgOVHRV
3WCGSsKYQjnhJajqBl60MSeFw3J8HPSmUHLrLhIAWKtzbmz7PsTyjZ7OezAsyoP1hbD3UfdNDvDK
iwSQP1vLhWqTzb2oJCuiONIn5eWlC4IkNmaabudykhsEMnrNZ+RhJ1TCfzHG2BtiBCmzn+3He28x
6qbhWZOIKw3V0rR/hXQB71hzvDgj9tBBIij2tPd7AAz35P52Ym50rwWZRW5Rx+SqnmGyrPEZub6L
y/I7N8HOX0Ecf5ZgrizTO4QYNJAQm3b0F3wJ27Rtmcrw9f3aeFKe/FfJMlu7DhFVju4zDYFS1KgF
T+polqwOCvzZwHJI4jXbWu0PkIGB8/jjebIOcb0RmVxSzsKGuh9XRKSRwxFhEuXDkFk+S3iIlykl
U5u6okrFs9QaU8DaVh050QMQxL8IQY5PeBc4cewB6t3Cax90u6emx1MVe4lyGTdCq6PQcZpwU1wz
6PFyMQhJD4Lra7bmqfOQZstOw8woscDjQQFMki8EMDy+HVVBuXc8YAjgBpdjmImJjv7PrJsjLtZd
luz7xTJ1jFGdMvOZHX+dj+pUOJSbfwTHzgJ2sYHyxZYYuAjpFVRl7ZtLwCtqzznXzKqLQFkaQaIg
rvtSIBB81l1/yqz9Keyx32jlgcI30D/4kDT4HWmnX6Bvm+rzKAQobO4qf1IjERZicXmy+9HHRPRE
T8fzVwJwltIb2Y3qKQie1K+RB0kfv8mJ7xOUHc7zaWRoXyeQHNu/C1l60T414lgNrVHwK+AMA1gQ
9Ijlct321UC7aBuUhfweqYwuyrptScA24NAAnqoLM0fcRfTzfvS2zP0Ju6JwvDsSCsEMBNz/xBAJ
ubSo+WcstzgxAA9UV4O30Se2GlQ8zzTh/BPlVj5IWOixCaEsrmexNcIFJmTi+yBlXfTo4bk7ByuN
vA+vCyeweFnf4sZm9dip+AK40KptiKBcD4TxQrorbcEDRgFRdj3f0PrlpgEgv5sblyX7ELMM3U8a
TiLHQuvuljTjnx2pzJpigTF3B0tnkasALBSboLcsldqo6Q83F44/ZgEKTD4Y7z/x3n53ZFFvvcNi
k1WbiZLnpvioZyaRfu1zoaeWEPeW2ZKTZa1egm0fQ71Mnw4bVAlKw1hGkJK3HNpoTeshKSnoivmt
EGUnwFCRaxxsmDfKBQAKCdXf11weAPg99kH/jkBTWsiX6OHd74QNQwcgD/duYS6Ctv5alzKzsgC9
iGuhCTo9o/B4D4M/ANgYfR9CeGQPTvCiRJ/sgrjOV8qHCIRws4C/2CqWJjs8NMUVzCVK2cmGHyC3
insLchkK9qlDzfXc1c5T65VIJJEDoQiicOHJ+XOca4EWWLNXjOQ3dQ8VeC+CVkXQ7dXcnYwOLlFa
LxV7Cu2KWq/LYWe1I7DpleL3fz0kWqQ0rAmpyQHJwsvWjEjBbPe+LITLzdOzjCziMJXDWIJ6VTj1
hBJDniM8LlCAKt1hgG++jzWIoOhHapwBuHsV2mEgR90S+0HS7fkpSkgYLFXCnm1on1GQpV3r+JbB
5mWtPd7LBid6dkiS8Zu3aYqcpxLcRlLmsi5MoRh8ceci/iFCu/KOegT8Re09YzkGVKPa3o0u+r9X
I7KpcOin8nAQTClTeeizk1khFS5wSdtYce6DN5i8npmgIQcUvjALaNA1RIoZHJDOdW5Z6bWW5VkN
IqwPperI6QXwRaZ2Z9f8xhUVT6ZnhxgsKCFfmiL+/DafsORGLXvogPK6+T6ECmJ6TAGw78LTukn9
e9RqFkaAqKA4sbYo89DG1awWOOVGWwEGlmM0PHTZGG/kzyERq2RE5oraRqjNCfrxhbvI40++YStZ
EustPJKOezpxJXCCV+HG+9xdzqcswaGjzBom
`protect end_protected
